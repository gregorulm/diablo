MPQ    r�5    h�  h                                                                                 �%P=�T ��W�����G4h�������԰;�Z8oY��m�VtK/����%��?oy�
�6�Ԡ.v��i J~����8^��l�i_#{�?e�%C@��S�=���9 ���tVF����\��vDXI��5e�v��*A��ϰ�.T�b�=1P��-��E�`��Q��h*}�>j�8�����!���樟��|!��e�N��q�ِ�����c}�Q%�IT<�k�rS>lΖ��g_�D�P�c��P��Ew|-5�̴�G)ni�tȠ-�0�����"��G^t;:Iy�f�*�ƋVQ���}`pd[E��䝲qe�w��{
u�� $P~�ÿ�&,������w�	�L?^;E���LI��J�.7p7�*Ϝ(@�$I��C�֗��U!_dO�A��I=i5R��~��a���;��P�hN�#7{�,Mde��l��S�.N8���M���+��俎W��>�6����]����&�M����1M�8�:H���-�	�����H���Ab�Am���q�aq�r�*qʼģ�BV��AI`��^N���#����B^�bg�S�S
���=��`m� �{0�Z9�Ǘ9��e:ӄx�\���62���\�jGU���q��ɽp��040�5�z
M{� ��Gφ��\�ᶱNtz����C/�j��=`��HNW]���梅��t�Q���,�M�5�`���\��H�PL��W�!�Ë���
`R{�X��O�$��>���L2�Ș��x��)P���/�8��)Y��v�Gm� �\��Ò�%�*�81�&4u���詁аpy�$���`_n�� *��(Y@�!��:�(�!����$�	�Sk���ޑ��[We�4}#|�Zk	"��YZE-��corh� ���Nu��4�S{|I�Y�$KQ��sY�Fo�>u"1�y���`���8i%�����[x��g����]"=�q�ߑW02�Rnx�Md0;���sv$���^���G���bSSˤ1���)m��K̽'=�����{	�֧/"_l�AZ�iԉ�qP��?�Gh��������cl
��F�~�t�5��vK����7������Ƀ+��	gj�7#Gڒ�,ò���+�A=j7?����a�|(�� ��u�����p���6��` �?�ͤ;��[W#z0}�x뜘pc����z�6�Sl��tP��
���lt�'.����Wp# ������A_ �j��5�,M�O��blgjr�´��6p"��U�
'��b�]�N�p�/SlM��3��Hx	��r�T�G���b�XL��z�/�y��1��(�\)&�q0��sG�%��;��k�?����,R��ۺ�}�E��ӝ�\5�pH@�WDf&B���k�E&u��HT��W~�:q�i_ H��տK.ˡ}��4԰\�N�����u$f4Q�j�����jUd��s���;kG� �=lU닿
3iJa<1���V���"x�A+��,�h�m��y�N�3��O�2w�nՏ��M/#G��4�B� ~=�2-��wK�P���ğ���/�(�K�5c���AWȔ9�,h[%u�.�"��ڜ�@��{1o���Q?T���$`J��O]����3�%[]�y�v��&V�&�f#&��[�z�4x�г�l�J��;k�ml���)3����4q����Q��G��u)�K��ʆ8M0W'�B"��E���V��(��#bk.����k
����3E��!ƨ?__�QjBM�t���K���d��k��d ɾg1�S�!�7�(zX��� 6N]ڥ��ʺ�w߿�ʵċ�~���XP���U�m�����p|`���6 �ɭҩ���=oh��_Kr5���nc?��Z�D<�ٝp�l@�7�jX ׎n5짭��O�3R�O�m�`��C�[�N�W�ȩ�E��QXokXTw�\�(���ĝ�ӹ�� �!���*J�vy�v9��ώk�"�FD`����*����4�d�Z5'e�Pz�>�=~e�N����u��cj(�00�,��ƛ"��y�jq�����<f%ߪ"���Q�͟�},#��É�}��<d���⇂&�l�q]�1��3�R��t�"��=;&`[<��l��������.�s$%QL�PI{�k���>S�e��)����*A:�aD7���p�B�_�����5
�O�
��*M��f�Vð3�t�kJf�Qۧ�rNx��?yK.F�)���![*Cy��r<������㟃��W��9�2���IH�s7��ϕ��UnYL��2Q�L>���R��J�C0ߋ��p��.���"�#@���a��B�y\�2���X��pٽ�Xw��/<��h�/�o A�V,\mG���ُڇ�6���Bv|��>���ǁ�}�l��5�aJ��Y�[�26Y�2V��F�~��,��>����O�ƙx��2P%|w_���q'�ɪ�E��ٽM�I_�R���B�I���r~�wo����ULf/h�8�d�s�{�ⱏ�ʩ*�^�9i��Z�qZ�盉���'H�D������T��s����ofE�{��927��d�+��u2���&�H2-��@��h<��w��|W���Ё*�"�4�v��(2ܮ:a)�u��s{ ����,S��!�җ'�i�mM�r�2Hb>�#�'��M�kŲУe!Ƴ�n5�N����aa�[Y2�	{77�N'�
�+9]�ם���wvqi#��x�|�oӄ�����E�3�&: �vDo%��5Cx~{{%�%ݎ7T�Q2�쬟�[�F9��1B�_SB��&t%]�������T�"g�e�I6�_��2-X߲�G��S�Rm��ʒ�
�;Ni���Y��3�S;� �_��=NG�9(3SdS�*	Z>�+U�9��hE�>���ܸ��?)��!$�V�z0J��Ww�}��";�����&���!r���a�+Y���8�1!(��j#��u����y��p2;�W�v�o�>�(��_�>b�s����ξT����$<@U]l�ͬQ9o 3����X��=c�������9;�eWJx-Cjt�˩��S��d}\���&ے�p��Zj���|�7��^�t�o����dN���7.�����-�h�X�%G'�[�����G��0Y���۬b=�P1LmLx��H����q�њ˳����[��B��q���|d�&f.���t<ֶ为�r��T���}f�V�rGƮLJ�]��4{n�Q�����,>(=��$�~ꓪgq��i	u����9^�G2II<x��^+&���%���]f��E���}�'��U�zP���Jzކ�ߤ5��%SQ�j� }��� Qs��� "kGI;)�AI�sc+�b6���`�!�ye�EZ�w���Y�<����h�]LW�!����-�����3�"-�Q^���X+<��cfb���Z/�l���$�C�_�!����ҵ;n�����������4�Ol!>1��{ĝY�@s��/����gPX�����N��6K w�x2@/-�;�,��n���VR��K� ������������­`�<�mї�o+�'>��	����E�w��bYe:b�+6ap�x�G��3�xz��)u1
t�u�b��ʋ�jE���i�Y3�8\���U�py�z��b�(�G*�O���ф�t�'���I�ߥ��=����DXW�pڪ����ɦ���d�,Q��g�qM�%`�\���1��롘��fL�&��RJ�����1���Ź��L����s�������yt��>/5y���t�� m�;�7Y����'%@��8,�	4��6������`y ҝ�ɽ�n��*���Y;�>�?����G��$m�.sB���u�ƻe��n~��Z&2{���E���cJ%w�;(��h��pQE���{7��Y�O)Qp��s4{�F���c�1��e�V4���
i@���4�wx��hg�@m�m	�=ː���U�2p&n���Ȉ�;eMZs�S�ՙu"�1F�U�S�Z1��')��ZK�3x�kژ,�	{��u�'_�KRAuq���P��?�'�Nڢ�}8�c��
�7�F S1��@�i�K/�i��%"��;�$.�+���	��haA#":��M���)��&"c�Q7ѿ��e߬�$�(��;^>u7ѓ��QH��6��(��"�"`��#������k���W5( �nڮ�����k��+�p��1���rW�y�����S����, jv��pL�M(���֤�gi�?�}a�Q�U�WG���ݣ�B�Y]\(p�<,l�����=�c�`���/I'�x�bc����R�/Q����<�C�O\�e�L=Ǯ�O%!�ם�?����������}��� fr�؃�5���H;	�D�S����U�`��<��jx~��Z:o�iZY�A0S���~�4�Z��7�&�����!�+u(���5jYoŦ�}jU�:�scB�v�R�) �3�ŋ�z��ie��a�V�]h�V�|r�>�A&�߇��(��y���R/�*�wB��*	oM*���-9UB�g�~X��-/9�K�
|��7�f���*ߒ����cL�Ar:9_�[ څ.�"�u���;��f�oR��QZ����{`%��O�̭;��%V����]U!�Vo�Z�#W�[ʐ���UmЮ�̥Q�;&�V��j03�W��Uw�68Y��Ge�-�G��)�iK����8(A:'�ng�T����}���ځ��3�.�����6��[�3�R�@@�:Qi���������4�^y�������ɹ�sg��x���<�%��<�3���[�r]u�L��Bw:G��p7:�Hx�NffӾۼ>��m� b�� w|�]R����ȇp��ڻ�װ�àr�I�����?������mٸ�l�0w�EkT����5�!,�	��O�;��
���{h����X�)D��#uE:/�Xj�T�/���2���:��N�e����:-4J���y���bT��I:±=/�D���`>y�?��&҅UZQ'�P�z�q��X�:e6y���&���2�c0�m,�!���;y*�Cq����f`�"�3�Q�����.���)�ʟ����������B�]��}���RV��=^=��[Y���M�S6��	�dVs��Qg��I�ݼkyH�>�`��r��)�LK�W�>�OJa_��2O�p�X�_Cw3�H,5���e:[*��f*��>B|3�5�k�B���>��m%��F��K���)�p!��XCT���Y��c��jҟ�j�WW 9�֮�j�^H��-7��̕��i�N�D?��0�>l[����%��Ck�����)�5�}��#���ۖ����7���1�\+Iٸ�SwmBQ/���ͪ���� go'm����]��+�ڃRM���e��㷊�Y;}6R���� �c�Mq;ѭ���!6��G8�]�/�ԃO�`3D��Mv2|�HV�^����E;k�H,z_a9�M�:� Z���ӻR3��N�RU�+h�2rd���6V����^��7r��2���bZfy����j'�9J߬���i�TB�`Щ�i���������%7�X�yC�-��u��Ɠ�O*�L��-�]�@�~<R�8�`�/�z����v�v�@�2w�a$�G�I�ȷ.��=,��˨��B�X�����mHΜC�b����B�:M]�qk�x/�R�Xa\�i��A���2a|Y�&�{��NI�r
�?�9X:���0ޏ���q��-�%��W0o�uIcE����Z:�Æv_bV%�CSE�{`I��)!��LOG�\([��9�J�1��S�&��2�K������gJ8�IQ�i�a�|X��G����tJhlӿ%���R�N��e�ԧN#Sviǵ�C.�8���nv<3M�n�C	�A�+0(��7ͺ�=k����n�A?�O�!&�\���0%���P�}o��6��<�z��&�l՜,��*7+��V��\��, ��(�XM��a��{�K�Y֒xc�
���#x�_5(�����E�I���9�_6ZU��*ͧƺo[G�°;���i�lz�˛sB�@�e��x(�"tTj�~���)�I��m��/_jC4<�wŧ7 *�/z���k1d��3�N��5�-��D�S�G�,-��ŧ�"���D�p�n���'�=���P,�kLӵ�yܙE��LAس�Z���qB�h�qӁy�g3��ک��<Q����-���"_	}�o���r�(O�gc+]$�|{I���,�[�(8֐$Z���e��q�di����8�^$[���7I7E繗˟��x�ɧ�ِ 	�5�� �U����gJ������5��S,�Z�[���<$ Lր��k�(�IV�^A�wc�6� �;b!�����G�w]��Y��\�x��h���W短�kH�-����&L�"��|^	:���+��c���Ň��g�s�U�CA+!�!;II�X{\�v	��A)���O'[w1�k���>@N�/�fs��iS�m!��	X6f|����
��;��R��`'��{������_�[���gY��b[���ђ��o��'��J	ؼ��`��.�"�e�)U�&�4�.F�3�����:"�E�E?�u��׈�P��Ŋ��<�~�t�ɳg���	뾫O!z@hB�ytG�G��ґp��w�tp~`�og��k:=���`~WĪe��7�d���޳";뢼�M���`뜿\t]���۩9Yǡ���A��a�R�(��G,��>״2V�	5�L(�1�N�d����_�K���/rQI���H���Pm�M�+���%�s8'��4+ ��X.h���y{�&��:tn��**��Y6�������L��.�T$���	����/Q�e��<ٖPZ�z8�)�>E#Hc%���vV���Sk���j�{��YۚQ�O=s�`F�#U���1�A�ϱ'@��wi[���ɿx�"�g"����S=���Gt�2+ n���C��;@!�s좼�4���;��ՓS���1���)c�$K��.���3ΰ	v�����,_�KA�hI��KP��?H�������z���7
}��F;5��j��c>~Kjd��m��
T����+>�	�����#�����ز�v��!X���7�`����W�(j�v�ku�r��R��=Wt��G��eT͚(���#�2셮<�f�H�Vk[�ޭ�h��jӚ��n�f�!�]UI��	YW&��N��Ϳ�7x� E�T���M���gČ�8.t�l��.������}��]�!�p�i�l5ƥ۩�C�~�?��y�
��L5�b�c��J�/]H;秭��^.\���'jX��J%�`+����?S������J}����=��W�5H�H6�`D�j�kͣ�{&���Oƫ��	~:�:��iU����P�����y4������/�S���VuLd�wgj~+��c�UZ��s>ʫ��G�� ��5��5di��qa2�݃8�V0|�X%�A!���⨞���y���5���w}����Z�M%J�]B��~s,@-��*K���W���f��%/��7�c bA��/9ڷc[�^T..C���T�Vӷ1��oa�Qu.D��` �vO�29��8�%Q�J�/r/V0�Ɣ#�1�[�׽jSJЩ�i� "�;�j��r�� C3�� 4��Ѡ;��Ô���G?t�)����8r�'1�`������u�� ��%}.���a��6�W3�[���~��5cϤ�Ö��2�A̯9 #�AX��;Qɴ�]g�Y�y�W����&����]�����"w����+��2��ɓ(ә��y%�mT�Ԁɓ9|0c�;���\��S%��^I�WFJrk4���ʵ?N����mL���Sl6��� ���k�59w����OTd�����ޖ:�9�a�"�>��E���Xe�_T-�UÞ���ҙ�Lg���ʎu��JD##y��l�҈��ݱX�DV���;r"�z�Uj���P��'�{zgFжs6�e���woǻ��^e`0	B,L~|��P�yE�q�Q���0%f�I�"%��Q����3Y�V˴����~'��^:����A��]�����G�RN��X3�=1�s[�8r�����x���'s�s��NQ���Iq��kT�>�F��C�)���ǲ���waz�����ap���_~hf��#�5 �����*æfE����3uk�>�͇�r�h�ܡ̚K�i�)�I�!Q��C/��`������,�9lLWM9����H��7罕,tdSͯ�k�}��>:h�H�P ��C����(�R�$(���O�#�S�v�8���w�<0=��Z�ٳ�
w���/|���R0�%� �:����m}�G��Kv��q��>��76I��U�m�y�}�W��Z������F3�h�%�(�����ƂLׂ������O_�����h�g|mR4�9õ�?3SE�FC�C{�_u�/����;�����t�-��V�U��h�LOd^0������Z� ����f���MHZ+I��S'��O�gׁ�p6T�|�Є7 ��0�7����y�7l]ފ��H�Xu(T��4^ˇ(_-;�@��O<�i9��K�*WJ� �ϣ�<v&̑2t�a�����?��k��],�Ҩ�/#��3n��Q�mC��ks�b��{�]C�Mط�k{^���$�$/d�����MFa���Y(��{�8N�_�
+s�9S��S���s�
q��u�;�2D�oI�:��E�C6�qix:��Zvz֥%��EC.,�{�e��*��G�Z�b8�[�M�9�b18E�S���&��K���҄�
Шg+�Il7��-xX�uG����T�c?�������N���O��5�S�Lⵕ���3j,��Ӱ3�U���D	Pe+�\�W%ɺt����jh��p�?��'!A��Lt30 !��I�}
/u��iU��U|�q�&�bU����I+�⥍n�۠'�-�8��j��S�o��&:H�͇$�����B&_�1xA���J��=as���PhU��͢[�o�{=�k��� ������v][�eeOЧx#�vt�jJ�d�|������.��H��K_�j�k��r��7_�5��O%��HdD"=����pT�-$�C�N��G��^�m&�=��t�I�~�"n�=8��P'�fL.�3��d��/�����s����C�B�q�76s�ǜ3+��R<̹J�p��N��BH}� crw*����]�5{$���X�.)�z(3��$�!;� a�q�0�i������^_��h��I22��$q�V Ё�I\�U��J 4���]�NU��a�B�J����ϳ�5�6�S�z��m�!�� GY!�C�Ck�V�Iq��A?�Fcᮓ6����5�!�����T�wNaY���aqh�ÔW">���-�ȓρ��"�,^$��w�j+�Hcܔ��"���bi�ڸwC��S!(Y���;$�B�/t�E������fO�t1���ē��@)%/&�����N�������<C6����n���;*���+r7�����y�Iv�m��ƨ����o��88j�rb�э��o�Z'���	�[�;������epS�!��i\��U��nx��4�*�u<&%����� �t����яG��.�������E�z�%��CG��J��-���_t��%�v���m7=1������Wn�M� ���R�J�vX��������MU�(`�\�C�ˁ�H�TB롎��dĖ��%RL'ہ�%��Q�oo˹$	�L�6��).�)���,���%;/͍�ZP ��~!m�`6����CJ%vH8"`�4��'����!O7y��[��FnZ��*���Y1����үY*_�I!�$cSW���8�?H:���e���4T:Z��Y�Dz�E��!c �䛱������f��ES�{���Y��Qf�sꖖF }>FD1�Ւ�;w�K��ivk1�*�3x�k�g]�yţ�@=�.�ߢ�r2��n�/W�1";�s'o����e �?SO)q1��)�2ZK]:�6�Ώ�	q�֧+�2_Ek�A���}�Pr`�?�w❄���W�A�
8mJFV7���*[>3JK��ʭ5���޼��+�F�	���^b�#�Y��Ý`�_yk���R?7G!]��z�һ�(EY}��um�H��s�����⑓�(��O8�h��#+䁅I8�a���������`��D��Z��ΡA����E����W��Q�J�,f��4<  ����M^���̈�gN{��������M6mÛ����x�]�;�pŶRl����d���e��ur���l���b��ґ�b/�_��b���yh�\������$�y%WP7��[?��K�]���,*�}�x���5.�NJ/5�?�H1E�Dw��&�U��V���a�x�~u�R:BڞiP+_�@ο|�СΔa4�7i��K��j�U�W˙u��E;9jϬ5��i�Uխs4����<�� �
uf���עi���a����mVk���+A�I�=�	��c|y+�����D�w��*�`�M ���㡵BI�>~��-%nVKdޭ����B�� �;�\��c�z`A�~�9U�c[�S.i�����w��{�o�F�Q�˿�F�`�9NO~��q��%L��Ǌ�{���VK_�}Q�#�,�[@b�qФ���[-;�f�����a3a�o�?�l)6��_���vG��p)�
���8��'l'���\�+/�9G��T7,.E�������_3�Ҍ�vݠ�0���b^�~3��N鼃��j�|���5ɯ��gB��4}rʙ��!��w���}�]��pջ��w�7��|�<j�D��t�����m����&�|q"��gy��QV�|�Z��2���Gr?<��(�?��W�u6����l�׺����?�5������O��
��K5ޱ�Ս��v����yuEp�^X`�T����Y��+�)�DƔ��:����cJ�n�y�S`q�Ͽ�sQ�Dш3�ƛ����t��KN�'v��z";ﶎ��e,k�RnX�G����,0o�,�rכSЪy`��q���\�Hf�.9"�,VQ�� �*���c� DX��5�9��3��=�]����D��R�㦎s�z=���[�8,�������U��./sU�Q���I�4�k/~�>Mb���)�.����k�)a� ��(<-pd��_�y-�~\f5�El��n*~�f`�L4��3PJk�Z��"f,�c3����KK_+�)�BX!���C
�s:��ҙ���ğ���W͙�92��`n�H�]r7G����_ ȯ��A8�M>U����=ۡ�C�6?�þ���l�3��#q��/0����1b�wx}���#ٮ~w#g�/7���}��� ҒH��?m]���Y��>S��#�RƋ�[���mp��׮}l}��3H�r�E��J�كGѣ�[��qGƽ�
���X�ʫOO����A��"�|�{>��z��EqB̽>�_���àv�V�A��ob�:��շU:,h���d��Ӭ��� �������
��!Z��S�'YbU�"<�8�6T8���_��� �]�5���I�7�,������cįu�Y���9����C-֌6@�0�<dz���ET���6X�ŵ�vaw�2��Jae�������'���,��Ũ��s�����:ϐm>��� boE�x�MS�UkVd���H���_�=_�-�a�y�Y�	�{��)N�+<
�Ƹ9N��׮]�.m�q�������o��3ͫ�2E�����:v:Q�v�j]%��C	3r{����_T��B���4[B��9')�1���S�I�&%���Tc����e��g�=UI��v�W�XpiGB�D�$Tb^2��)G;nN�X&��x��=/S�OQ�0���.(i�$Q�3�~��-	˨'+�m���39��V����$=?Z�!\.���0�~�c�}�oD�����(�,P�&�x�Ւ���+
��	�C�"��������(����x�����@���,�_�Z��y�8��?��Nx��ՊjU.�E͝2o���&�|�c�b���Qg�0�Ke�:xcgt
�J�4���c��4��#b����jyò�m;�7�T��E���(d�r���Wϫ�:-�P�IG8��(���X�h�:�c�$�a�]��=��P"�]L���yp��J+�B��NbM���B�y�qɹ����W��
��<G뿸Kw���i(XF�}�j�gv�r2L����M]��{����� ��(.:$����q�t8izk����(^�_v�I-?��o��8+���׮]�֬
oPE��	yU�������JDb��͏5�nS�ʋ�]�{y B�}���4kE��I��A�C�c�f�60G�SP�!�cu�V��w�&VY����nU�hi&�W]�굡3�-}���ܮ"^�_^?�F��+ͪKc^�Ž���]m��5<�C�� !9��|;��w�@ʬ�7���EL�O�.61�u�w @|/S��R[�I��#�h�AT6�����0+��;e���ƣ���%�����1)��M��Qe�J���s-���)ш�No<Ƶ'o�	�?����E�Q�e	��fròҩ:��޽��ۺDg�5�uטJ���r�{u��-�Ѫ�ɩ���_f�!\zv�{G;���H���"��tf���Q��V��=�d���Wɢw��A�m�X��9V��#����M�C�`�ʛ\*J�<�z�oKW�	{��W��'R�E��zB*E�*�$�?�7L�����d>���b����/(��8���]zm#���.��~a�%=�8�[4�У��<yq�<�Z�In�(Q*`^mY,3��PDN�(Q�d��$ޫ���J��z��e��e��l�1�ZWlߖ_�Eo,c��C����9:a�R�[�{h�oY��Q��s�T\F[����11ȉS�gnN��Vi�����x��Ng�m�>�e=��Y��	2�9 n��9��;�(�sb���jy#謯g�f�TS
��1�J�)Y�K8��))��iq�	l�y��@8_ �zAƶI�u�UPM��?�ޝ`+��ѷt �
�7�FqY:�`�jHFK�I����� �ʼ5�+��U	�ޒ�)#����X=�����$��RF7K�$�M��( ą�P#u�4���D�L���͐���C�#f������\��bDf������`���5N�������y�˗�W�<�2��G��-6 �Y��!��M��=��**gz/麮'���@`��]M�v��j]-u<p�#�l뾛������������.&���b4+ڑ��/�!�ӎɔ��\>��#��_��%�_��۷�?	_R�Is�G��}�*��MӉ]�5~�MH,�Dқ��l���y����SS}~���:ݿ�iK�	R�˿7}���Ϯ4�]�ȹ�������u�����j����ZUP��s�,N�'%N�u� �9�����i���a(C҃�S�V����RfA�ߘ�T�Y�.yF��p����Kw�3���]Mw=�>fB��~��m-�8K?�^��Yx�7?��/z��5�c}��A�Pk9��[�ȁ.���F{���׷�5_o�L�Q�����I`��uOI����%G٨��=�s�Vf���s#�G}[{�`����П�W̶"@;W�)�x���3<I��y��H��H�>@�G���)�%��8�3'��o�%���z�$���4�i�.+���W|���731jh�\�+篤��9����n�7[}�m�޷4Ś��bɪѥg����_Z�	 �D����+X]F8�ն�wK��ʡO�fߵ�N��O�d�u9m��ဿ��|�4E�"���gu���\��j�ͬ�r�iơ��x?%�06�	�sl,۾��c��z�5o����)�O
�;�*���y�/���=#�N�E��X[��T���τ�F]���_�l4��y�Jzگy�2�s/ �zw`���DLm���9���q�J+�F��'Ѭ'z�O�n3e�L��-�ٻ��E��p0��^,�2�phy{ q�&>�7�|f4�"[٣Q���i�� 7�Ɛt�~�H�n�-��(i]������UR��ꎎ�4='��[�X6�X�;�$^.�+�)īsR	Q�?�Ig��k
I>?sI�C�n)��3�hl7&S_a�c����p?Z�_�����'5��X�v��*94�f{�����3+80k6�qͽ)�^j��WټK=)�[h!G5�C��uϔ�4�%�ǟ��2W��9M�!���&Hr��7�k|�b��Z�>�U$��>p��>:��C���^Ä�8�^0#,9!J
��.�M��|���-%٩h�w~)�/�򼓤d� �
�iJm�7!�Ň��<,Mڴ��mv���Lj�H�=
V*}���,�����Enٞ�����?U��>҂.A��oOvd�r鞨J|c�t���;|E^��9ys_+L\�~ں�qM�v���>���t�U��0h��d��gDٱ�|��v5˥�]�F��Z7�։齙'�&[��V��S޾T��o�:]�[{�m�ܕ�9�7"J�P�b�~��u�r��^V���\-qTg@~�&<c~���SP�`q�������v�BK2H��a���Z�M�_~G���,����4�	����l[m9a!4�b*�䞓	tM�D�k1���*x2�Z������3�a�WY�{��N�/
a:	9I��	$Q����qՇ)k�/��o�� �F��EŇ��',T:��v�}%��C�YO{�t�����=f��Q�[�|�9B�A1.*�S��&`�,�	��B}��>�g{p�I�+y�ҨsXK��G}����s�YE�6���+vN��2�E�q�e-S's�˃�)���3?���Z�	F%+�@@��a�����Ȝ����?k�!wy8�B�0���C��}@�+��1��M`��8&�E����aE}+EK`��_�]$��#���p�C��e�>����C#���z�6�_F����S	H��<)����`U�2͘�'olD����;�6Z��ݩ^�,��k�e��ex�te�k�ھ���E���Y&��6k���j;��h��7�`[��8s�d:��m'��*�-Z3ɥD�)G����G�sg���^?���ۘZ�=nYpP�PL�Y�4�u�eβ���F�)8��GF[BU2�qą��`����%OB<�<a�&���d�in}�v��r퍂��n�]�N{��q����_�()��$kD���yq�>i�RT�\]X^�9�oRI(l��ʜ��̏��5VR��.%��ݓn;U�������J�D���5}�S��J����WK� =�����ek I��A5Jc�>6k��!��2���w��Y���hyhD��W��7�<ټ-xZ��7UW"^Z��m?�+���cRG��X���X��ԐߐCrڑ!T�V}�k;�s\	���G���^���OXȻ1�ĉkS@���/����A�D��~���:fI6�Pm�dp��(;��ӝa���|���/ ���������D%�\�BĢ��Cу9�o�1'*"�	)̜1�#�ʊ�#�e�@w����=I�d F0��d<�ەt�`�ur+H���"��n�m~���o�$J��w:L�\��z��,�G�XF��K�=>t�A��,�tߑ��=gm1��s�W$�A��kJ���l;T��Te�SAJM�`�d\�p����p��t��_�������R�����+�{��Hb�Z%L�E�������0`��׿(/�f���?ܾ�\[m|���`�ùμ%�Q�8��4<�������W�y��ɛ5q|nР�*���Y'���
��E����$Y$����o��.O� ��e�*��..Zɖz��E�2#c�0�'����q�\����2{#hY,<�Q\�s�2�F���|�v1�]0���Ň�S�i�w<� v�x]]�g�W����=�L\�X�_2\�&n���Z�;�\�s�PP���+��q�SŲ1	��)��	K��d���s	gܘ��>_�
;A���ҬP(T>?��흺�3����Y
�"RF�����&�|rKu��>���Tr���+o	�(T�c#��Y�94n���+�����7������l(�N�'7�u����яNxm���!��@�)�#��i�&�W��g)!�/��ұ�ۇ&�/q�l�.��Ǝ�W7��ӳ�b����| ����\�vM������g�07�iT���4�C���Q�W�.}�]��:p��ilF���\Y�ϣ�kwӛF��,�b��y���/n�����ɯ|�\��ظ�xǚ�s%��w��ڣ?dᘒ���b�}��+���*�Đ�5U�H'�D-I���w��?�J\�.6_~�:x�riF}���I��`��+4��^��G(��D���hu�w��!�jEj6���Uˠ:s�e�by_rQ� ������f�li�Ëa��>��7�V�9�)��A�=��T��M�ya��xш�B�w.�Ֆ�M\qB��~��P-#RK2 ��`��[���T���c8��A�B�9K�g[l��.�c���/�g��Bo>r�Q�e�w'�`�9�O�ty���1%B��@�_A$+V�φs�E#m��[�)ӽ;�К���S�;�"�+��3/��Y¢�s���ˏ���Gph�)3"i�qb8�ħ'�_�����uYV��3��ʺ�.F7���(1����3l!�����&Y*��l����)�R��T�����k�ɥg����;�h.�����{��G��]��ձ��w���\B]���:�w�*�*N�m%�|����|'g��T��4�\�r|*ㄶ��?r<�(��D$?_�6��'A�$��l������׵�)5
8����Oe�[��R����%��zū�{���GE��XV/�T>={���ǡaSO�:t�G�p�&~cJf�y�1���5!ȱ��ED�q������+��;A��A�[',�Mz��ٶ�:e"���J����/*-0�x�,]����/*y���q
�n���fLY�"���Q�m��Dɚ��K.�6hq�ws��ه����s`�]��Y���RBor��z�=�؋[�������� �!��y�s˲|Qӷ�I�nk�3�>z����3)��y��L5�>a�ƺ���p��_/�w��-5�=a�ѧ*��,f�,�*��3y�kq���XH�Y�ܲ�K��)��!C�u9�6=��/��2&�J0vWC�v9h���V��HMkw7��I��@U�1������>�����+CWƥ�������#�ېe6���0�����h��ȩ�٤�w�@/��{�q���z ���S��mN2R���҇�9��ouc�F��Q ��#�DE�}�(Ґ�E�($l� ��ٹ�љ��-��3�-����S	Opw����N�|�.���-����E����4(�_�ڒ�94��� ��!�����:4mUSg�h�Zdo���")�����u�ˀӡ��L�Z��щ��'aߘƼ�nE�T.����#��P}���I7}+0��
ƙHVu�d�a��8i�-<P@y�,<����L�8�{�݁��ͣ{uv�-&2��a�)��^��˙+�,��o�h�d�D���p*m4�|�Qb�\_��BMI�jk�K�>+ �>U!<o��~Z�a�U_Y�l�{~��N5$�
�͑9D���d
M���(q�p�旛�÷o�����bE�Y��=:��.v��%U�C��{L�ݕ��8}�s�[�D�9]�}1��hS��&��R�ޢ�����g6�qI��#�M�sX&��G��r�Z�ZTx뿑.��	/N�b����z�{Sb�+�f.�$w�ګN3�/	�ڸ	��+�3Z��u�E�"��eb���8?�^�!�䑴��0��
~�B}�P+���ϗ�/B�-]&�Ո��<��+��ˍ?K�����Ib(D��^����MQ����~u`�vHf�`_�*r��n5�5����K_KUd�@͓ڙo��N���QqխX�h����e �(x�t�H��i��G��T��+b���|j��	�c1)7p	���4�S`@d�s!�~G�!�-�5P�?N�G��4���֎?څ0:��+x�� �=	�1P�?L?�,��簙��W�8��.����{B�
�q�qGU���W��@�<=�.������S��U}�E�vr�����]�{��	��U�($
$�E�Q��q]�ipZ��7Tx^�W9�KI#���%�b���5�(�3���O��.�.�U����S��J�G�� b�5���S�9��GƜ��:� 8�k�T�k���I�B�A��}cr6�6�R��!��̿=�wI8lY2�l�d��hL�W����מ�-sӋϒ�"ԨR^u��`+�&c�P���%�S՛��C-	�!o����;�l�D���l�����O�17p/���@��9/�#S��HA?����ƴ���"6�,o���9vw�;ۿ��f8�wO��a[����#���G�; �(��w�C���~��o��'�|�	D� ��v�]o��c'eA����(����7���|B�p�1��u������1�z�(����ɟ�m�R5����z�r���G�H����G�X��t\��G���0�=���0W���Q���_��\~�s��뎭�M&R`�xh\�n˲�*������9í��M�`R�v��O8���נ價uEzL��Ⱥ��"L�)Z�Ҽ�/����g��|�m�9�~����[�%G��8X�4�}��D9��r�yg�n�n9�*�}�Y"9��	�������$Լ��uz�����훻[e��EL8Z������Ec��R�bO��o� W��V�E{�_�YG�Q�Ius{0�F�Hs��1�Q)�5݇|2�i�-����x8�g�S�tCX=��߳-v2�n�%/�;��ns�ՠ��袣J�;�S��B1$C!)O�K��}��ڟ��	b14�<	D_v��A��j�k-�P��?4��UY��ݙ�*?O
i-F����V�����KVe�ٻ���?ּ�a�+*�&		Y���j#i�>�t/�0AP�p=cu7x#S9>1�C.(���b=�u>���i����6�<2l͆����~Q#ܷ��_��RK��ح��M�����VY���/��R6��#�����W�	�����}�ڄ#* �����M/��Žαg0Re�$�����o��R�,P�i�]cH�p�]�l�7�ە4���r��)�vv�8jbjԱ�}j�/�e��x���68\ؓ]���?%(߫��b?������}�|}����gݠ����5�MH"�D�=�W�đ��~ݻ�	9�~&c�:�PiAVS�G��d{��a4�rk�~�П���(�u��VEoj �,�*<�UF�s������$M< ���w�!��i�za���;RV�n��<A��N΋���?y|׷�χ�q�xwi(|�1�Ma!��.�Bz�~��-�-"K���Cd]�m������m�8c�J4A�TG9�Ml[G�o.;�|���ͷ�
�o��Q�b����$`l�O�7�Bä%=�wǛ�����V��'�#H�[�߹�։oЕ�5�l��;���,v:3�4h �C�=����k��tG+O1)N�Լ��E8ou�',O�[[��p ğJ���,�.a��M����JX3����G���!� �sr�ɨ�*�K�-j��[��-��"Uɠk�gS�5eO!��Ĕ
�6z-���U]|A�լ�^w̱�U�.µ����l�eF�m��π���|��'���O���t��_�̶C�9r�c���?�����P��?4l"B�茩����$5�K���O�ED���� ڍ%	��p�i�*a�EA2EXQ��T��Ê,��|i���%�"�]�a��J�y�P�)��������DB�����f���W�<�D'��SzS٤��&7e���*����kʫa0�-l,�雄�y��{q�{+��f��|"��Q|���HF�B�I�Q*�j}��M�������]���U1R�d>��'=),[^�:��]��Z���7��N�s�3TQ�OdI]�(k�>�>�t�y9�)�q��M��JWa�I�����p���_jm��O��5���,Ӽ*�A,f�����3��k�o�����T8��f�K�0�)3�`!=�C��T뽹�j���t៥��W�?
9�����dH("�7�o��PǠ�]3it>���4Tlg`C�����,��ѴD�#��$�B�$H�~�B�(w�cYPٟ�@w4�/h.�(���� cZ��[m�L[�C���fa�*Nc�6���0��8���}}=����~8��|?����x ��i�h;!�n��d˱�WO���ڭ~���|Y�e����+�uEB���/��_ሉ����|�l�����uU�-Bh��\dʫ���--�1�\��)�[�՞�6gZm1E��g�'jg�SV����gT�f6��^���E+����y7�Z6�ƾ�ƴ��uB�<�si*-�C�@t��<��e����غ�V��v9U2~~�aWH��ܷտ��Ff�,8'�C[�̕��m/c4�t:b�^��OM�Qk�5{�yLh�P}�pJ��9��at�YN!{Y��NpP1
��R9?��׿	�_�eqz�a�S��s�o5��|�~E�K���n�:�S�v���%|�vC��{�TU�0�y�3�����[s,r9xfA1$��Sd4&����&{2�v-6g�56I؟v�ȣX@G�HX���Oˇ����l,N��;"US������"H�5�C3����zZ	<3�+wF��CB��	}�N�5��?�r!�o�8n60lX��nK}v�B��yۗc��]�%&8{�����q+�3��Vˠ;���i�݆�yI��[ү��#ֹr����
��_��%-����挰���T����)U���͎�o"���W:��l���Ӿ���D`�:�e�B�x��t(�P4��j��/۴@��7`�jJ�I�^�_7�������nmxd0$[�YͶ�\�u-�X��:��GI��Y�֩75�������X=�T�P�*L�W���Sp��t��aͳ�C��0B�Aq�}F���ǈN֩[�<�?(��Y'�:��)u}�Qx9�rcqy����]��[{��b�Dp��$(��$!�]���q8�i�>�k�^K�j�¼I&:瀕�B�U�P3�H���g�� ���ɗ�U������Juj�;�c5sl�Ss�ۋ�Ί�J^ 3����n�kvM{IݧnA+�}cMN�6� v�$`1!�mB�g�wq�YM=����1h�gW�-�r�v-nl���("�l^�!Wc\ +^��c�y�Ŏ^k�N9��F�*C�W`!� �sk�;��6@��}s[��뮗VO�[1R�����@�g�/cݍ#o:���4 ����6�(��ZO�Q��;
�(�r��Ŷb�t�>����d�ۨ�$�n�ޔ?�y9oM�'���	_�ݜ'�e84Ĺe��{�E4��6����R���Z���K4nlou��ˈ�����������'����-Ph��^GzG\*���ZGLYB�y���s=t����N���=������W�����I��s�b�ԳN���9oM��`���\;��mͨ��&L�zXÈ𖈍�R�a�����S~_�[�����7L���ȕ���f����/9�[�F���3��mr*R�Y$!�/	�%���8@+4�d������7�y���rnF�*1=�Y�Z�aB�Eῑ��5$Ou��PB�+���6��e�(���Z��Ȗ���E��cl���{�
}XR'=�4�{���Yb�QR�asVNF"���H1�e>�xȔ�71hi�����x�egI���%=����L2�v�n5t��9;�$�s��;�=�M��w$�S;�P1?��)�0jK��)ڷ=�:��	]�K��J_1*�AG���P���?o�I���跅~e
$X�F�,�р��F[K�u��t�F��J��F̶+�]u	$ƪJ�=#Dt��J̲��L�F����73dmT����i�(��?�cuقS�7���>�}�Wu��)z���H#顅��X�M�D����P����J`��P�΍r"�d�g���IW�=w-�
V��f� �]p��aMʽŸ��g��s�������9�v�����f]��p�*ql����P,'�b��a���Q4��s�Qbف�x�/$�k�N�%��_\�6�n*���>%�N��̀�?F�I�Θ~�}yZ��BUg�:W�5O�H=�D����W������[s~a�:�0'i<O�c�ſh���:A�4vq��Y�	�V7'��͗u������j��ǦE³U�s�7��؁��h� ����{���Fi��a����_�VWX�_�,A[�ߩgw����y�3�n���L��w�������M�M�O�wB5fK~�O�-X~K�Ӄ~n�������ȣ�c�%�A��9A�["�..U���r�ܽa��$#o��Q��m�D`G��O��H����%8)�����V���i��##X�[,��q'%А���z;���)�]�V3�Z�[���؋�(�O��G�Ud)i�h�u�U8JF�'Xͅ����kn�����@��.|������}Ơ3������3��c�j�O�E_�騡�����h���kɛ�4g��[ �
ކ㔅k)U�M����]��էtw\p�҇GI�/�0W	����^�m[�ڀ��|�+y�S���jf��h�*�:���~��rr�u���?���a���Zqpl��S�g|��+�5@�����O��l�#�K����D�KWe�e�JEܒXL��T���E�:����0�������3JKݧy{���*$ϫ����D�گ��U����q���7��'�(:zNT��2�e�`�����3;�eM0��,�D�?�y̢�q Vt���xf�f",�Qw�������@��l+�a��"����/p]�~����9R�zN���=���[9x5�	����s�m�:DbsAԏQ	I�b�k�i5>����){r��ym�Wva�����p�{^_����~�5��ׇ*j��f�(� Kp3�Zk��͎4D�Oϟ�hܐKKr�)NgI!���Cv�?&e
�-N���� S�W��9�O=�LL�H�<73"��3oK�f)�$_�>�f��G�G�C�k��/�ĸ�+���#]���X�����Y%��cه��(zٚQ�w�0�/#��C̅��] >2�ɂbm��<���M�{��F��F��G'u�ٻ���U}�S���׀�����v����s3яK��Ci�Ʃ����̱�{3O&�,�������|�a ���#�f��E�p!�*�_<W@��G ��` ���tj��sU�Oh��d%��ӘR-�LQa�����6���@Z�0���%'�3m�N��s�T$�k��8�[�>h"��ɩ73�\������L�u��+��3ˮ��-BkJ@o�l<t����D։��(���s�1�lvMd�2�a=C�k�4�� �a�{,|�ʨ6������m*G2E�b[�����M?�k»:������K���E��a�yY�O�{4�N��@
2UK9:��7��tfq&���X�yOQopG`���E�]��8�.:=��v�L%�c�Cu��{¶���:��.� �)f[.4]9�e�1�qtS?Q|&���R�Bvڄ��ԩg��I�q�C�wX�iG.�q���3J>�G�a'%mN&����0�S؜V����`�Đ��3pa�;�	���+Ry��~���{_��W����4?F�!�]��|�0G6|��}�r��M�^�����&S��~D"���+�׾�u���X��>k�'���F��vZm�"���W��UE��_W@�c���Q�+�d�3�����U��͉$�o}a���������N� ˽�� >eV�wx
�Btv'��8�!�Ź���ۏu�r0�j�aA�Y�R7&>1�\�щ�xd��`�4�vϗ\1-+��5Z�G�L������O�&Q[��!O�I�m=?�PSL��S�e߳��w��.�"��y����yB&�q�����/�Ce[�v�A<3�M��:�u�OĔ�}醙�Dr��	��]�l{k��w/0�(�o$|�V�� qS��if�U��^��qo�I�N������V��k�e�8��Bt�[i�d\U�B��	C[J0���Vv�5�I9SN3싽���(z� .�I�
�yk1�I�,�A�%Jc(�6T����!�[���w�w��Yh���Zcph��sWI5׵�G-i%s�H~Q"JPV^�|��+9"�c�W�)���I��ԡ��C�ƽ!�F �tC;k�+��x�O���:���EbO�U�1m�	��@pK�/?�;���=5�.��Y��k��6E�����,u�;Qt�2���m���@J�@�Y���=O�����_B�y�!�t�<o��c'[�	z�b�����=D�eww����l�ҕmg	��]�&���cuC�Q��[��ʴ�03��"ɕL������Dz�ک��G����4����tR%����BS�=8g*�䧱W5P`��_?��{"���V�)����M\R�`ͦ%\����(�ۯء�)�cOÖ�DRS B��g�/��s��]L
���ppD�P��2���/��,���N/m�l��4�n�j�%}O�8	HS4Ml�������Oy]z���5n���*�4Y����M�� _��$�MZ�+*��fx���0e����lZC�ޖ�گE=�cG�!�����2�M����{TgiY}�Q�Zs1�FG{M��1��o��{��O�i�����Bx��g��iŪ:+=����i��2� 2nPUm%�;b�'sNY�֓�����-XS��B1Z�*)E��K�4��a��7�	X;ߧ�QP_��A2ӫ�aB�P��Z?�񕝋���}ҷ�ݛ
ߢ�F�!x�Lfa��K̥M�|��uҼ�V+�3	?S���#Y�����ff!�<3h$7���oެ9�t(��ةut�����_���8�r�(�|�(믊�#R:�P0�HC��xϗR�v�+]��L\?����������|��3�WHV��x��C�� gI���Me�ų�g��a���u� ��;��]x��s�]��p��lW0��D�� q�����,v��D�b���s�/�o�	��� .\t��IJ�K	r%^�<��?u(�@gγcF}�����}�u�u5��H�D>��A��' �td?����~�.:I��i7h��Ŀ#́�U�44񏩰4�ҟ���^�Su���jvv�`h�U<}>s`З�6�C�� �56-
�XZi"/aUL�Z�PV�:�,tA���!C�E��y����9�'�fwߜ!�g��M����(B��~�*-��fK��ă���qj����#�:ci vA/��9�Xy[�.����Y�ט��S_�oo��Q����h0`"�4O5֮�xH%3���Q�r��V��!��C#��J[g����Ћ��"��;C1'D�l�3��l����s���K ��m�G�|;)��$��U�8%7�'�$���bm�fT� �O��o.����C���Xb�3 �}���o¤)u%#��`3��#�)[��ޣ��<�'ɖ�g	�۾��E�� �0����]�ʱբz%w�zNʍ��dOE��D�ӻ��ۖ�m�����6|8�
��GɅ�����\�.o���)rT`���O?pZ����u�l)�Bo�f`w5����Ov���'�)�8�Z����&����IEwXG�TOB� 
j���4����fH��J*J��jyv��hP�fޗ��VD8?��]I,��}��s�2�*'=� z���_�e�J,��H?�n�b 30��i,n���.�y�q{PI���f��c"���QrM*�U�����쉇`�Z����Zw�D��]�	v��Rs������=*�[��Dt�������o�Y_s��/Q$�IS>bkv�#>+Lo���O)v�3�ԭ/�_a����p�qk_௾��W5�#��*%�f����3���k"�#�)x�J����rK�5)i z!3g�CQ��a,/Ҡ��Xl�[�Wt��9����S�H��7n�j��-SFA�����L>����*��"��CI���
��!���S#����R�c�4r���̪�\ٕ4�w�r�/�)�^��F *sv�m���쇨!�ڠ_��vr��Z��^����}sM��PŌ9�f�1=�
�N�
�Z��-�䣹��C山�rO�aTP��
�|O+�[����?Exý%�^_�E��ju��Q�b�{�Ox��1�U$�h��d����S��g-Ω4��`�2k�Z����Ց�' xs�����:1T��-Ц2ؿG���D���9�7���<T����<u
����1�����-ݲ[@j�<�'��}*���%z�9���v���2�ÜaC��N�K���|V:,�.Z��0���Xb�A#7m%�U�5�b����M��dk�a�����x�F��&a����a9CY
q�{>GN�
�H|95k��u}��Յ+qA�W}��TK�o��}Ͳ?�E����1�:�lv/%r�CP5%{�8�fG�)����[�[L9��a1t�S��&L>���q���,�=gg{+I�ܾ|X��GiY��+24E������b�NA�5�13�EGS@j�7�+��~��M3+*�+V	2�S+-�H��Z7��鴀9��B�?��!��δ.��0"4�/�}�����AG��)���i�&n�������('+1�F�Γ�	��Z�,u���k��Q;QHQ��/��G9� �?_�	������y%�����2�����U5��̈́y�o�Ua��a��v{��S�˘xCW��e�;x�?t�F/��)��<,�y/��j�g�� 6j�Y�T�7����L�Ѥ�@d&�2�����WA-����0�G��k��
��߇х���k�bۄ��=��FP	��LPx�� �{�њv��N���χ�3�VB�T'q���XW_������Ǒ<���;����[_8\}�.Kr�Ԁ�$��]� �{F�����E�!s(d�$�	0��Mqn�ii�0ً��x^�m
�I`��6U��.1����>뻐v0�B$��@6U��8�d��J�ֆq0�5iGZS)�,��>���� )S�e��k�I��A!n�cީ6W���Z�!�i¿E�wzB�Y�=�����h���W������-d�`ϣv�"T^���Y��+��c>,���_@�Da!���DC^U�!��3i��;F���ʳJ�����nODo{1�c�u}�@KO�/zAn�Y�0����7�&96#���P�z$Z;��؝�{r�h�����m���tѳ�Yh�<���i���o��o�_'M�	����X�Rx�zea�[�9g$�PW��dH�P�9�t�M�u޵���z{�B���Y�1�.�8D���D�H��z}7���/�G�>��sTᩝ\t�[���g�}L=�OX�ߣ�W�˪��F���9��X��X?�?�dM��t`�m�\�I�����X��pђ�>�f��R�+���	'��{A�ơ�L���Kw���i[�FR��s�/�������i�0mh�(�h�åÓ%�8p4����ut���yؽ���$)n��"*grY����z�����?�$EF��2���{j�l�Ce�b�Vd�Z��X��oE��7c"<���@�H�ge�{rY�(?QH�^s�F�4���z1���.O䇭��i4��x���g���E�h=�����:2H�hnkV}�,;=l<s�M�q����-W	S�E1u��)��zK�RPz�p��	S��M�V_��eAM������P���?�6��&�F��X�;]�
�F��k��k�`�K�Э�bi���j�� �+[)�	Z N@eH#����%�z�)���Qxt=7�E�������(g�A^u������������[������@�#��*�����C�����^��F�6�ǍJ�|��K����ɹ���W�������Μ$��?� BU,�H�M {�Ů4�gAv0�UG�)U��/ý�]4u�p�$il�܄��{�;�>�WM��f���b;B�n�/ڋ���`?�%�\|��$$�ǆ��%����¦?�*4������hW}o�)����Ӱ��5���H��D�>L����8f��Wc��H~�=:��i2�$sB��/ˡpת4l�ڰ�+�̩����'u��SgoFj1e�{.U��s;�"�N
���� ������R�1i=��a�)�5�V��]��A�nw�_�� �y�K�d�4���w�b�=M0���B�e�~0>.-�K�Yƃ����>�����~��c$;MAJK~97�[؀=.ˤ��Maғ����;o*I�Q2�ci�`���Op�h��%.w Ǭ�-'�V�/{_6�#٭[��&���xІ f�}T!;��0_8��3����|����IG\ö)���k7�8 H'�P�,�a5v�[���A].���ݾu�3�3X> ����a����P�J�{'$�p�60���?��^�ɑBVgd@����%��{в�3mi]M� ՝swM�HM��&RKӖB?�am�}��8|�p��ɋOɠ���^[��8��\ r�#�}�k?�7u�׊Vِ��l�̨���ס��5vN2��v�O�������SA'��t�����l�E�XB?pT�Joû�=��k|�&?D���E���J��eyqm:�<�!���D�ö�8]��7�[��-*('��z��_�0�Ied�tq��O����0��,�����nZy�1q�j��~uqf8.u"bQm-:ﰆ	�s�t��0��M �[,�����~]����f�gR.;��=���[���/��+�/�9����s�u3Q?�+I�9�kQ�>f��J��)q�i�/.�-*a7���
�p��_��� PX5ݭ��=�*��f�sN�3r� k]�R��� �E]�)4K�U�)���!�C�C,e��(�;�!}�;���DW/9�wX�B{<H��7���ig�A�֯"&�n�>�d���LaCCFťe����U3-#Ӧ��,W�� w�����E�4(�ِ7�wE�0/�ׅyv���N� �A�?�lm�\��M�����[����%�=���!�1�a}������E��� ��%�qхh���$��e�5���#�O�D:��%'@|��6�S�� �EȜ� $p_�S�%ۍ��b@���1�*���&q�U�Aqh��nd��5��ٱ�)��}�B����m�AZ>�o��VE'{�y߄����!bTf{ЁL߿��tA���ɶ7�	����фu������$*�-x%@er�<*�B�80���Ⓛ}�J��tv��2O�5a�h��!4�ř���,r�ը�K��0�v��`�m �`�E�b�s���M5�%kx'j�*p�9!�AQ���˃j5$aT�4Y�� {ꮐN!�{
h\�90�u��㽏���q\U��	E�/g�o�Uo�M��E������:�)v7�5%���C+��{8�L��a�$�t�߾[��?9�ý1���S�=&����pCl������g"N\I)�_�9�,X�6�G�A����@�ſ������N\�*���n��SNҵ���<��F�b3��F�	���+?#��(`��j\��·F�1?�m�!��H���70�Q.j��}G���U����hX&��\�tW���	+l����9L�x�����0g��,����#ő�jr������G_�X^����%a�!�ZpQ��7�~U�:���:o3j�4��íD�	�sB���e��&x �t,���T��W�:�����E?��0�jqY�O�l7����ѿT�d��������s�-a�ݥ+��GZW>��K���ߞ��_�F��ۿ��=u��Pu�L�8{��VǙ��;�$��pE��n��B\��q�ay�B/ǹ�Q���	<)��m\˧����#}����r��*�?�x]�<s{!�d���/fP�(fE$2K�=��q��xi\�ȋ�oY^�l\�/�I-��z��s&�����������џ�ݚE�U�RT��QXJ��7��
!5�d'S���3���^9� $n��Uk��I.��A��Fc�U�6�����5!{�̿x2�w5�IY����P��h��W���C��-_�J���#"�wj^ᒰ���+�0cy�~�_��?%��W�ACe!�2���;!�&0���Nfx��8j�g;O���1�t��h@&sa/��t����+[)�El����p6>݇�ˍh��;Ǩ��hm˰c#���������3��l���Ռ��J��j�\o^�{'�'&	��d�����B<���e��g��������@��O�˾$��CFIuy�刏 x��5o��:�L�"ɋC��`[����z�#�G]J}���`�Đ�tH���s�߸�U=nX��ڿ�W�f��=M����"��(n�z�mM��`�T�\L5˞"��"ʡ�H�'ږ9�R��m�zWd�Z׌���U�L ��&����k�7�ꍾ�v/J�΂wFz��8�m�Q��9:��л%���8��w4�e�0D��uXyS���|�Ln�ٵ*<hY�T�rw�v�����$�^��Y�ܞC�&Ae�@��"Z�@7�{E���c���NH���/C��-�{���Y�sfQ�Cos�g�F�m��H81�a&ωB|�h�>i3F���4x��g�&P���=�G���Q2�cn�w�qi;@!sĜ���p�b䈠�Sl��1���);�KZ��f��[J	N�z��]_b�:Ah��WזPo�h? �j���G��{���h
U�]F��B��;e!KBf��E���+��W˛+?�	u����#�8��`\P��S�����2T7d��^+�/<l(B��N�,u�I�ڤ�ڹ�%����rܪ�e�#�<ͅ���>���.F�0�aY��B߁�Ws7�>���5�N��AW�"�nܢ��x��O �BwM�	�ũ�g�ߺ��D�p���lØ��U�K]�n<p�Q�l��ہ�z�V�^��3w��Yצ$��b֦��i��/5���C�6_�\�N%��P���yu%�]���i�?+M��z����0}�S'��|���pE5 :mH��D��C(�S'��jks�u�Z~�:�zi-��t�@�������(4�,���������u����yj�sp��vU2�sb]���Cy{= ������l�iX�a
҃��V�U0�A�(lߺ�z���y������wU��՝gM����` �Bf�~K�-���Ka3؃/���ʱ��.���1�c�uHAe��9��6[��.���Rͮ��	4(o�iQM��މl`���O�w��M�%)]f����w�V��ڡ4#��R[��ݽB�Ё����$5;�Ⱦz�!bT�3^��!�©e��#�`D3G*�)���8�8�x+'	������\|ԟ����q3i.�Ć�9gD��Z3������ �s����y����;��	�����r�Ɍ!g���Q��/$p���I�4w�n�B]��'՘�\wm�k���i��n�q�Qgm,�L����|�B�넩�ɻ���ٖ%��R�/�jrC	��x:d?&5u��3V٫Q�l�5������\�5�o���O,'袝��n����^�ܐ��E�tX=�T�<�vg���왡����X�Ms3J �yl��E���QL�09PD.h,����R��B�(�(��'��-z?l��K e�	�O�30�y(�2��so���N����@��c�{��~-��I�)��mQivސ�#�f=\�$G�Ѣ���Y���}atlf�&��;]���{��R��k�*G�<�g���@e�fp��K�ox允��(��a�
-���8"p,Ś����	���S4>��50��O/RZn߱
C��z��Z=NR�E_�!�^5�g.�s�����1�:�,� �Ĉt�lw�7ZmgCDl�}��|Zu�y~�A�s<_O�tX�hjZw	�(�c�����/��AC}�������f����Q�(W0F�S�7��Y&�B����$(�ݕ���Y�FĠ Em���,���Ķ�6F�)(&�M�������T�O�c"N��<��]��5H�����v0P��G�O�h�B�|����3ԣ�ܕD��34~��1p�i�n! �`jPC��j	_��O���N�"nz�HM.��63�D�|!�(ȼ�@*N{����o����8��ݪ�6�}��AH�9g~䐧tJ1|f������'�˅㔬�]z�➨�@��狵�?"=W�GP�r�(˲ME]%{"�<b/��o.���7��l��{�Zp�O��������DB�e���7ƌ�<������n��-�_ �#*D�Q����[���<���5����~� VC�8�	8b��s���t6�j�0���9�M�5�i�i�ހu���-�̤pm�%=w/�����şq/{&����DC���q��'RU�3�R��2 X���T�����g��b�� ���R֓��kdvG����)�|R�/ɽ�&Lo�V�0��sy<��:�߬�!�Qg��>���-�Z�g}�yC���_sK�|��X��S�[�T:.��lC�a]��/�7�w`��-5P�S��_ػ�Q��&UdM�o-5�?n��;`�/ۅ}9��E/QD֍�	��#��-��#�я�2/P����TO������o��d��?�k�d-\5�6�	�\-��Y*�d�ۊl�Ԣ��]��H���Y�n�_����nVFϥu�x�s&�-���2u���V/мw�nA��Sr5�
��!�ȝyIi9
����@z5,�EC#�:�a�ov�ȃ�^���.ZY�Ź��"}�}?8���kZS��g�ufͯ�o��R�E#�"����4�b��=��|3[F��oRf�t����mhF �J�IG
h�|��!@p6����G��@N�7>seIR?���!�v&�k#p�$W�M�TQ7����ɦ�0%�_ѭ�\#�4!��!@u}
4�������>�#C0��U\-�B:�!W��`]�kTf������]��q���Y�׆��XD/���n���8��;0�r.^�Y,��܉E<)!�h��d�tq�r����/�T�	vAvU�	>ܓ�Fl<�3l���O���k������z[�7�>؏e#��P�
�os3����9�(����GM�݄�����e��֦$H����.�(��*�&����S�ţ��$e�r�*�(R79j]6ƅ�?�dg��Z\�#(W��p��G��N�L"G�mN�+?5	�D����DO��<Y�P�7YpLL����=~�R����Ɨ� ����^��n�&�jj���2��3���+*�Ch�q.׍gr �����M���2xUX�E`�8ω����'�l "�(%e�0�e4�}��Zwk�;E7�������˟p�����y��(�EEZ�n���?lу�e���AE��ZJ��W��1�מ8=N��<�B���S2 Y���F�9�%�Hc��o��5��\ƁOSf/�F��[\̧\ʴ�/���| ���?��h[l�	�T�[%a.����cl��75��v�w|h��6�{��AY�K�ª� }5��L�����f�?�ߏj���'F���f��s���șs	R�KF�Ǌ�pxC?�ކ�m�$�������D�29쩑�G]��f����qm�O�2ڡ�?|�>jGG�ZB�x���;�_�K��@T�V(uz�;G�7�L.���S���,\b!��IeT�������懎'��3��~�K7$�!2"�fyŻ���r���������������C
�P߯&��"k��������;i�M�'Wl��s��(��-�XD�2�����b�3VCU%�'��f��k����D��z�0�1
b��{�Ug�tjx�Zg�<�(ݶ�I��6��$i���-z�w��'�?!~�0�!�+�Q�Y��*	�1�7O��IO��;W	e����	#!S$(��E|�v���\��l0�u��>�s#2��y��u
�S4�=����>�	p0d��U��,��ʋ!��z�Qްke��+)�®����GZ΢�7SXe��p3�陜'1�;�*��㠴CQ׼ٟ�Zn�)`�h�6)��4&r>&��%eŉ�fjv�i}U�|�>�7��W�U�d�2��9����vyj�5�b^s/w)Ʀ12{ݑ?=��>K�G��Sș9����_n�c������MT�7�u[��G�L�LOF-��6�؍ݘ!�������T`�M�m�����z������v!���f4���ݴr�j����i��t��+����$���ߛ�P�������3�Q؀\��MH#��`����Wr�S�^�-����3n��	�b�PnC��@՗����1��A��J����5N�*�w�d���5�ޯ(>�q>��2�i��$�I�(6�>�����-�_�Iq��n�]C����/e�Kc1L������f���/�_�/�1�X֖�����KPШ6K�2x\XJ�%��Sff��XL�p}��z���I�������7f%��X��re�r���7W��qd/��O$�=���=	�5#�cT^QOS-��������'�Q>�N�"�[�S����=���:^�|��}v��f���ǐ�-��)!������*�W��;(�U8f%fK�7!x�X��HO���aX��}�87dz_� ��t�o��*t��$�?�R�X+�GQQk�V�ݍOZ�RDH_*P^�)Ng�����\#ir��,���˦D�t����TBg�L�l�@��1����ZNA������t���?Y�~�p�k��|?/�2(A8	Z�C��\˒x���'l}F��A�%@n�7k�����(��ɜ�&Oj2�5xmE^@,Y������6ۀ�([-M��Ǻ�z��.���cw��|
f���Q��G�@S�(4�Ѓ�1y�V�@I��&�A4rѭ⎒J�s���y�@�
 t����sm����$�'��J���K7��;`ϩ��@�Sw��d���[�d6�Q->7an�{�`�o˅|�1�h�0Q����X��`-�1����}�{���a��>ψ`w��������˄k�����522���#�>�Y�?���&ᒑ��� ���S���٧�R�n޽ώ֬�s&�lϳA+�2�g^�߉��";n
��S[o!�!���y;��րi����Q@#z}����.VŕCBF֘���Q�h�Z���l"F%��*���Z|Qgc��f6hso>���"�N�����4��	�f0�||c���/)oۤztL���6m� u�$IP�
<$�|�"T!���)V���r�	�7'�I'�َ���j��#�4�$ 1{����(��j)��0nY5���#
�0�Q�Du⬪4�v���>�*0<�'U�}��\�!����)F�k=hw��$�Ϻ���z'a�=\X�;슱0���}��F�;Y�v仌,��ה��2��)�w�h�I&�}��rO�������%�v�PUQ�>��f�/�C�<���պ���;�g����|��>�\�#�M&P�-�o���e��9�Z�{18�6�M�Ԝo��e��M�3�ܽ�&U*%��0�9�|K���eч]*�7��6/j;?Q�~�[�a���W�zi��^���Lk��m�Ŕ?��XD��o� /�%ք���`A�L���A���ۂ���妰0r��� ^�
�o�-j�Y�{Q��[{��N�,~T�j�׶�m ���Ox�\6�x�^eE)e���9���KP�� k�%΂-����&5�Z@ �;.e������ ���dj�S�,��(:~EZ�� ���0l�g�7��O��Ý^�W�]�O�����8&.[�(�B����uY6�(F]s�%l�c,G�o�����2ƪ��S_�?ү�[�~�\s���=#��Y� ���?A��h�!�	�W[��y�|��t��lp�5�L�v�@h*���z2��'�Y����sٰ��d�5�u��E�a�J��$]���^�³� '/��oF�s���)�=@��aH����a�m����JتE���T����NuN���v����J��.�_һ�}�:�	�þo�y�7v��[[=�͈D�C�;�3��9{qH���o�pHk��0��Ԙr���ޤ!��Y����հbѮ��c]=*0�ߏ����b��oxC!n솿w����F>`*?~��'��<u.6ۂ�q�(�Ԕb^�r���,GՔo�� ���&3�b��*�F����XRi����o�܌�c�AsvT��	���{�MNZ���`Ϲ->ع�i�j��g�����[P4/Tz<�٦�B��#H"p�e�z���j6�!�菍�"�"B}L��(9&T����)왜������h�J�������� rbiOچ*�j��A���.����ah*+�����n�]�N �{0{�TW�"� Y�R�U�cx�d6��D�-�d�tďM��+$�πܬ� A��U�\X����w$��k8�ED ;_�~��(��O��Ks/��:�=BX��B��n���[<���<>��4,߭4�:��a��q�	VNw�ۼ�Z�|��:E�C����o�{Ȅ�Z������	���*w����hU��5^4W􊔳�$L���-��X��b���m8Jem+�vG�/�a�*���ֺώ�<�R�q��J��L�Y
�\�{#��������n{�``�v�5��(���q)�}2:)C����I�E6V8���� .$_#O�q��'��\CL��:8�K�e�Lz|r�܂��;���#/@�X�/f��|4K����s�؝I(�\�L%��f�VX��>}���AIt��8�<�1N�%}�O�$X9��*�B����Iހ_⯲h������ � c�^��Xq-�Τ�	jMU�QI%�٢P�F$;�
���Ա�Te���}A�f������٭B=l�ݫK�b*'�1�G�@� xcfP��K`��x�,�ڙ��h�Vac�>���B8c���jī�=�_n��3�(���f��=R:e����c|$�����:�R��_���^篢g��轑��@��,�٫���tf���g#��l��\I��YI�AԚ�?R�t8�J���d�o�7Χ�/�|*A#����eN�=ᒃ�~1 .7���3av���:�"�]�䙇(��Pɧ�x��  �mp�,�����}�6&�(�nMΨD������/|Dc_��g���i���%��g=ϯ��P��ڂ/)Z�"����VS3�4�u����Ϭ(��I��!�*P`J[˩��j顲�/V2�.yunZ��ME�6��\©/� M	{���Oߑ���=*6�l�qZCH��tg_������1\�M��C-o �իTX����]Z�ƞ�ޥ��&��jZ*"�;�'f+�RQn˒�@]b�"��k/��.��k7���ʮ��:��O�C��`�e03�;E�y�б�R�t��Mt��'ĵy����t�A��V ���f!�b�"e�����۞G�~�>�Q�j�W�&���;w򙝻I�i��p��9=T:�Ak�ż��8���Q�Y����sL��J�GR�30���Ou>�K|�,{���V��� ���R��� >]d�(�f��a">�y�
�̱��cH~�3{0�2yY�_:k�[��KQd&�>J��7�g��.y`v:�r��K&�{�UhSJ�?TwD{
��޶���7��3`��2 �S��T����oQ�d�S�-R�nz��`�f��.�|b�Q��ֺ�|}��v5-���uX ������y�q��3���)y�`��/>kxz���5���=YjOyYci�X���T�e[�3?�������Q�n���"�8�+z&U���U�}2r뤻��M�0n�wS�g�5a!�K\���i6讻f�@���������ٕW���,R��Z����Z��M�'�z"Z��� ����Z�gw�<f��BoRv��N?"��T�A��4� ����|�.���o��Dt���J�� 	fIdM
�Vq|��!=�=p�DL����7���I;����N��I���\�##�$���1�\�oN���Bv�o�0��Ѫ�1#����  u�C�4+��̢m>OY*0P��UY�����!>#g�=�!k�5`�g�����ΰ���^�#�X��%��o�y�Ԝ�3;����5��L<רY����)��xh)������r�y��&��QE�v��U��>��y��³�P�W�i9B��O����gm�J�">��#`k@P��o0�	�y�9�"8���g��]�a1ۜ2�e��s���/���%Bt*9��(��g)ӑ�^e��`*�Yy7��j6��6?e8����� WW"���>�O��L��mK��?�)�D�Z�!yйC/����c�L�Yk������r�Q�9��P<eZփ�^�[��Ljgza��f�p�L������-2��JL� ����Ԭ�p�rx�S�E=�LH,�x��� 	�%b������}�ZT[�;�"��"����)��7��[�(�Z���:��l�	"�����*�WY��k�Ƭ�Ş���=8��h�<1QB�����Yʕ�Fquo% ��@)o$CU��)�>UESs#��Cf�[�T�\QF�;�g� ��?�U�h�6�	�j:[�6��l��&lz^5��vVW�h>���>��;&Y!�,ţbs5�����5u��|Y�8�H��f���p'��ԃ��sd��.�=�\�un���a�͠*O��Z#���(a��.�(�bo�0�v+Z��|��0*.Q�b�Ҷ�:�e.��=��Uv�mW[ц=�X����F���F�q܃KÃv�H���DJi�,g�s��80b�m���*�Ab�$C���*+{�s=~��bqb��o��n�ޔw������*S�N���<�b5��W�-���3�w�"�|�ݫ�+��Q��St܄u�)t�����G�ކc=?E1�Q�c��N�#�Of�L�+H?,��0�"0qÁ����G:��8���ـ�
+�G��]�O}o-	<ů���F� 38��]����$O)>���>�s�+{!I�ޭe�����f���k�`	B"�N���#�M����C9@;�my~��׸���01r&p[�j���z~W��f�'�G�~��]�޳FR��}�ɹK(%�Ŏ��
y�����j�FF��O+�'BXCBMw_k��g��1���%e�J�S�!�8L�ߎ��`M���	5�g�Τ»eC}��`>�agߛʒ�{�1�:p�s���z�#�*����i~Y�j]�,6F�ѧ�p� R�	_���f�
����-W��=EF�j+�X��wX3���AٵΓ��pH���|u��m�sή�@����x��b�2L蜑8Ư���~�'�]m<92�!U?ρ�>�%G ����Vm�}�C_@x�����P�T@x�u-�(G��oL��g�&p �_I�!���<kT�I��?�暳��]���Q��j�x!Ř�fl��T�rY!@��r�(q�����v�����rߢ�=:-ʩ]1�+�I���|Mڲ����Z��+`g�-d���E���^ JbyRdC���թF��xC�6�x�q��+�0��bYYǈ�tt�z��<�����iȯ�J����u��@�
��ӂlJ':�)��ad�NLKx-<���־w������>�[t���e��c\��d�A9Q��v�#(��\G]�ppA�YR��c�1��\�ߵUv�tr�=��~f��pO���@q���ca��Q���X�X'=���ry,b6�3x2*ʤ��/Aj���F{�ŗ$O�fE�B�\��X�i���0W}�c���0�$ѷd����m<��v4~n��
�����6��}��B���e���+P~T�c穙�/�����ظ�y�ҏ˞��P{bAgj��#-�aç�x��خ����E�j�_����2�(����ԅOjl�8wUqvjp���z g�2`��i�GD�_�f3�~�a�2���,��A����mAϗY��gL�k��.1�h�����Hc2��TG��Y����3i+����J�3��F4��(��od������	"�@���8�3 �e�	>��%�D���7�JN���@~`DeI���ќ�1r2��I{I����p�֪��,���[�%�hŋ皋{�J�����K����֐����E^�Z9���x�_�+����o��q�w� �6ew�N�دk����+V���r�#+j��ձ����N�ڽ3�q`zVi,�	��eIρ��2� ���gQr��R2u|�R��~���Ӑ�u��:��ޙXc0��?Ś��r--������
k�Ȣ��UB��~+8�ci���28��e���<y89�`�P} M�V��L��#���zL���R��?jJ�����;2�9�����jn?�w�S�v���� iR�2�j��G�D�k�h����䭴�c큄�����|�̑Y`��NTی*Uq1W��m��J���i�G��YG��5�u+E��P��3�+q4����		��I���ޖ$G�@�Q"$wW�G
��S��ۨn�
2T�7Ju臙G��Lۭ�e/ؚّ!13��7�TM4|���浠$�؋.�,-��/�!`�Ufgd��r����J_�Q��꜓��2�?Lߝ�D�m��}k�F��)��M���œ�ա2g��U��=-��`���ّ/bT��Cú��D���/+��RW�,y����|0u�b4g�ê&t�)�1}��x��$�0���z���4@��+�n�}J"�9���a�JNg�b-��/�xw��8����9��[Ϛ�� ɳcwdF�m,?U����(M�kGX|]p�-�>Qc�v��׬+�0ngt��=�D~a4Sp�7�������ap��ʷ����%X="O�m��iĢ�%qN
l����F�/|s��]	�{	�$�_�Eѱoc�y"�i��@�kk���̲|?u$,�Hɳ�U��Օ��~�3�E����~6|�P�^�0B��ˀ}��|��~/Q�c"�Đ�~%��,K��yq�k˹gP��paN�Y����q�s���	��G��j�ϫ�v��2����ۆ�o͍jg�?w�v%V�Ay ⿩2;3����D���a9��ً���c`�X��O͛ћ��|%�Y9�?G�G�Ck1�d�"z��94�~��G>�Y $��.�+^�<���L3�(�4#�j����2;���g��@�-��EJ�3
z�����w!�D�$I��CN���@��ej���1��E��F�{�}e-�@� -(�sŘ-�F�Z��c�F���tU�r6�t/ن=Y%8~c-Ep�P�}���a�arg:��{]�X=���ok^���sɧw��<c��R�/���.�{��$�jES���M{��i:����aO����~�R$n%��50�J]Õۤ~5b�����5w6~NVàD�B�$�Bw��~��~q��c�����S���:�U�by�Ϳ�{�P��}^��܇u2��LW�uAI�K���-2je>�x�u2̓�VZ��1�ji�Hw�/v�E�� F �2}�(£��OlR�Xt�ǃ��ɜ�9�㛶�)��أ.�ͤ�|�V���;!wh����WI��pJQ栣� �(����r~�\��}.���������J�eB�顏1�
��S��}�e�B,�!O�N���W�:��R�!
�q�o��u#��~f�d�\օ�K�W�6\m��6����N1s\ �GdS��	�������� G��c�761��(v��6�Ղ���W8��K�6���wС"5�AKO��� n�1�k�U��]cٳ5ڤ�G&s����=�u�Z��	�|r��SC8��Ʒ6����荶4����@��r҆�SoY�*�M#�Ys�@���<�T��?�n���/�Pk�)�,?Z-����qG�.^�l�=#�K&�]��ms0�7Xj�-��kEh+�XEs��t�IX&*��r{$8zW\�1�"�D!U9�s��c�n�>�}�Mi�F�u)+�@ϻ�S.$Ŷq>��%��s=�Mc#� �YRYO'�`S����ڭ��?l2��O����D�4`�UI� '�J=,5��y6F��k�5���5d4�d�;`�����$5�A��U�-�}FЎ+�4�cR5JK����X�鎍YTsB�נ�����s��É�,�cb�`��-����5TM�.��烖��w� ��z]���rۣB	p�#Ϋ��Qz�Zj���{��m������B�:'���T�5���Ƈ���V�Ŧ8���x�k&��9[ �54i��*�g��i�tA��.���U�,��W�<>i�I1���R;�t��bmC���D_T��`W�ۂ��:�'�WPA �M+C%۹�М�E]gT^��dL�^�5P/f�u���ӺAI���7$��En�\/�����'z�jL�x�6G�T�Y�J���Α[��A�G%��G��e��I�K9����шs���A�Q�+�tp��e��u~&�^���v
�g�e:��c�">.��=��� '^��2C3D}p���K�߸���
HnP$��B�Ӏ(��*i���ilB��V�Ev��
Bʚ�8�()wft2�^�ҹ��7����9P+��+,��FM��(�Hp$�qq�eo�n���E�aR�,����(h��n3�.�=e���i���>��y�l{Jl~T�0r��-�2_k5�=�>ܽ�w8��m���B���X/Kt%v��䠚�������'�6'�rc�B�74:m���kX��a�rl��V�;~��+�W|+p:��ޟO޴L����vf�{��8����� ��ٍ��ja���"\@��?o9/�O&rH	+�����O��a<G��ˋ3�+}��s�;�
}<�&*�ELv \�B;;H��x��^�;�����?��L��3���V�˚H'�m���A�9�Q���҃׌1ណ��Z�=�{�`�q�Mp�aq� �m�t6Sq�s��-��Es��o����A��l�_�~Ɋ�.��o��߬��2A���-m{�YV$�o��Sn��<d6�; 1�ʣ� �J�V� �;Ɣ�h�S��|�R�H{}QAA5���(N��7���}s����] ���7�o�!B�q��~�
ă��'Y~}>�tB�O�bQN���W��:طҟ
̠�oPr�'{�c�Ud��ťCW���\}�V�������1������dؔ�	�'�DP��I-?������b1���v�wxK�M��v}�#M��;dݣ�H��慑�&8@"�%�=�""���^]h� �=��X�&Xg�v�t=<U�#��*nb��O��#�,O�'̑�Ԭ��s������=]�pJ����a�m��3�A���V�"�;������%�䨍�9;v�xׅ���Y�S.����;F�:��{K����vȉ�[����AݧF��h/:qey��,�H�-?��5�f�+Fށh������G<b�d����m*I�|Ȯ�O�b�o���n	Ƶwr�D����*<De��(<�g��_24�����I��w���|����<���Q����>�x�H)�MYm%I�u���o�.?N�Q/�k�#����j�+��,M��b}Ê "�>8(��8 ��	��+^���&m�}X8�<���7/FԎ8v�]@L�ʧ�_)$Ւ'�Os��Q����'u{�|@��}$.�s��`҅�7���,���'�}C�@��w��Y߀���-,1�xpd��-n�zǐ��� ��З0~>�	]t��F;I_���P�t���M�JI�
G��~M��3Z�F�z+�l�Xl()w]
ĠG|Ab���+����~0��1�m�R��L���V��<��212<��L8��
��!m�ф2�b?t��>b&|G���p����W@�4;�+b�\�$�r���SL4��F���@�׶��J�� q@�s�r�[��\6W�S(#*�̩���Ā�����7�W��Pt�^�9�ZO��S��q�9f^:��=��&��I�v,��`2V�v�k�pv��Z�sZ��t��_&�{-�88�W�>Ā�9"!��qs�:��,��'���4�M�닎�����t���ͽ�q�K�ھ�t�|�M-�����xl/�ϒ'a�¨h�)ږ�?uϐ�x�p��G4�mBU҃�'6u�,�x[y���twG���	r=4[*����ƻQU��]u�*7��^y�V�F�ӝ�cR�5O���!閎v��sKp���\�/wf�b���L��X9`��\-s���>�e�W���0k��hHl���z*j�;?%B�L�#H����z4{�0�vএ�Y�"�B��3��c�T
��> ԜXN.�Nv �?�:�4���"�� ��i�%*4�͜ҷ�A)�.���D	�W��i�OP�+�R;�Om�
$�C��D(�	�I�hۋ�sc��'*�nP����TC�f�ș��.w�Tg1n��
^scP�L�u�<���LA�a��*p�-�}��d�����6Y��zT1�
2xu�{�=O����97[�/�XT�%;<��:����UI��و�׍ѱ���)������ʖ��uG�^q��E>ѐl2�[x���I"����椭���j^���C<xp �ԏ�>߸a7�Y{�L��0�C�Y����b�2/��erd�76�1Z�J��N�Xt��%"�7o����J9��W��FV�˜_p�Ϣ9;(w^�'$���&l����u�_��Ed���y5���29`�ؠhl3�B���`K�EQ-�<��'�j9��~�ʐEp����?���,�@�\}%�MO��n{ ����o��0��IDe���$�~�GC(.(	9 G��E.�2�R7N��z,޿[� �킋o��XY���J���ǆ�fHB5Lz�T��6F��n3�+�u,ԦP��c�����g�w�P�+�k�M,��;Nv�[��E'�G�k��H>qz�-o[;]�0��+���S�̵Gǟ�H{��z���߯�ŌFI+_���m��\z��=
̰<J&�WXO�̡ubAbvԱFcy�y�f:�E�y�.�����4�$��H�s����-{��|��.�7~f�=@�?�_rӈ��	)5I{�M� >d��Yp��1�Uf�Ė�_��z���+oe�yn%��x���w�kU���y�'��j&!�;/�􂰉���؉QG�!{�\���aG�<�Y+]��/�z�4�3����|���	������Q<韺����b��˔��|TW��@J	JֽN��p۳�VZ���{8��ڤ��P�L{f�ۨ��!�,��� $k���L�h��n5���1+�[�g��|b����p9��΍4�<J�+H{V�f[Q�A%u���ߎ�AT�Ҥ��J$�.��u�\"R���j.�����E��z:�����( �qq`{2Q�㤐�I�='6�����_z�Qq����GhCCh7�E�K��L��S�q��ۨ}�/W�OXx�$�ep�K>���
�m�� �\:I%��@fȏdX��!}�ZZ��kI�\��)˓��8%��{�;����I�}���Fb��u��߫Mل��WF2c������-bwd�����Q��
�0���}눚���2����Ϟ���}؈\f#���rkE��P���BA�*�=>��#ܴ� ifǎ�K��>x��ݗ��_zLa:#䳟�8��e�d|��
��J����z�x/sR�D������͊�8��q��R��^_�M�^��^g�y�T(qUq��,�@�X�t]W���Og�<tl*5��� A����A�V��t/���g����og�>��g>D!�v6fƯ����yr3�)���/�^�1�W)��P����������7���E�-�/�Mt6d�c� ,�c�'�->��_2d��R`b�@Cb/c�Ò��AH��v.�K%s����0T�tb�>�k�$-�xe(�&C�1�����p��N����+c]�Þ�K������Y" �Q�jI���!˕�]]h"<"w̸/���.�7�SƸ%���=�O�V	��P���=�D�e��7�0�<����v��ȭ�c�ڵ�ƋyD�{��P��w.�_/s��A���П�\�V�Qi��Yb+�6����v�������l�����	���PU��돁,p��=�H��<<����Q����6�����k�0u_R�A$3�ϴ�u9z�1Ź�������@�%�* �D�RYS���d��L���������ެ�IA�ى*0~��y��:Q<a��=�Q�L4>p��n{�p�g`�y����XzhK��=ʻ9qSp�nT]�I!���D��>�y7g"`�d:�R�S����A�2)d0I�-x�Dn`��`�D��v2�򢧬Qgp����{�r�-�)2�[�o�5�.�[Rw�7�ڣ8�D�x߻��^�k^�bg�5,R��sPE�Y�<���4�̽��K�~�Ԅ����1�ׅ��?n��ψ����&;���g�2�;n���3ݏn���SU���[�*�1��Ƞ-oi�>]�B�0@�:�B�(���}<��)�Ȇ�m�bpZ����|" c��Õ��RZ�l�g2f0J�ox�,�h��"��s����4�����%v|6��k:o`�tƿ���� o�I���
���|��!�psc���*��×F7!�!Ia���q���8�d��#3$�$z���mq�Յ���fNl�0(L��.�#Dg��ˬ2u�lN4�ԑ��>5��0��U�!����!$U��k7yo�=�� \��t7�t%��I�Xg��k$/���9T;�L�uͣ�%��rܬ)�)���h���}r�:&����1v�2U�i>_�ʟ)-�v���O�f����a����0<>[��#���P��oW�`�9��6��V:j�}����i�
e�&3��^��ծ׽���*_�H��~��6z ��eTG*{2*7<�66)��?�/���}�򦯑W���X��5K�L%؆m�9j?���D#r�ǩ|���U�T��H�LO��e��1��NX�䂝U9�w~|��Z��1�K}�����2X�s�؉����4���ʨ"|`�M�RQo��t�����z �II4�B
���|�K&! �H��q��k7�A�Iꇎw�}Ž���J#��!$d�c�g��?���R?Vy�0R�d�zq#� ��r�u��/4�������>3*0 �U)/¯:�!e_�-"k�+p�����P�Ϟ������XQ�ꊕ�u�I�%���;�K���Uz�xA�ܖ�v)Φh�Ta�abrzí�ᩑ�!C�v��mU�W�>�z��(�� ���9S����%��W�f�'�9.>�� #0�3P��mo t��I�9_�q�_C�Tv�1����7+e�Xh���{������*	ղ��J��`���a�#e���*e��7fv�6�?50+�����Ђ�W�9�����F�LO0�m�d?��"D�y��pЉ�����čLy��ɋ޿$˽!�����-����R^lU��S)�j7(��_U��@^զx�����8���
 ��"��R��@ !xb�=EX�.���1�o\ O�%2�ɒҐ���Z$�:;�ؕ��a|�O� ���枷U6��2�(���Z|���
D�l���7(�n\�'G��;���g�����8���AGB�7��&[Y�S�FA�%�i�o�h������/SC7��Z[ɜ�\ג��d)�`]N �/�?��[h��	x��[�N���}$�X`zl�?<5�`�v&��hm��kz��Y���WHP�2�a5�-���>!E:LWlg͐줂�'�IR�S�as4��Z=�*�E�T��a��5���c�J�����������o�2�%��Tv���L � �K.!�����:`��âen��vCv���[�\��(A������
�q��3�Sn�Hϕ�v6��{��Ҳ���=B����2b��U��W�*�v�C�᝽�CbtG�o\\=nP�^w�l��\�*#i���><Yb��恤���
���ow���|�?���Wo�+�QwͫD�-��x)���R��|y`�V�E?Q�p6����#r#`�f�+�O�,T����k��QG���We
)�8�p!�P�W+��-m[}?9�<�5�xIF[:s8��]������B);��/sÁ0K1lʮ�������$xߚ�R`ٳ���������˥C	��l�N�'ߧ 4�r�1�� p+~���i�zNP�6�{�F�~e/�]{�F"&G�MG4��������A}
IL����ڔ:�BF���+r��X�;w�#���nAe�T�&����I뤝Y�m����j��<�Ń7�2XN3������F۳�(mH�k2Y/�?�@�>�0�Gl�wJ���_�~$�~z��)@TL�u�I�G�HL-U`�2!1���!�����T��r�����h����]���2_!�qf���`��r�%+��f��/���J�_���er�.�4F�����7���:گM�Gq�b�Pl�	-�L6�Q����b�3�Ceյ�0�sN<�BC������0���beH����t	��PH���(��:B����#�O��@�N��n�J��/�5Pa�KNX]t-��u	�wz��2����\[�����Tch�dWah]��̘(�rxG��pM�f�HCc�����˵a�t�x=�P~�Wpp[ͦ���x��Ya�A�藤���?=��i���{3²?1���ʰ�U/� ��@R{/$[7�E�{����i)�G�����ǲf�$ݞ*Ʉ�v�y����~$��ߖ�[���6�����Bn3��qǾ̍�~`��cs���;Y|�U}���yB3�˪<PŶM�U�V�|�m[��&غ]��r8j��ɇ"2���%.ԥ�i�j�+wa�Qv�h� �� ��Y2l����
�D����dz��)����J�&̈́`Yj�̫{��fY�Y�믌���1���QR��F�G1G��bY�cឿ2+���Z�^3�	443I����S���(�l��y@�.��non���ʢoB�=Gù�Fl-`����-_��d�<��8��;)�9�v��~��lwy�h����E���vƢ�%'�:�9�v~F"0r������=�+K[Ʀ'�y��3�b��2 �3^��-�\��lJ>e[��$.^��-J=.��� ���ET�8A��<6z���[Ĉ[�h������)����lw�H���z
v��\�ٌTFҳyS1�IS�䁗�H��5�7=�uT���jj�ϗK&�ݝ`
�\�N�L#�HaI���K8� �j3�9ϣ�g|y,(���-����k�����ا/	L��H3ǹ����R����O��iK�V�5�笤��B�v���K�c"��ԇ�k��Nl,���*20Ɩ9O�C�xw� IT&k�T�5B��O�M|�myE�I}���.x�5����
diV�]�^e�n?E��X
fT��=Z�p�a�Ү�7��'�n�⃱��,ޖM��zhJ$o��q��������`�6�k,'�����eU6���v�2�'�e�)�;T�>�8r��vJ�'���=?ԂW/���Ek����sz{�L�`�mJ��m�Ӧ��X�%k���5�խ-]��z��JC<��r�
ь��:b���!׭(��rAl���~�H����A�:��p��X�Lԛ��ꀔ|it���	�A+t�u��ق%�D�0a"1���n��9D�x&'�Rr���0O��Xaqޚ��	�3d�����;�4�<Y#��e��� �����H6�)���f;8�o�B�_��P"L.D�3� VxS'H�9=m(��ڑ5<93�8��h&�l��e���d�&��uѵ�m&FpQ��������aUSFkw�K�:����-"��;`A��-���_ɿq+����%Q���ЎXV�m��QV�f�&�I�2���2��6S*�/��,��PV�i;[�dh�ʇQF���65QVk�9M�(qQ?��ﴖ8Z}�qw��n��YՄ�B{�W�I�
�]�J}s=B��O
h�N�=�W?4��
�X�o�����8��d�0a�ڞ�WD�\�v��yw��;�1��|�u�dM��	�ʑ��P�՞D1���//281,�iv�1���l�&;t2��V��0���KN�>u��Ւ��ù:�C���� �]](�o��<�&-+��=Qb����{	�lrb�S} �@�"�`�k��~��n-����@{�5r���|���7ϓ Gy-��ՙ�� 10���E��;���y�G�$Y�CҞ�+֮;�^'3rD�4�/����z:��/�����@s��Π3���,����DF%�J��Nnڣ@Q�Je|��d�91e=�F){�uS����I���ߍ��A��wh� a�ގ����6����K,O��Z����MK���9'z4xt�9�>(B�����B����h9���,ej�6N�]�y>�9��S�Er�^��[����)!N��q3��`����9��SOI*B�d� �j��~܎u��@�`A[����ͨ��:o�K'�6��sRu�M�:$eNG0�FV}OZ��І�vzF�g�r�������k\ ½}�^~O׳uTċ$��*|�dTw)<8�KA\:7��{U���H��]o���8)�-{n[I��$��z*�Q�b8Ӻ�Q�@��8O�Zp��P �y౶���$�iȯU��n'O��DZ$���@o�5E�I�GcF���j�rK����o�բn�~���#��O
�kq*8���j����5�A|K?!���N �Z{2��]���tQ	�8FH� ���_�R��qġ`�i��7V�3�5�t9N�?rM�H1'�]�ctɂ�f�Qk~al.̙���H�0���O.x���
�kWݹ�G���p|?�Ej�v���\x_��Q(�
�XihI_Ұ�����E}�w
)�o�43ϝ�}٠s�� p7;l�@Ź��Ah,o�FM7#:�$�m�qD������р�H_�,y�:ѡ��7����A}������Gw���>����3�=Jgӷ@ Ԕ�0�H�rk\�E��^3�pŪ�o��xU�X�a�%��&���s����������W��Jr��jў�>:���I�rS�#�f~3���ޛ�t{:�}�v��L��6��V���W'�����������;�[/a���"C����b9�ȹ&�	��P�?�)O �paCt���Y�3c�/�/W�;ac�<k,���0#�l�� c?}) �H�+��s��;
�	�T�5�H��L�K#�bV���H��m�J��c��9E���'����YL���]������?k[p 0ѢG�"?qp�{�DSX�R��y@��\$P��MAӴ��
�ɑ�<����w���z��*��m�?Vk���Ŵ���xΏ��O�)��z����V��V;�='h�!Շc4��Q�%1�Z�(����C/
�(��}z�Y��㔰]�\�9�BM���[��
���Npo}E�B�v�O\|TNL�YW�k�k�
F�owe�:2�Jg�d�v��l�	Wk\��ũ˖J�D1��Q�T�d�\	�M��%dհ�^�P��}1��^v��29T��/QMMhJ�����;�����p������}&��!St]���h��_�y&?��=V=�:����	�FLr^I�S����rJ,�#�{� xi�R�n@��JrN�����v�#��?̌
�MV�?eK�:j��׃P7�t�\�Z�_��6тqU�^�F=�&�K�91ƙ�Ϸ���k���$	�s�S=t�0�&v�!>EQ8[@W(S��nޘ!!	�s^���/��ŊYN�I_�M�nQ�A����a����p�q�<I�!�F�?/MP~>]�[w�%7F'B�k�S��C�?8 \�M����4��vU~T'ٷ,�y�6��7�jhU�
4>���`��^�G5��a��!�Hyk�F�7�ӀQ�RV��f<F�$&��as�ʠ8b�}r�EZ�����ۯsW`�F>-�B��r�z�/��D3�KR����z�8��>"BU�f#��@��j�z�'�E܆��ڏ%�XB穧�&�T1%����D�;����⎏⫖ĥA~���Q�LHi��v�&�{�U�1w��TY|}�<�	my�f���E���.��ҏ�C5��:	�]�(sv�={D�|���.����ݣ@��_&��-)/G�{-�� ��X�;�/���U�N=������?v�\y��Z2�Ù�CU��Y�7'ذ�&C��/��'�+*⺄�Gy_�����"<��V]�>/@�*4I�u�ˋ����^	4ʘ<��,�5��M�-�m�[�^ө���	���N0�ەԱZ�;b����|Q��2�{�[0�����%���Q�#z�z�h�-5�������[�W,��p.��Y�0����J��;+jܴ���{��V���Y��db�4���.J4��د\�q�u
�p$�gޮ�y"����r��ʒ(B�aq�x2�"��r��I�c)6o�E�y#1_��]qAZG�r�*C%Q�3m�K�9�L�Ӝ�5�b��D�q
�/�,�XZ����;K�b�Ь����\\x3%#�xfjK�X�/�}ކ��	��I�~g��z-��)�%ֵ���h���M�;�~��8*���y������KĹ��cX��v$-����"\�P�Q��f�RP��߀-�������2����c�M8�47���z#ǍH��I���<X(wK�n��b%-���H�yH�;f�RzE�}:.�T`��Bs���p�sͱ���{[�|��.vW�?��@}1O_�5��2�)f�{D�_ �yJ��_���U_rɖ, ���.��O�s�y���1k	�P.?U�oPмV'/}�&z��/��"	�⑤EGѓ��U4�z��<)�]�/W��4@�U�����X�`	�LN�? <"�S�l���dMd�d�c�5����D4	CU�N�Z����Z�g-���sgʖ	�B{?˔��Y��E_��9nw�Z�m��TKh�J�5��=���k�T�������H�a�G�I���J�*�+!�׽_���Z�ɏ�Î>e��K3����Jݤ����t\u�����ǰFŞ&%��q��� ���;�(���qYg2jxQ����I�#6�yh�~��P{s_SB�q����WC|�jC�K��}L�A� ��^g[/p��X������CK�&�УZ��y��\Y�%��ff�5CX'i�}�z� t�I���h��a�k%�t�Tg8�Mx�rV��Kр�	�����b~�P�cϝ��}�-��d�9H#}��Qyb��	�b�vm��4y��ڱP�w�}q.�f�"��Kے�ݻ��I�{NB*W��wc�P/�f��|K��x�լ�
i����@a� _��n82J<ն���ex��G[�c����ي��u�RjVs��S�!���Սj��R���_�"^k�g>�6����mJ��,���!F9t�08�G�FgS FlÇ�����L�A$o�th�tz���y�},��W�/���ASǆ�$���͒� a��gZ��c���G��Rj]���(��g��lj�~�0�Km��,���v�6V��(6��M�Sֺ#�f��_�c2"����ߺ�/��,I �+C����]P� �_vL�R�Ӕ�3�9ܥh@�C�U�ܙ<�y2�!��`z~��tejQ�_�с^�n�f�M>�6C�~�K��J�ۦ>�£�pR�L�s�	Ut���&�+���8-bW:|Ā�)*!��ws0��A�����X�ۍ�M�o��S�l���/��$B4mqꐉ�sԑ�ѿ�M"1�o���&3��'���}%h�KL�?�2��m������4��#U���'�5z,H�y�p���_,<��f4��jٙݸ�0����qg���+��K4�F�U�Җ�R�E�8��6B��+ s�b��
�P��R����waeہ=`�T�-(g�L��L��h���^�,z{~��P"�B���#rDG��I[z�༇T �K�x��o�JYBg��R�iT�l��Jy���x�#����U�Ii<�׸� :��i��g*��j���A�7_."^������W-
i�E{��X�;2�-��QVC��D=����q���X"'��P�N��DCC� Ȯ���5�T��u��^���P�]�uztk�$*�A'C�J�Y������E����k�~�O�����vx�o[����K3���T[��b�/�%~��-������IK^����Ѧ�͒c�����ը����u\[6^&�׿���х@�C����c"�M�[kŬ�3{^B!C���p���)V���AOYP�?�tre0�V�T���'M���Nȸl�����J>�Ʃm�^'��p�z��J�3�W���V�&y_�%t�3�!Sw���$~ymè}�l�X��l��_�qd���.��j�x9�n�m�HlFэW@�T`�Z?���P�'�#9���~5��AH��m%W�!��0Ȩ=5]��9���I;iU���(4+��פ� �B�8)��h��
�r&��U���S�v��UU�C�>�ۨ�?�̱L���4H� �w�)���9��r>���#��P��o�A!�u�9���A� �<�]�����e����]�+�Ͻ���*5?�@���h����e�/j*��7��6?��?a��k/����[W�p�ŪZ���%L{��m�C�?�3�D�
ё���5�>+���p
L��v�QbM��ҿ��0�������g
^�O��j�<�o��콾�����<���)R���k� �
��_���l�$xѱE9��k�ԣ`�& {T(%�@+���Y�6��ZP��;>�m��N��*�ɰ�c�ϧ��(J�Z������l���Q�������{��gm��_w�����86���8A�B+�l���0YFtEFm#�%|et<;�o��Ɓ�j�ƺ So^�ҿ �[�>�\�zJB���e �?Q�^h��	$�.[�\2��Qv���l��Q5ɤ]vҚh:l���P��7�oY�c��x��
�5����U��q���'�4M쐘P~���s'?�����s�b*�=P�qH]���a�L����z�ҧ�U��$�&��)��^�Í��v'���� ��,��.��C��Y�:h*�ΏMĉ�v�.0[Mg.�Tw��K6f��%qXBp��H{�@G�Ԩ ����޴���i�Y��S�b���s��*'�y����b ��o�O�n��w�ڷ�V��*OY�7�s<��ے�G�)D�<&�w�d4|<_��'m���Q��A�Do)"P���(��ނP*?��|Q�?�O�5#�Z��ȂZ+�, ���Y	���,�@���8�%����+�=���P�}k��<A�P�b=F�8	`]3�Y��V])�
~�:�so��w���Z}��Od�pd��ٺ`�o�J������4C��I�hY�3J � ��03���=��w�9ﯱOp�DN��MB�a����S�O$�o�����ڛ�m�A��ǀ�j:��]�M$��g١�����%�mR��V�}��(���Xҙuz̛r�!,�գ�b�!8�Vo��;]~�h`pe��P����QXģ{`s(�����������}�Uɾp����Ն�kB�������
{�뾐�}�HBhsDO��N��/W�r�؎�
��"o��k1ٰ���AdMqR����W�j�\TY�;IB�E1/ ��0
d�{	���;�S� HG�vr1�1n[�v7&0���m�^Q3ޖ�s���w��Ed	��-q{nyFZ`��΅ρ���nQ ���E`���Ŋ-���ts��n{���Q�ge|y��[���w1}�U���6<��6��d��8_ Z���4_�n��J��+2�꽐�o���X�w�9�������r��JηK���\L��=湤8���/�o�A5��w:��Ư�(
}
q�D02�2A�:�I���67^"����AP9_d�kq	��:W�C�d����tK���L{ϩ��5��R�9�~/���X"�~�OLXKhM��tW/�jl�\$�c%븳f233X��}��_�ѻIu
C�Yz�r��%�,W�%5�� ��������`�貉%�پā8`c �h�V-L1<����Nl�Qjt�~m٧g󚅹hRa������!�}B/�f�=)�\TY�W�핒��y�*苐�(/x�!q�fq�K��yx&�[+��	��a$��ɖu8� Ɠ ������${δ��g��b�Rd���2�_`�"�t��+6R��_v�9^��g�";�ݧ��[ �,'2��rK�t�*��=�gp�l���}����JSA5Ē���t��O�V��p �ȸ�/�.�A�~ǆ��\Tk�D�Kc�8"��T�|��G��l �eу(a$��ha�1���lm�(�,%��>6��	(�#lM�������\��PcC$k��#����Wǝ]Ƽ�>ϐ��P��2�P[��c"��<��35G�^���}�ύ���J�\!��`����2�<jj��������Xn;�eM�64aH���\�i�$�9�{;����p�ke���6�QL���HQ�qg�^�(a�1��ܽ�p֥���&���u]�8�	�z�V���+�l"��́(���sX]���]f�T"5��/5�!.A'�7�5̸�F[�[��O�������gD�KeA��7�0Q<q�o���)�������҄:�D8��C�	����ׄ��(�IVV�����bMߊ�4��2c�k ���j���� ��s��_��A�#���pN�=x���=s�� �ܙ��uL�88>��e����R�A3�.��s�����ٗ<�ݖ5l�#� z��R�`s����d��
�1��jD�ڟ�H�NS�W5�0��_y}r,:ìxRQי>nޚ��l[��g�b2y�-��;�KJĵ��!�Sn�>T���=�}�<T�7%��`�I֘�S�*l؜�饓��dn~�-vr�n�`Yd�����ӨQ%9�
�2�D�-�$@� =��I���T���-���W��%�w�k/F�8�5j�1�v���Y+u���Z���	�uW�^�<�/�/煊@n���j6�:/&���y��2X���H�� anB��S��7�YT����X�iڸ��@K�@[�B��fZ��{́������j�H�Z��˺�"~:�%���B�Z���g���fn��ov�d�&�"�����4�Ӟ��|�۝& Eo|t�[�n�� ��I��6
t>|�l!�b�a�g��e��AI�7_ήI_��K�.
Ț�!?#1|�$8_1�U���Ř��w*�0�*��N��#B�ͨ��uZ�4�q����	>�lL0t�U�-��:!�h�a�kut��;zm¾��β���G��X%�ފ�M��h^�7��;�����S�^��B^�j�)"M�h��ñ��rN�o�5Z�����v�[U�N>�4�g-ֱtQ��ݩ�(������0��;>١�#:�P�Roԑ���93�+����(�3݅�x��de�%��wјS�+��&�*]&k�h�E���5Mte	k)*9)O7�v�6g"�?��y�����$�tWƎ�퍖���L�Dxm�5�?�j�D�&A�E%,�]�&S�ژ��L���y�{������m����'����^@W��e�j������*���b�d���Q-u� P|�����x6�Ea�%��Q�+Wb��� �A�%��&Zu�^s�Zx;;f��F�Q�#����E^��؜�:(rt�Z�y@��E�c�\�!aA�vP�PtiS��QZ�:� ��X��/U�|A�@��&V� ��{����d.��t&��n��ea���(�U���+�����m!M�,��G���67R�(7�Mt��d�b�Q���_c�jb�X<ۺz$;�-�e�L��� �KP�Ȃ��������=v3�˳ܦj�dy� ��ڀ�!��`���2�j��j�`^��Wn˝M�+X6��3�-۴���{�1�{���������N%�68F[Bj�H��gpɀ��p1�1|�l�- 	��\O�]�]K!��ś�_R0�;���Zi?�?�h�\{	�P�[��q^��	S�l��k5�òv7�h?P��/���|�Y����\=�:�5��C����v���a^y� �}� �H�\'d��D�sE�
/31=��_�+�{��a9��ː��z�n��<Q)K��O&��ݭ�f�v�\��O����.2EY��H:� ��]��n\�v`a�[rꉈ_����� hq��r��F�H`|��.����J��{|�Q�n���K��b&���X?�*�P��7���[b���o��n�L�w

�;ES*�c�\;�<J���JɄ.�ȥ�2�w/}|!)ɬs���EQh��U#O�_)$8���dJ�m?��Qǝ���#�PH�m9�+]��,�_ޣ�}�"[/����us8�>�١r�+�=��YB}�S<f�@i�'Fl08l\]�J��?��)�(���b�s�1<�ʿh��.�;���~`j�_��f�ĝd��|�C��2W>�E��-�7b�1��pp�� ��{�z_Q!�g�v�h�M~���]�?F�(��_����Z��4|
��x�c�˾�FW+CWYXfJw�����A��ړ�fa���勎�n4�m~�C�.Uɠr��2ɓ��U���B2�ۄ׷m9?�2j��?5>��MG}���?��:��_��6�uث��\T}��u
�:Gr��L�J���Bؼ�!���f
T/���<�����z}R�Sx��!�������m�Iw�ea%UMתg�J��Nm1�w�8�F>�9OB2@�n�Nb<Ug�%�� `����\�ki}�E�O�w�T�����:�Lo)$���\"I�q����>����E5t�:)��nC&P�z���; 䥶9ߍ�s#B�B�L��Yz[b��'�����QAqUޑ_���,
����(�|5-;�/�Y��j��K�V��W�H�VU��9���>��S=�8�D�jmQ���|3��	!�gh��Bҵ������%	��H��'��G�R��dĉ�"iŐwV��/5���!�i��)�ϊ,,+`��������(즄�S�!悉��<�m���,��4���6ҏ�(2Mz��:�}R<�[Ȝc�0>���/���(��Ƨ/H��J$P8��[���i֔�i3`�ܡ�
���q��Q����o!O3`����Ij�f��[�#���n�Z�M�|6?���>�4Z>���{����jy���|�id#6�h�� H�gɐ��1,�'��3)�׼�8,C]��~�4gb���ڵ�+"I�i��d�~%w�>2d]1�"`t�/�&!.,ӻ7�^�v���f?�OG�����v����D!��e,�T7�t<l����V�Rk~ү�ID���.���g�K��U@�5!�P5P�V�Vτ��E<b8�:�ih�_�}�v9h�M�g�Y�&��o���'�,t+��p�p��k=�.��P�
ūc;6�� n�#�(�� 陦xR�c3?���>^��o��&� z]�n�� %�GR�*m�/�
d��-5uU�B���*�;y������b��0'�pyH�f::�?���`Q�Zn>���G�qf:}g	�,yO���AÈK�Qg��`�S���T�w������9��c7P3M`�����
S�a��G������d�u�-AWknI��`��݅�����%�Qз��h��7�-��>�D��>�D���W`{&�CD���C��3��\kG�dp2�5Uݽ���>=Y6<��g��ᕪq�4Z��ƹ'q��z�u�5 �n!M��1N�ᄋ�&$Y.���2�)�b??���/nMLS��ƀ$@h��ȩbi�t��$"@_*��ѳp�FT]��9ȏ�B�_�Zew��v8p"�mM�{��d�Z�Vcg&Y�fYR�o���ј�")*ՇP�r4�|����W|?(+���o^��t/ς�yۢ tIS(�
���|��8!̪P�*,�T'�L�7��I*`�v�X��;��$-#|ܧ$�ȫ�`\P�~ET��Uf|01W��9��#�XQ�4�tu%��4:-����>�'0�	IU�b�N�}!�Ȩ�l �k�j��>���[��}��Ν��ג]�X�l���}<Ĝ�;��Q�~�d>����O=)-X�h82α��jry�����ω��vM�aUb�>���ԏ�?��8k������[��)-t���e�G�ō���S�� �!���f�f��` r�E�����4�핻���&������:�j�3�����[�O���=M
پ���6������%C-�4��u�l��p�b��dC����p�a��f���ˣ�f�0*�hb���Ǹ/1t-MB�<��իݙ�.��7�ǯ&��@������JW��YDna�,/N|��-li�-�0w��P�-��n-[�ڕ
Tc���d�Q$����u(�PHG�A�pq���$�c�+��0����t�!D=,|�~�^vp�m�p��Ca%�6�e쫈c�=�K���>:%fVBcIc�����Ԟ�/q����ʇ{���$ڬEF�P(�.)"iMu-�`�Q�f���?$&^�(C���I��v�~Ht��:Z���6��'�3(�B:˕�P�1[j~�8�c� �_�ۯ�O���ly�fy�κ�P�qq����O%��u�樄\�ސ��	#j�gJ�+32ྉ��ɥh4j�Źw���v�dB$e �?2��d��8�D(r�㖋c��$��b�zF�2��q�cY��|v��11-�a/�_�x����mG3�Y�V�c!+3tڪ�Ξ3�N4��1��ŗ����LGkRJ@��`��30�,�9�ą̫"D���gX�N+��@�~�ey�B�_1����#VC{yw��ݰ����<z)�>���U�wh�kp��a��1�ͬ��RK�%�MT��:P����Jj�9�Px����[�����������:m�0��e�/�N�Jc����*��������F[������[�N�P�3H�`��\ߨ't�I�UL�� 8�L�������u�Ć��g���ͥ��:�g ��3����㙂�u�L=:�G�Gdj�FS��O�����Wg�g:�����-�\]	:}둃OtF!TrB���V�ὧ)Y�u�`2\����[h��9�E�:��tN�)�Zns����z'a�R��u�϶.y����w��������7��B=C��u+U�P`�?��aZ������5B����)��:j���K*��݌U��+d�����������8��jbZ�ϲ�|h��ށ������W���m���'�	{4sHB�O���R{�9���iڿ=V��5T��@�d�ee�oWc�x�cg�kz�lkK���90���O�R�x&ў�R�k�$��� ��~W�|�?E����RGx��L�N�
~��i�q�ҍ̛�*�E�� 
��O�?��_D�������7��M�]-ƃ��,̃M4Z���$�oXqލ,�4����8W,֯iў���!_��0��aq��t�k�*�>�"�ː��J�:�T	i�ѐ��%"k���bek��M�����l&�k�X�*�%����D�����"]�K�,���r�R���w�:���($���rscz��~0?�{K���:Ɉ˟��4L���Pq�+�q������7�ĥ.ٱ��S�oa��C" [̔2�9���&�S������O��Wa`Dv�o-73��,�;���<��������� ��$�@6H���p]m;��D��4͍%�9L=f�"TpVG5�HKUm�[�� ��9��>���{�SH�ڪ�T�a�������p]a!�$y�呴�ÔS�����=p5����:+�A��P���ɮRi�j���)H�w�E���mļVHn+�5������/�_N���5��ɤ��V��4;j9�h�2� ��l�Q�*���(���� �䴥�}��
�im���<�X�B�6��r|
������}b�
B�bO�<lNI�iW��t�[*
��Ho��^��}�d:D��i(�W���\!�ʈ�#�1ܞ��D׈d�6�	�s��hC��L��:>��1IAv��bo ���<�����_\p�ZEt�
���̛d���ue�?�^�,]���~�x�|�b&�����=�g��C�%��/\YO(�9<�B�&[0�%�O���x�����kk��Ѣm�k#�|IebE�4��(4x)��[eq
+7di��`�z5U��AE��
�E�p"=�DW7��)�����7(W��b5�M�W,9�MA���$�q�0l��h��B�ҏ�,Ckѫ�þ�������N���8*�W��>Z�*��PJ����|���	kf>B��1P��7��:[)�y]�,X ��%�%/�Ѫ��I+��a�Bด�؈Wr4��(�]:~��(�D9rݾ���[~=�I�( V�":�<���0^L�f��_���k&��;��]$���ٞ���]�a@&"͠���1�9࿴&C����	[O*E�a�ax�<�|3-�9�z;��<����mw�v�] ������HR�*�}Ċ;T��ޒ���LʋQO+YV�H���m��ڭ�49�H>��݃�2���w������c1��3p����fI����T�S���g$J��N���A���������M�79�A� ���t�]ml�V5
'�­�2�Q���������x�;�V���;���h:���0��tHQ�l_�U�x(*���l�2�t}��߾6��'�g� �PB�T4��4
�^��X��}���B�G�O&^WNV��W[�بpw
���o���̍��!�d��7�v40W`:b\n㡩�w��>�1	;����di��	�<����:�ξ�Zv�J1H·vQh�ܘ{�dN���M�LC��	[�7m���E�!ٹָ�J萫 �]y<��m���&���G=�g9���,	l�3r(҅StH�\n����ȷ휡�
K���@G�r���)!/��l�#7�|�V&��N����P���Y��ZPA '��N�Z\�� �q��^'�E=yy&ܘo�Ck�Ͱ�ރ'k[>��.�osG�Atp�&@�H��8���W�G��8d�!+Hhs�Ĝ���-�T���SwM��/�ˀ,�V�)�����qbP��낎�I=gM�]z�m�%QR7����RyM��v}�&���"zI}R4�aȔ�z16%��'�1�ƍG���Ţh�hX����[���ĉk�c(��p�-T���HV��Qruϐ"�3ٯ"���յZ����&�� _}J�f���dV�����9����*�Qֳ0�v�)�Ufyu<K���x.���cW��j�a,	��ѥ�8��΄�����wtμ��o���j��R#����3��؝�*Ja���R8o_~a^�eg�A������Yc"s,/���z�t%^��#+g�l�U��/����A=�7��5t���҅r�x9���1/�`sA��
��ad�W�L���@���\y�����g��m-�(i)�p�Q�p��	�tm�I�,-Q6���6���(��1M��Z�ܔ��	�X��cK� ��.J��e�ǥJ[��s:Ϙ_P��I�X���ktW�D(3=�ӽ�   �  v  �  �  �%  �.  K5  �;  �A  H  aN  �T  �Z  *a  ng  �m  �s  2z  t�  ��  ��  >�  ��  ğ  �  ͭ  �  ��  h�  ��  &�  ��  ��  @�  H�   Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�� |d��"O
`�(�;���8���-0��1%"Oj4��ND^[��"3/9�0|H�"OB���H��*�ʞRy=a"O�味V�!X��!&F�:J�$���"O,��a
���C�Ą�M�"O,$3%o�-���p���+Ն�:1"O��ݢ1����`���y14]2��i�<�6��{_���c�H�`�fX�$Kn�<��A̼VI�xR[�)�Ć�pඤ�ȓA5��('nߡ4�� �)˩%� ���,��r�؊b#`T�eT09���ȓ!�b��g��}�8�F��-? �ȓ
K|m�ș�VṔ���2�%�ȓ"R�X�j�4JN�1�˘X�i����̹	_�jZ��1!g��zܶ��ȓgil,*�J�
j�Ne��i�J%b���f	�(U��:���G��$Y^م�~r�� S�%T"���k\�jx�ȓ|4�1�îJb��@ӵ�ݩn�V��/[`�"�v4�R�!ʎ<��M�ȓ`:��z�ؚh�J�Z��$HY:	��H��p�m�C1��!��B:��0��EnjZA V;9����J[
2���	��4'J�EA�IVW&��~�(aZ��ӹ�>� o�Y�|�ȓ�f�A�
Ο7�H��M�$�����mޠP����/���ANXo*�ȓTv�����{ ��-7�*h��I��sB�8�8���3����ȓNe*M�悡;������X�o��!�ȓ'lj�#F�m�+R&;�|��2)n�C��0S4���T:
b���:�0!��e֊��)��ͷV��,�ȓ0�&�8#���� ع�L�����;�P�AFd���,w�6d��r�EQ�( �gVlɦ�M,H��,DP���|�I	$G#\���ȓ"�)���E�B	yt&B�^�LɅ��|��B�,�r�Ռu3�h�C��'8!�D_��p-���K$��aU�/ �O@�	i�OOx�h��	:T�)�"��,n:�;�'�ś ֬y0<�Ɂ�މu\�	)�'C �8�:\[B��@�׵olV��
�'(��#t.\Q֕����c3��q�'�F|#�άt1�@+ 
�-W�Ɉ�'�|�Q��I�A��A�Q	5�d��'EXհ��IB�k�	K�PV�%I��hO�!�s+�'\�F���ز=����"O�Pr��� +�Q[2�[�_�� ��"Ov4�m�?Vd݆p:D�D"O�3��S�( ���1qZ��Q�>yG�'�j�AF�O��4���E�5�t��'Q��4hV�0i�tK��*��m:�'�K�N2��F!�9��hê�\����?�'%��)&Β�C´�;@�C%IK�a�ȓ`��s���8!m��Ks�%�t�Ў��s���Ū�1|_��z�%�"e:"���4D����Ƣ]!.�c׋X
[��Zu�����xbB�6����MT��
�� ؏�y2�*=2D�w���2��5�*��y�?@��2�r@@0�X6�y
� �E��U�x��\z��P+E<b�"O�0�䌆�n[�!�� �Tx��d&LO���h��Ԩx��E-�BG"O�D�������Mb��XL1�"O�	�F��;(�bhc�-��H \�"On%a��Y�l�{$���BS�"O�ఢ#̷F�0 �G+�VX�"O^���Æ�u�n���Ɉ: @�I�"Ot�!�'BR��F^�P:� ��"O�x�ь�(v(���{6���"OLH���Ti��a�dU*'�'�!���kP���^\��'� L�!��[5	�V����:GPƠ��e�Q�!��$
�
�"�Zi<`�G��.'�!�d)Bà4�cD����<!��� �!��1E)�)�ի�':昌�̘#o�!�dN�|4X�����W�M3��k�!�$��DX����-���VK��?�!���X���`# I���_#+�!�d�)%_�ʆ�f

*�P�2C!�$Yh�|\�`��� �Z����=!�ı�n�7F�0{�xu��M�<a:!��* �6Ҳ�]:�x4��!!k�!�DDL��y���Xl�Q��ͯYta}�>Q <hwR�X�%Ym|,[�NA�<��FT�(�� �J>v:Ț�LM~�<�"�N{\!J�#;5>&�$�Iw�<�GZ�F�Dzgჹ(�v!�t�p�<�Aj��e��,9��5}:�d��h�<y'l�]&
�1$�q�i9���c}
���hO��b��1^h@SV��>3��g�'�MP�0A2MB�Ni�����1KF���>��`���j���|6��s/�30�	��J�0H����+����glΕz�"̇ȓm�2\��L�x��\YwKő2OZ��<y���	 7��L���
u����a�k�!�$�g��e`	�9�i�� �n�➟����锅0�t�:c̊@����2���C3!�$�� �~��T+�6��uH7&��Q��/e���N��V�n5� ��)MZ�͇ȓ]�.��M�������@�IM�����z�E,f���9R��.9��s��)�}�Gԛ���$.3����C�y��	@lY��d%-V&Y����y"ݛVd&�������TPg���y���%mB�`��GS z%�uK@ȅ��y�葎�=��L��C#Ԣ�>�yB��l�|���i��?Ĺimޛ�ybo�o�d�Q���+:b|<�U���$�O��"}�E�VWB�ု�.��� ,@a�<�'jަF�7�ս}S֙j'.y���=��� d�ZP��n�9/�Vi*�SL�<1�鐡S�ʨ��E9��T2 ��|�<I�i^�%�>@ ��3o8��e(�w���?Y�W7U����)Ӳ!Z����z�<�G��U��j�L5NH��2T�,����N�����Z#�$[$�9D��s�ʑ8n�
-�Y-����/"�Iz���)�[x
@H���EA��d"D�x*螙HU���'^�Q�ƜR�o>D��[5H�q��iR��-��ibi/O"=Q6��\�y��bԺMw�հq�u�<		C\�z�WO�/��A�5��h��hO1�^0�"\>�T�'�
$��"O�  =�r��xN�1���>�1��IyX���q��<6�B}Cw�"tM��Q*:D�D"6�_m/t!�b�#��>D�����P
����uB7���O;\O<c��W�;t�ZMU���4��2�h9D��2��N*O��t��KԵhɶ	"��7�	]���'b�6y(6�mwJ����ߵ1�lX��*L=��ʂ�W�����k�1m ���6�\h�S���k�Q�%�)i�!�ȓ/����l�r����3��0cI���O',S����V/j���ɭ  �P�ȓG�H�FÙ�M�D�׀�2����>߰��,�TJ�I�w�[�v1D��<�����ӻ-����'�ۆ�>t��'Q�E�!���DfNd�W@�y��ђ�!�e_!�dR�^����;p� �@c�0P�!򄆗e(� 
Ãٱ>�TBGb�	]�!�;n� b.�6�I+u��G!�@<�Xce�1!�dU��	�R4!�DVD�R�#�B�E������~|!���9_�$}aFOڵL�pϋ�s\!��ܯRT4�&����$:���ML!��G�-,�e��j�і^=�t�s2!��$���Zv(M+6�*�l�Y�!�U�yF�X{�E�(:"��9Gl�|!��-r�<ate���(F�$�!�d�'J�L�W)J8l�*ؑ��I�!�d�G�X��M�L��I��)�8Bt!�	�z�;�^�
�� Wd�0s�'���%�=-+ΐ��-�w[���'�Nq�g��^|�EG�&q�"�
�'�����J(pUd��g؞d,���'4�ЃRD�#kĞ��t�U#V��<P�'�V�D�	<`����K��0��'WJ�`@LW��p ���s�;�G�<��+��@6ё�&�+�f����F�<ɰ�=N�"�B�	rH(E�UA�f�<!��6W\��f��6vz�Ѥcw�<Y)I/V�*�ȒH��^dPE��k�<����U��C1��ҤX��Ag�<A��?B�^�#�w���g�a�<q�Y�.�����1PO^(�R��[�<�Fd	xQR����O,�8%Hb
X�<�)G^��!�R�|�G`}�<)#�9�l�l��bi\H�v�^y�<q�K��s2$�0�j�5�@L�1�XQ�<Y]yG� '�ܶii��4h�j%!�D�
� ( ���6	�C�ªg�!�Ć#H�Y�2F�
�E0`�dJ!�DP�=���Z��8~���5P�!�D� �,��t�*�����m�!�+�|2��P��uصP��!�D�2��I�H<L�Z,pwL��p!�d�E|T��CL�J̓%�Ƣq1!�;4*�����[���`�G	�01!�d92�8��F�JH4�;��WW:!�3b���O_�73N�K�S�s�!�D̵i���ku�ǩS(n���8+!�d˽]Z�D[햻p��Q���T�!�$�i�<��mι �\a�-D�m�!򤆫	Ǆ�C�C�(��QE-�0Wi!�dªc�0�[�9�fh�t�=!�dK�]'�麀���}�J�*c��`X!�d�l�����b�⼻��@�2?!�� X,����� 	��+�h@��"O ���rZ`��G����	�"O�!��Nױ{��E+^9LC�0�"O�u%�SUE�{�ކ(/�� "O�4��j�WE�|3�ǅ�j<�]8��'�B�'l��'��'ZR�'�'�Zl��R'$�\P��'2U"h���'d��'pr�'B�'�B�'Cb�'u�d���ԾvR����E�tp4(#�'#��'-B�'���'j��'F��'/��2-��i�V�+���;[����'�R�'0��'���'���'Qb�'��LY���r��gW�"�ՐC�'��'���'��'t�'��'x!��JܒH�
�#���fl\ ��'���':2�'�'�r�'l2�'��u�W��>&adCϋ%D@=#��'�2�'�'~��'�'N2�'�ܰ��T� �x���6Qr�\���'���';r�'(b�'b�'xR�'��X�OɨZ��!��A8f��9�'�'�2�''B�'K��'l��'�dJq ` �9oQ/\��(��'��'���'��'vr�'VB�'u(�J�d�"�U�$����'���'���'(2�'Rb�'R�'�^H�F�#��sސ0�t�'B�'��'0��'��'��'q����,�ѲQ�T��7N1U�'���'�"�'Bb�'o��b�����O�hru�D�N2��R���!�� *�fy��'��)�3?!Կiڭ��M��FCp���`d�4�S��	��禹�	I�i>�	ٟ��)"H(,��E�N/kG2�J�ERџt�I0r��oZO~9�xU��Q�)ی\�~�S1+p�c Ù[}1Or��<��	�>0����U��-L,13f�=d|�n0Q��c����U��y��I I,DX��D�vp�$�[p,�?a���y2T�b>}�����͓^)
�iƢٻlR��U��"X�yϓ�y��O,���4�x�dT�� �#B�.�pA�d�[���$�<�M>y4�izv�яyB$u5n��W��!z��	���IE�O�@�'uR�'o�D�|�4!�?&w�Q�A�P�`�qW`/?���B������W̧B������?Q�b��-����� �DOv"�g�����<)�S��yb�^@�z�"�8N6�)�S 7�y"`~�<Dxe��l�ߴ�����j�?7��$)���@0MS�'�y��'o��'+ni��iJ�	�|���O��\��ׁ�hyZbY&~�Ԭ�aH/D�`�c���\�H s�l�t��);D���FnI�f�Xy��KAw�(sQd�o���&�<D�7��5Y��Y�o�w����IDc?ƈ3�f�s��d+��	ou6-��AH�`�R��@G_�\5�IQ�މnq�T�&��h��j�C-�MHWDM�t���EX�@�逤d�}�nX�!+еP��d�l�s=&�	Dlɪ �����	5x�iB� Vg��)ɞ"�C�I�:���� g�a�V���
�b�ɃK\-crePe��d풀� ���*��e�q�QK�`藭�X	H�*,�,)m+!d��Q�q�Z��ˉIx}f�H+�A *�,���*zj� i��yycT�
�`>����,3��%"�N�\�@�4&@US~�3�/Y�'K(� �/AןL���4�	4�u�'^2Ň"M~��30#��#u=S˞�C=�����O?:(��K���;C�"���O&�����Y̓�p�a1W$d���H���s�L'��BC�5��=���mB��֘~r`��>u��D�L�b���Gʮ'�� ��Uu����<SR�'(b�ħ|j��
�~b�� �,p��Yi��Vi�<!u�^,YX�:��'R�ʠ
�L�-����S֟|�'��t���l��``lD*�jɻg�0T�^����Or�d�Of�d�������O��e�h��C���<%�T���f�!�
C�dɢ�型|1]�"�'x�e��LH��	7��D>�mwĆy�2�0��D4�(0w�q(�8�t)��'�i�=��C�ӟx�	/�y[�Ƅ,d�T�cE�N�d1�Iw��h����(���X�+Y{n�EC��+V�!��#V���e'�j��x$"�a���W�����C�S�O2Xuz�\��ĀB��0j�p�'9&,��U��ճT�ø�JD��'/ 0��lW�#㐅�3��0pt��
�'�΄�T]!E�F�r[�S,�̃	�'_4��#Oǈ䶝��b��@X�	�'[�E���]=(�.�.ԄeQ#���y��ˎVA��aR#�=-�u���y�#F���c�M1#Դp#��;�yB)�Q�,��u���z�a�E�(�yb+V	��&�Ҝ^�t�Ō��y��@�ĥ���=P�\|���Τ�yb	_�ʥ���67Dh\B��.�y"g 7�� �ʞ+2}K����y���z�D&�83pڱa ���y
� 4�p)ߐ/��xR$��; rt(C"O`y��'7v����lɱB�j��2"O��A,O�x�K��7c�ذ�"O��F@@�X�a��$��ju�v"O�0�F4̞	��E�,��"O� b�/N�>�hbC�/,���f"Oh 9`�Ơ��ʒA�-,�j)ʓ"O�1RB,N?�h�2�!��%N\u�"O �I�'#�i����ي�"O>�i!F\�V@|�".�4P�"OV�F��8�l��/��G"O�tz�E�> �s�ēA%tDIV"O>!��HݹQ�����Ⱥ`ī�$"OHJRKRA�t`S&A�7u* <��"O�m�ċ�.�<�:�ʙ�t�%�"O�d�2h�+'����JN�0&�R�O��W�׋(��;6�V�V�
�K5�F�<�6��=%�1�E��4ӆ����NE�'���j�(�S-0��U�C��u����cX���B䉪C˞؈�۰+˜�������8\�\�>��<E�I޺Q����!\� ]�Ê�.�y�iT�H��h���َ���Fh��]F�p5O��j��^!-6��I?�4��)V�uۊ����˒=�`�Ӑ.!�O�hJ���1HP��# �tLX�p�#~/J)�`�%~��IÌ�jX��z�MV-2x32��!2@��`�(�o��H��U&/�F��5L(Y���
Z�"UA�a
Y��RB��"C\Lا�	`4�H3�F9�%1O&�QA�Z�a�����a��M�?qY�OQ4 'zyH�GK�P��0Sd3D��3jG�s��1���Y7��؇�s!v:3��J��t��=H8ʧ�OxD�"%�*���*Cc3w�c�'ni)��HҤh'oL(09.qQC*�e�@�� ��6rƅ ��7u$���d�2�A�Ƙ.	aКǩ� Cl��`�h9>�[gD��p�h��Pap���܃ _���bA@�LG�i@�a�iL!�$�s�� 	�G�A�B�9ǟ�`2"��p�DL &Խc���"+�1����)
���,���
�#X�S{� ��#D�09�M[�>h ȿ��%i�e�s��%��4m�����d�M��Or���gՠ<����_rb�LAd�'�!��kNl!2q�X���Tmޢ*��x"�Sǰ@�Q�.�O��(����nj<5B�ɒp8�U�A�	]E���E����![ט��	A���1�A@'��9�Q�H�!򄇚$FĠ�G����!	� %�dT,:>z�KaO�^�R&��z�O
,���u�-SȜ�5[0x�'��``S�V�n��(�D�@�̩�ƥ&vj6��S��i���US�3�8����L�S����/�����I�2�`t��\A��!�:f����1v:J����:�����I�s�$���jT��~�3�0XB�=	���	��&U���ORjiaaӞP.���E��	K��J�'#�����Աh���!���#q ޡ2޴{���8ň�y�4yy(O?7� �E��<�ڳd�h�3-ͺ-�!�E�2�8�۲��!>	�x�s� nA�ɶ5��K��#lO�B'��d.�U@զ��F	���'������<h���`9J�`���
P�`�'D�� N�wU
�1 %G1u0@�.3�7\���I��v2��0�ݤM7:u괏��	h!�$K�J$�H� �0)r%�;lb�V��<S�c�"~nZ�4V�B��7Lx�7eM�C�I��	ɂ�y����gްZ����8�A� 6|O����HZ>J^5Zb��,���;Q�'����s��M��l��2稉V�P6~�ҩ��VS�<�'!S���������l��Q�'Ȍ�!C)O�Q>�X fɒ:^��h���h���
*D��AH�tT8�zr/ϊkJ��Hq��Ot�IC�C�gw�O?�8ccN[_։ғH4W�l1�DZ(<�5/4W�d��I�?��0��ڮb��@�OX	d �U��� �@c��V8I�i��#W�JU�1���'7°J�F#?��,6����.�,p~�a�V>x�8��V"O�y�D��Df���!J�,7�)���CMS���$�s�0G�����Y�d��$��+>������yb�E�'���W��v�2�rg�����̟*U��i��k���~�<�r�rM ಶ��8Q|r��ōY<�v�<$`�u)�䈈P��	V`ĺAN
dA^�Lx .H�Qkaz�@!7vz���EI�j���bW`���0<�׫�=m����^�Tp�  0���	[1f�Y	W���y���
|%���qB8/���V�����(0���'��&��B�~ڕ�uU���Ɵ�(���6�H�<Y拖�*� ���ŋ�2����O}i�?�^}j�'n|c>7-)q��S(�"x��k�D�.40$g�;V7fB�IG`"�{��Rr����*HFu�V\�FH~Ӹ-�$吪A�R�Sa�|�?�A��2� q%�c0�!��EL�\�I����X�V�xс ��p,vd�'��Rx�$C�@�P	�jW�92|�#Q�'��t0�U�7�,ф��:;�H*(O�Yi�L��?�&�v��Eb[���g���d�I���3P�Jp@m8�	��yr�Ӫ`���9�ؖ&�F��<{W>�£��S_��9v�T?mkd�� ,��}޹���
�$i.T(�� ��w����dLW�US��� &S���Pc�}�P�J���Ц��'�jm��'
�)pt��{�1���-{JZ	3r�R��=����/��-E~�B��s����ɽ-�~p�bf��MAD�	^�{%�[?j�@C��P����(��r���)���r/B/��AJW�wNj�8�z��5Oz�qVK�4��	 \$t�i>鲑�Rsግ��m����Qk��$D�<9D�_������ѵJ�l0��oͳD���E�'o��q���~z��J��9��I��ɥg�*���� �x����'��Y���!�${�g7���:e�_�!���.��O�<�ቹ,ňA��V�xe���|�#?)BZ}��$S�NP���O��l*$��2���ȶFv���b�O�����'�y��ua���ӄn��|��OH�	'ȵo&u3��۵BC���4�`42d�ܲ";���g�X�v`�ia�"O��Ģ����>����ra����a�:��Ѥ�^�m��T?O�Β�O �ػЭ!��8(�MNu}a���=@�RӄYi��ڒ"�1ְ� Su͘扈��'��<���>��a��{1&���+�q����3dD�-;��݉5)�Y��1�X@�%f�	b�4уE+?���Oą��I�|�.�#3��_B:�8d�R8qM�ż����[i&(^^�O�����߶\�DP dfE����'�!`�H@�n�()%+Y��#"6
d�I1�MS�*����gܓ@Rܹe�%R��T+�	�ȓ2V�T2��;b}�=h+A�:�R�mڹ
�<�sC�P8��c�
%F\���@�_�4x�pb*(|O��J�G+g&�牆�
�B �����X%H��~B�	"�B�j���Xc@�}�l����'�-n�\�F�d�K��]��
�f���K�r3�'P��{a͙�k�5fN�[)���H�WV���J<!��>!pD@��||��X ��$h �OL�<�E ��ij,e��$��D8���KRȦa�7E��l��e	�J�Q�D^�"E�,�ĮW�a"`����"	lz�"
��<5�ːy�(�k ��<�0�,�O�<���k�Tu�#��Gs�ӑ�s�'p�H��d7���P��D2~4�⡯��j_,�ȓz!�0i�.�v����&��}�nZ5f�ބ2�}���i�v�ä��{��逽���3"O0-�I�.���tI��M"��I�]��r5���0>��ˁ�Pl�f�n]�ᯈ|X� ���G!�y��<z⼹��݁|����lY�yb��>*U2�K	n����!�HO���`>�h��RP�4�H��f�[P��$h�"O����da��V���=z �iþ�B����������O�e�څRF��.@����/��yc��r�t��/�Pв�X��Z���Ę�����'l�S�m�1�zaÁfWE���
�lJn|2���O� �x��aO\�<1�桒�+x� �B"O�e�1�[+x�ļp���Bo�2�鉁m	2���i�"m�\d��K�|��	�!K�N'!�S)�ƴSQA�	�����M��&	ͨ�*c�"~n�m�������=V����PHL�C䉉{�d�d�B�"�ġi��=���Sֺ���'��w�D����3!a@�@eU�� AJ5�7O�S$��-��PSĴk&eAS"O\9�G�"QP���&AT�Z��ɢnŠ���U�z��<���,b� ��U
(�!�d7PK$E6mD�Q3�\�_����O?HWIZ�^�x蓅�)ց�pR�<��G��8�ޠ���B�&��H�z�<	�!��8��I�̲li^��3J�a�<�4��1]&-À/�J��jK�_�<�ƠY�L��)���**��M��ÞY�<��b�2��!�M�|�Pi�-J�<��M�]�Ē�g�D�\���nB!��P�C"}ȀH�$	>�K�*��0!�d�I&x@��M���2!	I�!��Q�q��I�d�A�}�ܭBWH��]!���&=�W�]�� �h6�
��!���

A(@O	t�hu�R6!�!�ā�oa�~�PLӾ^K�9�"O`1�u�Y:^��4����|J��r4"O]K3-��RAL�Q4�2 ��(Ӥ"O>�9�펊_��l�F"\.8���J�"O"U ��]�	S�#v !K���K�"O<́�b�&D�`�"�ٽg� ��"O��Տ��z��h�BκR|N�#�"Ox,���D;(���с�� |��"O��0�X�S����� ¼f���q"OzH�����*G���oהR�:=�u"O�I�wCP�l�a�D�B�湑�"O�%����v)��;e�_�����R"O(��g$+u!|�֬ԔK^�;�"OD��ÃǿI,Th��쑳cYl��q"O �@"�d��t���Y�X"�"OHX�#dQ�E����3d��Q�,�$"O�i�W��K̔DbvB[���L��"O$�HǍ E^�{�!�P�����"O\����rg�B!J���-�t"O�ء2��01���o��[��p�"O$<2a�J�L�p0�o�2n��(�D"O8 s�LG������B�>�;C"O���V��G(ܙ;wK�H�T0�"O�(�0l�Z�Dк%c��n�xV"O\,�t��,$����b҄q�J�f"Oʈ�%�8:���c�����taxd"O���0�ǀ7��T��CҏQd�c"O ���9S'̹:a(�jl>���"O��ܬ]vd���=
,�`"O�����O.4}�ɱǅs�|��"O(,;1C���%pD�/gHqV"O��@w�Y�p���$6_��ra"O�����M(a��M�N0��q"O �0�Ôr�[X��,EN��"O8)���PY�)8D�U�P* � e"ON��� t��L����5�"O���ԋ�E���j�'�6,�`"O����R{X�0a�{g����"O04��e�::�� K�O��n_���"O�L�1C�f�a�&��;9m y1%"O�]F��\�X�а$<�Z"O� ��:tGј[c$lq���&c�� ��"O�c�/
�}�9��@�.V�0�"O�4��ݘ|:I�@�N�B1 "O
�p�G� DvU�0OPs�����"Oڍ�E��M���A̛Z'�P�"Oa{fE�*U��l�e��[�Xr�"O"2uc��4�K�.	A(�H�'"O�YK����:�3Ռ*472�A"O��j���!
�1j��c��Axp"O��ϗ�@�|}����_��ĳ�"O��aCV�P��PV�N�Jq���"O�Y�ϐ{��$YA���Rd�ʃ"O���W=0�ѺR��L� rG"O@�`'�Ɂ����bW�-����"O�dCD�7��m�7A��??ޤ�e"OTUSCL��'5�m� �K�lc�"O^����=F��F�-NB���E"O��� 3��t	�ڇL �`�"O�[��=�mr��ME����D"O�9
#���\�"�a���8��e�q"OP�[�L����G-�I�����"O�Wh��3:p@W��n{ yaB"O�ps'eы+	 ���/بK���	�"O.l�� �7|�jq/I8T��"OT��rM�h��1�M�_GT���"O�pHT��.
���Ro]�@G0�k"O�3��N(5Fp���^*/8�dB�"OxT��L&1�L��b/�AXi��"O2��"nY�s��"$@�*?��k"OĠcAB��b�
����:Z���
"O�{gG[���������hy2"O�� ��8%�,; 9��IX"O���엖+f�H�f��i]��"OH�[7��*E0���<%(J�+#"O��I�+�0f��=x�e�*\�0�"Ot���n�.I��١^��!� "Op�(��-:l�u	����Ѣ"O�5(���J$D��R�Y���qF"O��c�Nтr�ڲ`S��"h[F"O�8��(�|�2�U;(b^��"OEƩ.G��Q3.�t6EJ�"O<Q�I�=>/R`J���tZ���"O �ߎ��x|������!��R'~K�\a�R$B��t�LW�!�D�	]lp��_&���t(�!�,}��sF�LJ��Ti�([�!�DŬ8�l�]�&=0�yV臡Z�!�U)�\�R!bF4O����F�dD!��Ɵ~ˆ}H���j>ld됧J�r8!�
=;�~趡��Dݻ���;i8!�$D��m��%wP^�;eD94!�DU9m'��K3��;v9�����a2!�DJ�no�bUaD�t5���DmZ�,!򄊎&l���#ïv'��r�&"&!����bi"�.j����"IP�!�dP BM�%��ɫr��mY2X��!�D'g���p�����*f�D�Z�!�A;z�@U� �%'�e�4(Q�Q�!��,^Al@jʖ~re�A�_���)� ��9�&fjt=[c	��)��H�'$���A�<(h����@'�x��'kT�բP�6��AS�:;�8��'��|�g��m���rGMH�J�!�'�
�����]D�H
���/�2	K��� �4�eDYB�z�.uF�P�"O��`���.�t�6��Hf0�"O�@�3!N JE8����.(*`ta�"Of,�%��W$��!�n�bf��"OB���Y��qaA�*] � "O��H���>���3O"@�X��D"O؈�ك=q�HAc["Q�z=�"O��t��2Ŏ,���e��D�"O`	�%�1'��K�G=OY~��"O�i�d�ل=�4���KL�$�R"O�庲(B�����O�0d$X�"Oj�y5��z�3�G3'^h��"OfYI���z��1�/ÝÚ�"O���JD+v�R�#��P*�:,��"O�U���� �}��튏!�,T2�"O��toF�a�L�a&-ЉQ.ΥQ�"O ���ЇF�X����E$=u���W"O��d&��<�:"tW�`��"O��������U!���v��!J�"O�	���Y*�=Ib�<K5^�"O
�R��Pф����|��l(#�|r�)�Ә9pR ��:K��i�%؋^�B�ɥg�^(!�HZ?̚r���B�75BԬ��#\!��V�)�C�I!�p��u�"/�2��@�fB�I)"$�+`���}��٬xH0B�I
&U����.M�ča�܃{�C��[9R�T$ �'�!�a�tn�C�ɹu�F%y�(�?-Ƅ	�`�U;TB䉯��\j@!ֱ�B���6~ B��m�� ��Ö;s�a���MYB�I�u%�%��k#o��D��;N�PB��07�|�C��d�����X.b2B�ɴ�� Ba� Rit)����:)A2C�I���ภ�
}Î	�*�C)&C�I�{$Rd���J�b�!a��fC�Ɍq��!LM�p^�Y� R�öC�	/��YWě{ܺ��Z��C�ɽ+��Hb'�
�F� e)Y/*��C�I4u���-ѳ���HE-�C�C�	��4�!��ʼe$PYjC�N��*U#��nTrD�L�HC�	Aո�� ɕ.�`��	(��C䉘	�:��b��:_""tɁlݭl�rC��8r��ъ�6u{NLc !ܱX94C�	 l�y�5_3d ��iX�R��C䉆�b��g��T��Ÿs�ոQ��C䉢E�"�+f+Z�Gev�k���C�6B䉸?|.QI⯅�4Ɯ��6�@��C䉘7\�+2 �N��8�1*2��C�	�f8� Q�Q���*T<�(�5D�8#P`���l�����!k.D�|�������;�BJ�j� Q�-D�ă�l�?�`��v�U
��S��)D�����[;2r�r���Z��ljPH(D�,z�\�<�@��^�J����t,D��a��8a�!zB��(+x�)ʱ�+D��x����88dd#D`4�9�P�'D��C��)�=Q��;%'͌�z���'�
���lV+�����	
F ��'�*�*_�6N�
$��'R(�� �'�j��!��zTN�R�<8�$"�'�\�O7D� $��(3:2k�'~2�	�L�K0L����K'/������� �H2G;.Kf�����I��y2"O�yg�ƃ@!]*p��1RIj�"O���Ӣ�t��8�d]�RM�0��"O45	v�=J�i� �>B5d��"O0]��B�K���R@o֮;&�]�"O�x�Iۡ2���S-�A��]X"O�ܩD��s^��cËH8f�:(��"Or�h�U/FL��S�/T�"��Q"O`HQ����O#�M
��Ӵ!���j"O���)O�1��P�5���P��"O
����"����0��=!ָ���"O����	1�@�IF4�RM�"O��e�i��h{�G�4���Q"OD��f�L��9(@���a	b"O��J�-�/�T)�Q�W0\����7"OX�wB�=Th�HAW���;�L��"O$���_	oWZ�QB#��x���q"O`�3�̕�@���d�
j�Be�2"O����e�/p�18�l(xx��)4"O\p��:��H�E�� vY�"OL����2:�X�PܲA���"Oƈ�4��4[y	��
5�Ԭ	g"O6�@�ì2���֏x��� s"O	r�ꚴ<���f[(n�E�D"Op���䕘C9�����1���Rr"OV岳�W������)'����"O:Ј�BB/Bt���C�jp�1""O֭{D�i�>��7CW�O�l� "O��j���;a����]�?\!��"O��j�Jh�go�h�c"OJɛ��T��������273�m��"O���^f��q u�B�t.ZM�"O�shT2r0�f=(Υ��"O� ��V���[�Vv��0�"OzIC[4�i���2�����"OVEsKή!�$���Q�KG�(�"O���8u���Z��J�j�&�!q"O*iS�A3b�Y�'�W�x"""O�0;��WmÜm3e���5�ɑ"O�(Ѷ�.P�pX���E(r���"O4};u摪\���"D��ά�as"Od ��o_p�Ό�0o��k�ԍ
3"OF���eȎ v��;��I!x)hX�"O�����` ����]`d��"O�p��m�LE�A�҄Ўr��%ɷ"Or�A#ۉ�
2W�T	 �|1��"O�8�܎�G8�=�Ս�Q���J�"O�܂�C��i:���*���`"O>�2��v��|��ɘI��q��"O.5�Eϊ�h	v�i�J��D-x�"OB�Sq�z��J%ǵ��0��"O�1�% �=zbM�@�@4d�F��"O��B��Z�B���F� �Hh``"OT}���W��]�UI����5"O,�����K����EŘ�;�LY
7"O��±'^�<�!&Z�(bH�"O&xvLŇj���Cv�]U��X��"OƁ������H�ش���X8�p�"OH��L5�� �K��A$"OXHUgT�;MZ��A���q�(`:U"O�!����4��U��цQ��i2"O��z�Z:4���D
��%��hrT"O��*C�c�l�zsɔ�;�&eb�"O����%6d�$A16ꕨ/��ݒ"O� �	���F���1���A{B�)�"O`d�k�b�&P�b���Nc�ܢF"O.;1��!/谣���,D�8f"O6���)<Զ!����5"�:��v"O�IX���sJT����hpށ9�"O����ݸe��)AbW�Y���"O|���a@7"������*C(�H$"O"��D�	M�D�����L�a"O� p���_������ (8��c"O��S��ʇ^��0@2oǪJŤq�a"O��K�D����p�gP�e�@��4"ON�+�G��j@ ����W*�ZTY�"O�HZPA�/#��)��A�9�$	"O��#��$��P%T�l�R�B"O��qD�����I�d��X�3"O؅�$ ąUK��J�ͦC��Ř�"O(`:�[�!�A���`�)�0"O�d��
2iܠ����#^�=p�"O,��Bi4�l�n� AB�"OjX�dԤ|���x��%��\;�"O^�:�.,Tb�s�1_L��"O.e�d��-#h�ʡ���4Y�#"O��TlĭSJ�| �e�K��d�"O�+ǂ�740��C�r�\�S�"O<���y\aS���hX�"On1�QaɡY*��7��3ȅ�"OPL�$��)�)�|�Z{`"OԄk�m6b>~mk!��"����"OnQh�+�P��#`�7(iPLk�"O�u��(�-��=�R���K�j�7"O\q���'�y�%UDI,}�'"O�C"1�!aU���E��"OF��._8/�]��B�H�dXp�"O*D��,T	����P�n�6�� "O&��a�^)w�\��+���"O U`�
{Lq�*ByF�"O�%Se&�u�1ɂ�T�Dր�"O�=ã��:%׮O�	8�8�F"O6ٙ���"A��11W,3��{�"OT��k��@0�kLPt2�s"O��Ҫ
�_��]��d̕2���pp"O0�����B��=�@:��tZ�"O��!�մ/�AKE@��6� <��"O��p� -DZ�HJC�ӱ�ѹ"O"��(�5
���<�4�hq"O\4�f����QA��S�K�N���"O�p�0�E�<hh����/8���"O
0���W��'ԻK�QW"OB�{�b@�ZM�S�ӌ,�`�3"O��&�@�B��m
fW(P���:�"O�4Z��S�J�F���K��`�"O����>jm���_�i#Tm�&"OZ�'���	���DS��Y�"O�uZ�$��<>$p� ŕ ;�.��C"O����׾B����D��d�:�˵"Od��C
](�N���R��r�"O��"�	�@�ȧ�ƿ!���)c"O��p$�Ƥd{�܉4����:aJ�"O|c���nZ�)��-�2�I�"O,��B ˑ��QC���!N�J���"OP�Cg�o 	�O�7�C"OʱA'N��wmD�Q��\Y�xL�S"O! ����* x�ݠ]��ѐN9D��!,�H�m�Q;ܵ�6D�� ��b2��!XH%���_7�:eB!"O�s���I�*<j�)����P"OBE��I@�����"'��Р1"Ot"��9Q�$��m��v8d���"OF�s��P.�$����Ȏ (�p1"ONM�
-2��0���$a!���p"O��;���!�`�[3�N`���7"O�,
$�,/C��G��'�vE��"O����AF�/��E�,�T�XLQ"OVlX%�<l2\�B��/r��$"O�JՏ.�|�Aa�Շ��i*F"O:�(��H,h�I�V)�>"p�"O�� ��s�BdZ�H;���"ON���M��|��=<��M�#"O��y��1xP�9�6��Y�|�u"OH�5��W*�H�E�U�Y���"Ot��C�(�+��Of*Бa"O
I�D�)����%�2����"O�{ �Þ&���R��0RQ$�?Y�!�d�9:�q����f�aw�S(�!�˩ ���)ŠT1~�$����p!�D�;��eET���(U���Q!��<3��j�Y�z�2�����8l@!�d�Qv����m�V�q���61!�\�>-I2�ƖzR
��.
��!�$ÉK�l�b��FQ�y�`�ͺ�!���78���KZ6K��y�.Z R�!�d�10���9��ߚt0�P@.A�9�!�dەjg
 �tBǴId����N�!��$O� pa�	�<=��BŒ�'|�@(�7Gc�<8��"O�4i HU�i���R`�B�L�^�s�"Od ��,��#���J�&S��)"O�D�Z�9rHsu�{�J�2"O>���@� �8 D� Q���"Ol����A��L2,^V�Р�S"O|Y+�^�!lEzīB!�$��B"O��8�.(���B�K^,j�X��"OH�c�,Ӗ����E��p'I(5"O�0K�j��'��AB��č^� h;�"O�Lig��W���B��.~�J�"O.�bFCǬV̔��N�$J��"O^���"�&Y���O�9<hYd"Ofq!�ǅ=�X}��GT.���""O�TC�O�J�R��c��",~��"O��3 ��: �2���.C�uY"O���� ~%�${�E:z��A�"O�p��K�(s L4�#̳0��H�"O�d�@I�8���1�3U�"���"ON�� CB)!�������X�p�Q "ON��h� x���K6-]��"O4�YtB�27�y+Ń�� ��"Ob�1��J�R$|�#M<%��}�E"O��@oI>n�д���Ԫ¬}��"O�@�t$� H	����7!�@"OZ}8ЎO���@�5��q��"O�m����8�`
�C�`����"O��T�T�!g*@DV�LѠ��"O�lI�)B2;&�L�s���v-H��0"O��kS�&H��}��@�IZȢ"O��ZUFE8�h���M"<��G"O>�����259� ��$�z�x"O�j�C�5� �h�O�E�n̲ "OZXڎT���x��S���	2"O�  ay��ݧ���5�E�\�ZUp�"O<SW�ݸ
��#����@H9r"O�P����]Ք�1Ck�"3�t��"O~d�u�ٗsĮ=C�&`����"O�AkWdO�3-��i������"ON���G�*Q��ň�u��("�"O.�S���0pS� ��^�bt�l�d"O������U�L�b�̉0Q,�c�"O�IIV�M���5
_�_H�K�"O,%���S֌�P^aȰK$ܙ�y��Tu��� ��H�
�S�#�y� �=�@Us+S���\����y�J�-o���h�!�$8��T���yB��x=$z�+^t���)ٕ�y��d�(�Ł�5ePR9�)���y��[�)S(�4FIL�pAQ	���y�ú#y\[c�U�T� ��@M�?�y2oJ�z FmB�6�0%�����yRF�h�b�b���0���;��
�yb��3<�X���'\���a��yR��֞@U�M�%tؑ��y�>C�>�S�L�p&8��m6�y#ҥ} ����з;F�Hc�L#�y�GǌULP �(:נ[')���y� �)h�+#�N�Af��yVN��y�g�Q�V��G@�>�"�j����y�
��=�����͇:�N�D�9�y���>m����`�8�J�&�y�	D7n�|�s,PScT�ї��3�y�j(,� ����-txi8$��y���"zجKR,�l��Qs6I���ybA�?���%��kN���  ���y���KR�3Ңu5P��ɒ&�y�5!l�p�/�?��x�2G�+�y�G4(i�FkhP�b�K��y��؈UD�Rk^�+@�1R C+�y2��9�67fS=~	�(j�yң�v>)���`[�5[1��+�y�c�����^ۦ|�☌�y��@�G!�cO��V�"m�`BD��yBI�
 j��K���'G� P���ܟ�y�2�0��&� :*fݲgÄ&�yr�D(+xI��H"+���:��Ҟ�y��T�k:�3OH���lb����y���.0(PzPeS�b�F��q�8�y�!P"WW�az�	�6f�
D+���y�N�7a�����H�V]IT�Ͼ�yr����h!�:��:�!�>�yRF��,B�m�D��L�ai1���yb�͇r��AP�C�8H������y"D�
%�& �t�B"{�&��DB޳�y�]�(@��z���p%0����yBj�d{>̲�b�
g��-��_��yҫ��d��@�Y�r����A��yR��#=�2Be�ͪ=q���\��y�DF���¼a�,y�a
��yR��"��U;N�XY��b1��y�DS�{��U�g�ڲR�ܙ
v��D��L2X(KÌ5��a���L�8v�ȓo�*�IUdѕֈ4b"�� X3䔄�U�p-
�\�ׂI(7�Q�)��~�⤓'�P�Z�(�;�#� r0�X�ȓ'���g��e����v>�L��+@�A��%:k2�_��T@l�<� ���1�)ņH�j�p�5@"O��J�T�Q� ai%*E?W�A�"O��[W�� m��4٭2VN|�b"O�bc�-~/PH�ūCjتB"O@�jE�R�G+HPp(�9���f"O�)��!��&w�զ׺U+���W"OX�УG�H���C��(fN���"OHY������	�q.8v*<�5"O&��eS\J�y��A���S�"O����N<0&�ŉ�*y�v�"O|xRK2����K�0Q`�z"O�\�&��΁!�O]�R�|�!"O.d����"\s�}�w�@�CA����"O� 1�NMt���p�L�_��$��"O8)��ף/x��0*ٷR��hr"OViJ�J��`���:�I�/�Z���"Oⵁ�m�Iu|�FD/cШ�"Or�3uOQg/茑�e�L⼺@"Oz90v�X�T�ʄ)2�U���1��"O��C��\6I�X���e��L�U"OD]h�	@8+~=*�K�Pڜ��"O���%�֥?��)�`�/-`� "OL��s�ڟJ�Uʛ�|�� �"O. �g��$�H�FĊ�(�PhR3"OJ4�愍m�� �dE�<R��&"OD%z�E1+hδQpc�?rD�d�T"O�b�ѓ��ԀpK

��"O�ثMU-Ƽ��
[�A<�T�%"O^�/'{ ���k�<*:��)�"OX`1H���0A�b��A��H#"O�$�D�I�0��Ô�`]2�"O��A^�s؀��D52Q�X�&"O����G?8U0�(�lѫ=N*e�"O��+�Œ"��t�Q�T(F@�˗"OF�I��,1�8�a��N�gݪ�"O��;�K�O�D��U�� ! ����"O�1��A�2>,0��8I�@YA"OȕcR_G�Ω�ƙ3��u��"O��K�Q�Xn��ö̆�WDH��"O��j섰@ᆊ�@`
|c�"O2I���؏p���aV��5d(�	W"O�5"�X\�0xH�ؗg��:T"O!u98=��3�
@�t{���A"O���l_�),�Y���
VK�a�"OZm���A��A��x= H�"O��%n���)2��Z�0"DDQ�"OJ\����.��1�iF (���4"O`P��F(8���]�xa+&"O�A����10��`~͊\��"O��9�$,� ��F��2m�@��"O^�S��J��`�R���U�"O<I���*f��t� ��4�x�B"O����7=���Vc�a:b)y!"O�,��ɇ�i?��GA�2܉�B"O���!��h�ԁ&B��s4Q��"Or6y�B���F.^��NŪ-!�]��Z�QOP٫�&U�{ !�H/2ق�3��Y�a4��SGFG�!��F�(d��r� ��2Yd�%?�!�P���Fk�(�Q��!�$��@��Q��闄M�n�����9�!�DJ1[��1����7D�j���GF <�!�� !8�|��Fl�FF�&\�!��`��� �N���	�Mu�!��  ����]� x'��v=��H�"O�)��$��zd3v���r��%"O�����N�?b�x�.�>�xE��"O`阃�Մyy���r��1�.xR"O`��G3'5(��L�{����"O�u�Wꞹ?\�h"d*_�Qʆ �"O�xX�N��>V��IG��T�U�a"O~�kp+R��r�M[B>r�4"O*�È�j����e#��n8J	�B"O(�S�/�I�ʶ�##:8��"O�x���'�R��
P�4
f�""O$�ӒF�!X9�@1��L�^�<��"O4�I�+H���y�a����`�d"O��۔�1O � � �"��@�"Oxh�&��_r�SW/öp<�X�"O2� pj$�4<��M��al��"�"O|1Y� ֙x~�$[%�jW|�sG"O�Ps�V�g<�(�i�#aK�
V"O\
%��,_@H�D�W>g�`X �"O^}����=A��p�g+i�pbF"O�H(�/�5�@�2d8c����"O�M+�*�>��i��ͥ:�%H�"O���&�9hz�|bb�4b�&D�w"O���LLn�(�`��u�$�Q�"O�d˂��U¦ *"o�$<�~��"O$@;��f����������G"O\i{%A��5��0M_<WPza�"O���ҢY�p���cY����OL�<q"�6e�j8	7�"!F�P��J�<�OT%m�b7�@'U�l�0/L�<�e*n2.%�b��%����L�I�<1��*D" �q�D	`&�@S�i�J�<�2 ,�K��L�~�{�l^C�<�MUc8%a"hK��Ġ�GOX�<��"�a�So�p�={`�V�<ɂ�^6۲�FÝ�"��`1�Mv�<���23��8���O���EX�<�&��t 1����4�
#��Q�<q��m*�%�S!i��#�D�v�<��BN;n DQ�f�J4<:Ako�<�@"�;O5pY�ȃ�i��x@Q�<A�΄45<��@�.��s@�i��Jx�<��I�~��������	�}�<�3OC�k��}��-��Z"�K�nSs�<�������;7��i��кI�r�<�é�*�PԨu��H��$J�TU�<����*�YR.Ɣ8n�i �N�<i��0LX��S���h�0G!H�<1ǋ�?V՚q�/Ն  N���o�C�<1� �.qr�����?!Z҄Cg��B�<���K�Fu��S�7G��8$MZ�<iVH�<;3���r��5 P���JS�<�7.�%O��Aˑ�O�X}�f�	N�<��#.���S�)^<5g2=y�k�I�<y���� �8H˲f�0!�V	cA�<�E�N&�l��H�-?d.4I��@�<��	��"Ҭ96oΣ/��8'�~�<Yᤆ6.��ys�B�XfXhp&�S�<�6gS�Aº�h$�B�nի���N�<QE	C�?������	9�d�#cGV�<���6?�̨KCOQ�t�MFR�<�֫T�0��E#W�d�5�i�<�d�)ltAz���f��$���n�<�a��#F��R��&J��C�i�<� �ʂ��M �� ��c��E)v"O4akQ\�I�He�����w*O�d:R�� �x� �4u�L��'�`JG��]r��P��=�y!�'�Xݲ�˕M��@���F#~�v��'n$�+[�o����r'L�|䪭��'�y��Ɓ*A�"�̀n|u�
�'o���"=,��Y%����Ҵ��e��4(��^=!<�laD@��l��ȓ̼e����;v���	g�0�ȓv��sr�O5P�j8�6o	k P`��?��=��AT�Xp��A�w�@�ȓ<JpPs��� P*�@�����A<Ω�ȓd��s!�a�âCUڨ���Dמ�1��Dϔ,���D��P�ȓqW�P�?6���TH��.Q��n-�U��V�It�r`G�8]���j�����,�U�@� N!�s"O�H��[�1^��öeݵp�T-H�"O�4�l��&n8��e�,PҊ��"O��9���3'ر����,�'"OR偛a�إk�"W�qu2e`�"OJ�8e�T7�(��� N 	��+0"O
x1���3i��[�o�%2⮸ZR"Opx��/pv ���m�
@�Đ�"O��K�f�k�p{q�\�nL��"Ov��Z�J�K�+t�d]{"O��1�A�s��srk��F��A��"O���. ����:��	*!�Z�1`"O"�sq��!��¤
4Va(�"O��t��<3~F:���
{�jᚵ"Op`0�D0\�x0�Q�V5�m+1"O��� �N? dB��N�L&>�;�"O��o1T��sB7;x�M2"O�d�V��#�)Ò�5+ÎX"OD�"!�!�|��C����ٴ"O~Y S�_3F�ȑB^D��}y3"O�y��X�V���ۀ;�R���"O��H��C�9��R�Yw�P%1�"O"�{���+ ��Ѐ�U�/��"OZmC���!ف)O)�&}�"O�	Kt
E�$th��T�y�hL�4"O�\����G���PT�̱T�htS�"Olչ�;"�f໱C̎b�I�e"O���ʀ�N���C� S5[4B*�"O`-Q�f�\ؐ} %O[�2�"O�d��)CdQ8�*�c 5K�3�"O�u��]$#	z�����N�.8!"O�H�3n��9��ţflI6i ��3�"O�m���8C���B$k�\���"Odp�R�Ɯ*猑h��W%}�U��"O@�#s��/Q�ͱ�O `M��"O��f Pp��k̂-NA�9ca"O@��,�~V�زQ,�����"O6��s�I�,#��"f��Ȼ�"O�M�M�&z{������9T���P"O�D��o2(H9�ʟ�q�zG"O����*�D��O��QE"O"���㌄Tr�M���B�X׀6"O�`���2-�� ��j�&g�"}P1"O ��b�V=8x40� ��lr���%"O�<�P��f�*��O4<�2�C�"O����A�5Y���kU���=�*���"ORԪ��;����.i�*�"O�  ���Z�\y����jB�,���A�"O��J��.DL4:t#P"mvU; "O��� *ºM5رA���!"O�M�t��<���"�\�a"OB��gM�U9��I��{;�DA"c"O*��$	@4P�:sHJ& ��|��"Ol����N�`PH�XE�@N��I0"O�4��\�H5���=3���0"O���n�3'��yu(&�"O�t�I	�B�C�iT=��u"O(��#`�8~�I�w�[�hH` �u"OV���� s�$��p��H(`"O��x�Q���1R:���"O�$R��$]F9뇣��6x��"O�a�˃�
�Je����pE3F"Ob�qd��X�-�V�U���	#"O��k�(�#NV���A�*u�""OR��gW�O��9 *F�c�p[s"Oͺ��_�.H��J����`%��y*O�"%�N���JV�I��`�	�'�̴z�ږ
�v�+��]�w:�H��'�:Lx���+ �Н��b�0D�PK�'��!��:12�uQ1Č�9�h�Q�'��	�kq���p'��,�����'-�x��BN�z�.�[Sc#�\��'m@���H�[m��ɦ!gH`��'��N1
)��R�H/(!p�P	�'F�q84��s����!d7+^d��ȓ<���Bǉ)]��y�Ƿx�J��"D��x�ƅ
���!J�9���,D����&��q�Q�݊)TTr))D�`"v&�>q��ER�"@�,z��2��1D�p��/�M�xE�F�%ZT5�5E/D���"�~o�pc�{��M3�N/D�P�c�ߋ1��㇈�8n�ȡ[�!D�r� ��5�Eg2u�z�f$D�|Ȗ�[Pl��R`ғr���`B?D�t���&5�tUiu��D���'�=D���1�>�sv(�W���XE#;D�A�$&t���s ��8��c�4D���T!�0g�d� 2'ό�P\J�o-D�$��`��
��C�m�~W�3k6D�l�q�Y�2�"xkW�Ӡ+BbHf�4D����CW����\�4�J�ɲ�1D�d�Go@�p#8EY#�;Wj�j��1D�@��6Mr�(H4m	���y�P�"D�t��[�+��U��f+4]pa���<D���TCI�pc ҧ�B�!��<D�pQ�E\#`�;��ёl�؁0)=D�hP�OT�	����R�4��ѐ�D(D�p���O�@D �@i�3y�|�Y��*D�`��J*2����$���\�L���'D���P��(Htը O�.�2�H �1D����%7 Ac�� yYS�*D�d`�:-�c�e�z����`)D�T���ޮ/���[��Z�I��*��4D��SdJ�b Bl�b!רX�x͋�/D�t��"D�xKh=����C��u@8D���u�D"u0'L@�@�t`y'5D�D+��_c�c�AZ.'�@��Ǥ1T���!��4<L��R�I�eX�0"O\�K�
�6*��2�P�M�Xp�"O���۬sh�V�R2}���+D�L��uH��2�
a��QD�<D�� ,��L��[mx�,��:\6�x�"O��V�ׅ��0�ˏ?-9`@Q�"OR��P�M�6��(@�CRf�۴"O�	�%� i��3QOR� �[�"O ��qEĄN���@ծ�.���RV"O�u�
&�ܝ��-���AZV"O����
8J�PK��ߙp�,���"O���ӧ1#�``���Z�~����"OLUA��R��6p��P�g���5"O´�cD��}��<A�l�3Q�j�"O����J8c��pCta�&�Ԛ�"OҩGC>C�z`AYu8�B"O���+1W�Prq�F�c�"O��Ak�'�\�d�$TL�C�"ORB
����S�I_�;0 �V"O����'�o*d���T�B}@���"O&����J@��TÝs�j�i "OܤIg���yYxp��D�,�D��5"OΥ�d�υКd�wI�:�Ή˃"O\@���(tot�P`�?H��B"O�Q��@0Be��Yu��90�L+"O�l�"�øXv8iCG�r�z"OF��DD�^�b�Q�Ȯ#�a�q"OrU�B�4�@���o���� "Ot<�7+I���%��7u��h"O2��0㎙z�Z5AU&Z�v˺�h�"OԀ`u��_�Rg%2h��8��"O�(�d��#�2���T4zeZd"O6�k#�G�{݀Q���L� Lа"OXH�/�GIu"G�W#g,uK2"O���Q�;=H,S��IU)�l@�"O2��$YJ�Y�nĔd���"O`8s���9�a2gߜf_b9J�"O
�sF�^�?���;aE[��&	�"O ��E!u�-[�"T+e�\h�"O�y���1vB �G���t�j�{�"O��� L��a�J�İ?�FU""O.UB�P&|^*Q���%1����t"O�q��5L�UC�Z�gI6�2"OD�Q�D�!)��=ɥ�3w/�0�T"Oe7�QN�p;���?Zp�"Op(iL�6}K3�Ο� �"O0�q�G��\�t�+��E�f�Z1"O�����+fج2 �<�L���"O���2�ŽỲ�g�� n�`l��"OzĢ�n�y}:}挏|r^}P�"O&MC6dX)k���"�E�#D �(:�"O$e+Fl�7���&�n��W��yR��$����#�@�d��f�O�y��=5pxVK�L�6�)�����yBd����<U�ߓZ�b���]��yb տT.x�j���N���$(N��y�o���H�)�D�}�$���'E��y�i��=C�<F^f�E�����y2JŐ{\���B]: &J� �?�ym@�M�.I2EȚR���o�?�y�"�2*a)%�5�@��I���yB�"a����eʗ3�) 4'I��y2�]�x�H��2B��}�PG��y�h׿<�4���L�iQF4�7c߾�y�d�,esp1+�7Q�}[�o�6�y�5��Q`��7D��&���y� Y	b�T�٥��4�`́�+ ��y"C�jW x3ׄL�*�H��<�y
� v�#E`�/R�"�w���6�, D"O lp���e�1��L3� �)"O����
��a
#�`I�"OB!�7$χWJB�X1OHi���"O��`�$��v�<�j��X��P�"O(1�P���,;���`a���
�R�"O�`kG���f�H"�"h��ɩB"O��҄H�j�\���+ܣ�Xd�S"O�i2�.K^�� 	�*E�Tih���"O@U�U��R�����H�</U��"O�}
G���k�zaG�G�a�"O:u�EI�e��dߡ>��p"O�m���$9ݙ��Ř=�x��"O���e'9\���;�E@�b�����"O�5ړ��%,�HP�@�<����"O��4sHݩPƋ�4�1"O���@)L� �Eٲg� P�A�p"Od%�3A�55t	z�L��H�v�B�"O4�6�5��t�Ǎ1:8�)�"O�5�@-��4����FK�ZR(б"Of)�FHT7'�.Ezd��;4|�5"O��#�	)p$s3FR�Y�Z��"O����(Ӹ9��
��I�لb�!�L�>����m��JN���j@*�!��]�3��yS�f�44�H��
��-�!��ޒcg̥�U@�/3"���j5w�!��.h>��3�X�%�Läǁ;T�!�$�d!��`��9$>�P�Ʊj�!�$S��1A��W��L�q�ɢ%�!�dO�o�h��	Y�4ga�&܍B�!���w�,�"pL0��A��<8�!��Q�	:�����"|���s��!�ρL
�H)����F�DJ��[�!���"��3�$�>Xh���)�!��+�,ZQH
;N��VM��!�_�~$��C�-���'*�!�䛢F�x�)��!r���l��HB䉐��lp�ˁ`@18���8?:B�I-2�zUa�ȥHq=���
�zC��/i�`�儙8$m�1I	�9�BC�I-ޒJC(T�[�I+�ğr�B�	3 �8��r��=K��8 bgf�B�	$ZxB�����q�����l̸t C�ɭZ �%(�d�=/u412EE��!�JB�ɤ��1Jef�]�$��%z?LB�I4P��+EƉ�D�UY�_�E�BB䉚 H�S�'̘
�����N\;~�B�IM� �QW
ԉW�zɃ,>4B䉄):n-�f*�'�H�vI��v�RC�I#x�.�G)X�6��aEv3�B�I(1�jԃ���#�Ɯ�-ɩJHC䉣<�4�;䡄)qZtD�$�/?��B�	<7�@��T�ǿK=$�qa�fsJ���+�X� O��/��sW��S�A�ȓUf���G/s_G�	z����i��L:1��)[.�ă��Z+j����ȓg�d`Q �U�K�.ŐeP�=Ѐ�ȓm����T�b�,=)��$�F(�ȓ&���1�A=%n���s�A���*D�$�Ş�]Ϻ�1'D�!Z�+�g4D��%Z��zqY�I3(<0�N1D�Dkd&�6��;�(S�@�:��/D�X�w�R��Ɖ�2%�$b��+D��&KB�D��5�$����0���
=D�� p��ӭT4ra&4;�*\�A�N"O��
'� s�R`��#��u��"O�pZ�C����iW� s�J\Z�"O~����K4G��4J�b��
����"O��(@M݇1��$ca�Qo�mC�"O���B�'�艠�NӬP0�5�#"Or!X����&P�[w��"O^X�c�6+˴�Y��S^^Ih'"O����Λ�XBԁ�"Ϟ49Lp�R"O0��'��`u���$I�	:"O��{v��'j��P	࣍�L/M�s"O6���R�A��тޞF� x�"O
�'
^���Ѵ��՚�`"O��5*ߨT��4�rԓ5���q7"Ov,
���'ܘ�D��,�����"O�ҡEϙ)L8�K֚z�r�6"O`�!o(~���'&�|H3�"O�����B�AJl<Sc�/��q�"O��)q�ߕc���;�섅��pV"O��ApaIvwZ����Pe��,��"O�I6ϖK�2c�ԭj���`E"O\�1�<6�����
�����"OD���D- (�,�"�T�"O�i8�+�Y��u2�A�{����"O6����N8U�^�	E��^!U"O	s��)肴!�,��[�����"O��h�O��wh>Z�EQ*\�)t"O�,�`g$U��A��y��"OΡ9UZ�a�!"D��HLp(*�"OB��q�۬37�4Xd�Y�u�ӱ"O4�!��?N]Ѭ̤7�r���"O���B�6n��Y�,�%W�*�[�"O��6-á��y{gP�|�p:�"O�J�U�v�%���X
	o�Q"O��3�WX��h	��Z\�HQg"Oh5�R���q	 %�gS7o4@Ap"O���"E��@D�H�N�b	�x�"O�u��aB�EޚMӴdT�M
.8��"O����R������2x���T"Ot�cڄzT��GM�(�v�4"O$$�3h�\�&h#b����	�$"O��p&mE t'�D�di�^�Vq��"O�!r��j��4HY.M֜#�"Ov�����ER"Up!B+��3�"O��M�,t@ȱ����a�c?D�x��d�z��oB�a5X��>D�D�P�߆Ry�i��:u��`�<D�8�dA��"�c�3E��i$�:D�� $S�K�\�O� ���ᶥ2D��5�
67X�
&b��	C�*D�x�T�#R&�MRu��-Or�B��)D�@1 a��������Sm�`�$D��#h��T�4���D�1��˰�#D���B-42(@h�� %��@36�#D�L����+���@#�� -J�!4b5D�����V�L����$� bb��G2D�<�e���HTH�	W8Q�B0��3D����,S��T��F�� J�yP�6D�X �j�le�`c�L$�F�p#6D��p��$k6Z�;g/�'I�`��f3D���!�ID�U����t�W
0D�� �.M�qqv�As0�v:D�����N� К��cҕ5�*�
�/7D� �����Ar0ą*&L�(6D�� �i���Y�J�rU�ƍk@���"O�=u��>"e�O�
��`�"O�q��n�����O�Z�<��c"O�8�b��#,�p�+�M�?D�)��"O&X�#�%
nLP@Í��:��r�"O��d
#(�4}z�ʼP��}*�"Ol)�S	 ��[��OKŚC"OV�w������� a����@"OL�����O�d]ا�j��,�T"OBpPa͏�8���*�HvP��"O�* ���L�n �0郍]xIg"Oɢ@y��i  h�;#^a�1"O��c��A]ϖ�J��
	\�EY�"O.h��	h��	��4��<�s"O6�ag*ěuQ���	/2���5"O���6B�J�ˁ�O�h�Jp�W"OJj�F-Ҡ5��ú@0�0�"OD�[���vG�����=s�"O2$�ď7(�>1��c�:Q/��p"O�&�	��α@u�6TsV�x�"O ���@	�4���];4p"$��"O���C�/��\�6NM� QZ��""O�����һ{j4$X\ʨ�"Qn/�y��-��%s��B�^k�0q�� ��y��)I�����-T¸�@�Œ;�y�iO�1.�+'hL� �ڱ����yr鋥r@�٧�ń|!&��&�ˋ�y��Ջ|(T�b�	��D�0��m��yr��BZl-kS�
7��D	���y�M�#W6��Y��Z�8��ٔg�'�y2-W=l�xh2- >-240#	���y! �2�8��t.B�:R��`� <�yb��89�.���4g�dx�'���y���n4��Ѐ�ɹ+�ֈ���	�y�m�'1o�����*�=Qf�W�y��������AB���HƆ��yr`�T�TYh�MS�$�DM<�yRN��%�W�@�R� �5,P��y� @�jA�K6E1�����	��y�K�]�ᐡh]!@�4�	�e��y��B�a�F��a��6�z�3R��(�yBJ�a�.��4�Rk1f���yb�H��䰻U�S0^�Q�a»�y� \�{�����敢N3�f�ܵ��'�t�_q�Y��ҬR�\�k0�!D�`�鋮`Z�B��ԉ;�@#� !D�T��D�`F��+ ��/A��DZ4�1D��h�����nXbt��"�+a�$D���
A�(��ܳ�B����9s�#D��`���J]�)�$>��U9�A?D�xe(�TzθcAΤDh�9t*D��qQ+z1*�p�iW�sy�����$D�4 �
ߚH�TI��d�+�M#"%D���4�+o��jb%�,�f�iT�#D� �`�=`I����_�#0����.D��� D�j���hޠĬ���o-D�0�dU��<AW�F5ug�-�2k0D�����A`�ࡁ*�$\�B1��.D��q%l�k����"_ pD�kf+D�������$۰��W %Q���pb�;D���֧Ʊ*�J,���$6aP����7D�0+Ƥ%\W�)�H[�\�`a'�5D�b�I-8�d-�`!�*!~L9�5D����#(���Q
}x����3D�� L��L�s@Ȁ�!��B�\B4"O��#�I2���E�t	W"ON�0n�����d�&>P�P"O�q�S�^���ـ3��6 ܨb�"O�y��hA�P��	���M\`$��"O�q�2+D�.|���"O:Q�B�)��@��e�i�24��"O:�����P�V��&�%$��y�"O��1(M�rQ��t�#7&Q��"O\bg��f�����5�ذ�"O5���І-θ,��� �l�2�"OL�1�Ö�o�zi�7-����E҆"O:-˒��R�Di�bW�]]�|HE"O �ԁ@<b���;P+��tSpxS�"O�4%�S�V]Xث�)#"���CP"O$�2V��L��m %	�L��J�"O���ư%�]�2��5(�֨ �"OԵ��gl��"��B�|��M�!"O�}���6!n��[�e�3I0���s"OJ�h4�
�3|z	3��o.$h��"OrH��
B ��@�6 ����"O��8f�MxL sÀ�w|�6"O�� Į��
�`ďĳc��1F"O
�rd�G�S&`-ɤ�� J�Q"O���pe�TT,ԿnZ*5 �"O�TʗG�����Y]�4��b"O\Dj�ߣN���˞�z���x�"O���%-�9P#t`�dLb���&"O&q2����P�R��1%vL+�"O�1ʗM�<V,81Q����h��"OxD�B�� %��M�����"O 8#��-v9�2A�R"r�|�t"O�ja���,���ւUH��2"O�y{w�K���+��X��"O��kPJV�a�0Qƪ�	X�j97"O.h´f�!o�S`�ͼ!)�e"O�h�ݵ"�&p���Kn(S"OB@uE�� J��:3�¨r}��"O��+�=z��H� Y�ob�0�"O��I��K�v��A�!!�p��"O����
�@|v!h���d���k�"O��@�G�g�)k�;֖�	"O�����׀��p�4�_
Q��	��"O<���@sg��g#¡O��9F"O.�P�CA�#*^t
�!�g0�+1"Oeٓ7W �@��W����"Oyq&h��?��QP�� D���!w"O�H#� ϴ�(����|?�0��"O>��4���\�b�kS�0���r�"O��Ð�k֘��)o�H�m��y2,���B�0E��L��Ӡ߯�y��V:�P�%�@�}�"i �y"@ �Q�8�b �bo4H�5�@$�y2���z��)!d�
hd}�3�U��yr�?pz�^2,�rC���y�8A��HS��՘]a�\�#T��y�j�nЂha��ƥT�O�tWl�ȓ6|�`aG�I�����hܤ���c��RQ�׮.�9���F�2�t=�ȓ_T���S�$aC�Js�^a�ȓHb�f�
�vO:�P��ҍb�d݆ȓi��P�jj���J�4>h-�ȓUW4�s�#Ȋt�����M}7�8��6
#�ڶ	��t:!��@ ��S�? LQ8��H�#��A
2I!q\�c!"OBlct!�q�|a��.����%�"O��&J�7.X%
2�;>K0X0Q"Oz	Q�GU�p*l�1uf�7�v���"O���&$V�T�8U@P�J7bqP�"O�u��� QJ�Y�GͻjIzD:�"O��s���Nf^��F��t��%"O �FI�:�����ѳN����"O�$Y4HŦ;���ˣ��d��R&"O\K�O�89���耋A�j�LŹ�"O�-ش
\��	(��67L��"O�h��#ʜb����v�0TI�A�"On=Ia�))�|��A}=Z��"O$���I6�L @�q��@g"Oܤ�V�:@n�ԺGn��*����"O������D�CmلI��!g"OT���E�%-���[M� L�Ĵ(�"Ob��� �d��M�<�����"O&�#���4納a%��'R�`r"O�p��$+6Aps!Պv:]�Q"OZP����ܢ��v ����"O���DOQ�t�n;7 ��*��"O���"BLm(�$�2<�\q�"O��֐Q�N�aIڊO�H�"O��bvNE�R��E�ć��-�L���"Od�(��,i0f탂�U����R0"Opt󀭆�yZ��B'�����"O䜲���9)����P�D�b���"O��s.N�`U��ĉ�4yy+�"O��R��yf�L�GN	-<�8��"O[��!̅u�6�W�}�,�g"Ozl�A%y}64+@�S�L��D"O�ctf��}�%�VnI��<u��"O A2�L6=[��o��D߄��"O<d�%"5n
h�*ģ�72��E"O���� ��mر�_�`0^4� "O�h�"� Ah6��e'ӝ["��bc"O�	��k̸jJ(@��D�F0R"ON�x%*�0km,e2�T!E�&P+"O�˴��O�(��B?|�X�P�"O�X�-�!Q� ���<��r"O�<� HS=�t�@gEh/ج�"OP٫�G[U ��T��=��9�"O����N)
д\����7eG����"O���P-T�&��a�\?5b,�w"O>|�t�P�Gmf���GZ:G�3�"O� C�a��%ـ��Ȃ� ���7"O�	x$F�(</B�!��6?��})�"Oj$�£��B*�fpP�c�	5;�!�DS�z��M����ayRL �h�#[�!�'!B�B#.S9q��¡�E�&^!�d�(M��Ek�j-'͐�;�وQ�!�D��K=ĵ0����Xdo�>�!�dF1R̮heBV�a�Z% W�!}!�$ m2q�!��|H؍K�#T@r!�$P�,xT0��,��,LP��fCC�[�!�Y�D�P���&B5����0�!�D�	l��!��R�5��Ȱ�
$�!�D^�k�B�#Y�$R'j*H�!�dH\�ڼJ�	�D�=*	��"(!�N%z�L��"L7�|M˅(ҥ!�B�<{w�ԑK��)��a!�dšK}ZL�E���>��-÷�V�kf!���;]�\�f+U�?�|Z��qP!�� ��%WG��U�گk�&�i�"O2�B�G��i�lꒋ�<��P
�"O0�6jZ�3��仠OA<����"O�i�6ƊbP��ƭ��� Cv"ODm��˙�s:����,�+� �@�"O�@��Ff���s��.q����"O�
�����;T�#|�B�Ap�<A"*֜pb�pCW�H��`Q;0ɛi�<9��	/pP���@�X�u��y2�g�[�<ek�CT.��g_37��hQ�SV�<�U��2�Zp�UxT�QB�H�<1�d�7X�N\�C�(Dh�Hxa	�B�<�7��/Eb���O��
o"�� iI�<��Ɛn���y��\�U��e��#P�<�𠗳D�������jAb$��J�<��D�;8��
��եj]PG�q�<yP�@�,��pⱅ�r�z���END�<��Hؼ'y�`��+ѿ3~�(D��@�<���W�|q��ip���7T1�%{�<�$������I�P�X��t�<�aU�>@�5�Re̾"fV�H'��Z�<!f+	)p\hp��J^duh�S�<�t/6�P�T�YUmMht��e�<)7�K�o��B5f
S�Ԡp0�i�<�nH�(j~�����  �@PR��J�<���W,T��I<��ѓ���I�<9��Z&z �������|#�O�}�<YËI' 2���TN�[��۷��x�<� �ȧ)���")CJ��ѦMr�<v��k�$�Mrd	�$C�f�ȓ&к�X�*ǹnY�<���V$h
0��ȓ_&rmy�JO�~n��Z��TE�ȓX�6�сMF�f]�A*�@���V���YP`��?�`u��Ǘ��p��xM��l:$��U�%�@9��E�R�Z��v=�"��~�<��>,(�2'O**cy�T�f �ȓD��!�3~.P�v�F��dU�ȓlO�r3)G�q2ꡨ�-��z|���6�ۇ�؎mj���6iѝ:=���v�Q[�H�@�Xq� ˳7P5�ȓs$�P���@��dz'
*mh��ȓ/�2	[���#fu��l��<��ȓ}��d	[T(���͌b������Z�q�Z5� ��-�>�T�ȓnfj��b��Oٸ�[�������ȓ0\5)�
���� l�60V4�� h��A̚�@�<0�/A�D��؇�a�8���
}s
���W�%���ȓi�B����+V���m�!Y
���M�P�tE�+S��\B#�Ĳ
К���2l*�oN��RQ��,cZT�����<.To�pu��O�%G�����:����Co����P�U���#�PX��r��r�	�\�,�LX�v����ȓ\LX�i��ڢ\�.�z��
�hl�ȓ�:���q�Be���݅e����4/D���&�� �&o�>D��ȓV#�h�FLz�LU�n��yN蔇ȓA�����V�W�u$Ň�b|R�@�i�#k�b$C���	9�
��*�8����v�fA"#͊K��ȓ��Ȍ>N>��Si׿^����ȓXۨE�Q/'DnK^�&|:d�'D�� !�`�%X��0��s��Д"OJ=���ɖ|�����B���Mz`"O�| �%ͨ�NX[����pyX��3"O�˶	�����ɕ�G.$�B"O���#C�ӄX�U������ "O�MS�`�X%�Y��U�I���a"O���#B�t�h!����Qچ ��"O�XC�$W����Bg�	x�F���"O ҕ��,���6�W�T�����"O��C&�K��$��Q�-�(YJ�"O��x�o^��c�E(%`���"O$�(�S: 9jq��nQ�~W}�4"OB�w�N�SC�p1ůA;2P:� "O�`���k0h�vN�;n.`��"OddrebJ��(� KLR��p"OeX�$�9Ŷ�{d1@�1�"O��2����Nd6u��'̇ƺ�{�"OFDq!�:Rs"U��g��L����"O������"�䙭I��1�g"O
��j�orb�#�dO�K�tT��"OJD�6w*d	B�Ú4.�R%)�"O�7��72�̌�%⍕;x��0"O"��B�ՁzT����4Mc�zu"O�MA��_�T�C�Ըe�p�"O�y7NA�Lj�I�o� �YD"Oɳg���-���4�4��A�s"O��g�P�ol��3bZ�#��� "O�q�l	6l.A��X�es��0"OĘ���P	�ٱ�"��P�G"O8 �M��@ǺY:�I8y���)�"O�Ԡ��R62�A�`��|?,IѢ"O�	�Lݲ|�Jɑ ���]H5r�"O(E(Ƣʈ|�6�:2a�1nF��"O�H
aiү@�!�o0���!�"OdYYE�y	�= �űq��`"O\�3���d��Y�67�"O��)2⊍#�P��$�H1pހ��"Oz=I�(��k?��K"�O�R����"O��Ydo��L,�� ��%L��	:"O�����ĺ8��=)���I�T՚�"O�uj��2| (����!{uF�"O���Ḵ��"�͓1�hAP�"O��02)S
<�X�S��B���"O��aU���H	�P�P��(��(��"O�<Jt�Ji�t\�cBHcz����"O>9r���_"
����,��sd"OLaP�DJof\�z`a�RF�Ɂs"O (�S&ĭHJ�
��6W��J&"ObH0o�7fI2�P�NX=�"�9�"O�uB&�Z>TSx�)��e^���"OR�R`i&���$_D��xS�"OLMc��*kr�ģ�t���P�"O� 0��2S=��+ �I$.6�-q�"O����험XӞ���NB�65n�p�"O�£ W%"2�x!��?P��"O\̨�mC�@���XQ�F�W����"O(�˳$)�P٦�lu���"O�!����(Y�*�.mR@XBw"O%��/J��1�`̎�k3���e"Oa`�&��+P�U80��"O�9��M%!i����G�U)~�	F"O�d�V/,\��2���+��"O�TC�5�~a4 �+BB�`�"O�� b�bS|��D�_)k2��s"O� ���2K(. �5�i�(k(��4"O�)4�D1>Ƞ��ĜǸ��"OH�që܃���*��,I�>x�"OZ��ƥ�8�B����(:�t�+�"O^(J��F0k.�5Y�Mys���@*Onh�$.�@�!h��-0�\��'��p�	3P�l�E�W/S?��)�'1�|x#.;F�ݐ�i�%9����'T\�'�� rG�$�`J!I�l��
�'\���B���(�2�f��jRQa
�'�h�h�f�,�}6hF��:�a	�'�Du
QI����S5p��'}�<ɶe�#L0�IƉ�$5j�AB��u�<��K�X�9 "��������r�'R�M���J$Z�Ib�x��A9�'���q`�ǲ`����	>z�X$p�'"j���A�jEy�K?p?|�h�'��e�F��))�D8� �w�(5��'K@���e��J��0�GD�:�����'�LL�S#צ@
�$#A`�??�h��'0��B�7g|8kq�H�`N\�	�'��kUeϟo4�$� �E_$}��'cf�9�E_�h
�gτL��=��'R4���/=��墡�KT���',x�G�ݞ9�,�-�~b6���'r�Ԫ<0|�ͪ��W8��i��'�(�8�a	 &�zTÓ���>6�B�'�&�X�M�W����e������'����%_[��ٷ�ڋ�4�{�'W���TdR�ǦS���r
�'���Ä�4���_�bO��R	�'���Wr�5��d�8QK�'�4��w��.�]�D��R����'�$a	VA��L�!��8��,Q�'�ĨRc�*���#N�M��I�'��q2"���XR�;H^���'��0e���H�}A��w��t8�'�$pàBM�H�LA��� i�$K�'�(
�oP& �����/W�U�&(��K�a�a
�[�0���gK+K��방��O{┆�IW�>���-�����j)1-4�bՊq*\#�!��[!E�V٢%��p�t��	��B��,���se���uG���]j� �2��dߤɐ3���ykp%�C߳e� I9��*�5B4b���O�b�U d�1�1O�� ��׳�2HѠ�_6�4H�4�'2����۝2�,��5��6!HN���O�{>��aS�C[�`
�[�&��$�ρK��q�mV�Q�D"B�5<:�:w��]�tH��O��Sh��W����6X(X���'`�|���WT�h��=T3�����j.x=P���r��+��*lf�tF�D�F,t<��+�EK$��FK�!��΋��p�C�]�$����B�8������&;ܵjb�X�8"R��cX?�Ey�hF'x�' �*:�D `�ۉ�p>�#���m!�)�a�Qx�y �+�,h�� ��
.̂5yu�݄%�l���'�����͊#f�t��/]� ���K��d_~o.��G
IN�đ0e�8X�y��O�ۅ��� c��Z2B,��X(	�'��z�ј*��1��]���@*�*4h��1^�$��Uή��F�$0�� $ӽhn��h�"N�W�l�xS*Oи�DGV0)2���)P��@i̩Hqfӂ�ޮ{|�
�����t�q�'`P��f �I5�D�s`F�t�	�:j8xa��mJ��f��p1�5(�̧�(��� E��r|rǣQ��t��I��x�"P/K4�Ep�kU�F� b��B�hQ��|(�ej�>{o2�pǡ-V����6"\E1G�� "�|��pk�h-�ȓ�4� �6m:°Cs�XZr�|(�H��z�T�V�͸3h�9Ʌ��0c?�I�1�q�E˗�p�Ӓl�1"��F"OJ�@�ʆ{:�9��P�����&	U�F�\��di3�,[�k�J�ʄ�(O� L�Y��6!\YB�
 TL�R�'��`��(����(J�̰<<��An�9L�|��Θ��rѱc!�4���*�O�(bw��<vU�mC�0���w��W�{���ԥ�8l����ӓhl��7����-�&ѠdK����fL�9��Uo�<@'��~��LRT$ǯ���aP��}���)�CNd��p�	�]d9p ��B�Ƴ6m��.��qz�'�|!!�D���!t�I�儠S�,OX�ұJ�G��0����(5l��b�Į���y��d֑z�r��X�Aô1H�E�&8��z� ��nFIIiO3\M��S��J8Ǹ|�OԱnQ��q�����ȸL˶�a}2���z��mq�iC!e\��j�0Ӹ'C|3�h�+��K$�
L1�r$G0��ʲ'�5�fbY)A������
�!�$�'��	��Nj||�cA�N��`
K[{�͑�G9@��qP�S��y�o�)��  6�h)�f�A�_
|�ȓ}�: P���8cܚ���l
%D���爃�4�B��m��*��@b�
�?�>YС�,B�!�Ą7B>�q�fFAe��a�41"=��KP���Q��E;t�x��C�^B䉢ewd�rӉ@���(_=0��<	c. �du`�z��ө7�F`y"K��i���!_�o��C�ɷ]�ªmcX�Ct�C'b�t����<�f^���JL�IZt���.�s���`n��ϛMu���ȓ^��)Zf����0����)����ȓmQ�rȎ$I�x�N],p>���f�R܃Ņ�,%���M
�*s(��ȓJ�+1�<���t�#Ы'D�dj��L&֥�$(�,}bX�y5(7D�`s�D�A���db�����'7D���C�W<rJ
�a��$p2��V#2D�L��Ȃ[w[&��~
�țg�'D�$�`�Y�f�АT�~0"����#D���S.�"�x5��F�kM|Ib��2D��!��?L���a/�1ٌ�� @5D�P��ˆ#�Ht�t���3��#�B0D�L�����0Nl��ih�4�TO1D��j��C&�\����	�(��6�.D�
���%v �M�.����!D���G)M-��Qg�����c <D�H��k?��|A�G�V�Ľ�S!D�P���ԅt ��z��ďmL�y{@?D�di�Æ
#��e��A;�36s�̈́ȓR�bٱ�h���v�\RA<<��I��Y��kϣ_$
���%�s�Q�ȓ|��ZE-
1!>�K� 9Q�i��E�������&��Kц\�tҐ�ȓ	�p!���J+ve��S�ۏ%h@��q���H��Lh (�"*�!�`̇�a��i�c�Ψ4��!	Np�����:(�"��٤���gW��d�ȓ$� �;3��+Z��DHۍ8k����LC��gc߽&���f	��/�̄ȓQ���5M�������<KTe��@+�b�׹M�X����Bl��'��1��	X*4N$(tŞ�}H���LrJ�HC�p�HY�HK�%by�ȓ��3!��+?ӆ@��A��+>v=��h�Ą{2�C����e�M�:R��ȓm.�*��D��ȕ"��JX���S��e��J��
�z�C���!���������?h2His��%N����!02z��-_񎜩W%��4�ȓFWX|8�ͼC�yb ýpT��ȓt�x�p,C
|����ա��n@�؆ȓ�4az�΄�#�&x�f[�>e�u��hq�<H��!pՠ��Q�K]\���S�? >L��/���FA�$�P��"O��2.�\\\(r�@�76��咢"Of1��&��8p�/Ş>�(Q�r"O(-jc͔��D�����+5���Y�"O�@J2� 3 ��A�R9��9�1"O]c�H�/n֕���ɒ|�0ܰ�"O��
a송<���qTʒ=)�T�"O�iѩ�"1^ꑻ���.j�ٺG"O<��J��o�R+s���ZZ6�Г"O�����v�$%��b����2"O�=�c�rБ:U��<�$Q��[�<ɖ���H(���r����@N�<���R�j��(E� o��EH�I�<���O�f��Q� \.e!�/�@���5��"����#V��z#�'���#ǥ�R��C�	�g���kTi�?K��́��b/`�DB�1��4#�S���؈�@�	^�QPo�{�B䉡o�t��L�F�\�5!^%C�	�f�M�/��01�'�(:0��>YdG�'�4p��\�^��;qAzH<��cF�l?�%��O:��o�=?�`�����>���@�+�p=af��`��aMA�-* }b6�yX�Ġ�Cڃs]Z\¤�Zq�
�0c�Â�b&;#��Y��'��y���*g�\҇��=�1�$�ø��I,rS2I�u;�lPe��J�>=xV�ҍo�tI¦C2����"D�l����*���L�I��a�4O��Y�쭁�l�x,΄��*_�M�$�>�O�PF�ǰ_�",s��:X8>%)sO�HmG�c���Z���`��ٵ���rz8{6�-`*��zqX\	��d�@�2��R�Xp��7-ӱ.ax��  ��2c�o��QY�B!xT���`�%�Hm�)� )\��Ox��eIO	�<h;���GH@�ї��|�6��z���*C�,z�<��`!�G��Q5�LdoO����'��]����%��|�W 7zk����\$!��3�I|fP��_�^B�Q*"�r�'��WL����x�Ա�aX�d�X��TD�h��_�?��H�"�Q�F�T2ew��� ��"�� qb޵��<�FA����TS����D@Z2�i�@�D�j�*�x��TXA��J:q���eȎ`O��@�^�b: ���(��E�*R:���D`M�I���')$9��i�n����ŗ=kXIZ��i�"G6����t�~	[ĎJ�$x!�Dݵ+"����J�ABhH��_�5k�u�b�+(���4K<��`3��|r��>N��9C��<"���b� �PxR#ߧ<*؄`��U��٠���`�$��c`�I �9����h�鉶S#�A��J�QJsrψ}2���U�&�� �^$�t�FJ�8@x���cgZ�;������_��t��ȓx���N\,htp�DM�iN��&���0�#זp��#�3�ލG���E�D��Bj_�y�����I��yb��d����kP�~��Ŋ"E�D6=`�J^��	4+t)��O�7E�^L"�IG#J=�� a"O촛w(?�␊��,{nFU���x�V���K��y8a|"b��@���b��Z�[Re'��=y�<%T��F�
��0́0�X����u����ȓ+��@���?�Bq��E������ȓ'��(���!	cdD?!F.H����#H�`.�1�i�^x��ȓr�"q�G �@ u�n7���t���r���eCg�Q�`�ȓf��t3c#��W:��OH�FC�Ɇ"��@U-�A<�=�e@	G�C�	�o�"dw��}���*��]~s\C�ɴk!B�A2�]8���C�߾n)�B��+�Mb�/�`B�5_q�B�!o�	�KC��ZqB$W%�B�2c�X��CjK��T�X�C��XC�I#
[�06�yz4릧�9e�C��$� �B�V�(�Xa^~��B�)� f��Um�
�|��a�<\F� "O�I����Cf����
pTQ�U"O�ɒ�Մ4
 �6k	1/�1P"O�yxp�K:�\����T(@�"OL�R89̊@��*p��Dcu"Ozu ��P�ݺ��G&R����A"O��5A�l�����χ!�dS�"O�lpt�ȴR�8����<{�uAD"O����A�9����0�Oh���t"Oz�z��$�fE���${d�(�e"O�=�tbP�9D20�a�9Qrh�&"OJ�����_Z<T�kM�C\�1g"OV4�a��,x\NIӣ�YgL�\)"O��$H�,CE��P�j�v~�@�"O�i��1nl�(�éB�Yɂ�iT"O��j�� "Fȸ�*��&oH�!"O�P�CA�*��5q *ۻJ[�{�"O9	�`�S���0h�REI��"O�0�D*D�O��@')��Q���;U"O
{Qo��F��w�A06�hw"OH�nĿ6vL�`&�ad�:�)9D� ���кD��[Q�ɰx��0��6D�@�s�A���%�P-_��`��b#D�����)<˖�j� '�DSæ#D�8���P�]����UD��Ͷ0S��<D�Dx� Ŕ�9�1�L�'��,��C8D�̺�X�/0H�w
�'td�a9D��RS��ht=�w�ԟL�,T���4D�����Ք9�VX��:tTB�K'�3D����dƫ40\i�I�<�05�3D�0#��;ܸ=I��D�a���` .D�h��Y*����F�b.��2ea2D�$�D.T�f�dC���T���f.D���ceW�P�ve���0���q�!D����([�?�DɛCiǤbrA��C(D��'IL���)���Bz�03D���R���z
m�O�<|��Yr�1D�ā�N�'��p��̄b��!�u.*D�#��Tr̆�3�*C�PKԝQ�/D�Sq��7�V��n��	 ��y��(D�8y�)��L�NaJH�y�i�Ū*4�`�T�G�b��8��e˙R�PXˣb֌N�x|8V,/�O�s#:^"�(�U�@s�����'�B�qd+ 5��	��8ڕ�pd��r��&(���Kw�!:�G�?'TΩZ�F��!����O��s���xE��e�O� l6�W,`�$�e���
�C�'�
M8�ʋ����6��p~ 	pDHP�q���hܸ��s�@b�g̓P� u�T���]d�"��Q�����IQ�i�Q�H���� -V%�.$�TdǕ��b�+�`��d������5m[�0R<A���A�]-џ\�G'׶h�d��嚯�t���`	G���Q��`��S�B��<�}�Sc�O��Ð�~����<7�`j�Ċ3K<ɲ��\=	�?9S��ߚx�h\�N¸\!�9��y�<��h ��-ڮ��p-ݞL�4\�"H�)���m����ɑ��v��	�&&���n�4ڍ0f ��,�����X��`�gf�M7�#����s�M�'s��`�c
�u�Jh��~8��qT� #�8�r��:�Z��4�?U����H�-H�)��
s��#e�?9���@J5�&G>.y2 �)D��if� \i��d����+V�D�d��(�Ƌ~Hd�p��=g�B�IF�ɼ�b���F���z��K0i�R#ѥ�F�<	��@+Ij�v�Ûh�$u�M�&����mL*��f)�^����Ld�<��lܭp+P�T�ҚU����`YV���y1��}�Q�̝.'��i`�*��1U#��f�B�A ���M1�O��d�&6�tM	椝���5(��d�=n�@1��S���8���Yp�p���?� b�+�`�h�Bݸ���Wt<iل"O��rU��8j�.��aєW�nC��+S\̹�Vyq�OG2qk��b��$lۼ�5�O.`!b�R���+
^��s�g�C�<��KY�o������Q�>86�R`�^�:����<� �s�������+!l���<	���@���裂G��\ڇ�}�����"�,4���C�ϝ%I���F��_�0�pp@��v@�n�k� �����p>��@�y� �б��8/b
� ��C�0h���B��u��Ԡ�`�IIà�)l"�	�$z@�����B��m2eB�%�!��cԸ��@G���9A�L�U��h�mڣInx2��X�a��;�`،��O�^!�;4 �)��f@x�|Qy��T�5Z\��ȓ
Kpթ��=�~�S�#��0!F��dWk�: ��IV>c6�C�B��
Ix͑F�#�5�.���@]�+���X3��d�~؇�	0i5���I�:��t�E� ��LQ
\��j�)N�}it�[����I6�1Y���o�b�f�;9���4k�(]�K�(���� v�XH3�P25���G���!Gq����Ō&��C�	����(cl��5ڢ���HM wp��{
�1���bí��+��jg8�'9��Z�H�Y�m�<{X�,"�0}�!�U�U]B��p��F�ݳ����T�P�E�1�{d�<	�,E�`�ϨO�Ԉ6'���rJ�C޿lɰ�s�'��ik�E��iIlH�c�R>o�r�S�9��ɰ�y�a�S�lmqal�+e���"�@C��(O6Pk�!��R�niE��E�?l%��u%N�^-V�Xֈ��y��L�6�<$s�Ǫy���FF�yRm�d�~Y��ဟ,���ȁJX6�y�/�4h�6� 1# XKLP��y�g��l�.8�C�S�k
r�P�5�yB�K� 	YB��v�Fi���M�yr��O�hmi�%�k�v�W�<�y�.;�b�jt%��h�D$2'�\�y��D'�Q�#ʈo��4�ŉ	�y�+C(h-T�sB�)Z����5l�y2�0F
�Y'L�e��{U'�9�y��SN@��#T�T�)�N���yBOܸYպS�:Q���&ף�y­6��H:��<<*��;�[��y�h�=7���F�]�(pT(�`�A�yBY-��b��#���Z0b�(�y.�]�D�j���$�i���y��?)�F��`� 	�`l��+�y"�Ĉ�6����K�!�1.��y2�@�6��9��I�}��l�D���y�e4NR0��π?sB���/ώ�yR���@�ۢ⋕K�ʆ�^'�y���J����
��˕B�y��/���K7.�0�8��
_��yr�Ku�&�1E�ֶw�)�"��yB��-<���EIЎ@����U.�y�@	z�Ҝ˶EA7�$I�g��>�y⍎.5�a+t!$�y��\��y��śr�xK!l[��`�Y��y��׼;�f9U�7'Qz8�FA��y�C��[ L|!�$w@����V��y��T.i��qkD��
�e�H͝�yRDC9N�@ �l�xN���bܺ�y��^S�Ԃ�����|������y��E1�͙�l
5�J}��B��y��G	>���._�0�����݆�y�Z�F_�1���T.]�mqW�yB�ܞX*�$�`bJБV�ޣ�yR��m���4����i4�yBg
7)�MA�I	�6x�vU��y�܅rf �Ӳc���p�$���y��F�xBT�Á���j�xi�4a�3�yr�@�By"R�7uJ���,���y
� f�"�ĉ\��X���d��P"O`��׮P!)D2B�B����x�V"O )����g��ɒᄜTΆE @"O�JD-�3���GB�*+��$�"O���@�H,pҖ"֯�6��"O.�q�3C�b�2AaيZtr)��"O�T�rg��/r(=$FD:a}��Ɇ"O�H�1gF�V+:-S�&�`�j1�'"O��I6���;�0�6�Ͽ�t�zE"Oj��u�
2N������ʒD����yB�]3Q�J-�W�?��\�B��-�y��OtH�bZ4�J�e���y�0��4h�B<��ȳ͇��y��Y�s� ���!�|J�9Q��߉�y���o���q'OW�sw0��e�7�y�E�:+�jT���_�[��8�"�1�yIH#����bSx|��F՜�y�W� ���U4s��C��y�KX�KT�ö�"x������y"Cϔ>����5�ƀp�����Ո�y��ڷ1�h�s���!h��xc���y2��Rz^��4j�:�)
1N܋�y�/�f�2mZ����o����e��3�yR��3���#m<f�0B�폻�yr� �'պ-8�n��S	�)�P���yr�>�tek�ܖT|"�Y- �y��h�4�ycm�*�fԙ1���y���:��M��N��fZJ؎���S�t�B�ش@R�f�ˋ@:4��ȓsJ�����F�b��/��s�4 �ȓ&�=S�g�^Ѐ4�4L��ȓ	e@q���@�x0�0k�D��ȓ�l5S���2��Y�P�N�{����ȓ?�Z��4Ɖ ^*^=8g�/i}p���}p(r�C�9��`���Ϡ�"=�ȓPR���c�0da�X#��%6����^�P 
�M��r@f�:� �q2�y�ȓV��M��O����CG�N��`��դ	��hG
|B�LR%��T��z��#�G�,��@�ώ?~���#�z�ZD,@%��(���8'O�1��	�0�'cU	���!��1jP�ȓ0�ֽJ��W7��dY��\純�ȓH�l���}�8��U&P������`�Zv�X&��d��@P�rUD��ȓ0%�I؛�"T
��p��L�ȓUp��o�2e�n�)�)S��fهȓ�ɫ�B�b2]1�"��w����ȓk�}YWC,zD&�h�lԗ8���ȓ��ѥA����] ֮Fy��ȓ*� ��GI���,�c�F�q�*��ȓ�F��n�jO� Zg��,V��9��E��'F���n��NV�݅�5������¹XA��B
�a�ش��nb�y��Y�;	����A
{N���k���Q�Փ
s���O� I�ńȓ|�D�����K�f�;��a��I����-��]�B�˦ʔ@ L��ȓGff��ȍ#�����(k.$��_��(&�_{F�䇓+��P��}y2��D1?$ {��n.D�ȓ]C` �
�l%�a��+U+�M�ȓb�
�3%ʘ�)�I��X�4��n���CD5%X�Y0q��u�&h��S�? �-Bs�׭]�z�HdF�����Q"O(��#� y�Ɲ��îk��	��"O`�1#�5�|�*����i�:(�"O0M�3
�,51� e�%IH��b"ODR��א~�V鲒
�2�ܫd"O�|¥�E�)`xI
BOP��"O��x3Q�ͤ�ci��L'���"O~T�d�jQp�hJ��c"OL�B���c<��*q��!X�p �"O���@H�nLPB�Q�u6��"O�*�[ m�n�0��:#)���"ON �ȣ3������t����"O��BUjE�k㐔+������"O䁙�E�u��]PB�2>��m��"On@cto] ip�ѡ�M�7H�0-�f"O�ʠ�|<\k���-�����"O�P(��1~��O�i����"O^u�,��i;�Ͳ��[�W�� r"O&y���6{�,��8k�ļ��"O(��bE9�`9��'o8`�"O�YJ��W6�`2��ӡ|���V"O�e�D�ΨWN���!FZ�l��əs��7+��a*ȑW1�tsaMѳ>|0�ɰN�h�&o�:1��ę�n9T&�Dʆi��,���: ��H��
�<Ld@�V��?y.=���t��D�O^,���b?�+d�6M@�Xw�D>q�6A�$��9B�rih�O>i��i^s���S	����U4TX�P���^��q�H�����I�,�^�H<�}2QN2L��9JܔO[0�I$��ly�P�qR<iɀ1}r�!_�� �c]�b�\xR�
�7A�6M�:�x��D��S�0
� b�o3la!���;*����d�ںGx��ƱH6.H�b��1+vj�ozxT� ��۞�2O�3��|�'l�0��u��l٤�]61�@��'ݞ����}��O�>�@j�+
�h�c@�CR������ɸ�:ҧ�'8��O:8x�eʜ�4��)�VΛ'��H��i�N���ƕ�%���	;H>uϧ_x��aQ�_͎�Q�E<vԌ�q�E�.���̈��M�׮�\2���S aH�RザF4�B��=<�F F����M�ƨ��U������Ḩ��ߟ��ׂ\�N9�0�'�2�"�w@�কc�	Ǟ&Q� �'a��I[�TBb0�tc�8V�����LL���B5F#I6���g���d�?Q��C&�p�H2��&��z%�T��cHB�.$�|�i>�����Nx���Y��!���/`~��>���KX>5�v'P���Q�OM2g��M�@�6��3B�$`DxJ|��j��e;`�z��ٖ@�����g�	3-�"<�~�r��1\*�A,6GU�бz�	�:����<|W���Z2t��Ya��?�(6�ʴbu�"���i��a�b�GEx�`�猶:.Q�l�ᓸM��u�o�yV� �Ŭ��~C�I�X�"a���*�z�#G��HC�	9#.<XD�Y k2v��!��V�C�	G��@¬F�izF����A�g�C�	3�2��$��kfx}�b�+HB�ɠ`��	��׮�m'�	��hB�ɐ.1F�t*
�{)H0��G�u�XB�-Yfya�T,��u��!�d�;�>͉���q{2YA���WG!��W�b��<y�B	$Ӕe)ԯ�#0!�$G�M�ѳ��H�%��� ���4!�dT&I]:���P9�hI>Sq!����8�ṠӃp��]�(�/�Py"�O��&�sQ��3L�j�`����y m�p�"l�=qP��ҤE��y2���v۴�z���>�Ur��� �Py�J�+$Ɂ��O�cŦ��'J�M�<�g��[LV`x�"ْC)���J�`�<� �
�K�����J�O; �Ƞ@�Z�<�R��,
4�B��IZPr�UDV�<� U�v�.�r0[��_�D�)�%"O��Aƀ=s�m���ϒ3}�1��"O�t`��\:b�#�LZ+p��4"O�U��OX!4�z5@ኔ-L�)*E"O�,�u�5A��*�#�MI�"OB������A��i�>-��\
 "Od�ss,'!��h ��[�����"O�ta�ҙ��5�B)M�K��B"O�q	���/:'$�B�M"�pA�"Of�2pbS�4�6Sfm�/�t���"O:(�eO>u�����ڟoȴ� "O����@�*�0P�R�Z\�i�"O<��1�K;�N4y����HQ�LHb"O��Q�S+2��T�X'c�> 8�"Ohq�e��.\���+�s	:U�"O�p��L��R- �3t�A�<�4�K1"O�́�-�]n̸;���0Ǌ�H�"O��0Q�Wʶ|a�dW=c�v�9�"Oh����$!#�ʄ-n�z��q"Op�R�n�.
&��ɡW4:����`"O����btlظ���� ��	s�"O�� {t����ۛ2��i �"O�x��ҥ\
"�D�7<$	 "O2(W"V�,DQ���Kz��"O@�cvHM��	#��ħ\�N�Zf"O���t�;H�F��G�#j��$"O�U	L�z��@L���KP"Or�C�o	�*�`���6A�}hf"O|�{��:K9�t�G��*l!bPe"On�`�E�y$�|₌4[��Dڡ"OްB�.�L8��Al˪2R�U�"O�P�E��5��x�"VI����"Op�*$e�v�0��u�[�S=����"O���i��M�-���p,�q#�"O�A�&/]&J�p��3Hʕ|!y�"Ot؂ԂÅl���sA_��� r�"OHP��	�(Mh$AJ���P9p�I$"O,���'��T��҇J^3h8��;f"O�5�@�CV���;D*���"O�%�`b�67��@�bI��l�u�"O���V'�j"�x:���	�P��"Oh��F�#D?���f�-|@ɢ�"O4�bg�4DR��0�G
Q^���4"Od̑���v�)��ɘB�N��7"O)���`�0X�e䑤t���Xc"O�@	�艖LR453�(^�`��M#v"O�a���L]�j9"�,f��$k"O�X	!L̐Am]3r�U@�"OND뀥�j(�� +�9��z�"O@�ȓ�E@�(�s
N8nMD�0�"O��P��+J�,�/�;��؋"O�����/1^��`�L_����"O� �%���R��$����"O��3��\ ��,C�#�Z�:A"O�AS����{7�4������@&"O�l{T�3�`U�k� |`(���"O��4 I�w7���ˈb2�j""O�Hr����%pJ��q	�G�J1�P"O��k�$�vĘBh�Q7z��"O���VJ�8Ey�<
��F�*�\�"O��.��y����r�_�S�xJ�"OrHy"c��	x(dJ�����Е"OT0�tK� k�r &Y���[C"O �Z���rm��EK�|Y�"O� ��qr	̩��A�Ŭ�:d��q��"O Xq�f�t�YH�DC�fĠ@"O���#H�pG��v��7�:�Y�"O��X�c.�9��b��h�h�҂"O ,�Ҥ�+/̖-��]�S&L|{�"O�l �aЅt�D(f�a��3"OHY���E�LE<pA邪<���1"O���5b=&�nЁ%��^���G"O�!�7��/WoByA��	���"OR��"��}��i��J�+����`"O��x5��	I����#H�O�L��B"OX�;5�+'S@���dE�p�.���"O�u��Ńy5޼�!S03�d�"O`M �@G�=��qr�^�"O�A%���$q�O�{yʍ�s"O�5�!h8���҅�˩"�\���"O�@s��$�J��Ra�� �w"O@ف�fҝi��J����� q�"O��iքf����5�Ϸ.N�}��<D����� �P�q&Hѧ{�VI�Չ D�HaB��,\���"��]�1-#D���իJ5Ztb�8u�:��đD�"D�[��KF �g]6D���TL6D��{��U�_�@-�e�NUx)���!D�� �� $vI���Q�03~��A&!D��b����q,ˈd
0���3D�|���:�xE3Q�	���5�+D��KPN����� ���r��YX�)D�Ȣ�N�	�D@@fŌ>�d\�!�(D���a��|4��ђ�r͜���,D��;��V36l"�RvNJx�t����-D�+'a��lj��zc
J�Q�\8�ׄ)D��X�#]�_ANi�gƺ�H(2��(D��X�J�[�4XHႍO^�/X�C�I�f�!b�#�NٹQ@D;}gjC䉙e������9���c4)U�6DC�	�A.�$���(|����g�s(C�	G�"�@�] &F��2cݰZڶB䉟�x�2f�$ Xt�S��d��B�ɍ:��xFd��{�"l���b�xB�ɜa��qc ӣvT��`�J+4B�/[~�}� *V�q Rx�WL��l"B�	-K��2�&^�	Cl��W+�B�	OjL�3�	#��զ�F4�B�'xBE����,����6��;��B�I~F�1�B�J`&<���G�АB�0Z�)@%��,���C�F"D�VB�	�?�2��Âe~�EaE�?V2B�Ɂo�q2�N� ��C�KúgZPB�5J��ze.�������*A�dC��u-�͙�e�.OU��P��=ZC䉹okdh�ɬJ��dK�#	�p��B�)@L��G�S�V��: b�Y��B䉠[���� .���j@�~�JC��/����(�;`h�"�e
;!K�C��/`.{��:�8�g��E��C�	 w�T��ך^P줠�ƅ�>Q�B�	sڴ9gϙe��th���0I+NC�	�Nd�i�LǮl����W49LC�	�"V���nS�J�����9BDC䉾w����@)����y�DL�C�I�U!L�G��h�b]����l(�B��1u���X���69�"DfH�.3C�I�$�d����/O6���F�~H�C�)� 6`h��O!1��ňE=#"OI��o޾80h��T�϶I����"Ov�q�O��.� dA2̆ N�"O"��W!��#=����J^����"O)сȕl�H��
�,���"O�@����-��hعYvf)�q"O:y��(_�k��9yHėgBܢ5"O�]�� �,�XY �ُ-����"OڐC�@� Ek��a��<{U"O챉F_�-�����X�Z��"O0A&�W�Q�$4��Q�:�zj"O� Ζ-2�R��G�\���"OR���%��W��}I�-M�;ߘ�0t"O�S�A7��
w�^� ���'"O��Y�~2�t�O)��q"Oh�0ëO/�D�A���L�\h�"O ya(LV���)ܶ/�J�r�"O�E��oӜ�dܨ�-8�*�!"O�Ui�-��C*δ7R�a�D"O�����"��!��I�8G�ɱW"O �(�$�(Y-n�pT�P�
��e��"O\��u��!�2� �HO"C��=ؠ"O��)qf%^������](Yx�R"O�<���ÑM������gT��"Od�ٗlӂ(�R�QL��h=t|��"O�ܙ����@��d�I%'1��@"Oh���,�aӢ�>}��� "O�̓%�F�)ZD�c�M�D��0!�"O���R��"L�u��%қFY8"OD<��B��`�>�p�KK�=�"Ozl�Č�{8`���*6�� "O��pqꉮo�p3�kV�>��͊G"O~ 2i
� ��� %��,����'"O�M��5B|���3i��H���ȥ"O�9�L��Y��M��h.'��ڑ"O���ֹe�&u��AA9+7�a��"O��I��!R:�ȁIj�4��"O*1����]A�@��a�����"O�4�s��ku��B'U��\+p"OƁ��~f0M��H:B�ܰ�P"O�$9���lPL�c��ϓ+��A�"O�e{��?����#����"O�K�j���Ǧ�;���rf"OP0pt�j���4�҉L�8-A'"O&Hs�CO�O�|�	�h_x�p�@1"O䨢�.�P�X��pmM�a� p�"O�i:AoE�g��c�k۵Vt@@�"O�9B��҅� ��Dʄ ��"O��a��P0|�R�	 �?��Ƞ�"O��{�c^�PD�)"�IL�_�{�"O�q�T�Y`´�H��,Ԁ�"O�S  
  ��   +  �  e  s   �+  �6  �A  �J  tU  �`  rh  �n  u  f{  ��  �  -�  q�  ��  ��  8�  z�  ��  �  E�  ��  �  ��  A�  ��  ��  ��  ��  �  I 9 } � �  Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�� |d��"O
`�(�;���8���-0��1%"Oj4��ND^[��"3/9�0|H�"OB���H��*�ʞRy=a"O�味V�!X��!&F�:J�$���"O,��a
���C�Ą�M�"O,$3%o�-���p���+Ն�:1"O��ݢ1����`���y14]2��i�<�6��{_���c�H�`�fX�$Kn�<��A̼VI�xR[�)�Ć�pඤ�ȓA5��('nߡ4�� �)˩%� ���,��r�؊b#`T�eT09���ȓ!�b��g��}�8�F��-? �ȓ
K|m�ș�VṔ���2�%�ȓ"R�X�j�4JN�1�˘X�i����̹	_�jZ��1!g��zܶ��ȓgil,*�J�
j�Ne��i�J%b���f	�(U��:���G��$Y^م�~r�� S�%T"���k\�jx�ȓ|4�1�îJb��@ӵ�ݩn�V��/[`�"�v4�R�!ʎ<��M�ȓ`:��z�ؚh�J�Z��$HY:	��H��p�m�C1��!��B:��0��EnjZA V;9����J[
2���	��4'J�EA�IVW&��~�(aZ��ӹ�>� o�Y�|�ȓ�f�A�
Ο7�H��M�$�����mޠP����/���ANXo*�ȓTv�����{ ��-7�*h��I��sB�8�8���3����ȓNe*M�悡;������X�o��!�ȓ'lj�#F�m�+R&;�|��2)n�C��0S4���T:
b��'mў"}��h�/�P����RE3���I�<ђjŹqWq+�)K7����c���hO?物�6�r��N�U_�p5��0C��;� س��ܝ8ƨ�9�/ġ@(&�'2a}"Ɉ�B*8eG��6ʄ��@����Ox�@�'L^b>��.؇�vm��%@��!)Oz�$�X�&����JL�k�<!�||�	��y�8�)�!���J�gQ�4�>|9q,���hH>)���I��j���ɀ!�~��7@�yb�E��f	钥�X
�$��7��>YH�p��D]�OqT"�S1C�̽P%$D�y��� �М�6�?3��+҆#�I�=DxJ?]��(� X�R���!G;&�niӔ�%D�ȋ��J"x��ӱ�E9,Z5@ �`���'f�S��M�E�q�f�+s�R� ��Q��y�<q3���;�\*C�x�����Ox�<p��p�0�@�؃x1X52�LKt�<5�֪o��pwK�m~����Es�<!�H�+/T��E�J�!��A�EIk�<#A_�4���P�н%M&T�,R�E�(g�q(�!��}��0� ��LG{��)ݠة7��3K�H8�0�N^�!��J9|&<P���M�$� ��ԠN����>��ˍ6��-YZ0>T5�Ѥ�X����'���s�އyX��RԈ�U���)�':L�b#�9fk\��&$L�^(F����ͨ��i ����	����?�6�X"Oji�r�ѷ��I����z� X��"O��djP�%��U1Fl��B"O� �y�R	E���Q{ �(}�ɋ�"O@��2j* �d3��
�J��'mV��9:n�lz����ܭj�IǮr����<1��#E���*��cD��P�Ew�<	�G�4nz��ƓX�R!�j�'	ģJ��pҲ�[�b�0��}���O}��)ҧMع�UF��"-�5�Dĉ!m����� �W��/	mT�GI�v�
�ȓt�@�q�Z�N���rlQ�|�f��O���D±WΈ�5o�!X�0�6��3!�Dƻ?Aƈ)]is@6|�HP@�"O��ˡaD�\�=#�䞣6��9�"O��9��#Z��0��"+X���"O���&�����8
���tYD"Ojy����j�>��p. �@"O�	���/A����"Iޘp��	�8O�b�\ԧ���� �Bd�"�!=��1Uaκ!��
+)]�sт��)��q��`�3 h��'���4�~
 .��h]J�)�!^�T��h��,�0�d��u[���q�T&7u�YsS+Za�� #��)�-N���S�Hݍ,Z�4�*�>��O8�=%>�� t��50V����-8',D�Dɥ��Mq�����pb���\��hO?��0L�t����xr  ��.X���Ux��"� 5��paR��:���Z�yrE�7�8ɱ �_]3�0C����>)�O�xI�暽>�[� G�Ag�C�"OT5;��4s���c�a�X_v���"O�����Y��*ᨗb��W)���"O4lJaʛ!��	�!@���["O:$�!��TK �e�X�b�t���"O�31)I�t}t�
C��!r䮭Yr"O0XKCK]�],`�0+2I�R|�"O��%Jq���hs��H��	E"ONHi�c���KJǼ7n%��,��h�����[L�*S�]�[����63�!򄌧{ݒ�y�b�+_�4�r!BÁ]�!��ȷD���a!�1�M�� �/��{��$Z�n�(�c��eN����
.�!򄇾�d�����s����S!����������,�N�0eF�_�$5�S�OWhH*���J]֙�s ��)X��!�'�9ؔf��^�n%b$%�S��|z
�'�X���H�7�LY4D���	�'Λ�癃B�`iC-�'(�P�I�M�y��G�2�X	Q"��4���#�C��p<qH<�-O0��V[��`1�IJ�h`�O<(#�ʍP�.xH ��%M�ƘpI�<��A�� +3�R����y�O���3Ї�)o��JA���%F�m��'Hb�!�X�2L:!FJ�N���:��d,,O~���H�M�D2*Àp1ș@"O����,|Wj!������
�'5"1O:a+rnҵ|hz��s�K�[%��%�'^�	�4(D�_v5*S��Ѫ�?Q��S"Oj �r���1t߬I0�h���D4�iyS��	�T0���B"2;,����[�0C�I�\".(T�: �Jt��b�)-���<��,��)�1j�Z�z(8��ȉe����!��DD	[�d�X�#��k*���#פ�jWN"k�Ԙ[X,s U��,��G��9�\�C$e����ȓ�L	��-^`�hC�$�49����H*)�DB̤^�"0��F�Eᐙ������	;�����˖�L��S�? �hS��C�!�L�BcJ�b0�x)"OH̰G��*k	�I�i@ +��s2"O�Y��g_�&�L��.Q7?*��"O�\I�ʹEr��ҕL���C�"O(H�EeF�r��<S�e����i3�"O:�"DK�+��,�e��6s.�)�"Of�#�S󶼘��!z���Z"O�u�$�
�(�V�����"�a!V�'�Q����J�MY�ЛP���9
�j��6D��`��� y������ީmo���`�֏'���Dǻs�֐�뚇s�m�cO_=+��{b�!���W����GrJ�u��5�!�d��.���bE�*�ʉh$셸nY!��,.��ii���{F������Q!�DA�F�J��FG�c-���DJئL!�ŶM��d�rl�0oΜ��k߁"!��U)�.Azb��i%ֽ�c��j\��N����I=���N��3����U�U �B�	�KV$(i��РQ��q�PI�.��� �xb�r���Oi�\;��D�x�*�!����:�|��
Ǔb�$#<�����{�ِC/��,9PK�MZP��p=��ƉmW��e+���R8��M�IY���Z'BM�֢W�iP�I�w���R�va<4��Ȅ��4R�	�B ��e��X�F]+�x��ڝp$@$P��_�7�-��e��Q�!�A�J�<�@�ʍ�s'hp���j��'�l"=�}2N�!,�E��*@]�riҏ�i�<!�흀6Ұ���!� �J1�BAc�<)&�"L�$|I�/P�]�0�E��#�O���,5�6qI�u�њ�"O��*�m�5�vA�	^\��"O6e�a�G�����'�0G����"O�D�7��4'V�����+3EN,�V"OH�� I��+�XD���IC�T�#"O~����=O8�y`!�JA^$@�"O��QcdQ|L$�9FaQ+F�L��"O�@�>I\�o�;&���"OR�I��1���`ѓ)t3�"O�5+�d�j朐�o�b���"O��4Hʶv� ̈PHÝ~����"O�a�#/B�h҈X@G�Ŭ��P��"Olj�G[>��I�"ꏕ#�6hj"Or̓EjA	���5n��!U���"O1j�)�8X����	 q0ex"O�Lj�#Zbഝ8ecV>a�pK�"O�]��
]B�x�#,,^x�P�"O�A�,�+(ɚ4Cփ[�OƩP�"O�����3{��+�)*EN8���"Ov����?}�U���0?<PXw"O�d���� ��41&��:�P!h"O�Q8r�0MpR�WX�M2 "Op�!���z9V�JԊ��c"O~E� �˺T��y�e��*�ܨ��"O���4��s��a�W��5'��"O�����^.$ ��+`���:��Pb"OXԒ�m�]�1�q ��2P��""Oh��Q�˵'�>�A�V5p��d"O`����T jP�槆�,9�`H�"O\��ñw�����_3��0"O�H�
A�(Ęu��62lB7*O������w|��K����
�'P��HP��{Ti'IYT�&-�
�'C��K��].�ĸ��QM�%9�'����G�d�t+e]67:ـ��� �	iE&�L����n�4/���:W"O�GCU����qU.د �~i:�"O�TBb���U|�(p���+���"O<`+cC��3�"��Œ
�f�4"O,��gG;�v�S&�db��'AR�'��'fR�'���'���'r�H�v�"Z��%�KB��E� �'�b�'e��'�"�'5��'���'����Ϙ;���d��_"�6�'IB�'"�'���'&��''2�'u]�$� Y|��ps�:_
l����'2��'D��'���'a��'e��'?x8�"��*R�$��mj��B3�'TB�'l��'��'+"�'+"�''v5�N�`F>���@�H�8�c�'|��'+��'���'2R�'�r�'�8�#�OO4i�`��p�ƨ/�NL���'�r�'|��'�"�'��'���'�j�H�*@(=��%ke�U5!<@���'��'��'q��'���'b��'���a���(��q� ҄B��[�'Q��'$r�'���'1��'x��'��x"-P�b�`�3f+�?X_��p�'�"�'���'g��'��'U��'�����l)K!4�d�9B�XT���'���'���'r�'�'�r�'�(D�%nW�,�F4s�i�66^��rS�'�R�'���'���'���'T��'�dT2��Vs�]w�ڗdMn<���'7��'<��'�"�'���z��D�O���EAӥq{�a4�&i2�0 �Hy�'��)�3?�f�i-$	E2a3�1�n�:+래��A��d�ަ��IG�i>�I��MC�C7)��� dƑn%ҝ��GO�`�&�'R�q�iv��O�@{u���?���u���� g�8-9fU��Û�H�
2D�(�����'��>�{q�M�3��Y	�g[/k3Α�0ɉ6�Mkr��w̓��O^�6=� X�Wg*F���c�/%�"r��զJ�4�y�[�b>��tc�Φq�W~�����3z.���S�D�?�F͓ޮcD�>�����4�^��ݬ_���qM�J�H�X�葭^,�<)I>���iX򽓍y2��/b��2�fU4L �US#iK�Cb�OЭ�'	�6M��U̓����74I@�q���^Ƥ*�I�v��-��9 �&6WNc>�h����;��'X��1�<(ݘ�e̴F�����Q�@�'���9O iҥ��B�l��%VC��m�'l6��R��>�M��O�)����}T���,�Ӱ(�'�z6����e�IZ�$�nX~2/2��<葠ݦXy��,N#k �ģ�C\_�T��|�S���H�Iڟ4�	Пt[4O%r�!#7"�ex6\S�G�by�ӆ)S���O���O����䃯-ƑR���HaR,�' ��lg�8�'6�7-]̦]����ħ����@X~9g�,!T�HqdΖ^M�(��n�'����8G�l9�d��a��1���T�5W�0�R��
t#��C�6�v8툦&���S��!%{$�a�ݪU����r��:K�`���Ѝ&���胰�]'�;�m����4r�L��%�
���"H1Ha��Y��Fq��*��Fg�$u��̅�j��d1��nh����ǆ�Dy�բg�X�@�v��2ǐ-_R4��Ԧ](t�ũ$�ž[Pf�p"u���U�|Ά\*���3k:�8��h�{��i��˛�zSL�j ��*
��a�m�4���	wDV�0?�P"C�Q�K�*���N:�1���
��MSq�ƀ����H�(8J�4�UhN��'��'��'�I̟���e>)���@	4�P�J�+��f$(�|5��?y��?���?�e�d<���'x� <�õ�
e0�g W��26m�O����O���?q ��|�/O
��p��Yc�03 ��6!D�
D�v����OL�d�O��J`��Ǧi��러���?1�p
<>�BDa�)e�\������MK������O�b65���O�i1�}���ښ5�&d��,�?P���#�4�?Q��[FZ�:2�i�R�'a2�O����'`��� 茥��H�C��}U��ϧ>��$��������|�H?��S�Q��E�1ݩ��`Ir-j�\� ӊI��I��|���?��Sџ<��������˄{�@	�s��%^�zi�b�ȟ������@��Qy�O�O��ަ-�z�h/�S>H����3Z&7m�O����O~lQAB�	��ß���ן��i�i�&%^'����$�;��U�GKrӦ���<ɷ�(�)���?��O2�*��W�n�X�`�'��۴�?��@�mh���'��'���~r�'�289��d��\�w�	'��E��O�4�`7O@ʓ�?���?	��?�
Y%,1`�n�ѠgZ�dv6�Pb�i-��'���'ZL꧉�$�Ov�� �36��͛�@ًf>��(V	Ea��O����O2���O��$�Od�	�ئQc���!��Q���2��};�*\��M����?I���?a����O"�B ;��T��3��Q@�	�S6U�&�g}B�'9��'���'!D��.o�4��O�٘Ud�*�:�5� ��r��ܦ	�Iß��Qy2�'���J�OB�����H3{�$X�wÌ$y$�m�ퟄ��ğ��	F�j�	ߴ�?���?A�'K�Vܲ�e�Io��(T떞�Ȱ;��i��V���I2"A��۟����4U�R1�B'Ǫq��<��hW�iwPIm���ɢ<Y ��۴�?��?9����+�J�D_6�Ҡ�R�ԈāSS�d�ɤ4iT�Iݟ,���d�~�Ua�h��}X��D)x}�y�aɦu�A#��Mc���?A�������?a��?A��5
� ��U�� b�Ġ�@#?}�v%�b��'�i>�&?��	P�����%P�J��81�����
ش�?���?�3���<���'���'���u� ���)�ŀRi������M{����$.8��?a������I��� L��ဴ�v� eB o~�ᗽi�r��7XJ6��O�d�O��II�T�O @�$+ٓh`�22��.vle�W\���V r���'���'j��'�bĈ�*��U��S�
U1��@�vX,���ba�H�D�On�$�O|,�O��	ΟdcTP�Ј�cW��9�^����#m���I����I���	����I�������M�v�� ��IbB<S��P�/Z�]Ûf�' ��'��'	�	Ɵ܁tEb>1ص'�Y� �W�$_�U!�F#�M��?��?a���?�" �HK�F�'��hV0Z�X�0%�f��L��F
$)�.7��O���O.˓�?�/��|�,O 5���\�=ef��OI�G�N\Rɜ��?q��?q�[#�y���o�����?�k�d��C����T�B*�
�B�1�M{�����O�g<�����<�禝�pC�#Y�����u�� ��Lt�l��O� KP�HզI��ϟ@���?����� S�K�Fk�a��h�*ơ���O^�ӰN�O ���<�'����;�
�� H�|��� lO�7�� ��QoZ�� ��џ �S�?a����8�I�B�,�S�NߜG��q��v7��Iش%>����?�)O�I.�I�O����b@�x�)�6���B��U�# �Ʀ}���T�I�q�`��4�?���?��?��6��@�!��$ �pCN�l�C�I�^�F�)���?!��? ���MӗL<hu�C�y��K��i��K�>
[H7M�O����O�|Ӗ��O���@�V{�
�G;_?6��Ri��&��,u�HȞ'Tr�'����'�R�'&�Y7E�,��փ�(^LH�Q	9�t� ��r�x�d�Of���O�T�O�I��"/�>������Ǵ �n=�"��(c���I��H��͟8��Ο�'���J��x>}XGnD�RJ�������z�c��˓�?1-O���O ���Qy�	�'�]���Je����z�6��O@�$�O��D�<����F}��某�6�[),Aja��+��t�&D#�Mc�����O���O�A�E�iih���Q2�l��G!��.�jxR�4�?�����d'F��p�O!��'�����'��ʅK� t������,����?���?�ש��<�-��d�?%�À��hb*)���J�:� �|��d�O����C�Ǧ��I������?���͟���X�|�l���(fh��p斈��D�O)�h�OVʓR�b�ͧ��S�<�x�5�Y#h10Q��K�)�z6-��}��0o�ݟ��I����S�?���П �	4Tt�R+m�A#o1f8@�4E+�Ej��?��|7Vͧ��'���e��75X���F�lO0��� I�P���'y�'Z~�zQlj�T���O��d�O����Z0ՂźG8<܂�
Ák8�v�i���'O��Ç�כ�yʟ.�	�O���T�L}vE+b�Y�7�l2g�7(8��n����&.'���?������b�V(���C��Q,"t��$jTh}�+׳��'���'��[�,�ai�"�aH���>`�M�Ť3s
�1J<���?aJ>�(OIs��ǫ]�:�:5�Л�dh��¼ty1O*��O^���<q��-��iLyN�DΪ#��e8��W�?��Iԟ��i�	TyR�9��$��BDt5���s֜r�"ƞn������	ǟp�'l�Us��"�)� �p�HF�#������ވJ,R]mΟH$���'6�S�}2ʄCB݊�	E�-��*�Ꚉ�M����?�)O�0�B�C�S����Һ��fF4o�S�J�G
fA1�<)C��Z�����-x� �M	5w<H�j��A:
��_��@,��Mc�X?��	�?���O��@��6�h@�g�'S�Dk��ii�I23#<�~�1��8%�-h��	�i��pˀB禕���M���?A���2��x��'Ĺl�q�9��.�'��)�b&s�ڕ��)�'�?	�oZ :�|Đ�-�
Gn�c!�Ţo���'SR�'P�(+t�=�$�O��䦟�cG%~�xh�@E�
3�1���/�I-
J
b���I����I�5;��5pS�ܩ���^�۴�?AE�֛_�'���'�ɧ5F�R.(��G!M�NW��a#cҳ���O a1O:���OF���<)B�O�T_�8r��֖	��u#�2�0���'��|Z�l�B.h�`	�H�>����� "Q�b������IVy�%Q`B��,�.i�'�n���[DG XUBO���*��<��{}� K.�x�f�7aXah��ކ���O\���O4�}GƄ�֖���4�	;�i�Eb��s�����7��Or�O$˓�F��>�`��@�Y��/<��ѓd�礪�	Ꟁ�'�V�Cc`'�I�O|��_��Z6^��
91<w���&��'7^�[��T?q�U�Vt��칀IF2>c�tAR�tӨʓQX��f�i�H�'�?)��E�	�!��@�a��3�j��d�Ȯ�T6m�<��h���O1NP;T�Z�Up�&��
����Ir�Fd��4�?Y���?I����O�,^f]!�cѦ�����ۦy{R�!�S�OEb�) ��!q�m��b"�t8㥚�2t�6��O��d�O��:���S��?��'i��q�؍d����Uk�/I{j��}2)��ۘ'9��'DҎF�&�9qU�ԉH�*�+ԥ��]�6m�O����e��?!I>�1Z���℆-*^�q� V6V��'�v)��y��'���'��6%�:��E$=��E���G8!B9�����?q��?�,O���dX���?q���Q �5
YV$� I�K��?I���?/Op�pv�^�|� ����GY�H�r�C��<}U�Q�vR�L�	h��vy"Y�px�n�~��-3* ��yRd�=KF�K��k}B�'���'?���>�i3ki�e!o����?T,�o�㟀�	SyrY�H�e�1�'6�cf�ڟ<��}���/H~�ش�?I���u�<'>��	�?=c�bW�8��S�cӃ)d H'%�	�MC/O�
������4��V`*.(��aCF�\yf(�a���M�(Oh���Ϧa���h�d�`��'�\2���[�4��̛MT-R�4��dS+����3���8�2�;�G��J
C ��[֛&��rl�6M�O���O���T^��ퟸ!��ۆpp� �խO�z{��O��?��(+�Q�c��1X�֕@�F¶�:���ig�'K�#>Y��O����OV�	:O�X`K�K��Ј��>x����O����O�	'��5��H��KL�p�@��g��Ҧ��I��h��J<����?QL>�1Gd�i�a��-ivI5i����D~2�'?B�'*�ɛ<`���U���X�dY�P��F�(a�PHٺ�ē�?�������ɂYta�ՂP�A6Ω��	N� �b���	�\�	Kybc�`擗Ci��&#�{�j�Ca@� <��듛?������䒹XD�	VqD�0ңĤPݖ�I'5꓎?����?�)O"��r�SQo�\�S���H�bR�['"p4�3ߴ�?H>�/O��������s����Ȟ{<r����
��'�b_�d
�����'�?���c��@�#OH����K�H/�qבx�Q�<�g#=�S�����n�@1"e�(.<���4��$Ķ))�l�����OZ���@~bK��v�I�	����2bԎ�M�)On���)�S�*:��V��0�0�P�i
	*e�7��F�l�oZ��p�	ٟl����'�Ҳd�|��ѻ���sL\PRQ�yӨ<��)§�?�3슣XQ�2O�1��&@�]��6�'W�'[<��3�4�D�O��d�� ���Z�~T�hKT�́
�n,0�/4���[�b�������I�k{�uѱ�E�'����3S��cݴ�?���:&w�'\�'lɧ5�a%y[�!�!�1@��̰�`M����Ô�1On���O(�D�<�Ј��\
2�%w�
U���B�X֑x2�'���|"Z�� ��hB������+�k �1t�c��	����I^y�F�'/��Ӕ�`�4A�=G�lA�ޑO�듈?I������Ҷ(B���6��l��Z3�ĭPW��;&���?y��?9)O輢��Hx�ӱ3jx�󗤏 T��@��-�bU�Y	�4�?I>�*OF�T��_*\֦�a�@�D�`�!��"���'��X��k����ħ�?1�'L�����=2`��q�i-:Ɛyd�x�^��Q�.�S�4�L�\�X��G
�D|�hP�M#/O.�C�æ9
��B�d��4�'��!�p�8"\��c��q�ݴ�?	��Cq�������`�sGI�,>�8a�1��aݺ@m�A4���4�?���?��'O��'\"'�!q�	�`��!�D��h]he�6m�	5yN��3�ɟ��6@�\�����GC�.� �u�B�lZɟ���؟0�"���?i��?!��4,���sA��[[T���aH"j*�O������O���O�s�<�|�&�Kằ
0��Ʀ��6%x�%���֟�%���5��pȖ$R�I}^)�.�K0�(W&�cK>1��?����D^7��A���=���� AA�u�T�3�K�\��?IK>Y(Ot��mÓ}~��A�ն=֐� /^�1O����O��ħ<�3���B���\z��I�CȄ*�����6��ß��	p��ß��I/5P��.=m�$��HLЕX#��YƼ�O����O�ĭ<9W)��fh�O����#7f�ögJ�%UbUJg�k�P��$���OR�Dԗ}���$*}r�G�4}��o��!��@X�G��M����?�-Oh!�"#�Z��ğ��S�4�Z���d��U���a��<Q�h�N<���?���Γ��S�$� 8 �!tH$��Q'�,�M*O@�X�MZ�ub�������T(�'Ȝ-�Ƣ�n����3(�
����4�?�����p���DH(H��V��4��AAȓ��M�P)�3IЛ��'e��'���f:���OJA�EB�7� �+25zQ�U
�ɦ5r�a��&�"|��F�X�Sj�*a�	�*G�P��4��iRr�'�RGޯ�O����O��I�+�����HT��X���j�66�!��:1��?E��ܟ���U�) ���g�pt�u���]P�lZ�� K��0��'��|Zc>0�!�/	�5#�*��۶V���x}�#�*D��]����ܟ��IwyB,XrF�����6?�`(�8; ��$���O��D3���O���K ;��� ���8;݆ (�G�f2�	��8O|˓�?Q����'z�P�X0����`X�ṧ]-S�zI�_�$����&� ���l�"EX��t0W�O���G�
]J8Xac)O�_;���?���?�)O tzFK�G�; �湘0,߿N|��Y��.)��J޴�?qO>	��?���?�M���7#��}(d�3��^�*�T�C�y� ���Oʓ��ۦ���'/�4"%� �u�hߛ5�P���Ǉ'�"�{ �x"�'N�)ع]R�|���M`'�7a
*d+�����i��1V|D�J�4+��S۟����D�=��{GƘ�A� |b�-B)����'�2�5�yb�|��tb	�u�έ�q�ۃOT.��&�M�/E�?�v�'�r�'y���'��O0�c��E�o���(T苝k�ZE�dWܦ5�b�_ڟt�'��"}��?,���ѱ=�dBT��C4i���i%��'�"j�*�tO�d�O���J�X�9��9 	�E���[.Y�46�6��H�C��i$>9��؟��	-����0A�9@-��UރQ��|�4�?w�)��'�"�'Cɧ5&�>+��%�`%Y�d?�D!d́4��D<��O����O<��<�F�9xsR��𤑍=�lt����2,N�C �xB�'��|R�'��]?}��ah�����5cY�|&&����'��	�Z�yIs!إFժ�3e����O+H򢇒m��q�/T<-p%Z�'W\<I���Np�\�n�-N��K�{�'H콃b����M�c��*y�F)@E�<&2���IA�I�qS����E.�\2e�Y��<�;��0�rX�$D�>e�rU�rOL�}m&�B���yVL���T�"��t��q�"E�(B>+�"\[Ra��j{H����%�
��`A��f"q0� �P���	�Ϥ����o]�?����	��I��ǡn�Q1����?��:��o�-:H]A���.9��6-�|:)�҅��k� 16�A�F�<_ھ�3�>���AN�~�;`^:@Y�!�����pu��U�	X�x���3i� ������ �N|K~ʱb#L��ѐE�9	܌XA
�n~��'B�|��$H)a}�d���H�;Ƞ��a��ax��|�"o�W��$q[q��4���Z��C1~@Z�O\���O
��7E�����d�O����O�Gy&���Z�|��PB�UʬL�FE�;�F7�յ�l!@L]Ņ9u������	�YH�)�!��_/x�*�ق;wXp�޴w�t��Bj��}^�i�I?%�d�i���3�,uA�l�0�� �RW��4?94ȃ��d�'w ��I6��i�S剱�~���'?��R0&�KR�j��/�>��OZ�Dz�O�[���-ʭ(�Z��I�}Dj
��	�@��T П��I��I*�u��'�R:��Y�b�Rl��5&iZ��p�."J!��Ddȱ!�o��A�kJ*ΎyHqO
رq)���@-� �!��\27m�$��I4�O^{�'_�=2�*A���\}q"O� ��G��b�^���^�.w�0f��W�>�ɛ�i@R�'H�AZ(
�8Y��c듋Av�t<�'��as���gY:��$��g�l9����2� ���i$��'��,J��Ӄ$�M���h	�.�X�IˉSx��Jԅ�Q�ٚԠ��.�$��--#��!�÷sԣ>�"N�����Iʟx�ɯ kh�GJ&K %�A�P�4*B�'�����$ ��2�恮�M�# H*B�	��Ms�A!��gN�$��q�#��?).OB]�$�Ϧ��I؟��OҖ�@�'�(�°h�Q�J@�"�:8�.YQE�'�I�I��T>�����L�a�*ՠ'A�Z�@��O����)�S'MI����!h�8G�)�'E�8�ɧ�Oτ�pˑ=36B5�����-� �'�@��]V�#�J�=�A��w��؛֡=.}�t	�L} �c�B:�M��?��=0��b���?���?A�Ӽӡ w�fD"G�D��r�T��*MЕY^���MA�hLb�$?c�8�2k�4Ka�������R�֠�*�`�_E�����CL�>mN��
3C��?n*���g�ej�1�&l��؀۴�?�lM:�?�}�'���B<lx����J�|�X{�NJ�b�)�'���9���0L���ʛ"���͓�?9��iC�6M(�4����<i�f޴h�������?ʬ��aC@�(ҳ�G��?���?��c���O���x>]`�׾��e�	�E��b�A��49����\�e6�c'�ٴ&s��s���w�qv�Fu�<%(�Hƨ}:���A]�p�'R+����Ǎ&{s��\�1��{S�|�,\9�ƔZ�Ϲt.v��ɟ�`����GpabK��(
�u�#ð=^��-�r8��$�z�A\�\��*A:'�&�K�2扅�MCO>A �� ����'��^=
�4�����{Ty�K/+42�'t�����'�B5��]���$N>��$ͩ>afM�=��j�HA��8sbDWQ8�h�]�[D�j�J}¨O�7� Y+��D��.Hj'َ�p<	t��������4�	3 �B��c�=��:6�ڣD���'�B��S18l�VNů6q��p&kXP|�#<��4�to��	�|��a]3;��)@��כ{]�}�	Wy�j�_h�7��O.�d�|6�1�?��G
�'��5j@U��2�o���?y��p�!R%������G� �*���'cO*� �I�o ��U �%c�d��OP�Q����[��I
7�E(��#}�ԄP�DJ�6/v� �\�d�59h�e ��� R���6���fI�g��8�5"O~A3$���N�����eE��y���'[�#=����5r|	��(��v��j�V�gx���'�B�'�<�яM	m��'���y���'m�8��#���J`���$i�hp� �>�D��,Q�B�HJ~�<7�X�'���1q�\��!�ub�C�dq��OD*�q˂�[3R86��}��*����d�~��񧨌*3IL�˔+O4t��m�"�M��0���|�ʟ�I�И���A����� o�~���F�'џ�����6��a�7A��pP�.?9Ǿi�H6m!���|�,O2-���{�ܭ���X� �6T��%�_��h-�O���O��dZź+���?)�O=��ը�f߼T�����p	Ցc�j�[��¾od��
�\A$��^�3Ԉp!텄?,b�4�Bq6�롇 �%����!8����GL�9C�L���
T�0���E�O�oܟ��͟<��ԟ(��ԟH�O���A.T9x�$as&�A��&!	���*�F0��º!�x� �:WΖ��<9��i�\��c.]>�M+���?���J1a��HP��!HĂ4��
�?��;�4�r��?��O�h���M% G��G�Y�J�ڄeɎSܨ�p���������}4џl�U��J��p��[�t�m���?��[��?�
0�E��?�>AD"�]��?aМx�"� ��S��YR�X�EH*�y�$F?e�*9!�`ߍ}�X@C��x"�y�J��C�_(X�Ԁ��C�2=b��D#�9n��T�IM�Tb�C��+X'[.��s�6�j���DA���'7V���'�1O�3?A�#H�~P\z�J�0���X�B�S�D]9J��?])���4Z9�� A툎�n��E�&}r��?	��|����5@G����1!&����:�y�� p�9��b��-9�H���7�0<y��ɚ�N���ə1`MA2�r~���ش�?���?�"͔kk�r���?���?ͻ�j���G02��Mf�]�
n�	���B�	*��R��'A ���F�����K��˱g�eU�0�U,�Y$�P�ǋ�(.>| %�'����Fm�g�<�1�a��7
��x�A��U�  �K>A�A�ޟ�>�OĹ #đ�eI��kVd�J�ܑ[�"O�����9Hd�0;2�6���B�X���4�|�O콑���XQi2$�B�X��O�u��,Q�E�O����O���˺s��?���>���H2;�H�H*Fl�z�RD����$)���'�����"�*��E�w���д��
m@n�*A(�B'�U�Ӎ3,O��BEM5~6 ���fT��Pq��_)6�"�'�06�OV��?y�B�L=����� z`^|���5����͸/К	#¨T ��*F��5_֒O�nڿ�M+/O���p�R���Iȟ�Z�TX4cY5b �&�͟����rI�%�IџPͧ9ъ ���Pƀ��ȟ���YsY����i�5\1��%Oj�pu��x9>��J�!�"^�p3l��Fg�A�%ߪ�p<��g���(��4^���'���b�(T����QD.Z[
L�0pZ���Ir�S�O�b`�	� 2ʸ9�ӯU�RoJ����$-��|��iߔ�#�ܦ�R��R㋮R�֤���'��)K�uR�������v�d�C�}�"�^�U����犟5�T���0ox��'h D��I�bR��u!R8|�v�o�|�)�z}���.�\��s��00�8��>�a2Z�Xѱ�T'TY Xz������O�|�CG�^�pP����\2�sM����Ol$��?q�Rޮr�ne��@-R�X���4D���*F(Ж�x ᐾhINU��4O��Gzi�^����f�͹׉�:�y
]#cL�1���w1��RRN���yR/ ���@���2�� �(C�y�!�"�9Р�T�:q�"͍��y����F��QKԪ9ڹ�q���y�I:�:\�҅].�I�A�3�y�j�.7H���鈋N�칅	�(�y�*S��䋶�D��I�2� *�y�Ċ�B�4`3�ۉ�BX�4A,�y2.~�8��X"��(�I��	
萄ȓO�JY��@�2<8��7 �*-�ȓۈ|z�,
$� �gF�Y��P�ȓ =QhL��0r�ː�@�'h�A�ȓhDIB1j�/&�����49����ȓn>h�4`�<&&
������~�݇ȓQ(�p�dȋ�~�����6b.!��S�? ������p���A=�l�"O�Д�R*W^����ǘm�j��"O
��T�g1�x�a��&R9���P"O�=�gT�}��T;�E!T�93�"O�쐓_4t6()��&	�S�)�"O��3�6���J�E��c��XU"O��Ì&���"4�$��]�T"O�U���P�"��
%���U"O.�s�FMF�� �$܍6�����"O� ���ȋ%���b���A�x!��"O���U�����9��aJ�"O^�2D/ f��y(�OA0���"OJ}�S%�;c���"U�K�"O��`��2b�%B�%�,��t��"O��r��~ݸ���(��p"O��墖#_|�Xsa�υn�*��3"O,\;���a�Јc��4�!9Q�҅#_�Ԕ��͓+q��i����g�8U�Z Y0�P�FY - �MZ�O�v�Q1��E�"=���X��Լ+�n1{j`@��ɑ+�a�w�ǟ��$k����'hs�_;=Әu%�?k؅���Nc�6az<��@ܱ>m�Ma�m��C�|�b��#[MD�Ѧ$uX��{ �P� �h,t� ��'wI:P)X�F�,\+��_�v�`akY�:d�
���U�j���B�Q6���G���P��[��m��ggA�Z��ʓ84��O&xe��S%6���"�7�)O��!�U,m�nMV��� }���&�	�$hD
�3�,u�m��8�#wM�a���0qͺ��Aōi�gy2�]7�8��c�7HthrȏZ���r��û{�\�r���tjv��/�y��̕�Eq��Z�5,8�t��L\x�$Ucp>u�SǊ�i�axb�һ2C�\�j�� ��	��o��v�Ĵ�?��&�����R!���|��4M%ҨjSjP��$��`��8k��A(��;k��U���5~b� ��؛o�PRA	�*u��,�1{,�e[W��8qF)�Chv��êK�5�X��o��]L�T�a ��:d�'���#0��'��*V&ԑw�Q���g��q�'�B�u�	��h�u���Z7�(��$	;�f-� �4|��I��W�c���o� HA2H��#�O��:�"ո�?q�'3&+�J�G���0` � %1��5k�rj��{��/�HO��.�b�u3�z�1��#?_:��f�B5�~ʣ��-1�h8�q��?K��Pa�>��䆸aMȭ�1�źS�b����,/��PC�}2�۞sTP4#�
�,WkN���*�2s<�8EM#����|L8s�CI�q������>�d�)��r�KY�1z������p0��
~ώѹ�U�y� Kr�Y^@�����`^�:���D�x1��:�)�	ݭ9����(�8�@A�A	�3L�1�>Ń�h�2x瘡�1�
�<!$�?)w	R�j1.�1QF�+\0&O�W����Z3%��9R�"}���Ŧ�yP%�@'���#[� `�GբP	p*�!�2Gy�'S  b��j�ix�r!�H���H�U�ơ��P��"��tX��1+O������śkf��KA�Tr@Q#�Z�h�dZ'F�mV�ȗ)��Z�(僤J��y���r��y�����{cv)�� C��~b�C�m�O����;�v(��(S�*:�"��F�s�� I�n��*��UCQHӜ��'�TAU@ì}��:S#�4l6٨�П��BB+�
�P���cJ��S�����4{������y����$B�,��\:u�0�#�(�)7<"E�V⹟��%�		L��]������6�yx��  �HlA��Л- X�ɋ- G~������G7���S�;\tA$�\'Q��Txt�ڎ}��O���t@�'��	`?6�c�@�,�<(a�϶����rj(Z@~m�Ê	���xR �6?ѥ ���eTa�OB����`�M?1�&ۀʸ'���j������ [:�:�	d���16��f9n ���N�W�*�Bb �9#�c���I+�Uz�ԟ���rr�9u��	�f����t*��&��5�O��Ҩ*b���3�F�DyBG�/��pB�'�	�T�0Ŝ�aDp��>1�eh��ʧzc��9v	2f���s`��"7��ܨ3�۾#�!a��^��u��Z�����wdR���ݴ�"D�,�z�D$�E&��⟢�J��C]H���Kؔ  ��k�T�C��!�%~t#5�K!ӂ&�x�U��%K���w E8
�������([�L_�S:�*%
��PT�ۏB,tɺg�ۍ��3˓�6�RX��I��;����C	�}3<�j�#�e�S��'O��rlG�c���@�4��U�L�����)��� �>ڎ�v�!�I�a�txH�'�Q�|(����^ܥ��c�[>���{+����H� G��-�6BY�q�@���˘(
D	Fy�'K�,�2Ji�a�'.B�|��`�5B>Kh�''�9b"5ˋ���̨��(R��
�ԵBKφc����>ѷ��r0΍��e�e���K�OM�ɯ5�����9\ೲȕ�"bz�t�#<���y�ᱶ���b�z�X�ʤQ�u��N5:�4Qt��RkB�h^:M��
=N�)�o�g�'p�)� P|�eX^���@W���n��>���N<��2F-�O�I�#�|��������W�Tu;�=Y��`�	m�����ê+�r5�&���朱�7�0|<��f'G/"�Y�d�韜��3��y!^�|�N�K�}[B�PC�V�?ɋ��S�dy��p��IN�9 A�8�t�(��]�Js���,�&8c�$�$a��',t���S9HT��K���ɖɻ,O �<�P5caR1��.S�%r.������b���23�89{!A֗��� �fXl,1����W�d|��D6?�'gI�,�Hp�w�HS�h0�Rs��&�i�dn�&z�-k�m)|�OBm�DFӆ3kP�J�	>
��+�V�'|p�Fy��LT��H�="�HB4���?�ŀ0�Ti��a%*�sj�<���(ʓsuJU���,wδI`c��%���8S�D�![��p�D�$�M��Ið��Y�ؗ�Jw�F����+��&�\z0�[G�D���)�<)� �$f��!ZyzD�!KKF&�0�e��V�Tuv�W�^2�eb`ʞ!�~���<%?7-���#TJ� ˪��o��P t��`�%t	",OB��A��Iy��:�����.Ջi�BL!����~/�|2���=/a��#[B���/OR���"�4��'���po��{
l���F�d)���<�-Od(�^w��!�"[eF}i��AVnڊ1:�1+�i> 4��£!`���� ���6��?	R�<�m e���s����	�TX��+8i#r!�-��1G��e::��7�]���'x��j��e~���]��Iئ�h�#�����	T�7�!�Q̖�f�ryid'����<�|�U�f�%�5.�K�> ��Ƨ<��a�V�cr��'�}2��<���d�f���' �����¡V�,�D|�!�Ŝ��d�a�͔'� !�#N�B�pӄߖ*�LŠ�Ăm�0��Y�H1�'[�<b\w!V�k�g�Ob��j�|Z%���T�p�h`nNiҰЧ�T'���T#3`qH���O�X�Q,O��ʳa�!N0[�F������|�6H��5�"��`�峟�3*O�t"[v�rh��,ߓu�h������' ��`�٩,��tȥ���<���M<is�ҫ�bd�%J�^�ku�s}+|�'v�-Z7BW^�iq��vw*�h�#1fkj��1��6�@�蓇�f�ra��F�Y��m�į~�Q���'��,��dU�'�j�� _���;N��J�!,B>&L�s�����%�ɜͨ���D
yrJy���A� ͋��"�S��H�1
P��"%e����j�^��/K�2QP���O&���bݼ��睯}y6�#ɠ-�\*���ڟ�D{�������@�Bז�@�G˲�>��}��҈O����2
]*�n]
?�ē;�N4X�*D/	'��h�$W�J��'=Q���Kҩ9�� �$�E���18������!E��+�q���18���84꼰��!oEy�H���Sc�IX��]�a��z��!}���DC���b�#	�~��db���'q\1���0�0�(Fv�����!JVXc����%���0�����31�m��T.H3@����I �lGy�'s��l�� d�Ms �41U�(��ièuߊ����4G��@Q�e� ���|R��'K�Jh
�E��e�j���R]��>��V75�,�(�!D6.�,���9�|U�'&�2�W8F�"�sB)Y�d��)��'8�08�ԟ�8��$F l|0Ud��0!H���	T��)�v�X���	
��1���B�Ǎ,'�$�U͟t�ɧ�>�ĠC�M�>��q�#I�x�P<�Or(�4O�kp��z�/��X�H������6L�8����ҎWvV���D*/jI���j�	
o�Q?im�"�N����Sx�`�n�9)�-���> �8��F���f�<y���ݼ`�GM�`.�l��
����.����9J��
�I�be�D�	�� -�����e|�4p��5|L��ց�3B��?�
�V�2b�1a�-؃R�����*Đ!�}2ԟ�0c�%ȣh���פ��P}ؑ���̱_BQZ���=E��
я�(:��!��%����W��N�S��'w4,R�bĔES�	q0��N�B4*OL["��,SD:`	��=Mԥ5�	�[�>���%/�����]It ���#�Ɏd���T>B0���ZPi�h�r��o��X��g����O�T�Eҗ�~�kE�{0����U�h�����B�6�V���=��~���E�����?��c/P#Dyp%I�Y\DI�'<ʓ$����O<���	G�l���I�m쒴i��*rbe���O(x[�'��Q�#[�|O&y��'�Z��������l�7�L$`u���FY�c��E�Q&�Yp1O�D�U.���E R��zᔔ9��?�Q屧윭/]0	�s�]�o�F]��A>;J������~g���d܅j,�b�$oeL�1W�A�,��\:�}�-Ӻ�?�O�64�4+Z�0&��H�r�Q��cS#3�g�_��HO��Xe��;�Ƞ�qĝ� !$�Q��R E`���`�*Y����?E�$�߯5e,2Q<)&Huש��'F��qb��??֕�H�$q��JL<��J�R�C�OB�X���pa�w?�b������$�H��By�4���(q`R�ϟY���5�Fq���QRf'f����a�.�lE�_8����'I^tX���D��UH֭�zB���O�����K?Gt��A%��.+x����� �iQg��
ul`�Aį�m��Z�.�v�'+�Gy���K��J ={��`~�jR�N 0٫ ʓ7ή�<�; ��hV>���b%�2{e�0�'c�+Lᶐi2�'�ў"}�7�����S.CjY�u,���P㟄R3(

X�.M;�L
H����(}�KǠ�0�tMI9t<Q������$"+��D����N(���K���ʓFF�%~�9��?�����J�<Y毑�#�����"X�i�ȗNVc�IJ~2��|�V�4��X�$E���?�@�7;�`H���t��4�x�'2��ic�;�����bU�9[f��'ˉ}(<9�E*qY"��G�9뎹C��G�S���-�/<�d DzZw��q��y��աZ� �$o��s��Px��@�F���5K\#I ��1ď
�Mv�(�>��o������1$ *�� _�	�R�rq��L�n����s��3�H���Z�s���ic�ߝjOE!ťD�VQ�֓}�v؊�DM���qi�aj<۳`��8�����=,OrTY�I�r���S6�L3A,��A�>	�d�&XI�V�jK8�XF�v�V[�)-��������d��c�O�ⶪP� ��RS��$K�\eB m�.+
�	
u��<��\d@$5�$]�b�ֻ$�tT󆣇X�,�
O�D�ծT9oiz�`��Ow��/ʡ��'��D;��M�t����&��Y�K�x0�
2U�q�F�)dƪ�%�<�	��p�B�	$F��'3��6��g���\8A����o3D�9wퟱ<��)��B?ZXR��0D����ʡ*�x�և\ s�� 1H:D��H��ݙ'� C�Ř+B+�=P'�4D�$�$iU�/�,8�$��f����5�1D�ġ�쌜\#�{���t���E�4D�4pg���+H�9����3�ler%�3D��&OĄ/¨��`E�`?`�c0'?D������=�+P�P;8�F��A<D�����
J���X4��i�����d;D�L�3KW�&��b�5@�p���"/D�,)�G!�J6���|�li!p�2D��b��
;�"��ee��m�y�6j0D��Ag���N�1F`Brg���N9D�DI�$_�'WF� �N��HhZ��3D��`��{\r�`��?G���eO3D��{E��YJ8UxDh�*"՘1R�3D���`'ƪ�e;�����#�h.D�8�wk��\k�Z�ilB���n,D�@����,�`����zpDjuM)D�����4���:tM�����b�+D�,�'Ȍ<e�Xy��.+.�+eO6D�4����5SC���!��o6 ���5D����g�&{?Z�j�Ƈ,R�)YD�'D����;����ŒnĦ]��m)D����/}��p���?(>�e�'D�����]�:	{�a�= !Ā�C�9D� ��M�Z��H�O�#j҈�P��,D�p� ,Y�;Ұ	efAa���*D�P ��`��8 �`��qu`l �i*D���`��-�N��eCɶw ^Ļ��'D�x�BĘ.[��=PD`�4�j!$D�tS��Җ D������-K9��t5D�����(	��%�w�}��$�q�.D�4�v`$i�9	�Z2���\�yRk��:��q�	P0��ez�섉�y�.�Z蠹��͢q*d|+��%�y��4d]�|і�� n65(Ǎ��y�g�(Rn��F.?m5�Q��%�y§��mF�T� ��\\&�Jv��y��$o��� �)V�dS�ń�yB˖/pJ�:$/�(#׌�i-ۅ�y�L�����2נV�m!�	�E��yBg��s�ώ�t�l�dĕ�y�$$
�1j)ũdb�����N��y
� R�y�[�!�
�A�IW��"O��h�4z�x �r����4���"O��bu' �.�aF?w���%"Oj��"P�:�!�g��F�E"Or�j��R,}Db<��H�|I�=0"O�TJ �ѻL�����_a?�\IW"O^��W����Q4��:e>�P{ "O����x�2����~V4J�"O�=ɇN�/5���2���5
U���"OLq��I� ����΀�9L���Q"O��LO�1#4�`1D�m�J�W"O�)oG�!#ז(٤����"O,5�����-JC�"s��f"O8-�Dl�*|��
q ֹ^8���"O�Ly�%J�s�I�d ޞ
�H��Q"OXXN�(j��}S OPmKlP�U"Ox�Y��-EL�Uq�I�I���u"O��qf��)>P&t�C� _Ep�R2"O�-�dd���B%sECC@(�� �"Op|ke�ţN"0�$�U�h
�{"O�H�4��;)�,���";g�Z�"O�@���h��r�! eKN8�T"OB}A"Ѿ>�̹�� [;D�1З"O����QR�D�a�H��cD�i�GO�9ZS!Λ S��KQ07�bPP�"D��9sJ�	��U��n��G�4pc��2D�ШuO�7'N8�b�M >-,���o2D����˼.c4��voR�XQ@M���/�O�˓S(�C!�G�~�>��"��%H�ڡ��>�JI2w�ʥ`�(�4��a.$��9S �B�c_/fꬒ�B_���sJ��1��V|��ٖ��%�*]��uL:m��K�= 1� b	Q�o� �ȓZ��hj4O��w�]��em��'a~r��T'�a�A�*`R|C:�y�`�r=r���GQ�������yP&�
��0�Uu��F���p<ы�$߿'�l�)�o˳��U��۔�!�@�5t�*UN4F�"�ci��ey!��K�D�:�a� uRPY���-m!��?��D��A�j\�!i��-R!���xL�r�\C:��"A#ab�Oh�fH#YT�䙣l]0=8s"O��镨�7fM��+_E��v"O��V
נI�$$�G�U?P+(�%"O���7[�t��&�!�4qC"O>��R5tȀS6%�0]>R\2�"O��9�A�S!h8��)��1���A�'6n��3$����](��|�����'��]���*U#���f���%��'�ȁ�5� �g:�8��� |�yJ�'H���.V~�AU��5�@�
�')��,q�<T�Q�M�~����'u����ŌPX�����!��i�'�`�$Z�Tl�{��i�||2�'Pb$R7�1ޔ��k�&P�ހ��'��A���9s2<�z�e'2-��'�,���g^?j՞� �E��N�Y
�'�L��jѴ
��
r#ͅ�2�a	�'r|��
��5��`*�Kx��Y��'G�S�D
> �e2MQ�p�6�
�']
M)�B�.����(� m��Yk�'�\�����.%X�X!�(g�2���'@j��cFI�;�k`
;f�>����� j��!`]���i` �ē_Pz�{6�'Y�'�R�0@�+u ���bʓ�;&qh�'�>��D�B�Ay�Sb��(`s�'�&��*L��������dܰ�'̂��� 6spjD�K	,:\hk�'��Q�ひ;�90Ё)~��=�'���9q��6!�� 
Bq@�9��'_��rBK�.6����੖�<��л�"OFEt������h_�>�&Y+��'[�O����i\�!d����߆x��Q��	d>M����) "��ӧ(/MBlY±�:D�������9
"��) �X��9D�`�'�_�rg� �d���*}��P�1D����cգM��&$�~�ņ-D��ZЦ�^Q�aȄ=/1���7D�8H�(�)U�=���+E�Xh���6D��[��%&�H�re��~bP8ꃩ*D����ϕ�oV���-��e��K'D���2J�-!�}h��L!À)��%D����^��:�#É#RFIQ��#D����.W�`�%#��j����n/D�D0D��?<��
v%��g�%��.D�8��]�r�(���,����'!.D��BS���3k��i�HM�R*t�?D��i��ʆ>��b�/1�h��L8D��k �T0|۸��	�P�0d��6D�$۵̟��qJ�D�wg�9��L5D���f�
�sV ��/w�}��+2D���C��P:c2��$[t���'=D��#�!H	>Zr�j��`�@�ɴ(7D����L�)[�Cקfw�TPѪ��y���R�L�T�H[�	[���=�yr'� \��o�<�ܜ�$��5�yb��0<�>Ma奃 /�A����<��$	��<`�C�#����Ą%A�!�[ ��uB�JE�"�(1�
\s!�[6k�����'�PT��@ՃO<9�!��%&ڊ�X ���rQ���%)Ӝ{!��)d�p`��!�b&��A�s!�$C��Z���ύ~���:��H!)|!�DB�u^E�E��oK�=�EZi�!�D0"���-�-kL��w'Yl!���!C�0,q�Ŏ�Kw^�	���Pj!�D��*�w��f�D:��%�!�L5�8���ZCMf������!�D��n�0fd�b<JQ`�8!�D�:-Xi���6 �rd$�!򤜐NWpZ�E�:X ��C�S�-�!����h-)���la�\A��;!�D�'Q�y���(X&�����F!���%|��{U�
(@�t+��9$?!�D�:E��&�O!�a1�B^�!���7���&�
��q� b��j!�^�U�Y����~z�)�a�Q!�%a�����M0qìep��G�x�!�P�8���I䊢0�j��@�Y�!�d�8I���R��k ��h�%��.�!�/C)�U�f�Z�z�f�rw���8�!��\�`Ma�bSC���%�ތ,�!��ɦ:1�S�$J5V�+"8U�!�d�;wh�M+C�J%6�t8eK38�!��O�`��H�L�����n!�A�|�z0�Ԩ�HO��a��Se!�	�'���t]H@,��BmM�-�!�� J��F���E���)��Su�@=��"O0���^�a����&��"OFqK4CßS��	��OXH����"O��g�sh�saB�$/8��""O��i���V,F�g�(P?��9tW�\%�8D��'? P�da�kA͙�,���r
�'��QC����64��$N)�m+
��(OR�)֧A�pż2�
��/��x�"O:��U�ټHF�ڑ+׆f�H��F"O��0���<�j-;@��)I���ɥ"Oh�Sv#�0T��=Z�.�--�F�"Ob�iF(6��� �-�p�q)P�\8��p��$-�:�j�E�mT�x��`-D�pZP
�0yH�<��EV�3'�tC�$&D�\���� /�Dm�ҍR��0���!D�����/<d�Y��G]�e7$��1�5D�0��0=Gt�0/['2�$%P�4D�����I�׮fT�ᕊ�V4�B䉍\���ڷ�^(�p�yBhV/,��B�	�����#���M�I��4�B�	r<��l
���AwfȖ?ѰC��5e@��3oF. �A����+��B�I��qz&��mQ��B��R;�B�I�:9�S��][F��)�'�B�ɣG�6�0�OQ�<�����3W:�C�I1"q�xP�G�cW&8����Y<B��6s���a�ᎀt(�KW�C�.�B�I����A��ȑ(f8,�b��2HzB�	�U�h��6H�e LY�"AK�B䉑(/hիs%�'O�� Bd�� ,C�	�A;�����}����N"7��B�I5S�(*��Y�O+��2C��Z��B�	�F2�� cW0�!�fkO!��C�I-{d=i"��|p�Ա��Y�]��C�ɸ��M�5 ��{�U�N��$�B��!L�ʹ3u�<<dH���b�9�PB�1pD��X�
�VF4 4�ʝN�*B䉋n�(������9v�B��bB�I�B�M��%�+��:��=�R�(D���"ѽ��k�ɟ,b���1(D�����+p�RA��ۃ$(n�id T�0*����BpiSC͝�:�~u�G"O��f��%%������=J�h�J"Oz�-T=Q�m�u��j؎���"O��z��|��c�ED�A�f��d"O��H��>d
9��ɖ?Ӕ�[�"O�ERCF]��0�"� Y�I�"O$iQ���fB�p6!M,�� r5"O������:jh����^2C�Hqx�"Ox���䇉)�^D�C���P*1bQ"O ��ՌMZ ����1iڰ�"Op�Aa�>L���YW��BQ�A��"O@�`"/�4S;�ܙaI�4<p���"OF��� a�zBH �$Ô��"O�u� ?@Ħ	���>J��"Ov8�L�o��Q�m�*6x�C"O����E���*�l��(!`,�w"O��(�u��`1��R`#�"OF8ɷ*@�5�$�N �d��"O0+q��wA�|;��V�����"O�PJ��&B�a6gݛ|C*��7"O�0 ����9v�ӱl�JJ2"O�����1��x�d�P�^A2"O4�q�%JL������Q��A��"O� �mp�!K"���&��B�ZS"O~�Q3�ݤk�ji��d�'	���Q�"Ol4��i�R���B���%`5"OX�9�HA��|ca�DB��+�"O���#A>kSꂬ��j�"O�'�\���aW�T8Y�"O�x� M�C����ۈ^c�l�0"OB��w�Ϩ
�9�.� �`}�B"OZ�KUE\0h��h�*�N�y@�"OP���_$#) E:�o�>��`�6"O|��u	R
b���J����w��Av"OʁKŏ�\��G�R�t"�"O�pXd����e����eXPLs�"O���Z�Lƥ8cDܾg�FX1�"O~Q�Ę`z��c�5W6t��"OZ�aq�0W#&��B��
0�aC�"Ov�!i�$��1@!G^�]�<�"O�H(�dӡH��}Kad�8�tԙ�"O޽r��ɱ1O*�a2cǮ!�0�1 "O$Ip��ϋyhրʣ��:(�$d��"OzM0�X
'��E[�IYS��![r"O�BF�'Hz̘����Hӥ"O^�Zf���f���)�ۇx��͊$"O�XJ2H�vt�ǖFS��Ò�T�<a6�L�WZF���	�Q��UQ��T�<q�Ɍ	7�PP�5h�7uiP�P�AE�<�3�_,]q��� J4}�l�G�<�6�`��+�l��Sn��%e	C�<��HS*M� 0�BX�4ú�2��}�<���ͦ/ ~H�'���&_r��PKz�<���X�3o�4�F��Y0�=R��Gu�<)%aÇ'4���)6��C Ft�<��N�7� c@�)H���p�<dMH�:��)`��ť#�BU���G�<YFC�,6mB���1���aT��n�<!u���G��8����2����j�<�pk�0�&��b�V��); $i�<3E�e�.���&*2ҡ����M�<ico�<r٢R��|�~5 ԋ�F�<�0���% ���Q�ʫ0D��egAz�<�@��=[f�kR��1>�<H ��r�<y�-��:���j�kU�U�`0�2�o�<�$�/���R#T%�5#���k�<�&Ş�qk�%;g.�"mpNЂ���r�<�3��%��!�e��*3Qh#7D���5���ظ�fN�-#��ɶ�*D���v� �ċ @6t���(�(D�XQ ��Q�P1j��B%;F���%D��P�b��`8K�1E��@'$D�H@fI��,r�P闋
Hp 0g$D�����.Y��J%&�9q�H��o&D��wj/��� g�װJZ��gj#D��k�߅�������6����Ԍ&D�c&
&=����S�m3�d�f D��h!�F�u0Q�`���n�R�*�L<D� ��G�����n��q@�	��9D�H���~"`y����tQV�+�j6D��)c�>S%h�2F�"R2PݹUd*D��22��P�T�u�� p��'D��Ecڢ%��;��
��+D���e�@B@�B��-׼Qv�<D��hU�:xXQ+tmF���P��;D�D��@��NP1�b$�3��D"��&D��s�*�\��A��§K����$(%D�� ��B)۬i�vY[�Ǻ$�,5K�"O�1�D��$pZy0P�I7m��b�"O���\�ldL�Iw�%�"'"O2p�B`r09rp.�x�0��Q*O)�����~^��&�TJ��"�'�|��(&��CٱG�����'�uP�d 	B_�D;w�]56h>���T���d�$��8�1���[x^ɆȓigfC&%��.�R�G�+�Y�ȓk@�iyf�ؤ~Y�a�A�גW�]�ȓ�	��ז	�V��#LNxLه�Lr��B��0*⎙�n_�r�X���M]�H�	�7���e/S�!6d�ȓwJ�ದ��⅕�=� &n�s�<�B8Cc�8�&@��D �N r�<� N%c�PY����`f���q�<�K�#���уaŖ.�ZFe�u�<���!v�#u��"�Q�eCy�<�FJ��(���"���ˍx�<I�]�G��푓錈sQ��R��^�<y`U<}��'�v��(blT�<�gN@�m�R`��A5N�b'
k�<Q#b�$1��]B�#�X%x@�2��l�<��c��H�[�58J�"�e�i�<���2 `i(�oQ~��<�$��M�<�c� ��Z��t�2br�<�pHKKc����ΐ�P@�-��i�I�<�E�Ϳ�}�[(�`(W\�<����
�WKR��� I�.�C䉐;XP���͈�mm6hSU���5Y:B�	lmdpc͓d9bEЅ��F0B�IQ�,�x�	�h�>Q3G��|ҴB�I:����fK�T6��b���1=��B�Ɏ�$�Ss摹P���W��(:�B�	v� �s�`���ղ!A&�C�IQ"�-��f���Р�d�C�I�4 z�Qp����!�Fb]���B�	����~t��p�
#xB�I�W'��@��~|x���֖�bB�I�;ɐ�aOCP���CJ�k�,B䉦$[�����m:v)J�G6k��C�2=��J�/V�7��l��_d��C�	�B-̕�fIЕ1�ؼ��Lߚ)�C�I**t��  �v�t���\�v��C��p�"\A�$�nr#����B��!?*Ԍ�u)��6t�yg+XyBC�Ʌ+y�m��Ò�v9��q욳w"�B䉐`����-8���4nt%�B�I	^�X$�5.�C�.��d˻/a�C��vr�!���>*�`'0%�ZC�Ɏ�!X�ʋ\B�E� K@"N��B��/�\�2dE f몬��� �3�B�ɇ$�TPAr�
�uQ8ljWK ;T�,C䉪*L ө�,i����PB�wE�C�I�j���z��J��=��Z�t:@B�	5/h@ �rMA7�%s`�R%�BB�	�x����E��}���\��B�I
rl����&Rz�V��[�,�:C�,,���g��	��ʅA��tC�Ɍ�p�CuoO'n��T�d-#L�lC䉉�XH
�)2~}��S�Ȅ'AdC��	W�\�Bs��]����'ƐN�B�I�j���xB�+I|�ZG�ė#ռC�I	�
�q2`ɒD<����H1�C�)� ��ʔ!�J*��x�LA�$^rq��"OR�� �J�)E�8qr!�.@��"Op�U#�� ���Q�N�':��"O���1�ΜZ���5���
"O�z�`��Af8tx��E5���"O�d+�fU�Y�:�9e�ڗ=�.���"O��RE�\��{B�1i�m�q"O���g'WUi��C� �'q�|��C"O���痂*x��/U-c�t�0"O*������j3 �Z�φ8��Y��"O��q�˲%R|8!N�5�^qȶ"OR���e	�-cvt��━m��2"O�-��]=�NܙH�Ew\��C"O�YU-6Z�r�(�An����"Oΐ��خV�}+ aG#jYr���"O@<�Ŋ�'�}J��] Q��!"O���1+�LUZ�k !(6���1"Op�˴��9gn�y�*[Jǈ]��"O�8+�[&c?�����(ђ�"OR��c�B�>�����ϐ�n4XIX"O��S����Vt��:'�1��k"O�����"�~my �a����"OV|c¬�4r�A�Hƃ�
�y�"O�Hk2nJ�Nd��7�N=X��p�%"O<B Ǳ�fX�q%�F��0U"O������^����B�^�d�;"OZ]3��@�1q�eC�%���g"OE�q��B�KE�sڞ}��D��yb*M)|�����id� I��'�yrɔ��Xp�lW�\�����"�y���G 	[�$�=[vB�z���y�BU	3�E�!��'ao�ǃ��yB'̄
C��+�� ^J��Y�2�y�Nm�F@�K�*HB�i�0�ybMGXl\r�C�йĒ��y��I�b!��lD9�pP�$Ő��y2̈́�c�,����Q�{�#QaN=�y�BC�a�l=��D�z�^�b�f
��y�W��%�B��|X،�C����yi��C�6��l�D���ۓ��yB�ĺM�=2a�D�1����3�Y�y� �,7������)0ҝ�M+�y�O1 ��P�D�8���*j��ȓ0/��0��"'��Qq�mĿ(�ra��qL͈fn ���?H�u�W�>D� '-��4n�yn�TQ8z�+;D�|J7��r�P�Z.�G��uu�-D���Ӊ{�:I�cc��?�����,D��#aO�8s��C*��kyT�Ц-D��Xqh�;�`�Â/[&��I��o)D��+r�̬,u�Ъ&a =q�!D��'( �A�P ��9���:D��ە�ϙr�(�s��om�����8D�@�� a�r����M��,��;D���H��!:X��D�0Wv��c�3D�,�P-" �~ĉ%c���0ja�$D� YS��M������w�Y��I&D�� �@ e#��9CM�T+�1�ю%D�L�c%</.�B��3C�zQ�se#D���2Ƙ�n��a��Q��F�0G!D�$��Y�"�FJ�n��kQ�$�?D�D���D(�H�u�\'#� ����0D�����S} )'[	��B��3D����"��-�ֆ���-���1D�� �����$uG8l�!̓�����"O��Ԁ�y�n�22�x���a"O���"�وW��r2�Z�w�QB"O�z�䆱Z����.dv`ŀ�"Oh`���8ZY����ݘe}�k�"O�	�T#��m4��%�RH��G"Oځ���ݬB��XٲO��26�=Zt"O��J���e	 5i�H�I�9�1"O�ԁ��ٔG�*�;!�C9]�,�0"OD�w��F�b%*N>,8��"O&�e��(��P�
���"O:p[���d�<0�'J����� �"Ov��	��H�PV�]0\�H��""O���U��l�DI܁=��A"O
�2�ͱ3��L��jO.�$$��"OZ4XQǆ#0�DY�)��ěE"O�p+�/�L���z����p�h�"Ob#��U�f:r�0�hA=<z�B"O�HR�ܖDW$�Q[�1�,UJT"O��3!B�,&X噇�?1�-�%"O��86��~��ү'�,- �"O� 8�IB=�ve	�N;�$���"O���u���:6��1�9�t�C"Ox��f�W�!n�8���W����"O�eT��22�;6�3b���c�"O���Ǘ08 �QFN�p�C�"O�����_+0nM0p�H%I�*�3�"Op�@7�ѵl?(t�t ��ndH�"OĤQ�
ބ���a��3UX5�!"O,`��G{@������<3����"OD�����@�М逢̣{v�P��"O�<H��G�j�x�fצOk�m�5"O�h�W�Đi�(e�L�2i̜�F"O�lz��՛z�<�zD��55U�H�"O��
T�˳CC���b�,O�ZI�G"O�x���	�Tސ�:bc�"�U+�"O�H!�昜a�X��ȑW�~�"�"O��k��/1""p F��6���""Oĕ��m5} h�i\�[���#"O��,�>_=t���G6isL���"Of�x�c�!���R�,E16�d�`"O�l���jP�
G�S^�\˅"O���H�!z����
62_����"O��El��x%�r�� xIp�@"OJ(
���f�
<H�'�����@"OT��$�?b����`�A JE��"O�|��MK�ZQ�d�6 �����v"ODh3��i��l{W��}st1�d"O����.`�	����ti�Y�"O|�!DY%_����ML,�r@��"O�1E+�0xo����o��R�@�"O-���=2���[.K1�Đ"O�����
HX���$r��"�"OVPa`	�:26��j��P}Dt�"O��#8=Pc(�$g���"O^1D�J6j<��%9�Puib"O��h�D�B6���N.|�,s�"O\t�b��X=J���T
dԼ�"Op�y�K�?�e��Y)/vt(W"O�;�윽Sh��iE8H/��"Ol��JB�TY �4h� \'Ҩ2$"OЭ��#
�����!u#h"Ox4���O�mI��Q�i<4ӄ"O�̚#G{"f�$#�.���"O� �(*$f��%_��X��S�zMƉ:Q"ON[A� e�l��G�/.�I�"O���0��3;����$F�W� ұ"O�A��j �/������*��t"O�=�?���pǥë?���"O��S���3��P�f�1Z���
e"O���Մ�p���a��
�6��e"O�U�A@��k��ar�m���P�"OԝC�lK �*a� N�/�}�q"Of���R�v�a�O����w"O�0��^D/��;sJ�5%��@�"O�ɀ�o�i
��9�+H�>�P�"O����§A�Α��,�#�B�"O`Qr3d��@� �E�Z�.���I�"O&U"��Ͱ��{�(ՕLݢ��F"O\�ӂ��.C.��k��S$cİ)�"O�}pAA7 ]�Yxdř����q�"Om��,�B��S�&W57����"O��H���p@Z5$ת�͒�"Od�����Yya�"��&�v���"O��iw(�(��C';k��Rr"O�]��7 TVͺ�4ZL=��"O�lc�.��-$L�PS �*KRTaAs"OL�ጆ	2�`���!W5�lC"O� �V Y�YMR][�MW-G)v���"O�ap��C9l�P�0D�� $�(7"O�e�D%iI�����5�q"Ỏ��Xb�V�bǤ_�=� �"O��s���*-a�щM|��$"Oz�cgӚ|%��x ���y��02p"O i�Eg�����P����x��]�a"O\�!QO	�h@�Pe�ܕ_�LpK6"O�m�/�>R�r&����$�a"Ot���"n
l C"�J?V��â"O����D�)j����	UXlm��"O�QʓK[�r݂I �Bۅ8N(�� "O���.st�쓰!O Z�"O�hQ��'vO���!G�йK�"O���Ï�[A���/6��2P"O�x��łY%h��E-W�Y"OF���Hb$�����}h�Akd"Of�{�"��DJV��s��"K���v"O�-;�Cў4���	]�jЂ�"O�h`���2H�q�J�a���""O�S����*;��aC`�	�ޑ�"On�ʰ����Hi�a
�w��	w"O�]�E�Uqs2�I�@E'eK�K0"O|���Mܓz�~!d�ԷH>��S"O��i�S�'q��B�͛��}9'"O,d���]�~5^�8Q� q��"O@��%K� {y�q�!���<��T"O8���'N �� Ar��Q��"ON�0I��Q��p�j��)�*�k�"O��25��m�LA�ri�A�0��"O�(��LZ�H+I���}D�R"O��@��� @�>|��%��Onܓt"Ox4��Bejik��H���1"O����ѯx���Aѹ�e�C"O��i�U��J}�w W�h�d��"O����&�1H�蔎Y�����"O�8����.-� !łS� �H�v"O�*�a�`:h(� E>lH-z"O��1�Ι90���� �,g`�1��"O0Q0v�V���e*���?� M�"O� p +�H3W�y[@ �B��M0�"Orh�$�(Dޙ
�����Ґ�"O�A f+ԭ�&d��F�A�,@y�"O�|"��( �끆�`��xe"O,q֯X%L.�0T���t��ű!"O���fX�r���b������S"Oਛ�ہ5�bu7�������"O���$ş!|Νc�\w;@i2"OXa��ҲH<�pB4 �"O���.�_]d���&��ctU��"O�u`A��1~tRV��V��X�'"O,�QJX(z�\�٥�R� �� #�"O�䑄Œ�0ڎݚ7$��d���"O�!�1m(K�|�Y�,Iz:jF"O�D*�+��Wն�� ,�^m��+�"OT��v�,'� x@#j��SC&phE"Oi9Vm���xr�_��l�"O*���mY��� �4*�5�Cd"O��J6��3)��Q��	?ք�3"On9W��k��x�ߕ}���""O>I��[�K��EkCX�[�h�`e"O�̢blf̙�ѥ=ߒ �"O��a"�)p���@ŁF0M�!"O] ��_8.f����E,{�(S�"O|cA]�F��)*VR�]�~�t"O��"�+K�"
���� D�F<H�F"Oza���R�t;WJ]�P�4"O����턚mz�-%�[�C���9�"O �E]4BƄ��A��I�l�+ "O(���-����ge��F����"O�4�"�E$Td}Z%���)Ps"OR@R����I6d<�4#�,2y�4[�"O�RTc5�da�!.` ԁ�"O��{Uܮ<X�zA/D�x;�"O
���AU�"
��M��ey�"O�MIV��:&Vը5�B��U[V"O���wʗ biLD��&^;u�`Hx"O*ͺ5�ң�X�N�eʡf"O���$�H�|ܓq�@�4>���"O���ǀ�8)��5�roԴ>Z&�J�"O�`j�H
�$9((a�n�LC�;�"O�0�3)�ڬ�͝*^,�e��"O$ё[9���v ��i0D`g�K�<paV��L�0��,B&�}@��z�<���s�E�a�J+z��T�J]`�<is����	r��eo�Z�<��Ev�(��C�0��1���_�<���˙x�t�) ��o���p(VB�<���[=�t-1���>g N4wF�A�<a��M8'�P%��OJ4�e�]�<�A�\�l;�H��e�.3�w�<� �Г��̀�
��xr2Mx�<�G*Kt��`M��k�$XʓNWr�<у�K����@��0�|��2��y�<�r�=h�@k�)X�6qJ�m�{�<Q׈� 3φ�۱�_&�؀�V�U{�<y����X�֎�$]n@q�'�A�<apW�}�pw�M�G?bU��K�z�<��(P��a���.�1�L@p�<��
%j�rF�5*�P\�� �v�<���M
�1a�#�/	��i����t�<YW�_�V�|����{��qHp�<���,K��Ң�ĕ��q�%��A�<��!`8L��	�͆m)c!E�y
� $pzQ�%*�x�W��!y}JD	�"O����A`�^����z{N|�F"OI��ȑr��i��T�l��%"O��B���/Hb��G��$eMb�"T"O�m:��̰U8 ����oE� h�"O��g�&H���S���Jc��c�"O���E�S�r�W�Mz}|$ȁ"O�!qĊܟ8�hIS ꓱ��3�"O �:1J�$>��6H �*q#D"O��S��F�.<X�G�$j?Zܣ`"O4hy��9gL�
��Q�MC���"O�h��)ޑH���I����~\{�"O��M�(�@�x�#�c4!�q"OΉŹLN�����ۃ$a`��"O��Bj�ZK����m�8a@�ʀ"O� ��C%�����GL�PE�9��"O�T�"J�-z2������+]�f��g"Oni��J�'x��Y����r���"O܁y#3QV�-����ɓ�"O��䟱���[��Q,L|,Z�"Ob��fЧ ����4�[����w"O1h��X@�B��`nPm�-*b"OpX r�WXƶ�@�oYT�8�0�"Oޙʇg�L��Baw�$�@�"O������Z��y b@̀K����g"O����]��!��lԽRS"O0���k��!^
Ǎ�*$;���"O��Ѝ���P%XsG��9�iv"Ox�j��1�dx��戕l�b-��"O���(������J���<z�"ORyْ�F��%MF5e��8bU"O]�q��y�����0T�@�Q"O� ���Ѧ�-(sr�N��l�"O����	bf�!1wI��88�U��"O�=X��X��ց�f��T!Z�{�"O���� ��i�H�?1
\��"O>88S�Y�P�ʱ�IU�GI�5"O���R��& ��+&`e"O(� A�-Z�VĞ!������a�<A�dO��2�Z�SO� !#'�^�<�d�7q�\�p�\�;L+��E[�<)1`�d&���O4JOtۥ�B�<��US��P#�OݧY�Z�����f�<���a^���#�
�4ʒH�<Y3�+F7<���B�B�b@{�E�\�<IѨ>S0b�ܿ*Q��
HY�<�b����ha�*��(�%��W�<I��M2$7��9#�Ԛ$XP ��CV�<Y�]�_����こ���3i}�<��̈́�"�8�{p%�<�@<���v�<��]6z�;3��h�j=Y�N]p�<yp���o���{C�I�辉�(�k�<	҉ʻ�<q��Ë�c��!R�`�<A�F��C�c�-��,&�Ը�ȓ\�"���hg���skZh�8���K�ִ`��
jUZ�`�m�� �ȓ+<|!K��_�<n�<����+2�ȓz�Pۇ♏@�hi�s�˟<���ȓZ�b���T (�`���3"H��A N5 ���,\1�C' a�݆ȓ(D�)(0I@
)JU��D~L�ȓ%#Ȕ($�X�QqT���NZ9X��Zjȹk�R�J+����� J��ȓ(�䙀�$E�\��5S7�]�v���S�? ԁG��T�	���5��"O��%��&�X�X듅-�&!"O�	&��SG*����̦ ���"O�d�$Z'��Ӧ�9'w�-X�"O�Xc"a�PjY;�UT! r"O�YPTLޫR���$\F��9r"O�HrJ�!H���BV0A�U81"O�t⤤�QVl�����.��#"O$(���Q�>`4��gIE8v�I�"O��aAɻ9`�2gm���\��"O��2�=�ZI����${�"O�d�G)�X��"+�t��l	�"O2�����	5s6TK���"BM¼C�"Oʘ��*J�4\ `A�e��X!q5"Otx��Y2u'ZxkPC�5n|�F"O"})!gS D=�4��� �Z_4)�"O,�-��0Nڲ�P�4b��"OVѲV�Ω0l��i�$§|ڤ�"OH�q'4�,�+�#�F��e��"O����� \$�$Ǚ4HQ�B"O�ѳԄ�?����FV�=40�r�"O���5b�b�"}p�"~�u2�"O�i�"��v�D��"\0,d�}cV"O`�AcE\47�p4{����<KH2 "O�Q��1N����S��
M9�l*�"O��8#(�Ha��H��5i6\�ZS"O� 0�M�?����ڴ
 Z�HU"O�(e��'Sڵ�ta��sq&mSR"O(��ń� �q��eʐ2\�9��"O��3��.`���"���W>Yd"O��3���=K\X�Q�D?P�=��"OP�8���X���x"._%x����"Op��U�9HDJ�m�	�~�+�"O�XY�d8��D����T�4d��"O�e�`&[?2E�fH�B�ܨ�"OHXD��4?f�C�����8�*O�\��J�v��⥢�	��P�'��p�"M��z�6@��F�� �'W�����J���x#U�7��y�'G�0�%�)~�1���R�s�d��
�'�������}:]��H�v�p�'X��`���b"z��Vg��;�9	�'�N�`�nP���a��譠	�'�ZqR!NY��%iƊFV��M��'a�i05̂)#�=���J!{�Q�
�'���3�˓>���I ���40
�'��4�D��@���"�˩��e�
�'t	Q2%�{8���`�R��	�'@���C��7P���1�^.Q2&�H	�'�jդ�C3@Y�J�;��}��'�Z�A���!����� @�C(i�'���rr��?�+��W�	��n,D�J�G�:-��,*�G2"H�WN7D�t8��P6a�
-���Bo�A�<���P�<����@ؿm� �F��@�<�F�W�T���S�G�'x�����FPw�<��Z7�ti�d��w�2�	Uo�o�<��t��!��R&v|T�	u�e�<)�d���倁�!���Y�z�<��!�/&����S�j��3�bx�<Y1g	�p*�g�� E�RɃ���k�<I$j�:��a�K��蚳�o�<��Κ�t�C���L���'�n�<91�@4FS�-���P���[&��s�<� ��r�W�^f�P�� jD�<S'"O�!���;��u� �,��b�"OL+�g�2B��Kro��<����"O�{��
6��X"��V�zvt�"OLh��J��S�<?b�T�%"O���E���>$j䬓%0GTQ�E"O5���L�~��U�2��*Z9��ۧ"O��I�!F�RCl�ʐ����t�F"O���Ń��r��GL��FY�Er"O�1l@OH����g
T��"O0���$`$s��O|@d�"OFy��WJ�����KޤS`��+'"O��IP'y�b��ꕚ:$���"O*��>|�� �G��@"O�u� ��DuA('
�|0"O���m��dRB�h�O�� ��@��"O��e�\�� ��W�O�n�&�`�"O��Q�?��q2�C�.�x�"O��Ņ֣	+��Q���$����"O�%:�o���9`�E�N�4ܺE"O�����S=Q��tp �C��"O�M�oQ6A^�ip��4|�j��"O��)$eL+!��7!�(f��A���+D��d`@4h	c")��V��,,D��+6�E'Q�����?zQ"�C')+D�P�$�F!*0��I�E6���W�=D�pP����L43�*�1��L9�%<D���c�va���TL�\~��q4�5D�8�t�ݠ0��S@-��Ћu� D��*��T�nY(�24NB�ZE��+D�d{�Ϙ'<��8�!@f>D}Pd#=D���c�\�Q{4{�Է|�90@
7D��ce�S<\�aLE{]�,Y�C4D�d�լ�8r�¨!�_2R;��vJ5D��k�η<���2�Z�@��lr*OVq#�V'a�l����T��a��"Of ��ɒf-����%R��A�F"O*�T٤h���G�'3��
"O"pj$�!���kZ�i����"O�1g���"E���)/��"O�t� h�0�0h��Vw(H��"O��� ـ2�y�M�7"�9�"O�e{F��|!�3�Qll��"O���Q�C��c��ͫ�"OxQ6. �hA�(��N�U���"OP:)]%���-��^��V"O&-��A�ozzP��B�ό���"O��s���e1���)���ڀ"O�)PP�T�g�dE �����D�ȓ"O6��T	ܓ}�Q�a�$a>�@�"O�l��+\]���ku�%)b"O�M vZ�h2���U�VlI�"OV�Y��Y�sϬPxӅ)uA��х"OҌ�u�/T��1Vg�m6��H"O��R�W�4��F��a���&"O��V�����\±K�.�H�G"O���V(�[�<�d
˕��PA"O捰���7o���gL�-��h�"ON�bq��y�4,3#l�:#�2؛�"Ot���J��g����HȪ��N�O��-3vIF/a��]�DCͳb?$9��'luHE2u>X@S'+�b���
�'BPH�gW#@�����=a���s	�'3�Y�ӆZ�&<X�����\�*	;	��� � ��)��3��e8ff�6;�6"O����� ��Q�E3�a�"O�Ub�! � ��Qd� yV�8�"O�9J�	�h>�#�ׁo�h�q�"O��1jЇX���� 	Gt�Zc"O�ِ#�>vP@�*��K+Q�D�J3"O�UB��"�v�A�MYP�Ze1U"OU8�
�&R8y���I� �Uh"OL�bS�Z
��XI�KԖz�<\A�"O�QFGѿ��!�H#� u:Q"O�qS&��<n��cGH� ޤ�U"O�u��[)�vA�t]�uqR=
�"OT�U�S�v��IR<g襂"O��QE��.|�P�]..p9�"O�����B��B�� �7aLX��"O��z���8h��s��<~Ǌ�3%"Of�R����"ę�kG�`�i�"Orx�(�v�d��@X8z�Hd��"O�|Kt���m��y��"Z�C"O2�ySMʂ�V�[�lZ�
�8"O(�1p"L r�m�3���"O ��ٰh��ɭYP�l�0"O�A�k��[a&��tIM2QH�q(1"O"L���(Bl�H�Ȑ�>jl��"O��c*͸\9f|b��_��,w"O��#cY�;u(P�eɂ�
x��"O�CjC
㪖�z����R<�y�BƦE��D3��q�����L�y����f��b��d�d0 ��y��Nʄ�:�P /����g@^��y¯�"κq���Ʀ]8������y�$Y'+��i��H��Y�pAw��0�yJ?u�p�qR���e;6��w�@��y��"tAl	Q c��]<,Q�j�4�y�kچ)�B1spݯU��ٚa���yB�H��"��"�Ч�ʭ�yrӅ&wR��6,I�xk%���ɧ�yrDM�C����a�H_�,=�᠗��y�ݩ �f����O�m� �W?�y	�k�*�GM�?�Lh
 㔉�y��� K�q2f&T1'��!)$�yB�Еpk�M�A.�#"GX<�0˅�yRH��|S~]�w��|��+�y�(�?B���H�[N>�}[�Kң�y�L3��@�"ʤBc���'@��y�d�=$Ȱ#TؖA��E(��.�y"�����ٹ8�ƫ%�!�d��	�^�aI6U�B%�,�#3�!򤃪&5�ԸaF�!S@@8u&΁+
!���4yj�"��><L��<o�!�$�X��=aW�2�n����\�a�!�WO����b��A��Ab�ႌA�!�ٴeE�Ͳd�B(�,��g��w!򄆪d�8�`A��:l��CP���B�!��'5�� �D��?dLц��:�!�$	=�@���?E�`h�A�4z�!��E7=�rQX�Q$|�%���7�!���;��P��4i%�X@� Ć&�!�D�?bi�12�
�L#l�ӧo�8j!���5+ ���$~d��,�4!�D��渠�(�(t�}��,�#!�d���XTx�k�z�v$!�쐔 !�����1%�&_��L�K
�J�!�$�)�0��B�*%��D�A�/�!�� 0ī��8x�&���a��C����"O��3���6n�M�e!�~\f�"OX�r�hT&C�Y�e&��)��x�"O��v'��h�땩1����"O��a�I�g�r\k#iQ��h��"O|��U�ը�tU�è��^}�Y�S"O�D*U&�,z����d���to�T��"O�z�i�4N�܁c5K��Q`q�"O�}%,R/{~�I�RI=D\�Tq�"O:��(�#aR�gǈ����Y"Obu�D�X&D�(d�	�Zl��c"Ot8�O�70��%3���A���q�"O>�Iv�'/���Έ2C�P	�"O�ڂ��9^�ԡ-��\�t� "Od�� �Z{|��F�^�s���c"O��t�N,�����9��"O�t�e ��w���#��6˨��0"O�X�tM�4)|�$I���5S��U� "O��0�F@��e'Q\�:�*�"OX��b�*d����e�n�%��"O�x[�HN��i�4��:N��;�"O4rC(�/=9�e��j��5p�"O����`�챰A���h;�"O��$��{)��92�Ax�0�t"O��[�/h�f�6�	&^İ���"O��i�EԶu�%+��x���@W"O�0��տz�� `Ez�&�3"O�]K�nʝD0�M��$N3q�č�"OE�� b*LZ�����]+"OݲG-� M$1z��Z$HB���"O���֠�&i���
�Њwa��K�"Oz@x��5g��PTf�3jJ �g"O*�sQ��yfj1�E�	����S"O�L���E�88͂���K��MzW"O6���	p��
uA��fu��ӣ"O��Qsf "!�h� T�9�z<��"O��#��:����H+L��`H"O��ƁT�7�ܰb�G�'�n
�"O�(��hV<ծ2
�>K�y#�"O��"E	 n�4#s������"O��Q��X�@)��K#9Gn�� "O�M� LKr8���͝sB�i��"O��0�'�G2��""G����e"On���E>����0 ��#�"O�y��ɜ�:����G��[R�P"O��pKW����B�] u����"O���2JZ��|���ʹ0����"O8�L�\�����W+O����"OJ���gL(4N�r&O�7X����"O��c��9 (� ��=@$�T"O��� ʝ�p2����Va#��X�"O��Z ��X,�,�t�H1P$���"O<��-ѕi�H��#�U�D��*O�,`�K�'fŶŘ[
~��%��'�|{�$��|v��ҔI�'r1�Ј�'6.c���-��"���k�X��' v����ڙ~h =�r*EW�p�
�'�Vl�@�sx���n �d��Hx
�'q�1�ɏ�2-\��W��]�0|��'���I��b����OV�[����'B�� ����5FС�q��4[�M��'!�Ӄ��-�4���n�X��)�'���vÅ�U���ֳ(8��	�' P館�1?�<�W��5tQ��� ��)Q�ڙ"�vDč�'3����"O4��f@ +'��`���ح{,����"On�7
�pҵ �G�~#��I�"ON@#����XJ��ԇ�m��"O(��	��>蠁
�)�-{t��0"O�i��V�T8$����S�:��V"O�*% 1'?�%���j갈"O�p�(�)l��}
��r���y"O,�P� רy}hӐ*���Г"OL�����|��t� Ç�lS�}��"ORX����"p�"��A�y<�Hq"O`A�f`�����ao3�<��"O����!���#˚��D"Oh��iØ?W(Ce�J"`P�"O,`zcnָ59"���W�o�x�"O��J�!:�ȳM�g���!"O��!�b2�:6->k�zs"O(I��ϑ5YC"��j82�j�"O���N�VC���g�^
F�ܸ�"OlM2�O�R�B�0+M�p�E��"O��R�C>Ajҩ�	G����'"O|���#�� �H��;��#"O�(�y�H��!u�(���"O��H��CX����R�Hz����"O���I�4b����ϯ2r��"O��@�K�,��uu+H<gc�}��"O����ژ.�r��@��_�<��%"Ob�y�[�_�\�JR:��XP�"OPq����5p�H$��Ѹea�͠�"OPHʲ+�m�J���蒞L|�u��"O�X��勏h��x�Hd�D��"Oz�(�@Zzԡ���0N�D��"O�A��+эy:V�QF�O�UD��A"O��|
��A�i�<�(�!"O�ٛR�X���0���4rt"O
���oݶ3dJ$��S���W"O�����){Ƣ�^��\r#"Om�4c��@�ȕ�����D��)R"O愂���=*Y�*y#�=��"O|����ut��p��`��ջ�"Ox`��-l�~�@�����"O0��a-VI�)�A��WҐ*�"OPc��Ϡk��H -�G$V���"O���/N�|��-��.�K ��U"O�����	�0�\ix�k��x�A"O\��"C�L�޸Kw+� O ]�6"OΕKW��Ym��`�Ӹ')8y��"O�P�U�� D����`L�/'j�Pf"OP����#	�RI6�Hs,a�"O�mXÅJ*e<��c��q�5"O� 'ŗT�����ْJ`с�"O,U�R�ʔ(X�؆�H�ISt���"O�qCN����B��"^Bܘ"O^���G�"�l� VL�&ly&"OL�薀��<�X�����Y
�t�f"O�d��a�:��ƋS�$�6�g"O�+�*��C۲�ī��e��٢A"Oأ�@�3m��0k!o���
�"O�	��K���q��	U��v"O�U�5d�(*�����S�8p��E"OЀ:F�r�r�)��M7g���"O��B��L�i�f�c��cj�"O2H�م#��TH��;8l`���"O�|�خU���lL�CJ\h�"O� �QEb@���Qa�%9�p{�"O�	��.��(ɡ�`�3b���"Ox�cЅE�"D�0��/��yI
���"O�eȱ��9]�|-���A4=ΤkQ"O�4���Z>���ð�Ŀ4@��"O���7dْ7�z\h4,�-*�8��"O�P� j�0LK$���$6��s1"O������\�@Ͱ���']���U"Ob�!Ј�2r�Z�C�a�_�	BV"O $��O� V�
���?#j��a"O@�s�'�+bR���ɜ	|�rv"O���jP� Ρ��+�6 �0�*OT�ƍ1S*I����euP�9�'(Hfg"���X�F()ؔ��'��`RE��31��4��E��@�'���@C��:l��EP�`Y������'�\��&�2�vd��E-Ab�1�'�(��-%�HѢA:��R
�'Y=��M.R�xєI�	1^Q�	�'un�#ǜ�r!��i�)J'6 
�'{�	�w-��6j�i��;�����'X�c�l5"GIKW�T�%D���
�'����`�Y�XHZwi��",��'�Uʣ�)�
�`fጀC�ԅ��'�&|�Յ·`�M��LB$Qyd+�'�4�I�E^/1�P��	rl�@�'�H��r��[l<���oɤ8E�݈�'?n�	6C�=&�PS��R7����'}�P)uLQ�=��\�)s�@��
�'Lt�Y���B�?;VJx��E�y�-��@Xk�!å/x̡�,���y�G�-� �. \�F�SU�Ę�yBE>x�I��� CK�ɘ$���y��_�1��r�̙5�\�zDC��yړ(��]+:|U,���"%�<D�D�jU��$�#Vʈ��	y�9D���&�)X�J�+wAQ�f���7D�@wh�6<�b����Xb: ��4D��[�lXl��u{�'`�X�?D���jXu4�`b�K7{O~��1D� �H�=��Q�e*�#'���Ҫ/�	{�����>���*}��ʖ'����HKEPc}B�'e�h�v$�Z�&��5�D$ZT�͘�'�L���/�4@!S���'ԆQ���9�T��GƀtX���)OZ?����S�j���J4n�9 )|Ujd��\��>)���F$� �$�	� ��šB	[!�d�h�^鋰�9qj��f��tT��o�^��~2+�u��̋��I,}���A4�J��y��']��\�_Y؜��JA�IQZ�i��ݜ}!��S!&ICv�1!�nu��'T'!��֒v��G.\�{���;�'G!�dX<D�)C�Ɯ�z�i[rF�!򤘦���q�!Ԉ@c:�y����&�O(!�b��B��s�� )瑱�u�x2�'���7V`Ą:r�:?�&��. C�!��b��a@O�M�0�6�Ha��'̛&��'�Ӻ(�Ph�l�d���H�D�+hB䉠(<��U�@T(�ȋ��ám�8B�I�h�5#��� 9hy�@E�K���̋^l�Š��[S��8��(�?xU�� Uc?D�h�!�B=dh�"�#ٶM���!D)O."=�t��&;�̕��A�%�ٚ�
IҦ9�4�'��#���
\l��nQ 
�X��� \��N?j����'���t�����'`�'v�Pe	�Yv��y�ɀ�AɌE`g%$����`�9����s��/-�Ь[��5\Ob�p�Gi�����8@�ٓ�*O،y� F���m	@� �nuܠ{"O�Ѥ�׃.�E�q��%b~��*O&�����H�|a�t���Uu�� L��'�E�T⟻�4����]�Td	��0<���D.JI(���N	f:�dF�'@�!�$H�Ng���Q��Z4�Å�>!�d_k��xtʝ.I$1h祘3�!�D̄l���2�B�����ecM$u��Ğ)*A����6ғ\���� *��˙�c�9{�'��	�h� �C'ԌQ)]�<�hC�	#`�N`��k��� 2dV�vOT#<����?�"�%#\�,D�Rˆ9�:1#�`�PB�ɳ��Q8��U=�L(�w� Px����7�ɍn���+1j�	�`T;$Β4C��B��{#j��u%P�2ٌ�A�U.nYb��D{J|:��]W�r�A�N
r|����x���/q�2�,��@��#D�;���Gy�-%O��QGWXM@d
�"��K��|��"O��P���0�ZMZU�U���d�'�!�$M��؁p�BS�zr0<�@���Xeў<%��}ƙ<=֔����S3``�x�`KW�<��LҥQK�\�B�Ա�dI�PCF}x��Ex��ǓH@(Ԉ���\z8�ic��0>IJ>QeD�a_*�;���d.ec�$H�'i�	t�'
t%�7�FM˺L�g!d-J�q
�'�~��` 
�<`�\!��f�PH��'7xEY�� �'o��5:Ҥ�'��M%$����P`fJT3*�j�0�'����tw���ŋ�(,�4$�'�ʌ��X~��� %"�*9�	�'�� {#"���!bA��.XA��'�FlbhU'i��h��d�w�2�	�'�`�r ��63
�������gX��'�ƥ�2O��)���9ii���'���q�b�' ���R����ea�;�'�������)|:�����WV�P�'^I����>V��I��I������'D9�!�9]B�Ce,5m<�
�'�\��R������!X��듒�I�D x�"�5~�a� � �&��C�	l������- ��}y�@A*�C�3-��ّ�er|35�УpkZC�ɝirZ¡���@� �j�ʓ.7*�<	H>ю}RC�r@���J�,x7^�����yB�%{I��a",��r��yQ����yb%N�!��\�A�gn!����y��>�~�a� Ã^� ��7cA�ۘ'�ўb>�)�D$`����Y�2�����
5D�x�׌�,Wx,�Ql�4KsA�1���<�aB�\�̠�e���?$��D+�[�'Q?=�Ն�88��"Ɣ��±������x�HZ?�fA#��ƶO�f��c蓽�ē�(O��?�je�C|���YpiQ�0	�Q�!+4������%�P)0�ɻ�(�F�<9���z�a�*�t8�`����A�<aǈ�=/ZZnm���jbi�G}��)�'1�88{�d�4v��ـ��2!�lT�'��#=E���D=|O��;����W&W�Y_HC�I�^4�!�h��zR2t�Zg�㞀��V3n8�R�\��5���2��B��[�? � Âl��%�ʨi��'|n��V"O��Ģ��Hq4���k^�tЛQ"OH�w'��Vh��c� ���Yv�i�ў"~n#w<������@����W�.��F{J~���S:@�X19�FY�Ȏ��#�[�h��9�O�ت���5/�����;&C���V�')����Qe����e���	U�RU��	���=9�Sw|��Ä+��*I�I0U��Y�<ŀ�;/�1�� ٟjN&Qh�	R�<YlP�2"8���[0D�P�T�ʦ��!�:\��_6.<�:aF�	�ч�I�e��i!Xj�CM�UZz��� �t�"��Z��a�
6@.%��Z�'F�)7M,SL�j�i\/v��h�'�Ӳ*�qF-I0�Ú%�!H���hO?i�D��2,���0�
���V��E!�N�<YH<p�&ha6b��Bv�u�bM�<��c׳m�>�
&"?*�Q�F�[8�,P@���2�����*�)PfI`!m"D�����?s��if��%�;b�4?A
��*��5��E����B��9D�^���6�F�BP��/��A:�.� $$���Ȯ��U��%��UK�C�3O�T��.��4��E|���w�X.w�h@�ȓj0��J槜��p�Ҥ��"l6�$���ɑE�d2��N�=��
!�ͼk�|C�ɗ2��C���$9��YEL�j#>	��)r���psD�	a��B*�4^ �}B���R69v4�1ō	�B���`�=D�dYa	wJh 7�ɒV��� H:,OZ�<!��ըY�j�	"V|�H�!c�X�<)�bE���ċD��}��(�&�]��p=�D�(l���I '�6�C6!�t�<�FD�$��uY��@�d���rfϐq��hO�Ʋt�c�	��q�E� ��i��i��	�M&(�j�j�RM�'��G{��T(��(~(�'^��zfD(�yZZ���ph�gA�-��`S0o�X�ȓ&K����tZ諐,ݪ$�����?�W��{�[ekK�1�����/�m�<Ԁ�(O8��'m�'�X9����r�<�%��b&J��s�Ѥ$�;Uŗs�<��������z��<q�؝zT��n�<y���Y����Q�@U�p�hIC�<A��J�ul����@�K$E S�R}�<��w�b]@���&�����w�<Q!gΎU�TК�!U-��E#���s�<	��7Tt�#�FNG����r�<كB�#Prf B����r���$(�p�<D�6��r4
ֲ\Ŋ5b�i�<1�Y�e6��2&�Z�kd 3�,_�<4,?zm�$zv���jx�B��_p�<I��	#��	�qLɄG;��m�<�1&��:W����戄J��B��L^�<�1o�:t�d�W*V�i[ƀ2�u�<��N%\B�̫��߫�@9
䍕p�<9G�M.{)'m40�)��"z�B�ɭ_�v�eBֹ@�D��W"yC�I.#@�UP��"����焖�/�B䉊jJR4JS�|]~�q�1.�B�	��8��Έ�Dm���P�@0�B�9��+!D���.щb	��C�I�O�ޝkP�ܜN�V�ٞ*��C䉻xe�rWf�GG��Zs��d"rC�)� �8�lY;V�FM���͵N��x"�"O,����.4ОL;P�E�7x�݈"O�(�@d�3�N�2F�K\�-�a"OD��!S���p�Pφi�d`2D�h��(p*� ��`�|���n.D��6\�y���1�+�E�x�(6�-D�J��@����a��;<|�P�Cn6D��P�*M��(�!� �@\Ԑ&3D�X8�� �W�R����J�K�l�rk;D��f��&�x5a��9
�@��:D��I���.�<�y�&KY+$)q��6D��Z�<:��ɳ��d4��:VL3D�Pãm�)��P2Q^*:�D�ֶ;�h����̦���
P�1LO\�q��$^�\�c�N+o�t@c"O����N]�o��q��zh�0�a"Of�!'�%&�H�Tk�W�,�"Ot9���&��)��K�@K�)�"O�IK��՟Rwؼ���`���!�"O򩓖�ڎ[Qr�)U�G�̼Zp"O�`�``l��SQ��2|`��W"OL�lKN�U���# ]�V�:q"O I��) �j�Z�i6�\b��hr"O�AP��Z�����UD�c�� �s"O�XAtkL�%�AZ��q�(E
D"O4�2T#]��ؘ�`G6��P8&"Oʥ�S��Y�R}�J�%��#u"OV%C#��+!8�<�냘G�@I�"Ox��
�g1X櫎��%��"O�=���*P��1u�ǹ%���A�"O
E��摏Z�d�̀'�xe�B"O}��j�)D&V�ᒩKXG�C�"Op��� �D��ɑ�yO4�%"O��;#�W�zW<�{�'� O��R "O�eAu��oJ��W�#Gp b�"OXV@�5r��c��Ҽ/��ȋ�"O�h��埅hHi{� ��6��"OP|SP��#$y"uȗ$�&i���Ӡ"O6da���	T��4%�H�q"O��@��6z¶A��$!0�`l�"O�����B%*�J�1uF};W"O�m���B�|��y�w�jt�$`�"O���Iϸq@�}ʢ�Z=FW􈫳"O���GӁJ� !�D�*6���剏
�����Ӱ\������L�c���%�1;C��07����f˄4w���ؑ��c���n�D@K�dG��'S���
�M�H��C�XjB)x�'a��д�3]�	)�
9J]�}P޴�p@H6��#aP�+�@[L�F)�������߭}�m��	" ;>���_�G�a!��(2����-F�>\$<�gJ�75t!�7B�z�0�'�L� �3�0iqO���	�0�1�F������`x�F�Q�(��P"O�Hc%Hڈp���1G�0"c
y�򁌶R���@WJ�q6����+>�y�f!���Α*TK0��i?���p���@hN
ٮ}��F��~[��0�J*�� ���l�T��j�@�[�O�d��Ժs�ޕ-���ɲMwd�i�O�	Np�U�3-�Pp��& \�ȱ͆4@D(���l����D�߻�2a¢\0\*��<ђ��1V2ع&��J��;��$�ʸ],���"��	~X[��� �y����e�x�����]]T�Ae�sx�3�,�|u���'SpI���A�Ɗ1l��	���G�X�a�!D�<#�v��'<5���Ő�c��a�0V*{�B�c��Lx�8犔 F�3G�U�x��3LO���玨{�yCs���:U�Z�G-eRp\A4�ы	o�m ��14���a��6"i�6�g`��cu�.�	�1Ṷz�g2��y0�3� P�7*Ƃp��(�jH�c��0�"O��(�L  $�0.�8*���j�AK�!˺�P��B����3�(��Ib�\��0��[�H�@Aѡx��C�	�[��5:��#+��ǎ�&g6-�0G�
�Z4��#����dƐd� P��톥CI4)��VX�{�� B\�p�%�Цݨǚ3_4�Iw�I4	&����-D���e�
#A���B:Z|���+ʓj���u�8�#׊�9��(�FD`$K��N����~�;dc�M�p�X`���LQ8L�ȓi��I��K#r���k�!^͐a�ȓv
5[w�ړY^,A��)k����Q�1!o�;P�yٗO�<US�ЄȓAn���/�22_҈���?W.4�ȓN\����r�
t���	#~�ȓ/��L�bOø
�:�� M-0���ȓ{VƵ36��M���QjFm��w�P�0L=)z�,�>C���`G"O*-��X�|��9#e�(�FuS"O�t�`�֥@��܀�ʊgn4!�u"OSc�JǈU
�ό�%C��"O���-�~f4h���*"�r�"O��Jn^�Ȳ����
�K"O�|j�H�]�X����)6��w"O���V�N^�Xu�e�ٺU����"OP����O20��dㅫ�$2�ݹ�"O�r1酶Ct� ���y��F"OHt�� ^.�.��Ӌ�w��"O�zROR S�U3@���H=�0"O(��nݖ�I���"s�`��"O�xÕ�F�z��٣tf�:�L�`A"O8����#=��٤D/i�cg"OR�
��]L��JEnѽY0��ѱ"On}X�o\�3.e�ed,$L�W"O��S!�.��§D8;~�%�"OxS3@(u�l�E-�YO��YV"OV�@���6p䀔��-[�r˜	��"O�Ѷ*�2�8�hcᄂ��	��"O�0Ia�_.`�1�7��C��Y�S"O0-`�I�~��Ep3oT�6�t�0"Oĵ�6 F
��{W͑/*�eH�"O`�a`�2Z����r�J/�B�{�"O,�����CG� 3����fƒ r�"O�Y�U�Pm#��E���� !"O*@����	F2x!t	�>x��$"ON��7) Yp�Dڶ��Dp�"O6Ը��Y��Ҩ:�,
	���:�"O 2% :z�B��L���X�"O�͉�*�q�\�Ъ����B"O|e�B_O���9kç&�a1�"O\(Y��Y9oƥ����n ��a"O5����`ؤ ��BQ�O
�Yq"O��CO�6lf���c�N�b�H�"OF��%��*i��t�[�}D�"O�����]/F�d�1��Ј/G�8r"O�e���A+r�@��s΄J�\R�"O$xۑL�)B̙��ŐEc�,aW"O����������cJ SڬZf"O��5#_9NpdK�g��vL���"O�aI1�Ol�Ke��HZ���"O�@#�E�nX�1�Y8v0�Ib�"O��@ӫ� gfP)�@ �X*;�"O�Pb���;�mq5E�_� �6"O�bw���j���1�"O�D{��Bp�^�x".�vr#"O� N@��
�F���cQ�y�xX�$"O�`K�o 8fK("��bp"OB˦J50�+��_�G��M�"OP�4d��7�2��k��o����"OF�-��-��B7���cq�M� !�ė�o���00�WneR��R"O��ꇉO����0�ȁTj�I�"O���Ǌ��y~q��"m;H���"O�4�vdÅ)���S��!�,I�P"O��j\8J�x��`Kڬg*�4��"O|�BB��C��(��JM9�<ܡc"Ov=�'C�����E���TI��"O*i	tgˏ.�B����:ۢH"O�(#i� lU2�c }����"OD��2��$��� '�5C����"O��pGL�)v�8M�E���pb�"O�es�m�t,�9��T�}B<	`p"O��x��K��Z�4nF?Q;����"Of�Prş��)��M�=h��)�U"Ol(�%��*`�T���%���ٳ"O���U�K��T��*�43�6�ڃ"Od�#��Gb���JO?BEV�Y�"O�A$�I<0=d-t���ތr�"O��J��ˀk��lSè@�h�J�H��'TU�vR��Ɇΐ�h���;�'�Lΐ].)Z!�$�4_b Ҕ��Gi=
��� q5�O�I PN5�ȟ��7G�k���d��w���B"OHM�,\*m�>	!�)U�P����gT�j�̩�=����O��`���Ѐԩ�$�W(���yB;�eSj��DSG��?Q�㞥5���Dͤ>N��������Z���w�{��/ �$M�' ��9R�ނt6�:�O$BSt��'1��9����cz��S6�=�@���'�	r�h�G��K��J�٘U.�%m�"	곇��y�e�]Ͳf�] m��$y�!Q�R] \����s����
��n���ڶ�O
{�\���2D���ӒU���1�I�*�hܢ�E2D�����9���F��(�n�c1D��2/��s�:��oN�b�x4�Bi8D� 
��͚5�uqd�l�d�H�) D���Մ��}�H�q#�O�P�B����%D���dhȄ9FU�/P?. �r! D�q	��v���!�bP�7�$ö�%D�i@ͬE*�Y��%��(vք��B.D��#�#f(��!�dK�OU��Ё@/D�TX1-��JcJ$�ЉI�{����e,D� [6␠/�����.E=�P�
b,!D�kCiF��� ��lYNP1�J(D��I��o�ֱ;��ޑ(hA�"D��1��	�_�L���_#	�,+3� D�ؠ�W��:�a%��O :�:��5D��s'N�fm���!$X*��&D����)��5���E%�/\$@�a D��jB�:=��Q��� r!6�Z52D�@	���%1��Q�Cɞ�b20Y �c1D���dߵi�Ir��=dSJ)���.D�( @S�w��qpR�G�E�:a�j1D���r���c<���Â9wQ��)*D����e��P���7[�Ƅ�R&D��X2F�n�$�$���պ��'D��I&/�?S��ᲇɯb�40
��$D��q�M'a���� �>v�xtQ��!D�����*,qD,���ۘ�|<�8D�X���R)	:��t�!�T��3�4D�� Ĭ�qܟ=��pSa�� D�A!"OPL��ږl��P3B)�J��"O�d8%��CR��ň�"�$�(�"OFUpFď �\y�'f�+�]�"O4�p��ݾ"���5���&x��"O1x��H?׈����-��HH�"O8-P���d�B9xG�2|�D=�C"O�����*R���k��,��L�2"O�5 W�B��"����O�C�"�yP"O,���(�8H�h-`B��R�R�"O����+�J��s��/f��!"Ov�j�����wn�!i�N�+4"O��x.�V��ct-U�e�ܐ�0"O��b7�P�j� �j�8%"On:1�B�5�J�	G޺R���K%"O(��Dǋ�[��x˱&�6�tQ�S"O�)�/��И��2���S "O"���cǒ+��[��[�$qT"O݉��:��Q:viZ�R�§"O��� ٧;Q2U�%��
3� �"O:؂1�Ҟ6}��P���:^��)`�"ON�
W��d�vi��d4��["OA���	���ҳ���J� "O�H�B��+\���"ԑM9�;�"O�@,.������6(İ�$"O�u*��֍.O`��"c�I�~y�"O�9��U��8����L�a�"O<hz$�[��,��C��̅�"ORDA���-D`����c���J�"O$�1���yX
ܪ�lL�%˖��y܍r-���ΊP<�z"�T0�y2UÀ�Pņ>T�xP����yRD�Ul9�Ɵ(X�|T�#FV�y��(%B����勦3^IҒ����y2��2�H������Jh�&�y�� 9��x1 �KAqD!�Vi�-�y�BI7U>$�l@1B���M�yr�ظ]{4pA�bK	+?|q�Ł��ydݺ�J�[$� �� �C!ɤ�y��҉x�H�q�S�g��J�G���y2-ķ�`9� ���=�r�Q4�y򪖷Cs����D�4˺A�+Y��y�]9b<�N@9g�%Zg �'�y�ǯcHxp��K n��\I��,�y򏅱t�|P����5��Cs�W��y�fGrPBІ���S&4�bBҧ�yR�סn���U$H.'%Xq�qG^��y��ă++�Ja,R=F��u�^h܆ʓ=z,������"恁��_�~Gr��ȓM��]�&ٺ_����d2s� �ȓMQ����B�:s�������H�ȓ SB['�ڠ`�p���O�?�"0��a�T-x�%B�IF�Q%�U�m��L�ȓ24��y���h'n��p��}����ȓ,�PÁd��{���
�`][H0��'Th��Љȥ_>	Jj�T�Ƭ��|W\W��y)2�bQ+z��ȓH޽x��!dĘ�� ��݅ȓkitY��"k!�ŀ��	]<J݅ȓLfh8)���B��a�������]�ȓ ����,B�p���G�I,��Ʉ�?��Z�B>�h���w�X��ȓ$����l��M�.���L!P�.L�ȓ�*����[�)�ad�4*|��S�? P�����K�8�x� Ja���"O��QoK�*�hG�I=HN Q@�"OTH%)\sN�j���l1���"O���Q��8!�����'��'�� P"O�(���Q0""�l����l�d� "O�9�f�۽V��m�Ԅ�8��"O
��b�8j��3�e�A��H�"O�0#��ڻ@9x�Af�)%mK "O��b( ��(�߬Oi����"O�����BM8g���os �pC"O:RC�׬<�l���4(�܍35"Of��ֈ��n�a�# B<��"O��p@�t�0����I�-VF]�"O��'@�a���SB�7iC�!��"OBxI�Ϥu��!q�"^/MȨ3�"O��:��N y%����@�.$�\�"O��B���S��	B�mb,�R"O��J�׎tE��	bJ���!�"O�A�:�Lc�
G?.��(5"O�=:��$Q�����ТN/X"O���1��<^���3��F�T1b��t"O�]����fTp�ޚ!�EbQ"O�̲E(�3�Ry�v���a�"O�I���0��3Q,�,TM��(#"O�	Ȣ'Ѵt�s#�R�0���"OpѢ�1N��A�U�_�n��"O���E:Ȉ0ȣbҪ��`�"O�d�%�9��(��Z�b�Rij�"O@��I΅1$ق��.~����"OP�4C���� C�-q%�-�!"O�Yp�יA#��C� �$1@&"O8)���X��X8⊸' ,��"O�P�.�%�Y��'[�A��P��"O �VIȰr^�G&ߴ*sR��w"O@���H�Y�H��қ*vayW"O�)iB�# (�M@�Ʊ��"O��P�+�8T<�-C@�[!)墵�"O��qu`�!y�M:`j ��n}B"OD��c
ev(T�j�_���$"O y�$�!C �zE
�&�0H(p"OBD@W��#JQ�s��#�zP��"O��x3I�Y?N����:]~�@%"OF�[v��.�Lz�J'b!�(��"OX��'_�N��2�\b��ݱf"O�q"F�S'S�������{��y��"OB�s'��B�;����.A`�"O�ZvM��k8��T��\�h�ZA"O�(���-�(5XW��#Yf�"O4�)��d�A�!
�]h��"OV����::���Lٰ]Ju["O&�AV'Q�R\x�&��
���["O`� :����d��OG�LcV"O,��E��8}���q\�5#�P�#"O$|y@F�g#�T�^��j�N�9�yr��Lh�TyDC��"<�c�R��y��ϕ��r���8`|��f���y �%,�0Z���F�X�{�'ػ�y��"~x�� �>��q;(٘�y2o ���H�A,����g��y��ܮRZ��q�8��@�����yB�H�t��!���@>uz$��jҼ�y���-<�b�$��>��yP�f0�y�c� �Ѷǈ�A����$gG/�y��Y]ѯH�> ���iݶ�y
� a�f���M= |���8{tZiY�"O,d�ɑm*pӀ�G�oh�%�1"O�	:��Л?�"M� �!E[���"O��[�A�f�x���"W���j�"O�t�2/��Wh0���UJ� �'"O��xpc��B��Ӂ��6-� �@6"OfPXs�]��niR�_d`�r4"O�d���2z�T�	'~�Q�"O�th�h@~��h�qgfE���0"OT�J��SC�uaE�;6�س"O�QWg@+EU�=(��:pC�cV"O.���ޡ�
��R��4 �p%q�"O ǖ�1����Շ�|*�i1�"On"�a��#���}(̉6"Ox҇�N��r�y"E�1��,I�"O�)W@�=��89,+Ӷ�#`"O������.lT���2g� ��2"Ox�IA��O�*�����J��"OY��Ƀ�
�H��NӀ��7F	L�<a��T>M��5`��4~�m!�H`�<�q'08�#�� �Z���,_[�<��+�3.d�g��(72,@��T�<���;��t��T$I�T<�rCL�<�6�T,e�@`��� ,�1o�R�<�e.D�$R\]_�N��� �TN�<	�K�=\��$�F�Ms"�R�(�N�<A��* �Bez�̍TC�e�a�]n�<A狛?i���*�-�j�(y:��8B�+�^�#!͏I�@� Q퓔K�C�	�Z�,�y�`�<������n�C�IEq"4ˇ��;z,�p2LӮp��B䉪uV( �4炅x�����E( HC䉬t#�ȱ!�~Vر0��E3�TC�	���� C%N��=�cG>3C�|�n;��@�h� �����'zC䉔;� @��I����qA�C�Ɂ0�z����:���
 �5Y�C�s�@A��T�V����]M�C䉡.�$`2�Scv8aS��
��C�M������E�Ril0��K��B��$��y���0)t��R�F3fB��W��H0�H�9:zND�G��?� C��1R�n�a��/~� T(��>��B�Ip��  �9[?����/��S;4B䉨k*�t��iY<5��5(j�C�ur2�!h�bd��1��	�"G�C�i�%BQaӣ!��DY�"���6��'oks��E����~�X	[
�'��-��� $@��p��'�>� 	�'�0�7C"&��i�;E&���'�VY��'Fkl�D�`���`�'��7G�yP�9Y�#Mp�� ��'�l��@M4���zU�0_��pb�'3ޱ�dE��!Z@�+��`�����'h�����/�-��"^�h��DR�'�RYґ�Z,1Ẁ��đ?�x�	�'�f�"SF�t�`��m��x��P��'�r�Q�%B�Hyޜ� C=
�
�Y�'TPA��dm|��4���h���r�'����u��8���u�����'ݚ`�U�V��вE�8a�4��'�n�H��ͳ5��J��M<��D��'��t��LV>P�8���ٲ+=�D�	�'zmJ�J�3&�H	n��5�١��� v!�4���&�b�ʈ�hl�q�"O�ղC��*E�X��IJ!*E@�v"O���O�2'�� {�*��M��b�"Oʰ���`�qq(�,Z">x��"O|�qŐx~t� �g�;�t�I""O����P��H��枦O�L=#�"O�AL���\C�Pr����"ODH���WRfЋ0Iكg�.�cQ"O�a���[mPքP����/�4`�%"O�#iʪ�*b����"�B"O���f%R�[[�dG��.m*@��"O␲��/�~�9�d�.Vs��j�"O�l���ʅ�E���¼$ ��@1*Oqx ��	{: X;���!�=��'s~�:f�fv��P���s�z5��'�B�a�hV*9����h��9r�e�ʓ���1��&V��xE��U��نȓf`�њ���b��+4G�Ex��2 pAR�E
3�:��Q@ƳD�	�ȓS�6U�)�V�X=��ӱi�m���� �w��,}J��p%� $J�1!���xi����`>Y�5Fzb�1?Q�`ݛ^�l0����_�}��L�IS���O�ր��+K�H�^�H�f�k&&(J(O �=E��\'ei����T�E`0@�~1��r�����Hu���k�b�;6�@$è}���	c��� ��/(H�� �IZQ�G/�hO���nfy
��d��� �O�=�~ꆂܣL��5M��}�.�Ì_}��'���P�e
-�v��u��j��d1�!80t�Y"8�d\���3x	ΝD{b�O,J��2`N{���*WG�$*~�QP�R�)�'�M�*�2M�в��G��&���~�F3}mZ(Ѱ����@"�/H#;:p���P�94�����L�atGG����H����iP�~�8C��F<JX�����&�1�g�ʳ���~r퉁H|����N n�b��H
o�v�F{�O����%�5n�nx��E�
�>�q�R�)�tC�6)K�ؓ�ı"����fԙ���0>I'Əy�����e	cPp�cw�J��t�?��D�"Ub1&K�S�̫���<I���S88�;4C7?�r�a��{�V����>�S���T)"ɢ��A��~����v�����'�ў�O���cУ=p�h���A�l�كO>����I�z�S倒wX�d��(e��	U��(��j�F�5tUj7�C!Y��@���'nў�~ʳ*R"�TU��DC<��� ��HO��Q�Aj���@�^p��Lr��O��@�8ò��L�=b{ E�B"O�H�K�+�u��XZ���ؠ"O@������挂���x՞��d"O,����<N&�h��V�1����P"O`�s��c�P'���܋""OB�k��+�|��%��� S"Of�����1���BO�$(��03"O�b�n�(^"�90Ɠ:�h`�"O�A �ɖ0J�؆��}cX�i"On	!k- �۴��'J���"O(�n�	4fe�pl��b3���"O��@���������'m%�-��"O��Е3m
~�Ң��3e�"Of�X�D�X�h%٠�8ܴ;'"O��c�'��M��l��n��P�`95"O���s�Ҭuyޅ��75Ol�Eb�<�e땝B=< ���7/kPИ�]�<I��Û<��Yj
6,������[�<�Ƃ<#�4ؘdo2P��P��Z�<� R���eY�w���C�TZn����"O�E��f!2��u��KulM��"O �¯�'ZwVM��'�*C^�p�"O�� ��Щd4��;}����"O��bѠ��e�X ����g����"O4E��I�cVdl�3o��D���!&"O����_�kx6]1e�2>��T�"Obq��䀴q�v�H�d��t��'"Opg�� �bT�U"R <7��R�"Op�1O�+��)�R��s	�	;C"OjI����	 �܈�L� �0S�"O^���i�A��!�LR;^�Ř"O4�8���up���!oet��G"Op����w^y���1[�L=�"O�dP`d��Pi�
�rX��"O��g�_�^2���uG��>���j�"O���4��#t��	QU�˪3�$Ȑ�"O|}�r���s�j)WEگP�x��"O���"�4|O�yr7&�QAL@�4"O|]�o˷vO� �%=5����4"O�Õ��s3>h�qCI�v�n�"�"O2���	�D
��:Iڞ�ؔ"O>�Ǫ K�`:���a�r �f"O��g�����wF�YВ�� "OƐx��!}w��Q�%�/�h��W"O�mZ�E�^���4
�B@� "O���%醡>�,�f7Y��H#�"O�����y��89��	ul��*"O�ؘd�
�x�2� .˰H
"O��j��24,̀yF�.:!�#W"Oءз��~"x��NF��;1"O����T�/2ЊR�^+d�qd"O�DJ��ĕ-v`K �l�|"�"O��%�T�MԄB���<\ںxP"O���C7P(�s�n2��3R"O�R�*���G�](�"Aۂ"O��;��� �>0��n�&kl�,�F"O.�c�`J=gl�A�G#6[�"O�Ո��>;��PWCR�O���"O&5#߽It�I ��n���W"O�����(��8�1"�*��(G"O�c`��b&@d�_�7b@E r"O!� 2o�f	�&�L2�qa�"O����Dk�B��������`3&"O� I���� ����-+x����"O�YE���s�����?7�Zm��"O�e���J � ���!�Sm*�x�"Oh��P�/���g@�Gi��S�"O:$��(]>]q�}VA�*!�����"OBu[׬�1}�6�7�;�p�aR"O������	V�	�eb�$yF@�`"O�x"@��+t�����j"O@Aj���'D�t�ٲ�X
�X#�"O�0��i��n�6� �.L�d�DM@�"O�y���P-^O�ڵ@3��J�"O��aC�9�����
Qo���5"O|����N;J�Ԙ�����,��}Ѡ"O�e�lS��$�" ԫ�~�('"Oz�����qhT��.K���4��"O\�f��$�1R�lN/"�Fuc"O��%��+bd���i�/Q�n��"OB5m
{���rmS��h�4D� ��h	�dh����-N��Pc�).D�����Om�|#�i��a�3�-D�� �h�%�	3�(��!� �fIPb"Oz1+Ek���6��rz�H%"O����M(W`�`D��H$L�R"O�x�V�]����B^*�ȡ�%"O,0c�V0j3T�ɰ�A�%��A"O�Q�2gX�Q���(q���"O��`�S;� �(a��eV��;A"O��!���1�����VΉ "O�	�p����e�84B�۴"O0� �c�2Y�<;U..عhQ"Ol�Z��!?ע9�i\�.�(HB�"O���cP�g��0�E�+G�Dmj�"O<p�떨6�@�:��	] %��"O4�"��̀L�ЬÑJ�fI�	�"O>�²��7F9+jM��n@��"O�h��"�+1BȢFȐE�ܵ�T"O&u+��O�A����T�P�OŊ)�Q"O�eq�I�<���"�/jf�Jr"OL�Ib��!�lE��Pl��Mx"OjQp�!�*�H՚�k�%6�Ҹ�2"O��˳�, r���\9m�@���"OF���'hW�(��@�s��y"Oʘ
A�D�~��ݡC�D5Ci� �"ŌX�\��+��P�PN2��"O�n:����6�Q�ֈ	��?D�Xx��:>�$��OWK��X(�H=D���B&��_��!x ,l[�x!�%D��j4�F�;ty�a�ؔ 'V�a�$D�`9�e�+��{Ҁ�<S b�1�F=D����]�>+�m�ւ$��4�(D�PK�郠>����oY:4
4` M'D��6��6 >6�W���S�E�%&'D�@2��<J��ӱ��f(��� $D��s��"M��̛99��2�E#D��aé��t�����. ��`K=D�����Z�� K�+���it7D����ś1NR�J��4`�q�(D�p ��H�b\�� >���k'D��@�P�i����9�����'D�X1�)a��P���1V�D$R!��)s�ĥZS�6-�p��'�!�$�&6jH�J��H+p�(�HU��,�!�DF�e|xSe���-��ԡ�J!��3 �r�r�\�sY��#�/S�
_!�9(�L�BK�Dv��u� V�<��� <RnZpT���Z���as��J�<��� �}�4��'g�+� @��E�<)���]j�HѲ�! ��pn}�<��O\��#7���L}�����
T�<�� �7�����I���C�y�<a����:�ڄ`��!C:m��Zv�<�e��[  B D�,0���	;�C�wv6�p��<z�[���ox�B�>v��T1s��-!�-S�΅�r�B�I)@��0G�Ѥ|%�@�L��JbFC�	�Ph^���3�v�!�m*!	PB�A���4%Z�l�bU��$#8B�	�o�b$*th?QD,�Ս�7- B�ɖ?�������:s�z���
ɁV�C�	=2�ae��V�6AJ��ʚM��C�I�2�f��&]}[AJ�%M]VC�	�@R�8���,8҄#D�	J�B�&����-X�AYX���˘U�C��~���L V5�B�K�[��C�)� VY�/�B�Ueʟ\<l��"OR���^�
UY �,m(ݲ'"O�t�$g؟hA@�F���|&M"�"O H`�N�t��H�Q��R���"�"O`�4�C�2�	P��I��r1��"Om�4*K��1WȳZ����a"O½��)�.�B|AG���@U��x�"OLMQ�&4����"J
�23��p�"O� L�F���)�~�*0�"O�my�-�&e[B@K@!�'��	x�*O �`�`@�*S�т7��qD� j�'�
��c&\_*���3cXQ@
�'��뱌v[Č�#f 9	N��	�'/����'ۏmL�u9�Ɛ� �BPX
�'Y��PwCձz@|h��}�H 8�'���r���TX8�S��x&��
�'�b�Pp�ٝ4crl����:F8}H
�'2�u
Q��,;�]��]:z:�m@	�'94�����`�F�'��: ���'��5#p&I3��)����2�<��'�PM��JZ=B@`B/(���'�၃ͥ*�̌���0I�:��'�p�9b�[�2z����@�xE�)�'X*��,J���RM�C�x��'��)Bf@=;(�\�:Y�@�'���
R�=ĔaKU�I�{���'0�X���S�9<�:
�*\�pl��'�\����e|�ܳ3�X.J'���'��\bW�I�%��)A#F�v`�Ma�'�L�vC˫ �E`�\�mؐl�
�'3�#5�J-�4�	ÅW)_fb�'������V	$�Y�d�'\>f��'��('��~v!i�ǋWM��'���DIb�4��,�Du~D�'\����>���)���s��m�	�'��
����c^,Vm��s	�'�������7c�|��C�/W!4���'���WI�t됇��M�P��'�tx���WF�!�Pl��:��y�'��C�Ĩ\|������0�����'<d5�PB�>���a 
�Q��p�'���4"�^
�,I�C�f�
�'���0�� D�8�)�O�9����'`�!�/W�=�h9���?4�~�"�'�0���2tK�Tۆ ǻ+��(
�'|$��a��t��H6���&�(�	�'�Zݰ�����;GnԤ��h��'�V$zj%�0 �VEO����
�'���áY�Vg>ӣ���^8a
�'�q�E��<N�������A
�'�(I�   ���   x  �  �#  ..  �7  �B  �N  yZ  Sf  lr  �~  ��  Ŗ  ��  y�  I�  ��  ��  p�  ��  �  E�  ��  ��  �  S�  � �	  \ � �" w) �/ X6 �< �C PJ �P �V >] �c �i p Sv �| � 5� �� "� c� �� � w� �� �� �� ��  `� u�	����Zv)A�'ld\�0Kz+��D��:�2���OĴ���%�?Y����?�fY$E+F@�S�Q+)���W�Z%#BD5��F��2�˅NK>36H�cAՅg���+}"��	^�g��)K9�Ar�/�47N�ib�]�����Nɖp�2�EU�F���%iX�}�$�;g�5!�'�?9���[����cH(|ɀe� (@,�f��ÎСl��䇙uD�9YV��!A
7�//���OP�d�OH���9q&R$��=3
V��gc<�d�O����O��?�C�ށ�?q��?���Ҵ~�@�Dmϋ>�.�zǩ��?!���?����?���?鳂��ӄꜦN�6x�d��i�$b�r� b�8�J|�vAj�H�'s��@��T�ca������2
����]m�l�a����dh�hjU���pI������	 0&�ԛd���|8�`�4[;��d��y����d�I��S���O
�G�T��p� "X恣v	�!_R�h�nlmڣ�M�f�i-bij�f��1D�u�d	��;z�9#���-W��@��l�\0��ʔ��HO� ����+OL��i&kC.?���t�᭻.�����o7%?�CrA	`���b��)l�pP�

�$�n0�ش$\�&fjӬ�	[�|:e%H��Mk��ZJ�rL!�Ŏ�HIBа��>�MD��q��IQ6�<��e�*��1��';� 7��Ŧiz޴L1&	��n��[wv�s��<��A�G�0saD�\v��a�`�l��w�ٸ�%]�;�$s@�s�x�e���4�ڗ \MZ"�I�H�Y��PK-|¥�ܴW+��v�Pu�r�H�t�h���[�	�$�RԌ�B�(����=-ڄ@a��d�Z9m��u<���g�$���Z�z=�ǉ�O��@Ҁ�� `P�yHȌ.,��2�l�1ܰ�@���	ҟ����?9yF�I/ت�3����2#E��B�0K�~H����G�����	�O:�Y���X���T��U%НW<2-�ߴ�y�֜90R(�T��(Z�FEҵ�Љ�0<1�d�Z��Qju�޷����"����ʎ%g?@dY�a�y�ax"�>��$�FyR�T,��yz����^I��`B��?Q���?1H>���?�)O��O�pwRK�ʜ�c��H֯� 4��d�OTT ǩ6ƓO��9O�ɂ۟�����0��T;@��h�a��.�O&ʓ D"�h��i����z�qklO�g���#t,Z�48�(�O4���v�lu�O�R�X�RPj#W�\a����::�N�a ��(�t�[��ک^��I�=�i�%F̬C�X��d �	rd�Xw��aqj7\.�Ti��6�4I�G�U���� ��dO�=��Ky�� G�4=���7�A�"k��#��P��s�'��O���	��kA�
�
���Z��V��hO�IŦ��4�?Iq�i�D�yC�)!V�N�'"��o]`���',�	a%�!��ӟ��Iٟ��'B %�`�E�^r�U2��
���������c=�ָ�kK����?�+��xҢ65
�@��H�hU(���!��?Y��RBGݐ@mJ��G'�	K\�Y���j��@?#Tp���5� 8ch�"\}���	�t^r�r�+j�쀕'K^������̟�'� �b��.X��p�S�5hr�4@#�'�[���	T�g��&�XE�¨�0XL�Z7����Mc�iMɧ���O��	3�x�s�:{��ZW��T�n�%G��D�OT�$�<)/���(LR�	%@ҽ;���Pb�<Qv�A�j�m��h�c�thD���O��ޘ��E��rL0�5%�5����H#uoTif�l6p5x`��-\�B1ʴa�ȸ'�e��c��^7:,!%� p:]��̓�?i0�i��"=��2@-�����ȥ;t�`���B���'���'	�H��GR�DTf|�"�r���N>�$�i�l6�<A5�1C3����LbċHk�=�Ў� ��T�"����T�Ʉf�9�	�\�	J���aU�ݫ(�8���4�yKVB�X�N�WmH�c�ɛ�0<I���'D~�tkrO�b)޼����0�f���&�=�^�sB�V�RYF(�s�	%6A���BӦ� �4�?y�*�A|�%2�%�9(q��0u.����O��d�O���)��h,�)��l�:L.�M���j6�"�t��!�l�yTF�p���_�r�Pr�٦�'%��BT�e�V���O˧si`h���ʒp2��O`�$0�R��b|�����?���Ͼ���	�`��=�X�Y 1��O;�D5I(���"�h֔,�x�Ád�5��U�'� ?a�e��ѪCJ�f(�M����E]�)a���:���q�'��8p���� ��A@
��\�'(@"�=	�V	2�i&���S�͏F=����Es�^�O��>�D�O����<���ߋj�
�IA+bS
�@W�.@���x����M�
7�v�'騙���2r� �l�]��h&�z���d�O���܈b��d����OF��O��iށ���5��Eb���M�J9�"%lPTDP��f��IHt)�+M�ʧ�J��=�d�vϼ�S�A�C���lڥBި`
5o��D�GnG #���1 ͎F�Z�'-�j̚wl�ȼ��KV.*�Й�<��gע�M�ó>���@ҟ��|�	ݟ��ɸ-[ !Pd	V����f�z||��П��	�����s�g�DK�KUTɫ�)��5g��g�^���$�M{�i�nӴ�����	�|�a'�;[�ŘG��(����C��s]�<a��<����?��4Z���Od�D�O�q�@!����ce�9���3fOH����/�;v�`�0������DU�MD&U�u�Ōi�ddp�d̙o����/ZB`�0V���Nlb��!WҦ͢M�+��%�Ժ�0?I��+=Ƃ����ôN��$ۦ� ��$$����g�D�Ɛ�e�ko.���]�Iğ�&?!�<Qi�H~�e�U�Ըy�����T@�	:�M;аi��7 z�#�4�?�'.d�墓�W���b�;C)�5I���OF���1����I$%�!l9� �1:�&B��Tx�@�ߦ*o���Q�����؊�DŖ���Cb��b]����9v�<�P�;r�*H7��cn�q��A�
�J�k$k�Ƹ' �5���;��H�<���֮wC���Y�l2l��R�Y�	v��OJ��f��&i�%i�a��=�4���'�l7�ІZ����1 �;NRH9�� ?o��l�syb�	R�7��O������O��"�M�Yg�D�#��u��鲴��Ov��Ͱ�0}���&j�$#��l4��0o��B���v�R%�WJҹJ��Sg�ֱ@:�A�'[Fh��,C�s�|��R7��I�ĆD�E�2d;&�	#q����L���A6p�R]��e�[���'唥��(��V/�'��t@�2-�<r�$?)��@�V��hO���]8A̜��t��X�ҁ�؝5xў��Ɍ�M;S�i��'�⍫�Q��tL�p��1 �<	7~ӄ�Ġ<a�/	�����?9�����	2i`&%��aP�`B���A؍_G���g�\�??�AZ��ڡ?�y� �|�'P�"�)u#�Y?��C��^��PqĹ�Ţ��XI��fm��Xg�C#���1�4I�q.��5i�h
/ow�nH 4tي'k��y�hQ���+g�6M�vy%��?�����|b ���� 3j�8o^��b�G'��O:�=��F��ե�PE(.��k
.�y��'r��j�H�l�C�i>��Sgy�K�<�4�1�I7@ ����)+���ӵ�L܊��ٟ����u'�'jr:�`]B�a��0>0a��ɉ�*�|Ӂ��#KǞ	��2�r��G+'���?�b�)���h���;>�Ti�rIT+�М�1o�EY�Z�N�"�1���$�yY����ď d��J�H_�a�μ�w�'�R�'��O "|��F�13���c­@�H���:���u�<Y�bޏ[��T� �Cd�s�r�I��M�����*'�YoZ�p��� ʌ(�L�8j����+�>��̟L�n@㟌�I����e�+���58�~��&�Q��l�S��$XA�hg�B�q
Dc���
6��Ar�@O�wo�-�p3L��I'aXD��G�{�*��2�YN�t��!�0"qO�Ő@�'��6�F\y��2y�Ztywf��<����۫�䓒hOq�-X����~P��'B�('��1q�'�.7��8c��r"A׆*ETL@ч�>8�o�uy�"D�3�6M�O��d�|"�@��?r��0u;��� �Ʋ����j�?�?Y����������D�O�g�DQ;��u��(@A��G��H�O�� E�F3;h�2��݌����4s��%�
��n<�F�Z��  DC�O4�l<�H��SI��J��nl�2�oɝ!��|E{J?-xB���4�8ak��/ƮЕ�<�xr�Fay��c>�� ���	]�=y�.O&���ꦅ��ݟ��	�p�
q���0�IƟ �I��6M�8s�"ň#"ĄF@�J�'�0]��	̟H���ٳ4-����(O�Hbv-r@x�q祝�L���q@=v��AI�b�M^X�a��͐7�1�1O�|1S�]1g�~尴dI�!�N�уgk�6!�'NT����ʟ�'En`��w|�c�_�Н��0ړ���^�5�Z���ǚ�T����B�iC�I��MS�i)2	~��˧��-��Q�'c	�b�����͗
�& ق�1Lz�{�(�O����O �$K����?!��(����+�z`�
z���(��L�0j(���'c��2 ���^]D�RF�*^�4�fM�	GU�lyG��2u� ��n�P��Q��ʝ-��Uφz��[��m���R��'j6�XE�'��`y� E�03@:`���]7rIд-�7a!�$@�T|����[-G�ѻ�.�fE�C�v�����ٴ��		c��oZ͟͓Q�	Sg�/+UF�P�#<VU��ty�'�B3�dp(��
a^D\�5j�Eg��xT�Mo�����YN@�	���A=N,��V�(O����|`8��ҷi���	�8����h��[n�Be�Ʒu����+ n����|�I�o��������,O�$��m��Ab��?�$�|��'��d{�F���8P)�W[0(O|ʓ�hO�ܦ%I4lX�~��B�W	%̸�W���&*ON��T��m�	uyBR>i�I5$J\3�)L�0@zPh���I��ퟜ#ѢI�_�N�;�$/
�E��$.��!%
5��GP�}��u���uf���"����N5�(�����/�2���S#A�8��遮f��t�����Բ Z<9�v�z MؖW�I�星���@�O�un�3��d��O�Q80��!{ʰR��I-4d���L>A��?������p�H��V�%�A@�e�""Mn�t�|�U���I�����<!�O߰3�m�)�ܨ�!��)���Z�i�r�'�LB+ea<�r��'V��'�R9���`�K4�9�����<�g�]�)3~�*�h	O�5�)�X1���˘�~r�Y3d�D�s���j�-b�Cϖ5��j��$`7��;���!~T�T ���B�9D=,��*�т�*�'�t���@�Z%JH>Ƀ@�����|�<��L��2�d�R�ۈH�vS�Xz�<1��C"_W�A��G�G�����xy�+��|�H>�����js2����;%�52ݕb��Q��@���?��?���dr���O��`>!*d�T�I(L��Ę�>�XyE��>c6��� ��nRA� ��g�Uو��'=�� 2�a�-��>7����#X����Č�� ZJ��k��6Ar�q`딼��'�>����Ўtex�k��?���!U��?��iL26%�I���O�x��0'ǣ$6-�p����Q�
�'[�U�¦��6�f5�	T[��E:J>еi��R�P%��M�͟�Ń��_"�hL��ުC��Ī��',�I�L�	�|�E#��(g�����\?��-�����R���P'/'�}��G�$���#­d�ԣ<A��S�S�����R�,E�$bQ$B0^ .�pD�S1k�ƩQ-8t%DP����s��+EM���p���	��M�sZ�|qR
R�
�)��\�C�u�6��?ړ�'w�����բ��!��N�=Ui6L���i>}�45t"A��e�8n�Jc'�!9<�@D�i��� 4����ٴ�?����ɂ<$���hE@H��B��x��E�L�n>���O, Bk��n���aB�^,�m�A�dV>�sh��a�R�zc�5P�6�02b�X~�B�0]Ӳ�q@AI�b���F�Ӻ>���$�",�h����Ы�OrT��'�T7��O��i��K�@�S�W,tP�e/��R��y��Ʉ��a���G{h�F)H�Uǲ�?�v�i�6�6�Ӄ6�"�����'��f��/.Z9�'��'�\Рd�U���'h��'��J+T1��G�-	B��g�3Fl����H
C��P�f�LQP%��R>)��v�'�nщ��E��� ��[�$�r��� _���7o� xx�i�=ъ����2���2����<����Dѵ��Zu:6M�Ϧ��ɁQBt���J�gy2�'���4%M2�hFa��IF0��'/2�'���a�� ,y�@1�Ѣ��ovE��_����4,�֑|��/&1��W�����HU��!=��"�g��������4�	������ug�'9�<�
 �wC��q���\\tʧ`^LZ\� ���T���x�`�=F|,����(O.��UdY03G������2]��i��E�Y|�C�"�3Hl����#͚l����+�(OF�2��ʶM<p�Q��Ή!���2�L�"BFw���Ez"�	
9�J<���ʴX!��4ŗ�ye�C䉚��U	�N�
̹�P��SԴ�O2DlZԟ �'�(�y� �~���pm���c��:�X	��_�vR�����?IF��?9����dP��!Џ�6A8��1 �	 08&cB�C����3}�8����.���d�Ŭ�0��IPlB\С��
|�wl�#�>I�Ǝخa����'���(O���$�'�B��4�7"Z�J��(X4H� ��]��!�:�O@E3��N�?�0��kL�
�z2�'�����.Y���K�%�6 ��o�1 �P��*��^��M���?)-���(�f�O���@�W6x>)�$ �@m�msC*�O��䑆xv2�{�$P/'��h##K׭$̕��O����/Eİb.�bs�5@��>U?�>��c(��N�ڄ�b�! $A�jN�<���O~�R��?�@����B�0����S�b�'��>����d㉫j��4"�V.Y�6��ȓ|��p�C@7~�
EIӁ�j��9E2�#�'<����3+��?�Z�C��U����4�?����?!҄�H9ڡ���?9��?!�w��� gߒ~��S�`ߺ+���	���6.����"~8��S��	��O](}�!m�W?D��&h��a�='�iKr4 ��s��/,�xbB��E�h�|R�d�qߴ��04k���k�t÷'�5��o���ؾ=�2�O��3��kв�Ö\�#΀$6B�ɶAf8;F@åYш 17)^l��˓rh���Sџ��'��ؑ o��GYD�;�`ʉ�>Lk"�=�^p�'&R�'���O]��'�2΋�K� �GJ������T�6��=�`.�4J�z��Wґ	'��PoZ�':v�Õ�B>�\t�T�I�4$H�����ъ�6�؄���ϞD"9�۴lI�9H�{B/N6�vHٔ�P�b������=(~={������5�$�O
�d:��5�&Y�Ǡ
�Z6D���h�?�&$%��Ɍ���@�-�8��oƈ�!�ђi�'��6��妩�'���I�g�����OdTQ��Xv�ڭ��I�?��	��l�O��$�����Of�S�A�p�C띦/�b���ʎE�Z��	Xd���#�q��P��:��O��a�E���r��tz5�Hc��p�j�	xH]c�%K�*�1�o�(Oh���' ����R�G�?ά@8��I�>}0�h6��+�O�4rì��<�J1�dL%fv�y�P�'��$�r�S3H�!Y�����G�2^�lC���M���?�,��E00H�Op��ΐi�f)��[���#�K�O*�$ؤV���f��"R����
NYP�b�OS�S�4��]��/<�2mxuH"}��PSv���ҋ-d^�:����\ua�$�ٽ7ζ�OwxT2��R�K��� �& q�ep~�II��?���h��牿g��d9�,�8DS�|���T/D^lC䉈+u0 z�( %Z?�X��=��?9w�S�Xd�ٚDj�>��܈��Bo����Iןr�E�x�Ҹ�	ԟ��I��λd&��{�Ň'Z�J	���  ��ye��B-���&(

?�"�yG�Ç��'�](1�L`�3Di�< UF�@SNT i L(�ܬw�T:��Ř��OĈJ���C?� �p�,�,"�2 � % 8$Tv�'����p���O��=Y���.Ê�Г�
�+#��3bP)�y�m�J�6-"��� -]@����4��d�}�����'��I'��i���#[:t p�O&>ih�����!1T�}�Iܟ��	Ο�iYw��'����Z
���4	����΄9\�	#�c������z|��`c�@�<ip%�2���U�2��g�Dа��H�r,vt��
	"+b��A�LM$�� d�ɪ~�R��Ѡ1�a4 ͽ%/�q2t%�Z2F������Jڴk���Gx��&�~�H����*@�Х��yb�%�θB� M10/R���+��OЛ6�'��)8T�u�޴�?��4��p p�R�{bL�ԣ�%v����?Yb��'�?1����$_��?��y2�'�"�ДfЕY��{Lł�0<Y�ǈ�'�$��
��R��1�dMZ�{
�W|������LҶ���pB��a7�u��D�B���@�;�d��c B�^L��	��?Ѳ���w�#��|���\s��*}A���ٴ�?A�������V$,A!͝%m�p���
J�l���O�E�����M=p�$��'���Mx�PC�I�C�]r���1:�I�%�%���Ѐc�(`#��S��q	B/9��2;;�!1%C�0e=`�p��so��b�z��I���S�O��pXA�3e�R `�O�eָ	Y�'(���T%� ��ɡHZ�fYԫ��čj�OoN%H� P��XQb�7IƐΓ�?y��?yU�9���?Y���?��w��鉁��6B �٘�Ă�z�.��w̛*�f�Rw&ېbm.�(׉ȘO�H�DoOW?1�o�I{ƅi���*�L�����(g�>I�tA�y�u�0k�*/:�|��M	"@��I�*�:�P�/��X���\�5����K>�������|�<�Ԯ�jQȹyG�$�,�1w�BF�<�#�]�
>�h�!`L�'�4:a�CyR�9��|"O>��-ꤹZ��uIZ�1k^ ��'T�T���O0���O��)�O��o>U��g�i4J�3�a�-*Ze�Ty�F�V宭Q��[?�.4�F� P>Q��y&EJ�x��tQ�p��&�o8�Ј�u v(82/�|`�4P�&O*;�j}*��D֦B�`*�Ԛ#�Ե� ŏ7sL����'�j���\�d@ys��U� 5�ݒ0-Z�?c!�Ʀ��k��2(0��ܜbv�'��7-8�DOG��d�O���P]κi`���,��B�0���O}C��Ox�>uլ���u��-[t�,�ѥ�<6|*Kg^+
2$��� 	 �}��$��Z����I���I�
� ���ɡڊ3�m�AN�$*�j�k��N|9�`�I.%���Mx�I@��u���r8����\�Z�C䉻w�l�y��G�:'֠R �O�C|���$GğdSEZ	d�R�XtlM7K���P�;��>/��oZ�����Z�t����m^�f��*��q�����k�b�'�,�x	�YYjљM��'��i�4cT����ϊ�� �YT`��{�I�b}(�n͂$G$��%�J�
�2#|: dB�v�=��jD5��Ikd�s~R�Ո�?��|��铸T�Ըb �Ƽ����2΂	'P!�dʰB&�����[��LL㒍�Cџd[����{�� �s���'���ˇ���WQ�7-�O^�D�O�!�+� i�����O����O��]�5rR℗9q����"��N�����~ybB�j�2���y�)�)m��Rƕ6k|�y��	,����A�D2E@��Z�E֜B\�@���"��u;��O"��)�_s@���%�L�%�\�+�O\c>c�X""��kМ@�s �!�\Cm.D���u,_�֘A�^,r��,�<���i>�'�{�!��Kn���мY�؈Ig�˘W�d���G��0�I˟��I��u��'��4��U��'T1DZt�t�>_�t�8@���g�=3�A��I#�t�V�ٗB"�s�'(�(O�=#�A0Q
�:�`�1}�L���
-W��0pa��/fh�["!��K�dh{v� 6�Y���� 3� ���#R���,K�RP���'5���Đ4#u�E�vj���8�*i!򄄔Nf�x[�G�4�X
%&��J7�'�7m,�d��QY�oZڟ`��9�����bH����反ci�$��ݟ�%�Ο��I�|�"�E�\�P9��S^�����LR"i�*x<YsWB!("��I�~/���B*�X��!��&K���
/@�N��`��z�Ȉp�]|�Q��"$i�O�c��Z��F��a�!�Փg�J;D���E�έ,"4)�����h�5�<�O0,�I.J%���O�9X|x�:�G8�ΓOB��wc�����ԟؗOˢ Q��'p�@PeE�8c�eyQ�A�$@:yH5�'6b���!�\I�b��p�*����O�SP���T����/er�(��	����2o;�\;��	B0RQs`�S��(����T�ũ"Gq�(�#6^�:�a\���Q�?B���3�  qBE���=/��I:i�M��"O�h#o���%@r�� G�(��5�I�h�B���g�t_�]� Z4��F8} �V�'pb�'����%!�+s"�'��'��N�	h��(���-'���'�8=������v!t���J��9�"��
d*h�i֔n��!�dl�_�X���b��Mi���	H��Y��	׉��Ʌb鲠�'��EB ]9B�S3��c�@B(�O���F'~�1��U�?��%ٵ"P�.�!�У���i�`7r��#��S2Y�=�HO�	5�D͟�(<��h �5�c)�<.Bu󱎟��J���O��$�O8���?Y�����)�!6�٣���;L�X9C��]�B$}!$���mOJ����)c��yRJ��_^�J悑
K�r�V$�%]�\��'H$SHX����Z�X"���"
|�'x�D��+`�̤X���V����!���?��'������� �J5z��@pT�X�'T�U�sj�.����*�DuV�(N>A�i�ў�QD-��|��&[�B쨀:bbO�8A��*D�X@�%��~	�O,	&�J��'D�hP�M\x�����*��p�Ч+D�H�)^I~XӢ��M�
(D��16���x\y���K&�P�"D��&��L8����Z3d�p�&5�+�LtG��L���JQ�dNU;��Xc�y�͑�q���JK	Du��@�y�Ҭt]Υ��K�I��pJ�k��y"(��NOv��U��F�~���N���y�+�6.Ă�h3�H/	�J=���ψ�yR#̥<.� �����7���?�6�n����Nx���?*�,�(�^�j� t�"1D�\b�h�Z�lh`S,���--D���H̐a�B=�EcO� ���C�%D��QB��Tin}9���i�$�j�6D��H笜�*�m��	"�	��74��ó偺[~}�"�R9,૰·�<](��$�O@U 9 ��G�n�( A�*\Ul�;��ֿ� ��<l�KʍZ>���eƃ�y����	�&��OL���OD�w���Qr�L�`a�	hVu2�kٓ�u'K,J�t=�t$�6\Ve܈O��!�O�7�B����P�v!�X�^b�h�./h���
�k�6�1Dm�8�(O����'����I���bP)+Z��#"M�9X���a���i%`%WWd�!��Z�2�!�)�O�x�'�b���h�'v���De�Q��*O�-�'��O� r���O�ʧ TB���?� ��4�r��Q�@�8 IԄ���?q�D��sE�Uy� v, �[sƂ/w�`̧Tvl 4M� �^��d��`>�4�j�|�ْ��y��%e�(g�l�� ���>�y�):��
�%���!.m�(�'�O���,?%?U�'=XE����3.լؒ��P:)��q��'r�R�Ŧr�T,��eL�6������d��O��x4�(;5��z����Nw�(���U285��'�X����a�z�)�O����O����O6�)�h�����^� �T�b�4��@�&,J'^E>	z�I�Af<���'W�u��퉚'd
,�TmQ(e�(�cC�8��x�&M��k2 ��������t�L�tP@�''U~Zf�+�~�J�@:?	��П4��x�'���_ǈ��*GGNY�aǽ�!�D�x����P�ڌ,X��ѷe� �B5��|"�����7�6e`��J3�™%IE���c�DKD�ʤ��O����O2�)�O���f>�� �A<�-y7�K�M!�M�B*��XXl`�b]�g�t�D�(�@Ge�ABB-�Bh��<YChI�u��E2e��7	�t�T�$�:V��!G�:ʓr'���	Q��a��@CE'�1�� )iT���Iz�'��dr�I�'�`&�
�M�sB�*D��K ��$d7$l
@[�dY�Ef�<iG�i��Y�0�2�J����f#^럐�'E>�$2�B��Q#�a��	z��I	0��������/mQjp�r1�~�*G:��"��	��a�HU$��BO�H��iF|2��-�)���`�zE�aO�-Mv�E��nZ�Z�J%K�N7D8�ՈB)"{�d�Gy�)V��?��ݘO�ܑ`q��|�6���s�8�*O���DI<+�D1璗|B6� ��ܥv$�}2�<�Vdݼ`V P�P
/�&t[�dX{y��C�{92�N-��^>UR�΃�?���$D�uۓ��(!>mx5H�/��q�I���,k��W�d�@�A��+DX5���4b>���ߠ)��3�N�7��$��*n�L��S!d�*I{��:n�>$�A�9�>y:&�I֒W�PISg���c?�L���.��U4u&��'H�)�)/?� �m��8����'@ES"O��@7[	L���gdc�X�r�	��ȟ1���FE�j ٓ�ɭ\7��`��O�D�O���f�{�t���O���O��)�O^���G�� R�J3��@N�3�0_(T	2&�'��{��B!#YB�'��'J�y��d;'|rQEnI/M�6�c��ҭi)� r�dW!R��ī�hG�����5p���L�s���'WtH �n.lس��2?�0����	i�'��$[*�"N�.d��d�d�_-�!�D��)�$�/�����㢬�z(b�2��|����$�u[j<z�đh^���U�H�ѡ�l	� Mh���O����O8���?����Db�.3�Y�ˁ�C�Y����r�АKƍ|�\�'/��{�<Qb�-�p]�@��K�zGP�J�L�:!�lH�� �r7�-K��-� ���Sڛ6�7p�θ#V�|B���?���̨��q5c�`��[Sg���?����2�}���nEZ��*�mEO��݅�IR�'�̘Q��ʛqG2���aF,EX)s+O8�nZݟ��'��y0 �'q��'T�� M���!mV
4E,h�ņ6N�X����'��:wY�Y�b�ZH���D$P.+7Ԑ��\c���c*N�IGĭ���̿2�X�F|�n���EU!�I�$ ��^���p��Kcڱp'���:�0�%i��M{1N����'Ǝ���?���9�ݓT�p�z�U"A��0ƍK%)"����O �"~�U�?K�6A׭�%-`Y�UA���M��,Q۴C����-�@�)�	`���b�2��	矌�I՟��	�@�	���I�|�¯�<>��Sa��G��l�U&\c�'0�}�$��n|dmH�¦�^�
���h�R�X('���'��S2�d��O[GW�l�����-0�4�?��Ȋ=�y��;�?�������y"�X�T��1�JP$j�J�֣RL�H"A�i;�,ԉU��9O�D��ߟ�^w��SݼS�[�P�FJb�Տ&V.�1M�'n4�D�OB�Hr`r����?9�����y�q" M��@��>����L��WMd�pB�\�ɯ�V����<� ]unz�-i$<O�9x�.\��Z�i��Ry���O���%�'��+Uv���k�5�I���?Q��4I����:f'\$��.�;�?��k�џT�	�^�x�����?���En�;��H�\ؑ����d�"%_/��s�4�yҢ��?I��r�8�O�B�'����˶S�D��)O6OX�Qԗb@�w5O�h`�'}��`�a���<y%'I��ٴ+y���"�#����u
��g�%hn�>{"�&�OJuq�'���?*F`�'�?I�p"�iQs��v���D��oAd-+�ieꁚ�>OF	x��nӰTo�?���!�?����j�+M�	Th,�ˈ�aL2$�$��Mc`aˈ��&D�>I��O�Ơ�|���?U���$p�ڣ�]�C��|����
�y���
h��`T�L�3YvP�S���M���?���?y\?�	Ɵ`��M�'.�,f �d��C��=aj����ן@�I����	�T���<�Ik"5*~�И�K�:�(� 0�Ц��	[y�'���'s��'^��T�0���n�g�����C�`�ڴ�?9���?���?����?A�������c�@� |��qK֎.&@���<�L����
��E�^ PP$	d@��L����'WB[� �'"�'��U�B�ϥ[_0i���Õr	����i\�X�D�']�'�"ԟ��r+�6v�ᱤ�Q.c�X�"Opi�L��B7�0��W��R"O���W�2{L<���k�]�!"O�X�F�f�ԥ �	:��(�"Oh0:BL��X ��jU��<g���1#"O�(��R$j&պVAM@g^%����X�	���Iџ�Rea 7���!1.Sx�&<yA�܆�M[��?q��?��?����?����?��&�G�a{���M�,y�1X�qM�F�'
��'6��'�R�'���'����Z���BՍ�c@��g8r6��O��D�O��d�O����O�$�OL�ĜySf�X�]��%�͢�(�l�ڟ�������\�����Iğ��	r�$�Ad��L��j�>θ���4�?A��?I���?����?I��?��j�%���ƣ��,i@��24Q�� �i9b�'
��'�B�'r�'V��'�ͣ�đ8��9 �#�]T�t���{ӊ���Or�$�O ��O���O����O�8��d��f�Kr��#P�Ir��ئ���͟��I��P�Iǟ$���X�I�h���<F�y�W*��t��h�9�M����?��?���?!���?���?��ܟW�b�z�$D	�q�W�\&1��F�'*R�'���'�R�'(r�'\��S�/p �`5선&�V��栕�y7m�O����O�D�O��$�O`��O��$�V5J�ⶣ�/�(|��ğ�0�Em�� ��ğ�����L��ퟸ�	����	5Wq|��%�)6kPDbu�&^I��ݴ����Oz�����dhD��6Bu*d�������)k�h����D��
��"�du��� E�g)!����x�e��ߦ��4�y�W�0�S�?��I�1o��"�k{�ȣD �ej��Ë�3B6H`�˂ߟ�Q�K��8�X%�0a�D����7O�U{p�S�^�QZ��^��f�!��'f��j�	��Ms��]R̓�� B�xv��[.����D�O�D�����<���i�,7-}���O��0����?bH�`�N(aN�I*O��!BҎ`�E���擺�.9�p
�<P�� �9�˳ ��z��MTy�V���	T��~��1	w����̧c!Ƚ�Ą۲�?Iq�i��q��O��%�i>����ߗKȮ���ʝ(	!�P"�^|�ܴ0�v�'�LL�G@������@\�1��聽�u�d��(M��h�
ʜQ[�0:�-���hO���<��d/ܟ-)��QEd�3[(2yC4�D>��٦B1�;��j��*�T��0�6I-R�Z � D�lL3-O��lڂ�M�'��>�ȁ��_�T8B`Ϋ_��V ��h��T��+.?i���5��=�ԋ]�hO*���>8� �e��8	tԘC��O~����+����)�����ܒ J?{��b%U�\h���O(��OP�O4�4\��ns�J��2�@P� ��wi|�A'kW�;�)Q녵	�w�V��o�7�LH��M���uoI���"���}Bl ��j0T�����O���<�+OQ?�!`ӨPX��r1*R�x�c %�d�]�V� ?	���'IV����Y\T3��˺r�*�'"��!�M���i��
Ԭ4��@�'%0ҥ-�u�^ 8�l�!� ҃Ć��e�����/�J���xⓟ�SRy�0O@ "�C�}�x�t�T�H��'��'<�7}&1O�.��qՁ?�y�P�A �}�'j�I��M���i��/�i��j��eNùc��Mr����i��Pƛ�N jwMۥ_b����0���E�^q��NLk≹/�P4g_1aVFa�dK�&�R(�.O����<�N~�'��7-�|X,9%H�5g�2��1��������\�	e����U�Ya������t,
"mN�M���k<�`����<���W5�����
<*\��'�89b�n��@1R�%�q�0H1�'��ןH��ٟ8�	���	U���l5��S�P	W���2噆\��F�y��'Sr�O��s�D��ʼ�e"P 8} l5�%kT�	�CM��M��iD���>i�'����$"Z�3���<	���>""4���
�s>������ �?��!
� �x ��������Of��˱f��e�Ǫ-U�94C�� �$�O��O�ʓe9�����yr�' R�T�46�D� c�nASE�p |�U�0��4J����Op�'mȽ��i]�[�L�qw�^�����ܟP��h�W���%�Fy��OZ�Uc�,Ra��@/��[ÀEHL͂ƈ�\x��'+��'�����<�b��Eՠ����Jn���DM؟�Xݴ7�X�)O���'�I�<�"a���4�0sJ	c��q��Vӟ(۴h���x���6	�	f��O<c��͖\��ԯ�:���`."�>��4���#���O:ʓ�?���?����?����pX7��l�0�Y�"�p	�� *O�qn�<*j��IП��	t�s��k
N =섬�0���ZC2�Bsy��n�\�m���?aJ|�'��l
�>&hJfL��d��y4��%P^���ֹ��d� 2ȼ����	琓O�˓d����ŅFӺ	�VcD�z�(x���?!��?���?�(O�Ul�^����y���9th��+H`����� �x��Iٟ��?Y+OT�m��M�'�'�n�:�d@<b9D���_(L�X� F)K0Γ�?���~�JL��T<����|���)���K��L��Ǐ�����O2�d�O>��O\�$"�'Y��{����3Ќmb�G\�SA>��I�����(�M�b*ZG~��'�������O;�q�"�����9�G_ݟ4�'�<6�ɦ���zP8d� �{����7;C�|Cv��5x"�`Wh�r���!�5Em,A�'��^�Iuy��'�r�'��o�c�=;UF?1���e��m�2�'J�	�M�]�<q���?�����$jO�b4�|@uFR5�����DȻ��Ĵ<�F�i��7��͟�%>%��9!$�Se˓bΤ�����r�����l@	��E_y��O��sb嘳1Of��𬄡If�H3ר�<�9��]���	cy����O�MnڿL'�y�A�F;IФ��M�@��ԅ;?9���?�M>I/O�`n��+83W���F��<cB◍� �c�4�?���ߜjNHϓ�?�g��a��H���o~�W�K� �b3C�W�Py0� �g��'��R�pF�A؂V�����\�O\��AC0�����'��n��w�0r�iD(������NqzX��C�H㦍�۴�y�P���?e�	X;�x�'w��H��F�P~F\`��_HaJH����ߟ���sA���D����7OްPF`ڱY�H�e��l�����'�	T�ɏ�MG ���"yb��ϗU��S�J:"x���������Ʀ��ܴ�y�W>i��G"NL�7E�?Ҿ��,�O8���$)\�8Jᮈ�F��I�?� 4��2�j��a����W�M8�
3��FS�D�'�R����^'Na�,Y&`��%�h�d�O��nڟ%� �?Q����|RV#��<�(Z��Q�'�	�ad��?�u�ip7��O�|�D܍��d�O\���`��D���Zw ������nR����~\�J>	-O���O��D�Ol���O�lZ6��yk��)Q"��,�fE�<�B�i�
�'��'m��X>�	�`��논a���a�`Q"sv]�'�7mE�A*����'�Z�'i���ѲNh)A���D��]*!�0Tx'� \y,Z�X[ �3!��	�'Y�	p�dM;� Њd��TO� ��������P����`�'�z7���A��3� t�С�?hGTq�嫙�I�u���'l��'��'b�ɟ�MK��iv���danTk��ֽ�|��u+�e��az�F5�yB�'�Ri�ďX9Xgb�iC[�T�׿#��Ot/�`��J��Y��D
f����������������ȟ�F���B�ɐ�a����)M"�?��?�`�i�"�[d^���IƟ��'ݴ ��
�9U�9��Y�&Y:ak��'�ɀ�M3ճi��/+;S����'�2���K[>[�쁽T��9�B����Qr@��9�LI��|bQ���I����ן�[�IեQ�� S��/u��M؀�۟x�Iyy�bgӸ�x���<���j�O$�4��*ѣU�ڡk�pc+OFʓɛ�
l�(���q���?���,Q��9����; } 2���D*�e�1� a�'t�����]^ʖ���=��#'T#y�x]#�c� ^�L����?���?�������$L��>�*RjE�`p@J �)�<����<1���'���M릀$ܨ����
��)S#�wn���b����w�m�D�O0X0U��%>Sx|���<!A���+O�DB�d��a��M��?�*O���O��$�O����O�'nz�Q�t%����*�r}�!����P��O<�$�Oғ����O��ɬT���AĦ��y	ǨS$G \o��M���'_�	�?i��?�2u̕�Ht�	�9 E�R��9?�̅i$�
��M�I�*M@}���әE��m&�t�'���'��� ����� A�[t�� �'R�'[�U��0ٴZObI���?A������ʌ�* <4 rm�]��� �R[��I޴JD�&��OP˧A�i��ٲVݺ�ʡl��C������xkUA�7q0 ���dy"�O&}c�����$A����Ĥ�4Th�Δi���'B�'�R��<�UZ�}�B���<hB����Fߟ\�޴�P� (O��d:�I�<���!a+1�á]u3�,[F+�՟1ݴJ�c}ӴIS`J/8���OF�ۇ"(٢�F�ŏ(���!0)L>	�>�Z�ɖ�8|��O:��?���?����?Y�=͂U*e�+MŐu8�	�M��S,O@�oډv�Le�	�4�	g�s�,��3p�L����̢ G	�6�X_y��rӖ�m��?�L|�����р[u[�QX4�M�F�&D2gӄB�T8J�M���Ϝ)L�h�e�M�fi�O�ʓE?�YI#
#c#�(�R!�1S�h����?Y��?y��?1)OD�lڻ)�0�	�Zגɨ���S�f�'.�5-r�	̟��	~�Oy��w�.�m&�?���3�hSTO�?Q&��@l͵EH�� �o����)�l��Q�2���'��$!��\*���="�2͚�`�*��%�'��'���'��'>��D��!�r�c��c�HL��e�O
���O�)m�	(��?i�y"�I.7jm���ye�"a�W��Y�4n/���O/�	cI��y��'?�0 �iC* ���(B,�>dk�͏1F�����!�ў���xyr4O���B�H0��y�1�̰k�(`���'��'�h6-�C_1O��	c>�Ci�4"�ȝ��j���PM;���<Q/O�HoZ��M�'e�O��T�\�z�0PH��z�ĳs�T�����.�,�ҍH�O:�	Ӫ. P���:�I-STd���-y��ٷF�00�˓�?Q.O���I��M4Ʃ4��e@ڣ|<����#���'+��' �'%�	8�MK���3N��X�M���YY1�-ϛ��'0��`X��y2�'X��1�8;&����O�{ \�x�V9*�Lԙ4��-4=�ON���<y��i+3�0�j0ቨ$ozP���""�7�o1Op��2���Or�7j�4�R��)2��3�@al�|o1�M��'����?E�����0IƋ�"�	��)�$��6:��<���<+�0�	8L�T��c�E]�>�G{�O�$�9���3��� ,�؀�Ƨ��xZBY�d&���۴��i�<�DK��x����í�Rdr��P�?�O>�(O`�nڭ�M��'���t�J�p����vab����u/0�$��4q�`��T��O���N>f�Z'%s�P��� �4����[?�X�*o�?���?���?q���v�Шw%�~~�HS!ㅴPQ�0���O�l�(i�`��'y���n����äo�ت���2X5��²��O��oZ)�M��i!��J�y��'#��Q�����U
P�A�e&�h#�`S�����+[�&+�'��ʟ<�	͟$����Ɇ'�]27Ȏ�~��� 7LO�-
0�'Ժ7�M9(x>���O>����H��<Ʉ�ƞ})��&m�7c�rd+ۛ����i;�4F������O���O]�Պ�4`���h��	��S
��V%�ri�I)0���z��Ԕ#E�	$���'%ktKV ɨa҉)~6�h�'���'���'��Z��ٴK�t�H�V�tt���\�p�:�3@[?g�}����?�����D�٦9��4�"�j� M�0=�9�B  �<�V���
��<1��/���d�i�jLC*O���@��1�&1��aa�Du��!���O��$�O����On�d�Ot"|�UC�P�nU�L�d�H��	����I��Hߴl���'���d�y����F<3�T��R�۶V� ��>�4�i(7M���S%
8x��O8Mp�JO4<�,X3@X� "������X�L�@
Ҁv�O���?���?Q��hꚵ���%bRJ�!���|~������?,O�ym��u]^�I� ���?�ΧH�0$22ㅾe\P5�׾]Fި�'���.�MS��i���$#�	�F���`�=^F�R#�]�A�EA�nHW�܋�d�.�(˓��Tk��Z���jO>��#��)��������}�
�2�Y��?���?����?�K~�.O�tl�\�? 򤣃`Lv���[�F�4T5!�;
�ş4��X�	Fy2�cӔE��:HŢ��I��=,5*%iO���I�4�vC���<��?�hZ��]:N���/O�4j剙/`��|[�kV73� u�%.�O���?	��?y���?�����	��'���c�H�~��1C%��G/�7͂81n���O�������<����y'�ć�@8)`���Q��E���3a6���r����k}"�O����O��5:�׋�y�o���ji�$k=�\��AE�%L���$bJ�����?�'H�ϟ���&{���+`/�6gP\PYA��OĦ%����`��ܟ`�'�J6��a,��d�O����aa�}R�m�v�����\>p�D;�D�<Ѱ�iӾ6�Ο��O��4!�Ȭf��H��Ν�q�.p����?IV*T�mf-��MV�����@0�0�ڷa<扏,ܔC�nG�N{�Ĩ�T="}4�D�OH�d�Or�$(ڧ�yr�ŕA���Q��@/�Bxࣃש�?�E�i*�Qz�O��$7���<��կXӐ��,"��Y�v��֟��ߴ)����O��0�,�y"�'��t:e�S�/]r�{u�R5x�`p�� �T��Ej��K@�'��IП�����	����	;I��J�<x(���FO�k<q�'Ƞ7��6Rz�D�OD����H��<��<:��1�^;z�9�h�\`�ʓJS��f�t���F���?��S�(	qCC�'��y9'��Nݡ0�5d�p�'p0��g�J L��xR�|rX��rv͌:	:}Z�ڻXj�$�p˗՟�������I��$�	}y�,r��y8�;O�A��	!b���5���IT��Ot�&�	my��s�H�lZ��?�Q��Ux� y�` �/�^%P�ˁO��@��`���	��d��MV(���'����������u�|z#�.+��d���'0��'*��'D��'=>�I4�A�Sj��悒����6h�O�$�OHYm�1bN�?q�y"HD���`�đ`�Q�([��]��ڴwÛ��OƑHC�M	�y��'#鉀��#FH]2u�E$Vq��Z���?%~�D�1S��'���@������Iʆ�ൣ L�,{#O!�����ß��'�6�,�ʓ�?9̟L�z�1b�p��K�+���*�^���'Yh7��Ц�����'���b�F��A3�*A���aW,օ/&��ɝ+�*YC/Ov���o���am0��5=].�`@M+�X�{1�Y�G�~���O��D�O�#�ɱ<A�i�.x�3��$~)�}*��{Py��B#=Q��ǟ��?�(Ot�mZ�_���M�l��G�4-0I��44��N�"!��'�򇆑i��|�ѡ@�?�ɐa ���	�P���H6bҍ6�<���Yy"�',B�'}��')?鐑焤Ѕ��	��3Xv�s�#�Ʀ���j������̟�&?�I͟�����Y�/͝p�*y��	m�F�q۴SϛV�O���J�'�����ؠyϓ3��c'L'U���;sG��;�>�a�h�t�r/]�0q�h�H>�*O:���O6�2@�U���l�FO�P��RR'�O���O���<�վi���O��d��qF��!�N;��@��EsK�⟈�'�n7�ʦ%�����+c�-��΃�/�P�f�&1��'�< ]�f|�)��T�T��U�j����<I1J_ s�p��uiPd����P�ß(������	՟�E��2O�T�AD϶"����C@�j4�)��'{�6�
�+��	Ɵ��?��'#��9��� Ǧ9���,F�p���S#�&�a�hn(��1dc��� MU��2��Ŀ�|{샀Ш���H�Oj�[�d�D��Ky2�'/�'B�'>���:1Ȝ!ƁW����w����M&����$�O��?=(���')�Jm��b��1���Fy��jӐmm���?!H|�������R�P4�a���Ρ���1 ]7$O|M��N9���� �`�`�f�i�*�Od�
�\�ɵ�˷w��$Hfi�pb�D����?��?y��?-O��n�1�&����I\��W�s,�P#ԅK$f:>������?I(O(�oZ�MC'�'2�y#
��<�V�B�4]$���(����?I�EK�'Y0HC�����n���	��QrQ	�pϚ53�KW�GG�d�O��D�O&���O���4§GK\�)7刌,H-�t��-r0� �Iݟ��	��M�Wn���Obc����X/��B�h
�9툅��ϟ��'��6�Kᦉ��`��芅�~���0�����P/x(L��V	\(��kE�Ї}���rэ^�'yBR�x̓	���4聎\����L��n:�y�IM�	��Ms1a_A̓���O?�����3[8HAP+=d;��+O��:�6�g��IV�S�?%!-����a�gk��8	z�	QJ�r��k4o�{�l�t(߸�l���y���!hB�%��lF�"bn�3쉊����O����g~Bu��IHa&;f�����s{�|3�j��)d��ɟ@�?A)O�MlZ�_|0@Q	�O@�h�3KH8a��T��4�?��Ä,uf�̓�?����'����G�P~�a_�j�AK�ĩ�虀�Gݝcy�'��W��G�Th�~�b1���T8U&m��|��֬�2ǘ'��ğ��'���z��t���P��1F(t�$)mӂ$m��<��O�����`��4c|
X�>O�v�`��qK�#ej\���O���
ɸ�h%ڤ�%��|��'����
�4[���8D`͜	�
�������0�$�*t�$扄Uu�QWaR!�$( �{����?(O�oZ��M��'���4�|H窆�V늰�v%
Ykh�d�O �i@NC#-d�g�����CP8P!�B�<a�FщO�
Mi"�?�]k�,������ş���䟔G�:O� �����d�D��đ$�VX+�' �6�ݨ7���?)��?O�Q�Wʐ�zh�3D��b�h���'e�7�I֦�Y�4e�1ؤ��<���>�Dh��l�b�{��FR-�-��H$�v)���_�����D�O��D�O���O4��En��*ÿ>�rTs@��;p_Z˓ߛ�Z'���'?ґ��'9���@�����L28<(��X��ܴ  ����O��|�i�Z]��HC�
`��cԣf�J�鐀[���RtG�<�ԧ�#��s0�ŝ����!#2���h�,8p�E[�f�~����OR��O��d�O(�]�-��B�")�!E�FS�%(P��� ��,W���'\�O��
�w�$��	�u�ѧ�#0���%�бg�5�c� ��O@;�)ЇUmm���<���<u��XB���'Y�)0�#Uf���?����?���?���?���
� ì��ɵ	��\�Yr ����?���~J��BѤX�	����<�+�{��Cu�c��c���?��O��nZ�M��'Lh$d¥� �<�9|�X�B]N���^�c����〃�C����E�	�䓙��O�$�O���y�}�&bU3}oʤZ�LH
c�d�O��<	�f��
���'mr�O��-R�"&��FO<�[����z��	{y��f�h�m��<�L|r�'�ɺ&F�0�<�
�	�p�'a�=
}��p� 0��D����@�E6O�@�O��gl�/&������<*��r���O~�D�O����OR��HʓI㛶��G��CQ�8pPI���3~��b�O��6��By��i��Ź����/��@��p{d�ՄΦ�
ܴt��4��-��<q�D�>hi�~�b�Q.Oh��'�s.�mW��Y\�����O�˓�?1��?y��?y�����5`"��e�?�T+�*I�x7M�����OJ�d��F��<9��yw@HK�0�gb�$\6v�2U�Z2N�M`�ʕ�	M}b�O���O�0���5�yɗ�+��ܡ

@�&u$O�-o�"J̍TP��7�R#@��'Q�⟘���Dd����%��9�8��u*h4�8�	Ο�I�p�'87M�3������`O�"FȈ �ªbM���#FUY���dOæ���4Y��W>�kp��(OT��@ J�Ţꖌ�O��N	$�p���i��F����R�C۹���*�'�t����4w@��)�cW�Xdj���?Q���?���h���I�_x��C�lJhGt฀�X�U������I�1�Ny�'�2�|�5O�䰄胘R�~�i�B1 ����'H�6����A�ܴbe���p%��<���
�|ٱc�>+S8Y1LH5�2�(Σ.�e0���������OX���O���O��	6:n�q@Γ��4�Tğ�^�z�%o������y��';����'9��叝?��tLX�M�t�S�T�ݴC��� �O������b���BZt���H�$�H@��^�s:"4�sB�<� !L�K	���ĉ����D��r�P'"߫�.P�R�U�/����O~���O����Oʓ2t����y"����DբO��C��1�C��H���'��O�˓5���!T$]�VF[�2JQ�'�.1����v�uC��+��y��'\h@���ԄF	��^������6NǬZ|�ћ���>)�P���Ɵ�������ǟx�	���F�DbT�l�t���1? P��CG�8�?����?y�i��� �OZ���O\�;���R/�/����.L�q�H�����D���Rݴ�2b�El]��Γ�?�w߄X��AhG� m��<�UŇD~�\Cë�u���M>Q+OD���O����OZ��ǯl=��#��0gq�h"cm�O��$�<y��iC�)d�':��'q��eB�i�D�;}��2��'Ls�������pٴQh2����O� �+�.ށ ����ޔ-�^�@-[`iY1�ۨ ��	�?�҆lJ5mt'���$I�}Ǡ�!���	n�Xՠwo�П���ɟ��Iߟ$?��'>�7�֙ �ʵS���M�d�2���tVН�T����	A����˦����7/tͳ7-H#?�1�s�E��M�ֵi���񍏱�y�'��Ј6�V���X2DS��/�=)fi� .� �X)�����ܗ'�"�'���'�\���94,I��B��[4I��)2��o��)�X��矄�	^�s���	�<ɆH S�z=�$`=(lI`PGV�M��iV �D�>�������!�H]���<� d0E<���7�p��p�(��?��S��ˇ9`.�$�0�'��'����t� 4o�5�GKBLt��'�r�'�bP�kݴC�:���?1�~���c�Oܢ�^�1�c�-{YX�`��_�0�ݴ&�����O�ʧ	Mn�E�^3�z����. m�IΟ�1c
�B�3!��Xy�O������v�$�&`��|Y��ɀCo��A�mJ0AJr�'�r�'���S�<��I_k�)�J��]���z�&�����4q�v�B,O���(���<�p��0D.��'o�@����O����)�4}��pӺ�0�n���D�O� �Ơ��5��Q���B�Y_Jm`$�
$i,��i�㰓O(˓�?	���?����?���wŨ2
�+UX(0"�HT�e)O �mFyd���ɟt�	j�s�l��[�'"�u�[S��1ze�_Dy�gz��	o�#�?�L|������+��K���x@K�gs�ܲc�ͅ1�\d1�����D��SH6�@�d\�O2˓PF�`�J	4 q*�K��55�u���?Q���?	���?Y.O2hnZ�s�]���3�^�X�b��b��#�o��o�,<��ϟ��?�)O~�o���Mk`�'���A%�4F��=B�m��aQ<�����5V�Γ�?��y��!��4�����M�]'$�D@��	�:�,���?U9��d�O��$�OZ�$�O��D9�g�?  pJQ�I�DW"d)E	W r�'w��'�6��hB�˓�?q�yrD�$S8l��.F�38�1��J�;F�S����4@ϛ�O�(%�J]�yb�'�Hk�eք~�8H��Z��J�
�댔�*�Mí*��'�I�t����,�I$&��4�؂T0H96N�R}Px�	ӟ�'~
7�����$�O���(�v�M+>c�UےH�J� �`^wy�]� �ٴ�����O����&�.���W�7����@
� !tnY�hb�Qv�<�����h(w��!��P���(s?����>
�v����?a��?���䧬�d�ϦA3�>ujhxy�Ȝ�G�*t��F^1�Z�'$��' �'*�	�7�Z���Ǎ99.9���Z��hF�iyܔ��40�6�{��<�#-�s�i��d׫!�r)���b ��"�6�ġךTm9�L��MSR�0����Iß�	ȟ��O1����4����L���i3�Qp�'R�'+��yr�' �d֘
��Y;���a⢁�V��+TF�7����y���������	�*�I��O�W���1�2�O;6�D�`�N��ZB��RE����@'R%���H>.O$���O�IѷO?Q&�G�~[uӆG�O����O$���<�ƽidDͱ�'���'����!���e��v���$�<���i�7����O�pr�%�)�� 8�˃1bDd�����?)��E�;&��D����$������p��G����&b���aroZ���O4���Oj�d;�'�y�!�g�dZ�!� j���A�Z�?�׻i�2��O0��>���<��c�1K^xl���.���
͏ǟ��4���k�4�bȦ�d�O�x��I�]0|j��/)���˖���>"�/T�5�R�O<��?����?���?)�S�� Y!
w�F�x`�	3Hߜ7U�P�ݴ[�9ϓ�?9��r(�󤄢CZ�\�s�*L�E��)q�� m�f�iӘ��	b�S�?��Ӳ �~PHcH�$�vuK��J5.J]HB�Ϛ6����'�\��gn������'���$]{^�P6��2S_��S��I�:/�U�IӟL��� ��ߟP�'��7F�_��d��,���S�"�~%���A]"�'��Ox�p����yӈ@�ɘ6�Nt�ԨU1=�y�ҁ]OJ�p�GχO����O���v�ֈ�Blx֨�<���"a7`�"&�2��$E�=^Fh�ɗ����?i���?����?q���?���D�/
|;�EÔ�j�#D�<j���'V"�bӸqc��P�	m�;���b�|0M��� �#��ѫ����d��Ar��?Q�f
�
}��	��D�c����1+��H\h`���1���ө��A�D%���'P��'���'�"݊��߻z���g`X�|�0��'��R�l�ݴ;�H�����?q�����I�:������^�r�V���W9(�Yy�{�СlZ��?�O|�'Q��%zp���?��#�	V�Kܲ��2�5�8���Z.��ퟸ5�dσ�8�ʓO�q�U虑@6���)~��.�O����O6���On��\ʓ���S�<P(U��W�U*�c��a%��f�Ty��'m�ODʓb��&i»T�L�����)�5)v�(��6��馁��k�iMp����;��ל'�V���XOy�OL�P�6�3�� �!!�c���
TrY���	ß����`�Iş4�O�i��x��e�7'%j�Y�i��36�'�B�'U��y"�'Q��(g�)ڰ����2��`
]�N�7���#���d�\�����!h�������uA64:WH�)U��C�l�/3���D�ڄ5c���f�@�O�˓�?y�	��Yk"�81��� 	ȗS��2��?����?�,O�oڵ}oN����8��1
��0��Ӱ�����3{�`�?-Oz�m��M5�'f員��AZC��$����	�3S.��O�1�E�T�X@梿<	�'Q�vSa��y£�	T��𑉏�p�����/�,�?���?���?����p���+�J{8 0�-�2��=����O�an9 ���'a���m���5,� V���5/	�+����U��Or�o���M�Ҿi�:IP4c-�y��'w�}Z��J�FPNE6嗅Z�P�g��"L
��C�;�'N�Ο$�I៬�	ǟ|��3D�2`���P�3��Bdо��'/�7ȵ����O ������<��_	H� �E҆mY^x������Ϧm�ٴ	�����OT����:�xI�ơ�3f
�Ɂe $uC4�Sv�	�E�����^1_�Lu$��'��8�fӓ$=��Ӧ� l��h�'h��'O��'��S��9޴d`�1�'���KF��^�n�A�#
�z�������?�\���ڴЛ���Oʑ���t8a�ǠJ).��Ӣ���,�L��'K��\���hsHD�tR���?!��h�M�jX.w��� ��� 	��䟄��ǟ,�	ܟ(��b�O#�  &�گr�� �� #��dc���?�̛�ս��$�O4b����`	�:,zԁ�E�
�8��b����'*�7���:;�T�Ad�<���qv��"��Q���hA#��٣k�=Cu�����`��}y"�'��'�`�V�õ��$��P�t%I�F�2�'��I��Mk��<A���?�ʟ�0�%�ڷU6�c��(8v�kUW��'6�6�FƦ-�����'��T��: ��%�7E8L�q.�^5�X��Uj&�(O�Iˎb1���r�-�d��1�h��A�	1&��;R��d����O���O���.���<a��i$�1�i�.XN�E)3�.#��D!qEb��I؟��?y+O.lm�6N��}X��K�/0T�I�j�7 �T���4!����V9rV��'n�� �>h��敿!�剁<�FX)�/!d|59�W9~�D��Uy��'�"�'L��'Wb�?� ^�( �d��I��:�X��q�l  �<O����O�����O��I�8GFEp�O�5e�`R ��O��n�8�M3#�'*�I�?I��?�s$����(��ԑp��R@v�S9y����I	�Ѝ3�b�9f1 t&���'���'{@�pu��0;J�4��/��@
��'���'��[�Xc�4P^��͓�?9��t��EA��Xd�f�.���������$\צ5��4Pb�Q>!�G	j��1����3-j��)�O�����#��!6����E肚,�x���'�v��gnܦS�hQU��8&MpI���?���?���h���Rz��@&ŊyL�෪�7|YP�D��a���D�O�㟐̓+3@h 
��]b�D�WX�����MCҵi��6��!ټU��5O��D�?���q�V�1 D��Ȉ�l�Z��տ	]]�$�5���<a���?����?A���?A����q).����#G�ʡzdl����DԦ��dGU㟰����t$?�I��\Lc���Q��M1Sk7_�m�'��7m���yk���'�b��S[�d�5�>%hR`R����ᡈ-H��)O0U��g�k�,�rSh)�$�<Q"	�A����8߶� �����?Y��?���?���������d�ߟ��-&J`�#���iP�X��I�����ß|&��'_n7���!���f���j᜿\Yx����B+^%I�ș�g4�Iɟ�(4�SL�ZF�ey�O���n��f���3�Ԗ��9b�nC_���'9��'�B�'���*l}S�Ü+Ch��C�8� �$�O,�D�¦i��@y�'�1O��b��!e>�=�4�C�G]nd�пB7ͼ>��i̦6-��TE���	����O��3aR|�r�1Ʈ�O��(�!/SJ{��Q�藟1��O�ʓ�?A��?��w�a#4F/v�:b#���I..!����?�-OR9lڜ	s���I�Ie�Ԧ�/�ƽXDk��yo������<ɥ�i6����&>����H�k،@4:Q3��/D�di �U�_��)	�oyR�OM�-�$dp��'OB�B�ܟ�HɊ���I��uIs�'���'���'��O�剡�M�[j(V�ˀ/�[ LX0��V�<�.O`�d ��oy¦p�,�Y�F&X%�`��@��5��*��Ǧ=��4@�-@�#�<������5�E^<XՀ)Od�"/�%��B�ֻ>��P��&�O�ʓ�?a��?���?i�����P�c����b$߾ <%���X23�L7M��tZ��$�O�������<9���ywf�89@V���
��Ȉ����.�&�d����	h}��O ���O���:@D��y"gɈ��TQ&��3N����	�A���J�J
u!'�Xz�'��ޟ��:L�(hk���98�\!���ju�}�	��<�I۟�'�Z7�U`����O.�D=Su��2��N�q���#DAǦuG>�Д'��7�V�U����Ʌ�B�,�8�DR�8W�Xj���o��'%$�r!�֛u/8-�^�d���o�&���FT�<��It��C�,50|`�"�۟������I��\E�47O�E`K�2�9����;��'�7m�ieDʓ�?Y����yR&Fn��Jw�U1B��3+U�?��i2F7�
̦u�"���31��Iʟ����T l;@C)��?m6�/D�pQ�(A�F�E�$��'��'���'3��'����Ǚ!zx�˃�L+$���0U� ��4lg|(i���?������<�S���@�>�
E%����W����$̦	[�4x4B����O��4�ʒZ�<�ق�]�J<����f�, �j�O�6B�I�Uz�`�q�?N~L�$�h�'(���R��Rq���4~ֈ��7�'z"�'<R�'��U�0ߴ:�|�k��,K�X�%��Sb���Ν$fM�)1��?�������1H�4rJ2�Ԭg�N�Ì�<��T+��L=��Õ��<	��sJ�,���Ʋd��K(O������I�m�;f�]p��6 �u�W�OD���O���O����O�#|
r+2��c��Ql	ґ��F�$�������4^�D��-O��d%�	*,ܼL��&��nw����A�#t�t���D}B{�̭o��?���J2���Bi)6A���ЁK��Rh���N�L$30-֫��H$�,�'B�'\R�'�.8�I�>��U:`EM_�4q#�'��Y��)�4u:2���?������	%f���2N����!��NQ�I{y�z�"�l���?O|"�'b��� ��0B\���Q2z B�;@*�ȑۇ���d矈�é��ax��O�asp-�b�,�v�ޙ<+f�����O8�d�O(���O����˓9���NG�5��H*�
ədq���#w*vhI�^�,��w����D�צ�`��\�[Oȝb0d�MZ!�Ĥ�*�M�f�i���!%�B�y��'�l���L�E�"�k%Z�,�P�ީi��Ai�[�oJP���E����'@�'��'B�'���f'.�S���uT4Xw9=vlmڷy�4x�I˟\���?Y��y�'�N�=p/�x
���>*�-��ƬR2L7��Ʀ�����D����IퟦH�rR�Y���ř1��U2e
�4��g��U����^%7���nI��+v�O���?��Pd�����x[*��Bn�&�����?!��?Y+O��l�-ܩ��۟X��Y�1��
(6LIw�ŕz��i�IS�IVy�Hz�P�lZ�?�/�L��V���g�pi��itia�㘥�?A�Y�$xa��+8ĬK*O���;n��8�Nd�<����:;�8����zr�Ó�O@�d�O����OԢ}��'p"�z����aD΍��z����iʛ�cVm��IϟT�?��'�z������jT�s$���c�K���Hy��m��卉��<I�%F��*p��/�0���kV#v92������Cۈ!�B������d�O��d�Oz�d�O&�7� P$2r��+!�0MA�K=[�	�Q����4`_�����?������<�󂑱N�(Q���!KbTI��D���D]ۦYy۴%h���OS�d/
*l�Q��F�0X
�C�	�+�v����Xou�I!$��Ȼ`Լy$��'�$3����-7f`�`̒�Hi����'���'�2�'�^��ݴyhށc�u*8aJ�z$h�$�4$]����?��Z�P1�4k@��o�O*��M�N�9��P&����,��4�'q�����'Ǳ4�:��'�$���~����Ǵ���#��X�����'�2�'t�'���'�>��̊�=�l�T ��Wd��
�O����O�IoZ8!CFi�'S2���'2�2�z�b�3N��Q�e��'���>)�i� 7���h�aU
g����O28���@4W\�\H�Ӳ˾�r��>N��A�I&��OJ��?����?1�����ݪ�Mȏ�J�:�����?+O^	n;h�^l��ٟ��Ig��i[�T���#˸a�,ɳ�W%��D�<���i��7m�ß%>���:L<����}~��%�@�A(X4R,�JKy��O�P��aG�'���)b���MS,Ԓ�(]�u��D��'�r�'���'*�O��	��M�f�0���"˲Ot�j�.\0�X�)O2�d�O�O.˓f�ƯԖ�r�!�`d� �ےzC����*x���l�2E���q����!���C��m�꥔'���4iD�e�����O��*ӌE R�'����X���P�	����	f���I�>t�akC4v�Jd+���x��&��O5��'�����'��<O�qYt����<Ҡ��!D���tӮ�m�?��O����h�	X�b[D��50O.l�d� |L�bIZ�4�� @���OtP7�Kh��`F�!���<q���?qG`�x�^q�r$�D6�\�#*�#�?���?����$P�	2�e���������n@���3mV�q� ��x����妵��4�RS>٪�O�g���f���7P:�$�O���ޞM;�9����E<B��2�D�L����'R|�a��s��(����6|ٛ���?y���?!���h�z�I:6���;��B4 <QXR�U&n�t��M�����#?����?aM>��'X�t7-_�8R2����[�� a�Q��fgc�JMmڷu����d�����)�t1%�*/ �h{�����LY��J�(IF<:Ua�f�	jy��'g��'�R�'�R�H=6%Bl�V��15��@��I��8&���M�w �<���?	H~Γ9X*����f^��e�՞C��x)O-mZ��M�4�';�O����O� �5F��	/v,7�^��@G�l<�ssU��x �H!\�Bq��ʍK�	ay���s׼q�T�������Dě$b�r�'�b�'}��'��	��M+�M��<�C���JE��N�eo� �#g���?����?QN>�)O�lڏ�M��'M��;6��!y�*��,�"N����# �����?��d�="P
V��!����=�;p���'wꞜ��d�(N
��O����O"���O��0§2�D�G��3"�H��iY%7x��؟��8�Mk�&�O~�'�1O�5��E'x��H
d��Fմ q���OZ�{G�6hbӔ�	�T�d��?O*�$�&�@�!TJ��0JuJv��4
=ᒣ�w�Hq�q�;���<���?���?���/
�<�jv'^�\�Dh��B��?����¦�腥7?����)��z�M;sOߣ_;�Q�`Lʱ
�I~ybhcӔ mZ�?�O|���-T�42��<�<4Ҥ�J�bp��Fe�3���	<��D��,�#$�-�6�O.-`�L�(^%��3qe�2�ȰC���OB���O~���O��� �q+��(��]H�3hG�1���#�����9��O ���OT�O�u���wq��2��(r�jd��eX�k��6�Ӧm�4dݔY��	�PqbnK�W�8}���Hy�f=P���H���"F�H{�W����ǟ���ӟ��I����O��	��ȞB�|�Ec�,H&Cs�i>���'�B�'T��yb�'R�Z�.x�����^��dz �2p�27�����$����)��xA�!��e���D�XQ�3ED7+�>�E�[��2��}�.�yL�O�˓�?A�ke���1loz<hgL\?s�bd{��?���?-Ot%n��7��	蟌�I�	>�H���:%��*���R�n@�?�)O$�mڪ�M�e�'��Ӵh�Bqzg$�6P���4�ҦSR��D�OTi���e!8|��°<��'O}@eѐ�ԋ�yr�@�eD���uj�J}��B���-�?a���?���?I���}��
�̭y��M��+C��zY[��O�\nZ�I�v��?��>O4qQ�Ԏg�I�1n�}�^�C`�'.�7��榉Bߴ0t�؂���<A�c�F���h�(�(:nF���#�+|��������O����O����O����#�XQ�A͖N$�ukp(N�M�`�({�f�[��y�'�����'��]���Ʈ�Y��Z?g~�yP�@��4}����O��.�	�F�·��EFX�r눰i��tN�;\��Q۶��<I""��!��!C'mю����Ur�܅q5�Y i[�|���zH2���O�d�O���O�˓<����y� <Vh��p`@J3	�$�HC�޴& ��'��|BV�h��4b�����O��
��ʰ5�M`S���h�E�'�� 9re�<y��:Z	���YgS&�h*O��)���:��LS@�3!ŋ�|��d�O��$�O����Of���O�#|���X��ԠHU��*�`�q'pyB�'�6�p���ɟ$�<���
	0�5�l�C+��)1��?��O,<o��M��'y���D��<���r 8)��Ϙ�&� 7��� p�q�&5�X�[b�������O���O|�� � � �⏙4S�L�V��	5��YA�'v�Q�<��4zZ6�+O��&:ЎM�I�V�A�@W�3vL���G�oy�W����4?c�vI�O���	T�yZl��Ca� �P1s 7L~�Q��*[6H`!�o�<�'~�H8�%@?���(��
��(I�D��gC�.ld���?!���?�������1��o�Yd�a�'`̄	�4���8(l�1�'��d�<A�i̮us�#��(hb5Z cZ�žP�mv�*`���u@EK4O��D $i�0�F5F=^��&���4��8�g_,UM�������D�O����Oj���O���<*s�H'Z�H�ʂ ��t�Z9�r�Ɵ�M�A�	�?���?9�'��9O ��h�-9���m��"e��Q�D�W��˦Y@ݴD2Y�\�S�?��ӜY�4�2�s�X3�eǱ �h�sr����h�۟�+�̄�	� 	7`�{�	hy��'<bKWF��T��V�&���F���rK2�'"�'9�I��M�q����d�O"�����K�d�C�M�hu� ��%%�IQyR�r��m�?I(�P�舾	�m	A�7/�U�F�'��M�$?�:��P	�V��I�?U����$c�Z�]-A&��#�2Y�}j�#��bm�i������	��I~�O��DS�%c4���.S(����C3�"Ew�нXA����IV��y�+#6�ʂ�$N��eҁi���?1�i-�7�妕*��_���IƟ�$��2li�T��|ܐ�ဒ�8`("�	̐dR�]�H>),O���OL���O<���Oְadh���D<��m�4=�\� ��<��i��Ü'�r�'+��yR%ƫ�v���K]�h�b�k�i�U�剿�M��i���d&�)��^�)T�FM�t����[cT�@͆+��4�G$Y&0&����H��h�g�`��M>�,On��7x3>��5��`��(��O���O����O(���<�i�d�љ'���]���!R��:Ҁ��F�,�?����'��	��M�i����r�I��d|:����hF.L�S��4�y��'�0a���*t�	
4Z�t�����['?�ry�`CE�w���(�ԟp���t�I�(�I�G��ň�BrQ���D�|�h��,9�?9��?���i���2�O��$&�I�tPb�"��B��`�0[�z�$��	l}""j�N�nZ�?a�j�E3��	��ꑪA�u.�T��ߪ ���r�� �x�IE�Ǥ��I'���'�R�'�B�'Ӕ(��H�^O�m��g��r����'��P���شK4EΓ�?����郩T�t━E�d�x�aD�Z-5G��EyB�s�Xm�8�?qI|
��]�"��#זV@۰��-��HB�)Z�S�L#���柬�c��P�4�O�T�'�"W^$h�F�A��ʶ�O^���O �d�Or�� ʓA����6Q���"�K;p���XfΆ�l,�O
��=��by��oӸ�1�'��i��tM�@C�1���Ȧ�ܴ*��"��<��>�&I�
�+N.�-O�z�����C��.�a[2��OZ��?��?���?�����)%r�tӦ�I�x��@�s�
��6�'�0���O���3�9O��Ds��X����.��U�R�
�83Q�Wզq�ٴJm�Q�����?Y�Ӊe �]bf}�p�q��
���Ży��\�H�ݟX�!�@�XL�������~y��'!RF�8+�����8���֬;>M��'R�'�剱�Mk�h��?����?�'��.�mن�� >��E˰n���?�I>�(O�)m��M��'��S7|�{R�@��m\�SOH<VbZ�d�O���P���K��<���>�2Q�6���yb�J�ꀂ���6
C�Ɖ���?����?���?����`����E��r�!@.fؠ́�.�O\�oZ�=�&�'W��$k�Ԛ�_&S�2�)���+`��jTI�Oz�o���M���i��:����y��')4x��kڇvDfًrŐ�UD���T8q�VQ U��/
�'���l��Ɵ��	��t�	�Šf
(f1>�����viB@�'��7��ezh���Or�$4�9O~D�3��3��mj$G�d%�<�d�<��i�>6m�ß@E���h�L(F�Ħj��� �Pd^8B��-\>�	�H��q*��$pU%�x�'TL\��摲$/n�I�����<QA�'��'�R�'��S�kٴZV���'������N�Wϊ�H�����?	�R]����4oțfG�O���H��4Ka�!m� 9�P!���/���O
0�K�(<c1X�&$�)�ߥ�#��-J�y ��E�w�dЫ'��O�d�O$���O��$�O�#|��JB�8
p4��B	~݊�ʑΟL�IП0 ݴQ~0�'C���9v��H0e�  �ePgK�,�ĭ>��i0$6���j���@}�I�G�b�����fC.$��ǔ=�p�o�,�[6�L�	Ny�'���'!�,U$}�%Hq�U�\���Ƈ�!#R�'c���M[�J ��?���?I˟d1��J��=׬Lz��0νA1[�d�'�7m���������O����E�؏X�f�"�^��pk�OA�w_p����R5��$��.�Pu ��Պ�O*hBw�,	(�a-J��P�Y5D�O@�d�O����Ot����@����­*��J��ÕE���a�K!4�.���_����~�����ܦ���"+�p�!�g)Ms�җ���MCt�ixĄ` ����֕�4=@�A'kM��p�NE��%�g &H*�� g"���ty2�'���'���'�R�?�B4�� _���Q�j��rWBpŌ3GDZ�?Q��?�M~��?��';��	�����C# �0���iC�7�_���'��O�Z��@N@��~� Z����ƅ.ܴa1���?!�A�>x	Ӡ�������O���'� �I˱�֚h"��cCb^9Zt�0�'���'tQ��ܴH�踱���?��_�\6�6g�\�;�+;T����"Q���4��VF�O�ʧQ���z�,L�h{�D`U��+�5�X��6�@��0���x�/F�(�����<A�'��y:v�uJ�J� 	�uDP��8�Iޟ���џ4G��9OnH䋔-ibxpp$�;@�z��'�7-G�I���?9�'����3#���P�F:P~~8��K��f�v�&�m�&g@6h�dd/?y�F^-(>���Aɂw��gJ�Jq����/�I�ޥ�J>�/O��$�O��d�O����O����m��&v���>&P��.�<	��i�q��'&��':��yҫɋ^�bt3,Q��:<�b�Ɗhx�� �MD�i�j��)�'Q �;��K'C���irF��K��� 
X<?��/OVy2��8U�� ��0�ļ<1��}{�A"�mߜB��%��I�!�?9��?)���?�������������<I�	ٕ*�CjX�J�xR��ߟD�I_����$L��yq�4>���t���rtDK􍒧��6SDxx�J	u~�LW�B�t�3��ջT��O��NA,Q5���
ڥr� I8�m�`B�'���'���'+b�S�f�@�c�U�Xxx���h�����O����Ϧ��$�W^y��'1O���VO\'e�(�����r�n y f�O��~:��dj���I
 �XXH��xc��-Z��q��'Wr��$�L#:5�����t���'���'�2�'���'v0xЗ呫V1��!nL�P�bA�Q�'G�R���ܴB�+*O���3*�Ȕ#b���a�1!���Q�hyRZ��r�40���O��?eIu��.���$L�E���`�@B�0��Y"#�J��P��z�Ϟ�(o0�N>i��=*��x�,J�!#jmీ^�?Q��?��?)I~�*O>0o���a@���15=\����_�i��5���FyB�'��O�˓fW��Ӄr�
x�3iZ�u�F!��Q�7���KPG�P���v,�H���$t��t�͟8MrF
O$�Bq�����-�,����'��I�����������8�	`���}�Zx��Mx�I�#^i ��l�/N�I蟨�:��y���$}�b����!2�����Ԕ>���|�4�Ia}ҝ�Ą�Y3��r�'��U��bV%?ZWB�S%`�@6n�O��أ̐���Pb;���<���?!���]�|9dH�2��BG%ߊ�?i��?������1:�H����I㟠
\zFx���$����p�E��⟀�'�t7�黎�����I�2�a4�X�c�P��<R��c�0m�$SU��$?�B�-���L�H(4!:��T�hKY+ �썊w��OD���ON���O��}r�'M��3gX�.�{�A��lqN���"S��ʅym�I��?��'��Q�Թ{&�-3&���b�.���UěvChӈ�l�>D��\�UO"?�7�S��
��`DJ�P��;��M�E��-Y!�dL>�-O���O����O����O�Ls����S�d]����L(e!1g�<At�i�t�rb�'���'���y��S�X���Aᬟ/9@��H�+!�剃�M�i�v��3ҧP�,�n�i�(�$���0��e�0�sl�<����$2���nY0����$��{���@/m�*���C�B�H�d�O����O����OD�؛����x�2�D�H�$X���b���OH��P�����?�-O��nZ"�M�f�'��X�`�yW�Y�k��"D�l
b	V��'y� �D�O�,m8 �������H#q&�;�t�9��(*�"�'fR�'���'B�'�>U+ ��U��Pe��B{�8 �b�O��$�O��lڃ3PĖ'��Ď!_���!Oҏi��`31�^6���d�>yp�i�"7M����E����);N��cEB\�O#�a�a�
�Es��u�c�4��dH�\�Fy"�'~��'8ң��b�ʕ��X�4A��<K���'����M�P����?��?Yʟ��$-�N}Ό����JzeR�W�̕'��7��A���OH꜐��ܠ*���O�`T����b[�ת��D�zĠ���*p8f�O~�a�߶2��Ƨܮ{��`�U��Oh���O�D�Oz���˓]�F������z`(�p�BP��K�x3�eyaX���	S���d^�a+
�q0�r��VX����b��MS �i��BS���Ć�oG��(d"��~���'U���1�υ]?"]�Q'P�|��d��Pyb�'���'\"�'��?�����X2X�S�ݢ�r�H7,E���%�러�I�H$?���L��h8�쉭��t��G <@BC�4mc�F�O����'�t��W?�A���&Y;2��t�<��E^����Y��|x)-	y�	KyR�'P"b��pNł���<�,Q�/{M��'���'��I��M3Vn��<����?���ŝC�F%���R�e��h���'��ɱ�M��i ��d�|z�̩A2�� �����X��2�¯�Dtq��}�#��lA����<p�ń\��+ �g0��p0mG�T�I���	ڟ\G�9Ob�d��h�VA���81H���'�7M�*`]����0�?i�'ͨ-Z�̨yvEQt�� �<�Q��%��6�g�&oZ$�|zF�>?yE�O�X��``��Т�p1a�U�������h��M>	+Oz���O��D�O����O0��ŋB�l@��{�L��`��<a �i�h�1�'�2�'3��y�Q�q�( 9���"½�� �Q,剫�M���i4��1ҧ|V<4�bCO=K�>i���ܕvkbS��%>2T r/O��i���6���Ѓ�2���<�� ��u
�'���Y2qʴ��'�R�'���'��Y�r�4G[&|�L�l1*T
�B�ytlװ<=�����?Q��V�<sܴt��O�O��X�i�l���0��8ry�%ǟt,2�(�O�(�n�*�:u2��4�I���ŪB`0U\�P@ŉ�89i��"�Od���ON���O$���Of"|�-��L����G�E��:�Hȟ���؟�Q�4�:��'aB�N2c�X�	#�+~L��ȘA���ĵ>ᢴi 6���\Q�
ѴW��I48�6�!$ʑ����k��������c��QH@_c��Py��'qB�'~b��dr��X�	�,*�r1F������'�剗�M;r���<q���?a˟؁���J�Q#�p��kr�|��V���'2�D���MA�'w�RU�t�ŗP=��jC`�7AN+�ΛT՚�b�� g� �'S�t�	|��łP�|bd�$z��x���{�r93`K̞6y��'��'�B���^��Y�4Q�J�K��ϖdX�DS�JNc"B��2�~~��'��O��ꛖ`�.F�rd�1*ǘK6��!�
��P��6m�Φm���#,2�[:����'�;\^��Οd-���}d�Ls0�Y�.�����'�̟t�Iڟ��	̟8�I}��M�����ŋ3?�|�g�S��vA@�y��'����'��9O@��1O�8X��"���r���+}�f�oZ��?�Oⓟ�$ �,C"vo��F&yo�,Q��J�$��]�`�#�2�ɂK�,܉Ѫ�o�'��۟��ɄR��p����E��e� ͗�v1��̟x���l�'	6�΢$��D�O����pc��@�2�t[E��%0W6�,�'�6��ʦu������W&2���Eƀa�\�X �
J}�C<ICŉ�2Hx�$?�Pg�3K(���W"fY'K��m`�jW��5��ߟ��	ɟL�	W�Oe����1F-�H�:&��"I�8�?�R�i��A�O��$+�	�<�w(�ejV��6OH�E`ܪ�O	ß��4p��FAg��-2�$��Cd�	
��!I��2X����)�zY[���T{�C'@A�IAyR�'vR�'(�'(�A��w�ԚB���,� �d��R�剓�M����<����?�K~Γ<�P�"O)X?
`�F� �Pv��/O��m���MS1�'�>�S���8x��,�A.�&i�@�D�)A��9��iQ��-�
]�ɻ�A9��<Y�K�(���s��^t,Q�F���?���?���?���DզIA������a��%K>LI���IR-:S��O�#��Cy�z��	o�#�?�kN*��mCw] ����r���.���rL1?�D�N>JB�-� �ҽ��'3 �J�G�*��D�sZ�M�����?q���?q��?����?��iܢz�����G�;�&@���*/k��'�"mf�����%�<	���'r]�l�dpV#�͐�P�Ƹ�2�'��	9�M��iV��o_�0���O��Q�D� ��`���ڨe�Ip��$H((��m�7
=z�O,��?���?��	�(�hS�#1&XJf$LO��hz��?)*OHn��˟�I�p�O]�]��� O>�!�5)T?MK�89)O �-/�v.g�`l��O��g]ĸK�Nɣ9ϖ�t�U��exV�G��� ���VKyR�O���	�$�3[F�'���J!����C�Iݖ!��I2�'[b�'���'A�O��ɞ�MS��ğ5��uI��X0pBUpR,�70�j�I+O���)�	zyjq�R��nٲC�t���ȯ4&�����֦%S޴f���#�+�V~ROٓU��$3-��&�Z=a���C�^ �p�Fj�T��<q���?����?���?i˟`�j���]E����X�2�dͨ�b�J8����OZ���O蓟�d�O���5l�,�c ���-\�q�`�n��M��'��	|�ӡ򆉸7.���3ܲ�sc[�G�,W����	�e�,��;|��m'�$�'���'�\����:l�Ja!`x�´ɥ�'���'��[��c�4��8���?�m\���U��n�@�`�7C�B�0��X��	ݴ��b�Oz˧�A�4e���e[ F�+
@��'"v4�&��़�r���@
�7�(��;O��[��@�SB�3�$F7���'��'�B�'��>�Γ?@8��S�+0�%Z�`�1C�	�	��M+qe����O|�(�'��$��'ק0I�%���*m�@�I�M�R�i�6�W�1*0�d��� o^�X�XC2c͈Sn��
�)ad��6�P�$��l'���'�2�'���'�r�'�ժ��pe�U�G���wyD9�R�|q�4b%����?9����<	�) '��銁'߀j��DK��)��$ǦU�ߴ���S^�Fi��h�>��(�ώ{lb�Rb�&j(\��'"�r�	R��5r��|�T�,�6K~�A��/Q�T��1H�� 䟘�IܟH�I˟<��qy�"q�:��g�q�<��GޚB��(ր=]�'a�O��$%��~y�lӎYlZ"�?!!� (fʈ)��n��T�FÎ'.�q�,7?I��_
=O@�1��1��'A%'jV�57�\(g`��[�Ъ���?Q��?I��?a���?9��i[�����/ 3Z`���E�XBr�'�"�e�.�2�<����'x)�Gg�Ppt�5kX:S�t���'u�ɘ�M3�i8�n��)i�O~B �j�푰e
2T�^��s�M�*�%;aEP:5]��A��'V$# ��?�S�1U�\�'`�P�(K�{�Z\��ٱJ\^�*F扴����'D�z0�U3�d��hx�8�A��t���F`]8Yt(j�䌾+@��Y�~P��V9���Z"��ur�n	�����m��/����!�X"m��0qQ]�h���� p0 �b�-;���3KP;�h��IiZ@��5�����)<OL�����\�����  e`�r�"O����,sf0{F)l^��0��b���gD�^r��b��O-p�h�`��=P.�Kd$#xv�4pC���"�҃�=A,��6e�(>&U�v��4DB�SCO�Y?�B��Q2b+�� �+*��9�`�"*%v�����:|f����6<jl�D��D {'혰G6*%�p$��a@���hr�����O�����@�'�����e��Q���-��z��?Y��nWXb���?����?Y�'���N�t��y ���>u�~$�D��$N��I\�>�oZƟ���П\��9��'������s36�Fg�	@� :��'>��e�'bR�'
��t�'7"�HA�`�p^�a07GG&L���д�h�����O��Y�m��>I��yR	�,H&���)�za�8��B��?9��?���Ol��1(���$�Oz���O"-#�͑\!��U,�6� SJ�O���$-˒e�>����Gh�)��̄,�� �O�2Վ����?a!�J�?������AW��G�nM޴)#�@�8�����b�Qs̚<�L#�F;���$?ْ!��ܟ<�I�@%����"ԫ�8�ÕmCP8��O�ԟ�	蟐��ş@%���Op��,x<���}��M"/�\���O��O��On��?擡O^xk�-�8���C��[�rB�	ȕr�*'o�b$�C ����ݠG�4�8rh�����f� <��޲7���gnJ�jU���SB�'o$��۰�'j��d�41l,R��դ;oX��hG�^=N�Y���FŠÉר"�\٢(�V����S$�]��Ğ;������eQ�>��$ ��2`�PCf
�2>7T4��ـ�Jq�g:�G؞H1��(n���)�ɓ�8�,�X�8\OTD���ϰ>H�z�%<���=~�wJ
r����'�X�q�Ǎ\�Reɧ��1p�����'$�ݸ�oQ1L�!g��r6���'����	F5w��E�!�w*���'�$�zE |ԂRW�{��P��'J=�ri@:,���R�}��M��';�u2�恜2�&���Ul^��{�'z��d���j�Ru���e����'����ᎾU[Z�12�Ԗ+��P �'w����ʙ(F�QWm��q��)
�'8D�sFN1ư�k�aӌ`O�ػ�'��Qu�L��z��5_��A��'{@,	aA	-X`��go�9]גM��'.
�8sd�t"��A薕��I�'9&E�fڊu�\��"V���Ĩ�'�6���dK�@Ք��W�.s�BP��'���;�!Ǖ=v�;�*Y�i7lEP�'�.�c�*j*~]s�ǵ[{`� �'}4*��^0�i�
<GK��'9�ixW&�q�f[�H�#��'��P��>xe�}@-�#��}r	�'r��AG@�!;(��@�4/�l�'��dd�{X�1�  %�����'l�K& SC;��Y"�ξ��u"�'������M�l�@1a�_�0	�'ͪ�[s`
�`'��W��%if��'�D�[pf�e��DӇ�
<�E��'������Ψ[��m��CKu*~M@�'{�P�Shۗ%m�����wBά�
�'�V�qWFY�����]�S16�
�'N�UB�Ț h�:Dhf�GMd�S�'�X���cF'FM�V�6N��R�'�$Ȓ�\�2��0�)��7�pt�
�'j�,���F���;�����A
�'���.9cJ1�IR�BV�A�'�v����L b����%źhh���'�t��F	N3��Ёc��<Ё��',���*4j^��#��.S"|�'��� i�)�,�q�ʔ5y��z�'0$�H��ӯ4�(�������
�'�(TؑGG<"�ڔ8�⁁y
�	H
�'��1���a]q��M;��	�'}�`���
�k��Zz�X	 ����MT4�J��� �$���Y'_�틑�� ^�lT"Oй�N̗Ew~1�'��<�����i<ԁႈ�g��|�O?7��I�X`* ��9_.YR碚�"U!�䀆,آ���H�%?��Q�W^�$ͤYA�8�a�������dK� �.�'�P)����;�a|��p����e�|�`���d8t�"�uFO7����J{(<�2��({i��Y��O�hڀ�d�,ʓA��ĳ���*a��y��/��]r �he�8;Lऻ$e�AӶC�	�2�.�r4h� x��8��Z�s�&	��C��h@ gو���D2�g?����" �2��6㶨:5"Ob�<ᰦH� ��M�� �7C�F�J�p���6HkI�s;� �ቒT,��f��>/�a����!g����dڦ~�^4*�l�Q&uZ�N��21�E�#i�V\2Q&� C��#Q2��$��
�R�C�k�6l΂���-YB8�X w	٥_��|z@Y"u7���ph(��KQ�<i!܀X�x��V�M�NC�E��h�5G�-��(�-k��T�d���PG��'߂�8g��O���󔄑�d��X�'��LҪ$�>�3�EJ'T�����.�
B�R<UQ�P���0<�2�ſ2�& yÁ�*ls��z��s����v�ܪS)�����|m��Z5��;�h� ��-]��T�FJn<����b]���r$Мdvp�"'�Rb�'�bEzt�aͪt�х�`�'�V�� �$QW�p���P$d�t�ȓ	A��_#M��D�]�W������3��I�ˎ@���)��<� E٠l��x��L=�~E
�H~�<�!�� ��-YE@V+*�ٰ��z?�'ɫ �P�xA�%�<Q� ��H��-*�a�!��`���uX�L��Aj��@tꇓFS$��L_�:z��A@��u�����85�*�㥭@	)o���c�Ci�����%|�Q>I�`�H�<����I,%����-D�؛�L��-_��q�ؘLި-Jq�+D�L�ӓ4�y6+u>���##D�|�RG@9{WV��vl)�d%)��%D��!FL��|(e�G��h�@=S� D��1�q��tɗ��z�R��!D����R*f�����$���Yk�
=D�L+!J�3V[�I��ԭi]�p���>D��K����nľ� ��[�$�C�>D�$��mX[\�}� �V�?r�<��<D� �5+��i���e��PΒ��5�9D��Y1�C%;�*��v�L�{����I7D�@X�FMOAv�!��
�9O�0R��1D���@�1#m
pb�;|D�X��j D�,s�^�l�4��&�ЭA��+&h*D�	�Tn�Q�!#� ���'D��Pt�N'0м�e.ͰQ�����O"D�,����8�>��ዱ?$�;r>D����Å�C|ƅI8V��ܚ�e>D�������J��l1�A8�D;�J6D��:�,�(���$%��-L�{5(D��!�'��ls�C8n�$��%(D�8��,��Di��IU��F]��"c5D�੢�3qz��3�؀U����0D�x�2��,�y�gΖ;A\�#��1D�d֬�=QHh��f`�M�<�C�C.D��J�oU2Q��F�V0�5���!D�t"�#�/l�8$���\Y�̳dd<D�PׅO%kv(I�Ҍ�ظr�=D�h�*)9L ����`��'D���<o�°3��R<&Rp��o>D��#���2�p��Z�ą���:D���s��|�����1҂�94&6D�$��Ə�dP�uqDW?R�a���7D��JРK��J�2�4�Fe3D�<P�
�{���JլS�L\8(K�e1D�� (`3G	�'
�	�(A�kX	!#"O2��1"D4r�p�f
lLy)#"O����c��S���h�Ǝ�V�:P�7"O���t-��5npI��\�(�
��B"O>Ua�lѽ�,���!U:0`�-�$"O��0CR�_�ȨI"�_�R�A�"Ozq���v��p��oR T����"O&�`N�;�����&C�8���"O&`q�܌3IؽB�.ҿC�4h�W"O.RC��S��i��h��H�D��h�<1�B������A�4AO2����a�<1bN^:�������!>�`��b�<A��:�j�*��ˉ ������A�<���~f���BT-1�n(
Q�C�<�Ķc��	� E*I�V���'Jw�<i�A�+u���&�Ҫ>1�1StJ]F�<a�Q�F�� 3�8c�F�:�G�<酁
S�,�ʄ�`yĒ5�}�<1�bEa�x�c�V�8`@2�,�~�<��\�2^�`�Ph�70�`��u�<9�l~^�U;s��)3���1�%�{�<!��Ǥ\�Tq��J >x��C�o�<�A��9��P#wn\�.�QY瀉f�<��� 6��$r@�_3�iI�`�<9Ĉn �@�=ZHy"����z!��X�S��m��C�0�@����[�!���4<e┫ť�#mg�����-!�!�$� {�i�ĈH!}~��R�V�!���}Fh�r��.~j��H��Ɗ!��H�o�褥Geb��[6㊭5�!��U(^>�V.	�Ao��Q"�W�!�d393������x�䁁:w!�Y�<Р�g�D�A(��d��|�!��.]�}��$.}/��
하9�!�d߂@�����ք"�J��U�!�$�l�m��E�(�ސ���-�!�D�"g0@��.�	e �R��U�g!�_7-̶��S�/B�=C悑-f�!���3+Rf5��n	�I/D6��!�÷Iq���bV�N�ĺ��t�!�ą1g<B(�@�*j���!���AP㟢}J!m2|���z�j�m~�Hd�Nj�<���[4H�5(w�j�ua��Xf~rNާ2��뉅~���7fx�D�I�|G���D��&�8�sfF*`*�&�G>�p� �]�6�!�dH�99���� +ݎ}��C�t?�1��ƱqQ>]���\+�!��(5���k�' D��B��"��a��*^$�b6kt� R�O�u,qO?�t�6(�e���^A` azu�)D�\x���J!ܔ ȝ�����*?9�P�(���$�F�P�pAe��\�:,hS��-X�~�%Q�����P}�4�&��0J04@�0n��y��PZ`�1bUb�>�D$𰋘+�y�&��aT���c�<KD�맨T��y�$�[���Y�Ks~�x"�F��y�MԹ+5|���Q�ޘQB-��y��_�l�)� By;�d�1�T"�yr�L�zކ�ac�֒;T"�"����y��0c��۱��+a�x�'A,�yC����PY0/��Otqw��y�b�/)���3�N6;�@���yr�l1~�d!���%[���:�y¦T�;e��ˀ+�6}E��ulF��y"�K�g���y`^*8k�����]�y
� ��[�Ȏ�I�|�x��Ӄ��ɺ�"O�؃f�7T@M��U�`� ��r"O������-bYE�,+p��:g"Of�"HH�7��͡�S�*���:�"O���G�c����3f���&���"O�]�NF�$�T� oB1Qh�*�"O�d@��t�T��( NU�@�6"O
�S�.P9;�x�0D�R�PAC�"Oh܂"Þ=\�����m �w�d�1"Obm��˰+�&����E$?B����"Ox��B���7~�H�"+�Vu�s"O@�h�a�%B�D5u��4�T
_�<A׈!e�`თ��12��h� �U�<�C��X�<Aq��H�\����n�<)���7�����Ӣp�� �Hi�<Y aQ�A"H1��H�5���H��y�+]"5��A�BbY�;�=Un/�ybA��g�����1�:�St
�'�y�dJ�C R��5���{qH9S'��y�ؑ
t���R�E6t���@Џ�y��$y0�!�Fv+BM���� �yb�-���r����i���!����y2)߰��A���Œ=�� C��y�d��� &u>А�L�8�y��I�;���Zъ�n��$��	דq,�Q:��S3�zX�O�Z�:d�sM��=�Ȉ�q���B�	��nq:@/V�1�̱� ���jIVB�I\>�M:�#�J"l���v�BB�ɨw���i��)�4�p��U�D.B��)N'�9�5���$�9��Ӟ�C�"7ƽ�c����n��1���!"O��{�O+3R�sH�0�����"O��z��I�dj�+ǴJy�Mp"O�H����C�~�G��f����"O���e���<kTIy�&�Q�<���"Oȩ�uD�/.鮹�hَ���c�"O��X\�Z0�,�$��!��%{�"O+���!d*�����a�A�4GL`�<ٗ�5r��Y�G�#Q8��)��\�<����	!��K"���E�Uo_�<'�ٱ~��$��,L6;����Y�<��	+]���9��X��lYa�XU�<A$�ڑ$�J㰁]��P�N�<��\K� &��,$��r�GO�<)�~��}��%�� �����Y@�<��&H��8�&OKn�L��e�{�<I��,t�xIs#MF>.�Q��x�<�PL߁Nh�����l�v��a�Is�<�AΞ�l�W��E8�90��l�<	���H~ɓ��ޘ�
�y�h�<A��%h������A&�|�Đc�<�3g�/y��(jw���Dm��g\�<�G�J�c^�=K7O��}�.a�­]�<�i �I˒�[�
h�4$g�S�<�� �-n.�P���.X����Rj�Z�<����$���
��*Q��X�mDU�<�C/�	D�H=Y��K�5��h�j�<F圛_�m��	U95�(*��Qg�<���`�d����0,�Q	�b
d�<ᦉǱ(k�͓d�ӂ���1��D�<���DH��}SU������`qn��<���!}󚁓1�PcI,���"r�<��.J��PK��(��9@�Tg�<�kB-+�<�P��I�P��)�v�e�<� 6@jV�h2������8�B"OxT�U@�,D��{�H���"OV1�N�ntܽa�"\���v"O�����WE��d��Q>f�%�I}L��G���5W$��)����h9�@��yrDO3 x�(�6΄�l.�r�i*�y�˕#���=E�t�81��h��#|dSs�ű�y2�B�F�R�� %ڻl_T�.�+���6H^d�Ԭ����<) Bj�$�@"�N6� I�u"v8�� "iϹ0�A��+�Ctd11J�qZd�Sf�!�ɇēcv�p��Xyc�ԫ��ٻ:��-Fy�Dǒ���s��@+���!���7J�����P�7ߠi��"O�}�v����q�6I���i{v#�'�*	��S�)֧����H�
�RT��M� zhF�u#C*!��׀880�zrL�L�~��CA�T���Ga�r��\�}��	�/�����Aմ9�8� �D��n:>���[: ��� ��O5��'�M�-^�X�����8�������x2��a>5�w䇴͎������'|B�gK>�}iV�0�S�	m��Qǃ��Ox�qk�
X5��C�	�Vy5z ��~�*��
7�N i�I�c�Zm��؟�~r��R�(P�jE� �ÂA|�m&A9D���s�ͦ8>�1�2�@�|: ;3	�OZm���Iۘȡ��Ӱ<y@�ZF��8��((�Y���k��C��?O6ؼ�N�t�|x�!=x�Ba���4-�neH	�'L�5(��njt	`
�3i�R�9��$ݯ3�4+����c?MP�n�^��d����/|;�@9��1D�$P7���x)W�Q�Cl�ȸF�O��ע����T:*O?�D{�AP��9[Ρ�s��!�!��v�.hr��U/v�F���	�3���;?n���2�G.��y�'$d�lM"�	�:py�����0?�S�B�_� �W
 kP֜z�%6�JY�[h�<i�ޑV\V��u�Q�J���"�P}�'/`j��S:C�Dh��8ɮ�(3�F�&�C�I�!��*�ID�}x� !��iu�C�	�
���Y�,RO\�:���yC�B�I�:vD��S���?�!iR��.(K�B䉛8��I�(~� Ă�$<�B�	3N���s&	7�&��ٙ2C�I�}$J9@�� ^����-�dC�	2���1E�T��2�W��B��4� �"�!\�;56�FV�=$B�Z,��3ꛬG�Ф�Wk!]��C�6m���S�	�)
Ĵ�Ɗ��G(B��@����xqd�rc	�7`yB�I�*"�����E��J��̭Q�C��]���Q�kԖq2�������C�Ƀg �#D�2{fN��W/=�C�I�[�l�{v �.o"`F٦ ��B�I�kx�s���#�D�2�w�B�I�9u�`r�H\W,��$���mĐB��&h���0 ��6�F�4A,$�tB�	�	굋�3b�*H�V��r7�B�	 �F�5k��$ޱH7�Z%U��B�IM~՛��~g����-$@�B䉚9�튠�S�i�9b0⛃КB�I���4AReN;K=]K �W��B�E�P�A'�p0Bh�T�҅"`B�	A=@ۀ͔9hR�!�+N3>4$B�	�8���4�ŧ�Ɗ�igZ���"O�`���82M���M1Z�$Q�"O�ْ�#�:=�v`(��Y2}7V�@A"Oj�z6�ʽ$R sA�[�E#��F"O�)�4@*k
�ٓ��X
���g"O`�1���-w�Ly��Θgg�1U"O� ^tyŮ��>a��ƀ�v��l6D���ש_�K2*��$�
:)"}��F#D�(�A�D����J�IJ�d�7�%D�(��[��ܢ @K0����c&D�${t��U"  �K�$p��`��7D��k�ܞ@r��SF�1QD�C�"D��������Ad���6`
pn"D����ĸ=f��9p�1C	n�R@<D��(ҥU)d�j0�7ic�]Z��8D���7L�| p�0E�2q8N,Q$:D�Kb��e�P1��Y:g�
+D�t��'5� l`�cV� �����.D��:W�����i��ı`�i+D��Y`�L�FY��Է\씅�Q�'D��d�S�*i ��JZ`;qB+D�:P�O��z�i�*�z͓Ӌ;D��I��*k��l�qjBXA�G�#D����&K�Њ�/�=/�J]�� D�����b5�<)�@0�N�#�K?D��x`bL�S3<<sə!IZL�caM>D�dq5A�1lV��'J
.���:D� @5ș�p��Es�<�Jly��6D� c��76L4��Ϙ"oC�y�7�8D�ؓ�dΆQ邙be�
?�����M)D�Tq��
�fqYf䒨+nQ��a%D�|�VƘ?G*�]��fF'v~Bq�g>D�x�vI�(A����c����a�?D����Z�%1�l
$f�\v�4qn<D���9�TSG5���Q(-D�@��i�<H�J���EZ�ʔ�!�+D��z� m���v���?|��@�%&D�4����?���S!L˥[OD��G D�x�4 �Fȋ  \4i�5�=D�4a����b��)3����L�25Y�N;D��Yb�� ��Ñ,��f���V�,D���G��?��QƏ;q^�|�o=D��AE�P� PR�]zq�0`S�.D�P#�"�H�<)J�B/m�ȌA��,D�D���_'�@XSBZAݼd�An+D��Hq(
�K�5� �ҋ�b�g�)D�hrC@VdgP�"���.U�4M�w�(D��"�^SO
��sJXdO6%P�-#D�����W��"o�1JE����3D�ԩ�d��"���"�Z?o��*��-D���O�,i�ԥ ��Lu�h��0�-D��E� [C
1h�	,ΜP��`!D��pF�I�a�8��5�Ȍ^,�2D���w�ӗ@�\u��P�+D��"1D��z��("w� �iӄ<`�� .D� �Æ�/�d�Y��ְ<y��'D�L�b @40ޤ ��Q�bn��iT�&D�pr�?3\L(�d�*��1��H"D��C� ��@�P�(���aB�Eq� D�t�bOP��af��!-�HY��#D���r�W�'-����V�(e�V%<D�0��;TAz�(mڱ[e�<�a8D�����
�hI3=[�yj�(6D��;�<[X����lŨw�t[v(4D�\p�c=X��a� 0o�k��0D���O[�5(���6q'��P�*0D�pA6#'z���kC��D'�}q��9D��Ҷ���Z&����X! �؂�2D���eO��"uP�� �NS0D�D�!��!U��Kׇ�e�v8�3�.D�� �,�4�دimT��dO�Z���R"O���ˌ6)ah@KbO^�7ȵ�"OP��N\�-V�9��Y�r�"O����3ެ�AJ^�:���"O~���(��}* m����>%���T"ON� ����\8d	��Ɩq0��"O���c��fcDiyq�kj8L��"O|�Ё�z:B�i���h;��"O�5ijF0|��n$+��j "ON�!`���"��y��#�!����"O.}Qu�@:��ʴ�;��Bs"O�%�&jN+��<��������"O�Z�G�N�P�:o��}�V"O|5�Ed|��i�K9n�*�"O,�H�(�*xF4��e���{eHp�"OL�W5?ͬ��B��W���"O|	��mO2%SPD8���0Wqd3'"O�����>x�@lpi�iXI�"O�A�gY�1,,�4��e �a"OX5s�<4����"�� J��I�"OD�	�M?8�� ��VW�^��"Oإ�$�C�M@�Y��� n�v��"O0�xq���b�&DKt) "eu �b�"OFT�����M�|`�`�7?k�*�"O\�!�N�.>Z �j �oOڙÆ"O����3*��Py�J��#�R��R"Oxѕ���(���p��Z>�,yѴ"O�ԣ5����0
���\kʄP�"O��+W���!�L%�7Ζ3@ZD@J�"O:Hk�FVh8RA�҃V/tK��h%"O�Iz',�5I�lh�B������"O����!Q<1~��� 1_z�*�"O��c�Q�a����	Topz�"O"�����2r�aGc]�VX�U�"O��@��FP1� @��	�"O��P���l�.����U"v��x�"OP�R���#jIn(sD��/\ۊ���"O�XБM�+>V�ٲD�)���e"OM���ή꾤����X*&"O��Z�-MdEn�3�@ժ2Ll�b"O����l�>I�~���4�}r�"OX�A7��>�q`�䈛z�����"OTԢ`뉆R��=��N)s2RJ�"Or���S�j\X��Q�$>�H$"O�xR��R_��b���D H@�"O *�Й&J	"��	�Xz"O$��1
������Dΐ2$H���"O��V�N?�ܘ�g�G	@�b��"Ox��G� X=
A(J^;B�rp��"O(T��'Фb��h0)���ꭰ�"O���2�
�~���D҉ޮ��U"O&t�2+I7R~R���N�j���b"OL�i��SiPάC���z��d@d"O⥣q%�0B�j�%�T��re"O��P���q	<y�x9p"O�A@ �U}D"��O�]4��"O�թ�C��5$��$��,� �"Ox<�0ǏA��,��*�p����"O�#�B	-ۆ!�1R�1"O��hxR*�ڒ��lb�B�"O��ɐ�R������ �6��U��"O2�@�&D�w�|��.�oѬ���"O"�hS��	@��AvG�0_�RE9'"Or!�W��ST�p���Q��k�"O� �fa^3���d����"O:���%����[�(ys�"O�(�s�_v�Ȋވ|4�53��=D��w �ZB@���9���k��'D����L
5�8�B�f"�v�{f�9D�x��h!W>(�{�iݧ�Tm��$2D�� V RZ&T��/W'#lB9S�./D��BE��?3h$��K��;�Z��U!0D�t(ԃ\0D<� ��@�.�0�"ť*D�� �4I`�Pȓ��0	(.��2�,D��1�DX�u�"���3�: ��>D����ծ.�����a#HXӪ<D���`Q*T/��cTi�Vǰ)G&D���4kSV��a�ܞ|%j�qE�#D��bb���P����ءo�,�I$D�PC�l\7l���+�"��%D�08!N�o��8�&DUf���A�.D��G�$v��A���-*Qx��*D��'�=z�$���B#6��9��)D��ئ���� GA�E�d�'D�$"��L6~��I�AB�3|�L�r��:D��{RG��0)`LPe*�6)I��9�������+�`l�����!��C�"O�����G�l�� 3�I>p4�"O���R���p��2 ���J�B�"O��X#Ê�,���)/R�F�N�ʇ"OĀzQc �� ��'p����"OR ��ϝ0�L5a����}�x�V"O�3�� �pm"x��������b"Od��%D
b|�����`E�"O�@҃��/*�H"5a� ]��ke"O�X*�I�#q E�!+O%���K�"O�󈁚49P���o�5rց �"O�<���	h#�Y��DR!"O���G���;�\	��a�(�:1�"OR=IT�.;Ol�2���q����"O���d�שl(�H@�� g>�r!"O-�C�]//�Vx���+Nx�"O�9h��F�}C�hxƨ5`i�5"O� PF/g���Wen�=��"OPؕ8F�D�q e+WP 
d"O6���l��A"�!g�
16ؼ�8�"O"��7�V�	j�(
�ܾpgV�A4"O��3�kD�":�ݲ "�8¸��"O�LCb@�SȔQa�%.&�`�"O`����8>�:{& ��M�\�G"Oz�z�	!f�ޭ8p�tr�"O�੗k�?	��k4�غ�i��"O6M@S':-l�i���xU�,�"O�t�Ĩ �JUH��U�[pI��m(D���獱J�p��������C�,D��Sm7g�t!�OBg p���&D�`
P���d HM���K�w&d��&8D�� �l](��y赋
�ܦ�i�n4D�8{�A�Bd�)�fH+3ܵ�u'4D������ &�	g�X�.�䙘5e3D����s���j�B��~% ��O3D��(�`�!#�:H#f��ct,�[W&0D�p�2aS8d��k$�R�'{�s�h.D�H���Q�d?�%I�#�J�e�3h,D����	|����Q�"eʍ�7�)D� �2n�?���/�z�EK�.:D�`���#?�~y�e��:<V��d(:D����I�	 ��{��9z�zY�E�<D�� &D�W���x1A��& �"O���E ̮H���P��R�"O��;���7Y֘ur����@*%"O�H�g6c��J3ꞽ:�D  "O8�W�M��,��`�TLv4hC"O�03A�O�JVr����\�|`f���"O�!a$¥[*�$Q� �7Ga2�"O<@A�ҁ��5��i�Q�-�T"OrMs����1��H��.�R$"O���R�fr�1����sBYS"O�e�e�@&��@���E�]�
�"O��@5!ێ��掑�i$h<;Q"O�u���=w�����h/TY��"O�%: �Q13y������p���'5N�����)}����K˷u����'�}�r�Ps���Y�L"}5�1�'����$Y��lsgd�phf ��'��E����s�J�EB�j&��1�'���Y0,S"X��_+VX��'e�+���!&Y����5V/2�K�'zL��$ݷg�$a��RL0��'��i0��Bl~��Ɍ�I��z�'���C!kC�<x�@�E;Do�l��'��wk�|w&�2�D�;��@�'Ġ��!�I������� u�'�r���./�ZuC�X�v��1	�'�|(C�`�g���h�.�o_P�B�'Cޥ��L�T�!y��2vSp-��'$�=[S�Vv��P�&]�d�@�'cTu��N	m����M�/#G�&;D��`�7?�̍Rd I�Y�,pi�H7D� 3�� �
����ȴc����"D�ț��X$5�
��q�t�!D�$��+��R� �t�O] ����;D��v�sH�����k��'D���Rj'͕�aW<�搫�f��yri�${@������v���0�) ��yr���f� X�F޹�uk�kX4�y�F�e���3)̼Z��x�B��y�B(�N˱�C/�~$����y�,>(@�aQD
�}��[7!ϫ�y�랠q&��'�Zud]��֫�y��T�*�y*��ȜX��ׁ�y�o�)F5(\B���(��Q�o�
ػ�'q�U���ߕQBeː)\�;qP|��'ɬ�%*ó.$�8�e�/	�E�'�ԉI�Ĭ�6�+��C�$L���'At-����X�Pغ�/Ct�@�;�'-����,="Y��'	6��ȓR�PQh�U��P	 "�-V�X��+�N�jEO��{(�gë�t��U��\��A�*�?QL"��ȓY(T]�7�ؕR�čku�߽+\�D��8��Ks�8��x{Ո�	<��ȓo��1��M�W���* ���B�L��BV��#��~�����gA8j��$�ȓ�5� ��
JW� �� �2~��ą�"�U�e�L�OH����
�v�B�ȓ�l�jb�Tn��P�����I�ȓ��|�M�Y�� �b	�(�^���1�����+�>K�f�upC �������C��X�`
�?CD��ȓD�|�Y�K��^��ς��h���IH�����@�!�08cr
Ԣ����S�? v�6��f�P�A����6��"O8��Ð0{������5ЬEJ�"O��#�#�3��ʔk�����"Oq��&Y#:���sȆ��\�� "O`�a�%v����-4�"O~x���̘B�)9�眆qn��Y�"O�Z4C�#�1�ڠn�
��$"O�4�`�&�ds���k��!�"O��z�OČgj(�	@����"O>�BCO&x�0c�ÉlBR�"O�Q��#4���5eL 3���"OH�S���Q����e���iw� *�"O�� !�6y1VA��C�_d�- �"OD�3bq[�#��B]�9��"O����@f�i(G��1:��rP"O�I��X|����1 �r�G"O�(ٓ#۳n7�;�P��h�"O�y*QaEK5�:�Z��"Oc%*��1Hj�0�/ĭ�|���"Ol sa�'�����Ӽ��Z�"Od���UX�TD���Q/�\yF"O�� �L�*�\@h��67��<�E"O�cJ�P��5Aҡ3:��i��"O���Ӂ�GP^���&+M8Z�"O����K�{jl�"W���f��<
w"O~D�%
J�lD��M�&S��<8�"O�����F�[��AV���H���u"O$�`iN<(j|YS��*�%AC"O��q����D�	睓&�(�P�"O腑
�5�4p@��&�x�""O�5�V��1$� ��m��X�BP��"O� їD�?Ø �eϚ�v-�l[�"O>Uɲ�Ǳ"�l���nS6{(J�y"O�er�e ����KƗ8����"OP�ȶ�Zx���rI�~?�x"Oذ(v���X"���߇w��"O6U�u��-0=��Z���<bl�ɳ�"O"�)�@�8��0�7n�>Q*@s"O�⦢ϕ(��ȱ��֩_3��v"OX��'��~��͸�iQQ"TT"O��b6��weh-뷇q<f��"O*`��s�F1�&�m<X؊"O��	b -7�~`�"FÙ6�9�"O 4�w�_�$���#H49;
��e"O�ᣒĒ>��!PugٽN�ģ7"O^]���0o������u�n�`Q"O $	��4��	�Ջ�#���W"O���$ �	X"����k(+�2rs"O~�2�O=l	�� ��;��8�"OV��"T�T4`)Eq��uA�"O�s���dϒ�B7) �\>I��"O����e�,&� ��(F�k��]2r"O����-8c�5��j�7�`�r�"Oxh+��#{"�8@��)>��t�<Q�Q)?�n܁C��h�D��Q�<�Ak\�"fJ�Xqa��3��[7�K�<1&*��,v�آB9C�f@"LK�<�j[Xo�%@���w�EA��J�<u��7n��A��:C�P�I�k�<1%�͛$=���e�B�_#�DI�e�<�Ҁ�g��$sg&[Rd�s��^�<����R*ㄅ�=���nV�<���I (Q�D�s�D�'h�y�<��T&tj��;  ���U�0n�s�<� N�zw#Ł�<���@<I�D��"ONexrbD!)��9��IS,���"O����!��~��I���v��Q�"O\��N�!�zBjF�}Od�"O�a`)S+5�L�"㋖+�`00"OJHr	�o�*8AD�	�vq�"Oy;Q�ˠ�$�˵���x�c"O�����\�1���O����q"O��z�D�uI�E`ÁE%$$ZW"Od}!T-��~9���� �:�Q�"OL4����!���X�&
x�3�"Ox$a�K,�y oPW����g"Ol�i�a$6lfY{� �P��@�"O���S��=��܂1b	�>�^�ڲ"O��j%f �h��`Y�A�&h�[�"O<��� ��{����� ��.e��2"O�IQ�nj��+3TR�Q"O�5�w-�-͆T�.	�7>�Q�"O�
��ȇr?�`����z-V��"Ol�Pd��<�Ĥ��J�����"O�t���-*X���Dj���j\�"O@U�#���6�E��˲@�<�C��#��ź`
N/C�<�QE-MS�<�4!�E��DH�$ѩ�U��OD�<y�*�D��C�Ҿn�Ph��n�C�<Y�g����pmM�S&��.{�<�,��/���`�*̼}��3"x�<��υ�B@�%1Ņ��$y�TRV�r�<QT��
n~��� aNy����w�<���*,H���)�&h�!��k�<�6Ǚ�C���B�鏣#���ҭj�<�5�\�K��(sEDT�u�͓�/�d�<3�S�\9�$�Y�1(h��J�k�<qC�(6�96�M�{��kg.	i�<���"�.���
sQ�$��b�<�fV-D{Vx
1d��n�t��SK@x�<����r�ڨ�3dԽ3)9�N�u�<Y� �3
tm��]:a��ᨶ�X]�<����x����m��I�`�<ٶ	��~4�r'o�[��вe_f�<����k����OC�ʴ)�id�<�Ō��n�B-I�`T,\��;fN�_�<1	גO���Њ���1LBq��g�@�h%E�9l�DQ��ș|���ȓ+Rbp�!�\Q�i��_��d��ȓg^�|K�N��\�T�����]�*<�ȓ `�U"��ľ|m�,3�a8oІȓxV�4Iw.�1w�Y�!ܮ$���ȓ���S<N,�R�.�'
$贅�U�^"ԣׅ��R�T�R����9P����?r0a���%BԆ1��<��0�@%�n[���	: �!�ȓn���-�"e�\�{ŏ��V_���ȓq�j�P�
CG
��A�� M��ȓ7l�H�Tm͌d]���������ȓs�J� �8%p����#ҿ(��T�ȓ*�N�8��N�VZ�@@�K�
�ȓnv8i�����ј2�C��I��*�@���u|����?m R ��n�jL#ՊΆ*�v��tc��~�ȓk�d�����AV�u0%��MDv�ȓa�����& zm<��� T*2�t��McPhX�぀ex�`A�Δ�;�t���sg�В`����hs	�#er%��S�? �q(�"Ծ ���F�	�Tp�m*�"OH5G��W?���@�ТE�1�d"O�A� �V\��Ԡ��]		Dj�r�"OT�[��	y�,�*!D�7�IJB"Ozػ��9!�fQ;t`]*��`��"O�p2B�E�X�ȆDF4�.�q"O���w%�����y�Í��0��S"O�1��B�v!�W�K��.�8�"O�Ċt�@D=�b�J�B� "O��adb���H4�TcڑԈ$D"Od���̂q�4�@�5`z(��"O��Z�M�h�*�L�,��Q�v"O��@C�-4�伳E��8�fpCC"O��1lͫ<���DA�\��aqR"O�L��L1v$�n@�Yd|"O�T����	*�2�B	�AKdq�G"O2��a	TIĨy3�`�"Hp�d"O��K�;Cf��W��IA��"Oݪs�>ф��%cy�4�sb"OB�9DM���I��A�_�(,�4"O����'J&*�>�X#!�+�D��E"O�K��(l�Ȉ��-�=��` p"OV��h�\*؈����mz�@V"OH@p����TɃ��_�Xt"O J�:P�[�'B��`�d"O �+�bJ'C��y'Oִ	�ܴ�a"O�SiO$��(*n�!tr�b"Oָk󡛇e�.�J��B�v4,��S"OFX�1�Ŕ�~�酯��{x2"O��i������H��t"}[�"O�����̴������4D^x�8�"O�]�",}��`2`�) �l��"O�L�g-ۉ/�ލ 4�B�x�v"O�걨�U��qh���!�N�S"O�Y���� 2�rTx5Ȝ�T�ج�q"O*D�t�Ѯp@�xw���JW�]��"ODL�#�6����*��ec1"O|�yՋdb�-��L�T��l:�"O�I�Rm�#W��5()_f�́"O��x��mt��X��{E"O���1ğ&8���JE�S�lP�-ʣ"O8!K1kF=�H��bҚJ��ڀ"O��j"�=?hd�&C��C4���f"O����A��b�E���"O6d��ϗ�s�F�B���%r@e "Oni�ŬE�6Egn׾[�`d"Oj- T�#~�ƍ��,��H�<�C"O�����T�[�P���X���EK�"Oꕒ�"�A��)�ɮ���"O��Je�� ��!��-� (皜�"O:�Q��M:0l��:#�	�g���"O�}�΁�:t4�b�+ɢ��h�"Ot؊�hF�츻vj
�h��0�"O+�C��@h7� m{� x)�t�<��^��d�jSb	��# �o�<Yp(�-�h���X�]���C��m�<I�$a�駃�'9�p����<'dC�I�g��U�ݶS���v��F�C�	�&��W������c�w&B�Is�	����m-�0��]�"�B�Ig��X�$"�.��|0%�h��C�u���8�O�b���tm���pC��w���k�DC�*>�G�t]8C䉗0�6��L��N�03���U/ C�)� ����S�6`�U)J�$��"O�8��V�9�����G8s|�"O�p�� �,�I`�9C�m�w"O��*��8��b�EM22\�Za"O� C`Y���ـ��Q�{,�0��"O
@�����6���烑ABt<"O���`�?U�(��ȵw�hH�"O,p�ƀ���~!"�&O$}�H-��"O���(�4(����80��u"O���։Ѓ&U̒��	R��sV"Oly�a��#}h��3�j��]���"O�q��D�_���oQ9�ZE��'bPЄR�FGZ��c㘭e��e�	�'�� 0*�LȄ�0�a��a
�'��{��M�x|��W�ҥ\f\͊
�'�l��'i�	P�mȱ�O�by���'>�@0��#���ɁJ�(��]�'A�0�͟�3d.���h�?2�b���'T4�p�^��@�B�-.�Z�'YhT���F�B�P�f�,�����')��
%&lX�'H�+N<MH�'͘L��m�9X�p��3[�JD��'N�X�[3�dSW��<z�'!���q�m�s�{k����'��!������6�Z���H��'�z�y'��բ���e	 {�����'�z�e��
Xeq�@�x��Xb�'����V���{�DQVe�(C�MR�'�ث7��
��%�%��Y,A�
�'l��
:]Rl�:P"n����'A&�PY>`�܌�d��ktԩ�'`���f̅;<y ��TL�
j�T�A�'FN8��L�Svf���d$����'A<�{U��Kh�t[�'k^����Ib�@�D+�<Q:p��
�'�(��m�#Z\K�I��]�Zqb�'}
������4u�D e��g����'���`�[�z�v<H�cV�]G`�X�'��<��)V�x:����U6G&5��'7��P�&�0<R��y�hlq�'�N�sw���f��H4u/�i�'N`�N	��� �m�W�x��'r�
Z�*"���`AIq
�'�t�s M^.~>�-T7��Y
�'��E����G����60f��Z	�'����C*JK|{D��U�d��'\~Qpg.� �Z��t!Z=BsL�	�'i��B�ߏ1*Y��U�/�̬	�'u��Hd�I�c(�R��[z��`�
�'�D#̯ �nI2�����'G�y��o5,��{1���m�J���'��:�K
;�1���X�m��'m ����+�&�@pό�i�,�'@h�	i�%E�:�ʷ�4[��
�'���a�=,ʌ����:���+
�'� ����[��t�A�H.�A	�'w��;��_#���&Aϻ+v�[	�'���T��O�
�:�,	* �-��'-f] ���8�X8+G�M�}ߪu:�'�����n�/X������|�� !�'0�<�wEE���1��� �l����'
V�pp���,*��h�#�c6��'�ZH�C��;Q/yX�h؈)rT]��'5��g�
j՘��V#&"0�0��� ^�1�A�i@h 2�_����`2"OP��D��+�l�f�����"O2�����!U���딙&��b"Oڴ�ƃ�5,�VdY��d�"O"�� �ޫknu#�ȉ"y�M��"O��+���[�pka5v����"O����%���! @�"eT�U�"O�M0B�[��2���5DT��"O\�B�g�13�� `��NU��"O��������T�_ߪ]�S"O����W7azz�@	Q�s�I2"O���IP�'���A�h
�Y���A"O��3��	V I���N�F��"O8-@����$����%\�9�a
p"O��Aԫ) ��HuC��~%H��"O`�Kٻ��A�p��B"O��J=_�@	�2A�%:��`�"O��qV�ڛyoF���ͣ;E�[�"Ov�٣GX���ad'��<W�ġ%"Ou��D�',�XK�$��r��{�"O�(0���,���B�ے�h3"O0���E,�꛹Ÿ́�G"OP�cR)�7��`�!	Ռ"���"�"O�Źp��=^^½B�_�,�*��1"O(p�+E!1�� ���{�,"�"O֑z�e:#��٧fF��8`�"O��iZ7n8k�%�rj��h�*ODЃ%,���R!�K�,_��;�',��$
�;̮��ᅜ�;�i�
�'�f��V�Y����Q��(phC
�'m*�b��!w+��hBI�#};v�[	�'�`"���z��՚�g��^P���'䎰BU���K�@�/��a����(�y�I[�pٶ��T����"b����y2$B�N�E堅-^��%>�y��H���!AbC<x-��!��J �yr��+��{VĜ3v͎\"7+��y2aޘN�Hh$�^v�x���/�y�
�(~.$QAC# �-s��.�y��
�qf�"�F#"���s�hH��yR�f��:��8kV$)JSiŴݖC�I2C��'I��P׾\�� �A�TC�	�#����Mڹe�J�� �Z:C�Ɇ\�ܙ�Ɵ,_.k�'t.<C�ɚ�^������26 `�B����C�	��8�󫚄r���W�C�3H�Z�+&��W2����
��B�	�B�DԚ�.ɊLV�!�ՅI;p�B�	@���;7J_@O~ՈV�)l�B�	g8�� ��=z���ȷm��C�I�s�5	��3�@ZVA��hC�	�|О4"V��D�@q��$��ZC䉅r.�y3G�!�>�8!B�;zC�	��(}�U!޶C_9(�ޯ%�:C�<=Dz�3��lD�R������=D��b�
* A���,.gf���0D�DS#1a�x�1/5eQB��f0D��qE�O�E�q� �9H0g�,D�����p���Ձ3`���h*D�dK5#�8����&-�8[�����o-D�xqb.� D(��9Do�ڈ�S��,D��'l�n� �V횢S�h����+D��I��[�])����kTn�A�5D����O7R`R�I$�I�:|�1D�� :1�s���_�>U��ܼe,��"O4��a��+i�n�.��3��!i`"OTu�fd�3;pd��F�-MJa"&"O��� �&���A���L/4�Z$"O8ȹc���r |522%G�3��� "O&̡�&����A�Y1p�d���"Or�SJ�x�pT"c��.~
${b"O`��Y#�XM�v`F.Km~H��"O�@�o*-d�*e`e]N��"O�M@&#ֈq�n�I�Ω<LJAG"OP�J���x�1�B>0I`�I�"O�8�@�x^���"\01Y�"O����S�V� "D�;�.`�"O`racH�`栤�j��l6�eS�"Oh�RD��)�l8v'��'�@p:�"O`����������f�=�.q��"O��˧L@#0>���D���H�+!"Oz)�_�wni�g��8&�Y�"OP��ˏ�/��m:���V���C"Od���IZ����H��-@�~�C�"O�q�I]�Hv�T����\� �a�"O4���,.4(�pK�=_�L��"O���lC(�	1u̯�1��"O&q�
�,Q���!��J���`"O&�Q��o�,��7�(u�}("O܌�yk�X�&Ä�7hB��6"O�	#���2+\u���Er]���g"Od�p�ԇ~b}�O�R�A2"O,S����ekh"��
%a���R"O�E٤�
 '��3�jX1�V�`D"O���mݪo��L�7���y�H+&"O�8��d��f��sv�2/���X"O�i��r�e��!�:Vq��a�"O�Ͱ�K�X�<��@N�=oX�Є"O^���/[��P��!;J�pv"Oh=�a�
=nș��ϔL'�E�p"Ov�����=Kd�� �:?,�C�"O%��F�4�~�ݸ^� �B4D�LDH���N-he�.J<R�:S"3D�(�&��&:z���l�����1#/D��R�h�6Ѵ]� �^�I��ɵj/D��1��k^����Ȩ[<��cK-D�ty��A�6°e�!�Ҋ3�����6D���EiF�A�>p�"cOH���*u�5D��1ת�'R�����@ �d�R�1`3D�l��`�]�F��*H�!-0D���k��w�&ܫ+�>�<��v�)D��: ��U�6}AdU�� �*'D��J�+�$g�dH�\�c"�|�j&D��S�O4�<��Re�RL�A�Ն"D�l@Y���A솆bf5�K#D���t�W�p	t�!L�A�N�0$K!D�T{giG4A >a(I����$`�� D��A���^*r�10�	4Uh�t	�,D��ʱFU�u�� �1�Z�f~�Ѫ�E'D��HF@�5N��U�E+O�~��Ǌ#D�hB�/�^�BCb���^e���3D��(�J��������h1�͠�,0D�)CcL�� 0V��D�~�9�.!D�	�v� caA���Dr��>D��Is�΢[�A#�D�-S.N��f�<D��٧��?QD��ɂl=r�4�Al;D�X!sX<2TCA�I8�4M&D��hT���|\����,7l��%D�� �L�R0bdZ!��((�|���"O�X9b�<� �j�!�!x�p��"O�TH�̈́7]9n���@6E�ʘѷ"O.��5�����@E�\�Y�P�X1"O���S��KR�,8d�ś(@t��"O ���C�e����ƥ 3P	'"O�4�6�&q��;`ɓk���"O������, �	���"d�N�4"O0I���yP>���L�=�"�RA�'�ɀB �#�@�# 60Q�>{E��]��t�GC�������_)20	�3J*D���	:�d�����S��h9�A>D��*�"�9pT��J�b�̨+��'D��	�EF��\p0B_�?�����)D�vd� ��ݰ3��*PD���	+D�`t�Mf����!���'��=�m3D�D���Ʈ.��FD�u}��P�1D����%q�e�oٙu��Mx�:D�0ӏ�-#���ą�������;D��9�ʁ�B�x�!� ��NLP�e.;D� (�5
$D�A�U#�*0q�/.D� �pÜ��8w��&2�"���+D��;�.�UF���wO��ؙ#-D�D˃mū)���aeɥ)�<�l%D�4���x�|� �]�3�H$D��q%D
z).XA��vF�$p��"D���A�Y�Z"��SK	M�x�bf"D�h��镳S$4�R�I�8-�K��!D�|C��5�\m��ƏH[
L#�l%D��'�Bz� H��<I����(D��i0'K bւ�#� �7:�Q�F�3D�,)AAC1k�W'�9��$Y��TC�.Wi�%��!k6��� �Նi�RC�	=`Ȍ��I!7��hC�BT@C�	(�l����	ASpT�C�1�!�DC��0�j��k�b����Q'R�!���}�*m(SaV�X�pAD�2�!�ۂ1X��Q�L%}�^10v�+e�!���+h�K��֬w�f�*��aa|��|�h�Yq�%h�VMy!׉�y�˞�G�\b����p���:�y�
���X�F�@ �J��QF��yB%��~���r,�!p��q˃��0>J>��#�7�H����Y�`2V1:�*�`�<q�MS)�v�J�6-N���PY�<v�>%ҤbE 4PX�d	�oX�<��.+-)>m�j
�z+:� @bS�<�J�+o��D�Ťұ@���`#��Q�<Ibmڏ���D) څ�RPJ�<	�H0v�ꖣ�$~U��[k���?��_�O�` ��7H@�+�h�g�<����
�6��e�!-�L�Kp'o�<1��V6"�)G��X8���h�<�����}��p9U�ܑqX֨;���a�<��m� �8�.ِ%�r����Ka�<�e/U�X��Iq�⑁-��t��df�<��AF3j.��)&N 'kq��铥X]�,�IY��X	�A�,ڊ"p����6J����8��CE�Egl�x��M�Q���ȓT��vG�1��Sφ�'``��	�c�(Q��j F�&W��Q��n�h	&O�s�"�Fh� _d�ȓE������b�$ ���ȓT��{s蘄s����̮/`�u��S�? ��"��\&=B�MC��O'^��y�&"O�dB�$ۉ<@H5XT��VH����"OZ�j���36�Nɛ�k�[<@)�e(7���hO�(f&V4͢� �IW,] �"�"OZ%$��lg��)wI�7[�.T26"O��11�S��`��G3/����W"On������zh� (��^ݤ9�v"O�EYR�V4�]�4-
8�,��"O��H���2qW��R1é<��S"O�����[¸��s�O�r���3"O�m��؂C�z��Vnفu*>��#"O"1�ać�X�HI�D��Bk&E �"O*��Cg6�pČ3
g~T
�"O�<����9`W��"Q�#�&as��'E�O*�2�H"1���f�HFh��"O�1�d Ր��(U,=�m�"O��+a��fZb�{���?X!v!�q�'�ў�#I�v�x�J¦G8|��A�s!=D�t�P�R�_�ڃ��e�b%s1@5D�@�	�6�2T���96�bX���.D�(�5`�&�P!YphO]����(�	@���O��10gت=�|)H�ǢVF��	�'y����t��U��"��N����'�nz��,C�.D	�oI)E� u��'�$0��+؏T7d�3��&`��'�Иi6�����&I��jTA�'3jxU*_u�~�Q�Ȏ�qk,x�
�'�^��B`O���"I��.���O2˓��d-ڧY�,�¦B�
��`��&M�fE�'H�}2a�A,"����7��������y�ȑf�u�1)JA �!�q�A��yRFoi�<C�J�aIuY�ϝ�y�b��-�9Qd� �i�X������y"㕜�(8�-�<  ��)W �y�FݽEk����G޸;��,���\��O�����\l��C�U!p*�p8g�i�<	�U�F�x��gM�)��Y�gKEb�<aG�5l�P���N�u+W�.D�����ڱ*.��b�BP��1�+D��ЇcˡL�f�C�B *c2�jv�7D�܃7M�0�E�s��JQ��� 4D��h6��~� �#�A�8!��s�<F{���P�~H����ܳ���c�U/ ��d.�S�OZ��/�6_�T�g���g���'��8���ʃl�b�杇eX�:�';ў�`��YXn��C�ױ6��K�!5-&L�ȓN�Qr�L+EJ�(pɝ�-B8q�ȓ+ڌ��@yZ��+�
2!��܅�S����`/=:�K�*K��!���s�$��K�?\��p�ݲh�LQiV�#��<A�ʞ
�ܥ��$�50�(-�5�H�<��DF2]Y��.d��� {�'�ў�'j�:���&��0��Wi�y��7��8J��\�PUJQ9�K�{�\��o��b�@��c	"%�''ع�pP�ȓ	z*��2˒�^H^a�ԍ�[�~(̓�hO?Q��>^B�X�N�O|�e2��>D�t�!eǜV�ڰ���Βuź��D)!D��x�o\#;�`��!�����1�!D�4�'��8���RfE,ށj�n?D���g��T�B	�#-yp�8��!D�x�j��iu�h��N޷ <���<D�,�!��S�܀��A�9V�$D���G�D*t`�-�o�a�q!D�� ������`l��PS������!"O$�'*9q��yI�+L��&#�d/�S�'a;p����F��G�)DV���ȓ"���j����\X�����ɣ0T�ȓ8B�SQ���d@e�^�����Y��TӴ���]�3
^"5�"��ȓIpp$���\;{q^P1+֢�eΓ����<)���Sv`{�%�"O>:��g����V�TPġ "�,���	Z}hϓ�hO��#��8	�1 sȑ`��&��'P�B�	�g5z��,ޗH����G�L�|B�I9��J�$ߴ{8֐��˱/�JB��68�%Q��]lꍋqd ;����?	�S���ĜW�epw�3�������G�!�D�5F�,ĀL�@������&�!�D�*Kƴ�R� g(� ҐM�!�DQT�pX��Z�_&4!��?�!�dσD��p�,� ����/z�!��K�/m��#�e�F���MC�-�!�D��G&��C]�3�ّRL�v��`��I��&�Q�����W��(Ę���OV�=E��- �MR�V+|��� p� �y����5:2�9B��)H~T��!̿�yrd�-fG�=(�EI;W2F�q�����y�e@�w�T#��!.���f�ۂ�y��A4�:y�N�^�J�Pi>�yb��0x{*��٩E�V�3�mX��yB�ձQ�6XStɴ&K�4�і�y�Z�p��,1�R8O�<���Љ�yR*[7stl�۰��tx 9�rn��y�GBJNH���F=erڙ)�O��y��2d�|�Z�ٴ\�����ڝ�y��6V �i�#ά��V	��yB���,F���7E�2�ru�%�Y&�y��G5[��U�N��'H���HS�yb$�0	�� qD�ӶG��1�	��ybȄM����/ׇz+��
�.X��O6��v��^�d�G� 6];4"���C�<APF>�� в�.O�*e;3���<)������z!!"TL"`�sMIx�<�1a�E��l�Qf�h�^0#��O�<Ir�Q.r���y&�@�+9R�DD�<�PjD� �RQi���>"᪖B[h�<�P��'4�x��Ε3<��T��b�<����>�00R��A�Ԩʕ��Z�<I��?�n�����8GB��BgL�@�<I�]<i��F�g"� �S�y�<9ć%Hl�u-B��^a��Eu�<q4�^�m��@��,ƲX�mi �n�<��!��oH|�I�+W�[�]��l�<ѵ�/�v���K%L�����O�(��x�mE?E鈠��D)AK6��C@�y���j`��Ё�7D uᥫ��yb�T��}��+��1��$�6l=�y���/�Ye�� a�ıFK�y�ݼm�pmQ�Jr��h�V�X��yb��>Ci�� �H�l֪�U�(�y�]�>bOԧf��iY�HK4�yb
��h��qb���M9e!�	�yR$K�zj� 7�z��=�4
�yr�L�,��ps��2q�ء#n]��y��aj�`�F�i6z	C��y�E�b�X[P��AAL���y�M��l�D����E�qP�M*�y
� Ȅ��#Q*hԴ���F�2%�� h"O�yP�X�iPl�z��͔|��iP"O�̪dDٽw6X���:g�� 3"O���myp<Q�c
1B���"D"O�qh��C�����C� d����W�3��<E��'YP�X��R&#:��*���r>����'(�҂L�x�Re� s�V�b�'���cV%5��HQ��P8c���ʓAx��1cE8��|Zt曄g+0���8�@���bC�gMj� �'�<��ȓY� *���NM��dJ$|����;sT١+�ez�i��`B��ϓ��)��\�@�gTeVĠsu���B�Id�ʇ-÷}����2dϭ>����?��0�@{CdИ�@���xhz��$���bq�͊X�`� C��%?�lQ�'$b�'�P��v+�0�X�᫟+A� ��'d�Y��+ڃ-�����(�Ơ��'Dpd�D/Vzq�%�9Tȁ��O֢=E�$HO�(4���H.t0�q ˗�y�G�>%�LsaS!�LPc�����)�O}���6V���r��� 4Tް�"O��I��2J�:�͚/�� ៟Д'W�y�J�sbX�X�'^bm�Uc��y"dJ=]���:�Nͬ\yd�r���)�y2]&A�E�7	NR�`�	UIȇ�yb�P^\�t����tf�u!D	
���O�����8hz-{��;P��xcD�J~R�'A�\����v��Pҫ�\�z���'�|�@r"�%7u�6�V�Z�4��yr�'İ�j׬	r�����W�a�'�F-h� ��kʚ�@Ư�7OMfr�']`-�6(�iPYȔ>Z*���'� A�CʱO�$��#Ն B��	�'�h}i��^�,��,+��Y<*ѐW`�<1FN8i��LrG�W�.�(�CU�X�<�W�L�2Inʣ��-p����y"NK4I�n��7EQ;J���L���y��(�4m����j��Ũ���*�yR#�� �(=�&�̥4������y�j���e�H��
<Ap4%� �yb��qt0�Zv�P+�6t�k��y�/��HpL,*�O� �b��R���y�́:Ps��q�&�~����`
ŝ�y��LM��		�*E{����o��y¤ =S T���Ӊ'Z`�R��+�y҇ҵu�&�r��2&�6l�%���y��V"��1��R��5��	�y��->Z�A/O�z`�aEOW��y���7X�𓠌

zP��Q�G"�y�E�?�P�0�N�k���� ͌�y�㑙O������v�R=��X?�y�7�p�U�P�>l^�+��"�y"L\i�D���O��'�H�y"��(�L��&0�DQh�Bݰ�y�eס��@��8S=&��sB0�yrk"E+�}�0 �G��*�� �yb�'}�O?10'@�	����jʳ܄��3D���D�DtDd�z�+H� Gxtqe@2D���4��>�*��آK�bA  =D���%,��k�(0!���/�@\c��%D�����$h��7�Q/w��"%D���J?M�J8�H��ʃ���ybOԀ1:THC���{qE����ў"~�S�? ;ס��$'��+�A1H��f"O^	Q�yU~�kCR�{{f-I�"O�	*�(�	jS�l���]rUs"O�QXM��#�,�KvM˽i
TA�"Or���bP�tl��A�Q�6���!!�'�O^e���ںc�ʙc'L��D���Cs"O0���W#y��)Zը���Luh�'�ў"~�R��<�湪$!J�8�^u��{�<iV��82YrU��A�pZ<m���L�<�p홾ul�A�fXs�XP��"�@�<ф,��V�L<�w	Q�p3F�Y��@}�'.�y"�ۿ[��q�H��~/�	���,�y�j��w2Tpa���}~�A���y���,P�,�K�	��n�>(p��U��y�(��2Zt؃b�ÆR�� �F��yr��8b�$��g(�2Dz������y2��:d�`9 ��
�;��y��͈�y�gI<y��1r��O%E߂}C�+�"�0=A��h��b,���b�/+��:d��y���T�'�n�
7���a$��뱧F�BwN�8�'�X���E?���B�E"�2�'z`6jʛi�1�A��%	S�R
�'"��(Pe�qTp=����#SO����'��,�T�
�b��I��?�fp��'��4�
6��b�$A����'g촢эC�0�@�S�S�tAv�I��$>�'¸���n�(�PTP@��Zb8��z+8���B�UhR%Hw�B� j�l�ȓ8�Z�����+T�0]��T-UZzH��v��ewM.A����k�/=�x-��=�։���4��2m̓2��U&)2+�&v�:�{�E�W��y��V�v[��P3E����c@��	^�'��Ț�EY�G~
j+�8
�&�[
�'�l,��ɐ%LqS�%_48Cb�
�'��#�IS,�����lŤ,���y	�'����d�kt���)xX��'�T5q�e�`!��6r���*�'�X+$M?%%J��+��aH�-���'�������+���	$́�W�������'E�I$�8L��zgI<Q�~a��'V
=ڳ D�]	+#��>Z.Ġ�'oF���LJ�`��[���5��ɑ	�'i�䈣-F�<��Q0իՠ5�����'-TъЬ 7g@~(hէZ'_Ր�p�'�$�4#x�б35�.) iɌyb�)B�+�@��!�	����'��:���<�-O��=ͧ%�Y	P"�{\�PA��(�6؅�g�^�Z�X�&�pЌ�~?�D�ȓ;�l�c��7�L*��#g���ȓR��Se)�&�5K��p�y��͂<��b0zQ�7*7s2&P��v���3��8B2�iA��bþՆȓV =�c�d)|(��g^i$�F|����b6�Q-n��HJ˽3�4C�I�L��M�QeR�BR@���8R8E�	ڟ��'��Z�b>�	�*�
\���ЉT*P���BS�B�ɘ~w����_�z����Cd�]��B�I�)����AB�r,��	qNG.�B�I�Jߴ�r�e��\�}��i��)�j��<��<����c�p�s	��NI�Q��]�'�i>�Q�	�Sby����4��:#e-D�<�fiC�cW T�b��v0H�6�,D�iT�"�f���ږo���!)D�� ��s��)7$�1q,�9�fhE"O�K4�¡!-�T#�
Z�4ꊑ�0"Oxy#���#Cb���4I&u�6�'|�O�J��Zr�ȴm@�9���0>O��=E��I�omD1��Ψ^Ͳ�FM�y�/�x�|I[�h�f����0���'��]���'��O�Q�&R1*�(��p�T"OPi���S)m��V���p8'"O\ܰ�i�3�5�E �@ז1* "O�aж��y���q�/�$�ZE[A�'��O0�sd*:7��jsIԩK^�͚�'#�'2��[��v����e�% |μ;�'�ŋg��!մ�SEE���P�
�'uEJ��l&|\zѫ�*`iVp�O����>qƈ���+�*�#HرuH!�$T+%�����˸O�`�I�GO(0!�FDú���Y�,]C� (!��',��y[�R�L�K` P�`�a~"P�H�m�%\�J�����&k$P�v1O�=���Q.^�9��,��i��E�?���?���?�*Ol˓���Ԧv!pHr�F�@��k0�ߊy4�d2�O�q�	�,x`(N���#C"O������ m�	��?�2��"O"A�FD-rú���^k x��"Ox��"�:2U�d�gŪ?s.yc�'���|r���]H�� Da�2;�^��yB-LJ�pE��,B�U��R��Ӏ�y'�2z �DQUI7J�*���%?ܡ�d�L̹�B
�1D�f�U១]�!�$J�f����F�<g�M����!S!�7`i0�4ƭ�X��!S�Raz��'��S��H��F$<8X!��#ccr���f��E{�O��OP��F�CJ��![ac�N'n1C�"O��bmM�J����睜J�Y��c�<A���?��Ş��9O��P�I�(�b�%�sR���"O�`6h�!{"Z)��:�A�?�!�䝀h�yp�$ыF�vT���"�!�d�-nz�d{�%��(a@ �"Ea~��'UD�c��ls��2w���S�f��O����Q2"@��"�.'�.����W�D 1OB�=�|ztYq~횱��3ST�����<��F�	��(Lr���&�PL4��� +�⌁,/i�=q����}�J`��~k��rD�0X��h�Rn��i�ޱ�ȓK��	NZ1��d���`$�����?Aeӫ@�n����!8�4E����l�<��.K �2y�C�]�48�=#0�e�<�`����l�釬:�M�' ʞ�?���?���?��2_�x�t�J!)F2���)\�Tp�I)D�����Ԯw���R�m�}�^ �,(D�h`T�q���d��	b�E#�&D����֮i�`����YQ���%��C���)�O8U�#O0_��BE�E`� p���<A��4�����J9Am⨐5+�,\BP��'�t�R��!���huC�Eژ�C�'���''�X`�F,e¥(V�0�Y��'��E��,Y�m� }��y�"2�'���X���H~�aC ���E���
�'"DXIe�ϫnEb�аG�)9�R`!�'3�ͩ�Cf @drs&;[r�p��'�2ݢk[����
���L,1��'O�eB7��!J�Ō�T����"O������i00H0�̕	`(��"O@�y��8I|��4	���8�"O� ڠ�M� (���qHܮCl����"O�t�U@��|��@�h=IMH��""Oz ��kV�3Ǌ�1��S-O42U�D"O<l��	�x�93�i���"O~���P�1c��9G޻x��Z�"O<�
���290^�QDE��-Bܡ�r��O����� gkP�aV����t٨�I�+!�$+�p�Մڿ5~�L#��ˏl�!���n�����L��T�E����!�d�|i�	yto��Y����S��j�1O`�=�|�2nJ�2���$�!F�t��Q��f�<�%� �n$�� d�c�Zc�<yw�G��S��xn��#4�I~"�'w�{Rko�h��wM4p�Ä�yb��1�>�Q�s�8�ާ�y�"�Q��E�"��S� ��q����0=9��'N F�D���g�Q�u�1O���y��)�'G�X�5.�.<��4�`B^	��Dx��)"I> 7�y���6��H��NJ�<yp�!W��dbץ�"�2�q΋l�<I��������� C�BL	����<�Ë�#�~�kV��8IoF=A�I~�<�U+�> �Dt*eN�-�<�s(U�<	�c#��-J$��'sd�!��kF�<��攰T� �$��_��d��%x̓�hO1�H�㰉��_�Љ���B���أ�'W��6ӈ�B��^��Z�Hd�_,{�<���>���(14���� $j7����`�<9MA�z��4Y ΃�E���S� �B�<� Q���t ��Or��3n��<� � ���	�FNL�& ^}�<a�jK3'�1������>�z��Cs~��'\�O>��sv��x��T�H9ȥ����>���Ox��TM��|ߊ%� "DN<ZU�!D�z��
�b��rҭՠd_Tl3D�P:����	i��"���K��&D��B%�S�Xp/ˤd���y&,1D��@��ڧ�.�+�ϻ8l��2�*0D��b�@ǡ=���Ή �����9?�H>)��	ƊG�9��(^<ƈ�WF_,���.�O��Q�֟3�%"�!Y�r^nz�"ON�RR�(R2$��a�1`M�t��"O�)�F�ϰ�����)v3vy2�"OD�h�lE:�ԉ(�N__u�P!R"O80���
*�L��Ȓ6kg�%s�"O������w�nq�7�� ,DA84�I��LE�D ����1K��iE^a�@�A �y�@ظrk�4bC�Z*t���­�y�G'bn�p"��Aw��̏.�yR���,Ь���.5rye��3�y���/1�r)�� e���4&O�yb�«W�����W����ӏQ��y� ��j�����K=<�0��Ymz�O����<1L~λ<�d�E
V��h�{�)Gs�hUI>�.O?�)C������ɵE��d���;23�C�	D��	��I��;#"�I��эL�HC�I4�<�R%]�m�$$������B�	�N|�xW��,6�����[T�B�ɀ7��q��g/MEҭ�4e�	��B��-�|��A?Fqv�cA�16��4���4�'���ɒ�v�;҉Q$[E"����
�{U�C�9_"����!��I��C�k�hB�	�]�z��jͳhi��/B�	$~��Z�iJC � R�;k�C�)� `i��k(VK���W������f"O�}�����,���w��"O�H�VbV�'�8ܩ��S1jk�0�"O 홷�S�fx��q3�J0MZ\Б�"ON���m�V%�qH4KҳfR��"O�q�-!U�$�"�HȪw��	�"O�����w��Ϫ���
"O��2g�S�rR���S ��!�r"Or�	����TX���w$_��f�{B��O`��6��<E�C��& �-C0!H�E[$���ybɚ*^pњt�L��%X�C
��y"��}-4�8�m���{��5�y"�E	 E¤�J� e��/��y��	�����hő�bW�y�(Ҡa�8�*��ڷ
ʊ��#���y�	O����#�N4G��#��?����<�(O��O���L���r���x(�Ï�!!�C��ϟ���$ď/d��{�-�FQƼ��&ah<9珒��b�a3���+ �\��oEK�<q�Β}qH��Y;/d�7�PE�<��D;j�; �"�Ġ�~�<�+ҿI�>ȨA7%>�u�Q��|�<i#㊊8�8j��\+g���ST
R̓��$'�'u���v�1�p`2t"Z�Nȴ����ʟH�ɡ^� й�@��r|E����5]5���s�,���c�82  <{':��H��Bw���<TFlC�P4v��l�ȓ}L��C��c�r �W5�ZE�ȓ)0x@�c��	�(��I�
x��ȓE�l�h'��P`�6��]"���ȓF��4K�A�!.�i���J./c.}�ȓV&��YBhP�(mj��C?p�p��H�iZ��C�J��T��YHȆȓ'M��uM�|,8I3e�ܧ.����,����GG�~�x���-��%�ȓmg�("e�!������~��U�ȓd�v��I��{�<�P��]����-l$h�ËANyE�Qb�Q���~Mi6OӠTT~��1ȃT�$,��L�ά��JJ+B4���2��|�ȓ7�dIa%� 1l���UHMND�ȓ���⃒:A��� �-S��ȓo`.]5�Ģ_����6��Q'D��SB��ւ�h�ۀm���h�����]QbJU).�+�]<zp��ȓ�J�����(u����#+ p����ȓe�($r���ty���V:�f�ȓG*dhQ,\iS��b�V�`2,��ȓ��`��&Fo�AB�_8M����ȓ�P�v@��wa0MS ܰS{�A��\�x��G�.���SS0/qU��#�&����'
Q��� � , �D\�ȓ��dsԏ�5*(b�
o�X��ȓz*���ҮA6M�6@�`�rS�І�sd���c�)d(�a�ׅ!w����n�c�.�9!�y���=:7�ȓ~���W�5��%�ǭݐ&`���)҄�Y�>�򈺄��W�u�ȓ+���K�"�����H��{gD��ȓM��q��~�(] �,��u�p4��U���@ ,�����W�U~ ���Y0TM�C��/{T�&��&��ȓM�-�WH�p�Ő!�b��\�ȓ<�@|W#�-���D��Q�n��S�? ������7�HHBH��P7����"O.E��ښt4D���m�l��D"O���l@����p��=|�9p"O��{Ë1>M� �D8S>^�C�"O>1�"�NQ�z�+��1\qHB"OT���nAGf�m�5@�&7�)��"O~��6%�ac���Ο7+��@+�"O�e�,N�jH������R,��9 "O�a�A�_��F䚧d��/,	c�"OJ|K�/��7J(Q���bp�hS"O� �a̍�5��$�k3�T��4D�1b�X#eOH	bM�>A���D�&D���� �N8���'�iR��J0D��!��b�.(��o�;)�D�
!D�(�g�	k��}��b���j>D�"�C� m�DX(q!�(�t��d;D��س�V�o"�(p*�'i���K%D� �e�P�f�8�;�+Λy%y3�1D��S��J4K�Д@PC��<"�!0D�x�����iꢋ�$"�lӵ%;D�$�@h^���AƦ�\���e&D��I5�ݨOE��*�̜rbz�8R�$D��0��nK�5;r�\�J�|\��-D����k�$^�<�K@�_MJ�9��+D�ę¯,a����t�7v���u(D��r���9]t8�'��(�ܠ�)1D�8�$��>����A���0o����/D���V�� ��L��G��o��-���9D��[g�� 3cԴ�-�	c,ČR�6D��I�(�"U�����Xh�(�.6D��d�:����@!@.��C#3D��͌>a�>�cfNQA���1D��ed��q)��s�Yv`��y�<D�����R`-�aX�*~�٧E,D���@JD+U��UҪA�Uba�2�*D��H4jY	�M(���5U��CpI#D�,0e`�6H�pc�1D�`,D�LP�E �R&'���b�4'Ҫ%X!����ugN,"�\�n戴sFΥD!��ٯ�t�B�-��i؊�#�c��d*!�D�4�@�0e���u)!��H!��֧�h�*�`�B�;ϕX
!�dΉg���)�OK
f��ń�)!�V�%�l�?JZ�����!�$ 9T���ҤCLa�$)���!�7IFr%��d`Tb�H��^$�!�$O�w��LqS� ���鱠�,c!�D� Q����uMB��������z!򤙧l�FB��,�b��tKW)4!���1�g�0a}��#���`'!�Ğ/=	�P�Ɋ-^��(��&!���*6 :�B�`��E��}!�d��b.�Dy��)>��7��-�!�$Ρ�"A)��٘H�r�)w&�D�!�D��z'
с�ɦX����O�!�d��l��Ơ QdĚS�Rf!� *<������"92����Z4!�d��zϼtc��/p��8��9r*!�ЭWZ4�ʡZ�s�2h)��^�!�D߀6FJ�jэӍ �a�I�6?�!�?nx�c���E�� �%��FW!��\�� ���E�/�N S���!�ă�9R%ۑ`2#�0!���R%g�!���4S�Hm;���h����SJH#\�!�� 8Y �\�!�X�k�Ƨ��\�#"O� �Ū��z��Pr���T���"O^=�Uᝓ|b�	��O��<��e"Oٙ�OW�"��T����1qq���"Oj�"3%O86MR�S�&q�2"O�A��%E9@��QNEO���p"O|�Ҷ� fM:1�1��d6��8$"O��0�d���j\QtlC���"O���PH*` ���$����vX;1"O*�;R.[_��	[�OͳE"OL�cק#t����X&N9��s"OFLI��ɨ;�T͊b�������"O���%NɼCITq����&w�N�s"O�P���
�����%Ɇ����"O~h�1-�5l�1���Nt	&l�\�<A"��,���1Ɏ(;=>�8���r�<A��ȪX��A{g�ܣzff����Fy�<���_3	x	�V�¹7'���Ew�<)�'�4��a2J:I�("��z�<��I�,w�D�q�9G���2���Q�<��O�0LLP�
���-�)�A��K�<9T+�,�*���/g����.E�<�G��)'�=!0D"�� ר�C�<� n�tH�a��e�\:�H�{�<����$&#�HX�~��H���t�<13e�9_@P9�D^�q_���	h�<Qb�;L�Ј�W��>~�`�#�Nn�<a��G�mS��v��70���S� �l�<é��
:T3 g7
�䫓�O�<����n�H�,�-������M�<I5JRMv6��]X�8lA�SF�<ɔo��,N�ʂ	ȏ��X� B^Y�<	�蜼]�"���-��P�X�Yv�KX�<��R5D���� �!�j0�5A�S�<AV��0���Y m��G�­#���u�<qiߙ4�X�$!�^|��`
]�<��C'I;���� ١>�BW��V�<IS���W�x: G�G�5� F�T�<��aN 1^d� Gב{o$q���F�<�&&�&b�D���
�l��"���x�<q�.޽粕��
Ϯt���)CƔr�<Pg�<;���"Y%ft�A�Mo�<�&O;(vn$��hءU�D\�֥i�<1卌7]c�!�TN��c->�j2`Yj�<ɦA�zd���T�x�fDjC�K�<��A�53�b"h�5gP��Wo�<�D�Ż:e`|8�S'q�0�`��B�<!��;'�E�%�<��8w�\B�<��a�O���B�_�D��R�	�<�0$�kGʅhT	�"�䄹�O�A�<���6Y��dkF@��tF��0f~�<A�JF�����I�e��z�/�r�<���K
c�хG��"�@chf�<A��ք! �q0�K~&�م�I^�<��lJLܾ)h�FB (�2�x�m�]�<���*'�Z1��a�83,���R�<ӃH%4�$�BK�U?�䳦mPK�<�V'M-f��<Qcl�-@r����H�<�6�F1\BQٖl�<�.���K�N�<��X6��i���ܑc�R���Bf�<qA��N����L�Tp��
Fl�<�P�����y6�
/�Yۃ#	j�<�B�ed���4cٽNU��`�d�<�v.��M�����7{L�1��%�e�<� ����`w�H�s�8m��P"OF��ª"*��Zgl���.h8�"ON�z���c�T� EH�{�T��"Oj!0H�"UHb�2��Ч�<`B�"O� ���C���t�E74u��"Or$�����`p���^�̶�
�"O���DF�]��딷/Մ(B"O<���D98$`���>�"�R�"O���hM�E���:�(_�'�(�S"Oi��ʁ<n}zʉ���1"O�])�X�o�25زG��W��Ɋ�"O���GN��.&z]a�@2`���� "O5��f��yˑ��+Z��yeLq�<��K7 �pc�Ӑ�yR	�E�J�H�ȷpY��:a����y�ǞDx�a��m���P�yB�� E���e�o�ZQ��)���y鑋tD�h����kKΡ+w�4�y��L'D��03��c܀E@V�ɸ�y��u-���%VX����e"�%�yb�M�7�l�&�M{����̎�y�C/|�l�A '�Fzvȱ��	�y�
Љi��%ヲ(	n9�L�!�yr��&)�y �E�������y� ȴA�hO�8m���'�7�y"�э-��|���ң7�y��痡�y�i�l����w���,ޯ�y��ۙ�,spXD-��JC��yBjG�& H��5OޚD�nxGU	�y��2R�(�1@M=��T��/�y�)�$A�5�a���X�稏�y��#=�&t����<�7��yRf�&Q����	؀Buf ��yR�X2���W��-9�eõjW�y� ރ4��G��3��=q6h�;�y��:����j͕{��pF� �yZe^�}��*^�n��1�рڔN<B�wH�)�.!`m��A��1��B䉊D~�� �ܘIl����NS)lB�	
*%��*�)�_�����T�"S�B���Aq#JKԀ)�����ԖB�I�,�����R�R��G�ԉJB�ɝ��=��Ǟ}��d��B� nU�`&��z����gLV��C�8&D�NT�X@>L;�ᔝZ��C�	�}�����,ULk�GX�E��C�		x-h�����%P"��B�C�P-�����S�d���� �2e�C�I�z� Z�r��e�ߐo�@B䉂J��
��$'
H���h^4yW�C�I=/8��W��'�@p]^'�C�ɩ,Tx��椔<<����eF+S��C��#&���0��څt|���M�?{}lC�ɦiB<�I[�N# �Br�Ѥx�C�I�n�&���B����y�g�=P0FB�I�D���1��=�ݰ�!�,x<B䉴S��qV@Θd�h����&$PC�	: �Ը���V��^!��M*EyDC�Il� \3W� 0i�DaIC0�C�ɩ��|��L^te�CT���>�B�ɏ'��80�U�(C�.o�C�	�>!�OI��Z�8�$	oPB�9�0z!�(gA  x��!�$B�2Jll�P�:Q�^xA0h��ViB�)� �����(m=��[ /@<��r"O"�9�%�Hkht�!��(9�T3""O�\�'ܕPE�9�ˤ	9Jq��"O���s��%yjx�`�H8�!"OZ iGGS ޜ W�]-F��2A"O^4DQ�\(:��9}0&�A"O�Mi�)G.I}�M����')čZ�"O� )4��Dr�2fe.N��I��"Ob=I�)�1Zx���c�l��|�3"O !m�֓^���1��%o�20�"O�D�c@D�z��(��g� ^��K�"OBe��3P>��T�``p�B"O����Ą�R�= �)��b]�iYb"O��s��]�"��0�A�`���w"O�<Z�H\�=\��0' 8��L3�"On ��F��X�R��"G��(�;�"O�đa��C�*5 R�)��@�"O \2a�˅a����74����"OV� '���QO���5�4v��""O���4#,"ܺ��R�?o�DCG"O��W�י1��R1�4P�"v"Om���9��`��FQV�4Ѹ�"O`�UF��k����R�^)	�"OTIRF�I�>rv4[0)Ml�c�"O���GetN�{�`�%�jd�"Oh���F�#�9�A�Ҳ.�����"O�%QdKE/_�
��.�7>�6l"�"Ox��t�]�L���4�Ȧ��dc"O!���v�<Y6�O� �ve��"O ��犹r֎�3�`ϱsX�4�b"O�	�W ��9����NB>Q���qV"Ox��ѯ @2wv��9�A"OT<s1��@g�e8�o�(�LQ��"O�(a��?p`�aUɐ��a�""O��L?hY �[��&k���"O8� a-8OB(���A�x*w"O��CA6�t�[dJӗy�̩V"OP@�(�~3�����B���2"O0 �4K��`&Z)�"tH X�A"On�AP��@	���O��Z�"Oڜ�.���B(��6B�T:�"OF�Bj�WO\}Xp�
3P��Mh3"O8��ĀrsRI�u����8��"O�k�%�|����$T3��ä"O@Q��K$���bF���p�"O꬚c)L�[�e �_E��Tc�"OHh�-�C�r����	%]����"OT	 ��<s<б��
 �����"O0���V�V Huo�\@TT�"O��)����p:��t��~7�}��"O�4���	�� ��[8����"ODı�'ٝ"F�l���	�!7H"D�D�҉Ra�􊶅��#|���e#D�B���x&vER����C��qhׂ D���ׯ��#����K�B��(h�C�	D���b�V�@��)V��A��C�Ikd̩Z�����m[d-UT8�C�I�P�zU	�:A5�Y���G�x�C�26z�k�e�����Ź&(�B��sl��F)1�A�G�VB�2�Q:�H[�L��gB��S$B�	7Bg6<ِBTKe��R�HB�3%�R#H:Bp۲�ڞB��.	Zh�1*qv��i��9uB�)� !�E�	$G��@���R)m�l�"O�4B�h`u�	��&�01��#�"O�kQ��焍*!H�p��8�"O>a�w��SŁ�L<(�r"O�9!R�X:|��(Ձ	��#�"Oޝa�F�.Kܜ�B�F��e�l 9�"O����b�  K���jTo�|A"O2�)��ʙ`�&�i�[�`0�"O¨� l�v!	&*R*8�8x�"O��P���-�(�W��`.С�'"O� ���;�9�F�I,(!�"O:T˶�V	�n���ە.��"O���*��mY$��Cڌ~���v"O���CM�%s��8��ũQ�"�"O�A��Ϗ�AU���̞<jl�Z4"O���AgG	g{��ec��b�rػ�"Oڄ3��T��$��N�`"OH��1&�?Y�(�����6��[�"Orp����~��ir�`�E|jٲ�"O�Lxp�U���q�s G$l����"OR`�D���t
��!��`R�DBa"O.q��:p9����B�_-*��"O�} KҤM^p�R �<�y�"O��I���|Aڗ�g� �'˻�y�X�S�ɹ��ƣp\0��$���y����A��Q{q��d'~ܸ6�́�ybo�X���	X��`�&[��yb��&�,�q�D���	�C��yd��T�"h���и  �<�1KG�yr��23�6�!TFړ�r�p��=�yr�
,b�l"�,M2^�A���W��ybm�0I��M�椋r�摈`�
.�y�lE�p�x�AŁҪ|���#�yb��&o��p7R	�� Cc��ybF�$Lj��"%����B΅��y
P8n�� 'ɒY�#�\��yDʬS*��s� �/�	�����yr�4B̊��Gf�{2���B$�y�"��\b� +ʈA1�e�"L�y�K d���3F�A�6I�_/�y2�U< bT���ߪ1�yP�?�y2 ��-���P^�<��5��d֠�y���D���˦#�9~��/1}��ȓ{��1�O��P�Dm�B��+0�h�ȓ7�!K�$V$z(y�ר�4��ȓ0��̙ͺ"\iA���g���ȓ6��]� �LGs��8�/��'�t����XP�%@�~����EW"d$��1���cGnQ�Y@g!&��Ȅȓt��H�j3�=�KR���e��.[���2i�	k\�GA�+(vX��>���qň/v��8s��Z��P�����,Wn��jZ�{R�Ct����8&�0�$YF�PMG̍U����_�X����+qd$p��`�����zl��f�B6j�,��&	r:n!��~��xs���E��U[7��y�]�ȓ=��E
v��WD+�e�����ȓ,�>�X�ƍ+oA2aPp*�Dy��R~ ��B�QR���A�A�M���ȓ7�I
��Yt�� ��׽����ȓ;�F�������Ql��xg@�ȓ>Y���$Tl�T�I ��U�ȓY+bpz��	M �[G菝9��<��S�? ,j�e�;��PQ���2u��uRQ"O�u�R
�<C.!��@0Q�bp)"O�E����]W��0LO��~�q"O�,�+�xD~m� BA����"s"O\�7m]G
i�#jL }���A"O���+�5Pʉ(�)����ti�"O�P����'�]��ٝO����"O�S�L���AT�O���"O�}@#����{�&;3�$��"O���/�<o�=�S"[�x#�"O
p��ߣ&��1��T����v"O��3�B�̀���q�u��"O�AF!
H�ր��6m>�q"O��
��iٺXBN;%V<��"O��r��E1A?�`p�MV�Y@"OFd3Lۦ;tf���L@Q<h�4"O���$d�����ta:ͺa81"Ox0��k�[h��)���b̕�a"O�	Lժ|�`-����n�TA "O��q'mA6S�4�RS
� +X�9�"O����C�b�C��,X
��"O�׊/*��rצ�.@D����"O����B%-�E���%R41"O�(dDˉBt��b&�N�E�"O�(����F���;դ.�`� �"O�u�4�ơp*�li���'*���"O$kqd��1�Q��"��V|�5Kp"OιS���.)�,�Sf̨r"O��� ��q��TҀ\�+\ƴ�"Oh(3q̘27~!�V���8s��6"O�cC�£����T�i,D�U"O���2O���h%���)�Ne�b"O��0�
�eyT��B�vp�("O�y����i��dH�b	�SSQ�S"O8�ʒ�V�o�
b�!�r1�%{�"O@]��"�Y��2%O��/��!Q$"O"���B�$݋��-���s�"Ov�QC�^-
�����(߼C�d��f"O4����L�Je�8���T37z�k�"O��b��I�x��� ၧz��5�b"O�Yy6	ͩZm"U��)�,*�Vcv"O�M)�N5NTD����w��AC�"O�Uء��j�h��e���q��"O���3�U#`Kt�'bZ�4@Y�a"O�]�mȷ~�F�E��zp\aS"O<-����!�$����R�4x5�A"OT��[���	{�lY�n}�"Oju1��B$����1,Λ��d۴"O��M�u��q!����e\1�"Or`�`�ݼ60QeA]�"H:p"�"O<Q0%��\�,���/�y�T]�"OnEh��T=D�S��8��$��"O�P`�ͯ�~�d��=�`&"OZY�U��6oB�8�Aś"�EQu"O��r��*�� ��ɟ$0`�x"O�њ%�ܝQf���(!+'Ęd"O�I��J��9;'@�$VI�"O,��W,��^�U�`@?@"��"O���2��|pȭ+`ԉ��́"ON<i���8c��3��
v
xBc"Oh1�.� ���k�KLwrb)@����D{��	V�]@l��2K�Z"5���4{����G{����q�I��	��U��]�t��B"O���e��n└��C;mV�,;�"O� AࢌZ+32����^%a�p�"O��ۓ���W&h���fITЄ�q"O@���.Q�bͮR����1���"O�ip��%b%j ;ѫC�Bꀘ��"O6�2�ǐ83��hyc-P�>Bt,��"O&\R�j+����r�D�<9$���"OB�9��F!WI�(��6(�r��"O���a���:&n�30ЮQ:�"Oz} �K[���!@�MLM��`A"O���C��T��F�. 
�"O�t���<
����,I���"OFLz�i�#M�� ��aK8���q"OhtC�D�	�d����I��;�"O�|0��#��\r��پ5�C"Ol��b�߆@�(5s��Ap�z�"O&�����)͎��(��djd�"�"O�{R�C�T�����ǉ� z����"O
�y��FM�sԯ��E�ƑH�"OȽ+�)R/k�Ak���L,�cF"O6�(s'�:-��I�I�.�|� "O��r��[�����ΏM�v@$"OzS珋=��xj��k�d%"O���N<��xi��ў�\ �"O������<5D�UiœN��px�"O�0��" 
pr��R
"�LD�&"O889��GmY��ãH_�$I>�K�"OV9
�O%i��@��m5^�h�"O���Ԍ0jfQ���|�YC"O��oA�duf�R׃�}�iig"OR����j��I�
=UxV�9�"O֠�1!�g�8U�,�5²t�"Of����="<�%��e�����"OP,�`N
�
(����ß������"O����PȀ!��L�f�h�#2"OT�C��`vb=p��À[�M)B"OTY���(-��2g'�nZ�!�"O����A�@v��1�M!�x�0"O�h;7�>jT��g
:�:}���'�1O�a��i¨V.���H��}z�x"O���N4h�]��<2e.��""Oh8P�U/T&����m.nر�"OH�J$Fܤ�����}'�%�d"O�����\�Q��H��2���"O��7�?�� �Q5]AJ��U"O,x����(h˵�	�)#�0; "O6 1��U-"d���A�0zfBY3�"O��s#L��qV�� �
�m�v5�"O2�KT�N�r����䁉�" Vرb"O��y�(2���s砃8�<�Ѱ"OD8f!�$>�hp���4|���"OԕP�NV/��RaNN#cwܵ�&"O��0��6/|�s��jqn�*�"Oʐ���&l���Ql�gXI{�"O�5Qp�_;
�*�L�fZ�1+S"O6\zan<��q��&zTR-Z�"O���Si�l�f���B�M)��)v"O�� ��K�e�X�ΰ{�.�:�"O�P+ �3Z���@�Ⱦ��%G"O�%d@�pp����)�"�Ct�'�1O��S�ck0U+�$ŵ3?جh�"O\t�U�G��0D2���=.��G"O��
�%ֹfu�D��8l��z2"O��ZХ\�9+z ��91�ԓ�"O��ʇ������^�i�b��0"O� `�[g�I/������^U�r"OV阃�Y�j��U��*������"O$��MY*;ʡ��'F	�0;E"OxIu��z\�Ӫo��JA"O�Њ'*�L���dhc�u��"O��9�umFɻ��^��n�X�"O���E�v�n�ӳg�A�����"O����b�J����-q����"O�@��k�$���a�Z� n�"O��:��]����
�I޺] a(u"Op�jӨ�#>V��^���'�\�!�Me�	�$E��]��j"d
<j!�d�*'��!��>{���S�L�!���,�6]��^"uT�Q�R�ɐI!�$�[� ����+ Z�`{7B�-�!�f�i�+Ϸno�ls�A�V�!�D�b�y�T� b�qR��þ4�!�$�f�f�cU�C�W��S�*_�x�!�d��+�F��NR�?�j,�ǟ�s�!�$ca��C�}8��c��`�Y{�"Of��m�@l��[��Y��~��1"O�ٱ�X%��t��+��� �"ODQ����#e?^+��s!�G_��!�Y�?)B)BF��N6����!c�!��$1�D4E��$A��yv�V��!�Ď}L&����:$,�9�`FDj!��U?1 �ة��ռ/�]hcE�(`!��,���c��s^��%J\�_�!�D݊�f=0r�	�?<�lЯZ7!F!���IZ��*u�R$!��!c �:�!�²$���!�BC�~ؔq��V�!�Ď�h�J	E�jg�P�p��	v!�T>)�`H5��`�ո�-ߩ^!��E��r�G�'eQ�9��n�#7!�D\$y��apgV?CW$��@�*K�!�E���lI�`r2}�uN��!�V������4mWh ���'5s!�$��tU�C懤V^��3g�?nk!��]����1��<,ON9JR�@�VZ!�d\)a�������`I� �9R!�$H,fǸMs�[
z�0#�ND�RC!�DHA�hq��S��"�#[�(!�A�t<��4hRW l��%��B	!��U-�"� s�C�Y�P�S��� s�!�Ŏ3�\1�0C\�9�l�
A�X�!�!�$Ь'*���/ݴ;ܠze���a�!�%1�b����T�5��������!�BX ���o��q� AXN!���]
$�t������JN�P!�d^ =5\��%`�`0�� ��1z�!��Ėa��E�-� ���!h#}�!���v%A��O�5e��y���S�!�|�l��&ݏ?n���uY�'�!��/ N��:vJ��{_��ؕ
M$Jf!�d��j��9+�_�JK.YR��fD!�$ɨ7��}�4d�(Y��S��+L<!��_�1sգ��Uz�;��
�(!��%[.����Ck@�� G�!!�D�V^��p6kԾgJ��Hf".!��ٞ]��=@clެM�Z�!C���!�d����]��-�>��"<��z2��=��� S�:Z�l���ηM9��4$�;Ƹt�P�YS�<�N=(���K@�,UK���P�<!�&���:Ggέ'w&����K�<� �ỤgF�F�^dX+ʻy��D� "O�]�@�U& IBT�ɉ�l�;F"Oĸsw�
�o	Xe"����� ��"O(�2�O��Od�[�"�R�.�Q"O^�ZvO]t��X��<E�y�"OV!�"@��4�d����ˮJ( ��"O:��T#	��p��%�JVpv	�"Oq��a^S�$����s��*�"Ou�wL�;���T�T5o�hS�"O�;���#M0������x�"O�1��C�	yj�[S"޹h�(��"O�l{7�E%%W�}��!�3{Ҁ�"OX���Ȟnzxc��֤QW�<`!"O`�,-(@.���Sgb�3�y�$U�w9"l���8K�����y�n֧S�q`VHэ8В�y#���yN�MqdEӵ&�5N�8ꂤ�1�y��M-iT�w��+U�4�h��y�M�6�X�C�	,|Ra��ߪ�y� Y9@^��!�ݞ$Q^��c��y�S�OePx)��J�T9���D�y�'�O`V���/� �������y2ǆ�9�b � �T�.�����	�y"懳U(�,�J&n~6p�w���y7z D�7ꗥY�xt�0��yℒ�F�xȷ.T�RM���_��yҭK^�v]AQ�W/J��0
��� �y",W��A7	�5r�X�Ƭ��y�m:.R�97'�kt�����ybn�T�n�#�'_�V;,��%k�0�y2�N_��T)˗Iu�4��ʎ:�yRT�)��2�ܓ@x���χ��yb�؃��T��" ��X��B���y".�3YP�@�'�C�7���+cч�y���h0�D�Td�!)7$ [�J��y&D�Z����V�UC6����y��  ���O�$���"-�*�y��X�e�Ձ�'�pi�ѮX��y�)�*	Z&�S��f�t�a��y2���J���6� P�|Q0�^��ODqbp���(�L4@3���y7�hz�*��0�Nm��"OV�8tᕭ-�vV�CSdM�����Ъ�d8\�s�>E�ܴz��4�HE�X��.3QH܆ȓS~�D#O5bT�4��ށ��d��y���BQ����˓$���`J��+��ёogP4��Ɏ}��l�B�	�h�R2�ЭDz��Qaʋ
 ����7L�*$¡���'��$�bX �(�.�B����(�n���S� �N� �)J�$�2X[#��d��+Fe����VZq1�n܆v� q��|�ڬp���g��E8�ѦK�z<��J��~��Y2m�đdGεB�P�T�yҫ�%s�H(���C��AA��?9w+��@�Z�$OB�Ը�W#�	;@�_^#n�(��.q��%���S���B'��Q(�)�&O
�*`y�n]�YB|!n�i��h��3��$+�K�!=�E����e�?Q��B�lLu1�"G}\������F���o��|E���^��y�*K�7��yp���G�hm{��-��h9�ބq缵1d.��?����O�\hg�*<��8����ڝ�p"Or�P!��?~b��*[~�н�7�'��a��T����gϝ
~2ax$W�țC��&M�ܝ1V.���=��M��`� Y��	�T��y�"	�[�T���[*[I&	����xߡ'�h�Zu�;9v<�d���OȘ��a�GGV���j���O���ҵB�Kv�|���TK H� �'�T�H�eU�%ۀh�׬Mˠ]b��&XZ�a��ȗ}����S��yb�_�W��q�ۯqa.H�	��y
� �Dx���=#�|��O';3
l��O2�1E��%y0Ɂq@+,O�}ے��LA�YAGH܊}!�a��'�F�S�I?nY�	%$A�aw�9r��*7e*��P�Zh<A �_.����@êVA��&�u�'!
���ET�O7պ�ǘg.� #�M�3��Q��'a�;�@V-	]�0�2�##)py��'��)�oC�_�$��AJ��4/N0�'��pӄ�]�Z�rF��>� ��'���bK�4C���q�MZ�1����'A�x �G�V�FE*��e� ���'�j=��n�#9Av��w#�*]��$�
�'���g��o���u�T�<�0��	�'J�hI���'b{��yE�O�>���	�'Sn� �F�5i�4J�c�(2��Q9�',�P�b�!��&�!����'��)�Pτr�d�@�n��+��'܈�v�6p�i�c�7�@9��'<�� �_�& ��N'�Q��'!L9i�#�\�t���aT`�-��'��P�F^.D Z���H�cz���'G�H����in4yQ�G�X�"��
�'� Pei]9m�Y���ޞ+�64�	�'���━՞4�pC�q5("	�'y�(ZS�هe؄	��e��X��'��� 'h��:<�-pG�D�Y�>��'�n��p�يVa��xp�GU���
�'��T�UNR>MF����??[z�!
�'�xl0&
R�r���1I��d����'�x8�[�e=r����(����'�`���f�=�fl�Vi��}q\��'���ia��r��$�%�A���q�'�vȣ�$O�t�%�T	 ȅ�'^����-�7�UC�
�8V��H��'�<�!�=?9�\PӬ�V���'}P��%f�`|:�OэG^4��'`�;?=eJ����S�$td��
�'��H� &�6�$i'��Hn�
�'Ineq�a�p�I6��?\M��r
�'Lѡ�K��aZ��R�I�0�	�'����Z�4'���$G�(��t2�'^�\�!�	!�%
D�#,� E��'�p������p�'�j�J���'�>y��@�:i$�iH�ˎ�`�$i�'�<����L�_���Z��=*E4T�'����!�3_rЁ �&����'���Ja�	�0����צ_��'�2 �CLl����_�C�HK�'�&����9u��Q�'��E,�;8�d�(#<q0�x�'v� 0P���E�l�3Ś�zm*���'$������|�vl�K���'�4�
�_y��8KƁ�6s��	�'zx1H��6�����CH
��'�HEӑ.���6� �F�$-1�'�J����KH��'�H�<����
�'-�yʒ��0R̚)�R�D�|)	�'Uz�Hp��b���!��D�Ԍ��'J؅��d��X�L5���<�X���'�� ���{Ӯ�	IV�{OP@�
�'�@�*��++|�hpd�/i&L�	�'zH�;ׁ���2�*[�k����	�'��1�7H��4��;Fǉ�ȭB�'�`i�e�	�ʸ��
���F�y�h�N72�Q��/"��� 1@�9�y
� ����J˺\^���@T-L	�ru"O�\уlV�h:@i��$N�j�$Y"O�,�f�d|B$�u	.` %"O�d�E␑g��c��/��DZ�"O� A��D��4Y���G��XS"O�9�cĿwԨ�U��W��*@"O�-"Wd@^��V�7i���0"O��1�._� r�}����.P0�"�"O
�(�ɖ"CH�a36� 4h��"O�x�%JD�V����J6P9~II"O����@^o��Qa���(%k�"O�81��V�c=��h�h�uH�p)v"O��%���%�:}B7�]�	P��ٕ"Oθ�TNL)c�R%8���i9,��"O�= e�'\".LJvO�A �H�"O�ћT��U*�i�O	w��Q$"O�9�d���P`ΐ�t���[��O�,�%�&�)�'G��-q'�K�\t�HS��]82Ƅ	��?�-�͉F��9��[�tw���'�lB�Cw���2H(��#K�3d6��;v�*�O�kť�@�]r�YP<hueJ9{0B�"O�EY�2�H��TC��+�&��I?+��|�3Q�E�3EE�6�4���^{�B��������-�ZV��>>���
�JD�r��ӘW�8i����0:,��w�B'_�C䉜5���zB)-1�I��CA�p�S_l��v�%\O�����҈kKؙ��W�D.80
��'�����i���9��X9�ԉi�
�(ł��'�v��u�ʡQ4�c�'G	x�\��	�'W���Â�%JB�hH�c�Cظ���'%|�rFX�J�Y�IZE=T��'��@��ҷN�t��B��r�l���WMf]C�G�|`A�D\'u���q*������^w4��ę��
�ȓ.#B����jn�U+`�q��1��V�$9å&+YL�(5��.ܢ��ȓ�"�`ᆎA�тR�I��p��@Ѥ Q.
G��E�1�<���p�<����Lw�<lҵ)ϭ�t<�ȓ	��`✙??�2�ʈ�*��I�ȓ��(0Q�� FS6�e�S�]`B���_��}�-<hx��@EӺ'-�$�ȓ
���*&��<�Bt�b�	1_E��ȓ.8=�ȋ1vt�]PBl4����1�1@w �Wy�����7������6�R5;�C0"��<�����
�z��)�S�:��Q�EU�$�ȓS���SF\�xv9�� <�:%�ȓ)��x�V���?�Ȩv�� -�%�ȓ]��0gd�I�G���V�J�ȓ1ޔ��"�[��0,1��	��-D��B�ӝQ��D�I��,�Ǣ+D��Beb<2ЀcK�1��kQ�%D�,���@q@�Ժ#�R:Tሁ�p�#D���ݩC6�8%&�3�|���-D���P'@Eh]ʷM�~�8�b�7D��e��m\�*G�<J_J\2�E2D�xS�
`n-�G�ہ6��[0D�`�9&��|�%%ն�����/D�T@���M��)c� 2�p!Bc�*D�H��/Ȍa�v�IW-P��*
r�<D�8@�\�R��hU;t��sB?D���!⏴-2t}`WQ���� �g9D��R��	,�rT�K�1L̴ѩ�B6D�� ���\�%P��C���
�(�a3"Oڼ0G��	�����B��@`"O�9�0y�����YZj�h��"O2`� �A!;��y��O��(J�HS�"O��V�4gԄ�tN�8%
5Hc"O,����{p�X� ��=v�e�D"OJ£ �0��+u.�)hk�m��"O@S2#�)YG�<��E�!�-�e"OT)���9Pr��'Ľ�IqC"O�����QDj����rI��ɒ�+D��p���%�@���1eg)D�g ��qf\h!G\�<�.��3D��A��Dm,��:��\�Vަ���'D�p���[�]64��4]8o[��p�a$D��em�K�) 2��!�D�$D�h��mR��B�˒,$V	�K@4D��{ ���I2 ��4T�90e0D�@k�FF�z��mY�X�؉��=D� Q�����q�e�80��� ��,D����eΫDF&�9rbƈV� ��<D�l���$Hxqq�N:j\�`� D�������T�L�c�C<N4�S�%D�|���X�&a�s�/�"-�q!9D����ꘕZV� F�ܐ<��a1!6D�p`���.�嘗�=���S�5D���DI�;
�nū&��3`��D��7D�L�E�&!�|�W�X#мM{6d3D����`�d���C!�W�4���t*O�I�B	�v5DઃP�M�\p7"O����M��PZ ���Pq(ɔ"O�q���,H�8X��XiR��'�>�86e��٣F$�2)��-�	�'�\�RI��k�	RC:/lV��'̹2�/C�vԚ""�'�v��'�
h��$�0I^��"�(`Fl�`�'@H��&-\R�r�E�=YR��
�'�Hq*a)M�~yT,���F�E&P5C�'��aHe�h���_�,�ș��'�(A�V@�kQ�yz�n]�'�L1�'7:$�㏐�bA��j2GȌo_��i�'� S�*.����'+O�M��'�%y4˒�o�c� �K�e��'*��G�R�!�����5ll���'r�qa1B�/�̵[!�H�]7�,�
�'ࢁa'�W�j�R'L�U��(+�'
(�5���Vy+�T$s��ġ�'X�M�E��p	������{�
���'��`80���+&�L� ��t*0�'�� ��I
$�F�rpf�%m8(��'�=���IHx�'�D�r[���'�^��p�C�F<)g���|����'����C	HR�a�*�k<����'�x�*7�	�|\,5���aW��h
�'�)hr�H�q������A��'>��ͭ(��M1A(_>y{V�
	�'��r����^D�����&r�&}��'�&@�L�
a�`pf�v�,��'��]��Z�W�QX 犪9t(�b�'N�g�Q#$~� [7�6Є�S�'*2�B�a���Ł	%{�&Qh�'m��k���'�z�;�G�� {6��'�`�R%��n�2�1��G�ypN�x�'� ���@�e�:���ڋ{*���'O5��\PG~����1q
h9��� .�C�d�	{����I��{� �1"O��I��^�R��,X�F�9Ed���S"O�U��Q6D��Ik���Yd��"O�t`枹�
�ȃ�N���A�"O.� ��/�F=`��<��MA"O��AkY;������ j��v"O�Y1�=�V�$$�Q�q2�"Oh4[�k�8]��e��̓�E���;e"O��a�`�"9�9��g�H��"O,ic��!��㱋�<5B��
"Op�p���%^�m�djڴC� 9��"O(Ⱡ�1��|�@�9uʮ�c�"O��p�M���|c�@51��)�"O��rP,D$j��m#� �+h����"O���`�%�HA1�k���u"O���R�Ik���3�C�;�\D�"O��8�j M@X��wI_�)�`	2B"O�$%k�K"l�����,рA�"OH��_zzܔ��	>Or��R"O��8q!2T���8��7(�h;�"O<(�K��x�p10�@�­��0"Ov�q���W���C�� S��B"O��h��0q�@8������PA"OY�B�]��-`�,J�,���H4D�,��dH�i�s0�2"��d�(D�����Ѐ_\�ೕ��<�:|���$D�Tb��5eY�ye�P�_1(���d1D����d\_0x�d�5
 � J.D�����A�z�Rpl4�3� D�Ts�d���v pcG)V!JA��2D�����V8@\[�I��hy3D��R�� P��UAH,($Hɸb?D��തD�`��!��eaH3D���(�;R|�9 ���,��|fD7D����G�ĩ@��k�:��'�b}�tJ��7a��)6��e�pe��'��0����
֔���i��t��'��@!.B�a�uaʌ�X����'��S�đ9Ϥ��`ȩC"��h�'���G��3E�
��-�	�!�	�'�xe�E��rw�
ƤY���'͸�c�n��Q�z,Z�$R,\hz���'�"5තC�o��ps�E�I �Iz�'vР%.X�n����d�׫@~<a��'8:�*M%c^� c�΃�@*"1q�'��
v�G�"�*4k0�Ԯ8�.��'G���J�	��diu�	7` ��'�l��$��7BV�хhV,)���'�j��"O'�4���Ā�'�	�	�'�Kf�[�2A�q��"ax��H�'C��VB| fѻ��[�y	�'Kp`p҅�1U���S���e*�	�'�9 0/L#H IU��(
p�	�'z�-��Ǝ[��TQ�)�,����'�a��/E�\F���Ćڇ��$c�'�HK�nW�=��s�膨-:@�'@|�1C�^n|���V�Q�X9��'�ʸӶ%]"0���BBBe���p�'���3��N�Go|�	�Ӫ@shI��'�Z��҉β*@-��!H^��'�n��t	]�5P�����s\0�
�'+���@N�qX�Q���&e ��
�'��5���,Eyt �o��ZMC	�'�P���W�hb#i�	"���� �y:U�Z�F�>��V�+%'�y�"O����MS�+��-�m�8�j���"O�Ȫǣ�+i��j$�z�ı�"O�-+�
8�c���s��(�"O��ɐj�\��m3� �,E���2D"O�\rE��랈ր�"�����"O�lp5��1u$�����.,q"O(!�*�26��³�ŵQ��y��"O�d�^6�xDуKدz��q"OB�
#�ř`' �3'J��
.}1`"O�,H�D�/��YS�E7--���"OX�
ThV�H�R��H��履"OfS6�G����`ǫ3@v0)%"Od-����<]�A��+a~�"O�5�P���6��S
'l*���"O���wcR&(����C*,.Y�1�V"Oh-KU���|�1�,�/Иy�"O,ţ��I�.�t1��d Bx��"O�e9��R`�K�Lכ"��c�"O�����M#B���"@��X�XT��"O��pvI�=0��2cOU.F���I`"OR� �Y�d�h��P�F�c "O��2nD'z�(iH�� �3u��8u"O6��AQ �$���nڃ���""O���PP3v,��֌E�����"O�H�L=r�h�J��`�{�"O�A�Q�Z�^'�Ub���F�.qS5"O�ERp
�������m��.�h�f"OH��R�1ݰx1�`���D"OJ����:0�X�  �P�V�>��`"O�TsvH�."tl<��h�Q�q[�"O
����҈�zYcG��=_��1�"O�����(�6��% xu�ݣb"O�D�B-�<��YN��\��\h�"O�(���e�`�����Hu��"O(�RB���x�t�ӭʁRvx�R"O��2���V�*U� ���w\8��'��8q��	1�z�iC!$�ܬ��'lf|�%Y�m�l}*��=���'
�xA�� ���J���r0��j�"O�83(j��u��T�S*&Y��"Op(ӅL�oG��8��ϕ~2��"O��!クVp�h��NRZ�:��"O����Ԕ|n���fE�N)pԑ�"O@�YD�ƑHI�`��(T*N�c"OB�24*P}�.-
�G��ix ��"O�z�i=|��s��A�{�J�ʥ"O��rH�' ��A�օ_U|��Cf"Om��'��9���T��)�BL��"O�<s����E�G�A��Ӷ"OT�;`S=�"�s�e�_~8��R"O
���	/	^��G�@e��X�"O��h��G�G�85��Im�Ti�v"O����F^�1`�&�]�|��"O�ڄLU g���ѧ)F%^��"O4-�,��2 T!C�j�(��"O�h[ ̑�a�xѨ#�QO�1HV"O��$��Z�I�P��,�1�"O�L��F5]��C&ɖa�\�q"O�L�$�j�l��b�\/3�Ԁ�1"O�ep�l]�^�Z�	䀊�*�,�Y�"O2��c�7/�,����$i2�"O� z��2m�d��чF�X��E8v"OFu� ��		�<l�U�s$�Eq"O� Ƞ��a��5�R�`�$�f2Q;�"OdT��ў*�<U�g#K9>g�#"O.��s�G�c�.��%LЉ
g����"O��e� �6������{!|SR"O����N�o8L�#�	�O0I���'���2R�K��Ԃ�GҷĬ�0�	�+��H��j�k$�ȓ6O�=���D�_u�l0�X~Ņȓ<��x��M$�N�����\��Ex����0|� C�֑:P�		e
�u��O_�I�e�q���)H��C��ϊd&R51�&�`��u}T ;���a�S�O�
���lE�@ T0�m�����42��� (@B�S�O��(���vc�h1��\�	�f��hPRѪ�|��S
#wd@�0e�6	$���Fj�^��Dx�k�\��� �0P��@'.�96tP�y��@9}3!�]�dE*t���QF��,�"埓�Py�/K����2n��b�pɑ�^��y�#G�P�
9��#�pW�г`��yb��b`5`!-��d��cҸ�yr���'8��� �~&���$M'��'��zB*܋Ť���b]�&�J"�-�yB@.rI� W�%����bR1�yR	�I�9{�#?�^d��G
�yr�M�T�la�CH��D�׎���y2�ۆ�t5���[�X��$w�J��y2�^@��x�&��#H]㵧^��y��J�J,��r�����H��B����y�'],��P#����a:%.)Y[�ȓ� 2D�U3��j�e��,�ṗȓ3L
,�QBQ%s�\���emV��ȓ�02�ž`h������cG��ȓV[Q9S�� ���*��)�BQ��OJ��Ză)u�:t:&)�� {����6:�R�ǖ.y\
�$�{�HԆȓ{�(�M9�=x#�g�ze��Rv�Hq,�b�\�S?+�l�ȓ3����ӕ<4|����/=��ȓy�p�R�a�# ?Lh��2k�"���wT�%[�(�.~�3�E�9&��ȓ<n����Ŗj��i[T@(KI���'��<��ޮ6�آ��ms�h�ȓ65�IH4�ʴE�� SoX+�~5��J��At��|�X�`�.�]\ڥ��7�>�� b��|���xЦ4�ȓX�|��kٗMVD�cΏ�n�xD�ȓ/�$9�3�G�i��y��L�H���ȓ'�6��T�xE���b���Ĕ(��P��Xaꝳ�|<i�l��,l���ȓ!X݋e�)`�\I�f� ^~�$� 9�t,�<�����&Co\��͜@P j=��u(Ѩ"'�T\��K�p�b@�V�uF���� L�P�ʼ�ȓL���#��yP^p#��E3
!�$�1�^��$BZ���X�L�S�!�D˚vK���%�L�8���[gG'!�d�S�T��ʘ'�މ�"$j*!�č.F;��%`1$��!��#�?E�!�\6Ѷ�bb��4n� ��(�Y�!�d�$5��a�AT�?WR;���=�!�b��m��G�T�R�����ms!�߿�
5�� �1���ޏ a!��02b ��DͶ[t����^J!�d
dN,��#K��	X����,SJ!��0N�p�W��AAС�G�H�bc!�$�:F�>M��G@�	Q��ѹ/a!�� D���[�M���VD�	�m`�"O���`I�ukB��b��M� z�"Ox��"b_0�Δ��@U�&����"O�uC�&�_<"�h7����"O�U����z>��0ӊe�~�k�"OVX��L�8H�X��-�2p4��v"OA(ƄWp�d�H�
E_��:�"O*PhfBZ�]6���_$H��prS"OtH�s�U�P��MaӌE�J|C&"O�Z�{%~bs�ג	�@	�"O��J�Ĉ�u��{c��q��1��"Oj`3g!�$W�-a+�+A�>Lz�"O&��A�ƙ.�R�����&^ir8{�"O�#"ī[�Xv�Dki`��"O>ـ�Đ~p��S���N����u"O���Yzp���0��;�^�{U"O�m�1C�5�$�fR+V��z'"O��'Xyt�񰤯���)��"O����mн�Rh��N	�~���#�"O���b��Ol�Q-E�U���K�"Ozy�R
C�M{*�p����Y!�"O���V�B�K�>P(�L[m~H��"O�<��)�� �v����y����"O�p�#i/a��(p
�=�`Y�g"O�[�+D�5QrܣRDH�a�B�х"OtI��gJ�W������D�z���"O�lh��N�,��$rq���d9�"O���	 	�,\��c�3qu4��"O̋2,�'2�QB�Did�5�c"O���R�.c
�g2[\�zW"O�C�/^;4�A�r���*G�u4"O0��ݫU�6��'P�8"^dI@"O�-B��́s�Ьs�b�	c�q�"O2�!�щKtv�R#��ߪ\��"O�db6�ކ+i����V'2Һ�I�*OD]qTF¢k--&���N�%3�'3ʔ���=P��;ĥԷE����	�'Z��褯Djz��Y�őrj%k
�'�͛�/�<�"���ă[w����'Ӹ�Cő'�u*���-~/�Y�'/�X��S�ɒ�#�O%?S�X�
�' �Q&M	�D����: ״1��'w�%���Q,	�LiP0DJ%v����'2�+u$��&���/Ե=�v�Z"O$����.R��r0�L�d��"O�����Cu�u�Ӎ�-��2"O�Y�f��9�PRoD�y���$"O���ֆ�	( ������by2`JB"O0��O�/4�֩��`��q�t��"O��G�ԥ,��I��E}pB��"O~���k�>|��@{&��f�R�C"O~!�B�ȃA���ČNo8`Q��"O���L�~Nm��K�$'4�;�"O�� A"�dƲ�+F�ܙ&
$��B"OƼ�0a �m��Ki�87�j��p"OxM�1�O�
V��	W'�K�%��"O9 �nN�5.bͱ3���&U�"OP������䵊p�V�Dű"OrE�6�<���cǈA���x4"O��bd��
r�^QX�čG���e"Ot�	eB׆&������L����"O �����
&���֭ P64�H�"OLpDO@�$)Q���}�)[�"OI����ZB$�!�;XiKD"O� �X���M!Y�0)���m �ң"O����AM4�ID���F#,3�"O���)E< �q��SA�,���"O���$իA�θ�0EF3@��"O���i�$y|�� %Z��I6"O�����V�2A�b�bS����"O>�!�ba�V�� '���G"O4�RҮ@+2�����OD>M[n|
@"O8�DhާVV�P�ߛeW� �E"O С��^�(�����G��r�F�J�"Ox�x���H\Q��E[)8~���E"Oй��D�	�,�C��*s4�"O��� bA�P��(Q�bNV�x+�"OV��šܟ>��(����0ވ��"OƸp���vL�xB�홃Pf�i*�"O���`F�0\�nq�ĭ���@M��"OFYZ��X=]I���̉?"�i*'"O��p �WX-0�K�lj���f"OJ����<,	
c���ZfX)�"OxUړI��y`"�c�A0�V"Od͡�AG0Y�8���ˋi+��3"O���+��:�TٸD!�q'�a�7"Ojd@��j��`�g��+)C�l!"O�q�@� �d�@(0Ӥ<��"Oj U�2p��pR��lꐩK�"O^V��j�9�Ř5*����F�<�pC��;�� ����d߾yX�fB�<!��ۼ[D;��0c���Y��Jh�<q�B�p�p�����|Tȍ�C�J�<��b|�1�aj٨]�Bya��~�<��G+W�*��@(\�Q��ݠ�M\{�<V[�.��H@K��S��8�6w�<!�J;N��mP�"�a�y���w�<���N�!R�ՠ&� i����Y�<���ڰ2hz�!�kϽCa��p�YS�<���i��a�EB�T�|�A�a�i�<鴢ݵ
��T��`H|;ZdI�d�<�eR�'��bFOJ�Il�����E`�<�b�N�Dxr�i��(���3q�Z�<A4���D��dևݾU��e�Y�<3)[<i߼L�Ь?V6��7#�N�<�����ah�k>5�-Bb�r�<AV�G9<DkW���B`��_v�<�S�� "�:���L��I�G�t�<��lU&^V���b�)eG4���@Z�<��g{^0Q� ��"D@�Z�<y��D�q1FMZ�&�8*�<��� Q�<��I�
��)ZwJ��q��س@a�L�<�aD�;����F�|^N�%c�S�<�e���s����PD�p!aP%N�<���+K�z٪�eU*H6�D���S�<Aլ�9!�&�ۄ�$b%\Ȓ�mg�<���C2zcV�#�G�.TB�%�X�<Q��3��jR���p#�Y�<a�pI�Ƃ�NOV�@Wn��o2ꔅ�|�Z���GS��DW/I$�Ȕ��/�!P��2!{bT𤀎��*���6��A��8%8b� ��Y2�.ć�-�ҥ
�CZl"-�bߩZ�܆ȓ%��rw͡��Y��
�t;�8�ȓ+.��
S!Ŋ�h��F.���ȓ��1z��L�cu\�g�^	?��@��2�a��e@������D�HX<�ȓ6����+n���p&"]�c�fE��S�? �xj�.��Y� ��c?u�zl�s"O�yQ%jG�4T1!H�A�2�ZS"O�K4,C?v�#���($���E"O��RD�9U�>���8��4(�"OĄr����r�j|Е�ѯ7�0l�D"O�E�'�ʢJ?(Qb3잯���i"O�@c�8R~<� vh�/4�2ݑ�"O����$� ,���G��@�ތ��"O��I�	5\{��&�v��ұ"O(Y��z 0�HQ
}܌r�"O�("r�[wb2�)�T;�\�#�"O>8��F�hI��m#yTxX%"O*kUn�	%>P���j��/-��e"O�8�v��>{E�HBg)�
L����"O�`Z��׎M�H QU�:���1%"O<,�#,�5x��(��-�5"Or��æ���Ƙ�P�(l����"ONy3'��&Y���$	O�4���ʒ"O�܂�߇T&�@Qq�ݴQ|�(c"O����O�h�؉�]�)o൱�"O4D��Dڱ4h\ !ߋ!ix�p"ODx�2��22 ~8�R�VU�[�"O���Ф��7���`��I��l��"O��"S�3.|=���-52���"O�<5kR�XtL��ua	�~4p3�"O,{���)���sG�H��Ԉ�"O�� ¬*X�s�eӻ5+����"O`�0���X8P0Їg�x N��"O҈�tB�8>� �C'����p�D"O&�JRJ�/p�ܻ�5�4�A6"O4�e拘%��PBէ0��ɋf"OR����hl���fd�x���"O��!���F�=�&�����zV"OZ��F�h�@���-I$�+��'O���i�4�S1�Z$}��)UD��3��¥O>��d�O��D�O6ز0��O����O�8�F��� RN��L^@�Hs��Z�)��H(/����Ɏ}���p4A��K@BL����b�Zn�:"��'#/*Hl5�l(���P���8���06�.�p�Tʎ�Q�������M�������O���'J��᳅�ь��(�w,Ԕ]�����?�
�*�4�H�K��)�� �pc�N?�2�L�?[�FS�$��Ř�u��'�V?��AL�l����*�g�X�áC�l�&�B���?y��0O�8[�o�?Tl �hP�l�Ό��g�V�� *�ED{��H4�r�����g�{�'?�d*�I�}@aυ�I�z%��'c���h���0OJh n�0`l�`eS�'�R0Q�8�f.x�~�d�~��
	)����ЛR��l�E��0+�B�4�r"=Q#!ϿJ[�x�%�M��^�iQ�B8�X�ٴZ"�V�i�rQy2M��4�I5�S/`�TL[�'��0�ɦ�BZ���;�M�L<���/�u /I>6���d+�p`�ǓO�`*�i�����(4"�q����I���Ͽ�t�NM�Y[6%��YZZ=��G�Φ��Se� ]��К��F#py��Bǁ
JHDʕkʥ���s�����h��������0��1�M+�ڟ2ߴi���&"|n��-j�+��ߦ������߬$>��X��?!(O��d+�IR}S�H��,�@�ښ_�ɹ��7�(O�o�6�M�Ke���'f�Թ�04��"[T``� �H>�4�Cǟ��	(S�N��F��֟�������	�u��'2��!�0l�2�L@�����/��=w�@H�!� �x�������n��b�Ν#�'�r����d���ڬNR�<"�	��|0x���Z;�l�;4%{��G�P��8�5�]���L;0��"��1�U�n�T��p����k��$��Iݟp�'����)G<�<��t犦U��ێ{2�'�$�����r����fH#Rj.0�5����ܴ���|b�'��D�a����L^�R�N��H�P2V�u��]�����O(�d�O�P��,�O���OT�e�	��*ueQ�'MXa� �8|@�sV�̉�����Sz~��J�P�Q� ���"18Q��	��QQ8�%���	^����-�@ ��h���3g�NgQ� �tF�O�M F�Î2ў��˪!��0�$<l�� �'*��T>��`p�:,��`�
W�I�, D�
S�л6T��B4�U�@�	P�ߠ�?նi)�6��<y���&Fe�F�'�rT?�+ j2.��q�v�7(WT�災\������?��#�`�����O�g�? �t�R�P�	3(��E"��O��9��� -��P��M-zc?�J'Ú*h�ɁV�B����j(0�B�h��	��M�&��\�"(�ر7��~u䅫ݿ9���-|O��j�� �/�qN��� �~�0��� �M���i��v��;V u�u��6�����J�2��Iן���^��[�I��� � @�?2ӧH�>X�H��dѷ�RJ��c�'��5o�,��"<�{�_�zA��A�M�(�ÁM�|��ć�N| ��#���x�R�C6�4���ZMrhS��\=�̊t�ߚs������IU���$���_HW��ȓaF�� 
�-[ށ���B��M�ȓ�(BabV9Y��+�&�A%�؆ȓw����_�&�¼C�L׷Q���z u�C��dW����X�F������zD�h��і�� j-F�b<��"` ڕ)�'`�nћ�ύ)+��Ն�)���V��@��H��ӌ�r��]��R��&o�L�(����	�ȓR!�Y!�o�6<�2�Q@l:;�x��ȓ�1��D�f��lѣ��S���ȓ8E�Y����m��a3f��\�ȓn?����@�:[JQ"��޺݇�yz���`
L�zp����-�9�0݇�OOF���tɘ�@��M�%�tч�%b��D��"����/�jD�a�ȓ~�XUg	4]���D�~�)��/��xKDꒅ)Ɩ�1���-W٨��ȓf�±##i�*�2nݑV��T������W͎=tA�]�ṗȓv�8�RG@�:�H�AW-K8�.ՅȓlE8Z���V�z��M�]�&��ȓL�4��Z�
�=���J?~a�ȓ(�pA�b�>Hp����8��I�ȓ���Q0.ؽ"nx���LY'�΄�ȓs@^�Q�'&:�5���ß7p���9:<p�f�2I�i��R�GG>���	�8���-r	�a�''Zd�ȓO44 �Ӛ;�V\{`)D:3�5�ȓ12�����	���2$��6y�І�]Ap<���Ȣ邬�ٲ熝��a�ݒa�#6x\��oޱ%S� �ȓ[�4��FH�+Q����Ƶ#WЇ�ba�{� R�!�@�9��H/�҉��t6 -���)N�!I/�m�b��ȓp�ک@P�>xhh9�D47Ύ���y������1��x���Ԕc ZX��T��ia�X�x�QH=�B9��=ynE��G<.��=b����i�n���_�Ψ���DS�E�0��2ƌ�ȓW��A�X�T�A�I"8,�Ʉȓ0>�]A��1����v�]f��Єȓ4|��cՀG�h�ӑ�T�[�~��ȓp&AS�oņ�&�1�Y�9訄ȓ3-x4��ųy�z08Te!����S�? ,%�$A�]������
|6&�CE"O,h!)�5 ��R��@�M"l�""O�Ń@�6F�bRV���dw��C"O���AE×P�|I�UL�r�  ��"OX|�Ѝ���a���2�ҭ!"O�蘁e\�p(w��;����G"O�����=�����
���p��"Oj5j���=� 9!�JԬa ꁀv"O�MX�M��A�hs�jԹdDb�"O��Ò#�*W��� �j���d�"O��$g	�{-l��a�s�>hu"O�SPi=NY!tɖ�p٦��A"O�X�@@�42�����ݘ]�҈ٕ"O���l�'6<� ��;5��\0!"O�L�q�
�T��JW?	0�@4"Of�!GY)x��ʇ�H?����""O�dC#jG������^�%���1"O������c�������^�Z��"O&��`�H={L��b�N@�P��'�<`��&��x���8d��'� \:Y�y�M������# c�<�v����FY+A�]:X	����ʔy�<)`.G
lRl�"+��Chqc!'�~�<� �@�^Q�z�=/��ы���@�<9S�R-#������ٺDUj��f�<1�P."�������H) I�q�PZ�<AE{�Ț`L[41Wh�)d�KU�<��J��k�E����y�\Tq��w�<y$m]���8��kϙv�R|�U�^�<IT��J��"ܽ%�vD�ef�R�<��*�Vb袰�I�� iQ��V�<!hۆF9��c�ƒ��@Ia�U�<)𢅺g�z̨#��
>���3��{�<��*��-#Q)0���f�v�<	���z̺ԩ� L(& t�G�YL��hO�O�d����2����x�����'�t�ɠ��p���xĦ@�Fu&5
��6O��≁&�urC�̓q` �K"Oҭkd`��6L,���F]��p�Z�'�Fk(�	JX����A*z�Q��ό�?�`�{s#.<O�١�F=���S�x���M����&�V��*=���,D�T� �,~o<�p�.�Z3�$h4�,�	%���S�\?4��l��A1 Pi��K=^��B��wή\ dl��*���	�)�nb|�s�i�'d�𙟌�sR�D��eZ�B�v<H�b%D�,s�&#
F���Re$<���o��[���9ް>���n��T�W%V"[V$ ���X���B-�-��$\|�E§��sR���흀i�!��T�/�� ��S�Ai��25�|mS2�?�)��7}� (�\*|Qb�C$D���5�O�)�e�p�<A� Xz��ןtb���s�X��� F��	ڗ���t�e�`�7D�p fF/�5 HBziړ	j���z���䞾J1��s&�f�`Q��F�a|B�O��	�C����A	v�VA`gƷ]�TC䉪2�x�I 1K����k���b"<��Ov"~��_�$��4PӋ�6h��lc	F�<���� *!XXq��(N�J0jJE�<���L�&�c��)y�`����I�<�$iS�e��	�fڢ-d�\	"�p�<��))W����$�ĴP��cż��ȓw�x��aD[h2���H�ntb��ȓeP�s��'
�J�P��Y�����ȓ+y*%�Zz�	K7Ή�	C�	��S�? ���](|�p��lƬGj��"O��D-��)p��@1k<A�8 p"OL$�eS�a}&UJ$�O2r��"O^����8{�L��Sʊ�D-�5�"O��3�'S�>���$X��Th%"Ob����&���ޡweę�"OT�  �5;;��zB�E2!]*|;�"O6�K�\���ʖFE�p'\��"O"!���>I�.��V�6K<��"OL�&�ƎMC|�3@I=#j��sV"O�$
P�.B�6�8�@�5g\�"OH�wk��w��y�"ϋ:tI��P�"OV\���1 �T����[�<�Jt"O�Ј�n��Y���o�?�Fd�"O�Q�9dN)Sf�[3D^�uw�h���0D��  G�DC�A!zb*��ȓ2W�Kc�S�`���Ǥ֝E�X9��E��xSW�=��R��W�8|��O���3�ķ6� ��m��;S�ԆȓA�A˰&�KP�Qab�b�`��v�&����C�i1X�5�H��ȓz8qۂ�+�hд�2���l���U�F�p���sk�|1����!�D1ע5Ҥ\���q�� ��c�Ġw�C�G�~�[T��
��ȓQ�}��ӏ�V�f�Ӕ)ۺx�ȓjLm3BU^�-P�
�~|����,\p�*	�>�& �7��C�@I��5���'�׍X�Tu���ҳޠ��m��=�Jͨ��<yTe;գ8D���@M˘%7dܐ�  � exG�#D�(#I]�_Bʱ@fd�ـ?D�$�(ƫB���h"-U�|1�t�ҭ9D��249n��hy�E(Z}�6C6D��i�¸'.>�E�����t�3D��"�pz�ؚ��"K:l�C�1D���H �l�8g��m0��s�/D�,jՊB�/��ty�i[�Y��@&&0D�4�&�&'o�t�$m؜UU��3D��@��_�r���-ѹ��a���1D����
ڋ}k�h��c2��	�� 4D��s��F���k$m��"�P�"g�=D�x��eR�/D4$�q���Ac�!Eh<D�P��K���t���Ԛgk��a�L;D�x���Ѻ2�0O��MR2%9D�X�V��?Z�=Rl֬,�\Q��5D��xơ�H�4 `k_(nF8�#��3D��!C��$��=�uě�i��bA�>D�`zG'�0��Ha`����'$1D���éN��A� ��p*U(.D�|ї-��X��Al�@ql��1D���&�td*vM�aN�H����'�~�Y��D�Q��lD�*��2�'�\`$�T,s��eC$�="�'����
���0Y�d,�tz�'��(J�O*3�uB��R�l����'�����
6\ܸ�T�+$���'��T�(�xҘ:���yQ�y;	�'��Q�'�3j���s�ߩl4�p��'�x R���,!�Y���Ѱa}>�+�'e@峗�3N��eB�֫\�̜�
�'�&P�I�6U;�$���3"_�ɓ
�'0p��FJ�:�a1�&F�I�	�'Bh���
�U�C�@3Ij��	��� ��#����4�3�EN��>�`A"Oh����ZW�͑pO�!}�LQ�"O椁�%�G�}�w.K�Hj��zT"OHq4�Ǣk?
��al�?y`d��`"O*Q`�D@<=�B^�NX"��"O�yJ'I�[���6߿wKPi�"O�1�d^=#Kn��d�C#F4�w"O�MJ���-(�����y΁ �"O�e��V�z���n��Q}�t�"OdB2���.��0�r��	Ry�H��"O:QV��"($h�*���__��P�"Oέ!R�]'%�$�Sn�$9}]T"O�̓���
`RjQY@� l�	�"OJ��CLY�*��@�e�nd��jC"ONYXBH��1��� g�	ba��r�"O��AB@-l�2p��T�U�lQr"OL���05r��"�_�?\���"OB=#�8����B��!W4�Z�"O�A#w㞉u�L���d\ �Bx�"O��#�̒�<k�!��C^�3�&�"O8bP���Ѭ�7��?I}��A"OH����E��A@	{M��"O�����T�@��t��a�"vn�(6"ONL ��8q��b !ڄ5YJ ��"O�q)��ȇ+��H%n�r:��""O+�ŖX�VU�䬐�_;�e3bD�p�<���\�|X΀����<Gt�:�"@u�<��˔_@t�*�)E�2�z��� �Z�<I��1Q�BaPc@�bJt I2hO�<q"��bZ����,�CۈȐ��
N�<ل�J'��u�ri9�� g@`�<�q�,   ��n��8ыR�^�De�)ODDzʟH�7?p��tc��:,r%͕&��aC�6�&�'���'3�)�ӈ2�r�H�0�Nl�J��1w��8�iD|�1 l�5ǔ�cP`ǔ��OV9Bu�Y%i��(�ӄ&�`3-Q� &@�sa�\Ę��O�rh�`�U��)}.D���M�4@��(�Z�M �����ON�D�O��|F��h���ty��ܿb���#�� �y-������R6�h�j@��-���by2���:K������H�,�����J�wFheb�'��Iڟ�	ԟ���S��픈j�
��g8b��1Ee�(@�n��A��n��%A���ގ7��U��	oxaBt�Y�F��Jsl'#�]��B�5sJ,��3$7�N�����ǟ��'&̀V�؈`_\M�c�H4���sN>��P1�H���,.'X5*��Pb��t�����?���ќ@~�h�ׯ�a��HQ�h՟��'KJ��!T����O�@s�% "鎀SE��t�Q�d�O���
�bк�9$��,(	l�c��9"�l0�����r��() �ԃ��T� �M~R�43d�ѕGƧ)��i#(��i�ZE��n�>K�.�o�C���)���@r!
�O*�d%�'�y
� ����7\v�E3m���&"O����W�b)��aL�6 �T�	��h�n�c�@Q�$�Y9�!�/��ya�'��X�u�4�Q��H!k	-rƲ�;�OB�~k&���(D���Γ$an$ �a'�~��صl*D�4�d"G/7ÞtYr�ݼLE�D�'D�h��퇕r4�0�@%Q�5�+�3!�6@r��V�ڲ�ܕ���GBA!���.C�>��q&!(h�jsJA�`9�	&'{���DX9 񸨓�3�*0�&J'+!���5�TeB���5�*{!��ٛ찕�KK��d"���(u�!�d±B���f��v88�s��*\�!�A#"�=;&lW9ip(F6.��}�Ǚ��~��F2�i�!�$�P �N�Y��4�ȓ;q)���.RDF�T #�8���I��!_0:00 QCV���ȓx�^��i��N^Ы���Qt���j^���g�(�<���@�>��ȓ8k�@#�Y�����"�>28E{�����4�Җj[J����D�9��=�"O.5�pk�:B�p��O�>=�Z�j�"O$���L���`Cb��T^��"O���"oO�9`�����+��咧"OL�I�NC�7�.���A�#�(�s�"O�͓ -ėm;4Гł!�L�1�'/��"���4#�(�م`;e8њ��=#�N���)��7鑣-�5R%��;e
�ȓuv���T ��n��pK]7.��ȓ~���'ٰe͌,ipƗAl���ȓy�(����� c��x��	�1A�ه�{Pj��D��S�&;�b� ]%���V�3:j4�cg"Rl��:+\x����٫#?¸���$II����;;�H,��̶ 4�5�G�a.�)���X����?�����@Bm�=;Ft��IJ�xK�(BJ��*�l�2�bi3EEݏU��`�0gEM�'#�Q��!�"q���Ї|�N�jc��K޴U�'��Y��iqE6Z�
��p��~�'�l���u��V�>�)�ʲe)c��#E��@6�A�@]�Ie��P��D:����BG�lxb(�O���'���1ƌ�e��dYV.ѩ���*,O$tKdb��a���@�O_��S��'�b*+SD��@��2,����"^�p�BE�^)D��3o�b^:%���i".}IE�T)�1��Uqg��}Iw"��%!ܨ��=O�<�BN\�dH��h@E���@��d��!���8t���?\_��@���Q�Dؐ����hD��	?���Dͦ]�,O�O�ӌ��Ak��/�V�b %�j�\C䉓�jБ��	����x��EvL�=���K�j�(5�˜E�*m�or[��E��ԟl���$'v�Y��Y�����ğX�ɀ�u�'k6�h�f�T�L:�	N}����H_8�d�)�>�Ж�J��3Z�A�	�@ޜ��h�n����'��?��b��m���)��Vu�����-��������em�Į��T��'	@,k���?���ds�ؒ�AS�ܕ	�]����i�G2D�Cs��U�yK�oД��0��O0,Dz�O��Y��XVI̽t���@M�������- ��lA`Z-s+���I������u��'xR6��p���~�VQɂ�*��	�6�Ʊ� ����M�x��I��S%��B,��(Ot�0�"�"c���X���Y'V�ne�W�A�mT����mI=eV�k�ɛJ5ܜA�{��%�?1��{IN� 銱Tn��͕��?����'��>G�RW4�
V�O*p+ B���<A�706�X��բx��YZ��@yr�n��$�<y5b�au�F�����1�.a�5+�"7�H��WF�{�6Abb�'���C�'u�'���2��!���]3S�!�ħ|��_z��x��4Nd���m3����Ώ%oȚ�-�D=,�ȣ@�$+��h��W�L�0p�7�ԥ_KLT`��\�'u�a���?����N�`�X̀T�$D��ɠ��
��D2�O<	���E/d�,(5F̀ s:���'��ʓ}P���3v,�ՠ�"��ݖ'U�i���'t��_�4�O����'�t8k��R0�6�J"+�|d\�P�'Ύ��3��t;�!J/{t4��*��|��>�!���7K舡�U5;�6-��f�|	��M�/ڄͲB��	Kp�(g�Y��H��X��LT 0)�q�������4OJ��1�'������S�? �tz��G&T\����2#N&ȹ�"O�TY���
.�h��r	��BP\t��I��ȟԥHP��n�h���a)0�L�8�c�5{�b�$�O1��K�}5L�i�O��D�O\���O�����h&� Ka�	�L^$����N�Y VP�F�B?#rJ�租�~v$�'��'V���J�3\IBc��::��ɡp����l�@"�2��`�����)H0s�XN��H��A�\�~9���+k(���e�/?I$A�����S�'L�d�� ̊�a�
r:�Tc�_>/!�ē���\����:7�(�RΊ�?G4��|R�����o1<��j��}�@�QB�G7�b ��MD�[� b�O��$�O���O�a>a���Z����+)�e/~}Q� ŏ��Uf��0/2�z��Z���Oޠ�fI+C�ȐCK���v�@«����)�g͍�lYk����EF~�-Q��?�B	�Wb�rV���b\"�ça���?ٌ�$3����9���o���i͞z-��Q�'�@�`Ɓ�J����D5��=�,OԠo��ܕ'q�d�#.�~����d�ү�6q+�@ؒ_�d�1GB��?)��X4�?���?ydm�2SR���F� >>Z��A��D&�4U�I���"w��!��D1��OhX�@G%y�Y��B�J�˧x�j�
�B�O�l���Y����E|bT-�?���O{���gl�{�d6����@W�ԇ���	=�u�T���a��f_-!�����RyB�\�L]�o�#\і��E&��d�On�d�O���OZ�'�?!�O�x��M�6$��'�mr p9+O��!g�ĕL�'�V���DI���
�`��!�����E��'�F��	w��f��ɈE���pN=TS�y���g��Ը���I�/�b�D�O����O���)D��9���z�g��&%�M;�/J֦�	:ବ�	�<�B��rnz�=��OX�Nڐeq��H�H�Js�0��%Ѫ�	��?�4gH��yұ���d�O����O6�Brx�� {P�+ď^(W,ih0��O`�$0@����r�H� �?7��P���'J�Z��F�N�H�tH��7�����'lfX����?I#��*���T��Ox�)�Ҡ��@�Z����<y���V�[矘�UJ�O��$U)m8�������?7�[�<䔝�V�&'�L����*�*���Φ�Γ{���	�ّ�<���?���YY�y��i���6��H �ŲMG�q��'�&����?qv����p�tK' ��?�mZ<A�|4��	lU��S-��q`$MzB�G��M#��'b�Ő��?yv���Sܟ����A��ѣF�K</��a*�p�����4y�tݚ�'B�}�b�i]�6�����D�Пd�g�O�QcEmԿDv�{ ` �Y�8LC")�Φ��g(���'V8��y����By��Q���h�=L{��I��\51���"OxA@T�W�zB�0MH �1Z�i�"�'1�'<맯?Q���ih���jF�`����cѼ ��<sܴ�?A��?I���?)���?����?	�O���ħ�'a�)���B�r��Iݴ�?�*OB��O���O���|Z�#\�H<�4�A
�1��n��,���[�l��͟`ь�L<��$�GB���&�P({( �C��i}��'��� V��Y��p4�B.m1�H1H<�	���c�*އb��*�Nݰy�D~����?1r�"�#h��<��
�59P�(0�>D���q�ć2�x��@�0�Qb�?D�2��n�|}�rH[�wnF�ڗ�<D�����2f��PJFm�&5�@b�:D���&OU�`I�ۅ�Uv ���8D�T���SzNB�p�g�9���"�:�?a���?���?y�I�'P����ъ������`d�3=���'��'"2�'�Z��'�'� ��1D�0iW���V�Itt�s�v�����O��D�O����O����O����O�hK�A7�r$�ʝܨv�X�y�I韸�	ğ���͟<��џ����"F�o�.$ R�K#����pb���Mc��?���?)��?���?���?���A�[@h�"�C��:i� �^�.{�F�'{�'`��'�r�'kb�'M�H%��]!dA�#7Q4��UD�<;[�6�O ��O���O4�d�O��d�O��X���A�� �4�9RG�R�fm�<���h�������՟���П��"(��3!I��V,Id�!]
� �4�?���?���?���?���?!�&B��E$��4�ؐK�NH��$�i���'��'��'5�'���'���[fEJ/���;F��M��]ZRIbӺ�d�O��$�O\��O���O��d�O�Hk�X��@�q�%nL�X���æA��ߟD��ݟl�Iß��	ß����(��n�~b���o�>0D�qc�.�M����?���?	��?���?��?Y!������Eߪhz����= _�v�����Zy��ӵbD0@Ҧ)�Q�5L*/�8o�H������I�?e��~��iD�n�$7*���	=�,@;d�]�6M֦����d���i�O�1zP�����DŃSД��iY��\q�#���f@b�DH)�f��a�����=�'�y␄@A�Q�5J	GZ���"�?,O�Obam��q=Nb�� �)�@
ٕ� � �G��{*�0�dq}B&y�Dn�<1.��T0 ]�[e�u�R�k�Hh�RV�<i�� 2�}�$#?�'3
p��vBC�y��1�2����\(ʜ�F��,��D�<����h��D�N�15!^���8'$U�Gy�F��7����ߴ�����GĒ	D���6�˜�$�	�B�Bhzӆqm�����R.\��o+?I%a��\HP��^���(`X�3�>��X9q'��Z��=1���d,�:w��)�4&�%s��೤�T�j-.�L����>̘'��l��+��B��5Ό����b��z}�h�L]m�<Q��)E �X${����,E�m�7&�9Ef�ք3/���s*H(S	ͬQy$�1��C.�M#�	�%Ib���k�'1�X���_!X�L �BO� "���5���L}���[!�gj��>/6��F!9�c�h��F�;�)����z�i`�A�kyFtZ����U"������7dC4�]���2�H�pj�{W�RbGט�AȀǀ�1��дcL*/b\���ԁ_B�s/
0t���b�3��,��o�6��<#��!E�]#A��3���Zs��{���E�0��X��.�#���6��,qg��B�jAkЭcD��f����7'J/2�ΔU��'x2�����6MzD�CmN_i "Ǡ�J�H��X9Uj�p��a�:9�D��:��0$���8A��2J�xP��,Z:Qf�*0i�j�y	�)��Mcv+�OԶ$�ĎޟX���)�N�3h���Q�I�}�0-(fn�L���"�-�s�F�xG�хl�ph4H�%D�*%P�/&/Qh��hQ�c$ ��\��1R�ˇ-,�E86f�ZM"�y����ؼ����Ħ��	� 24lŨ&��%a�jI�2�\͋��˟��V��˟���BHf�$�OŔ�1ƨ�&8
�f���01�'�b�'���'H�\H��'=B�'�B�O�r�2&�/�ص�#�`���p�|2�'�RG��b����y�O�ĕ���^X���Rd�Û�Y����?���P����?�(Oz�	�O�/\
N��u�.<���gS�}cN���O�$�1Y��"�����?�����&�j{��X�%��'�B�'�2�'<�t_���O]ʍ�u`��T{�8�D�.R϶���'�h�DhW<�������C�A������E���VB���O����O�1	�e�O����|����yRŒ�`��0�f�҃2�`X�aLN�h��D�<��W��'�?���?f��
1��9Y�#��19�	�1��\��O.*'�Op�D�|�����1j`ջ�K'>9�$̃:�*O,���/O��	؟��	ן��IП,�P.G�~�.�k'�9t��0��O\(V�l<�'���'��|��'��hϋ#����C�G�h�B\)U�#3�6ѻ�%�����O �$�O�ʓ`�Х��O�r�"�)|�p��F�Z)|��-O���O��d�<����?t��q� ��Sy����̡7�y˦fBKy2�'���',�	�$�Ҽ�H|bTnQ]@ �%3f:Ԩҕ�%�?���?i.O��D�O�D8���W�0�e!��4X��p���'8�Y�������ħ�?��w��U �,��:�q�ߠZ��I�����$�Oh��݀kJ1�l��z޹�p�˅>p�Ⴅ�˂MƜ��'��O�ʓ!��%�ÿi����������D�&%L�h%��o��[VB�rB�'���b$�)��g��Z<Ԃ��д�p �w�d~�,��(�7��O,�D�O~��Ba�i>����9G�<0)�lD��DE�7�ݟi�cASy�'wB�Ϙ']��.f����(�&�]�� @Oˬ�M��?i��%� U�b�x�O
��'#N�Kg�԰v92��T��i�Rx��S���	��3E"%���@�I\�q�'c��%)�#ţ0���#7��t�I�FXL�K<�'�?)�����ӊ �$�s�hЃl̪Ġt�O�<XD��O�I9���O��$�O��S�����.�#�l��Ĉ��H��@��@.)�'�2�'PrT�L�������Ӕ3f��Tf,p�l�2���T��c� ��ҟ���_y��ݷ(�T��]?gzBF��-*�<�2c��L������	�D�'���'��S�O2�tk�/�\�� ��%����<����?q��� %p��E$>%k�`��j�؃bj�� ����N۟|�	��|�'m��'�X����N��8�S���El�,I%����?q��?Q,O��0�_`�Ꞔ̻:K�\c�O�r"���&�{ &���uy��'��k ����5,��Q����uZ�k��]^��D�<�W�խ4��]>��I�?�(OƨcF�Q��h'{op���'gB�'P�E��V��'��O ��Q����J�a�]I(��B�'j��(@e|Ӱ��O`���x�'��ӗ)G:�C��R�&4Aw&�Y����YԔѕ'cb�'���y��'���{��U2����-e*���hӂ���O��$B�R�(%��ԟX�	0,��-��C�xH�h�F_2�6̕'V��'M�4q�y�'2�'
�m#���83 ��`��2?\=R�'�r#��O���Ox�ħ<qũ�m�����^"
��Aq$��?���>�.��<����?(O����8Li	�F��B\IP�9KL���g�<A���?9���'r 9h�R���2,d���J�:��]�M��On���O���?�S��&����3��z�D�6��4��E��I����IG�����N
a��ݹ��O#V[Q"	g��P�<!���?�/On���6'*0ʧ�?��M e�&eH�BH43̽Q&/R9�?Y����'��I<f �'��Y���ǷP,Jq@�IS8[�F�����?�-On�$G�@Yd˧�?����� �Mz��O�v\9ŀ͒�,���ı<�\X�'� t���c��(�B٦7gz�ڥ\����~����	�����韘��Xy��� x�u��/�6U�A��!J��	ԟ�
d��*y�b��>	M�a��,�D�������O�|��O����OX��꟢��|"��LP��d��wU(a�
�����b�nL���_m�S�O�b(Z�#��p�Š[&����!)uX��'B�'Y+�T�����I�<��نQy�P� P�kR�k	 �nb������{��럠�I�<ѱ�݈�Vix��zdT��ggB������l��ŕ'�"�'?�$J1x.i�Q��NS�H
E�м]�	��Z��+?	��?�-O:�D��&m ����U� T�S0,�?Oz68A!&�<��?�����'{R�AD�����,�:
]S��%O_�x�fA�����O���<���E�O�p��a�6YDA��.˝?�RY���?���?y�R�'��i���ʽ{~$QC遲6��{��%S[HQq�]����ȟ�'�ң�&0�S��\JP�ɝ)L���?"�V9�F��X�I{���?Yĭ9 ��P�Oڍ�$��/;��Y��O^D�l���'�]��I�m� M�O��'��$���%
`B��h�׃�&]�Ox��_�U�(���ԟV�C�
9H<(�OƔC�&h[�$�	.6Y�	埜�IП���ay����H�p��-n�6%�g��a�џ\�r�Z�t��c��>}��KM;^����)����G�O�\�C�O����Ox������|���"�b RЍ�
�d0K]m<��<"�X'�y�S�O���E��������թ :/���'���'�f4��Z�����	�<��$�J�De`���) �����e�|b����JDe����I�<�Q(��$o�[�Rmv�[qN�������'�2�'�2�$��.���w��vZ�JG	��!��Ɋ%�퓖�"?��?�.O�D23"��dLh��y`3��	@K.��b�<����?�����'w��Ë?~)1 �3o}0K&�ĻtWd��H�����O��$�<�����O��yzEŘ.zv�b�l̜^�U���?����?ى��'���x�H�0�.��L�G��tCD6-�(Q�_���̟�'�l�Ce�S�� �ɷo1<); �PP�Ψ@�������v���?9�C_;O_�`�O��5(F;y!^$�+�3�8���'��P����%h	�O�B�'��4	��y2Ƥ�DK��v �dP�O���Oq���ԟ�I��	�(=��	vؗ��P���Ɂ;\���˟P�IΟ,��Jy҉��A��A��-�y�b=��n4�I��|:B`ʛ%�Db�b?���NelMҔ�&�Dac��'È��D�'���'.��OE�i>���+Ɋ�!�F�r�贛��T)fd���@4�Pf1�)§�?�҈X8W[$]��
r�r�z�kO��?���?1��a�<��-O��OD�Du��CW�[�v�����S��[á��j1O��	gC8���O��D~�tR�#��fPp+A�_z���&F�O��䎸2�0ʓ�?��?A�y"�J?rk�r#�Ło�@�����#���<@x�束(�Iԟ@�''�O
g]�+��Y��a팵;�0	�T��I����	W��?���
�=���D�� ��](V�D+���#�_~��'b[� �I�V@4\ͧ�*ܨ��U����#`P�!����ϟ �	�t�?��� 2T)[���:E�kg+g���5�м.�8���?	���?y����D�=np���O��.H��)�7�mFZmsCE9��$�Op�`���&��H!�	9}+�47��|��BP�_�Z��F��?�����d�Ox�"��|����?��'?�T@`a�X��5S���&I�ѻ���'
�)�3-ݹ�����3F�t�;
\��r��4��Q�����|�
��	ʟ������Ny¸Ĭ�uAZ�"f�����T�#�СY(O���C�0�p5�p�����/�ֽ�7�Z�6O>I�$��L�B���y.R�'H��'���S������+%dO�3?>���l�0O��C����y ���`�y����O���N�kG@yv��;S�*�)q&�O �$�O`�$S� h���|���?��'o۵@�<���+�ʏ.��Z�N��^L�M~B��?y�'z�8p��2F:إh�M�,v}����?��	���O �$�OX��*�oԬ:�\��_T��� �X��p�!������?a�����O�P���<-X�@I7���>�[*бw��<���?�����'uB =�\����E
:*Vd0(L<���@"�����O���<Y��wyX��O�n����Λ:t�jTb�<6����?���?I���'0��0��L� 8�-� V@�06H�EM�8Y������$�'���d���h����Z�nTg�4�ZIw�����Ia��?��	R���H�O�u`��T6��=�V땣P.p���'�BY����yF%�O���'���IW̀���E?jX��(�#~��O����tQf��t�ԟ ����K ����6�C�%nDa^�x��q|������I�x�S_y��S�5���
��]�ؔ�òf )W��I⟄�t�%~[�b��>A�f�Q�X/�U�be�^�j���O�����OJ��O �D����|*��р �x�!J���6cՌ&|�q@C�'�4��6dԮ����V��0K�Q�G�5HJPY��ǣB�:���O�d�Ob\7��<�'�?���y�`E>w)�U�p'�E�q�G`8(���<���V���'�?9���y�A
<{�� `��y-���֣�?���-/OH�$�O��D>�I)�I���;�,�൤�#<�n�� Jmm~��'��[�|��
�%³N�F{�Q��E�6�8�c��fy��'��'��O �Dʀ�8tH��Am~a �GƢE����k�8kq��ǟL��ly��'�ּ��6�v� ��	�m`!��O�ELQ��'�'�r���O�A���n�䑡�T�}��▄�'1����<����?�*OL���\F:�'�?��"��dnDa@ ����
�?!���'%�8'w<}�I��K���86�44�����^%���O$��<q��fZ��*�����O��	(},�	��IޥRO��?����ɔ-�����'0�?���L�L}� �ӵ�%��<f�I۟X
ǎ�ԟ���۟����?	�'f^��c�=D��љ�)^�=���U���,��{Ԉ;�)�C<�+�aT�.�f��E�t���䃀 x�D�O��D�O����<�'�?�%aIF��̀�K�_�hM�'��?�ã��GFJ��<E���'�.������s��]:uJ��YY@���'���'�R	�(-:�i>��	���̓/*�
RN��U*'$ÆS�%�O-�Ʉ5��%?��	ɟx�I,x-Be���CNC��P��<=�xL�Iğ�ˤB	 �M����?���?�dQ?i͓d	�@
%IR􄰐�D��n�8L��/m���kb����ԟ��ן��z�D��vE��D�:z��'��9,����'���'���~�(O����m�ЌrM�z��쪠,ƣ%������O��D�O��$�Oj)�j�Ѧ�A%�-�����K�4�����X�	���ʟ��IzyB�'{��O�d��!-� d.6��D�#(�Ae�'�����1ob�'��S�:�ذ�ߴ�?���l�Θ*�mJ���Ei�,ơy�1[��?���?a(O��dٌ5��O��D�F<�����ב?0�I�TG5�3L�OB�$�O���2�P�m��D�I��H����DC*~�d h��:d�V��	��\�'�]�����'R�����ܴM��y��g�Q&d���/X
�B�'~��V�<�7��Ox���O�������DI�}�43�H�t�`V��Y�˓�?��������L�X��@�B�|,"'���2��L�O�
��������	�?������������kH� 'ϻ`����C������ʟ�'���J�S���/h��5`һ ���H�D��M���?9�klN�����?��?���?��
ÿa߈<ȴ�ށq�&*^�?!�����P/P������On�DؿU,�����.s�5�­ߧ"�"���OD����Ӧ���ٟ����p��0�&��x(a+����,�mhʓc�:����$�O����O����O�m2�$M�a�7CC��v`�L�Ln�ן8�	���	���)�<���h��T`&�	�Lĸ8+DKH2n�4h����<���?)���?����	ˢ9�`lZ�2S� ��A�&�~-�&�	!^di��͟���ڟ�����$�'k"oƓ����U &�B�C�Td�,�ѶDY4�����	����������؛�MS��?�'a��tc~))����8Z �ReM���?A���?�����$�O�%zG>���$�O��Aㅚ"�HYy�B��NT���MP�d��d�O����O�QcE�Xڦ��	֟P�	�?�tO�0L-x�Y~��j�]Ο�	}y��'W�xP�O�B�'R�A��O�t�cϋ(@��117���l���'�b�'�DH�Ѥf���O��D�j�	�O�h�V��-R'���A�<I��d�$���?�(O�I0:�կU%蝹�- 6��Y�mH՟��d_/�Mc���?����*���?1��?!�! v������19�qc���?��������yB�'�8�� ��رð���,���sӴ���O��D�/���i�O��D�O���O�`��m&H�@�0�)5E.ڔ��Of�$�Orl��kD�u�:����)�OJ�D��KY~R��B��)�����*���O��h��A��������ȟpH��8��	[�2�3 ��KS�ɱ��-� ��܅|-.�au5O��$�OF���Op�ļ|��`��Z���`7)�j�m�1M�L�;бir�'*��':�'��D�p�Ү�%P2P��r ��Z\T@5Lʍz��<���?���?�� �1�E�i>��$�	b�%{s����1����?����?1���?�������O�JG8���'	=eL0e�@��|r!�'�O��$�O���O��D�O8p�IѦ��	����C��9n����G�k=8D���ğ���Ꟑ��ky"�'^J(�O��I7A�F��3��#t����s�Өq�M�3��ןD��ޟ���<J�a�۴�?���?Q�'0�&p@w]���q�Q��`V�����?A/O���	-p�˓��4��)[�.
L�L��F�H�A���O����O� r��Ԧ��	ܟ����?�Sڟ��]M��8	�˅=(/,
d�jy��'�
l�X�����O
�� �4��iA��2s������O��c�O֦=��������?���\��ݟ����#����Vy  ���G䟘�*�럀��ry�O��O��M�W�>���7+G.���^>3�6m�O����Oj��3g����d�O����O��d��s���׫�ahnH8�22����O^˓2�P�pO~r���?���$�2 �A��r���!$��y���?A� #k���'��'�b�~2��� ,�0K��`d���ꏯ���CW�@2��p�4�Iܟ(�I��\�	c�t�ȊA0J��@,��&�����T<u�a��tӊ��O$���O���O��I۟Pk��Q�4u��F/YFҶ�ƗzK�	֟����d��ݟd����&a�-�Ms��ˋ04�� ��i�\�*�#�?)��?���?����D�O���;�dxæĜ,Rj�$k�I�Ƙ1���矜�	"�����ҟx�'���c��4�)ܨs����������	B��s�d���OΒOf���Oni��;O����%6�b�j��F�l��<�	Ο��Ilyb)K-B�B���D���Z4n[�P�裗ԓq�̅�&�<�$�O���ߊ=���d+�ԟ�eȧ`��L�F��f#�6Bdr5�'�ɛ[��xش��)�O���L@y����ظrG�g�NA�'R��?9���?�D蝜�?yM>�}�Q�ێ~��7H�J\I���Nꟈ�R���M���?A���E���,G�0ҋ��~Э9N:y���٩���=� ����$!3Eͷ����_
v��mʀ�M[���?A�vq�G�$�O��I,,�AZç\ ��ШQ��-9 �d:���!T����d�OT�ӮO�H���O��RDj��^�~<����O���)�d�I韌�Ip�	�?�)��%P�2兌 4s聕'�6 �'���ܟ��h�
1�8���)��"'�ۃ$�9 i�����?y���䓅?q�&|�$)U [�2u1u(�.bS�i^�?�-O��$�O��d�<	�D3q��D�S#�Ua��_�LrN���W9����O���)���O����f�D��0�����޿pt�a�2��` ��?A��?�(O��*���v�6Qh�)����p|���C�2o��������&������p��
}�$�'�r����h�ԝ2�M%ao�����?9�����_�n,e%>���?Ɂ3��K��h�̈�CdN$�6�AO��ϟ �	�	�	M�?�!�]l>ȋd�;U�ص�)�OX�C��:�i'�ǟ�ӷ���>��i��GM*q$��ˁV�'}RI	�m�ɧ��Q>%�^mچg�/~@�Lu���ٖT�IA�t�ߴ�?��?���r��'��锢d�佃4*��)�&�1j���N�yr�|��I�O��Y�n.
.Ƥ�'(J�31$(����ݦa��؟@��;0��}��']�"��H5���+��X��rP@���O�t7��$?E���I�6��!��)��[Z��kQ�B�>ŸP���誡bY�ē�?�����D�4]�Wa�-]�r�����).��/O`�����O�ʓ�?����?�*O�y��G.N,*=���&b�xh�a��o���>���䓪?���%kR�0t+��
� �䖀2"�	�l��?�(O��D�O6�����@��?	 Cn��gp���M�����1ϲ<!���hO\��� N���G�?��|�"�:z�p��Q^�����O����OD�$�<��@P�O\���2���N��"6��4X^d#R�'"ў����"����ڟ̧%A��E@* +��@�
�A��9�	L�I[y򡙌.�����dw�9�F��_�8��D)K�\7pH��*�IΟTB��埘��W�'p���񎆇�R��sad� ��y"
J��7��|����\���� $S��4P������<���
nz���?1�����,��U/��"m��"��>�R�_�B�'��I�?��'��	2
��PF	�7�H�Qr��-[����?F.̂�e+�)�'�?A�$X�x!�D�˼-7nekDI�|H���'���')&qX`)�4���$�OP5����ꊕY�cͽ�F�	��2�	�#��c����ޟ<�I�]XY�[�rѤ���H3F�}�I՟D�R�ݟ4��v��'d�'W8I�ӥŒ!c�P+Wj�A�NQ�`Z� v�j���?Y���?I.O��x�Ңt�t�W�
�?vH� c�\#S�� &������%����៰8��^�h�ؑ�J:��9�B���%:c�8�I̟P�ILy"a]��|���.%��M`"�H#X%.=Ya)��3�	���a�I��I= �R���kKU(7+[�er����Y��˓�?���?y/O�@�&�K�S $v��P`
�u%1!l�.Hh�I��%� �	��Q3I9���n�B�'�mvl�A�ԄA�����O���<��l�/��O��O�� �S��&8�jŖh9FQ���-�D�OD��\�qO��SN��a�N�^Քst��9	[����<�4��(䛶U>����?�:/O����?(2B��"�����Aj��'2�'E��K����R�oIE���,�ب+ 3O;Ri�<e7��O`��O����a�Ο ��I1]o6�"�@ `�&ᒑ�Z��P)%�S�O��M]�Oކ}�"�ܝ
�hH!'���7�"�'���'^4h��'�2_>����<���V�YC@(���B�5~�-z�c��b�iC'Mw�ןl�	���`����dI3�$�.��h�#D؟����p(|��J<�'�?����$�94dN�g ^_�Ti·.�p}�I5[,jc�����\������	g,@�E��P�F%�?~F}�5 ����Isy��'��'��'��P�͂`4*կP�`؀��4MY�eQ��O�I4MX�ED�^���	�iǊuDX<k$ޓL�DP#��ltᅡK�"���"	F8�P�Q���?����?�K>y���?Q� �$�@*ӥr�ʨ;��"O/Ե���'���'j�'��S�?}���?iu�E,W�YQ�I�,;�%���K&�?�����?9Fɟ�H���sфU7\��!H7b��+���xB�ӆ �&��#2@H����2�'X3����g."?)S��Ym8aa��3���Z���E�'�\�r���}h���DMU�~ܱ�H��x��q�޲*��M��oj�^(j�I�۰���n�!%�nA�n��l�Hd��դ�N�Ai^��ȫ5
�&7 ��3���Gק-�U�B#M</���� ޴BlL	qNS B�l���-�3|�bF�>;������@�Q4��X�X%��P�LZ,(�������?1��?b+B�}�X�I�oT>!���jV��2�$0%�9���&*V�4�ŗ�9�"=�����DA�+~m�q��oj�.ʪH�����L+�т�Aǩ@K�����mm(�O�����'�1O���x(���^JabY�`׈&�zC��1W!����=X\�rVo֣Ma��'rў�S��I1AfH�B@�@�&���H��&5ը *ڴ�?a����f�"���O�7��3��]���|��X�,s#|cs˒�+��H�4���F�y�S���i�"ዱ�:v�����8@ {�4T^^�Y��ʸ!�d�r���So�?7���%�J8jD���ikW�Fu��ƤQ��?������ĝx���(Tz�gN(9�5�"���yb���u��D�Al��+i,E�Q�&�(O@�Ez�O�F�=�����Ȗ5�8�	
"I���D�O�a��'��o���$�O4�d�O�8���?Iڴ-�\K�A��%Ӕ�Ǒi�JL��I�O�����)]ֲ��d��_���DR6V��Cף\��$`4ĕ�to��Z�\R"1@�I�=sc�@4P?#=!4�T>��;�+L�n� �Rt#y}b�~y�	�D{RP� ���,����A<=.�� D�T���#|�B��1y7����I�Q����Sȟ��'����	@Z�X����l�~�R�.� ���h��'x��'��L�@P"�'���@6�4 �#�->�Tآ�.ZO�^�&�[�X��q��5*�l���m�XD��N�=K$����O9uX8�����2��%�6�ߡKv4��䜦2����!h�t|���.FOЄP��%%�(���#����6������w�0��-�B�<1U#��l&��`����B�L0pk
���l����|�'�I�^7M�O����~*T+�`2b�{�$�+?��'W�B��i��'B��'��	K׎�vW�I4��3?�<�T?�ʑ+߉!a����	�p*eA��.�L�u�u� �����ԙ��S(wQ%��S��`Ȣ����j#=��(�������(t}�y���5�쵂D��n�!�Ċ�1\���-Dr�JaP��O<�|r�:}R.��	� 6��Z��`��1q��E's���n��t�	`��#���'ћV�ܜx��,���	)a
�u{r�/z���$�eӮ� �� Ro�������)�s�@]($
^�
H̳�J��d:x�Ѿiq
�@K���J�J��U�c�8���RB�
F��] ��W_H�H`D@��5r��O�9$�"~nZ	�n�0K�
��E�fţ�`C�	,'���񣌮�J��c�E�K&�<�F�i>�lZ i���Ј�0\u�&�^�X���?i���+&��|X��?����?���� ��wD��!����bPгE�>��,c��M��dR
~��EG^�|`�3�tL��c��� �2�Y�G0W�Q�G��͉�FU�� �����	�~�ź�(;G�����֔[t�F]�)�I\؞��3�D����/�2Ȇ�Z�!%D�8�J�6[ȴ��1�Ė�HvO�U����m�	y�4[%��\˲�C�
�=W0E56��-C䟰���D���/�(h����ϧfZ��"��o���R��Tɠ�1 ���%2
�H�ƙ�4 �F��OtI%w��PX��A:A~Tcu��ОBŲ�#��&0�U��+�
 B
��WL�< �����O̅A�܎6���s�
��1�Bo�&�y"+A,ö�������Er�ǂ�y�w",��qE��$��C١�~��h��O<)+�"_Ѧ���ҟ8�O�-��"��/���.щ��� �n�3V ��d�O��$�U�>9��?�����
M��0��Qc��*"5�h�M��F�~@Ez��G�>�(Ie(쬑�� �j[��߷=O��P�`����`�/?�����o�O�D��OW�kC�Z�bK����q к�y�����Is��,�fHI��p>a֚>a�m�g.P�(��r<
��#��e?	��An)�f�'�Y>�kG�͟ �I��#��V�T�]h�Y�-Dh$)0�>Z��iƮ�_�|�� b
�F2\�vk�?1�|�1#�橫Qa��86�¥Q1_01m�BY�,s�͆ev2���B?65"I�d��/iz�avÅ�\c��� U�)/�h#լ&I��@"�4A9��	���S��MC�Ə�Z��@�H�P]3�GU�<	�f�Ow�1Kf����!��Oi��?� �i>�mڳ^Zm�A)R�}�^��D�6|�p=#���?�Rk)Q�0U���?����?qT������� 
(��]�Gw�9�'�V�,��}8��y0"U��C��1�8��r�'g��2�FЀe�6�H!�\�W4��qD@0JơȅM��>Qz��N���(�	 v�y�C�}� L�3픨g�6��OL@賯�O.�nڴ��Y� �	f}be�(,��a��З
vQ�/E�y"�S1�M�dfN> ���%�pF5������dz�Q����4ξA����6y2U�X9<��$�O�d�O� �A�O��$|>eK���;tD])�oK90J���J����Yt�$��|��܆%�`$��h�6��d$bU#Sd}�S+�y�,��i-uE��㉬BV����5' �3���X木����<5pi#�'��u�e*ƕf�J	�B_3�`���'�n5B��7z��� ��1]Lu��':@6M)�d��^=T��'��^?B�a�;���� 	�c�v�a��!6(nt����?9�n�J�[ФH7-� S2V��'fJ����� |��ؒ%�|z�iDzrhϪ�����Θ-q��Ȳ�*2J�������,<��9�鉙~���O�D�O��'r��ǥ�<Nޢp�׌�IZ~1!��'L�O?�$ҙ8̼x��2c|Q��]/#=��hO�W]��A
]�0Esq�X�pQPxk��Y*7��Ċ)�B�o��t�IY�ԀD����'I�"�9z�,Lj��@#q�)*�cǱ ��KΤԠ%��'���M�(�.^�C� �_|��2������CQ�f���A�kh<ѢT-�5/Z"|�1-��aP�
5q�����-���o=b�D(�)��U�@�I�� �8w�5���c	-D�#�)#3���)�a�6l��/*����S�A�D�'�f�
W���t�⑬��?)�^]Ɓ� k��?���?a��u���O�.�� �"A�
>a]6qY6��4�R<��&$�d�W�S��a(���-ExR�ǖNH�M����Q����ԇ>J>�����9��y���Fb�aۯ�(�)���u����(O��3�K�|1�����Y8M�й��]���q��O�m��I.5�`���T8L9�MY��C�ɛ69�E��Z#��s�	5B��d�i>�$��;v�C슽ړ	�H1p!s%��=�`����,�I��p�I
^�����џ�'����������Gu����*M�����H��Ę��Ne�(Aw�͌p�p��!�_�}}>27�W�u���z�jE:�)��a�?K ��Ad�u�'��R�/�0U��O�%zD)��7#=^-R��IC^���d�W��?�EC� �fA���T�݆�22#�t�<����oV:T�f^*}^��C�g?IuY�D�'���k|Ӻ���O��PC$u)q.�+&,fy���(����J �b�'n�*I�f��A �ۣV���%� ����wbD�A�,Ɉ�X ��F7T"=�SD�"1Θ`�F�gO��Jc�̔I� * j�Shz,�1OI8���M#��t:1��OT"}��#�4����σ�G�x��ÅY�<�Z0H�5��^:I�2�@�%�_8�1K�����.MR����OVl��e���ذN[��M����?Q(�Tч�O�dgӬ��o��')| 'S	(��H(pǊ
M��8y��ߺ:�E���0�sӲ����y< ��pz9y��i0 0�5��6D�p�C6'f|����iT|)1ϑ=d��b�
� Җ�2�4,!�)�	��S��M��o��W_.���ª'�t��%Zx�<���M�Vy�ᐣ͆�1M��Ӗk�z��?1B�i>�l�
Y�����E?}�n����k歘��?��N�ҕ���?���?Q��"��w�>�
@9`LIT��<.(��+��ȟ�HR�ʔl�xʁ�'���w�\�b���9+�����LW��q�Y'r�p�3��^��dTx˰~R�e���'�^���-N�X��A���Yl�˪O��j��'�,��D�'X�|�� .&Z��G)O;!��T1�ȉ�)՜C<=�����W�N���4��O����Z���X�X1t6H�1jM� �8�"��O����O������$�Ol�ֈ����%���馪ִ�@��Þo�<�K���]�j��)ن��Ox�j����&�v�+�؜Z�OߟI�@Q����J��I=w�i�4��9q��.�����I�l	�@��k�)���QE-B�z�i�%"O2�����!��YrkH�5v4\���'���<14CU2L��)��!ӕ*ft�J븟���4��I�a��i���'���� <h� F4i��� A�wa�	h`I���?���?�'Bԛ>�R����$6-X5fO&O�����"+A�|�51g�
uᒩ�3}<�Gy�#".�af��P�
�a`�Ί<�B%~��)��-���E$2�� tG?ʓAv�����MC��i�b\?=SLY�k�܉�F!�C���90��3�?я���'�"�HÆX9�=�+��]�	�C��ͤ�Ha���1�ܠ#��d���b���!�?������*N���$�OZ7�>+��P�C�58����+!����/ >�8�����08��m��d!���:�s�� x�������Q��'���Ӥ�i1��8A�JM6-�!{��i#C��1���h˅��s�ҡ!�:+�r�1�ɗ�dgPY[��`�:�['�'o8�O?7��k�iv ��C�XM	�V�]�!�$�9d֜����B�b���I�;qO��dx���$�i�&İ"��'/"�Ѩ��CT:����O��$B P�Pۖ��O2���O��Fĺ������+�?;2�a�H.6�6xXҌFߐ�� !RD:��K�ώ���'>���H��OھE�Ɗ��Q��-��c��4��8��7c߀��׫���N�z�bd� n��˓9��puL�_)<Y+� ˲hv@d�'���j��Y�z�-�+e�����K)g�
<�ɕ�yBi Qp�1��´�b��dC{�(�Gz�O9�'b(8�/�(?��݃�@ۋ�$y��,�'J@��3�'7��'��:?���'��I��p��x򳭑&}��DgM$��YS��$`JH�wNL�X<���TB�'���P6D�t)���"? �����u�� �Z�l���s�(0�S9:�$����\6��i��ˁn�$E�ڼ9gn�87���1J�O�d�<y������Z�jaR'�Q�e9����'B*lO!�ۍf��dN�5%4�<�FC:����ۦ]�	Ry�_0��6��O��D�~2eH�r�Y*5�D3G�b��&C�6S�LH�'	r�'"��R��@�dn�B�&	k}���e ��ܯD! �مi3SE�<������g��w�\���i���0���?�����6��ZǄŷ�J0�&�+ғb[�I�ɍ�(��L�aO�r�ڤ!T���C/���%"Ohh0���yx�d��D�D�'���'��@)'vH����_!ukiP�'2�Щp������O�ʧ}8�q����?�4 ��}�˕VF��`�Ҽ?d`� ���V�\� r�^�3�l��`�H6��(d�r ���\cA!���*���'�!��	ٴG�llz�*�Jx�!�� @Z8j�n�";�!:�($�\cǜ{Tb�A�(!A2��h�4�شa�J��ə��S��M�!i#6Ģ�z4���5�h�2B�v�<� �S<q�� !�U��bPR$�m�'}�#=ͧ�M��G
�8Y�p.�Dnn0��͏ ���'��$d4/��'���'~l�����R�\/ mh�#
=[
=�A�d�l�愝r7z���޻an�h��Y?)����Я���UB�K?�@
C��p����(B<J/H��!� ���dX?�SbMo�D�r/�<��*�>B���J"�tJFuc��	^}rgW�?�&�'���iD@�4v|���ݤh���'��iЗ���AM�l��J$oj�<��By���ԓ|��ÕO�6��j�#�Rʢ�C���DA���'�2�'(n���'��8� 8s�䖂�Z�!�%Q��|�A��=7bX�i2c
�t����+��'�AF~��B�+S\$sv��8����f���m��m�N��H���ź_5zѰQh��<K�/Gh�T����n/�	�t �"X0�("���`P "O�\jT̖�<�����EJ�N��"O>��QI>O�d�E�!G��8��O��>�6oA�`���'�S?i��	�pR���"O_�^UC�6p�&4P��?��ư�"�nFG>f�z��K����j>U�WLZ�:�
�;�PF#Vu0�n/ғUrA*�^�8����+����![�>a�$h,B�LŀJ�hE��V�{�@���O.F�Dl�,ld��sٵED���m	��y�iխ(v�����q�
�&���p>�Ǜ>��#]��T��#�R�iC��0��z?!�oRQ����'��P>9�R�ҟ���֦q��2 ���UO�
M6���In�"��Lo!$��&K��y*�~c>7P�j?|l��[�x�(��95��&	��_5bxb���(%�,������6i�!r�9�HٗO�:�ڂZ��Mn����J>E�ܴ[j���A^�[$^@*�ᆺv�V-�������c
	3��r�D7a�D�Ey"�+�S��*T;W��(�HM�ơ�H�d��O�jsѥB��D�O����OhI���?��'�t��dhǕk���E���608@m�|�f�u�k2�y!3�~
F�	
1�J��ݫQ|\ q����n8P���t��@�}g�좓
�~B6h�1>Bb820�<���4�a�]^r\M ��	S}B��?���'5B�.Fôrp�Y�L0�(��VQ�<��bǠX3�	�lz�1�.Ѽ_�@щ�4��Oz�@���cy��J�CߗN��lQ
vɜ�E��O����O��D^<y����O��ӈA�,��xӶ �FT�|ό���,
(n�B�z��'�r5ۮO�@A�ɗ[�͓���K�f�B��'��͈��#!(<9��ܫN���N��a�8D����6����ʚ�p �}��"0D��JtJޚmDP����G���ꯟ���}�ՙ;4�7M�O.�ĺ~��i��j�uᐃ��;�F����7j�|x�v�'3R�'���5�'1O�S�D�H�"Ɣ ��5Q�6=�#=�c)M{�π ���vb�/G�R h֭�&������fVJ�$c�O�l�JA�D�#ˈm�u���GndAs�'���C���?�ƽHR�,F8A�iO�!��#��M?Jʨ�ؓm ,C��^A�V�i���'�哽Hk�L�IҟpoQl�T��*$��T���ᑵ�F�� LPb䏿p�(K���mx��K��#���&>���[Se΁a���6%��)�A�C���*?c��Q&��w�P�!dc`��5f/�-#P��m��O�B)�u�M��e�[K>E��4�2ѥ�>f���s�'[�S����ȓrJ|2b!�^=��g�J�<~Fy28��|�۴/���Wc�0k�=+T̉k)е���'R�~�H�ц�'�R�'�R*lݍ�i��H��U�G�V��cL�m�$3�U� �wĊsQT�:��5,O��O#m��I�.�0[�h�U�t���@d�T}��(,O��(U��@ �)�%ӁF0�p�]�"!��Or���I�sɬ�H-��#��ەf�,:�C䉁oP0�$�-t*4�U�G�Af,���"|B3DC�nP��e�7Y�>����(�HpK&�3�?����?	��z�d���?i�O���tNR�6<���j�Yͬ��e�S&o���ղiE�}���-n�0�G~�h�h-�e(�H_�.�d��v�˟l�As��^}0��YN�PCC>u�bqCsτ�㞼�g��O� �2�D�K�$�� s�����_��y"�H�~�Y�+_�:����y�T�K������8K�d��𣘾�~bA`��Oz������9�I���O44��l�>&\�U@�6zt @�"� ���O����5h� ��
�'|�S��HԞ3���]�|�yS����HOAgl�N�Ƹ*��H'i�R�y W?�)c���2P��O�6
|�#(=ғB�Ԅ����(��쩥X�v3ڙFJI�����"O�{'Ǒ�t(�k�Ȟ���q�'� �'k�0�f�X7~HdB.�br���'�]�B{Ӕ�$�O��'<�[��?yشV�QA��?2D����a��th��R
JE"�b�Z���*�`h~������5v�}[��ɒ�Y� tٻ���M�"�ҡ#7���У�6LV�ѫ��37�0E��E.
o���5�b��B�4��/L=9�l�P�E��MkC�ٟt�O>E��4T$RIұG�2k�Č+4�T<-�y�����I�bA3#H�" NH�|�0 Gy2�<��|Jݴ�*l+ N϶ry�m��R+F�nXZ��'��$JHa����'�"�'X��r�����qP�!ݺ%F,T�w�_�^a���V�<p4��DO,}���QGoX?]����OF�B�큐�9r6�¬t��=H"�I�}���Ѫ�^| ���k����V��9�3gR/g��I
Mٺ�Ȃdې��	�e�	\��'߆�̓�p=��+,܎i��)ɚ�a���t�<Q�N� ����7��;l��3�J
u�"=ͧ��Ne��ڷȈ�n��<��:`��Y�b��mL�����?����?	�J���?Y�������"�*��mLƸ�3��[�6�¥鈷#�$�GK�$s�|D��#?�BV�^p��e= &ra`��TB<Ƅ���Y^x���z���e�Ԧ	���Ƴ5�"�%���*�O�6�٠~.��@�@�[���5+KN!�$C�n�!-Cı*˗N�b ���HO,�-�c���i�s�>4���Op�o�P�I<i����4�?A���I���HE#Eh�4�8̂�A)z����)���d����#;�4�W�נ{�8Q�gZ%p`�i�O������lئM�D�2m�0��H"jc��I�[�朳��I�� ��	?�,C ��#X���U莇1Y��3����=���N>	��������	��xW��
㎍,�9�$*^�!򄑒]~�h��3�N̙�蘿J��hO�C��)�d�;���C��`��'G�wC��FC�n�����\�$DA�(���'$��f�x~��kD,I��pZT̄!ijVQ�Ǜ`��P�tn��E�܌�e@���$���m�E�7YUPh����r�=���i���e�NqZ0�&[V�qJ�-�
�u���o���eɧ e�pEEԩ.[L�1e$��%��Ox�nڬ�Ms������\=?v���Z G�&��2�U�~�'�a}R�E-v��\�0C���3� N��(O�Ez"�O/���1i�1[T/ο%{�̺��՗Cn�8�����hO�Sj��*��O�o?V�0q%�#�B�	'�� �0��vnAm�v�b�����4��I�Ub&ՒWK"1	Tz��X�/DrB� _�p�q��M���)�#Y��C�I�N�0��`
�t ��+_�I C�(f��k nV2���k�/oC�Ɏ=hRY����-m����*?\B��#	�`8����UIt�� M�g9bB�)� *͘��X�r�S6��@}f�0�"O���#��8��%Td���C"O�u�N?��8!����C2�A	A"Oz��n��~�=@�"�,���"O��p�ζ
7�u�#ϳw��!2"O
`@��X�D�]D� ���"O8�v�99{��2&B?�t�"Orp�M�ZT�1����jiu"O�����C"��Yf��3/����"O> jHϫ9����R��	N=c"O�D���ܥX^J��w����,+"OT��0���,���#X�Mv�1;�"O�C�@�\�Zh #�W�Yh�qyr"OB��@� �.�����*��~�^�B"O<�� �}N�@4H��	��<0'����(��L�
�)�#�$<�Ӏ�$N�=��a�!*�Ɲ�aꙔy�0g�_���x@=�T�!��R1+�R�:���.| �č�_��]�*��D�t���^	@�؜�U��p�FCd�������|�&�!�˙�9CD<ba[{��\��nC'r�Q�Ǭ)�H�S���h
 l�R' �#pܲ,T�6>ؘ�栂�.v�:a���?�C�M)j���p��l����c�6hѴ���6#>�4�/=�܉l؇,��5�@�٧K��͹C'X����+2�#��\�8B�a��EH�}� �ӡ��0��M����C�k��`0�ƕ<��x��_�W�B��iR�qg�4��)ke���i��@ppƔ�y��@�^�S�,D�֩�1�vP�C���	M U�aN�&@�& #�*'��ܘL��I���(J�0(�B�4*��Q�ԀB�R�r���0*�}ۂ����V�B�L�21�7$�E�b���Z)h��U(H�H:�³a8m2u�u/�y���	��S*=ay��^#�@�ɣ�H�oG���P@G�V�J1R�G���B��v�(bT"U�#Tp�y�+��jN���P�ǦV�P"U�������g;�ђ�e����5{1F�~�Q����*U�c2���$�F���!cm>}�L�f�6<$c�OX5^G*@��k����:�#C0c��m��ă6H�� ��n?��[,&�]��� �N�v7M�d(6�1,�S���r�|��e-:�@�LU�����eX�}��y"���Ph5)�+[�m���H�b$�(h��>)���(�N�/iII1dgH6 "�ډ�R�愑G~�PC�R~�'�(�y�P1{TR!�&W�gX��9�,B�V�ۗEգl~	Q&e�b�2�!U��2|YRj!�V`Q��Q�,B�SI�e#1�؉$l���I�gG�]���4j��`��I_�'�(�í&���� �C�?s@����[�1t��b��5�<|��Ջ^0��[��"q�L6� H�gU^7��s��*f�p����f�l*��ǯ5FU"�CC'V� {戀&��'�4Cf�A�df�
�D��p90pr,��c�@ꆆB�$/ة3 ����,Zq	�-hd0� "�]:�Ԩ����#��ܒ&ƃ�&*́{�(̘���	�ka8��先� q����� ��\�\_��x�"��j��xq�`�̵��
( Q�A���xv)�(ZR������Y$X�㒢�
��`O�"xn���b�=*&Z�8��
�~�G�X\#RݳR"�	������<��	ԩ^�Lu
��K���Hè� j�B���t�H�#o:dAcĭ�+T�,���`��?������5E�*�je�]�$����2�65�q�t�?�ȝ1")K�)VzIpc�[�LЎ���
"��I7-��=K#��7N������z+�U�E+�"kr��G��8u���W��X�4xRRf��_z3Gظ"�}���'$hr���'�?w�Ы�P�x��p��^�.Q��Jե
�~!��7a9?��
�z�T(2�C0�:���O��\��O�����P�
4�@dauEȾ;�8�ٰ*�6��H#��VW����I�	�K�?�W�(,M���t�Vo���9���[�a�� ((x0M�8�����:b�2����)�9�!�%!:PZ�oL�=�D�r6�B�.*\$KPF�{v=p�#�gm:t��4cиإ@h�r�,��Z^�p�@L�[�:�:`$F��M3a�
�~��8S�h�	6��K% ��rȲf�TU�0C�<T�%{����{��0S�`����?S�1 J,]�U1q 6|��0�
�C^X�!ە �m�� H�K�|S4%�,^�I!P�$᢭іU�bY��T�3.���S��.s̎�[ck� a�Dah�=?��
�LX�7��	 f
�2(�� ίqɄ�[�^f�PuPsy��) �Z8�6+Ҵ�Z��� ����'�D`R��(}��G�,L�S~��Q5�B	
�й�㭓�0��egh�U�&��P��<CJt��5)�l	�ޭ�#'0����Q�$���)����}��Mx�薧| 0a(C�2Kb�w(�A�z]�g���?ͧ|��Q8$��$z&Ih3��0Md�Vg/����@�G��@��F� j~���!�Y.>��X�O$\o���'�$������C��`���΁�M��kr�4(q���z�rD����1����5����J�${�6$� �Gp�:$c�^�y�|L��1�b�yu���^Й C��
M%���̰V	 4ѵ@�S4�`D�Y��(+�@\
�	�C�$���@� b�yeǕ�i4����k�`�B��T|Rݳ6ᓊe����vǮVo�uHՇT�o �Xf/ȸh�d�J�F�W%��!T�H_T����@  Xp�b\F�T�e�>�h�9:����k�3VV�A*��y4�0
��! �J�&ިe��Aݻ*�8(��l���D1B%mȅ�B�b�)CP' >,V�x��	Z�pⰜ�p����!@+i�fuk��ǔ!M��B#d�O ����6�r\�$�>90����y��
%�v�)2�D)	bMX���UJ���B]R�|[c�����u1u�T�(�Mu,�51ov}0qIPX��@\�T�L�6O��x�T�uY�Y���/T�Е�O���R�ȣB0i�B$�/&�R�
��^8(˔����/I�
򬄨2��5A�đc4���
Ev�2�ɑLX� IJ)fÉ�|�B\17�̌H>9m��Ɇ	)��X�Tb~��åV Y��A�GA�y?�kE��=8Wv%��${p��cX1PkjԳs��"_��mJ0��4~0�!#��هDJ�{�J��V7h�.tƕr���@L�sO<!�@H�	���.��:�l��D�P�4���^�t��2�z�����ϝ� ��9@w�ʁ)&��'h�*��=H2���s� ز��z���a�܂%�� ��6�p8aE�Qw΄�� �ӛ��$��� ���Sنp�@�$i��8b�ߊ!���9�� "�	!&:� ��{qē-h+N-�S#8BGh,a�I�M*�V"�;<֐3td�T���;�Ē�k-F!�3�:FOxYe:OF\��M�=$�kWB�Z�kEÄ�{ݐV[��܅(B��ğ� �%�#�Z$�N܊'p01nUQ�a�v�� e�`�6#@�W˲�;�%C6i��Jf��6o6�*��85S&D�n�a�$�sl�h���Fy�]�T�˗d��5���Ec�Qʆ��Lʢ@1��� {?��xDfۧjt�I�d��d��1�Gc�Co�yږ�N�1 �AH :��r��4C\h�u�Y6��K��Ȱ�g$(y�[ T�Q�戊��s�+v�1��(f��}�s�X0N21��G�j��*�M��9|�Qc-t�-A&�(f��A���yӈL*҅�}�$4���^oB�Y��i7W� ˧�2T�Q��$'+��@u`K�~�4�A�_�jH�y�b)�5Q�$�Oäa�$8ӋD�aRM�fd�����d�@3�D$eFmÖ�~����6�Xl2���5jC|��l����οG~�	0�őDB8Q.�k���ST��!�q�&�0���WHO��6͑Z�����";sz��%Z C7>٢������k�gӸ6�M���suNC�4�J��Q�?}�}a��c��[i�$���*6��٣ 	���
���fH�M�6���
�Ұan (]m�4���6��������������D��D�	#�(�B����a(EJ��T)��>Ic��>����$��Q"�ԠA���19���)�SVeR�M�~�&��$
2ذ 'g߆|�W-R�M�X�p� �8]N�I�k��a:��ƛa�)�JHi>N��d#�q��#�d2X� ��#�I<t-H� �AMH]ӥH l2T����t� �Kd�7R��f��/&�*�4�Й_�Zh�wD�=R���:����N���ȅxK��%�Y�yH�i٣6���p�ɖ��$J"<�L���LL�ps�
��<��,T*$����'5��� h� 9�\�:�a�ML�`c�����LC	?E�Qb2��>Z�4h���aW&��$�妱�w���*<��ql
�y�'(:��l�q�`j�$��0~j@��ߧjVB��f$�H��
gG$g��M�Ve��lHvTJ���-3t~p&*ޥm_T݀��&F�IVn��-3����ߦ_,l� Teťc����"�8�J
J��ٹ奆0;�jыd�D�����l]�4�c��X�Q�;'Θ7PXؙ'O�e3u�:t�}@���&�#v��5T頁W�� ^D�1N¿s�8�E�����h@�[F8��X��i�)���l9E��p���Ŏߕ���(�ȗ]L,/Ia���"&�@	 �eT�
F���-i��zЄRZ�ɰč�b	����(L9xa�N��3���<4��ɀ��)���E��FՌ	)ɟ�kʄB��?_y��Y�6��Ő�!L����a�Eӌ�ߎå�ޞ>&3�B\�L��a��!�$���#���1/­��7Y\<r� = *�n�0�P��A�_���:�)\]��-����%6�L�u�	,7�ҡ�e읃K�`AC�#�\����i|�Cg�ӹ]ݐ��#��%�.���}�y ޼CZ���H�H��\��aZ�����'�έ�D��=�揟�(��hjGD��sl(���E^�pd��f-�VϺ��$U�V��xG�.h��5Su�ʓDJ騱垌pxho넝2VE%�f��OM�Zr>aq!��`Ԃ!��3W�2����� �Mǯ�,;�,�M��b�+�ɸ%cG�$'I|��D%�M�\1�4K�Hһn�� �7+	4P����Ճ�B�0���/���dC��LY;�{��9j��0ؗ�Wx��b��;&XR����M�4D;% G�*flY��T�`�N���]>��uA�
P��}kYw�0|S�²	≂�"�)��lH�'>8���*&`x� �8ʖ,�B°���QB�>A����Qp@�Ҿ:��aq��������%��qI<�룬�4�4�I/^f@PQ�R�
0oK�t�@dL��7-��s����z�����R@^e�2˗E�i�g*�	�f�juD����[�Q6`dh��%�$I��e"
��i\�f���w��tZ����C�^��C �-~q∙G�,4$��E�]�n�����y@��Rカ\������)Z�u��.T�cX�!����8|I�e&=�V�QV%� Ld�㧄�n�OZ�2A��l$�ХJl��3��/���VrӼdy�z�8�s%B�z�:\
�K#��]��`��$d�G냠>;vH��t��tN�**�ܻ�ap�t`���2I�֥)�E�|��e�.�Sc�K�-�lm��E�z*
��$�T��ɤ���oaR�WB��:J���O*���� �O�p� �E71*�ʒ�$;�`a��5�f��P�((!��a��*�X�PRFd��d.�>���Y.<�=0EE�Jt�]谊�m"1�`�A�Q�Md�Y%˪[�0)�'-��pú�F������u2�'D.�r�k͡`@�����W�.$���J�U��}X ��;@~�!T�H=�2�H��_��ԭ�#��jv�	,d6����և�y"��d2ԍ�2�S�NMjy�
çw��db���}0�[�ʧE�ƄAw�M$����g��:t�lbN�v��b>yJD��ټ�̉%h�-�Т��q�p�-�p��	�;��Q�A�ԶRs�iI{I6��K>yr��s=�\�S���:�%�P�D?.x��c�7:_� ��.��H����	q:�x�<��q��H J�<���R�f�Ys����Y5�%��4S�b�Q+Odt��d5h�X���̾H�r4��L���4G\;�� !�	��]!���䡟9Jr��;g	8vqO�bt�
+Iyx���)2c����a?��C<S�L�q�h�
�bЅT%>:�iT3��\ɘw�  2��Zk���W$�78źt�b_<��g�P &����W�]'V�(�A�	�#8��
�x��E25L¾r����%����w���*���x�J�=��P�3 �@P�fP8��OPe��� 6��Y怄�?��r*8�T��'ZnX�P �&zi�S孃�L�,�rE��H��F�zX���d	Ws0`�:C
��8��|r�i�OrMW�V/7��AÃ��&E�4��D��p8r�j�*޴=ˮPD)�K�zѹ��;5�x#g �9t�� ��ːx�CH��� ��-Q�q*����L��C<���q�̐_��	�b��e(�*�����џu#���ф�y7G �v3�!ѕ`K	h�X�Y� ���>I�ڞ4y gJP����J�htv$㦦3^�� ���=��)�gưkg���*�����ꝃjs�'�Bar�F�;�\l�a��c��L<Ѱ�� �"7��'R��4��)dĚf�%s$ iJ%�I�y�@)��3|��V
�	M��7���&.�An�d��˓D\��#�V+��cOѩՐ8Z`��<5�:B�>0����I� LL��c�!P&��;��Q�Ӝ bd�M&����	�]�^��m��FqY�D"�O�$`b�]�r�h(
�i� .t��r!L 1^�9G!T��$����-� �C�r�l$*��N!-p�=�¡�8N��-F�:�Z�Gi�QT�U"GE�+�J#?��"��H="��B�8(M�&*^'���ݙ��,�Ʀں k��c�C�=�ءAȃma��KR�9#1���M����f�[8%g�)� �Qp�/�4Ǡvf�����:�Q��!F�ر7>=(t���.(�gL�gؒ�IC�N��0��0{��H�gE!Cj�$���+8n)��imEshP�8@|�1S
Y�|mFRB�du��c�L�94�qzff��y-��hv'�!:c���cS��C�/F�?g�Y����"#�JH��l +/Ӡ)����P8��ʑ����8�
�-�WI1�p1�7�9�f�i�(#L�$�(&d�c�ǘQ�xY��2�~7ͅ�t<�`�
-!N�Z↓�q�dYa��Z��Ah���09����<aЄQ08��7Mt�b��O�\��m8@$��8���	7�i]����?�F(�ץ�e=�����7���sJD|\p(F�\�(Z��H#���A�"�<*?�)Of��5Ë�6$К�NX&C��\�SV�^1�`01���YR�*8�`Ѯ���'^�����V
�za�e�1���C��˧Y(x㐪�Y�8���2��T��!B7��OP��p�<�4��2��m�aNM�a�6�c!�C�,@�c��a�B�(H��!����� (��S�<.Y���_�f�4%�#����\D�D�48
ў,�g,�*N��T� ��&���M0aZ�ό?��,Z��H�*� �~e��Յ+UJ<]	d���?�8����PY�b%�RE��#� 1c6� ��BJ�wb\`��U�~��	3�Ȥ�f��
��,Ɩ#z@`ySn��o�X����b�d��Aʛ�r��ȿ)��%he���Qqo�1/И̃�i\T��9aK��`-����>+��1�'�� ��I�>PgJ\!�R�op$�h��	2l���C���&f8����	R��)ߨ1#�'F�M��R�q
t+8�V�k���@?&�{��2F��)��OD>j֙���|�U�7H��{�%h��,ﰽ�W)�/�|�W!܀3�<��a����	� e�ml�6�>U��C J�(P�Fb3��e0�B_�_D��`B4l&ў���,+e��'�x��Ƞ-�a�1���(S��E�F�
2G"pN<��-̔"o�x��L\� ���#%�P2�jb�H���K`����]���èq��sWH����dJ��v왧/"?{�1����iݲ4� 
Ɯ~��s�>� c&F%f��͠�f��`h�s'�R�4ltDZ�ݍkj�L�A&�=s�:�SF�%g���3}c�c_\�"����Y��|u�xb&�Q���۠�Er�Y�o<�)	�&��'x
xp(6:���5�H�,`�%���@��BA�s�>[����"F?�y �(f�UyU� ZD=iEa�+����ѦQx�ȵ!U�R,�R�O�8����+!�(@H�B�1U;R����M(G�F�`!o�2q��Yt���7�QZe��(��y���.�&���,��2�O���̰e��l5nĦO�E�!k��N�`̐�#�'w>���F���Wf[�'0r!�'�� �ʹGr�D�G:�@Z����O�~�b���Rm����ߩ��#�W�w��:Ŗ>Q�>9���H�bMY�s���8wF`�,���U�.ޚMoXqa*��|2'/8}��A�)
v�S(٥E���QJ�y�@�<��Y��ɃyP���,Գ.PV��0���j9��f��]�H%�r��T`SP���p<�qȚ�ZФ��SG��x���ҡJTX�L���nc�Mb0�
(Tx�����H	�u
N�es���z�E�ēS�� ��=p�.�h��y�8�<a��x�>#u	��:�����b��o�8���ڱz���C®�y��ݓc��<�S�UY�S3m����5)��J3[:��O?�?ҸdФ˖>1Yc��6��C䉨:T���iÙ'�>�zP�N�|�C��?4�T}q��N�<�,5�r�Y, vC�

���]$�����Q�B�I�-� �qHΛ4��(�0�U	t�C�I�s��e�G)�~��8F"� �C䉒.(��f�+�zX{6M�0 G,C䉓<H|� ��C ��X�iÝ46�C䉄UZ�i�"C2^v��� کwB�C�	?`�A3�
�l��y���ZhC�ɟ5�꘩b雖c�ܡ@T�ٲEfC�	�9�(��*1�؉� �U�YVC�:�i��F\uL@d-!|(���"O�qr-ѧ!�
0c�D��Cv���"O����V�U����	�W3�Ay�"O�̀�����m��&�P8=��"ONC�@Z-V�ŲFD� j�(�"O�����I'oJ�`h�a��a��<�D"O�XÂ),r`�e���Ap"O )�+��HX�c3�j�T�9t"OB]zG�L�B:�y稗=]�Ը��"OP��J$M-)��"J����"O�Y�`ߢ^�Π��g�,-m����"OJ7F^�a�y��H@�;o�E��"Oh���ODP1�A��"KL�0�"O�xc�"F�P�T�2'��v�����K�!'|rE�$�O.8K1��gԨ1	1ɗ�>	�!9�"O~�V��G�n8�!AќEx�"O� �B��T �E�W�["�0|�W"Ot%	CnR1RN14

��|�5"Ol��'M�7��H��)ɭ6�����"O�ъ"52ʂ<C�H��s�=��"O^�m�"U���PT�	 b+~@��"O�%��K�nFn�����vfA�b"Opq��Z�*�+%�0x��� �"O���'ҾKW�p����+�Lu�q"O��Wꊅ9��᦯<�*DR3"O���a�F�MN����ׁ&�r��"O�u��E��ԁ�M�{�8���"O��ǍN3��SUj�V�<}9"O ��QA���x�Y��	-���@"O>г���+2�Y�������YR"O�UA!�S&��ӕ�՛`B�"O���e�/	��m����g�He��"O,�ȗ/Y:Oڔ�����8�I��"O�(��P�,��m �
ȷ5~Jh��"O��j�F#�"3i�nr�Ѳ�"O�TR� jH ����ƾ_[�9X�"O��)F"Ͳ���R"I����"O�� 1BT;���D�}4� �""O����U�1 !�G�8�l!"O���#H���Z���#b2R���"O Lp#��{PI:.�+����"O8��E� u`�����F�*�,��"O�$���M��A�R��=��[�"O�-P0�ֹ9�t2b(D�!��]��"O�YI���ՈY�GҀS:��v"O*U+�[F�J��q%ޡDRe�w"OrP"g+S�A4�0vcLR��"O&h�#JߞY�12��X�`�#"Oj�i��W����#���!�x2�\��4��K^u����<C�|�w�E#���Q�I�9�pY�@̾s0l���?Kи�ؗK�E����3Ӧ?���� �',�q����E�v-[��#G�
�Ja	X�gǒ�H1p`��@�dp����%8�,X���n�J�P`�E㐴gab����ʍ,n����ߕ�퍟^y� I�+ȉ	Q8�iF�E�1�^��c�D����K�f��b>���S�&dڕ��ݾ) �q3E��Bt�@$��B�����6�
<�1$�XB
X�g(1:��H�a��0jp�jBDרk�N��^�T\V�ߺ��̪�`�K�m��P��iDHϘ�����e0�� �@G�R^���`�����H���X�FP��U��
�Lқ4^�́n�����R+ ���) ���&V���%È>^����FH�8(���+�2��䘒l��A ��MF!��gƣt��"dѡY�(�`L H?��倢��G��-�� �OQ���S��ko�H�w/��W��p�ID�x����w��TX5�?1�,u��Α p�H��FOC�q�����Z���	�9���?�q  rd0���iD6rZ�C�>�́����>����~x|�q�"�n{DM@����9 Ec"�	mJiC�C2��R$�P���H�tѶ8&,��{��D`$�7ОIe[����B�����Δo^, �.z��[^�Y /�t�T��h���ژ����5$����C�D�Hϖy��L��Xi���ܰ\�6Q�w��;d���.��z�,��a8� ��D�;`#Rm���v�ڽ��E]:�4�2*Ŧ1i`)k��͛IT��J� ��l���)Z�OHF���)5,9��]'	p���C�9�����weL���)�T�ڠ��K�\��V�\(�bAH��:��A��Je\��b)V�! �'2��P(g"�#�\�Mȍi<��
F"G`�tz4�8�(�nM�E/H�8 w����QuY�]R�(T�b�P���6�?A�h��pa����|޸l �O�)�HK��X9!<Q��O�@���K3e��PZa	 �C�z����>��� ��PS	:vvyk�d��<As�A��bc_	28!����vZ�I2/K�N�p�'�
/�##M��$����P7�D��d{���W;�q�����>}R�M�"�W({��p��#>��"g!�'j�I��$ԟ,"���蘾qQ�LB�S,����&*(��C8l8ڣ>�]6c��uy�C�<���f���d12�M�GO0%�'i���B�(��e�8��]� &� E�L�Q�+R���	dj0� ����:"$yTn��k��&TY��QS��h�hQ��@)�큇T�2�b���*pAH?���s
�0����69sd	��G��*x�'���&G� ��a�u��E[� �2 ��}�@�Q�ή(d����0h�b�#�:qv�̊B�����z�7#:?���l}��Y�	��!��'�JO8��"o�$b��RĎ�o�|Cd+M�/а�E��8e����5�E��|� �u�ax
� �`���x�l8te�"�`�;��>�t��{�4��sf�"Z�`0L����x��_(
r8Y�N�#d�Z��E.�'Y��B�I��U�}���X�Q2MR2����l9E���T���iHė�~�A��D�r�> ��$�DQ� 1�� e��'	�mCf &J��cQf�' ИE�|��:Q�Q�*M�;ㄹA4�[�B�¬�	?+�Ż7�O��|"��A_�I�l�|�c��4�N�@
�"����B�P��XJ7�1	$`�(� �?ӧ�@� Yy3-�7t�,l@�cC,N�T p �dS	T�>�2jI��G��5��� �2!��̑9a�D`r�Obd�|jP�A���A��<�����c[�0#F�I*^�V����#�I�L!9��"����aau���e˲X`�	34��Qs�\��MtӰm[!��s%b^�k��� ߟ�ԟ�I��@���$s*��Z�'?�'fTuK1�3�n��k�S��}�`��W�KU��9�	~Ֆq��ˁ�B'�v��?~G8�!��O�(p�|Re	<�I-^��;C��}��y�sAU4y�4� dM\�w<���A�8�TD��@2�'}�$�`�M��,>蹫��g����#H <Fİy��.�DD��>�]7gH+�J�m�i�����2�ƀ�F�4X��J�T?���Y�D�4z��p2\�y���$��ч	u���SrG�Ȁpk��W��q`%�==����E����2�����[Ц@K��� �i�U��	��<���eC�� ��a����>IІ�o��(c��_��yPo���I!>�w��0�QawE�[��S�z���A��r_��Y�M��@⊆�U`]�a�_�u��5+�d.h�Z��e�d���O���`� �X-	���5��f�*H��CV�ŲɰHX"N�d����d�3`��OqR%ͻ!��Ia�M���J�^���>��A���M~&�`�3�	GJ�q�Rd���գ-LJ�h��ʐz�4�橍4���%���~r���,!($���r��2�Ƈ?7@�k��D�e�v�I�і��t���!m�������C�}��5�Il�ɞ)�l�3lM,)N�����~�h�j�(" yJ��	Ԏ�.�4Bv�X�>k�������AL�#`Ϝū3f;x����c���XW�
*��Il�	5#��I0�H�]��:#ϊ��X�`������:f5��ǡ��Zd��CR��z�ʌ!R�Q<�y�f�9 M�������'	\x��^(�Ҵ��Au�<]`�4o2t���N�v�z9j�憇KL�F{�;�����i윴e��HHц��C?�Eˇ�eh�ᑃ0S���c��44|I�T�IZ�x�"��"/����35����Vg�ڂ�j�F�2�[��DPf?�J>a $ӝ%\���R�K�Y8� +��H�1+x#��VY�f�V� BX�u,�}0�4$v�?q�}LԹ��,[1A6���5�عGyZ���{cI35��1�RD��~>tL�'�@pP�N�T��c���h\��d'U���[E�Vh.���)�	�{Ҩ�E.X�{�(��,��1�fGX0�i�h_<e����2���hOkL�;W;:qX'�ԍ0��x��I�B9
�ExR WA�S9��+�|s������S҅i4�|ȴ��GKў,��'!t��pi
m}�~ƀD3h��>�^�qE�z�� �cX �g�U8W��Ѻs�h���u�]���]SzL�r0�N�!�@5��VO� �b��w,!H���OL�3%��)z9�h"kȍ(w��#�(@"��I3�ne�ׯ��\����\�D�?7-I�bR!!�]A�y8G��	zQ�쒤/Y�"�R #���10�!򡒇�f=P�ŀ��=�M��x�ě#w�¼%?�LA�,F.%�}�E%�@[�]�e�jӜ�ʡlR�o9��OQ>Y���I�;�H�!�`Ȩ'|������iu�W��92�a�$/�ȑi��_�b��9���Έ��OT� C���:i�\�J|Z��L�8�&��$/T�;�i�<�#�a\|܀q߬I�P�bêW]yr�%<3&@��K���TY���&J� �@����'B�C�I`��T0���z
8��
*T��uJ�:t��5(hx%?�LYVd(X����������<�L[Rl`���Rj:�I�թ��A\M#0�| ����/pbI9&ᅵj�8�@d��G�џ��!툤WV���|��
Dr�B�H��ٹ?�^51a�C�'p\�
E�I[)019�OËf�l�p�'�LAs���y�*�S���6q��A
��d����F2s�T*�
�-b�I�|A�H�B�ޝx>6qCw�K�~�����k��܋�k4W���gO�<�Q�,���ʹj�(Y��A�P�9���x�M�҃��*��a���.l����͕/�*8��Ղ%�4�h`�ڤs��]��Oڭ:6E2vt�`����-�d�ѣ͊�0=y���61�2����i��)PU͞�op<𡣪�1a�1��~�T49"�2r4Q���$t��4`��&���� л�Ox��	h��k�$R+vʹ�3��>Q��T��p���A�p��QDi��tUUB�b)�n'�L&�d��e�
�z�3k�0`er���]K�vѨ��Wx3�R.�1,i�x2���H�b�B��9`fܹ���23��)�p$Fd�:0�nֽ[�j��D	�?��Л���X9N����86Ԕ���O� pt�ɕ>U ,�9����R�>�1�7lOT�RbͧwF���4 C��T��� ���q/�"4�B�	=G8��A��A�И�4LY�>z��(i�O_:6q�7
�&s��>5�#� A���2#��1�~ł�+%D�8f�Ўi�l�a��9ȲA�篍�#V욲�F<�`���$�Oڣ}��z�"�Y�$к
/� a�^y�$��� ׈���%\�O�Q�U�2�� t�8��(Ok��,r��kԉ&��8s�N��R�����i�y*��V�M�U�ؙTFȭ��/\�W`�X��d=,O��YCIO�b/���ٚI0JI��2oNfY�!JNq�4��7H�T��4}����%^�ͰK��fb�h�O�Z��ܴ,|H�nO5.H8I�$�x�̾*ܐq��A�+����-�/��'�f���1Or8B�ܒ&?���f+ �Q�,�d��,k��@K8�`�tCsS���������6�� 33mQ�p���s+\���nӁVK��z��R$�| 2��5�O\Щ,�V�\B�O[GupTzv��DrPW�'7�$�0"*�B�*E�Tj��[�蒤t��'ER�{fg͂
�3�'��J3еD����r)rE3��V�"���s����'�NtaӅ1eR�b�S�J�|�sP��s.rY�9p�4�0�GG�>!:�"��aа��9��d�oX����k�\K4��9f��m�:�� �Y����8>�Ԑ:��Ɉ�:���ڿu�H��7F�˘�*������=�C!X<UH`��%�#�$ȝ��Q�F��8��iX~��@��r�Y�?�U�B�W�jZ:u�g����=���Cm��	�p�I�\��Ѻ�Q�;�0�beR%�j�'y�$��n��u�c�:G<�I��WI"&2��Yw]>A`f�աD���э�<����3D��H�g�*5êp[�%�+O�uc�'ƭ4���P7����˓�h��D6zJa  �&
��֋F�:�!�W�J��9�Ȫ
3��mޒ
�D[�cO���4���p=�'��',A���,�D��G�<c�4�*�
g�۠.?��� �Z~�<�!.~J��ȳ��M�aQ#��r�<��A��!J�X�k�y�����NS�<�B�S�?NHu�� ?�Dh��R�<�Ӂ߳gEL�Ą�v;�%����P�<s���0��Bb�W3"�lD`���L�<q 5H-�s,��f���L�<��BЧY��J���f0dyc��I�<9�A�1���R��H�\�;���H�<YfC�"&�\�����>V#Xi���y�<ق�C$
>`�"�D�&[7��s�<9������x���A&	KV�Lh�<��@�5��h�E�.�jeR�o�<��.M�NwP\x��V . ����_�<)R4^�Cj��2#�hGF�e�<13"T/|(�q�������N^�<	�)�,�֔��AU���@c#�Q�<a��M# ��Q��_�|w�8���h�<��aQ�@����t�R=}Vغ�N]�<f�U�
b����d����hj�]V�<I!Ɵ:o�a���5'ĸ|�fWT�<q�@ѓۂ�'�, l.��`�e�<��HC'9���7*��H��<���}�<q�֪Le���Q�^3$���b�]y�<1'뜛w!���%A2.���օ�P�<�ʞ �t4J0IC3֬�04��L�<��`��^cT�QF���1�u0TǔG�<��O�a��*����QD�_�<�G��M�������W�(����R�<I7$75�V )���L@��	�CCL�<��O�;F�b�"	O���]�<q�)�@܊�(��E&����RIR~�<ǮC=�p!�"	;�l#�mRr�<���o�yhwcպ?��aP��k�<�6��W��0���Q�t��%HR�<� R�wg�(�✙�a@"O8�"�'��X.h��9B"OR�G
x.pa�� A�&Y5"O:�z���70X�"R� �ġ�"O���Rb��a��J2��F8�""Ov�5�T�[�<�e�	�U,f�	!"O�ZD�߁/����E�@0!\�q"O��W�W0Z��v��9$��
�"O�b���)Q��Z7&׎	�yxf"O�MQ����l��bF4uM�0$"O*-�#��$r� lz�/c��X "O���!Tn�K�aމV:@X`�"O��0�n
�#W ��á�6�Y	�"OV(���ޒ@�z��E����ZI��"OHْ�kF��3c��d�@yC�"O��(�#L�ya5��� 9���2"O ���Es���:���[8�9H�"O�d���J+�nص	�}xd�O�<Ѧ�~�x�GL��Bvf-P�DI�<PC��T[�L�&�/5�^��.F�<�u�Ǉ|d�,
6"M+���k�<q���
��(��G�Z���'��e�<���%= B�k�H��"K)�"�AK�<��:f�a��4��؛��J�<�S �)pB��uXx��I�<aE� ��`c&)I�H,� ���D�<I�� OQ��.ۊz��[��}�<�N�EqZ����uh�Ȳvh�a�<YP�X3t�8�w��;$2l�����I�<Y2m��f�tX�6@��S@>M2 o�`�<a��؋�x�w��i��L*�JXt�<i%�A�)�\�dB~a*�F�<Av�	4a�*��<]���N�E�<Qw ҙeըX��L44:����v�<y�U��ĊWT&~| iQpF�o�<����5�6o��xQ4��j�<1��ڕ]���Cv}����C�P�<)WeЬ5��q`��ϔ@F"��Ug\u�<��)5�^���-ֵ�a(�'N{�<�f)�ek~C��ׯ6����Bc�<I����+�v`��ȗ*g�L��B#�a�<�O��s*R#i��^��QdWa�<q�j\2q ���W�S�!Y�Q���F�<��e�"W�H�AZ>]�xaY� D[�<�PB�*e����ц<�F��U�<�硒.:��ݹ7" 5mo���G�'jv#~�0b��;�l<�æB�hD5�a�k�<A�$Q;}�ܳ�G�7K ��
�Kg�<9-ˊyo!i� 4F������~�<�M_4ܰ�e�Xn����a�<!c��%V�Vy@QmA*m:�t��^�<i�d��u�BUb�';,��1L�W�<����v���yӀ$!A'TN�<i�I^Z�v��a��#g�� �M�<��ǽ5Nh<2$���L'��(W�M�<a0�L�%,^�+ ����pX��b�<��������"ˊA��hS\�<�E/"4�LC��q�nmu�QZ�<d��EbN-��\	a�Z �@EU�<Aom�$Q@҄�mAM�2B�I�<�c�*}PH6�Ԙr�l!�'��]�<��5y�P���Ү�J`���<�A�?N�誰`I�&�4٢4�f�<���W���0�1jA�Fx�bPe�<� ���)KX8�؅	�6E��C�"O���PBK���Y�G\�X0�D[�"O8�	6C]Wb�ѳ�S0"�4�e"OV�SKֶҸiR��J�I���"O윙aΘ**M+� Y�w��d`"O*��� ����Â�ǻc�Yp4"OH�c��.�x`.%I�Q��"Oa��*U���J��Z���
"O�d����Vbx��j-z�i�"O�\�`a�8FO�A���H2�B`T"O�!���D�N&��jńR�L&"OD[�$Yk���PV�L�w�|�2"O���򥓛m�n���蘸e���)"O�tȃ��W	��6HU�u��Dx2"O
��/�K�����E#��\s0"O�|Hv��	����բ�?�R-p�"O �� �P���˶�Aۊ,�c"O�eqr�_f � j��k�ʁ��"Ov��AJ�.w�F{�"����j�"OȨsq�Y4<_.Ԣb`���ʆ"O܉*��HI&v�y��րb�T�"O@dɁ�B
μEa�]�4���x2"Ovd��CW<frl��2T��b8��"O2���+��1X~�ye@�8K�X s�"O���(U����F���OA��"O�-h�o�/8XdK��{Pr0�b"O�-���M��@���H�0�"O�-�d���fz��ʄS���pU"O0����Bb^@��g�
@���f"OP��g"�<��%z�F�� �"O��(4�����M��D��U�pa�!"Ox�b��L�?�YS��#(�)"r"O*AI`ۭ;��(0�A(7�EZ"Oa��,*���Bde�z�����"O�³�/lz���#ӉRxD��W"O��n��8=���]�4��l؁"O:���e���:����ݱ\��#D�(�b�tX� i�V)�a�S� D�8� �!~�RЧُ5��2�!D���N�*a/傀nY�.��lHp�>D�Tceȱ/`2u���x���#*?D�@{�f��?TmX�
�)\��Ăc>D�TG
ߺEdp0��mh,��0D�H5%JB�L�S�6<�*� d*/D���4x�"Į�Kt�#f2D�L�7C���)�'��LF ��/D�0!D�·r70D�N���¹ʷ�/D�L��ńjWf�ҦjG%M���M/D�T�d$U�D�:fą�YT���u�,D����-D�!���PJBL����*D�T�C�05�p�� /G��9$3D�X�$��t��s�N�S�РYg)3D���G�#QL�㭞5�̳B�0D�L���~���ģ�uW@꤉.D���6�y�hP�'�� �@cR�(D�l�f/Y��{�$�/}t�A)(:D����bZ��S������ щ+D��jF�ߏiC����R�d��-5D�xQeB�r6�����'PL�c�2D�$X�%]`�=�R$�6�"�I��0D��x��?9U���P���8�j�9D�l��fX�d���CĎ 2�K	�!�_5ͨM��B�.vN%�N�0)�!�DG�a�ܐu��8Lb��;0g!�� "daV-N�#�.�cBL�K���â"Oz����B/�:�A�
:��p�"O&������@���e��|�B"O�a�ܥG?e�n�8����"O:��dOoJ�M���0r~�5�a"O6tCgj���6� &ɈfRLH�W"O�P��Ar;��C3V	x?�K2"O޸P`���K�!8��p{�"O\�sG�D�@�UJ[�m)D�X�"O>9���+���ɑ隟u!NY�"O�#�$L=/Z��#)� �&�"OZ9�!&�8#d:8a�HE���%�S"O��CU�
37��c�&#�6U""O����e�8�����Z�~�
�"O�)�� �>�hЂ�P�a�*$yq"O M�C��$E&��s�E�
Ҥ���"Oz<��	S���F%ˣ%)B���"O�$��&*ƀ��r��B@z�QS"O���v�16�(Ɋ��H����&"O� ,�%[���1�����"O�i �B�]M�����3&���"O���=~�(�d�X�^�8��`*Oz ��"I�0NhH�vm��L��'�^Z6d�0x�4�w�QR����'����,�0fб���Q�58�P	�'�z0rfL�=[��#V 1xlM	�'�A��'X�:��*F�&RѨ��	�'��T
wI^'*,�` ݋4Ү��'�d���	���
�Р�=+�'7(�iG�ؒN�eP�-Ī	����'���vʗ�nH� _H��'�J囐,��$�% �zP�<�
�'4����m���ēm�0P�
�'��9�a���AR�$�?Te��'a�u�N��W�q��<w��D�'AF��ddM�n��3a��p"����'-�i��#5p!������<I\pB�'p��+��K�?i������#n����'��!{�����ܑ����.I����'�08�� 0a��2΢�J�'t���gD�Z�N���4o��k�'7�8 �M�M��j�,(Xv4�'�����0��Hѻ"��x��'�T�J<2$�=��a���2�'`�a`�M�Ud����D&T:u��'�4� D�*xԫ8qp���'���1&	�F�	��؇g��"
�'���g	�fC����CgHA�	�'(b(�G����"Uj�[��A��'G��@#n�w˦9;��~�8��'J�P��η5hZ�2#g�6y�D-a�'d2���A��OtV��,Q. �
]��'����cؐc���:`KC|��'�Р�0Bxm���w�A3v�(x�'9ԑE�H#}nȰ��D�@�'��:�� :>Y&�*�īmY~�y�")���vAG A�\�_�V��ȓ\��&IA�Eh�gC�2bu�ȓ8�=��)a�yDOؚ9�\фȓ:��� ծ�q2���ʁ0oV�ȓa>�z��Rr��7 Rq�P��T��u��r%`TQt�
.=��	�ȓr?|u�!J��j&��x�`�&ELش�ȓ.��Ms���B��CG]"+gLl��S�? �]H�+�?\�m"�n��]��""O�P���ŵU+��fnY���"OV`�OV�c(�@D��RA�"OLL:/`�H���M.^��I�"Oj��&n�}�&��$�V O�|p�f"O4A��6�T��l
Ve��pv"OZ C�K@�3�"A�ԏTZ�M��"O ��P�װ�.�[FD�	�4ٰB"O�)0�k�B�V����_v� �"O|���1U�sGC �^r��"O �{bmU�1�fd��+�tL�('"O:Y�E�O")�v�q�hY ����g"O^̨b�:
�4M�e�<W�6�Ju"Ov0U7b*�k֖�,��"O&�9�/,"��U�c���~sx�8"O P��$;�H)�iB�]���"O��V%ɨ:ǘ�Zv�'e�x��Q"OB��B�\ 
������ /�t�RF"O&\[P��h� x�,=��9��"O�P+i,np����<���"O�4I�iÓ��2��\��"O�pX�m�c��l�B�U�_��4B�"O�`t�f��hЄ�/M��	�"O���F��^�
gN dz���"O������e-��OL����"OY�LШ�R1�凘�h,� �"O�0*���(��3G!��"(��"O�dwc� \G1!�m�		�5�G"OƘY��K�P�*����c	6�À"Ony3	��jR������=�dy1"O�-�FUV8�H�)�b�3�"OD��cdJ�~�����Җf��e�E"O.�i�!�3	����7��8� ��"ORyD΄47�4�g$��Q��y�#Y8g�JA�� ���dX��y'K;o��٘����P"S�N��y���+�D� e���x��2@��y���2��S��]��:���F�2�y��^b��ĢU�7"���Q�V��yb��DQ�!��R  5&�P���y�@�?a�tQb�`:q���Ê�yb&� ]�*�	�E� ,P���Py�&�:L��xC�!3�@��g"V|�<q�V�Xp}7k̔\:D�YBM�y�<�4B ~��Q��g�4-1Ga
r�<b�]�[�T��֠D<���G�p�<��f]r��f�
�cHh�Z�b�k��U8������p�Q�ۥ;SB�$6D���vi��z�z@��@�R�@�5D��9�Lvd-��KF�8{�@z�*'O�"=)�\�X+�u�Gc�B���ه�L�<�5�/D�q9� �FV �C�F�<�w�:)R��@-�-i�@�!$
�l�<a���'A���'��p�"��G!�h�<��b�?zV͙��W�w�dd���y�<AQ��F�Lj e� [�b��n�n�<�(�[�^ �aY��Je
�o�<�$nߌ���P�0��Ð"w�<���� Nk�hZv
�T,����|�<�PkՔO�!3"�ս{�x��WC�{�<�W�F5X���'*��T�w}��'[����.?Sg�}�ř�X�0c�'C��B��IL�:��Ҥ�=� `�'T�˥�:�f\cHƜI����� t0iwE�7}�ŀ��*�����"O��CƒJ֐3u��3~h2��5"O���*��n��C���Q5��"O2@�cA��=f�$�����_�1�"O����ƒ6$RV��cՇd1�y�"O8���A�����VYs"O�e1��G�R�R��W�rsR)�"O�5C��;�8���c�2\�C�"O�5�j�A*� ;W��#c�H��"O����L�A�����B\\�[�"O��r@��3���H��X��"O:ibt���� �"�F͉4� a�"O�y��]�1��91����X��`"OąJ��U �>I:R��L��= �*O�q�*O �5��ʞ�Nh�'0f���R��Q'W8?yX�'ѱ�n�8|f�6M�>i'�t�
�'Z`��l����X�LPc5�͓�'�D�K�%�=�|� ���T\r�9�'Ȁ�3fE�I�,�Z��=}2���O@��D�%W��p+���@��(D��}r �<Au�Ԫ=/�D��ƛ�\�����a�<atlL�x�$�Ո�:da6,�\�'a����n�4�P�%(��@,A��y���8tiP3��t)�=`Ԉ �*y�=�O��P�<ٴ�_:N<�+��^+G�<��HQ�<9	��O�&��ӍЮ#��)���L�<!Q��"h�,U@R��>_�a���I�<���M]�V��ÇR�OL�B&iV�'#axR,�l+~42��_ۨ�Q'�$��'����S)����iU�s�Bh G�W�cn��	�G��J����iWb��CS%,D��ڴpt!�d��`<����%� U	�
ԚM�yҦPp�����f����9��K|�pm�ȓ�lHK��׳	�l芄+̑)��-$��хW�ا�O�d)��G��?7��B�Q�BQ	�'t�(��bH��"`NN�i�h�3�IF��~�X� �#_
sh�AvA��p=�}bdȐXv�)`�����E�5�K��y����(�ߝ{&�Q�s���y2jY�a�č�P-¶s�h�Ƀo���ē�p>���W�FCxy�&+�6H�>����T�<q�ߖ3��!��R�nf��p�HI�<�f$��}S��A6
X;c�ȁH�CC�<���{����T�Ү^�P��3lF�<q�璅^FV��2�.$�s`�A�<���)�
����(|���e
FX<1��~��Q�c���3��d�@ ~�Ɓ��Wp�X��=5т�9�`�yX�!�ȓ-ǘx��M�\�֝��C�50�I�����X��7l�z�Q��׫?�|��z�2yH�#kz��QG
%4�<�ȓu�����]j��i�L"B趁�ȓf�[�)�{�N�v��+���ȓ_�z���:�he�L_���d��F!4� �l\�#��%�`��J�ȇȓL�������!D����NB�V�Gz�'NΜ;UIHF�f5ʶ$��c��%��'`�}�S�ͷT���C�ON' ��'��HP5eƒ#��1kv匱Ff6�
��M��{�Kۃr���G#ZdYE!�b/�y�γ3��Y� �5�~	#ӆ�(�'�h#=%?)y �9K� �6nL�^��"�5D��
�Oʬ�f<	�ϔ�f� Ћ��/D�� ֡�t�ʷ_ �3�*���V��D"Oj!� ��*`LST@�7sɨ�E"O4�`��L��ԙjZ ��"O.$y�gȑ eB�qN�6QD�k�"O04)�}�V-1F�����Od���]�� eʓ·�G�:T����:L��l}����m�6�����I�n�iQ��Py�jF�`)�+SM�Fe8���|�<	7�߆�Re�eoF�mPD��"F�Dx�l�'�dzA�R�_r�e8��ۦjF��*�'��:�뀠EGhc���%h_�ݨ��(�S�ԭƱ���eNխ+��*�d���y�G߬5v�$�Vm�+w0y���п�~��)ڧ. I�s�@�N��h���W?0p�؇ȓE��4���\ z.0�vh�`� P��!/�hH�B"wJ�L��Xr|iʇ"ORrL����s��бO�zp`q"O��S`��.�8d�Q��%� ٚ"O�1����\s�ܳ"�O�e�ZY�U"OJ`k&'�ޕ3�냶?Y�!1�'*ў,���4������V)u�	[��ih<	�!�p����]n�iS���W�<ɵ �x�ZB��62@����I�<Y�Ԑ<����h�0	���jQ`�O�<�b��v�B x��B��az�
�K�<�uQ�P}�I1��pdR�(�I�P�<٤���7IFU{0�Q�	����Gk�`�<�5eX>����bԑ9KƷ!!�B��:[�d�=+R��eI�aw�B�I<#o(��SBZ-������C䉷&�6Y+���)R�`�) �Q�jB�I�/��su�/Ϟ9��A��*B��(P�!�$��3�0�$��2��B��K�J��.S�x�j h�Z2v%�C�v ����.\�*���n�g��B��6wp���m]�m�
���DO��B�I�z戜�f)�(�
�U�RB�	�Q�5�d�љ'9��aa�6AB�I�y��Q�5[���QhM�C�I'�z�H�j ^v�sCB;W�.C�I.	{�L0WąN����"@Q./C�3@��%0�"�:W~t5�H�"��C�I�q:�Q�S�W"*`���#X+�~C�I�s���J<(����#W.4�B�I�:p�P��҈�D�ì�'L�hB���
�*�C� �����Ϩ>�&B�Ɉ(������(J�D��DG| B�I�S����)�ZF�<	���T]�C�	�8l�(�4����N���# �d��B䉌z@\ȸ��QT�*��g�4I:�C�	;<Z*mQ��W8r���%3OJB��&=l.���\&lB�a�ϕ8]�C䉖{���b�P�\�� ��,�:9��B��7X\��%��:��x@��N$\�B䉛G�����S�Wo��JP�R��"O4���5H6����%Ƞ"O�L��޼q(��c��N�54� "O��p#���!��@O�y���je"O��:�����X�[���4)��rw"OJ�fÌ#�eH�Ļc"-��"O8�p�̙3�U���e9�@3"O���T#��j�Д�*�)�M��"O�	��&�7G�H\���?�DA�"Oȑ�w,А�4�eg"r���I7"O� �IStD�r����L%R9�8�"OD�pl�
`�w�9]��F"O2a3a-1���`2����9�1"O��㥥�#�MF
'Y��Ï���yT7l�p2�����S)Ђ�y�L�,ذAG����z9k�/���y£T�h8�l9vG X�&���y򧀲�x��v��R��9�����y�Θ�q߾]���ݸM6N'����y��K�v����d#�]�V)ƀK��y®V7S�,��PA�Z���4^-�y��ЯC� ���&K�p�*S�yl�R�ZTq ��F��݂�����y���4���DG{�QS��yR� 0cj�J����YJ"��!�y� oU�Ɂ` �RV*�{�bB��yb�Q%Έy٢�[4R��H�K��y�nL]TP�´���3�&�z�M�y2FZs�a"Q@�:@�=ˇ���y�鐊��=*R�H6n�0�&/X�y"#��{��H�a�� fP�1f�R#�y2�KNQ�FH*{�0��(�-�y¦�%2�~�h�hR�T���#%ċ��yRg ��8�8�+ F�p)�̓ �yb�Y�V�l�#�h��Dl� aC?�yrdعq��٨�^5A���� ڔ�y2G�4�Ą@d�B,9
�`T���y��B�J:-S'A. .Y�c� �yRn]�"�1��H/Q����y2jǭ���ItB;,!z ��yr�˟�ژ0 aH��^�u���yrA�1	4T���*���A5��=�yB�G�5[�}�䥁�.5yT�R��y��^1��P"bL�;��((!���yޢ!L ���/�R_�trPGG��y�oN'veL[����gĝ"�y�hR
�yi�� �u�I��=�y� �����%F�3Ex�Z@��yr�U>J�Ҝ�#�CU�A`��y��7VXy�6 ߥi]
 �pM˂�y�b��|��3���
�(�y���j��a�*_�.�`)�ؠ�ybb�z�(��$F!8�2h�AɃ�y�	l=	dȐ�<�i��A�$�yҧ�>��%K��<;O�q��ܛ�y���?����&�)5�p%��jщ�y"Fg�嚢ݻ~��#?�yRbѮ�<��ka����c��yb%3 �=(��5�Ф�����yrG���D�-	�*�C凫�y �W����g�4/�Y#v�X�y�ɏ�N��J�=�D�VF�/�yR�K����#O�9�.��B,�	�y`+r#­���7��Xb���y���;
��[��
)���˱�y�ƈ�itȠ�6kզ��{@ē�yi�1\�Fԑ�F�'Ȅ��F���y"e�>Qc�,��'�L� �p&X1�y�֚g� ��f�yNhP5����y"��S�h̸�mP	)����&X/�y��μQ��}��l��/�*H��?�y�"�9|�r	zA�Ya�(���T��ybO�2>� �1@�Ț̅)���!�'�`�8q��r<@�3hԓ|Lu���� i�������'�%T�ਜ਼""O*]�4�XmXЋ(�(#��( 1"O�=rgQ�B��`R��V�t��"OT�	HY(!���x�&��}P:�
�"O�ݨ6/��b4���e�!Md��7"O:m��[�B��Y��$�:	ZZu�0"ORX �j]�;k -3s�
3C����"OF���R%H�� ��5Q�����"O��Z6@D;*c��sCٓw�Vي�"O(���C�4D��[�߷ĺ��5"O,�b�Ę�d�z�cĮs�ް��"O�9��?)&h�o�B�r)
e"O�a��#�dJA	�C��Q��"O4���I�l;R4p��@�)g41Kv"OР˗��� PR�q)J5rx��6"O T#!j��@��	�M%�Q"O�$�F��iN�-���W�DΌ��"O��@቞�bL� �uJ�0 ���"Ov�X <Q�<�S���a��"O��c%ϖ<TSj��e�J�]o"��"On(��$�r��	��f�PP�p��"O���իG**@�Pʤ�ڠ7Lq��"OX��H����Â8-$<Ҷ"O�ɰ��@-1q�t�؃1ʉ��"OL0SNU�O�9��K�P���"Od�S`�g�r�C�9㤽�W"O �	Oo~<�eD��6��%"O|��2��'��m;3�e�IQ�"O�KWd�m+��c�"3,�P�6"O:݋d��
�2��$=h���"Of����_Ϯu���Lg�>(X4"O�� K�T�P�j�я�x�hE"O� ;q�#�<��#.�$A��"O������5r��X�⊃)� ݩ7"O�(�S*X�6���[q�Xv"O��H"ci֩�gΊ��x�"OD౰O�:|�X=�F�HGӨ�r�"O�9�T�,��C�I�c�L�1"O��ɖ\�$�h��7���cF"O�����c�t Y���4L��዁"O�1qp��H��i�jug���"OVTrC��E}�rRdΡ1�L`�"Oh��Hȶ#C:I��{p@��YN�<��J�3|��5�rg�/KB�t�DK�<�Q�N�7�LlQ�ˀ'�L�8��J�<�dӊ]	�K��ͽj�дQ�@�p�<��+�0:D��cFc�21�&��6FC�<�΂1R,x,��5P2|D�QfTi�<!2nG "�]Xu��<�.�褣�b�<�5o�T=^P��g�rb ���^F�<�2b�F�d�sEV�9��B��\�<��ÃI�]� ,�Et��1�
R�<�A�Ԍ�3D�';���!�!\S�<�!fQ,P(;�e�,z��}�⌒O�<�tAF����g,g�XY��F�J�<i��S�9dhuI�+ ��Õ�K�<e�
]���k"%�0s��c��B�<Ya��9P�-`�J҆cEҁ3&Y�<��!�)��Z�gV�h��%SWJ�U�<a	�]5Zɢ�L�5�����Q�<�u�A m0���2���bU��G�<A��	mUM��O9M�|]��$C^�<�3����|�rg�3���@A�]�<iNN8iU�bs��2��Y���V�<� .�7�7Q�D$��̈��(ܱ�"O>��4�~t>���.a�5"O�������Ъ�L]4���"O<J������(���F�i@�"OX���"K:ƀi¦��,;.t��s"O�q���ˮ^c���S���zhk�"O�hS�+XW/��ZR  E�n�p"O��Y�A�hڦqKsn'sF�Z�"Od�p"��7Ѽ!g���>m�\��"O��1D��(VV�X Ð�FM$t�"O��CRbV�K�Z`��U5rD4�	#"OxL��m�<Pk��{B��Q:�p�"O`u��i�E�F���P�m4��YU"OV���&Q�Xa��H"H�X	"���"O´Q�	��!��i�,��#`��"O���H�I��5[��R�>�`�!"Ol{�,&AH�0��-�^��"O2c�	@���z�lӖUk4��"O�XR�.�Ut�I��E�mT���0"O�-q5!�,Pêِ��?H�K�"O��rv��=+~���q+�3d���
�"O��R�C�k|xsI^���"On�я�5wy��dU#K���"O�E�d҈X��k�m��'��r"OTpj��F=��Ss#�	��l�b*O��Rg`�;����l>��'a�0�����i��S�����X�'y��x�����J3Ú1%3�'���`B�S"%�Vd��ߖ��K
�'���T-p>�U�Dˌ0^�P�	�'����nF1F}��q��cp�	�'S(�$I�rp��f�D���	�'�V`Щ��S<>H�f�GZ��8	�'���d��JP��+sO[>j{�[�'۰4
%P�<�#C�[/�4��'������]/�(��H�
DX��'X�H��̽�$2�H�9B2�:	�'cbP#&fV3C��d�D�`�����'M�}R�G\.���G(k��X�'~h	�e䘤��a�%Mrn��'���K�)"qx4��퇴}�0��'�VibC��aW��ŧЯ ��A(�'
~��B�25謍���<
���
�'�hPh����j$���J��
�'n̸���؜)
�=0���U��@

�'��¦�H�5ZvpVa�/Q��-�
�'R����-��\�FҮ\��e�
�'��(�0�Xu���Cp��	KHĹ�'�.���!��@>j5ے��a��	�'S���䂈*#����!jѧt�nX	�'Έj�ǃ�J$|}ဍ��j�"�P	�'�R��F, ��b��a*��Q�'`X(� �]/|�~�����n5|��'�]Q���s� ��
�_A��*
�'3�!���*cn��p�E�!���	�'�P�C��_f��p���D8�b	�'A "��RI��4����:m�i�'�� ի�
 A8�v��8Vl`�'z�HJ�'��n�˕���:O�I�'�< 0���,�����1:��
�'X�T�$�ʇ\V�i��Y�1oj��
�'���3���̒iqK�l�9�
�' ���N�(r��b��,1
�'k���J�A�:m8���"O� b����@=tD��� �R�� "OfDy!fۍ �%Z4�Y_X�<*"O8�i
F1b�`u��<��T"O8| ,E�"���OY�j�~Ѣ&"O0�Q�[��zcѯ�� :�"O��(Ej�?���viֳj���t"Oҙs�A�#$��\����4I�Vyv"O��)�i<-.T�R���+0�T�)�"OV�B/�-Mhd��b�N�I����"O�`��J�(O�~���B��7�҄�P"Ofx�w���%�b��2�8R�"O2����M c>�(���5���za"O"���e�4Rd
���`-f%i'"O�mC�ᙳ626�Qa��;f|:g"Ohݘ'#��-�5S6n_SX���"Ox쯚<Zr�`C3$�*���H�u�<a'����H+�KR�\0CTo�G�<�' ��$��`�mG�+��j�HZ@�<q��ϐN�	!M�F�r)�D��}�<���=Lf0�@�eC�6@r@X0��|�<	�O���(a%`�h��v�}�<�'�ͿD��a���W�?\Z)�u� A�<���Hy��i����6=iR�4N�d�<�a��Fi�bk��j�����d�<�L1QRh��C��k�J�d��G�<a���G#~�؃A۞r��S1ːC�<�a�=>���!�������@�<���d��$�J\z�� %�8D��2�#Œ-��O���yS�9D��nF�Y'<hS'G�I��1#��5D��Ca	�Q���RnF�QY�҉5D�HV�ތJ ����X*��3�1D�dۑ���"װ�rqʖ��D���2D��jV��_\�[aɓ E��4b�I,D���6�݄y�n���g�.
����U,D�8H���2�F���.Jf,q&�(D� 1CY�<q�x�5n]
�N�( $"D�H0��H�c�\z2O�+�H�#U�5D���E�h��sց�-d &@
%m4D����C�;z�9I�N!+2���aK5D�<��V<��Q�=+�H�K&D�(�.^�.9*�� ,д	n�${Qf%D��T�F:�vy��g��=�,T�7J$D������f�B��[!�a�*7D��e�H$e.��b�lZ�+��9rO5D����F@m�@!cӤ���D�/D��j���i�Ph�W�ծo���0k3D�8 a��-BޡZ���P��4D3D��I��"t��,�.ؿ'�>��r�;D�$z��Bu�,){��"��\ZC�-D����I�8>6ب��\�@�Ĝ�*D����쌟5��:�l����LxK&D��91%
�x_�h��×�;�`,��(D� !DbE�s.��.ˉ�n��',D�����Y��;qN��5�X�(�h)D��+�I�0�2\�!Y�7�z��%D�l��*�X h�D��#�jͲ��$D�J�Hg�Բe�*~���F#D��Ӗ">e���JS�؈��$ D���ᆒ8�zBD��u��꣍<D��(&�[�R��(�u�W95A�����9D�h���pn����W]4��L3D�Ђ�ԑ�Έ`� T胶�<D�lGI��2/B���D�;0h�`/D�� ������l��5�$��8 2��31"OL�a�hԹ+Z����M�:�Zf"Op��ѥ�=GԀ�MT2Qa\(�"Ot��pg�R���@�[�VD;�"OT�"��&��pJ�Hy6ܑ��"O6e`��q��� ���"�"O��t��0X�ؔӃf�"M��Х"O�a��#F�y~����ӊ0\U��"O�e21�G�\��!X�L��Kf��1"Ö���ֵV�~y�f��& 	�"O\E ��&䊭��)^�J�T�"OR��/�Y�vkS�:��"O��`n�!�D��F�K�v:c"OZ9�M�_v��u&2���*W"O��aVܔ%*����,����"O |�ЊN�≉E��t�
��"O��`�F���丂��&O���	c"O.��vH����Y�d�h�R�"O@�M߉z" \��:u�:�j�"O0a�i	�|4�S%��o��d��"Ot�"�%��y碸�N.h�8f"O���B%��$\��pd\�Dw�x�"O�u�UK3�H�2�ʤZ7j�C�"OI*%�tg8�@$�X>�*��W"O� ��� 3n�%3lZI��a'"Ox��w��r��e[��K��1t"O^:�

M�+e,�1=��8D"O��V��
����q����̒�"OBi�Ջը�޹��i�1y21"O�Xp5k�& �� vi�l�a��"O���!��3h��[�b!jF�k�"O^��_
����T�0i`���"O��#ȝ�AϪ�����>e��"OD��C�)nc@qPP�x@����"O�|H��J� �6�ibCY8a7\I�"Ove�ď�+\�v��GJ�&�܀ "OlM�r+�0�R܁!J��#	���"O0����8^��O߷Y� 5"Oz��R�����1�( %�%+�"O\;bc�{�|���˚�n��� "O��Y�.![��uj"y��Tc�"O��B�(]���s�H�5�!s"OܕS�"�Ƙ,�6#<X�αʑ"O�l�5kR�%��!j���I��p�"Ov�[���d���iwa^0���r�"OY�C��>}��3���c���)�"O��r杨/�@���9�T
�*OX�2�Z94�hHa�1fdj}:
�'�X�bi]Eu�0;@�q��h�	�',����W0!:�̿mq�c
�'b���� e���@��O��Ī�'F�H�wQ0Iȭx�lϩ�<���'��X:U�Y YX �8��	bF{�'�p��'T����4%D�k�<��Gґ��� h���	'萷Zl�Ņ�r�活!�E�J�y1�T?M�2<�� ���j��E�i	�㗀tx:��ȓ5}��B&&Ʒ.84����>��Y�ȓ�L飑g�,!z��-�E�^��B0��cF�o�������(ȇȓ~X��Eɱ
"�e�#A�&��-��),f�G��;	��0y�FS����ȓC�H�a)͉a�l( �� ����R�XU(�H�0Y�n�(�O >R��ل�S�? �q�`�V�%Ɗ�A��@��f"O4Q2�:L����&�9	�.�"Ox�
q'F:
MFH��EH��9V"O�%Ic��o�pD���C�0�"O��B��������2��%�:Ls"O�����ڲ��x�b��I]v2�"O��`%�M�����0z&UIU"O\�A��%'<� !��X��b"O�)�K�~D1�q������"O���"m!Bj>�Kƈ�B���"O������8��t�'�]�	��"O��@�&��q�Vf�,`��d��"Ov���g@�9]����Ō96�d��"O�Yk���]N��V/t��)R�"O\���B5��HشBE<U�ĭ�"O�U���B#,��(C�P7S���t"Oz�9�ɞ"h�I1`�W��F��"O��ȒŐ]jNQ[6O�  C"O�ѻr�B;�2Q'��j��Y��"O���B��q�Xa�>E֢�C"O0-���"A�Z�H�
�;6|D`�"O� �"P/����Be��Q�"Ov<a�K�*��̐���)|M�`��"O�L�����p� G?��c!"O�����,��]1���O����"OtȐ���D�n ��I��n��b"O��=?�,D�#���0�"O�196@^�H��8�'�f�,�C"O.��%�K�M�,�!������P"O�e�"��.�t[����`k"��&"O 9���0�<����2ck��� "Otq�w�ݝQ��
P哷ky����"O�Up�ڴL�9B�Q�+rpT�"O��0���os�Q�WH��t
�"O���e�Y,@���L�	&w�qC$"O�(Cwh;�D@���!��X��"O\M��K�T��F� �\tˢ"O��j�{ÐL���)v��ٓ"O��C�**�EA�`٬z��a"OT0��h�9&t"�R�d9��5"ObH��j�h�å)ˈ ҕA�"O�hk�JX�֠0@�U)JY#E"OxPS��Z9:�N1;aO*�����y��Sj8X��.!\��Y
�!�y2��,T½!@DȺ\�Asf%���yC�M�����O�P���Q?�y�J�!�4���$�w�X�1U^��y��7���/�8L�w���y��Ư@*��1Æ�t,8�7��%�yRK��`!�&�B�m��3�Ҋ�y2�ݝQ\�<(्�oz�r���yE�'`\��eI�/��1��j&�y���U�h����#.:�x@"���y��)��Q�
P=,_�I�i�<�y2�M�SKt=��C
!��maf�^��y�l����2����
ϰ��"�ͩ�y����<��Pp�*��rh0���!�y�(��j ��fY��A�"k ��y��
! �ȴ��{���r��yaõV!��!��Ü^����'E��y��%"���N�;Q�f��a@���y��4�l�Z�)ƯY�h0��)��y��A'p�D	�O��3P���yR�� ��p���B�JoF�`w��-�y
� >В �D1^8��vꈍDۊ��"O�L��F�GC
��6'��A�0-�$"O��B�-eЖI��k��2͜D�w"O<�ʒa�%x��Yj5��_+0��"O���#.}@���p��c��V"O�h���ƣp%x-a�C s�ZI�"OZ9S�O�vLM���C�� "OT	ID���}����P.W�Q�Q"O`̋E��$b��U���-:���0�"O��w��<���69TFuB�"O��!�lIͪ�sD��Q���"O�m(A�ݥ|��Rf�;L�����"O|��Ǌ$���!B��lz2���"O�s�^!k�ũQ���H*M�"O\����*s�a� σ�Zk��W"O�1kC��)Zx��,cw���E"Oj|d[�|��0�uh]�
Zr��"O�hҋB�*%�PӝxITA��"O� �͜�c
;��0>�J��E"O^b�k�/��ԍˣ;8 �: "OF��P��3q�V̚6+P��"OZ�QU:�V�:6n	%]�|�a""O�P���rʌ�6�J�:��"O\	L�RQ�Hs���d]�u"O����F��9(v���kD�N��B�"O�ip&|@2��C�����@�"OQ��I-F���'lSA�PJ�"O��u��1]�݊����k$�u�"O����#
�-�&D8�@)6 �b�"OD��F䓴�B���M�D�z�3
�'��1pцLsBp+# X�o�4��'�X8��]�:�`�hbh1w�5a�'��@�b_�Xq��O&D6��+�'�����n�l���b��'¢���'��1	�^gEd�C$���;�'�H� �%[B��
Q����P��'!����a���! ��6�Ju��'��s�nJ��0�)S�0���'lN8	Bj�-3@R�9ֈ�=~4�1��'9��JŌv}��H�5`�v�[�'��	��˒F�8��C��S^e2�'Vxr��@�8<�"\&Tɜ}��'���3��h�x�p�˙�E"\i��'肵Bc�۟k����
��	�'}��C.ay��7Iդ�bp��'^���F��:��fI�-����'m��Ha�¿:qV;&`
5�8���'A�q�V�ݕKH4�+�/t�mb�'?4e ��۞?���b��_;z���'n0�0d) s-�����X&�Ѫ	�'�H�(�
[��9�dˌIA��'�t;�"�VKp���C\(�0�'j�E�!�*����WE��&@1c
�'SF�U#J,~X8`�Q�A+i�T��'�n-C�ҟ(A���i��'������5�dLs����t�R�' �t{���x_0أ�������'�N$[��@-ir�A@ׯ�}Ů�*�'� E�т� �s�/�4oܢD��'�&�ۑF������LKt���c
�'��QO�+>�ր�!���]6f�i�'��H���V�lJ�p��,*���'�4mЁ�݉V�����=)**��
�'����%A?$T��eL!%>l��� P���,�|��B�&$8�S"O�X[#BI6>�����NJ��"OE���L��у� 1:�2��7"O���6N�v7�$IT�xp�"O	�@F*!�L"�&��I�XY3�"OFȩGNF���Z��=jk�P�"OƁ�햒H(��Y�k`���q"O�DY�d35]��bJ��~��"O4�9PMwpA��&�*.���2"O��!�ډj��ukpY0�:���"O���!?L��%�R1!`zM��"O��p��� BPm��ǢDk�d��"O.TQGeGL�������x1!j�"Ob�y��2���3�F3?��@�"O�$bMF~O��ڣ�����I��"O�Щ��Q>��=[4
L E��ɱ"Oq�3B�q'�L�|��,�v"O��v��5 ��|�r�����"O~��g����e#��7켝�4"O������$r�tk6lL�J�@T"O���F�T��̩K�5�� "O޼
WB�.^]��KۖwH�X�"O8��rD�1h���B#��Jlj@"O�Y8c&Έ;��"@��ЩC"OL�"��G2��`\
n9|��"O�篂'A~�:
��h��r"O��aFM$b��B�H�>���(�"O̔��f�9oZ4�-B� �4��"O�|��ՀW����h� #c"O�a`���$oP��4��M���"O�񋧌�A�p�caG_��d1#"O`) ���%��0V @8
��J�"O6d�.-&A7o��@	aU"O�%�����42�M��kE,z�Н��"O�a�`��`X�;#��0جM�"Oj��e��]�Z�@���(� "OY���._��@�3�īz6�J�"O�){w
�_c�X��/F3t�4�"O��H&�:*d���&B��g"O�,�k3��`r�?`�F�g"O�i"� �X�Yw���T���"OP�ѧB�}��ٳ�,�"EL~�Y�"O񈢀E9J'f�<Q�C=0 !�\�#$^�A3L#T��� �B[� !�y���t�Ȭx���U#S��Py������Hud̓-)$Y��:�y�P7\Z	zWoׅu�D�J�&��y��Y�iR�ɤ�gNL��ʂ��yA��_b�e�E�A���bg� �y�Ri��|3�K�
����ūL�y���t2��%8-jT}X���+�yb�7n?N�1�m�$�P�`�O(�y�ɔE����E*�RQ��*�y�%�+�8�Kt!(F����e���y��G&��b`�>{�����Ȇ�y�0nI���oA7qT��j�)��y2�G�M��Ӱ�ܱ`��y#è�yb@P=P��irGC_��Z������y���:Z(�휘T�(�R �y�@�8pĠ�[2��I0���6(��y��VW̮MB��Hyn��c�֐�y�ß�J�t(�RȖ�J�����"
4�yr�ƳcV��V��y_\��6��yr����HcZ�j%P��M���y
� ����.��&]bt�@��\ic"O,���3���%H� �`!"O@}��F��"�ޱZ �Y'���D"OJ����4U`(��IS�&�� 95"O|40E��Y����)�/Fh<�R�"Or�å%C�l�L���`1�<��"On�`@(ފ��s�N ��T�D"O����Z�S�ā���M~�S"O����.�?�)�פD�tR���""O��e� �%B��s�b��#"O�飄A<�2HU#p)�T1�"O�ĪR�,� ����X��� !"O��C�%�V�� ʋ�v�a"O ɲO�~�kCXttJ��"O���C�_�±X�DA�|e���"O:}�d�:�:�s���S�|x�"O�X�6�W�^�`�)%�~%15"O�<c��Ę X�(�Bd3���j�"O���Ã��	b���㛆x�$��`"O��ڠA�/bXd�+'�E���:5"O$I��l)����>8�� @��y��E x$�IӶh�DqO��y�S4a�ex�&�g��Y�����y�*����S�Z!��p��yb���a5��amL1�,S��^��y2h����$ E�@&Z	�rD��y�LT�SB~�#��0��J�yҬ�	Be��a��J�f��Q�)��y,Ѿu2.�s�$��X���N��yR*�;	��m�d�^;	��(;p����y�cI�H����C�μd:/^9�y��מݶ5�#�-
�%3�釪�yRNE�6+~M� ��(rڌ9��y���5k4��� i�8\�� M�5�yR��Np����D<��{1� 3�yMx�T�Å���k�<�ࣚ��y��@��E�`ލx���q�/(�yB%S�_������0x^uZǏ�<�y�`<� RlQ%�v���Ȑ��y"��2�,!���f&�Y��?�yb�P8��p��._���a��yb�чKQ�Q�`A����Ȣ�y�$::����`�V���)�j̷�y"$ֈr�;#�B�����2�y�)�<l�|ٔ'ç��x�!j���y�@�����I�C^� �o�"�y�	4#��0&Z4=*̹�ԁ�yrG_�It,,(gM�+Fİ�M[��y�d\Iz #Q#��Z��yqi��y�G�b���Hݥ$�^-�&
��y�	?I��IS��w��`%��y�
=z��1&H������O��y2ғ�49o��0,0'���y��^;P�H�o	��9��Ш�y"
ߣ!�2��oQ�T9�(����y�@W0e����J��@=�1@��6�y�B]�/hHM�vK��(ɎdX6h��y�A`���Ӥ��"��|�EkI�y2�� Ғ�7Ϗ'2e�̡��٣�y�o
�
Q`u�)a5v$���!�yO��1���\�&X���v�+�y�(h|��P(*@��Kv*��ybFJ�XPv1�	���<�ŦT��y��M�`������tY��$��y
� �X��c|�M˥MK<@l`��F"O8�U��]���$nK�O4l�y1"O��C#ΨO�8!�d̉K��(H�"O��(�ʍT��ȏ%�4q��"O�}�A�k��00��U�Nq�@"O�@"K�1��H�$=q�-��*O\	z"/J�_rdy�=S��0�
�'>����#B	��a�͋Ehy�
�'���R�]i��K��.�q�
�'�m��b�K��h�̚�q�ʱ*
�'��A:��H;"lt�"��T��t��'��E%e�9b��1kG�;�Jt��'GFl�T֕���������'����5��G��c�M!���s�'rP82'D�ބ�"Ý�#�
I8�'�>1��A�eX��q̏+���'%��*��P�
7t�i4��Medx��'��ҕ�?*n���d�-sz���	�'<0X���<x�ܤ2�ˤY��(:	�'`�dK�H0+�X]�A"LW����'�H���oY�a'2})!��R�MC�'(�IY�DI�Q���ra��2p��	�'�D��v
ٰk��idK�
)#�d��'�~��W�)
�����w9RXI�'�l�(��ĩZ`�Q&+W_K��r�'�ٲ�"�*}�BI^O��� �'��\�@G�<P����"�E�����')�%1��:ҍsQ�L�Fʚ���' ��ဪ�4:��ؕ�S45� I�'��yj�ՙxȆ|+� O)O¨ �'�x�:��?I.E�������H"�']�Lg�J�(��Pأ+ڮ�,u��'u��7!�!ĚL���
�=�5;�'�\aÁ
H��K��S)wx)�	�'S2�*�N�:��yA��$=2b ��'��ujp/<���(�aD�kyx���'Ú���#G<i�R(� ��������':P�F��1x*h�����'(O�9��'�n���-����M�&+�U��	�'�b�bd� \�2�x��������'�2(#�⟷i�j�I���^��A��'�V�9To=z0+f+ج""�k�'� zf���Y�j�9e���ཡ�'��ق��hA���%��l:>5��'O��!���w�L\y��5�0;�'��[UŅ�4Q�0Jamƽ4ܸI��'+�HIeE�+�^�ڡJ��+p�d�
�'ްi$B=�I[Q�
*P��

�'|�������V��FށB���	�'�<i�2�͕ߨ�@u�$=��`	�'��\��C�P&0eOS4]�
�q�'}H��!a6%�p���d�W���R�'ߴ�H1�P0����7��Ulz���'��]#��� �>=3�#R��-��'^F��L[�xB�hR-LYh���'_x�h�/g4�b3�D�o"@���'�aR1�. Vd�3���li�5#�'`��e�Lt��s@�D�a��'iq:��_I�ԁ	��@!U�����' &$*� ^B�a���Aa�Yp�'����2��v��x����Dyx ��'̓�@�-�Z���N59�N�c�'�|�蛰R��j��C�6R~Y�
�'�Xс��ƪ<`�3�lڌ#:�I9	��� ���5ϝ�[���� W7
P�x��"Od����\�F|�u���
EJc�"O2���Q�}� �Ps�J7"5"��C"OV	`����l�8�B�!�lQ����"O��@E��T�^-3A�		i.�b�"O��PdjљYHȨ�Ȇx"���"OX��lS�ƹˑ�D�x�Xc�"O�y#�F5q���s�S,K���"O��4��:}XUb'E�?]~�1�"OdDC��3���i!D�!�z��&"O�Q�/�c	�ɰ�`��*Ŷ)bb"Oj�H*�Wl�|bƏ�~�a�"OHTP�@�%]	�t�`�ZUv���"O|jdO�},R� �5��  "Ol�A�&ˌd%�!��P�r��9r"O>0���J$&#�g��X���t"O�((���	0�!���21&��¶"O`U�Iƴ50$9��R�P ��"Op�U�U�!;HX�p��7�
��A"O�pf�E�@��9 3dXC�8e��"O0�@�	�ܩg��7y�Xځ"O�#+@V��*��9���"O�8�7��aLb�(;A L8�"OB�k��;��9��3V��(�"O��au�˓j	z��e'B�-��"O�q�f�Ɇ=�q�S�'>3� i�"O����c�Mp�[�&®U&�@`"OF�J�/X?-�ܤ`u��; u�yA"O���#Ä~o����Iy�)��"O~�@��:e�K�ƳYw����"O��ÍI����8%A\�s�4Yi�"OH�9V)�4T�:�i��\�U���R�"O�li��q[bL�cm���Z@XA"OL	�F1�p-:�L'4��2u"O�I6��!IR@pG ƥ&��t�"O�e��ßD�N9zd �b�>�Y�"O\Z�AɷE:�P��-Hx�%7"O�d�&���(�#�Y�xT"Oxȉ�ȋ�,;�"B9V�p"O�tőK��Y���+O2�e+�"O>d�C�1*[���@��c+��1�"Oԙ���ҧ0�,X�o�Jn���"OV��=/�h��m�v;<D$"O�lx���8�<��L��b/d}	"O܄yp"p�(�,!H�"O��1�ՠf����_D�$"Ol!���r��;6��'���"O|��SJ]Q��l!C��5)� �e"OV#Ċ�3��q��"�
]� �SG"O�ls�:�������'[JU[�"Oj����:Wh���ӍS1��Ö"O|8W�O�ԑ�́,Z"���"O�d� hj�xWk�u��`"OT�ؤ�^#%NB�A���ge���4"OʴP�Y7F	qU��V��K�"O0q��A�6�@�pu� �>��"OT��%T� jp=�UO��{%:�)�"OH͑�%
=c�Z�ك�^G� p�"Oy�sM�#eK�ۭ.M`H4"O�eco�)�P�A �mI$ 9�"O��!�)F=y<� �۲9E�Ց�"O]�ş�[��ek�.�vΐ5��"O@�6�X�rـ�MT���S"O��A�.��alb��� P���#"O� ̡pa��+!l2=� �b�"O� �1đ4����W�|�f�:�"O��ʦD�&a<���Giڲ�.8��"O*Q�O��U�'ۘa�
���"O�d����7w��D��&rN��"O2��S�[��E�N�taj]�D"O�y���ٞ'E��񕦛;}P�S"O�1!4Ϙ1,����$V�T�^L�6"O|1�4�őK���pv��9��"O� ��K\}Ը���8PfJ��4"OQ{�N�Q�t�@
��dg�հ"O��1�C`�����<t}^5�"Oҥ�C�5>�0�`��N &h���"OH$A���f0�� �zO�,�"O����׽</~$�V揗_����"O\u�5LF�F��}�`%Y5Ρk�"O�-�%k�Od�ҧ��R6����"OF��*C�5.�eQ�N�%4'v�)�"O�9WM�f���	@��.��X�0"O`��C� 8m�Z�X�-�#a�r�8&"OBɘ���XQ��)�m�c����"O�4'w��A�F
=#�R {"O��q���}�v0��?F^��T"Ob�J���P�mJ��U6$:�H1�"O���f�>�N=� M�f3�x	 "O�Ӥό�xH�#��|&�9x�"OZ�E̘,P*��#��l\�"O~=���D>Du�siTiI"Op��@ӷ	�4���	� N��"O
���Y�$(:�@�]��"O�3�Z�!�Ēc狏n��8��"O�C⣜$s(�)�:~X��"Oh�8�g��<e�Ȁ>B|���"O��4��<ڸ��%*	�5H5"O����7]���#V�L�R�b�J�"O~��p*΁g�������:7u���%*O����V�*eP���4��{�'lp�pah��C�^t�B�+M��'j���ޢ's>�x�aҦ�f�K�'9N����"|x�`�놩Q���'K���Ō�?�T��ː�pW(�:�'z݀`���o�������4�[	�'�>���9y��y	ĥ��w��5 �'`9*�-F5
������\��
�'���P�Cݚo�$-�"m��m�P�p
�'&����㛊{}��%d�	P�h��	�'�Fʂ�M2��<+����:�
y
�'~�tѦФ
Ő�*ٗ3�j�h	�'�(LL�3�U�H�&��y��'�z��e�DO�B�s1	�"^�b�'ʹS����d��7)D�0#�'��`ڗjA,rĂ��̴AB,#�'�$�k�'X�j���!(��9���C�'J�A0� �nS6\ ���g�:�'�a��
C�4np�Ɗ�Z^ha��'�V���A%�N`�Ux�ѡI��Py��	z�"��Ki\�vd�u�<)�'�yBX�%��"V�i���p�<��+@:N��FS�jX�����i�<�'�Ҩ5�,�ҕ\�Z��$��g�<�T`C�_�i��e�8��gQM�<AtK��0�hIY�&Q�K��	uRF�<���ԭ�R,y��/Wfy�e�B�<ɰKT%^�N ��	)i�P�`�}�<� 4�*)� h�$�"
ćs.9#�"O�	qbH6 ��̣�(�H�.xS�"Oj̻�J�=w����f�nu�tJ4"Oj�3�$U1M������Ouab"O��UbF�w���2h�8�R�Q"On���1/ra�l-c|���"Ox�r(
D8l�LV�Fp4�"O�(�2�N�{�P=+g	M$p>���"O��SS^�B*"� dkɵL���s"O��1�.�L䊨L�~�jdY�"OL��Ơ,u����T,�qT��"O�e��dKT�p	���N�`Y�9C"O0���^z��+�b�d�E"O��P��1Q����kھݞ�)�"O|ɸ�&ѝ+�$�v�=X�B�ٓ"O�a��A�$�� V��^m�e"Oh9��X (�8)�pOށ]RnP0�"OΘ���4`~��Z4H�G*�k@"O~�HQ�Co�$���f�7)5t�"O!yEeQ�u��9X���"d#.%��"OH-0���J�$}1B�͟���"O��#��aN\�y��5t�l�"O����M$$���C���$)Bd��"O��J%�ɉ�L�@���^��%"O�5�U �,�)�(د) ��z6"Op@NH�(�d���hB�QCd��Q"O|ha�ן*��͂��x*��;�"O�4�͘^�6��'L����"O&��Kٰ0+F��l ��w"ON-`��j�B�*!'W,A�>��"O����/n�*x�GeB�#��e"�"O�A)�OY�(�K���AP"O�%�CB�]�P�v�L=c�����"O æ�[C�H0�`�[���b"OF��sǏ?Q��Œ ��t9����"O���])���A�\�R���J0"O�m��iJ�=V�LK����q��ّ�"Oz��r���nH(�/y2�=�"O�(U�X%iHV}[en�?�	w"O�$`�d8Tx��#&n�T�8�"O�@��I�7�*p�ɺIݼ �D"OҽꖃU**������>_^t!�"O����[$F���2�j=S�ذ4"O�p��H#`{�)JP�q���h�<Y�ڙe�@�R���$G0(����L�<�qM�@��`���	&m��Z���I�<ac@ɼkc(h�� AX���g�]�<!���
�2��B i���P��Tr�<��V�̺��2O�}�hȇmFV�<)c��p�j�H�,`�X�R�<I����:��l�Ģ�J���s�D�<�@*�<�4��LE�[�5 �QA�<���3oP�2@�L��!�y�<A c�o�HȤʊ�32����x�<i�.J
����ޅQ��i�e�y�<�g�A�B�hy� ��@����T�Q�<� ��21ND��h߃b�� *W�<iCo��N��(aDD�z�\"0n�T�<)�i&I�ɺ�ϋJe�u��I�O�<i��D�h���R��Ll>�jSK�d�<�r�T����ԉ�u��'�K�<�&�q4�aԈB���h�GH�<�mL';r�}�o�Q����t	�J�<�TJ�CNxPka�u��U��N�<� �`A�Ȅz��IT��' ����'�.�<aP/8
A��R�̀��E�z�<93�D�FQh�0�-
9S	\!Q��y�<����V��c�8f���0�I^�<��,Z ������� �J�0U,�U�<Q$��:`@�a� NJ9(�D�ҧTX��Ey�&ך6u���$�i^N��n4�y�*�j��� ���d���ᷯ����O�~@��u$�+TdX�P�I"T�I�<9���v��\�󣍩Sj�8��C@�<UJè"�p�sRMإN+L%�1D�|�<yp/�?\����)ԤC�0�`�y�<I�b	T���k����0��4@�~�<�GI��V����1r����bL|�<y��F7�2Y @�T?K�n�2���m�<��G�T5��"�{]#�P�<$�5���hֆ�8��3��H�<�w��CQ$�rv�)n���+�M�<�A�K�v+�T'��J�����KM�<)��ɑ.�Z���I�+d��OYE�<�c!G��8���*��xq�A�<t@0N��������63�l�d�E�<���5�֝i��X�����j�A�<��b»7��� J,@:�icL
w�<�2����@AR�*O�(�v�q�<�"��,VC�X����</l=�qA�o�<y��ęVh~� �P�Aw�m�<A��O�i���ѣ���8dYDM@�<!�,�=B¹�`�ܖ5@��U*�C�<�����Z��x�6.��~l�T�"DV�<�f`�WL�d"��$)�d��l�<��jq�$iq 
8n> �FcSs�<�!���a�^���e��Jp|x���u쓾hO�OS�Т+Ƃg�fY(��V&e�J�'Uў�}Z&bO�2�K��H��!r�,t�<9��W:a_xe����6R~6tز�Oo�<Y�֠E�x`����(3�����i�<����	��0�����#��e�<���V0h����B��e~ȉ����w�<I�lF)>�mU�� Z�<ۆ�s�<��)krZ�r�G�3c[xA0EMDX��T�([�ޟ#pYZ�* �NT�4D���޿\�� ��Ü�,�T�s�4ړ�0|��Mf����V��]�ܥ����e�<��Wk��y;5Z�'��x�p��m�Oҧ�g̓2z��`��بj��Q�Ө]w���I�bkSg�� %��q�*!��Oɳ�y�f�3V��a���l�:,Rg��0<���D�'P�(��c��F�.H�F��&U!�$�Vr>5YK�8��,k0c��w`�O\��D�Aa�l��D�.x�du��	�<!�$D�z70lBC�N�cX�ۂ��(b�<��ȓ[A��آ�y��H�Dr�D��Ʉ_�4��<!�����Z@��T26����䔪��'�az��B�J��q���]���d���X���M���imc�\��ŀ�|��Ū���!��-T�����.���aC��v����Ó�ŋӛK�NC�G��8�I�d
,T�4{ L�V�DZ5NI�PNv4
�'�!�d��<��T��B�E�ĭ�!hqOdO�}�v�S�Hd��5���*� �5�A�<Q�$�3��1ө'F���@�f�}�<a��\�C�ٲ���!Ɛ�ЦFn�<1�,ylqr�� �L ��am�<� i��˜q@>i:��b�zm�c"O�T�$E��+A��٤�Խ5��U�q��o�OtN�4�K�@tt #p]�z iQ
�'�4�8jӟ{���*¢��
�'��١ ���,&n�D�%�r`+
�'"��d��pJ��f��,"u�a)
�'Mu�U'�2c��q���!���
�'l�x�G�8R�D�J�*��+[ X�	�'�v������H;�Ș�Nm�����'���F��8��q��j�`��'y�ʳ���h9��  ə5[�X�	�'�1s!!�X@ &�%\i �)	�'�ش�Rԉ,�f��*ԴE��{�'�Q��bWijȼ��-�::3mY�'f�P% ȸ@�͸�L�;'��9�r "$�hAd��0&4�r�f�i��R �=LO���>���3P�8ԓ��.q�~� f�Gu�<�_�(q��F^�\zlp�K�X��C䉰^B�B�&$p)�!�+F�BC��,�1�Ҡ���B|W���'�a}BJ�p���&B*n2�K����$0�S�)�>W.�/,Z [b̝==9(�C2��u�<1�
�c��٣ H�"#�<0��OG���0=Q�+E.� �r%$\7���C�<I,��z/$�kp��0IWd`GbJ�<�aaM��ҴA�kQ)p���#X��hG{��)�1H�]9�舛`x����ۺ@��C� W�u���]�@
�Ҵ�X ����0?([���Rp�Һ�PTS� �e���(���$�)�@��ڸ��|5L�!�d��)M���S	4�����@�G�!򄌞 ��A��4L�^pyd`_�7h!�V��.5��L�	��)����:��$�D��h��9x!g~��slD��""Oj�#�%�'Y�=:rh�6��x��"O�����.�I�(�9v`�u"Ol��F�NJ
eBE<8n>��"Ox4x�$֢t_t��S��3��kB�'�˓��ɓC������!M����%w�7--�S��MK���!H,D�t��7�4�	�V�	L���OB��"�h�]A(`��x[@��
�'�z�#���#|�`�Cb�C��,�	�'�PYB�,n�Թ��� J���J�'��ۅ'L�A��P�b�8F ��{r�0�S�x7�9�0��_^�t`S�<chC�I�?�5���E�}�F�Qj��d�<�˓TvY�*Ɖ$9x���)$����zv��Q�k_��2�R�"���Lp�ȓ-�r8���2,=�q�?>Pd���`���c��?��� ͳ����jwf���)E�% 6gG�ö`�ȓz�%�@�wjH��Z�h5�!D����׮���%ih��r+D��X-I&��ؑ�$K�R�H6(4D��I�ȧw�(]R��/OX ���1D�(��$O%<j�Jv�i��)Q�0D�4 ��Zr��B&��l��c�2D��i�nE,^HZ�Ϙ�/wPLHf�5D�X@�
 �z��B�q�� �M'D��@Sf�e��`�1.Ѳ2��Ţ`�%D�L�F �fA0���0	���l)D���w��
0�zͱ1n�$w�q�o4D�d��V�;�dɹ7�˟-_����/D� +&�ż7԰��$I�G�����8D�� J�J�Z�A���eHa��mї"O�Q�E+�b y����*J �0"O�9�s*��x+~hg��+
��"O�e(���/��d)q�"=�԰a"O�r�ŏ�`^��C��ܸB�X��"O�d{v�s��A&��A���F�^�<��eкlB���F�/F!iA�p�<��@J'd�t�%�N�7֞49$�i�<��K� ,'�P��G$ZUh���l�<��E�#
��I��%��9����B�< +�!"���A&ٟ|?�E�Ǭ�x�<	t
�2Ia�h+��Ȟb�R��Vx�<d�vBj��a 1�ܩ� x�<��*̘Pv�2��S��a@�
�q�<	&eʍe�^\�f%H�[ @yx1O@l�<�W��?\-!��E����!�R�<�d�?�j�d��k~8pPG�TR�<�X��b�1�tH2$ï
�rB������:bE�e	s�]�;�hB��<�,�!Q!5!����㚠K�C����!��� yb&s�"չyZ�C��;8���xL�$e�@ꗈu��B��;X�� ��0=�u�B��Bx�B�I�L����ץ�����J}�B�I�Z���ALM+ ��+�@����B�ɔc�6Ye���D4X88�� e��C�I��XŻ&lo%�)"F"_�VjC�	�,2�k6�ֆ�z���,؝f�6C䉠(BV��	S��R�`�gֈ	�ZB�I�Xd�C��,uBm���T�@B䉸(�̐B��)�2�Qů�1\�VC�	���3��5pa
�r�C�5q�=�S#�$3���T�*�C��7@%��y/֐>���9p��iTC�	�RzB�Rg��,C��U��e�lB�>S�~�# �[?1�V�*�mݼy�B�I-'�Ԁ;���+y�� h�k3�B�	�Ck��C�k�-+���%p�B�ɫ �AҰUf���ۑn=*�C��>pn�@u늺3 �9̗I �B�ɫ,b����GG���͋1j�76vxB�I2��5�hZ	J���@�D�mhC�I,F��50�둤W��¯��9X�B�ɨ!�J4�2��?ו���oDmr
�'_�a;���:n�`2	l�"l:	�'�@�w��4���шP3a3��r�'E A	BOH�>��3�%C����ʓO�0($�=~�l�� �B4ن�(�m�2�U�6h<�!�'�	}`�t��{�uP�dD�]�j�T�\k�����>4�1iH�NZ��Q�a[9b1\�ȓf ��c�c��5%3I���'0D�(
���/�u�Gf�9��D`��9D����ȍy���%={���$�,D�@���
&1�[� �~��9�!I(D�����Ae<<:���=H{��j$D9D�X��"U0��1��2jl\���5D�� �J/�T�B�U�@>��è3D��X ʄ�K ��:����?OErj3D�P�wMV� �p1�!�X$��L��C1D��E/ׄ3 LK�m
*#���93D$D�tx2O�L�f�b���{�L��6�-D�,Y���Q�����"O�
.f��7?D����,"�M)�I2�nٳ֍=D�� X��A�G�1��IAB�i�����|��D0��'��"����qj��:�<i����y��5i/�0TB�l쉊�nŕ�y"�˓F�6�+"�Թ*�x�#	�Px��iz�h��%>e�1Y�@0~V^���'��`@w�B'\��0��CPn��q	�'�0�Yʆ�-�L�m��k�B|�O>I	�5��ؘ��՝Y���6k�O::ه�M���;+*����a%X���Au�'k�x��<-¬�vF_6k�@Y	� ��HO�OeS�O�}��w�x�ȱg�t�\9Ȉ�SM��j���GgK65�H� ɕ�z{�5�<I#�"����O���㔀G�V̩%Ģ@t�e�'����+�J���I�:����G�i���<1�S���"��`�����IpZ�iO��E{����B�0��M3��W71Rb���̯�yRH�*��4���0�������'�(#=�'�yB�C_���a3�	?(H��	%�Px�iS�<�עT�>$is�9xD2,г����Y��~ң)����/c:BP� eF�sF*�	r�I;feJ���c�4�S�9_U�h��=<(��mZ�Q��6�S�O��<���(�b�h@�κrz���'L��т$���* !�;�p���'+����ʀU���`�X-Ғ\*�q+�7�T;`�1�-�U4I�q�5G�!��A9�x�&�(��Ѳã,�Q��D{���� e�ڮƄ(�"ťR�
1:��5D��z�d@�.4z��4Q���p�2}��)�SK�����	 ���m֮o��B�L����fQ�e�����D0�$/LO��Pk��
����d+ʹ(t���f"ON�(��ˁwL:H�� Q/E2]zp"O֝���T߼8�o["Tc��1t�>��+ҧ<<|���ͤ>��)ЀM�mzx�ȓ+���0�	T,轛�!`��ȓY�,0���#0ˬ�b* p>(���M�w��v.ECA�n\x1�GA��ē�hOq�Xa㒧�L�������O3bѫ��'$qO<���ةA@R��R�\�;��z�"Oq���̅���v,NF7*���s�'7���9ot�����r���L���B��#E�@U�$ ���\��'�ց=�0�':ў�?����x�����k�
4[Sj=}R�)�>����M���U[�^��ؒO2U[����ކ=��Ȁ�o�_Kl=" ��=G^�<Q��>I"�� ��A�/@Ў��$�Q(<)ݴ �&@IC(�<j�8�$�2~xy����	��MK����u��i"R٣�޾,�L���hR�M؀3#�;$�ܙ򯒝~�6��+�X�<�xSD*D�x��k� p�B\9�<sX�ã=Of��ēu؞�ۄ���m�D��H@�.���>������"[
l��l;G��҆�	��yO��>�R���Һ4�P�Q�(���yR��",� S"�ޡ2x� Ý2�?i��$�8��'�k�� 84Tyl�2�V��%?5�!�DA�H�mAVH�3.��y�&�-t!�Ĉ H�LD1�([�@K�u�%����z��'��_=��3�A�������\�0�Z�"Ol�c
��e�&�e��"+�Ⱥ�"O.�(B�~� ��1"4PQ"O�A�G6�N�j�.H'B���S�'�Q�,�'ʱ��]XB�Y�K�6|0fM̂Y�R"O�P�K�;�Vt"� �xA�Ѐ�x��'��*G�&�쐒E�O�Ү��
���y
� ��x�ʛ��1� ��nDA�S��ϓRў��*`e�˥K�8h�@�@S��u���	���'?b�pt`��g��Y�Z
/��h*#"=D�!�d(�@	{7LVھ���
H�m��|r�Ov�I�"�\yȁ�����A[�K 9�n�T�'L�l:��±_�B���6:N��/4ړ�0|J�"ƞc�`��pU5 �0�Wfa�<A�e�Fb��A��U�x9��q n�Y�<���c)RD�fN5~��H�6�NT�<9G!S�hڰ	�.U���0�aGS�<�1BȽ\��3�Hǂ<�JYzV�Y�<�k� ���DIA�L����X�<�!nLd�Ɠ'	����V��M�<�1�J[����𦉣vuBt�Ȑa�<�cגk�EJc(S0doUZ�<��ɼ <�"'H4u� ��o�<�3�3�0�����B�R���'h�<	ϗA���I"`ULw��#�k_�<!�h�:`�ļ�2�:9���^r�!�D�!9�Pb��PK~<:�ńm!�$�$x}�g#6[,F͚CŜM`!��Xa/Z�w�ݖBD�Q��D��<b�y��O��Io](|B�/��FMd,�ȋI�C��z(�]c�f��a�8����?��C�	�4�+#�2֐*@���&
�؏�d<��]8u�
R����'��}���"O������ U��-d��q�҅Aw!����P��e�A	}� ��! �Y!�$����ٰ�c�� o�>z�!��S�*wf�Z'q���)pD�@ϓ�O��"�Qr�nX�� �j��xH<ɒ�ǉi��E�u��0یô*�ty��=�h�s�gJ�f� `�7�Ӥ+zC�	#<���u�?D��Jb��fC�^H�`��7a� 5����B�I怸�q@�17RX��V5P �B䉑N���/�?c�DM�2.�NC�I�o� 0��-g���*E(U-��C䉹;�b�7��.j�Hd,R1戣>��'�>M�wV�- J�P�cW*+pRAs��7D��K6���)��0��5���z���OlL��JBx�93���aOT��^��* �3�>�l���/伲!��<Z%�B���I[���Mk��d>�	�7k��2�o:8 
�O���E{b�xaD/A�@���r@B6�U9�y� �6i�8�f�F8~�AS�����<I�'k��ҟlH��(6$�|9$IʀEuٛ6�-D�����]et�8��II):�Pw�?T�l���ŜV;��Ť�+��`S�"O���C��4��I�U��A��	M8� �Ç�;y}9x�Ӱq���1sE9D� +O]�T�E$8Li���2 �<�󓁅AiF���#$3����@Ui�<	3�D�+l�Q� ��l#��r���K�<��&�#_o
9����KX��f��E�<�f�L�bP��1P�v��I_�1��x�?y���~*��ڊz!� ��.h:	�v�u�<I�B�1Ui�5�U+�Ԗ%�"i����IL�S�O����/f8��e�{c��""O0gɳ{���KE�Ur�/�y�	�%u�]R���p�"�ɇ�S�y��0zT��(�1k���'���y���fƈB���f�|y�W ��yM��U�$-1��[�sVZ�� ��y
�  b���| ��!�M/���j�"O��FV�7���8��M<'H��"O0Y��3�t�@�Ա?&��"O�MI��
%����n��,�(��"O� Si�#��EBt�R�+6"O�@���b��xx��C
�F�� "OBa(�osXd`t��*�HJ7�0D�(��F/�dU�0��{�z��6e0D������~��܉�h��:R,�Ԭ;D������<�JZ�t�2��s)Ot�<�.;F��)����y�%���Gn�<��Jj9\��4a[G�������D�<�5�L�B�d��A��]���谂�f�<Y�ቦH�4	U"��e�<th ��k�<�  M$�ub"��\��@��B�<������A��L�L�S6,|�<�t+ғI@@�����k����t�y�<ٱ�OGM��kؙW(����s�<�5� �?�*5h�c��s6Vqa�/Ro�<97�P�fXz #;&怀� g�<��MC6e�X�D ǔv͔�@�`�<a�'>ڦ%� ��w�ܽ��,�g�<�G])}v���T17,��e��`�<م��E���0��F	B�| G�^�<i�#آ9�P
Die�4C� \�<��(&+<a�#����}B��V�<  ��:���e�8jIZ���Y�<��@ϴA�x��T���7F�,rBq�<yt�Č�c�H���9�X�<	fn<�2�K2̞=�2d�C�W�<�等�#w�E�AX'P��`fȑH�<���\�)@�����kՐX���G�<���Z\� �@�tԾ�Z&*�j�<)cc͇`��tX�e��{�����.D)59�@p6Ύ��>a�/9� iJ�e�
�d�H�<� �C�Щ)��=��d
���H�<��.�q���e�5R��9�I�B�<���C��|�@�^�BU	fFOk�<ɱ��>^�����a	F��qV"X�<�#]|����AC�YTp��T�<��	��]7��� �����y����P�<A�/̔���� 
�QWR�<A1�Ÿ�r� �'JEd��'DF!�y�
��j�@}���C��w����y"	=`O4EX�֎(���	�y���=p��g���"Pa7C��y�Í�F�&ܹ��8xZD�;�yዀp 4t���Qr����p!@-�y��7_l�pR��M&h*�-�f�yrK�w�|{�e>�컆���yb��(T=��I��?_(h.*�yª�8U.]�sF�:��� n��y���?{^iiv�h�� ��y�Մ/M���ǔ� ;Ȁ�M�;�y"&N%F�ޅ���2SR�M�'�#����d����H�tr7��w��$a�.����s�+UP��'JׇO��P�D~����	������A	N%y�'��v$��'v� RP
�+=0��дQXzt��E�����#�L9�]w��U�' W�d	�蚭Xt�����>y֝b�͗�e�T!�h�I������G*�p�h�U� ��<�$_n�t���m�
d�V�I�2H�����O�Ab��IL��˔ !ς9��5Io܄RQ�@�W�j�4�0F��H���M�I0�hB%F0~�s���yO�L�T��$Qn�A!>��M���d�'���2�#9�P��oV�4`B ��+��)��	��^�vxCFD 朁B�!=�@�����0hR,`��/�j����%qLVIs���%#����KF�:��'GHi�L�'E�e�sA[�}�)Y� �I�ʼ�d۶8��\C���dh͛nO�M���x�)At L�؜�V��6��8tN�?�aN�C�d�T�ƫ�;wM�<�cO�C�d�T�ƫ�;wM�<�cO�C�d�W����2}F��݁��i��"X�SGG����߁��`��/Z�QNO����׈��n��!U�]IM����׈��=o$��hA�(DLPB?�%���=o$��hA�(DLPB?�$���:g.��eL�"LKUA=� ���6b܃!��k��-$*��P�Ҋ+��c��#-$�u�S�Ӊ+��c�� )!�r�W�ш+�n��jt�,"$3E? 9�]2n��l|�&)(<H3>�^0m��`x�#/(;B74�P>c����ZM#I�R*���a��ד�#��[M#I�P(���e��ߛ�+��]N!I�P(���e��ߛ�+��]�_��g�t����_B�������Z��d�p��YB�������R��j�z��QL������Z���'�Gn���f܉��Yʹ���-�Mg���bވ��Yʹ���-�Mg���bވ��[ɼ���"�A����8�z��w�蝧[������1�p��u�ꐮS����:�r��t�랭U�����Uk"R1�T�����޵Wi#S1�T�����ݰPc(^;�S���۲_c)T�{����!��ȶ��������Y�w����"��̰�����[�q����+��ǹ����ɂ��^�s��N=ӱ	٘+О�`k�%	�h��O>ַВ ܕ�ic�#�j��M9նѐ#ؙ�el�/�e��B6�s�X6���m�$�g��yf�r�T9���e�-�n��wk�x�S<���g�(�k��ti�x�S/3P�y�fF$PпfLp&,3Q�y�gI*]ܰ kL}($ <^�w�nE"QвdGz. 9�z$��aj84�O�_�O7���t+��im=7�L�Z�H0����w)�im=7�L�Y�N8���|#w@As�m���Z���K��#�yOO|�`���W���Dq��!�tDHz�`���P���F|��$�zN@~�L-w}es���_����K+s~gs���_���	�F&~um{���_��� ��N��^Q��!����^�����N�\R�� ����_�����K��QQ�� ����Q�����I��/E��C��b���'^�<�ܾ-F��K��m��� [�>�ܾ/E��B��e���-W�6�׵%Lژ3��~���U�g�>�$�>��v���	σ^�j�>�)�8��u��� ňR�`�6�,�9�����s��>k�m�X�� ���s��;l�d�S��s ���y��<k�b�R��}���vP*CD����M�U��ϚmJ\%CF����O�R��ė`GV-DC����O�R����hM	["IO�������"��-���Q"�������*��(���Q  �������'��(
���Z,�����Bf��61m�������Ol��32o��������E a��88g�������L7g�j��۔������y�T:e�o��Ԛ������|�\2k�o��ܑ������|�]0o���\J�:�o���J �	�]��Y
B�0�c���L��]��\H�?�g���G��X��Z�o\�3k��i�z�8)��ڥV?�dW�;b��i�w�4-��ۥW<�fU�8g��`�|�?!��ҭQ9�gU��Q(t����;�6��(��P(t����>��5��#��Y.q����6��1��'��X"~�f�Z�;�k���9LN-J!�h�Y�>�i��	�2AC&@(�o�]�?�i��	�2C@ G �g�U�/���rV�ߒ��<J~~�#�u��wS�ٚ��4Bv{�!�t��yZ�֚��:L|q	�%�siED��Q�[ٛ[��u����U�dIN��W�Xۛ[��u����T�gMK��P�^ޟX��u����U�fKM�z�޶�N��p�E��~P�24s�ݴ�A��}�N��~]�<;}�޴�K��}�K��t[�?9~�֣�����{�<p�%z\�h������~�9t�'{\�h������~�:w�"|Y�o���^kփ]�5X��ԶO@*��eSb؎T�7X��հKG!��lTgیQ�?Q��
޺BO'��mTgی���x�õZ덽�W�c«���z�Ʋ^�Q�dƮ���r�ȼU僵�]�fģ�/�'�1m)
��$dQ�
n�'�/�4n
+��,m[�f�"�-�4n
+��,mZ� b�'�(E����y�7~@3��{x�|��G󹘱q�=uN;��v{���F񼕾s�;uH9��ys�w��H���82�T "0u0��?���v*�
38�R!1u0��?���v*�0<�U&7p4��>���w(�40Ｅ�	D�S'��C�-�3E�Ӄ���K�R%��C�*�6I�ދ���D�Z/��C�'�=L�ډ��� L���wy.+4�
�gW�n������t})#<��`Q�l������qq$ 8� �oQ�i������{~7�.uzK��HC���U���p<�#utE��AI���Z���t?�&r|O��ND���]���t?�&�2�a^}*�F�7S�M!8�#�0�f]p'�B�0R�M!8�!�9�nQr%�H�;\�F$>�# �52*9Dn׵gO.��>�44ٽ2)?GlַdH&��3�9?ӵ5,<GlַdH&��0�?7ڿ> 7���c��k����ޱ��������l��d����ܵ��������g��k����ս��������h�⾠�c�醡{A_�ɭ���跨�f�膡{A_�ɭ���ལ�k�㌫qKU�����
�⼥sK0K4���J�|?I�����tO3F9���C�u5@�����}C<I6���M�|>D�����~F;A���m�wx�/¥|�H�ۜ���h�{u�#ȩp�D�ћ���e�|t�&ʭu�C�Ж���e���H���w2)�����G���: 	�����B���r7,�����f��j|���L�~��'g��i��my�����M�~��'a��k��av�����K�x��*m��a�l�'���oM�d���b#�'�϶�&���oO�a���i.�*�ž�#���oO�a���k-�-�ϲ�,����F��\�+7J��ʱ([�6���G��W�+9H��˳*Z�4���B��S�%:C��ƽ$S�4���|��Eb���9H4����T�w��Md���9H4����W�p��Fi���	3B>���^�z��@���ג�o�F-� &��u���ӕ�h�A/�*��y���ӕ�h�C!�/�
�x���͙�m����y�~1c�{�Μ�g����p�y6d�~x�Ǖ�a����t�r:o�qv�ˑ|>��\�>��-����_{v5��U�0��.����[~u4��W�6��&����Y~u4��={�o��M�؛&�D��	*D:}�j��E�Ҟ$�D�� H7q�f��J�֙%�G�� N0v�d80eoE8�/@�/<��w9Z1:cjF:�/A�*:��q<^28bjF:�/A�*:��w;V:0jb4Q}@�'o��I��*(i�30RA�)n��E��)*h�10TzE�-c��F��##a�:9\pptl��q�dhM�#z1!��Yuqh��p�dhM�#z1!��[vum��w�mbG�*r6$��P{b�n��k�8*^�"ueӔT�L�n��k�?.[�/yaҒQ�H�k��c�1 U�'reՓS�K�i���[�۬��l�Fu����L�[�ٯ��i�@����D�]�Ӥ��k�A}����I�X�y4`7�#��^�:g����v=x4`7�(��T��4o����u<~3d2�+��U��6l����p8}1e28L����g~ LH`*`��3F����a{%IIa(m��
<O����d!JKm'g��2F���7���Y,G�Q��`M�F��4���^)B�P��dH�A�� 1���_)B�P��eJ�E��9 8��E)� #���S�|j��TbB9]��U@���/�0���ǆN,6��uɘ�u�+�H(�űAf�
�x}�H�zH|�(�,S�Xr��>R�t1�!��B�$��'��R��<���,K0�� ߩE��3�a�)) �D;�皝@v�Iɣ�=6��� N����c��>,q�(��"�PR����N7>����K y$<@���0-~qɥ�R�h����$������i�1O>�� n������W\�,���ƈ��	�&g�����(<6�H���?QZ�D�oދ+���#s��aB�����d����rh�>0�\�Q�A>US�hzV/_09ꈑ: J��A�N�R�2jr�,�#nX���50d�U.@�$󆧬|���U��ې���$��.532��o�
n_/bm@���ۘl%��n�5+�V�
�ŭq�������{�B�4+d1ȓ�L�S�#D-�xn$҂`��2��5�e�8F܂�&�033�5V��#���ym29�R��04��P�Ş�E�DZR(��mƎ-f��b���<N���eBj��	�jxJ�!2Č+Np�V���Bà?��6��251���%!]oV�9�R(��!������ܐ�<@�!T 
�"a.�ߵI�L�M���qR�-E��-�� �O����N�"p�
d��*��A��I�kB��$��;[�8�O��0Ynha�U�yCx�lZak�q� F-'܌*�/	�r�<Q&��i����T�r0�7ٞ6+���U�E>_j�{J�3�M���ś������
����Od�9aO��_�V�ځ,�W2��SG�M)4��3$���l5q5�ؼr�μ��Û�:F,�r`����f/"���%]��r�*F>
��Bc�-xN����(݌��!�A//6O��� ^^h"��ϋ'~�� ��Z0{=$p�J=Y9
��f�ƈK���A�7d�����A�i�j��'�V�׻��mS$��$tz�'����	�8�� C�E7m� '��Q��I�m��!A&� ^2m�◟g��-����d�Z܆�x�ωX�HˆK՜�y�-�5����5Hİn�P�)ç(�:��ؤV֘a�f̉�<��McP���w#�mR٦o(�s�[4*b>=�#[��;��^�/D���
�?E�-�ЏԱB��	+u�� ��@>P���K%Eh�ZO>�G-P5R^�,)j
�h���
3oh I�%͐w��H��+2����6aP�PY��<�!p�iQ���7u��� `��	��p��d|�t[G��p���ˁ���D��j>�aN���&l�<�~�Cg%	��������s|�0"5���tT��ҁቒQ8�!
���߃RGX��h�e��Y+�e��o�Q?y3t�����5B��bb�߱E�� k�o -��mK�w�])B"�/t(Ji�u�G�
,�j�`�S��8�"�����QLhy�!n[�#9����+�8,��IEDV��} �#�;�(��"���jq�a�xRC�X���8(ˎk`�YʈOnD����O^�)g���?ys)85�C0b��2�x��������3(�3 +ҤC�/��'�N���X�,���-Ea0��B���y�d�O��rD�S�*PI�nЛ%J�$���ڬFi"���bU���2$�0O\���P��64����A�m=��֋���xrC�j���^�uRL�fL
�N1����ʆ�L:�IK��oĢ,�����d���޶q[ `��K��yǉH�`�d�0��UG��T8S�����>)c@�O��`a�@r�6��L�.
O�)끯_V	y!��R�xʲ풠�0���85 �v�<����ۯH�'�*�g��+c^:4l,`��3�ĉ�uj�P�4N� �����4��M ��ô������&W�L��Wg��|b���!Fָ@�pX��U8|r��w��`f��d�:z0�#���HQ2���J[2�ۀ���4cP���l�ҐHP&�� �!J0MXю�'�$���ӻ~Z0���2�Lӡ΂0
��{�Å��0?���ѹ.�-����*L H�9�&�	�8���!N�ꍂ�E�rn>-�@�A �!���+N'D�qWf�����JE�r2�l��ԓ��C�m/��`���0��x��F5~TekEǊ&�^���\�8��3B��m� D��i~�LÕ�C><'�|��	÷Z��Ж��5_�*ă�"6i�6t�',�j��ι0��LҶI�v�䉋�Oʉ����	@��cGϜ<�\-���]�{o�d�9s���3��0�<�R���#4fRe�)�=#�z�S�B�ϲ(z�Դ;�P�+W���OzuHC�A�%o��3G,�H�С���6 A�&��q���o�$�AA �0��C�/J�F����� pJvW��:ƥ�W�x�� �a|R�ۉc��-�Ǆȓ8����$M��!��B�IXƟ8��
O��QbI��d��Q�Ҧ��ÉZ?5E:��,Ҳ	��<)�E?#�P�ʈ7$!40Zw�ɘߘ' 68JW��ئ��7� /IF-�6d��E��<���ʦ�b���z(�*�G���YI`�,A�6�G@�-rWx@s�*ؗ?j�"�S,|>�J�����u�'�UH�jA�r�P����d��B@)х5�qQǈ�	�p96!K,���j̓-�|�a6K��l �O*3��Jr��##.A���'r�b[r|�QiC��#>����2\�l�)ჭ�Rd��
^�8aR�u��q8��y�l�t(�B�h��\�⩱�0X�r�)঄-&b��b!T(]o�z���m�'����7�@	� b�`�*\d�a��M+*8��(ixh(��iP����)NU�3ぴI�6(۳�U�T1R��T4=5hӴ�18aLјu�ߔ�6=P��@�kT�\0w#�q~��ǀgи���9`�"����$�h4 �mʓ	�l��R�+������?X���hDOЉ�Asª�Y;L�n�@��蠎�5#����e���\���@����8!t��
�U��h�_�i�dE�%d�ʐ
�Q��@�g�Q@D���Q34�&�!�ßz��iW��?s6e��j��z$���GJ�5wJ����'҄?���g�?ғ�5V�4!�)�ä@�/ �!hr�ߦz�qcb��<F찲�^  ���'x�4�1��?ODՋ�OРh@�m� &��U��I�����|����(Mdt0G{���{�\�򎞆~;&�g���Z�H�� V��2�.��Fj����%��]�2��C���
|"�
ÓX���)­9?�������c�x�96j�:ݦ!X6! (hz|˓t�h�&����ݙ5�Y�Xw��� �7h
�I�����H-R�Nͳc��1A�̠���Q��&�z5=9���;*L��(s��*�n>�'6.�i���~�^q�'	�B@öc���̘�j��[u�@y�@@��ħ��8���0�ǐ
!|0B��R"d�6�z�ƛ�bdr��!p�"5Z�.�*��O�� &&Ɨ;�Ԑ��8%m URq�E�1��Y���̋)Mµ��=H83�k9?a7dL�N't�HF׳*��� B=�w��i9�F�$�d��E���@�YtD�#=E���ejU��=H H۞I��%�ȶU8|�zpBդ���Or�X�@�+K
u��=�'U���(d僭}�`�"��*?��'��ѐ5*�Pv��cj�4��\����ژO�eۡ�F0t, �5Ku�EJW �6�nSג>���>�2=@m(y��K�F��)R��4++<�CT��%�:	B�.� #pQ�|b�n1}2͗1A���U�H+0�HQ�R�\��y��ͱY������/b���JqU�dR�O�#m���P�J+"�)� ͧ�ڈ��[	�p<�g��'�`�jDk�|y�KzX�������
� ��׉v�f �k�
$kp��#A���a���u�tB≢T>4ABWM��R_V��R�1
bc���rƏ�|d%R�#Ӥu�����3H<|<4&BT+8�e����m�<Y6m+��0��_3k���Y�l�*e�¸� ���ӧ���$�1.
R��4C�)t��M��4�!���s��L O����k�FK0!�!��Q�;7Vڐ䋬����E~v!�]3,T�۰���"Px!)��|!�d�/d�0i4  :tb�e�/��,V!�d���Ƥ[�L%?Z
����Ƀg!��4G�(�(���oB,��.[6yU!�X�D��5`���1 �7��4�!�d $�DEjC�X;c!t�1��j�!�Z�L��� '�j�r��iѳ�!�]/)B�X��� �M�n�AGe�1�!�P#��y��l�:P��6�!���X!�%����9�3*!��$w
Ȩ���0 |N����Ԉk!�S� �݀u�ێ
h����#!�׎g��@+1oq
�dm��!�Qtpp�I�=~l:�#�A�!�$�F:�ՂH,Am i��#6H�!�Y5)��X�wc
 5Km�׭
1�!�$,����ɡe�6�{4)�u&!���bX�eߔvJ2ѸSI�B.!�dD0F2�m�b̀UC�7hѴ�!��K�mQqW�)L"$̋s	]3h!���"j_�:�Lh9W��Q��$P
�'�����*USF����C1čS�'��ٲ�F
b[�uxtb !:X���'#|�;�B˞ �l�ȴN_!
��	��'���! Ěvt� ��7a<da�'-j��
G6=���0�ʠUj.��
�'e�Dqp�G�Ե��@�qF �	�'����iC,�<�	`HE"a�\9��'��H3�.M�F�la؎	P{�1c�'B�}�c�.0�=��
ÜL����'�*�A1� �Mw�T wH�Gp��`
�'��|��E�&b�q	B���`����'+T���N�(EK�щ�NE�N�(�P�'�Z�0#F�Uj��RDb��',L�c��P�cK��Ѣ�	�|^�s�'�*5j��y�z�+Ɠ3/2�P��']���&�ħ~	�`�aC^��`ȃ�'�8M���)8��Qzw<i�'.&�CwD�QNxT� ��,~2j�	�'���fO
w�6!"�*ޜm�����'�d���Y $N��V�^YL�z�'�85[�*�
~rz�Bc.HP\���'\č�PKP� A�V]�4��'�
�*�eXh�8�U4_d����O��QB+��*^�i��O�~����֣ ��@�V��/8�
�Q����$D9�a�Cth<y�œ14HCJ@{b�X�a=�~R���S Ȕ�CD���1�ҩ؆�1%��	<2@ ��~�y	.�&Np����,6�@�YSF&�OԜ���92�"8�V��?L�	G�ƮQ�9ip킳i���ГA�s`�:�l��((�v���`�/���wEp�I�IX�+� q���7��2�.H/;�2�%Eބ!�� Ц�.!�����p`RҎq�Jg���̶���seTՉv�M`���ϴ���seTՉv�M`���ϴ�����>e��`�P�|�Qf��]����>d��d�W�t�Yn��Y����:c��h�X�{�U`��U����6m����y��A�����( 1�O�����y��A�����(!0�M�����y��A�����(!0�M�����ŞD�F@��rΜ��h5"V����E�BD������j8p,V��ϔM�LK��qΟ��b?u+^��ĜF���@�#~Xw,�t�����B�#~Xw,�t�����B�#~Xw/�rƢ� ���J���p�>���2�?VF�� ��H���{�7���0�6^M����B���u�>���<�1\L����B�183���6Ɠ���"f5/=�183���6Ɠ���"f4-9�60:����=̛��� e0(5�:5>����!�Wu����$��9����)�]z����(��:����)�\x ����/��>��� 6���4V�b�/��v�� 0���?Z�m�#��s��<���9Z�j�'��y��/��G(xh���4\�� (.ێ:-��F(xh���6^��&/&ӆ2%��B+zh���6^��&/&ӆ2%��B����i�{�U��LP/�͍ߑ����j��X��JP)�ǎߒ󧊓d�u�X��B^ �ăМ������sU���{��E���	~��T��y_���~��D���	~��T��y_���~��D��}�y��X��tS�m�F��4��n��r��W�m�O��=��l��z��Z� c�D��:��m��|��_�e����G�!���2{�U�B�ӑ���F�!���2{�U�B�Д���M�,���:|�Q�C	�֖���L%��|����:�j�}��?��\�(��}����:�h�|��;��S�*��{����3�c�u��6��[�/��{�}�L�1 ��*��^�G��S��|�I�9)��!��V�A��Q��~�J�9(��-��X�O��[��u�D�=���S���E�)*���?���[���L�&w$�͈7���Y���I�#s'�̈7���;�ū�q.���.��0m齆�:�Ĩ�q.���#��=o鿂�<�­� ���/��2f㵊�1��:�^�('�����<c��|/D�3�Q�"/�����8f��{(B�7�S�"/�����9e��s!H�;�Y�2}���$�a�٨2����6�=|���!�d
�ѣ<����7�6w���.�k�Ѧ>����3�<|��|RaX��t�Z��o
�NW�6�tZi_��w�Z��o
�NU�3�|PbR��|�]��m
�NW�4�wYjmY�܋V��a�1�ǲ���fY�މT��m�;�ʳǨ�m\�ӋW��o�:�Ž̡�i^s����d �@�B�(uܸ	s����h-�M�H�/pߺ	s����`%�H�H�"|Կq���\L#�������������]B+�������������[F(��������	�����[F��:����)"��A'�`���:���� +��D#�a�����9����&-��K-�o������О�o'F\���g1���0{�ɡߞ�j B_���b6�=v�«י�i"B_���b6�:~�Φؔ�objw�I�|cO[�v���hgd~�N�~`K_�y���bllp�L�y	fJ]�s���bbcfT�N��S 
k+R�/�M�k[�B��P
k+R�/�N�lS�I�� Z
n(P�/�M�kY�G�CB��"jj�B4x�
t؆��CG��*ed�@0|�
r݌��LI�� %mo�L=r�rݎ��IN�tw�e�s!e��$�n��ͳ�t�ut�c�z+n��.�f��β�t�tw�e�p$b��/�c��ǻ�q�ws�q�xΨ�x�24Aa� %�kr�sơ�x�?>Me�%�hu�qŤ�q�42Fi�-�mv�qA�f�����~�!�����"C�f�����x�-�����,H�`�����p�#�����!I�lɲ�&\G�OW=Dd�Nf#���!YE�LR5Oi�Cl*���#XE�LR5Ok�Gk"����C��Wp�(�+a���0��M��Pu�-�"j��8��@��]{�#�-e���2��J�/m�@s��b�w�Q�^�Q?F"a�Gu��`�w�Q�^�Q?G!e�@r��e�t�P�^�Q?F c�/��A�bN8����=��}��&��A�bC5����0��s��( ��B�gD5����9��v��+��;����+��c%��+�����;����/��f ��(�����;����.��f ��,�����3��3/�c�#Wb����̼��:!�n�#Un����ŵ��?"�h�*_e��������?"�v�;`z��߬��	QN�m���v�;`{��ګ��UK�j���q�2jp��ԥ��YG�h���}�6z ��X�<��O݅j��(���r/��_�?��K؂b��"���w+��_�?��K؂b��#���r.���Q[��cM^Qx�5uʝ0��VZ��kDT_v�8vΞ2��T_��iFRYt�7~Ö=
��XR�s�Z�Z3��(U �˾<z��x�S�_0��(U �˾<z��{�V�X7��,W!�˾=x���Z���r�{P�?~/��=CW~ɜ��}�zQ�>~.��1LZv����r�uY�<~,��4I^tÖ��z<hQA~��\��ۤ/��)�<jUGyȇT��ݠ,��+�=mYHt˃W��ݡ*��#�1e�u<���w9W�(��垩��~6���y7^�"��ꓭ��}4���q=S�/��햮��}4����C�D��8���&,"H\����A�F��5���'/"H\����H�H��7���)!)MZ����DQ�n��p%���D�=C���Q�h��r$��	�N�0N���V�k��r$��	�N�3K���]�`�9��|KE�p��ל���)��8��sDJ���ڝ���.���4��xHG�p��Ӗ���%���9��w�s���ox�Fǁ�M.�Etv�y���nx�Fǁ�M.�Gws�q���er�L͋�E(�Aqq�s�7761
WZ۴N{�����B�g035<TQѽGr����	�K�o9?:3[_߳O{����	�K�m::=;��>�b�{xs�q*�E��5C��;�j�vw~�{&�I��?D��6�k�wsy�y"�O��>I��63n�X���v�sW`H���O:d�W���~�{^oE���L:d�R���s�vReM���N:d��f��tc��@��5��4k���j��qf��M��5��5k���k��~i��M�
�5��7f�	��a������*/�i;[Ň0H�������+/�j>\͍;E�������+/�j>\͍9F�������3R�@5h~8M*��R�w�4R�C2d~6O+��S�u�7V�D7ip5D#��Z�u�4R�x�9��A�6U)��u��@�r�1��B�6U)��u��E�z�:��O�<_#��}���K��<H�q���6j�x�%1�	�zOH�p����1m�z�*3��wCG�����1n�t�)4��wBE�z�~@$�ϙQ�����'^���J~A'�ɑX���
��/Y��OyH.�\�����(S���@wH"�R~3���T�$࿥����y�Xu8���
Z�'伡����}�[t8���\�/촩�����[t8�k}Tj��6�!���{1ӳ ���l{Qo��>�)���{1ӱ���aw^c��1�,���{2Ѳ���fpYa;D4��T q���؉�5��2N2��V p���ݏ�2��1L3��V p���ݏ�1��9D;���"&���Lx���kI�^Ҩ��!$���Bu���hK�^ܪ��'!���	Lv���bB�W١��/+ve�!�1��NWф:r�/襕s`�"�3��NWф:r�/褗pd�$�4��F^ێ0{�*ﭜyj�+ަ'y���^�5Ś�U�RѦ'y���T�:ɞ�S�Vԣ.r����Z�3�R�U֡/p P,r�V�Na�yRq�=�-�&�'?d9�D�&�����Q�n�\4JdW�Ji�aj�	9� 5�v�"F=z��Vi�<I�R�b�I�i�0%
��O���$hԪ�0�6�!�t�����M�D�:) "l�":@,G�o�R��#�;H\i��ƍ���v�T�8z^Đ��;j�l��Zk�X��G�;JZm���ͅy���l�8{|%�c�\�ȭ;A�ŇU�\HR�+V�?%�5x*���^xH�H�%f�l9�B����ɊJ�r�B���>��dN O�lY��=.N4��aO�H��dj�i��ݻdR2?��D��:�ڵ�d��<�tl�=Ì�V' W �e�3e���S,�?e�@Q:A���0}�t�ݓ-����0wA��1&�_23�н����h$jD��(�6����ܹW����b�%>�B�1cL��ƵSg�AX�\��4��1k���SƘ:v�����$h������!��-��k��Y
 ��z��p� :��l�HҴ��o�Cj�k�L`�O��GAe�v�֥%�ݐl4l�����j�lm*�H�(�Bx�fO��BJI���W$'������6iB��`e9ov�������لd�/S>����95P���a�K���p�Q�M41dp�;LJ��2�M?�œ�%T�t��	pAe�75K
%Ӥ�Y�~WVqGm߁\P;c�0H2���WU����`�&��u���ӂ2��X����90<򥹶`U�w(h��Ix��d��iXu����5��T����63�� Tr"h��[�=(��`v���`%ʴ�Ѝ��R����S��b���O`��D���`$c��`�\�i*����+>�{��4V�.yY�%#s��9UU^][u�SSSzBw���BDS�S[N}%��QYj5:��T�h�@�I Q�9k�Eϗg��ɏU�
PAE��0W�\A6��U�Q?���)ܩX����&�2Pޞ�dJ��Y�ح���H��MKƊ�1$�J�J ��R�*1���P�g��1���,��3�f/gq�1��d	�_ 4�X��k��b�i3�8�w+�H�j�P>�		:H�p���`��Ո@�ֿ2ZtI�	6,/t�ѷΝ�h�S3aĕQ�KV����G�F�꽹ª>���޹q8>�� �9�2 '�L�&���C������c����!3�9S�R�l��T��t��\ZR��1pF$*��� S���5i	� � L�u���f3�IB�>Y��ɉF�j(�;.n�պ���@�	�06��p�d��M�&'Y6
t�'@=�0���h��Q�&�L�������"
��4�f�n>u@��bG^�.��Abg
z�D�1"+p���G�&r@�Ƞ�O�N���7I��M�e,�'c8��U�U �Q�ԫ�%\��m��;Z�J��|:�CP:�y�Ҭ �t\Hd��T�d1JV�ʜg�.�rVT}���(w�瓸(w�|"�x�
�'A.,4N�����gVޘ�'�=uH̒��U�{$`1jV�Mz��[�yB��ٺ��ءE��(��Hŉ8��8�e #,
�JĎ�J�R��koY�I;3H*%z"�.1E�MypHʀg�	8wɟ4�0�0̀�7鴜�@BH s���P� kFppA8�I�MUJl��AGFs)U<32���';�8 ���I���q�%,."}��C�#����
A��.�����)(�|{Η�-�a~��{L�(�K��yƺ�QfJ�����n��m�P"o�l��ېk鈴���ģ{ž����O�5�!�J�WX�i��a��v���c��>'<�MIt
J9i�>\I��'{J�[�C�d�p1�t&�G�B`�PAX�F�1Ij�DT  - ���$��R�Y)V����3N'e�I-d�ڥ�"�>�� �4B&��zf�\#B����ȰK+M��"I�;����.�&H��db���ҵ��O�a��J��i��PP��$i�ƕ�ToZ�:�R��f�M�2�|U�6-��L��I�3JT.k��@`c�V�l�н��?�EQ�$ME�R;}���y��'���A@��3�n}8�@^�6KF�T��17� ��R��c$�:@��<#�j@�tQh��4NL�#)*��$$Ȉ�أ�G�����g��OM�'�ó�ݦ=�v�	0g>�ԓ�B#�����l��Ӈ�I8>c���N���)�!���{G�����	-/���Q��ayrY�MZ���DP�b-����eGe��Ȕ��ON�C"I�jX|T��X�I]�����9g&������b���$�U<M��yb��'��DS6�caZ���ɱ1��}
������C��L� 4�	��X5A�"��0�	�a�Ҝ�AC�q��a��

��{�-;$"�Q�Y7B�2�8G����5�V�2$H40H2.�x�'��1Pn�6A��5a����s$�=���24��0�兾G��JO��C�f%3�mL�YZ�[d!��C�Th4HW�0��,B�D�A����!?"(P�c�T<X�Ĉ�J������XR}����'At���ަ%	Th�i"��'��E�LH�D�����4@,�q���>���F.�?]3�b��;���nFB�'C`躢f+|`�"�?@Z,��Ư)h����V�S��6'?nms%T�8�x��r+L!.�q{��@�xb	�8���@Cύk�@�Bd�� �0>Q6��#�D��M�:~�F�Pq��M]�����O&���E�t�$e_Gt�H��b�L������̳�(M��a�a&�%b��
��0L�o�~b��o��6S�ih��Y��аD
�}�ҍ_{���S�%�`�X���
A\�3����9$1;��F�f�,l� d���=I��2 �z� FlÅHH�SqY���P��-8\�K�/�0S`h,~6�l8��B����W�Y*6$�#�ƺ��y�=މ!�ǆ��]�U�BM`�e�c�H�jp�QOڷ^/>��6ߦ؉�DJ�'
n|H�)P��,9����ѱ���C�ň�.">1O� .
&4&Q��H��h�4	��ZJ��#m��a�@�Pm���uT:�hO�@���D�A8��盧9-v}H5��U�`����U�c���b&IS��I&D�����Ɣ5F��W���S��T"dj���bT�����R��� _�@�ɰ��H�ΐ9�`���$�+�ƽa���	�xM+��ى9"|����0c(�5 ��%1@'�d���QW"R�I"����\�p<HhZ�r):	�D��R��9q�g��a���y�K'��6�v!��E�-_T0!�,��33h�Qdq�r�#�иr��3����ʗ��D��!�&�W(&�ҕzG*R�z��C��nj����q�6��1gνV�z-Dz»��K���΀{��
�`�Z��W�.'�d�z����r��@@v
�^�$�t�,m�*8�R4�5dV�V��$�H�4m�Ty��狭��lP@K��hO �EM�Ppء��A&%��2@C N��@G#@�_�~�R	&��`
O=E�b�b4�P�	�`4��B�?��O�C�%��͆�/
(��g�� *�2��a�ay�ބ8��`��Ά"�>A�1CJ ��M�Ȋ%��3� @*��[�v����	;5x�dF��v#��0�/�{z���C�׈CaH:��
w������ɶb3{��['Nr��bP#Q�y��YK�Ð�aנA��'�-1	�g(?�i�Y` �'��q
�N���h�'3=�r��6��ѻ,�e�=�S'�i��yz��;��}	�c��,)h��BN[,n�.�ѣj�F4���B⇨(����Ojh�%D�RV�e��M[�0{x��%�Qq���UDU�-�y��� FAz؉��P;r��C���[�x)�aC]�D�y:���pj��8P
Ǐ3���O��1 T:l����!ҧq�� ��8c���ct�� s���'��ٷ�S;�pɑ.��.+7lP��O\�r�Nȣ� �תݺ�|�2����&�4�Q�>!E�>�7�"p�]bӂʃN�`�Ɍ9xK�	����'2%�$�$I �N��|�	 }2$Wd���"���B@� ��y�� 9*P8Ć�	���I�g#��T�4p���Slr��4�%x3�Pp����BJ0x�F?�p<ar��*&ڹ�v/���f�[NX��c����?"�m�6IdEH�e
&wP���#�& �� �Њ �\�B�I�_HB���F**w��h��ϥV�2b��`�O墤A�%"�U�a5�S�o IS�G�Che���@�B�M���z���{G�i8�+�
x���Tʈ+W����g�>E��'u���'d�!�@���=�:�	�'G&�����b$|XW��=`�l���'�V��B�T`N�!�F#n���	�'d�ʲa�2��1�g�V�f��y	�'VD�i�'�H�P�� Siz�	�'��"f�ưYC��p��V�C�'�k�E�qǮh ��	C��hP�'f� 05��S�\x�D҅GI�r�'�)r��Q"����ߧK�\p�
�'$ ����Z�����4��8�'[�9[0��VS��a�(�
�2�{�'��y�j�*`�kGOI�X����'����~���w�!Q\H[�'�fI!�C\!>�I�v���r����'ݘ���05�p;��b�"ڤ�y�D�G�\s&7ZG�k!G	��y͓�>$ )H���J�ǈ��M��C�6�F���N�)-*��T�^-pD�C�I�d:���,�3A0��6 �1KvC�	!JY�P�B��'W�+a�P�L�xC�	�B_J���i�Ĉ��k�$)�XC��	d>~m����|�jHr�ƽh�<C�ɝNPk�Cͮ� ��1�%��C�u��YS�k��{yU�����jC�	�(�4�M0=���@b�HC��pՊA���z����U&,��x�M�7�b�E}"�
�^�i��^wۖ=H�K�t�L���ܣT�\x���t�ֹHO����+o>h�!�/�L#V��g�Pl��jV ��;9���⁕l>���!�1Xf��e��,N(���<�1�ם@K�l0��#}��	7P h��h�2w0$��O�����yb'b��?M"�L�G�Y��Z��S��^�M#�dC��}��y�B���ģq��8��ag&_"|�"p81I|ܓ�0|&S/������p��fE��~f���O��x��ʎ����	�4qTN])kz[�(h*�;i�	,i�8[��U( ��S�ONH�nxLH�B_�I��y��4��I���)�M}����L�/#4aⲈ��U�<i�,O��Dz���ҋ=|���d�|�V�A�3Y��GY����>Dy����`���+	5����T��0|�ԫ"w�hӣc�z 6<�dBx�'~�"=�O%j,ҢG� v�hI��L�p��+F���-{��ue����g�	7E�X�É7Aa�I�7/[X��xCd�-1��b?ac���?�c\%X>�qC�I�9�P���l�<��c_����h�(*�䝶[4��4���\Q\�:b�� bO�m�>)	çj}@���M�CƠq��O�$3.��{��@����Y�x�\��[��� 9��R�'���72�Ib��e�)§ �he�!��-��B��%Ֆ�ΓX؊ ����S�O)Bq�`�F���� �|��x�T�h@S�(��|5��WB� fB�H�j!�v&~�v���<%?� �)ґ���P\p6Z����:"ߢ�X���e�0�����m�\���ڴ(��]�3�9p��ȓ&�H���W�܍��-��yb��0�
�QE�De��<��Sc�e�ȓ]�� �(8�^M�$D��%�,Ԅ�O��d%� G��Dc�ߢi���ȓ��i���ʣy���T
�c>~��ȓ@��A�@l��Ҵ=�X�ȓ>�Ա�T?o�����Av�Lm�ȓO�\��Ԑf�N�I0ㄜ6��J��pϘ'�k�����ȓf~���N�t~���W�!�P��ȓ%�tIS5#�XlZTÌh�ȓIVXx*�nYI���` �E�fԇȓ�@�Q£:����G��l��K��� 5��%-b��IU�|bVQ�ȓ&%�H87�ز�4��6�ؠB�Y��/�]X��T�P*r�k���:��фȓ.m�<0 ����5x@'Z����U�,�7�W�`��`+B�tW5�ȓ��I0WE#�.�#��NQ�l�ȓF6nA�#��
��h��`G8hA�ȓ+ܐ`��C	4�Z���ԑSʈ%��2��	�PlT�q^��*��/���ȓ4�,1��=`�(8� cJ2E6 ��St���޳$.b8����~��ȓ]�I��-M�O� ����ӿ��H�ȓw���kq�I�^��4��)Y2:&"X��N5 �"ŗ�Bb�uz%g�36�ȓ:/��iǪ��M8.���7=w�\�ȓJ����B��,��`�G�0;�����(t��gV�S�H	�AIĔ�$݆ȓ$�`��ch�5K��R�)����ȓ}$v���F�
���'��k��a�ȓ[g�hpc/JU\�
�E|j,4���@�f[�I �(�J�:��d�ȓj:H���!�R�����nӾ8�ȓR;¡:��>�,k`o_�>�ȓVҔA��@�~�����t����ȓ&Q�|��Œ�J��F�Q]�=�ȓP9l1$�Zx�����V�$���&���Z��\�qц�Bp�2-��>4nĹ�m�[���Q1��X�����w
PZ�J� #B�=�܅ȓ/�<Rw�O�h��P�{¤�ȓ"��a��C�V���� \�����WPbT:�������1��V�ȓb�5�Enž=g5�pJ�07bꌅȓp[40�G)&>�d9�����]��4S�����  D
�r��ԲJa��� ��Q�D�nXi�Eh�nj-�ȓ;���
�d�=A�`�:����E�ֹ��+W�E[���V�ȉ$@G!9��ɄȓA0��*gҪR�0i�dP�B��}2�ȳ���D:āU%N �\��p[��"p�_�$�:�9��:V���ȓv|$���ث�|l��^=V_���ȓ,v�P���Ue)��^9w��A��W���*׼D�y�cn@b����ȓ,f�I��߲0*�ӣ��1N� ���	G��q��4H�d+Q�۩o��8�ȓy����ї�� ����#K�>���A�v� �a٦����۟R�ͅ�\|��6UD��iB�@�<�����S�? �8��ȵ����椘�vQx�"O����H�t�VH����5�w"O"Q���8<@�� �Ud���"O�Uy�C�&�:�s�d ���P)�"O�AQ���6�VE�vj�.D��$��"O�-p��ݓem6I�.����%"O�}�s�ΰT���ʊJ�&���"OtE�q�F50	0đ�lA%�XL�"O��0�iQk�ȜZB��|� 0b�"Oj�&�~�\P��'ߟ0�ޔ�"ORm�C�޶X{֐ZVD\��>��"O���V7w��S��6�Dy	�'3�����8 M�@���}I���	�'�rD0�mJ
9���c�� r��A�'`�������!��9v�� ��'�R8I���?�ʙ��;qL���'��""S'6 q#��y7�3�'��4zS���Bt\ �Q G7i�.	2�'¼0��@�q1"�@ѫ��`�����'�.���[�\Y� ��� T�8lh�'oT�j��3~���_�t�:̠	�'��laf�����s-�4o>�l	�'�`"C,B���z�@yG�Dj�'���q�Vm{�HKF˹H~�b�'^~! �T/��D�V���B�C�'�5�$ Y��l�9C�� �.���'dA��+W]`i���@�s����'�|M)����;b1�b�F4[�Z��	�'���tJ�5d�;��+[.�`Q	�'N��A0F��z1���a�X�N���	�'X�	pU� =���I��K?>����	�'�x���SE���̚-)�`	�'#J]��ڵZ׊����7u�U��'��t���⬈bo�Zj�!�
�'':�s%T
Y�� roO 8 9�'��yW"�+@�9�c�`�$}�
�'�R�B���t_ވZ�#�8���'�:�hUMн'����� �4�I	�'s��څ��h�tl�0��gIs�'bF(�H���ɉ�ǘ�yk%y�'�
j3gN�lO�A���udY8�'��!Ys�ΨOTP��)V6l��*�'�J�[�F8�fu9��U�/ԡ��'C�MQ'��.I E�s��QI�'@���K�&�����M��q�b�
�'�Ib5�߃tt��@�e�i�-�
�'�"�C��(+ۀ��&�ڥa߰i�	�'��m��.�k�@|�Dˇ�TGv���'�bIÀ�V<!	�LM�K�j�2�'����D�R L=�VN]	p�D����QQ+՚X?.�!�K��8)��\���p/��b�(P���A�Z����Y�٘d���kМ*��d��;81��({Yh<����H`��
Y�])���U�&i�& ��5%�H�ȓvr>���m"�p�nϭ ��ȓn�Z�����2l>�4h���B�< ��B�Yhp��A��qV	�r�D�ȓ7�Y� .I6�5���64���ȓ1�����E����W�4�~���I"�� UMM�f�v�VF�x~I�ȓ]tX�s`��2C�Ր�Ģ�.y��:��ģ��U*Q��8Q�[3p��	��F�D�3L�Aߠ H��B�7� ��S�? �L(Ջ(���r���((=@�0"O1������yQ�D> ��0�"O�t�ңVr�r��5��i���""O���#)�M\�q"u)F�~�:E�*O��C�g�y1�T#�ُ`�@�
�'�>�2�G!u�������=�[�'l��4�� Q0�,@R�<M��i�'*��)��(X&����@>�y�IA�	�����h���=�yB# ���HU� /�p7aX�y�K[5(�|�QA�?:�Dq6.��y�H�IpfЖ�V����F�$�y��H�'�&���D˚/�.�C��H��yrD��pVj�����	c�̠	�'��ؒW�T eѮa�s� 5	��m�	�'�Fl�B��0h�2г� �R����	�'����K��t,1�`��53�����'m�u������q'#��#����'���8q�OG&�@�� �L��'���2Ą�-:~�a@�̺"g�1�'��x�g�ŗ�8�[�B��+����'H���CD�n�tc޼+<ZP�v"O��YVk�-@�� �V o-��"OJU�&LK�
�|1R�C�r~d=��"OZI:d��	Q�T�[�)�a_�ȉ"O�4�T��9 k$)Q��]�f�,%9"Od��`�Bäእ�G�`�"OlQad�Ôbf��d�	`�x�p"O�<�i�N
T|�ea���1"O�4�gC��G5&���-P��)�"OP�e鄆���jgf��5�BpkQ"O���Ů9�<� &ڟP���g"O 1��1"Z�X7���͋4"Ou�F�M(��ROS�l��"O^��6� �30l��$�(d�W"O��[�"N����$c��`��y;$"Ot�ّ$�Xܸ,)e m�����y��[�	@� Z�`ƕ]@p���y�aĝcjlp!��Z�L�aS����y�ҁF4b�
�f�n���Ï�yR���$�"	#�
S��@��ᅳ�y��[�#��;`H7\#�͡!Q��yB&�(0l�X&c��e�Y��lU!�y�]l�p5U2M��a2 I]�y���an����/^!B�2A�Aڢ�y�+�v��0p�E�t�ZW��;�y���HuYUaE	A��!�v�'�y©�>*)�܁���;�N�C�JW�y��A�hX	:pf�$9H�)���y�S�n�x��ɍx���d�E:�y���8�y��Ƃi����#!��y�N <HA�q�H��\چ8 n���y��3.�x��kL�X-4�g冮�y��6U���C`�Z�`0����y2�A�n���a��]W�(�F��1�yBO)��=k���V����ybX2r��P,̅G�4IS�M��yr�"gd�Av�H;iFB�YS��yb@'�4�) k��+#|1�;�yr��!s��yh�%l�nE���:�y�@_hf���+߃/��tIp���yB�.����!U�U�N���yb�� +�T����(b�	�w�Ԧ�y�ǔ��.)zt�C�_y��R��C�)� � DF�U����_8����d"O��
7�	��N0q(��b|�0"O��",�/s�4,@�@��:��0ȥ"O�ɫ3�D'�@H�5	Z#4��b�"O��v�ύX�jAx���0���:�"O4�X�!\�D|��2�h�i�Ѐ�"O`��a.u���S0I��l���B��M+�O�ĉ�?1�1OV�)&(�#g�Hx�j}��H����=H٣2�Ă}Щ��mF	6T�(ʟ&�	�%l�q�w����b�Vb����3Qs6��I-��jT��	M&p��Q�$	���~�t-��&S��W��x�v��0>tdqKY
N~e��48�l�v����)��O��$d���(!IP%-	�Y��O�#�썐�#�[�I���?qL<y��ԉe�4I0p�ȾC2H�:s�b��զ�3�4�?閺i�b�O3�4P?��W��H�aפ�o�)�O��\����i��y��'�H����ݍR��a �A���4���-�'�D@��Q�͛v� �Ѩ��(ORYe�03B�����.�AH�'�uXT�BEQ���铱��p��t�X� 1șB�{��Z��e�]���ˌ4h���%��vO4���'5�p�2LF�j���A̟���qT�>	&�i�nc��?��3�0�����D<5�b�?�?�iP�$~�,�nx�4�1oU�7��OW �]Tk$�	�2��3���O��d�%w�DD��&�MK����2TeF�a�4]ra�������`!�Xj�ȝ� Q������7�򝐒$�plv��@��~��Q��Ú2ŶM�үѽW&����R,Un�8 �D�*�rbk����up�Z�ϗ�}�Dq�SA������?�������O���3C�2d�в���,w�ݓM�x���9}@��c��>f�z����u�X�W	�M�-O0���e����	~�S�?%l�Dp�%�â� K	�5ځi�>2��Iܟ\Bbߕ~��5�N��@xX���?3�=�G��|�d��rTD��5�I7[���o�_�Y�����Ǘ�3H��H��m�n��U��A5<u��OF"���U�~�`A��842)#H<�4��⟤p޴C>�>-���l[�U�t�P�X�%�k�T��=��-��F�� �#��9B�0���G���x��z��`m�㟔�ٴ�MWaD�r���j�3˰`(CƙfV6��On����\�'	J�z爒�V��pC�79�0+�Y�A�(�
�.*��Hs�N�g���?�rr�J fv��+W�
� dK J���*1.�#m���1;VK�`��	+0��=�<����g�݊"�� �c�kw���R�$4��h�i9�ʓj�J�i>��ēh�f�r ���U�q����3%x�Ey��',���2=��� ��dӎM[��>���i�06-;�4�L�I�>�撇��3��_\z��i�� ���nӶ��D�O��@cj�3	N��A3+��ub�ْV㘐5�,%�Ҧ�ǂ)ʎCTE��U��ā�1�ɼ)�j����@!Y�����Q:,��J�<8sH�����!:n$PօM�KڶQ���i�qO.u �H7{ ��e��]@�	��A�$ �"�x��'�D�I�� '��n����p�d�#|N��`���:$���	%=�\q��H���j�+ғR�Q��i����'�D7m��%?������Nѓc �  ��      �    �  +  �6  �B  �M  �W  �b  �l  �u  ��  f�  ��  :�  ��  �  &�  h�  ��  �  1�  o�  ��  ��  5�  w�  ��  ��  �  ��  { { L" /* : I WR �X /_ oe �f  Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�� |d��"O
`�(�;���8���-0��1%"Oj4��ND^[��"3/9�0|H�"OB���H��*�ʞRy=a"O�味V�!X��!&F�:J�$���"O,��a
���C�Ą�M�"O,$3%o�-���p���+Ն�:1"O��ݢ1����`���y14]2��i�<�6��{_���c�H�`�fX�$Kn�<��A̼VI�xR[�)�Ć�pඤ�ȓA5��('nߡ4�� �)˩%� ���,��r�؊b#`T�eT09���ȓ!�b��g��}�8�F��-? �ȓ
K|m�ș�VṔ���2�%�ȓ"R�X�j�4JN�1�˘X�i����̹	_�jZ��1!g��zܶ��ȓgil,*�J�
j�Ne��i�J%b���f	�(U��:���G��$Y^م�~r�� S�%T"���k\�jx�ȓ|4�1�îJb��@ӵ�ݩn�V��/[`�"�v4�R�!ʎ<��M�ȓ`:��z�ؚh�J�Z��$HY:	��H��p�m�C1��!��B:��0��EnjZA V;9����J[
2���	��4'J�EA�IVW&��~�(aZ��ӹ�>� o�Y�|�ȓ�f�A�
Ο7�H��M�$�����mޠP����/���ANXo*�ȓTv�����{ ��-7�*h��I��sB�8�8���3����ȓNe*M�悡;������X�o��!�ȓ'lj�#F�m�+R&;�|��2)n�C��0S4���T:
b���:�0!��e֊��)��ͷV��,�ȓ0�&�8#���� ع�L�����;�P�AFd���,w�6d��r�EQ�( �gVlɦ�M,H��,DP���|�I	$G#\���Ex�%*�S��F�N�~e14l&#��0ɠ萑�y�O�:\q�8P�� E*U�æ�y��X���}�'Gӑomr�c5�y�O\)𐥀��̩7�.���-�y)�*{r��ܱ'F6��E?Q��E{*�,������ ��z���_�a"O� I2�ú�]�s��J����6�S�ӡ*�ɒ�wF
�ؐaF�S�B䉵�:TQ�(���*Ċ8:`�C�I6�~���j ;A]��G��+%B�I�FA�ٓ����+��ʷb��C��>@�B9��ϒGA���&a��'��C��;,��#߁y���J��Ǚ= RC�^``±��9:����T���5�B�.5!x=�@�rɔ����X�9��B��N��yr��+H|)�$'�I�B��j�P/bX� �O�4P�B�	���Q%�>���A8�B�_C�yV��<h^|S�瀉,�B�^���XsjL:l>ђ���I�B�	-�X}��i�2۾@B��{K|B�ɩ$�浃���1_�D �d�[�u�6B�	�c6�X���d;���m�3fjB��"p�V$� Z���� 8���� �q0#���U�>�@Ò�&rlQ"O���d�NR�X�aM�+*$y�f"O4EV�m��T�UW	)�`"Ohq�7ߴe�Љ�✚	C�(��"O)��%1�BI��l�_B�q�$"OPp���U�mV̢���ђwJ���yBoƛzt^DAR���	������yb� mǚ�B��O��ҁ&_��~��)�'a�(E�s�'-�p���ϋ@D��FxR�' B\B�g�		,��s(D����	�'N��yV��y�8����aĺhp	�'kZ�)��[�h�`#�� YSʬx�'�Vy2�@K4"��=3e�דd��t��'Φ��tk�`�
�ZC@�=Y�X�	�'| ��'�l�F0{2.|�,0��'a�J!]f��{�k�<KLyǓu~�"<i���b��;"M	.��ء���m�<�v-]k��y��?�����g�IO���O�t��M��rYC��1�ؐ��'-��ڶ�	�d���c)�I�h����~؞LATJ 6��r�H�}7��0\OT��y�N
�lc�,��)V!If��]�y���#L\:�〧|�����J%��'qў�O��,�A$�BP��*�xk"U�'�,�� -������nJ�Qc�'\a�!P�j������*fC5�E��p>iI<�W!��Ջ�L�:2���j�J�<	�_����m��{Mnh:�/F�'�l6�:����>Z�8�Xc ��s������]���:�OVQ3���6q�԰⍗,�^D���iś�/0�)��PU�.4�Y��N3qzw�#D�0��gƃ���F�B�Hp��_k���|��� ��E�����FB0Ec'ۈ��?�'XЌ+�����Ĉ��9�f(j	�'@|�9��W�\'0�"#��G��ʝ'�'��)�;�&�P#bPK�Vm�����H��G2V�h`��C�X���C�.��ȓL�Μ�s���XQ�\Jg&��H	��Z4��QWH1,�Ũ�o�&W�t%�ȓl�9�G��{�	�TeLv]��?��}aҏP�-=�U����]ޭ'��E{��(ش����LF�E�	��y�n�4x� �$B�I�Y��a��y��mc��"EOo��-�6d���y2�Yr��1 ��%\�h��uKQ#�y�CF=c�!�%��YĀ��7����yBV�rpfO1dRe�0�T��yb��OS:�Y1I�.q=,��F���ybe�A}���O�vh�H6���yR���4�ly�C�M�m�f�fO֕�y���$�D�1�۫i��<��ۖ�yRKKDF0@��:N��[sM�y��n�+â�XԽJPg]�0?�.O�Bg+�[I�)&�Ur���x�"O��	�B_�hWz��0���o *�C���7���pKR�I0.yi�^�Y^���"O��Ғ���=���~��Tr�"OU2�oͫI���Qp�Ԥ)n
���"Ob�r�'ǉR�qau�ȍ_h� ඣ:4�R��O����zR�R�d@X��2&$���/��� �n�P4��0�0��sק��B��>e6 �2�#��R������8Q_���p?��N	f�>��vě�us
��tOK�<�e��[S�}�~\�e��`�<� 0��#اV���"�)6 �����d0\O&u A�2�����G��<��誀OB(�� &�����_˾0���D�<�Q�Y1dp��Q%D�3C��f��'L#F�%���,G��ÎYa�y[BE�^��C�ɵN�����B�T�\��mސO�pB��.5��[2��e��2ca3%ZB䉰[�J�Zg-Q5H$F
�c_�#<!1�'7L\b��\k׊�C��SH�z�'g��Bw���
ƚ�c�����A�'֠��Bi��.�4�K�"4P��'4y�%(M���1+��9w�Y��'":���c
KΆ��ң]"Il�����Afyr铆]EdQ��F�TE�s��,j� �L��I�s��! ���U�0��D���|o2����O�� ��
o&���D� "�k�"O��s$��t�Kv��7O$�uA"OҕC� �\m�M�6�Ֆ[�l�"Oth(RkC�&�\a�s�1V��%2O�Fz��I�, �h2�잁o;��c�I
!��]QX��r�
�u��I�a��V��Itx���C�L>1Yr����4�s�%D�ț3ɖ�^�ؙz�΍;3̺t�1�)D��Ac��6���*H9�����G:D��1�ݟfB.�ps��:�r`7D����hY8��H��P�Ls��X�!(D���n�5��0��'f��aZ�(D�0G��W�F]P�N�y��0{E�%D�h𲈆��bł������@*"D��`͞�I`��`� L2�m�!�$D��J0�.��' ��3 4��a!D��a���f`"#��ʵ�P���>D�h��
�;Q��J���j���� D�@{Wj��Y���*��(R����A D�D�B�Va��IW,�y�ǥ0D��ip����\|I��b>-��d��y��ɱ6��{������`��yrh_0�<�W�Y�	3�����yB�-�z�XB�)��(􂛈�yrn���,����)j:y*c�M(�yB�#jڰP5f��q<҉�B���y���mTMs�Bl�̼�����y2�[:H�ȩ�bR�hҞH�Ѐ��yBK�*jpl!�A�)�0��l��y! �K�Ng�iQE∃c��ȓMFz�HF �5��)Q�.	�(^B�ȓ����A
�j�識��R<{i��ȓm;9[c�����Y�!�M�M��Ʉ�:��݂p��2��!�&�c�6���Tn��aHH�%3�ղ�(��rL,�ȓYY��§���0�`Q�"�U)G7�<��:��$S�`F��A�w��y B��ȓ"����4��;B`@�T�F~���\��mS0��c�P{U��_:T�ȓN�b�YS���WiLQ�#	%xn���P�Q*3�Y+x4���N�,!�洆��nx�fn��L�����	?%GZy�ȓ*�nT�f׼#����s�W�]���:�	*e�M�C8��Q�ʛ*QP4�ȓ�<m�W  (e.�ID�){2��ȓ��Q���88���1�/أr����ȓA.ʙ3�"�7XL����B"D��L�ȓ{�N���]�L$��"`�R�#K�p�ȓ	)ʈ9�c�I�T��@F�Rߺ���S�? �1R$e�3�d�� U���"Oa�$bE�>;��Y�z1�HX�"OBy��F��!�(�!a['J�z4�$"Oj�ʡ�m9�6�^�>f�M�v
0D�d�"�ι-D���#6=j�� ���O����O����O��d�O���O�$�OF��6	�+�mC�Eځ1�"��'�Ov�d�O��d�O����O����O>�$�Odq���^s�j�Q��Z#B�A��O����O��d�Or��O@�$�OD�D�O���æ�Np�����x4V�3��O>���O���O���O6�$�O���O��YQ/[!V!���C��Â5���Ol��O��d�O���O����OR���OF��T�ߝ
/�0���U1!�"Q�#!�O����OR�$�O~���OR���O���O`}i��8'�x�s��bN�d�F�OZ�$�O����O��d�O
���O����O(�	b˧B� �sށX� |���O���OR���O��D�O��$�O����Or�A����?�����[V�
e����O��$�OH��O���Ot�$�O���O��i��_C�Zi1�n��`��O���O���O����Ov���O���O����'K�  �*�:�2-���?Y���?���?��?1���?����?)���)��h���d!��"h���?���?����?���?	��?����?��Ɖ�rr�t���2)���0�\�?����?I���?����?a��v��'���Wf>4)a�ß� 隵х�Y�x˓�?a.O1��˓SN����.1������9��G4e8����O��nZʟ�$��
�O�Qo�=4pa�P�S� �R���g��L��4�?q����S)\\��?��ߣ\�0����C~�*�/IN�E$n��$a�A���'��Q� E��ʝ�i�0�y�M��x����ү��7��1OX�?u ���K6��=�"�rK�0�m�d��қ��yӚ�L}���I�|���' �;0�ٍ%,��XD�K���Z�')�]"B���y��ĸ4�i>�I�C��Hɧ���i������K0���Ty�|�D|�dL+�󤇔`f��vN<<a�ոA��-tAx�T)�O�o���M��'��I�N�h�ת�1�n�6�����
b� Q��z0~9�|���y6�9��zdҀ,�+� Y:�H]9���)O�ʓ�?E��'q�d�C��-ޤ�6��o�x�K�'x6͝�
��	,�Ms��O�̱z��O���Z'�P/8s�`��'��7�������/gi�|*��2?�F�ßq$�y���cQ  ��lm�\�$��t	����Ԋ$��	���A-E�����mK�^f��9n�.t��
��%�T�S��9G��e �ڷD����AQ�I�7lW$��-��-qM4��Ч�/k��߽P�X��F�8� ��>V�>�2���V����Ŋ�
p�p�Å�Ѻ"gPY�%ꋜR��`��R7F�v}˳���B��ID��l�ZP�!��:M"��y�,�'.
�! x��䌻4L�pw`ͅw���x���,az�h�G�m3���*�=�&`��Q�%HZ���芣Nϰ�ũ�j��I�Qc�V�|�ܴ�?���r�4�:ՙ�\�\o�aJ%����kC�!�M����?	p���<�cX?}���?�����j�f_}�*���H�#? ��i��}R��'e"�'���O�B�'F�Ӿ4�1�V���dtT�7�N��T�	�4g=,oSq�S�O.�˚'5v��˱���ʙr��ԂWgH6��O\�$�O�ax��<Q)�h����8C�?��1�E�y�$$)_���'���(�� ���O����O ���m�x���[�ny��O覩�	(��<����	�����+�$*^�V%pQ*גv���貋^5�XY�'5H<�k�(����O���O����O���Gڢ��A�t X<���2F�"m���?����?�N>���?qU.з6�b�%�vf-�j�p{������Q~B�'���'���' |{4ޟ����皕V-��&&q�~�(ûi���'w"�|��'vBϜ*����ܴ�n}Y1H �I�<لcg4�Q�T�Iڟ��I�����K�@��Ο�I�/�v���h��X����I�Y���4�?1J>����?�vm�!�H�&��X3膭�}�2�5\�U��y�v���O$���YC����'j�\c�,R�.��x��fz�����4���O��Ċdy>��sӪA" ��B ��R)x�Lр�iA�	:l�Tqi�4���ʟp�-��dR,v�2Mc4(�cb<҆.������'�����m��)*�g≢[�{@�i��hZ�m �7�ȲD���nZ��|���������|�3`K�1�'�u^�E�B�U�Xs��#ս��	ԟ����?c�h���Œ"�O�Đb��4��th۴�?����?a*�zn�����'��I
�o\@9cgGR�.a���eEI�,�듻?��D]�<Q��?��.��e`P���A�
X�M:F-&)��iroAC�O���O����<iP�W�#��ӡ��>_�Hl�r�>u�f�'��p�y��'���'Y�Ʉu:f��e�4 ��@���X�BÞ����3�ē�?����?�.O����O�����ϳ�Լ*7��wU�5��%�3Q�1O��$�O��d�<�WlW���	Ű�f�$�	"N?� �`�2m��I�t��̟l�'���'e������P�ISc��1[l�Ң[�\��ٟ\��Vy�S�n�f���KU(	�+4��Pd�W�n�*(	����!�	���'��'������4i�`�&4����е1�����M����?�(Oȴ�G�p�۟@�s�u�@.D���q� �t�`�r�p˓�?��"D��|���n:� \�Qa�Ȩz�Z��Q���P��Ǹi+剋����ڴ`��S��h����Đ>M8�Ï%��$)�CI�}�v�'�� �/$�)J�g�I>.��sÊ=63&\C�ߤ.��6�@�Ma��m� ������$���|�Q����MH�+I�\n& ���?�&&é;��Iǟ����?c��	�[�\����D�F� 貅�]�s�4,R�4�?����?)�bW�1)���D�'a2��.@<@�(Ͼ[Ӏ(�)Ń=�0��?���"���<����?Q�����$^L*��� �� B�pAq#�i�N(�"O��O����<��G�-6����>�`�b�I �ʛ��'*B� �yb�'4"�'-�I�rvApd�*�d�8�?1��Dk&�����?���?�)O��$�O���D;z~��1M44��"łY�:�1OH���O��ķ<�5����{/���d��<ȹ�B; ����D�I���'��')��ˮ��Hr^�i��)k)M�@v�u@0S�����T�'H�k��b��S��(9t��1�v��O���=�beC��M3���'���\���xH<�����|�#`N�O��ɱ�O��I\y��'�hu�cZ>��I�4��-Z������@<����8�8�}T�D�G�'�Ӻ���1'�$A���>[��qq�HZ}2�'Oa��'R��'�2�Op�i�k���̡���Q�_�P2�c�>�(O �Z��)�)�<8���w����ؚ"��/���ą?���'Z�I�?A�����'p0X&���A��+$�ƈe0$t���>i1��^���O�b���Pе#���F!.����Ճ�x7��O�D�OXhR#C�<�'�?i��~2��BU���Q�()Y3֤q�2b�4�-�ħ�?!��~��M�U��)D�s8i"#����$�|.pʓ�?I��?A�{���\�$�Ъ� K7�\	��4����B���AV��h��ҟ��'��Q�3�N���^������	�N��@�_�$�	ʟ��Iz���?)E�:,�8m����mc�������0:�by~��''�[�h�ɱ]}���'Q4����J	)�źfJ�A�0oZ��,�	���?)��M���5����zG�.@�t	�V�X�f���"�>����?�+O����sӈ�'�?�#�ʏ�0�'��[���6�S6!����'��O���ߏ"M�$�'�xB�iߺ��0`ܔN�j�� �Mc������O�9�%&�|���?)�'8�H�Jqd��T��)W#�� ;E���O>�$�.j�1O��>@�P�DN]b"��1�� "wd��?A��@�?	���?	���(O�Ņ�X����\�rl�`[+|���̟x��,�$�b�b?q�rK�0����L�DO�Q3I~�zq����O����O,�$�����|��L�Ȉ��h�VP��(�Y�MAc�i���2%ݵØ����D��H�#g �	�̥w�܈?8��o�ן��I���ۡ�Fuy�O���'��D�~X�0����2�ݩ�: �<�f# m�O'�'��D�����c锥"(�b�O5���'=@	�DU��Ip�	Q�`�������0Uu&�;�,6��'�D<�®���D�OP���<y�0�H�갃΀%�<#��
X��.�-��d�O �$�O8�`�I>N��`�"����Aj��Υ�x���9�<��?����$�Of�5c�?���
u҈�s+u�P���)zӪ�d�O��d?����\{c�Vǔ6��&��`��:5@k �?�����4�	Vy��'��A!�V>���]�f�a�aT.*Tt���Î/~���Rݴ�?I��'S���M����@������U��@b$6b]��n����'��LR9{���ܟL���?Q�!B��Yk��	�jP:]&�)W/��'Rd?�P��y��n9�DN='�N��Rʘ�̓<���ӟx�4��Ɵ��Iby��O�iݽxso���aS)O�x����g�>��dB�e�h�{�S�[����vM,Z�D�ႋ^�2*��l	����	ß��I����[y�O��L5���M���Tӑ�F ?�46-IWrD������H�LI�&^�T� e�tn!p^���ڴ�?����?!P㘖��4�~���O���[���d�%JHu(托h&4J�y�JF=a������O���8%7����K
|k��s�.��������,%��'ab�'����މq$�I�L�%�𔠱�B9��Ɍd�n�jrH;?a���?�,O����r�Lۂi[HP�׋��s<B���<i���?���'A2g#
���t�V��
vf�n�x5jS�S���$�O����<)��!��L��OI���/cCl(��h��`�%�ݴ�?����?1���'U��+d뉭�M˅�˟+5�`�Ā|��D�Z���	�� �'�b�'���Ɵ`�իD�h`X�2�� �
��TL!�Mc���'�ҮG;����K<I�O˚&9)왇W�~��]ʦa�Ihy��'�b0��U>�Iϟ����5���A5l�Dܩa!��'PU
���}��'#��
������|Q�Ő���*j,Ӡ�&��7��<���E�?����?�����*O�NތJ��#���F4�Sڧ��I�X��!\#/�b�b?-x��*u,n$��狧��5`�|Ӵ�jV��O��d�O.����L��|���[�e{�� `��uC #A�P��2D�i"!p�� ����R��Mc�? x�#ǆ(@��%��(μF��)4�iD��'q�Q�%��i>��	����/b
ݑ���wʮ\+c�A�*�&\��dЗH�ء%>����X�F��Jp�@E�l;�C�e\�Hm���N�iy��'�"�'�qOf��Ҿ)�≛��׆M6��C�]��`���Z@��?i���$�O�Ҧj-Rq��K�* h�ۃ�F������S�$��ߟL�	K��?q����Q &x��H:����B�&���]X~2�'(rV����$g���'W}�Q"�
�(P��a�B��DQn���L����?���`����&��Պe�K�I����-�}άC��>���?1*O��d(0���'�?	¥� beP��l�)U�$�3��S��V�'P�OH�$�<K��d�x��,R¬R�%��rӴb	���M�����D�OJ�!�G�|:���?I��QȀ�q�J�_MxdӴ��7#.�����OVQ����U�1O�S)��!�eH3x��g�A8��듮?�CS��?���?����)O�N�6 &btk4�ќs�A؆�d��	�t�q��+��c�b?�xq]�d��e#!D�C��e�lp�l H`l�O�D�O��D�����|
��M�h�Xc��\�\��P���*9	��i��if�D�������dD,#��`5�\i�U*!&Ɔ�n1lZΟ��������Ŝiy�O���'����c�c,ǀ.w��#�	أ>��<�,V6A�Or��'���&prl�����lͨM���B��f�'2j�ف\�0�I��L�	vܓ`����0l8��&e��F�0��'�բÏK����O\�D�<���j��K�jø%�Ո@力5�����8���O��$�OP�����X�4i��^�H��2o�.K��d�Wj[9>��?Q������O��1�?�"E��R ��P�I�at�5ڴ�vӶ��O���,�Iџt���$;V7��_�{�7l7:�(�K��.�������	uy��'c�D��]>Q�	�/	h�0G�b\,u�FN-oV�ڴ�?ɋ��'�~`�%�ņ�ē�@iJ�B�T�p1c�͕g�qo矌�'ob�GQ��S쟜���?��d��(_���x�%X0b�p,�v��>��'�2�Ā7\��A�y��`!̈H-L�d�՞g�����[�@�ɴV��t��㟤�	�|�cyZwm�	0g��'Te!�AEE:A�EI�O>��V�k$,������Ŷ[��X`�R=z%���-�_j�f#M���'���?I�����'��Ƣ_�8�5i��c�vI)��l�Dh27dY�1O>����~,�ZF@Эd�H����]H���4�?����?�ШE=��4����O@�	&'>ٻ l��Q ��a0�
j`Ƭ��y���[�8��$�O��I51h.�3PB�z88�wJY$&�D��K)OZ�$�O��$'��u��"��.+�	�U��R+�en^�V��P~��'��X���I�YW^$����T� �S���#	*��6FyB�'���'�O�@�G+�!ap)]7	$ �1c��C�K�íyh�Iן��I͟��Iğ���U��M�pKC��J���R$!�Ҍ"A,T ��V�'�2�'4R�'
�ȟ�Uj>	�B���a��߂LD�m3EL��M;�Ă���?��X?�
��8�M���?q�c�4	; ໦��Q�<rS�6�'�B�'��ܟH��EAܓ!:��SBQ�L 0���g�VMmZ̟��I�D��+*j��ٴ�?����?���5���Ǔ4S��5�6��%
�<)�u�i��U�T�I9x�8�Sԟd���<a��s��q�d�Ѭ���ӄ�3RL(ٓ�i�B�'/�e v�i�Z���O~�d�>���O���b�G�D`̚��9t���8oQ}r�''b����'r��'���
�OH�':�K���:I
�E,�&m�@n�t@�Y�4�?I���?��'�����?���_�֍8�o '?dn�Z���?#���R�i�4����'�r�'��P��O�Of��_�9�i�̊'���C M��6��O����O�uHPɁަY�	͟T�I��x�iݍA�E�"� �6Ɔ8B�Ѩ`�'�	(��b�d�I�,�	
������E7,����C�$es��ٴ�?����8{��'Ar�'�"a�~��'��J��M�Jn�h��a��ѩO��0r1O�˓�?1��?!���?q�N^�b����ɓ4j���h��j�6�遺i�"�'DR�'-P����O����X$:��� �Q29����A�C�0*�d�O�$�Oj�D�O��'.'��'�i�"y�j�&*������)-x@
rӮ��Op���OJ��<����>�ͧV��$�SHY�c�b��M0x8a�^����ٟ,�I˟��ɐu6��ݴ�?)��8�jm�$2t�����Ƕp�����i���';�Q���I����Ɵh��<NRI���4ua ���@0Z�n�����I�$�	�\��޴�?����?���\���C�G�f�N9�"ǌ_� ��i"S���Ip,�M�i>7�RP�����G��9�1�b,��X��'�RbФa��7��OT���OR������'(_�]�#�/>a��s���mX��'6r.\!k�R�'��,� ��ԙ~j�n�B�,�׎�.Y8���a����{�4�M����?A���B���?��?�� ���r�.s�����S��f�۪LY��'u�eɜ�������O2�i��\�'E��!wC�+YH�C&Mv�$���O~��W�G�T�n�����͟p��Ο�� Y����e�[ƋBN� 7��O6��^P�S�T�'>��' ���h
�E�*a&�<O�����i���p-<	l�ӟh�	�$��#�����Q0�&:(���R�:x��B�>� +v̓�?Q��?����?�s�  ��E� s����D2���
Э�-S��'KB�'`c�~�-O����#ys@x�
��������[ K�`$1O ���O4�K���O0�$�|:� �^ۛ��?��͘��K��ճpK-gЮ7��O���ON�$�Ov��?)C��|��-��4��A2�nG�H�=���!;뛆�',�e�'�rg�~�r(T�gK��'|"�Fc�e�E�G�x���$�,2��7M�O����Od˓�yBI��|�M���pA����1+ɓh����c�����Od��O�m�p��¦����`���?C���U�n�X�V�r�$���mˠ�Mk������OpXc?���d�<��Iy�H�4d� I�D��C�e
R�`��d�O�������)���L�I�?������W��P��4;��ĭz�zH*�d	����O���W`�OXʓ�Lhϧ��S�0���R4M�����46�J�fx��l�ʟL�	ϟ����?��Iɟ��	4L���y�o!ӄ��bc�;Uة�4'�b=),O���|����'*� HP
A	})Pd+d��<���"!h�:�$�O<��͝W�	m�\��ş4�����	`�L�u2k^��d�r�J���!T��i>E��џ$��9�
=�"��%ؐ�ow�-��4�?�
O�x��'���'{�~
�'x�IĪ[t�	��6��5��O6	ؕ2O����O���O��'�?1ǨA��>m!���e+��9QȈ9��i#"�'L"�'맖�d�O���l �+B8T��*4b���S0O���D�O���O��D�O6�D�O���ONЦ	�&�ߒ	KHU+s"��d2й٦k��M���?���?	���D�Oн��=��L�Q��B�j@Y��,2��L3��CǦ��	ß ��ןx訟bU3��증��ş�#$�=�V`k�ՌK��4���:�M���?������O�U�#8�����|�M@Jd4QqHP/t�`���aӴ�d�O�d�Ox(�s��ۦ-����	�?1`3�h .�s� ?�Z�x�H�M�����O��2p5��$�O��r�;���oV'?�B� ��՝6�č:��Ң�M�,O\���n���꩟N�D�֝�'v�Qs��1etnKਝ�Xd���4�?9��	~����S�'S"����,R���g�R�n2@��`�ݴ�?1���?��'P��'�R�X(k��"� # ��rOD�:�6m5:�$$��S����s��.�qCC-�IM��Y����M���?���#�97�x�'&r�O�ATR	1ؑ3�  S���B�i��'��J�:�i�OD�$�OUa��6���f�
�~K�,����I??�R@�}��'�ɧ5��|�jx��$�*64+�'����Z��J�d�<���?����d�/]d��/U�3N��b�*Ib5�"E�~��?�N>����?�TEׁKۢ@��葈#�Б;�.�9cg������D�O��7�i*m�\��'8X�l(w����l��?��'���'�'���'�\ȝ'w6k��� ���+ƍ^#6m�E��>)��?����򄗕l���$>��O��Dp�n�Y�^y��,��M+��䓮?!�
��|����ɪ��p�ŭ�0@��1�gg^7m�O��<���4F�Ou��O��x��.�v���Њ��R�+7�$�O �d�V���$:�T?�'�5�<Lz� R��L�u�t�f˓T�J� �i1H��?i�'lc�I�@���١ɔ�m�!iM�#o�6��O6�D�6�-��)��b� ��
Ў[��q۰��\�fo�coZ7�O4���Od��k���Ls�8=�xɑF,/L<;`�N��M{����?�M>E���'��x9�d�� n�!�;*̜ܳ�gӦ�$�O����In��>I��~�Ҽ5���qӠ-��	��إ�ē�?Y�ύ:�?�/O��O���38���2#_�;�r�u�	�7��O��g�N���X��D�i���h�'�LTq�@�&U���e�>�2��<�/O�d�O&��<�E���@0��C�@l�J���<fjt��'���OܓO����O�=��� 4<n��Q揋-R>eZ��O�x^���<����?����d���(iͧ-,]��ïw:�L �� ;�,��'��'��'��'J�iV�'���+M] <�G�^���4h�>����?	���$���X�'>�
$���6� �^)v����-�.�M;����?1��:���2����	e�
!a�1A%�1"c��!s�7��O���<	5eÎF��O�R��5Gذ}�@@B#��t�-� �0��'�i��k���'�q��z�kݼ'A0�Sg̜�k����i��	 ����شN*�Sӟp�� �����i�,EscK 4G�d�.L�J��̣۟�i�͟���t�O"�e�Q3*=����HX�m``%��4'*Js�i���'���O��O��Y�X��Q����}����e��Am I����������;�H����5��q�OX�z,
���z@0mZ���ϟD�v�����|�L�|i��Mw6T�b,��[�t�jrNfӘ���O����B=��$>��ן �ɢgT��ӄ�6#}�-趢�-V ��i�O��� -�On���<9����p��R�Y/h�zd��)��5\���d�<0���?����?�*O��r�.]2p�#iW"F#�Yz@�8�%%�l��ԟ`�	F��!rvTi ΜYװ�+T'K<_�4�K��S̓�?Q��?���?������F�%4��г��2pJ��nû�M+��?��䓓?��%ڹ�`K��ɲ�H�
o�12TCI�a`��p���>y��?����d^�r��%%>!0
� t�I��Q�F��i�!�^�@O���i�ҙ|"�'��L����'���JDC�g݌�aI�%4�JM��4�?)�����:p�(&>Q���?�JdA�%<舋g���+6�2�������?���<,�Ex���qP�:]���{E@��Ec�ui��i�ɜX�� �4yz�S�<������,��2E��o��L)�ӧOg���'��m�<�O�������ő1�����ˇ�N��21�i@�A��r� ���OJ����bT&���I�&�(��$kHBR���
�$R��zش`"�Ex��)�O�ezS��-.��:!	��OP�G�6��O��d�O�ܠ(�C�I֟��I^?F��"1��9� Dr����z�c3���<)��?���[��m*Čķ8y���#�[4V6�Qӻi�҈��?�bO���O&�Ok,ɣu��$�bI#u���S�����|c�����I՟���%X7h��g���po��|p���@uyb�'���'��'���'��궩[>qb�b�Ɓ� .D(��WdD��O>��O���<!�"i��)�1t�N [�%	%
���	�E��I��h�	�(�?��-�g���4d�x5(�Ӎ)/��
�Fб����OX���O��$�O��P4��|�i��u" ŏy"lj��H�L��ie2�|��'db��n����O<���gY�[R@)*V|�s�F4#�ʸ��U-q�Y#RDK�
kl�r��V<�ZA���4v������[���B����
a� �2e��N�<!�"�l�����h�h�c(��c�ך.sTTȁ��o~�A�;V�I��@�
L��P'dǞ �h�`鉈d���A1�՗Z��XS%�=�vX�U�t�wjۊ`��h9 ���1�N(	I ��P���*}ᙢl��80\L�p�I	Bh`��ڦ#dq��K2cZ��-dV����<��)���?���? ��l1�"�&��f%��ȡ�C�[�M��sgR�^:0�8��*�nc>MK�Xz�o�s�B䣂.��d)l�v��?3�~�9�j
��d,�BۈTO���H���ɑѦu;A>�"}�r�\�W� �����D�����-�I�F�����|"gC1<x#�d�8��@��\�yr���bJ�%���b��EQc���y"�'`�#=ͧ��z��9�s���t�T�*BM�i�D�b�-��8&�����?q��?�s������O��"k��� P���C���6&]��5�Vp�]��䄦d����I�0�����g�FP�e�I�u5�T�W���(z�N�>o�Bx��Ɇ����LCw��1 M����$��O0��/���'�<$@!ɓ(U��phd-�ڱs�'�I��0$:��VE�$�̬8�y��e�>�Ŀ<��M6Q������*�����Y25��:�L�K������>o���	���ϧ1� MJ`܆	��eBW%C"�M�
`RN$bb�
�=	�\j"ˀU8�@үD��(����45?�oZ�t~Aٷ䍿:UK���u�r���7�r�'��u�(�jFP�|�"ɚKhb�p��	�2"�)3gD� #�c�k��˔B���M�$�qML�q���z ��BL@��?�/Ot��ԂI�e�	�O`xa��'[�H)wA�jc��p�ur�9b�''2G�<�`@P�ᕫ00t�(���O��\���X3H$��*�/�48G(����4`��sl�J�ȸ��P�O�`eY���wt�P9�/ԗ�RN���r��O��%��?���D�{�P1ѩ��e6�`C�*D���I�@6�#p��1m(�f�.O��Ez�Z��1�G��)F\X�T���7��O��d�O�����8�8���Ox�d�O�NbrL�E_�j���A�Tn�ya�K�`[(y��Z|}1�d2�3��˸5z����$� �s��,G`j��X`���k ����|b�ϤF;f��� �d�� `�섆 ���O�`������4>�BN>6� ��F�
$�Ʉ��&@��M7���b�o���<��'��"=ͧ��xR$ �	�>lȲK\�M����V	(D����?a��?�ļ���d�O�'ljD��LԈn�.�
Z�*_��1�h�^P��>B��
�'�<����<%@򯌩J�A'(M{��S�k^���P���\<x"?�CM�	���8�F�` �y��O�|��	%Ӱ?!�7b�}2�dO�D��y��)�P�<�L�	!n��� I���~@���Cf�w��|���,"�6��Ov��ѕ`�X��@L�r?��L��j�X���O,��%C�OP��y>���JN:nV�����j�Z�h�I�\��8��EA�$&A1u%�D�x��71� ���QH�H��*\��� M�}Q�ud.	C����I6=���-��I�)��@U�L���TΜ�5!�$�/D\��"��!j�4��-�3+!�����)�G"�0�px�7(�lan쒕E�b��l��ݴ�?������Н �D��Y"6@�f+���L�rc��B���d�O����N�
�*%.i"P��5��g��^>C��y��m�厱0Q��!gC9}2��Qa~�� ��!�5x��S���X�%!
����Χ*]p<䎃�Zd4��Pꄼi�2��O�x���'���O�� *41�O�V�rL�vB�'w�@f"Oa[��W&H�����M)��Li��'@�"=��J��c�\xr�54ހ��n�-S���'��'l�ҥ���W R�'Z��yGGʞ;��M��.W�Ph T W4Fhl��+�/��u F`�.gdp�bU��(񄖪c��pY�¨#��ERQ��,�1;gOD�33�;R*��"ɤ�����:�$�Z f���,�]�P%�"��xU�<$�8�"�Oq��'�=��d�-z:�ZA�φ>�tA 
�'|��4}T\�kϐ8,4��O�UGz�O��'~��@$ΒG�zU��Ch/�11	Jb�h]D�'c��'�"*nݽ�Iڟ�ͧrPE�iٰ-ƹ�c.Yu.C�P�T��eؚ�X%HCA�*'����3dL�9d�⠲G%8���s��'}�L�hĶX���O 7Jv�����9^��*�O|�	8\��܁�FST�J�L�A�����O�q��ɻ�����ET2a_�V�S� r����)�$Ť �����Q�?�*J�Ɩ�%A1O��m�m�I�WC����4�?��X�P�@����[�d������0��)"��u����ϧi�*��VѾV�)M~�4[$h _�*�N��Q{�<)����O��-Z�-��B�*���p�*t\Z��s��}�c 䞊.V��?yыҟ��4B����'�l��Ɍ�?ݠe9�%�}g�\B�Q���E�S�O�"�"H����"�֌q5�l��'K�7�$Jj��	e ҼTI6�""�Y�g����<1��P�GL���'��]>�B4ɀޟԢ򆗨�@�Jbk
cQ�������(�~�1& �28ӧ��|B� oS8J�,C�-�F�7o�_���?<���=/,$is���^\�K~#���4��~$a�7!}"銋�?�4�|���@�82W��
���E;�y�-��MpܕP�ǌ;�2m�6����0<y�	�}�N��5K�~��X� ӯO����O��Q��K�m�r�D�O��$�O�n��WTj@2��x��5�N�E�
y�,��C�8��L>�։2s�`
�X0_0��(�|� ��V��9d�T�?q��'�R�h3�3,���*�^(a�����I˟��2�Eޟ�>��y�����<#����%��I��M��Z*6���7]�p�(� #��͓�?)�i>��I\y��[���!�F�� ����jD���'���'����,�I�|R�J��u�����8%��B��l�Y�E���>au�0IF���2K��T�#�J����\���U��$i�]�k۔y�i�'��z�D�'�������S��CѡF��?)��@�p@tC 
�iqC��?Ĉ��ȓJɪ� ��-��w&߮t8q�<��i��'��K$!s���d�O��h�Ζm�����Yt^T����OL����Iɟ�Χ:��5�%��� @����?/
٫�̒C��d�2@֜}�(�b��ާב� 󷣟�7˦̺�/3y�~��@�K��mQDH@��H���ʮu����I
E�����䅣{r�
?�ÒAa�p��C/=S@�2t͎X�!���7���Df�"Mܸ���<�!��C���+��)���	�K�;D_��� ��	=������|����)0���Ds��"r���$1��^y,��d�O�]���L	U�4����B��	�A,�|�/��Q��ݰ(��� �oQ>���p��>�3��,f��FK�=���ަ�(��J|Zs s�5"���vF�� 
D��j,�t�v�E���O���9���2d��*���@r�����(r*jQ�&��v	:Mpŏ���ax�d%ғ6 d���^@�r�bFJx��i�2�'��e�� Qjq���'���'K�����g�B�W�vm�4��	)%>����X�q6Nغu6� �䃥�1��'oH�bb�_�B@�)	���/Ov��@���&� �"�y?��JQ�7��O�Y�S�`����V|j��t*IJYTL��/]~̓I]T\�)�3����A���G�Q?d�F�8l�!�d�,:�~1�� �&)>�ÖkȞG����HO��#�ĉ�>��PG�޸0�8���&
�R���=[	��$�O��$�O4Ĭ��?�����4J7B`�e
g�)/$"T�\+h�}�6F�&�1	��hA�W��<0�j5��k8���D
-ze�|��Z�|ҮA��gGC��Cd�,0g��R���f4�lz`�U���dQ[؟��
_�L
�x�e�k> ҡE5�O*�O�-��Ν�q�������m�d}0!�d@��&��QR���M���?$aģ��c��!h�°�����?���/3)���?��O�:0�1#��]�0����\u��EB�|d����R�8��q9%B^3�p<�e �H�<H�GC�O��l��"���؁�E[Q��pǓ�\�j�B2�� �hO�x�V�'�O����ګW��){BNX�|�����"O� ����b�t���][dtYO~@lZ2,o�!!#���:, i;'dݐw� '�lI����M���?�-���[ad�O�%3��	��(�	��mӶ`�O��d܉�z��/m+,�
��9�98�O��� >�RbG3N��
D��?uز�'۠�8Ȓ)N�j� T;R�hٕ�y��c�[&V8,ɭ;+�p����3_97g@2*芙�O�2�'�ғO����`�2#�舠���0����3"O|X�nϖ4�*h���,C�Hh��J"��|"D鉓S�x�rb���Q?���B�_�PҺy1�4�?9��?ٶ-35(�B���?����?ͻ������ yQ����B��L.9����N�:!:� J��+��OV���3G��<�1B�2 R=��@��=m�j��5$F��Xp%�+w`�	� �ѣTIL�}r��]7lz�I_�p��O&+�9�eA�/iW��@�4"ݛ��'�n]P����$�O.e���2s#�[���X0����D74�8�]��y���9n�y�s̙+Y��ɒ�HOZy���O�ʓ�4\���
r���Q-q\Z�P�H�,U���?a��?!��h���O��S���8�ءREakp�X�Y�|ar��c+n����-67.���L�H�'sP�m@~S)K�Ę�9��4�V� �e��IW$R�D%N� A* �]A�ȅ�N�N$�)�=�'ƴ'��r'�^�8W:�`��_p]�ɫ��?9�$�xg\1����S�¤a��f��&��#��,�(s�ٟq2�xAc�,�	 �M�J>�bE.H�V�'^ҍ��y�a!C�D_2D��T�B!<�2�'�����'"?���@�\�}]�I��'O:,��}��]�{���$�<	�ZГd'ڐV�F~�i<u8��W&���XıcO��Sj,i2mT�eB^�т#R�u$)8&���FY�5��CܓS����ə�ē&M6����c��bf�)c�͇�v	�\����7cr�J�&ؾI�X���	��f��6%M���M���P7��1dG�'��!�7�fӄ�$�O�ʧG%V[��n�+e�6|�P�#�H�:V��B��Ov�/�@����b�J0dίL�D�O�SZ׀�X�nmp�b��3���H��e��?GxE�F&J�{��(�"A�n2h5"Bᔅ�~�I�>ⴜ��͜�@Ĳ������99��$�O��d�ON�?=�I���t�P	f5�*�	ʟd��I;T�`���JT9`T���2����c�'l|R'�����`��;_�,���fӰ�$�Ob�$�4�F�v.�O4���O��4�5[��J+}*�h�`��Āታ	֪E�j۬O�AE
χ]�1��'y��i��F8%�(�ʀA%�\�d� �� nZ<Ji�ڗ ��)�q���s�O�l��BS�)�X�:��^�b�$�� ��f�`�,���|��lً"��G��� �U~�E��5�dL�u�J��$` �$�^��'k�"=ͧ��~���R��_�E<�q����h��p$�<cxD�R���?���?�׻����O4� �|��KL�k�x�-�7-s&q�⃭+�����N�3�&���aR>A�|Á�	�+�D��'�+FrdX7��+j���fD��u2X"�J�]��]�a�ݕ[''�6d�#&�	1.ح�g`�)�����*e\��(�O0�������&
-rq	���9gS�C�	�hz�$�@B]1lF�ku�.@Ьc�$�ڴ��;���0�i�R�'������n������{�l}�V�'�"�B����'��	ٜ'6(Ph��M��}��iD7��@�#m�7B���(W	܎ ���@��M�'`�s�o��y����7��.K�X��n��:y��H��W/E�>�s⟦���bش'ݖ4s�{�ʓ�?���x���AV�h+�ba�6�*V��
�ye"i`\,�ea�SӠ�r�����x�`�p���ц���PTIнXt��3'7����H:�l�쟸�	r����
?�"i��@%;�ے;��if��7�"�'�6���/��vx�=��T������OK�(�Z�ӣ+�mLDAAA;����>	p�!vt:���k3Kt1H1뇈(�@����=L��!=�Z�;�-�W>Ra���Ӻqv��'�t����F�ɧ�Oq�xZ���@@@�N�P�'�RQ8�N��xZj)"OAY�lĀ���D:��!}Ġ�:Q�Gs'B�4iS �M{���?Y�yZ�j%� �?����?�Ӽ��N;7�~LIB����"�S'и%0��`iʜ ����2*�&G�@�����?}bE��%�(�Z�aÞ$�1A�M�rv<8Q���f9�L`ޕbʒ@y'b��Ӡ�p��9�� ���!B�@J2�E$m�tɠ2�Kp�%o�|���|��U� y�.�)u��ɴgK��y��Ȗp˘��֨�qh��m
/��D�b�����|�+��$Л����b�.9���Ρ�P\��*_�',b�'�&֝ğ��	�|z��J2M�4�CH7 ��4�eg�qx����K\����~��tsf�iD���١r��g#����Лg �6$�Z�*�>LO��30��n�^MpA��f�\1�H��I�r�5�Op���Ӂ8p��@\>O�b�"O� P1PG��jk�X{�ޘ:���g�T!�i�йi�"�'fV��HH03�@�7���P�1�'���3y��'S�+"kl���F�������	�x�.YPD�:.P�Ţ�!�+��:�,�H�'m
����[+Y�)�eYw�����k����/GmM�Cb�;:"h�*��5g]�<�=�6���bK<)�
�� n�	��G�,��$�)J_�<9"iS�|bV��b-��k��
f<�նiM�q��G�qr,���j<\����|�êB,^6��O��d�|��?�D�y�xh��D(jФ�H���?��9�4��Ș����lÚO69�a��/'��"�"}R'���O��b�0#^ &(Ë.��X6�>yPLPǟ�I>�ʖ��, �,җ.��PX�E���E�<��T.t�T��,��4U�t�z�\�����pܩyu�գ~p�,�W�[JDmZ����֟ 
1�H�J�&����4�	���ҷ�K�&6�Ab� \�1|�[�c/�
+]���Ę�M��z�� �A�X�!qO��jB�'I|<��a� 3�P1�IN�Ț���'��N����L>bGH%_�BX
B/Y=@ԕ�eIr�<)5���,�ڡ eC�6`�q�'M�o~�%9�S�O�� ��v�)#F��	*
��-�<+.�A��'@��'�"���;��?�O�8�WI�5\��2Jƚ���1BO�K��}ꆭ\�ϼ,YcLԀ��#?�Vh^ M�x�Ҥ�Q�g�L( p
EU��\H��V�Y� �{g�
:Ϛ�6I@M����o<�I�^��DPg��s�Җ��?L�4ڧO�O�$���/>�Ukʪp=��;0�G��C�	�[�.q�%үXC���T#�Kіc�\۴�� C��:"�iOR�'�"5[b�P\��H�u�_�f�8�	��'�b/��_�"�'��I�j�r�`W��P��	�R�t4�wkن>)ԁ�M'{����S�$��!�.��I2D6�X��@�i���¥ɓ-@���[)=2�+�ė:\n�أ��6`���rN�"!�_�~�<�rÅ	+\���MX�q!�d�ͦ	����8	$��8��;r�՚��-�	YO���ܴ�?I����)��;`�DM�1����	�.H�P��FS�R�����OP���٬���A�B�#� �3/H����Y>-{��.���'�R�-Kw9}��B�/|LZJ)S�@%�De�/��K�GJ�_�
��'?o������0�p�Q1"���O�����'A֓O����� sJ�u��f[�Rjz�C&"O�@yWG�9 ���F^_4�)Q�'��#=y �H�u�,�#&%�vۖ������1��'���'k�Q3�R���'����yG���;X��Cg[� H�lµY�� ��H���G�2e�c>�O @�� ���F�R����3��L:`���@\��㌀�Jbq��'�,+��o<F4Ғ��Gl$x��!�D�Gh��L>�!����3Wm��
�(��@*�x�<)Ԁ��Ȁ�ơB�KYt��gCGq~�b<�S�OKbM�f.W?@C�=����N�(A����H���j$�'�b�';bw�%�	��XΧT����t�< x.��~����D2o�:�x�oJ� ���$N��:E~�	[<b�����ηf�0���DA$L�0,�����cIN�cU)O9_/�D�Պ�P�@����d�e ���煬W���7�� +AM�v�
ȟ8���`�d��!<E@�@HB�|G*���v.�0�h�5�@���\]����<9R�i��'< =r�h�b�D�O��7g�9����$�Ig�q�2��O����a��d�O����`�h��L�U�����/�M ��0 ��15��A@�<�)��g����O1�R.�1:~D�b+�
�z �-C�����BA�4�{��'j��:�(F-Y�鉏{b#���y��xG��f�(�xf�C u���3Ț�y2��X?lY G�
ju~y�n�9�x�,r�`��TO֟j��R�KQ�tI����&6���?��l��h��L���1��hԮ1i�Y��.	�[�:p����/���'���&�ì.N1�.Z5	����\r(��Ij�4?�E��,K_��2�>��J�X�r@y� �,����u!/�뎘?P�IpB�f��
,Vh$�%+U��l��é8}��V��?��y���D��;mIW$G	@,�0�eI��y��׀(r�`3	_"Ph��ɋ*�ў�S#�HO:�id�F�L��k��$��h�@�Aߦ��Iџ�ɍ%���m�ϟ���՟��i�a�t��Q�|�)���p�"p$EI/^�(�8Vm�0_�UA֮�A=Ld�|2��>A&��6By�7"�
����S�H�P ��\X��jQ�@�m;�A�1�>�M{�`d�A� a�,$0�A8u)�&TT��5j����WP��)�3�[�|u��q	�!b�1��(h�'ޘ$����
n��piwH-����'��`2��|2L>� @�������M��oZ]�'�ۓ��2�On�D�O���Һ���?ќO��;��� s@�Dj�CD8 {�����S^�T"?QHDC�A�xQ�#?����lM��{�
V
2�q�2.V�ց����U�Xm9�GV�-��){�)S����wܓ_ly�c]�Q�����|u�YcS�t�.�n؟$�'&R��/~����MN����TV>]G!�^�/��E�KH�{p0JIS&1O��mZҟԕ'��`�pMnӆ�d�O$�B��1B��5B%Ƌ�-a�y&+�O8��zo����O2��u�F!�&�1a�E%)
�(�X�`��N�,���,M�
�,C�g���O���'��uf����2v2��2G ر���^�iu*��v�U�+��!{'�;Q/,� �{�	���?	B�x�ȓ�3Ⱦ]�qI�>���Y����y��g�NX����;d����x�h�z\��:{�<@JS��/L�vYq��'�S��y"�YdT�ڤ
��O��;Geբ�y"C� J�H,�Dk
%L���ab@�yR�0J�RQBu��9�r�0f�O#�y��-4���eO�e�� z����y�FUbf��1da�
e�ح0�J��y�OE"��{&��V�2�sa޷�y��_1k�:9	3#®�VY�b�-�y�o��Q�N����>|k�a�e���y��H�?��q�6GΦt�ڔc��y�-#3�2yR4#Оx�.��`
�y�T�a�P�@��B"5؄b�Bʑ�y#%/)����)޵b�j��y�׵etR5������Œ��y�d7~]B	2��6��D���Pyr��9z�,�!V�I�uA��;OM{�<�� x��kT�\�-UY��\@�<Q��ӟ�2�X�(�B������y�<�t@�C9(��T"޶��0�`�Y|�<��
�QRȖ�s��}�ufNo�<I���{G�y�GU�`�z�*B�<��^�a�\�1�Bߓ0��q:
R�<y��˹�z�A�e�[}�QJt�RS�<a���f4ya��3m@���@��e�<i�b#�5J�>e�  �e�<i�a����]Z��D5iV�swd�<q�Fs����7B�QF�����E�<)�O�.	\��� +ۂG�4̉ӣQ[�<P��z��:l?Q碜i���_�<�$��;T���5k�<φ��ELX�<�E [�Q�H�å��7&zHk��V�<i����,���2~؞|pB�I�<�'��KR�`�)Hrl�v:$B�X�ؤ�Ѓ�%�Z�{��}�TB�I�<���#牗a�"����
rk�C�ɨx�J��e�_u�`Av��k���=+.�#4"Δr����)|�B�{��ȺSX�:t�	+�1�S"Ğ7l��9�Չ׺7�%>ʨ0��J	2Yj�öfȫ!��z3�Z�|�Sg��r���p�eݰ���I,�|yð�T#8�vi�u�\c�ʓ�ء��3�P���^0�GyR�P��n��PhS1� 9B�e�1{������F)J�pw��F�S�@��~����+�'�f5����ff�k���F~es�dF3_?<<3dn�[8�;u�ACƬt���4�Љp��ʑW�1f�B��H���Wj,�=��w�|��`ʒ�y�8��A��U�N���l*���s
N>��`�*�/_�}FמSd�:��P�"��'9���B����!��P�t�5MV�S:�&�V3:�2�F��	~��[���	)��Fx"Ɋ-5d�U����<;�|��⟋S�,�S�bV����#@F����bÀ��\�r�) ,�a%;F�D��+\#4�H�$+-ʓ�t,P��M�t߶Hc�f jJ���D�2qε	�a�V����웹^ t-R��]�4_�Ia�n ���U�IH�#��2k��@�E�g~L�[�EO� �
�I�X���F
	ȴ����#B����E;(��ђ�E�-�ހ9  �;��DJ-�����y�gR,4ٸ%L�?M�P�[��ł�0>	�Ɗp�}�5�&?�;��O3��Z�ɱ~���!D����d"#����2���aV<� 8;�8y��I�n�)��ؠ�$�\�Њ��OڐǀČ7Ϊ�G>)�z����QL��9aHL�,��0[��E)3�4���f�/7�D�W�J����E5vk0]�%.C�>ؘ�Fy
� j�vD@?
�H�G���&�n�Q�N 	�����L+��Ijt�<U/j�rLPJH�Cɔ�fg�I�v����U�z�4*N)u'~L�����e`r���q1O��ˉ�D�|���80�	B! �
�A�`Y�-�����##��!�� _��
��� q�,�~�9�ZuQ��#�vف�-L�C�L�)&[�Ӱ�T�'���c�U9m:����ָ()���k٬ƐA���ɺ=�ꍦO�Ä�Q?����?Q=��Xe�?��RgD4 	�@�2�),H�,"�/G���Gx��1��E�i�2���}�"��t#m����9Җ%࣍kZ:B3�����$=)l�x�ҙ~�'����H,�yp��'xD^����E-��R̚�g'�}�A蝪9����,�J��9`���BffY�P�1OX�`u�CF($��'��AB�I?}�>��MX�@��;��:��	,�bF�Cm<a���O�a�$�U2w�=h��|�'Ԁ�u0+�2l��Q�'��;��I��`E~�OQ�<��ɨ+̠� ��-��7�}*q��^��h�)\��9u�̇V�P�#��cL~�íG��u�ƪ�R0]7][J�H���,3IJ�"O�a��Q�i�¤H?IV��Z&$!��ƈ�j̊��`�L�i�`����A��.�[�L}sfh����:��[3a|r��%��٘�癍m��$͐6cP�`���ٔb��+ю���v3�$� )��<Y���ef��SFf�[z,�CE�'�H���hShK̍����"_���Z�S�ֲ�N��d3��y[��Vx}rMe+��0�e�a����M�b�p�@ ���e��y�ΞO���'K.����C�}�i_��g?Y�F�5�(�{S��0�N)H!TL�R͑��J�y�P��6�ƜP�(R�V�ʧ4j�b'��%d�l`K	I�;�b�E��͟X@���d�u�G�On��Ɨ|ch��0RC��y����[y��� �/c�4��3A��~��$R�/[ �b��|��u��<{�P�"�YvNĔa��7���7O�'����'�I<uj=����
V����h\��ŁT�Ƴ9���ba��<, ��k�%��b?%̻_I�{wϔ�s�F����U�XK���'&�)1�Ɍl,��f��Bh�=qU���A_ bR1�bJI�b�Qӭ��<$.3m&���$��?u]��瓞����4΀+YD��3���Lݢ%����Ox���g�#���:�o�DIƋ�|jŪA���(b"j�$q�(88�ϑ,�)U!����C���~J?�~��nZ�fJ�5I&O�j�-B� SM��h�,I� z�`Y$��  �0���hj>5K"G
�A��,@��O�t&�k�<2�X�/N���&�8���MQ�Dʹp��,���8�bJ�I��ңm�� c*V�`�L#�̍4[8 <���2r�r�I�υr?�Ӵ<퐐A�#]>����5��.��K���a4L�Op6��]��s���hO�0�d�c���;@N�4^�X��TJԸG�&1��cܹHti�E�O�<`1�Q�\c�DB�C:,@m(!b�O��O؁��AI�xS�Ɂ�9��
2�Ƀ����t&m�"��#/�l<�#{p]C�BD�M�	(V��dz�����D���L��"�<�H�/Ϯ�3}�ϐp���3�)����3�5�Cס���8wC� e໴kM�dp��'�(����O��4��O
��VS��ٵI܇w����d���#�c��Oo6̓����b�'�<9��)�I6b�A5��:�.x�Că��y�#P���C��0<���J)�^�A!0>�,��.��Yi��@5�E8d�H ���/dK"�	�fG�.���+"�B�>7�e�W%2Z���˾&z�xR�|���>z�PUm֊"aa�T�$}�Fx����|0�{$�ˎQ��-��� "�yB��C��a`�$f
 ��ښ{��Uȉ{b�|2bEsfe�t*�`� /*.m�N����RR��{;x(����1��9���ee^�����r���J	�m�~�;ե�:���kP�$}r�[�5�.�kӠ�)�\(��e���'WI��nrS�@f	��V4���Zi8a}RCm���E�B]r�I��]�+-T�p�/@1�Zu(�-ǽ$:�tF{��Z+U���	T�w���\)2, ��&.��S�i9�A/��(O��Sd�07�r�+"��2��2W��O���ئ!�H�SL+�<8a����$�/M�,�ũ� 6��l1�ݔ\��I=�(O����I�8����fZ�1!~(j��K="���%پ�Iw/AE��A��4�eY��Ks'Q:1��g���/N���<L���6���	�����gʐW�����MԠ%�:��?�薏,�̺��Iތ1G���<�v �L��Е#�����79�dʋ&c��'����J�F>�݉�ʤ!�Hej�	L0M|��)`K˿X��T�0�
���Z�/��S$&\�5��,�e�C;5^���va\��To�=�tj�λ?��:�uW�[�rb��'\n���Ju��T3pCm��'�n�6j"5���	�u�:�`��$#�A"V�	Oy�����������S�S�-#����2<g��r #Ѻ&����d�.|K�k��1��M\�Lɷ�]!.�TP�0p�z�@m޶8���'`�"}�'�:$�!.Z�3:��2��,-�xH�'\r!ʱ)�? Mk��%9�\e��4�6D�so�-�x��DV!�l����*p6DYP&О�a{Rަh����ʅ̟rtGL�!�s�f�̽˕�2D���Kәsڄp��K/��a=�I�w�DC#����>��alLJ�|� G	�C���Gl D�� ���rڙb���I��	��%R .k���%�|�`yr�ӆ=J-�CfP�	��,��i%D�a���?׬��u�K�'#L��c�u�����늵1:N����*qR�mD=#ĖAa%j��]����D�
T�4�a&Q�v*��"���=\JlI��6,OT!A��;88�ږ"���% E�� ]҈u�ѡ�+wde�ҍWH�'tH!��V�"/ݓ��Z�@��2 �~���1'�K�nQ�GAG�剤nI^��A�%q��@a�ώ}�̢<��(��,d��8I^ȝc��M}�oQ {��H�F��n� a
��HO��𦟈>�2����ɀ��Գ�+ɱL����&�iX����S�|W0���	#fc� �
�.90��sMS�����w���1�/V�p.���W 7���*�?<
��� �H�D�R�JI�<Ð�v���S�#?A!J���z��dߔs4�Ԛ�]ĦZ%FK3	�\]�5j+v)�(�V�2��5����5#ư`����)�.�ɷ�|��健i\=s֦V�K��ʓG.�s��I�-.�q��0mGyD�?v����I�c���ܸ�ybq��3�	�!N�̌IL���O�pIg΂�a,��b�J�<$
 �QV�����
r�)�@NIM�3���X��`�p�N�vQ�wK��4���&}1�����(20����4`�~]Q�gۂA�� w	C �a}G
3�l����<]R��	2����O��2cK\.o���-_�y�0�ӋN�
��Я�s�xh3ec�L�C�I�Nꤨ�fH�+*�j�s�	E�eW���^P�Pˌ��2,���W5��tEz�5*!A�2$� }��;�I�\�P���m���S���c���	�s�>�1��Ģh�4� �gȐ&��@3c�S<	J-���'���ċP(qZ�P�E�U�v)�q@?<�|�hwޙ����"O�d5b�F6o�D���E)�O��5�_7e�hh*��'{�L�x����;d�A+ܻ��O>ؙaJכT�#'a�Ĉ�i�(
�	��d�rxW ة�^ݑ����=y7(���$ry
Sȉ?m�I�n4Ҝ���ؐP���1u�J�iW��wF��xp͜�#�
L��%WZ���Ez�a����i�2C0!���0V
mٰ�X��4j	�a�X��HN�mFR��:B�RXvHTc:DѲ�Ʈ�l��'���AÆ�Z;>�"P-يPA�C��P��$��ܖJU��
�'�*����� 4�W�D� �X�/̠yQ&A[�`( �剞p�D�(�|�J��h�S�Z�����+��p���)7
#?� �@�-�]���-��ӡSK�A�ffք$9�|�a�G:��ށˤ@�bnƤd��}�e�W�<�g}���}{�|)@�պ�F����ݗ���[!2,��j3
�,|l�e��ӯw��\I5��!�@���Z�>V6��۵�� 5_>�t�gm#ON�[��_9G%^�``&^
^:,B�┞�򄑹8�ty� �j�3��"z긕�%�T!'�1��B�(����ȼt�pac$..�(�a��<Rj��FvƂ��6�"�O�Թ��/\�	k0._�U�(l�S�ɝWMx �&FH�1y:����"�1-¬���L���=BD"O�����2 (9�q�#.l�Z\�X��֩O��a�>E��m���&��$U�CDU��yB��L������r@��y�AT4��U�N �V�`h=�yR*��d�!�nA�q��q$��yҊ {M����E$�� ��y�OÁ8�FЉw�];�,8�'�3�y���`Z������8Sb	�yR�W����Q׍Z� �v%�\��y��w�\�"A�����(!���ybiG�q��I�Ɲ!Dw(ysNH��y�@�P�T�b�ߘB�������y��D�W���j�lN<2���qm��y��8"�n�ת��K�T�sfÌ �y����'2�� ��[(r��McFB8�y"��X�P����>^���ᥤ.�y�?(��Q!�0V f���J�yBN�} � ���S�����dj7�y2fѰW'TIP�_�D�d9tG�y�k�a�nUZ����9��]�C��3�y�J��"�\)
jK�.	��ز癑�y�읭rv��1�DE�W��1P���y�n�G(�g�Ô_����y
� ��1�@�\� ]:KI%f|q��"O�ՀgI)#�9�K�%{�\@A�"O\���%^����r��H�X�{'"O�q�UM�4T��:�v��|��"O\9󷏈�%+��s.�v�Vt��"O6P���=t�Q	5Kޚ\��-��"O���䙼i�EC+�Y�x���"O��;ä�D�8ա��׹)�@}[@"O�����,.%Ȕ��II�{| t�E"OXZ�o�u@̬�sCט=c��`"O�9�b��;gM�Ar&d�B�����"O�P�sK�'|����)b�X	��"O��aSEO-/��|2��^�Z��"O"��a�+�4��񏇤km�q�G"O�u"���9h�!s����Ilh��"O�4J�C/9sx�;!
#)HS�"O�@;�ڰT�qk��i���"O��Q ���M҂�F_�n��D"Oj� 2�Ӫ7)&��W �Pw$���y2햗K�"!J�KK�|9xVB�y���&<��9 e¾I� P���y�l��}zd�:�%�<;�
�q���.�y�NN����섃[Dtڢ��"�y��E�0�f�ƞ^Q�)I��2�yR`O7\�mi���k�%��f^�yr�Qxp@7��h��!9�ܒ�y�̂3|��ڇF	�^ 
���+��yr*��'Pi�J0P�8���#ݾ�y2�Ҏ�F��@-@P@D �Ê�yB
�+T&����4Ai�(��`��y�Mĥ]2�A�l�Q�<(Q靧�y�F҉s�,@jل@��-;Ga�>�y,�Xi¥�G�:
�1	�#P��yR�
�dY���B܎$$��C��&�y��ɚ^�=	A䞬",�YY�/:�yb˞���ٹB���D��i���y�Z!�Ti ���,���$�yB!%m;H qe�+��5�	��y�⏪s\��A��3 u�H@c�'�yr�ΒpԖ�0@�N��iۧA��yBC��N}����MրDh�Q��ڀ�y�Y{T���U�5.] ��L�yRÄl����/�"��'�_=�y¡�=S.6AѳfC
^��0EN��yR��q�t�
W`S�Q.��pFț�ybe��{q̅��K^�Pպe�*�ybEXT�����.V�"!s�A\��y[�{��(�&��Lۼ��(��y"m 0�@y�!иJ'���CKP6�y�.6��t(�&˱?&:t�3&�,�y�!�*T`�8g�2<��2��S��y�,Ԙ8�T9����A�썣����y"-_�sϜ��Te��80�����y�/�:�MQ@6T�a`��yr��Kra`��5-JMѷ�]$�y�G�S�ك�.
1.��4F��yB�Y�̸uwO�&��\@�E�7�'~ў����I��D2e92Y�$eʖv�4�"O>�� ��gJ2���RJ�~��0"Op��A�$r�ԃbCW/�T��@"O��*����q��I�a�+4��۷8O6��DU�!b�؀bNW�8-L�A�·B}ayR�ɨq�L|#!V����R�{��B�p�0���gޫQ��a��mӼS��C�)� ~��5L��[ft`�$M� ,}�hB�"O&�Q`,�7/<��\_L���"O��	�D��uݒI Eb
�"��y�"O��%�:O��7���G���"O̬�Ïɠ2��i����*r�@��*O�(��fMR�θBpN\�.b���
�'?����m��P*���@��*@bРI��E{���mM 4�`�J�X��V����y��]�8(�\p�b��a$N�(�y�JC�#��e�vo��D$�*p�O�ybFR��qt	�j ʧ����y2,���@�gc3r���6����y"�W�d��8�KQ�?r$��J���y�g�TKE��ΟD�ĩ���yrn��5�^�YA�><Fm���Ɖ�y�M"6Dz�Jc.	4q�$���y�M�6IHJ-�Ã[0XݸA���O��y"�F�����X0'�&(P!�[��y�Ύ/^�襋���G��eV��y�*�2e,��J�j��/�TH%�Q�y��]�w�T�R'P�*}eC��yBjY�c�p��G�
��m����8�yr茍E'��Ƀ��W�����yBj�=v�)��B?{b)�R�y�)�,zL$d) C�D'ʩ1�CW�y�AV�r�����	A�)r������yR-H�Z���D�6�8��u/��yE��e�x���@?����bն�yi�"#"(�iҖ8���cd���y��X V\j�
�@X�&�n`�t�V���k���Ow���$��[���dL\=2�u��'��̉!�"hj��jՊ5����}"�-LO*�FZ�Iz���E^Y���fO������+���Sf�\1��XcC	h�<q�R�2Gb����ح���Xb�<D{b�ˏ^�4�ZD:��sP-V�����p>y���Q�@����f������i�<ٱC�{��Mhы��;~
M2p�TL�<�jY�3�TY�ˎ�{�&Y��M[p�'�Q?�إ	��#��;��d�U�4ғw�a�4��-Yn !�H +�$	���[0�y��S?{�ؔ*��\�!H��"�,I����~�S��y��K�*��6	վʊiJ5���y�`��4z��pFO�xw�	u@�4�����> b�cNT��6.f�*C�UT8�� `� �~ҩK�c�����_/!��J�0�y,79l����HS_t=�F���O@�D�$�ӆ\ {)���ZݺQn
��y��Q�= :���NЫE�1�I���1�O�Y[��)O��9�a�
Af�(�"O�H#��F:M$�}��X'	�c��d>�S��1S�hd�C�l�4�S�Ӛ(rC䉸@jD��-\"Sh�=�$�+��B䉱p&�DbU�ڢ'���˧���B�	� rf�C��j�tYQ�(���B�I�p��EϜ�?FM`v㉪)0C�	2j�J�*Ĉb9<]z����$C�ɪ�Y"�)�x�*=J��ܨ�=YÓZ��yA "8�2��0 ��ȓI%ȼ�R�S�oX�#Y�(�����&.M��Z�X�   H�e�ȓ'j���, �m��C .
F�2ɇ�8���TVe�peR�ra�E�ȓ	��p��3(|Xq�揀 -��S�? Ta�%� u$�AV,�P0Tk"O�Q�eV�&)�2,�)�9pb"O�T��̎�9� %� {�V AR��[�OX��$��/ _v��&a�k X8{�'��8���JW@���F�:)�	�
�'Rx�kBj��S�ԙ�=-&< 
�'G|d�!A�sB� ��/��"ؒ �O�6m �O�U i߬.��{��A.J(RQ���'���;��0��M�R������>/r����eg�Lxׄ���2�Y"�(���x��I�i�*�jP�SP�$
�!��`ZPa�s�Δ!,"�(s
@�VTp<�ȓBϲ���]������̀&�(��GT��W�
�A�f��ʊnL��ȓ�`Y����,�S�J ����''ў"|����$��x�Ǭgp\�"IOd��lZU�'K�P�匟k�*�AE']?����'�|�!�Y�v��e��՝�@��	�'E�A	a��Xrk �P4:�'�~R0(P)���H0L����}�'BQh�)R�m��%j`�ՋjdT��'��Fˁ�r{�X� ���4.��e��y���(be/_(�(Gd���0=���Bd�p�����z��"�yB�4<ܾa	�
�D؛d�»�yr���L��B��B7�E�§�:�y+�d�օ�0�P!>uB��Ҏ��y�e��)���2U�=^?n�����y��9~鸧�I�QJB����G4�y"*80FyR3��[��a�S �(�y�b���$#�	ќN���2�H �?����*�j]��ጘe.hr�Fh�H ��1Vµpc���"G@�"m�����ȓs0�2疬I&hz��Iz�Hd���f�x�A�;`��!U.b*h�ȓ5>XdR*�$dJk/ן�����Pu��O�7ܼ:r+ڑjlن�G\a��O�<X���!�Y>���ȓ-�v�j��%�Qӡ%�3��Մȓy��E��O�r|��rNR��*)�ȓx�<4q�-M&xp�lAG����l��ʓH^�e@ABT�&�~�)w��3t��C�I[�\��f�0�`��Ȯ�yRKN�s�lK���|�d�[��/�y�G!v�2���Ŏ_c�je*ϑ�yr
�g��E)2��[;���t��yRd<sq����Ym�(+e[�y� !�hZ􋖀X:(2Dh���y��ݵ3���R'��H�RyP�B��y��۔d/�ŋӁҨ<X������1�y��u��0�*��@ļ1�AJ�yR�Ķ7��$V�O��x�0�G��y�&��<���e�ݱ8�EPp��y�a��"�k���"H��bI&�yr�1F�B\ɠ!4��hb�gN��y���a�h�A��Yc���u��y�T-v�ѓU��V���"tgڒ�y��K���X
�2R<(�1ӯ ��y��/ra��Zc�� Gn|HV�D7�y��U�S ����A�3�es��G,�y�/��C)���#��?3z!S�.B��yrmIt�L��9�ȩZ7�6�y��?� ᣷�4;��  � �y���Uwȝ�� �kt&�9�n"�y
� ��[�h��L���;�n͑? I(�"O�ٹ���h>\D*�>o�
�ّ"O�����.y� �i1��	��UY"O8 �@��d>�xB�Uw�	@"OB�����?5a���a
QsJbQ"O��Y��()�8�@� qk�AF"O�A���	�s@� A�$޼yr��J�"OE��J[f�nW9S\��"O,HC2JK��$�cƆ�L�d@e"O����b�}�$��
,$�t"O>y�M�7u8���&�PvH�#"O��V�ߖl�,"�ő=r6T��"O�T���E�p2}QeOT>2E���"O�@�a�H'n[\�N�{;|��U"OT�p���f�ڐ�҆�	.�)[�"O���*D�u*��V�0%B,�)�"O4A��X'O�	r�n�
\<���"O����C�3���A�����"Ov}�E�R(oH��V��`�~,�"O
)iT�"�����بB�� ��"O�"�(йo��X�,�#q�51s"O��xk�I��H`EQZ$ep�"O�5���yh��BK֑Un��s�"O~��
�b(hHѷ��3j��[�"O�U �*<w��6��$T�t�"O�yH�+[hՈG�M>U�)q�"OBi�DH[�o�i�2A PQ ��v"O0$X�EI�U��x����v��r"O&�z��Q�"���C��<�"O����kT�{7m�cު���"O�����>.9lU:%� 0M��x��"O�ɛ�V�q�B;B�\]kV"O��A��ӞK�x��J��E���C"OLͻqJD�:��$��QM��2"O���GY=M@�7I�9,�"O�]鶩�
SXĄ�R0m��< P"O�0b0mS	8��ّ���5]��"O��9S�ԝj��<��-��b2ޝ�&"OʸXdI!x�B;��VDƒ "O@�*2��yT舙r�\�����"O�ja�[3V�В�FD�}X-�"OjH�!j�=��9����(l�ј "O�2��gv:�R��6�M,y�!�D8<��`�*]U���@u+C~�!��P.Q� �0m!1C%I��K�!��,v����b_5\�0d��+!�n�sNN�3�U�!!
��y�"O�I8�����81�T�2�>ې"Oj-�Ė3>�0�٦��3޸Q�"OH�4��j�>4J d
,�4Yb�"O�ٱ��*>D����4}z;�"O���� 3�$���,L�/a�͸u"O�R&�	�nٞ��%Qt`<�J"O���n݅p��% *�Hs�H{�"O���"�T�E���H�
ƀ��"O"�p�ϱY�h��扐�6�zȓ"OBDPB%�;��8�)��"ՔZ�"O���QꚲUf������.f˶�RR"O�0�CK "X�"(�&'�q��"O���&�ӻb�:ax�ΉA�L��"OЁRĆ[o��
�֧� ��"Op��T�R��8ZfOˆT�Xx�4"O6]z'�B�x.]WE�5p�v�b�"O�|!���%!N���!���� "O� Ԥ�h;d�	 V��b���X""O���⃙�7�4˔#ĝM����"O��x���]��� A�> �.�Z4"O�lK�E�?]��$+a
�*м�(C"O8@[âʑE���0тQ�i���C"O����[@�q�P��x�Ԝ��"O�C�i�
���֞�ځk�"Otq�戆�8-D9��B�<ޭ�P"O��YUh��Ύ8�e!ݝ<���R"O�e��DMj(p���>*�H*"O��Q�@RBx���o�l�Ҽ#q"O����K-y�5�S���/��4��"O�pr&N�X�0xԯ70��|��"Or� -�D i�������"O�ر�ѷ^�����8C��p�"O�G���]b9`�OU>0P��"Ot��ƃ߫R�Z r$�ƭkݶ��f"O�pY�� sځZ�)]�!n�=c4"ON-+��8Xd�lA�H؏z�h�"O���f+Ģ���)�y�ػd"O*];`��]�"�X�I@�i��=c�"O�1f�]�6��K�b�]�U"O�Z�5'묨�Ce�S��xQ�"O4���U?�Je�A�D�?b\��"Ovd�e ��tr��4`�3 5�8S�"O�a�g�TS�l��.K "r�	V"OfA����I�h(�+I)'����"Oj�Z$�Ү`�ɲ�
�M
``a4"O&�3GD�4i��)%��e�.ᚣ"Oz�#5_�>�͓���	��t��"O�,��*ܰG�$�4
�(�.!��"O �W"���P�	�	�@89j"Oh]`!�}����R�[/e+���"ObX���J�bb��DcO�sH��"O&$�������(^ ��2b"O>5CR)�Zn���UO�? ��hc"O\��@�R�0�MRPNTV��L�"OxݸVf��R���s�N�0q���ZC"O68Bh�>c����$�A	�@1��"OAu�}KY
��KÇAb�: "O�8���Gf�����Ǔ$�p��%"O"��w�,�~A�Q�͂\�T"OrM��	8w�}I�f���`t"Ot���u��i�%�tɖ��"O����
�0����CD�w$h�"Ot3���Ip���9e~�I"O�L�F۰~Uڍc�5-a����"O�m����Rf���&��?KgT�҇"O|��!�0CD��RB��+8@���""O��i�q�h}{C�%L0�0�"O^ñJ��c{( At L�P�]"�"OLqj�'�6,�n�Ccj0|����"O\��w�T-�2��f�?o��#"O����뎘L�^|���I��2&"O��Pg&E��)�c�-є4 "O�p9Ph؍W���-+���2"O^���)�2/S~���&�""O@58���[�$a0�ӱ\�uY�"O
e:��f�����'h͐t�T"O�Y�P�U\�}�B��N����1"O��AqEځer�ScJK�lƔMSp"O6�b&�`*���Ӧ?X�@A3"Ox���؏ �()T*�%W^���"O$U:�� k��	0�@2��՛�"O� �БŠ�?u�*����!k>���"Ov��'%E8$�A�&M�n���"O�a*�mZ#?9�lS-Ƹ[ʒ\S"Od� �H�E�룉��_�5c "O�]; ��F��@VIP����"O8)�A��4�ܒ����	��1�"O��C��"2J��(Q63��Ḕ"O���-�.{tB�X����,���"O��Ѓ�lh(����8I�\�"O�yaN�8|�����S�x˸hT"O�S����lܘ�8udЗ3+��D"O�DG�)!B��2a�0Z"�4�f"O(���	ދZ�l0aV����)�"O��Y�60�"��&9�\Ԉ�"O��a�cрm֪|��f(��@AF"OT18�.�*v�H#�((^4	+�"OF����m��|!P�@�K�`x��"O�3����2�,�h��L���R�"Oji�n��� <�N�;s|h�"O�u����l J �۬r\��C"O�ݢ�A��qsa�z�"�B"O8�C�lpN�A-� N�@��"O�s�/��8BԳEa��dk^�j�"Ob *@8VP �rc:�� "O"$�wc0����J%�f��"OX�r˖ j�xY �L aRb"O~	�C!S�����nZ)[�x��"Oƙ2�	@�KE�v�Ҁ30(�y��c��/eF�Q˴�P��y��ֵ[3^�@�+�\%��AW����y"�ƶ{�m���ļY:prv�Ò�y� T��$��J�'���aN��y�O�6�.�2�H�"d�DI���y��ܗ\%xeC��N�Q*��9T��
�y"-̨QM�u[�x�Z�`sO;�yr퓢*(��3�ں#F|�A�+��y�'%+�0ɪ⧅� ��	Ǌ�yr(G64 �I���B%�5
"���y���n����
D�J�@��р�y"���*��V'���g�#�yR���kH:A�IH�K�����M!�y ]1(@�͠Ӣ�3�|L�6E�#�y�B��%>/X�h#�\�y�/�Y50e��δ$@:|�N��y"�T�V���sڼPLhF���y�R�y!&�%\؝p�K��y�ُ:�f,��-�Q9@�7�y��N�]��%�k\�v�U0a�.�y��V�N �	�u����0J.�yrcD�g�*�zX+D� �2��ȓ0�ݒP"ޙ/̾���cL_"��ȓq��1�GU3x�Vႄ����$I��4l�	�hPzH�T�$W"r��I�(e��-��\��^�J��ȓ06�a�ȅUJ�sၐ"~��ȓ8X�	J1���t�T ��� %��OE����dpiB�N2t��ȓ +�lY�J�Y69��kH��x�ȓxf.��� �U��ixu�_�	�V��ȓW���R+A�4�b`(@��0���ȓ���
�~�8M �L�v�&��ȓ�@ܱ0�.(
L���ȜU��q�ȓ�$�ZI_�	���A�v�V�ȓ,�B�æ׳h��ĨdWtR0��S�? �H&/�<56�ذ��5���a"O�,҅G��y���V�e`c"O��R���	���	�mƨ9��Tz�"O%������D�b� x�1"O̼���ղc�t��m�6 �$}H�"Oތ*�#ߔp���4*��*��]9�"Ov� F�1=�@,P�N���c�"O^z��
q,�������d�r"O�����1��]S�R�*��xs1"O:��R��J���P�	Jl+0"O:iɔd̐��`��K�v�rQz"O����@�"y�U�v�@~��h��"O`�H�Q�{W�5��Bå=�fU��"O�*�FA7��(��KӮl�"O~��r*�7_.�PrBA�_��	d"O�`�D��=*��y�@��b���U"O�\@��<���h��15"OL�4(��\�B �t��I�hr"O��+�'	W��I��M�#��(�Q"O���Β�m����R�^u��8��"O(q�pf�G�R�	&L���t��"O��y���41�T�%^�*�|tQ"O*#!F4h �҂��9��0�'"OB�STg@����`�͎�"O�mk삎
q�5B�kC)��H"!"O��C�Hm,��q3j�BӨy��"O������9��L� ��@!t"OXY���77���h�i8��E��"O�=[p���z���rƉŗ7���("O��Z�.�e.�Pe�%V�ɘ7"O�1�!�շ>����I���%�"Ob�8���n!`���-��y��zE"O01���4
ۦ���솖���"O8�sN̺Mn$1�PAJ�X|��34"Ohs m�#�8j��;],��A"O`p��C'�h�Wl� W�d��"OJ����n ��U�մ9�b�� "O���Ќ<6hv��,]��s"O�U���+q+� ��ߎQ3Ƶ)"O*�p!
��ue �����B$�$�5"O���U3.d�����o�<�"OFicB�]�`��f��E^�H�"O]���&��q�@[�v���%"O���G��b��D��MϐoY T!�"O�	��O���6�3qBz(��"OR`�ϑ�\�`1p���=�`�C2"OR��RKѐ@��'M�VY,��"O"X2����X-+��E���E#`"O"T�����v�hU�X�����w"O�$ cJ��vQ�T���S:>� Dp"O�ظ��H?L�X��N����Xf"O �P��#�(E��㘁#1��7"O��T��:8�#��,�T�a��(D����ML�	�x�&̃7P�r"k:D������$�T�r	�7�}3ƈ6D����.m7<�#��}���Յ"D���eƆ"+|u�	W\��z6?D� C�KX8��9��/T(�F�
�*>D�\���Եp�TDzb���)��<D�8i���6Q�$ap��uj 8�e�:D��*��rp^�Q���(���7D��8 �2iX8 �&�e\�1�):D�$�s�U�) ҍ�j�)���i<D��	��[�v���Y�����:D�� VRBJ<NqIe��/[�x9��"O�� �U��[�n�0>�`F%D�dr�'�]�P���g�)S��Ć"D����J�X�p���>dv�kB�?D� "@ʔ:���AX,���a=D�l�$���9R�,B>����!D�@��F�JqY+u�,R!��QD� D�P
��A�~>20�R.�5�����?D��TmŪ)N�Q����g�|@���=D��!W�(}r`�K
:Ոh���0D��c�����FA��n	����k2D���妇�r(����E,�����/D��)樚��F|1*4kӀi2�e-D���6��@>j���։q�>�a'�?D�l��ѩV&fЋ��R�/��|H��<D�����J�ek�q��Ț4ČY�>D������f[6<�3�ֈ�g�'D���2�ʵ�S 5Q����;D���EI=i��(���<�ڜ���:D�\xV�(;H� ���7[�L9t�"D�(����,H֑��E�n��%.D�,�ԭ���U��Q+aZ���,D��J �^_���bN��vyrsA=D�̋�$�?��`�� �|\����;D��8�/W�&9�m�+�K1�@�&:D�8���,����F�,d�lP��8D��Y�Ȏ06��9�!�/q�R�7D��1ĥՑ��ģ���/yn�$ D�P��M@�Q��j1 VT�`�>D�������J��h��H'�n9�@7D��� G� &��:G%��e2T:�6D�DIq+؁ ��[Ƈ'L�8���  D��� f֤�aP��D�;}2]�D;D�(��J�����P��ji5i5;D��"�Ñ1��\��_� 
J����&D���4aM-�*̣���Av����8D��R󤙍^A��3fL_�a�Z����*D�HJ1A�,tKj�#��o�P�b� 'D���S�d�2p���p�rCO$D�L��U?E{�@3POT"=��`&E"D��8���k�!T'e� ��#D��`�H�? �8�8�͑%|k��Z��.D���T.Q�{�q�0��?�}Z��!D�$x� Β@������Wt�M���;D�гR��c5F��ʊ|��$;D�����1l�4 rn	2vA['#;D��8�*��G��t�`
�[aq"��8D��"���e"~�`b"D$~F
M�C�4D��I�gF�H��x��EP�� ��i1D�h��/O�rK2��K�*�p8)�.D�$�E��.)����F|�p�ȶ�2D���V��i��.�n��0D���i��@��LI���P�+g�)D��JF��?� �
�P-C��&D�x:q��h�Nt���R�.�Z��9D���`��
jĉ���2.f�g�%D��S�#dا�T�&���CP�%D� � �U.i��"�g��=v����F0D���öi��X3���+K�x�D9D��i�#Z�N�θȷMَ"���O2D��;p�� }~�"b��� ���Ņ1D���3�^3��)VoR3����R�/D�@����	hڀ�a��}X�<�uG*D�`!�Բt�����m�2T0n܀�H&D�� ���8?.	bd��9=U"OR4��k ap�Ɽ��`����7"O���G��UE���$Z9i��Y�"O���F��f�)���t����"O20��ęG4���b)�?�y��#)`h�Ң��B��b�j���yb$Z%2��b��@��>�t���y�?l9��$�	@ԥ���Υ�y�@"Hv�)J�j���a5bՔ�yb!۾N��q����S6t1�I
�yH!B�ԡQ�M������I��yr�0�����@[L%#j
�'����L֥+���Aa�Y�t�p��	�'	
P��#ʪ5'*E��,��9�0���':||9��@�¼�G�]]�|�#�'���P$�q%v=;�D��O�X��'J���F��5:�I�s��p1�i��'y�s�J����E�PVQ�'^^�H'�3T����G��^G��0�'8�!��<&'��� \��k�'r0�+�g\�S@���F�C �8�S�'lJ����CQ��C@T�\��'z�Xy��F^SL��է\=s��uk�'b�� �=B��0���
o�J$Q�'��"��I&6\�+0���d��a�'�*�`2̞[-���v�ϗ����'F�*c+׻��$�&&�oy��(�'�d{����:�3<~�ؑCD��y2�ַr��]�D�	4t�Z��ئ�y�I�Q��@�䜘}V�l83i��yB"!3~��ӕ�߹_���:�D^�yR�1e��� KY$VY:Ug�W��y�I_1'%)K �K e�������y	�\�eiSa�6�����(�yb��a��(�!G��@���ǩ�y2��:�zMj��S{Q��R򪍜�y2�ׇ5���祈�x���2�X �y�a\�5����hG�s������ńȓtЬ=#Dܳ!��)��a��wjȨ���A;$�ϭo�8���ʡQe�� #�$�#K��2"�@�L{�q"O����.� U
��!���8�}��"O�ظӣkw
�iȧ�r���"O��Q�ϊ�C�	q5E�9t.N���"O�բm 
=�zhp������:�"O���N��5U��zP�H�4�j���"O�M�u�+�vKa�\-�|���"O4jG&ƊbX����K�}�I��"O�ܹ��;2O^�� g�5/�8@�"O:y7��	I��):��#pd`�"O|8���FM��a��-�q�g"O,�@��ܒ��|�6A��@�(�"O6$���$3!th�a���0	ܔb"O��3"M+4[�9i�g 3 �Ւ�"O�3���W�$�a�f�P�d9�c"O��d�=E^����%O�c��$�"O����H�7!!)���A��X�2�"O����E��7�K8X��"OF�Q�C���:�B#"O�IW/�%� 	���3`̬AP"OZ`+�Zk"��&l߅T�`�"Ofh��@ZP�*@ޑoS��J0"O�C�a�&��s���-Pĩr"O>��֨�7m��k��NCX�B"O� l��C�nk�,�)k����"O� k�i�OO�ȲQ�(�x5��'YFx
���	@��+T�^�_�D�p�'�dC4 �E�j\�B��n�P���'��k�OԴU��w,�cv�#�'E��פ�OSh��ɀ�[	�'j���C�D&J�n�+�޵��'z^�S1��-&(}��ȁFLt��'Ѣ��� V�&�z4cĽ�ʡ��^�<$DE�R!r�0g�L,$���k�@�<)�l� q������#W�Ux�<�b��"�$(0��0N>i�bXp�<�Ų�� �G�)L%8��ƚx߀C�ɅD��%��Nљk�8ᡐJE�je�B�3�����#^U�4ҧ&^�B��B��5 �j4#����� �p��B�I-;��Y�WA�e��ha��يe��B��-a� �4�ۨik�:/���1�*D�T��ʁ.;���J��,g
N��E=D�Dh�On	�ِ&G��v��A"':D����#r�v����M8��I�p�6D��H��V�h<�g��72�(UH7D�@��m�䠕m{������;E*B�=X�Aq�R�D�"��Q��P�HB䉌1����D�$��̺��NM�,B�	+�R��E#�9XAٖ,P0*nB�I�!���@����L6u��C�	"w����r#�'Zdȕ�eE���C䉿5րm�4D�!.V��7-R��C�I�-GTu)���y�q��]U	�B�ɔO��cR�(|�8�V[�x�RB�ɣ*"���W�Z�-��]3N�|B�I�+9.t��jT�Q��u@���&}�xB�I*&�hS�GV�I@�j�4�"C�IJ��͐���g܄���
�-`C䉄l���´oɀK����2`C�	'd����gݔlz0��[%-��B�	�qȶ��p�yp� X��W���B�	7Cs�Pڂƈ��(9���+8C�Ir0:d0�ʜ�+��D�����W��B䉊A��Ā�"=���a]�Mh"C�I�ror{0R�"� ���%�B�I�T��:�
��5��ei�G&B��B��k�������5x���%�3ԲB䉒y���I1"�� � ���E�--��C�ɛ#�!��-͵^y��y'$_;�C��:J<��A�G�=y��PBN�g�:C�I��< � �8t��]�錐H� C�I�b$���Ãͻ�z-�עM{;�B�	%u�� :�i j%4!2��k}�B�	?J.����j��P��9w��B�ɔ!.* ��
1= �E��*�t(�B�Ʉ_�Z P�f�&b޸	�W�u>B䉢t���av!�>[��9�R��6T4B��4o��S�	�^?��U�A�B��2rF`��m�(�d	��R#Jw&B�	�?
u�u�gŚ�ud���*O왪ei�L����"׃w�z<	�"O�!�%�c�T�Fa�40��4�"Oj�і)	̔,7!�6&��jw"O��t�`9ʀ��	�9��4"O��2��((x�
e�^�'$��*!"O��̈e}!�d㉷+B�Z�"O^詁	J!hx�!F�Tz�C�"O� (%�d��Hy�/�!p�[�"O�m� ��a����� aR"O���V=����F<�2�XG"O�@��ݘ>]��cW�E}L��"O�ub�F"D��X�gf�2Pn�X�"OZ�yWl	(g'�)h�RC{
��1"Of|{�@P9Y���s5	��P�"O�E�&-��&=4����ht:�"OXMj��Y�|������E�b(��"O� ��/� <��0UǮM���c"O��A2� �C�-bϙά(:R"O��aJ'R����0�u�X��W"O ]x"��pۢA��I�A]\�!�"O�T	uAP)r�rt���"���B"O���3j�2�ȭ�3#E�L01��"O>\i�df�x��Z�`j�10"O�ѱ6��<�|*�d2���J�"OT�3�MW|0r��đnȰ�{�"O6)��!Z��;�`R ��踶"O42F��
-J�3�@DMXla�"O�� ���W$B�B�~}�"OHD*K�+!������1x���Ѷ"O0� ��!�y��Ҽ�|-��"O�XᗃH�b0�m` EY~�(�"OdQ�`�DV��2%$$*�n0ٱ"O�M���D=`��%��m�{h����"O��̲҄"�+N�3�r|yb%GX�<1҅�a��"��-;I^��f��z@�X./N�82 �Y�z�8Єȓs��}� ◽�n�z�@�ae�|��1��	�˒7H-`���A	3h+����M_L�+�Q�:�Zp&�R_�х�P�0�$�߼+p��y�g�^����&�§�Q`ׂ5��ύ-�r���(�����lI�t�(SP��(z��ȓNg��+d'W49�h5�V�ۢO+t�ȓ(0iQ�*TIB�*���2?Ɣ�ȓyU6U�r	7�H��#i�d@A��wPl�H�,V�4�a/ج[9���dT�g�ʘXst�ō�U`|8��U�0	��A\�*B�c�	#��̆�rj��S�h\1����:S�p��ȓ*).m���ӆL��zb�ĝT;J���3���FAth��cb��1U.>a�ȓ�ii���.\��Bn�^�\��9u��g
�/?��5b��5�PȆȓ6A�D��O�1B��L*
h���D������	Ua\
�Cќ�lu��5�&��!ک�qӍ�1(`��l#l�:3�³p-~ ��+�m�ȓl�R�`g��JKH��t�Ĕ#�]�ȓ�B��Ce��)(�Y�"S�k쩇�/�1-؂*�8 ���/[�m��N�2��:��HR#�Q�F���4�J�S���/;���&F sf̆�]n�ő5b�����c�dr���ȓETEj�#L	�P�0*�(T����)+�5y��6~�Va��\�`�*���� m�U��$+�����ߥ&��Ԅȓ*��@8w�ژW��$���L�`�ȓ;N2@cb �	P�<��/�$H�ȓ'��0(�L�,����B�r��܆ȓ��)�P���Hm��I��Q�@P���ȓ�jAȇ�5L��qgG�o�\8��S�? �-�t):Q��Cu��qE:�{�"O�*�<���P�!&#�@sD"O��KΘv9fqx�焍:���"O���w���`��}i��Ux:a��"O�j6�ҙ��1X�&[�B[��9�"O!"�
� m��G��!KT�P�"O\!�ѧV�A��m@F�KD�ݳW"O��wHUQ�)���F(G�>BD"O��X1�-.zd�ء�8+����"O�M��jW�"���ޏ
?H@E"O��"�b_	ve A��H��Ԛ���"O~�:�m�*f�1D����5`&"O��(w��o��I� 
e�"���"O�kC┃)m����ЛSz�0aA"Ov�B��H�]g���1I�-����T"O8�R�OΚ�zЍ߿d�n�+T"O�\KrJD�63\ ��ȳ����"O�hp���$�eK��ǀ1Ԁ驅"O�|�	И
l|�HE�Ik�8���"OB�S$��?'����(��A�"O�}{Vj���6�0��"{����7"O^�h���T,�P���ҝr�t�8�"O1���A�59v�������x�6"O|�Pa�����z�J�>�8�h�"O�5[0�
E�Bw��%O�,���"O�0���!T����ѨH�(��pK2"O��8�o@ p;����%Q�Ҝ�
�'�
��󯑠h6�E $B�}f�:�'#R�a�D��{wU8��mR��P�'�j��TA��f��{A�ֵ0��Y �'�x�1��l��b���$0=��[�'I4i�#^0BV�@iD�,�:�A�'���8eJ$
R�4D�x�<q��'v�AP��X�Y�$��s��g�xq@	�'�Xͳc�\0�v	�HަPY�'^V(��a��u�2�+�ϕ$/}����'��X��Rw8�A����ٻ�'�)T�X�y�����!:��:�'����]kN�z�D��J�ј�'�"�ᓨĂLxe����`��'�2y`V�9w˚��%�(J	�'�x���+"wTL����$nO�)�'m���B�߷YK��bbC����{�'$r��p�]6S��I��J��Ď`��'z������-9��Pxr���,u�' �X1DM7Q�� ��)ՙ�n��'���(v��}W�����L�����'��4�����=>1Y!�$0��݃	�'4@�:CDOK}�Cd��S":���'H����V��Y���-LG�(
�'�<�H�'��;ˌ��cb
.�8�	�'��Y�_+^	�TK�@HB��4	�'�dU�FaP�n����3�Q>���p�'hZ�@��dA��s�#e���'�p G�!v�X�#P3]�nhb�'=��[��Ԁy����Ĵ><�'ҩx�ɜ��0a{��G�� 	�'f��h�N�8#���`E��'FUj�'F�I���<l���z��(-�5��'��IZw�!wV�ě�,
&���'�F�&�N�T_����t{�̱
�'�`Q�Î�.r$4q�`OƘp>��
�'���U��v�`���
2�2E*�'�n�ib�I���Y2��e����� ���,�%r��7v�u�%"O(��hV�M��݋��O!�(���*O�x@��#��(�i�]YD���'���!��,j��"0J�S� }��'�`��Rh���H₥\D��)�
�'��(�ãV%I�&�R��A�(�q
�'�"x[r�L{�0�Rr(߮e�x�X
�'0�A"�[
ڈ�ڠ��VV੄�z�n	��Ɵ$SV��� �s����n��8��F�3`�{ ܪ%`��v�>�iׂ��uG���`��2���ȓ{�}Z��G�a��X�B-ϲd����ȓ\�����d�)j�T �!ՇU�l��ȓ4����J�7㰑c��ٺk����g�z�SGK����+sDG�l��ȓE�J�e�	4@���q�D��+K�̅ȓx`��(sNAaW0��Fʝ�xv�<��Ϧ`aP%T!G�P��ǣ�d����<���@�<wF�!��
	<����ȓ����M5���؎� �昆ȓfN�����.wE !��W�Q�Ƅ��W:Q ���,��Mz#�	5x���(R��S'/��Q�dP�@H��Ɇȓz����'_զtx+��C|n���@��qIX�ze��X�"�1����>B|H��n�� �|�fR&;H�ȓ=I(l���6i<��!@�),��@����k�3���E#XSk\��ȓrz}��� ��,���ENQ���l"��Ə��wz��t�X�&����ȓ8�M"�X%F�ҭe�	"\܆ȓ5�D���� t�B��qmI�\��D�ȓ_Ɗ@+�[�<���؛w}���ȓW&�B��P#N`*��6�� �J���YW@t �@L,}`NH�N��-MTM��?z>QZ���(׸P�t����H�ȓȸ���(���ٔ�;N�l��d� a�'X%,�	b��e�̇ȓj��0���)�煟9�z$��Pª��`�?#*�af4ZP��<�eQ��&���xt��t�����Joܼi�)Og��� Hũ_~z���F��(�$�M�Бw���5)��Q�r�h�F�<6�^�Ԭ�(S� �ȓrs�h��E�(e�è̏Es�y��|���9vb��`.�qB�x��T�ȓ-x�h�=�-�1��[fx!�ȓf�vx8�]<�L"�k��+ ,��ȓp��0H��L�P���A��k&4]�ȓJY쓔��,e�D+��w����5�r����o���䤐�:��u��gVܡ�߀fw��HC��i�ȓ	z�4:�lC�'�"0v�A�c����{���q��w_*�C #�N����/lԴCFj\3�09����%�r�ȓ}��2�#H�`|2���o�^ʼ�ȓZ�@�mi�h#Wk�-�r�ȓ46�2��	3�H����9��P�ȓ~�(�C�!�;k%<-��������_��x�V F�	z�ЩP/��K�؅�0��e�d&J�l�^�)�DF$�%�ȓJ�p� �]ys��H�w����ȓl[ֽ���)c� q�"������3T(��̍�;�B��݃;�����S�? ����Ŗ3R6ya�b�Ԕ�"O��S��g�n%�����	ZQ"On����VbSnE"%�I*$��ق`"O|��`�1}��XQ'�D�{�(�Y5"Oֱ�2�O�0x`�ŴD�*�:�"OV��g _ d5����b[8A�bD{�"O��ÁbFFt6����q�J��"O�!��e��:%�^�M~
��d"Ov���C- �����c�-$"OJ��&o^=I���O�B���"OD=a �V�Vl�LA��WmNI�`"O�%�W	��┫տ�"�"Od�!�(Štkv�%�/�My�"O��͗�o
y��#�"JW��zG"O܅!W/�F�4�d��%<Nh��"OP�8� �C�,����;���"O2! 9�XU�a� $m����v"O�����2@�4�ҡm�~ xB"O6m:N��}"�)�w�_2FqZ!�s"O��!Sl��DY��
�F��B"Of�	�@�_�|����:`V�a�"O�=�6�a�*�B3�I�.�6$�1"O�H*���*ɰl[a��>�e5"O�ܚ���2.�(
".�3k`dy"O
�����.�0lS��b��2"O����*Պk�)W�H�Φ�@"O��	QJ�e���&+�B�^A��"OZ]B��\xElb�	�.0��h�'"O�iƣS/4�����h/^|Z�"O��xE�p�Z�*��ۦ(Q�YX�"OZ���N��t��mU'nFTx��"OpA����Fl��D.N����W"O����o۬)��!3g��4���"O�E0&ٰw��t����6�8q��"O��:�MF�	u��ؔ���:L���&"O�P{�T�q�@Z#��]��"O�컃Wt/44+7BP3Ƙ��"O�`s ��b�����XE��'~��vm�2'7�\R`��^{�]j
�'����/�y��Ȗᕩ]��hH�'�|ƫ�a3lxQ&�UI�
�' y���g��9���'S�D�j	�'YHq��k6kp�`�斈|���0�'��!ؓJ���b%/Aμ�C�'�`�R�^�Z@�l�$n��;IҌ�'/x��@�Ҡ@�Zy*ӊJ�4�¥!�'���Zw#%l۴�b�M�2+l8{�'�"(��%X&}Ef�sg��5�@!�'��L��$]�g،	+r��v+b���'U`��V,��_;���Ƌ�j��mR�'¼�)S�ۘL9f�s�D�e��
�'�z�Ba��#]��A�i=4��<��'�� �W�C:I(`@!̒-�H�Z�'��U��"����9q�݇(��(�
�'@u��J"+��y�65�8@�'���rg�ľT�6�x����#�l��'c��z��$@���p�H+fx��'�)tF�R� �1Ь� ^��ʓp4�@b�C�,��d�q�� ���ȓ06�M1�ܼXjQ�Ű�4�ȓ	s�c��nt�fө;p<�ȓ_d$�j���.P�i��νc�PT��L�@�y0���Rz\<:�P��ê#D���IΞk!���P/\��0r�?D�� \8&	�\DI�W�@t̀ڀ"O�!��̖�"a$�Bl�R<�1	�"O�g��0�R1�v �6'z%i�"O@��+�-��,����i�!�"O��(W矟*�85�U� *^:��k�"O.��Ã?W�1؀K��W�F��%"O�yɄ�Q�:J�IU,��.��"O8�)e� l%8y6��q��ܪ"O^dWhҋ4ܚEk��M�8�N��"O 0S�^�*NbQ2%�1yp�&"O\����� e��`���ZrV�(1"O�wo� ~[�yOFG�R���"O�}��K8���!�#��9��"O؃�#�_	����BN0�l�i�"O�}k�% �0��qڴ�O A�Z��"Ol�C6�9qz0�`���7+@�5Pf"O<�#��١I)�lje$rN~��#"O�)��� r�d��X8��"O��÷ з<�T�gJ�X4�ɳ�"O%�pJ^3�1"��վtA|���"Op��E�nX]9g�	�1aftY�"O�x@?=�T�i"�ɵ]N�,��"O��j�(ߠ�d��SkT?8�!��"O�<#a��iU�i�@�_� ��)"O���$O�=f,T�S@�DD��"Oj}3�?SR�٧�DZ0r9)C"O�`ӓN6��F,�"��"O\!#�-�2O��%�b*�9 8`xY�"Oځ��Mغ*�&T`��ѤV.��:�"Op$K�E�%(��,��X�N��}�D"O�4��曲
8��΁�-D��"O����I#�֥���N<;;�Y��"Op��AE��N���#5�ϊ8�tU�A"O�͸0/�'P���yP�M�{��١�"O.�Coޤ1��	�be�Z��"O�(G߀U
Q1���l��)�"OԬ"4�Մ->�R�H�)�:� �"O��*���'C��0x�(�s�ș�"OtݠG&�Y�4P`���-G�x��"O���)\���b4eק2,0r�"O��9ЄI�g�>��=$�"OP�!kЙww|�����K#r��E"OP�k�)�ƐI�1��p
	i�"O�}��%D�l�v�x ���,
�bd"OL�))�Q}q�p]d뤽�'"O�%�4FM%.|i%.�
\vh1�"O4鋶)�r
&H� � �!�L`�"OL��3f����O�p4�|#�"O�X5O܄dZ8�Cݮ(>j�!�"O��6��<��$c�:$^�k�"Oz�R��%�Flr&H�[�X�#"Ot
�iޢ[|x5�7�Ny�4��"O�I�vLQ;v[jIs�ژB����r"Or�,Ul��%�ϋ$� ���y��SK��D2#�TLj0ё��+�yb/ڐc�r��5�ʲ&Ѯ�A�[��y"� �$�� �%���E�Ո�yB,���zy"5�7����Ë�y�èxP%�G��(��1��o��yR	��_��Kcgۇ$`l���
�y���u�J�
�!#/�4��4����yrC�SmpHӕL��"ܒ�33�,�ybFXr��0N�61��p�U��y��H�6VL�����6�B�3�����y
� "��fkʰf���[1�»4����d"OJk1�Զg�X��U�K�<	�E"O�=�fdJ06�|r�E%9�Bh#F"Ov0���K8&Ŧ��eV)4l�v"O�����PA�$@·�	f��}�"O��ڄ�W.@F�� b�#]�	
F"O���1���bѓc�tBla: "O�I!1�@�vެ$`s�N#9?H`*�"OT�* *Pn��I񀒊G��9p"O`4�d�,!�m#��I�e(3"O*l�1��z��=���8	��D(q"Ot1I�AP�B��ѫD@��$Z�"O�Y�AU9'�4Y���[����"O�9�Ѐ9=b>x�"�aT3�"Oؽ� 4\�łA��$}�"OЀ�U
P��H��.��p�4���"O��k����N.�L��͓�qy<� ""O
Y�,� 6�1b�ADk�L�"O(U�E�������g�f����"O�����H�]=.%z��P-gPP��d"O�(Q��G�r�m� ��4�(Փ�"O����ρ/\rE�iG��]�0"O�e �!3�&��	o��is�"O��Y��.Ka �@2�C..�z|��"O�}�`��G� �(A�{}�"O����6۾H��M�^��ݩ�"O�������G�X,M�a��#D���ԎV�j���H5�Q1�B���*?D��q5��lS ��a��Q$)�V�:D�TZdR�@�y���+258�H:D��bD�*��  � Ԑ2�]"Sm7D�p�P�a�����lP�E(�c��'D� H'����UO2;�޼�a&2D�D���\E j�*#E��2��l��/D���Ɗ�'3��DH]�"О��/D�p*7�M>V`�9���=��yU)D���Ήe�Z`���otԲqA)D��'eK�̑���8q4�
(D�j4.O�o2��4�]Q�Ph3�j$D� ���ȋU�Z�PFc!l�fp��"D�x��:6hP��dCG?N�y�Ɓ"D���B.Xnd(�@Z���#D� :s� l�Q��6n-�])ק/D� �6���-�J����_��i�j,D��1�K	�
8�=+$ޯ}7.��)D�\i�F]W(�*��T:� ��&+D�(Q�8�b� �O��̊d?D���Uo�	�>m���J�prAN(D��FB�moҰI�&�eh�9f�%D�)$n���j@"G�9u�Mٶ�"D�����K����,��H	��bp� D���fBM$;�ʼ�ec���8� D��Öו4����#�NDv�	�#D��ك�Ù$��!f�ح�F!Swg#D���F/$<���b&T�$˱L"D��pA�
*���C�>��2+ D�T@Giܪ<-��P�MR�hqz�?D�IK� <ظ
�U�~��)>D�t�q�����B!	K�jdV��S�8D��i�&�1[kJ��'�۟y�`��aD2D��8s���(�vQ���=r���r$.D��S�l��3���b�#�,D�8�Wly�؛k�u��A�Ca(D�h`f��^Jy�"��
Z��:�"(D�� �����d�,t���K C�tZ�"O�m�A)�2V�B��B����s"O*��"�֕p3���w�� �,���"O|��f䈢V��p���n���"OB�����E�¥C����7"O��J�#�.z�bŠ'.�BA��"Oh� �i@�}���9P��5|ޜQ�'��;�8��j�r�$(EjH	]�h��'���?���d�5P�<�v��
?Z�P �g:J!��M�:�z��FO�V�E���wh!�$�+�<��֡_
���:&f���=E��'��i���
S�RxѶ��%s$�X
�'t��JVA$�[֡J)
�r��}"�)��P�G��	��f�|KU����B�!��	�� w�x3������� �=q���$9�*�#��pK a�%��@��
O(6m�Mz�`��
��9vO��I��:pDaxR
�10x
�O&��hx�+���>��5�yr��)ac��{��7h,�%I�E��yGE�x�@�)7�CZ$4���$�hO"�dq���o�'6�p����'d�0��FF+ú��D�	/��m�%�;f�@y:P(��B�)�$8C��Q	+R0CtB��dP?�Ѥ�9�,{�Dʚ$�B���Ŗz�'��x¢ёm�%�jao6XCC��;pO1OX�',v���H�缃�ˋ�#\�5��-�4t���HA��<�����+!�xh�YDљ�D:%��	Ϧ���T?��<�m�������Պ|~�u��Cw�<�2�C/��S�YA�٣F	�q�<���7?nhc����P���	k�<��\�q�=���JR��R���(O��G��O�s�$;3L�ۤńpd�O��J��Mi�$͝.J� HS�ԘY��V�)��U�s�B�dzT@��mȱ^��*��)�O��Oܼ���\�UH�#N,H��"O�  �оl�J!�bBV�oJ)��W�&����'_���ږ��-XV�0C�TΉ�ȓ�n` 5D�k��P�����2���''�t��Ι�8}����B!a|���d�<�!!�
~��)cf@K�>�r|sV���<!�J`h��dF�FR4�G4�l��y�(�;e
Ԟ��1��l_+^۪��`vh c �I�V�L��K�)'||�ܴ�O���'��zdc\��4��a޺B�
�'c�1��J7l��R��y���K�І�I%fo���(\Gu� ��A�`�=Q���?�i ^)Z��Ż1���쵋�/0D���E˺L�KL`��鑤�G�J	a|�|r���ðH�=%<x'Eȼ�0>�K>Y���%�,-J!掛l]�д�Q{X�\��[�\�vJY6w�*0:�+^%D4�GD=�i��#~z`�	\��' P6&�����L�s�<9DJB�j���I6�ٳuq��c# S�HO��'��I��M+��T��Y��	HH�^qHv >`���7�)��<�vfݚɦ��GB�.W�n���ZJ�<��N�$P�+�+�(;���҅�C�<i�@J�F��]��C�.�h��3���<�.O���>�cA�u���X�m�(ׄ��$x�<Q1��y�^\��KJ6������p�<	A!��B)�X��/ao$�#r�nX��Gy�gފ:Ab1C$	߉^z,"FIS���/���j\ғF�/���r�G�78�D��� �r�U��FHî-},�ȓSk0����Oy��hU,;��oZZ?a����	Fԧ� ��PRh"Gܼ�a7N�8�D�h&"OV�;���Ĭ����xr��r"Ox�`�°2�����!A��×[�0E{��)J�&���;�	S�6�PeC��7/�>���>�E�%E�� ��.��n��Iwܓ�hO�O��8�&�m	20�%OW�*8�'�� �!,��_/�`��$}�zقN<��'ߛ֙|���˓�F�$��<���r!DڤK�
݆�z �8H�Fѯ-���TkٛJ�~��.�IL�TE}BDQ&B��� ��,`� 
/M�yb�#%\����ؚ��ɺ�D��n� ���$'�O���J���W��{���);��'��}b��>$��l��Uf�j�SW�	j��C�	��� 2��cT�Y$��S�C�x��Pi��ݚ���f� �&�VB�	?��p-����XH@ @�-N2B䉊#c����9Zv�����l�PB�I�L;�\����C6�)����|v4B�	� KH�)�� ���a��-usB�'x|i��%��j |qt�=Z"B�	�K v�+E�;���b偪1O6B�	iT�u��H�Sk�9S�^0m|B�?�P�p2;�U�@臼R'VC��'O�y06��7Y��y�7���B�FC�I�@�bE�m��oQx����ȩOv"�	��������A��X1̑Bs#K�5�d��"O�Ȫ'�A+d�\�
?1����"O�����L+@��2C��(z.z��Q�x��$Y��O�r4�fȍ����IU�_��Y�'B��)��H?+X���φ�H�<��'CfY��
ֳK�B)�k�?"�i�'�e�ԋ�6<�1�+V�ɥ4D��F��5\���f!W	O͆��% /D� j�7�PyK���.[Z0r�A!D�lW�9�ްSEm�(]Q�Q�=D����A,��4$'�2D�� ;D�h���Mz�0�O��IIƌ�W�n���$�	H�'b���Ц9�B��p�̳'���I<����i�68%�R@(n�|����I7!���,Q�B�i�JE�)��M���)!�D�A�02un�/����&D��P!�P}>.��fIG !"H�Pb�O;!�.':�'l�;,bJ]��.�/]�!�䇂$ŀ�jq!Q,�䤋� h�!���3!n82EI�f���ǳ�!��!e�����&l�S�s�z����p?�S�+�����W
<K�Fo}r��_�,c�"}�U��?0��2�o��Q 	; ��l�<1�-g�c���3������Qe��y|RR>�I�\$8%-� ɖ0��ՋL������<��N��1Z͓RHO	M�¹��%GR̓��=Q@f^-QM����(��@0�r�EL�<��MߔcV�5+O�^��"�DXR}B;O�˓�0<�gJ��]���ѱ�/]�Б� E}�<Y«@�jO�ؙrˈ2[$̩a�.{�<�0Bƿ�zx�d�>��y6z�'?�?a�#A(>j�H���5�\�"��<D�c2K@<vl�ra��g�N!sf.�$=�S�G�ЃNP�0�c@�˟~t��ȓ4}&�1$O(f���*�5m���ȓTc�QA�h�!:�	����B?�|��$B�B�K	?<��APJ��I�����I[?����#aVt��CD�@��B�N]�<9�̻~��}��C�I:^eÐ�IOX����I�S�? t9���.x�z1�ʁf"�[�"O���� �\���='����"O�q�K�
XZ�j�/M�|s%"O���!�n�i���J�q�X�F"OT�r�J��[Д��F
�lq�@�&"O���V)�[��ʋ�����"O��@��I�+*�i�V5^�6c�"O�q�$��#a	��Sŗ,��U�C"OL�i��L�}�Y#.��1���T"O��D#�,��T�_�#Āx��"O��I�*؅*�~�9�. F�VŊU"O�	�G:
�p��焹^��<r"O�A��D�;���3����`�"O��� k��zA�] �i��"OL�kGo�3=4��"n�*lh"O`�R��z� eq�l�=n�� "O��*A�_�m:MA��*�Ѹ�"Ob��b�I�*@T�U@�%W�d�Rg"O�����!6b�������(�{2"O�B���/a���4�K&��}�!"O������0m�ʑ`lR.0��A"O����<:p�	]���;@"Of����^������5E�p�#d"O��;��Ժ1��=�I�*E6Y�u"Op��#�([�:�@�5Y��|p�"O�����K�
�>e0�G� ~��R"O�tcCG7 �0�H/k�Q�"O���@˺2��p�]��*(0�"OF8���[H�i[V"� -�R�y$"OJY���6z��P���r���p4"O��� +@,�0�i��̓�"OVŲΓ�',�/��16�nw!�B�8	FIB�,,��Aל#�!���i�u�� ^����"��5E�!�$żL����ǡ��QɄ��O�!���
|p�\���g����!�@����
��5'�hk"�0x!�D	� �1� ��5r ��r�%�!�D_�G�\� ��Q��!����w!�dǽC�@X��C�/I5{-�02g1O	��I�5hh�C��E6}1�:`��	���F%�q�䤻 ş�)i!�$ڶ ��#
D#@8 D%��S�!�D��7�0Ex$m�|�n9��oU:�!�dKq�\x�������s�nͧF !�U�:%��9q Z����ف�̛!� �Y��8�n_+l�ƽRЌW^!򤜀E��h�V�GA�N�%�OK!�䁥B�9%�â��D�
�R�!�DT9��'G�T��������`z!��^15�r]�N��f�¥Y��Q�k!��'R<T,1�-i�<�yD�ڀn�!�&#e�pP�ͱn?�p/G�!�6|��y�P8�E�f�ٷp!�M<(T� �B+	�>�I3��!���#Xs�$ç{�NEH����
z!�dE	s��5Q�d�*�e��ji!�
8�M��ԉ��۳j@�k!�DD�H�b��GjՐ��1+T(�1CO!�D]0���pG�ߢVRT�JqFA Q!�����Pb�\ @��y��۷ .!�X�5j�)�D˓4F����I	��{r��<:��D�'��ZG$�	��ԛ��Y�= m��.ۭuEv�0`��O��ȓ@�&�R����J�n�� j�>Ihe��h�$zZqO��Y$ҽ,�"XJ�'� U��e�" ��m��Ҳ-�<�ѧ�Q�&���2T�s�|Y�����|�mzB֧�y��l�L�҄�/�ڂr�=���|��i�H�Ѕ�/�ۀq�9���|��n�H�ׁ�*�߇w�?���y��l�2z�>�Ηb*����2��.]ӆ2z�>�Ηb*����2��.]ӆ2z�>�Ηb*����2��.]ӆ2z�Dh���l��yDڦ�NAw�@l���n��{Dޣ�HDs�Bh���k��A٤�OCt�Fk��0w�
w�X�׷�;��f�0w�
w�X�׷�;��f�0w�u�\�߿�3��`�2-���1p\:��;iC���&͖�=zT=�
�<aK���,ǜ�9xT=�
�<aK���.Ş���Z�x;c��_�]��*`Y���Z�x;c��\�X��#jS���_�y9g��W�W��#h\���P��Rl�<�pwG��!��"^��[e�7�wrE��!��"^��Xf�4�usE��!��"^��X���:[��$T�dy�Q��K���2]��&W�`r�]��I�
��0P��._�mp�_��A����o�7�%˾6ޒ��6s�M��n�4� λ3ڑ��6s�M��n�4� λ3ڑ��6s�M��k��ò.-2�����e��#�;��ǵ.(8�����m��)�;��ϻ' ?�����c��#�7��ɺ�,}cY�Ot�r|:�g����#�,}cY�Ot�r|:�g����#�,}bZ�I|�xw6�h����$�(~ԝ"�� ��T�i�f�rz�DNޗ&��*��Z�`�l�|q�OKْ"��+��Z�a�n�u�HCњ*�}��1���[�}�|{�}��1���Y�u�qv�v��6���^
�v�ws�u��<m��A2��(n����ы�;�e�E5��+n����ӏ�>�`�L?��"f����ӏ�>�`�Lm�_az��#�_�h��wu-�b�Sjp��+�X�o��yw,�g�Wgr��(�T�f��yu!�o�ZgM1u-0Z����w v�2� J7s(8Q𸂋~&s�3� J6r*9P𸂋~&s�3� H5w-�P�ʯ��/Z��Ȋuf�ᬵP�ͫ��!Y��ʄyi�כּ]�����,Z��ȇxn�믶R��wD��E��y�m�{h�h)�3�tF��G��z�n�yj�h)�3�tF��F��|�g�rf�a#�8�~O��Q_{��q��F[���53d_Ru�|�s��GU���71`ZUp�}�|��A]���8>hTX|�98M1t����֖<�c��Y98M1t����Ԓ9�i��S24A=����Ӓ9�e��\<=K6�K�b!b�����<���sk�F�n+h�����9���yc�K�`"f���
��;���d�L�e2c����]�"3t�����=9i����P�)9r�����27e����X�'6p�����<5d���%Π�>���X���ϫo�熏!ʤ�?��P���ʨm�〈)¬�7���R���ʨm�る,���.K9�W�I�t�1&���'@3�T�@�}�3)���,M3�T�M�v�>(���	'��Mم�s)&����ߏ����I܂�y#,����	ޏ����I܀�~+&����҂����Cԕۙ�^�Z>� ��������Ց�[�T3�,	��������ג�Z�\;�,	��������ڙ��"6}�z�����D$ň�~E���"6}�z�����L.΅�sN���.:v�s�����E'���wO���(?$����7Xs�E��=Guz&Nɞ)����5Xr�D��8Cvx+Aǖ!����5Zw�@��:@s#K̛,���߅�C�����X�Jv�rЈ�I��˴�\�O|�x׏�N��ʶ�X�Ix�w׍�< 	K��Ah��]
W�����2.B��Hg��]Q�����:$
O��Dm��XS�����8'HjF��FɌ"�d���1R���q`O��C΋%�c���>P���veD��AΎ �k���>R���p`N��&���]���<N����"���W�
��4I����"���T���8B��	��*��Ԫ��R�ցQ�gNu,�c�}.ӭ��X�څP�cK~!�c�p%خ��S�Ҍ]�cIs+�g�r$د�#�<:ۓ�bHrQ����Z���"�<:ۓ�bJvT����P���%�;=ݕ�fKsQ����R���.�63���rV�6�������U���[�;���ʅ����P���qV�<���ς����]���j%bv�'�U�WܕcW��K�?b-jq�"�P�SߖcU��N�2m-k|�-�]�Rِg\��G�:e(n|,�Je_����~�,�Q&����(�MaY����u�)�S%���$�BlU����v�)�S%���$�@o�+jc�2�A�*b��Oϣv�-o`�2�M�&a��J	ɪ~�#ai�8�M�&l��AĪs�-ng�ʥ_@q��M�if�����ͭUK
|��G�nc�����ͭUK
}��C�kf��
���ϯT�<6����v��x�!�EI�x�5<������v�/�OC�}�7<����v��v�+�IG�v�>5�P+x�b�n�T1��pэ��P+x�b�n�T0��sҎ��Q*y�c�o�W5��w֊��U.}�%8CE� +'q�,�e��"9CD�$(~�,�h� �*6KM�&,{�$�b�	�/U0+�5}��q���� P5.{�7|��q���� -]8,y�6x�{���)_9#x�L�W*�'	�� Ω׽_w�A�U*�#��ͨԸY��J�^ �+��ͨԸY��K�]?��>�>x�;���~&V�|R3��3�0v�:���v,]�s\2��3�1y�;���w,\�wP	?��:u��k��PL�C��T५A-�p��a��]A�I��Q㧫A-�p��a��^E�N��Y믬E.�r��`w���
�����#�䃄Z�{���	�����&�烄X�|��������)�Z�q��_�,� �عk�9}L��_�,� ~�ܼl�0wF�
�Z�)�"|�߱a�4pA�
�Z�+��?N���=xJ��[�ú���5F���;}N��R�ͳ���5@���:M��X����
��2�Uէ���r�G<��2 ����^߮���u�E>��<����Y߯���z�L1��= ����Rӣ��~�X��`��!�Y�ʕV|��q�T��`��#�Y�ϓ^u��z�]��e��#�Y�ϓ^u��}��򺉓�,�����ھ�̒������!���Ա�̑�󽍖�"�����ݹ�Ř���&�e�9��E(�C۾�SnT#�m�2��H#�Fؼ�SnT#�m�0��O+�Iհ�_bX/�j�C�L���a4
�� ~�ռ:M�M���f5	���,p�۳7F�D�ʗn:��$x�Ծ4@�D� �@ ��	��-�?�sG�/� �@ ��	��(�7�xJ�%�/�O,����$�5�~L�%�*�M�c8s�����t��%��w`�x�i5|�����y��(��zj�r�d;~�����y��/��qg��n3yA�Uw ��-!gH��wTS�[N�Y}��!-mO��xPU�YL�_|�� .jD��zPT�[M�]p;g쇺��P�������T~�I9d脸��Q�������Qx�@3o䏲��W�������Qx�@1l��h���r`� 0w��)S���O�o���t`�'7v��,^���H�o���uc�#0w��+\���@�b��&�q)��54٭8x1�,�H��"�v!��?>Х?}5�-�H��"�v!��:8ج5v9�'�O��%�s&���F]�04z#��9���1����C[�75y'��?���1����HP�><t)��<���=����G�X��!���p�����vG�X��!���u�����~@�_��$
���}�����{J�S�G��%�"�MK/��Q�B`�@��*�)�G@$��^�Hj�K�� �*�GA&��[�Om�M������t$o�:�SF�{2!1�;�����|,g�2�U@�p;.;�9�����x/e�2�[A�}7"?�;���� ��!M�3�$���cG�ea�TR'^�4ƐCS;>r�RF̥t6�cC��5�4��K<I��"I8pp%Ϝ�m=���`+СR��Pbd�P��e���	�r�`I�#H8�	n:�����"U
���$�A�I�7$��Z-�pΈ�4(�0$[y@T5"��e䈤O��r��&��A�S �|CdJ�0�IQ*C������͆F������6Hz ���
��X0t�@ޟ�aj&��	�Xw�2��V�=��� ��2c��p���jѥO�P�aa�H��cgԔ���#�L�$��� ��9}V0��
����$V�����C��"ɼ���Y/Bf�I`L�>;l�2p,Z
	����Q�V������  ���#�S<U�*|��#�j >**�;�a 2\� ���GI:a���sB�W�Π~B��Q�Ĺ婃�0�+'/�L34H�.��_�$6�p����1��-�ೋR?�y@�N_����mG��i�m[)Mz
@�$�ӌ/z���d��֠��Dg�O),�Вg�m@�ם7l�8�p��H1��GZ�`hD��O�-sS �@U�m�EOU�~��G�@�@$E!�'^���8+9,>CPy�F	�?P���s�3J��� XϬ|��`ѷe\0�T��y�)�e��ke���1M����[ȢX�& �4`N�e(�2�:e1����4��d�I,\����'��  !^�nAt�J�gk��Z��)&$�V�X�H	0a� Jf��B��uj�l�
0��<C�K d���[jߤ"�L�S�ɱf� ��=F��n��R�>����!_�9����B� lC]h����Ս"[��)�,]�F���2�ѧ�ZErR #2� (���5�� A��!�B���Y�Rs�L�ĵ0� �"1�*4�Eiē2��<�'��("�
���RS�!��)�!��}( ѲmXu��?�(�1��FIA' %;���<U�h�𠣕��\���^�H���jƉ=Jq(���6/��I�d �>�a*� xn�M�/�'���j���,K�ii���C��YBU�EH�z�	�<K$�%nR�p,�T�U�� ܮ �3�ã�Ms��ĜM�lу2$����'��=+��u�0ޏ��C�Z�\a�l�e�h� U�UZћ��	C�d�9A��a`6��7��1�4,�a�V.��y�f}�R�� �p�y1���``2������E�(4�r��Ab��i�46J����ߒ#�vy�� �N][s�Y���b�]�<�o<�B��oj�1c�@=�e�f-0sB�����3=P�]g.��O~4�pӽEp��I�
_4b=�f���>��'�G��I3���؏@�AgDB�K��3c�C�M"<�b�N�h:�0�n�1B8(��.Q�0��J~"@	&Y��Y����ةm�����G��F&9R�$),��#=��m�x�jq�#�M��9x"	T|�jI��Z�?�rY�FHA�d�4�4L�l¬�&�l��N,܎Mc�gn�O(X]�@�o�Z� �ڶ45��р��%!ҍ�F�D
ER�I#�H*^Q�`���X��kLC> ��{��$G�a;�	I-T.XX�3�J�f~b�'�X����ɶ�ا%�V�x�'�|���?����8!��P0װ,�H�� �8o;8���B�������>	��=yぐ�V�Q�v�	w���3ҍ���\aeA��jf���xC�E��Fá*��$�v�����72i�aȗ-QK��#��(o�4ekrχ3�j�Rń����>A"E��}}�q)'Aפ뢨�'U�D��g7�bZ�-�n�yRE
�
pI����%EЮ�(�ۼ�0iJ�5���W�Ĩ-�|���h<��^�/����F�%�NI�a圦h��͂��lw4�bU�^�q��K�.,�����璛'�J��\�j���D�L��F��ţ G����<)�-͏S72-��!���ܕ@���4ev�R�LM9KH|�A�`�D�X\+1�G�A�����R��d�D4`x�=	��FFX d��O�X�����|�;$� �2���|+` i��
�*�kb�)2��ۇb��0�uz����+*"!A��I	-X�I`���c� X���'A�<�F��Z89����*@$܂���n���	�ӒY�|����kL��Ə�R(�M&*E*�ҞwBf��s�A��3 -~�K3$@�9��|2M�+�o�?�����'�1��`��� �o	�{~�- �LϥL���a��r�����7��@����8�'ɼ�8�� :v$	�v��)P���"b�*��u1Qn�u�8TRXح)�B����ei��"i�(��@֙P�Xh��8Ī�A��O�k~�QE�� z5��&n� Fz2�E``�J��S v�h i6I�f]yT��|z<(U���@U۔˗Fgp�Q��W)b�0�	ԴL�b]qT���R�2M��GF�JGЭsѦS#3f�u�j`���I���Xj�A�'��XBa)�z��7��&@�A"q�щ!�@��z��Tj�aݧ�� �)�j���O$)<��*��ØKu�Ts�*(�X�����2�R�J�������#�i�A����S	�Sr���-:8��� �
*?���� ��x�:�ӃiB����㩏�Xf�g�p=��j0�H��#M�R�Db��Q���V�P�PG�/�4�����6��j>,z*Me�ã
#dNuj�b#5��P���Ѥ;;� ���%  ��N�J���l���x�����IK�d�gă=Z�<3!�F/��4���K7��d^UFU9��ȕi�|؇��|�|��a��>�X2��X�l�`��h�=-(�/��PFBہ;��9n�0��a��oz��bEB
0c�~$'���jd��� 6�BR?����9Y�Vd)&,�e::|�2a)�ڹ�a�O�f&����O�'9��ީ�ޱ�Q
��b>��Rc/�r�ײ=���h�n��L��� ��҇r�j������[�i���X���/dy��Q�ܿQ�i���kLYN��tؤ�"�H��͘�	�vp�4�O�
� 2�Oh߂y� ��HˤT��kP�?A%��(b@,��y� ��"-�$�3G�� �JA�Ǭ�b�̀:~��h�.��#<AfIN�n���H�l`�4�oF`��L��JN����VF
)��'����&�ʓ*�|����}�4\h#(�;��t�6��y�����0����w�W�']��1�Da%�1�С��G�`�z��B4`��d�O�d�`D�x"	<�2h�S���a�3�X졡������r, �!�l����$$<�	Z��-�I�x�x9+K�u����4���اh@4��ph��Y�h���+�>~	���2L�6/�0Ԁ�*:~���׀�=(��A�"�Y�l�����<z���R�6�yE�����Ң�Q�vm,8q'i^U�(�g/ج( m9G�r���q�}�����O���dO��T[�!^�He�P��L�����2E/B6p��TFH��š�H�+V�2DC��IgQ�� ���7`�=/zN��l���b��;}vћB煚>�p}��N<'����W�x2C��{GHQa�oA�s���Ci�=���c(�Fj<��'ٸ9��}���/%�8Z "�~�!vB>���h�k����`E�M,ՁC*	�d��z�P(���U��jX#^�����8���k҈@�� ��a�M�,��}"�Ҧ�At��@	\�����mP�@"'��|"%��kx3 �7K&L� #�ݟP ��@5
rU�4"��3��ʟ��F������^R>�۱D[�Z�����#N{�Dڥł;G���E+�n6�̰$�M$_P���ͻ1��q�
�-Wj�",����i	�!m��B%,q�<eI�\V���D
,q.m@��\-O���	��.���R�Rg�������F1.<���̙��9}b�ɔ
wZp�!	�!�\QB�ᅬ0=#���Z����'fJ6'�:	���~�|�K��-��KS�L9 ٬x���9Gt�CI<�TO�r�,䂧�%����`Vf�#��<�$L�\⟌����
-'�q�A��tO@�9R���
��N�q�#߭��`��'�;�0�|�>\
��*�)�'+&D!�����;��(4&�"��!�B"�)"�sAʉAd�L���*'�>�][U�Y��QN�N���nT��C�I�b!L�pu׻%_�I�K�;cvP	&�ԈW%t�C�%�F�n�f��?�=�$�ٜ	�
4�喝+n�Г&��Mx�ԛ�IJ�����*Z-uz9�����Tp/_���JG��c��X���A!)�赻b�C�!� ����;�����Ǯ
�T��z$qEC�|R�Y�p	#"�"�"OX���d-[/L��C�&D:-� "O8%��"��
�yAĎ*v0��
�"O&a:�$I0]8�cC 
%*m�C"Oq�-��%�$�>8)2"O,��Q'�.c���6��
{�l��"Oʈ�u�.i��}��@7H��t�"O"M���vFQ�u�Y�?��y	R"O��p��R���S&�%�V%��"Ot�d.τ�&�xs�۟K�����"OH����u�\u�Sc�<�Rd"O�`���Z�ܘc� 	p�"O�ٙD��EF Aㆇ�_�dݺ"O  �aC�T/��v%U,��z�"O��pkɫT��yDA#"i�Ԃ4"O�|��i�/pL�L�4R�_JI �"O�4���Og�v�+�y�h[T"O@Й���7�,Pх��.nH-�f"ON��@(��$��D�f�ؓ9S�XS#"OxؐŎ�ZJ�AP��5gX|��c"Ox��a��MZy�u�P�U��hr"O:�ғ(�L󬑰�N�8Q��Aك"Ob��2D�#T`ځ�Cb_?{>{w"O&=hf+?���T�&4x�"O*<r�K�
J �u����G@�r!"O�E�ްޜ���À�Ľp�"O��+c�W����1Q.�@ĐD!v"O4��#t�I�N�=;J�;%"OR|��׷-*�eC�kǤ����"O4�����i��jB�^�b�.�yR���a��I,5�ؚƆĴ�y�B���BfY�̰����"�yb��<&�i�FԐ
�ސK5KE6�y�(=b��&�E4?�yEE
��yҋM6]߰��J0[��,�4�1�yr`D�cj�����Rh�����yB�^�LP��)ن,reR�e�7�y��^V����̊~���s*��yr�P�t������)�F�떌8�y"�q��$����V�� &���y���N��H"��>F'ެ��IU�y��TR�m:BH�<:lTi��)��ybʶ��1��)�����y�Jʳ+.�c�o/����N��y�&&*�����	TM�0!�4�yR��m7@p*'�9q���j0Mؿ�y
�  ��2i
�b=dY�r/�3\�j���'��0�ō�p}"z��Eŷv��#fA�w�tաg!N�|PV���?`�j����Oj$IЁT�`�������-4
����Ė�txfc��~2��"O��0P�C�Kx(�b�?3��L�`���<��+#+��+éO� a}�!�.�h���J/34��M�9L��
�֙:�R��.s�Z�˔�.�`����C�11�2�M9�y�"�;xxf��fa4��ex�
���xT�Q����CJ�0y^�e�-ִ,�H��k�>��	���2�h]���T�R����3��1{]�a�m�.�D�;���B�葊��0"��2R˘�s�aykcBH�s䤗���=�C��2ax���po�
rR�r��id sf�O��b��@�����a�2b|���o&�ăd��੕DN�P�%��E�o�]�D|�$sۤ1�D��}����0CJ�eY:�hg�[�NԄ��'+Ȟ	�tY��ʙQ�1x���O��9�WHV�\h��A5(Q�v��	!X�t���fU�EqO@�p�#�;>4�l��mG�W�dᚅNUq7���##
�|�"���[�T�0�#�9;?�@�P�/S�x��%.���św`H�W����AD>������'�XZ%@	�kL��@�'�����28L��sd��7~��u�Ā�� <��DZ8B�u����L�LKñ<E��Ԡݵ|��i��ϗ�2óN�:�,P���_�i���6g�u�џt�ڀz��=��$۟doڽ�g�ΑuW�ܨ�e7�m!f�h��5	7ʌUjIA \f���ن��rW���A�'�Mq�i٘n��	a�E��Db�J3Q�v����2��@c.�W�N��5K�|��hj6h�[j�-B�N�\T����h$g��8!�B8l��4A�Ⱥ��iB��(�;��۟�m�71'B*�q`�BC3�(�A�!9�;&�V
���,U�R��Hؚ:���+���b�Z�0~�����HQ9"�F9ZP.P�N4�wH�>��K�U�~���Di�57����AG�5sV�)��O�`m+㋘qBU��}������$U����YCM�Y��� W
߫^w���BF	5c� �]0�p��ީZ�ȐB�H�3n��U+���M+e��V�$1s�M�x2�iJWFZ�4t�$r��L4V]���'���-�PsGɢ�ēL��\31�O�C�
�ɶj���9C]0��ј=�r�WQcĊ¨^��Y��(J�lt�44G� �ҵ+ޕ�����ˇ�KZe
�[��1��Fħl"�Ҷ��V��T�7� ?!��ÊW�|�POÃ%�܄�M�Cٛ�J,&�Y�d��(�h>��=�	��.�P�n�1)�����h�	��3a���"�	;���0�ܰ�0�(6.
�,�q��
��x�M�g�Q*�����%[��]#�7O�� i�L�i�5}�@� E�.p��b�-F�j����Ę]��Qz&(Sr�Q�:4BX1P,�6a1��B2$D���#�͌qc �0?i'��0&x�seJ)�^��4��*I�P�Q�F�R���rHL�ڡ��-�1+x�C��(�@���͜(L�@�	�BF>V]�aYPWE�f��7C��h	Bq��]�bM TM׿6��.O��E�7[�����EX��:Y��e0���p颤�Q'�j�f�Å	���diW�	z���F�8]��uP
OצMQ�Î6U۪�bw�"��P�2
=`8!"$�.���'�:H�a�I2�4
K��!V�ӓ#G���X-'���`���4��7�/A5j��Ǐ�
7vi��`��~`�2d�ֹ}�h�83�V<��G@ƮB3`���/�5z)�^lZ��6,G5:���Y�8&xyؕƅ؟\+�P�<��	�b׆XgN��fLG�<%�i� :"K�cny�w�%��i9��_����Bv���{H�Yr��X���%��.bjm�'Z����#����_P�a�J^0Hh��*�5�v���e˩���٥�ŴI�(T#�W�yV��:�ʛY2Jp��B4 �~Ͳ��(y�6�f�Y�t#\�p$
�R6 Բ��S�eL�q!��	C��;-O�=	��݉W,�:$�������|9f	y��BII p�đ;��	��#p�$И��P��H �3
_�=dY�iC�H
Q`�<���C�3P4t�����X#����Ͻ
�˓�j�`d�O5:�8Lb��T���IQ9���� �P1U
�Y�rD�t��!B8Ԕl�1ǝ�,N>���@%-2�C-Iv�i��$��
\�R��=ބp����)D��xb�ЈIe�yR��W��0�z���#Q��t�Ov�x��Ԙ>�T��(��6�6=P��S�^�����.k�`gʚ�c�tm�'���Aڼ�1�&� t��)Z��{�̡�-�fc�0(Ǫ� f�fM�O��q`N`9n���D��!pl<�T  ]��X(��F�F<�Kb�Kb����e3z��Aē�${z�f��Y��X փ�#pp �+U��*`R\9���!B�g�9T���r��2A�'��a�EL�(`�p���OXdؕgϸvt�� #�;Q��Xp�;�GP>l�0�:�@H��Go!&g
>h� N��Rl��G*!�$�ie%Z1�yZt��>v��'�qBD�_��5�Z�@;�@>L���㗎яVG8��q��5T�̄#D� 1�a��FXC�n�;Ek�h�@�����nE6P�بK�F�
4 ��э�\8��)�Bd1�lA4��10�Aʒx�:�9��O���g�:_����!���	�[=x�
����H?I�"�+3/�<f�"�53t�ĭ ǭC�0�b�C�C2_�=KG�\t�.�k�o>`�6(�M<y�&9 m��G���h�@��!��2l|�cfX�~��=�� )�U`#fF��MSįt�]C� ���"�qÃ܁4�"�� �J'̍�C��*�1�f�B�*�@�a�]=�B�aI<�$C�:7r���C��3$�HXX�a�;'�ʙJ䧐� �!�#E�V�3�ܩE}�cR�Z31=��C
rLT�c�"|L�i��ƈf;��I��U�y���f�޵w�.,+r��d��'��Mp&�S9 8�rC/��>�dݫ�n�aO8�;��T��ՙ,��Q�aȃa�B!���*\�B��2�؆l�(8fi��f�Љ�5��)��u���b�H9��ܫ^�L�� �/O`09aC�4U����"F�W�պ��S�<�YsE��o-h([ŀ_-Kg>Q�!�1X�����3V	���T��>Kt&���-����Kl��Ad�a�F0�B�l���d�>N`*vDc����~5܌�SO�&�ca/D�{��P;V���M�Ѥϻa/�6 �/#ےU{3��<6��a���?
��z2M73)��s����ih���x5ʈb� ԰E��y����c7 E�g�,}�#�8�z0�o�T`�zv�-�&$�!�ŭ��P�Vd*SYx�8��C2Z����H%jH��BE�u�, ����/�T��[+PYz�HG�°ynx�UOI���|Q��~�.�k�O���҆�4(�:iBw�)����a+`�L��4N���Q��/�4U�$�ԴC�%
<�r�2����2]µo�CR����,,�pm�w	s��7�P-�p���
�Y�A��R'�u��$ۈ�B}�A"�+9U4]� aZ�E��ر��4"0��C��%�A� �Z��XI�1B��8R<iZ&��!�@)�
�J�"v�dq2�1"�	�6�l�Y�"`�5LO%7,Rq �f�$XHi\tD��7H����H+k��l�j��M��扡Q�xA��K!^��	�\l�ΧW�����ԩ'��d9"��u�(2���UxI���La&2�	�,� '-T\A��>�#�فEGN��2jN Mw���Bl�g�? ٫�@���je���d�,�����H��*����o��'�p��"P�K�4D3�̐�V�z�)�Kw��"�L�W��}:P����������Q�* F�	θ]���iQ�_=I
�$T>-���gF���yQ`�U;&�l�Ȅa�sa�bQ� �L�;OGJRYc��^+�YشsE���!���h���s5�K�C��aQs ˝}x}��G�e+�t �1��yP�%Xv�yQ���F��I� �{ti�%����th��0
f8���H״mL5���lqh(���	X�x]��������F'Ƴi"��5��u�	�f�Ir�A׈H����C��A,��h��]�@t���aΨ^=���B�P��Az�1O�ʅ�܏G#��U��EXu��H��_������4��!��K��t-���5��'�:=��k&bL[�#�J��B��C�Uw:0�ŋ�"['�(�u���$ 1��� Z�8�5� Y���J a�O<$�e�� ^-� �;j�D� �×i:u��z��@��
�wp>�'� ՙ���f��H�"C̥*�dq0�+[jA���,:�hx���X����"?� JJτ"c�AK�%�K�j�a#ȣ��|X��4^���dF�'2�4�
N&k� �C��0&���>�E	�@�<���x��Ct�dY���p�0�K��2 �	�_?�C@G�\�Ω��GJ1�0�r��W��4��.��<s�6CߥX@�к��Ӑd�ة3󇎖f;�}�e�ʭ�����C�v�y��E* ��;�-Cr�8��W�B�L�b�@I?V��*��#@��2�rO�?���s(�8Zud�N����)���s�.!X�'��^�|hHAi�' ��o���d�
Hv�IPΟ:}�����ڮ!9��K� \�&�,I��:g��0�?%�y*�Ӷ'�l�3&kP	'3��;B@�$"� U;bN��c��h#�n0$��b��[���ؠO�Bw>0�V#By}B�~p�<�3�@��qq/�,@Dq��d�h��k�¥p �06J�ً��y�V��&��	Zkc�[��H���U�n�ιH`�Ĳ2@���7>��9A��G�F�`�&�a�сDDJ9*X9Tn�Ukĩ; F�LN��g��/s^𠖯֢������/m��h�&꞉l�t�@o]�>f蒆*H�h��������ـS!��j��\�'��:VE	P����VlٌG:Du�JB.`]0�h���n͘�P�#��?	�eT���ٶ,Y�D;L]AC��fR*ɂ׌;,�	"SN�"@���ݒ)�~ِ�b�7�nY؀:}�����׫�����S��ɕa�t50�e�:t�` �(�)l��86c����7�@�FLFu#�`���0�r�\�z� x�4o�
�`�ցGP�ɒˍ�z7��6䄖*o��(�#ڭh���6 "�t1�FF*�|e����=���9@m��dv�(5� ~�>����\���V'�T9���+;�)i�-��`x|�85À��8���1�и��(�GJ��;�#��\���(a+9�p\I�DN<�?����
����ɛ<��)3�$î~�P��@�T���hS�ܲAN<Ĳg���RQ�p(H	5 �!;�$C.�\�������DI�g�P�����	x�����IX&��\rh1i�Y��hO�1��;{�)�"��44C@ C�R�O�=j N��~*TPksd� 0�$��dA����}�'aEr�	B�Fʕ���ʦ�!���;&�*��e��5�V ;��� A��M�5�%H��s��X��O������
,5����-�W@^����O�	0{���:�m�0�UE��oD"?Ȋ�F���H�k�(�D ��LolʙI1���L����">ʈ��=�����P� ��I�: ��߭b���P�IϏtu�D�#}��^���~����#Y��yB�E�J��t�B�ǺU�c�#C�P  �ԟNp" ���Z�::�z���N��$BRܓ	`�I�=7�D�phɝx>�m�I�|� �{�i
!�CoG</�X��O
L�0ȉz9�E�@�)+�DuX3:+��U�uᆂF��l��/Յ1tZ��
�z,.P	!�ʮD9.��#f�D�^���7��Z��'cx���+y+>xi�C�-C46��SƁ�D�V��;YcȀQ�Ix�N�RR*�6M�u��p����O��L��T�6a�4��`W��?��O��LCF��2K
x��"�N��B��d�� 8���'����؟q�ƕ�$+L�Z<���?႙#iךe�j0JGg�<�l"���<KQr�0�g��(���
B�ȧb�$���e�t0��JX�%}�d�h2�O���+�܏Y�,�֤_	;8�%�\PclI= `@hCI�6~`$���ф7ˈ�sa ��7�a��`DBV�R�*�>|�j�Ŕ+ R�aŐ)4��}�*��z�� �6�I� �4�x�I�)$�}(��C�F��pc�����:R#�>�A����y7m�$=I�,�s� )!|�r�
�&�p>�Ջ]*U�n6-R8��@d�M.��m�O�?�����E�����oٖ0����#�,:��4 �-��q1CK�;8�Ī�\=t��ު2������A��� �?�1�ޚa�|����<T`:A��@ ��9�KG�j�� .ox���a�Jjf�h��dc�1�hP�����$Ԓ�bfQ.r��t9�L�#����	�z�x@�ga̞�R���P��d�竆6y��]q�ٜ'���KeH��np�׏_�&9K��Q9d�ܤ��ݷm��M��*?V.�{�mM�_�����(!��P"1��r掙�-Y�}�H�R
L�#��K�ێ���T�$��P2!�ؾu떵�YD���Q@Vʅ������ӧ�Z�D�hu��9\O�%���Q3^հQy��& 9a��Eb���ČA�T:�!�!S#MXԉ�F	�H�`sE!C�d )Qb�Dj���D̀4R �q��%�ȱ�֡�-#��riI3}�t1�y)I��d5a��])k��"�/̠E��(�O@M���ϑ3W�9p��* �a;���-<�i� QU�-�R"4g �q�bcN�5Z�DxD�P�ԍ���,��aÁnߤ?yR�S�/\
�-آ��6���0�+ ^�j5����N	y����#Q�����g؈]��i��	0�j��|$џx3P�M&5�a�	<��șP���uB���'<<�$nV!=0DQ�'\?����2I�|-�AC��`(��4�������V�I�l'	�� �)��8��V�����"��:И,I9N��bgB+�����bcX�x$�UڦEHs��8���kC�͈�v�r��O�0H�өν3���X!X^DѰS�3������j�Ҭ��%�9����͍>q����VO��^SR��#)��O>1F�.�B�c�O�o��Li��Эa�d���N�<"��)�F�L�C��r�W/�R�Gxҭ�6M8��
�b�*HEG�_�HA�d��F"�) �
� V�|�O�%0���U�v0�u͔5H�P$#��خ<9���@�b �Go�4�Ŋ�Q��hO>�٥��@��#1�#C�V(�A�� ��X��N4�(,*%��$m�Exd��	#9��H�m�b�QҦ\E�J�� �q�1�M, �&�I�$��q���	��D\�df��g�F
2����P&�H��]*�&�*|�|��p�K,tL`�����S�r�������j�d�<>�>}Eh�)i6�E�0�,tNf䃳��W�b������c2k_9OØ}t�L�4&~���[�$�汣��EMޜâƣòUXB�8M��y��=�p��Od5�Ј )=��d*lpP @�������#�%B���f�l9���� �(Op�[��T�P�
 ����HǨl `AF� �Hc5���=Vx\����v�c��x�����Mƹ�N����S�R0H8@�
S������j~4�sae�hO�2�U.?zdH�"ۜt����W�U�z���)H��4��ܞy]J��I��y`��89����V�0�!+%��?�Ya�<]A�J��G���*�'�[�1���IQ�Q�l1qè �R J3ܞn�i�T}��i0 ��Ԅ�p3� �~�G_��l��4V
\��G?����o�ʧ>��I@/
�x���Y񮖆'J�9� �� Ӈ��p]���şA�
���C8�b��핈ܢ��!L�?MܩFa��y�mZ
zΘ���c�3ʓd���3S�C�;U�t8��G%�,Fk�3�4���%̅�dx�qk ����O���ɏZ 0�e�_[�T�֤�8	����R��6����	 uX�țue��i�h��V���;�O������"��5 �)��:�:��0�.��u-�y��!���O�RƠ�=l u"'K!2K
|��R&��MR �Ռ@vs� ��NŗA`��O��J�<8�����ؑd��*O�娆��6⸧(��鹓�^�N�Pɉ�kE,���i��:��T�Uk�Z��bk͞t���E��wָ����+b�Шb�$�\	�'��LX���OQ�̓�������M�T�l��$%<Z܆��O����љQN|T�qቜsPxS��!�}B盁#��$��EF�ir���<�<��%H	7
T@T�&VPa~R�\;��)E�Ҳi�Z1�B����Oī�T)Jɢ�bM|2��/�B,33	��8Q�an�b�<Qg&�/N�,���+SFT$��/�G�<��o,�5Z�/��M��õZ~�<A����$(b��ʞGJ0�;�'x�<��eW�+���iR�RJ� 3f��o�<�FD�W�:)�V�W2��9���l�<�ǈ��"��p�R�)�HcaeWm�<�'�V�H/*�(n�� �Dk�n�<Y�GC?m��L��oS�;��Ʀ�]�<�ЃH��|(� ͖o�P���Bm�<QT�0��
�F'��l�a��p�<	עݤNJ�B@"��)���e%i�<� G,D��\�7�Q<�ʴR��Od�<��ō�6ǜ���Z�%�z��G͂]�<��LQ��D�X6;z4y��ܹ~�!򤞕t�n��@E�a\�=JB�R
^!�$�5o���i�[*�Џ�0O!�DQ75��0'FQ""�8r���1,!�d��i��y0hǫ@��VDћ!��ޜ8gvŻ0��PD�@��e
!�D��`X~<�4�N�P�4��%1-!�U�9J6��b'�Z0���1@�!�D4ް�a��Vڔ�ِ&J�v!���[��wIV�1�D���&y�!�D�(v�1:v� �`��\p�j�"O:�at*K����j׭�>_��H��DH�X��tcGB�A���AOZ,q�1OpP�WB.t�V�q��M��x�a� G%D"�J�M5}�.!��<����2.*	�eOI�H��a��#*��'3(��>��EH�ܡ�ٸa�D6a0��O9}b�^	m�dpw'>�Z��o�.�a��k��� [�t!�(,t��X{'�>��<%>��`�v�53��_?6����&Eu�h�"3O���O�"��@����C�C�r��q@������3p�qO�?��� �����F�>����AEZ/Y����Ox!9��t>��Ǭ�<_X��k��F��t�hFB�[���<=(�Ѭ�J>��R۾yȀ��yѬQ����>����<�v�"}Z��~
B)q-B8+��P�ȰҁĦE -O���O?7�ϐ �.$I�^s66a�B�7'����HOQ>���̙�4u�U��{����O�MDz��iެ)�.��N��r�����$��|H�#=I
�'r<Ոe�ǵ�T��d��8���k,�	�?)��ؘOX��>��U�3�īq8�2�#�4����6��a'\����M��D� Da�J
���GFN7F��Im�(- R�ԟ1O� d1��Q�]|��#�K<S:��"�i_�=B��/�)�2��5�&&�3
�r5�p�S�sM�!"��C�&����\�d�arD�+[&�P�MvqO�P �O;��-��O�dX������7^�~����yy��p��֋����S�O���Z�b��@�ǝ&h�U� ���0&����S�O���Z f�f ��f$ ,�p�d��O�����?y��QZ��xR(nxZSBf�I�e_'���I`y��iH�.3%x�/C5�8ċ��
 �!��Ș2ڀݠQ���5�Փ$!���1@���p5��h�t�ۥ�Һ�!�۷=G�ebGi�F�5R�.V�I�!���_����S��9ᤍD u|!�$Ԣ�� ��d��L�W���W�!��jA =yŅBU��	s�~M!�S�K�bM;���$����Û$;!�W�yG�t�"N�-f�!�¤N�-!�T�B�^�BO�0mYX���Ü��!�!7f���5��@D0����7U!��m������.b��#� pR!�8|��X�V׎:D�����u5!�D	�=F���Üc$�	�T��g/!�$���Ι*�G��r�}Q ���!��J4Q���G圈1
�`�$Q'�!�dߓ	}����*f���s�֨!w!�D& erl�r�� ���s^!��+-��e� \�j����g+!�$ٖE6p�I� ������B�o!�$X��`�rA�2|�h8Ȁa�8!��:^X�8� �r�D�#���u !��6V�����̂p����lY�O�!��&j��;���B��Q)3�F��!�d�q���7ۜ}�*!��iA?�!��/-���&����&�B01X!򤃖gʎ�3R�C��L�ND!�d�;wJ���lD7m��R�<!�$ 
5k�@y1�=$����ME(1�!�d��s^�p�M��7A�-9�/C�v�!�D��~�����3i:(	��ci!�d(d�Ƚ��$ؐ�\�i��*T!�$�:|��-�&(�@���x���!�L&BOܠ�5�0;��]��:���Y�q>\�:6=Um$!	BB�y�]�uy Xf*��Lp�al�y��Z�%�l�j�n�;f���#��y������Ak�*TnrR|�0̎��y���	�� �UgJ-l�����^%�y�&g�������U��q��I�yRj�?�@[�FOb%�!��y���S��8D-R�oP�mk��j!�'��X��
��pQ� a�O�}Zj��'�t�"Pz��G0P�����!D���F@R
��,h���lJ$q�J!D�ti�埗al��wFS�`�Ӡ!*D���RK?��8C n�(l���I_<!�Ũr�r�(�ۉB�,�@&ʚ="3!��"D���c��\�/_\��SF�}B!�$B=~^����E�5Z&P�W���r:!�d�=�B;�(W$DGv��Rʊ9*W!�$��61U��,*(I��KR�!�d7I�\���@P�s�0 �^�!��>JQ�1�l�k89X%�9 �!�ĹcW�"UIN�=���"���8r8!�d�i*\an�#=7�!ǂ�	(!�D�O�j�U	O�q�ν3����|�!�� �1臋B�H��	-�@�E"O��(��Os,\��!P�]�"O�飄�Z���T�6�B?l#VѢ3"O��!���4h �Ö���o�yJ�"O^8{�	�Y�t�Y��P\����"O�@KN9 z� �7I�<&-\峀"O¬�GdG<_����N &�l�"O\H��*H>��孜g����"O���agY$Ed�a��L����`"O�+��V[���!�X.��k�"O���q	N�U�Ɲ�5	ކ]� D��"O�<�ł'8�LأEX����""O��B�D�^�F��e\
I"Y:W"OnY�bM��S䮴�DS2>ܑ�"Oލ	�a^2io���5vy�v"O`��B$TWl(J�P�i	��x5"O ��b����[e��4�t��@"O�`)W���,��.�#9�-��"O��T�S���z�,6���s"O��0���{�~m�P�M�P�x���"O�q��Q}-��Ҡ��W�D%YW"OX)j�Kv ���D�����"O�m�+.	����`Ǯw��uke"O�홲�� ���� M�n^ͻW"O]p&�ٔP2�$*B��0p ��"O�ř�!�4)�@�Κm_����"O��bދNצu�v��b/�e��"Ot�@�#�	`l��OY8;��\!T"O�,��)ӺD��raGR�����"O��е"�$L~(�A�_�^�����"O\IH�G�L?��*"*�E�@�a"O体��3c�e�%F��'|��A�"O�{U����E���� +1"O�i��	L���҂�.F� ��V"O�|pe������*QD�l�"O:�R�.�
�1��%
���'ʀ����`}�EW�_���	�'�0٘C�Fb�1F�M�l\��'w� @BbY�y�|�s���#	M�',��F�� rfaa�
4 �潩	�'D�P C�,|0��˖�͑%�\C�'n��g��1qeDxL���Բ�'/�9�_�s"��zf���� ��'����Ad�����Ǟ//{N��'$fI���Z�f��A"��V7QX��h	�'���!�ǐ��ܱr�邐G"4�P	�'��A@&j�1A;���+;3�	�'�6��d���"���
�8%��'���R3i��io�m��� ��5{�'aN��u �M��6N�
�jdP�'M�x�D����Y�l�x`�h�'¤���7���btD<uB�$��'�ڀB���
sn��D�O!��b�'�ؘAv��'����m��I���3�'� yaC���0F ���ʸI��'�Byk�H�2c#|1��`�&
Az�	�'8��`�� �|S�t"!ֽ	��'ZLz��(WF5��ѴxR�k�'�IR�0C�q��	��r�
�'N�i��^�jWp�₧�0u%��Q
�'�(��� O�v��Ūl��	��'�1���$H&|�6�N�l���x�'�.�见Ȩ98�����a���'�d��ᎾK�H�(%L��W������� jP�S��>Iq�K�	�	���D"O\`�'8�M��� �z��"OpX�i(F];g���-�"9"O�M�D�(���3��gc���"O�	P�@N[]#V��7
\�"O~0(Ê��	��;�f
;o@a�"Op5�ᭉ�l��}	��,Vݲe�B"O�mI��N0l�8ebT�"!�%Z�"OH\���I�>�`y@FD���T"O(ظe��&t���h�j���q"O���FG� ���"0j��`@)�"O0�1��f8x�1���O���"O]Y��š��,	�8Ͼ���"O�y�m�#<9�u�A�8}�Z�9�"O&$!�*��\d�	P��"w �Dp�"O�4��_�6z����²*����"O�tC�@W�0F������0k�"O$�Za#��bu͹�홛_7F���"O� �w�P~~I���H&$��G"O�j�kG4n=��#��%!^q� "OH�V�,X��tH�˘}�t��"O�Sq,�>�P�)�'K=,�;�'���"V�{��f��h�` "OD- aƜ�9��1�E^0u�����"O���)kt������Ma�"O���G��.B�Y�3>�*HS"O:��$�Wf�B�:v'
-""O�`��Ӣ~ȅ�`'�	6�JT	f"O
�*U@+SD<zG�Z�p@a�"O���cӎ0kjD &�IiP&%P�"OP� U��&mΉƤV�N�$u�"O�pi��ʚI��Q�D[�B� w"O0uPƦN�v� ���⊺�(m�q"O8p!L5�|A�n��r�����"OZ����Øxo���p�;i���"O�LzBdƓ!:Pg]=YȰ`�"ON��r� ��x�&R2 ʐ"O����H%2=�XX�eJ�b � s"O�=�w�Ъ'�B|9&�EkF&�(�"OL遆��r��ucA��Zq;"On�	 !΁[m�6L�Lv6�'�ɤ�� Z`je�R�7s�=1�'�H�`eĈ	!#�@X�&�?]0��)�'�6$j$���e.�����9Q�@J�'c�q2g ��Q�$�{BPw�B�
�'�Dӱ��x,xQrM΢h5��'F2`R���wb iz�)pi"��'6Q��M�:A��*�-�����
�'4T!K0!>%��s�D!m�bd��'I�eS0�7t�.��%�Da��P��'i����A�[�:P!u�U�$�A��'�Fd������闗o�$}��'4]1��G�}9�Xc�A�$R��Ы�'Y��'"Ssz�K�.ѮDyBU��
f~ճ��M�~�H H���c��ͅȓ?�\��ޘ)�5��T9npp���_�T)��Fk���	�&�\@��8H�����MuN���S�}����p�氓a�_5�r�O�(T���E�v��V#45p����܅=�����n���X���f�G*h�u��D֨��񈋥��QićK\h���ȓY>�ЈA�ŜR���qF�>2�4��ȓo7�����,3��5�1���[�Z���S�? B0pn�>)p���ǀX`@��"O�Tʶ�!m����ҍnf��(�"O���$6sRH� F\`n�RT"Olp�	4��E��bJ\���"O6�a�%F�iS�Hy��حD[�ܙP"Op��"ܟPR@ ��f��jzR��"OƷp+
�8@x�Ӭ\A��@"OHe��F��!��iQ ]4w#����"O�$Kh��Yi$P��n���%�&"O���th �(�$�9�,�6`480�"O�ْ�/Ǝ]Y�-3'��N"O����^.I�R��
Ӥ~�$;�"O$80�g�5xbQ��1��m�v"O��B�   ��   �  i    �  �+  n6  A  �K  U  !^  �i  r  {x  �~  m�  ��  �  7�  y�  ��   �  F�  ��  ̽  �  S�  ��  ��  ~�  ��  >�  ��  8 ! C $ �+ 2 b8 >  Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�� |d��"O
`�(�;���8���-0��1%"Oj4��ND^[��"3/9�0|H�"OB���H��*�ʞRy=a"O�味V�!X��!&F�:J�$���"O,��a
���C�Ą�M�"O,$3%o�-���p���+Ն�:1"O��ݢ1����`���y14]2��i�<�6��{_���c�H�`�fX�$Kn�<��A̼VI�xR[�)�Ć�pඤ�ȓA5��('nߡ4�� �)˩%� ���,��r�؊b#`T�eT09���ȓ!�b��g��}�8�F��-? �ȓ
K|m�ș�VṔ���2�%�ȓ"R�X�j�4JN�1�˘X�i����̹	_�jZ��1!g��zܶ��ȓgil,*�J�
j�Ne��i�J%b���f	�(U��:���G��$Y^م�~r�� S�%T"���k\�jx�ȓ|4�1�îJb��@ӵ�ݩn�V��/[`�"�v4�R�!ʎ<��M�ȓ`:��z�ؚh�J�Z��$HY:	��H��p�m�C1��!��B:��0��EnjZA V;9����J[
2���	��4'J�EA�IVW&��~�(aZ��ӹ�>� o�Y�|�ȓ�f�A�
Ο7�H��M�$�����mޠP����/���ANXo*�ȓTv�����{ ��-7�*h��I��sB�8�8���3����ȓNe*M�悡;������X�o��!�ȓ'lj�#F�m�+R&;�|��2)n�C��0S4���T:
b���:�0!��e֊��)��ͷV��,�ȓ0�&�8#���� ع�L�����;�P�AFd���,w�6d��r�EQ�( �gVlɦ�M,H��,DP���|�I	$G#\���ȓ"�)���E�B	yt&B�^�LɅ�4�� ��gëF�ڙ��n��R�p����?�  ��[Q�q�oY1]N�$�u �P�<�0�	���)���eL����N�<��*�%[�J�z�D�(lf�䀅t�<i�*I3ъa�n�!q���H��@p�<�/ӷ,X�C�ni����\n�<aS)Y%֌[�eʱ�Xp�Lj�<	�gA m�&���nݤ,Y�%`�Rd}�'�D���B���A�փ+˪Z���I�W�\4�u/��z,���bC�Ƀ�j]*b.�y�8Fh���B�	*���2�W�X���)dc#��B�	BY�pRVz�D`���Y)���>9�c"�'}�2H1!!Y�~O\@�R�4�&���w������
%`d��I�2=�<��'א#=E���S:&`��#J&�ja�K:X-�ȓlX��0��CC�}�B6YXl��ȓVp�� jЅ (�A2nF�W����L��A+Y����y�*�!v$���� �maѨ[�.8 �mIa�(<�ȓ/L��8s�A-~(X��R3�愄�����	�8�Z K&�ߛNBa��"����wi�=[;�8[�]����S�? � �fZ(�D PA+ֽP���"O�H[&Ҥ_��I%ˑ�Y�"�;�"OfPYDaB-6l�my��τ{���""OЌ)�������r�(W��9�"O�|����*^|��/�iq�B"O�E@�B�*;z����I@�]Rg]�TG{��)Ș����P�؆���J�>�!�$4,��(�����l�����s�!�d��	r@)�,ʓ>����$�62!�d11�Nd[R����H����!�޵2��9r��A�Zvh��)�"[[!�$S� ��qHӽ}P�����C�dv!�DZK�2�a�-
�p�e򑏒�9s!�Ď�*�~���fW��`�44^!�$�T@n�%��5Nl�D�Ɓ5P!�D�!F�m!�*W�M5`	� +�V`��Y����G�]9y��s�D�>N%J��6�O�T��s�κ6�@qa�U'	�ܵ�ȓ(ߤi���GB�	%kס2���Gz2�~�gjg'� H	y�Lh
'Xy�<�-�" m��5bE�g-V��0j�r�<yB��$��h3W���]<���mTl�<	F�I<y�$��aD�	X�i%���<�����"d=97��
{V�)v�Ɩh��B�ɹ+<|��FEį,xX(�+D�_.Ԣ<��T>Qc�kЈep��2҅��7L (zf�)D�(�5�٭oJ�����2�&�BW�-D���e�P�4@mRg)��-{�p��(+D�,8fN�7c�X��eZ#�X|@Тm�p �]5f�۠�?�Q��gÈ|�qE}r�S 
�Hٷ/Ѷh�b��o�u$�B�I�b��(bD�1
�M�P(ܖ
��C�	�"r�U�@Y�p�F�;5!6r�C�	�`�Z�ŭ�6z=$����|��B�ɟv^�9��	�G/!b�핳f�B䉦o�Ձ�i�l �\�w�1J��B�I�C銹1�� U��gH�Fi�B�I-G�L�Ӏ�
g:h�r@�P-<k�B�3J�C''ȳg� ��g:+N`B�	�l/��3`��q@�Uy��\�6B�I�����A?Y��@�[�v�LC�I�D�08��,Zz ai�jx~
C�	G���d�ѿYڽ���	�B�	�q ��A�/\�{��aX�Y���C�ɶ9Ll�ba���=�h���I\�?�B��z0pbS$��V���.[�L B䉠|T؁3d5���jX�4)�B�y�� ��ꄘ+ܘ����r�~B�	�)�RX�"��
�H];��xZ��=!	çyS8���FP�Z���n��'��=�ȓ�l]
⬛5~͆��Q�4����ȓN��ģ���M�ne8�c̑P"���S$p��Ъ>+�m㣏z3�t"�'3 �D˦\P�i%�Ca���C�'I���%> Lt���*��LK�'����p�ծS�*z�ϵ��}��}R�)��Ӳ%P�E�g ͆A�� x�B͓	�!��4� �2���_��8�W!��a{��9�IK�@��d@@3���pЩӼ ;FC�Ʌs�rlk�	�nDS���
��?�S�T�8�DIp,=ی�`�gL=�yB��?I�L���J5rψ�qa�ʍ�y�jZ(���$�!:��7����y��T�c��i�Ύ�f�*��7��y
� �-)���}��Ɂ:"�0�p�'�1Oʬ����KvbX�i��m�j�#�"O��3�x��T�K��<%)b��[o�����-���)� X~H�6�ڡ"
B䉻(�N�
dŔ�7�0[���6�8C䉜^~�L�A�.NV�lsŬY�t�*C�ɇ^��GƇ Q,��Q���Y�C�	�S��� ��3�x������h��B�I+N��<񵭝�[�B��R#�%.�B�I�j0���@�	"*�U����C�I;`+x�w�S�W����5-�1לC��&+;�x�S�/̜��!�/bNN�	S��h�]@��S�'��&Y<%K�&���yr	�0���@ͅX����&�ē�p>g�UXe[6�K�!�T�h �W�<	�H�g*�\RUDҥ6r:*Ml�<�'�á=�	�@kTP���(ͧ{`��XG��w�� +���/b�(+E	Ӆ`��4�˓�(O�,[&(�Q>����R7 �����"Oj��R,�!���fCWh��D����l��OR�X��hq�fF8?��H����;1�А�O�y��	+yC.0$ �\Nڡ��
�0����O���>�O�L�l�¦��?����'T��!x�!R5ז�
B �]؟��I���)��n����ѬX���N<i�4��$1�0*�؈��^�N,�8��U�3DT,��I]�'��DFK�r����AC� �Xsݴ٘'c�)�3}"oQ�s�b�C��_�!�c�6Аx2����t-J'���Z��P�O}��Ҧ���I9}�c�l��B㎁X�t0�j4D�|�a)��b���!�v� ��2D����㓾��`��E�
ت�g�:��hO�1���U���s4RX��� o1hC�	 ƠLRШ��f
����u3PC�	�i���	�Q�As�X3d���LL~C��-Z���*e.�t��`s@nE�2MBC����c�m�8'�����K��w��B�I�7J���FLP�H����u#C��bB��^���(��O�K$r���՝c�0B�I�$J���T�sET�&h�!FS�B�	� d�<��m� p�D�(wVfC��;. %��^�_�`�s�_�3�dC����|��7
��1V� t�C�7l\j\��	9	�PhS-]��BC�I�i��A�b�W�2K�+ ��L�C�	�-��(Q��I%z%�whD��C��4C�����l��@#jq�aGA��B�(%Al���7�vرE�_��<C��]r����ݦ�����Q�E�ȓgm8�
��D�tSh���N�n}��B��);�MD���yE/�����XL��r��'*Hn������IKRЄȓ���g��F�$a�K�)oر��m�n��E��3`Ml���Hj%$9�"Od@ѣ���JZi+e�[�f�su"OSŁ��B��Cbf��Q�q@�"Od��
P%���d�T4����"O�bRe�3*4y0�A�3�Dx�"O\s�� I!NaA@�,-:@�"O@p����=Gu�\Kϐ�b�rT�"O�i���E7 ����rN̖y�(I2�"O��&��ʈ�w�djx1��"O�ix�#� w�(�ـ��5x����"Od,;@�O
WI����&t�l�r"Of,��NM�:��<���.�\e�S"O� ��ž*�Δ��'�ppQ�"Oj #��`(����l�k�:%Z�"O�Y�@�@��x��/ �zēB"O�1�R`�����G$S�*)XF"O|1a��>7�����B҂J{$aB�'*��'B�'T��'�b�'q��'��x1hD$�ZP�@G�}"�t�u�'���'y"����'��'T2�'�pdk�H�j��L�S��/'O8DJ��'���'|b���4�'�r�'��'����q("��x�@�Mq2����'�r�'��'���'���'��'�@�+��A�wC
��R��5^� (��'�"�'�"�'���'x�'L"�'�:��2k��~*���o�S/l�2�'���'���'��'72�'e��'� �C��!Rd%�)�4x��H��'�'���'zB�'*��'rr�'��b3��;���3���i�h �R�'�b�'(R�'b��'-R�'���'��Dj�F��(��q�6�ǁZ�5Yb�'Z��'���'��'���'S�iL&	,��ࢀ�!ɎI���E!>[��'3"�'���'��'��'Q2��O� !��Ls$�����4�'�r�'���'u��':b�'��
+M�-�gѾ
ۀu���� "�'b�'�r�'W��'��'
��$<���V�. �D,FT�2�'���'�b�'Fr�'�6��O��$Я>w�`r�ä<��\(��ߨv�h��'�bQ�b>�FZ��*�
�H�:sIłl3h������t��O�(nZҟh&��s�hA�4�FTS��8K���~�����i�r��Nț:O���2?<aa��.�ɯQOV���M4m����yюb����My���c�L����T4aȐQp%k�&	�4K���<����}��G�p��f��/{�Z<SP�E;K0
�m>�M�'��)�S�E��<n��<����	B�vD��N��e�	C�H�<q5h�7F��8jF웰�hO�)�O�AY�(��O�ڌ��p��)�9O ʓ��y��e���'���Qv,A�
u�Q��K׎Id$���M}r a�j�oZ�<��O\�PǛ�[�	��U�1R}�������M:) 0�$.�S?#�(�;8/���,'�ڍk���/�t��bLB�6I�IZyr������"G�v4a4��Y@4 w��Z���ڦ1���+?�P�i	�O���X����4]֑!n���dЦ��4�?��$��M��O���n��R�	�-�w��Б�gt���k� 8�ГO���|����?����?���z�:P�0n��*��@[Ə)u�^k.O��o�0*D��I�l�	�?���y2��8��q�d���L�{@I�Y�\�ٴ�0O$�����O�D{Î4��0��k5�.9%��*�Z�(`�<)1�F"�x�B�
��0Cc�H)%-�tIbc�"f]���ː�7��.�*L:$��h����T�����G��2h��m4�-hۑ����H�tl�'�����Z?���[�d�{g���<� ��{!����y:bm�A_(�MR��y��� kك
ب �@�#[��a:�)�
8�N�	�
Ts����E�� �l֙>�x��C'�!�p0�O���#��������$�X@�$Έ�6p�S��*N���H
s�zx���4��\l��s�LI N�3A\���dN�k��X�O��D�O��d�<i���?q��|��N"ro����C�<�$���L�&����O���O4�`�M���i��"r�h���a)Y��`q��Kx�j޴�?1����D�O���\�w1��Mt��S>PiZ���B:����Ǧ]�I�ؕ'�x�Sw�1���ON��ƸX��Z�Y��8h��%�����i@�	˟,�ɝFc�c>%�I�?7-
-�h� �ɨ,�.逌��S㛶Q��(�oI��M�4^?u���?eA�O�t��(B�j�f���'�(�NL��iTB�'1$lITR���&���$G^	Z@�_"i���y��Q��m��Ɵ����?uyM<�']��(P��h����ѐO�F��¼i��)[]�x�	ן��3�ş�E%\$\�b2�:%#P���l#�M����?a�)�H �x�Ob�'�p��A���/�M��&ܕ9fm�>���?	n̓�?����?)Cf��{�0��SU}\��S�ÉZ�f�'\���#ů>a)Oz�$�<i��Wk 8c�!�V��`�F�k�U}�#� �yR�'���'	B�'$�ɵFg>���ȱ�)���P�a�&ԙ@%��D�<�����d�O ���OM
$d�6��9���U��n͂mN�$�<���?��?q���J���i����ֆܽ�$����1Xz����`�6���O���O����<q�S�N���[�L%i��q����4X�@`�L���	�q��0��Ɵ��Iٟts�I#�M���?iS�ęJ��	��}ʪ�k�ݫ��F�'��'�I��X����~y��O&�3�̕�^��IrwK�LUp;��i�r�'���'
�ѹ�$y�x���O ����l)�@ʝ7_y�$q@*��C��Hy!Pᦽ��oy��'��A��O�2[��s���(!mȂW��,�"!7J��׼i$��'����*iӎ���OL�$������O�Is�,�86�$m�F=Y4f�8���g}2�'����!�'$�Z��L��R-(�5�Ň����#�^��֫�#`f�6-�O*���O��� �d�Ox���`i#!B.~�T��B�n�^�<L�	^�i>M'?a�I mS]�PJ\�\E^�����4O
l���4�?I��rڴ3���P��i��'-b�'ZZw�Lqi�H��Tr�|Zj܂`��bݴ�?�04�p0r,��<�O��D�'�ҥ=� � 2v�Q��ҝ��(k
��Ǻi�rJ�#uj�7��O���O��D�p���O��	��R�*�`4�$�O�`
,\��_�ȺQ-?����?	��?��?�5g�U<��hv䁱<z�x���
D��i���'qR�'C~꧹��OX�!4��,'�~� c�?wL��'!�a���OX��n���OlʧF5ʀ7�i�fՉ����,���CS�p�x��gi�>���O��$�O���<���/f���ˢ�08r�WL�^2���"T��'{ĝ)#�'"��'�b� 4G7��OF��6=v���"��H6�qC���Ky�Dl������Ɵ�'���.���X���0&>v�(5�Q�X0�j��X&����ȟP��ȟ�	�o��Mc��?Q��B�����t���qA�Q��'nV���'�����C�No>-�	xy��M���B%P�J����z�T��NզU�	��k$�[4�M����?a��J���?YWi'N���6�P�k�dh�"�U���	���!�	�ԟ���矜`�Gv>M��Ќ�F��B�xqh�KP.J���%�i���z �y�F���Oj�$�T�I�O����O�	���:����m��	\� ��M릍�T���_y�O��OVl�%
�B�r3J9��J��Q�e47��O6�D�O��aL]�5�I��L�Iڟ��i�a���T>k�f�iV蛉?�&��t�|�T�ĺ<��"A�<�O���':�ꔩ����LK�n(p��?m�7��O��Sr�ͦE�	某��ğP�����	�M�z�K���NWNL���YH��i�$����O8�D�|���"�:pJш�$�z�TL�<�R��tKO�h��v�'l�'�̱~�,O���'9������KIT2Vh���2���:O���?9���?Y���?�u
�8��֍F�jrR�KS-�
�X<H��C"�6��O����O��$�O���?���V�|ғjqO�)��hӛ wN]r�/�4��'f�'3��'���?1��6��O �$��~ [�&��J���?�$t	r�i^��'{X�|�	�h���� �	�H =pw�Í�B�@,��d.��t�Mş8�	˟L���v�Ĝk�4�?!���?����j�+�i�2X�8��5V�Z�°���i��T���I��<�Sӟ薧��4&x2�`KޖW����B�W��J9o���ɡ?)��4�?����?��'���3~�e��̳W�r혁f	!V<z1\���	� ��'V�i>�ӺK��ҁ{�Nx��oG+4x�P.���Q���M��?����b�'�?!��?qu��o�����20�6���>2S��R�-�b�|�O��O]R,݈y帍��αHrp�` �I!�6��O��D�Oj�y�)Ҧ}�	����	��$�i�ѨA�R�"w᝴=a�I 6rF�v�'9�	�F��)��?���"� ���,:�(1�t���T����i��޼`h6��Ol�D�OB�A���O��'Η�_b����;O�!3�i:� U>�y��'�b�O�r�'��$����憔�X��-	E<m�y�H���M���?����?��]?�'>��W,)��XVF�:��1� � ��XA�'b��'(r�'�2�'��ùd�6��4}��+_�u��d��k�&�^ym���IʟL��러�'("�������.�,���+d°���2��6��OP��O����O����e�TloZ����	?K��U�M)d4bE�5��Vx�)@�4�?���?�)O��D?;���O����)p�-�xM���c�6�O���O��d��x:2n�ޟ`�	ڟ\�S�@�$�سb�9lz�RUa�+;s@`
�4�?�(O\��ֵ+V�i�OT��|n�/A��B%84�*��G�$Ң6��OR��߽e���l���I�$�S�?-�	�f��=�Fj�=m��+D�Ȟ!1"�Ob��ׄTc����O���|�K?	
"l��z�xp�)\�@���jS�s����������	����?�#H<!��C�& yp�_V괥cL�#ZI��i P���'�剾�H���dǉN�XcE��8��Ux�� ���mZğ�I��rF'�ē�?��~��:D��]a�E�}�֔r�(<�MkO>�ł�x�O��'���.Q4h1q(��5�SĘT�(7��O�rA�v�	ԟ���~�i�]ò�������u�إ)yJ�����>	gh����'���'�W�<9�3V*!��91k6 ��6:�#K<9���?�O>1��?i�-ͅH�(�# ��aV�-2�
�?-��͓��D�O��d�O����͓�0�zp����6W>8
�iJ��Ǚx�'��Iԟ��IПl�bOr�LY��ەs�X]귀o0(����	���d�O�$�O*�9��dƝ��\*ji;v�غHH�(#� ��V6�O��O�$�O���,)�I�z�h82kQ��,��!�J�:6M�O��$�<���>7�Ob�O�h�S��(u�Tb�G�u�Rh���6��O*��Z L��6�T?a;���,6*^U��v�,	���S����܃�MkZ?��	�?�c�O�౮�0|�F����M*wW�;�i=��'S:a���'��'wq���+�䑍�~X��^�FQB\Kֹiת����}�T���O��d���'� ���&|i��a���HD���&��M#�4W\Ba8����S�O�� ̠=������sâ�ȖA^�Iӌ6��O���O�3�iEQ����N?9�̆�~��co��#!@p��eJΦ�%�H떎g��'�?���?	��ѧ�����ѨUH�z`O�2$8�F�'��sU�*���O���<�����h0A���j`aA��5L����Q��	��O˟h�'
r�'7�Y�d2�W�Xp%{�؇-*�0�.L��j��M<���?�K>����?�s�ڽO|H�:��6��!�˗��u�L>����?Y���$U�l/���g�? � ���Y
w���Ӏ�s���Y����ޟ�'����ޟ\���������9(�W!��f�itFȚ���O����O�ʓi�䐀ǒ��@Ζ7tN�1q�]+#����	L�H:�6��O��Ov���O�d�G��O:�'FV��g	�y��@딍B5R�H�2�
C�ny)Dm��q���R���//��$�ԑI�z<F��#|�� �w� ���-�~�Z���UR|pz	�'"LÑ��|Y�Ae		.J<��5^���'%�S���B�̆5((!D[�sF��QT�M'$���� �?C�aB�F�5&s�=:��W�@���;N��� վiԢK��!D; �34@�/]����>���t�1Z'h0�ᑈ>h4���D4�$�X@j�]YpEܓC����0��D��j��'"�'���h݉�c�RG��bfF��V�� �sm���u)����?�@�	���|&��b�HĿ�r����Rp0�ࣧ�55��h����?h� �aQ�	��>�����H�c`ƓS���C_
��r��7OO���/?�S�@��S�'AT�@�%\�k���Oy<��'֨۶m�?U,ͫ%:}�Ⱥ�O��Ez�OP_�HG��3h�(qr%�q�M�Ч�:d\�ؑ��ҟ��	����2�u�'!B<�͐�I��;а�ʇ�ߥ1�<�y6��E�!�[�%>H`0�:�|Y8bn8a�0�O0X`�H�8"�鈶 I4J���%?�rf:�O ��Ȓ�5٬u�Ǉ*q���q�"O��[���Gў<*t�?�:	����a�_2
�`f�i���'�Hl��H�"DY��(J��]#��'���ڇ(�B�'��i��2�"�|(O�9/^Ix���&JTQ4\��p<A�g{�<1D���S�Im��h�-�|��܅�	/N�.���v��_NJ���b1W��U����1_2�B�I�Sr������p�6,�b��	��B���M�� �0܆m�"��Ibx�$P|�d��84�i�r�'���c	���I3A��Q�OA�RȈ�I ��8�����ş�w
� �TZ*я-J�i�S�$^>��G�?O#��pB/ Y�#l1}�`S@�l�h�;w�𙒔��O�$i96 ��o�>�@�JP�p���'�.}8���ɧ�O��В�aS6�|�[��DgЊ�X�'�.,[֥�=�xZ�/B&em܍��Q�He��7.�0�"E$���g��
���Ot���O�H�d�M�w�����O����O��=IR.|��N�aRP��`�<�A�Uϼ\���O~�Ѵ�1��'ofS��^)��Z��n�@1a�
�fV4��!��O�]��Ƹ��"��xt/�/�HC��W(	�>]J��|�aW(�?�}&���q�ʳ(�ahceV� &58��2D�\2�"L�4��|8$-V�b�ƽ�#?��i>�%��z�b�.VSZ�ڕ�N�b2��	eG���IȦ�����ӟ$����u��'��2���Ԫ�%f����b�>�(=z�@�bɊ�"��4y_�p�+��1g8�F~" :	�b�r�jU�`<>��e�'A�n�!���-]�xYc�^Jb���o;��s6�Yiܓ^Y��i�ƌ�hN��$nT���T۟��2p���Q�C:|P=�u �W0B�ȓ{������� P�@��߱A숰�<��i��'��}X3.p��$�O*��F`+>��9����i�A@��O��Ċ�.��O��Ӻ	�d���D7_���!���Xh$4��I�m�x A ��\�`4�dϨ��O�ъ�ȡ7x@Ast��[����&��<�����T�@���CQIH)J�	àH�?'E����{Ri���?��xZ�x��&��U�&�GΙ0L�X��BEX(��.�Rp�E9҄��XՄ��=��&�,�bUK��J�����EBj#�'���Q�db�@���O`�'y.pe{��t���!��:Ot�i!p@�7bܗ����ɣ�~6D�e�4���:�A�?��O���k�
�	cpyH�[E+�e�O��3��٬����E(N�r��4a�25(8�*��˭U����>�'%<D�M�"� &P�Ky�4�Ɇ�M���i�R�i^..��S��8d� ��v!	18 1O:�$�<Y�����y�����o�pMk2���d�axs�$mo�<HhC5lB'�Hi� �\�(}���۴�?����?	4&�0H��R���?����?a�;2�pd�UM,�&|����RI��*�y�"���<S����l��9M2�uܓB Љ��	R'VHI���*�y���D�1M>���ϟ�>�OhL��nЛ��h�q�c�~@"�"O썩��ġu�h�镍&'��C���L*��ᓄR��z�҄E�� �A�%��9D`��:I�������ݟ�r[w��'��	ؚ�)�I�K�~���h0?&-��^�B��y�l�K���@�k�'���ǫ��5�8`[�C�8"�X�XV�D8u�b����ɷ[�(
ANەRvJ ��+�%�x��=�U˒#QRm��cC)	��r�%f?I��<��?BDX�:��5ۡ��'I�$e���GU�<� ��𗏍P���`T)A�u)Ԝ�%�Ğ榭%�L	4����M���?YbKX�M�^`�s��`��*�Ш�?Y��`sLxY���?)�O��(5��u� ��S��:$Ÿ+-r}�D���k�0�gF%O ��G$M��:1� �N����ʄ"�*�K I
t��.S	�@�.�	���Ɂ�ēH��B4����,�д�ȓvP���rB�����MYT���	����V�9�d̲��ұ$Ұ����'X<X��}Ӕ���Ov�'��(�n��%	�~�-�cLM]���X���?ign9��`F�ɑ7n�X�:B����n�T�P#�X���,l�B��-K=��%`��Q&�zQ�ă�*!i�����B=���E���{S��J��H�.��6-<DA���I�Da�Jo��mZ矴��卝K.���#굸R��^��?)ϓ&]28	vG�@�P�k��٢J9���HO~��5�>o��S�mH���L�$�즉�I� ��<2*�*f���h��ȟ��I��ݳ��L�|qW'�=��l+���$]�`r��CJi����r��>�S��	�s��Q;�A	;L?��慃	�2�x�hQ�qX0cw��uE"�(�hC�(�O�b�b�����OtN\���ւ4n��e�I;]��'3f�������BKd &��%
�v܃�/V� ͚1��5x��b�Xiw'ʠN��)R��#?)��i>	&��C��4�=pЭ�&N�� L��{��Pꐀ�ßT�IٟL�	��uW�'�R0�`����F7 �y�Ə¸E�L�S���&h}j�!�J��<�((<O�pcBU&;lC2kr����!� ���M�q�H�)���Kx�����n��Yc�F/{�5�U	W��t�$#�O�,�W�+m|��� 1!g@��0"O<��A�]�d���5$T"@r��DʦA$��cP����M���?r�?���� �0|����I�5�?a�P�n4���?!�O�t%!f�B�K�@��Gϖ=&lA �Ъ�d��w�1(��9
4�Ԩ4��#?�ץæc2T�I5
��iȊ%Ѵ�ٲ�0`���E s���3�m� SB�C(�
$���;4�"�ɓ}]����Q�	U�^�"Tŗ.\��¬R,~fB�	�-h�90�����2��&ZB���M+�F�kH��td �['�]�����z�,lh�i.R�'��S�}������)+.}�戝�C����N�E�� ����8�쐥,�T|0��L�Gn݂�йt��I�|2���v��Uz"�����H����K���4Cm
��C�%F�drPڪJo�$[���i�Q�Og�<:��L�,�������6t^�cI�(`���O��&��?��#"�x�p���&y���vG#D�d�Ѡßx\F�؅۰8@�� ..O 9Dz�� 1�]j���`V f$^5qͲ6m�Ov���OP1�"��Lt���Ol��O�.M�E��b8b����mل[���ӄS/f*U,�*X�^M1�����1;�|�zݙtj�Qel
;QL��pH�0U� 	@��O���6�ά՚�O�R�@$j������ɳ{�HKd���#���h% M�Ř'���H�S�g�	�d��H8�MB�o
BE�a,	qrC�ɪV|��3�Z�V�1�ĖNp �ZK���X�	�L��tB2哈dx8�ǰP�0�X�C��$��	ԟ��Iȟ$JZw(��'��	�8�3��,)x�M0@΀�A�x��RMQ,AZ���4|O�ys'�!dV�t���͜�bU0ah=*&�{W��v�:\�P)��(�RAF~���;{�ڕ�	���LtP���k�ɒ�6�a2"Z�7\� m���	�y�H%F�[PCِ,�j�9b�ʘ'{�6�*��R<7�,�O��`�A����v �; ��%�'_D8��'[��ir�'}�5�BPJEc�6�p��#��rX�z�$8|��|R��BU�p�L-5$F~��"x�(r��_�S� ��*��Uc��/
Y�T�� E 2&U1�U��2E����c�'�4E���Yg��B�>����=�
�q�R�P@{��V̓�?�
ϓ
wT�`B�7��Q�dT�e����u���/0�$�a�Z�R�t��t�\�#��U��:��Ҭ�M���?)�6�§$�O�h�$�V�2u�I�,�Uڰ��OR�$�6I��r�]8?��!1"՝f�����O��S�:�(���
�
9b�a+3.�'C�S��Ɂ"�ܒ3a�$��Rf�=Gx�8�R∽7�S&s2Q9$D/cv�֣@�i�]��$��2��S��+�\�1��=*�0E�	e�,�ȓ.�i�������)�M�1�T̈́��HO���A�.�LT²E�3��-)4*����	Οx��u�E�����������i�ͻ'烙jH�2��*SP0��N�&O��v���4೅*<���|���>i����}�6���[j�9UK* z���n(���(&�ޗ[��k��J��S�C/���8��
�9�<��%�-X.8�TM5�I,Z.0���|2�A.x���)e�V�Y6H�@Eٞ�y������ĭ^>"hX`3��2��d�B�����|
� ���%H��+I��i1�;D������tI�F��O��D�O��Ă����?��Oz��;t���682<�lK�� B��Q��	�W1R�ca)_�wj�TF~b�ǛM��D�̟+7���3a#J�X����ˣjC��P"��v&���������_pD%�d��΄�2�(�'�+_-`-�2�*M�l�D��=i�4�?�,OB��-��/ΐ Rg��4�6�P��]8>B�	"\�D�@��^��(��ۑK�b���4�?�/Od�r�'���1��矐��Q�T1B7C�	W��Ze�^ԟ4��N��������'w^�h���;wmSNR�-J�a� !Սs�����kػUL��!��@:u����7�6N�-��� h�0�j�;~ �cV&�� ��"��T���򀁜�T�Pj�J�T�I�V��d�T�I,J��yi���in ԰�
�	WB䉌�Q�5`B/&![&%��_�""<q��4��Yoڗ*�t��JȐ��S��?�b�D�����M���?�(��)�A��O lq��_*8�=!@�Ɂ _�p@�O:��5�Tsa\��M�!`G5fG�
1֟˧M]��Kr�� #*]Z&ږK�@�O����J�	�X��"/FJ(��2�C	�|�nAC1.�����J�+q~�
��^ >���cB���I����O�l'��?Q�QEO���ڄi ����w�"D��9ƭ�PJ�3"D�����) O�}EzC��-���g��qk��c�R�Q%�6-�O����O��R���AVp���O��O�
����0�*I����L�.Q�-.��,{�����V�\( ��/�?���fNO�P�qOZ�R��'%��;����g� ��7@0@�|H��>�� 0D��L>��h��M&�
'lRbhT� �DX�<Y7
Q�J��ʙ������Qj~�(*��|�H>����v%��S-��*EjH&fiY4@��?���?���w���O��Ds>�f�XBM4�*��&B��(C�V�h�Du	�CW�u�#4���������D��),|���?��E+EC�����i��_���1��kMt��êB�OH���ߙGOqOr}i��C"M6eQGgԫb�N�rdE�F�r@3�O����{� ��uˎ�t���z�"O����+�-<zf�r��ɳ{�E C�D̦'��J���Mk��?��闈A�޸�F�Z�[u��O��?��6��p���?y�O� @ /iP���@�P�~]�v��Jކd��T|�h��ʴRB�	w��M�'��l1�4J�����e%�q�Kݕq�y�r�:mA�7�ٲ
����l�' ����l�'a�|8C��"��Ĩ�_�:��Y�'�f��&��;P6��4'Kh0��'J�7��[LВ���9A[�� �#dH8�Oɨ�eG�m��ʟl�Oۚ	)�'R�A�FBH(E
@�Q�)(hNh���'D�aLm�rY�c ��<:����D(ss�L����I �^$�3aޔpǼ�H���1S/��n�q C�P�Μ� 'TW�h����b��4'p��!_��@���K�XYZ���P���'�n����?iL~�L~r�B�� �6�3c��)X��mqC��k̓�?ϓ[�Y3��2mVabaʛS	p,k��4�2�EzR�Ώ5�xh�ᛌFM�es��90��6ʹ<���Н�����?����?��Ӽ;��3r�[J��k�̌C�y�2�hQ bS �ʔC�5hdV��1-�Y̧Z
�m���p����C1~������ٓD΀�MJ��"�&��<H��
�>I���>U)��>K&��1T<�R�B@-/�  A���n$*�l������	J�O��3�$� W�`Un�h$���f���!���=G 	FD�[�d��&,��A�I�HO�i�O���>` �J� N�;@���8��eKA���8���?y���?�ĺ�,��O���uW�]s#�ͪv���ʎ�0��E+���:�~cԈU+:�0�	C��Eq ]� �	�:ވ\YQ叝Jk�x�P�������2k&\�@� 	�a�bɗ8P@\YP�	��Ѣ��Ѽm|\x�\jt8t�ޗ��,>�O^����9�xa!�,�K� iÂ"O����
u�h,@�Z�e�Q+��$�Ϧ&��[4�Y��M{���?��)N�j���kVCI-'����?)��8A��*���?A�O�$����֕��#���d��M��e��Lۑ��R��|�4�6�D���f�?>f�F<j���9V�#xy#B�e��ҰkIZ%"�;����ֺ� a���O$�(�K��	P�kц\�yrF�⧍%D�����X�C�F�1c!�2Y#t�7�!�8(ܴqT.��cX~0(b�N�+zZ�YO>i`�8p[���'�P>!q1gS��$(�H��z� �� p�������	63���H�긙!Bn'I��"�);-�H$�O����i�w�5��HnH��ZL��!�ߑ5�Nܲ4,S!Ok�1"��̧�عP#�?�!�G�{kxh��Oў_[^��!�.}�G���?�7�|���l��9A�ҐnfD �a�9�yb��Y�|e���˛S��s��;�0<��	0pmF)��<}�2��T�A0� A�4�?����?	��Z$>�ȹ
��?Y���?�{�? Xx�S��$B&��
�3�f���%������P�H	�5���΂b�4���>8rqO���F�'_��@4��
=<���L�:�:-�"d9���:���L>� "ϵE6�9�N��k��l�Ga�T�<ad��6+H�8E�۸%������R~�e7�S�O��U���25�	�G��gܰ����3-U�9��'d2�'��t�U��۟�'E�l���I�a�n�Ђ��3�A*�Z�,����i̒��BPFW���O<H�cW� ��0yB���OO�Ł��Uv=ѨF�7C���ğ�O��?�,=:�ԭ��L /������"�����?����o�`�g+D�y5L��m�J�<��D�6��TB�0�fj�́H̓OP�OxE��QԦ��Iܟ8�F��
+H��q�H�0�,��̟P��w��џHͧ+J�x��3�����޿B�|��S6]<��ʱ�вUI�x�Ҹu��a1C�	�{��	RR���V5���\!e[���;�`��I(�M���iZ�Ő1�l��`m�+Ɩe�5D0P�I���?E���H;\��L�15.n��E�[��x�@xӚL��?m��� �EW�N�MX$>ON˓|6�`'�iJ��'}��F��	��]
�@]pZ¡"c��o)�u�������1Vީq����>�ޝr����i�|
dh��2@��ôhR#P�o�_ ��<��8N��]�U.J��c?���n
�hň���{x	���4}ReQ��?��f�O|�O�8%rm�)�e{Q�̷r:>�B�y"�'.�y2Gy�
����9��f�@#`"?��ij6�#��J���M{�В"���2�Ճ9{�m��������Ԣκ�&9���H�I���ݘNqԙ��'"�tx@a�S�t8���<y�e^Tx����ág��t�'-~���S�'�I�����d�2��b��k���kч$�l%������Oq��'�Ȕ�s�
?h (;�L�Z���'B��� c�VMCV`�Or��)�O�PEz��		�n����i��,mq�‚���G����$�O��d�O�����?�������L^�!򮈌$�b��J+ �k
�'�X��6C���";'��%�
+�x���6��uX���U+F�{�h�!���B�W?a��.@v������V��q����yr���8�
L۰O���#�BT��'c�\p�M^�M3��?A�
`Ht�"!ƠcX��A�����?��qfp9b��?ɛO��2����=yHY�&�6K�0Ҁ�]_�hل�I�L�����	"pp칢�N�@P�h:p�$O��1��'� O2+�(Դ*~
�I�]�RS6���"O$��"�G� �1�%R�ICO�yo�1̼��2}�j\"�Lë7=b�d@��.����O�˧ynX��Ш͒'N�:M�*2��X�\��i���?Q4�^�$VPո��X21�tY��T�|��n�cҁ���K$���m8(@	�����ɍl������1Ŋ�K��F�B�~
�#</�Y*��@2�����Ze���d/R-�B�D�t�O8,���^sr����f���O���,G-I^F���.�"L�w�'Ɣ"=��U���<sC������9	� �i�B�'�r"�	�*��a�'�2�'7B%l��Z�nxqbb͇t���
٪2~:�󀗌�?q���� /��|&�ԩ5$X4pJ�5k�$���RŊ��ic�r���(�?y�͔2U���>�O�{�H�("�T�6�BB��{�ɗJ���|'�2Tz5��$t Y�wjǆ�y�r�d��,jtf��i�����W���T�|R�(p��Ӣm�d�����K�=���mМ+�"�'2�'d��������|0!
�*�^�xQkؕ>n1Kң�g���	���  �������7J8�ck�D<�@ ��L9��Q�2�;�Af����	>��?�V�ԌpX8�� �ƣR
ă�+�H�<��札��a�E�{���`ǥA�ea{L��i *5z!�W���q�f��y""��vR�S�cڜa�~`�P�X:�yB�	���AL$W'��; $�5�yr"��;�2xaѢ�+G��됆޵�y��9�T8 @�D$��.��yA$X���f[��8�{%@�$�y��?T����&�^�<��Y�$��y
� `�qN՗0��F!�[����"OH��fO�yd����A!�"O��#mW$g����'2/yZt"Ob��$$L+4�X���N�:|q"O�ڤn�]��@ׄ^>L�Ve��"Oh�%O7qE�y�t�t��5�"O`��[�Jc��At�H �H��"O&��Ӊ׻j���-�<�ui�"O�8ꂅP��:I�)·+��I�"Op���.D��St�"H�<�T"O��P�Pi��':�����"O0����t���V7�v�x�"O�L�A�D� �~�c/�m�H�"O�ZB��=����`������P"O��b�o&Vm�<:�R$r��t��"O��r CU�	r���!LK��Ӆ"O�pG�?p�xa9A�?]�"O�47�Q<X���	-0>��D"O����B_źt�Q�.e5۳"O�������D.l��e�5cT"O�$����m�WaO�����"O��ÑTU�!�?����"O�����0	mr��"��4�l��4"O*�2Qɞ0g[.As'�j����"O8�P��=PJ�Y6G��j�6!@�"O�)�����+�\�iNR�Թ��"O�H#��ɔ��gΩ&|x�s"O�A`�'�%?�%�D=ae�8w"O �Qf�м	�9����D�*��' �Sb��QhR飂��~#|mq�X�Gn|��'�������l�fŹ�G�3Q<����ĕ �e�0#�}�'_�K��2�t�ϑ�y+ʜ��I6O��ֹiL�YU��2|�,Tȹ�ˁ�<`�B�߾��3��|B�o����_ y���	�O���ݞT��I-O�pj�۝,_>13#�ۉ�
�{پ}`bN��S�����S6��xExb@�6,�sb�(}`Z��P��M���ң�Nma�� �P��I2����Ð+�z��5i	�5�Z$�U��9p�x���7���'~�q჋U ^�����BNh`��(�Ok�?ku��caRc�h�b�V D��>����a��Fk��|V�U�(��)��8�A	�)P��I��3�0<��Α.
pN�8SF�OD�@��ʴ1��`k��/�d���k=/%�?���u���a��Ŋ<Ta��BN���	"C��|�wF_0@�L�S� 
�<�' F�:R��!|x@`�B�Or��	�O(�F� \�B+�	)4�y���T�\h0�i�h�1%�VBv!��+�0<)E��6��D+֯F��!��'%h��'1~6ͨ<���ċ�Ylm1�+��S��*lŧ��9�!�''�QȪ�p�4 r��O"�zź�étɈ��$�-@�N�IB�'@�\�2!:	�d,���`}Z!��H��  s�Ô0 h$U��l�.K��'瀤�P�֨GD�{U�"x�,	�J<I�2O�X���4����X�U�� .?qD��	��P*R���Ua��@1$���E�Z�A%"��e�I5(��	�W�t́�C�(��u ��I�9x�{aA�<h��q��`O'�y��'<ʵ�aW�Z�Mig��'w�����L[�'�ў�];H�=Ңß�V<ݻb�C�K�L�ۓ;�lt*�kٵI>�x�-�ykf&c���(�h5X r��Ř�Ƹ'��^w^����țs�J5�E��5���h��"��T�|ñ��/��Op-z 뛌c�d��e�~��u�ˁU$ȻB�f�.�b�ŀ��~"E�:��1Ys!m��|r���
G�d\Fx�I�q�b�@��#.~�Ə�
x�S#�AT���i�����g��ɱi"B0���N�;J�	�.Y�-f��"*�
���'�4�O����%`{z���^}��%	x}��4�?��LHQ�@ɊO~��H@�5&'%Q�]Sq�F�<#��R�Y�-p����^�a���^3
"Y10�,)}t�J��UDh�FEO9g�z���C��?A��V�.\�24�i�t�H��E�|��M^˼c�V�n�Y�K�	���׮J�'m��b�F"FQn�ϓIa�����A˼8e�O Д��T?Z�4q�ȃ16~5�	]	~H��QA'<9Fx��gs�D2ADۓ0ؤ2��Ҝp�{2�[SĴ<�'�-֧u�Dڡo�X�1��ʬeL����VDY¬چq�xѫ@�v�й+�cU����i,�O&���ո8�Ѐؔ��~@�ԑ�mB	��IX�� BTK�ie�DbO?���4,�k,:� ��b "� >�8��� 7��wN�p=�d�-eG���y1 �3m0��c�W(.����%c��1��jy¨�"��k̟Bp;��A'����Oxxi���VI`�Kfǋ{�x�d��=z�����O`�Ib��HS�-$$XA�+L�vP�@q.��M��`
;���Q��D�;.I� ���8�"��&��XJ&-�em����R�E6�T�m��$R��Y�nM[�(�I5oQ���?Q��^�J�"��i�,J� ��g���Cc藴l!�T��Bт$�z�!�t~H��'�`y�en[�A`rtj��En�
a0��'Yf�I�WŸE(���8�db>7��?�xv�0o�3B�FNP	D�[�'�a{�@�)jhy�Zc��X�D�H>����6T�9 ����(�d(��#?qD�O�����E��u��y���ý)��-�(Z���c9�t�v-9 `��;��0�'-��?h����c�Y�]R�$�P�f|���'���'��1���0���4;�1K©>}�i͜ix�C��
������8P��[��׍q�<��O���uߴ=�Z�I�T��(�!��>��P�5���?bА0$"ݫB����GS�Y�')������deZ��%��Bz��2��}S���'w�7�0sCM'��3?a��(n\�ܨ�.O�ht10��C%v�X���IA:������D��g�0x�B���*V���QANE
=��1
O<���,��
V��Iu�-k%�41(�ɗ�H�[��	)Y��-i!�R�*��i�@�'�{��F�p�H�cɤ �����ِ��$�O�`�5��݊i�\�r-������95��Mdk�) ��#m�, �.�QGb�46&� ���~R�Ȕ��L>�P��3{G�,z��Â/(�c��$�(9�s�؂g�<-�����	�7hV�Rċ�{����%�?p���{�n����$ϖoi�i���.�s�1bǍV��ij�X<l�ȔZ�"�O��+�%l�p��GGq�[�4�Q)���@�/O�M���WŦ5z��~�gT��`�O�$Qz�$��7���5Aד`r��0bc�'#�<C�C�;)������Yy�v��O2]�A)���PVk+U"��@�'�5Y�0�U�iJj�$�����'28��e)�<��,��nϔ
6�������w'ݲ<o�M�d+P�:�8��S���yg-X�ns(i ���<�
��J1�?�2��A�����'��zg-X�	xr�ڋ4M��1垈7Vb���SV^�k�m��<�5=��y�BV�tx6x
�3`���%;��>)�[6�R�H��Y7D���p�ʃ�@����ʣl-�tAp0O<�`Á�Zk�=��ڟp�a)O��/g����CB�l�*|����A+ΥDy��L�o箴��KR�l*}�����?���+�R��'�%1��l2��ک� �!ŜO�]l����d`�$N!��+����!� ��Q�Ġ�T4Y��FI-=������	�:�BAHc��l:�짿�P�Ĳy+�,�p��	H5�[�,���ۂL�8�ߓ\(x�BvoL�!w��!�L��o&0%ˁ�I�ĉ1_LaH�'w�5vߟ��s��.rj�� îR��� E�C@1a|��	r�����0��C! �ۦjN�=�^���B�c�<p�'���B�O86��\r@g�J}�'�R��"�gƊ��SC�&��9`Ң�O MX0U,FO�)7��6��w�'C�ѳ-��y��t� U 2f^�Y3��-Eo�``p��Jě�`�,O�榡�gy�-�/���4
�_:-@%�N�"l�"&�#�����"t�¡갵i��)��w�@A��B���-���nh�C�z�@k4F͢	��X⢉F�0<	V�N�T%�Sb�%�*��4`�� ,��PC�<� �àA�SR�O�����(3JxJ%͊#~; � ���;��=q�g�\�G�ĿK��QR��f��1VaX�kBL�ٴ��>e� )k�Y�\f���瞑JCJ�'Xd��߸
A|Z�X,n���DzM�l�lp��`�>�pS$�����6��¤@؂1ܭ2�J$�6�5	Y4(��f ��E��+����	=+��R�M�d��S �5X���o�ʼK�4Y��
cd��)�s�9�c蓥�bi�G�L>6~0耱ɟ{>X�'�=$��a��.X����H�8ta��Q0� ���V'`�G�q}b�/E6: y���%k���'E�& �Fb��1o l�"%��jMQ�gB؞�3JS��yw'�Hq�����ܼh��		)�b1��O �M��X�H�|��M�8�H��.���f��& 	���cըg�R#=ɓb���h1�h�D^����b�S}��� �&1���-m��-��FK%�?��c��M��5O�i��	����?� �ЕÖfE:��(`�R3���n�2XҭJcRY�lT�g���S�s�x)�- �(�W�5}�
]ઇ�2�P� �R ;U���@.�x�I(X������#��EF3Xn�Uℊ%}����&0�|��������W8�����	N&4,�5"?�OLiZcT�2�����A23��: �@�x�&���.E/x%�5�L�'�d�gɄ[~Ф������ݩ[����oL�z��qFz�� KR���Ħm��|�3�E�����l�Iz@b�2 �`��˻N�%�8� Bշ71z��	C��|)��6h��3��0�OR B��6MZ;t���Xo��#!�� D%���<���؈� 'n�*p`$d�o�ȉꅅ-2b�F�@���@�^l���Ǉ�,;ʴ`b䘹c�E��.^�'9d�{?�)O��'����l��%��8���H�&��3u�'9R�rӷ���� ����0�k$�g$���ǛK�
A��c�Hr�O�&��6�$��y1�IE�q�Bj�)ّ7�3�+�y�"�=�Tm�PlHr��-hE����I�G?-!)c�xÖ��3�$Ő��0P��5h��}2'O�<IG@�:hV��[wr�'t`� E���.�� �X49���ߴT H�p�m��$�&�H"T}��&�<ɢ�I`}"���s�T�V�].:����V4��$H�6���
#+�rx��*���D���;C��)Y-�x1(K�B.\�KH>9�(J����9
�N�hM?��w��s���&��T��dxO�=�a|�.ӓP�wOҽP?d�a��7u��" JH1O��&(Z{�'��I���Z�h�D�=�ֽ�T�"F�*#>�Dc�1M�æΚ��C� D�<9��Čl��%� X��r�&����'n�$�YY
�I2Hh06ū�OʀH5f�A��}�C�P�W$�ѳv5OVa���4�yAj+�ʁJ1�'y���c��E~.���a�J�y��'�XuC�>�&��0i(O�رEBO����``.awluP 	�=������D/����"]jj\RÀ?[�E��I�
`�w�v�c�GD�,�he��ؗ	8VH�%F�MµJ��;���g��:�,��_�C>ʔ�W��S�'�ͱ�A=A�Qه��_�J���Ol�a4aV�W�e
(£j�XD�	! H��`Ҍ./<=�,@�Ud�-y�q[�l_�Xd�3�ϼV-�lZ.˞��c��8�F�oZ+e����=��R�BĈX&s���v���h0�<�WMM �d`5��..g�ً�۳?U���D�a��y��R5oZ`v�].Љ'^��nP��2ƍg�g}�n��@���W�<iв�"�U�khy
�2NP�o��L8�Ȑ+
h�I��Ȗ
�N0!0nʤ�M�fM�{零�җ��D�Ayb<��3�wm�����,�T����f	�u�
�'�I#���$v���xu3VȏR�XQ��C�1 �l7M�.F�����'3 +@$�)_�r%�[C���	�'���x"�6ZK��ct�	�J���qU���M�Bc����qF�o�\��Z~J��F��)T@���o*!���=��Y�R�y4�xk�ُ{'!��?WH�H�*"`h�L]�t!��+\��c�-ux)W�Q�3!�$4?0�,aP$UDk�eOq;�!�	�!_�����0`�d�N�6�!��
s���JD��{Y�drFF�4m�!�R�Qb
D��a�8�2�E�*b�!��3�`�3*�>��]P#��k�!�d�:F��-Rs^D���%FF�.�!�Dm�081d����JB�	��!�Đ�p�"�cX�:Rm`T���}C!���5>t%Z�g�1�<e03'L�J)!��e&�A��R�P�سfA #!�D	�a�)Sc��$=l|�Cr�R"V�!���6�����J�B2]K#�Z{!�d�2<���[��W�J/�=8�ϐ�ud!�ď �
��,�0p�Ƨ�dj!�$Fg��g�"x
%'Y72`!��TJ���#k@�Q�Jh"��Xv!�d4#��0"��бY��[C���!�d
�0�z���M:6�\e��R�"%!�	�ISttk2kE���5����?!�$\XfI��kG�JqQaß�g(!�$I�k{���!�)=�$�۵;G!�%Pd�'�	@ݮD`Abu�C"O��S��7L�&|z��]�Ol���"OT��®M�Wa���d�F�f�Z�ar"O�i����k��#��7=߰�"Olm!��ư\�Z̹�G2��}��"OR@n�Eb~L`G��r��u*�"O>���A���PUX�%�5fU���"O1�*�	m�8(�#%�/N�����"O�����Jؠ��D�C�pYc�"O�y����3z�Q�#��8M�"OdT���Ů3�0��B�0?���C�"O* �G��}ҕ F�0�t�c"O�H˲A��h�N1���	)J���T"O� �ɢ���T�b�	��hThT"O�D!�$W#
m�$Ifd�B�H�Q"O9�&�ݠB�٘�)�8X��"O�� 7k	(���u�_2E��w"O�D2���j��T8ug$&�y��"OX���	
�~��s)ǬfV�Ñ"O��C�.�}����
�$��"O<�#�!�U��i)�D ��Xa�"Ozy���.%��fE���*(h�"O���D��(���
�c�E�|�{4"O2�Q-�;O�z�y$�?p�l]q�"O1!&�1U�ȹ��ɛ�
�N!�"O��j⭚\b �	�Q�w��bS"OJ�Kcf�	
���q��ɸ�!6"O,m�G#ٹ=��jVE�z^"H@d"O���E� `�"�s`jөb��S"O�BB��1�����ߵ�P{�"O4���B=\�=@0ȅ�C���"O��i�o^VN=:��ܹ���"OL82��Z�M��$�4�ƨ)�@�"O��#�(B�P:td�p���j�"O~p��l�N�Z�jAB"O�P%�.,���ZQ��1*���@�"O�h�cI�\v��a�*ڼ}�sE"OT��W�c���4�8x�)h�"Od����|40���V>r��(A�"O��HF�]�A P��s��(<�`9[T"O�� ��mʵB�6�0��"Otȫ�lK6�"��+��$i�d�"O��pî�
�.�;��LR���"O�@h#�H�p��\X&���t�h�{p"O�%���(֔hⰁ�D�h��"O������S~�Ԑ3 �/�ց��"O�|��G�S5�<C��F�<�F�z�"O�(���E�w܀cQ�4
� T�3"O��䇌�B�Zٙ���`���	d"O"�s��b�d,zR�	%�l}:!"OX�{!E�gE��H߉Y�xm�$"O�]�!�.9�x`[D֝�j:s"OƬS�T3
�<��f�_�P�D��"O��Zի���F��&n<`�Cӻ�y�R�	l~�{F�ӈ:~Ԛ M���yo
�PmV�+Pd�
5��S�eX&�y���0%#�-�qO*yX&�{��Z�yҎA�b���s� �[�L��y�d
X�����g�Jy�E�Ϻ�y�ђrL.p"$fN4�f�1읦��>��O�ٚ" d�$��Bf�5�r"O�mؑ� D(!��Oê,���i_�tE�ܴ5�2���i�)N�M��.Z�N�����?I�F�-�8aqsNW�P.�����M}�<$�����b��h���S���4�չ�B䉾9��T�w��(6Y�"���2H�`l���ƨ>in4�(U7^D�EI4B�!���O8@ P�ǬF���ϙy���6"Ov\�Q��� a��h�K?]H)E"O�����5�رq���>%��@a"O�}�� �Jm��gM�+�d�ab"O�;�P���=�� "{�
��"O�iR�#�$z�R���J?p�9R`"O�S��f�6����X��i2"O���4��
!��q���	H�1"OV1R���{�9�q��6�m.�yR��j�Ĺ�ҠA�BT���[>�y
� ���b�_�m�7ȇ*K��U3�"O�9�`��^N����ǜ9d	8]�"O�� GȌ�s���
Ѡ��~$�P0"Od��!�P>I��O���:���'���U��P��Ģ�$��D��N� z!�dB�D%�(J��ņk٘鸴��#[!�ӋiҮ|w�� 62hQb�òM!�d�/M�޴#��Q�Jx���#P)F�!�dԷJH�hvoX�Q˘�T�T{�!��T�|�j��⌺ZP���?�!�d�v�a��@�9:M��y�-�=�Py�_�)���T�G�R�HIQ�)�>aI����X�Eߢ՛���q�l���3D�(�,��`=��cp@�AH��)s�2D�x�@)���ʲ�x��(1D��p�M	%��B�F�27�hp�B�+D�\h焂� B���m�!a`��T�'D���2�ɔD�*=�Ǳx�>���f'lO2➰�7�вF�YAÐ�"5ʝy�!D��˶HX><�J�U�S+D��I��L"�t���Rτ�*�m�W���w!W39\���	x�0��>�­ك-Z��8iGzB�'��M�T`w_:x��V���i�'� �F�-�HBr��
�Q��'ia���K��� ߕSW��Z�&U��yG�;3jt)ֱ3��|i  \�y��ю$����B��%�f�@0[��y��#u���p�D�RDN.�y����)J�,w��	�+<0�=E��g�`-#��,\[BU@��Q�u5Z��O�=�ң��6� C���_ �'��A�<�,�a��2��=|h��Bx�<1��hJ���0BX��l*Q�CN�<��M�>wr�t[p&D!�h���i�G�<�Њ�P�\B�\�܁��N����'F��K`oR%z[�qj�
9z 0
�'x�qأ ��x�r3Dc3���	�'0r195Lɡ+<�)t*��D��'
�S�كc�����FҼ=����
�'�\1�H��!JqE�ܫ2�0��
�'m�e
�i��ѩ�=T�q)
�'�0A�@a�W`��
��	
&	�D��'�̌R�拙H��T! 	&-2N�3�'����an,4KHX#��(��,���5�S�To25K�-���P�H���
�yrm��n�n�i�!���R���mƱ�y���C��uFW1�>L��jĽ�yr�αV~kG�]
��� �O�O�=�O�<��"����)4�	*���+�'&�;6�>8<%�c/ω$ժiv�)��<�'��n` �M�L�tY;���r�<Q�B6E�ћ@͎�(U� õ�q�<��#]�~�2%����\�0�C�C�<��DA� ��p�P�#�5@�b�I�<it�@�8U�Zr;�mD�G��hO�O�N�+Rd!���`��*�� �'��)��J�NW��3�
�7�`0��/�H��	�Jy<���_�r�d�f�:e��B�IvQ	RA�8:,����`��5��B��>u�]��ʶv�\9��d�9�B�	�&c �Ѐ�&j�DT.܂L(�B�I�����CԅQ;D��G�;c�B�/t�>T{�̳26L�Q4@�q��C�	�!�`@�6  }��b͗&x�C�)� "P � �'( ���E��Xg"OZ��3F�
o�`%��d˽q��9P�O���dP� ��aa�Y�}ꑻed. !���9=�-�g��p.���aČ.Tw!�Q�D���fTU�BIN�!��张P��G�Z$��j�ι
�!�dI5#6�P�$���
�-f��#�S�Ojz��CIB&w�p�p�F����
����*k����Bg�����k��	�yb���L�b�!#
���)�����y(<oY8������@��6�6�y� 08��X�{�yf�����O
"~�˟8h�a��ʛ:gf���%%DF�<1!�ƮU�ݱ�*�:$��ia1K�A�<A6�A��!	��?jJ�Hw([G��@�	T~"�C�r{�蒑�į{���p�Q:�yҪQ)����'�.(~]aA�B/��';�z�旑x�:��5��U\�쐥����>��OZY�uB_ 9;�A���'1��\z�x��*�'֚�����!�8:�� ـ؇��V}��>!E��(������"^A�x�.�z쓛M�˓#�`-I�G]�P?��A�-��ϓp��"~b��_�:"�����_�8u���syB�'a|R�C5��]j� �~`�!«ű�0>�H>A��	�'�x��!*����A̜k�<�FV�Qƌ��)��z�N�(�m�g�<1�%D����$&��Wx	H��Vg�<��Q	���b��?ɋ1O�e�<aI� q�X(����kSr�FcBe�<S��[z�(A��G@���Ō�d�<�bI�In�D ��wcW�Bj�<i�*W2���3�ѭ@�P�0�f�<qd�Z�d��0� @Y�2�B�ʶ��b�<�$��3��1K��k���JQ�X�<i��I�%�ʍ3L;jVx:g,�{�<���!=]��Qs�R% ��g�u�<YwȒ���t	^c�h���p�<i�-C}��A� D�(Z�����g�<	1%q�~x�7�E�'�l]�Ɓ�n�<i� �!jK�E04H��0�6 �e�<�4�e3�ɴ�N���C��J�<Q%�N.���ψ��Uy7�QE�<)�F37R�1A���G��=ɲ�Z�<��[�R~Xa��iI:o�@�0��V�<��팜*��9w \�NF�`f	�T�<q%Y�4�膉��9c��#iHI�<��E�=G@ qã_7H�h��7�	I�<I�JG:b��:�.Μ= ��bBC�<�d���Ax�LITUQf��PH
A�<9Q�8?D�i�g�=89��Dd�<a���w)p���.qk\�W��\�<i�M�P)Y@K��:���Wo�<�ġȈ)�d b�AQ&�	cD�j�<�S�`�j5�ᧂ;P�*�1�Rf�<���G���q@�ڮO��F�d�<q��iε�`���y�4�K�z�<��#۽h�0Q�A��o}f� ��[u�<Q��ǷWe.@�,�Mp���o�<I��j�R��c���U���j�<i�.�8.4�}�b�#-���#A�P�<��k؀G��Q�6�L�gJ�<�q���Њ�Ϙ\�"%2�E�<�P��J�hi��O�m�왷�g�<�g�
�D�l��(��P��Y��AK�<� �|
U)$�0�)�X)V�yH�"Om�A+��UT�A��;J�e��"OVxp�M�ݾs�v$"�T�y�X���Z�b��@�� �ܡ$������q۪�����:���酅�4:܅ȓ,UX �4 ��(6�!ˆ���I���Y�%pd�����Y�B�ȓc�-��U�6��y��D�g�6͇ȓ�, &f@~�����e��T��&$B���:&��z5��yI�E��+�� �"�.Pahy����*/`��ȓ 2u)�OK<*Ҭy"dO�cbB�ɗK�,����H@�Er)� oC�I'�ȑ9Q�M�:rܔ˖F�<;��B䉼{-ʄ���WxC��S�gA1$�B�	�;Z��EQ& o~uiB�߸&�B�ɑ��H��5J>�@;B�ޜp�B�		Ip�����V�E;PݱղB�	�vԑs��_'��i�E@��B�	 4.�0Wʊ$:نq�n�8˔B�	�e�6��UB^3��eխQ��B�ɱ|B�ŁU�J�dh�W�T[�B�	:n �zE̗4J(�XFkH��B�I�O�֕�#M(n��{�d�_%�B�Il^�� ��b� �2eFʠB��jHH�c V9dʼ�� f &B�I�E�~$�w. p^�d�����0B䉲l}R-��&A3|���@�G�-� B�� 8���a�މ4�v�CG�C�.��C�	�6��5�DY:���F ��C��0_ �H�aT�'�&Lq%�W��B�	�r�= ��]�A��\"5#(<�C�	SY;1h�����	�rB�I=_	tHzDF��6eb]kc��#�C�ɶhw�(� �T�T��!E9��C�	7Q�-P��28t6!��I�2��C�	�I&v%� GB�+�$�xr�7�B�I�H��i�h�QbY��i��5jLB�I�+�A�%҄{��:��D�h��C�ɥj�I��KW��H����ƽe��C䉴,�8�x���Jv�a1cY�no�C�	El}b�M]�D�]�Vb�Mk�C�+R*|����M�@���R�jTBjDC�.3M���6	��A!���07�BC�I��rQ��D[�=�e�|�C�	<��dl�q}�i[f¹[�8C䉀e�в��Mд5��K��pC��2�v��*RD@��A���C�I@�l �) 7Q��c�͍�2��B�I��� ��ϙr���%,L�C��C�� "�$�����>*��=Q�.<^"C�I����K �Q�|�I��F�iT�B�	�'Ve��k�9%�UXFo� O��B�	�2`j��8ߴ��C�Z$8C�	�!B���h[�+hƘ�w��:,��C�	/v(���U�P)�ިR���>��B�ɵ���hE�H�,�� �$+�8>�B�ɫ1�9Z�"�5�� ��݇e�B�ɫf�Tmۅ.8����f�>�C�F�h�ըE�L��@��^�0C��4R�^�1�-�cz��˘�Mg�C�=<LB��T�"a6�b#��(�C�IV��l95��p�f��v��y�C�I�pHd)@lY*S����	p��C�)� ,<�G���eT��xJ�"OB�@ѡ(���g� �R�bq"Oh��g֪uN�x��E9W~����"O|�5�ɞX
H�GK*b�0�d"O��C#�˽\��E�K��?w��AD"O(|8F��E(&̉k�X�T��"O�Œ7@ǚGJ���oP.	�@rd"O���Z;Q\�X�ԣ�) ��"O�,C�zG|����=�z)��"O61K0�ڶ4Mش�.��&�"OJ�ao
�-F4�yF��,��"O6e��ꏟK����#�o�����"ON5���дa˕w��"O��uAZ\����jud��"O����&��q�D�pWc�"OV`c�HC�F���$
��N��q�"OVͫΝ�a2�Br���@<���"O6زcfD|�V\�u'�WW��ۗ"Od�C�Y�>��Mأe�:X݄���"O��{�+Õx��$rDA.6¼�)�"O�	A1��~m ��� T�T�1"O���u+_	m:-�1��{O�|
g"OBT��-2Y����k�UR��`�"O�Q@�ė�6uX��Z�2�9s2"ObD�a�F?_��##H+)H���g"Or� f� �[�Ȑ��lX�CF�Z�"O��YKd�Pԑ6��a/�6"Oи��M_6?�I& )]7vEC�"O�Q*dD��_4�-��/I���B"OV�Aǐ�N�<2���$ �"O.���C��y�-"���`:"OV�X�K�#��4� 01�BD��"O2Q[��܊jR\��A��D�9�"O�\� �C� $��0`�-���"O�5��o�?o�mQ @BAl��"Oڈ6��h�&�"N Afp�"O�ݹg�<+�de���Տڈ1�"O��	D�Y=+���6Gòo�ά�"Oj�Ƈ�3)o�;�kJ'���W"OB4r��crjQ���@,b�sS"O��P2a�o_<�÷�_r>��"O��#��՟z���B��ՓX�P`20"ONA!ף�D��A�&E~�Y��"OZQ�c/K�?��l���1z\�,�3"Oxh�U�`!�v�ڹ!��Y�"O 98uE[����IP@��b���@"O6-�fa�.t�Z�����BV"O����CS7U��@h�.!0��tS"O���	*xG<�����;���z6"OxP
1��x�x
d�N��܊�"O2m�Qj �yI.�k�͝�6:`R3"OaaAhC�B���'E|"M�"O
h�/��>��y�IɆT��"Od;��
�1#�T�0�J�?d8YF"O� 숵F��af�9OD@��"O�� 뚸�x�H�āp/��	T"O����1j�2 {��#A6�"Op|Q��%j�h��Q7Hy9@"O^dW�(`$`�B�0�@(`"O���%)�Y_�er�i��I� ���"O^��1�e������#]��k"O��,K�;�N���ץH��X""Ozqq͟�#	�މ,�nxk�"Oz-P�#�Dx6�]a"pX��"O� �k��T����K�B�?vl�"O|*�_��Nx1� эd��3"O�y)֨4"��x�/zS2��&"OZ��&�.8w8cp�RXb�{�"OЩ��c�#`Fm(���,5����"O]h#���^1J��W�Z� a�"O0���d�85��)a���00�	9�"Oxu�wŇP>1��h�D���f"O0�XAn��Bc�!��u0��"O���A>H_�иtc��pd0%��"O:p؇cM6%�V�Zu��O��yr+Kv��"�$φā$�K��yR�?ZQ˃�������&/�-�y�E*e�n!���p��5�Ul��y��� ��MǥV'E��E�y(ŭ� MK��Y�CD��4�6�yb�(�!��ɜ5:/����J�yb�4�@CF-C�	I`HJPa��y�ꉩR$yy���y��٤�T-�y�E��)ڜh�� ��D�	!���y���S�1TNO�s¤:pe�y��fI~m����f^du���)�y"�R%��e���6���Ǣ
�y�N΂&� Q��.&�|��N���y��אE��:ҥ]�HLneq���y'Q!�����
Q�����'Q�y���&i�@����F�D9@F�#�y%�/��9s$�8qT%�I�1�yb)
3�議�$�FjԹ���߶�y��;q] ��w�э7_����y�C��(T��r��� �zpQ��[��yRD�p X��I�e(����\��yRϕ�D�R=k��^j�5���y���l �P��aZ+��.ޖ�y���>X�TӠNCZ����y�*�f�fY���E ���>�y��-+�XR1ô6��x���_��y��"{<�B��]�e�NQ�GG���yr鞽]a��@��2c܄!f��y��F��x@P�E?/=~�B�&G)�yRLC�K�P�[5�ݑ.HT�;G�9�y�$�N}�[��΀8���8wIH��yR#�M�D��G�31�p�g�3�yR_;32������ iH��a�ި�y��I2z䀢,�r���QD��yH��3H�9��Z�m�n��0�2�yr��3(R%Ak҅vf�) ��y2M��d ��v���l��0Bp�P��y�cH�
�e��%vc����9�yb��G�.��B!J�<a6��C����y�d PU~1Z%F	�-�85�"��y�i1�MH���-�5qR(>�yBFN�.Htcr�J��`�y��"�r�&g��}��d����yB��&6]V4@�'	nC�i���y�7"�v�hᭅ�tӀA���#�y�g�4{�)�HD(l�-*3ˁ;�yBH�Y/�a��C�o�^5�⁀��y��Cbf]b�dF*k\
#rC��y"*�E���r���;P��?�yb��C��+���|�l̡�`Ղ�yR��&���EzкE9���y�X�R��P�3�N,K�g��y"O�3���A�f.�"���7�y
� 4�SL�''�����%E��ة&"Op�1�kA5��mI��E�֡CP"O�� �@�T�2���C̗;��=�T"O�@它!	,��{��G�0v��"O� [(�b
4��F	)�Q:6"O�*Do٣8�@�+��7r��p�"O�x	e���w�P��䃿^�0��$"O�TBԅF���yz��ѥJ�t�"O�� w�V<s������W��*�5"O���+�LO��y� ��n,]P�"O�XKT�,�����(Kv�,�6"O��3�Nͯ'D��XTk�|V��"O�`�OP�(�H �*�6@OP� "O���1g)BG�E�`�C���T"O8���� !�h��g�>��&"O�����y�b��á"Od|S���&N����$K/CR���"O>,R��)�&Q#�Ѹ�aj�"O���	�0��K�k�2���R"O��UhAR&H����Վ.ǐ I"O�4�(��`��8���Y��, 0"O���&��$3~�p�*	�{��:�"O�u8bgD�ᠨ�e�|^�	"O��)�h��!xhp!���`a"O�M0��y1dM#�E� -�Գ�"O�<�W�	G(v������0z��24"Oj��#/�e|%1��M4��T��"O�x�gM8i���I�o)Rjh݈�"O@p��! �M����ѱR`��a"O��9��\����eh�G�e� "OZAcZ4}O�� hכ>P�X�"O.iJ�l NM\�������aT"O�d���5|� 0s�)GA�USR"O�ss��F���G��pH�w"OzyЬ˾ { �aB';.�f�8�"O��Y�O��bn�Z�
����4"O`�(OX8x���O,/��u��"O��2U�˽��C��|z!�Q"O�UӤ�:1�r�R�BE�Z
ذQ"O���� �GdL!�!��
�G>�yr��a#��)�!������ ���y�I��;V�!��D��5�U��
��y�I�����	�VX�c	��yr�[���J"ϵ�B�jc�ρ�y�o'+�F�y����5C䤎?�yb��h~���"�!����t�N �y��חV����bI߮k�����͏�yb̏'g���פ��_��%��\2�Py��]�9�&A+0	r&Y�N�h�<!���e��U�z��k�EJ�<���;!����l�*O�u�E��E�<�`�-*vy"���r���B�Wf�<7�RF�x��J	�bذR/�F�<y�
�Mz��v/��J%��P�OQX�<q����:���2Ⴠ-��]>�B�#3�&��� �*��y�ъƛ �rB�ɪz�\Z$��.dO�Q�0c��a�jB�I.5�4��1
�\��y�
ޠ�&B�+2���7(G�@2�T[<7WB�;Y�΍xQ�5H�LB��N�C�ɓ5��LQ6b��?06���`�� ^�B��5�.�R-�3]�@}I"��y۞B�	�?�n���A��u��l@�
�2m2�B䉐�H=��a��&�t���,{QDB�)� �z���@�6x���/O/Z�9�"O�\(�.H�G,`-��T���"Oj�[�h_"/����W��$���˵"O�(El͒b��t����a8��p"Or�Є\�y\25r�����ţ�"O6��#H̘��uj'y��'"O��㰭�y�0\�%�.O2X��"Oz��-�Y����(+>��s"O��U�\��FQ���Բ7o����"O�P�c�U=&"��p�BU9����"O����]�gZ�'-�Q��3�"O$` C[zø���+?� ���"O���a�>p��Q��9=�n|""O$`@���A��{�IfAxd"O�H00��/�2�!UOP�@ �V"Oz�K�D�e�ā��+�X��"O��aЉϭcˤ�X��O5~�!�"Oִ ��P!V��(�����Tz7"O�P�OŒ&OЀP�O�::8�'"O:�P�+�.`W�Qq�ˁ񖅫�"OP+�*��:k��)�0'�ر
V"O ��$��dCF#�*w��MɱkԖ�y�A�AQ(X��=i����*�y���!R�����&P��p"���y¯�6�|4�c �<9�5+@&3�yB�[	u����dk&0��\��]��y��J�=������',���` �=�y�!�. 0#��\1�j4k����yrh,7�@�Qn�?.�h�@G���y"�׊_L�i�@H�o�BD{p
J��y�I�-��Y�0�$4bVL�Hؤ�y�a�Y��q!���$g�1!g,���y��N�k |@��^�R3h�ض�E=�y�nM�h�ׅN3Myz�x����y"(V�n�N�8vMQL�Q���y�Γ=~S�"7�C��Z���;�y(N�
�l2�# �.��,p��	��y�N�_��􋳪�0��ၣ���yr$�+/w�z�Aӏ* $��1�y'�%E)z���d��U��P�aB>�y�ыB,�5p%��N(���̟��y�iΉz� �x�n�8L���3�5�yBiʂI��Cao1*P �0@(���y�ݘ�Ա�(E�+�@h(��¾�y-I�)���b�'V�"=�]�f���y�e�x��}�����sܴ�����y��F2E��$�ȴ�J}*���yRg� �X�s�΂u�@ �h��y�#ҋQ�ށ�^�Ba�kތ�y"���*]#-׏\)*���^�yB'�P�����e�dYi4F��y�(ӽk���j�6	D�����y"��*iZ�����U���{@�3�y2�[�-��@C���O��D���y��ߛ��)K�+I�@���0GL��y��V�! �d�8�"�I*���y�#P8}���ڟ2Hr�Ӕiߧ�y���St�B�"z���:���y�n] � 
��W�v�ٱ#�H��yRG	�N�2��j��i:s"
 �yR
]�si^�X1툜0�,���<�y�j�((�9��*S��*��Ē4�y����*�(�ʄA�E��IkQ틅�yRe�+{�p�T���CO��$��?�y
� .8"b5��D��G.X����0"O�8��bV�]���Pf��$-���jW"O�E�х99�Y��L��j�"O�$��q!pI�e�3�TT"O
䀓Æ�:��z`K�&o�Uc�"Oh|	Ռ�?�D�PԫX�`��:V"O�`��퐃R�b-3�>�$��g"O��B$ăo��k��{�p�"O*)�u��'�$鷥Z�-�ڀs�"O��(��>��H�����3¶��"O(��O:��4j'�Ϋ	 ���"O��K4���^�d�	҆��Q���"O�Q
p�F'�e���PQ����"OaA�]�2 +���UH��c�"Oth�
�42F CbB�(7��7"O�5'�ݝ8��9��\�q͖�
�"O�ebw��;;r��R�
�\���"O�}B��!*%�2�L�|�@"O^\3E�A�G�S�V�) ���E"O�
���+=:�P!h�� lӢ"Oj8��U�bX�p��L:b����"O����r�<9q.Ëy�>��1"O�1���+/��b&Ga�(9p�"OFx��-�+Z��,�	Ԯ\�t!Q#"O��82H1d���1*�*b�Li�"O���[y/��&IS9|�>y�W�q�<��$ZQ�z��$^�),��+p�<q��X	P�yنoܫX?�LR�k�<���3GL\`C�&����c� _�<q��ku2�N�
^�ju�W�<�ԄN�t���j�MևsHƙ:��<T��['D�P�v�js���%�D�b��;D�40��>;<�RE ?>}&����7D�DxE&�@��C��\3�"y�$�4D�l*"��x�<�d���#ҫ0D�P�댁�&�kcةz�N���i+D��!S U�7�zu�ҌS�C��ĈT%D�(�5"^�r�KV��#=}�4s�a$D��*J�X��83��T�^�Л5�/D�(��� oh����h�v�~�R��-D���d��FNм����D7�q�6D���Ɓ�T��4K`�4Z]�-�i D�DaS�S�'����ں-0�i��&?D�\����+CJm���O��Q K;D����mL�l�ɐ�oI+K� ܀m7D��@7��$��l`���.\��%�#6D�`���K?�i��Č~��)�bi5D��B�K�0��#�@���ap�3D��qF��8!p���eZ%| �$pb�=D��#%O�32�l��bW�y��405m8D�h�㖟$���1'�'���ʗ�2D��G�S+;���1���2}�f�k��1D����i��5��5Q�K�HM�f';D���dM�iؐ<�ԣ�A��9D��"�X�v�z���!q��}z��:D�p�矏5�̩��B�ɳ %D�H@0�ՓSϲ���(f8�@��&D��󵏓�H�,)�
��:/&��'(D��� sJe#�f�eY��q�%D��ks�Ӱ�^q���
@.�L� �$D��P	�a����ɗ61����!D�,z�h�`�|��TE +��%:D�H3��׍(b4�6�@:0W|Hk4D�@��ѯq~��`�]�UL���2D�� ��i�(H�N�0��թ\<4A"OhB���:b?&i�"�8m�(""O>�;�
lJ1G��&��"O��P�I�m�\���"��{�"O�\y�Mڬ.R\�葳3x�R "O4x�C�F����I�,D&a�@"O�\�שކd�y���S�4UnD�T"O� ��N�	T�^Ij�枬UHi�c"O^�a���	p���*��$��"O��c�)ۗE�h�)�揊[w^�{�"O�HѲ�!��Pg�]"&^F��$"O8X!vt���0IV?-|XL2�"O( �b��6t������	/wv�ȧ"O`%1�C�B�>1��� v����"O�����S�θ�M�Xn8��"O` �ao��_�M�3+�>qG�=8�"OR���+4o��$��<u���Q"OT��g'�4:]��*�1lv>D��"O^cc�^*xДItj��7�����"OF� Dg��a���i�b�q��"Oȵ�S�ޓ��� �!�Z݋D"O��c%M�l![��L���c"O0} Q��g�d�����dZ��Zc"O�,���W�+��t�SN[�JT�["O��3�V@�	-K���ф"O��'�̧Knb�ƍ�z��|��"O�|�P���B7��:@���rậ��"O���b�5#�ސ��=>��-�q"O��!��[�Xwڐ�%)Z�O�B�`�"OD|� ��	��I�t(P�8�d v"O`�Gi�-H���hO�l�q�"O�% @JO���]q%H�qr�B�"O� +7!��E�"��fX�k5�ȗ"OPE���B ;�.[+R��h�T"O�����8E��T:v���n��Hs�"Ohݰ�)�)!Nl!@a/�MxP2"OƉ(�� QM����.^�Th���"O`�@�t�4z4	$1U�T��"Oi�s�ܻmc��pK�8��@j�"OR8��͊=R���;]h��"O�`����/4�	�)"x�1��	O�O<B�P1��Eh �B�'�� n���'��<���6��m�sB҃�~5p�'.�\�1+D�Zւ���N�6 f���'�ht � �M6���1��"�H$��'��d�Sn��ȂV2�ʉ�a��g�<�'�/ �тTfC)fPDq���Vc�<�����6X>d!���D��}H�-�^�<y`g��`����׌<\����-t�<��(1��}�Gˀ$C���!
n�<y�Y�;��`���|�^(`țe�<�d+@q(�A`@�9vUpS�I�<Y��H ���"��e4�ܻ�j�C�<9��C���I
򎞸_G� ��$�A�<A��X�>��`�"/��=����}�<��ˍ}2�4�1�ԟ��S � p�<��.�Y�������J���.�g�<�`M[5TZu�ʀ�"q+com�<y���"&�*7��� E�h�<)�jA�d��"V-]�v���+A&�J�<��.*i���ԩRI�?36B䉠F�|pN�:��Xv쒉z� B��=9���!���m7�8{�m0=?�C�I(:ͨ�f�V��3ya�B�)� ~\P7�V;B�$�r�;V��L��"O>��w�	�{�ڤr#�F2R�Z19�"On�(v�ǅ`K$������A"OV(RFB����<� ���q��"O����ܵ?��2��F�4N6{�"O��ÂnΝ	d�9�F,��:�"O��b�/�Q�Z�cr#J�l��x�2"O����a�g��볡�$m��� "O2�P��L�CS�ER5 Q�@׼�x"OB��v�.4��˕I��=�:\��"O�aC@הPX������)��yV"O����.�'xfl2f��@����"O�14� �5ȠpP��0H�@��R"O�a��@�C�AH���r���"O�L"���9�\U���܈w��3�"O�qB3�49����Q�{>�Y2 "Oh(Ja(�~���s�W�T֡Z"O�y{�*ڎ/�
trd
��dY���"Obl�����I�6aB���/��x�R"O���I�vm�$	e� u��qP�"O2(�RH����:>�$���"O�2Wj��JO�����4��`1"O�$pD��#����lK������"O�U�fI8�,'ˈ�k��Q��"O�]�3NR�z�xa棈�|�,a �"OHu�4I]T�ԠJ�?���"OΨ�j��K��8(�J\d��r�"Oy�'�P�s4eJBϋ�H̀�4"O��9!,�+�U���Bi�C"O���m�fx�<r�n�M�%�u"O�<t�!��a��v�  !"O�p�׆Q�1���4��5)U�"�!�dH�Ul����� W�5qBd�213!�da�i���W�"��(��Z"s!!�$�7��=��)I5��� QoD-H
!�F3`�����2y6Fd�5.C/L�!�DL-gꥰ&�G�M3���&�S,>!��H�9W�`ؠՂ(��pj��!�dR30��Ъ3�ѩWS���HКd!�dx孑�g���y���ɟ8�)��gB��;"�WZ*�v���7�\<�ȓIҶ�I�e�9��q��>`� �ȓo�U�0�O9B�������V����C����!/�8��- ��3����C�J+��>�`t�S�I�]�Ʌȓ
�r(k奒�\k&��w��9�&���9�B1{ӯ�3����w��3IR��ȓv�4���GL/!�D�i��,��Q��7��E�U�A��(���p��@���2�F;���BPFԇȓrl���I��:a8h(�#�DjH��h�����@,�����#����l($9�'n���D�s���΀��7�Z�hנ�3Lb8;�GO��ņȓ���*���T��mZ/��@�z���W��:gT,"*�ABf�ő�m��<v�1����Y���)֧RZ�ZH��/����/(5�4+P̒�����e�FM��G(TM��NӯC�B1���h�ɧ��+T�&t2�A)�&P�ȓS�*!��N�kW�����X��4$I#��RpY[�/STS����af�H�$��,2�vcw
�E��h��F@�![�M��,d:V�u5�y��S�?  u+�E���A�Ǎ�(b��q��"OHE1�o���(l4�ɓ[�<�I�"O�QP���t�8x8�ϱ;涅"Ofh1�D_�i0D���L6DɊ�	�"O��0`��X�������l�����"O��Zr&ľ煝�'�v8�!AB�en!�d��K���q�T0q�N��eI�6Sk!�Ć>^D�Ö�Έ>�,�r�(�� -!򤁺2��F�|��4�7�]0!�D��N��S�&�3u�F�" �ֳh�!�D\K�D	bHS=u�h����֮ �!��[���Q������UZ0	�|U!�d��s�������}�$�'I� ^U!�$җS�,�"��h�Q!�$Xh�ht�Gn��TZ�'V7!�DC6j|-:"�7��H���)!򄄷u�Ըs/&JΖ��e��(T�!��'8k�#�J��z�֩G?!����̹r�X���p�4�N�"!��;t!Y�ATb��D���'<!��C�j��@8�튓f�JM��i G�!�P�I4ـ�&�3, �ȧ�!���-<
�H�/�P�i�FG��g�!���M�Hk�H�/6�x�$��,b!��ʰCnf����H�	��H+d=.R!�L�NN^�a4�RU�"�i�54!�ȑj�R�T>x��h�5�U)_$!��7W(,I����J�^����Og!�.ۚ�Kf�.c�`5ys�M�&_!�U�)�L��I��=8���,f!�׭S�����I�n��I��]K!�d\�?��`�lX�I�:��߮nc!��W,1:�9� *�8��E�,jH!��ϻG���P����,��m�.!򄎺u�<8�f��]�Dmi"��!�D*A�8�+6"�]��`��Z�]!�D����@sVb_�V�<�#��:|�!�d�:;hT�ckէgC�+׍Л�!�D�&;�l��ʽuY�2�� ,
�!�dη%\��2ᦂ�t�x�p3d�[�!��F8E��uB����"���"��[�!�ܿ��yx����Km���u�H�'�!��1+Ϻ@��� }�Uap��W�!�҃[�=��₠_n9yTg�U!����"$R.ܴSup����T�!�$�s�8�;4+Pz9ȹY�Þ�A<!�0/N�㓨Z�V+���O�O�!�$����!��ہhX�c��2�!���%?�\#��k�P�LY [�!�D�O2v@2���'��"f�*�!�d�3A��(��	��2]�$�7�!�Dõ=�!C���.E����IE��!��H;'=�t�[��̿�!���82����(�+i�
��密�:�!��0���Hev�|JFO
�\�x`��ox\A�.]�n�}���+�"���N�|,K�D�y�U�I*}E�,��/�R�Rf �\x�$�D̈���ن��)���l�����H�,�ȓ{(tiu&@���H�0��#;T-��<.��)".l|���
�AX��E���c�^�7�!���i�&P�ȓ7���6��.V`=@�G�XL歄�lH���Y�G�*X@ǩ u�L��S�? ��3o�'@ް�Tn�S���A"O}˴�v���MH�C�X*�"O�� ٠hm!m����"O�]ٗ&K'Ȕt���ҋI��y�"Oz�Sba"MD:�P�AC%>�2�"O4������D����ӡ#�F0��"O�5S��&�X��-�V����"O�Ęfd͛h��awj�r���C1"O���ۿ�����bz��SA"O�#���MDA��Lz��H�"O�m�G��4eq�FE�0s"��5"O��C��C�d�r���!��"O����� E�2����]5EE�u�3"Op(�߼%��Mx�cW=E;b"O��b��G #J
� ܻa1 ]��"Oj�7�A3L�@-0U��Kn�@w"On}9G�4��b�K�=��PX�"Oz��C��B,:WM
�t��*�"O��ǭ��=��EǢe ���"O��CF�-��$ �	ٛuQ"���"O(h��X7�@��7UB���"O�T�'M�$&�(�`��'W=����"Ob�8#�J�
(��tሼ;ٺ�"O4YǩL��&YCcƸt�����"O�X!��U�2&F���.\����"O0���i^����G-+�Xh�Q"O �p��F�b��m��O�-���#"O��R�$T;Du�D�
*6�(��$"OZ9hs�]�z�0-	��4R�X� t"O61�D��$S����'m�6i��$��"O�M ΍�����8F��Ce D���pC̸m�F����Nr]�ť*D���橅�,N\{�,G�fv~pS �+D�܃" .P�� 3j��|��a)D�0���ş:Sv�pELBN�&��C�%D��`�Twp�$��
U�4B���yBF�M�l�	���x������y�ͰVS>f�͊����y2 �28`h��\:b\�c�*�y�]l���Y�f�}�V�h��� �y���#Y���8BR!t)ҭ�")���y�aɫ`� =fh�Cߞ������y2a�"�$���:"y�Y��y�CW�4
�d��I��(���y"f�7����V�m(�pA�V�y�8_D��v��d��y��߿�yl���~�CmM�uQ�@��l��yr�ܪw����m�(}��8���y��ܴ����W�o�>�8��	�y,�FD̻a�Ƥb�"A�`�	$�y�-�����5(E0fQ����j��y2D�h
j±�^�cW����m5�y��
o�֤�5ꓵE�|]0'�-�y��'e��(i��ԭ����e��yRʘ2H$$4̎;A"9c�N��y� R#qzp�"u�F����C����yr���00T�{��T�)�+�yES�@���ٴO�3�����FJ��y��1�Ĵ�ȓ~L��'#݆�y����0�45sf`���Ҋ�yb S+�٩p���rs$@�v)5�y�@?�)�
� �0ia�n��y�,U�05Q���z1�������y"�@!dt�tFZ&k=>�
��^��y
� ZTZ3ѤY8�k���$����"O�E�u�f�	�@L�Tʊ�`�"On����X	y�&psա����C"O�q�uK��XR��S� ��:$�p�"O�2G��&�^�ہ$J��
B"O������A�DA�ըG�x0�g"OT�ڵ/S dQ���@�d��$"O4%�7��&ff@�u��6yŹ�"O�
�Ǝ-U.�����,B20�v"O�cHL� fN�㕤�7B%�m�S"Op
�l��5�*��1d��O*@A��"OD�-,�|CU� �
�T���A�i#!��-9��h"�)�2S�Jເj�!�D�,D\r�OY�9�H]�0�\1 !�D��x=a��=����g�>U�!��+��)2�h@n�4	�ց��!�d�"eA�Qs�͢�x���玭_k!�$L��� X*ӴDy�D5_!�d�w�e
�M
k�����K�\!�^?(��p��^�&L��H�]�!�$יS澩
�l�2L�j��$�@�G�!򄇵"�� ��j�' ܜ�"C��),�!�d�=g.���MQb5dtځ�Ѓ�!�DW�	H��a��k+B�3��X�!����������iڸ=�!�%!
�h�EX�~Ԥ�S�I��J�!򤐩�)
�a4�����Y�!��R7��\���F�8�P�e����!��1g�����(Th�y��Ձt!�Y�N��0���dbnKuOY,+n!��t�h�`��)+b�D�0A�!�ә}Ͱ�9�"ݯlV�x�B�O44|!�d� K����Ε�f��(�4�!��;�� ��ʏo8�-��E��@!��X�[��4����p%E?O	!�DՏ*���
ń/i��%	ao��=!�d��b���ò�<>�p��@�	!�DΡC�* j!gU5A>�85M)D!���605xA#���>������+�!�D�9yl���D�Z�T<eJy!��6x���M',�`��h!�C���Y�� �[�y�
T�u!�$ٵT�1j��J���9���#�!��g
t ���\9CK�Z�!�����'e�{�Lē�IЏi�!�$
>\�B ��C+�HQ{��@�!�DN�8v�,(R�1%��A�h`�!�ć�o�B��&'�I��9U�_�/�!�d�:%�r@v�˳P���vbP*�!�d>PP��S�*Y���p���!�d�1afQ(��^�Z.ي��V@�!���H��P�ǂCFdd�QȔ|e!��x�t�*�"��c ���7F�
t!�=@�l�n_�KE*ai�GP!�D@�|Z������J���SDK�XL!���)]|0%��FT��z)㶃;�!򤘍5���i~��|)u�D�J�!�D�{�4�Q�"@�Lܡ��<_!�S���q�Z�EIx��(�&!�!�$R:[���"�i�f9^]g�Ƽ�!�D��X
a�.z��zc\6O<!�$C��>��CeXL�r��B�|6!����1�Њ��j;�1���(:%!�D	Y��h��+%��p�Н+!�� u�CA�/A6��r7�#:�p�"O���u-�<,�x� �0���@�"OnȚ�k�?<;�����6:�t!��"O*�x *�d]���H�8�HB"O�pH�m�|?�@ �*׿v{ta�"O�93'�D��rY�腈<r�Hc�"Od�" �#z<$��ř\`��2G"O���$Z�����!H�u���4"O�ԣ7��x�n�����P�*�o�<��o�I^ ���
2�F���*�e�<���� omaGd�S��S��b�<7J��L_F��T�ê%���R�F�]�<��Ҏ`�6l�� l^
����R�<���'Y����a΀C>�aY5kKM�<Y!��D�(�CT΅3]���
¤�`�<��+L�o��@��үY��e�E��t�<2�5�D-l*i��ʏ�7�ՆȓK��c��;=���퉽�Lq��m9�8����<"�a� �:�~��"��.[�l�R$�@?��-�ȓ@鲘!�C4"����}+A��B�@m�#�	#��p"R"�a�`�ȓpA�t�Vl�.|2,��f� u�����
�`�;�Y�Y.�C� �x
�(��p�h�csȝ�MԘ!��#ԏm�b!�ȓ"��8��d�50�@�6�[Ι�ȓc�6�JB�*o�sɀ x���$�،�w"ȭcNf�2��;o�^��ȓ	�t���8ri����KV }�y�ȓ3����r�]}D �f�]F4Ņȓ:�#�[
TM{���=e��!�ȓ]<۰�bX�3�n��O����T<����e��@G�0����j�hEȃ�_
e�a�!�2D0`��DJ��;��=}"q9%+�qsF�����fl	^���3"#C-s���]4DuD�æ@2	��n	&Rdʡ��!�6�� H.*��h��	R�1��d�8���E�"�.����@���ȓ ��@WN�#T ,U`��h��� \d9{��W�.�@St���� �ȓE�% F�	�$X�IJD28ՀЇȓ�����/���ePe%4p�,��.���BO�fҤ��g΍&XI��3ny�$�A�{՜�	

�9��=�ȓI)z�x� ��C�rL���R�fх�6�>d���Q�|e�	�A�{3p�ȓB$Ρ���Ì�ᑠަ��ȓc[�Txq�Z�M����`-��i�ȓ(��0�5&�Au�U�oP�pr��F����;Ţ=4�71e���ȓl?1Q���	wl��sKH2�̅�]�q�3�ͣn��D���H�S-���ȓM}ش�֦Ǜ;����W� ����ȓi��]����b�1t��_�h��
2��R���9�r<��e��A�N�ȓ;�H���P���K�0�0���Z �D�4������( ߘ(�ȓ4���6���0�^ �[&p�d`��4���'<l� "�$}�H��� D��@��'�N�ڢ��)5�Ԁ��$�&�� $ʵ8;��`��(8�vم��luC�%�%tt���H�#^��E��=���+C��k��D�!rP�8��S�? �¥��+#��#�*Ј[��0s"Ofĸ���=4��a('Ro�N�[V"O�l�hY=]�AP�I.�>�2"Ol��Ac��"B|�ۄ#�V����"Oz��FͲX����M9m����"O2�)��*~�@��!
������"O(	�a�-0��Y��˘򠱇"OdU!� _��P��v��k�"O\DX�l�9FH��qM�He�3"O��0wJ�qQސ0��UG4%�Q"O�DJ�LS:Y���3���{3n� A"Of���i�; +���vM��;N�{�"O��[WI�(*�>͢C&ޡ��P"O-Ire�	8q*�����t��"Ov\`�A�hWLٔ$�-r`(�"O^i��J�d��4&�ib�#"O� ��\1�Lʖ�5+[J�+�"O� ٗ+��t���Ё=D?��Q"O���G�F2���`k�\RVp;�"O�\�R�	+)N�2�ѡ�4�s�"O���C�`?p=���W�q�z��6"O��u�C$q؎!��ɤ[���7"O���v��z�N��K�6�x�#"O\q+�ܯ"�v�@uJ�8<ŦI�W"O��E@��F���	��dE��"O\�x$@#O� �ʴ�ͪ/�$,�A"OL��Q�
 ���E��%�
mu"O�YGX�_���#��&��AB"O�X�Ԉ��g8�"B�̬��hJ�"O��p�
;UzbTۢ@:K|����"O� �J�
8n Q���� �"Of���P9���8r-c�[u"O���s�#Y��	��lT5{��e"OKW��+r(0%�(i�� �a"O�M��M�m̚ы��>����"O옉��L֖DZahJ
U�(��"O�2ŏ��l���F^�Wz��"O�xqE��d5�ĳ�e�9[l��"OfQ���\�xe��6EDڬ�5"OP髁럯I?b\"R��*H���"O,<��-�;�iH��V��2�"Oz�u�9~���y��Y�BPqc"Oֽ�E��&k�Dwk�/oN!zc"O�]��bE,KƉ^3\��8"O� �@\#}}R`;`�?Ra8��"OVE�p���jM��ŋ1a����"O�1�!��sR!o#"�"�"O�91_"U4*�B�J�%iX5��"O�x�SNQ F��2��
g�Bx�"O�T8��\!��D)������`�$"OF-�D�@m3�I�!����Q�"O��)Y�?��֊̼5� ��w"O<bsNaV�)$ci���G�f�<Y׷}������ V�+�	�d�<�b�� E��J�+���[��F�<�Gk��nꁊq�ԇ*=���l�V�<� �C�R�n��FX�i��P	�/CL�<1$�W�4�I8d�#f�|r̘]�<��h �VDP�/���&�W�R�.]�ȓ�dx�@�;d���G�<w�����.�yr��qA�b�
3'*���Ź�y�oJ�[�,ag�Lg��Af��4��OE���R/=E�(x4��#�Ho%���ȓ^�����8�z�胊Gz�a�O ��<��� E@W�ɝm:q��*�-���"O�ꕂT��hS��K�|��#�"OX�$k� i�i_0pi@0)��D�d���'~� �S��_�N�R���?[�q�ȓ:I��`��G/����	ؑ%�n��O��(?O��p��Y�<�rO��?��y��^2sꀰ��)$��hO��ɏ�p��s��s�z	�s�3p�Zb�0���x��h)ã�)p~l 1&W�,B��>�AV$U�A=�Ց��0@��C�ɋDg����=��ak0�Uz�C�I����[B+�b��9��KG?�C�I"u����W�E5 �V Z�*�	x�C�3y6�t��h^��8�+5(P=j!�C䉭vJ8�7����^�q��̰w%(C䉍1sX  NM&^X����]��C�I�[��#b�^},�z����~C䉯_45(���7� P�@��T,�C�EWĝ�V�Z�_����M݅L��C�	-dI�W#W�W�ԕC�ܖl��C�	�(�a�����f!�b.���B��8���B5�	�N	�=ٕFȱ%M~B��T.�YãLBD��Ԭ]|B�	����%� \X�5qFhR?,%B�3W���hǲ$s�y��CF�J��C����!�g�$�$ ��C�Rx ����<���X�5�5�Rᙺ{��̋��E�<��fF�)8������o&�q�W�<a���A���OвM̈́�3o�|�<�!��p������s�|��
�A�<�RdǓE!�=�"d��M��e@�<郡��u�|���N��:�m~�<1LTIM ��O�n;�U���^X�l�O�@�4(I�R���k��
�xQ�"O����oB/xFxrƋ�#.�n��b"O� Yq"��W���鰤P�@�������=\O�0qC��$b��p��[�n| �
OF��A��n@c& ��^���f�y�/�"s pw�[�.x�҆�ݰ<���,6�+ǧV���)���T�0�!�d�DaTUH��f����t�Ӎh��IN?������$��9��Q+Cǒe��>C�	�J9�A��T[�8����x�d��'r�q��A����`��;:l�`�'� E���V�[?�8`,�V~��Q�'{�C�U?a�RxF*K,#�.��'�vHr���c��Ÿ���!*BJ��~�C
n��Ƭ�l5�j0M��O<�=�Op���0K�U`N����q.L���hO�\C��9):������D�$!�&"O�`�n��v}~)"a����R�"O����j�?.��8IZ�"���KU"O�-�d�R���N�-zZ���;!���,אpv�AaL)�ňƛ%�a��蟀RҨ�!�P�W)։ �u�0}��'�x[GF�Yb	���6������7�	���$U������^�ND�<3�B�ē�p>!u���p�X�r����y��Z�'sQ?�� D;+�P��$��NCF����,D�t�4BD�*�B$�����h��,D��fl�?4~ȕ�a��:$��ux�,0D��0�m��pL�3 �AS�qhR+D��C�(4�.){��_�B"6@�֊'D�R%��\�:9�4�!L(&��%$D��zSl�2~��l[N�!�G��>��d5�g�? VjS�7�	��B�%��"OX��d���n�8� ��1X4e�V"O���&Hԝ^z(ܘp��J[��h�"O��*�6��x���F�L�fx�����(O�|9�IrDG	<ie��I�>O�p��l =�Q� 1Qn��� ;QP��=������$D���1!�G�@���z�$�6�y�h��Od��K�,5'D���'�yrkF�	T0�5Y0��j���yrBU�^�\��3�D>#��P����yB�7wr5��.��+���Η0�y���Q��m���o�~�Q����y���H��t
Q^ItX��A��y� ޭYE��@��EQK��Ж���y��eXī��<G���6�[��y�+�5$����nŕl��	H�M��y�H��P\�QH2��Op��ȳo���yBd0�R%��%�@6�]��+��yrO�H�z��"G]����1�yB^7�����D�*�k���y���*쒽��݇�%;$*���y�'�l-\�#��"L��y�IH�N��࢈0���:B�Ҕ�y2*�?u��-R�/Ԯ,AR��V�y�&�cb���B�jt�4�э͞�y��@�<uŅ�s�d�B�HF��y"/.Hm�Q"rKq~.pˀeV��ybћ<��qc�
f{�{�,<�y"#�7mXL!���d:��p���y2GT�N�*�0@�R$	�`��G'�yB��&ZF�A �w��T�FM��y"Ej�r��F���i$c�ϵ�Py�NK�����V4fc5rbD�NX��Fy��׌�2@u&��e7b�� ���y`��-�n��f��mFr�����5�yҌ&4��D��̜m�������y"��++*�{� 3$���jD��O�=�O��(��`�.HxR*Y�v���'l����9�!�Y)f�f�$D������u0(�xA��*b3f��w(���0-�t��x����.�������O.�=E�T)��<�Xzȗ�$Ǵ� E�$��>aJ����Ê�2&�U�� �0ON4�d�/D��JGo���MHP��'PXT�Aց8ʓ�hO�ӭ \�-1ai
�W@�9���frC�I�~�B��)x��y��̏c�Nc�,F{������x�xq��g�7j��4S�� �yBń�B�
h���^�L\!���y�m�y�tA��TO]���ø�ybɐ�Q��CulŭH�,}��,��y� ��r����aE�9�J�\�y�צ��[GAUf�*�Q�E��ybČUTʜ�%��]άKU	��y�̈́�a���2��O�l%R�lɯ�y��Z$m��X����P��+A���yB���RT�)���r�,�rw)���yR) ���Af�z���&l��yb����%��ʍvh �
�P��y�J��H@�$aQXx��RkQ�yB�A�?�`�6��FpJ��ϵ�y�OL�|��J&-�$�d�$-]��y��ނj|ʝ3�Ȕ��20ɗHF0�y�
{�ک;0�OY9�9��#޴�y� )J�~b�JF�M�2��%I���y
� ���� ��m�ƥ�sXb�h"O�����_9Mր��R��� %"OK'�:�h��aP��-��"O-c`��w�0��;��Y��"O�$A��^�B����[�x��]��"O��c�iF fj�<#��w:�� "O�k��aM(}B�4v�AW"O�`�c&V�R��3#��K��D��"OT��l��}�´�`)�7H�"O, H�oț���EF�x�T"O��#����j�t1{4be�vi� "O� ���V���ن
�V�H��"Ojʕ���Z��dK�f���+�"O�{GB��z�h���F����9"O�r��̂qP8i����5ۘ�J"O@91�DfEh��r�*z�>�@�"O̀D���L1L�c��1YU"O����mժ��8�w�s�h�k�"O\����\�p8	�)S�:xC�"O�TX 6Y�>���H! a���"O"�J�F�	i�h02(W�Y24�d�'G*$ad˛+�]��)�0�a"�E.�$�ٴ�C%C� ��'6��u�.I���0��&e��P9�'�2���F �L��d#�H.��[�'���Q�_5�V��&ᛇAt�J�'h�����/ɴx��`�
�'c>�Paǿx�H1H��G+�)�'\z(�@%��.$���b��y����'�2��f䏁7�i�e�Ӷo���	�'�L���Ӎ�vmz� \�e�Ľ��'{���#�2��U�4,܆P�����'�t,���D�G�b!1�K
?e��|*�'2.��b��'A���CG��2X�@�r�'�P����";�ށ��j�]_�=��'�Ta��L֌d�`q���U�XeC�'5N��~��� /QG�괘�'�ePW��x�Zw'�B�Pś�'c$ԙGJ 	4J���ѭJ]��H�'�L�@ř}!�p�V�,t��:�'8��2�f�fU���e�3^���'0!)6"?�D	Jb��p�ƥ�
�'Ś��7�\!p��}�f`1�
�'�8�����|�0�Ⱥ:B����'�)��	S�*��)��m[�3���'�г��Y�bPz�3�&�8�0���gO�I�a���g�z���>��c! 	�wJ!�D��0 `�#6A;,�8�镈Z��3Ҹ�!����S�Odȭ� !�t�p�$R�1����
�'~��AC�&+0`%8W��<1�p���R0�2zd�%��~�?c�|� ���lɯ�zU� �{��HA))$����Lڸ	=fݨEkeֆ�'MYLϬ�����aǁE�,bB�(��B�d�F{b*ýEe�U(A�S$��N?9���̋�"4���D�1�ȸU?D���&c�+vr�O�'F<��a�`@k��ŬF�,$�d
��C��Mӂ�M{�|[�'L�8�0L���C�<1�\dM���iI���������7�ɖ#�01a ��5]�����hO�L�2�XL6$���aubDؒ"�'i��#S"V�ei<`���`$���fԨ2�<A��Q3����`�BH���x6��!a�\P�������/�	2#�L�iaL�9F�&5в��R�O�t�t,�[�iZ�B�6R��
�':6�:���r�RH���ܐ"���x��S�gDXr'�D�O��)n�h���V�$��] ��_/|�fIPTE)��|2a�	� X�uk	7n��(�MʥJ:�y�����X� تx�d��4~�^��mO)l��>y�	J2>p�!� Q�{�x$ar/�j�'N��s���fx� �A�n�� rD��R�,}1� ��K���~�qKxA>����;P,		��>��`�k�����*/V@�%�SH��M�ʁ+�!���Pu�� ;��\�T�]:��Rom>-λ�Г$A3Zְ�� �{����9&\Q��D<��1��	/�H<�����^� ��V��b)�cu��!�:�R�'��,#�H�'���;� �8���BY 㤨#ד ��{����-�Q�#ω\=�L�G���p� �)n�x��e�&zo�d��V�U�L��&jכX4Q���0�O��p2Y
Pd0q*9�I( 7��X%l�v��h��D�D�B�cHW��Q� GW�K��"��˒-�>���ؙH�l��T�K �p?�4iϨ4�aH�V�TR��-L��R��^2lJ���H�SSF��ĉ+?�M��)T�PZ����2C�`�b#b�(m�bSK�E(<�AY�
$�RBʁg��4���n. �+P <)#�X�JȂ[�-��?(����`���U��i!�䓟|�^x"�(4��!�'�@џs�锸�dȠC�]kM)���Q"�a���.?Y�@�m��|�{��صi�؊c�ͦNچt�@=V-��Hc����_�f�:E�
�j�{!B�>A#�*\L�6#��纍���,S<Z��R�D�i8xn9o�%�)� O��ҖF�h��K�m���� =#�s#�9I�&����K~%��bA�0���M:��D�փ;(�Cc�9H�.��� H�.�I��pۣʖ�^Q��R�Ŏ�
��~��B�:(��.�yM(��fl�M���@i�"�ة��D*l�4d�dJ��S���Y.�}D>����C�J���'`ze!�Ȉ1ي%i2���h$��� ��� �ِ#���1,�)odYY"
ҧM�2{��C��<³a�>
�>A�t̒2� ���/!>�yb��c����䖣O��C�֣�y2�ZoG`�tM�5.z��*�2d�����W H��8k�b� x�V	��a�PIz�ڌB^ݠG��Z���D�	`����WC��p�6�2�A`�N�� �$[���b���r��Q�ˉUF��R�n �0��n�0^���u�}5�E�׫;ca~Bk�����*̊���D~�r�B�BF(@H,�i��X!�DH��k֮A%z�zt$S!��!��Ňz�h�:t�|2�X1%���)L �@�i�f�0�O����1*�q� �
2��xc��2eE�vѨGn��`oҜ8�ē��g��4����4ѹ��.<O���eD(�~��gˍ*Y@�q�=OD��G�Mq���B��B� �����bC��:Tph��J� i�M�2���+��9#ċ^�F�(���oQ�񤛜_6X�I�l�Ec�8RZ�aʬ���DR�ʘ	��K"&D�)�LZY=J�y�MGf��d[�g���a�ܝ��_��B(z��A#>�a~���K�,�ũ��>���3%�-{'�l� ��3s���ۣJ<S���b%
�dKg�L?;���k���|(�'�%Z`�Z7?�]�VgQ�y��]bH���0�N�#��	#E&M�F���B��6L�2D�I�}>�"T�ђe�x��o�"I�������u�@��<��<I .ҍmh��N43%*�{���V=k�dsӢ�?P���0��kr�k074->��(��*� �9}�	��9�Hݳ�ʧҰ?�d� qi��cq'G�$�D��I)y\%�"�8|j0B."@�����/h��sQ���u7h�'��]iD$˛>�R�KT��D�Z��}�U�%�:�.�8GH�lL���i���{$�!��X�Ƭ�D$,�ŧ&k���9r�'l���K���!Zu�D���Ο'��d�6L_:IqO 4+�kۍn;P�XNW_E�\�v�Ojx��jĠt���j�%�5B���[m2F� ����XJ�p��h�����I�* �$�΄�m%3 2-�@
g�zRiL�r�pY��ɖ;�F��Y�%?D|7E�7?q�L�3	T-Q���p£�$rT`�s'�>�T�BuY'=Dxj�E��;x�h�]�zY�+$ �`�f�mP���DՆoV�5�'E�4S�|� ��ڱ'�(hK6n�
��T��׉VQ�[�+B7d�>��)��U�j�8�%�0&�*dcFn����0n��2��-z�<BA&QW[��=l@+��S�k�:�^�q4@ ���¡�1L�ᚱ�ĥ.�8��KD%:�PS�_,rX@�,S�/�@\A�CM�'1�}Zd*I*P�1��."���q��D���JU�P�7���z�k�c6�mBDJI+S�-)�ܯ!���QVc�Di�����O�^�Hs �)A����'~�pѹ�Ը�o��2��PTg	"X���ɍ�?��-`�K�Cx��h"%���ؤ٣�^5��)�wy���bg��v�ą��%�>-g�	�,c�X!,.�d��ƝJ"J�G$5ꡲ�,G�|�1�Ҡ&�Yb#+Y�z�`q���O@�S��9p��(  $ׁ25޵���$�����$94�� �sj2UYw��|�v���)��V)Obm�GN�o�!
�p>��	N�K^��ghءP8����̘͟��z��!ru�+�J��N��H�b, �	R94]'�P3t7�m�D)D�����'39�\�s�Z4[�ޙ�2��=e
Y
�cJ4<`�iӵO�*)�@ʧ+��O�����IL��V썓ؠe���'٦q�A˼jK``ѳmџGjPDɠ+�x����oǔ8��&���6M��-�,�E!��ꐥ���S�}פlF{�)%�Pu �@ĸa����$K4*��L� /�R���ti�8&��C���,f�!򄍃/ jMY!��)r*��ʖ&Y<U�0�"��4T�ׂ�,id����L�,&fYy�5�jޥ��ʒ�V(��b5���;���9�*+D��gC�3GN����=�teK ��|9�k�� [2������7 [���,�eE(�|��O�Rdjƶ[��q��]G��JE�'^F�K7�@>�^��g�h�? RȊ�5s�-�7�ӓ&Pz�H���.}��m[g��0|�(Qb%�	�p<��GX�=�<�b�h'n�*V�l�o�"!&j�-Hz�Y�M��u� E�F�d����tG��N\A�uh�%}�L=����u��e���0�4i�ˇv��iu@̆P�V�qg@PR�n���'��U�p@�鄛r%k����IU0�T�Q�p��5i�ST����-�9Z`ԁ#f,4��0�g�w���R�o���m��^�3Ϻc�L��Ӑ|��5�^9<�C���w4釭0?��.^.=�m��B!
 �����n��"�P�,�}jw�W�2~$ۢ�]�0��C��J��|bsA�1*U���U�N�=2�D���g�'[x@��k�$�=/,kg�ВY0�O([�_?�P��͒-R�PJ@B�2p���4+7�]�s��
��  �_9^�8Ad̢9�4� �O�mcԌF�%��h34�^ f�������A�v81r)M7@&�%0fo	>�QoZ&G��������yW���B.�98�]y�ܢuL��xr(>4n�akV-X�v�����#��g��ɜv?�����'�z���ˁ"���y�O`�`�*�@F�$*��_�?}��e�'G�0D��:p��j�$�<=��7�8tAq�S4��8�tÓ��9#o���$�(�(�!J14%ȉ�D�6Im����+G�>� 4�&=7�'�8�D�N�8:�P�d�;��J��EL�\��3O�����.�$��L��!B_�Y��J��'��2f�W
�̓�m	7Dc��p*٢e�6�!5�=Zۚl��ȈC��=J�Q�諕�	�Ec��@�w�@8�0�#*� �8��ɑFY
���'�����0?��CaԼGǜ|xUk��yp1۴zl,������zQ+@�έAl`��7fC�}��!�`ʗ��!�D��1B+��P�,K�.�H�w�/\O4���B	)]�)�C�R�TĘ����V�r��A�O<O"Bd��L��-��u�V����B4\��"JQM�'SZ���Y#�4�聪�L��k�{r΁�O��"	�[Ši�id�@W�҄$�D牃�����!�!_N@p���$o�b@�j�iL:��'o����ᄖ6�1�0�%*�J(��]/xPT���^bM�bME�+`���'�H���Ӕm#aͻV[�``e-�e��ԛ�L�/
$.�`�O����^LT:I?���"���j=��A���M�fAЎ+�bH��V��M�3,�00�ᅜ�N,���)���M�#^��8CC*Z.V*b��b;�
S�1�8�����	Sj6<ؑ�ŨKF�,��꘺u�d�D�O�c+�m�w�?9��+��N��H@F"{h~U�CC�t�H���g!�]��'6��c�,�q���>p���򯞳>)qOJu�7/Y�6d��G�H"J��S,Ux���1a.c�r�@���,a>��ƕ��	� ��R&��b�c��fRey�Ȟ�b�v��\�rp+b��ܴg�́Q���({^�q��@�a�[�)\�P�$�ڧ��#� ����2`�ҽ)E�i��03��gʠ!�w7ֽ�sKN���x`F
U��C�ݺ?��8�K��"iօ��
8�����]{ʔ �$ �2QCb��%�?_����w,HL oڬ]�l,��KT���/�,p�^�z���w���7,<n�v�ywh&"/l��`��$uT�&i�u��#?i!�]�'+^�s��<��$V�6�L�1���5#r���N)]Lv�#�.��gt5)���=�Ƹ��vݍ#��ĚXDĨ�!&ϸ2�b��B%_��P���A�T�.�ش����'��bC�M�(���� q�&arA��"7�d�4kT�*����Gi��I���q�b�79$\��bL̬~���d	��!&�d��,���7������ 0�i*Ui�1�U���=�� P���:e�Y�X��!0:H�کRd���ѡ�)��@bޙ��&X�$6�,��-MMn�dY��śhl�-["�-��h���"RH�3ړD|�0�E�_c�]�D��I�� ��0^?���5�ٔMO����N�F�8�%cϜZn�a�D$كM��04�N�S�b� d�6y�۠��r͜x@��Da�p�����ࢸ$b����k�+�*-AcDW�s��t��L�y�v��2��1Mb)bWo�%K�8�W���(�"=a#�סs��@�t�z�x��J�i�N���mI�c�fM`C˅��'n�x�@i��fޤ��So��H�R��P�O�RmH�M�Wp��CI[;��X�e�5Q
q�q%G�;����,�6fP� aS吇Q|��s	;��O�
�ÁN(2Y:WꋲxC �j %)C�$0�4BR'v��ӗ�V��)C�> ��ⓤq��$���~�.]�@����p"���b� p!��*��<�	̥gK4q�m�UF{�,Z�`�0
5h�;Jjp)��Y�ʮm�Q�#P����d��C����'c�(2�HϹNzXAqd)İQ��^1۰9��#�?��٣�E��Q�͛�o?џP�W�OFx�7�͆,(�����Ñ���4p��b�\��I(a

0Ȝ�.�uw��yD��b��M�OLE2���b0,�YC�R]5�H���H�v@]�@��a6 �q��\7� Xg�Ԥsoj�
�BS�q�h�M<N�|K�i�\x�W�!Z����)���y��)P�[��`��Dʩh�F��/5�X6-^�M�XU��	c����0O?7�x��2��++`�{��L�:�f��'�XU�@k�
ga�!͟�X�F�5&���ۗ�ü;���0���E}��^�e��!TL�L5,"<)���lc �Y� �.D8�2�Lڡ��ekP�ؚ4
2���	/X?�;�*�`l��B%nJ� ��B�	�l��R�$�*y����1��IBdB�ɗ%��kv�P6�zIB�+�}rB�I��|�93�U"*"~���62�NB�ɀE�i����F<��M[�.
B�ɹz�|�1#n�R��v�W+�$C�	�,��yC�+
��Y���Ֆ8�B�I �\ԘӤ�3>�e�P�O���B�)� `��2��1q�'�%dR��"OЭ�ԉP�aPRL�:'S���"O��k�	̃ dt�i"N� ��"O D� >����� E#�Ȼ"O����+��,���(�_.�@J%"OL��`o��5�B (%]�;
Ys"O��'��s�*�qD��:q�8�"O,=�G��U^�@��\�>y�)�"O���OB=G�4L����TW�ESb"O� #� �2Nތ�A�J�i+x�;�"O� ��I-�h�E�^
�sW"O�	3%�>d}�XC�d�o�(�"O�Xڷ�JE��c��B|}{�"O,��raW U�uIC�NR����"O�ia�l��C):�����)c�Z�"O�����E� ��9%a����0��"O�QoԻt�ȨRaJC>3�B�bG"Orp�4jK��$���ǢD�^�8w"OJ۳��(s2�� �̴S�Xe 3"O�p�EV|��]���k�䴈@"O�����Xu�p���ٺG�%9�"OZd�����-P/I�m�L$S"O�z�%��h��g�V.j\X�g"OXͨ�	�c(2��ժP���\ۃ"OT�pp�� ;t�0�՞{��:""Ol��Ɵ�{A>m��� ANH�q�"O��a�'k�����4'?����"OԤk1`��Px>CQ"�Z(Z��f"O��CV�2h��7�K�>  �X"O�QB"	#`��XP!�O?|���"O��`��_����"��/(�T��"O��j4��4m� ��
2sRx�"O�1"�Oܳ4���'��\	h)�"O�}��DA@�
�Q��Fe*�"OR��'C#j����X�7��+�"OU:����y����U�	���V"O*X�ָ4��1�T����$�6"O,������`�+ �P�L�h��"O���Fĭ,bd�Nʵ��8�C"O��ɐ��
z��0���<�p#u"O^-c���!��4����>(�8}�!�D
�a^~M�� 4 Ҷ)KX�!�>�$T�dD�-�"��"G��!��Z�c ���Ϗ�iC<��X�f�!���Yx��	�*��㐈�U�!�$̇G��u��#6�i�(���!��-I�r	b����d:�=�"'ɩq�!�dK�.��[Ѧ�?�y�G��%n�!���I�R����2D��G���џ�Cq'y��>yJPcC�A~f(�5oP�,�n( 3k6D��� .J�HS�L���	E�l�S�>�"Ҏb�F$�G�x��)�6Fl�1aDysڱU�H�d�!�ȔzS
xQ0�قp
���ݒ&G��,� ��:'I����'����kZ\���T�0{
�+F�%�t�V�v^iH�{��YN;=(^�`'�%Ra����8�)xj�)&��)�F����hO��̎x��JI6~��gب�A���s��U"�B��L�����Lp2'��$5�9jq�E5=���o��O�x30ć�B&ڐ��G�5�ȟ�)#Ԩ��i@0�vt�a)̥�y��+a�$3%��7	���D'
�"���n�e�L*qF@7��hi"ԟў�
��J��H9B"_�$PEC)�O�� ���AH1y��� ��P(bm��uJQ�bH؏g�v�@���p?q0� Ӝ�������k��Lp�bΚ�1f@��0+�{�#ԯ�Q��x�@a��v��	b�`�(H�\t��"O� ���a�=/��,U	,�޼�'l�r�n��k�H��R*�
}��>�ɕH��-2���h�X�"���26�����S���kVeүe�p%(����OC*���R�Tz�ɫP�W�#�fu��$C	M-4�1u��>	�t-D}��؀��=�_��9�����O4��Ͱ6I[���&,0AK�C��>� c`�ļyRP�g�M�liDB�mT��W%��p?q��29����f�O��͸Fh��h�9��n�k���d�Y�h�v�+&߱>����aFڹL������0m�H=���oS6 l�!A��q�<QG	5�,�7e��O��SQ��}��(C�ˠx[�ب�@�6��;$7ܤ���"90-c ����~���p@Z 
�mX-x���T���p=f�^(g(�+$�S(����!�#JD%C�߂{BR�wB��f�$�+b�D�#����q�\���,"�e	���1�эoM�-X��
r
��=y���8� ,��xP3 B�N�+@��1��qu��4V ���_�v��DK�ON�R�`)hC�'����lͿ���y ��:BBE��a\�n��ȃ���l���7?���f=���Ap��պUmn�Y�0NS�A=�S����L���,D���Lֹ������Pl �a@.�r�k�M�?"�ԑ2E&� �м�R�8��{Rk\+Wc���O0t� ��+D��!��N�>�B�K��'�"�+Ǝ7W��� ç�B\� b�1 ��D�N�(%<�� ��	+@,{)��;�d�j�C�	ґ�(��"��j��)5璷&9<�3:�ɓ��=9��P�~�h[ �*>���1i_�P��Kq��:0�
�RC an� �R\Ɇ�#s� �O ɑ�K�.}t�@tNR�]j ��P�Оl�:Ԫw�V�C�:��U�ѹ��kC/~|�XTޟ�E��w��e2燐rt��Fk
 e����'��ddI;��/:�,��l	�|N-RB��A1�ݚGC�ÈLC0G��'*��Qdcެx5��'�~� 1���%	��05�5!��Vn��L��LaF��e+�IA ���[���&tO�U�
8* [8,PmpO�&3�������*1�R'ʇ߸�Ӂ�0�qOT�� �
R�t,X�i�=^ �6��똵0�� p7���t�D��]�6�0���QO��e�@�}OP����
�f��W��[ ���[�>�� �G�y�,��灲~KT�O�,杆J��m����/�X}����kD>B��b�Xvn�	t�E���ѬB�t���a��*�>V �Rt*a�ՓQ�85-ʡ*�|r�H�2�����6L~�HDAR��<���6N{� �ᓇI8v��TJ%<=�	a��(BBzl£�/qJ�h�#�ٓ0`�z�DG'>��y 	�WOr�� CN�9��vj]��ēp
�)�;3��"
�vz���'�P�c�,�+�")�҂ՠ<�\i��G�4z��i)�l24����&�-�r̘@g����!�v�+~f����{DR�I�h�|��'F߯�z�̧��5�(v��T�GR���o,��d� C7��G"$؉�5[ AҤ�[u�����q�"]ZD�@�-=R(�D��ޜ!#ȡɅd��Gݺ�'�d��A���q��!Xy�XK`�<}��T�B��4��O*��q�ʏ�l0�E'�6��Ycem x�D�@�_�(0hЪŎ]��xrg��DX����\��I�P���p��8/E( Ҁ�B�.݀8�'��m��x<P��D��RU�8P ��$I���hK�r��Q�$\�J����:�3U��:"K��$	�L�x�f�]�zX��'d��t�d�BjJ�i_�9�pg	|I䥠�L)��|�v��{\�)��s�H���oP�!���ɭ���2��K�ޜʲM"�Ofu�.VN[�X��'��Q$�"//d"�'H�$ؖi�4"5 f8�bb�v�\0R�X$L* u��@��( z9Z0�	��'��v�	�Rv�{!<���Q�'M�|��K��}����N�M�6.�	Yl��R;���	@g�jI�����.�D)���*�Z�	��9k�@�bM8:���@�I�f�@��
\`eN�<a4��T	�V�X	P@�R��#6c�<M�t�" � 
^Ta�nʾe?���"�.����&�XI�#L��}2,�Xhxb.�=	O�`�D!�����u�����H5VNR�0@Ϡ9��A���>D�|#��� ����p���'|r�����%h��7���Y�ў�韂p���i��^���e�1����A74$&5sE��0-cB��h2x4T�B�S\6�b�� ��(�ga#���/��`]���SK���<�I�[���P��=�.����1��%�	cZ���#����,�0P>�eL��1���t��u��$Y��7D�xd�$�b`�P��9���.m��%j�NS�R0�t֏jixQY�	�!1� 5��a�b���F��f��.�+�*e�N K�Fa�D��"m�}b	�dX�Jۤtޒ��瀁�K�" Ce^7J��awجz
ԋdk2ES�e��'rӈ��Wትpۼ5�0	ʃ� }��h�,`�2�=�$��k�2p����O�4��X�N���
q\�T�DS*[8	��B+� ���*C0����'����)�39��Yjt�+	�8�/�.%۳
]&A(ƌ��/Z	6������. ���ϞS�ЈĆF�\���2 	 �E�[{,HR���ze���Ѓ�5T܈�'¦�4�Ç��J�4c6�ɁO����!�W�ӥ���%4�D-�4�
9�dD����W'�n�T�
Q zLP�.�qt�z��͉D�
mce�.1b�ܒ��O��hO�a[�<F�J=I�M*����3k�76$u�w� c���0m��"�:D�� H�Ѧ�ͶJ��3CD�uw,��ǫ�l��`�D�ڹ0C���'=y�Z���)��H��z�%i�
����4Ϟi@/�W��C�	5F� YP2�V��p��AɺR�|m��$�ni����r��c�lv�ݛT��9X�f���<�dR�X��0t� T���k�b@���z"hU1>�ִ(0���K1j%x�GH��@���L�g(v��a.�2$Gn ��M�\��p0�����dL96&��+شK.���O�1O*��b��
L�Ȉ[�ΰ��i��8)+����;2!�12K�.PG�4���J�,��U�Н�PxBc���A"w+E�#��$�E5K<�ȉ�Z&v�^򌍰F�Lx�Í�
��e���|4.Ŵ�y�KG�b�4�!"�ӊ&�$�3DC�3��xB��x"V\{�aB^� ���&k�$�W�Ŵ*�,�����P�
f���"70��яn�IV������2j�	[fHʷ2����D��1m�%;��44�� � �� ua�9ZtO�HsV� $�C���X B����ćT<I"p ԎHA�'���q��9s��pբZ�\hX��N>a�b�!XcB��/��"V@����Q �1�uft���CC�F�<]v��B��9-y�l���Zw�~8��E7�O~F�رea( �7#�����Ff�!S�чQ\cR��^�`,m2e�ºs�'�-�yw��Vd"ͨ2�.%D3C+_���x�_Q�<� �E^ F���#E2 ��pL�Y�ɑfH
�[P�Y�-��sRr�y�Or�����^r�h� 蜫94�����'s�|�])<9���C�.>�v�"s�D�/�V@���-�PR�l/1�^���ķx����a���~���$K�z�
5CAW�q���⑷(G�'p��1���5-J�����2�x=p�M�g$ E�4O��:)�$�!'��5wX\Jd��NFz���' ̅���%#N�B�݆OP<)�q��
fvmj��U+G��q��R�ҹ`��%X�zdK�NP:9��w�|��aM�D(��;����I{	�';e��E<��DXFW1X���C��XV�p�۴	���"f@�6_�p4��+˞)u$�� J�f�p��o�㦕A̘����.�C�!\O8�;2%�;m�N�)�"E�3���x��o��\�`,�]F�׭N`�L�f���<���E�u���0�T^�'�"Ap�dQ�BKEy��I $̞q��{Ҥ��e�.����C�!��	j�Ȋ;Bl��<Q�b_�0�$=2pDŀY�5Ѣ�ٷc'�P�H�DV���?�hK���[��.tFÆ�O,:����)�  P9���-8���.Js�pQ�7�yGdSi/z�0���)D[���g�WE�I�S��8IKNs��g�u��"F,�G�YR��:�r	g��"f�jp`4�iIb(���$�>�!4��Φ6��~�i�c��Of �hb �8�ژqW+�n�@!�G�ŋ$��#���-6q�Q[5��"�,�H�<LȀțg ���p5�Y��>�T,�?~	�a9��J�Pl�i���KŖ��� ���,��(ԋDlA|/npCd�T�Xe��6��'�
�0bZ�g����ڣ�t((p(�+�]YF�i�dP�٫z���1q�\�3z`�r��sՊ���Y��ƙÇ�+�MsP.�0S�n-SK~n%|��r�^<�<�;2oO5@Pa��F)��јs�>'�d|���ŗ"bā�4w�E��D)�j�̻k*�%�c��d��d�2J\�92b��Ƣ�28��xƊ$+��!г�hF{��y���:��N;N�T���^��%�Gݯp.�6-AH��\� �7����.Dq�<�i
��u7��>(����W&@xu���� �����Щo�ti
���S�n)���[�HV�f�y�ٓ9��:f���hU;O�`���o#d���A��5�uW�Y#eL��c��ٮ(Cd��X�Xft-C.�:��*� �j�n�`5m��B%M-Ck��z���Sj�<8�m	���w�6ͤ02It0p2���v�u8�Z�'������#d�x�A�0ƶ r	+��'p*���FJ V\��GC�SN�()Ag9	d�xy�e�/x*A�J4�� ��%]J䲷BPK�,9�w��=� ğd����L5Y2m"��]�B�)p�Kw�҈(cŒ������I0}S�}��ڏ<��x`�M$0[�0��5~e���s�e7�XRe��}Q�e����;��L8���%3[�8��4�. Ђ�Ä|F 7di^F-(c��.�8"?Qp*�8%�p�Zcj��B�G/N��I�`�!��KG/0%dԪ �!�-C�뉂C�v�r�bG.L��i�`��'�� (t���3#l��Bf�3}��d�p���'�< �'����t;�*Ή6q\�p� ���ޜ�D��Qک�Q�с]����P�͉O8.UA��)8 1����
�҄��S����?	 gY�M���E���3E&D���w���aZ�ZO^tb�æ8(B�1P��9J�����1F L�SݼCe���[S8H��O_+bx�����P1���%��H���z6�;�Q�g�'Ui����~6��u�A&-��'E7�JLY�R�Y�X8bϼ���mD�v$ͱ��� "��ǥѴ�|���3�R�#bJ�4�ttB�V�{LrQ(�	(�Xꡍ�(X��A���K�Q!���w.�b���K��ӵ	��:U"��hJ�U�:M�Xw�@��w9E���t��E��h�
�Xc�#�8�0R+��(Ov+ԅ�k��h	��!�>� rk��AZ������^|LI���Hv��6�J?�����+/����I�}�Y�����z-�扦LLhA �Ǯ�jMɖKe��0��		�"�����-(���s�ؤC��\%#�J���c
 *Yzu��z}r��� @ I�*���I+h}R��)��='�	`p��/3�*��'�&�)a���z��G�52�ˍ�?+F�@��G�Z�`C�)�&���)�	E������T�-s@� �LaCg�;w!�D�}�R��A�ęt��D�F��]4!�DV%rP-�檌�M��J"/^l?!����%�DӰ���oR-.!�� ~ z��C.M��K!
�6B�]�"O�x2�̊�rƌ�� �[1cJ��"ON����G%���PЍ1�\̱�"OȈ3R���&@�ł:�N��"O��C��ϳK� ��e��7-�`as�"O�=jЎ	4`��9���'�l�[C"O�A�3��4�:�S 
1f��PA�"O\ �g��n��$I�C�3�(|��"O<�p҂ޱ!�<�����4����"O���@�m��}w�E�F�&H��"O��[7��>���BR��@1s"OftB���Y�Z\�s�%A�|��"O��sp�U�}�
��&#C9#N� "O����k��h�Q���=C���"O�����(�1�/od���3D�Da��B�X�����:Ae�h:�.D�d� ��F;b�C�o� Y螸Y�,D��Yv.�x���"�CI�`���@,D�H�n��"c�9��5��F*D���`�PL�����_%� u���<D���nϣU���+�DW�S� q�#.D�T��mڙd���8E앢B�h���*D�(У&��/,X9��cօd��@��&D�<9G���2��Y��ˁd�ʄ��$D��S!�\�X�$�1����̀��%D�|�� C_�������`��1J!D�h��M���B��̷� D�o0D�ЃV�'?n��Cm�U����%D�LQ�D:CL�CSE9��YSg�!LOҝ�ҁD�K!�K) ��xx��J�Z�Pa�[Cp(�'4��S��$%V�d�	�ύ� �P��&)�+ASb�O̥��mx�O�Z����C�,qE��ŉ�n����5}B�˓/�dy��5�Y?�'��y���}L&�E���=z�E�'���k"a/�)�'*�0�Y��>(�����]���lZ2
��O>		�'&�F,���w�V˵%ܠfe��h�M�ryBw�1#��'�x�	�*Dd���D8C�t���\�x���Ӻ:tk�ꦕ��:�N��8~��p�^'F��� >e�B�a��xr�0.k��S��R>�y���fK
������EZ�~����'S��gǟ��D^z�O��C�k(1vё!eU�N3�S����T�S�Ȱ�������>
0�M1_�D�A��e�JxpQ�  ���<yA�O,��h��E9vbUؠ� �.!����	v����M�.mZ��H�������<�M�y�
p����~ʓi�Y#�'�.��	�',9������=^��d�`"�`H"��	>?ٺ���M�(O��7�S�&����q͝>?�Α���>&��cROJ*�?���<���!�Ƞ�f��#3�r�(Ӧ�@="�������	w�S����N��0�	�^�����iU3!9�L<���"���G�V�1CT��L$P��5�V�����O�`*��'���՟�;��� �,|~��2$��ELn{6j��~��ԡ�7�&�T?)jJ~�s L����`���<��� ME�=�`2�(�vݛ�'�<��|�>��4gܐ5@�y�/�,4D R%_�Lr�	Q۴>��	���x����3j�8��%�'a�-�2��a�,�:�O��P�ըN��"��I�#�ziI�'�Dq�f�9LM�1�kKz�O��1@�6nҴ���'�����BH�cۆm�6m�Y���rƴ�?�'m��U*Zp�d��1
?�b�'�΄���
se��O�
.�p$�
�'��샵y��$D�w�BXH�L:�y�%ê6	(L3ce���`C7�G��y2�ΟV���ueA�)��)�	8�y"��Q�v�@�	*MK�A�G'6�y�̓)g0�8���ޤ/�]�6H���y�V B�Ό�S�	$lȩ0�K9�y�a�w���
��L�dM�Ա��@��ybB��&p;�"��'Q���Ι �y�)��w_d5
���,�����!C��y
� ���+�~N��B]�,�ȗ"O���v`W0 Z�āV�,H3�"O �
W#�<nDD�#�K�8팥s�"O=b���M�4u�T��|����"O*�`��P:sl�Y�'I�"T.\�w"Op=��j�2K�I����#.�:�v"O�,��F:P�uf�	C�t�J�"O�i�
�EQ�`��#���q"O�5q�١d�I�3� l�By�"Ov�Y` Z����é)/���{b"O���2�т2�Vpj��\�x��6"O�)���O�~�q�)	!s���"O�1���TrY:��Ǚp* s�"Ov��Q*�d@���n`���B"O����/FFS���R�!H�i)�"O��tǌg��rF�%eX)G"O<Z�+�_.2�����aF8�H2"O̱�f���pjR�y6�7TRHx1C"OTӬC���r.�G�\i1�"Oą���C����/X�$o��"O� R%�����.�:x<����'; ���M�HER�`��I���R�'���4eQ%hyj��I�B�x��
�'p�I�r����I��J�A�h��'�J8�H�}\���3藘;kx	�'�h�$�1#�i��<���^�@��T�8[
9�`,��A�Ꙇ��6��эN*H�����C�ˍ0�'\����+^70�����L��'L����X+w�!s�/Ǿ	a��'�8D�E�V/��}1To�;Q�(q�'�h�{F���@�Z��B*'`L�
�'x��).U�>-��a�%|�M��'��H�J�7�X-+A����q@�'�h�@'�21�֡;���*$��(�'�T4�}ï�'��zy��1�'$r�qR�k�؝۶��|�E�\�<�oD6|�yذ�D�X��<�� �T�<I���&^�����C+|	Nݚ#`�L�<1��S� ^�=�f��>��"6/YK�<��?]�&�s΋�;B(�  \�<�s�]9'6����Z.J�4�
a�<AS�!佚D��>�"U�6ȕZ�<�&��9y\l�ET"!c�kV�<��Lߢ#�t<+��(h��U�O�<�eء����ǟ�	 Sd�L�<Yҁ��ZH�=>
�
;1rv܆���A��`R�IWNp�b��72^��ȓL1�jB⋻8k�0 կ�,^�D��|�p�ڡ���g� ��� � A2i��bD�s�!�/#$ӣ���60P��n*1"௘�T�S� ��U�ȓ<h�F����8Qj$<_^��ȓn�qQ�a��:��#��O6P1:��8�����S�t��6�X-�ȓ�a#���?>\�!��j��|s�Յ�K�Y96��ur�]9$�_�4����+S�c�͑*�� �v#�5SR���ȓT|$=�-D����C'S�= H�ȓ2�6����|
� �A��]3����F�Zܻ��S����� f���ȓoj@i	��ղt-Xtj1KD>)j����I�d�c��/X}�u�F	Z8P�0,�ȓ)��R��7r�����M�=/h&���S�? ��Z4� �9�8dh�� �>G����"Ov� aۮtK�X�S���2�Pu��"O`	e(��C�$PǦA��bY!P"O��;l��$�B{�Q�"Op��҆S1����V�d��,�"Od��M�5�� �ʊ��L��"O�����+2h�Q�I���D�{�"O��j'�@�_gve�P��\㨵��"O��XrH�,Q�t9AF� ���"O"��!ܕx6Y:E��[@���"O�d�e��]l�p����2X��c"O"�2q��>@�r���#C�P�@�R"O��#���|�V�����H�p�"O�,�G�<(k^���!дF� 1��"Ot9�%m��2V�R�/�6Y��˴"O�0�u �-{r6�E%A�`�ĭ0�"O``(ǁ�=�PȑW#̣n'
`;�"OJ�zq�0\w����j��2�"O�M�眭t����%�R:�`Ը�"O��{�IĉA���� �b�,���"O�0!NJ��Ι!��:m�ry
u"O�C�C�H����*�^��,��"OE(����k�� �Q
|��@��"O�P)��R���(@k�44�N	�"OE���A$6<�|c�<x��q�"On�H_G�x#���"��Hc�"O����צ+Ԓ�+�̄9 �F �4"O�)�D�E�uJ����&�I e0D����F�*�N���I�}�
�)B�9D�t� k"6�!�L�(u��8S�,D� ��I)gqDC�&_�<�ҼQtE)D�xpE�ڊ0'v�ǎB�`Z���(D�4�pڒ(Mx�3���6^�����H9D� ;#���h�Ze�ǘA��y�8D��GY���Q1�k�|5x0#D��x�BE># Z���N�]�"X�'"D�(���7�Z-�W�'7����!D�������|$Q��;�$���?D�䫥��"1�¤A��^��Eh)D��˕��#�2t���H�,؈t �!#D���j�/+����a vL�,D�����V<�-z���-V�D�;u*D����H�	�hA���"�J`�A)D�ػ��D��B̪U�.|�1�(D�t5`T�k�^�;�IբC[��F"D���t�G2)�0UB��S�t~�A�ש4D�L�i���l�* �Q�/�A	�*4D�8D	�F�͒'�N�hH�ј��=D����T�h� ��̖P�e�6D���@���|�xE9�ω[���s&/4D�(KP�ΧZ���se�̫;^FY�1D��k2�'F���Db#N�r�4D���,�$����E

�gA�:c�0D�Hp�Ŗ!q��3�-H��� ��/D� DO�[�U �#		qf����8D�d:�!P�y�9`hǛM�2u�� 7D� ����o�x�h�Ǌ��@�i5D�`"��X*��ct��.�¼���&D��z#(�|xQ��ퟕ���eJ7D������7R��)b�]7x��芇�(D��q�JU�!꜋�P%z����&D�Ȩ���Kݘ[W��dLH�is�%D��:���rZdXI���\~ �*7�"D�\����D���iMY,Gk���'h4D�� zRbH��[�ЌQ���	=�h�J0"OEʕe�LY)��	3���A"O��"��7Hc +6�r���"O���F1y��+Q�N<]R\ "O�e�� Y�\G��cf#A�x��A"O�ٸ%L3?�q�"]�@���Z�"O�]ڢ)֢q�E�������5"O^u�2b�
!*�`s4�iwDQ g"O��0P'�8���Å+%��`"O�dk�aE#2�>I*�!�/�詀1"Ov�2D%WL���XF�=n�xr "O<�qp�W�m`'K�0l0=��"O�+����d�N���:�O�*3�!��4|���L�v���$�!�!�D�h��L��V��8%�0�!��:K�ԡPeV�%�f�	���!��5px���]���t-��Z�!�$����D�F$<�D=���w�!򄒦i
����_#��Smҷ_�!�[sz�Eb��]�h>�A��I7R2!���9	��,QS�+�|��Mh�!���0��t�vQ� �@�[Ȝ)v�!�Q)L�>�ҴݺQ���W�	;�!��#)�L��HA-jf�*6�]
tb!�F�W>� �!��tƊ���!���4r i��S�,J�� "}�!��L$>��6��2m����-m�!�$N57�5�e@Q�'�"��DhW�p�!�΀�F1�����P���W�Z�!�K�BI�� l�0)�^9�!�M�)�.���ʤAb"��ċ�4H !�)��S��&&I�5ȁ*\�s�!��&�b �2DP4	���3#�!�F�w�&lAp��T�F�c���V�!��^%t�D�� �Xb6<˓MM�r�!�$������Stl��L�h�!��ę>�q�)I1*��Tl{4!�d� �z��sI�zi�Q�bk��{!�$
9a��Bԩ\�=[l������=�!��K�(�� �F�)N���r#Q�_�!�EΚ<�*��)�k!�QxW!�P)Y�`f��kRY�pǀ�-2!��#�u`ch�q�����X/0+!�D[����P�Ƌ���`C%��1!���/E%P=����e�l���d�?�!򄕒V���r҃�
S�ܤX��=~�!��@*ĀR@H�,�8	�v����!�/��4ʶό R�:}�FI��9�!�$�	W�Z��C"A)'hx��V�B}!�$��(Uʭ�ah .|h���f�V
!�ɧB��� Gd��`eeh�!��}P��kј&�hq�F�R��!�d-t�|Q� B��\�~H3%�G#�!�$L�{R�h;�	��[��x2����}�!��I'I� ���\�{����$�^�!�D�<�2�z���u�LeH�d���!�D��} Z���EP~����E�YP�!�䎺'�`
`e�[��-S �A�_7!�dL�<G �  �Ay�0}��ɔ8hA�T�3�7���S�=K!��:�)qT- �}2D��!c�0���=?)�Oq��'W�P�#�&�j���C��0	�'K�x���M�B�����=^���+�O �m�g�'H�OB��)��"L����Ь���'W	�'fvTx�f�9����F��U�!�{��)�i�jђ���oz0���P�)�ў�@�R�O*�-��ő�����qdW����~��'z��e��+����&�=J��98��hO?���=���c��vR�1�h�z�<y� ��CJ1�WIN�oT"�`�Q?q��d�P�'�(Y��`L*����/�Ht���d9�S���$S��qgޱe���HE	������<q�yr��O�r��A��e��,8�ߍ8�ў"|Z�4J2v7�!-J�Ȫ�WM�bM1*ЧC�!�D�y����#�8#�n����ʬF�$(�	�<�A��!��P|X%+%	Az<a&���5�^Ѕ"Oԝ��Q�W%���ȁ-�\!U"O�!0'`�h��e� Ü��b���"O��A剚ri��d�J?�����D#\O�m��c�9�ƀŢw/@���'���'6X����E�T�DLh�C@[\���
�'T��e�6���!!IVR�j����D�	�0|��&�N�S���L�n$��� T��HЎ_r�ܠ6
�53d���b�1D�4��%�d����(�$_�fᄂ0D��DlΙF~��У��p�Cᣬ<�� B�jW,Y]�(0���[h�F��w�h�
�Z}
5Ƞ�c(��ȓs�p�ѣ�YcF��C�#�	��[E�u1q�]8U� �ViS�6��ȓzȨ�HT�@�GMZ	s��u��+��9�OЮp�L(��IET����8؛�p�E�eP" ҷ�ǳu����7O�\��i�j+&u�q	\�#��|!�_�<�?ɋ�)ϔs(��ɓ�$�ᩡ��_�!�� ���I)Y����53~({�^��E{���D�	�D�JD��>#�I"���C�!���Oh�T&@�@��@ڡ����"O����5*U�!!/�>T�u�6�Iԟ0G����NZ, �N5m�L�hvl��yr��:{#��t,
-l����f�I��y�.�	��A�u�^�p��C�?�M#���s�@�8��B>��̲�*��F���'��N�O����d�X T��p@��'���@a
4.���s��*k�\�`�'�X��"+ƈl�q�#��.�k�'"T���)�q�LP��c��X�"�'	�	}���ʢc��f �x��%-�d���g0��hO�өn
������= 	bф��=̪C�I6V<� �E�\��lI��;c��$?�S�O*��wF�9uE�D��n�6�@�j�"O��Vn�����B�]�Lf����g�x��?�O��s�=W498���
,�:�y��K�$:L�'%E�-�ژR"����'a{�߉q��ň%+:"����y`�	P*�t�E	�7���!Ac�h�<�G��?��[3�M=[D�iT#�l}"3�S�OWvh���ǣ(�|<�F�U�T�'ot��%
�7h���G,�8`�!�{28ғ��'m���KSj)YJXx�B��<l�ȇ��?�Dc�/u�1� �9!@lr��O�'�ayrO݁nf�5d��(g���V�y��Ӓ/�$!cɃ������K��y���Ox0u�eяH�Vi��y2���HF�PD��|�������yb�	-M�t��a��Lȡ#��y"ǐ�^��ԇ�#J�����y�h�z�&�x���nL�sG �yb�<�Vqb���0���� �yB&]�v�Z��'C�	4��:qjO2�y�쑣\��qUBz��9ҁ!�2�y�jX�'� D���H=q� �!&���yn7y���C�@@�^���"���y�
�^�����T�Zu�`I���y�lډ�ER�k��[J�5x �Ό�y� ���u�>+�P�gnͪ�yR��6ߔ`��<��jW%��y2c��;��m@��� �z���\�yr��A�fhK��U'1�iA��y�+ȯ�Q��.�c�tC �l�<q%��B����w�� �z����\�<B�'��i��Ϻ2���`��X�<7�R�-D�4cwM[�x���D��X�<i �5T��u!a�Z�[q��붧JT�<�5k!fq��(�#��8� )&�Q�<A�K&	o�0 ���E�`a��&J�<qu�&9�����D��~]�H��o�<	��>@���K�LȨ:�8� �!V�<!1��g5v�	�O�!�6XXb�Q�<�f�/j�t�d�kK�)�4+�M�<Y����l���D�A.u��Əq�<� �97���J''�9k+�|��E�f�<ٴǟ0?jl��1�5i�*5�I}�<	�"��lC�"�0N���i�g�{�<ie.�=\�P�ğ�&�f��G�t�<1�&݅Jr����N�g���{DBU[�<y�e�z^���A�(b���C���Y�<��&̠d�FU��l�
z<�q�sɅ_�<���L�B2�@&��N��e;֡�\�<� ��r��W*j���@	"6���w"OL(��㖜`��-� ��4Ҙ)C�"O� �� SC���Ҏ�h���3g"O�dZ��^�
e�\#$f�90$���y����-"�2� Z�8i�c�� �?����?)��?���?����?����?	��� ?�rS�іn✙��Ѱ�?����?����?�'�?���?1��?#Zǎxf��[�����?����?)���?�'�?���?q���?���B3*�H���CF\�	��#�?���?���?)��?���?!��?ف���E�FH҄�E&|4�4��f�?����?Y��?���?1���?y���?��!bJ(!�/�2q~���ᢁ��?���?Y��?���?���?����?�7�X!z�&���B�7}�4�k�▸�?���?����?����?����?���?�$�(��ؒ�g�//�&�@m���?���?����?!��?���?���?�u�H�g��\���H��x��ο�?����?y��?1���?)���?���?)&F�w���i�1u�z��2`E=�?y��
�4�?A��?����?���?��Y�9�A'��չ�Ɵ�& �����?����?���?A���?A��?i���@%a������G�%	�����?A���?i���?����?���?y��K�\���AG������ ��D����?���?����?9���?᧻iAb�'  �+�Đ�8>J\Zq.��3t9�0"�<!�������4F�:�ːF.z��U� 
T?�M�թ�x~�is�Z��s����4.�ʘ{�fg�x1�Eр=}�����iz��1,X�(
�O�����V�3&�`�N?��a��9NvܛG�
�_I޽Xs�<�I����'W�>�S`�ItH�p�J�1S���Qa#��M5�	h̓��O�&6=��m�Ɔ�"Y���xAB�mRZA�Å֦QXܴ�y�_�b>I��ˌ�hB��*&$v)[��5*�F`�Al�

��	����bm��f�D{�O�򡅁<�8�T�&΀W�H�v��Ay�|BckӢ�
��ƸK�@����b7�[�Λ�l�b�l��O`El���Mc�'U�I��HJR��;)D��C�=zE4�v���eƮX�(��|R5%ǰ[�����*[~�*�kv|�YU]�k�RD�*O���?E��'�|Qq'�� q� ��b��cb�x�'pn6M mX�Ɂ�M���Oi&�1��8+l@Zr�_�*	؈�'N7m�ͦI��b�h����*?�ѯ��8d�izS��\]4�HT%�?@b��Fe�5$L,5ˍ�4����'M���&R�6X��)�5͘T�'�:7���1OJ�)3���~��(rp�X�"������Ȃ��'x7���̓��'���S�.�
�JF�i�4�x֎ӽHk��0��އB��L�'���ZS�h��z%c�t���K~r��1Ͱ�D�ɲb��k���:&�\���''�'P�6M_�=p�X�,��I�3BK�m먊�B�f��?����'Cɧ��'��7���E��3m�Lu[��DA(���U�¦��3��'���I�X�!��-iϼmk؟2�ij�Eq���TA#d	0#.�q�	�����3O��Ĳ<	.O?�YC��'d���6�,G��t	� 3� �Mc.Fg~b�|����<Yu� ?�X��r��=aRi8 ��#�y�Z��۴p��f�'m��Q��D�yr�'��Tz��٭O�S�!�.mTrͫ���-8���:�aH%ў�SUy2�'D� e�ԮF��ە�H�u桋�'��'F�7��(�1O����ؠY�T�`�H+��%l�R���,Z�O��n��M��'�OG�������X�m̒dy<���%�X-<��m��[��hX�O�)Tr�6�Y�
/�$��[I��zP$�g~4��@�6��d�OH���O���)�<����&�m�� ��dU�V�2�KF)M����'!�7M9�	)��D���7�E�7uP#�<R��U�⑑�M�ѱi�u��.�yb�'Y:��4�!C�D-�G]�3"ٯG��0��_�Ee����t��'���'���'(Z���c�:Y��#��3��} ✑�d���4#ob���?y���.��d�Ȧ��4�֍y�P;(�%P�-��XLش��f.*�4������&���� �GN�H��X#I�;1X���2X(�䄁%����DU�R�^�O���|�d�V�Ӵ��&y.�`S O$�~5����?����?�)O�o�P�@�̟l�	�r�Ƶ�U័�̯h�2`��	�]��N
�I��Mt�i���d�>��H�Ð��7��ͱ����<a�<�U C*8H��*O��i��O �$����O�SF��gY�CO�+S�P=�3n�O���ON���OT�}λ~�`��
�L"\����0	!���7f�FA
'���঵�IE�i�E�����t���,��D� �uOz��4rɛFq�����$4/��O� �@���h��P��d��ϰI���M�б�(ʄ>��O ��|*��?���?���..>�BfP"�����D���x3*O&al��T��П��	i�Пp�c��xq� ��7S!| [4KY�������}��4b�����O���	U+�pSՇE�6� �g��*\&a�R��,d9�ɗE��K�)ļ=ܐ�%��'d9���	k��w怖K'���'�R�'s���\� �ٴzGb�3��h����A�q/`����	]����L'�����G}&oӦ4m5�M+,ȹFz Y"�_3	5���=X��<˰���<I��p��m��E|� y(O����� R]ʅ�,y�bI�5I��j���=OB�$�O����O`�$�OP�?iH����<�a���d�ܡ��Ɵ4�	ߟ��4R.|E�'�?�W�i�'8(u{B��_:�1��n�)8���X��|�p��m�ş�r@U�a�h��ʟp�J$B�����_dB~a���K)1%�D��!j��i�'�.6m�<����?���?�1�	O���UiϢ`�8�tA_�?	���$T˦:�o������`�O�2�PdT:�MZ��&jr�O��>Q'�iT7-(�4����:a�`N@�LN���2}�ġ�T�7��x��"�<)���z��2��L,���{"��3 wzy���
�A.�,*�Þ
�?���?1���?�|�,O� l�%.U���O��}�����eЧj�z�*�m-?��i��Oz��'r(7T�[)�M4#��q�JՀ��ˊtb�oZ��M㑌�84 u��?��=��5c���9P��A�`��w�� �=B��d�<���?����?	��?�,�bȁTje%:�3� �D�D��G Ҧ�A)���	؟�$?	�I:�Mϻ�ҵ��&̘������Ô�N�%����oӞ�&�b>���bQv�	�%�ၐ�H9���S �ߘ��IצE�D���3I>�,ON�d�O�i�Ĉ��VjH��A�0Ŕ=����Ov���O$�D�<A��i$]� �'���'�V�8U��?�b=��M�O$Ĉ���J}R�i�(�n�v�Ɇ{z8r�E�?a�A��ϔu���I쟄���\�%o�`G)AVyb�o�Qɒ��u�h�	qj��j�3{�����N p���	�@�Iݟ|��^�Ocb�js�LR:�1�BK[�eT�,��'5�6�MYZl���OF�mM�Ӽ[�GN�%��q�$g	$��)	>�ɲ�M�2�ib��	�^��ȹ�'�f��h�8�(φjM��ST#��6����$�'H8D��P��X�4����O.���O���OZ�Ȕ�F��1�ʓy#D,��.	�	9��3u�f�˛pK��'�����'�~���2p̱)C`M�o%�m�� >�պi�@6-$�4�����O�8��HS�2����VJ�>c$lq�(Qz9@R��O��3��c���b�2���'�Vї'S䌸�F�<+�ll�ǆL~B����'n"�'r"��$W���4k4�A���d\���B-�5(4D��b^����t����J}R kӊmZΟˢ�6qM�A�D�gv`��$�;~_����p�P���L�*|Y�ˉ7r$�I�'�0ם�߹�UG�By��rT.4uz<)[@'q�8�I� �������۟����c��ӌ0�I�E��pd�:�?����?9�i&�;�O9�%u��O,�ؖ-��l����!�z�`�L2�$Ц	`ش�?��˗5V�j�͓�?�u�3,$>�"р#G����V���}f#�1�1j.O@�o�py��'���'��c�)(W����DG�Ŗ�Pb 0	%b�'P剄�Mg-��?����?1)���k�:�𑮑h�`�a�&�u~ҧ�>a7�i��76�4�z��(_6p�S�3w2�Ǆ��N�6�ҟ4%�%;�<����ҥ�3wP�ʓ���G�@�<g� �3��\��/�3�?���?���?�|r)O��o��?Ҿ��w�ѩ_|`{q�^H�dP�
�ɟ��I�MC�B�>1d�iMV�і��.,���1�'v�$��f�D���6'A����8O��$U5cMZTX4���{�˓=L%˵�ӓBH�Q�Ё�,yod����i��	şd����L�����Iz�D����sq&L�;�x �FY� �7-��G!����O���:���O[nz�P�z@�����>.� ا��M���i)�O���(���	��'?O�=�G˳/�iSee�O���u1O�<��C3F.��� �Ĭ<	��?1�C˼ F���(B�}��������?��?a����d�Ʀ!Z�$������ڟ88ь�¬s�g^�r�b���  B��v��	?�M34�iI�O��[�)0_�0K7�.w���s7On�$bӎ�)2Ǒ#}G&�'4�tnJ{������'���"��V���{Ӎ��?B���'4��'�b�'��>]�I)�T���3��a��%�2��Ɍ�Mv�Wr~Bnm�l��]:EB� EGH5xP�U�6�P�6��	�M��iز7F <o�,�:O*�$W���� 0�������Ⱦ>�J%�֪�+n\��2�7��<����?	���?Q���?ᖁ����	�*N&
z�����DJ�� �??���jJ~��0a-���󫋳���%A�c��	��M;��i�&O���$�iE���0��@+ބ]Q�
l��H�*P�|��I(�u�4ۡ�^$�l�'/��5���|!��F6I$����'`��'2��$W��`شe���la��*�߲JO��W�9s���̓t�f�'��'l��g�f"}Ӧ�m/[����Nҝ*������M>� �F�ކ-��������`傀P�t��2I�My��O�n�2s��l�s�R{�Ѐq�N$")���`��ݟ����<��V��3�tx��L�.ؽHS`M�4�f�͓�?��)?��G����ɦi%����@�D���%�D�U�ʄh��ߪ�?�OR�n��M�'c���a�K��<	��C��A�����ibv�Yՠ�>/b�� �?A2y�F������D�O��d�O<���	;��J���e�|[2F��>���OD˓0�v̈́�Lb�'�U>��u��![��yC�[���`�u�7?�W�`(ݴ{����6�?�j�GhPJ �ч[�qs�젰��妥hU��21(�j.O�iG�%04!`�_%8޺E�>Ӳt
�+	�����Z�S�M�z(��!d0A�N�4�˄�=%����n�|��r�^(0F�RAĕ����25*֯w��#?� BW
 ��hƯV�W�b�3�l�Z�܈u&�:d�U���TI8�Ad�΂BS�x#��U.B<З�* �p��C�dAr��> �X A�<��� ��T���o~�f.Y�'��=��B��^�h�1d�w��ҏ�<�Y Ԩ-3��:dզ���d9�H9c��Y�:;Jp�	�2Yv\䘳�D0
��O$�� �d�O&��F3E�
���	U��z�C��۰��95��O��d�O��O6���Ot�DB"W� �Ā���b��R�~��![�C�xmZCy��'��'���'��ZF+<�Mcp��>p���"�ǘI�D(���m}r�'|��'LB�'��ek�S>%�I�}08]���W	4�< ��={�,A��4�?�J>����?9'x?�e'����&�1E�r逡e��tХ)�Ga�Z���O����O����O����O��d����ĉ�������{� kQ)G@�	ϟD�I���+c� �~�2-IN��лW钐Eh�PZ�c
��!��۟0@ ��ȟ$�ISy�O1�i��R�O��H�فH�hP �gӨ��O�ո��]�r�1O���,!��B�%�؅A%hT�eӄ�V�i�5��'��\�L�SGy�\���$�@FO�hK�h�02d�(���M��̃�����<E���'k�z�D�J��L�=N��� &jxӨ��<A�+�3�?�����$�O@���4�L��L��T����\���$��yRʓ�2�����On��	sC|U�e �	"�ċA�N E�hPmZ���!�ē�?a���� ��!2���΋_�����QQ}�'�ט'��'"T�&�G���7E�����A@R�Nq`x�'��'l�|�'m�@�oZ�Q�C�+�8YFn�SvH%q�|B�'L��';�	��R���L� c(S���<bU&֚q$Yn�՟t�I��D&�p�	������>�t��'3��$!P��i��cw}R�'5��'��I*|�(�O����Z}�\����'��h9/J���7��O�ON���O���O�2_���I�/��ap�Ì�x��Aw�.�D�Or�(��D�)�z���OX�)�26���-[�����5n�> $���Iߟt�WlJF�S��b�H:4��k��'� ⅆ��M�(OT-@���O����O���|��C�'��`1���H(K��b�����I� i%�S�QD���ČY��{��Ϋ~�l��?�I����ΟH�Hyb�'>2��#Lf���b�,��9�M�6L|6MʡqR�"|���=3���G	�>� 9:��u�w�i���'���[):����$�O2���GV@2V�ٯV��ȱb��{.b�ġ!WD�ٟ��	ϟ\y���ް���ϑRJ8*X��M��H��!+Op�$�O"��(���,�ِ/D@�܂	H=r�d�dQ��B!/�d���|�I�'gڸ���ͪ\ь	�P����t�2�B��]�������	W�����	�rJ�Z��P0Z 8�kKN�1@:�@�Jj�Iȟ���� �'mN�۟2�Q���X*eCP�)k�)��i���'$2�|��'%�a�:�Ą�G��h�Q�[{�웻I=�	����	ҟH�'HBpqQ_>Y���F/��;�ɋ�
���.ĜW���ٴ�?�I>���?A�����'�:�(#L�0%B�'[L:rL3�4�?Q���䓠 J�'�?����2P�Q.+� d�g*�\
�!�3CQ�g��'���'?��I6�T?}+������Y�1Hچ�eouӐ˓ND�|����?a���?	����Ɛ8be)ɺ&�ʍ��_�0��2�i���'��lf���_�LZ���s�˓>��*�!�r#�V��X�(6��O����OR�)�E}BT����	�#\���͛�p�.����%�M+ I��?��Z~����O�1H� ;A}��rĀ�3B�C�����U�I���I�{���O<�'�?)�
젭Xc]�<o8IPQ��-QU�0�i`��'+�I���9OP���OJ�DI�2�"�%�sɣ&��<1����Ìs�*���]۴Q%��S�`�IbyaG� ����ANU� �~` �M�o�7-�<�����D�O����Ox˓_��h���*
�@�5#��j-�[��C5?�'���';�'��i�A+���J�t�ԀC::B0*�Aj�8�$�<����?���Ć	xj�E�'E*��� �Q'bE�p��j�hh�'�'w�'�i>i�	���������X����&
�LZ�O����O
�D�<A"@R_�O�@]�a�<��Xǈ��4���l�n���O˓�?�)�D��1��C�=�8��@��T%X!(#����M����?9)O�91�^���s�=ӅΉ�����@ǹH��ˁ�'��<���?�L~�Ӻ�E>i�r��u�SE�6]9�M
���'�$��j��p�O8��O���J�"�1t���+�- �W �L�ldyr�'�Ҁ'��>��i`�X�OъX�:�bv�F�2j�L��4,d b'�i�B�'WB�ObO�ʘ)�J}�r�haDH�D�!+ƅl��,��ß���xyRZ>��O��������h���SS۲�x��Pbb����O���̀H�S�Ԓ>Ql��UplM�/�*<�xAǆ�n:�$��4�'��DB&uR����ȳ_�څXp��X��6�'��H�[��r���㟬�b�V�)%$<aq	���-�gO)��� :궡CS��O���?I��� �9��.g��I�pl/%�4m`)O����O���s��OS����V�T�q��#�B�KV���2&&�	ٟ(�' bb�F)�)E%Y�`���P�r��z�EP�����'CB�D�OJ��α6Ҩ����� ��а�ɞw��� �&B�apP�x��'���Ɵ��1L�}�D�'��"�ɹ�(��C���M����v�P㟠�I���WI�5��O
�� T�}�x<��(K7 ^�+�i�R[���I x��Ob��'�\c_�HٕLŊl���ڣlK�>n5;M<���?��'I�VDlT�<�O�ĩ��À�%^Fi���Ұ�ʀZ۴��䚔{��Plڻ����O6���E~�mԖ>�\�jD
���\1�����M����?R���?���D�O��sӾh���ڣ]A�0c�b*�����i6Ш4�kӂ���O>�D�6t%��s�����g�P��0l�Z&FP��dӤ��0�O����OV������g~�
Q:b��7�Y�0L"��÷]�>6�O����O,dE�
G�i>]�	՟dS4hU�K�E�3B�� n�Eσ�M��?9�K��qQ?A�O�r�O�l	��:"[�zD/��1h�[�iQ�0G��I���)0�	�>��<:C(@Q���.]�n�H\��O�u9T�;���8�Iʟ��'���d�;((p����#�~=Ij���0O��$�OV�$�<I��?uBSy(TRb旙<���Żb��x$B�O���?I���?+Oz�Z���|�Ҧ��ww�$�w	�-H*�j�&�P}"�'�r�'���П �	!����O������6$Q��UI�J#�O��D�Op�d�O����!B�nݟ,�i���!���~	��hV��r���¦�������LyZ�M�4�ϧ�򤰟\+�I��V�1`�E�S�5@��`�N���O��D�O,��FN���I՟h���?)��iX�6N���
b V`!�*��M����$�O���!:���D�<���A&��K<TA���VoL�!��|���D�O*��&jW��I۟�I�?��lJ2��A����
|�`��( ���OBA#4"�<�(O��]�+��D;$*ʵC9 Pį�(^�6�Z>!��HmZܟ��I՟��S�?�����|�I�#�4�@m�r���ٗ��:K`�\�ڴH������?I/O��#���O�\�NZrB}!��R7o���pӡ�ݦ���|��3G�$ԡ۴�?����?y���?��P�ڠ3�lї@D�Po�Fk���'��I4�v��|���?��6�(�ZV�Qw������M 90F�Ї�i��&֒; 7m�O�D�O�c�4�O��y�%�
�V�h��R�¡X��0s1O��$�O����Or�døh�Tt{sA�4A�.����0]��2I�����4�?q���?�]?u�'8�������GS�o��� �_Ҍ��'m��'�~m'�'���'l"A�w��6�T�o�����ӌ5��H�C�V��]m��\���<�I����'��E^6���Ǘj���īI%p�|\1�ϏS����?Q���?Y���?��D»=���'�2ȋ�⥘φ x�^p��9M�t6��O���O~��?��&��|����~"���m��Dh%HА K�-˂�M���?��?i֠� e؛�'J"�'I�$c[�f���s! �L��@Po?t �6��O���?A��G�|�/Op1��&�E<i�2��lL�5eR�`���M���?YQ͞�o/�V�'�R�'�t�Od�@ڕc�������p���;����?q�S��?.O~![�=���O�|�`�f��@�2���Y����4,2�Q뗲iER�'���O�D�'0b�'q�����z�,����)L��@�'l�� ���O.���Oy�0�������΃R�b���dX5K��$����{�9mZٟ �	۟��WF@��M#���?1��?��Ӻ{Q�<To��HC�_A�f�����٦�%����Jv���?����� $N��0!���7p�iI���M���_#J�QǶi[��'���'����~�̅1|�fpsN˄4G��[1"�����ݙx��O����O@�d�O��$�OD�K�'��Q���AU�]�(1� ���4s�$oZ՟l��ן��I�����<��ct"��m+"�K�pp��
����uLD�џ(�I���I����!�e��M㷍ٵi�Ԃ3�O�f�Q�,L;P�V�'y��'��'�������~>a��*��m�*�j�<o�¬ˆ˖�M����?����?ђ^?������MS��?��!��df AF��������Tԛ��'��'���ҟP+�j>��'�6u �@3vp��!��]>���2�`��m�r�'�"�'�|����`���d�Ot�D�BPD�bP ��q�F�~<,ld`����{yr�'A���O�bS��s�N�B�	|P	��.7ɢ̘`�i��ɓu~�DS�4�?	��2۴�J�\��݂&�v��ԥ� �9%V�p�7��O��$Fp���O.���O����V�0�@! �BϚL���4rg\�2"�i%2�'��O��D�'��'�#�k��K����PҎ'* ���v�(��W��Oh��<ͧ��'�?�c�F�H��,<�RmR�ǖ�#���'�'�����t�@���O����O^���6P�1�U�­�i
��aT�i7�'�x�⟧���O����?�h��P#s�(Ua��!)�B%Ilt����K$i�Йl��������	>��)����$1�,�Ju"�B�4	���>I���<)/O���O��'�?)E�]1>��B�]�<�"��%�18�(#ֳiC��'�2�'�z�'��D�O��Q3%DL�(���W?�lٙ@�ƌ/V���O|���O���O,�')s(-��i 2@J�aV=sQ*d�E�ݎU���D�d����O����O*���<!��F����'����%�6�X�e�Uw�[$�iAB�'���'�D�D�V�XR�i?"�'H�\*�(L	z�ʩ��D���RR�c�����O>���<I�~$�	ͧ�?9�'p�`i3�E�bH|�P�Ùr�a�4�?y���?1��b$�%��i��'n�OH�\
�̙�qpR={a�� ����'`Ӓ��<��>���'�?���%2���� ���J�*JXQ������b,��i�B�'�\L0�p��d�O����V���O��Z�ϒ8Yx�a��p�ء��t}��'�\QZ@�'���'�B K�OT�'F�H[GG�z�t�P"�MG�ƈlZg��`Y�4�?y���?)�'Pȉ'bBD�|t���'��?b}��g�<� 6͋�l�f�/��.�S���HGfF/.	��`��\7��u4���M���?���@��(���x��'���O"X���X�t�����@;�,��i5�'��l����	�OJ�d�Ob`xF�"]OfT�j��dq���ϦU�ɋs@���}��'�ɧ5�@C��^��A��_��#����L�sRD�į<����?aK~
� I*HU��r�aP s�����愵[�t�Bc�x�'���|�'��dڔ2�d�.�'v��u��&���@�c�'��	ڟ��I埰�'ʹB�Fo>I���J:䡱��`w�Iapb�>i��?9K>a���?�'�Z�<y� Տָq)㎛�>�~D!�T���؟���ß��'��JU�<�5Z����fĄ�5�d+�g>�"8n����$�@�����1"f�\�O�0���y�( '���5��i��'�I�r1�]XJ|����z��^RX��E	$^�,��@r��';��'>�d�'�ɧ��A�l{.i�ਂ�C�1o����]�42OM��M3BZ?q�I�?U��OI�͏���a�B�~��X[��i���'f,5 ��'Oɧ�O5z���
��JqK�=P��۴�@�t�i�r�'���Om(b������*d)�b2���E탻�M����<yN>1����'V���g�<��#��S�
ò��F�fӨ���OX��S�$Ҹ�$������0��z�t��g��YEz�+q�^:f��(m�C�	�=�t�)����?����Ƽ:TD��*�,��ɔ<�r�.�M{���Z:-O�A�OxB�|b�H�v{�sG�� B�hy��i���?%,��<����?����?���[ZzH���ia�q!r�.��YB"�T'���Oj�$�O�Oh��O��{D���Z|p@�*_��P�1��� EƅR����	�����Oy�.)Mb擯%����ug��n�y�
T	 �j6�O��$�O�d;�	% <�*fx�@��R
wZ������'a����'�r�'�r�'=�e̝*����葯��VnvXX@h�?h�8�H��(�M;����?1�QL\(���X�*�b� ��P$E�p#�a�	1o46��O4���<�@[$2�O�O�b`�&�U�Dl�QSs'f�0`���aӦ���DW��3?��]�Fc�`%p�nL�|��ݓE�j���O��*a��O`���O<�D�N�$�OkL4� ��%�ݸ"D�ps��-Eᛖ�'�r�͐�O��>B$�&�H��/ȭ@�L�S&$�;,LlʲWa묄R�J�1svJt��Gé2���w�#_Ϩi���o��`�,͠|ڬ���O�XV�a�[-�y⍏�� d��"	F�26��5�JX�a`�N
�|2 EK!u�b��/��:��H��,~�D��!���p��y���;`
[XǞ$��Ƙ"K�RA9g����� �N�9XA�����m�<{�\D���#U�](_��yv	P���\*��F�-���8`�Lp�H?t+r�'j��'���ȟ4���|
�F�d���y��<t��[��Q�/����G�P����>A�����O��z��`���Q<�A���y�t�ѴF�-��9G�J�����ɷͰ?�!�!� X��.�,D.�uB���q�<)t��6R�� �N�B��i0$i�=��O~���O_}2�'ƒ�q���F��ܓ��Q4r��'}�l�O���'��	L�|����eJ]��^)sT�uӦ�$�0Rb��V
Q�r\B,a`�'{���W�sӊE R���^��6��Lm�H�l�0v"�a��'��p<�-���@��Ry΋/L��ن}%RY�7�͡��'#�{�能W���V�zx�K����x|�����A6�>qh��p��T3O.��x9$�i�"�'��ӅX�p����}��=P��ѲG�]��럎m�$|��۟l�F'֝}�$Y�O��J��m�S��S>�:6�M�u��t�2䕀"��Y#�?}B@D7�9��	�l�ĵ��)6���b!A��)̲�_ ��R���	��M��i����ƚ@
�����ˌ�o��X#��O���$	S������
:��Ĳ�J	@�axBi!ғH�
m2a��$j���q��)]�f`�5�i-��'s����D�.����'[��'���w�"�����)"5&�[�K�3y�n	�b��=i�#���O�����;8�1��'��側ȁV[Ű����kƀ�PR�R�n���`U�O`��%
�����r���T�Q��i��A(l�&8ae�|�gA(�?�}&�ܻ���lBf8�i�Yn�R��(D�(sw��1o�:�q��:J8mȷ�3?��)§Rۺd�Ɛ�,\ �C#P�,�g�9U��}���?���?�������O��S%�ĹQc��E�ȭx�ƓN!����Ɛ̰?Iq�K7���2�K��23TP�"̪B���_1@�B؁�I?�&`��I�G�n\�&��8F��"P�X
m�n�O
����"!��1�� �d@� )>D6�C�)� ��p��=lB��!.I*�
 ���j�-:����i��'*"|��A���x�jՈ��ZE�'
҉V-�"�'d�)�1�U�b�ە(g��#6�'C,P����/>��E)�_�O��Ǔ"�&02�ģD�樐VN͟ ����-qz���b	�8}8��1OT��A�'�6���-�ɓC������+hd�Hۗ��.x� �'����
��[�D�b:8y��KL�B�ɵ�M6ꏈ|���%j@ iنHɰ��<�+O@p�偎z"����O�˧�<�H��H���S2I�A�T�ےE͊Q������?�D�ȠY,h��Ȉw�]R ��;p���h�d,D:йQ@EI5r��Y���߳��I]�@���c��w�d99�eŪxN��~J�E<:g��z�n�F�
���o���-d��-���Y")���jd��G�̥Q�AL�e�!��^9��f'(w�@x(���{�ax��7�[)��!�Ǧ��xb�A��
����i���'��	�-��m���'7�';�w �h���Q��*�:�A���>JU��D	M�q�DBo?]1��OX�"�LYa݊%�VK\)u9X��h�2b�J�`կ�)W�9*T��7�q��O@���7k=8��
L��Ĩ3��N����|2B�.[��hk&n�&.,��9G�0�y�	Z�H��$hY=�=c��V9���M���bq���`�C?*mP�)׃1�A
�@�O��D�OR��ZպK���?Q�OH�t &��A�)k�G�B�HL���G�xrj�Pc��,~�����^
z�`���'��P�I��VL 9��B]�x�F�Ɖ �?	��'D����Խ>b\��6��'����'��p��p<�I&����y��>�I�:�U���������h���v����D�Æ7�"u����0���X��X�I���ܺ_���'�`w�G�8ܙ����-
���O5O����&F�z� �%"lb���_�S:����_�B�p`��p<9bN�؟�����M���_�	���(�d�U�W<:b��(O���4�)")O��BM�<ZY�ɂ�j�~�4��uO��nږ�4Y�S�>bXQ�`�	�,��ٴ���"}^Dl����m���Z��� T��p��D�|���S���'�����-�0=�1O�3?�6�\?H��suc� '�>����{�w*(�s"C=G��Mz��~�O��uh �؜w�(0����$8k:��I�L@$��ORp&��?M)%���1�0x�@�)"������:D�h#�CG�Pz0q�����1`e�8O�xEz��T�a&�Õ�X;6�"hQF!I{�N7M�O��D�OT%0���	2��d�O��D�O�P"+<���tl��)f�ԍw�%��P�A؍6c>�O�Eya  ���Y�o7${�q�чM�ɦBq����|��\(l"D��憱uO�$��n�'F�ʓO�4�������k*=(�	�x���[�XMu��QX�Y�a©/� JwM,,px��'��#=E���W9P��Q�	^�:<,ܸ��-�P�ID�H�C�2�'��'��]�d�	�|z��.����e��T]�����h����F�+G�P�x���V �'~c�hb$F�`<��E(��w�;w?T`����)��	���?!A�Vx�$@"�Y�X �4(�	�S�<�d�V)_},��$Z+�t9q�/{̓r2�Oص�`	�L}��'/���#O�ZI���D��*m�5@��'�ҤXE�'y�)Gc"�������t�	taE�_pٱe� >2訛��$�B�Q��-�,`t�`h	c0$V`�\������8
� q!�ЮT�T��A�knF|2a��?�����dM!o����r�F%�N�{a�߻r�1Od��><O2ա#�:3��84HB�ybO�(nZ�Q��h���.T����f��# 9��nyB쉛��6��O��ľ|����6�?�Cr>�(+D�"����n���?!��Zv�������d�� ju�[G���hP�H�<��ɏh\�#<���J�)`L yd�O4?�ƅ���P|��ʟh��'p�O}�O�8��
�`�Zu�ˣ�JhP�yB�'��y2녊P@�u��N����eE�0<Yw�ɡY���Y1��1PfX遑ؼw��<�ݴ�?����?����]v�ys���?���?ͻVV�B���P~��M���<y��94��mT�'T� ��7�1�0O~��ʘ�~�P�B��&|8�|:7���5Ɍ����7-^�ͺD�ŧASq��O���f~�މ�4��DT R�Ş|�	FT(���|�ˠ\�J�{��̄m�BTRU���yb��2��-ʤbu^�1d/ɠ��ąk���� �	�DjS�&�İ����9`~*l���%e�@e3�i�O����O���ǺC���?�O�J�
^�~ӆ����`IUq��ӄ�x��S4���r�K�b���闒w)�t�
�'��尦K	xDN�j�!Z<x���U)E/�?�V�'����p�M�e|���F	((����'������g#V�1vK�s,����y��3���_�=�ܴ�?���-â� R��H�ڥl�6�D=b��?	���+�?9���d�_�2|9+��C�#���c#�X��d�U�TBs�P�隫��0�'�u7gC��v-k��X��#� � ���o��}�v�\8�L0g �O̼&����녆5��,�ƕ�/{j<Z��?D�X8p�EKR-Z��@+ON����=���ߴ)��d��N�L��D�ʄ3�� �<����7��&�'�B[>��E��ן�j�دV�Բ��W��$�Kv�Q�|�I)Ң�H񨌥]����)�|
��S�b��`c3@L�<�0ţgn^\��I��-3���e�)�S�Hk6��"̵ ����ڱe�h�'@ja���Lʛ�r����;�Ӹn�=s��^sD��6I�,bddc����fx���T�'1y�8��� �*m�b�3O�tFz���� Y��3w��9D��Y�l�aQ�'d��'�����KN����'f"�'�nם-��R�-�IΖ���� 9���0���3B�B���� ����R�g�ɸE^�!'Þl4��5aĞ1��1�RF\�'2\���{|�|�;�3�$S�!մ�����1�.�q0��*e�$��Q0d�Oq��'<�E�	׮����d�&q_��{�'��tY'�F�j�G�4�~��O�)Gz���۰~	p;Ĥ�
:s&O���vAx���O���Ot���?������g[�xX���؄4-*�"6�P��,	�޺Y(�yA0��.U�5��GǒJX4Fy�^�~j�YRX�{�,�z ��+^�Qy��F	s�Ѳ��ު0wh���M~�DEy��K6]l�e-yY2vB��X,�@���a�%6h�V�ƅ��I:ت�aݎ�y�� 7�B��e��$r�,V�)��q�<�����\��o֟��I�
�|���g�*z|�9B��P˖�I�X�q![��	�|�f���&���t'�`�"����
�5Ce�8O]�3�$��]0�
��К2��2/�*��x�� ��?�w�x��F�r��e�55 Igo���y�Ƭn�$��R�W;��*wbL��x2�y����ƪחv�l1�3,L�v��Q���$�w��UlZݟ���k��.t� Ps�y�D���ƹ
��Z2�'Q���sh\0s��3⚰gB�T>��O�� ��%�`��G�2Pą�N�L�#;�r�2��G�D� ;�D���'�Ms"#����N>��F�)���R��)�!�M"�������GZ�B�	�J��)!���/��_����~�'��HzR��n�L��⡋�y�,Iөh�<���O��PN�'��O&���OL�4���gU89Pډ���-3�X�Ԋ.�I�ݐ���S:��v%��}5F�٠LD�6?qOh�1e�'6~<`��G�6�*d�_�d�8 �_���L>���%Oh�׉� 2V\��HS�<a�� BftA��s����L~r4�S�O���Qb���:��q��EG�8��������pd�3�'��'��ݡ�Iǟ,�'T��hB"Ô1�Y{��[(�]4:N�����PX�(P�A�7<��)�`��N�,84���o|y�`���>���P!���0GU=��A+1M�m���Ʌ��?Ƀj]#I��pKD�26K�L�ǘK�<��,9o4X����B�m �Z^̓=�Od(�6�OŦ=���PP&��_�� ���3n��c�h����t��ퟐ�'|�<y�	w�I�v�4���@�c?��{@R�L����D�85A�O@|'F͚>�d��T��3zЩ�W�'l�l��ZΉ'!�ᩇJ�?���c�+�>� )�'0�����F9����snG!�h�	�'�p7�5 "Ԁj�$ْY�\ѫ �'$1O��9�FAӦ���ן��O1�H��'9Lh��el��sW�_�	3|�A0�'8�&Aq�ŀ2�9�T>ɔO��y�H��� D�[����0O�\���c+(��b,�)D�z�]�%:��5�9G�&��`M��f���O�]"a1O��O�X�(Ɉi�<MQ��U�r����P"O*a���.����P��M&H r�'�"=9倾x^ �Ȇ.#&��S�<PQ���'N��'���s���{,b�'&R��y� X�S�Ȁ;x4ZE *ٽjY�M� ��.\��p�'�t�P4�������L@|C� �J}J$�[� Di����#3�I�X��8���|b͝;�x�W/[>P�����%�6[ޓO��ڠ�����1@N�d[W�8��-A !��D��t8Æe2й�� O���'��#=E��N
+I�rP��+9�B���2��}��oO����'8��'8��'���'�r���@�);
��ϟ*h$�r�mK�{g\*!�T���c�.<O��#�` 9�����6b����U--�)���\+�݂#�T�5Ԁq�Q��2Qh���ė�23�)Uꋀp�V����[��\��'��$�D�O���0���O*Q �O
$X��dH @�脪w1O���D��x��AX�Gʠz&X��7iȈQ(~���ƦY�ɬ�M�"�i���W�z���4�?����.h�tʝ�\����$�TQ���?)d����?����.��pf�'N�8AT�ј�)ϮT0�%��������}p�KU�/�J*H��σ�\?0�D�ً�fW r=r�j�C	?zx��0Poͣx	v�#W�'_JV8:L>��0L<	�@�&M:�ZE��py�4���^L�<�B>2���ʑL�z�|y�YG<��i1���r/�'^�`C�?|�<�(�|�m��~�>6M�O���|J��	��?��@6�2aKp���6�C ���?a��B<�C��<6|��i�M1�*��' E$@z��I�X��1M�M�&�O>�r �7z�͢��|����3ge�Q���;a���өsh�|kQ�M�Iq��`��V�I��'��TQ��'�ɧ�O�l�K��&�Z��Q�^�S����'��(��GB)1k��QJ���Ó@푞�$'�m����#L�"A�����=�M���?��.p
F%��?����?i�Ӽ�r��2 >��6L�-I�D����9:�B���E^5\����7^_$	���L>gŕ�w�B�F���$���H�Iv�ed��0\�PR*ñ*�d��t�[w��Z�c'6ɰ�w�Qi�#Z��8a��T&r[e(�䘳T"��L>R� 1=K�0qs���iO(|�aM�g�<�%���t̸�{"ŀ;X�Q��SO~�;��|�K>���-&��)����Y�<Bą��X$LȺ��Ա�?����?	��%��N�O0��w>�I�-�'��t� k��/�]������y22JǞ�T	�3��8�<ɖ�Y��`�Z�䁵$��s�dRͤ�R�n�-T��Q�#]36tY6JZ�� k�&+�v��1eף}���$"�@�I�`K�O���D�&N��A OL5p���h�o !��]�P𧌾Z��yq��#2^1O1n�c�8�jܴ�?���?t( x�"2���,�Dv�I���?���-�?!�����$�:k�a���F>t>8�L��$|��%�8�Iv��(!r��s���\HD�ū����@h Oal�pmS�s�t� ���2����7�6��-Y�"�J�X��l�OVdl�ٟl��z�RA���$q N� ��Щca�Y���|�	ğ�I]�SO�	�VA�9�5BelZRSC�ɫ�Mk�H�!,1�}�'`�4o���p�N �?a.O%8�D�զ�Iܟ �O)&u`t�'���򈐲�*��E�Y[�E��'��J��)PT�T�S,���h�O�V��5^�>��#J[~QtѠ$ƀ���I'�j��B�G(��U��;	���(�3.�Ա�f�޺�C�7~_�)��NUdԱ� �~�$W������b,�q��D��Cp�p��m!�dK3o�hzU�@jΙr�I$�ax�,�$�j`h�$�4Ɔ@���%jߒ¼i���'*r�Z7htx�`�'b��'��we���9Kۚ�9ӌ���������w��]�WKU�ne�c�*d1��O��#��X�+�xĐ��`�h���8E"R��	_R��9�Fɘ0<R���xB4i�R���H%u�0P��eO��O>@�������1|���lR�6�HK׭t],�ȓ$n�p��׿jb�\Jqo��n�l��'*:#=E���]�{�.ˤ�Q4��͠U
ém��qTn�+J���'���'�,����I�|��Bܦ]���4`H*S�*���	WH�~��u�ЈXETl�N"��<�m��^����C]*j�)�W'��9��m�F����<񡇂�#,v9*��7����U�u��Y�	R��� Ղ7;$D�i6d��*@"��� D�t��h�.c{��!�Ɣ;g���j1h=�I���'W�P�df�x��OX�ʓ�ԇ����@�	!ό1���Ol��^�99����O:�H�"�����7�@��p8O���ĢP�z��Pp#�vn0U�'
4�L�h�ٲ��<��͏�0+Ԡ"+��88�4Dq8��p�
�Op&�[���2w-��x�o��_},|���(D��!*��չ��G��$�J��$��j�4F���q����>2&Q�J� ����<�K����v�'q�T>Q�sB��B�ؚJ���ɖ=x��T��,�I4<��I�pa�H�S�tT�� ���c芄$.��jF��ٳ�>�q�ٕU ��<��1�H�Ha*U��H';:�B��u���Nr��+��	V�U�ȉS�� �Z����W�+�!��6}�E G����|�����&2ax�=ғX@F�#��Ѡ_���R��(�b���i��'h�BP��
!���'���'9�w�,I��C�<�0)���](?1�A�D�3	U�y2�
Gjƹ�f��
`�t�P��'Bn���A����/.}j�i���7:l���|�o��?�}&�+�ɀ�)uNd���[��a"N<D� Q�!�8$
V�bɥ/����T�>?��)§m#B-�s�
�x(�8����mfv�о sz����?����?�c��n��Oj�$t�V�� V:	h8i��Փ>q����ٻui�%�r`-�OP*`䍎N��EPDG�J��Ssg�'"޴���ڔra|�&?2�\�V�n���I�]�.���`�aR�-BL�Y��3U0`ٷA��y���7�H	��i �1k��ȝ��'�Rb�<l�=�M��?!�IB����Qm�5�u��'�?A��`���?��O�Z,[���cLU�q'ʜME�!K�Pk&��X8�����?��*1B.)�i�BZV�[7�
2^�x���̦Q�B@=��#JS���@�6o�|Ts�eC�+S!򄀌	�j%�WJ�)���A�o�!�d_�cS�W�ǲ��A�8�1��1�I�~.09�4�?����	�b�������|��4f�Ig���%.͈b�����Of�� �O�b��g~,�o�H0�0�B�������#��I{K�#<�*���)I��y��D�@["S�-�l����;����':�V��'���D�J�+��l�!�7
�2���)Vp�J�k�9aaxb� ғ9�!:��E���8#�+M&�1���il�'TX�,O��*��'�r�'L�w��@�ѳ}Պ��B䖱x;�A@b�^�N_����I%%.�0#@g�(|�e�gA	d�.���p&��p<9T 6[
��s�U�KvHp�ψ�P��'q@p1�S�g���<b�],t�1�և��'�C�I6"���O/?p�����-(��O���"|B� ҃.��b,-.m�@� ș�B�(_���'?�'X������|�*D�v��;'K�G}��;@�'҄6͐�ia2���NB��0=a��ڗ({Μ�"O�&c����B�7\p6�B�c_�, ����0=�R!��bT��F�%��T��$O=�l�I��M3��iQ�Q����I��},��D��'O	+�D��&.D�|Q6����,�)�5$߰(�)'扏��$�<�`����'B����w�^��1L�=��Y��a�C�'�����B�'�	]+�n�"��=Z���N9���
<L,�/�<B|���I�KD8H0��Ҡ����'
��j�!�j�ȸ�'�D�
���sت1�ɐ�ē�"�j����1��%w�~��ȓ r�ݡ���9|W�1��ɥ9-vh����V��>k�v�)�l�4$��b����'��9X,q��d�O��'!�Ph@�P$p�T���t&��J9]�(�i��?�GF�!� �k܆of�|�-�������Y���l��-��>�6
�z��U�Dᆩj�������(D��]���� 
(▁U�T�~�'A<���<���dqӢ�"�S�&�1��hО,������!��b�,��_x�\�3gQ&)d�d!ު	n�	��)O�FzR�� h��w��m�Z�r�-T�3z7��O����O�ђEfE4�x���O,�D�O.��Z�|p�t�D��+k��X�	f;�c��!�-8<O�0)ų_��[3k�-t�eb��$ޡU��y�h�{��E֭M��m lK2��O�} V����� ��a`ԭC�l�(�)uN�_tP�ȓ6/���;�=�Oڥ(]�]�'�N"=E�D�
Tf)�W�$D6�1W A��| �N8x���'Vb�'^d������|2�=�М��º�4��G��1��p�ǂ/|�˳fB
/>�������7*�3@���n���͜�(�I���N"t�]J�-�$m�Bg3�8�LXB�hå�|��.�X��eO���	��i�&R�r80q�W�j����̎w�<���"'8@5�3+��
ƢKq̓LԱO2\X��S��)����c�:a�v0�FC�i�|�YA�����	�_���ߟ�ϧB��P�� Z��mP��W��M���6��p֨�PX0�&WZ8�d��DU�i���`@,�j ����� � ���b���7�P~b0��fú��Of���'�O�A���T�h�(
t��'K݈�B0"O,��c@[�J����(;j���O�m�s��I�Қs�&���h�,U|�c�t2����M���?�*�^��p-�O���׃ =z`AW��� န�'-�OH��E�D "y
#ˆ�G���ԁ]�k��x�OA�>ոa��JD��dܬ^,��'V��2�Σj��P��!��>e�����U���'q�fd�2�מ:8$�J3��>}����OtLR5�'~
7͌�A�IX��a��H�@�Lܶ�J�Kݶ#���<Y����<qRd��\/ P�(ʫur��+F%\[����$�q���qS.�'t���j5�K9!"�l��������Ad�4v�b�I�����X��?k8���pm�k8��f`Kf��\��%p~"h��,������L>a��y�:�D��>(�0��h�:��O��hO�����-�H�gB�tdMX�B�`���P������d�����?�����-ȃ�O��Qg�&"��x�'<2��Eݿ!��M�X,A��]A�O�8Dz�Z>�'�J`�`S*h�(�*��U�;㾡��'��=�bj��8��z4�P�'�4��m�2)fG ����'�:�[�OSr�:��,�,�!�'t����BEd��7(ϡY{��	�'�����2zP+$��Ml���	�'�< ���Hk��=S��	�'K��)a�(r��� ��]�'O ���'��FKVd���aA��!����'���k�^�9x�
1��	�n4a�'UR9Ӂ� 	*�ʩȱM��61�x�'�8]�˓,����g�(�"��'�]YB�qV�6 �.Oߞ�
�'I8�2�A�e�|�v����Y��'<,U�s�$�B�BrH�W��̈́�i"͢�,A�w�`�
$_�F����V�{�*��oE��#o��5�|I�ȓM�.�Ht����H��	�Pb̈�ȓM�da�E�
2jJ0�Ǜ{ �� �Z�2��F=ܐQ�c�[��,�ȓM��m�K�n�0�xL̈́�c����W�P#a������#n��E��z�����fQ$K�T��☟{��,�ȓr/pi8��X/6�M;6oR5
"^Ԇ�aG"uB6�?q��:�L� ��(�ȓSl>�Zp͍v����(�
��Dlq�H�!+���$+(&`f]�ȓ_7"P[��W�p�h�A�N�N�:��z������o��.;�%8���](<�O�H~`��! �,7dJy���\d���<A�����O�ջ�GJ�=@w�G�) ���'��q�@�X�*w:d:čK�*���уg}�u�v�S�s�����O�d�.	����Rp����C�4w�I9I,�m��L:�&�� ��S�t���oZ�L��]J����ul��s� �$'�nB�I�G:$ͱU�T)�N�
4.V?g��$Z����P���a���~�#��u���O'z���L�Pc��H%b�j5��'�j�ZFc�7FLܠ���=Xra�����.<�i1���/^�����-�_�Y��k�6w�Lݠ�����':��q��KR�( �J�Ko p�Ó0(�}ІOQ�:]x��]A�9��@, ?�[�ω5 qj�*��,��� �+J�Qq��e��HQ%��g��H"���:-���0c6?ILAe�JUK�i�i*$������T��V�u���&B�+��i�%5���s�9TbԔ�ȓ�D�'@�_.`�s���)��F�N���
FgU�����p�<�4/Q�|rR�8Oλ?ih�7@�5D`���eݳZ	�p��HT/<�BP����)Un<�����E��$�lDn�P����0h[�'	_ BQ���7�	0)��j���(�Zy��D5i�*���G6�F�J�d�HYP	�T��Bck$|�m�ŉ	p�`ȐA�t6�@�ďȆ[��0A��'Ҕ�ROՃ�XA@Q��J�^-��O�����Z�]@�X�E��4��x��>�O���s�iԣ`��c�ϥo�t��'
,5:'�ؿyX�0 �AL���:��B�3b�����U.��)�I��fh�	q:�� ���4,�y���v�:> ��O���0�Ņ.�����Zq�i	���%D���T�0V�Ɋ�E[ N$, ���R7�ў���>\�B��@�ܙ3��a�$O����&
eΝ�t�+@��ъ�
�PZ%�BAȒ�L��5�.L`P
�E�k����?.�!3��9:�^,c&���3�J�Z�DF>�:�����$F����M�S��%�bMHl��T�'��P�!򄙍f��T��(j @T�W'R�5��j�G^*RУ
�O"�Y��3?a�ɛ8��|�'�ȏ���8APa8�H�i��b�R ��$�p���U��H(u�C�(D3 kʙ1������3��RC0����E�Vq���/)
�C� �$|�,�W.?)��F���[D�<���!M�^�'����v�����I���GC"-�"
*G8y�#�'F�� �?TR��T��-�p{fl^�HR^�A!폨���+�\��ݙ^74q��/(>v��C���0C�C�ɹ�4|@�AA G���pf� ��p�#��'4��̓A��O8�����s;H�q��|"��X	�HA4&�	7�*t`�%�}��HN�q�N�+S��o)����an�X0�%xB;��Ϙ��h�. �]� gP� V�7(�8���	���`�E�U)��6L�}ۢ�R+R�3�e��qz�D!G�Κ�̼*��ē����G��!e�ծk��(���N�d�b�u����`�;{���1�dܦc.P�Z�'�!�f���A�;S��l8���d>�B2�\�p�$�=~Ȁp��#��@�O+�	2�,QY�(ɲ&����"ߧM�D�Cd���-iƤ�`��|��B6,�}n�B�}R
ۀT�҉S�ޯlT��䃂X�ȒFT�"w~�b�J�%���_u$Ks�̝=u�\ɆjSiZ.H�U/Q�t����Wo޵,(6�g�'���d���q0�$�h1ŝ�H�Ɍ�x$+G�	.��`
�z�L<�'+�#F���L��o04�@r��0:28pd����>9��k��⇴}d�`lL�s��b��Q�~I;�OƌAF�c�H�禵λe�69�U P/�> ��	jd*M���%'68"f��&q��=�A�^�b�����$"jl�σY$�� G�&�O��*B#8��mQ)M(���tϜ!�XMpˑ� X�ЀJ

ẅ���$w1�	��ا�I��Q+B@P��Gr��M��c-�6bU(HJ���@f�I�rm���$��2�ɽI�&�q�Fѵ(�.M�Ȑ2`���dB<7���S50�O�=f��_رs��(?��1�c�ɓ!�J���gX���{*�@�a�v�U0�k�9_.v��_67c2(�6C�<��CH��?ɤ��,����i�@t���I;D�(*�g�+��c�(�o�kL��@o@�,��IP��O�9O���VE��� �fI(l ĉ�h.��Oʧ�M�� �#v����'l�,	���S��Q��H�_֮e��(ڲ`�Zl�4�M<.���<���L>&����[(����GH����Cl�#{d`Zʉv�;�daX�K��E;%�@��r�U2������o���*8��k�5�Q*��%�HeaSL1�'}���]0��l"csr�c��=v��Y0��d#�r�ʧ>��q�w��Z�� 7A�&Pxe�68����!ePSDh��yrkA2���ɲDclވ?	�p�΍_�=�<q�ޭ><JЉ�&@����J`̓@LN�z6�зMf wc\���HD��c[]��fPv?��$�\��n@#6����5A���^��Cŉ nS�*rB�:7�՚���zԜ	�2�Q�b��ͣw�NM̓f������O�My����͘�&|���(L�^����Ś�0'���͊,H31i�/>l ¥ꁄ-�I,�`�y�������hΌ_Ĕc���shώ[̄�b	ǟCa
"|겦PR(J�Rb�_�N�T#Ӧەn�
T#���eF��I��:�|�B�]��ywϞ�Kq���#�Z2j��|����oj�z�'������Y��js�J��P��W�P�Kt���d̓�t���
�vG����՛<���<Y��؅ xb �1'\�	tر3����!}I#�<;R��y�	�|�R��ƏC+�6���7@Dᢱ�՘'������.4I�xyLZZ�{�A�L����<94E�h�\����S�T��Q@�1a@n��& �O��[S�8#�K�[���(���`��K��e� ��\ ;h`TH'c)�I2 �t	�g �+�)8��:�'2>}����,�l���hG��IR%��'.18��v�F�_v�ʧ�.��w�( ���A	9z&�A���5���Ŋ?Ԉ��!cK�yң����剭l7DɊ��'L���B�D�D>���<�F�T�����rK��(� |� !@_�c~ڸV�7H͒�Ȳ!Wk�
)r\��!jQ�rK��D�+/����E�#��8,�̰�0�L!4SD0q�G/�&|�%��N��@7M�Q~���d2�	�uOD`ە~:l����݅��%���_�j�^�ȷ�I���%��`�g�*"�ջ���z��IT�$��D��$�Sb�I�&�A��b�hꤦe�Px��+D�E�#|:R+F�����:���U�\9e�ՈUnP�hE�B���=�OE��W>�p@�&Ƅ:r�1 �F�!/^9���p%�l�'HZ�䔱+0>˓v��HB�A28�P\��CG�Lp�1 �y�KW��0&��dd%���%�?��<�`�
&1�e�`ڈy���
��O.�A`�c^�����M��X����D��	˪=_����?ը�g5%�T=p&#��H�&i��B�Z��PQ�@�#'�2���e�O.�3��?� �ɂ�m��7oδ�1@����i�,�t��OɃ�Hң|t>��ٟε��{���4P@�7/,I�\��P�;�?I�	4����I�W'"�,�"�aQ�$|R<!�Z�d|����!�<V�i�D/�Q2�b��	�O	��s2?�r@�c �L%m`�&��
�>I��D2�?q0)�pr�ڐ���?�3'��<涉��(R^��!D��)�HON(��G>�hO�!t��
g��%�GhG#?�< +�� w^�r2�N�9v5�w��6��H���)r�;>�x��G��&(�'�æ1bC˗>/���2vɔ#%p$�q�$6�_������20���7-�+y��Pm��T> XNb��!!>�IV���ɧ �7#*y�0B�89Q��b�A���<�4J�y���yj(Rr%���K��iĶ�e����sd��ᑞ�iS�l%Gݠ	4��s�56v��VA���GyD�I���	�N;ʓ� ��6����ts�B(�6��d&2��E��e�1J�ND����Dl�'��\���$45v�fg͜3�jEA ��9Ξ�I{k��Ӻ��'t�v��s�$Ԉ���	gKۍ��t�#��5qȺ͚GhL�06�ܪ�_7y]��ˌ9�'��	�o�rW��!7ZV��7N�֢��2c~I�ai�	>c$Yϓ2����g�t���E��MB̻chY�4�B�I#b�h�IVy2tyb`I�tM�*������1`h:!�J�7�\@�O�&�G� ړC��X��.�+�.�ۆnF=7n��&
H�6���gFFy$�zy�oV�-hQ>eچfVHH��sF�����F@'6�Dx�̖�A
�b�I~ZP��������-q��Iԥ��B�ө):.��͎y?9J�<��.��%�V@��?��Ѐ�L���Y8:�ː�,.79
����Q��ᛁ�C�Ly,��v끃��8��	Ur\��U$(pN��Z㤎dG\���1��Y=eH���B�+8�e�҇˥29�PpB�e�hS�	��](��<<O
�(Ө�>�[�q�x�ksc�y������!0�T3���v��p����M>|�
�;L����Ff'?2��ь�7*�n�Gy��?Ȉ�pȳՠ/4���%�͇>ߐ�ۢǞ�HO,�kԎ�hf���S�/H�l�gW��3��ch���l	3���v4K��Fx�O����Q��2l�f����?QᆁCW�]�>j(�S'�Ӣ5��t��N��꧎Ru:,Xw�_78��eAS�����?��JX�(�.���+M&�Pw%�z?y���*1!�
�k��Pr!�L�n`�?(�vmVK%bL+���*2��5q" j�n��ƵD}�	Z������8ɸ��ۧp-�4�D��%	wn��Ԇ��[�|ӊ:�&(ظ �~��R��^m6�;פ���B��<�p��F�T�M�O��zC��* )�c��1^#�"<9�c���p��Z�~:APf�PٟXkq�{-���� q���M�>֖��Wb�<|��<$F�#;#�({��ʲS~J��h��-�X��C��=i�j�A���8�ւՊ�ܑ���9T]�A���i%H������uO�ls�Ě$}�� �W����}�AJh�	�G|�|�EZgͬHг��8eh���#�	h0�!�(Պ|�h�s�ŏy���R6�B�������)�'c����m�7H*��@����p���\���U�h"v���Xt��%܁�G�3)�IFZ"6!��" ��@dR��DD��"8��Q>bhء�Z;W��+��:��p�$�3�|�ҴK�6.�:S��a��V.I��@��_6�`�O�H��� pA�t�'?���|b��9A6�ň���8H� ��(`1�)I4Iy��4��{JP��&h6C�E���\ � ���u�-��B�,�������D�;��lz৖#A:��r�Ȑ��It��!�J�!�F�|��>�HQ�=J'S�U*�e��)U�Q ���ͣx"5!�N�?RD�Ol�����*U2��π�I#ҝHa�,��IY��Y)�aZc�*��&�.9J�e��Q���F����萧�H�]>t�8O�O;q���1'��eݞ���R�.�^���"O�h[%&��y���A�O�=?���6O��"9x$��O�"~
����р[U �C��G�N��̇ȓi�4��2�VG5l(�tB��$:a�Oj�R@� s�H���.q�z$a��d��l�����!��]}Ԍ��;ւ�µ��G�!���	!D�ȃ���Y#p̻�*}E!�DOK v}��FڥS�R*w#I�P!�d�b��E� AV�����@;+!�Dփ'�$Zv�%��Z�(S6 !�dP�>"�|�%��c��񀩟9G!��\�^��5*U��'��D���*e�!��L�t��p��Sb�LX�b,є&�!�Dƹ�|Mk��I�JBQ^0Vy�)�ȓ`Uz�10�A�`1�,z5j,�bх�[b(���N�F&xɂ���J.jŅȓ_!ܤ�@j�R��q�E�Bx�H��c�h-�Vo��XT0v3d6���S�? l�Y"w��ѣ�Z08|��"OhA#s��|�>iBe��Y��@:�"OB�#(�'R�:|�C$��1��4�T"OMV��-j}����ژ{T"O"�cË4'����!c��yՒT��"O\Mɖ��'[,0��,AY���!"O�Y�d��-4��䱳,�>7~|��"Op��GɟP�px��9a:La5"O0H�tʇ}�Q�g�?6�EA"OZHZ��(h�@�J@.v�)2"O�}q�ȕ�pֶ3��"8*j�"O8-�W-�@Wl�14P#o6�K3"OV� ��:`&�izt�ۘk�4z�"Od9"B//Z�!�W�O���"O�L��l!欹R�D�"��"OX̊����p��
Nk`���"OJ�9O^	��x�n��6rX�&"O�`��(3WH���ͅ?X�t;"O�CQ�E�F�"A���@�oR�H2"OFm醯���i�"˓�虋�"O�Ub�Ŕa��X�K�u�m8%"O0��];��f�4F,��iF"O�x���)�r)1A��esp�7"O4U��>x3������h��+�"O�����>�Ѓe�YRpeY�"O���2�K1$F.�8*��Ը�"O�}����/42���O6����"O��)�EX�	o*�p�&I�v)�"O�-�㯁B�~��Z.!��1"O�XP��D���Y�A҆z����"O�`���y��8�4'L:��Q�7"O��x�JL��8WG�5nLm��yrDQ`9��ֿ>� {d_:�yREX~,��ca��)ֲТ�c܂�y��$���b#癨ln�e�䉹�y"M�Z��q��˞^$uy��K��y��b��1�tWFt=s�/_�y�E��Jc�.L%��mu�Э/��B��<4p5´-��
�j51Wț�$��C��-L��zvK�.�4��,Ykf�C�I5t��уE�҉�$��C$#9	�C�I�J��15��/u8u����A��B�I<�z�kPd�|�N�s��GN�C�	"N�V�Af��=-<�:� ʙ9��B�ɂ�p9hu�� ?�\Q���Ɂ}m�B�I�t�(	r0�V�kW��w�H�}NtB�ɪ_�-��%��L�)VXB�~�Vh@����`�9Q�LB��\��0�$�4�"��� ݼ"tDB��3�TH�s�"B����!��\E|B�	�u�����������;v�
B�	�S�������䬻�"P"SB�	�q�1��Í^cx��,�+��C�	���MZD �Bf��"'�u�B�I,c�!�D��
�1k���p�PB�	*�0��Cdݮp"$��p��w��IJ����H��jƖ�P����=��]x%"O8�Q���$6u�\z�mF�(�2L0�"On$K��n˔��LY�)U��"�S�I��RB:� s��7�je���C�!�	HAp����	�t�� a�-�1-ɚE{���'��!#Ոkf4�;R݀�P
�'z��
VH�^1�XSC"#j�`
�'и�q1�Q�{������P�	ۓvt�0AJ�� �Aw�B8~@��df��4�	�"O�)H�舗x��|sw��T��D�0"O�H�g�X� ��H0��t
�Ӣ"O�\�������JJpS�s5"O~5R�虠. Ѐ��@"9=r<��"O��p�Y$
o��vcc��d�G"OP�7�*Ru�Dx5a��w�P���"O��R)	�}�F�aℤjH\t��"OZ����7�*�Jcg�B�tP#"O��Aa�)Os،�Ѧ�Lh4I$"Oԩ(TH�$��y���)P
�z2"O��ˇ��6ʹ��L� 
"Ot����9*�5��iJ g`���"O
43���3�b�X������p�"O8���+i�p(� �R����"Oh�rV��$�Ѣ�����$��"O���w��1>>D�R��HzQ�*�"O�ʐJ�n�`	bu�6eI�,:�U�h��ɔ>��dk�C _�F4QFJ�>@W�B�"*8���
R��:���� _�B䉓,�
Y�o�+\�H�%h�b+L㞘G{J~b���"D<YsA݈g7T�2#g�<a�&8㞅	!�V�HJx42"�Vb�<�� ^�����8P� VDb�<���Z|@��ˋ%����WE�<qAB ��zu"�d�	;����֎�D�<�R�/�����S�"|v0H�M^J�<	E {�|Hcd�P��iJ��[��hO�ON��˗��9T�T��JN��-p	�'}����kY6(A90uE���:���'"�pC�T��iӴ�>T�@l+	�'�1�4	[�,��4���߫;�) 	�'w��B��D�T���7J�ҭ	���\ (A��TT�hx��C��a�ȓZDu��I�/D)��C���p5���ȓq�K}���G�O�`��'fazr��DH�ɔG�`�#vAۧL5��p�9D��f&ŷja�����'8͖Mjs�1D�\K�
ǎ'��N�0s-���'f.D�h�QL,Z�>u���M�I\p�jT-?Q��:�'(f�%I��TZ��Fƕ�,����O<�o�s��`��a������ON���' �'đ�[G�K#���a�D8=�C�*.4���,@�d�bi��|���ˁa�<�'C�.�*A��H�k��:� �^�'L��'U�O}�J��ˉ\�����*h��'a��]�Э �J(
��`��!��O�#�u� %Quq3�Ë�X?�U���N@�<��
��~��ު^��"NVyr�)�'q=$�1�MH�ynh�R� %d�V5�ȓ\Sp�F�٢'��T�r=$���Ɂ'��D2V�-�L)�HRK�R���$��l?����x�u��OD!Xe0M�Gd�~y"S���<E�$�>wm�qD�5J��!L��y"J��-�L�Pvh��~Q���7C��y2)��p��U��Эgi��Mˎ��sӜ���ȳz`�k�0@?D�A�"O.I@�Z/%&����j��l.�˧"Ol�s��	My M�U(^ q�^��#"O�/$���@Ɗ]�l�w�P����'���'���gh_!!��@�bǞ�@tX\��'I��#+.�a�a�S
�\�����y�/�#i��Qy�D	n��Y��Z��>AK�,`��ד
��=IqΚ�b�nQ3��o:� V�����-�F���L��O��0�3"O�=�6*�
j�ag�����!6"O��;�lH������ ;p�<4Z��!�}�����Γ�b��A�릸��	g~R�tL�r�*<!Ǥ���,�+�y��$T�jD��B����w�ϣ�hO����փA�� Z�'�!����G=�!���~Z�+ԇ��:̘}�"$�@�!��i���)u
�R[�X�a��P�!��ڇJW���B	�P/@%����Z�!�T�h�Eb�">)D��V�ˑ!���%�N��J�:,�u &� +}!��[�4��A�B t�0�k�eA!��	}8jq��9t��,�' �4�!�d�(�>a�5�z �/��j�!�;8�D��va�
R8�qsn+|}!��6O�
E����4�j��]�e�!�!:�|5x�F�1v�,�5O�`�!�$ށ_
�*�)�"М��g	�!�D=v��
w&�����Q��]�!���/-'0�s ��G`���$1 �!�]�,�n0{�a�vl�TۇaD�!�!��ɓX��)�7�η/�
J&�)ϑ�G�do�8�����h�Z�xi�2k���yB��?;�0����J�S�AB���y��!������Lp6 rD^��yB �&,��(��E?���$͂��HON��T�'xf��LZF�Ny���)E��]x�'<ܕ��+N X��9C��>�*Db۴�MS��)ڧ(�&�(��DL��1f� ��M{�f	������<0��FH�<��&���^��Ȉ�%��e���C����V��Uz��x����" �7|���{"��� QMB��t`A�Sc ��ȓ*�P���ͳ0k��r���'hZ�ȓ90 �Ȑ�� 8^9��X4j������?ѧ�V 3na!{�2i��
����'�΍�ʂ7�<՘��=��p�
�'�vT��
@�'�0��3�ǀ,*h���'a�E�u�3V�p�k�4T	i�'�,���!��q+f���$��'!N�@�'�Ȱ��&e����O��m���'z�R���8r�[��M6e�FH�}��'}���+AN�2m�P�O_׌���'�������"iw�U���/T�Ԇʓ%��X���U�zA��@��(�ȓ-l���M�z������E�ȓ+�8�B����|��f�0[��L�ȓ-,v�#ˉ�7FL�;��	�hs �ȓj�*j	0����!	�!� �ȓ)+~|����a�ر�Q�N�T|����vP����3� �
�N�8��ȓ6�<j��ŠN|(
@IR&� ��璉�K"�����؅ee�ȓi�y� T�6,h�y�G�e�`d��2'~�2�,ްF����i�#��^[�<�.��h@e-�"/��ez��N�<��J�s�"�p[�oN�	��I�<�"��>m=�L�,��1xF�F�<nT�%�F8�ɮ����4���<��D4r��ɀBIH��-(u��v�<aaKΕ"�Ɛ�3�fIErc�|�<!ѩ�RK��8�-��p��\!W/|�<i��$P�(�Y�+��H�
�;� �c�<� N��C�H
���e D�5�J@�r"O���T�G�8�����Oűl�>D 0"O�T��O;m���*���$W,�pP�"O�t!@�d��S�hO�J���"O ��I��I�01d*�p����"Oi'EY�`�T� �(�O��z"O���0��(a�lӧ5�$��"O�`��8?�FxQA)L?'�
a7"O*�;����JD� �����"O���V�8*줘��ą�Sd=��"O�̫�球h�FD
Ra��X陷"O��h�l�B�l����X3h$�y�"O��rc�:H��oѴ>�`}��"OpD@��1�<�î_�Q�8��"O�eI��a��Ųo�^h�IK�"O�(+�aJ-C� ��ډUH��z"Ob�zWGW�2�4	�.C�,��1��"O��:��CRT�¥�R���jb"O�� 7OZ{6n���jաR}���"OfX�iQ��Q#
TmC�d�D"O"x�1�N�0�H��p-2��A"OH���N͟$��%*7��,o-`��"O�|4N�� ��)�/!"�×"O�(�Ř$mp�Ua�e�]3"O*�j��^�Ng"(9��.\��	��"O�����/�bdÆ5}UH�iq"O�Y؃�P�sJ�;3C�;X�@�"O�H�&�L�:�H�Bi6����"O�=����D)�� #k/��	1"OF}pd/�i��8+��:xzd��"O����>�đZ���&o��H"O���9JUY3扡nh��X�"O����
^%�<y�䆱g��
�"O�8[���(��#\$If<x5"OL�)��T7"dhT�2k�FZ���"O�}8�.(nI���SL�
dB�L""O��3 �V�t,I^r.y�am߄�y�/G�j�i��7*��l(эR�y�f#kBtp�C�L�� I���yb�C*&!���әO`Hcw����y"��7����k�I���X����yb���c;�q�@��T�x䠃�D�y"!:}~�ث�FY�L�dh���@�y�%K.F�ȘۂD�H�VZ�b��yBn��4:d��<�,T�����y��C/�����6���땥ך�y�䁫 '���U#�;6a A���C��y���8/<8�9��R 1�&%3�Ւ�y�gE�Ț��#̗:  ��𤒬�y"��b8��y�g�"5G"�h� ��y��G0cV�J�ƜC�nɈ0A�yr�	��I�J+S����N�y��>1rP+&�үta�%ʗĘ�yr��dQ|�⫘%Z�VYʆ��yB�'Q3t���z] (JE��y2��=j��#�Z�Fc>��$@�!�yRHe;'"P錜?{J��AN8�y�L�D�Y�F@�9;��`D���y�� �%{h�����;B�|)DC��y2�T5+pٓ%%�2b����ˬ�yr	���-
B��4*���#I�#�yb�c�r�y��M��<�����y�O��v�2a�䠁����#��ճ�y��U%Z�Z�Ó
}j���+9�y
� �@����x$��\<6��\#u"Ob�J�� ��y��Ӳr[估v"O~@��ϩ'X�]ᣮ�</HZM��"O�8��m�|t���eWl��"O:A�C]	S��]�U���ڪ��"O��U��?M(H�r�v|�B"OjY�kP�@��f��^���3�"O��C�1<.����o�.7�x0Ƀ"O���a�#0�D���""t�*�"O6us ��U���гM҉��"O6��F���e�PP��:bʔ;"O`ZP%+dfȡ�7
�>s� ��g"O@irFJ�,\ڨ��h�=��,;�"Oʙ�ⅰeP�gA�x���2"Oy
���L�9Q(�@�B���"OR��b��T~�@Ȁ �Wy�y�"O<Q�!�ɓ ̤� ����t�]Y�"O�@�2G�P����GlD�07"O�]�e�	Q5��@�/�!]e&�˂"OԩEk��m�P���㝌W��zR"O��aE��8<l ��`ϚT5"���"O~X��+Z�F���P�%��d4�"O�q�
שXSf�bE��r!��6"O�Ek�����3c_�C��%(C"O�T�B+���x0��<+6e{�"O��ch^����.چ &�0��"O��s�]�e�Th���<@�"O��qR,����qH�n��`*�"O&,2�+ʾ=�Z��tN�'�0�Y"Ob���.Nc��DAE@�"��x�"O�1XpÂ� ~M2�Ԩ��""O�ԙUk�C�ǯ�D�\e p"O�����y����.\�{�X� q"O -ag���Q� F��O����"O��K �T�Qr��`�K�U⤐I@"O�ɱRT x �0�d��<�L�K�"OV,�F�U�Q�Z�3�,_.���s"O�+)N�#c�-A�,��H�1�"O��bU�:��U�0y�Xa�"O8���Ow0)s�d�v��r�"O�A��&
e������1�N\�c"O:�x�/)�FoN>��c*Ob� 	�qZ�XP��7����'쒗�Hm;�8ibb͹R"Oj)sb�B&`��h@e�"U���kq"O @��,�"��S���x���S"O�� ҃�6I!�X�"DQ�ymT�R�"O��dL�v�d`�� PT��"O0SEjѧV�fd0���O� ��"O8��mS�R߸* ] W�>��"Oz<b���1o�bPC�	�O�V"v"Or,�B��v~v0���J$r|H��"O\�1 Z�"�.MU��CzZU+�"O��R'�.%�y��K�^^x��"O<y�3oJ\����"AvP�"O��0�cl\!�%�C*q��c"Ol�Q�cڹ}X]R��S�elfL�"O\�Zr/UUD�ȱ�!S/i`�QJ"O����+k�le��ʔ�A참�"O��*��r�T|��Ɛ.Κu��"O�q�ίdp�2�w�f���"O����S5lj��9Q ��Gf����"O
�9u
*|�0h�$�~r�c"O� Tn�=c_��T
A�+>ȹj�"O� �,��Oф{\�| c�\C0�qZ�"O�
P�җY���p�Ì�;)B̈�"O�䩖
 �<�y��#y��"O�%����K��3cC�X(�:�"O����aζE�X�p����9+ "O�1�L6�t��1A�;wZx��`"O0q�RJ� ��	0sO�uDd�kP"Oh�if��,Uib�2�?�mP�"O���HG	A�ȡ[��W�Xx؊"O&$��7m��#F�,g�vAY"O��8h Sl�xk�BA$6Įc"O��ѠI.�bԚ%!��
��e{�"OR-��֛ B:Ȑd�M�,P۱"O�LYJ�3$z�rG�ުB�
$�a"O�H���HOvN�8��
9H��÷"Ol��M9k4^-�n�Ԝ��f"OHQ�A�ʼf�"���Y�"��"ODd'�O0/���$�|�M�E"O����A�9p��S/_�_��K�"Ot�����o�d�Ӂ��/~8tA0"O
����qPTE�0��(`��4"O`Kcd !�*I�@nS"R���"O�PAkЩuVlH��]�_�v�H�"Oh@��K@��1��,@�a�B)��"OʐB]S����j�% ���`"O�9�m@a �)
4�	�MǎA`6"O.գP^� j�����f"OV%H'�@�E�0�C��ΦT�&�1"OU�s��JЉB��\/�f���"O��22�6A�:��T�bk�	B�"O����˟"�F�Yd�Z��l0k�"OX��B��+qֹ�T��� z�1�"Oz��pė%1��1�V��B�"O�y�C)�'Qƙ��LZ:C��a�e"O\�n�-}22�0F��n�;�"O�i�&�k[0q�KG�4$�'�d�e�
i���B%Jۨ]����'jNI�cW�(�0ŊCU�UN���'@�� �S���2U�Klh��'��S4�ոR��@#o�=0�Ls
�'
l�A���/��kGm[!6�q��'�x2�e��%���E�P��a��'/`#2�D�+�d<Ѕ���Z�I �'!�A�AR ���o����I�'��K�<q�e� ��*�'��Qpq�P�v�,a��P�l����')>�Hģ�J
���Y�fT�h�'�P�j�
^��p|��I^�W0�r�'������pĄ���UԐ�i�'�"U����\c���.��ct,���'��ڀ�	�h���/�����䓫?i��L�� &�ڏ~��1�h�IT�m��7D��B2�X*A�1��� (B|:5l(D����aJ�v/\�<�d���UM�<1�	U�����(26�(���NK�<i�q�NIQ��9*���oO�<	Q��,�� ��8G�2�"ON�<�Q���U��{E!�.d!�%��\�'axr�C,�Ja��/�|Ћ(���y'�n��A!�"��=��%��yjˬ=��x�%N-�(�����y�C�O��s&��xP���8�y��-�8�{ �ܺ�J��E'�y�Ȱ'J`2����=ɐ�K��y
� �a�s K��F	0�؋6	,�O@`�t�,���X���;Ҳ`��l�Oj���O�����$G@�i!�AF^�9�b�ڡ|j!���;��yr6��g[��2wf�$}f!�źC�RDR�,��WL\,�����;�!�[E�T]��Kצl��qG�]��!�d�<	��I�A>-��!3W�A<�!�d58Т��G(b{��ᆇ_�
+��'.�[P�2� ����b�+��'�!�d�%^1ҘA�a/oH�v%�l9!�D^!qɎ�C�#zK�-���E�;2!򄝝����G%K�wF��{�n�8!��	7&P�B�܅T2ZV ގL�!���;
��
S%¿4&p�D�O�!��z�d�Z��J�)�V�2#EÔ��B�'�F�􈀟1��pT����L
g�'�O.�}��2k���N�}]�ykFm_=zxȓ�D��9f���zƃж>��-��8���2g-
 N�N�rdӳe�5�ȓm� 1 F�(����a
�cc�5��g�-�7��Z���SEJ�L��ȓK�P�{�iI�M�����!p}��lV�ࢅ)�VEkr"C&~%�h�I`�����?W`��y�d=]bE�o��V�B�	�v��Y�ƫ8�6�J�E�4zR�B�	�r	�4(dB>d\*''�  �B�I�;��$�pC�'�̡�	�T�B��	4�bAUhR\�yag	H�Z�B�	a$\t�A�	�U��Qq��V�B�I}t����'w<��q �>Wu�B�I&k��a���.m�h���B��B����ʯ7"2�Q�L�1VHC�)pn��
֋A!���0�F�"C�	7�u�'%��"�H��t�P��.C�Ʉ�xݨ�@ i>A�SGC���-Yज�}}�fХ)�BC�I'˦�?X��
uED�	~�L1q"O8]XA��h�LD;ƃ��qkTE�U"OT5�goSF$�$EW��i�s"O*u��|�L����;}�����"Oz툵(��"q�)'	M����"O�F�p��IJ!n��t�ƨ�a"O�(p��9u�h@��5�F��"O*�R%�б5ȠP��d@"*���q�"O^����ʰ��f��U���"OZ��!��/���!�u����"O"	�QG֜%�n5�V���KoR$��"O�p3"!��t��0�  8����"O���b�Z�4�Va!�*,,:���"O������1��ѡ�	��@��d���D"ړ��$R�j�P�����+y�UQө��0u!�$6(��L���3��+��/�!����{fKN?�^`���P��!�[;Cz��8��K�v��%c�*!�ĝ42�����@ �~�ʖI�!�d\)C/B��V
�:z>�RAJ�8�!��W��ˆaڌF����1��`��'/ў�>ըT�3v��D��o̱���N1�y�$��
�����)�3#�ڍ�1N��yD�-^���+�/��!��H�[�y���J�(r����f��@Ɋ��y2#�"sZt� D�Jr�`aS��y�m̷M
`s�/M�I���PC��"�y�B��g<(�k�'�M�H�Z1
K?��'�ў�π ������;���1��1}�6"O�YScΔU�^��C
�'����"O��� �D�e��qP�B�4�hi
"O�Dhr �R&G��dzS햝�yB��!#$��^3�\8l�T�y2i^!|3�]��h\;����4��*�y��!+���A��Ic�9"D���y2�լF$�v��n�p�[bG��y���%e~�f̎yd��!���y27��x�`�y��cċ7�y��{:T����u7)S����y�+�@F�x��УrH�*�+���y�L	<
 ����S|B�{��;�y�	����z�KA(rf\XQ���<�y�g��^kzb�O��[N�r��](�y�g%F�x�B���K�|� ��ȶ�yҩE��D�ȱ%4���BK��y��M�s� �+q�*o��)��P�yr���To��3����s��jM�y"�'p�2x��Xės�J���|��Q�%��>��R���zΊ��ȓa'z�h����qh�
�A�^�l��Io��h��$��4��-����7*mXB ��LE!�D@�
�pQP�ȌL����[!�1q2�E��mO��a�tK:<I!��Z�Z 
 �E�]TJD��H�9�!���>�u�v#�,>�SfI0\n!�@�E���b�M܊�ô΁�vZ!��Ű$Tbm��K[����@�O�j�ўp�ቋCy�w�ҤF>1P��O�&B�Ɋr�ڸk3�����3�aK��C�	2`"DE��뗾xf�U�1�Y�e�B�ɬ���CEU�zx��E��8�C�I���lɂ�I�|	a����cHB� ����	�(|�μ�"��<��C�I|+�)H 蜋J����
�C�	�7��:g�U=Hip�zQ�Ne �B�I���xH��E��K�c��B�	� ���BE�s�����H�l̀B��r�zAZTmȴe�p$��!T(o�C䉉U�� �(H�e�Zx(�����B�I����s��\+>�2A)p �C��/@��򥋱d
$�bO��jQ�B䉋v-�ܛ�/L�T^��+2eضn<~B�	/��1l-b�S�	�0\B�I�g
He�Wd�����s
�*��C�ɾ|���[q��>�|����JJfB��+����-�1nbf�*���U``B�ɚc�"�krc�[xNL@g/W��4B䉈�:�� �8��D+�\�C�ɀSA�a+a��^�\����Ng��B�����eRC�d�z���5��B��6\�b��&�Q�J$���׭P�|B�>x�Mi��W�֑#4�һ=fB�I)q�а���]�Q���*�V��LB�I�?0$MS  C(��U��n	�2\B䉃}5��[��JV4��	��LLC�	(j��b�^�f����b�5�C�I8X��\�Y&�-��ߴ@�B�	�~ܖ���gЩ$2P(��I�D�fB�ɳE���
0,	���z�ϒ,� C䉐'��E*WjIh����#�8$`�B�ɖx�b�i���hR!i�&*�C�ɲt��kΊ&3\��8�AˎG�HB�)� �UڇÈ:y�LD�ѫ�$C�x%"O�f"51�`�ߖc)�ɹ"Obd;d1 􈁏�-3
pA��"OLM+pޘb��
�Ā�a� <�g"O��E��s9�i��⑵���b"O`m�e�E]p��t��e��A5"Oda��T�nV�����#-< {�"O�DPSD�.ԼQ��c$0R�"Of$hH��m P�óg@.�$Y�"OPd9ƇX�^�*m��˅	���p"Ob� ԥ�+3�>}�e�4H��"O��eCBarl����[�U�.$A"O��ã��D�)
F�l���"On��B�C�p�ʗ*F+T���y�"O�U���1D����=KǨ}��"O&4���ӪS
�	��]����"O��ZĊ*{8Ĕ����5]���t"O��yu�-]�hH�5B%tJ&�!"Oh�i�r���X��\�E82,� "O`"Cn
�tˠD��et$��c"Oj5h˹KTh���	Ցr�0���"O`t*�`�<���N���	�"O^�i��S�o��Ӎӎ\�6� "O�KU�5|}Ԕ�u�H6Gd�E�A"OB<k��*�M3��_1,��v"OR�E�T��,@3 �i��i�"O6�jw����"��2(�ޜ��W"O��B���e*����m�$a!�"On4)e�*m�tAԭޘ[Ī|��"Ob�┬2)�$���1\�i�"O�Y!
�9��E]�:�H�"O^�@rㄞZnf!��&�7���"O2�j���9C��ZXHu�Ư�p�!�_e����CG#eh�0(��hA!�>���Ն�G�u#�'Џ>�� (IlX9r��	hgR�г�7�y��D2�d��e��1gH�C	�yl�7 �d�	h>�Jp�$���yrϫe�`X1�ېc��L"�cS��yr/��5���+,%��`7I��y��=.��s��lp-��雾�yr�Qj\�QJS�Ӑ��;�k���y����p=B Ct!�	z�#�j��y��L���	k"Dݮnb�Y9dJ?�yb�W�+.� 	�Ju� �s��y��S3+g�y
�� np %{Rlޢ�y�F��-��hüC��pq�۠�y���lJi�1銨G�P���y┶B�	q�ł��H[!#Y,�y�i^g��q�	҂Y|Z�� ���y"j�$��<�`��A�q٠� *�ybƁ+5T��+D�;�D�뇆��yr ͝c6x}��.L�I�Ă��y".��<��MQS�4
Ea2�H�y
W.{��҂�y�6��T�D0�y�MV��Ҹ�0)�uKv���Ȭ�y"��H>�� �8p .���V/�yR��:��I� �ڡU���:��F��yR��>N$lɲF�/!_����-؏�yr��3]� ��v.�>�b�kuH��yң\0��d�0��r�K5�U�<�G���ܕb� �x������Ec�<�#�4)�V�Q�ϳWd�(f]�<��h�@(�� ӭL4�ɀ�mYm�<� �)��ꏧ���B&A�-e$��H�"Od�+��*�����3s:����"O&����\�}�Z�Jr�'j��)r"OP�i��3t4̑à�>ؖ�A�"O���mE9_�ٺ@� �j�u"O�*�"Q;}=��PփH($���e"O@�a�i�� #��`bǷ{z(+"O�@�!W�t�P�[Ţܨd���P"O4�7�[<@��$��L�o�T���"O�� ��F�*��	&�ͩse��˂"O�d�/���r�P�%l|!�"O���2�:*��J]����"O$͋��H�q�N�`Th��"O�d���#D� cfH CSN`! "O�C��<|����j�[_ ���"O�K'6‡�Ϗ�ٙ�"O��c�䁉[@y�,pG$�1�"O�1��F�m���9f�/Ҙق�"O��`�C�0�"�˖�:�B�0�"O �����iܢ� J��Bİ4��"O��/N'dTP%A�)ĭ/�T=�"O�QRW��L@\T��M�Zx�1@�"ON�q����Ss�D&�x�hlK�"O�!@g�M�i�nyȆe��N�f�k"O����K�@���ɅD�:�؁�e"O|���l�&V$ݱe��@m��"O�-ykD��02��4#�ɑ"O����	�6m~R:`�T�r}0�2"OL!��������EA�����"Op8���_1�d�X$މi9��C�"O��&ˉX����t%�7|p�+v"Onq�5.X46jЃ#ȧ-�VA�"O�I`+�AUL9�F)�6m�\ ��"O�yh$`�Uh�g��&j|be2"Ot��}8= �ړJ��bS"O�DIUI���0�����
� ""O���3���#0�5� ��?5���"O�M�e��5���f�E���U"O�ڇ�4a��؀5�RB<�S�"O�� �U8H��m�$���y$�i`"Ot�B�4H%�A*��R4@�8Ez�"O��A�T2L0���T"O:e���F�J{䔉`$�I�"�"O��S4�-
��8[R#S��V��a"O��*��M��|z��V# ,�`(�"O���G�M7bg�ȑ$ �r2r,�e"O��ӧƓ��8#��Ѿ0��"O`Kad��<�|�i��!`J�i�)&D�SB����Y �G�Ըɤ�6D�HhW���q2Ř��� -E�<XS�1D��q��<ن`�0D "U@\`;�"D�<[E�n�VUH�+��,|�c$!D�|)Vk�B;z�#��ϖ0�j��K?D� +�k�������F�6����;D��s*V�&Y(����Q��4(;�-D�|�,P#F	���e�O�"f\�rt�6D��(1G�1g��y�*O	(.5¦$'D�dÀ U�5X������hP�a$D��҇$H�q�ؐ�V'�2�0�B�(=D�����4A����nP ��u8T� D�H��"M>F���ҐiɴL���ⶩ0D��0�E�;�1�iF=U1�T e,D�0 �	8판� `qq�l��! D�PKCL,R|Zx򰇟?��d�s&2D�� �Tȴ.
2��UŎ�;sO���"O\����1u��f-ɸ~E��9�"O �a�����Sw,8A�0K�"O�th%SS\�*��S^�P�"O���K�!���2��,p���"O
{���2Jj�:C�׿V�F��q"O��1��C|xQ��$Q8��"O<9���ǭW���P7h	 Pr�"O�SԣL�G0m7�39�h���"O~�f�	a���&@�ܓ�"Oz��WR�`X��
��C�6X8
%"O���/L�,�h�!�c��@h�"O"��V:R*.=��V�*ꊤ�e"O̸��F�*����cA��4��"O<x�Ůs��ȥM��7@�ɰW"O�p�_p����A�2&Ƙ��"O2�su��@�)��֫>��1Q"O�Q Cꔷ/�\�ۋ1��$`�"O:���ɖ a �)C��1l��@"O�S�jӧfN��Wd�#N,��""O�ಠ��m���rÈ� sΐCt"OX<h�dV4{>p7��_� �Yf�"D�aF נO�~��KE��u8��!D�4)p��i��]���K��i��?D����G�{#�}c*�%cJvM��?D���Ri'~�±I�9W�Ȱ�=D�tx����[�F����=:78؈'�:D��h�#0NՖ�FZ*���ul7D�\r�#H%�D�q�̮+�ȁC�4D���ㆾIv����L�)#F�2D����JF�^$Đ�7�.P��]!D
5D�p���I	T�<��/�B��!�0D�<���!~@�3�^�4�Hł2D�l2�� @Z�����h�0�/D�XQrl��؀@F*֚�vh*D���D&��u@��%��'�)D�А�����	�K�~d�XBSO&D�t၅�&D�jQhG�ݎ f"D��I(��+[�U`b/F�Fv�h�'�=D�$��f��F�0]u䃼#���Ig<D�a�OG���0���P��|!�M8D�0��� �I��	�c��y�L���7D�\a�Ƚ=����l�;
=+0E D�L)v�āM��A���\�"D�$��bW�8�Q�ժɂO��u��H D�|�W�7V���D�0
��I��!1D��x�̄+"�4����>���N"D�<�ϔ�'P��̍1_��h��>D���dލd&��t��X����,<D������6&+�t���E(|�l���L7D�d+d�3+����4��͈B"0D�0��
I���Ł޺^��2�,D����	Ko�PT�>ts�Hkp�?D���UNۄ-���,(C�<Y��;D���tc��0>���7�ƈ��9�.D�L�T��w�L��i�`Gx�9�-D�0�֤�f����cB�� �!f*D�|�mB�*
�ˁd=E�u���%D�̙��*NϜD#G��%,12�(�#D�� �-K�"ly�M\.l7&T�%-,D�l�1!��Z������Z%7��m�i-D���WJ������Bڂu@b�z�� D��� �]�̶UrE)�g/4�A�:D����B. -R��E���b$�PYb`8D�� ��A%L�.YU�E9�π2�d�q"O���%7:��h���ʸL[a"O�0�$?&��{f<Q���Z�"O�!�n�+�`QW�Y�u�����"O� ʤIW6L���𰃗�<�(���"O�qQc�l�d:���4WJHC�"O�`���Z+kp
�ۧa5N�T3�"O���G��goґ��@O"i�葐�"O
��0c�Z��� W
&`ȡ҇"O�|H��SxԄY$�6
�t3�"O �ѢE�|��m��t<j i�"O�-�Ā�"!@u���H	$JEr6"O�h��g�/IR��(wE�97�� "O��y�)^����D��@�(hU"Ob�{!kܜ�.�J�h�2Wu�m��"O�bROD2̈́ w%"6Z
M�"OzdP�P?��X��&�uT�a�"O<�q��t�Q1Ѕ�VQ���"O�����"�@K��X
O��J�"O� 7�C3Q{�b�PB�kw"O$`3Dȧs�ٺ �O�>H,@0"O�!�Ħ���>��p��Q3N ��"O���d��"o$Zp���ћK�x5"ON�q ��	���K���\ ���"O�A�DoP;shl�A����bF"O����V�g�p͙#��'7ܖ��"O�9���(=2�5`w �̎� "Oh@A�ȁ8|%��r���F�i��"O8�K�"��JA�0�f.2��d�#"O\2�,)�eQD�ۭ0^�,@7D�X97��p� ��C9���w(4D�X���Tm�L�U��#��<)��3D���L�?nTm��$�谧�0D� h�`G2-�(�� �'Ǧp��+D���O&��)�g�4B������*D��S�Imk �wg�8�����f6D�̊/��I�����S�r��`�75D���5�ńN��A�J��1i�e q�3D�T:�Û8�\� ��?�	ˆD3D� �3�Ӭ����l[�oֵ��b0D���I�x���� 
�Y&�5ؓ%/D��q�E�>�ڵ#+�w#�U�	/D�4j���!n�K�#��&�΅��?D��X��U��+�� .�0��n!D� �O�`{�D��ީl���b�a?D�,0&A��s2 m��.�7w�qjf�*D�`s�g\�g�`�Z���8h�e��#&D����U'.hQ�L�x�@��!D�P*R��1���X��Ё{3� �A*D�434��}�H�3�ۢ!�
5hS�+D���7���,|�tAeiZ;<J%���(D�T�4�J=Q �q�WK4` �`�&D�X��r�j�s�χ�Lծ7�ZM�<����l��@�ӌ�1��Y���^�<���]M(�8��JRѬ�꣦W�<�$#�.�Q��a�.l����XV�<���� =�|���p��婇�g�<���C;?~Hzd�� X�혶/D�T`�jԩ^��9Qȇ�y��!�:D�pi��@�9)� �� D�X��m
�8D���c��L_�8�A�­WZ�5��!D�(3��Q&ǧ@�ql<h�a� D��0��X�ec�T���3f�>D�d�Ʃ̢
����� �gq�YC�6D�� j�Hg��`�����sA�};B"OD��%"B���q˰���1)0�!�"O؜�ƋUC�|ݢ�c�s~并"O��P�A�;���v�?o[A�"O}Y��	!�:PgBR3.P0�b"O�`j'�])>�c�@�	Q9~�""O�Ձ�Έ�n>Vа7�Q�5+4̰"O��W��rv@�-{y�b4"O�R,�&`����h� ^Ty�r"O��
�~�"r�M`����"OTA0C#�s��)�ET�v�p�"OV� ˜)A�$�҃R;�@=��"OV��ŭ�V�zAX�̞�2���0�"O��f�;Y�^���DD�����"O4-a§MfA4��&�R~��
�'�f�K��¶s�I���*����	�'��hS�d�V�{��p�'��9��Өsiz0c�<Dv~!�'�8� �ܽ^�h⇅0?���'$�\x�o[#4��+����; j%�
�'��[T���k�D��`
ͩ*�`���'�0`���"qrp�2�*	�X�!�
�'q��t��3w�Q�w_���'[���_�=�J�	�V2i��$X�'��q�f�PH ,A� 
`�VU��'[���Q�%-�r�t�ԃg���)�'�]l��I�����+[��X�'�E��o݉Ql��i$Ï"*-�y��'$8y��l��y�,z#K���H�:	�'����ĭ	�5}��Ys!�7|%��C�'��9aШ�*;L�Q�m�t�
qs
�']�4�G�^�lX�LrS ��:=��'����L�=I�X�q�֮]|Ԝ8	�'�0�E����s�bFQ��m�':8
Dj��[$�%Z�-T�S��Y��'�Na���� �J��B�MpЁ��'��� �'��`�d��A̋;��(�'"0);���"O%�}Y��Q�D۠,"�'Q*+�S![
���;,����'Vl�V��D|��$ݸjV~h1�'����G�L�" �N,,�I�'�TPBt�!u2�y��Z�]��'Gv��Ui�<��2��
:G����'�h-��M�4�ҹK �;^�P�'~L9 ea��L����+l�e�'���C�4LL��X�F%1���'��19f��tw�	jAh��"N�d��'~Π:�C�7׾q��&�j����
�'�$`�v4Ъ�fyЅ�
�'\�8��+��u�`��`D�\�>�0
�'We�G/D�B��wLx�	�'Y�����ĉj<`�p
�yG^T#	�'F�����RL����`聰i(�'��}�&�(h����zlz�'xʁQ$��S%�q�g�V�'�lH��'�j��!�N`���(�E�22F���'R�N�>	�0#�J�v����'(��@Bͷ7��PI�q�ll;�'�T�z�,^:N����0\}l���'��P#q ��F	�չT$ؐO�����'���I�'��H��Y`��9�%A�'���4�I�Q�4�f+O2H��	�'��4��,B�HƩ�Ģ��*O>�@�'1�xs3�Ba��!��-�v����� ���E�3�����@H�B�#�"O��Qi��^M��pB��"���"Of�����b�P�2��Hl�I�"O�(
4�D�J��WF��rx���c"O��B�,M8Snj��$���rlq1"O@x�%�=5��"�b*��%��"O�QD�1Z�\l�֠�j��"O�Yt뙠=���KGe�7.c�8��"O��#d�A�c>��CMiM��j "Ol�h��
x����oL$DV�c�"O���1��4��u�� N*�S@"OQ��n.]��H�.�/.U��"O�=@��3L�t��P���&p�f"O�, ��؇J4$0%�6F�ƈB�"O����`Ї|�Qsc��N�b�:�"Ò�d�V�!@(�HB	�0LoB�2u"OAc��1���2�R=_�i�Q"O���'��%|̤�w�.Xܠ�f"Or)�nȴd�`�%̍O�C'"O�8!�G�
���N�z9P���"OX|&� ?�4�Rっs�z`"O֔�D���\�H��� F�L���"O���ۅtt.�	�����q"O�я�Oqh8�qAޞ ��bS"O
��P� �5�r�7*́l٦d�"Or�����G�FD��)ͧ}����T"O8"�C���⤉��C��4�P"OR9h��#2o��
���H��Qh�"OF�P���_��r�Gާ;�n�b�"OXUJG�3=@��I�Ӂ(��1"O���rB���
C@�'ג (S"OF S㗒O���["�YϾ�#�"O�Y���P;��	]����+ZU!�d�\& 8��̸�R�z����eI!�B4B�^cҐ8l 1{��6v�!��Z.Z?*���<6Rf]�֍��!��M�ܥ�ԋR�:��A�`����'� 9�@�5&@�0S'��:�V�c�'��IX�����Jtk��u��]�
�'a��-7'Q��
��t��j�'$�m�L��
r�j�GK�W{��"�'`�j�	08D�c����T�	�'�Ԁ*�4-�@��̒ r����'�z{��ܥG�1ա�U6:���'�Va���O"*xPa�w'VI"�b�'��æ�=u�P�6)��8?`t��'��A��.w�z&� *g�@��'���1L��[蘸��ѻ)��LR�' z���IG�gʖ|(E��UTXh�'ݪ�!`�ӛ_̀��4H���X�
�'@Pv�� �lل��7}�m��'����1��N8��E
�a=,E��'0��o�*^����a�����'��ɩg��Ѣ���[��i�'���"!��+Vt������1�V��	�'�-`�ʋ� �	��A�L�8�'X�
v�T�U[��#R� ��2�'�VL���(���".Fv.R(��'32�+�dG�&*�a��<?ʬ�'U����aC
���_�4 �m1
�'֖-��f��L���&�˟c��	�'	�� PK߇l����)s �11�'�ؐ��aˀh+��N�m���0�'M<D�ԣ�d��cl^�ze\�H��� ��mN�m�c�f�7d�x1"O.�c� g�b�'��2�"O��10���p�	0Տo��$� "O���!� $散d��bS�P�S"O&d� oV�K�:)�Q�4`5��"OD��OtF�5!���:}��"`"O�mhvLߜv �G���8(U"ODDcn�;���(t��1C�N �U"O2�kJ���a��)�ѸDV"O��C�ґ%��)�D/ܖ.��Y��"O���dN�T��A#W��
BZ�QE"O�9Yc�ߝ��#���&K��i�"O6�J�M�*w��%˓ǚ�f�c"O`Y��ȸ5ENTk��M�E�X�0`"OZ�Y(�y9J�1�]3���"O\� @�^�a��4��dOK�����"O\�B1�V�ud�	l@#Xܝ3��2D�����2w�F�qq���QߦmR�E2D���$�;R3BD��$F"=F��3�5D�4���!gj��&��FC:X�#5D��ǔ�7V|��m��'�(��'D���*�	�|����H�k�X�e1D���j�d�G�ˈIp��q,D���$K�v�� �EE�(\�Q��7D�,����6U�s"a�/P�6|�sB7D�0���/5+0���+�" ��+D�Ȫ�n��h9���i>^@��'D���V����`�ڳ�A�c%'D�0�G�A4Q ��z��ֱ*�P�x��%D��@Cm�>Smx5��G��6J�Q�?D��`�0Z���O�4h�=���;D�`���k��J���2kR���V�'D�`�T�T+dv>|X��N5F���%D���S��R��������|���.D�(0@n�HB�� ����uL+D�����٭;"��:��F���4*)D�,	0"��t��TK��d9V��c�'D�(s1T ʴ��Vj_�#��0r�#D��S�
X�	���{���([9�����?D��Sa-H��pɖo]�~����7D��F�A�w��	���2Y�-	C9D����$�(������2b�3��,D��@�,]=��E�b�$��C,D�$�5�N!-/���ڦY^�����$D� �ʔ.s�D�q���	�����B&D�����`Ҵ(�T(D� 1��E>D�h�3�ܖ8�68r%>w��"�B/D�$��x�&x`��A4,�����%(D�Ģu��Q�آp"�dB ���$D�����t+���t�<����'D��
C鋟NX1+�"�`���eC$D�$@�T*I4�s�Ղq�iC�"D�H	r���w3`��@�E8���*i-D�l�b*��K1`��2������W(D�<B� /e�e����[ۆ�C�1D���lRl��9��&`��0D�$�HV��Ma�j�=hG1D�|�5C�4��� �ĘQrVD"W�,D����U�}�rP�� <�H�)�` D�i&M��~��QaH�0B`��f#D��W�B1Z`p�%a�=@qZ��$<D�tjF䆖#z�%�DI��#�b�*Gc9D�4�Fܔl^쐁tD7pBL��"D���G"ĹeR��X@�ցb��!�?D�� Dh����beJ�� a�9w�x9�"O�,��֙	�2�� �@ڒ��2"O�Jv�͡J9�8�!r��"Ofc�mӾ*Q
�¬�>B�	:v"Or83��-��Xy��V����q"O��pDI�,�^հ�C�\�0<Ҵ"O� z���t��w�/	x8�Z�"O���Ia�<�֎Χ1ohZ "O��9 ��

e�+��8��I��"OJM�2B�w�HudŜU�\Y�"O�X�+X�(�"]jX�r"O�aV�)x��2��\@v8�5"O �B�(]�q���a�]�=|��"O�Xb��(�C ��k,�y�"O���͔��� �Q$���3"OX��p��i�n�$���_Dhd"OlX�DʛD�K^�vBN��2gπ�yb�!]�V�jѪ֊i�`]����y�N�r�De�2Ce�1c����yB�X0��0��oX$n_� �D���yr��2�12�1^B<����G��y�N��T��%��j�xb 
º�y��?l�6y��gF�u+�i�I���y��n&XR�\#j�F�ɇFO2�y�DB6S�0�`���;\�R�
i���y�@O�;Ll}���K�S��{0G0�y�j/x;�̛���a T�4�]�y�
��p���y�e[��X�Ӆ��y���>Z�( ��W�΍��h�yR��W�\qRfɎO�@qB"��0�y"�ޣ3��K�I&Y,�2bė��yRm�Hݫ��ΗC%T��A&Q��y©L�6��	A��>Jrara���yE�(���E��<_�������y�	��,�x͘� 3@��S�Ă)�yr�7ؤ<N��#s��w���y��J�k���b!�"H�����yC\��H����R�H �+J��yBe\2B������O�<�ح)�;�y�Aիj�|�;�)�"b6�Q����yᗶ��%X0���j@�3AO��y������N\��D��&~!��m���+��̓'�@pC��!��,b�*�r�Z�0ߔ�PM��$!��[�R�����+E{��k�K��M�!�J�aQ�k�_b1�#kJq�!�dݏ=�pX����ZO�� d��!�䉌Ah�5�%F�+o?��6��2t�!��'5�2M�҇Ѣ�Ժ�!ɖ�!�D��R�(�f
�|�4 24C�(�!�$lϞ,� �@8u �/ز�!��/qʙp�c�#O,X#�D��@�!���	)�iӄ��^^����Ƹq�!�W�`%�1�Tcνc����cM�Th!�	l�����Jٵ�ұ6m
`Q!��>J�q�d�uj����,�	�!��3c\�Q���#�:���KC�!�/zǼ����fUF���	t!�D,r�j�!�3lŹ޶Oc!��D�9�P�°NV0� :fO��.Q!��i�����X��0b�I�=8!�Dڜw�8I�E�#x.uDb�#q�!��ޥmGD�1�NQQ X���R�!���{�, �6N��3d)cġ�>f�!�� ح��.� >F�a4�
�h�$"OL��GH�v���0wM]
O��e�5"Oʵ���ʫ8�4��v,P�u��}�2"O�Y�a���Ɇ�@�y��0��"Ohmq�� (�x�b�U	%���6"OYc'#ɛ[�|qr�%��q��"O�, RC�:0[�	��/p*q�"Oyp�Ã9]`��hY�G�Mk�"O���c
oV����i�CZhW"OTkb_U��1K��	ޘ�0��}���7�i>9p����X`�u�S�;5��
3�O �/�¨B�L�6�uJ��ɡJ5�H��#�����V�)�6�v�E�MC�F{b�O���ɖ ^��Č��H	(T��O���F#b����^;q
��h@�Twh!�ɩ���KT�5)T�Ys�P�V!��^1c�)1�Gڜ���� �Q!�D�(CV���[�]��qb�F��?_Q�@F��[	<=P����pEv�j����~�'LVl��JɲxvT��'Q4F��9�M<�	�	 e+�Jy�i2�fF/l���nwTLHkԵg^��l�
��'6��v�)ҧ1�Jl�GkJ�]	r�R�P��xT��W@�Ӂ��Abq���\ ^�ipe�<�.O��%>c���R'�,6Z�5 K9��zA7D�H��EבR����3l�qZN���s�D��=�O:��V/ܻ7�$<`�m��(��a �"O
�1�u%� �$���`��G�'�qOa#Ud�?s7��:s���u�����o�'ّ?Y"H�mN���	�H6T��
5D��j1`S�
��{!EX����1o-D��ʰ���,�` ���R�m)�.?D����c8���$fU�wBZ�y��:D�P�'{��T�В-��9D�xʠ�R�N��Y�C̳\O� ;e�%D�\Ya��p]z��3��:%���.�Mx����G���9�E�+ =PA�ȓG�NE��Q���F.E2[}�axdY�̄���wh���MR��)0��٦h�B�	0'��0ᶠB��a"�*�6��C�I�m���E.����#T��hO>���
�7^��!�	�o�Z�J�f9D�<P7�O�+�j��8Q� ݘ �5��|���IrǑgf�uA!��&/�awm'D�胴i�=:�TIЧM����;$�&D��Ӣ�V���qHs'�<K��B��(D�,���5p��QF�U9i�̻t�1D��Ӄ��FB���E��n*��S�e1�"�(O����s��M,f���8fB�2WC��a"O\�wꃔCˢ��Fጴp��8��$2\O4|�T�U�U�x��O4R���:�"O�y�B	P�@H�!$Z<S_>�u��L>Y�s���&����4����2�*�O�'�2�A����+P��`m�,o� ������'�8#}�'Q6�р)@�,�2���e��<��'�<�0A,ǎ)F-Х�_d`Psڴ�~�$<�O��
��͞[�S�$�?`'��#��`x����H!c�2ဓ���:3����%D���nƭ:�6D
#b	]�,D#D���siO�^��U��䆥��â�-D��T�ГQ�|UX-� ��d*�I�� XD �(v��ٲQa�����h(D�8X�f���0���;,�9��n%D��cA/@�03�.�f8j	�@�%D�� �t V&�-MrN�R�K� �ޝ�@"On��ə�w�Z�z��,E��š�xb�'T�5���#��"�A�D�.���'8&<J���PV�7#�
:�#�'����w�Ӿj<0r�тD���2J<��e(����	���L�7{�Ԅ��K?���IԬ0�����m<�"5`e�<���-[���Z�g-V"A2s��`�<ij��[`dhk���9�4�4��\~��)�':z�xs�L�@@���$�A!{�J\�ȓ�b��DnJ8@Նu��D�]��h[�y����<�}&�l#�$X�L�t�hVGڠ_����g;D�haW�\��tRv$'j} �S`I|����IvNd���>
���d�Zv�C�ɴr9�dx���.e��L�dl�2�C�I�*�0��L�<B��1d+	2	��B��vYQ��e�&F���F�>:jnO��=�~zש��N�	q#ϺelD�R��s���=ys��2N@J	�3`S���D�q쓞p=�!Gī
���Z�	Z�+2�|���E�<��@2Yo¤8�)޲�p���,�u�<�p�@��� ��'c���I$��o�<�@G�{���G& w��q��P�<1$Y�>O29Sn��T�XI�%	P�<�e��S�V��e� ;-�\C&��L�<�g�V�@ ��ڐh'ɡ$,R_�<!� �4]BU�C��"Z��MR�@�<�돣+�|�dU�b�H9Q!Kw�<ه�\�l���{�-�>����*Yt�<Y�l[g4���qJ14�t�V��o�<�d�H�J��:��Q6ۦ��E�h�<)$e[,I]:���nɭ`� ��+HN�<����,Eִ��͓�x�N8���t�<Ӯ^*"�`�.�;JI��� �w�<Q�ck��� *K�=3�hRV#�k�<�q(đ\T�l����@L�p� �Si�<	*I�+��C�J%wz\��h�'��x2j�����m�)oF}�b�,�y��].U�8԰p�ߤi,��I��?�M��'��1bEB"����EN��� iY��7�f1Y3��+GJ��0d)�6��O��Q�*B!6����e��Y�8vpX�HFy�ʞ�`f��O3
v0����y�!;#��8#K+$Ԓ�;QR��~��'/�d �:�Xr�)s���瓞ē.�H �Ӫ�y4��x���6r�mZG(<���P�aC����Q��[d\�'��ɿK�>�e瘸z��H�G� S�|c��(?A�+�����K�-Ǽ�e5.�<d�Ʌ���r���L<�C�^f����ǁ?)]�d٢�PT�<9�g�s������;A�@)�휌��	W����}�o;#�؀�Aɀ&Rj	��ș�HOأ=��'3���
+j����V+f��EI�O���D�in�(��K�n|���U�"-�f�'�O?7m�)[��/m�Ⱥ"�ƍF��u3�OV̐`/A)E~0�J��QTuְ� ��?��|"�O0�#����;��C�Kսh̺M�a"O"M:Ec:*P@C�L��du��러G{�'p�FBG���g���A�L���O�	@�y�>���O����*���*���8S��ae �Kg1O ��$�=}fx��A9#ABaa�.�`,�v�'�4�B�4vX��u'W>ӧ�#wc��)(�"�f>�JqCR�](<��4��A��K�S]�T����1C1"�͓Z�X�<�{�'g��(�o�lZ�x1�[�`�.����HO� :M����7�0�X�ρ�~��@IDN�<!M>��O��R��$ݲ��3O��*�\��"O2D�6�9|:n�A��"x��Uf"O�PY�Z�I�!�%&u ���"O�X!�Y!&8*i;�K@�r�+e"O�B���3b�\s֪�."8�H4"O�]���F����-g	��I�"ObI����$�$���_��Yð"O�I+��ʐD��-A(�k�^���"O�,�+��s���F��*[�Y�&"OJX�gj˨w�8��� TH�r"O�����N�ax6���@!��`p"O�MÐ�V$b$P30h�/gz��7"Od����̇Ja�ݱ�&K�ƨq�"O�0�B����ÒE�9?��9yg"O:�s�ň#�] ��Bj��a�"O�q�V��	G;�����j�0��"O����⟗a�Tu�A��C8���"O6��'K�i�56Ǆ�J���"O5*��[7o��9�'օ]$��""O��ۢ%�Uɾ�J�K/>�z`"O��[�R�\Y�\�t�	1'��"O���'A14�@��ߡL `y�"O�ě� ��1���:��"O�����\��
�u;�"O�4QP <��\�q��;��2"O �jp�h.�t�����L|�Ჱ"O`�ः^#H�@�0��9g_�p��"O:�B6��=�}��DT he� [�"Of	�7%�@�@U����e]��"Od8�3g�E�,8p�"��4a����"O~HywHR$$��} u"1@���۲"O�d/*��Q����s����b"O %���ѝC̔a��8�|�30"O�c��2*qz\hêO;S����"O��aWy�0Ab��Gl��aa�"O6e��]�_�DP2CU�[����"O����1#��� ̀�WY�zq"O$��]Q�<�5@��w4&k"OL�ᱠ_�pa�))GNM].N�jt"Oщ@@>�ص����� "O��G��?7_l4`�l�9ftU�"Oʬْ�0h�<��B��zk�=��"O陵����e���;g���"O�e���L�D���/Eb^����"O>D @�&L	 O2W�P"O�L0�MT�%d9+uG%E�l�'"O����:�d���vb\�b"Ot���(&K~z�*@�\�5~�w"O�X�W  {+f�p���^����"O�����D�d��f�Fu����"O؁�W	�;�z�s��~܌]h"O�('%+?G,��Ga��2-ن"O�Ч$Ӳ�4��u�|ʎ1�4"O6��Fĕ�_� ����.��C�"OX�J.�M�8!�vF�;��y�"O�xH����"e�� �N�#6"Od�bWI�&�>���'ަb��@�"O�L5��4{8Mi�'�/r�°��"O&M��gM�"6&-���
�`���cp"OH��p��׎��m�;��p��"O*�P��W�w;�8b�O�8d$ u�"O���g�6b���F���c�� �"Oʱ!�O�e�9�7n�6R����"O� �Q@v�A�4fT!+S��1vA�X[�"O�Pi��ҺҘ���E~����"O�����8�$�I�P�
܁"O杣�(^�Yڅ5o�� d�S*O�}��.��2Rf-�7-���9	�ܰ�����<�Ms�*�=#/����(�rHS�l�G�<I�Ň,�,�7���SVD`���W�'��-��hˎ\�]F���ʦ}���b���)g���%��yb	t� �R�C�/��(8���x��R�Vh2��*O�}� ��zS��c)	Q���!�`�� ���Eb�K�*�DC�-/R8�I�X"&y�$�CO2\ц�9`Sp�(C�Oώ��VHX&P�����H�m��UbuL�cVte�$ѯPV�Y!i@9�t���$<D�q�JԴ!ʎ�w.Ȁ%H<�,4��O8u�'�\q�\e#Z�>	9mM6[����SH�!B�&��Fg/D���Ro�5T��x��Ş9<s�^)�^m#��X�T��h���ī$4�b� d�J})�A8X�H⟀G�?�g~��ߢA���"��U}�Qs�?	�+�.G�ܩ U���<D�_e<� ��ߺIV��y�O� Q��h�#/O$Qa���R�.\�ǃ�*8Zֹ�d'�?Ekޘ�#�$/�d��DX>@`ʄ�K<9�R�<T�	s���)4|ۥ�Jb&��<ѥ.
a*�
�c%�	]��y�(��}��[�mߟ|%�Y3_���~"�ekq�?�)�)z3$ ���̈́~�!�R)��!���g�B�+��L�O>�G�±*��D�|��~4ll�ǀ�W`I`g ���Wp� �Z�2.�\d��e�#z�{�O>�ScLF���ԛg*U�"J�O�y�K�-&��I&A�,����3�*%��'M<!2� � �8��Oq�6!
�'�Jֺ���d�a $�Q"�'��Ec��|��7|N�(�g%���I��@�'bHE���/}"��kD��o&���HW�u��8���78�:���]et#��ʍ��xp�I��*Г#&�;�����.�O�<rwNR����f��3ry��'Q�ѸF�6|u�'F��ZT�\R&�hR��L��u	
�'*�S��M+Z1T�;D���q�^{I>)@F%r�PC�/�':T�P�"�7X���ya@��8ǘ8�ȓΖ��uEf"@i󥅂1Q5���8��P 9G��O��3���k"�A#�C�$Eh�"Otr&F�P���+=�"�V"OV���\Uk�G��W�˗��y2�R�p��Y�&:�ҵ�d��y��M��A ��Ӏ���I��yB<y`�+G@Ѳ8��� a��y¨ D�T8�4M�`�3����y�� �RX��BQ�t,��  �y�f�y��t��&J�t uʛ<�y"e�0C͠���%ئq.��T(�;�y�eH�3�",�TLK.Q\z�1�-��y"�w,��T�@'e�f5�B��y��D�T4��䈍v_�!��Ǐ$�y�f#l� 8Z��o����-*�?ɖL ����DJ �4+�����2����a{��UC�H.�~�J�0��񫥧 > (A��.��y�f�
/�������" �d�e�O(q3� ��6��������t�j��w hC`L@63mv��"O6t�ՈIJ�����0O��%d�5]��|�>O� �DQ�^D1�1O��21�@L��ӕ*�KL�@��'���Ah�lpLݒ3� <���@��S����v��.>�����d��GV��yB"��(��1�L U��1iQ����O��
��I7�Z��6$�/H%��U�f���J�/D*I�`�*Z���b]�@�fA\���<���{�n ����%!�\��/KYy�,V��P�@�K�*i8},��O���"&�@�sᮏ^�"TJ��یSXA��xH<�
�.9��[SM}�8��$A�U��Š����8�G�B:N�$9�
X+3��{s�>Y�wΨ��u�էP�D�a�	�wˎ�y
��5J�M������a`:pO8%q�I�mL�P���@
�C�$�R�đ�?��i'�)���W�d*�,N��z��X��|"?��f���pY����f�bU`�π `q�.ջ	\�`m�<di�T�xQ$��62l`�ڰ�'m��S�ހ�Ρk�d]}�H�[�O8p�n�*&�~�#v�]�7cq��	e�D7��4!j 8o���D�
xS�I��D�x�� �V����� בC��}rGl�z �s�ڟTOZ�t��h��A �S���ɂ`7}?�`-Ӏ�B�`�b�R��!dÔ�{��'M��b֡�&
�hsB��3&��HQC͂K��y��@J7'�(C�(
���ɔoKB%h�������d���i�L�s����� ��?��/���իt;JL�C,���d�mC�9R�
�`�^`*�����ĕ6@Ć��t&#<Odi8��N&Y�a��+�1:��0�Q��
��[&\樑�eD(�<�d�I)�0�d���Ԅ1�kԪa���ʅ(]0�yb�[Qv�Zg
6_�H�A��I9.�5)�/t� i�(�WR���J|�>yW�T5=dE�B�b]���n��@�K�(PYF�����#2~�p'B�2eZ�I@�z�CG�u&�&�j�ǟt1O��{!f@�`�"h�blP�x��I?f��@�OG�'��LyV
U����:�����@<kj4�v��$Yhk���h��"MDԤ1@��'�jr���b"F���ѡR�%s�'��;A���`���@L1V2)����@�X3�Y�B�84{�l�A�&-J�6��!�I�w�& �u˟aH<Q��ܠVb����� �R5z!N\2�%*U�X
,��9�j#���q�]�Sh���Т��B"᎝ݼ���4�"���)W(��R��X����w� �<�`J����E�+*V(X�g��8B�h�#L\0��BB4x�*�q��K"�	���j��$vL�r�%Z�#�X(� ��0P!\�>i�AT)tR��`��(�,3e�&sJ�H�
<A2��Q�HD7W� Yq�Sw���+��v�\HS�K���<a#%�-�yu��w����^`?Q��ө^�K6����b��p�4��q :c�R�PЯ/�`�@s�K�L�2p[�H
Rn�{�G���x"�	�<x9)T��l��y��D�f��@ѡ#W�G�D=ʖ�MKZ|*fI	�6lM"m��a���ŧ�y���P��XBⓀm��5��l͹հ?1�
Y��,��$�'/ <򄬋������(JGv�s�B �Nʰ�ra]�ɁI��6=�қx�������Q-N*Q�8����;��O pbp�Ǵ;�J�� �ا�
�;�%���~䂴AA�{�LPQ	V�<H��J���"�,��<1�K��5?ޅb�&�q��]�E"sy��Eα2e�
�D������g$x7�ǝ'/%�����ľv#�l��'6�Y�G��/Ef�ܠ�I�j�.�;Ń�~�^���O�Z\�4i�?����}i
iXv�H�xQ���Qǈ�l��b�'��G�$27n�(�A�C�|с�O]�p�dUc�O�'���Q�E�Q�~D�C�ǕN~�Z��>LO �)ԃJ�>A�	(}����ǉV�N� P�$2ޓO��d���� U�!�>�)"�@ U��������л4�\?Ϣ`r�A� E&\y�.�JR!��A<+�0�P&�J�̓�m�Ma��\I�ɏ0�"T�}2v���]�Խ���E�(K�\�<I�Ӕ1Kb0����nE{c"�f?Q2#�l�Ұ�W:}��� }b��ytɌ�d@l���3Q�!���f��2	J�@ԁ����y{ ���𤟻lQ��tmL6�<q��@>m�Q���6��mPqO�}�uO\�.����,��m��d�2 �;�\8�t*�xb��:I�L�g�B�<_�%"6aǭi'���l�;pS �೅\�crԚf�ٻJ�T�s�E���Iz�i�2��P&�)�%�@+�8S�	9D��ЊęF��@vI
 #��$s���J�Q�M�d��8(�-L�Vd��i�H��R,�B���'����W=l�p��B-5E�X�ߓ-о  ���^���ue�F 8�ڤb׆.��r��cTR�x��Or}��K.oa)Ó��8F/��PrN��̍�/� ��?a�E�31:L+!��8V��x�O�$��a�[	Z@��bp�ȫ_�65��0{aX��U��n<1'`�:��1�����Dq��"%�qrp�S(޲k��u'CZF��Y�Л|Zc���ǁ+"hZ���Fc��'<��r1��uJ�L�G�O6c%B0Q��v� G��3��Ot�0g�H~1�O���W���X`$V��PT�'����^	AS��n�}q���{�]��+��cS��+�&`�ג��<a���,'����|��4�'d�&~�<��W8ZL"=!�d	��)ag�mY�� ��A$N!��T0C������Bq�1��9 �L��cl2OX�:��Ӓ��p�H|�;B��|y�fǮadȴ9�HϜ,�
=����=ᡧ�
��L��#��l,�U�I�|:pЀ�M�+9�Ӻ�s�Rf������&Ǘv@��:D�>��8FI-D�l�!��U�=���I�*��=KC�<�����!���k�l-,O� <5��,Z:���J �	�e�}3��'�acNR/�\JA��#NobpU�Ǝ�`B#AeH<A4͈5�	v��j�Tc�s�'�Us�GÏaD���~��K[��&�0�Z*�s�<!TI��`$hYZ�F�1]B�����\BV$h��5�>E�dAG�G=�]�1��*R����:q�!�$�6V�Ld�$/\�.""YBჭs�	�AYNP�`ĂGx���GU�k(�q�'�E5�\�5�?�Oh�7b��U��l02%��Qh�
Ga
7Q��h��'��)iq�*LRRPYP+E���*�'C*,;�ϒ9Khc��J)?�pli�'0jeۡ��]�������*5�ij�'�x))�[�A����"1��S�'L�5�b�_�v��FǏ2$�Tu9�'���9��Ә��� ��Cz��P�',(������y���6D&�"�'ṮFO�*F�X���$����	�'\�8��D�`'ɂ7DO�):2���'�t��s(C�͌�D�2u6�h:�'���ц;�,�F�����'~Xa�e+��c*��:QOJ�	jt���'B�EdI0Nz4����9u�����'�����jː2����g�43&�`�'�"���)NZvf���cҝ*j���'v�0�sJ7V��-[��5	t�5��'��2T�
2�%�%��+ǖ)R�'� 刦�ԡ,A��	��	I�TE��'�p�g�ǠUA��J�Nܲ8k����'��̩�k�?�ph�5'��=L@ �'�p�ZgoG�v(i
 BF4BX�
�'����l�7��z`��'%��`�	�'������Y��X��ˆ1L\h��'"2�Q'��\��b��.��9�'�T�1P/ۂE:RL��	Z֩�	�'d`���eke�KS��R��}P�N"D����/@?��#�O�?|d�U�<D�HЂ�F�N+����
Q�l;�/=D��d� 0J\�5����%,D��
��сR�,�!$��N��ٻ'�*D���4a�\ɮ�����8k�b�t�&D�أ�l�-�tC�]���P�$D�����a8��Z5���O"D�,�D��7�x�
�N>�5D��!��q�z����L*E|F���b>T��xA.Y�z����&����"O���0.Ƅh���)B�c|Ds�"O��s��0x<<�v��w����"O���d�ʌlג�(@��7{���aB"Of��2b�c�@e��L��p3�=h"O�M�!�/l&`��5	�#^Cr�1"O�L0V���k/���j��R)K�"OцT�+W��C��E�9��a"O�$W��-j�ͯz{T��!G�Z�<!����J��U�AfI�gg4���[�<!�'[�Z���6I� ��aB�V�<A���?r���B
�z�4AI�H\S�<�&�1H��:��I��8�r�C�<���ځCq�}��"�� 0����_B�<Y��L�>�G�Y(b�� n�|�<�pE�!\=�k5'��(����C�<q�B��:����&M��**�OJG�<`��CU@K��{nhHy�K�<񁣗�zH&H�2�L�d�u�t�	F�<q����(��$"	��<Lq'}�<� ~0S��T�C'�%���T.0hʥ�"Oz��֬t�|�&bK�7Gh���"O
	SA� t�!3�N�6LZ [s"O�Ly@��#6��ƯF�WLA�"O��JA��+�萐�Y��<y�"O��r�IH�DD�C���p����"O�d�����/e��r�G��Rv"O�� k�2}$���Ӟ�xR"O
Z�U�p��5��3�^���'�hk�D����i"y�Pǧ�2��ӥ�yBl�Q.*4qQ�����Zk�0�Ob%:V"�'�T\`��i	�@<�@
E�݋{ *���"m!�d�>Q�ya!� 
���Q#w���#�nX�E���P��G��'Ե�U훜,r
���*e� E�'�����|�8�X�̜nE�(���q.F�7�ҏP�������b���9&��,��5]}�̄�I2R�H`������C�L)E�N-�E	A�
�&�I��C�<y�HSZ�.J�-�&bl嫃CC��}p~�  P�<��I ��i!<�8�@�M�}�@�HL@�o�!��;M�|���X���d�E�4,:���4IƊS��rAX��D��'Ңt��f����3�h�]��0��'8�X���`�J����E���h��d�Y��5F@Hӓ�}
Q%S L-p�5kF�B��I�[�jX�`ʄ��y����/d�������
,�%��K�<1��5I�t%�
�3L���B�B�jT�<���R�A�fH��h7�)E$�yw�WԄ�"�G";0���X��yRMbb���Ā�li�%PT��`׌�	��F�lO�O����ƯmM1�¤�>^��%�F5���;c����<uNƏ0���3�>��=E�vP@�(��ڂ�n�<���ۿ����U�-�:x���|�.�,D��Z�y�?
`h�f`pz����zל̊��=D�l��.ȣFx�-Ң��1�F�R�W4l� JL�� E�m�g�$��@8
�pFS�U׈ A�A]Y����gK������sJt9h��1e��`(F��8�8]�P]��9)!U���2�Æ�G^6D��ɡV���
W�$D]�I�Y<I�Y�g1��0W��	��B�Ʌz�H(�ϕ�g���� �;{L�O�������|BH���I�'>2� P��U��N�	Vś�-�!�$��5�J���M3J������t�vdx3�4��Cv�>�F�Q3���L�<���# ���u� Ԓ�W�?s��$�[9yP(�ȓ$���CIWC���s�ɳ����6`�P���^�]C�\Yc�.5{VD��@�@�Z'G5d����5�ǰUƬ�ȓJ$(��G�E�pn�3�ЭKY ��O��%ٰ�!I�xLa1C̩G�,��ȓ[�L<Q���Nsh�x0̏"/�$��j�ƈ��A4��1DkH� ��U�ȓn�bg,ej���B�TB�$4��sб�JS��%�SA!�2�������C�d��T`�����ȓv\TIZ''S�rܐ��<?k���*a~��GE��<�H"�N �T����xV� z��'P@})���3J�I����6�2ѓۓi5z((�Fئ�~Rס1�l�`$ Z�����	�y�)�wh�0���Rʮ�9��ϝ���#��U9#�8j>����q̡�s��!"��t��a��C䉌^�B,S�6����k	�-����k�0f�:�8����R�?�3�`)��jq��]��������d�b/������
LC�`0�ǩ�*q�k^�y����
�!Vx�PzBEB*=1Ob�����5`H�V/ܿ|����iѐ	io��u� �	7�P�|����{0HH� LL�l(:��Z~"A��,�t�@d�'���ì~�J� �	�G5���)O�1���3 ��h��m�꒟� V�Gm��L���Dcj��GMA�H��hG�B�x
� ��0$�_�=���*��ӤHT�iTe�F��]���'6Qj@�ԘCP��p��ކ9����O���ʌ�'h�����F����$ɒ�Ҹ����"�^���,��a���26䝸�M(�����N� � d
<�a'?*�o��H�* �W*J�XxѢ��y�'�*�꠨ޫ,;j]��3�����(|r<H�/�
����_
��dU>0�� W��<���*H�x%`eD��4x(\��My���"���� ��:E5z �}�����3�8iEDO�`���K�S�M�@x�E�^6A�B≻∵P��A耉D!�.K��'����T
,O�����ٹmґ�I���;5Ҍ�))\�t(�5mˤ4���iDШ`��A����'�V
>o0����
g��*�.x4f��K�8D���^�Pf�AB�ģ���p!Q�4O!�Z$���RgB����3�-�"��,l1�%�',Hx��iqER9��,�Fn�:N�h�C��$�Ol8!�E�I��A;:)@�Ů��H�2��'�x��D▕@���E�k�'�eH��#^�F����ɛ+���8
�'��h�"��tQ>�R��
�a�Qk�'D|�����b�S�O-�z2p\�5e�9��	�B���y�䜥>�Z)B���27m2uJ���_�gk�p�4<O��o�.`���F�
� ��S�'��#n@J�f�02�6B�p�k�U$^�� *�HH<�W��mo�����u� ��� �]�'t��)Z�h�b�~b��X=	��!�*k/ڄq0 Ul�<!`D���@w�� ���3ܟ�c� �r;��P�>E��/�4 �4�)EG]�(���x�eM�B!�ƹ%,���Η�)3��ՍQ]G�ɻ]���+��Dway��3xv�9ǖz�A�դ��>��D�Q��뙑�؇�A>O���r�IQ�D��C�ɫ/:�!�`b�'���C"�R6Y��=a�*�dB$�(�I$��(n��uq�&v�l�����9x�B�@�(�5�E$Ez,0�)b�$�^%R�y2G���)�'< �8k2@іGr�T��h�0p|���
�'����WE_��d��L,$[�O2p�F)�4 .��D�*h���AT+��Rb�	�����Ca��@%�S�4̆�cQ�ߌX� �b @�'�vC�I�@���T�G�
��C� �O�zC��;sD.Yi)!*������FC�ɞ@t�r�J6XAXq&P�K�PC��.0��ڃ��=�"�AH�$9�2C��1p��A�S�)	��;��L�%�C�	�4׌��5�e��ze�����$��5Ո@�dML�Q����K�j�:�$ϐx� �:?�h#�5.����������O���q�[C���>��vi�Q�ЊpG�(+k�\�1�1D�t����*6T�w�B�TT��'��Pa�a�>X氲2�>E��HN�?�����V4y&`��ׂъ�y"�1Ґ�c�A�~�P��'��;��	���"wO�u�ax�#XI��Zp�"z�ZX:G���(O*��cؘɸ'��L�Ѭ�'�t	��i�4�I���u*8����@<Q�e
>y�ɺ��)<)�����Z����,��Z���QǙ�nF���O�R�	�T�6O�W�����ػ�y��.����ߜ8��X�q�	�?��b�*�����4��I�BR��Cg�_��rB�"ņ�tL�4y�ᅅt����DH�tJp�(� �M�Ս �-}n� �
�Q�(XI�L��#�FyJ0�?�0<��%ϥ`Ƽ@�!LZsI�!SE�� L0L�@/�HĈ��<l��O�Hr�z���t����Y��p�Ѐ�W/�x�_�(6��q� �eܸ-��,T�}*p��"
�'�����Q &���X�"!t� �7���D0�.���y��:�t�rF�(�詡-��?�s��/`���ڷ
 ��/a���ʗ* �$�0�(r�	Ǭ:TU��H���{b��4�0yp�Q˦q�Q'��/9}��"��K��2?�N�&@�E�ϓ1&%�a��~�
��Q�c=���?)WG;"lTb+"ғ�����Ϛ�Nݒ&�L�J|؈AO�agP�n�� � y�*�� M���c�)R��'"�K�'�T�f�'>�=� �y��H�4�� pf��A�r��G"O�0� ��[�p�Z
���$��'p���u�F�a�J��O�.E�M:j%M~�3�s�0��6H�TnN�x���4�ybMѿ�B�X�h�0I���h��[���$�"j�<�s�BE��<ibg�(n��ӥ��VCyh�d�px�p@�$׳ zB�ZIհX�8�i"�K�m���#��1�!�3N�(�P
ӘF�B���*�ў�§��%@:���i�/S���A�R�<��hw�!�dX�8��U*��	oln��S���}���q�������|��S�S���H=e��U���?��!��1�n9 �`G.E�.�ca��Ms���'��M����?F��y�J��K�#�nRh ���c��p?C+PP,�QAh�4])���R��T8��?D�tx��ă �wŅ:z�i�&b.D�|�pH�o7�,�����g��9a�/D�|�7�\�D���M�I���H*D��藯�~	����Z�Tri�r+D�<Y�̺KX�*Ao�Y��
��"D��jU�~�+ǏX&s�!���; !�߾4(=�$nI2�����I2w�!�$>k[�u�'	!b�b��r�EW�!�D�k��A�QH�3@Œ��!���� L0��;�
������!���P\$���Cݹ�R`�%b�39c!���9�6�s�־Rn��9r�ߦZ!�3r$�9��0Fy�I �㇒En!��C��I땊ܹp���b�.1�!��[4#ڍ85�A	% ~���	�<!�d;7nⱈ��P�w,tIz��޻R�!�Č3��P���J����E�sP!�D��a���rrhK�L`w���W!򄗈Nf��֧�
�$􃔮�}B!��T
�A�AH�Q�+�?Bj���aG��� 	�z���"�E	g�ȓ@mr SRG�8#������w�m�ȓ.6xz��ՅC��)р	�f}�������΁8��=+S�j<��ȓt�̄z��
W��5�;񪥆ȓ��9�i��|�T̈4BX;v`}�ȓZ
�񠐈��u�D�pBJ��+^�ԅ�6e��h%ǔ�%h�A(�	���ȓ�\$�BhŤ+6A��L[�9�D��ȓBb�]�@)�����K��0Y�N��ȓ>A�T�6!ӱ!4e)��ٲ$״X�ȓ$U���d,h��ȔJ� 1@ ȆȓW7�\ȶ�B�NLp 1��81�����V�Ȉ���4	��e��3V�d�ȓoY�ɒ��7v���6��-W�Hy��B�q˶�߷�c�I9�Ѕȓf��,2b�� vf�Z�O�N�,�ȓI�P�@�O,"�q����'1B���!+��SP�7muXDaq���8�x��N��J���$�3�䤒p����j��W�	M��T�2i�	v�׈xD����%-�a�,��t� HzC�T!g��X2�J0w��A�/�$75HzV�ͥ � {�����-Id��C䞰_�����+�CߐPH�ǎ�M�߱v�~�Kd؟��i�7�6�*
|����Є�	5U�R��@�U�8�~�$�[z#}p�T�~��H��8L�ԡiуH*�J1�/�\Aj���'<����S�Q�`���;��ܛ���G��5*�:k�5��)iʄp�!_>�ȟ������+�q�k^�R�����A�Hh��I(��A�7�ۘ
�>y�O��:0�Po]DU�G!�4y�Aj#;O
��y2�i>E�/8xhb}QE/B�O��ˀ�*�>�O���e�~����/�?�6��"O����C8l=��b�G++�� Z�"O^`�bB���<S��7?�%2v"O� t��k��W���UŽ36��h"O�y:���h�,=2�9r�"ON4�"�\�%�ґ+��1&�j�X�(E{�􉑏�hDz �;����B�,M���'�?���-R�i�e�fR��>��� �	D}r�O��T�
�0�;��M��OF#=���	ւP�<A��)`/�d��OT2;���Sd����D�PR �)9��Q�b��F�z��Dh4ғ�0|ʕ��]Ȇ�3�AE,E�a"-�_�7Mў�'?������4]�$ݭ{m���<�����^�W�p�5�4��\�W(�>z��J��n��6���(O�d�!d���i�6`(� &��x�oB�8�l��K>	�O8�n���1.��<;�鐝Sh��6+R{!�R KH~�#t*ڗ#NV�R��ԫ�!��R�*t�Z�L�� �.Ł��E<n!���$�R`���߫N����c�	.Q!򤎗/�\�F�W4x8�p��I�3�!��G%e�,���Ȩ+!z���1 �!��/���y�灓:�IEGV�r�!�Ҵ/�:�ئk��~��BH�T�!�/I�!x� /!�&5�g��//�!��Z�	;��%o�� �R��DL?g!�d�i!n};e�N�1�N�{���Ws!�D��TW�a�� B8A���9TBBn!��]$>����%c�R�R���^U?!��=pA�YPF� ��LW0f&B�	+�\����#��@)��H�ƞC�	%z�݃��
�6\9"�z}�B�ɯ*tDՋ�G̪k�R1
��|B�	;R� \KF�֐(��YHS�#);*B�	����� +h �)���.B��!Z�� ��H�����i��B�	'����ha�-E�\7xB�"c=`I��ߐ��� �	�!xB䉍c��ܳ��˲IO���pď�	`B��D�F(ae�<G��9Ѩ��c[�C��>p6�KTn�Z����Ϝ
p�C�ɺk��YJ���&]�°ȣ�-=D�C��df�E!�M�4�R���a��DrC�I6QZ���GM D)"����ZC�	�|���c�/Z%
a�p��g�]�$C�I/�X03`��>:�x�F3[`B䉕�8Hإ��-G.������MFB䉅PP��oO�.(�I4i�@(B�	�z��8g�M$=$Ȭ�m�r�C�	#F?8��F���ytA o�B��2PT��K�5��(��M�;#�B�ɤr��x��	͢��P��J�t��B�ɒ/]ܜ`�)�*u�A�'�U,fB䉃;�~���F����DsB��X�C�ɏSČ�Isa�o]�����R�C�I�l2HBpL�X�D%94��B��J��`⪗1f�m�������D@�,}�#)T�mr�h�f͒!�� +x� �Ņ�XP<e��lڿ
!�Қn�*$ �K�R� D�sҜ�!��� H�IK�j�+��xplªP�!���%�r��Ƭи+�ڴ��8�!�ʽ6�rx��� w����Ŵ:�!�	(y}�J��Δ3L�1
6�ՙ+"!�D� ���,�.K6rM�F�T>\ !�"[KXt�BC��fPxu� �`!�$B3 �ޙ����5?4��0̟�r!�Yr*X9��J�?3��xCjC�K�!�� F�
 ���������S���A�"OL ���Á��K����0��2�"O4#�NR�,�di� �ݷUs +�"O")#`g0f��]`�%�6r�~(P"O����.Z���Q"�}�J$Z�"O�p�8zQ�@Z���-/���"O �
������[�/� �Z %"O"E�b ��g�����g ���"OxQز��+=��u�4Ý��I�"O@}ڀk<((�i�� u�@��S"OZ(�`D�wz�� +�+'q��"O.q�R��
��YF�8m;$���"O�Y�#E� �IK�jN���ã"O�ak����	)�Ȣ��O�4��r`"O8���%�S9FeKw��nh�*'"O��Y�^4b��X����:T�=�A"Oޠk��άe���A���	'"O�q$�1p��P�Oԭ}�0��"O>-k���)Bz}!V%T�q襈�"O(E��#C!1��Y��EI�cF%C"O ���:RRI�e�C_�x�"O>�Kר��!�� 0$Ke�(!��"Oʹ�+�'�Ы��hȸ��"ODa����"�$V����"O���<%]�Q"K�H���#"Ox�����QH(�`2�����V"O"5�u��xP��1,^�eh0��"O�8�i\6�:D� K\|�hC"Oԩ)3�K�;޹p�X�zh�@�"O��q��4����+c�\r�"O|�k�»p�ᗈF�G��AЁ"O����6ܐ����N<��
p"O9#m@�>�Z�S@k߻o����U"O�AQ�C
	Z�~$��i���n�cF"O�M#���vC�u�Q��50�Jv"O�! W�<k�]Q�蘮o5�X�"O̍"���'e�t!��Y'd*�rW"O��B !�n����&才=`,�p"O�,0�h�#3sfP궄�����"OV�zaD��M�ʉ#@�2K�ڀ�f"O.�[uH.��$���{� hȳ"OZ�[�H��%H�ƍG�&�б"O,Xď�!>�#�X����k&D����gL�)������]'j�H�j!D��b�J�Xy���R�R��d� D�����:��%��N��b�*p�"�=D����FӇA��@���Rah�}�g@'D��� ��[y��(�E�l��v�'D�X3�[0SyhP�!�����;D�`�w��h��uK��܁E�^��ȓr2t-項�(M�a���71�I��/'*t�w8��4�ڊ-����>�R�!p%�%�`8�I̓]}�ȓ<�ʱ�"҄Ij��!м9� ���X���OiAn΀n��I�ȓ�$m�#N�A �,�ǖ=�(��FR�1��e�8i�4u(��=w>d�ȓRZ|��g�Z�p�����y�l��t*�� �ԠX�D��Ƙp(^������6��G6�+5h,��ȓB=�'jS�b�H��U�\��^Ԫ�37�q���0eP��͆�{$<�4E��|�ԘВ�N�\����)Vr�@��/M�Z(b�B%|���S�? h�x�m�.-����6�p��"OZ}[��N0�)�u���@�"O��ړ�єN�֡��S�E��p@"O��s�_�G�Vp����2�Va
v"O��ARDQ�l�d�c�OR�|P+�"O,YZw��!UJ*�qb��j����"Oy�Q��t^��aR�,E �(�5"O*PZ�(�h�Lـ�<BA�P�"Of�b� +Ί�(g�c2����"O�i��ґtLPM�&*Sl q"O��P��60u���9V�4�g"O��8kE�X�803)Z�+�(���"O��A8���C�4��{"O4�H��ˡn�ق`Ō=&��Xے"O�w�d�T���W�X�Za��"O�UXǈ�����P�ju�q2"O.t�X�`���ѰXSb��J�<���I�y� "%/#�p�^�2B�)0�p 4꓋^��9��%̉4z"B�I4#��FkJ�@B<1��V�@C�I�nt|��7egz�:@g�� �4C��h�m���Wo�
�z��@�Vl,C䉓�i�T ^�vsި�n�+m
C�	򬱲ԮS��P��͞�$��B䉎��Y2�?��Q�͜�a{xC�5O�(���٨ ��S@猧;�XC䉦u�6D��V�k�-!ȫ_C�� 2���3��T@�'�ӗC�C�ɚ�T�6�����Ti�E^�C�� 	�'��%4�{D��-
h�C�I S,�a��
7�E�4�O=�C�	�6\�C��R�H����K�NجB�I���)L�K�2�(���

�B�	�V�Р��ˀ1+��0�O
�f�B�ɲw2X!��Ŕ)7�Fl3f�F7X�4C�	����0�H1f�L���8bC��@��9�'o�.
��)����,C�I7�ұSU�V7i��XR)�L�B��$Ra�4h$�E5=3�h ej\�e��C�5*g�P9�&I�|�td���W2��C�I6�0<�L@��&�c���$�6C�8�^@�v&͑t�V�ff^�2f�B�Ɇwt*��
�wS8��'�צ�|B�I�j��1BݾZhS�┰H�B�&o70�:��VA�h�D��TzB䉪5R�3@��|�0H)7�=6�C�	��\}b',�$��u���RIjC�I1>}X�ز�\�En�1H�F�9~B�	�Lr C��6G�H� ��2�C�	�)� ���]�P�̲�P0*�B�>��H�a�ƩX�H(�+ܖR�C�2!������N�x;$��>�C䉂&( 	ٓϋ�7b(�2"��~��B�67�lhX�)l��8�BӁkĄB䉉R/���'O�<W�)"K�2e�B�	�y����#$L�d��Ah�&,�B�ɒ#�d,��M��|�� 7a��nX&B䉰:A�5)�P'U`)0� 4#B�I�=���3H�,e\6�Ҁƃ{�C�I�B4�Y�1Α2a�\�s/�O��C䉶a�΍B�s��|12�A=@��B�I�/V�|������S�k_h�xC�ɘy�ptc�)�%4%D�×�?hbC�	�f�V�2��h�T�P�(C�)� ���Bi�._�SuEˮ=�z	KP"O6i)Ţ�j���z2�Z�{���"O�`��T�#���C��c�fE)"O��	.�x��y�&"M�4�����"OQ���+q�*�`1K��x	�"O䙩FJT�H8$!��'`Dp0�"O� Y�B�	�x��Ơ��9%�2"O��gT<�����(�J!�7"O�E��HW�xt�3E�$=,�A�"O>mҷ@|8+�l}:�yU��k�<���G�p�KB˂�4lA�nm�<A!�=��0�g��$3���;օBg�<i���:��[�aR%	}$<+R��b�<�S��7�
	A#�{la��N�j�<��
�8*��s�,W~�4��6��~�<R�8��E�(_�0!�P13 Eb�<��A @  ��   6  *  �     �+  �7  �C  �N  ~X  �b  Dl  Ou  �}  �  <�  }�  	�  ��  خ  �  \�  ��  ��  &�  j�  ��  ��  2�  u�  ��  ��  �  � J � � ?' +. 6 �= �D #K gQ �S  Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�� |d��"O
`�(�;���8���-0��1%"Oj4��ND^[��"3/9�0|H�"OB���H��*�ʞRy=a"O�味V�!X��!&F�:J�$���"O,��a
���C�Ą�M�"O,$3%o�-���p���+Ն�:1"O��ݢ1����`���y14]2��i�<�6��{_���c�H�`�fX�$Kn�<��A̼VI�xR[�)�Ć�pඤ�ȓA5��('nߡ4�� �)˩%� ���,��r�؊b#`T�eT09���ȓ!�b��g��}�8�F��-? �ȓ
K|m�ș�VṔ���2�%�ȓ"R�X�j�4JN�1�˘X�i����̹	_�jZ��1!g��zܶ��ȓgil,*�J�
j�Ne��i�J%b���f	�(U��:���G��$Y^م�~r�� S�%T"���k\�jx�ȓ|4�1�îJb��@ӵ�ݩn�V��/[`�"�v4�R�!ʎ<��M�ȓ`:��z�ؚh�J�Z��$HY:	��H��p�m�C1��!��B:��0��EnjZA V;9����J[
2���	��4'J�EA�IVW&��~�(aZ��ӹ�>� o�Y�|�ȓ�f�A�
Ο7�H��M�$�����mޠP����/���ANXo*�ȓTv�����{ ��-7�*h��I��sB�8�8���3����ȓNe*M�悡;������X�o��!�ȓ'lj�#F�m�+R&;�|��2)n�C��0S4���T:
b��>	�����R�O����Ί6h6Z��q�R�y�I$m��d���>a/�0����m�Q�,ێ�Y����*�.�\�§�@�"��ӆ�<D����o�!o�(�Kݷ#���RҌw�|B቞Kԅc��#b�*�m�Y"���"�	�4x�+R	OTL`r��:|��B�ɒK;�Ѹ�/��#�`�ꛍ)��<��\���L?���U������j>�dL֣4g����ȟ:/�}ϓ��?A��+a��M�Ӣ�=@�q�*_x�<�S� T��X�J°_z"�)�Ëu�<���Q�
���є��f�$��Č\�'L��o�Of9��`�.0q\�`
Qf��i��'m�d���R#h�4�,��u��ّ�'��	x�)"M<Q(ғ#*��R��~�6`�j�<��� =�4�0�D�w���.��<���r���$�%���_��b���Ɵ�>�2C)�|��?yz�xjUf}��'U:����m��5��<z=���'`�{��+?D�����vx�L{�'������c�8�]������'ˆ!�ݬ���`��9����'&��tF
�i�l���UB#"�(�"O���vL�,=>h�M��_��"�"O�u�C��6�d�*Vk� �(�"O��zE
l�N�J��"�.�X�� �S�Ib@��"KJp�(YR�ˎ�zX!�$D�p���/۴��@���(g�d�O�㟢}r��H�r�,��$U�A�ЗB�V<Q�S�? �M0�ûp�$A�KS?�����3Ov)��ZX�T3c�V Xp��iKP<:#&@y��7�O�7m�1)R�
�ӤB�#���lPp�eO�9e�� Qp��v/V5\����P�I�����O�^�u�H����R�A!kt&*
�'��lQCj�h4�YHe�s�5��'E�0��xTٰ4)y����F�<�t�ԨQ�dP�ART��Bc��]8���䁙U�<{��7}����<�O�批{�v�Hp�۪1Yd �%�0j��B�	C4�SI(V�p���ǌ(V\B�	 ��Z�b٠sK���r�����DE9vJԲ�(_��`�RbC,>��	_���6� �A߼���"J�0���V"O(4R�jX=H�h D+�6!�'�|R�'-N��g'�к����AJؚ�'������Ej&�)2ጋ�'��M;�'�dQY0L���P�3ϖ�E�:��7ILh<i4'�/A�z���T�\�����IM�<qB*D
V6SrO��<*Fx��,[F�<����xѯ�Ndũ5�G@�<���R��d�gEA( �A�/�x�<��#[u�m � ^�W�� �Q��n�' �O�OZ}��'��P�jZ�'�H�B�'�����^�x��ɵ7���AŪ5�!�d���lH��j[�j�f�j!	�X�!�d]�R�Ft���]97j)��T0:�!�!,8�)*�M��D��V�P	:��D{ʟ��B�4+ڽj��_-(`��G"Ov�	pf��IX`"In��'"O�i0F`^�/W��X�j�.��fP�Ѕ���tZ�G\�p�` �
B/=�#=ɏ��^?�v�Y����+D$#��Y���Qs�<A��r����U���j��V��M�۴!ғO<�i>��B���HhZr��N	XIu<D��p�$O�Gp-����)Le�We��H���6�n̈��.��4� � �0j�\�Dy�Z���'��'7\�*�a��RX֑c���U�l���'��Ը��*XAc`�R%��zJ���'�ɧ�O��9��,ZF�����N��
�}��)��ԙ@������q��J�28!��V�t�#�X���+�'��!�$A�P�6eY���|�Xr�Z7����s���%G+)�P�Ba)�����#��}��dԄS	n�8b�Dݡ{�v��gf��B�Ivz`a@ �!B��W땵��t���'h���@G_$.g�aZW(,yH�"�'\(Xg�WI��jF�����ӌ�dc� �=�'b��������Da�Ȫ��Hq����|�V����4���㟥;.�bܘrB����<�
�Q��T�dw��`�	D�&��J��1޴��=�d�&'7�k�Rh����G�<��E2]7��@�9�,قG@�'l?=R�eRFT����1^D�� �>D�X@��	� ���U�<`�b�>�S�)�'�< ���N�a*A��o�U��`V��&�Q�8JŐu�ܠ$3��C˜x`��8T�Ap�U
���<aI>y�yb\��@g-A��]���
C_��`5$�HI@j!Q �Yf�u� �����0<���$ϝ	s"Y����.Q��,��F�A!��,_��� rdC}6��Ԭ��ب#x��}j��Ѹm��i"�h��S�F�c���~��}��ħ�?A��Q®�8נ@mt�I�$�z�q8�� �1�-ʼV<n����%�X�y�|�i���'U��8	g�ہi>B�pD ݠs��!(U ��x"gD�ho�YI1�]68G�dRTɘ2��	R���O��`w�a՚%0��[E�|�H	���y2�[14���J�35X!�S�/��O 4G�$R{���WD�.����#���y"E7`�$���ȇYA ��� @#�yR�Ѩ5<�fB�H1�"r����c�l���쟒*�4��6�Pb*M�ȓn�x�C+-RqBx1E%٬���ȓ28�����ZRl���/��<n*���I�<d.	1�z�ɗcH9^�.�	��O�<Q��Q�C����u�صY�����mVW؞�v�|"e�W���[��̥^�B�p3���?Y�'Y %d�?���0Ǖ&-��:
Ǔ�HOȤk�O�)h�2�P�҈;�M�r�'0�ɇg^����Q��1���F C䉱ơ�'�Ȧx�I�􂃲	+
�>1.O$@�p�&�I� c|L��ܒ$7�0QubH�=��|�����E͡^���"��s��M�Be��XF{�'��'�l��5�O���HÈj�DՁ
�'D����սQ��L�t��gؾ[��d ʓ�����?i��Šp��7+�!�]9X��PCC�g�.��c��."����Y��`��`������Bq	��F|�ӡg��sO�w{Μ�@&�3YE�C��4t�Lb��L&8�Č"4�W�S؄7�9�(O�>�nZ�t��t'޹�|�rQ�Ё,q�B��53�٫f��f�P��͚`�b��<ʓ}$�H2���GLT����>_�F��ȓJ�BL`�% aa��ֱc��ȓ3��@ؗ�ͬcY ��f� .W&RT��a0�b�"��ge����(a6����W)a�ȍ�Z0b  �ֺE��ȓ7��m5��o�L �� ���p�ȓ�艄Hզ:C��;����@�⤅ȓО���`��.�� MJ'�͇� /%!w��a�����ؘA(�݇���C���Y�|�S��ҹv�Ќ�ȓ����sc�]b�a�7n���I����&ϐW�
��D@��j�E�ȓD)6�Yå�9]E�|��*nJ�E�ȓD���c��ӫInM ��[Et^ �ȓBк`rĄ�z�<@!���X����u�(����_1��VO�4ഁ�ȓa��lh���nV:5c��TX�b���H�xE� �pO5��&ĊMBN��ȓp�0h�/"js��*���_���ȓy̍����aDtjJ�� O�t��dƠ53F��41�U�>RԔ��u%���P���V���e��7.�ȓ�*�C�N��f^]!WN���~�ȓ2�V p�@(�(��0#��2t���&<I R@C�Y�H	���c��ȓ1�v�ք�%>�x��1�3U9���ȓ�Rl�3���gȱrB�0Ƽ���}����jII���yo_�C�Vi��4X
��S���AЖ�٧aŪ��ȓ@��V�^�2%��ɡ�RJ؆ȓR9���4�߅"�ec��lȓ�^0ې׀+�1AIӡ�,D�ȓR�21�I�&y(�cK
�T�1�ȓ+��Ѳo݅M:.����dD��c��q�� S-+r�l��OZ ��5��S�? j�1�C�kW.���Z|�d�#�"O"}Ж�Ӥ5�(@"�6�q�"O�ͫ�н0�A�4��0L�"O��Ig��.W��H@�Dl�}��"O�0+p��!���3�#Q%bVܨ�B�'3��'���'��'�b�'(b�'�z��A2 ���U�؉N��$�'a��'r�'0��'9��'q2�'�t��%G�
PĘ��/�$ =�@���'Y�'��'���'5��'v2�'�]jէ-�i3��?0x�0�'��'��'���'��'4�'���zT� fF��W�%&`��C��'���'�r�'l��'2�'X��'�&��$��)"�Da��	l��u�'�b�'Zb�'���'G��'�b�'/ι����>�И"㏚��z��6�'���'���'2�'fB�'{��';:��A�?z��0�$oQ�\e����'��'���'r�'hR�'���'�b�a���GcJ��A�ʠ"D|�V�'���'B�'��'���'s��'�H�vnY!�C�D�u��s&�'�B�' "�'�R�'���'N��'��}�W�ìP�����[�YI ,I��'�b�'I��'�b�'&����i)�f�7/�*���ӹGI� �q�'���'�"�'��'���'_��'�r� 	B�p�NHQ�����1K�2�'z��'�r�'v��'��7��O��$փ	9���)�(FS�u٤��9�~8�'��U�b>�#�&+�,�jk6�Ȩs�$�����Rl��O�PoZ{��|�!(��`�	�d�J�oFn��ʠE����7��O&�B��q�f�N2�c
�k��Ov.���HL�&h�Ӧ��;�H�z�y��'��c�O��(	0�?RR��R/�9(����h�攊�=�S6�Mϻy���,9[��;F"˱s]�͘��i�`7�l��ԧ�O����G�i�ٴ'Td��"!��%k!�13�@&`��B���3N��=ͧ�?Q��<A� ��ٞA��+s"�<�+O�O��m�n��b� kF�U�Yx�T+gS�^���c@r�� *�I�M�@�i���>��$�%K|�h��6��#r�t~��j�4je-�=��Ou�����A�I О9+�	.?|���`�D7x���'��	��"~�U�"�;5.l�%Ô���h�Zq��Ņ���d�צ��?�'	h���խZ7�ЙSO�   |�>ܛ��a���ĕ�z:ܴ���I=	�H�p������'@�9s���볆�("�s�!��<�|�<)�/�#��eo�g��9�&Cp~2�x��U�@�O�$�OL�?!@�'O2g6��v��N.]{5-C>��D�����ܴj����Or�|q�lգ��E�ʟ�<F|xBs�9�Xi��\����EO��İS�h�a�I\y��1e'��3�k��#n����І�0>��i� �x��'�p X�i+D��i��O��� ��'f�6�0�ɥ���ަe�۴T9��J�q�Z�;r/]�]�p��ƫzĘ�������S-X�,Y�)ߪ\G~�� ���)�+ZXQ	��ìo�j��0g	M���BEd�
_d|��/�����Xaq��M�9&�S�aȌ-��*�`<?K��\0��@�,)
9|��$NM�j�hE��b�j �@A�Vެ�P#��@�8�v/',ȥL�%&i�Ua�5p�x #��@��0��ǁL�P	�	�9D�Pĩ@��7g �Ĩ�c�;l����G��`,�F�I�|Q.i��gR�L�����Ȑ���	IՐ"auk$�Lk�T9(ଞ?~�,݉SeW�Pΐ4V˗��ҩC�+�;��$B�"|L �k���6A���f����Iğ��i]%�a'?���X��4D�t��PT����E�:h�Μ�>���f̓�?����?��mA�UF4���^sz!�G�Jߛ��'����Q.�D�O���*��ƂL�Pb�	�d=P[He�F��q����6�^b���Iȟp�	uy�.H�h�1{�a��^EH`��=OL�	6�0��O�d*���<��@'KC�5�s)_9���DD((���<!���?!���䂊�p̧�\��)?���3dH+B�J�'���'c�'��Ɍ	���3�8� cƇ,,JD�rIQ�99P�'"�'��P�(�v�G3�ħL/��S@�YO�����Y�y�N0Pq�i��|�R��2�$?���,�V��WD�/�2���B�6�6�O��$�<!�KH4(�O-��O�V� �~��Ԣ��+����#*�$�<I�C@I����U�c�@#�ʲe���N �~I�&P��i��ߜ�M+�T?��I�?�r�O�M��cU/ h���7Ҥsмiw�I0t ��?�g�	:m[h1�c�.^�*�!��Z"h7�",��n��h�Iȟ���ē�?!BkO�v����b,Pl\}��1c����S�O>��ɽO�Jx�u�X�Q��T�1�E�	�`��ܴ�?a���?�(<��'��'X��ؾa�X�%�!o���GA^<O��O�Eu���O��$�Oh���F%d.J����H:�`ZD)Q���I��P\��}�'wɧ5�N��!�Lz�ϐ�Q�¡C'[��q  8�ʟ���Ɵ��'\Hp�v��3W�t�J"U3�L0��S�a�O`�D�O�Obʓ�~�&�Z�2}f����XS\HE9@��K̓�?����?!+O�����|*��G�Qڍ�3iV�t<)Bc�x}��'���|�^��KA��>��G�q\~I���ќz:9�2�q}��'�b�'!��
tԒ5�O%�h'� ����U�x>`�1'������i:�|��';�$P���'q��s���Q@����eM�YP*:ݴ�?����DD�)��˧�?�����&�:�����~�(�4cM(R��'�2�'�2����T?�	�꘻*J8,Y5��;W�`���n�X˓3��B��?A���?������Ҥ�6�?p����#D7<#���A�i��'QB����i��e�����6E�n�P��)))��Ɩ�[U��'.r�'{�dW����ԟ�c�J[�g���僅�h�0q(@ρ��M3���������3"B����'D��]�&��-p��lZ����������tyb�'���'��d�}j
��p���=�ޭ+�L�FE�V�|"�;�������OJ�D�y�h�{� �N�6���kL+9Ţ�lZ̟T(��NyB�'5B�'ɧ5�Ᶎ)�0d����J�
}؄����č�e�6��<Q��?�����Qw�¬Y7�D5[��D"P��.'|�`�+Z}�V����b��ß��	�b������w�Z\a��f)�g�]@�ݟ,�	̟h�'��-@�ҟ��x�#�9��Eaj�a��i�"�'>��|2�'?2'܉<����<b��)��B:	�\��4���˟����<�'����Q>-�I�l��5��
Gъ�v˂WՀ|Y�4�?YH>����?����'��yA�jڧqH��9u�>7-f%rܴ�?	����n���'�?�����*>p8:�N�Ah�٩�e�t~�'�B�'hN���T?Y��aJ%,���g�Fl#@-q�6ʓ*��|+��?���?	�'����I=Y¸��V�/Pe$!� �i�2�'>��6�����"Ү�M$Dr�y&�6<���K�H[$6��O��D�O�iVD�i>�vF�<Ǫi���˦Baƴ�u#��M����?���?a(O���<y��Y|�����=MN]0(n*,K6�i���'%��j!�O�)�OF��\2o\8�h^K<��o��w�pxm�͟���GyB��~�'m��'�ba�ǓF��`��M:�H4jA�v���D8䦭%���ޟD��{yr��#adu�t`Y%z���r�C�~[�7�<���䓨?Y����-�v�:t��]a@�V.��vd��m�n����Iԟ8�'�"�'@1���J���d�� ��eP.�KEٿ|3b�|��'r[�xʤ.K���$�e��ɢ�Z�x���E�(����O8�D�OD˓�?��_���j��R�)RV��*��L���#fX�B�Y�X�	˟��Iby���!�&����k��rL0�0�z3`ɂ@�����I����'�2�'O>M��'��6#����RI��� 5@X'Q\� n˟�'�R��y�Sڟ�I�?�5m*�X�"Z�k늉�t"߁w!�O����O>�+1�:b�1O�S3HRJ�U��lFl����2\h���?�DH	��?���?����/O�lG6@R�oC�l !@�A�rI���'bb֕���*�y��Č	&|�p�&I@?g��Q�C�-�MK'�Luԛ��'�B�'e�$�:�4�k��+!�!�$!O�(�<��GN���n�"_NR�'�r�'U��Y>ŗOBXkk��|�����C<i/��X2H|����OP�dҸ[�S�$�>��\�t�Fd��VD�w���.�1O��2soKZ����؟�C�%Bk[ֽ�E�� z�%y�b� �M���q5�Yw�x�O���'H�	kA��q������Ǐ��v ��4�?E%�!�?)-O���OT���<��� `@.�5��L�
a�A��>��M@1�x��'<��'���ϟ��I.�LF��;fTb(:��΢x����wNIߟ'���	ϟ�'F��zGH>�j�T�u<zQ#L�D����̲>���?a�����O���Ɗf��D�sG��!	��T	�-]�fǲ��'���'��U���@�.�ħ}y�@:a"W�9F��r���%����if�'O��ȟ��Iivځ��t�	ǫ����C�DD�*�g	��6�'��P��!�W=��'�?i��3e$�~$Z���l ���G
%]��Y�`�I埼h�+E�&?��s�E��삸j"u���}�,���gӔ�Yk,�C7�i�|�'�?��' @���'�����<7 �q"'��*g�7��O���^2k�:�D�q��?͔�M�C�/(8#CN��*���"�EŦ�PT�(�4�?����?��#Ɖ���@�K�� �L�L.~H邡V67(�7m��Pm��d�O2�$�O���|�'��F��oP�!�#�d�(�!&o��$�OB���&5�%��S۟,���f�X@���4�@!�NX�� �z۴�?���?��J��No��F�t�'��D��Q�`�PC�.�T�ہ�U�O_���'�$-��U�����㟈�V솷E̲���ޮ[���p��ގ�����=�� a#��O<��?��`���	4iQ*+��Q�`߶X
j .O��D�O���I��\�4� �$��\���z�$y�D�ެ)ܲ��1?9��?!��?	�q���i�lm��Eŗ/����'k2s�ݡ2�t�X���O����O��d�<���2W���'**��hd앜y��͓��.:qR�hF�i���'3�'���'�P��O{�����O
;��2Sd`��R��A���ڦ=��ğ\��^y��'P.�K�O~r�O��
��H6�x9�UEK�}���P�i���'���'����Fe���$�O��d��"�(�O�|�$�p���-�����/�����I[yR�'�U�Olɧ��4D��`�M�EL4|��IG#m�"Ho�ޟ��ɓp�s�4�?���?�'���Bi� @�0Q��d^l��Mݦh����[�$���iu\A�I@�i>A��@��H��=�T�F��2� �d�i���&�g�����O6����	�O6�D�O�%��4`�Iq�ɔ�$�Z��
��=TcD����	˟�C��ⓟ��$ �j-����늮g.�(��m�����nZޟ|�Iҟ�����M����?��?��Ӻ�ҎY"�0p1D�]`l����Dm}�Q�t��F ?�'�?����?i��<h7����c7T@H1�baBg����'�n�aehӼ�d�O��d�O��O���7D� ����O0�|b�A�8/��	�1�8��|�I������(�O�n�XR��!P�0d3d�B���I���-��7-�O��$�O6���w��X�h�	:�`¥I� D���7Jv����fk���Iٟ4��ߟ��I�	��U�شLx�ڱ㒃5�^%9�(�9��-0�i�"�'�2�'"S���I!ol�s��-�$��!��-[�E=k�(욶�i���'���'���3��m#�i���'��P:�F�%�A1�]��4��$qӠ���Od�Ģ<���f̧�?a�'��-s%���c)�)˅�
vٶ�K�4�?i���?)��_�=Ѻi2�'m2�O�\���֤X+�-���<���v�Ӽ���<��ms~Χ�?q.O�i�έ�PI�y�*���`b�%��4�?a��q�1�"�i�"�'$��O��D�'T6X��>�r����xH0��D)�>���ZvJ���?�����))�t��-P��)Bo��B\����?�MG�ٲQF���'�r�'����O���'��T2^5ܩS%�DY0���ΐ�kK47Ȓ���d+�4��������l`\)$� <~)ڔQ��<[I\�o�˟4�Iٟ$�`)���Ms���?a��?1�Ӻ3��pD��ES��8$��!ᦅ��Hyb����yʟB�d�O�����c�()���^�f�4hs��[�8�o���ΐ��M���?����?��]?U���&x��
X�5>����=P�`$�'6�P�'��'*b�' �[>�ѵ�ۗ=�p�!.Q�/������c+��rٴ�?Y���?���[.�}y��'�<�(��ABfP��Ϝ,Yڡ�ѽ�y�'��'HR�'a�S�zܴ5����	�K�x�6�T1cG�Q�i���'�b�'5�W�����hm��NH>��t��,`a�!p�Âd�.��O�D�O����O���� �@l���I;Oj��@��#�%�0��EQP��4�?A��?a/O��D	��)=}MB�`z��%�$�<�r��M���?���?	!+����'���'-��,�7e�$�^/�(l3bI�y�h7��O�ʓ�?GÕ�|����4���h&u���Z����Ub ��$���M���?�d*@�Y?�&�'��'����O�rF]�'�`L�a
��.mx0�D�F�2��?	5HD�?A����4��O!İ��H�qC:|���ǐ�\�ܴ|R�@�i���'�R�O:���'�r�'�l��f�)�~�+Q�Y���EcӔL���Oz�D�<�'�䧶?Q�E�$�d���J�s|��2 �=I�v�'���'��a2�b�����O��d�O����6Ma%�� {��xB ��3�]�c��M/1O��d�Ol�������He�Ő�v*�cܧx��4lZ���8Ձ��M��?���?�BX?E�D����a��T�D�A�W(j���'���;�'��	؟��Iß�������a°�l��#��8��4��kB%u��ٴ�?����?���:�SAyR�'Z����>1���/��h����9��D�O����On���O����,��n&
��H��߿#�Yr���)Zh���4�?����?a���?�)O��DB�|�	G�op��� �D��(@���|��nZԟp��D�����)I���MmZ����	����#5j�(��p`��)`���4�?9���?�.O"�d؅|�I�O���H�(M�v(��IN�ط���7��OR�D�O���� �\n��h��П��S<J�4K����<;�¤B*;P=��4�?�.O���\�Z$�)�OH�D�|n��Lݺ�p1+�";p�H�g�r��7��Od�$7��n��P���T���?���Ȧt�A:P?.�s�Z+P��<R]���I�\����џ����~
��%kL|�1���L��'�L�A�c����M��?a��r�'�?1���?�si�8 ��0��ҦR�y���
V��֌Ʌ�r�'��i>�'?U�	�F4Ѡ@�l�x�EGN-LF����4�?��?��ǌ7d��6�'��'����u�e��p!Z�h
P� ��Hײ�M�)O6��[�M��?��	��ɍp�40���K� �z�!� �X�Z��4�?IP�P]3���'q��'h�j�~r�';�2n�x���
�Ќ�$�����",��D�<����?�M~:0JO�<�Љ���d �]�'�Ƽ Q��
�x�'`�|�'a"��B8J$12h�|��Q�A+ϛIr`ّ��'��i�lZП�I`y�◚A�f�S/u_t|�D�,�����K�Z��?���䓤?���ld4u��/:�1��ބ����@�ӤHMh�* Y� �	ʟ��	Ay�	J�}�N�J�zd BX��F����h�bJ㦡��q�ԟ��I�*l�=�V�ֹ@�X@

(�ȤD�ݦ��֟D�'YbM+��<��OJ��Թ	���֧�Z���K�cF�d�bT'����̟����y� '���'$@e�
9�.e�� KG��'��Z��d���Os"�OcH�Mf�i(p�@�~��|���Yy��ynZ��I�=�	u�)�S0D0�c�<X���æ�ۭ_H"7m� �ʁn�⟬��ҟ��S��ē�?1�ӽ\|��c�̐o����C'k|�F��K}|��i�O0�9�@ӆ�:�B"A�qK=l7�6��O8�$�O�L���T�������w?� �� �ޖ�lu��)V��`�i�'��p��'��O��d�O<��i��X�T�
'+˙}W���ͦ����>�D�"K<����?�M>�1[yeЁ
��Oc���ݞ�4��'��Hj1�|��'�r�'��I�o�$8G�ߍ ���k5L>D�B�O>���?����?���md�^���p5/Բ ��Ā��?�/OZ�D�O��$�<9cP�;�ɟ�.��q��Y8K~��w�ϴu�	���	{�I����v[����k`��Pnϙ�^4��e��/^L;�O����O�D�<Yv�ߏv�O�( #P�o�P}�s��t��y��*p���d<���O����ev��D0}�'^�6 ���;��	��Ӣ�M3��?�)OB�`���o�Sܟ���#^�SpIX��DYS���1%VْK<����?�"A��<�I>�O58����m�@�B6�D)&}��ߴ��d�!P4�<mھ��)�O���S~��a�R)RRh�($}cU;�M{���?�c��<YO>�~
R�E�z��-�t)8d�-R�$�����D���M����?�������x�'(�Q3!��+��hr˙�O��%8 {�x�aT��Od�O>�	�l2^�#S�r�H�赠B`r�4�?����?�f(>͉'#�'l�$��&�z]��ϋh�:�@3o�1��O�Mi��#���ON���O���W�@�x��PwBK)��������ɝ>�n���}b�'�ɧ56��&�5z�ぅ<㜰(�����D߈]V.�D�<1���?����򄊞L*|�+`M�58j�e��,)L⤕���z����LF{"�O2�r1��0/OP!x���Z�4Y��im�V���ǟH�IZyX'#�$�SD�]R3�Y���|��AT/���?Q��d�<!��=��h�CQ�r�� jFM4|;�0X�Y�D�������by�H%��X� �̑7���kT�J1[����q����D{BR�h��c�	W���P�X�* As��4՛��'"�'iB!Ư:"2�'��' ��]�x��BE�zD|0q(	8΂O��İ<p�U��u�W�R\� b���H2Ä�Mc��?�Fǝe��'2�'����OqZc<�1q�Cҭ$� �{�,�CS��8�}�U�d��H�M�C�7�r�14蔺L7��N^�A-��'���'����'rX>e�p�X�;�hÃ��p����#������ġ+r�b>m�	�T0����Փd���7@�I��Q�ݴ�?9��?aq�36����'���'M���u7O��A>�%;4eWu���
F��M�����. �?�����,��l�D���f�DY�c�3-�In�՟dh!l���M���?���?Q2T?��q��	q�e�,m/4x��+�-{"6��'%��(�'^��'��'��'b��>S�:�Ʉ�?H�T� �T9Xg�г�c��d�O����O"x�O�����x�E�G�=�t��,Z.Ż�(��P���vy��'��'��'��ʢKt�x���	"v-༉��^jp�ʧ����IޟX�	ʟ�IQyr�' �؁�OG}ZҩDLZ�ոP�8U����d�8��O����Oz��O~��8Ѝh�2���O,�h�+>�P`����t�Ŧa�	şh��my��'1��O�r�On��& ƉI�Cè�Fzx��a�i�B�'���' ���#`�$�D�O��쟊	�b�n��e���B�y��i'�PϦ���Ay��'>Ƙ��ORQ��s�~�����$�R�8�K�6`5ig�i�Z�M�S���cc�F�'�B�'=���O���C𔘘��5+݌̉��J��?��c���?�M>ͧ���K��yff�k�̱�ӛ{�6�C�8ߔAl������l���?��ݟ���4�P�aC�
�H��EHQH��S��T`ش3�������|�O~b��l�`��E��تqb�w��2%�iFR�'="n�R^�7��O����O���O�.�:�^�����u�6�D�[��'��v�@�)����?q��ղ�I����,e
6��#6.Ke�i��_�D9 6��O���OB�$@�4�O�A��U��B��3���].p�@0]���֬i����H��ɟ��O ОfQP���Y,$X0�Jب��juӰ�$�O��$�Or��O&�	أ�M� �A0�&�{����Ь����ş��I������X�O�z}��g��!��?z�b�S�BA�b���0�Xզ�	Ο��I���	oy��'@�ۘO�����&B���Sׅ�		Q@�.iӰ�$�O<���O��$�O~}���ͦ!����H���G������b�*Q8�����M����?Q�����O&=��7������[��z��A+"���j����hӈ�D�O����O�4	�%]���	֟�I�?E0�+.#���Qi�]R�Ɯ��M������O�i6�v�O�in��&��sč@�g�#o����4�?��;l�,ѽi�b�'���O��$�'���&�_��e�%���V�>Q�u��!����|"H?]��B�6~-v�H�ߠA���4~��8��Φ=��Ɵ����?���ӟ���ܟXlZ�t��U��}�:�bӁ��`z���r��|�O��O����	�r�J�^���٣�H�6F%�7�O����O�]�Ʃ[����8���4�i�����[�<���"�*�s5@ [sw��D�OD�Ʉvy�?Y�Iß ��"n�rىעܳ'B�KC��~d�0�4�?�J�j���'�r�'��B�~"�'=.�Q�dB0y���23
J��#�O �Z�4O��d�O����O&�D�O��ɉP�8H�� ���h��Ɂq�ʼs5�Wæ���̟�	���j���˓�?Q�� 	I�hN*	���*�H��P�`,��<����?���?I��?1��;���W�i9s�/K4��!�Ί!}m X+#�u���O���Of�d�<Y�����'zY������������J�)�Pl+�Y���	���	�D���2p`�@�4�?a��lN��f�2��j�.��{eY�i���',�_�����U:H�����f�F@Y'��7�4��6�ǘe��In�ٟx��Ɵ���-;�l-��4�?���?���PD��Dǌ��n�i�DZ�FIt���i��\�0�	�,���S󟰔���4b��T��k�$|��x�	�<8�mПH���e�mbٴ�?A��?�����_Ռ��W�NMH�Z���
$vl+Q�t��T?��	{y2Q>���j���O�
��i�2���FePH���igp)�p�����O��dퟀ�i�O����O�;G%�0(ݼ�����;��R����B�����&���w��H#��r�Q�^8�Pl�q T��M��?Q��/2Īe�i`��'���'�Zw*�	@�˔~c&-"���%%�x2�4���O|]07O�������@�K��F�����H�"��%q1m���M����Q)c�iH�';��'u�꧟~r�]�c�iQ��A�y�٩'aY��M��/��D��?a���?���?�+�Z(�d�����-l7�ܩ��N�KF��mZ�H�Iҟ\�	����<��6bT����(GD��ʒ˂-}n���)K�<y,O����OR�'�?�6f_�z��6(U�qa Sr�9?�^����if7��O��d�Ox���O���?tɁ�|R�Q9Bo�l�7��(�TL��(Bc}���@�IƟ�I�H��g�<�M����?i�� I��	�Q#QDT����(0g��'�r�'��	ȟ��f>��IX?�T@O�0���D;� �P�R���	͟���ܟ$b�����M���?����� �N(Jn�����(g�)�C
�{C�V�'��ߟ<��Ow>!��Ty��MkQ�
�R��E���P�k�@�̦U�	���В`]��M���?9�����'�?Y�lχE��}R�KݦK��x0��y����H��C����Iby�O�.^�G�\Z�Lس��Pj"�"$�&r��U�UD�V��t�d�T-7v8�ҦL�>`�ŉ�ES����e�
%H�	��$���]�V�B%�"OxX�U�'W��ñD�G�%���EW�����=_�@�Z/Q�6��
�-C�Ba0G
�[$���5�@C�\Im�Ah�q�3f@\���rL�!V̮M�D'[�3]x41$I�>���o�U@ڕX�e�A��%��N�+B��`ç
��w��H�0�  O\����$�Htj�O����O��$�̺{���?1�OV��a�����rv@q��B*��ATŝ(�jId��;��<I��D%�Ф�!AóO�R"[�^賲��.2���G�:fay-�n���܂S����e�}�p��rZ���vӞ�|���$��Y���r�F k�N��w�
�y2�\ Qx�覆J�]9ҕx��Ǒ��'Ǝ��� 	��Y�'��z���dkp��S(Y<7r�'Mt�ئ�'��6��%RA�ڐ}t�<�Y����4,WDE��?@2X$�#�H@�~l��ɧ	��u���2,­��̦��U�	�T8r�KJ#e�� 3�*&O\��a�'�"_��K"k�_m��
J�Rl֌!��(��b���Q+��2| �0-ӿx����(��C�4,T�x�(C�AGtIFG��u�������ĸx�)lz>�	g�tH�H��H�'���зo��YS�%����'���ZM.6^�a��D,��T>e�OM��C��Ӹ��I�S4ƌhH�d�u�Խ_�PE�DH�G���Xpn��O!q����D����C��$�Op�}J��cfdP�C��:�	�*C
�jL�ȓ0���P��|M�@����qD�d��	:�HOp��M�>=����f���1�D|�VF�ɦ�������I*l�P;���ʟX��۟d�i޽����<1�A9%)�jt��H�#H�<\]�f��?!�AVCS¸�|&���qЏ\֤�	`E\e�M3�e.ǐi��kW�?����44��>�O  z�Dހj�L������f@�C�O��2$$M�i>�G{�Ǆ�o5CJ#zO�V��:�y��ʮ`�ā�S�ٚy�2�p�M��D�L�����'�	�[�|��O��|�Q�햑e3�y�
ʙn����	ϟ��	۟l�Xw1b�'_�	�0J����j�b4�d��OǖUB@$R��z���hE@-����$P�L���FB�!Ct�c���KgH]x�͈�yK� [`b[%t��$��y������-9���:�K�7H(�Y��'c�����^���NۨD�d���EJ!�$ضZ�pl�7.V=7�T��@>1O��l�V�IE�ݴ�?�������OJ-n��,վ<. -����?A�n��?������Bf�|s�.�W@%�2�*�,���	��Vj�5(�:{�b���ɶgZ��9��ۨ �4����?q�H<I�Ñ*)�4I����(o��!���'�����{��'v���Gר D���
 �j�Q�'j#���$5�Hi��k�t����'�7�N24����Ŏ�^)��.F�"-�O1�Q������ʟ��O@e ��'2Z�@R�ĺo��r��Ӛd
<��'eK11���T>��8�
!�05�d�����%>���O:u���)�3� ��C�O2:��hv舙Li���>����П �<��K�_�
�C��jhmY#dk�<�B�><@��V�ru��h��ɉ�d��2���eJ�'B���C���'��'�<p�t�CuZ��'A2��y�/��bvl� _PE��:�:�<e�
T�>�$�0a��19��|���?Ul r�A����A����.�5�RE?�t���ߚ6�����IA5s��%H%�B���h�FZ�9�z��شXX���'>^��v�����D�O�}Q�M�:��MR��H�vd>x	0#24��t�3���bGGȗn`�g#?�2��x�DV���ʹ$ڑ�0���M��Y`V�0p���k�\ɟ��	۟L��5�u��'��0�N�#��}A~�R5΄��L��6�&R��8��Ͱb�����D�y��ً⋁�5et�J���_`��E� ;�X�� Y���I�@v�'�١ۯA0pX�,ɖ��baO��?I�'t@�Ç&zY��"�⊭t4�9
�'�,a1"�K��d�E=�@�`�y�bz���O8PS���������,�(¤1w���a��t����ӟ��I�{ ��埸̧=s�᱑�Qg0�)� �A8�&K(���53n��3%�ĻZ�~�X���;!�\@4iK0��xڄt+�,*�dS�[P ��� C�@�
�0��Y�!����촱BhF% �txH��
H�!���s�E|[ 48v�[0��Y�	:�I�#�]��O���|�6����|1 � J�8tӤ�Ҙ#�@���?!t�ϫzF�IA΄�NCР*���ɨ|��(u�d�1�^�Y 1�o^s�R�]Fj�c#�ӴE^5Ar�B���z8�*p���Bq�Oc9�}YQ�>���Xߟt�ڴV�>��S#y[��c���5��m�b
��,��=<�`h�o�$V�`�Bt/�PU�ቬ�HO���cK�ްd1d	ݶ�N W��ŦA��ӟ4ϓ)Gj��F�Fԟ$�	���	��uw��_�������=5>p3ÃTa�`��Ʌ`}�e�"*t쳈�L>A��CH=��tژ2�e�c ;7o� ����{��E����� �}��.?����HV���s�@?_�Z�Qd���'�R�q�S�g�I#4a������{<��5��!R��B則"�|��!_� ���LX���HO�))�d�B���G�H{�4�[q�	pOV�i�W���$�O`�d�O��;�?����B �9�N��J_4u0؉�X!���!�vHѓ��#��=Yu�\3 ��#��j�������b|��0�D����T�ߓ0Kt�B�M_'��б�4bT����M����r)�(G ��{U��-$5�م�Ij�ɭU��A���F�W�ʍ�!�~�b�pc޴��$,h�ִiG�'�B�B"�@��5�a�n�!�R�'r"�E4wB�'���ջv��|B�ʸ&��\1%/{����*�p<a�C�e�'��\�f?�4��� R'����ɚ[@��$!�$��N/�ᡕ		ƽ!�)�-�!��Wc�I8��� ,����&m!�$��I��D؟od�*�������6f+�e� ��޴�?i����ֶV>�d"iSH,h1MS�ԽY�����O�,�'ܟ ��&��'��	��;�^)��-i ��LD*x��rA8�Q��ѐ��S��0B��`)b� �I��[H��O4	"3�'��Ԛ�d��o3x��$���������'���'1�|��C�l&l�%!��$F@T
Ó`%������� 8�"s��V�x�QեC��M���?!��i����?���?I�Ӽ��a��'/��k�P�jn�8���	�')T���y�(�C�ˈ�H/�9*�G\T �=A%%�Rx���ʚ2��H;� �'�  *���� � 0�)�3��I>kXHCt,�)0)����,��K�!��?C[��3 သ[!4x���*��	��HO>�c�%��0[܀���@0�(F�X�߂9�vc۟���џ$��2����ON��_���6�ECm��_��-H� ���b��d4b�$IfВ������`ENv؟L�f�R�������W�k�2�n��~�L���O ���O^��?��B㚴@��Q�F˜9?I��"�$E��y��۽s�p� �&���Df݃Ә'E����$�6��o�؟L��U���UgJ���K���|��	��T���ޟ����|G���M�Q0Ʃ�4���	�}2v�*�E?:��|95��TL���R�$��#�&�X�'�R�qf�j4�x���Կo!����`m����⟐��� v�8%�V�y�$��̊Ng6��Q<Od�$�O��"|��	Y��B$��o��9�f����[G<y�i�eh��P<81ZiT��%"9�Qa�'��	�&��X�4�?�������6���]8�l���";J���t,ӧ�<���O�5�`�V?y��勰�_���T>a�O�l-YP�1
�򜀑c���jl�J��@¥˖~4&M�w�6������ �Q� 4��h�P�"۞���	�t�$�n�)�+pZ�����)�إ���Xo�~B�	s>X�p�F��4�̵X$��<N4����Z|�'�l�X #�-"�"Tp��ޕ���v�v��O�dj�L��c@�O��$�O��4�.s
���`�5,�.UwԔ)�((W�*YK�C�m��H��A�u�,b>�+N�H��ŕgZ���գX�酉W�3	ֈ���Q_p��� �Â^�8�>��I��PW�4�,��T?`�Y�D�����c�I�)�3�D�Yt(kD'-2��hc��?�!�ؐ+���@1��]�9�$͇?��I��HO>���L��-X�� ��`�Y�-ҖY$vy��$�ɟl�Iȟ,��,�u��'4��q�D�W|�!3 �
l�8!f�J��Mc���>(&�؆��8���Q񢘇]L,�C�l��A��Й��&j��棎$#��(��i�H���I�&��@�L`���A��=�,mB�@�OLalڤ�M����Of��(���; ��2�#�z�<��ԧ$D�hPD��3�F\�b��U(E�0�I	����<��KT�U�f�'\b L ;YLT3$�<��avA�@_��'�bp�#�'�3���c0*�^Oܸ����a�R�)�ޥ(�,�U�'�l}+��N����jچ��䙱	�Y��Q������"�=-�� ���C!w��'��ɰtC`m���M�vfX�p��*���I���I}�S�O,
���SH��y�mC~o`q�	�'��7�>ޅX�/�e'> *�n�$�<�*�"��f�'�2R>1����şd`� ��QR��B'���I�ğ(�I�2t��S��]'<���i&	�?�O���,[��sw�(/�iS䕢wH^�'�@��ţr�М��)A��>��D]���,�%)2!����(}�R>�?aR�|��d��8]r�e�P�l��jUo[�yR�^���!6N���!�ʎ��0<�1�ɰ"��0r��n�e�U�Aipsٴ�?���?)�hبY�p���?����?ͻ'��\�R
���yg$Ȧ�"tx�*¥Ҝi �W�Gf\P�Q����'w
\�c�MH�<aT��bi�1f�
7�����&uդ���Z�-��س@�u�e�}"c����I'f�ly�rJK�@Zu�-	�����	�T�<�i>%�����O�H���/
Q��"A�O-y�-Y(U�Q��xE��'Gve�&�3%3)�cM�lv�HA�O�y�'�f����|:Uh[��@Gf��'�(Y;�9F{�w���?Q��?��	��O�Dt>������\ؒr/�kL���cM��m�\���7��>9�$�> ��igld���*�����H8+�a}��G�?���P�,Lw1�E�Էg�@��iޛf� ��O���+�I�=T�X���{ �@����2I��B�I.h"@�uC]*9��츃K8e�b��C�O�˓,�~� ��i��'�j��ݷ=)��1
�5������'�R���e�"�'��I�qT9��)�B��
�8�9;e$O��!�V/1� �!cd
�t�����h�ٲ���6�1JD�'t����M�%
Ҧ��R�m����s�Y�H���3+TS�J����S≟Y�f���o@���>.�"C�ɾ9! V(�'v�:x2sC�@UZ"<���4�0nZ*[]������(�T��Q�t�&��5�S9�M��?y-�����o�O��Rca�"F}�IVO �+X���s�OV�d�S��6m�� V��e�Ƙw�"ȓ�ڟ��'j�r����Z��KucʎDl�O¡�Լi���
�N~8K��xyJ���*��a��u�K���1U��Џ\�"�.}�u�(}2!��?��|���k�Q!
�#�쟺]<x�3a�
�y��+����^�}:`�F.�0<���	�z>��2@�I�k)L��t���U(�i��4�?a���?�b�H?N�0���?���?�;w\�qe��*V��rB�O*XHT ����gh�)�G�1s>l�F����O�'�ԑ�0G�!��Qr��.]�Ρ���1)�e3�U�uTlKe�P�YbK?9ن��""���F1��S�%Ȃ<���0$ؾ o�/��$G!Y��O����ҜsU(@�0�U�6o�4�d�Y�p	!�8SJ�A���k����L��	��HO��O�6�U S�Hgd%L�F�j�cK�,�6�y��?!��?!C���D�O��ӽjg�!�ĄU������ȝ�R�L���1�<���b��1��*�w�L���i�N�fC�ɞ`���ۡMՠg��p�)ŔT�L�Z`��O�	��)� �y�ĢS�r%B$��f�����7"OD���`�
#���Ie��w�������^^�u?p(����l���У�Q��%���s�$Ub�C����I�X<����ǟ��'r�E��x�	U�`�#�(ב��͒��R�%w��d�j#�O��X��J/�HDD�A6cqB4Z�'�`H�؉'�nqc �Ɓ'fn���6Jx�I�'�lE؅��x��P��3.���R�'|�6M�]��qBg�*24YJ��I�1O�q�'DȦ��IȟȖO�=#��'{�k ��0�!ID3�h���'�B։"$��T>�r�^�	��hH�"�br�\�O�u���)��#}"R1sց́o���Y&h^���'�d����ɧ�Oƶ,1�2A�"lk�,a�����'�D=����;H�CCM a�A Óq���Ҷb��_͒��mx�\�Z�����d�O��d�K`d�8�k�O��O��4��2堇�=9��I��ڀ?���Ɔ�3CZ�8���M����H����|&��SW+7U:Lc�+b�&����� F�J���/?țv�Z��(�3��"h_��r���4<��ۓl�)0+`n�����d�O����dο:e��V�)-�.�P:!�$�A�tc��cȈmuE���ɤ�HO��'��3�Z�]�D\ix��^%Z�m��Ʈ'g����ɟ���R\w{��'G��-�D-��띶:���d�źq�����M�
Y����o7��"���+w����oJ4��7�I0A��9K�&<|O�D�ǡW֊�@��'����5�׿?P҄(�O�1V",n����a��a�2�6"OF�� 7x=�,@%�S($�Ȥ�d�W�-, �	��?��6+�ɺN�7IE2PQ�>!݄�����?q`�N�?y��?� j߫5�dq��
g~",��5�,Ӥ P�`w�X�p<�ĦE�\�N���$ѥZvɳ��ƉR���RIH8������ON~��I�IB��d�On|�'A����Rqz�h�AU�:ȩ�'R�'�O����O���Ob��,�3L��%�e����H�O�}m� U=.	�	�	k�+�O�H�J�4��d[P�|n����]�g�T���� ~���lR�I�tI��d�L���'ۨ	���'K1O�3?��jL�*[B)�5d٣%��]Xī�d�� �q/��?��F�#����F��8ajl��i.}���?yg�|���%��br�@����2��U�DX��yb쑇&j^� �	�'��C���0<��0z����/X�/�v��0��C�� �ߴ�?I���?�A�\1j)R���?A��?ͻE�� P!�cHpKή0�z�Q�yr�õ��<����6z !��
SQ�9�0�ܓU�DɅ�	�M�4�E-\����5e�&��<ф����>�O:萍�<m�F�O�k��i�"ObE����6��T.�3�Bc���ى��ӟL�\�3@�B lʚew�C5%�tՐ��5a�2 ������Iɟ�;Xw��'���f'�}@@��*�(؅/�[\<��4Op�!S�H�=��p��,_�	q�����Q�6�!�H�=�B6�#�v(�"j�W�h1�u�'���N�(n.L�K�&Y������ybgB��֑hcS�+��Ct/���'�^b�@�3O5�M����?��L�Yj��V�R�*/�%s����?�mZ? �0x�	ɟ�ͧ��d��W�	���s��/D9�b"%"����pt�O�5� �a^>D�4+6�D)�a�'G�y�����'��a�.�+/������[C0�+	�'���� N"PG����I��[\j���'rz6�!�	P���r ���6l��*1O����J�O��$�OHʧk�r��x!6�9��]/��(u�ݷ1������?	1N�`���ǃ"DI�08Ҡ�'���@����<x�~�j���̕��\8���'O  rH%F������j9�@��%$��ʧ	����lO�@�(-)�B�#Hv��O�YZ��'��6-c�SU�%wd`y�BM�mf��\)��?����䓫�'r�8(�,M�q/����*�x�AK�e���'��'�"�Pt#I�c(�3 �N�ƅ� 6� 7-�OB���O�0q'��)�t��O����O*���͸��TD�Pְ
��n�"c��k$��UX�L�6ʧs��)I�!ȡ<H���4�g>M��I�;Ü�Ë��q ��o̰>�e�IP~ߘ�?�}��՟����/H b3O$HdX��ȝ/�4a��S�? �	P�!_

�<��b��QB�đF���ێ��?%�'��)Ku�����Z�T (���߲B�Pءq�'n��'1b�}�1�	ٟ��'\���K���:Ή�c���v bȳ��d<q5�.q0��`,�L@��Y�d�p���r4�a��" LQk0��1Y�T��U�
��
�]\�+pHW^�A%'ίVҝ��1p�2o"~�����S,(�hH�<y����)b��l�֟T���F]s`#���lh�s��C1^���񟨐�nGԟ��	�|J���ӟ@%�L�uO)c��n�C��}���$O�0�D�3����R�``�S �v��x2��?�?qO>)��Ҍ[��ɧ�(5Y||�t�<�SNGO.�3h�9o7L$�#hh<!��i��@�&���ty�D�6Ņ>f�j�y���9g6��O@�ĥ|�Ҭ��?�r�S$<�3�H0�h�2�[�?��2dT�R�����򙟐b�M��p���0:s� }B��,�O�1f�	�����?���r��>�sb�ܟ��S�'Cm�=̟�LA���W��'u�l4��5��|!c����(l#�O��'gT��ɦ�HOP��5c�0؍�E,$]d�u�c�E��I�4�Ɋ|�Q���G����IΟ��i�5S7������W��h .s̓$�ZQ��	V_��U	��<�N�"��ձ,�l��l4<Ort�����N��E���:d�����d W�	;f�����|r�� �m�Σ,�������y�I���
	)��U|r|��
�3��T���
���,�>���?���@�ǀBq:H�1��O����O\�$T������?��O@�y�s�H.h�"`�� o]��
�d�
�����5e_2ܒi� y�XwKL�P�D9��'56�2�	!��T*dDա��2�@��?����䓌?)����'nL����\���3E�6[Np�'.D��&� x2���>l� b���OP�\�^L0��i���'���!%�g.�p�$�
@�4�(g�'B"�T�1@��'���Qv�|b�H�9�`�Z�g�.��q
ӭ���p<���F��3�L�0�vٶ���/�����	�9R���S~�I5u�Y�3���q(X\0񬊌N��C�I�#ub$knE�_�>sOI{\�C��<�M��-�
)�p5HՇO�-�qƁ�w̓ ���yֱis��'��h������P��H�b޶�"w���!X��	ݟ�i���|�<���dF�r
��W�vH�5Å��r��9�H�Fx��4��!s�,� ��P'Q���I;c5����O֓���T����K"Q�*e��=X"pC���O��C�JKR ���/x�N���@9*%axb�?ғS���r�,��%* �_>%"�:!�iQ�'Rbo��y,a��'R�'�b�w ����ʏ8AZ��s� >-褰�d�%2I�y"�=w�LT��@L�4��qC(ָ'�,�	�,RL��'$ϸ&^.H�cO�
�\1J1�|��O��?�}&�����G2y�ni����{�FM:D���!ʑ	�d�����U5>�9��4?�B�)�'�x(#֠�+�ԡ�"m���I�% ~�����?����?ư�x���O4�S{��[#�מG�ִCe�C:N0*��2�"�I�W;�i�"�G3IY��ktmʱl7,C�IU;>�ٓ�ūpj� `��*
�t��Ub�Or����12��X!6F+���t�ɠ��C䉓nw�z@�ׂ~�޵�1)]�'�@c�HR�}"(�t��7��O��������?1�L����@�,�����O��sPN�O�df>]���$�� &����&b�<�d��U�*%A�'/O.u�3&��KѶO�кF�8z������e�0��'�������?�-O��˥
��4����J�<s�h6O��d�O��"|J���/T~�u��V�?�<�:6GL<�D�i;D��*M6�0uZ�GYVb��қ'���7��	ڴ�?y���ɟkwl��D� մ��D�͔�����IWPT�D�O�x�	A�>�6��K���%��|�-�P�ꗣ�U�z!�MW��5�p�>a�����e�Dƈ6^��L��j��q�~)K%/S�!�֍qcJ��Zop�{�>��T�P�ߴI˛��'��:y��F-��`x��a�H���$�O���۞}<��S�3���j�E�"axb�"�S�? D���e3|���ǅ�
?`�*U��ަ�	֟��ɓ:Ԑ�i����	�|�	�ߕRc�@�*o���cF�lv�ę0��2f����P�h�P�QuHc>�O�q��.�2k����nM0��CD����ʪO���O�����Q�θ!!��M�L�Ԉ�-R��Q���đ�[6�����?q��l��,�@B�7���#EH�!��Y�'�0ٲR�Ef\�|��� >4�OF�FzʟJ�SQ$�q� � ;�ѩ'��:]���M+��� ���?Q��?Q����d�O��S )�x'��>Yw��P/+��"F�@�Tu��C8;�m��w�f���Ș'~�訖��=�Bp�ڊ}�Rqqc���\�,ԅ�	���Q�@�`�FusP�G=���)tc�O`���I�]���A���  ����V � C�	�3���(�	պd����7�T'
�$b�T�}�	-6��O��d��s+&T�u���Lp�#�
]���d�Od}�d�O^�da>I����Od�OzL���#�.�v͊h^<���'�P�����1!\6�͚�?s�ܚ�B���p<�cX���&���72���Bc��[�:�J��&D�8�b�ҕ �FGų+$U8%�9��jݴ"��*өU�O��آ(Ω)��Dy"�iGR�'��ɓ:$H ���n�8\;�K��hz��")��������c*ʹ<݊$&������&&P�y׎а��'�V9��ȤO.%�s	�� :� 2m�2D48�.6��,J��JK!5�9h�*O)#�P�'h�#��:A��`�d��3�	韞m�dA�%<xk5����~���IM���'�: �g�W|b���L;�P݇�ɂ���<q��䙻$�j�ae`{����'�}2��ch\��ׂĹ`��E�����y�
�Z�D�Ue�F��9�v��y��Z+A���ȵIvB�h��͍�y�H�Z����Ӈwy���o��y� �"Q���"MF>f�9fa��y��Դ ����BR���E*S�y���� ���o�Q犤+ң���yRj��sx,)b���>	L�.��y�	�\��9��	)2Z�<���&�yRNA����@�PZU�X�~~�tB�'��c���V�e�(�x�Y��'7,�
�GA�@՘U��qM�<�'�H0T�I���0k�%ܔe���'b.�Q��!ij����SO�1�'(�	r��]$F�X ��KªM��c�'��`�NB8��r递9�*��'F�CVO��Ua,��R��]�n���'����4g��!2F��$O���'m�=;�˰#8����ۨG�����'�,���4ut��(abM
���	�'����4T��s�n�7
N�8
�'��qM�8~��W�J5{D�![	�'�z\���	3�,���<nZ���'[����۪wW���$�_�\,��'`�C ���@@��X ���$u��'{��5�T4d@|yТH���٩�'��"�B�y��S�#�y�Y��'J��d�4a"TD�N]*p����'I�1R��5~�!�`��:vɺN��A�ɸ�ȸ��)���-z�v�' XD�W�O�4D.8��D ����@�XEP3`��B8PţI�=l��1Ɖj ���"Wȏ�D5���~�<Y�-["0:���g�� I�|��d��)n�%U����O${���,�L�j]�ӈܐuR�e�4ώdG����I6p�G᜞�P�1���N�}����gn5}�&�7�2uE��(_z.5y�'�pL�劓�l�Zm�+^��qT"O���U��:7�J	Htg�$a��z�"�^}RBQ�C4)�5�չI���ɟ�I�cщ7��W9v����nǯr\��s�KF!��G_��������T��DW�X�h�b�ۙ�y�;OtD�ф�#l^���d� �S��X�p�׺)��|�ukE
	:� �#�>O�LKa�Ï�Bi���O>}��]�|�L�kc�A�>\2���J��$��E�r���S�? ,M2�� �X�ӥ Ӭ.'^Pz���X�C��^��p �>A�Y��8�鰟��o��\?�� ڭW�<t@T�5D��Q�P&`���@��tm�J�<1�
d �e �O�^�����i��@�&���\�rI:e���)+�!�#F�=	�!��L�2�f�Y�e��Z�H� ڒ�JP����c�iI�"M�Y�����N5ʓ/�Uk�*q����A��$����I6�P�� �,F�1"%l�7LK�P��k�	r�~��ף���i�(	�i:��"��:�����PΊ��VKL5R$B���"�=���*$H�3�T$H�zA��I�Pj�Oj�9%ih��o��gҔ��NFv�<B�	�=nhӇ]%����*ԟbA,��g��v��T��� �0jAcE�E�y̻�����(P�?�.yK��ɀkX(1���D�����@�B8��kS���$-��� (`yr�]�&ʒ���4 8�:��,z�h���,$�6 ����V�H�G)Of 3�	Q4�,��VN���4��ǡ���4����;X�4!FF\�)�:HU@Q�o�~��!�'��4ysI�.���YU �*1�<B�Ob�����}�r�;�*˽f�.Hbԝ|2��\q�/G�Jd�b�[�j<4K2"O4dPQ�W* LJx���S2�Nx�aIR$Q�x"=i�+ f�<���!	-�<��w�sw��*�|,#"�Z �� ��iU:a�Dظq0`��&�җ$�<J�|h9pJ����DN� r(���	E78�e��!9�"<I���!b��g\'J�┰�/�c�'6�${�.��w�����
p�+�O����[!(���#B�v�y1s�̞  N���éK3a|Bgͬ{��	ab-VE���h�-��͸Sd�0fVb�R���?<�X���eV��4��A�*Ú��k�@ؑ>��=��ݤt�мȌ�i��j3���sΙ�Nx<��a&O�9����8�u'�_�3N�r���M�0�:�w����Pd�&��}K!戵@�dt��4Z���s��͜/��ӧ�'qǬ"�W��W]NtSn>&�t���L�F�R�E�5�&�a�G��{K�0h ��1�^UY��d����Q�NկBX��*��$y.���5*~�f�D�n �q5N/I��/��p/Of�Y�$v`t8�+x}�k�b�ua@`Nס��O��kt���s2��8���`" � �|a��X��'�P1��dЇw�<!��T "�P���Q�'�&[�̴ʷ�[�|�����@�'�����,�Z���`d�C����g����~�{B���<1`$�<=��yiD�G�gd8�dl!�'5!�9+'�Pe�@I�cdT�`��xlZ'edh�)��S��Ms�ń �t`@���x��� ��=�L	ФAT�8�C�J/ ����O
U��˭!�> !�ը|FV���	9T(F����'���CbU��ӣOC���&`�H����w�t1&M� l�` R���*Ѐ��)b�c=���I���53�(x�dJ9*�d\�D�O�|s���P{"��`b���U�t�=Q6�u�i_� 2ܡ����)x4,X��FEqO�x���b{���N��eɪ|JH޾x����O�� c&mc0�F�tM��Gl)��X
0b�t�-1�yH�j�F�j�J��؎8DVQk LZ��Ʃ�J��.9F����F@�D�E`�!��k�OZ�S�xD[�F؞N�ƈ�d��?��F�������؃!-�IƂ#}⏜�C�J���'<Xb�j�돒~����ҨU��pr���H�+c��O,�Xa�AGZy0#�ݫv�����j̧6>��Ã�HZ��B�����à�[��舠�ƺ+�n��|B�1�=�O���>�bDa(A&%4�Ɋ�O@�E��\Q�)N6��dS@���Hy�tZv�q�bD#� Pa<qOk@�{��y�1	�2C�=:��G�i'�c�<8��W�-��4��`��Y���+7�l�t�r�J�Dv�aQ(�9Il|�*�U��9c��2�"���ʟ����Hc�'�\�h���9[�|�kA��w��'k�s���q�m����8s&�=:&�y�X;']�H��/r���g�m �r�a	�+��x�F�kr��X�[����Uś�y_�x7���Ss��qE��B� �g≷~T����#W�Nk*ŪaE�
9���F-s�%�6�Z�:��!Ň�^l��0#V�Jc:���Eh�I��o�1�`��b���{t/�!�$Drӧ�N�,�*���w�I�}�O�0А�\�*�����<~D�3�i���<�+�[ \0x���C)sنl8�˛�B!<���|�D��>�#&�Af��[DN�f�� G��~�c��"C��:b��X�n[�AL�j��q��롂�!�&�����:T��fD�#g��a�K+����G��O����!y�D�n�U$.�*���uRXIQ�)׵u�B��0gU�u�ڌ���6!b}�'D	�y���:��HR�%υ;�6c�OʬS�G�q�j�!#�X*s%~9�����I��?q��N�6��5�N-w�D�t�l�-mLt��	J�X�$�"��r���F�I��0��wH�=R>�u�'DT�E	K�\�4��B�M��G�*`�p��K�Z��Q�j|�z%�&F,'/��*��O���'�ĦEq� MBF��z0C�4):���e,����a.O$��'��t������'�z1�BEȊ*v�c h$ך胵a�n�dW���1i�oܔ�.�f�a`�<��i�K��#t-A	r/�T(��<Wॡ��\b���!�&A�2�O�%�	)8���IGk�ZD.$+��u0U1�i-W6�XS�þf�`Xr�B7'�v�vmC��y��'S��T2�e<M��O�`a�T���|c�5S1"%℞>�"�'&bEH��7l,���s����*���#��r2���|0F�Γd7���`n�>[�,�?�edC��?Y�J��G�e��N
 ��i�r��>���cslL� ��6ƌ&�O��I�9��\�C�ɺ�r$PƮ���ɡՎ@�~���w�	�F�=�'��s&W"%l� �ā ��h���KgD{�Q5�D>;p�S1�^<H�^���ٞ4�1O�=hQ�L�O����˚wR4��$�'�(s'�[n�ijgA��G�j�j��ѬO}��:eȈ<��4S����&����O�����:LOꍪg#��Ma�-I�
Q�
����|�=!
���Έ:��NͲ�'#h�Y��2.��5�
ҐF>�	�'�V����,"I�|Z�VPHx��cU0;��� ��܇!h��=�O~���43��#s�I� sR�$��0}�<�0Q��K�'�d����'�?1
�I��P�So�0����_̓��1����?K��1���d?���?�ɭ���Ʋ6�	x������֒v>z��	.V��x�!	�,ϖ��"I
�]GJѨ�
r�����dَn�!�q,ЀT���~>���{g��ۗh�6,�XJ�V� �l�O�YH�F�@'l!�s�˜=	6l�&��0������|�~:���7|Lp �A�?��"~n�!�� zE�gu6
e�����fc�$L�sRoS���O̵��4YJ|�1���_"������Ak>���G׸'��A�'�D�����>^	X/O����kČ%��*����RhD��HO�<JWG�&N���鉎y�8���Ȃ>��]b���y��3���HO�N��E�"Թ���gr��]�Xv�p �j	
M������x�7��7JB�ũ�d��)�S''��8#��kM���j��4�"�ۢh8J�J��k�M �Qp�0!�҃	8���F�,�Ɂ��pj�ώ��4��E� X���V���
��\�8���T�a?yPgF�tf
�CP�@}���_�>��g�,a�|KT��u�������=V.���ɗ ����	[�� Q�Ad�,��`iO���҆�!�򤒅}e	F@.�hO��X`܈�T��D��8��0�d#=Q��*LN-�FT��: ��'pJ�I[5/|����! ZS"�X!�T��/�L�'�z�{r ЧA��J�*F�3σ8����F��a���%e���;���2]8�`*m�tH��\8��'t���#TA<!�W�@�9���;��ܷ&�N��O8 Cs���/���"�dJ�3�����(�@� ���-���4߻a���PYu(��7I�E�'���	�^l2�i��09��)����"��QbT��Cv���)�3��)�]>~�=�dm���;���%�g�/?�s�9}�d��9�tAz�'pRhp����  >��r�kX�6:��i��`�'��ȗS?i��\�&�̓!�8��œ'�e�5�Λ��ɗ'Ϟ<��AǴ�M�L�Gx���s~2��a��9�DH�2c�-[�}�b �f���<5Nϒex.�I�}  o�<Ѵ'Cl~�,̫iQ����+�9�t��P�?+ؖe͍J���Г�<��)�����#�.��'��8(�MP�7� e��.ߚ~E�L�ag��r\�{/O�s6���1I<����eA�ndT5
��L�IfH�q�^�<��ND�t�U����z�'�N��eڢ��lʱ&�-�]a��є��A:u��F~|��'�.��޴B[J���՛�%m��i�N,)%h�>�R0��k�Q�\�"g��)N-+!`	���9�hD]yb�J*��t��L'<\�2�i]�'�x�a
��-U�}��X�
_���'��_7;�:Q�U�.vjDH�
�k�����6U��`�N��t
�Ѹ�G>/�@i�?��O��㔯�#4�"���+�=#��>j�
*S2�ؑ��'��p������Z�y�ӊ8������	Y��W�kQ>��˓��'ql������"8����/�[�na���O|4�5E��:)~����$�n`����?/�8$SO�nH�(��M��B���*�	2{ʤt�쓦B �С ]�k.J�s�O�D%a��G�L�Ex�	wW\��#��]v�HƦ$���O?l+n"�I�g$�,�p�A�,��'��-�t�Q�LZ�����R�xs�{B��;oZN�bk@��:��'A�"TH���D�j6�ؕ��;`�uG|R<O���X�ex�ʉC6��׉�<�޹�a�M�W)��2ד8���ra��6�n�*W��&]��\� /����H�6J��Gr��C�E �v �<��'�0����P�vT���
���sa.l�T1!CdA��?��C�/����ti,7T0#GlQ���Ѫ��`�y���M�;T�qk�ȓ4�Ox�"	�HA��T���Z��	%�(��X�#�~�g�\�46v��F�<�����2����5Ǔ:��=+����?c�<���7Sl ]aN��[ǊTҳ҃^�,|1��5`��q���y���dA*�s��*�́9�bϣo.�K��'� ����'�k��V�/��u	4#_�d�X-'�qO��Hk�,9��˛8�LA�$�*~�HI �g��y���J����4�@`[�������=��'��If��²dO���Ǧj�����3K\28Ѹ��B]����T�׆*=\� fU�V��u� -U���qg\������h� ���#.I���?�0js�,��9Ack�X�0��"T�t����R�� �@x�Cr"O�Y�D)PШY� ż/�r�A"O�:R�HȢ�x`�1	�.� 5"O\QIs!�aj��t�F�_����'"O�l��ٱkZ�}���T8}�فu"O� <���O�A�6`7$V(����"OR�A�ؑW˒��w#��I��k�"Oܼ	��ͥF&����d�so*�IC"O�8"���C���dš1yL��d"O�LB��e!�4���K��Z<�W"Ohm*�Ŝ
5�U�hn���"O��"!�b��$*��TT��Zd"O����ȇN�Nu!G�p7Ri��"O�dA�CV�]��88r��/`��"O|� �k��a>~��F��,�a"O
��MM������P����V"O����WMhq�B�zh�ȃ4"O�P  �ɝ' ��z�-E (V|Q�"OxE9�E/v�I$m܋D&�sc"O�i� V�'6���7�y�|�b"O��b'���5����`�,u�<=�"O�$I��(YW��E�ų<L���"O�%ʅ��`LU�-� 2#\�"O�E�AGڋ����vJ�+��3v"O��,��?L�`e#U�B/��(7"O����IM$&q�t�K�QI�S�"Ov�	��M� ��bN.?@��c"Od(��*|L�P���	6:��"O.�;�#�n��Maw.�ތ�F"O`���ϙpEbpYE�X�g��-�"OP�ȥ�)[C03���<��c"O��抗J��*$�*Q�Z�Qs"O�hv���'%n`�0���I���J�i`�G=0��	S��=�&��ȓJ|H�UB��3�PI��E	Oh ��O(t��n�6�����?A�=�ȓ1ׂ���+�+*p�h���;0�v$��#�����8Vlb�`��к~�J���I�"{�m��GT?4c��O�<i�C��L#~�9�G̼��ӌ�G�<�T7��4@"�;|\�i��D�<!�� j�Z�R���31���2mJV�<q6�:D��R�f�5Av���'��U�<�w��T��陴*T��(Q&�N�<1v�"'j�9�Ffװe���Hw�`�<�g�Y�A�z���߫k�T�v��^�<y�'J�?wj)𮒍gǖ�!aJ�P�<	�ʌ�wހ�p�H�>��P1⢃C�<y�`�V�8���#+88���~�<ď��*̊��Ʌ9x�� �ŉD�<5f�\:ȹ�k�:F�ai�<��QMV�R�̟u؁�p@�^�<���Z�k�4�( �)���V�<ɢ*�+F�V�bFk�wn6�:���^�<IO�4b����'��;e�pUu�<�wk@|\Y�7k�&6z�����F�<��)ʵBzN�h�ț&'@��A�o�A�<!t�J:;�l��nҪM��hi��}�<�7������/hX���e�<i�H�68n�ȡ.F#p2!cd�<Q�F̞J�:4 Sd�W�;� c�<Y��T� ��KۙF�����ȟ_�<ysg��p�H� d���X��^�<�C#ٔH�f���$���B� [�<I��:����eR��j��p�<��c�&����C�2>�V�;�em�<-��ҥ�B�b�~��sA^3�����O����[�Q|�J��bk:��ȓ<H�d�/�n�@�"TO&�p��S�? v�#��:���Yo�T�F͹�"O������4��%��(@,���n6ғ�h��d�=�V��d�<2�`��'+�!��)I�R|�1��|��@�O�4Hx!�V6,�)ƊM�(����G�a{��䀝f5~�ۻvՂ��d��)!�#O4�����D6-��C���I�!�$I�E�*P���Y	1:���R>b|!�DD<T�m��Y�w9䜰T�ظ8
�gh�'"#}
�'4��$8re��I��K3���yb �14+��	�H;Ҏ�qό=��xX��BV�Lp��zc�.#�x�ɳ�8D��@`'�w�(���	��jV$���6D�H��/�:m��l��Dן��qhs# D���bه�`!�f%��R*����:D�"�D��H�<DP뇯(�|���`9D���c�:��r4%��~`Z��8D�`��#�>�y(g-
8R�ޑ��F�<Y�&2�O(죢!�5�ĹH䊣#1���f�	n>����
=��8E.�6z�&D�%K8D��'�ɲ/28�d�ص	�2i��g#ړ:Q�?�(��'t�F�X']a`���-D���4lHv�4���L�_�60b`j�h����T�BdB� kW�}�(F|9�B��
99,"�,N�.*�x L�9[6B�?�@T�1��"�f�x��(��#<���?!a�`׸'�v�@� Xf�KL F�!�D�*��X¡a<"��h�w�R!�$�=�~�É�$�� CPc9-!���KM\��@<i�RP{��4\qO���Č`t8�+�O�O�:���ݽy$!��D�i͖�#!-�L����El9|!�؁v��1��!E%��sAŸ2�!�J/���8G�;c~Y�vd!��1 �D�p��	W�����Z-!�����eӉ.��-Zr�-?!�K�41��	I� Pa�BкH�qO`����
�,p��!r� ��U#$�!򄎎Q��X��K�r�x�Pf�z�!�]�E�Ƅ�ᡒ9l��PpA��b�!��h�1w+ 	���Cna�!�[�b%l��䭉�H��웥o�E��	m��(�N�x��p�v�K�T/�&��"O@�DB�Ī��3�	�;r��"O�ۦ�bW�<��Lɍ^��x�"O4U���U�|���O8LS^�õ"O�`t��+UL��dJæ�A�V"O$m��/�|&�He��18��9G"O���&?*E
����AJ���"O!SqB�HM�m��Ú�5�����0�S�'-j�a:���*9�"i:g�%:�8���'$Yp��,2�H�!!��t��u�~\���^�gFm+c�K$��ԇ�c�FZ\�i���k��[�%�D���"�� �B�L�]��$�fY6g�n��Z��)��^�>ܞP�u�S1[5�}�ȓU��}��#^�9�Z���NThm�ȓ[!�M�r�Ϳ3	��scUF�oZ��E{����9�N��aA�p������ ��(�牁PH�5#׭R�l?꼘P��U'B�ɒ)�ܢ� �1%	ͩS+W�Y�C�ɠM�� uぼ[��Кt�������d7��+� QsաQ�%	�0�#�
'FL��b"�E����ǀ��G팰Mi�8��S�? �u�Q���.+�����E�<A��Y�Ԅ��9U��}�dF1Otp�6H�u0C�I�M`�8(A(I�^��E�V�3;��B�I�z�*��Ў�M鴔�D�++�B䉓bJ�E�`I�  �� �B�I����"6��I��;��)D�vB��$>�VQaRD��<Ѐ<	ѣL��C�4�0i�v���S�B�D$1DpC�ɨu���3���/V����Jr�R���� ko��y�BQ�ƨ�p�6K�C�I)�B|[���!3i^Yr4%��^Զc�|�뉫1�l��fW����e�&tu��>a��iB0u��0��<�b�D���=W�
O�ݳ��P�^N.-"�mC��ၴ"O���6䉣B��� ��R$�K���y���4wѺL�°SJ��Su ���p?a�O�
W��1MU��3��72��� 1"O�ţq-ԐH�H��-�4_h�I��'�ў��_*]TL����}�ƌ���6D��T�r)ʀ�2G�b�hx`:D�
�g��S�8���H7O�����$.D�J$�
��b�(���L��S��0?A���=�"�	�W �S!e�6�L\�5Ñ\�<�e�J�jb0s�hؖ.Ȃ�jՅ[D�<q�ɚ�;�0�"�.���z��u�<����G����Ď�v�L`Z�i\�<y��S�(}F%��S{�����Ar쓁hO�O1>���ĖL��Q��2����'70���݀ubYx��ALT9��'�#=E���R/�Bx9�`%�|��ō��yBV����YI��EX�J��yρ�����%�<jE��-��y2a� 36����H̕
JV�+f�)�y�FH�|�{��Q����UfЍ�yB��br����B�uG2�:���.�y��.O�䊁"��v�Q�����yR�ҽ1����m� 2)]��y��`{,dc���f ���2�y��(߰��fF4c�`�B6O��y҂n����1�Ć[��ex���7�yFܔ� ��
� ��A)�(S��yrƛ:_7 ���eә��t�$�	���/�S�tOG�g.�	>ux��tl����cE�C�"v�H rb7h�T����ߍ~2&�8��8��?�+F���[�v°�X�i��-�f&"D���G�7 `"�ʎ6��Bg"D���)ӡ_&�PyC-�H����3|O��N<�e�3y���cGӆ*)�(䡑�<Y�k�c��;�b��xJ�L�R�5,�25xFi.D�T���Z��4��C�p���j��*D� ���,5�\(u3I�����(D�t#!#�,W�8�QA֌J�r<�1'�O��'���C�
&.+ְ����b��ݴ�Px�� _��)�"G�Ta���y�I=U���i�A�'�iړ�3�yB#��>0�3�3g�RX�s���0<	���	74 �9�Q�2f���t��q"!�$ѫ�|��g�;3y�<����6O!������'�8�Zf'ِO�!���ԉ�L�V�� ����!�D�pV��:RjZ	�s&�G�!�E��밬J&#�@���ʰX-!�du̔Ɂ�`�=I�8�����G!���k��xx�Kh�M��R�?!�� ���N 3��	ДV�.u$��D"O, т�<A��L[&M
:�� �"O�0愛!V��1��A2����"OX��B^2D�-��W�9����"O����&��<��Հ��^S��s�"OP�bg�U��厾V�N�R�"On��c�4��!�홠ߠ���"O �;�K�3J Je�jF�$t�ի6"Ov	��	�EKV��+MF�"O�a!�10\$sA��>�D��"O�킔�#aBp�҆kňZ4�ո�"O��U�رwc�w�˞-��`��"O�!hc,ޝUHZe���d�c�"O|Ԫ��� 	��@��Ɵ3V���"OX�7�A}�R=I`�C/��#�"O>��'HM(~�� �3,c)�i1"OXE�p��H:�[q+�n���#�"O�dw�V_} H���P�.�X��"O*�9HR9DPb� #揱�J�Z�"O�8Kv���H{ ��0�|U�
�'�<X �(|d �@�Ёh�9P�'�X�z1뙍!�1��A�-Y�P<:�'5:E���-T��햃L�8,��'6Ĩ��~�<<h	�(D~u��' u�ʊ�!2�	�!ٸSHҸ��'���ĈA�h�N-�G'��FpE�'c�,S'�-���I�I�**��c�'_��AM�#^h�Q�M)��-�'�b��6�ߧ>��	�LC	���Y�'����G�E�dyj	W�P��'ؐa$�D��%�4��.�jA�'x5(��P���-�	�8BwșB�'{1:k��2�Ͳ�ŝc��y
�'MA���Q؊Da#��Z8f�	�'�H(����%m�����#U?Y1`� 
�'�xh�OM�<����U�F=z�d��'���B�C Y��U�nƍ\W�u��'�5�EQA*�[p�Ŀ[H<��'�*H�G��Fs����\�L ��j�'ʹA AE�
)D-���,�d���'�j��6-��+M@(Ck0$�ͻ�'�:�Y�kR�1���� ��H���'��2�ik�ڴС�X�/@4��'fx04��s��0KH���' l�R���}��!�N��T���'�<�����0LsDP�P��/�>U��',��0g�<2��S��t����'�8͠q`�!�08�IL6#�Z	Y	�'�r��q�"_C�(�A�p >���'b~#r�Y�*[�A��'�e�H�
�'C�pP�ς�.�v�j�Kl����'��P������qՌu���
�'���'MOI���dY�p	^\��'�,���C�<\��с�ES�ptj�r�'P�L#�BY�/�;k��c�'X¤�PD�&�J��r)H�d�L�'w�|�d 	����PJ� �2wU�<�P��R!����|5K��Y�<`,�az"嫠 Έr�Q�r��T�<0E�@�,0(�M�o��H� ��M�<Q�c�`d�AHͽY*�ӕ�E_�<#U�M�yʰ�͹Yf̓�LI\�<���J�X, hU͉�-�#��V�<1ҍ[�æ��G��$p 
�n�<� nHP�N8:�q�vm֨a�d�Q�"O�=$A�$�)j���R���` "O(��Wg*'Lh�'*J� e��2�'������C�^D"'�|����V�<I�IO/&�`Pk�aε&	��ҳ��T�<�'i�3���Yp��
Ƣأh&�C�	�?e4�Z�`Ѐjx�+"�m��B�ɳs��ܳ5��Fh�Q���4�B�ɉ�^�Ѧā2%P��Ԗ=�jB�ɊF�I�	Z�F/�!8#��&MY\B䉃K��}�p�Y?��yc�É�B�I:W�d��î�8��Q�N0v�C��SѮ��w� /P�BB�Z� C�P��cˑ�4��d��LY�B䉒#d�9Jb�ҋ+.i{��@9s��C�I�[��e�ₐ�PP�(	c/ۖ^BC��� ��D�?��JE�#,BB�	�
���i.O.6�B1;���f.B䉂oF��b��I9?n��t�Ή1�C�	���DJծJ��HT/N�/�C�ɴvF��`&�\2B�D���L�HB�I#Y��a�"��1��}�d���y�Q�k��<�%eͶ#s^��C!.�y�`�D���S_>qa�3�#���ybo�8[��pbt��/i#D*�oҨ�y�+\�e468S���	]D�|Rc�4�y�(�,KT*��f���較�慜�yc��b���2����F��ŧ���y�a�h*��Y�cN�.?"�9�'���yR�\���3���6e
Q�L��yҼ���a��"o�4����:>�2͆�=�b|�Hٚ<H�4�k۝�p1�ȓ.�,\H@�
�2)^��c�;K>��7�X$ w�Gcc a � ��'�F��ȓ��R �K.O�u���YLh8�ȓ+�@��b-os��ӄ��";����)�@V�T�Qw�%��HC�|�u�ȓ'~4�(@IN9��4���,�:��ȓ[nT3��5b��Q����8�,�ȓ�J�z&iD$onh���e�w�^��ȓ^����/@�`�V���`��ȓ-����0GϪ2="��f�XQ�l��7�j@E��ArA9�� X�T�ȓ-�ֽSRE]�\1����Z�j��-��
�hiCg٤T��U�_,�p@�ȓ����Dy�<3�B�<m�L��G�P��'��	҉S@��8)����@3�$#!a�;p�QcB�>oZЅȓh�>�1� 
z�����G�䕅ȓw��݋4(�'a���m���p�ȓ"�a��R�H���A��*[
t��})�X bT�vҜ�#��-�ȓ8,`=y��.A|J���
�݇����!��'�pZ 噅hHd �ȓ�nt8,�k&y;�o\|���d5�3ʌykn�9�ኼ|.�(���P�ai�xd���)6�䠄ȓ���B�@�sj"���:W,�E��=k�4�0LYs��tH ohl�ȓE�����N\����(�+��%�ȓ�©���d�h���/�=6ԨɆȓF���qH����YTA�ȓG�,Y���K4i���� F,����z�����y�Y�0o]=%�\���S�? ,����ڬr,�Պ�h	<y�\��a"O�	�w�ړi��\�狔/mh�j "Oj�f��jI��(M�n�`X"O�d�w�hPvPj%�3�ܭsR"OT8S3��F=*�C��>�ɂ�"O`-��ؾj����â[ ��T"O|�	7�\;�`E�V�(af4`U"O�t�0WS�ryʖ�T�>�x��"Of��6�=|?��"�B�6�� ��"O� IAɑ;PF}j��P 8�V��b"OS�eIo����� ��&��Ei�"O��wn�/p]j���9i���@"O���b
	j�*�s��/a�(�"OF�wf>)f�[�CA��I�"O���5�Q�D���i��Nj8��"Ot\���(c�����<B2��I'"OdlA� �7*MF�c���8�~�x�"O�x(2�"�QO��w<q��"O�)�U"B�2�l%r��Īgdj��w"O����*W>sz
Y� gP�h�ڬ[�"Oz��ЁZ�����KT�Bpk�"Oj���GPxP)H'�(Z�E"O>@����{�#w
W!(��"O ��E&@,m�hX�6J���&"Ol0Cb���Tc���&^���"OVHi�%�DFxa�H��)�،�4"OX(H1���2��%9�L�p�"O&�Z�ŷ8�|2�՟h�2p{'"O�(���l%0#��#��2�"O��bG�3^�b���!��z����@�<1��P�2������"���~�<Q0�>�(hy��)^ښ�P!�y�<!!C۵{�`�ĥY+��X0�!Sn�<чE��4��Ńf�J�K����b��f�<��Ť]��=)�J]�3���J���K�<!w/�q�0 BS큯 �p*䡓S�<i��^�N\j!�T�Ө#���q�Jz�<Q�,J�����@:&��Iw�E}�<��n�6R`6l[B��5"'R����@Q�<��ś�(i����킷\!���	
L�<y��D�:z�Y� )�1r3���IYE�<�`�M���$g�JQ�P�bWh�<	C��6@x�����1�_[�<A�I	"n()W�<i`V��#��U�<���_<�9ڄ�7��0�#JU�<����!�Ȁ��/ҡa�ˑV�<Qs�Y/Y´`�Ə�+�0��%ğN�<IuM+m}�\�f�'f;���&Lv�<A�B:p#^�y��V�f�\
��Y�<��U�?Uj!�d�ș|�h�RÃY�<�7�*vzY4$1�{�*�O�<����낵P-ζ�	�D[J�<ᗇ�0y�D����M+'s���eM�G�<IdT�[�A�V�(,i5 2J�C�<�Fȃ�*6h�e�<�&�Y�<�S������Zs�s�j�C�NW�<Q���@�)icoL� �ɀ��X^�<�GB���
�8φ<_�-�E��c�<1&�L8�	���¸Q#l�_�<� ��e���$�^�hu�'�PD�<�d����"��!�Fy4#�Z�<�PI~�d �4cդ.R8�4HW�<�.*Y�0+5,Z$�J�y�I�]�<	G/&��`	ڴIfV��#�[W�<� ~A(���:1�Ʃ�%NG%�ԍQ "O���&�3a�|{.�.��8ؐ"O����zTp�%MC�Y���QR"O&Y ����.�����DJ�a�"O"�H�+D���!U���~d�8i"O��2��ńx͞b�d�6W ��b"O�� 
�d]&R��c�"O�
�F]z��3�)XJl��'qP���@94KpD�p��N��� �'nBtk#�� �@���^�I���'�a@�D��n�`�'U.IA�Y��'w0!d��op<L9TM[�/�8Ѫ�'��4Cw��^pMI#A֊T��<��'Yh	���EDDEI��0568��'��p�M�P<��U��d�k�'v�aN�0m�Y�eg�Ǩuz�'�|��AJ��n�B0d �)�'���	A�)^�~9�dA�[3f��'BJ� @kM�qq������J�����'"4�T�/M9<eh�B͹FI�@+�'� �K�M�\��̢��*k����'S
d#Ta��*Z������_����'�Y��N�
S ���'�Q�6�
�'v�@���ʨv��Kf�]�]6�B
�'��� ��ʱ]��\R��8f"t�y	�' ��]�z)�e풹h�lib��J�<i��R�=�@	���3hz8��ZI�<���U"ـ!C��,>���pR�[�<� �"*��r�ֿ;���8��@Z�<	7�X�Ili���=H\
�hU�U`�<qTi��F���Tmٻ���BA�E�<�G�Z�'wT�v�¹j<�e�A�<Y���i��Q�A(�f�(����<yVaO�<�`� �8r4�9��{�<	�@��\pH�9A�1φ��+�P�<���$G+����eܨRs��"�GD�<Q�!�#����
�R�z�J��B�<1�F��uJ1`p�X�2��2��S�<�c�C�69VDk���cr"��pa�f�<���M.��0̙�->|D�!�Zd�<�e`D9|��E���ňZ�<��!c�V�<��fŕ|�d@��螬g��6��\�<�� S�.�~��*�"4�!h�N�W�<��	���l{ �� ��+%��S�<)F_�����$&ƙ!���mKI�<�E$'7`�:1�]A|R�ɴj_m�<9��V�d�ѷhƊ4�����}�<A��GT$n���Q�Zp��@
^z�<1��� �h6��W�4�K�y�<I��Eilap�/�NS8�Ѣ�r�<��E��|�|%� 
͑�	ӃE�l�<1�D�@���x�)�8]�f]���g�<Y�� �wW��LL7qB8X���Fj�<��	�#Ro�Z�Na��+!�l�<��̓.t��cw&�HH$��J�d�<��޽�йp�)ɨ5z4X���w�<	׍B�hǼ��⤈,"��h�vƊJ�<�6�*�T�i�L�%U�L]�Ƃ�M�<q�� �b]�A`��ɕ,8Dj0A�a�<�qIM�|j �Y���t��9Z*Wv�<��#H; mF��bK�6��Q��W�<��LƵZ)Q��9:�c���Q�<!��L�ب4j�}А3ԧ�M�<aȈ>|^������r�MO�<� �Qk�H_�a��yХB.�4Xc�"O��z0�T�>�����l��3�"O�)�q×�����T�*��\�"O���F�K�2�Des�m�t�-�"O�h��@/[�,��a��Ok&� "O4��'蟺"F���QG��=f����"O�܂�cV�R����t%��,�d1c"O�8��A�d|�heo"wmV���"O�hٶϜ+?\������"^��)�2"Oh���LR�:XL�G$۷�p�#"O����� <D� ʦ��-F�<8�"O��B�[.�`�q"�!Sf�UaB"O(�b���m��� Š\�&�v���"O��b)�nx蒂Mɼ�k�"O��-̈́*��ũ�O��j�>�"O"!yĝ8wKw�Ǭt�U�"O�y��m/v��Aق͞�=]��"O�͡%������eϰBF֭�T"O
TZ`E�N褛���|�֙�"O�%��� r֬�idI�]�vp��"O��(Q!��2��#�G��2X �3"O�rqM-A�e 2a-�L��"Od�3��op����{+.�Yg"O\�2�bܦ�F��M؃`>����"O�tE?�XyFMO%}D"O��Q�Y1fkl|���I�6�̘�"O��ps&��3�p �I���"O,�ҋ�}�,������xn,D�lkԈ�S;���2zq����$D� ��ՇTUS0�_,�h� (D�$��,[qan�3u
�!AR�����8D��hq'�,*�Y�����x�á�;D���U�40�&�)��,�hXS�b?D�8�lǙOg~�Sb鐾ep�t�>D�p{��K�)�l�������,p��:D��;tf�l,cA�ȓS��\�֪7D�L�`O0$ 4�`��qy�����5D�����,C�i�5��Z4q��!D�D#��G]��!�VZgD��p�!D����bЕ8t(d�sES�d�Xa�!D�P+窜'Bpި#�R'��a��=D� �T�T�` ���쐝W7��D=D���m��/�,J3�M+_��7�<D���oT� м᫶L�JL�"�&<D���2�^��P4��E?���Kf�8D�����}���h%���U���)��5D���F7y��p�Wn��VI��J4�'D�h�WK�}O���s��2	���P`&D�t�Ʀۛ~צ��A,kWf4��.D��(�D��#l�����*d	J8�k.D�hs��)|��H��+�'&��x a)+D���'hR R$Ѹ�	�g���Q�d(D�(y�aG��HiVI���NE��#,D� �B�r��bC��pNQCo=D�Hb$�P�\�$��21k8D����|������3���J��1D�p��螫 cjQѓ���7)��b��,D�@��ʛf�R�T@�(Jڠ����(D��sŁF�e�gFM'Z�1*r�%D����l�U��I�UA�.9Z8j�)D��)�.Bxt�TE�խx� 0��)D�d0�#��n�B�Ca�H0A�'D�H���֨]#����!U����F�$D���l��k;��K��^: 1��n$D�� �Z����G�"T���%mL�]W"O漳dA�4B��s�%T$̰A"O��Sq匊-E;A��L'0�Ȃ"O�qk4�K�ε�f+��ѡ"O����I�
��CD�&&��"Oɚ F�9�MC���J��u���)D��@q�Zw��x��Ƕ�ؙ��+D��r�1"���Z���ң$+D����%�'0�<���hUJd��'D��#Ss`��B��/�
��#D�(sun۴G$���㩔D�6h���"D� ���/5謴Jo���.��!D���ő�E�:�C���MT���L3D��2BhB��u�@(�y�R���H2D�$z늾�4���M,l�hlJ��;D�hxRE�>(�a��H��vdd���+D��3�J�'_A��{�I�jp�-	�)D��P�����Q�T$���)D�5�uo���'��b����w�%D��u琴Oh��`B6nTr���0D�����:#��5���C�l1* �-D�������f��86�^#rn���,D��񮗤yHr��F�t�yx�a'D�����5A���T˘��\3��(D�Xh�&N�v�R���OD�Yy�"&D��̞����/��(�ʜ�@#D��:S��8H�$b�",F���p�!D��0����d"$-"r��?�Ȕ A!D�@����@�	!�8~P�" D��Y(��5t`����vTH��3D�|�e�.���U'_3<r@6D�����JѬ���c��!�sB5D�웷.�/j�pb盎K
���$4D��@%�(.�F�h)�G��s&�'D�$��P4/�:��KC��V}�!D���Ug8.�BsCܶY�!;`�)D�đ6a� D�ܢ� �
 �j���o&D��)Ċ+`�\q��̒�X�z�H/D����fVK$:�{2��6/x�[��*D���C��XLd+%�5���8��(D�<y�ՊP�����"at$*��%D��1MզH�(-Q���$ :�;7�?D� ��)��(��!�R�[�O� �!�!"D�8y�喸tÖ���&Z�����l!D�,�F�I:Sv�qƈ;j��%�E/>D��C��8�[��J�y�W)D���bl�B{ƀrg�A�t`Ł�(D��9lC1�=#B�S&�5��)D���ݱ4۞��ĬQ*��2�'D��xF�&+6�8��ρ<�0��+D��QCA�e���Z5K,|8٠v�=D��P4�͕"��k�:`�Ѷ�=D��M�B}���� J�
m9?!��Y�q�j4�����7�S��$`�!���%��T1� ��"��HpPmK>H_!�Ę�CP��Q�!�`Ebᬃ�z^!� .
����G�30�tq��A��mS!�d�b`�+ŏV.z4�ecҦqf!��¨H�A#̝tg�R#b�6Y!�
�Zc� 3���-X]|���OX�V@!��9~\cRN[=@�(h���D�7H!��̓EWl��u/k�<,q��8�!�䏨8p�D�W�R.I��Љtb߈S�!��M5a#�5C����
�b��&��1�!�� �P�W�A�&@�Ĝ�\l��"O�(ϳ =�q	t��8���"O��C�N	+>�(ը\%V�5qf"O���	,rɼ$ypH��>R4��"O`��c�� B�)8�a/���k�"O<��C�̛n�  q���;E�:y�"O�����E�Q�~�P�x̌Is"O*��ƭI�_J �Fǀ��a�"O֜x�`âz���������q"O�=�qP�0U8�j&��z��|b�"O�L�
%��T�R���v2��E"Oa¶���8B���A�mĠ��"O��x�A���Y�����nn�!c�"O�}�`O�'�Iy�
��d�0@"Ob�Ȃ@X�9vUk�i�!Vf$`�"O�Di�M!Pw��en K7~q��"OL���0�r�YrC��B
`��"O����n\�4T�[���W���"O�\J�۷�$�h��S9�HPxt"OzԨ��~���3��
	�h�;�"O��Xq�
3,��L�>?�z��"Oҹb��B�C3��;,(:�"O|�b䧁�H��i����L���J"O
�A��Ǯ�Rq��Dm+���y��J%Zϼ���� w�� KH=�ybk�h��i��Dε:��0��jS�y��G`8j��)�^�T����y�,�)t�x���BN�̀3�dƅ�y�`�1_�x���e��uK�s�J�1�y�燔&0�(� N��a"��&�*�y�'К.����s��6-�m�i=�y��V�TĠ��e�+R�1E$�!�y���I��=9e�F;gR4TB�6�y� ��~��e#@eP ��{��%�y"�آ����7(��&dC����ybI^mh ��Ä�͸!CVi���yҊ\LP扲`�X(|��\xf�#�yr��"��C�̐<pP"�%,��y2��?U($TH�A��`��$"�#��y��A� c4`�EP	���Ә�y�� H��⎞.7���2D�G�y�\B>�YgB�1C�815���y2��,-�9q�J�8 �|UP�FM��y�,�3Q\���V����/�'�y⭛9u���c��2�bG*P��y��`���`D�cʼ�y�fHO<V=3g�5sx��񢍌��yrA4;����Qm�8@�JR�@�ybnԈN^-��� �+�����`+�y"AJ*, ������\!��R��y��H1`}�Q�O
~�@yW�y�m�9� t�dۧ2���a�L��y"����!3����"V�D"�yb�%����$ �vń�sD��,�y����@�0)2�]�mUj�[�
���y��X3�"���hCR)Sw�$�y���)M���eF��2=h�I�J\�y�*E�o��XA6A��.�ᦌ 9�y�&��(�����"��"�!��y҈�l&�%vOM6�4��a�\��y��ˋ!�0�31�]�]���� L[��y� ��gk�J��	#YDؘ31Â��y*W�H��D �/ԈR����l���ybM�h(�����1OXA�Ť_��y
� �H
� �I���d�[�^�lP)f"OF�{Yyu�l�BD]s�-)�"O��i6aڰ0>f� ��Q�Om��R�"O:� '��V;�hM�TP�["OT�g asZ�0bIvt�"O:�ċ�w�̬"&��<\�"�"OR��Un�$BaP�S"䉸!�|�1"O�5Z��#O�Ƽ�v	�� ���"ON���g
 TR :u)�A�����"O��kA)�2b�f�pH�2��H�U"O�a���Ӛ_��mc����7�2�X�"O��s�߁t��[%F�4oY� {�"O��QC#S�8dZ�d	_P�x��"O�}�s�σ3l0����'77l}R"Oq���K�!d�硑-/Jx��"OؠI��_1��M��$�j��"O6$�r��v�~�{@�"d�Jx2�"Olpe>c���h�a�E8�"O�Y#�BHt+0U#�i%^܌0I�"O�5���@(]�d�Sc�"V�rDK�"OFd����Nf��R����`"O�MS�^�
tı��K�[CxܛP"Ov��ڎ=Ԁ$����F
����"O��i�O_�)R�Y�*�	0�:å"O�J�#�*��v�I�{��)�s"Ob���h�f���[�(�(H�H���"O�lISo�&��0�JV�[Y��f"O� 9�&�((�q�T�WB�|:"Ov���� ��:�
�'ZgČPɱ"O��Ɔ�$I�����	�%�Xx��"O�h:��ɲkX<b�dI""O���d�_63�f�жj��	g�qC�"O��`�q��#��]}�@[T"OԴ��S�	���p��/^��5"OR�Ʌ,W�C)���t��6ְh�c"O2�I"��%c,��#JI�Hϴ�Y!"O�Z�ΐ�<Q1���P8��"O���+�	���+g�(+3�`�"O�k7�÷w�mz���|0T0��"O�Y��P��Lǫ}l<9�"O�ḅȚ#7p:M@�K�of�A!�"O4�	��g; ����Bcx��"O��Ht�L�]yD�X��j퐆"O��Y�
�/sP�9��A�w��R'"OTa�.��R���9z(�=X"O�%s�#�d��#���
�"O^��mUL���,��}�Α��"O�ਓBYv�
Ux1�͔^���9p"O.}�6�گB�}%��~vH&"O:�D ��`����%�6q���"O��!����ht�oe��*�'�RYC��;_z���e%R53Wn ��'=������o�`Au �b�t���'�h�`ć6t`r�����\���'����d�¤	��(��`[�Ob��q�'�"���*ƊH��CG��:��
�'st��qM�<��I��X�1�� 	�'=�q(b�U�0�8� �j�(-�ٰ�'��
$ی6ZX�s
��敳�'���C��Q�0��#�˒)$�#�'����$�)��c��D#��}��'�� �4iƈ+)����6&1��'Lb��!6{��{�j�0��T
�'�q
޴FҜܰ&#�-�.��	��� $���Y�[D�+D�7c^Ɉ"O�pr �4���a���RO�]4"O%������~x��cRr4��"OUi%,C�@`xMY�&֕@a.�QT"OPD�#��Ox^�����OLRtA�"O,##�#�����ԟfItr"O	�f�2,_L䛱f�SJ�`�"O��6@�3�v��V�
f�й��"O�)jC,@��0�#�Z���$"O��%�N5B�y�!�(q����"O�� L�*�5b���#*�^�{1"O�Q ����*�J� m4�0L�f"O(���%�-!�p뛂�PT��"O�Aq L�������.����"O"i��MD�d���ei�����ܑB㉿r�x���%��`�G�#>B�	�&�����Ҥxsukb�J0d�NC䉷o�v��U׭a1�5a��$C�#(f�]6Gk��q�ňY�o�JB��
b�dy��F�tp�R�=\7,B�	.Fͩq+���|d!�`�I�XC�	
��Pz��K�-���T��4�&C�Ip��Zv�E�xk�Ah�����DB�I8X�B��s�͜p�8�P�]2P�(B�ɞ>r����/�ܜ�W@ք7;�C�	�.v�Y;���>�d� ���]RB�I<G�.A
`Ô l�49ꗬ�854�C�		5�n�����M����Ug�I�|C��gv!��tz�sD`O�.�4B��Y��qxe��v�<i˅䋗-$6B䉞/b�����P?q/Z�� �ɐ2tB�	�Q@���oZ#,�, g�(gHB�	="0�t(Wh� eX�I��WJdB�	3���d�'��i'��3>B�I�FE"���|:Zi��j�L}
B�I(�*��-�7en�P	F��kB�	�'�D�U��wO�h���i�<C�	&n�$=�7�J(}�T��aW�,�C�I�XzYR��vX��F�S;'R�B�ɞ�~\���Q�'����C��6�fB䉔�<aYUǕ�b�X�kg�t@B�	+JT"Xk�G��F%�N�j�B�ɸ&�����=E�P�����/��B�	"�>���O#X����[U�B�>L��I�"��	���Y��<#"O���T,�D�l%#F�I,{�~�;F"O�=����#Y�!cP��F+��&"OB���\��B(8�*-Z8�89q"O��˶h�
W���J7P!:�#1"OJ�"�.]�H\P<)����r�E("O��d {���� iA�!�t�Q"O�E��M�+]԰���~�F�Z"O�$�B@$|(<�z�(��_��-��"O��ҵ�C#2i{e�9+��9'"Of��2Jޠ)��c�-�0Xx�"O&�`*�"���I��!u���B"Ozt⡪\��(Z��D
q"OF���D�~ �']�o��2"O�T*�i׫)�H��/Y#*��ݣ$"O�L �X T3���p�c�L�Ү>D��K�'�2J���i�	�+N�� �''D��[�m	�vͪ� ��-j��K3B%D�bǌ/��L�p��x=N�Z6k!D�����P�a.$��N��j�#g*D�� �%(�FD�,QU��U*|ዳ"O�ȓ��ҾH�*q����Gj%�b"O��
��1�����	A�P��"O�u�s�/[�ڹ�k�? �qP�"O�� f�	7y��C�
Ւ��7�y2l�fW2�3C�R��*�Cۛ�yb#�+2�ڔs�٬o��Jv�ؘ�yo��I�
7��?T(\��L�y� �6��آ׬�9��`��e߿�y"��_1���C)���(�g ͊�yB+0\$���2�Dc���yRG&A�n���V+�\̐���2�y�o
�Δ[�)�"�,� c��yB�`�Y��@�Ԉ�`�,�y�G%���RCB�%�0)����y�ȃ�\D�VO� �'�Ŏ�y�X�{�ة0���%�%��޽�y⮟�9�]u�C��\��3k-�y���7;w|hr�Ƙ�H��![�F�:�y�f�t���3S�e�*�N�"g	*���C���h;���A���7n��������勵i��0�P�K�|Іȓ���H4�]8X��q�GBP `n��ȓ�n����R�^���Ub��X����	81y6�җZ�H%I2�ҙx���ȓ6�@�	��_
|�����!5zʩ��&J|  �W(pJ�lb�ǤE��ȓQ\�@6�;J��p ��#VU��ȓ$פ5r5+�"B��ud^!O��$���Pb@�O *H���HG��'�U�SGER�H�a�,��ȓ��ah�xy��ä���E~��ȓaX�A�'�;��2�ѐ
�F�ȓv/�H���$9���$ �j
D�ȓxi`!Nkrh
Ѓ
k�>I�ȓl��X[WO�. �2)�R薞0�FL��u��u��g�>i���!$Y����ȓ1�6��4O�$U80�QD�Z��ȓxah`�H�Nz�7n� �ȓ��Y��gZ���0�'�0L�ȓQ'�%�b镊>��`��	 S/䑅ȓr�Npb���Eϒ�̐�qG�m��IG�5�!#پ`���@��C�`��EE<����E2E̐�D�1{$ĄȓVC��Ӏ΂�O~B���j@�e�����>�`�-�p9�&ţtlNE�ȓR�Щȗ��m����"*H	]}>�ȓ3璱�� ԪDG��3�C1����m���B�ƨI��L@B��n�L���u�|�R!�<����
G.:ެ-��,�T��䔲J�&����1�j���}��Y9El��NBl�g�K<��jF��H�c�/0�IWk�=-����gr@4{ ��,q�R9�ӆñ=2=��$����F��L�慚&1h�Ƥ��"�𜳶əga�`�!$�+^.�݄�z?�h1��8o���yR�ۥIPt�ȓF\6ܡ�$6jnřR�Vpvq�ȓ=R,�7�y(��Iv&�HW2Ɇȓ+�DX:U'�2qI�5���I�� ��b�Fx`gMP��*Y��n)=�ȓ~Ǟ9Yg��%Qz���( bv�%�ȓF�{��0ɰuR�A
7T�B���MU���-U�Ƅȳ+ &��d��S�? `��MK�L;�`�|3���"O�P8d�� ��.@+w;X@��"O�,�I2n�`��B��0Mb��"O�*�6(�����B�{O�<�C"O�E��'�+s�n�u�@"x:J@z"OL�	�^Eq1� d�"Ol	zT�8
~�[�ާ7�J�+�"O�]���?W�ļꠥ:.8�h#�"OV��nW$]4��Q�Br��"O��ڔ�O�{���g��?U�i��"O���f�N�K��ӣK@n$:�p"O����㔼0�p�I"2DR"O��K��°y�a8��)Y�()"t"O���тxp���K8a�v�%"OD����).��!`�(B'X���"Ot]�.N?}ؙq�W/]�<,ȱ"O���Ro�8��Af��n�(�b�"O$�2�.S~����UDQ9�nru"Ot�������\�p�2!�d���"O*�D`G@�uϩm��"O�@Y!G�\��]P��%F9�@��"O\ٔj�;!~��:e6��i�"O�]S"��L�`UyՄ�5y#�m�4"Oz0z�
�w@j�P��]Wh�`��"O\9K��I/K�k�%ـ0�PQ�"Ot�H���.�ԍ"d��\�r��"Ot�S��k�b�`�#�ޒc���yR��L�A ͒>�^��"���y�f�#>��U�H/W�$�9c�@��y��]
6-�  كQ��X�#���y"���x#1@P�D�����X��y�E>	WN�z�/�D'���"Ą�yM��$Y2�DI�2]�G���y2�_73�̹��W�Ap�����y�m�:~f�ݣ���7P��hX�K�	�y�r�БD��7�܀3cM��y`;h�>�-��'�P`ɣ�X��y�L��|�6�L2�2��$�
��yRG-]�F<@�a ���#���y�	�=7��\ٔ�l�!FU��y�8��!��L�O`�-:��G��y�C��X�K�#Rq|p�.D�ࡥ)�Rh�Xk7bջ5hܜ�6D��8o�xҲm�;(�ș�5D�$
s�J����XE1�li6(D���B�Zj������ s�A%D�T
�.�L�i�`�cJ��+��#D�@9n�_�B� ��
�o�P��"D�PQńG["��9V���i����E" D�|с�J�����E&L�p���D:D��H�H��GS^dɤ%�eh@�&D� �6l���X8
3 �#��[#$D�H���nUA�$	ٙ`i �X�#!D�p#�nH��m��SH��Ve>D�+�Jhl�kh�3Z��\��&D��P`ˁ T#j��F�_�y3J%��#D�����)����&ܕ>w�I�d"D��0�
������Q�EՠY�S� D�p� jG�j�	���)!F�����,D���3/�&rd���B-j��֨)D���rc��2�fE�wdԺ7=~y��=D���0i֕!��ä��9�^�� (D��뗅�{00�4G�=FTj%� D�l�F���[�1�T�~jB`�>D�� �tb�M�"P¤�H>QjL�U"OZ���^��8q��7k��}k2"OV���d�Z��YR�ߐ4�b�"O*��+�mo���4��,9���"O�� e�Ê=�A	��|S�9�"O`\j�b�\4�W�
%H�d��"O�e��� �̵�PBX$\)�ei�"O��(�ᖋK�P��@V�?t���"Ot���F��� N;Xrƴ�u"O��H��
v�vO�'$o��`�"O�x� 	hߨ������zhp��"O���dC�8�Q�s��#IbH|�"O��1�;t��[��]�!��eC"O"]��)�=`)*�[Ѫ�D<�|2U"O>a�EC66,R�j�)#	�"O M1u��J�jɑ�f�����"O�5���}���v��\>L���"O6P�0"�bb� (5Ֆ5�\�a�"Opp����h�4�0G��V���3�"O����H�t�B���W�5�,���"O$� r�H9C�~T�G��"T� ���"O޹�ƁDt��iQ��=��e��"O̴ZT�8*���a��>�N���"O��֌]u�!36(wdAP"O��!]Ҡ���C��9�j�RF�1�y�M� _/`(1�Í0�"��eR0�y2�̝];�P$>_�٩e⎘�y�X�\?by��-�'�ظ�k���yb�	9,���nÍ|���B��y"���?�D�i�I�S|ج�kV�y�A�D��Sl�H+r���y�]�7�X� �H����#��y�+ς��$�.C��u�E��y�,Ԭ6�1��W�J����SJ�"�yr��!������@�*��n��y�c=%��H����8i�A��N�yb`͏c����Aӌ2>R�' ���y�mѡe���"tFO1#��h�v�χ�y�JS.y�ix��V�!�v�˕�.�y"�Hq;ѐS@��
i�Vȏ��yR��E\�Q+G�4=���:�IS�y"� <NA64Q���F������(�y"i��Je�ҏ�m���3ˆ�y!ӵt����Wi�W�B5��D��y����/��"��	�R��w��,�y�b��?v���l���L�r����y�,˟7M�Ɋ�眽Ufi�C���y��jni)Fk��tJC���y�E�u�e�3.�;��p�r��yR��:f���c�QX���"���y7 #eˁ4Un���\�y��!'L,80�Ont9�!)�;�yB��f�`��ˏC:�)��"�y�'F�4l^�:�J^�6_̥"W��yb쉼��)�0쓄*�ک��7�yb�*�<�ja�T*���@�&ݚ�y��X��ZyIo�f�C�#X�yR���l�hP�`�̑D�M����y��T�9׺ ���<z����c
�yR��S���2��*�R������y2G%��=#� �UK�`���ŧ�y'�J��yhvf�K�$�k�%[��y��! 3Ȉ�ua�?>,4݂�̆��yR(�U���Cm�6V����fG��y
� p��#w�p�s�.�"[$Ȕ"O��DF)\���3͉�]\�	�"O������0Vxti���̝8SvA0"Oj��aʗ3�^�k�I�P?��+%"O���Ԫ��j�m��$�-w"�!�g"O�,�fF�-^��z�I\�Y�XӀ"O ����ǆIX%	���)P8���"OD��B�rd�A�ƠT/���`B"O���������S���o�|Mp�"O�ŀ�8�`�Ʌ�ZSC��"O�+�i�5"=.��R�hd"O�݃ ᖈt��ڠ�7nu����"OV5�_��n�P�d)��a�"O�� ��b��J^��@�"O�����b���"�ć�z.���"O�y�0e*Yt*���bl�s"O -p������,��m��f=��01"O.�kR/�� ���뇂�uAe��"O��Q��ʸJ�$��*��_&�aF"Of<��앲�ڈ��Ɍ�E(�Ej�"O�YZ�ߕ-Th�5h]�L)��a�"O�(��o��l��IGF:e�@`ʤ"Oh�k��� SR��as$H$	����V"O��#h�vB��C+ � �"OX� ��> H*�B5�N�s���"OzM���Мi���o�?8��s�"O�̀����$��/.ۺ��g"O�Uyg�E2b[�����I*�6�C�"O�-h3B+eA�,N&��5"OtH�KS0	��!;�ķjrjxW"Ot���-��"�q4Iۑau:�I"OJ��ck[�T-iaǛ�-t�t�"Oj����o�ryZV��F��= �"Ol��IH�Q�ސ�&�:)�ޘX�"Oj�9�cU'�*h�!��n�\�8a"O�-����>g���լB�t��"Ot�0��g�������d͜yB"O�Hf2:0� #T�@!k���2"O���+r-�X&��D�� 6"O��*b	RF�T��ƕ2�^��E"O��ے��X�ba%��z�0���"O��y�n��=�)�u��w�Da�S"O�$���!긚၁1d�N"OU�����i�]��F}���G"O�bwKG rpa��2ckT�
6"O�8���3@"��B���e���3"O�њ��D�rJ����I��%ѷ"O�䃃$� �E����S��!"OL]R��J6J�R}�7��;*m�s"O������4�@�㯕��
t{A"O<���r��X�դE>b�t���"O�b3�/���;��ו"��)i@"O��k'�9�i���Lx� k�"O���e.�)����6&Y`+�"O܍����Uzt8�R�oV"�rg"O�e��H���Yc#EBOd���"O�(�@Y�|0���Q�@6"5��"O���7��N\P��va	Gx:���"O���`��%`mjQ3ՊY)Ә�Õ"O`�3���bR0��
߻��Q�3"O��uF�%$ekc��*q�ʕ�2"O1���P�ƕ�� W9m��S�"O܄2'�:�	X��\<��(8�"O\����\.5à�s!�NMМ�-�y
� H|�e�S=6jhÐh�\��1x�"O��XT�Ռ$jZHIRhж�F��a"O~q�l�$hrŁ�ۄK8(
'"O6�X ���\�hł��,�\-�C"O$�k*H7�b��V�4�\uXE"O���JޒW�<�qeO�|�|S7"O\1
�G�NQx��E��[c"OH �Tl@+r$����W�k��Ѐ*OXM�W鞸g{���vCI�M	����'��8�à�v���j�0 � �'V�4Z��]�xq�G�/����'�t-�ᩜ�3���A�CX!�tȡ	�'�^���DGt|���B5Eϖ�A	�'�|e��6-��┴
�x`x�'<8���I�q"u�S��t�hY�}R�@Ux���_n�b%N��0�.>D����E'�R!��`�{�i<D�l��G-&'� ⛭	��"s�>D��H�NƁ�X<�%O�&g��ÂD:D��`�g�<�"Qۆ�U��=@�i-D�`���*�n�{��Ն:}����'D�0k�e��,�`��Q�'�T��R�������7e#S�R
oR�
a� ^e����-��5mT��1� #�v<
��I)��}�IB<�q"�;��0އ%*.�ؠ�~�?! �<%>A��6B�-�D A��Fic�7D��:3��|
ى�e>o4H�p�ʕ���'B�LѶ,۲mQ�i@�G\-4�,���6D���6?���� ځV�$��ԍ�O�C�I�s���4G�1��hb��^�[�\���1���a,���k
O]�aBQI_Y1!���:t�����K��Ԫ���a��L�G���G� �7��pq���r�2�{�K��yr�]�T �t2ئgb+���+��c� Γ����B_,�t�@�uK�!����Mk�J���E��m+5�z� PJ��1���x�Z��G}���J�#����P�茢T����p<*O��'�^-2j�{&H�`qj̹G��	�"O$Ha�(̅��(�ʝ8t���Y�>��'���%��?���	��5�A`� v+�G&D��"g��{�H�e�R��Fe��G���'n���xb���|Y�s��HLX�sd/ɑ��x2f��4� ��ŏ��H3W�O�u��I�հ?s+��6���(��t�DJ�@�W��p�їx"F�'*��K#
ř;��)�A��y#5�����E5�A҆gU��y� [<��a�A`W�@�X����ȧ�y-H .E���e� 00)��N4tь�<���Ov�2�j�/T�|A����c��M�s"O$�B5`ֽd��=�Ċ��x��:Oj��d׎V��h� ��н�� �W�!�\O����P�j|*��E�%#!�ē���՘I�4vd�1�C֊��x��I$B,(�$B�q�`1'{V�C�I�\��f֮"�������v��C��,�Z�r�a�z�n�j��B�%b<B�mG�T�	\p[�_	@��C䉲@�@)����n=8���@�h����D�<ј'���ـ���L��р���]	~`H�'�a�ŏK��Pa!d�>�0�7����O$#~�BD����tB��B�����Prx��Fx ��X�R=qZ$` A����d�"��"}�d�X e�4@�j7~�r�aÑ\�Ƀu�Q�b?��PL�Uo��2Y;�d�c��+D�� �I3�@/i�\9��H�P��ʇ�$�� ǉ'��4��� (ӊT�AN�Z�@D�1�g������H���F�"���U gL:X'o!D����-E��j�"�f������>�O�Od ӷЙw���8���PE�R�D���D��.�/J�QBa�<������.�'$�6�)�	�>RJ(�r-J�&�������kZ!�$]�Oe���s�'_�d�1 J(O�q��I�hO��8���*�^W�<3҆I����d�>A���=C����k˓
mf�2�dJ3D]ȝ��hO��(�A�X���-�v���2�1T�	7��ɧh'1�6�) �Y�%XL�X@dK�+�$�P"O2$�V�݈yp�I�A];r20�S�,*���S���ЩI�B����C�i�0C��S�4�p�"�&nvBiH� �G�˓?��I�߸'��Y����&�
�&�SS�G�gE之wg-�O�	��8C���q�̨��eޗq���x��9�S�ԫ�0�V��S��i�"�
���hO��D#�<`���"X9���z҅V�k�n�T���<y�O�s0>���`�7��=��1lO����
��;��X�b׺t�`�{�p��=E��4�؉�A� =�~�VF%Jޙ�ȓs�ȘY���fID�ү���X�	N<�0���F�S�)�di��ͥOӧ���&g�-F)�M�6.4%�ת\!�yBM�X�j ���9/���6�B�y2�P�8�4u34��6)B�$25��yr-D� ��`򎏾$Ơ��ÌG([���^ZhZ�Y���g8:d#�&�EQ�`&�%�(�7��Zv(D�&�<Y� ^;`����?yrg�hp�U	�6fD{ƪҌ'z5�'/��ip���o�v��|Γ��(�ǭ�zi�!Q��Y3Z���*����x?a���Yh�L-�aר���jD��1I�'D�	��X��r_��H�&H.���U���U��j*O��=E��ǡ@b�
��[?E������M����a�'���3�bU�YS�쑧�ALh̺I>q�n��yP�Ď&F���AY�ܠ���l��BD��8a�� �6Շȓ^0d����"���!W�>=�&1�ȓO;>�0%Ξ�Aپ�ab(�<jL�'�ў"|���� f�J��Q�C)"�B���r�<q���4���K�/��j�)���o�<�&���Q��!�!՞�dR�mC@�<i��&i���"�Ʋ#4��qSx�<�$"؉U)r�H��12�x� ��u?���3�I	��֞oTmP��ʨo+�C��_b�쨷��"�6�r�� !ؚC䉑b���R"��l$l̘7˂%�l���2}�=l���Z2������M���'��z��p��g�ƵZh<}���K���0>��͛0)Z��1�̸O���6a�R�n�L
��?O.8T��f�5{O�x��1D�hcPd�*`[��q�M���t��a/D�hʷ�KUN��e�تw|� *D����A\iܙs�J�<\��)D��;!�RF�j�Y&L�zԜMH�I-D�X�d�K!^]x���w�5��0D�����HS8���V�o�vUQ�L2D��3�G�@�ylѲO��(���.�It���kê�X���8�,z��H�@.4�\��Z��ek�f��/&���IID�<QNj1�-j�k���|���JA�<��N@q�� I*���i@�<A@ET��< �

B�X��r�Ay�<� �<��Znh�΀
8�E��"O"�����U�Fd2�c/f��h�i���Gy���i�4D�`o�V��(�۫m 8)A�'LV*d��-� ,��m�j��Q�ON��$T�'X���u�٤Q��խ��.t!�$V+�n%�Pn@�CBe:���"r�!�Z�?N�mj�4����iP24�1O4�=�|�EG�~a��
ߺbE�fb�<�BÂ*�&��:P|H����t�<9A̙��<}�rkM6Rgܱ�W�[�<�2$��7���qĄʖJ��T� �S�<��J@������a��J�͐H����<�פ <(�&)�3!�m� �!{�<i�A��n��=���ۊt�z��IL����?)A���k�`�*!�G�tŶ���m�<�#k��i2�)�ւ��Mz$�zc��i�<�� T�<q� �Gܒ+�ZQ�EQ�<���*u.�(C���S"$�A��v�<��`�'����6�G�8�Er�<I&,��W�N���+T��/ZB�<Y���(' �uA�`��82��@�<)�۶�Lٳ�����I��Ȕb�<��(���zDݓŐ��rAU�<�3`��N���CC�p#�H��j�<!�\�J�IS�Y��M9�Hf�<�P�ӡS�r1��EèhA��ȃ�a�<�3A�1x( ���aE�S�2宇Y�<���8r��x��O�{$���H�}�<�'m��<�)���5�! n�y�<��Z�/޾���iC�qvU���s�<9�j"�:؛@�J7y�|ya��t�<��`\����&U�x^�8�A�U�<���H?&*6������H�`"c
x�<�$�ؕ/)<5a�D�E��t���p�<)waڻ��! aJ����Im�<9T�Xe��W�T�?I,=��B�i�<Q�'U�p�*0�B�ß�l@9���<�K�~ƶ@��'	p�8ԉTS�<��I*b|HP�*�@���p��h�<���Y�~��r�Wf��1)��h�<�aFI"IK�h��"z8��~�<��S�>�n���ta���OHT�<���V�cӖ52f�c����ૅQ�<��)X)�b�*�"8*��S ��L�<��B��S_�:#L�9W��Q�L�N�<i�l�v�v���b_84`���mMG�<y	��o\�Y���IA;zm9�hY�<�A���vU[WK�1\T��N�@�<�Q��K���t�P")�!�`�~�<9�)�<.�B�SV�˶M������P�<i"a�C~Πځ#��4�.�[fN�<I�k�ga�eD
��!׎D"s��}C�fХVSh�9T�/LOT� аIw��0�ײ��3�"OFlx�gK�,��v�^�� �"OޱI⩞�nn�Ԃ
"�"��"O�x�狏?F�Z���PT����"O�OY'�,Dh� ��-�@��f"O+���Nے�2�g�%M2��"FQ�<Y���	Q��sA���t�3T[�<��C<lr.xYD`ȉ�v�k�Q�<)U��Q��ܐ�@�O���p�@�<y�C�EV�h����!^�a���F�<Y�Y6,c��a%�/�&�`��RZ�<�T��nDZ��u��Z���%�i�<� ���M���ի!o�=l��B�"O��I�j�|8�!k�Q�T��"O8�[&��=5�̑��H�8��"O���DƗ,�i�a��'�� "O<x��n]�F�(�GJKT�Ap"O��;�0i�v]��*==f�E#�"O�3dmF-!
����%]v�+S"O���N�m�Z�`�i�y_�t�'"O��C,ڃ~�¸h��C�%�L��"O��R�gPH�>���	*� p+�R�L��$� &��|�Ū��6	�MA�̈%��dD�<��掶s8�p�ᑆ iL-�(E	��#E،r$�P���g�h�E�7�&�l��2B�@]��	2Q\�9f�J�Rq�1Eߺ:���7��2~�xakUG؟�2ᢋ�)徙�`�:8:��i�>�*�(��4���K|�P�"4����%E�to�iAD�@S�<9��F�h����J���(iG?��SAlLd��, ��퓤���Zd�8nlؒ��)k�B�������l@<T�Ȑ!б+0�p(OXDYp���Fȶ�8K?�4���`������R޲����9�O�qZv��w�-q� �,˲��
#rFQ���X�$
v���ښ��`�m�1B��s�ޯ<iQ��i�h�4*Ӳ�QC��I⓲<x���$I��Yb��xN�B�IKQ�ղ`��6a�L���K�DR��
Ѻc@��EZf���h�Ψ�Ȱvv �"��JS0��X"O2}�V��'& ����?892"3}r)	�q2tdZ$>����."��8��a@,c?L�R kC8<���.#�����F�"����bť	�)s�M�
n!�A�iOJ�3SF(����*G*�!��!�B�jG��4�mI�1)�!��+ M0��͆ �m��M��!�DOlւu��E۵e��1e.��Qr!�dM6G�L-�$]��	C��X7#`!�$ף!2la�l�e,Б�%�ÿ=j!�d� Ҳ|X��V60��j�L�#uB!� .>D��i��!)���i�!�$H%_��r5�ݰg"إ	�@�	5W!��"��2BĔ&�E�5�E�!򄈌{l�h��N-u(����Fj�!��M�~f(�&�Bx����A-u!��� ��W�	4C�캲�DZf!���u��H���V��d�1Z�.T!�$�"J �0�k�)�$ȃ+C�6B!��)��Ջ`E߀[ײ AJ�K,!��0wG��0�ح���行� $w!򤖳pN����;�(�`�S`!��N%Z�n�{b�//0���d)O�K5!�$�0 ��\�PH͏R"M@��3,�!�$��/�,�SU
|M\�P�%��;�!�$�>\��ӓ'R:v7ƀ8��țh�!�d�9�LĒ->����T�N�a�	�Yq�AIs�1��kG��ں胃���5�Dh��'p�%$I�,!�TMHǠ߻1�fX��'�n$����O�V}�&,ϐ1`���'��4�����T;�@�7)����I<�fl�>oS��b?Ii��3Z���#��U�q�ֱ9WN3D���Ow,�;t�P���8!O���b	9irj^`�g̓�X!j7��+����j2xa��I�'��b�,i�0��(3 `d�!É �Va����}r��!ۘh CE u�ղ�W'�O@�K@�!�P��.E�|�UkDo��Ƅ�a�ם�y���u)4nȤ!I&�I6fQ>�ZcTՂ�	(�4-1�CZ \���'�挠b�S�`=��%���[bQ>�̻)U��2�^7����K��r�٭q��My�n�b��)C�𻴭�mj��v�?|�h��>Iݴ��6���?��_w[���6.!�Iԧ�  �إI	�=UB�bv�5��-���'����I?<2�1k�a�DI�E�5ݐ��E�2��A�i��#ZޱB�MY�VP�1)^��韼�O�XВ��y  �c�����}҇��3�e7�f��aI�8�� Ӆ�G�����ɡ�ލr��<K�l������,J�M]h��">�?�'"�s ��8o5��0�������i��3���s>� C�7ZN����ē�\p�"�<�'BxN���D��0R�	b�.`}���'E4��Pʘ/�yY��@��I�B�����Qf&t|��D��u�cC��BQ`*lT���>!RE���j<�GӬU:��`@�u؞`���i�(8�ɗ G���P�X
w�r��II�4���sB�L�
i�� '.;x���3�K8#b���O$��Z�i�=L�����L���"�͢[O�O��Y�4'0�ud_�*]�T2d��6e�jZw�M���X�Q *��bȨ��Dnۆ=8H��A�IK�g�DǭegJ\��ǥ��7*�5K$d��43&��3c��#?^�X��0`9+[w��O4�]57=�@�R22D�E
��Pc��K+aU��ɷ_-���t�#={>��po��(N�T�5Y(OV0��
����RDlݽ ���R0��g�O��ѪON�B����vO�Q��]Ϯ:�'h��I�BCH�(�:e۔5�C���#|�Q��Gq4�mX�9��8��z�N����'q���>q�߀H�:�%G5(+���_����͘~ |��Քݮ� `� +}܀�g�Q�c��K��ƒA�t �%ѵB1Y��޺�a~�c��f���ZjX�yx���b؟ >��ή7�����/3��1�#�����U�G���飥1>C�G�?	b�q�!P�ܔj@�8�!�,"�}"���0E�4�@�Af��b]�{b�I2�id`Ƽ/%�i:�OD�8� A[�Cl��ap }���Ʒj���چ��Kty��Il�±���Ov}6gҶ%���0-V�Zk�� u�l8+N[��f���'�|�-��'��D|a/�J��8G��A�b����r���ۢͥ<auץA��5.�~�U#`H� '�f���edX3n)�� �ŋq7x��dI�w!\��c��-4���2�,8`J��'iH9�E���uʚ�S?�����X� ��vs��ځ(�(H]�%�J?ƍ��,���qH\�K��� ��  -d=�`�� ���	�%�:���2�S��r���gة��tB�9@��q��'��Y P��^<Y_4P���X�(c.�{jS�p�͛M>q2ꓛq���|�	u��T�p��$�2��&�ȽP�\CT���]29�$��G'�#r�D��2��1��%�C��.~vqO��m�W~��<��M�	��r1H�0K1�T�#ft�<IDJ߲�xq#TD
�2x±���<����5GB����	�Sl�����6yz��[ӂ�|�t��$�ċ�;O��������>�5:��'FRMks��E�ҩ!��5��hۢ�[xm��AThݚ��'����hPz�S�tE�2����Uu��3u�F��y�*D�Ѫ0VO2<9��4�B��%���<E��':�L�6�ѰrKX����Kl$t��'I ��SiD.}u�ʰ�G�L b-�d�:�B��7�o8�H{�œ
d.����:r$��%+<O����D_;v,��O@�ʔ�	�Q��:�A��� G �y���~T��d˜�Du�5�7-ʻ��Er��GM*�)��N��<$�&�$h*XC�ɝW0�L[�n�'���e"�Y�{B�5���D��,�!�#O$���������0����!�� ����2u��̱����$T$cM���g)�m��SR,?1wJU���z�������8$�f�CW>Qⲋ�"D��'&XE�6����H%���md�$��'�l��M	 S��|:���?��!3��V?qے
ʦ!LM��[r�����-O�������`���܊CX�\Q�'3�$���6TR��3`vd���Q=_�x0�G�����lvO�I����n^Ժ" �A6*��B��%[ �C��;#�"|��JT�!��m�D��bZ��0!d�d�<�����f@�F��-s���x�jAe�<q�P9��P�S�2.�5RH�^�<9R��sHBP��*w�T		5�_�<QPmMx�؂��A�'�r�`LT�<�$���5	�H� ��\�"��bDN�<Y4g̖����n]>L��:�/NW�<�d슔^�nl�"ӹS��"h�W�<��ְBP���^�h�EDe�<Q��ۥv�� BG��J@+���{�<� �:b�\�d2+ѣa�r)c��'�XY��)�Ovq��D�{_�e�h�+z�by���'Mry��������l�B$RͣF��>y�)�2";��R�dS�>�
����R\�<q���R�&	x�C�x`8PfC�Z}�@Q��+3 ��q�$[�O���2E>�)�92���C�`C|�w�#Ra}2��gM��	�L��-+�� l�~���`وA��)��O��~�c��Hr����{��	�"lפ	'+Tm��HO��2d����O �(4�(�b`t1&���̞�jњ A�ЪS
���I�7k���ķf%^L�� Qv�6�̝��{����XL��Z	�t�7iڽ��=��M���56vx\c�F���'���h1L�6�@ē�h�-�ʮO��X��@���@1O���?����e"�UyL~2s遡d �TIA�.3o��(��Zlx��0����<r�\/$��Qz�S$H���Q*إ"u��R_�(IJe��T� ��&Ur ���$T_�2��BۇBa*y�#��.�����[� $�%Ͻe�N8�r�-@���C�dX����:�d!Z��,;�#?頇�-b�t�hFH�hQ��1��X�'��5�1B�"h�A��0�xۅ��.Asrub#��)%iV�Sd�� ���*dg7�O��3BMX s|�*�aB�t���䑟�>�,��'֎`g��,�%>�Z*�?Jf����A�<��!"2D�� P޳\�K�/�*�Pcϕ�Z��I.L���DB̼T"n�}B��+��$l���M�]���V:ys�����\SA� �|�4=S@/W8Q�b����>i�@^�u���I~�=i�㏉n�� 8��Z##�(�[�R��$y�#O���aiV�ټR���$�1 �@XSA�^�gDa���O`��jsN�6zf����ˁ�0<	�qw$��K>9�fO6C��X��ߐ�l�v)�O�<���A!D��i��`t�	��Gn�dA���{��T�W���Cæ_!������y�o��z���V��Izr���y���;5(�*5cW5���%��y��ђk��� ��R�6���P���ybHg�X���*2���-���y �	4�� ^�,j���0"Ȏ�y��� ��ZՊ��^��S�y�(�!fb4%Ef�#�x�s%ǩ�yr�.#V
`�Q�'z��z����y2'2$�,����<l�0����y2��5))`]�!��+	�WҪ�y�e�k�|�[�U�P���ފ�yK�VEh�����z��ȒcL[�y�
�>l��鋱b��#*���y�^��M�������?�y�T/_{<;���tOz�h���d�<��IՖ9"�!S�Oڻ;"!��Kn�<�UCаE���[���4f��b�\C�<��a�IBtQA��7�b\J�Kb�<	4n�8f��Ѣ��I3��!aF	\�<c��U:����.
� -�Ⱥ'��Z�<���-����̕>�P�b�K�M�<� Q� ���0��+����׃CW�<�@KI��L��� ��(��v�<�Pe�z0֜vJ�N!:���+�h�<��&��x��ѻ��X�[ԅ ��a�<�c\�,&r�H�%����FA_�<Qc��Y&duc��H12L��@��^�<��䈝�q�E��Tj4��Ěa�<q����R�ɞ'�4c�M��C�	�)G�s�Y2_r:���f�P��B䉌f�zp3Vc-1N6�1*ϴ�B�I?-a�)�3��>&�0�*�Ǌ>�B䉽D	4a��E� T5�˕�H�=��B�	��1��56e>]`Ff�7@�B�4��3���3.�$����J8EVB�	s��e�$�,BvM�r���C� B�)� "T�c�1k������)t�M�"OR�!�|�Ġ�(	�3��"Ox9�E�2b̒�3(]�jx�� "O\	���3���[�&0}�����"O�i�OȤErf��'T��Qr�"O�l��S=Q�lu�Pk�����"O
�˷IDi�b�*�,�/���hd"O�����"Mo<��w�y�ݻ�"Oti� FWC0��q�OV#Wk�@S�"O����Ǭx�|[���6I��9�"On@��i�]���f�ԨdHV"O
<x6�ٕ���+��mm~�+"Oڙ��lӹ}����ީg~�a�"O���1�Y6<B���3p�\�[�t 0H�/'�8�%��|��,]O0��X�%	�yD��h�<av�0��-S ٧xr$)E&ɦ��I�N��<`*L���g�;�|4&�؁+�}���
6�����l���ʡ�ұ(6"s�iZ�ٴ�G� �B `؟���ĕy<�	����k۞)0
 �I�B|�g#�>�\h�N|2Gd ��Th�I;T�jFNw�<��jO8���g�3<�c5j�q?A�GX;&��A)_���퓉XW�<!�AG�4d<�z��	2�C�	����J�ƍ�1Nꑳ��yObu�(O�,��N5q��M?�a���,ii>y��1{,�`�.�O���\1vH�RGǕ0)\uѦ�T�>b����U�vqX��)d��<K@D�2�2�Y��& �Q��b�N�N �j�S[�S��(�`�
=y�f���k� �B䉡r�E��gǌ	�4�ㆆ8c��	<?>jP��@41�Ŕ�h���ӓoP�eR��f�@;=��u"O�I��	�7�f��b����=}��;/6$R�k"�����Hw��Bb֨�:�,�b��Iu�c!Z��A0�-�+vermq ^97!��J�R��w&��\`h����ϙ 	!�đYNH�!�a�O��Ȗ�=K�!��Y\��+!	��5�ܳ��e�!��	T�.��5����
9!��nptw
�Z��K�gM<!�ŭ'O"!��C�S��1��m�|�!�D�e���/AN����!�U��!�$�f���&r�T�隑�!��E�D�.�x�%�%n�E �e!�Z�p�,Q�SI��M����F�B�!�$T�Pb(S�N>R�w@ێW�!�dW#`S�}���F8t��Ǜ.�!������t��dD�a��O̒oL!��B�<yBVƐ}�>���G!���_���٠HV,�L9v��s�!�1Ӏ�a���#'�8��F'�?�!��P�(�J���FKF��d���C!�$Q�<р�k�2o�|	9t�]/ !��B��y�7���m',�J4�*X!��2M�|d��ɄO6�4�ӔC !�d6�ZG��	-�p3&kF�<*!�DJ'<��U�# �8���_�|�!򤆄]k�쀷c��k�����H�!�䁾esr�V�;~D1�� (p!�D���-��J��+����i��e!��M=�0�3gCL ڕG�_k!�Ĝ˨�h���⦥���1;Q!�V�"���BT@�k����eT/h&!�$�	�TKѤ�$j89��ܼ:�!�d�*?�q����'2��HQl��.�!򄐼�9t�6;O<��k5'!�$�C ��T�6ul�$�ԬC�!�� 
5���˭~�0]�į��}�$����#=qO�����Y����S�zknu"V����$�26b D�x��fE�w�$X����=�,�ƭ��^l\�Sw�ux���f��`.�P!��0Q� m�F<<O�X	pl
�R�*e��OD�+��Y�Y�p+�eI�Q��8��"O(����+8��H��Z�t��07�|�dڒp��pW�|�O���VD"d=��ˁ�U�2����Z}:Ӈ�>Q�h��H��� ���^��p�.� �ĝ>�U����� R��V��k�܉	�*\�c��'J�a�0LE����U�"�9��}R�I`
1/f	�̓�V�d����-`f�%*��X���$�B�	0-P�d��'��Oi&MytE�#8*M�'� �a�EL�q���bF�BTB	�'EjL3fh�1\��v���)�N	@Q��5`��IIC@�n�ƨ�®�Aj�'�1��ih��7 �z�˖ӸT0H�s�'������W�VH�I:��/ܩLQ�l2a��Z��aC�@��$0|�0��L�� ^!^��x��љ|�H`@��!�ɾO#$�6 ��?e�R�VL��Y��Q:�F�c�"-!b9��_x���F
1@E)���a�`��cD �bF]&��Sq�~"���O Q�O��۶�Ϡ)yx���OW�]�Ua�"O�ij����2e��.%�,b���&Dھ�{ /җ웶���@iX$Ô�I�V�@�����'��8�Jښe�,���ɀ=#�����Y�Xa+�I�4P��� b�biPC&M2
ɖ(S �Ō�0?qS�=]Ҙ��GЬD!Җ�o�b��I�L�6jN�mڗ6���A�+Љ6i�����B�ƍfn2U��/�+7|�C�k]����>� qql�]7z����?!q�˞8�%�7�'�yR�E�=����t&}��.�yBo��m�A�ɂe]�Y:�0E����H���l�f�q��'!�š�h��v`%����B�?:Ӟ�XV�:����r욐t��u`ৈ�c��K0�'��y2V��)q��u�?�N�"�G� �C+՗(f���:���ٽ@�V��̳W��Ć�H��`N;}N� 6��*bʤ�O�ba�ΪVA��'K�b�9���u��t(�K�9Z��܅�f��b!��2c��`�Gg�"R�HAVI0�D@" W�\�~&�쳤�?7Hb8���;�Ȩ[�!(4�xᒯ4|��iA)�^5F�)�K+/��I�G�'��q�p��nF�C�6���0D��B!Νs��p�g��x���z��.D�(1�R)����9���qEa#D�T����&꽩%
_�ʨ�4l>D�|#d��G����ɝ4f����?D��i�C3[전�V���T�(��c�?D���0�C7Tm�]X�`
?F�DIfd<D����@��J�(�@.�� E����;D�hs�a-f"�]SɉuS�]�r"9D�p���R�s52�5����P@%1D��J�g�ovࢢ
�b�2�k�I/D���%��)�m2�b$o����B�,D�x��ǧZ� i�É�/lrIH5�9D�0�7�_�Jx�I�r�ϰF�zaX�
4D��k��w��T�@�ȍO?HuA�
!D�܈���gB8�CJ�r�Ts�"!D�|9$J��T��Uhe*D�g(�`e� D�`3�!� \�`xAE�&)#�e!D�t�i-x�JP���CN>� +��-D�`c��?GS��K�n G%�0y�$D�t��@æH���S�Ç0冸[�)D��i��Ó%d\��D�#;��Y��+D��	�CW����,���RD9�-D� ��m��wD���ԖH,	�%*D�����%^
�̦ �A�%D��6�Z
��â�6���#%D��8�mE�Q��-�R('+R��c�%D��IP�֒H�d�1ӤŨl�R�V�&D�� �´b�S�,(�a� (J�HY&"O��k��_�Z%��`�/m���"O�ܠ����jo��N��}���d"On$�6�Q�I*B����|b��r�"O۲��Y�:.D�(q���4�G"O8�����%H�s2隄H��=���'�P0ю�d�dܘRӃ�E7L�����8�|݇ȓ������q�0��&(Ж���'�q��P�,6ɧ��8t/�w�l�["���{��b�"O��D�I���`�
M,'d��q���ZH�  ��)�����H�PN�%���y�ō�'R�����g+Y���=�4.����۲F۳t������	؀ �閟4��)�0�V�D��?qSb��]r�<��l�<���9��X螡*��I��ӃK&�T�3@>�T�
�s �������� �<�4b�`k6l��F�>I�N���8+K~�4n�@���`م%&JIe�QD�<� �NT|d.�挒o�\ l� �O0�aS�4x_|�j�+ �)Ե{Yv�b�O�*��ʑ{�� Q�o�D���0E�'V�j�Ɨv�qקR� �ڜ����&R{r\Y���]?y_�E(@'�>=�"?� L��p��j��؈�X!�ń�V�'/�qx�Kݓ`&~���,�!��R�_�6��V-��]k�
��2}�u-3�Oh!!"�-68"2J��!�KQ��h`�ԟ/G,�' He�b�� '��`%>�!nw=�@���X(��F�8D��W.s�<d�P�ٜh�r����<����#a�U�N����Oо�"U�leGL5!��(���v 0i��"D���QU��i�G�Yh-�M^)����0
�-}�3�	04�*�QqO�(<|�*��̴����Ę�6�$�I�D�\�<��EBM��J�L'OI�����bv�ƈ ��`�_�
8��I�J3L���G��&P��8��ȣ<�l��@h?*C�	�y��D#V#U(T/���@T#�z�'�Z\�W��h�S��nW<��E�T@��A�J2)����ȓ�`�)㠟hPEA�Cnŵ6"O�h���B?q_�+��A���YR�"O��#���"|S��)bgT��"O��)�3?�i4b-l"q{�"O���P��$�3bˇ=�J�r�"O��)�)A3����C�@KX|��"ONu�5�F7N�|[��#~��"O>q�7
�27���$�P�W�:�+v"O$�I�@ �G�Z�נ�+,Ң��`"O ���Ƹ͆��O�FuVAʵ"O�x�g�67*��Pнr4z�P"O�q-Z3Ja���B�2���@�"O^X�6��2jX�rP�%E�� �"O�1�e�Ȏ?#:uAf!�	s����"O���� P��  �$z����"O��)�c] W�t�/��T��"O\�W���5z.�2 �W NЎ!x�"O$b��Ԧd��mq���QŘP�"O������[	D�Y"�;��#S"O�� r�ȯ8��q'C��BxZ@"O\�#�e�#:�J��a��r��A�"O�$�7�P?9@d����a�#5D�����"$�Y��\���)��2D��ಪ;��h� ������iA�:D�<�O�-��A�b��Z��t �6D��
eF(y��	�sV�"�.xJ��6D�l���4c���ЀC�R8lXd7D����6z�~�����-��b0V�<��P��	�:h`�����b!��}�b��F ���?�O�>Țs�76�Q�A�\TX!���,9F��ys��OV8�U����0|��(H�8���&�U �l)m�⌉��'�.hJ�A�P�����/~�޶�
b�'6C�R�摓�?��`�* ntj#���k��i͙"0��� Q���Z��O3W�֘�0 BN����.UH�0�)�'f�֩�3� 0�B���6p���UMG�*N��Q-���mW/�^�vģ��ԑ>�0�V00G�^��Q�P�-00�KE�sE�a`� ���)�''��{��Sn�XS��w�Hz�>wkb$2�V��{2�OaRX���N�
Y��晫Z�v��e����Ot�Ʌ�����i�b5��*ٛS�����2S�R�2�y��'w$A�揗�!�BhS�D$u�t��
�'Y8��4��	/R�De� y@Ls�'�ؘ�@Î�TyָR��P5L�4 *OP�=E�4(�_�}8e��;>���é�!�?����/I�F�9���I�j��g�<E�H�ȓv��M��/ٟ�~t��˹.�>-�'�ў"|���QrG���a Tc�<4�₈�<)/O���<�f�A�'2��9�f�Ir�~Иr���@�bxlں'�.9!R4�)�禍*��[�Xa���{�D�d��O������
V]Ȕh�-U�z��'����D��@����	y�|������hb
+l%(��e�,0jXH�'��IX�)§�(ժ'ED��4XF�'_2�<���D8��S�y���а�՘CW,u��HS4��`�׈͍JX�%�����PZ,`a"�Z &�t�[Q�N�\���"}��^�-���?��OΊ,����|������y������x�N�7hA-������gܓ5<��9V@��,����=�(��24�M��@�dT�X*%�t��¡(D�h� �5U���pq�K57��=��N(D�ٔ���`@���1-��剄K!D��E].~(x4��4Y��4�!���N<��Ig��U� @�B���$!�$I�8B�[�&C"IJ�nÿA�!�DL�k<�x�c�6��t�(�!�$)mj���/ɑO+�,B�M�S!�D��a�Jd�#�������F�o!�$��B�ȍ�c�$���XuE�w�!� /PnDٹD$Jk���p�@B�!�dġcOv��5(�Z�����S!��8�̈���*������)TW!�M4/��f	� N됽��B\�G!�d��t��A�C��<,6D+B��>BR!�DλsX�!�CNq�ʷl<c>!�dΉ9�D�Y%"�+
[80A	�n�!�dY�;\�rG)m@�9�W /�!��<g̱qE��2!���Ul�9N¡򤗒p�dK3��0�։�e"@+�yR��V)���a��)�prR��4�y�M��`�PPy2���v6l��A�O��y	u��`�6'~6��S6F�2�y�Bؤ=�t�!��5qb���E'�y� S�.>4I�'$?,�HK���y�@��C�uأ[��@Y)� �y�)F
c��k��ǡ)��P�&��yr�,G����ą+�F=�a$J=�yb����~��d�J�q���_�y��o�z�P����a@(C*��y"��MPP���+�N�hD"�͈ �y�,�(�F9���@9�!(ҢI�ybG5E���EV/?6���A�͍�yr�ۅ��M[A��
IP�pց�y��7q�T�[�hD��.�f��yU�e%�B�12�Ju3�i��y��іLw MaUe��)sj�h�aG�yR�G��c�M��(���V�լ�yrMK/?���0���H��ќ�y2��Z���;d�Qa�\]�D ��y2g�~}x!���"gw�p�"aս�y�(��*b>=��	=\	B:2Jƽ�y�E�(�pMkE! "=v�Eh����y
� |X���5?��1�#�˷!��$"O$4)��U2\��RV`Gh���E"O�4ôj�&E�z���ō�}L�c�"O6�[3+F�tψ� O�C���r�"O�Dh3'[}~����/x���u"OZ �� îD�Y��+�W�����"O�}�ت �	r�꘽)��$"�"O��4�G�/��Q�o�?(��(s"OcS�H<xZm�Շ�H�V$ҷ"Opx���گ<ߴ0�� ����"O����]�Og���
E�d�{"O���-�%SM�L�4�R��⠐�"O4mI���! ��y�w�P�U$�D�F"O�x�N�.x�FH1"��"OP�&I����ə��$�H�"O0�s����,AR�2#��]M�Q�'"OP�+� �7v�Kڭ':��b(�,�ybN�3��# �E��8�ȡ�y�	F�-�ȨЧ�ߧ{�I��y�SѸk3eC�rO��cTO�8�yr`.H���\���|��ո�y2�,t>��BD�I<�V ybա�y�aU�nZ �4�� 8C�S�A�:�yB�/2�fp���@�Zb���y��ק ��Ag�ӄK<��J�+�y��-?Ɩ��#)<��j��W��y�r���Ä! T���Q�۩�y�j�lf�P��ڣB�Xtҥ�D��y�.]�+l�}0���>z�h1%"��y�+U
������9j^�d�3�y�)ZL�ܠ�n+��ـ����y�)�����CՂ�&��Ն�yB� D7R�{B'J�"��A����y�!��/Dq��I�
H�6 F�y"�״Q6���ƶ+?4�y��ϫ�y��T�SS>E�J_�+E4T��.Ȑ�yB��-J8�$�PH@�M�r�z�����y���</d�i5Mױ71Zhs��̋�y��A����7.�ȱ��y�*�V~�"�΁4�Ρ�Sn"�yR�
/p
^�9�\j@d)vK��y2M�J:�Ke��d�2¦��>�y�$	7w�,�q��Q���J��y�o��U .-.m��9�d�nԄȓ�|`��D	��>�D��g,��ȓ@D�� NΝzЙ�M]�kD̆ȓ@Zh�� �?#[�)ᒠӔDw*E��$�4�Օ��̐vC@6葇�]��9���4ʔi@hδy�DP��K�0��t�V�M��8�	3b��ȓ"�Ԃ2H��"�9��iУZY5��3���$ƀU���J�|���ȓ, ]b��&T$���!�z�\9�ȓ	�nP��&�23��U ���,К��ȓ��1"G-��Q�%n�g��M��ts2��5.	���;���!����lA�\�~c5�S@?ZA��8��%a�/pL�bP�J2f�$��*M����&s\��J�ꄾ@rHȇ�e�b��h�&J���4�
�4��Ʉ�Ӻ�a��F�Zl[DE�q��`��j����7n�i~��UN��0�v��ȓ%x�:����U�̵B
H$ϔD��;�x��RjO"S�. �Oۏ7:l��S�? ި��"\%v�Dp����,p��"O�@��ƙ���b����i��t@r"O,��v�y�d[ �1KȪ���"O��@KҌNv��֏H�����"O�0s��`
�rUl2�h"O�U��k��3>��W��$��B"O�D���П���"���.(z�"O�8�� >=������ڒ)�� ;�"O�MA5&6����I����(�"OdZp��Nz�� Թ/ʺ�s�"O|�X�BLh�D����f��L!"O� c��[�>8 ���DޡF�4@�"O�m{a�Tlt (�@+�R]�t"O2u�c %5g�x%��M�ظ��"O���I�U>R�j0"ǈb�ưˠ"O�PA�ą�m 	A�@��^U@P��"O�R�A�/n�ă2��ZJ ��"O�)�+O�Ux��Pr��Z!t`S"O��#д)T�p�P/X$"O�A��MKc(��B���i�0"O�lZ&W�@ 2�̘�䬻�"O������|V��C���91�¥"ONMyBۂ@��#EO1Z(�1"O�5��-H��!���U:@���"O����U,|�nm���O$ClE�4"OpĹ6�W'��x3E��W�e+6"O �h���A>ؚP��!ژ��"O\| ��	? �r�4��"OFpIVdф5Gf=2��I~�1�""O��@��ަ�����צ���"OL�YR`��F.J ��5D�'�y��E��ni�0}H$�#U����y�
-R�����.}������;�y��+"��↠�����R��ƶ�y&��f<nD*��YCC��Ar,	:�y�	�x�d��ϐ;l>@X�LE��yr)@f�|A������K�y�����<
���
�(C%L4�yB�_�"j�x�*�7���z3Ϟ)�y2#ݰ@����V*s��M����
�yBʚ3BZ���l�*hz>8ЗI��y�@7~"�3b��J�d�Kw�(�yB�&l��S#�F���ٖbU�yR@)e��Qń�; pyb%���y��5��zcb ?���d'�>�y�c�� � @���@�څ)��yR��$��,��jK�ᙧ�yB�O�&)zt0ڑaT��jO�yR�R�O�*pP%�E1��1�����y���6� �7I��� l���ë�y"�ךI�8 �e��)'�|y"%��y��x(�� �?]�%!�I�6�y�C�%�y�A�AA&�4�a���yF�%0�m����7 9�-I �y��5@C��s�Y�2}z����y��C�
κE���T V�B�K�IX��y2O�y����ҩ���̥��C��yҨN�|ْ5��RD���H@��yR��!-*��܋)^�`ǥ��y�&�g��5��-3	����%�yB!�bp��\�J8̭���؞�yRg� ]z�� ��-��K�'�y�@�"
lХ�4ʛ� ��ç��yrA�v(�� �ٿ=����
#�y
� �P��F3Y���v�>z-�:�"O@x1�O�l�
(3�c\X�ճ"ORP�OQ�|y~�8s��R���"O ���LF%Q��L��@M�`��"OvQ�%
��Y�f��El�a`�0�"O�h���s$F������k1��C"OD@A$�,S���S-�9)r�Ȑ"Oؠ�&�D=�Q�4�.�}x�"O�mz�c
O ��"Ko�
+e"O�ɨA���`4)2� G(=����F"O&tV��bC����4����"O�`�qƉ E��3W뛇LE4��"O��#�J9bO���� ��W4j!Y5"O8�!�?�8��'"�!*#$L3s"O�R����>|�h�g<@�(F"O�D��	W\|���kX,���"O4lb#%DO�n!��/χvE�݃"Op1�q�]*Z��(����!U2v���"O&WK
kD��C6(�A��dw�<�s���!�>}�G�b�6�p �G|�<���-�l��EܶЊ�P�	u�<A���4F�����8o���ou�<yD�`��L�5oFrZA�m�<1�,W �h$�u��Ff� @�`�<���&A���u�չ{؎��Ԉ�W�<9$'�   �`   �  "  #  .  9  �C  xN  zY  �c  !k  bq  �w    -�  w�  ��  �  G�  ��  ڮ  T�  e�  ��   `� u�	����Zv)C�'ll\�0bKz+��D������b�&D� �y���yfY$E+rT(b��L�dmb���������^L�L/6�nm[���a�Tl�;#l�M���7�~ ��'zo�s6e�,H.�ū���z�Jd��ŐkP��C�,R����;�Z$�&��.A	 O���D_h�V�cִ�"�8DJ�I v�H�cI ��'Z��
&E�ov���+`�ιq�G�O��$�O���O��r$!��	Π@c�W�j�(�(�Oz��˦�7�By��'�R�[P�O��'��	#Àg�|:S�
�o��t�F�'U��'sb�'2�'t���D�J i��t� � 3V��K�4̈i3�E֓)�ͫEo]�Q���9?���:z�d�\��o�-,�1z֏'֔��m@�3
��'��Ĕ.�'Y�xSR�f�|+��<�e`�r�Hu�CJާ =�첀@����(ߴ�?���?a��������u�EJ6��()���c��1��]��A�O��o��M;׻i�B7m�OX�o��	Jݴ?��X��M�!ڄ=��fO�Ck쀲��G�'JP|��鉴eÜ�x��!5wB�I���%)<���3w�7i�H�6RS ���+s5V�!žk�:�3UH6�M3C�iD�7�����'L}�����KU��!��Ӣ$�(H�V6v�lD�ƱX���$������Ƭi��H�;�ر�i�p6m�ͦ�)�B-*��ǯԧ�^�[����ǠE,wX�Au�y�0�oڧ�M#�B�; �8�z�0��ܺDf�?nr� ����-�6$CU`
}���J3�	"c��a���C28�&�s�"�m��F*�R�����J��U�9�9"6� �Oeh˰̌+%��IV�ȥ�M3�)C�n���#Dɒ 9D��?��B%��Le���n��C�2�5�[&R�T�^-[R�'�"�O���m�E�4=�E�[� H���6߰�j��5K¬�Ag��E.��'�btٴ�'y��'�x#Q+��~:d|���{Ӝ�]���Wiǜo�N=��C̓/�z��DR$~W���u�S�,F�pa��%F�%l�Ȋa镔vH`��	.0���5�I�=�8	�bh��vuMh�A��rD����O��4�D�Oh��<y�^j���5�ц�a�)�$? �����?�vǩh���K>Y��<ͧ��銇/�� c��#_��9�3����?�(Od������	F���y�!D8\h}P�JC_5�|1�O��?���M����V�����A��9�͙7�/��_TuA3/�6Sn�l�Gї	�H\�'����mĸt�-����>4���`�-����TE�1�.a�X��aϜM|��h�@Ⱥ�;�.�ɮ�M���|"wjC����! � �z��R����8�?Q��)��E��b�d�$)�]��C	���=a�'����h����֦-��p
L�a>���L.y"�q�I䟤�'6�Iaw�'���'�rR�t��"���`)��8�TuP ���H��(��Q4���⫉?bzHa2R>��ӵ��'ȺT)� �.�~@�X�����ƫ�rw>,���Aд�`0/B�D�^���F���Pi����p�[bGV0��,�ȹ	Z7��Lyb�5�?	�'���|�pc��� �'1��1�4�X/:��'�I�H��O0}���e�a�*D�)��i`Y���ߴ0W�v�|�O���T�< ��%w��u�ʄ�5�z�X�Q�6S�4z�O^��O����)e>��!\��rQ8T�I3H����tR'~��@ɓ�u%p����}���ی�$n�^�K�K�-�D@b'�U� ����$&M�
P���,Bל-"�W�\8�`J�l��=a�)]�BA>M�t���o��"& љ^�h��8�M���j��vK9�����zv�4#�$�.{���@��?���0>Y�g�!O���w
��z�F�t��J�I�M�g�i��I�1�l�x�O��_AXpyP+��^ 4�F�	�����O�ؠ���O���OZ@ �M��3z�(�F�?����֢ș<��:��-'h|���?X0%���D�����x��ϑT�*h�?3l9y���H���L>��b��B!L�*��0���"�	�]W`��T˦M��4�?�ak��0V�TyGрS�i8�ڹ����OV�d�O���)ȈE�X����Iў���Wy�1O��=�O�|7ퟱ��ݣa��F�N���E)�,�o�iyB�7-/�0�$�'��Q>u�`���<p)X)!�>�A�G�5��<�Af����^��`ȰI�9+>� �(�>uh�K�8�O��Q##��0t*X�3�GQs�$ 򗟌3T���:X����!\ ��(���@��CAl�?+&��4F��a��$:�h�7��W��VKt��ɍ�MԖ�D�i��Ry�5��*CB$C���1��'qҔ|b�'T�V�h�� �=w� R��D����ؓmO���O���I���I��M3�e���Õ��?~,Ly:E�͔bL�)�i���'�R�E��� G�'�r�'5�=�ܵ	Q�ڭQX���'iG ���S�@� �hy{���3M�&�`�ʛ/ch�S�?MꃔxR��}��� �P=]0��EPmAzH����>J�q��A7t��d�ŤD�Ӄ>�\䑖`wލQ��W�,���SQ�H&H�z�9�#�ަ��U�h����O�c>�D�O>��� �q��<UG(
�/�4?��D�OT�d�O��:�3}�f��UJ"�B�-�9_�yb���,���Q�ش�?3�i�"�O��Z>9���I�<�*��h�8q�`�Rcت�F�Rs���I����9�u��'���'��T��(�3<�:qk��E�����,�8sx��3��8SS� �D~bos�I��,B�.v1VI�g#�L��͕F� �{Q��s�Zp�edg�X��*�N]�OT�(�[��]�L�%P&1� K��_�G~�FDz��	�	B�*"f�s�m@�j�H ���;���Oʒ��c�L�`�(^Hd�Da.���#��+������4��dD�=8�lnZ�p͓���ã��/U��>�^pE{��'�TL�U��s<
"0�C<#2Ԍ��� �0�a�l��� �CC�q���*���JdĠ���F l�� ���K�=+@�prɓ��<]�hᚇ���#����2�'iY���VN�6˸'��MK�8���<�Qc��$��G�U%R�0�QL�	c��OB�ƈU�W�!��F��^�eB�'�d6���k��7���Bz��*� ���o�Gy��Q�v6-�O���	�Oa�F�_00���*�cT��O��$Q�~�p��l3g4���F@Q�jE�y�'H�%��6��8b��v����pj�N�@�'���`�Y;b�Is�޿,(P�i��ۊ/s��#�Z;q��[![���������,,���1'��y�@)F��7��D�a"�;o{�3��+�l�ô�	|>��D�,*@ѣIC� R�m(��?��?	v�i��6"�ć�x�Nظ$�G[�`K I��|�\m�ʟ��'� �ۦ�O+r�'l�]����#H���w*�?Q���B!.;��U�C�� �d`^,a���O{��Iņ8��']�yWb�(	*`����l4�!y���-GB��D۶CO$�V�.b��dU>��G�T:T��Q��3�(H�w��pP���Y��!m�%��DE�b(��O��3�d[�!��`�!�ț����RG�*ϸ�dD{J?��5f·v�m�b��%s"���F�O����e�޴���|�����d��V:�`� �N�~��	E�K�11p�����2����O*��O�d���?)����t��R!!51hujS�J��>)kA���%D� j�G[��J����!H�3�&EbCp09�
�Lݠ��$È$%K��!w�ʎd� �Z�*�`�'��,9�oV���@&T�w�@4A�`ؘ�?����?A���S)R�xh��Zw6��8�%<��-�I�T8v�zlƋ>�n`u�؎tfZ�O��o���'��͠Ӓ�D�OM�GK�d�<#cTr��0���O��Dt?^��O��d�P�:�؅$�@�Z�Q㊀^f�K�H/�lIPj�&"��iW�'��O�� �f��akr����C��>q�F�%Y���Cۭ %P<�V�3O��Y���AIv��{'���?i��i���!�F$�ѨQZ��(�f�0=&��D{����D72�� f�ԍu`�0��M���?�÷i��]�T�_�Ԥhkצ�(}ANA�(|�L�6����b�i���'��S� =J���`k"�"�T�h�)"D�� �)������U���'��[>�'��1	
��"��'X1!z�y�O����'��Qb�H��������P`�ٽ��=��j'm>ʵ�F���c�M�O��o�H���� *n8җ�E�N_ͱAGĊz����D{J?�AE�;+b��k20D+ç9��b���`rӖc>�l@� ��h���a
�-�t���9��۟<�	;\ap��ßT��� �	ż#UCسj,��B�e�4O��ٸ�ɘ�`YL��Hcv�P�+�\=��(O�|���ӕK�Pus �˶E�]��I .{���ч�Y-=�:�Rr#Н2�1�1OR�� \ 0�vl�\�Ua5JuӤ�'��������ȟ�'l(�0d�$�>�ʉ[��$B���=ړ����	aR�d E	_-`��w���I��M[��i��DiӢ�'�z*�������*X$�Ϲ �j�E�4�T�B����?i���?!�&����O �D�OjPl��|� ��e�&(̱9O�f�X��FD{x��F�
*	zr0�UN2BPBɪ��R(��4�eM�h����6J�ɀ��!�dc���r�X�>h���Q����k�֟Кݴ ��`�'r�I)m�̘��L�E�0G%Z*Z�D|��Ӫ@��[�^���T�w� �{��'F�7y��n��MK)����������<��*��-�I
��K!%�p9��	ݟ�'���'�)�N���aN�l!8t�`��1%�`�PM��';�5�'G@(t8䠓�e��<��%��� Vh��$
2C_�&��n��۷d��Sa��4�.���J�&1e��t��&�)eG�O2�nZ��$�-`K��[g��&q��4I�]��'ha|��I�֡2�&�Xm����.���<���4��n5-& a��KV��p����cۼ�ش����O�o�� �'���ٶ(U�:D�B(� (���B ����������$�"8F�Q��(�5P�8���<G<��u�3@�\٨WaN�pD�Q�O��3��@��8�@��~ ����λ+��px�>
����B+EtPl�֎S2���W2v�I&e.,�d���H��)������dg�yb`�|N,1������?!���?Q��I
�צuA���C�b�i�*�e��'��	꟠`�O�˓���n�[� �²�\�pw�%;e*�	�?���?��GږL��"Y��?����?���y���V:�T�sd��vF<�᥈�<p�fEC�"�9#�b�*1V���4�)�DՈH)X$) uF�r�F9\���H��j�0��#]�X,Z�aY��� t��}Y��m�u�B`3>�������pb��OJ�84z���ӟ�F{2+^��P-�E�"b�Q  �o=!��!?�t@��I0�1#Jޗp<�	�HO�I�Ox˓�B �'���.
�n�at⚴a� *��Sc����O���O��	�O�$r>S�"5�jU��N5����A��R��C�I���� ��OFP9$4P���TgF�@O ��bψ'@p|1���@�4Ͱ���ĕ�FV��5�OBH��j!kp�%l�m׬���"O0qQ-��'y�5�6�A\ʸu�|��pӺ�O X�b���E�'�>�Qb�����իF�]a������Ot�Dc>��c;D��u���ZB��(���(>7�!Z"�S9Mg0)����Z���`%S8�Q��J�I wG§Z�j�$�Zc�V
&�s�$�1���Pa��+z���\�P �ԲORT��!Q ��DDզ�X)Ot=3��4%�h]J���
#(��u�|��b�RD��$%�_���6��;�έ�?i��4�(�n�/�9�0�߻$�T�*�:Y- h�۴��ؾ���n����	}�Ĉ�����&��<"�*�Voi�0�B<^�"�'�f���h�h'=_&P���i��x�4�׻gd��� 	d�a�S��k�I{��s�ީ=P�d*Bu�OOh}�eϋ1L�Xr��X1\����O���$�'P67mV�Oz�iЂvrn���.?{x���3`C�yr��&}���M1=Ę���k��d%��?y��i��7�)�(O=ZY#�*ٲ@~:@Ub>k���o�(�������.�13�`��Iן���۟��;	d�Iأ����@�@H���Cd֙��h"����5 0��P̧#�l�i���P �ӯg�rX��'�R�l���0��MEjͼ�#%�B7M�@Ց1�~�lXZ��λ�"E�`�:t��˦~H�ٴd剷t���$��g�I�x�YP��C�e�x�[3	�:�T��OQ�Ef���[E4�a��82ȕ'�"=�'�?1+O]
��K��H���;604��P�E�c�O0���O.���˺����?1�Os�ŉ'fܚ/;�"$��j �s鉛4-�х?pG�#�	�P"?��.�Y����*�x!Ȱ���za8ԈPC�=\��1k�Y�?��0��15�	ʖ�4�I�� %G��?lf1�K�U�X�s*�O��D�O��\G�Ԥ�
���Ud����3��
5�yb��*,E@�O�g|�!�
U������'f剝4�����8�D�BX���v���VZ&��sA�/6\�d�O�аv��O���i>��U�]w�<�� �X)GC��'�r�@�H�3_��rP�?9P�A��D̒|�DI�u���EW�xȁ t���Ȟ��T;����t4����@�!�
��3��)�'��Б�FH���<Q'�ܝ|�MQ#Go��U��ÄF�	ן��	�c�(d!�⛘b襩�$��.H��d�ן8��Y�����q%�>e����fd�OJ˓"�5v�i�r�'~��i����	0~Ј�Q"�5\<�e#��$l�$����C7%�EH�q��?H`�(�B��+k[��#2�#� I�ȸ��aI�mR)�T�	\~R"�R��$*S�J�j��Pr��C�,��ʂ6?����v�p�����]��]z0�UH+�<�'�����?Ɋ��y��Hա� ;c��%���>pࡳ�b<D�P"&�� �B"J�ax���(9���>qC<7�F�+d%Ӊ1��	F��O����O�d�	J����Of�$�OF��t��Ar��=+�X��С��3�����4am�яܡ:q(0x���6��b>�AH<�­ήΜ�b0 ��1�����f8+"�;4b�����%$����� ��S�29H�Z�w2Th�9=� ��G�?ք�������<\�'/ў�贈O�I�:�fᜄ#��8��o�<���'r�Ac�F��
}���Zky�b"��|b���P�e�횱�H�P�R �2�H��̟$����O�d�O����Od��m>	Ҷ���]��@"�۪�<���8s��V�R4�V�b,��>��4
�����`��]ȧ��*V���p͙�U���\UѦ�k0�Vm;&h܈.i*��VJ�"��'��d���uJ��;7ĝ�� oZB���'12�Ih�'����)�}������/t����	�'��q�	�W�<DR��֐ l�P9J>�0�i@�U��B�,Z�����O��#�V0o�\��K���p�B�L�OH�$ڤb�����O��S�Xwp�[u	�؀d#�N@�bM��iv�-��
&Nrr�qGf���O(��� �+Q��! � "�,�a
8C�J���J�$-���Ɩ��|2T�J��F�K�{�O	�?q�����\	V����e���8�@2O^e��'�a|r��.$�\{���KX�5��� ��?��~�v��Q��*vA�36������'H�ɂ;"���ڟ<��W���H�wf��F?$���z^"���(ʏd��i��?ae�G�e�~|8U�ELX"���ۨb�h�r���ñQi�%ȃ�уI4@��&����=��8��A��(�9��A�2,�o���!��ӟj���Q�h�.�e�چ{������@�!��OZ�� ڧ�y"DӇX��;c��[?��<�̅ȓ+P<my������y叕�d
EB
:ڧ��Tsqb�̙I'��2���	���Iޟ��dIF�a��d��ş��̟��;{=x5A� D�������-����"��aD)�R�G����2�Ţ'��'��-�a�I���:�'�'A��TRBo^�'�Fd+C-�;WGB��d*��(�B᤟��n]��J�=� p0w��/�B��6,ޔ��ِ�'���=(-����O�=�s!�
,�>pi��^�F0Z����y�b�Cn�33(��l��� ��$_�����'��I.ON��*Pʑ%�T-��G.�����͆`�m�	���Iٟ����D���|J3A�7L���7$8I��+DHٻC�Vi����2Ic�T2S�-p�LJ�i�� �A�nz�x�Ǝ8I�p�+��R�l7"�r��C48�����D��	�VD̫~>���{R�U?��d���ÉlYN%�t*���Ѐ��?i���)$�ApFŜEa��u@/#[���\6��9uL�/,� }���JA�ɞ�M;�����(����O�21��Y�c 8�TPRa`�&���'�����'r?��*0n�.���b��=���r i�*�}��`����$(�oD4D��dD~B^�3,�=x&#�DOz�" �!9�\3��|$�C�#�?o��(u�5Z���`T�lܓL�n���ߟ �'�*�1���}�j,�q���t�t<�L>�	�_5���aG/|扨`	�4�꽅�	��?�S��c
�C!�	����d�͟��'�R�)p�'7B�'���;|���@yta��h�i��8XD�(V ���	ΟX4��r�*8S v4�����^��)4��=g~�)7���I�����lKK~R�C�5���3�],�����(T���.�|��'PI��S�D�0�.<���?$ ��'�]`��?����d�H��dW5����EJ�2j��Э!D�4���S�qAP,�T� 9y�.�B�G=��0j�>��`-�3)T�Բ��9hLXPkVC�O �$�O~���V|ܥ3���O���OL�Dh�� �'T�*\�Te�4B����\�G��#���~9��  ��:,c>iK<�`k�� A�N"w�t��v)N�9v����͓ e4����Y/`�DH�Cb?��k��g��E1�wK6L�Ĝ)D(�1���wH����d/
���'�ў��f#�i�8���	/`~��r��l�<���V�"j�U
2�N�sK�-���Ny��7��|b����*�b�Y� �(�z�9gfG�WLR���\� �����IΟ��ܟ��	�|j������Ӵiח<T��0�.�mi$�A���#~�����
�1�
Ԫ��	J���+!�Y�%U�y��Ph���VBg	uM_0w6�R�F,8���*���i�6���{2	�4@�\|AԨ#]��Q
�Vu�X��?q���1�4��A��ڐF�,<8��٫	�ȓ?7z�aF��7M
��Go���\d&�T ش�?!�Ox��V �~�1.���%KN�q� Ah É� �X���?y�B]��?a����$�C>E�xc��<���ض�D�i�j�Д^�(0@�T�� ZT�!H*������l��q��Й�F�s3��3ӭ$X61hd艤x�5�W�
�ʈ[�v�x➰قn�O�d;?1�
��	�|ա�Уm���F�Ic�tyT�3W(5B2O?hq�B�"�Oԉ���O{� �!�	(l�̓����`N���<�ǥ��?����?�)�pH�5��O�@ْI�
"vQ�Jm����O��d-�F]����)|D�KǓ,N���O��j���Ic(JE[b��$��2��"�^`k$O�>E�d0������n˰H���q��?ec����Nx����F�&�(���J-?Q��ş�	�Oh󄝹$����b�C�i�a�F�<_!��P�e��a+�H�?L�n��GO1Vџl؈�)O� P� k_=�L��"dʱ@R�'�"�'t��!���6�'�B�'P�.��(x��I�H�fa"6�N�f*��y�	�,���7�$X�6iW�i�}�ɫTW�Y�E�H��(a��I��$K�m�p�Ĭ�9|��������m$�'D����`E[ʼ/Z9��hDϸ!���D�A���'DhI����?9�����"��Ș�fv�M���ߧ5bC��Q��}9�!Q	x����*>˓=y���S�ԗ'����-�#O���{�jҚF3��H��*m�Л�'���'��O�R�',�I_��E�7�� \M�Z)�)����j�⁋�&̾H�j���B5�[P@�"0�B� N�H��)`*[�$K=�ȁ!��U� ;�bL�Mp�Y�Æ�( �➰�a��o���@mތ��9�AeJ
nJ�D�O��=	��$�ވ�aĥùH��x���:�!������YGj@U��8�A˟?��'�l6m�O�p���eS?)�	�gD@i�D�ԧVE��	���<)#"���H�#�ݟ��	�|�I�Q�d8�À�O�)BE䘆sܱk6M��>����` �4���/$8�m��i}B��0��D�Ĳ�hX	);ԙ+ʊ�7�Q1��G�;�`��d%��'�L�x���?)�Oڽ��ַ?���-��+���8d��'�a|��	q��*bi�8Ec�uk�#�'��?YV�'��$�I�!����cڙä=�����$L��$�O��$�|�u � �?�W���!���cMh%{`)H��?�&ђ1r%B[�0��d�D����aR^?9�OȄ\�g��@,��;s$YNW�e�O���� ũ �b�V(�?���[�Gh$���%��$+ŘFm��:ƩEzU\)"�Ə��d��(�b�'@�>��S�? �y1�h�x��غqh��
��	�"Ol�	��P�l~Z�Q5�D50��Q���!�h�J�A2��y���5Ӝ|��}cd�'B"�'l2A�N�h(��'�2�'b;���/A1����兰`o  (�\(�r@[�e�.^6��e����1���OV�Z�`-HʁKV��	Sg�ұ�I�1hda��G8We� ��g�4@�\�J?�@"�8nh�ݧ*�L���O`�x1�d��r��'?�R����,�IC�'>|Ӧ�͵@,�� Х��s�:izW"O��rU�� �� ��*� G�m�uU��Q��4�X��<��e��^h��΅�EWz���!Э'���+����?����?��������?y�O�PD��֦M��h!��<�lM#��sw��7̉�`����P�-0�џ�����0|�Ef�͈6b��&ݶ1�Fy��똕H	�  'k��s/Z+K�f���DU�d���P`�B�s�b��O 8����C�'"�I`�'a�|a�5.�T�w"@!w(�ȡ
�'�x y�ǋ�$�f9���4k^��<qg�i�BU�*uF�?����O`1���ʜ *�u��7k�&I �e�O��$Id����O���^@ءBDQ.{���a6���Z�<9e�!R��:�Gq�e!2��J�'����-Y�^6��b���LNŻ�O�3r��Sq�L�Z~�I��f�1�����F� /f(X�=Q�g�ߟ�IQ~�ǉ�A�Ȃ���T�A����0>�C�XB�j0@qb;2<-	� �K��D�|��ip�c�*ڌ�㠯X�q�|���@y��j-��' BQ>E:j�ɟ\xU���6�B��w��^2�trsl�ƟX�I	T�楒���<���|M�)�e�g�ę?�!pgD<~���r(��KK��2 ?!�b�`��xgW�h<4�įWHC���v	G�r# ��'mP���L�Ex����lȚ|�$�U���Iܟ�D�1O����k�����RFCW�;� ���"Oԥ�W��=S4pQ1�g�l�������&�h��E0���1Whpr�ʬ\��Z��'�R�'�2lЋv5t�YS�'B��'��9��x�?s6Ƅ��í4t� S�R�C\�Az��@�J*X`�С�"�1���O�0(쁰+F� ��^p��@��V�ܸ�23)�@��Ͳ%D��L?�(�,��e8�杻Qzy�"J�;$x �j�:7V��d6?pJ�쟼��`�'���Ш0n�^��+�m�p�G"O|ň���1|�9�@��O�p���\�ڍ�4��Ľ<��d�K�t� �Rj�	an��tOJ!ʴbK�_3"��&ǘ�"Q��D�U�����C�QdF�9��P���i��G̽��2I��Qb¢��?�����?���?1���%��	
��#u��"����g����]��JW #8�I�FغV��">!G�֢w�J�Q�O>�(r��m܄A�Ƅ ���S���l�.x�,A�%�����#�	�MG��D�Ob>��"���?���ӌ��pm�$��<�
�z.�(ض%�#O��m�&N`��B�1��ɱ<����G�����ܼ~�ʓw��:��?)���i��d��D�O���b�;��1`��Ɖ,�`�١��Ov�J"��q����X�+:@
4D���d�i2]^D����\�-/����O-��D��t�d�Y�l���Z*k7�9�ĠR[hU8L?)@�f��d?�� A�G�h��9c3�v��S�c�OT�$,?%?��'9�QA2Đ`��U�so��K� E��'��( ��6)���!�K������LN�O�����A"��%��U�����'���'�ݺ'"�����'�B�'����'��	� �������#(�(Q��;(؁�ϙU����Ȇ6�����'��d�t�TR.�sd� &���ʡ�xH�c,�6>���(�@*1�O�|:࢑�����v|�:�O�TMhE��	˜��'�����?���g��2Fa
�� ȥK(B��*e D�|`�,%nT%�&E�B�r�K�O|�Ez�O�RS�\�G^m��1��
Y�@��C�T�aPw��ߟ��Iԟ@�	�?���ʟ�̧8;:u2`	�:�5iPH�~&���\8%K���0�P��h~��L���	:���H�`A�>��d���9��Q�@bY�}>��@j�t.���i�	W~QI��L�+��H��=
4)��`4X�)�.=�b�	Y�'��<�d� .*�Y*w�7=3���'ʊ0�Wb�9p��س�e�>&U�*O> l���D�'�4�c� �~�����tkʊwäAb �M�;�|��ʱ�?r U'�?����?�r��h��rc�ɉ"W��C��*�h֝�L����@�E�W�(T��F��x#>Qf�X-u�	�]�\����\5z�`�Bv���E[��An�0��� �]��yS�b?�	/R����Oc>� �N��0�hv ��<]@ u��<��j����g�j"�;'	�f�ܱ��I���Č�: VIf��P��Ub�nS"A�IC���������O�D!��Y�E�	}��]	R��~�Υju�	�/�Y�ɑ����$�رe7��F�<|�v������� �RN�eF�<�X�b�Ǖ�/��=[ݖx� O	'���qfL�d'2�f�
�"�8�H?��L@�oz�Ȳ��U:2�*mȤGy��ᦧ�Ot�d ?%?]槀 �P� �rI$�iB�^�@&���q"OJ���J � �zv�Bs��g�I�ȟ��8���pŊ�1��,ZW6��@�O��D�O�Ԡ��1���OJ���O�i�O��ID�C%��Rwhĵf{���,ÇrD�Xa��$q���ń ���'~��O
l;cC�'�b=��{��[�#ͭ#~.�C��1k���i�\)?N�S8P֦���¡k�d��x0�"������CN��G����	��LE{5O�zt���T�B�N�=���"O�7lk��$�bʥa����'<�#=�'�?�)O��1]�����#5�!��&	t���ԫ��"�'�'���'/27�L� ���ȉ��b��ݪ�d��O��X�	�)���2�E~��F0I�X\��փ7,[T�0d�$1����B�����F̺aЈ�
e��Xm���RR�F��H�	�?i^�A��M>d������"`֍�	|�'��(��),�|�V�"zՖP�2�7D�����
Uƭ�\tx�2�]�z��	�Mk���d˝yP�OY2:���
S�$�F��� 0�m� �'�&y���'	�'�P �R��1>����4>m�#�㟲xxƭF3��i�7�Ƚ{3$��5�I�8�ji�ad�$]�����K�r�F����U82f��gȪN���R��0|�DI"S��#H�qO*��@�'rb�i��4�l��KW[��h����F���l��D�6bYp��9h iƈ\����� �O>�'(�a��i<nP�U 0�G��\�/O��D�O����O��ĺ|2���TbG&P�����}�DsQF��ONUF�4���2�PBw%��(Л@� ���'��L<F��O$�7�Y�ԍ
�)l:PQ�|dh'�i�*��d���'E���'��R3x�ݨoC�n������P��pӘ�dP0v����`� �Y����u��?λe󨈀qN�Y��c��K�l=�4{&��O��d_>8����K��?���?ٛ'-�ْ �K�(��� ��g	.Ha���?a���u��.��������fd��SB!A�OY�-hƩ֝:ע�ÓjS�äE�OX�ě�?�8a�	����?9�'�jPl&&"�����҆Td�@�_/{���	�d�����O�e�g��O���ɪO��s��ГG�I	I|@�p�;�H9í�6%x�m�<1�c��0���"�H�'�?����ze �0c[�Ų0�56օ���8PQF��'�
����?����Db��8'&��?�m�0-�j\xP�ҫS�X��j˾+׼�"����M[e�' Lm)��?�� ӬW����\�	��� ��.[L\���W�M8|p�4�l0�'���Ѻi�*6m�R�dş��ѣ[�?y�3�ƛv�}�gg��蝎h��6��q�yn��?q�4Ul���i��ɤ~R�'j�IK��X�b��b�g�Q�ԤI�"OJ�U�+N�h��؝*�����i�R�'_B�'J �'�?!����i9$8h�,��hxbQHfL�Q۴�?i��?y���?���?Q���?��O�ٳ�h�882,��O�A�xQ�۴�?q/O$�$�O��$�O����|
gc
�T�R��g	r�y��$O�\�V�'���'��'���'x�>1��22.5�EA�a)��aE����3<O��'������~>P<;��	#x@i�4�?a����$�<�H>�'Q����䘌[k��4��"^��ܴ�?1*O�����?9�OA�\" jۍF$(�@O��ƍ��'ƌ:��Y>o�D��
�l
� �'8>���g�T}�h��&* ��'���0$.u&��'		G�l�'M���A[6�t�sv(_}^��'S"�;c-߰H�`5�u��5G"zpb���p�R��Õ�U�$3SMƹD��xi'��Jr��"ʧ:� ���.|x�
aJ�6FN�K��'�O�<����H,���EV_&x
��ě���5A�Ȗ�c�:}�0ǐ�bp))�(_*�DI���@�5&����ΠWzl(XE@�.�&��#2��\��F��=�J1�M�N�a�P���k�ș�B�%���1NQ!c*����iU&mA�4X�!ܯ�$Yʖ���[d�4=��4���A�ƽ��K��Z���R�Od�h)�4R�iI�"ei��#v4�"%�'�B�Y�^r�T>�,W�<U	T|��� ���u�E&� (��;�S�N	~H����'��@�ƪ��h�\u$�$� M�OP�&�b?�i�@X#n����N�,D�h��"D�\3b�� VXY�d�?B~48���?O� Fy�o�$a1��S�W�d��Kg ��
�fIn��<�	͟�ZQ.߁s�x����D����L�#�$�tÞqY��7��5G=�P�<��,�lX���`;%���3	�H���@9��G����d�46�`��m��51#T#P��K>	c���>O(��lD�_8��9pc3G�E�"O�!a-ʬE��dC֢@��Z ��>1q�i>1'��25	Ѡ5��h"�׏w�|�{�l�.w��K��å�?���?���:����O��Di>y�%�)��-jG ǓP_��e��/<�C�	��� ����ǔy�C��r��PB\s<���ijt�����Era(t�܁@��I%�p?AFZ�@6�՚�jY�NG�"Va�h�<���Z���ȳg�6F��)@�TJܓ\2�V�|"���f6��Oh6�� (~x��R��*i��f%�:Y4ڑ���01a�Ο��	�|��F��$��*P�P ��s�J�0;K`�q�",O`�R����fsx�Hu&P#-��8��/�;Yay�jL��?1�>�P��!�:�X��2uV$@���}�<q���s%.�ↁ�+"t���m�}(<�tAݶY�҉� ��6*@IjT#�7�xm�M>����I˟��O����i�����X%L�<Ӕ�1����m�ON��J#t���.�$v�U�׭^�)r��O~��q<�\Xs-�W��H+K�kp6O����̛���o��p�B�FػAX�	�"cT�tH���������Ѐ��B6 ���E)�ēu�l��	��MK��iT��~J�O�J}� M�>1Ӗ˒ TW�<S�'f�	韨���D�'��V�����P�xØ Y�
Ť%�P������Z�6���|r�S�Ж'���`��F�8��
?>�#ƓCP��nZʟX��֟S���;jE0������I��L���l4SR�A�~R����;P��Z�$Ա4ay���B�*�cjw��-i�L����'Ąr˓8."�a���2�4h��Z��P�cJ0�$Z���L<���
/����4�K8/C�ۡ:^!�ֻ�4qSwj٬h��![�eZ��&.���Sr��(Gr9�6Y�W���9�����
g�� 7�d�r���?����?����?����Fͷ&A�5�0z��I�M[qt����'^�m��`��Av�:��շ0�^H��bō�x���~R]�C�!Y<��OB|E�+����~��W�^�4�C@\2+�)��H��y�^)4όȺ7��9$r�U#F�#��'T6m(��E�<t��lП<o��(h!3�J;����0℡pܪA	��?�f���?a��?1C��]��pc䄩T�d��N>8��[�F[�Y��oZ0LkҧW�-V6#?9�K�Q��QGW����!��Ҝ&8"Uҳ�X�5�E˖�˅��@��if����έQ��'d����3��v�{�6-�y#"i��I
�a���`�X�8��P�'��'��'���'\�i`��e�hZ��m`s8��$��o�j�I������?y�׷x��u���ͩU?4���%�p|�����J
�\n���0�	����=qB��o�!���ń_M�8A-�d:^|A��?�� ��#�<I@�f����|B���D
�%K���0&�:N����x��A=G�*����zmQ?��"�i���z�N	���]i��)��RN'��IǾ#��Ц&�8:|jCf�xW!�$[�^�
��ƀ���򪔀"���F{�O�<��R�L3n��U�W�O�Nݱ���b�87��OP��O	�����~��O(���O�Ǌ�0�8ek���X|.��!��0d�b�)]�~�i�Ꮱwu�X9��|��'���n�`�L�$D>�[l1R�T�IR�O0��(xAf]&W�Dc��E�!��X�K?�)�l���yDF=2,Z%Ib
X���pq���AD�o���k����?9��M����|]�� O����p����'B�'�Ҙ�L>!�F�K�h 䀄$��l��{��Ϧ��ڴ�?yD�i���O���Y?��V�IV�|�2����,��}�r�����	IQ��'�b�'J���'������S�&f"쑠HQ�k��H��!D��Lt�X���Kr��d]�~���<1�A lԬ���̏9�@co��D ������L�*�.۱/�r�c'�u�v���N4�I}JP�ېH�&Z��iVp]c�d�OLln>�ē�?i����'�\�z���R�2����ē+|���'�a����F��������8�!�_Y��O�l�(�M3.O�Z�I}�i�f؛HH����Cn�4g�
r�O��DC
	����O��dȶ%��4��+N/^cΥkq�$i�U{0bJvZd0�r.�B��m�.��OTl��DO贁�l][��-@�J��rx��bC�ޔ���"J��F�h���7\�\��{�囈�?���i3�6Mu�2��ήt�\ᚶ$�<3��yb"SSy��'��O��?�8��h�劣f5p�����	���CC@���̝)Y�}"��[�cΰZ ĕ��M�'P�eۥNp�H�D�O�'&��4)ݴ7�Ԣ�oD;:p��te�/6Ht��'���ϓy3�1c�"�plpÇ�C�����i��r���.$4Q�h� B^�'��I��ߔ6����'(�,Db��cM�&~�YqO�:r�Ln�4��ДC�+r���B'�+�ćW�&<��	�>R�M�iשjW(YS�<.!�$�8�*� %*�jV�Թc
9$��xbl+�DCBy{�k�ql�l�6�B�G�zF�>����?��	�OuH�����?���?�}������h��ł=8��E16���U��(�BBg*�`��Ts0��'��@�>���vEp��`,���2��Ӎ_+-�$��?�����<�صB����S^���=� fe�#,E�1�֨2���;Q�ԐYql��M#ֲi�2n�$5Y��,O7��:�|\��.hhXA37� 'z��5��{��dX�p0�`����}�S��T��K�& }��j��o�ٟ�ش�?��������(��U�a����� ��h�/M�/��E���Iȟ��	>�u��'}4�� Qb\�R��Y��+�y��)p���=sD�u*DM��<�@P�T��òdF~BJ#7�l\��|�1A#�2۸�KsH�'|����W	W�	h@K8�܋�𤜗;��E�㤉�'�z�cŹL�i���'Ƽ���+
q���Z�9f�0��D�`!�DǛi������4OZ�{T�Q $qO�m@�I%�^$����6�R����c��$LG��Q��.`�*Q�	��<3� ���	�|�7�(EP@(�RL�[�j�cÉ�9 ��̹׃6����C\<��b���ORԣ<i�
 ����������X�
�:^sF�a*�%�F�a��_$��(�6GH�-�ޢ<������IV}B��`�������R*~����'���'Ş�@%B�$��8�D>�J�'0����e�"|��8 ���l� � �[�N^�]�$p���M����?Q-���Z �jӖ�����;��z��өI�Pe	韸��)d����M�S�,O��ȃO���0iҎ�OH��у�x�@�O��h|�`��L�ĸ1t���> N�8@�xhV5�?�E�|���c�-2l 1Wg��RKA��GS,�yR�_��Թ�$M��A��#���p<��	�4��J�ԙ)cb���$��lU)�3�iC��'vB����H%�'Y"�'T�;g.@�01�77F��`�Uy�	r�X��ɓ�Y��b���x��I�O���s�,B�b������ىR�מږ��#Rz:���#<�A�LT.��O�($��z�!��焜Fl�dj�ϴ��I|k�'�"�S�g�#M\M:P�ͪ1l�їH��U�:C�	49]~�*W!#��آ��S4$t��'��"=ͧ�ē0Nt�I��Q'~�E�'��S��!:�𝋷�'Q�'ub�q�A��֟DΧ5�>�g�\23��i� B���x˥hN�y�����ׯ=LFp��Z���	1��;M���T;hФ�ŦX�����+0�͈� elD�>1�kʳX{�As�78�x�{r����$�	��p?��*��2�-y��X������o�T�<1�e��I�@��� An���#!EeܓH��6�|�'�2��M���J���I/ゴ�#��I	r�'A4+��'��'���K$��4��x�d@�{i*�)sFݷ/>D��Ν�{�8a�E���F~�e<N��lR�k�(�z�qS�:�T`Ǖ2����o�7͘x�n�-@q��(����'��'p�����P���'m�
6-�{�4��;n��Q
�g��'�쩉�Z�l�'����$���m8�ȥP�^y&0�hǂU�qO6m<*b���"�d�O&�:�l��N��	B�'�[��Y����6�D�Ľ<���#'�f�'�"�'��4O�b.���޲ 'R4@�����$CD�lq��'Ҏ3�����"����1��,v�����i�:p�������	RbC�5V�'X�%��"�;~�1D���F�"x*A�ަ(�ԭj��]&j���@f
4~���u�,s�O�5���'�6�d�j�ӿw� ���Y��-�a'_G���(�	o����v��0n���8�ʟ���O����D]���4�?���i��H�T�A��67<\�[���<9�عl�ޟ�I۟�c��m�0��	ݟ8��՟��1+Bh���̾ĕqu,A�T�8e��$�?�,x
��RW�V� ��1��)V��?��K�'r	�a�$D����*�d�Q!g��w�%JB	���m��S9	s���w��897-� p����ȖI�Ұ���\W�	�K�����xB+�1"`=����h؍r�E��y2�6g�☈���2p�d�D�&�􉔚HO�)�䁊*��Ȝ�gc��z�bP$!�Т��6��]�I���	ϟ��Xw�2�'��C!|�nLS��N���%ɒ�b@����K6��A��G�m��9(fc�J�n�R��N6"��q�e
ӷD�,��/��?lLH	U5{�2D^(\����dJ����^+v�1O����P=0�����%)Pܜ��ƁjҨ;�O�:�-�E�`����EHx�6"O��g�Ĉ2�(@�pƈ�M3U�)�I��M;M>1p+Յg����'�V�O�E!��)C��F�c���$�OV��7I�O���g>�P��	�M�
"�Հ+��x�ǫ��,H��%�

Ԗ�rG f���GBL��x��#e�ψ^�D��Qi��{L�E��
�y �XD#�'R�9���5(P�d�I��>@.�Ǌ�8�����+�!���	g�n���ދ1���w$����[S�m�q�Q�4�h��l��ݜY�8��M7r�]m����IR�$G�˛�-�7Q�j�RB˟3s�8��৑, �V���O�%J��
<^�Q���ұ�O�c�D뙁��p�W�W�H�{��$��]��k�˓z:��:sf��(��9�A�T�ѓt����t �xRi�)�?�2�|��� ��rT���,}X ��!��-�2"O��3��N�vLt����2��ڢ�'�$�<Qd�ǵ})R�F�ja����R�|6��Or�d�O���H��V��D�O�d�O���I�\H(7�'Y�NX��V5hJ@�O<�F�]�j�v��|&�0�wNT�n�j�KU�R�hE�WI]��!9&[�����R�����)�2ѥ-]}D
eRFH�e7��@1���	e1��L<YԤ��#)t���"��zg64x���o�<���
,�40$#ܟ�xh��'@e���G�����x�	ԡZ���Ђ��0b��`K�O��y�>Њ�×u���O����O�����?Q���tN�.rBH!�fd�#t[��SG�
��![��_ vi;�B�5]�`���I�U{LB�m��X���dP9-n����`�?��D�t*Vm�)B�A�s�'�XR�.�=� )$F��r!���ħ���?���?���I�"�d�#A&@W���c�J�D!��:Y"�����_L�8���7W�qOb�mZ��ė'gc�c�~�޴d�B�0�P�bv	���2\ �J�'���_}��'��ɚ�[E&U�6+�:2>�K͙/S������;x�p�fœs���R!C6��B�1RG^|6��ʚ1�6��ҏ#?��,��k�=K���q�Z�����*�hÀc�O��ľ>��T�îER֎�>N�,s�Ci��?q	˓G:�spŏ{�̕kw��)t��)�b�虪�`^�l�Z#
[az�)�?�(O��C� �����'G�ӗ_lV�o�pT���eS�DU�i+C��.�h���?�d��q�����A#&j�#]3|9�F���� ��J�ʕo���zУ]��ē"�&i�6���-ʭ�l۶=Ӌ��T�r�0��钛c�����Y��ē4�������E��i=P�)�C�+�P@B�Ǎ�umi��5$��r���4�
ݐ�iԑ(��Ur5�4O,�Ey�Hq�N9���K�C����gcH�~Ծ�m�����֟��wԆ���	ß@����N��oo��X"Ǟks�Y[c���,�a����0��@�-*ux��F�m�'���$3�z�&g(+؎t����=��JЮ�W* 2p�F�+7��83�8	�����R�ټ�"@ҍ�\q�K�)��)T�׌)�B��(�S��O�)�Otc�l�qM����7IT�@Ξ� �%D�؉ ��y,j��JԚ>��#ԡ&}��+��|�����ĕ�4& �ai��P(<d��ˌ`F\�A󫅪#�<|��ʟ��I؟X�Yw�'V���d�!���\��X`�#`���"F��	r �8Ӯ��"_p0�NƵR����$ق17�$(�_�&��uPӭS�7zB@ss��e/6U(@�S���������SҔ)���M)gT٣#(�9z6�A0���n���'
�����j�>�A�]�>zQQ%�(�!��ыw���"�K#n��k@\�qO lT�ɫw��y8�4�?�شg���1س���!5�T���`G*wϤ���O̓�,�Ob�Dv>��0��<��(rKd�LqÀ살L'䡑 �:�=�mDG�Đ�d�=]@�<�!�#�X�0�o�w�(۔D��w�|�B x�>Q����./��`R��۝5Fآ<a#��ܟpJ�X��0\ϾQ�hV*l���v�=D���@�D�p�ܤ�C�ϱ5GLű�O0���c�2CV�X'R8CkP��Cj��E�ܴ$�h�&fK��M;��?-����5�d�F)����=*�<-5,Y�f��,l��X�Ɇr�J5h6I΢�F��[<�<�9�
UR�x(�Ox��#��7<����O/'I���M<1�+^(�h���ÞM�ҽB��Gr�8,��Dj�,p��pM��GƆ�?~*}���Q�h��4%�H� ��O*D%�b?9�jӾod:I� �c�̫�O5D�h9b Y��F�J���E�L<��E.O�uDy��
�w��Z1�1��,[8E�\4o�ß��I럄�%�#\s8�	ӟ4�I������lۘu#���>0�n�K��ǜ(?������t*U:�H��U�d���c�p�'g��\�2��Oj��cjίX6��+ć�#Q�|)�ҕ�vh��$q|2�4h�&<��>�k'MD��y���M:��5"�9��)�A��)/]μ$�4�Ad�Oq��'m��) @ǙK��D�w��!IZb��
�'���BP H�?
�ݾ73�:I����4��Oޡ���Ʈ
L�	�Y�j5�S�ݣV��l cCП �	۟|��)�u��'B�0����Z�DԒw��l�<�� ���
u�СD�H%]򨰁�,?<O.l � X>��A��C�>@��#ciNto�I� ��3k>���5<O�Y�$��?��):�d��L,�q���J$�B8�O���d-�!(zЋ����)n�\ke"Ohh`ȔI�P���`�,�4u�F�d��q%�,p�$֏�M����M+��"x�����ڊXC&0q��B~��'�BE��'��1�-�#�'I�':q�ɇ9�.�Js��*6�DA�
˓Pg���>I��!>lS��t�J ̀tX�����O���O����ε9`j�jA@�2ul�mK"O� .� B���'�z��d�����
O��"tÉ�x~���Do�d��n��7��O�s�K�Ȧ�	۟��O���A�i���F�/Dq� ��FH�Г���O����&>X6�	I�N�Ȳ��7_`������'B庰��*f)��A����$� +S����N��\~ʨq��xܧb�	� �2bء�5��:Nxe%��c��O�&�b?ebB��g(���D.�8Fv����%D�l�a�\#��!ԋ8}A\�J@�%O�pGyb�=�u�3�޻6��	�#\5����'�"�'��e05A�]���'����Ò�3ْd�V��2I��!p��(�H��e����	w�P��|�?IF�R�%�<��T���x���;�F�wn	���3J�^ 0���=G�}�~*5����^"k'(���8OQ��Y���@t���$yt���Y��o�-)@�Y��ފY�RPWAѧb! �r��?��dI�f�����^)9p�Ob�n��MI>9�'��O�(D�D	d�ft�d�7~����ȢA�H�	G���O��L��ۉO�jlQ�Ņ)l� J�'������_�'M��n�(�pZ�'7`u���6W��UQA�����'pX\���<N��� ���|8���'���D@�F"�YG�Nt��Z�'B��P$'�K1h �CŚq�  B
�'�:��5i�18$���C�m�~�y
�'7&�u�[7��1�e�\5��=�	�'�j*fă<�@E��L�A����'���%�дI��'*z�c�'7^t��h�y\��3��j-)�'|����f�@�9���r��-��'��3E��pRq�O|�N�)	�'�2���!�Ҵ��Ðm\
�J�'{vມ��R����g��� 
�'�ᙗa��'7>�x+[�,%�XP�'�X8	��|�s��Y�����'0CU'��v�`��˔cĸE��'$�=B�\-5>p�( ���_y����'���ʑ�#B�e{�k' EJ ��')��Za�2y~��i��K"&@h��'r8��
�!(_��r����@�p	�'�n��B�/�BXC��:z���'O�P"#5|�Ѱ�&�5\��	�'����bN��X�4��KQ	&�0�'%ܭ'g�*c�r�C�HȐz�'6���g��)�(�Jt�P�	+�� �'R&�� '�5��8��Akc����'�	��T5IU���0e���`İ�'�N�b�b
1M�+��Q�'��T#��K�lF��`	bL�c
�'0��$EϒZE�<��_�sȉ 
�'���1ɚ-Ksb!&�T)~:�-q	�'����"c�U�|�`
�o8N��'D4��
<+�!kp�̆c�Z�R�'��JDI�&��%r��c;����'���$�]g�Lx���X�Y,��)�'J2�I
K4}B����Xi
�'��=Bp
G?Nx�XqeS
s�6X�	�'�����a�(T�f��a�͓eIܽR�'rP�EGTS��(5�m��'z�����)�葓⭂<	��y�'m(��r� �O�~-���6T/L��	�'��Q��D��`k��reȋ�����'�Myl�
�ֵ��kĭ,j��'��}�����'h��9�l�8S�!��'S�=µb� �rM�g��)bdE;D�Ly�+/3�5R2"���e�-D��0�D�c��+dmլoFt��)D�3`c	�U����A�5�:,H�O(D�� ���t������I�n@�$6|��"OF���mT� �8��X�\kN��"O0���+��
6p�Cj�.f􀃗"O�8�e�v^]�R+�q/�ذ`"O$��E��1;��|c"R%{D\;"O��3�'�	P@)D)q;�9�"O\�@7C�^ؒ(D*w-�0�'"O �9� �'U2bxⶦْXq�U�"O��ϒv К~z.�:͏,�yR?.{�-0E�Q��ɨ�g9+6!�J�1����3�Ј=�T�ia�'9�!�D�!d��]㇮�2��m�1��NX!�䙭.Ƹ��F�D�y�Q� �p!�Dհ 0�I�ɍ��BU)��!�D M� @D��`�����J�;�!�D'_D��0V�+�� �N�]�!�D��%zb�j�L������LW�u�!�d�Y�Z(ѣ'�"�T$��b@'�!��Q|�����g����`	-~!�䖉G��a���.0���.��Hj!�ߥ~uĀx�nO��h���ªBg!�d��B�)��I������_;:V��䇛X��8��Ɵ0l��K���yr`U-lݬT�C@�7e�|���O��yb�ɩi�]
g��7(�(��o��y��]�l�sQoU7c[��U�B��y`E�.rBt��ZhZ�%���y�E�9����鋻O����U�(�ylT�oo�`P��3Gg��Pvș�y�@N#Z2��"J��7Zj\�UB��y���"rJ����B! N0h�����y���u��TS�I���ϸ�yB� Q���{���X���F�y‌�%B&-Q��=[Pm�%D��yr�G�t�9bfI�L�&D�&�&�y��)�~l�ë��<d�D���yBU
/���.�Tن���*\��y�LC�S�����JE�I��3�"Q��yRiҭYY�<H�N9�r0H� ��y�-]ɰ �7e^ � ػCә�ybC��;��&#�A���;B'�%�y��\�(ZT�B���2<ײ|R�\��y�S1�j�vnJ�9��iPP�[��y��TzV�����7帜�FȆ�y	�	����%b"^9��g5�y�Z)���)Ҋ�[��r�\�y"� `�0���W�( �S%����yr7����ƒ.x��g�#�y�
(;Up&��ow8�������y��^L��4��e*f!����y��N	?N��7�� lX���3n�)�yb p��a�RNK�e]���Ҥ�6�y2N#=�6�BA�^�^�@@��A���y⫉�QK��oW#GkHa�`�>�y�� "gn�kdn_�9l��!J;�y��l�6$��/��.l��r����yr,��,fy��K�
��� 	���y��C)^\=cgדVXlKS�
4�yBd=Ut���6��,�=�y��tC���#�W�p�c����yb'�2?��ȉ�" ��ܣq�� �y2d���PE�#8�3�璯D�����BZ`M�5�]�C�J�K��Ʈ����ȓ,��ԛx�Ԡ+Q`�!�hi��S�? d�`��	����P�{�k�"O.f-��c<D��kJ�NXs�"O�mJ��&f�T�C�KҭO���"O��{�س.wP�0���Й�d"O�M���ʥ7��3�V�F�4�S"O����B�Ĩ��矵:�X���"O��'�3<� ,�F�M��I2�"O䝁R� 8$�� "��[*�9�"O:H�<E����  J�(����"O.��&-��>y�lQ�$+A�$Q"O^آ�Z _pL�󃋈'�Z�۵"O��T	"Q����G� \n=("Or��d�ҿ|����a�z-H��r"OYy4�4l�,��7a��?���"O�X��̆m'��u�T��쩴"On:���/J�x�#e"�-����"O��ukٟfxو�]Q���"OL��OQ7T��2�M$Kr���"Oje�� �����ڑ��XT̸"�"O(tcUk_�Y��똇@R�1�"O�D��K#��K�JΣ^?�0�"O�����I�kߊ�"�'�7.��v"O�՛D&9X�)�'&zE<2�"O`c�iH
~2� ��?�$#!"O �qƅ�63�Z�	����%�"O����l�P�a`EI� ��"One�P5Pd~A��iɪ$�H��y��$=�p�h� �m
zq;�`�y�b�p�r���ۗM݌����� �yB�Q�@�P��m��T/4\����y2�
knh�`1�_:H�!��Z�yRo?;Z2w)V�<����slG�y�$�&��!L�$iGD�j�X��y�!ցC7C�Ϯ^0 Ȩjщ�y�m�.Ru1�
�I֜�R��y�O5M� ���\#1.�S�f���y+cĵ��������l!
�'��
��>>���E%|� ���'�������67�LMU��(e�\�	�'��l6�q$�C%��ibD���'���ŢB�4�T�ĠU�	Y^m!
�'�
 �0-�'I<*H���ǡM�4��'<~�su?b�<q!D ��?uP�	�'�~�*��ݷ��� 60�B���'�≫BKܒ.^v�˓�Q�\ݱ�'G��f#�W���p�l�H�l��'�
��f��
N�V}�3�� U�����'2A����4,�A�o_$_亨��'�8�Q⭓�9�if��bT���	�'ޡ2+�
@��²+R�F�0���'�v�8�������b-�*H�vM�
�'#0�,~uh�Kǳ pqÃ��!�y���x!deA -�=,����J��y�ŦQ����#�"\\tjU��y�:%P�A�/^q�$D\��yMϕ%ZF Iˉu�d1S��y��nDTr��pa��� �y"KE.#z����f�Z��L�y�a�
��B�W>ZFp�,I�y��	3�$cG,0"cB�3'�Ñ�yA�:���h��,�� ''��y҄�;,�SD�F�w,�� �)�y򭘤)PZ1ˋ�/BR<Ѯ��y��<M�jd`G�&OѹS+ĺ�y
� (�{-U�
���CrJs"O��:�X1s�2���BEo@D��"O�4��g�BAש)Y*Xѷ"OUq�
{� �z�iB�70���"O�ivO!%�H��HːFL
"O�xZGL�{�^i�6�q ��h�"O��8rX�(����`7��d��"O�%���<^8!���)C�pp�s*O���r�Q�D7l�����--f���'a
x�G�®;:�=��,��։B�'�Dq(�A�g��sei׭�䄣�'�8E�V��a����&X�f�j���'D��qaN&ɾ�;�D]���'���*3��4k>xk �;P<L2�'#j`��)7�6��7I��W�r�'� �r)N'r�!�f�\"b[�`	�'h�#ǅW�\�
%$Db�iK�'��S0�J.]����Q&XL9��'d"�Y0 ȻZO���ų2\�`��'�$�Q��;)}д��N|KPO*��!R�[f0��R��(J��$"Ot�y�fZ�d2@�Y��l��"ONQ��͖�~� �'�<<�f(�"O|������2���H�$A�,�Yd"O�3�ˀ�`a�4���	0<4��"O���cM�x{��?2n�C�"O�Ѫ��6T��R�*R���
 "O�PzAnѸI_)�T
ڙ?�:	�"O4Ի�%�D�ʄ�ܓ�<TsR"Oı0D�
y�Pu�RW�f��2"On��2�Z���Y&7+���"O"Y��ǑL�>=ʇ�����"OZ-b��9L��i�u#]�5]�W"O���Iܼg4�a�JwZ�ͩ�"O����E�0Aph�S�;+O ���"O����G�N&搨�g�pM���"O�S1oKA�8uS���B��+2"O�Ȩƣ��q��A�D��u�Tsb"O�(�N0sB����*1���'�جS�]	g>�h�E�$+�J���E!n'^C�	�Ut����$=㊍ӗa[(0�L#>��q������@	Ǧ�ʢ�'��ÕB�yR˛8�D0
#"!ﴜ�U�2�M��(�D�'썶���s�|���ϟ��F�sd�*A�fEʅ"O�a��n�J��`)B�\
Qn���]�T0a[1BdR��t��n8���ӥ��&}U�A�"i[@�>�O	8A�"jv���ֈ�;��%����;ش8�W�I�������(�O)�§�$
�c�#
��M@C�ɞI�(P�_%H�H0�+�^�U� ��cӤꊕ���؎/�ZC�I8�$�"��?r�4=	�L�$.AX����Q�l���!�BóOdMlk��~B���Y�|1�ª_�FE�a6�K��yR�	N�7$����s�⋫�?q��=0�-C������ÓS`0��$BԵk� �]��Ї퉚6�!��O<:���2A޺����)��e��!w⃏x�䬅�*�B���FI�2�l��W%�,=���>�1C��9A����:e��E�~bF)'&7�a��o(��D�J�<�"�B�z��'�5|�	+��iB(%��#_002\Q��'"}�'�8��c�.����ЮT��F,��'�z��H���͠Qj��6�I�nC`�(�� �Z%��iǁ��n�(�vt�Yir�*L�+@�isP�hg���(P�)�P�jc��$�tp1���bh,�Av�![ni��!P'W�ڈ+
��=�*ms ��sW�L�`fx>�l�?!��M��T�"�P6Cg�u���<�)��v�P[��ǯ�T�d��B!�dׁ��@n�զ\�]`���?S�v�e��6Xl�q�%6�x�1u�� �ٔ@��2�P��u%�O̡��"O�����c�tU�Nʝ?��-!��O I3rFG�la����'�2RP�?�TE��S��%�Ƌ�T��ZǄ�P���@�f4�i�&Fۡ\�by)fe�	���F#��7y��1'�w���㓪_$�TA���[R���.ғw��Kѧ2 * @���d��ubV|ʳ _I�, �!��y������a�DJL(Z"�X�#���?iԁ$ą�!ʚU~���A)ެ<�U�X�J��!��ŔC䉏-[���k�$ZXD�Qg�cM�ٰ��vL��I.��;��8�@�(|j�-"tX���L:@tЬ8�ˑ	%�3�9�O�1��!��z���s�X�J��H!�LB�2�J�m�09��U͔	DI�V�U���#?ySヨD�ؐ�Ћ=l!;3��J��l�q�M�>���l͋:_���$�(L�l`�$I�Xj^0�t��?���.��4�jW�'z9I�/"�`�<I�+��`��@�!��e{�Ùæ��19v1_QX���d��n��\��"O��YB��<5�dp��b��l����� ��|�R�M'8j�˴�i"P#|r�S�H�0�W�4��r[�i���M�jC��a�\%�&@
�?��q2���Jz�7M��D��H`�c,NfPSMǪ/����zrߣ"��k dU�]T�-b!/7LO`5�.�>
�����ރ{��B��g����Q "д��`�ٌT�̄��5{�:̈�&�$�:�ƽ+��c��;�έ�Y�E�˜-RX�CFyӉO<v��+9����fdJ��n���'pL��@O�8e{��L)
�P�LOt����[�7�N��ڴ"�>Q
�O��p�k��O�D@k�d�M{ m�'"Oޕ�s͝`5,<�f� {� �*Զi;.�R���g�l]b�4u�Z�*��d�)&����-�y:0��S& �az��,=X���-X��1�e�	<7���DeQ7�@�Rq%��o��r!'�Oʜ�Ue+L!��#��R0��p���Z	�.q�ę~���FF-bM�N|z�ɒ��@3m�'a
$r $H�<T�����W#Oz��R�ÝaU yp�lH�?��5�C��u���i@u}��vk ��$���s�bphg�R��y�ET�T�:%�6�аG�<��娛��M�.S������5��u2s��x�'i�l1�,Z���/��sJ�TAӓU�сD�)*�K�`�1P��$����l�$��7g�4l�L��NF��aI�7^��aw�O�*�6`�!�N'��'��`�#�F71�T}2��V�~��t��=+�I�߰q�Ǆ'�B䉽yt��4O�V�t8#�&�$ؚE�G�a�4i�NO�p�6��T�O���q�9 E�#��٨!���Z̆�(D�![Ɗ�)���1�X�Y¥o�/D��� ���=v�J�$C�T"?	���"ΥB��^0T�Rf��� �u+8j�)2��W�_��]�Ʃ[�!AV�y /�4h���ҵM�:����L`�j�V���˲��<{r-�<ɰ��;�-��o�&�k�������!��J��j�[��+�T,s�"O:�WL��R���H2��* �x���K.Y�T�(7����H�һi�"|�WR���*�
��4h)S�r��9Scm,D�,����.���ʤc�0/���֫n�Ҕ�G� t�����.<���X4�ɬ�Z�h6aD)*?��є˖8x/:B�1.U&!��.�n��Cq��TB䉴fF�ݳ��)_��B��_<WG�C�I�<���"�M�0☻�ˬ]EJB�I�֨�j�K:B#��st�����>!0j�����O7@mD"E�M�� 	�_�[kB@��'������  @�!�'G��X�H>!�/W�K.Y���cB��3��'q�"�sb �)#�<�����34-��<o`���B��$�LteҋGS�h��!2���r�u@��?��G}"ˀ�n��#�*�#s��9�	S��$:�f�|�C�ɐzjl*���]B"i2�l���ֆɎ��!,�F��h	0�QGC�;�&`XGK��;�,q��v`������v䣷����6��'����CgC�}����d�?S�\����N�r9ہ�ϣ*�a~��A�2S�(��F�P�]��s��I�wi�!Y`��� _�}��I�� 9�3OX�f|���O��HO$����A.4 ��#�i����W>��%�;	�N�� X:\BTcF�*D�� �0��m�`$��H	�����i�,b�ԡ (�q�̐<~bic���i�Q(��Z�t!�8JDG� h�L=�	�'4-S�Ã���!�s*N�& d�I�%�<�D��'�%k�	R����I�_��I7�	��ܠPaٻm����R�%o~��)׷"�(�R��<6�ykզϷbhD��!�Be	`��g�,�O=놤�*?H �5J�+޴1�`�	L�<邬�
� �1Z�k^�0�O^$�FC2J~�bIÎa\`Y�'�8�AA</�A�(��J�6���A�#n���%,�Pc�����}�]�c
��R��G\�5�0 �JL:B�I��P��	��$��!����|be�s!m0XJ��L1b?�#N�~Fzb�ܳRu:���Hɜ+Z^�ل����>	�ձa�,�yR��β��df�7%����tbV)MZ�Ѹ�$�f���͗n��@,9φ����`W"�َ�d��o]���\�<nć{܂�'?~P�kCfЄ{tza�!y9���-�v�SA�L�e����' ��-�	U��5[BAɱ>�p Va�R�O�v��H�5N@H�U��"*�"O�Q��U�L@`�ӭ%�-�GUy2	�7�mz�,S|��䞇#�v,Iթ@�K�i�iN2��~�ܔ;��a@��-�Q;��\,>�ā3&E'T���B��'L���τ�l�V�	6À�du)���KSr�`YE.(�2)6$�91j�"��"�)Q�}'�C��:OW���V-	��09�wBZ�`��'��`p"��	�m6���@�X�XU@e�� H]!�$�6Qw�)���i
�S�cN�!�$ȬG�Iӑ�Xvn�#4"f�!�\7;��Y��OJDx1[�O#of!�����"g�;[ں�tŇoe!�Ĉ0�q�E��7Dض��v�ڑ	:!�D�^�L� �
d.1&��A0!��2i-j��p-��R�t�3"X� !�ĝ0�Eq�� �P�3`�!�!7�(���E���(�-@�C�!�<�(��ShZ�w��+�T0^�!�$eg��/�	}j�h@�Nf�!�d�~�&S�G�5P\Y�@�h�!�D�5V&a���.!뤁0�!�}�!�d�}K�(�H4��|�T!ĥc!�$�"is����@K��� ��fJ6wR!�$Z
 �h�H_�D�,m$I:�!��#>"I�5f
7İx�q��*�!���U\F��2M]�$#�*$� �!�$3s�0�C�*(�1ѫ��y!�P\)���!�@ʂe��9!�dXX>���Ȑ?F�g��9|!�3Z� 4�WBH n�c1c@0L!򄀺2�D�樒�Mc`���X8V�!�$ϛAS�(e��4j(8�Q/5�!�H�Z����0��{��L!�DڤYօ�'m��S�$��Tg��,E!�Ā�J��	�����`(�����	zO!�/�� �S�H�h���+KH!�F��@���CE�ei��1DI�!��g�-� ot��E��!򄓭4�d���)U#~�q���N�!�$��G�1�f�� �x�%��)�!�D��L��E�� ��)-椉d��!��ys�9QC�K(�`B@�"2]!�D��r�&����,.�`�趄JSD!�$͕+brp���z�0�c)��%!��UP��;dW*UNJH2�(A�v�!���.=�D�1�L�s�����m�!��
HSΏh�u��V�9�!�DA1ZưT�s�M��9B( �18!�dY�8P(�À���)����(!�� t})��#\� oťz@QZ�"O�y��]" ��0"��=�VyR "OD�N�X^�esp��#E��TɄ"O��VE[0YH�8DjR�d�td��"O�0`'�'d���ņE�,d�a"O`�6gZ�hʼ8	#�REމ�"O��
���'X1)s��W�~0:�"O�#W��3e��|�Q�R�e�^H��"O�%!�`�"�B��T!�I!f"O.�`��]%nz���cJ"��0"Ov�aiH�D۴r2c�'u}\��C"O���+ i?>e	��%!�4��"O�=�!�)S����@�(H�P"OpX�&j�� u�&,E�b:I�d"Ov�[��Cm����B[�	�(��"O~�#K�1T�J����
2[��4	u"O0;�,�kJ����V�^$aX�"O��a���74�v��lF3��w"O��;�ZM59�6����V���"O�\�6�Ȼ�����M�]T���"Ob��6�ݙ-@]0&g����i�"O�Pۑ�:ik���& ������"O������<�p����3S�A�p"O�Y��r�0�k҉[���v 44�@�pJ�;(R����V��𝢅�>D����]w�0Iؑ��9o���QĀ=D��a�O8d�������H���PE�<D���e#�1� E$�µV��p(9D�ۄ�4<�����@�.��2f�!D����U7WE�d 
`M��A��4D�H;�b��E�dLK�Ι4�P0f6D�H2���~���2�ƢnTE` D���ã[:�q�1hn(�	S�8D�ܪ���+"��`qBA�I����E6D��43��]�$��g!�(�F�5D�(�
Z.24��Q6��%[y����5D��(���v��@�a׏)��ˢ2D������`!9%-B�F?b��UD;D������,���́**�u3�B8D��)�ɩ�BYP �-������6D� #a�C���V�5;���2D�hPT��=.v�h@��V%�Z�ben4D��@�%�	g���h��Wl��b�.D����Q�HS�)Ʉ��K2� a�?D� � Ɓ *�~�ґ&֟(��-�g�*D�h"d`)kaX��'� d�=Ja�'D�԰R:V����5#��UQ��V�$D��ʲ�&�ɦɜe����,0D�DJ恉�?�2�Be,[5�6|��,D�<��	d�ְ�F��e��} �#.D�У�ER�T�&LQ�B��3z�!��9D��A*�;�L�
�� ?�����D8D�H۴�ۧ`��=����%I�1�Ag4D�L��[�{	�y�e��@�ĽpbE?D����$T��i�E�?�r���b'D�(�n�v���B��(D�Ґe&D����Fn:��%�F�33�H 0D�R��7F�:,z#H�^`��r#D� ��P&#���#A�28l:k��;D��r(I�Mڡ+ro�Mpq�:D�L�kZ�Ϩ%�U��v�)&A4D�(8��H�iX��ߧ}ٴ,�QN?D��$B��(�<��g��4հH:�=D�D��-B(u,P����&%g�U���>D�� ��H��u��X7�%-�$-�v"O�� ȁ_3�g�<�:��"OX�q7��z����#F�4^rV�b"O.�k���{���B����~� �d"O4�s��0@��2�.B>Usw"Ori�FO��u[�ޒ|ڼ��"OB�F��6fry'lǱN�,䀖"O�]q�lT�z0@���_�)�lµ"O@8�Ce�4�b�334MZ�e��"OU���Ѷ-P��L�0[r��"Ot�RK�0C�R\[c�9N�D�"O�C�N��_"���'�?3�RS"O^��5�[(sp����6.����"O�@�D-Ro`� �2A�"O�48gaĹ*�\���	,'�PV"O�}� �64���H�"@� ���"On�(������<`@��Vs��C"O<	��P4|�X`r�1)�% �"O"�`�cE�LY���13�,��"Oh��vf�.h��g�
'\ ��0"Oj�Ӷ�]�7��eha�@�?BB)R�"O|�!�H�$z8��B���1�G"OH���ܥ��@(&@D� � "O�5�S
]q �rP��F���R"Ox1�ႅ���x��c:@��"OJ\�� $4�q���� /3zX3�"O�h�PN1.ۜMrG�ν,�p!x6"Oꠁ'� �"���ߡ$�����"O��R�ӵ^�>�c��@�xѠm�"O4hGl�_�B�� ��;�:I"O*�gfI�<�R!��/��?����t"O"�Y�{�h�`��--��q�"O
�x��& *4rҢ�o:l��T"O���T�]�#ě"�Ԏ3)pY�e"OV�����I��F���A"Of������\��q�ۺsB| !'"O����M�t
x����4��5�"O�[Pi�O�S��0��ڳ"O6�t��	`ٓ�!C(>�vp*@"O�@�U�C�t�zaʹ�\m#�"OZ!J��B"S'�U�4@/6r��#w"O��R�E�=2� �@��~���a�"OfElF���`YX�P��u"O���K-:8�؊B��.b�]�1"Of}1A�,�2|���v0L�r�"O���#��8Î��	��y�"OdM٣(�jV �чS�g
􍳖"O��vbR�n��D��M�o �"Or(#���?.@��1��H�0|�2"O��Xr�+� ���)@ Z.�q�"O�ceG�:�JYB93�&���"O�K����toJ/�`q��"O2�*���]����휆X`h�2C"O���I�?H'����"��8��$z�"O�MɢS# ����Ε�}�6��P"O.X�GB�b�f@�t�Υq"0""O��
���/�ʅ��f�yA��"OR�)ӎ���H ��<3z@@A"O��2�ЀG��k�d�=i���"O�0y&W
=d�@a��m��P�"OX�q!��;_X�%�g"]&y�q��"O�`H#���1�ՃƇ��\6<�U��E{��I[xq�P�����oy���Q@�lL!�D�{`�CG�3?2�{5�ųH!�� �� v���`�q�"���"Op��1#�!y�>���@�1?�z��"O��#�I�~M4�殔�4�00"OеR�њ�f9�� �+R�fd �"O<ljAɸ� I$�/� ��1"OV�F)Z2A����4-��"O��� L��nݖ��らC���"O�T���'%��pa����c�N��F"ON��I�``2Hq�.u�"�;"Oʨ!Wc�W�q��ԭ��T�"OҀ�@� �NQPdE^���3�"O��`fm	�v�f%�'%�i��@� "O"��t�؍T,�M	� L�p�"O8+e���FB:�z��� �V8�v"O�Zbm��pZCM�	>��ū�'SL�gi��v2�d"�g�^�N�0�'#�����"�����
E HY&���'�E�G.A�n��Ś"�X-@�:��'X�5�,^/@��S��4I� #�'p�У`�3Av����
|h,e��'���)�:\����	�A�T@��'�����K��~U3R/L8.L�)	�'��j�����ZU�0ŀ�-��0�'�m0AD-J�R�p^�+i����'���Sh�4�
����)0�"�'�`��4I-
�D驷�B6UE���'��쒤&X�a��z�/Qt�T��'��ձPጫ,7��Q·�F�\hA�'/�tQ@�]�K�.�$*2��'��`�P,�MX���A�+
&� �'��|`�k֨os��b�ʆ�UB�'d %�$�O�~���"y��Z�'``)B�U"L�B�-�)8�~���'R��[���$x-�N�9�^���'Ä���b͋.
R-@���.�~,��'*\B�*%#>��`�ζ6}0+
�'K݂�ި1l�y� �XAO�<����&f�R=���5������S�<�$˰H��R�/ޢw�d�3�VI�<1����NbP����9dE�,���\�<��+�1X^��'O�1r����!_r�<��'��?-<aFiU�>X��pn�b�<aCk�S2�PtϬ����EX�<��bK�n �h���K�2�
���AET�<��9
߄Ph���0� �ڣJJR�<A%�b:�a1�Km�H�B��N�<1�'T�Z5��$�ңH�Bej���G�<��-)�4�+�I֞HM�董�T@�<a�>5´�A�q�2���a�u�<Ն� y;[`IVQ&�8���p�<!�J;~��T�CZ�D�(SJH�<�+4)��ku��;~.��qO�^�<A$��9j@1��S�L@X�X�'QQ�<!��1"0�eP�8��(�K<T���Pa�@z�Rhw��	��#D��QR��R���M�]W�Y`�M!D�XZ�,U7p�dJ�'I�!���ի1D��YuO1!j~t� a�A(�)�!d*D�Ӕし �:�k5,�>�V��+)D�@�5d��3G����̲l�Js�1D����ϕ*_��UZ@J@�rI{5K0D�D@Cf -!N�2��M�>+6�IR� D��#�(�,�xАƑV����a$D�0� R�Io�,25��UA�U�$$D�� l�(�D�)P�l1#޸n�(��"O�*Яے(v�Z�/�i*�"Of���jו`I�M"Ed��65p�"O$�0�a��=VNa�h�40�H�"O��)�$��|t�	�F�N�l�
!"O��1�-ܻ=`2M�E^��*�"O��$�C	,�FQ�'Ô#�@�2%"O�l���J������F�Y�"O��3!��=*���ᇚ4����"O�)��+�h�,�w�J%`�l�hD"O<�F��R���W�[ T��#'"O����E�}D;�h8���r3"O��K�����!�	�L�A"O&-�����;����!*q��E�4"OVq����P�� ��iB�^ܒ�"O�@9�g���(�R��l���E"O������x�Q�ł�{Q����"O�,Y�j�3	�"!!D�"5�|�6"O6b�
`\-M�m?d�Y�"O
(�F���Qbx"Q�W�a3��i!"O�-r��e� J��B�htőD"O�Stb���a (B�	�l%Ҁ"O��2�N$�@0��E��܊�"Of�1am^�p%�bf�)q���"O@M��,:`�$�
��1"O��B2@Xr&juQ#���%�~�{�"O����G�H���9��"�N�Q�"On�3�@]l��"׊�akr	��"O.�r��V�Du���2�Z�eV ��0"ORț�KڒQƸ邉޴?� �E"O��b1 /���\���q�3"OB`f'�h�б*@���]���jE"OΡ�r��r��a@BŽ� iD"OLh��G%�r�;vaP�\Q��"OĩX��}Fd��� �D��#"O�q���6�r<"�L�nI�x:�"Oa���jҘ-ʂ�"+=@�:�"O�� +άx��A� )סk��=s�"O��a����H�W��+���xp"O������\D��ͳZ�����"ON�+�['6�ZQ�C«4m*�"O��qa��s�z��"N���"O��Аŕ@�&y�#4A���R "O��y�KT�6�6E�򇛓j�|�)�"O��X1)��0�瑅8;�`�"OЩJ�ڻ]k}��I���v"O���iW�}�����m����"O�}Ȓls�՚ ДSQ���0"OR��a~�h�R	ڦ`�8�9�@+D�0�AJ�<	pLux���s6ɓx�<�E�lM�	[����b^_�<�W��PLb�"�J�Z��g^�<YĢ��#@"9��lBy�RDr��a�<)�o����:!OإU�*�,�C�<ɒEҏgS\U;`@�1��APJ�~�<Yr�P_i�|�`i��b��g|�<A�I��rɨ!��Y����3�fQ�<y��,{1�t�2�/��bBMMO�<��[w���Ã� a���G�r�<���/h�\��'F�9~��z�e�V�<����/���bcǴ ���YCI
O�<�0�T��jTJ���3��䁑iR�<�T1aOZ jW�1(�"��҅�U�<Ia�ѬZqR��u��/l�d�c��U�<� 8��%����HQ3�=R�D\S�"Oh�0ᗩM񦀰���\:Zh��"O`��%�*5�l*2铦Mİ�2D"O|e"��LȞ͹&n�!P �"O�t�u)�gn,��M�(=*x=��"O��ڢaU���m͂Ym���"ORCk��*]M���}�%�"O>�b��KsPm�B���	U�i��"OV	�ŇίtR؂���9nH!�%"OH�hcD�5|���w+҅wZ���"O�x���Q�l~�� f�11N�Y�"O���aN� ��Ï�9���W"O�I��o�)���&l��$�FP�1"O��SA
!/��1��@�:��H5"Oغ��X#PJI)��B?���p�"O�}�g@/i���%h�5o�V�Q"O�!7�3ΚQ q�!4IJc"O���L�o��X4�
+xƈY�"OL��-ۦ&���P(�mMf!��"OC$KWT��\2G�"J�61��'��I����Vf�x��?N.��"�'N^mҁn	�P����7��J;���'j
m����f�����ȸy��P�'���ʡ��N��(��os��C�'ajt8���a	���D�:g�V���'�!���K�x���E	(T�"e�
�'P:�)�Bn�#�G6RP�	�'r8Pr,�9��3k@0;:nqp�'x<�Bw��c�Θ���JSj!D��k؍C"���`�>@L��H%!>D���C�ݻq+�tpV茒hv܀"!�'D� �� ƬAh�d�$��,1>� zRC%D�P�'R�ʈ@�&
��D�q�&D�,"3��(.ni�#�OP�d���$D�P�4�W.G���� jS��9� D�x��i��13�Y���=IŒ�(�#����6̩�
_�h�(��H��aT"O(��I�:����G��aA$�X�pD{��)�8?R(0jnׄkL8��dϠN!�d|��`yWE�w5��R!-^?e��/���Dʇ�j-�(˴`x��f@os�b1O���V'$k^�@a��?K`���"O�!
S �"j|T��c/�A�ڀ"O�M�oЈ(�j��Ӎ,<X �p"O�1���	�<��d�ߐ;"���"O�U�f�C��ȖMVu�&��2"O"���f���F�)Cj�<r�,��'��S'�.��d�\4���'�-� N�t	p@Y%e΀@YXA��'��X����[&:=��� g#�)��'b�p���ߘ>���b���K����'���1sM�D�0,9�W�W�rE��'�I"=(]�gL`��m��'^e�o]�+�:ux�ς�"� ݀�'���5�h��8J�ɓ)��Q�'S�Ӗm� �B`��k	D�I��'`��*�h�_\t:�e]�me���'f �"�啞r�֬Hf ͌f����
�'��Y��`"��j �Z3�@��'����o1��I�c�Tް��	�'��i25�f)8� 6]��	�'��@�֪�7h��b��S�(&���'�JIP��ز6�2�g�+��x
�'�l��T ν�>t��� ���Y
��� NmѣN�]���фKV.��80"O� "vA�G�� ���,F���2"O�ԡć�Yx,R���/�Ms�"ObM�PLշDm�t��ɑ(�L1�"O��E-�v�<��&�Ն.±3u"OF+�a��f��f�	�(��u"O�q"R�(�����ݏ}$	;P"O $��*@'.j``�JY�t`�I g"Oi�����i�pCI̐]CV��"O��j'֨_��h���c$P�[�"O�p� K��*���	�%-
<�<X��|b�'o�	����<X���@KU�H�p��	����4T^H�t!�:a����i��V�h��
SΈ;� �G"b���O#R�E} �h�$	�`e%�6��D��{�,ͩ"O�$��L�1�:���=}�ZXҲ2O(�聭� _�1O?��M0/N̋�R�-�Xa��7D��*�"xn�
��P�e' �pu�0?�G�i�Dm��ɯv�r$i6C	,�U��葝Z������3s�Uڗ@�:����5md���$`�B�
dT�9�iqCh��dL!�">)QA�p�O�\�����S�4=U� �OP��y"͟'��%rA�գ^�,�P�&�~��)�'$�$�4�a���R��A�Lx"��ȓ(.6|[�M{�P�z��1Z]��SKpA�v�= yb�B���m���#��ܳ`��t��Ԇ�n����ȓh�=�
�:Z���, T��ȓV&"��(�p��T�ÞT�~�ȓ!p��B�X�pp���T⩅�W�0! ��7e�9��ݫ�r���V�DQ���,0)��GT1M`���w��}�4i��
H~�4���v�̵�ȓ8���J�O�V�[�Gɪ�|y�ȓ<��Xӫ�x��r�*l��K<I9T�ʓ\Jv�RP�F{K^���+8� ����}0�b�Fܽ	,���
�d:�.v7x<
G��{��I����!��gMn�2F3G�(��Q�^ha�������d��DT~�Q��Ls�xR�M4��A��lm�q�� ��%��8xS�M��b�*�eL@9N��9%8,���ȓjW%z��W�%��=z�a�	��U��P�F̐"�_�5���C���
n1�=��{+��$[�xN쀷._C�`݄ȓ}�*1;��'3��@ T�w�؈�ȓL�<�	��ՠ$0E���FЅ�33:��r),J�de�5��
{q�P��;y���.U�Z �Pg	4��L�ȓA�L8	B��ul�m�4a!TZ!�ޖ����!�$�ǚk�!���NDt� ��-!����gz�!�D�%����`Ι%J��"��@"�!��ٳ|Ե��*�;x��w�<Wv!�$:"9�4風�i��,@����!�Ă��n;f�Y�o} �S5��Il!��<Gi6���P�Xg�����#X!�](`d�R&�mTx}�#a�Z�!���W��[®�"(��`~!�N�L�bT�k��4!��y����n!�AE��f�NPիsH��!�D�]�T�i�f�e�f
B@!�7W�qH�0���G�<!!�� R]3E%F��9�1�S�b��P"Oޭp�N��W:�#�͗S���f"Of�*�R�fl�����KC�4��"O��y��`�01�u�E0G֠R�"O���7	 D�i26H �U�9S"O����,�59����p��P��"O^�8` �
Q������N�"y��"O�\S��2L��3�.��1w603�"O�1{s�z�T�j�̞� JjI�"O��"�aD�^#�dz��N�#=졫"O��Ғ�~p��+��;��q"O��BC!_�v��ɍ%3��7"O�)a�PT l���c�P�"O��� ,��������#�)�!"Oօb�(GX L�֜��"O�p0�#1$��2�˦;�E2W"O, 蓯J�wR4��bջ���"O>,�U(P7n�`�3���-`�"OB��@/�?h�[6n@�AѾ�S�"O,��K@ � (97�V''Nl�"O�)YĪ�goF9`a�5 l�B"OX�9��V-֘ �ʰF����$"O����(C1y�aH�B��eIS"O	a"B�#�}�e�j9BAa�"O֘[�l@7Q���p��!Hbe�4"O��kc�	#|�$�� �U>6���C"O�ջT��	(f�|K�hR�y'��`�"O�e1�^��TqfGGc�)��"O�
�I��@���s��2jڹ�`"O���N�u�n8xA�Ѱ(����"O�E���V�%�|��7�(!7@(�"O�L �խ0,�`�O�,8����ʦ���4e"�⭄�,��'�R�'b���ɟ��!\���I�e�`�!U�Wj��		X��PWā�0���&"|���u�\��L��g۴Pd��#� �h�н�4oǜ$x�F�~���d�
 >"���ʕ+9
�'eD#"v��	�>]���Ʌ�M�GG�~�'+r\��۶�یF٠�b%&Ɍ4TZe�\8�hO?�ę6 �4��p��5'ph�G��Ys���ش|���|r�;>��V�Ђ'�1�p��b��R�,��aT�x�R��Vߟ��Iϟ��ɓrp���ϟp�I�}̦��B�@UN=kQ^h��{w�[�3تe 4e��g�U�%`"E	zppk7�&ؘ�XWc]61� �ٲ��I12��F��L0��F)Fi����-��H��#ʓu�<���Gi��cU�f<���h"�,���M�����O�����y�v�	�L7�Uh��\8+x�j�"5D�<���6X��X�������  e?�"�� 0�vW�\�"Y�u7�'��O���	�圥>8��S6������{��'YX|���C8	��El&S*�}�p-��hapŨE�{�.Pz!�Wn�a�R	J9:�Q�ت�hH�M�nds�DZ�%���!��%:������ٰ>k�,i�� ��ru��B�4	��������"�i�n�$>io+G�T����{����a�_�_��������?�|*)�R��0H  ³��Y�����h�1�p>�S�iL�7r��#�lS�C����ʞE4 e ��)�M�7�N(=���'	��'�����-jb�'ƛ��E�(Rc�#AF:�QFCׯ�,d�W+95� �;g$�WZ�-k�-�r��+�(�|����5vA?P�� pB��p�\)Ku�o�/i�^�q�AI��� 2lZ-K��`r��E�8�@T�-�1H���
�K�.�����[x�hoڽC�^�db����ڏ�i;��"!�?t}�֠]h�j���'AR�Ih�xM�����;�w�Y xGy�/eӊ�o�k�'�u�&��|����ֈXr:P�r(ʳkm��$�O$�	��4n�����O.�D�Op�;�?�ڴx����r­f���K��X�Ɛ8�-&  �X5lVW�@�J�H�U��Ɍ�b�����|���E"~�)� �^�p��Ӻ-~h�ˈ9
��ѡ�	�^&�⩟FtX��A��,�f=����2e<���C�.�`��R�'�)S�'��6m����Y���ID}�4	-��"�%l�*��tO$�y�+�(9$����a�`	��jPs�LEo���M�*O�d�&��<i���#�:��e,rI07d�'<\�fV��?����?���&�R��?��n��R���M���۠��<�0i9Ab�&IX�ȱ󏁢%R�<R�����f�R!N����l�.�p��d_�do��
b��,�E"�~X�S�����#vI(���O� z�hf��?ZTurː7U��D�՝>��i��٫uMV�z��WfD�$�(��oM���j���O����O�O��S��  �,   �
    �   T)  �2  V:  �@  G  �M  `Q   Ĵ���	����Zv)���P%G�AC ���ײH�Ąa���8F�t��$!�~e�S�'ll\�02���ň
�,�|��h�\��)"O0� �����$)2U/�1&���f-���qn�Z�ZL�r�؛a�
����	�n�
�*�;23�m��.���v��G�+U2�$���Tz��R��أ2,l���A	+���ef#;n��"R��zk�X����@I�\2�߭.=���`�'[�H�)�D4=%vMaE�� )��C�)�*t,�#%���?���?)�<$���O�x�׮��
�X�X�O�0 3qy�%�p>��-�S�	��X��oy�HC��p>w���v� Bd��f���c`ayr����?av�'T(d�`��=�PCg�=��%3�'>�u�J\>o��� ��&8P���41=���~�		�jUV+�9:h�ZAo��o�4T�S-��Ϩ�����Iџ�Y[w���'��醮JN%t���Y񣀹M_L��ƩXE���D�+!�M.S�l��Ɏ/��(�U?��}r
U�?d6���+�fM�S)�zx!�$�1^�� 4-��t7JHP'�Y>[!��E"v�%ӻ6��Dp�ĩk%��Qf�f�|B*!��6��O���?I��2Đ1%�R����� �M�B��?���?��(E��?��y�O͐����:����է�"$d�}���$�(�Q?m)B��zUԭ�_�")��4ړS_���<�� M����d�H3���*t�pr�"O��s�ɚ�����!
�Э ��'���$��#�/�ꌡ���&7� ��'���Fl����O8˧d��k��?��N�	SZ�)�E��"H���&.ޛf��"��T>c�x�!��"��`:�?���c��O��K��)�!HEhv�ؙJvP�%�:HBh��e��	���S�O��š��Ŭl��5p���-�!��"O�Ra�J'm��p��L�.T�,:5�	�ȟV��D݁  �y�/�<?��5��Q��П\s�Jļ���������P��kl� *Z�&	+B�n��D�0CG������BJv+��B�vT�2����)�K�'�.e"M"� ��"�O�&�s�2����@N_d�J�\����B�0�}	�����d�*�H��-�2(�yi�f�6Û�'���S��'��H �;|�'���]z?�)پb�tX� ��-=I��Ԧ��ϟ���c�)���<Ѷ�A
�4@e�P����{�2$��.�>Q(OF���R�D�<�/��h�ҥX��Ƹi�-��	����?q���?���>����O�$}>�!�O�t)4gف-^zi��8k6=�E#�yx� 醥���"�$_$�`뗋�&O}6A00�?�O8Q0P�'�Եه��#2ԍ�A���d�1f'0D��і�L*	�P �V���Cu,�J 3D�T��k\
���r�ɞf< \��M�>���iV�'z�L���'\B�'��I���j�p��D6��i�f曖��3EB�'�-TI�B�ԟ�0B�j dU�d��x�����ɮ �Σ~2�&\�0]L��Te(>=J��I�x�'�Ĵ9�W�>M�ED�4k�J�&���'��ׁ:D��� �' =H�����7;�,C��-�O�-�'�N�(������鐳f��+��I�O^]���ܦ���ן��O��D� �'m���+�@1�UO{k���-�'�6��9_ߨ1pK�U�:��B\�<;�9[�Oj��?����j��yZ��K�#R$tR�ĝ�?�D�S;�Xhy�cO>O&�\���4X���C<h���.�|����Gu���kޅK���Ϥ�?aD���L#�4\���'-��A�'G].��ΖZG����L� �H�ЬO*��O����<����?I�TiD�k�)т2�[�I�"��E�vn�j9�v�|��'(��'��d�O�I�ok�9�����T�n�ڒ�ܱ,2UnZ֟����Zg��5柤�	ϟ�I>�u7�'chYq��o���k�!�p����fŢ<Y0)�HaR�@��0<�Gb��F��p��ϛh��	Fd�Ay���8o�8 �V3kax��ҿ"5�|�5�(�R�a`"A2����1j
B�#LO�Y��+
 �����	vt�j�O�����>�zPM�� c,,q7���Y��4�<�O�0cA�Z��(�Տ�n��9+�	�5,S�!xF��O����O �$��[���?���@�T؀"�R�f�գ �ßS�,S�*�_�}���S�0��|y��̩q�"?9WΆ������	|2��Ǡ�6mѾ�+��< ���1�O7Ad��KUʗ$K*
�
?�����D8��`펴5���8B�F�NfH�mZ����?����䓦?y��<Xp��W�8I�mYT��Gu�]IԿi��'��$2��S���i多7=JM��4�?aӻi�\7��Of����3����O���n���%� 0��ceX�N��]q����K����8����%m��~̜��G�s�6͓�;L������@M��I(�Qu�±�hO@5����g5���N�^-@��SK�&F�Z� h�*%�I�H�,�@�� �(<ö���hszX�=Af˙՟�2�4o�O���$�O'DJ��ZtDɻ'kZ�9 y�R�$-�i>mEyR,��]��Yp5 C%�F�T��,Ͱ>�c�i�(7�ήW�
�S�ӽ#�X��r�		��8�'���#*�>����	�ʆ�d�O���P��+>��ھ0���`gڦySTB��3A��4���bEL�?�l���O���?}C���Z8 �"��c 	��_�?1��]0`�$�;�F�J]*q �.	5nY�A�9Sz��O�(��cϫ>l�8{��1���0��'8��������~�D�D*�HrE�c��NU��ƏA?Dh�O�d-ړ��'μ	RE��zv�X�W���9ZD0���dѦ��4����*�1b�7&Ў:��@+�&�3 ��v�'��o��R�<��'E��'��Gm�)�ɓ�Fqõ
,#\�F�.
?�;��n�HeK�BșA�l�%�#���S��R��\�+�\/�B��X0vLبQ֪��QϺ�"�=YoQõ�_�t����)Hu����$�}|�C�9Ts按��I�P�=�\�$_f��p"�B��j)�!,�^�4�)D�p��e�/�HH�Ŋ6o��]�d}�J�Fz�O�'YY��DK�c�ss��,b�|�Wϝ�,�v�Q��'��'���~j���?��
��?�BP*5{��A�ьuV����M��T1S�@�L��Q��I�a ��z�.Ǟp��s�e��HHY��V�t��8s��Ѹ =F�����E��	ct�ɰF��$L�Dq�L�4��K�^!Ҷ�]0��m���MS�����O��d6�Ļ?=�!��3x}�D�m�%mS�=h��7D��)��^;E�
��H�ov��	Fev�\�D�Ŧ���4�?a��i�;7�b�Z���O^���d)q�#�h�t	�S'D�\�Tusźi2�L*��'t��'��u3a�ɿ�tiR�BV�j�Jum�?	0u(k.$���J�n&���2�hm��K���8��Q�V:|�����9Vd��x5nß%@�)��e�� i���G��P�'��4"��{X>���jK� ��ș�A��r:��x�>D�hy�$�5!���P�఩��:�O>��'!�mx%T"ZfqF'^d'@�O�c��!�IʟȔO`=�W�'��*<n@�a�N@�:	��ˋX�7��y@2m ��>,ި� �.= �l�4E��pc>���Z�Rh��ٽw���{�fQ���6ʈ��NEzfnQ�@L�I��%�Z����W���<0�A�G"�V?$�Y�Fـ5�*�dܴy%r�'��)�i�O��ɈH�B����*�}j��ԭ:��C�5p�H<S�
�.�t�3��2u�"=1��,�pK�Ȝ�\��80#��1J b0h�4�?���n8te�N��?i��?i�b����O���"���{�xC�	���'�MXy�����p>��o\l��sH΃p[���֠^QyR"�:�p>��͛��e���_*[p֙���Iy�A��?S�'R��tAK`C��1�'+���!	�'yl	���K
k���ʠo�&#2� �ߴ^G���J�I% ��qɵ�٦m1�TRu-'�����Q�i�I���	ğ X\w���'���ΰUli��׍(Z�)s� �D�<lړ�R�c�6]�І��p��kO=��H��DW�b�k+� U�B�-�7L�;��[�=�H��C��4��TS	(ѫ��fJQ�TH���O��Y�ݸO���#���2&�b���iUA�<�B�٪F�@`z�C�O�@��&�}�<ѳM�%���pA�2)��2EG�y}��{�2�OR hǨ���M�	ڟ��'5@����|���`g�T� |�o�m����ן�I@q��۶lKٶ�0�*�?�';�
��Y�]�`�%��x".6�{ȅ�E%R
w���1�/̫t2~,*f�}�=�G�1�d@p��D	j}�'/�?��I�	����3V!*h����\#�hp "O|(��օ6�B�˦���tl�Uj�'&�{�
�c�1LH�D�H�*�H��'h�G�>������V�3���$�O��Sg�K�D�����|�f�����B�[s���:fݾ�)�HQ9��ɻ|:�':��#�O��ܜ{�*Q3\���'�p�h#/��5�D�8w%ٕ0,�L��	G�z��Th@��m*�4�c�|~�UNF�A���	�@=������(ߴ�?1+�$�;U.%j��@)Q>z�Z���0�!�4�����Op��O6�$O�MkHW"o����Qj\�Zyf��cN�ۦ�&���	��ɿ<����ڕe�&N�~���13�Ë72�f�'�bA=�L�q�'&��'&�G|ݭ�Ɋ�0��&�ڙ۳��8!fx� ��3��Ƀ OӠ��,Z1@���u'�O��\�?��_�83V��b��
[,hj��H'O�0��� #�҈yP�� 6�\�O�h� ̞"��|I�?O���i�#E��	3N�!�*��[�ؓ���O��n���ē�?Q��~��[��$�0	��r��MK��'�ē�hO>iXБx���94c�Ƞ��Mo�vxJ4'��Msg�i*�7��O�(n���l���?�O�| ��8�d��9ڞe[��&te*��'���'r�y݉���dΧ�Bsf����͸tC�:0�4+�!xD����ڑrRX<��Ͼ�pYq�)�6x@���E����,�Y젴#V"�:��&�8Y�L��ʦPK�]�/V��<�P/B��<� �Q�ĉD�?�h�����nL�Р"Ov�1 ���h4�����b@��"O��cD�u�Uz�(ėi+����U�XS�4��}g�!Ȧ�i$��'|�IHM��]q��@8(�	q�ě�>�f�!-���'��&T�>B���Sp.ڭc���-U��#%�+|�\��A��[d&�I`�E�������+}w�āŧ
7id�=q����x��w�COmLȢ�W_�H���C�e'JH���6�1ODX���'4V#|j��JR�49s�����ɐ|�<i���,%���i]�5q�ep�hQnX�0�O$x�N��U{�œ�ִd ��P���� �M��?�-�\�P�M�O��D8\b6�J䇗�(�ܽ�b�+#~�o�{�$`���$tD���c�;H�,�鮟�c>Ţ4���z�,��͎,5��CG+�����M�0M�2PS"�!C�� 2w��`�O��$ʒ�\�I��P����0ݰ�R��'N�ū��})ɧ���$bT��w��)��ȋ@�e2p�!D���f�E�t~yC�e�V�̝�p�$�ؑ?�cA��1�rP#BiO�z:���#�J�M���?䪘*0a����?���?A�����ƾ�Id�N�\q�j�1�LR�fƂ�'V����/u�l{�P>�<�u����茲��D�O*N���
�n��@�	�L��Ԉ� 	�Mtf��(O8T�+˾3�R�!աES����^��j�G�O ��I�x��p��"=T(ę��Q$�C�$dd ��j�!O���gQW̢6mSs���Ԛ|��sf$��b�>g�`�h,� A5�Ȍ}+B�'���'/d�ȟx���|Z��,��&"��)O��6�	Sֈ{�A�|Ga}����D�ڳB͟H-���(�1���5�[7�����'4�A�;L�u A�H$�h@� �+����"O\�� @�U���RC-�����@�"O�Y��h-:9��;�,�QY�S�,2�4��s��<+p\?e��nb���!`�tb�f��My�$���҇�؟���⟤C� �;KT�8��Hɣ� i������+�Q�z�����H��L8�hO^p�u癸N�bh�"��-�>�� b>=XQjK�;��ݒs΄R��ؙ�-ړ7V���ܟ��}��ɵ͈����c��YAuk�W}�'x�|"F[0Y���㍄��J"
��>�b����r��L�e	�_�0&����>y���{����'8�[>�0d��ğ<��=J�R�����;O0���c8,v�8�4:�Z5��a��:z���)hBu�0Y?��|���\�3I�����׮^w d�E���?��b֐V:Q�v��=c�x�ȴ��u�e�g�1��⦍��~^d���~�8�"��O&��W�'�B������Ġ��s'�5�д�V�J��{C-;D�L�5aF8�t��U6)Kx) �L-ғ��?I��	�g��,c䤂���9�풵�Mk���?i@j�@i���?Y���?�c����ֳj��u�5ȓ!{ �%Ӓ$R�P�娒<b���$�U)���Jc��H�T�I?,yL����6+���sk�O�L"	�6̒�"Q�Q"GߚqZ�ǣ|*�𤈘��˥�ӵJ�)�d�[�G*�I�N�(�$�O��D&��Q��Ցv�	kr.((xQ+C��F�<9���hQ����f�(oJ�H' �˦�Ì�4���Ļ<A`�f�a�R��P�,
A&�G"�#wS%�?���?9�\)�N�On�Da>Q�'�Z�G�hLssO�"s�n}�g��]W�ܐBh'�z�Ct�@�ZaEB&�=PD��I�)� ��0-�(\�%���0l� ���ϱ$�v���:�j�b�OT�B6b��	=hl4(���� 9�@��C"�}�޴�?Ɏ"�s�44#�-�<�$�z��-p����u"O�h;��õ3�4`B@���E�Z�`��4�?�*O�嫔�Pͦ!�	̟��'p��X����&۴3ʑ�e�,Ln�>+�U�	ԟ���j��}q$ڞ~.&� �@�z�j���ܣ%:8�b��5hfB戙?m\�xTE>�d:<]c%�^.0H��K��m�0Q�cұbk��\�2j����EZ�bqT=ID�1�G ��I��`�pЉT܈��T/V�7b�q��"OP\b� �S���t�LCt�R�'�x�-�e��	j:hT���[�t�l�S��QA�i���'���P��X�	���6j_�:&p���d��]�^4��W��M�$#	�d�F��ҍ�t� X;f��q�d�F	D���Ou�K�-� W��C1N��b��'�\��r�#ՠ�Ӯ�01�������8 >i�}�M�=7���EE��J�q��?I(X��(1L>E��&��Z�I�%�)\�@`"s��>�!�K�}j��񏗛A�`A����Rޑ�h	��I�`�n��@�'W�nI�g(^4�&Ho�㟌��<=\	)��ğ����(����u��5��ݽ1�0`��D/a����d'�_LA��; �T�Z�k�(v2)a.�J�Z�M��ē¨��N*u�`|��	_,"���yPjǳ�8(Z��=-�>��2JRD����'*�j����F��~� X�$m"�B�e��P�h�p�+ӂ��䁗�b�;LO� �`���׿K��Dے)#Lx���"Ot�!n�?�X��.>dq&Q���i�:"=�'��cG��B1��fDFq�a C;KF��S��n��b��?���?y�����Ol擀C.�i �)���x�ɷ�^�h+Z� Ñ$��8`-��JB2���e[u�ظ0��I�$�Xc��J�6��@�
�l�:0a
�Aw�<��������4rNt`��t���Φ7R���5j��nE{u�A�FgR���.��3 ޿f�����B�2�m�ȓ$���y��� 6���
2�`�a�' �7�:��\1\8�o�����Ih3�΃gܐC�gԫ"Ua����!�S+�П������k���=���
3g)x ��S�#f�]�}�*Y��A8l�o�'�28x���;SM���1_w��5�S욆l 8��t�ŗ0��=�m��4!��i��D��=��H-\ߎѠ�T
c�!�\�a�|�RFj�:6"VQ��Av���'���s�X�q��Ȕk6
9��L���'g�Q"��a��$�O�˧zL1*���?a����p�H��7�X>F��L��$��/Q��вH���T>c�  ���uM�!����D�@��O� 1��)�'..*dU�e�Kŀ �E��A"P�����S�O��z'nG�����Hɩn$�x8�"O2y!���,pŪ�
���Vz� @����ȟ
p3�e��	��ф3ю�ҦC��������2	S9e�n��I����	�d�]w�Zc(8���.yn��bS̜4n��F��`{�h� ������I-.��Sm�'�@����,d�Y@r+�>JҤ�G(�;ɰ嘳��$��i�b� "���#iƜ�E��Ԏ���M4EX��'ejP��sBazR�ܙN��h��N�"GZ��b���y���[E*�7單�ْ��;�M��i>�%�4;�[s�y�b�.
@p�H��,%{d J���ڟ4�	��	���	�O��dAPp
����v�K�f�r������C�(�e��$@2O�*~�t�2.dD�`�*`*��B\�
�<�`Ed�Rv�9�������b��%j2tr򀈟/v����g	7��%�I^yR�'�B�'[q��]�h�:X�22���w��X�7"O�%5�x�B|H�F�f�6�c&X�C�4���Z��cOU-a�<E���u[L1v+aӴ��B'�9�-	Q�ؠQ����"O���%�
ZҰӃ�̾�ض"OR����͖YR����"?1���t"O� 1��W�~�8ǩ1V~X�b"O�I)ׯÄ%�����ϲ2��s�"O��r#��.U�yZ�/�r�I�4"O~<���UQj��enϤzZ��"O(����5{��;�ۮpQ��Ie"O`1����4�.p;2�K0,&i��"O6=(EL$0|�b��Q�*"O�:#H�
JT��O� �xa@"Oj��aE_�U�L����-x��"O�i�h��upHB2�ܵow��c6"OB4`�EԿ{�xx��Վu�@��"O*�ѐ$ȡf���k��μe��"Ov1p1-�= �$ܫ0F(e�p���"O���� d$tI��⋎��pY�"O*8�!o�9idt�[�"D�4`��&"O�MSiR.2��M�1��QJ�ͨ�"O��P�ԲY���j��O:Kb����$R�3�����T7`�� �1!�3(�D��T�h�!�9f^B�С�8/�R��f'�!M�a�-�h�1a�Q>˓i�q�PN�pv��`�JG���n��zu*�
>���ۿM���5&�'¬�7��0>�3��cBx�4�Ο�2�Hex��0�~u �7�X5�J�Q�J\�G����ɢ�'!��K%W��\����M$X(�bMǼ�CH�R͊�9�:}��ι�H�Z��Մ��?"�)#�`�
-�,���"Oy�u"�W��\��A�����iB���BAxQ�����eF��u�g��7T��EK@�\�%f$�2�7J�vC��_�(C1�3w���8dJ�T����Ts�8q��:Z�ʉA
�k�qi�隼L�a�E ݘn����IW�d�2 Bh�u�t��՟t�2(�7�asӫìw��P@#'D�� b�pNQ�$q4pP��Q�v�(@S����II*l�D,ف�����E�4��<y�}��Q>
��8b�f���y2�?</2���@٩E��R�K9~����*S�<�SLQiź��K~�=�J�!]~���m ]qhp�dd�\����B���Ԑ�we�0M�B-� 4`�y�C�;�ƙ�$�'3N�Q�ȣ~��v�,.xq��V�b��qd�n0I���Ѭ�`1��LɄ!X�k�/e�d�#h2D��;� ��x���q�D%X��2`B�<I4��!R`d�wÐ)y`5ʢ-�����	 S�kj�`�`�*�ʨ*g"O\){	B�_��S#'ٍ.  ��Å�' e�1Dur����	2}�1�1OxT�n���b����H82��_!��W�9`��r"�U+l�j�h6+<��I��dIg�^��¤Ư&3����Ò%�E��F8� u�b�����	4yB���
�)N� �#�Цi9a��Y�(`��C�&Uff�ۖ�:D��A��J���S�n��}�����+}���"_���'-�7v��\���?p� 	��F�vk��h'�	2,�B�	jvd�ߊ\��L*�bF�E����oW&1�ʓYy4��L��r����;�33�\�J[>Q�Ċ4D�9��1�z\��)L(�*�풰y���j��D���>	v�bj� tM�
��z���{� \Qů�(I��|���F}�J�d���C.�X�M�?jo���e��=`��8�&$\OFi�c�ؑ%�z\�&e�gZ��ش�D[�^6���Â�4���I� ~�4��m���YI��E� �P8���^������@l�<)��ٺ}N�](�-��=ՠL+��_?qP�JO���aR�-�~p�h�|����\���K= �CB%�r�<iW�]�b�3D���M��i%c�V\%�#!�Ms������K?b�{�*�:%�PQ�%g�^�	B�f݃�p?Y�����he��i �TQ�
��=%���v6� �����%�S��<��E��4�H�\ vm#��1�O�=`CEB�t`�f�&b]�=m��oJ�Z���c��lᢀL'3`n؇ȓo8���暫��i�c�G� ������dJ�3�r,А�B}l:�'-�T�����?t��⠎�l�(�ȓ����Q�S(lG���P��C��a��/9����ܴRV
��pl(�����'�8
3Y���X����A��d�~��b,Č��mQ�ʂ
J�DL@���L���y��E鬨��O�4��z�CH�L�����Y�#��H�	U���O�ʆ�?Z��:�h�1��÷i�����L!_����*ӏ"6  z�"O C�琽{�hm�0l�1M��&�Ol�REo��A�F�h��%aC !�q��(�DU��+ī&��} �#����"O�yS���`)�R�;U��S`���0�~Ӫ��`���q1��O
2�x�p�,\b���ER����7�O�-���-P˰T�e��V��������ѰC�|�
�i�nG-O�j(���3^F�8��O$r#��E�7XH�>�g �#N�|D#5F�0y4Py�W��㦅ɖn��j�f,b��}_��K��Zd�<�an]@���h��Vs(���Ia?�7�L;W���B+U���1���|Jf��-���aq@��*&	r�<9@R.+���G���~����ƚ#d�峀-� �M��K��^!T�YI?��{@�_G����@f �Su,�p?�_ �����%�<�l���)���u�[�B��F�UvXq�鍑�p=I�ѱHlP�:E�¡+j������L�'������s����B���Iشc�ȵ����� ��D��'Zp�w�8Sh�!�w�ƅB��S�'hD�C�
	�Kw�d`��"x�:�t�O��P&ɢVl��e�4P

��	�'A���bve��hg>%Q�A���p#�iP���H˷��}�qO��R��ь0��$����g�Td���'Y�-� O��CS�D�P���v ̒`)E�R�P:6�B�.%�x�b�<)�����
t���O
�oF����냍�Q��A2E��>�$p�d@����r�&�:S�`6^�"��ܒLE�4D��(aI�$�z�����)��".D�����ȑ�!�M�Pv���L)D���eR74�0�qS�M�!129�%;D��j!�N�$�q�� 
a�.�*��9D�,rI$}�d|�G��|d@��ˢ>�"��p>����f���pDO
r���YV��i���3lޒ"lL�)� 
�xl���Э�3E�4eδK�"O�`a��T({�����7K:y�7��ݲ��X���f�O���6(��_R��F�V�/�<B�'�:U8S��&j���6�ݢD�,B��C�s�kN<Y��>��F�e�ъ�I܈��m^`�<��O��2R���I��a�ȌO|�+�(U1/n����2@�]�RW�W���7���z�셥&��8a�����ԭ�q�2)bw��,�>��/6D����P�[�.%�D"|X28���L΄%)�#^ޟ��@ �kH�C Jb0#/Ŕ[0C�IV�,2ЊL����"��3E�42d��C-��Ѿ0�d�Cv�v�g�O"��f"«��Lz�.ēȡ��#q	(la�ͯ{��D��W�%KP8���66�����bYn0zDX��'?���������� k����Q���aIƠ�fT� ��2�����"s� 1`���<'XD��F��Px��Ft��%��=�)��'��u��P�e����e�ʨn�R��č��8zHZR@�6�I�G��<�yR�߲~c�J7�H�B�r�p���%�,�3.܁4S��(@&�'i\Í��>!"�?*!xt��t7&apfGuH<A�ǒ=�x���F�yɒ�X!�Ѡr�,��7Ƙ:9j��$ٮU(Ǔn�60v�ː4�v����"<O����``� �(�*u�������s4�˽p���[@
/p?�(�'�ɣ�H�O�b�A�`D�j?�|�J>A�hT�*��}�6�J�<�"&�Ӣ�)��,�~=��f�.{ TC�	��Y�ɺ���SKW.0�.���爕{A��yT!���� g�2�g~Ү�yq 4�(@:3غ�������yr�Ug���ɇW�Z��e�K?GL�Sq�ٚ  �}zѣ՟�y��Ԝ(��������) 9�@HB���=q�*g�H�7iӉyQ>u9!�X�$N���(G(\ X*�"O���$τBF�l�.>^V�bD����U=��rf��|�
�|
�jI.#��l�P���|[j�a4
�b�<I��
�Q�0�@�_ �|��'F��q�A��S��y҃C	L� ���;x��I�Ǔ��y"���h"�&[5{�N�����D!vY��������b�P:��0r��+C!���b���C`���iq�R�!��l��l�1N�0G�&�s (8[�!�dvS�	3S��$.�=
d�C�I�� y4/L. Аuy㏝>Q��C�	!B�j��*o=X����Z�ka�C�	Y�15��&,�mCCɗ�!�䆆e|�sl:L_�5RŴ�]�!��^`���G�NT��1�֞C�!�@&e����2	!NL}c���!��4���)�Iժm���r�!� b���	1�T� c���!���~�<����E� �`�0RdG:�!���F�j`.R]����*Q.�!�F��f��f����1*ٺ�!���p�Y�튏J�$ԛBhBr�!�D��G������'F(iЩO�	�!�$�.h#�A޽&���yc(V�=`!���8��� �K�^�x!�ə\v!�d�)�*�%.��ZEbB�a!���Qe���Ӎ�*e�6-@[�yK!�D�2h	�I��E�>�|B�lMO�!�D�'�	��]����
*�!��]�6{RCdO�*IǢ��J2!�d�"�jyhd��I�=���Շw!!�dցH�vԪc���"���ϐd!���#T����wB�7�$L!��љr�!�Ą�������.#��)c�	�>qk!��S͚�j���%�R���Oƿvp!�dK=&>��Y��E6��p�`�_
!�� �YP� �'i�6�z�)��_tz��"O����ZNUn���鍮Er]�1"Oxɲ`a�+ppI���:�Z�@�"OX C2��.�Bq1O^n��p)E"O���Ч]�Z��蒣A+7�0ݩ�"O��Y�aI�3��LdC�(��a� "O\#c�Ģd�E]T��PA""O�8�E�
l	�G�	<�vY2r"O��;`�~0I���,�4�y�"OY�g��ʸ���#,���i"O��V"�!q�8��"��;	��"Ox��aȓ�r08X"�`J���̋%"O���0b�S�0�£g�nIB�)6"O*�#f�{�$L�Ń�|�d� �"O��4�7.un�*�
��l �7"O2$
�h�h$�,�1I���hx"O�	V�Q�d��Ӣ� �^��"Ohy��"
g1��f
��lA��"O-�G��-e��x��%V;����"O u"�.�=�DI��ϰ�慱"O�����}FZ丁��/Q��e9&"O�y�S(��w%���Ц�6��b"O�L�D��n�|�%�)F�z�"Ola� l'7�Lz���<��-H�"O��kf���3H��Z�i�
rj��"O豫1k��Ft�7hI�D�ā�"O�l3�'+/	hi#(S�16؁�"OB����Z�Y��\�V/݋�(��"O���Qʌ�e��e���M Qk�MP1"O��p�[�2�Q��>����"O  �`�_~?N `mJ}�R���"Oj��&�2S1�E���_�$��]��"Oz=RA��Iݴ��S-2Cd10�"O�a���SH1�ܙn��<� "O�� �+@!i�f}�#P;!��Q���	}A�I27��>�Z	�v��m�6M�:�(��ͭixV}pv"#lb!�䕻@3�b��_nX���t�W�:T!�g�D)sV"D ���#D)EF!�$�8}��J�`� .��P��ۣb!�D�i��P�'����q���'Z�!�d�}4��h/Lq0z�ݸm�!�wm��1��- �pA���[�!�Dڋ.�-��剽!��Y�$Ҁ�!�$Y'&��kC�z�.�т%��,�!�d��w�XJ!�:H�t� f>|!�I!=�b�4��xXS�Q�g`!�D�WH�A�Α�Z��	0E�-VA!��;�|���IK/j��!E'9!!�+9'�<Z��>�(!BjǊA!�K�j����T.B�LY��Be�!���T���ec�<���
'��M�!�$�?�(��&l�3�|�K6&�-n!�̤\��<3*R1�=�r�?T!��GY�5�r��,Tp�%)O!�D�<�~��P&��[!���'"�!yN!�� M�05&�A.�%��/L!�(s�<� ��@�bn�042!�$��bp���F,�V��C��F!��ԁ3�6́)^�]�L��-�85!�d��U�� ��B�A��|��fI�KD!��9@�}��R4Z�2�H�ID!���9d@E�� ������ݷG4!򄖜F{��ٔ��-�na��+K/ �!�d3T�uq-`����'�6t!�� N͛�����H��W�>�(��"O����$�;T��qs&���	U"O�l��G�z���X���/K�	Ba"O�h��Hآx�ʱ�* �Qv�	��"OTh( &B�_��I��GQ.XS�"O^Lk�j��3M`@�* df� ؃"O�PӅ0�p��W�3�T-�"O�]q��U1֊V|ln� �_�<qkA,X���0F��+U�A��mJu�<هalwL��H�$AS��V�Yp�<�5�X�4�R|ɳ'��F�bP"U��D�<� �
���U�S�R����IVB�<1�䃮�Pܱ%g��R��]�F�Du�<P���-�����dT-u6��G�z�<�i�2��{��-��{��^�<T��'~N����[�,^�xxQ,Rs�<�5&P�Q�px�c�K���yc�Pp�<�b*>B�z|P(�<J6T��mDo�<a��IoM�e��K&R��3 �j�<am��u6���%/W�k4b�kw+Sc�<!-4Qv��R�T�"Ev4��_�<�F-߅,X]�-�Ib�.Br�<y�J�[���B�C�/:RPB�&Jn�<a��4TY���D�=[9�P�E��i�<�A�H�~���բ]g��tK�l�<I' �?����`'/�k��j�<�ь�i lC���.��Y��Q~�<���ޜV;��9"�.(�l����Zv�<�ԍ��Q����W���溁yR�Q�W��pr�k�X�H���S��y�8����$�7QN���s���ybmПt���ہkD-Bf��� [�y"������7�˸.L��PW.߰�y2�˾� )B���-��5������y"��_���0���1��yT���yb+�A=su�+4���ӥ=�y��P�d�d��*$Cv�8�S���y���j��d��;%�x=�3hW*�yrF�C",�T�e�����yR�Ʀw��\�a��+Dzd�WD��y�$�R��n_�b8��O��yr�ʖچ�ȅ��=`�b�Dʤ�y G�#��; ������&֚�yRo�B�1r�ʗP4L��.��hOh���dj�HQ���n�XÓ�܎�!�H�O�kpnI�<��,6�ʙ`}��=�Oj�V�
���8g�c��': �%��
���Lk��D���-��$ɰ�,D�piWc�Tr��c���#/��*�)�hO��
۠��q�ϫR�1�����\B�	9e��-�e��-q�܄ꂬ�� <B�	 Az
�ЋS9V��T���ߞevJC䉔;����(��WK���!��>D�B�I�$���9Չ��Xy�wB�V��C�I�AH^$���V�@�r�1��ؘǎC䉆�\5�� ���2ա��v�HB�	�E���"Vd�K6XHY�C�	.B�%~� �V�4'u�E����B��N�
�Z�*C�|��t��D��	�B�	3B���W	��y���+���B�	�&�D����TJ��2F�ܴr�0C�	�L���'�?N�v%��.0� C�	=n��gS8cz���@X��C� #1uҦI>A��z�T�F��B�)� ja떞.��Lz��̻S����"O�d�v�ў,�ޙK���Mx�Y�"O�x�r�?�δУ�&4�F�J�"OnL�B���@�$Pj�BU�7��b�"O"�
@��/T�t�Ra$^b8���"O��A���K<ZS���'��s"O��i0�ݙMw��C��
�a�ꀑ�"O��b)/7z��� �N�0��"O}����%}t���Ζ9m*	�U"O������B�>�L�9�"O� Z�.�.|���FD�c�s�"O���	&!&(��EE%#�*�za"O$�`�E*s��Ԧŝ'\�1ag"O��BA�D\[�)�Ƅ�lD�Q"OVh�Q�,5_p�P���Q�(���"O��kczj��'� W*��R"O�]��ɩ|�>�����2DMbc�"O���V�ť)����١W�@�U�'��''��J@�]~S��Z'�����X
�'������3;�J4�qX�px��}bO��O�Oh�zs�����B(�1X��=��'�x<!	\*@��iIF��8R�f�*3�,��>�(t�����ɫN��G�Т�Ї� �Vd�vmДN�^�5�!*v�] �ȁ@��M��P	����?.q�`��5�zĆ�	 y��vf&?9Q-�sݶ��4,?2�LɸF�k�<�Ϛ2bY����AǸ%+,Bc�^�r�{��ވ�ȟZ`zUL�d3F�qw���tr�"O���/��<�0ѐQ�V+.��1q�'�'R�|�'fN�A��U	8�p���n'@c�;
�'�!��G��<�`��0�r��ڴ�Pxm�!(�z� ���9� �N��y2�Tk��H��I,'����&�yB���A��ޤQ��I�ҬF!�yR�X\��4{u�.E��h2bQ�y�f�)_RZ�x�ǘM���q����y���INraF�(L6��qDo���y�f�[��l���>��a��"ݓ�yr�BՔYq2n8�E��"��yR�"u3�EǬ*���p&ʼ�y��m^j��h��#ٶ��d��yb���S�t!I��+�2� ���y"� R�$���񾠡B�y�̔6�8��s�	�ֵr"FU��y�l�n�� ��8z���K�F�#�ybd�q�0a����*GV��L(�y���
P����.ܚ=�REA�����yb)��{G�}r7�;!�C�f���y"C.�T��g73z9"��y�4��I&^�1k��ǡ�5�ya��`gF�sҊޭ#T�x�����y�R��}��#��ٶ����y2�.b�Π�ɇ ��E�3�y��U�B1�p���B:U���5��y� Άi���!���Nt:��׸�y���t���'鑝�A�����y�m�!�H�:R띻=vN���g��yK �Gjڥ* (��c�dcFf
,�y�l�,.� {bgFzB�1����y¥R-�jy����ox�t����+�y2�AM��qi5ʕ�����dQ	�ybJK=H�m*�Μ�^��z��\�yB*��~��䑳.Ҭ[%�ٸr���yb"�&Sǎ�#��ҿY�:q�d �/�y
� RT��D�5L�5�b)��K����1"OF�0��ƅ7Q~���%��bH�S"On����W�:�cO� �����"OԙZ��R�/��X1�\�`lb�e"OV9�e@<���c����d"O�����%e���d����Bs"O֔�.�
d&�x�� 1B׌11"O�1`��5M�鋰E\.A�XR�"O�$�1�K�4�����5!�N��"O�9���2�,Eʠ�	n��(�"Oz�ك���XĖ!S%�^�f@��"OB���PW��P� n��Cx�p"O�P�g�::�(Z'��+{n�ܓ�"O�iB7��"%��ҶDN<�e90"Ot��5eU� �Dx1IY3^��M�"OF5*�Õ�bM�A��-��G�L��"O�-ST�X3t�*�#!���$��9�"O����Ql��g���d����"O2���%a��y�J��^2yS�"O�}�aE��9n��e��O���"Ob����ԜW��d0�l�9BG��7"O��`LU;
x9�k5@� J�"O�L��ܑ4�d�)ӪQ$`!�G"O:8`뎨:����_�n�d��v"O��)�͐�0��$�e*�/c�4��#"O�iS䀻#��1�	��v��Q�g"O@�r���FzZlc��O�%�B!�"Oz����&�)���>o��XC"O�e��*B?DZ
��g�E��=�a"O`���ԙ��e��J�"��O�y��Ƥ1%�0c���;Q�.-����1�y�/�r��ے�E3E���i��yr!F>�.���g�DEx�Y����ybN+K�hz�M��<J�Ru����yBOϚ� �$��b��E�P��yr`B�"���I�M�v��,�yb�	G�&�b��H	S�*A!��yb(?�d�c�I<P� ԃu�H��yRL8Z��Y�gK�d4����yr뇲$ T  ���0)������e�ǣ,yzqZbk5D���BԵ_1Z؀V��+c���A�2D�����eMVzG � �Vx��F0D�̋�̗\���5��:��4�Ѫ,D�$��݁TN�p�J��wn/D�Ԙ �}`mɀ&U���<Y%C.D���GM�!j�Bè�U�Jpq B9D��
s�� ������> 6����8D�T�4��9Hu��k��L�.LsE%<D��aġ�\ @Q3�Yt�	�'�7D�x��Bّ@Ǭ����O��|��3�7D�HZDO�/��Ԁd␎<�T�j6D�|�Sf�ty��gC������bo.4�0�Ϟ
yg�@���Y�f��r&�U�<qc�߾?|�p[3/* 쬠U��E�<M�}�� �ŀ^����F@�<�%���P�ie%G9.W`�%�}�<S��r����V��CE�c�j_d�<�Q΋4gk�Y���ˑa�l���.�b�<!���5)8�	CuEz,���6�Z�<�����p�i���
]p �r�B�l�<Q��T� b]�V�	?KnEHC�k�<i֌�=x� `w&��|�hJQ��h�<!#�JD�z��dϸ2�^����N�<ၮ��'�N��ھK���AM�N�<4���9��HD��W��_�<i�&C�{x�X��`Y�~�ճ�[�<!�C�6�^|Kg�M�0Ǯ�6G�K�<A.�(`
����R�AY�,r`��D�<�ER��8�����	���XY�<�'�O�+̂���\�R� �PS�<��e�,���h�9V�����O�<1�l�x�P�@�4O" �d�I�<�E�%��\�/�-lb<KETz�<�4GZ7+�j�Y�i�&rܒ���Z�<���Ҟ9�H����d�r}J��k�<YR�`�� P3(�E[�xzj�a�<��	жZ�8����̟�4����D�<�w�!?[�U*g��pv��) �~�<�b��6��`��_�U�>i����v�<Q��='B��aԫe.4�Xs��p�<Iր	��ȨbT
�y&X!@�ITm�<I��X ��׊�� >�x@ހ�y�	9�(I���O�wb�uk���yR$@7"������Z�~\�8�M��y".B/�bPb�$ğf��	(�y�ꍓX�̱)c	�[���T*�y2�kr�����X�j�c&��yb  �F0F���mM�IA� p��Ha�<�b��V	ˢd� {�T��%$Gt�<��*t��i�� P�M!S��m�<�!ոg�YYq�A+R`x�HC�<I��"Y-vax�T�w�����v�<y2��q�,B�B6[�����+t�<I'�E�x����h��=-�`+6D�� ��k�g,n���v�R�(`"O�Q�e��?$ʼ9Q#ҞTzn52%"O}k��|�>��LI)a^�`@"OtA��ӡx���
3u�J;�O#D�|`5��x}aW��Mw�d�F D�0����"3�69�Aa�4}ȸ9�,"D�4c�I�%��� FU����c?D�<�b��Y1~�v�4P:��b�@?D�D:�M�6-��qmM�u^��7N:D�t�,ʑQ����v(˾VR�/�y�"vɪ�S ��#�a
 ����yҦ�������/ń�X��B�yr�Q�׾�����)���&Č�y����Mh!#!��q������4��d(�O2����>6��}#��9�pa"O��yD� 7y&&���B�p���"Oư����|p�{6������"O%91�_;�x�'��=#f���"O"�r᫓z�މxs&�|�ȕ"O��aw��dD�R@�@�x�ʧ"O��#��[�ht��S%���[D�|�'�QA���:9/@@B��%Y�!	�'��I0���J�ܵ�ѬX�PU޴�'(��7��0-���MZ�r-h�9�'�i"c%�~� �AՋշ�=��'z0�V��E1�Bt���BH���y���.�viJt���}"�`� �yRE�b�zAk0m٘�,��JD*�y2��2� uӁ �\#@�b��W�y2��O#��A���&H��I�&S��yb�ѝbj��� �ȵ|ډ#�S��y[&_z<#�+\1д�`&"��ybO� |�$ Iqi��ٲ� �9�y�u;�R���1~l�Y�u���yb�!ʠp�r�n�`q ��M���$&�O�^	JVY�r,�!y���'@�{�<�4��ZlY`l��30��r�g@u�<1�C m`\��E���Ȋ��y�<�R�L�}ͤ�r	](p��qJ��
`�<�3��=:�Y�b��&yh.ĢB_\�<Yc���Y0�ؗݛb0HR�`JB�<) ��T�PK�	ѓy��,��E�<!��H�O�4Y�F�y�X��@d�x�<��k4�Y���χD�����|�<�5a�8�R���yd�-�獜B�<y���5H�]SwEޕ6?B��.A�<i �U}�����N%-,a ˙f�<�p��I��@t ��A��Jh<�2L_8�� �і�
�����y�薌"f���1n���V���ˇ��yц$�b$!���{m�0�倆�y��E"U�b��R�	�d��|�a�(�yBG��9���t�Ʊ0��)ժ��y�ȣ1�4H:W%�^R�aYA���yREӦR�j!SC([l����L��y��j� ���h&P�^!��@��y��@�<Q��*]3F����"ǚ��y�,[�+�V�X�]7�R�#�Eۛ�yB'&����@i�+P�10�V��y�َ���Z��W6�!�W0�yR☢-)��
$b�/>���/��y��xn�s�/�:!�,��FS#�y�	bD�c@ɹ	�npa
0�y��o�lh!�u9�IB M[�y
� �P�4Cp�ɉ���2R�qZU"O� ���	�2lbn��Q) -x�"O�`	�O�L�8��GU�%"O�Q��/հ%��čH"A��y�"O�1�w
�B)n%Is�C2q�8Љ4"OQ�p�$a���c�]0�&hIp"O�h�c@ْnJ2�a�^�D�Re"OT���ҁ.�R�[��*{�t"O@�JBʀ".����OD�[��a1!"ONEƏ,br]y��\G�\��e"O ���+q�a�o�F�ʓ;D�� ��
I�t��P/ݍB����A
9D�,�C��@%P�Z�۸ax��p�:D��!+RU� �����
��H9D�����|�� ���*�* +�f8D��Q�F%`b@Q��H�PiHL��'$D�8� ��+}�1P��E�|����� D�| sV*J� 4�R��y�PR��*D�t�r(�){d@��8O9l�B�=D� � J�
�:X�� �))�X0jQ�=D��	�E�q��(��i:;*�FH7D�$�B�ʵ;����D�����7D��Q�l �T�ŐY4��a3D��x`�́6�:���� �c�X�!�O>D��@C�Śk=(=[gM˶P,�S�?D���d��9i�N�j0lH��l�3D����(�A%�DxTlD+AQ�|�C�1D������<���A(`�l��� /D����hJVl��柖]ܚ4�+D����o�0O���	r�]%@@�<�e�)D�h�B��VdV���	�mxؠQ�:D���ˎ�X�tt2��5F�H��#D�!�OP�f���Dr�,8�&>D�h/�+|�2�0f�A)���p�"<D��cH>Y��)X1J��as�8D��r!+�\h����>���i;D��Z�-0g$��*�$I|��A�9D�� ��H5����*�� pfe,D�l���Ɓ'�R�eZ$$�|��"�4D��h
��������?_d쐆�3D�T�-מC�v]�GT��L �=D���3cT,Ok��p���k}T,"��-D�(
�h��H�V����P�jqT����,D��
��^�u�xc'� Y�,P�V-D��{b�B�;?���#/pް	 ��6D�, ��I��)���"D���3D��h1�\�.�*�[V늣2�d�`0D�h�Wdƞe�h�2�bjt(�/D�ȑVe	c�r�l�*����-D��'�$�����"I�s�}� G-D���o��H�����
C -D����H\�l�P��#l�!N��09�@+D�,����U"�� �#{��j��(D�0�`�=����$%Q�\���&D���w#�5l�����N0l���q�i"D��(A/��yP	��@:n��JW�:D�����Ra��}ɶ�@�^���F9D���a,Ӑ*]�p�[�gtj�;`�9D�|���,J��T��(j%��8D�@�� 0A\x��L�)�YQL9D����X&{_��	W��e�8U
PI9D��3L>O?@أ@V>
"X��a7D����)��3� �G��2��<:��)D����iB�F]h��@���J��vC)D��  I�qNG�S�#�� 0+��"O9�F.�,�aAU��Y�"O8�{��YY�ބ�ǭ��u��"O8!��f��#Yb��s놐c���[e"O���I&)�
��ԩ��5Ѯd:q"O<���EƇ�Q�Ti��5�R���"Of�Jum	�*�|S	��@Ÿ���"O���f/�$\��@昀?҄`�"OR�� \٘�:�$��64!�"O�!!���6�=��ЃQ���ۥ"O��wgƠ? 
���Hӫ=�<u	 "Ox����WP
���sܴP"O�<CG��X�w�ŸSl�R%"O�8���шZ���s5$ON����"O���VJ٨k���/��xѼ���"O*��J)b}��bRo��U��x��"O��C�+����q쑆Y;l�%"O%�L�1p30Q�d�]�;(��a"O��ڠ�
U� �8�ʃ�q�&)�Q"O�G��.�x�q��>4�ye"O.x�b�}����H��yR���"O��J@�&2�NT�F�G�<{�"O�}Iq��,���c�:V>Z�"O��!��0��`K�A��SW�U"O@�[�`ƨf�L�����YNt耇"O�`r Ń7�\��+݁YK8){2"O,��V�ߑ;�Ĳd̒�I��1��"O��Y���.ɞt�vj�1#���*"O�Q�Gf�v���O��c���"O� *a�3m������(_V �"Ol\X�g��a&"��G��Q�����"O0��`�8CwDp`����T�NX�<�3o��)C��z���#d���aA�O�<!D�(R�B!�g��dP���J�<	����j�������/���j F�<QAMQ�<�kf9V����!�f�<�5FU	MӐ���		Vձ1Md�<AUń�t]~$1%i�T*$���Wf�<a1�(��H�̑b��XC�_F�<9��W
&��Qᴭ�\�>����CH�<a�gʕ��!��%�8�8�D�o�<�����H�E I�>�a��Xo�<чA�i�ƔYƭU�v���_�<!׏��\sb P�MK�:�3#[Y�<!gcܩ�N5I�呲�ś"-W�<���Z�"2��H�T��c�/P]�<y� �k&�̓!��q���Ba�S�<Ap�����{E����
���M�<iE��g�H9c�`B�+!��t�T�<�3G�LWF�����V����UP�<q�
H�F ��#���h�@8�4�VQ�<i@��d�hE��=+�j��i%D���&Μ1Ԑ�� �>]���q�?D�H`�K/z㾹��!^G�r��?D�$3&��(s����B7j?b���=D���'���"�V%
�l_�Q���)��9D�Tؤ���B��Qr���&C�����5D�0*0�� 3֪E���Z��H�D�3D� �1�܀rɦ����_�b7���&�=D�&��

� !�I%h�����/D��a�,Cآ%���
�N��q!D�<��޴:TFd��Q.6}n��ł4D�p:F�-1��Y��dΔ\< �6T���6
�(U�(5*�]�GL�1"O� ��;��B�:AS���2�±"O<���7�z�R�N�0ȼ�:�"Oh�Hf�ƑQ��Y�c5��"O��`ؖ_BPc6m��E.�,��"O� :���
3AY�Lˎa�p�"O�=
4�!m�H)��77Ｔ($"OJp�dK�*j���x�g+*��	J�"O��IV!A�Ήb��ML�m��"OR����W�h-���X S-<�Q�"O��d�Ռa�hܲ�a�'G�A�Q"OV�0��U�0P�f@O�4 ��"Oj}�P��jB��ۥ� x\� C"O����4�vѳ�oR��5��"Olu@����r��h�	 ����"OVa�_j`ppQmT�~��c"O��&a���er��; ����`"O��Qa)��!f�I(׭�AД��"O^�zҌ�*�ީH��5�z`�"O��ʐ�}6�#�@�p�^��f"O�`��W�j��5����溁˂"O�lA+}�b%ɵΏUCVYAF"O�Uw�R��	�E�K�S��� 1"Ol�hD(��6}
-���r��C"O�h3�c��.�,{�K�`�	�"O$d�!�1.n�i�0�N��Ĉt"O��c����-blW�<��Ƞ�"Oc���',�Y��W
nL��
7"O@9���#��{��A a/0�
�"Ofy������j�NH�f�`��"O��ꇄȮMu��+�CM�#��ye"Oȱ@�aÚ��h�-��Q�B="O���k��f��{�A�L�½cG"Of�┣\�1K���pa+ pAX�"O�A-�ARl4�A�	t��%"OJ��r&�2l�$�#���j��"O���M��R`@�D��u<�L��"O��1t���>��(��)�d�:�e"OZyi�ϋ�����a�"�zd"O� �[T�D�r������P"OZ�:�����U��(Ixñ�"O�L`��:x.y���ƴ'uB�r"O���.+d�8؈����@@d�4"O�����
D�ȳiԎ.@��"OL��aNϹ�����-�6i7����"O��ϔ){)��SDlD�ZJ  �C"O���E�a� XT���V���[�"O�h��N@�`𜓐J��9��H"OD[���0A\�+R �2��hp�"OXt��KK�\"��RnҏgY���"OE9�#S���y�bl�^C�ī�"O����J�k>x"�
D�R~��""O֝sL��^ؤ�a�fE2d	�V"O��,\���ec.~Q�Q�K
�T�!�ݑ2C�0K�!�a�ƜR戆.[�!�$?$/\�J�׷�n�T����!�D�he�ܳ�˄)>�P�TfI�,!�䞄S��H���Q?*i�l2EoI>�!�8T'����"�R��i�v.�K!�W(<�Ph�@�Xy�l)b�E�!򄇖v#(���iȀY�R����M�!�עoXάBs*5F��E���է9i!򄔭rKp̲G�Fq�.�  XnJ!�1`b���cˍ't�]c����N4!�d��V)���T� ҂�HV�j/!�� ��������'m	>���"Oܡ´&��K��8$�02P�4"OƐ@��7Gw��)ʂ��fm�"O�f@@�]6.���ލ3��"O@�:�A��V,���!H�ܺ���"Ob�+ֈ��8!܁���5>�0 yf"O�+m��W�$���(ɒ`w��A�"O�L� ��"�v��@�Я7��1�F"OJ@���Tg��c 0gM"Ojë�� c`(��
[�L�*u��"O���E���D��!+��V��[�"O2�Xg#!��l2�"�5>_V�"O��FK� �i:c�N�`Y�}��"Oj�E�:!�DX'���W����"O����eҦW��{��5?���"OP�#��L�m�I����Y$���1"O��z �לGIBM�uo�B!�`x`"Ol���"Z}��`�nI~��A�C"O�Y8�=d�~S�CO?k���s"O�$��M�Zṟ��"�~טp(�"O�p)W�сnW8P���Cdn�Ö"OX@��԰ײXX��X����"O^@G�H>���ږ��G�2A�"O�q�jZ�`��-�P+�6rDM�Q"O��A�/��/s ���T�SQ99T"O�0����+x�c���K��B�"O���)�g�1+`�|z�"O��@_*<U���)K��+��$D��;��S�R�И
2�+d�@��M/D��`C�N����u�(_��)1�h,D�����]%^?�bG
�Y�$�2�/D�ı$P�L;pH#n��\�^`Y�+D�$yU�)o�4�"n��D�G/D�@zvh�`� �`V&�)A(���/D�p�F�<*��b����O"�%�G�8D��˅�$��95K�3!*�a�u/6D�������s�j)B�h��(��3D����Kךja���4�C�<P��"1D���qƟ��,�a_���t�0D�Јsd��
����ߐ$���7�+D���׫ʷ@��#Ԟ��'&D��ɐi]\$��ԡ,�~����0D�(Ё���<�����R�f`�b�.D�\@��J�<�h�[c�"y8t:��,D���`E�;7e�����;c�l�n*D�hB�eq�(�ɑv������&D���¢�H�$���-W��$���$D���� [�Ƞ[��O R����'#D�`C�:clh�R��s���e6D�ġ��2�>(�`L2��c�l5D���b�0T�)���*Ѕ��'D���So^����r`OƗj� 	A#�#D�0!��	6��Ȳ���, �c%�>D��jR��3(V ���bYN��PPr`*D��rweJ	z�B� �ɉh�����*D�����^�r$�1��6��pI7*OF\)�oԀBz�'�بW��"O<0	 !U���*���uv~}�G"O�$�'G(%G~�a��X�|a҄�"O���G�x ��pgP~��$"O<�򵌜�]-j�À#��@��Q�"OZ��ag���8���rP�:�"O�3g�;R<�"sЙ8���""O�	��FN������\5����"O� ��
�'��8�*�i��+"On�h#(#h���b�į\�b�A"O@<86.� �����C�Y�q��"O��K�I	�^��(�VE�G,N��"O��T畽I���C��:̝�"O���4�I�u���@����ޥ��"Oة�5�\�z�������[� !��"O�Tg_��h��1�`�Pz5"O�,���Ǽ�%h˿K�	3"OQZs�5~�4PP�ϲ�8Đ%"O���M�68�R
��Kj�(s"ORD��BξdjH�*W�Z
uM���"Od���MP�y�'QI�l̡�"Of��4�����('���l8"Oh ���>c:!+C� ���'HDI2�dʿKv��#����<���' ��I3'K�@$�� �_��
�'2� ;��3MU��ceC�^�h
�'x�x�5 Y����ԃ|�p�	�'��aģ� q�3���a��*	�'��<�`�K�9ހ�Cd̠]�q	�'�J=�ҫ (�U�#�ʯ 7�e�'It����o��U�硃�f<��'Ď��AF/��HwO�)_��ܠ�';hP#c�<:a��)7��?R]���
�'�xm�&�/7�0��C�4���	�'lc���o*5k�j�2-�`QS�' �`��,��ٹb��'���'դ͈t
��XZUp�X8i�n��'�̬�t��.g�ʩ�QoG&^�б)�'�B� :7��qa�ͨ\v��'T�bm̑iAJ�Ȁ�PB���'W*c���'D���I,� ��'-����M/ljp�I?	�:$i	�'�.0�S�S<r�̙�kt+b�`	�'�N�3`�ؤA���D#��4�*h��'�T�ZQ�Eu�<%��iR�,.�A��'!@e��֋X/
�)��H[�h��'���æG�8�-�R	�N[�\@
�'٦ؓ�Ɂ�$���r-��VτE�	�'V��(3�ٯ{�J�%�аTF��'��-��=>�Pc#F&7�j��'B,�6'�.pxi��(p�'�L$��
h���㌋'�p k�'�p��:0��`�@_�!�Z�[�'�hr��I���b�.~���'�4����٪&�8��\�x�]A	�'_P�-U��V�O4�Y Ek�(B�ɞ4dp\y�
A�<��Q+p*V�t��C䉖%p� ����*�H�-P��C�Iu�uK�GŅg�(Y��	�5?NB�	- @Wĝ�XdQq
<�,�	�'٬��e��1��}2��:u縅	�'������RxL��w�ܭh`BQP�'�^	sDk� $��͛+g���a�'�p���\�4Z�З�o��ٰ�'��qB�
�+��% g��n.�I)�'��YA��
?�����(0�"@�
�'мi`b��{>���c���!�v�;
�'���щ�8��HKд�/;x���'ˮp���F/���7�	2+�$5[�'�v�t�C#�fQB'��9nY,��'9��m�d
f� G�9i{ƁK�'$�����,kvt�Cq�Ϯ`�hI
��� �!���E>���c��*�� p"O���P��xa�7�j��"O�zgAArr}�u Գsc����"Ou� ��^u���)D�$h#"O.����ǫ��:⍒#;���"O��䋕�8���+�f�m�L\A�"O|�`��]���eRW����p��"O�Հ	YB�&iK�h�4A���0"O���`#�&H�9c&ӺG�@�"O�l;��^|#t�A����\���
f"O���#�'ONlu")�N��6e/D���GïZ9��ؠ�?d��C�e.D�°��*	����Q�A�-Q>�!�`8D���C��$;$�`P�I-'��y�G;D�p��Y�>8�4�@����)sC8D� ��
�m������4ԝa�8D���*�%-��#����g�Ν��6D�X�C�B�{E.J@�V/M��cC�6D��/
�U���A��5`�*i	��*D�h(2�Sq>l��̋�Cb��9'�&D�@��oK��x��F� U���a��#D��ӡ	J)��<[e���q���3%�#D����֮\Y�T(݈_��A'� D�{\I�2(4M�;�ĠS0�?D��9¬>�0˗(S���;D���m�$'��eѳ��$�ؼie�7D� �d)��$�P�R&�.'���@�4D�\Bs��p -��Kz ��6�?D��:�ˍ\p+��QM֍���!D��rf���
r�-0Ä�>��QC.$D�4pA�C��MXpa+q7޹J@	.D�T9�['ڬY� %�:u�e;gH&D�$R'A�F���XQ-s ��K1D���O�;�$H��j	�bO�-�3�*D��z6�A$.bHK��u���&D�0��OیF�l�q& ,b*�[��7D�P�J�`�ej�F*lJ�E;��5D��p��٣t�z@� l��d����6�0D����$�D����`�9#���I�o,D�|`����qn$���'j� A�<D�,���H�T��-�&Ɋ���-9D��b%�	1�h���Y�
 ��+7D�X �,���X�5�Y(i0�{0�'D�L8��D�����^���R�(D�L�Ǆ���X���=2� �2u&(D�DZ�!B�n�r ����D��2��3D������?ZB�u��H���f��46D� �@(��X�8Ir!�g�3D� �$�	g�J �X{�
jsA7D��j��@K���P�C=X5��05�*D��b�ҧ#cީ�P'��	��Jr**D�в
M��z H��V�,`��d'D�xy�HɻZJ|0h2�N��X�*!D��	t�Ȍd��(VI] ���t:D�8Ȥ@ D:y����?8��-@�3D��i�%X�X-  2��.�&�Rs�.D���V����L�y�ަa��@��� D���E�ސW������|J��"�?D�\�4�]//϶�����7\��V*O:=R =��K$0y�qw"O��-\N��1B֑Q2R���"O��q�H����xE��Å"O���!��m����6�֖Q�N�[ "O$aRE�� #wu��I�@�4�(�"O� lD���˷�M2l
�[�v��@"O�<+t� )[f:�8�G�3��@�"OH�)%̋-Y�YʷfB<���SA"Ob�J�O]�T#�03��[{�~)�v"O�����ͧ`��1�)Pu�����"O�y1A�@I�򰲧���F�z�"Oz(����P� Z*K�p�q�"OdA�g�6ya�@�����0Ģb"O!�7	�;:/ր�5�O���g"O��v��E�"�*�LħkE8pd"O���E�J�fy�()���#y9�"�"O|�B %�Iw�eLD�z��"Oژxb�:p�L:�j��+\��"O��Ye΁)gخxzv��;3�t�"O�t1�mU�#\�9%�c!����"O*���A"x����u!��̩�"OL�{�膟+ ���O�(M�恫�"OĈJ ���-(`̛�F���"Oj�U�U�S�p��A�8$���"O�	��ME�
Dd)s�b؁3��"O����C�B��Y0�B@�գ�"O��El�i�z��Q朎F�n4��"O���Z�(]Z)�4E�)����"O���J�2^��!�IӘ7��)�"OH�ᑁFH��2E�D����G"Od�B�j�!mXi��k��:b�!��"O�T�0�ʁ_�<�i�*�RI�\�U"O&q	RkTC��@���/%��"O�Ay'(8,���_n\��"O|�ďK�(��g �q����"Ol	8 �P3P���I��i�� B"O��I��/a��IR�I],D����"Oq;G�1:e�����> �t"O�"�	O��D����Z떙�E"O2��_̒�)gw�y۶�U>�y�� /P��2MB*X�d�PQMў�y���3b�%s��]'[�d{��y2�L�D|���!��I*v�む)�y�e��PP%�%m���s�4�y⩂;��M#A��2(Xf����y�̐�/ΰ�"�+�Xc�!����y��	Q�ݡd�̏K�֡"���y�E��S1���G*:��q����y�ς
���㍍.M:U1�L(�yB�O�� 4P�G�Ux�Pp�����y�JA�Z:ݱ�"ԗJo>�*F��y��Q>g8mp��I@�)�E��ym<��1��O�,`��Ĉ��y�Y�,L#G!m��x�F���y��H6r!������D��@'� �yRJZ$~��9˕���6�����	�y2D��+Ѽ�A�Ƒ�{��u�b���y2�ה�1r�Fix<�����y��ޛC���V� \�|iqvFK��y�ݥ�X8�&'!:i�y2d@��f�[�n�91֬��	��y瀗�  �P�HZ"h��Rl���yrڍ`��}���Y�(#�B#_�y2/�5~Jq�C�RX�ܐ��լ�y��HR�|�S� <Y>|\��(���y"#�+HLE�j�=|<����V2�yڵw�Y�oCw������σ�y�	0T�����m���CE�Ω�Py��^�4Y�'-��[���s��Q�<� $-�eƔ9a�9S�φE����"O0��ìի �x{�d�22y��"O��� ڝc������T����P"O8�`�>#A� �� s�4��"Op|afo
�*0N��k�8,�`��"O���ʙ��Z�4|ym��"Oz��E����>	�V.N�,�qs"ON;'	Т�A�E��l�J]80"OLXѡ ,|/�%fX ۄ��"OJ��v�Z#k���BE[+c�D1"Oa�eV�vDA����.idk�"O�\���	�<�f�P*� m@M �"Ox)����K�f|a��������"O���&�*�ک:�nҪ;R�U�e"O�@A��ˌ7iBT8 ��@+P���"O�LB��D̉V�F(Jn	�"OX`��ӕM�
L��\��"O�5��@ӰZҊ�â�>3E����"O�yDV�YԮ%X�#�\D��k�"Oh�`�J9D�[�BAR�yp"OQ���	13T��a�OE���"OP�yՇ�x���D�Ni7����"Orц�P�\| B�ݩgӢ��"O��NN�`�x0�1��r���1�"O�@d���DJ&)�q��D����"O���S���ɂ����(���"OM��A�I� �S�<��m	P"O� Ƞa�:,�9��[�=g�}C�"O�a��Ί5*nAA��ΑG��P�"Ot�Ja��7�j��B��!s"O���r�H�N�΍;� @:���q"Oz��1�HL�+�`��k�@��"Of0p1�5-�^Hӕ�R�8�*��e"O����m�^N���3�\�8�B�{�"O��h��9��8XR��-�~��"O��C�k��~pRqnK�L�P9��"O2��g;t�9�kK�v�I�v"O�4���%XNh0�EL�$cN��"O�`W3��Q2^���yy!�dA��nY��bܩQiʭpWiM�xo!���7̀)XB�QBh޼�g'N"e!�$S�w�9��h� UU6X �&�v�!��#GGXy�@�0�x�	�ڀ3�!�dI7Z�QA�nC�_2�CFd]��!�հ=*�Scd�2#�䋐(Y�!�#3+d��@���z!�LIŇ�3tx!��̈́&d9���G"U�b)˵D��6Y!�G!j)V�B�@�Z����l�06X!�@�}��MX0Eٛl�$2���R!�$�1M���!�� e�� a��z�!�$�K�R=�%�4?��"�/Q�^�!��8Z���q$ś]m��S�NM�!�er�Sb��mM<�8գJ<�!�D�\j�}J� �,W�)���R	!�dC7#<d� iT;��I�ɞ�[!�$ی]O������$=��iԈV�4�!�d�(��b�.O\�y�F�_�!�!��-(ň��F�TV��a#IX:�!��P�]
�J���r��!��^D!��,e�X��l�ܱ����f�!����8�Qҁ��D�٤�#�!�G�[.2̐p�۳�:<*a#Z!��7*�\C��M:7L�G�!�Ã/��eWj��j�<e��d��8�!�� ��AcJ ;v�[a�� BJ@\# "O��Y ���I�����善%<�)1"O.V�)L��bTmP�]��lScmV\�<�"�P,b����h�H����Qf�A�<i6k1LD4�pNH
�JPP��H�<����*FP8F�j2����JL�<A�4�����¾S-b�S��E�<���>'��ۆF�%S��#��@�<aW��A-@|`���,����}�<�G�߷M�<��l��o��20�|�<�G��g<t��a\�1�x(�COw�<I��e|�r�֡�΄[�@u�<��Y,3(�7�NE9�-�2f�g����'vֽ�d���f�.�Bt�u���'^�	�׍�Yz�`tM��r�¥c�'���ƏY�A���i�$v�$8{�'��8��\M(S⒅C�D1�O��=E�dm¼0צ��5Gj�	���1�y��@<T�4���.�E��l8dGA�y��Y�V� I�h���ps����yr��J-0g/�o+0U�U���y�GZBHH��c���$�M��y�B���x֣�,S��QNՊ�y�3E���ԝ%x��򰉚0�~R�)�'⺭���RT~�xT�ǷFU�5�ēM��6�+]�x�*�K�!VW�(�M0D��j��pQ⥱�A�	���`g1D��VM��:*�YL�{�z���m+D�h���,p�z&���_��#*D��A�e��k�j5��E�H_ �Ia�;D����e�F0�5'A:>��	��b��(�O��DâT�R����N�أ'%U�3�|��x�e�2͚u����"���0.X��ybf�$�Sc���h�B5E
��'!�'þ"|%	V���LJ�r;�`G��a��&�O� �m
�z"�h ��3WP���>)ٴ[��d/}2��Ƙx@$�`O]%cB�\��d��m��D�* N�!�ĉ��!@�����ً�'��	�,�)�L>ysb&C.�0��O=W�"��j�e�'{����; ����� Q�J��ҁC.Xu�B��!+Zy� +μ	_V�+@�-Ӿ��dQ����(?1s�T;U\Q��ݰ|m�0V�	W�<1uA~�VDs"M'[�|uIT�D{�<���O�.l08�-Gw'P�#U�y�<9Q$T��F���P� c��˱J̟�'��V�^@}J~&���A]����EN���xs�'$|O�c�p:f�ϰ�C5��G�\L��j#D���槞�Y%n��5��1[ T��"}��O�6-�<�p�r>��?	�ՀQ, �]!S	�	 bN��o D�HZ�i�L�%�%`��-�d�<��hO哦<���C@�έ=J
�"�X��C�I�K`:s���\y��ɇ���bX�"�%�S��?VᚌA>�uKsA�v5l�3�D�<Y6d�%d&��=&���ůQt�<��m�Hw�T��Ô�F�3��s��hOd�T���T	D�~�±�+h�8p�G"D��H��p���7%��+q�?���<���8k�����+"p�h���}�<����>P��q@
c�o^y�<�AC!4d��b		�V�sL�v8��EzRHBA��xyF[4 aRT���y�,� ]�I�e�"|�A�\��y��É<"V�(��C&�I+V	��E��5�O��H10�
t�b%P7�as2�'���� (�� �Oo��q���%x��XE"O`L�r��4?w6`�
退BQ�@D{��iF/�����_�J��MH#%�!�Ĝ�t���#&e13=Ƽ�eN��J2!򤙗s���!�C~/�����4:!�}nz��t��)!����l_�0'�*�O�(ؓ�U(�x��T�=a��"O�<�0�˫B����a�`f�"Op���`����x�P$��3O�=E����!1��X"hF%3�4��+��y��	j"�t���'z����Q�C,�y��)Q	��(N>u��ŲmhK����ا�O1z�ѕ�C9���37!-	���
�O����@��ځ���!t����%�����y���0��D�yI!,N���$*nC��a��O����[�%��d��
�o�N�
b;O�b�,ק����/hJ,}#Q��N�J,�lùu�!�DŶp���A�-1!��Pe
���	Ix����,��uX`I��F�>]�aH�O8D�xr�Ҫ�H��뛏vR��A�#D��0��[;}~��f�u���k�!�OXO~����>er���?W�]��"Oz�#c�����Xr�T�Da��<O�ʓ��S�$�|�$^��zd���ŘO�Y8�G�(�yR�� ?�*���aį{Tꐱ� \���'��Z�S�'OuBU	PN� q��o�
 ��yGz��7��;��
��6�*P�d)�����d쓬y���O��k�"l֬�4K8A&0�h��'��#=E��U|h�K2��+$�D�8e�� �!�׵2f=�dƙMv��Q��(�铅�=�ݴM΁�Q�V�Z�;�*!fX(���	dy�Ϛ :��af�E�Bga!�@���O"~j�iDB��b� '��,x��Uܓ�hO��ǟA�ā�rO�� Y ^��S�>?Y���&�"�Ŋ��]�2���U�	���Fy�)�g}RƊ$v��h:M	6i� �je�F+l)�'�a|�M�+�nm�!�<"4쐸%HQ%b����ԣ=��BH��<�p��V}��§�k�<IV(�}��W��U�j�2p�<u��'e��4qWj��G��_,���#i����h�|�� �r�XZ��L5�� �I�<y	�F�.#�\�q���ɃnT�\� Y��	G�\��˄(��i�&ӱ^� C��86���W�`R�"�+`#�C䉘[x&d�u�S/d��#���ǺC�	P  ��#薞.�)�P"�"�C��n��d:4,��J�)9i�%)�C�t�
�ۓ6ǼA��C�/E���N�Mݤ`�i]�rFl����3����c'��F�#p��熉${2!���TU�����_咹jE�� W�az2���j���!�/W��1���58�!�d�7��!)��K���ʱm�>~�!��0b��D��I���x���B�J�!�$� �%G��w�YP��+w+$]��'_D8����C:B���>qQ���
��~LO�!L,��E�:���O��yr�Ų���[�g��{�X�b�oS*�y��X����Vz�R��V��4@�')�T!%*"a[��z@�P5r�1���' �9㫚�r;�0��,��Vdr�'�j�@ΘcLd-!��D*4Hqh�'ipD2���u�D�R(��8�Uk���huR@�6��g��x8�&�}��S�? �) �m72��i�BT�wX4�"O�ڥb�'	��F"�R�];�"O�u�R�v�z]� �<�$�� "O�D�f��r>dB���h�����"O��6��n�hz��1b@dr�"O��儇1$�&�I /S[��8$"O���#�F�P#�QkWT�HP�K�"Oz؂E��SD���4�	��U(�"O��;@�l�@慖�x��"O�����-1ҍK#�V��q�3"O�m�4-��\�
#��
,riu"O�E���0�2��2��%H�}"O�K �Шql�+�(�;XV^(P"O�-�#�ju<�'��&�p|��"O�X�D���L��d�Z�r�n�!q"O�
R��/{�f��e�YEp"O~d)�H�3���XdJրj?`��"Oj�Z��K_\}��)ۣQ:�C "O��Q����cA$��c��a�"O���
Pv���b����(�ą"�"O���P�\Y3�[x����"O�	�"��}�G�M#i�!8r"O��r�E�&�d:&��Eص`t"O\���J�s{��r͜q���J�"O���̖&|^�q!&��E\� p�"OL�ð-4gXh����2oѢ�"OnH#�E��F�ऑ��)"i�\��"O$�ң��$2�1��A�:>���"O���ǂ֔P��Do������"O�mJ��84Q^�t��o�u�g"O�0�DJ�5.�	�6OY��"OZ�(f@.L�J2A͔{:���!"O^���ȇ3{+��b`ϼ�dJ�"O��j�I����i�L�m}��B"O*�0.Q�|���#a��D,�y	�0{j��I���+6����X��y�W/��}`��6���;�k[��y��%M!:��O� {�D�$Jٗ�y� ���Ы� �oWXl��HC��yR柽gq�$k���z��tJ�L�3�yr͒#ШAW(ϒyh��Ro��y��e�L��r�I�
X�R�O��yrd_C�쬘T�ͣ@�z��c�
�y�a��~T�J�CAL-Ҩ�ǉ#�y"�4_瞸�V��40���H���yR�Տz�p��qtl]8�C��y�蛜@���5,ϼe*9�'C!�ybK�@@���#�[/]���&�]��yB$L+:�~���ߗY�J�#@�����O�����sQ���k�*V�2OB�	F��&f���O(W���t"O݂��@	9
"x��im���"Om���(K�:|�ℽ�P"O�|Z�/�)c�F�1� �N�0��"O8���̕�b�K i=:P��"O��Г!�B�\���LW􄓐"O6xQE���9�g�On>�g"O�j��F�Ju|<�&Y�qoD�V"O.�I��	s����b%X�y[���4"O0tX�iV���WEPr��"Oҽ[g�ϓ{��Q1�`Z��@�"O\@��H N�=Ä,L�VY$�u"O.TBϱ�$��������""Oޘ�e-8/-@�I�e�	{�.=�v"OR�(B��j��	&BP�"O� N�2�ȸ3R�@`�2f��PC"O�+�Ơ
)�0K�F�;}��堶"Oꩣ�H9�B<@"eͷz.�(�"OJ�P𡇂n͸��2�+2�� �g"O�8�C��A�޸�1���"�fyʇ"O�$1���.f�Q㏺C���z7"OR��F씤�核�E\>%�Q��"O�ڐHY2�� �cߋ�����"O��z��z���`� U�l�R"O�Ѡ�m�U���Oq�}��"O��`�I>Lpcr�Rgn��`f"O6畷2,�hC&�f�H�cL$D�L+ë�i.�49�꒵A�N�Xs�/D�d�"�I6�!&��\B�E*D�d��J3e�\���?���ÒK(D�hQb*��Tͨ�	�
ߴII|��&D�����%WB����z���'D��@�ϑ�Y&t�F	�=\�!"�8D������{�X`Ei�^����r�4D���*I�v��5`��Q1h^��Is<D�̻�K�96�*X(P$��8��Ѕ�'D�4('��fu�l���'�u*�J.D�x��E�,���R�E�Y*h�X�B3D��+cb�,*Ĵ���6 <{c-0D���BOc�a�r(��q]���4(/D���q��lɸ�{F�?�pq�A�#D�<�Fc��+�R���V��6tB��<D�L3^�ڭˁϞ��HrEo�^�!�����;+X)g͌� �/k�ar͞)x����^(Z�^����
=p��|��[^h<�eȏ�>`H8I�DU�2�$����o�'����S&��eI���Ճ�V(�L"G�T$j [�"Od��hA0��$�E��p�'�l�1��%:��,�O?�
f�2	�:X:�m�* Z�ݩ�/2D�(����L;�sK�!��񺰋6?����I4�5!7O.�b���@
��5dX%@�X��'&�X�)01$�<  ���pZ�15+D>N�i�3�NC(<ɀN^1Gnt<Q�l(�!�A$X�'��{&(��B'���}�&�ca����ɨ:�l�kD�Mc�<!���Sʖ=�&
)};��[���<!��Y!n�H���C;}��Ʉ��)�D��@��(�@-�`�!�dš�bAȦ��/�tM�gͮI��ɩ1Y���g_��x���dSp!��O��4H�a�<�0?�`��{x<�&(C�Up~�)�Z>$�V���vhæTrz�!�>���4lM�\:��1��4��F|�S���)ˇq6�ɹ�F�~b�d��p�:=1r.��nla`�R�<��EO��(�EO�_%`=(b��<Q�d�
[���u�V!��ۖ�+�'c������78�����P�T���^��c0@Ԍw'�drh� y�%@>@7̈́�N�
9:�����3�	�YZh�9%n�$�.LA�
��V
���d�+��؊CmW*l�]c�c��3ԹsP�ˍ9�x� _�>B����w��}0�aA�;91�͇�az��dɂ(��cJ?��ɛw-�݀f�ߤ%�Z�¤��j�<�t˘ Q�U�Q"��t�C0@O̓u�0#���M���~��⇻%�1�cLT'TNK��E�<!5`�$8��#wkL��^x�d�?T~�xң/}�-���I�A!�X[T�S� ���Ҥ��C�Ʌ�&��r.�V3~l�eJ�; 0�UP,)놀I�i�H�c'@�q����ƺ{�T��lB6}�ĵ`(=LO��A�a<o�� �.]�0�M�0�@�o��a �"�p��(�c������d�^�����l��`Q��)h�1O��H1�k��I��h)R�� �a�M�ӠR ��&G�,�$�(��
��C�I�H��J3M�E���j�@��'�R �T�� 6��Th��s�c�%�'��ݢMs 8CD�@�S_4(� !�� �=󥅲spJ��E�.�zb�Y#0\^ +Wg���T�Pm��"��NLW�'�|�c��	%�b�ڦ�?wI*��W����"��\�t!a��8�R���#%?юu��.���#i�Nx�Q���Q���XsK/�)CӤ8�5H�!1%h�7R���8ӫٮ�!K���!!�r�%I��ɮrO�P�s�H�Dn!�䋅.�k���+@��-��C[��P���2�\�B�iY��
|��BQ>�&>�ݩD��й�m�+X4�z!��IeC�ɼt2h�A4.ܙZ��xq��Q���+�C֛G�̵Ʌ��uM�<(�I�j�i,O�1�O,����}��&�j�7�'i*	��ɉtY<�Q���*iv��Q��'x�cV���]���R��:R�i�' t���V6!9v��f
���.��x��O�Q�\�&�tjJ�I1�$(Ń���:yƬ�KS�- ��(S��M
>ܨ��'��T��EA$|2��%�_��ɹ'��
Tl�7���[(q�����y���'8�S���U�m��	�d��=aKGB�<!�[�>A�Zӏ��$�32�����s�O�3�,}��NS?%τ-��:<F��;���Z�Ь�EIh�p���.���dQt1�X�`���Y���9�ɂ�P��,@פ�)A�f8s#��E�"!�/�B~B�&OB�t+$v4�%�P
@�x"t��t�d.[����EH�K�p+�AT�m�F�'1:y�R��t�f�:�[�!�m��3����7}�pI�i�"���k�&֝0\�e��IǑ7�b�z�J���M���t���L�s���"�#]w�H�c �o�!�7D�|!�M(c�� rG��l|C�axޘ�g& p��1��ēB�Ոd	�ɟ5b�X(� �#x4U��	��A�ӘL�̝(4�EI�*͹�|�Q�G�J�̑b#�|�9O���G���bQ@U�_�m^B!���� ��xK1o�y�� J���'#9l��LH-tH
��Ȑ
x	��0��6�hAV�3N���Z�P!��ŗgOH}Y� Ę�X\��h@�X�}�P�����Ünܖ�x���5`��e��BǄe�(R�Z�����[�4�
TLؖ�V AU�T�^ID(����?�>���U��<��ƈw!�̲g�Ng�v#�ĢG�g�I�u'������&x�>h��	s3�٣`�D
E��0i��P�S�x�7�=dJ➈����@@�)x�*�.� z�#Y�\]��!$�=}�lǳ:��`[c���	�^,	"�LG38���]�I�xM��#<R���!aj�+��0�@�)�p<�T)�&3$�1q�iY���%-�F8�r�S��! �P�G�0M�rN�O:}�Qi]r�mͧ-�L �BS��b#P�V�N`�K�)lHh�@�&O�d��+܈5�\As��>�@i�7Q�2Bߙ~Zy{.N?�p�#���k��[�q!z`�����F�OF�̧#h.xz�M1����*V�u!|��O�ɳ�U�*�Z�P!D-�'c&�U5���h�`ID��j�m�6�2 �-�.��S��M�U�A�t��a`kQ�Uv�z��_�hbW^��it�мs
q��'�X����\'ha&Fo(i�O��Z378lS�W!l}�g�̖U)��j�gUpX�+\�|��\95��0<��*�^��k��]�3���52u�Y�I�����$Pk~���S��Nv8���[��R�aD�	&�?c�2�Gz�韆p�#)�N�'}<(KU�Ј{��h�Ɲ:T����Ox����L�v���C��"�'_��d�SP'}��V�0\+��nZMtb#����K���@�熠O>�(�|2*�PƁ�w�7C�J�HXY���@�>���1��O�@	r�"aj�҇#��"n ���'ԭo/>��R�ұ
2vQ3�FP̦���M�?X�Y��ɠO�4D��8J�,����#H�pD��
�4`�$���muY"�Ò&T��g�N�'X��f�Q�@:&�X�i �PҡG8��i��&�<(��'v\5Z�"Q�"mԈ������ԡ U�fA�C��@I��	/�(���ʝ'�4Mx��%�\a�$�fH �'Ҙ[ ��>���ȃ�D�	���£��hBܣ��?.@���-?֌c���2��$2��4l���J���z"�B6�gı_H�$R������fEru����;c����Ϋ��>!F�P)`�)��%D�/ڲ�B�~�l� \A��2,�D!��Θ)+�d�֍�W�$E���u;���) 8��#�-�y"ă�dS.���[�\p	���_J( ��C+^����.H�i��#�ӳ/��Ε�X*�ዴ�!�r1�U�N!�!��
,��a�h�4(���q�C�*�h����7X�HU��
�A6|��ҋ�
-��}Gz"n}X�5_5{G�P����Ұ=�Fo�(E����*� ��M����;Ƙ���9d����r'߇:$��� �IX��J��e���	a���D� 5
3�,�I�Gc��Q�搢�tݱӢ�71��QrV?�Yӱy�0��%h��"�	�1S�<᰿d���n����ԒT��pp�G����K��+2�<9Q���/��}�=� �h�r���?�$���d�(`�H�� "O�|�*μX��i�� j�(=�E`M�\��̓ej�L"h$���[�I>ғ\�J(R�
0#��<ZF`��I��eȭx�йP�FO�U���D[��h9W��' d�PU!�	 H��d��d\���͂4��<������������3&�y�GF@VW]�c_>-�����D0ӷ�ڄ�(?D�����=C
��Ύ,aB�,pF�qӀP���Ȁ}H��ѥ���N0j���i��-��!�,t�����*.0 (�'�N|b&b@�'����3 M/c���rm��?q�(?�X�Bf����I�r���k�OH�N?�KcI�N����d�O���׫�Eb�)�BH�y����n�e�Z4pt&X":#���$�$�I���p���bC���a~���D�3�D "�ԖYm� ��+��L���j_�g2��ȓ8o��K���S�t��FP�8�� �'�������5�v��O�>)���I%f���ʰq�z�)J D���Ee˾y
08BT �%>��5 5扥>��%�'C| �b� vO:$�1(��>��%��'��uq3A)^P��F��0�<�
�'�rP˧d��ZB�S�P+G�N�	�'��I��'�c-z��ڰ9Ud�
�'����&�&&��\�1NƏ4�X�	�'�����1A
����(�[�F̀�'��S5hI
}{,_^��s�'w����ЗE��ŁQ?�К�'l�����	4٨�"V��M۞�j�'K>�h��M�f	>�p�Q�G�A��'�j,��$F�*S�-� � H8���'���B�П6�X���A;2LN| �'66X0%��Lt�+�%�^g�<�A`�]ӌ��R�f��#�k�<��"z[>�:��D�,5��{F"[�<Q��02�Y��L�ҽ��͏x�<��i�	_֌�#!�]oިy���{�<�aN�A�ЋUnk�u�r`t�<��HꌙH1�C	0�leP4�k�<�"���8Y$��Nȇ@��*��a�<�Q���☬J�@7qO\�G^A�<��n1t�)���%%F�Xb��^P�<�7�O6�	
q��"gx�U���L�<��g�<�MI�'�[`�%��
a�<i��,Lk���䧛^����Ј�i�<���1uX1���:Ι�dkk�<Q�@/����R�=oX����TY�<�� r�:�qT'���#dTV�<��E�h�-���'�@xP�M[�<iҠF
��� ZY}��TJ�<a�!H�S�r]�g���9?�8Wb�~�<a�ɂg�J�F�i�i{f%Uc�<�M�
��h����I� 	��I^�<�E��Cj$Xq�@� �>��E�1D�{�%��7��3��.� �ġ.D��ӵ�ģB}"�9�@�:�pԊ/D�4��bק]|"�i%+E�vƴQP(!D�8*r��U�젋���3*t�Z��!D�X8v/G2$ HT�H<iX��3�<D�,� �(`��D�K&r�|}� 7D�D
���I�vU�&fgN�p��i0D��{��͝L�$�(dIK=�ư3��;D���T�N�"�uo��r���u�8D��u��#,�z�0h�4Q1z}jv�:D�`�1?A��r��ͼiမ�' ?D�db��1�^D:�$��E�peSv�<D�
ѯ�,�P��H	�\��a�'D���Tʕ� �^)!��ƿX�<i[�I0D�� �8�� S�I�؝ �m�U|��"O����&�%B����I�r;�a1�"O4�#o��#��ɁS+B�z?��[�"O�D�dϓ�nt���U 4,J5��"O8I�pi	uG���τ(-�(u2�"O��FM��4��%Z��Ĥp�"O��wA�sz�As��S�]����"O�ԩp@ͥ(����ڨV`҈҅"Ou%���C��)aU�Q[�ɋ`"O �*��tnDM��[�5��DCc"OΜ�v� %c�����K�9�$1�"Oƈ{ �ꨬ�	��K���"O�4;��Q�h�����7�|-�u"O�A:����H�p,�wHpI4"On}�X�S��x:d� epѹ�"OhH�4&�$��h�%ꛀc��5�"O�U��c���ƉBi�hd1W"O�@S����G���)4@.L)�"OF�Z�,Z	�ā�ۡ6V��"O2p�@̗�}�,���b�<X�ڠ"Ox��D��)�@��`�T(l�T"O�`pv��.�`��&� z�"OV��"�]{b.�H���"��AQ6"ON��U��.au6M��+�8l�2�C"Ot�p�2�����@�8~	H5Z�"O"!p��$~"ʔ;E�צ&��3�"O�5ȑ�F�Y�$5�U�M��haa�"O\�R�f��4Hq�pCZ�u�*	R�"O Ló,��K�u��=)���"Ol����!8L��3a�� �����"O�m�&h�H�8Z��ۖ��@"O����D	(
�@��.^r`�P�"O��� �I/��<b�-�^`\ �w�'��ċ���B�(�DI[��]��ؓ*`L̇ƓQZ���ԩ�1Uں5Sr��Z7��E}��M��C���@q�6�Ѷ܆y����0/N�!�DٸF����8�p���>
��D.IP,�s��/��)�'96�J��Σmrpx���S��ȓ aL+;6��=�D*[� ��'n�];��մ4)Ht��;���Ǐ_'��a1&
 Z���F�'�I �o�D�Va��AtL	ЕCح9x�X�'ۆ���#tY�4Έ�F0����$��!���$����O
u��Q�fQ��p�Ğ�`>Pb�'d��s��sL�%�Y(��'��`�_�/��P�O?u�ሐ �l�`�>[/b�*Rb*D�@{�N�/֝�aF�9�j���=?)��B�|
�#k>O ,J�� ^ܒ-i�-��8���'p̹��P�mW��3!�w5d\��������E�!:V0aG�'��i���)�B�k��۰���q����:!�N5iE�_	~�te3V�P�T��@F:���}���y��`y��P���u�-�\�Sq@�<B� ��^5*���.U�����R蘢~b�ꃣ,b0Jef\>sB�9�@iKD�<i6�
VJn��� Vx��ڗ#��cY��Q�fӢ| ��Ͻ\�z�H?㟸��`�!S�0��J�7��R��2�O�QbQKA�hNh����3n�6�J�I'"r�\�6  ����6i�|��C�ռlj� �%���1c*���0=�Q�N�K���	E����b+֞P_��GIq+�T�i&D�<;�J=w��M��F�@(t�Qdf+�7B/`�1�&
2!�Q?��MJ�3
\ʣ�G�Y���"D���q�ØJ�؍RC���}��Q!*�[*���>���z����Z 5bi)��
,=s88�ڗ5!�$�m�f	!�i�Qpa8��Z,6%�F�4���
ݴń��p�%O�C+G8O��� D�� Y3�X	��'^Zbt�F�`�lZ�}*T�ˡ�VZՋ�5M�z�2� ݦC��
� *Mk'H��T�1ҪD�&w�)����$q�5��R�w����a�� �N$>I�c��D|U�!aUM��@y��?D� �D	2B��gjT$ �8hq�FN��1�/P�}�R�� �5b�|b�O��q效~�K�)�6<�ʢ"O�"�u�E��	�>aG$T��,Ϡs�4Ia ǘ5y�|�C��C6?�뮜r�';2U��'�-��c�P��)�CIdd���O�p��� �v�P�vl̈́>N�`����[L�H��@Ux�Pa"i����8��2#�/�2��,a�ᗠj��8�Bf̓>��:��Є#td[�HY.1���J���"O�Y�vD�*����OW*^�f� V�n@PP�`��+�`���*fc�QE��w$tQ{��<��yS�o�W>����'Ӑ1�@��ג���C2J@1X��������ѭ�Ȗ><�Dᔁ��`	,ғ&y�[�+I(~6�#�BG��}��1p)d�{`P�"���B�?l���_,u/�u����k4��F�[�a}�chVq�0��W��pJ��C��'kzl��"�~�ܸҒ��)J�b}�䦇G���
�:а�%Y�S��D�5�ǎ�y���9Hj�OW��IR���:�@��D �;��@ �J�&@�3��4�'�y��[�|�'�D�@X�Y%'Η�y���B�����+��=���U�b��(
�d�S�;�Fi�'C��#=��X�H��53B�V�t���#v��r���iWH�;g�H1�r�Y�d�ҹs͋dx��G�0s���2�m\�22ش�	�l�6�HW�+af���Z.?��L�?�ŧ�Jߐu��N�+P�8��?�p�'��`c�ޛ��[0Ŏ�m#�)��=�(l2㊐�r�x!3a�Q�<���C��1� a��0L��#�鈟�䈂~Lb��Wm��o�x�x@�_CJ!�d���1cP�A����d��.>�A_2r�� �/O��ٲ�ϨOZ���iZ,e?�����iT��q�'o6A�v ��R��u��qU�SGF����i�(w��xi᪀�)Ċ�����	�٫���)	���A���,�O���BCY����.UbQ�K|*��*��j`�B�"D4�h�WF�<A�`,*����e�IQ�@ k�VB��b(L�\�	��e���8D��'�Ȍ#`�92j�ua1fR�C
ظ�'\R�z�j_�]]�����
b�eE�&��=�Q7{2٫�*A��F}B��"\j}�bBV�nD������V�jL�׉E���W�bd�W��AҜp��5\rpď��,�iGMT��y@�� E���=���)v'��# ��oV,  ��57\�J7��{��=hn���.�v(����� ؓ�&�ܼk6 �58�lP��R�O� �A[y�7H�4�C�'�Ȱ �H�1�Dģ1j�蒄C��A�U�<
3�����YѮɸ�?�p�"2�Hг!:���k�
��Q� 2�iQ�l�`����K ��q��"���0<AD+G4jU&(��N[-����#�Y�⃃�|����ģ�(T�����7�&B����\��>q���>QE;�&� �KԽ@���X�ˬX/�]�>���P�_�FےȒ��ȟ⩛'���\�K�G�#'XyC7�i�έ���d��O?7�H�E�x�Y���(}�0牜#V�4
T)�]yb� �"~�h�}&�	�
�~p�����e�
����>�����v �� O�z�e�%��E�&	�8Ѽ�#��=R~�1R�ئh���^�����R+̐l=|�9�R�
)R5���bD���Ó]�N8���`3�O:q!�Έ#�|-"`'X)r!�2C�	���1�gE�P��2�@T��!��y��� �q(l�ؐ�>��π'�^ĨсϦ�ȟfӅ�ՙA���0��  ��v�i��c��x��Ot%zU&Я�8H%>7-��q��d����^:�Cd�Y�Fo�9n/}��J2Z���p��Qf����&\8Q���WLr9��*��o������0`'ђZ��݅�ɡ4��`p+�LZ9���� ��pQ@!��$0��@�W���� ��"4��Á���@�	TO1s���s��Df���!�P7B����@��[�lТC�QA��!����rblU,Z1f�	�Ȉ��(���"�Xʅ8oaV=�&G	�i|��i��ĪB��,�QhAƏ����ͮL,��B�Q�ltԘ ��*��O %�sï�n����N䈰�:\Odm�`���6:��VɁ�fԋ�Kգx\��0�o5D� 3
���z��'�Hx
pM:|�4�Vj�0���z�{Z/f2aq5�
J��G�P�C�@�&>E���!{����/پ��$�'L D�h�mW�}���4g��bR���i�b����A�^EXy*�-&��|r�O��g��
��$-��#"O�X�si�2~����9ag���N�=��0ۧ�Ўr���S�&J<{��\D~rʆ��J�B4��
\�y�#n�4۰=Q�K�Mz�y�F��L*� ұ����o�t�c�K�3d[�p�T�ݚ[�����)�l�:��K�DH�B��]�d�㟰[���8P0��UH�x�:�RM~
e쎈7��4w�XЮ$4�@���B5k�#�)�0Y�6Έ�X-h��O�i�-�︧�O��T��P�j��|�pm�`$�}��'����Т5B�����'d�(�k�'̤!UXP0����RG:�I�'d��uL#`7l4ѣ�؞SC�l��'��+�΀�K�)��	H���'�"x����;L\>l���;\\<���'^��R�U�$�RI_5/���#�'��ǆ�U�DHR��Q:2����
�'Q����fA�}˾��C�, q�	�'&�d�ĥ�%�:H��e�<!�����'+p	�����~M�A-M�$A����'C
�k4ö>�V���L��0���'! L�2F��R��W,�{�ys�'S�y"N"TX0H7��e�l�!�'�&�ʱF] Xe*��Q�O�[�v�p�'���ϐ7V Xآ��FR" �2�'Ԍ�����bQ�����	�'`�0P�K@]<��ZQ��:?�����'�ݐ�*S�*iJ�����z��Pj�'K�yJ�/J�D���Q'��?u[��b�'Ҡ0!D���H�ڹ���LbY�c�'�L�"ԤJ18��z�W#ݱ�'�T�L�.9����C͒L+,��'%�ieI�.#�2�X�'�9 ��	�'�T��S�娓][g�$��'=�R'�ؒS�^�;��J&]��'�F�g�""@���Y&Ca���'�Jd9�'^*"����
�8�����'��qD,Ќ_��E��
�*gڑ��'���ۤG�����U r���*�'�֤r��ڷt�Fȸc���P3���'�8����4WΜ\���EC����'� D��	�-m�I"�W�m���S�'���8��K�VZF��"�[�ZX�;�'��Qx�h�j��䘕0�p�
�'F��)�S1P᫰�M8%N�9
�'�, �ЏX+RQ��g߰B��P�''�̹c��	f��I��$ɻC�`@�'|���BZ�]V
19�l�?6H�x�'���3��v�b��[�9���r�'�R�r�i:PX�={����=lP��'�fтt��v���J�"}H
���'�69b`H��͘���zKx}Y�'I]c "dOt�HQ*�~Z=�
�'0�����9*���`&�ijp
�'B�$��Ax2�M� �
�|.�L�	�'�>�@���H��"�O�6` 
�'M��;p��G� 	J���
h�%�	�'�z�q�fH?0)��;0�Z7E����'=��%!K-4��MӧaH� �@ ��'=����o�R'�D���@�
$ S�'���c��\;�(�À��
��'϶<Z�eH�^�ܠ�So^/z�J���@��491�su��ϓ�;o�U	T�P:s�U@����s`-A]�S�v@�6��'"��ӈA耠��=<4����� mw����y��Oa����3`ٰ�nB2цЫ5BQ�M�OF�H��'"�~j/O�S��4I��ғx㘸�P*T,�t`qٴ���şd�����m様O�2�SAI]2"[2�K�D�JLF���O�`��	 ���JA�O��L��EX2U�PB�������^��$��%n�y)OQ?u�"��r�=R�"R�HH�E%7�?0g��u)����O%�̪�π fi�D�-�0��bʂ 0@sVjֶN5�� �')�(0"C���|zF:��	��Zo*!br��s�L�A��*�I#ޜpG�M�O ��4�L�	���,�)�f%��x�ر�S�`��h�w?i��ZL>��3�7~3�ɡ��s��IP�Lpӄ7��L?�r�x���O���0�/
�q-�8�ЈY�W��#�OXxy��)�'a�"J�!ѶI�\��ӥClZ$�iGx���B�E��Y��ɟC@\p)��l, Q��)�2�;6�O~�4��(Za�n�A��I��0|j�$�p���
�C�u#��t*�p�2���֝'��"��A��Əb���i�<�0�(�Z�S4��<E��kZ�4N>�[��C����.9v!�Op�-��%��b��D��K)4��9����ŋ �,Pܲ	k�4;��\��b�8xf9���ax���IУc��Tǚ*%�:��F���Y926
<At��Z���h���e�Ǫ����W���04�E6T4�#Ь��^	��s�*��C"\d�Pe��0|1 � P�z�yc
Ca��.Kԉ�b@�{�и�1��!0mv�%����T>AI���!��U�Cj?>Q�,]�n��=Y��O��DB�B;#��X1��H�JLX���%$(�ᓢAZ���R�ْr������FB��4x�D
~Φ����Íp4�C��"MIĠdN�N�p9���%DC䉩��1��1w��u�� 0u\C��;��|�Qf��&�MI0P%FZC�ɗD�<y���3i��IP��όJ:C��=e��<�wH��~���	��M�{��B�ɛt��L*��\�7&dE�6c˗$
�B�	4(4x��P�$=6��I<{bB�I�Rդ��7$ѻ.�(�	�C�B�I=����
M�/��̸����ij�B䉚$�"a*�j�'�(� ��[�"�bB�I�D�F@Z���{e�����1�C��>���n��F0�b�T
"��C䉃Sю���cH��1a��S�P�~C�j��a��H��1���P�NbzC�ɳ,��!T+M>{	�R��V�C�I�Zp�M;v�N~�ޥ2�Q�<�:B�ɹ*�B�_�oc܅Q��͉F�dB�I6;h,h�dƯ����P�4�C�	41��I�����\�v��C��C�>=���$�8*�{e�L�F9�C�"��3!�Q�$��M
�#SbB䉽G�^�;��T�Z��J`���L��C�I�Zf&�0&�l�ɱ�  7��C�D�YSą�;G�N�C=D�<�!
�'}Xԉ��gw�xkT�T�:�P�[�'�<�9q	�:L8 ��1�T���'z�KBkF�"FYp�	U0��a�'8N����_MU.���$rE�\�'N~�I�*��.�Ęb�ˡl>���'�r�d�-7�002A��g�`	��'�J=9&�����	��Js(b�8�'���iW�^����B�P�},�c�'�4����[�N�tMq�h��z���'E�l(v(�Q^�@{�)� Il�ea�'Q|%p���$S28�KȽD.�@��'��=��,c� ���.={�%J�'�|Z�B�pۦ-;e�.x��C�ɼQ\n8�S�]��B�9�C䉧P��M�2+�R ��r���2F�NC䉭B�\Ej�ό��ٰ�E��yC�	>��� �E6�D3c�͝R�C�ɼ;��y
4%�Fs�)���A�Hh�B�It�4*�OË���c�>s��B�Ɏ=�M{�BÇU�@q�'�q�B�I�i��9�@�R��ŉ'��ޡ�� ����,� +RE�j�c"Ox�l�2B�hz�*�@v8��"O��p�ЮLM�)jՏ��� ���"O����n	l"�r�T#|
���"O
,�(�����R��]	�"O��4�X�s�f4�"�J����"O�9+��ɑW-(��*�Q"ODlض�ғD6$U��ΩY��a�"Ol�`F	�7���1i��.W�P�"Op�b���gXТ`�$)L<d�"OV�@F���7s�t��a��j�Dm�$"O�h�s�F�^Q�b�>�hs"O����Q<����o��G�^���"O�6✃($� )���Bf��"O���j�g��Ps�+к&n��[r"OLT��*M�UB�1rʘ	�Ƅ�#"O�m&m�2��0µc@�\�5��"O�t��)F��<����r*�I�"O��Sa�Ŀo��0bܭ96|劣"OR()g�(ux���rb�(�*���"Ovݣ֯�3;��Ca�8l�\�"Ob�{�M��W�lM���Hc��M p"O����lW$�Mބ$��5�3D�L:��	��}c���u~E�.D�D3�G�J��I��ǉ�S�PQڤD D�xQtC� /H�h�S�҈'jTjC?D�x�I��,ˤ��UR�+��1ɷ-8D�l@Dk.<�J�$	QP�h1%�+D�d�Т��t4�fM�gW!č*D�d3�m�(`l<��F"��]s�)D��I f��IQx݈5I�#-l-��l%D�EA�
,v�z4'C�F:5W�5D�lq�Cզ7��pR�@
v8�IS!�4D�<�M�Z�^(j���5�����b2D���-C��:,��]�~8n+D����,X�r�T�C� ��z`�w�(D��k!FMs�flQ��#���%D��8!��,*FE#��+X�!	�=D��k lG�u|v-Y�D0 ��D1��&D���lJL��Fb. ���P�&D��ѩ��?t����݀ ���)��$D�\��!�(y�)���T�!D�C�'�POB ;6&�0 � �f%!D��Q�*K�|�`��lܳg徔Is�1D��+���=M���)��`�L�R�.D����%���`�Kb�t	 �k1D��A�O(D�a�c��g�Pq2�1D��Ô��9I����EǺ	��y"$*D�����8c��(ȗ�&Y�!��.<D�`3A��2ت`�FJ� �� QA�5D�|���Ͱ_��á26#�1D��9a"C�T�kP�S=@u�a�V(*D�\y����X\�Wģ[l>-�s����y�� �N�P4���DbЩ��_�yb��?_���*F&r1<آc�V��y���6?8��FH,X� �j"!U7�y�I
4�h�Z3�-H���a¡���y�⃡:P��qmCC�@)5���y�
�?';���nپ6���AW,�9�yR���+j�	�c��E�M��i +�yR��Aκ�JG�8A0������y2�W�'�<8C�b�&~u������yb!�Ԍ�PW��%8�t '��yҩW8�$%�r�J?�X(��@�y
� ��W˄:���V�Q|��`H5"O�T���G�6fE�5#O�sx�ey%"O��ۄ%�%c���p���\lD"O]��K?5QP�Q Z17R�@"Ovl��mα(��l ��>_50���"O����ɽ[�F��B�G6 �J"O�)�$��'uipA2T��9bX�b"O<|���F���1ˉ
g8�r�"O� �Qo��$ �]z��qY �p"O���c��iS���􂞑q��8"OTP!� �"W��ʅ�MuҲqq�"O6� ��A	=�j�� 7�X��"O����@�t��9��^)m&hAP"O&�I�SY�$���2��h��"Ou�
-��ܚ��p�l�"OD��3��+��@h��nR�"O\ i3��Q��mb��#8VDk�"Oإ�׃t��г@�d+�XT"OԌjB�@U`P�Y��GE��"O�13�ь}����A����7"O�l�u�Y��K�T,D��TD#D�`�e\36\�$���KQ�Eac "D�$��dƠ�ҐK'��au��b<D�8��$\5��%ptn�<�Ҍ��6D��C�H!5�NP��Ʈ[���q�4D���J;>�Z�p��I9s7D�1��1D�<�3�L�u�x,��"�:Q�\��!D�(s�N�x[���B9�D�u�?D�X�7eÖ@���4IA�p7�Qà�<D�Hr�D�1hd�Y!�B�k*Q�ӈ:D�`���%�
9����8خ��Sd:D�(�v�S�<?�hf��"<|A���9D��QdЎ=����m�9nj.��E�!�\�L�Y�4C6`��ۦ"��8�!�DN&^\(��&�[>
w���6��1H�!�$ĕo�@ �ٳv�x�(�D��Wp!��?-� ��4�ҩs�2�`WI�+7[!�DȬ�����%R�-͆E�"��/e!�9S����AOQ*?��ŋC�Pg!��͊ج���*�V���Ia�!�nF�%��'0����'M�̬��k� �ёsdh�9�+.z��ȓS_�\�d"U"����C���ȓ+�*yb����e� 5bj����{��z0�F
�j�6��n���ȓ
��2%`*��B��'�(��ȓ7��0��`��i�	���m,R���E��	�oE���x�Fv�蜅ȓ&uB�nШT���7/�s���F�\:��H�K�1���~~n���BgN�V�������&JdT��V@�S�<�t��K��t��!L K�L�;ĉ�P�<i)
�Y�%�����x�V�<yU��	+�z�J
 ;(��;f�N�<I�f��{B� �ɤ;� �� ��F�<YР?[dUA�Idr�ɲ�w�<���Q�Jl�CCb��չ@��s�<!��W�sD����N>H�JD��k�<��@�=�DHAFE&J	
��d�<�pM���~}p�(F �Y�@V_�<Q"_>mJ��Рe��u4>��Đ`�<Y�,��M���"u�A>�>drw��g�<�b�):h��펍�R�ɌY�<1'kZ�'CR�@�dQ�1�V�ė`�<� QRW*ѧ"W�T��C?z�R"OT�� �HR���憓���r�"O�)��/v`(��U.p��(��"O�ueg��;�ȡ�'�28ꝑw"OJ�[�o�>�18R���<��"O)�ak^"�2DYt/Ŵ_�����"Ot8��iQ�WM`s�MB+4ٔ|�p"OH�ð
͓S�^$hg� Ҁq��"Or�b��5;W�ݛԣ@-A^��ʔ"O���ƢBlG@%#&�ԀnD���"O��t#_�PH�����Q5�x�T"O�!ڧ,I�z~x��a+ңZ�z8`�"O�(���ST��!�lÆy}$]��"O�Ѩ bפ=Ԗ��l�4RWX��6"O�$�#	�r���U��-����e"On�R�� N�IZ�,��/7ָ�"Oz���٥/�� �+�]f0��"O@I����<}۱I�e( 0�"O�4+r�]�-��8� �ñ�Y7"O��P��R�=���z�~�d���"O�T�q*�a�&pS�A;͢\,�!���94isV��4C8�!��/! �  ��       m  �  �+  �7  �A  �J  �S  &^  _i  q  rw  �}  5�  y�  ��  ��  C�  ��  ȩ  �  O�  ��  ��  �  [�  ��  ��  �  a�  ��  ��  �  7	 � Y � �% �*  Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�� |d��"O
`�(�;���8���-0��1%"Oj4��ND^[��"3/9�0|H�"OB���H��*�ʞRy=a"O�味V�!X��!&F�:J�$���"O,��a
���C�Ą�M�"O,$3%o�-���p���+Ն�:1"O��ݢ1����`���y14]2��i�<�6��{_���c�H�`�fX�$Kn�<��A̼VI�xR[�)�Ć�pඤ�ȓA5��('nߡ4�� �)˩%� ���,��r�؊b#`T�eT09���ȓ!�b��g��}�8�F��-? �ȓ
K|m�ș�VṔ���2�%�ȓ"R�X�j�4JN�1�˘X�i����̹	_�jZ��1!g��zܶ��ȓgil,*�J�
j�Ne��i�J%b���f	�(U��:���G��$Y^م�~r�� S�%T"���k\�jx�ȓ|4�1�îJb��@ӵ�ݩn�V��/[`�"�v4�R�!ʎ<��M�ȓ`:��z�ؚh�J�Z��$HY:	��H��p�m�C1��!��B:��0��EnjZA V;9����J[
2���	��4'J�EA�IVW&��~�(aZ��ӹ�>� o�Y�|�ȓ�f�A�
Ο7�H��M�$�����mޠP����/���ANXo*�ȓTv�����{ ��-7�*h��I��sB�8�8���3����ȓNe*M�悡;������X�o��!�ȓ'lj�#F�m�+R&;�|��2)n�C��0S4���T:
b�D}���%���ƨ]�?�Li$ �B�%����
�	r~��*gJՈ\��B�	�2Fl��J�4m�x�����\�RB�	#a��u�bY�U�����*\jF.ʓM�}2�ۿ:�h���4��<�A����>��O8̚@�K�X�>�"��P���=���Is���B�53�]�'a��,_�����[;Wt��F���J����#(Ա+���(V��y�}�h&�~t8We-�(O\ń�Iz@}�BB͈$Z��N� }y�I_��,qm�8B��q	_�w| ������x"�	��4doե?������y�A�s�T��털�P��㉔�(OԢ=�O����e�9
H"�m��~۶E2�'�|����� �T|&ǘ�tl�����)��<�e,�Q�xIPDH.<�T����H�<��$'����Q Uk��r�DB�<)e��{�A��1�,����t�<�T�8�9���8n�.mK@'�o�<�3�C�a�����Z9K��� �u�<�"n�8�Z�ˋ�=p����t�<I�5f��5`X���-�b�I�<���O8J��p�A@]�+9����BG�<�pe� 4�ּk�JTq�n؀�@Eh�'�ў�'-����J�'%Z�x���:���	��?ɡ�AF!�����z��0�A�J�<�d'^�'��	��j2A� ���	O�<Y��
[.�A�$1eGR鉵M�I�<�'�	m��It�^������FFH?Q�'>N &��}� ��u�^ q+���ΐ aD��3���F{���v��q�獖����K��ݩT^�����ԟt�)!Bݛؒ� T�*D؂A��'�I�4��+rX��J �G��x�B�g
�ٰ���A	:*qJ�O|d��&�I���I]2STb�9�Ҟ~��hq��Dyb�i�i!%�0v�~q4��1d��p���.�O  I�t��T	kK�d���"fQ~`V�j� D{��)��y���,W�R� ��⇠*b��(˓PyL��4�,b�Pk��V
\m����JP	F,!m����GD�{���&�����'rM�VÄU�B
?=�P�b����O�b�����T���Zf̸�,\�-�h�a]��y�L���%�V�PRF���8�IEy"�|b��.��[���2&�
���>9
�,����酁r�Ċ��џ5��{�ȋ���I�Kӎ��)��gb�r��[{,F ��+\ ����6p=.�:�J��P[0P�ȓ,oR�:%C�dǌh�e��E�l���-U�%�%D�?jjf�H�%�'�B��HoZ#T&�1 ��Ds"k��C�		����P2G��( +�*�O�mI��\6��*40�x� ��?�>�p��1D�4ʱ`����I#c
��5�2@/D�Tqk��rH@�C(~���Kg�+O��=�B�uCT8K�CH�IH�`�OQ�<a�R�3�xA��ā�j�s��M?1�u H㞢}B%6�Z����AI�t�#4!AqX� AU�č�*冀2B㜎�fH�Q��!��ݜ`�6Ph�DȘ����5(�JL����y�V�1#��3,�h �I�O1]�D�'�a~�A5���'ˠA�dhլ���=��yb�)IQx�a-;@'(���@��y���-o��E�"(�6?�y�e�KX�U�ቫ�H�2��(i��x�#�c�L�ӁE<�y"׻G���# -q���(��	���,�O�ZaeA�h'(+֊ &9�\��'��	/;����<�"+�+éQ�:C�	�D�\ꤊM�n����50�r�>!��?N4�SgE���]�V�֥J��C�I�|�-b����8p@�2T#1��$g�D�>E��͝M�t��4� #3h-���S3&�yR�	�1H��F�
.�b�$A�V�w�a}��*LL#��9�
9���+ܰ?Q�1O=�,θNs|���P��<��"OfYI��h��]68D�E��g�'q�xbn�Ju�a��(ҝ,�l��ǚ�y�4/��$p�g�$3�2x�ǥN��y��'�d?�S�ӑ��Ԙt���LhK��ǻ-�"B�	1)S�iB�m��up*d�᠆ O�"�<��pD�b��*]s�`'*$SQ��y'��<E�$W>|��Ү�?^�;��y�ٜ|m�)��[4��p��L�yR!�.?VNpx'�)
R�Y�b��*�p?��Ov� �@P	:C�yb��� 4��"OΜ"�l�[�p53tLɌy%"D�P"O�9{JO�&�P�[�)ҙ*$l<D��H��n���:sP8Oj(��#;D�pі(Ʊ,�Y�NG�>��&�.D����d	>FF������x-ip�O��=E��d��[�8���k�:v�
��F�a}"�>�F�\�;��P�
�#GdҠ���HD�<$�_O�T�
��6X�i�%�~�<�W�Wm��=q�Ú3+LJ`�JMQ�<� \1�J%��hQvk�"\M�] ��ɸ)���DD�ZN�`��rBm�d3gg!�D�1J���)_�<uĩP�"f!�$A(0���� ސ3HԊ��d�!��A�Z�Hi@ш�,q���:�@�<J!�yC��bVƁ	y�ƕâ11Z!�d>	�n���
�I�0��&��<j!�d�P��	��N˸uJ�T��� NqO��=%?�v�S�HZ��롏ˑ�̔р�(D�����K ��	/t���gC%D���n1n�-�t%��m5!��� 8��룍 �����< [!�$��4i1�w��	�0D�b)	�T�!�d̈́4Q��ʴ Q��@5�T�E�,�!�dU�=Ӕ�
�&��X%�''V'�!�D�(9�ܹ�)�;%WF��D��C"!�@'],be*�K�!�|x��BJ!���ϸ�����=�\u�6(�>!��Q��+K.������*�!���N���rs��0����\[�!�|!v	��'6���@�N2)"!��I�#L�����%�dE����+!�d�*:tyQ�@��'40 ����z�!�$�6�����#���2�M�u�!�$�	a58q��:i���E	 8!��Ԟ<�Z8��8���mP!�5j�Zܱ��K���Z!� �f�a|��|��Q
v|D�B �0�	��^	�y2H�.��Q�t��&��y���Q��y����>��A�-��}C��P����y"��R<��8ă^�|���ό��~r�)ڧ_�:��'X>7�0�"�ɳ �ȓ?�x�@p�W�|6�!��T�6ćȓ:Ɗ�	"H'���SΪ,�p�ȓ	#f���� m$�@���/l��ȓg��@tk��.�@��商ir��ȓN��Ec��./���[�ǿvh���ȓC����RHn�*� x,�@���P��G.D�!�ך0��t�ȓs2��!�B	&�2��a�,70�ȓG
��ɚ�x��������l���k�R������:N���(
S���ȓ]B�����8&,(a� ��=jy�ȓI��u�܁M�ԉ��f@��jه�"�D)Y2��)�^IqЇɱ{�����F�@�M��\��+u銱*�~L�ȓ	��*u@X p�q+� �B{�x�ȓ��8!���_��+�^I
�ȓ~u�O�;�����ᔰ�'{DВ�
P�K�x����h2�Q�'Wj<� ��,ZE��:�M0��I�'hZ���i^�["tHQ&~��X	�'ٸ�%�[H����݌~3K�'�V,r2lߖ�6���%�>�R�'m@���5�U��Ȫ5`Rth
�'���rJ�>#O`#�O�7y�U�	�'�,݋���H5H����Y�ʜQ	�'���`5�ΉLk�a��N W-���'��E �l��'B�̂Š�D=`�0�'U��k2�W*:|�ԏՀ;���q�'��4`Bc��\�ፗ��Y��'���t��AaUPs"f�d�I�'���xw��?�� hE

&+]����'?Z�4�CH(��J dR6
.���� �I���9R'��Ie�R�i�ŁU"O\5��3Z��5�E.M��p'"O� ���?u��,
D�(�T���"O@�Q@�P'r|�9U!�
ʺ4:�"O���%T6n�JԢ�ܠgD�;��'Z"�'Y��'z��'��'M��'o�i�d��x��qpt��7u�$81�'R�'���'��'�b�'�"�' ���B�Ȥ@���̿SBh���']��'��'�"�'h��'>R�'!�胒�H6��U
3�P��'��'�"�'�2�'��'lb�'�(��e�9qh��`�D������'q�'?r�'R�'z"�'�b�'��{�kR�.bY���O>C�`[r�'�B�'b�'y��''��'�R�'�����G*G��4AY%)��S��'Q��'	��']��'!R�'��'5NAS�	Z���@��!T56�IQs�'���'"�'P�'���'���'�P1$JRC�N�7@ӫ,�tm{��']��'���'/��'cR�'�"�'S:tJ����J��Ց�Ύ4j�6m1��'WB�'���'"�'���'�B�'Y�4�L�!a��0��F	����'��'���'���'���'"�'�^ͳ��
�D��V��%��rB�'��'��'�R�'�2�'/��'�&��� �=r�Ċ$J�7���u�'��'���'P"�'��abӰ���O��@`)U�FBb��%�6�#��PKy��'��)�3?� �i��Sg m�V�u#ϗk=0[���%��d�צ��?��<Y��i���z����L%G
9L�L�Bn�
�䙳/��6�9?yEH��E2m�C�6�dm���x3��� H�|���H�9��'��X�8F�����I.��U��t�X�J��.�6-ϥl�1O��?��}a3��PՒ\YW��v��\���'�M��iB��>�|�r�ֆ�MӚ'D���2��
k�*ȫ�f�
j�`�'i�-�v��6l쑱�i>����V�z�ㆺ\�Uk� 5	�>�IoyB�|¨rӴ�e�D��m�L���2i0��"�8-6�(9�O�m���Mk�'����.q� sV�8��11H��B���9qx�T���^�NE�|2�솗�u��OB5�i��"᜵������@˓���O?�	/8W�l{Հ��1~܈���"}V��ɺ�M32�LO~��j����3�
h��;yqF��2W��0�M{1�i��Ӟ,����<�2�S�� 0�@Li����ŵm�4l�A��,��a$�t���Ϙ'�^�	b�
O��0���4,�@�O@n.w��x�'k����J>�@pЬ�-% ��zPf;8ʀu�'uj7mG��'�b>U�G��I悄S�ұ2"�b �ȯ4��M�īBjyb���*32k�
ݧ6�x}!G�ѐp��ʁ�A�|�����
+��S�̋if
 z�끈f2 �41���x&'�=��8�"�(Cb��Њ��E1�Tہ�˜4)�$A�,���˔�=dAc�L���'~��A���'JHq��~k
��e%H���0�&Fx=�F�L.N|��@F��JzB�� �ax�� �E������0ju�����A6�Y*�Aϋv�qC&�X�Z�h�l�>>���e5@Az1��+�,�N19�bA�q2�����{ɘXy�ʛ>V�l;��L-�?q��K�0 >!�DG�?Yآи�F�'���'{�'���'94��v�'3 ��/�0r�Ƀb(�$�n��SI�>��?�����T�M_
�'�?�+C#Vt��5�ۗeNti���߆4���'��'h��'�D����D�4c�����'kLl��d
�X��F�'�r]�Pa2��F�4�'��O8�H�Q�hf`�r�F�y� er'B7��O��D�����'m�`�:#��
HH�� P�;�&�nZly�G���'���'�$[��ؒ0! �:g�=F��J���z�7�O��D�2F���b?����0J&(�$��4AW�y�4�R��O`���O ����V˓�?���' 
ʖ�ҬK�:���Ń[h�蔼i���'��S럴���]Z�\`�ᖼ''��xFm��M[���?���6tz�K+O,�d�O��$���S�ˈ�2�1�q.Ȃ=�*�'a=��}ܦ]$�\��۟���/#�hA��Q�%�B�t��q�ҵ�޴�?i�����O����O�Ok,
>�D8tǁ�u��UɇԊ[/�ɹ$���Ihy��'�R�'��	3���r1�V�| �`!�/G܉�GKgyR�'2�'��'"�'�\챶a��EfT�V�_)0�JIa����Z�Q�t�I�(�IGy��Î��)�z�xc"9�$���؜D��'h��'�'i��'�Y���OR)�B�ʣ*�"�(Ơ��Oʈu�[������H��hy�>���d��/�tL��K��px��o���MK���䓽?A��E�A��{"��#/0����ψ��e��(�M����?�)O�T�"e�|����?��'xG:L���@ XR(�!`���nI�� c�xR�'��	]=�O�S�3�!uN�(pL��/U�7��<�����?���?��R*Ok��Zm�({�`I�`B
��eI
=��V�'.��	I��O���L��'�h��t�c�X�d5qQ�iX��;��'.R�'+��O��	ȟ��I#?����`��<J�(�"��1�$Q�4&��娏��i�OT0�#H�&ݫf�>;�`}��aRϦ����,�	'#�*��I<ͧ�?�������s�Ph���w�Q�@2\Ȣ�iZ��'������|j���~
� ��x���Q-.Y���9_S�eb�iC� ǿl�剝���)���n�>I���;
�� �����~�AK<)���J~�'���'�剿�ll�!�w�c���r:R[?�hO���O��D�<y����T�/[O6pz�N�cL�����M�������O���y�'JP��ӟ� ���˴�j� C�&M ,j��ib��'B�OT�d�<�G��������/t�A�5c@%1+؝��f(���O6��?���,���O@�KW
�+uÓ׍�;H�~�Ss��Ϧ�?����d�7p�'��E�d��-A �1�@ �°3�4�?����DПf�rx&>���?�X�y>h��
D�B�2���b��ʓ�?���?������<��r��-
�C�z�� �&��MVl�ty"�6�.6M�@���'��"?AE�>~�8�����'��}������	��I��PBO|Γ��i���Ѣ�~JB�����l/�,aݴ) �����?A���?��'��?���0�t��Lh��"v䖫��D��  �b>���$z�s4�K�t�ҕ��C�(�Rܑߴ�?���?�@��O����'�b̑VeN���O	`4�P�W���7��O��Ħ<�%X?�I͟,�	���9�,ٕw����׸ͮ`Pj܇�M����
�Z��x�OV��'Y�i�ni[�?%���.�����i�����$���I쟸�'�@���������
d@LC�"�;V�O����O���<����ɿUYm0w�i�P(��.���M����d�O$���<��3���O�\I�b!�1@��(Q6`ʩv�.�`�4�?q����'��P�@�@!j��	k�.g�~�+ѫ�Cw* U�x2�'��	㟈�v�I���'�¸hb�;:�}�2���UN���u���t�	Xy�fK��;��i��2H ��*Z&ѐo�����I�@���[|��ڴ�?����?���dZ�!��MޒC��!J���$2YX�KQ�i��W�����o	�Sߟ����ܴ��C�Кk�ج��$G�s�0o��������ڴ�?a��?��'����<�*��3��<�
`�AJ�)V:�ST[�t�I�?x�H�	�䕧�$�~z���*5)�ɜ�*�q#�-��A:�c�M����?���b���?���?)�
64Ru�SM\-cņ�p�&)����{r�|�O{�O��;^J��Qj���k�͔?X7��O����O�|��������8�I\�i�l�]DTӤ,]�S~ӊ���<yA�<�O���'�l�,*�b0�f��>��]8d�n�7��Otă4`I���	ߟP��֟lɯ���7Ej��1t.�cu�iC�_�T�����ϓ��d�O|���OL�?Hp��%F�<h05�Ԧ��R�EZ a�Iey�'S�	埐�	�[�@<qʤq���=[鑇-xh�	Ɵ��	ޟt����d�OULX-k����E%Z�5j��L��VQ8#��Ϧa�	�������IyR�'����O$�d����a��
,�)0BR�x���d�O���O��O}Ys�Bm����O萡䫔�
~�I	��M;S�h��	��	����	dyR�'�f��O�"�O�Qz�@Dt�!JQHEkRn�c�i
2�'(r�'!2��tlw���O����~ຳcK�_,� ��IR��8��Цi�IZy�����|��?�)���.O�T0�ɳ+�4@ٙ�M���?f� *����'���'����O[r��;\R��7#� I%�(R���9p_���?�K���?�����4�z�O�����=3��]S�R:w�A[۴o(���R�i�R�'���O����'��'�> �Wf�����sb�(|��o������Ok�i~�ï~�M~��� }k��կ8&8��HY�-�YH��i���'2Gî��6�O�$�O$�$�O��C�F>�ŋ����c��a
�S�qh���|bA!�yʟ����O����hq�M�����~�	8wd��l���K���MK��?���?�X?���AWM�:6����ê�c�ʱnZƟ��fb}���'2�'���'��E�?i���H�Q�xP
!�p��.]��U�am� ���O����O��OZ����4Ib���$−@^�3��pK��?����?A����^�:7X�o�4IK�CՎːZn�XӠP�.�h4��4�?Q���?���?9/O��d3 ��<�6���\)W<8�9b�_ƤlZƟh�	ɟ���؟`�	?h�f��4�?I��	#89*Q$H������̐Ua�=�Աi��'�BU�`�	�{ƈ�ST�Ą%p�n��Ԥ�<&|�|CE�<���'���'�RE�L�7-�O��$�OB�	��p6�����[�R�)��AM�<lZן��'ȏ���D�|��M��0`I\<���W��x�g������˟�Sl��M����?9�������?�4�
y����� `��j�*e��ߟ��oܟ8��Ey�Op�[cPl�7e�*��Db�9�Ms��U�V�'HR�'r���O4��'�2a�7^ $�ό�8Q��Մ6��7��#� �D�O���|�L~Z��2���K@�h�V��Tό/Lzٰ��i%��'�bdϵ.�7��O^�d�ON���O��������_7B-��O�)���':�	��Z�)2��?y��-C$�;Bw%��@����i����F�6��O�$�OB� U���O<�33���:�0`(��>
(�[��#�k��	�p�	����A��Ǆ�F�(؄.ș_�^���e�f!t�l����OL���O.��O�����֍f�R9�/0��HK�K�")���	Cy��'���'�'�|A+1&j�l4� аj4dגXؐ��܌�1�i{�'���'1BX����4:��Ӡ!P��	 B�|�s�[�_�2U�ڴ�?����?�j\��Y�bdh�4�?����HJơoT�;E�L�`�<p
t�i@��'��S��	$A �Sϟ �|)ڹ�5�\�n���TfR�5�l�������H���Lhݴ�?y��?Y��~�Ҍ�̙�D��`�iZm��T���i�bW�l��0��ܟ�����42}\yC#%ߓW̪�7� s֠�n����	Y�P�ش�?9��?a�'�R��(��%a�ϗ��LiA����X��S�@�	�Cx���ǟ8�IS���~�2���<��Ĳ����Љ�0�Q��]�A�:�M[���?A�����x��'�Ԥ�!BʽS��"��L�e��iږ�y�^"���O��O>���)G����@+7�5�M�B�z��ش�?a��?������O�����i�ߟj&^d)�(NK�(��A`Ӳ�O��sf��@����Iɟ|�Ǧ̙9�/ P��U @:ڴ�?�PIщl]�'f2�'�ɧ5�MI�J� g*=-��=�Y����@�I?�ĩ<����?�M~J%԰7*���c01OV��ӻr��1�F�x�'�2�|�'�H�SB�`8���T�l� ��a���P5�'���埘�I۟�'&��c��o>�Â
U:a�B���I�Q�2��>Q���?�L>Y��?qA����?I�*Y�gl�g�U��U����|��Iן������'���7�;�Y b��y���A��"%��S�،n$���I�$9���៴�O�i�	(a���3�����yy'�i���'��I+����H|�����ā�7�,a`TN�ٺ�R/É'�b�'�p��'"ɧ�)U�L�푑l�2S���ӅT�	��Y�	��)�M{�P?��	�?q��O9
"�J���f�--b�kƹi@R�'�$�K��'��' q�
�zG�%AH���g�4t�uxp�i�����`�t�d�O�$�N$�8�	:2�"���Jq�AS�M'���ش1�ĵ����S�Ob��Ǥ�v4B[�R� �f�P�wM&6��Ob�d�O�X��D쓑?!�'�bM���^��g������4��4>��S���'8�ӟ�b��E�KJr|{vl5�`	��io2�\h7�O��D�ON�OkL"��	r!�%�t�Aj7���&A�B�	Ly"�'���'1�	$ռ����ˤ����?
���+J����?���D��97,�\+�a����EDR̒wOz���$�<���?I��?A��(����i�2� ��|o�$	�I�F����wӌ���O����O��$�<��wwU�'_4x@ᆩC�fjLX�����cG�L@�\��������Iҟt�I�.L�eX�4�?	��j�����4>&�ׂ �/�N�:�i<��'�Z���� w:��Si�.2|�H���y1�3�g֩xL���'�2�'�m��[�b6�O����OP�	��j�.��e�ڠQ��)\�V�ʌo�埨�'���H���Ē|��M3��N�&(�,@nY�鸱*�ۦ���ܟ���\��M[���?�����'�?YT�t���#�O�?h�(���2O�Iޟ�8�Lٟ$�Izy�Od�'Y��H�N(X)F)��F�"E�D�oZ�����4�?Q��?��'�z��?�>6�h�d˙���a㈙w�Uȇ�iK�#�'��R��H��C���5���8D�\��l��	(�Mk���?���KT���i�2�'�b�'HZw>�%�5 ���\ȣΛ�)b���O4ʓ/�������'Bb�'�j�`�2V���kfN��t�2���fa� ��Q�I�<�m�`�I������鬟4�RHʜ+�qE �BIQ/e�7m�OJ�j�>O����O~�D�O���|�tBħ0,�7��=��M`2H̎Xː@��i���'F�'� �'��$�O�H�U ]�5�+K5p�@-���ѬX�D�O����O\���O�˧u<&�0�i�T�֌F�G��0�BX�w�4��v�v���O����O����<Y�S�z���k�M9p�$��A�34�ڬ��R}��'��R����S�<�'�?IS�B�s�fF�y�*���ۉ61�F�'>�'l剉Hɦ0(��+�DҾ7� Q��1I�N�;T!��N��'l2�'����>zmR�'�2�'���g�)a&dܺ��h��`��OB�>�`O���<��	j��ug��19�ޥ���J�7�f��!���M3.O����̦�I������?=��Ok���NI�AɂȞqcޝ"��#�'�"�Ia�D�.}.�׬B"��B��Y�t��䙿G���'���'5�t_�$�OT�\�ԀSv2t����+"��Re�>iV�z���OcT��cN):(�%��I�	+��޼%�Rm!�AA8(#0)��&S��8mzQi�f��z���H�KCG�\_��0��w��~���2H8��J"?��Iؤ ĺY�@����GوtR蚏[>*|;���/��UM,#���%"��M8��H1���k�8ӒJA�o<��U+F�7Wju10��(#�<�ӓ�(2f˚Da~�	gIN$�*\1Q	P�q���TGʇZ�8�rϪ$#����꛱o����BP���d�O���O!�+�O�d}>����ݩ�.4K�&όg�)3���0�t�@�чH0tqۓ=�����͝��% e*Յ"�H�Ù�:������g�a{"�վ�?��HzP�$�ýl"���ؒ"�j1#��D4�`6�pY� 	�ID����`�Ԇ��X���ɑ3U�����P�m>>�Γ'c���'���,v�X5۴�?���� &|�-�-a2&�b��@�C#�Ӂ���?֔�$�O����*d��d)�|2����d�w+вG �����u�'�������r0�,�e�8ƐAd�^6/�Q�xӲ.�OT(F��n_�j���R
ݙJr"�� �y�gƓd�,cc@�~-���3i_/�0>�v�x�nF�x�̺ $�q�x�l]��yB���A"��?�/��@9��O���OʭcfkW��~�94.��aZ���^g�F	��l��hN���I�>�O�1��(K�E�����H2f&F��1���e�ſoD!G
]�#Ͷ�S��?)�E^ M�6\�Ԡ�&a'�X(�bZ�����?��O�O��'m���J������d*��-X�'
6���O��=������E0����B�����'I�`;�V5�Q��N75Lے�'��g��a�F�JP�'@��'i�Nl���	ԟHA2���s��2����P�3����ܪc�X��])V�2�p<Qa��+
yR	�oL�>�4|�b�t?Ia�ޒJH��C�4�x�vq.�7��8}E&<j���~�H>�?���hO��P �c��AY8�kbGG�(�E�ȓ|{&ɑňgA���d��Z�F�2@�i>���uy�i�i��7�^�s����HYba��I�4.�����O���O��@��O��D|>]ɠ�C7�2-z�CK�S��r�Љa���E�^5����a ��yrJP&jZv��g2?~�2�dJ1u6HpʸY��ـg�0)�ynʸ�?I�q�-���<s1����8Vؙ��:�;�x�eb��l
�tc1�:Ad��ȓ	�q7K�	�I���G�y}.�͓|�&�'	�	/h��L�ߴ�?!����	̣���p�-H�"�`xѱꟹ0�h��S��O���O�ժ�Iڧ.�0x0&�2�~�p�t�#$j�f=���L�P�DA���(O��v��]�&a�瑏mx����!@w�դ%G��ˆ��/$��Lps�I�7��D\䦝����ԕOy��*���!��I(v�X�P'Q�7�'���'������I<�~h��N��'�V�{W��0�����D��&w���g )+�8��WP���5f%b��4�?���	�!u�Z���O���Zw���0�!��p��b����(�O2b��g�'\ ���,�� `����������؂��"~�I�@��}�r��.EԮ?�����j�����OB�&���7�\�q#�?d����"O�,��I�;�8� �-���I�HO�)�O��XC%S���(�݌Y�>�r!��OL�$� ���y���O��$�O��ĝ캫�Ӽ�Ĉ2� �3���8�Pl�i�J�ʣ�"!!V�3���_����'R�Q�8�4C�0p��r4ԗx���!�OSxA����Q�~�a�5+Jk�4�ө_�9�p�E�`"�I�-p��p�ӴU�
������!�I�n����؞�wK�l���c�N% &8�c$D�����a�D��G�k]���3)P7�HO�#��ԙ*�@�m���v��q�4���@eo������͟<�	ɟ��N͟����|z��Ān�,T 2�=L�D����t[^�r&�I/'���ߓDBdsiI=nKF(YNʪ��$3�@�G��AK�\��<[0σ)*o������O,�n��I���,Ԯ^�C�Ԅ{�hB�I�s,~y[d���&Y�V鑊fB䉀Q��Yp��S����G��X�I"�MK>�dܞEu���'RU>��V*�gI�estlM	�b�ZըB �8�������+v��`	�&t:�YR�A�!��+�ޟ^4Z`�U�C��9b& 9F�C�剡3B�4"�	�z�t�[uX V�����E�1���s�$�3 e3��ҥ�P��t�H M+v�&���t!�O>�F���ąp*��t�88��l�6�C�y���D�Cr�ݗ7]�]�Fl����1��|U�xeI�D�-P���ZH��%���y�G H��?a+�M����O��$�O�$#�×�{�h�)�M�F�:����^�ͻ��m�J�7h�0Sc\��O�1�EQ�(��`�2,تF�f�5{Q�1�!��9�R	CW(ƉV��Ԣ$�܇�$��1,�7r�v��߹�`�qo0ь�9hv����]���0�I���D���C���XA
�DDv,@�@Q*/'�b���Iix�<����Z��uP��;r���#�^l��H��ßH�d�A;��@э�ZEvm��' ܟ��	>4Ol���������I㟠��5�u�'%L9�hA��I� b����~2�W�.OܤXP��l�� �U5*��)��㎞}�&��  d*�Ś i�;,W,Pئo�<g��3ړQK��CW��
,�����#U���P�Y�Vp�I,��=I�O8I`�2��\;6X�$"!���h＜�PKX/{�`�hY5��tFz�O_�'��2�j|�f�v`�u�=8p�be��@�E�Ox��O���;jVr���O���U	$��$Wb� ���&��\ҵ���V$�T�h��Bw��X��͉1�n8Ju�%CV,;�a��[=�!����&�j���#sJb�������ơG>w�@A*�&'T�V{$D��1�	R�k,�"C�'$��p��*!Oޣ=9U�]8n��U*��Vh�٨q���<y$�i��'�!0�hn�d���O��'A���cH������gM5o���!D�?a���?у��&�?Y�y*�hU�� x�5	PS}0ӑ�ɢ*U��z�(Xj1@B9Md�T�PI�'� �X��LY�>�!��:n�9SK�8î�RVH&D���G�ދx��$�F ��i�FB�&�O:�$��"&��BR�3���9%���#��c��P�K���Mc���?�/����3��O���OeY���R�n�R��S,B��H��28��6�|Fx�҇J�6����9���IbS�p����7�)��(���8�7��'75VDH䊛b�`a��B�S��?�ү[?$���c!��8��'�u�<�ӭ�&I%>l2Go�	��Ʉ��p�'fn"=�O��}��%�<BKĭ��'G<�l(��'BH�:E�����'���'��w�M�i�Q��	j�zX9g�
�&0��i�B��L:E&�O"�Y��R0��3����XBu�O�(�"�'_δ�1E�22\^ܒ�c�'H0�X�'�����B�a{B�A�k�>����R>����CO�2�yr���o��l����3y���u&�.nh�"=E����#q�
6M�n+xat�]<`G���Ӥ�b�&�$�O��D�O�%��O���u>����O2�d���@5�矛.) ��C��6��|����$:[��`;�%�h�9��u��|rdH��?���i��ѻ����U����/=r.�C�'��aI�M�/��j�b��-��<{�'hjP�M^��BP���\:%�0�'#b�zt�M�Mk��?�*�6lq&���z ^KÎ�%I�)���'I_���O��d_�l&��� �|r��Зl����D�eͤW �\�<i�L�R�O��E3�DC,).��R@ ���0y���&~�ri#�'Rd8UHQ�/z5�B�ǿ;���ȓU�����Z~�����i_:Z�����"��L=����	3x�zb[Lu��ΓC,��9�iD��'��b`\�����I���x��ܾR�i��	 P����W�Uv��>}0��|ҏ��g�����7�
<jƃ(8�s��F�l�Э�0VRZ�S��?�E*T�`�h1��T�$҉pf�X�J�*��������L�Q{ ��7`�*]*�%�pF��yb	(gU��a���V4#g���OR�Gzʟ8���Xp��u�aV"D����O���'85��n�O,���O��D�C�Ӽ�A��H��J�.�3ے�w)�T?Qb�[3v1��E�'���7%�7	@<5�R�ŖLwT�ঔ|:�Ukpœ8���`W�Y���d���' ��#�[s�lP�ɘ�n��Z�'��������=	T�iD�)wfS����W�<!��L&X�D(��<#�̠�O�=瑞"|��×�B��kA�X�b����	k0�"e-[��"�'yb�'�rtP��'��1��1�֫J��T����<r��a�鏼bfDĹD� ��FYJד8��H���b���ۖ(>S��Ka#[o4�rS
��[����$[��lv��uplZ�dq��+��$���c�U����?���s��B#V!y�n�Q���l���Q�M8D�����L�mё�r<��t���O.ʓg�T�0d�iPB�'���C6�(��ނ7�ޡ��a]�2{��r��˟�	ҟAA�ҟ��<�O�I�{<���_�i>,�K��$J�Rl�?�p�K��DpJ�+ ��U0t!%ʓ@R���{�O*��G��6�x(���T;_A��S�'c�Y�և�tt��/[7_= �&�'����ϥ��3��S7RÚթ�'\��a�`�&�d�O��'D�N�����?q��h
f���$g��Mj�F��5��ք˪�?y�y*����+ċl��p@R�U�^���l�>Қ,Ex���'��ѐ� ^�R��C��")� ��J)�+���O
%�M޾Aw&���X�T�$q) "Ox���Fb�X�2`Q��!*q�I��HO��&b���oII�2��_,n�b)�	����� "!p���	������:\w��w?.T�O�-"�	+��[�Ѳ�Fί�pD�"CаuQ⨁�G6�����#�X�<� ���M�p�̑)��b��ɢ š*h<���^B>�!��7<`�I�#O�ȬۋyB(�v��$sE��#B���ۥ��~��+�?y �'0����&pD��fRO=�x�	�'�0(�lȻ/���`��1@�v��@4�S�O��qr$�kӌu��ǃ�;I��r"ӡ)˔e 1�O��D�O���+>~����O���2�=�A�O&1�&��Rm�ɹ&a��!\&�S��'FXȠ7�(�?���*h�c���I�$��Zq8�,���O\�� �9)͉!���#�H
�&"�$�O���?y�ʟ��(����
* $�|�(�U"O�M�'��
2����@�"^���
W5O�Q��'��	�+��^wh��'u�Ӥ *�e����6[�&�j@�ݓA-��"dǞ��@���|!&���L�<�O� �'c��:M�w��s����R$Xe�?��UI�7k��Id@X�fJlP�$/ʓJ��I��H�V�����B�j5��*��Q�$�*6"OU�H�t��{���*�lA��'ۨOp�1�R� �jS�Z��xh�;ON,�#Q�Q�	˟��O�<����'r��'�F�P#H�=���bk92At�
ޔ�,p����
٘���'�9O�C���F�N\�C��m?n����c�kh]�+>6X����XCCh�|G���#l/�(BB
s��(��R�5¦�'xZ6�N֦Q�Ix��?�慄Z��,���R�Ls*p�A*^�<i���>�/��X�`#�0lw6��	�i̓�?!P�i��7M6�	'����O)|�ƀh�\�6 s��[�DF�'�����q��'���'�4���p�	�br�}pU�F�[������l���	;WLm��'8�	��CTfb�a��o��i��'�p��e�_�h(E��N�p�yr�́6P�IW塟p2���O2�D,���O>�D�<��n����3��d�xi���x�<A��.R�>dSE�'��}P5�C�{�����D\�K��o�������5'���3�
B��XE���������t�.Tǟ��I�|
ԭg�����4�����h�*,�4�?�Hp��	�>���"�͉�����j�����ˑ�4�:j2�O�d���'�n7-޳DʝI3.�) �D!"I
9joZ��|�'����?��IX�$���eI�5vaX):�=D��Q��$j�@!በs|���e}����O ʓ.�f�k#�iQ��'�����]2AW�#�Z�I���WY���-��@�	iW#)*ܒ�C^���q�S�� �W ^�X�g�����S�����(O�I3���GO�|�A�(���Q�
�|i0x�#E=2�����	L=���IϦ��4�?�*�~mr�j�B��Q�BU-$�UQ��O��"~�@+��*F��MlpL�b��/G��Ą�ɫ�ē		`�# m�l�R�jׁM8<t�:`��f햼�?a�������O��d�Ol4
Q��?6�}{�D�$ ���kfτ�&
benZp�S������}	�%وkԒ���.+FF�U��iM�S��?9�K��N�J� ��1�X���@����B��?��O����O���ƙH.b=�'��?a�\9�0O��d4�O>��.Ǆd���2Dȯ` $z���?�HO��@����C��2I�vl����=u�	�Ы�E9j�L����,�	��d�Xw���'󴁭�x�Ь���� |�Հ��:F�!�O:1jB�6�6��aO�U������O8%���'#je�S�E�%�J�a�T���'Lh�h�a{O��u�<d��Ph0�Ð�y�JA6PO	�%i�C"xx�`eU�#=E��'�XZ���t���	TDQ�
�'�.Ԋ��ߊ�5��L�'�B��
�'�`�2iԮ)�B��P%��&� ��'�����cN�\����F��%
��r�'&N�ps�L�Xu&�"�i�,C�\��'-��:��]�?C�S2�.[V� ��' �0��$�Pxh��"HO?E�̅��'�֤f�F�/� X��+=(F"��'/NLxf�]a��ĉbn���4��'9����W;w(`�����o<���'�F����LD�"��B�?�xa�'���%��B��@��ፁ���	�',��BV K�Em�HcS�IB�	�'n`14�	 AO�!C�B"H���q��� 0(��+������e�5q �*F"O�%@UJ��23���*Qdx��D"O&mpOӫ)fE	� �6I[���"On�8��1?J�"���,J�nY�d"O��Yr�Qb�R��jY�si `�"O���$�G�m4�j1��3S��b"O 8 ��.�Zd8qh�3%,�(2"OT��D��A�
���T MFPL)�"OV��$P8~�%�p/�-�Py�a"O�%∺i���a��G�(y��"O��RW���O��� @�V�rxb"O�� ���0QN�P%��HԬ(�0"O %���`锬��� ��m��"O�Q��'�mˣ�]�@����"O�)kF�q��S�35tL��>a�D/l�j�˓^2d��`ފpr� �	J\w���	�{���%kkJ�Iy�ó��"n_��zв�
O��RG��|hE�C� �zA�"�IC��)ї݀h�q�.��D XKE��5a�:r�<��p�.��@H6Ş�~J����I�@��\1��G�<�c���8����u�%}��	ÉoL��p�;v\��	;0�0��� M��as���~��9O6�A0C�d*D����) B�]�p��T�f�������'��)��\�/������o7�Ű�o�4�i��P�Vu�2��֐X���T?�+�	�c�Є�w��-&~��F�\�Ɇ뉠_���S�+��0�iG�}�$}z�
E�1b8��5fmv��#�T>I���%��	�.]�s�"]نʄ16�#<1���S��\�T� 'hĄ��%����G,D0�.�1[�RŸӉC8�y�J�y`B��&El�� �sa˗$s	�VdKomd	�%hPW6|H�5�,Ŷe��N6��<Y�@M	=;2���)գ1��ʆAj~"�C��"����N8��h��;OBf0*��/=�RfjC�V���� l�"k���G[ %&6�3�|�]�J հ��H�nJ�	6ҚL\�ą�	�R��L��.��*��W���Y��!R��=!.xAS%Ў?E�h���T?�A4�I��4(��
�#�1u�4 f��x�<:g��P�W�#j�hD�~���0��	[��iW���WJ}2FȪw��M�=E���)VІ0�̜.���a��`e!#O��0��НP�����9O(�qrl�
g*���L�.���x�E�t�2\" %ΎL���'4�h��v��5�D���
���@G�v���в��h|2Y%�F����{�O%B�ӣM��"�xt[��<�	k�*�}Z4h*ւW���'��>� 㚖�R��`��|��,�v��8@��h��ԟR�	�h�V�y~�9�L]CM�˔}�R��q���2м0�����g�Hrhɻ~�^�iDb� t� ���a�"]R�ӧħAh@�$D�b����� n���Ja�K�8����<Ie�[�x%��b>�@ѯ�'��h�J��7��ٳ��)T}�Pz�����OR�i�&s�䘱c��ż����>H��Y�%N�/��9�x)�7�7ak��S��q�g�S��Ûybl�˂IF�݂Tx�E���G]�Uz�M�5�8��#��ldEx,��$�_��Bs�F���) ��2p[��^����t�3g��+��1K��NM$K��T"Ć��CX�5H��ſ7��E� �\��;�mN�4�Z�yG��~��I��1��#��L55�<��2����	O窨3��Ķ(��"�ʸ҆�<�C��QJ6�+���O+��r�M�f����l�^?Y%��;,�1G��'����o�	-H���+�=h{����?Hq6�҆�	{�>��cʾ'�0�]v����FY����ᖼ}��c����}��˕ ��_�n���Ba>c��'z�V��&��P\>�yKX-Pj6�r�{"�u�`8ٳJLI�d�����[�'~8t���H�v�%a&nV����K*j��ʧal�8I�Ď�;�'��32��i�C���7�&pG�c:���t�}�Tk!��O�jʧi;T�!a�=ڔs�'��*��=�\�f�AE�]G��ͣ)�TF|L&��V#�()���q�dL&��@��.?� �s�����E��'�!���L�G��AC"G@�l_ra��� �)��%{��dd����-�yw%T_>��A.��,�����@B�BT�U�SYdR��6CK�[�$��Ϙ��� �R�K࠘��P�L�
�����M�� ��"M"GE�B��iU�r8���Î���p�OA�]yVdb�"��������]�j���ȏ�l;��ɨA��e��M k�Az�-NOi��X@�I�_\��'�<������1��3,��4ꚗf��	HDh�5dut��#�xk�g��v\C�O�)w��$�\A*��Aa�@s.���篁_s�\���4��p��9~��Һ#@!���Ȓ�y�.��%gn��O�(��j&g�LN|Q���mt$�'�Sv�� i|4�$ΣbzF�ć�<� ��ѫ�
=��ڋ ��1iw�'��%���]屮
#�67� �{*�q�ҩΠrc��A ��,`�Uaq��O�j�&_ �BIQ��.���NS�0�L	xr�_A(�v&�\j4d	�Ą`�S����ߟp���]:58�.��x�:b��Ѷ^,�"Q��?
��iȟ'�'�c?����� a$�Y�O��x�fa*fcB)=s��H���HOh�'�_��a(bkR	}���J��X}�ىC�ҙn�z����@�l4�����䓀?����,��B���!y@���VC��.)� ���J*n�A����'�'\6�F/C=K�N�!�$q�Xh@I��̓b�D]qq��U�����ي ��)�E�5W7<�[񀎍^���
f�=O�DK�Kڹ(�ʠ��@C�@��1H^�$?�����4էO~�=�1��5;?X��0'C)���1�C\�3�]���5{�:�e�"6�(#X�9D�)Ol�=ͧ2��D�I�PS:��-��_
�i��_Y['���ΰ<��q>��FJO�d��Civ��
Q��Гō�
JZ�O����J�Z(�������q+�Б��>a�)��d�N��fD�cb���!�G�Ę�gF2Ũ��S�O>Q�D�	[�O�����q!ҵ!"Ï�$�U�i���7&T�v�Be��R�D=
`��������J76J�s��ŌSp�0t"����u�d��J~���|�f�ݎ*� ��HI(Qd��W8���B����
$ �������u�8�=��d���@���F~�0$��N�7�B�h`DR�/ax�)�%6���
V#cҤzu+�0U��_�E�x�d'�a��ٴjX�On�PK<��uN��@�l:�O�����}` Ղ���%��H�� P�E�U1#C!�`��P�-w�⌐t�@��V5���ݠz0��(	w��dE�*��+A�7�>�k��$z�`��Q�!�]ʅ'ܼ~:�)8E�(&~4Dr��$+6L��r j�pN�.8� خ�dI�Q%�`X��ˌG��ҥ��6�F)��F�2/����?��N�<r���zP�=��{E�Z:f%>�����/�ay��4LJ}�7C	 g��0�/��f���b�1t�(��ǃd&���>%�y�KG�B\x=JbJ��&d�����FX���GT���b��2G؈O�	��އ%���@R���>!�'*���B
,f �S��N:�C���
k�����������6����I�7~"����tj�ii��<TQ{�/��$"��>��`�R.±G��(1��_ ���ҕ��2u�C��	g���@B�Z=Y���W��>h��Sy"�|�#�4@Xy��P3}J���A=8�Rl����-���⌫_l}ڳG��ay�O�9?�9��o��`�a+p^t;nΫh���9��)��D�G����L�S�\��$ 50�t9 fދ(X�b��S��$�<��r�/(�Rd;b��<�`�۱c<�aI��5
k}��F��y��\A%���R�^����I���tPj��u18��'Ή�0=��	��!�!.�f���i�)�$Z�JA��D^bqO��Oޔ��G/t����XL5�T���	Z�ʕJ�b>�OX�	���t��EM�=��LCtA���Ґ�'z�O؄3w^nr铣o
�K�-Z��\7�9B��B�-L�s��a�a33�<�E�B����H��'X�M"� qӮ�b�h�<hPT��+� ~�S�'���ET=u�b���p��`�`����yR
y%�A�åUbl�$��"��$A,b�.�8ki&�����A�S���>��HEK�g�����=i���H��4T�8B�K�|�4Dն1����e�	���
�H�	�Tlg`���X��$��#Q �y��֋K�r�87"?�T���⛋��>��ꋋ\�l���咏u�p�R���~Ā��J=�?YSW	E�,��C�>O*TЁ��o�'*R��3��5K�l�@�6D��1��	"Q����ƺe�6M���,k� R���<5^���B$E⤽����AĪ�S�-�.
� ����C�䝋"
WnpK�]�v ��������[\R *@�V��d�s&:�4�k�2m�	R2B��lq�w[#�!��:~� �f�_(W"�`0v��P����� h��2�y�'(~�0!�&#�8��0������٘{s(�p⛚0�h��P�'��(өw���02�@�;�Х�RC�,pTtj@`�<A��[-D��Sա���M(���A�'�c�B]'P���1��X2����d��{��c��&h�Rܚ҉WYuv���@��j��d,,�\���;��8ȕ�F�Fb� $�?�O��a��]����F��u�N� ��'^8��aZ�.d�0[S�-`�� �e������d��[G���T�B�������%f!�d6l�E� O
�S�<Iz�C*@z�`���I�Op��{qăD�ԟ��yu���D����K����S��}��� �6G>���/�th<�	J;���R'd��t��0yB>��D��m
�t��(x�p�ֆU$!Q�(�6m����1����97���e�(�O̸���;�I��cW�����1P��T�J�v�c�	��k ���Ol�iÔ	���!� ��b� �GxRD ^X	Ѐ!66�\�ATI�=�?�'[6 rpO�=lm3􏉊n���S�?  L[ G]!^��$�0���z�"��҄e�T�3�T�J�z��"o� MY��9�(�B��}�FY���w��M�"O��c+�����юu2��џ6B�h�L�/?N��[!Q�z��)��(O�Q!��?> �X����` 1�0>)�n�c�3�K��fpVHA��Px��d��^�O��ho�4tXd�3:�O4�5�O~��dJǅНkxh���0-��i�wg�p<�ʒ��{W�	��ߟ�IJ�! F�"�2#f��st�  �"O*�[��M���2�k�
N-E�Z�uI\:f�Q#~�9���Ģ�*�Y��9�Ɣ�Q�1C�:A�%Hܖ?�8�d"O&5���) ���A6�%"��}S�oB�{��0'P)c�Q!4E�U~����(O�$�r��#A�z�@f+Q!��}9q�'I�	"��ӹK�H��9IDt�RǂJ'N�#W�^S����@LG
5��Շ�	,�� �Ѡ� �.8����$�z"<��hK=<6�B��Y	v��\sd#;Y�6��4y0���;cF� ��		pêB�	�R�,0 p�^**��\		YS��)�1d�z���&�<X��1��PQ>�R"�ڰ'�u۞�3U�&J�bB�ITwL���&R����dh�5y���Cq�ЄhȺ@a�`ƽ.F�X�Q�d>M����#|@���W# ��Z6O� �`��d̂��$��g�!^��2��g�L)�7n��!�d��2�Y�H��`yrƄ�p>Q�J	l+)��ǵ3YˁL�Z�'��%�� \�5Q0�˿f	���|j�FN
&QTɁ����i`Ĩ�͇b�<�MS	H�.><(�p �.=����AK9(1pU�ŏJ9gB��З�ͿqY4�|λM��I	C�D�x�H؇�}��5�ȓ5���ȣ��p�l��AdǊQxz�Y��ۮ|���	1��|������xҋ��$C�`��K�S�\��&K�o�!�$Їt%�ī�C)e]Ҡ)7�-B�!�0W�ֈ"���op�)��('!�D��2OZ�j��~c
%Е�7�!���!����S�1���cP��.w�!��4Q��X�7�ڛ}$q�J��!���C��[�a
)_�>q�3阽�!�B'
Ӭ���A�G�D�"�ހJn!��&K����$��� ®A
	-�!��#����E���=b�K7�!�.��]���t�(�u��>�!�䘭-�u�t䇈V�h�d�w2!��ȒJwy��@�n�t�y�ƹy!��C ^�YK��V9M�+Ub�0?
!�d�'<��rDI"a��r����!�d3�(}��#ٺp�4�%H�y�!�$��Zf�[G
�Fє�C#,�1�!�d_�b�B��*RR�4�
�#�!�$
�K�ڭ�e+�W���j��G!򄊡k@�y�/�.%
��0A�� X#!��=m���E�S.��Yb��		�!�DÚF�i�(�51Y�uA���.Q�!�,�
ij��1lA��@L#^�!�d����ɠ����l��r��B�!��L�	��	��6���m�	�!��n��@n CX �3��+�!��l�|\p��#%9��ӓe@�[s!��t�DN�5ƞ]9���!���Ȟ��ͥ��`ق-1s�!�D�	WM�"aD��b)�q H�]�!�$ݣ|���&� E�Tل�<�!�dM�:�~�0傀A��0ǧ���!�x�u��g��1����<~�!�d��o�8d*�%�9]h�B4g�!��ʂKZ��@�J��Q�.�A'�!�րw��( ��	40}6�iׅ|!�Д���*�-\m*p;�d_&7r!���kw�\�#�E�apxr���a!�d�&N�H%mу2��˱l��.�!��n�0DҤ��+\���
E4!�� B`��%E�o���˱�&���"O< ��#��t�d��5�:HyhЕ"O���k��\l�-�ČM�yh����"O0�q.
�to4ء��I�XBl�"O�0G�-'�!z�½6K����"O��
�*�	�T��!��DY� �"O�`�C�.D��1�I�G �:�"O�	�����(�����%6p0W"O��d"�/QF(�^�|�e�"O����͌�|��q�ƒ��Yx�"O*U��H��)� ��� �VE�p"O�TaO��%c�+�0�C)�-�yҬ�:LT�|"��@)�H�S�Cԙ�y�.,%�V��L� �Ai��9��B�I�3n��x�S���b�P۶B�I�Rd�c���¸��&��&�B�ɳ/g������
���a"�Y;؀B�I�BC|T����.�����#��C�Ih#L��F(A/u��27�.�\C�U��@[ �o��a�JQk�B�ɟHd���A@$&fV( �� QTRB�`��ŋ��Z�)�2,��!P1�(B�ɖ y�������G�\�5�!n�8B�	'x�XR�K�Vq��K�� ��R��h��0 H�$+z��Qռ���3�"O����H��-����/m����'r�P��09�<��gcL��(��'�
��r�I�(��C�48�ʩ��'��hDԷqB A����-2�B+�'�R�k���@����7��)�'��eR���]��L���ٵ1t>��'��� E�B�U�*�YfO-<|�*O��=E��h�;����,G�O��q����yBe�lUD�+��,pKPܳ���y��F
2���:��3���ׯ���y�*Q	T�����	%�����]*�y�F6@lpuӆ��*��F���y"Bߩ{�^l�p��	��0&� �y�e�;X����+��T�eT$�yrl��/��@��LÇxŔ�bK���y�LA��4��#2f��i@�a�!�y�(��"�hE�[����s���y�MC�I4҄�V>������v��I{<�⇼�P�a���! �h1���T�<���ȏeX�ʁ��?ޔ�u��u�<�0"
�;�j�C�Lj��GiHq�<	V�ŕ{K<�3�ļ}����mTi�<�G�P/�~�{�gٳ9�ƈ�V��c�<�c��C���A�P36˃iY\�<ICa[�zbAF�$�,�$�KU�<	���wT��s�զF��*l�P�<yj�P L顃 J�U�8��G��c�<1��I��nP{CG2#H4	��z�<�BBZ����D��9@�iC`K�k�<م$��q�v݉��Hf��f��c�<�u�B�=����/H����tI��xbgժqJI��GR�q����a��M{�'����dm%A��01�؉!(a��'��z!�ʧ&���W"� �z9y�'i`��腹c���SE�E;	'�ɳ�'`Թ����8>�}x���,*d&���'��d>�)ڧ����Ys�xj���j7��ȓ�q{U���i�i�D'�`$���'�ў�|�w'�n��(K��J5ZF�@* �h�<� �k��&Lü�#S̕|b�°"OX���O@&��B��љ(����"O��+�o��;��庐#F�e�H-��"OXp5V�f �P��g����6"O)�T�#�G��E���ZD"O��K�6T�xk�e݈�B��S"O�Uб���M���ۺ[s�]#"O�q��O]:8�PQQ,�'gZ��v"O�%�SH=�t$��aQ<��t"O���3�M�l`r��w�ёXP�TS3"O`��EX'��� �<^�i"P"OR=����}�r`��I	((�"O����º �Xs'D�_�jL�G"Ov�H�Q�%��e@Q`�B���t"OH�FEU�k�P���h��F#�Ĉ�"Od����I�$����s�W)w	(�"Oe�.֜9j�q�eD�=.�ʢ�i�qO��)�3?����QE�xR��)O�;�Ps����'	��u�6y�T�C���-�U:�'��U��00'2Q��[�&��d����y�7�
���c>@��P!��y���+�P�2���z�gI ��yªP8{��0���,L� MfO���y2�ͨRK��"�hK�<��I9%�Ѣ��'�az��^�.�����-R�2�A���x2�% :��`l,��uL�_�C�	��%�"ִ��L(E���B���|\(�b�+Ü�s��&6��C��<m�Q��C��*�,+%(
�e��C䉬@������X�h��l�4 �C�	�k��S�lע�`��d ��Y)b#<��	�R	��K���K��G������b�8p�r��T22%�-g�@�ȓߞ��Q!�(IV(�x�b�P"����|~���O ��gH:h�@�e�~i��IQ"O���t`ʳ{ª����
�Jv�r��	�)��>E���RX�ZA�6�%{܌�Ԣ?D�4ye̓7y�A
�Ys����D�q��mZ�t��O?�а�~�Ĺխ\(�1��<D�(R4 �Y��ӱ'Ѯt9�a�<}"e��d�a{�#i
�`6Bh��ⅡS�x�p�<�����7����jܰ�����"O�`�v��=v����3��XAU"O2d�a�h�Hr��F�<ݑ�"O�|�q��	��E���|d�	�"O�����M��x��ơ9b �"Ob)yDIN u1��h&�;+r$'"OH��+  +�D�qP�R�<�F"O�u�%�*vbH0B7_���2P"O&1���C%Mh �0ơ�1Sd�`"O��� FU�:
x��4�8G�"�"O.�[��U�P��+G\p�"Ov���b��"Ě�B!&4��`U"O�:/"<(A�M�>�@*S�3-!�$��z@]��-�Z<��/[�2!��ԆG��p@�&V����/4�!�ĐL��xʶ�N}1ڼ���ŔX�!�Ć+p�VL�T�O�& �る^T�!��$D��*���а����It�$%�Od8�j��,Pe���2ƨ%�B"Ohp!�#i�q1f�ʧr�h��!"O�����7>yg�E�m�JEР"OZ)9W H��l��J����;�"O֑	���zU�f��[uJ�`�"O� �кP�W:eT<��F^��aC"OBQɳ���K���a��~o p"OZ�H$��-8�9`�J^�x�"O:���*�3Z%��)�q��P�"O��I��ߎw��IfC�1����"OZ��؜]\"χ?��,p6"O:��f�9!��YY���.Qt�a"O�4�K$<��+�f��6"O$(Q�hI���M��zt`���"O8I����F,O%np�k�"O6,����x�p�%NB�*m�i�"Ox���kK�X��T솆:�+��,�S�'�A�Fb�~�rR$C#aA^B�	�f4Ċc�Q&rO��A�KrYRB�	�v���fg׬N��$1��d��B�	$i���Qm�&FtP�#5C�-^P$B�	'��� F��G��b���4dC�I;V��8W��J8�%�V�*R>C䉰�J<�GB׍��e� FӔ �xB�ɾS4J��&���Z!Y�I�a�C�I\нZ! �H�X�"��E�B�	�5�:���,�!�Q"6�݄c��B��(2��jQ@+ �@у� ��C�	�G��=��H��\~���4��� C�I�� i�3AW�P���dF��t��C�I�muj�@��5�� �(�#C�B�b��H��%�Y�����鏘O�jB��/7�R1F����k�,��:B�	
j\���N��1��R�\C�I�:M�}� KenT�e.ƕ!�nC���  ����[˜�a�n9S��C�Ɉ��acff�)'�9ڴ��� 'pC�I=vj���I�+���Z�ԛN��C��!o!��`e�g8�P�cS#j��B䉚E�J���E-���h�k�V�B䉠6�\���8'��b2��8o(�B�	�$�t����0<��y*qH�N�jB�ɟl�`�@���d�C��H�
epB�	�;U l��҇b�I�+˛K�LB�	;�9��J :w�T��g�"6hC��'�΀J%�O2PL��h�-EʂC�m�8ԛ؀$vBh)DM�x�JC�	ih�b&mH0	��EU>��C�I5����Q��"@�*%�C��.�fɻ��)�ܡ�%O�4�C䉮f�D�:����;5l(Ȓi��KttC�	�?���`Ø")�I1u�=tFC䉼y7d@Y6�
��sFb�/?����'��4�FЧg+���l��8.,��'��CP��?_�j��RZ�*��	�'��)k&+���Ҵ� W\�i��'�v����L3_� ��CO��L$���'�6�A2톙lyȔ�4V�21H�'K���#$�``���]�a�h��'��qe�] OX��b\6'��
�'��x�RnB�)e� ���=+>�;�'�̉sUB�&�bl�+�;c��r�'F
qi2A��,��C�O�.
p�J�'e���UIL�R��]R�gC)#����'�D [�M'(C8	XuAI�h�z�8
�'�°�� �P
eBj+5\&��	�'���R4h]q�<�x��R4&k8���'��RV*��+b�BQ�5h��u�'t����`X=~ܔ�2��9_N�|#
��� R���YS*&#�͜B����B"OR  �%�1�6���lJ4��y3�"O����nX6&/\���(1����"O��:�5��L�(�l��"O6�#c��%5�j�!gAU�N���9!"O"$ R�A�}��b� �|����"O�,`�	&.y��Ю�.��H�T"O�mzv�tl>�[� ��u#"O���q�46��d��D�d�!"O>٨#)�gA�8h2��hb d�"O~�ӆ�LZ��)� zCb���"O<=�d�u^<B���$
a"O@���f�(ՒL��@
�n��T"O(]���G��dmj�A�9�HIp�"O^I+� �%B�	`��X<'{p�z�"Ol�Ju%Fj���q��\�|""O����B�|�PK�K��"�§"O���2.��T�
͢`�B�G�ָ+�"O0a�؈p���Hs+ܮ��`҃"O^da� &����u��:�*œ�"O:�`��ŴrJdL	�*_�w����"OP��dn�7��T{���t֡ha"O
���B:(�U� �U�6 zW"O� ��L� HT2����� "O&��QD]���۵�ݪ;����"O��:A��1����(޺*���"O�]�q �2����vs>��"O����֩k{��/�.0�6���ybcQ6k2p�"Ŭ"�l��e���yb��C1l�{��8DC�%)���y�h�?ߘ����A�9��11��y���/V���[D�K�6�&��E˿�y�7?:�)��W<2.R}B�

��y�ȿe"<�E�&��	p�S�yrG�#Ȅ�g�X����ӆC߄�y%6o�^|(3����a0�C�-�yr �=G
t�J���$�Aq�k���y�N��)SP4 ���>߀�@R��y2m�;��@�	�� M�!����y�HFNh\���
E��n��c��y��I~���1����'R�˰�O6�yb�ے
c. ���|m[U�X��y�D֗U��MQE Z�z�u��-�8�y"$ݘ�J����*bj(1h�I��y��K����Cg��VL69ҁ[�y�施Z�P�a#��V������yr�P���ʕ��JEL�a�/P�y�ǁ�>/�D�eH�=���#nI5�y��a��g���;�r���h\�y��ަwx@ ���G22z��St�yeF6��-J��ӳ.e x����y"��?Z~��!4�n���䓒�y2+�<~���Sv��14Ԡc����yr$�4�
�Ct���p�!��X��y�Ŏ&��g�)l�F�V�yr���"�qŁ��0�h���y2
�*��pD�3!CR(�(î�y�A!���`�K�5������y�!�=Rh쁸WhѮg��s�� �y�Iݦ P&�ic͂���I��y�.WQ��KRD��;��7�՚�y��׍xPfq�7Bۦg���#g���y�JUI�YaaJ�\�ޭ��a��y��Sk	[� 0T8�5X��V%�y
� �Y�������.R�mȘ�b"O$U�c�C�Jt�V+��r�"��P"O:	�ȏEr�Y
�G�'E���"O����)E�G>��J�@�$0����"Oƀ�3��:��0o FyF���"O��j�A	l���㇎�"pOPp#�"O�ɬ�Z�=�A��5Q	�����v�<�2�Ȓ!Pp�KS�y�(���j�<9�+A�(U�(�6+��j!h�T��Q�<��Y�F�VP ��� �@hfIY�<��j�>6w*4j�@�~0aR{�<�M��\�cT��AV�S!�x�<�[-bh�0q�:vH(��Et�<�����hqJ�S�}���EE�<6��yy����GHeL�e`\g�<�P��;ql���Ɋ ^�N���e�<�4#�+��-��艼f/v  ��j�<q!�ۈwH^)�7#Z�:��,c�<�&�F�	�('<A�e�<aw�\c�X��C�ז4>�@��e_�<Y�@"l%���!��gV�@2�X�<�oX�5`�d��L�}�z%b��OR�<).1S�Z`S����2�q�h�<A��Y�.`a{ W"o"��Qa P]�<y^��XF	�58�a�M˓DYH���B,�}J�c�:\~�y:*�_�L<���v}����;��T�.U�YL@�ȓP�f���
�1�N �4lG30�RP��j����C�I�]��dõJ��^%�цȓ}�^�*dXi����A�[�:���B�� ic�?(��s�HUX����ȓ Dą)6b�$j�(��ve!.
6͆�*�.q!��ձ`TDyV!֞��q��
�N��F's�٠1�U n�bm��jR}��O=f����I! s(|�ȓ����ޓlѮ`(1nM|�0���e�첷�̵��|��L�uWf��ȓnAL)y�'E�>D �)�/� ��s2�E�^KP �B�1K�Hy��.�ۦ�[��5ؕ �-��Ѕ�HŲ`@BO�}��)v�	 M�le��K� 98�F%�A8]�R0�ȓN�D�!$��Kӊ@#�A�1!�<���~�z��7��2R�ά	¦��2-BY�ȓqB��d�I+M��Ia�@Z�a,�ȓW4 �I�H�'�<]�P���A�4��|.d�# ��%aV����XD��i.�}�GmS.v���z@L�>S��y�ȓ*��}s���0��,R���P�u�ȓI^����E�+N�)@��C�8��P�ڽ�'Dͩ{�`��6�N�9�0�ȓTN�	W&�\İRF��� ���T�.�R���]�H���J�;o|$��ȓiH�����+(��!`��Sr��ȓ�D̲w*W�h=�x�`�>1�������X�מ����B�/y L�ȓ	^d��a�C��(*�n�	�V���II�@��@�
Ay���nB�%�ȓR�¥2��Wj��<�����> �ȇȓT��%�#��-�:�a�)Ί�ȓi�JQ��H���|	��> �X�ȓ
�q�c)D/T
I�v���v����&pƬ�ԯ
�`	��XSmĂ1��h��A���ƆL���� 2^�u��S�? ���x�du"��j$p5"O���Eμ)Ԃ��F͝Jø�"O<�[�-3�4���,S�B�����"O�8˲lV�;��˂F����i"OZ<C���vR����V�{�೴"O ��A�ѿ�]�/��$�@�f"O\�
⎑z�X8捅$�P��U"O\y�p�	�}�����^F�l-��"O�,q"�O=�����q�+'"Ot,zŀ�'+��a7��c_x��'"O>0\n��[�쀛$_E�5"O:��p��)*�͙f,�^�=
"ON�Z��R���m37�A�?� �"O�mHf+�C���g�;f����"Of�	$� |A���e')�R�a�"O�T8�@��Q��cA�h��� *O�ڷ�Z#�!� ��W�p�J�'O�cӀÚtҕ�'�ʠJJ����'ZTC��[��P�W�	�+ ��
�'�|�f�;r�^ b�BֻUi6�[	�'Rt�!��M����	���=�	�'l*�����~�*Š6��v�Z	�'^M�T�T�N@��9�i�hx�'TI	�Z�"�e���98�H�',L�C!��q�	����y�%��'\���j
��b�卜xx����'?Ԉ۶�:	��Tð�Φm�x�'a.��7��2m[���E�L(Rx�	�'��B�!���-\�6y�'�j���� @��j�Z�Sy�x
�'̎B��}��P%�ͷ=Ȓ]s	�'P�0�х�'8�8�Ap�L�?���	�'&�-�oƾ��T�&�'?�\-		�'�x�_*I�s�+�Euy��'�����IPi����B����'|��An�p�(��-�:@�z���'�jhk��@�-�a�ɥuܑh�'�(�Q�eK"%(в��1���c�'EDcTGŲSh�p��խ����'���3�喋;�$B�g
�=��� �'�.,��a��NAI2D��jJ)��'�"�xeč D�4��Î7o}0��')��"��%��)��Hut��A�'�н	� �4��8�`��q}2!��'!By���Én�8$�-�q�0
�'HQ�i/�����j-NU�	�'����ִ[���UĈ�3�L]s
�'�ؙ� /�2�b��TҗW/PX��'.J�y���2t�Ҵb#�Q��HK�'���TKA�S�@�ML�y	�'���q�M��p� ɕ
[�H�*̹�'b.�8p�x��L!�� .Am��i�'F~��d��XUh��N�/A�q�	�'َq��o�:u�!c(����' �ic���-��9�@�P۰��'�^ S��q%z �p�5�����'�L� Ę`Զu"��3�aa�'$�q�W)ʧOj ��%2��p�'���ٚ_�5�g!�"%3Ty�'�D��c��]_\�+!E#e�p�Q�',&�#2�
%-��e���<)��'z�Yfʑ:>��ݳt��|8���'�*��)�:)P$��Câ3K2�z�'�(�C/ѩCxP�N,*�>	��� �С�.3(Qʐ�YJe;$"O�|pu-�M���qbE��~��m��"OR� ,I�W<l�c�c�4l�$�Q�"O�P���3��Q�)۵fN��*�"O����B&JU�D�(D؁��"O,�*@��n.R�������晹c"O
q� H����ԃI�W�J��%"O� z�H�b���gh�T�NA0T"O8 sAN�0up�ppag��z��P�5"O|���LN�n0 ���W�|�Y�"O����Z�?�2iS��� I�%�@"O�j2�Z�eA��C�j�LG���"O���6h��2����J�1D���"O",`$T����]�YS "O0$s�
!'�Q�B��z>��$"O ��sA5j$�5	$!ɰA*@0�"OV9�G��A��Q@H<$��"OR�PҍG`L��g��=%�J0"O<dP�n	�<g�Q�	E��fI�"O��d`Ӂx¼ġ�. Fn8!�"O�AQB��_q\�s�NB�FSIp"O�s��)r0q����kNJX�"O$��%k�1���IĴ	�f�X! 1D���#��Q���!}�YV�4D��"�G~� ��VHDF�51�M7D��F�F�q���z�$�
m_D5yuJ5D�� �N?��鳪 �4�")�+5D��0r��g����ݛ/7�%��h2D��KV��)y��8@�[5"-���.D��q'N�$HV�	H5�MO��I3�+D�`x�köC��9����^�� � �)D���d՚���J����}h�3D������o򑪦�זYO�=��/-D��b��0�L�"�U�ct�ӧ*D�3��A<ĥ��AR�b�]�!$(D��)C&��D��A�Ӣ��#�.�2 �&D���H0yɳl��� IQg &D��37  )m�>�7��b�a�L.D�hk� KV��"���D?��%�,D����%�(@�(���S(۴< �/D��Hŝ�~b�q#C�nv�|�R
-D��s�I�+Ϣ��@��9Z�t�3�/D�h� �\�V���b k�`��#0D�r�ʃ���(S��)0lRq�2D����ػR��4�$�˭+�D���:D��1�n�d8r����"C�#$D� : ̒�=�*p��I�f�`aX�l.D�[d�ߺ9G�tʐ��+/+�ȁ�,D�PC 1sb��
���QΝ��,+D�$r�L7!���*�ףҬRC�*D���j߂i���@���>ݮ$��,D�@;�C^y��\��i޵,���5�(D�t*dO
'u6|����=Gj���j'D���V�άl��8A珛�Q� 1��$D��q�MY
R��Q���y� e*#D��8�Pdp6��3aԡg�uj')5D�thBK {Z<��P�{H�h�M2D����ܬ'��2 �?A���j �$D�tX�g��wj����4�i
�
5D����1�T ⴬��A�r����8D�̀ϯv;��b6*�ohe(Sb5D��A�����@�̩c$]���2D�P��L��lc��pT�I-yL��3D�4D����%�0��]�vUrhvIq�1D�� �H����/K y��(��-U�x҃"OMz�Jcָ0i��ՕW��ۂ"O�zAa��n��� �aA^xJ2"OT�pP'�Ƒjs��5l�zE�"OLIbWM�	"�� �u��dР�"O$�(gaz�6h���	d �"OLܒ)�7F�tDx����X!B1ȇ"O����n�"T(	S'��
RDk "O D��#F?MyT�y�ƛ;�9��"O�0��Au�p�R�E�C�QK�"O��
��PK���B�5x�K@"O��N��c�d%q����o�!"O����tj�T�HeFT�A"O��	c	M�>HയQ�/K�x��"O� j�B̏M�h�N�76ˎ%Ð"O���֮W�0�؀D�L�(9"O�9��E�"�Ƽ��&\�)CV\j�"O�����7���Hv��8c%Dx�"O��`ƈQ���h9����Nh| "Or� M.{�d1[B������"O�����[�n*j��Ҫ��t��	+W"O��+�G].$��xzE��Gy�$�6"O�Luً<��I 4�
8e2p��"O(R0���x(i���30|���"O��J靂_8l�V>||M�"O����V�]Lű-͹^hT�"O��_�]F��$�I�c$(#�"O�i��&w5�3�h͓kh� a�"O�x����'�����]�H_�	؂*O�$Q/�	G����ď$�>�;	�'D�TC1��[
�{DHͅkh�
�'��!��P�8@!s�C��.i	�'x�pBŖ�B�Xk2��X0��'U�<	�V�/Qh�����tB�	�'\��i�#9�Z!"q��.�z�'�H�$.�D���C �� "T!	�'fx�(��~�T�����3u�H�i�'�(|h���n��T�8Yj@��'H�T:%,Z.jw�����e��|��'��ʣ�
��+��α{�Q��' :���PYY8�����{i���'�V���d�:p�|MC`��cW:i��'�T�j�j��'}�zb�F`�����'����fFOu�̠�YkL���'�9��bIL"����ڜ=�L�2�'94A1�D����)V�P<4Z`�#�'��]��o%D�Ԅ�$a���i��'�vTiBj
�Y�H+�,P�}	�4z�'�x)�m
��L�� U$�|%	�'���������#3�����'��q0�E6c*\h��6�t���'�P�BF�k���{R�ǜIh�(�
�'�P��OO�j8�|� ��C�T�R�'�%�
�3P�p� �J�Fy��'R�s�K������c@	D⌀��'�6��dI .��̡�I�;9�,|��'Ҫq���݇|K< ��iۼ,���A�'I�R2��*�ĵZ��]z��a�'���oL"1L�`�$�(_�A��'�f�n�j6a����6O��T��'N�����-}��,g@�,E%�P��'a��Q��L�	ˬu*6'��5ʠ�
�'u��ʒ��d�\s��3N�\:�'�f�J�B�GE��
��6���h��� t��@H�J��lh0$�>+��U8q"O�=��a�0w��q3��p�6m�"O�M�P�ɫc���w�Z�k���"OҸ(��)b���"J�T��$c�"O�9���;wO&�C��`�D(�Q"O����f�2}� ��g����"O���E��&�ƀ� �4@:Y�"O��B�/���\��נSKz�1�"O������C��aٖ��8ЀrV"OL��C��-�LAɱ��d�� �P"O.�)W Qm.���
6u��h�"OlY�C]�fxD�B2Lk�8+!"OF�qṔ�f�����N5�I�c"OF��S E����D`�A51�"O��Ǣ�1^p����{����"O�$�
@�2w��#�o�'�2���"Ol()��0�$#R.N04ɞ�"O���֎�p)"Ac1��>	�5h3"O�=R�O�?O��x��ǅ���""O�5`SG�I7^�!� pi�v"O����"���X@(7HÕ4T&,	�"Op�q�h��]��F�!J��xX"O��×�Y~{&�
�$Y�IA�
�"O谺�Ժ,�L@����<�¡��"O���U��;��#7���ܑ`"O�0�1
�0��H�H��9��"Oy(7��7�yAH�*bʈ�[v"O�Hf��?P��r�@����C"OY�U���^�:x	d ��X��u�"Oh�A%�J4o-��[�� �&�!6"O �:S�ȥGP|�Y�b�����c"O�-kT�%X�$�p�*C:h~
���"OH�H�J�v,�`p����4o�y�r"O�`ʥ�C�w�Lx��*7I���C"O\�t��$U�n(��X3u�T"�"O�-b���T����xt$�R0"O��0��/����$�-s�	!4"O}A/�4f��q�-ilX��"O�̻!�6P�L1!1ǈ�7Z�=��"O�dy�IZ1���Ŕ(Nz���"O�X��F@"<2��%�#��#"O�Z�Jñ@����c�&��4I5"O���sF�2E�Ւ�C^F�����"O�<is�Ɍ7�D���7x���B"Om��.�,!�����C%`t��b"O𸀢H�>�8;���]f�B�"Ojբ7�Ƥ8o.��� �/)[�1c"O4��L��F��C�'Z�qZ�'TXi��:@�HCҭC$m��`�'����(��?���@U.d��,��'�����i+
�b1�6TR�'��*�*��	AdȻRm�|i�'�$T��
B�LG�Ppu�ÕP$09��'5v���͋-#;6]�thJP!|l9�'�� ����h����N :���'֞��&�A�_���3�ǮH�:mY�'�Ҩ�qA-��â�'M����'1h�4E� x	�oQ�u*|I�'d\�7a_/]� %9�Enڈ-��'��<�C���{8t�z�f��aV�@�'1�e3$�R3�L���F+WJ� �
�'�X�I���T�p�����R bIC�'p�h�J�Qb*��6�Y�O#��'���C�$�m:��O�4��S�? 6-��CƸG�|��JK1@��80'"O�E�T����X8��i�64`;�"O��Z�A�+fUFU�ǖ	��X"O�l�kC-Z��xp���m�l�3�"O�M CL/��і�A3N���z�"O���I��N��h�()��pV"O�H����=Q����N�:~�E�"O��0�� !*�t��͒�hu8��"O2H�ƣ�.��5J��,ck��""O|M������q��DW&l�"OZi�u�7�NL�C�I�RƄD��y����8YeB@�`�@��EG��>�6B�&��b�H�:T�TI�v#ŞI�&B� S 
��K�,d�R�#�IB��"e�Y���֎����A��`�C�i��%@­O�]�´r3 v�nB�I�w��Я�;Ą�e * NB�I�L��h@"F �L���-,�"B�I����7�� }6����Lkz,B�<gKru�q�Z`�d����
P��B�I� ��$�#> ���MF�H<�B�I�
̀m΃shDm�$�!E�C�I0~�4C�4&.2�K6p��C�I�B�.̻��ٜ*6�x�e^�9�C�	���-:�
��V��c<0�C䉾�ʑ�4# �/T���ãXGdC�	5���Ӗk�r��:D�Y�39pC�I�x���hd	<)��m��X��nC��������,Z�1����7V�NC�	�s��yz�B����b�(%�$C�I0:�B�s7D KV�`���2>8�C�I�/��S�,�)jr��Ӂ\�!�C��"$���i34��g
��m
�C�I�A�4qu`ݘ;�%�%�[7r΢C�I.�N���B*@�r��ɗ�s��C�	1l=���bI��Ll��1��i�C�	��hq#�^�~o>!�c�T�hB䉀? �E�Fm\��4[�(���C�$l>����N@ ?���&ܙ!��B�	�]��}���U��}��L��UPB�	u�8u��jȏn��-s'B�<*�B�a�d�T�I���K�*���C�a�D�`�S�o4� �E!H|C�3<��tK M�V�ȸxFL��dQ|B�I�Fy(r��,]\�@µ~h�C䉏|X)h�n+g����q�nC�I>lX�����:a���bC�ݾ8�C�I4� �;�ӞN�~�ñ�	5��B�I6*���V!�:�Z��ަI��B䉍��V���ˇ상y��AV�*D�̸�C�&A�AhB� 2!�h��%'D�����Q3����a�$��=ّb%D���!!���.ar�ⓣ ��%D�`�CA�&`{je���E  )%���$D�T˃ �x0Lmh�͟Z>���h!D��[@��5}��I��G�����
!D�T0�n� V6usH	�$]9�i D�d�2��5f�K�K���t4D�l��K@&,dr�і�K�u��RJ&D�p�c��*4Gd�����R��|�f�$D�H�q�ؑe�}��ӵeXd�2��"D�`�o@%��@H�j��2�V����!D���UAB����"ˈ\� �jvk$D�@z�i��6d$�E��}�"0��H-D�� �;�f�Q�D��,�6|��i"O�A��K&�4���eG�J#�Y�t"O �s� �V0��R)vH�k�"O��tm�k��h:����B�"Oz-���׎O����ʐ f�pA"O�K$V�<�1�T�;�h��e"Ojec�S�<��4�( Q4"O�Mk�	�o#�q ��1���u"O�9���v���9�G�d/�e�"O�D��Dр1�/���yJ"O&�(ኃ,K@J!�u����4k�"O���욢!��Ԉ�d�G���"OdiZ�]�d�%8\U�B�!�$�o������5!n�z�k3F�!�$R�n׶-�g �e�R��I��!�d��gD�qׯA7;�T@J�M�`!�$&��I���"5�v�[v��-�!��U��2,��ɀ�d��a�#ԫ(�!�d�9Ay�5��s�:p�b%S�!�DN2y���y��� )�53�(��!��&rU���w�e
�F�e�!�)MO��P3���+�����GY5/!�$�[M6����G(j��`�M�8�!��[~IH9a�@�����V�~�!� ���(�^�R��t�Jy!�#X�B# �&8�"�سTc!��@0`��?8�F����	MT!��Ԭ��A�6=�f�{�*��.l!�ą)\�H0���<�A��x�!�dW%#�Z1ju͒�P��yu��->�!��d��O�!r�n�8�B	�!�D�;��� kˢT��`�hƣg�!��I$3��9ca�>\g�$��_�!�Ǿ<�(F�ڄc[�[!��\�!�d�:�B�J�[>_�"�١$YxO!�d����J��� H�%a�[9!��ӏ{�b@ʃ�Y2���q��:T�!��k�!A�?�|����)�!�䞸|T�P�Ǭ� c���J�=�!�+}�X+��z;`�x&Iǌ�!�$��`��������툃l!��E�b��-�$���Q:��'l�?�!�ē I6�Q��ʄ�*��&�"r!�X6y��ij���@�£��3`d!�ҹ8���	�%�T�Ġ���_]^!�TRR�]�E%ő.���Hg��?\!�d���8�ͿJ�N�{ak�8H!�D�7(fA2��#M<�:�#�[C!�D�9����ɵAJ���_;z!�^�3��A�Ik�:+�,� /!�D��o�|�&�z*�r��Q9"!�$C
Wjn08��/X-,��\�J!��L1	-�]S��=IP|SF	��!�V�0��!��5	�j���"�P!!��Ȱ.��T�@�j��@j�lW�(!��??�����W � �+��#!�$�=�Rd�w�8إx��K0.�!�����+��!��P󕥇$f�!�f|V,Y«_.3�������{�!�d��:J��Y�"Z{@�7eרr�!�D�Bs}�tg�"�����р8�!���xy:%�D�9�ؽ�@�M1V!�D�VM����'��Q�a��|n!�d��x��0�U�$,�
ͳ!�� �lۢ�_sz�	���qj� ��"O����JM�ʶ� �VL���D"O�\�RM!oGƐ�Q�Sv2N��"OI�6
�I���bLQ4I0���"O�us3m^>>p������r1��h�"O���3A٦U�0�AHIO����"O���S�w}t���!��G	�|X�"O�A���;d-�Ga��儸Xv"O8W�4��)�O�9H�h3���H�<��Z��Bd�0B�:A��Pc�A�E�<Y��K�O�@q�(U�n�Ԃ�k�<��-A-52���E��f9B�����_�<�&J�'��I��L��A��GE@�<y�d�����^�/�=b$m�p�<�D�����T��4O��ҧFn�<��NT�D�[�E�5��p����N�<IG ��	��81
h9ؑj���M�<i�'M��-�b��6g��@:Eʆu�<���-��Q!FW/_���r��K�<�h?�(� ݧM��-�U��o�<	 &���Υ�#��*���Y�D�<�_�.�i��3+��ѷ�Y@�<)q�B�6u2��®ؒ1!��_~�<�2�H�2-�I9����cĤ�U�<�	�i��= �-�m3�E�Q�<�v�UU��s$��=��Dc���I�<!!�B�k�0l{� �C��S'C�I�<1DGƖ�� �"��Q��I�<鷫WL��\x�g�$���[�<Y��Jv��E�l�(�p�Gb�<����:3N,��לd��AQa�t�<	!.�1t�03dF\���i2��G�<9�ҨX �QĂ�Hk���3�C�<A�Λ+R1�(gm�F�Qy��M@�<�wJǩp�X�Eh�?��Gd�B�<�$��2!Bm�agŊ� �@�<!sj 2Lna��$�C�,��T`�U�<�A"A�Z�8�2�	�N���k�L�<)pa�7� -j�FٍO��
�C�F�<!dj��>9����,���#�Y�<�ď�~t�Ʈh�,���H}�<����nC<���R�}���r�<	�惶)%F (���i� mqg�
p�<�gH�`Q��H5 �|q�In�<	a�F9���Ag�.ttq(2ȉ_�<��גG�"DZ`��J
�#a��Q�<q�`���2���8��	 .UQ�<q��P$$7J�hEP
�&�j���u�<���	}��8a�L�g"l�x�!�p�<!B	�6D���dt��q�VC�l�<��T\N�H� D+����b�C�<Yׂ��]��yY�I�.>�c�G[�<�Q�D��|ۡ��0fԬ8�d$�U�<ٱN�J8��U鍕#���)��]�<p̐�w�&��a@Ў:��5yv�FQ�<���Y=�u��Q�vՆ�PKZT�<�Piʥ$���6�R��.p��[�<����t�)�։E�t��qєf�L�<���ܾ,p���ш�z7����H�<Q��R!v|*���l�E���F�<y�lݗ*kJa�6�,$�w`CI�<Qc�	�e|��`&jy`5r7�AD�<Q�-�ɦ��G�]k�)vF�@�<	2腗(nuࠏ�=�H�b {�<� �	S��;r z=zV��I��Q�'"O�p���S+a4M��B�P�V�i�"O�xq��'u���1�j��|��l>D�@�¨�!�ǡ�����J7D�:�Y7-�B�x�׆{���G$7D�Hh"��	r�@��u���[#Đj�i3D�TK��"�^x�ŦB,q��h0�&7D��@�!/�pO�In�뇏3D�t+�c�Ѐ����AjU���4D��B�2CP\��1��j�.i���%D��ca��O�X �]�u�-arN$D�4BF�<`�f�!6���AL*Q�f�#D�D��)O(�8�f;��`��a"D��*�l@	��DZ�B�$���G�,D���6��QK� ���ب2�ޔ �(%D�8z��\�EU�HV�בRtp`�"D�<@�	D"Eցȧ!�46r��5D�d�dOL�b.�IS����fjSK5D�`��l`������[H����2D�p)㊎�G������Z$��0�.D�D�p#Z-J,B}+0e�o����!�,D� � m)+\��p��W$n{`,�'f6D��2s�ɜ})>-B��%O a��3D����
	=5$���M�8D��@�)3D���a��3f�H�����$�g�0D�:$�
}Z��k�*��j�R4�3"D��w���ee�!���C!,��!D�ت$�B	2]K�����:��$D��krD�+̆�YAx,
��"D�py2lI =K���7��k�<Lz"�6D���@�Ґ4�x� ��
C�d�0�5D�t�$^�Q�②��C�7�ZPq�6D���QlG�Qd�3�(��)�R���7D��`�N�y�\ ��4:�x[��0D��[�L�8����I�z�tC^<!�D�{��piab:2�L*��4oO!�$T�W����M�Ij ȃ��0DE!��םb���%N�FR �)��r'!���p�A�Eʁ@l����-/!��v�1���1.x�y�$/�!��
%���l՛ (>��P�;@�!�F�:��(٠���9 ���J�=*0!�
�.! �古+�,���;!��C�s���#��	-"!�8*"f��f�K�$.HvDFJ!���d��� u�]6N�¥�\�w�!��ӁT(A8���</&�[��1HB!��#E�Dl�C�.cNJ���"#�!�Đ#��9��J�i�)�RbX�H�!��D(�0�[�ƣNe\;�Ɲ��!�D�{���i$���oU:IjF��!�dɻ)���2�*�Fqi�f�&x�!�$��O?��ڶ.�;�йGƈ%b!�Z5i����e�kq�]���P59Z!��@$q���vk	8S;���T/�!��\"Ug���b.�F"�٪G�H=|�!��ͦ[�����+X�Z�g�:Os!��=�rfC)8��A�mXS!���}�*�5!\e��I����O:!��Q�!ֶ�H���&-er��^��!�D�8u�	V)S�d�
���a��!�D?p��0�� ������AX�Fz!��-��\��)�;(�� h��Ȭ\`!���k��t{�j)=���c�A�$_!�� ^�h�@ޞ-�,<@6��,vZ���"O��15!_�p^�2�`�y�l��""O �Y�K�(B�e� ƃ6l��is�"OR�$O
�;�FL�e��5)��}y�"O��GK��<3�U�A�"O��R .^�7��Q,�4>���
�"Or�� ��4 ��b�-u���e"O�X�'`��lj�*ݑu�4A�"O
�`�'�1e�1�#�?E�x�c"O���I�V��)�d	��D1��"O��2�j�?n,�}06�9N�YR"O��A�� s�]���c#j�"Oe��AN�3j|���'R�� ���"O4Z�b�l�$i�&���M��"Oz塱�͚.�$���⛭.PH3�"O���E�C�w뾘Y���(����V"O���%�5s.� ��/�Tj� s"O$H��M�Bt�LC���	TS�D�t"O|��7�Z?2��H�m�,/TQ`�"O�� ���R[�p`�,Q;Nx��"O̅h�I0`�^�Q���i#��0""O��CЄ�Z���H�N��={^ {A"O9��M�]���'M��4Q@V"O�4:�ᏤEڱ��aA#�� "Ol�����G(��3�Ǘu�@��"O�t��o�<i"A�/�"�$��3"O�]��/˛J���I�iY�g�V�Q�"O䉐�[5>h ��ƙ4f�<�hU"O�	6G�zv"Q���R�}����4"OH	�dT�Vp�҃ҍDC��IT"O��N��``@y���&�� S�"O�%�ס��2�p�+r������"O���u Y�XP��\~!�"OD�35�M��M�0K�|p5#"O�m�΁�F��$B�I��G���7"O�����G<05RlQ�.۝�\Y�"O���Wl.�T|;���91�ڐZ�"O��(�/A���d-��j�"O��I4΅`��m��l�-��5Sr"Ov��C�#�X=j��`˶"Ob�k�ԏ	��-k�����A@�"OT�&#�1s�8��O�������"O��A�m,�����''��y)�"O ��W ZVl İ�.�P���b"O��)& >�j��c�&;�D�R"O�QY���;���K"!մ��t"Ol�	Ջ�	2O�@��۴C�<�Z%"O�@�a!Ϩ8��h�H��t��Ih�"O^����G~�\��)P����d"O�l�U ����I+�$��"O4�"��  И�	B�T��\uP"O�0����&>4T��h\�P�j%B"O\TpF�_	Yj�����x�3�P�<a]6,�.��ŋY�=k�Xx�ORO�<9���E8�Z�bڞv$0�
��<�D̀#ϚL+�Ci�pP�T�Jx�<�D`�&h�\���\9J2<$�t�<�5G^�E$�չ��1
�9�d�T�<�Q��X)z�QB�J�2���(�k�<�q�H�p�͋l6lI�gcf�<!`F�`�@����n�|���^_�<�m��-d�n�?W�h�a�G�<YbnM�	5@ ��%L�DN�8
�+E�<�2L�v�� ����<��t��C�<� �Ļ�lD�0�0�%�X0V{0"O�m:$#Աq�<i�$T�<\)�w"O��1FۮD�@`�a����@�%"OB1��&/V�Kኟ8j��QR"O��%�Ś�VI�E
=��C�"O|�B�mԛF�� cҽXЀ(0�"O^����N�)B1����hbݱ�"O@H�j�&z�l���LQp���"ON�jC��� :,�,�n�)S�"O\\8a�ŵ�hM"+�]?bhɖ"O���6K�K- U��
MԆu��"O`��29����"),q����"O���A�ղP���
��;���V"O.�-�8Θ�#��#�z� �"O&��$.i���� &4x@��v"O�(��A�Z��b(�&a��g"O�y�c��4)�TAj#���(��"O�(6J��r� p����R��"Of�#U��(� e����%��z�"O����h�so�p�f+.���rD"O~ͺv�1E����4��){< �"O�As���75�"��&��}v�9Y�"O���bŐ�f�j�2�\�bqv�'"O|��Lݡ]Tz �G ���̶hN!�DƄ@T��5-�.����C�( A!�d-��1s�J"ko ��,=��D�����f-R4|,`�0�����p�ȓyY��!fޟ3���A�+��q-(��ȓ$�E)� �]#@�����%۠܅ȓWtD	 #`�,Z�iI�!vmn�ȓQ��T�1e!wT��03hۚOZ���v��jpI>6X�U %).~�l<�ȓ+^bq�׊A:,ʸ���hhEUC�"O�����C}fΘ��Cl�aȵ"Oj ��	&q��ӇA�����1s"O�CL798 uǅ�*��m��"O�![���>���FI�G���P&"O,|yr�/I]n��4l�3��U�6"O�D;�K�dyP�@L��zE"O�	#T�^�_$����ذ{���3�"O�p�K�22��ӕȄ���)�"O5�GS 0IǊ7HP���"OpP��MT�?�ze �&��	�|=1T"O(�R��!&&��c���+H��1�"OD]Q�˟� ����E��>+u���"O���QMr�g�Јo\f|#�"O���Ug�H��Ss�[�ف"O�d�!��b&�0q��yH
��"O�1�6��D��C�g�\-��z"OB<�Q�Y�h{T�Y�ր��j�"OPx.Ľ9���˒9� E��"O��B�GVu���T�(��+p"O�P��L�&F���ق��{|=��"O<�ق�N���z�OQx`\�"�"Ol-�A.M�b�6����)EL��"O�"cNɋ8����� !'"�x��"O����Bҍ"8��hg	�.���*@"O�LÔ+�9D+N�2�(
�yA��#"O.�9GD � gHXR�ʂP(@<�6"Oh��GE�Nj�� g϶6<x�A"O����8���q�05Z�&"Oڝ{ �/���tlTN/�7+D���4eM�U� �CF�KU��x�%D�$��˖���U�R�=�bM��O%D�� �h��k�%6�X�rHC�dpy�A"Of ˂�9/Դ-"��ٱL4PA�"O�q��)٫qrd"�������"OFȆO]�y��qӡڱj�z`� "O�u�ބ�6�{��N$g����"O&\�%�7�� O����]��"O�@ �O��w�رB��K�h��"O�(R�)��0�2��|!���"O>�&kĮ�^l����qN`["Of�� �^mY�(��kOb>���"O�"5#W,rt<}����˖2���"O�4*ËM�B&�̪ kT����Sp"O�'�� .F*12PK�<|ɲ��"O�qv�C�*-�����O�^�6"O�`ۅF�/�U��㝜f~��!"O�������ia�c�7	�	If"Ox�Z���9-�H��01�<Ԓd"O����%�8zG��� AH�3S�i�"O��2�I	3�>h�@��36�	��"O��$��+��ձ��Ϯ -�D�t"O�l{�EZ�0����TM�'8�T�!F"O��IPN��p�ɪ!��,v����"OT�be�534�D�4�[z$�/D��{�a�zͫ.�/�N��F-8�y�oC :�����������"C��y�cِX��!J�Gҽ.�2u��H
�y�A.fvX�r�� [|�p� ���y2댁��chњQ�
��W�y�F\�K��!��iF�J��0�$#ٵ�yB�Y=fk
�s���:<�xJTb2�yeԷ^�|��EC�R�c��4�y�o�F�y��߻z�N�
���!�yB �#|zL�#��0*d�$��GP��yE��x{ M��^�t�y��C�y��""Kp�P'j�(vT,�A`A��y�H�"U��וK2�Z�-� �yb�^���zrbV��1����yBl��t&T`����� iA@,9�y�oM�eѤ� ��L2*vm˷cH�yr��@An���A T�	�N��y�*MP(�����:�$��%��yBn��F�(�HHA�/���pU� ��OJ�~"��rx�
�dܻBL�$.�
��ȓrtZD" �j��1���+0��(�'|ў"}j��\�
d��T%�H��0c�h�<���!i�D�K`��47 �rNQi�<���mFF,i��5VL:�/Fe�<iE�A�z���j׏G*�L���c�<Q䌓�^,��
F�A�Av�����Hb�<	vnhVn�� ��	�*��0cU�'��?��w�L�1E0
��W#Ȱ���<D��k��/S�]Z�A��/����e9D�lӀ*J&[�n082�ӞB�n�E.8D� *6!l�La���'����G1?��{�z,���$������Z|U4؅�I~ybM��I�N�
�BK�I�x�jGL��y��Q<��})�A��#u":�yRJɺĦ���N;cUR��f�5�y���t�R�
1�V[�TH8F��y�bMPD��.*Nb�m��HC�yb��Lw�qCf��I$��͖�y�%I�*���p�X<�����CҴ�yr�U%D�����.�ܥ��ݤ��<Y���ڰMX�����[	M����+L1!�� ���+B�8�9V#�&q]X�p�"O`�#E;~`�LA�b�	'E䜋w"Ou�ġ� "� )a@�}�
 ��O��=E����$Kx����c	��1�
D�y�e,r�dk! W|$Q��(]>�yBd �O���N�mZ$*�m\�kz:�r7"O��RK�?v�)����+m|�!"O�pS���c�R �5$Ife�l2���H�O����#��7�Rm�μ)n.�P�'j@����|r�t�A�#�ԍ�ʓ-́���M��y{��W'��ED{b�'|��(I"0Z\�+G'Hu����&O��AJ��ZYJ��S�]��8 W"Oj��xPqYE+C�ZoRRf�'�azR�|�͜>mN��R�L�3J��9�S���y扭XđB�) :>�$�0D	ԣ�y���p��)ñLX, $aX�b�y��=]�(5a_q�`La5�ў"~Γo��UpG��Pp��ȶ �)"��1�>AۓG���0�\�;�U˒lR�f�~�����Q���$�
��Q#.��E%D�0�l�� MHdr i%�ȉ'�(ʓX����'$�|*��m������#����I]N�<�s�F�nǎ9�S%%w�$����	;:6�?�)�矼Z�jN�8��a�6�Q�'�(���L"�$"�O�l
�,�2hVl��C�G-]T%a�O�A{��'�) fc�Wz�!C"P���x�'�~p�^�-��Q��O21�L\�������O�=�Ozt���h
��T��$�#;�t��'`���+rYR�j!��$�$���'h֜k���
�@��e�h㓵�31xɁ`lG������F��*D���m�!b� ����!6*� ڔ�)\O�b��ՏVU�t[P��gn�MA�#)D�����G�9��JDb��B���i�g2�I~���'F�~h��#�Y�V�@��/��H�ȓ+{ ���@E�ݔ-)@��,jO�!�ȓ �90��� MS>����/䮀�ȓ`��%�Eb-	�9P�/�8+P�EGy���M �j9]�n�)#�N9i�(h��"O�x'��5��|C�ňrd6�`"O��[E��g�, bwB@8<FX91"O0L �фx�ȩR��>|/6��gO:�$�',����d	ܩLK�H�  �9!x!�D�%*#�И�ϑKIh]iᎌ�{�axB��:fr�`�U3$6�	��G�WVC�I=Tw�!���5Le���<i�T���'Q?��O���B���ϛ�e.�RGk4D�в��ǰx��5ąY�^,�U�apӮ�=E�ܴ7�rE�v�Z�Rt	X\z�E��D�Np��"p<̊Ga��b,����s��3ѪF��b�!өy���ZG&9�eP��哗ln*9)E�¾s�ָ)6A�$>�	2��?)���:�40������*�OyBFȗ�O�IҔ��]�%�׏޴F j�ra̕���ȓ��SCi^�P�883�Ƭ6ln�c~��'{J#���pvhH@�#I��ۓ��'�\woԼ4d�q���<���S�O0�=E�d$�X��<U _�j�t�0��"�y2C�Ĵ��*�.]I��Ap�?��3�O�u���+���G�B��\�6�Ipx� a5��c��Y����,�i��A,D�T�CI.l�A��8�d�(��Hh<�6�?l&�)Q	U�YH��4��N�<� �"O�?|�����X	��ܓS�i1ў"~n�6U�l�g2��)�0�N<R�rC�I�c<��I��W�-g�(���5��C�1�"�it��.i�F���Ҳ]�HC��m��(!rF
#��a�A��8q�C�I"A���B��3IZ ��tl��t�B�	5J:Бf%L ��Y�ciM%��B�	�:OD�I>��i�eK�i�B�� 8i"�`�Q�A���"ٟ[-:��$�S�OK�<Q�l���ŭWU6��t�(�yB�X}`"]�ք(%��u;#Kߤ���=�O�hC�� �N��͕ld� �'X�	�6�4Ijgу?�0����	�H�z�=��~������z�`X����1L\E~���< (�QZ��D�}�Yc��E�LJC�B��h�f��ww�tpD��*�p#=��O"}�uk
6�j�R�#��I�(T�tH�G�?�B��C�L���<�y�2�=E�ܴ�
���"n��p��!+���%��x�L�*ilz��g�;�����*e�9C+[�/��X����1�f\����E��FHl���Q��wOP���d����G�����c�n�GA�\��4Dt��J��`69�$��b䄇�$=>hR��H�D��2B��=D7mGxB�)�dKǷy@n���N�v�<�f�M�<�-ǏzB�A��Oee�[SQ$ո'���x�f��@׉͜\�jŇ,�y�O80E�|8$�O]~�ĈG�y��ڒ#��9H���8>��������0=�2l�2'v��#��.��ä�4�y�n�/��.4�Բ��S��y����V��К'ퟯ3Rxi�2/$�y��Ą����C��/��t�q�G*���*�OUSS	!��y�Wf�?6����"Ot���ᏂX�bI�q$�$�Z�%"O��P
��]GH ���I�N�����'֑��Z2�C#4�gg�(�9a�&D����ܱf�ňGV !8v�a� }��)�S&\:N� $��A%L1�"�S-Q��C�I4$r�y��&J�6���ݭ/��'A(O`��f��`��"��Rw���Ol� G&ڑ2�4�jE�G.ق��Ԍ`!�"0���֭�n� �HbG�4J���XEI3,O�I@ŉ'�*���b������J̈́��k�'8H�d�gk�0�@N׷Z��	�'��	d��1;k�� ѩǳo�}�'� �2��	�3���اn�:�S�'3صA��D~���ïk���r�'z�9#J�q�9���". ��9�'�����(8a*E
׊P� ��Z�'V�u�k˚7p�$���� ��'� �闡�G���`Z��X��
�'b�1�f�rdH�u�>G:�
�'CDDB!C�/>��UI�l�}��'F����Λa��}S�A:x���'v$h:B��gx|���n�,|�	�'�Ҥ��E�7��	[Rh�>-BiR	�'����n�W;�yٱ ��u[�'34E�D�W8�:�F�yS��
�'�x�P��Y����c����)�'�L��MA;9�ȕ�*�	kVp|��':8����6�4�"V#�	o�x���'���r���8	*�9K5=q`^q���� ����H>��p���7C�,��0"O`�y�lF�p���ڳk���R��G"O���I�3)�$ �)�'q��� `"O:���Y�-.������Y��D0�"O�m"3$S�8X��ɛ�"z���"O����#@{� ���R
J\N�c"O�A{���"f^%�TN���Q"Ov���S]B��IK6y*<K""O��c��[�t��k�eK�
 ��f"ObH²�C-z��9�o�Z����"O�
T����+��@�i�"OP9��.Ʉ3�(�R$C"l2�B�"O���nçFL�X[&Q5L�e��"OX=k!B�h���A�EXn�B��'�V�5
��	�������k�-&ڬB�'��XG%B*�^M��o� 0�1�'� ��4�y=X���t5����'��ܢ��N�0M�c��k,���
�'�DЊ��	Z�x��L
?d���'�"��oF���Eೠ�d����'0�@�H�+��a�BX����'�N����] L�Ȓ�o�6�C�'�r�Q�J��+_"�U�=O)��[
�'��I�mȮ~�R���`�>E.x�H
�'e�Y�R�^2$w�Y3D�<L��-��'��}񴀇?����	F��`P��%��'~�
 ����h�T`nH-�y���.hjV	qs��'s� ��9�yG�M�x�yG��h�)��y�?� uk�����p���?�yR�23FPxq��,y��A��A��y�E�V
��[4A58M�X��B��y���\�L���L�2�5 4$_�yB���Q#�\'�Ւ!T�@9ģ��y����uj�HC�x U�$C���y�OB�qd%{�K�[L2!�F�#�y2�XN��$X'S�zXӆ�@��yrgߠ	J�)�!ԶO-�P[�����y���'zX���h�0��yY�ꐉ�yb��=�&Y��Ǆ�(���:$
��y�	���H)�E 5�,�C4M��y2��^1�黖I%fͮ$��"�7�y�g��V�R%�K�^yd5 �k*�y2b� XӸM{_�|XBNE��y�I��=��J
����]��y���*��bG���LFeS/���y�C���.aa��J`��SRf«�yRI�� �\�r��D���Aq+��y�'�X�	��D[y�=���Y
�yR�%������h��ISߒ�y�i�$�j�-F���X�Q���y�R&L� �di��]��K��;�y2'u��rg�F�L��yb�yB�̠����A`�=��R*�y�-� -��rbb�9Ty^D��+�y�Hx�&��Lc�ܡ�D��y���Gd\�sBaE�JݾDc�L��y�ֳ.�@4�Ǒ�N�0p�Ĭ�$�yß����XC�BFhxC�c���yª�	�r��ŇN>"칹Cb�y@ڜJ@�7�Ό'Z|�Î���yB���5�vƁ�.�k��P�y����4Y����:�C�9�y�f *OD8T;'S	pu�+����y
� 1��#��2�y˖M�#J��@Y�"O�MZE��22��*Y�����"ON�����+n���BL�"u2h��"O|�R��`>�=�6�*$��"O6i׺y=��B�;�(� "O��T��54��d�W�����Rb"O2Ĳ��Yj�+v���9�|�z�"Oִ�$̖9�P��(�<�P[b"O���m�wm��;�F�~5�"OL�R
\�1_����KSu�j�D"O��y�DX�^����)W�+ǘ��"O���ц��|<y�S��i�|���"O�|G�ݛ���/*�.�	d"O��bV�i~<�b&�f%�S"O�cׯ�!o�� �Al_�ԡ""O��B���3[�qp`T5|7�!��"O��a�$N�y���ȋ�HEZ�"O��i  �+,p����T���Y�"O9�m�M	
y���-	u��"O��y���6u��Q���}���Y��'�~ zs��_�S�O�\��,ؘ1�|�Z��.R��"O�A{���"R�ɲ�A�,4xifZ�����ּ�`��	?f݃� �>j����!�� H��z�Ϛ<c=j�T�ҧhy ����
�xіP�W�F�}�x�B��K�<f�U�a��tB��J��dpj#�C��ldBs�Z�eN�X�j�g�O�,�c�	��)0��S�E����'(���ܵb_�X�Ri��Y!`A��L��eCV%���?�f��*��\5��>�c��?fj��R*-5(X�t��~��9U"�
�Y�'���Jm� y�<[�:�T�3,��P��$�WA�0r�ĵ!�'����D�k�LDb��&@. 0zN>i���C)(R�ȫ�Tb8"�$"� аCXt��h� Ho�,µ��pӦPp&�i�<��阨, �iC'�4����t��]zF��A?����,0�Ȩk��R3TQ(+��0CNq�ej��I%e�ˑ�2�����;4�0I�I��f�ǟ?��y���2 ���iq��1w�����xc�	��r�+#ן�+Px,ԁ��5K�Y���I'C�a��	97L�i�c���%A�$�,<,A��Oϑ@b^		�,�%ZJ��B����!tF��q��zr+Պ&�Tx
Q��U3�Ka;��T6 �+��L<!�V�	�C]H����	i����i�\)$L�������;,�	`�'�RA��nR$u��sG�$O�  Vn6^�"�;�(8q� 2��OK���<����ϺMx����˷S40��4O�IX1jϪJ��d��B��[D$�����TK���D��U\���$��^�l܂ ���%#�w{*��D��h|~Ѳ���<	A�I��H �ϝ�I
E��ϔo�<I��V�� ���Ŋ	�(�����fܓc��qh�,�:�ȟv�#�h]�oLj��q/��'��"O�T�2N�$d��a�9#�A�$+�<	I>�a�>��	7#��q�# ���0l�©�q�<�6.��[�����
�Fp����l��E�ką��	@�ŃTn�E��Q���jAN��8k�P|!0nZ��ybI]K��Hx�m	]����W�*�y"� ���V`8��#��@�ܸ'���+��yيQ�'�lcLc3�߿|�	cuJT��Ҵ�ȓw#����IF�;Z}���O�Pl� *�b��=�nܤOܸy��Y�TB�&N�{2���$�0r(�{�F2D��z� CDH��4���A�
&i,f:�0D!�H�
�'�|�A�j�'�h����W�k�hh1��z
L�9
�[V��#� d��I?.�$����t}sދ���	��0sq�W���;W�[�Gl+bɒ�A����t�*Y��yŜ�#���%T�n���)�q��N� |�<���^�q���_<sG!�DM�d$.m{c��'�b�y���/=�cbR6���\1j�YLd�1�r�̻.pi�d˕'�4l�%Ϝ=��A�ȓ-J$�haA4!_��z�oO7k#����C��U+>���/(���+���/��i��O;ONur��g�`C�I�$hz�bK��U�h�Aڜ��Ǐ(�L�(q����=� BL �(�@�Vm��6-���'��}@��!(8HDo�Q� ;󨙦7\!j�!@�#-C�I�C�lj�k�g�&%kЉ�'A��x��$��W�r���S��¼BT`��`v1#D�
��#<I�P�ڣ~Rs�^�T���+�w��<k��+4���^�d��M��F��'�ب�0f] ̾�;4D�8[�P��a͋	f�]H>����O��	W�٬
<\z�F�6�&���Y�6HZ�f"|O�@؁��*��"�e)��(��i:�k�B�Y��(G|R��??�b��D(x!I�Í-LB.8A�W"؄�I%nP�z�����4�:P�f�)
mX<ꁆ��y"۽]�hh�a@��r�HAAŅ��'$XL �a�i�@|E���״}��d��&M{_�b�h��y2H5	j��J��t�z�"lGx�d�`��,&y���>�;ܞ�cѬ1 �Y+��3�P��_�����a܌0#-�zX�n��|��Ș��Z�d�{&̘Vd���Ύ+_���ĬV�=a��!Q����2m�O�x�J�d�AI�U��� "O�X��G4�
��ȧ}r4�W��G���E�?�h�
<yR�ޔ?�!��
hW$�v"O"9�S��  芔���aj�!X��?�n,0��(}� =�g}\"z4�4BЉB�h�(V��yB_��@�V,G�m�H�wG��M�ӫ��KՄ�`�M5|O�)wCD |�J-�qiD�}��l�'�'�B$��ϧ|���ߝ4�=��e��܍P�J��!�$\V�X�j�h�15y�iR4)�z7� �c�Ƹ#�Q?)i��,]0E���NU�<ɪ��8D����I���B�Ua��3h����0ғ�RP��m9�'l�XBfL�k���CH��Q�؅�}nt��aȌw��3�ƙ�b���W���{��hg� }��9Or�x�SY�$�z�]�pD��#�"O:�����<`&J�y�CUh"8�3��i2���Gl2+~��!mDGx�"d��_�$؃�C��5�*PP*(\O��H��M=	Z�"rP)[PV� ���*P00#�t�,�$E%$�d%�0ffx 4�*��aq�=�I�U�xSn�*%.��s�C`�eCh)cU�{nh�bJ;0�)�ȓh�Ҕ���͇x�Ґ��"��Gz)�nL�h�\�g�)Ps��s���$�� ��z���Wx%I1j�9�!��/�f�/�T��%(X� �dђ��,ܞ��QO�
Z��IǓ,"nX�C���:����A۱n����ɡ;��ڲh�����ks��R��K �K�/O.6��$��l<�A�B�L�����]($�겭[�I<\,.Ū"���6(��O)����|"��S�AܐA�Nɻu'����!�S�<Y��]W:!2��*J����4IV�a��e� �&d>���m��L�n����O��b$@� 8%�H�7I7Y`�8�O����X=nI���QB��y��;M?��ec�L��p��L�T����$Pw��iÒC9.�ѰR�Tq�y�hC�;)���D՝}uG*�5�52�o�(���4�;y�@+qO��*��0��xyw�-%�����|b���#���FmJ��h y�OOu�1��=B&�=CKTT�%�	�)y���#"O�ة��7TѲ��$JS�5��N��P��E.m&�T����IG���H�X�e�G�ZTXE��W|���#NXb0bN/3�=0�bX�^�H� �� $��b�@� ���%�M�HI�
��#4ހ�P ! LO�B�@�H�)����)KE� �ET874r������)�PTh�"M�p]!��V i���j ۻ1�f�cB.Q /qO�=׈��U����k�ډ�}��"J5-|}��-�ALZ�aʖA�<�e�"*]��GJ$��A0��_҂4��Q�y��Q��'�%D�,O��K[� ����J�{�ޅ��"OT|�ѯ��`�` b�'}��@�i:�}8���L��d��ux��뤍։|�N}ZF�E�OЪ���=�Ou�f%�4��}�FKZ�&�p����Ԓ�@-[�!�d��{���Y���Ъ&)f�C���^2A3��z��)�@i,)� �
3CD YB#7�!�/��-ѓ��{�6�9�Ȅ)g�!�� �Ԉ���u3z����[x���"ON܈�[��L2���;Y�P1�"Ob�	� ���	)�%*L���"OD]c@lӚ������Wh8��"O��+�"�fk���jY�H�!"O�]�a�P;D��$�۠b\���'"O�u�Q�		�x��g%;�8ã"O,�g�� Z�q�f1uB((3C"O逗l�5�"�@e;q=���"O��$g�J,4a+v�9���"O �z�
$�t�ւڐfŜ5�"O� h`:f��D�D�QYШ�!"O�U����V�\D���1-G����'� L3�R�_H<)H�T�B�&a��'�ݚG�7`�T(�.�?�VL�
�'�����RJ�{FNIF���	�'@�D�J%Vj�e5�:�	�'Qp\YC)ϭ*TMӅ��&�N�*�'����HK;^�ހX˻H�"���'�t5�C��RWa:Ձ��6D���EI�)��T�P�X�]��%/2D�h��'Y�A���&�y�xHRÉ3D��#�)I�;xr\���
,�e�$D�TKФN X�l�P��Y$g��h�s-"D�D8�D^,^�P�f�T�˔�s�c<D�4qB�/	��Ʌ��X�F�PO!D���f��D�h ��ic�$���i?D�*	S�ZY32���xTdj�k=D�08�H��	���KѸv8�m�!L:D�|�'"0E D�V��og�����9D���U�U�4<�S@��+1�`�yq9D��Qt
��
�����΋�\���a�:D����5h
r��DiGd	?/o�}�	�'�nx1C璇fQ�8��˃� �}2	�'d�vLG:�fx�F���T*��A�':�(hM9PRİ&lF�X<`���'��U3r��B�zu��Oӧb-���'$@3� ���� P�gm�U��'��;���5�@���O��PL�T��'���P��+Cx�b�^�I��Q��'�"\���e��d��ѹ}��%r�'�H� ��8u@��Ҫ��D}Ą�'���A��~)�H!�,T�6 �p	�'� ���5^-�Is�C>-�����'����uhR�.�TQ�φ�I�Hdj�'1J��V��"TE��]Me#
�'�z�2�g=���`��J�c
�'��@Hdf~�5�V��kJ�<@��;D� 	d�������5Jݶ:B�P�v�2D� �D��O��8���3�`���d.D�dr�@4��с��ݯ�l�3 3D��B���!��)R�[]r �3��1D�� Ph�/MC&�E�X9R���"/D�غFM�i�~<�U��a���#�*D�h�e )2FF�s�$)Y�dXq�-D�<��*=25(U�@��iŪ���+D�Ps�&�L�)w��G~� )@�&D��k�)]2U�� W����`���K9D�D�$ꀁA��	ʄ才z�+�:D��[�HUH�����I�\���v%4D�ܸ0��ee�d�T��,a���'D�ty�"�-!f j��6�F0�U�%D��A����Tb"JR-��ۄ�$D��R��F�g%�Jt���+?�u*��%D��  (�#�����;���.�>�*�"O�Y��DM�?�`у�B_�^�% "O�x��֡?e�K� 4XPe��"O�zw� 2p�8�MA5)Ry�"O�y)f�ȵd�8�j�J.[,>4(&"O�9�c�)8ƺ�)#J�=�`}I�"O��J�škF����=q֠��"O�0�bmC�F|x��V㗜2q�"Onu���2+>� !�#�58Gb9�$"O�,�j��"(��I⩅�O2	�$"O	��
$A�P0�f�
N3��8�"O��6�\�C	Nx(�י��}�"O� ��_624�`���d�<BA"Oؽk�憊Q���#��3v4�Z�"O��(u���b�Tl�S�K"jɾԸP"O�� �֎Q�h�	�+�%,���"O8-���W� 	�� ��.`�8�%"O��hi_.�LB�IUH��`+�"Ol*S+Ǥ`}D-� ��
h����"O��2�Ŕ'���`2gU�T�J]��"O~��&GB�jK�E�U&BW����"O@�A�Lq��da��2Ȃ��6"O��P��D�T��%�t�E"W�HI:t"O� ��@��B��$�Q����A�'
����k~�S�O�t�Z�_�Fթ��u�0�u"O�� ���>+�%�U�!b|�`V��IQ��-X�e��I3�L1a��T��Z�A��=���ƨWcI���χ!�(:���A��i�%B\ikp
��Py#A:s���Ї�mN$	e�H̓oF0!5� �v;�s��_}�O��T��F�`�j�J�BOg����'�āu'�%#�$l���[�n�@9�kA�Z^eZ�����?���"�̑UgT���>�"���>�v	[�^* @0�F'MS�����U�"��u�'(�й�H�ml`�*ϲ,ǂq��D��o��a�f�G���0�R�' l�C��3�P-�$�O7��|AI>�ϗ4��di!⦟���*@'q����f
	1��Ѷ��u �؆BQ,��))��l�<���z�~
��\���4���x�\i�g�O� �d�:��[��B?I;˧'�Z���w��D���H3�M�7bڗ,&>���'�ȩ��,U�J��a�灊�y7`=�5�](�F��D��'|R�"^�µ��T�O�i�g�dF�!Z0�kU@�	9��aآ�0=9��Yo���`,��`a �Y2�y�!h��4��X1e�$.����&���j�+\O��c����/��Ā0h�9`9��|�Ϻ<x	�g	Kx?�G��B|��A ���I_�7���,2^�q^���q��a+�`��''�-s1%\�]�:�rfNؚY(�j���0W��s���JQ�U��O�X�Cu6��A�č�\I�qZŊ�\D�P�'O�����3D��QMӛdUH���cA�_9L%{�N���$�z�8������¸Z,����I��Ɂ�az��N�̴��T���b�^�l��uh�ȓ�.S>!��:D� p%(�=/*��3 nO"���y�M<�I�n���N�k�O��F�\o&��� Q�q�R��'��y��/]a�b��1|c�Y��٦	�֕%�\���Y�j�.��zNZDB٨]�!h/D����!�F���R&L
�̀�˗#�=ȸQ$�ɪg�����=M:oH�4�t��z�FF�G�����<�����e��b�/t_�\P�{�<�GފhZg
$u%�b�,�uܓ�3VE�>�R"~�� � S��E��i������O�s�<��j��X%恓��`���X.�.z��y�%x�D+�(��m�N����4;��ك�ny(XC�	+~ʬ�ZFʙWž��a��2]�̰��l
�b���A�;}��Y]��qEx��=v5����^�K����g�p=��%R6;���iF~��a�?s�i�K�5q����{��#W��~� X��	bM$�S0��y`L���Æv���L�ѡ�:Z^l{2Y��*sM��jq�Q���.U���� �W�j ��R�"OV��5M��m`��dˈ&�h�y�U�_�\@��O6&r�'�z�1�\��{�? �@�#�����A� ,��"O���&Δ�%�l����["}K��[*k�P1�*�[�d�Ƒ�����'��:D��dv>1kB�I37���'��e��۷|~�)`�ɩc
�Y��\�U�0g�Ӝ���#D�R�QMȅ5Ԙ��Y�y��{b-�l����-��5�P�Z5���r/E).F� r2�9D���1�)0�狉|�������O�(�T�՞@kC��i/�(X��ݗ ����F*���c�S,-	Q?-yt�T�x��5ԍ�߰���COE!B	���3���^��~R��C{pm�bdֱ _���­� '6D�W����h���<@SŢ �ΟD��!y���E����,���iD�8|Of2s�`X Ӿ p-!G�ig�Ұ���eF|���]I�Uϓ6*�q��+��l�D#�JB�zJ�-��	�b�Ha��O��go.�e3F8
q�ͻe)���ϓ�y���(D�ST���7�"qXp&���اE�o)��E�(ڧ!��q��1ra
9���$Oɂa�ȓ7D�৭�0�TzE$ØL���@#�Ux��D�I����Y����D:��x� PS�ջ��&D�T�u��g�l���$-(����*`ӊDA�cM�k;�U�ߓz�R|���Ѡ^�����������퉐p����!T>S������dŢtDbl0�a��y���G�b����͞n�65XB)�9��'�L����C��G��o�_��1Ӯ��6A��0fg�P�<�S働s�e`��o� U��J�>]*�8�'X�􉕦H��	�)g�D�v�	�֭�fM`�C�I�W���d�`¸����)��7MW8a����b�7��=���D���Q8#s��K���N���#r;f�j��-ft�r��^HVpcC�4/��!��<ff���i�4��tC�O@�\�qFx��2Oz��F�T.�16�K��l|� A�>[&��ȓ<+T<��f��W�zTژD[����K�Fz�Ӈx���B�n3����Q��W2T9NdBA厢Z��Ői�t!�=E��Lx$br͍�`���Iӥ/�*q��^O��@��Z3�$�A3h��'�(̓T�![�ҙ��=A��έQAB�1�$�3\f9R�� T��<3��V�&� TQ��i��qC�җUm�9�E��3U���
�'����Ōۊ@eƭ�U +r;|!�b�.@H���w�O���c�&��Y1�M��x+�'jX�{�H>V���8�k"Ά�Q�f��q�,�[��,}��p��"h�*�(��R2j���&%:D�trB�<=�p1�$�	1h�����OP��s��G� ۓk{rD@�[#-[��r�޶9R���I.0�]��ōiyvLص�ƍ�A�aLb~��ꥫǏ\:!�ԑ"����W�F1B$X�{q��N�OJ�T���&M@i[e�c�q�,buBΦn��0a�>�X�r"O�̻d,��rq^�����3��v'��H���G'�.x�h ��'v�>���I���#{i���o̘\�.C�	"r�����Ň��,�r�X&R�J��?H�Vh��/Ȁ,=�E��4O,�K���`�A� �@+bB�m;��'���M*N�
 I1.S�[]$p�4�CC���뵈��8}��~�}!dE[;
�;%��5SF��D}B�GZ�����@z�'3��́��I�eT�|�*�`!�5�ȓ{h��ӧ�c�@���G��Y��0�,J�0kƢL�<o@ӧh�*��шY�m�t�`��H8�h�rG"ON`ɓ+�
6�D�:��sa���SXU��f�":���1�x�W�q�:i�egƃ~��~����$�0(�F�9b�P��hI�Ew͒u��Aj����n�A�DNI��~Q���$5��G~O��pO�����	52*B��TE�QZ�h��!�Ѿavv)���|Ozؚ��&U�	 �5�q��S(��xA$�
K]f�ʥ��8�&C�	�`�4�����H�+� �C��	`{ƌ��b��(�><$C�)� �L�cE��\ kVL�b.��jE"O���Fl>���s�Z5V�b�"O\�jdl�75 d�#$DQ��\��"Ode�ҍJ?�9��t.`�R5"Ox(�����)��h�<
`Պ�"O�j�!�T$}Xg�L#��I�"O�eh�e�q�
�QE�F�qR�"O ��B	�(��)=�L�Ja��BN!��:�����$�v�(A���!�$��uGԉ�! ԨJ�dEIjGA�!�D@�h�e D�F����q��3�!�°
��: �&���6E�12!���F�����̏}x�=��GL�R-!����Ś�+�}o��9$�̬7!���vhp9c�M�mO�5
F�ٿ^�!�� Ͳ�{`�	�D<m�b��d!򤇕thh xE�єeNЅ{�* �r!��H�r��ń~���d¥J�!��^e.n��R/���Sa�L�c�!��I� #)!x�4tSE�C�!�>r�1CTK嬀���D�mL!�V���{�%1%Τ�p�NX�u>a~�lU9�ތ�K޸|��t����&A�t��&����g�)�7-Ԯ|�&Y�)��>���� ���5& l ��8�(��c*��ʭQs"���B|>-qЏM�	��]�����Z�)������� ��5�?�2[���i���N�qmZ�O9�|爃�פ�����M#�	�O���O�|�*�ҙ\Mj�����C���f��*r��'���N|�����)�BE�l�p9�����c̸�~��O��,�|�#��;�	W&�ዏKڎ����̢����#G��Y�S��gߪ�"�E;� 8�'���V�~���.@��~�Ӻ�?���ˮZ,�IT38�^��E�p�<YG"�#9|zt���W6��h�E��Z$ɂ�8q�6 R-*q�����4E�t9��B����[i�v�zdeG��)���-���/r޸�:��o+B�_�uQeū��S�Oz`�F���	�dp �;Q�&p��'��ݐ�oF�2�ɧ������_�C��вE��-�0��` �Hl��3D�-��~�%������$Sc�l���Q���O�x�t�Pa��V�`�T!t�9P�\X
C�6���܋r�R���J�la�T!*�9z!J�w����B�H�y�n�#���r�m.?)T�9�p�peAf9�@]+���*��GQ �A֣�ҡ��A!�h\{I	w������D�:z7��5G�F�xg.�9zRdCd�!w�a�D&؉�F!�Ă7�������]e��I�I.|���ʌn�z��ç��d��#u��H��k�15����K��e�\���-O�>�Sႍl*v��H��`�fY�����:,���BG?=��.O�?q�i���$
���J.Lur��O��$lr!i ���]��0|�R�:�x��0�k��J,�r��,:��I�u�V0Å�O#2�ڔ,�%��@2w�\;�A"�<�霑s`�x@&)����b���=�&C1����$"OVŒ�bܾc52%�󌙣`ü�{f"O8��qe����19¬�obz���"OdX�DD�d�B�(�%�+Sx��T"O��4bބ�ST��FH ta"OR�04Ƙ>5�RY9`�ƒ����"OhE�H�>[��Eq%��l@�ez�"O��!Q�!���E�1���"OD�6����(�b@�!��T"Or��#֊e1	E�;h�X+G"O��g�D6u��h �rIxc"O����%C���Ƌ�\U0�k�"O�1���-=t�d�`��
EZ Y�"O�<�`IO3�DE����N5@APW"OrSa�&,��M�U6!�m�"O���˒�R����T��7���kv"O���c�	J4�����L�"O� �쫔HW3X�.�+�@H����"O:���a�)Z�<	b�e(�]�U"O���d�[P��eP#�	[�I��"O� �mP�^��Q dg3���Ӈ"O�aI��@2�0�xS��< �j���"Oi{p%B�#e8�@���9<���T"ONP!�o�a,�k"D�'�I�"O��%��p���
R,���"OZyʤ���fm���B�2d�����"O���q"���_�0���Yv"O���5�U9j�\e&U�vh��"OJ���ϲ4t<pH֩e�B�A�"O���@�R:GnNE+ф�"�Ҙ
�"O�u���'M�}	�#�RP�S"O���ulJ0��%�R��g�>�x"O�Y�hJ�CB����BE6r,�ص"O ��c�x56tq��}2ܠ3�"O����h��p��L�v��|��9B�"OȜAb
O�|[8d�a)PP����"O��:�#�rR5;�A�Q����"O����>���6f_*CdM�`��<!$��7
�$b�,@�/�$�`�s�<��<P� $	��u�-i��E�<	�&�6EΉ���!BhȨ��YC�<�6�S36m|̳���1��L`��W�<��7kp
Axb&ٌG))p��~�<aTl϶k������lh���u��|�<)F ;�.�� IV���;���{�<ifM�n�:��M�R�Q�C��P�<��gO "�k@��-<H�j�m]J�<��L��v��3A�'&8�H{g�C�<�)�D�x����I=t)K�(�x�<A�/�:<�@� 3�
%t��tŀI�<RIJ+Z;8-��hʤZ|�	�q��|�<��eA�1H�<b�j&�Ba���
S�<�G�_�}�H$8RO�.��}:��O�<�&�	����bH�W����$MJ�<e���!���3.ЍJ��2S�H�<�� 		uܮ%#�eA,��G��<��C$�<��d�ܱFP��x�<-�@JQo�� ���ԅwA*���y���0�`ʅi��"G�3�P��P)��1B�4VX��I�ʜ
���� �f` ��@�T���	 ��}�� ��B"-�`�%%h�����NF�%���6�����U�R�;�B"](U��0�&��Dd�F�t!����F9�� �t�[BՓ~Q��`S�����ȓ<( 鋓	A���Y����4�E�ȓz��̈1ʉ6#����Qf�2�&q�ȓO�	:W��"}��a�MTn"}����]�S�Y)�������x�Jp��u|a��F_(���P��,9����r��H�r,�B@��{C+�<-��ܥ�Q�\t���&G+�ȓ3�Ҍ���\2w΍�Q��k%���]�ՋC�=��{�������{Ƥ�(�O��e�Vt��eΘd�*���~d��������$+p�ԇ�6)��ࠈ�-{ZvЁW`UZ�>��ȓSh�Ԃ��\$¬9��G�2i `�ȓ8�`�ʢ┤7�e�gޥ4�
��U:}���\���*67���B���E2S^�����5�z]��S�? �,S%�@�1b00� @\�w�8q��"O�t�R�A  �搳 N�<�C�"OZ���j�=a��x*��M�f�y�q"O\�p��Pin��qJ�P��p��"O佘b�D�ŀ`C ��e�"O�\!R �{ ��4$X:u-�@�"O�{rD{u"�X��\BY�"O. �u���a����VoИ<<�$"O�9#��K�"�-�@���#���y2 ��2�8TA��@p搝���y2C%uB!���l�4	�%� �y�L�l�y2C\-L���G5�y�˞_����To�J�C�oɗ�y�'I*j�F��6,�@@혿�y�F;�V����I;`J�17����yRh�e��B���6+p��&�y��~(���
ݥ~J������.�y"��y�j%�bD��{��5���y��1'�,���l��nu�	���ڎ�yڌeu�P"(&�!��D3a!��=\B8���.�#ܨ��;Qi!�D\+"`(�W$֘Ka�/Ʌ^!�DE}�)��D�@��)�m�	vK!���{Q��m\E�p��B�1�!���yU0���V�Vޠ0R���!�dǉv��1ku�U_ waăo�!�ʻ-8� �W�ՖUۺir`��u�!�Ė.{ �P��>o�`�Αd�!�7L.�aTF*q��Ha#.W&!�d�3N����o��*�8EN��I!��>uGހ9f�	�n��]�f$!�d%~���ـ��3��Dad���[!!�Ą�$�I���hn�݀wJ�<�!�D�w	2a[��C�7�<�BJM�s�!��&�$ P�Y�T� �� H</�!��6�(��\'>��h��
�t�!���ݮ��vOZ<>X�>D�iEm+�Lq�:��ᷪ;D�$���3l8�����_n� �A�5D��1O�s��≐!
��$�8D��ga]?W&�Q�⎴(m|h�F:D���e��/s�8�8�/�@���{w�8D�:���i ��0	�k�&*�BC��=��C��^c����g) _
C�I�81�dSC���!��9�+)#�B�Ɉ����e�	�=w0�0�A�g��C�	8/ �v�$b�L�[!�]�p�B�ɑu�t�ᤆ�4�Y1��3c(`C�	
�t�H'�_��.ǗI��C��v �i��I+D���J/�.�B��7B����K/3�-���-͐B䉅E�-�&SF��pㅨ����B��?s�Y[I\%bx�U��6B�I*1���:�C�?Ja$�3U�,�"B��'iʠ�Xs��"�8�Y�P�r�B�I�
��U8B�ֵh:��s���"*	�C��)ifjI" @��ԫ�/��P��C�I�/7���D�#^�{Ы�(RN�B䉚u�.<�*�!\g<�  B�i98C�:j@nHeF�_)|�)���B䉻F��	I��9�pԻ�	ڭO��B䉄N9�u8�"�?V`XPz�
�&_\B��;w`֎�jW���(��PV B�	�A���A��8x"&���%�@B�)� 99��H�e���{A� �� �"O\��R�W:BI�<�1/@42��q��"OU�uoI3�}�PmF�(��UB"Oİ@�*NX"��ࡉ
<�$�S"Oވ���
ga����%O�T���"O��B�ǟ9JD���J��C�6"�"O$| '�,�<'�^��@"Oιj����1{F�ǝ��e{"O�A�C�Ŀ>?��+`]�\����"O ��&�Z�P�aE��F�"O4���K9)�|l��F�%qw�$��"OF�S����D�	s Fp��c 3�!�$�!
twX�U����VBקA!�d�:2��`al[�V�ĩp���e�!��  ��q�Ƃ�\���֫K
�!�F. �����'(�d���F>p!�֡[z�*���=^�����Zh!��)S�J��&b�Hdމ��ڼ$[!�K��}�&��~�qS@/�S!��Y-y�<C��)Fm����E!��y�Ȑ�CT�S��ᶇh!��\�^Ay��Z)w3n�a&�?!�DÙ |�� �Nh���3��-y\!�dߘA�(���O�!�P4Zb�ӷA!�DC�P�Ñ�7�D9����?1!��Z4^2�� �.�B���m=@�!�>q <�2?qJ` �PJ�!�D�F�=�5�Y�.�P!c��n�!��Ŗֈ��4��0'�D�cV#�f�!�JQ�Oơ�6�k�B�n!�d��x/�,��#H�%�LɪԠjf!�DL�r���+��ۯ��3�̈Dt!�ā�n���觀ðh�@�*��M��!�dZ�jP�q����;-s.4�0��#5u!�d٫v�N�@�	xV��aQ� �mk!�$�3:���(W	�"9R�������~\!�dŏZ����gE�o/�)���.}�!�$N�3l�����%B-�y���7�!�ć�E��S�&�S�\p����$�!�PG��� `�ރL! ���i�4�!�ں��10��-8�u��D�!�����l6%�'
+B�B����!���;�x�`��5�l��U�Z|!�$^�F�$@���A�X��@R,�"u!��	_:�i�gܘL�-���W�|l!�$�mI:��$,=m��sIÌeT!�%o��ʵb�9��${�H�O!򄁹}V���nS�}��S��"�!�d��'�����J�ew�}���
�!���b��|�g ��/c�y�e�8b!�DQ%\S ��r"zMJ�ΐY�!򄙅\� �  ��     �  �  �  >+  �5  @  TJ  �R  I^  �g  %n  �t  {  X�  ��  ލ   �  b�  ��  �  &�  g�  ��  �  2�  u�  ��  r�  ��  ��  
�  M�  � i  � �! &( )  Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�� |d��"O
`�(�;���8���-0��1%"Oj4��ND^[��"3/9�0|H�"OB���H��*�ʞRy=a"O�味V�!X��!&F�:J�$���"O,��a
���C�Ą�M�"O,$3%o�-���p���+Ն�:1"O��ݢ1����`���y14]2��i�<�6��{_���c�H�`�fX�$Kn�<��A̼VI�xR[�)�Ć�pඤ�ȓA5��('nߡ4�� �)˩%� ���,��r�؊b#`T�eT09���ȓ!�b��g��}�8�F��-? �ȓ
K|m�ș�VṔ���2�%�ȓ"R�X�j�4JN�1�˘X�i����̹	_�jZ��1!g��zܶ��ȓgil,*�J�
j�Ne��i�J%b���f	�(U��:���G��$Y^م�~r�� S�%T"���k\�jx�ȓ|4�1�îJb��@ӵ�ݩn�V��/[`�"�v4�R�!ʎ<��M�ȓ`:��z�ؚh�J�Z��$HY:	��H��p�m�C1��!��B:��0��EnjZA V;9����J[
2���	��4'J�EA�IVW&��~�(aZ��ӹ�>� o�Y�|�ȓ�f�A�
Ο7�H��M�$�����mޠP����/���ANXo*�ȓTv�����{ ��-7�*h��I��sB�8�8���3����ȓNe*M�悡;������X�o��!�ȓ'lj�#F�m�+R&;�|��2)n�C��0S4���T:
b���:�0!��e֊��)��ͷV��,�ȓ0�&�8#���� ع�L�����;�P�AFd���,w�6d��r�EQ�( �gVlɦ�M,H��,DP���|�I	$G#\���ȓ"�)���E�B	yt&B�^�LɅ�4�� ��eëF�ڙ��n��R�p�ȓp`@}bŇ�=�$�AUN��P����Ii�~��T�w��5-�u���� ]�L��;�>�̏)?B�"&�;[^T��R'��p*��x����)��6��e�ȓv: ��@OL2$��	�Ǝ8@Ć�_��U��+U�Eqxy ��"4���ȓaq$��̑(���ВX�C�d$��GȄ�y���_���ȶ�\1UB���f�AD�R&�
4f�Q0�a&[�H�ȓ}��+䈃5m�8h�1��	~Ɇ�ITy�GE�KJ�K�M�>yR�y��̈́�y�W>.���+E$�H�s&+@���'Z��Fy��>a �/F@����C��L�XCt��E�<i���_�P���?l^���p[��x"o��h�ΔY5+��C����ͫ�y-L>E�Ӏ-��rc�cb�0�� ����$�1gkDhy0n�U��Z� �j���3O����  T��&�ϙF)\m[�"O�I�H*u�4P�Q�۳�pd�0O���D $,�e���=;/�]Iц�(xMa|�|2k��6��m�A &C fz�J��yk�4f_P��C�v�* ��y
� L�yԅ�!�Z�z�C���p
"O�M��� n�}����.}T�qA�i^ў"~nZ�����c.��_���	����w��C�I��4�ծ�8.�� �J�2�B�ɫd��袔��x�x5�$�r�C䉢=���ҵm�&IT-� f��~}�C�I�34���j����R+|��"?Y��)�7I^�W,��cLԻ�H_ ZJ!��}m,qa�a^ hSU�F>&!��B��Y2���l4�
*D=3%!��
�;8��$e1�*1�I�?!�đ	,k }Sm�N�D�!����!�R"P'�\ ���]���Cɒ�sR!��LgL�s�ө�d�0�ӷL��O�=��!@X6-Џ@�D8T����F��6�R�d�!���E���<CڨТ5G� 5���=�|�*O���(e!��"fH[����D�:�!�=\��%i���!#[1r�Dߩ mF���Ov�=�O�`�`��ǡcƊ�saԠ	]� 
�r��<, ���B�����d��m3| ��(,�M�Ԧ�l��|
�M@�"M$�Dxb�I|���IL0bq���f���́�4!!�䓘Y;"-
s��? ��:�럂K�!��1���A �mn��v �{�!��L�.]ḏ�Ɣ���)ҡ&t�ўD�ᓬ#%� ���ӀC�̀b�)C�BC�	�LQ
��ֈ
=��yP��r4C�I/Y�0�j�-��a�љ!&L}�B�I=Ɩxpan��b���R�]����U?�?��j�� hFܪ|�d��b\s�'��?�[�oO�`�[�͗;~����6D�81��D#K�u���&F��Q&�t�<Ey��ӧHܘ�*p�_J����N�Q@C�ɳ*�����b����[��FB�	.N��]S�dZ��%B��&Z���d!��3]5$	�c�̣Q�H�*���*|�!�Z�Tಡ؂��xoH��b*Y�Vax��ak����iˁ"�T@g�!4 B�I"S��{g,������g�/��	��?��}�����A6T�Ar��w7�s�iܶ@�!�$��s������7\%��HސWx!�d)S�P�`W����Q�Hw!���Z�h3�*Z�b�޽
a&���!��<Gz�lrւ>���1��,}N!���w8���7�$���䕂-!��I�=6��J"͓/Æy)�Î!�$�Z\L�*q �3��P������!��
9"����'˽z#�!: �m�!��þ#Xά���@�-��GԟG�!�W�9q$���Ӿ!���
	��!��Tv��(�NP�T��Hʪ5�ў���:>��pj½&P�H���,ELB�-k@��@r�ȲF����%�W&6�{������mOD�̹�_�tM�5Q��H��y"��x�J} F!65���R��y"�Ҹ1�$��PԪ5qX����y�a��I��9z�k1#�P���C��y�C�O���W� j.��J��!�hOL��IO�3�r�A�l̢K���)5n�:�!��Բ%".� Th��1��xvm�+m!�I4I��؋B�bath�8��N(D�h逎 ?/B��(D�=i���%D�8a�N�!ӄ@�d�O�6���Ҷ$D����P+޺��a�k��\"!�� ��@
ʷ�P�����B�VT0u"O����̞�e��<U��PzAv"Ox;�ԁEy���R�\�,��"O�M���<O��E�1��M��g"O�e�$�Z������6,WXt��"Ol`�ŗ<�z}R��QwJ�D"OzM�Ҧ
.�h���c2F���"O�ٰ5Df��`I�00XI�"O�iR5,X>��h�,b8�4"O(�(��؇_�<��H3;��9�"O*��5��G���S���H����F"O��pW�pr��ZGő'(�@�2"O�	s_XGRt����Z�YѶ?O��=E��dS�h�X�r�Dk&� �B��y��-)*���O>R6�9QNß�y2�Y�N�tP��I,�|�elô�y��M��&��D"o�jQ�2&��ygYOR-�v�#$��8�j�,�yRB�!�RX��@�	a �ea�����y�GY06 J�1#X�+�� �P�Σ�p=)f��>a�<O��
a���0��a@�E�<��Yys"O2`"�I�-).�=�7��	`��L��I`���	���%J��Y=CF*跠Us,!��2a��"���,\�����*!�'m�t��(��v{l��Y�!�d�:�2�IM�5b��ؾC�!�U�h���z		���S�Q�I�!�V;��vE	�sV�1���
+TvL��B��=8&	@6x
��oD=O.��ȓb0�JB�\*U8�84�25��/n��%��2jpգb��9Mj�	��]sV4�p&
��Ayw�K�S�r��ȓL�]�_�F�z���C�0�>�ȓ3���BD��	f9e�#���ȓ��
Ƙ#g�q�"Mbx�����p�O@M�q{��8{����ȓ7U���B晭tgmk�J�V Z�ȓ:��A t.m����m�!m����ȓp:2�+S"�2vt��#w��w�Lx���0��OҮYT�u��OZ��������������K 2l�ȓteV����9�|��R�#E��\��Hd4�36D2��]Rf&[�$|��pD�ٳ�#�>�
�V�G(t1��G{�4A��IߐeŌ{p�ȓEP�J3IT����!�l�2��E��Hւ rS�˿f�r�y�mU7a� ��,� �"�G#y����u#�)Oߠ؆ȓ~5��g'ʹGg���p&S*U���ȓm�%{�	�$�|Xk�(��Q�b��ȓP�9�Q��+~�@�1���<��i�ȓhh0�bN+Cf�yq�1)�$�ȓ�8��c��42~�Y��}��T��7W�0�IK�o�lhi�L��U��=�ȓ?�n}�Ա�*pӖ@N���ȓ&h=���}8� *W^c���v�n� ���/�4{b��lj�ȓcP*��uJç?�f�8�h܆�I0U��땩n2�zb̊~v���ȓSI�Lx��P8'����Q�-D�X���*�&`��ΤH� `�D·�R]���ȓ<"�Y1j�&3��9b�,Y�[�$L�ȓ?V�����G8�A'�ZCb���ȓs&��l��t1��f�>j�e��S�? �c��E&O(�iԯܧ�ő�"Oh��!*B�m��,� �Ω"�Qf"O��� jDJ��+5AXIIA"O�����7]��,�F�5Y?�ԑ0"O`iI��U�l8~m����?~)�B`�'���'���'`��'2�' �'�p��m�|��yV�M�0��()��'�2�'��'<��'��'���'�`Y�7���H�"
�}a�D#��'_B�'���'$R�'�B�'8r�'T ���ҀR���D0^��e�')r�'G��'%��'���'s��'H�e�׀�q��+�`ȓi	 H ��'dR�'{2�'R�'�r�'Z��'b����F�O�=� DS�]�r����'FR�'Mr�'��'V��'���'�+�戞G��p�ˎ	��	S�'P��'���'�R�'q��'��'^.�qu ��y��Yp��Ҭw��`!��'"�'��'��'���'�b�'�5*�&H�YW��z��A�K��hY��'���'���'�b�'���'��'�V���� �>�	�P��;2����'q2�'���'B�'(2�'1�'x���/�2���k��^kBe���'���'���'?B�'���'"�'��=�7=���@�NU�\<:)�B�'���'���'#b�'���'6��'�T�
u�3yN��h�&s�
�x0�'�B�'�r�'T��'�2C}�D�D�O�DRwO�oP�t��n��(ŧdy��'_�)�3?4�i��H���@c0�#T ݏߠ=��m����$L�y��v�i>���M����f�ԙ���D��>0�R�  -����'��"¶i�$�O�R�昅b�r�`Ãׇ^��T��,�M�^�cF �Iğ��'�>Iz�AB��x�ӤՏg�zL:�F �M�5A̓��O��6=�x���]p�d�"*�x���ئ�`ڴ�y�X�b>��b ʦ}ϓC����X���8�I��C��Γ���3O��N��)0��4���;q����f)D�`c�*��~��D�<�N>A3�iR�;�y��Sh6� ���_�$	B���F��OTY�'�46�������Ν��0��ǯ$l�Jb�Ǚ	��I�_�4(8pbX�0BVc>�i�b�غ[E�'e��&��)H\Z5⃭X:r<�DV��';��9O�1�O�>�:D�t*�# ��#7O�lZ�(�F�N7���4��qҁߝt����9�t-�6Ox�m���M���L�z,�޴��9_��AAў޸�"H9/5J��O�f
��uUd\zQD�g�����^'~T0��îi����Xv&��3�:زm�>r
J�@�	uH���"Oj����X�0����)��|R>x򔃇:M��s��Y:9�Z�i�d� A-P�s��H	ᄯ�v��D�s���&��$����%��Iw�c�&g�̸ӢHW5`������҅U%��vI�>'�,�c���e/T���a�,s��X#K�/2�p��#$�.�
���9T�(��H9sBH\�.7��O�d�O��e~҇EIU�L;��^�<����>�Mc��?�
�l���4�>�������O'n��%�1�5)��M���?���b��$����M eP>�=�F$�5�\�n�,��"<���D�'���h��٦AR,��b��Ge��AE�`�
�$�O^�$V�`�X$������	�f��ȃ�E�1w�����N�"L��Ё�O��$�OxxX��D�O�d�O��1�d��{i���K=��k�N�ަ!�	45&�4xK<ͧ�?y����D�)�|����A<�*�-$>A���S���� 5ڶc��������gy�� (Y�,�q���u��9��K�����,�D�O��d�Ol˓�?)��g	�	��3��8I��Di@�B���@̓�?a��?i(O>�) ��|"c�R,��1�G��� �l�J}b�'�"�'B����(��%m�b�;���&!�+�pc�ȥW.���'�"�'ir]�\Yg�ĉ�ħ<LB�8)�q)e�F<7��Q�i	�'���� �	1v0Xb>)pd�:-j�����ϕp[�XH b�>�M{��?�*OJ�+GK@V�ğ��s�Q@2L� Vw�е'[�D����#}ӄ��?Q�� H���|B���nZ�0_`�2)�"��y`���4��7ͫ<m׀'�vJ�~����F���AUK!���j͵_�Ș�y�h���Ȏ�n�<�O��L<!�I//����""Y�j�$ �a��M�o%�M[���?	���ⳛx�Oz);Ca٦3h��)��D^�0�yÀ`�Z������'��yb�']������	Ob�Ȣ-�C��B�`ӄ���O��N$��S䟔��&��Ah��I�}���hi�_ 鲪O��d�OD�9E�$�O2��O"��	K�^Qz�A$��QqL�ͦq�I���d�H<�'�?�����$K g�f�ٶ�V$rЛr�Q�G�ܔl���Y�!&�	����Iڟ8�''��3�1�^���]S�Ƀ�	C�t8�O4���Ot��<���?�g�,O�^H+$�2h�ɓ!� (b��<����?Q����T�@p�ͧL��e���Ӻ/��0%G��0�'�"�'�U�h����A��~�������3V�(j�N�fe.��?A��?!���?���($���'lҁ@�`rjd�t�V!Ns�9�Rg�A��7m�O��D�O��?�Pn��|b��~�X�@�hT�ǩF1D���b��1�M����?!���?AP�ӳN��F�'�"�'��T&��{���2���k�1���N��7��O���?� "�|����?y���|n:� �8�E��;zp�;�'P�r$�JU�ib�'Blpp"b�����O����)�O�i1��](/c�|;֦�wK8x٦�t}R�'����Q������O�[(ID,��c�S%i�Ċ4%�)g�vk�w�
7�O2�d�O���韂���O��D�i@�y���J�>�j��_]��o<<PY�'1�i>��|*�~n��g�����D�|�B�9A�i��'�B(ٮ9߮7M�O���O����O�P������h=�:�����+u��6�'1rm�8ab�����)⟐���OT�A��+q�}�6�	�d+�O����	! I���۴�?���?)�4��`?1L�36a�L�[V����Hd}�`�/�y�]����˟T$?�*!�ܞW���{�#�VT������%L�b�O�ʓ�?�,O��d�O���7����>@Q*i���-#;��A6O
���OH�$�O���<	���_x�)�e�!"�� �g�e�g�Psb�6\�H��yy"�'�2�'���a���eZ`�$�X|[ c�\���Q��i	��'JR�'K��'�-�6.f�r��O�A�(����%��6~�A��צ��	����	Py��'7��d��@�ID'T�Lً�F��hL�V�'���'pBoB�(�6m�O��O���l��̵M
B p��R:Mn�͟|�'��Ι����'#�i>7M޸+����f��	 V�|J%��&a�f�'�R"�;H �6M�O����O��	�������d{2���%�
�`�'�Q�>�B�|�O��$���r��~���XQ +�؉n�M�0P�ڴ�?���?�'�b��?i��!�X,q��S)i`х#�fj��P�i�愻4]�0����O�	�Ob�p��� w.D�0#ܟYS�ո 
��M��ǟ���(5�Z�;�4�?I��?��?�;+&��Rs���Wedu걦�.f��n��ܔ'eVpz�����O��$�O��zr��
lY���1.�7g@���k妹�	��إ�N<a���?�O>��<�X�.޿O����$B�R`��'	�Q�'=��ݟ������'���H�nn�Q��:\��8��K�YpRO��$�O��O���O�;ᮝ)��Sr��w�bTy�]F��<���?9�����D� �ͧ&��ӅOܵ7�Y�.��h����'�B�'��'�R�'G��'��=1�n�x�����%�d)�S
�>����?����$ ��&>�[� �-d�貀F�H,.!�
��M�����?��4X=͓��I0����� $�,�S�k�j7��O����<р�L	 ݉O�b�O��͚��\�;M�!���F�%�8mcu 6��O���ɝr��$)�T?]�aG�
)x#�'8!؍���p���d�p�I��iL�'�?���8��	ɶ� � ��#���Z
�1e�6�O�䎴6�@�,����`	�&�>F�0�*��2H��ݺ+��6��O��d�Oz��	Z�	ٟp�P�M�kF�s�ŕL�~MP�LQ�M�&	F�?�*O�xE���'ϮI+�k�Vś��T�b�1��g�����O$�$Ͱd)(�$�@�	�IC$r`aD�=�Aa��Su��lZCy��'����'���O���O$��均{���ck�5*�5�dX妥�Ʉ�|M�N<q��?L>��A���K��G���P[ㅓ�_��'����e�'��ڟ0��؟d�'9�H��@	r���Q���G.	c6�^�Y��O�D�OO�d�O.4y2�N�\2,�{�
�@7����ڹ�O���OD��<�� ǧ���1�ʝ�AE�/ZJqW��;*���̟��I|�̟��I�
��U���Qh���F���M���μw5�h�O��)ֈO�Uabr"E(���aY�h��t�%R#*t �A��2#r½�w*��f`�D@7J��X�j ��,���j�-ɝY�R`!Ef�Ia�	��AH�����(6��aj���t�Xyq�%)o0���c�� �@���[v�J�˨O8 �s�C�-)��e��Rb<[Ǆ�%9G\-�ҥ�gj�P���Ķ{P�)2E8<qB����N������H2�a����1 ?Z4y���#s?���d�0�v��a�
�)� Y������	�X�	=aP���
ԄU���c�֚z?r�+�cV��@�9�N!0� ���J#V7�I"��ﾩA�CU75	9�\�20"v�[�SS�u�"� *�(�M;Yrbe@��+5z���Ғ~��'.�4�Xu'ݕ`0�L�D%��Vc�yڂI͟��<E���D�j�Zq��"^9�͇ȓa����4�T�)�ޕ�#lC)��(Fx�� ��|��x�<h��JZ��D�T�N_d���?��ŗ<��k���?���?�T��8�4�r50��¡=Ⰸ�#C-l�2�F�ڟ\�PÐ_�L�w�_�W���ɫI��uH��K۴E��%������<V�hRK��Kz�Y���?�=i4b��X#���E�S=��5N^G?!��䟠��c�'��I&WQ�0���pXƩ�f`�'T�lC�	>7X�Ȁ�-���A��X�7nRh��4�L���<��	�x���N�8�zȀ��"g�i�u��H�b�'b�'34���'�27��X��N2^�$�QFA^��)y��YY�T�pGQ@��EL6<O��8��Pk���c�4?b
d�Ӥ�-#�P��w�J�'[:���@,<O^���'iB�	7��t�3�����3� ��rpў�E&�<ӦQ�iI�������y2�O�� ��O�<���AO	�yBda���d�<e�5+
��'-�^>m{TC$w�B|L�~к�֙}��m�Iş(�	)H�؇��?A�B�q�� ~̦4˕ޟ� $�;c�֓f޸Y�%X�R2�1���"g��؛`m[�,X��iWV�
�L�3�<ոR`��{���p��'R|pI�vqO0���'�N#}z󭂕Y��x�SK��K(��k2o�I�<	��O�tűU�w<&�!FȄF�DN<�#A���)�98������$�y"&��7��O �Ĭ|jQ�M�?���?a�WD�H��c�I�rh�roRz��`��]P�H9'�����e�2�?}�|��~P5� a�![��t�ggD�t���뇻T�h3���x�2�� �����h��I?��Y2G�,x��)�(qXF��6 ��"�̙�W2o4���O&=µ�J#e�f!r�bF�ْh8 "OrU��SJ��7����8��ɥ�HO�	�Op=���x�s�^@�ƭz�i=�?!��/��@$�)�?����?y�H����Or�$� q�^���oզ$#���N�v�����4^)&1�Wb�G9ikԌ�?�=�����ٳ.�53�0���HQ�����D���ݓ��NX�T���{
Q� ��@R�C����To[�{���jdʥ� :��"�O�5ۓKI}��82�B�>��.�ybd�M�x���d�8���čY�X#=ͧ�?�*O�y�Ə�ԦaY��ۿtfT����<Qq$�Qҟ(���Ɇzje����|ϧs�����ҍ��� !�Ș
�ɻWqV<��nQ�QiZ��Ӌ̳6���� 䖟L��K��]#N��3��˓���
�f �2l��oM�_���(��� ����d��h�@}��y��Za�F�J1�� Q2�I�FLS�'oџ�*` �I����;G|6��0j-D�X��[�?���ٗ)єl��d[Pq��ܴ�?)(Op̒$�\���i�F_>��e�(j�,���M�!�� Z&ͷ�L���۟��	&V
�z���X���ƍ��B�{����"�KH�h����N3N�E$剥v>R�ZqM��$x�<���*^�B�j�������kȄq����e��^t��#¨�X�%���#��O��E�d��-���:�$O�MX��1'��y���f6�Z�+� E����IB0�0>�P�x�i�	D?R$�抒�6��$`Q�-�ybMIt�*7m�O`�D�|� ��?���?�0�B�=�Lݫ��D�y����G-����m��>VH��Ɛ	rǘ;�]?Q�|��2��)ӧ$F>[?�!3� ۽a͢�Qk�+}%�dv��!k~m2���>�n_��$8�N,d0�zWV8
�f�е�Op�&�"~�	�jB��kc���l�p {�+�;hY(C�	+e/Ιi&AZ�Y�Ё!��	>R#<���i>��	�r$Zq��aF-}8�C��6'�T�Iܟ,�!�9	m��I͟���֟ �[w��w���yeU6Y��y�C��;a�'�lq����=� ��m�HH�DʙNm�z��O?���>J���2`�\ɸU�?@-�1�F�$,�	�Z��y�Iܟx��?˓�?�+Oj$���7�2I�2�׵C|D��"O�(�P�tpf, fH�-ea	B�P}�'`����$��,�;]�Y��T�E����"ti
)����?���?�ҁ�1�?i����T��?���-�, �I�&9�<�i�֝m�j`��ɹm~˓mn:�����3J�@<I�A@�P�vD��AJ��ۦ�ɶ�K6iZP{��FVc� ��9D��0W�P!J��8���?>c��UE6D�h�P���v�*4ύ9V��A��s����}"
�c&��?	+�@u�T��
2t��DK�.N�~A"��E�(��$�Od��U5D���z� T"9�e�wMƷ~����OI�HDD�Y�*����ٵU;@ᒏ��M1�I��
��$���/g�1��c� }1B�����,�F�H�)�!L��qW�'�'E��;����6��-mܡr�Ͷ��A��!ȑg����h��D)�+W'(C���")�2|l̊AO+�Oh,'�X��Z>�.L2@qS�C�ji� X'$L��MS��?�)�^�iSg�Oj���O8�¶�G�jam�%��5�񣳁�[���0�`��l�S����'t���W2'��pr˜�v׈ܹEԔ.�zU��d�7� i�kć᨟�0U�.��PD��	a��3χ�EfS��'i �O?���t�����砠q�/��8�!�ğ,/"z�X���� �RO��z�T���4���ĝ.8��j���J<d�!ЬV	u N��O`8�1L�F�r�d�Oj��Ox���y�gW�0s,�Y�`�?���O�7F���b{^ b��1S��*��hO���-ր8�ظ�z���j��LƟ@�p��-�]0t��P���	$#N�=�`�u�4�j�g��k�I�I����O����O�Y�l��y�E0��8��>qɄ)ᣯ���yMH�V2 �Vn�*;-���c�m/z#=���?�,O(!S�L�ЦQ��'YT|Τc6�XR:i��OY՟\�I���s�y�Iן$�'{=�	��ןl(a��e�2�R�JDv:�Ç�8�OV��WX�� DD9�%B�5���A�>���'U���uP���͐�>�o�~����G�yoq��i���y ��A��y��׉|���A�@��wˀ貏�?�yR!#�I�6�i�ش�?���i��"��й�lߺu���*�e��E��`���O����Of� �b�Q�H�0R!E��@��|z&�`��eM#�msPb�D�'b��Y��&� �
4CA#2j�O�
XCRBRx�91��\�)��䙃��퓠a5 �cd	�?[J<�Xj�B�I�D�i��
�`
��s�����D�b�IWV��@(ϐK&|PE �t�P�I3iv0�ܴ�?����߸E(���Oj���6��h$.Q�����R�P�]��/)�us6�>�O�1����-�z�!2�+v$�<�v��=r�p��sfmkdD�(_�݃���'�0�J�!(#�xh��&��RX�����'���On�EMVm@����N�2�"O�`��@�e�N�34b,��3�HO��OJ�#�ћ|v��P�� �Zaa���O.����Lʘ�k��O^��O��^�;�Ӽ;cE�.�:=㱯Q�t�:�+
��WT�d����(,�ZUa�<x�Ș��r�Q�<Z�JG�h!1K�|�JQ��M�9e�t�8�!��Jߞpc'jF����5�X���U#h��I	/��y�E�ŸO$�5�ð�p��-0/���Th؞�{��Zh�Q3D��#��:D���&E-q�zu8k�*°���HO�6��ڸe���nZ�93�P����3��"��X�r�4q�	֟h����d��şH���|`+U�HD�� A��'/�T�����_�M�MW�*nB��	ߓ��嫢��'U&Lx��&)��8q�AD?h<�cBf�.�~��C�B.��`��}�|m��Y�Zd.�3TƐ ��Вs�&B��?d�� a  ��%�L�`�� 0dB�ɑe��<�$-أ��¦��W��	,�MsL>�'��Qa�F�'~RR>��#�ɒ0�ZQ��'�w�Z-{ �	���O���O�!�5E�2a\�����T>��-K�H�J8��j���X	�7�3�Zl���+��{�мʄ�iH:q[sh �|�k@(��=�ġ%��i
��h�'���2��h��#.86����n�">���"O 0��/�
J��c��A�.�a| 6���mD����D	=���k�0{�DF�=~l�lџt�	y��)�<E�'�Ҫ1k�l�s�Ñ7)?(������:�T��UɆ�U��򱅂�Lג��@m�h����+J�ܪQ�֡&&���O �:-lu��`Ķ(������G�D��������X~��5�I����w3�5�Ыڗ.�谉�WQd�$x2X"����s��r��ɮo�k�E�6 �j1)�"OF��m��M��M��㚘��z����HO�Id��BRh�}J�q�ƌ
p������OL�čj�\�K��O��d�O��DKӺ��Ӽ�D��CQ:4�fMʀ|i����Z�IѼAq��[������).�|U�'	qQ�v�{���16Tttt5����
SW���n�YRqyWfc��S-O.Ì��D��'�L��^�Y�*������A�H�X�'�����'�2���,O,��<���2,��tQGM�qlQ��m�T�<y���;�)y&��m�j����G���ݟ �'O����/wӔT����;��Y��͘<����O����O����84\����O���X�-fz4�P�<a��U���D�5U((u����(�
=,�NtZ����O�m!�	I�a樭�����@D��5�]/E���q@��a��H:S"ڇX�0Qc��\�&t4%i#���&�bFc�R�&��!V0��V�܏ؘM����䦵��Dym<^t�O�iY2�C�vܪ�s��/[_�����
�0<�����g���,�+�4���Xl��ѦE�4���*^m�������d��9Z����1o�����O�QrD����'�R�'��86�ړx�r<o�/��Ir�����@)M^�YB�	����딫�(Oĩ��nN(�pX�i!:�(e�YM�Ĥ	�Վe����Ք��hZ�I�t�%��{�%��?Y!�iOZ�(��Q�w�,|j����]E$@r���t�N�D%�)��<r#�8��a��
~.�kb��x�4L<I5�ӟ"�X�G,K�w�t@����<�V�ośV�'��_>����8�I��'Ő�y�fQbtm��n��!�.\=�I�Ie�S���ѕk)+�H8U�<KJ�19�EkW�O?���90�&��dE*N�
���D,Q�x�#S��On�&�"~���m���h��9�X��G�F�4C�	:��<0�h�P.�B���)��"<�2�i>���
"��s��J(2�~�I@��+�dp�	��b��Z3>���IȟL�	��AXw��wJ��P�#cV� `C*U-5@ ��Cx�R%�O��;pg����!<��a�$��>���	#�Z&͖Y8b�Н8jDc�ɚ9s�b��YJ`fDƦa8 ��}~
� �D�&%گJ;0�ⶀ��ݰM���OpE���'����D�pdBE�Q�
�L���j��y�!�sNL���3����WJ�F��Gz�O&�'�rq�t�`�f!��	���!g�ߝw�ȡ��I�O����O���|�r�D�OL�@�xp����m6%{�
R�y��a"ǈ/x�d ��[+� ��ćB���O�Ġ�"��!��! ��ǜzͼ���Cɳ4�>�[w��F��8��2UJ�nںK�Nq���G�	�I�F��Ǧ��'��a8,!Hl�<����(=D��
� ��O'��KbD	�ȝ�6?OD�=RA�1����Hۗ`����g�<�T�i��'��� �j�(�$�OP˧Rbri��D�P�p�0�.:AX���`ƕ�?Y��?��!�>��ɂB4g��EA�(P'r=pj��K ���j���@�!�&.kG�	Fy`�;2�jxk��>@N��U��3P"4��s�F5VDܸ
F�V
;���[�#�mGyRn�6�?��)]2B�u����4eݼy�5�H<!�!���`��;���6��t��e��,�a|K$�� ��Z�J7��F-0Ń۩J��L5|D8lZꟸ��T��hO�S�b�'gr.�<Y;8�A�2D��!�v䘊&�\t���$��s�m){D���iO�t0��w��3*d\r=���ؒcqyB�$��@7�ۛ�R�87"�o$D:P�
ӸϿe/t,��Y�쟕.�(��C'5P��a�9�ɧ��r� /t����SԨ��n�y���oY��#�9 n��*��O�HEz�Oro��/�(�Q�� Sϖ Xa_\��',b���G ��'���'ݔ��Ɵ�ݚ:��r&$Na��	4��Ђ ]�<�!
a ݝS[�j�m�?q�É�4�1O��vH�AҜ�7�ڟ9��.�>P�G͟&y��@ik P��O���hp.�]��EiJ�sY$�yt�G�q)�樟��"��O����
�z�C�C�V;�\���«v�TB�	=����G� _�b���튀IL�
��4�Z�O�Qh�F�Ϧ�Y⋣$�.�Z��VG��MR2��ܟ����t�����	ϧd�<-��ޅLD�(#a�I�m
�BsbV�4�l�����/$���� 2@�����=e���I��ζ-��g���Z�+1c/u$2��A��&HB�e�A�K�@�t�t��S {�buӴ�J�䇿O~U��E.�AS�"O�DQa�S�@%�c��2!z��q"O, g�B�I��³gی�up�1O҉l�X��9�T��4�?����IV�M�&!�A�R2��sc�6�$4���?��?w�R��̘��I<L���S�"�o�px3U��U�Q� ��+�'QN�i%�
@Q��͉S&�Gyb0�?A7�Ӝ8&V�K`�͚\��i��lB�ɰ {:9sş>^�S��
	�.��DGU≖�9�fJPĨɶ�G#`�&�I��LX�ٴ�?!����	��lo����Ot����VmC�-�-*Q�)�t�G� .�hr��6��m�Qb��|~��/�0��Mց[�1���%�X|�tC �v�u�pCL ��s��/c[��bG]>V<���F�8׊�Ï��;n˲�)���>!"h�8�̓94���Ƭ��?�4�|���'�\8*�`��ɊX��h�i�<i��1w��qXҪ�t��+�ob�'�"=�'�?�a�A��g��,F2,q+�(^ �?Y��)�b�q�C4�?����?�O3���O�6C=	c�W�y� hi����n�����}2_2��-q �	d�2E�vm��~r����>I6�(\yjRbѨN��ْa�C[?y��Sҟ(ۓg �z��
�dP��H Өg �I���B�"酅S�VL 4��#{����)�';88�p �iM�[U�B�Q1J�*��_�����'���'�2N�G��'~�I	"�m���̷b���eͽD��ٻ�$�mNǘ�i
�'�1�/	�$8�&�P�aR��W�!�h��G�]�	S�y�@�ͽ><Ub��$��O(\q��'��6-ߐdUbFはl�ީ)D&d!��-`ϔ��p�DWپH��(E!��s�ޠɆ�w]bH���-*��e�f}d�i���'���b����[5�B)�P�\nq�����L�����2c����<�O�����ъi�q�tM�!���򤀛]��?���㝉ڐ���j�7Vd�E�9ʓ]����ɋ�H��m���\�H�GL[3s�.=3�"Ob�`���M0��p�̃�_G��y�'��O4�XD�Ւ'��eJA�4D�}��;O�0��9����$�O#��bQ�'���'@6�QF�;F�f�RS�����keJ\P��J��ȵ���;��âVP��s�s�H�3@J�"#����K�7��$cH��uz��1�ãG�Z�@oN���K��ǋ"Lpt��O�.�t�a���}��jϬp��`��� &��� чX��0����MkCS��	7��� @%��OD�0��$��nK:ú�+�9Op���O�⟬��!�  d�M�W	�p���� �Ff�'J7m�ߦ!�ɝ�M;O~2$�+b�Zi�w��7w���3�� �?���U���/o���	쟐���\wi��'��x!��ȚXw��˴�8=�{�'t��rl�C�.(�-� E
��(�>�ф��'M)@ Y"c�E�1�u$N�4��	�T�$�l؞  4ϐ6?���I�KY�Ի�L=D��b��-��Y�->vKr�hbE��HO?��$���SAK��P8"B�/o4^u��$B��P9�!R�i�4C�	�+f�(��J�m��)���Ϯ%�2C�I�Kѵ�` �!82��'��B�ɮ$xp#B<O<d�$�غl�VB�IA�((��|�l�wI�PlC�I6�݊�.Ȧ�Z�J�d���B��:����͇��C͘�pB䉟+��4	�B��>���j�i�&Q�2B�	N�2��Ckguxa��!ض,5B�I1�bm �-�3�\=��Ă2�B�IlВ CNI#'~��hD�¿+�B䉶%��ѪB�D�1U��	@�B䉸h>8�� &R>���I���3Z�B�I�5"�$�\�#ߔ͂dbR%|�B�	��p���4D�bҎ��2tVB�IlHP��eGK"{��آ��!-�C�I�8�r��F,7a�H�����C�IHj�E�vʌ�v"���u��+H�C䉓�6�؄���u,T�7ƒ:l�vC�ɷR�Ia�O�<u9 �VK�S�JC�I�	������͓+�Э9�DM,��C�5r|�=3�#%5��*Ck��m8�C䉪M���*��ڽ[����,�$r��C䉤au22�MJ���(PϜ�C�Ia1 �����<hd�ԍ\H�C�g<HpA�5:=z�j%&�>Z:`C�I0,��P����wBd�L�n�VC�I/\�]�@���%�}#��X/!�RC䉚^5�jՆY2~��)b�ɣn�nC�	9޸�*���BtA�ƌ3W=C�ɛ?u��K�nξ8�B!����T��B�ɿzIXĂ�$�	�Yp�Ɖl��Lc��E��'S��ɲ�hOP�c�D�O�8��#e�2�h��'��|8���>i�Or9XČ
"@F��ȱ
X�{�xq#"���?`�oX���V��	n2Xk�g�ppE��
��p���J~��ل#�W��d������'.�I=��8ڡ��Oծ%��B�L���͓]J�~G�}Ռ�@��3��5�S`ҳ6���S�=�M�g������}�uH�Z1	��7F�=����C/�O��#��S V�dj� T�0	Ȁh����V��`�'���� L��m�2!f��� �R6O��XCD�2'�60��MO�����ɬu�d)qfg j���@_?��)эG Z噴C�RX��;Aڪ���E�	��(��iG IY1��n= ��$Z�M4ps�͟)3��@��Q��d��H��M��
O����Z��|Z�M+��,5m>8[��H�d����R���P��S����7m��;�dr�.Y�(���C�([�;S�)���p��$%��9O��	��]�_O )[Q��5^��e��FE4ZT��$:m*��x�ʺT혐��Ɨ�<B���*��;V�'�֤hÌT՟�v� 7�P�ڙ'�L��"�6�)Q��G�~�b<ي�d�)"�ZeԎ�e*��J��B�g�󤎭[3xP�F��&k>�J���w���!%�D�j��'�ڸrs�����HH���
ts�˙�e��Mf��OhYk��Qg;�8ZR �6%^�HJ�韌Y��`׾E�"@��Ig�$�B4Ĉ�J�v�Y��'��dx�K�&zM��U�c+
M/�NԐp�$�w�Cʼ����j}!��ߟ(�*���!]ظ��A;<O:�R�]X���I�7b��x��
�S�L�ǧD��$c�ck�\s�d���$��:�J����\V��D[� Ej�>0�<��@͑;ɉ'�"X���7��h)rK��`��O���%�xD{%o4J\����'�\ϓrF@���̟[1�Xs���e9xEE|
� � 	�-?#l1%FZ��$ڀ,�A���7�1�$���^�	��Oh��+O���"��>R�@h�P$�(:1��
oBp�'�>�Ok�A_��1�D�;'�`�y��=/������'�^ӧ�F�|ء���?m��%g�~��A�XAX���C޾y|6-7 �(p� C�_[|yUoG�ː����L
���'/���N~�k���Mە��d� 9 �/�"��V.K�^��9�!BֱhG�\BЩC���(ǖ]@ԡs��d����'�Dɬ{}�~�j� �GB$�J(��P�t��<�ˋ}RJ	�<���ш����')'�HO�HA�m�Cl�ك�탠v� ��͛4D]f 9��Y>	(e�xZ��D2)_���5\.���6��I� 'Аh�=R��_h9��ɓ\���(�V�F�R��U��>���'��:�4/Û��Y�(�f���~�7�O���GE1��Z���%�B����'n���BҲ9��@����jV�)��ù.FB)���=OR�!��~8��f,�ʛ��Y�x$�eQ�O뎙�|"�'�T��b@23���F& 42"�Z�{
9Qf
��
�5c���ӡm��y��<�5N	q)81sʝ�&��9� ���c����Sq}r�	%H.�֝r�'P��ycF�@���!�6p�t�)m[�wv`
��ή,�i3C�O��{�+�O�N��/�p��Vx�J�P:T���Ol����_��J'�R�H<��@A')�<���4�	5��S���'���.�'{g8�cpe��]�R�R��	�3r���D�&g���C���9l�ѓ�ɔ�cf|�Q"�^���3Şx�xBGV
��/s>J�x���?&شm1cK��3�\���D
[B"=����e��d&L�L�Q �
��?��6Y��!䠅)m�s�B�t��	G��Ik'�l�d�JS�0�Gz�%�Sj18f�Q�h�
�� ���M�r�PFG�5h�L�V���V�[�|FxZw �غ��њ �r�F�8}���*H��O���	0�O`�"`�2'�@��Q(���U
FB�^!sF�j���O#J��XЉ�3jԫ}`�m+tn�+))a{2M�i��z!-�9 1�	v�ڵ)�B�94/Y�g^��f�A~r`N�(O��+W�)	5_?Q7�CA�7m�?[�td�7iE:Y΄å�clqO�����1v�����+K�	�҈�v.���'av�S�HćG;�-���ָo���I�'�>=�Ed	�'6�|���\�p��i����%v�;�"E�6IZxh�%Q_��}`�/ё#�Rj����f���u���Q�\`ӧK>�Th��Q{MЉ9T%�H�%�F��lQa|�;0%t��39J� }ӶC
:[��RB��;k@��`1O��'�����mX)Y��}��HH����
��=�Ԋ+O�A�����,��Z��A�ܾ�I �Ђ��L�%a�sb����AG,*tQ��c��7�3��j�nH��,*Ľ"��3xT����ϯ"f�'p�i;r����4��S-������<ͧ<�	a�ԣh�\�+�� }�(��k�0FΛE�=eb��9����)ғ��5L����E���H���腉^�C����'�{̓����$�t*�c���.g��	DM2 �C�R�������b�)�5C��+Q5X4���|�'\�+���x7>9y��XbhX�׈g�B���ņ"�d��ei����X&έr��Q!�UZ�@"���,R0IH�'�Q��U)�3U�Z�B&���l�0HJ!�m���C�P�:�=x��W�`�!8ԛ�y�d��HAN@t���u��R�1(n��!�B�3|���jĦ�G_X��T���ɀ�Gv5l9�&�B4w��G{�� F�f�!��E�&h��#S+X!b`b;2X\5I��;�I�F�~uˀ�U|#2\��K��t�(�k��G�L�\4��i��S���9h�
�дW9��7�0<OĤO���mˮ]qb�W9���g�(4�|�Gr͙���a"FƎ�c"�I�uF˒+��pK��X�X����G>o���s����G)o�$��#qb ��<^,{��9�M�� E�f�Zh��cޕH�㆒p}�J�^s��Bv�w��b�*G����d����rd�I7�d((�ʁ4#��C�*��'�� ����ў`(���T��
scQ��>��el�Ol`I��΁��Lev�<�;y(����φ[�� ��N{�ܓ�ʑ�:<�m�ۓ�y�%J�ʊ�c���;?�.@!�Mʁ�y��8ʓ�u�_��БoѲʷmƎ04�AӒ�$K�	a��[G�'��ђE[�7�6D�,\:��2k+!m�i�0-�_�<�"�!��牖OS��ae�3*��I���98h�c���j��Ma�,��C!pk&�R�����(��#M��jP�Fn؅J<�q�'�Ǝ
�d��}x1��beq�$�D��yRE�g�I�wl��JRM-�WK���Ri�0)� `�E�̨m\�*,�|�b9��6�81�>�֩�4N��Tt��5)�%k��4�Fm��c�EMWjX��k$����%k5�хV�d �/�k~j���%>�I-2���I�b��K��ѧ�剝�n4zU�6��8 ���_}�">��+̭/j���j��@�dpP����<��$T�ͺ�	���7I`�t�a�Ȫ^�Bd�դ�]n}�'=�'��dˬ~�M3+R�H�Ñ.���!0��<�&� �dq:7�B2z�� �p%�
���Xw�2K���p�A�2��6Pj�	��,��ՒE�����`g�=%��tP��&��lG?H�6�Q���OXAi`.�6!1qO�52j��X��� �͊�X�xp�"�i�J���JΌ�<y�Q�GX��
�#��y��D�R%�.$��Q�c�;(�F�@
C�R➠�)Z�J�v�"U��<	�Z�D���5(��%Buc�3�|�T*2�^� 	��$h�z"+��x�JD�/���
'��8}���J�Y��4���ը ������O4Ѓ�J��6�ƲST�Co؛Wq�|ZB�(P���A'|<�zkЗE(7��O6��ΐw/����
% ^�Zrb�;��=����
�զ��+T���
����V�rC����hO�)���ֶ8*:������j@;G�<��ߙF*����H)�&$��%�j�±�yk�J�bQ$	-h�aT�@�}1�Q��$��0=i� ʌ|3(T[7A��9,`a0�d���&8ZxY5E��,``2�t�N��1�u�OZy[1�i����RBL9z�̈�,���A��DZ��ډ*A��y��O��)�W&�Owr}����7x�[��<���ēr��y��'"6��g���6��1R�6|��g�k��-��!����d¥.���P�Ă	��֧uWE�0WJ�Y2�SQ�x0BböD��Q��]?L8̵�7 �"@L�&h�`�e6OfjK8G(dGz�!Nm��ܰ�ʆnH��q�*(������-k��7��κ@C�i�aA �	/)Y#oD-�`��J6D��0=a!i.n���9m�J���ӛ^�FLi��0�,#=�`��%���û�M��B� �>p[�(�$�.,�`�E�Qr~�`m*��&�Ssm	7S�r����3(Ӹ�mZ*�Փ�ĸu�RYq�e��i�	Sc�MIa͉�U��dȒ�&"u�#=�S�Չ_x�1��y^���,�Qyrϐ7 ���z#�ϓX��Ubqj�'�M� S�|/�O���q�0,2*AA.�6ou-Z��]��	�&�tX���#]t3�pI F�	��c��8��TB3��d�"J	h�	�������H�F���B�m�"�i��W;>�a¯ɱ��cH��}���t-�� ɓ�K�|̓���qF���3kÕL���� GZarB"Q�w�m�>���x��&��OBݺ���-C���#'.0� ��i��`�a[���R�R�3"�"�4l�0mi���:j|UHwnP��d�G~B8H��[fE4������D���d�%T����&��:SqPC��!��i(�~V�$�V��rP���ߠ&��c�'<��Ku�ʹv�R!hL\8RI;�눙���i�4$��0H�'�p�J!�l�a��i�}�lD3uDE6�4؉׋5�OX`��a�>�6�@�-�Wa�p��Lӧ^>$���_���{��,a.�W�ß$>��'�Ĉ�DDͅl,z `� ��(�i��Db�.em F��i{�
�6n(�7��)s9ʵ#C�ͺXofaGL ���Lr�ڭ��n6q��2���	��O��`���Z ���G*]:,�U� h�,n����v�z���R�<i�+��<��'�ω� �"^�d�Z���6	������5�O��Y�D�U��	X��,/�DRDZ��#h���P�A	/�&��J}���ɂ���2�J-3���f��Np!�ȴQ=���dF��)[C�ހ%�M���O��+�O-O~zdD�:u�.l�L��ox����Q	Q��d�S�,D�������qyS�S�w�� �fA��-n�o&�4ŒZ�g�H�(���݅z5`J�L�0��E�-xD�7���yB��];coT�(|f�p�� �OL��(�-�H!���0e�ި�s"O>��B��30�8���h�]Ȥ���"O*�J7֛\�P���	���*�"O�MHA�	����IOA�EQ'"O��q�G�H�m�"dQ:.Y��"O���d�	��x�6S�A}V9 �"O�) ��F'x�VA@;�f�xP"O\�e�F+uⲽ�� Y>fr�]"Ov���
)2(jEO�+;�� �"O��᠏SnN��@� �)�0�@�"O�IpOS�<� �٣ej�j((D"O|��B#������!X,k��L �"O��Ip$�2�*u��ٵX���B1"O{�Ɵ��� [_!��)�!Y�<D����U���Ƚ�x��˃g�<2&3�:PXD@����W��c�<��M�z���c��Y (�-x�l�{�<a$�������iV9)f.ݻ�H{�<!	<V�z�sƖ�����b�<!t#G6��杖 �FM+&�w�<�6/�
h����&W_� ���Fu�<�3I�r`|����N0�	2̙q�<�7��x�T�h4ACt=�*�j�<� 
����I*%�]�p���H�Qd"O��۳�#@�y��& ��"O�5����H�=)@�P�@��T�v"O�̲@BQ6��Q�s�Ą��k�"O��p�N�= a@�)�O�2�(�"O,������X�w,�T��2"O�����s����D��$��"O�}b3G��(@��c�(�ܤqg"ORl�2	�Y����2�Z���"�"O`��荨3���"r����"O<X���V	B�֤���R	O�RI�T"O d�Ga��S6Bm9�M�e���1�"O.rb� WzƝ
��	u��YX"ON1���=����1͖?�&�#�"Ov �
�yd���G�x.1��"Ol�D��2O}x���	�?w��Z�"O��rU�J�2�C G�Sc0�"O��Q�σ*�L�P���}V90"O0��P	�
�}���
:?zܡ�"O�P��w�T��gU&��$� "O�!ԪK��V)C�,�<|�"O�cҋ�&F�u!�Aĩ~o���2"O9����8_&���'~jl�#�"O��9U������7 ���b�0�"Orm���(
+�x�0/T8g�QY6"O�9� ��>�cE��Y��ms"O�2E��*?h��u�[2��D"O�`Z�N�	F��n�&�d�#�"O,0�֣S��(���;j�aq"O��!�-�D������z>v�js"ObM��E/y� c�ȡ]��A�t"O��`Ƙ�}|�:�E-B��}�"O� �"��&,�9�%��}�Iʳ"O�)��l�P�VD�M��)*�"O��k6��'�V1�����8XQ2"OzE�bh�������>#�` �U"O٪��e�-���0E���!"O���T��[`��	@����*�A"O~�X�b˻9徨�,�To2��"O�̹�%�(J!��K���*3‰"OH���6d�����v��U"OZ��K+@���"���\�Y�"O�L�Ǉ�tT��A7�T
@����D"O8+v�D:D	^�&��(>HiE"O�	�c�G�>;[!רԀ�jha2"O0�*m�*>���'ቜ[����u"O�ؑќG�����B��٘�"O@��̰v�I�Wh�;{�x�"O�=@��VB�DX�h�\�����"Oؐ�p@��'�=ڠ���j6"O0�����&�����0�x�a"O�ܐ��&d3Υ2Ʉ��8�$"O�p���T�w*�M���9Ǫ#"OD�"�,$P7�aX�&�Z�Q�C"O$�EH�T8���W%MZ�Ը#D"O�m�&S�_�ui��0�ȨYg"O ����:>d@��0��Ihp_� D{���^>2<my���?+�䐩
�	�!�Y'�G ��;���I*�!�Y�JvT��5�̿#Ě��W��!���R�H.2Q�H`��(R�� ��'�R�`���@H�9m�-2��Hˏ�d0��"��x]���N SI�h�"O4�hwhS�d�8����$/��3�'�ў꧙ا� �iZ�%z� 1&�!UCM��"ON=p �=6]��$6?3~�Ŝ>9�x�:"� ��}�0� =>,���xe��[���#L8uR�ڃ�lG{B�'��%���?����D��}�3��Dc�O̜P�c섘T�ty(�֩pVdub�'�����)&%��HÉ���w��'7l�Ձ��$*j<{����G:�0��'��,�eл��%jD7n�v���'b�	�աH�O�y��Y� j�'I�|�QD$"TR$��j^[�A��'�*8"e	��1Ǩ�):8`�'K��jg)_OZ���
�‐	�'d��8�Hџ�x[� 1[�b|��'J@(u��%�.œc� �~��lK
�'$�؂u��,_۾51���y-�@
�'���d�1K��!��;n
�(c�'n���#@�R���Je�׏f(�TI�'b�H�BE���e[��@�0�6��'!"[&��
gG�`�_�-bj	�'W��S���b���(s�\&����'�p�Xq�!~M�m�2,(qӦY�'D���V�X�#@]#>`5��'�0�ٳ�N�%��Q��Ѡ� �9	�'���iB f�J�3%�~�J��'���R�j}���%߈?�O�HF{��M�co*�����%�h "B���yb�X�&��Rr�&���jܨk&x˓��Ӻ3����+C�����BDe/"�;'���B�ɮR4��)��X�*��6�G+8����M��h�ㆃ�!��mj�&��<Q�D ��'���t ��86��L���ݺ�\	��(/D��z����8 ��h����Cф.D�����Y�O� 5��o�"Kv8���.D�r�i�0k���;֌V9pi��1D��j֤~j^�HP����5�C#D��Z�������ᤣ�q����ū#D�����а0��̡c�K@��r��"D�<��IU�x6�����
N���#O!��u�D��d�>E���#��@	&;D\��5k�!��DA��D ��mYA�K!sw!�dbI�I@&�ݳ.�ؠz�(_ayR�1W��)$�_!~'�]`2iЈG0BC��<r�ds�eG�0��Z���*q�㟨E{J?���32l�ހV���k(D�딶	�r�[�	<L_���d!�h�<1éN7iGR��4�S�o��e��h�<!e��6"��Q�H��\�j4Kbm�b�<�CN�<43D}i��״m5�(3��Z�$4�S�'/�<)K����!�nĹ�#�K�Y��'�&�����9���!d�Uv�L���4ZD��ҭND�<�!�Y�y��_��p8��í�-�VJ���`�<9P�Q?Bv�As0�K"��-hC�]�<�ģ	�.�cS�G '� �c�Z�<��ďU�.P��M7#��zu��[�<Q� �&��<��Lq�ȥ(�.Y�<I5F�
p��l��I�~��E�R�<�̐�q�NU!g��3�A#c�G�<� ҶDҗ(!�جh�$�5TbB�	��\��D�ɤ*7���#/S?9��C�I�|o�;&AS�Sb�\���{��C��&d�$8�#ۦ1�������"<l~C�ɗ R|�PD]U��<(� W�+�lC�)� 
�HU�!��1� �`����"O8�H���\<B㢇 cȬ`��"Ot���D �8`�����ab��R"O UR�*Ҵ�C�K �$X�d�	u�Ob�ARQ�ZI���C�n�J��'=�<��l�1�R�8f%��l��P�'��9�t�CC�~10WBD�c^�u`�'��aABG*+&����e�<�y�'���NŀR�"0��,S(W\�r���'�X���2�R�� �Q�&^z�
�'�F�3ɐ�]ԑ�F"[�#�M����4�S�$S=I�A�A�ޜ7!dt���y���E�j�3���6���`�뉏���4?yI<�����Ibi 6��zd�틒k�!*!�S�>�!"I'NQ����/:k!�$ڏ,�tb�E<@c�}����Ig!� )0:��B�M�\F*��K%�!��P�p����J��ꅹ��sf!�dŢ�栐"�UY�bg�©f!�]�^�d��3�$-&��	�`ɣ<X�IH������S�U�jLz��r����-*D�$�t���>d���ܮb+�1A�d#D��V/L�4j�g�%=�$;��?��0|����	�`��"ڢH���X�"�A�<�ˍ�3�nd�S�^�����^f�<���di~�a�B��LatE��Bd�<A��@�^ꆠ�g`�%;G�IB7F����x��k����Ǘ:>�5�BN���y�L9A�B�hF��0?� �Ņ��y��L�8�v� A$�>=�!8�'��(O��=��ڟ�򵍇�7�8 ��ᘼV��ᐦ�g�fC�I(.~���CfJ�^���6]X"?ш�iE%?��tz�e�x�ƆȎe"!򤏓x�!��Zv��`��R�5����(O?��WI �CZ
݋K
��:qrÄ>D��QW��P�d ���}I)uㆵo�qO����x(�p��-�:w�0Ȗ�Kš��	)Z�Q(� a�ö�DnC�f��+�Ŝ�-�����X :@���F{J?�Y�*�� �� "��ȤUC|�b��;D�� 0�NKht�z5G	�XN�<��,D�"vl�PŰ�[DDD�&<d�X&D�`�Į�7���bA�i(̠"�#D�l�R�ܣ6���*��޳33�9)�4D�<K�!��g\v�*Rl\��y��4D���Bk@'�0�h�HFSX�9���/D�t 7��5!ܶUy�EG�X͆�[3�,D�HFA��i��d��4Aj2��&D�t:���.�6��d:���$D��A��תV��3���
:W$��@J-D�B�S�)�\���G�\#�M��,D�H�EW��	tiG_� � F�?D�4;�IF�2`�t�d�ƴR��k�D<D��g���&:i��5J����C�-D����c\;�(���ឦln�\#�(1D����M�9k�Z��ai�tQ�u�.D��;�ǆ��8t�E�w��*�C?D�l���c���)�aKOd�: f>D��b��KE�8�t�\2)�jً�.=D��r��"�F C �G���p��<D�ت��-h��qB���.R��C%�-D��h��O�
MN�h%��0���(D�H���*�fTJƃ;i�vD��(D� �g9 ]��օ�7�\P8P�'D�� X��.קr��u"3���@4�w"O^��X�i�D��6m���q"O�A�Wm� ]c�,`�a�$o�\�"O�mȵÖ#f�s֢���S�"O��ZGΓE����&ጅ(��hx"Op��"�1i�E��M\��h�"O���/V�i��K�Mͼٸ�9�*O��8s�]�M���3*�2�(��	�'W
9��J߿q�iS"�Ai !��'���,lV���.P�0n�yr���J}���ТI-cvȠa�E��yOæh�0<��g�H���j��yB
A;D��II�OJ�����S� �yb&�|Jy:�'ֈ�H2���yBZ�r���Yf����iX��@�ym�4]�j	ɢ�
,=��� l[ �y���)N#~�ȵiKbE:���5�y��Y2h(�L��gS�PLt� ���yd՞�|y9g���~L����$O��yB������a�MLL���#��yr��mr4�p���\|���.��y҃K�u0�ä�\����@��y$�S�v���ɅP�����yRIR�D&<�m�X�Ԛw���y��� J>	P�Y�Uj
�!-A��y"���tA!!�L[�IgV��y"\6�x]B�j[3��x��M;�y�ט2�jeU��u4֙a hW��y�d��C�~8� ��ty����Z!�y�#�GPu[���2i1(� %���y"�A�	�h-��EK�Tz\`Hc��y"E;�;��6H5�)��ϳ�y�%�ܒ�O�?8l8�U���yRlS� Y��Q��_�f��$�G/�yr��2|�Y3c��[�D,��M1�yR�4pv��ш�P��D
#�y�♙?34)#s��=*�� ��
�y!\��R�IΨ<h���C��y��[V|%�w��3A��Z��G�y��,x9I�BM�@���駅
��y"A�-!W���<�80����y�	˪>:�XꀆY�g�6\82�H��yR`">�B��#�`t\XV���y�B�]Dj��3�_'��p;CF �y��	�^$#�A���� 	�$�y2��9�$j��)�������y��=
�x(Af�	�G\��JG �y�A)@�X�ga�2�*��v �	�y�/ ��R���L�	����,D��yfG��1���#�tZƊ'�y���!hMJ}
��ڑJ�5���y�"�B��M�V���T�D�O��yR�D��x�ڦl��)^JQC���yR�c�f]���/2݊� ���'�yr�_�;�ʸ�f'ՠ$XRq������y��7ch��pǧM*-x�`�k��y��i �RS�(X�9���?�y��$\9pA��(�AÔ��6�y�NCyp|bf�S�!�ĸZE�5�y�jB�y>blK���O��Bf��:�yB��)H���bW�I	|�����y��ϥ~���bā�^���rd�D��yrg�(-�6 K.�Fa�4��y�GK+)^����ڇ+6;��K0�y
� 0pذO�p�ܨ���Jnrh;G"O@�	V�X�O~�RbT 1d^�R"O��P$��E�x(��J;Eʡ�$"O�Jakpv<��3�I�"O�3 � �X0J�hW�@&��:p"O4u�7�L5u͔�sOK�bP���"Ofѱ�'�$Z��ȂA�F#s�b	�"O�]@6�Z,.�Ç��\��0�"O@�p�ݲFGغ�o���=�D"OHmKeF�2T8ɨt�G�<��"On c�!��X�d�I�R:d܊�"O<�PcL�$V�~x(p�W�O��%
�"O�i��@�G���ЦR�3��Ea"O�"��h��e�x��D �"Oh%sA��0O`N(@bD��Y~�d�"O�<��:���F�g��i�$"O�
�S�R Q�E�3C�����"O���6i�GhL�6@��V-|�K�"O��G�E��|0G�ζPs���"OB�ǩ�n����ֱ$c0%X�"O`5���j^�@V;��Y��"O�m��LW
,ax�� ڂ)����"O\耂ι*�ʴ:��ӟ�� �C"OJ�kR@J(1#�IQ�$%U�l�s"OJe��X7+�Ջ�f�=V��w"O�+wd��PvN1k䆎��Ց�"O<my7���,�p��3&�:9Ei"OJ4�%hN�b^���%��e���F"Ob�z�,U�Wt`�����S��P��"O(|S6�	;|ض}��k#i�$�r�"O6UP��Q<�1����3�2�#�"O���S]_���*������"O�L�BF� .V�(P)��t���"O|�;��>cΘ���� |`�W"ONE�!h�<~ p�&��(��HJu"O��@�*�#-* �5��t�A�"Oz�2I�%`�x�D�r��ɪ "O��Əƺn�d�e��,X�NT{d"O�<�0���p�8@FA�6|�E�"O]B�حn���Ȱ3*��	Ys"OT5����>i �����l�"O�H�p�ֲ(�qqaD�*��ԂT"O�q$�M�R�v�z��,M��:s"O.����o�ɡ�lļ@����e"Ox�kb ��(����b,�!e��3�"O�yC$Z�S���0��J~DP��"O� P�+�/�u��˅�@]���"O���o�IX��g�^8@0b"O-J�h�94�R��Cʏ��.�"O�=�" ^��5�E��.����"O"���h@�FJj���GU�1�mC�"OX����6n;��0�e��>T�g"O`Ia&��9~jEы��V����"O	PB��=ulq�����k�"O�is�g��W-�1�4J�^F���c"O�]�.G8b��C).O�q�"O�q��!M b�X0�֊L��h���"O��Ғ��S)���� �|��Q"O ���1z����.@6�¥*u"O �S����ȇn��9Ol=�1"O�S��.(z� U䊝\?.��g"OF�4���:PZ\X��"y�L�"O���猕�/L�X��l.\��"O.�IA93{L)`d�'$"��A"O� ���w"T+Y�ҔJ�"��
.8 �"O��iSeH*o��PA��=�d��"O�qCƃ ��u�`�Ǚz�|!�"O(4R5Ďb@Z��éy����"O��{3.P9C����m0��"O�u�4i<����a�Q�d�f���"O�1c�(��i2Z�������g"Op�i�B�X�qWc�6)���3"O�d#�B���9�G�]�u�L�$"O�YRanȿ-�8�C0�ʊX��"O X��!ȍ4wbej��[:A?
���"O0�� K��$�Ԙ	2�#?�h�'"O����^�c��E��.V��E�V"OLЙRØ��|�p��;��ɛ�"O�%c�g��x��A+蟚X��D#F"O�a��ò<�	��	\[���"O�@[!�L.{;<��Ƨ��]G�h"OX����2<vޑJf�3~�)*W"O(��w��|�98��ʔs�����"O���P�̢6�h��!�'���E"O���'��(p�����o��#���"O,Q�Ã.��9��-W�;���"Ovj�)�V�" /�1v�T'"O�qZ A�?�1b�lإ;-�4�"O�]:���1��C� )J	a""O�Tk W��e�0cA2��:U"O @K�@5G��}(�� G�xq��"O&IPd&I�G���
�b�d�ЬJt"O�|��'� |H�"S�SҎ�"O�x�U@@:uMX�����AZ���f"O�mQ�L'��R
L�n�R<�b"O����(��"��@�IԻ6���R�"OXMs�l��4�e�J=i�"O~�e�,��q�4h�.nǢuQ�"O��blJ7-n�p�GL{P���2"O�q�gm��T#��w'ǾVo�к�"O�в��oȰ���:iV�"O��6���m*�xJ�Z-b�0A@"Or�����9WEؤE��u"O.}���L���V�_�w��S"O���!�V �	���@�c��}sC"O,L
&fW|�&l����;v���"O��ړ9)�l`_�qYT"OP\�6��Y�6��%)½t�ո""O�4�V!H1r��ņߩU��8g"OZ��t��*���D�܌��lr`"O<���؃	�
8�&�S��N�B�I�b�,�
5�6C�=Ѳ�A�l(�C�I�b*@�o� ;V��Q�C�Po@C�;/�ȓ�*S~ܒЁ%
VxUC�7���`��c�8p� ��;9�RB䉸1��}�d��a��t��-B�I0i��]��N��>Q�Ը��{9�B�ɣ=�8;�W��Dِw,�P��B�ɨ}j1���6O�\� �cL$iH�C�Ʌ&�N�0ǩ�)B�5
o��C䉭OشA�u	�.�� �00[*�C�Ʉbg�2b'p٫��2P��C䉖)�|�s���b=�,� H�j�C�I�&���p C�
�n1Є��Qk<C䉞x` �0mI�2_( �S�,�C�4��A$j�m�B;d��E�B�	�B��a��^�L�N�����0��C�ə���٠��2Hr�jƻzsB�)� h� �\<^ql�g��[�֜CQ"O�I A �V�2���<|6�Er7"OpzҪ
�?޸EA3��rx�`��"OiH���1X �/��`�$p"O&���*fe���u�ЊRE�ije"OL��W)֗Y1�����ӆ��)��"O.���`4���x���j���:�"OdI��GF�Ո����N���t"O���s���z1���d�hlK�"Od�؂گT�6h9s)
?b,�0"O���v���N�bd�d	İ(�}��"O栀!n�2�<��aE�J�n��@"O�)��	��B�PB��s�`��"O�C�Jӆ]�i�Dc��h.��p"O�D�᧕�!d6�0h�0���PQ"OP����X^�3�;��ab!"O�h��S�|9�f�)vp���"O����C9Ty��8���c�"O,9As��4l��J�n��)��"O�Ր��V#�*��s�J�a�j��r"O�q��IT.:5D�2��۳��!q"OV��I��;Wn���N��t"O��� ��=7F�ybM�H�C"O��2кyU��@m���̙S"O����00�zYT��*kx��"O�}i'�˚J�b��PB�v��Р"O*�����67nx����%�x5"OR�;G`�;@�!x����y��l��"O �Q���/F�̪�.X�9��� "O<:/�Q7i�N��y��mڙi�!�d:!���"��*��c��!�D�1=� !�R�ڷx"J��Q��w�!�0Pt��[�%�U��P5i�!��ܐk��Z5�аp�4E3��0%�!�d�޺���?H8�zvo�+�!�� L�ܼ��(7�(�7��Q!���`v�:V�57%X�j hW�S!�P�~�3�^���fɟL�!��N�2�p��`&�$BVA�R��9?N!�dr6vyd���Pe�e�BW!�$��^�*$��Y�L��0���J!�
B�@1�u�&mó��A�*C�I�"��G�Ȑt4��A*�%?G�C�	�+��U�n�&��T���	:�:B�ɯhp>\B�A�"��0	U$�%j�PC�I�lٵ�Ɛ0j���0���f@�B䉅x���q��7�T�:5KŕLgB�I�r�(8��,u����c��Q�vh��H�>ș�C�i��� 2��;%����ȓ6�	�Ϗ�%���'h3\(؇ȓy�\���Ď!�125*BM�,��^��S��$��q��K3l�=��R�\�'��re��YG�P�ͅ�V���q1�ƺe=h�1�F3��фȓ���@�����0�ջy�`̈́�,�V��g18b�-�wCς�`���� ӵ"��l[l)
5$�7]�����oA&qpR��-�f��$=!�܆ȓ4㤄�w%��(������;H���0f�ʭ�䕣���j�4��4��\A�$tƢ9�rfN�!�фȓr�HayZ�&��sRֽP�8��p��+c�$A�p�J�O�5L��(�ȓ|��C�0u! ٚ2ɇ�Mzх�S�? $8�=�TX�DW-"NJq"O��"�,�P�E���Hl�ӂ"O��!4Đ�Rym�@�ڵ��1D��(��T�g~}�d�+i����u�+D��W'�&����dL�3�(A'(D�`��H� 
�E���J,XR�0Վ'D�P�qh�q@<��F���r�L4 U�&D� ��E�Ryt���i�+a4H�h��?D���c@Վd5,H�E���+�( D�,��ٲjS`ؐ��_'5\i$�3D��+� 3y�hJ�dѷ`{�!��0D�h{"��`�V����	N -`�!D���,�Q����� ��<�8��:D�$��C�'3N8��bS-\���B�3D����n'���`�P�W�¤y��1D��I�OT'Oh�i��(Πl 	k��*D��ѐ�N�䄚��('�<9s)(D��hP)7�� ' H<�@St;D�X3�?b\e#���?L=�4�W:D��I6Ȝ��0�A�@8$�n*�*9D�piEm��~��RW��![L2�f8D���F�idK�H+
_>��"5D�Hk�ɬM���P�&�R��X�%2D��Y�8�h�+�`;��9���.D��)��l8Ĭ���]�H�ӎ7D�0��m� 1���ơN�<f*8�e�5D�<��FD,+�ܘ梇�K彩���>D�� e�R�=����-GF�@��<D�p���DKlPc�MҌXB^Iq��8D�@C5�=���Q�[29��yУ<D��+#�;X���C���VOё�:D��K ���| \;uE[�cr�|��:D���5H�*C%�+���N��#�N6D�lb�Dګ|���"d�,�L�V�2D����ı�z��&/�`�hqE/D��)�n�' !�@�%�K��N�S��.D��!�HQ&o��q����mx!.,D�p����/;a9�F�����"*D�@���A���"I#TRĹ���'D�8Gln�LC0��.=����'D��haĘ��&�:�!�	>kzQ� j0D�Pp��>�)w�^}�H5��".D�`�#E�(t�� �I�M��1WD>D�t ��ԅ:�L�Y�%� n!��D)=D�$�U�J[w43���4��xYÅ=D���7jԸ���q� F�	�~�!&�<D��"@
V
�D3�kH���&D���Q�!���	�� �-/��b&D��y��Ävu,0�&�*O�!S�9T��x�ψ�Ђ &#Ы\�\�B"O*�1��A%���bc��*�  ��"Of1K�a�xM��SfO`�\�Y6"O�E�GL�
0��]i��������"O ј%"N� ���*Q���G˴�	�"O�ݨ�ޮo��Ic)��f�и�"O�tkփ�$v�`�(`�ˁ+�C�"O���􂈢=*x`"���n�X"&"Oe�u��~�j��W���8�ec�"O-�0�)r8h�r�/��Y�2T��"O:��5k�3Ff��6�1 <Z"O�8��؝G�p��I����"O�i3 kàA�� 7-E$$�����"Oz �7�֪��aP�-��Vl؇"OJ����ۍ��Q��S�Y`8�a"O� ~d�wOB�+�0h�r�
Ox`�"O����T�6�J@�s掜w1d��"O��R�+��&H4U���s��@��"O`���m_�2b<�s��;�ҙ��"O�Q$&
RxP�+c#� T"O�!� �̕%�����A�R�)�"O��2��#�r|�ǈJ�	����"OHH�Q�� %�v��$��P2l;�"O�C�b�����?K�`�G"O0Q��Y	x����� j�ų�"O��g�(�y�"��tZ dC"O�u��D6��Pk�ˑ(%db�qD"O�"�A܎3
̺e*υFYlPx�"Of�a1��5<L81��ήuBbt�"On����
+v���@%/)�|ZW"O�XQ��ؤj�*��#IU�>�lI�"O���Fŗ5zPqHQh�a�!8@"O��;@�[�G���'T�k%y��"Oŉ��R�\��eIs��w;�41"O�tTn�QIb���Q&UI"�)�"O�X�BEE9eW0[S�	mCށ9�"O@�P
͢!�6���ޤX?Dl9�"O�	pf����e� e�n�*"O�J"�	8­��ʟ+�Rh��*O.�	b���k[��uĘ<3���`�'M�IE�- �
y�ub�0-Rҽ:�'g������8~�Adk(���k
�'�th�%�ҿw2�N��I��U�	�'l���C����p��+E�Zl�	�'����d�|n����.ϖ�)�'��yf��`���"�\,���1
�'ބh!�G�B�=P�'��ޑ��'����d�T�
7�4�P�=`��'X҈�p(�?<��k��W�a�R�j�'Ǽ�0��:/�����ɏ'_�tH�'В�:ֆ��8��זez ٻ	�'�j�	S�J5�a
�nD�r�Z�`	�'���%� $��9	�g���$�1	�'+$<� +P���nG��6���'����q��J؂��j�
�'���Y�&��/-$ � /���:��	�'<=�E�
4�`�2㧐�L�(%��UK���č_`�
��E"86-���a�3��}�&�BT�͒N�q���E��D<ZA~�
D!UM|Ԭ��LN ��X4�R�r4�G6��m�ȓZy���B
1�$���6m��`�ȓ�᫳ Ќe�Hi���ԱW�n��4z�=�d��!��%�#AJ�u�E�ȓ�~���g�k�Qf��^4@ل���
�L٤KF���QeB�
A�ȓ~ݑ2�F48�|��Q��O��m��fʐ�F�3���a�?yS�<�ȓ.�j�`�ؕ*'�<�*_7�����K�1+ �F!lP3q(�AS�	��ar�h�GֻP�@���)�:iఁ�ȓz�#��E�( �=�a��1;���8aH����ɦzc��t/������ȓ8j�ce��O7��J�d�{q�ȓP�q�e.�*Fp
��em�P��!h| 9���=/���Vo^&r6<Ņȓu\6�Cr��"Zdʹ3p
�P�d�ȓQ�|}  ���p�S�J�xV������#�V 
D��L�
N��=��S�? Йk�eQ� �ԁ�KC�^�r�93"Oʡ��i��X���\�JCh�S�"O|+�S�\��6#Z�g;��K&"O�y��D�>∰�^�B,�"O�0ic��7Z$��m�"X�z���"O�e'��:|g$�����pc��3"O�(I�7�} ���.$V�U2�"O��� ���'({En0fTɀ"O�t
���E��c�֦]pH�"O
�9���9�"ع�N���JY-�!�Ě..t<��� �2��#��Fs!�DկS��)��g
3�$P�XE�!�՞D6>�������!K��(Y!�DS�<�����;T�(�!S	xQ!�D1FK��{q���΋0 �B�	5"+^) Fd�5��\z����ni�C�	P��!�S������ p	zC�	�T��:��*���C��#sB��-Nۚ�vƄ�Q����L�.L�C䉛5�% ����Q�oA2A�bB��3^ p�PG�N�~is���"�RB�	�
�@�J�k�5K�l,p�u
2"O��ڄA�ʠ�޿
^�!�W�@�<B,�L�Q���9����c$A�<�t�4$Ġ#��(ֈ)���z�<�h֎(>��L�5{���'�w�<I�E�#�t���j�HY!��Gt�<�I�.^1�L�b∐v��a��%Xm�<Y��V
5jѻ�˟�
7I�(r�C�I"S�D4a�C�# C�P�SB�I��0M`�<vF6���럽E�C�	>=��\
�-��(hx�"^#{��C�	�J�<���_�DX��!w��C�I�G$y�׮Q�yN܅i��RDa�C�	�8�X,�qd��+f��&,� I;NB��8��[�M�
G��5J'��!�vB�� U?D�H�/�;'1�%�R�X�L�B�	.Tt,yc_$�m��D�c��C䉻!�*�H$(�%��s�NUL�B�I+518��.E'd�|��eL�*T�B�IJ�`�I0$[�[Y���g
;�B��/�PiCe�����H�Ao<C�/	�I��">=�e���Z�+qzC�I�7�q�]R�qC�φ
_����"O�`	TG��D� �yQd� l��H�"O:��BF%>�ڝ
��@&|c�-�""O�����/x�L3��1I�p�"O�E�ԯO�q-�˥-\�h�*-��"OXm`����d� �2c��x�:7�8D��!b6=�%��+V�MV��l)D���c�S� VԐx#XA F�Q@�4D����	���n���T� ͛E�2D�`����'2XD��H����R�0D��!D�:��ԙ5��%2����E/D�ly�ĩY�
��J%@0d��D8D�D��+ӿ0F�{�H�d;,m�D8D�h���֛c,����n�f0a%�;D��w,8hm�j�
��|0`sE�?D�!��S�\�����N�L�X�!9D��gl�"�>�[�R� ����<D�T���IuU�q��A��1�1O9D� @a.@�9 9T�Q��ј��1D�T0�j�e�D�w�R|{ȕ9R�-D��0��F��({��[$D
�-��1D�� (�y� ��0Ě ���-oPqcQ"O` G���T��`���B��MZp"Oܑ�t�2<i���"�ژ��"O��D��5m�T\�mK�E��@b "O6��cL�/��ܛRƍ$�N"O��ҷ@�
�*!+�*M*~����"O����dؚEL�\c��ӭ��u�u"O�*b�'*�$4l�;�����"O�%� f�9�9�l�%p�Ѹ"O`�ykM<��(�/>c�mY!"ON�6h��R�N��q�aV�]� "O�	qT�:}(�����X�U��"O= �I��.���D1`K���"ON��g��\�ph��mBPC�}IT"O�B��3W���2��"k3�
"O���Q�$�=X� �GRo!���0j ���\;h����n!�Ņ3�\�#���~#l�u`ȌoT!��U�,��(@#ɏA����lH!� �4l��L���d]H�Kd2!�d�Xs���S���^�h5��'!��>!Ta�Шֳ�H�3�B�"!��K8=#���%��FЀ��3p�!��hD�P����H����Z!�!�$.L��EёML)F!�Wj��A�!��6�p�o��@��ۇ,4!�4IX>�qHεh����ҌN(!�$����r��Z�5�њ��64'!���Ȏ#!TǞ�HED�6?!�d�NS0dɅ5f�z]X�Z>@�!��D�g&$�x��X�<9!g+�5�!�$ߔb�T�
�(�`�ɉ��T� D!�D���7ϳ�&�,@�,$9	�'��s�n��/��h��M�<)��'k�I!��	P�^=��-�!q	Ꙣ�'�Ew�K�<�����5?�MS�'}B)z��O�hP��N�.''�y8�'^�b�Jǯ��ܚpOL�ТT��'t=���� ��E��&Q����'h^�d��s��H��$K�t���'��T���V�o窕PQ�^3q����'�^���]�J�x+�:d.�I��'�@���;�d���Kc���X�'fp���)X*g�-K�M</��	�'��F��F����Y�'@� ��'o��0��
Rg@d�,D�t�f���'��X�ҙ5l���Q��Uv��'ĶL�5M��y�����ǀO����'�Lh`�UCur4A%][�`@�'��C֣]��L�c��	>&��X��'�r�b0��	�(`I��Ȗg���'Hl�4�X:x;g
	��X�	�'�A��)�$Wb������ �f8��'"1P"�4J��5�
Y��'q��c2�*�0@#ԯٻ.=�<9�'�~��椅~��t�G�$? �!�'<���O�(k=�U��ꑟ6�'�()a6J��(y~�@��N��'�4X@:80@�өp�DQ�'zZ �4�ʤ:A�U`�A�k[��'^�����
t�|�� ,�84�^���'��,�C�)M�=)�n72u��
�'��\J4���o��+��B|�b��	�'���� ��_<�|�%䉹"Z�-b
��� bm{P�,!�d-���D0�E*�"O\�"��U/�6Q��ʑ�fDpX��'�F�ڳF��be��j���ze�'�����JU�ܸ$ဩ�RU��'�b����D�3��4H��Ǫ<�@�'� ��` Q8Ҵ���٢L�|0	�'�t0�@ A�8@*Tz��$@	�'e�xI �*X�����'K;]F�DX�'�,P�N~2���M(_趬�ȓP��x��C���Ƙ�5�� iK��Q�j��~"ĺ� Qv�ȓ7!�Y�&Ǹ&n���#l��0c"\��S@.b�ʀ_�2�#��"��i��g��q�b�
r�85�b�A$?���r�@9wC�{����egXe���f�j����*
Ƣ�	�\�(ڞ�ȓ�< %蟔|$�LA�F�p�i�ȓ����%���6)ġ�Bg�E�<��0I*�锋A�#��&�'X�Ԅȓ
5����?X�zE��#
��8����L9q��J�D,2�-��l7-�ȓAc��)���G�<�)T��B���7
�i@�%����g�F�������t薁�7��m�qL�#�r=�ȓ8ءŦ�*!N IgA��K U��x]�$q3���q������ͪ��ȓ=��)Kǌ;�����B� ��Մ���Z �̼=�v�2�@:Z��m���Ɛy��ÙG*D@r��&9�ȓ��Y����S�#G$ۢ+��D��t��&��M�*�[ЀH -�̡��lavT�g�ΰs"0�Bf�^��q�ȓ?�(	��܌g��衷e�@����ȓNB:�1q͈79b�@��O5�PP��+�L���4/��!�f�'=+p�ȓD�H�c�K�5&��g�]�ID���!U�p�C_k�n�� M-�ن�q��`c�Z����c,�x�t��ȓ84��������@rl�3)avu�ȓ1���s�ع"��p�g�2=+�8��hm<�E��#` P��a/i��܅ȓ*�@,�!-!c�tÂE�3^���ȓ>u
H�$�Ġes#�� /c�~��ȓM�|aע�h��J# ��R��,�ȓmf����Eܽ~�>�� �	�3��L�ȓ9�3�ğ�����Э^��d�ȓ�
��5��|��P���٣,㆜�ȓNޕx��� �r@��&_:G�I���T5 �8)^Dq��
R� ����ȓ5j| ���3N^�R���IӸ��ȓ,�4}(נ��I�t�ѩV#(E�x�ȓ-hY�%�֔ajP#�Kk�-���v��5���R ar�A��8��"OF J��G19�b����T^>px�"O"%� Er�;B��+$&�1"O���%��<z��죧,�?Z,���"O"�h�kZ�Q#�Y�Ъ��-1b"O-��I�Lȁ �.O:�T��"O�$����@V4F��Z��'"Ob8�!���5�V����˻*�ya"OZ ���I�%z�а�l�#2��Z�"O�����C�Įy	�,�r�L �$"O��[���vv�)S��+*��aIU"O�����%
6Y�4�E!%H.#�"O� �lrŬQ�8�<��1��%���"Ov�r��-��X�'�!N�F���"O���5�7D�!1c�F�-�ir"O��ŔY�v�a���O�x99�"Ot(�N�����3���%�"OZ����)H|��.ؐYp���P"OFCU��;{���@�Γyn���r"O�l���L*���R�Vj�@�"O�c�oǨuc~���<;Lz=��"O����.{�홀��4T�}(�"OԬh�KʩbN�y�B	��
(�"O(4�w�`���
gL3�����"Ot�Br���os��@4fҥC���3Q"O���(M	�hi���X	_�p�"O��;��a���h� F��I��"O� c F> ���ńA
ze�u"OF!A�_,Z�dإ�@�%Ld���"O��Q��ȼܡ���P���Q"OЄ�#D�w:\�s$�:{/s"O �s��r.�����v'�1��"O�(���)?7X�QP"F-o�x��"O�]@P��1��́�`ŕs�<�f"Obّ�OT�6;8��NN������"O2aC�c�Y���\��X��"OP���!{��B���/��92"OX���).�,�c� ��Se �"Oּ"7	��"|�r�eK;[�3c"OҘ(DlK�H|�Ԅ��k�
h��"O��㷫�|��1��$z�0�c"O��Cd �ajR�zp#Ѧ5��RU"O�X���	�i%:�X�!�
���6"O8�R�-E�%�8A�A�N���0"O�I�c��(!Nv�x�_$rn\ 8�"O�J�F��\)\�HtLL'T�$�Q"O�=�/'F�&����{�b2�"O"�Hs.�wz2�R��'��0�"O:)�-��qLd�!��X`�p��"O�t�F$�"Ic�ن �C�"Oʑ�2fqkF1��N��V���"O\y�7m^�\0<9귍�Cڒ-k"Ol�Dd�a�)�֋�>�D�S"OԑЩАh�D���S.[�dK�"O*�ZSo��x�V�կЌ(?Pi��"O``Cd�\�I��i�D���j-<��G"ODM�Pf��kS>���<<����"O�Qg��#=yp��ԙ:�d�@"O�lR�,D�^�yK篛-q	�"O9ɂ�W,��5,��[<l�c"O�,��mM�\/Xl��հlQ����"O �bae^�f�&-��i�%G|��"O|�6nH�`H�u���,:�{�"O�� ���8��+�jZ�Q2�ae"O<���"O�]�����CV^�E�0"Oha ȝ$K}� �⍒,J��-c�"O��vCB���u!��=sE!�d��4귬G�j����' +r�!�A�I��h �Aɸ,\ |�D�4;l!�$�k��Ƀ�M�?PT����Bj!�dN1<� -��# �e���j�b!�dϷ6i�M��oKgpx� �ٙ8�!�䅕/�0�c�H,V<z��W�A	t�!��(gH��F�>rW�)��C\�p�!�Dva� ��OE�H��ډQ�!�dP�7LJ� 7L ��Qb"B� �!��  �Z�*	.#}�mZ�g6�!�"O�� D�0~���I��D6n��K"O|+�B��k<�4��Ţ\�"O�� `��f�^0[����ߜ<��"O��cϟ$Fj����q3A"O�	�&Q�"X���:4�l-�g"O�-�߷s\�a�bJF1X��D�%"O��o�.����6C� BZ���"OT@��-��X�ZXs�pEf(�3"O� ;W�ėK=���夁�N?xI@a"O&�����}��MA@!M:PJ���"OЙjD�B�Ժ��JP���V"O8���H�pc���&�FsB��4"O`�0���n�!�E�J��|1��"O6�@ć�qQ���0��>*����"OpACCJ�,�:���*fv�!"Op�@Z.6�l9%)��t�b`"O�h�QL��o�����'�;X��Q"O$`�A%A6�A���r�J��"O���G$b��a�+�F�#�"O��P�ԇn�R ��dN5CSr�C"O��`�	��k> ���m�3U�d� �"O4�hȂ�HFL	u�A�Ju��"O���F��7~F6�C���]s*��W"OH�1$�/$<<c�!�C�0@�5"OL*j�2�~�I���h��,;b"O�(ʧ+P�8�N�!�H70���C"O�HT��l>��cu`�)}4�c�"O��k�+��q�XT�����r|�w"Oz�;1��YF5!�Ģt"ONlX�(�1e'Pi�UϏtA2@:D"O�HrO�t�b����lV�UG"O�1��G�R��t���Q�j>��g"O"٠�6�D�����W7F�2&"O�	q�,��s]����U,L(�0"O����ċ f�\�0pE_.tT��"On4��D�b0�򗨝� "�A�"OZ�0C�j�`XafI�%T(k�"O01�EAQ5BisABH�^��b"Ot#��[4!�9�TOȽ��"O�Up�/�2Q�����y3. �"Ox��P�L5`�
5�3k[�h���'"O(�aV�#�xU��ڃ�q��"O��S��?Fh1a��u�"O(��Ņ��$��i�e�P>8���"O>��H��I����G$]0�HC"O ��is'�i@Ŋ$UL��"Oh�J��8%`�B#P&���"O��ț/Ьu�w��S� �
�"Oj�sC/��AC�x��`>�*<2b"O(��K�NȴY�i
2�"�!"O��p�/�I���لC�I�F]I�"O��1҆E']�*m���Ѓ>ΌH��"OJ	��Y�j�i�&NE.`窩��"O̚�IF�Ҝ�C�'1�h�i"O����m&]NXˡ*�����"OR���(G�acf�ȉe���#d"OJ��Β;Ԙ�F�D��=QD"O$X��E�#�����B�5fF]+�"OfԻǅ]�X�x�� �];p^��#"O���0柭<&p���2�J"�"Oe;�a{!�'	 |L>8"�m^F�!��Z���1蒏B-���,R!��g�¥XAMo��("#L[X!�� P!ӆ��5\�$���ߜ(S���"O T��=y3��v+0RI��y�"OX�d���k�J-�jO0t0z!�"O0�����eX��*����!#�"OH����,sa"�v�� s�޼��"OF�K�Pq�L\�Uˍ+*�,��"OL%5E]�L8�Y��ɂ� �"O.���L7:<��{���+=ΐ�A"O�"�M�*E�l�F�	;�mȔ"O\�S���2C��33�T+t��@��"O�]�Ui�!/��u�B�F�D�A�"O H(S��[��"����r#C"O-#�mQlw�Z�B��(,��"O���.P^j`��#�}��"O�%{ĬH��q)��S�P��"O�� �\�$~b\�m��i�n�!"OpP�r.G f���p[>�^���"O�!�C+������QZ��s "O�����Ɖ%�މ bVv���"O4	E�X�z�<Ĉ֡C=kD�%z"O^�1s��5Z�h�֥Q4z*dT��"O0��v���y�-!&�u�V"Oh�QC(�$ة�e���~�`"O�8!�� î�S'��#G1z)#�"Of0�j�
0(Ä��(~,�QB"O��2��1�
�`�A��1����"O(s�D��J�\@��oR�&\��)�"O��r��O�2pHsAܝb:N���"O��aQ��5P��� [U"���"O�)ItW�I1�m�Ư:o) q"O:��W``^��c�Nڳz��g"OP��W"N�:D�#��3
��["OvX!4	�Q@�Y`L�7`JIi�"O�J�ۍK/v�a M�*yb����"O.�#�/ R]hZ�� };6DI�"O��e�/��z��N�CώMK�"OP9Ƭ���vt���ԫ<���s"O͒s��%VX�v)άQr
��"O��`�hΘ�f;��a���`'"O� @@Y�6@:q���Y:�D$��"O�b�-\5��Ř���r�x���"Op��t�� [��(�È�l����"O$��L�/ ���H�$X�\�| �s"O\��@J�gbjp�[�)Dz��"On�Ó�$ns��P��Si&�e�a"O�%Ů	"�dxa!�	#�b-9�'�j �C_�@.	b`i t(tT��'���"q@i�����A�z�!�'��kwE'!�(h��#dn|��'��|qe� 6'�
�D�D���'��ĩ`%�U�ޝ���.h,)�'��%H�D��ptjG���*���'"fԛe�AX+�4s�� �
�L��'�BA��Ĵ[ h��I�-H\(�'���w�W�����c蜳k,���
�',>��GLB,,L��s��S	�'�n���01�L:'m�t�T���'�2�#��1HHq3[TFl�'�m� 8�{SN�W��<��'�`�!3��x��KC���R�8��'����vQ�X���9c,եU&P��'}>I����q��(�mȍL�<���'��p���.f���'�2��tI�'��5 �gˁ:�ep�a�"�P��
��� ��T��!$U��(_#��QI�"OX,�U���9E�9@&�i�9S�"O�r����Eke��h���"O���4�Y# 3�D�>6�iP"O�t\wDZ�M�n0��+"O�e@�j��:�Y٦-�ɜ��2"O8�;�Oϣ^�5ʠ�V��j��b"O*�R��!~��@��9�|u[�"O�!"��h��7#��%�e��"OD�X���{�r�ÀB̔u�!�W"O ���/*.!i�&ǳ?n��`�"O�����P�R����>XO���"O0!C�/�ڴ���2L�d �"Od�-gN.��#Y.8.q�b"O�p0�U�p��8V�5?�\
`"O�a��GQΠ��#@�/�jH#F"O4�aU�H�M�����H�>��T"O"��v(M%kʄ�a�
�%n�Z��b"O��Z���N�򄁇
��l�s"OF)K�Á�~���nQ?M&h�5"O�R�Y���u�s�8F��P"O4rU�6j�<CT���M�4yQ"O*���` 1�Xi9#ED�%���"7"O���P�ǚl4��EV�HT*��"O�,97⊴Xn6��dѪ'�̕(V"O��p�P?"Ŋ��7)�;N�(�	�"O���4�ծV�Ԣ�NA$��k�"Ob�G�0j.��'�Ґi�T3"OD ��%K2���^�v��		"O>|�b��9��\CC�Gc�2�QF"O��{v.T)iJ���Ɍ�?���Z�"OBāb�ѓa���g+��<�~�"O2p�G{tz���JE�J۲��"O0%��։9j�����Q��QH@"O"�17.��G�A1���y[��B%"O����+�?�8p� ݭbS��1"O�Ġ�Î�R]�=��^i��q�"O�蛰��P����y,���A"O�E�%ޡ$4�jM�=�챃"OPHsIQ;�U!0	�6"A|9S�"O�@*TIǈ=���5?0>9k�"O:5�aJ�	&;������o9���P"OhHI@F�ā;3eǱ>�HD"O�yCծ��ᆝ	�DD*C����"O:�+��Ƌer�� ��
X�t�F"O���r�D�p �ci���̄�"O��ӑ����Da�g	�C��I��"O�Z��	i��\a��H=)ڮ���"O�e�����j;Za	C�؊�	�"O���tGOZh��䒪,۴=�W"O���ŭ0"������w��q1"Ox��`�r��Фiӗl��hQ"O�=c��O�c!�h�g�	�
���"O�0�G�^<X�HɄ�� bR<w!�$!�݋E{�C�L�N*4�z�'C0�05D��E"e)�$6���'[�<��K!B����Η�e� pr�'A�4z�HY��<���l�qԾ	s�'Pډ��'�3u���cE�S7X��z�'?P�E��\���ξO���
�'2�k���Rkz}� �ӊ�$��	�'�<�{��0\6�2AK�zFr���'{8��(A �D�@����T�'e�0��������ÈM،0X��� ��ǩP�.������(N�L��p"O�Y����"5񎄧d�yh�"Of)�S�Uي�+���g~�tj�"O,���[mK`�2�)z�p"O8]i����c���)W-�Sq��I"O��U���F��j̀>2���c=D��:��!p�B��U�|�p��+'D���b�8[P�#��M ��2��d�F{����:j&A��%�ڈkC-�*_2ax"�ɡOӘH 뒋'ԄP����L�B�ɫ'|D���~)J�ӈ��_�VB�IO�~�
�!��B��ٰh� G�B�Ip���ٴ%АUǮ�@T��+d�N���'��WC*xI@□4F�b�i�$:C��6��"�$�[̶(9gb��zWKB����� ;k�Z�x�Q�x��H�Ac�?�y$�S�p��d�S�3�i�Uf�6�y�O��A����R	�<*����y"!�!$@�����=X�:ud��y���g����Q�6�Mx��#�yrA�:oZV�s�")��q�3���y�b̪W�-�K	)~�$٢�H�y"�E5>�>xq#��&��"S��(�0?�(O�D	E�!-�$�Ѵ�"S�ū&"Or傴e�0e�֭�%c�A��bf"O�����U�0058����l���*�O
��$R�=g�9(C$��}7�Y��A8
!�I��M�c�ݜ)7 ��� �,!�+;�0$KE�/�H�lΨL �C䉨*N��rE_�SlB��e�σcZ���$3ړZQ��1�O��g���a�S3h�	�ȓ�,r�aW�?h��@�V�U��,�` �R�e=e:��ӧ_��P��0���SC�wP�ɕ G6#���?)�\i`��Aح$�-�����z��ȓ6��)�2����y��a��>z ���٠�ElU�n��&�\�nzՆȓS���f.[&��pC�V[8X�ȓbP����������
-0�u��pUt�z!�VQ���$ފ�H��ȓ{``*�� 1����a�O��]�ȓtc�h�-[/d������ 9挆ȓp4��$�S��WnƻdH����I����HD���гaà12�ȓV�Vt����s
 d�f�7H�z�ȓ㾱�֩<e]8s�C��$�JP���Q�I>$M�c �b�)
�C)@� B�	4N������K�E��Ŝ�a�#>�e��u�X9�2.ֳ \�p�ۺyW�C�ɫY�x
% �(*j$	�B/Y*,��䆧�(O?E9�~-D�5�^\;d�~�<-��a�  	K.ph1FǕ/�\�'��}�	҂}.���j�B�Xk+�?�yR͛�9Y�,��%�?��1D��y2��#�� "Rj%��9�" ^ �y��̈́!���*�#~sl�3!�Ĳ�yB��77y`!8�푋{j�u#0�U(�y2c"S�K^~S>����	Ѡ�ȓg�:�)�&Y.nv�)C-[9,��ȓRr��KCB��H9���T�0��Mc3܏9�DӕU(E��y��F^o�<y��u9��r��	��(��a�Box�L�'ք9�'�UD�i����k/��K�'��MU��'ꔙ�0�š-Đi��� ���"�׻�e#ѠO�V�dZ "O.!�Q��&t�������7����5"O����@�+�.0۲f�=M`vd{"Oи1�NՌq���+ c�X��"OntX&N�pZ J��.��M��"O������=X�t�� ����9�t"Op$XrF�4!�*H���7���`�"O�AjF_�*R��P���^��"Ot���1K"tB2K�$f�&e;q"O��c��?P��6$ρi8��2�',� �f�D�}�N<C� 	�^��u�
�'�d����3���R7���"]�lC	�'�\q��8R�\q""�'X�(��'�`� �E�m[��p�×�V��$�
�':��bO�a�^L��αIsnX
�'561��ڧ@�]��ܥ<���h��)��<�`�&��1:Zg�X�ɔ��C?���)ڧ*��`����?M�y�Ƭّ˪̇ȓ*~�����{b�AkbT�Cd]�O����I$���`��o�2�Z3l��\3pC�	<=6�ʆG�!H���ِy���,��4 Y�4�!c(~�X�P��*\zB䉒J�.�X��;�(�Q� !A��#=�Br�� �
hy	Ԧ�#E�Ն�g���X1�X:X vu��M qr��ȓG�$qC�!�� "b��-OtPr
�'�`���'ƍ:�2���4	�'%z0��(�<!�c�U
=���Z�'�����	�/t�4M��3~\�1��6�T��`���HE��n�(/<�ig�*D�ԩ�+Z�R�BM��b�������&�$�Q�b>uk��!0@I�`��()�4`�%D���4�n�� x�,	A�%��nӚ�=E��4?���"�$�5bZ|#b���b)��D�'0���G��%*�\C��XJ>�.O|��E�6A��3��'Qj�逊��{8!�Ā 0nz���/C5jn�jCi�7K!���wC�\´#��Rtڧ��*�qO
�=%?�@ ��'�>1S*��T��%�"D���� �'}�m��2^�h����#D��p#�O�?㾜z�,Z���b�K&�O@�'$ƙ3ŢP\<5�u��[&D���'�� I �-t%�	�ub��=���'�T8h��=��m0eCD-�.4[�'�r�Srn�9m<�s�RtT!����;,O��o����Ej��"O�ԋF%؅*���&���H�e��"O҅{�+ǋ/�-3��.��[��'�����c�6>/���4�3Oa�-�ȓ9���5�͊�r�i�e��B8���#���4j
�
Zh�@,E*d^p�ȓ"��2�� Q^��P@�ɦ]�D��S#0�d0K�G2><D�vgV�U.B�	0q���) nʓk��sϔ;B�I�oLS��γ��� " ���"Od�j�%ݒ
��qE�2Mݸ	×��0LOx�k%dG=)~�#p+�;+$2�y�'>Q��1u���a���a��XSX���8D�(���N(�1B��;[X����5�8�S�-���!��>�����0$E���ȓf�6�a�+A?k˔�VhT(ᔁ�ȓ.P��UH��h
���O'T�K8D����$q��G۵c5,mF)2D���.�/nD91�ĩo�h�"$D�� �삦H�6ׄI�z�=y�"O�9���N-Jt�@V@L�n��K�"O�Eb%��2Hܬ��oT�R��	�f"Or������6�0<�r�,���ӑ"Oި8!��%C,��Dn@�(�B�"O$���޵J2Jɀ��_�{���b"O� �@cɛQ�\�$l�鉴"Ol�2�� or�łpLR5~Sd��"O��#�f��e��ӥ@�`�"OBy) ����Ԭ1T.\�`"O�)�n�u`��J�N$aL<��"O�m���J��y��I56@\���"OҁSA��"pɓ_�j�4$�S"O�	(�G��s�~05�+
V�D�B"O�s�%S�a�l�XS�F�e[�`�R"Oȹ�t�0�9�a!D4"�)c�"O�J�M.�����D�؈=�"O,�Y0GL2u<΅��O�rﾱ�`"Oj](�k޸w�r�eC�Y�V�2�"Ol������G� ٳ���G�� �"O���GJF*�y��m��*���"O� a�(E%o1�-�3�U,�Z0�"O�� RkX2'�0Ah���-����"O�]3�)A�,���D�`M��"O �$�D5=��A��άr���@p"O\�r� `�.i�ݔ1C��"O�T10G��W;�4p!�}�EE"O�yc4�F��T�

tS�"Ob-��9<NY
3gơw�x�yP"O�"�ŊB#(��,��?E�M�7"O��bQB	*F3� ����%� �p"OtH�!@Ԍ8���C���4�"O��rv��#,� ��"�ɠD�ʥq�"ObHS�Ö�~Q^�0a��7����"O�As1�U����3�J��C"O�P��=3����f��{��P�0�'}6}`�f��?vE�c�I�vZ�ȫ���<nA��'�.`#��.:�Іh�87��Y�'�up�L�d%Ρ:���8G��X�'r��vDW3�j�Z2���!��7�p��*�f<[�:�!�;|٦|K��!X�=Ad
 g�!��f�	�@�:c�1��/ը)�!�ܝ?���!����vl�&.�	/�!�O\2����˪A�ph
�̐�|֡�dB#~~��$�U5GW�����%�y"%�'0y�P�.�C�Tqxa�,�y�B��M<"�����G��ICgǄ��y��){*8(j�IW%i�����k���yB`ȆpX:�����&l�E���y�S$!"�P�D�)&hm�%��y��1g� ��*U0=
������yR�ĭK��I�'��(ު�i�Ν.�yB��?$#�Y{D&\2�8�I�B���y�HO�	�*������	�6h�� �"�y�W *�L�)1�]�h���\�y�EG�	�H2eK#Q40z�N���y�eJ�(%0�p�M'��	+s�S�y�����8���}H�16�E/�yRˁ�<����-�j2v��4���yR×3�T�u��j��L��W��y���DJR��+�.���AH��yr�E0�;W	B^�MP$+��yAZ	j�!h%`����l(� �y
� ��7��X8�(�qb6C➝i"Obu���o�x9#���|��U�0"OJ�K�cC'g�S�V
b��#s"O�t9A�ɒR�����ЮV���0�"O�]{w	D�M�Z�Ė�(�L}�p"O"�dgɍi��	��P7!L��"O�݉��&3�e�P��)O�Re�R"O�ڷ�+g+x�����gٲ�xr"O ���O'1w|]ʡi
];Ha�`"O�<:��A8Pt�}���#&N����"O�� �H�}
��C�o͐RpU��"O,�P��%��C�.�+]X��"O"]�#n��]n~HՀ�5&Lpa��"O����@i���a�۝~���r�"OP�+OA iZ��u Ҡ�F�s�"Od�b�bM�`���*��N�P�ܬ�6"Ob�	S��x�@iQĂ�lf�IE"O�p��+�N-.���!��A� q�A"O>Ģ���'H0N��po�4x��� �"O.�����pOv���n��,���q�"O��ૐ>V�h��DL�"9GxQ�"Or�Q�gO_���l�=|1�hSR"O	h��W���V�GW6d"O��y����5R2�0 i�V�p�"O��ף[�o�Lu괩�=Y2�%��"O�cAMȘA"�1h�!%�$ �"O��ʃ"��]�F<�热D�Q���"ͬ|�B����F��蘍_u�)��U�`$�*�D��y�eC�L�3S��4M�mR��Z>��LT91�@Ü''��q�𙟜�Đ�����+gS��1�#4����h����.����0ȁ�m����V��9r���o��<�&ђ,�Ҹ*�
�P�q��e�AX��i�Տ$����k' u�<z2ä��m�� �=����j�!�4B�	�c�dXzÍS�0����M�N8�'��q(W�l�TH��֎O�n�R�<�`�ѹ��FE/Di����@��B�I�������P)2��\ (���@ɞ9:��(���#B���!�*��!��ɶi�� ��*A�SL� ��z���
O�B2� f��E�rF�/h�2�Y�O��� &�+j~���MBf���	+sF�Ht��T6)�#mQf���dф|tB�T�N7Bz�)k*�R^��*"��Ediyo�;g̅2��m(<�fS!16�%�R�͇
�@��C@A��H�F�P�F��PR���8GS���p�3a�S��D��㌐�k�^貐�͢g��C�I�L�����G�P����"��CD��$�!��E�� Z������'}��0z��p���n*d.`-
W�ިG�l��)1�\I���(1v�պ�G�#=��z�� y��z�GݮqRe@"��(c͒0�'ڪ4z��ڈ�DJ�T��ҧ]�?���E�N�l�x2�uJ���+�/>$ ��"T�^n��T�K6�NT�r荱N]Lѕ&�J°�QS��E�H���?Al:��ƀ��~�^�S�+}��>.�*�`���,�"̐��>�
ԛB��	qf�y���e�Qx1�0-7��!K�S����ȓ^] �;��Q]�r-[l�\*��ѥ�>P�f�Lɘ['����� <��S4�X8��w���:5� ���ȸ�� 
H0X�'�tI���6lK���K5V^b|�p��eu�m�f��H��x;%����rY1�G�oB����Q):�[�)X+zЙ�1?LO�!�T,�<�Z��p��m�`�CeڞQ��H1�l�y�rܐ��5=[��q�K`�����S$���KgOS�Q����)��8n�`�8{ORhv�T�s$�x��Ur�*R3�6A�vG�?��6Ms��)X�c���;�H�6j�!�DM�?~\�qү I������9<���s�� �d=���K+[tn�k1c��<zZ��OQD�ڃ�y���P�HE/�';�:6���p?a4��	CX|���P�X���Zu�%u�b��w`��8f���H�Rٔm*�ϗ	z8e��>[���2��$��w	��7��<�Qs)L�}/��®8 �ȁ�ӠV&0`8��B��(����ŨI9�!É�J�a����]RN��D�7�&̸d�0LO�u"���D,�H ��,�zY��'K
li��ڀ �|ɉb�VP�AZd$�C#�-,��T뉨�0R2� 4�^���+X#g������_8N��.ZU佋��ۈa�pّ�!Pt|����8n���Xf
�MX	"W�^Rꡫ��	b�P�!dT�U�� ��wf�:F�X�!bݭC=d��'��h��ڌ,J�1ѯE:RN�@g����D��^�#Aew!�Չ��=@�`X�_T�8�bۜ�
�'�v5p�l�Z�,aJã�[��y��_�f(S�\�2]23CX�\��M�����0R�3�`H�~� �G6Sw��҅H�4��ס� $*jD%�o8�i3� R}���CC汒��ɑ7wVjeGJ+<YZ|H�ߨ~�� �ģUr��ҳ�e���G/�3zTh��نy�����M��T��)N�Y\��dE�+�p=@&D::�֜Jw��9 L��b�oR���i��*@	qX��2�r}��Ae(tZ�](T5a%�ƉdWlA�� ��q�����w1�u��*ÅR�8�k䮎y���%G��s���r̓�D������^{r�@�*�	'�&�3T�O�|��5�էWH�D&W����r���f0�ȡ�l�Q�d��[�R�����cA<`;�1+��iۮU��ܔG�HQ&���K$���7)D�?�qDiՖf���Bعy�Nt�	ǓD)�r�!Jj6U5�	9qRx�H�B@�4��Xq��W���[We�G!�*S��e�dȺv]f� $��n� 1#�^� ���c�;�H��fM2�QS%��P��P��`׋1ډAā�6S^ ;U�J6)	z��'B )����U��P�B@	7ĵ9Ҥ`ޅ0��ݲ5k�LCr
�9�=P�!�O:�[���$���$R|��R��4A^`��զM*��ó[��ܒp�I�k�@$���'� ���ͯ
b���O���Ϊ	��<RS��r˔��4�I�l�`�c�C�;��80�k�3'`,��v0^OHa3�F0*[�(�D�2���dյ4t~8�Be�VEJ
�/Oԅ�F��)3��hP֡�<c(���'�`�
ëɅb��[6�A�<:ܝ���Ǫ4��T̓d'$�Sc�9�eL~��j�	��F#��B�/S�e���ā
n\Ҕ����8�P�Z7*�Z ��`ƤLۼ�ڡC�^�A��D�	|p�D-�*�.��<W����&�r�
�b��D����׫+�`�K�&9\�R���W0��t�S�C*�̈AM�*gz�Y�H� 5a	ۺ�
V� R6����S�	�-`��T�ِY5���C�Bb�0��P.=�x����bJt�(4�J�I��2C��\��G
5�:88��Kj1 �n�V_`�(I� 6�P(�4�'$ls@	־MC"�������B1�n��D�>r��`X��,a&jC0	W<HH4�sG	����Z�"�1�'�K�9�h��D�H��#�OΔɑ��,F< �G�\��Ksj̙� �J��N{�a�q�>0�Ь�-S,F?<�$G\Z��{#���F�p�Y&J���#k~�-��'�F��(��`A��S#A7`d*�a7�M�"4zpۃɔ?�$�S�ƃp��b2#Ƕ>�B��+S�b`"�y>�~|�K>y2�����$	:��tÀ@�v̓:��`��@ٴ"�~�p��MM������1���%�\!��LzN�C�J�0��m�NT1V �ܹt���w��܆�IL�P� IR)X��)1�˩-��M��O	�<��U����²�z>�0�(\��p�jJ�+��q�t�E�/���f�*X<@����1|z<�Ɠ2���	�O�i2�]� *�`Q�$+���#��8�棝'�uh��ʱ4���y*��n?�i�jcT�(#��%$�y��^%-PԄ1��QQ�l��ɖ)nȄ�pȁ�O*�p��M����C�TH��_�d��@N^�96�q�$�Pl�E{6����򉦟�'�M�D\�7�NPb#ڠB�\r�y2d�!@�t*4a_�M��}8#H�7C�O��u ���y���
�E� i�����[!�	٧H-4P����9<O����&;M(��$�]Ht%�p.Y�8�X��þhH���D�����y܌:��	��%��G�2\E90�O/K�phF�G=B2�B�	5g2ґ3E@G�j�bH��Y��>Qc���PfL��J6��ʐg��)��Μ(��D�e�P �T�O��r�I;N�H�H���R:|���S&Z�K��Z)���&`J=�����`��GM�1"~�s ͑:v�@�O ����@[�g}b-��vA��DǾP�Ӈ�'��'^���#�oqT�{�˂�*_� �S]�& 1�χ�y*T�xp>u��DB�x@��bM���	tάS�="���?~�p�"����B����mP"a�r��w�'y�"}�'�Ҩ�УH�h�PL�#�-`+��
�'W� ��G���݈��]$]W2-ڴD P�ĢT:Tک����&�p<9�eHV� `w����0t�7�H����k�z�����p|��%eÊa�R�r$[w�M GO��FkZ�i�8�e�	Ev(��ɢ9b���vڻh�>���K0����d/ՠ"�"�0�A*D�("רD�)vXj��n����OH��A�%�����JH�d�#n'��[B҆L�� F4D�� R�0=�f�u!��
��`qC�4D�X��	J�
�֡Z"�F�{���P�'5D�x�C.#�E�����kj� �)D�|��W�X_�!�Cʈ0N�tSd'&D�|ɀǚ==���b�I -㚈�r"D�X
���U�>lS#* \�<�sr�"D���@熺�n7�<��4�d�R}�<�0@�3$�jA*�9-�ɑ5��{�<i���0)Q"�\:Q2��T%�Y�<� �-B�b�>/��P�@,Ek���"O���@B�e$r�B�@�.UF��U"OL��'���A�6�I�E�~�`}x"O�H@5�� Z�� $M_�;_xz�"O�������8��,�%A4�D"O�5��K���i��l����U"O<\�:��� �K�Xqh�6L2D���D����15�ɛ*�%��/D�jf�8,�x�C���an��;��,D��� �Ж~��Y6� �+�D%s�b!D��a��QL�1Ճ�7"�XŢ:D�x	֯gܖ��à/M�Rv`6D�l�c[�[^0�7$ؾZ3$hi��#D�T:�C�6���$e�	b"��2&�#D��c3	L $*л孔%���e�#D���rUQ�x�{�k���8�>D�H��H�-̑jv*'+>eHg�)D���hR$�6 ���4YlN�X��!D�䓲�ə �F�{E�J`�l��l?D�L���x������F�n���O/D�X��h�fP �b"��,�, s�K*D��ca��K���X�u�8H#I(D�����' ��s�Y�?�8y�&-D��3��������^F�ط�,D��!7GQnk�����W��)c'D��;��G S.X�r�o >l&9��$D�������ؠ*
�j�!��7D��bVL�TR��򵅝�_��*'�5D��Vm�<�у޼]}���u<D��蓫Ϣ$��g8oy2����'D�x���=)�(�Iቚ5D���#$D���	�gF�u���[GH�yd�0D�t �!�e.(K ��#_�q���2D�pc񤔌!D)��KԽGJd:�7D�D��MA\H���KR
=�(XQ�m/D��5Ł2.�8"ϒ$c:��&*&D�ı���L.�c��v�L��w� D�xk&MR<IC�0J/O'}�D�8�I+D�#�F[�{Wb�� S,g�HAye�)D����k�0`��	�ZuPB'3D�d�Q��7Z<p��L�	L��I��,D�hK���\��H"�ف8	�� �m(D��#p��X��Qə;��h 7�)D����� P4BA1��/{�<�U�'D��"��
Qo�lH��кl�|�S!&D�lx�hL*bx���(�7�0D��
�MB7ʶ��4^�䩑�.D�,7ܒO�b�"��L�:��X�$-D�ġ��C
C�hS2`F/l��Q'.D�,���Z����9���0p���� D�\�a� ��$HЃ%G�q3-D� �#d;/b�X9��~��Ea0�>D�g&�#���d. \��Yk�!<D��R���48�t�b�xl�J�E=D�����R}t��F�xY��/D�̩�l�(�2Azr)��3��,D��6�L�m�D�X4$��6:��K�(-D�<B�?L*�3�h��k��'V!�$:5��q򒤃�'=4Q �`Y�	�!�DLF�`	2u,J)t��S��!�N�`0uГ�%�D�kK�{!�&(B����D>H�1�
�KT!�dH��
�s�[�~�J�w�T�M!�U&`H8\����#O�1�����!�� ���'���Ñ��_ِ刣"O��ۣ��"P�Y`���?h��s�"O^E[�����A�τ$.a�MI�"O
��!��b��XQRnWT�x�"O�xc5*Y r֪�(��\"�b�"O��)EjH�����QK�> �$�Z�"O���1n�$z jM5�����"O°���-G����j&���W"OX A��I�-��Y�B��%R��"O���V@�l��h���LD��"O��isE�g��iXe/ɣuUf8	A"O�lQ�Ϛ�K�ͰS��HWA��"Oxh��ڽHk�q�O��FW�� �"O �JU& ���#Sh��](�8�"O���ˇ�
 H���ĦO��Q�"O24B%���B)��)C���!%�L��"O�(1�A�4�Y�@�B��$"O�P��%�.a���h�.���"O���0�C,P"t�]Ԃ��"OVXh�D��
}��Ƣ0�(���"O�V�B�{�l���F�1_t�a�"Ox��R�Z�q�+sD٫&j��b�"O�t0 M]_R�mۆ#ƻW'
�ط"O� �cM��j�H욡�A�X..5H%"OT�w��K�B,
�O�p��%ɐ"Orq��K
"�y��1y��� "OTT�+Z�%���s�Y%�~5��"O����Q���`��)irA7"O8�1�FJ����6���uBL��"O�����}�
p3���H3	��"O�U���g�rd	m�e%��h��dȲ}X<���X�+φ8G�TLɟ`$n4�˝���L÷�Y��y"���(QMY& q�.�'�@ạ$^ܒi"�'��P��� iB�UpvI��V�P����C�%4�D�ER�)�N��Ԇ�('�.M�GI£^P*M�R(ĘIk��B"o$��<	�oB0'r�M���
&ZE�=<O�A3ư�K�!B���f�_�bP���u�ω:�YഊE�*Yr�26%+$��h�΍�xq�畬X�fH�=}bI�*Z���ذ.H8d����.���>���e�;<U�$����u=�e0q�?D��BD��!>�03J��v�Ub�䚯A_^�B��6���y�a�$R@��>��H��P�E�:N".��t)�cU��Qr/$���BdϩCr���6��9��a`��C�\$��b�=j����؄r2����e;\їk��Sb�"n�l8���&�,xsPu�� K;"�v�B�M�_֘��-N[]��VJ����l��'�l5���)|����ăA�(�L��#�#Ʌ4��(�I].!�FXr�O�8A>�p 3h�|*�h�
m�-hGiV �ޝ���a�<Y��ҎL�Ƶ�Ĩ��t�[�A6R�0٠�8H�h��L>DQ\C�����?FUP�;([줘 �˶[7��AR�B>�I�,r^ڰ��4+^�@��;��@�k� 
�i����g��`	'�*�  ��-RQ��{�MQ�o�(:$fA)����G!O��0� �L��ꉜ��Xk�F	n$�T�D$Lڼ�&d�'D~n��6��_G,mP
��
�e�] Zb=�ub�(:ڼ�O8�Z�ĔU}�]C����$���CЋ.#�\HQ5��6!2�@��f��HS����D[�CY�y��#q���f�����E�Y=Z]p%Z7)љn�~��@��"[���%עp��@� ,�7;�>|)rg�gK�M�gN�G����@O�X�G`V�x�Ą�P�@<���||)���9�aR�@�bT��ր{�֨�?���L P���!�$ȡ�̖K��pb�c��i��(�+s��o�q����NN�B�@S� E-l��ܳ��ۈY�켇�	�"��CD�5@����(� B��'�F��C�F����_��r)����7
I�p��8�
��K��"u ܿP���{W)r�<�&��]E64�t�N�p�`'N�Mf�M����0OX��b�ᚂs�F\�t�'\G�Ӹ�
�3�{��
��U�X��� c@�6
�.����9�O21hv��T���"K�/x�> 1���!~��tʕ���4�*���.��Dwt$��
�$[���s���|�$�=�À�2H1H�7h9�d��d�n�'|�B�I"���v-F	���g��р ����'PѶ]�m�.)SB!!��Ώ_r)��Z��\��'�6y�bÔ rxr�.TzB%���.5Dr����s�P����z�,E��#U� lD
'��|T��͓&.���3N!Lb�EEp޼k�OP�����:AL�!T�]�ҵZo�-S�{��F�`���]�w�J���%;CK�$��X�ę�?���a��+v���0�Ϣ�`�.�p>��)��~��s�E�P�иk��)_O����G7'�:�uI��]X��u$O*gs`H"H?V�ʌ@��X@��j&�>	�D[J�f���&������F�']ju0!��O�p�y`��!���3eWE�9y�
�:q�"��3��F����l<`�n�kw�Ì;�N�0DA�	/����D�br����C(B�
4����t�F瞲KC&�J$L�0y!b�0W��d�1�$��E��dVr�1iV�?Mcj�ydD��k��X�׮F�=;���'¶u0�dI��Q��kǆ8ۘ%����EE(�Ȥ��M�0'��e2�Q���������
~�#�3��اG��}�$y��d�E��'�~�1�mRf9�ՉCaǄ���ɄH�:�	���9r\�ޞO���c\9N�����ё4(@5��'j�ŐBF<9O�h
�Lϻ���ۈ�dO�m��𒥇�>@�\RRl�9���p&�/��\����a����qQ$��Y8P��n/d��!8�n(�)êv�xb얹G�v��

<0���Uc�8�l�S�j�~����cۘZ<蕋�;B�n����k�����_��x�CD��P �1ӥb�gT:0�D�Q���2D�QשE���R���	L|�j3�Av�L ���-󄑩5K�1w鄑��
AA_�Ks��;;�T s��a4��f)��}!U��ɜ�N�ԧ�Z�e"�k;��0%)	�
�.۴M�z�;W�ӓ�8Q��&m����J;u,)�*���I?� L;�G�2�-��6N��=��O�ؔ�)R�ƅ�Hy��MD-v�${�'/|����e$X�5۳dͳ%p�̺w��^�u:圲>O�8�㉁	�v�rH*{��b$�֊�$�,t�����hA�Aߪ4�-��
�d���ک�y�-ʂۜ=�p��A%�!��A8Ku�E"�%��h ���'�0ѯ� b:	CW@Z�xir��a@
�
��2v�͚�fǎc�hAOA!d6��/~dh�@�wJ��y��ڽ�'0�� 
�3��@Ċb�\�c$lζ>��5`�R�<���H��D��L�3L�:y���=�J�3���7?��)Z��|r�O�z&(����!k�@��F%���hO8�ҳ��������?S��]iDMë;�^��U7@�y��4 �L
�ZHJ�؁� �U���Cx�st�/�I����;tC�m�`��iQ��V�a�66� k4�L+�e�P(T� H;��̲D�Șh�@ŚHZFT�+^���Ih<ygGݬah�pҷ��(o�F��˅�uu�7M�L�\]{%��~p��.�9\�޸��/�7S�Z������y�G;L��9Z�L��]̊�3D���?�%n��t�� ��JK�}�I*�KJ'��0���ΐL��@��KP�@��\H�IN�?��0��*��|:��*�Ĕw��	{s��S���ѣ�֧M�џpj�M=i8J��Or��n�@X�Qz��+�MyF��0s4H4�X&aO�����d����I�8�!+�Aє5&�hClӏ\N^��D����)���e�`�B���]��2�G+)��(өF�N���>4��1f	����7p/�@�"�#}2i�l�N����5� I�b6��O�v	���A��`�bg�-3��A��'���;'��?;���'���'������>v����S��x�db�iʊ����ǜ ���;�� H�� ��>��e14�3�	z�����̗�x���%��28���G�{�p)���'r��R6OL^04�Q�.U�si�ԓ���k�J8��S:�v!;�#-v�X��I�%����U�_�<1�j��#樱�G��+����mQnܓ�r�����W�)g�S� n���/F�iz�袥cEf�&C�I8�(� ��f� �10��QA6��`��
��q�O�`F��O|�H�`��<^ع���L��<��"O�U�rH3m~p=�Q�@U�$XJ��'�68��GW3�����
KV�@���;-�L�LC�m;!�� �"��dB	31b$I��J$2)!�DϫL8 9b��B7`%�}�`�3!��׆5�x}��_�c{̨�wmٕ.-!�B�$ �U�F�[$k`��c�߆�!�D�)X-��pGX�iu>��3i��3p!�$6<
޸"s�O�ex�蜔'!�C~�9�OñbiY���8�!��'�"}(�4wђ�EN�d�!��_0�� Q�f��Ń�C�!�Ê���(��ӵ5���7+��!���l�<@3 �qsZ<�Ck�k!���n[��yg"�o�\3�^1�!��>H!6�0bE��hD�+S!U�#!�� �m�6�S�R�N�Y����I�"O.T�k}�|�ytX$#\��q"Oj`ᔣ�?Q��x�c�$2B̫Q"OA���B�%��Ř�@)f<f��"O&ܫ��){�B&��u�yZe"O	����5D&6iIBm_�)^@)x"O0t��&�	
�D�ԬگnP��QS"O�aA�$I�j��\���¨r[� s"O�t�僜1U�0Y��Z�t��T��"O!1��\�m�@i�'T�BrD<�S"Of��1��[� �`%C��l� �"OtIY�Ɍ�1����f�`��t��"O��X'�U�"v�����5�n��@"O�!�v��~E�V��L����"O��bբ
>J��[wB�6��!9�"OP@�R��<�H�R���a��P"Oz����7��G����w"OR�C"W�(!4��r��a�*O��ʮ]�xjmX�aHM�	�'��v�N>WS�"��Zu�@y
�'#�p�"�B8{.�9h"��Hd ��'����G.3�,l����?>��j	�'ڲ�;�bΞL��ؘ�IL e��
�'���!R��yf`Mر�� q����'`�)��+j ����B9k���C�'�D`&��m �웱��%~���'�����K�k�|��QX
�C�'Z|ܐ��&y^:���F�r�p���'L��ծ-5̙R(T7F|0��'H
!{���wm�i�.��;2�;�'�$0Ģ�
L�q�Q�70�$�+
�':���¯�+=���*F
�1���
�'��AW��ѣ�`B�c���
�'�\�b���;2�]�iT�]`�(0�'�
%æh�A�1H�&�@�
�2�'�:]�H˵^��pp��j�2|��'#�$�Vm^���֎dۜ���'�("&
 3��<IP�\�f��,[�'�l ��.�B,|9
�E��Cy�	�
�'���B-L5�#W倍SԜ	�'m�h��l��O�����"��e�x[	�'������a�R-eJXP�i	�'�^x��k�3(50Ę��"_z��p	�'4�A� /T�b�� 2��z#j0������K�
�!���5�6<@',@�$rx�0���B���A:a ����I*r���?�;$rz���]��H��ҴE���S�Iq=�h�e`�$.ISTˎ�U@��)��@�a��e;()��o4$���O�.�]S����~2)^���'¸O$@yd�5($�v�B�2�	@#`BG��!�4��7 m�7�<;��
�MзpKX�jR�ۙPB��o����ń73�����X�fP�=(���T��t�JqB��Op�I��'z�ڠ'�b>u�'����p����苗�ӿ���8�n���(� nξxh8�S�|̧T2��wd�������B	-���B5�̀~Fd<)O��s���V��/�h�]�!�]�ptR|{q%�$A��e��<A�ͅ�@��|���e �d�:NC�� �G2z@0�>�8e<��<�r���!l4<�������� CŚ�<��f��	�l�I>�'��O���C�E�cu���D^
�x��HJ�D]99F���� �$�!BV={z|�F�DJZ� ��!�	�%,a��V�0=tpc�C�yLd9��<����>9���s������i�u�		G^Lz Y�RJ�� ��t�`ą$7 ��W�h?��DS����&���D�6A�����e߷9�� mt�>A���?	�5��c��8qY�L�KP��b]��A^��?�%�D}��i5YM�Y%��K�h�.h"ES�AG�YL��B>K�j��	�5��E��NBbIs��W��8��ٸ
��)�'��	 f�(��O�h��(NOi��E��8n�V��ߴm3�Ʋi
D�*�D\w?[w������ L���������5�1Ƥ�a섰;X�l�@�O�]��dL���OǦʧD���!��cZ=�U+�,>�LB aT�~0L���\�`��#�d�d�O��O�H����՘��E�q��кi���ĬNN\�a�'g���m]>}胄�}An=!��E5H��a©�>Izc�tb��Y�ԓG��\�@P�1 �4�b�z��)D�$i%-a�K4�V�?n0��=G!�Q��,�pc4�q���Q>!�dr�d����O�E6�$ҐMƺ:fPB�Ʉm*����T61��r��+uB�ɥ*�PA�Sx��t
b���2BB�I
�~u���[�	��X\:B�	�q'D<س��J���q��&�B�I��TN��b5H���B�I#,��i�2o�h����̠8<�C�	�6��0#���E�
EC�.r�X�Q/Z/���!�sb�B�I1�<̚�ȑ=y���yv)� !̈B�M�����j�-d�R���	�s�C�I+�!��Y!K�V��dkL�.C�	�J��pj���@�D� $�9
�B�ɲ��y��嚫0�8C ��~/:B�	8����0B��Y[�AO�c�TB��0E�����,_t�dE�.>R2B�I�	��[2e[�U��;1(H�{ �C�I�{vtH���V>/�l��sm��2��C�#(m���%� FX�Rb̦�B�	\
\��$MS2h�\����&d�C䉬3p8�Q��,�B�	��,C�	(.�"��w����� ckT
PC�	�(ǌ��r�ԘQcx�˲ �9�C� 'x!�7 �(t�\�3�Y/m$ C�I!+�,d±��Ê�h��!D�#�Ρl�\�w�F{�y��?D�<�k߭��܀W��A��Kj8D��0�E�v������%~�Ac��3D�Ѓ�'��Ty�؁���-�T���%D��[�/,x���h�F)qޢl���&D��gF!H����/ƃ3pnH��l D�,À�:"f1��	'Y�3��=D��3���1������HI�$;A�8D��z�jQ�<�$ k$lH$ި�wK+D����'ȩ8�0�ɦ&zl��6D���� � /�������:���ٲO7D��J�)�-wPh��b섡?���R�,+D��Z%
	�v@ի�C=͚�)F�*D���͓�r�A�G"WDx8;�h(D��zpN��Z_l, uaJ'�:�*C�:D�h���̗&�T���E<l:�Q�U�9D�@Y��q��*�ߖ%��M��K6D���$���k��^�U������/D���g�ҞJ�$����v���ʂ�.D�d����o�t���(0��� +D��a��ɲ������s����E(D��@�K�g.����DY�9c�cV�$D������@І%B%j�0ٲ�S�*O��ے�U<xfn�� \���I��"O�u*�F��h��	��۱a�"yɑ"O%�oÆ`a��`��%i�6 �'"ON	C�$
�+n�hHì�Pye"O���[>v�|B���r0TpA"OD1�5nU>|<��`�I�N�X�Q"OН�&,̇�fM���[3��КB"OČ�rl�)ƺ�`���.89Y"Oh5K���-t?E �ǫn�&\�C"O� F����JuU����	J����j"O 
�fK�{�>���O�'�
u�"O(��`�����B��Uڞ��"O0A#1ǜ1��t)E�M!���P"O���C�(0�h���Q���"O�a8����4ih0��`'Rpr�$"O���n���yU�xx|�;�"O�� GfR�\a��6&Q�u^�)�"O�}ض���>�ށzf�]���4Ӵ"O�M�%$�3u� m�6D(FI��W"O�-
5BK�5hZ�HC�<؞D�%"O�Lz���.Mf��$O��& ��0"O�L��P4���0�ɱ6=�٫�"O��iB.Oh�����Zx #B"O���Vݒx��S�E 7S:�a��"O&@���^"�ȕ��#T]͚ ��"OZ)Ң���)��qv�A�`�z���"O5+��
0t�D	��]�
��1"O�!*2�]*mz�I���Qg5"=S�"O��d��8��8H�NI�C3έ��"O�ۄF]�/���qAO�s�PLZd"O8<ӤkJ@Ũ��F���"O�5�I�Y�������<o��s'"O��#L��Fа1{�K@�cZ����"O*�3�ݬl��� �&GR���t"O�S�eC������?���@"O��(���&[<<��S얡jT8���"OhM�E��̂,�("�����"O�y�@�8u,��+1Ɍ��P"O�\�����b,`W�@`��"OD �$Î_F�9P���}�hzT"OA�Sh�"V�R(kei�<�T8�S"OT����U�,� �H��@nM�"O
��v��~�H�[�E�%3K�H�"Oڴ��mE12V8���m��<?��#"O~�(#�֚r�r1K��۩^��=@u*Ol��3+ƕ����5u�,�i	�'e����L<5��t��H��'<L�`b�]�?�V�ا�l>H���'[��
#���EY2xpdh��'��t�v.�V*�(7$��u�(�{�'`������4[q�Y	ov�]r�'/Ҡ�f!�Og��cgQ	4�޸r�'>l1!V"�=��4QfK�;�&t��'aTqP ��FV���4
V�,��D��'��E�ӫO�,�ڜ�cߍ.b����'������� F�ܤRe\1��)�'��1�ǎ�h`upE��~ˤI�'4��Q!'�2[Y h�d̓-vY6���'�h�sA���0����,F5Z����'� x����Ar$5�P �@��0�'Ѐ���S:_K�0�G��0�2�'76ly3D,�˦)�.�,4s�'2�}�l��JK���`�T,"���	�'�r�W�1�&�Q@㇭���P	�'\|X��E�(���Rpݺ~y�	�' ���S#���h@�ÕJ��tr�'fdA��Ùay���A%B^Z���'��àb�	sbN\s�.�o����	�'(�<��ܐFN�� �!J*3�d�R	�']H `v�αdI�0�.�.���'�B�i��R�Cf�r��J$]y�<K�'O��e��F���H��*}HPP��'�@Y���Z�Tyw��.mEX���� z}
�N��y���i��H0c�i�6"Om�C�� >����	%e_��*�"O����X#z�}to�1z�܁�4"O����jG�
�n�ӄ-�D�d!(A"OB4�Q�{��"2�#�
 	�"O�eJӯ�
,2���[r�����y�Ο+���3��P{{xp�V�=�y�,íj��Z�cѕw�VM��
��y��T�:	�l3��y�܅�ƩQ��y��Tژ�sq�F5?�8t�F��?�y�Ɍ>����!H�T�u��؄ȓ0iJ�R��K�u�ԡ�%[*���ȓZ�~͈�W��xY��G%�lE�ȓ�ʝ	#�{������M�\$�(�ȓ\8�]��λN/�UO�5=ta�����5�E��tʧ)�����ȓz�`�W��*�(�g�q<HՄ�	���C���WB,1q��� ��}�ȓpy�ơ��a��	����'�� ��5D�� ��W"fH����߹)����9���J�L=��pGIvч��L��ⓥ?�Xx�r��29�.ćȓJ��q��2�֨��C0G�n��z�NE���$�m5Õ�s�����.U#!k]_^궎�)����o�����O׶5�F����Ѻ.�V��ȓ� �0�`��]����f��z�����E����nV�AΈ�V��ȓ5��Z����	 `��C��	[���lc���R�� �]Y@M�j�jY��~;\2��2N&����ւzU����>�2䛤k�zU��$�BW���ȓ&_��9tl��f���fOp2Ќ��T��h�*���k&B5OR���T��xv]�S���(E4|��l��\r�kA�dیPR�g�!^�ȓrB<\@wF�??�|}*�iB������vt� ��,�&��7���r���Ǆ:\rv��Rm�>F}LP�A;D�4SF�JW��F[�Tt��>D��X�]�E�=��K�j��m(D��S�鞷t��`����d?��x��'D�,{!��88 j��Ņ�l�
��R�2D�dH1��'"���%� �\��)0D�ˑ#˘v��p���$s �P��-D��s��دs
xyb�#_��͋"-D�t#c��pX^Yu���\
0��+,D�(ё�<��T�-�	`�%��+D�xж�3/E�����ĘW`���/D��j�e�S�6�zs���uB� %c-T�|*�	O+3��}�7��&U��=��"O�QR	���a�O� ���90"Oʼ"��#O'ڭ��A�����"O��
3/��hy��3S!�-T҄%8�"O�ź���h�����O�Vl�E"O�3�E�/K�h� ֘x� I�`"Or]"�:j��Y��
��d�,��"O���7�g��ys K6?�Bɓp"O�a@Ai֜5#^U1&���A|�Ed"O��#D��lȤ�X`.Cst�r"O��� L�>e�~��5�!l�di�"OH�A"+�#\��z�a�<���H3"O֥��DJ_[�|J�N̷jh�F"O*���'�g��Āf��1]l9�#"O� �](!�ѮN��%j�Μ�\����"O��C�_����5hfm�a"O�eHP��Y��=y�@�eS���"O�!JgOҬM�n h7LO6�tG"O:2N�.&�,kE��0H?�I��"O$���e_80��Չ�ƯG*�!G"O�!
'��T�|��@���y�"O̅94�6\o�ܳ!C�
�3�"OƱqq@� e�}�4�ѡ]�褲�"O���   ���8D�����'_[&�{���b,*�� $7D�� �L)7L�#-Ǩ�@��R=de�Sc"O~q�&�
�0���Mb��)�"OfH�6�\�>�`r��J�J}��"O⸐���(PQ�\ �'��U9�"O���	eD `8��=Wq�(Z�"OJ�� N�40� ���[�y1ԥ��"O��H�D�:d�T�[�l�c0�|H�"O�\3���75���KЫJ	�9%"O.Dc
�,r\岵³[�X�"O@�ڒ �K�S�'�0Ȕ"O������s������

d����"O�)#��5�P����;���D"OVPD�%a0����2=z��"O�A	Ҥ�<R���cF:6w�=�"Od񃐩W+e�CT�S"sa$}��"O��2M͌�H���^!/��z�"O��*��_�sV���LX*>8��"O�4:%,�/N�(aƓ�T���"O�ؘ���&DO��1UL۽2	p�c�"O0l��cL9;"�=��̦vɚ4s$"Op�F���0G�Ĺ<¦h�"O���ѹP?İP��I;w��b"O�0��7d�زR�_�o��7"O��h&�P.���?3�z�r&"O�%�P�+2f�#��E���c�"O��06bԍLN�<x��ЪiV΀�"O8y`Q�"wL�j�J�*=��d"O��c��ߺJ�&Y�@֮#�ĲS"Of���f�4@@Ҍ &�}TIJ�"O�񡤞�>�J��uot%�!p�"OZ�Xef��R4T�v��n����R"O�����l�p�a�g�5D�Dڴ"O�)��)�6:��ɨ����K�"O�|�ȝ">$�S#���$X�"O"`�RcA�@\�*�C�$2(h��"O�a���̥[���2"Y�O�bE�'�d����E=���p���t0�m�	�'AڬA��@����9��e�|��'��`����#r��T.�=W\
�0	�'*Ȱ�jޟ|�+D���Q��Y�'`Us�ɂ�6 ��³��?�&A(�'z�T�5ǁ�SS�4�Ug�&B�Lz�'��    ���S�<����G��b����4�v�<��cQg8]�g��a� �G��s�<�����D�s����m��K��^k�<�F��?3�PHF(և:%�X�A�J�<!$� vݸ�3a)��hMj�.�J�<Q�#b�
@�"^:(9� 
)SA�<����1"���4GP�({hyrP	��<�ЦѶhΎ�0T�D4Or���\b�<���	-�h�ꓬȷ@����.	f�<� p�G �50�\U�K���"OvY����s�f`�� �/��c�"OFDs�-թ�%�R���=3d<X�"O \�d�2�����b��õ"O��s��	O:�$��a^?
N��"O4��G&�i�T�;�`�"v���qC"Ohl g��Q��u����a��d��"Ox1sr�֘?�|!��֓B��0�"O����䅌q)��Y�.A�?L�p"O~9�e��-#c"HC�o�1}��X6"O@�)7"�Ѭ]�Ԯ�1
�(Rb"O��Sd 7`��@�G)Z�HQ3�"O^��� ]1
P衹���(ߠ�#C"O�T�(#&��I�t햖nd�(�"O�ͺ�a�N �Hp����HS""O,�˥��0&v�q�M��Y�QqR"Or����T�g�x�f&tPX t"O�� h� 5�"� @��R��8�"O,q�3-�6I�xa�Ҭ>�����"O��	6�N��d�x��<��"O�ś�H�N�q7�ۣ\�3r"Oz�)Sf*~4&l �I�-b8�5 �"Oİ T�H�|Ў�A�h�1 :��r�"O|-Q��M
p�\j�aR<s+I��"O<�1S���p����V��L��"O���E��"2L����~�AX�"O�8kq��,,*��`E_�
f�R�"O���u)��A�8��DI �����"O���B I.|$�4�׃�
S8`��"OV�p����-�p�P�F;1�E��"OV�9��Ӷ@|�l�F�iH�S�"Oժ�EO	�.UI�P��.�C�"O4X
`D��[-�����Ơ,��Ic�"Ol��D�]���f�ڭ	Ă3�"O⠋���~E���[�1�zlA"O�٫���:U�n4�C�
.A��"Ou:Fο#�M��G\ -��1�A"O���`D�Z���C��P�n��4"O����γ2���%��E�$�z6"O�MHt��Rl�Q�
Y�s#Du�"O�p�B�xZ���*h��D��"O0Ir� v�* �6�:ٰ�"OP���-�SK���6���&u�"O�A�4n���2����S)�R�@q"Oz��A�D$}��� _tð"O4|�wa�m5ҁ����+
D��"O������1a��N�H(Hٗ"O���`/|� 	9��-�P"O"|���M?Q4	� ��}�����"O��r�,�4@�L��5\� �{"OFDäʙ=6�tɀ�l��8���"Or�Gm[vub����DI0!"O08 �E&Wߪ%j��S;Bw\`A�"ON�S�Λ�%�>�K G��h� �"O��B�$�>$P�L	�=��\��"O0	㤂�V$�qj鄁|Ȕ��W"O��
և��S>�=	s�Ҟ_�8%�!"O>5K`�M&i� �6i�����"O��1��	�%ʞ�ӆ�#:$A��"OR��*��h���J0�V�u�Ȓ"O|�1��'=ĩ��ӣp&@K�"Od� 梌!/��Y!�̐�r��*�"O"�X��*���EZ *�fhB�"Oލѡ��-,��XB��H�vt�9��"O� �@�Ʊ�.�V�L,{L��"O���D�}��I1 �=�ڄ��"OXB���=}��ks�W.2vVHku"OL)��m�8@�p��H�wT��"O��#��):����5HעZ�ve��"O X#)R�93��T�ح�W"O��rD�Eo��pň�h$QP"O !*�Ǟ�C�̋bDV2Rx�ذ'"O�}���er���ߌif�*5"O� X�Z`N�Y��%�	t_���"Oj�x��L=`��p�v�S�T^,���"O�!�+��<Z�:C�׍Fa��C`"O 	���ѬF��<Q��9/RL��w"O�m+0��S���OBjCV`zp"O,��@�B�-�|؅�٠d:\e�"O1�҃ɾA�4-����
H$舋"O�
�/������
˽���"OQ���l��	t�`��"O�%��,�K�9��Xp�P��p"O>-4jM9S��}+ >����R"O
!���		=���%�K�<E�0��"OZ	(�*��l#b�ʑg��"O�
����jaZu0J0��p"O�m8�`,E?0�ʥ�R�90Z�K"O&�H�MN�.P�Hy4�T=q4�}I"OΌ#E+A�[�F��׃W��n9ڀ"On�ɴG��(��`"�� s�d��"O��z�莫UID��d�|�@P�"O$��pK��R��,�i�`�&"OdM�� ƹ�%�L"l$�H�B"O:��e�K;u���狉3x4��"O��{��[�'��,W*׺s,2�c"OΕ0�ׯv(K�j��:�#�"O��+�Bʍ�	Αz`X�"O�dXtjI�~ʨ2&�JZ��]ӷ"OT�y�M]�Z9�ā��N5&��"Oj|�!*�+2���S�-,���"O���dy )_
��k�BX�y�M<�8�n��S�V�p�߹�yh8\,����r�JЃ��Q��y2��i8���ȵ$�N�d��y���Xqz4)��ǦJ���be�"�y���&<��/ǖKwP���yR�߰f��=�뒮C�<���bJ��y2K�@�TBQ�:�Vi����7�y"���]��=Z�o	)c�����y�+�B͒0��&�z��p�c��y�-��)�cюJ1"�L�cE��y�īX�2��¸aP,�f��yҫ�Vv�X�Ǘ�X	G�@�yR�6�XM�
N�A�X!���%�yB�ưf�JE��E�#D�F�ЁJO=�y3TB�Ej�?`v#q���y2��+���6`��sqI��yҀ��.W����&^�:I�P��,�y��Դlٞ]�B�5N��m��ϕ�yRė�{��-""��s	r`�n�.�yR&��_�$5:��X2D��y��cO?�yR$L$y�`A�J��D�~�p����y���15d�0�*��=�"!�P/P�y"N۲+�@�	��șd=��[E&��yb�b5"�9V@��^.!+1�y�G�J��+�/\|y"�iECY�C�	� ��!1��5ךԐ��A:�BC�)� t���,�|j����?����"O��%�>=ؤ��V$\,�2�a"Orl�n�$5�t�J��N:JZ�"O��"���p�Rv%AH�	��"Ov�����`ڒ`�N(&Yɧ"O����gXH�҄�؄|�.D��"Or��EE��d��)��١X�txC"O8I�����x	���v�L��^Ȼ&"O2	��S�O�$- ��A#� l�p*OhL����o���r����BϞ���'G�H!bCפv���#(��;��-{�'I��I�LH�2pԑKd��=9�
�':x1�m��<ElE+S�9�V<��'+�����­s��\9ff�����'��S%č&3�]	0萼p{$���'�J���EX�>Ƅh��e��q��� �'�ZCɛ7pT�"��˄��Y��'*V�I��^&�Y��g�0��t��'����%�̂\iB\�6+�	3�@X �'�@���׋O��lʶ���9�����'�|��w�G��)8f�ھ"� c�'h��ɕ�
�]z0U#ħǭyW$���'��UHp��/`��x��G������'E����� ?s&�R�Կ�^u��'n��2ER�n\"��E7
0���
�'j�${3N�ʔcc�
�J� �'�,p�S�M�.���E�;rf���'Pp�P&�ٮ.��C�/�3K�X��'jr]i6ȏ Z1X�I�Nt��' ��q6��7��)J��ɘM|p���'��!�%Y���"�o�-<�4���'!���LN�&��Q�'�P0�'����5'R���Ğ��|8�'�H��M0^��7���$X�'�*�A�9'�
���ߛ?���
�'��&厒"��Pꡨ�,x&�	�'SV�Jr'�$6���V�Z� 	�'lH�q'3\E����B�#W@Ry��'=B�2$N��9���0��p�TI��'�Z1�B9�\���B��}6z��� ~$!PM� �Xl�����}�����V#\��A#M�(t���E߻Qs�ȓ^'0M�@��	V �I����-a�	��<�
	{��Wc|�Q���".G�Ԅ�{�T�Y�d'/��]�tj��eqꩄȓ-�����,�/U\���B0 ,��ȓ2�t��Ӯrp�#�	)P�u��M�^��Ѭ�=
�,���ɯ\Z���ȓO�F����*_�ppV�C%�D�ȓo[(��'b��5Ӓ�y�CG!U�5�ȓc�`��!�+3��+��`$j��*����$���,��Ӏ�v���4��(���'d7��c'�Ư!�hd�ȓU����� +�@c��2z݆ȓu��(*�+�{F��&BzŇȓ6l����XZ�s�W�r����-I$|�D̓�LM p�gm ;����KŢ�ڴN�^ؼ��wĎ�<����"툍spD��	���@�HO-譆� ��L�3  Y��P�)�8�6��_
�M����MZ%�T@T�ȓ%�@L8�+Y��b�Qь��[����ȓm^�I �I��|?С�#)^�Z۲����Al�PpE��1 �4�en1D�� 1j0n��ydP�2�G�0��Y	�"ONYP�n_�R��+�+\֒��"O@"�& �)�
��ve�����3"O %;dUF0�F>����"O�T�T
k�)�D�ZsX�r�"O0h����A>�`�-s���"Oܼc'�O��f��9g���"O���bE׭SR>���▂ZI.�u"O�L!fa��b���Ѣ�B��&"Oƍ�t`��m=�ಠᔬ]�����"O���m	=q�jT���ֶ�}�"O��Xѫދ׾�k��
4�(��g"O�%R!P>���CR�� Q�Јc"O��C(ÆL��Qң,��_x|	"O���#ŌY 0q0���'e ̢R"O��iyu��:�C��.PZ �"O�|Q��48�������oA ��"OT5c��G�ju���!�DO��ce"Ob[�%!��)8�Ь>0��� "O ��d�8����A�'Jn$+�"OJuJH?FWz['N��2L�u��"O�-��T3X=�dU!"�"O2����0(��5H <0��"O����-�Jt�4���S�z�$�"Ovmɂ��	/"M�է���V��5"O��CB��?-��k��8��Y��"O����LF�Y��I@��F::�D!��"O�����@�
[����V�
Ɏbf"O�XI�#1/�03K���أ�"O�8Q��[��*QeA�rXi�"O"���E��W�D�ʳ�ڈcg�塠"OU{�c��0$ku�G0Y��8��"O,�B׊�$��ڃF:����"O�(����0<r�K.v4PX�a=�7�zH�lČ+�E�5.B��$�ϓ|7�`�Fl�3WbR��O� Eh=�I�mń8�?E��D�6��]'���$ӠH�ē7ZLF�`K�D1�nɧo��V0+����~� J+YB�)��M
Yv��p�(ҫ`���5�'Kڠ�u��'� ����f0T�9A�:h�Rġk�r�a�S�����ƈ!TB��	'�"jTm '{Դ�WG�;]��$� F�Dz�g�}t��U��П�Ґ���N1�q���/�����h��(-��\p\~��B�'�8D��Q>���O��iNU��)o�-�R�/��̂���:�(��ƝҦ���#}�r@#�����CC�<�L�;-��9���}8594D��0���}J|@��Q�&��	�]��܀��F-���O���ѕK��8�lІ��<�-cFˎ�$�r�"�Q	)�Xe�sK��f��,@"�(���"�5��0�b%^䔍��`��]t�Ĺ�cO3-'RU�Un��	�M�E�[<>��O��許 �9KyN��w��I,B̙A��
p����T���Z"�92a��_#t$�����v~�zC���1JW������@n�E���	�?7��>�2���;�
(�a�Ҽ82<���C����V%ypf��>�����6BM��H�e�V0JA�?D����֋?�x$C'��"z�:R�D0D���UkM1z�rt˗$�.sq�`�6� D�`���F.���L>��XA@:D�q0�U�gH蜲F���Y�p�8D�x�!Մ$KU�V�@�!�0t!�d�=V #s$��{��2����#�!�Ǯh$��r̖(AQh�C�M�!�#����F�%�-��ʕ$E�!�� i@��(1)G�5mHmҰ�Y��!���s�)�h�q1���ꗹ|!�$#*j �iŚL�^�X�K
�$!��I=!�����2.�����ϣX!�d��N���B�]��(��
0�!�G�EQ�`T1u҈{����|!�D��R��%� S�2���sǎ�!�� ���vJ�$[�jQH����G���"O���i�8�;WO��8$�"OT8B�5$B�+TÔ(�N��r"O���MG���#��9|���26"O�����0l[r� pD����"O<��G�C����_O�y�Q"Oq2�W�e���"r��4/�À"O�� *)��m��EK�cp��4"OP}�
_ww�1�o�
Pp`3"O�P �ҷu).)�e��&��D�"O�K��×3�fU�+Ww�J�Z�"ON����ݑzך	9�M�>2m2"OtQQ�7pA���֪��c;z��"OPa���O���f,��00�"O�XkBf��<E4�C�Kw���'"O�YcGK|g���]�^��!�"O,0���#i��8�M�n�bP"OP��OL�E+l�c3�U���"O��9S���n�����/>�T�$"O�� 
ёDtF�e�R�t"EPT"O��"�4Aޱ
�낓d.�9�"OJ��[��:D��&���"Ob�CD�e/Mh��L�
XN(X�"O@|8�/^���R�R�wT��2c"O؍ʦ�B�f}^�Ѷm������"O�< G�)!R"�X �
o+��J$"Oڝ�'@�9��I��⌵� �"O�$B�ȏ7b���6�*�Rˣ"O��S���%Ep�c���F�,x�"O���eo��<N:���R�1|�S�"Oʐʳ	�?��`�E�R�ul���"O�A�4"��]�tdz��1�:�27"O�42����Z�$�;Kҵ��"O�*�̌.`gZ��A�M*F"O`�K�%	�_`6��d��!L�m�U"OX@rDY	� �'A�޲x@�"OL�*�)�P� �/��X��e��"Oz={A�φ_.�1��V;I����g"OQz���@vRg��3v�f$�"O�U����H�E�k�|��li�"O:�Sq�E+H3��ӪD���r�"O`h���O����	�!|t(�y�"O����P�0u� ː!ocRI�""OTD����>Fģ��,(j��A"Oc �NWv�J�怵a�2� "OⰻV�Ӱ3�ҹ���*o@�=ۦ"OhtkτuްXk�F�*�{�"O ��eR,Z�)wf�bn4@"O��e�KQd܋%(�1I�V5��"Od��Ӌ0�v�*�H��m���x"O�t"�p7H j!Gـ1f�]"�"O�pXè��E�~E�t���'�j��|��'Ƹ����݆e��A�JVj-p�P�'{|0ٕ$�7+����3^����'%j@*̊kH� $��P���	�'���j���.��Ȑ0�K�n�0	�'-6$˗�!'��K ��z5����'�Z����΀WLjuH���q��{�'{:l�c"�9N3.L�FF^��P��'Þ�zd�tu��ud��Ap�B�'��q�NTeJ`т��`7V�P�'���(�g�d�wQ�RU����'���q�ǒEy[G���Aު�Y
�'���/�~)����\�2��$h	��� ��H���:OJ0ʖ�
gQ�YjA"O�(�
�0�G �CQе8"O~�۔�N8.��Zd�M�B1c�"OT[�`\?	�jQo��T\�'"ON��%�E(eH���@Ҡ=(�"O|���Z�80*��.H��܊"O��9�]�h���J_I��!�"O\��Ղ�%N`	�郒q�r���"O�y�U�X�=B�=��K?�n��t"O8 �&�F�A��:�ǣ\jC�"OF�Ġ��X���0��X2��"OzDQ$�.Oؐ(��EV��5i"O��AeI�G Z��&�(Ow���"O���šͶ4�d��%#PT���"O��G@�XC��i��εc����"O6�
䃊�}e$i�a"6#���a"O��t�=fS&�p��� ˵"O���6+�?������� )Hf"O�9ӓO�Zк�h ��8� �a�"O�+�iP�7 �F�ȩ�`К�"O����6Ąs���!�B%�t"O(�2��F�0���́}���7"Of 3b��9�@���,[��.�A"O-s2�]���"&�ӧv�x��"O��V��	��vI��[�p�"O��iDFE�&�p�?0<�a!�"Oi)��?|��`���9�t4"O�T+�Z�$K��QP���i���q�"O:�����v�q5̈�G�p)�"Or�HRaK!T�|)�"�F���T�"O䰙C/0�@MX�菹o��,&"O���/�&iZ�8t'����T�W"Op���D�E ������5���j�"O�X��!��.?�L��͕=���qt"O��a�Jd�p�K����+�`P�4"O �'���j�A�1G�)Q�rhR�"O������:fh��f�{�8��"O0p������Ã#̼\���"O6��ǡAqlcK��92e"Ot���m>PN���(�e�x��"O���7O�Y� 	W9Un�a��"O����P�#J�C`(8:R����"O�4�V$Y�D���G�On)��"O�@@�G�K����<H!D��6"O���R���$12�('gn	f�Q�"O�ʲC؁Mvf0�D(�S%�,��"O�e(#D8'o�AI��~�����"O�KV	Rw��[.�Y�fLJ""O���SK��[v�C���&����t"O�9ĂS�� ����#Y��Ab�"O�D+�B 9!̰▌�$'c���&"O~,�eI$9��� AЉr6d�2"OL8v#Pn �IP��ļ��@��"OƩ5m��@�F�kƮ �x6��`�"O�]��U/(zy�����dD	�3"O��I&�P�����%��aDԊS"O�x��,��$u1T&I�Z�r"O@u����%�	a�	�A�x!
s"OP��j$l���Ùd{�Aw"O��F(�O,�%����x��	"O$ ���&Dez��`	8��R"Ol:5�id*aAt�ț9���3"O����K0\��k�k_%E񞝘�"O
��A�(SEhՂT24��s�"O� �1�VA\�O�N�BlI0t���A"O�91w�OGtr���Zdj�)�"O�L�3kY�6��-����
Y(�&"O>�) IT�7�����	C/{XP��"OBU��*�$?�����.٢0(���"Ob��OE3�R��এ�K$
P��"O X��Ǣz^�xiÅU�|@,�"O��#�(�"C;��PC�D�� �"O>-�nͷ-p�c a�W�ܜ�p"ORdk"�Źw/��Y����"OΩ��!M+���C�ݢ2p,92"O,�ag��.F��#�+	-oL���"O�%�pǖ�E��y��KI�Gw�4�"O^��Gc� "���!���X��A&"OM��M�ZWJ��TGE�sNɐ�"Ohhd��j\��P�X�x��8�"OД� �Ў<�!��QMH��{�"Oq{�Ƌ�7����+,�4�)�"O��¥,I5=ȱ��X�W04i"O�I�S�%X�D���>Galu �"O�Q���EB��0rA0pZ�"O����Qx 2pEE,]T��"O�	JՌ�"u�%{�cʋD����"O�=ਕ�~˂��qB�C�"�"O& ��"J)MQ��Kဟ;~�鱣"O��B�B�x(�E�0�X.Qfm(�"O�xqhT�hq�g�:qB^�W"Ob+Ƭ3͈t#�&�:><�4"O�I����ڶ���D�-�fI��"O�%�2�Oli�3A�4Z U��"OZ9bG��A$��,�L��Y�"O �.����V Ap���ka��l�!��3d7*%@��_-H�	�CHƒ6�!�d1 Dف�Q(E'F���I��)$!�d@�1� 0Y#,�H�lp���Z�?!�d�0@\$�C˙�`�qB��|m!��1��P`L�/iy�x��JA�	X!�ߒ,�6��TiΥM�ds��ȱB!��Y=�t ��ӭH
�=����B!��W�<���J�� �=���,̀%�!��L<��Q�$ph���	�I�!��e��0A�ON�@�,ǝLP!�C�M��p1��$:�PXz��8P!��qE�c��H�.��,����2JpG:�t���B9�����	֤�I���3
�t�c��B��\L��,Ն<��I��{l�[�f�Z`h�ȓ3,2�hf�[��`�Յ�dr��èԃ�D��C�,%�ȓ;墀�k�o��Պ.�:~�P ��2\���lΡ�h�"p���|�bu�ȓVj���wh�Y+@iX  W�6=,�ȓKx�9`R&L���1���ȓZj�a��C9�����) <�-��+�qRf�_������C�g��܅�15�uV�Ā�ꭡ`C[*/����D2�p)��'wI�����$)��)����*R"qR"�&��чȓ	�R�8u�˘-�6��醡Ub ���]��=[�	�m�yжG�B��1�ȓbf ��-j������0��ȓM�Z�	��-�Dի���9q��ȓkm�51�[Q)LLZ���6+�Ņ��N�� @�?      Ĵ���	��Z��	�3V���C���NNT�D��e�2Tx��ƕ	#��4"�V����c��mZ�V�D3%K^�+$�ʡ�ښ�ePĩ�<w�����`#�Mc� Y!��n�]��i�;F�hxۀ�'���H��,�ڰ"�Ă18��pY�n� tR%�2�
dy-�!�dp� +}�VC>�*�#�SGt��֣M
K*��(�;`��X�'R�D�C����Y�*O!y"���`���_��[6��)*-��-���pۧd�m��=Q4+C���ɶv#�`	IE����n�ن�ȹ	���Ѓ#�'Q��<���A�'C�$�fl����f ��L�D?	 I�U �Y9pH�'*	�4�B.�e?�u��~�,PH<yË��|BH|���U�9����C��;taN�R��=[J��)Y*��I�'ɐ�@FΒ2��I�(�T!��Ϙ ���pː0tl�P�4@x�I1�?��[�kIH�$���`�oWtʓD�$�Geڡ:@	���6s��ɢ��i�G$7��ۂ�K��'F��"cB٤F����/� Gl� ��ɖ"�'���T!�
:��OPU:F��"�&
�#9J�Q�H�<��� AOʶ������ы�U���Xx	�g�w�P��4.&`UEˁr%�p�4��������)*(G��O�j�}�|	Y�a�J�	��?���"	��]�rgւ�$KW� �o�4�BF�:��`�ڵ�֚|b'�l���H�'\Ȫ�FC�ʌ0���D��*+O.�0�^��(OD3J<9W(�u��Q�G@�=U���a�Z?o=�
@O(�!�4-��ߕ+"�3GJ�k���/R�q�Q��`�apX���-� �'�)��`W�/{��dދ�4����.�6D �N&�qO��M<u�E*�D�M�<
fN��t���� �^=�LX�L�A׾S��0��ϡ>1�9�w�DУ~"�a�g��>s���Rb����U�,D��A��   �� 8�Q�Q"O|(���  �@ d  ��gb �  �4�[���.�Z(���;r���I+�Qf�'jnIa�[�?3��J���M:V���&V����;v�y� H�o�I��ß�ntd}��wIb�z���|��,I�ks|aG}C	u�O���p*�2E����c�MQ�:�r�'2��H���`��b)HP�0�h�'F��5	�YiJ2r�ZE. ��'�1�v��p�+"Y+ST"p*�   �  �  A  �  �+  �5  R@  XJ  �T  (]  ,h  t  �z  S�   �  X�  ��  ߚ  "�  g�  ��  �  2�  s�  ��  ��  =�  ��  ��  n�  ��  ��  }  �  | � v' �- �3 "8  Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�� |d��"O
`�(�;���8���-0��1%"Oj4��ND^[��"3/9�0|H�"OB���H��*�ʞRy=a"O�味V�!X��!&F�:J�$���"O,��a
���C�Ą�M�"O,$3%o�-���p���+Ն�:1"O��ݢ1����`���y14]2��i�<�6��{_���c�H�`�fX�$Kn�<��A̼VI�xR[�)�Ć�pඤ�ȓA5��('nߡ4�� �)˩%� ���,��r�؊b#`T�eT09���ȓ!�b��g��}�8�F��-? �ȓ
K|m�ș�VṔ���2�%�ȓ"R�X�j�4JN�1�˘X�i����̹	_�jZ��1!g��zܶ��ȓgil,*�J�
j�Ne��i�J%b���f	�(U��:���G��$Y^م�~r�� S�%T"���k\�jx�ȓ|4�1�îJb��@ӵ�ݩn�V��/[`�"�v4�R�!ʎ<��M�ȓ`:��z�ؚh�J�Z��$HY:	��H��p�m�C1��!��B:��0��EnjZA V;9����J[
2���	��4'J�EA�IVW&��~�(aZ��ӹ�>� o�Y�|�ȓ�f�A�
Ο7�H��M�$�����mޠP����/���ANXo*�ȓTv�����{ ��-7�*h��I��sB�8�8���3����ȓNe*M�悡;������X�o��!�ȓ'lj�#F�m�+R&;�|��2)n�C��0S4���T:
b���:�0!��e֊��)��ͷV��,�ȓ0�&�8#���� ع�L�����;�P�AFd���,w�6d��r�EQ�( �gVlɦ�M,H��,DP���|�I	$G#\���ȓ"�)���E�B	yt&B�^�LɅ�4�� ��eëF�ڙ��n��R�p�ȓp`@}bŇ�=�$�AUN��P����L��p���_�a�)�Y�!��-��u�5���o}�`iF�@A�p �'Cў"}�ɃJ��ӗ��GT��DKKv�<Qb�ʚ\���'$�QI���M�l8�xS�� 3�L]`#"��m�d���$�O"1��}t��qș�A"F�2�Q1�9��*Bh�4
�=#�����A��]�ȓ}�4t	$e� z�`��՗f:�ȓ\����!�U<Ed�`�!K�fVI�ȓp�Llk�%�$h-�(�e�}.Q�ȓ�@!xdOZ�Zn.��!�Z
�:�'Ua~�O=W� q# [ 9�r�������yRjK�U��ᄌ-2$,-����y�I�2�[k�!-\��"3�y�&�1��e�a��*r&qab�E>�y���
F�:�0���q�܄�!$ԻIj��=E���`0ze+S�h��$H�w&Y�ȓASN�5a޵�$��'��\����3[�)��G�מ0���r(Ȅȓ?5t����һm6�0ϝ�f*.��ȓ)����`E�	&��mBS�v`4��S�? *8G�#'��v�^15�\��w�|R�'��T;B�I�%�j���'��M��'0����*��0�0@ `%0�����'l�@�u�N�`|�}��n�%�X��'-���@��5�Ж�[#T	y�'�ư��!ȧh�J�����B0��'	f`H��GM����o�:¾1��'5^԰�%A;t�A��wZvi�
�'!l�iT�ݧ7?�i�	
6p��$���(O`E(A�V���+��ۂɊ'"O��e�@�P�X�S%�F)<D���"O���	a�-{D�[�Eέ���'I�	 Cd�!c��0"��ʀ�x��C�I8�h���ڏib��9sJY-~��#=1��T?��wo�+M�2�8�l\�2��%G&D��bӈ$�|����z���`/D����\1��A�*�|v��(Ԭ(D���5�Ɲ[d�)��ԩXE��Br�)�D9�S�'9�^����bk,�}�r��K�<!�$�92`h+�UjATa9���J�<��5s���I��I�R���)��|�<9�̆x�l�kf"�ν!Fy�<q�-�(
qI�I[�P�^xY2��Y�<Qt��3���V<X���҃�Q�<��$O4fm4��ON8ldzi`�.�N�']�x��%>
k��]�]��H\��yrl=n/LCw��8�Je�����y�ʞ�a"�@��Gy�I�Wi[�y��>��J�/D>]�\�('��7��d7�O�"�nL�[.��+�k��U�b����t�'���{��IjE�̭R��P��ʗ~8���ȓMc
{���>p�4�C�B������	v��?���.B��h�lG�P�����S�<A�m�8PHr(��@G-o������M?Y�4�hO>;��U�|�8��4N��`��ݛ��"�O�Oz��ㆈ5�&��hިBd���"Ol|�@O�kW\��!+6G��u�'/�'�xPp�X"}j�3P���,uz� 	�'�p�$ˈ5C�!�4d�@���(ORT
��@.���*�AQ�ؐ��'�"�I-�.�r��BXl����/� j���OJ�=�}�$e
�6�H��C��5;ڌ����o�'�?�b2�(o�"�h�-=�͢Pc:��gӾ��$ώ *h� FjF�YI�Y5@����=E��']����ˈkZ�|㑯�MY�!��'r��V���\�ڑ�̺v�jP`��i��~ҡO�{1�x#N^38�20ʙ6�yrj�3f�uRCnK!���`�,�N��<{T^��F{�����:%����(ċz�	I��yr�-���n�S�;l6$ 1AA��x(h�NOT��C�I(sAT�1R�Q�
L����<�㞈�D�)RL�,
e�qX�,#S�p�fF�#5&C䉙DgB���X�<UൂfI��>�E{��9Oܒ�EO�PZ��1�A�.d챲v"O�� ��$��,3ǏD)?<�V�|��)�	"! rFڞ4fz�� ØuI�6m �S���ě�&� �Bqh�%B��1`ϭ.!�u݄��wfY=�p���� 2M��w�'D�����̘�?^z�˕�G�,� fJ&�O��'��)S�^�\�I��*9_�%�	�'vf�{�@Ȃ=v�DV`V�<�^���'ԀmHd����ɒ�ގ#����'H��s��Bs�q2���Z�r� ��OJ5�
��3p�iuoJ:i��������Vx�� &�x�XQ������?9�dYs���:\O����O�IQ�x�����h��q"A�'�'�F0�טM�6P��3j�h=`�'���@:`�9cO���E��'*�tc0%Y�t�)���4�Px"AE�H�t0g,��b��G���M����?E�=i'I�.�|L�Ѩ�,'�Nh�!��U�<yR�ˬ4vnu�3��*R��Ak�a�v�<���D�<|	8e��'(y�9�a	Dt�<�SL�-�B���ϙ�U�b![Q-�r�<apD�|舘�BIE�2-688�HJ�<��ʙnx�5�F� �N���Hz�<��'ɴ'&Bi9!C;e7ҹC�M�x�<QЦ�7rr��͕4et\5�1���<��\-OD�A�/�2&T�����Zg�<�#��4%p�pR7f8��^�<�qꇔJ���kP̊?FzT����]�<��a�qsn5�MZ�98��W�^X�<�����n��5�$��Ep�<!��Ԡ%��l��\?l��a9�@�<I���*t���6eO!:¡z�i
.C䉸xࠥ:��O�9�p��$φ;1�*���O���b�O��D�\�@aFl
)e
�aF�!��P�@���W��ap��&��{��K}��)��IK�8&��D���z;J�4���hOj7�+�Z���i��v�!֭�3HbP�ȓ]��a�+аJ����hZ�h�ȓ6�V�pg�\~�����;L"����n�@Q�l	� �PH��/Y�.�<�ȓNF��'bѻ5�t��Q�I+g�fE��)��w�����B폣+c�%�ȓOa{�n�U��L���69FD�ȓy�l,Clks���"@ȝ����4�����K��I��*,{�хȓ5h��Q!(N.I���s�Y�?	\نȓeB!�%��;* ڡ��,�+,k���FoJ�����auOP)c��ȓ:TX	�'U1O��"Q*P��d]��X	�����Ъ�\���*؉4�؈��Ц}pb ղ{�>t����0{Q	�ȓ �v�+S){4TQRȂ�*q�ȓ��@h��  e�z���,D�b�$]�ȓZ���@:(>��f&�q���ȓj\�y�&˩a�T����8����qn�{�ȱ[u�J���/a�ȓ6���{g#�7����S*_ղM��U��A ���,V��*a)�>����y~�ͺĨ��csyj� Ԓ_R�ԅȓU�BD!�J`��e�v��@��ȓ�=�GQ��=��c� �����Y9R�s�E�fl��a�9D ��+B�I���O������N�9�^ͅ� :ƑC�T�<x��q�S?]\L��`�Ƙ�Wꆪ8��c�	:v�\L�ȓM��T�n,OZ�
�e��rWl(�ȓu`8��zr��!��kW���ȓc�J��џi2��2���"�t�ȓ8o Pc�	*/�)`�,�p������lZ�� <�p�͐u�<��2��qQ��%wK�ի֧�'?g���ȓdu�E�,]�6L�C^"&4Jh�ȓG���%�ؑK�T��ԡ�9���T0p$c��	#C@����n
'�X$�ȓ~;�I��"|�z�GT5����S�? ��+��8-x�@�GT	b��#P"O��Q1Ϛ�=!�]c�+#�p�ȗ"O��"������)��mw�)`�"ON<`u�(cȌ8yG�)f����"O��e@�L((i��w��Q��'��'���'���'_��'V��')��SK�QCTJu�''2-�V�'���'�2�'���'U��'��'�B�@�ᅶ^�hј`�V�ɜ5���'��'�"�'��'�r�'�R�'dNi����P�
���t�x����'�b�'e"�'q��'���'��'�JM*��݋1�L /ݗ\%����'V2�'�2�'r�'"�'c��'V�� +8�pL�'F�٠��'���'���'jB�'L��'<��'���˅I���*�hdD�6�'X"�'�"�'*2�'���'-r�'8 ���[�U�ZqiS���XA�X�#�'B�'�B�'5"�'�2�'K�wzTR����Y�FM��	s����6�'���'��'��'b�'���'�8DS�NY�}Z�-y����A'�QI��'�r�'�"�'�2�'L��'-B�'�$��ʉ�I7fa���M�5���'���'�B�'��'��'r�'��y2ċx�%@�ůQ�Ba�'�R�'�"�'�b�'nb�'���'�l)0�ς9ԴX�D,�xS�'���'���'r�'���d�\���O��
����| Y�)�����G%o��Iҟ8������Ѧ��#i�2�잹M-*4�U�ئ_�$�Wٛ��'�ɧ��'Z|7��s(,hb�,u��j7F�JҞ�mZ���d��Ҧ��'+�%_1\���ś~J%&W8� U:��>cV�!�`(	v̓�?�(O�}z`@�s��2��;8or� �"H�$C�v_���'�X�mz��[����"z��q"�P�0e$Y�MӢ�i0�d�>�|�g�	��M��'%BC��ϛ*��ȕ�O��*�'��<�R�Y�`��ea��i>��I[w���%�u�D����wb&�y�[��'���ܴEb*,�<�D
 l�tY�P+�t$h=ӣmK���'20���f�v���f}�K� ���#@m��>r`��q��-���߀3r\�pp��sp1��� ��i��	�X�\urAN�',;*����1xj��-O�ʓ�?E��']2A����d�n���oB?m,�d#�'�
6�ԍrW�I��M��O�yR�Nĭf��e(rZ�h@���'/F6�����Ɇb>(�mU~�Zo8�S@��3%dr�(g�ѩNp�-�q\��iV�|BX����I�T�Iޟ����=_�6!�,��B�&�Ay��l���:O�D�O����ą�2$�d�E
.Bʾu�@�	)����'�87�C�}�I<�'�z��4������^$#�L�JQ��.S]z9�" ϏF�2=r.Ou�Ԃ���ݣ�����|�.�x����p�P@Q �;=�8�d�O��d�OX�4�^ʓ>1����ybk�I��I�蘢x�*%	J��y��i��Tk�O��nZ��M+��iٖ�	�%
�[T�|3�c)��U���(L���:O�d��:��t�G�?�����V�A�2��� D	�\a篈�~��\� �P&j��qN�l��8	V��9d�5x��J�0���	�K�f�	'+/꡸U��0�*��^K�����F'*,���L� �䬊S��}���0*As����ˡ.	(�������uK�<��LJ���U�m��(m+X�"u&ӟrf�`���4�T��m .\{��'g�`�D����Ҏe�n0b�$ԑn^~�&��>����nK8qd�mk �Q�vXl� �U�Xgt�{w�n���$�Od�dX8a���%�����|��1W��Q/�0?!j]��.,5#���>Ip���?A��?A��ɔV��a�-��8!:5	��������'�����H$�I��h&���4h�xy1�Iǝ<�n`r��L=8��Rj�p�<����?�����$��l;��!��#\�1�O�"�&��Cy�IҟH��Ɵ8�'H2�'"m���8i���Ac�!�(��E�7Ϙ'�b�'h�X�X8%����t�k������*sVpA�)����O"���OJ��?��6��O�4䊇��d�����Eē�>�@�O��d�O��d�<��#k8�O��@�%�`��ek���6I��R�Mw�2���O�ʓ�?���E�V�~����g����Cɔ�Z���@�Ӧ���؟��'�pq��+���O@����Q��7#���Jяޓ7v�j��i�	ʟ��I�p"|z����ʌ�`�Јp Su"�B�h�\˓XnJP($�i����?i��6�	,i��ܚA��Smn0��1y�7m�O��dX����S����ēi�$���C,{�!� ��>}Z�l�(�@���4�?i���?��'�������i��@[��,a�q�� �%�7M�66h�ʓ�?I���<	�@u~l�t�g�zE���ܝ'(�y��i���'�r6�PO���O
���	�=�q�Z�q�v�D��'?��'.�e[�yr�'0��'��ڇ�X�8єΌudHX�4�p���DT*3��%������IYy��ͭ����G��1�Lq)ði{07�O��j���O����O �?80l2aEJ��  ���zn���"gU�'�b�'��P��������tb˕E��"��K�^aP%�',Y�b�L����I`yR�^�\v�擎y��i���,|�` ��QbV���?i��?�*O&��u���4X?��%�}I�=���A�>\���@!�>���?Q����䖉3"�<$>}�� :�b��{��d�S�#$��`7�i���'��I��0�	�K��b?	�`�4-�i�ݞ-_bxbb�|�h�D�Ob���O� S3�S����IΟX���?���B�Q>���쇍c����*��MK���d�O2�@�9�>��<��A@cf��+PF�����W�v�'�-оRk\6m�O��D�O��i�t�$�:H�1*�-0,� �s�ڠCk���'����s�R�|�O��'��s�)Fyő��\�[DN�mڴff��9�4�?y���?��������?1�[����,��%
�5s��R^��YѶi4l���'
bZ��R�ğ�zL���AƁF;<,�QӓNH��M���?)�h]�I���i:��'��'�Zw�A�WJK:}x��rm�/Z%P���4��d(Dt�h&=O�S�?��I۟D�g�,�\����~��� K�<�M���	�`�Q�i�R�'�"�':��'�~�l�]5���##��v�ibu����H1����Oj���O���O>���O�|�b�5c���D��v�@�>�m؟��	꟔�ɚ����<!� ���*��Q a㚴v,��
�<����?����?�����)�?Ӧ�n�v?�h�2�P�	�Ыq�D�"�R�4�?����?I��?�(O(��V)e2�i�5ꠉ<v"��CmÄ s���O���O�$�O��/�8�m�ğ��	����  +��O?��R�h@�b�n��4�?1��?�/O��	 6���O��IJ��)��˒�VY����O��6M�ON���O�$W����o���������뺛d��1��]�V"f91ԍӮ���<��VFP�ϧ�?�-O�i�h�+�'4-�u�ME����ڴ�?��`�N�!��i�r�'�B�O|�4�'��5AV�{M�`)��/�p�Ƴ>a�Y$�Q8��?�(O�� ��C=�����P&�:	�BK���MK��U��F�'�r�'��ԯ�>.O�i�'b�	N޽�(@�A:�A���˦�$K!���OUB.9E�`
�*��D���1��8�>6��OB�D�Op�@��Ǧ��՟��I֟��iݹj"�!+2�����v�>%�
gӴ�`��\�B�S�d�O��'S��2境 �
�Cwň%����UHy�L�䝈`�^mZ����˟8�ɯ������իQ�b=���w䐼w�^�GM{ӄ��#�/��d�O����j���O�˧h�Z]�Wn/Gf��􁅅]����R�б曶�'h�':���~�,Ov�d�"��		&#߰=*��ȁ] ^9j@:O�˓�?a��?���?QD�#���Lȃk����@��	r*�#a&��zZ7-�O�d�O��d�Ol��?��&��|���V@� A� � �P#�Cɡ)��IӟT���H�'<f���=�I�`C�,����R��!�B���,@lZϟ'�\�	ϟ(�q���O����H3G=����l�,*H�ŵih��'�割puJ$[O|�����ΐ��l݀��;����`�dP�'v��'*���'rɧ�i�2����ëOլ��4 $I0��R��CO�MKS?i���?U�O ���
ih�p^h��1��i<2�'`B�2�'Eɧ�O���� �/L7�@���b���4�����i8��'nb�O�0O���ΆOW�(j@)ϐ��|��/;N~�mژ4-���	Q�)�'�?Ѣh��u���AQoR�n�R5��ؠ-d�f�')��'T���4�,��Oj�d��0��U)TMB�Dɕ�G}��t&nӔ�O*���L\�S����˟<C���%j�ЀoW����ia����M�������b�xb�'p�|Zc���a�B[+�llڀb��2>�1�O�@�0O��?9���?9,O��`�ꔼP�2��F�9`i��L����'���	��<%���I��@���+����V�r��=��NG��%�$�Iɟ$�	Zy�,��3�
�!:`�
�oŽ 6�!��n��$����?�����?���r*I��0�	�b*��WB9�CK��J�r���]����ӟ`�Iy���!o�n���Ҡ&��=&��d��#�p���a��z�I��d�	oƊ]��[����Y�Nyh`��4if���#ꋌ:E���'\2]�ܹ�����'�?���Q���NZ2[��q��P�� �%�x��'���ݖ�y"�|��D�p����A3���
 �Ⴒ�iO�		;v��40��ϟ �����'c��H;@�ԧh:p����#(ϛv�'BHB*�O���E��b�y�vۖ��J� ��ּi�:1�t�����O������&�D�I���d��M(MXA���6r/�-aٴm\\�����S�OL�+�+U�����s�t1X�j[#9�T6�O�D�O��P%�IJ�	�,��W?�PcQ�S��z�$�*J�ֹ�%�_��f�}&�8��ꟈ���V�=�wK�&'Z�`[够2@ne۴�?��O��'���'0ɧ5�A=!�f=C�`��{� x�Ę��$ć?t�D�<����?����Z+;x��s�I��b�Ȇ6ZKP���F�I̟��	I�	̟����r�^�`G����d��L#bwxX4�Zȟ��'�h� �.��WV�a��,��oX�ϕ-��]�5��rT)7�Ֆ$�99�
ƪh��v��_��	�"�Ԇ)����H���O��!�]�F�}�Ъ�>%"\ac�K����N�t�z
�艁_���a�I�̹�#K�ۊ���)�b��"��H�,K&4Y:���
.GZ�I"&F�*�Z��ĝ>���H2%�*~J�	b�Ji�^p�Sc��|4�Tk�Ŝ.?�  �kF2)�iGbֿs<.-c D[�p�gŎIJn��H�
c�	�!�t��P�­=`���6mR��'ՠ`��ƣ^���4�D�!��9�S��~�/��h���7�\Q;��q����e�>��B�;�j�J�i�:9B���+�uW��8s��!+�π j`k"D"2rl��j�7E"j�A�>���۟h�<��Qi��]Ba����&8�l����Y�<����!�($(���C� d��)�X�\c��D	8$윑G��;m�x�R�� {��oߟT�	�� �%��=J�8���ßp�	Ɵ�]&m��5���3E{Ĉ�D��&;ъ���V���0k��l+���ӫf�g�i�L�框� ��x��H�a����u�Qm�����<��	��̄�Y���Oʹ�1Yռc@5o�R����ߎ`�����E�&�'�����S�g�	�S����И;cz�H!�\>JV�B�ɆFќy�ሺD@�*Q#��i`��
v���Sn�� �r���!�e	�>H�N(В�
"���O���O��U̺���?A�O����_1SU�B$��3��+ƃ�.�x�/R�J@���فvٸ���\�`�r���'G�����<Q h�:'B�
�]Z%���?��'nTHj�˚��B �e���;I.��'��)@$��T�N ¤��?�tj�yR#"�	?a��O��X4�(��D
b��J0�D�bm2���OX��O�Ol�$>�����y��9K���8Rm.9l:�j���X�Kx���D��`�����Y ����*4@�Ѓ!ebӂ�HF#�`N5�Q�Ȱ_~̄��'uz����?�*O�aP-]2����"C�la�9����#�O�Ěr+ܴ"���g�;QG�1��'7�!pf�W"E�r�@��D�Y��D�<�s�����f�'��Q>m�2����l�S숐t����b@�s<��K䟈�I�>Cބ8��ܧxD����?�O��4&�2%P�����U8g��=�r�'xhu�sΒ�OyU���ڿ�d��ė�
��a ,�$q���_f�I���6TbL]� �>�"�ʟp�L>��g^���ِg��N\�3�B�<������-|�8�B�C������$H�X��e���Ʀs:��z�i� d�� oZ����I���3WFR�Q���	ϟ��I���s�����
�U�n�VݍvQP��N��,� �`��O�Mi�QA�g�ɁYp����|�z� ��C�HP��G	/�> �D.J�A���f�2+��O��ŉi¼[���)|�̂7 �5k�8����T�5�'�0���S�g�	�]t
�[�Cխe���8 �ˤ'4�C�	Nc�t di �]ҨCFM�9��Sԑ���z�	%�&P#-�2Z7
\�@�6A>��!焎K2(�I��0�IΟ_w���'��iN�%�y��ZLbGA��rb�`QOp@�=)l��PaѢmF�b�BSc!��<�H��XG��j�@�,Yנ����'^����-�1��l]�gޠl��o�p�!�X�}jX�0a�S�fü%�a���a�1OB��>٧����v�'��#JE���:��& i��l�) j��'���!"�'��0�D][���[A�|��C4R�\t0$��0c���7��&�p<I#�͉xP$�(��*ů,8�EY�$I�?�y���+O���V�'�PO�ᣡf��Ĥku�Y�jv�y��"O��"�{��� ��ae,���Oj-mں$|���Q�]�!Ly"`�E֩'� ���6�M��?�+�����.�O���`V�Ba��ሜ:k�hc.�O��$�'� ��'�C �(-z�����'��ID4�R q�l�:o���S�OD�(�V��aj_B�!�$ޕ~	xc5��}�<)zd����M_�;v�Q��/����P����0_2�D;�)�S�~В�H�ő�no��Y�. �3:B�2	� �#n$�ȹ��B8����a�'�v܋q�Ɛ{�1!W.�v��I�Ig�����OZ��L�%����Pc�O&���O��4�樛���=:bH�%n�m�`�#�gã^Y"3�Kݦ��!�Z�aW,ȕO0$b��ĉ�N4���� XzҰ�U��4N$D���5fP�	Q�[s� �|����i.杰b�6��q.�$;@�zr���;�H!�4&剓j4���O���L����=���-,K"���4
��4�T�I��hO�S�U��CV�݁
��H�������;�� hӸ�����I�?��E�t�'�,ዷ*7/��Q@����Y�~�ɑ��z���' �'�.ם���	�|�s�w���ɕ��6Z���J���E8���b�>pkAnD4�Z���3����Y���?-# �0MD��6|1�Q�F�
=��j�O�1m�;�Mk������O����;9�ԛ���s�Y�
9D��R�KU
5J�P���W�yA7�I'�M����d�6S"l�ҟ4��$'�N���'�R,�E��[EX}�I͟��Ƭ�ӟ����|�f��h예x���[)�EKٴ	*Q�0�	2�|,�c��+EZ���	� H�ݒS/FiD��y��aKE�G�k1�9�bȎ?&�y@���9�sM��W$���&D�O�%�� �-���JeV�s��� 8���"Of|r%M�18�JVU�#��)c��{����lӦm�j.�x�X�.
+`����A:�$]�+��n��L��e��eާ�r`,@��P�RD��ZLp�D�}B�'UJ����U7�ҟ?��)��S�T_>qK
� #P�dK� �0�X�;#�*}�(aD-zt$�Y��:cf�
[�t� ��7D`�̧���;F�l[�bI�T�h��O�E���'74�O񟮬"F�^�nl2��U�b�Pb"O��c%�մD��Б�2Z�T���'PX"=�##������ e��D�P�(83�V�'�r�'�|ى��U%��'����y��Ӣ	0b�C�'ַ$7$1ruAN�4oؓO��۶�C1��'�h m�:"�z����_w��$�� �^����(��!�3���
������G(d:����ڨ&��d+?A��[��>�D�O����Z��Ȕe^/T4p��g�/7BC�	�j��t��a��g�rt��O�p��80����$F�J�8j䩔0o��偲O<�k��?6�P���O����O& �;�?Q������ɮ�\ �U�#@U*=��́
)��M��K*l��s7㜫D����ɻ�<Ę&"@�ui�D	�&(�Ų�B�kg,��c�O/x4��������K�%��$�I>��K� FC4��a̜�dJ^�8t'G�Q���	(�M[��i#�O�-�~ڵě�P�$Q�B�Ԡ�qld�<��ێ5���I�)
�]*L�)���{�"F�'��I�.�(��4�?���7!��$��yG��ز�C�X�������?y2c��?���������3�|���G0o�nY��'?vC�0�G�?���R���=��X*�BZDFy2EH?&��u�1��^�[�DԴ�+gV(9� �@���P�(���O�UGyrg[5�?q&�x"#!�2�`H]#8^�1�ǜ8�yr�٧jR��QϏ�
PMi׫ŕ�x�f�iV@ͼk��"!�t�0!�1�$�<t�4mZ៌���D�b�� �C�A�Î�5p��<�2���:R�'���b,�;�7�t����|+�@�{�k�Z��Sr���Z'�t`��>�Ub ;��@�Ä�B����2�R)�ug�@-*��X�O�k�лz�t� �E�#�H��3�*}2����?I�|�����&d"ܡ���$O�.d�Q-�;�y�j˻&~F�ɒ"�2J��Uy�J���0<	��/G��Z���}@y���B�#�H���4�?y���?�U�1m*N���?���?�;9EP��c+"$}��
r�%@ұ��y����<	��c̒�k���L�T�yP��d�[���牀i��`JVd���	6䝃�R��N>1v��>�O��%N�O�:10bِ�R0i1"O�����W��]ӥaD`��P�V��x@��4�D�OY��$�0EK�Ě�Fr��8y���O<�Y��O����O��D����?!�Oƴ� �~��|9��դ+��8ZW'ޥcH4�A�N��3چ��!�'� hvL��jG�����U���l՜U���J
���B�)+xQeʙ�@(Lh�=	�̌� ~����G]1��z6M��v:P��ƓZ~�EQ�n�1"��p�s�ʁ9��	�ȓXo��ف��n���,ν-΂��<Ip�iZ"Z�dP$ ��M����?ad�J&!Cv\`�c]y��/�?��z� Y���?��O�Ј���w���@�
R]U��x�LU�Zt��I�xz��d�w#؟
v��Q�-D�S�T�ȓ�4O(����'�R�'��hةw���H����"�AB2C��I�x�?E���-28^�����;rȣR+��xB ~�,%�*N/��u���B�jj0�3r��O��v6�\9Ծi���'��L�&p�ɒ`�U�bf"9�� z�� h��I͟`�Ao��t��k�R����q�W<��)�|J�CN!H8�D��+��Lx��%)�~��)yC�LT�� m̴T �
�2:p��$�	5D��ڴ�i�őS�@�\<KF7'��SҠ���m<N��I���S��.q^�+� ��@-2��d��m��ȓ6���̚O�*����h������4��<Fz�O˧�	6��"u�0P�۽�6m�O���O2���g�?����O��$�O�NC:e`Q�!bݮz�4���	�wh�<Rw��(Li���A�o�R 
�d#��g�Ɍ����^�CoXD�GO�;!�p�#T�a0�I�k���#���?�*�O��V�Γ�ywN�=WHl%:�AS�#[�AaUပ}�2��(��j�Oq���'�RD	�xdDt����-#l���lގ&]���C貉K�O1�(�`l�$F/�I��HO�i�OT�`�L���U�n�+�d׵Db�q���RX��R���?���?����B�d�O.�� PP�'��Xb��<������� O24����M8A��Z �E`�'E�y�&��}=�6���"�4� J�[�$��%��^Dtة@]�R�џT�.ͨI��耀GctU;�M�Y"���'�O� j]�VnH(w3�Ux�̀@�v���"OX3g�[���#�S�������Φ�%�����M���?id�2$�N�1f�q���5ϩ�?��& A���?)�O��	�R�C��@���!t�`���	�(|H�����8񆕢cџ�3�\ R~���BG� `��C��T4 ��j��ᄑh�	n? �-���4�I�$�X�ɫ$6�2�����4�V=D��C�ɀ(�4�+
����y㈈.%Z�B�	?�MC��w*fy���V��g����Ba$U)��iC�'��Ӣ����D��k��i2�\0U2v�u�	���e�S[ЙrbE5%�1��T���)�|�c�Y�s�Pu��5q&��w`�m��f���)�<}P�
� :E�-�;q�`�F�55�դ`���RL�(u��E��(��R�ZQ�I^�S��Vm���#�b��Cт�D] E�ȓ�f5#�THZ���C�P�����HO¬��!@�rʆQ�ҌgG�E���ڦ-����|��%1pt�0�$�	��i��HF�V�鑆��ITd���M�j;���牻	�@� ����i_�H�Θ�"Z�8�J6<O�УAc �4v`	��U[}P�4BD}�Y}X���|�R1-Ք݁�O�Q��d�p�@��y��LQ\`�LP�[f�D��ş4���G_���t�|�iG9?`�@ì�|i�j��Y�QxѮ�76�B�' �'1bꧬ?�O��W��t|���wDZ<Xm����g�@m��0�.��� L9\)��Y%e�_m� �c�Ð=�j(���T5�):�A�;����cˈ-\H������O`���O��D�<�����'���d�[;_�.Hx��,42a0�'0��ǐ V>�/�B06E'ޘ'�듡��_l*|o֟��9T�l���bM0|��Rr�RZ�I���	韬�I�|�$�@2
�F {Q�>Q�K�1K� 5����H��% h8�0�@��8W�<!N2��<{�G��[�"��fE��E3�U)�����x2���?�C�x�C�f"��i���V��bB�yb�D�|�"1�w�$�ƍ[��� �x�{�^\CDL+� \[���"@@E�A�%��R-\Am�ʟP�II�D%�5x"�I��\�`l�p-�!
ʒyÁA��n���'Ǩ����'1O�3?A��ڛ;k��y�Rز� ��u��̯6���?a�Dƞk�0y��
)=,
�:��8}�8}�Iܟ@��̟X�r��\��0|	A�*�2}P-�W̓�?	�͘����ۙ���A� 3b���I��HOT
Z��	�@�D�2��w����m��џ��	��3�������柰���ߕsvM���ˡ&��:���	��"T�H%j�Ƌ(,��
ք@~
��|�q�>�Q��z����C�~n!�3�Ϥq�e��'�)]�6��/Rx�큔�����ʧ,�Hu�7�~���e������)R�ۢ]�R�6n�3��^�R��)�3��և'��#�;�*�8dB�4u�!�$�+Y��ȰT��b[�q��C��_n�I�HO�I:�$K�8u�2������=@G���r��%Q�ka�'���'g�p�u���$�'9yL��ǭ��q3�,�A �4UN9�A_�|��U)4��-h�A�Ø3��O|u��l����
fc�%#l�]��ϡ#���P�+�:zC�3�U�q�6�&���t���P ���cX<,E6����jB�,pA�'`������I�X�D�͌PWִ��i��0�!�W(l8 �zg�X&6��(g�E>nP1OhoZK�Ic@ؘ޴�?a�57J�B �Uͨ����֒$atU8��?���ƌ�?����4���?�M>Q�J��B�­q�J��
ư� D
P~8��st@=��
"�}���X+0��QS�@���'98K��+k�'��[�1蜽�t�OIH$S�'���M'X�$h�4B�?{j���'�6-B�8�͹B�+~0��k%�C
J	 �Oz�!1 ʦi����ܔO���i��'M�ٓ� %!@r}) f����?I�(�`�!�J�	jd�!��i�2d􍀲\?�O|ڕ;g��A��{g��G^�<�M�34H@%?�b�x5/A�DǶ��%n���`? ��'�������4N�f�:�C�#1�p�O�ݨ5�'YH�O�\)۷��M!�@�J�9&p����"Oj��AY#W-�x�*]�|y���'5�"=y�����Lq�'Lo��)J�0I�&�'�"�'���7�G�B�'����y��K2������G�\}p���R�<�v��7 ���rGo1��U ��)=�DVgO�G�V3����MH�LZ��q���2F������ ;��蹗�^<駸M3���޼�0���9r�Ϙ�:>&4j�Q�i2�'9.4J�S�g�lx��@`D��[Ȭ�g�ۂh�B�)� � ����2��ݱ���*���j��t@��4��c��c�Օ}���$-S�2�: �FV�+���� N�OJ���OD�$�պ���?��O�h�c�)\�YfxT�z��xP#�q�����4K3�P%)�%Bџ�rwH�2zَ��G'�2{��dI���:�Tä��,VA��O�RR �oZS���M&�I�M��`"��w�p	cN�z6,�*M�O��m���M�B�+�ӱ8A��W���mx0����B�	�
)���*�d�ɣQ��0�jb�4�޴�?+OR��uk��Q�I��쯘OE P�t��*��鳠�Âd�R�'�`��'�;���ǩ(�"�"FΙt�����*T�����(�=+(��@W���?Ye�P;&�.@���4Y����
 m�h�l�
v�7+R�`pڴ-ސ���VN�n��A�	��M;пi��F�nJQ��ǰy��s���	�D�?E�����z�Y���Jb�S�o��xRds� �KI�D����Ea$f
�e!�OZ�D48��оi���'2��)LA$(�i!0�ݯ*���gձQ7�4�����|���,�4*��x%qW��3I4�y��V?1�Oq���թW�&�_����FK��ڄM��:�Hυ5l��ۄ3������\�S�k>�"p��,9��wO&W�)��!}ro��?ɒ�|���*ߨ!��`Fŗ 0���v���yb���`�P K�B0�b`�ůG�0<Ir�I2X���x����	�ޮ)��4�?9���?M��|N�uh��?���?ͻBRh҅�ķ5*�i��! ��-�C"�gԔ�3���>+찁)�*��OY�'�Rp�� W���b����)��I$<��q�mG�f:ly2��w���K?�mZ�b�8睆\�L
���5A|FY���ƒ^�2��M>���ӟ�>�O�q�Aآ�.�gぼ:M�T`"O����锻 �bb�׿jT@("��Ȼ��4�x�O���s��=�R�2I��zM �W�Qj�.����O���O<�d�ǺS���?�O2L�kFʛc�,-1�醬x���p��9F��E�R�)�H�u��g�џH�dү�8Pc��ϧ0[��EGj �j@4?��k�V060t,m��eN��ŀ7�I2�� ��E�o&J�Q#�Ǵs$����+�OֱnZ�M�����OT⟜���%@��E/_�Q
���2#�!�dƭ �\uhւR�0QP<!��n1O�n��Ė'i���-v�(���O�[eƝ�w�]�f��� =+Gd�O��$Έ9d��D�O��S@�*����D$;¾�b�%e
��Á�E/E^��2�*�9�p�Q�eҧ��O���U�a�fקC���`#EA�*$�1�E��-(�� �el "7��d	n��	��"��n�r�|2M��\x �d˚���Ct�V��yB������Ȋ�CO���t�0�Oޣ=ͧU�!�>F��*cJ�f�I���f�'L�0��q�6���O��'~�$��@� YsI�4|��1,E�z]&�R���?��%
+Î�ڴcF�w���p�o��>w��1���?��	�/��q�f+�+^U����̎A\�t�r@���Ճ.��J���(y��&�
 K��'�u:F�DC���{&"JLoZ(�O�����'�ڒO��B��j��T��+N|���"O
= �	X�N�r����7qlU��'?�#=IA;֐�B�!Ѷ,ڼ�Ӡ�R'C���'���''f0�W��:}"�'9r�yGO@�\�����u��h��E�n�<t�f�(2�6]�$�č`����T�	I�`�\�'.t��f�m���y��Fl}�Q{�K�Qb�`5,��]�8��FU:ĸOs���0̐�<)fY�'r��jƄE�:�4Y�ߴpb�'�<Y��S�g��+�����W�`ú����E�g��C�	�ir�49$@��n��HҨE\�L�Vޑ���I�I(���dnK�|25��*�G���C�&T�w�0��ן��	����\w�B�'��镀f3@=k��ơf�F�s$&�5j�4�XqO΁
�BN�p�P���9Ѣ-C��	�!�dBN�4r@B'K��������. �� [��NՐ�C���ΤaC�\�ɇ�q�.���Vi�J��*�n����<Qa�i��'cBTxB�jӮ���O ��cT�{!�5(�ֿeU:���Of��N�(v���O��LM �I��Z�u�y��ĀAD��Rg� B���E�SU�lH�� Z�'4޸($�x����+Z�ᒊ)���ɧL�T���hE	Y}�B��V���{�J��?�J>9�iO�V�vI��� +�����^�<Q�nY4J��]1⌛�P�$1�M�W<�U�i��TPb)Q,���	�"3+����|�#̥
%�7��O��|��i�?�U�K0��-c�������͎�?��b}��������g��m� 0Z� G7ߺ!�U+3}�$��O� �b'F�.Y��A��>�0`:ט>	�F����L>�
U��M�^�UK�F���oP��y�f�#���y��������0<���)� �풰�S-c*��H��03�pJᄝ�i�����I�i}�8�#��`��؟��i�e�N��4�V1����8IrQ�<���K�o�Zܘ1B��Y)�v`�|2N<a�+�-�k���^-�ob�(ic2`��M�x=(�/b���}�L<!�Ù4,����㇒0��8ZD \ ;=�� �<�7�Qǟ�>���Ol��4���A���(B�����9�C�	�
SB�A��٧E��=:!)ي���0t����O`剆n��4�����s�hm˥�ѥQ�yk��{(b��I������\w���'��Ў��ժ�E;��]�$l�?�V��U��1y���c�'�dq"%�^�4Iѳ@��S�R5����h�)Ґ�ئ�0>)VH8BH��@���  "�'��t�~�	=�M�g�i��X���	u��s�9�MBc1tu��_�&_ܩ��pul � ��Q�#iʸ��<������'��x"�m���I���9�,��O-Mq�b�u1����П���;}��<��ퟌ�'lB�-��C�P}<p�f�1�|�WA=-���񄖃CH�OD�x��K�0#B\ڪ>�Y ��'�ʌ(��n��'�d��R�2��qĝ9F!�J�'�T���I�Ф�fc�'U) 	�'#�7�!E��HA����Bׁ�!or1O
XP@��ᦑ�I����O���S�'��X�E犏>�*e����;��M���'N�-n_�T>�=?:���H]!~���qŊ�$�΀�O~AH��)��=;���5��<X�H�2��D�/�h�'������^ɧ�O�|Ṱ�5n{�:u$&}B ��'�r��U��v�r�a�o�i,����=Ñ���p��=6*��gGB�*�������M���?Q�P�v��?!���?�Ӽ��az.�gŏ�$B��c�4��'�<�ϓ0�6�yD�)j6
pSQ�(UR� �=�ęsx��B��З4#h:q�S�@���h����C���)�3���J<p�S�=�.�Q�ݢ`�!�dR�f,Z�0C���Pzs,��8Z����HO>Q�FH�d{���Cd��7�rM8DJ',�L��i�ٟ`��ӟ4��4�u��'�2�>�R2�<o[��Y��	!{z�;�e^�"7lx�Gc��6�F�3�1:�G~'��!�Y�A���lm3D�W�[*"!9�'�7|�RsN�>g��%�F�>�<�l�#�
_'sP!Yf�#E�I`�(��� ;��.H	��@M:���
gd�7)p��ȓl��MYgjj- \�(�:WS��<C� ���mZ��I� ��ؠ6�-x/B���nL����ɟ  ��������|��۟�'��kA3ˤ�9P!��z��cG�<O�����X�;��p@�i��gF�Q���(J��x��Q��?��xrj\9D�t�9� �? l�Y��+M�y��B {��0W�+��<�ծ��xr}Ӭ	"��	6��1	w�+5�,̉�"O��Hb��e��Mq�a�8.�J(�B"O���ښ]��Q��с0I���"O�  ���8J�¥Xv��}�B��"O��#Ն ���ȑ�A$D���c"O~(e�݂`9d���i�)�v H�"O���W��|���JCK}���!�DǱ'�44	��{��SA&Tx�!�DXL&FҒE�^�>Xx��B"�!�J�p��C�zE����#�!��V����B��0^Q��m�wz!��W8X�^(h���:'{n��g�ɣg!�$�,�X���G%��CU�ׄF_!�0L*D�#��B�0�!�^�L=��Y	V��P�B@!�$E'b ���0D�t�F�B�d]~0!�d>AK��"l�<�{�C��n!!�O�Re�d�۰��%ya�H�:=!�Ӣ:'���K���c�a�4!�$,Y�L�ZƦĦ9������y)!��!n�i1�	�.�����3�!��E5P�����)F�rUp��UL�!�$Ьt,�� �T&A�F����)e�!�d�>X}R���L�Є���ǋ{�!�� x���FƲ�x�B!���jsaS�"O����-EdP}xѨD$2n^4�&"O�\r���[�ݐ�) _���2"Ox��1�U�K$.y��yJ 5ٱ"O����4fѴd�D/-�HPq�"O`)c�&P������&`,���O��x�=�)ڧi��$���Z�MH2�넀�`�|��5C�Ik��A&�!�72¬�O\�c�B#lOV2���38�\�:���)�(bV�ɛ�MS������4D��p`��C\���c`ԖQ��mHQ�ӪO�V�9�-��|��^2�lJU��Jx�@K#�z�H��&v�,S��>��P��4�)�hɸz���SÀ_��tb$�F=J�)z���4�a�C[���=I��i�t7-8u���"�˕:-��[VjFp$�|����	8L���� �i�i�� ͒�Z�!��C����D��!�a3�@"Q �ɁNED�'�Ш�ԁJ�K���blӈE�0���I�Ţ�!����	'ۦq}&�Iy~F�c�Mh2�H�r�:�a�Ǉ����������p���J͆��L0�,�P�&Q)*�mڥ���'aɧ��B*'���� ̫@���
U���p6�\�M{@0u#�����Y�E�ģ\'Cv�ɩ��4#D�͂��JT}�E>�?�Ɂ���ëM�h��V���8T�ݢr�_�U�<���	567���f�/6@��fȧ ��8�0n�k�F~r�|�>A��;�,�ض�K�a�����Y<[<��s2)W
Cl~�b�� �?Xċ��V6'ql����ل��'#D��
�Xri�ås#�}����ēgF=�o��w#P@ �
[M��a&�@����3p�ݨ-�a�(I�d
�:�.=��˭QR��曲԰<!U��(l�@4�+u@���@��65���"T`� �P�X�J�ay��R N"N��Ф�6��	�4��(�,B�Ɉl�:`�P�ߠgj�����Vj���:$z�0'��#���$�W��ZqS����O�&X2薳�0=Q���(�,	p��$<���%���~��Wbʿ	bs-�d�AD�]�2��,v�d����N�i&�'� ��oC2�m��B�K�Ld3�e �Ʌr��6m 6%aZ�D�e�D�?�V!�`��u��,��J�4���q�eU0B���Ys�ނ+)D D~�w�∘a��7?zR؂�D�#�H��O��ӗ�4GR���I
z��X����R��P3��V�~������E��*� 3���_:�M�� �:g�Bԁ@�A~4��F��f؞<J��&_(ذ��51�������#z�)gT*�q��O��^ Rz�[�X���$ֲSV�A�WmK�uf�I�r��%3���
`��܀!6�k!N�m�֘k")�5w�'��ҥ�^�f�I����AB��ͯ�M��/�|�n���3�D�Pp.�X�H�mP�2Ua�J�@�����9�����F|B�eމ	)ĞS�N���aW�UFp�$�<9q�η=��L��Rbrl��J^����=��X#��������k���nT�-:�=�DFDx�@`i���+o8�ж�ߧ\�����ɑCZ�6-G
#��l �m�4#	BD�����P`2J�D� �>��c�O�f � `�$+c�	CF���@�I� )�F�ke��kz���`�~Y*e���)�I��y���YV�:e�Ѭg|�7�ZghB��2t�T�B������K��1��@i��@������O(��T���j�1��DϦq�� � �R� ��%�ը��.|�	$QZ��&���t�oØ� O:�BG��[�뚩[j�r��]�07H��<�%�,n9שFz���h�j&@�L�����DM߫&)6` ��ԑ[���BM��؟`18T��o�t�k�f˸*�PC������÷fؾI�O�Ts��&+Rt�D&�*g���Sv�@�>��$UNl2���{�Z6��k�t�F"�
'��Q��~Kl!i�jE�4X�Aeȩr�!Kt�Tg��xbA�a'�ڂ$��霐Y씤~kx����	�x�@ e�G*Z�P�鳾i^�0 rFL(��JAc��M�5ϓ#f�n�+�{r��4" , SF�@#�p�����Y FI�	�f����B�%@���#����4(ɪ	�X�9��Պ!�U�L�R(����i7:���D�;�N�9��/tv��V���J�T��E�D�{`�PE�i���s�H���>i�dR¥�s�ֈ �K�q������)Es�N�4H�8�1�i�}� в��8�$�Φ)D�OT�	��M�`�Ol�02čERB�(v�n �"Kڧ"UUs��GQ�'dT�1q�R>ojc�$����Ү�;��tc�,R#�๲�O^�͓�?�i����֦�Z�ua�$B:��DP����jCG!������� i9F\�v��ƱiP� %��r��^�y��D�[5�ࠄ$z�p�a��%��|�Q�!N�8�C��7a�6�Z&�'h��1Sf�!.�ޡsn�G�4r��\?s���'���I�����<E�,W��0u�V]�g�ա2��Q��'p�8P�p�7�B���� ��TZ8�x�o��(%	��'�t=�3�-�y'��7@�@�SW��e�b%�C�߻�HO�<������C�d����Ӻ�wKN(tfPA��G�$
��p�Oa�EatH:� ��B�1'��M��$�{�� >b`��2��#��Վ+pKq�i�L��U� �!$�".��|��u�i�Z���|��H���bG)R�?KJ���Z�Jp��nl(dwoX+�@	Q�|8�� �>%D��W������P��A�'�>���?��R"���'F��(�V1�rf&���Z���>J'�H��)W F�z���)y�p���	�:phGl�fJ��9���,(,�"Ö1Q���f6M���*P��M�3Z$E�&E��)�4W��	�FЮ��%��D��t"��L).�����,�#B�<Q���!@��`'�H;8����wDQ��Ms�����ޕ?y�6-U�G� h��q���>�o��0ZAq���p2���o���3I[8F-Z�p0���//��	4W���~R����0i���6Yv���"�:5y�BU�44s
L�a�.or\���	=�F8i窒�B�\|P7��%<�r��M>Q+O�O��,"�	γ��dkDo6d�W"�8�q8�ϋ&B6F��
�1�d�tB�7l��G�D��pJ���9p�-��b��=���#�S��gɶVs<��+F�u��NE4-.I���Z5^�3�}B�F�Wp�ya��U�е� �V����'���)t�$�^8Q�cZ
DT�&��ΓN������6t�u� ��g*tM�OT�z)Ŏ3���h��R3�fJ�7R�nڼ]m��EbV�:CL�sqɧ��)m�t,HaMx14r���9b��Bע����QG�L���ֹ&�rdѰF� 5p�T��n(�l�irW���O��kv��٦i��@	Q���e��j<�ir�����=�Q������1G��C��K"4��FO��m	�!��8O�%@�����-�� ��@_tM������0dy4�Z�3�~i����M;8lk!��'H��`��`^�d�ʓ^O�e�$'��'W\�0�i�Q�B���O���-OLxx'�y9�<�����HR���A�Bd�b�ˀʋ�]b81�B�X�,eC&�L(��!�S0C�.#<���`JEb«/5�@�jI0=kJc`r�HMz�XțDߺ����!%�L�p�m�}�j�hIOb1�ap��.���<�{��M���a>��q-ݿM���"��|�&�x�M�YW����	&iyLJ�d����ñ!H�?����q�E�::�AJ�W�'�@���kS���.;�	�bN��Y1��>|��"- ,�'�	�@0t!I��38�VM���$!6��'��ܛm�){�$���MiȄI��ܝQ�̒��x��>Q�`4;(6�#^�8I�D�j�bP���O�a2�A��tpN��"&5�h,��&	���V5��)�>���C�<F*�a'�EY��0WJ�y��&���2SBř,����o�;���"��^�I���Z�����m����>!�M
n���2Q�D����Z�\�� G�(ip*$�5�H�)�<P��<m#����l�$�y���.@�]R�+ZN�nxɓ���'�~Y���>-�J#>�`�1j`��f��>�L���I�tc�Or�q$͸YF��C7Ȋ�0��1$��<��:I(�:q�t0�)eH�eF�L����S��T��"~%�`�ĸ>����4Xجk� �(n�����:�
	H��ݚf������O��?ɷ#�~ZA-��|��t�uO�hق����T�(Q�Y#�ѿi��"?���Ѷ[��q����D�0�D��Ц5؊�$�z��GvP ��O*$���ڸPHi�`A:5I	7�R"H����Ei�i: -�ȼ[�nʞ���Yg���2݊����<�L�d��ѕ+1O\�6���٢l<��1&�t�J(W�"�I�RJ��o��Qpl����J��Ov���I֥>�l�C6&M t��	q'aG�N�ȸЯ��1Hƥ�&����źv|��KM-y�e!�f�W�\��d�W�A8�Ր�A6R�VG|�a��qaV'���D� ��]i�M+?w�
,�p����6t���t[�%�9FH����-V<*Ĕ���FG��hO�q�`6O�e�����C�6^�,j���'	�ѺbmW�]>�i�M=O�%JC㚕=v@�;[�:���� �@�� ����$	Γi9@�4;O���ʴD�@�gyb�G�S$�|؂!��`�k�j:}e|�Z�}�FO9:�j��iq����Ms�I�O۞Ir�B� ��JaC{z8���G��D��T�4!����s}"H ��Lqq�eҹ\yNP`0B�=
.����7W�&��)O(�ğ>�w��Q��6��r��;l�j�iQ}�6-�/@p���O��򨀐)9�}���|Fy�m�M2�H��	֭p��&���XFO�8PE��9�n�Y��P� �Fغק���D�u�̀>Kę�օ�5���B �'��-c
J7���Q�w�Y���Q���B��	�O�t払]@���d��!��O�Woݍ�"��8�U�M� L����R���Y�m�]�����}�LG3�1#�'�J���n]�=O���~�Ȱ�K1 �Lqy%
/R�������M+��	�M�ƃ�R?��5���|�I,Y���}�R)ˁAԔOٰBTl�֦���K
%�0��N<���}̓�X� ��M/@Oʄ;����(�e����)�M��Y�0'���/,O��"���$p <R悲U~�T�G�䒒��U�C�i�����c���3o[V;���ѭ�%Q�R�j���@�����΂�2�n��Zc��<2s�^�)��Y�
��JE��6��sG����'�Ey��ʜ�ħ�<U(6�?�	���.?f$%{�����K�c��O�lт�}A���Ϝ�$�б�'�>��.V�*��H�1؃G�L��c�ʼkbԩք�ZC�<z�4U��]���I�i�<g���C˨d��ۄ�HYZ��u�1l���H�e��H܀��O1����S�? 	r�rd�HFE*�&�{�J��`'�a"C.@�$Ԅ���c�[X��r�k�
I��iԩR�T��$+��MS#��&�?锢�� d$�;��)�:�T&��?�x��獹G8�"ӓ6��q���̣ckLW1OUȍ�ǈZ�1,�a�h��bJ���P�̘>��'E�M٫����[h�O+xC�[1An
(�wj�#��s�}B�#>f���EY,E�+�l߉��	}X�a��)b9.����)5�8Ӈ�ϡ�M;A�im�|`cB]�q��'�a��8=�vjV�M�	�N�i��;v~����O��֧�O��P���z ���A�D��s"S�n�C��K1H�Vl�t�Ǐ�H(�m�[�@H<��G��Ey��$I�������,�`�L7�y�5)���Xq���"zE!Ћ3�yb��b����2w���ʆ,��y"�����%
97D\l�U��yr��E���hF�"14�܈UM��yr�Z�:3����`�M�l�-^�ybB��=�2�k�J_8�!b�U��y�A (��c͂/�~lY�"��y�f��j����(�"%FUF����y�Ҿnz�]�HK�U�Mc���y�׬w�v%&�ߔ ��k��ycՊ-3Q�KRz6��/-�yBo�"�K��Sg��i���yR��\;����E+WH��;$����y�������ۧ咬#o2���B�0�yB �$�Ԣ�5�hUsJV'�y��݇	�v��R�M�J5�r �;�y��α)O�PÔ�M�|M�1�R���y�cV
Y�P�#��!e�A�q-F��y�eA�'���'L��M��%K��yA�Z�(!c@�˹���ڥ�қ�y��UWy#�Ϝ����(�7�y!ѽF�|=B�D�?���f�'�y2(��"�tYk%+U�/5�u5�y�j!l��J@�Y�j�����F��y��"6���(gɴ|���R��y���4I�pѰ���X�$U�A���y��ɳp7��Q�	5@X�BX8�y�#�{1�u;e�܏{ْ`��bC$�y�N^�Jx�R6
�JA���'�y�^�w��@!Ǭ�)4��k���y��,+���ƈVL����
�y�����Q�`
�z������yr.^�	+��@F��u�r�z2���y2�đP���g�΁rAh���隝�y�NA r��� ry��Lp�j���yR�¢)���RU(�0y��
�yR��?1B,�v�>|J���"N,�yB���w���:���<�vŋT)�y��C:2HD�1�̯��x����y҅E�^�
1�v�C�
���ӏ��yApd���ꦸ�˖;�y���J����2%G��L�d�θ�y���*ﬠ������2�d����y�ϒh�5��lN9Ψ�ȓ�H�y��T��9z��'b9����y"S�5V,������m�A˛�y¯I��A�$�0r� IJ3����ybbE� �`ApH�a�Hc!)�yR�ʈ~�pLҥ#�	Z��=y����y�$Ũ�����,��C�02��ў�y�G��$3l�H7#J$"�2�D]��yX�g9�(�tሰ�,���]��yB��w�DP*9m,��A���y�oG )p�����4)��-ܢ�y
� �<���ےk^���2 O`�D���"O2,a�n��F�"/��Q��b�"O&�����v�(�f���Up�"O|���,U2W�V���'�*�x5�C"O4ٳ���1�@$Y7��^8��"O�a"����4�#ԥ��6��=Hp"O��g"GS�Xq2%B��:�Ұ"�"O�AS5G��;V�9:����1"O`١m�U� E�# ��@T�""OB��A��=U��8�!<8|���"Op3p#B&3�> *�)X�0�a5"O&��-ږ�p�c.��)
�"O�u�F�\�1m�p�bź*S|rE"O�d�� *��P���1oN~MI�"O�y�FP<������i>v��D"O�$5� T�Dx��݀t<r�"O6ɠ� ��gt�z�τy.�}�F"O��K%���_Ͷ���ķH(T1Q�"O�0q0��vH��)�'\6�)�"O��(��]A�����D����"O0q&�ٺ�dL+%B���b@3�"O�MY��ȶ~/���&��&[�r�Z"O�\3�e=���۔iؙ }f��t"O�pQ��՚t,~��h�j�!�"Oy� �LI�!Bç�S,\Qu�'X�R�-@ZT�D�+���?[_f���'��"��.$\�9B���Y������$;�!��l˘r�F��rb�Aю�ȓ#�BdY��R"8��l	6mQ=�zt�ȓ7D��@��:x�(����&�|��F>D�B��vb:����üR`>��ȓ_����--� �j��igd��IG~R����T���΂un� �]��y�뚪x6�a�`�t9P��P��HOj�=�O!���a-	�yy�I(g�!SaPm+�'t��z��B2R��a�� �DՄ�'�,��3�		n�	�uʀ�h�.Ŋ�'9��%��1t�̄�uϙ4]�6A�'j��ƭՠ~�ѣ����h��'��1I�I<Qʘ���7�L���'
H z�'��{��1�JӮb20��'�Nh
gEJ�y5�!X����'�&�Y#m�vs���e��>��d�
�'Irh�G ��= ��' &t�
�'��y��@O�o�ؽ�pI��yt��'����� 0�:0I0+�#.��0��'ג��u��C�F5���ė i�1I�'��)�̍lm�J�jN>���J>	���)Y�+g���pN8��1��5F�	Gx�t�c�ٚ{�|�	��6�� T%9D���(y���
]����6D�x�2�V)o��� |��ٚ�I�}��W�V%h�&Rut$�`v��GW -�ȓ�p��`�*4mz�*'�Y�Z�`�ȓ~��䫅䛬$�L=*6�NV3�(��}���XRLX���`@Ti��P}��/ntk��ߴ}Ql���
�(�tU͓��'*�?q�t���4�2�O�?����=D�����W�B$cb��1.�K�N7D�hQ,L�|�.�rf �K�D"0�4D�<:��Y!-̠Lcp��P^h	c�4�Dr����xT���������W7C"C�	U��a�煚)~�^����S0\�JC�I ~��<b`
6~�pY�eCR�kitC�)� TI��q� h�� �ptm�#"O���,�_m��if
R4D	ve(�"O���Ms��� �*n��d�"O�X�0�΋fv(�K���d���
"O Yв I�Y�e*q����`�"O�4��o߿��EkЎ �z	!�"O
����������o�U�2���Y��G{��)�ù9�M�`�Q�v)P7$�!�DO!Y�Hey�!T<hkG(��qj��4�戟8[S��|�\h�q�L�TppL��"Or�24��&<�%�G��d���;O��x����w,Y�%,*�#e#-*ʐH �� D���IB7zx�͡��Fb��XsO!?I`�*�O����`��lH�@&b��,�u�'=��D�4bP κ����`D�����Z�hS�Ά>��r����^�L��ȓBEtu3��ƫ|��Q�\t4F|��S5��İD�ڸ%�~]��"�TO��=�~��j��0�(N��r�Z^�<QV�T�ݲ1s5�Y�?�p�r��<�5
q�>-j�M]�v���9��}}�)ҧ1�M$���K|`@5�D$&��Մ�'�����ch��*���b�>8���Ol�\J6�m���M�
@ިB��#D��Cq��it�99 ��&���cF�!D� �&φ:W2L0�͍�;�(��U�=D�<�%Gѩ����̜O����G'D��2 Q�o��]�%��_��CT�/�L���O�00Ó
��C��h�N�z���������5H���`�@I�0x��ӮĈ+m!�F�"$��ap Rw'(0��كgP!�DOQ�8�V�C		$�љgcҊ;�!�_�l)d�ɔ�v�8�{�O��a{���N��X��5�J.�*X���ٱO��D��Q��h�k�p��RLƵ]�!�č�S,T����>����!aW�"��}�<A���F�����uG�tCt�:}��)��3ql5��ʝZ�X!���	 42�C��^.���O�?8�h}��h�%~C�I%|�z��M�&�8����i=PUZ��-�S��?��n�7z�0�c�#^i�}��g�<��$E<�x��C�k7
9���_�<�t	Ҕy��Ʌ��:nvDK�m�Z�<�cM��.U`r�ߗ>4Pؒ`�}�'g�'�O�=���V9��pH�b�6���O�|{��Z�dɬX���#{H�y��*��*�S�'^T�]����0Kε�w�7�\%��Fz���#�!'�ʌO����b�$�!��8v�-xV͐Tļ�b�:E�qOԢ=%?ys����f��|8���?D��y�cY)$��[��A�9V�X�"D���1+�ZR�¨ �x��C�%D��&�H����v�]�d@Ԉ7ci�	�\��Q���J�A& �kbǚl����	`�=+TYx5��+�{!���o�^,��8��e��w�p�B�I�('ح�'��~"�J�F�`�e,S�dt%p� ���y�Ҡ=̆���ŋ�X���q����yr%����&X� xW#O�yb�I-4�Fa�噚H1�s厊��yRK
�*��c��?sQ*}˵�0�y��Q�rÖDڶ��x1���ҧ�yb"I�3
���MDpXn��F'�y���,w<�JDoEל� ����y
� �Uӕ-O�,	�6�JM��1#�j���	D�*���,Orj��� q!��:=������u<x8�4����hO�|�@��	&Tx�'��!\���'���Ey���ܵV<����oZ3|��@I�g�:7m-��r��\B!���A���PCJ�;0)1D�8�G#�o!�`��b�8i�r�h10D�������2�q�tJ7]�n�@�1D�� C\��>��J-x�0��
$D�tj����0��CL�#
���d!D��0cCJ�s\���%�,�T-�>D�,�g��3�V��D�&Y�n�0$?D�\i�ʎ�5��H�v�I�Lۂ�XP�8D���4c�!�&YzGO܄acV	2D�8�'a��
�@����]�t6�"D�,�A#�1wrl��b��m�,�� e D�8��MXzV�帒�58���D?D�H�u�l8����i�CB�u��*;D���Sh�Se������ s�-���3D��e�B9"��@!@b.<Ⱝ@�.D��q�雋|��x[�(�LԤ��*,D�x��� �u��h �wHČvF(D��K��Tlhu�W쒥)���ń;D�� O����Æ-~�l��i:D�Ģ@�I�C�`"MЃ^�v@�DK,D��KPMʉ1"�i �?���->D�dٗ̩MhbѺ�#H ��5�<D�h�!��i�R��v��'Þt�4�:D���C��K4�����]�P�*��8D�`AB$��ʎ���P9~�W�6D�p�g/�+}x�9���K���� �5D�XX���!�<���������'D�d�&(W"pq�H�������a��:D� ���Nw`��F�@6]@�L+D�pQ��N,R��1�@�GE��8A$%D�\���C�4�NQ��Z:�lӑ�#D�ܣ��Wi�,
1�Y�9�l4r�;D���t�P]0i�q�K�v�~�.4D��ə�UXD��(��E�\hi��2D��[EI	93��(
��m.�IP�0D�8H�GT�[����p�
.c?��h��)D�({��{~8����1wn�Za�:D�dK��'��l)U�wqU 8D���l�>�}9�n�5M�ɶ�6D�pC��Z0Q�X��d�Y<q�f����5D����)P��=X��قBCZ����3D�l�U�
w�&���)܌x�f�0D���so��^T�H6c����H�,D�8 7J��?Ѐ a��5 U�y���)D�0(�"HA�D"�P�.@��3D��q&D��*$:d
/*�S �.D��:�d�a��pA���t��ڗ�.D���C+_�z]���Ǒ��Y�R�8D� jr��Yx:CwD�?a}���3�7D�P!gBߟb�P���	 KCd9gk9D�P�����q��kڣK�@���%D� !FQ�| ��dU�Ui{!�$D���&��N@&��r'A1#��p�'D�p{�m�5=^š7��t�x�8�	%D��K4��?�q!G��+yYB�qs�#D�lH�%:G�,ϛ�rZѳ)!D��O���b$Y�X;T��CE>D��ɵ�S�B�|4b�cB�p�:�i��8D�@�v��=��|[�	�_i.�Ň,D�� ��;ƀ�%pr��`͓.����"Of�Q(�,~
�����L��#"O�P���-:fi��D�}-Z��&"O���PEDj��v��B*��� "Ot���!KI���J�Դ:�1��"Ou��	/Q�(6.�8+H��"Oh��Q#Sg�8�Y�"	�o#<�R�"O4ls�n��g��t�u *�<� �"O�� ����4�ʯ��i9C"O��h��H�6���'˼����r"O �à�91��Q3���Wg@0rV"O*!��"X�>�2�%����,´"O�ܺB$
#,����#�cEh�x"O�]�2 ��=����,ߕp��"O(1 �X�H;�ϐ[;����"O��"GÙ3`H�� 
�0 �y�"O�eA3�ݖ~J����$)ϴ�"O~,�$�Iǚ��A��\�"�a"O��H���RM�%�$��;@��99p"Oj=Jg�}j*����N����"O�%�%�سd� �$΅L��L)C"O0Ѷb߸"�T��M��0�S"O0S�mC}Ҧ��R�y�anY�!��z��t�BkS�Jo�-k`h��`!�D��41:D�3↨GU���6(J*�!�� ���)���O�L+ӧ?�!��\�D^��h�ʂF�i���7�!��!E&P�K�����3k\�[!�DM�A�8���nݶ��-��J�"O��;�*�gz�Q��
)y"E�4"O� S�d )n���#�Nh(D#"O�qT���b!�%�^3\H�"O̭ʆ �>A0ƇN0��k�"O��r��$7�ցZr�	@#���"O�7͛w�f�3v��pALA�,3D�$���$@��T�@(C�<���+D�0j�lR��.��s��D:h��&D���EX�.	�g��&o�Bi��	#D�X������]93��	Pu��C?D��"W�W�S;�A���	5�}�P�;D���.��JhR���?O|I�3$D�� ���R�j����F�ر( D��QRU_��J�j�XDn���L=D�4��(3VvAHs*C<*���(��'D�����\!�(p�oD)��i3� D��Q�)�dJ�*0Dչ*r�p9p.=D�$�ဩ%V�˦N��t���6D�|q�'�&_�T�7[�����4D�xzVN�7�fu
5�ՑH����B�0D�xHAo�&ʆ��`��z�<��3d*D�����"/.(���Z�P�[4>D���1d֋@d ���WI�^xᡩ>D��C"N!��ж��hS�s6�<D���A�0\�)!KY/$<{�n5D�l1��j��!�`�L����9q
4D�H�
7T�Th��̙{A4�вO2D� �wC �yR���8
���m.D���d܄=dȵ�D�W��q��+D��ȇ�� �Xj�&�.���!��$D��4��J�����j�����4�!D�˳�P�bb��U��.�|�*1@3D��ؓ��=*�á�?/���D�;D�Ԣ`�Im�@@HLؕ`�C6D������O�a�s+��}���2D�� �@�&U�p�%٠R�
���v"O�����V0�Ȣe�
�V�L�"O��S+�l	���F;Y`�@��"O�ۢ�����d���V&6-B�S"OV����.ns �w
��j pܰ�"O�;�� ��akW�^! 6��Җ"O0���:��dS2FY�d�S�"ONx�A/J�:�~�A�∉_6h$"O�Ut)�U����Y�(0�"O����h̲6  3�a��"@Ҭ�t"O�!��H	.�Tg�%׺XӴ"O�%X�KO�Q+�<���˺'@�"O�a�'+�KXHX1A�M1���"O`SCۢ:�&���E��Z
q"O����)ѝ$�ܠ*'K��wtȈB�"O6�PS��@[�XC",9`�I4`�!��˹S:�Ha��R�c�T�3�!�d���
i ��N�Ʃ�'��2�!�Dҧ@V��*B}z y�Ã\�I!�db[��1��БFmv��2��;R7!��Z�l��0iQ�pE�%����-:!���>1 ��a"	�=�I�0Xx!��2i@}���;!�<y�E�``!򄚡36XQfկ.�2`���nY!��0N^fq�% "F�@�j`m�T!�$��i���$�Ջ0n,��̉�Q!�$�5]Z�R� �0]�
1��5A@!��'�$��H�i���w@ӲR!�د,Ɖ�P)P?W��41���#s!�D�wTF(�R(%W�=��n_�ld!�D���m�K 
������� 6!��B"``�	�6�R���UP��ߵq!��
 ��\���D��,x���P�)!�DH�V[�d��+�8~5Up��D�!�D4��q�O�:'�p5˒�Tz!��R�h^E#R A��u�C��2�!��K�=����N\c�
Bf!�ĉ�<ݺ��P�ذ6��-`!�׷(�첰c�	J��Q"F�K7`!��;U\���IH�5�`���a�b�!�D�".m�M+A��HqĠ�AG�j�!��\�5?�3#��'Tz��LU�a!򄈢�r��[��t%��eQ!�$�8"T��B�&F�>p)tF�6;!��+P�ԉ҈Ƭk9MC�*��v2!�$��Vb9Rb�+ �c�ǉ�|!�σb�$�թ��,���f�ר"!�-h��,R
�Z������!�Y T1�̹1���5����FbT�s�!�غ~F�(� �jG愫ѣ��!�D�,Vf
ѻd�����H�9n�!�d@�Bǎ��U-@��̞c�!�Ҩm�l���"�U7�T��T*�!�D_�������F�X]�nʟ\�!�DHQ�Ι���(b�*�+�l�%J]!�$�@d.BF�P�U�@L#fl��!�P�:Y�x�$���~7ʁ�ᡔ.:�!�D��
�phf�/*����!��Ƶd���	���.*,L�F�U6�!���7�]���A%`��B f�:O�!�d k=�x! j��	j��O�6�!�D�� .
h�.�	pU꠨G���9*!��:Bz ��@���c=�Ei3jF5!򤜟|$c��Q$i�*=�2�đ !�� L03��
����D�]�b�>��"O�j�$N��� ��x�n�I�"O��=�}k�I�k����E"O<����Y-a�A�2n�Ap�̊�"O�Sw
�)E����۽UÆ\�"O���0M�>nJQ�ǟ}�bEp�"O�s5��- e�֎�)�����"OZ�S�j� ���@�n��s��8��"O���q�[(8䜌��❔����"O��P��(j��[� U?u��y&"OA���!�: h/J"6lH	�B"O
�Cq��`��1L��lBġ�"Od���G�Im���ƈ�y�ʨ�"O.d�0�Z��Ԁ�`�M�l<)�"O�	�ѡſR*�y��Ão`�"O�@��`U ��Q��̂(����"O���e�O7~O��qc]*�Ac"OB�r"�ٿH>:���^,Y���
�"O��"bz�T��
~��<�Q"O�%
�L��N�t�Xc\
zɶ
�"O��e��;�B9qa��4���,�y�KI#�0Q��>kh��ٍ�y"�xS��qG�+Ři�p��8�!�Ȳx@��3�/�j��2NK5�!���&b���" dP���zG���X�!�d�}����qL��]�fu�"�Ca!��
�xi6��2BL�p�x1��F��yD!�7%!Bᱲȅ�&�8�;5�(;!�е9H)���H8w�����)�:O3!�$S�ewHe1)�%=l��cH�:!��=��Բ����SXH���	2E
!�$�<ΐ�bs��IL@A�Cu�!���]���� �.Pq��1X!�$
Z; �96-�.,|��c�73!�R�eϐ<"�ëg�4l�*!��Œ"r��D+H*! �����ɓet!� -�l[��O;
�Ғ+�\!��!���;g���S��d�S�S!�P�Z�J�Y�Q�7Vк�*Ì"/!�DQ��|kePvu�U��L!��0H��8
�����p��(
!�ČL�h�Q��TRH�j�&p!�QyNlK���Td8P7
X4C#!�C��0)�슪r>��e) {!��M�uiH�PB�Ҏ.Ƙ4�t $:!�$H��"I{fBF�$
.(�W��+y�!�dLY�u�n�7�̔�e�hZ!�d_�d��maă
 �Tě����!��(������th ga�17�!�0z~���c�T�)�����9K!�d֭c��;D�F���MC�T!���-��q�
v����L!�!�L�<?�2��ԭD�-yR��=a�!�$� V���c3��<��Z��V=_!�$���҃�I�s�J�02*W�	�!��3�=�A/��-H
��HL>X!���h1��bd̅��%G�~!�۶l�% gO�/:.N�椗^!�D_P>��r��O~��26��:�!�5}���@�ϵ8�����W��!�dM�W9�$ß8�EҢ���!�$��c� ��T><�~�X�,\�!��8���Ub&m�hAE!�+L!��d��<��K�2u����.G4;!�� �\�ꅆ}��]�#!�mt��"O�1��S�(���:"AD2BH�St"O�1p�
J?XkbX�'@��}�"5�4"O��jd��,�
 ���Ua�=��"Oε�B��\E$t(�NY�q%�pj�"O�����3�>�Ra��o,��It"O ��-O n�1�j�&
?���"O(��ujAJ]��Ѯ>�"O��"f֜4\sbH�G3�h��"O�����6�Pl�h�	F1�9F"O&M��C�\@�	��1��0"Om�� ��� ��"�8�ld+�"O�����,�0� ��s�p�8"O*�YWM �X���
A���i�<�!"OV�!G�.O)��ÂW8t�:W"OF�3`	җu�0iz�c��o��a�"Ob����#;Ix�"�ݯc$֘Y%"O2x7�N�	�\���#z49�"O�e��+џ6g��c6,}[̌�"Ot�XR�J��
��j�%V��i�"O�"�
ѼvfF�*;*P>��"O�x�q�	�=ؚE�1��	<�+�"O���A��i�����l2Ƈ
4�y�
�^���5I��*3��A����y2΋�.���2�_$%�Hae"Q%�y�
L0~��a %Pr�) �²�y�K�-	�D�3a�*.��`@�۫�y��O�( �p�1�����F�y��=vp&В���,,�p��Kˋ�y�1g	��XqNJ-'��G@��y�ރ)V�0���/9,�:5fV0�y�MD4| ��d�C� zJظ�h��y�-�I ��R�˦'f��ڄ��y�(ǵ{a �J���:k�������y�$�3C�:@SE�>a� �S�L�yrI($\}�%U�R[��̕��y)��VȽ	s`K�3T4�#�*�yR�%le�F.&?x�R��«�y�&��0*X� )Wq��� 	��yj��h�}#��82y�Ma�� �yBd��fl{pB��-���1��G1�y�C˺��WH��p`��k�/К�Py2%�=(���z�D74�x����y�<�"A!�6�zGĵ'��a��L�<�V�e�`jd��8/C~�^d��&n�X��C��-�L!i���n� �����@�ۿo���lT�ԇ�i�X���	s�v-a��!B��ȓDhx �Q�~8�㥋�x#���T<9R� ���.G8�RF�U�<Q"�ֈE1:ـ���1gV���g��l�<A�n�b+ΰ���"��,)�*�l�<�� �3k�D<���Fr��(oe�<���
 ��`q���,�@�W�]�<y$�	�G��LJ�
�2J+ `^�<�O���Л'K���i�Clf�<I3`��j���E20���:���e�<Y�'԰p� �T�\�i*�"b&�e�<aD�4LT��6�	:{�ڝ�0�l�<1�*9/�x���4{��貍Se�<qp ��j"X5´�Ǖw����-e�<�@B�O9z1��-�y�+_d�<Q�(E�p���#�&<������MW�<y#�=0V�QG��!��p���IV�<� y5
�xrv��1�Z�h]z"O�����7zJtb&�D�R�~�"ON(�T�]�7иCՇ85����"Ox ��Ľ7����Aǜ0F0��W"O�=A�Ɗ~�X	 �%�:@�8F*O�T`���Q�N��#�8̂Y�
�'ڔiG��K@��K!ϯc:i�
�'��SŖ~�b�x����c�z9�'��*!��	S�<A 2UO���'{(�S��չw�d�P�I#.�8�'��:��(a,%� ��I����'��X� �Cq�����H�oÐ��
�'\�ي�/�X':aL�m>�i��'P�Gn�.C�T\K�aé6�%8�'�^|�U�WK�`�YѪǵ&�����'>�U%��ba�J��N	H���'�2mK���#W`F�P�� P���'Xj5q�:Y���ÀZ�qM҄P�'8�a���ʃP�<��E�y��:�'�Μ{� �/��8�@C�w:��'���p�eO,o�Tj#Î�q�<�'w����m�T�"bb��1
�'�ř��\+J��X�AN A>Q�'���c��E�45���r�"�;�'�>5��f��P�>��,÷j*"�"�'7�Pr�g�;,Ϛ� �f�����'���2���?E.��,WV1Lؠ�'�\aE��f��)eL
<B��H�'?�!��E^�qdBH��1�'N@M��E��!�4LO���b	�'�R�	$��c&ذv�Үa�����'*M s!�$�]�T��3]�xݒ�'B����}��� J.|X�<D�P3�K�5��1�P�Y�i�����$D�PPMG?Q��
�6D�r`"D�,�GA:W&4i���[�+�.�� D�X�D%�����Z���! D�03�՝#GJ��s�R q���p��#D�S�Y6<$����b��LIE�6D���d$7��ē1�J�δj�5D���d �+J��!F1Zc�ѩGG1D���BC�.oLءqiB0�D�0�/D�4h�H��"����+�6���a�:D��ՀI=�޼Z�a �AI�1�$B2D�����`�jUpv���I�C;D�<�֟t�v��v�bO�i��3D���#�M�.e��-ff�u�R�2D�L����$`���w�ټ
fXi.D�|#a-2�i���'y�P�;� +D�r3��\�染M.0�۱�)D��uV^��1z�ˈ5Mp�P��3D�D��.h�1��:P#�����/D��÷�W�6
d��RJP���*D���휵rK� +�m��S4���'D�tA��#	^h<�W핈4R8l@��;D��FɆ ꢙ�$+I�b]ބ�C&D��*�.ʄ=,�GG�)o�@Z�$D���#C�G<��0���Bl@�`��!D��:���65n�y�O�+e@����9D�����t�B��KB w<�!1��;D�h�`���lhã�*B��m�D�6D�Dy��L@��)�`c�'�Xxc!.9D���5W7:�2�04�ϟJ�$:5 "D���g�܀>�\�UIϮc��8�S�2D�� 81@#�o��q�#FaL�tj�"O>����NDP��T [*p��a��"O�y�f �����_(E�@�"O�0A�`�26��2R�oY7"O�,��#��M9�G�)_:�2C�8D����G{2�Uc���1�<Az*D��cl�*)x�����z�B�&,D��8��)h��3��I��G�*D�ī��P<%�@$��@Sx�� �$'D���	y�4�a�c������%D�(�c*�B��`g	U�Ps֙���$D��@U)�/�ƭaB�M�p�0F�"D�t�O��*�}�n�4�t��E&D� +u=_d� 錑r���j��&D�c��O'X4=��iλ֘��h$D�H�%Ǒ�`�j�K2��s�#D��#�*ŝE P��O$e�4;�=D����e
#e��K�%K:X���'D��8���7O8M���S���$D��X�B�2Ek�T�1�F�8���Sd"D�h��-B�zܼp�2)�X��d(R;D�(�HB�L�d�1�aY
�+��8D� ���~�Q�uHJ�J�H�c�7D����n�x��hQ�&V� Fi+D����.L8Oc$ĺ�dB*=Q��z�#&D�|C����Ҍ܌ O��˗�&D��p���l#�@�%`[�=��D��j)D��)q؄de�5	P`T�4�j�`�&<T�H��쁝:Ɛ����3G���u"O�D��4�
��"G}=(}��"O*5h�C7 2Jp$K���tX!�$��і��t(ڼa����$ЍpB!��1R�P�
���ᲀ"��RH!��4;/���&�H	�J�	��E�4-!�D�nH���Ƙ[�^�c5�ć"!�^�S�82v�b-5A�l�m!�W�u}z��`���8@xjq�E�9�!�$M;�BMj�]�*n � �X�j>!���|���0陊B��Y5dޡ;!�D�>M(r��.�->E���!��W3!�DV8���@V��J$L�(!�DH�U{&"�j@�	lXiR���&R!�DD+A[� p����d0i��ؤL�!�$�X�,	*#�G�Ҁ P/�!�$�&eA(ɹ���6{�M1�MZ4c R�)� 
��Q�D(�Q��_ڔkt�<D�������f��4�ʛ{I� 8��0D����*νz�LuSVe�^j6�zF/-D��{BM�-u�С��Ą0&�E�ҁ+D���PH@�/�J���EX lDa�u�&D� S�F��~߮�7Eđ-�:Y{$D��a��!pm��宖�w8�7�'D�0Y@)��z:V1��#S�f�21�r`$D��S"2V��!�2G5)��;1C7D��S�@�Nf����P.3C�(�DC5D��s'��!��DIm��8�o5D��X$��;U�&-�2I�5
D� 26�6D���,�Y��u���t����M4D�ܻ�'�}>*2�!��ti�m*�H1D��c��_�!gX�[�o�(���+�4D��2�A[V7VQ�0�a~���2D�$���B	�8�wB�#M��r�a1D���J��HF��4Dٰ?��N5D��:�o/����&W��̒׍7D�� z�A��~A�YU�ϬX�Aj�"O
a��D�	�2�+�)Ы�:t�4"O��6�9�N�k�O»0{�b2"O�-Ӕ��a�}3vM>̼�*g"Ovx��K�d|:�AB�0���"O�pB� 5�5�q��u�f��%"O��Y�	�4a�,���!L�C���1�"O�u�TL�T�ؔ��1��XR"O鈶�G?;HՀ%�P;1��4:2"O�3$@��]d�A�&J���$��"O9�W��;����+�:�> XT"O���
1UQ>iS)�:Y�A"O�m�奟�Cv�=3R�� yJ�"OT��a@��|rZ��'��q���"O�d&b1x�hR(���J�"O,=��#�,`4n� }�0��"O�]oT%$�@$�ګR���a�0D� �$�T.Q5���T}�����<D��P�J#-���+R
9� �W�;D����¹D��* Ɲ�udz4@�:D��A7��Ah�Y!p,�:Md����7D�<!��(�j�[2!�"Ģ" 1D���.Y�b�J8#���2'���x��.D�h��L�}/�sTl��l����*D�80qk��R�ī	���)��$=!��׷����Ř",
���M�&L+!�9���� �ZG B!�/f!�d�8���v	"���fJ�.�!�d��.*�%��	�z|���7V�!�ױF&��D��q܅��k�!��а���Ȟ�s
.aa#�P�@�!�D�ch۱�	qj@�� /�$X�!��*	.�]�3M՟jX�Y�C�2�!��_�� �K`X�`v2�
�"��Ag!���ڼ��'!�$E�C�7P!�F���J��ۖ4\N��U�I!l!��w�<8�f�3p>�C��5d!����N��3��L2�$rŢ��D^!��wc493�FO�~b�A!�R�M!�d���Ԉ^�A���`ˏ�j<��
�'�x����ZW��*Q�]5U�l�	�'�8�¶f�<��(��� ����'���	wn˴i�Ɛ���.uL9��'k�Ac�C��C}n�3�,�S(�Y�'�p�B�&T	N�ҽ؆��y�����'�`
B!��U��S�N�$�� �'���[R��#t��gE�M�6|*�'��!�5f/�t9zDe3W�u	�'�8� ��S�S�ݹK	�*�����'B����2�ܰr���Kڭb�'��M�$_DR aS�I��� �'b�)��L� �R�����0M5d5��'���.	�N� r#E��{�"�8�'�d�[2�V�4!��F$oѺ@ �'3��9Bɔ-A󮬃U�h��4"�'U8p̖7.�x�X�Y�4��''% EΝ�d�\u�%��X��Q�'o���B���3~���\&M�@��'8��ӆ@I�m�]�³=�uZ�',�10W��� �饨���8�@"O*��A/�� �깊u�U=С#t"Op���G�jJ\4h7��q����"O�{5�فS��\` K�h�@<�w"Ov�Ui^1}©����6&<�sA"O� ��8A�^�7O��j�B�45��cW"O�=� #f�Ж��55vx0Jw"O��q$�(i�����/�=�W"O��+w�/kwNQ����y��p�"O�AH�n�(((�X�G uxx#�"O����LZ�dV�4�GǤψd��'�t��'�U��&����D�f�5��'gh�X�ׂ?.��2"�Zph���'GBe�7( pg6`������'�&E@�E�̝G?���	�'̄P�� }�]�$`�9� ���'h��B1I��#]���^ò�"�'Pbh�%��/w��D�!"Q�Hu	�'�dI�M[�l}t� ���KWvb�'Q�u���+w:�@�	3A��I��',��y��Y�V0Ha�̃-ࠤ��'Uv=�qHK�%[��
�W<�"+�'�z���g	M-.�R�g�$KW:���'��X��-�PC��1%�/8м|�
�')-X�gˊ>�V�s���6��){
�'�l��D�O�D{#'�>��hI
�'�����?��])��G�K��4��'ώ:�JN���-P�>��Y��'�>Yi5B��w�T�q �A�i�X�'�>Q�b��8i;�d�5h�\)��']�؃b�9'4����Z��,�'=�Ђ7�B���H�IƕX�=i	�'L� ��{��ų���f��1	�'~�]� k_"O�I���O43Ju��'�R�٣�6")��94�ۆ=/J�'2��S��٨] p4�@�	3��C
�'��ypi4S��#0N��5I.)j
�'�
�aqM̽5����� ��dԆ��
�']�<�9g�*D�Y��"OX��(��8~��#"ږ=!2���"OԜz�Hٻ�Na T!͍f\�@R"O� ��&@�1ʤ 	u��7"OVHbྲ�٘ej̀4����C�G�<Qp�r2����^�t$�KP@L�<���[aw:!(@D�5�&P��d�<)��<���(¨�.:�$�r5�Wx�<iSI��(A"�����;FzDS��Vw�<�d���4c.�B�R�����y�<1�(�'[M�	i��D1e�9	CSx�<��_)`������'#�ְY� FY�<y2�̷2�z�(���ά"��S�<��G�5V1A-�#\~8��H�c�<q�J�&`�4��F�R�Q��	�!�U�<g���Xc�X c,4f�*�8��x�<A�e%6Z���H+I�`�[�+D]�<���P�4�ᘤh��Ȇ�BZ�<��a�6Z'��#OE�8@��KR�<�� <ۨ�9τ�~�B	P!lx�<1Wʂ�DǄ(F�<M�x�% P�<7� _�H��X �fp�G*�O�<	uo۷2lv�VEl�L�&��d�<a��S8>�8p�/A�C>�p�a#b�<QWL�'⦵��ܷo
��m�e�<�1��:a�BϷՐ�*��e�<ᵀ@�-�Jy�V��;P9���d�E�<�oC�"�|�Q��b� �s�	�1�y���bT���M��j��=�Ő�yB��7~���'�۷J�f��I܄�y�&�mF��s�(ƵVy�e[5��(�y
� �$��L�^KV9 �_�ʐZ"O>�� f�tL�Raw��""O����W؊Z��04���a�!�b�<92��<I�E�pn)z6 QF�[�<a������XPj�$��$R'YP�<��0<�Ƽ)�灣�^<	�CP�<� �5��H�d�X_j��0��M�<)��B�E�A���9}L�K#DCH�<9d(�)O8F�0�	�53x|��(Xy�<�s�/���+��\���\�ΐv�<QաWf���X������Ǉ�u�<�Ǝ�x)���7�%B,����p�<��)�*�xۣ�Z5q�\��D�<wg��xQ������.���� �Y�<y�@�D���`��Q"S���*OOS�<AI�a��4�D�Lb�r��C�[L�<�Gޝf�-ӱ�c��"�(F]�<!נ#y���P3�C�a��|�4(O_�<�V:e�M�LZI�2���CU�<�ڸVQ<���dgf��"	�J�<���!+h)[Q��0则aC��H�<��M��6::��R<F���a0,Ap�<٢�^�q# h����5o[�Y�Hl�<1�l	�<�\��@T��J��P�<5��#,�^���Ȯ�p�L�<�2�L�:�
�Fӭ�X�w�H�<a���>=�
&���W V!��(�K�<A���s��JQ�'nz� �fO�<Q�%���M���%^2�;��v�<��"�2(0�	�-%vi����r�<iN�$}6��	,�a��_o�<�� �K���T��m�f MB�<a��_"Q0��
�[|(űG�XS�<��(B$T]T��WÅ))�����	�x�<A! �=�Z��צV� �1Aq�<AWbʬs��@��: ��0W-�i�<��bK$u"�Bqa�;4�����MK�<��KŴ%4�;�l�74�f���M�G�<�昦�F<�6dG�E�DIT@SG�<�4�����ԉe�J�Pm(i�!���+4����Êo�=Z���*	�!���.�N�sV�_��h�F�^��!�6�-�,��D׬��C�d�!�D��_Yr��6-W�!�P	���-�!�d��u�$%*�I��lz��$)E10.!���q�xA�"��`a��b�F }!�ߤ)D@�aeJ>O�D�����$zk!�ХI�RbŁ�4��0	 
�I�!�]�=9h&N��F�V�0wI�y�!�dX �FTa`
N�B�H��S*@�!�Ԋ6����Ś�M��v� p�!�DM{�1u��M�d"�ŀ'N�!�҈j��`�P'5PbT%E!��Um��{C���(z������!�)o`�FM�tr<݀�U�@�!��+O�.����ԗ}T><�4�Xw�!��YwcԤ؆L�i����&�Id!�$B�^���+F��.?��9���R!�D�9Qd�)#u!��1=L���c�`<!�D�btf��ǉ��/3ހط%fQ!��X�!b&��x�aa�+�!���Z�R���O�&l��h��;�!�Ę!F��JƮJ2p�d�){�!򄃋~�JP@�'L �8�A@hn!�� �l;��ȢDNr�cB�W��L�B"O6)�p�ӵ9�x��l^�{<%�"O�����^q��m�9jm��Ip"O2�xC���yb'_�iЌ92"O���<&��
�/ߏD"�	p�"O~P
o]� t�������
`��e"O���wf [� ��M����̡�"O$<�d�5**��b����#"O,�C ˖�v*�uJ�օj�8��@"O����/��]H�(N�B�eH�"O�@�",��H�W莚݄LAr"OHh���w���2)�\�2"O��˓��rȨs`��M'�P�7"O�i�1,�>N�³/W�"p�t��"O|�(a,ϑtT�=1s/�4���@"OZ�pC큨R�P�b�C+A�$(�"O�����a�T��ņ��_���"OX�jF&Ib,���ˊ�k��$[�"O�5ՠP/� a�K
�**)�5"OTt���[�7S�hP�IU)��Rv"O�T8-)\LjD��̵=�d@A�"O
�
�
�$f�3F�c���cr"OE���̙:���! �<�90�"O���EɖC�̅�����;�fq0"O�!sf��;yo��ӱ �6��ճ"O��S��QNX�Q2 Y��@0"O�<�bꊰ8���B�0g�$ܲ�"O���Ǐ&8ή�a�������"O�T���
�qGr�a��×$��x�"O.����881� ��g�����"O�Hw�ӭ}���@f 	 n���"O�@�� ��(B6]J���F�yٗ"Of�A�N�'r��`aBO@I3����"O.t{��.'.��!V��'m87"O&H ì\JB%f.?�$��"Ot��6Lu��Y�,�!F�@��"O$�ȂH�H) ��F��Nb��"Oܺ��\[�n��'A��[A��d"OaA!ꊠJ��03T�y�t"O�%���B�_u����dV�9�"OE oޗT�eX%���>�,4��"O��)ӭĔw�:��;|��4q�"O���e�)+����!�Y�s"O*��˛�*�@�/S�עp@�"O��y���8'���
(şe�,�	�'GεrcD�h�@3pdF2^���k
�'�zM�&���&<��K7	�A���A�'x��#rDɮ+ٞ��f��(dM�u��'��hz�$ʇ4Fɺ��
W��q	�'x$��կ�����W�S��h�'X�X���>C>Ƶ�C�<{%�YP�'��)��_)K���n�~�f���'Pq��	+"�@��剱w#�j�'˄����U�Q=\8R���o�``�'�&#�Φ>L���Ő7r�\��'Պ]rb��8���"ap���']��P5�>|��"��hi"�A
�'��\��E&~�X�f1]=N���'~��Z�ύ V��
E7\O�\��'�H��g��Z4��cd۟U�����'���	V�	:w{��20�¿��uY�'��q[�o�1�|�ȄJ�Ĉ�'~�{�ΫX�nX��aM,{:�� �'��-�E5t�u �.��l�Ԍc	��� `�����	#��\�B��72�|��"O��3 ���@I+&����"O��:�D�c5�8��Q���RW"O�T�H�:>0Ab뜬a_h��&"O^�0@��5-F!{7kG�p�2l��"Ox�`�.J;hBi�6����"O��2/F�`~����	�).�H��"O�i���O"�Q�'v����$"O�=��aF�Q�� �O�Z��P"O2xq��ש}R~�AH��r"���"OH�A�@봉��-��)\����"O���&�<P��m���=��0�R"O��8v����I�a�J���"O�)�c��
��0AS�Xb�ī�"O�5��۲�Hܒ ЂD�9�a"O�1�lɤv^�噧�;,<y��"Op1�����Թ�P`��t(h�"OX��L����V����v5pW"O��;�n+s*t��Q�	�����"O*�YFbރ8��*f��:z�JͰ�"O�4��D�p����ۜB����"O�j"�]^�aa�IA2GP�ٱ"Ove���j�#kI�f28|�"O��L�=>�U��l��A���"O�Mr��/���ʗk]�թ�"O�٥ろ`�����
� {�	�"O�sV艁 N��p��3a�r�"O�Iz�o\<u�ЊC�JU_QIt"O���w��5�&�����YZRD�"O(p��`)���Y�D\�trdt "O^%����)[�FY�r�N�` 
��d"OJ��`B5�M���V�O�8E�q"O�e�uϊ%L�!`c�:+�H ��"O~ݩ��H�����~�jj5"O�D ���gZ�����!#n���"O����k"�I2�� <�A�"O�|c	��uWN�PNM����1"O>)��ԋ.d��-&G:*	k2"O�tR�/�&aA�xq�J�|9�s"O�d#�օ�e ���ucDJ�"O����+��ԃE&I�:M�=�"O����Ɏ�"�0УQnI�x0"� ""O�����X$G~f���C�o#��*6"Oz��M�~�mN&><H�"W"O���� #�����*i�8Y�"O�� �F0\L�ArF`���s"OH "���KvB�+Rc�mL9i�"O��b�� ���rd/��n<*h��"O
y�3�%*�ɫWL@8f+����"O2e�1��i8v���k���l,P�"O�0i4��	h�Hk�mV�k��A"O�-��Ú.?�����+_�B���"O&�R�gK_�Xt��9Ϙ���"O1��!*)�>%Ɔ�>��� "O�x��ac�(�Gќ.��YR"O����~���%��7�����l�y�A�7����1j 0+S�a��?�yRAE�$�zt*rg #,�2$[�g��y���9hK�ǥ˺����B%�y2FΎ�B����M�|)�d��m֩�y��V�X��a���9l��m�cNZ��y�Έ1L&	�GV�xD U�����yR���(E��q��t�0R���y�J�f�f9X�� �,q1BȘ<�y
� b)�W�
�&L3��͛D9���"OZ�
��?L��ؑ�<E|��r"OP5 D%�,|,�[LûoN� "O�hq
�<���:pD�(gĜ<0 "O�QxF�J�
���XPD�&�P�PS"Ol��C�R�cڀQH&i��>��)"O��
8:���1�1c���"O���2-I;�:��G�U�^��D�6"OzR��9h��K�Ϙ"=���Ц"O��&&�l:Q�	k���k�"O2�@�jʿ<8�5("��#�T R�"OvD�2,<0�XT��g�aϾy�S"O&Q��(�I\����F�B%t��"O8�t�Nz�z�r7ǈ�H͉�"O�ѓe
خ�4=�B�F�i�Ե��"O`�{��W�R���g�����"O�x�R&�Qb`M�1+D�j�����"OP�3�]5Vd���#6��ē&"O���IĆ^3@8�ew�b�b"O�F !I�6T�Vn+ �pXqt"O<�2�f^�3ܨĻT��� 	�C"O�A;����"�����Sa�Jh�c"O�|9QjO�% �!f�4.b��%"O��QB��4���Pu�4�j�a"O�9$^�H��@4��K&mТ"O�e���=�l18�c�	$�Ma "OpŸ���RX����!�
;���p"O43t,��s�����劷e�)0"O6��0L��I�������@%"O>���?Mr�U�-�/����B"O ��7Dׇo�J�	�6���!�"O�!K�)�r���{�O���$�R"O8�Z��ޱ5^��S�֘/��|��"O> �A�8s�����l�<p��*W"O�+i����a������Q"O��)Q�N�l���r@jJ6v�I�"Ob1��8�2ջ6Z$tb.i�6"O�t��I?:���r�C	&i�"O�����B�t�V�XWL��@g0���"O�9���5�1���Q8(��"O�lrr�fٞ��I�*��=�t"O�I�K�]��"��S�G�4$cT"O���������b�AI5/���e"O!B���5���gK�^T�v"O�����Z�y�I��M�����"O8@���ײ�v���f�}���"O���(�}��W�q^�-�"O"|"� �Cx�\�e�^�XU��q"O�t� J�$:н�T�Š8T��x�"O���H>l�BՋR�7J1["O�B��'`: �� �����"O�	�ʜ"=�,����ۏC�0�2�"O| �cMM�P �UaT�Bـ���"O�`2�G�Eq�T!�%E�x���"O��آ׆2d��Q2��K� �f"O��� ��4W�Sf/��K����"Op1!��>{�ahg ¸�*�"O�����ޥ���O�W�z�ڠ"O�t2�+ҙF?�4B$�۷]�H��"O��� :}�h1�'�Gr��@�"O�<Q�aF�.��� ��n9��F"O �IF��������ԅn���"O�@r���o�:��rM�/���z"O��8r"�>,|���͏�{��)��"O� .�hP�� <� ȀQ��K��]J`"OH2���?*�ȪvG�: ��l�"O���vo�_ކ����_(q4��Q"O���D�`�<[r�J�`$B0�"O��S��ʅ	��yAmT%}�P�2"O�x���.�2�9�N�m]p5:�"O�HZ��N�b�S��\�<���q"O�������3�Ȅ�֮��g"O2\�,طYP��aH��Ӯ���"O��h#��<��,��î�����"O2�b���a��D�0t��$Q"O\A��Ɋ'*q�0�I�#Fhe�&"O��K��]%B��%h'��n��8��y��H4u�0&����qԢڐ�y���+	l�����y��q��D_��yr��b>V8k��БA�JX�mY��yB&�>B�̴�%��H� �b�S�y2�f�D��A,�?>v���R��yR��%�Xݢ���%�����/
�yR�?t������-d(�4	��yҪ�*O�,�S��I����dl�
�y�I�w9��`MRD�Q�0�y�Q����N���� ���-�y�)�%O�	��N��tހ]����	�y��\���9h������yRd��
9b�aY>fX]�t(Q��y�3}�0�Ѥ��eڌ����6�y�*u�rUZ�*�&b`� �#�y�,Lg`i� ܱ~���S�B��y��O�gR�@����@���4�y(I��\�p/� ݪ�;!]��y�ƅ����(dN�/q��:G���y"�N�c��k��7��KΗ�y�!Zr�0�$(�-����L�ygF)���"�dX���G��yK�F����wGߘN�Q0�	�?�yr# �B�M�p���#C�Д��'���EyJ|2��ԫ<����%��Xi�A�7Ä`�<S-Έ(SZtHd����P��σ��HO �}�G�z��`ZM��ځ�K�?��ȓ)LҥA�/�'(�49�]�(|�͓��?�u�Ժ?�}x*�_�:u*�+@W�<At��P~�He�+d�}زcVJ�<Qg��~:�@��A�N����uwў"~�	�JMzQ�� 12����_����#�ɑ|K�l �M�p����[6U/B�ɰt��ӋV�w�L�80)�$>�C�I M� ��pL,s>�:qKT/+_tB��<�"��A�V�d��7"��B�	p*u1�)ȸQ��y�D�N�gf�B�I��-�5�Y8f4�lr�	�d�Z��d:�&K2ٳ����d��8�&[?���ȓZ8ɛ��G7.�<���djf���'1j�Gy��ɜ���a��&�3]c�Qi&)�:|�!��L�
��R���t��i���z��'�8��dQ�a�64�C-����0�R��}!����W�9<���  �<�ȓ��2ю�!B�D����Ee�����
��܈&�l�x��@<;R�ȓ*��3E�6�����	ٞz��P�'�ў"}�%da�`p;�ܛN�\��C.�{�<)�B�� lp��A^���K�t�<�T�\n�"f��"�Z)G$Ct�<����87��@���<
�d�t�<� ���'�N-���^u��HÌ+4��P�B.A�5� +ډ=��Cv�9D�dҶ��C��;ǈԓ	0���Q�*D�hPAI�'*&�@��U��uRp�*D�x��I�Z�� ��O�(Lr-3�B*D�4��:$ʁ8�D��T�4%�W�"���<��!�N�PPn�;A������h�<�`��;1�̹j�ő�cR�����O�<���D���mk��K	�¹�NM�<�FP�|cB�'�X0tݪ��K�<�5GD�zM�N�;w��I�R�D�<� ���z�{�f�4��� #Q|�<����fL��⚯X�R�Z�o|�<��	z�
���,-HT��гa�t�<��bٙ&Db���L¥��q��)DG?����.]������-~`
!s��ͩW*4B�ɭe���2C�A�V���͍G��C䉷z
m���X��L�-H�ͲC�.*��`�	%�"�?�C�	95��1�@ˇ��: r0
#?R�B�I/-�ڸU�C��:u��[�B�	�sƞ�8'���@o��B7,^�"<9�'��?A"��V���`-ߪY8`o=D�d�f�������e�Q�l;D��CЁ��%�� ц�";Ar<�o9򓥨�Bq�NN�u����"��,�"OYS�/�2[���!�` +,Ќ�"OX�ק��5j�Y�b�Z�@A3�"O�Рp'�N�vIV+2'���"O2q�b�� �Az���m_�t2�"Oz����e�� �$!U��"O&	���*^��`smτDܬ��g"OTiZ��H*(����M՜�r�8���!lO��)�ʉpP��{&��P�"Qi��	��<a�P�Bx��!��<	��y�)�{�<9�������Ȕ8q���-�����'n��P���Z $H����5��;�'�(�l؎i�}����)��2
�'�ll!�E%��;$�V�N�v=c	�'�x|�b�N�|2(���0E6^%*
�'�ZYH�@�bAp�9+�����O���&<�& Z���]`:�[V�UW!򄌻i	r������\���L�!�d�!�e��m@�+�F�#@i�F�{R�$�4.�XH􀌫�vd{��(�"�$/<O�C��|(K`,sv�;�"Ob5�Pƀh2X��
Liʁ�"O���pD_6���	�44� 40��0���i�VUi�� ��ǬA+zPB�I�+�dH�k��J .\��*J�c�B�� [.\qQ��Zq�q"��1P���T�I�e�q	�H?�2�)�i�rB�Ip<Z ��)����QFG�c���|y���~*��B�5[w�OR�!��K�R�<% Z���Q��]e��y�TʒK�<���.�@��1l&{p�Q�.�]�< .�]�(b��N�ŰlA�@u�<	��V�9?Dt��C^���� �Be�'nў�'#qĕ�$hV�Q�T��#�U}z%��F�p�;a�A�S�$�1��ڿ&�>Ʌȓ�,AcT�آ3�l���oο;M9��q6 �o�Zl�Uف�ֻ0�:��<���	8$!���5)�8U�|Q'�0:�!�$O�aĝ`Q���R�Zu&B�C�!�� ؑ�!�ߝ1��X�j]Pơ���'1OD��&�eDY)U�� #S��#n�˓�hOQ>=��b09�)c
$�FeBc�<D�D��/A|O����J��a�	8D���T�<+X�hrLe����@�v�`����G�fe�UI����9��
8x%�B�	����@)�e,�كD	ȈSI�C�	�4V�`a�:z���ɒB�PB�I����Ђ��3(V ����e���&��P��R�N���u�֨��7	)D��[PJD0�(��j@^�`c�(D��Y�(ڣA�\)o��	V6<��İ�����?xD����1�����n�B�əHir�೨�S���8'�@�`�B�	�}j.LH�M@	?���B�D���B�
>-�2�e�(6�Q�7��O�d��hOQ>QЃ`$���$Bͪ�.t���9D�x�bΞ"U�X�l��H9p�g=D�̊�&,:4�PS��
����";D�����=���[����|":D�t�v"�<KѦV�	Ҽ����9D�(BE�=WT�w�2z?tY�-*���^<8FNU�q��D�P��<�ЄiQ"O�xzf*V���թG����z�O�<t��,��@�` bA�52�J ��'D�Q�3��?)r�� �)2DE+�''8��N,��� G��&�^( �'�d(F�'<1�LHŎݫ.��1�	�'�0\��,8c(��$�M�8F،��'.�����&N6� �oP=,�^p�'�f�a�F�a�����#�"GBt�'�����F�z������,*8k�'��b��Cx�K��^%�r�'V  �O�3U�z2�։���+�'��}�0D��̔ͩ��E�.8�
�'�z)3�R+buԸ�F*�5g�.�2
�'| ��X�)�
��C�%g�ʔ;	�'r��k	Ю
�N���=dc\X	�'+N)�fNF;4�2Yq&�X�����'�\1���}��T��	Y�>���'J�
����0�D��JK(W�uK�'3�y@ �����i���G4@��'	 �q��9$ҽ��gO�G,p��'�D�s� �,�v}����<���'W�%CJ�Q bQ���x@�0�'[ę
�N�*�%�I2��s0��z�<���Q8H��ĩ�)ZL��ѻ�J@�<�DЦ-��) ���nҢA���}�<A�!�$GSa,\ip�9S/
{�<���z�j��f��~�p1H6f�w�<��B�?�ڵ"6%��w�؀p��Lp�<�c ڍF��	b!єs���pƭ�m�<���1)\(#e<fZL C��i�<�ʊ�R�t�U��<��dk���b�<��KL�e���
N���e�[�<��(^��*�~0��82� m�<p��9Aʵ���N�ͨB Mm�<�S	��V(�#��:�pZ���o�<)��K�y2���( _�4��h�h�<A�8=�4<�IK�<x*e�L�<�Amô+�x\�s)O�k�a����F�<��I�lNY�� !h����]DC�I4n�(��(�-O��6A��x�@C�+���2T�E�D�5ᒛd�ZB�)� �y�F�Q�{Wty�%sZYXD"O:����%j�}��c�Wh�d�V"O��+#��6.%��'�:e����"O����,�vm�Ɵ�xdDM�'"OF�av�D�}o�,��U�F�{�D�+R�X���U�a�R����HW1O
U:�A�;�.�84C��\i�"O$�9�E�,��h0��&���S�"O���`O!}���5n��=ZVD��"O�� B/KZPR�`�o\)EC�+�"OH��$l^:	 Gj�ҭb�g6D��i�#?
¨��f��!����*O���֫lD�\Ǎϗ�ܙ��"O\�xGN�l3>УcLX�*ƨh�5"OL�s�<uҬh�)�)e�"�"O� ����8[�9��hB1y���:d"O�	�Q��{��ӑ�Z����k"O��3��{��pƅ&K�t�0"OL���7 *��p���\�	"O4�!B �`ml� ���}4��u"O�T0�#����%b��eS�"ON������p��L_LDx�Q�"O�|��JP2�\ D*Q�ANvH6"O�]�� ^7�xE�����#����"O6���]:i�\�ۖH�Y֬��"O���(
z{|�R��o��y�d"O���n[���\�����bH�u"O�� w����*΃2�B-��"O&��0G�I2!Z#�H�q"O�EQR�F?m�8	��ǋ�}�0h!�"OX8X�
��D�|`����lNP!�"O�9��j[��<�s��Z\���`"O�g�R��;���2V���V�'g(m���
�"%s��\mטG�������퉡t���z�J$�rU �8D�@��'�		��b�	&�<�)��ل<z��0�`N�E��pK��(��wb!���$�^e`�%�5��]@G�w��|RaA�cP�%��Bט��5B�S0�ց���ְtPmJ�,�F�<�0���)8nd[� 5O�����̙obJ$���p�����ቼX%��O0�ʈpT�U�7�v�+�%q�����-5�HV"��a�E�61�@�v�6��4�M�w(h����W�1AtĠ6���TM	s!z���45Hd��I��H̐8�BV�I�xm�Ok�	N�%���6�� ��?�!򄜇ex��i4F��x&�;��	��U &��@`V`@��8w*tȀ�Oy��Q�Ts0�c0��G}�A�\����T2�<P)�LI���=1c	�F��P�3&S�Gvv�)�k �;���=?�����'�ҳ���>���˚?{l�E}ŕ&���k�C�� ���i���'�8��F˨J!qQ'�F�'�50���$m���T�� ,���	di)U
v��*Z�o�^ ��M��p?!w��!.<|m��yǲ�`��[8paD<�#�F�m⇌Z�c�[�FE�(1fYs��Ѥzö�������Y�D����.B�<����t�<)!��9p��D�� QՐlz�/�3��K'��?<5��$�L�S9r��`�3 ңW؎PQ����@�h�8Zy ��@�6-t ��g"�d�6,v��'E�b���GR [�d�2�|r0�(d�W O%rA�	:]'�|�t�N�2 ��B��R�������J�`��ȃ�H(Q�DI�*K�}�86�X�\Ƙp�"B�&����JP�a��E�lɦ,&d"J�3{�!P�əZˀH��!"����G��]ɐ�
a ��u߮\��)�2;t�`���'t�!a		�(�;s&2;���4m����0�!S=6l`��ɀ�J��dc��H:�c��V2;���D�����Ȉ��ִ2�Z�s5�%W>���fJl���]*:�&�ʑm� Wl��$��+f,�"�Uz�q��h�� G�	p0bGY"&�a��'���Q�ě�.j0ɵB�Pq�M��JH�5��ơ
��:�l��@���.�R1���
)�ÊR:(Z��� `��0
Q1?�(���!�h�L0��C
ƭ��錼i6EÈO�^�(�� ��9N����F�7������	ؑ��-��!؎0��VY-�up��:��I2���& |I�e�Xp�����
 �&א9HB@��^"�E W�
:�
���{Tp@��C	��c1Lbb���ǅA�f�6�,-^ȹÓxw�m)0,�S���Kө�&��lx5�_�q�<P0����5�^�z�nO�Vq��W̃V���k�	�-#��D(��^	u�,xXU+�}q���e��	�����O��a 
�g�ht�H�3hH����^�}j�IqDT�<�@Ԡu \�*=��"�R�)��/�TI�qNӼ1F��p�ʅA-t�B�N��$�+3�ȑX�>̺��[�D����fĒ�剓m�i`秞D,dS���5�p�f�ux�m��y2N0��L�gn2�ʩ�R�L�-�~�a��x��	�i.��®ֳ��p��@����� �!ɤC
K��I��ʹjv �Ĥ_J'*��/�5�����BL��d�i��-�c��w��\�qȈ=&�^�#�b�2I���vD�f�'�	�1!��x#Y=n�N�	�/@�'NΙ1!�S;�� �L�
?���u��$"��	�Ý�Mc�'W�C�fE�D�D�8�n���ػ|x5#�VJJ��j�2O�T��ř�)�L1�P�� '��(G~���.�Di���^=�%g�%p]ɇɁ����q�$��f��}�Ļ���2�iBLA�iTE��� ?������S�#���E�{�l��3
������I��`�6���96eS�8>���F,{H�k�؛dX$U�C��p��1���m����ի"X��*�m7%A��
��^�:�aU>i�8���Qb���A��)!P�'�P�6�N0u�q0�C�4_�<A�m�4k��S0G� ?a�%���a��l���2 x�MHp���[�4A�͍�i�� A�ѓ9	����Хsj�a�2��3^
�s�λ A�_V8�p1d�vt���*��8[�Mi�!�;��1�G
u�@��#���H�3��uq��תԞ?V�]A��:�˒:T�����l�D�Jc�
=6�T�I˓R�0�2�`T{n�2�]�pډ�W���6A����n_�o���%�x�x���X=Z���f-O�^ޅlZ/`��k=uи�Qf끹���zWH�?�*��ѫ[� !����ɭu�괡�Ø��Á�fy�R��"Eu�<����_#F�`��>b�Ԅa�~�"��5B����&�M�Bz� �G�Ҹ\'B�<��F��Nr��&я+��%sdCY?�C���5�d`y��X���x)s��?M�`{SHƖu��!����`K�$�-W̓��u�ə%CZO�����><u�(��0=11�Ѽy�Ƒ0"n�3��dI����|���	݋&���Zs�̗&�x��ĝBN/3��L�L�?�2�1G��ai��A#�D���#ba��o(��P3��[��ә(�r���AR�;-�ᣎ��e�a��y�����扰x��`9��&	��! ��F��;b	�K�؝�F����O|��[��N�α��쑉>7v�Y��k�mq� ���NyhVHI74Z>ݩ� �T��	3BH���iN4º�R �DCh��r%*G�x�PE̽Ho�$�)n@����/k�a2��ċ"2L|����Q6|�V>5S�f� v^�bgk�6�h(�sAH�Uj�xׅ!w�����x?: Ѕ˔縘j��ɳtDα��C�^�D��q�K�@u��~:C�֒��1pL��ګ9j��[B���sv�䑓�Z�/1a�E��Tt�X�cA�%Z�#
ʺS�����Ŕ;j@�U+�)9���+�nM/qJ^D��	hL�r�j 1����u��*((�?!�KU�6����n� 0謬��O����+�]��EI2��(E�0��'OT�#jB��~ ��f�"g�9��O2�X��ͅ+GȐc��Ɋ����y��n�mu��2e h% �B&"O�I��T5	�|�
0��Fs����:��Fq������|��J
)�!YCǍ/B����P�y���3>D)��͞$�Ρ{�Ɍ��y��qAxՙ  �m�ɒSb3�y2���@I~}�iV��k���y��pd�5A���=V���X?�yr� �hL�0�`d7*x��q�ń�yrJ8Lp\ʇ+BQP`�!����yriHycE ��D��Ԛ��à�y"a�089����2Z����
��y��	) ��p�I�"4��m���yb�D�_7*�c��krh
�GP��y���dMA���Z&�YT�O��yR!�#L�\:c@��<��t ���y�&X�(�F�Z��-?0
�
��P��y�lJ!na���g[�\���w#Z��y�,U�h@p@��H���CP&�y�`�T�:5q@�4d\�9�j:�yB��S�L���]~�JS/ۚ�y�a�^��Bm� b����u�Έ�y��5X�p�Ѣ�?f�P���AF��y�풣QL��
�b�а�;���y����j��	�r`B0)�-*tO��y�N���x��62�Q��Y��y��=2���S	Є�B���=�y��J�dR�<;��B�����0�$�yRJ�"�� a�o�,Ѯ �gʊ��y�l�L������TD�h�G���y2NG�-l�ɺ���	|�&=kW��yȋ^ļ-�g˰|��YceW1�y��0!X�p8���r��2i���yR�ϋ&�~��g�G+s�h
�*Ő�yb�E)�^�;".�+$x� �*3�yBD[���@��%Vx��1'N}�<� �Ps���	`�xs� 2/f|�q"O�ųao�W�x�
��/4��"On�r�ߌm�*���]�=T���"O�D���/%�̵�gN�1�͑�"Obȣ���
�#a���Ĩ�%"Ob�R��^3:���g��`�*"O!	��%L(�	��#s�tK�"OE�������u#�q��Z�"O�JAfU��X93��@M�҈a�"O�A����-���{@�$w�e#"OJ�W�t+���`͈8YP�
�"O@8���8� i�j3B�؃�"O�CBO��~�8D�E+A�G�<��"OXq@���7*�L�)B,�f��q"O�t�`%��ChM��z���K_�<a���6,���۹ho|�`Ca�T�<�ӣ� �PqISDޏN�a��R�<%��:�*�w���u�|IBƓg�<��CE*��@ S ��&(ϓW�<���*������R|�}HЏ�P�<ɴD¢5�v�`�o^r��=���S�<���@�Uc����N�EÆ�d�P�<�fW�S6�=ӯ�Df�"��k�<��P3,Ryp���S�0�j�<�1+�h�<aR�
><<���ԥK}�<��)��B� -J &V�Y�T]
��e�<�㦀�Tj)c��1���C�Ņf�<af㍒FtR鈖�y�ӆb�<���<-d�t�ʝ��蒵ir�<A�/_�}�&�ŨA�.�*�e��K�<Q���D� I�"�J6{Ba	"DX�<Y��w�IZ���#���Zl�<!0�6�mQ��R�p�H�P��i�<!��^������G0O�2�9`�m�<��+3[��b��JJ��+�B�<�%���F���@�;=�TX���P�<�N��V��q��Q��H���j�<Iv@�6���%f��l���XChUh�<��K�FV@Pp��(B1�D�Bh�<i�k����EP������
#BXd�<�Dk	 p_ZՒ�皓7}�*t�<�%J:?� ���h`�3b�H�<�&����Ag1I2�l��ȃ~�<Y�m�	���mL
�%��_]�<qF�ų8�����5!��g�<�6�ȍe�ZҭݠG2���hv�<� �H�JZ�7��A#��foY�<�&V��}��c�:v��oI�mB!�W���z��3t��8a�N5t?!�d@쪭�U萑S]�*`O�1!�$�+g�8��� XD38�
�ُn!�$�1h���OH�q"��	����!�$��C�|�UI�- �ء���p�!��V�V��$�ϋ�a��4��S�!�H�T��������@{�F�l�!�9e�x���	z�pi��fѲM�!�$E�h�jp��Zn�:U�Q/tI!���#�f%��h���q�ʹO!��N�h�n`z��EB���Z��|�!��;V�-��cN:8x0I�s���Pw!�ċ�Ia`�@�g��-g(����;^!�D!v�C�V�T��A��:!�D�`���R!7��â�O#'!����:e�5*��tF �13��,~�!�� ��⣉_��>��r�'m��+ "O��2fiS�z�>���,ʷ{���"O@�bk�4�n9j]�_�����"O���FF�)ۃ*�#`�	��"O�Qp��_�2�񀙱*X�x0�"O���]�X�9yP��{+�X�"Op@������س
��7f��V"O��u�G���5CC�:@ ��3"Odq����;dZ�qIr'`��q"O�ɒHۮ���B�W�*��4"O་����[`�����(a���"O�u@thR��+�6\ј�"OjY����p����j��:�#�"O��@v�$Q��Y')9IHu"O4{d쎉r��U
憛���q"OX4�"��*u�|��"� +h �I"Oh=kM��}BZT��CP<S�$��"O���7��2�ꠊ��n"��"O�`�+���q��Sxy��b"OL%���w~~�b���Bh8�"O�5Z���V�T8V�)e� �"O�iaQ���PLr!(�4iR�a t"O�5���^,�f����)y���"O���H�k��H�S����"Oh��"�J�"IT������]?!�D�2��(#�H�IP5+���r!�$�%̦�����$�ܡ�bh�+c�!�b׶@�e��,�@�xC��2^�!��U<y��B��W�a��ؠ��+}A!��ì��([X�����y�����'H�Q" �������5vdea�'����Dg�f��XR����8�N��
�'Œ���gV"��'F�>B����'�|c$���Rɀ���D�-��'���pq&FRX�d
� �+N���I�'쨘��O;��k %&w��
��a+��锃Z�R�i*aG��q���X�O�"l	&W.56���l�"O$�sGV�)l��:�`ۈNtA��,=sl媲fX*	��ȴ�x��S�7�T�X�yBn\�W��T*� Oqc����-�?�p>9Ç˶3�L�+�(U�=�d;����A�V���.}�m�@�`x{���i�,����'fB��P��(�$2x�+�]�'�fՂ���3��{�5�nي۴P2=��N��r霡 �6a�}�3
�!�\�&��%KԙIR��`R�G� ���a kX�V�Ѵe��"mj�@���4��E���KQ��'�y��I�1�4��ЈY�"k�Qc���yҷ�D]�h��a�$��,�m"Zܩ��7)����C3O����FQ�bh )d�2(�DLH����φ1kdx����s��۴����{��:N���1K�7f�d�C DrH�;	� g�����i��G�(4*�'�?e��!8f���~��$p��38���Ǆ2�~���d�$��O����Ҁi>LHBAJh�*��IF 8�fú1<V���G�=P*���u��KC�8|�~2�(K�.D8vkG ;HX}��dT%���4N�d�h8�sd��8E\iZ�k��L�4pP��8NPu�'�yg�Řt{j](��(��Dk2��+�y�g�E���"��Z�{0H��IT�;tl�2ċ^/Q��=� �Ry���D���juo }=t�!�W?���R�7�ܤ�c�N�h�`�(�Z�I N�l�p�h�i�*-jc��*1:��do�C�4��v
����Dڗ�MJ!�X����8�4����&xDĸ���J����so�)
���>aG�οv�6;GM�!u:y�tJ� t���K��S�q���0gSN�b"ת=s�()S���$x I��jעp������2L!�� ���3R_Ɓ��aF~��4�T�<�OR=I�j��E���uO�W�� ��B5p��!UXl��/�)c|x��i�RnB�E/~�^�jV��L�(,@ՁG��b�Ȅ^���s&X}TI��ɖ:@*8��0�n��Ӫ�<q�nї_�i�G�-�
Di���3�U�U���uy�ђq�sE I���[�1g�\��xw�O�H���"<;^�*u�A>t�,�^��`�k4��q :>�$(�S�Xy; o\&�����O�;�Y���S#D@�R��"j;���3�Q�H�k���T��uu�{��\k��dL�Z�4��� �c�~��҆�,�и�U,��c��+n*�B��
]�*��1��0d�f葢f�-���)әX
(�օS��>}�B���$��@��0>ei�/�x<��*VN([d� ����mG�A��0�B��Dd�,����mǲD��(�"E0@o�h�L��W�`s� ]I#4\�U$��(���z!�Ɍfj�T���Q5�F���
D�FX��5� @��ZR*�&L����E��~}(֐V� A�d������b��A#w�lQE��%JP`�کO� ���{0�9
T���ZH�l2w_��8��_kt�B)�>��ٸ�%�f�����WѦ�ӟ'�v�w �S*L@F��	%���)���x(�Bu��g �`�H�s�џ�b��ֶ@=|�
s͞)��i���tYcc�+6jn�Q,
��Qow�d�j�M�!;�-kB�S�Z(������k�Ȣs�O/XaV�z�M	�.���I/�4!��BB��34�#�"xre��A�"\d��
�B�\M��0 P�.�T�S�(A�C�i�TjO��$qВ�E�L����ҟD�|�C%U(��OmEbڱOv ���OP�J��g�O�"H�`ň���d��L�4�b����^�D!K�h���2���I�<t��%I�qO:����
D8�&J(WX�5�Q���0.�S��$S�C�^�>eZSC���xq�J0A1\X�%�ҝT/P��+q�h+ cϺC��1�@�]
�*�H���=�Q�߆d�8T;�BU�~����Jї��uxVMô -Z�G�ȯE�Y��Ka�"`C@��x��
�
������CP0��0�ԡ��-�Y���YH<$,	�|:�qyAE�!\2�q���>PI�đc�]�8��C5OY��U�	<�aY�� ^6�m�dE]�UB����CX#z;��cG4-!X�:w��'o��yrg�4,#\�*W�B�n���CB#d�y�%ض&0u3$�9;(4���ZQQ�Q�⒴D=��ˣ ��o�5��Ď��2��M�- ���aD-VQ����Ƀ�)�>�� �8Xب�%O9�4�#aBD��B���"�t�I�t�ҿ)^�����9�p>�s��3یŘv�e.v�s��SU?�&�5fbA�\�3���ѷ��k�xx�&��2ڡc�ٟ� ӦE�2UL�}��Eb�2�3�"O��Q���"}�D@%�]5��mH 噘BD`�yb�	�S/�]�̞X��Y��&�"��[=`�(��w3N��"$@��p�	i��3�'�OH��As���Yo�� E� P��2SO҃Ȑ-�`&މd]r(JuK�7�6��b�Dy"����� Vi�Mw�p��
�ݨO�9k`�f�L��� �2����Um]3i\�a�<T�9���(�(\i�&��5�s>�O`��#�_q�� a'ع bf�`��O`���ي>��)A�#G1���!���YZ���sL\�01�S�xΐ�T�
o��I��2�zB��1I�x��d\�L����s��>s�d��\/N���ҳl�=y�O� ����%y�(�TԤ����3� a�l��gޔe��	2��UKWIR�+��uAĠK�J�:퉆�K�W�(}��h�G
�$���S�i��i%��w�'�J<d�L�a�-��&kv�Y��P�04�@����A���1$e>��l�H���� ��Hjz!b��<D� "���*�>\a3(A�s:xT�$�7?��P�N�|���	�/%C�~r� T� X��t��=���p�G]l�<��,�?f�f���#��g	�(����͘'� �ըR`�g�I�$X��m�%t� �Ȑj��*��B�	��:��m�N���F��U�C��(�{���=s � J�6��B�ɟ���j��ZR�ʝ�Ï
l��B�	$&\�9Idnx��8��%�B䉦v��Cǟ)����4�ȾV��B�ɴ(�ȁ���M9l�p�C�bӨ@P�B��0����v����iqsM��lX!��"@k޹�âU>p\� I�j�Q-!��f+PP�F^�a:�eh�*�(!�d��(�
4�DP(N�F�kw(VY!�$
���%P�Q�4h�Fȟ[!�D�?}���@�J�u(������t�!���;.�RIp�A�2�XU�O�o�!��La��:�	�\
x��C�D�C�!�:W��v�5U㦰�&A�  �!��.�0[ӍS�r{��0'�ܝ7n!��O�\E�Ν.����o�<h!�d��k"��٤*�o��ED
�G!�ر	�V�cW	�,7R$�r�7�!�$W�/�,�[d�HoD@�b�Oɂk�!�$�
�򭈵)IgC����-�8}�!�D�-Qp8�GMG+'X(Ң� �,�!򤒵,�>�5F��&�}�1�O�!�ĚH�x�F�-�ѩ�R!�I�4z�5�U�4�!����!򄝢t�8�s	L�("^��t�q$!�Ӟ6F�8򄕺
~-�T��= �!�$�!U�L��Ę+�P�0��_�!�� hp�a��>��i"���
P���"O� ��
�P��Q	�o���"O���
�J��as���H�|4�"O�<��
�.f:`��(گUH�;"O�)��!�;��܋�U�W&����"O��p6��9�iKSd�C*��"O�l�4��xY��G�+oZ�,!��<� ���+82��N�,$�!���h)x]��* -}�r����!�5Y��%���E�<�q��{�!�d9��SN�0�XZU'��{�!�$��F~鷠ܲu�l�U�4�!�Q $7]�"��N�HuZ�%�c#!��a���  ��<�RQ#RD��u!�C+;b���	�V�H�(BԘx�!�D��kbP����g��-�A��T�!�D��$�|�+A�T�8w�@�!� 
!��U�/��L�ײj{�!`d�̾!��R�r�|��Wj��=��`�"�!�$ӳ,��(*Au����N�u]!����Q�ħR#[m.ԉ�� X!����xx���E��Б�F�I�<�!�^�挚uūb�Ы	�n�!�$B�`��%�V����R�i��S�B;!�!�(\X�G؂Z@��g�
d<!��Z�pFjY� �ɏKAʡ"�K�<!���f�H��U+ԭs��Q�e��2�!�$=���7����`�!��`!��}�
�*�S5G:���L��!�ǂcҜ�dD��1n:ac�Μ�-�!�W:@�L�"sG��`����� 	�!�ĈW��Y#����UztEK!�;a�9QY��c�K��y9Լ{V"O��Ib�ޮ*�x �H�>'�0q*Ox�[b�_'��$���H�=�hݲ	�'{X�S�+���X��!
%/hЉ�	�'" b�@�1�, ����S���
�'w.(VJ4o$�y�F�,IBZ�9
�'*���&Ā'0j�#��ݻU.DPh�'֢X��l*�VL9A8NBx9�'��8�򂟖e�t��T�t��'����F.A�U��(��F�#g�
<i�'Hh5�䎂�c��LIp�����xy
�'����u��c��Tv
pX�',�E��@�B��aEF�c�����'h~)�#�ڲA	�آ��7]�8���'��UI���"Fz��p�&��H� )��'	6aÌ#h=2.�4�*d��'($yZB#�;4@^5��ս$7l�I�'�m���м4������&)�ܹ�'!&�X���hдXpBiO��2�
�'$�z�H��d��J�N�$��'_�1���C�q��ؓՊ���'�~�C���2��<B�6iH��q�'���D�u/n���1��1	�'�j���STt��#�[�	 �'"��H �҈e ɳ��opҔ��'���R��n�8�H��Ϭ��`�
�'E،2W%ŒD�ݫҡ�/�c
�'�� �#�ѝW�֌0�#�����	�'�Td����eݲ�O��})��s	�'�f��@]�/c�+ܔP�Z	�'Ǌ0U�n��H��+��S8�$�''&��͙�pؠ2i��R=3��� ��`���1زc���2�@"O�%Ӆh�fz ȤL�7{"�R�"O��@6�P1<ڕ� �";��x�"O��r�P�B h�K"�G�;��ib7"O��K5�ؿ�}�j��pJô>P0)��q�^0�TK�45IL�`' =s弸�ȓV�&����O����Fm�c�<u��6�h��`T,u�r$�A�K)}���  z�܎PX �qœ�(�n����m���]�:�~U��e�k2|,�ȓ���ٳa���0@K�B�B��a�ȓ5�����(�a�أ+ud��[��-Y�b��S�X�Âh��n,�̜T��M�c�Ԑ���G�8������	����2h���	H���;���� ���l����p!� z��'�vd6�����7|�q�Q��8@@�B���:>�y�����0|�V˘(�����S�4A15`�R�~����l)��(����|و��3K��9� ��>	sGր}r2b��z�NJ>2�,��*­k�d`x��Q�<�3��Z� �nڌ�v=����:��H������֬m`��$��?:��c
*-]n���&֊���?ɮ�ؘO��9���	ti;Bi����X����~�[�@2�C}>�cd�GB��E��]P�c�%�ص�T�%mb�R������!K�[�C8��)�ӷR}L��&��:�ҡF��W���'8p��c͢E�1O��0lC�FHn/�����>����+��ts��_<J����蟸Apɕ4D,���/D"�>�:��i ����8��O�Y�''���A��=��%� ��E{�_}}"X���'~����E	��i��ub�J��4�>���Ҵ5���*7F�()W�� @(ȘoOaq�΁H�	1ޜ0���ԟ�	�`�0f��S���rOU_�X˓|[L��J~r�:O �A�kڧi���L�/�@�f�'��y�&�O|= -O�i/��&r�P�!���&�J�E�e�Hh*g.����&Q��$?�SR0A��?������\�h��H
G��B?qD��LW������$6m1 !�5C�H-"tTL�#?tv�O꬐&gN�~�
� N��>M��Ct�����	"�ʐY���<A��K�#&RF9}J?�A���&�����0v@Γ�b����<Q�y*�qO���#|�̌��J�=: ��G��y��0|z�a��Sn����NC� �N�!�w�'�L��S�2�^�|�'Ԭ��a^<i�
đm?��qE,��H!�D߷	'�Cj_�l#@�`2�Z T!�$���T1afY6������7d�!��]�7���QV�S�,��٫�P?Q�!�d��)k�QB!&�(���©�h!��2_0M��0vK�L����'I��!��lî9�郣@-b!`�'�B�#�#ԅYݐA#5�ّ>l� �'{�I�b#�UfL�`ބ�I��'C��"�(P%!�$��'�* ��'�n�ɑ��`o�	1��7N5+�'9�vkD�M�2M�FٳEi�;�'��$YR.E� y�Ó�Q ؉��'a����d���Oxp�(G��y��8}L�G~}�<�v�b�<���RE7�Q,�:k���di�I�<	�����Nj#���1D��j�B�<i�nK�]��|R���,Ʈ�m�<��.T�!����J�&g�n8��a�<q�&ѴbJt�eO�!0�t���CE�<�Fó`s��B��pI�|y֣�D�<I�͇�a�r�02l�se�I!�KB�<ɢ�I�_�آr��7+��dF�A�<Q0͊�!Z�쩐�:�X8)�o�}�<f�.k��
�b #a2���i�w�<�@ͽ5�I��G�3|�x��Hm�<9���h�t��ؗnHx���r�<�4��x�x�:���Lz�L�7�E�<� ���&�a�R(a�M�j\�aq"O�=q��?x�ȥ�PD�ZnQ�V"O8�����L��(� F�3Q���"O��`3�
���$��\*>��#"Of��3�_�Tʠx#���ڰ`7"Ol8����S��pR1�T()��+�"O"PRD�G�[.��j��I+5"O�M��
My\UjS����h��"O�e*C`� m��C�o��?��8�"O�p�Fc\,�<a��O�nx��)D"OV����@�8YfL�tAE
p�*S"O���I��3 �ü]@R"O�ua��Ǣ3O(�a��9��}��"O�*f�ٰ
ԡ'�o�^Qd"O��C��N��� ׄ���v��"O�̨��M�MnvA0Ɓ�f4���;D�Pʄ-E	|�bYr&�K]~����c9D�P���+ِ$�Q� R^p��i;D���0��%���Ӣ,v�1�c"9D�|j����U!0B� 'T��8�(:D��p�
�B��R�ޡ%18�s�o7D���Ѓ��ڡb��RL92�$8D�����ۊn�f�
���T 5D����x|N%���X�I(88rDg%D��д�̐�q3R ��^ �SE�'D���`iTO�Q� l@;%p�	C�.(D�$�U��/x��RO]%\ D2��+D�8J-�#=��`�f�;ƚ���(D���$a�.�iz�_�%.3B)%D��".�2����E��}���7D�8a�$#B-B�� 7L��`���5D��;�l�$TR��ؿq@�d��� D��@����O�q��QLr�U{��"D��꠬;|渁K�LN�o�|��3D��b&pf�@�*@*Y�}�$?D���ҋ)<Z͘G!A4��%Ʌ�9D�@���T�3n]�>[��V
8D�@��+�]�zp[���w����(6D�D�@,ԄV�S2�ܘA�����3D�l(Ї�69x8����(KYB!��P>\�<��F�3_��Ż�-?6�!�:K*�Q1L��8� �X�T[�!�$��9�da(A͒	�����ғ3�!��	>�`�yT��9���1�*�?Z�!�$tth�Rh�$谅�o��!�D�p�
Ȩ �
_�KJ�hB��y�'sJ�B2��"c�8*W���`J	�'j�$�B�՘C��)��:����'��J5�(E��4�Frm �'���Q���:�Гj� ��4��'C�� ��I|&er�MX>l� )��'�4x 6��?���"�Ǐf&���'$"�:�D�R����5��:�'��u��1Q�u��K�4��M��'�� H�f�":t���$\	�*a*�'-C�aN�=���â-��\q�'���AF���؅ϙ6)S���'g���!
�[�`��U�&�\x�	�'�]zcN�2_�$�[u���3&����'p����Z8 B	[�J�0%�h��'Y�07�^<~Y���B�
$� m��'��iq#��֌Â��10p `�
�'M�$�UE����
B/E0r:1�
�'�X�c���T��6���l�]���� �L�@�?g2�D�"� �xi�a�g"O<��]7n�J���� ,2^�0�"O~�J6��^L���W� 'C���"Of-IP�K������*� Qj)x�"O�M����ht>�8"i�T1��a"O��Q�Ý��ř�
��?����"O Ie�[(���/��"��l)3')D� JӅQSw��{�+[�8�DE1D��h���l�(|�GD>N��͊�d,D��臂@�w���#�3W8��E+/D�����&j�HD�%څHr����J,D��c��'��ir�4y�`�25M=D�,qfN5�28�&LK:R@��&&=D���Il*$M#a�֚8f��d/D��3�M�(]�	-��z�4�D,D��@@�9Hܠx6l;*����E�4D�x)7EI�m�j�hǞ3n�:��2D��y0�[d4ܑ"��F�e�vx��'=D���WB��Q ��[�D^bzL�b:D�X;�^b��p'̓*��I�F3D���a�B�t��.<(��/D�h��	��f��)�f>
<0@�/D�T 5��/]��@P�/j-�!�R�2D�(�����s�8��s��o�1F>D���k��u��x�W�\7Iy�B�1D��iS�RWL�-Sgh��ہ�#D�pi���`�Tm\����,'D�,�ш��tW�m�g˰F��Uo/D��`q�?j�@t�J1E8���d-D�X��d����&-�@f����(D�4��+L�U$��7
@;�<	�)$D����&ؙ9�x4j5���i�LR��!D��YD)_Y��rfG8F�Tx
 �2D��
p���(3�a.\��볡>D�X�C���T�Q���6j��l��;D����f!:m�89E-^`�05�5D��R)]�H�h�D��1���&D���h�1��f�_�u	!�I%D���j��N~)�1���O����1�$D�dh��ū�F�Yfo�(pؤA6�7D�����22���� װ\c�L;D�p�/ .3���H�@&NQ��RJ9D����#�
6�n�K�F��Gd0��a-D�4B��/��m��L�x��\��#=D��cA�x`�t�dn�S�&<�G;D������}In4�4&�&N�\���;D���1���"`��h6Ö�Y(�*,7D�����j�r�AG��w
�I��?D�`�`]�t b4'�����A�=D�T�s�J�e�`"��Xrߺ�!��:D�8'�2{�n�a�fW�3�ˁ�<D��B���'4����`GڷJ:�PC� 'D�HС	I�k�H� �V�G�l�A��$D��n�#T��ą׎o�.�K�b	@�<��! �N�B�B�mE/Maf5�«Az�<	���z^�ꆧV���bЏ�x�<�E�Z
:,m�!��2�&����Jo�<qdo��*s2�S���v�<	�b%=�6����ܬ+J��$I�o�<�E�� ]"ֽ#�DI�A�<ARb��Sq:�0���"�`E��!Uz�<1��ǳ2�<8�G�@4l$��S��t�<���?�q�sh� �*IiƎZm�<��"�%�x�X��N�V?``��i�<� ��{Oé2G�Ÿt�=4A�H+!"Ol�Q�-[�t;�5�Q�J3)�Y�"O�U��$�dւ ���L�#$>�d"O$� �F ,t�j�+SmزF���1"O�|a%�Ɍ��,�Vp�x"O�Y�A��$n��9���W~s�!a�"O 
��G
c���4x��$�2��y"���O�ՁO�}�5�"�G��y�E�$6�����x���_��ya�>���	4��g�QA�B��y�
�]��p��& �ڐKAf�4�y"� �F]<Yz���q�P��-\�y��� 3���%�V��P��ϐ�y�!BY�l{��>^�uyOB��y�HT#1�$��/�pL��B�5�yB���d!���S1t�������y�!g��|Ia%� >Ԝe,���y��2W/��a���Au���t&��yb��6����;,
qz�I6�y!��N+���/�ʉ�$'���y2�K8c�P4xv�޾&7raT�V��y�l�fیQr�!�&J�\ )`�4�y���!z,�a�Z�7s�:1m��y2�ŁAa��0�OF f��pЭH��ybH�:*ڀ��7Κ�Y�(|�����y�e�+��������!2s	��y��[�!���2�pd�ɸ����y� 9&��j"iD�9U�D�1K=�yr"� `
e
c��{���k�!�yr�~>|m��� �d1�a�� �yk��a Ĺ�CJ�m"����5�yk݂rY̬�d&c��)��M��yBLN`������y�cr�J��yR�]�c�$!�&ʲR�h����y"DJW�x��Š�Q]q�s�%�y2.��N_�hd/P0}��T�b!P�y�@
H���qK��pX���y�oH�1�H�j�hBut�!QW����yb��!*����o�H$S�M��y��U�T�j�c͛o����K��yR#T�/����Ɯ'rem1$�F�y���g`�}����/ L"�J�;�y"��5 @  ��     �  �  ^  *  �4  �<  GE  �K  �Q  VX  �^  �d  k  ^q  �w  �}  *�  m�  ��  ��  7�  {�  ��  �  s�  ��  k�  ��  ��  9�  6�  y�  ��  ��  �  J �  Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�� |d��"O
`�(�;���8���-0��1%"Oj4��ND^[��"3/9�0|H�"OB���H��*�ʞRy=a"O�味V�!X��!&F�:J�$���"O,��a
���C�Ą�M�"O,$3%o�-���p���+Ն�:1"O��ݢ1����`���y14]2��i�<�6��{_���c�H�`�fX�$Kn�<��A̼VI�xR[�)�Ć�pඤ�ȓA5��('nߡ4�� �)˩%� ���,��r�؊b#`T�eT09���ȓ!�b��g��}�8�F��-? �ȓ
K|m�ș�VṔ���2�%�ȓ"R�X�j�4JN�1�˘X�i����̹	_�jZ��1!g��zܶ��ȓgil,*�J�
j�Ne��i�J%b���f	�(U��:���G��$Y^م�~r�� S�%T"���k\�jx�ȓ|4�1�îJb��@ӵ�ݩn�V��/[`�"�v4�R�!ʎ<��M�ȓ`:��z�ؚh�J�Z��$HY:	��H��p�m�C1��!��B:��0��EnjZA V;9����J[
2���	��4'J�EA�IVW&��~�(aZ��ӹ�>� o�Y�|�ȓ�f�A�
Ο7�H��M�$�����mޠP����/���ANXo*�ȓTv�����{ ��-7�*h��I��sB�8�8���3����ȓNe*M�悡;������X�o��!�ȓ'lj�#F�m�+R&;�|��2)n�C��0S4���T:
b���:�0!��e֊��)��ͷV��,�ȓ0�&�8#���� ع�L�����;�P�AFd���,w�6d��r�EQ�( �gVlɦ�M,H��,DP���|�I	$G#\���ȓ"�)���E�B	yt&B�^�LɅ�(�t2Q-�<Fsވ��C#E��U"O��Ӥ�.�ȗ" �d��"O�t���[&q�j��WbԱЎ$&"O�\�Λ
v����E�v��dKs�$�(O�'����7\0&(��#V��7�ą�o�y�we^�[��ѣ��)I��q�ȓL�b�2&\e<��DS�V�����<�P�Ѳf�bС�e3h٨��K[�<QU�zd|�:`�'Xݸ��$��V�'ǐ#~��D��i�F=���Z�X�ȜS�<�ѫ��uĢ(񄕩v��S��v�<i�芓b����C�;ȉb��Q~�<I�ϭ��1@���� ��@�~�<QeJ/=�t����΁ɗ,�C�<!�B����� �!x9V-�ڦՆ�T�B8���ʦ������d���ȓ"rbЁd �i�N�5,��0����$���C6�۬_Q�gA�h��1��	O��e�����1$�t���Z�  �e��>D�����Ay��(�$Y]@@x�<�q���OSt$����Pyձ���Zq���?9L<��C٤>�B�x�hNXS���U�C�v"B��?��_�2@8�Á�"�0�
�+��E"�T�v�>� <�)�j9�p���\d�b�K�"O�O
Q}�3�Gu�Fh"^�xb��T�7qO��DQ<�L�#	��]�����!���a�����Ν;��p��b��'�l@�ق��'��'��4q�}���j�!�4oȉ��Mk!�	�`QC���	�y��_UBlC��9mY:�*�M�G��E��C��9d����K9	>0�>�6�xjƀh���lYp���W�<��f�vT���~�°�B�^Q~2��(�O>�Y3e�:]>rE�~Φu��C,D�4Q#`�)i�4"����6d�*D����C�15�Ű6l�,09�Xv'5O"=�tk��l���Rdl!2�v��\�'�$����z
f��*z�с��D6��d̓Q��#~�@�i`���5AM�o���WBXA�<s��}�*j ɘ+'�\���b�@�<I�At��R�@E%G[�Չ�}�<�ի��Z�<P3vDT�]x*��c��x�<��/mo���@�M�!20$Mt�<�:ej"��f�Q}�T(gK�<y%/��X�FI��ѓ<>YI�A�I�<����}��hy�fƺs�8���
�J�<��"Y�qPPQ)0�J9�T��#G�<i�(oc��K@j	7SΚ��dE�M�<��եRX�2�V�fH<H����C�<5E�Cx������!�Xy&�Q|�<���	'yV��6
O)�\�z����xR��;�D	e�ԡ�tA�v�h��r1������	)�>i����!n���:f�(W��,9z�i���Z �\�ȓS4A�"$�R��.g
"���u�rjrf'�~�0ΐ�*D�D�ȓ���UDR����p�)ѡ&��u�ȓ�v(@BV�+<Y0×9��̄�'J�)���RDc'�8P�Dńȓ|��r*>{u@\�4��*Z�� �ȓHQn4�'��h�̴�C�/(�ԩ��Q��5���X6%�����T�z�0"On@��۠N��p�p<U�h�P"OF1��"�"���'(^�� "OH�s�o�dk�|#R;LI�"O����ߏOr�hrrB�8h�^Y��"O �
�� 4�PO�8�r�c"O���'kX�IW�4[Պ��D�(c"OZM� ��crl��g*Ϡo���B"O �*Ɩ�N�����E(@(��K�"Oƌ��EWx����*I&l�H�"O��bC,�(>p�o >1wZ5@"Oƥ�p��6k�<-� ��Nl�@Є"O��T	&86(�fnuz� �"OF@�qF�O0��g_qW�m��"O�ىs-C�x%��s�?+����"OY�0ԋ`
�|�U�Y��̜��"O8�q2�@v0��Z�lF/*�DLjt"O�� ,P9Y��Q ��M�\\��"O�@�P˜6Vxn�F�]=BK�E��"O�) ��CQa���:Ϡ��4"OȴjqX*��$��+Ǯ��1�Q"O1�&J��pA34��D�D؃p"O�U��!�)%�2M�Ъ�3Hc�3�"O�A�ˊ�Ԙ��o�8lt�0"O^��=���q��bo�u�6"O�,�C�.r�8��?{3z��v"OM�Ď��P:Mr��P3����"O� \�kF���@4Jq�E��"OB�qO� )g�}I�M_%(A�m#�"O��οs$t��)%ZD�f"OT����ĥ
�����oG�BB�0�"O�9����gG����1-�y�P"O"`�%E^�.R�l�rÍ<�My "O�p�
f����������QK�"O8l�5%�,u�Ӱ �D�2l��"O��l`�PDȓ ƆcT��B"O����8E����=�&Lj�"O.���;9ԼxRI��3���"O �canTs�q�L.j9��"O���N�e�*��g={����g"O&*�Y����0�O3����"O��Z��үo����!�	m�(=�S"O�]â*�f�J}��J��`��*1"O�:��׼�؄1��(\���{B"O8���,��B<��$�K/-��U��"O ��v� � �~(2����Plh=��"O�!΋"D����`�Yhr2"O�<���/W���
)��AC*OhT�PD�c��0lצ}jȓ�'�`@���\��HM}%6���'B�eC�C,Ša��+�P�@�'�����	jR4x�.�Uڀ�	�'t��O��'��kT@Y�G<<�+�'�������2x�d��4N�Ĳ�'�TEz���������A�	�LT�'I��K7��G'°�O
J����	�'�P����G�+)���R-?J���	�'^
	*#�B
/���Bc@_�4") 
�'����Ȉ^&8�k"��oG��I
�'i��q6��9�(p�P�c:X�	�'��mK�6<�<�n��]�䬚	�'��ıW��J�)��ƈ�]c�8�	�'��B�ˉ�A*�5�w@N6���'E�XJ�"M�t�cr�ɽ$�a(�'~D�2"�;i���Cުe��̩�'�q:.�	c�pA1�A�[	b5�	�'+�(��'�����#�V����	�'I�Yi��
�U��P;`	̹H�R=��'k�}(��O�PO��q�^>�@�	�'�2O�Z4���*75�E��'<����R�bP� Y�D�93�pA�'�N�jQ@�#n��!�H�;T� 2�'�(hY�Ȭ���;E!�f��<�'1z�ZՆ�78�a�L�8[��(��'�r��C��(��8
�@V/�X1�'yF����)��D���U�B�x�
�'B�Y�C�C�g�h��&�U�A?�\S	�' �,P�OT�o0��3=��A	�'̊`��K�j�a�.��<p$	1	�'�U�g�6Bp�E^�:�x|z�'8�Z��d�
�R�2�����'�4��%A�J�2EI4kO�(��tY�'0��S5J�g+�R �vxؠ2�':8�����A(z��G��u��`�'��R��Dml�s�G�5)~� �'��`��&9�=Zǉëf��Z�'���H�;}��b��_4y�
���'ˀe"3-�?G�J%��n��D_.y��'>\��� f�,�,�1�4��'tʕ*IK�H��)���Ǎ%Cf��'�����F:݄uR�(Ϲ��L���� 򩰳��.��ۇ�І0���%"O&�S͏:a}�0�B��&I��'O tk�N��'��@�Nܮ-�n���'��t�&R
ZEZ��O�x�(I�'�(�ڒ��0^���e�>w�t�����?A���?9���?)���?��?���".p%�#͍(Y2 �b�V�t�����?����?Y��?����?��?��'���eN��1��e��O>d��@���?����?���?���?i���?Q�Tm8�	��<T\Y��ȳu�@����?A��?9��?i���?����?�=�pQ���4i"ڜ��N8^k������?!��?����?	��?A���?ͻqIxi9A��$��6�O�	��=�$�':��')��'��' B�'���'4�e��G�<�F�"���-�&�'A��';�'5B�'�b�'���'O��p�(�[�b�q��\9��
��'���'1��'Lb�'���'��'����q�ґR�	��;T36!�6�'��'$b�'���'��'9��'����ԴY}T���?q5$���'��'
�'��'kr�'?��'˪���*���C1�<,�"EH�'�"�'���'Gr�'�R�'���'�����C�!���ծL���ڣ�'!�'��'}B�'���'��'/��m�uϲH�c�kD�I��'�"�'C��'ib�'qrHm�V���O��bL�Q�\ȳ%	zT��	Q��ş��������ܦ�� � %�a���X�56�yq�bQ����Nq���4��M3Z�4�cH�М��%V�Z�f�iV�iMB.�)��z�'�"Đ�8L��b�������`�[����JVA����_u1OT���<����I�(Xظ���@�g��BU��!fq�n�c�<�Zӹ�yGǏ�I#�Eb����B��[�g��3��6m���̓���i���D�<O�xZ���AD��"$�#nĄxu5O���d�.Gz�)jDl(��|��5u���Ey�(�	u�E�Xu�qϓ��4�dS֦	K��-�	�UE ����2Kx�������@�H��?��Y���ܴ��V3O2�:l\yZ�Bحo*��9e.�=(OE�'�T�K�;s@�L����II9OF��Q�'4� �	�,��U��m�&B���QS���'���9O:��r�K��1;si��1O��l�`$��(0��4�*�9��̌"��d��b]#TF� �r>ON�lZ"�M���Gx`�t�@{~B��$ �X�4i��%?����)]�S���i�m�'��`��U G�6˓2f��#�.�3�dW��]�e���
�B�qZ!�$�e��[S�G#]�Hes����{d��6o�>2u^|Je	V3]"�Y��8j�^\CdêN��34���o\�8÷L8C��"�.'|XR�	�t}<q��2=xQ�1C��*�����F"w\@�� �,�H���`EL����-V6fy�dǫ1��E��^T��D�|0�DCpdE�:盖�'���'|�Ԉ<?�V�S�׈1J��B�+�ȈRg�צu�I�dHg� ؟�%��Y�IZ�K�f��#�2L�۱C*H�F��}>z6�Ot�d�O��ɘO�I�DRFˊ�?��\��/W93�&,�ҫЃ�M�E��?O>E�4�'����cB�0���v��Dh�i9�Lx�B�D�Oj��y�n'���I矜��z>���mS�J��Y��-H���'��'1b�"�U�h���|�	Q?a%��,~�ᓊ]^&4`�����	�j�LQ�'�\�'�?��y�^�X�Rq�Bኰ0�t'fM�	�n�R6�8Pd_G~b�'���'c��'�"�IËҚH�I��F;w!�$3��8�q-O�˓�?�M>��?�/*h�
� K?3d���O^�t�Na{�.Q~"�'��'�r�'���1��'.��dC�o�, ��,�VSCEEmӒ�$�OT�d(��OV��L�VU�׷i�^��5j��e���� ,��N0&��O���O��$�OR��ɼt��'�?a嫟�4O"<8�'I`ruI�z5���'7�'���'�¬y���ē({�l8D���䡛����f)n�ݟ���|y��H>:�0�Z�D���l`�i��&c��[N�[ ��[�G�����	�^��#<�OQ�h���F���"k��lg@�I۴�?)�_\^����?�*O����<��:����Q� E�)�`����oZ��8��S��i�-?�)���4F�U���
��p*�$u[x6m�.�h���Ov���O^�ɤ<�)���!�%�8L�xR`�-C|b�86�HȦ���g��0�c�"|z�x�L���( !%�<��ĩ�	�� �iY�T��)��Qğ`��Ry��'�$9崜Ȁ)K7I+(p`�J,�l�<��ڟS��O�R�'����;�ڌS�EY�s�xT��$$6��O��ȅ�o������	H�i�qc�I�$�6�{v�Փ ����fa�(�� �&���?Y���?!-O����6yA^t��E4R\laV� Rp����<���?��S��'a�IrӪ���	��.𜤪T�˭~���[��"b���?i��?�*OF�b ��|Za�D6c[p��q�� [���h�a}��'���'��Ο��I#.
��t���.=B.N��������'���­1'9�G� &t�R�`�.�z���\ ���]=�
�rGH��:��p*83��?�Dz�0i4u��d������qb�)siʻ�U�5.]U�hQ�ğ$�����ܴ���a���Z1z�JO��Q�U�'̄pj�b�1�,T*��U�V R��
� �Q�O$� N���X�\D
Â��rc�Y!nǫ&�<-��K	8^�Q��aN)��H�q� n���`2��Ov��O֕���ҝT
�ñ�Z�\$���i�(O���9�c�%�`������'���?��/O :]H����w+�8SD��nM�b�c?�S�$ܐ"���'^��B�MӴe�����S��,)���]-4�I(���O�5��]<qxڱ;R*|٫��ϧ�y���BʘXZ��	|wư�K �O�TFz�O�bc�ꂇe8��E��#x5��RP�'����ckT���';�'J�~�;}���"�!I�p�pE�!�X��6��ŃE�+J�}9��'�R�Z�`�M���H��^ �����1y�U�DHQS��iA��7��T��}�'q�B���;V�Xa⍑`���0S�'�N�À�'���,O����<�D�_	�x�Xs��t%�vM��PI!��6?�R�+�
	/c"�B#m*q_ΔDzb�O(�R�H�����M!�]%#��d�jH*�:�C�ℕ�?����?a���lQ���?�O��u���"Ԙu��D�+*���T�.6Pi�4�X<29�����'q�ق7IU�_ԀH���hC`"���0�dL���fY6x�E�'�lL3���?��
�C�db�OE6fTMi��[�<�B�"s�,�,�����S�<���oL]���T"T �CI��<��i��'��R6-r�$���O�ʧI��1���3):by���~�P;�R��?���?a��O��`����ШC"q���M��Ԛq�ߋ)��DN
b�&i�(B[���Dyb�ԑc�):GL�T�f�L`�x9��֢B�U
@���6��s  �r�Ey�כ�?Iw�i<��'
�S�}��A��ؔ:9��
�?����	џ0��ß0�i>�E{�㒗-x�L2�MQ��V��Q(��0>�A�xb���H/����a�2���+P1�y��)�J7m�O�d�|*��3�?��?q�C�]�p=0c�M~�U�*T|������W�(��S�H�*��b>�$V=V���	h�.L����)ARb�:��ľWN���N�.�)��$�R�Ƞ,.q�G�6Y&\��H�(ь�	���S��?�C��|64��c�O�0\�85`�O�<ɶI�
��a��Ж'Z��,Ps�'�|"=�'�?)@�	1vN��3K+S�8�!���?���:���4ȝ�?y��?���U����O�я!�8(�Ϟ�H�E-;��M�ٴF� In�	J����PIrF{BD��N���e#'�Ib��]s%l��Wf��n8ưq ��?V����O0V�<y�FK8q������(k٪`j��h?!D�����7}�d cD�Kؼ�a�#n\�ȓ:�:�0u�]�p�kSM!��Qd�i>�&��JbD�M��FA�q��P��4]+��q�/5�?����?Q�)=e���?i�Ol$4��#\�k
TLY �'Z�ŀ�B'	[~y���]Qr�qa#5,O8@�aiW�*�(T!["�B���G$J�I+r�8�T�⭙qX�D�Vd�OءnZ� 3v��ԯ,E.*!��5o�zB䉊_�����E�r?:�cB��d�B��7�N\�&N�d5,�G�l~ �	��M�L>�q�W2"�&�'��U>�s�B3f�x���*���|�P�ᑹa�6������I�l�	:��8@��-��l�,Ħ]���	9uΚ��$(I�@9����	5=�̍H6�ޗ,���H'�L1;��K��Հj�,��;?�Z�!p(��#�b��+ߜ{�61s@K ��G�^�r�y����K?��	.n��q1gJ�'�8J�S�Ya��[�ԟ�F��w�p5*�����Kűu���	�s;���{Ӟ��ÄJC���b�W�`���em˼undl�.B��4�?I���?���6cZ�3���?�������C�b~p4�f_�����	\J~Xbu�K�Ck4���F�)��q������M�\��iZ�J�A�`���x� X��<Q�̰�*[%=�а����e� �S�-/��;�T13C�ˎ9�)Zt�W�K(X�����i)R�<��X��?i��9UC�ՈD`97�=b�'��<����䓬?a����O�D9B�/�(�l8��0= h�+�y"�'+�7�R��'�����?eZ�E��L!Z�c@M� g�z�q�*D����ɢ^���R��ݟl����l����u��'��ɗ;]�Ä��c�F���*ո�~2|¼�e��v�����v�\����U�31:�r#�S>(@S%L
���;"�޷^��3�w��l�eQ*Mb�WoT�x7���.�Ry�I��=Y�鄺C����ޡ� �;q,�k�<����m/>a�G*�%r�v  �L�aQ���v�I�o���xݴ:	
U2`�-~dP�҅��d\�i����?���?��iԅ�?Y�����웈H��݈�T0^@�����}",Wl��.vE�v���@����� JBr�9�W�f��y"�K]��.�j�$��)�0Sv�Q�I��*��G��ʃ�?���i��E4�ä4�����- -��
�'�.�`r曟K��!(�ѐp�&Hz
�'��q�A��i�* z�CH�B�;�'�z7-4�đ���n��X�	I�� `� $P��2��1~jp�ֈ�4����O����&]��9�ԭi'41�[��Ȓ�O�ڝ��'lp�]�BN�6j`�����>��!����;|5V�(��B ��3+�#=�6��2�I˦ęW	�1�&��'�x�O(��g�'�z"}
rΟ��VU�g$�ysh!&��R�<�w)�`,DM�aa� 6&�H��U~2�i>MO<qWN��`�x�C�b�+�N@���<Y��. .���'8�\>�s)_֟t���<i�ɟ<N!�Y4�W�K�r�r�ėO� U��&�s��q�/O�SZ�矄aУРFdf(0��ʊ~� u(�kM/T֑k�B�5ib8�,O?�$E�D�N��#'�*$Ai�3���lAR�Z��O��nZ����O3>��ĉf��xPC��%���90�W�\���O�����9�4p��!e� �ca�D��1O��[�'>���'V��g�̦t�е�5c��o�~Jt�'#B�Ηw��V�'bb�'��Cb�y�	ڟ��d�ݷj���MLpn����H�t��/I�4��	� ,TI��K�0I�$�V����Eծh�:�i`���VO(�J�J�?��� ��;b�������5p��XC����I�"�$?|O̴��V��q���jr�"O�5�	�~ [$��8@���' �L���Ĕ|2	4��7�Ohf�s�/G
Uj��e������O����O�uZs��OL��c>��rcU�%�,��G"��2C��Ѣ�=V[ġX���x�l����R$��4�0 1bH@�P�#� ���7X~i��D�3����pA�`D{�A��?���i�����
^�	^��i��t�rp�	�''R����$qn�hy�-Sl�0l�	�'/(�J��M��y3��[�-D�h�'c076�D׷.�dn����H��KD!0�.�2bZ�q�"�F�7��ek��')"�'��`�\�&��S�DV
E�����@�U�׀t��e�T���;q&@2��m�'��l�V�CϊE�G%׫&�{�.�-m x�A�mL�N.���cP�i��ѕb֧�O\����'I^"}���N�Mpd�w�/[r�QY��O�<�M
�ʸ�4�F6r_���āN�l M<�3�K�H��D���`�}(����<�񈛸/����'+RU>��G��<��ğ���'z+��Pwa��	��9�!D;���J�S�����-K3��$f��+�Z��R�<�S��?����53���0�l�e�t�Xe�Y\RY��Ϙ���r��Q�Ys�	�- �(�	��y¡B[(�H�Ĥc�r\Q��M�O�AFz�ORO�'�PQ��J	ȝ��#��`��'FLM��Ď^8��'�b�'���̟�/^�F�eT��@2u�	2iN��ʘ� ?��[!nN�dUT�P��?�EzRk�;)k8�PV��:���%d��Q�F�q��cc�p�LeB
��Oې��@��]�<��'SL�k7/U JDi��	�NF��'�
P�uMa{"	�!-����!:5眡��%լ�x��'_�E#�mO�r����5?X��1�!��|�N>I3��+�&4��)�ph�w��ً��Һ@j��'���'Ф�b�'�:�e�@K�6V��sCHR�K-+���D�<�i�I��A�ʽ�%�]�{r�IG힇�(O`�y�O��Q�=�s��!Ӣ�(X"�qQ�P6�$1FD�L������(O�) �'�&6-�/x���T;V!�y2Ueɩ6a!�ߥ.��!`�%�^����։GY!�������'	�2�D3c�Sp>�$�Ѧ!%��Fm_��M���?�-����&��!�Hhp2b��$	�0��C
�OgT���O��D�2,Tl��ebڳ!���Iad� e���O��9�Qǎ�+{����̉7%�*����DJ�.�� <���aP�"�8�ZA���d�JOUrd�+��'�H
!����i˺�����I?�H��l� �N:���P#�>x,��"O���g��DP$E`�9���$��D{�O�0Op�y�#Y8]N�l
e/�;&�Qc#=O�4������l�OV���'�'���'T����U�?/T���)��omD�aFD 5)$X� DJ�ؙզ�O�K��(z�+N�0���f��j��py�×"t�:ds�U�zD���4�~x�l[�d	���U�k����,�"�R���h�RIR����'^`�O?��5b\�q#��~C��3�`Ôy�!�$� D%�� Uƶ�'�P6+q1O���I�����	n.��Va��.�1�oJ�f��d�O@�$�=���D�O"�d�O4�;�?ͻ'�|e�Wm�4^*�{G�T;3ʄ�y��'�B�ꦧ֭KAJ5[�jGF{�ˇ`P X��E؆pڑ�$V3Ab�	�CF�:K�� u	�e)�C�B&���'�N,2T].$g��K�茜";^��6�'��B��'J�6����<Y���F$��D(�G�!-*�1�È�>�!�!�qӲ�[�,��Bc�=���Gz��O��U�@�Bgء�MRW�pn� 2r枻|D$y���)�?����?I��`���Z��?�O��)�ꅰ �E� �Q��(F���IK���4q�`���'�t`��>Bt ����G=!�"e��o5|�*8��f(MߢD�^��0<�������4jڄљ���%OV׍Z�vў��2��hqq�
?.�x��¢9A���ȓz�(�ɂ��A��ڠcL.9 %�Sg�&�)§kJ���/D:Yo|�z��Ӆ{�fP�ȓt����dkZ~��QBQ���?p�i��)� �s���)%��Rf�<RfH��}r ��	@�.B&���'P�B�N-�ȓp��%���hcr�f(�ךa��[�2MpPa����c���C�J!�ȓZ�!P�
�$M,T�&D�� �\u��It�ؒ�Z�A$5Hq��$��ȓR �E���^�S(6�SF�^w�ȓ
��5"w��%�u�$�\L��]��FFm���-x�4�d��r�<9@�R�c=H,;B8=�R, ag�o�<�V
:9>]��$�}���â�i�<��/_�[��@oۼ����c�e�<���T9nt�m	6'�2���f�L�<�f�ޓ/,bt`E
��$`���t�<�EK�/�Ic����	|.�*3f�Y�<	s�ם׾�ҥ�T$q�� �0�X@�<�� �8i���Fm����S�)Oe�<A%N^�f��5!�'Y�f��!���I�<I6�C�G�H��O�B�}��n�F�<ig�˰g�DP��Q�ڐ���V�<Y��ڙ��p{��B8J֢QH��X�<i0_�t�V�3(�77�:�e�V�<�� z��z�@�fÆ�x ��T�<�3A�?{�٣�D&�����H�x�<��O��x3��́ab ��r�<1��0���b�H5VѻF#�U�<��aS37ܺH�ue�d�D��P�N�<�p�����t@O�	l��DN�<I2���B���@��^�p��1 �_�<y'MW�_
���[��и'KFS�����$�;2d4{#u�⒂Iܐ �m^�\��͘0.B�(r��$��ꏧ7⑚Y|
��b������A�D�$\����1�:~��p��#KQ�X��W8P�TB�U�xp��
q�m@��4xp	S�'m0 �r��&Tl�!�g}"O�Y�N�˷�D$P2�"�f��yB�����ز�Z��0��	�M�'F Y۶��G�#_f`:Ǔ���z���`y@� xi�ن�	Oh < '��D3�*�e_,�[�ɛTiJ�Ē�P(R͆�qN,EÔJ��m1���ьڔ}���>�2m�u�8�C
U~�����T��*QIf$:��Д�> 7kB3�yr�_'5bՁ���2�6.F7*��tP�)F=8jp��"��t���Y���E�>��#��Ĥ:	V�R�8D�
��D=uc��E.Q�	�"�R�u�0���f��}7�$4�M�a�j��њ{�ޙ����E���D�N�h�џ�xcfÇ_�챓*�{���h���x��GD�$��-�`�pvN��sO`�rIG/:`DT��'�(g�.��X��'�R}�D8�p��8�B�������>��R�ٟL.��Xr�K����B70D�`! �ȕV7K-Kb�,;r=���P�Z��倦��@I�^�q���OXT��J�0�� Pp�?;u�t�'��ħŚ�-ɒɉx�p0c1��m���uHϲli����V�L����'&�ْ�,�s7���t�^]0\�)O��r��Á�xt�t��)+6�=���	�r+6Xig�V�94���#�K6H7mu��H�(�&~�r�	e��h(�OP�ha ���cM<g"\�"g��~����O��aL<�&���6D�������2� �/Bz�(eK$|O
�ϻ6�fH�.8�:}
BG�?-���?��3�I@?�B��YRʙc�.$~(e�΁�Ktvm�W�I8�p �G!S�4�l]��c۟
eL7m��+�Jų�,�FN\2�'0a�&	�=ё���\�R"��&�`4p��9}ـ�S�? �1#�_�=h%I�%�z��);�W��D#Yo�ԱpF�Ɍ��ӧ8���cQ���m�&��Oż]Bb%�"��V�=Ƹ���CWY
��� !\ti"'�Lq�D�FbߊZg�	�M�2�ӓ�����3LY��"�РQ����b͛(]�8���/��=!ԍ�#lV���Ē'�tDӣ�4;9l[��	e�'�>m&��e�ȊW+��RVN�VvD���e�nܰ��D�"��O�ȞP_��Xƅ�> Y ����	���C���!;�@��>y���.~���"�"�h��D�7z� ���=N�pX"�'faa�̎�q�����Y�	ɼP��O��N�_H:MJ�ҟ@3��hb��)�6�
���f�
�&���2$Р-è�����*1h�G�	A�Q��9C=����T6L"<q��\�s� ��7�П�p=)U�)(sPusբ)�R�(a�2<��*3M7�Z���Ɋr3�ur7&�tp0iT1a�Z	BwK��O����A�R�	��N��1��Y�88�h`a�1(��\zT�Xq�v�D~�P#K��@;��
Dʉ���W<�M����Z`��#֘]�H�ap�Gk}�U)�F��G��~Z�[g�@D��ēc�$�1���O8����T�����D�)�f�z@W�(��F�W�M0��#z�I�G7�T�T��b�N�7�cs%��f��BK�m&�z�IQ	V��:gJ�qT�>.L�X�P��q�T�44�c�B�4 `�E��_�Q��I��xrcD2t��W&�"_l�ҧRn�F%qeL�K����w��\Ae���X��x�qQ�;n�B�r�M�'��E�s�P an^*�@�"f!�x �c�#�3s�Q� �K$�M�w��n�={�t��]Z��|0���� �ӏ�d���ޡ�EC��Of���f����aC���@v޽�h]�OS����¼<y�G�5�>L;��K+3��Qbe/�}�'�0僤��p�P��ѮU)D���۴�yF�~�ڴ&��6��`D~@��K\��0B��[����a	:���1��H�OUN�Р$��nC��)�~Y�1���'��Z�J�!
=!�D�+(&|��Q��\����O0G��fJЗh���M�:�;N|������*BBr3 �O�ш0�售1К��J���u/��k ȉxv-@)�pd�bk�w������'W���W&k6f��^i�&m� �h^�bu(	�MYџ���M�$�xzQ�Łd�6d��Nʊ[�P�B��Z�)`�n�k=^ȹ�O�E�dP0�tU "��|'Z�9�"OBXá�˙37��`�z ��"Opt�7���h\����E�>�D��"O� ��f[�H�8�"�E�,$�G"O�A������%*e�ܨ$��1"O���6g��lˁ�O�x�4y�"Op�J�G!�(���D30�r'"OZP;��݊l�KE�Uu>��ѯZ��y�[�'�����N�Gf���Q��y�m�R�(��"��;�p�Bi���yR�D�x:\Y�%�]�A@����(@��y2&�	o��Z�[848�́�K߳�yb��99��l���C�Z���j	��y"�Q&r]N�x���7�PAt���y�C�0�,%��̧%����c�W��yR��"�QY����r�x�`*B��y�ȑ�*�J	��E!Bߠ��b�Ѳ�y��. �]K���:L�\"��ɀ�yR'W���(�竖�E,�JՄ��y�"
)3YX5�W�:��q �a-�y��!;��4;�ML�0�����F��y�O�	P~�;�nY�%�J��c��5�y���7Oʰ;��"J���%���y�@�� unm��a�wư<rRgѥ�yb ,6x�����9Fc��a����y�B�S(��f�'b���A�y�ᐇr�0��`o�,���~W؆�O%XH��ئV�wj�P�x�ȓ6o�h�Ӎ�&�Y�s�ܕN�D �ȓ�L�rd��i�|�Q��|����p�t���Y6�u�t�� "�Ԇ�Ɯ�Q.�v�����Z�r0�ȓ]}�EzF�29+|��!�
�)FV��ȓK�r�PD̾ZF�� ����,��S�? ���!�G�TK��Z$>�����"Opx��;�Q+G;t�xj2"O�"/��6��[�Z�|�$i�"O�hQ X�� 	4�U����S"O���҈�}��9�8����"OP<y�@Q�(r�e�hM�\Aa"Ot!�w�T���I:ue�.F�	�"OTa�Gc#z�8��#��w(�b�"O�Dx���.o�8���,�%D��0�"O�P8'��#��Y���c�Hl�"Oh��N0s͂�#/�;�ސ�"O�͙�+I�j$��1]n&~�:�"O ���0WC@y8ǆ�	|���W"O���b�/a�(��V�3lC�ݱA"O�@s�Z3Z~Y+�D
�&��d�"O^�bN͠C��S#�۩o&��c@"O��2c��vG���i�3$$��v"O�Er2)��	�m0��7e��"O���ޝL~�"3�Ĝ(�nE�$"O�l�QO�k
�h�o#���s�"O�	����x%�P��Y���c"Ol)� 	 #�q��>S�T��""Ol,��Ѹs��\2��ʃa�4d�w"O ��ᩄ2{摻�Q+B�
t��"Ot�0iVF�l����F� �����"O���l�%r��T\I�4ڄ#�|�<i���.ވ�B����I�FS�<Y��;��q�p�N8#�u��D�<�aKV�NR}Y7@����(�k�I�<��c�g���X5��z��ث�(�Y�<9�ãf�DD���Y�P >�����Q�<�Fɗ�=�
R��fUJ�<AG$Z.Ժ�*C��Y�˓1�pB�I1b�q[�FаL��tI�fO�{ �B�	a ��!���8
Ij�8e�9ZLC�	�r�;��N�1�n���� m4C�X�Z횠J@���pL��(C�	gD4]����W�d!�kަU��B�	�
,vu:AL��[�JX��*[g�B�	�v���2o���q��i3a�B䉑����� �@m�5�Fh�,�B�I?a\ �P���j(��#�V�3)�B䉫*�5 `Q>+�����Ӌ`�*B䉦>	fA�RP�bҮ�!e`,4O�C�ɔs�,���4E�p���׸��C�	z>�j"FP08�BI�;V9�B�	��R���hZ*V�>��"��d��C�	��.ݠGbC�GXލX�F�7�C�~�ZD �[I¥� ��/�LB䉳�D�����u�"�	mB�2J*�<���3���s�
�3âB�	f�FA`0����=�E�k6�C�, �8	cGC��1$/]�a�B�YF���Í��H�a�EY���B�I:u�W��-&�-�4���BdnB䉭F	���&�%6�:0ʱkK:9�^B�	�R�r+O��T$s�-�6M,�B�	Hk��X�
�&Q�.V�;Ӷt��"O�Q� F���®��s�D%�"OT�����+�N����%$��Tr�"O���Z�����ˀ je!�"O\��EA�.����H2o�\�X�"O�d��	�L����F�;_���hG"O�e���]7P�r8�c(� pި��"O� ڜk�N	��0-H�g�'Fb�x��"OhIH��N)_�5c"��Fٚ0"O29H�ߎDS��5��ܔ�yB"O��Ӭ�-b
R�`�ڌ!�xIX�"O�5�/[ {6|�SR��o���g"O��R��!?��%�W���O�耰!"O��CAcT(;�^`ӆ�Lkִ��"O@����އb�t���
S�\X�"OvE���S�l〼�K
�+S�8�4"O��kW� a� �LʈM�q"O: c� -�����6�4�a"ONȠ�CƦP��5�$
ə(�=�"O���d�1~��M��i�4?�`x"OfXB�%H4t�=�"��I�r�+�"OV�x�M?BiΕ
b �R�N���"O$$��Ä�EX����
�HS"On�����4n?l0ɢ.��bjB	b"O0Yd�S;W��љ��&�T���"O��[G���"$�*��E�o �:�"O&eCȋ�z$��)�(wd<�C"OZAR2H\�g}(�P�_�PTb���"O���;�����EhP�F"O8PȔfܔ��0�A�{���C!"O��Jڙa;N���qqD��B"OƘp��'.����Y�b��P"Oz-�EaÄi^���/6����"OhM{ׯ���vhP�%V^REK"O��C�F!Y�J�:+"`��"O�����,�� �$˭u��H�s"O�XZ��^��%R�d�z��Tʁ"O�%z��$i���a�ˡ*���d"O���ɜ�f��勴�H�ww-R!"O�u���,q�� �.?�9R&�E�<�!"��(�,ȫ2�i&�D�<�r�43�����FW=$:n��n�J�<q�͗�@w2le��=H� ��FD�<���Hq�J��^ZRf�ӓ�@�<�uON5p���j���'T�p����|�<Yc#����Ag!V�PQ9�M�O�<yG�*:�<dY����2N<��J�C�<��'Ɗ�<�Z��ݽ	�2�� �Y�<�7�����xt�Z�?�\����Z�<1��C59%����	�A-����KTY�<)�G���z'BU{�����JZ�<����%e��!5пG���ZU�Qٟ�E{��I��9}�ɉ��01��Ś"�%(k�B�I�Y>8�h�@J00��qq�I-�rb���뉇zP���p��C~,��3�I�6/�B�I
wQ��så*a�]w�79��B�I,x�1��֙/�d�P��@Z�DB�$| ����G:	�24EȞ;WE�B�I"-t�l���[Q����BJ�o#��'�ў�?�צWZ��#�=p3�x�
)D�p�wn��ƹ[Ue�4,���V�:D������N�C���$JĆ�ZPb9D��R"�˻R����S�B�h�"#7D�@4 ˯A��Tm�,�J�yQl3D��"����]�ǨM:ZFBͫ�/D�0bBF	V�Di���آj�^��6:D��z'JؑZ�t� &#��A*�<�$�9D��K`�Uшh�%a�3 �� �2D��@ X�@�X�`��<I ABa�*�OT扱Y��p��A�g�Zi��;��B�	������K�[_Z���O���B�)� X�;���PV���ՊU�%;*��#"OP��SO��) į&X𕛠"O��8��R0����ݿ:e���"O��C�4�Va�D�ƙGE�k��Oh��� i�A� GY�ւTxWB̔�Q��D{*�
p�������U1�.��6	��cU"O��'	]TZ�R��T�T�(�WY�@�<!�'|���ቀ�a�:�S�c�$gvt�ȓ4,�e�,B���v��,r�$�I.^�1Of�E��O��H���6Zt���7hP�GpM�'�'R�'��`$�K�Z���	�Ŋ�]Ƽ4K*O�����73�9�&�a���)�!�a~BZ��+�i����,�F�:��0�w�9D�,�b
Ҥ��L4g��Y����9��M���i��T�J���O4�$k�lGx�!� �y宙ɂ���3��UӲ*W.��=E��'���G�F�;&޸;�7S��Lj�'"�p���J+d~>M��*QF$I�'������(�Rm��M֌<v�(Q�'�l�(��C-O&4��N0�ҩ�ʓId�iR��|��dK��j�~��=A����KB�]x��`X4Ok&������y��j�����I�-��GA�O�	��HO�NTh��ǵN`��(Æ�
5!�D�b�����3ri@�`��ϖ^"�f
O �{�eC�8��q�K=k�);d"O~p2϶tɴ�C����Y�4�Å"On�IхC��� ��EF����"Ohm�O��0���s��Y�}c�\��"O ��r/Σ.��1�N�a��x�"O�I�@ƍ�0��J��R�dD� �w"O<H�&�ӂ:�!2dn�7c0�<�"Of́¯��q�R��4DߋqL]��"O p O�3��L�Zh�A��V!��#5B�zre�.��%�G�*!��$m��s�
�b��(���?$$!��� ~|�� ��@(�V4����!��F�h��UH���."p��QNθ`�!�D߯B�d<�W��
.���Q�ٕA�!��ݧg͊4���F�0x� &�(f�!�Z���(��]u�$��dJK�!򄗟m`e� ��Lah�
W5/�!��fc�D�Q��
~T�	�i_�-�!���pd��L�'0��aQO�Q!�dQ�.�]�r䂘6&��U�,�!���Z(�Ҥ�(@�SJIC!�D&W�PY���>�!��˃ T!���|C!1��A+85�F��$.!�ٯ����g�9Z�́R�[=+!���#")���˄
�r�SK��!�0b�� q#������'�N6�!��L.-�|�"�߶ �XT�f㜪-�!�ҟ�+��ԍ|�8!�E� �!��e���	C,	vYԚ�@�g?!�$sep3B��8/���S��oB&h�ȓ06�H�b��IP�����7y�L�ȓt�إY���1��D����4I�2��ȓȾM��@,f�Z�b	ҋ�<���-��0��"�̘sW�.�y�ȓ �*4p+�Q�M3Ձ�����"<Z���ݰd}�`[�N�nq��ȓ] 4	�G�c뀡
5C_�I,�0�ȓ<�� ���	��oZ�Y�x�ȓ�x@1�-ϰ{� ���K9:��݆�S�? >�3��LM����!��#>w�tb"O�`�w��
�k��A�@��4�!"O|2�l��r-���՛M�R�"O����a�mBD�Gԇ�L���"Oi	�ЙX3Ȕ�A�5r��R�"O���f�������R���Z�"O�i��V+!���PMނ�����"OƤjѪ/|:]�Aϖ ]y�C"O@�ٓ�[<���qD�X?F�=�"OA&�ږ*J�u��*Ӻ_C��2"O��iC(;�h���\�D�"O��j3E�����D�Tz�"Orȉ�a��P���'�V� ��0+�"O�0��R8{ޞ�y��)kμ� �"O�@Z2F�c>��؇@�6�<��W"O�ͫ��� @k���!A�<p�"OB K��I�[��%��Đ�"O  �����X$[`k ����"O���r��7����	G�`���@2"Ot�YV�Ǹc6,�H�G_87��铔"Oڡ�աCng�q��e
	|�H��"O�ݚ��7�8��$�8C�=�E"O�0�g��.G��+�	��`unEhd"O�Xٓn��;(�=S���c����"O�쉒�����g��VG>Hy"Or0��ΠdiP��iS�UF~ŉ4"O2a����@~ Tb׈�:e��l�"O��15�8"�&�&%�{��� "O�y��Y+N@^<����_`���d"OnXi��/�<x��zp�T�`"OV}8�.��H�l�Cħ${j��K�"O��r�(Ҿ!
Yc��ɣ2�v�C"O�p�򀒼+G��r�	�*����"OʼɒjC�T<�cfM�
а4"Oh,AU�ވ~���HL�p�Lq�"O�����~�0���Y�,b�%h�"O`ӰO�I�&���N�ZT�Q"Oz�+#�[�I\@�#'.�.4L%"ODM�r�H�*�� S��y�%B�"O^�z��_�_�h�5�l.�9�"Ov9
�Sk�4� 
��@۴�k"O�Qh� �V�xb&��ȥ	�"O�����Z�W]R�� 2�b��"On��. {��	�0��Aa	�'�n4Am��%^F� � �*-!��'�ia�K|�EkA�^&+{�*�'��Pe'�kل)� k�(���''F;5k˞}�`�!3��$��I��'�Щ�Y'j���A F=j=~���'\���`HȍC����A)4x���'�>00�J�7>]B���!+[D���'L:q;3΀�K� �f�A��ޑ�
�'>�,�ƣ9J�\T��G�6B���'�\����^�8c �Jf�
�{�Z� �'3��a�.ǂg9$h��ʣ+S�͹�'=ĉʃ'�P��	&�*03�'����#I&r���0W�L4O�X��'�D(��5y� I�g�ŷ-����'7��9Q��)^R|����$c&|�	�'|�`IB�#�.���.��
��q�'��Dr@�����4��0l8"�'��	c��-	���J�2R���'�"q�!����tIé,&&\���'��� �#(�e�S������ ��"�A�Fo��cd��r"O6;��[*~��upWdL��(m�"O�e� �U����sa�7*�~A�`"O&t� �$B�i�&`ߦZ�t�r�"O�9�JJ8���N̏K_�X
�"O�#�&��U�&]��P�xjL�C"O�����W
�w�J4Xtƅ��"O����?rn~��5��22e�a��"O��A"��!�~�BF��X�>��"O��)q��5fVlT��-�9J�4�k�"O�͙���"(�\���+��}��"O4i8�߮f� �@˄�^�d��"O�@"f�&$f���SZ��9�a"Oz����Q$[�7o�f�� "O�P�e�+7E< �F�
=Z��9��"O��E[ێ�K#H�v~�]�"OT�Ō� dD�|b�gr|3`"O�9�#EG�%�hUi�׊2&��'��A��
A� �8PI�h�)-���'Y��B�,P5 �j�j�L��O����'<���D� Fj��F��
G�0 
�'ǆ��LD�r����D���B�N��
�'p�l������
��2�J��
�'$Z�3��c��0J��]�`i�	
�'	�X9���V}�h���(�N�z	�'��t�E��=-�V%�%��ŀ�'=�\0D F�!�1�_+g���P	�'&͋�/����f���		�'���	S"� �(��=LZq�ȓpF��C��-HZ����Z�(�hU�ȓW̨��"L�Pndh�Q�[��z܇ȓy��!a�	U>Q@�mPW\�=�d��_�̣1}�@`�ɞ��&��ȓIX �#��<ǌD@���{�r=��>��� 3뛉&��G����ȓ#H���⟵:�eK���{����c�t�b��,�.}!�	�`�~�<��M�Zg��Cfk�A^"��Jx�<�@	$gA P�p 
�>��F�<�E���-�t�h� G/�0�tA�y�<�Շ�8c�*Q���Eo��	R&�`�<3�܃ �j��� ��zk\e)�Ηv�<�T
8F�|�`/[j�)��r�<�g���4�4q�E���yɆ��m�<�7���Ɇ�=�Yt��M�<��eE:�"P0�d��O�+���I�<����t,���5i���V��B�<�G�ՉXt��ǛA����K�@�<aT�J�h4�)r7Y+^�u��X�<�B�ر I�%C� �/b�)*���~�<�Q -���`��IM��!��q�<��c��[ж��נiU�yI�ɛg�<�Ջ< fʝ@�g C帘�H�`�<Y��#��"U+�_���a��^�<��3g�"�S$�5�̸��fLE�<I�����R �2.^�	���1�C�<�&F�O�0X��@%�̤Jrl��D��y��!	DL��H�Ng�i�ȓ�y qF� �^iK�煒AL�=�ȓy� �蓩�`Q(8���n��.�aQЅG� ���ŌAQ�2��ȓl1@a�0�܁-7�u3���%�nԄȓ$��xk���[B���a��K6���T��-i��.u�3�	�>x8h��S�? ��CL6)�!����2΀ )�"O�4
JI� ����Q�L��B!��"Oh``��.<���� ��Y�Ьq"O��cN
-!�D �Iݮ�ȶ"O������{���րYl4���"O��Q�c��^<�A[��^2�y2�"O�8I�g�h��I����'Ez��"O�L�PN��)@ّW�8E��t"O<���)̠.�E��k-x?� p2"O�+S�914)��ƤW����D"O�9��I@"�� P���E���"O�+�Oa"m#@JA/� 	�q"O6A �,�"�@�t$2��yPc"O8��:���N�9vm(�"O*�{��G9o��e)f�F�D*��0"O�	��ѴuB����� �g��Q'"O��;&�K*>`�e�rOϼ�����"O�I�BdE,V%AË�8K��b�"OT4��@W�I5dp8A!K+aB��%"O�����B�SB(`с��
I;�Ȉp"OY!��	�[4��R�(96� �ȓ(~̨ �c>4�����P�����"�^!i���E'��2pc�@
���Y�yX#JC�}r`V�J�����6R��K�3�ꀂ�g]=Ҕ�ȓJ�^5�D�� Dz�$(50�Y��.�Bl�T���s��0��
��J��ȓh"�Ⱥ �J�5�:(
)q|��ȓ{��%�`�E/Z�\I2ƃ�"J��̄���u��._pl�d�(��L���u�5�4�jJ!fwx���e�&��R٩I��J����"�����C����� Rnh-���\����ȓ'�|Ȼ3�����13`á��x�ȓ%���ǉh���Ʉ�vA�ȓj
�ŁeJ!6U�E(�(]/��+А��3���6�~�k�.�
{&�чȓ�V�1� @�pn�핋��̇�U*t��c�7����# �a�Ti�ȓ:�-��V��0y��U���ȓr�4y@�(�!
<@�Sşb۾��ȓ} �<�te�49m���un�o�dP�ȓ\�t��#�6u���Vk�9ԄȓC�(Txa��3*R1�B�7R����h��@��D��p��S+3�l�ȓZ0m��m(>v���`$�h�H�ȓ'�xj�I�;nkBC��]s�����Es������}�n�2��#�$���*�;��L�����C;�A�ȓ/?�$�@L_�xa��!ǎs�h!�ȓ ������)\��&bI=Rʅ�ȓKb�ljb@A�A3�%�c�Ճ �ȓ��Iu'�B4�YIp�W�3�V�<����$o�Z��Ñx��C6a__�<��A[�X���$Ay�A[aYZ�<���5M�1��#1�(SA�R�<�cHߝ}����5bJ�|���F�<�EM��*r�E2�+�?dw���#�F�<1 Y"�D{wP94j�"CB�<a��܉G����ԅ�-{?`! bEc�<���B�DE�)�f%'T��p��DzdB�+B�=�5�e�.7�(�ȓwzh�%��2D�����l�"�,��ȓ�Ё'��1c�4� �7߄��S�? $Z ��&	v]jB�nl���"O�C�K"Ft���1vfp���"O*�K3��|�	���d9~�:�"OhQ���o�Na��L�zF�Y+4"OV��QA_1t��P0t��s��z�"OU��&R0� D�r
�8>��{@"ODT�a�U%x�L��ȝ�h���"O�gHm���+���?����P"O��q�?��}�t%�o�H�`�"O�5{!,�;3��V�(.��y�"OT�q�ɟ�r��h��.!����"O̅���ˣ�A'�	�T�I��"O\�Pu�(��d�* �Q)�"O�9@�Ȑ�L�
�Rgh�"���q�"O�`�PiÃ F��iZ�aߢ��u"O"���ȺQdF\�(�8.��e"O$ԣa�Y2�2������"O�`��L �#��PS�>��� �"OD�+W%�ЭK��N	<�$b5"O ��@��k����N��Z�\x�P"O��P�>&,Zəg�?*4�`�@"O�)R�̑�x�A�+72L�#"OT,��b ¬��$π!���1"O�M(D�0��c��3dz���"OlyA�	�x�xԘ��F2?� �C�"Ob�� a׷m(�%a[\Ԟ5�@"O�]��1;R2%�r`�a����"O�!ɐ�Ņg�9�A
#{�x���"O�aw�S;�H�"CՖg��C�"Ob���c��R �P7]�$�a�	�yRaY��^�C%�&�-����yR���5��z拊�.ȩҌ�5�y�MjU���ϐ�"�\@A���y�#*�ݹ���rA���,��y��7"4I�-7#ؑ��̇	�y�

	A`N���kE��*=�u�Q��y2BS1/M6�X�$M���`��j��y���\t�4�=�(`�6c]��yҭN�r�R�J�$�0$h�H�y���&|d�0$&�"Yg���D���yR��N���c4
�[�Сxdi��yR%��f̝�p YL��)e ��y��@^���i�U)��0�$!�y��@rv�P�$Y9
�Bt(sA݉�y"OH)bl؁9WL�8|D��C�[��yK�o���s��֥/��l��׍�y��!F6]�aJ� q ҭ� �	>�y��(=�pp��b1���(] �y��$vtX�E
 [P�C���yҊԃoI�A�#lқ~��T0Y'�yB�;���R�ox�9���%�ybK��"7���4�� x�0���GH��yR		�B�ޘS�ń�v�ReBA����yR/�
���"	�g>Q�0,�y�D��18���A��)ԆY;��	��y����RA�ȡB�1���&�'�y�Ђ&��DްH��(N� ��'x4\��CG�MH���e[�K�,��
�'� �F�W1QW�l#Ջ�U�=�	�'&��`bʵ�p:�=S����'���u�H.3���W��
��Q�'�,d�I%�X�!� �`h�'���+�d	�Ū�'ƅ}���
�'X��J��(#b^�s��<<4dc��� �T���� 1:��wX��$�g"O�%p�ڼ[���Fg�"���Q�"OXJơ8]��qcƀ�D�N�Ɇ"O����$�� ���(� T"O%����B�&�	�B���""O�	��IK4�z����q:� "Ob�0�	�Vb�{��֫Fo�t��"O��0�� NN�a�,��U`�"O8B<юU"��tAz�js"O �37�^�j�F "��L*z��"O@Q䖪-14-���^�w�`�""O��!���NF��qi_��@�{�"O�la��������Y�(�1R"O^��� ��m"�摆H�8�)r"O(!�畷}pF�ó
��He"O�d`���YpV��'���R?f@�D"O�(7����� bӷ'"�1"O4�aġ���x��b��6�z��e"O�!w�3x��@*�nڀ$�xP��"OR�`���G���*�&˄�B�"O"�B A�k�ؠ{bj�e��J"O��ʕ�X]�R�I�hO�b�\P�"O�𴃝�NF`@����v3E"O�h��lR�YU`&f2o����`"O�4�2-��mRe�]�(�R"O�)�W�M5j�d�+acq���0"Od��ք�T��mY@l��Uպ�T"Oj��	����2C%��<�,�q�"O
�ᎹA�@���c�5�D���"O\��GHˎI4�%����^�@� "O�}��#u������z��u��"O���dJ�%ӬiXp���n���"O(-���J�5�,�W��#�B��"O��S����1�V�Ч��(Z�2ق&"O��&��߾�j�ی<�܅Z�"O��T��DW������x���'"OR,�G�����'�U#dvI2�"O}J�$N�R<�A��xG0@�p"O��Ǒ�E*&�
q�;3�d(f"O
i1�� �+�`�
^�W6��"O.w�ɟVO����Ħ/�B�"O�!!�R2=vd�CI��l�X�"Oҵ@��L(���Q�枽g�DmZ�"O�� '�B,tP�2E��D}
�b"O�&�[Nj!�'+FV �!�"O�djvMcv���(�<`0���v"O*=Y��_G�������:+�i$"O��H""��� �bi J��"O�<�bb�5]a����B��("O�QZ�e�:7&DҀGء7�z�9�"OX�ᯀ ��yu-�`pص��"O�\0@�Tn{r��E�+!\�A��"O���CɋY[ܽH���+X��@V"O"8��ݗ)�#.A~��c�"O !��!҆'��iS2/�3fh��"ON�Àčs�~Ⱥ�d]�/V��; "O"����m�`���O+N��T�$"O�hHg(^ˈ�
��
11�ְ�3"O�i�Ä:�9�"M�.BP�騵"O�1��;l�x9��+�,r)3&"OlT�4"#`A��d��"r���1"ON0�3�.^��g�͔"!�) �"Ov��U���-ҿ1�C�"O�a��< ��Qm@�!����"O� ^�`�������Du�(�P"O��bk�4c�)0�\�L(�"O(�0`L)}"ZXb�;m�D�z�"O���O/u;�a���I��-@"O PpH��"�4zb���$�|��"O�yC5hсn?���s������"O��qM��Ȍ"��ݹvwaۣ"Ol���ݙ�j���� 0l�A۱"O�� ��A�Q���f�q(�"O^ِ�ǋX�PX`H]�I��	R�"O�0J !��/�r)
C�='D�L��"O��!��4SdJтde�IFl2�"O��[���7f0<�#^%l^>��"O��u�Zoޖ=�bU�EYd���"O�%+�W<T�!�Sˌ $ޅh2"On9%d_JE��aӉO�;>��0"Ot%S���r�D9�F� o��3"O��A�O�}�fh�F�?���a�"Oj=K+� �dY�SdR�s����"Ot�Sv펂,kpC3��?F�4�"O<��� i�
p�bȁ^xd"O@��nD�W���S�KD8p1�1"O����aNT�n��k�2L/��[0"Oʤ��H�T�Ebs	cpZD"O<�kf$��� �hL�
">��4"Of��퀔ܪ0[7Nĕq�(!"O�TQ���a��IB3��N�I��"O֌3i�1�"��*?0��L�"O��*W=\���vi��0��%"O�	�
-K��#F�4��01"O��������$P�G�.9+��"O�-B�锐:S�����vG9i�"O }�`Aŏe��M��e�1J8�Q�"O^�sdG�?x~� @��O�\J��U"OHѠ� �	��%�df��>J�1"OԸ`ƣ��ZQ2�dA3 �G�<����i��3`�^Q�eCr�D�<�D�
1q&��a�G��
L�HC�  B�<!�a�%TH��w�3�m"0Ji�<1���5K��|h3
\W���Ǐ�b�<񵂙�~���[@�;JHx-P� �\�<�#I�!�vE�k�7E�}j�Io�<�M]#j�J�� )-�����l�<��U7:b���L#5���䩈`�<���F���@���$<$j �X�<i��\$�`�Q�]iZ�%!GS�<�"/�g=��r�|R���pTX�<�e�/	���͟��ܫ�h�R�<���2��Iꆱ$��s��BI�<�vD��T�{�ƮDd�:�bUz�<Y2�_�CV�RQ���/C�PT�r�<ACƯ=��T:ԆS37������k�<)��,G;@p{��kx�p��J�e�<� �
![�~�(g�1Ɯ bB�W�<��Q�[���!,ˆ2�4z���S�<�c+��pHA�`��{L�(Z-�I�<)kǅd�=k�>R�2�LC�<Y��X�)�H�
���4Y�5��Fe�<�)EI9@	��w#B���m�<�4nYE`Djw��rWAs�F�k�<����:��`�В�N��@�
m�<�Q���YӪ|{*ݙ>�e�Ak�i�<Ir�Ӕ�t�k&a_<?�D`��{�<Y�M�yT���� ?r�v�p4�B�<� tA���\���7�U1D�A�"O �zk'���q&��8^(�"Of��u$׳ ]�be�Q!byF1aB"O��AG$��8��ӸTj�\�a"O.t���PE@nHB+�-3�����"O��	����PŨƉk��C"O�Q�v�LT!��6Q���p"O�=�2��)jb^��MT�;�­S�"O��iCM��f� �Σ��2$"O4܂��ZvU(})�1$���G"OH%����@�4���h5ez�p�7"O�ݺW��$:j���!�[�"O�iD
�c���0�L?*�a�"Oz�:�c��ҽ�'ԩ[	>l��"O�Q���F#�j���
l�X���"O����o����T�RG͏���Q"O��[��);P�Y�eg\\^d�2F"O�����>��щ��$kD�0�d"O&�ˢ�E t@��Ɣ05��"O�,�f*J2v�p�Ss�@��"O�A#�;��$R�]NޅA�"O ��+��S�H��k�Fk
��a"O*Aq��M�(}���W�>���"O6u�T�3UVT�d�Z4fM��"OL�¥F� !��8+���1A*�%�&"O��qo�W��x���Z"4B8�T"OxQ�� \�e��d`���z�l(��"O2�@P�a�^�k�o 7,���8E"O`Ek�/	!P�K�.؞AT�JU"O�������ȸ����|m��h""O�H
@�\�(ZFp�fl�$|[�49�"O��@��U�U�Ӫ��<��C"O\ڣ�F�
�ƀ����e�N��"O^�)ďߏGC\U
Ӧ��vԒh3�"O5j�BB��(�܏lȆq�"O��X�ڵ_�U�M�n���
�"O��s!�Z8Dr��Td;_{���"OH�rL�:�UAb# ntr�Z"OrxCE%Y�~���ΐLq	��"O��!7a�,��㢢5M^ƭ�"O^(1�F>�������~Pj��B"ON�"�n��g�V�7�VfP�%��"O�ba/^�hs��z!�Rb�l��"O�UBZ�w��!�wȄ5V�*�"O����G[kܐp4��BH�"Oby��A�zp�@/�f�k�"Oh �A�V!B��@�C�SͲ���"O�����¤C��M�
�,Y���S"Ob��3	VAs����(�J��g"Ov��Ǎ�F����gi���E"O�Q�7c�\�1�F��ΪXI�"O�Y�CˈmJ� vf\'L��X:`"O�LR��<^<x��r'�3f�͙�"OBU��Y/��Ēg�T,��	�"O~*0bT-��0!I�O����"O�`��s�"@��(^�(�"O�,�ugL�[8�4X�#V5�l�"O*��PƜ�,# e�Ԣ�W�d��"OP��%H�%�n��Y9���g"O@�&�Q�,�IX�`�;k=
4�"OVL����g�{�� �|��|x4"O\����f�T��.tRL��"O�L�FA���|x�E�IjK�U;"ON���A
&��$�ԔQϲ%r"O� �e���6!�jE�a킡5��Das"Ob��� W��ɱLW�S�"��"O������Jb(��劀8�R���"O@h(AeݑoLNp�ʀ�w�ҕAv"O�Ҳhiޙ�BV�O��ڣ"O@p��#Ph��0��s,�-��"O����+G"iU�	2��R�DLB�"O�0�E;U�R��AA/0�j�"OJqq��R�k���5G�;J&����"O�Q� m�i�DA�P������"O���F/H$ᒹɢ*۪a�Tw"O♻G��7�ց�dY�Yd����"O���5����M2��� OLD�"O���դ�"b�I�B�E>�3�"Ot�3N
�*ȉS�˩.^��W"O��k6HC!:�^�� ��m�	Jr"OၖT\���n�L3b�����"O$Uk�ũ:\�����T#�v50�"O�AR���ZT��ʈ���"O޹�'I6ֆ��?��(��"OTw�#3l��5�Ǥk�¸4"O��`G͜�zm���@-F�<�R`"O��1�Y�j*e*��?a�"�C�"Of��eHM�D���v+���u"Oz��w+��/^n��c%�0Z��l#q"O���HV�&$��!c
�9��a�"OV5�D/a(r�h:��3�"O�8��N5`P�Ɂ5����5�6"O8�e�л	u`���(��rlvX�g"OF���� �F �$ʡ��p����"O���V/L X���"����N�A�"O��b�G�7A	P�"�"M��"O,h�g4����㟩5���"O�!rcfԚ`Nq:@K�!�@�!�"O&X�tH�{rPE�o
 h��ՠe"OD�%(ޖe
�yTcܡ|�~)�e"O@�+	+�� �AU�Ҿ�a"O��z�#ÄX��3�P)̎��"OH1��O�gP�e��)S����"OD	&��f@fHk��S#v�
e@�"O:�ɕ&�3c��
�`11�XCb"Oԝҵ���-��� �<E��"OD�; �yO�h!_�k���"O���`'H<p�;�n$F�b�Z"Of�"g_�&�L��CC{d2�"O���C���b�-�_٠H�u"OVQj1��;a^�uk��|qi�"O��dʎ.ڮD���Z�|�pH�"O�!@E(K�ĩgC!�ؽ1�"Ot0�� ޿����4 St����@"O2�J�P�t��U`�
Cq�A�"O6�0�G�)@_����cR�_6 )9""O�l�1e�I�}"ŢϢ,6�H�"O�!17��������Ƌ$P�	"OR���HWlh�fo��88 �c"O�`A�^�8�xՁ@N�2vN`A��"OFtp�@ڈ_� ْ#m�G��А"OP���K� �r��L�W��P�%"O�-�0�8@���!��:S�i�P"Ot,(���Q��j�f��i�@��"O�#��NJ�pGK(`�,`B"O1�K��d�l�@!$P:q�J=�b"OR4
�)�	?��e�ТV�*(q�"O�a�&I���Ј�i��T{�"O� �m��ȕs�2x �#*3���d"O���TK%p�L<#FlC��Z�"OX��p'�;�F昙985��"O�� 5���1upD�p�Hd��B"O�� A:A_nik�aI�T.�Qz$"O���NƫI����#cԌ� |AF"O��z��ļ6p�pt!�0)d��0R"O�0ضG	�uH��E��G4|�r"O�[W�^�4`(5��'�����"O��+��@� �+fF��9(�"O����
]_�����_d����5"O��@�Ʃu$�D�bE�'��d��"O�����A�x�$�`}+�"O8����ٱ2������6#�>d�"O,4i$^�e���{�m[�-��!S"Oz!(Z%W��BB�K��P "O���fc�8ȳ�SL�1:�"O�19a]Y�+>F��@"O0��$Ϟ�B��q-�d�5"O���aN�v��Q�
�"�ڠ��"O�Q8�I/1�1HѮ�8 ���ɣ"O�8�[�]��A�� Z��l�"O�,�N�Y�@�e�P`�u��"OU%���q}R3�S�mC���A"O̙��
��;���Z� �R7�T�U"O���Uň3*V�؉�o�?8 �&"O:QA�*%�6D�V�Q�r���"O��6BM�i��@U1!�^XCF"OVܹ��L3K8L�d��"ȑ��"O�����!UR�p"/C�V]�0"O�P�*~A����U���kD"O�8�HۃT"
� T�ːtnb���"O���ujԦ"'ꄋ��75Wl��"O
��N+|zFe�	�/WEb8�5"OJ�����:�9�"�ոu�؊c"Oxs����`�2BoʐF�PJ�"O����[b����al�8H�m��"O�(��LMI�*�2��>Y¶x��"O*�A3H��\ؚB�ɓ!�IJ!"O
�	1
ƟN���`mº?�vȣt"O��A�=5t�Z�L�;�6�Q�"O��e��>�c���<3�P��"O@��D��)�>)ؔ�U-GV �W"O�J��ƭc����C�[x�Z�"OȠ��ڷ7̜Q)����2�شyA"O���bV�=�0|b�g֬ t��c�"O��kq��:��`���Si0��"Oȳ���=^~,ْ�Ι�?h@�w"OLx(�!F�z@t�22�"UQ.�X�"O~�{���:�U�ٍ4���T"O4T`raC�v!��aOY<�"�{B"Ot��:V��M�����5�"O�H��珂E�])�o�>y��"O��
vk�#��x���cH�5��"O�|ZЋ9Vs��C�̊�QP�A�"O�t�5���(�� �&kP�Y:��r"O<�!^Csv%3A��7�qa�"Oݲ�Ι}iމ�D�,�&��V"OR�QS-P6|��S�n�_�R)��"O���dd�mڬ��3j�ZF"O���2�R�V	�vj
([��|{$"O�xiE�~�"�����"O �ˁf[%.}B�C��B�@g�di"O�pz��9�.`@o�2���V"O� �Q�`� �Hͼ�K�����TZe"O�� �e�%(=V%1DbţM�,:�"On�kU'�3�u�֠W=Mz�p�"O6��6EF1�I�헕�ؼ"O��Q�Ʃ1�1��*�J>�Z�"OH`0I�?�(�jU*Ȣ�|�Q6"O씋f�W�N %�C�2|ƭ�"O l{�׻dg�Ah���d�:�r"ONP�1��<}��h�!Ąk��u@&"O��d��4�Ԑ�D�דm��It"O8��1N�]B����^6��1��"O�����L�?gz�����Rgf��s"O&������� D�@�B^ҽ��"O�(�˒+<ͲPH���'\xk�"O��c�@�&�m!�@.5�|D�"OT���
X?,���
�Wސ�4"OX����I�Th�FN�P�.�c"Ox�꙽#uJ<�����,�If"Ot�B��M{�1ʡ̛?~�*q"O^P:���C0LӖ���I��P��"O>�"��� �wAZ�P�y�c"O�(�e`��Q4pp*�OZ�{d��r'"OF�S�EW4���/�8BrH{F"O��[<,[,�@ȇ7I��M��"Oj�R���W������Қ0q���`"O��!�$�0����Z�k���s"O8�T�6"�j��F?^�|laF"O�m �o��*���E�V)m|�@��"O �rCa�-'yz��� ��<h,Y�u"O�x�g/O+f^�ig���>��`�"O6!��F�U�t���oÑ��1X�'�a�S����.I��N`�YB�'v��#O�������мH��q	�'��$A�aB+䄑�͟�s���	�'�0�cSh�]I�5���C����'�����!d��E�E��A�����'� (���J1�Nu��N�h���B	�'<�h��C2	G�<�g�ؙ)�-J	�'�@h�oĤM�z\��D+��0
�'�����J�w,L�K���a;	�'���9P�H�,��D��Ȕ5",8s	�'PPD�F�O���kP��0K	�'9�E�� x��	GQ�&Rpj�'8�!���b��!9&�(꤄˧�yR�Rpnt� �*� �h�V&�y��	^~^���I��ْOȚ�y���
;i�仂E��d�*��&��1�y��O�n�8m����p�Aif�̲�y"F@N=$B&R0I~��x5L��yr�N#K����`�B�E��)�q��y��Ǎe�6:�KG�,��d
��y��y���c��	o*��Ǘ�y��X�G]�9Hqh�I�P �W�֧�y�/�7�R��@�F�*�{�G��y�m�4�4L�a�9����b�ː�y"�--NEHf��))�:�9�W�yB�r��E�a�ٺj����@]��y�Դ}�0ѻ�o�9u�P�0��ч�y�mԖ��x�)�$fF�`A���y��е-�@J"�X#g��I[vc�=�yB�)$A��  �Q�l/:�p5�"�y��ˁ�8�@��j��Xc%@��y�'H�&6��e��4d���tG�6�y2�X�9��iȴ�IHR�"�`֒�y
� @� PcW�M��Me�l��	��"O�}�v��5z\8����=M���qa"O�MP���@�V�H>��"O0!%GT&k�8-�U�����yqW"O��h�o@�^U"�O�9�,���"O�,�Z�uj�%�ŏ_�g�~%i�"O �qh�,9)����&�$}c�"O�Y�JM��z��p���|L��W"OF	s)'s�.e���7\ɐ�PV"O�(���̹�ĕ����"O@�p IF8x��q�UH T"O�,�DJ�ltd��r���J"O<���#��74<�1"�(�nŪ�"O�D�RGһt趀���+d����"O�i���J��ͨr�Щt<"`j�"O�YASj�������^��C�"O�x(s�}@��Fh�-�0�$"O��wg�P""3�`��w�\�ɶ"O��9  өs=bL4� 7��M�c"O��ç�J<ds��!kr��3�"Ox��� ּG-�A�֍K&UU���e"O~yJ�X�I��٥KYL�H��"O6�Yl��:ˢ��M	u\ D�"OPYa���#�P�i�hD�R'"O(�Z��V�ypu�M��Q�"O�(�@i�n�P˱�;�Z` �"Om:a��C@f�i#䑹VWb��"Otd���7h^�H:�NS�Y�"O��{��� 2|"��ᅕs��2�"O�A���Q�������Z��"O�(��(�3T�����XA�"O^�À�](ځ�F���HZ%"O�(Jd&٘h�L%R��p�P��"O�KtF�7G�n=�d@Xz��0�2"O@�����b�-�$@ m���N�<��kӧN_���(�t �m���t�<� 5�,��w�4^D�֏Zv�<!1+�#F,�pp-��0/jmA��M}�<	&̝2�����	��8�u*�N�<Y7���p��P ț�e��yjJAN�<���|P2bM����r��G�<�Ǥ�D����ġ�����B�<�W^�-(�@�(�� :#��A�<I�텣q��Q��@Nd�TC�A}�<�A��V&���@E��*ɔ}Ғ��_�<IrK@�HB�bW-T)�r�w�<�g�U��i��n �z1jJv�<9��]�V[�}벭�W%�tz��o�<i!b�*J]���g��?� ��-Ov�<����W��݀T��9\le��jl�<��29�`%C����r`Zs�<1��<zY2�3j".`���	{�<a4H�4(�pMI����}^R�ꢨ�N�<A�Å;r�� w�ژ�d �pnXI�<�u`%���%,�V���a �~�<D�SwE�|ӕ�X�/��1Q��W{�<��!Ǒ<dJDf�}�:`R�j�P�<�B��b�N|�qό\otX�W"�J�<I��� T�IلΈ�h9���I�<��A�*"�Dj��Ep h�j�H�<���J�"���{�),J�XPd�^�<���,Xy�<��hI2]}� "��X�<��ìH8|!���B�n��k�<q3�> �Į�/' СG/ZP�<� �\���;=赲"$^�;��ѕ"O�K� �>�n@�"�>s�~��"OH�$DHJ�Ř���F��[�"Ot�Z�JT/&�,��d �|xh԰"OM`I�O��)��(؟bdB���"O�dX��]o�Ӆ��F'�� �"O90e���62*�;��]p�t��$"O�����3��4��*7���"O�\	W�p5h�$���f*֐�a"Oι��� 
��h&�J���X�a"OB��qB�0v�1�Ac�?1C�ؑ�"O$�#r�
>R�z2b���"Ox�e��
v' y��#Q36��Y�"Oܵ�Q	QikBe�V���Z�i�"O�x
��G�����LR?��81"O摐A��)iZx�����t �"O>uؕ��j��T
��B���0r"O�$:���!����E�"-��eC�"O�i���WD����$ۜ�"˦"O��a� ^;�fbې	3����"OPHW�l�B��qF��A��"O�)����,�Z�D�h���`�"O(����<|�Ss͍8�r��"O�A �+�'0mpl*��D!o�9�"O�̀Č��B;�١�P#Sd��	�"O�UAriܐ�����Ly��y�"O������$L����	V�晫"O����k�25:j�#���$�87"O���[��LAH�DS.�๺F"O�8�rd	p���pУ��o٘���"O�q���۴Ly>����T���h3"O���A�٩�N�bՃL���h�"O*e�Al�3um"��@�=;��p��"O����ɟ!�4� NN:K�d�"Or�+�] /i���Z*��ɒq"O����+�<��+ŵ��T�-D��@#��|đ� fI	w�)��*D�X���G�X1b��
-A� ��M#D��KЙO�ػ!��5�Ĭ"�?D���6C�:π�Z�H�'�P)�a D�H�
�ZY�Fb�7sV\-x4�*D�踐�E�R��eP�V�r�`*q(D�t���,Y�xHo�?S� ��c�$D��z��د`�~L�#+ڪq�R��E5D��!'Fr��9G�8�����>D���eƲ4~<�'Wy��@�P�'D�y�߲PcL-�QdS�{o X���&D��@s�څY ��肤])jN.�;�#$D�Xh 
�e0�D�&Aj�$�ua&D�����o�<�h�Z�#F:H�3 8D��������eiU�� ^�J�+D��Cn��L��yإ��94�V=А�(D�<���A=R��V!�<%X�ǋ%D�\��[)R9���,�0r8	)R�?D��� cٴ���ټlܥ�D*0D���e!Ley��X���_�(��(D�hr�*Ax��y�B2{�>���&D��k�8p8M� H��,!�g D�0��B �i�pp�&�
QF��Ӑ�=D��;��0�,��E,��oGp��:D���gǋ p�n� ���g�@t�6D���`D��5�%�[�gb&؈a/D��1�=� ���BU����2D����3G�^�����;T���1D�� �1�B�P	jN
 k���}� ;�"OJ��		]�,�c&�(q�}s�"O<�����]4<��w돼}��}P�"O4$�Iֈ4`���_kz �"Ot����(l;xx��ѳ/ ]�P"OƵ)�k�X���DQ�<G�e��"O���ۂg>�D��C�y>l�Y�"O~��@��]�>�0��2e�2] "Oh��/
p��X�@�0k���:�"ONᥤ�?��}�V�3���õ"O(H���W'��m��N�#��X��"OPL��L�mv�iÎ� ��LP4"On��ࡏ�-~�iŧ��T=*"O�`�4�L9`X�}��� �Z�NX��"O04$e�vL���DD�Uw���"OP���ͼB��5�۫k�r���"Onp����'i�6�8�KE+ �ИZ�"O@l��%Y�sAJ$`�i��V�x�#e"O|��Aa��{Rܑr�1f�@���"O��1q@
6+��8���t�ֹ(E"O^Uj'��K�Xt�@a���D��W"O�[&�G�`��])�n��u��Q27"O.IZ���9��H�5d^�p�� �"O��!��wW�c��1i�j�I"O
�1T �/NT%�U�۵�JU��"O�јQl��R9�E�CM��Jw���"OLhq2"�>�6M���3�"��s"O��i��ߥo-^�xGO�1F/r�	�"O��p�,U:^�����7p]q"Od��e%\�	��yb�k><js"O�-��h!O<LB�!S�2��"OT�y'�ݮ��<x&�W�M��I��"O�QU�ptB�����(��ț�"O ��b�Hs<�c+Y"{�� �"O�v��}�ʑ5�Y�$<�hT"O��!��ʧ'lh�BH�k�M{P"Oj�6bY1L��i#4���|P*�"O������*_�h��#ax��p�"O�b�F�X�mXV��P��y"O���DdK��DYhG�Y'zIDq�U"O���ă��0 �L�1G-��p�"Oh�sEˉ�HKn<P���.��P"O�0fcܳk}R�L�,��H�"O\b�Y�Y�e��*�' ���Җ"O��&R��}'�R�/��9pE"OL0����[B�A�T0��ɳ�"O�+AmP�
R2��$�:q�G"OƑ�s�\7�2�{�!�-�p r�"O�yq�+dSج(@ g�h��P"O:͐�o��h<2`L+��+�"O$�)�D��9��!Sh�����e"OTс0��'y��"臱U��q�"Op�X��ђ(76y1����wmV-��"O�Z����u K�'Z�,jV"ON����]+z�P�Θc�Y�C"O,�T�������z,|�T"O�����R�KT��!e`"O�C�M�@������ 7�t�D"O�1d���l�d��Ì�`�( r�"O*<#��-u����6kצD��a�"O� ���zZ�mk&�#<��@1�"O$�z"e��9��YS�c /#�
H�$"O����L���!����d"O�X�� ޱ�� īqq���"O� X4dJ��P�s��P�dJ�R�"O@<�"�A�$�fy�5��a�0�X�"O(�R��X0q�����P�)�(�r"O�	�d(^1i�V6���w ��"O6�q�ͧ�~U�6I7R��("O�Q�#�҆8'�)ɥ!:cc�[R"O>��C@��t�����j�(��"O
��%
�
�9���.,�jU"O~�H6�����;G���u0�x"O����1A0�jո%-�Lb�"O1It	Ԇ��Bb�> �|\"�"O� ���
 ��H��)��(2"O�9rg�/�dUɤDE�8`4��"O���a��B��'�zX)�n�<u!�DV�3����&`T��Z�k�pB!��#Y֢}�/��-�Z��I�y9!���5>h��&cU�5�\�d��I�!�DB�W5dEp�B*h���ծǇ~*!�d܊ �h�E�T,ToT�7!��3"P GV��y�7�P�=�!�d�_��`��R�E�$�S&Z!�D�<y(�-cC�I�*��&)S!�d�3F�j ��2�}���#�!�� E��RuK">t��#��0J!�D[y�@z&��49p�q𥔗8=!�$̸E�����'WVhd
r�3!�!�d�@Z0YR�ԟ"K4�K�dӢ�!�dL�s.��`'-ո��ra�Ԡ4�!�dZ����c�H�"l|`U&���!��a�u"��@�f4tMy��
�o!�9QdV�8r!��A��i�]�u�!�d� (��������0�����!�y�C�j�~�є�Ia�!��߈0��!O��#�t���T%�!��)��,r�I,u������66�!��t]d����<�B��^�C�!�D��Ԃb":6qX��V�\��!��=J�xv��4�F-YS��B�!�DD�X�b�z�G蘻 Y�Bq!�$҅s}�,0�� h&A�t	?.�!��,�5˗"Dc�1��eA
�!��Ոc��Fl�r�Be��풵QY!�D_�k�rܑ�����0;��
�-:!�$��o�\d��h�!�ʘ+�W `�!�өj�p�#!&&�pH��)�)Z!��:�����C�>1�fyIC�A?!�d@mPy����XuL�I���M !򄚛^�d� 䏽���y#�.N�!�L�Q��"��S�A��	Q��F�'�!��9m0�Zt恑P��ɱ��'J�!��*!+��A�I�}��H­�y�!���}��͠��,8��p��!g�!��Βl�����ʚ#]�0�J��5�!�Պ�F���옌_��Y��2+�!򤂔l���f�\ {��� 뜯h�!�� 'Wf���B�O���u	ѧG�!�F�?����Ό�i ޹�W狚�!�d�ټHv'C/aVz���!���1+�=���	'=��+5oM�mv!�$�Zh
<���7ơ�2�B
o!���C�\M�)��(9-Z�oR�>�!�Ď+EAr��>�E�n
a�!�d
6R9�``V�(���`���!�Ē�@�N�ұ�J�^�)�`�,�!�� ��.=D�Y(O՘����i��IZ�S��Ms6-X�9є3�_����8ta�g�<CV	�T���DC�[K�5�0�L�<i �_.XѶՃ6a�1:�59���D�<���{ڦ$��h�/xV:(�ˌA�<� `\>`6��5��v].�pAfJu�<�t�ƴn����שC��F�W�<�􀜧-�I{�k
�y�  )A�z�<����^p����/�xLR@��~�<�B�?51���g����ҔbSœn�<y�B�
V�d�&.�
{,�5([_�<a��3�eb���B(L�� �ȓR�倗�Î:�jXB�Ǵ]��|�ȓ#G��3��@�h���4Q�t�ȓ6�� �O?^l�	�A°�jI�ȓ���E�ɂF�:�a
'p�Z���"%*̱�#S95�.����!t0���n�yXqM�-7 
�i5ꖞj����Ij~��>���]	U��4��K�%l���F�<�..� %ۓhW�eZlɗ��E?��'�qO�#=q�����v+��rL�4�`LI�<YC�L�U	8��G�X[�U��VF�<�����@�T�Q8I�6�V��x�<93j )+z��0��1�����p�<!3B��	���#��B�s%�$��p�<�$
D�fzP��S�@)	*��K�q�<��CB�wňu��)K+W�^�a��QXX��Fy2�$2��6
�e:=Y�f��y���Ȱ��FT^��ĩ ʄ�y2$�t���P�lA`��8��<ً�o�b��Rgb�d����w!�Du����������D)M�-a��O����lG�_��
�G��<!�%+�"OR���_z�@-�B��R�ʃ"O���԰)q�����¬�*�!�DI
n�D|���$�d@)qF�3�!�č'����+�1nvݓS�O-Bw!�$I<V�z��E-QeQ$M���
J�OJ��d3g�P�Q�K!N2)"�Ow�!�%��)�,��"���a�"�!��Q?�Q�� Ǻl�V�"&V�uk!�]43�R$;�"ӺY��:�CإxN!�FA��t��':s۰M�UL��K!�Ċt�1`���ň��֤&8џ��=Q����� .��8���*�KE@`����"O��J�-��]赨wl^�?PjP8��'���B��	1�b9�,)F����s��7!�$�P�Y	�H�x�,���;!�DԎ	 H�J � @��9�J�x�!��	U
�	��D ��*QA�" �!�0.	���ٞ��Y�n���!��O�j��tE�&QJ]�f.n�!�E�<|x�4���E���5��!�dW*� ��9B���)�!�$U�xf���șjWr��d�۞q:!��I�+lKCV�������`�!��ш2w�	A�� J�����LH�!��_9V�N4R��5
���6�J#H�!��ÄR	�	�&���S��D�Ri	�t!�؈z��m�&�G�,
�Wh�`m!�Ы4wH����A��!�1h--5!��41i���L��B֧�3-9!�$����pf":�6�qT�D�%"!򤖡l;�B�� ��quG(x!�� ��c��ȅz<���Bv\$Yp"O�Hxw�*q���E	�%,0l+�"O�yj���*u���6�ޮT �d�"O�����Q-�i(t#ʌt���`�"O��A���{�!��"r���"OJ��K	[�Ī`F���`�"O^�S7
��)�-U-E@�|Ҷ"O<��p�H|��Ay���8&��-�G"OVQ��ώ#�&��0���.t��"OzQ��G�9
�� 1ÃB�k�
q�"O|I�'��>KN�i@'��?s|n�j"O�qa�N>j:8=�!6�^]��"OX�y1�Â8>>����¬Ei@���"O�C�E^�vY� pg�˭gL��� "O��f�JP/�����ܽKC��ؔ"O�M!.ǃ7��<��h�;|D1Q"OI������*q(� ���`�"Oz�('�ҷ)���)և,6���p"O���DL�:�H�`fN�m����"O�5���@,�<�b�N�i��5��"Ob�aŬ�&1�l	����r��Pu"O�uA�g�nL-��<��t�"O��$C��< ��뒈X~7�l�f"OḢ�ǽ6S��["HI�!@��8W"O�!���i�H!���̔i���#"O��f��RZ�Ə��$���"O
��&fmS^��S���n�y�s"OU�d#F��"qXa�}*fQ"O&��1����(�Zq �o..�
E"O�!H�	\�q���x�OPb0F�5"O8�@S�^�2�$qb��7&F@f"O��Aզ
gpy��#��p�<�`"O��p�ᝥk�Jy��b
5Pє�k�"O"��v���r)A ����!�e"O0��#�n��x�!�O�^�zX�"O�x�A�S	6c���5��7��A��"O8hKPm�	v���(����0D"O�8q�+���d�b	=B�M�"O�(Hp�	=$t�e��&OІM�"O�p�!�5�^,���
����"O�T�&LD�#��ajw�%nt���1"O�8#�咨��b%��"�p,#�"O�� ���u�a�4�O?U$%�r"O����F�*6eP5�a�XB7"OX�b�ƻo�;.�$�b&"O�M+�N��w ����)tHhAF"O��r���_׮��W�� Sq�X�"O,�bcM�] ��+g���W|��@"O�ಗ��2�f���jT@�`"O�E0�C�P���h�	�'Vp�	��"O�h��+R-~69�կ�.2dP�R�"O�lQq�B
o��`ą0`��R"O�[T�ϊy�`F��i����"O�8ģ�.<6 �����:��	cC"OBxY�Ɛt����1w��Z�"O���1Ĝh�
��W����"O4�	�"�]p�"éE!n��D"ONhqq ��d�$��`T���"O����K�@�\�s��Ȼu掉
�"O:\{��	�V��F
U�Ц���"O�q6�V6
�D�<&��{�"O�K`*#U6�����?5�4�Kv"O�EsdP![uP�)�bT� �f�3"O\���ّ/nȕ��� �=�ݪ!"O� l���U*%K8Ԉ�KӋT�ن"O�q�:WY22mWr�x"Opq0s�ŏ=�B���l�*"@33"O`�F��x��T"K�_�~}#�"O^ c��
�D#6�!�X�l�X"Ob�Y� 	Qo������u��-��*O��5A��w:AHG`@,n�<=3�'d��d�)=k�#�J�(1��� �'�tl`�-�z)����&��e	�'4v]+���#�JF�������'S��qJ�"9��͠�&F+�����'�r�3BÒ;5:,a��p�!��',8	�d��H��� TmW�cD&@ �'{0���۰�)���9`��p�'��`�!�
}@mSW���N�`�
�'���g�7�4� ��H�~tm��'�iv��
<������;0�{�'ϒ9��XFڑZG�����	�'����c% �pFZ̸��٤	9�A�	�'���U�A�FA��3�nG��z
�'�\��%��>�\Uce�0���'�J��̈J�vE�f�}=Ʊ��'�X,z�9<��:��H2w��-��'Mڀ��جe�̱��`_5h�,H�
�',�9P�E�>��QX���h� uS
�'{� �%EF!�q	7�ϿO����	�'Aat���dI�t��,K��	�'Ri��շ)�z�1b w�P-)�'��|h�"�`l�14�̻k0D���'AT�n܉pv(���@Yo�"
"O��Pf�Z��f�lbQ3&"OT�0���;�F�x��2)��"O�� ���?��S���*,
E�ɝ+<��  6yelH�1`�B��扇S/�hj���f D8@�]?pB��>]������yu@!�Ǎ3
]NB�I$L����W2ׂ)��܉t�,B䉷W���"Mӻ6� lҡ@�m	�C�!�}*eiQ=x�l`�/�)��C�	�L�zʣK,EN�J�d^�6��C�I�\BT]�amș34ⱀ��4I��B�ɛI�jՃ��ai��k0d��f{�B�Ɍ&�<e��O�*7��Q"�җP |B�ɉ �&h+�9|B<���E��6B�I[9Fm�lBQ⒬��#�0C�ɧV�|X�kD�Tpl9o�<�|C�ɑ]y�͐�m 5L	�8E�L@��'��Q�ș=��90��S�}��Zde�;k��ub6�G�>:�C��]��1��	R';�ҩ V(W"��A�ծ��L�"��
c�v)�A�:��Ąrq�0�s�´ u��1)���a�C	
��Hz�i��.Z ��4)���eڇ���e��X��e �L���	�`�]9����Kׂ��$(P�u  C�ɶpY�5xc
ГI�աM&@��B�	6?s����B�\Z���^�$��C�I#F�R�a��9�#� i9C�I.�ͻԬ!�J�r�KOir���0?ip��(�r�k�_�>L<��YX�8h�OԅRg�ٲo���R��)�4�6"O08Bbqlx��!{���P鉆�0|�ւ�=<���N���x�\U�<If"
�f�rS �/4�Ha%ԕd'��Dyʟb���V»@����g�?Y���qT+D��X�vOj�"�	�m��qi���kb�O��=%?��FGRg�Xt���F�^\��&D�܈T�S&A�	�#ӀB�:���b.���<� �(:�j���l�y�_�����"O�p��
pU���D�[+P�Pd{7E�GH<�P���uT���D��<��c&[�<	���T�*By~�;'���<���3ʌD��	�U�lx+Ƈ�Q�<��E��o���R���z�E�<��$�HA�E��AH?}̈́��W�G�<��ǝc��|*��#p��Ų�ei�<�Q�� '2 �Ōǅqk�1k$a�`�<�$��R�*Ik�B΀L<���.�_�<Y"D6�6���$�WDX�s"�c�<Q�A�9��
7�@���0�ǎUE�<�d�;E���ԲjU~��I@�<�Q�Y�c�Z@
��G*HH�x8�G���P)�셤Q�a}C�/N {�[1q*�h[`�D�y�D�����'@�� ���S"�Őo� �O��xy�=\S6i�g�3�ZY
�'�he��*N�AN�A�⡓�#���ᆪֆ���1�d^�-0�Nߝm�bm��'AL��$1������9kR.߼6Ć�Y��!6���ICil-b��1{p��	>ް���
��:SNi�Ei3l���-�.�����t�,�S��O}�uc��$�p� ���R������P������:I�Bat�'ƕ��	Ϫ���d)X�e�|�r���FM � �`�"��`6OF�A��y�$"a��8�|���10BmT�&��8w�Ħ�v�C�EĴ���'�d��-�fg$<�;i��$P�F;X�$@{҂إH~����	G�n��  1�hT�,O�����H�	ÓJ52A�0Ȓ�t��"�ؾ8Ԩ �Ó��0U鱧�/t��˃�O28I�`(�|�7m]�r�]Y)F'J(ʬ;͡1��Gh�5u���i��������;p~� ���0Ŧ�kd��'FTjC�V1|�LZ�,�C(@2!�"�M#���K`�]ۧ�BH�$�x�f��Ч���!2�a�I�2�$f�.]L0�A�.�t�����V�d�$�/%��2�Ǒ(;
t�c���
�$�U%�	"|�)�A� 7:`ະ��"ZT~�X"'�#֛Vg� ^:	`4kJ�N�TcT�O��9�F�_��)��ś�5��`вi�ޜ���2��|���	VX�nͩ*��d鋶)n2l��-sօ�Љ��� �A1�9��"�
�ֽY�M.u(Qs-��m-����)�[�'���;��F�%�n������t���� ���f�p�K�)
��Jwl�<���PM�#�h���m�.v��܃����~��nŗX���0�Z����P�1k�^p��Jx�x�T㘵$�W��:��bve�"�y	�OPġ6 ��,�h0��O6d3�/�lX���QȦ˧ '�00M� 28�])q S>B�6����`���&�1L7�X	��Q������(~d�5��	1m�1������(i&�����yg�&?�4���Vt�8*��<�p?���9�� J�M����F'[�*�hP{��H	��|��/�/k~��¢-6%��� j�G�'��h10�#�~�X��9�,t��$� �
�a�(׌�������d��TAp/A����R�I�!5�(�G\�K���0�ϯ$��yROܙJ� ��� H6:(b\��#Z ������~2c���8�/>@F� B�d�<0艁-�]�@�,��@�3`�_~�y��Í ��lâ��"/��p��_?y#��o]y�Xw�ԡ��P
 Ҭ�0/3jތ#�J8��@���(�v���"�N�B+@X�B�*ð@c����|�	٨fv�9'�A,0�5�$b� )3�,�6�n8��f��Y��Ò3S���i��ZjK޴�ft"�-]����aT��a[]n%���{���I4�3
�M���#��q;@�ɍ�>A��J�&Y�dT(��P��h�뒶�,i�u��
%�1Z�2ao%J�b���!%2&|�1@V%-���J��d6�q�"䡛2��+ˆA��I�F'�#�%UdJ�B���a�m�`�Ɏ/�lq��/1�|daA����eT- �Ā��f�*�<���Tҟ�����ʴr�:U�� ��gD��h��ɋobN	yĈ�(M"d2'YP��&@��h1�*ֲg�L��F�	������r	+V�D�|nⱑ��l�|	@�ױa�B��^���{�xm#�'�1�%�iĔ��0o�/oc洳��"F�a�c����6����;��хK,�L���h��ٱ hV4o�����D�<�j�9�֝
�b��8KN^��a	FQDlѹ �I ���+�T��ң퀋|p�ѩ	�W�X�(� �)8��H�֢����.R3B4l�nZ������OA����M�Q���;����kd�����H�܆L��53�L]�4�oz�9�Uc�s(����d(���*3g�Y<�-��		:K�lZ�Xc��c��:&�X01Q�>�ݜY]�ذ�M�j�\8��V�,P��=	�z+>�i�'�|͂ĥ
�8��.ϒZ�,�s���K)j"R�V.#�(���4��1����aܓVɚUB���**|Ivd���H�{o�������y�$�&�@�'WF�ڥJR�Vo�"]���O9T�S�댽^h�ģ�6.��h�'4��r���9r%�0D*!�$Y��2$$
�"lD����n��z�P�m�?6th���'Դ�WA@�~ �[��.4���'�,����U-K�< ��O��R�',n���3{�z�I��$�$�	�'nڡ���U��P��U�7۴�A	��� V`� K�i"v�I)�&t_¡�V"O��bdET��ceH�2�1"O~M���E�9��< �H��nx��"O�I��i%%�(�9Ӧ��D�9`"O�D�*O9)�Z�FR(�H�(�"OF|����i��}Q片�X��"O&��Dd��"a������`�"O��s�Ϛ�t 츑Ѝ]"~�r���"O,�����x�Q̕$I����*O�+�hڧ*�� ʵ�����i�'�Ɉ��Ȳ8R�×P��@l��'X�	 ��'$��Cbڷ�� z
�'_$�W�]�L����� �*�3	�'E~ q�F�E�� �U@:��'�HAK�&���J�0B�Z�'��9��c�ii���E!:���!�'�ā�&���>Dtf��;����	�'�<�c�(�,I%�&�
3�qz�'����K�
6�(piv�E�6´\��'<f踁M�'T�॰eJ��"L:=C�'�:�i��?�%*�??a��'������ w�����OA�	�]��'w����ˌ�/�*	X�N8.|�
�')�Av�W#�܌+��ׅj)~�x
�'~D0�Y ���	։<V�t��'���	�f�E���r.�!���'�Fb����N�����7x��
�'��@��K9WC��IU�	=u?�%b�'�����1�Xx�T�b�|�H�'6�5�E���+�I�S��d��J�'��Q���T3��P3!��.�``�
�'�u�R!�3����R��7�)��'.>�׎^OYj$B��>]> �P�'a�����8��1V�3J��8�'��C@II���\�w�D=��'˜p���P�B��Q�b�4c�'8ʄh� kA��n�*�:�'t�� #�/`|��w��#D|P��'���#�^M2�CW3����'��Y�"@�$�~|��	o���'GJ)�bmԵ4��ŤX���{�'�ՒǄ�"l��=5�߬����
�'����TaE�	��qcЉ00D��'@�mB6ƙ!�6C�S4��ܢ�'
d\�U�Z���mG2�ܚ�'ضT�ݤd�zҀ�~��H�'�D�2+G�IaмC�bD�p%��'0E���@�ћ� ��i;�٢�'�؉w$R�lrL�po ��}��'��uBf�]J���"��Xx
 ��'���#�(
p����$���P,���':.\�R'T�)�f����G�c@����'J���	�Y3�u��X���3
�'���
�IT�?����,ΏO>�I��'_�1W�d�N-�u���(}.�3�'^�Q���:bS��ZE��*Z��M3�'ˆ(a酫2�8�����/�8���'�|��򀎒|�d4��J�?ڔ�+�'ئ��҇��1� LX!
1�L�
�'�Z��E��66Q���W�4���'mp��r�m�:�B�_�U�D �';������{V�����B�P�hl�	�'g�Tq0���R�cBA��1	�'�p��D�Y�d�bc+B�8��� ��� โ��C<W>b��@�ăY��"O�U�ɒ���(v����MR"O�ܡ� �*��ā4"�H��Y�"OV�#eC]��Xz�a�h��1G"O�`�U�W&�S��Сp�"O���giA�Q��X�xXBP�"OUiTǓ�
)���䮖��6�Y�"O�0Q��L
���B�Z�r1;e"O�<P�L5Mh ��v�V �uc�"O� ��m��ht\Pql�D�ؕ"O��s��L�#Tz�U$!v]�Y��"O�ař ¡��c�$JW�hV"O��iV�%cTY	AG��L�@"On�{�f�s��]
���:�3�"O�4�G(]�i�X��X0.�\��E"O
I�R
��k��ܯ��DkA"OL��S,�-tq��`+�,�#�"O܌S�B٨�`t���7U�Ј��"O@�q��:d��)��A��{�r�jg"O2�)�kF%�I�d�6~� �JR"O
%���M�h�ZPYkXK���B�"O&|��ۨu�l���
�S�p
�"OnĀ��0/��ٰ�ɽn�l��f"O2ĺ�Ѓ5&]X#�ԃd��7"O����О=��Y��'�?<�ȉ2"O,�c#D��6?�t�h��t.<Y��"O�x!Ek�#�b���7q u�"Oz�H�-�>����^W����0"O�`'J��h�4HQ���k�(�d"OR�Q�]�|/�a�$&�}D��sS"Odd�J��:).l�U�ϰn�^�E"O�跦�!�|��ϊu���"On�(�CϹTn� !+J�9U����"Oz�I�16��4�G��F�1"OD�@�G��0([���O0�� "O�ڑ����@a��[�9���"O��k�ʇ�mM���QjU~�0�"O�Q˵f��ؠ��Ot�l��"O��S�Œ;B��ڗd@�G�D{S"Of��@@A"O�����������"O6t2���/�ְ��gH�hk���"O����FL(�nux2f',�м�P"O���تe2Y2��!h�,���"Oؘ�G�?��a��"3� �s�"O��vN@H$:pe/z�P�:�"O��*D&��~NlA#X�T@�@А"O]��O������5�)�"O�=Q�N�gK~ac��F��� 3W"O$�Y��ߥ.�l�!=h�f*�"O�](t���~��� �o*3���S"O>�q&\�9lR���ީ[��
�"O\}����@�6q�!"Ǘ [��H""OvX�BBZ	Z�lmy���uyq"O`lk���ߠ0�E)��� �J%"O��VK�?b��.�|`҈ڂ !�Ǐch�0-�u$@�V1�!�dZ�>/��#'���uf>����8�!�䌅@�n�@���k0���2�!��������<mV��E�)�!��=Q �!��ǐ�XC�$�W[�!�N=��z���DR������!��I�p"&=�3,{�`�O�3~�!�P�J�J��n�<_L�(@��,�!�d��E`��+>�N�	Ů[�W�!�� ���3)yn��`lW�{�\��@"O�ђ��MB@�"���?��p#"O��B��Fo`��f�F-.����"O$M`B�=��ڧ��5
��IaS"OM+��ƏR�"4�Ʀ�+��ye"ObBG�G���D�ԫ[3�:�"O�����9>�Dq�'��0/6�ˣ"O�c�@ێJ���q��@:Qd�9q�"O`��iK,;�rmY�V���+#"O8s�ɒ��fA��E�%*��5��"O�|[��ޏ1�<	;a�Llؼ��"O�s��Q	j�v�a�HQ�c�t��e"O��+'���M����\R�c�"O���A�@�2�Ttiڠ^n�<A�"O���'�$� x`"KZL�E��"O��*�6Z,���3��� Q"OU��Ĩs錱��Yl��|�"OBH��
Z�o�p�r�d,t(bM��'�����J�kX����G�t1V���dq�X��ckg�pZ7#ū;N�ɭ��0��ٟ�d p�R�~n���D��$�'F�f64uP���0�$B�ɱv�Ɣ�A\�_^�qGְN�c���j΅ѥAUwlӤ�^0t���iܘ�?�Qg�?�Ά��i!���'6��c$�WX� ���F�-1��`WD�ҺT��ӻj7�q
w�F,�T�;�-�4��&�[�݈����}�B�	>�1�ܿZ���Q�u��"=��ğ}�8�F��O��HPhC�~D��Pp�8fа�BY�z�2)*Q'RC4�ɩs!-"�ـ��'�P���g®2ViȦ-LF�h��4^�d�U�G�ܰ���.���Ł���u��7hm� ���K'B�xQh1���� �B�(�- �ɡ�lŅ�!�D^�C�.ts�IF�N���� ��Uy�� $m�4@�d���K���9U�A�&`K�)F�M����?��AK��;�җe���kp�6�����ʄo<��y���H����O�h���b��8����n؟DJ��ڦ��M�G����ɞ_��kE��D-?��@��D�e	�����7�����G��r~��B�'g�p"A��z�`�����7�l8�ץqN\�J(�l�n(S�� �zM*g��������01��kgڃVj$�C�@�1�:�n�~��PC���r)"&�\gl���l��?M Ǣ� ~g��KM9�1
$Q�5��x�2,��4��q*�"B!�^�*D��p`��ށ�&U�)����H�L�GI�)`V=���0(C��j�`A�֟�.�b��((gܥ@r�ܺqB���0?1E.w��C���-��dV63����~�.� ����a�O���]Kb=q#��;�ڡ�c��+��qa�1�y�&�::���C1��-f~t�w J ��I�\�Ը����B�ax��߿:�p���0"�>;$�ڸ�p?��U�|��X��^�J���: bĒ_Wƴ �*�-#�C�ɁW���B��E�s-Lܩ��A�t�6�>i�/Y+!qN���$�&k�<���!|�!��\+2����4Q���P�ة�撔����/�~���?2���ȠF���}c*A�Q*��&8�P��S���\��90��&/�ў�2ĩ�����d������u��݆E>�5H�	v�RUpG��?�p�C�_�p�Xg��q��ŐÓ?04�!�V65�mG�_�C*(anZ�G>(����þl�bE$Ox|X�B�?��f.
>h���� 
�H��G�&p�����+$t1!��"�!��^.��Q�#��%��QG(V�����x��Bm��x��+���*l�x���i\�� 2/@v ��9�ıA�8[��r4�º-�^���'Y������;3���J7ʅ���-�R�߃�n���X�q�H��)\ /��9l�-ycz	��'T0�;�%�=0���'�ܩ��/P<���!��U��Ѝ�d�/y����M�?���A(Qz����<Yt̙Kd�<23�9���#=ti�eg\�A��sC��3�49�c7O0��R�$[�9�7��~�� 	D�iT��ФK�3b���	�&��P�削J��Y>z��̋��	!;�P9�-�	
צ�ǃ�8�=CGc� C�	�M����o�<$��4�%Γ�Z�������i���#r
ʁ[�:��%��)N��֝�;���nZ-r�x�9�<XF�J ż� k>r@���'��RE ���lh���
k��<9P��k2,����MGڄ�f/ r�͡6�i�(,�����Ex��0f41 ���Y��EB�C��hO�p�b��C���I�u@ԄS׺�a�>mp$,����N���Cp��j��v��O��̆�I&!��`�`&C<iYR�j��7+>f�I�d6̃�U����	+=�	˪^(5�F�?�K�� �n:d��D^J��e'D�DS�rv(!Ƃ�0B����c�'��1{{������q�"�&%\�DL��U�FB�)� ��PР�.�A�%/i 8�"OZ��qO3�tdЂ$ƭ>��]* "O"���c�8?�\���Еg鎱3q"OP����B1� �1�7x����"O��@3:֮��IЭj��!"O(���HW���`��K��<�D"OܹPR��+;��y���W6z�^�(P"O޶0��.D��5�t1		̝��"O �ӊ�5��47�Ӧj�`��"O�����C"�P1"��(����"O����F�%A�j���ȏ
x�K�"O��Qo
���	�v�b"OVبT	Ҧ]��q����?D�!�"Oڸ��U�uap�{�-B+C���p�"O�]���L�H��M��0W���!"OjMici]ɢ�����aIn��g"O�UH���G3%I�*K7Xj&!Yu"OT��N6�Z ��� �,}���"O^��l��
@�Ђa�uQ�\w"Oh�y�I��1���~�"���"O�=i(I��ls�^�X���"O������Z��e���I�MCd}��"O���`2ِV�[%fM~��1"O��z!(u��\ �aL6$<$��u"O��C��);J��/̶ �g"OHpɅ� "?d��W9�`���]��y2N¹@�TT:f�I��1$K�y���c,84ГL��a�c ڵ�y���g$��y�o�cXJT�2�Ȯ�y���R. "��]�-���:�F��yB���!.!�c�)$�� �W�y"�#,����`�6\���ԥ�0�y� V�K�򡊶���LI:d�T���y���xY���BH�8���!׉���y��T�W���U�O-X�h�j���6�y�U�[]�8�W U_��4sQ�*�y�D��p���bC�d�@�ם�y�f~�:�NUa����JL��y2���k���jb��)i���&EP��y�D�
" >���K׈`}&��ӃB�y��	�=9����\Kt�Z��Ԝ�y�C�n��K 	RK�m@a��0�y��1Ò	��^�R�0�Ӣ��yb�I�>��H��\�L�u-��y2��?;��! N۶_Ƕl!R��*�y��F��م)��L!bT��nV��y'Ý>)��p��+F�d\���9�y���� C0��S��/d�s����yB�=MB(k����&:Nx�wC;�y�غ;������ʠb�7؜�y���2"pswBU
(�\��B 9�y�.�2){Nu��Ǎ�_�lh!qf�y"��?�j��f'�UjmC���y2A�/q�
P�I�E���J�O-�y"�^��|b2(Vx� ��d��yRL�B�j�ʸL7h��eC[��ybh���j(�8�������y�/��>{j��F��(yC�ٿ�yB���V�i�V���k"&�y­^=ڬ�1O� r�B#"��y������`�7<�z�i"j��y��;fP�\�r��$L�^�[с0�y�(R�7�qc��U���б��yR'����ª:QĻ୎�y
� �(h�ț)�L�9ŉE�f��"O	+��>Q�Lу��H&;5\��"O���`�"X�X�S�"׮{,^8Z�"O��@��-�
؅� �\d�a"OҨ�&�&	���*н%�n̠G"OV�2p��p��=Y�oG$��<�#"OJh�ɖ'��3�V�Mrx	�"O�Xi�.\�Id�	d'U�K���"O�e��I�?�)12�0G!3�"O�tJ�/�-O�!�cJ�0��a(�"O�x���߯O�v![Fa�34���j"O�#!@+�8���@JzX�"O����nQ���g&\�0�$�G"O�pZP❊f��A����T*����"OxXu+� ظU��O���kB"Ob�	"��d> �RD&ɉ6R|���"O�����y$� ��EǨZ E)!"O��v�ǿi��l�r$^3O�5��"O�Ip�W7{��8!�X=o0.��2"O�-�[6-rQ�!ˎ7H8=��"O�0�̆�c앨� ��2X�7"O�<R�'�'���c׆��B��c3"OZL�qh]�|%Zܹ&C�M�x��"O��i���@��5� ����"O�a:���*B��j1fSC��!"O2�A��@���ӂ�O����x�"O�y�0���X�(�� ݣ@���"O l*w���/��\k�T��"O(�(s��8=Kf� G�ѷ,��D2�"O�
T�=�4�SƦ� �؉�"O�٩'ʶ^�� �wQ*a�1g"O�H��">9���I6ǜ�ZD�A��"O�$h���]k:����R�!�}G"O@	I���Z�ڵ��I�H%�'"O���+לN_�#�Z9��!"O(��)� -�Uk�Ɍ����"O���ᡜ�@���f�: @���"O�T#ÀܯH{�(k�
�6;P�Ӣ"O<u	w��+"�����C+TR�"�"OV@����Q��Q����4����"OΤ�%��a��z��M�t���	su����,��D��8K#bȕiY��9ߴ=���@�� 4�B� �#����'3 lH��AG�O>�b��1u�p���
��a�3Fh�hCGH7.J��H<E�t��9FJ��xQ������bRІ֜�k�$�d��r�4���S�T=`jv��3"<7��Y�"�@�#v��ff g��T�1+D�L<�OwNݡE%�yD�3�,s�2`�y,άs�0dç٠|
0�D�<�@����y�H�'z��0F�阧��5#ΪV(���� {�r���=O�b��ȁ]1O?��.�J���񂈖�.�+[�{�PŠ��,�)��H �鎶aO6Q�vÔ�bv~%Ʉ �1O|
5�O$��jgA�+1��}�0BP��4��y"b4�6��U��.v6����43�z�����>�5�&.��Z�B�_Y5ノ�j�@M��Z�"~*���;zJP	[(r�lv/r�<�An]�n�\� ��"ao�]�B)Sj�<Q0L��u����
V9t�����p�<�Ʈ�
pj�� �C38���ӧ$j�<���55G(�	�#+pb�S��c�<䉑5N��P0.�'�H\�  b�'�x�gT�5?��P@�D	1����~�<��d�l�jp��/��D㕨�l�<ɂ@T�zY�Cr��A2�<���\�<y�*C�R����U��d8��Q�<��
Q���e_�����*
N�<`H
��H�$@G-+���ˇK�Q�<� ^�	���|��D@N�l�̵�"O*ؚ��J8
�����J�IRE"O�Q���*��T:���*K:8���"Orp�g�F({��}�se�+)���K�"O>�j3�D;�����M��ec�"O�a���A�عh�b�1vZ��D"O��G͜��@Ȳ!jU@Yp"O���$E#xx�p`��a�|(�"O>x�F���:�^L��nP�bȻd"O0���l��4w���!�W$�:dY�"O��sSCܔw�$ԻP�R���E"O��j�`��w�)s���
�<q%"O� Qc.�5M�6�ru@=y:(z�"O* ZwkU�5gd"�G
��H��"Oz���a_8�{�.�G���jc"O���ō@�\-����mV�+��B�"O,�c���"��a���Z+`���"OvIQG
ܣA�����G��F�+"OJӣ�)�F$b�(�ik�f"O T��KK�{H�=���Vsa.\��"O�� ���B�Sfƚ�	a�|;"Oh0�F�VA���/D�HF"Oh�9UK �w�e��""D�ّ�"On�)��)��xZ2���+�8�y��˧&ƺ����?W �9�@��y�>��DX�D�9�P �.�y͏:W���Iq�t��"�y.�;;jp�q��ۦz�~hYE$Ӕ�y	R� 1�EQ`��w7��k���y���7�$�re�ݤ7q�s��� �yR�L�������&a
	��Γ��y�@�U�V�I`��y����@-��y��I&ʘ��ct��!@����y�.W0u�TcH�}j,
@�Y��y�+�66hh��2��w��Q9��D)�y�o�/vM4$y�%Ǆa}B�3�����yrχ�~�z���l�0*@`�i�jQ��y�ƌ?y�ډ2t!L�HH�P'J�y�lA�>u$����<��X��V?�y2��!!^"� �k�|z7���ybl�n�i���90��ˠ�y�a��,�N,�#��C�(�w嚜�yB�R�(��Ѣ&?�2��ᗺ�y�O�
ws�X�B�7p|�`�:�yr	/z=:�@C�8����?�y��\�g�\���½l���@���y����Dt�R��<;�]z IW��y� 	�%;�m��H�>��g^��y��wx�P�f���� �����y�Δ=u��٩� ��d����U��y�b�g�`�C�ǁ9����y���&j���@��>2������"�y�AO�e2��f �8�*d������yr�I�����06�B����yr��t��&�A�&���r+_��y"�	��1c���h�p%�򡘫�yB�ƜX!��V�P*hT�A�X��y�&�	h�m�D&�����s�ŗ�y� @()�tt@�D
q9Reprh�y���Qڍ��#S�8٠���y2n�V, ١4��a�*B��#�y����s��kA�^&,��El�,�y� �G��ˢ��D�H�����yb�80ll����ӄ?�R\�t���y
� ��Xb-؏K�}�1FNIo�]"O��ْ-G���O-Tt��a�"O2�O�fu�i�#d].��%z"O����L�!s�x�कG&��a"O�${�B�,�%���g��Y�"O�ij�	߸f�-�1b��o�P4�"O �)R'�RZ5�[)8�(��#�O�<�b헹lT�Fˎ�7��1C���K�<֥M)'�`E/���� 1JN}�ȓH҈Ȳ dԩr�D��#.I)$Fd��9�������'�}
c'��-D|���3Tv��cF�0sZ>H�6O�%M��|�ȓWXP���B%]f䩥dơY`<����X��MC*]sc��AG��ȓ!4���D�y�`Ȃ��@mk�ȓr����s.��G���A�!d�ȇ�	���'��HI@7��P?�Ʉ�A!��B9ꄠ!0O	,Xn���i��US���g�h��iC l�ʡ�ȓ^������3���y�o9iи�ȓT�R�2���r�V���*�z��@�ȓ�h��㟃-']i6B���L�ȓS~�)���nC �P5 ּC4\0�ȓN�R{�G�';˔�2��M�'�����o�X�p(O'%z$c��d~���ȓ�a9��ދr͜���c�@Їȓ8$�@sT
X�!��{`��
hI�0�ȓ+�,���.$}&,�T���b}��*�jq3t�&{c��ć+a �ȓS<Y)�$Z>~�B�Pf_�4t�u�ȓ�he+�I�"������M���i�ȓZ�h�"'@J�3B%��XB���ȓlI�j-l�L�gh_�Z~H�ȓ.���*箄��2h���\(_Pp��P4��0�b��"Ӽ��%��*���ȓ-����I�p��i0)S�T�V�ȓ#md\su�*Hq�$	:7~|���j�8gF_yz�B2M�:*�\�ȓ3��M@D�w�V����ĸ̠�ȓ}��xC�Mœ5�2�A#k�77����ȓ*�:qSI���<��a Ը
���ȓlKDe����i ����*��ȓ.���jH׸hN4J7@M�dx^���qJ(����_�Kt��喨"��ȓ!dT*�ΆF�JU1- 31L�ȓ��+��iY򁃃a�;�X��ȓA��DAc�.^�=���TJ~A��d�ëA�w��\Y��+��S+@4�g��%9�ꥋª�"|g\��ȓ/rjp�F���"`|[`f�A�"�ȓ��h��� ����a��6(5�ȓ�>�!�'�5%�r\ q�@l7@q�ȓZ# L��ʹb
�<��^�i�t�ȓA�&MC���7u+,8���ג�3D�x{R�P�Ep��^�I޾��s�2D��`��7?��&^���B��2D�6�(3�ؔ1#��=	h4,�䥟Y�<��-S *���d�Ӑa����X�<� ��3�.q�*C)���i�JW�<QUǏ�F^	�

`B)P�<�F`�7r0� v%���hlҧMGO�<���7�H�B��û0w0x�H�<Q$c�$���6��<9d��!�M_�<��U�3|&M�dN|p0�'r�<� t�"�OL�uѰ��!�>���XT"O��$C�/NY�q%]�/��AJ"O��cfɖh_�+�-Ұ1qN��"Ov|2��2}�N��5C�`RIh�"O�L��'v8�Y��	a@l}��"O�(����!U���@W�j'�M2q"OF��#��)Q��J��U� �$��"O<]�K��5JP�n�=Tֱ��"O����:Kw�0���yi����"O-��+��U���&3dp���"O.X"H����F�*Q`�"O ��pG*n�
��L%1�b"O���5!����lbƆ?#�H�"ObX��6�:��Ԋg3�H�"O(��K��qド�6f �9�"O}�'��,"�0�s�B�7]	Q��"O���<;��P�H����"O���Ü��@��^�.�$Y�s"O� ��d�*V ?(��\�u"O��K�$��\��SB�"aN>)�"O�� �!��qL��u�q7�T��"On���(� jà�Y ]�e#����"O��s�K�g���bcH%F�ҳ"O�5[?;�4�ҒM��Q%����"O�dBSeŧA��z$C��Lr(�z1"Oh�y�	�-{�"�@�[�1��"O���!���s�N}�d�{Q3�"O�	1ǌ�7a�҆�W>P�F)P"O��5��%:��8�b������`"O�I�eo�%I�r�q��*���
�"O���,�&h�|����5R�$iC�"O��R��\H�(����۟����$"O�#R+Qc�����S�^�␡5"Ot���+ۯO6� @
����k�&�y�F�O�~p"da�?L��G/J��y����AO�qgKr,X��"љ�yRO� "��	&a�g.~E�1���y�`��Q��q i�03L!�;�yǍ�v����1g}k�I�y��^���@�0�L ��
2�y���'g�as#A+/��\��gۻ�y�U+	x�u���́PA�1zW���y�Ԩ.�}��G�}�DH��I�y���k�0<I��C�l6��T.�yÚ�DŖ�)�*��L��"�C�y�OɆs�y��N�?�9Rd���y�IѢL!�pp@��`�FK�4�yB��V
ٺ�6��\�VgK#�y""�r��� �)	�}ZD��%�Z�y���lR��tGrd#�&��ybc��0�k7I�\��R����yү<6[��� T���@ �y���$���g��K�%���yB��L:<=����a�7Ŷ�y"o�.P-V�2!޼���VHY"�y2����6H1�g�#	�d�ِ���y2	L1)�!2V	�-T���$֌�y��J�zp����q@��I��T��yR�µkh���M.9j�� ��P��y���
�0��� ��E�|9��M�?�y"��͐���ǆ-	��` ]8�yBL�!
2�qÅT�ʕ�0�Q��ybL!p��@JrĕW�` F��y��+^�bX� ��J��xx����y
� 8P��'a�<���^+#�pi �"OD��V(T���)��Tw����"OL��!�ۧm<�|0������7"O�=x�~#^@�҇J�S�<Y�"OV�ҢD��>�L�3&ɲ�l�)�"O�!ST�)d��5�b��={(l!�"OU�d 
  �?D���2,ѿc'P�f�P95qim+D��+�㋅_dRH�@�E�ڜs�M*D�� Ύ	B:a�dI�<����`2D��³�
^�ų��̛f����ɯ<q� }8�4cwХ=m�P:G$M�����-,D��1�ɁT*(�#��-wX�	�
8D�(S7
��)7�Y��(�m��j� 5D��1U���S2 ۇ'/P�d$�P2D�h�3��Im����ȗ}R�V�1�OA��O���UBG �Du�)D�}R.�!�"OK��~*F���ƞ|'�X1�"O�qXq-�?s����-{�0Q�@"OA�R�І|,J7KMs��|��"O:���4$��iڢ�Ҿa�P�t"O�I@�(].Eb88x��
�LP�+�퉩��~ꑢ�}`�8�p`N�u��=�Ԩ�y�<�"JǨB+@Ց����Z��` Sa�<Qb��-a�:=#�@�au�<ɵK�r�*ـ,/��k�s�<)1�� z������&}�\`)�?T��$�O?/zF�U�
>�2�O	U�)�'?���f�01�x(�������@��'�MB���F��j����H���b�'a"쐲���AG�4�F�-,��q�'���'�4ΰY6LM�ؘC�'�:�h���� �2c�Z�A(.9i�'\:��M�?5�p��k·b�D��&��r#�I�?��Un��	;Й9!`�̟���X�?���h�.��2ņ�@
�j�+W".x��5Jv��蟄��@����fË6`�c$ړȬͧB�,��Έ�C��z��@=|{b�G|��1��iqeL!an����iO�MuN�A�떦x��H�'�ֲc�������	ϊ������t���'�1�x�
!��f�(��98f$�"_����	��0�1�/A�#ZM�cg �������wy���"���/HJ9^�8MK���$V�74$���Op��|B�o�	�?���C�s �� �2l�%ԣ6
�����9���	>C�'!($���+��b>��$��/��Cο+U��(g��X���:d��A��,��dkL�0��9��"�S�r� Ly�"��s��³E�]�`�	F/r���O�S�SN~�� ͪy�Ą��s��a��@�y�A�>j2���ag�@צG��hO\�G�T��c�
 zT�U�R!@b2NX�I�2�'02J������'�R�'�R�O��kʼ6P���ƚ��n|�F�V�0vd|���-&
���K<yۦ�K1�?#<�v��4y�^�k��g8B���@'Xۨ��jۦY�f�FB�o���O�M��J���D
�Q��&f��l����84��ɡM�z��O�=��'A.U)�&�o��y
��=�HԚ�'ް��-7|��SK���Ĺ��b.���Sɟ��'� ���M�gM��K1X!wO��ʔO]��Vv�'���'�B�OL��'j�I�� ��x'�w唨h�^Yߤ]{�V1���:h��$���'��X0Bءw�,<���ۆ_ �UK���j!�Ƒ_�dɉvdX�f��q���0�O�Q��'� �2'hS����
ݼ|$�I��'�ў�F|�iΧ:�RYc��I�LY�PǤ�y2�>~`^L3�D�J����+�
��$KĦQ�I[yR�� ]I"b?�+��S�[����&��6xa�IFy�'���'	jJ���->l<9�o��vR�f��#��I�e|�a`��̅�� Ё�@�'�l� CJB�;�v�3IQg��Z��g�I��\�+rԭkM� (��l>�
A��	ߟ�|��oZ�SXԌB-N�p<r p� �sy�'0yB�΀z��٢r���kH�����ɠDT��c�ǻ
Z����d�<�3�
!�?���$�|����?��"�I	����Y}�����?��ҳe����A�a�&�a���ug<#}�q��	f]жJσ��c�T�<"星ZŴ�y�@��
��bB^�>j�>}a2/?7{��:��b�sפu��k���O�d<?%?�姀 &TZ�튒N��Pr��gcThC"O��ȗ���I
0PI'�27�C��ɬ�ȟ�=��^,G$����I�Cϸ��1��O��u�c���?Y��?�)O��Ȟ5e ��#wU �j�']�]pT\XҢN!8!����ݳ5�W�?��}��ٗy��j�c�,������D4F��%n\2�1)m�n)�ϟְ�>����G� H�4�ΚB�J�9u�	[~�	��?I��hO��/h`�x��MKIf��R��Y��C�I
�a���-w'@̀�U������I�����'=�ɌKk�ۆ�M#}O$����݃F���3G`��t��ϟ���xy��$�֚#�h�k"nV�r@�d����kc��
�@
Ҫ�U�A�iP4�ۥ@u�'T<�٥�� -�tQ�dE�9T�य�?T�N}�IÁ?%����e	�z��#?D������HَmD>�R������)�蟼F{��ɧW�>���oQ [Р��H�"7VRC�*���r˗�!�vUaahM09x˓ 5���'v�I�&"���L�$s>�S��4q���+W84�R�r��Oի���Of�$�O�*Ӥ��-\B}�w� �Nm�B	}>��AcJ@2�ŚP�,���[j/�2U���N¯k3�,kA��G��Q���w|��XwX�z�N�#�'W- yڔ�� �S�'��r���?9��d��ڈ��Â�t�*|��O��$?�O�ax(�=d z��\�#�n���'p��h^����J�X��h�䎢5�@�'l��'�R�'�W>-�	�|:碀�%��� ��D[� Ky�Ž�'Jў���&�#z���YS�C�>�vm�0'"���O0b?��ՌWc���C�ܡo�.5JEN ?i7�O<1B��>��yb`��z�0��ă��E6	� L�-C���d�N����-}�9�!~����H�Z�ڶ��":��O�$�x?��9O�t���Ē�t�S=|��A�#�x��If�O�'9l�Y����XĔ��4f�h���R�'4pJ�lQ2�>���&T�"ȧ!T6�2"�	.,m���(���OL�O�t�ԕ>1��i�ԝ�&��&���q��c1B�i+O�`k��>�&�S(!�4��B�ǣ��ܓ7MQ���b�'2��I���<��o�4�?a��M^B!cgԋd�܈��d�2rP; 4}R�Ȭ�����H�N!��ٸ?L��!hP�1S��z��'ʄ!�B�ȅ��9O����O~���3[�e�Ї��i*�9��'+�m�O���O2�$�O�b>�9��H�0�U[� J$nfJ%�'D����F��0N�u0Fɺ{.M��aeӤ��.�d�J��'a�Q>7-ҵA{�h�e-�4B؝I�h�A�Idy��'�2�T?{���:D���Woű�u�F�"D�`��
�G�<-Jbd�R��%Qg�?ғ�p<�#O�$�̸i6�ˀcC�h���`�<��i�2D�L�����;PFz�M�_�<	eݶ2B��W�ɮS�X�4l@�<Q��4> �Ad�P.k]	SԊ�x�<�e�ݎwt�"�"�B��2F�|�<qC+�|x��Q�l+ܨ*t�z�<�4���}0�)�g�D\�b1 �t�<��&�T���T/ �U��T��&s�<�CÉj �l�@��	R�Rp�'T��Š	�F��#��-�,����gWv�>��BBd��H�"O¸"�ݨ(xVl���ѵUS��s��d��t��:���r���)AM�O�~��B�=���ӑ*I�`�z]�ơ���F���H�(����F+Բc �XY �YJ�X/D�TȪ��E���3��% 4O�2?�jT���T<خ(�t��e�$I�E�=~�f�a�l��D���E��'1dr���f��W�^�.�8��޶A��&��='9��QTg�5h�2�� �[.8�:�$�O�A����O�c��gy��&�^L����,8(��'�*��X6��Ex��ĩ
�1]��[$��!B
�B�-���ēF��I���S�ZD"��/�j#\Xs��
9d�5�ȓ�F����-|(ubf����I���(O�(qK5�����Ö�4!�5 ��	�M����?9��]�؛ nݿ�?!��?Y���Y a#E<�Ԣ%� ��{"D����'��9Z	˓.���������񁦁�s��>Q�o^X����IG�q����P�˾O��Mhp-ʩK��'��MX�S�g�I0{��1����td�$���`B�ɢ��ly��1ۚ����-R)��'�H"=�'���h�r)ڭ9��X�!��ur$�Q�P�*���',�'��z�E��ɟ�̧`"z|X�#P;u*���!��ೖ$�^<a!� �U�"��G���x�O�F���sS�SL<�Q�QPs�a�C�
B��@҉Y2�	�p?!f�]�z= '`7��q+FC�<y�$�i�̢T�ʌB��i���gܓ^$���|�dD8�J6m�O�6�
!z ��h�7d�)�%h̕{�l9�	֟�k�KX��t���|�$��� &�P`	��� ,+���p���1,O<�9���1�f]c�h9E9n�j�7;|ay�l��?��>����5e�4l��$1��L"�p�<!���W�n��RbL�.�Z�a��i(<1$�ݠ'꺙������-�w���V�4rJ>)����?!��?�*�"i0�h�"��AEV�8,ATc�6<y��!R����ɖgZ����q�S�,O�h�@�cR����T[�x��x����O��dm�%�)�D!��@A�rC�x2 ���?iї|���/��c��0)@�K`��ڀ���y�o�(s"��� .�-��8�Վ̐�p<q��;n�"�0C��?�hP���/J32��il��'����w��4���'t��'��;c!��k��M�K�<����]�"�3�$ݠk�ayRoѤA&4�f蕤 �(p�W��'A����Z�����*,��6o�Bq���'�d7o���L<!@[��V ����x��,��Fd�<��f-,en1U�ڑ.HLxGnd�D�J�����xR��)M�x��ШLv�KwM\N83�
�&��$�O����O���O��t>J��X bb_
C�hY��Bl�B��#o��#�'�~��YZ�!�..x�1#�&���`<wʡ3^�l�#�ѵ9I��Ǡ�O�����e��,aPLY7:� ��D�C�0��-�@@�W���Ғ�ѐ㞔�ش��>�VTu�i'��i9��*���/P�;����s�����#�O�����md�D�O��'{�@��ݖE��I�o)��4��*NN��x���3�d��N�c���b��SI�yK���qRݫ���.#��ܢ��ɿc��HR�'h~��\�d�rT�1��&�0��Ec��B�j���\4�SbJ�%`��(��lG�d�Qe�M���&���ʇ�ktHE"ܤ��Sߠ-XU�i��'��S�p�<�o((�&�h��0Df�����D*ȁ����?�1�K�/��H�%���i����	�~���jQ֠h� �HI8��+�x��)�Zpʠk[4E��P�+
'����}��X�Q�МPlO�g�:(���U�hˉ'��u`��r�ɧ�O���Ӳ�_�7���K���"���@�':���֩¥ej*)����
e;����uhQ�\��*TF�%@��ޤ񬀒��ӵHX��ğ8��Ɵh��韔�Iڟ(�������Y�z�$,Z/b��9`΂����t�"'�z�i�8����O���a�w~��FQ�I17-����	��.U&�1�G��@�r��p�*��XB�|0Z��OL�&dd����·Z]�}9�l�22�8r��^͛V*������&�D�1
�\�gy���b=Q ��xJ�+�����m�S V_y��	��x1��|��ЫuX���E���n��~"�'>�7��O�ʓ�?I�'�?�O��:e�׈��$P'gI=����'-�pwpa�.��������	��u��'u��'�L@d�׻v�u� ��e�& ��C��v�=c��S��pu�N�Q�eD~rH��.�x(tK�A�����,��<���cc���t)L�y���{�&~Ӗ�hc��1�ȓO��@��) �x����l�l��s6T�B�o�mZ�d�'���']�'�X9C���#f��:Ș5X��S,�Ob���O�Ԫt�:���?a�I馹-]����&݅7��8"��?g� �'rwӒ�d�<a�H��d����'q�&D�T&�m�G�[;K֬�FA�+B����O-ӷM�O�d�O�A��ݺT�d���0O$7�$Wc��j]
���	���Ņ剀�h��. f2U��D�1���e��lžE��cV�"~�Ƀm,O�m+��'#�7��_?Yхυ:�h��A��38��шC.Ho?���?)���$��-&��!�C�'`��y�%�9Tf��O���W&>���Ͽ/ʂX�K]`���#����'�B�l��D�O�'e��(�4W�����ԈO��0V�6.T�Mr�'*�o��W����Q�׹e�b6m�O�˧��)@�a�!���ζQ�� #�	�
��'���8�
JFؑ����2;�h�� )�=k�4��Ȇ�1d O޼iP\�8	J|,O��]�C�d�j�J�m�D��F	�:�'�2�'*�П����`�Ɂ���ˆ�#<v�Q���+z��ũ�@�I�{�T�i>5��O���Mca$L�`�,�r�N�
C�0�)�E�!��6��O��$�O^dA�BH�l�����O����O��He!ԩ�5��\[,���%8V\PW�Pi#�lX���>(�HtAb�(��%(���8��'C�L�q'I�7U,���E�(O
X�3FF#L�	P��v�8����:-q�D��F�Ƽ� ��j��Ů�(���Ɲ30�LTQ�`�ܟ��'g�����|r���'���@do΢$���)� 8!�2��
�'*FYB�"W;�-�cb��.!IJ����4�t���>)���l.4C�Ԝ,����K�b�$�5Y�"!"�'b�'/֝ʟ��I�|zb��-��L��A�RҭZ˚�|aL����� !�P1F�D�����{p �tH�;|�Á&܎ET����a@�{Ό�1g[ *qY}� �w�6'�H�cU��$j7��A�c�&�<0������l8��g�+��UA��� u��yG氇ȓ2D�D��n��@��W��y�=q'�i��'j1ɠnfӰ��f�*���*F'�����	-qJ��ǣ�Ɵ����Yº���ޟ�ͧ�dȚ%N�7'Q�U�'�B�B�:4�K�@�2��D�	˓+��i����3�5��^Gx�8i�f�u���i��`]����Êo
�`��d�"cbN:}� 2	]���u�Q�ĥ8w���yҤ �&��d�7���#0\��Px��Rk���+���/Z,��aRÕ�T$v��|b�:F&t7M�Od��|��ܶ�M��� �8��I�l���ݩ6\&_t�'ۨ`Ђ�'"1O�<q�O4V��	��dW5x0Z(�e�w�	?]��"<�~��0Jd<�u�1�j���l�v�`^��r�)�ӵ���B��2�RIb'��~�|C�(Y2:#��[��!Zg �9&\��Ss�'�r����	����DL��a����'��'Zay� v߼T��[1t�I
�j���y2`�-K��D�3�64��oI
�y"��k��	&/@�,�X�j��L��yB��eI��BA	����`���7�y�gg$4��F�P3����
 �y2��&UA����m@Z��QKΎ�y*��JO�i ��V�)�{����y�ޥo�UF��)��u	�Ǌ=�y�·:�4�ȁ��n�i��Ԧ�y�͘�-]R�R���>���$�yg4������)M5�u`��0�y"�Q�EYS��7L���)ރ�yb#�Ouhɇl��NZ�l���V��yˏ�	j4@ĉʉG;��b')���y�É"���҂@�7&��w�3�y��L6�D}ȗ��1����Y�y�͏=�P��D�w踹�f���y�ش'	� �ֽ{A����N��yrM�-���Ǔ� ����D�R�yB��8V�H\Av���{2�,���yrB��j0 9�gѭgkP9£N�)�y�@�>[���e
�.a��9í��y2�'QK��;tF՞)E��bRM_�y2l!g`ֽR
Ӑ/z����y�ჽ �p��ݨ>,0��S�y2��)8�|�K���b��!6%[$�yr�N?_���ӪUb��%����?�yR�M.�ZD ��+Z� �١���yr��)�9�a�C$Y����	ϛ�y�爃*h���2��܂����y�HEL�BXQ�΀�~&�d���y2�֪Ƽ:4C��>Y��I�y�X@�l1g��w���P,��yb�0J$��J��q|�	�aኊ�y��5~�p!�[8�ic����y�$כ-j�t�c'��9V�%X�&�y��r��8�����8�\�'=4�X���*P��d��>^�@
�'V��EVdHmۃ�T <"����'�� )��ؠА��mZ6!"1��'���Z W�1�I�B&ݖc9�`Z�'�ꕂ�oL�T�8\�R(F�d:(J�'�pZçT7Z��9���(���H��� ��0��B�ah1vc�8�P5�"O�ePl	u��Yiq��\�DP�d"OLtH�%*w�� �fAL�[\�j0"O��ċ�3<O<�Q����x�X�"O�!3�
(��G&�/n
��U"O�XwNQ2��!�S�S���Hq�"OH���,Ί�� "U <UsL���"O�����P8%���e��Z�̨2�"O����g�S������*ea�R"O]�Db�m�,��F�C;QB,�"O8�����r`�bփ� /�l�!�"O,�;���&'��`T��!s���"O�$a[�E�1,�s3x��P�|M!�ȴK�Hi �ˇI�Q��R5M!�$� G�P�/ҢR@� �� )I!�ط,嬀9D��#���1�X�Py��O73>����`�q��*$j���y�e֊I8l�2`��&]Z��Ǆ�y�P=	���q��2
��$:s����yG�_V��p�M7�l0�#�N�<�E/�ofD8D!Hr��A�u��Y�<�G�ƅ3ѐ�3��-{���T�<�2��9+��0�b�6~פ��b��T�<���]�����q'�6N�ZaKMP�<��U�� rtB'z�bA��a�N�<)�!�T8~�KP�F�ȅ �C�<��1q>+�Jė' ��e�{�<�eG��?�z�fR�ls��[��w�<i�a�qw�(�QmՍu��ų I�o�<�HO�Q���2�>cB�K�Hk�<�VܟiR��$i�Z��P3��~�<q ���&��d�"G�_����W@�w�<qrmĨ>�M@���;?h�u�礟\�<1�+9+��!�K;`요����W�<9͒4
;P͡�a�56�T�p�^�<)4d��[�V�qU/E/~�:\{GM�Y�<�po�&HR�	�Kp���E.�J�<aA̳`��P���*BF�y"��o�<�#�P����m͌J���yBGF�<��l�,Y��#�2���"	{�<yE�ݿWw6����&���b��w�<�c�O:kw^\�w-��R(���/�p�<a��-(�t���/
Pv]�Ek�p�<���Ff�s�ֺ,E� �� T�<I�L�-���qI7t��9���S�<9mļ
�@b�K4/$.Y���N�<	���T&a8S��"�~(A��Vr�<I��^�9���08�V� �"�V�<)�͌- �n\b��)H�j���iS�<���̸^]0�&V.G��Ӵ O�<y3B����1#�d��L�G�<��� [���Ӈ�C+$��-NC�<Q"�<�0s7 ܷ*���b��G}�<��(̣j.f�K��|��d�v�<��خJ�.�	 $�,�,j��@q�<91%2r��YD�=��xq�
D�<A3. i�H�
v��|��&GB�<Q�n5A��� WHP�p��	Z�<٥

�b�]C�� 8غ͐��W�<�3_�_:�}����"i �����S�<	p�$?x!�RD�(�>%�2��S�<��j5l��4
��0G���hIv�<)�hX#�
��!)˵r�L}h`�W�<I��ބ')� ���/��96�T�<� fa��&/\�=��JX�qXn�@"O�YHq&�JV���^C>x��"OTò�>�L ���D@�r!��"OД{�T�ʜH&�F�G��M�&"OR�k`�G�	rgF��T�s"OH k¢�`x5&�+ڼ �"OxA����q\����-%�L�"O>���Z�Cb�0U��K��5�f"Ob; � �!�xL#v�ѩܤ=:u"ORd��l��n1��y��SL�b��"O�P;���N���aA��G��)hr"O:����ЖI?��0b�ț����"O�*3�(r�z}s�����i�p"O��H�W�<ے��zs
(��"O�	�$f�
4f,E��ǖ�q�$�p"Oi�1.��X3�S 1U8��"OT�J���9�ne�ń��BK��"O��
ף�u|$��w�E-'�8)a�"O���`B]N� �p�G��}�^`�Q"O<$���] �
�B1��?r�,9T"Oܤ�do�K��`#eדdS�P��"O��fO�-&@�%���Z,p'�,;�"Ol���K�<�B�25�Wl(m0�"OL �5ʆ�D���Aπ|aZp�"O��zF��R>X�V 	 "M| �Q"OTň��#0!��" 6e�h�K�"O��H�y����'NM�A�ZIR�"O��I��5j���H�L��"O��pS��}�|)m��p�r�Id"O,J��	(HB��Ҝ|�����"O�dp�.9F� ��A��66q84�"O�t1��F&�H�#��|��`�#"O�yzw��6��t�V��A��"Ol!�6��#aD�p��P�V�!�"O��mY�t�*]�/Wl���"O�=�$�P�`6�,��p�NR�?)!�$�  �h���ňc��E�̓!�D�	*m�X���_�-���N�"�!�$C�c>���4iDu�VC�7T!��
�6BJ�F�=V2��b!./"!��M*y�Z\�ë؍=�f���O��q!��4e�D�i��@Z�,��dz�!�DɊ$�6�y,��"54���M7{�!��?b
�`Ə=��Y��A�,�!��7h1�員ޢ�!k�\�!�Ē5-d��u)�(��hٖ��J��dZ&���vLO���cN�y�.W,X$��Z�;�OF-
�����'�t�H֏ѝC)�9J1�&we���'�N��%ϗd$T)���}�A��'�b��Cu����FA�p�lC�'u��#$�:����M
j�(���'�	!� �NMjuqWD��u�$I��'�DX���81�	�VN	�sw�D��'�QX�l[7/c^P3Cd����'�����M>R�p5��	^`M:���'x�`̊t�h�E�ܿW��Q�'F�e��&Hd�jgj�S�v�!	�'<�I���J�<Y^�R���L����'>rm����-7G�aq���z>�Q�'� �r� 3r��L3��˄mK*��'C��ig%� �zABV��8j�����'q�Mb�L
�XM+��WY�FQ��'ڈ}�vjV�Lw�@Qt�
V0��� �,3�`�/�ⵈub	1u>���"O�ᵆJ�e	��C��'%��ie"O�a�'�U�)��5 ''�d'��{"OT-KDEDl�]ɠƏ�a��U�1"O�9O	zZ4��ê�B�1�"O$���䓋Lj%s��� F�~:"O�ѓ�"O�1���Ek�W� �g"O�QP��%0���"�*K�[نc�"O����ę$TL��i͡>Ð���"O�Y�c$����.��c�Hq�"O������_�2աȊ&�lc4"O�8PШ�(�r܀Ҭ g���"O΅P��^Zc�T���j �YҰ"O���U-��T�8��e�[�����"OR	�w��KW4�H�8�,P��"O��y1hW�\T����S�.��H"O�I��*P�T�c����p��""OF��GM�sڬ�����(�0g"O��9��R��H̚D��#]����Q"O�� �� $�zAע���HIu"O>5�͘)Z��	S��x���"O>	i�OK|2�A�r�T�6N���"O�$�GM�\��XD���O���C�"OF ��M�"V9<�y1.D�2�H #�"O�`�1J>�0�&dX$=�D��`"Oʼ��Ag��� �B>v�E�q"O�d��$F*X|&�qE�Qo��d)A/⤃�c�wd���.$<O\-�!��J�ܴ���8 ����"O� ���#z��!��@PD�'"O�PAP,��f�S��9_L.l�&"O�H�ue�[*B�p���S��#"O�� ��]
u���"��	��L�"O���p�$���b� F���3"O|�!��� �b� w��r'"O2��@���&v��Q��ؕe�v-J"O ��a�xҮ��%��;Kf�M
b"O4hp��&=F�
��*j�h�"O Q���ɓ{5YPƑ1Lj
�(�"On�����-}�=��[Sj�:"Or�3uFځ�[�4	��A��"O�5���̓�Ԁ#�KZ�`����"O����["Uk���KG1+���#�"OT�5��e��xRj�#w���1�"OfЊ���M��A2��N�l��"O�%���W��h@qh��_�&Xs$"O��Շ��������:~��a�""O�*f�R�~*�h)c��$q�X��q"O�es�#]���y��3?. aT"O�ds�ٕ��Ѥ�l� �!"O�@�0��5��bRO��b"O( �mR�Olt1 �1�F���"Oʕ��\�D����v��	���c�"OV��WC��p Xtz!�_�����"O�a�UĄ�A�D�#�$c��DI�"O�Ӡ�T�8oL1!5�M�^��*�!���(?��WNF�)����l7!���T��<�Eo~�܄�ԁD�="!��+�Դ���_@��h�c��!�d�2�`��b>���!#��:m!��=u�A�ǌ�#�2�8f��Fe!�$@:M	�4LZ>vS:]{4��6Ia!�/���#��ÏG$tKE/}Z!�D�-ghHq�ӫ
��qiC)��4H!�d^-�2y�Ă�� z!��-n�!�� ����:�0� ���&�V A�"O�kҋ�~HqQ�W�f��Isf"O4I�a A��y�ә}�$��"O�!���^-r��kԨM��ye"Oe�t!d2���
�'-�Rݹ�"O��r�C�%:�CT&/��trG"O�=��DS�=
T�H6q���a�"OhiBWI� W������>�;"O���cD�T`�$�.C!�"O2�j� Y�4�Q��kO�\$q{f"O��nɤ	�B	�p$@�}�|�2"O��""*W0�W�'��<��"O���4n��S��� �d���u�"O0=��E�,��EbWD	�ȡ4"O�,pl "�]� �;7�:��A"O>��Z�*������c���"OL����>��	!���o`6A(%"O��2���{�x��c��KW����"Ol�BG茟��}��gL6	q�q�"OD�s�̙;�T�J7a�3"O
0��
8�T[��V0OzP�"Oԁ��G��7���ݯ^]
�+C"O�C�Oʂ;zD@�R Q`�\�$"O��JBj�:X�Ĥ
!@�-S�h|��"O��v/֒$�e���ye
�O�<���)y<��Ӈn}��)*��r�<�PC�3
1P�߷l¤����L�<a5!H2L��<a$�18 �|��d `�<�S$�4=�V)�7��(8��i2`L@�<�����\?�H�DV
-����P(�@�<)#b�
^����޿Z�Ʊ)�S�<"��o?��Ս"k�t��&�w�<���ǲ�(�b��ܺ?"��fȓp�<ق�ג5������]�)�B�L�<y����x�@��-]|%��~�<4-I*\����3Jɔ|�x��Zy�<Q���0�Q&*Η8b��o[}�<�gL�X$��Eqa�&��X`x���]�Z�!��2�x���غ�j,�ȓ�8�˃�#�j�+ϯG5�Ԅ�	H�2�@�4�X�P�G-B�j@�ȓ6�L�5.]�_��q �⚍a�(���;�~1���2�a�&��1����ȓR�NM�D�"\��Y�G��J��L�ȓ�j��a�N�%��$��ŉ�c�\���&�$��"	��aAr��4��P�8s���(zG�p"�Ɛ�y�r=�ȓHҊ}�a���3)Z�0B�+3<H�ȓr��aj�o��ܐ<�d��5mȅȓ%t
�H�LC�3��)�tl��G}8L�ȓ${4�I��� ���Rs`�B͛o�<�3@��DT���vDKtF
I	��o�<�U���Z�D;ס�-Ϣ	q��Q�<1V
_=l� I���؜1���qQ�n�<���b�F�2�n��KY*͓"��f�<�� )r*<����6@���@i^f�<��ݟD�ld��H*�������x�< �a��=I��f�ǰdrb1�ȓ	�`Iito�5Hh0Ǌ<x���=��5��HHDՁb��Y+:I�ȓLby���(B`�Y�1_�x��ȓ �L8� ��A��Q�(SJ�|��L��'4.��U��'�j��ȓx��(���"c���g���E?L���S�? R� c 'zjY�a.Q=r.���"Of�d�?��4�w���k�J9SE"O��`��C�a���z�mF��!W"O�����8���"EK_-v8��&"O�tC�@�bδ9+ Ԣ;l�ij�"O��0���ܜ*��T82QH��"O�� Μ�}E6��7����2"O|,2c!Z� yNy�'�L(G)���"O����Z�8���&�+DH�� "O�s��C�S��z���& SQ"O&Iv+�7K�У�jP�����"O�d�gn�+Y��A�e�_����$5D��ж���vE"'n e^���C3D�|r��ƃG�2 ��b�@*Z���H-D�0H�d�]�,<�E@Z�B� �j� 7D��qF�_�@}x6M�n���@�?D�x����*��2��U>��;6�)D�dsT�w0��X�` �*
V"C�ɫ<�И�-�*s[�2�`P6B�I�B7�!���H�5)(5ɀk� a@B��</���"���6^��DgӔ?�XB�	*��PQ&�.S<LU�C��wk�B�	,#֔�`
�8f� �B@f!�d�n|���J�z�LKq�V�g�!���|ܸҮ@�7g��9��W(�!��_�	\&Py��0Ud���R3l�!�dZ����ZC��76'�m���v�!���"	D�@�/X�Md�� �5!�d�%C�Z`�I- �\�:��E$  !�ԩ�����kY%:�誒�:{,!�D�9��f�g����&�I0i"!�V7Sv*Pv�J�	�H��AC!��	#��3��g̼��U"�j!�$�>�:,��kرw�X�W��r!��S!U��Љ�V���Qa�pd!�D���`��j�2��tI!�C�Gp!�d���y�����5~@+bFY�:�!�$��2j ���Xa�����B�t�!�d�u��d�G �H`5�V�6!��(�tm�rI���ᓤ�f�!��?_Xȹ��	f9�� ��~�!�,>(<�$��e0� �ω#!��^�ec�qشi�>u�e��L��!�!�J'�H�"@,�z�hl���7<!��J�z|$ �Q�x��ɗ>t-!�
M��#�$ܣg�&���Z�_}!򄚒g� �{A��<@��Т�`�}u!�䘦B�ڵ�V�&,���5mV�!c!���c�p�	|6b9iǣ�z$!�d�0q'B	��L�)@��1"Ȑ!�F=%B&�"g^�]۳�E�'!򄔚�z�����֩��"O�X���J�0C��;E�J�W"O�40�a^8?^8v�X'���"O���0ki#�l��j���"O���p�ԩc�p�����/�092#"O�#��U>
�~$��#Q���PQ�"OV��hD�gf��T,�g=vͣ5"O�#�L�%b��2A�樛�"O�1���7`|Z�����f;b���"OjE��aZ&(�p+˂��8��"O\���G�$3��и�*�9L���z%"O8 H��Z���ۄ�§}��:S"O"�@��	�����A����A"O� �Qq`���xO͖r���"O�́���8C��kB=V�٢"O�Eb���+H�R�Ht-��+�$9"OH����:W���ѥ�} $9�"Opx�u��V��hPC��$崜�@"O���,�H��8K�
��ksʉ�"O�q�ǃt �ZB���"x�r"Oz�r�'�sLfT;�jC51�*�P�"O��!J�B�n�j�(�.Ŵ���"O�LF�Gr�2��#�Щ{)�d�c"Op�!��3OA�%��8��ҧ"OD��'ɂ�npB�J�KO�{t���"O��˰�!T
L��'�(�["Oh�
��-*+���'�^��s�"OXɛrE�H���.�L��"Oʵ)�e�h3�	��e�+ߐ]�"O��A�6���SD�q�zA&"O��1��D!���x�F3<ȡ��"OF�c�g�<��`U=�=A�"O�Aa�
"%����͗-z00"OTd��=�($����)	����"O��S�JȾ@ݬ�9#g�l>��e"O-[v�*���t�^0]bݲ�"O^ӄ֭>��e���%#�"O<�"� ��8j��C$���P"O*)�ہ|�؄��&6�%�@"O�T�!. �Rf���d!X�U�0��"O����e$s��X���<ocΨ�5"O�L�NѨC�p���C]�XI�"O�]¢fD(k=|e`,��r��j"O(u�uH#U�P@��ôr(�a�Z'|��0S�T_�LJ#�:<O�ً5��+y4��S?Yx�e w"O(XҦ%W .�V SF�cƬ !"O��jTcK�5�"AA��B
'�t��"O��3oȡN"q���j��"Oz�"G�W��0�&�L>$<`�"O�!A� î�:��d R!Q�z31"O�pa$n�	L5�BN��]u���"O.Q�㤀�i��P0��>	��9HS"OD��Ɏ��V��ԪY4�Y�"O ixU�.r�&aQ�㼔8f"O�j�hI�4x��� B/*��!�"O6H�qhU�CQ"(k�-�4Pe����"OZ�q�BG���� :	��@a"Ory�lջG� �J��?~ ��"O^q�%D�?!�p���ߴ!��9�"O�p� � �>��`M+T�̨�p"O��Z��.$pW�R����M�j�<)���0u��n[*����WIg�<�sɃ6��1ȁ).�D�r��`�<����G�������=bG��Z�<	&+Lb>�4�Q�Oz�%�q)OV�<I�c�.߂����C84͚ɉrJ�N�<a��V,d���15|)��a�p�<�0'��E6k� �q�h�<Q�SAR��"�TS���8sb�g�<�+6$D(��&O�E��ɴ�Be�<y!]�<�<��Vˌ0JL�!�N_�<�C��b���J�f��A�k�^�<Ѵ�=�l-x5��7"�@���V�<�b�V�P�Z�9a�V�mt��oLO�<�) �'�������"�n`0s)Zb�<��A9D�P%�B�@�n�~�(��J�<�QBM&\� (�GI�25i�ˍn�<� ��y�$I�Kz2`"g���CQ&d �"O��7/D����`�,�#B~U��"O������<>ڮ���6F'|�*"O
��w�
�!Q�a�ak��x-|HQ�"OD`��%�l���ٷC�����"O�kV)W�zջ�%۱��ԩ"O��A�;�PQ!䈑 ��(Hd"O����S�!@���$z��]آ"O���BD�,<�D[�;x4x�"O�96�Τu�����R.+�d$Y�"OBxZ&�-.N�ADc�'\1�!򤒅W�:0�D��#|G�p��͇f!�dZ5=���DY ?a�pĈ� 
!�D��X�tqI�h$�a��!��܍)��� ��-a�|󄃚>3E!�$�c�f<:aɃ]��5S� (!��ǚC��c��y!���~q��""O|�Q�g�U�@Cm�lZ�Uc�"O֡�V'#U��x�͓2Y-���"O���G0�\`BG&��x��ag"O������.B���	�dR�z�45�A"Od��G�(*`)x���ʇ"On���_�2Bj�9 �J�.�Najv"O
���0D�$m9����_>jqz�"O0`�r��6_�x��Š5u�8��"Oḥ�C�~=���6@S�\�B�"O4��?V3^����g@�U"O�)I�J�6*p�c��W[�T�"O�M"�:*Wd�P� Dܠ@2�"O���'�q�Da�A��U��=h�"O�u8 `^�+�h���0Gl9�C"O��Ð`�yp�s�ϸ��"O5S��L7r2����M]#!bt�8�"O�A�]#\��5B���1CB��C'"Ob�3���=�v	 �f��g��t"O�t��M1i�9��%Ӧ=��l�"OVXIG��1@��Q��J-t4�*�"O���*I�(4Hy�p."W�H�"O���ڢ$ʤZ�gZ�E�p}
C"O~�!G��4E��%���ڎ�E"O�K���s��8OB�6�P=�`"O�����V=w&Ґ�d�Q�����"O4Tx4���O���Q��ç.�4��c"OJx����3^B���O�P��e�"O"0��/ɑ~*X�#�İ)C��1"Ol�9w剁2��Uj��E(���y�ꍪ�6-S#�G)"Z�����y�� ��aqB��;$Mi'G	��y���u��&�6�����G��yBn
�q�0��Ղ�:P�m2�f�8�y�T�w�(A'[6)eX�KC���y��i�L��s@D 2B�EbZ��䓜0>9��25!�������N�ƥ��
GS�<i$IY��	��J��%~��ReP�<��	�QV�CэJx�j��J�<Y1��5�����[pZP���H_�<�j�%fX��\��Y��Q�<a�+K
?�����G,�a�%YG�<�`�F�~�.��G�ߥg_-#��h�<Iq��Y��y�B>�Hي��L�<&G�z�AA�TY���aa�[G�<���M�j�������	I6�V�<�ƍ	hX�W��"*�8 a#�P�<Y���
8]25	���)B���gd�<� �����֍Ե�'NK �)"O���遇�l�!M�;*��Y"O�����o�T9�ЬǧnYt"O$R�
�QIzՁp��g��0y"O�1���Ģe� 8�E R�@��"O渑����6���Z�ǔ=Ti�P"O�3"�;d1��(�Л0pZ9*�"O\ա�Bƪ�rq`��A�a����"Ol{ҊͅqO�qa�E���С(w"O.$���]�<��D��Kk��١�"O�p���CIr��RşO3����"Ohб��^`� ���cO�� �"O�	�2���Es�R�k/�xs�"O�т�)M��nS��,]\9y�"O��!`d��S�$��s�^�O��� "O<�١�Q0{�@�Tl_�R�8"OL����#��$�&EX� �mѠ"O�415B�+��c�-=�l�K�"O~�Є'@�H����o�����"O.	1WGޔs��DЏ�Vx�"O:9�i$rƹ�c����`�g"Oڀ�S/�-wX(*��[� �Xt;'"O���
�A�ț�π*���b�"O��i�癁I���a��x�"O#��,��	���!�Y�5"Ö�e�կT�XXX��N(V�L c�"O�@��:!�h�G7����"Op���J�I6�A�g!T����"O6iS�h�e5�8� ��3�aH�"O$e���vD�\��%��:ܶp�f"O�u�ξye�EC��Q64-e+a"O�l��a�
��IAQ'�.mj��@"O��`L%�G2Y�\� �"O|E{���	ޤ��@Y
4ТI@v"O����"Z9�h$ۑ����Z�"O;���OkĬ���F<xfM�F"OP�PŎ[9!�i�#ͳV(`�"O�4sGbW>:8�уl�q��hs�"O���C̰|�B,��׽z�<q�"O���l���a���T�TzP"Ot������tq�c��@�"-�"O\�Pd@ݢ5+t �cc�(�V4A"O�<b2�F�V�rt4��*�PM� "O$X���i�Z�����~��)�&"O=:�f�t���QW�[B����"O�rF*�}��pX4��S�0�[�"O�X��EP29��hI�B=V��lcd"O�\���#F�`pf�٭%�Fȸ�"O� ��ʝ"����,ߛV�q�"O& s ��9O dBd�2w&���"O6	�G� gj�Q��ږČ�!�"O��̟$n$9±#�%��@3G"OV$Q�G�*�u���ȣ�"��s"O(q��k��9F��"��-��̛�"O���KS�\��u�bH k�Tb6"O�3�I�F�`�{��)�&t��"OƐc���;�����7Zu�r�"ON%����
!h���!�V��k�"Ox�x�C)Q�(� �>����"O��Z%#̔[�2��O��m�&0x�"O�l�C��pC�)X �ʒ*��+"OpX�q*O�6��1��wVp{s"O((0��D/�� `��n�S"O(���e�:.��m�$��@�9�"O� V�Peɛ�������R3�nX�"O^i	�#�i�� ��
e�PD�"O�ٲ�ͨY|�E���8"�|a�P"O���d�ˎ	O�� �EM�d�j5��"OBdz����R����t�0��5�V"O��֥R9HL�y  ӫQ�n�"Oй�mȥ s�ј4�ڏ�rظV"O�ѻ$mq� �3��&�&��"O���g�4t� � l�RUq�"O^���̤+��ٰ��H6'u�mɧ"O�LT���!�b���	;o��P�#"O�q�UMMQ���Bq��}��Yqd"O��C 	gwDe��:Qܤ�#*O,���O�-~F�9�In�L���'�$$CQ�7l��Q�W�+b�2��
�'U��c[8�q��"X���k	�'���C�M. m�L�FhߪWS�� �'Đ��&jѧg=��	���z�JA�
�'W�Bwa�r�R��W.uP&y��'c�0��UVN�35��j����'�<,�bH0r� �i-�Բ�'/u��)���`��B c
�0�
�'��0@�';�ڵ�F�T���':�D�T��#4*�AE�_�=�5K�'����[z}�e��y��k�'[~��S��}�>����U��5*�'9°b�2� ę����٠�I	�'�����D�aX��1vi�s.V��'�}���O�&��4+�"�Vq�b"O~��-0q�����V1l�{�"O��f��I�8'�+r���"OTp["A۝+u�1iW�t��A�"O��SvÜ*la����@�P"b"O�]�2k�Aq���ccX0'�0��"O��F��2Us4]kr 'q�9�d"O0I6j�
�� ;o_�D@˲"OС3$�4>Қ|����+�"� Q"O~T����v���+Չ �B1)�"O�|K���66{���A��`�h�ȴ"O�L���Y;�FY��I[z�JmS"OPc ү>B@�[�O�-OʸA"O
�V���PA���4��*"O,�3�RD,�t�ӡ�
Z@>��!"O��cR�#6�p��g��j8䰰�"O�y��/) k�ˇe�-?1q�*O0����K���k� ��e<$yP
�')bY17�A'��}a��� XK��)
�'?lQZ�&M�1Y��h#��I�h$�	�'ͰD򶥆~\M����j�9�'NHy�*]�O^v�c�̗�
\DT��'w�P��ITm��"��{k����'鹁%�7F�4�6��r6޴J�' P"�DI*Ȏlh�ĝ�6�L��'����/e<X0�T�{�Qj�'�� �2�dZ�r� �U��1�'Մ, qO(Y�r��r��*N��us
�'�T��φ�\��x��ĕ>p�	�'�y���x�@x���/<����'/�mef����DHԱ.Zl��'e�qrB"ɞ�<���XY8�'�x�ѓ�P>g6Ƞ� �(��(�'C`x�`F�Q��3�X@d;�'1Xp:TMъt���+#O
~�:�'�LA��ʖz/�Y2�D�+������� �|9`Nڲw9"D�c$�
TM �0"O�M��J��A!�u�!�6l��	v"O�\��O�;�˷���j�A"Op�en�9ki����LE�֔��"OU0� �		��p���8I�� ��"O"��G4Nt��q�F�I�v"O�%z5�I�7�����ޙкY��"O�T����T(��iA�R��z�
0"O�HȁN��B�"2�
�F�����"O�Y`���Wrl��1�
`U"O�M�q�	�t�Ȁ�䄙����"O��k���o�t}��*S1�h �"O6��f�� ���I�HȲ\>�PS�"Of��åE=dM�<����: �"O<�x���<� ��7C�;"��ԫa"O��Aa�Mwz:�Ɂ�D(�h�z�"O�[�"�5` 4�x ��":�"O�����?K����ʏ9�D9"O�� �(e���BCi��l��"O�Q2T�ѥL1�����܈&׆l�"O>y(eE��B�8a��/1$̄q&"OL:2$��k��A�oZ�x���J�"OjP�Ga�:���l¡\��02�"O�lQЁ��
�Ҁ�P)�,y.�"O2|Y僎^AJx���@h��"O�ma��Џi��P炻9`5Y�"OH��Bt>��r�^9ID�c"O
�B�I�9�ȆdT�O1�ؙ�"O����'Q�nu21�A�tO�<�"O�|����> 7�L*�K��(6�"O�!�*� Az���'VҀ"O|)��O�)��=�5JVX<{G"O��P��Ѷʀ���I�a�b)��"OґB�nޒ���1��q��9�"O6��r�Y8�h��J�,��}Z@"On��Y�8�R�0aJG�^[��1�"O�i�兔�`).�b�C��F�)�A"OV�䨃��23ڃi;Θ2�"O�E���f�t#v�!%�m��"Oxa+�#�(g���K��Ȁx$�$�f"O���A�P'{����P�f��4�0"O04ەk�+;
`A�C��iȲ��f"Onxj���7kz
@`� ��9M��j�"OV��A�@` � ��C��@�"O2����$ ڕ��n��qZ�I2�'ў1o�&���"%I�jfrk�!4D�"���f�)�Ѡ�8O��a�.D�Ĳ�%ٝUn�A� ��'�yi�/D�\�q��z��U���E�|{PL D���Sמo$"�˓��{��I��>D��HU��&���rхPD��@w�<D���F높p��a`�`�����'D�t�֨�=]��s ڰ*�lj�� D��h��6��P�,+�	z�i)D� 	���3 Q2Y�p�N�m��aX�,+D�H�����vv�(pG�̭ �ѵ(D�tH@���D���E̷r��@u�:D�������ڔ�#�U�s��]��A,D�hhP�C�^i��bT9��!j*D���d@��.�D�³H�;)�Ւ)$D�P����\����1wn���P"!D��x�.�}Ծ� b��5T��=�� D�\����e�X��Ï̖9�U�`d>D� a$!͔=}��� ؆!��0Ȃg!D��  �y��eӢ1!FD����{"O�X�M�42p�s�C;�x�{�"OB�X`f�*��/~|�I�2"O�=ؠ�I�{�V|�h݆W�� "Of�SE~BXm"@�I�U�r=#"O���T�	���5�Wd�)c� �A'"O�;rB�b\��׬��r��]��"O���&.�1zq@�Pk'l�"OJ���S�#3d�K�
)Nj���"O�$�0i	�}�@	3�N��fBr<��"O���։�2c~x([����$*p�"O"l�O�U�v�q�l��|)���"Ot��aF�Z�q���1]z`�p"O  x��;U2d�1n�\�D"O�<��I6	ؤ|`��[`��"OP�s4��k����2AD���"OJ1�b��]�p��b��a��"O^	��?�������<1�� "O��@��HuP�L)S �"`Ѽ�2�"O��[��!Kpp��{#�$��"O����H��=2 �:�np:2"O��)vhS	.P��P�l�S�؝�"O
�a��I�c� #���^��$�	G�OZA�E�'dPu��CM�OU~���'��=s1N�(lK�(AI�[��l��'��1Gy���F�:Ji:�@ ��ᅋ�a�!�^�q���ҁ��h�r�SA� q���'��|��9+�8��W�����/��0?!���xKP >�����L�b��<b�*O��*�m˄(���(r�D�H��u�V�I�����A�����w��)�Q:Ri"O6��Iѯ;���;�!�&/�B2�O�����S�Ph��"�02'"�:5�
�P�ZB�	�6�|�D����1Ӭ��*>V�'Wa}d��
�����Bj��kV���p?�O���E�n��[fI�s����"O��0����=O��PE��"O@QY�c���0�J�^��P"Oz�Z���Olw�N�jx&(��"OՁ�@� 5մl�#	[g0�c"O6=�Uj�4v 2�X��*`���R"OT��⦄�_@\��N�HxĐ�"O*`(2��z�ơ �G,=���K�"OB���.�z	�����F��@��"O\�A6���m��"̉o����"O*����G7eߌ �5L�.>��x��"OL�P���*n(��)4l['^�p�k7"O��$�O�?ݰ� �	a�Rh�"O 1S�%��)DБ)a$vI�Y��"O�Ÿ��*H�`t)`)�
H�!�"Oz�WE�^�E��j@;-j���!"O�	ӈ8_L��BD�ƭV����"O��"�"��-O��A�#\ ��Tё"OdY�3�P�~ ����,"S"O~��rIZ0B:9j��:H�R�P"O����gP�=ݖ�9����DJ�"O��hCG��V'� ��߾rZ|-c%"O慂��ߘp��˰��K��"O�D��ʏm9�m��;�Ή��"Ǫȳ�N�.8�Ԓd�H�3�@!��"O�)h A��
m"��/Vi"Od�����']�6���D��`�"O�h��CH	7&�ѡ1iG(<��H�e"O�L;AjL����aHI�_��@"O� ������W ��@g�:l�hZ "Ojĩ`(B<$&�jg&E�fjf���"O�d��T,� Q����'SBp"O�4�w�_=ED��ɐB��$�b"O�p�f�Y�%n��獃��4��"OЄ�mј@�$i1%-��+ .}H!"O�{c �0�X�N�1lT�@"O:�RoP��й���L+C��"OD��'�����pV�P�=XT��%"OȜJ�`̔|x��5J��l��"O�����K�uJj�/BAW�H�y����	�B-[7��	��q���
��y"D�7�&�q�É�t�4���Q�yb�_Ǹ�� 
�#)d$�&�M�y���8`>V\�@���au��pE$��yR�Tݶ}��'۝L�Ĝ`0C�y�&�'�|��`N�,3(8`�@�y�$N�J&����+�(���� �y�D_U�\(!CB�UX����y����g��ũ�	P�B�eҔ�y2�G:j$��ʯ�𔩄���y�� �L�2l�����c��0�y��{��A�IՋ�H���kJ��y�!F/���+�c�	N�h���yR���P9�(�;��br��=�yR�7hx�C&��Lq�χ2�y�Ϟ��n�c���M���w����y�a�2������Y?F�tҏ5�yRHH:�B���@�0U �I1��yRE^$x�4b��	RdJ�"�*#�yR��6:�R�25�[ 3_D<P��'�y�
�$!� ������<����yr�ԫ�X�#��P�-Ko�*�y�d̊'�ҁ�ք�$t��jwB���y�!p��i*�"P�g8��s��y���]Y|�X���g�viI&f_&�y�Lҩq��պ�FȖ[0�<J����y���X�a�O!VvF������yR���(�F5�`�E/I�]��
��"S�4f�nZa}��9OF��S�o�FQ�B�ĸ$�"�@n=��u��l� ��CA�2�qz�S[���'����=\�o�%a�� AC�K��6�ɶMi���7*�O�h8��>�\�]5NX�����#.�KH��갢5\< ��ia�����[C}�'����nT5,!�)H��ʴ�8�N��~2�'�'�"��OQ��§�țgP�����&L��X���ʦ%��4�?A1�i7��O��.�b[$<���1Mw\L4�@�-��}�'�X<�� q�:��$E"R� ��U���1��*
W��f��G�M�_	�j0x�&�?��kљ^,�O�aҌ_���p���e�^`��$\6�(�آL�1O� +$j��Yj��S�5x2#պ`F�	�M��U�!7���׃W���8�����M�6�Is}�Z
TsC�����.4|�HEy�Kn�(�D����m����S���Rm����HR�l�
\lZ��ڴ�?�'��)� ��fF�m ��BQ �hp�UI&f�Ab)<Oj�dȲ+�a@�F5"�~h��/ǣOXRL˶�
4!r�A�۴=� ]A��^�v��Ղ#�}_ʨ"�!����ñ@�ڄ1BW	V�^D�钁�&��ЃbKX�C�`��6a�zB�l����O��ؔA�� {u��b�m�$� ��ߟ��?�O(|��"j�ҵ{�Cε	�$+���(,O���gF�1�2�����N>x�w�O�o���M�*O��3�kZ�Y��DⓅ#�Q��2	k���7nl����I�y`ƬP���'Z�^IP�%B+��6��C�6L@��Y�s�.���C� b(�|ȴ�.�m�.�!��:E��,��9r\z��W����TU��R!֬S��5Q �i�Y��㞘�4,�OrmZ���OnX@��:m3d=�`!'fX�K�'U�On�=��4,�p� �[��'jz�q���*�McP�i|��ЕBA��@��^��p��Q>`�m���0m�ܴ�?�,O�ʧ�ēo���ׁ� �����P�g]2���oV+Jz�J�HQ�:��51%�ߍU��җ�Ů����W��9`���*O���^(�M�u%ΕGqؐ�v���uM�`*�!�DP>LQ�aL�b����5� 8pyP�]���p�(�1�̂Ѱi
,�+��k͛v"�<%?y��M�`Mļ9�$t�d��6𜰃�bU~?����S�U&���+�r����8��<Iv�i{~6�7���S`��=�.�{���.�Pha��1��I�68���4߰<Ij�Y��E�*�6�,�Z��Pθ�0��ؕ���dן�M�#�?]J�#��zB�O:$��ɂt*�� `�����sjO�����%�V\���ă�eA��t-�%�6_'°�-O<P�G��<��� ��2 i*P\���1L�O�l�*���?�����Ȟn�D�U�LGp�]>(����	b����O� g��#��QBp�6qf���h^��M�R�i���b�d�$�4�i5��fӬ}��  �      Ĵ���	��Z��wiD�:\���C���NNT�D��e�2Tx��ƕ	#��4"�V��񄛎z�m" ���T$�3F~,Q$��2~J�@�M\h@� s���Mψ��n̴'c���;p80��'gF]� ���}�V��ʴ����ś
?�]�/BNy���8��"Bm?}���w�t�q�ھ\`6�QQ)����;'�B" "U�'��1!w�6��|h-O҉@fC�?\�p��R��e��t�.�+�%�L�LRZS`d��6@�l��'�V����CbډOٺ�#�B�(q���f �-&.�(�j�>�Kf�@�O6�ēU�xҤ��:��T�ڬ2��P��G��l��$��~��G-�,�7�x����<�HX�����1�Ɍ]b����H��Fq�`�A:��/|���k�?U�?�:�U��DЩE,��& B�ڳ�.��@
L��U�4�|i/���*f��<�Ro�7DU���W/�'E���b�dCܟ0(Ǡ�0t�"}J�O�.rZ�D��,K�Od��'o%�1����W��Q�$Ô-v�<=Y� [����B�'�y³�m}��hô'\a2� �W�r�K�^�@�P�1O	:�M�2.�Oa�$l*��Č��?i"͆��b��{���!$���rVA� C 6E� �S�Y	��z��A�g�牡�y�*�
Eo��l:�I�&��QW��1�z�3�8'1��b�Ɠ��O��x����[��	����T�s�X�Ӎ�5j;i`�a+�D�<w�ۼ5j�<�4A9�ď[�d0�gܚ<Z8Uɐβ9��$�)�O���J<!�Oh��V�$$��k�'@:u�H�U�ֿx#pqC�"��Ap��eΔ�XeX��gR>�1�	T�.|n�����r��w�͈M��h"`ѻF�u�'6�dY�f����{�jE�Ɗ@�Iih�Bю؏#2�|��\�}Θ`��1�OL�ږ���1O��1ԧ�;3�u�� 8Ŧ|@�� ^��B��l & �  �R��D��lC
��!��yBO�'Nl�
�B�9o���*2�۸'��CS���KϠA82Ɔ�N����G劍Z�F}r�#����	�]�H$rcF��6w�\�с�; � ��=��1,OX�c�`�H-
uP!(O3P��J��Sܓ��π �����}FE��b��R"O��8v��E��[T�l�˷Q���ŀب�y��Ć��g}ʟ�Ű�.�� ��x�udI)'$   
    P  �  �%   ,  �2  7   Ĵ���	����Zv)���P���L_zX�R��4�M�����+F�'��L>�V �?�敊����qRj�H�<)R�
��ܩ¡�/CH4(��K&o��a)�(�M��Łt�����G	��9 �C�;W`d��6I:W��1�ǤyR��7,���,�)��"φ�;T��N��[�.�Q�����ʲUI��A�)�kҚ�q�+ǒ>��|���FB`Uh�L�pN�� 	������Qh��d�F#S(#@�d�OV�D�OJ����?�'8i�^��GEۓ�!xc�x��ɄZ#���\�]��]A2*�4t���P&E|��	9k������'MNM�e��vi�Т� 1m�I;����l��ȣ!�
�:�j � F��$ːY�3'8D����Ys�p�4�\#f���vӾ�Dz�O��'H$���Y%e��Ajd��	�Je0��Ʉn/%;��'���'�2�i�I�I쟸Χ|b���4|M�a�޼uЄrT��4�R��	���$�,T^s�D�	O( LQ��*�Z���ɽ(�V��T�$*z%������8��6y�f!�ȓm{�R���Y[�-k��O6[Kdt�ȓ->,P*�*Q�f�9(�E\�"M��'v|7�9�ċI���n��l�	oZ�I�*v5��V>v����Eצ6����,nb�'����xz��ԟ�����R���4��2e|)ۣ�I�U�΢~�`�G B*��/��J�*��p��[�'i:����ts>!a������0Ŋ
c��p�+D�
��X4EL��K���-@�8`J(�O�}�'�24z�@=<�$l���K  ��O�=Ԥ�Ц���՟,�O�i��'e��ɸtڢ�RT�W�-6�])�.��K.�6M��n�B��&�|�>��ǎZ^��@ N0>7|���K����1bc)�S�O;,�b#�3e�ы�
�o�K��?)�؟��M>E�$jN6C�l��Ti@��ْ���	 !�d�9H����Y�s�L��&�?!����*��i[�|��"������$�<g�*�o�����,H�<i�!����IƟ����?}�i�i����d��b2��1H���Ʃ�<I4�u8��{  �:%�B�ҥ�S����:�¤<1̚c8�fBV����$m��%��,p���<�S����@
ӓtR$�u�
"GX(�EŋS�tl��x���s`���R�jiա�(�d�o��HO�9�$��f�����ܸf4t K`ޕn9��P��S����O��$�O�m�;�?i����GO��?y7��@S��Q� 9�XQ�C��m��}2!��~�	�6Q[�
3H��Wj��>)jBğHi0e�%�R�C��0B/6PB�/� �yB�݅��!�g럀.%�S�dH4�yN[�$�hL�� 'ĭCu,[����UߦE%�hAQ��l������'5B��K�>I���� "���oڲ^�z��	�8�ɝ[\��	~�S��M�&X~Y0Wn�:$:4�{��A�'Ap�2��Ɇ2c��%[�NV�KѪ	ʣM_�|bў����O��G�T$��t�u`�L�T��Ŭ���y⩋�v:�L9���D�Lq�������>��qbI��?�p) aD#2(�!�>a��"�F�'�R]>�0-M�����=yh,�!D�Y����P͒�ܴm�����J� nNd�O�Z̧I� \����$�y)��ڳA���9��������x�27��w���D��e�
)0��	sO�z..��T�%�r��?�ӓ|��	F;9��s���x�N�2���4�\B�O�6��4��	h�nݢ��Ӏ�&"=���Ӧ2t���%Y�5����fA�ː7�M����?鲉��vA�-����?����?�F������;&c G%�pr3K��0��)��cU"&<�d�q�f�8��3ʓGK�Mp��-����e��d��L�7�-Y� ߦN)t(����4o�+F�1O­lS1g'юS*!Ѐ^�Pqp�O^��IR��Lk@�;&$��;#)ׯF�C�I�|��ڒ`\l��@P�I�b�6��b�����|��'�율��v��Re��<�<��$�U2�'r�'V��'�?���Q��+�I��MgT�A�Jaë�Gv*��ӼC�Ԋ-��#?�q�,#�>��a4Kp��0EE@�A����e�+�Ҝt���at�w&2Y(QA%��3���x;����S1-�|�vț� d9�cۓ�M�����˺3+O�˓�?�R�+j�ŏ�"]§%����'Ƭ�=�S�?���|���-e�4�y���D�3op���'V�7M�O�u6��bߴ�?y���?�16D �'��%iU4A*��%5�8�m�1�������B4��əy��H�' ñy>����O�xS���*2ޖ�����1:8x9Z���D�g�)p���,� )t�D�n�خ;π ��s砃Sr((��چ]n����� g}�@�|����?a��iut6��O��.`F��̆�Oyh<z2L��w$�7m�O �$6���O����O��8���S�G9e_�9�lרg������x2o.��|��'?��'?��]i�P�l��u�5����9�Z���e���M���?)���U#Ô�?���jx�����p�^��7j��1���2��i.`�QBH?l����'��R>������@HȲWL»B����B�}���H�O��8Zw�?���O�����xA7@F�e&�-)�L� 9 ,d���OflYv�'[V6�fy����dT���F�t�h�Z����|9��c5"�>Q��䓧?y����O�M�h�#L�;�ڔv�`����$�ll�^�i�M��	�;{K�=�6�D�  ��R�ߋ1k�F�'�r�'�@��'���'Wr�`ݕ�	�%�,3���7uF6=١�^�֠�ٴ�?��k��*8��fWax� *)��	Q�^3�F0[T�����O��+�[ 9�����I�}�ѯTeĭ	p�t��I�SE˓eq�'���'��$ k�R��c��w�5%�݃G����'�"�'�򀁿��T�'�ҥ����_.ȵkt�$�D��Y�`�7-�F}�^��q�����<��LM/V�ܼ��J۰������.#�t�BUM���?i��?��V5��O ��w>�mX��$�%K�1z5�Pn�!�1{�Y�I抄a���83����S)P�Q���T��T�Q�R� �3�	݊&߬x#���	��+#�%j�i�K� Q�����Ob��i͏)����ejZ�3�T\ytOLܦ���S���h����F |� ��%Fܶ *ĠrGJ��yB��2��9�&H�y���pa#ͭ��$˦���JyN�P0Z6�O���?�s"* ��~)zt�E'(��B�j�<��O����OhH�$B1v `eSuE'�Ȓ󢋎�����w,���
�>}Ԅ,�7C�y�'��EZ��Ε<A(�+��R/l�Y��[?&�RЪ�<{ԦA#��(�*-E7�O����'~�#|2�,�+����A$\�=�xJ!(I�<�S��'= �A�GK�Q��q�#HX�0�O��x�K�r��zbK1#.�h0P���'�Ғ�Mc���?a(���1���O���.������)�:�Vl���Rn�:V����!GS�{��A(O�Ģu�$͋�S-1��p�I�7�<��+�E�qe�S��l1�.����Y#�޶��O~y ��2�^(yCP�c��]bb�'��)��s�ɧ���i�&��,K�XYo�F�8����4D�0��Ѽ2E�X��EϏ��i)�!1ғrv�?9At�@� v��1�dK e\،�k��M���?�F�D�.�̙���?a��?	3��P��ƌ��7JP�������;$H��V��@ ?�OԍpY�(f���P�T7e��i�V�����/�O��Kg��%��|#��R�r�d�b�T� ��M�Oڄ��ɭo��)`M�2���4�&�dB�ɓ ���0!��"VFj�'��8o�r6� `���4�|�)σ �~��s��+���*�O�*�%ɂ�)D�z��i������;g�|�Ibl"D��
�"�>��$cQ�F>a���$D���u`�N�:��#Y���!э4D�|'"Z��@$yV�_7:BD�cQC.D��+c�̛KZyE�Y�m0x�Q:D�L�s&tD����F.Y��BE%D�$*�'d4�$��*����@&D���孂'0���O-��%�r�/D��9���PT�8B�I��n���0�'D����'ǿ-�J�B�D�=0��i�'D�0h���y(��TC	c����0	1D���'�
~��1��&�N4���:D� "���s*y��m�6��)P�o'D��┢ښ9xhU�ǭK�)$ȵ2g�%D�8p#l�0n�
Ș���2WGv�Hu%"D���%�����	%oAC2 ��6D�ġ[�I����d�N"_H	b�3D�@v��a���1�$�l�Ҩ��G%D��`��M��I�/�.������$D���g@�
sn��Sv�چn��za!D�4���;���k�Ҷ!�v�.D��(D�5Eu$�#lж#��р�o&D�|@"ˢwA�@�`�1����q#!D��jW���}�0���A��'d,D�hKU�Ľ���&�yD��E�/D�� ���iO�ɐ`$�N�cX42�"O� HE�	]�u�t[����"O�=sj�/&^PQXV�A�̮I��"O��)�U=�l�Y�햗C���I#"O�<# ���%g*�����;Q�qb�"O|�u�è�:��u(Qټ�H�"O0�B�o�4*�$��O�nk$I�"O�4hm�`ؑ�G���0��ԓ�"O<j��6`�`)�N&(ƆPZ�"O,M)UA\>|����1��0h�
�"O�����?f�F�Yvɑ�l��A�P"O�m�F)J��ت���5H�ꔱ�"OZ��a��P~ �� 4�l���"OF-%�� �3�N�4�:�q`���yR	��V���䜻:��zc��y�%�|ʾ�0bD0._Jd6��;�y�*B		���*M�,X���bg�0�y�%�6�yC !M|Рa�=�y���z�d�f��F�s*���y���nŎ���*�\��!��y�ߐQM%��J�j*L���N�y�f��>v����K�e����B�4�y"�Y +y�E
���+P�1EG�"�y!��=� ���B�W@�����
�y��](�>D� ��8 .J��$As�<)��>���I�L�=�@Ԣ�H�S�<����RFl��'(�f<��{�<)�ƈ�l�!��WY�~��Sʟy�<�VJ�.���/SQ�����I�<yC�F�E'.�Ab�%0�Hf(N�<Iub�5x;�q��Z#h9�Hxu��J�<�ւ��� 4�4��c�$G�<QQHK�\REkZ�w	ON�<q�-Y�Q��|B�Xb%cSTA�<��f���f��#� 0���Z�<)���c].x#G쌀93(�5CR�<��%ρf�t��&�>d���s�k�<����2��!ʝz$c��p�<1���(��RFA!��mQ��p�<���Քj�^���a�<��V�LJ�<q��p(�W[�N���q�N]�<ӥ�lf 8@�XI��1�B�-D�\P���L����Ï���1D�$�E
:H�cDU�Ģ�$D��Xb��m��DA�*%��d-D��h���a����.�h��@��+D��x����
� �ѵ2�V]�7�4D���.�)��y�J�$h�<ŀa�?D�p(@Ά�JbTp��<�@9��&>D�����!R���H�'<���7D� "�B |-�(���-#�6�H�0D�@��c�jH"�IV�B�q��+D���&\\R��F��9 F�q��k&D��S6�X&r(9M		μ�ʓ�(D�|SebҊ`�����H�-�B��e�4D��R6L
k��H��C8$|ਢ�8D����U	k�|9���O+_�]�W8D�Dk��+;>�1҅L̑rNt0IQM'D�@Q�� �e��B=� 0%D�9�c��2)z���7�;` #D�d�Q P�T:ش�&T(xg,T�U�/D�`S�%���0��L"�<*��+D�<�C�
pi���!^J9���F�)D��S��}�]flɻ�R=�$�"D�� ڥ��N�S��=��j�V���[Q"O�iP͟12S��	�X� l$"O�y(��*���`���4*�"O�-�%ȡMM���eȆ c����"O` �!.�,U�D4�#�� a���9$"O�@#3"�S��(�e-˟.�.�"O$把�ܶ}�l��s>�I�"O��0�/�@�0&���Ic�"O�)[Vk���H�C�� �uX%"OR,���b���+���|���8�"O�ѱ 4Z.�2�	�M�Du�"O��#��!/�R��� 	��u�u"O��s$Ǯ!�h��MM�bM�G"O5P�����P5O�w��֍X�<I2e])i�4����;<��܈��R�<��ڂfyt4k )�>�.��B�	2fD��&�o��I��H��B��3�8��dL$$�]��!K�]dB�	0�&ؘe�;��Q3��E�PB�ɠ?�X@n�e�4b�B�
�FB�I���H�Ď�:�"��b+N;�(B�ɮ~�h}(�(�����X��߽	i�B䉶q�v���l���X:��\�Q/^B�M�j�(��XV�Dzg�"RVB�Co2�9�#�8t�X�D
�v 6B䉴3�d9hg*�{YH�9ġ�_PB�zb*�+�E�6�Ve��/ڶ.�C�	'E�J�#�Y R�������G�.B�I?	�ld�BA3]M �B�sY4C��}��ݱ�Ё0�Y d�_�C䉴E�r��F�K?�i	U�)��C䉸���ƁS�C_�))5#;�C䉣�:����:�J� 0 І ��B�I \q�X��S%[v�+$�d��B��O��h�ġ7

���Y!xC䉹G��H�r ��젃��ԪB��6�tZ@�0!֤�P��-_�BB䉋X�F��NI�[�r�� I&S��B䉶~)�<`�g_�\�n$lLg���7?>%ZA)"�YсM�F��K��Z*���v �9'x��A<D����Ƀg�$�3��I�N�2�J0'D��YE��<EN2�CևݭI�xk�A$D�4h ���3%e"w-Q^�<���%D������l(f��p|�襤'D��9���G�$;�(%c��I��#D����C׹A�H�B� �wnxj`!?D�H���Ղz���a�lX @s�1D��0��tZ��C�&=ߖ�ré:D�h��ש=�X�@��2�H)H$F%D� �*G�T�E	�E_vV�JB&B�I�tH@��jRT�!'R B�	�w�8ʦ
����jH��B䉖C��@Orz���E��DA�B�	�G�@���7�Q TΌ'�C�	�m������0k㬉��BW�M�C��!r{n��6p_�%��9D�B䉀t"T�w�Q�j��F��@�B�I#^}�=8"͇�V�|�0&�ilC�	;B�l��w�X��=ɕ�J*C�I�Q;cï��`��'�آe��B�I5st��H� ��c�&�0��A�B�	�g�2�3�O��w��C�D̡!�B�I�o�qقƃ�Pz����>e��C�)� 8S�P�o(j`�͌
N���""O�m��-دB#8�P锰J2���"O�e��Kz"�����/�̹�"O ��Í%G��Rr�w�`��B"O&�uQ=۠�A�C�J�:�"O���dNI#s��Ѫb����<8�"O�@RB�^	/�U��A9'��Ԉ�"O��@#�Y�\۪�HC�P2t��%�'"O�9cR�8[:}e,��© "OB�9TR�-���`c�D .�5;2"O�����j��@we�#z�t��"O`,)c��  候2�K�W_>�"O����F�R�跀 [q���V"OX�2 �9g�^�1�Kgb��"O���@�:l������5\���G"Op�*���v�jA!
!3C��I�"O���k�yb�ty@�h����%"O^-R��[�{r��fG��䌐�"O�e��W�ұ���� ̜���"O�90	�!R��9���:f��	0""O�2��
R!�w�C8��8+D"O�	r�%�7|:�勂���\��IÅ"O�<Ct��50�� �K�'���z"O4 )c��vl��@��
u��"Oe�m q�4��5b�14�l�)�"O����D�54�W*
U�Ե�e"O<�B(۝b����<m3�2W"O"��CׯE������	4�2"OJ�X��9�ĸ�� ��jBBai�"O>�3$\7����"�\�j۱"O�X�ua ?9��e#���"O\=x'hK�,x6t���Dgi�L "O�EX�N�t��(P���]�b�yS"O�����L����cٖD����&"O�4�6�Q���Q���>!_����"O�
G ��_�Ja� ,Qx�{s"O(����$Q��P�J�E���$"O�|{�`%C� 8�����H"O�l�B�´jV�2��,/3FHJ�"O�ps��P]���b�H;E"OVar$ƟF�&(sT�Y�6�y
�"OB���"�-|��B¼L��*p�'En���iM� �&@Rǐ<PְZ"�G(T�C�ɞ���p�GѤ;Q�A�d�P�$C�	>Au¨�0��>9�X�㓍�_�C�ɼ��9��o�x	=R�i (��C�I�6���ABO��!���Su�0C�� �����l�,B& �+���ex
C�Ɂ��xq�PU�:�0���@C�ɾ��%���͜B
�"�*бx��B��6,�g��>�8�'�O1.�C�	�Ú�q��7M:��J��E��B�ɔ�b�IP���a�0�2���/=�C��S���Y���ਓUFT�~z�B�	�|�ҽ�$�.e��Xa�&v#�B��$��D(a[Z��͸���40C��8h�輓��_;e���j1��#"B�I�lK.�P�"��S���c��W�s��C�ɮk'|(�`�6J�tyF�Ȅ'&�C�	�N�H!ŉ���(-]t�C�;��a
aу-,����#h:C��`�p$r�@0&��dk"��/H[C��

��-�(L�ȴ	ub@=2�B�	��HE�g�품�Q�5L�B�)� F�Q�*Z�+H����8$h�"O�����S�o�ZP�$dIS2��%"Od�+�K��P3�H�"���8$��"O�p�Wk���̅���7t�FP"Ov�A�ᇷ"�������={��)	�'H�p"cҤ�&(���ș+���'��X��,��R	\14⍣xj}1�'�Q��NE�2[B��@�t�h�*D�$��T�&;��jtn�S�~d:Pi-D�ܪ����\!�!��B�O.|�!�$�9sJd����k�8%��"тL�!�g�4�{�HG�C�Nl�T!ډzt!��
1 [��P�f�^���p�%C8q!�D�QO�@H��=���zA��!�$Ex�"q*��ޚJ�(��='�!�D
�IR�]��Dͣ�:X�w	צ|!�䌛Y�z��^ 4�zpqSKԥ	H!��0lR2hҖH/c���I�&,!�Ǥ"���W�2
wH�����J�!��M�T�1��(&�a8g�E�-�!�d��C"|����5\m�gˌ1�!�d]cDT� ��"�4`�o��v�!򤜧��u���`wJ ��/�!��\;�*�`BF�gnش�
�1L�!���K��0����eXxx��FA0v�!�$��\�2!���;;ڀ�'��0k�!��+)ж�$���>1Y�e��6�!�D��(?���)�8��,ʷ�K3�!�D��h�J��ea77� ��#F�h%!�Ċ!��8!�˄��0�"֜p0!�D��[�#�|0tP�D�Y�>�!��پ�t�;T�X)@�����a�!��v@�J��ʷR�<� &И\�!�d�(l�,�*�K�`�L��5C���!�D��5u��� G� Ԡ��S�%!���F5l CqA�/P朑�e8Q!�$��W�5�dA@�H���%��\>!�0hQk:q6)ajʁnt�"O�%!�́;*n�!	-{{����"O�4�lZ�H)�x�TB�
���t"O��q]	J��F�����"OD�3���j�
E�?MP�B"O" ��;���W.P��f��"O�X�gJ'>�8M��)����"O���P�ʳ@��A�ӌ�����`w"O�����VM�hY"���D�:p"O��K��Y+X޲(�v���l�8�yb"�:w��J'�J<T|BH�ᣎ��y"��x����hT#|9�n�/�y�F�	Z�9��K�0�X�� ��yr��@c�����+kP���Z8�yF�5=���&�#z�VJ46
B�I#SPzd��֮X�)�%�4,q�5�����O���W�� �(��Η#�"���"O���,
�!v`A��T� �T1r�"O>�9�i�^�� %ĠZ����'��I�톧5�`�.!�9Z
�'�	+�@
F ���̞��'{��ȣ��B��#�	�Y��Y��'�� Ꮒ ui�1/ʥ?�0,A	�'%݋�k�_�Tı�!��@m��	�'^�� 䠝�W�@Bj� ����'�Y�գZ
�\=���"|-�X��'�0E`�Ώ�)]�}y����҅�
��� ���]$5Y4�s����Nu�"O��΅�D�~h�N݊ڬ�2�"O]㵏��Q���-9/|r�"Of�!R�J�'C$9�J�+��a�"O��ҡ�0:on|� �=o�QaU"O^I`*�8νh�/^�|�.Q+�"Ohd�%�\�RjF���ό�XS"O�]0��V�d*$��d�,��D�"O\�&��
㞕� hX�Y�Jd��"O�x�0�K�X}h1��<(}�P�"Oܹ�&lO�j`�����XD(�"O>�hf��(}3�"��T�z(`"O�}�Ư,!lJ�rC�F%
����e"O�E�f��5m��y#T"���3"O`��K��\�v@�'$�j��Q"O�����L:d���64�>��#"O��N؇FRh����f�i�"O����X�f>4�J�͉�[�qk�"OD�ɨB�Q&)�>10�;n!��(̬cp��fx�#�,no!�_�$��N̥=� �����"	!�'K�m�'O�
�`�B�'�y!�;d�A,�9EJ\t��$l�!�Ž��P�b;4D޴ۢE�;�!�@�N-�PP��ɟ�}
��H�!�@�Q��+�#�$p�=���!��ͮ&R&����Q> ��xi�HA
!���0�j$C�1q�E �GU!�Ē�l���k��8B�e!��-�!�d�j$`�퉙vx,�ADOT>J�!�B	���z�=N����ΟHё����	�>�V)k_2�\��m��C䉔+ꔋ�Ǎ	W>��7�ӜB=�Ia�E#���� �t?��RS-\�n��+ю7\O"���y�b��\��q+�öl��U�3���yb��jS�d3���6fH� �����'�yDyJ~��h_�WR�P��ɫevХ3s^z�<���^��a� 'k�(����l�'z����ҽ:4����.,�@D3Da��$�!�[&XF��WH9U�T!:��C�jٛu���Rg�	�A��Je���&��r7�4lO��l�G��<��t��g.|.�
�3D�\�B-�~l*@ �,T�bF��gj.��L���'o?d$ۇAW8w˾(bPc��^"���r�� PLˋ��%ji�E��}�ȓ9Z�y$C�wR��	�
ъiW����&Đm#cb��v���1@H��H��Bf ���M2j���QR�ۼU�؇ȓ/�-��W�Xj��j:`�hć�i�b���� ʄ(qBʠ�XЄ�9����
��uPǀ��t��ȓR�.�����9��@��)}���ȓn)9K�*�'�����s�l�ȓ:Z���r�W�j2p���K%~T��ȓ!����gIV�e&�)z`؅ȓX�5K]�s��1)%�ߤ4�K,D��I�C^78�f�B��;? 驑�!D��I�|̊A��F�uߘX�2D�0Q,��P,,��mO�_ bhXr�1D�0XLD��!ЬO؈Q��)D�SIݽ�H�2�f�q�P���L#D�;h�B%@�^28`:Щ��?D����
K�ԲŮ7;��[��+D����K	04�@����s�%D�� I��M�"�r!Q��4r�n��"ObdaE#0�2dzF�E�I�L3 "Oh%���&^a�0aD6Z7  5"O��:q+W9W&Zy�B/N�j:�ђ�"O|mp�%�fy0�`t--=N�-�"O�Y1�ֶG�H����
G
��"OP�h�0o��!�)Sc��Q��"O$�Pd�Q��#6��XހHz�"O�Lba�S�I���Ye��+	��UPv"O��1���Uy��HѦ�;VL�"O*��#�7@��y���RN�)��"O�J����^�J@�B�OlAZ�"Ob�zf K$f�>0���	���"O^!hè�\��Rd�J(%Ӧ�{"Oୋ��C�CҖ3�CI?=��͒�"O�,�%�`�.�Ʃ�^�|���"O-���܊�$2��^X@,��T"O�У��4�p��i6S�!&"O�iU��V۰��2�X�Uئ}q�"O��js�1����fP57�$S�"OA��' �mF�0���U6x�:�"Oȸ�TJ� p����p�R;0QR�"OF1`�hB�Gt��)ś:�1$"O骵�2�N��#��lؒĻ�"O2Y�.�a�Y)D#�#MȔ��"OdA2BO�	4^��䂕^����T"O�8{���,k~,2�A�e��X�"O��Je�f�l<�5�� y:x�E"O*��2�G�T�bPxR!��G	La�"OR���Ԗ)3.,�g"	9���V"O*�*��Q����KE�,�"O�`�V�~�V|{�o��w�"dIe"O���Pe!�9� !�06�T��"O�٢M_�	2t�"�����p��"O.��@�ű3F&����*1A�"O�u)4��+��ٰ���_t�h��"O�h��X4�P���H]��xA"O�<#��N�]'�DZ3�
��`��"O�y�GM»p-PSw��&A�a"O��d¾��D
u��5�"O��;r�����[��Y���F�<�8B䉿0�"�W�lN:!Cu/�!w.(B�I:<��}Ez���wcB�	"Th���;
�JUcE�mg�C�	�EO|h`�P$lV��>j�VC�2u�`��r���7h4@K&�D�_b�C�i\� �  �      Ĵ���	��Z��w	�;F���C���NNT�D��e�2Tx��ƕ	#��4"�V���#o�m"� ��3��D,��j��Ljc��Pr�²V�9��b6�MK�͍�J�.�,ÚA�;lw�����'%4��ŧb���9�(�=.�I1b���a86�Qy�M��\�X��`�8}�oנ}�x�� 1�$�q�n��2v!)0���I���'A�A↤C:SD��)Ov���N-�J!QY�D��-#^\F�0� L� |J��!��y�E�i�I2 �@Sd��{��H9��{6 	���Պ���&H3�E��V�' (<��fR��'�$H�/���i�$��Ǣ� `tM��N[����X3� M��"� '_�e:BC:�)��_2��Q
S�u�8�d�*�Ma�$�=R�6�'�c4����#��h�2�J
{^�@ȒQ5Ȅ�"�,D��&�D{NK�U�V0�M���nCq�� �9Om���.W���b�L�&T]���'(��uN�>��3��c$f�j?Y�:O��'�bz���	M62�h��ɒ<���@%�'}".[�p1=�I>�A�%6"oZdu��Pc	��n �"���x�f6�_�<Y5/A9{��S�� ��4�OR����Ǔh�l`��CG�E1v�y�#	Z�"%�6���܃�'�����	Ay�Okxh�g@���Q:.�R�̠ bXxZgbh�ɔN}(�I�C ���7[e`��s2O@�r-� lxq!@F	�ءbQ���f�Q��k��x��g��uz��U�JJ� ��7�~r�d�'\N�%�$�'!���#�(r�� X�hW.
 plpB>-X�B'H��P�|	ǄƄ'v���SR?�z�,\�<>6X	��2�\�BE�4�V�*�<&���'�J���~C�'��Y�,ߺ��jS����
(r0��Gٍ �j�5��``��$�DҠ� h}�b��v  �am�(ԯX�G�ق�z]j��ȓ�J�  @�?�Q��r�ȓw�@e  @�?  �NM⟼;���X�t ���>S�b�S@�?K!�d�+��(B�[\�zt;�.�}�a|"L$��%S��ID1`�B0q�	*p����Lo�ʟ��	Y���*G*R�''R�� �8��AS8.�J8v&O%��cB�'1O�3�>��(!��=SV��ʏ����㍄	�O?�� ��JQN�>%
а@��7c ݉%	
��\�$6�)��|�q	V��(   !
  t  �  �   @'  �-  �3  >:  �:   Ĵ���	����Zv)���P���L_zD�R���\��Tx��ƕ	#�e&�T���Y�k��(kw�,{�bHA��$D�<RG�]�QYh�@�3���*�K�!pO�!he�Tm��a�1ɨ��I����@z pg�9��\jI�/lw�� !�^	!�BY���Ǭ[�<14�,> E�!��>MSV�uN�O8	a��U��9su�¦O�Z�X�#�0p��`�+4��JH-4�t��SI�!5��� RA�v����>���'0��'�v���wA�3<BI����j�vp��cM=��D�3 ��|B@�)<�
��!jG9a�bH�%����N�+��|r��y���3���=a`�%eΓ��$�'��H4LO��qA�!�޴`��W��@b�"O ��O�rG� ��	���׿i�
"=ͧ��"l��˱�ůxH���②yc0�CC�M�O0�Ȃ��?���?U������Ol��0U��D߁<�X�G&ͩU�zݰ�	�?��q���"�J��&|��t�VBޒeY�	[�ra����[�rg2�Ϳ�2!�$��',� 1�Ŷ7NtC�I�@(j"��<�&d)҆�E��B�	;����c��!j��C Ðk���ʛ��|bL��7M�O��?���
�-	�(�,I���D�tӺE ��O��OH�+�'�Oc���HC̲��߽a���`D/�Q8�=�v��I�O��)���o�rX'ǋ�6X�0���d��n��9�'A��K��Bր@��B�s�u��u����E#6�����K��6r<��I�����9�6�A �>Ow,@��{��I0;�J�۴�?q���I�,%�`���O$�d�00�Y�7�ϙQ�̄21D��-������<���'j�y�AK����[�Q�I�zeZ��iltGx���h�%h`V�Fm�E�u���"��[�`Rn9���6
�����̉E�@Mk`AKAD.��9>��DiΨg���K�	�<Q�v�EzB�1�'O���0�bA%��٢d��'D�=y��i��'nx���5!���'J��'��T��5���8�(]�N�k6@I0����V�|2⎺_��m��
JB��UeФ��d�0	�|��
�W��x��C�w���(�
�;���3_��2LO�LЂF2P`lX�m�&M4��"O؈���T`��8d�$A�(�6�i�"=�'��Eע���O�&=;���#�A�E��i0ӡC3��X����?y��?�"����$�O��95|�$Ύl{����F�$�	�`@[������l���	'[�AK1I��;�z����.04���.62��r#<�iT�R=.���a��_-eA�B�ɴU=�E����%y_"yP'�C�	p���q,L�M����rkC�����'�ܹt��͟0��矤����ԩ�e��A"��׹��Al�Xi�`���|�I�+^*�IV�S�O��$�+��J�eW*P� �Lj�'��]����#<��L��P�p�]Y��Ŗ'Iў8A���OrG�toZ:G<����{d: ����yč9/� ʒ�t����˓��>�$���2�I�lR��E��4��U�E��>����6����'��]>!�c�L����?55N����_�M6�ULH�u�t%��48�MJ��Ü�R��O�\�')�V�s��VE���:�E�!3Q���T���P���S݈P2�e]��F��nѺ:���A+͠]wz��%$��K��?�A�|����Dߪ0h��	�
&�A!�C� ��C�I,TV��6�ס)�h-J��-�p#=�r�S�U]�0�ާy��Pc���8� ��4�?��/���Wk	��?1���?q�np�N�Ok�^��,1���H	�N)!M�w�:�8 �'T$1��^be�u\>�<��٨3�Y��eE�h�ڼ!����1�-[vt��h�V��1�O���xR��S�����4��=ߠ�� �&��	!H���D�D���*�ǟ�j���+��7^����9D��K�@�9Xyrj�J p@ҁ��{���Dz�Ox�'��!�$,���K"�i�unZ+>����'l2�'��K�~
��?)G�۟d��Ѡ��}�00�i�3%�ph����0fy��Dc�d�Q�+�||lL@�M��;p�Q*q�}s ǂ�s�4��X7�֥:�"ת7 �؛�LL�jB�K>��Lğ	�훛wC�x�I�6J�43�i�++پ�Y�4�?!.Oy�;��<��?K�ū
�%j����=
�0���'�R�Wr��?q��Οx�OP����

:��H��䞍[t(zеi�2�m�(�$5?yF��M���?A��##�S-a7�p�#C9J���Ӧ���IG۟��	�XY`��4&��PȥG�@���"��J�d큡[q����C&fl��9�+�hO���SO� B�~	���D��c��
�� �P�3Ț�o�`Ee
��lT|�@,+�D�i��|"�@��?I#�i1�6��O���Q1>����5Y|���'����7M�O���6���O8�$�O�ʓ��h�ф�0Ks`��#ǯ@֢�ї�x�-�1 �b�|�'qR�M�B�m7���YP�Ŀv��$�[�P�SNA��MK��?���z0D���?��D�d� 3���,҆`1�e�"=;�iu�u��Cn���'&BW>�����2�V-5�L�	�e0+�",.d��a�f��h���RH����U�V�^��T}�W��F����#�O�Yq�'U�7��cy�����SR�/[k���:"�P���>����?1����O�����ī4�!bd�M6}�z%���DXҟTm�j���?�����X�0H���Q�C�>ak��B �M����?Y�%N�lX���?����?1����E,M�4ucb�P�M+�|!�,�\�@�o����O��?k\%��L_��0<al�>a�����Ý-�������|y���9Wh,���*�axB���-����-R'||�`
Ԅ��$��HB�	���?���~��6qA\�C��+�^��✞�M���?���?�7��|���?Ar��|�&�@�u��$RV�5<uBy�� �'��F�>�+O��O�bW��íQ;kIT��'ɘSPF�QFڿRp!S�D����IΟ��	3�uW�'|�5���P6�]	�(E84f��q>d�Ё&� '5@jM�i�Q�K'	��?�Gf��]��u�4eQ�t�6��j�Q����8'���N�[1�D�����*>Or��Prְy�o�4����-��6��O���F�ܴZ���P��^�T���1�E:����t�d�G�J�e�N!���7E�,�'��6��O�˓7ߪ�Q��i���'U�	ɬ#�$���/TI��H6������3���'�"�߉o���PKS����kr��%K����؉�Մ�!PAñ��%��=��k�v2�Pp
Lw���D��I�,��x��hfD�`���a)��eExR���?y��9V���"A�:Lɔ<��T��B�	4O0R7$M�Z�Pk�
	krJ���j~��a�|��AL%?uA[c�_��D�3s"�m���T��s��jW�@�r�'�%9D��$��H�f�2}y�P��t���g��#��S���Ny*��b>�"U�M@�(x@A��>�����B��hyw
�w1ԖQ���Y"�5N
ތ�'/�Sq���o���2<+�A�WZ(�	��J�$w�)�7^D<qD�J�h5�� �̓��h�
�'0��Ip.F�~e �Ĉ6��i؉��q�Os�҅N4�P	�.ԼY��0�qӢ���Op�[d��*H���D�O���O཭;�?�1/),���T,��K�`ˢQ�\�'Bnث�)���W*� 6�pdC#-�*_
m�'�p�
�@�UkV�N�� ����"x�bܕ'�2�_�azB�߂j�
t��XD�����y���..�t���~|xA(p���M#r�i>q$��CքI�粡��I��Z;�(�##O<v@5h��Zɟ��	П��I��u��',2�~��f&Ģ|G`�k�ǥD<�l0�s͢�c��L��KņA��?�ɗf�r�I!��$���+��P✴���t�P���.U�p�`���X�cm��G�W�6ɻ�ƌ,-���"l�r��7m�O���D�ܴ/
�	���U�H���$kl��ȓd~r����EF�ǆc�u�'�87M�O��%�tm�չi(�'��iФt�H�Ҁ*y��`�R+=ݛV	>{HB�'p�F�����T,�ԟ�q1�Ŝ��|�bBlM(g��di���'P0�yqu�"�|��l�Y��R���:\����H�]�Hz�)��	���F{��?Q��S�7��my��ȗLm��A5�K8N�C䉦ot�V�A�T�lH��L�e�r��Df~2�d��}aꞯ,Dfx��B(��$��N�xam՟`�IR�$�U��'k�u�e	G62�v�0�@�R$��l������Ob��g�eB�0�,H�l� 01�N�1�|���T�J"<E�T���V��ҿA!��A�@;A��?�$�|���B�l9�f� �y���Q�S�B�I�A7n�"���G~�4��K�F��#=i����[IJ����2	����.�B�Y�޴�?	�\��Vͅ��?��?���j5���Ok�"��PB��(8�^�K2Έ�X������K��Z�E*��8�6_>�8탽!ǉ'h�iel�g����F��<�d��a�nU0A L�[i�LKSH{���@�h�($�H��Bú1D����/ET�Y:�j�<)�C��p��ݟ��?�O�P�3�Q8v�l���u1~��'o���J@�ac�ѲFF�m�X�ܴ$���ꟼ�'����e�.�Lh5MT�XtT1{e!&H�(B�	�B|����QNyRbPs��C�ɲK��Fa�
:rd������#�B�)� �Ͳm�����b�P+t@�8�"O�����G����'(b�4���"O��+5g��U���À^dA�D��"O^%{"�#vB�Qi<I�u)r"Oz)���7Q5�`i��dr�A�"O�,#Չ�w��+h]�Q��"O̜��E�(*|�����FC 8	�"O�D�#� Dv��aᔑS�*���"O6@������ʰ`�"eRI�"O���L�&��
���">���k�"OL`d�Ğ3��tjd+�b䌬�&"O yc�wc*HItj��qv �"O�8jdb�Ne�����;Opr�`�"O�h�4����H�EO7a�F%��"O� �4o@�;ێqs4OQ�B��"O½Q.b�$�6�	���Y�"O���	�Ӯ�ʓ�Q�{��X��"O\,� ��:)H|�ȅ/Z1���@"O:$C����}j�a�vW�~�$8�"OP3�H�t���cdH�r�H��"O��rb�Ü,/��1��t@��"O|�`G"�'r��9�qm_*=���"2"O�9�6g&��!0r쉷y�f���"O������ɪPń\���Z�"OF��CHM�@�Ԅ�GZ6/���$"O&��uA��o�\\J��Ŋ�n�E"O89�-��F���¦!3�P�"O֬��$Å�.�4�B�F�

$"O�dSbΙ�q���Wg��B+�"Oa�h�?�>�`�%��} � 6"O�2g��=P5��WL��"O>iq��� ��C#C�!Flr��"O�A�`-�kfd`@�ȯT�t!�"O��Ȏ�f���F�,�ysW"Op�s��Z���	c��D4x�"OJܢSE��F�H#��!�&��"Oz}`�'T�\1�N� ��I��"O�����t�퐣�8F=�Y2@"O�8�c'��P��)�N�o��q"O��س@���|)R�2@��"b"O�`�c�ͮ��jBJgiڔ�$"OhQ�t�Y�(��iR	�;}.Jm�B"O���4�_:=����0��4"O��bI*_����R�0c�h�6"O��9!��S�^�X� �3td��d"O�tJ�c�4�>u�&�C:h�(�6"O�D�����v~���&$�!c�́b"O�x�)��8�U�T���c"ONp��(Q�N1�$�Mu�8K"O�I�i�2v�¬��	�<||�٤"O�I+͏z��YbȒ,#Pс�"O<�	�D�$\�j�H�(���"O D�G��F������?RY^�c6"O�mSQ雦Pq�`ȅ}T�8��"Ol=������v��(H���C�"OƕbP��:P�b�K��X���Q�"O�ZE�ȃS��Y6��&�����"O���B��?�:�2�mͫn��xP�"O(��D���vP��B�kڦ�"I�"O��Ҷ���e��9 >��S"O�bu�M:$�4�!��$&��jr"O�ɐP��}�0i��L�R/rp��"OĠ�֦N<V��R��3{>��u"O���V�EA'ب
�4'����"O� ^�[�,�!G٦8�6A�%S~U�"Oj�I��Ln*|�$!��DvRi��"O4xJaK�����UX�E�G"O��3*Q�1P�Ub�@	4"��9�"OV���G�� j�=���'֨��"OL�X')�\�T)
�$7R�hq� "OL��G�I��R�[�$�5u'&15"On}��� r4�a��+�+��W"Oh�;@�M���Bԉ_�Jy��t"Op��EK�>�U�sS�`�]�`"O���G�X1h����5�֐\��E�W"O^5�R�,D���'(H�M��P�"O�`j�g�K.��/��{eNlJ�"O�a� T��XD��K8VPÆ"O�eӄ�J�WG9��j�ؐ-C�"O��"b8i�zJ��M�.�(홂"O&��"�W�L�[aƌ e>�2e"O
qXp��E�R����G�m�|�"�"O����	g����[�x���"Oz��cJ�D$��a�,L�y��"OF����T47����ٌ2�f��"OЁ�oM �`s�m�F�2"O�hc0#�i��������X�p�"O^ȢG�B�z��UJD�5l@�"Ov��#L�%U�����,n���"O���$n@�S�.hJE��	����"O����L��
�)�3T�0�U"On�Q'i�;8h��ʎ\\=�"O(pj�lC��) *�
Q�\�"O���Qjf0S'��6���s�"On���f��C
��[q�X�4�D�3"O����*�K���h�.A�� Ӧ"ODeH$�@����D��!�< T"OH�g�
�e�:��2�B �`h�"Oh�Ґ�`V��xf�T�ft��"O��;�b���<�A��>�H�"O�U2����z�Z%N�Z3E"O@�3�Ԛ�$�v�T�^�\PF"OZd���˲q3b4��ID�#��p"Ot����L�CZ�4�Qhθ%4P��"O��RH�	 ��:@�
ۀ�Jd"O^ �i�WF@}��ٛ1N���"O��[4C�; ��Z��@M+1�"Od%{��H�<#ݡS'�t)�hk�"O�a⮟�&٤�X�#dz��� "O�Qb�V�J��}v���"Ot� �����t��d�eW؉*E"O���#N�ly�����K0b��:�"Ozh+�To�2����	7>`�:"O�9pa��o��
���6!��:�"OɈ��luL���-/�x:"O̡sUĜ��8���>U�l	�Q"O�qɥf�5<�
��f	�=�1Qr"O\��ࠎ`��;g����Y!0"ON1&Ǟ�@K�nB�)H�xv"O,�q��R��p�'�_��X�a�"O ��N� r�ԡ��,H-Q��@B`"O�ꗏʵQ�������(�>iR�"Om���CQ��Yy3���F��$j�"OR�W����:�z��,$6@��5"O&Ի6�O�\����E\$�"Ov*�I�;z��y
$�Q�/|���"O������U�¡<B��"OHM����F���	�b�s��X�"O� ��`�-��3f (��		"��"O����]�%��M��,1Ţ��"Oc�f�OM�lP��u{�"Op1:B̓�]�,��̋�VP�hh�"O05ATF�^�����D�D����$"O��!eY59��x��l*�l��"O:h���=&D��ش���[�b�Ғ"O����oξ~x�x�-�3@�"O�8@�M�4(F�eIvc߭g�<�i�"OPb�FS�F,]��,�;Z�ț�"OP�s�a��W��$��4��Q(!"Ojɒ���(����0�^�x3"OੰĈ�r���Ca�.��H[u"O���r N���$���&�@��"O�@r�
;�y�<m޲�X"O�����N��̂��&`X��B"O������,zL$���+�",B�c�"Oqqr���H�P0�R*�V!�!K�"O�P`F�˷He��	��!h"Oppc%O5?��3�(��	�m$"O^�DH=>�rk��Ղ#�M"O>}�'_�t���M� $����t"O,���oǆE05��7Y.<�Kd"OĴ�pE
�~m$)�`_?9��Qɑ"O��q�aQRs,�:�@ݮww���"O �)rgWO��x�A�([o&D�5"O�q��mU-6����@��4�S"OH��J8}�6��@eF�j
�(��"OШ*rB��?��s�E�)ռ�J�"O6����L�l��󋌄.pN43�"O�a2J+"�q�$뜇Cn�sw"O�5(��=.rL�kc ��H�T8�"O���M�9z�����N+~Z����"Op`�7��"-L��B��U�e�2"O�IxE�,��0�H@I���"O�5��
5#�<��AT�.��ٛ�"O����աz�+�Nu�E���}�<ђ#�zͺ�k�,���u�� �v�<��iX0�<�3��w�.��6�~�<9V�͜x����E䍗\L����y�<�ЍQ.[�1Q��S>i��!Y�Nw�<���=Q���+�a�c�>��"�N�<����;9H� p��
cf-���^I�<A!F�0	�ͩ�]5$��l��EE�<q�ƎQ�AC�Ǝ�A'\2�$�K�<��^�*pm��#�W������I�<)�٦b!����@}�z�{��
B�<9b���=�b��i	/U��$[�<4�^0}2�U ��
�	(�@�֩V�<A��I,F�����N4Ag��� �o�<��4����`^� ��ȑ��h�<y��h-Ҥ��� � �I�M�<i�A��)v�-�A���_��E)5�[b�<����5#�R�*a��:��Q���|�<� ��(b
:�"��]�IPL�	��_�<���dE����(\�"���X`�<a��+�tz�e�/�(�T�g�<�i�!g=��Z�ןI��2V.�a�<��!Ȧ̄<��m���!�-�U�<W�ج}�T](��[�'�5yC�L�<y�	�n�TA���T�z%�!��J�<9!��@1�`B�(�>	��HB�<�6�Ōos����7�E 	I�<Y� �F��ѐ�&Q�p��2P��`�<� 8�cЭu�rP��	�p� �@�'@hq�)N�+]���%�>a�4�u,_�pB�ɋR$ ����r�9���6 �B�	)P��
R�{�`DC�F�$}bB�	!g��j�Ԅ���b��lx�C�I�l�DQ7�QpwĠ��J�="m�B䉉�zi��/=��H�W���C�� a�@��4L�S��h"��)�lC��2G��C�R5@Y�pВ(
>6|B�	7 �l%��J�#Y<@tIӣ�8ۦB�9f�@3��,[�:t;R�A��B�;keH ��'�/}fM��N��H|C�I
.��r�Ů)&���$	�xzC�	~�P�+���&�Xx����i�"C��Xu���;1�8:�둮= C䉃kT�q G"�.n����
Ѡ4��C�ɧG��(Ԫ�p9���&O)z�.B�� ��<٧H��u��� )3�B�ɬF��z�"[f��I��
�9��C�IO�����ŰuH� z2��<��C䉑��:��	:j�H2���x�C�ɩ��{�,�,Tv�`F�=�HC�IdLn�*���<=�UG�Y��B�I�rVp� W�s�R�!��Z��B��+2��`��W�>4"����ߚB�ɪe:@	1󉇂r�,��悗}vzB䉜>��e8D[�Z6�
 :<B�Ik��#�H�@��Ȇj�vB��A�x@��Y6u��<��.��4�tB�	
h��'@N�}g
\�/sdB�I�2�ͫc.GoĲA�PCB;,�FB�I�,o��a�� �4�����h��aB��sۮe��a��悽�5ȑ�tO�C��6|�>�"����I3��*��C�	2gE,x��,��?vTm�҉�	QN�C�I�CH�a^�+�U꤮�=�C�&H$2Q���÷��y��Iѫ.ŸC�%T�x5��LEe���J�0�%"O����C�~�F�N& g�Q@s"O����W4�Iw�8qLz�á"Oę'��>53���� �e <Y`�"O$����fq`p�`ռb�°*�"O�@�哚@t�$ɕeY/�Ȍ�2"O�H+�'G�p���
$`���"O�5���SZ�6٨aB�r�le�"O�TأgқX��i��F-֪�B�"O�a(��_z�}I��;n����"Or(9�퇊Up�i�����\ݲU"O�4���0��@m��'ى�y�e�&�u�D�4E��y
LL:�͐�
PQ$+ޓ�y�$3��lz +M�x��/ݽ�y���;Yx2��B��[^ňbiǒ�y�"*p +��F0�Jw"B��yr�H?>�����N�H�F���yb)�o�ƹ�׀�r���$�y����w�D8�↊��d�q�k�yR+Ey<Z�{ ��H�>����yb�Q#Z���o��V�����܇�y��+;��\��Hŀ{۪A���D �ybf���\*Ư�($`y�VD�$�y�Yd�����"�@9k�(��yb�A<:fd��RJ�\q�����I��y�К��	C��
�=R(�� ɤ�y
� ��ðF��?���)眡x��9Q"O���HĻX!*E�J	�r���"O�-A���"o�Ri�7@�i
"O���f��4�|���%Ḝ2"O>��6�1	|f��"���("!"O@�J�'��xvZ$��j	�V"O��CŌ�?����C��s��i�e"O&�r �ˮ��:��@�����"Oqam\�j���qW��'��E
�"O���4MK3@ܠ��a�G��T�0��W���Ӗ5�L����_K���$�JC�	( ,�9��*A�t���㒷3�\dG{��9O��R�(�m�Z̛ÇͤQw�lP�"O�P��͘�dP���D�!42i�2"OhњWJ�]FR��$&\E��-A�"O����� 4XyK��BY߶�r�"O� [`A^�p"B��]�����(D�t�&�!e�|��S˂�E��fB�	�S-�	�b�A���0W�M�liTB�	�:l-�V
�.�z �S���$BB�ɽd�����%BoZ<�#�C��C�ɠu�0L�f��)Г�Y�*C��/�HK�e����m	��4�TB�Ɇn�.|��
.Z����+��oq|C�ɭ>����;U����N� JC��30qD(T!Ƚ=��=Äϡyt��D�Pf2-���F�|�cS��g!��?S�l(S�A��0�.l�-�Ic!�A5֘i�j���RG'��U�!��u�者K�]��%���j�!� �fQ�%��
z��C�dU 2�!�Ǆ.^��µO��|2���a�1M=!��\�ld4t+�ᖿu�Y��Ũ�!�B�8�@0s鏳MO��a�A�Q!�$�1/'V)��m�587։�����O!�ĆI�� *ݮ2��tU���7H�B��0l�tG]�y�x��E,�C�I+/�pht�!����į/dC�I/(VJd3��e�H���ܒB�I�Xd�Q�`��!I#-X?'s�B�I� ��p �*��� �$�<	evB��6AHb�c$b]+I���P�^�?�2C�	&q�Ld`��X)B)2Y9��14:NC�I�l�.��QOW G"*2%H���C�	*k�$u㶦�?	�h���ϰC�I�};�� r�Дe3H)s"͌"KܔC�I�A��ڤNF�xE<e<�B�I�J���b�+V!^�ǧ	H}TC�ɔ�t����^�F�"9Y	ta(C�Il+5#�$ӹ@yP���gZ��B�'&���� ��},4!@�[/'�B�	 Bq�E��y�����l�r�C䉅%��!����%��z��8C��;o|�=���Y7Д���C�w��<�a$O��0�a��3FF�z0b�E�`Y�p"O=#2'õ;�& �¡�$.,�(�ȑ/!�$�6@�`���15艙��U�O{�z�CQ�$�Ò��V�)����S�"��ȓ� Fo��TW�%�G��<�=y0�*�S�rl"��5��/pv,�S���E?�B��j ���1�-C�&a����d"=��'d��Xg�M&YF�]��l�8�"O��A Ʒ�t���n��f´�
ԹiS��	�|�(��w� W�r���H��A ��$3�)� ^�ل�ޱ~��J=h09b6"ONa"�-P��LQrj�;DL,-���?�S�9L��2�A��$!y��+3�*B�ɧz:��sK��%#g. [�B䉔<.��:���cQ]�eS-LN�B�	�{VT��bgņ�DY�V�MtXB�IA�8�S�5$�nщh��clB䉔V4���"I).�$��Ҥ�S�fB�	]���W'�</D��6��5<B�ɇ.(�@�H@��a]rg"B��4')�K�	7��(�q�M�B�ɨH:M�`����P�$#L �B�w�^��R�N8k��}�/�>!pB�7}����mJG
�١���g/JB���J�따<��C6-V�g$B�eC.�r����٣�&��s�B�ɩ`�R����qǞu����r
B䉮CJ�xt5�R��U�'E�B��$\�(tՄ�H������5�B��'�d��ۄ�D�d���h0NC��bNѡT�]�8:��̏�p\C�	�Y�EU!.Z	��۪\�C�I�P��ሗ�C�;�,�#EJ4�C��'16� 3F��1{(ً��X��C�ɼ}hd�8�M�yC9�����C�6D�}2�L�`�<\�a#�t�LC�Ɂu�����KȠr�2�S���*E�NB䉗 xT,ٲ	I9�,hp��=3�&B�I*\�Ⱥ�c�&���� '�bC�I�b��a9$��&��!�M�NfbC�	�2�L4	�O�D���jq�W�T�\C�I��.T��.�(�z�gԧSuC�	<�|�v��$T���u�O�r��B�	�z�5j�G�L�b��2���B�I�`���z� � 3X�@���zk�B�Sr���g̠T�.4)u�Βy�B�	K%�:V��Mw��b�-@�>̀B�;^ĵ�KK��}�" /Y�NB�	�t��Á@P��v-p�G���B�	%4�l��X�x� ���TTrC�	x���04.îP�}(�
!�RC�#20���A�?�����H�
L^C�	�4TXp�� �.M>��١Cƨ&xFC�1GH��!!�G�h��'΅�C�
�.�2��X8d�0�1G}N�B䉴?����΀:�Ԓtn��?}B�	^�^�k�/R�j]z���<�C�ɔ^4�e�(c/�)�p��{��B��
|�"�:��H�P}j� Ī�*T�vB�Ʉ����Ъ�?�^��(��r�pB�I�M�=��H;S+�������(B�R}.T����k��e�uC<� B��+v���9�؏~����`�Vd�C�	 (�D�Q�d�"6�F1���JT�B䉘U<�<���ו|&us��J*�C䉪J��IaR���v���:�B0szC�ɐ#�T��NW�p�\9ǋ��C�B�*]�� !��
���p����2C�%�U`�e� E�f񋵤֨]s^C�I�t)�͛FCtI`y*�h�H��C�	,}
��@T暜n�`e���_Z�C�ɉP��T��"�
@�J-���=N��D��-j�D(�bL�g>��eO��!�?Z��a�`dA,
5\d���'P�!�� >��MQ�_`����ӑ.=�K�"OP�Ӧo����w�l>���"Oj�X�ٴZ  �B���V&jq�"O�		Gk�)�-B��"\�t"O!T
�����ϔ3�q��"O,Ѡg�  �      Ĵ���	��Z�$I7=���C���NNT�D��e�2Tx��ƕ	#��4"�V���$�f��m�tT^�0"�6;�2�#J9̲�A�e%g����lS��M��'�:���R4{�ͭ�F>>aI��'�Fxb��G#}e>`�u.�D��٠���?"�^��g�Iy�����K?}R�[1$�1�T�>o�L�wED�ʤA�� �(_��'ޤ���	?s�h�/O���ǀI�;m��@�V�P*� WU�0�/�4ֆ�X�R�Gˎ�W�0��Zf &WT���=}�m1dӒDۃ���ʵ��pW�<�f�J�=*"Q�'��)c�X0V�''�;�f+�I�>���%]�� U�G&n���@�PL�z�$�$	0w��4�q�;�i!+8 �kB3a�8C��Y�R�%5�4� �'+�`�G΀���O>bcA���P�KӥيZ���F���L'�h1��Q'VPZ(�N��#�9L�<��?OR���"2�(���e�'��!qd�'K�U�S+����S~�a˛h��l%� T�PYP2�zOYq��+#��M
M�DS�4+���<	�O����@:G�V垯|��IƧıM?"�C_���$�)�(Ȕ�|��K�i"| L�����O�6 ��NR�6t�f�9sZa�1N�d?�1O�D)e���ԟ��jtb��l�����>�4�'-ר�x�8J>A���&yL�$�8!U��/8z�I):52)��!>�⸣R�Q�_?,�;��a6�O�O�A�+��gj� ���4P~	��O�<����T�ē6|H��n_T����u`�+��B:����68�yrO�>0�$j�/�-oY��k�'�fŃ3�;[����ɻm��(�w��9G��X�LA�nt˓+���c�u�t�%)b=�d	
x�Q�3i�F�E�Z�\�b�j f�'8
E�kV���'Җ0�*�Z�n���֖����k��5!�d[�v �  ��:�x�bM�o�,���z�T�5J��	��T��S�P�Ue*�#&�P6S;@�	e����8o$���sh�)q�칓@(���$L�CO"�=lO�tqkL�^���	X8(ur�;G"O��n�S���t�E�P0\x��Nf���\���k�Ovy��h�iFN L��u��R�i�O���O����t���O�B�LMXr��
�xyJ�J�)��hG�ڤi�����<$�l(��i͘z7��*Y�(   !
  t  �  �   @'  �-  �3  >:  �:   Ĵ���	����Zv)���P���L_zD�R���\��Tx��ƕ	#�e&�T���Y�k��(kw�,{�bHA��$D�<RG�]�QYh�@�3���*�K�!pO�!he�Tm��a�1ɨ��I����@z pg�9��\jI�/lw�� !�^	!�BY���Ǭ[�<14�,> E�!��>MSV�uN�O8	a��U��9su�¦O�Z�X�#�0p��`�+4��JH-4�t��SI�!5��� RA�v����>���'0��'�v���wA�3<BI����j�vp��cM=��D�3 ��|B@�)<�
��!jG9a�bH�%����N�+��|r��y���3���=a`�%eΓ��$�'��H4LO��qA�!�޴`��W��@b�"O ��O�rG� ��	���׿i�
"=ͧ��"l��˱�ůxH���②yc0�CC�M�O0�Ȃ��?���?U������Ol��0U��D߁<�X�G&ͩU�zݰ�	�?��q���"�J��&|��t�VBޒeY�	[�ra����[�rg2�Ϳ�2!�$��',� 1�Ŷ7NtC�I�@(j"��<�&d)҆�E��B�	;����c��!j��C Ðk���ʛ��|bL��7M�O��?���
�-	�(�,I���D�tӺE ��O��OH�+�'�Oc���HC̲��߽a���`D/�Q8�=�v��I�O��)���o�rX'ǋ�6X�0���d��n��9�'A��K��Bր@��B�s�u��u����E#6�����K��6r<��I�����9�6�A �>Ow,@��{��I0;�J�۴�?q���I�,%�`���O$�d�00�Y�7�ϙQ�̄21D��-������<���'j�y�AK����[�Q�I�zeZ��iltGx���h�%h`V�Fm�E�u���"��[�`Rn9���6
�����̉E�@Mk`AKAD.��9>��DiΨg���K�	�<Q�v�EzB�1�'O���0�bA%��٢d��'D�=y��i��'nx���5!���'J��'��T��5���8�(]�N�k6@I0����V�|2⎺_��m��
JB��UeФ��d�0	�|��
�W��x��C�w���(�
�;���3_��2LO�LЂF2P`lX�m�&M4��"O؈���T`��8d�$A�(�6�i�"=�'��Eע���O�&=;���#�A�E��i0ӡC3��X����?y��?�"����$�O��95|�$Ύl{����F�$�	�`@[������l���	'[�AK1I��;�z����.04���.62��r#<�iT�R=.���a��_-eA�B�ɴU=�E����%y_"yP'�C�	p���q,L�M����rkC�����'�ܹt��͟0��矤����ԩ�e��A"��׹��Al�Xi�`���|�I�+^*�IV�S�O��$�+��J�eW*P� �Lj�'��]����#<��L��P�p�]Y��Ŗ'Iў8A���OrG�toZ:G<����{d: ����yč9/� ʒ�t����˓��>�$���2�I�lR��E��4��U�E��>����6����'��]>!�c�L����?55N����_�M6�ULH�u�t%��48�MJ��Ü�R��O�\�')�V�s��VE���:�E�!3Q���T���P���S݈P2�e]��F��nѺ:���A+͠]wz��%$��K��?�A�|����Dߪ0h��	�
&�A!�C� ��C�I,TV��6�ס)�h-J��-�p#=�r�S�U]�0�ާy��Pc���8� ��4�?��/���Wk	��?1���?q�np�N�Ok�^��,1���H	�N)!M�w�:�8 �'T$1��^be�u\>�<��٨3�Y��eE�h�ڼ!����1�-[vt��h�V��1�O���xR��S�����4��=ߠ�� �&��	!H���D�D���*�ǟ�j���+��7^����9D��K�@�9Xyrj�J p@ҁ��{���Dz�Ox�'��!�$,���K"�i�unZ+>����'l2�'��K�~
��?)G�۟d��Ѡ��}�00�i�3%�ph����0fy��Dc�d�Q�+�||lL@�M��;p�Q*q�}s ǂ�s�4��X7�֥:�"ת7 �؛�LL�jB�K>��Lğ	�훛wC�x�I�6J�43�i�++پ�Y�4�?!.Oy�;��<��?K�ū
�%j����=
�0���'�R�Wr��?q��Οx�OP����

:��H��䞍[t(zеi�2�m�(�$5?yF��M���?A��##�S-a7�p�#C9J���Ӧ���IG۟��	�XY`��4&��PȥG�@���"��J�d큡[q����C&fl��9�+�hO���SO� B�~	���D��c��
�� �P�3Ț�o�`Ee
��lT|�@,+�D�i��|"�@��?I#�i1�6��O���Q1>����5Y|���'����7M�O���6���O8�$�O�ʓ��h�ф�0Ks`��#ǯ@֢�ї�x�-�1 �b�|�'qR�M�B�m7���YP�Ŀv��$�[�P�SNA��MK��?���z0D���?��D�d� 3���,҆`1�e�"=;�iu�u��Cn���'&BW>�����2�V-5�L�	�e0+�",.d��a�f��h���RH����U�V�^��T}�W��F����#�O�Yq�'U�7��cy�����SR�/[k���:"�P���>����?1����O�����ī4�!bd�M6}�z%���DXҟTm�j���?�����X�0H���Q�C�>ak��B �M����?Y�%N�lX���?����?1����E,M�4ucb�P�M+�|!�,�\�@�o����O��?k\%��L_��0<al�>a�����Ý-�������|y���9Wh,���*�axB���-����-R'||�`
Ԅ��$��HB�	���?���~��6qA\�C��+�^��✞�M���?���?�7��|���?Ar��|�&�@�u��$RV�5<uBy�� �'��F�>�+O��O�bW��íQ;kIT��'ɘSPF�QFڿRp!S�D����IΟ��	3�uW�'|�5���P6�]	�(E84f��q>d�Ё&� '5@jM�i�Q�K'	��?�Gf��]��u�4eQ�t�6��j�Q����8'���N�[1�D�����*>Or��Prְy�o�4����-��6��O���F�ܴZ���P��^�T���1�E:����t�d�G�J�e�N!���7E�,�'��6��O�˓7ߪ�Q��i���'U�	ɬ#�$���/TI��H6������3���'�"�߉o���PKS����kr��%K����؉�Մ�!PAñ��%��=��k�v2�Pp
Lw���D��I�,��x��hfD�`���a)��eExR���?y��9V���"A�:Lɔ<��T��B�	4O0R7$M�Z�Pk�
	krJ���j~��a�|��AL%?uA[c�_��D�3s"�m���T��s��jW�@�r�'�%9D��$��H�f�2}y�P��t���g��#��S���Ny*��b>�"U�M@�(x@A��>�����B��hyw
�w1ԖQ���Y"�5N
ތ�'/�Sq���o���2<+�A�WZ(�	��J�$w�)�7^D<qD�J�h5�� �̓��h�
�'0��Ip.F�~e �Ĉ6��i؉��q�Os�҅N4�P	�.ԼY��0�qӢ���Op�[d��*H���D�O���O཭;�?�1/),���T,��K�`ˢQ�\�'Bnث�)���W*� 6�pdC#-�*_
m�'�p�
�@�UkV�N�� ����"x�bܕ'�2�_�azB�߂j�
t��XD�����y���..�t���~|xA(p���M#r�i>q$��CքI�粡��I��Z;�(�##O<v@5h��Zɟ��	П��I��u��',2�~��f&Ģ|G`�k�ǥD<�l0�s͢�c��L��KņA��?�ɗf�r�I!��$���+��P✴���t�P���.U�p�`���X�cm��G�W�6ɻ�ƌ,-���"l�r��7m�O���D�ܴ/
�	���U�H���$kl��ȓd~r����EF�ǆc�u�'�87M�O��%�tm�չi(�'��iФt�H�Ҁ*y��`�R+=ݛV	>{HB�'p�F�����T,�ԟ�q1�Ŝ��|�bBlM(g��di���'P0�yqu�"�|��l�Y��R���:\����H�]�Hz�)��	���F{��?Q��S�7��my��ȗLm��A5�K8N�C䉦ot�V�A�T�lH��L�e�r��Df~2�d��}aꞯ,Dfx��B(��$��N�xam՟`�IR�$�U��'k�u�e	G62�v�0�@�R$��l������Ob��g�eB�0�,H�l� 01�N�1�|���T�J"<E�T���V��ҿA!��A�@;A��?�$�|���B�l9�f� �y���Q�S�B�I�A7n�"���G~�4��K�F��#=i����[IJ����2	����.�B�Y�޴�?	�\��Vͅ��?��?���j5���Ok�"��PB��(8�^�K2Έ�X������K��Z�E*��8�6_>�8탽!ǉ'h�iel�g����F��<�d��a�nU0A L�[i�LKSH{���@�h�($�H��Bú1D����/ET�Y:�j�<)�C��p��ݟ��?�O�P�3�Q8v�l���u1~��'o���J@�ac�ѲFF�m�X�ܴ$���ꟼ�'����e�.�Lh5MT�XtT1{e!&H�(B�	�B|����QNyRbPs��C�ɲK��Fa�
:rd������#�B�)� �Ͳm�����b�P+t@�8�"O�����G����'(b�4���"O��+5g��U���À^dA�D��"O^%{"�#vB�Qi<I�u)r"Oz)���7Q5�`i��dr�A�"O�,#Չ�w��+h]�Q��"O̜��E�(*|�����FC 8	�"O�D�#� Dv��aᔑS�*���"O6@������ʰ`�"eRI�"O���L�&��
���">���k�"OL`d�Ğ3��tjd+�b䌬�&"O yc�wc*HItj��qv �"O�8jdb�Ne�����;Opr�`�"O�h�4����H�EO7a�F%��"O� �4o@�;ێqs4OQ�B��"O½Q.b�$�6�	���Y�"O���	�Ӯ�ʓ�Q�{��X��"O\,� ��:)H|�ȅ/Z1���@"O:$C����}j�a�vW�~�$8�"OP3�H�t���cdH�r�H��"O��rb�Ü,/��1��t@��"O|�`G"�'r��9�qm_*=���"2"O�9�6g&��!0r쉷y�f���"O������ɪPń\���Z�"OF��CHM�@�Ԅ�GZ6/���$"O&��uA��o�\\J��Ŋ�n�E"O89�-��F���¦!3�P�"O֬��$Å�.�4�B�F�

$"O�dSbΙ�q���Wg��B+�"Oa�h�?�>�`�%��} � 6"O�2g��=P5��WL��"O>iq��� ��C#C�!Flr��"O�A�`-�kfd`@�ȯT�t!�"O��Ȏ�f���F�,�ysW"Op�s��Z���	c��D4x�"OJܢSE��F�H#��!�&��"Oz}`�'T�\1�N� ��I��"O�����t�퐣�8F=�Y2@"O�8�c'��P��)�N�o��q"O��س@���|)R�2@��"b"O�`�c�ͮ��jBJgiڔ�$"OhQ�t�Y�(��iR	�;}.Jm�B"O���4�_:=����0��4"O��bI*_����R�0c�h�6"O��9!��S�^�X� �3td��d"O�tJ�c�4�>u�&�C:h�(�6"O�D�����v~���&$�!c�́b"O�x�)��8�U�T���c"ONp��(Q�N1�$�Mu�8K"O�I�i�2v�¬��	�<||�٤"O�I+͏z��YbȒ,#Pс�"O<�	�D�$\�j�H�(���"O D�G��F������?RY^�c6"O�mSQ雦Pq�`ȅ}T�8��"Ol=������v��(H���C�"OƕbP��:P�b�K��X���Q�"O�ZE�ȃS��Y6��&�����"O���B��?�:�2�mͫn��xP�"O(��D���vP��B�kڦ�"I�"O��Ҷ���e��9 >��S"O�bu�M:$�4�!��$&��jr"O�ɐP��}�0i��L�R/rp��"OĠ�֦N<V��R��3{>��u"O���V�EA'ب
�4'����"O� ^�[�,�!G٦8�6A�%S~U�"Oj�I��Ln*|�$!��DvRi��"O4xJaK�����UX�E�G"O��3*Q�1P�Ub�@	4"��9�"OV���G�� j�=���'֨��"OL�X')�\�T)
�$7R�hq� "OL��G�I��R�[�$�5u'&15"On}��� r4�a��+�+��W"Oh�;@�M���Bԉ_�Jy��t"Op��EK�>�U�sS�`�]�`"O���G�X1h����5�֐\��E�W"O^5�R�,D���'(H�M��P�"O�`j�g�K.��/��{eNlJ�"O�a� T��XD��K8VPÆ"O�eӄ�J�WG9��j�ؐ-C�"O��"b8i�zJ��M�.�(홂"O&��"�W�L�[aƌ e>�2e"O
qXp��E�R����G�m�|�"�"O����	g����[�x���"Oz��cJ�D$��a�,L�y��"OF����T47����ٌ2�f��"OЁ�oM �`s�m�F�2"O�hc0#�i��������X�p�"O^ȢG�B�z��UJD�5l@�"Ov��#L�%U�����,n���"O���$n@�S�.hJE��	����"O����L��
�)�3T�0�U"On�Q'i�;8h��ʎ\\=�"O(pj�lC��) *�
Q�\�"O���Qjf0S'��6���s�"On���f��C
��[q�X�4�D�3"O����*�K���h�.A�� Ӧ"ODeH$�@����D��!�< T"OH�g�
�e�:��2�B �`h�"Oh�Ґ�`V��xf�T�ft��"O��;�b���<�A��>�H�"O�U2����z�Z%N�Z3E"O@�3�Ԛ�$�v�T�^�\PF"OZd���˲q3b4��ID�#��p"Ot����L�CZ�4�Qhθ%4P��"O��RH�	 ��:@�
ۀ�Jd"O^ �i�WF@}��ٛ1N���"O��[4C�; ��Z��@M+1�"Od%{��H�<#ݡS'�t)�hk�"O�a⮟�&٤�X�#dz��� "O�Qb�V�J��}v���"Ot� �����t��d�eW؉*E"O���#N�ly�����K0b��:�"Ozh+�To�2����	7>`�:"O�9pa��o��
���6!��:�"OɈ��luL���-/�x:"O̡sUĜ��8���>U�l	�Q"O�qɥf�5<�
��f	�=�1Qr"O\��ࠎ`��;g����Y!0"ON1&Ǟ�@K�nB�)H�xv"O,�q��R��p�'�_��X�a�"O ��N� r�ԡ��,H-Q��@B`"O�ꗏʵQ�������(�>iR�"Om���CQ��Yy3���F��$j�"OR�W����:�z��,$6@��5"O&Ի6�O�\����E\$�"Ov*�I�;z��y
$�Q�/|���"O������U�¡<B��"OHM����F���	�b�s��X�"O� ��`�-��3f (��		"��"O����]�%��M��,1Ţ��"Oc�f�OM�lP��u{�"Op1:B̓�]�,��̋�VP�hh�"O05ATF�^�����D�D����$"O��!eY59��x��l*�l��"O:h���=&D��ش���[�b�Ғ"O����oξ~x�x�-�3@�"O�8@�M�4(F�eIvc߭g�<�i�"OPb�FS�F,]��,�;Z�ț�"OP�s�a��W��$��4��Q(!"Ojɒ���(����0�^�x3"OੰĈ�r���Ca�.��H[u"O���r N���$���&�@��"O�@r�
;�y�<m޲�X"O�����N��̂��&`X��B"O������,zL$���+�",B�c�"Oqqr���H�P0�R*�V!�!K�"O�P`F�˷He��	��!h"Oppc%O5?��3�(��	�m$"O^�DH=>�rk��Ղ#�M"O>}�'_�t���M� $����t"O,���oǆE05��7Y.<�Kd"OĴ�pE
�~m$)�`_?9��Qɑ"O��q�aQRs,�:�@ݮww���"O �)rgWO��x�A�([o&D�5"O�q��mU-6����@��4�S"OH��J8}�6��@eF�j
�(��"OШ*rB��?��s�E�)ռ�J�"O6����L�l��󋌄.pN43�"O�a2J+"�q�$뜇Cn�sw"O�5(��=.rL�kc ��H�T8�"O���M�9z�����N+~Z����"Op`�7��"-L��B��U�e�2"O�IxE�,��0�H@I���"O�5��
5#�<��AT�.��ٛ�"O����աz�+�Nu�E���}�<ђ#�zͺ�k�,���u�� �v�<��iX0�<�3��w�.��6�~�<9V�͜x����E䍗\L����y�<�ЍQ.[�1Q��S>i��!Y�Nw�<���=Q���+�a�c�>��"�N�<����;9H� p��
cf-���^I�<A!F�0	�ͩ�]5$��l��EE�<q�ƎQ�AC�Ǝ�A'\2�$�K�<��^�*pm��#�W������I�<)�٦b!����@}�z�{��
B�<9b���=�b��i	/U��$[�<4�^0}2�U ��
�	(�@�֩V�<A��I,F�����N4Ag��� �o�<��4����`^� ��ȑ��h�<y��h-Ҥ��� � �I�M�<i�A��)v�-�A���_��E)5�[b�<����5#�R�*a��:��Q���|�<� ��(b
:�"��]�IPL�	��_�<���dE����(\�"���X`�<a��+�tz�e�/�(�T�g�<�i�!g=��Z�ןI��2V.�a�<��!Ȧ̄<��m���!�-�U�<W�ج}�T](��[�'�5yC�L�<y�	�n�TA���T�z%�!��J�<9!��@1�`B�(�>	��HB�<�6�Ōos����7�E 	I�<Y� �F��ѐ�&Q�p��2P��`�<� 8�cЭu�rP��	�p� �@�'@hq�)N�+]���%�>a�4�u,_�pB�ɋR$ ����r�9���6 �B�	)P��
R�{�`DC�F�$}bB�	!g��j�Ԅ���b��lx�C�I�l�DQ7�QpwĠ��J�="m�B䉉�zi��/=��H�W���C�� a�@��4L�S��h"��)�lC��2G��C�R5@Y�pВ(
>6|B�	7 �l%��J�#Y<@tIӣ�8ۦB�9f�@3��,[�:t;R�A��B�;keH ��'�/}fM��N��H|C�I
.��r�Ů)&���$	�xzC�	~�P�+���&�Xx����i�"C��Xu���;1�8:�둮= C䉃kT�q G"�.n����
Ѡ4��C�ɧG��(Ԫ�p9���&O)z�.B�� ��<٧H��u��� )3�B�ɬF��z�"[f��I��
�9��C�IO�����ŰuH� z2��<��C䉑��:��	:j�H2���x�C�ɩ��{�,�,Tv�`F�=�HC�IdLn�*���<=�UG�Y��B�I�rVp� W�s�R�!��Z��B��+2��`��W�>4"����ߚB�ɪe:@	1󉇂r�,��悗}vzB䉜>��e8D[�Z6�
 :<B�Ik��#�H�@��Ȇj�vB��A�x@��Y6u��<��.��4�tB�	
h��'@N�}g
\�/sdB�I�2�ͫc.GoĲA�PCB;,�FB�I�,o��a�� �4�����h��aB��sۮe��a��悽�5ȑ�tO�C��6|�>�"����I3��*��C�	2gE,x��,��?vTm�҉�	QN�C�I�CH�a^�+�U꤮�=�C�&H$2Q���÷��y��Iѫ.ŸC�%T�x5��LEe���J�0�%"O����C�~�F�N& g�Q@s"O����W4�Iw�8qLz�á"Oę'��>53���� �e <Y`�"O$����fq`p�`ռb�°*�"O�@�哚@t�$ɕeY/�Ȍ�2"O�H+�'G�p���
$`���"O�5���SZ�6٨aB�r�le�"O�TأgқX��i��F-֪�B�"O�a(��_z�}I��;n����"Or(9�퇊Up�i�����\ݲU"O�4���0��@m��'ى�y�e�&�u�D�4E��y
LL:�͐�
PQ$+ޓ�y�$3��lz +M�x��/ݽ�y���;Yx2��B��[^ňbiǒ�y�"*p +��F0�Jw"B��yr�H?>�����N�H�F���yb)�o�ƹ�׀�r���$�y����w�D8�↊��d�q�k�yR+Ey<Z�{ ��H�>����yb�Q#Z���o��V�����܇�y��+;��\��Hŀ{۪A���D �ybf���\*Ư�($`y�VD�$�y�Yd�����"�@9k�(��yb�A<:fd��RJ�\q�����I��y�К��	C��
�=R(�� ɤ�y
� ��ðF��?���)眡x��9Q"O���HĻX!*E�J	�r���"O�-A���"o�Ri�7@�i
"O���f��4�|���%Ḝ2"O>��6�1	|f��"���("!"O@�J�'��xvZ$��j	�V"O��CŌ�?����C��s��i�e"O&�r �ˮ��:��@�����"Oqam\�j���qW��'��E
�"O���4MK3@ܠ��a�G��T�0��W���Ӗ5�L����_K���$�JC�	( ,�9��*A�t���㒷3�\dG{��9O��R�(�m�Z̛ÇͤQw�lP�"O�P��͘�dP���D�!42i�2"OhњWJ�]FR��$&\E��-A�"O����� 4XyK��BY߶�r�"O� [`A^�p"B��]�����(D�t�&�!e�|��S˂�E��fB�	�S-�	�b�A���0W�M�liTB�	�:l-�V
�.�z �S���$BB�ɽd�����%BoZ<�#�C��C�ɠu�0L�f��)Г�Y�*C��/�HK�e����m	��4�TB�Ɇn�.|��
.Z����+��oq|C�ɭ>����;U����N� JC��30qD(T!Ƚ=��=Äϡyt��D�Pf2-���F�|�cS��g!��?S�l(S�A��0�.l�-�Ic!�A5֘i�j���RG'��U�!��u�者K�]��%���j�!� �fQ�%��
z��C�dU 2�!�Ǆ.^��µO��|2���a�1M=!��\�ld4t+�ᖿu�Y��Ũ�!�B�8�@0s鏳MO��a�A�Q!�$�1/'V)��m�587։�����O!�ĆI�� *ݮ2��tU���7H�B��0l�tG]�y�x��E,�C�I+/�pht�!����į/dC�I/(VJd3��e�H���ܒB�I�Xd�Q�`��!I#-X?'s�B�I� ��p �*��� �$�<	evB��6AHb�c$b]+I���P�^�?�2C�	&q�Ld`��X)B)2Y9��14:NC�I�l�.��QOW G"*2%H���C�	*k�$u㶦�?	�h���ϰC�I�};�� r�Дe3H)s"͌"KܔC�I�A��ڤNF�xE<e<�B�I�J���b�+V!^�ǧ	H}TC�ɔ�t����^�F�"9Y	ta(C�Il+5#�$ӹ@yP���gZ��B�'&���� ��},4!@�[/'�B�	 Bq�E��y�����l�r�C䉅%��!����%��z��8C��;o|�=���Y7Д���C�w��<�a$O��0�a��3FF�z0b�E�`Y�p"O=#2'õ;�& �¡�$.,�(�ȑ/!�$�6@�`���15艙��U�O{�z�CQ�$�Ò��V�)����S�"��ȓ� Fo��TW�%�G��<�=y0�*�S�rl"��5��/pv,�S���E?�B��j ���1�-C�&a����d"=��'d��Xg�M&YF�]��l�8�"O��A Ʒ�t���n��f´�
ԹiS��	�|�(��w� W�r���H��A ��$3�)� ^�ل�ޱ~��J=h09b6"ONa"�-P��LQrj�;DL,-���?�S�9L��2�A��$!y��+3�*B�ɧz:��sK��%#g. [�B䉔<.��:���cQ]�eS-LN�B�	�{VT��bgņ�DY�V�MtXB�IA�8�S�5$�nщh��clB䉔V4���"I).�$��Ҥ�S�fB�	]���W'�</D��6��5<B�ɇ.(�@�H@��a]rg"B��4')�K�	7��(�q�M�B�ɨH:M�`����P�$#L �B�w�^��R�N8k��}�/�>!pB�7}����mJG
�١���g/JB���J�따<��C6-V�g$B�eC.�r����٣�&��s�B�ɩ`�R����qǞu����r
B䉮CJ�xt5�R��U�'E�B��$\�(tՄ�H������5�B��'�d��ۄ�D�d���h0NC��bNѡT�]�8:��̏�p\C�	�Y�EU!.Z	��۪\�C�I�P��ሗ�C�;�,�#EJ4�C��'16� 3F��1{(ً��X��C�ɼ}hd�8�M�yC9�����C�6D�}2�L�`�<\�a#�t�LC�Ɂu�����KȠr�2�S���*E�NB䉗 xT,ٲ	I9�,hp��=3�&B�I*\�Ⱥ�c�&���� '�bC�I�b��a9$��&��!�M�NfbC�	�2�L4	�O�D���jq�W�T�\C�I��.T��.�(�z�gԧSuC�	<�|�v��$T���u�O�r��B�	�z�5j�G�L�b��2���B�I�`���z� � 3X�@���zk�B�Sr���g̠T�.4)u�Βy�B�	K%�:V��Mw��b�-@�>̀B�;^ĵ�KK��}�" /Y�NB�	�t��Á@P��v-p�G���B�	%4�l��X�x� ���TTrC�	x���04.îP�}(�
!�RC�#20���A�?�����H�
L^C�	�4TXp�� �.M>��١Cƨ&xFC�1GH��!!�G�h��'΅�C�
�.�2��X8d�0�1G}N�B䉴?����΀:�Ԓtn��?}B�	^�^�k�/R�j]z���<�C�ɔ^4�e�(c/�)�p��{��B��
|�"�:��H�P}j� Ī�*T�vB�Ʉ����Ъ�?�^��(��r�pB�I�M�=��H;S+�������(B�R}.T����k��e�uC<� B��+v���9�؏~����`�Vd�C�	 (�D�Q�d�"6�F1���JT�B䉘U<�<���ו|&us��J*�C䉪J��IaR���v���:�B0szC�ɐ#�T��NW�p�\9ǋ��C�B�*]�� !��
���p����2C�%�U`�e� E�f񋵤֨]s^C�I�t)�͛FCtI`y*�h�H��C�	,}
��@T暜n�`e���_Z�C�ɉP��T��"�
@�J-���=N��D��-j�D(�bL�g>��eO��!�?Z��a�`dA,
5\d���'P�!�� >��MQ�_`����ӑ.=�K�"OP�Ӧo����w�l>���"Oj�X�ٴZ  �B���V&jq�"O�		Gk�)�-B��"\�t"O!T
�����ϔ3�q��"O,Ѡg�  �   	   Ĵ���	��Z��vID�:B���C���NNT�D��e�2Tx��ƕ	#��4"�V���Yq�m"J�ν*W�X�}�]3R��)�J��&H��V����A��M[�%S��뎁�w��;Z�V���'��Y�����?�C$M;���G���j��3�G~y�d�3�8�`E�/}�ㅄ8a�*���1`�<���ڇ.'(t�I�f���'ԀB�fh-|��h�<���]>rd�d��o}�R�T}�X��m\�* ���'�L�J���T۸E�'_JEXǎ�1/����O�8e�,�z���k &F=�8��&@�*g0��W�>S#�"F��)L<�'-�>x���I�O'�Ea���aR��PU�� �� �'Ċ$��ͅ�S�'���� �.u��O�$�9গ�D�����͚�
,J�g_6KN�K��>)�I�cX�&�,Z��W�cF��۶���qA�韃�b}A��'�H���r��|��'f����'�2B�k�1�6M�S�/`��-2��O�D���7��'U:�S1�����Sy&�p�\Z\#F��7�<P+	;C���O�m���F�O��'��xk>�n���LP.�7F&؉��)�(!z�:Di���@&:R�g��e�اLv�I_ ���u�Z7 ��t�AM
>-��ѓ�[�DѨ�Di��W"<02(O��B�P4��&P �Tu���z��U9'�I���)��� �
C�	3T�%���i�,��f�'�\�C�O1h`*�w"�<�!
17:n�<��9���&�J����ޛ���S�[�b��dR�O�LRN<y�O� �bn���:�Ё�&6r��Y�ϡ-挺����	��aN�:J���a�?��$Ȝ5m������'���"!"+7�zqc@�,
\�,O草�ȊM��'O���΋��JL�-��c��b#�
9�8y:!*��E�B�%�PyDbW�A�rb�x�1]e��B�aGj��
WY�z�L��"Oj���  �?}��)�+@x:#㢐��y�b�,B d  ��K%D�@�th�\N(�dI�����1'1D��"5�\�[K8���*�2Pw����D/D��R��E�~AɁ�V�zh)�-D�$�P��	F�v�8��(�bs�*D��b +?�u�mN�*�U)�C(D�8�"6p ��!@��R�\�E3D����$ /(��P��@(,��,0D���1�V\��:��s�>x��a-D�p�6/��6ΤQ��K&�(���l)D�X   �  K  �"  -  �5  T@  �J  }T  �Z  a  Tg  �o  �x  $  v�  ��  ��  B�  ��  ��  1�   `� u�	����Zv)C�'ll\�0Kz+��D��`���b�ƦY�y���yfY$E+��[�J��F��c�&P9H`Ha���͜`���3�+ԧk~��pE�� 2�U�%H���Lr&�I�t@(��,E�WBb X�	�`^�ً�)�+�򍃃M�u{�����I����;����'�?	��͘PԨơ�wO�p���ڠP1jxj#BO�ZӨ3T��LYI��6M�4J�$�O��d�O����:�ڀp��0`���x�-��9N���O�o�epBH�'s�CX�R`�d�'����e��4�'��$Hi��韒A���'r�'���'��/�=�uw�$}Jmcq��S�6Hi0j�WL�P�ZA�Ҥ%R�4@����ɁO�f�<��m��(d���E�M�d-���7,0��A�OF�	w�M�p-xe�.BvQ`�'M2]`+Z\������pI�����A��&�'�2�'��O!�[>��;Tΐh��P7R������km(̓�M�жi,�7���a�I�MӶ��g񛦆�ZP�˓&ܪ,�=��F�Z�>��b��E�#=!�N���Oj���SH�cC��qp
͙~��:%(U0�>���h�#"���ߴ2��Flӆ����|�"��))���.��_n�Q7	�H�x!�\��N�!<�<�`D��
d�U�i�4�����$L����e��nZ&6�\�i�R�HÐ V5�a�'�;̵!�d���M��i9�6�܈$�ꔲ�@ �)H�z#.F	~8�bĄ,0�n�s �$V��)�+�/F��J#�nLn���MKдir`����ݷn�$�A�k\��<0b��*��1jDdO��5�D�I#8��6톹�(�a"B�0b��9!�ǝ�|Xb��>�I	J�D�r���=^q�-��L%�̢d��z�	ʟ��I�?	��e���c�A�L��L��}��a�dޅP� (qi�d���IByR�'�2=�H�d��?,p�蛆�T�,�>e��NIN��%	4�I4�W�C�4�E~B/�4~�x"�)D9g�����@�4;�$���
*����I�R������bۨ� �)VܓoVV�I��Mc�_��8�M� ~� Xrc*	t<Պ�O����O��O2�d�O����O��>��L�HL�iN�%b��E�UK<��CզE���2�ДAS��<Y�ł 
I�M���BF�ǟ`�"6�O�˓����?!�F9)�bI�cc�m�4	��?��1t"IuAЭ�����
 ���P��3�/�Ѝ3� ;H�0jf��A��'��@׎L���ǐ&C��)�/q���FH�>���C���Dj3�V�X��J���eҝ�	/�M��S�|�R�H��H�.�,Ko�p�D�ןl�?q���I1cEƍ�qg�Z(B�"���).�ң=	�'t��o�P��ꦙϓ>V�P{r�i�H�"KB!�	�H�'?���5�'�2�'�R� �&FW�ZihA!i��H���+]t�;R��Dp,�s�hG��,�O�Tz�	�'��`鴧U iq�4��*O:g�p�;q�y���G�V���
u�]���/وyH��c�B���֨�ɗ�8 �S2H���M��\��@�O��I#&���R��W(٬ ��m��I֟|�INy��'J��K���c�1SR-����';z7m��1%���?�'�xX����W#�*�,lz��0�ES��?����|�O�v��a�A�.)2r��:<�
ȡ�j�g��3�H����,�a���~Ǹ#?��)��#z���j ��UU�L�)�2x�r!�7���#���up
,��O��eD������'$�t�E�J��"gI���}�#,���?)��i�h"=���"�&xp�Y��jAYԂY���6G��'���'%�\iVD��eX�j�NڮL֬�I>�W�i�6-�<�C�H&v���ğ(�&�Xzi���õ����l�ߟ����a&l���|�	\b��G�L�*q�I�j�XCRq� ��A�j�:ug�8t�����:f��8[fĘ��"!˗��o��l��HT.R�J��'#����@%̑�9��)#��
'yA�����Ӽ ��f��1oZ��t��J�I��DF�xdj<��i�cyB�'
2�'�a����)>�:ɠ`G���h]y$J0��?� �i��+���o��d�p�*Nbi�g�8�n�>!*��?�?����	+t�t�$�6Gy�d��)Ӻ%m��&	���O�"��O2T9S��6qY��\!��V>ơ� z��ՠ�jS.#��d1b&[~r�X>l*�Q��! �x�"G͐&#۲�k��݂,6$ ��O!��6�1W%�h�djI�O�ĐC�OH����'�@7m\_�b�'I�����E���\R0��*H'����Y�ʘ'0v!HQ+Ë���!%瘱/��0�(O���E�O*�����i�N�Ė�U�I�-�<a�G�W"�1R���A2t��ڴ�?�(O��SV�䟆�$�O��D�<q��؞|d�� �(�vUxԡ/�*;�@m�U�� � �)��E���(���݄�ē\z2iR�!����%�dR�i�!W=F �[b���6WЈ�
e��,��� ݔ"�.G����K�;X�8�$� 5@6m����S(@���'���'��pr�^X�Q���0Ț��'{"�'�b�'��W��´J��T�CW��'lM̸�'�(6M��i��#�M��������)�� �{'��  y�ͱa���Œ�ʁ�������\��uy�R>�ϧq;��IA�Ѣ3�lp7̇�#�:@��ƽ��B&C��H�"�C�v�����s���K�K�8
�h�*�$�
Y��W�i�^�g-ip�Z9����d�Y��;����K�-+�4�i� _(�栚��џ|�ڴ0 ���Ex��Q�vx��@h�c�*\�?����'�t��#��L<�p�3�
03^��ZH>Yd�i��6��<��jCI��I͟T�5(�0Rs��T�˝>$�D�G�E�H��Ty���	矰��0s�I���S��ܴ�y� �,BD_3�.�zV͋�4:�����'�f< �G:S~�x�r��-}����˽��YjAn\���B�cv"?&(���8k۴r����' ���ǡS^S��Ȳaԥ0 �#S����ɟt�	D>EJ��	�� 1�!k�LI��;U�7�Ov�m�N�V�pGS"���k��J���ݴ��խ%i6l�d�'��t�O����#��q��)���jQ¬��X�R�'���xr�8!�* �	��3�z�
��	 ���cɟ���Lн�e��OV+3=�i�V�<?Yb!R�F	�S��� /Rt�/J����SȥsE��?EhEЊ+�T�3�A�FS�U�n9?�W(���شV�>I�'e����5�]g�d0�dD��TG{��O/!7�F�3��@��A�I��T��$�O6�n�5�M�N>!��٤B��K�m��h���1k��h����'��ɠU�4�S���I�H�'�e���!a�p7�MN�|�I�M\>Š�M�Mİ��d�ʘc����?��AD�$R�ɉv�8�j��׎D���r6���q���EN��&�y���`b�)�j�L��	�O�^�sAѱ�yg��1�G(śX:0�m˓	���'�<�⁙۟��J�L>�����pxq%&7�9��؆��'Xў�O�>D��#]Z�	�"J	+-�����?�U�i��7�+�4�����<�ѩƁ[4�����l�s�W�L����i���'bP�b>Y���
Q���L�mǰ�:ŏ��.�Y� �	$Y?Lี
O9a�" �a���=?B�<Y�J>����O�BD0�^Ff�	�N�Q��\�-��1�
=H� ��%��8��.F���&��)Ѭ� Z�����G���`��	���شs����Gxr��M�Fyң��.��@.���=��y�l�	l#�I��/V܄B�*�<��P����'��	�q��B�4�?���:���Ze2�%��Q�Q=Д����?����?q��?QE!��#�����\�<��w����fX�H�^I	�Í�:���8Ó����� 2*	h�%�34����pM�E�6�H�G(rR���G�z�8Z���O��oڗ���I
S7Le���Ӫ@�>=����E�|��D&�a(�zQH�	D����`�57� �Imx�,�޴����g�G�����5�ypG�i��eb�v�k4KĦ���Fy2]>�L�-�F�40�0�c��@�psfa��ڟ�]�t
C�-#L�������E*wa-Z(C��A�u. �]���b�������h��PHB�N���yt�<��)��̓c_
�Z�M�� ex�!55���`�!��t����,����O<m���H��Sg�Ab�I��R ƌ6$�:��F{J?�REӼ#7�����\��[T�&ړ�?)c�ip�7�%�DS����pD]A�>��DH�WF�l���ĕ'�D�+3�O��'�Y���� >d���$ +G����ϛ�,{\ԁ���<("�h��[<S� %�|���W�g���INӰP��v
��C-��p�d\�U��H�1�C�D��  w�� t�T��O�Ε�Q��yר�(2�Kf�Y�6��lAa�^���F�<�Gg������H�L>�c�g�@ʓ�\EH %X`i1�y"""5�ũ�L��l*q�)���?!�1�������'&��A��.$�����7�f=PU�'>7-�O��d�O����I�O���N�YE깘c�оX� %�6�;��˥d��'�}�O�]�,"�M�%k$Q�H�EEܰ���"QH�A��)yf�B�'\`kы�<	��T�׋R��XcDK,!�H2C��D�	� �l9����:���J�V
{�������O<�c�j��u7��S�ZY����fܫO�����d5p*�d�O���/�$�<�}�5���ta�!��9y�PņEy��'�7��O:�N���ָi;R1O<P�.�l�b�lL�2�l�g�'�������|��Ė�<����%6�Q���W'
4�a��+{� ����Xp.���f�2>�<	qeܰL��#SDͦ�pE�;�ΐ땣T�f͖C�]İ�cW*A�dP��h��9	7�'U���}4��/�<�F�$�%��Mc�����y�I���j��(p�se8q=зƶ<	,O �=�'^\��eH^|�9!��
z|��#�_6��<		y)���'�I_���'����������Uf?��=q#�'��l��h&а��7�)�ظ>�� �}�gą�Rv���q�F�)v:\B6�Ž����*>
�ɇ.�L���QH �&(��@r�$|!�O��s�N��~�
��lD�`��@�O�X�')6�g�O���Fc)c ���y�n���#.��y��� \�9�"C�bA8�j�	Mz��?I��i�7�3�SC�"�ig�C&����iI6�l����9%E�l�u��⟐�	ޟ4�;{4���cX!cŦ�1�̀�u�0-�D��&R�UKu��\��8�i̧��>�|m�&%��` ��������N=V<�x�S�H
fx����όf�'��/r����/W�Ж��PDM(�� �	N~����?���?Q���ktJ|������ ��Ө\q!��˒i50�9�d�Q��Œ2p��_����S��'��\��&�[$:DiB"lt|q�u��T�E�'xb�'��ݕ�	ڟXͧG;<��b�>L�T����w���V���x-�U�'�%[��YtOּ]��<�$d1�d-��� �5@Ĭ��i�bЉq�"\{�Ը��c��(�4��e6�kր�+�^�A��T���J���.�6�� ���̱��'Vj6YF�'�����(¹l�8h@C3LT�(���:D�HH5�9&��8�vO�8*�	�c%���ަQ�I^y�ύ�U@��'�?A�(F�ai
�J'c_+\r
��w,B��?���>�,�J���?�O9����6J쑴�O�Wﶠ�����R��I�_<�tq���L��q��Hr�'�R�ZgDhZ�l�@�e����eO^�]�񥝆#��H���=9* A�W^�'vx�����V`�<91gǤ�Phs��&��`)���\��q�pZA�1	6H�
��L\=�X�#0�O���I7mQ���`�vyd�JÃ�:����$,U6\mZܟ��Iu�$��Ha��
8-��0梋�s/�h��@i���'>ěd$�ahQ�dO#=&|9�S>9�O��@���=j1~0����7g�$��O�@���Լm�y���
Q䪌�	�ޠ�����،�Z�(L���	��~��'�>	�,��e��.DS����@fI��5��N(�X`�@ n	��F�%�G�n&ڧj\=X��ߊV��A�POԠ,�S�4�?A��?�B���#�����?���?i�w��pR�X A�N��D���O�KՎE��P�x�*��Lt(���8�Ot�'�= ���2Y�@Rd�G9#/��¦(T�;^�|B��D<EʦDz$�ۘO��'�X���+�c��h�"N܉
�n�Q����\x?����hO���P��:	��a�m!f7&l�&)-D���p!�x�A@�!�\5���,�<���i>��IkyR�R�B��A`�0yF	a�OE�0�.W�-��'�R�'���ϟ(�I�|B&E]��>`*�p<��'�۷4HBta��
3��u���δLV�2`�	�lӞ�9fn����7ᖄ5W���F��g�����eU&Fz��Y3ⓥZ���Ye�&�7���@'�֟;Q�Xx/ޮB�������̟����g\&���K���bA�"m�ba��a�ԁ1� �f�u��C��'��R۴��
� `2�V?A��ei�+FM2y�]��G�1{J��I��$q@�៘�	�|����0zࡋ���
0{� ���SĨ�	��Mr�JI�.������qyB��D����|1^�i��%�Fu��+1�"KP�A:��E{I>�?�����ē7��3eF�#�*��Bf�
�'�a|B
�.Q�L��d F���R�C��?��'8�l��@�\��0Ѳ�Ȼ8��������du���$#�i�|J�C:� ǋ�z^����7 ~Y���?)� ��{����b��7/�`��F0 b?�hd <D��%�5oT�Y�=?	��\�h�W�tlVM蒊ɝR��"4�t-A�*>H�׀�58 ��ԝ�`����O:�d)ڧ�y"
I�V}b�)����`N��yr��*08%Aی
儜�֏���OV�G��a�)S�0�P1���#����?9�����ݼ2N����O��D�O�˓Sb�`�k�M"<yB�HB9Es��{C@�,�~��v䟼 �4D��7��O��O�B5F
�"0He� ��D�����(�#w| *�'><K�	�WMV�_�1�0�%��I�/��[0Tb1�å8q��3���O^�Hr�D�����D{�#LF���b� P)6���a!P�t�!��ĩ�,0ؒ��:b�ĥ�G�� ��1�HO��O�ʓ(y~�R �we�,��"�<=���߻Ep��?���?	��G����O��m>����ܺ��F��x�����+ ���BȌ�A,���`��Ű<��ރD#̌���^����柸Q�r�3��3|�R���X�'ayΉ�u6�=�"2?P``���ch@����?Q���)�9T8���"yZ\ xIw%\��ȓIr��F$7�����S�\���'�a�4�?�/O�m���XS���';>�ӑ =4���⠉�M/��1�'i������'��	�&����QNҚk^8L1	�''HP���6jq����'�>w����
�U��ҍ���6g`�1ᕶQ���o�¥@���{����e��`�Q�1��eʌ�d��L���'<�I!���e��Yl�425���g�֒O����I�}r�"DB�(F�i��Y����D���� �H<X�D��m�5�!k�O�������?�����5����	@�
H����������W�Wd����O�rmT�?��]y��Tv�Ի��Od��?x`j��Q ��xe�W�D�D��fD5?�L�55�@5�����3c�k3J
��5��:���O[��Cc[9e8�h��.1H�?q���I�XF�t:O������qv���&��=ۆ"O�Ȩ�X;q.�,˲���P��aȃ����h�ܰh1��o�ΐ`��� '�h!���'2R�'�"�
;�V���'���'�b9�d�0��ػc����=hB����Jg�Nr�ā	�a"��I!)�1�̓O��G�\�mm��RM�42J�g�5T�e�5`@����r�c��v1�D��EɅ�~
� :eش.��*t�g�J�1��'��	�>*t�$�OУ=YG��CI����/�r�a�˙�y�*��e��D�~�Z�"tn����M�����'��	�2����D�ʼn��QN��M4I��:h���I���Iן�������	��0�C&��<��0�f�3[�ܢD��j\����\�+�+��2a� �B�ƸwF�չ3.��"׎990�=�4b4�'@���SX�v��gǖ	B��MJ3��?��i��"=���޶Pu`G���t_B���Hc�O��3�m[p��Q���
I�+��|Eh��8oZYyB�8[�6��O����:Mʰ�vM	�-[���!*�0=8V���O� �a��O��d�O����+ 2>Z �b���a��P#G<,U;�	i�0kvn�M�<32^ꪠq eԪcF�,3"�Q:$��\� �)Q�xX�!�NX:��DҤ ��c���'�i��]�D�n�F������'���1��I� iQBb��=)������O���ĄߦA�c%�u^L�����"�IRB��2�M��[��c+e�6M�O��d�O>��Ң\1����O0C�A��Y5.B#� {$<��O���^��3W�Z���Q��c��Sb����5�:8!�BD4�zsL�&��O% ���� �,k�F��$RZ�O��<Ռ�4���Ksk�6g�����O����'����<	�D�mv��Z �����j���|�<a���*~�x�Rɑ]��X���{�'�T�}Bvn��J[taJs�V3[�~�zCO⟬�I����I�.E�,J�����D�I�����[�=0�v�[S��5����O�vA�Ur l�$�?�Ηa�x�|�<96�0[�}�D_=F��U��a�PJ\q�Z��?��/ip���|�<�&T<%a>�2�د(��nȟ�'&V����?���$�>60��9������gF�~x�C�ɷXJQ��K5.>�0��­>�H˓Q*����ߟ0�'a)�����~�� M�<h�F /�,隦������'��'X��,���|�V�Oޠcu�؎ e|1ڱ �4������!ewy���8.��3��I� #ƽ�rB�>��1�b�hF��Q��J0*t�pr�(�5A�%�&���D��q�&�T5ĸ��\�2Gdx�g� ^��dK��#�����&��T(�y�LF3[Τ�ȓ$ZJqH``O'm��-�#�2Q��)$��{ܴ��8<����X?���nJ��cFD-M�|8c%N�+=���I͟��o���	�|zQ �7�&�R&L��)QP����D8�* O�bEt��S�NWbi�ቕI�J�X�J?�ف�����R1fM�8�~5�� 0�R"b�.O�ɹ��'2����z7�O4Z{LP�M�8.@:L e�9���O>����$Mi�pS�CE�Q��Ӂׂ;����O2x���YjL���)%R����'��ɪi�@ٴ�?����	M":����ը_2%�����+m�x�t螆I���$�O(��aD}�2�uM��-6.���|�ϟBPs�8���BQ� �*m8�����ƅ`����<�DF��(��4�6��!�]m��q{%����޻���'��>��r�J���ӱ�0���)��~�J݄�
Llq��C "���S';'�2�D2.8ڧ�����-�=���a�OC�+���bٴ�?�*O�i@�������O ��<�#� K��{d[�b�x)b�BlT�8�'gG� &�o��	􄹍��y§�.Z�6@ͣ"�j٘�E�q�44�W��-���\�30j�v��C�Kq\,��nY����`g!�,$W2�� �.�O���.ړ8�Дk�m�Xx��@�O�jT�	�'gB���5����H1	�T��(O�1DzʟʓS�hm�b��
���B½u)t�y�ܻlǛ��'R��'>�)�A�:��a�@� \!0��|TX��QiI�x}6�0g��9� x�d�!��ODyH�e�>Р��s�_9c� ZAU(W
�]B��փ�-2G���op��?F	�/s| =c����!�I@�Q����������c�����Y��T�6�
a�!�ԫ7�� :�"O��[�g�!
�H���1Z@�pҞ|$�>�/ON1JV�)qs���a�^9\Tb|ڄ�ǋEp��<	���?���s�����'�v����\[��0�%�-�h�24 =� ���@�"4џp�R��W�ҐUn�'�L	I�<V<4@	�KM�H0�	Íb4:xFrE�/�?����59E���2�[k��Y�u�}�'�a|�-ņ$q��Hp�ndݺ�,���?�4�'�4���)8�(uC`�WEma����$C~�S��P>q��~(�!#�W�Dr���ɨ<Ӓ��	��T���Yg�0�0/P�N`�� a���O���aBŅ`<`�ۀ� I�A!�O�|�$�P<���j�wT��
*�S�4�Zm���ߢu$h��bP�ww@�F.���I�HD�42O� �=���b����R�K$�b�"O�|�èϼW���3$�
�h.P�I���h��r�OL�0F�H���ax$�':9���4�Q���BB��D�>����'�ڵq��<D�D�ՁʅC�h�BeY�?��=��&D�X;��϶1��cp��4>\�;�%D�;Rϊ�oҲ��B  O�m�3�%D�,� &A�})��Z1�?b��9��"D��2�ُi��<	R�C����6/�<)˗v8��!6f_�7=b�P�F�f؆�1��7D��vOW�C6yr��0_H��E4D��qD��3�4�u�B�'/}�S'&D� s �Z*TF"$YSEݜkI��Q�"D�p�WC� ?,d��ϼlQtk�n=�O扐q�OT]0f�A
^��偒$���A�"O�4���=WQ�ը��)��� "O�رu@�&L�)��O�}���`"O<��2�)%��5W�`�0��A"O*��g��)J�=f:dxa"O�A�5C�<3Ķ�aMFF1^�I��Io��~*4ʝ-�k�䊮	8�`���d�<ɡ��)b� ���`U~��""�W�<�!n��Q�={��,A�n� �mLV�<a��Ǝ����!��$|��#��JH�<����Wg�8�r�\�Y8z #�m�<�,��]q���PO[/5"��!���`#� �S�O'dy��
&8}�l��%ֆ?f2�2�"O�ciAtT 	 �k�����&4D�TXQ��2:�rt"H�?�
e�!�3D�h�5���b΂E��)U��f3D�x�RS2%��I�o��)�#44� RwGM��
@j��: ��%���|t����-���kp&1i��L2�'�6b&`�;j����O�wĝ�j�@�y�O�%e�$Ȁ� h����	q��'�b�W�P�%FGC�
d��c� Q��)��i��'�̾\��Qi@!���(v �"Ժض$����i�UA���%\�'�"��$�!O�du�E�=3Q�(�3#�OF��/�S,Ր���֥Fj\�
Ƌ�4~P��0?��A��0���2���0,.i��QLx���/O �JP�A�HP(u���.��0R�`J�k��L���� �O��Y���'1RB�]UN�(�$U��.(����)�R��x"�=ځ)��o��X�!��d6����O�������x�%'C�y00a��'Yr���lr4��^�x۸)q�ƚ	'�.��}� I`G<Rǧ_�v���<9Fă���}~J~:�Ob�����1tj�"j�>t���A""O�41F�وz��#iŜ"�l�{c�I��ȟ�5@�+$۲4вb��xO6�����Ol���O�����E�Ú���Or���O&���O �W��{���鰋�<�� 	uB[�J\}��O�9ϊ��pM��@o~�'��'>0��5�N+K��Y�F�=
�m$�|+�M�X~~��2��1��I�&Q�.x�J���Fʞ���� E�R�2��3�;?�1������{�'��T?�jQתW�T�n�b$�ط.�!�$W4k�T)�c��#*�Ęj����*��|:���dH8���9�#��b�I���'XS֤ �f�]1&�d�O��d�O��	�O��$w>�Y����D�)zb���HMS�)I��{g��7��E��M-�UD�
� c�x3��X{̤<B���=���:�C^[�Η�V>̙���e˔�2�)�)��X�I�F9zIЀU�x��B�Џf=4���X�'`�t��!Zxu�U �L&D`�8D�P���58H$X��#4F�R1(�<�f�i��[�|81��4��i�O�S (~�y�׫^1=�x�x�<�F���&P�����O��dV�

�s	�(-��]�a�%�����XrP�bJ�(D�$�e�R�T#>ᦄ�=8S��TMltR�X�t%Tt��"�.�.�ҁ��;���pҾNM~�<����Οl�	w�'7��bA
[�V ���[6"���'�a~b�;r��2�H�P� i	-��>��V���bB$L0��!���'g�ӑ�>?Q&O�ɟ$����X�O�G����ݜ�L��D�,
�A��M�2䐌���)$�l�g����9(�(D#'ݨU1��"b>��eI�b���_�߲Ȋ3�y�hxb� �$��p�ǴzD7�\�  � ��8�ӥ8ٔ�He\�č��G3϶�%P���O�S��O~
� ֈ�g.xI�4+ԭW*C ��j�"O4����.&z!�ɣ3>B퉋�ȟb��c���X1��c���B��ׁ�O6�$�OT9�7�B�Q��$�O��D�OR���OF�����\dSpa�1z>@2���	M�@����2cdEa��=c�����'��"��[�R���:Ť�E�-�1I:U����)�+UJ��I2�ې��I_�n�FL�H�0�B�>SUJu�&� v�`SAM,?��M�����T�'P�M3_�0���g]�$��Ց���#N@!�	Y��r���N�UJЏ��#8b�6��|2���D^����a  <�)��2I3��+�B�1����O����OV�I�OL�Dr>�R@JȤ(8I����-�J�c�S�7Y� r� 	��ո�o�!0��1E�-�7�@jD�aҦ MW�r���ʏ&�Р3F\<Zm��6/G�,�hDEy��F��?1"��	��  �
�f��:��	�?��$�$z✂ωw؈�*!�S�	�ȓ?X�`10���x2M�db@�\X�!�'��7M�Oz����&_?u�I�|"���	
~��sLȬp&h��sʅ����fE�Ο��	ğ(��fσ\8$U�pN7@J���p�K�����ټ{08U���ߒg�N��#k�'���҄�/_��r�J��40t��ƭS�K�"T�#/rV�p��C&u7��F�N�'��� ��?��T��+]n�� @��F�ܠ�	,��$#�Of�XaK�=�E `��>-�(%�A�'@�ʓb��m HȚr����,ʪ'Pڄ�'i�'�R�'S�W>��I�|� mՑ72�%�穙-iY:����EyB�@��'F�"=9rmѲ� Y#�Q�Y�$ɴ,����'��	iH<�7!�O0�'~�1�$a�)��p@�ݪ=��q�i�B��Z�<u���'���'y�d4F6$�2��M�g�$�H���?D,a ��y��$��|��h�#uƸ?7���5VA�?���GWK����*\������<�d��<�]w��'���'���,*F�	�oU�U��'�X&Fr��R�'���wDB4OB�П�^w�b� ��GgܳU�Ұ;�M�m�.�C�|s��I�fiù�?�_w���'��$�O#��``�<,�`L�	����9��O��˒�'���'20Ojh��֟�^w8��]�<<�$9%�/m��9�$ː��6�g���On�d��s!��� ���?� ���`f�1I���[������;�Ńq�)���O�d�кS��yB�C�_��T�i�����FF>LU��x��r�Ƒ�s,�+Lj`6�
џhRB��O$��z���O�R�'9`8E��5XnT�J%	ЌKR�}[��c�$�¶�m��Q	J���Sڴ�R�H���:�?��*5d�����Rt��=�@,����֩��=[�>O�7M��?�oZ���.O���%N������*J����JX�H��C�	!gq�};��1m��t#� U5@~�6��O��$�O�$�T���'�2P>7��K� �;ңʺ H����O���'z2�'�r�'��'N��'�)�-�.eҐ'̸{/�|hC)B�\��F�|�'��O~�O�ݢ G��脝��eB�y�8��4���?9��x"�ۤpD�1۲F��sJ��q�&���$9�OX�"b�:k�0�( �T;��֝x�'��m�%�K�YG:pH����h�����~R��8Y�J50V��n�N�*��͸�y�,\�4��%�T�n��6T�y/�}O~� �(ݬ1z��ڤ���y2�1:kB4��T&��)�SN��y�<z�69H@��Ж`�����yBJC},#�ڥ���b����O$�B�ۘ���u�(sf.(v��k���;�Ѱ4��v��������yb�A'C�A�����"�`�p���6��'A�i��-��j�E�1����c��%��1�h%T�h9`i�#�����b���� ���	�~��p��5g`4QK��36<b�x�o� 6[ �E��^�A�����$G�!IC�3K�}�'�|�(3��>��)���٢c�2��dk�'���""fջTe&Ur^��ش-Q������"%j�X��+H+\��]ٲ�'��A�.�r�T>�KMR)��oS)A�XbL�1-��%��[�4�S�'l����ŋ�&�vݥK�n�'�P:�-�O"�&�b?�+���_vmciJ�����A=D�|#2g&T+�mbA .�xQI�;O�PGy��Ҝ4���M�X,�1����&-:�mZ��I�XY�kI*[5 !�	����џ��Q�F.�hR�-I��`ԍ��2�A�<Y&�UX��SV#�.�>�i��R�1�T�Ua7�	�"W���K4��@K<[�������S������8�	�)�3�d�)@j����n�0l�� n�!򤒋'M���D�ZJ��x��7��gk����W�I8�@�3����Y�G���k+n��)�=)�u@���?���?q#��F�$�O$�5'b e�b�\'7��R�MH�N-R����<�x�	� �	��'�D�1Ɠ��� ���I<��-	��@��C/rN�	�cV�-���	��p?�ҘR�.ܚ�+F�-�ި �S�<�mӕDH�m��@ɛ7	�"	�W�dv�6�|r�G0��6-�O�7-
�Br�A���n5h�j���NB��	ߟ Ð&�����|zro럘&�� VA������&�żKݸ� i',OұB�$Q�;B�kaD��aD���D�1g'ay�B��?��>9Ƌ�/�&A���޾c�n��u�SN�<����N��I<NS����f N(<	0�Q	|���R�O=4���`VI�+B�xI>�����?)��?q)�� 냂d���MM�=���r�c�?ߞ�Y� �ڟd�I�tQ�l�	]�S�,O�%�Տ��:�~h��A�cєh���xB����O��R���� mơyD �*��u��x� 0�?�4�|��$��2�����ɬP�� �M�	�yr�O���c���7Ƹ��5 Ŭ�p<�@�%B%�Ph�3�DC�"�60�F!�a�i�'���n�!�֏�ǟ��	꟬��w�TX@�/��p��j�#M�Vb���T�:,O8h��7vߠ�vnQV��З�d]W@ay���RJ�E� 6kt�a2*Z�m�P�%��A2��Oq��'��Ѩ7�����׈��0.���'�ry�V��\݀<�gP�&9�L�����4�O��c��G�_�l(`��J�m�b�I�6�d��1@�Ɵ������?E����|�'�tYXV/�=*qbx*�ށ^��k�\<a�)X{��բb��"{�A@�P�''ZŅ��x��0Jg:q�.av,Ȉ@&����⟀��0pr��h�+4�����c��h�4�ȓ`+ęPe�۫-��,�G�;_စ�=qT�i��',�¦�n���DbӖ����	_w>[���	_{����a����?gDf��Iߟ�ϧ|�mrva�m8ʓ}`:x�-F�ɒ�#��	�L���W}Z%�R��#z�q�	�=�0%)df$D̭K!��iOv�	��?O.1" �'4��'�N=�5�<O����J*Y�$���'>���wݦ7�m���'ޘ��'�4��`�/u��ѣ��W�<T)���!�'���B��o����O�ʧ� 91�4"�T`��U�w��u�rƄ���#�'�BN�LH�� 2���s�M�O�SC�t����pyЇ�S@,s�k���ē�X�	�Z9��D�Ԇ^�i�0�q�����ӗg0y�]g{�#G�Y��O��1&�'�.�O��.t�#�O�4�=b���T$�""OR��%T�A��8Q0��D�L����'���<���B"*��p��Ax/�sWGF>{�(��?A���?��� �?1���?i��ߵٱ���GAvA"�Cô�N�J��O /�\PV�[�BX���O3� ��)�
�i���DB�U1�x"#��l�xb���Ay��a$䊚Ua�R���4*� ��NlE,t�)��1W��ż��L�!bN��ǩ����1�C�*e�6M���a�ɺAhL��&7I�����$w���acK�d$�񛠈	 K�P��i�(��D!�?��c;�d�m��-yf@����pe�$!2�d�OL�m��L�'B�O��X�,�A��U�����	������ŲB�ŉ"�՜�?9��?	��>���OT�$�Of�$�Dj���ÁJq�~x`֦ڭ?��T��LU60<"(��ǞVxeÈ�C$M��w<{�%9�JT���e
�#�)r�f��g/����Z��7���@��t�DH4��Ƴ"��D`5��6r؂�(���< �*�'��7����Oy��'xBm�"]�LUR���;��0�`��b�<�d�OT�����P�S��HlZ�5fq(5�],I�Dt�M�J�zR+O&���Q�Izy�.�b 7�O�6mZ�B&� ��R4UF0jfF�%Ҧ5��ȟB����$�	��XrC8j��C��w��n��>��ɹ�vNLȩ�N!C�n��䗂(�T<��+ʉv�$m��g�#�H+R`F�l�(��P|�r�'�D���������۴���Z�}If��,nT� �S����I����?�:��;�<���R�4$�uۑeЧ�B�'��{r��tbb�qR�Ca.*-+ؘ.��5B7�v�6��?�%�ie��'g��x�ʽmZ�n681%�*N|HP���3t��t����?q�"H�'�p�JVK�Zq�f�'��Sz�Dn�?\�V�iR�56"e�ce���AG����ƠA���	ܪE\��j���-'	��Sb&����'J<1-O&�%>��'�� V�������=O��5��^�S=��?�����d�O��d�O���m�����9u�(�
�@��%2��!�:��Rr��4�N`�'�����iD���z��LQ�>�ʽ�g��C�F�'���'@5�B���+���'T"�[R눉oҹ#�
ۧd�����˙5�BX�� B�n��un�5$.d,XB��"}"+%�֘��♇NkF�K"�ګQ���Pc�@�8>�y�AH30v{���>� D�R����}X� ��2aE@Ɵ�'v�k��|����'�]�G��.��CS!�`!
�'�\�a$ݡu[� C�J�j�x�I��C��4���$�>q���^;JL�d��L�f��g$%7�`��f ܣi@"�'er�':H��ҟ��I�|��0V�A����u����qG�P:�b��՟.���S�-�-g�rF�ɺY�t "�@�?K^��n�,,=|���G;TG`B1@	�8��UÒ䚑(޼ B�/G��4
�#X=~o��I�Ũ+>V�:"���y�|Y 4 F��|�P5B�EYL���ȓO>��q���$�z��LɌ58�=�Q�i~�'6x��v����g�������`н}���CR�N���3c��	����' i�2�C�D�L��'Z�Ht�]�����II�:=��'P���qǗ��r�3'���KC,fwN`�`��{7�RD$��]l�{�!�_�'x2R��3��?U�=abQ�]�U�%k��J�PU��Fu��R����x<�BH[H�i��Ev�
����5Nn-h"�y��eAW,���v�QG�i
"�'��5Hdz-l�FZ
�Y�!��p�DS�.B^A9���?�7��*�?)�y*��I�;*J #q�\�=s��9Т˲t��Oh�0�)�4̮�a�o��e�������/˾O�-�'���O��lx�	OW:ms���6-�U0�"O\D� W>&� YȆ͉.5)>�A�'f�<!�X�R����Z1D�����  _�J7M�O(���O� �A��n�d�O.�D�Owdۖ#ԢEKR��;2�ҤS�gj�8ȗ�5��j��?�ŚrD;�J�D�2|.Dҵ.��0�8�7֯..Ԑ�䠊�f�b8s�	��o0�A�!�i6}����B=�DN��*W�B�v7��O��+
!ۭ�h��(�	�TH�!a�AT&��r��o2xC�	��ͯW�L� 4�P�~�Z�3"l8}��=��|�����dѯ��B�%n�a�«���19�*�OPd�I����	ן�ZwR��'L�	�1h����Yd%��pB��-G�,�᥊�l�B��d� (�J&lKΚ1I&(�0+�txb �2V�l�+U�S�Ųb��u�|{v�6J
�eKM׀^a`pP�ፌ&6�d�r��(Ʌ�8Fؽ�R׹+�ͳV-#D�@�v��y�P}j��Ř�A"�	3�M�K>���gᛆ�'�F*L�Z
�D]8c��{����$�O���$��O4�dd>��tB�OO�i�akI��d�ٖ�εF4̅	��'��y��}f�L�}p`�Wx�1[��.��<����� �N������1\t�1��Ԙ(�|ʁ>D�,��Ά=� �	h�t'v��<���f��:iDb1�F"Ȱ�b0���5�Ψ'���u�\�����O�˧i�v�1�4!��9c3oڥi hS�(�~t�r�'��gH.l������!�$�b2�W�!�h[�_9��/%�6ې%
�	[�} B�S�<=.O�j�üD��RWBYqKl��&��5?4:�;.������Q��2����ƠjxBZ��?��h�n6힭RX#�b�,΄qy�i�
l �ņ�}�&dr`�
��[S�U*8��a��I.�(Or�`�삖K�0�����-���q�j\�����O��D%{�R����Ot��O���wJRu� lӴv�@`���:BBNS�o�Ґ�ԋ�$9��@��t)A-�B��UM��΄2���j�Z>r����&:�:ȑ�i��P�AaC�B���g���3,-��L�ƨ��+�n�f�t�3�/�\��c����"b6��æ��	�)���iݹ%>��5V,Q4`���Г�J�Jՠ'P�v��?��?�M>�OE\�`�(X�Z]��K���s�Ur�H��y�'�����On�I�O��xXZ}���B�L��
ߟd���GMY��0� �'���'�b�b�9�I�l�'D���+/_?�Y����i�h����	�֜�D��!��&N�oFtF~e�H�B ��Ԏv�Qe�)F��=Ӈ̈́"�r�0Q�'9����q�X9C�U�$T��OV5a�e6)wzhY6ޕR�lP����"vr@eӶ�o�h��!�q��*rOjx��n*7�M���'��'�Y���"?�!�F���I,���{� �>/O�%�޴��S�9�Ec��ߵQV��0WiL���➜��ɰ^T���' Sh�^�X0�vB�	�]A $+�HY|2Ii�FUp_�B�	���X'h�*��|�uޅ*�dC�	�lP��E�o���Gɤj� C�I
�(��V�v��	�%I*
]�B�*mK
�	��ÑC���'F�+U�B�I ~��9� ��r������B�y�bB�	�L` ���@�\Z���'x�@B�)� *�!w`��:dJIq��h#4��"O���T�'8�����j���"O�PX�ʄ�����hx�l�0�$D���ԫ@��`�[�j� �`��+8D���u���P}r��[j	9��'$D�9G�A= تU�D�^0�A��=D��"Ș\���*�Z4T��D<D�3S�B� ��@�5L��I�d,D��Hd!�i��`�����6�V�<)����U��yw+���tkUN�<�ciY�D}�hR�˟k�������p�<�$�{���`�?ܨ��Q��R�<!&�R%u<���T.6��Ƌe�<� ׵kvz��DM�*v�n) e^�<A��0S��kY����q�r�<yR���
\Z�4�ɇl4�0���R�<A�)��-êA�� `@�	�ȗH�<Y�%��i#f��*����F�<!���	jV���=�xaA�Y�<�&��99>9jeK�|K4i��a�<���9,��X; G��w��9�g`�<yq�%BvXj�΁1���HB�\�<�f��yb�D��Q�.t�O@\�<	p4T|ܬ+4 *���0�L�<	��B�_1�2��>F��q��<����ȵ"@�5\���(\@�<	2(X����1�`�q��y�<�U��_��dO�7���t�x�<�&Y#8��aBM=%�ZL@�[^�<	�h�
Ԥu�9)�FhU��\�<)4	F[�]��,1-����V�<�V%�j) D�p+�Z��A���U�<�1'*��3�MM�,!V�_T�<Isi��%�ԋ�G6^M��p�AT�<i�R�%=neH! �2X����ˋS�<�V����i��9o��SwJ�M�<��)D=!����/�a�7�^b�<�B��5�.ij4(�$�`�;%�\�<yR�:Y�P�[�IK>8%��EXm�<Q� �'��	R��A[�du��F\O�<��V�!ؤ�Ы�c�H �Q.�P�<�PFZu���/�=J�p�{�RM�<u��O�^i�t�\^��؛�h�b�<aP��@ͤ��ĕ6N��{�Vb�<!@h�9��K�dƐtG�i#e�[�<)���t���&!�y�H�#S*�Q�<)n��|Ti�%
�	!�T��+KS�<�"�Q�L��c&�]4��L�<�s�ʠ_a,��f� E�����i�s�<9��t���Q /ʹ����P$�f�<�f�ܙ`�D*g�Y�.>LnP��y�d�Lg��`��&oН�&�F��y�hY<AV6�a���"DX��B��7�yr�I�J���eV4�>��B�	�y��F�p�g�ڲ-�*� GE�y2x���������Qc��ye�>t:���U��ȑa�L#�y��G"3h�� ��(G�$-a�I��y§ŵ��`0�g<2Z��a��;�yBd.z]jmz0lݞ,欈��N �y�n?p���G�R0:�����y�'��Y
��)0D�"���.Ԣ�yR�^$x0B�Kc�M-5���g�C=�y�$�-	bș�NL��9J�fԿ�y
� ��cd�B�E�$^�K�|��T"O�Zt W�������Z�H`"Of�h�C�wJ���"N�h8�U�"O"(i�&X
b��1�Q=%K^�!"Oz-j��@���냭Q-i(��"O� )���vz�(����.U� s�"OP�C�D�K�8�b�E�р"O� 0���)W"�#c�-C[TPɥ"O���ҼU�T�fl!_Q��Av"O
`�� ����D+�E#8��"O(��"A�8�p���H��N���"O"M��bZ�~mB���H�8���{f"ODi���	_�p���E.
aH�X@"OP��e��4ݶ��g�s�x�"O4D&Jz,��G �b�4i��"O�yb�$�5x���d�?��Ȋ�"O
��Vr��ر�$��$ϐ �3"O�%2u�ٚJ�Ȥd9c�`]"O(�@��Y�Cg�uQ�J�)�XA�"O|Y b(5o����)˟e֐�"Ot���P����$.J�7�\Uqs"O�Q�*z2���S̎�bC�h��"O6�����_�nq�"��S�Ĥj�"O���jXd��R�:�!"O���ܥR��l����:ty��q"O�� e<�49�G��i�|��"Ov)��N�U
Nus��G.*�8��"O����� D���·z$�h��"O�A[RK��T���Hd!^�;N]3�"O����D�%�&p�jA�0�aPG"OX4�1+� 0S�I�����q��"O���A�{] �7H)J*5�"O�T��%8��5i��E=|��'"O�5��D�/B�"5&ې1|���"O���v�a�� C���>
S"O�=�͓���$�K����1s"O�Y�T�O�%�8J�Lͺ8���"OX��GO
��`�d�	��)8U"O�����E���ƚ#�8"�"O�� 	�t�F$��A�^�0\�`"Odd�P'��I;��a_���8-!�O�GX�T%�?9�"ub1a�V!!�$P�^ft���_u�Xcboҹ!�d�"�ِ�$�� �`5���C�Z�!��5������Ь+wj<9Ţ�G�!�dŖ\�X��FN��$`��PJU�!�$�/*���1�0�^�B�`N�9�!�+��C�္E��T�S1T�!�$ڸd� �h��_�eP�m׉�!��)4��p�4&V�u�V��E��	�!�dL�4J�OO�8�����K�V�!�d�*��=�g摈pWF�6)�(2�!�Ċ+,B^mi�L�J �q�q�ػ%�!���y@����Tu�ZIcPÉ�v�!�̻T�\��*�4p��4��=<�!�$S�OX�q)%I��Q�a� �-s�!�dV�Cx�<jc�)kI��#�Jd�!�$O*<
Zt3�l�+)�Q�ģ܉�!�DP�GhR(��Iŗ�X��%L��!�d� ���",���Yb����	̡�:\f�S ��b�l�I#M̾�y�!U* ����J�/;��&_	�yi��'+6<�w�ܚ^:�
G�đ�y��
>�5P�M�Ym1@f.[;�y
� �}�p	��"b�D{1�H�C��)��"O��'c�y|`�{`jܓ;�h0[g"O���$�/I��	F/��$��Tx�"O"q�P㑠^��@��D�7?Hv���"O�r	�`dq1�� i=D0�"O�H�EM+i���z��!`���v"Oб�ϒv�
��'�X=z+����"O��Za�a��C��N^Ȩa"G�6	!�d�5C������A��:���}�!򄟇RH6P�H��l��/W�=7!���E�8�Zr*�
�1���}&!���<[�0����+'��9�un�+ �!����j6lU�S��\�BU��!�䇟6�@,  K��t�r����HN�!�?L2�PSkC�q}�I��F�25�!��Y;��5�a�$_���+>y�!��!H.m��e�K&ƁP�yI!�d��o��pp�hEɵ�_$=��5�ȓP���5�ڈP��ѐ��\��Ņ�9\T�h^�֪��e�S�lنȓ/��L:����V%�F�&Bm���}�r��*x�z@K��H"�B$��;�aa�Ǌ,*�B݂����]r���ȓjfd�Ɖ�)&]�4��-%����I��h��(�"A�ٹd�O�z%n,�ȓb��d�!�z�$�!c�ͩs�jȄȓMˎ)�#��=v0���+�'S��P�ȓT��d� ��2blچ�>�|�ȓVu��pPŝ�4�f�z�D!3�,l��{^��p�%2�"8���ց;~p�ȓc�rٸe��6 �*$+W ���ȓ^�� X�!LSZ�!C.�mg��ȓ&
�SN�(�l��A�����y�ȓ}_���T ЍO��<��#]TKT�ȓb��� &��;Cܾ�Cp��KXd���tY�4LM&�T;v嚖4����l��dt��f#D,��_Lm����=���%ʓ?�����S({n�5��%���䐅a�i�,Cl�@���q(�Z5�8��Ѵ�ߌefdp�ȓf�2i��/׺<�	�&9�q�ȓ ��B���McB	C���4���S�\l;����>�(܈wcJ?<��ȓcl�Ԁ�)!�R�P��ę� �ȓm�`�ӑ D�F�*TȤ�̜�(��ȓ"���H�#�4�f��YͅȓU��¡׎t�H�(�dd�ȓS��y�F)�%2��k �y����h�<�"�ݓ.g�4pd	\���-|4�5��J��PTG�BI4]�ȓe�d�U��ð(�G�ۙ#�L��{p<dQr��IR�`�(ߒF�HC�Ʉ:9pQ� ~\�(�!G��,B�ɻ!�H���Y;�qISرn�6B�I�A��銃b�\;�� ش�>��ȓ> Ĺ"��B�h>!�ԨV Y�Շ�d�:!�d�.B��⥣>qV�!���)����!�@���A9~4����C�2yS񊏝\��`�5��P�$���*��}���D��2D����هȓk �����\��=# Ǭ`F���ɫ]����3/�1�.�9�ǘ��1�5&�l��{�!����5P���)f܈�J�d^!�65���ڥA{\�3Ĉ^#?�!�� N"�ƳN�*y��rP4��'"O�Y��@�@r�A?HD!�"O��S��u� ݂4o�7X�J�"O��ҮƎe~B`X��^�^cNȂa"O��JU+�3�JT"T'��o'<��X�<yB�0p�����іMf����VS�<)�j�|���q�/ʻ�$�#��n�<��>9�B<a�=8�� d-�Q�<���Q�E��q#V�,0(b��T�<��'��eM��cH+'\���LZX�<���9FR�r	�)�0��ЫDX�<�Gf�m��]��/�&U� �)�
Q�<!#��Z3��p�A�o�m��ll�<aB	�?�I2҃��J�zb�Yh�<i��r�p�M�?��#�O�?N� B�	�6^N�c&�Y���p)0��N��B�a$е��F���I����"?!����(����0��n,�dnP��z��A"O$�s�f��	�&�ĆQ%�ڴxb9O69�Tb/	��O?���M��(A"=�5�;3m(�g�=D� 	Ҋ . �G�
	�^P3 �>qɘ�x�VI2���p<�Ƥ�;,Y��bPL˞ �Bbt�pX�� ��� ^��x#�I�;1��y�o,.��E��������^p�ҭ�
A���P1�.��Dx���P�4�↭KUTC���E��t@�jw�S?�RUI��ybj�D�ZY2�E-��y�C�[68&��I`����0$c��|��9O��[�l �pP��ڥ2\��1"O�Q%��>Cb�`�lπ[挍2�chӄ�c`P[���tÌ�&rG�-���ʕ�Xg�-���=�q��2j�`�c�%�!T�)A�	��=`ڵcŅMx*�{ĉ�2�x��J�f�rO�qd=#��́��'O�bw�;k%� P��9q�4`�g�ƌ%P�ͳ"N�v:�:�"OB,c�H�T����B���`u ���p��F�Z^,����>�z����w�]�W��}�p���v}��_=$1�P�\�?�\�HaO�;q�(o�f�*���O�\��p�'�v�hGA9 ��A�t+�58��:�(n�c��G$��f0MkεZ\.]I��&.Æ�D	���p?��$Ag`1!�Ø(e�"�rT�$�I$
�� �:	��`F,�J.D�������)�~-j�'Y�;��m)�"O�IgO��R&ƈ��'�|�� ۳ �4v4)(aj�((�(���=��>��$)���C�υ�b>‣g�77C�I���3��Jy�
P*�#��͌u��#�e�#����ً���Q�p�RLk)����oڼz0Dh�6�O�҇)R�58M+��Qی袤@S�m�N������}�0���8�O��{�o��>'��jF�P5�*R�I��*����Ϡy�N��фA��/�D�q��� Hjܛ�g1J� C�əuȊ�[2mI=Cu@��ĊN�m�7I�7˦,�c��sX�S��Mk#�^$p)P���J�;V=��/�~�<���*rT2|��M�	܂���*|y�a�5�4q	�*
��p<aQÓ1���6o�J��d��N��p��O�Z��`b \R�����[�[�� 9��L8&���'aS?�<庇��9L�b�����6hٗ�V#$��HW�E�B���ұI۞\��!8��L�:l:���}����P���5����B�����J�.�����
6���1 �:(�lX���)~1O:lY���9^\��a�O?:Cx�����']�R�����,`�g�W�
d����8%<%Ұ��sU�i ��εIZ��Q�[2-{�I0Ua�*h\nZ�����'�\ifn��/���E�����D�<A�A�'|�����P\��3�j�Ѧ)����w�^ K�o+X���1�B+�sîL(�(�-3=��y��ԥQ��鉉>�r<�R��8lFz�taʽ	�\Y�E���W��p�B��F|ܚ͝5��?�dV�(e�D���WC�p�d�b��UG� a���2�Z��8�l:��̨p}HL��պLz�Ȫ���/6$!�œC|8rc��ed4)��N&!��<(3��3gq�XDB��0��&�7�'��ɴ,[�)����g6�80$#�NPDC�)� ���p���K�(2:�삤�iPn�2T�J�!�IGB�}������!��z4�� f��B��S�azrn�R�ΡBѭ֕(��7���m����יq�XpPB�R�;ch	لO(�O�b1�7o� ��n�/J��ӄ�d�
(�҆��06Üq��{��N|���{�h����7SlH����h�<���!>[���U�1%|��/oG^��S�����+�P7��[��e^������:�vx�OX90�!�"�,D�Dr�LQ�+p�mɓ�S�\'ԐyD"u�)�p��9�t+��
�Ȥ���	('L� 8$�N���s �LN�����v/�8�f6�9`��J)��Y�'3,[5��6�
apc��b؟H�3kI�>�v��Ń�Fxx顶�"扅f8�頴����t�j<�6����N�(W|�*7C%Y7 tvΓ��y",��4�܁	v'6P����u��(K���@7R`7N��Mã�����Ê-;�)�v�����ꕧlH!�PE�� @CX�;��!��ˌ+��l	�<D�ju�["d��p��
���O�X����D2]QP
P 3C�A�p�'�.(),��� X9���%tMNS&�%Gan,���iv@D���� E�X����AVv��"�PY���qC�a�1O@��sG�A��0fa,.i�m���ħj\ȁ�� Z�'���v	ƂZ?l���a�xe�֜E�`8@c�I����B�q6��X�����l!����'($Q�Q`X�u�,��cH�3�����'�D�ӧ�k��y2�
�,�ƙcߴ:z4Bp)�&fU`�a�(S� �G~r��$cJ�*&��-l>r�O��0=�U��*ߊ�ဣG�;�(%��"82��͙�z�B�x�n�p�)���'Є�갏ۈN��iV`���ư�	�'��T��E��@��m@ӡם�~0!
�'�����	x���q�ټ�`�	
�'n��A�7a�)!X!4E�'bzX�C�V�e:���<Ib�$[�{��q�ayR�`�2i�֓k ��Q$�9��?QT � ���2�l�-
�8�fN�	����&�	K(<���"�Ua�a��	%�H����t�'� �z%�I5v�&�>I�����
o���$�q����-D���nZ�Gfv��ϛ	��0�A���<0�+Ȏ0��M�K<E���E��쉆�#0�p,X���y�bZ�JD�4#�u� 	Q��d��0t�`f��<����)V?~̛��7�4� b�a��d����NoN�j�%Òu�W?���4'2}�^��ēt��×b޼*P�����G|��>#xR͙SM�O c�[>�E&X�kᚽ02�&Ϯ�T!>D���wc��5�.�`��497ҘQp�|�nM���_��`�"�i��)c�s�̨��ŕa5�IZ���ew��	"O���⪛���(b�s�*d�GEK*m.��)�'��a�L�;s�R�?��3�?)���V>C��QBP�˟&����I�n��r��_*�\
��3*�%	��0!i�����U� �8���ArX�T��@�99�������r���L,ʓL�U��H�y@�����XGr�۩��PCQ��*�IT�7� V"O�
�mV B�֍ �J{�YkN�`Zf"@b�("�u���q0�D����%�� ��C�"��0W�^��ȓB��x���x��J�l�*���W��P�C#� ,�x"��N�����0�YS�Փ*HR��I�S,a} �$k&X���&IHZm�D��5R�
��<�~l���Ŷ�D���	�8e>m�rÙ�tB���a��+�V"=��
^�r�e��DCa��Y�4��|�u�\�sW��&B�v���r���E�<i��Q�����!�,��r���h4h�1|�.����,o7�-F����vP�j�{v/F9`��j�'���@(�6J��!0C�tH�����?��HͰ
�R 1�B����	az6 BH�2J��|!��L�X���$ƿe�����k�l�d�I�eY� ~$�G��*<��rE6�OV��%N�g����@� 䮔�6�Ib�xrܛ� u%>i��+M��&���6 �i�TG D� �CPf>�5[֋إI*�"�<q�dI"&�H>E�4�*{����Ar��-�-��y���2���&\l(R�1CG�ʸ'�ܙ#���� P1�pC���!�<Y��2`"O��� �u�����H�Ax��"O�er1C@�?(ɨDH�<H��H"O�55M�8����[�0Lr��"O&�ہB�<%�rda'cL$��mKV"O��+t*V�
�PQ���-=�U�"O�F���b����m��PI"O��#�"̸I�rEO�i+�t��"O�I@��y�(|�ڗO����"O�8@���1�Ԉ8�C�1���`2"Oz�(Ą!2�Ѕ���(�x�*"O�%���B9<@r)#1O?!��\��"O��r+M')r�E�#!A�n��"OR�s$��Q�T9�s�[�E��"Or�uK�0�Ƚ�1EK?k܄
T"OHΗ1�X��a�� �(��@"O���%8/��IV�ћ�᠒"OlPpN�(:*��b��v��<�E"O$dj�j�4/H^(!�` �]vv�;�"ORX�*� ����e-�x��ݱ�"O,q_%[K�(x$f	+M�N�t"O�.i�����dƤN����"O�i�b���1
ج.���c�"OTbu#�%Qd,�2d��0#"OD�1�]�K����f}JA�"O,���f�<.��uIf�ќisP�"O�E���ik�КG�P1H�#"O�E�NQ���p7�sRU��"O@��W�|��-�`��S ����"O��ɒ��&ph��V4�&$"O����O�/� �P�Y?_��йv"O���Q��]��x�G1;�ȒC"O>Y��,��*m���� Ȉ_���C"O\]2աҖ$��"�Σ!-���"O�`�X6Q0J�*B�.'&|}�"OxR@ �O�dh*0r��"OB��W�
;�f�)����@y�4�"O��c�N��8�l�"�ow�X��"O���,Y�@Ɇ��0lA��`"O�X�g $�B��U�J��
Q"ONhb@ �{R�B���&o���ѵ"OH�Ja*�s�.�ȷ���t�"O�$����.���+.6����"ODl�BJ�@��s��[$N	V��W"O��	4�W�clHػ1�3JM���"O�1�!Q3^؊l���7v"�}�a"ObySQ��������M)�ڰ""OV5��h�lP���f/Q/a�hY"O:i�Ġ�S& x�fK@G�L=93"O��S�M@0��q���Z47��P�"OL�����������k��"O��>X��d�7�,;t�$�y�k[�.#�=JEH	�9�d�3�J���yB#YA���ǠA�����P(�y���c"�h�U�N�|�)�����y�gʿOZ�1�'�z!�`{GÄ�y�h� '�@R��F t
0�Qm��y�GǤ_m,�oJ�:$��@���y�%�5Sۆ�h�mм/���	w,F�y�F��~'~EJ4��,�����*Ƃ�ybnD>�d��H��#� ȱ�O�y��< ���X7N�Y\��`�&���yb-�`K��z@ᇖ%��K����y�+�3$�HS�ZЪ4�7e��y
� v� �"4�	S�ȅ����4�'��9sc+I�Nź��g��;��9ٔD��=�������1ˠ�����pW��8J��RVֳ�*m��`th`�NJ%N��t"#a.J�lC剿rH����BԆ�f��ą�:y�*B�I� ZJ��<����EgT"VrB䉨k��a�K�;K�55.�2)��dn$�aі ��?�B蓧"�@�!���>�2%���Sx������ڷ1!�$M�b5�fM��c���"i[�t !�����d8���?z��"�>�!��T ,���{����p��B̤ �!�8;t�cMޥ@j�mK�I1�!��=hU�����A*�X!�@#!�䜁��j���6(��<;é4
!��YB���B ߒn��Q���[<5�!�� [��	��4
���U//<=!���39̌���MK�F�ke�7QH!��8��T�ak�/J-8Q�C(K�!�O�*��Pڀ�O�	
�I�N��Z�!�B�N6B���,��	�ι0�	9 �!���#��1�Y�X�����.��;x!�ā�o	�`��+Ϻy<8�a��}K!�D��d�t�z�d��1�ɗNQ$",!�$N����hWn�O��<�bl�< !�D� �LDe	�q�ư�Ek���!��P�L�x���?W(F�H�/M !��5K��,�҆��7@�*�!�d�]�P	���J5��n6$�!�P�<6�A�s
�N~����N�Y�!��F�X��M �Z�$�����cҲX�!��  K�Lp8Z��Ѕ�A���!�d��@T<!Y�Jv�X���(*�!��- ��3�E���,$����H!��&i4��e��m��8؆ Ǎ>�!��:6�z|��f�Ol��*"�29�!�ăA点
B)D5A���u�KX�!�@�e�d�@E�1xhU�N�w�!�d@�_{�t�⢚�^`0TS��Gw!�䐃	�*�Z��PyF�KG ]TT�ȓ?���ЈV�����e4���@6lp��_��f� *~t��1�0�1��ԣ�x�pC�9��@��!:d��,�2�֘��mC8tp�H����ʐ��Nb���#E�̄ȓ:K0d�Q#�TЈ|��L�O&���I�`%d$ʂl�8ieD�F���ȓZq�(��W/ ʘe����u�t�ȓ�6,Z�/�fʜ� �C��+̲���6���z5y�~���� �H���^=.M*ւS3D�J�#�f��[�t��M����J4s@sRh���0���Rd��D䊱B��-æ�(4E�݄ȓjJ�xɂ�\�Z!��@F�L �p��~}���QmX!W0�YŨ)��݆ȓk%~	�c9����f�Ƀ.l4؆ȓ.���e	��8��͸`*�@-�%��Jb�@�ãc�n��"��<D\��A���X�#�vQ���Fj�Bм ��5�\�n�Ќi��ˊNy���ȓR� q�Sπ8D|�mY�e�/\��ȓu��P�ǚ�xjh�b�IƆ7�Ѕȓ&2�X��l���E�]�L"(��.��ద�
� �\�FG�a3h���S�? rhQUm?���⡇��!�. B�"O����
݅ek:hB��+c��s�"Ol�D�:o��,����A��+""O���4d�&�(�B�+-�R��`�"D�h�5�G�0m�u���S'.���?D�d��#���4�d�w3�2D�LֆZ#m�U����
�0�!vE2D��#�$��9��1+яN#_Q���b�/D�8�f�V��r�8�Ê!��M��+-D�(��QjؾQ*��>���%D��P���h�le)�(�P�d8�tC/D�������4��M�k+N`�fg0D��sc�S� � ��d@΀qR�x50D�pzwe�$8a�����0�>���/D�P9 &D�:�\��AJ�f�\	n/D�\�À�^�>ط��:ՠ��g�,D��!' ���a�F���K�x����&D�PxPfç�v�Z!�G�q�0;%�>D�d�G#�Q�l �3�HhG���rC<��(�O���Ȍt��c-�;��!@C"OD�ag�r����#��0�\I�6"O�m�R�3��a2G�&^�Xق2"O䤊e�ս�s1G&;��3�"O���(H�z�@���� s���P"O��@��I6]�W��F��+"O����"E?l����c�އ�����"O�j$)��V����C�/}FE��"OxP��.�	\f����ã#�Z��"OT���+�������(�f���"O@`��f˨@��\��AحP�Fu`G"O���$�p�|X�oܤ%��83"O&(���F�GՊ���m��v�v �6"OnH��;
&��d
��pڴ��"O�<��H��T.>�l���"O�-`tᆑ}M����'۩jxV��""OL��$T7��
�f�)]
U��"O꽱V�� �'�P�%+(L�b"O���3�K�0�!��M;^d�y�"O85Sv��	_x4oS����1"O\�����z�Q��k��� "OP��%��4[z�QU(H��);R"O�0�cC4�@Qۥ�����ȓ,( ��#�G�e2~�!T�:�x��7�a�� �8�K���R�ȓZJ}�E�cl��Wb�&A�"��h��u��)B!����fn�e�ȓp�X� ��H���@��	%`���Z��q��� &�Z�U�n&ĵ�ȓY#����)�/(u[Q�� V��T��Ui �@�S�b	���S.?��ȓ(�LB�b� *f�b�.	�z�J���2��<���!\*Yj�B�|NVU�ȓ������]H.Z�l�ˬ��ȓp.>D�r ެB���t��8*�!��@h��P�1/P���B�	W�p0��2��X�+Cb� E��8}z�ȓQ������O�@�aE�ǜŰD�����(��!�y�f^�~��ȓ%��*�h@�0׮�:�䖫L,A��^�P4˂�A:��A靻2+ང�8�`�����1G|��ف4)}������OҼ��Q��Ȅ3zLE�ȓ-
x���ˍi���r4lHY��܇ȓ� ]adL��G�Z�B"��)�����S�? ���El�C�,,�	ѹZ�L���"O�x�b���iq�HT�253"O�y����	3�L��4.�&:���"O��A���>.�6AcQF��#�:y�"O��#�`J�\�ؒn�-=�9�"OPI!�"�c�:�@t�͈k�>m��"O��٦��.h���W�b�@"O°��,U$!@��T���B}|�إ"O�̩#H��Z�+��9�xDi�"O��[�e�.O��:���No&���"O�%i�O�!�rj��F*ʨ��"O<T��!L: �r�@D�t�j�"OJ8�a�[28��8��"����j�"O���A�=�x�"Vb�HoD0��"Ol1�`@;h�8�bE+\@VX�P"O��Xg�H(G���I��B= ��V"O��H��]>2��hピ�cٚݒQ"Oʘ�񄓘
$x�� Ov�|Bb"O|��gΆ'9����H� (��"Op�BL��X.�b�ϧ.�(�Z�"O|��"����.|! �D�9����"O�l;��Ωy6^R��3#� }�#"O���u���$�P�#��Z�o�`�`�"O�D{ť@
.~��-�rʎ2�"O��#7-�#��t�.	�f�"O��i��R._$�Y�f�_C�D	"O��i�
�*[�Ta!��>��kE"O\�g��I����:�Hxc"O`9[!�D��(TB�J�C�.d� "O��Bn�#�$�{ M 		�|�d"O(�d�E",u����$����a"O䄣��F,8�#&�	;�� 0�"O��Xk�:��Q��O��A�A"O ���c�@=L�2��]�6R��"Olk�J�V��ᑠ�0N~ �s"O�x�0k�6!E@��7,餸��"O�U��Qch)��䔭�>Ԓ�"O$HZC!�U�*�ʦ#Op�4��"O�X�@�E,���+R�.ZLY�!"O8큶$�$zz���O�mY�"OPxW���K�$�Ң��*<c��P""OL��sJ̑H�:@���R#�8��"O~!��#H,U���P��K�hb]�"O�T��D��pO��S�O�� ���"�"O�ҷ#��+���K��[�c�V!j�"O\���n%פd��O�-B�p��A"O&��v�Eo�f9��� KsT��"Oz0���+['2UA��ѻ]��"O����.���K���#B֍A�"O\� k�E�~����̈́q1� e"Ō��%үr�]!�Iհ$6 �2"O,��φ�+�b!r���=��S�"O��04�c��8B�K�Q�Z0�E�N�<A�L�74j�5[
���B�[�/�L�<Av/A��h�ӥ�`g�q���K�<Q�:��+���==�$��m�m�<I�G)Za�ې��%/�:5p�f�k�<Y�J�vL���m¡Hr�;w��g�<	��e��g���]�x��֪g�<��ω�S�4��/܍��	x��e�<�6i	�>S��:W�ӕtz�%a�<�ǎ�Oa.�r�A�N�L9hB�v�<�d�[/W`�	�;^8�Sf`{�<��WWܑK2E�Ţ��"Nt�<� �Q�ע�Jra��#�%��	X1"O�T{�BK�$r*iJ0LQ��\�S"O��3%�ȅBΰIk��G���h��"O�u�2lֵT־R��-\sV�s"O��EĊ�-�DdZ b�'RW�UZ�"O���OY��+���M��'"O�A�S=�a�.�*R�n�`C"O:�#&K*$Jdq��[-gD���"O���FI��$�Px��5�e!�"O4#���y4�d٠AG��,�6"O`e��֋B"z��6��'��i�"O)�P�Fx1��@N=V�.�p�"O$��'iP���Oӂ(L"�"O$��掀2lzh���	, �"Ofh�V݆w* �!��ەX��Mb5"O���W,�>N�dT��+#��Ƞ"O�����*��m#"bڄ_
�[�"O��!����*%`栓<dִ0p�"O��A���9D�,s#"
o�܍�"O6Mx�g&3�H�+�`�K�4(�"O��F�C;�jhD!ʦ^���"O�����
j-��P`�6ro�(�w"O�4����M}8�[���^e2@3�"O��@�ߋ���X�D���i�"O �@4ƀ95�$��l����&"O ����0Gx�#�֐)и0�1"O��eI�F�y�JO���D(P"O6a`2ݨ��� �8|�z���"O�� f��3����sND��4 �"O$���a��(̘� ��+�$X��"O�<s�m�tx�Y���ݡ.�vi�a"OJ@1R-�=z?&a�v���>�G"O �Ӣ��a�80p�i��wct���"O>S�%�Nj\I�W�_XR��s%"O0�81B�/|?FE!@H\5Q0I��"O�k$嘤غ'�¹X8����"O�쳄ˀ:^�2��oѮ8�L�h�"OҌjů
/<��X�s�ԍv�X��"O �*�9>�@ �0%W�b�(`A�"O��[qbM��.i4�����C�I�!�N�H�I!�._�ѴH��� �!�N�d\<��A�
#�u�AO�a�!�d� U��3�g�*��SPlH�t+!�䊉^����J�8ͼ]���b!�$]dUT��!〞p���(Em�I
!�� �dA��ɖ	LAm3sΏ�>�!�$�Pi `�۰~�B�(4��IjC�	��&�;"�Y-\�S��םcMC�I�|bbB���4��`σ�"��B��(]��!ZwB��b�h��ViM1+5�B��:}{j��o
��5'�`�PB�<t��8�/����)J`�ց[PXC� ld�0#KܟKØ9� OW/t|XB�ɿ2-�m�KƖ([�1ZTG�*#�ZC��
�!��*д'���H@��2*C�h���q�ʕ[.Ry��˒O��B�7p�&��G��{
~����t�B�I�{I�ř#i�s��
�(|�B�I�^Z�tZ7�D m���2T��6$�C�I$�f�:1!�
n� # K�$tC�	d�,��Y>C@����0y�ZC䉋"�\A�?	���CwO�=}�B�I���0Г�]"w�X�p�bo�C�j2F�`���h0�ʥnH��B�)� �0�&�D�^�*݁р�.6΀k�"Ox�	�|������M��@"O:�y��e�8ܢ!H�o8��"O�P�!�%Y��x�@"
�\Q�"OPA���5p[���6�Wo����"O�|r��\67`u�/�b8$��"O.@3�iV+�Jp�c�GC��c�"O2Y+cI�N\�a� Y�hx+g"O���6��q�VA2 '��N�H��d"O��
��W'W��Q�3���~���"O�	A��@�\>�Ly�呁�H��"O�x��bW�`�|(7��R�е��"O^}R�*�Y��;�nP �0�P�"O:X��8S�v�0�.Q�f�~Q�U�(ی��4V��$��̨�8F��cL�B�ɾDd
�rt`�T���"5.~���O^��D٨ �H|Ʉ̨L�tSr��&'!�D$�\\bL˸34q��	�X}!���VTA�Q�I)P��/��Py���`�������� #�%���yҮP8&*���e��z5����R��y�+�`2ȡЄ	x>�S�%��yrF�ox��p�ݯ$��	�2.պ�yBLQ�q��(	��L*�  �@_�y�f�6�6�"��H�v��p��#�y�H3I�H���@�kޜ���ą?�y�AܱhR��C��d�ARD��y�j��d��-�V���	��$�/�y�� 	 
�k��JR���p�G��yb��c���02f_�F_�8I@ŉ1�yG}�� -ۣ<Z�� � ��y�*�5?X����ڞH��h��y�큖Br����틞qg`P1�OA�yR̕�x�\�t�m���5 ^5�yR'в�
���ꍱs����ɂ�y�1sH�4)�(E 7��ᵥ��y	S	 ��!�� �)Kd,�u����y�NG�(�rP*��

kV)	զ���ybB�Tn���"�{1@,���y�I �+	�V�3������^��C�	~�@�j�M�4s��!ۓ�Њ<�C�n�Q���3_��˷"Qsk�C�	{����bg�+Wn�R%�Z�$"�B䉳U�2@1RgʶAoJ�Kr��4U�xB�Ʌrx@䡃��/q���&MI�"*fB䉩[�bP�A,�	]��4�dh8B䉏i&~�Sc�t�^�j�*��w_�C�ɮs�����űe�,�z�LO7Y�C�ɉ<�6�� @?�D"��bz�B�	.����JH|:H�A�O,�FB�I"����K� C�� ,���fB䉨4�l9�De�2V�,QCM��a�$C䉗Z0�j�i� Sx��5F�1g�C�	����b��:�"�I3�D>��C�I�q&,Mr�o\��AA �D�'jC��9Lf��FF]"<d�ǅ�	�2C�;���g8FR��'�4�&C�I�*4�"7�ώc��pY� �74�$����D�84O$QH����A��mӅg̘,	a~"!�M?A`��jg*h�ܺG���@�<tn�k�.n����M��#>��	 �8��%YCE+>��QҢH-�����z@�ِfNΗ37��@kI�Px��̓V��<E�4o�M�ι�&M�:4y�+��y
� ,� �U
G�R��?R���>�f�'��@CK�-`��:�� `y���nw��ɿn"b�ؠ��J�ɐT�¼�^B�ɾM.�<��@�!e���*����F�\�>q�%�'o >i��K�.*�Da1�e��5��ȓ ��xp��]�ĕYɔ�
�����hO�>u��ϝz�V����4�\�P �:D��"/�-``�D�&{�|���b,D��S�I6<�vLKE$Z�����,+D�ȱP�O�j\����LC�@��g�>D�\��س�<Q��k�>�QT�"D��Ѓ6�\Q(�$$<4=b� D��87��Ʃ��jS�{����<D�L '��=�V�����i֠����>D�t���Τ8�ژS�F�-c-��B0�=D���5�ٴNqz�������L� �O?D��Kq.�#|���!�
v�AH�:D�p�D$H�_�~p3���6uޤ���5D�pS�T2$	�љa�I�Ɣ9�2D�0#a"�8���b7O"�H�I��,D���E�h��=Pì<0.M�V'D�X�B��}�*��"�PI�d� �#D�hZ��T�H� $�P�d�
�zL"D������,JuB!�B�)L���#�"D�(��zf�E����j��$i A D�x[FI�'����Fl���K�D D�ȁG �xLK���c+�����8D�@��
_Ha������6�5D�г7b�k��feR�'KV(�R	9D���F�z���ؓFQ=5�	v9D�|C�,�Y\!��,B�+-��2��5D���f�3/8��s!�W��P�R�3D�L�C��;.�t�
�҂;� zq�0D����b͌�b�>���Y��$D�����
4[�Xp��Z/��@�B�!D��+��y���K�`Ύ ��O:D����"׶�8ѧ�ʧVr���6D�4yp-.����F��$&R4�!5T���B�	M>��5"K�|���1w"OL��Q��a�X�Y�� �?�z�z�"O�+0�@$'^pp�$��r�����"OHu��c�,tP ���e!v��-!��!`h,	�R=g��VKͿ[�!�dZ�Uhh�!J��'�>dò��[!�d�
�N r��Z$dJ��0+9V!�19� ��+`S�]�k�>O!�d�z��p�6{I��k\j�!��8B�t0[�'D-�vu��j?�!�$��%ꐨ�C��@u��[�!�d��k��i��+\�J�4 Q�	�}�!����(|(qa,F:��� eC\k�!�d�{C^���섴_}�!�bɘs!�dD=K-���'dU
jb:�YRa�!�̶>��E�N�bi�ӓ�ɸ�!�D�(���1�A�*`fh�7iV	tx!��~k�U�r�B�7K�MP3�I$b!��ћC�JX���ء�~5���ؽ[H!�ۦ~�H@ ��H6`q�t��~+!�d�;# "\з�D&K1R��aR!�D^>4Z&yc��
��P�񠗇W�!���ˬ��g�n`�aH�YP!��!9�L2w�	-I�����(!�d�t�d! ���}A�]���
�%!�$�)�pX
s�W�'NQ��ͬ9�!�� R����]�k��Ҭ"i�ar"Ot�ip�ʧ�.��B��BZ���"O�5j3`��|	�7C�$I��g"O�� ҁƉ1�,�p�A��*���"O���&�����ԛ�&�$y4T�6"O*�Z���F{�őĊ��qY�t��"O�y�֣k�\��7锄UIz x#"O�z���n=�T�c'��s4bA�"OAq��&|J�p��&M�,��'_�!Tќ�S�R>N�ڬH���A��)��87�>���O�1B�n�!'��aB����q\T�r��3�ʠQ�f7B~��zT�9*��B�/B�rQ�L�TF?jx}S'�.��e@���Bt�qB�q� h�c,��	bWa!��$�d�����j1n�S,ؽ8��`S��R�ʕ���Jz���O���1�	d��(�#gpA���M�g���c����IWX�0� �.Go��AR�(
n��r�#�?9Ʒi�N6��OX�oڠ_�a��4�?�(O�N�P�R���N�
0�2������'����A�ṿ�ȏDB�0�to��2�`�Hʳx���S4'��1ڜXpV,����M�.��נpb��Rށl���R�\ƾ��T�ݟQ�Te�E�آ���v*���'�H@[��.��g"�S���x;�e�Ux|0��K��^�<��g؟��R��b���`ckGW��DƯ���4����@ڴo\���i��Ipg�8Y!�1K�6���k�Ѧ�� �$�M������|�M<!t# �V�@'���3b^0D�^B6����#R�R8�o��7�@
ϋ17DtRc�?�����a�D�Z����A9l���i�L�LV�'mڝI����JԋcO 2Ѧ�q���Z���PP�F_�hݺ4ˇ!Z$<���ǳi���[���ϧ<��k��M����2G�
)�"��u�Z�B�a�K?���hO�c�#`�) �i2Ù�lj]��5�^�&Oe��Oj��p�Xъ�M�uTeI�25$E������D�ey��lFX�L����-��e��&5��	e��.H�2�=VZ���˓�P�bL���l ��6#�f�I�+̔T1G�.1����GB������iRƬp��pz�����~�� � Y�2 �p��<��OA-��F#�
���s�#J}bO���?�P�i2@#=A�OL SFl�U٤'�77����7�>���)�	�
��h4�/��0����R��P�i��7��O�im�ğ��?�OH����U�AD��~�:Q���0u�� ���'��N�*B��l� 
�
���S8t��C�bB/��l�r��/0����*$\�8����	/ߢБqRMݖ���Z�u۠��5�*v?D�Yī�"O�fE�$뗤]Pt�*���'?V��*����	U`:�����9[�i(҇S�gё�X�?��O����D���� (�h�ͳ�"Op�'?P�
��f�<�v1��O�n�
�M+OV;3���I~�S�y4��F"ư}{�E��dT�s���@���S�hҢfI�&]����_,F%q��@�C]J���-0(��LU�N��֕$]�Q��֎K�j-�Ȩ'��b�z�Cѯ8]��f ��A]�Ya�F�<���b���Ft����d�#:���l��$>qo�"r�~��CE/3jC�"�=OT)�����?�|�/��'f�D�8H�,2��u�)�p>�Ժi7J7p�<��/
.6��dzr��N�4YW�Û�M����?������'$ԑ� ��   
   Ĵ���	��Z��viĎ:B���C���NNT�D��e�2Tx��ƕ	#��4"�V���Yq�m�Z�l#��j�d8�&Bd�����i��g�x����M#S��8��
4c:H�;=�"d�@�'�����ٚ*Ш�&�TJ��\�u�6H9����I�!l�A@̓���I>+"P��5iJ�(g�b��]�&�� ��#^: �_��q��̍P|ta�!�<�b,T�/�l�A�J}�앮h�`!1��<	5|Ac�j,�"�0)*x��������	%mʠ��ş?%`��ԛDLkՌ؏Y)rI�7�6Pŀ�����p��D��E჈3�Rj#T�[Fnq>�a(�&En��p� �3��ڐo�� �W���8�$�|rA���}&>1��?PX2x� NW�8-��� �O�%ܽ�,CG���8����|rI�+��pGѪw1Ka�yC�ē�Kߝ�ēf<��f��j�I<��0r����@��z%�9�
�x�\a@ ��?a��0U�x&�0�A�X8H��O�����ЧaC��ao��u����`[�R` �N>T͈6m�2x&��Wh+i�6�Iޢ�zs���F0FmԹd����f���X�I���	.8�V̺1����Ă�|�"H�a�T.�R�[�f�,����(���y��*lR���Do :^V	�hɔP�bc`�=��9�h�s��2s�H*I5�Αf��@�8O�`�O�
��E)"`
5B�*���V�@����V3Q��cŜx�kx�Y�EG1r��i	�+���~��W�'� �%���'�ʅ�r!�2�\ܳ��m+64wJ+Q+*:>��)����z�ƙ:�П�ա��ٜ>����	�\kcjF�=%���7ɒ�[��'�%K�e�"��h�L=`e�d�	q�r1�-��j���`�)�Q �M?)��Oz%c��H=%�1O��؎'hx9q�E�  "�1r���2!��'��)�@ ��	�dB�	 D� �  �c����ybn��yL�#�B�:xc����A���y��p��J3��n��e�']��y��������J�<;���Zw��3�y�
ґ_�-��n��"B�@p�Ӄ�y��M�_B(Tb������Bi\��y��� *b>Pc���M"d:�yҠ�"JKfUzƊ��2ī�^9�y��'s0����8�(�[�CJ��y �7^�8���n;&TB��IZ��y��T�za[�U(   
  �  j  �&  O-  �3  �9  ]@  B   Ĵ���	����Zv)���P���L_zD�R���\���9��ƕ	#�e��>���x������ڂx�'iLZ�<�ɋ�P4��wC&9��4�K���b�� �p%�%���]	F����(� @PP��]2�E���W��Xҵ��7=�ig�W�N�f|p�cGv�rkΊ@��uHT�� 9=��6��!��|����Z�6����
L�b������
!�|� ��	�e!����ϒ!6R��ý� 3��1�?Y���?a�N�n�O�Y�@�M ��y�+�?d$�s�Ly��ɵ�p>ipn�)2�찳�R�:��@;��Ey�*O�p>�@��:�X(S��<B��X{�b�y��]�?�W�''��h⪔���X��X�[��Ȑ
�'q�ȱ�+�#v|N�C��z"U|�%Dz�O��'������"�zAg�,]���� �6X �B��'IB�'B�z݉��П��'k,  ��(CC� )&ƒR܈|���34�.�I���x��ov�����S�y�tЃrC�c��̄�	a���$���V8cn�g䴑���o�p|�ȓgL>�p"��-��s�V�Tv��ȓ��Uu��$[��z�Fx]�'��6m9���z�.�mZ���I~�`B	r�X�2��&X��"�����鄫��|�����(�G�ğ��<��P���X%\�\�l����-i�$�G{B��.���P)�ƌ�ᔅ���J`�z���2V
��$�|�O�~,Pd�N�v	��t|��'����m��8Uf,��fR�l�x��}��	2D12�����CmE�08�,�a־i��'M哻�|��ğ��H�:Aþ��+�h��|z�M�M�W��,�?��y*��O|+%(ƆsW�p"�H���XP�'ż���� =O�r��3-�B|�e����)�� u��$s�)�B0ɘp�+T�4P`"���2�'�,%)R��6G��,�V"FX�#=q"��"GNuP��aS�kg�ۺ@�\P��4�?I��פ	�Fdш�?����?Y������;1�Mf� 4/
B�* ���}y��ݧ�p>��߇{���4�Ip(�� �yy�G��p>�QE�@D<Ib5$�R���ʚxyR	Ր�?���'�x�"G��s���f��E�KPt�<���@�Z�EB�ܰR�����Wڦ峋�4���O��1� �zp,��+ݲN���R��!~�DeJՇ�O��d�O��׺;��?Y�O�&���Kb�'�J,+�Lb��+�5g�'�Ѕ8�'!��LC6=�
��`�^%H�@-p	�K�@5�I�	v`�����l��A��aX�8,N���'��y��o^�ʠ��u��9&�p��'s�%	'
�0���*͂#l�M��O�}n�i�"@�)�	����Uz��'6J��q�K��'�~	ac��a��֟`����ܛ�ߟl�<��$bJ|����'{���s�BT�l.�iF{�̈́�����=�V�c����% � �8�ɉkH��I~�O�����9`
�����Jg4���'�$��a	�:���KW4�S�Bh�	�6K xs��)��)���f��I�͈g�i%��'�S2֚��I� pH����Ը��� Z�\p�����M�'g�(��X͟R�T>	�|���Q���`l�W�ҡ1R'W��?!gH�V��Yz�(P����T#t�O�2�����J��pRt�	ǪѰ'�'"����ɧ��2��h��a�aySO��X�b�Гe0D��ل$�kiB�{��Y*Ox����M.���?%�RU P��6�$H��J���M����?�A�x�����<�I埔�	��u���5��3Afh�0Dܩ TĔ����t1+�+,@��{��*�Q� :�b"e�(�#A^�~4�iq5G�.��S�̖<�05�$Ŝ�e<˧i�����yR��6��Т�C�~ܘăF��򤋫[�g0LO�`������[��!A"Obœt�.�M���Q� y�9�imp"=�'�䓗?DL˕P��4�S(�=�5�3�
-�lhi���?����?Q�\?9�	ߟ�!Q�[6]5vs4@�<J���*�+�D0�Za�K1p�܂h/ �D;7�	7�T��bڵ>��Ѡ�*nԪ���f��\zR8�#�Z�>��5�w*ԷEF���!A/�N�$������O��xW,Ϧs������ abA��u���l��ė'Xt��Vy�^���I���:�b�(��`�"����Dx��?Q�g2�韨�)�O��'^�@�����3_��lą( �@�e�i��s�H��)?���%�M;��?�����A��[�H�H�@���5������N���I��X�T�ϧˆE+���-w�|� �Q�^��m�r�,y��o�89D<pC%��hO����"P�r�4Iƣ��(/x����躃� �鉷/�O��`��ǻaN��hpчh�J�i�|R(��?Iq�i�X6��O&�0*ސ��BA�6�yă-0,B6��O���?�$�OV�d�Or�o�0G<
0�u12��F= �Ӓ�x��i�b�|b�'}��' s%�4 Rc��-)M3�-#0X��J����M���?�����ѯW*�?Y�x��G�*a\��hW.S�J�e�7�i���v�+&� �k�'��^>����$TU0��a�'��q ����ԆR
����%bzQ�0�X爟`T� n֓2�u�c��>I��I;��Od51�'�x7��Yy����f�;�h����2"��� 	�>1����?���O�<y���Z�R��u�a�ߞ\A`\����xlZ~�I�?}ˤ)K:'mf�P�+Z&,)�,U��M���?��l�L����?��?�b����d��VmM1��%Ø�pP�Զ�+p� �ě�(�@)3��5��(��n�@�& �������[:<ʓc嶜s�$2��}��F�IV+̀4�i���:D,�'�T�,OV�%���̟0��4��!(�?=���E�.I'8�m���|��џ��	'N���S���	/"m��ӷ|��5ʓ'N�1��!c��W�vЊ�49���]yR+�~b���ȑ)��� )Ev]��M߮@I�yB%�
���Of���O����?	�����l�h�8'��3;՘dၐ,b��e	L�îm��D]�ay�����I�K��ڵK��w�3e
t�ni2 ��9=ޜ1�̼s���ʚ}�'���p��W�n,BP����u��E��(	���i���8��qYćs0&D����-k�p:�#D�����I�a�6���̏'3Ґ
te�>�A�i��V��Sr̕��M+��?��OȪ�a"H�i�0,���ֈ,LFܙߴ&��}:���?��3�N�H�H֯�HA!C�ַ>�\q����������%. ��j��XU�`��	*J����%����SJ��g�3SQ���V�(1�lL�A�+T?r�3��2�w�pD�����P�Z���.3+�Q�G'�(K!�"O.���
�%R�E�J��p�G�'�:�r��qp�T���`�4'6���'��H��$~ӂ�d�OJ˧85�1 ���?1ġ�0�r\(���<�f���
;�����=�4�ؒޤ\�2�S���IV�A)���M^De����w0��d��^P��bC�JyA�KuL|a�P	)�3���Eύ[u��ڗ�.K�����*Z��dLj�)� ۾}ZC�!�2Em��Q2��:�'K�}Q�E�pE�j
�H�����$ @�O^����fȲ�;�ǍA���N{�����OV��q������D�OP�d�O ����?��j�����Ʌx�:�����&$��'P<1���RDˑ�j��TzBm͏^�(��)�<�ol8�$�fJ�f���A	<=W�E� �ryf��?�"�'�	��O3��T�j�'p�Z���'���4ᗨ=��p��$p>,��ܴ_e����h�	-^�t⟍[8�����цS安cA�1>K���I�D�����\w7��'1���u��-��%ڇDװ�J-��[���AF����ū/�JI0�D5��.�⥘1�ߵ$
���6AF<�[FO��}U��b�*G�)jGC���O�Y���'רP�r�ߜ,<�z��{��Z�r��d%��g��MC�I�G�Y����n6X�y�!�c�<�T�Л:�(5�`�@	s�h!'\\}�Ff���<���Y<73���'J"ڟ��$
�}�����c�R!�s�i�ΰ1�'�b�'`��r������O�	H�^�����n��)����zQўXx�"۵Ye���6��"E$j��`�ӏ2�];Ц�z�t�c��4Z]Rh� �W[�'j���`>9��N�e���Y�ḽ�2X�F�(D��:WA*=5Z���j�Ve6!�3-%�O4��'ÆAp7�ׇt��&oS�F�B$��ObL���X��]�	�H�O�:��d�'��3��)�KQ�R|բb��}L6m@ )��d*�|�>�G��7`��q�����)dj�ß$A��:�S�O&]�L C9�eXU1U�F"�� �?Y��|���Y_�2��B�]("U��/h-� �'�ѲtE�A<��,ȧi�J���h�O�,a�G��?)Bmx3�ң��L�t�j�Z���Od�
�ϯ���$�O��D�O�|�;�?��^1��#K
�Q�ȁ����]q��a��f��_9{v�y�T��L��	X�E�2a$�S�+˝u:��i�Θ�\")��@+�l���^�U��$�:4��'L	�R�'3�$κ#@�� S���KC�T�ɪOi�$�O��(��y�B���D`z�k��M�!���#1.�P�<9Ɵ.b�����FA4��a������4����<��)�Y-����dÜU���h h�,QR�I�L�9�?����?���v��S��	("�0�d.��X��@�1[���`L�"{$D�X'�>8E�]�6�\��OJ1օP)��9��C G����@;4ZU#���Jy�qdNB�~=Ĵ�c�[�;��8�{�ڝ�?�� �=H`�\�����%��|��G	ۃ_s���'P�I1�u�X�|���^wd�Q�ӕs����7��1Mj�+M<����?ɠ%\�<YJ>9�O����!��Z��V��`���r�����Ҧ��Iiy���O����?Y��k��C&	��&޷_kD�WJ��P�gC����🨒& U��ӓiB����P/�0
�dHQ\8�!�����}J^x�So�*�hO��+'�S��s�m['20�S�-��c��*n�	!����uBp�j0�R9ix� 2�Av!M>��G��� �4�1��H"�n�Y�>x�A�^(�KaU���	M8��{�@0'��Mɧ���4�
D��@'��4��|ꢟ��{� �.'�챘��Sgaڅp ȥ>e��=CB8
�*�Wnd=X�f�C�'�r'n��c�<����$�`��
�'J}�㉞�#z�)(��<Yt�,x�'8�C)�F"�L�Ɖ]r8�
�'I �@d��<���0�*�7�J$��'�����xv��ah�!9h�
�'JHy
�K �+���R�3.؍�
�'Fͳ�ዲ,:�Й%.#��K
�'��
tO�axflq�G:Qx2��
�'\����Mh�}P�e؅ Ǥ���'���BGm��Y2��otl��'(�5Q#�H�1���X��8X掩b�'l��`GL�-���@�P9DV,X��'��k�E.;j�HJ�K�J�\K�'� ��C�ܕF$�|h3��;8&i9�'�^q3.�d�����N[C*��'s����`�x)�i�}l�պ�'Ќ!癪�0�a�d[�L-����'v��FˎdX�)�,�x*���'m�-ɗ��,�)QP�Q�uM6�H�'�"ܑ��K0m�cbM!`V�q;� �=��'��>�	�l��b ���a��Q���.&k�C�+s�f,�������Aaة|�Ҹ2e�"?��3�9�������:!�44۳�@�%a�P���aa45ٷ�P�e�Ks�Ш���4|H�I
���S�mI�7D����-W�pe�E����ypA1��(O��{tI��=\r"~R��V�e��|`��Y�j�ʔ��a�X�<��"*�B�[c�^7� �WI�7o��@U$��u�R@0�y�}&�DU@�8L����Ш�H!-+��($��=*аbҬйc>>`��
�zG��ۧ
fM
�9��F؞$����c���h�F� a4: &�6Ola�W�u����q7�n�=,"4�Hw�Nn���c�#�NC�I�?�
�#�i�D�y�P�$\�pR�h���$�2�J�oI�h�Ƞcw	��k׀�F�ܩ<Y�9I`"O�	�p�Ƽ$���c6I�<���w�Nwl�I�'D���k��=��ϸ'X�Y����G)���sbǓY��̃
�h؆X�bD5:�����
�Lc��DP7�@U�W&� N�A��h�J!w�W|cP8zᏐ� �̢?)�̱���C���6�' Զ��Q,��VH�8qƼȅȓ0���tI�;t�����3o��'Xj��UJ��ZO�@�'E�0\Є�Ӏ>T��R'.^8ڕƶn C䉕-�n=ÇG�M^B1S���*D5�X�F�Ƴq�x��-%9,�@PK>�)$扤|U4��@-&c��1�Cľf��C���<�4�X`�U�p�� �DS�Ҥ�2��E�Z�	�g���2��'������6Q
�ՅJ!��\�	�n����V�H�n�
�b��B-/|V	�H@�K}��v̀�nh�$�I�<��١C �����_����ώY�D�z?d1�ˏ=s7� 9p 1�'^��А��^�˂�iB�2w0h�ȓMh��ou�a��o�X�Ԍ.{�q�U�'��(�Q�g�.[����)
F�F����ۋcV�C��p�	�h�H��#�2}�����送H��ы�d����YF�1�ց�Y�z���;LOe��ǌ,����5O�,Aa��Y���I�W��$�!Q"OZm�e�)U��
2-����Ӂ��M"5~��B�b�{̩�4�]�I�X%Q��D�6���дp܊C@ةs�8���̿�yR��K瘰��=6vP�jƂSu~P�p�+��x�ag�0��,9S��k����t2�� ���CGT25צ�q7��jx" �"Oz��@�y�b%���H.  �y��_�a�����/~��� LO2�O����س�5<C�5h��P�H��f"�O(���g�
;P�y��d�h����J(#{j��������Ad���.���	$@a��ԠP5,f<�hՅ\��>bI	nM��P�f�3��]�wl��-H���#�wƔ%��$�Tl�f�<Ѳ��*l����F)V3�P(��\?�BM'j��F�7�fh��g榣|�����m�@�c��
�:�M�a�W�<qF���/d���F�pFl�[��JG�
��@�Ǝ�M�ʀT��TI?9��{R�
�IK��Q$��u~���kқ�p?��bI9Ȧ	`�(X�p%Y{���Ut�h"ˀF��
U���'	\lQG�'���c��X(>;%	���[�����@+v
��Y�0kJ�A������J�=O��t�oC
y�E�G�X�|6!�Ğ�~��+��X0����Ā(4��)͒���AdK_�bC���I+2H��K�c�v%B�KC(p�!�
�8&��S�O0YzС����Y� ��aƅ��z6M*4��28�H>�ɩFq��^E�]��XyV��^�5��f+9X��3A�ߪ<��ŋ�&=b�B���(3$~��Q-Tl��\��F%��)���?o��1�^X�Pp��QaY���+9�]oڍc�l�2�;`�tc$�7K����ȓ6�yC��<���y����u[&Y�j�f�aubǣ�d��0�Z�)�z�l:ʧn�
š�a/��s��F�>na��$j�"���w�P�B��U9�8A ��=R��zݴv�4� c���S$��'u�y��D�d�.�Y���;��9���]N6ո�e#4�= �eW���l�׊��J��1@'�R����6X��z�_)XKd�b��_�ȓU����Op���@N ��)����,y��p��i�Q�//�j�K�� f ��"ON�dW�n����#ќ_�by�@�O
t�E�>�f�s��2gL����(�vآ.ڍH���BØ%}�Ȝ��"Oha�Ȓ{���G̾� �{���.ɬy��q�`��u&4T/0�O�r���p��x��P�僨G|dda0�'L�$���  Tei�0Mā��� ��D�q֖< �@H8������l��I�h\�5�r�)&~
Q�L�Â��FXq(X1W��a㥄i��Lh�G��*�8ؚ!��!,����)3D��h�l+{��@U�O� �A����١K�=j�1�Wz��4k��}�Q>���́)���L	?B �;D���&	�&t*��JE6���#D-D����J���Câ��
C�,D�X�˃)���Ӷ ^�6����-D���ˑ	Q�)a�X����/�Ov�1�������%96��cEZ��ل�"D��� ��JH �y` �;%�i�=�M����CI�k�O�`��W
�>�� E  z::Yz�'� %�R�VQ����� FĶ8/� $�V�$��'Ƒ>�@qnU��L�1/���iv�ϕ:g<Y�� 
������T�h�(מ]nZ���d	���0>�1���W���ȃ�`��WK�a�� j��!=����!�O��9�-)b���DȩO����"O@5���:X�*`���v���S��H�?��(	��h�O|��	��#��P�䛠l��P�'��\K�f.����:���J�$�a1����La ��I��(��	6=L�$���u*8�!�̋i��C�)?ь�"b�6ȫ���Y0���	b�l�be+p���2�1,Ot��ɌO�� "0�*06�1��'�! 4�8j�6�3�lP�xʥ�i"jkD���֛k��1��L��PxrN���"P
HzX@˛��p<�"���w�ADʈ�J ��4&Ī_@Vd�sf̓�VX��Ê��y�k�oZ��8GS$[�Pwh.r>&q��mͭ3�4D`�mP
5�� ����>9D��_]�A�Fm��Wo�QH<!��A!u6�U�ԃ9��9��[�@Uo�UN<��ǉ@��1�	����z1c:���J�)`����64�T<�兰@� �����ږ#M�d/ �+�aV�N�`�Q��M(<9����.���!�QSj���`��\�I=���d�ܼ3ȸ���
/]�����/($ ���Z2 �|	��"O� Jt��/?|�
I�pO�(����T_~���Ӡ�Mw�y���B�	���k �2��0|u�1I3��O��Ɇ�?d���P+p���m� �b��Q6}_��
�
��)Z���1��qUb�1� Y3���'�����8$ ���p�ĳ0�L�3� _�}'N`�'V�u�B5��iT�DU��'^��JK�t"�)shR�j0���>�P�
,-��qzuj �(�܈�s膂4�p�qF�G�+�^���"O�pr���$ep�Q��6��inGlx�JV���X����� 0k�́��]�0�U����8pN!��S���eG	�<�0�mN�{E��[�vU��#|O`�BW5|:~�;Ҡ� �S��'~�@:��O�Y��V�~�P��K9`��E"O\<[Qo]`��q��I&r��4"O4[��V"h��1��b(,�;"O��1�Û2D ��� BЊ�"O@H�ƍ��1�
���\�("�#�"O��"PiT&W��<��bE�0h�;"OP��N�?JgTa���u�Q "O~qZE�\�x{UG�?x��@"OHI��j�	E��-;V��8��"O � �j�<�
d��c]B���"O>����ؘ+�FdQ���	��sb"OJ��TA֜5�H��$ԙA8���"O�a#���45nP[��A�/�-�R"O�<x���60W���a�V�n�X��"O\��q��ZBܫG	Z�JZ�r�"O�"5)B(%'���v��^̛�"OHj�zn�y YFL�CG]��yl�6p����΂5l���2!��y�Ü")�0Ը�HP c}�3�K�yR捛d4��AQ���L!��	�'�$����l���A&�["��}B
�'-|\����4�x�@Ph�# ��u��'�xiz2-��`�L����4:zvD��'�J@�dc��w�J��t�L/�d	�'�r�����!O� ����#����'$�yc/�mA=��T��1��'�tLH�l 	{��l�V�ҁ����'�d5"��.&x�摻SN!��'$��!�׶|����e\�q��'��	S���$E!@"  Wnl �'f�pfB�;�܅�E�D�v���'mF�!U�-���sD-w$R�	�'�d3CN:�<	自M�`��<
�'&��zM,|R�JG�կ-����'J i��.��YU�xj��ߥ#�H���'��Y���"�2鐄�K"\ ��'�,$�2��y���g�+Z���9�'_�h�TVs�F��K)?����	�'$l�b�Ė�={F��<"��U�	�'��)�%�°5R�$XӁ݈�B���'�V���*���u���#,*&U��'�r|*�';$q�զSb4��'���q�ߗ`��){2�ǰI�L�z�'�Ys'�U�=r�Q#���*��' D��1p ��7��'aHH���'���@�b���w�>��p�'�&m��A�d2J�q����Lt�'�9
�m�M	�q��ՁFn�t�	�'V��+J	yp|4N\�T�'�Z�05��>� ��ע��R���'�R5��j !{4\2�J!��QH�'�y�+�0�`�9��ݥ ���J�'=H�`eC��{0>�U��jj���� 4� ֌�/0ZY{�Ij�e:�"O$��U�ܦu�P� R�*\^���"O �(#�G�J�L�P3잹Kv�"O<s�MB|��<z��^�c!� �"OZ�g!ΙDV��BbG�i�
�1"OJa15t�B� �'�>.��(S�"O8�M=0FyS�G�	�F��"O�=��(�6-���S�L�31"Q�"O��jV&ڞ{ւ��q�(.�%�3"O�G��?�D��"H�jrm""O�<#�N�vbdR� y$��!'D����A�%�l�6IU�JD�c�*D�j�W)�r9 ��Ҩe�J�r��>��	 ��-JT��@��b��X�'-�mb5	��."���fז0�ح��'-�Iy�L��]>�R�!�~a�
�'�� ����G�u�."6� �P
�':���a�
@�ؔ�.ڏ<f�M��'؜ݢQ�-Զ=�p�"$�r�b�'�n�r���|.8�G��h�h`{
�'���""$֙;�ʚ!\P�0�'��hK�h�&c���:�B��b��'O �����M�T���(�04Ƕi��'5�a��ďp;�Aϲ&��Uj�'�0��	J+^�b��BU�L.�-Y�'��y9��_.(��j4LGK.��:�']f�yd���p��AcN�L��Ik
�'�"�ѩQ`*�z2�ԼX��c
�'�T��B؉;�	�a�;G@>�`
�'��� gC�)��$�	�BZT�
�'^,�i�X��v��@� 2m ��'ĺ$b'
F3cIXd���C 0��K�'0���d��@�pM˳I�/(�P��'a1��H��q�©C�%Fb�8
�'k����b=̑Ca�=^��	�'�^�&�U )p|�7�&�B
�'�:����	9G�1ѱ�Ů/a�q`�'��Ȫ1��:�pQ�q+'�����'q p@W� �\�D0rF���,�@�'ײ+&� 1 ���1�I�
v��'W��I���Z8�q÷�[#��@��'�qQ��-u���צ��O�(9��'b��C�@MT�)�wI�KO TC�'Q��X�"�F-
�&��@�|���'gL��wN(+���0�ň-}�$�'�Y�F��@��U%,��mJ�'����E�J�Zi��
��
�'̨b�Ħ���)SQ�[
� �'�)��,{�E�E+��L��R
�'�Ā"c(ͳlF0�`[�D�t���'�ބc�ô�@*U*K�;풐#�'~qh��x�v\���9;3���'�䢠��RF(��c͔b���c�'�@ �uM���H83�A�a�ء�'Nd�k3`Z�t�p���N�_.���'I&؋������Ǒ�?���
�'NLa �F�g6���c�?i�@�'�2��U
A�6��c���	��}�
�'�t�yT�_�a>K�� ���	
�'��������1�5�I.}���J	�'E��F��Ms��×E̒n��1"�'�<}�����V��@"b�n%`�'ը0s �ȡu�]#,D`� -��' � ƪKo�E2�\9e+x@��'J�|3�������K1V5���
��� ̡�t� Fӌ-��Ɔ��"O�<KuG�5k���JŀĎH�Ȳ"O �7(��zT:e QR8��%"O`��@��4�R��9�/X1�y�W
bU���%�Yv�$�흏�yɅl\fL���H6b(��2�=�y���4&~"p��s.�,(�霛�yb�E8����#N�f�r�Sd���yB�D�F�� w	�&-=���!��y�h܍z��� %
��j�X$�@&�y2b��Ps����E�mE�LV��y�HϻE�Ft�����N�Y��]��yҏ̖<�
�Sb'�1�(�t�J-�yB�?_ ̘�-F�6�������yR���R�f�3�oZ��3�Z�y��th�9�k�) T�)qH��y��.:I�E��cˍ{�q�W��y���=&�, a�aR��C]qhB��$J�,d��`��\"R�	��Y�C�ɥjR�����H�)�ݮ ÆC�	<B$�����8{�֔Q���$y�HC䉪8`��Ab(��kX� �%��+ND�$@B��h�E��'Lih���(I�Q��D�AA2�O��O�S`iH�e�ڈ�cËK[����"O4m���9,���3@O�[��*�"OHhàl� zw�����G;`0�c"Oؔ���I%k�� T�_G��A"Ox�U�J;b��Q�%� �m��-��"O0��ၔ�B'��b'� �h��0�"O���gM�|���M��5�
lQq"O��3��T�M3ڝN�-&�J���"O��(E�.����G� *� "O��"''D:�4)��3S�<(�"O�A[��\�2���rE��"D�zuȔ"O������֐��+��#�����"OHaфᅪ$V�����
L����7"O<D0w�L;2Z j��c�R��yb),�А�2 ��"fZ�rG'�y"N�-y#�5adJ�$r�+��^��y�a�g�ĝ�J���H�؀����y�횊FTz����\�2Q�˰�y�.�"GJp��wd�z�L��y���9��1�$ɟ�hcޱ�2��y�N�I��.C,0lT�aɕ%�y"��"e9 ��q@2<Vpk1�_!�y�+g���Qv�H�0r�h��ݭ�yr@{(�m�VI��'�� �\�y��Y=fl��Nتt�R��^�<	�O�8�*"��8_���xgB\Q�<��.ށ�A`G�z�\=�A&�R�<�s��8�5����&�Z��#˖O�<I��X�[�H�������)��VH�<�c�<+^�<#R�9S01�3�|�<!㯑,j���G�I*M.��$�N�<9q�T8X�*�RJT�K��D�B�<����	iNXVG 3��؇�@�<�"�\s�Ő�X�pJ\�ڄHz�<��ͺ��C1 ���G��{�<	� ��z�� HCdF�d1ʵ���O�<	�;"��rro�j~BIZ��H�<QV�ެJ�H�q2A�H
�K��Z�<�1�2�s��vS��r,CX�<1��V�ĽSE����S��M�<A���&�2���>yh��c(�`�<� ��y�W�,FxKG��9Y丹s�'���<�@�A#&Ԓ��١c��5���\�<��❈2�I��Y�@��y� ��Sܓ��<%?YQ֦/T_���!L�0U:���j,D�̐2��+������qf����8ʓ7�h��dΓ��� D�1�aF�\{!�Vp���,$Q����%Rd*I�O�=�v�#Z�`Q�R�[q*E�'��b�$;R/�S����f �]M\ز3�!D�0;��ѽL�0��#�8�Lp��l �ɴ'�Q��bL���e@~t�4Iň&�)�!"O�aPo��V�z1x����퀳A!ʓ�>�(rص�t�N�	�*�Q�Ap�4a�ȓa32q��.O��T@G��>}�xUlZ{(<����#H0j5�r�ʥ� ×C�<Q��R�"12L� D�,��DI�<��jV.RH*&�V��V�����M�<�qmH�hc���7ŜJ�tP�桗I�<y�	��-���\�F�4)q���E�<�%#:���Q�q[�Dc'A�<�6�V�@�h������0dE�<�K��=��$Rdٿ�\���X�<�l�$�mH��7k��j��QZ�<�gC]�:`6�r�D)!.����O�<�#�A'l���pF@��V��� �F��<�í��٪�g��Y����b��z�<����iXE˂h����!�%(�s�<�!�׳tzm���˨4��H�0�Gp�<yC�6�f%)H-,GT�@Nm�<Q1'W��AA��(G����q�<�ǚ�a�07��Pܵ�TK�k�<��˕d�0t�'j�[ )0�d�<��'�Y���ڃ�ILdf�8PE]�<�JX�"�RT��$@�rq��*��GU�<qf�^�{C��R�o^�X��B�I�<Q��<t>���Ղ_��M�+��Ї�d\�|��^%8�ģ �pD�D�ȓ|4j}��fX,��lR �"Of5��,
fB��� �Dld�P"O�!�S�=N�t`��h�~Pt�Q"O~��aKM"&<�w�ֿkO��Q�"O�tcpƔI���b��̺7=})"O
���� #i��2v�F z��e"O�����b��mJ�M�����"On��@��U��� $H�2��z�"O���'��#��W�,s�"O�ň󆊈52,s����p���3�"O�"�C��*�+r���a� -�e"O�]���Ve�ؕ�!�M;C�U�#"O(4�NA<�ji�tm�(lP����"O`����Qx�л�����=8F"O�e�q�C�4�$(#�ED��B�2�"O�(�c�ѹ.*x���s�x�A�"Or�(ת�g|����ؔ�M�"O6i
��<
�8T�"��-Ո �"O�d���e(�cw*^7O2�s "O�8���i��곂/Chl[�"O��j�����蕣g��)��"O �r��Ȉ��D����=�fmq"OA���
T�PB�`�
f�����"O`  W�©o��`�f`��H����&"O�a�0kǠd�[���G\��"O*�هOO�n[�e*��U���%"O"���'߭��U2b�ˇe����"O� ~�Jw�L�K�"٩& G 
MU�T"O��gA� %l�J6��;H��P "O�����F�R
fa�0/�!ZH��i�"OjTk4"���*�k%���)*�Ad"O0� 䙭_�Ra�2�U82�d�: "O�9*&�Ȫ+�n] &�� TT��1"O\ۗ�@�*�"�h����y�G"O�l�6#یI���ht-�Q�j QG"O
$�Dg�Gs!�RlԷn&���"O@	�@h�\�xAҀ���)r"OƜ�e��:q�гe�1w��9�"O|Tӗ�N�
��W\l�)�1��E�<!׀��q�])�G��4̙%�T\�<16
Ϗ<�4��m����`i��<YUEVP� !��|��OS�<!`¢G0�[�EZ�CK���R��M�<ɡ,� Q"��� Z�hQ�w�G�<�%��   �      Ĵ���	��Z �I�Z���C���NNT�D��e�2Tx��ƕ	#��4"�V�����8H��m�H�uX�Օx]�LV����E���XX���	��MS��2
����+�hЯ;X:vݛ��'��"�cěP_������T����vH�!di�%ay�Ϯs�V�Z�%4}��HE���BK(h��v����B��(��:��M�'!t���)Ͳ\5��r/O,��`B!�t�a�X�D��-�
dB�T�Q}<��AM�sd�l�'�9_��ɪu�PP�d��r��S4׺,H"�V�Oanܘ�A ��q���-�ni�O��x`��5YlOR�cF��&*�StV ��mO4��Ě�)�iK��I%1l��Wb�}�	�mi��æx⓽:�b}�T�� HB�P�䗻���'9 �)b�0}�%��lFu�L>i`GL )l�='+���Hc$�P |��:��q�I�'�t�eE#�Ě'q:vd�e�O���3mǈ�C&'j�N�"�I�T	t�#fn>�O����	�hs�'b U��o�*E.QX����y������y�����%�HybAB�O��S��ʑY#���w��m�Ǡ=T/xq%�R� {������%dX�=������'�¥M��O�q �$A�����爆TZ�,Q"�]�,fj���`ƀB�dو�'� �ɽe�9�UV��ө���c@�E44���T}�2�jN9
i�'� ���%޿��5!v����<��	� �pQ3�ɺ&�bE� syR�@'�d�DyB@�r��IX��iG�#z�.	�Ő\"P���8��H��xr��?y��t"ժQl?��à,��4��,S����X��3oH3�N�c�l�3���]7Pw��[B�7������lY|��!↱z	�4�`hB�m 剙*� ��R�!�$Z7��Ҙx��٧W���"���?}��i��H�u�J���
�.��SF��R
�h��5v"˱Y�\�v�I�a�򅙁fU�cD�C�ɦ.:�  �'<�c�dG�1�5XU�ϺAbƙ�Ó�hO�8y �M9*�+1)]��F�"OP��K�s����%�O�i�5Oޜ0,1�)�dS��co����x��FߌT����ȓmH���EO�yT�)r�	{c4�'��#�q�ݪ&��`I���l:;]����l������)]�v�z�����(�CuK�J������ȓ.	`x(���Q�
xZ�E� Q���^d6��   5  �  i     r+  p7  �B  �L  �W  b  
m  w  M  �  ֕  �  آ  I�  ��  ͵  �  U�  ��  ��  �  ]�  ��  ��  #�  f�  ��  � C � u �, q4 �C �Q �Z Ka �g �m �n  İ���	����Zv)C�'ll\�0BL[H<yVCQ��F��e�P(������C�<��	��e��A��+O��$���X@�<�v�C��p�TJ��izsf�a�<�&	�P����w�&H�ؐ���e�<�0i�������^z��B�V�<��(��Fz,Q��!\:�\U�N�R�<yӅ�I~��3��,}��٣�JVy�<a㇊)nt��;G�ʏ���b��Kv�<i�B�r�8��L	�W6�}�=T��zf���R]��0/�6őf?D�haV���  ʔ ݿ���1D��[�
(m����@!\	{�� 7�.D��`ƭ�}`|��a˚t���Q3)-D�[2�ߌ=�v!����ɳ� 8D�t���O�u|D�Z��Y�P�1c��7D�LÐmֱlGfPb��U̮L,�0C�I�[mH=�W�٠d��C�l�&9�dC�IMM^� a!1�>�Ie�?`'�B�	5Jy�]��tn`���JF}��B�	�v�6��V�+#*t�c2H�`��B�ɦr9\�{��*v�h��⡍��vC�I�v��ɐ�ƙ$�P(˅��=EItC�I��9��ǟ l�����&2lC�IO��P��(����'�lZ@C�I�aS����k��p,rI�3%�`B䉅%���Gk�S�X�z'.�#�C䉙U���@
��K�V�j6.����B�I6\�qi��-d@��4�\�Y�B�|�d���a϶l	Ҭ����_��C䉈-�I�����NL�,�ب�E�8D�l�C�*&�n�h��Ώh�YS�j!D�h�$�$!��0*$�b�p��� D��3�X(q~T�אFbv��K!D�ȩrMY>n��ڵ��$V�$�P�5D�l;'N��d�MJ�6[EHS�%D�����£j|)��f�}�� �L?D�,q�
ۨP>&@���S�b��K� !D��`��F�h[�D�!�Y��dZ� D��i��J���ˌ x�i"B 9}R�)��*4	
p�׳[���0��4GV�C�I�b@t݊/T&#�V裂iG/E�NC�<�T;�%�D�>,�D�5{C�	%l��,٦ ���� a��M�C䉟wƜ@�G�ǚ;�,+�C�J%<C��J�1�P��P�J,	��B�;C�%����r)՝���LnبC䉆`�t�;���0�:!��
�H��C䉨c>�ّdeVC!S���0ѬO����_ ^J��6��Op����
�lab��
���&L������-C�f"��"O\{e���9����g�z\H��'V�ȁ�M0��ÄA`�A�� *4B�	5X&��ٕpP�����
�z��'��⟠@*�b�nӘTp0E �l�H��_�~�Ʉ�qPLQ���:s�T�pv���YĤ��?�w�'6��1W
;dd,QQ�>wt��'�8�m(z����c��[_`X��!;4�L[�� V|��#/�5ۚ���vӾc�\�S�gy��ȴ/B�jgbD�wޢ��2����y���{��ea�h�|���r�)B�J��#=����k.�P��gޡW��y:��Fnaz�Ы��')�Gf�ZN<	�E��;*���p�'rֈڑG�/3�&P�+Һ#��=�y�EB���π `a� !B�a��	�(�-3��'*OTM�l]�Jz"�4b�!ȴP�'mH�a$n {\i
��)fe~��'�d1�T�x�A����I�jT��->$�`S3��<�+�"���@:\O���<��'Ť̳��H6|��1�ƫˀ3hx�	�'μ�¢��Q:��{�e�2-� u+���Oz=E��J�01ꭉ�J@�S��1�!a��y�I��l��gH�Ic�yQ@���x��'�2�#R�	���pg@T�[�'~A�_�p�ቃ�.:��(9��hO�-�E�$)�,�ZlL�W͌9 ��'g1O�-�7L;7��Hy��K���ɷ��dF{���ɈL��yQ*�.I���0j[��{����g�"��$��\�@���96�����ɬ),J �tǀ�M����
+b,n�=�ÓM@2Ȱ7X5�rl{��7 P��3J7�ty�A]oG��t/8�V`@&d8LO��d=�D��Oj���	
��n���C@�	Ia~B�l����_����c�"�2	��Ρ�!���"}l����n�rp���
�!��S�68R%�/e�@����'nۛ��)����
\%;�D$+��S(y��c��:}2�)��16�v�+���dtL1�pD�(x��C�I)�Jh��J��y
0����c���	�Qj����	/Y��e�$o���C���Da���de�i�Q�?C�mUd.D�P���
����o{�x p�(D����ݹk[�<$���e����rG'D��өX
���	��	Ͷ`*�,"D��� �E�s�	��ȃ�l�#3D�,#���\���Ԯư\��p@
2D���4��[.ԙu�����(A��0D�� v��! ,7�ޠIfvl��L�Vh<��+yf���cлcPD"��\����?ya慻O���A2鞸6�0����R�<)¤�m90�xe�˝ѐ+Fl�զ�l�G���>E��4E:���d�G�­� �B+(�܄ȓ8�.��W��z�rq1��%h�=�ȓ~�}�@J�;ufu
�Ǡ4��M�ȓ.T
M!w�̋f���psD&L�ȓE�f�*Q�T�P֢���Ĝ*H���!6�	��4�`�0ѫ�>*�}��c��,�c��<������T��l�ȓ*�f��o��y��*G��6%�܇ȓ/��``BJ��J�h�lүy+ ��ȓ���	� Q�a�����jG�sY$�����)�dL1�l��ʄ���%��0�5�dj�;|=�Y�G%l!x�ȓo��,q늌'���T�'+�L���W��Q¢�1�X<�ĥ@�YW|���2Pa��cG�=)b}լY$x�Nч�w�<��eY?z8D�!�%��M��8�ȓ[��B�펭	�NxI�A7s����p�X�"��_: �n�@�K�N����q9`�2,ޞ��B�սmty�ȓ��XnK%�Uh%��0Y���ȓC�x������*�2��(���0D�82��k���*�o$K��%�T�.D��*"��a�X2��Ē}����%lg��7<�S�O\P ���	xL�*���^�jٱ	�'��y�Q,DOw�uYt�XK-��C��?�C�'��X�� N|�H�+�>6�B���Ob�?	�O�P�9���=Ca��c�.#����� �ӗ� 砍A�ߐUCĽ*"O�Ȉ�oԅ6�Ꜣ3�Z�|�p�:�"OƄ������HY�a��;����"O����@��u���Y@��ifH8��
O�6�J:΄�23HQ�Yh䜀��f��	{x����-�!"ނy�A狌$s�`d�4�O�O�p�B�Ґ ��9��Ի^َ����'�!�d����řEʅ�K��4��,�^L�Im��H�x�kd��%H��c�,p��i�""OD-2V��Y7k�za�%JW��'��hO�OT<��&K�M~�Ѭ�DҬh
�'DI�A	;H{�p��3�d4D�8�� ��s����(�~����(4D���5N+� �C
W8V���E�?D�0����z  �c�j���z�j�O�7�;�S�O~C����	��x1C� =v�^숓"Onmd��ߜ��a"��	�
1�S�h�	P���Oن���I�;h\��M*]�8�q	�'�v0���⏷|$�h���J�<a�.�0L����fN\�����Hܓ�hO�O�`�'VH��u�*[��:,��'2��b/�0Xfe«ݣ]�¼z�'o�'��<D�DX?!@�Ӷf�,���ľ�$�f�!�OP�Q<�qP��CkjH��J��2˓x�ў"|ڰ�_�|p�j��q��	���{���<!��� ��1P"�D1Xf���aI�y�<�E�1�$81A(I��	 vc�\�<AU�޿GڲyxĪ��"�����GY�<y�LX5K^�I³F��2Z����؟̖'@ɧ���[�%̱0��xH�����հlX!���4OK��P��ѼM�Vey7���vC!�DI%X��Mb�iL/.�h!�D�!J!!򄜆&9��9��-���-�!��$LJjI��l�&r�}�(˵~�!��\�2F�x���?j�IB-��9Q!��b�M9��޹:g�yj���ZP!�Dڶ=�68P��xVL`��L�`A!�D���$Q'qP��EX1!�$�hi
���X^���@�Q�+0!�d_5$�څ�DF[&�xQ�`�/!�$�-|Nx��6�cI�@�@ 6!�$��(��a�af�.<������@!�$�5`uqR�{��z���1!����\�$ I@�d���ȝ� _!�D7`�\T!taC�ƌ�E'.!�d��g�T�A�<����2�T�
�!�D�a0�[S�G	~и��"�!�DH�g��5{�oǙz�u�v�	�!��F3�^Ux�NK�%y�`��,ߵ8�!�?�`���E�	]��)cQ��	j����zh9ڴ��v)��s�+�,�y��y8�� jB b��������y�C<�I�ae�"Z]���[*�y��&�T	Y�� �X��Y�G˯�y�J�Grr%��� LyI)4A��y⯁�-ߠ�j�N�.B5�\z#d.�y�ō[�lfoX*3v��Šv=B�	QU�ٸt�T �P��UC�I$Q\R݉t["����.�<��B�:y�} ���P��&M�?�B�	}�du��/τ!���УD�l�|B�	���hh"��V^ ��n;ʌB䉊�(Y�1��$���$-Ýa�C�Z!p @.��-�
)i�䁭3�C�)� Hs��&E�b5�P�J��ҁ�7"O"�8�	N�H_�������d�"O�q��٩~NzH�1 ԕB֚���"O��C��B��0�Eߚ�2��"O���CJH�@v�	WI�@B�'�"�'��'��'PB�'��'�D�� �ب@l���TF�.3���w�'1��'ZR�'���'��'��'L0my�OS'|�8��ht=i�rgUʟ��I����IƟD������	�x���̓m��H�n��U��+������,�I�,��ʟD���� ����i�������cˢ9P�T��Q��	ߟ��I��	ş��	矰���4� �r��1���OUT�s��Zşp��՟�I����������(��ϟt��l֩.��	�s�-h��Mp%��ß���ӟ���ɟL�	�t����D�	�#εp�L�b�K�Dy|�Z��ɟ��I������x�	埀�I˟ �	şh�J��O��Xh� ��T�~��ԣٟ���ş���Ο�����`��۟��Iٟ$	e�Q-m����ſ�D%Aw�Oǟ��Iӟ��I������� ���0����#`�5=�U�d�x�@�sŨVퟬ�	��I����������ß������A�2�(cÞ!H,�I�U��I˟t��ܟ�������	�����0(Q)%-ZtyZ�C�unP5N�ן���������`�����h�4#�v�'��"G+��t8@�,'r��B�Mk�	����?!)O��Dئ�� O��h@=�R��ĩ����>z�ɂ�M������|�'m6휃9�*Ԉ�dK�[`ԡ�*�S�X���O��%�z���O�TԈ`�C�Rvl�i�Z�������u����X�a��,��l��<�����D=�'e+z08')��mh�ag�؊dN�LC�i�$��y��i����4cl5+do�BȪ�k�M}��@Xش��&6O��Şz�������<Qd�'t�6l��ɏ�hK.���M��<�i@�����Ę��hO�i�O�����əL4��b��@�Ta�0O����\��T���' ��#I0	����u�z(�
��UW}i���m��<��O����(�
l�E�ݛ��1�����ؖaդ7 �B@3�Ӻ2БrP�T0������ �9)Ƹ93aEy�[�<�)��<A��*Y0"�If�]�z3@���<���i�l��O$Dn|��|�3�K3%�>�Ȗ�
%ˬ�JפZ�<Q$�i�6��O�ԙ��F�/��I�ev`E*�-�z��
���z�-�f���&F�h�Ny���y2.x����\��f�F7h�i��O�Tl��Ƭ1�I�����@�'\�����=Y���-C�|��M U��s޴jɛ���O�������|X�ǅ�>^��Yy���c�-���K����-�<��$@�yPY���W4����d�	Z�R�:�'d��O��p>a2�i����v�';*��wgC A��@��r̐C��'��6m1�����d��a�۴����P�UI �"w���X6��O�2�ˤ	��yB�'��p2��Ӻi�BV����;�56�J�&�@�@���le����y2�'����D��$�5����u{�\Xt�'���'�7m����*�M�N>y��l,��e�\6)o�!13���+�R�H��45��&�OAD��၂��yb�'	P ��Q�|�"����ME" �f�O57������͋�ХxgcL�U�K�&~�ҍ�3#F0~=�ix��Q;�l��Z�^���+�e }�*Qؖ��#{P�vHҥ(*�1�+�W=��Ӕ�H�b�-jbcI��1��5WD�z��U.��XY����o�:��%e�<¡�*ϔ6.���*�+X]f-��%��<�#ϥ`�z������(ʌ�m@�i|LD��D��h}ys��~�.1 �J�q �y�cԒ=c$�oH$��z� �"�8�9����:T�֠K<w+���#L�w��C�)P3R��E��,ĉ���?�6��O����O�i]�	`�	4#I�]v�ԋU�'�N�'���I؟�2�X�	۟�	�?�b3+?Щc�/]R���/���M�/Obt���������R�������'��
���WHY�Ԩpr��ܴ�?��u<ت+O�i�O���x�� ?�<i�C�O�T��Jc��Mc��Z$,y��'��'��K/�4�R��Ԯ�:G�h�mV��b���Ҧ�j�Lay�'4��Ϙ'�d]�r����A��f�����@�F�6M�O��$�O� H�P�i>!�	Ɵ�j��0I� �����Vd}Ҕ�+����O��dB�1O����O0�D�$iش��6)P7rc*|u`+^<o�����3�M?���|"���?�-O��h�-	sR�Y��⇍-�K�L��7�O*���d�Oz�d�O�ʓ��0z�L�b��S��ڪ9�jdC��c��'p"�'�B\������v#I���s0H���=�dŵjb���������|y�F�?@�S * ��s,�Nj�!��I��(K2��?Y��?Q*O��D�OȋR>�p'=��0���E2#�%�"^�@��Ɵ��ITy�M�����
�(��կ}��1�$��d����������I����'���'�Z芉��b����M�8N��2�
=/�7-�O��$�<e���|��O7B��5���"eνz�새	�QIv ��MS,OF���O�ҧ��?7�;w"�h��v����5���R��1�n�!�M�Z?����?���O�P@V�ַ���s��96lS�i�b�'��;bS��'�&� Y�� L��h�D!]�"2l��grӢ�8w�Ӧa�	ǟ��I�?U{J<�'z�� 8 ����P���U���p�
�Rŷi�:��Q�������3�	��Pk��ݶ��0kB���JS4�y�hC��M����?��L��Q(×x�O�r�'�F�0�jãNX�$KQ�ݞD�\*��>����?Q�*D̓�?��?a�A_,D��Se��R�PD�" G�W���'��(��=�4�����O�ʓ,Dt���	�r\D�x��0^�D(��i��m���'�r�'��	�,�� 5ra�Y
�ņ�ɰ�Խ)��'[r�'�R���O�R���t�0���B)���4�%JjЍ������	ޟȗ'nb@?va�	\�v�����[.݈��3v\�F�'7��'�O��$�0.�&��`�i�����	D0?{ sQ��	��[�O��$�O�ʓ�?��C�����OL@��KA�([����k�"���i�Ǧ��I~��?�Sd2>u�$���d^W4z�c �P�A���hV�a����<)��2̊�J*�2�$�O2�	˼L�d�&/J3[�z�#�DX�8�>)�r"%k��EC�S��甕tt�Ⱗ*5�,P�S�����d�O�t��!�OD���OJ�����Ӻ+E��L�^E3QN��M��)�Wa}��'v�A�w�V�꘧�O��pv)F[0D<�Q�p�$Mk�4a9������?����?�����4����3#�-����:�6�Eg�1M*V5mZ��$�E_1O>�I�E|>�A��t��l�!��X��4�?y���?9WR���4����O.�ɐd���S �	bش�R�dߏʠ�y�/Ե,5^�����OV�	�Il��hV�!�B8��C�$e�<7��O��q��<���?����'��q�v�X�	�,up#�n���#�Or��0H?d���ܟ��@yb�'�Bh�� "YV�!�ޡJo��G	A�F�������I��<�?���8g��0G�½:�,9�Jm;���G��{�!�'�R�'9���`��~�qGP�	�,���ֈ������-�	�4�	u��?�qȉ H�!nZ�d�����'	�>��l9D듊?������O^u��A�|��]K����/? ڰ����A ��v�iV���<qa&�T�V�9SsMI�S�����X�7�O���?�AIF����OJ������[PG&E�"�("$�@J���nR`쓶�͙:g��݅9��4�e
Ǽ�r�hÉ�:(��?9�g��?���?q����.O���7�~ѢJ�0������.A��Vy��Ђ�O�OO\�S�/��QؔF?;Y��sش._ y;��?���?I�'��4�����FVq� -B�ssb���$A\��m�3#�2���1�)�'�?��E���Y�-�z�w	�O���'�R�'���X��Sğ���g?�#�0�,ЉA��!y�� Պ5�1O
%`$i�J��L��U?)ѨT�z������W���P"�Ħ��IUy�d�'HB�'<��$̹`�j�r�^�.��"�oo���f���Ӂ3?y��?�.O���
6FBll���lتD��N9@��a!��<����?i����'�bIפl��%(���$R"2��[�9#~t(��=����O(���<�~��O��]��i�B�-huʗ�?���4�?���?q���'��0���M��;���	�e*!����-h}b�'ur]���	;2)��O���]�)VpP�5&W�t<�҄���Q�"7��O�����2g��,�D�5�؁�n�����GQ>r�f�'Y��<*T�I�d�'�2�O6JI��g�0X 1!�+�D��7����ubʹ#�bb��G�ĝ��Iwƒa3�׋J�x��'M��E(z�"�'���'���Y�֝>S��A�7����`�`L�8)�r��?��₎�8��<�~ґ���@��T�Q�
�� �Jզ�*�\ş0�I��@���?���d�'b~�!�NA�\5Ҹ�k� J��h�:1;�I��H�1O>��I/K��ic��
5�勖Ǘ�3Ͳ�4�?���?q�J"��4�����Od��I�z���C�{���R/�HӶ!k�yr�*[,H�\�d�O��I�R�4U��،\xY�"��-,p<6m�OZ|�b�<����?a���'��!�d�+t:��2��$(�ɨO��Z'�+.���ٟ��Iey�'��� ���23�}�E�T,X��H�M�%	�I矘�	�d�?����(5�b᎕F�\�AȂ2��A��FW���'J��'��Iȟ����MJ҃"�:�*WÛ3>��h9 ����I�����V��?Eo��'!
]o�:"��D���"{ Y�a�H/?����?������OP�7@�|b�^K�XH�'�N��\�F�_5<�*��i���$�O�C�`ĢW��'���7�U"XopT�%�޴�:�4�?�.O���`��'�?I���B�ٲ��y)��I�����Aa�66e�O~�$��r��M��T?�Џ�2aF�h�Ȗ�>�8y��«>�����q��?����?)����#�̒>�Δ�E�٫)��x U���	2NR<�2�)<�)��
�PX[�.��p� S�S�@��6턼X����O8�$�O6���<�'�?ч���\9��C��ǳ1��Y[ ���"m���w�L��y����O4�"o��Bg�4n3ۦ�����M���?y��x�,�p��i���'e�'�ZwȂ�[����3�n%�Iނ?��;�4�?�+O"�Y�9O����������[�� ��"uo�"eR���J�M;��_>�u�i�R�'-��'���'�~
� X ����T�`��e��mV��+!�ib�?�y2�''��'#B�'�b�' ���W)� 56�ca���*.I$ymd7��O����O����l��Z�����P\3f��-D�pdce'}��tS�.d���	���������	m���4/5R7͚�uА}����G!����η\?EnZϟ����������'�h����fr���iSm�8 qԩ�p`��?����?a(Oڹ�R��G�t�'s��cd��d82��A���!*�M~���d�<a��?��h4}���)3S9R�����,rf�{Ud�E o�ß���ly��3�N�'�?�����A*
�H����6�3I�֌�թN�����L�I�H  D|�T��y�ٟ�y��ݹ!����NQ�M�D�$�i��I�L�Qܴ�?Q��?I�'V��i�]h@aϙav�[ a����+��x�*��a�Q�5OF�OV��̨#٠�ƯA�.�L,4L�z �i
\����Ӓ�$�O������'9�ɟl�T������Y3�X�a,����4P=�Yϓ�?,OT�?�I���83S���y�T��mx�%ܴ�?���?��
¼x����'���'s��u�H��YC�:G�??7Pt�A��2�M�������;bg�?�Iğ(�ɤYZ��;w�a�bء��_k�<=�ڴ�?1p�G�F�'���'g��~*�'���&���u�/'j�z�O����:O4�D�O���O��d�|��j�|�z��Qb4R����G��us6L0�i<"�'���'f���d�O�y2L�3(�Y��8C�.D%n�p�'����`��՟\�I��h���!�M��d��<\"����U`�j.v<���'-��'��'&�֟���~>W�+��))��&	���
V%NO�1mZ��P��ПX������I�wV|�ߴ�?��tJ2��򮏦s��d��W+kzR�qq�i5r�'��R���	�R�~�J�D�$s��ayb���>fm�R���?��&�'j�']"� N�7��Op���OL�ɞ02��p+���Z��8��W���5o�П��'���B�����|��Msr��\�0����ńC�-J&Y릑�IƟ�!�n�Mc��?����B���?���?+>�)SR�[%[�$2D�=��ҟ���g���%���a�	�?�4�CD�x8rf�9D]��晼�v6�O���O��i����O��.�N�Ё�E#36�ı2��M;v�lZ-���ߟ����Ē�$�'v@�x�HP�M8�eFAMJ& �A#f�p���O���T=��lZ����ٟ��	���Uc����l�~����E`җR0�7��O�˓K����S�D�'��'b�i�@�]� n2YKg�;3�%���j���D�;_��n�̟��Iٟl��'��ɸ��1����i�E��O��c��>yl]�<����?9��?a��?��� �����"^�4Q�G��T�|ɋ�M�#&/���'2�'���~,O��d��e%��"���I�4�W(I'j%>A�D��Ov���O��d�Oz������m`�\Ѿh��)��#@�5�M����?���?������O|��<��6CN�$��H�58(p�D>�M+���?q���?�GV?�!'�!�M[��?a���O1n�1�Z�k]
H����93���'%b�'������*X��d�' ��	d;nE H��3]��Q.Nm*���'�b�'1r�ˡ p6-�O��$�O�	ێbP�`a��$Z��Ą]�v7`o����'��A���4�'	�i>7�,L6�DA�~��R�	��v�'���5�,6m�O~��O��iퟴ�$L�|��앙r�V�h�G�6���'�n�9��'��i>够�!r�M�v�!�"z���;e�i��p�{�z���O^����R���O���Ol}@ -�6s�:��v��{#�͙5���	�@�GyR]��3?ͧ�?y�M@
v*\ i?�TXcŎ����'!��'��Dh#�?���O��D���F���v,���!��b�F����aӄ�O:���˓C�Sǟ�����q,ƾf�^��捯h��������M��>��1"�x��'r�|Zc��SPa�$_1�yq�]6��9�O������O���?����?�.O�� Q+Ƴi-2As�K-'?‐�HT�!��1'�����d'�������g�_.@o\X4���{��B��H�~. �	Dy��']B�'剠ߐ��Ob���$��owv�j'`�!~n���O��D�O,�O��d�Ob�0��O�Qb0CKk�X2�R:}?�|��L}2�'���'��ɒ]�~�QO|��F�<ج��e�y~�#�,��>���'��Iџ��	Ɵ�Ǆ�����u�B��R�x�£oL}.8��bC��M���?�+O:�qRL�i�S����R�:�Ó��8b�x�$ֻY�^�RH<���?��@�<�*O�O��EЁ��8��nY:����4��H�DĂ�mZ�����O��)]~r�k
����0D��%�'�T��M���?��/�"�?aH>�~ @JEG�0�S@��4�O_ަa�����M���?����Øx��'U� ��� �(5&��w� H�H��pӌP���O��O>���'h���e#�4g��턂57�1�4�?����?1��0:��'�r�'d�dV(th�,��,Ʋe窈ZW�=d�ƞ|��5}�2�����O��$n�ޕ+��U�C)��H҇ʜ#2�	lZ����΄"���?I����;�F>��ɧkI��!��w}��UI�'3��'i�X�@�2��M���`P�Q�~t�K�g��qtf �L<a���?�H>i��?	3g%/����P�9!��ye��:Q�>M������O��D.����a�$�'��:���V>؁S��S"�x�'���'��'���'� �О'�� ���1�33��cDfIX]�sX���	��h��]y"��pd��f��˴P��S�aؕf��A���ߦeD{��'<�q�'�BڟDD��-�:S:�K��j���ɂ�i)��'(�	�VE<��N|����1Xy~!�V�Ⱥs���0dR9Y8@�>���z��ax���?���e�&� =��选K9�ɫナ��M���?��K��?Y��?Y����.Ok�<5���숮|x�<��fĥi2���'1��J�Fi*qC�y�����"J���-A�E"T��>�M���
Zܛ��'��'7���>�(�n��эՇ�:������Q!��M��ʚg���jL>��M��(U�O������nV E�d�Z6�i��'�b FV���'$��ٟ$����
��K;fv���E�@?vn,��6�k0�|&>Y�Iş��	�Y}����;6�fx�B�@��a�4�?o��Dc�$�'��'h�up0县q*�4k�%u��㍴>	�(+&��T�'l��'S"Y�*�)�(�r`[E�{�p"P�~�,@�J<���?����'4�Px��2q����Q��>,!$�������'`b�'��'4���#L_�)�*5��)U�D8��A2!J�a8���'��'6�'��'N����?�M�`"�|m`���I7L�FD��K�}�'R2�'��	7>�d��N|���W,�pዒ���]'Є(�NY
 ��6�'A�'A"�'��}�}�DίFH  ���N9?~��{�>�M+���?!/O��B��c���h�ӫF' �W�	|1�%:�b�f��pJ<A���?	'��~���I��a�e
fg��'|�jS
�E��&\��Q��&�MS�Z?	���?�)�O��ٗGĸ}ZD0U&�\�0|���i���'�.�����iD�D_$�0�=8V@1��-ܩ'�V"@g�6M�O����OR�)�T�	ǟ oڗLټ!cP`� w��ȱp,_0%�憗��O>)�ɠlQ��ʤb_'ɴ\�D�^�y�>z�4�?���?IԪ�=�'V��'k�d��c��!@��1y�pG���3��O�Mj���O����O ��`�ހp����[W���I@���	->5��K<����?AM>�1T�+5d��I�@@����> �'�ҵ�=Q���?!�����.���r�X	mRHm�ƪ'(hE��.�a��埘�IB�埜�	�<���Q��A&�Q{ �qbN���+��ß��	џD�'�x@�@t>�B�P �����&۰���>!���?YN>)��?a��Bo}��ƒe���g��`-8���nR7��d�O����O�˓��d�4���dY2LXTe�5��8
�ʡ��+h*6-�Of�O���O�Mٌ��ȽT�by$��y����2+��M[���?Q(Ox$A��j�����ӹT)�А�!�3R�0���	(4�QH<i���?���V����^U��xːΜ/��ԋ�- ܛ�Z����B_�MC�]?i�	�?u��Or�b��[�ar��VJ����iMb�'����i��&���SJ�*�0MŹ��ڎ&�L7��O��D�O���Oi�	Ɵ0Xj�)׈��.¦%���&����Mc�N�{���>�d�!����o�(�H����ؓ_�Dl����Iȟ,����d��~���'���B�q뀴P�`��UJ�E!ӏ$���<A�A[��O�B�'�"n��hz�L	�Af��Q�.�.
�7-�O����UZ}�!�~����?YO��@m��m%���Ec�r���6�>9�E߯���?Q��?���?�a�)9��T�܉u�>yd��&:T���?y���?�����?���r���s���N&ax�on��^��ѓ����R�+ -#�8%��Y�� z�HJ-�*��b�$KU�x�E&�c1,�ad��,|�Yc����Sp����Q�n�ƤK�BT&4 i���Oe���=9qď Pj\���J43�tEI&��Fܓx��(����'w�2� S�gE��9�����ǖ1��|BnE��b���o�=�Iۤ�"�~dّ�:G�nm�"D��wNh��hH�'��
h#!jr�'�8*��up�P& 1���u�<F�$��c�Z�>���X/U����G���*�y6�? W�����pǂy����O�՚z\j� s��K1�=�4�L�tM��'�r]�WeZ3z�&�`ԆA<�9)p[>��O�`�@a��0��z#�ڢD��8O��6�صd���CȘ<(_���� ��]��ZEN���A�$`���ʐ(� 2��ƀ��ɔ#Qt�BM�)�SJ|4�c�3�@�j��[C�	މ2HZ-j��ٝt�Rd)笒I�l���ɗ)ƨ4q���%hj<�C/_J�xm�ן��	ן$���M�y�I���I��]�&�Z���vۺx�d�9�؜�.	�)��	��1�2�3���<��qy�C��Ol@����$V�-q ���Mo��Ko�(R�&'�3��Ǎ	 ��CK"O4Ƞa�?��$��Af�Oq��'�����R�KP(PN�*�V���'	P�ɗ� �N-���� n����O��Dz��ɟ1u'8���e�Q���$X�;�@���	TF���O����O4��;�?����@��'�̝�����`���X!�	�0qё.�ڌ�/ �"��yr�܌otVЁ����|t��վl|i����/l�mä���K�y��l�~�j�cA�4�fPp�T<b�5����?��d+�I�}���`ԌU&����v�B�)� ��f�B�L��ï�;���QA�D	Ħ��IpyBJS�jL �'�?`�J���qq�[�<#b�+�a��?!�!�@���?њO�0%X��	E"���c5�mZ�%���*S�B�R1Fۄm�:��$��|�����IvtI�3�e��=�tA��I�(�"�Ѹ�|�C�'� ����?a,O q2D�tL�m��ʊ������*|O���4��d�N�H1P	%�Rt2�OFQm�$G����,�8?���Ҫ[�F�I��oy�D̤{Y7�O��Ŀ|J�$��?�d)n��'P
����̹�?��b<����*�O��P�$ ρB!��PQ�9��e�w�ݬ���3e��˗�� j��x8��@t>��D�	z�MX b�o��C��%}��?q�y��$������%G�0)jD�
`���y��7Y����I(#�\�%���0<1%�I v��m�l��=ʰTY�i�+Z5jߴ�?����?)��
�^)����?����?�;aӘ(�FjO�kА��� 0�(�+5�@�]ݶ��ŋg�8�a�i��c>�O�ૃi-l|����43���j��%�8H��A̮.-��ccI��q�(%�O�p�dG)<��$�33��e��-Kg��21�����|�dҊi�b�a�AȻg��0���y�̈́-z� �.��n����#�E���Ă}�����|B��HDh�Z�FT�� 䍆VN64E:c���'���'Hj������|�"��j6�IK�ӴD�,�h�(:�2񩦥_�Wζ��_UG�剤�����D���)1�
7%�Py��F.
ozU@���Q���2	˓_�p���ƝF��=Ц��9�Asc�dy��z=8=���[�"� a�K�@��P��Q��kUÞj�TAI�C	��u�<�@�i4�'�@;�x�|���O(͋�H�rTb(��bG�i_4 :2*�O�����b#`��O� E8�<P���P��a,�%8��1i�{�b������H��x��:��O�a�W�Ĥ1j�A��m���B
c���爐5O^����<^]�l��
�M����"!���M�R!����pkτ�g�li1��T!|�!��'8�]�Q/��<߄��D)3+���D{�OoF7-V��E���N:rb$�X�i�ВO���`�Ҧ�����O�=z4�'p�0 �@�/��q���Bl(a@��'h��,�
*%@�<��C��1S�맶�I�}d�}���*Q4�L�!��+>�vͰD��EJqw�L�����[�ȅq&��0�)W�i>��m	T�(��*?��Q�2}b��?��|���*�'<$zq��gˁf"�uk����y�n�
.
�p��G�_G:ū�I��0<q��I�cM�P��	!J��b��XX�U1�4�?)���?!�0"����?���?�;t�XX��I�,�h1
'�1."�m3TJ��BP��V�F6��!"Ҿ��Oe�'�b�b�b��f������ȳI��
f�'RN�I#ui��z�΀��* ��O�'2@�%�Y�QP���u�����#�D�u���L>�a�&Cb\I��W�+�8�3��D�<����:=�#�9K8�;!�\}~¨5��|�I>YU�z���fD�z.yK���z���	����?���?!��~����Op�D|>��4A��r.D��r ?a�.��p�3\)Z�ɢ=JH�*ORx�4#'&/db]�(_JzlIs�Ʃ4$*Q�A�[�	�0M���Ix�L�A�(~� ��ŉrebu ���N���B؟\�tjE,�H����
(v��p�=D�̉U�\2΁;%O�H�ސ�#�-�	��M+M>Y&��>jn���'8�XU����bd
%��1Z��'�x@��'��3�.��Ktƥ�pM�1rD�1楋&q�t��!��^���x��M.%7f�G~�g	;��pWȂ�t�)�2� tȔ����E�Ɯ	�L�����$�B�DYD���'�Dy�i��'?�D`'�Բž��>�� �'�BM2��,ap��A��ۏ����'s�6m�'D-6a����R�����V�6���O��: ��������O���0�'˚=��Ν�J�U�^�)�����'8�M̚m�������B�S��X>x���;3�Y�� W�n��D%/}��L�j��(s3#�?��j�7F�ftѠ�'�lhP�)}R"A+�?I��|����Z/'Q��b��cu�����^��yr	/�4eч.��K�&Tz�OB�D�ў���HO�9��'_-��0c�gٗaGʭ�6��Ӧ���̟��ɨO:�[���������i��r4,ѩJ�))�nϝLǘD�%�F1W��A�'�P��Nۘ��k��`��gS�E��_�����}��yX�S$>Պ%���GAܧ]�t$�'���!��M���:IE7$8LH�7b(��E6$<��L>�&�˄L��4���AA��,*ie�<	���XD�eː>�2�ҁ�Xg~�$)��|�I>� RA�l^K%,�^$T�=�TO)��%S�b�On�D�Od�dú���?Q�O�XBT@�*rt-#�b�<!�J5T.v�(��fۯ�0>�HB7F��.q������H�H�0B�����{���b���hO$ѡ��i����ΜA����3��F"�)�O��q`
�O��u$ԆRi�0#�"O*s�
]��hu-�T�\�{����覽&������#�M+���?��7>T��0U�
dS2�R+�?���o�4��?Q�OJ��ٵ�E�g�JD*!1B������
9�Δ����'��'ͣX1�#?Ʉ ُ?��xg�A�}����K"�X�f��><�ȥ�pH�M�����L-[6j%FxKF��?��x�	ӱZ'�M��u{�)��-��yr!9��3�,x�NB��A�'�L6���Vr&�W0[�@U󬍵e���Ob�"��������X�OQ&\�W�'����ӜB���K�)Xb݊�17�'���קR��y�o�J�����oޜt�,]�'���^<8e"x�LT0P�p���d��CϾ��� �,M�v�@9BZQ#%��P�*��N�B���Q�B��!�:}�p�T�~ȴ�'�u���h�ɧ�O$|hA4��*��=�rE�0�d���'$2�M1����_�a~tZ��i>����D�#�<�qf�?��h�
�;�^`m�֟`��ӟ�HT��N�i�I���ɟ�]�JT��09�}�b@�$���c�'(}�!��{8Y���L>�f���	g^�K�h�/ؘy�F�\����#`�T�,M#�i�sѾ0�}&���$�[/ �T��HGh�,Z�ʚ<��Dl�<�)�3�D�]�^�a-�5�"Qxsfgh�'چ(Y��&^&��y!Ƅ4&Dq�O�MDz�Oc�'}�̳ԯC� ���bU"&�@�05�,H��X��'d��'��g�U��۟dϧ'��իtm�;o0N��Qg��҉J'R�J��<RU�@+*���i�h�P`N�%p��90�K�,*�c�2=%8|X�A��5wl��D������B� �ib%��e�,,�%eߕph ���'�����V���4���V�n�H#�! �!��8����W�9�̹xBE�`
1O2Do�J��̬U�޴�?���z#\�@!H]�W,e:�:i�$@��?��L%�?�����T�P�{�J�k�(��^���{��E��B���V�{u��V� 
obRs�8��L�#I����ybN��}��0�('O�vuq��2g���$C�������>=�Y�՛|�.���?1��xb`��q���3���*9�1QS�@�y�eH�,ظ��28I��ܙ�O$�=ͧR��&
�>p�j �Gň10�69�s��W��'�4˱�i�@�D�O>ʧ}��z�9��0kpʋ�3p��Q/�m�������?�@GY*�ҭU���0끌�;_p	�����ɑ2��R2�«M�h3t�ɋ$j�t鲭qe��%IN�#Մ�`8������Y�r�'$�*��`�5��"�#S�#�8��OT���'�,7������I�'s� +�b��r9Da"a ݱ2�X�<����<�eZ&.�X��Wo���G�z
���dTR�'_�4b�W&�n���!C����1�i�x�$�O��DB�?f$���Or���O����iW�R=U�:����O�	6�y�E�`G�	�'��h��������fR�Q%k�3h- ``��W��A�Ö�d��P0�ğ�03~�(K|ܧ ܴ,��O���Wk�U0�JP�\VNACN�[�^VF���|LJ� �&ݨW*\��6����0�y⪟���K���7��L�ŬZ$��$XP�����������\�� Ԥ�����48"@Yb��O���O��E����?��O��PQ��\(@=�b�!zW���m�g
M+`ފ)ǎ���'M���$	�J=�f�T41��c#��
@)"-2	��X�E3R�6H�퉑JK�LH�gS/�b �D��;Њ4I�E�O8���ɣ/�f��3
_�'0�􍘦e�NB䉤+���ar��S>"0�Q�%)�b��J�}Ö�'��7��Ov�D�7w���*��õ���F
�����$�OFH����O$��f>�S&∄�2@GO�&6���r7o�n� R�J���y�J������E�1Q��RӅF�81^}x�O�77xȐ��ƕrg��A�¬u��%Q�OԲC���Htƅ�'Q�[��O|!%�`Ò��U�8�P�P�YV2��I4D�̰�蒊;��c�<�`1�0KܴZ���8�fh�0�kT*Y�rM�<���#_ě��'��U>9P���0Ф&�9q���$��=�I�R�������imPMBІӼ���ѥÂ�8ȕO��5&���*�&Ìb�i\6V6�'���'|�r����ڣe�ԙ�*ѿ��J�Le#t�'7<u�f�d�O`h�t�'� �O�h�B�����2	�rt��pp"Of�X��'%��(U�P�fԝ1A�'H�"=��=f�]C���wtz�ʣ�{X�v�'Pb�'�t� ���|�"�'�B�y� 0��F�0rw��Hc��A9J1�"3�	�vU���D\�	8h���uX�z �8^ qO���'�����ݗ!���a"ša��!�s�+��Ša���L>�VhRy���fD�b�l���CQ�<QŊ�$TE6��F���r���/�V~�b!�S�O�
p��j�'���z�.T
0	XY���'�b�'�R"d�M�I���ΧqH(���Òľ���0b��� �'�~(��K9�a{���Mq�1��ӦM������=C��`p�AM�C0�mڕjͱ�hz���_�'�4�ƭE>$b�1}f�����?���i�F7�O
ʓ�?����.@�I��(��S�Dtz�-A6�yX�1�tT�.>H�t� a-�͘'S�7��O ʓ;����@�i�2�'|�h�G-�d�2�!!!�V$���'����D��';��ZR����S:����6���O��5�JC�l�s&�/���f��G�'��#�ւ#���C.#K�@�@�V����_	<讔��ל�Aq�-X3z0Y�=�V���tKO<w��-:X葑Mg�@X!�Y�<�ѡW�3�}��DP�rV�KgMo<I&�i:PI��w��:�_y��D��|�*��g��6-�O��d�|*d��+�?!��)�vI��ȦL�$�C���:�?�aZ��������<��,�'�|(�c� �Ut�`%}�#U�O�ƭ@E'�:Zx��@�N����3�>��Jܟ`aI>�z�� "`|@���`@ⶄ�A�<	U��>�r�ö�@�OG�%�2KLe����DϫT��E�c��9�z�� \�o��n������ß�Š�5�P��IПt�I��杏Ot���Q�Q9O��bt&�[i��a�()^����L�Ro
@�5��O̧e� 6|�ڐLFVgҁ��@�rZ�
�g�4;��a4!P!o4:� H�W�4�����rFN�ywĈ{y�Țwh�a~]�#��YM1OpM����E:�RԭJ�I��zf��YkH��6�$Qʐ���/ �Mᕋ[�k����'��#=ͧ��f��|��[�r�L�2L>�rF*Y�C a!���?y��?�����$�O��8S]�� q
��e:��v잋CQ�ѓ� ӊ'�8d��[\��-1ף����O��X����B�*T�
�2@/I�m��5�)=^���ط�N�2�t�5�i③�,�%��'�"� �Jp6i:l�/r��x���?��'o$P
�D	�\��Ձ�c
OS�T$���u���[oL�x�����,b�E'�I(�MSL>1B�Vݛ�'�"N�~�,ձ�EW�U\2�"q�����'a�41u�'��=��i�W�Ow3�#�N���Ԋ��H=ݲ�p���/pj!�p�\�aPHF~��8����C��,A�$�&M �
GdŽA�>e��Iсf/(�h�̷I7V�w��Z�/��	�I�#8�R�싛"���9�@�-$(B��v1jT�5=^�Q2�� jB�	��M��(ڙ8��lxDMQ"rzd��"����:#d�㠲i�'��
w��p��?L���t.$������t����x�fO~j�9��KG2S�+��C`�i�|�� O�V|���E�6"��Ů�Q��ِ4	��MQ��`i �N}�� �aO�I���OÎ��0��Wfl,��c^wh���N��xf��Oc��?�9p
t}v5�u���j�Ÿ�d%D��#��_�9E]�����
G�ai7�&O�0Fz����c�E蔄K)<(��KJ! z6M�O��d�O��Hf�B>e��d�O����O��)�����N�*���jM�[cd԰A
�y��t@c�6*�$ G�+����!iQ�d��a��)�84�� یՓ'���Sz���	O�6a��`b���Y#2�O�Ժ�Î�;!݅B�=h�A���c#�Q�P�'��C�S�g�	�JLzع�@�>�(���	.�C��'hbU�V��%�Ѝ�E'�.^��%����x�ɥ}�԰R�
cV֤@5ʞlҎQ�S�I�[Y����ß��	���Zw5"�'Q��hp�#���`�g��w�z�WL�'P����A	�hp�h�F�'1*�0�-��u�x�&���:Q@[��tQ!�
d����0�4�Ks��B�8�9�|˚�WW���6��-I��!��Ư~�ĕs�4���v�㟨����C��a�A)�-�X*e!��y�Ο<u��A�4�=�F8	%����'\7m�O �S��A�ҽi���'-N�Aد(ڼ���%S5۬Q��'bn�*V�'���6��a�%�n��@H3�.�3�.
�mAFx@�^)}!��)4/O`�'�*Y��� L�L@�m��Θc©,�f�&tكm�B��Sf$���� _��@H>������PH<��k��EƼ�@��"$�d���U�<	g_�O�"8��H��{�b�2!G�S<�i=��Q�nSH��c6i�@�Tyq|2��j�V7=�����|*�D��?1��愻p��r�=�t����?���$(xR�i�;}�x	��Y	��4r��?U�π �q	`�ٓ��M���G�l �	a�> AI�<a�����r��BqB] s�01���S��Ӯ ݀���ml�+�(��'�ؠ��?�����OBܪ�N�>�N���Z�hS��ʃn%4�����3m.@Pä��Zf����;O`<Gzr��&��H��a9{�H5)���e�H7m�O��D�O:���k@����O����O.����쀀�L,D�sRB�|f�E�	͎2���"����d��)��ObZ�'>��H�L�5�	��N?-TZ�$� ,�� d�B��H�"O�J -�H?ŐdƂz��.O�9�r�Q�r�8����%d��\&������Oq��'mTh��Ȟ6MƉ{� )q̘)Z�'ǘ];C���"�N�i��"@e�3�O�`Ez�O^�'�lU�'�۰d�`˛#,�9��L:
|xY`�'���'��}�i��� �'���a����fU�V"OOu+FT`��{�T@\�7�\�%��Lz�GX��� �eѠ*����V�W��f/9m��s���\Dj��6�n�:E��dƷB¨|	Pn^�fȘ�z�dV.�>��2�'u�7�I�!�?���I�3q�I�A� ����͐Ue!�Ćz`�YS��~��� " 	XD1O`oҟ��'2�� yӔ�D�O��dƚ�o^j��Ǭ8����d�O��$��h��O��S�[1ƁX��ʱ�Zl���q
X�2��ZC`92��IڜŸU����O�pc!L��e����*B=py�g�S�]\:��eL�zQbe��ߔ��=X��^�YZ&D���;���Y��{���o�韼��`Y�u� `j�bM�&��
�jy��'|�O>Qp��Ң'���@2��?���c��5���ڴb8�G�O�;������[�X�����$B�x*H��d�O����|��Bآ�?����l���jV�e�h��K��?a�F��y�阧� a�`F�8��q��h�<� �,}r��y���`J���H9"a<�'a�l	�S��E�T�
�K<}�!^��?�p�|��t+؛hL=������@˃��<�y���1��Љ���o��myt��0<Q��I<1J`0D�%�VP�Ã�*����۴�?Q��?��� � �ڠ����?���?�;s����đ6ʠ(���_�ߞ�ʢ��k蘜)�*��?��������O�$�'�j��Cᛴ�hX��
T'{��֪ˣ	xv�C�����G��H��'�|:'�>��<mXh�`T>a���R�q���K>���R���>�O������2Q8�]$1��b"OB�ZA�ܺPfF\�d�̸D/pE���pC��4�ΒO�E�6$EdXJс���P��d�fl��!UE�O"���O��$ºs��?9�O�r5FL��N��*U���	�$A^�R�D���ѻk`��lM%~*#?�g�ܺ,9z����)~d�ө	s�p4Z�F�@�0�RGD��5It�i?2H�$Wj��'=0H���@�>�R�#��&Kn��ο�?Iúi��'���'zb�'I�\>�#�%Y����$��6��{�g=�OƒO�e�dhG�Q�v(p��#`	 ��D���	Sy�É�Jr\7m�O��d5?f��2��[��d����"k2���O�1�R��O���a>�K��%b���:][��򣰝PL�A$��n��l��E�4x��������ĪŠ�Wdq��K�4KZ��C��*����)�����������1�k޸�O���q�'�O^�@"0wg��g�˸D$�@h�"O�����]��h�ǐiēsOqoڞNHŘ��H4l�;`C&�`�%� F���M����?�*��$��#�O���7�LOHy�vOGi�h �L�O
��V�]����J�;��1�4�	�5#����O5�>j�FyhC�ļ�`���ؘ*�'ZƑ�ãY�1Ԝ�����?N�G���=Y�պ G��|Ѝ�o�H:a��?�*�b��JB�$҈'z�#-���ɬk2��GCBA,0ʳ�H�-!�S�k�0D�+=BF��ӱB1�axr�-�|z���RS٠ir&'�2������i{��'��%מ#4�EA��'���'L�w��	���� n��<)4��O&tA��;k�˓#��ӧ�b�g�L�ޙ��Ŧm�>����dɁ�gK<d���>kh�]
fd(h3q�ʕ�O~X+�m�R��=:�?{�F�����Ms(O��Ӥ����?!��?I�i :���j�Ըm���'xx�bʈoy�xɲ�؉8`���O�FzR�O�2U���i#���S�HI<&0�<���,6TP9�o������@�	�2b�O��D}>-��%�;A��u��gM)5���Еc��iT<rg(�5
� ��dPH�G�=V��(��k�89x�*�|��y6뀪L̽�U�ݛ���t�	-�����%s *����@/%(��$�O�Pn��Ms��d7��+��P���L�XM3���@:�C�6pcJ���Ɍs��e�Ǉߎ<�rc����4�?),O��`K]C�t�'���f���\�tt���A4K����'��I[�|�B�')��Q�e�luȦM�o�*���V_kБ�O67�D�@��G��hiD`,���8�s2Y���k����� � &��[�`bk׸l��\jQa�b��֧�*גA&���և�O"InZ���D�+٤ѹ��I���-��aجt�1O��D9<O:�B���Jg�,�1jI�A�P�3O�Hmڛr�����o�!�4��Haj��	fyb뒭s7��O�d�|�1���?QA�̶r�.��3*S�喌J��]�?)�6��uhS�Ġc/�)R��u�*�P˧k������WA�T���M�HݧO\�!�4,��%+��D�`a�EܧR��A�:��i�@��o+J-�Ov��6�'1O�l��.ӥ pY�@,�C����"O�T��KF5F�x�&�P
�L�p��'�T"=�f͐_���o�&0M\<z3�V[a�F�'!�'�r`��'���' ��yW(��r:DiCZ�A<�h
���%��,[�%���j:�#D�v=�`A�|�Nύ1����d.D�p`�0���ť'�nXi0,]=x���(F�lZ`+�����Ӊ1�����2�ڨ�ɓZ����ǣڌB�E�1�0�	�@����|͉%�<��o��T@Q��H��y҆�<A �p�������h�	��d�K�����|�o��j�A�2}�|�Rǚ1`.���EI'r�'7�'fםßt���|�B��$�+ҏ�ȄYYV"^��*1"ʧ��>ä40���T�ܷL��k��|��sb�&��>93bԅ�h���.)h��d�ND���ğ̸��Kv~��"H(,%���-��WB�Ʉȓ)��l:P'Ōta� zg��;?�6��<���dU^�0`mZݟH�ID�Z�CVX	)E��:���K�$�I��d������I�|z��U߲"ӛ��ۥ&�9D��ؕ��G*�4NǈVx����fBP�'U�7�]!k�exԩ҂	.��+W�܏1�Miः5`D	^B�џ� 6%�OX�O�S'��5< �HN�Pׄ-(�"O�L����4�h�����D�v<H�Od�mZ
9:�X0o���hL��.���b���� �?�M���?9,���`�O�h�K &8�6�q�4,�pM�� �O��d�\XM�1�Z�X_b��1��?8���O��?���Rǫn<���V=p�D�'���9��%M��ɣ�G[�W:�1q��Y�tWV!äb_������dm�&���ɮ��S�'m=�
�ύ2[0EF��&a�1��,J�;C�͜Vd��1���l��$��	��HO��z�.Á��y����\uN�cS���I�������G"đ3��ğ��I��H�i���" >1t��P$ B�h`��R耕R�@p U��?1s�,�N��|&���U)P3��]#�n܎�D|�̇�j����c�T��?�B��8�<�>�OM+��Puʈ�+R-��[;�<r�-�I�Y;����|�LZ�P`���۳\3��p�ˑ�y��#j��!���T�*%�7�ծ��D�s�����`��ƞ>@R����?��q(��O<>��ړ��O����O��ć޺����?�O�&P�դJ�4p2��2:�\2�FV�lM��jO'Q���%,O��靭�N�r$�şhOT��P愐i��YB�	�2u�@�C�DX����֜w�r	�#.�1dH�!���|�h��p؟h" �E�筨C�F�smr�p��9D��Q'!U'=��*�C�3}@���<���'yU�!$s�h�D�O��Rm�*VE\m��ڗ"����0��O�D�\����O��S�a)�y"#���:U�J�OdQS4@̯8���JS�]F���7�'�<���ʃ�NmX����Ъk�Й���J�i���aG��/O�����E�.o˨\��o�f |c�y���?��x��+R��	��D>Y��
f�Ї�y�-A '��0'�I4�������x2�~�f��A?��{���c��GK6���}��n�@��S��o��'*.��R@:��Y;`��K��|)�'e"jS�5�.�����L�|�Q��&+�`�����0i-�1tGQ*���e	�'G'�w[�����k�P�K�<��+���OB�-@�2BH��$,���I#g���Dn�)�ӗj��$�V,\�<��0�U	N;��C�I��\y  Ǥ�Ҭ;�e	����|�'�(Y`mP1aJDi�(�D�"�`Ӻ�d�O���φR	�`��O��$�O��4�f=�g�#m�~�r��#�:x�F-��IH�(D��X�dc>�O�L�2�B�=���Q���+E�|u��F��*��`΄�MCWN��N���>�O��c�w/�{rS$9m>���@�%;m6���|�h� ^D	���
3$8d)��yr�	Z*�Cɵ0IN��ì�	��d�m����#�%Ӻq��(�t��T��cT��GJZ��u��O����O��$������?�O���p��1}P2	i!�b��ӳ)��x�&�h�����5j*�H3�����0��'���� d${@h�d!����(9��a�V��Ov����6\o�	W(,3nͻQ�^�t�!�d,r�h����.$�9J%�Kp�1O8��>q�Jp�v�'�R����蚕���dak���)5q��'� |��'%1�~T��'��'�cv́xPP�H���Qj�+Ǔ$}8��?a�E$g1��i�FȢJ�� ��%t8��У'�O��'�Lz�jY(/ڈm�����{�/*D���#L<�91�"<O^���C(�(�4Q)��Չ@�CG.�e���.H,�ȓC�R\�3��#F$�H���;H�����8�┏(�&��3�@
/0M�ȓ�2m�= �v�wiC t�:��R��I�T�J����[�q�dY��[5�y���
�_o���ьɶk�p���C;�`��ī=���B���D!T���@�
����S�`�������9
�M�ȓT�丹�ɑ�/)lm�R�G��0,�ȓ<4���̊�Y$=�Q�� 	�ĄȓH�v��7��)Ĭ��K�J����ȓ#�XЊT
#]i"ݱ�T�1�8A�ȓ,��y�ʛ�����b�A�^��L�fH�Gl�)^����u\���ȓ<�\����4e�	a-�@����W8F���㓉:n@�X��$~�0���qBL`$�Nh����S��8|J|��}�8��Kˣ��5���#^�|�ȓr�~pP�Q'F�#EJ�%c���l� 3C"޲J&JUxQaT73ܰ�ȓU,�U��ϕz���#���>N�`��ȓ�p5���X�ZL�C���)��}��k���Z�	�4Q�'��0�Pl��h@�:�Oҝgr���ɵ1�l���:J �H�*{�l������ȓ<1Ę(�F]a�.�q��H�=�u�ȓ$U���S�����p�:���C���P��&�8�
�6� ч�IF�0Dk�^���#HԲB�q��-��M3�?8��C����6�PP��n��у�*C�ʐ�Q!U#-~��<ɔ�
�dɇE^���E&y��[B�@��H�#�9��J����ȓL��̒�WMMU鷦���l�ȓt�N�b�W=�8�� Z��T�ȓX�:Fo�Jk�,�Q�E� %�p�ȓt�]����;#�|��G\�)+D��%(�~�1&�ч0nar���R�g����<h��0�L Bj���P�_6F!�$_�L<L���4d�j�V�PZ������;I��HGnρf�`�	�>O��z����\x	�ǟLmP��'����J�ڡZ
3�	�F�&PMZ�IA$F(I߮��4�0)$��$G�s9��+CH���%��%ٽ#�'�6�Ir[�;����w&��;��17�	T�c�~D��g&p$`أ�à�!�D��2L�w��k�D3����p�D��(�;O.к©XS9z�J��$}�'��y'��񰦄&��"��x�b�

ql�`#�<�r�H�GS8�F���/�4K�rM�� ƫ@�4��U�'�9�M�x/:�)�A������%��3[Ա���R��	���O�9O����Nɝ:����Ŀ�F��e"D |T m�w��YC��jT��PxRb��(��#'Z�K�6�$/�$���Q��/y��"J�rm�j�[�8���p�c��ň	�u��ɈS��-ت�kaJTs���R�O+"��`��ݽ5�n�����p8�D͂@#J�S��53�(KS�/I�-
���|j#,���iU�;��ܨp攻Run�"��!�%1q�M�'�n��U��	7%��@AHY-�$ݕ�MKe��A��[��tV,M��g]�fYt�X�q� 	 ��O2ם#b��3&A`�Y���?9 ��JY��0�o�B��op|���M��R$�8_Y�a¨��H8O�يB�30뎚�{*s�^OS|��ꇱox"��!1�T�0MЇ}.~���������<[��{�G�D���J/}n�÷e�'�j���I�<�g�?x�搯��ez�H(}��i;� <;%o�2&��@Nۀ3���ѓr� *'hҟϨO�:��[Q
{����O�8@ᖅފD�B�4��h�'������yr���8��p�J���Բ|(�I��I?t�!ѯۑdl1�7C��OfIq�(�cnɨǪN�cI,�`���r6��K��e��%�6r���W`Nv���lW�IcWm�3~��a��O	�d��-�2]��Sh^:�����){:���1��C��tSd�:�����+��_�:|r��X氩�����5��% �u�OtI��;dRF�T)$4=� Q�'��;�0�A"eԎb` W�2q��I���O�Q��{�oCNM8��I�#
��C�oʛW{f��Ħ��tx"��?��ɩ� ��<O�m9sj�.[�P���:ulU:�E#4GR��1���p�Q��&��e��g!N睺x�,%bTFQ��,EX��#<��ˏy���y2�S Bm�+��S���LL�%�!��Y_|��K�`\+j?�-QGቚejh,p�R�~6�eɓ�јT~���<�K�̙�8�x{��]�~Q.\!c��y"΀�s��D���ӧT�F�ɉ�xjy�}r��QKRI��N-N�d�`A�{����)�6,&��pelZ�H����c0ORH��^Sζe���Т�>XA��g # �Y�~�hU�C�5�T(;RiF����V?�Gy���T/Լ�EL�Q� Pf+¿W�.�H�'�� Y�N a�2��O�Խ��D�j�ɽS�>��O��J�"���݌Ɯ]���7AuTi��"�:x��F}b��h�lPQ�w>$�1P\��(W%�,{� �=r�Lu%��-y�8O�8���],[�2�0�ҟ���t�бF�H4�g��:9���q��1��"<Q$Ώ�'��*��˱1���k��^�<9� �yVM�$��UK��{P�� -5�舕?O>a5lN�C�:)����?M� ����O+&	0���#Fc��{#-]�;)M���� sZ�<`0��wRҴ�����Z��<�s�a	��>{.�����q�����D����ϼ}��ASS)J�j�'�(O2�B�����q�'Ϯ}��L��'�t�Q��	��X~�s�/��<�'�p��XF(�&�h٪��ɪ}��\��N[�!�H`�����O���3�ڕXn���R���P�Oɀk�������l�D�?�=Z��O=U���S�'v�<�#��9|�a;�!�9��ђ�����O63VG
0��=�rdSW� �!�����ݻ�>����ʪ� �%�����
j+U�� �4�j�&��O�q�p�y7�ѠX]Ƒ"��c�4QC���w���m	B�q9��X3u���y��4�GCA�z��Z&�Js=L|k�O�.��cߪ%"��3��ԗ{�p讟V�<ai��̣W���0�w�S��r�铢9tʘ"��1f{Np���Y�@�;A��5�ږ=�z�AC�T�J<p O��l�Ǡ7�O�E��M�Q�x�#���J��=���O�X46�ς��Ml ypU�����:��X
�"�1-�0I��ʇ*Q���'T�ͳ�U�){7錺W�2�Y���`����&��7ΩyE#�u��2���)��r܂h����U�]���X��	�`�|�9���=�nJ��Ӟ_�܅A��$x��E���8����M8d��I0D��QR��L<�G%\ x��8gfH9�|�qS/f}B��s���⋝�:i0�E�&Pf�Z�ؐ��?���(͏S>�b2�E�M�J`	��'{�hBS/(U��5KU'5t�䈷��tuR�P�Ucy�'�?��}��'��,�ԣ��
�y�P�{d$�
�@�q$+���M ��	(+|,���J�h��( �S0@(�����ג/���dH��j(7��HA�Ӻ�`@��@�8���W<2��'���~M9�M�o��m�?��叐-/xej'-^����v,����_�VIE��H�!�|��/�5|N��P��h3([�o_򤻂��:h�!�Ρ�(O\ka%��$d6Y�F� -�� �2�ՑV�2	JFn��*4��S�2nS�)��D����h!�09��*&�3�*�{5J^���cweɀv�b0xg����p>� OR.��A��z#G����Y�'!8kY0!V������*�5���F\�ћOik��t<yp֡X�X���Lc�2U�'�U`�a&��z��N<���F�
.Xcݺ\��t�Ke�	%��L����3jU>Z����|�&ފqx0���:Q,z��U-�bw��e� �f�&���a��&x��G�U�x"r�^J�$�]�v,qQ"D
n�acm�$S�F�{��
Ԡ� #Q�H0�cT�7ۼP�Hz�'n�Uꔨu�X�(٪)��O`!N�Xcd�埬8�J���⌘�y��$��3it����O�v���ʑK�>}���0E�-�d�
��� ��W��֘�t��4�CI�=�I��R*H�IS�^�z��ء/�Z�L#����T�h4%>�CDB�?5���%
1�k���">��TB�M.,Obz��Y��h���h��f]��XP`�Px�c�"��
���bάaŦ���_��x�b�C<iv�[Th"�T͆�|���ڛw�`h�L��<Z�pv��6x�n}�K<��L�-p���d/,M����@k}�OQ�i�b.�X�`뵣�3.5�/�"��i��%�>���6�Bjq��#f"�68�RaDy��L�SL�����W�a�Ƅ���S���u:��[�JLx4�f�<��}�1��l��Q!�������2�|���1��4Ó�%B~I"wd�78<��i�Q�˖�T�N�P�Lˀ:q�6���@r��*D�Ԑ��æ9@�m�����O�(l�aC��y�ub�l�?��)�3���a~ay�F�8b���Q�o�?OC���0'C�^�*�0NH< �p�x���o�4�!��� ����3=�H|���O��#,.��uPX�j¢��u��)�+�-/�O �WG$����4/���fk�>�O�@�bs�ʛ#\h�ƌ��h;6v7��;��n��iHeh����ቿd��!tlG�O���0���Jl�IBC�x�d�-;����~n:2�c
`)~<0bT)�6X䨐C��A���#s�F����� ��p��~M��j�%P��1Q����
 .��g�>%>��W�3 c�h �p`z��Gھ �V�����.z�|)`�c�V��W�*����l�&t�9��aZ��t��Q����K>as����-�74�7枣1��O5�3qu��2̙\yQ՘|ZwT`���X>~�q�+N8�Er�OX���+����DK-��@g���V�Fj��kq�Հ4�1V��
�h�n�S�O�tA�$��tQ�o�C�T�TO>��D�+:��측gt񪁊C�}�	<4q����{2T��b��N,,�K�a��@�T�$n�&0N�@R�'��A������1�>Q2v�ץ)�L�'�y%>Y���$�
F.��0퐹Iu'|rJ�'�lt� UuZN�r�d��C�z�@H>q�l��z�B��V�X�PR��Mܓy�AJ7�/U�%E;]��՛g)�4�@��Ui@��$���G/O\
p&T3n`]6��&2EJ�3ԓ���&d@/䊕Bc����΅h�e3�?Ypث���	q�d��N�A.5�7��������Q�ʗ�4����ωL;��D@X~�'>̤����>/��.��[L֌�*f*�h�.׍�a~��֦1����hC�0~�u��E��x/�b@E*��'��J!��N��� �Mq^2L����J�h0"���H��]y '�� x�F�-���x���o��"��i6�P 
��g����1�{P�tSbk% �y2Aܽ]c�лm\W8�:W�:cZcP�TW�=hác���5�EFeL�2�ȡr�*%x������8H���)��:/
<+�� '#�	w�L.I�2 Q֪Г�0?i��<�܀��)�N�
1 I��Jn,�p�:]���$��>1�G�S0C�	�`�N_܁�!F
�I�`�` ٷ@�NpA�G ��O MH�C%CI��s�(�'�i��C	_�`�B!�l�GȘr��Py�DHB&�36Dv y���	G�џܚ����KY
�G-������3E�>�V�*9�\�0���in�@�O�Ŧ5��%��O��ѷMÏ�M��g�"4����F�Ȳf~&G�Ri�(����4�r��ϷZ��Y��\
?}��I�@7Z�}���ic��a��<�H�aF�OX�)�.ٙT�����w��j�ҷB�P1UoW6�A��rh����\; ����#��A@xzpHb@�� J
,02���G���b��L3{�����+���@�O �"HB�)�@Ƀ)R�~����		 �rM�B�Jm�G�N� ~6��	P����@X*&t�ɂ��~�1ل��x��� vH��lh���׭%��j� �k��u��j�
��Ip��\�Ҧ�k�Q2��ƮR�n6��/U�T�1b�8Nn`�lZ(>�V9j�Aޕ8�]�������Y �1j�l��I~i3N�`LАj��?��ii�IR��:P�!P$�<��n�Q@���w/0L+ӥ�q��QȂ;}��u3��.&^a�RNXu�x:���9a,j�z̀�/u����G��'�ª�GQ)��Oh}�����I>�c�B�HΝ �i�,^��� �x�'�bD�t�9�$�b��E�ĳ�4;E�ڥ�L
L|LcuA��\���׌N�"؅�@/��49�	ϓ\4\y;��c�\�CȐ�(Ċԗ'��q�'��)V7OyC&�Iq�1p *�f}b�r�e^�;n��w�j���
�@���B㉠�0���}U�u�$$ޢ���1{���AY��bQ�
SV���T���~�*�^�]�r��q���y2k+q"(
�d#$�����]�3�#ꑂ`�F1@�(�^~؄���L>)sʎ@�<�Jh��x����b�<q��@�."rm{�F	5,)���]�<)��V?�|P3���0�p1"���]�<)��~�� ��儷h �!� �]�<y�-�=E/܍n��1Nd�T���W�<���!�&tQ�������ϋI�<9����`�1f�!Y�p��K�H�<yVCXB�@�+Wq�q(шD�<!���8b?�,��T�0du��GA�<Q2.�/"��Qq�A�E�nu!�%�G�<�wZ6]@�����2��K�G�<��&����j
,��7�k�<�B�C�A�� G��d(����^�<Y�)=��ۗ��R�(�sq�~�<�AIϳx|~�`���y��Q#��P|�<9�*V80c�� G�Z4�₏�y�<��
�eN<�iD�@5AF�`B�r�<����%�8@1�C�3N��ճ�m�<��5qgl�A(,V覈��j�<��U;.�U3�B��Mh������a�<�w+Ş(���_�&�����N�C�<� ���v�A0���9c��1a<�:3"OJ���M�#l��c&N{�Ҡ��"O�}zŠŌf���sP�0OپT:c"Oؼ�U�<7P\�4"�1��y3p"O�lJ�`�-+�\1�#R�A�0��"O�H��N�j�
m��b�:_����"O�5�Q�P	\��p�.ή�,!�D�KO&ԙw��	;cl%����r�!��ܭ7�R+R�"c�xA�'FOx!�ĆJ�����f�+R~�G�	�^!�d^5[��!)&+�Y#��"Եz�!���l��Mk��	|d�X��nA� �!�40yD��@�pW|Ȃ6#J�n:!�d؍4��řF��(G;rU���RO!�D��?��܈��"8�0X F!�D�1lr	��-i-�8Yd���u3!�d�|�|��,H�c���Aʡ?)!��6��H�E�����P�r�!�$^�Ĝ�D���a� ��U�}�!�D�QrTpx�8Ѥĩ��K��!�D�l�t�R�5L��a��x!�ć�2��C�/ �^]�&��H!�Z<;,Xȓw�	� ?vm�c��c!��,@>�	�A!F�>�	3�z/!�+n�
�H� i�h�+rCA�!�$T�/zX���<=W�(����84�!�ޮ-����)P6		��C�m�!�@Lq����&vi^qӴ �>(�!�d��8����O^�eT�Y�AE�7k!�$S*f�4�C7�ƙ��x�G�W�^]!�D�)XW����'�����N��GT!�>*\��4DKQ���8��MJL!�Z[j�T��@3[w���� M!�D.=�DEA��Q�:�0�J�-�!�>W��P{eF �\�8a)��.#!�S�y�������_�B�I��S��!�V}�xrbH��^��	�z�!�d�d��E*B+ԞO��`8�]�c�!��p�����*�3Gt����&#�!��8M�@�P�?}�	elCR�!�d7P�P=x�oJ 1m�B�닆�!�d��S�"̀��|-��@�7�!�S�p� J4��Sͺ9�WmJ�c�!��'-��cɁ�L�p0�����!�D�"����5-� ^� �Š�T�!�Ă�V-�x����}�A7 ˇ![!�d�;#Ҥ��c��B���S��*H!��4x��Ǉ�!����� �F!��t .��4�O$�HӷnӭC!�!��K����R �m�:�!���^2�%�B���O��B�&�2y�!�$��T�8��
N�L��ѣ��!�dT�qON ���_�`ƈ=ӡ��!�!���f�>X�sE_8)��$sӉǾ�!�D �f�"��$ʝ�4������!�d��k�zy��R�d�Uc�>+b!�� {fX�2F����V��%P!򄝲�^8�����#�ޠ����K4!�$W-N?��b��Ǟq%0`x��Y|%a��O��7IF��IFaܙA��k"O���r�'����`�
EI|ф�	z�OɆiR��^� r��2�@���'pҝ��� �o�r�Q�͎I9~M�'�t'�܎	7Z�!�Y�8��A���� ֱ�Č��S�X�CњS�4�rG���>���C (����FL�#&�
 ��d/!�dC�?ЫFʓ8S �2t�"l�nPDx�'�@�95-ň� ձ�J$t�BU)�5qA�>!�n̒F9:`�D珪E}�д�h�<���:G�
ͳ�H]�/b���qB�K?ɯO*�Dz���*
:�h��)��ѢC���y��  ���\��X B���'y�V�'<���K�|Sh��`�y<z�I>I�e��b��>%UDK,���u��:".�dhjV��xB�4>0�e#�<����|=�OX��3?�4@�&p7�跥$���p`�YA�<1ƉD\&�
��;o����̚���xBFBEwLq���̭@�\�롍�8�0<!�O�c���Q��,������{�t`���9D�TQ�JS�g��ҮM�V�V��9}��)��);�|�y��os��0�e��I�pC�	�R�DMPvJ]�C`�t����/x�X��hO���7m]M��NR�..0�kF�YA
!��`L�I�@��5���ɠD��B��x�/c�N�����'*x��at��xeC�I�P�t�u�UE�NH��Q�L�����"|�fR�x�RUnˈc��=x��HS�<qLY�.��$�u��Ah��c�CAP�Ʌya{rL# ܀`��n���Ȗ��?�r�m� l!DJ�!m�bp�6`R�b0d]!7"O("�ӧ%�
����ϵ.�L�q2O���DR�V%�%ǃ�5��P��!T�%$�}"��D�E�W�W�*�AW�ߡr��n$D��HD� �V#����G!t�@�G,'D��R$Ξ*n�������,�4X)�"8D���@g3 ����^(qDo1D��H���q�&UKPk͔5z§g0D����#�3�\I�ʹ&(D�R��,D�`s%w,"jA���{�@�
vG&D�L)@�L��h��ߔDYZgK"D�� �B,>��� '�	��� ����l�cǅ��C�^pP��B?����"O( ��K�Aʬ��
S�.r�D�e��D{���R�zڮ�Z&���F��qR��Ul!�DV4�>�#;�L	��
�.Lj!���`�p9�H^�)�F1�A� _!�D� ;r��a��P�^�q��0@�!�
1��r��,��,�Wv��z���6|�l��&�H�R|u/,"�!��şf�Lmq#���xUs5��[�!����$˃%2�R� �^:.�!�*C�fy� ��;�t�{����D?���X8��!�E�6aK�Qb�C�-	�dy�H7D����B^1K�$��".2T�+0�4D�8���K&s�8Cw��3v��Cց3D���rg݀Y*�ȃ�&I=$ʾh{�cu��E{���P�C�� �,�>? ����,�!򤛩>� �)�OR+Y-��pq"@�\�!�Q�3L(�� ��{L���֔g��z�@�Aј�AKQ/-�4���J�n ��F�9ӣ��0>wD��uA@�A�V5��W�p�����:^���fm�DF����_w�I�& �v���!P��h��q��ת�!��I��կxz�чȓz�

�G�t�Y�\@�lՆȓ7JN�N�xLhCJSA��=�ȓ��ѢU�t���7)Єy��7��WhƠMwj�@�bB��*1��S�? \��叚���A���Z;�L�����x���Ʌ�o�Ę�<j�\���J��{�!��I�8�()��]��zd�D&Q{!�KXh�&��~?�`�P�=q!�DW�CL�Q �F�]3��;Ơ�-��6
O6-K�机�N`	"a��`W|%�"OzeR�(,I����ɓg¡�V"O�|��i�9n�򙻅FT:O�H��"OL�PEi��U�X����)s�F���"O9 �L"sU�ձ�K��p���	E8�؃�$!�&�C'h�;��%� D�C���7��"S94���!��h��F{��iĿ^w�@�f˼r�����,�0n*�{���:x� @�AnW�V:8j��Hc4!��8`>-q6�ΫF�(�S��["!���8�$��U-��?{\]�2ˁ !��_l�5�u�����aSj�~�O��=��l�1�ڈ ��q�V,�<�V99!"Oh�1AD�;x��9D��{G��"�U�lF{���#đ�4锜EPz��̫�!��{8��PD%;2��R�aY�jΑ���I!%�h�r�ˈJd�`e8ܖ�>�4�h��������#(���R�{7Daq�>��C��q�!o�I�P�sC	U4�1�ȓ*ނ�� �I��x��$Q�0��e�ȓ�
��@N� RTx�ş/o���$N4�7@U�r����	y�}�<��%I�A�<��!c���lH$�&T�L	����0�k��
X<�@tG%��ȟh�Ce�P�LH( s���L"���"O��e�M*_g0�����>x�I&"O���iۦ.-��(�$�(��A�"O<�9s�B�~E;�㌉m��(�x��'�N�0	V�fIV  ,8�pY�'��A��H_�C冈)��:.T�	�'&xrG��2ҞT��kȯ)P~�q	���yrO��eS��ED(2j�����9�ybE�Zd����a �+*�h@���y� ͽ���/��Ǡ@�N���ya9Yʶp	bG	����Pc���yF��$�F�Kġ�;E����L8�y���/x��-��Jl
��gC
��y�O�~���*�k�V����e��yB[���M�M1�z���L�0�y"�po꼹fƞ��4ěp�*�y��Vf�A�#��^�iP`���y"o� (f��q
܂F��
�-Г�y�iZ�7�@q�`Δ'�\D�@��y"&��(԰�`
�)�L*��?�y�t���V��

���%d�2�y2댝*{@`�A�%��I�D ��yR=tt=Bŧy���
'gL�y&��Y��Պ0H\&og�mS�!ͻ�y���?m�1
�J�
P�5ꅯ��yҨ	\̾�J��G����HZ6�y�)̺Ga����#�o'LA1G�y���uD��5�A�/:R��`�P8�yi�1c���c�*}��p{M�*�y)�*�_5~���W���y���#Ru����@�.t�l݀��2�y�`D��T1��DO�){7.H��y�#�:_(��ۡ�R�;�n�6��-�y�	�>UH� U G�ɀ�.��y�!T/k���Y�f�)}�����߀�y
� f���lC�����.@<4H4��"OT԰��C�z�JMJ�M��I�Y�"O��(c`G-F��r4�͐h�|��"OL\��O�31A�����̾[.�� "O��!"� �d�pJ͚yB�` �"O�,��K�Jn��9��XJ�L !"ON\;uH
*#�~e8�$Q��N<�G"OHݸ���+����!���u"OH�S 
4~wJ����	\���"O�T�S��$k���@'��(}��� "On�CEH�5���p�_ �P��7"Or�Hs'�"'P�y�#��8'�Tu��"O�l;G&T�VR���GΉ �h4�T"O~�aA�M�Y�,ʗ��(��Q9�"O@��r�H��HSPEĕO��4K�"O�a��)T��%�cc�2 !4"O@�	�O��cKX���b�?q�&���"O~}I���P=K��aQ����"Oؐ�*ʕZ�HЩ`ڗO0�CB"O���B�n� I�~,S�;D��ڌc�p�`B7Ip�ֆ+D��hU94����NDK,�b+D�<@ � �\/��Ń�'^����'D������t\�#D�4}�b�&D��a��2	�^p��BP�.f���s�%D�0���f�z]�`)�o'�P�G/D�4pFBƙb� ���D/7TX�z��-D���G苕/���x�E�M]�@���*D��2�<|Dԡt(�! y)R#+D���4�,����FE$"${A&D�H;�_��ԭ�p㟤;���2�%D�4!�d�@4�G��?r�hA�T�'D��)K�`� 8��$�N�Zi��&D�� ��لh)�8�P.��Hv���G�1D�|r�C�od躣(�Il���/1D����I:�|+Wf
:�c��-D�D�Dos�x�gܺs�(��s�9D�,��K�G8�ܱ�䗝lXk�"D�x�6ǝ�.�&@��OT5lBP��6D�,#ŊÒ=���P(�;9��: `3D����A9N�ڙ9Fk�s���	tI0D��q��2"֩h�C�D��� �+D�P�WBQyx�01&�!�dE���)D��X0�I�ӆ�� l�*�l�D�!D��z���A��"C w�8*�?D��s��'h��P�0#��D=p��%�+D��bq�C�E�!����rF8� �3D��f�YW�� ,ի:���2D��#Mϔx���G�5� ����P��y"�X�suv\uN�/{eF�hL���y���6Q^���"U�L0	�D�yk�.d����5)�jH�e���y�'Ԉ7tH��ӣ�vB)aUm��yBS;z������G��[�$U�'Z��84dY�2��ܺ�V�W���'�pӳ(�lx�+� 2M(	��'yf{4N��ph�b5 P�W���'�Rc������F��Dh�
�'%kr'�%bH�s�Z�I��,+
�'ݼ���a�)6x��9fOѵF1@@��'�%8��L�IX� �
�?r�'.�4�@�ȱ9䚜Ƞb��h�~���'$�afU�,��՚��\ 0N��'4n4�� N�6�p ��G�[*�}J	��� ��c�j6;�,�2��D�����"O�	1
�H�DD�g�E����%"O�,�q��*Ve����*�6P��"O\��sm'*��E��԰m����"O�I�7�֠oR<(t'T������"O�jcC�7 50`�>�:��"O�i[3�*
�qK#ꇎ\qh��"O�I����� r!�G��"7BAa�"O�r����yu�p��č�\���v"O����b`�� 	W��X�"O�$aub�_͢�j1Ѳ0�T��"O�x���1kbD�`�_�*�Ƭr�"O̫$�Q+x��`nV�^�6EqC"Od��ȍ(��]�5�XDO���"O��0b�p��Т��(B6!�*O�q� oAu�NYe�^.���'��h���'C
T�+�t�H��'l�������]�zE�C�R���
�',t�f[tb�S�D-	$�#�'��<0 ��d�,����|J�
�'.$ՃE��K��#C����T#
�'O���B,��{�BY�"#P5  0�#�'�>4��_8H�l43�#ɂxvZ1C�'�
�y�B�
@'��cu�Bq���'�H��٦	�tt:P��a��)��'�,��@ N�
Q����H:�x�'�(9�	�ka�tI���?_N�c�'t���!C	�fh!�G O0>���'z�{�f�%M:*հdF��$N��R�'Ar!3�l�\��ڣ-�d��[
�'���C!d���~%	��V�^|,MI
�'�x�UN�.]L x��l�F�I�	�'���)�����F0Y"O������'ȠTZ�c+���"�}�hu��'}�Sw�B|HfX��n�K�h5��'%Fi�t�.}��Z�`<J�5��'ԩ�sX;<7�H�qEU,5҄y�'Z^��c�0<(��%��4�4��E�<a2䜑'�px���Ȫ{�	"(K@�<ـJ0h��"_�)��(�#��{�<	�c�0a���3���?$@�tQbG R�<��Bκ>�H�SfiB�!A��F�h�<y�@#<��(� � c�|8����g�<�v��.S�L��䈗����c�^n�<���+7�0��]A��	E�F5�DC�	�5�	��@"F�>�b
��3�TC�I{�B�`4T�����`xDC�	Y�؉q&g�,��"�V�QT�B䉍U��zgO����IɨB�	�*�*�)�"�%X`h��ʞ'��B䉠r}�}��'Cy�.��"�${6�B�)NE��a���8�ɔ��XB�ɷzX*�j��4��Huӆ�tC��X�2hI5K�y���ЄI�C�	��B, D�� ���¤#�zC�;L���DCP�+Py��HRB�ɎL�����MB<o�������ѺB��C3�EK��J�3$�)R0����B�	)1�v`qw[
��Q�KʈJz�B�IG}��pA�K(P�S/�6�B�	�b��[�*�4��h�˃~$B��)o��8��V"+
m8 '�
rFTB�ɺ[
�C�`Y08��Pt��4B�	�s1�B˘k�@����e^�C�)� L�r�]�wF8	q���&�|�V"O�0P�'<F��d���L×"OXL3�D�$к9!�H�Iz<�@�"Ob�
�Ȏ�?V4n�xJ�8�"O������g�Π�s�L9���:"On�P@D�$6���ؒˁ/g,L
�"OƸ ���QGH�2,	:��1��"OI��gG�`�,i5� -hl݀�"O���`DB�w\`Q:!��&e�e�'"O�|�2`\�s
�����?v�=A"Oʵ�b��]���;!��%0L2�"O<Y�p�X?�,�v C;}��H)&"O��@IY!.5`��oK9�	��"O�8q���Kt�se(Z2���Z"O\��7]��D��R��K�:B�"O1���:K�"up�e�m���c�"O��׆	k\�Y�$��%���Ƀ"O@y�Gd��c��@����<�Й�"OZ��w�� �v���$@�F9`혡"O��W�H�$�t 7���=<\9�"O���%*�?�J �PdZbZ6��"O�0b���/�x��⎗2Z���"OZ<hCD��7e@�ٖ�5$Y�2p"O����#d�̝�%~*VERe"O������@%�q���FY�0:t"O�P�W�Rs0Y �Z�7r(�q"O.jp/ؙ16� ����0��'"O�@�e;ZDl �Ck��D��"O�Q��ͯY3��۔	Jnk��B�"O��!+]�*�Xc����N{~��"O��Hd�(K�PJ�hY��ɴ"O���o�S� Qq�P!y�d3�"O.D#F�J�x�Y�ף�azI��"OJMг�-��d{�cM23)\�B6"O܍ɀ@�W�����k'>]k�"O��8w�4Q�L�E�@ `h�"O��A�i�߶ I�D,#�RY2�"O���t��g�(�Pv���\q>)�W"O���㧌�cה��`�СW�4�S�"O��#2,úG��X؄ I<F��H�"OhAפ�?ibtd��φG]�|�"O��+�"\J��q���4@B���"O�pc�A�08�|��v���4:,u��"O�Q��i:q��$�'Õ�Q��9��"O��EiQ s{��X��_�J{�8�"Oh*�e�k��!j4�13cЙPE"O�i��b�)(��j�C����3�"OƜ0���d�έCA�A�L�$-V"O�m�P-A/7L�q{V<�P`A"O� Â�ɀ/+�M�F��5����W"Ox�[�����ք!�쟅X��Rb"O�;��}>L�{��-{���p�"O�q���F���arE�K��M
'"O����K������:=�����"O|M���:o�05;�M�p����s"O8�㠮�3v ^{�BIs�P"Or�y�/
~��}��$B3>�̘e"O,��t�JKk��@����*D�^j�<Qqi6�������#r�ډ��Ia�<�f�Z�3�ux  �g`���EV`�<���A2t(�"�v��x�m�[�<���D��E��4�0q� �_�<a,ҊI��Z+U���Y�e�<��J�=
^�H�.��k�
Yv�<� ���'�|�z��s���j�9�"O��磅9x"0��0�%�����"O�4�w�|�����X��C"O��Q�g8�`�E�'���S"O��ʇ��"����$U5~ ���"O��0�ǓZQpr��9@��X�"O ����L@K$c�HW�}"�"O���0�4" x��K�jS<đ2"O&I��ՌC��<�DȘ;GPT�"O��ҁX����hӝc?Z(�"O��+EÇ?�@�g��<0!d"O����a����Es���	5Hh2"Oh	Dj�
Sځ֋��=�.(�D"O\I��@y�j �a͈� ʲ	0"O��P��Q�:�d�i��";�0��"O2��̀{�8=���	r�\��"OX,)1�ܓ��	�'�ʮ!���+�"O�9���:��1k'���{�ui�"O�ų�N��g���g�61X���"O2�ѧ���y툸�$���IJ��D"O���n��z�T�Q�x�V"O�����ܣ"�j,d ���.p)�"ON�y���.n#�,����U���a�"O~�Z���Y���)P͏�M�~�H�"O�:�Y��M�tL�*i��0�4"O*)��ΛP.�!���*o $8��"OfX8�CZ1P�2-)阠4H�l1"O"P
�.r�؊QH_�V3���"ODq� �]�lA��@�1AT��&"O�|�Sf%`�y3��/	�[�"O4%���v�.�鲫�L�"OFDRS���Br����䀢բ�""Oj܈�A�&cX���Ǻu�h	��"OB ��U2&1.�ӕ�F,%�\I��"O 9G��9,�d���+˵J4�JU"O��RV>���!�HJ�."�"O���%]�C)�TA޾]��q��"Of��gm�f��E��`�w�帓"O�ٱQ$�_"^�n�[T9��"O���P���y����ж\P���5"O,�H� �8���u��;x<�pV"O�!�D΃+4�8�``5�ek�"O�i�w��t0�$��5�a"Oh�C��ݬ~��պ ��?��e��"Od�"p%�� ��	��P�	�4��5"OX1���Lڢ`�F'ͭK�J��"O��&�%Z)�t�5�ߣ}{��t"O���P�ܐL��q(��ʂ
ю�%"O���#Q��% �FX, &�m(�"O�9!�͑�&�j�K��#��<�&"O���A��#;9X� V�	~�D���"O\tÑ��;S�BëK�b�@y��"O\U�@۝w�����K&U�<��"O�HS��*bh%�@�ٯ_}���@"O|��_2"b!�1��a�U#6"Oj���Bե>Z��W�dO
��5"Otȳ�C����p�(��t��}�"OȀ��+�yLh�@Ü	A�ebF"O�(��]�m��pҊũQ#D<"Oı���	�2� *��|^� "O�X����A|p��#���Q
�@�"OX�q�x����� 4ੲ�"O@�k�13��9��H�o����"O��Hus�M�uǃ�m��ms"O� �p�u���	�:��G��,����"O`tR��_�4Ԁ�ґDQ a�@x��"O��a�D-k8Y2�hP�7����a"O�X�O����(3�N�\��eK�"O<����Hz_�h�6FG�ƁC�"O$�ʱ�De9Ԭ��Í�fZv�*�"O�<"��Hl0�����A�Q�l"�"Ol Hr�.R3r���֌sB�Z1"O��B�-�`e���֮�
�A4"O�& ة�Ơ*�P2���z�"Oz9w�&nWPY�$^3J�����"O�Tyv ��.[
i��҄�Dو!"O�8�B43����(Q%L��d�6"O�آB�ǯyh��AG�ԕ9^�e��"O��[���3)4���%�6e摉�"O��#�mHq���nP�\H���"O&�+F��P���H.��}ۊ �"O�U��ߚ~�4�5- �.���"OvP�ҫޮd�)��~�,	��"O8 	G�5(o�"%��<���"O�P2uO-.,�}@���6�Ȝ��"O��jT�ʠ;A��R噷e}z �"O���c�K�o|���B�|F�!"O.e�R.�=`#ڽ 򋕗��c�"O�1P��[Bqza�G�P��`��"O���b�>	�ü8�@(�A"Oq��N��#v-յ@�0�hW"O�5�A�#7l8I3�L_I^\dc�"O,�B�-EUm�q��@�qb�"OQׯ |8�e�	���"O.M`ïK�'x����Aڜ� "O�)��	Ib�.�x ݱ,��a"O^���0\�ycrO�2��2�"O:�Z	�� ��ŷ ��<�5oi�<�3�Аv�d�weU%�]��+�o�<ѥ���Y8pU�W�Ҋc�T\�V��g�<�r, `�6a�CAf�e9��Sf�<��K?=ꞹ	�����Y9l�b�<���ܘ�nx��茆E�����[�<i���N�`p0�ܨ}�i7��c�<I�dY 17���Φk��PzU��E�<9 ��h���A�&_b���C�<q���*Ѵ9:��P�'Qj�9d�AA�<�լ�,>���� 	>d��uH�<�^�~Y�:w�ٹhD�t�P�k�<��H*J�P��j�1ed�ܻU��m�<�aC8[��9j��۫'��P�L_�<�&N/"�r����&Z���;��UQ�<Q��K3�������J��CqJ�X�<����?�)bA*V\�P�K���~�<�뎏D$v5��&L*cV��%�a�<�G�r��H�m�[�d���,!s!�D�'QsRq1F��=z
��F�6Y;!�dvU�#Eg�a����%mL`�-�ȓ=0�A�톪7Rrap[�[C�@��F�"W���a�cW�D!T(`Q�4D��@����!�fA8�j��?���(�d D�48�IO�MJ��Q-��0 "]�s%=D�xq�
Y�����'(���b,O�<�6E��.TMW�Œ)��y� �U�<��ʃ!3z�r��G����&݀�ȓέT�UeA�(KF��t�lY�\��6�l�bEF�Xh&�`�P��2�ȓw64 : �&Bv��XC-���Y��S�? ��Qc��J���(�JM"��( "O��rǅR �X�P6 :$"Fp�A"O��B�ن�t��$���؅�a"O(�k�]#Y�4�)��C5;�Pc�"Ot��Wd�N��|�R��r�ј�"Om�Ef�0	�MgdR�f�H�"O��(�`)OĠ8X���=���"O�A� zJ\�Rc���>%�O�<A���C����@*	� MH(��Tb�<�D:u|���G�c���P% N\�<i���4B�h��-�K�2�"D�b�<��ʹ-�`M�G�y�P�Rv��X�<)f U�����fP&�P��%�PT�<�˕}������F#�rR�P�<QD���{��)y�D˗Xf�qJG�WN�<Y1�Mƺ�c���M8 �h"�S�<��K	17l0���a�n��^h�<���?ǚ�H!c��X�lD��Sc�<1g!΁(�N��po��*��僐�b�<!X���pF� ;�L!�#�7,����_��S��_+w���H��5��5��~8��3W$�8XP �ƥ��ȓff`B��F��<H��+
A�$��XO�YW��A"h���c�/
��ȓN���N��\���P�+�`����3c�J������=w�!�ȓN\���c#Voέ��M�!����
줅ӐkL� ���kJ�|���ȓ��:jx�a��oy��էl�<��.�,x{0U)�Ƒ,\7m
fM�Q�<	��@�hf��k!��-~����R�<ɃL�o-d��[>7h���V�Su�<�&��=f�|}x�{\�`x���j�<1qG)�"� ���\p� ��|�<yEM?G����Ugj��c��w�<Yr�
�Pz^�Ap������q�<)�K
�Q�\`��jI0��ċ&�X�<	U"�'xA�Aѩ������R�<i�N�"U�u��n^�m�<�8C)�Q�<�*)8��i�W�T�jC��M�~B䉆��b2�Ґli���:rHB䉷4[��0��S&	]�l���B.i��B�I�I�X��A@�C������=M�C�I4O�A"cK�0�v5��اC,C�I�^m���ÁäKj�¦���\[<B��-l&�* 
�2e�H���L�.B�	5��A�D�l�ЁcMh�jB�ɶ'IV1H�jG�*8�=���LXdB䉬U�j�Q�2�~���j�s"xC䉂l?��Fo�H�(�pf�,~rLC䉷'��Ds`����
ہ:y�C�I�'��u�0�Ҭe���C����C�Im�`!����^R�,��Eըi�B�	�	��k#,z��j����Z�B䉣&N�x�U��ɔ�1��C䉴:=���r�O^P�*��8G��C�	$4$��"R7L-�Q�.��C剢Đ��� ���k��
,�!��׬on�����\-�5F�T!�@�u	ᩌ�)r)���A5!��i��ؓp�H2x��i� A,!�;c��' �	:��t�O�v�!�Um �ႫmʲQÁe�*j�!�D]�<��!3��
�Zx6�Ԯ\�!�� �d��/�?)�\���M�9�rT� "O�h�t/��.U�C&��^���"O�YKg�م^���B$'�<�4�s"O��w�	-�2������R6Ѡ"O�`�A��1f��q��[#�d��U"O�H�A� @3���R�[������"O�`0O?�F��P&�
s�N��"O:�r�FMW:� C��/J*�K�"Oڨ�pJ[q���BT� �p��"O�(��J�_W2Т����lwd���"OLa��\1#ĉ�7�Z�+n����"OVy�oL;��ehX8~�V��"On�Ȣ��_��H���VL|�!"O�h���;z�E@��S۔Yp�"OV]*��'�X<1�O�_�j�@1"O�Ա��¡�Jy`'iX�{,�""O�PHWHX K��Q���)�<��"O����(��T�D�@�I*F~�I�7"OqRnU��kB�/v��["O�����A�nDQ�e�Ti6"O�DP3�f3� ��!�Ak�]:��"D��6B�3�N����Hd�A�a�4D�8B2K�LE6n�-�xyw�.D�,�eJ�#=VD8��F:����+.D��� .�W/���A�L���G�+D��R�E۴v��*r�����K��3D�ЁaFӔf��U
�fZ�Xk�=�#�-D�31	��0�d�з�Y�=e�,D��"���
�����/��p=7�(D�� ����q�+.�%!D�aS���T�f��$/���c��>D���h���ظ��X=�Tڒ�;D�Ը��	�
�������Qz�a�+,D��rb��r�� Z���*�^��&a+D����ԪG�!�!-O��
��'D�����&��=(Wk�"Ͷ��r�$D��q��B��$A��%��t��EH�!D���
�8J�c-����"D����H�Z�Թ*�i[�1`]�'&D���w��&�\TV�˽6H�an8D�X�*�;6Z��q�I�vz��ZA&!D�z`��7Og��1�-_l����#>D����F�?LR3���L�h!ڣL<D�|Brㄦ1���Ѕ ��&B9�C-&D���`��%�>`1���9� 9��(?D�$ٴ@�o&�U/� <��e�1D���`��0���"���p0�`.D�r��>F+�4��'�	p`Q�(8D�\+ҡL�v���
>sI���Ƅ;D���mۏif����G|�*��K-D�D҃����\�Z`Nؠ�a�� ,D��*#���\��]�e�V�5�R*D�8@���,����eh-��Qwh(D�����
S��0��иxT�;T�'D����F�q��3�d�?;z��'&D���'.�v|��"cd�~��|1h#D�\b��!��q3ŏE)R�<��P�?D�Dk%�ڃ ���ߤ,!*K�H?D� h�D�/jҤSu
P� D�� �"D��C�GA"$�d���bH3g��+��<D���P�"�yb*��`@�4�;D�tKekN�[� �(2��a�V�i$B:D�xP�j��&�:���e� ��ah7D���C*��3�`��s�Ɩ-X��'�5D�� �Y"�I��w�x��┮s�)�"O�����@�(Ŕ-ⵇ#o�zِ�"O����ܘ^NQHw�^�B�|��"O, �r�2<�6�G� �J	�"Opa E�F88�.P��L��'� �A"O�}ۀ�A�\�cԫљ4��}ZT"Or��Co�>GQd��2�4�FI˥"OJ��LD��=i%��T��m�s"O>Iqa�]�Iz$��j��-P�"Odq+n��Z�A�䀇E�D- g"Ox��b�r��#ƂK�ؘ�"OtPA ��y8��w+Ӌ/x6�;�"O�E�Ɛ��r�%zs��#"O���"��ʡ2d,��cd�y��"O�`��<��ڶ�X�tyXC"O⠋�MO~��b�ꇹWC�YT"O��[r)�k;�X�䆓�0����"O���� �H��4O��Uf�Y�g"O�XD�Vs��i��.SPD��"Odl���0{T}��H	^=�uCc"OH�P��%/����d���Ih1"O�8�֧/Dz[ P�L�
�1W"O|9դ�%��y��������rB"OJD�����W\x�S;Tn,3�"O$�@!협`{R]q�ƍ�gf�"�"OXȆ�52\����ȸX+8p	f"OP��7-�2@-�P(��C#~��"O��#A
W�{�d-���"v��R"O��i�e_TVZUPsdݳ�v�"O^���+� >0"C�o�l6"ORPZ�[x����F�Q8_�t2W"O&9� ��d"B-��j��3�n���"O�qr�NϘu�*U7'�1��8Bu"O�ˣ��:Q�8��PިA
�+$"O"T1��^<%�m`�ƈi�ا"O�y�ۭ=�E1f	$,c< b"ODP��{FDI�.(v|��"O�p
D!Q�	��5�+^�5�>��"O�Q��Cs�F�Ie)Ŋ!{�5�"OL�A�B4Ud�h�V�Tsd���"O��K�A�/Z�9 ��,��5��"O$p�
�1`.@	�jG!vЩpq"O|@B@�s(~�g��xbH5ؕ"O��3�[4O殬�4��s�:�q�"O���)���3$��'�t`��"OV��P
]���2�"�:��2"O>�@��*_kT)�VB«~V)0�"O�xCtLF�4�:1�[�C��уb"O����eئg�HE2T�|��81"OpDs�M�,-Κ�z�-Q?H��U�t"O���M�/p���0�a��d;�"O��v`V3@ `J�L�C�D(�d"OBL;�K[�>2xR�j��Z�� "ORYgQPD�x�T�1��"O*�;��\
'�&l)wH؞)i�@P�"O����� afi�%�%@F��6"OP�@�O�� ���P�@���S"O@Șf	 ?���&��Q�%��"O��1SÑ�R�� B�W��ě�"OJăԄ�=�T��3+ʶH�"O,��a��q�d�S1��.Z�4���"O�(�6ϯVz���eG��Pz8ӥ"O� ÂLm2P��B�_3�P!v"O�yIK[1h�jmx�V�s���6"O� jLסыO��Q��+��m��"OJ�Ac���~�y�	�v�SD"O��!N4-E�y���%I�M�r"O�d�s�*6rzI�� �,>&XZ&"O`<��T	?b���.��b��ȱ�"O�I��^�I	��@�?	zp�6"Oh����
W�1�#eS)As����"O�e+Q*�|(�(��Ka�08�"O�PS�(������V���p"O��'��.-��(���!��"O��qd�b?�0�㖲r����0"O4��c�Ҭ d��v!��6�Z	�"OJ�js��/+$��6:φ���"O�<�F���@Z��H/�h���"O�}�'��w�|ArU�Y n�\�!�"Ohi����!Y~j��ǤV�V����"O��`��JW
|� �Q�~H�Q�0"Oލ���ס]��q3�`��Nx�2�"O�H�riJ�9,0R��B�q.����"Ot�ɦ��Q=�rV��^�0U��"O���7-�^����!�AQhTD"O ��v)՜c�v��'9Y�E��"O����<\����� d=&�[s"Ox�P�I�/Π�p�
�+6�U8�"O��0-�v���#8$�\�"O�X��l��|��e�փ�� ��L��"O֬�S*�=5f�Y��⋧Y�v�!"O��C��o�2�a�����1�"O`�'�H
���i���6u��̋�"O~�gȟ�T x�
�.�$x@ "O����E�D���%N�,���"OT	��kW�i��y�S��"���"O����*;	���I��92�vi	"OQ��O�X3��9T��X��d�c"O�<u��-��h�E��3�¨�r"OXU�'	�V�A8E�6�ոS"Oj$�&�'i��IB���(=B��@`"OB�"Z"���R��'�yb�"OL�����c�t�3�"�m��y�"O&�"6���tVH�b��t"O�P�q�6�����7x�z��"O���`Ȉ�+�H�3��a)�"Oܽ��/��MKC&Ɇ\�� 0"O0uj�5����v��A2�$ZV"O(�x��M)>���k�$r(�"O6����v���z���Yf�`"O��sw�ӷ	�~LJW�	�kHly�5"OبKA� UU:q��(�)�x�1"O���U����v����B��=#�'Ht�0$���l�CF"�j��A��'���"A�N7"��ѥ
ܳL�E(	�''@��q���ʛ�l�`s q�G$D����EX�GJ�"��4�,D����q	>L['F�A�\�>D��`A�7n�=�R���H)z���>D��Y&H�f���@֬v�LU��/D�|����8z @��]O���!,D��"�(�)(�`����ͽ#���q�,D�t�Q"ǕE(��t$NȬ �C�6D��+W���(����[U��*wf/D��7�3>�B\x��=�dT�B�+D��ţƇ���醫̵w����a!.D� 阞h���'C��P`��-D� �"#-0���C�	�"������(D�� �T�5��.[|�$�E?2��"O�0x��@�b:Ĺ	3ͺ.ϸ��S"OJ����(�7���yt��&�.D�@�N+5i(�
��X(%�L9���+D��zQ�^�ϖ�C��S�|��)D��b��k���#�щU�<I�'(D��8�#@�\����`�`�"D�,:��āc)*�)�m	�~�&@j�,D��`�[/l!@*�̂�X��R�� D��s��6 �D���n�;�
� `E#D�\��ƞ^t��TCH�k(� s�$D��KE�M�`p-�c�Z�:e�U5�!D� �Gc�t՚X��m�8
�����<D��
�a�3Ae�ib�D��s�}I�j9D���##6tJd��)�[ў�r�*D��+PO�S�а��}�@A��5D�D��̯�б�E�8�8�e�4D����֟i�F�	ƃz+H1�� 5D���p�ŧ=|�r�$=��#R�.D�DBD�?��$�d��� �S�*D�p+�nS]t�b�͎H�9�D�<D�l��.٫8�LE.�s���kvF?D��`#�*4����AՒ��a>D� �#��@'H�w��85�I�eI<D����,�t!��	�җ1A:Icr�,D�p�5���.3���]�.MЕ'D��ch�|@�L2eϑ!�ڝ��(D� ��I>>��P�0O,p݊4��,!D���む6;@�)��)�
�zjË)D�T#�c׹3^0hVO
54D�s%D����L:bR��
���q1!�XCWrC�b܄,;�h	E���9!�Q(!�Ȝ� �R/��Q��I�
!���w�-� 	q���[�	�
!���t���n׏*�X)A��'q�!�׮?�,K�m�KlPf�R!�DE7c��0�$��$Z���"��@!�dE|69���?L���f׊Z�!��j�
���n��c�������!��Ʌc����%�?&Ξ�a��>p�!�]&*`���Mד#����(5�!��iI�̋�aZX��Y�Wß
�!��<1ޱ�
�#%��̂#�P3`&!��;"m��s���)�\�S��ѐA�!� >i�T)X"��t��ȡ��7!�D[�+�z%����hb���9l�!�Dʤ��Pt)�,gD�e�C��
'�!�D 
~֥��o�7A&RelW:k�!��֗I����A��^	��*���>!�D_*	D�at��9)������!��T�gv"��n/u���BCs�!�ݎ��X��H%/r@U�4"ԬH�!�D;x�]�$Đ�[��y���N�!�زU�Z�H��WRNr�I	͜#�!������K�ϒ�g *��N!�$D�vS.�@���g�q�/�!���.X`����ؘ8B�M�c�q�!�$O�O�D�'��h9>�F�"Xl!��Y,6ќ�A�%�8,6�Y
��^�"Q!�d̃t���`E�S�#w�)���S�K!�O�%z�����sb����	x!�G�C�M���ΝK�*��*��!򄐴t|
4�B�C#P�P�p�[!2�!�N�*��y�F��Z��}yrH�L<!�� ����1tv����f6�х"O����
u�Y�ƅ$l���cF"Od�S+��@(�5��d�����s"O�pA0��'&a0D-c�2d�!"O.��@^�(�T�Shѵ8:`��v"O����<T��	æ��NW���D"O`B�Y,tؠD�ᢟ�U��a�"O��a'ƚ$T6�I��-j?�x�"O�ɣ����R�ⵁ>/pH �"O
�)�*3��Q��˔r�k�"O挻�3v�ȍC���Y�0r"OPd���F�'�s�*X�(���#"Oj�H��6����Q(�n��"O���tk�.cÀ0������K#"OX����Q�4y6��*^���p�"O
��BIh.�Q�dK�7��\rR"O����Mǀ)Q�_
B�\���"Ox��	.UH�U�L�$���2�"O,̠�$ԫ2�.0�A��9*�""O��{��E���H��Ɇ�r��ر�"Oh	�1�A�51�ș5�J���"O�����H>:�#�'�5w�͡ "Od�k��΍<����S%ō+>��б"O��X�!�&��1X��Dd(��b"O�U��a�`OH!�G�?Jћ&"O�Ÿw@��B0qaDa�.�^(�"Oh5"$DJ.V��	fφ?��H"O��⧭Y�;C��ʣM�-�4�"O!P���r7�br�+����r"ON�bV�DG5L��ě&e����*O2<���5� �`!��64d�X��'�褀�½e�*Ix�+K43;K�'B~�c�!۳m��]R���%�
�'gv���K�Ʈa���K��x�'�,��1(�����c,�}*���6T$봄��TK�AyS��67��ȓ?U�����V�>l����tx"�ȓ��$���7��!8G�F%*�4�ȓ?k�Zg��G����
�#�6q�ȓhԂ� ���K�d��Ƨќi�a��.�@�@� ��f����Z^yP���K�X�3��V��h�BD� ��|�ȓz6�`�3*G�ibf0��	��FT��'!J��#A�3bh1W+W%m���	�'.d����*6��Tbso���� ��'(J4��$N�Wgd��q��2�
�'�0�b�a�w8.�c�Ջxz
�
�'���A�G)xv��E*e�8��'��t�_�]1�H@�X�����'���82�4�Bi��T�x$3�'J��x��V�pN�  2.��kܖy�'b�-A��k#���A']fb����'S�u1A��)o�� �b�)'v�r�'  ���%6�����'���'R����6��Xq,�U����'��­59�tC��4Q� �H�'��p%#�"&@Q@�F�|.p���'s���ҡ�>#�h��G� ژXs�'l0����Ę8*�PS���0}�!��'��	�Q"īYNPKG��!�D*�'���)�Ų�RQ��Q�m7��
�'�t���\$h��1Z���S��Y�
�'�4y�Տ�9��A��^�N|	��'�μ��m�0=k��h�%�(?�y���� ,�Jj�&T�ȫ�'M�ZBF};�*O�y��nO)y^��3j�=@@l��'Z�a�%۔>��y���#p�%i�'���� �%	����!JϨb:�e��'+�H��.���2c�gû��Y��'�2@�Vb�<�����-�l�
�'j(�QE�&r�*p�J2V��ɨ
�'�~��cȚFM�	ŌR0 �&�:�')�t:g����rȺ��n�L�	�'R�{T!��/.�����_�f��P	�'���kE#[9���ǁ6b��8b�'
J$�����^h�� �R��}#
�'����T�L84��bq�Hr^��	�'r��Am��x�Q�SxP ��'Ј`��GI�|�9�S!ޞm�hs�'�5�S�ʝQT0�R�Y�7�@-3�'�ڵ�`oޚ,�܉ @_00�	i�'�4�2�M\�hr�YKD�Q# �
�'��G",�.ɩ��M�(�
�'` �1MѹQ�j��ē����
�'� ����;ϤٚRI�9w:��z
�',@]1 Z�!���� $ ��j�'�Jl���/Dv�!��ڄp�l͘	�'�X��"K+�.�׀�
}�|%��'P
<��iïG��z�N5q�JQ��'�u�����,/,���_@����'�2��L��>"Tj�eؽ��'I��6d���,�0�Ϣ�!�'���ȰK�,9,�-��I�d횹��'=@d�W��
%���Ԣ��D&�'�`�+aAC
=�0���J�|�Xy�'���1��@Z�HEBL�y'F�K�'b�*�*-(�F%)�_�y�q�
�'�8�ECסS�Z4 �w�((a�'R�¦@�)�ة�2�Fk����'�$q��[-..C�m�#0�ҁ��'�T��W! �,����_�";���'�n�;`DXY?V��g����(�'�
�X1� �q�y����I�'��rT삄3�n�ǫ@}adHB�'{z�*Co��(����zm��`�'�$=�G�E�'�J"��|�5�
�'����[�|�Ac�z�|�K
�'�<��KI J�1����)	霍B
�'=�5���ox�qJ���E�	�'j �*��ۿn��y�TH�+J��	�'ʊ�RR�	�<b6u!M�Jp	�'ؐ �&#_�J>Z�0e�$`�%��'1��f��y�|��Ԡ�+	T��:�'Ά���Ԏ9��d��!%��S�'%&4�dG:H��\j��2����'�Ą����1O�1�3�F6�9�'A��rE��4H����#\��Lx�'���A��d�����.�5�hQ�
�'����i'B��d��pM����'i a���N�V;��)5♔d�{�'{*=��M�n�X�k�aƟ\9�0��' zj��_�CV��	%����uY�'h�����=z�P�f�&U�J�@�'�а��	�h=Д!yT�u�	�'i�)EK�#Ic�L:�L֡Aݜ�	�'� qs�ӱ*��)#�A����	�'�T٩2퟿Y%�ZV� 2a�թ
�'�� �i��^��C,3���	��� �!8�C2cn���n�.7���"O��Cg�V��Ƞ�7��#�"O�%xs�>`�K�i�/��H�"O��W��hL�)�Ɔ��U23"O�+!�Y�kpq���!���S"O���c-����-�q`��D�B9��"O)�M?o�P�y3BϺc�x1��'�|���.2�Q׮�+m����'Uf� $�E#"f!�WNN�M�]{�'Ehq+ËK�FD�
�Ǔ�Ki��A�'�!��p��S3�tN\][�'G��`�K>n�p(2�f� 5"\��'t��YW7Є:���X��'�t�C�^��܌�>H�"*O����W�p�|cņ� $u@���'v"X�.�l�b�t�����m)�'	V(��S�,:���4$D�Y��Q�'g|	0L�L0AzdJИ~�&p�'����BC)9��ɡ�bĠp7D<��'��� �	�)}�	����=3�����'9�Uz�"׮[<����˃�*w�}�	�'m��2&
0$X�C�%��d��'����7㜑i����JH�"��<��'vԥ�e+I /Zv �4��&�Ay�'�Z�(�E��ذ����P��'�f��S�!�t0�d7�f�P�'l���CO%(���`C�F�9	�'߆t*�נX�~����&�Hq��'j�e�!&M�u$��y!AJ4qlް��'�(��&�3�<YA�'ؕ7�F�z�'���A��]ɅkX�D�\�8
�'/�t����@w
����7n��$�	�'a�ɦ��
:��D��By$ "�'B� ��$��+���X��Ր
�'�x��JJ��dW���
�'����ȒJ��%
��9_��L�	�'�Ҝj0��.{���!G>R�THA	�'�E�Q��z ,ї�]P2��K�'�&��cR�_���v(E�[R.���'�$������T�x��FV�<d �'F^��e�x�@AkG8WK1
�'��y��B,x�d���?W�.4Q�'�A��C'M�
�qCѐBM�)3�'EHٙ�X�U�>�Aq�=��]��'n�aP4��!(B��#��2.��@�
�'�� �@!��0N��ɣÇ'�0�
�'ߤ�z��2�r���!W�%��)	�'4\�0Ea�)W�%bn�-h�1�'�rx)��BIڐ@AAز%�rQ�
�'q6���R�v�Ȥ!�`_�3D��
�'ل��IؠvĨL� ��+HPS�' X��Q�eH�7M�0G����"O���T�/t�X��C��g�$��"O`�$A-� m����� ai"O�`���ǜ@�l�� &�'!�Ѥ"O�� �
�1r�*I��$[�!��rg"O(թj��Qh��փ�Wh*��C"Otı5���E��`������r�"O���7*8�N�Jg��	sǸ]a�"O ��CFy�L�5�;��hs"O�TC �׿Q��-9�&��L�H\��"O���ALLL��!wEZ*ǤP�%"O8ݪ�C�1:\S�DQ�
I�hJ�"O�4�g�
$,�> a�\�uE�l�q"O� ����Y�k�pe �D�'m=���"O��L[�8l�R���Ǩ�˧"OT�P�b�@`U3���f�� � "On�Q��O�]���x�`�>d���"O(�a�C3�8 �S��3 l�Z3V��E{��I��V�ڄIƂ�5��8�F$C!��W6E�)��e�9��}����t*!�D�=`h͸D�M|-�Ũ]�4!�A�Bt�� �N�~1�b&��!5�!�8/��4`��0vҢ��2n!�ԋ5Vh������"�]B��Dg!�ę
�t��0m_�xkP|�M��c!�$V�L�^,�ro�M4	
ի�I[!�d�r^���o[,1%x�ʆ>W��`؟��0a��?�h���'�<{Z	�Ce��G{��I���^X$A��؀���X"*�܄�-�\��х~R���*ùE�Ƥ�ȓ_�ّP�E=N�
`@3��*_�*M�ȓwW�H�w�]��R���ݨt	����HO$	L��'�fو���r�z�sw�1r�1�'��� �͎W�X�Y'�K�gΤA{
�'8q{�a����t�eGҺ[K�U
�'� �� � [�Ĝ�E���T��a@�-��OX��˦o_�xӒ���k>��H"E!}b�Rb�(Z�ǆ:[���ʧD��'H�#U!�O���McP�[�D��RE0q���"���<������*�ɀ�̉Qg6�#a���Z�p9Ju�I�<����O���!p/P�gǜA@�w�"@2/O�m��O,O�g~B�!|@�"2��e������������\�W�{��Ӱh�r8 GR�o�+Х%~�JC�IP��Qk+�G�H��99� O��	O��0*4K�
l��O[�?K�) 'A0����6/�h�K�͏�o$H�i�旛�l� �W�'�Ĉ��U\^z���`��P�&oX�<Dy�B%�`�S�GRd�.����ְ�?i�
Vo��LP$֚$dpTp2���u| ��>)��&�S�$�x�G��>!@1a�^VpY�@���~�,ғ�HO��x��ӗ1
�8�[e݊AB"O@�a�J�zA[	��M9,#cO~�����g�@""D�*�R���8��'*�|BN�i�R�� ��.���N�yB��;+Z�I�D�->�ne��%U�yB	�����k�KK/G|:a�mT-��O��~��឵�R��u$E6��b�M�<�t�ٵz����M �,�2uh�r�<�Cgϡ :����%sʵ�0h�p�&�d��hQ�Wd��щ�2rݾE���8LO"�d?�$J1`�)1Տ�$0�Pb�ƽ/����D{��H}��kA��lz7�@�'YZ�"O$���-�Q�T�cj��1��[��	w�OS`<��hՇA��Tcvp*�'a�1��a�����J�5���'`�Ç�n����N��c,��P�'N��G��@"64��.ϋ&�.eHZ�0=Q��䌖_�����L�2L�PS�ÎK[!�d��Z��5X�MM.I�<���lZ1O`0Fz��d.[�wbH�TCJ1
9�h��oϚ��>��O�p�u�]p^�BA ،0�q� \O@v!��.�L{5�\��X��"O�Т�@�\�bS� �Z(�u��"OL�x䅂�{P�`���ӳ|�,$�D<|O�h�f��p%8Wo�*$�`��"O�1BI�0\�Y!��"�(�
�"O��'��=����(|�r�:�"O� �����O�?�0����2��HF�IVx���w��G ��1gCCe�f���f�ԣ=E�ܴH�.Ձ!ҍhf$�u�,['
l�ȓw���`���`�Z�s�
��cM>��\�����U�B��ˡ�T$s�>�����0A���(ɫ��,5B���hO?Q�p���E���x�O�J���t�"��V���O6��k.8�\�Sc�ì�@�'?�u��/I�̲��ۗK��H��'���se�ߺ^"�9i%B0H��<��'���`4�!���+L�vX �Dѯ��>�OdX�Ղ�uX��V(�1'vW�y�b�=�x}�� 00��H@�9՘'�ў�'�|rR/8u��� %�)nƸ1�!�2lO➸ѥC��L�!��K/u}~��/2D��Z� �N�`qJ� �)�\I�D�0��p<����<!�>���A,y# �"�EY`�<�P*\�\`�	���A&;|���c�_��Y�ў�'��@�Ŝ%�����8��
�'����ޏ2ܦ	)��Ɣ�*#�2OR������� �EÔr����\����
�'/�`��%�8KL�s��B/Rb"���l͠!1�D��Y�I,&��Pn���'��>��[�����k�x��г���U$C�ɫE���)�>r����i��5�B�I�[xɁ�ʁ�Itxl�6���Y2�B䉲 h�]��L�<42m�'V�9��B�	�;t����kˎ /��aEɕ�[�Pc��G{J|bA�BJ���I�ݘ{��k�e�<!��9FՐ9#%�[�3�����_�(OzuE��O�Q䧇J��� ���+ P�)"O��r�*V,3�v�8�H�R�Z���i�(#<�-O��?A2w�[hN<�a��"��Q;@)|O��%��ƥ��n8:��ƈM$U�y��%D��z�59�ąb�.O��`b+%�O����O�8s�g���e��&�Seq�F"O�9r�n�"/�D k+� ~I��)�"O��%i�"(�Q��R�o/�l��"Ǒ����?�"3�ْ d8���O��b>�C�d/ICąh���ݼ�a�M)D� � kB�J(Ƞ�w/S�r��DB��4�3�S�'=�&б�N�N�z����Rf�2U���P�'�� �dH6p�x�
��(`\}��'��$�6O�f��̱g�}!�'}@����_-n�h�#�n�& f2��'�
5�C@9N/Z����	0�6x �'`� �[�d(���+E�-��'^�Ɋ��H�9����ڮ$�(��
�'!�I���
�|�4�C���������*��XND�A'��1����'/C!�͇ȓ8/^U��Ъd������*����	4�pp�O�=Q��)b@�L����q��
!G!�}%�§nм�'��}�-��,���{��x����y�DF�zZ��ÏB�J��:����y"�4�^�!�e��C�[���'�S�OB�z��X�5��*��8m�����'�:5
d.!"]~��gkӑ<�ȁ(	�'��0�@E�d���cD�ϱ*J\��~��V�vYpG��B����b�]�y�iB8Hx��-]�'�T<�Q��y��'kR�Y"���)1��	��!�yrh�z��8�A(B�_�
�q璊�y�Ά8~uL0�gCT*]` �[�F��y
� P���p�<S�)	�#�x+'��C���Iǘ.�� ��úsw( rկR�g~!�䐃�\�ڠ��?9s���d	�$*j!�dӣ\�ʤ���PC��aw�3e!�M�g\�و Mq�|!C��%2!�$�����qp�ƛ_uF��7�V5B�!�$%��9�`�� [�\����'�!���(�����$�*<'*E�����nF!�DT�i��P� 9r{�a�A!�D�;Y�P�+�e�~U)�o��k"!�:QW�}�s&�Ua:\��m�	!�$�8�p���L2WD��Ì�#q�!� ��,��aA�$5���
��!�K�Mw^@	œ�k������_�=!�dN���D�FC�.$��@h�Ï6�!���xϪ����	�z�@Hă�[�!�����&���`aBN�NQ!�$��`����'�6�*�'ڀ.F!�D6o��ܱ��بb�(M�ɚ,?!�DI�/ꨠjsDL1�8�#��Ճc�!�^9p��ԭ�7����G��%�!�D��:J��A'c�:Xâ �E��fR!�d�D�l�����a��M�&��eF!�K>��IS�.@�t�ma�$�t�!���M��c/�\Zx�ǃ��g�!��L�8�
t�;OY�H)�ޕ2�!�X4q�8I�G�0���+���!�N���qC��&`�JlypD��v!���f�b�%�.O�Zً��Ďnr!�d�4�\#5i�
�%��8�RA!�'�P,�Y�腩�9u��RN�X�<��,z��"p�M�I�9�ʓM�<I�!ľ4}vM�� �N�x�m�<)f� C�&H� mŹꈑ�w��a�<���X|t╩ߴVJ�x�Bh�R�<	&�U?:�R��C�!|Ш��SD�<�sCM.�q�'d� lZ���C̓c�P"0fU 88�(���۴~]�}�<��lQ�g}�Ha�ͽa���S�W�<�Lݛi����!I�Td!���<ybjScz:%�����Y���ʰ�@]�<	E��
lm
����13�)�we�l�<ц�Y�b]�c#��G�1"��s�<���A�$�p� �D��xL���t�<�vg�#�Ќ��g[�L���PFv�<� b$P�ء��L~�ș#ex�<䯘�>�ޙ@TkߙSJ����{�<�D�4�-Y�N�8}��� NIL�<9�"�<S��x�!�Px�¬�`�w�<�À 4r�`5S�,8�㨒U�<9h�I6��9���wNa�E�R�<qա�8 ���F��=h 	���@v�<��E���r�)�➶�B�(�s�<��a˼n(�$H"�ӷU��ɢ�
n�<a��l��<1�"��#��y��d�<p(�\P��\�l���e�b�<��`�2|tRi��d��ui���FB�<�1��g`TXdL"k��@�E�U�<���,n��У��}P�����Ry�<�3��>.�#R�S�)�Lh������_�"$qO?�R&�9_�J�0�&�� �`���s�<�c�;/{��J�#H�\8�H�r?�3'�Bd�P��"LO�=f�@�E��iZ���'1�DS�B�,�#�I�zS)��n]�o��q��5���B�F��	��44�
�h7�[-aV�O�q�el�{���qSB���π ���Ly��) �ļ��u��"O:�q@���p���7d�R�"�S1 ]��J�Y:t��h��ת#(V�Y�%л~fi�F�ܓQ�!�D��a��ȳ���pPRuc�#Z�D��b~�Q�N�j�rT[��'L�<`�%K�$"Z�JWo��X�H��čw_��C�{J?�R��R�x�g��uwb-���hy^��V�[��j!�'GV2x���`[�kL����	�`b:0�ݚ�?���.�F�&Q!ԍ�'��mE��آ�Yd�~r�ۦ8�̹��-��]b&eOx؞���U1Iɮ�)��W�M>�٨� �c��D�*v8`�x���,,Q6 ЊKQ�J�#�v>�ٰ��b�)�*w;`�l���Z7�L�G��c��*�ʅ����Օs���RT T;;`D4�� ��3^Y9wn\�|��fةM7��	�=�p5R�`�8i���Zt���!v
����O��Yw�P�;�dj��;l������>?R�D�U*N��A��/K���s#�C�T��D`^=�𒤘(�u�Fp�\m
p/��b@9�� �#���'p������Pp<!�gѽD�H-prG^�隬�Q�ǒ#|�cD.��%s���{"c�iը ��Wqn�����'04\m�v�n�nIq�H�+9�@r�c���Q	r��D_�U8��S�1��hP�c�GN��qP-*sLO�@bv��0s� ��<FZ1w�4�y�E��6��h�F�
;��7�I9����"�ڠk��}������N<(0�)� ��?��D��Yt�E�1х1~@��A��Opl;�g�����
��-�	;���ZoL�9 y�TGF0 p�{p�H)3�Ԉ�#ᓗ
�f�,�`бM��t�����ޔ�r��a�M�־AJw�A�	��M� ����x���Z�p��� �_��x6�JF�	�AC��$pT���"¬ְ0)��23N{�gԺ?%>��AM
�G���Õ�"|L���"B,Լ4�b$_4.0�إA�.w�dS(*@�Y��B�]���g��%F&�⒄^7+>��5L����<����3c�	
���u��/�lI�S�=1ι��O��V�����V�>��ٸCȺ��"�s�*D�E�O<�!��G��2��i��Κ���{����}|tpr�O�5>���Q�:�d�<��Q�*�����'t�Z�s�鐢@������Q�RQ'���
)z��N�8YeȔw�^�c�)"G���K�$T�L9��0������%Q,�� �*� Hݔ�O�� �ʑ�L׀ ���ދ��qBu�
�F�)��-	0�z����H��};w`<|�0	`�� )���H�q ���'�T�'�INuzԭ�����+T鑃~?�p�G�L���e�Wa^΀�#-%$�~���_�li(f�M<��q2R�8N���ݱ_�Yq�&�7p��@��Ry��q3F��1|�r�h -��<�`�w-��biV�-ޔ��S��~��Ys6F��x�d�$� 0�& Y����O� �Z�ڰ��d��%N�(~�:$HPNԫjN4PP�A]�����B �@���O�`!��6aP�YA�|D!*6!�$�L[���4��g�1�	���c"�P�e��h�B�$��Xk�*]O*��q���6)<q��44���e$Í�~tyc�iO$q��&6��H�Q�ݏ)mK� vV1R�C�V���mA=97����2�}x��2J��H�DQA�O[�~ud��'��vlY��P�R�D��T��)p\<2p&Ɨt=�eoĺOR<��� i|6�ǢY��� 7	K�U��(��M,�tLhr�V�}QB�ꜫKEذ)U쑄'b`��GaФ�ډҤ$�W�YpR�=�uWi�p�<=9��3B���� -FP��&��uQ��Q���9�6=��6	V�����@�1�	�'��qS������Y*n�0&�O,q+�jƊ&Q����׋a��h�b��@�~�B%[�\ |�`��N-EK*Ɗ'T�����H�6E���T�v�
D&"�� J�5hT���! �n�0Qt�|2,��o�8ATbҫ��|��鈒#$F�[�<ۥj
!
:��iH�"%F�p��M3\�ЌH2@�Y��Q��u݁1���4 ��4"��&Dv����$#VpA%LA��"<bT�p�d��I`�莎a��Đ�d�+��`��D���8�K2��`��/�f�r�j��_?:�tAS�̅���q�O+[��{���֦�����?���r� �>|'d��R�t`������	H��/Ժ�,�iW�	Z)ޘc�@D/$�P���ph����b8J����� 7�ʑiQ)ڽ\Fy�q��^���k\���ŋ1%���e��I�4�ޡ��۾THm�)O��b�Eř'�����
=M*q�c�%\T�A���PB�賄R�b?�H�����#�o��r�l��̆�L2��B��b��L8�Å%N;dk��YQs��2��͆4Fl�2Eޚ=�'\�(�)X�e[���5��_2��ԣA-��q!��qFC���5S�M��bq�"8h*ĳ,^�4�����mv/��������9#��\/x�
a�
-p
�܃#kJ�S�\��'Wl�{��_\Y���eBޯ�\� W�ָN������*X%��BqÝ� �X�;�
@/sk�|�%e;ΉYD81��n����� gӐ�[1n����a�s�h�&� r�)=@���ab�?t�n�&ߣwذԒs$Ɋ'��K�N�n0�=J��,8H���A��ԡ��h[����RJ�	�L5qV�Km�4��4k�Y���'��|�vSH�d�l�"r�*b�Q�-�j�RE�H 6�Ot�p ��j9��@e�]�d�(m�D�	`�lڗ�j���L��)�������zh��jF��|�r��f ~��SŘ��Jc�˹��I{6`�
=R�e��)1[�I /�hYV�C%�@��E sОQK�J���!hMU�ֵ��m��}���к��8	U*]�;�9q�q�|b磑�&�D�ϓ! l!*�L�g�n��a@��V�%a\x~��5d����;v閴q��W�?pc��:�>�c��'� �H1�H'<p�(B�ѻ3z�c�i.��'�"F�,RG�t�̐M�0��#�uǃ��rp����)[��谆��`h�@f�Ͽ=&���5�I�i�>����b��o��T��$Ccc�<@v��9(��g�&?8x�ր�"=�P��qT<i
ٴ.�Z��^�C�`��M#zx��|��&OeD1g�ܛJ<��-�d��u��s�¹�d��{����Bnר^hFY�]�O.=��l,�n���s]��J�D+@,)`O�1
;L�pBeZ+N��Ez�N�#�����L,�����8Yt͎�"ԙW���'�I IH�B��l1��ß|�(1P�@_&��!�M�*�����O�i��$MR�G�ǘ-�B��ѫ��U�(!��>���WU��qJ�T(Y���O9~7���NK���\9�u�N�c%
��O|\��M��~�N�6BP�<��@��%;�U���՞e.���nϕ~��![V��xU ކWW�p��,B�T�r�eOU�epe%�'�yRm�#_^��@5�UP�X�#�àP�h �Uŏ	(��0�g�A�N]�\Q��@�bWt����#z� �T�ɖ3�Tz��G�)����f�
� S�T�{��D���҄)`H����с1�D�w�~16q��F��SMԏx��n^O��i��9H�9�cY�/q��{C$��}�����Y��O�t���#R��w��� �%��#��bH �`�);:6�a�K�n3��zF���M+�G'8�n�S���[�.� �ЋQtp`����>&�~���/hv�;c�<�Z��`�5�	�=��zu!�\��N#&z����Z�V���,N"�$��"�֟|
i�U�\&��(����;/�h�� �P�[p�y�#�0����	x q�%g��\`s�
>K�@�茓k�
�����PRFBH7Do�|�$�M�I�,�)R%ߥd!�d#&i���wiф4A�����",�h0 �8��9(fBb*��B���c�a�(����dL0�L(�j��r����s�D�$c�Od��1(Z#b�tXK����N4�T7j��fM5u��L�t�PD�l�e�PRH�ࣃ���`���P؞pH�`\��f!���[�Ёu�@ry��IG�L���E�Ϝ[��IT�V�p�a~�
�C�x'�C�-?4� �I½U��CP�H�,���fӇ��F|R�
�w ~0�@E�"}h�x��i��֥�){�j�&N	d���5A�LI��wI�>Q�-�-��U*�T<O�z@3����t���Ҁ���xQf��<v�`S�,C�$Ƒ{�d{���3�4p�(�"�";tI��lZ��E�i�E��@Ĺs�xq�m������>E�k(�,2<h!S6�ک<4\��5�Q��Bˌ�Z�ayr憙�+F�l��$�1!B)�3Ƹhǎ�1e�-7n\����bl���̙�V��z��F��"���߆Li��VP,�t��E��|�6��d��Q��騆��>Nc��86㞲L�X!P �L�B��Ć�c5�	�4�� �X�$�U=Ii��Þ2L�R9�NHJ�V���FC�1�T[��دI�� �2}w�lrFWg�9�����B���#kj}�a��`u���~��㵯��0%�6:�I��`I;X��P����nm�?ArA\�HZD�  ���W
��X��Ky?����s���/F%\�7�9J]T�@���Q ��`�d8'Ա�&U�G�b��ea-:V� �@��:kD�)�/W�Y ٪ߓ|>
�
㬁�gPT�G�77�������=���
(R����Vd�p pE�=ƶ�"�.�nl���w��xر⃎S�n}����eW�}I�/˄����4ڶ R��<�f�1$�B�{�lm0CJ#'������C�(���W�7߰,R��<�l6j5�h���5!�04�$X��N�S�LE���O�4R#���(��tӲ��v�UX8��t�w�~�IB�A-e�*|�E�M��T /�'��rJ�\2��	s�t�iN�,f��I!$�J�p#"�7J��x%&?��'����*��8�9���	jH��ؙ��,��A�CK���aNM#:�^�IU�\��f��H��� �shEUw����FL���1�-�*Q�[� �I��h��e�����BeH0R-���>Vp��@޼.W�K�`UK��x��%����B�������&ܬ8�C���a1��/؈xo�Ɇ�	�a �L����G0HR��m���-��ybD��$%�����]ڦP����@(db�(n��9ȵm����(	$LL3C"���J[�Q��ہ�'�
���/)i�V=8F��9HS�г4�49g/�#Q#��K���g��ϓs�Lb�b���\h��ix�Q.ޫE�@H���
��J���,ªE�90��S�K&���Ջvn<���H�V]��՘D@P�A��zz�Q��J��9�����)x�ɰ�֞y�P�2*��]|���Q�~�ɧ�D�*�����'�z!�%z䩋�������;�t�����C���1�K�[�δ��+G+�B�iK?�����L:�j�����&�Z�ŝ�lN�FE5A��T��A_�����:����T�-�Nti�����A�M�HmӲ˄צ�:49~'F���تk^t�ТLB�B.��7�D;�����*ňvX5"5�ar�I��0<a�`ʩb�� ��J�N�s��/<Z!�Đ��c �X�0�N�Ӣ���+T$Ѩ���uSi��/?����4#��ٵ5�\����@,�X��gZ	���f4�L�'�"�*TȆo�r,ɖh���߄�`ڴ|Lx��� )V�aɵ��2�v���n��j�L-�2�^].����n�DI����B�'�n�ې�H8	�� c��Oi|���s�?	������'.�6���:}l��!u��Yf�Ğ:���S�ׯ�; "�P�H!�ǘ�a�6)��EN3(��!�*|O�<S��@61���J�.��)k1���xB`č*u/��2`�ޱ�
��wD�44�ؘB�"�-��9s�zD D[Ӭ��D>l�R,cdN)��]�{m�x2$J,[���y%��1ta�9��imj�Hu�H�64�͕�O:vD{AƋW"�����R/�F��4�6ln�`�	�
< =ɒ�TI7lh+�'�Y����x�|��F��9?�,Y��I�����/j���˃)��M۱�˺��k��(��\���C�l�h�P�KϟQL��3r�X�v��Qb���A���)��8#ƌIJ�k^�de�$��R����0�L,}���	a��m���g����'
;_�6(X�Q��г���w������	c��q0�(&N�nk�@��R1�L�3�Яc�@m����0��<��X ]�>���wz<K��X���^-Z2��a�3u"V���)_8Zl����e�ޒ�c�;�|��/2���&�yb��pY ���9yDMPc����'k�c ��2,��@�'9v��� �� _N�2�`��'ˠ���$	�:���(�ƍ�6�5j�L��I�̯�|!F�ISk��u��	4C֤P�93�l�;7L�	�i� �	��I.O�@%��n�5>4�ֈ��p�Ⱥ�O��8S#�&�o�N��/������϶C��0��$�O 
�@��]�LM�ϒR'�� Ӌ��E ����딧7��b�	0��f�~�b�)�ᦉ�D�?i�HЌ}
�!��"t@���#�а=Q���1znhZ��Т#��+|m:"��]Q��s��c�
����%%�*H�5��;� )��ΟXZ���_R�ɚW��%`�A���渓h�&X�Db����0`D�R'�@�z�Dh�c�"�zC1�,rDU#���S
�P"�'�1يӱ��`��T� Le8�Db�7/�b���:f�ĵi�M�ey8@�2�<H��{�\��u:>hK>YD���nٰsi\dßw0�C�F	u�*Y��lih<3�'��Q��k�J "7�ģfi�l��+�7(��8��E�v�R<FF�]��UÒh�n�P4J���!el�|�]cִ�Kƈ̮nb�\ �ɗ_�ވ�04lO<����Q7��:7��h�àF\-(H*8�f�^�ڽf��h����C2k�4م�\�k���F]/����  ���GQJ1��m�9(��i��ΊijJX�$�S�@8= � �[
輈�fE&J<,�)�E�^��a-�}�vu�IΪ&2Dȉ�aI��H�ߓ�btP&ˁ?VA��R�2���(`�ԃ�`��bI8��C	�hdHkA>	@u�`o�V�:����E�)����Q{��B0�
�ht�]�ȓ&Q���Y�~�Z!"H{sl�y� Rm�4���. �$��gǝ.U��)]�j���yqn��1IVb2�(]�n�L�a�g6?��" �'~�q�P-Zr�����t�A��X���C&d�es�J�f��Չ�	y7�Iv��?�I&�;��<`��K�I�>p
r+�VC�� "�ꈾ2Μ�ǎS�|�Ob��1#��?���R�(�,I�����9����s	٭q��݊�'��t٥�
�� {�K51Z�)�rH��__����̰F�i>m��N�4�
Q��MM�m���	%]*H@�r.� ��p�D�6'��B�I?��b�&"�|��%k	��I�4� �cU,ܵ���}2z����z��K)J�Ng�\ы���=@L�H�dmx��@�$�-ݛfA�1&U�@�+Q7T�0ƤKz � �5�~���{5*A�}&�й`E_$N`OS��r,��.$�\�-�8cp�ub֦�O͚x#D([k�*�VG&dnh��� `����Õ$����խ*����%�����U-��� �v:���`	0S�B��`���X�!�$�i?�X+��~t�D�_*k�qO8I2�o�5�0|�0�W��e�e��Y���2D�m�<�Ə%�T=�N^�Q�+��Nk�<ab-M�7��EZ&ۻ~d�����k�<I��"\m u9�-�4(�2) �d�<�&c��3$�0��$W�AVȴy�H	e�<ْ�J�X/t�B�,�|��D��f�<�ٲ`\���Ur��hS �K�<y�¡=��i�@]
�P����j�<a�CM�G��H�q+�=Lt� $Do�<A�Ӯ7�J�j�*�>8j�t0'�_�<����x5#� ,&�H�K�HDP�<YvhU��!+T�-0���QC�K�<��C�:jbi��/�Kl�t:7��X�<� ��aL\@�� �5��Ck�L�<��U+RN�X��P,<a(���*s�<�v��d���[�Tʀ�1F�m�<�ƌb��8�d�#����n�<��)�;:�X�kM 4 �Iҏd�<y`f�#}@TB$@��"�����e�<�(K*^��-RؗE���Sa�K�<a�׉�p( 5`�6�Q[���K�<AQH�+&��8�fZRp����R@�<�pm���q�H�� E�R��X�<Y�i�Ap�@��C�=%FX�p@s�<�eb\
;7:丁��9,;�9zD�d�<�V ��!�V-��oݓ,��X�#@�f�<���L���7�&6���]�<��:Q;�P)�ʛE�D�"���\�<QpM�>��b��|����Yq�<��n�#b��ebhE�}�^u�c`�t�<a�&�1����	;��a[� ]�<��R�oB�D��MX�ե<�`݅�
g@���dƋhr���*nR`��P+�˕�=J ]�'̕G��ȓ=��<���yN	���(p���4�T)��DZ4VXPH����DI�y��(���t*��c�Ǖh`����qi���9�,���S'����O5�d�q/�@���Y�ń�p~�%��%$j���%�7����	�++�ȇȓ2`r��#�1Z�9C�۸7U����l��iK�U}h�1N:(��ąȓ�ڜ��ɢm՚�H��מ`�pQ��5m���Wǅ�>>��)���q���I�~wX�����9<�4��t`�&"��Y�=hjԥ��S�? ��@�H�Z���%�ɏs�^�X��O����f��Oz��V��D��2N��d� �^�~X��IP�����cR*e�1���0 �~ b�U=x����Msh<�VB i�Tdj�#@�]j��Lk��U4��JeM������ '�Ӹ>��0�u �=[r�E��%p3�C�II�Tz7�P�b�
L���E��Y�T���s���* ��~��$ ��N,@�ŭ|}�ْ�9D��I�m]�B@���D�h�@= bCwӴ�K*3�ગM^�Bn��Q�̵���3�`x�u*� U�1ȡ�ܛi�qO��j`��j]"S���]�x�p��9ᰬ��-�%!���׿��?�&Y�?�hESL̽@������ٟ��햤1���4O�YJ����X,;�~U2[w���K?�8����2�X��e�,���e(lOb����VU��Q������ރzJKс�v�l��p��(���W��1�%@���� ��z�ġ�w�j7�aج����E: !��D_.{Wl3�{�oW�)��M܍F��,�!Iѧ'�tի�@{>� G��,��l�pCW%EF�VM��qt��r���9h��$Eo��\+7�'��D���� OV�&�5sp�iS)ǝ}��0��f��SGN)�JB�5�b����ʢ
j�`)Ed�S�(�Jci�ݺ���&]@y5$ը��p�;:�,C�%�$1%*|�b�Z	.B\�#oS35X@U3"�+���bAD%>�<!{ӥT�0! �(c�� �������l$��@2�pi �b>gf�< �C$�~��`Ժs�~0���Oi�zsˎQF����4Z�h�!�'Ю5�� ��0J�L�e��H�h���gv�rsk!0y�t°e�+A�`9� M?_YV8Z�7O؁z$*��}���%D����� V��y�s�.)!��#	ȕ1�����Wg�!�ɗ���'e�#�V%��pɑ��j 1�F�6�r�)H͠�X�!V�N�
h2�E<�Jl�L��`l��T��UU䄱�����`vaW�J�t
�E��9�PX�L[
b�iH��.HG�*�c֘<!4m�`/�B�`����!@8v����R��q`$��J@�4J$�כ9$8m��o�B��3dN�4�JyXdW�7�` �	L�2E��1�KU�A�f�!C�q��<r�d��7�XQ ��|�%�P��y��	9	~�c���[R.x!!E��#~���s V�1��1���C_��IZw �,���rb�I�1���j�:*��  Ǌ'J�(Ic�L�<�˂-�!t�p&�����%~�@�$�ӓ7� "�o��|���x�A͢TЈIu��U���7i�g�:���&�:d��:`�(9cь@�4�A#�ժC��c�`��	�jO�D6�A���I)��D4�U�0��+"�~HQ�
�#��8!���㒀jүF?(�R�+�8E�&հ�/B
;d�0�0��r��k;�&��3���	64�*W��:A�4��so��=i��#ҫG�L��s	׮P(G��>s3
�JT�U�?�h������v*�kף/C�@��c��dp �]���`�kP:V���g�rx��r�f�q��=��`A�v:dHw��g��y����\Љ�'��q~��"A�<�D�y�-�En
�~I�8�TKZV ���`]2[�8�g�ɑL��Ex� -}��UN�0~M�0ل��Dz@M�k�V����Вzn	���N���E�Vn�o�	��G�KqO�L�s+��#x���/��7~<��G�[1�}���� ��j���|`��P�.��|�P")�MK�/�m��@�C/Kd925&N�S��]���Y�2f��)'CQ1��\�2P�h�R���G
�no�@у.�8e5�&H���\kU�ت�☫��/ 9�T�ʹW���9i?D�Z�@P I��6�@�R9��Y�F�Y/"@��j���`P;>R|ճ�
/K_��
m�:���S%��h�d��Y�5�ȸ�@H���^5W>h}��,�mh�E`���v�"����G�6�����d�8��'0��q�-��Z��,���N�Y�p�"rcI�f��'��)7bP�`���\�2!�׀A�}�Ι���rA����	��7L]
DZ��S�6Z�2)���'�н���<,�R��'�&�M�7�L
i	t����z�RaRB�P4��z�ViBR��4zqȰ�`��v%(`�u��&`�j�"7���B�X	₆]�Yj��,sX��c����w!0T����ݪ]>�a`���>V� ���Q���aui�;�l �C5}ҪR�ct��`�Ǫ�%x�J75�<�&[,�v��q`´s�ZH��BĐb�T(���,Dp4|C�LD�i.@1��œ)LZ�R�cӚ��ƍ�	#���h%��Z��D�VΘ�S�ƬQV�x����ů9�%�d'd ��	�2%6HЂ�A��W�֌��q��Ȏ���'����ӤJ d�<c���C�|k����:O� 0afN3E��8TA�6%����Dn� K�Y�L*����~v�ӓ,�+g�8m�W�O����'=;Ɗ�R�J��zA��j�A-|r���,Y��T����^&~9��/��-��h����5�(�0��GJ:b��"�I�m��2��7�p8�,O��z(L�K2̔��d�Y�k	�� �d9�Y�3F�"q�*�[A rE0�A�]�=cZRW�ӽ�(WD�6�i�#��v�>�1���V��� �
�!w��{�ޗlN��a�O� ��ܩ��L;"�Ϊp�J�c%J:�ġ2��
�!��zw�[����@�
S�Pȹ3�8R̘)����-,�8ݴ9t�9�����jS+�*��N��F+��.�|9r�,\�Q��I�)W���R���3��Q:���a���U(O,�b,�%S���ݨl�H���w��$+B�͏If�p�� N�D�@�2)�2"���H��lya�H4,��42�̍Mn�l��@�<����<|`�`�7#�D�fA�4q���? ypBĦ��C�&Nr�8�@��#	gR��PM�>hq���nL�3��8���3��J��֬F�8�f����O�?��%�T�H��Π:�bG$�a�!�1-�!
̬�J\0��𲕠(�	��(5��%c�Mͭ^`��� ΢7�;g	���ū��<t��\B���uK	
�Y��P���'� H3d��"򺐣U��=�(h�Ӂ6N�B��9Z�=-	}9��W*[I�8^����#.EP��r�ˢK����;O8��.,P�8�\wo��"7瞗"xLpI�B[*�X��cJM�t7vXJRgE!���ɕ:��p �#�妥�R�OP����̅t6ll
��Ce��a�M�7n�n��fJ��y�6�)tfڝ�M��M^x�\�Ѱ�P'��Ӣ�n��'��X���W�yNHJtX+~q�e
p�޹?�d�:�'ĤG6����X'����c�*vPp�#Y)}t�e0�8:�~�:��G2��yP��ްr�>�h�8�n8�W	�G�'�8��oY;F�B���B�y5��K���9����H�bAx�[�	1@�z��C+Ίy��H{��8-�<c��W�>�����H5eKj��	��Ń 36�"l	�h��#��#­]&?��K@I'd[�Hv1X������!dӆP#7������r���\�y�`H��F�u��"%}&-��KQ��
�1�R$��$�Y�M�����@���M� �l�po��YƧ\
�<�(3�
�	��5q���e~��3�L���k��aF�]� �P������|��u|��x�c�;V>B��M��?I��Ɉ33^�5�����3�/Q���ECUe�`oмm8,�e )N]0��a�'
�݃f�B!,^���EÉPi�@/��my0 ���A+J�P(�#�-$(��
nS��RL��c:T�F~R�%Y�V|�b�c&	�4e�lJш��՟��02nS�J\zЋ&�IMP��A���"�8	��G<hC��d����SNVl�Ӏ���M:���Y�<h���d�]V����۲!ףn%�l(-I26}ִ�a��;-t=�F ��pP�ܠ�d��"�Ą�%D�i
�#�e�+Hp�B��	LUF ��>sX���D�-!�̌謟���@� ��ѢU2!��mB�K$�~"�ޏ��)�oһ^�&Y�B�O?���x���M7K�%i[
��7*�4`��=�ƥ�5,Ԉ�7Y�6���/��!!F�"ϴٖ�(O�*�e���#��E)u���������:a^V�"��+���J��MK��V��kS%�9X%jVnƁ(m�a�`2����%�#d�`�
ۓ{���;l�viY�X	�-���E<q+w��&7����iІx��¦l��(��4c#hh�� �<'&ѧSV�QA�"���'�܌I��G|R*��0�6�����2}�J���i���jL�j(��3"��O�QKd*�7G�m����8!tl6�4X[D
(}2��-��N~BC�ד$uI��mV��R� ����<Yb'P��~�P�D�S۴&J�nڴ]�
�{1�@.������e��E2���o�:x3DM����o�>p#Tm+,O�����%��M����|��<P�,�	Zs�R��\��m�w��c�
���O����,¼NE#�w�VlZ-=B���
!�@�����GY��$"�\∲��P	:H��S�)N���e`N�=���3�D/?�J��d(ڳZ�����I�'��H��烧�� !�(�K���э��+��\���� LQbR�*���F��/���I����c��5`�t���i�=n�����lON��%o��:��P��LB�r�{FK���)�G҇c�Hp�#ݲ[���89��`� �C�b�S��?=��F)P�|�b�֚ �T�1D�q��������=N���X�O�ú6�X�}�t�G�����i��ؗ���Kx���Y��M߼˅I�0�D��G�]<',8	(qo�[؟(c��IN�iY�H�˷ub��gIE*�Qk��
u��xCw�|�B��2�ѷ��X7�˷��'��읒 �~�{ҡ�3�����DΰvI�H�1�ɇ�66���Rv��%or`���l�;gH4`u �[�����G�:�jX�C��W�<w�٨B���l�0dF8ɖ�^�#�D��1��=jE���GAۼb@�	���	$�"����+x��$��Li�C5&8���¤O*|g~�x �����?���ѱC�Q�3��s�U�"��8���N� vЖ��Θ.SZ����"O��4���p�]�ʟ֡	��Z������B#r�l����*8������$ ǎV`8���$�6��nS�y=�|����.,�9�nS�m�8���Η^<��
`��&�4���|;�d���O�8����=`2��"Ɦ����W �`��ɦ>PH��!Q�Rp�I��4�9��+R�mn��0
U�*���A�'"*�0-��&��
�LQ�"�˞G{�%nZ�$��8P��+/Vtm�(����ā�[�
$�F+C�B��s�-?A�͡U��2aǕ�w��0�dK��&��Z�P*t^�q�Oɂ*����d�ڍPX�����2�R+؈OD��`1%�50��@�m�(������d�Q4�GJ�1O����A�mO��Ae@�?y�f��ěZ:���$X�U:�7�0J�����<jC��I% 	�>��W#7��S�AܣI����.�6���Ĉ�9��B�R��`���اV���PX�/B,�iP�i�0�TJC�|�){ ŉ$?⩑6�3L�<��a2U����T�rГs��
�ҨYE�8O����+�d(7F� ��dǃep��p�Q5B�q'��H�|$PV�0��! ��v",4�lgw��(�+�?R�9�"L�r�D�u�B\�V�D�F-@�e�ް�I	[�T���k>g&Ȼ���H�$�}�B6-W8WjP���  |+��(��=9�^�3���	wڧBݍdr�ˣ�D�f x�`�I	4@4����+#F.��Պ9G���d��L���	�!��W e�@p�BH�QK�tPիUw�b%&	<W¬�f)L�[�f�Ck�G�����(n��<�ߓ9_ؘr�
=�˃(!k��d�]o��7��d�X�j2���-A�9��&�"xZ�)��U�'g��$��\j�$���@�T�.���N�i������ؐF����;3:�]�R�O�aE��3
uӰ�R�O�t�^(�um�x�F+ˮ(�����I���LE*��5n����ˉ�
��%+�%qg�LÖKJ�<����=I:��U�#5?윻S�ǟ�ҳ��^��<r�88�Ll�ҭ�(<K8��!;������O#�DSъ�fZT����:KLLI�nJV$36��X[��됤�v�d Ų�O��1˩���9�]1l���9""� 4���1�\<��+�" � �a�+���iP��0o���b�M�0��*�_Q���`a�XQ��D�G�.#����剱=�bѡ�/B�5&G ]�d�RȰ}oแdϏ�HS|*�5,{���_�J����E�  [�@��G��~i赑\w{&��7j��QƋOL�Đ%���b�d��l���Q��3�$���#2@ܝ��������Bd�K�d��PYAL�>�n��$ƿ&N�,B��J��u��f�~���N����w [9�DuKFǈE%. ٴ��>��[�i�4c�l�(��C�|�g@�9��tOǟ4��g�%
�aqǤ�C�*�a��~7�~��2XC@����[��]e/Oň	���K�P��^4R� <�\w�f9�g�;R|7�)y`��,y��8{ �Zh������8Q=؉��	�y7zQS���T�>MA&鞔z�C㉄pv�H�a$��y��Q��Lݺ2�P,@Ǉ��D�D�w��y���$�u~�\��OXm��f9B)N}�-B+t �[��D݈��;e�X����D��Ƶ(�8R���٦�׻:�j��6꞊BA�u��:l.p��#
h����$GV&�xA���5X��Q[q�Ծ"xh �bΔs�uõ�5�^ɯp5,�zqK�tȤ��%lZi������ ����3q���d	��-�"O�ds�/׋l�e�'���W��YH�K�R�l�p�F]�x��Lx�j\�b��t{���f�Q���
�S��Uh���X�+'�Ŕ9���T�ɽk���f�p؞<�烍8f��0s��	*
Jͩ%�O�S�n�0r
5 - ��U�U�\��i��׎ ��@+��\L��EhO�W��O�k�e��9��̭8�vL"F�d�>���
D�Hp(����1����AIX(G�Pd�'�Z�����K�;�&%���-4w�m����޵��1b� ���Z1t�=��˝?��:C�M�<�9׮[�N2���C�˭3g���a�0p�	�ăJ�;�����Y����₰�6����ܬ_pE�ȓ.I�j�m_��t�e���'B0t��Q(%��MX��YL#Ҥ��*N�Z_���\�� ��%@2p��E�\)�4hDb��eX�_��ɪ��']�Uȕ,���L5�tE�<]�<U��G\:3R��)@�
�V�8����\}ĭ;3% ��x0,�?Q��<��-tк� L 
c����*Ǥ	.���A��X�i2�X ǉO��U�v�*�J�D O9�B�yR/�%�X���L��+��'�H���*͏A�8��$7�y86�Ĺ	����G�J3	J�i>�Z�C�,�4�PŅo���ɘPD*���I��R��D�t��C�g��!B ��zD�X��+���P�I���#�g�X��|(���r���ޑ>�.��ϟbA�2��dQt8Q�@D1'��m�r�'��e�RV�8�OV�J(%2b���h|�)���0�n���Ⱏ@�́�v�q��'g��Q*O�ܬР�H�,c�a��'�b��ℓ<-��id� (Ѥ��p�:*K2�ˁ�ߟG�|��/�~XHY�$<����tf,��Ŧz�"0��>���&(��#@	�И��@�'�!�N�NWٖ�rƔsAqO��!#�9�0|�K��OI*m1����DS���`g�<��aώ�T#��ڸHi�=QQ��g�<�%C�
D�����G �l�1$�0D�t�U
(TH����Ƅ׬,R��(D�����	S�D�1c��Q.M��yB(�c���`	L�~�n�&�!�Z�v����>D�8�h�@�cH!�D���ڂ�>>aD���@�\!��� ,A�n_�$���m[#�!�䀻j�~=ɂK�.�����L�D�!�d���PL��.�o�.9"�ʟ+[�!���9D�u:�GR�$-p���0O!�˗CW(�:B��*�����I�k!��2q{v�ɑ�Z�d�3H�+&!�D5T�j��%k�R��ذEN!�""�n�x��S�,��&�q!�$�9l�����{7&���K�,0!�R#8æ}J�aŵ@,\��4���!�P:Z>Yf-V9?;X�b��I�!�D��mĢ um�I�L��#�9�!�!-ĘXĥh.x�C�$\!�D��:@pp�Z�.V�-�y��yB����E�Ԫ�/&	�͝��'�P9���EHI򷥌��T�j۴�tI�(ɠI����ȟ�L)t�J 	�����
(A� C�ύBF� ��kN~�,?��-H���V���,>z+�tb�躟���LT��M�����a���~�P[��%V�Tt��M.��$��<�`/;��S-w����רK��#'ڟrO� �����Z�jsb#tmѫQ4`Q
��T�$��I!k�Q�"}j�B�`��:WN�7>�$�t"�ҦE ���a�e�<��P����3V�X7���x�����N3q��L>�� lQ�F�������'F��=��C���'��9���#���0Q�(��Ͽy�tp[Q�x"�K^?QAN�`�O�왨�e\$�Z����:;n���O �(��T���y����'B�t
e�P���@gO2^l"�n�N���j���S�O�vI���� �p�0`N�J� ��Nה+��c���ç*,��E!S7����,Z� I����� H����	H
,M �l��P;�B�S��O�թf�Ţz�1O��i��W6r�*�E)���[US�����y�S�O�8T�5E`0Qd�Yaٴg�H���T>��'WZ��Zw.-����^���i��&�|��"/�j�L5J���O�>@ЀŖ+Zt�U���(e�� �C�Yn��	��B�*@�?����� >T���+g��J�G�$ 8��_�<+�Nh?!	H<E��C��P���!�&a���J��U�M�#�]�2@�4�'�T���t�O)�P��G���d_;h)Vy��"_���p�@[�^K����B��H�>���d����C2T�&Q1�%��K~��Cv����< K�HR�#_����G=�$1���SԒ�At'�%��rl2?9��Kv�I�$8��-����)X�h�R >�V"O0��i-Ett�	E��yW4L�"OPph���(4�r���"d��I�"O�M��K	a�V�ᵀ��#Z��`"Ol(�$HT�JVAA�*�Px5"Ox��i�_
mZ���� "O�Tuo�ID(�s��IR��P��"O^�1K��p��	�W/K�MrB᪡"OX�sL'A}�m�'��n�u"O�)° E(T���ۅԺ�� ""O2$�F�Yf�d��Fэ��5:�"Oh;7`�rj�mҒ�M2;�R	¶"O��㱊ďe<�Az�G.E�a"p"O���$�s0����.v�F<K�"Ox�:��K��z��WEɻC����"O�f�xh��BG ��cR"O@0ǮN�MXp��`�p7��{�"O���T�A�4i�wi��l,���4"O*��2Kצm$�D

<�qh"O���/�&f6j�B�� ����"OL�s� ��j�*4����=i�6�E"O�����s��)3�S��};�"O�d���R-d��a��=`�P�+�"O�ջS���JsE��9h��a"OBT@07l		/�[�ջ�"O�9�5o�N�P0Zp�ľ7�dy�"O��)C�شM8���.�a"OQ��#��R`���e�"n�(�"OpI���6��)��B��4a�"O\-:5�&^"�؀P+�0r�d���"O��-VM����ۏI���"O�(�2
�I���c��4 i�"O����В%�3��z�D��"O��8�.Z�#���Cp�ґHDz�Hq"O�iX��
�A���p���/�1x�"O��!�% ����m�k �-Ѕ"O"%�����a���|~�V"O� �6H�d�&x��4M�H@�e"OQ��NM@0���G�B"O\$cR�ݪF�B0pT��+_B��v"O~�À�&h����ټ'H��b"O<d1���Yh�� D	*4�3"O��P�h�di���"�h��d��"O��ڂ�&4��@ŦŪ�ZXa�"O�l:A!D�%�@�3�Ӽ��dyf"O`����,�F�1w��;��8�"O|�qf�N�&�����h�T��"Op�b���H������C�qO�0s"O�&��eVX�䁃�C9���R"O@t�r!B+oG��w��>1�f��"O�ta�_'2֔r�O 2ۣ"Oh(�BBmc�s�
���ț"OX0(�#�9��b�TM���e"O�Bh��1v���gԛ`��"O��7��w}��!��;��E�w"Oҡɡ��.������Žp��4+�"O��p��eA���$�.+�2�"O.�y����`�pB�����%"OV��S�*`�pLQB3VlR���"O� D�R BD����� 1&fi��"O�0DD�yg"d�PJ߄TQPh�g"Op���E�A�:b*�)7%�@��"Ol�"V���q���v��6Bj��ڦ"O��Cu���lI�5I`a�{rxi"O���3,A�1H�S�)N?|�$�E"O��xF�C3�M���)3��$Sr"O�	2S(M	]2��HR��L�9�"OP�b��-� 1�˥q����"Oн��K�`��i��+jMΕ�w"O �g(��H��g��{K�@�C"O��s��&����"�ً36|��C"O&`�� �0r�}��;"F��"O����:KM�i�P�N�v���"O���b�(W�,�4G!�D��j�M�<�"�NXF�����A_@����H�<Y�%�#e���oJ�cRx��ÊB�<1cf&C ��$#RG`�-5��}�<1��
k�h�O~x��pċz�<�1� 	 �t�ȝW�� p1�Xu�<I���R��1� b�O���Ю�z�<�C(Q^�냦<R�n�EAO�<AW�M>�8�D�S�R-�p � �e�<	Qf��,가�VO��0��3G@�I�<�A �(�L�spLF@��0*�l�<��!�)N,��&L�y�F��d�<�W�	�X6`rECL�Z���a�<!�旔(�B9��n�����
�^�<a� �O��τ�?o^�:��a�<��$>�N�1##Y�9�zm�� KD�<9m[+i��	VhԎai$ya�o�E�<�򅒵dX�ua�/��A���C�<A�ԚfC~=��H�9	��ృf�<�tKB�a@��w$�[2�X���]�<�CX�\��� �� � \���p�<Q �G�	���"6��4����p�<��	C�0x��co�!-v��sei�<�M-k5-��]�\Z��b�<Y�ȁ	ON�A�!ˢ�����-�a�<i��5�ͻ4O�6n1��I���F�<���S㚁z��ܲL;.�G��I�<�sK �P��9І0k �l�7�G�<�X�[X�$`���2`
� !D�G�<���E�3=�p��BɬZM4$ċJ�<��!ڐt'���c�E&:q�}b!�^B�<	�d[� �0�A@R%Aj�!T��A�<)"�X��$�� F��ݩ�*�c�<�	<,�fa�}24�]�f�!�Ѝ	x~���.LX-%�A4B�!�d��-mt�to@�jt(��T�5/{!�Ċ$p���E
*yU�9f!�4v!�d­LyX5ITH�SN$��ʞUs!�$];�F��g�N�<3�娢 �0Fc!�U� nx�r.Y:��Ľe�B�gN�A��_�I��`a)����B�	��vH��ԆD�HyZ���
A�B䉯j"�I��͕�`
��q,��u�B�
6������0�T�ΦTf�B�I�}����؇[�����gқ	,�B�	?76h�1!4\�� PB�)yvjB�0�0����E1_��5;�!N-0ofB�ɵf�ȇ�H���C�H�"�bB�	��ΈI�IT�_`M���D�!C�I � 1��B��2�P�L�	L�C�)� �bݚ\�T�x�	�.8�i"O(���)k"tj�脠}����C"O(]A#�ƀs�n<���5�L�"Oz�5��Z�8h��ӵB��i�"O���I�$���!���<7����"O����E��P[��6U��=��"O�x0�ј	��	1,�^�@�"O.L�!��G��򠀂�w"��"O���U�@)Gn �8P@ַiL� "O`���aƱ>y�,����Ek�#�"O`� 䏃�>>�bQ'�-WcRܡ�"O>		�kA'x��3WO�zE.���"O2��)�+;-B� �+_����w"Oja(SK��{R��JrJ�,R����"Od��"�Z�+2]�V�N7���8e"O�M�ЩۀM&���.�#)M,	��"OL1�,�	2������L7جJ�"ObH��%Lx��w�̶|�&ū�"O~����O�J�
`��̅0-�	
�"O�=��畐+e~d�g��$Q b���"O� �f��-w����O0P�r�"O��ء��ߐ��SG]�k
�,t"O���ca��E�Hk�c�d�t��q"O��э��y�D"�A����"O���� ZwX[����]��"O���b��Q���1��n���"O��{�#�8r4{cm�<B�b�ӆ"O���χ[���g)�_��"O6��7^+(�WI��P��z"O�`��L�@�!�h{�NL9� D���Ei�GI���a�3v(��2�*D���Y��� 	�N���Ce)D�h�"i��`(�����W�=�����j(D�l[�o�Y%dᚣ �t�x`eG&D��ӑ�V�P�,l��������!D�x:%"Q��:$ZE!�,20�DC�i"D��yFF_#��	�AҦJVUa�-&D�,���[o��m2%'Q��$��6�%D�h0���.peZ}c"��$
�5X�"$D���a@�� S��̗&�����4D�D'�*9,��dZŞ�Qw$2D��ˣ�
�>�	�pkp�Q6�1D��A��B���,[6Rvt�r�I1D�����֎X7Ɯ�7#��`�hH�.D�<AˆWb<5����w�,���	*D� ASo1Ϭp�ŧ�$����(D�����{�~,��J��yT*<D�4��W){1�I��&<{B��$G&D��b��ѝ*�E�D@_�bZ��3�!D�<���Voz}���($fU´e?D��kqhL�"����SJ��n���q �9D����6A�,�(��T����j9D���kE����m�f)����7D����f��\F��r/ȵi�v4Z�b D��h�@1'�%��dƶ�X �# D��"�@V�K69�Ǌ�P�Ҳ�0D�(q�c�
7����M�CHtPg<D���dfRv�ލ��]8��uC�8D�\��k�C���UE['+=��ӧ(7D�4Y�U�j� �x�E��4�����5D�H+�'��gv���)�B��U��A3D���*��,���%MK:K�Q���y2H�)
�	0�� "ƶ�%f���yBa$���b���p4�ޝ�y
� $�PM�f��{v�H&��]�"O��k�GΈ��*�� v��Q��"ONM	���4���)`.W"���;#"O8y����r8�\{7��i~ɦ"O����������[�.�0nYf"O,�k3�R?�jx ��̼]S,dR�"O�=�&�ՋF�p0�R✼@j��+s"O�	P�w-�<��T�J^v�� "OFYK$cV��N ��r��5"O�`��d^{�\p��&��d;D$i�"O(�q	   �   +   Ĵ���	��Z$�wHU���C���NNT�D��e�2Tx��ƕ	#��4"�V����c��mZ18�4��YX�ik���pc��(*�vpP�.J#�Ms&���n�.ԕH3>i'�ѝg�h��	ڟ��6-.)� I�
ц-.b�b6�=$�t�B�]���T)ҝa�y�M��9F�ԥV��I�K�4��h�󫐪AF6]�4��7A�	;:��i���� �L�nЉ�f��rZ���'��E.Zj���B��	$#0pka���]���s�<}�g	�Y��$?}R�׹T,uR6�X�<z2�^�����S��e��E>�xل�[��ē{+�1���*H�\c��jt³l@]�2ߟ�~���ha�=�F�2}r�T�d��H���0}�˔?hL� ����7�1�W�ŀ#p�(Fd)��|T���]?�?O�����׿%D�՚C+p4�Q��`�`��;}bT0F����(!}B�ػ�t�-O̴��߁	(!0�H�Q����p�'�|��#�(8%��A2E�+��O"�@�� ,�,�ǌ��5�!�t+�>b"��@~b
8O�@��ں��9OB���@��?e�.����l�&U�|��F2�? t��L>Y�L�1&d���Or��'�̭t�D�I�J�>����&� �~��G�.��^�	bGN�N���!��ݖ{���J��B*|�^�Ĉ��m��a�O\�Q"�qB���O, u�M<�󄄇2VlA����U�����*DQ�	�\��{�M<���(7 �P�t�|b�8����GH=IT<��U���t��Á"Y�I"$�C#>�����8+�*�)v����F���)����x%�qz��bb�3���:#c�����]T.����ŞK��0��w\�y���̛n���Ė�M��i�'� 59�C���DL�Ȫ�BMS�i���gÔ�<U��!�����D0͇\l#K>��L� 4LVy�<1�f�<TL���E�.@�)Ht�C�S�	��'�*x�@ ������`�
c鐸Iǉ�K�<Q*��y��@8��S
j���̌~�<�)�=d]3�aV0HM�=2Uw�<�VfS�0d<p���/o7:�@a��Z�<�J��]3���&��Z��P�c.�\�<ѵ!ؚ{��D:q�\�t��sw�@a�<���F�9{ �яRp�+�&�A�<�� Kx��$�f�c�Nf�<��� m�%1"�W%F���CĬ_�<��a��       c  �  �+  �7  �C  P  �[  �e  Do  *{  ��  �  W�  ��  כ  �  \�  ��  �  2�  z�  �  s�  ��  5�  x�  ��  �  N�  -�  _ � � 4 w �% -, q2 �7  Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�� |d��"O
`�(�;���8���-0��1%"Oj4��ND^[��"3/9�0|H�"OB���H��*�ʞRy=a"O�味V�!X��!&F�:J�$���"O,��a
���C�Ą�M�"O,$3%o�-���p���+Ն�:1"O��ݢ1����`���y14]2��i�<�6��{_���c�H�`�fX�$Kn�<��A̼VI�xR[�)�Ć�pඤ�ȓA5��('nߡ4�� �)˩%� ���,��r�؊b#`T�eT09���ȓ!�b��g��}�8�F��-? �ȓ
K|m�ș�VṔ���2�%�ȓ"R�X�j�4JN�1�˘X�i����̹	_�jZ��1!g��zܶ��ȓgil,*�J�
j�Ne��i�J%b���f	�(U��:���G��$Y^م�~r�� S�%T"���k\�jx�ȓ|4�1�îJb��@ӵ�ݩn�V��/[`�"�v4�R�!ʎ<��M�ȓ`:��z�ؚh�J�Z��$HY:	��H��p�m�C1��!��B:��0��EnjZA V;9����J[
2���	��4'J�EA�IVW&��~�(aZ��ӹ�>� o�Y�|�ȓ�f�A�
Ο7�H��M�$�����mޠP����/���ANXo*�ȓTv�����{ ��-7�*h��I��sB�8�8���3����ȓNe*M�悡;������X�o��!�ȓ'lj�#F�m�+R&;�|��2)n�C��0S4���T:
b���:�0!��e֊��)��ͷV��,�ȓ0�&�8#���� ع�L�����;�P�AFd���,w�6d��r�EQ�( �gVlɦ�M,H��,DP���|�I	$G#\���ȓ"�)���E�B	yt&B�^�LɅ�4�� ��eëF����n��R�p%����I�= j���ML"H^��P�E6d&�B�ɍzD���r.&r<5�f�_��)D�DƘ=#���)��Ľ&�z�Q��Q�Q�"~Γi�p)y�-^��0���,�dn�v(<!��i���!�$����Wf�ߟ���>j��C3�ǟQ�ҡ��� =*!2��ȓ��R`�!]�r-�p�-���'�ў"}S⊣<4,��`��F|�Sb��T�I�|$Ex��D�ˎE�ƕ�AR&@���7�3�y��לs��ۄ䎍;����U��OT��D�"���2Wd�	iyd��ʡ�D,'�p|)�l��Y��M�w�]x�ZM�ƓQ&,��� J�\�� ��+l1H�F}R�6�6�Hs��bd��2�/n�F�F{��'o
m�UJ�6iƅ�ʍ�TI�02
�'�6��F�O�5��˨M�d���'cP��!O�����)X�@Jb �,O��
�8�R�ӥ��O�0��6��2ȇ�M�u
�	��^P�@�r�Тq4 ��2�X�1Oغ@3~�8��@oJG{�<�� ɔ���fR��m��)�t�l݆�A����PGE�Y�n��u脍8J���S�? �����W�p5|����[�Yʺ��"O�@��@5Q�����
���qw"O�����[�\�80#VTƦ��`>O�Շ�	�l�����ʆvzP%�"�����	N?Q
�$\6�*��ͫ3�X��r��%U����	A���L�㈐�h�fUؕ��0r��ȓPb3CLE���[ā������X?��4��S�O�P[�C�x�0e�9f�$�"OܐԈ	 TZz4�ÄN&������A�'��7�;U��l2GKįS��P��K�)!��vc��x��0�6��VM��s!���y8b����2�����&\�a~B[���w��)I�� $�9eH
,�r/0D�`K� 4M"�∉%i�Y�I,D��P���1������z-��:%G:��m?�ÓD�Nl�l�:$#��pq��d1,��uɛO�U��˓�B� wkT �?ae�'���	�G�q�� BgL^-r�<�I㓲���(�V�G�K�9S�E�1)���ȓƴ�0Ei�X�!+QꔦҒ�D{��'�*���7=�� +��p_�=j�'���`��~��K�ђy�Pd�%�S��?��'���SM8Z#P!���
[�<���I�,�p�{@�n��q(|�<�B�m�4y	D�y�Cg��y�<�Pj�6I0L���Q��C��s�<٢���.Y���f�ܗ6��`#�lŪ-��t�=I�S���̢	�
��f�ݠA��B4�ùV;a}��>Y��9'G�0m՗�*��a�Hy2�'.�A��B,U���Ar�T٠���yB�O���ȡ���7L(@�e��fSXC��Ć��E����t��2kJ�(�S�O�\	A�Ǔ$��Y"�E���Ka"O�h;Ц�� B��5�\�an~eA`�x��'������� �pr�_,ٔL���M�d3O���SC�s
9���ҿFL���`"O�AC���}�y+�dT-C�[%�xbX�%���e�i�% ���`���P;�rB� O2O�*v�%Ed�R�a�(fUX�"O��Ȳ.Z9U�P��B�e$\q�S"O�1�gb��T~�9%0!���C^�(�'�ɧ��x2 �?<������t��y�����>Q�O,��C��uUTXs㦓>T�Q�T���'i�y�]=Z��%Q����D�Z���Q�yrhY
&�Z�頃^ �[h�*J����?q^P	�F�;�����<m!�\&8���Q�,[�9ⲁQ�l�_�!�Dگ5�|���9Q�f�&�0]!�d��� C-����P��|tȵ�0Ot�=�OG�D�>iV��.�
�#�O�QF|MٷK㟠D{��I�,\h~�㷯נC
>�S�
�+�B䉓$�ި*f✴g�8HU�½Q�B�In�Xq��♥=`�����(C��hO,e�>	S��pH� C�݊ ���2�[W�<�⎇�ns:s�Ê ?2�R��T�<���I�)T�}��כ@��m�d��SH<a�jO�8��Ś2*�3dQjh4�	%&Q���	ǓTXQ(��a
�W��'aN�I��	M�'[���	�
"^��H#(ڠ�ߴ�Px�g���CϹlj���`c���ē�hO�������ޠ`��5��
E�.���"O�0�\z4���%�1��pq�i���Z�v������m:"�9q��i�!��ay�"˪��0���y����S�? � 1ք�-sh�x��b\�"���`����'ўʧ�6i��֓~���as)�>q��-��V��y��U�c�Hii�a;Z��ȓa�¨Щ[Lr^E���Y�'�H�ȓa���4��G�&�z�$S2/�nh����$-�S�!��Q��D��F�c&E�VB��6�$�g�@Œ��#�j�<!˓D����n�:x--B�C](-}����IR�'�H�#�'h�,�sXH4h��M�N�nD�d�eHV�2
�J���-�_�<�#��QZT#Q�-?�R�[Ve B�<q�f.�!�.��Z�~lKsl[S�<����<	k¤�B)D�bZ���WOS�<I�$.n+\���mJ�Z���r�̇�d.ў"~���\�d8�'�@9(4p����fi6B�ɇM��i���"T(�*��E�2B� ����Q!gPЅx��[2F�(B�z��"o̘5�M��A�Y$B�F R͋�oʜe�حa���J��B�ɿ}��5{�'K
s���"$$��C��*T�ʙoD�|s��E F�-��C�&cҊ�L��"�-{���3�B�I)_i eᤥƞO �廂艼0)
B䉂��w��[���ض4��C�	#/���y�W7fW��S�Ǆ<F,B�I��Y�'ǜT��e�b�B�I P`�Q��P�B�
8���2XRC䉳ALF�Cd�̟
,�3j	�4�C�#P|��XC�s�F�"��ڟOg�C䉅JQd5;�fլ)ht�C ܡ^�
C�I�'28$&�2 "�hҢ��e�BB�I�L����L 9Ӳ@�%��Iu$B�I�0�
8��,�ry2�� 4&C�I�tq��ѣ�0o������8U�"C�Ɇ@͹�BUq�M�r�Ϩ'��B�Ij�}�B@�#A~���f�c�B�!-��q�cH��u��?Q��B�I9x%�����`E0�B��"Ra�(�` 'ʬ�9���7��B��OL�H�&G!�rY�Ƅ̀>��B�ɼ �����DM�l��@W`�qY@B�I\Iu*@��i�B��O�"pWfC�	�)��T;���t��m�R���o�B䉇(��HV&�"z���iדp�$B�/\B `��Ֆl 0l�f
W%#9B䉁N��3��]��ָ1�=[��C䉯5$�m�2��c:�0���Sh�B�I�p]xt�0\� ���� �N?j~~B�I��@a���)Cˁ/	�PB�I��|�Q�M�q~�p`��B�8B��0 p%I�	�U0U�"��'+BBB�ɑ]1�H�4��9,�ͣ��"0sB�I^�N�"k�?d,ʔ�R�J3QAVB�9���A�һ	^|�)��!��b�X�i��./���ƾ!�d˘f�bQx*�/P�Jw��?R!�ǰk��#�Q0y)�!b�ڕ"]!��U9r,�i1"G�	�]H��@.6T!��!v~�z �iҸ���=!!�$ӗN�"9��CF�!Zѭ؛@w!�3k��!��D��g�t��J��!�DX(0+(	qݦ.��u�!���!��I� �Y *�%$���	S��D_!�����&��3J�&T�'��=#!�� ���E�3@	���Q�R��,��"O��.��Q���i���'T��0e"OlȠeG/T�
�[Q�M�[h��"OF4��_�U�l�9C��f�	"O����"�i�C'D�2y���'�2\��	ҟP�I۟��I˟��I���!�AJ�:
�0bl \<ҵ�	��I���	ӟ����@����	�2��X��Ǻ,�<���Ė7�2d����X�I�l��ǟ\�I��@�	��L�	�p�@d:����c2p2'g�eܠ���|��ៜ��˟�	�(��ʟ��I:!��{"ƒ��P���]�~�A�	��4��⟰�	ܟ�������h��73YH-*�c�'F%����}�J��៰���\��؟��	ӟ���㟬���vaPU�a��u�����Y�}����IƟ���؟(�	ş��џ��ɧo�Z��0�ބG��(��-һ#����ȟD���H�Iş��	��L��<�Ʉ Xt��g�G�f)*��F�T�����ן���؟��	ßt��ҟ����t���87p���f�9�Y�#��I��������Ɵ��I��8�I͟ �	ϟp��40Z4�  ���A^�$����d���	���I���	ӟ\��ҟ��	џl�I5j�C�	}�d,3â�9k-b���ڟ���ß�������Iʟ�	����	�E�� ��&����Ǘ-�L1�	؟�������⟔�I�\��4�?i�Q(D��ɢDi�!�ŀ��,_|�r�Q���ICy���O��lڳe>����%V/0�
Gg
9a��[F9?1�i��|��y�Cy�H�ë�?7�D$pw	Q:!�Q'��Ԧ���	���RC�c���.�$i	@7%B�R�Q����Ot���k�� ��<�����'ڧ�ܲv��EU��H��Ijj�P��d�����?��.�M�;Uԙs�M�w>��SdԤ$W��R3�i��7M�է�O�*}(��
��y�(�?4�A��.A�9)�e��y�<l�&8�rD݇B]ў��@K`��#� #ǀ͌+�( �7ht��'2�'{�69;n1O&���ƕ�q ��Z7Z	�K�B"��6����ݦAݴ�y�V��c�N�S=rD�����5�N�B�(�Q��Mn�a�|B���Nhra0��;^����*d�:��B(ކvA<��+O���?E��'f�˓�ލPЄ�cE�Q�uw4���'Y�7�B�����MÊ�O�:<��ț��Q�T�%"΄3�'�6m�����I�m��8��9?� �ƒ<o�yٵ��<h�V�x�OC�������J?���4�����'+(�ܣA�Ĵx� �c�Q�|<��'�j7M�={#1O��i,��D��@l�c9D�¨�	�A�Tϸ>�7�iL�7�r�'>�������ˆ��h��N#Ǥ�"��ޙI�4��@+�>	&%��>dZ%����x����21�˺]���
�+J:.c�-��J�'��	n�I*�M�珀�<ytJ�v^�)�vX������<��i��O�9O��m��M���z���A�=� l���՞��x�Agڳ��QP���\/�n����?���ź�`�~�Y"��H�T�XP	�ɔ�D�5�U�v�p�IUy�X�"~��ض
*h�F@G%'���&��N�>�FNܩ�����=$����! ��͐3i�� h@o��<��OLo=�M��[��	Z�<��>n`�\���<�t�_Q���	Qe:v�X�A��3����4�F˓�?�6��$���������<�I>�s�i�&]��y�S>�X�'�����S4hM�p8�n8?ISY�p3ڴp*�&7O.�
��@�w�N�9�dƛP�P���#��Vv�x��g�����D��9��`jSj�L�^��˄	��Ҡ��d�����蟜���P��?��O��ɏ�M�c-��^��͘�J�~��X�JN&2�6ϓ�?��i�ɧ�O�>!�i�q��lA�c���R�����t�0!l�91	�`�`d`�L�	:�4�H��Šx��'DRh+CfC.p�5��JԪh_����'e�i9nߟL��џ���� �OPĠc���%K���	O,�zk�0Q��4O��d�O�����S���R��yE%Tk���*Aq 
c�4O�Ơ�O@��|�������Qs�@�Γk�f�̂�CO��jEIj��tϓȬ��� T�U�d hM>�+OX�D�O�=BR�*��s&�__�f��$��O���O����<Q�iU�q�'�"�'�$�1T�N"B�4���ʸZ��`�U�|2�'!��r?�&�dӔ]�	Z}�K%7�dL����_�p���
C�y��'���Ú	?w:�HY���3JL��'U��D�t��/�t�����o:Fa)c�W˟��	П��	ٟE�D�'�T �`,�=�p#f�$K;Ĉ��'��7��'��D�O��l�a�i>�]���`�VBZ�G�\}�� ޳ho��	6�M#f�i�x7mJ*nJ(e7O��D�%�|T*�c؃yI|�#&��9d� �RT�J-r֚9�B�(���<1��?����?��?y"D.R�}����h���J��$Ц���x� �	�D�'��	�Ob���j½��=#g�EO��Ӣ$u}��p���m��?�N|��'��A�˼g��I�ş�#t���	=�����P���20{YS�#.j-t�O˓S
@��f�/��$I�OM�w��Y��?Y��?�%�E�S��Y��)�4��Pͻ/H���mڼ^;D�Hq�L"͓�cޛ��'(�i>�ٮO�xnZ��M3"�Of(��A�ߐJO�h�GX{�	�gm��~g����?��G�&�m�!�Ր��Dퟎ��q�? L����'S.Y���-<4P�P3O:�D�O����O���O��?��K�!��0���/=X�:b�h���ȟ�#ش G�'��6�?��I�R=(}b�gK�v��� a�9/�x�Ig}Rn�($l�?�k΍9G���ʟ��P����hr�*�cǨ�*xMӲO�%��E{B�'������2�M�;T�p���O<7X,�Ça�@%��h�4*_R��<����*��h�h}``�"Ä�c��F~�-�>a�ie~6�x��%>���Vo����!�z���%G�\Ya��P�|,4�3rM0?���l�L�Đ �����l@�+��T�����	1)O����<�|�'`n7��Y>��cL+:m�͑�.�,۲��4�޴�����'V�7�F�dS&=JfGχ0�8a�R�,��qm�����  '�����z�&��k�)`�<?�%%�M�@5`�Q=*��e�e̓�?�-O6�}RB�Z8D�(xz�ĝ�P�P(9�%��Λ�+�Θ'K����t�z��N��x��@h�/'��1cE�dδ�m��M�'B�i>Y�S����������7c|���g.�:-",�Â�I/�p�}F�H���]9/Y�E{�O�fJ8E�0���ܘ���!�U��y�X�X$�(ݴg�2$�<AWEIg����P+\�Z�`��I���?yN>�6Q�<��4h��:O"�6
ȥ�Ul	\x����~�*���?���ɜ8�(a���P~��O&y��X!m2	�3OY��7�8x��.�?�b�'�2�'���S�<��k�.�ʍ@�ix����៰:۴Ip��(O�tnZj�Ӽ{ �I+$:)�"��lv�WET��ЦE3�4qw���Z<1��0�'�r�
_��H��N� 8�����G�d�PD>��)1�|rT�H�I̟��ٟt��ܟ��H��`e6au�>��1Q ��oy"�r�H����O|�D�O����?��}��-�|�Y��,�����'9�6��oڼ�?�����*������@�` @�ET�`��H��y�n�O]��#ؤ8���N>�-O8 1coڠYY&����	{���B��Op�D�O����O�ɾ<a!�i���'���7J�Yl����*ķg���'{j7�-��*���MѦ}�4Qq�Ƃ׿\;��hE�Y�Q�fMPQ�$g6�����$1\�]k���D�|��\���m�>4�gdѾd#�d��		�M��'���'5"�'�R�'��ـ�섩@x�-���kt�����O@�$�O�8l�<T�u�'7-�O�˓ �D�#A�I�h����Ħ(B�h��'e�ɽ�Mf�i����B3����'��睺Zq�IYpfԡRQڼP���AvN9(��9aJ�(��|�X��������I��Uȟ��a�p(H�*3$\ � D۟P��`ybEgӊ����O ���O&ʧ_/E�Ʀʪ
�@t�BBT>w�ZD�'�`���giӠ��IL�+�(�+�Ӳ5�����nܺo߬EY��[([]�V�_�������䆵l�re�b�|�%��a�IQ)7�<SG�Q�)���'���'���dW��2޴j�Pmq���3.�I�ƪ 5N����)����Ȧy�?��Z����4w��CV,�� "��Q0�B�sA�iʈ7-Ӝ=���c䟟�#���r��	��"Syb$K� ���kPD4=h2,�EAU��y�]����՟|�I�p��ʟ4�O�x(ӣ��b�p-�VlۃT%��X��`�*5�l�O����O0����ܦ�]�
�P����,�ҽZe$ӊ^)h���4y��$�OT�S�'?�L��+��<9C�=]UT0�&˪ �YʁBV�<1T%��~�M;���%����d�O��Ċ�{DX\Sf�Ĺ,�(��灓+�,�d�O��d�O��9����2�y��' �s_��e QH2p�P���$A�O<@�'6�H������Ŋ {  ��#0uq0<��͋O����OS��S��]qF��<��'r���%�?y���
;�:3�O�E�� 2��@:�?i��?����?�����Oh��U.T�L���2PR�=B���O��m�#Cn�ɖ'd�6<�i��"�	8=8l-��]�"��=2�z���شEԛv�h�0%w�[Ip��6"p�i0�U"7�`Ѵ��a��y�'ܖ��9�6B�L�IVy"�'�r�'r�'s���7 d���	�d�`�pш�剓�M��2�?1��?aH~��t�ꆏ͕d���r��H!J�M��P�$h�4'�d�O"}j��Ի"������&�0��Q�1��e)u͙���d@-FC4q+bT�5�D�O0˓n���K�؀,���c���L�X�����?���?���|J)Oވl�i�L}��#2�qc�ޝz��cL�+R%*牧�M���ĭ>!��in�7�Q٦%30 U6)chx��\'6Y�(+V-!^�f=�2f!?�W���m"E�F���dklQ ]��Ӡn� t�x���>�d�O�����S�vG����@C�&�>U\T�Yt�2�.�M���Ie~��p�v��<�P��7~���!�#�*B��7�y�Y�(�4�F�'�T@0��G6�yB�'0*0���Y�??\����
�P�DB�HՓ���:�.O\ў�}y�'2��'�ؒa���G��.y�p�'�'@d6M�2}�1O �i柰kqo��z�\*��	�`�ԕ��s�O��l��M3�'�O���l
)QD"��U�j�(T���~ͦ� �Q�X�TQS�O��IU���*��7�ğO�4����^D\-Y�瓽5��˓�?y-O1���/�M+��G,�N��G�l��F�N!J����'�&7�O*�O�9O��o�9�:��܊9�j��&A<�
���4�?)b����̓�?�t�Ϻ){�5�c�GB~
� @�z��X�!�[��؃�������O���h��� �ޖk~���4Q*1�5����Ҋ/�	�?�'?����dC�*yZ��'��\�xB�@ 7�V	o���	G}�Oa���'|�yB�A��y���Ju@��
�Rb�d�''��y�T�Cb��Ff	�{s�'`�i>��	�`T��ɂ��T��8³MO�P�D�	ٟ��I��'%�6M*Ci&��O2�$��psF��g,3h�d"��5#��⟔۪O�lmZ�Ms��'Z��\Y���ݑ\�Ryh��H�n�ӟ��e�^@� �Gy��O��H�``R5Dw2�X�Q�n���D6�d�)c].Bj��'���'��џ�ʐ(ջf���T/ΣW�� ��`�Z�4]�X�i,O�Xn���&��f2IXa�O|��u�0.E6�牴�M[Źi�"6�[�>�F�0c:O2�d\�\�#U��a�d��b$��u��+ύu2�Q�P!;�d�<���?i��?i���?��� �'R�Ua�LҪU�.qP����A��`�ڟ���џ<��j��'"�adX=z�P�@Q.4g�4Q%ϯ>!��i��7��֟�%>��S�?=�l jWؤ� �Ғ�pBvm�>A����&o�py��. й���ڕ)��'�	�I�� :GĂ �d\�r#!�n������I���4&��6Z��k۴C6��;�Dx�������sEC3-��"��'���|�O�6���j�j�o�<iV��g�]jHPm[�]m0��E���H}��Iݟ��բ� 2���b�ZyB�O�L֘���0�AK"X��7��?X�I͟��Iߟ`��ԟH�	ŗ�M됍�3�BqI�!^.}�t�**_�؛6�'%��r��Z�7O���Iæ�&���qF�>& ���1NI��hK��?٫O~�lZ��M��?��s/��<��B:N���j��e�)Ky6٢Q(3Ax|�q�ő_�Lu'���'���'�r�'V��Ɗ����#��T,7�2��p�'�2[�`ٴʹp���?������F�6%Iu&�8g����!�!h���'R���ִ�$Ye�',�O���*�%Q�|P�.N�>��M0��M<���`��2b����Z�`���sXx��A�p�ɹc:(�p6a� �<1�� �(���Iٟ������)�jyb��Za��a�v勓�ŏwA��s��=r\ʓ{����'U�''~�Jb���	�ew~���䄲j@2M�Qb�#�T6���=8jM���$񥢔-&XZ�d��Sy�AG=�p8���^�Z�J�����yX���	ן`�����	���O�s�
��S�MzR/�pi.��eh� ��!�O��$�O:�i�|Γ\��w �јC��a`49��u��� lt��nڃ�?�O�)��j�ɓ�g��q��7O0��6�>u^q��҆-���2�8O6����� u�N�<����d�O�$��*O6�ѥ_��e[��եV]����OtM
ǆ����'Dp6MF���	�O��d�@G~0It%ϳ?�T��a���YJ��ON�DZs}�`�rn��?y�O�-IG-�4(آi����4q��U�56O��䕶+xyp�M�u\˓�j(JVvq���l4�dQ"�S�xL��(�ʥȄ����?����?1���h���D�/oBh�#��L��IQ#M�e[�����ص�"?�iu�|�w�N�;�G�:h��^����'�<6Mզ���4sM�)�D
�<���-�r@�w$Q�d�p�" ��[� �`ť����`���!����d�O.���O`���O���&�걘��_t�n�b.|�<˓^w��FƔ����'�R?�d��'�Rk^ Wk����"l���3�jˤ/���(�f�&ja����?��S��ԁYפ�?
W����]�}Y����m�w�'E�e a!��<�5�|rQ�|��z)�6@��fۚX �Q/l��OT���O��4�ʓ,��	��yR�Ѯ�\L�� ߛg�|C����y�'t�⟸r�O��oZ�Mcøi�:�B�Q4�I��J'ʈo2F��#�Q��y��'ߌX�[7(�"7Y���Ө�5�C.&�Yi�W�D��	ؑ�y��'���'�"�'�r�i՜_JP�������΍3V�R��?qѷi^��s̟��lZK�I"=Z�M�T	�u0�$ұ.M&�-����$�צ��ߴ��W�
[�`X��?��G$.l1����mbj|�� �(<W�\!e��	װ��M>1-Ob���Ob�$�OL��@j��� ���<=��[���OX���<�0�i�Z ��'Y�'S�;*lf������LϨ p�#	�m2��A�	��Ms�i���d"�)�����E�չ[���[@��4��:��8�<��o8>���2#D��R�V�XI>��D΄�p�cC�$��]����?����?���?�|�*O��m�xW�T��IR���#�A"���@�Uy�bi����#�O�Pn�;>�j��Gn�%f?��!���) �شb��f/ӆY�m�'.LfmN��eG��n�剣WO�u5�-��ʁ����|���'��'���'@B�' �ӛJ�����%�h��B Q�����4
s�]�'d��	W˦�]�A.�6f�-W��	�eF�M�4��4a�����Ox��|B�'���]��"@͓T��94h��u��y�qh�=��͓_����𭒹��H>�(O���O��`Эէ\�b��D�ڂ`R�j`��O�dχ3��у�I�<AV�i�)��O���'��������iK�,��ڐ�|��'L����Viv�
a��Z}�f�&��l3����/�외�に�y��'ب ��[�� Q����<q��ta�
�ڟH�dΰrq�yGD�eKZ�Q��ߟ �I۟ �I�dD��w
r�	p,M=q*X�-�
����'�'��6-H,��m6�f�4�	�çĶp�L�b�a�i$�@�?O��n���M��i~���*М�yb�'-�l�h�:D�Y�� P�+0�DK�,���D�{�.` �`8��<���?���?����?aa�I"6��QSp%�>Y�>p��hФ��dIۦ�1d�ퟌ�	ٟ8$?�I I3�;^~�ĩ�0Cpx$z�'JG}r�b�
�n��?�H|��'���\ R`�Ex�$�R-�mZC��>x��1V�����
�o
I� ؘr.\�O˓,/����OMT��9ዔd������?���?9��|�*O�n�3A!�m���5Y�$�F �q�E؁�t�$צ��?	0]�D��4}��Km�,e��o�-S��K���WaTH�0m2�l�2�>O��d��n���;Q�
���˓�����hq#rBE�g��`K��]�]O�Y�d1OV��<q/O?9h�恤<
f��V��0hs* 扺�M�Ѧ�@~2�i�����<Y�?�̄bL"�&@���J"�y2Y���4]����'?b�y�j���y��'�b�� �LF]j�̙�> ��
���1v�@ ��V�ў�S@yr�'$��ħ�W����GZs��4H�'}�'��6�=]�1O˧Io8A�(
;S�,h���Ý����'v��}��6�m���	_�S�?�.4J�F�Q�M;\�R��J�V��S5F�*5(J��&2?q�'i`Dt��iG���)r:�$V�Da�pRG�U�4�*O�d�<�|�'�6ޢH�R(���5-h��DH�rG�-Zמ��)ٴ�?N>��<��i����6%��؋Ђ�:4��Qgy�"��8��4O���M\)��f� 9t�ɧzѬX��̪ �,	aI?4�,b� �	yr��(T���d����4!��:�*�P�4a�b��<�����w���1nv� �GxB�l臄����mڞ�Mk�'�i>���ɟ\��g@�KR�	�  >t�@LfJu �dŢ.���=	T���Ħ�CV(&�������'���@�O�q��vhE,?�6H���'�RV.��9	t\��ݴbO�U���?���9?dL�Rf�T���cUG��y�����$�O`-�'X6���������J��I���;b�X�z4 ��'��r���rGh�6^���Ce}�����s%^����³cbT0���2f�XD������D�OT���O���+��c_g�ءc텤#����ӹ�?�׵iE�ٱ�S��Jش�?!J>ͻ!^��0N��eZrB���BJx�j����g��nZ�T���Hs�,��=T&�Kq�T,*J1�̆mE��Y��/D�1��g�y�Ioyb�'&��'���'�2&�(-�>���
<6�nXS��5TP�I �M�v��<����?!N~�t:�hk`P2Ò���HմztTu�Q[��P�4ś���On�~�i��6�Q�(P�/�b(�G�6KƜ�1�=A��x�,�<�rN��w��b��K3����D��l�da�w�	&M�����IȀ*Wb���O ���O�4�4���Fj �)�G�3s��рq���qĩ��yR�n���˯O�Hn��M���ii��{F�t�6+H)\��5D��*�~�H�'�e�q��!��@W%{,�	�?�1\c���)�HK�"�.\�1�ͭVZvx��'�2�'�R�'��'��ڹb���,z.Ah�BS7�>�qD;O��d�O��lڵ;l�IܟH�ٴ��WD��$�R6n$�x!�1[��0�u�'@�ɛ�M[��i���B�>]��H��'�2�H}Wx�K��8X�nD�qGS�]��D8f�ߢx	�����|rZ���I̟P�I����rړy��P��/,l-�Kڟ$�	^y��|��I)"=O��D�OʧAZܛt��16���iֿڦ��'��4��6k�Q�	C�S�?I�g��9I�xӃm,B���q�֒�U$ϭ?�� �'�4�ދ ��`��|��ݳ3���&�D��nq� �P+qR�'z��'4���X� ��4c�H�슋����1G^�hJX��t~�����:��\}b�h�(�d*�7�xx�4�q!@�x�����޴6�J|;�E��<��.݌Db�E޶x^d��*OtQ�E	��r�T�eC�7�,�2O���?y��?���?����򩒏)��=9�!��@#��� �4#q�l�'u>�	ӟ4��d�Sџ̳���Sf�("�E	���>SS�E?�F�k��hmZ���4�*�	��1B�	c/�Pi�ꭉ&� ,hMz��1K��$ٚH���QCEV�`�O���?	�)8�]���
�p%P���fO#_J ���?Y��?A(O��lڞ��`�	ß@���b�d9��OT�_)ܸ��ʇmS%�?yFU�8�شۛV��O���=.R��݅s�I: �ڙ=u�$�O�]x�%�,���d�<��'E�te�Cf��?Q���*V��a�K9V�����?Q��?Q����ß��ՄR���c�B�"&��i
���韈jٴ{Mx��'{f6�4�i�y���(�2�E��|��Cv�X�شy��f f�p;Ҩ��_(�$�ODİ4.	>-�0}zw��_����ah_�R�b9A��\�ȓOd˓�?����?���?i�v�H��`�//R
�B%o�<���x-O>�m�y�"��$��V�s�#U!ߌ[��a�M��fzr�ׄ��S�i
�1�� �ЦMBI|����ꣂA6]G&�g/��p���;V�B&�P��$:ڠ����	]̓O��I�P,b�nV�n������ �ZE����?���?qsC�I��f^�T
�4�~Lλd� �$����Jƅ�\�%���֐|�O���D)�v�bӠlڑIA�]y���)Xj����&�*لɖ&k��	ޟ�30��i+EI���wy��OG"�X	%x)-�cT,��
�O���T�I��\��՟@�	O��pOxdk�+��K��Iȑ��4�>���?���9Ûr6OJ������%�8*�h]!.#X����1at�P�n�%�?�O-n��M;�'R���qSe	�<��YE��� B��ʀ�4���!sgν!G�L���I� p��0�$�<9���?A���?ِO˖����%Ƅ�V��E��?�����d�٦-ʇ,k�P��ϟ��O�*�v@]�U֎!���K+n^ ���O �'�6-��yH���'�
Q� c���s����hi� �5�huA�h���l��+Ol�)ײ�2�3��!��ڕb7� �F�67C��#!-��.�8���Ot˓�?�|�,O*�m�$d�)�A��p���jtB���йHB6?q#�i��O|5�'n 6��M�(��&���EZ�C;�YmZ�M[���j��͓�?���vz��X,��D�]�\�h�D�Sߦ�C�۷���<���?���?q��?�,�p�2�����+7�U1!�T�x!*�} ��c������$?����Mϻz,�`Z6;p-k�O�pd��U�i"�6�Mǟ�ק���O&���ٷ_�Ȩ�'�B�V��R�V��S:mٟ'����!��]�ƕ2�|�Q���	�����
% m�S�Ɂ�J��C�W�������	iyb�e��9�4OB�$�O,`JfT�`�25����K�0dI�"���O4��'�H7-ᦱ����$�7����͊�Ks�h��a�g����O@ع��]pn4�T*�<��'1�!���Y)�?�&�� vO�����E:�lT��R��?1���?����?���I�OP�ZBe��l��{�ɟ8U��p��O��n�y�(�'�r6M>�i�a�'Ͼm�r1�V�8c(Zp�ҏu��,7���nZ��M��g������?�v�3>�P�z�q�`M�(|Ֆ�0qkٍf#t��*�D�<����?����?I��?��+��=B䍠�hD(Qz�䈒%ٲ��즩�3og�8��ݟx%?�	7C0��3��V�>���Ci,�0H�OZYm��Mc�'�O��$�O"d��R"�@�*Ri�3M�p�"͑�N�X�S������f�ʭR1eDP�Hy��^/�D��@� C�0�1��Yu��'?��'x�O���+�MC�K�<Ahҥu|�a�(�<��4x#��<�1�i|�O���'9�7�Aަ��4?��=��G#B��� ���?l��I*ƇE�<x��Γ�?5��3G�&݃�G#����T��"O8Dc�6� ����E B�|̓�?����?���?�����O���b*�*zIC ��r��M��'�b�'��6M�� ��$�O�LoZ|�	�l�R��c��HE�Q*��F�O��e����������޴�*�hƕE��8ϓ�?�m�=�D�g�H�<����
kܐ�I�oM:~wv�IO>Y,O��d�O�$�O����ܿV�6M��LM��U)�K�O��D�<9��i*
$Z��'���'����O�vR�c�ln��p%d߀.�Tk�O|U�'��\k$� >D��*���Q	�4�9:�I �Dǲ�w�C!i�(5����Q���d�>twF��7����耩�ēJ�JX�bcӌn���pꈑ.8i���'nb�'�r���O��	��MKW�(�@I[Ѥ+VS�}�A�$%t��'p�7�>�	���$ۦ���81
��;�+"W,ܔ��ό�M�i�>�ʆ���y��'��(���ܵp�P�q�U���G�غ�"�"Y>���R�`�P�'M��'-��'��'���["��[7����d"���:(�4j�4(�BΓ�?�����<����y�bG�cz0�9�Q)8j���O��Bo�6MGԦ%r����4�v�i��iЕ�O>y���8rkX��A��8��`�gh��,<Y�u�0fQ�$&O���?��M�x@���E#��� �l `����?����?),O�8n�&���	��8��?��D�Q.ǈm�fH[�� Y���?��S�D�۴1����O~�-��$
!k>j
`�b��:6����?�� N��T4�4 ������R�S  �۴1��PـbR�q�n�r��+	�lr��?q���?���h���d�[`P�����YSػF��_p>�$Ŧj"*?r�iib�|�w�ָ�U)�z��Ū1$
C1��I�'�p7��ՑڴM�<00�ƅ�<��3RPlf�@�qm��*��՘zoB�"7E�J����!������O����O~�$�O������vJV�x��C ,�!L@ʓy��f,�&���Of#|��%K=X���;�_� ���80g���d��uBڴ��T�O9��M�03���(B�p�Ġ�V��2N�T3�=��I�u�+�/(����|�[�tIgJ mfxٱb�;-�j����Пp�I͟���ɟ�gy2l��Mr3O�|ôWxxf�"�L�223�	���O�l�O�i>Ѫ�O�n��M�½i��Yj�i�r��E�I�>( UX�#GS�,ٞ'�Rl����r��	�?��_c�����!tq�	K�ᛸB����'�"�'W2�'���':��<j�N�-%9"`�@�I��mM$Kdb�'�`r��A&ɬ<	v�i�'-�� ��2��s���9*�2ђ�b�O �:�֠���	]�L@X5O��$�4F@��!k�w��ERW-H��UJS{�Z�S��7��<����?����?	�#@D���
A�&|���)�?�����ͦQ�������`�OqL+ GD�X���KI�:��	��O��'xR7-�ۦ����'�F��>m�V�r��A x<����O7V��q��[�T�*O ��X/I�b�z�+%�d�S���5�H�]��8��EF�k�L���O����O���I�<Q�i�P�G�P�,�  ��#9�X�"E���̦��?a�[���4
�޼ c�
8� KШ������if6-�s��9*����1��1<%`=XT�AZy���(k��`��b'�P���yr[�����`���$����O�X�7/S.L�δ+i��|4�Eб�bӆeZ������s�'rV��wH|X�D2fv<P#aG�"[�a��n�o��?ɩO1����C�W� 3�� "d$�Z�&�: $$�Iq�0O�ը����6X|h�@"0���<���?��#@�or\͚�$�=V� 6����?���?A���DҦ1p2�~�L�Iɟ�
����bd� .�;�����j��_[�ɛ�Mː�i��$�>1$���@��J��=q�Ms���<1�ri���P��=*U(�/O���]��L!0�:i�w��D���w'�!T}��p�"O �Z� $F]�1�QG\��'��1d��"�2� �'[;�,�ML	FHz��ӥ��U���� �?�d��'�%q����)GȌ��OIRʉ1Q���"=xh�w���d��9W�.1ӲI��~���KƅU��m��m>7����J��nHP@���3CȸQ��7P�.>����&I�L�X��$X$����X�-��$mംL<A���?�M>���R���j\qH����&��i�RgY
W2�'�R�'>B�'��'P�P���C߾qh��9~2&,	F%S�-�Ob���Oz�O`���O�EYbN�� ��ˤ�ի4}<�j�-�n��D�O~�d�OV�$�O����O&�[r-\�|��A�▨xj=�t�ԦI���?����䓹?��	�`�x~��a�!���j0���b,�y�F�i��'/��'���'��1�U2��D�.����P�B�"r���w\ul�ݟT&����ݟ��Q����\1u�S*����$#9��1Ra�ߝ.+�%Q#���S:���Hո#{�)�������&#�j˒�FZ���נɉ3!�D�  �h ��{C�Ċ���s�`��
����K(Py�8�����:�t�e����S�R�<2��H�↋Y���ڦ.y;\��S�[.w� ���/��W�:�p�D��`UD�@�e�J�%(Mc�0ыP8[�p$��,�: Ú �&������?k�a��,=P=�@��Um��%bJώ����?���?���x�{���UQ�d@�Z:A�RBJ�\�A�cQ9H��G�zb>�O�[t��	��i��߼f���S�UpV�������r5,R��q��'ؚUїė�L�Qr����R��F)y�
�'��\���|�����'j�e��d��=6�E��,J��0b�'���/KȠ�S䇖#n�0��On�Fz�llӈ��<Ɇcí.�@���v�0T!@�}id�:�e;�?����?Y��!���O��dv>�8fM�%"�\�shM�x��1Ai�w���2�d�(	�L ´�'�@I��$�D��2�K' М�dB^	qw"  +'��(��$�3�?9t�ϼ2p��!>��'\���C_
xt�axХ!zKF�����?�Զik�O^�$�Ob��Ѧ B���=���+��0c��#D���e�,^"��y�[Kۘ��4�>�	��M���DG}డm�ٟp�i��F��]ǔY�́�06(P���OP�ć|����O|��k��(�'kD�
S�'�R�9"�:PV֩����\�	Ǔ=���8��Z:����O�Q��ȕid�Qw*�7�h��'V8����NS��`ӂ�dZ�?2���'@Ȩ]81��N&D���?q����m'�5R*��e f���

�XE{�Ob�6�;c��`v�NT����	��K�����<��N�=0����'�V>)���؟,Z7,��F9�!�^��	-i���O�8'��B��x����:Rܡ�R����4T>Q�fe�1�����O�r�JTyЪ*}R�S=ļ����[�J�"�`���M��(�:|��0���z�)Z}Kp��Wf�6�(P��>)3�՟(Y�4|���'2񟮤*��5	&d���6Z�<����O���(��|LŶ&�>완
8|���;�O�hO�IV��E3ݴ��2�^��e]T��]��\,� ��i�b�'|��Q1ҼT�%�'!2�'���wf�3ѫP/K�>m�H/L�h���@�'%�
E�%M�h��z�˘�g1�LM�Of �E���	r�(k��� xL�P"bK�j���c�*g�����&�5��v�~�����$j���*x欢aDXcI��z7
�.*�ڴ|7剻PX����'�B�'X� �&@ �h�e�G�YpF��O�x�N	�W���)fj""��h┟�Z���4�ķ<1P�5͆M���$]O 1�c�ߎr���#�*���?y���?����.�OD�dk>y�I!C�n�@#o �N��qI!G�@Ā�W�H�� ��mS$��0��$U�]���hv���l:+�:o�:��t�L�7N2A袭X������ w����D�l�xx��67��l�P��l��4kdᘷ\���$�ƦIx۴�?.O�D'��6m���ծ�]�8-hsh\%tC�		w����p��>6X'K�)
�b���I�ğ��'�$��e�b�e����@rD�?ј]ڥ,ҏ�%.,5(����OV<�ŉ�Ov�dw>����3HԠ$���7歫��/=q� ���51�l�IZ�güD����>"L�9xg���~���*�T
$��d�r0�y��V�<���JE ޡ8@��DD�ظ'��\�T��'
|��j�<<��z�jF�G�^�`�'�0� �H #��) o�+=H&$��'w�7M�
p#�LQ5�F�)�2�ؒ�Πz�6�ObŹb��u�	@�Oab9v�'&�HP�	�!_�� �u^)yP���'�"��i <5 �%��8DhHPg��9i���'��)�0#��kg��?>�tHD@�[j�G�H�����
�`P � }��y��	Ǻ�aJ���t� �h�P2��րM4bm�4�Ǥ�� ���d�O���|��䤱���y*f���\�l���{���O���� �����n*�yʂ�A�g�I��'y�#=y7�ߍ}�(��(;.�Z�!I�x����'��'IBM���\!��'<���yg��QǬ1�lβYyl�r 'L�mԜ�i��,���(0,�w����q�dΚ	ynQ��N�j6HɄ��� �A���T��E�MBV�9B适0
�'�^���|������;/�d%��F�Z�>�q%�*�M�U�iK��֭��,O���_�`ޙ˴��&1>�E����YJ��=����4Z�xZ1P�8&84pč����M�Ʊi��'��I1��OG��6?璈��FJ
�xx�W�h��h�'����˟����Zw+2�'��E�3&��B�U7z>|��6U9�$dκ0�uX���p=�A�I�AJy���<�c��)�d�Մ��#��p)=\OB1!Vn	6��D3��L>�.K�	�/^��Dm�&�m���L�'P�dj�ܙ�%�A2�&\���á�!�px���Qߦ=�.=�t��F�1O���'�	9JlىYw���'�e��L1ĊA���)+�D�E�'��!��n�b�'��)ݩ)u�x��|��ޮ	�>T+����m��-2�ʚ>�p<ab�Q�~
t�&�``�!�63T:��e�X]�  Bc�>O�T��'��'R�vFT�yb�L.�������I����?E��D߾a��y��X(�,qA�5�xB�`���K�F
�,�*�*C�M�E�&=O,�9�������?������_���dM�f~��g�е^���{�JE9]�����O,m���4,Ȳ�7-B�P^Lu��_.���R>M��"�w}j�!�c �8c�4}��J�s.J��Ŏ�2r��dk�A?�pȓ�G�;Y��\ϧcIb%3�+�*L�Ƥ2&� f�}�O�IW�'26�Ӧ���e�'�`8�E����d$CS� 5�>h�<����<y���*~�~T� ��	m��YRB�c�����>���U�C�p�8��b挻[�j�
�Oz�d�O���7'�+�����O��d�O��; YdTCv*iK }���]���	�y�	��<�w��=�
�xBߘ����eEJ|�o��T��ɘ^)���A^l�l��F�S#���M>�C�Fߟ�>�O�=rC�D�@.nx�DL��~&��p "O,h�dIF�B}T��Ԩ��+�n����T����S�&B���{.�P�#��(�)�a�?K��H�IƟ|��柈��(��>�9�R-+�H�c�7<~]�0-W�	�A��&� -�qC�嗬:��c��dЍdx��bg��4Z���8\���d�E)8N� �%j\,R#��eis'b�4&�`asÔ��1�C+`6
����*y�����O����O^ʓ�?���lߔ+y��3��l�ʣ��>�0>O>a�i	> �����W��@V�]�ya�6�';�Ʌ-����4�?���jy�)##سi-�g�Q(q�����?Y�B���?y����*L(�9��a\(MrY�!�
/r�+$�Ɉh�U �͍��^Ի��+�p/� Ack�U�E $��=�=���ޜA	��9�A!$��Q��;1�.����SnB��[�b�O��<�1�S���j'�(e\���LG�<Y���?a����U�9����V;I%����1}�!�d�̦��E�=Ld���t�H������'��@8G�w�����O��''ٖB�)K~l��O��IQ.I���	����?ap�ր.�v���S;K�왣��2!L��@�t��SSX��D��1+֡�����E�8�v /7 �����P�D��' &TS|��1�X���$�J
�!a�0hV<�s�>�S��q�49n�6�' �&(�Y�Q�@Cj}���ɢK�1OZ��,<O�1����Tt��/B��G�'ih#=)���:&�d� #�"����nĺf��k���?��B|�j$�9�?���?���h�NڼE��h��*�3吅C��D�xUZ�M�(��ڒ(7�+k:擬��Q��[G��2�T,r��N�vB%(��٣N�������*7���B�a���O���E較�J�W/�8:V�G�,%F��3�Q#"���K�<�ޟ���?U�?��Lh�@�w��҃�Vb�<��߶d���rd H�L����t~"
7ғ.~��'U�%*�:���ڠ6��P��%7?�C�I/&9|l�wK�O�d�`vdN3��C�l$<a���x�(����Le˔C䉃#�����Fp���Pb��G�B�INಭ�n��"��&i�7}DC�	!_\}�&S%)��+a@F�z3�C�I5s���-�u:���FXJ��C�I?SG�I����5�ڳ� .(�C�� 9`xy��
�O�Qj����_�>C�	/XjHđ������{��>C�bx����낑kY�uYb�U��B�)� �J�'��
�G�8�D���"O��H��|Szq������@�g"O���P���H}X�����zj�i��"OP��KA�Y/��%kV1G��<�"OJ���͐�!�1�
:�ɛp"O�� ���~Ўe;�I޷9}Rٓ�"O �i�.3�(���	G>o��� P"O���gl�@X��ߝ����""O�1��׫>4�<�1(�.�"O\���һ.lt��mҢ`� \P�"Ox�(B��a��;熨_���*1"O����S(U�Ld)�`Y�q�Hy�"Oz�*�̂1�T0��6A�b�r�"ON��E)0V����B)�5l&��4"OܴJa���s�f10B�D?m`6�p�"O��b��	�n y�ŝ
S����"O�0�Lܮ��v+��pC0��"O�1�-E/~Y���L�=2� '"O�4{�g��p% �iAj\P"O>$��a�5t{TVc�E8\P0�"O�<��Z#V���T�֪
�R� "OH�������B�4}|-i�"OJ��J�BS�9[��R���"O���g�؞�Z,��T�;*5Z�"O����l�%Q������
)l����D#Q]P�����"��͙5X�T&-�ShO	Gr �6#��?���@�i�x���t,P�ԉ���18�pA�$G�u�H�ц%T�(�\��K7t�r�[#��:-�Q���']���S��A��Fhr`d�9dB��4g��%W�Z��!@R�P!l�M���[�Uj�ȃY��:Zc���#ß3\ޱS���?���s�N'lO~����E9����O��N�fu�	�	��A��G�W��e�O(ā��6/H�֡̌N� �2�D@�<�%���>�\���!��}��#@"�8�1t�E�N�����DP���O:��cDE� ���(���~�bG4OT�
�N�"�< Å�6�:��g�	�&9^m�Peā/����"���&	j��ŖȰ?ц -r�r٘�Ñke<L�� -��� S'���p<�4�+��1Y��J���gC*����I�f���A�8k��	����+8�-C��
ᑞ�
#j��I�xU��
� P��>AL_M����Rڂx��A�L�Y�'A�t�� ʹl�,����pI$�C��D6���t��n�i� @�*�ioZ0<N\y���Mr�I-	l#?��CL�g��������j�����[?A1OΗV�8�ZPc�'&����%��S�'n��3B <[r��'�ޠdi䎎�}���?���T,.y���a�ݓ�G�B�jd�% ��(�1RL}��	 R�L��p<1@��"j�H��#N�p�&m�i�-+�CW�C��	�o�v���_:�)��0;��9���
}�I�☘�.�Z�	�'J$��P u�~�%kuD\�n,ڀ�>�p��c�c�¨`������Ny"����$�O.4"p$�=q�|ZČ<?�"=�u�'� ��t�ɺj�uRa"�6�,Q޴�9[SHݕ�LŢ��S�eJT �=)g��0�yre�0@��)����J�i&�_7W&�D�2�ɚE�T�&�t�um� ;ў Q��T�D]�U8�$�+bZT[ 0E	LI�{� �� .��r�'	��ra�2��i:����h �I��c�`��,AǓF'��Z"=��Iz�Ξ�����K	 (�%�'��	���Oӧ�O�fH#���(�eO6ymʄ	�S�7Ҡ�Dz��1�v��/��v��ѡ�;��$��y���u&�_�X���/D��� 	��r����E�������^BŪ!�O|����8h�J��b���J�̊P�i�= �I	q�L�S�K��
�:���]tB�P1�T:��TE���+�O`�nZ3zr�P�il�h$�F{2��#�U���,<��x"��9Cp8�� ��~��g�S�~���e(ڗ'ª�{D]�q���>�p<R��Zhr���) ���A�ضCft����pTqOr�	u�d�|�Zb�@$Q!F�+u`P�����?[�B��8�EE����D��yy�Cۿmm��'�h�yV�P�u� �"��G�&�������I���	rO��Ft���K�s�v�Ϛ�XA2��p�J�lV�[��
Hæ�QFγɚ̨t����On1IT�D	��Xs��5"�h���E���u׈iR'
ہFJn0IP�4�Q&���̈́ *7�0I�\�
�L�i	[џܲ�'��	0�2hyЅ�=rd�0���S�3���%��G�H܅�I�Υ�F|�%q�(�t��M�S��
*1��)��6�	u?������OE�6�݂Ԁ �!�F��\{��9��X��P ���ɌVG�@�f��}{��d$Q#/� ���ɑ/31�yk�@������\y�1��?��'k�DQ,z�^�XD'��(,r�D4�,*HW���q�&��46��V���5�R�ݘ�&��O�AL.&�\��� ���I'H@П�`�E10���
F��4�E<ړeH͚���*%8X��ߌs��%�T�Č��O���4�	z�" ��4b� ,��i׍{�� �'%i�pA��	����!��n��+D�Լ/ǔT�AO��&V8�b�&�Is����5Zy
9q h��p1W�_��������HO����Ҹ��ǚX���aU�P��;[�b +�E�:��� l!�I=�M��%kN��1'�"�X�o�,��|�4M:"�������ګF���m��	�@�v
���]y���<}y�"?�3&�9d��sf�K��8�����:�6�\�?NL|�dA3�Mcb�~ݹ����Xm�D���!/"�	�G��M�nY�ѮX�q<Q���*�@���p5�
��xr�3'��䨸y��i<� z�RN���{����˂�U%H�urq�U�,�.��G���<��"AG����&�^My-I��(�$���"`0u���I�d���Y�T�`�D�͋io�x�҂�>
�H�k ꝅQ�t4��!+�l����T�F �XDW(��y�Ʌ@B`�Z� �'2��T�-U�Y���LP�*O.�ƲG��dЖ-be��'��z�"6Z�����m[	w���x�'���@ql�.[J���o�/~<q����m�F�kWkO�><$�ǦΌm�DL�����%IGv�f�jW웖7#ўyQ�R}*<��[>��+�K�W�*����sx��� ˦��J�;Zx�����-��m���Hx����jޑ����i�tȪ�3dٲй�D,D���  :��K�hQЦ +'�g��B&KW<�,�ߓA�l��GҕC<�"�MF����I�N�$\;p�Cb^dC4�Y�/lb��y�n�;qN��ЅԶX��eIV!�z�||�P�L�+�l��J�$��1����J%΅����yM�!#(��/�tx6��"0�����	��'2=@JX	)��h�D�S:�<4M�1,��Oޱ��Ģ��ۃSd��I9G"��wi��� )�+A�Hi^�}z0b�'��X�AB�8�j�ҁE���0	`���H�F��wGD/aL�b�NN���dU�<�Dܹ'��p&N0V��#g����4��l��C0>�YI5�r�iH�L�&�?�qĖ�t�1!�e��t	�m��K^�lXJ3� 3�6h�	'�f�8wʙ�;84��+ �66mʬXgN8t/��|��i�&��O�m��݄y�����W�\ˑ��0�pxQl�+q���b��ו\I8p��WE&���	5 V���
L�dh�@뛙RY.Pd>��y?���u�`�'GzL˧K�l���_���@�}Kr1����:8�d#ǓBY�,���w��pE�Y�^(�@��l�,���>��FA
ve�e��5���ʧ"��1��/���	w���p��>�"=�Է	� s��NQtd:Wg�<y����(�B�Tzxa�Mئ���'�~AC���`Xԁ{���Z(��4��`���?yߊ z�U���;=<�({&l@Ӧ�YH_�J5z���6%O�j�gyb��~y�$�UA
, AW���A�ߓHX��Y��A �sу;t1���%��퉦(���.S��j�*=�F���!ݟ�0�(ڬ&(B���c���3��}�E�ќ>�]�$�xR�X95)���A�J
k�u��BR�ge����	�k�(�oz�Ir�e�	Td�����-�0+BGڦ��DM�A�ae�ɌH����H�Э�e��W�t�a�)ۑ����S�\h�ٰI~�Zwr�Q�J-U���y�c�!@AN�b[H�>Q�B1��{�k� �N�`��W��0���,����e��+�>�)�v��00��8߲��䚞O��}��dl��z�$�*>u��8�	ǾN�� 2��>�uf�=�C`�S9�%D{�.�'�*P`Q$��O�b�BY�(O�$÷&�Z^*˓;,��'*�j5���^����P�yo�m�����S��%�'	�K��~��"��7�89�+*i;�y�-�\Ax�ӱ���	4#>�1 ��	�hT�<j�8��N���D{"
X?´Q�3}�O�)���
�(�z�a�HR�!Q3C��"H{�1F|mO�z�H�3,Z�0�p��!O�UI�	�H�8&oˢEV�7홑j�� �"ЈO��ٶ`��;��7-L�3n�D�oA�9���w��<��}����Ρ>W���w \�s�ڢ=1g�|0"�)�#-y$��\{}��i�I eژ�S���@[>IA�	�t>p�+YP*���G�;���J���0�4��/\��Š��OĪ�x���h����'lR SbH�B�
��쉂B��?B&2A(6�Ӻ�%A{���+ �LI���_?;��\�"5�a(�Y� (?�'�?*r�N�Q��ٝv�	:�����d���~���"��֐���d�=$��O0���ስZ-�\�B�
�):���i�:�R�����0��9O�Q�FbZ��y���D��"�',��)�����:�"��tOԻK�Bx�V�Z��$�

wD�3ړ~A�ɐ�G�^�D��V�D�&Mta�,۱L�~e�a�O�4k������Q�����q#CT&F/v(9B'�� ���>w�Dd`�j�r8�Pr��+�Q�T�D�HTb`ϧ=p��a��S%;�N4K�O>샏����y�`?�8-"q)B�6r�JuD��6B6����I.���V�<9&�\;���"� �"@�� ~�29t�E����;$�	��M;@�
�|�d"v�ʫ�F8�;)�Bd]�Q�pX���Zց�q'V6-��)�,�����G���S���	���'#
���n�N�⥘ҦW)hn*�8�i֛F�Ø8����Q��
�) �ʚ�hORx���@������+|[j\�!U�W�� D�J/A�X��=��`�'N��"w��A�~鲇J/��,�H2g�A�<xEh�0�P����WUP�pF�J_�@�5�|B�Z,_
@���u7U�/5cÁ�C��{C�`�f����	$<
���D�́c���L�\@�'W��5b�JM+G�r"�ۗx*2%qA�LC�U�����Z8��ŀ3A]���s��:��ǙA	�aB�b��V��}Ke�gӜ�:7 �hT��"F�/)���q��ݗ	�ѹƬ�#]��S#��x��6�:W��q���j%�gϴo��>ړ(;�p#��;��3�Hh�;�lG�]���D�P�]���h ��;��O�S�'o��]b�!����!Z��x����V�P`�4���w�x�C��|!�LS���MЈd����T��H����2�~�7E�V�6�'9Er���Γsd��ħ���$�ȓ�F��j�Y�|�5��1�$l�ȓl�A�c Z�~o4�+�h��J)B"OԱ#d/�6 �69����nMz9"Of�3F���^LU:���:�ɠ�"O� i��ӨD4�򅪙��r��e"Ofى��ϖO<j��	���(�"O:,bխU#mT��s��_cR4�$"Oű�g��?�f|�I�"^�H2"O��᠊>.�0	��IL�OZ� ��"OЭ	�� k^�1��V(]J�0�"O~-��@�*WD�p��M+;�L�"O��w�L2>�I���#��q��"O� ��$ѓ%(^�:0�ٚJ�2=�"O�=@�GLh�9׆C�P/�P "OjX����(� �Jg��C��X�G"Ol�Jg�!¾��t�)EL(�$"OtxYh���d��5G���"Ox�p��V5��P8�'X&�"O�a�p��%(�i�1�H�%	�Y�"OH�e攄b\Z͈�� ���"Ot���z�rԸ���2��H#"O�[�"ȢYi^T	��Uq] Ec�"O�� W���[�D�"f�Qk�"O+�(�?O����5��;TV���"O
�96O,%
��߆�|�b`"OVĊ���q&�@��B�;�b��@"O�X0'�$mpP���C���0"O�p���;h�؈i��R�tq�IxU"O u�s�X�h ��g�	EcV<��"Ot��ǯ�+D��9�u��1K��1�"Ox45����{VH�7a�,t��"O�ᰕF����ǥւo�4P"O��C���3]��$A�&�*!�����"O`A؄��7�N	p�&��Grd�
�"O�$�tiA�i�������y\�j�"O�(�PKN$7���X�%^{V2���"O8��F�@� �RԚR$�7Pȕa4"O�L�0�0Y�u#��&NRuC�"Ov�Q�-ZH6��� ��+?��n<D�X�N�f���àm�&�q��.D�����_g��퐶��<ޕ�r$,D���4��+q�H�@�L��@�.(D�d���G3Jh���G0�5��!D���0c��P��MS�e	\��d >D�t��l$�m�PI�>8J��I�:D��0�YN��4�/��r$�!i$D�˦�J�N?~��U�R�:MD W�!D�X:T�ġi"�,����	R�Ԉ&�?D�L���ԁ�E�fִ�1�U�QZ!򄗋eo�B��B�8�ɂCݜ*�!�� �-����2u��EӕG��V�`(�r"O=�v�/�>��)>�:��"O�C�O�A�5�ת�x	��"O���C@[?Y�������&��d�"OvHs���\�:U3���%Q:|�E"O^5�O�'(�H(��$�=4�f!�P"O4�r�a,x�zH1 d+�\s!"OI1l�b�	��C�a�B�A"O2�K���<<�Y7ȕ0�|��G"O���LӱS�R)�6*�o�0���"O��ۦaǳhZ�3h�_뺡#�"OJ�P�N�|vΗA�e2���y�_�\�D`��K�)�:Ȼ�(B)�y�kҲ3�%IϞ
�`yQ�+�y"�ϣ[�f�k�"F�jW��y��e�DH:RG�U���/F��y��	|G�Y[�(UB����?�y�kY�)�4�B�/�=�29y2g��y�a�7�d8bH'RB�+�@�9�yҮ�\������[A���y2�<{g�4�AnR�~9��SA�Z��yB%v��|
���"�b9�@�ޠ�y�I� ��|AV��+mo�d⢢^6�y���2y� +���sjl]8�)��y���81*y��E��j�.Tq�Ώ�y�&��DA��"�!_�f\~�!���y��ޜV�*�(0��tv̬��Iʾ�yREϛz�"}*�O�n�p�+t��(�y�G�#HF(Ȇ-�a������y��
*=jE%ՋYn��v`�$�y�j 2��7kU>T�m�GK��ygU�bV�� uƑ$Z�Dx!����y"f�Z(����W�V��'�_�yO2^�����/��R�<9 5ʆ�y�W: ���GNڸH:%�S�K?�y¯[�(� ݮ8.ڹBѦW��B�I�|z�r�e�[��	K l^0r4�B�	+8I�p���A�P��h]4uQ�B䉀�3ێ��jڤwD4��`^M�<��	���uK��i$���HB�<yЭ+S����	�v$�"M�|�<S,ˆL��LAb��%�tT&�_P�<	ɓ1\>�C����)ڣ�D�<كǗ(<����O�� ��o�B�<�	Y"3��˱�F�i�^qx�/�S��p=�J�]~0�J��=ᖤ�gFPH<I��:�&|0jңIdi��≠!!��~��p���kA�E�� ?p���G��4$@�2+U�o9 �Ձ?�y�aKcb�k�J��d��p��J��y�gO�琌i��6_Y�`����!�y�f��a����O�m�J��b�yBH	0-��e�0�)g�B%�"����y��Ԯp��A렅�+���1b��y�&h�������o�
I�"�	��yr�1{%2���E�n3⌊% ��y���6�S�j��kƘi{�3�y��)�'.�Dcu��8��y��*V�L��ȓ)@eJ��R0,����®8�t�ȓMXp�BB' �U����2ECv, �������5J��p&����ń�p�'��m��&O�t9�U� ��}�ȓRBF��2�=W��h�0Q4��ȓi�}R���K��XI�b�/4q`\��S�? Z�p�j[�[����)q�೒"O 1
Q�K�|8 ��m�HԀ!��"Or�{D��8|�V�׫}�ܰ�"Ov|���ČI���tMÍhM���"O� �%ͺcUL(E�О6,(3$�'d�	�ozt��0o�Z�s��("+�C�I0mjب#�$�� +0!�'.�C�ɒeh���c��!�4������TC�	#��a���Ċr�Np Abɹ,��C�Ɍm�4����[({��� &�<��C�	�M������!�l� �ѻ3��C�Ƀ�J���L ^�^��E�óc�vC�	0m�<�j���Wf�[D��m�B��3Ik���m @M�]�dj��00ZB�	`vY#Rm��C˒W��ܲ��'6,(�e�
9
u�
�"P��I�'-�]�rFT?u�Ց���t#�Q�'�(8�r��r�J-��mZ  ��D[�'�h�R���C(v���߀f$��P�'ňRG�N�������]F��'��9$���>�L��W�x5��'L��Y�F		ygJr�]�|��p�O���$�Y���ŭ�5;��Ƌ=a~�T�ܹ�/O���d��5#���J D���tM*Yp���B��Z� ��J�O6�=E��.�n>B�3��.Hq���蛦�!��K�v{��x��p�����	d!�D	0�&�����'g� såW)p!�$[��bI��_��\��!��|U!��ѴI�f��nS�'6h�C2?��� D{����]�L�T?$���4D�p��Ç�;��ӓ(�nO\���f1�hO�S�ౚ�k¬*�lM"g"Č�C�	 Y��k`��"�fy1l%`{&�T���(M |8�iԤs@5Y��/r��B䉆<<5b�Z)j�q�N�L%�B�	�K��_a@���(=]zW�'��	�E�5��B��=̖��'f�(��B䉳
B�Pq��+�tT��B&cS�B�	)tjZɩc�ѣ8��dp���B��� �qC��CZTҷ��>08�B�	�4!��(�A�2�:���j�!4FtB�I{^5A��[�V��#��O<�C�I�{~���sX.Oإ1S,B䉁�� �t�ƓSe�U�Ҁ�0u8C�	+[Vb�;Q�X�o$V��3��66�XB䉫7:��A���bR�3A.��L4B�I�{��8�Ѻh�={�拚20B�I's�D�fÚ4N_�${���F��C䉩pf��q��|8bL��F�VÒB�	,I���&c$(p�G�
.�8��D#ʓM�z�B�'jM�)�gĖDW�nr(<�a'�!�Rq !�;{��<���w�<A�Oqo���v$�:L\�e��IIw�<1@ ��$�4MPQ!5���#��~!�䏎����^	����Z�B9!��x)n�+�ӧ'hbiqp�/~,!�d�=�0��|����Ť�)�!�d��k����P�D�#ˈ)��"�1�!�$�c�|�b��?�Z�2��?t�!�$@��:��@��;�4r��
l!��"%b���f۟���C���K
!�E9�� A ;�|��ƈ!򄂬��`��Èm��H�"�"葞܅�)� �	����"���˄h��d �h%"O0
t虞A�Rm�T�ŐRH�	"O �Ф)Ґ\%Ҍ
��y,��	�"O�	��	�b=�����i$��6"OY��-��te�����ݚ�"O����E.=J��Eˇ\*��"O� z�N���N4��-�����"O�]9�@�~�tQB�i�{��E��"O:�1�Ú���j�JHfTę!"O���HϮ`Q���� bx�3v"O1�CMW�1d�S�h�L�tUD"O��9BI�6�<ĭ�X���sd"O$�*᫉�]��XiU� n`��p"OꬠӨJhpEe�H�4���"O �S�O�	}qH�*Vd�@���A�"O䰑��Zor50Cɏ��fAV"O�1��l -xxX@ f�EWE�6"O>�%��osA3�W�<��C!"O��"�	Qf� �6��
63�� #"O ̱1G�!
R�G^�=Ş��S"Ox1�!X c���_�f��4���yr��o*ʙ &hZ�/���A�[��yҨ�x-�D�$t[�-�2@$�y2�Ҥa��r��
p~�0���8�y"ܝ,/�Ȫ"�C�vj��8ǭW=�yB�_~)���NԍxD��� W��y��Z?)�/�"�$��k��y�'������H���)���y2���P����)�B+@�+E�Q1�yr�-�xYQ�*�8@��IB�'��y"͛�%�H�ħQ 8.��8ZZJC䉓7h\�I*�B� �zC�H�KC�	2^@L����4qy���F��1;$B�	,}9`.�;DB�85���>�VB����i0�$^)���V��A�B�ɭYv�d+p-U(��u��U��B�ɋt#T협-")��,�aj�2H!򄀆Z9>A�ϓ�<x�g&�.hD!��	���Y�gF�~N�1�d�5a�!�U��tm�&ib5q���Gv!�$��Su��hT"��5wTh13��b@!��(]�P�T�N�^�t���fR,0!�D�l��jfhҰ��hTO�eH!�$�T�b��`&CF�"�J���+P!��:*f.��ς'c��a9�ٓ*H!� �� 
��T��(�`�B�=S!���WD���h��|��\ƃY?9�!�$�q��e1��&(@^p�X�"O`�F$U�B���������p�"O,�5G'y���f/L�1��|95"O�i�0��4��>�|kҬ�BA!򄇛a�UK3料(�H�%L�
|!�dP�X�D����ˊ�D�SP-X)~!���xV=���C4QZD�c+�8u�!�d��Mcޔ��kS�N��Q��#�!�I�i�����<]&����(|!�d~�C�U�K��p��M*V���H�"O^\���Ne��I a���l�B"O�����v.���� Q'�x(�f*Op����#,l������>k�7"Ox�X6I�&��P#Dϋ'�"�A%"O9��D�pA�Z��!`�jt�F"O�"���.�|,��X�F�<��$"Of��0�Q�� �I{�虂!!D�� h���Z[�x�E���4�`"O���c�R�'*X3E���Or��"O�x�tl�f��e�Teу>Q�(��"O4��De����r�cĦ8�tE��"OPQE,
.C�lA���A�b,�0"O��+4A�&lq�����5%�T1w"O��@�H"6�$��ì�-�r�"O���m��MPZ0��H�
�B P�"OjQHd��"�.�y�$ݳ]��%�A"O\q+���b$���#JE ��Q�"O4h��ʓ"�^q���B�"<b�"O|E3EbK�1B<�#(�>Vא�`�"O�U���ލC���G΂s��v"O��2�x��lp5�_�x���"O(�����L��'�����8�"O��)a�o>����[v,�ZW"O����+���}���0lL���"O*�s+P>���+&uP9��"O���/��2�<��I.T�Bm	�"O��Z6O]�da���e(��8��5x�"O����K�7(rT�@p@�*.�F�j3"OVC�A��2'T��6`�Odz��"O�(�0��8?^hmRVз8I8hSq"O�iB�б�����L�AЌ\Iu"Ò �b��6v����>fD �F"OR��q��e��ŒvΑ�Jq�"OZ�&m�W���p.�g�r�Q"O��b���/S���ae�[����'"OX�K1�"�l҆J�q��q�"O,e�'#�;3�h�rèJ�0vJ|1�"O�)!��Q��0�c��o.��"O|�J��ї�,X��QQ��!@Q"Oh� ��XF8d`�O���q��"OL)����y�F���@��ֵ�4"O��1�H	\zy����C��A�"O(�	�J��z .�Q"/N,cؔ�I�"OB�(�[))�]R��H��D�*O���@-�$X;h��'�e��@P�'lf-����8��#�h��YG����'���e)0jΪ�0�΄�QW����'blգ5�[�몉	���:�=z�'�`��`�î ��x��i�9V����'� �c4jO�J�[1�Y���x��'}��D  ����eT�Q~�p�'L
�Q�M7q���(�)L���-�'�01�%¼Q�V�z�!��CQ�UY�'��`��:�ɩ��ǅ8���J�'����i҃\��x��1hq3�'��DZ� �+t��Y�-�/YF��'5����
�� :S��6C݊8��'jv�nB.=��� �̒.oy�X��'�I����?�&Ts�o��2�p��'��� 6je[�Qr��>1W�1��'����n�\t2�֪Z;$FJH��'9�\@�j@�/7�����A�����'�:-��*�"g:��ԃXb(T��'�5��� �v*�<y�"�!v�C�<I���$/b�s�jź/i�l��E�<4	ӝ�0��`!_(��RAm	j�<����g��ȑ-˵\���be�]�<�# Ӫo��p�ɀ�:�B �r�W�<�&��5eX��o�/m�Ĉ{�{�<!7/�o��:w���:�P��{�<����H��bˍS>��7�{�<� �+"���1��H'c�=c�����"O��
2.ԑ�&x��B�qT@ZC"OZY�@��kH��P�8[X���"OBK6��2����b��"@���D"O�Fꨄ�g�G>+(ܥj5iP�p�!���1u6~$҅�߹Zؐcӧʁq�!�D�v���e"�t ,0d�L�h1!���A9,`��!ώ��LCT��Q!�$�58��C���?��RR�F�u!򤉢ff�QR񯎆L� �X��8j!�$	 7������?���;�D��=y!��u��\q e	�8� 8�p�P�E�!�B�Dq�ikΔ.�n�	�����!�D�q.�Ts-1�i��@T <�!��I����
�g��B"��*�!��|ab�B�E�B�b� �!�D�wj��0��G (��\�aӑn�!�.�,���-��v�`����^��!�K�c1|��Ҥ��P�֡J٤-�B�	0^I�Ȃ�H��Px�ٔ��YB�B�I"�ܫ��� {&q�怟�2�rB�aZ������\6�(Dƀ�ǜC�	r;@L �)ŗJ��`�V�:*vC�	->��JK����PlC�I�v��%���T߄,S�"��|6�C�ɈkuH����3vL�s��:��C��~�����_�&�z%[R!@MK�C䉅>����#J����B����B� J�,�R�"W1*�X�@+�#><fC�	��ѐG���|�bǥ��q�rC�9%4P��@�W�`7l+Bh���*B�	�VE@�2��:H�d����B�	'\�P�cUH
)k|�3��X��B�/#X�D��"M�$	��G'+ؤB�Ɇ
fp�����3T��|aq�Z�CDHC�	vB���&	�	hӓ֑lƂC䉞^�rPj+Ӟ~𠌡�U�.F>B�	�`#��
i����NLˈ���'�2hQ��i����G��5_��	�'��T�f�\�R=��n�/F���P	�'��2��i2��F'ԍ�ָ��'�6\Z���4��1���hj	�'�h �G8���Bм~�8	�'yDɩq$�%ox�Y3$V����'YP$s� �9W�|�:�ݺ~�z-y�'w��t$�M�ꘒ1+�c� S�'�`�g*٬B���� N3r��h��'6v �IU�bm�D��k���
�'�T�:w���4\j��\�h8JA��' (����%(tAxF�$vL09�'c����9-R�:1 E ���'$����L�lqqՋ��xzK�'�� g�#r����
w��P�'�T���% ���J����6�3�'�vHʤ�7p⤌�#`�� �L}��'�N��5J��A�rQ!���k
�'������7L����(O#Y�2�)
�'����мl�t��q���}�\��']�����V8"
L%i2Ϛ�w�4D����x��ҳ�G�!��x1gF��y��&D�I�׎ؘ����fւ�y�	 ������6.�zQ�m��ybd��1�|��'Ž7vԓV�G��ybE��n�<E��m×Vz%і���y
� <Ac3�V2D��Y��E9Ѭ���"O�X�3�T&oô�34��a�4QK�"O�-K!ȓ�=d����F]�E�Bg"O�T���*H/�L�#���j�"OUS&�n�+��d�>�S"O\ys%�ЈY��ىb���F��<�G"O�
�J�a�P�%rl����"O��3pC��q\IK�@H<B��y"O�0�Ҧƭ�N��jH�H���:�"O�����@h�=���Us���"O 1eRI�٫%Aی[�ᩒ"O|)p�E&!z� ;t@QS"�E"O\���ʎ�:�
����&S,*R"OplY�n�8k��	�UfL�cK���f"OЕh��RDUh�RŊ�#����"O�M��mѸv`�m�䎗M�<H�S"Oh�w�ڳ4H���A�0X��L�"OF��̿Wrv�A���R�;"Or#Q*)Z�P@f\s�V��"O� ��R! �e����zq"O�����2@���#Θ�S�8���"O��9S��@bT���K�Q�Z��"O$�Hv`�)S��T#���	�L,p"Oڴ��B��/7Z�,�2m����"O�T{0�9�h@���ƖW^��g"O��V�2jV,ѓQk�A&� r"O��PcD
G��� 툾P�,j"O�i�#a�w<�,���J?4M��c"O΀��d3g����!@���L��"O��+�F��T���r�ܞS�Ԑ1�"O��� i�,�P�� @<;���qt"O~<�@�V<ft��*!��Ȱ"O��lNE���Ѵ� �c���"O�u���} 8��&=����"OD5��:=���FƓx��L"Oܝ�q�[�"�X����>U><�S"O�A8�璐v��������t��a"O�B��Ŭ0�A�'K�<�@�"O:��1������0;�n�"Oh,�)���-�<�t\�3"O����,�x��ѡC^�h��A
�"O�D����,4���ҡߨcz�(AB"O���V��.�n�K��z]x�"O�1���6�(� �J�2���"OzL���qk����%{�b  �"O~ 9��Y�r�Ȓ�&�<��`"OPM ��F�P��eE���<��"O��[!EճPSn҄D�%h�\��6"OrqH�e�2"Vأg�	�z�.�HP"O�$��45�X���V�gS.��t"O��x�iG�T0��?0���b"O����/i"� �`��0�İ�"OYX��Y
�|��H�s���F"O�2%�.g��10Wa�F�>�V"OiB�.�PqvE�/xK�rd��"OT��rlֱ���S�R;���S"O�$���Ҩn��iQ˕:]�H�3w"O6%(]>6o���/�؆"O��
%c� xhņ"!���"O:�W��(�#`$M�Q��P�"OV}J�	S+.�Ƅ�~���k�"O��RC}��� ��v0K�"O�i5鑚j�p����C+!�!�"O��B���y�(�"�Bm! F�g_!�� "�9w� �31|9��fX#QZ��%"Odݳq��xx�=��c�;���"O��s6�I�u��u1"�&=��B�"O��K��-)|���ʹs
�ˆ"O(�c��./�LRG�'e�i�D"O����4^z$(��ņx�`��"O�u:���_��!���F1m�L�"O2�I���p�x�1S�� m���"O ���:;$!葎�`�����"Ovt�AH�u�֭а�G:P�����"O�����0{�(h��_3F�j)Yv"O���E�	;r}��\w��3"O@��Fb��E���c)�_��""O���$��,_2� �"�Y5n�`"O�Ԑ�ϙ�k�ɱ�N�B2\1""O�xc�!��<�D)�d���s�"OBA[qǂt��@{�!��(�ā'"O$���C�F�����?�j���"OL-�b@of � �.)�[�"O�eI���B���k�fT2��A�b!�$?*�Pհ���QшQ�'�/v!�Z���V� X��2E���e�!�D�!Bc�= ��0*d��/ߖ�!�T���)#oÇ
|�r �T�!�DP}1j�:�&���6�S�$7H�!��ӏ�N�K�l@>I�p�@�/o!���
��$��"sHt|�4oN�a!�dFj^�"��J�C*ԥ��Z4�!�D�dĈa���:K ̄*FF�o�!�$X�T���p�d=Lx���UG!M}!�D�>�P! ��Sk���W,�!�:C�@�Pf�%DQ�¢z�!�<�� tL3������+Z�!�dF2D��h�$��/:�!�d�b�p���N�RgKٯ�!�ę�}�a��1H�M���Z�n�!���0
���)H	&�d��	ڌ|�!��Hsw����	]?���hZJ�!��5�RD1�ŀ�K�.���FX��!򤔓X�)J���wӠ�� �X�!��>N�7�D2�l,C#�d!��e����C�Vr�(ҝX!�$�)�^��g� j�P��QV!�D� ��4ؔKY#6����T�m?!�dسS���Z'|��6N��&�!�DĜB"b����>?�0�7�!��]�N��+Cƌ��x��uH�+Mk!��ݸ}V&P��aĮ �Y���;!�d�5|y��J��N�<��Xr�&.�!�d J��ڤ��.e�������!�$$Y��K��܇^~�TӅKU�{�!�Y�O��u!�Qqv9ZMT&o!򤙺IL`�[�O\I�xH�Ϥi�!�Ę?a&0,X�`�'qC��2U�
�y!�$S>&ɜUk�-��r,��@U�C�z�!򤊟/�I���42�P+v��	�!�Dύ7�.5pO@3*h���bV(CR!�@@1�U�9^��Wb_)�!򤏁�bLS�a��mX����O�0�!򤓂+/$���ĉeMVD��	~!�d��X$�	L2La�4��#ay!�$ڛ!%���cŨH ��Q��[""^!�$Q$[�2���2��c��eO!�d%KʕK���-��kBu�!�� �%�"��^�&ˢk��n�4��"O�X!���F�䈲i��i��t��"Od@+I�87b0�f���,~��u"O���S	�Iov�'��Pi�"O�#u��PFĹ����7Wܲ|Ӆ"Oʙ���1kUd8�$�/� ��b"O��q.RP��B#�P�s� �zu"Ot�@PKK6d�b�
��%gz&EC"O��ֻN �Z"�_eL�c"O�-,��Zdz��ߛw�Q��"OPa���@�K?��g�E�.��`�"O<�x@��$��Yi҈ K�\�ɢ"O����_�pۜ�X�)�2��U�"O��vƳy�(L`�ꏵr��23"O���J]��I+��҄8�x�:C"O��Y���y�L�
a��a�T�XC"Ob8p��1bm.�`���S�h�"O��Jf��>�uYR���T&l�a"O t�椚b�*�*� �2o�eʧ"O�QS��8C����*�00�"O�u1��٬�����D9'�tH�"Oր�`"UR�܃6c]�c�<4��"O��� �*�L`��"-� ܡ�"O�P�&D�͔pS��0��5je"O�L;��DM�P�
̇{���"OH��� �+#�09�T �~�2�Qv"Ov�)PG�kr`����
B/�lZG"O`� �J�n] c�	L�h[U"Ot�ˀ�R=d�xсb��=/�Yۧ"Of�"⓶k�*#Z����"Oz4���Hl ��4,�+g׼�;�"O�l�	Ғ&�hp�c*ĥ�5!S"OPIK���~."�s�	��Y��ڥ"Oe���;+���q�	�)��x�p"O"}@���R�n-��扅n�t��"O�M�F�x��Š��I�*�����"ODEk�AF�N�k�	�}0��Ѐ"O �p�i�<"m�,�H�z�T���"O����ٺrz&�Bu�U�3h�Z�"O��ـ�F�GN$��E��8UJ��"O
���/ԎO]B� ��0E��y�"O��2tE	x��VJӗ����"O�X`I�[皼yr��m�
��"O>1ʆH.�Ь؄�7�ܙ�@"O�P˒�K8"QPHS���'z	"q@"O��
Dڀf������ݤt48x�"OH��S9�x�c���k�0إ"O�Ի,�~�2� G�P5-R���"O\Y��X�zm�$Q�䕦W�yr�"OB����m���s#�a��\��"O6�;vL��,-Qe�
��%��"O<%��,Z:�|l�Aa[��&���"O|�(f��Lz�`�c`F�,���v"O�yD�
�r~���W�ޕfW��"Oļ�Df� z˲�2�(E�B�"v"O.yca�������],Ij���"O��sEY�#�b��(E�O 0x�"O̼iTH�O� �au�d��QP"Oxl�%��^�>y�
��D���D"O�H��(��6�S���>M�d�:"O�}��śQ�8��	��8Xj�"O�C#'�xv���W�qȂȹ�"On��%�,U�f�r�ͅb���"O0$[aOD�]��b�ЉQ8`�ɡ"O� ��1b��N��(����9-U�0"O����:kJ>���
�u,,�P"O��yV���a{.I�� ^�ԙq"O�UۅR�D!�F�R����a"O�k���;(Iy�'Ҟ���"O�|	��Ԋi�p��L�=� �`p"O�ī��W;:Jt�s��"p
�B"OV��֪���Y�qa�2VV�9CR"O�����]���:qa��pD4��"O�]�#�,i����ȿ.�@�*O�a!��Î[�֩oF	Z��
�']�4�5��8���q��7�ֹ�
�'�r�!C)E��A�w�*l�
�'��bɑݠ�b7B�$~�xx�'�)07bӒE��"��P�l
�-3�'�9EM.ol=��J+f!�E��'h�AT�+Ҟ�cgO1^L8Y��'3z B�
�v��٣��=U��y��'�30�&G���hɻI�`|p�'Ab��&HP���vJ�x���'�t�%'�F�n��5��"KL`�'�H�1�ԁ\`d!V�^�}��@�'/&x�#�	�lVZU��J%r��'��c%�+�buI���<㔁i
�'G��c���R�VDY�� ����'�XIb���7uFQqBkD�=���s�'#2S��G�.<����dȂ(�����'#�=�v���*b!�GkP�v�i+�'I�:E-°h��١"S��
 	���|2�ӴZyx��<�*�êB���C��9;�Ƞ)�i�3Zz�U�� 1ΖC䉳t����.�#! < W#�~pC�IZ��`��"�NE�	��8��C�	�w��� �@�`
�p B�|��C�0,���T� � �9�̖9�0C�I�gF�Tr����1��B��߆��=�.O�#|���2�� Y#E��C(�� aCH�<I#�Y+� )*�ݛw�xTZ���<Y%&ƋF�Hy�fiJ�/,I"D�w�<	%CFT=&-�TL�Y�j�yCM�l�<�'�d=�e��V�"�0��&��e�<��[�C��$ڦ�B�E%��x/�a�<�v�O!@Lr�p�2l�8vJGh�'�?�;G�#a�z�Qlr	C�H�"S�!�D��fD�����/�|A���ױ9�!���>M���R�Ȣ5rbФ\|o!�	�F�@0�A��P�$��Q�Ԩ9y!�[�,���k��	H�Fᳵ�"R�!��;E�.\���݃n�� B����O�!�DT��x]ie�H,d����2f�c�!�ԡ��y�wlˮ��xA�
&�!�Ĉ�y���עK�P���<g�!�$� at�%�c�I�}ȵ�^6M<!�䊬&*Xm���;D���RPA��NX!��V�"�Pd�L�Bറc��C �!򄌹�H�k�숋/p{�I�*�!�Dƀd[�=��Qf�G���Py�k��5S�I����jq[��.�y�	� ���F���D��F�U;�y���6+�fa2'h��u0�D�"� �yRH½����׉�o�`����ݝ�yZIeܹ�e�*\pT0���e�(C�	�3|x�_9&p��F^�`I�DK�'U�I��.�4��ͻ�,�,��(���� X�MJ =�z�ѦS���"O X��4vzH������Pc7"OX����u�^Ti2�ȁyt�D� "O��S`̷\�rMX�����{�"Odib��1 W�DR@ �%Jܴ�k"O|�;�B�Hl����$:���xq"O�P��JΉT�8)�ӈ[
�8`�"OkC�ʺ,r�ж)=�ze�"OM��@�: x@��`IV�b�T���"O���� �>s\�����V�S�"OL!c�`�+B6L5�2��%Bx,d�"Oy2 -՛\�������K Hsv"OX!�����B��Z�I��}3Z}PT"O���@��M��Q�&T�n+(�A"O�D�$�#�>�R/ߏ. Ĥ��"OB�9#�Bsu��%̏�,��0�"O�`����Oڀ�3ƪ+!�@t�""O�@�7� @x:�����m��"Ot��C���P�� b�Z:�9j�"O�;g�ܕ_%�|��܄3�����"O��@��.&ܲ8p��֘ dj�3�"O@tk �יT�}�6�K�2N����"ODEP��5,�.U�O@�gB ��"O���s���X1f����J�=$�B�':XC��n�`A�.�4��P�'}D�����-j��l@��<'���s	�'�4�(��k��L:�E�!�|4�	�'"����Ӧ�Ze)[�����	�'+t}���^�4�=���(Z;�<��'y�������?\>�S�C�d�Lys	�'H��$�*�"�k#�O�&��_\�<�-�(Q�r����	�2���C�X�<	Q��|Q^`2����C�P�:�.ZO�<��䈮{,��a���"󮄒ІN�<I"ձ=F����5� ��1�K�<A��[���]al��wn�M����A�<!n� *v����!>�I!�HI�<!��<=� ���O�������M�<�6"�u]�l�`�� �xӰ!�F�<)��D�q�6Y��D�.�@�0o�@�<I�G��Xھ=�di&-Df�zp��V�<I1	�	`�^�����0p��ċMSh<!Р�{-���$��;JQ�j�%�hO���i).	���d*)E�BQxb�Ӌl!�d:9�"gχ��E�q��je!��
`g��x�ɝ�TȞ<��� �>x!���`(̉�3,H����'�F!���0��h�O�?�~�h�Ǐ�!�<PS�Qa�ą8C^�`���+!�dB�tF>�R��0.�<��K!�D ���!婀�~?����%_!�!�ҟB~r�
�`O�L�CDA�i�!��Ђ&�h�fNK�m��c�' �!��S��Vh߼mz*Ё D)�!�+�\��#��*x�x��iT!Y�!�$L �Ƚ��a�T� ��g&M#S�!�qN�3Ac�2� ȩT��U�!�O'�0I#V*ʹg�ܽrA��!�֋B_ =��m�3VK(�EA�:�!�V�B�B$��aοG��0����bM!�)k��	���>.��cp��!���,�� �.| �/�
k4!�dR�+�8A�ȎLx�!�S.ػ��T��"�i�j̝Y)�M�3��29:B�)� �qC1�%&e���pj�>��m��"O���G�-V�$�#&k��e���U"O<�9�(��9���#�L��%�8t�`"O��*2��!M�qᇥ-�QD*OhIΪ	�@Jȕ�q���'�f��R��3x��0`чܐxal9�ϓ�O����Stf-
uo@�mz�d�\�H�	t�S�$��x����>4�mB�[T�؀��5D�$83
��0Py�S#��xC�Y���>D�$����w`@w�߾o���Tb'D�P��%�M�-���R6k$��r��&D�@�Gٮ@LiIf^+ =L���8D�p�G� b"�j�\�e��|+�	,D��8��߇5�&��7\�",����O���d4?�IQ�J�b� ��3Rp^��%bIR�<!Ə[��P�g�2n�9b���P�<��P�Y?愚p�&X�L(R`�[I�<�0)�H�cG�� r~űJG�<�M�\I�I�� �P!�\�<q�d�<�Pp��@�c� ��`BWC��l͓?���5�Z7v\�K��F�CAX�'���i>5�'�Ju���úQ�6����͎)�<9�'F��
C��|�Z	�b��,{,�`�'�&D9��Z�5A�i�,+��x��'XZe�#�B=p�  V,
�(�k�'�xL�i]������@�����'����[''eDP1���,\T��Y�'�N,S�ȴf6�S4��V��Z���0���R��Eh�rTh�����"Oܑ#�lق;��5��-Z�r�q\�@�'���c�O��D`��ގtӊ��eM9��x�'UM�3�,t��r�I���0Y�'~���U�-�LX���{�1�'��V��:
�Y8RFB�	�0Q`�'&�X��#_ 
Q1R�7 ���'�՘&���Ĺ�u��
�'U*׈݆T�q��@�m�ڥ
�'���u��)ZM`���k?F� 
�'�lh��خlt�p�%vH
�'�Tt#�]�)z��B��8@Q�@q�'Ǻ)�4�Zwf4���a�M��h(�'z�( �ة�	qA�B���'b��妒�)Q�ۑ�� H��P�'7�w�ԼT9�@;��<v$r�+O�˓��S�O�t÷`�|o ��$I<Z�D8��'�
�1��?�h �@��a�RJ�'t��i$/��j�M�4�E�QON�s
�'�h��o�9k���P�Q
N�~����yB��B1�
0a�����ĥШ�y�+��U�K��>�mh�J�k#B�ɏw���bG��%���A�	��D��C�+@K�%۔�BPJ�1p�㍃u��B䉨k��{�'C9a�����F |�B�ɱv/�;��n�*-��N۠] �C�� r�\�'����XQ��ؒe�rC��Mtt}����4J61r�՟��g�	{���4Ȃ�"� x	��A��u��yB� !��d
��}b������D�<)*O�"~3"ʿdY`Y�M׻(� �#a�P�<Qr.VQ����%�7E$H�ENM�<q4m׵=��%2rŞ2h�.�S��m�<9֢�=e�$h�@M��ͫ�,�M�<�2�X�01��	�NЯ(��{ak�Ky2�')ўd�<	f+΢!��X#a�]��#5�]�<� n���P�y�v�bk΂~��=���V�h���Ց�ĭ��
SN�n����,D�h0�N:c����V�OnWdi
�F8D���7��w�P���IB�@�A5D��Zcjӯ{5>�C����5,j�@%E3D���R朶� =j@�R�q�8hQE�)�D�<��]`h�+\<=|fq��!j�T��ȓJ@�YQTAŠ�h��4�K�iPD��H����8]9�8�K&|�eð��&"?\ņȓX>`�2e]��K�B&G�`��@T�X�_�U��+�C֪�Їȓ&k�!�!ÅZ��x�'%+s<���I�'���RT%_	B��)hġ�O]�� J>���D5?����1eX ��3��/$l<R��@�<�'�JY'i[�-_������Łe���?qÓf��A���ݴ[A�8u%QY��ȓ.M�H�L�_IM�i׿p�ʄ�ȓvZ�,���SҘ�Y��ڄQ�1�ȓ#����.�(ޑQ�?)~��`�R��Ʀm�-1��X�s���ȓ�
U*w'��q���Z0�ن�P^ޔ�Vd�Q�=�g
J�:��Ն�HBnm�E�S4;Ĉ��R�����ȓ\��Hu�T����K�jԳ&K�x�ȓ�.]@b.�X��t[�C�1zf��ȓ3z�0�Ҧ
���eD�+~x�A��K���Y C�o�]�PC�"8Nx(��{kX�� o�&?��8y���'6���ȓ�,d
��Z��J����j9��B�F`�/ ���&�͎��ȓ#�y0�'5��L�G�
? X���Y��T��$�'�T�Y@CM�<Xt��_C���"V�)p`����/*0�y�ȓ+�4��˖�Z>��`�(��J�І�G�':�M�� �p�E"�+�4��g"O`0v�
�>�yg��Q��E�"On@���'m&�ɳ��׽7J����"Oz`�@
I!^���J1c��@�"O:��� �8q��H�f$�3G�d�s@"O��Ճ6`�^x9W#߹.Ԡ�O`H�
R.�.Lq���2]�b#�6��0|�� ��^w��W ��w&���m�<a�&_6�H�n<>ٔ���P��W��C���;h.t	d��
jjl��>D��&l^�b!�)���Ũ%S�@�D1D��Z/�V`����G���4�u�+D�C���g�(�	G���o��T�$D�Li$FU���0Á�=(R�[U7D��p���8%�I�2Οz�]���/D�h�����r�^x� ��*rQ �za�<	�r��l�'�A�	��q���yٶ���&�&dyW�!J0HY0cW�$8�܄�o1�}�v�ʖM��%�@�ٍ$�5�ȓ{�A���@�Uj�SaD5b0p��ȓ0ߔ)��-@�I���]���c�X�9�hU��`���]�HC��2r�\��"U;5�AwG�0�%�ȓ/��C��;}��EɖB'�L���
������F�UQ��R�B�����-Q8��L���JG/ޠ-sTa��u���$n����e�v�^�9��Ȇ�	��tS�i�PNքq�	V(I��s6�����B���� �Ҡa7����$Μ�Hf�D ����A�C��L��S�? A��db��RCo�H�S6"O���jp�j�� H�d�x�"O\�#R#�)��13E>LʘuP"O����C8S�,��!L��jM3
�'@�Xg,�0K�j�n��X9(X��'�\���e^�H�����W�H�*��ݖP:2 x�ӆ hb���b�!��ʾf�z�U�r�Z�V#&�!�$��}���ÓJ���.�4!���*3���2"�W}���Ђ�H���
X%1��@�d�3����y@
	������9sXʥ��2�PyҪ�:Ah� ����qDꡊu�[c��,��ryrd�� d}�v�B>o�ByZ�)]$�!��(x$YYD� n� ��.�l�!�A*Ln�y`�	U'PQ ��U�2�!�PJ�����,Pr�k1iھ_�!�D_"|�j��d�D�E�̜���Ƃ �!�S��z`�`*"լL⣧�~)!�d�
�����c��8�p��H�����5�g?QU�E T\K���/�����h�'%ɧ��(˂D�T�hKeKǥ36�a �#D��I�[�	�R�:�D~B�¢+D��a���I���h�/�{�XhS3�$D���tA��I[��i�%/��A�PJ/D��r���b}�2��p������:D��E�������88tU8H;D�@�C�&\��4 e��lDN1�խ+D����V�~	i ��c�.}��*&D��1c��K�҉��IS =�6���$D��W%X�3P�8��аZ�])��/D�0�fD(@d�
F.�d��S�&-D�[�a/p��� @(��fx�g�9��� ��\�I{y2bՕB4R�ဈ�VU�e��EU�.!�$ݳ=��T+5�Nv62���d(!�̰�4���ˋ1GGd88�J$�!�$�ef�)3C��\� ��D2|U!���?t�����~�2����-PI!�DAX�=��U�I�ԡ	��ƴ|,!�Pd<���E
�)�ҽ:��5���)�,O��	1��Qs���E�з��)q�B�� r��5�Ci�k�Hd�D���=t��O:��7LOΐ#�)_06�����>d���"OH��cdŲS\�8QM�O5�x%"O�d� ��,����v��0u.l���"O
]P&%�&��d'�nq�"OE�%^�8h4T��h�3\����d�'=�}~�G��N�l�`n�E���:D.��yҬ˼02X��P4af�m�Ȇ����O��D0LO��8�n<G��q��4=ւdA�"O���g�7:�2@��Ǎ9����"O
��,+�������<�����"O���&��*'n*�JfF�pk�M8�"O8�	�?��!�e-([(�h`"O��í�G� �&�ky����"O<TPE�ًe��D�"7wx"��4"OdAb��V�{P�r��[.
�2��"O���"s76��`&�!/��8�"O�4�Df��g|���ϕ35�jX�g"OF�@�+�:k����1��a8� h"O:lZD���e��p�b����M;�"O�3�Gϛ �Acο+�B��"O����� ���6�U,9���"O�-Ct"U6H�`� Pvm "O� ��� �E!]��mj����xhej�"Oj��@-������*�Q��1�q"O]�@cTΨ��t
wO !�%"OP 23&ɳ=%��Z�j�5����&"O A
�܁p10�gC�9/���U"O$9У�� ���b�2tlT""O����ꚋ{���!wU�Y���t"ON�kw�Řvi\�A�e�Rn��U"ONY�m�o�iEdЊ@@����"Ov�dA�,{�#˰4�D���"Oa�b�&,�<xۆKZ�j}Y"O��)�zh���'�-���"O
�`OM�>Q�m#0��`c� rg"O� �hN�&��y@�@����"O\���ծNP��Q�����HD"O�,k�h��X(�����5RPX��"O�lC�L��V�f���D��{P�QA"OhxctL�I����$�:?�	B�"O��ɅMG
pv� �&♋Y9��W"O��Rr�O�$��.D� �""O��S�"< h�C��?+<��"O��{�#�2��*��9m65�4"ODȰ	X$h� ���'ە��9�"O��)1�N�[s�m��G8V�:I�"O�TI��M�~G�a����8O�"e5"OThȖ��h�X]�S���K��]��"O$��� Z�	v� s@�L'h�8�jG"O�1����!6����	��B��"O�M�c
m�Ėu�$�X�"O^��BH� u,��k�G�ă�"O����a +Q��",M��Ae"O�%�1�ơyE�L8K�TR�"ODm���3J���U-��zIz��"O��c�L��N���L��81��÷"O�	0'H���~�"5l@�v)FQ{�"O���S��$t��F��6x�(�"O�\ԣ�_�(�Sʈ�y:�{�"O�p�I�3"�\�fc� s�XE��"O�2֪�=��p"�,�F�0��"O����W�~� x3�Ԁ
0$��"O�K���#^+���qD׾@�J,)"O8���)�-r��2�A\${���$-D����jE���`��	<�$qs�k*D��K��Θ8�(�!p� >��Ԉ��'D�4����
<��S�A�Tq�Q���%D���c��u-�9!%�٦;���@��"D��`�/E�mg�2��'#Vʲa!D��rw�E:6���ǮхX���to"D����?Q�N=���ϷY�0eۓ�5D��A2��?4��Z.Ы�G���!�$U*k��:���Rl\⒇��S�!�D�_�X��ڔpj�3�E��6�!�d�!xT�!�)ۼp�JE�w�J�a!�ա98�,y����`�Q��&�!�D�4p��Q�^u�i#Hޱx�!���R�0���:R4%bR�Q3�!򄂶@pĚ@a>HD�P禉��!��&=bX��` �5"�EzD��9H�!�Ĉ$@�\=��+�*T�QGMҞx�!���o����Ǩ�D��]j���
�!�DC�1i�� �ŀ���Q!�� 1�`�ƌ#����C�T�6Y!���0,"J	*ȑf���@}I!�Å|5:��D��O�]���^�!�� �!�F=�d����1�hl��"O����ȖqB�%�DgN�G�^��"O���L$#,���%� ���"O�	�j�Z'�pI��9wݮ�H�"O��K�)Vč�L�<��X[�"Ox���#əX�(h ��C�0Ә՛s"Ox<����i�lQ�S�A璍�"O6�Ie�2L�`)�@oȁ�`�1"OtԉW�G��i��Fv�q94"O�@�	$����Ċ1C�1"O@�p�䐖�f\�e�Ҷq/&Т�"O`�A��e:��d�$��Aa"O�)H�IF$$D�V�Ӌ��L*�"O^�Z��.9�����������V"O��*�U�U�&ӅO8�MX�"O�`��&_�pPM"��Y�����"OH��Ŏ9U�,p�-I��6���"OX��@ I��y*#A'�X�4"O i(0�۸D.�񰐪O�� @"OX�2��*넝J�N+`;�!��"O��Peܭu��J���8V`�"Ox@H&:�PYC��ԍI5`\��"O�,b�m��
<����%� ^0��V"O�Z`�Ä � ��G$��B�&�"OI+�-T�̱�s,�~�R�z�"O�,B����[��,V'OdBu"O������	Z(L��`�%[�p��"Oڄr�$5{���y��M��a��"O���c�-N�s���q8V��B"Ov4� �7Rv���
;�L��"O��qѣ�$z�9�®�)��D"O�1z��4~��31.^���"O�A0�k	R@�8ʲ��*�>�b�"O )p�ʎ�؅��I(a��h� "O:2ѥ�@�P�`���vC� V"O��sEN"?��q2�(QX@��"�"Of�Ja��%%�t��ٙ=@�y"O0��E���V	i��Y�zd�P�"O����b��U�`�R�M�q��[3"O>����5+*�#�N#x����"OJ��G G�]� �ʵ�E�H���"O��c��@�0C��0���"O~����=X ��@�ͭx�>�"O�,�N�)>{���B�hä�{�"O�y��aY�Ba���Z�	��C"O�5"g-b�*X�"�UQNy"O ��EUs�����,�
� �"OH\�	�>��p-Z)	}��I"O�)��ɇ#��H���Wt��#"O�LHf��A�&��3JBd9�ْF"O���"��2hr��Uh�"Mt�Z`"OJ�����	^��@�^) �l�"O&�ॅ�YPȘe&�4z)�Q�g"Ob����I�i-�������!�C�{�=Z�mT���C8 p!�D��67,��pE���b�����Py���?i����g� X4b���\��y���0V�RMK0�S�MZ�@ o��y�a���41�c�}�.$(P��yR�$��H�I;v<,<ɠ��y2�Z�'��q��-O̔i�P�ϋ�yҮ��H�c�k��x���Ҡ�y�n^�	x�E��c�,f,(�:�!U�y҃H( ⁻�,V6��xڲ�ҙ�y
� �=�kOG����F�}ENe�#"O�5�炟ui�lk��˱2*�`%"O���R��*�9�F��D0�=��"O�ꃪM%G��H�����9A"O�5 `�?R��]�@���
����"Ozk'`U�<N JQ	��"��"ON�B���ʷ!]��ܺ�"Or��ȝ4A���@a��L�x՛@"O����?g��)`D�ߋ̲��"O� �����T�R�`0 @�o����c"O����_�nٔI�ӬTj�P� �"O�р� 6�(���U��\�"Oj����
�kNu���:�����"Ol��%O�IJѱ��#��"Oڡ!E���-B�3�+!����r"O���`M�sb���g���1q��"OtPX&�F5Q�Ƚy�*�.i�,b�"O�U�LC�s�NԨ#j���N%��"O,Ad��b�$5��(~��y�"O���r-ΣI��Lcŧ�9H���f"O���#��&S�-8��R�x����g"Of���P�4V�0N����*O�K2Ȍ1�hH�Z7c�~8��'*�r���'���ؕ�P3�ҡ��'�8H���zRp%��t��'`*-��N
�	�x�����s&����'�5��ju~\�EΔ6���8�'��T��Ȍ0�ЊE�����'���adMQ�Oi��Dc��U�
�'?j0�4�v�8I)w��\����'�(�`vB֖��k�@�B���'>�(�7,�3�X�ՠ����D��'� �)�Ʉ�z�c��/R���0�'����Fg6�U�P�^W+P�h�'��j���	&0H�p�#҂_6Q�'�n1)�	��7>R�����]�2�a�'�f(X�+ƍEE��C�D2w����	�@ԝlM�5j� �+v�漅�(=Jp��k�5_�1�g�U�`��ȓQp~�X�g�T�E>N��ń�-�f�������ABD�|�ȓ�x]"��,��tY� �4��I��.�(T��8g���� �+BL��f����J�r�RE��G�S��ȓ�¬��A?LP4@Ao� "�Ƭ���<�{$�'�J9�M�3s�|��+��u3��!0���-658��ȓ(Z��Qe+�+ߴ���̥s�e�ȓB���p(S	l�����O��ȅȓ{�|�'GNI.^%j3��q�"D�ȓ���r�lPtA)��u����6��� 㐄u��(@� :��ȓp��!G�6T���բV�Ҙ�ȓ8�k��)b��
U%C0���ȓO�h��O�muf$[�T�K�Ɇ���(��
#p�2�z ��u��}�ȓ*s�5�4-�%w
u����x�y��9t<�RjӇ�����B�8kX�P�ȓ:V�m��OܛR��5��$N�
YV��ȓ4ml-� �60�*���F��0�D���Pޤ�1,F�n񌅠&ȍ+6=����>b�{��(ڠ�9��L�h��h��<� )����8݅�.�{Q"��PHRiR�e��8I��S�? ��d�J,�E�D�ӡ'�$YXT"O�C���r�,���&�d��}`"O8+�.�Et�9��l��m�"O����1vJ�2��Z�7�R��`"O��2��&��ri r>��"OL�R�*d�MRubZ��&"OF�h���7 ͐ԋ�E�
9kR"O��P���7Lö<C�!�S�hXR�"O�U��*��:��5�g�̷�`l!F"ObZ1DY�|�Q"E��r�B��`"OtJY��
C�Hg�e@�"O\�c�� �&�����ETF��"O�T�t��(	,ش��L�D*�9�"O�
G�O��0�ү�K&n�U"O|A�"?Q��RQ�V5��1"O
��P�N����YyT��w"O|A�
%���9�O)0�����B�O�~D�E���N�{��

7f(�	瓪ēb!�L��6gs�<@�
����ȓ3_̅�waR���)�JD:~f���.���ҟou�d9sOV�	�i�ȓ'��d� ��mT��Їb�><Մȓ�̱�a��L��iN���ȓi;�d;��)^u��ê(�����1x��`�<U+�hw(��y�d`��E[|}�p��F�,��)ŤJu���ȓ?�q�f�2=��ccK�$�D�ȓF���B��I�ڭ+�[=�N�ȓb�h$�����@0.i���5a^���b!�j��*U
�µJ�4
�:�ȓy)f}q�Zs�VIq���x|8�ȓ%O��z�ˋh'P�X@hIn�J��HY��ȢA�s��Bt%�/8��ȓ׼�@0�j���W�t��0��&b�`��6�tA�G�-i'&!�ȓ%��Q���:<>�x0eۓ.�t��ȓP���O�b�I!�]����ȓV��k�O�f���b�_�l�&��ȓX J���]�v����,U&ê���h#٩@�Ri�xB��1�p�ȓ�t����_^Z���,�M�б�ȓd�Rx "��,S��b�m�B
p��e�>�iQe	QD�Y�3��θ��GN�C��gS��j���&
8��ȓd\���aG_�e��Iw�X�(|z���b�b�pAݺ<$�	
J
]�j�ȓD1dp'�D�I�0��.� ��نȓ5v�9`���_�n\��cӅ3�^��XeV@�̉�~.�2�^N3����PL:�S�
=7�� 
öesF]�ȓ���3�مC��u��E�q�\݄�OC��B��فSڍP��lx`���4�Ơ#���	 H����ǝ
P؇ȓ�$y�f(ȫT�a���3i<ԇ��TEZd�Js_hh�����+�j`�ȓ1[�`9�#�rZ$s%'N�غ�ȓ'�
�*���(��*���!DȆȓZ]�H�u�O�| a�E���N�z�:!�(�T�1)Auv.0n�P(<1���>�"�(���$e��A���\�<9%�.l=�Ղ��J�;��(! �U�<@Ɛ�0��푁���3�P���Pi�<����#�q��԰P��8wK�^�<�soY�x{n�
�
4��� )B�<� ܬ)�AM�98m��+Iv�"O��*'�Q�ͨ�c���eӖYi�"OP�R�lG8����br�.��A"O� Kg��;�Б�!#�28*����"OHU��父W��ڃ��3mv�C�"O"�j�*���
�2�m%K�l�"O��Ye�(̈́�PG��&�e�`"OHq;���<�ܕ�熋KhB��"O^� �J��x�A�Ne[�a �"O����n_�G���P�O\�#A�E��"Ov)�(�b"���.3�5��"O�<9`�P3s:v{GN(|��� "O(�H�!��K� ��W�N�~���`D"O�tIbD��hx\�Y!�Fi#��cQ"O�h���)D��A��[#q��"O\��*K/�j��daCr����i���[�R�d�ҥ�=���f$�=�!��E:<�q��8�NA���Q�F{!�Ҙo[�*��O�����o��5�!�$ nl����Gr�Xz��q�!�& �x�Z�%��uю��v�KQ�!���(a��uCQ��Ȩ}bЌ�bt!��sVIaT�˜9�(t�f��Oc!�%���%<s�X����bH!����6���L^�����a�!�*ax��B�T&1[�y�©��*�!�d �96R,2C�4_FJ�Hׇ9�!��W�1Ƙacr�Ǆ9�M	�Fg!���Q�,��t��8MJ��F��60!�Ė�T���q���i�D���!�dR��
�"Eo���ص�
2�!�<i=z�Z�)$@x����[�T�!�$���A��i�uU��XW��:�!�$Z�O5�|җ��pp�UP�j\b�!��6��[��R�`✺S�8z�!��@|�Xe)��S�}�bƟc�!�C�% �i� �F�o�2�@C2�!�DQ7	BX����=��Y"0�?q!���e<ib�B��Ei�?!�ͺ��c#����s���dr!�d͇t`�]�����tP���J\!�B!D��Q�c��=>��Y!���q%:��!��'�8�`s�͋^!�D�Z� ���t�"�m�T,!�d���ptf����E�Ѧ�#>!�D�%IU�p����b�����㓿4�!�Dڬl�<���K���PrC:�!�$R�<ޞ%�4��9�RHrMF�n�!�$�D������Vh�] ӡ�5r!�d�&fcl�QL��Cbx���t�!�D5sj:%Ȳc�4���� �2o�!�$�9�Qit�E�4xF�Î�	o�!�D
�Otv�9`��aN�Dx���!��׿mx�� ��{����ˈ�P�!��4^�Bq�)*����F�Zx!��������˜3�T�!@��5@!򤄆B��D�#i�z�b��$�Ug6!���Mƚ���	P��-����n!��R/sF.�2��N�h�b԰�M�>4!�D�<%�(����C�8�q�a!�D��
1����@u��V!�䐍||H�hHKivh�(#�Ζz!�W)/�n�j�G�p�{e�B�d�!�D�8Z}�&&�%\PН�T�!�� 2x��A�65Ġ�wA��<��"O��R���N�|Mk��1n�Jh[�"O,L5S��h��ӃO�L�H�S"O��c�oČ�^�9va�.~��1"Oh\�@dL =�|%+�K�	���"OH�1,�&[�&���H��b�i!"O�-����0�9?oz��-	$[�!�d�3�)��Щ&aU8�kK$p!�DX=pRf���P�4�PMD�FE�!�dH9là�z�N-k�fts��ĉ2�!�KX��'ںw��<٧�.o�!��5�$�Kr��r�(�$!/>a!�ɩC�V���j��B)̱$H!�E.H�.��$�ץs���"g��:!�ċ�(�u��.��x�l("�ոJ�!�$��8v��x��>�b�q�J�*�!��
�y^�|!m��a,�*˔.�!�C�hAjA�ZyF��)���=Fq!��͔L*8AV
C���$�����6�!��4B
X���/ts 혲i.!���� #3g�f��LL�{:!�֩D(0�`��A�^����%QY4!�҈A�LR��Oܚ���=t?!�Dܛ:5<��tk�"|������	B!�͘%|d�0'щ"A�U��MQ!��#.Ɋ��"�H u��4�()���hT�eoм|��}:B����i��S��9C7kЍC�RL�C	r0���&��|���$`�����ڕ�ȓ������(#�cU��U��D�ȓ8t�yh�B�fH�p��s*�ȓ0	�hq"�F���ض�DCL`���(�G��6Eh�KLrl]�ȓ�px�.H�x�+r��c����G����}h􈓶�B�/��ȓ!��K����=sB@G\?.ZxQ��a8������vɹ������,�ȓ��ЛCg=��BN�:4L��F������Ut����Y�HW� ��T%,��τ�V�Z����2&f`���K쪼2ū=K).Pѡe�!� =ΓS��أ���X�(
�U��A6`���N��AP&{@��퉉=�> �4Ϩ2�0�*@�q,��$\�XH3B�8� B�	8��hF�`
��(b�ʇ.\$�!A���/��������~�`�ۧ,�a[�j�;%SȘ@Q\B�<a��H�9d٫�#ݶHtz������W�������|~'�����	1�2|���p��	T#9��C�	�0��ŉ��6��j�+
�~�@`Z��[C�1�Oa�6
�2`��e�,er (1��'e(��?����w����ɒ'"�^q��@�<ASd��S���0Ƨ��۲KIJ�D��N��?u83�,#b�5�T��f��Upm1D�lZl�50<NHI%�>^й�@,��.�����A~�@eF��@�R��ҤDe�!�$W@}nx!���+�b�֧O�$%2X�tm&4�Ă��)���&k��w��*O�@y�G'�ɯa)MqգH�ϴ�K��2�B�	��DP�F�{ʂ}���J�o����ӎ��I�s%RYQvl��O�8x�덢���r��H��\jsǇ.$�Phi��.����!��.����?2
,�fM;�HL`�&�3�'w�zb���H�{�%Bc4���)\L�p�'9��H�b�B������oN��wd��ax2�]�M �O�Q�Ծ~��y!I�E�G"O� \uRTfO�^�z%���,3�
��Ց��Rf��w�S�Og��� ƣ��� Ō��|���J�'1�ɡ�AN�M�ܸ���"'�$}:�y����%��yR%��jFxK��͢7��A�H�6�xrE�>h��Pdď�V����n�04(lUO�HJ�%�dǀ8�b
�gR�԰��'�V5V���8���PP�A8ȹ���/�!�DT�{'��B�CP�fr��� �&�F˓A�q���������85n�Vi���=8:az"���$��)2�Ӊ��{NXz.1O��cW�8<OPYkR�@C2Y�H�d�Y�e�$(�S����C?�<*#��'�<틐#��6��(3�O\�ЉS�(M�/K�r�j|r1�	M~Bj����'�v@���r2wg�	
�'��Q3O�)]�"�*QA�;�d��V��@2u�"�S��92NؔKX��n� Ԃ������ȓ6�$;�g3,���0.V�>�'�DKX�(��gM3@�2���5����e�.4���я�eh�QQ�i�� �:6kM���B�	����𪊎P�>�J¯^�S����dǨ_x5%���GR�c��	"Rb^������+D�p�;mT$2��W��� 5�ɫ\��U��J|�W(�.:��u`����4ӎap�P`�b�P:�J|Eh �$Ta�),JZ�5�҉P��QJ>��I�O��D	a'���f�ϧ�X�&)���8V��B�(��I[�XPc^|Qz���N�-��	4�M��:9��)�����pbe�L2�ի��M'�ԅ���9p�\A2R��:f��ɚ�& ��هDitY��O^�[c��)0܆89���$��T�f"Or���ƈ4s���	Rᙓ0�رr���f�L��'D*�0W,ˆ1�A����1&�ą�	�E.����7t�Q"�fL1�DX��o�b�aSg_e�$�#&�2��$���܂0��C**=)v��!M5Q�8	�H�	�D"��R�c�N�O|h�˂�]�e�H�c_&\���ܴuZ��9j��м��)ps�?��}̓?;�s0��5Ә�ۓ�\8h�~B�.R�wje�qaO�F�@{�͝u�<y�.�Q�@�T��O��Lcrf��%��$�O�.KZ��T銵$b<̖O��4�4.��ʦPI�i._�$ɲ7� �OA�U�� $���S/	8:��C�%�a*^�	b�83󎉨�c�8fY�H�;H�}r�	#��L��N\�NNtGyҠķ:L�iZ�a����T����LH|����xG� �����ɉB3\Y�U"O20���3?oN��4h�r>����� b:�,ۓ&�N��},cv��p���0u���}λ5d(9��5[�L�YViÄ4٘i�ȓ�;�FޚKb+w����dq��1@k���Ć0q�X(@O�|2�&ޛNn�0��#�6`l�ś ' :��I��9|O ����@�w��܂7Yz���%G�9C�C0`�z]�%��{@�a"�ߙ2f>��d�������^�:���/Z/��O�M���/���u��]Z9[`�0���L�H��P-Wԥ�K׆#�|C�ɤ!�Q���ZP����kN�8~lEP„o������*)����s�%'�I��(��vޭ�G�,��X�OY��l���8D�X�4-�c8�A�)L����V7I���C���o&��t�irr�iξg2�*�&"�	�k2H�R�L@+��8�k�0�2���N3r��19�	�9n>P���e��V��A㌹F9� ��S�	S�i"���82K��9LOI���%)�(�'��3�8����EE�0
N��gG�����.�)@$�/���K���X	ޙ�1�$e�Dd�ʉ��y��՞#䬄{4mY��t����
�V�	2.J:Cـղ@�֪�hHq��#E\c�ȼ���C�Ocv\�ֈЂb��y�X�<�7(��
���dm:�aҎ�x�f4�@��M�P����!�$�����mUx�L���ԠJ�G@h=y��nh���I&����I��h%�Y����']����¬�/P]x������OM�`��hJ���b�\�&�L�poQ?d`X��)3�	�j�0q:��I�1Z��a�!{��,��K�B\��cw%ĊY�� Z@NC�S7�q��c�<I��J%A��㥈U3/v�ի��Y�U��@"$�Y�Z�L��'���q�h
$C��'?��;"~J-�r	���,מ�T��m;�"O� ����m�+"N��%�37����Jޚ�L�"��BW�#Cʞ2���-Ŀ)'D�0d��)F��� DgL�\I��L���{�$OE��\�A-O蘉ыY�11��0��G�;��נ���%XcCZ�A;|��s�'i�a�.��@��,=��P��$� N��aC�/T��Y����Z|�h�D��5��}k�"�c�𤹖��Bڲ��"On�Y�J�hw�� G��#y��-+�F�t�l����s��$�g��!�d�y�
V���yר�#�Vi��'I(8�h��D�Z>�y2��y��P{�	��D��L���Se�űJH�w�j9b�kIRj�|�OF���D�d�1�|�yS�<Ȣ]��(Ǉ+�a}"��S��)g���{�z8 P��( ��U��̀Iy*�jǂ ���JU���2�K�2!�ѵ��9ǒ�K��,�3��JC!L	~D~yH���0%�<0�Om�	��� k��U���@�V�L��'j��HՄ��
�[g�)Ilx=@�'L,�ِ��gu�����Eh��D��H7v-�lY ��XX��[�y�[�x�Hة�bV�{� iŨ�u#�=�W��OdQ�H�W��tHO?� �E�Mt�� s.�ZZp�s��<�O��e�Dن5�����I�5��(3�x[�-ؓol���� �`y��L��W�I*���!�ةCz�к�"D�e�D�����9�!��7�h̡���D��1��A�2}!�߂�|��c̟>Q6�������'4P�����S�N�(�$��m�ܨ�	�':RQ�f�6a&�z��7([�Q��'��� ��g\@-sV"Չ^e���
�'�� ��3BT�q�ȁ�}��@�
�'�����w�.pf@�%ftQR
�'O�9H��zD���M��� �
�']v@�������9���$�nT+	�'�X<HJR�=|(IsO\>a��P	ӓ��'�����C�/&u�BG�=}��dX�'T�xQ������h��D2,��'R��@����}Q�ٍH�<i��'��$���\��<*���>6ؘ��'U�� C�Q��8���P�0��k�'b�	��^N�H�Р�Xc����'U0Tj�m1��� ƃV� ]!�'��p�����':ف�c�@4��'�́'O�Nظ:dڋ�>�X�'F�ҥ�G /*y�/�$�R�'8�p�&C�n ��QF�1����'~쩋2 "3���F�2=�	�'� � 5拈E`Љ���1�����'E�0/�$d]Yz1#ؿ(P!H�'�V���!2�|Iǡ��&<z�'�H�"���jM&��掖<F,i �'�^���سN���y^Y>�H��!D�(��(X���[Fi
-!���YM0D�`��ΤS���Z!q`�qg..?!
�M��p���D	Y���	`�oa�)��qa�����R�D��[x9�C�)D��ri��¨IR�U�\c��g+D���D�ʕP4i�5i�}Ұ#�;D��Y�f�i���(v��+����*O\<���1X�lK�B�k�<�[�'-����P)���p�(I�HBґC�'���X��j-�M
!®D�I��'[N�P���_=�MZD힎� �h�'b �ϟ�� �����'*F���Q�n�� 0 յx���H�'�B��S*�PS�}�'OĪ�Y��':�����.%~*h�V&DTT�p��'[ Y�F]ipp!A6cH�V���X�'����5�_8:a�e�D,[��	k�<��"ž) ��k �>�8=c��\�<� Q*�۬y���F �><B�� �"O�i��̓!+\���M~�@<Z`"O$Ii�H��Z�c�fZ�|���b�"Ov����)V${��'2�2��"O��P�*��fl����T�޽�u"OH)0�&���b �Y>\h��"O�0ЕC%OZX)Z��̚J#*`�"O���ώD��,S�J� ��"O�t�T�OG�8;c.^v, �U"OZEH�!賒�Z]��h�"O0:@�SC
��f�=5�x��"OH����k���!\�,j�"ODM9�ğ|��e�O�9�~4[	�'�Ġ#��Qt@b���@`�'d���,	)(b^��c��/Gݒ�c�'���� �=��x�.0��m��'�� ���:7���qd�/�J��'�(��?�#6���#ѶQ�
�'�R� �.�B�0�@1��ny�)K�' ��jD�ԅ����0B��S]��'j�yx����2WPd J�'-2(��' |<�u#��.<���N?D�b��'�@	��K�_-����l��E!����'N,�
��j.�P��>3TJ�'DQz0��}40��S�x`���'�
��CC�(���b
3B�tq��'�n!� �/z1��a�\�>��T�
�'W����@V�[vz=�aF�-���8�'9<E�Y>yFqP$��H�.C
�'����'p9���R���G����	�'��m9�`ph��	¢��mQZ�X�'��(�'�i�`=1��W5q�R�Y�'�.4�/Ʋ9�����6h@�R�'��ػs�ӂe��]��I��e�����'�(0P� �_B�Œpȉ�^HT1�'m��
���
��@�ŉS�I��(�
�' h��<�B��d�*61��	�'��Y����72X���Hɦ!j"���'�0�c
ѯct@��pu��yb]�@<`1�ąJV&��#(�y�h���`\����һbL+�'p���L�/K|rԫTT=��Yz�'K�d�4�I,4m�cۗ,���
�'��m��ܿ.P��2C�/8����'�T���@�Q�Dt2�]&����'6��� �܁exZZ��9.(� �'��e"Q&K�
D�!n�J�P`�'��p�O�;��x!f�%:��=��'w�'�Ia���bC�%N?�"�'~��n*`!�����Ȫ]�
�'��@㦙,-�b�h�N�YN}
�'2��v���N��W回P�"u��'�R�q���w��VI�
0��c�'�ƌh��$1�=
��Ʉ0��)�
�'����&.U�Hx���ϱTE�
�'��YS�L!az���,ɤ`�	�'t�= �m"!P` ��%~T�	�'&�!W�	V��Y(�,�a�ʠ�	�'�N�;��-c6� i�Z����'lZPc��]}�P\E�ѷ ����'˪a���_$���+	�mX��'�ޅ��Q�D/~�37䕌$��\[�'"�,�U$�B���I�`#�Ry�'��������<+vm���[�/���� 
@�A��J�-I��US� ;a"Oj�#�K�j�e�J���"O���ˁ-N�Ճ �S!$���c"Oh�+4�)C fTZVe�< ]��c�"O�!r�QF~5����!V ��"Ox��b�I.X�2f�.0j�"Op�"�b>_j���Z�Y�"O<��$У Rf�QU���33�P3 "O�,��L؀yd�h�F� .��Hw"O��a�lK�k������y(�+�"O��AR�P�A��HGG��rJ�"Oj�g�T�nd�j6c»-"�h��"O��p` #~U��HT�i���	�"O�!"���*E��7f �c"OI��j�5��$�f% 'v����"O���%"�F��e�`$L�E��`@ "O.�R�+�F.R���A�I��M�d"O4��f�a�d�T ���vicP"Of9����cn�{��׵�9�"OB�T���T��a��P�5"OV� �.F�R/8�s�D�%��"O� h�lT�b�)�
�VI��+�"O�:b �UF���0D^�8yQ�"O�}�t+Y�b���BSCW<>(��q"O\h�۠E*vīV�9wB�
�"OBL� �Ğ8�Y#Q&�$o<!�"O��A���&�m�#DC�$��R�"O.ȒA#�Ă��2�Y���s"O�]Q2Ğ>&T�`A��3jW6�� "O��B#ؙaip� &��OZ(�I�"O�<r�i׳)�BѠ�&
w��C�"O����$y�,��Q�S�cVX�"O��
��	&L �ֆ����}@B"O�Ћ�)N�4��ED]�DɖT��"O�Uȗ.�"_������<���A�"Ov��3�U�4y5�n�,�)�"OR0�����Z���G	8qz�I1Q"O251�JA>krx�z�/j&d��"O�s� v�T�	��/5�"6"O�M���4��ag��T,B<�u"O�m�t�īEA<<2!�5t04i��"O���C��ބ #�V� �%kf"OZp�B�F`"\�P������C"OL���0�m��CHXh$"O��?�U�扽B[��"O�u�፞�u����F\�mN�ղ�"O��hqꞷ:�H]"�Ć3�{V"O.����ӟU*�|qV��!8��R%"O����}N���Wg�7<a��"O��@�	_{�����'ͳ6+T�"O̱��Z�B�T��	X�Xt�""O�q���<Zg��2PG�.e?���"O�����C/d�x*��2�N��2"Ov��*@�]kz��'A�9�)�"O
8�e�?
$��8"��i[V�[�"O^ĉ$f\*[��QC@�_L� ٰ"O�MGFE�0�����Jصl�m�g"O� q�'��%�$%��$��ex&\s�<���;VW�`x�
U �̙�@Ci�<1&JE\����E�99츴��`�<EG�hm�`�sn�-Z�Ќ���^b�<��U0d�� +)T�-{#'�_�<���w�0\ǈ��V�����Rp�<g�<Α�2��! �$n�<� qQ��,U��
#.�(*��ѐ"O��10�
�7Ў�x�,Ĵ���Jc"O u�����w�eaGʈ�'���"Of�Q EP$��A���m*Δh�"OY��N��1\���Q.��n|�ۖ"O��ӬW7���M/itY�1"O�!1��=)G�����^�$"OnՉ�BR�E�F����<K��T�0"O(�q��}V.�AÜ}�h��"O�� �α&ரiS�%��"O�i�+�U��Rf�̏z�d��"OP*��ÿl��\�w�ύl����'"O:!�d.� �xRAA0[�4p�"OL�AZ6�5�� P�f���"O�d�톥
hTP!N:[�B"O�9��D�� iem� \���"O|�3�,� ���P4�Ы1s:x��"O\Q@4F�M�:�ڐ�ƞUmG"O�l{��/]��4(�X�}�ʩ��"O�����?8К-S ό;'|���"OR��e��0Z�hs�M0I�$ s"O�b7K�?@)�
�m���Sq"O�lG�=��}���5�4у�"O*h�2n��#�|��
L�nۨ�1�"OT��'+	#"`
5i	6���W"O�l��΍��QqW�6XҘ���"O� 0`z�{�#Z_Ԗ���"OH)y!ކ�·����`��"O�{�"�a�*=���m���"O:�B�Q�&�d�bŅ�"`�:p��"O�m1��ѰS�����Y,h�Tx�3"O*�I&!��t�^B�ӥa���y�
�>�L�+����\��E�e��yb�58��q3��.x�L:f�Y�y�J�!���BĎخ�&�2U����y2b�6"�:	�5dЇ>n���,�y��W�f��I�!��,`4`���y�l�4�%�#Y�LԐ�`Ɉ�y�	,\�^IA��W� �h�Q%�yB�/vH�P�F��<�0��K��y���mN�q�.[�/[L0���ۡ�yR�\dRE	���.}̐y�*���y���R���G�ӈ:>���y/HfO�arC��=H
=�Bd�3�y��ӵ���y�I�GQ�-���I/�yS�d�|�S�@�nI�%HJ��yR#��l*F&�,���"��A9�yR�A�T~( a+L�!@ A
5N-�y,&H�eI�ɐ<W�!�WG ��y�֫u8P!����T��)�[��yb�W/ea����۴6	~��c���y��h�!X�{�����+Ӂ7�j�(�'����%��emԉ�BKԵ(�f9�
�'L�tc�bL���I�Qʓ�#���	�'������`����a�8	v��'ѱR#A u4�0d���e�0��'RvE!�
4|Q�l)�%�Y��'�hR���3�h�2� ]sflz�'�Z���U(#@��2C��-b�����'���0B��Gll}ȁ��-'�l��'���5D�� 9�,#!)/��Z�'��@K���
$��l; �R"k$��'ɖua���)G4����ı
�'<�$���bR08r��91��y
��� r�yU$O���ے�r�Y�"Of��Q�G8�̨T�C�L�hȷ"O��+��1	曁��:g"�@�U�4D�h၄!q�@����
�	�p�9D1D�������ʬ����R@�1F#/D��jp,V�O(Qar�̽\�"�R .D�$Zq���jZ�����K�8*:D��h+D�x`[7!:]9u&�DJ�ՠF�+D��PbH�P�!���G�+�r��2&;D��[pϙT��4A��D>��o6D��pլ�,y��Ã$=���P D��z�"ѸP�آ��ߢ2PHq >D��Ο�−�O�5&�L3�j>D�q��5R�*���H�Sr̀�6D�P�A�K�o�,�ۇ�8{�ް��j4D�d���?o��yӥ)A��k�n0D�\����,8�.� ��ӊ,�x�ca�*D����':�u����9-��]���(D�a��C�|AN�IC�OaGڠ��:D�p�n��W�zefҢ����<D��a'dH�Z���� �FM�T�;D���h��`
~����S<�F�`��7D��0�"J*-��ti��D�@�6��2D�$2rK�(��4��^�u�C�0D�,���3r�@�p"C�&����.D�T�'̴d���:C����2qڳ�7LOb�)�@�{�:���'<`Ҝ҇��*W(�P#���'��zQ��}��F�J�k�Q����R.�"}�'����g̚�T�԰�g��.�`d �O �q�l�S�O��P�MC��薜!�����'n@����L���؀��Y�lH%oB�<l�y�4+����v�Q�K�4r��S���e��d�N�^����)6BN��q&�&<��Y)P�qO�(�*�)��O��� �B�Z�K4�Ԗe��;��1!���.�Zw`�J�'m�d�*�B+�~�`@U��O�>Ƀ���B�ƅ8#X�J��Dzc���Xa8}!���	�1�fY:2j�K��Pa��Q�/�5�?��Ez݉�O,��|��P	���: R�:�H�H`O����i�����T%d ��l4�g}2"��"�����7�
d���-��Isn��?�J�-~1��c4*U�.(�˒i?�a^#���h��$;@�H�q8�r�G2H|�e{��
2��0�?E����.o��{ģ��4\f�Y�m��:�yr=O�a�.��`�Od�Y����LQTذ�B�	]��pС�Tu?�ҦM�<15�Î�~��SL$1q�̚��"��eB<@dd���dR�<aA���~2�SYy�d׃sd��� A�6��x�l\]�r9lZ�^B$�'��7��?=Yu�W�G�t�V�Jw^�� ��U�zQp�O��	�A�a���3��<P�.������/�)~ɼb����ɩ����'7�@ڷ$�))�����4��O��+&�ivn���e�O���>^r̤���B�a�v	)H�G���.�G�*��5�,�>�G,�tC�����(������\P�<���H�F�J-S��#{'��s�
L�<��)ۇ-�t�x���p�eKSJ�<)C�E)o�(W��1G�%�d��I�<���ΌK^^��+���hI�<Q2응#��P�f��Q�2)��Lz�<A�b��$��Cw��vZ\�
T"�A�<���'���1�#�;��2��}�<��a�3w/n����G�:�Bm
2"|�<!a V�	�,����I�F@f�-�y�<q�A#n_�鑥�C�.�YKs��t�<���:�Fd��`ٴ
4��E%p�<)�� fߖ����	�*5)�E�<i%�~LIW��(2�rF^\�<�#�]�8!�ُ%�"�'"�W�<9�2}�Ȱc��K��|��k
P�<� �L�wƒ;G���Ѣ��6�J��f"O���� ;���Y�≁;g.��u"O�E�Z	��y���/�ZMq��]D�<)�j��5.�	�5��)��%9F�@�<9�H�^M���͊�Ke̘�3n�|�<Ys�?����䍏�*�V��*\A�<�'&�ⱊ�;_�䙘���}�<i'G�Rqn�äG��e� ���R�<��hT�6��y!Z�EO�����i�<����햌Q���}�V,���~�<9�'^/JIF �CD��"��Q�O_�<�tɗ�K��i
$O�M]��� b�U�<aC�-C�\в1/��,��g��G�<�ҤҪm����Q�܄��@�+�B�<Ʉ��6�p�i���(oŖP�R���<�.�9�>�Մ^�~�6�QS
G�<	#kX�}	�E��k�Dd��C�<iD��T�2ԁ��Xݠԋ�kLJ�< .H0�>Q%-��y+j��W�QC�<AE�̕5�����!����{%!Df�<�f�NI��U!�:��%�f��b�<12�&T�6)��ჹB(�3��EF�<�s'A�y�ЫT��8I��U��C�<Y��A�U0��K	,<�lăr��@�<a�%2��+bh';��$a �s�<�3Y�c!x�sN�&Y��y��Ps�<���
��%lU;��5)F�r�<a�ĝ*Ō�$+E��@X:WA�D�<�֡X�F�TP$Kv4X� D������*ո0i��g� %2�`9D��@�K>�b�zƇ�F�Ĭ���8D�H�SlF���ljƈDϬܩ�E$D�����ȃd�Xi���´/c��pui!D��ې.��I�̙��B���-� �#D�P*�j:^q`��7LƫKWNiid�"D����jŖ9'��`��=?���@ j D�<���Vkx0{2F\�u�8)�g D����I(٢��NW	��Ts��?D�DA�M=���ĭ��U[��(6�<D����bhS\98�`ӱ*�j�y�(D���Q���f�t��LҜ
���0�E4D��c3�Hz���Q��_�6|�T=D� �&BW���)2��p"4�à=D���F�Ը8����3!�$}&��G�(D�l	��UQ�6�p`œk��9"@(D���g(��i�����&����%D��C�*J	Eq���P'ѨČ��(D���v$P9�`A�O�I�"��j<D�|S���Zǩ�{"�գç9D�L�v��lg���m�7��9�a6D���V���h������HR�t��e6T��j��	� F�'��X9t{�"O  ���t�8���mV�i.2�RQ"O�a�S.�S��\����!�|`�"Oz�d$Sh�ԠE�&��h�6"O���$�r��6#ޗ}�\S�=D�"�ElJ��\�݌�Cv":D���e�D�H9��p2�KR�ܑE�9D��� � ���pi�;���P��%D���k�6�
}� ���@1�D"D��s���:*\�� (��U�т?D����X?`w\�j���7K�`!�`� D���������=14�S�#�>Ţuk>D�\���,C�8�C�O�J�{4F:D�� nѹ%	5^�Y+��G,1�⁂�"O>葰B(m�PH�Pgl��ؑ"Or[�呒$Ez��֏sH�1�"O�i�ɄM�!@�mF�W��`�"O�� �'�j&�CmJخ��P"O\h��'ʱ'�jel{�� K"O,LA��ۡ6���"cȚN��� �jd�J�(q�i�%蟙,)4m����=�4h@m�1B�OK���@���,�����Y�L��B�jV��ȓ\�*�AϞ�J�"�ȓ�'����A'*���g�	$�"R2(	lÞ�ȓ%f�#�f�C��p �"�+
���ȓ2Zi	��]�n�d�� &1|�P�ȓr�T�A��=/x�S�m��Z�ȓh=�-���:&���������e�ȓz�����C8.O(p+WgHP�fԄȓO�ȑ�ӎؠl��jQ+�Toޑ�ȓe� )"��I{��R%�4�tT�ȓ{���FC�������s>����]���
��1�ǒ{P��8:س�ٻPyf�Y!��}0̄ȓa�|�� ��`��'L��$|�ȓg��5XՃP�V����3(�@|���Iʠ����$V��@�dD�v�M�=y�������z�&d墒� شTS��Ρ�y�(M�?���Ñ��b�~�Ç����y�� k�<-���V ��c�H��yܖar� ��Q�HȀkvɄ��y����0]� ��9�`<����y��̻L����9�1�p��~�<��B
z���A�@�<rd9�`&AW�<ɷ�R-3�B,��ȑ�LyB�cB�Q�<ip�έZ|bd� 1�,0#(�Y�<ϓ�:�XÅF�c2_�<)[�w��u�r�ј*�Qct�@�<iQ���l��
��܌�U��W�<� �ߺv�X[�CJ	 zZ���n�<���8W������_F�#g)5D���h�0l��c�����p�1D���ƈ��U��z/R�rAL�Ь0D�<���8s\�z2�;-�$�*OD`�&��e�>q��I��A�����"O�}@�׶�F�ĭ�)e�Qk$"O�T;w�S�>����Ԅq\(js"O�P;�Vi�JDɠl�&d lD06"O`5��J2���+�
-�1�5"O���s*�"M�F�D�)[�zL�b"O�)�pj�pؐ��&._&+� ���"On�Z!������4�Ww�:=#�"O�H@�Ȇ�3)H�DӰ~�~\�6"O�=
&I��?k6� ���"Fn6u��"OR8��BW�}�z��@mٹk��y�"O�m�C݅'�pi���K,IaJ��G"O���BĮu�@�A�P�f�]�3"Ob2�S7,@��Y��� ��a��"O ��!��"�FeQ	�<O�T�f"O�ig��]@4�y�Hǟ`���&"Oj���N]n��j�h�� ��Q"O�iT���(��!A8��*�"O���囐7�z@�a~����b"O Q����^٩��5�8�	�"Or:@Eb��$��C¶[x�$�G"O�˅��	���3� � pRЂr"O� >My2E]d"L�����C���"O�̛�F8_��ia�%a%��"O~I�5/E�z���OU�wp���"O��l�!>�App�H�va��/"D�tcF�֞(�M!�a�D0ir�
?D��)&� ^КL�m�����3a<D�H�$iB� ��8`F��J���2��=D�|:�d�Z0�с�B�0C�X!$�<D�`	�c�?����򄋖_�h�%`<D��B���+�f�J�J�0ɤȊ��:D�����}ք��kH�e��=Yq)%D�T�+'B��p"�@�+h� �h�!/D��AՋ%i�Ԅr�T�V�<etI+D�����\p�fh��HE[ת*D�<���Q:�d�Q�	�����)D�\��J=p���%'�e��#D������U�*�i �%~�0����>D�L�u�ŊT���!c��
pa>D�x9VDF�j}I�!�A�O��U9�l/D�h��&G�d��%a��E,D�D�mއ{�X�cfk�y��!�)D���r����ҔK��v��.1F!���g��mk���� �\����G�o!�]=�T �bLQ���R�ՑL!� ��1��	-~��u4G� h!�D�*�iJ�l4x�hH��EԪ!��cҼ�2%�
v�����2�!�䒬d��a���xlj�Rb*Za�!�$�	h�}���X�8}���q�!���sz�����e���W/ 5�!�Ec��=��:h��m�*�!���V�Y"�&ݽD$���2�!򤅭)��HZJ���N&P��hc�'"� E,@y0`��4�̞^��'��X(�
�VQ[��L`���2�'�܁��� aԒuZT�DX5X���'0�˂�Q4���to�x#`%h�'�B�3j�.^�v)B�
�i��%R�'�x	U݊���1�62�@�'�`D��M�%�a�������'�
���L�\)��"UAR
Tp�'�n�Х+@���垺@ɰ�h�'-P��c�����7�X���' �����3:@�s��n#�'�.�y���2�\5�Q�F��h�'Y�d+��FvD0aI^�p�l$��'�8=(�.��q�2���ES���'i��xT'�'S,�;���F88a��'jRy�r#���v�0��q�5I�'�h�`���8=>�g�H��
�'?����!�>8p��`��rH	�'��!+����z]��xd��#l�|I�'�Ha��I�1�t����ee�8��'��a� 
�.��)d;^��'�,8@  ��   >   Ĵ���	��Z��w�D�8,���C���NNT�D��e�2Tx��ƕ	#��4"�V����cV�m��^�9z�Э~�vu�֌Zr�p�RE[
#E*P��M[��AX�nE��$- RO�Y�b���ן���&�9@*�{��JU.I;l��$�Q�p�Ӊ^-{���K��g���e��	����3NX���H�o>���d�=O�I�nI�|IĪ�ʓ��x��9���'p���S��b������6��	�q'�);�fט���	%��'������`De��v����Y�r�$����dh��>�f�
z
�x�H<�uG��$-�Ocr��0m��pV|(*�`��|��'�@( �$�H�>�'�N�*%��B��'������
`�^ ��B	C�b=�S���82�%�U�'+��?K|$R�_5�"�9"�$W4�2�E�CYԹjI���%�̛VԀ�kM��$�t�g���y����rZ0TĨ�l��׌�?�R�Q�g��5'��i��P�o�ړO�h@�U*V�9e�P*e�D�yPW�d�`Ջe5}�U��P�B�'(�	<5̩�)֪F�
���8>��ԺR��>a�����^��B�`P8>��a���i`	E6{`�}�O����㏓�E�r�$�^*�(El��N�6�P�)U�@dН'���H��E����?���M�X$(��X)=dj@����
��ʖ�S=�]�'쨱��D�J�'���y�OY��y2��"��lJ�	��ԋB#���N�I ��Ж�|b⍛!��N>i���.�~��w�R�Y?�Rd!�(�d�p�$��U�oAf\b�|OPU�F\��8�2��4f��}�,Eڄg��C�&L�DA4Fv $��	Ґ)#����+�A�dF �8�c4g��?��_TOt�a��A>sH\���Pym�	��U�M>�A���0��!%��ڠ(:jf@�']1 wȄ)��D �	"��7��r��I�f��Īb�ށK���(�0u��gـl�lq�`!D�l{��   �D�x�	�XLv	P���k��(�7*�?*
���ğ�J"��џ���� ��"��4Mv�Iu��%�M3�w���֍Ϙc+�	�b�w��`ÓE�Z0���"db)�/O�|���ˠ&H�|`GDи.x�}���'[5�(O�p�'� Q���ц9�@�;�l�y��?������?Q�����O��0W*����E��섂���`R��O\     :  �#  �.  �9  �D  �N  �Y  �c  2j  up  �v    *�  ��  �  ,�  n�  ��  !�  x�  .�   `� u�	����Zv)C�'ll\�0BKz+��D������b�vgى�y���yfY$E+�\a 	 ,�V����*L\ ����4s$�U����.���1� ����ц���I��=6���`�� �OοZGx)z6��M���Z�Ԏ%�D�S��Z:���ٱ.��B���:�����0g�Vg�7[,m)�H��\�N<�a'�3V4p��U�� �T��d�hĘ��"��XlZ�F ��IΟ���۟��	�n���qA`P`��$hՏN8R ����h���!����h�O@�d� �'�|��O�xc��A�g�Ё�Uj�B��ԩ�.�O����Ȧ��	֟���۟�&D�;�\Q�Sn�t���>�6��� 99kb$Q� ��;aKt�h�'	T����O�� 	�t�aE�P�:����-P�������e���?��D�=0�+¾�yRH�O]��C*��|��#�*܏�?aŵi�R�'vB�'��$�'���鼃�/X�_���8��/^X���Q��K@���M��i�j7��O�ѯ;Z�h� �if-!�l�,EP��PE��t7"�¯	VF(0�¼<�ش��V�'(��@e�6t6 ��"`�6)F,8Xw����5YpJH"5
�a�I���P;=ʼ���T���pF� _7M ���;ٴ���8�T���M�/xH��J �N���p���b|�=ɐ�i�B]iׂ^�D�}2ѩ��'���l�`�:�;Aȏ��۴<J���jM���ڢ���`����1�P ��>��A@�kӀXoZ4�MSRk^�^��`�
+��ɖ�� I;j]����V��8 ��6}x9�C�%��@(�/�o �V�oӾ�lz��ԡ�?K-rx��Z�SD.�HqI��*�⁠Bo�
3��UB��EA�<m�(��Q�aՉJ�u��cݥ(�'�O�4�����Cr�yH�B��@��"	^3`h���O4��O$����y�W�B}��c�	�Ox� ��4'L�A�)A�f�yYb��O��d��?�
�$�O���O�%�������8�l�߼C7�*'N܈J��5)��̓@�_G�`Xq�Y�y9���_y�Y*nD��g\�f7­�7���0<� �iy�L�<����z�'�\�oH���%�������H&�h�	����'B��^>�X��	�u�IcF�X���'�d�� iF���'-�����a�O��@u��/x��k=J��A���'��I;f�v%�4�?���7�̉FHN'qS>`�F֐���В�'�"��ad��#n=,VP�E�?G*��}"��0B4av�Մ" �jӦ��N�?!N�6@A� �52B ļ5�� ��9x�5�, �B֊N�)Ո�g��O֜",}b����?y�i�:#}O��@�%ڙ7{�ۃK˳8�X�B����'Y�?�{F�_1�� ��X��� q�S�'D�nӴ|lZڟ�Qٴ�y��!~�d�f��,�I���?������*!���O����O�˓~�����	U��*4@ʫf���<WF0�#ǵv?�SuH���)��H<�W�	>
�6%�j�����ޟ@�P�0PL�Q0��-ܸIgĭ�t�'�dH�H��D��w�X)K``���D�6/ ;����@�i���{� ��I�?A���(V1`h���h�14nu1��?�(O���"�3}�@�r/>I�hC>�6�*��5���^�aCܴ���|��'�򄚼S��$���ރk���j�u��lx'.b}��'��V���O��I��K-E+��ʄ��,0�(H�2�aR	]��v�	���C�H���N@�'���	w��~��X��i�R,���O�O��1�k��A��P��苋n�� j'*Iٲ��=!�ƯQ�J��T�6;�B��VP���I��M���I@��� ����ІNÐ�#���2�Y���?���0>!ǀ�F�Ⱡg��G�8�{���H���M۳�i�剙2.bU��O���
#�a�o?c��}r0h��Oc��$�O�x��O����O%v	�|�S3h��yC�89��0��c�� s^�S��Kl�1���W31�P���Y>3.�2  �>pQ㍏����Ԁ͏H(�l�$!� ��#���'���)m�F�a� �Ĕ�
�t��t*q�
@sd/A�M��˓�?i���?��'"�;l�ibҴ�(��<�<ٌ�T>-��4VU�,�R,BC���3��V�Jx��F�i9�I<��T� ������Ij�t�
����z��h��	�&�P<�#AYanb�'����J�;{F�q���M�r��ů�����0Q>����4ގu��o��)
�U�Z~���k7ƬQC�B� ^��s ׹�0�K���d�#��OIhSdf��HǂW�|����V�)?ɱ�Ο�:ݴg��O�1�n��G瀕�����d�>b��|��'��'���'��	�;��iZ�hדm�����F0Xq�����$�pm�Ο�ݴ�?1��5;J���&Ϧ���3����'e�'�  �Al<R�',��'<�ݰZ����7-��3BP��1RH8��NO�H8�%����PB�R>I���3�'ò���O�/MP��0@ޠx����s�W0/ٺĹ��160�IB�ʎ��Z�\>E9�7�"�]�wx5��I��=�	�!lZ�Q��	o�4�$=��ON�d�O�i�D�V�a���.D�S������O����O��$:�3}�̄�J�x�ȷˀ+A����rI���$�)�޴�?ar�i�2�O���Q>���jI:]z��r�눛	K�@��Cض�LL��n���	˟,�ɽ�uW�'s��'ڴ������C����GA�T�0�i���,�`�9T)\<�`֬��f�D~�g�8xì�t�Y/S ���R6��Jv�gH��rB��M���H��]Z�nǪd<N�O�QZ3��`�PlZw�J~�I�'�u�҄eӪ�Dz�ቆ}Xz .�&dA��N?`q��d7�D�O���~b�u�ФtY*����$-�~��J1���ۦYQݴ��D�4Kr��m�֟$�W��iZd��2OD �$��~$F{��'��}�Њ%���af$�,+��4� �#�Kΐk��C��$+z��g)�+r�6�ȍ�$I�ks�D:@T�J�x����+H�� S!�ք>U��x �]�|'��Фh�)�M�@����'� P��d�v,�<)�oS�#�����3u���Ԥe�E���Ol�+��6�᷏҄��U�F9�#�'mJ6��0�i��b�(aJ��X�fQ�VEԝo�Vy��*� 6��O�˓����O���D�K+�HY)�j7s� }��+�Ox��&�p���;خe�D����X��B�D��S�t���B��I�hs�)�U�]g���'�4�jaI��,��E2��ԅo��<�C��-�4��˝ ��+L 0ҭ���#�✁�����đ'
J��}���G��3��t� �j�૶�]6μa(�N>=�C��n$ju�fm�8s���`�5��?��iz7-8���-
�E\�K�\e���/st����iL�P����X�?5��ßD��}y�^�-���yTN �l��8 LU�S�&e�0O��W��(cU��ӆ�I'X>��ӀQYҜR5ᰟ�0`HL�?�Ҍ�^���E�# *�x��m��$�]RQ
4'�L�s�r�$�1J��$��w�&t��mE�@�LJ �N��D��D�i0|˓2v���I�?����>�*��Cɞlr=��X
z�� ���)�t�U�0c ���z����O��?Q��M���}Ө�O��������x"�L�&<��� ��@�(>@�p��Y%,
0]����?q��?����?�����%T�NҖ��e5t�\���L[�/�|x֫�68�I�dH�l�v%�)+�v�\MQ��L.3����<E����@4�n��&W�I���ZCV
kX�*�� �㞈�E$D
_��(�wϕ!`}b	���7��D�Ot�=����)S<9pt��;>� �cFCj!�Al���,U�n�R�aW�^��'X�7��OX�I=���ib�'t���*�3QpP���;��`5�'�B�h�R�'�j�)fs�8���\�!�ђF&v���/��b����L��+
?葟�1�`�[Y`1��mѬn#
��4D|�*M��12C�ِe�޹�g��8����@���Y@�p�� �'.�!%�>qLꀻ�+��c?|-sH>q���)��_��Y:S!��p����Ū�1@���x�А2h��~��5ءCX�y���(����a�'�x�7ef�&�d�O>�'<\��O6,Ӧ/�q�T�e"�+�p�����?�1�>�?�*Ot�Ħ|�Op�#�%E1#�
�9J\�S��l+�.&�t��MN�L}Q?U�X
7�6��#�+l��p��>?��G�̟��ڴ
;�>�ϧ#2<�X�eP�C^j�`g,�Z����?���~��!R�C�x;#�R�'g��z��c�'&$7�
ݦ��|� N�!y��#m[>gj�1s�Q��MS��?A��^�[��ѡ�?���?i���y��Ɩi����5閒r���v���F-����?!%Ä\�l�!/�Q����ЖE�:��'�.��i�W����X��{�E8��?i��c>c� �c�^$��9��W'
�F�1`����@(O0]���'3���?�O�yQ��J>?��i�e%��X�e!�	f�'��ɼv[�ذ�"��,�`�IZ�,���4�agӠ����-�O���T>���Ŷ�(�+e,J�.�XCw�Xl����q#�����	�4�I2�u��'x�'�����&`����"����?:|���/�O��`���hi�᪇,U
ظ����^Vt���c�5I茭��֣^EIS�ɏw�n�ؔC͜W��e��f��^��1��O�m���HO>���dR��بȿb|���_�a��B䉄0�H�"�K� dM�ElI����Lݦe��M�$�i�哖Tb�P
ڴ�?�'%�i��I$BI.\Huo�M�������O6�`>�0�o\9v�]K����&&� �����ȆM�t�<�a��R0*�%��[�Q� �v�C�|�(sD~��b���U�H!�8(+�@�G�[Ng��S�c�pn��8��r|n�����M�\�0;��@<r؅	d�O�"�"��q�:��,�O ��ddW�3��XS�8)�v����<���4�(�m� �z�P�	��7D9	��0(��TX�4���O�MmƟ��'O�SƟ����:ҬsF�s��"1�ʟ$�I�EY�5���B1!��4=�4@�á�*-�<��?!�-��!c�1g�K�a2C��l~2��3����g�B�n���#g"�"�>�X�)L@�
��O֔}��b�8"8,dIGϞNw�}��OzTȲ�'��6�[r�O��'\o��a�#H�.da�.�Gʠ]&�h�IٟT�	^�O�8m����-l"�9c��5/-"��L>)+O*�$|}BV�P�'5�`����x�t�0�kN!(z��IƟ���̟��.Q3W�P�I�4�	ڟ��;&u�%	N�P�7+�m��PqB�i��ȧD�e��D�e(�W̧R܉'�޼��;���x�	BG��k"�I
3@�9C��3O�A��E�.+�:p��BD����d"�
<���;D�6]��R����OD�$0ړAq|��J�wDli@lb�:k�'/����ܽrqq�o�	W���i)O48Fz�O�2[�hy��L��v�]8">�!(%)�\#�(j�j�X�I˟������i�O���>!%D�PI��UPUN�? ِ�0��4\�
Q\���ҩ/� @ ����=���2,X8)�	-*ڑ�3��!$�lz2ċJ�'IjQ	�k��^���1���{�$!pϧ�?��i06m�Oʓ�?a��?IɟefU���@�o�05��ث0�'H�O"aK���ͬ�� ��9�,� �|b�ӌ�lXyB
���7M�O4扒S	��B�CU�7X2��זl�d�<	��?A�O��$1�aC�'��|��#�/��)q�]4��aR	��䔙��J�&��£�LC�'����//��E�3m	
���r �H���ۀd	FG ���JQ�'��!��A�;~d�G�|��A&�?q�if��z>�: ��6M<���1K0�$��G{r�۲u��p6����<
��+k��O2�=ͧ?ț���-M�� D+"e�|��e&p>6��<i&ӫ ���' �Z>�h6$ߟ(��`M�U�Pk�6�}Y2�Q՟��I�r<����Y�#���F��M#.��ʧ��'��a�E?�a��O29���EI�p�ŀ�*=:�}�7&,]�a4���Z<�B��r~b���?9��i��#}��O���sgX1P�"�$Oǚn: x���O�<xdhѹ. X�� �G��*�b���#�M5�i�1� �Xb�����=�6�iƀE�3z��d�O��D��W^Q�bD�O��d�Ot�d`�9"J�4*� j���O^��a:b�>q)��D�#�@��DS��c>a����+��Ş<0|�B�W�
�h�c������l�QD�2TL�m �,P�<���;�-I���K�� ��{ޡ�� �U� "����'�r�������-O�1���'��$�?�Ob�'极-�P$����
`<K�O6D���u��^��P�Q�Ũi�+E�����z�����'_�	7����'K�k��$bQM��OTh��I��D�	����ʟ�ꯟj�$�Or\�f�ة)�diE��r?X��у@$�&@�ʊo�2`��� /Q��x���d%Щ{c��H�)�d)�8U �1�qo];3bT���B\�}�(	�Fe�#�> $ۧX["�O<�ǟ����7�pv�]�q�.j�2��x��6M�O�˓��.�<.O&�w��r�D|�׎M,P���!�+;?��%_��xl�?]���<��)҆a���'���GrT+!��ty��'��6��O���������}��P g?s�уr��L�D�O�q#�G�OT��x>�)c��,5^I���!9�Ha����T�9kʍ��kR�Mܸ����ݻx�1Y��؅���G�o�`9a�Z&-!(a��o
�zm"���J̏NeJQ��
�'�4����?��O���Y<A2�u̎�@Y^��a�|R�'	<�j�nI8�@�nU��}���2LYM�rD2q��>S[�`e [��?9,O$��Ak�Op��Orʧ�F���K��ċ�dR;v&5�׍�,]ܾ=k���?1c�_N�H���_"l�\D��B^����n��o�(5��q�ΗlCFQb& !��䆆�X4�5�L$aE ]$�ΠVH��
ƨs����Oc>lIS�8ZڊQ������i��O��2�'���<���7f6�S&2P�dXh5�I�<q¡��,�����	O5:\����E�'iL�}Z%�B(t|�	�0��0bϮ�[C�Kǟ��Iџp�	�1�$�z�CC�H�����Iü��FE(�"ta�(��r���s�SK�P3�-F��J}�V/�� _~��|�%�x ��m��1[!C�gr�/�j��s�1Wv�9E�z��I��Ws�IIy�$ݛ�5��8�4�T�y���ڣ\T ����'5��4F�����OB�=����32)b�R`�MC�A�y�Ї,��� B�7��%:������Z���t�'Z�I�sw��I�!�
qX���D�����6}����ɟ��	����^w���'	�=Mٺ��B�I{�L���	L��}+�� :��!|O$�҆
7'C��w�Z�T/�\I�7��l{���5K�de1�̉����Fm�'5l����X��\����V +��A��?��i0h"=I��d�1#������N�~0b��/���'���柠��y��.-UԢ'*�r�}�U�q�RMa�J�$�����4��iH� X��oZ៤���B�`�JW�M�m���"R��7�q�I韄(�L�L�	�|�e˃�d��XQ"��ԱP���R-($��D�K���J����$�6�I���U)
��s�Y�@Q| ����0h.�x��ο<C�<*G�+/�Hf_7�
�Sp�E?˸'�)���?9�O�`�N�WF%z��@� "8y�2�|��'%az"(�t�"�#Wk_�o��S3-�'�ўʧ}L�V�0wn��k1L	h�&��?a*O�i�"f�ڦy�IʟL�O<�0��'H��d��>�����
�m�`���'�B+�{Į���i\�sڐ�S�ԛ?�#uG�'-��lI��R�WL������&@F4s��D#<��@�B2p �҄�r�!�%� ��M�܍8�Zi�x�-�r��	��S�Oj,a�I.��h�g��X,��k�'������BB�:� ��y��;��$�O�DFzr���*չ6�)Ԭ���Z*e�>7-�O���O<���L�#����Oh���O� d� ��!8WX���.!B����t�(�����jJ�ᓆ�|���VufO����-w@ w�V�`��y��6l�rE�@�.!H6�Y�Rz4�I?��*����=� �;w�Ƨ��<0+�&wW�|YvC�\��']2����Ә�?����?�Vh�vþU"3�R�lX�M����?1���?a��?	L~�=�0�F�@�x��P��7���}�4�?ᇳi
��Ow�$U>�KrZ$~�ԁsoޑA�Z�!g�~�F�bD 
ޟ@�	Ɵx�I�?��Iן��'V����"Q
#�������X���4�_\ORQ��r����ґy������ŧ,��!Z�%B2, `�I9K���q�ܣ\hȔ�� K?!��)�����"�[���b���+A4
�@`�Ú*Cժ�!$�''��	g�'=Blp�lݿ*08�WH�#N�����'?�U��;�����ԤoOpQ3N>YW�i��]��p�����?��M�+Y�)�Xp(���f~Ĩ��?A�Mс�?I��?���Q�T�TQ)e���D(ѶiTʬh��W���r�M�����x��I?o����j����\�yʴJ�- !���V�r�iE�v�e�V)X��(O�����':v7��Ŧ]�I&PlL-5�Ӳd^F���̈́��)�'�"�'[�'�>�c��S�7������ڕ/�lEf4�U���)���Җ���IGv1a�	E�.��1����M��(���_�r�'W��' �D�^�8�B�P��qm7�Z=�Bk[�{A��'ǆ��sMX8:�zE�E�O�$����n�͟0�97��A�~h B��D�璟����$�θ3Rj=�	��nY�>D�="��O:
��	�s2H���$����!!O��d��:%"���O �}��'ǰt)�dA�Q�֜9�Eͬwv(x�'��M��\�hQI'�j����d�W�O:�$D۽^q }��ϳM%f���S�h�����l^4wy�x�I�X���4̻_3��;��N�e 	t�[� 	`GĆ��Mc��a�l�
��=���Il��P�M�;j\��,U�@�DX��\�D"�!X���s&$��	���ޜ�M�8)SjI&O�%�tzشxR�F�'J��S��'u1��Iҟl�D��X�h	�}����.��D�	]���j����(i���#--��F�Wn}�d��nZV��?��SNy��5i���;����/g���Ƨ��Z ʌ�5b�!U��'X�'���]��h�	�|�lھ0R��䃓'q�e�"L=m\�B0E�Za��(A �YI*`�0�մ0<��<11<z��PS⋘<<����'�"ev��d��.!�����ߐN����`�z��b���e̓y���r��(x�qXg�ڏLD,A�*�ݟ��L`R�s��-O��1�έz��8�ȓa�tT�(�
Fj��r�eC� RM>��i��'uF@���>!�͂� ����gM2Q�Q���O ����?��i\��?���?	��N9��)J�ć-Ia�D��
��D�N���k����A���8r�	8�]xڔb�/o 	��ܛx��`�R��<x��`��B�#���� �Tl��ǁ�v���t����O��l��MS��t{�p�c��xΈ� _��ΐ�/O���1�i>��<�ӥӑH�&,` ��(_Mj�S�j�M̓�hO�S2�M;!�P�t�跥�Y�^�su��+�FY���	%��$�O~�'-�:�;�p�(T�&׊`��F�=6.����?��Fr�t��܇+k*<)���D��^�T�@-G��ĸ4� ?U�p��皒t	��G��=�Ĥ�ɘ����V�*8F�Q6D�*�B��=w���^bP���G�����S����$πb�hӐ�m�ΟL�Oh��Z24���C!�t�f��#��?hu���'�	��h����>a��TK�š�������yRA�^�2�B�ܟ��'����'�V�'���O��⠭O-/|j��cL }�v��N����	ǟ��ɱQ�:a�t�Zܟ�����\�	��s�ċ8��E@��\�B���CJִ~��(�Oh]��ќe�擟qOp���ɬut\ŋM��2m0���m?TL"$�A�hـHl�$�lc>���ET?��$�%)¬�bǏӏ8��Q�ë�`]�6M�Fy���?������|"L@�H�V\Y��N�8���p5�C��_���	�4F���{TUh�M"���uoS&���'��6M�ۦ��I�M�+�F�ɭ|±�GV� �B���8Ԑ��(?�ـA���?9���?q��J��?i�O�L	��%ȷVY4�0&���,9
��ܣj6^��C�>�=3�R�@/џ��h�Ze.�R��ʶM"'"�l�B1�f�,L�*�p2�=rE��&kڏmE�DSG��"Xv<	�+B)X/�\�ê��]�e��'���IG�'>����_��{��^ ����'�
L	$�р+� ��)F��S��Vo�v�'��I�LsB�z��H���61V�ӫD�Gl���rf_*���d�O����O��$w>M����MAF��b֮-kce�)dB談ŕ/si�z��Hy���G�J�c�%���(d<	�uiʀs�USq�
� {F�@1,����u-,�L��!ZWܓ	V�T��Ɵ��'0*��T�V-r4=A�Ow.d�*H>	�+~�t���l��-2�1��ɼ�y2�Y?�eh�E��E�8��� ��4�'j�{��'���'哘A��	��,r��:x���v	, �������5J�X��x3��">��%J�/>��)6ҧF�_z�ӣ쓝5�� �U}~��ԺT�zF�9H�l
�M�a��#��>jct�''
�h�S+۽����g&e�rH�מ�?Q��h�"�)� ��dc֖m�t��8A���1�"O�I�w��hA�@*f)D28.FhA�	�h���a�C �7:�6�R���ٹ
�Or��O�DE�X�*��O^���Ot�`���f�Y$+�P�$�W/�����{�R��"ǜ-1���:{}�b>�$��򦊑oQ�QI)�����!A��9'`����ҌT���"��/A�u
��~2�eL�$^dt�;-Dx��
N�c��,��+2�%�	K~B�w9����tD{�C>[�24RTz(:� M"?J!�䔠B�&ɉ�اf;8Ĩ4@�5ec�ɧ�HO�I�O6ʓz��p��B-~8�)Q���i����$i�������?i��?����?���������������[KfXB�+]m-V���G������?��Ж�I�os�U��NC9�Ԑ�ŧR�sT�)w&E"9��3��A�h��;7#��r���� 
�qO��qV���MJP 7��E����U�V��'�ў�Fx"��8d�Q�U�I?vl<�[2�*�yr�ޏQfP�XG�6:���+#I���Ee�F�'_�	�?s�m*������=v�m��z��mK�/�~����O8�x)�O��b>-{F�^�p�n�Jv+L�Ho����.=
�k�+@)[%���W��=�yG2I24ʰ�M[��.�ٔKO,�l��f�e����o�.���)��F�'V ��m�A�( x������'n�|�&
�� <��Z��Jof���O>A�K�@��b;y����L�i�(��I��?قJ�8nZ�y��暳R��e�����'4�3��'���'���52| ��ɻl>yr&�=D�`�2S+� z�BE�����ö���r��,-= �AJ%	�9��i0ڦ���|����N�-v)J̉珛{~���o���p��E�,T�)[��� �)������b}���� Y�oR���`�`����'آ9��?���i|����I�9u�0��!x�0�A,D�@���U<���Qr'T�B��� -��)�>�HԬ�O�n[�
��:Z�Uqe��Ox���O��D�� ���,�OD��Od��oޭ!F�Q=�i����P����Lbi��xF�Wh�� i�,�7}�b>�$�ؒq��6�*U�aV3u�m�a4	/��2m�nwf�+�ܱI�\B�~�T(%Z-tp�;CxxT\�3G0��c�L>L8�Y�	K~2�ؙ�?!���hO<�f�	-c��Gg,|��uEB-D�d#pO�H�ĤbEb��j^��:�m�<�d�i>���sy.���zA��5_<L��CEQ�%F�	����o�llӅC�I�u�2eZ�?�|:ļ�b�@q�P(II�p��
i��0'L�k8D��3]4u��h��&�N���˟����"\�kb퐃X�m��Y�G�"����Ԡx��ݡAPʤhgTD �j"�#[DJ7�ǀ��0���H9l!�x�"W:-��3e�$I4�rѯ� �Ji�"	%jUqO:e�4�'b��iG�c�����^�=�z-��-�f��IZ�� ��E�8�"�`��ۡu�<5{��&�O�Ȕ'}n�!E�o�p5��]Sܕ�.Oδ�7��Ov���O˧	|$4����?��8qMVH� KWtLYS��?�ׁ�	|on4 &�E?=�귫�M#���ķa��Ȼ�mK�0��@
%&L� f|�Γc�^Pr�-˿cBN`j��8S�,l��k�#	��A"���&r���C�IkL�á���y�����?��������D�3G�5n��j,��~X1��!D�DW"ۄ)u��kG!΄1�+	L��hO��D�����W%�uH'��ED ���hI7a"�'���!?1���'5"�'���O`�C@`�� {��,~%|H����9V�D �A�r�B�$
�4�D9�1�?]�}R�J��`�2!�����OC�nn���� �,�\�*�	���Ɍ^+ܹjE���~RoJ�A��5��5��$a������8j��'bў�͓.bꌉԳ�Ih��a�&�P$D�\����r�L� ���`�ɑ�`�O1Gz�O�"S�@b����&��2�����6:B^�"w	\ҟ0�	џ �	�?�I����'-��y2��
���AjŝY��� �����sb�٦+����kL�;���A%�Rd�����^'Fx��yF������<�����WX��ӂ� -jj�M���d�55�B!5r�T4R"�A,�NH�B��#/���X�'�(XP`n[�ֲ�c��� ]��'y�D�D �vHh�9I%%�NJ.O&�n���\�'�VZ2�~����T++kbt�����aU�P��?��j	��?���?V��I�J�r�2�u!�\)Uۼ�]�lrx���	�&�� �(l��#>�b�@5>�, ��9}��+���3��8����~������Cx���%�ۭ@X���tm$-D���Ovc>���		Lp�A��l�
�g��<�	�<�L� �R������%a�����	����@r�$�_ Tuֱ7g��6�	p�����ܟ���W��텅vb�' ��d��qV,rbk7T� 0��'�ѱ�cM97�ڱ@�Gm��/_�����W��o7N;LU���٬�yr��D�:���д'DM
� ɉ&9ܠ��h�+tZ����x�ֈ�~��u+�(a��� 0O����'r������S�? <���ڄV���[�n����F"O�����q�����a��`T퉢�ȟ݃�a�#\�v��8In���.��?!��?A���C*$����?���?Y�'�?�ʋ
>���+!)��1��Q2"�3?�d(�1	%&�2(P�,��E Zȟ���>�g�*9.f)��� SZ�9����6����۸S� a�E�Qhp��O�R������,�nL�2��.Dp�y�-׿Z$*��'�������?���Df���"�<b�q�2�O)�hl�K"D��0v'��Ga����x z<s#��O|Ez�O|�W���tNH�m�ذ� ��Z�\���b�C��p��Ο�	ԟ��I�?��	���'=,�С5K�=JH����ř;!f��7���q�0E�F̵y��� ��2Ot���*��Bpi�d����چg�A
tH��N�f� 98bb8]t�"����DH ���$�"$#b!�	h�I�r�*l� )��=%���IW�'9�����-"�VT�t�;83��9	�'|d�хKLxX�׈O C�D��(O�n��l�',����p���d�O��ӣMt0��j�&���%�PA`��s�����O"�2zc��AT�?�ƸR���
`5����@�5�6=2��˫l �jtG��x�6�  剙5��=B�eF�>�X�� )H��9Q�e\�y�3h�6qA��a�U�h�2m)%���c�p	%C�O�u���U@#,�i�X# :x��/�]�<A'bO�E�h4�u��7J�~��D�MRx�h	+O2yz���9�"�I�p�0��]�4����	�@�Ia�T�?i�d�f
2ᐂ�H5z�-�S�-�Ds�>)㥇� �9;��/+�xJ��,�	OJBO��p����+s��$�4� �G]g��nZܟ B��D�<�����0�I�?-�	�<1D��DÆI稁�_ Ν��2��ܴ�?��K��?A�'�����M��i|�)p��ǤY7$�Vsq/Y�C���x"���p���'����f9O��]ܟ��I�?e���<�Ε�q���)_!�㕌@%��I���arl��?ɑa�Xnz��43Ot�q��ΊX���1 �U�Max!����O䰐��';��>
���n���������?i�c�ڙ^36`b3��B9�`#D�[��?ٵ�ٟt�I0BLb����?I���gn�a�r���GC��~�q��INj$jO�M��'Dl ���?`ˎP���'���O>p�H�+'Be����y��Y6��岜'������?Qg����a�����?EnZ�e���� �G!`1p�Ӗ`ޡ!&
��M���'�y*���?9�/����ٟ0���}�aS��;�vȲ��9�I��4&n���'� ��V�i��7�������(�pm�?���F��D��Z�� �OD����]�M��'3������6M�?��O�D��;�Tǎ]����	��ė7�*C�	�DU�P���E��у��=7-�O����O����c���'��V>7-�=e� h�A�q�R�1i����v�'�'\r�'g��'���'+�I�1_��;R��X�D�A蛲Q��'J�	ҟ����T�	�ؕO��%3��Ps�<���l��sR�{�H��O��$�O�$�O��D�O��'m�(1�C̶We���4$B���� �O���=}��e��=�g-_�KX��p�[4�M����?	(O�����~�^xx��BD雾zG0!��7�Mk���<aH>Q����t啖(~�I����]oh@ɵl��y�"#>kh���
%	k�������y�?��q���`$��ybk��tm9�O<f�
`����y��X2v�ޡ�c�Y�V'��	�㞄�y2�L�`63�ΔUR�LY�%��O@�!E7����#��N�@aH��x�S�� vҮ	@
5j� P/��r���떚>rj��Ą8u�ڙ	��&o��u0�оiX�O|1��Z���:צ�(��Y��@JI���)u/v�ffZ��Y�Vo�0� 36�E�fr��Y1i�e�.@i��-Yw����`W�/���0�h ���`jue�[�@@��	�6�K�  �z DȀ+S� ��¨}bT9; ��>:l�	�aF�<��x+$���*����i�-jE`J�-,�X�@$l+���6 �Of���"r��d-�|�'pFtг�۲m�(��3I�p�~�)N<��m���O"����F�jv6r抙�g��M;M<�̕��N>�~5NN7D ����SL(cC�Lf�<1�/X�d1�`�B'z�Q�Я�d8��h��ď^��"r΄��2凕�(0�I�4�?����?!�	�a|H,���?q��?�]�L=Tк��!u6,E���TŐ�Ìy����<a�� �#��8�U!������D�V��I�{�|�����1`ܸ;fȘ>1����C�|H�>�?�}&�hB�V,:���8�I60����)D����g��l!�/�'4�h��o*}�!��|JK<�c˖JF���͇�CI>�����=�x��G��?Y���'
��'X���������|��$�*q>�ˌ�}��Rq�H	�=���RQ� l�qA%.���r$(�;6���M�C<I�V�&����1'�*+��b��%u�hm��+�p?Ѣ�P�B�V˖;�,�r�IX�<��)�"0�T�;��b�԰�S�BWܓ��F�|��	M5(7��OL7m>]��dCJW5/��Ո�H<�6x�I�Q1�ϟ����|z��Zß�$� ��Y�8(���ZP�:YIA2,O��1��Dʔ0#X0��/ױ��� ��e�ay��_��?�Ð>9@@!OB����W4O�̱t��z�<�r*�4��)�"L�.]�1��p(<�bCB5(0�X��ɸ#�6�PB�4
,U�J>��G�;���'�rP>Q���֦B����u�����ݟm,�Lx!EU!�?Y��0�M�łǌ 45;�։r��t��I��WE~�q���Q2�F>L�l$���	1DTY��xR�C_���
��x'�d��o֐z�8pp��S�TcJ�vs��+�+�8.��@���ēyu&D�ɝ��S�,rY��#
F�Ju���EZBi��u��ժ5�D2Pz�nMrĖ���	��(O����V t�S��W6bQ��wb�M3���?��.(44t!��?A���?a���ӑJ�*����ƣB@��t��
ϱ��'�zġ�0t�瞐DCvlU�>af0��>�qɕ@X���w剦6��i#2#s�
%s7ˉ:D�'�%C�S�g��<!�)۱��pmL J ÚpUFB�I=� ��qI#�@'d+��w�>��i>q&��#�� 8��A�ċW�{
l�s�*ĿZ88��Q��?)��?�������?Q�O� ���@�L+�/'w�h4с#��xrG7:���u�_	
�������D���'�8��'�,�bĉ�J�.IDYR o���?���'\�Sj��2��e��ޣP�$e�ʓ0��!(ơ?������/����=!�i��'�N�"uj�6��wӈ�h��5i���H�-+m�ZD�������
����	ǟ��	�J�*���J�~ej����Pd��� �uzܲTj�lڐ��c��c��D~GZ9k����C!���R��:3K(7"ͳM�?VU�R�C�+țF��iH-h��|b�=�?Ib�i76Mj�2�i�~'�X25��>._l�rQ"Sgy��'��|2�'���'�����c�1�"��>V1k�H+�~⟠3���̟�'��ɳ4���9ׂV����}��$2fʏܟX�'���P�x�����Ox������6'o�&�PBْL���1 3TH��i͟��	�>ؠ���@��Eq+O��D�D��|�];���=k�klM��ē��'��'��a��)�%��"+����耀��'=�P�E,ɧ�OѾ�����O����F?F\^���'Ú ��(�4N0�Ec@h�85l)��|2��	8�:s��Ӗ01�$,�N������?���?93�8E��,+���?����?�]�ĂpiN�@��Iڵ�L�#DԴy�kA���<aMzub��L[�"Y������X�G�:��	)P��a��T,�!ǎE�U���R5�|�E��?�}&���B
�D�V5P�a�i�TZ��;D�@�c̓ {H}rdҸ5�@�>}';��|RK<���L�'���h��[���f���="�bX*�H�d�O����On�	�OL�d�O��h�ur��憃�5�xŹ���B�>\x@TP��Y��k�����J?O�q)&�:8�$`��ˠD����E�sP�cS(N?!C��37nT�7 ���@�LqO���f��2)(�f
&3]�DS�&˯\�R�r�,%����ß��>�6阕S5��`���gk1����n?!	��qΨY�
�f�}Y@��&��d'�|�i{��Ym�Oy҇�4��7M�O~6��e J�(Ũ˛'/���pH��
���ɟL�Q%�˟��I�|7.ƭ;��sJ�O�ح`�= H<���H�+:By�GL�ay��D�dW�<;�)C�F����{Bi��J"f�
� d(5¨��9D���2}2�A4�����&@�J�K���nC�Ƀ}�>��E�Hh$�8�!�NC�	�?��0Ѷ�I2�&3�oNh:�(��LS�	,gvН ߴ�?�����)P�h�6�_�Vت�3�	(�:��SR�������zA̶S+8���8f�r֏F6#���~b 
�l�D��k� 5�,�@i�	�6P��ɱc	"Cz��طJU�8ꖩ���~t���J�L��$◞J�N `W�H�� ɹL<y��П K>�~��M9^�h%��8~����f&y�<��� CN��L*i�4U�p�_8��򤐖.����@H�w������;="��4�?a��?)QA!{� ����?)���?�]�l�q�d��%�2=#��q��I�R��z���j3�(6Qp�3�[0���
���O8Uµ$�7�������2.?$v��1h"(�P��?�8��#��c��UB�S	���3�\��{�? 0E�#�w*a����;h��m@Ӱ�M�2[�Ds���Oq���'���ʘ�l2���'4� �I���_��㟸E{"��?	�l��E�p�[�GT0=̈́	��bAl�$�U{ߴ�?��i�B�O��tV?ͫ�E.:�q0Qa�1`|)1��<[(TK�R��?���?q��:	��O��Dl>q��^r��dn�_oR]�&�_t�(�#EW8X��L�f��k(i0����A�� �]*2 ���$ҵ�Ip�/*,^%rs%0"�]K��w������ Vo �W�
0�Җ��^�F�`��O���I�y�\��Ɉ�eۨ�ʠ�P�]C�B�I4�Ji�_ �:lܢC��R�>�	�M�J>�$�I"}��ĦU�g� `��2�մ��}�\��?��=�y����?ٞOR>@�0g��=��-�u�Q�E	��&��UT*1y���He�aS�lY�^�p���C�H�'n2Aa�1*��̵���;'κHb�A��#�f�R�Z�R@=ጇ�Rr��<��۟$�Id}R	�qzx�aG`W
N~��v�(��'*��'�(�"P!*�1Âc1��P
�'k��0� �O�V<���A� ��PB"Z�� �D��MC��?�(��;�!i� ��gyQ���֨X��Y�%[�R�����ON�SC��O�c��gyR�+ 7�p"���&E���Yq��2��n匕Fx�����6c ��o͸.�|q�`ś���rY�������S�'kp���W�l���p��[c�P����!���8T�Cd�KٴP���5�(O��a�eփ�\ȋ4��*ꡲ��W��M+��?9���~9���/�?����?)���-���
1`�� �;X�>���N�>;̀9@���:�Je2vʃ�R������$Πh�\-�I�s��Y�JV�j��
� @��U@$�7ͼ1مH�k3��$h�V�'+j�[�9�f}������HW'��R�fօ��$���)�3�d�/�8u���\(Xf0�X� VZ�!�D\, �ĽI�94F��k�oL�=������}�Ɇ^�3`�Z�f{6a:D��*ecmp���7S�^�`��?Y��?�p�����O��Q��kfL�3�vH��j
�2t��ӣƻQ�98��ˌ�z,��	*f����=p(6}C�gJ�tH�so�!Z��AƟ/zX@�h�:�Q� �C��������i��K�8H1H��j����Ε6�8q�ūL��1�%$D���&Q�`�lvL/��F>�I0�M�L>qօ��F��	����%��H�7c
%$$�x�$ڎ�?a���"�0��?���`�q2(�K�af�E0@ �I�#B�`�޶0�У!jV�џD�a��@� x��4f����4�յei������S}n���U�i���z��35l�P3��8�ɚ6U��ě�M3ߴ�MK �.v��r�B����r�K��#`ԗ'駑�O�
0�L5�������,�f�c%`�O��d�����%��>��A� #��Ac��h�r�H�#��25��O|˓H�fպ��iF��'O2�O�qsq�i����*ZaI���Nھq��O��S�Yܔ7M_,�0���+��f�*�󫟼�'����.R*F[h�#�˧,��U&����y<U�WfS��K�OV�')�(��EG�M��\�!��O�m$��ƃ�O2�'�b?r��6=˼Ѳ�#L'P�;D��hǥϔ=-�A��T�4E�yq,OIGy��i�4\���HR,���_*5d��oğ�I���S����E�	ݟ��	�����>�&��eF�-�@Aا뙝$/�� �kR�ax�pa��l���Q"�]�'^�FIH���O0tA�b�3FF���]�LTx8���s[�<Sw�ȐS�]���Wt�t1�j�Dg�=�6�] ��*��� _�xk�K��e@��|���?�}&�0�GKI�P@�3�
��<�ì'D��P�,
5E�	f��aa�ke�'}�#+��|N<!ǧ�8�tӁ����0K��Rrz�`�ߩ9��'���'�ם̟����|*��]�_�H��u�:��!����u�M]�]�� �Di^�#*�qa#
P�_��<� �,�N���=tW�!f�\	@��.��@rt'ҙY��c��,�Q`�/�}�/�<IxQ��L_��^q�����ş�Z��VA��EaT)?�� S�:媤��U� �i�J�Y�u��v�t�=A��i��'�R`xgeu�F�d{Ӕ�3��*f����%Tc�L�BY������b X��I֟�ΧE�ژ)ƄPϾظD]�D҉���y�F,��"��b�v���� ��Oj-z�ꎑHF{lD�^Ӣa�'%@����ᇕ��H�z�
.E3�?y��ޟP�M�p���H}�����䅃�T����4D�L°�"�!��Dɾ\�gj2�����E�,�貊��Fvq�#A���&�@�⇖�M����?!.���Y�FwӔ�P.B����7)� 
ª���G��d���_�ꙣ���X�����?�O+��%,����6me�칃nB�f�OD$�0]�rb �1p��B,��|�D�N�V���1�^ǹa[�lR�	�$ܔ�d^�)�3� ^�bcñ MR�gÑ���@�"O&����#�&����B,MS�H+%�'�p�<�\��h�����,K�
��pn�2W��7��O`�$�O�� h�7.X�d�O����O7F�k?�ܢ���Z|t�z`�02����M<QF�2a���|&�,�m�2>��`���Q�;"1���Ѫ ��)�`Z�`������ē��Y 7���9©N��i�eM�
��'��i��S�g�Ɏ%� �&�ػHG
I`/�Sx�C�	�l4Q��*ؾ��5�#d�7r"��'��"=ͧ����J�H�L�&�	�gۚ}�Q���~ȡ��'��'�b)h݉����ϧ��[�c)d�\�#��?^���P!C�CU&,s�I_�)^ʼ��B����O���G��x�QHp�L�C���a�@G��6��h��B����?I��K� �ƭa̪i��xD�Ʋ@��������L����O�V��v�(P΋
P���'��!u�|Z.���&3�(s�{��l��$�<9@
�ke�ئ��bR�~W}c0䓡��|��nנ�?i�(=�-���?��Oҵ�Ѫ&��,ұ�ڨ!B���� FL�r���䜡���!`�џ���\N��2c��d� 9��o�0<fTdg`5c����C�\����n��;���Gx�P��?a���$�4Y0Pa��
+\��g��{�qO���7,O��HrC�T�@ �d Y�y�
O�ٺ1���6�{�&��U
�q��*k�h��<��-���S�ԔO ��r��i&�$aBހ6�8��2b� {�`	�f��O ���Qȹ�d��yr"�A����O��S,k���@R�P�,��D�W����O���)U Qj� +�k����>��7ۤٓŪ�?�2��۰ T�Oi�3�'�b��ަ�H��_A��%^�m�je
-�ǐx�"�ಕ��� �<h!�p<1���6T�`�0���t,ą����M�e�S�i��'��#[��@����'���'*�;u!&��w,�/L��L+J�Bo0R�Ьtay˂^W�5��w�F�1�����'1R �p��J�o`!s� x�ʳ��,p��Ov�����ēb��Rq��V	�M�"��t.X��ȓ�p
��۱|y��[C��`*��O�Fz�O�'�|A����V�r��Vb�2u�	,� Z$$,���O���Or���ﺛ��?!�OD��J#ꉳd[��S��w/��1R���<˘ 2�c�GX6d��� $]k j�{�'�L�kK%x���+Y�h�q��$ٰlKC���֌�l����Fm�'�f�q$�G�q�ɺ�  �+K�|y����?Y#�'����è��XP�Q�k�03:�d��'Dاd�IQ~�zh �0n�ڋ{�o`��O��@6q�F�'5��a�{�8�k��\a0
Ë��9���O�T��`�O��d|>�R�Gj,��Boաrm�7��/�&``��ˎN�.�
N[ưhSb�L�A�Q��`�kǎx��\��m�l�R�O�8�����R<$������&Y��|� m��Q�@��J�O���O�����A6��) Ω���W"O���g�H���d�)$�̭�a
O�yڃ��PV�R�Ꮻ'��ШQR�@���O�m^�O�v�'��S>�谯���(��ɴ-q��
���=�vM�`.K��?���h�Tl���ۼ/�x���)E/.J�:�l�%1��򨟨0����r�%	��D��}�Óxb��<f��9�q�I��M�`�Ҳ$~����/��X[w@��ȗRv�P���O��y�M<��%�Ο�iJ>�~���2��I�@�0鹵Oj�<Y�l�Ro�� ��)%��1��N8�@���$ѧ9��tQ4CC/2<�|p���7�M��O���O���h�)}B���O����OGD^׋���6,9qjB�Id(] $c� v2�#��'������i�L��O�ȕ����rN�RX�`�Q�L���!��9��!V ŁF ����/�Ԋ�2z��]#e�6���ۛB��;���R4"�ieT6-�O��0�Oq��	���Ib�P�M@d��-V�,��uѴn���hO�"?y`�W}8tZ����n�\�҆�l��T���:�4���J�����T��.�@tO��ȰBp)��w�HAR�M��~��l�	���	���H\wPb�'��-=�Ye��Q��Q�ԂZ%1�}��B]�r̌�g�P8uHt�c��T+YiX��X�b�๺s�
�p.�Y����&���I�-ӫ�����"҈7K���A��T����o�YK1O���*�+�c�(R�d���`��G��rl;�O��1�Я\�"*��A�&%��"Oĝ�d҂vc�� D��&@P�D��E$��� d�ʧ'�����!۹1h�:PA�6���=�ۓ�|��L��=.��QW
�q�2ͅ�k�rP��HC.uNH؊B,�-q�Ʌ�8�B�"ף؛}'TR��?�����S�? ��� ��7�҈X�MZ!I���E"O.��5蔿_@�J�oE<Z:��P "O^ة�"w�u(�o�/)�Ԉ#"OX���Nkg����S�%�)a�"Oܰy��P�ܐ��e�d��XӠ"Ox|�/�:ɨ��eJn�e�B"OX�;���<��r �˕��e��"Oxyt�~�U{d �,P�����3D��cb�e��y0�MR��bL4D�\q"��\3w.�i����-D��ЖE]x+bY�b˴;��e�4�/D�DR����0�z��@��ji��X&�+D�P���3d�x8ӅźD���1D=D����ߊ>����l�V7��3@�'D�XȰ�O3 �p�$�%B9z�s��&D�\-�?~����_"7�p@�N&D� �uf.}ԑ�Q���xSŤ%D�����
3x�x3v���T��#D�LJ�k˪���� :\w���	!D�T�V��;k���BD	�N'��0�!�T�Z `$���ʃW�x�x�L��)�!��[Ō@a��G�>=��8�!�$J�2���ZfU���0Q���X�!�$�p�& _�:	�Y��In�!���{3���mA�V�d����._�!�d�#�R1MȂ^��\��[�z�!��W�i�KU�2���b�@�!J!�D�_�Tq�G	�P{P]hTO^1!�^R:��4C �Nrl��Mk�!�䋷?W��c�@��V]A �ҦT�!��ݎ8�4eZ��A4MHBwK�!i!��X��<���7KTP�6��7]@!�DB3~�,��d�,&�yx�IX'u6!�I�*?��: AĀo�0��k߉�!�A'��1!�o��YڼP��
R�H�!��ߒ8gj�Ki	zD� 񃍑a��$��,���R���	`���@��y����v�����f��>�ydn�8�yr��
^��� �n *T��eB��yR��!'u.iT�"L���S�'�y�ET"DaP�����@v�����y���.f���	X1<�������y��$� �s��� C��� �ȍ�y�"�y��hk4�	8�⸂����y���3=�.�[��ўz�&�*U�٫�yR'��g+���e%Y�F��ocE!�dT*���wD����Ëzb!�̎R����D�Q�2p�(& �11�!�D1"�A"�ɗ Vhn'�;
z!��;�F�p�E�M��I@'�9>!�$^2!�&C�	��s@֙����8!�J�V��!v�Ŋ_q�TS�p-!�䂨	��͒�i���+���:v!�$H*,��e ��9��E��~�<�q��8NAb:�D�i[�%���Q�<Y�A�4$:�YAfN�X�RS�4D�����s�|a!�c��x����`�<9�>���f�ՃN��$�UT�<�w�Bt���z�.�V�,T*%�O�<�f̄t� $q���&��Pl�H�<�R��V~������==�,�Q�fGG�<�b�N���XKb�7.���9�*�g�<YFJ��}��X��	0y�i��F]�<�1n�c�0��%�&`,0,D��B�<� ��1 �F�C ��baE�K$zq��"O�%�4��7VW�P6�Gy:Y:U"O���Tؠ<&�q��B�g�m+"O�jӨ؉��EX�M�/4�@9!"O��`�c5'�8i"ңj-��ZF"O���3��=T���K� 6MQ"O�	S��T�x2�R�
W��]x$"Of�A�>�⹹ªN�_�l�rB"Oи��&�%�z'��0"(�4�U"O|�E��L������><ݨ�"O(	 
?,�˻l�q	t"O�Z��UWB�U����%"O�!���ݫN=ؘ"�^�,��١!"O"�)���Y-DQg�۩q��d��"O~�� ��۪d���ҟ`��,*D"O���a���i,6�� c��2�"c"OvI�S�  Zo � ��?g��P�"O��Xbn;U9$��U9Eި��"O�� %�	�.��r�K+*��%�"O�ȸ�T�.���0è$Y��iӆ"O�B�F%%ˌp� �	&x�r�`""O8En�%8�%طgF"Ъ�c�"O��!�6l����m���r�"O�<�r��ن����g�d��g"O,��BL���Ң.-�V] `"OXpӆ�`Ut���-"�@�a"O4�s�斝)�$!��X՜ܩ`"O��G�	=P�,�h^4G� t:"O6�94!S-�����h�t���Ҳ"O��k�ׄ#���!/y��0D�t� ��	�A���#�T�
0D�P`�"�6e�8��&ɓ(^}��j-D���U�O,@H ����'���Y *D��i�-ڿ�QQ�D�{041#l:D�D:$h\�2��y#�׆>�. ��2D�(#���?��"����ك�"D��P�N�&V	rW$X1&��0q" D��GI� (�ZP��L��G�W�>D��Ǒ�U�ڔ�f��
� ��3�?D�tI�f��B�\L �i�-W�F�f�0D���b&jŐ�!�@�+#�B�ԥ!D�tؓ(�'�����k�,D�> �Fh?D�Xh�m�5_I8��v�U�&dT�i��>D��z��A�x�@�sm�!�d�{��:D� 0iH� %�d8C��L��k�b>D� P��ķ~Zd�3��kc�P�G+:D�����dl���B�P�%�-D�� ��Y�z�"����m���1��,D�8��G�x�5_Q���ӊ�J��B�ɞw��̪ $�\���ZA@U��B�4!<d��4�|�aa��:-n6C�I�pg��CO�9<%@xb@�G�0C�	�v�ث���[�F�7Lנ|�B�ɵc�xmy$�#c��0����
$�B�ɐ%��M�&�W%rxzԀY�4Y�B�0
�ܵ@��\C^ �����5�B�IwTj��p �:E`�Pr�@�>IG.C䉗_E�(���St%]�6則�C��5TpNA�Ӄ�&g��䛐Ά�-�C��2l>�#E�vg��x%��2W�C��0QYȐ{�
�N)���#MX2C�ɱW+*�j��.\�\S�Oۢlz�C䉡)����VLX�x��ѧM4	k�C��0gY��K�/tj�A ���?bpC�)� !`j� �Z�j���,����B"O��8�E�g|����#L�}���2"O�u�v�ҰX�n0҅ ����pd"ONm�KU�Xa��[���S�"O����g�3����n�1W�^8qv"O�1!�''�=���l�а��"O<<p�ŧm��iJS"�">H~�`�"O`��B�@�j�p�`�7Rd���"OF����H?7sP�k�`�f��0ӕ"O΄�R&Ƃx��Q�N�?�y�"O��KnZ!02b���M��}y�K4"OP��SeF�~ݢ͸�l%n(��"OT��K���ƌ��F��x��"O�Ƞ4m:(=���
  V8H�"O"���(pFzL�Q�ʘu#�mB"OL�C$M��Ҕ���?6x��lF.�y�	D�:�,��1Ǘ�*�9��J�ybL̡X�lĥ:!�噆(A�!�d9^<�AG�h
,����N�!�D�1+�j4s��~��$�D��  �!�d�;��I���<��"#o�3a�!��� j�p��-E�t��u�!�S����ƅ��A���`q���j!��A8�p�X��R+�����+"O!�њf����#����W� �w;!�V7/��1�эX�~��!�3�ҭ(�!�� 1a�G.��}rƬ��([M!�ě�%� ɘѠG�``��Á�/!�d��Vز|jĆeARyU�0�!�5~�I���-,n��/�� �!�D`�*�K4���-kr~y��"O6��e���W6P�r�ƪy��\�"O���bK^d�<�bD"ӭ(ܠuK�"O>ȣ��G��3c��H��"OD����0���xv�Y����9@"Ob	��a�*3ƌp$LԞ$�	�'m����<��R+A~E���'����cB� ��I�1�E4}�a�'��@�kW�Y�>���h[C��U��'�����l�3Bs5p�+?J����'�����oݤiO~,򩖹�n	Z�'e"��w�@r��l`@�ʄa:����'����$\�u�L��'�� X�
���'yN�f����ER7LIy����'��A�A���vjM6Hł��'e�]I�/P�s$ !!����t=��'��@蘜>�f|Qc/\�PM�0
�'���s'f��(;^�s"�N���	�'��m#$E�~��B��7j&M�	�'�������'w��b#" 2�I(�'�������e�x����E=� �'�RIIC�K9�L���U.;��"�'���
��{��`'oU3Ҩp	�'�#��R%ia��2��%U@|���'�e��T�GK&I�q�ýM��d��'�0�L��D���˰2�$��
�'zv���M�Q4ڭ*��)��e*	�'�t;��C�vr�k�<��t;�'�"%��B��\�����(f����'V�H \�I�ZHz� ��^隝K	�'��l�+r�z��^� Es�'�*�	oP�i�V0 ��R�9��c�'�~<�AS.9d�2��:$)D�S�';n����_��̺�@̛�mk��� �A�s�A$�:�!`�Ҫ�^cU"OhQX��W&ʰ��F�+v��[��'���P�肍�V��Ge��o��q�A��F�R��1'v��ȓ\_����=xl�K�AяT���"�j����Q�SJ��X G�'ւ=��1�T��`���b�A���H��5OL񢊄	V� J� ~tι��nʰ���)[\���K�G^�E�J$�ȓ[f�b��+ܐIS��_�i�̉��]C�-���D�|��}�s-�)&#*܇��Z�P���8iDN��!�;bZ9�ȓ&�$�J�C��h=&d���%�
}z�CC3C��{�-H*j����O��Mr� �Q��8���"M[���ȓ6�,����KL�<��D�s�d���!*�l��-��!��	���ȓ?��(��K�k��lA@ӑ�F�����!���-\-Xx�Z	v=��"O���������?/� "O��$N�I�+@�I��Bs��y��8-Bt��d!Qڜ��I��y�dXqoT!��ȕG��`"
PF�'�ļS�� Z��A�ޓ8&��sFH;B�C�Ɏ��\&:&�V+v�Z<Fp�ɥ!���a&aQ�)�'Hx���&��j��|�Ï1PQ���ȓF�4`1��Iq��p@n�5g(��'x�I��/�#2ۮ8aD�'�Ƶ��oҍ@.P]���<V�~,:�8,*�Zp�Řv��b��&<��e�J�n�� �	���D���k��S��a�E���J���X���7�Ǡm'('?5��iV��хՖP��A��N5D��3�g@1<y��qҮX� ���yу#����?gm�4�a��"~�	tp(���@Y`����������Mi��z8���ׅ��?X��ܴi�>�G�|�ѓ��;<џ|+��Y4��yh�&=��s� |O�m�w耚}7})�����0�q��{�xp���؋]���D#�ʧ�T�DD#�Cٛ4辠��o7�	�o����q �����oܧA2D�(1�d�93n�	!A���R@8D����g؝a�� ��EY:�.mcrG-L���"��zٔ�ќ'��#}�'������t�ڐ˱��C�
E��'�2UXr	��q��rP�(H�;ٴJ�.�P+޶�JQ2<O�+S��^��9 �!��'wi$�'�>%���� m��!R��X��t�v���}lAC0L��*����Ѣ_�*��~��q�z�Bt��K�V;��>��'F$���3T���1�%r. Xa�~2��9,:���)�@�@�<)�.�I�v���"�>=��ɒ6�E�"mb���eǋ/���ї�)#^�E��'ER��(MB�zٺ��M�C�Tв
�'����H�@����)T&�l,�V�/_���
��{Bd ����F}`˟u&h��([2)+�4K�X��0>Y��I*$@�L���qi���.�8I����Y
��t��_���?9E�?m��!3�h�(`�p��2�R�'�f Xv�>Z��Ab,��@�Om�E��&�(D���P��5I!.���'4pY�	A)�:��T��H�����4n�0 
'�B'8ʝy-O?7MZ�B�!!Õ�i����(�-�!�d�0@�u0Q�Ų�)�<�¨�/O*<�\v:Ð�N8�p<ɧ#��O�@X��������s��l���I]q�e�4eL�v<�u�������e�d�P�IFth�GT7Y���b�T�l�e���dط|����e�ݝ[U�G��7#�乳/#�nD�ଊ/j�>4�S�[�p���fS�sp�ҒNUIY�!�d	8)*���D��*���$A;uY�ɐh��1Ozɑl�$��yi��S�oRıR���ħg�(!a�V4a�*PY�ոF;�̇ȓG�hi��ΡE�`̙D�1 Odyz��΀VZl[vΌiD8n�<�� <�'��Q�ث: F�wg�6�'2�Ȱ�VG�"\�$) �,�^��ڴ8Yv��\�ޤ���ۻQ�dG~�	�U�(�*���I�3#���0=q��_�$ɘ�C��o���� PY�W�I(!n�TH@h��6�.Ց�5Z�����#6"ArT 
�LQ��B�p�vb�LP��J�P��(0`'4g����`ӉOҘ����N���e(��怫	�'WƸ1P��%70�C��̈�ra�#�� [p*tKL�Yڴ`>eI�O��!�a�dQ�I�^	�mI"O�`��C&UOԐ����!-̰�i=�`ɦ�
r�r<z"��	޶����$մ�������c1�Az1oM |�az�	ա8�����"�J�&e6	�}(X�������J���`�څ�=�O␐���}l��ca�HG�8��d�hn8�/i�L ���/V�N|"H�x�K��P��:��t�i�<�� �?]���� �ꤐ�N3lH���A0����Fڦ	`��I�k}b/	�,b�$�?~|%��厁�y�	ɂN����wC\Gx����<�M[�M�~��j��
�C�=��HB�'��0��_[|�9�`Ř6S�#ӓ�d�p�fD�	<�#��^�]��mH7Bĉ�G���J�\���Dӕ�a��IT�P��/p��Y�L��ߘ'0p�X�H���q��@ u8���tⓧkr�c�e����pfiϱXC��'y�Ԃ��	f��ʠË�E��}��JH=��a�bb�,z<6-^k�O��dBڅ[�,F�'����e �0�ȓQ0V��C�Vyx�I$W���o��t	�.�#�v ��nإ[��"?Q�K؂w��,yВ�0�CY%&mR���0��H��<��1h�N�>AK�b��ߧz0P��C3
=0����:6x}��	�Gd���&DĖ�b���?E�c������p�{F�:N�l��)nӉO��@hA*���ܺP(��e�H<��'7T�֊�>P�Ё�s���t�H�J�8��
�׬L��4"�>�OΨ�r�V�)�#s�� a�b�8�"O��kFK¦|���Y���O�v���i��IٖK�,�p0C��ߞtXB����䎺#�μ���0&1h͊��5$maz@�8����Ņ�NՁy�r9�6�U����S��rݠ�{%-��J�����ʐb��&��}�z�����5w�!�$��x���"�A& ^��=Y�'a��#�
YT� f�VG����'�nqH6��eL,����A�����'��8hu��	 ��J�>�f�ӎ{B�W?83ay��:!Mܝ��%V�4��H� V$��?���a
�#�F�0# ����y�=����](<9G&��k�����柖 Hx<x�dy�'�"��R��	���>��ROH�'�T:���"����uL<D�|pr� �^\h|vʹA���ZG@����F��K�� J<E�d�,,J��m�8m�r��y�.A�:
�&IE4̶%@�o	���d�U��1ْM��<Y�K�0�.e�QG
�@��|Q1o
D����3�g�ZTxV�8ChP#왹tI�᳅�[���x2��	!�(ѥX�N�`����O���')��@���� l�B�'HY�8#�03yj�۳i�6l�¹�ȓ0����	�5
gZ�������l�۴>��l@p�ҹg25mZW���G��4<7�T�+x��Qc󭆔
�4�ȓoa��Ce_�8T���1"��� �䉣�'I�N��كD�-QS��g�'�L�(B,�4t!�a�j ���$� �SKLS����H�)E@�`pӉx��
�K����@�	��ar�{�R%K�m��W<����#I�d�0�Dy��);R$I�e�������+Y�$L��=%����ۻ'v|��bD��
OB�ɾ!K�4�d`K
D�HH
�#�<R��\3���B���� �2�·)՞�h���D:4a���Q#H�XP��d��yb���[��D&F~2ؼ����l�a&��b�#��~{~-S�Oᑞd9��} �4|w����%5�O�i;![�l�ڀ W�7>�.7��.�Ī7��12u�q��R��>A����fX��W�g�L�KE�]Y�'o�!�r�X�#��@��#� &줔O*LĘKU:$Y�L��fC�e��`�	�'8��y�oƏ""�\����'xf�*V( 90��r�i���蟞�[��@c����Ǆ"@(��!%D��K��� q,�,���&(eԌ���R�DOn�ݒ|h�VNݨ[k,�g�'G�i�1EH�q�t;�M��kW6D���MQ(��� � @�����F�� �T��>�������?� ��@G�[)}�0�d�7d���@���,4����կ�!�|%>�����	T4Ѻ��4@`��N/D���S@}��'��"E~A2v�<Y���0���I>E�t�f"��+c8�h0@I]��y�ǈX�R�A�0Q�2�lG>Ѹ'։
��'�>�Q�Z�>>Q�Ώ�D��+�'=��c �4��(��AG�Bwrd��'��8�h�7����&ѡw���'� ���
�g�69���Ǆuj�=Z�'�m�G�Y�<pɚ�n|�( �'[�8�:xg�cӯ�1Z����'�d��͓3x���u�Y	YK����'��m�U��B5ha@��^�L�V�r�'Jvd���@���B%���Rx�P�
�'�0,!�]Q�2��#Y�Bq\lC
�'���r�J�^N����g����'�Ly�B�K�DCl�AuӕRJb���'
bE+r �:`�Ee���=�����'Q`0a��5b������ z�� �'���k���6��X$��Uy�]�'��q�p$��S�\S�b�Od���'�$l���$��bwOP�p�Hx��'| X��DP��<�FB׃mU��;�'�ъ�+|cƠ݄h�$�b
�'�
a)�oA$?j�9�1���IO�0��'��C�-
�@|f�q�>`�+�'�~p�"�͜b,=
1����I��'@��F�J�e�%�qF�'}.la�'Ä|��֓C���:��e��H�'��t:�lR�p)ԘeS4gi�Q��'t��i�(Ǫq��eR@��'�����H�y��4r3i�O~�!
�'ͺh��L�~k9��·���B�'�"D)��W^�$�U�����'p���&���6XT-^�I��Ĺ�'��Y*2
�u�tE�+7��t��'F ��R�I*��r�N\Uêm�ȓ9�R%p&�Vx�r�Q��<���2���
�X�l�f%��Κ�;�(��%�@b`���:* 1�R��&��ȓE9�Q27dΡ>���¦l�4��U�Ja�HM:���'�S�d0 Q�ȓ
�4١��uQ���w,V����ȓM�]�"�K�x�2\�g��<S��<�ȓ`
� ��Q�L�*���6}I���Eٞ<ib�O9^�Id+�4Jb����49PD�L<����dj�)��Q�ȓp"�Y�d�1W�,5h��dT-�ȓґP�$C*�n9!�D�m�фȓj�j��iR�s6 i����f>�����l��Z�B�*��#��'%�X���#)�Y᪔�>+*�)�W(|� ���,Д���F*]Z�}Q"��#2���ȓLpA�f��@]�,I	�*|�ȓ8��s@O�k "8J���(�Fɇȓ_82���Ƚ k�أ��4��Q��xn�"�� l�l+�-ɹ&�x ��S�� �T��VR��1�C���4A�ȓQ^<����.6F�!��
0*���}o�q�⊫O�ÐH͍v݄M�ȓM�ld#K�;m�* �a�ߋ4٨��ȓf8D2�IF~�����+�*d��Y�A!s�Z�E�  �O]" �U�ȓL8JC�P�i�)eH>r����S�? �$!��v����P	y�8yx�"O8��@/��v���dT��4�2E"O0�!Fgʯ�^�S�%R;-��;c"OB	@p� ���rQ%Fvv|�"O$83�ʩ}8T��k�OΨ"�"O>]n�
+�\�QLF-*�ف�'���S���e3���vAX�i��bZ�w��T�K%�<��l�����g�;(��b� GQN��ȓMw9�$��W���:���8.��ȓQk�;t���Dq��6�	P�\܅ȓ+�8AH��� D�ćω��H��J��C��)K�pu�a[�~*J��lb�)o�v�x1��N?����w㘩��'�
`�Ȑ1�<'�фȓ�T1����/'`f��d���7RH�ȓ9*��cP��84^eh5f��|�,L��"
�%�B,]|�`@��5�8��ȓ5F��f͏81q>4�#�RE��d��UPRN�Qz�c�M��"��ȓ::1S5�g5�P{B��U�l��e�(��D3u�
�y���J�E�ȓcj�;��
�7о5	���) LȆȓ	d�z�%J�&�|%Y��H;��ȓ	��9�(�9<�rs	Ҡ��u�ȓQ��8	�2Hj��5(!li�ȓ
��,@@�G+o}1��4O��ȓuD� e�j�v�j�&��U_�P�������jc�:%W�Ѫ2���kE2I����VD�D��r��`�ȓV�(�����"���u�R!c�$�� kR��@���[��[��$��.��u�H�J㠼�W$�	�$]��z#p �u4h�� �fI�p�D�����	Ac�i��A�d���b��(�ȓ\9����+Ž	ْYC��(��H��]�������
jvP����'�|��ȓ>�����J���(O�wbi�ȓ#��10#�Y�=�(m�C�7uZ܄ȓ�͢�Y>a��� ���hؾ��	�'�r]K'�Ȟ~��PR��̘Vl�s	�'I�q��*>�8���Pt�!h	�'`}j�B^/0Nq!�
�51?��c�' ��9��B�hK��ȃ�כ!,�Q�'�\`��b�h���8`�X�A�`�'{�I;��υb���i��6X���'_�|��n�?,$�`b�$(��x�'3vM8�� $!� �YB�L>(Z�<k�',�p�o_.,K$4�Q��$$($<"
�'�pd@���4(氩�Q�^> sP="	�'�� �Q��"��X�g&܅�Hmi�'SR�����Gr� 2ר
��c�'e<$c�(JɌ�Ɖ0Tb��
�' bXF��#����f
n�h�2�'uT	;	-�B��vfƘnpJ�
�'��$�T�6@3�GA!7,�	�'浐��H8��`���X (e����'F�,��}h��L��"�h�'�2C�A�,X�ъ;��ec�'�VЫ%��C_�%+�	K9���'�%z!��)}m�@yw���?�2Ti�'y�|*k��9:�@��N����C��+.Ϙ̺g�@�Tkx�4MH@�C�I�x���U�R���%#U+�:"ZxC�I&5AHX�#�-)��)X���v�6B�)� �P�%�E�z�����c�V��"OX�a�k׫aRv���,@�n����"O%�fKL�|��-�S��֐(��"O���Mբ[и���gR16��Ժ5"O$8�1� J]�ҧ%Q�{���F"OH4�hA�5�m9�����Ts�"O:}�Cb���ӄ�%��u"Ol�;�F�]���cN�,,�]�"OH�y���(?K�1����
r�[�"OrQ�̞,B�nԉQL�~�ޔ�"OJ<��)ΒV�\�A+�2nN�P�"O�5�T�I5[8�0Q#���qR"O��	 V�@�b�΋5�D�i�"O�C��9~U4l2"h�!�����'�h��5kZ�� ��͒fSP,��'|[,�M�RL��ʣe��d��'U�����7�� L��U��K�<i���`~�"�I�:[�! *�n�<YCP�G��L�����PHXK֠�n�<�s@�8`Vd�����	��l�<aB_��UH��]����c��g�<�W'N�n���G+5	^5��o�i�<���'{,L���;/w�<bT(�^�<�cD��7�i�Rc�4:���	ƣ�[�<9���3X��@\0$뚨A$�[�<iTOɝ36`�2D鑬<��7˖s�<i#���m��a�)߼ܨq+_s�<��#�RfJLzg�sJ�Y��I�o�<Y�#��]�>U�&l��c� {�i�<AN�HZ�p� /��BT��ʴ�TO�<���H"�Ԕ��e3p���@�q�<��ʥN����qz�@�1��c�<�l��G��1�v�l>�u��W�<�!J�+
�ŎL�E����K�<�Qk�0�M��Py�<貥K�<��/R�,�=�@�	 ̭k���~�<1�D�7!�V����=`�6P�ȓw�����)9��d�GI� i�O���d�i�u��Ks����ۥo=�~bY�|q�&�;3��劓aW,V�>�u�#D�4"AG�z����@b�#��!D��A��%>���G.Jz�=aR� D�����ys��b�W�@Uƅ��<D�0�E�=	�8y��i��+��8D����/�6��	y��=H��\	�,<D���3�C���p;*��h��Q�%D�C1̀!��ICf�L�TRx�hTe$D�ؐD&�*lj�A+�"�sX,0R�>D�������H�"���f���;D���U(ڴl�X�E�<����4D�P�FC5-�G��A��U�bK=D�Z�e��N���$��G�2��r,)D���$E��5���Z�[nZ:�%D��K�� 	lJRT;�/^�<tɉӊ!D��ڦ�W$Jv2`�b���2�����1D���gQ�E�uY�Pe��Dڥ <D���+"��e	���G� �)��;D�P�d*�S��T�P	Ə!��Y0@;D��SAA�
W��@�I�2ތy���:D��{�b y���A�,�[aa:D��I����>�����l߆]h6{P�+D���	�WE0�Jd/=*��! �*)D�4��c�D]�#�Bާ<���Y�)$D��
�#^.zX���	܁!x�R�%D�� tհ�	�`�m�6"��Ҵ"O��s��f�1B"O�5��Z�"ON)�'����X�MQbY�Mر"O��f��`O�
D���B"OȰ��D� u����0%�(tbc*OJ\[���Xb�^g,���'hT�!b�"U�J����[,P��'9��s���I[�� K ���
�'�d��g��K��	CۀE�L�'�蓇�-)��M�D���l%�(�'�Zd��K�l�@w�O:��P"O$}�B�ߨO�\� ���lo@<�#"O>BG��#E�{���Z0@��"O^��e��R=|���,�gX���3"O�H�6b\#ns��X�n݋tP�)�"O�(�+Щ%'X�Qw/��jk(e�"O�`�B
3�"�J��֩*�}@�"O.eR�B҄#�tCa�I�hNp��t"O�-X7 4h�M�%�YF����"O����e�5�F�c�fY0;B�y�"O�l��hA$g��)@�G� ���W"OV� �ި�깊�H@�p�}�2"O����7[�Qk�'A{�|��"O�e	eGh�ƀ�;]sP�z�"OTZ��S�+|�2e	�rar��"O���J�
���*�$��<aTU��"O�mx�u�pC�2䶐qE"O�A�_�J+$�r�٪iw�-Qb"Ojit��!ɲ(3�`�ik��d"Ol�2�D+$�{ mɷ�XjS"OⅣ��*a��Q�k�z��$��"O"�q'�Ǜ,�b�P�	��;��k�"O�哥LZ����/��q�8�ˆ"O�����$a��#z�����"OHq����0RO$���-XF�J�{"O���.H � 8�
ǃ].�(j�"O���Ãmf�QjA�n��HS6"O.��ŤY*9��C��L�Dh�Y�"O��O!#�=����+`Ne�w"OF�i�bZ�Js~�za�WET�C"O�yD�6@}���^)��R�"O
1�"��|��RĀ�6)��2'"O�d#�	L+t� ��h^�L"�q@�"O<,��a_y�^�*�m�4%�	[ "O��4iM�B�*`��Ο3V���+�"O�F�5�������q�,��"OZ��d�LrHxr���)��}k�"O2x�
_�:"�F�f�Z=�g"O�h���#m.�qVIY�z�q13"O�M�'E����젠�V"g$I��"O�	�v�C��G�H'>����"Oz���Jd���r�ʆy�Fp��"O>� �-ؘcp����eZ�>�����"O���0�¥*q$Yóm\�Ou���"O�MFh�}��T�t��,�L��"O�y*2��
'�����O���y�"OP��m�'T��wc 5@XK�"O��;!$L�Hpiă�^F�i�"ONe2��!*�� ��˒b�ȡQ�"O�eg�jRr��E�/n���"Oh�3���1���ǤY��9�"O�37��
���e���i��"OD�{�
3k:�=Hs*�0k�|-�C"O&�q��
M�� �̐5��R�"O� ^�h&fzr��^
Y��"O��aǘC�0Ղ���
�b�9@"O����C�4�t��R�?�r9�"OtQ�� �e�`�	I�\��9:B"OV!뒩�'|�t�#@�����"O��	e�[�9�!x�(��K�Δ�"Od�bb���褹����s��`'"O0�bQ�����G��=���s"O�T�$��0Q2�����q�*�"O�I��N�}ڌB�GM�
 d�"O��3����,��#�!N:�C�"Od �B�*y&��fI�!o�V�
R"OƐ{0"[�`�fU�(��7��ػv"O@E*4IN_���Ph�,��"�"O2m�5Ň)n+B1�D�:�q�$"O�4�BG�"k�XRB�+4\��"O�a���������R!>R�"O�a!�.��.�Z	�Pro��Kf"OBXꥥ�([u�`[��K�SQ���c"Oj��
$XP��S�N>�Y��"O"�BG���E�P\�C#�~4�(d"Ot��+�*�4p�V� 6�C3"OvD8v�XN�5�G-A?s���q"OB�A	òw�80"���ʠ�ö"Ob�Iʈ�l������q��6"O|rʍ>Y�U#�E"Z��I�4"O��H(�ka��s׉��4�R��"O�us�Pf�If�E�F��$"O�0�w��|8ީB���u��A"O@���ԗV�
}��">�ȵj�"O6���faP {F���\�jY:�"O���%>61p�j��q��>�y�d�6d
�h�l:s�e��#�y�z+¢i�7D��jC�0��	���y���ZO� �E��{AD��y2��+�v�%İS�� ��ߒ�y��H�8s��0�*�Z��Ա����yB�:<�
�83�#E�B�{��X��y���4�l�r!��'4B��y�߮�y���o���{�D^%4���i���y��EP����nɴ'�P���%]��y�!C1Px�@��
/o^ܸf��y"ϒ�EV��c��"8���rJ��y�g��<��u�ǩQ(����A��yr��,&�5)�W��"�H\;�y#K"��@e ���j!��:�yr���;������w�u3a��y"�]tv�1*%�Ů&���ʧ�L�y"�¤,@����c��0y3v#ؚ�yr�p�6D�<]h������S��i��'�]! '՚:�P5�`�4Nݘ8��'�y�T(�+#�1hd�]��<A�'夠P�k�9�lL{$o~k��i�'P����G�s��9��P�yШݳ�'u�r"�X�p�ZS˅�\L����'���A��ʝ[�5y妒'j��`Z�'Hj�0d�Q�aT���d�V�5� )��'s
�q��Z���qD&0�Ĉ�	�'d��C�*���@�M�-Oޠ"�'0�Y��2w
z�q�I-���+
�'<ܙ����	/���B��|�^��	�'�ᑗ�C��M�o͇z�|���'��	a����ۑ샃[� ��'C6m �Ϻu��|9�`�=_������ �RQ��:����Cə�h����T"OΈ�����V(@�t�V��"O�Z��L�J��QgD �!q"O�ْSa�1�xb�1r�zp"O����A=1�� ��E]-a4 �"O��X*;��yQB�B�oEܔ v"O>X��M6I$��$G(rh00%I�<��K� q��:�K8q-�����~�<)�j����亖L�2bU�P@�
Qw�<	��+8;fDQ�G`�@���J�<��j%p�(`{,Q�>�)yRgZC�<i����h�e�ecS�{�`���Q�<WjŘ#��%(ܽ"�,��BF�|�<)1�S <*`l��A7,�|��c�{�<�%��ތ� �6��P�NAt�<QG��T=4l!Ũ�L
X�s�D�q�<󧖪#��qUC�0LXTZ f�<�$�K��>�[�	εo��ex�%^b�<�&����E���Nr&�Q��AX}��)�'/nr$��@�?M��b��Kz ���f�A�J,F�HZ���h�HI>A�g�,��V(�#hԩ��
�D.���	�<�s�Z�%R��r�řDSt���d�p�<!5��p�a�ɏ^P��b�'Y?]�Z�F-A��i�)�dY�Q0D�p�w�� Gb�5jU0J6����*D�Su��>d�0�.^,n�H�pL=D�� �� r���3���0�>��C�<D�� &%�:@��a��ŋ:�"�0vm<D����ӛKa`�97C�-6�l�p�$D���SѾ;�-�%�x��$D�4��v���4��i��2� D��Q&hݘl*4���+\��Qy��9D��C���.yfL���HG2p�U9C�3D�4�%�ĺ8��>B`�9Qe(7D���b��i�����8J[µ�c�7D���Gi͋�Z1b��9o�����7D�Ъ%Z�\�xC�&k����)D�����R/ĪM��ϜT����3D� r��[�� @Y���ր��3D���4�B� l�V���a�p�#�4D�H�� ʰ`�0�6�T� L�)��..D� ���ߏK�|*�EP'Zg0Y#�.D�p��$S+��BhҗPKH��ǁ:D�p*��T+�B1��ꓪ� ���i9D�����G(X��"\�6��*5D�P�f
Y�O��t9�&0��h��8T�Dr4&��)�B �ՎּJج���"O��`�㗙lk^5A��ϯ�v�aA"O���7�'}�捂g�45V���c"O�5BP���+�4�'�8AV�R�"O^�[�bҧ_��t��%�\��q�"O�`�q�8	�p!/��"�2!�B"O���.U)j�Q��#�ȳ"O�}0��@0����L�p�T"OԜs�*9L�}�ҫ:ʤ�"O|���T�L�Lh���$h�N�a5�'��d�'zZH �c�s߶�эX�_n!�䁐c�
���ټJ�,}�;gaQ�� u��~�O�,�hWT =��hÒ��^��\�	�'.�UC�e�F��iC�.�U�@��'�v��D/M�S�O����.R�fG� ��E� �Z �ȓx�ʰ���A�I0pѐf.T�b���'ᾘϓ�0=cMP(�dp���IuZ=���u�������M� ��0ƪܥJ��eZfaTR~�Щ�"OV���MlL���4f@���	hY�ش��O���# E�]���w�( M�'���ro�0o�`�6(�!�N���'�D8Ey��i6�J�6�� ��fB�l!��F�v9 ��E��i�R�B3`���>!R�ƮTbpd�D��>�x�c��W�<��=)�D�Oؾ��u3�nK�<�H�5�83#�[�<��K��G�<i�ǹ\����/9t�q��I�W�<���W�@� ͑0���|��T��U�<a��ݺr��0�N� �H,��OMU�<	�.�1��"@��9[��e�vWu�<&j��rpHpq�_b%�6&E��y�I�ʭ�P�՗dMu�⏱�yҬL�
�\<��a��W?�X	PL�3�y� �_�Y�t'�UY�}��߫�y�J,�D����Q��X�`��yR�h��Ժ6*:<l��f����yr�V�z��	�JFb�h�e���y��I >2��%n;����/^��y�� /w�@c�Rf$ ��H�y2!�)(��5!�p�TiiS����yR-A�e��8P%U%<��ibi�y��w3�칢��1~�*+�I�yA��U6�B�	�+��ْp
���y�)DU�X�e"�P�`9��培�y���"���a'� �h����\�y�F7��Gb״$=֥H�C;�y�l�4����dF=�J<ZdG�=�y�̗�AT��Dːm���(���y��D�̽�lٳʈ�㢗�y�ԑ"l�Kâ�䴛���y�K�(��E81��	��ػ��O��y¥<k�F@B`O�y����Y2�y҉$S��'�NsZ��b`�;�y2�O���(�NƢ}�P�"���yr��͊x����^ɶ�PD����y"�`f�@S�W(��ł7]!���&dxAɧ��23�°BR��	`�!���/yJ���*�3A�d\`5��a�!��L�:f|�ʥ�ՆY}V�HŤͳ\f!���'4@%S��&Ő`�B=_!�DD�V(z'C&0��9�D#Y�#_!�đL�dP��b@�\p�/W�NY!�D�Oz�-���ߝ:�~	8��(-R!�d�>#�`|[�C��P�"��푥=J!��)Y���$�Ɏn��88���9�!�$ �Pj��B�&=��h�w��#�!��[P�b�e��)��1Q�)�I]!���g�h<;6E�+��YE�֬z!�Ă�>�6\�ś�9�<iqp�ADb!�$�%�F�y�OJ�m���a�N�5a!�$ۜi;�y�'������JD��=B!�D�td�)pA�۠h|%e�2�!�D�3$�)��7MR����'>�!����2�`O�4p`ӃV>c�!���4Cg6(�T�mAfp��㞙@�!�*�;��Q�Bٔ�q�"T�~u!�$�w�a�3�Õ˸(��o���!��Դwm%������*��1f!�$��_�"�Y�G_7~�e!���N!�	����Q*��A{a����!�D�8�l-��;�Q�sA%M7!�� RGm��g�� �oHs��c�"On9��U�,K�-g{: P%"OHأ�&�S<�!y��+-A*iA"O�H�p%
hI�`F�C�E��"Oй�3��JTz(���,
��8"O��	��rk$P��nW(f���$"O�5��QCmf��GĖ9a0!e"O��e�H�T&��r��VN:�B�"O؀ڱ�9\Q4t��F��f���"O~�3�%�N���Kӹ~�Du�G"O(��'��k��AJ�̻P� H��"O�-�$J�3��l��������B�"O(�B�L�̸��H�{�ހ��"OZ�(ӥ�b!��!錵($ȍH%�'a"�]``��Ri�:H9Byq'�	պ�Q�kݸL��s�&���O����%��$�O���[�"�`�:BO�2i�,����&}E��ZǨT
8�>�P(<�O�|x��əR���k�O�"j�^QQ`m�5{��E9�E�91����/[�6�ң?��Xʟh�Sj̈2Hۊ-����jЀ)ʞ!�۴�?))O~��.��|�C�7&˒��%]�͛˗I?���xvld A�+���r�aRp	�i4`7�iQ創:t��Xw���'��"�İ���8i���J5+�0�.aI�m]8�?��?�ߍm���"�`��S�Bl�5k�-*����v�ВGtx�"3&T'5I�iYQn]�(�Dyn��W�M��`��; i�R�� M��]a�٢<�xuZ$.�3Q�����"Q�>��Gy��<�?)�i�7��O��j��H�
��/o�*@��2^ ����'��O��7�hov� #��PȒf�0��T��%�M���ih�v�9\�1h��Z-	H���P��~2&����@��?Y(O�	Y�$�l�  �Q-�eɷ"^�_OЉ�6-�A�Q6$LB:7��E�h�{C��׈غɟ���wf� �U��Z(^i(ʏ/m₈ ޴mИ���-ʣ+$�I�T�P*� �kJ�5ڴ��c�8�\c��qg��6z�Ś��4���ش\7���I��M�U��� ��1qk&�H%P�#�l��2���?Y������OD⟘�'��#4`��N*��c��W�/e������ۦy �4�?���i���OX�ޛ7�8��6�I�tp�ǄB2����Iן@����+]62x�	ПH�	���_w��i�|�*�Ô�H�l�``�cl�pf˶f9�ah䮆�1h��ņ`1���O���{�	�� �.�C���4]~=3#���(t���S�B�1�Ԙ;��3d��a�� ���% Ӧ���d�)E�D�Rn�=qԪ%P���#q�	�sKF�$x�x%���I��0�'P�u ���8=�FM�/4º5[�{��'3r�kB�њ2�����@Ov�Z7�����۴���|r�'���øM1N�k2'�Tl�0ID�*|b�8~�d�O(���O���7G�O���O(t���W�l2�􀠩u[�})�L��3120���w� �0�Ǒ�'��|I0�V�4�Q�����W�D��e���Ln;�ES�QygP Q� I-q��ٵCP�qS��d�K�"dQ�� B��O���5@09��]J� FLWlIDk�X��oZ󟔔'���T>a���{A�|��M�pP���'0D�$C�%��	<�AA��Ļ%(O2�?�i�66-�<1u(�7y ���'1"_?�Q"�ȹ6�aa�"�|(�{�x����?Q��)B�)�����d�O��'N4`�M0v�p� �N�'0�0�Fz��ؚi��&� ��O"8�#���~K������M�P|+��D�)�R/bӢ��}Z�����Iƥ+�`�R*�e?����DG	_xi8���#~
��G�O��>�Ѱiq3'�Ʈ�*�d-���m�У"�?�����T�ID�Iy�U�X�� @�?   =   Ĵ���	��Z��w)��;X���C���NNT�D��e�2Tx��ƕ	#��4"�V����cV�m�#G�4��`g��3tdp�V	�/s���8f���(s����Y�M�������>�EZ�,ψu���I��.w;Y�G�X�eqfL�`�݇^7R��C�*��d��iB�����N�d�y�L���äp���i�~�����E�k&,O\F�+2��]��V� ��їG�^k�G�>���ʩ6f�pЀd��/`9;a�O x=&�� Ǟ�K�(�Z� ܛB�c��C�ۢ|�}
 ��@)��@ M�,�O��hE��H %�8�ɉ(	4!�'fQ�hCP`�p�i�h�@�np����5#\E���X�
㪔��l<`��E�"�F*�c��AL���Q��"�N�J��QD��>��ė��`����������=s6�EU>X�Lj��j��l04� FO�q��a�$ #)��y�U//�2P34J��Y��  C��?Q��"e�~&���b�p�M>���1e}T�Q�U)ۊ��wM�1b����b����I�F����E����
�'�J\��i#j�����(h���hᢉL
���A�RVy"U�Ln����m~璽Y��TR��?� q��U���	��^�48��xD�T�G�bE�O�@H�%H��{��Y�
̸Y��h��������,�H h�!.���&��-X�~誵!�I�Rr�R�T��ŀ�o�tZI�x��W3ǂ牶��e���#�t��"GF	F�G=��B�J�x�	'J���&K$�dA>eDҡ7H��5A�̫����G7�Qx�'��(���r�&J�	>X(�& �<@:�P6=�\y���d�
��Ь&� Ay#c��D�Jdˆk¼ڦ��b��6;��3fE_�d��WTz��� @M�T��� -E��u >}Y�D0���Z��=�S�x"fS�Ga��PB�)J���Ve��؀y9� C;��-��,��� |̓b��	��5-��{��HK��j����yb+Z] d  �O����WeR�K� ڡ8S�t`V�O����`��d�O���I�eB\y��6<�m��;RaZw���$�U�Lx,X�"�v�������f�*)c���Qy�L�2Ä|둬ҡO.�A�����Óc@���')@�P>��K�O�B��W	�gi������I`�����Ioyb�'�Za��\Z�a�b��z���'�b���%�,   D
  8  �  ;(  v1  m8  �>  E  �K  �M   Ĵ���	����Zv)���P%��AJ X��ײH��a���8FĐt��%�@e�S�'ll\�02�&EV�+~�@����<K><�5"O�4��KX�s�P��FA�0L`I"�l�!��A�*�-gx,Ycħ�#\پLR�i�b��GD�:XHR�bTo�/c���ʂ��	C��I�hˏ&��|�@���RL�GI��r����"J $�#�N �l�Z���+O�2��ܠт��dtxֈ��4��"��"M�>�[���@���pq�\n�"�>�?����?��L��.�Op��V��
 �D8��
�d��!*APy��F��p>qƆ��0`�"�0	��� E�Ly�d��p>a�	Ԙa���O�;����_Ky��
8�?1��'�&5h���,?W���Q��z�Ի	�'T���(C�E׆��a��<0��4ߑ��Q�u�J�A�En~,ITE_���P�"	^F����0�	��0[w'R�'�󩈪aRb�[$^�X��u�ٸx4�`҄L*�������dGX�T{'R)-�<8��1I�}��?���*)� P���-*�E�*!�H�.5`�&�
 �� �λt(!�D4K���t쇃.�a��CD!�I�M�J>��bU�=9�f�'2ןf��Ҁ3�z�+A`�;q�D}Rd�iB��s��'/"�'�BpKf�'m1O��X���]��h��>�hX�L�u�ў�K,-�'z��:�#�,`�����7��D� ��4§i�\�a-ʮ&k�}#�KP=X	,Շ�!�ĥ�ýh��!ڭQ��E�!�O���'��4I��F	J}*����?���`�O�{�DئE�	ş,�O�*�Z�'&�"�T�
�
�aU
m�t����B@�7���aM���3�|�>��	�z@
���C@���|�c+;�S�OD eb��1P���!� ~��×�'!�XH��/ɧ��LѰ�޿',����R�ɪ�*D���B�1,|�����c!�`��,ғk��?�P���/������9$pȫ��R��M;���?Y��M(��h���?����?aG��V���-;��,� `�f�C>{��T霨��x,g*{��V�`u:�/����[up�O����I�0;�V(5�~9#$�-N�Zlq��B1�%K�*R�tU�O|��� l�	�{�=B�D�h`�ZE"�E��˓b ���	+�0=�!��7A����ER�4WR)90%r�<��$J2��z� [0��T��-�Mz��4���O�!Y �M$pt�0��]
��ס��qє'�OT�$�O��
ʺ���?	�O?����}.(�����s�6l؀H�4^<+P�'֌
�'c�Y��Q�j�Xc�[�s�J���p�J���j`����Y{�I���!7n�Q�'��@p4��qGD��򏍀�4:�'�¡[�F�`���##�ց��O�yo�z��
U�p��	��`�	IꗍMNJ�y1gйb���Pa���A�`���$�Iȟ8�$�ퟬ�<��@:j���O�#p�(�3'�@lvG{rȝ�����)�FEW��\+�-�2�x�ɥAx���n�OH�A���s���J��ʿ厸c�';dX�� �+K8R0À��a�M�.��I�n�P�j�V�Q�H�_��0�t�ƿi���'���.a���Ɵ|CU�M!^9�pΒ*�x����*�M��E�7k�];C#��Y��� ~Fr��W���O�P\(tG�0ޮ�Gb�4����k�O����J=GG��
���u���!��˺�t��<�-�p̑���sP��e�>{.�ɛ��O�8q �'�7͗ɦ��P����s�0[p��]�����o��]���?9���?�(O��D�O`�D�R���Q!�+���	�gR��IB� Fۦ�&�P�	3��I�<�������\�n��v��(RAJ��YrX�ŵie��'v�#0ဵ&�R�'���'���]�|�F��C�LHړ�ճO��:0�Π��	`�>���ʁ���]�n��$`�G�J��,�'nϴ[=�I�VO�m���Z���E���"D@0�r����L �1�P'5/TʓM�j(�ɲ�0=qR��##+��x��d3%϶�$B�I�GJ̥A��R��\��Bε"�P��4Kב��s�ENt�A���2���l֏y�B��P�����t�����YZwf��'}󩀤ur�̷��x�w
���5�S�/^��d���DA=/��EfD��qC�9 N�}2��9�?1���#r^@SN����EE&�!�(2�!!�=N��aVn��!��&]��3T�D�� u��� ��I�M�yR�'�?����?Q�O�X98rC̜wCJ2#�^��[�4}�����?i�r�5s�&E/�b 	5cF("��aTn񟠡�C�ժ5D�88�B�!�
��I0Q�.kD�a�59E�O){E"���- m�? ]9�ZmmL�䁊�!�&|k���y�N��=�C�ݟ�c�4z�O��=��J!r���K� ]("����ej���$0�i>�Fy�"�>kT!����[����ջа>9F�i�^7�D�3&B��4ωj�.,��
;It�4�'�2	c�@iӸ�$�O�ʧU?�p����?	R��#9�$y��
(H��H�]o�&�ʎ� A�Åw� ��V�O�ST�'	��1�$�Jc�*�!�$��u�@y0��mmr�0�i�;!Δ[G-���8Ũ��Ȩg�iB��V�r�ꨡb��O����'0H�O?版�>�E�.$$~�	�^U�<ajޗ�h��� ˪�r��S��H�'�#���:����T�q�b�!���$,�&�'��f�+B�<+��' ��'��c��i��Hg�J&�����
K䠂U)N�B�b� qI��(��@3H� �'�O�������%K����a��aJ�q���^|E���Xoh-�B'��j���Z�q�F΁N��~�IH��5��L��m8X�>�'e�����az�B,b$���_�~�j�A$�y��	Kk�hZ�G^z}T���GX��M˖�i>m&���ՍՏK�Pa��b��FP����&1����|�I͟��	��u��'B�'m�$�Wdİ}�<��fڐ}���i�0S����\"Z����C� ���F~b�Q ��Q��+����mz��W31@�e3�(�k�ؙpP�T����BV*)�\X��
ӓ0��'�XX����T,@œ�'��ТDl�g�\1��i�ON���O"��}�!z�JP�a�-i��- �2�>����K�'��eH��h�ҙ�T(��V�!�0�l�ӟ��۴18���'�t6��q-8�mZڟ�����n����� W�.Ԫ�G�R�H6�ȏ}W*�$�OP�Dژ�F��tgO�H����ȗ&�v-���Je��i5��C��h��i	`�|F{bL_w�Q��9{��+qؿ+����!A�?ui�7f��$�nq�#O�v�樺��	W�>��~�OE��SteC+�勅"�iI�q�'�ޅr�h��F�(���P�P8;
�3^�	�|Z<��N�F�8��Ac�W�\�N�<Bйi5R�'s�5q�p��I���T��,��� �L%w�T�͗��MS���&Mp<ه��=�~y��Ψ54$
T�CʘOXT�V�N�Tl\�їM�V�����'v.�1@�J�����ӆa�ؚ���n�x�}*a �3vU���d��e��PT�E��?Yg����8��|~J~r��~ȄG�@D0uJ�*����DX!�y���C�����Z	 ��L�Ƚ�HO0F����fu�Ĉ�f�k��P�d_�=��6��OR�DL�</�9�dG�O����O������K�7b	0V�F
��d{ I�6���3�U�tQk-�Op�����!'@@eD������Z��yֆ9�Oꀒ�I5C��X����`�@�^�(�c��O�D����B�)�JT�`	����[T�C䉄&(���UdT3l\ ���6�ZL���D�|(ҽ6�9���Ҳ)��h�ҋN��Q
�+92�'h��'�̟֝��	�|J��ٙ*b�q���(il�1�Qn� �	P�!�!~��@��.� ��攝v�<!�a�!���&`ϑ6����D��~���+ßl"f��G3ͦQs�K�(��<�"�Nޟ�jc㌱��P���-&f���,F�y��O�k�C6@�*%(�$(@$�y��A���&�ݼ)S���oD���QϦ�'�h�%A%�M���?a�O�mZ���h��J̚	/�
jڴ��Ȉ��?1�J
��򋂄oI�j���/9�O��jF㋷+��-�q�:Q� y��ͽ1Ԛi�+�.J.�,�F�X(p/�`B[w8�� `'�c�.���R K����d�<2�:§ ��
P�[ 8"e�B�fȓg�<Ȅ��"uD�4�A��U���<��䍁wE΀jŢ� ]����AIZ-%��([���O��ĵ|2�b��?9��GE�}{r�˞Uᄅ8�On�(���i]ʸ����89�*�#�Q�5��H�5c�~2.����	Va�L��,��8�0m�8b�<�	�q\q��E��MkTjA�3���%��%Yf�x%4�4M� P�hܸ��]�^˶�3"��<4aR���?���i�7��OX�OZ�O�B�󐢞98��&�Nz,x�TR� ��{y��'R�'�ɧu�'4+�iip&YU4��S�����<L6�D�OV��'���ʟ���'44@|81
�\�ۧj��^{ �ߴ�?���x���,@��?a���?	�@����O̜P��;o��� �X�����FFC��%�	Ѻ=�F7M�+�X�)�#<Y"FP""�P�3� �Ur\|���V�%ع#�-	2�� 0v��R�ٔO��,R�+0�2�����x��؂e�<�$kƟ��ӓ#�Py���%^
Lq`�U���b`�csIŒ_z�x�Ů%D�n� �HO�i%��+��a���?x0��a�K�u/��@Џȶ%*�D�O����O�;�?������L$N��֚7�Pk��==y$}s%�k��BN�)uT����.@0z��剐k�N�A�J�.�0m��͗u����/�a��0��_/H��qxD�A9��H�@���0c� h��O �� �"�C�g2��s�m˶��"Ob$ۀh�S����Ƭ�^�v���"O^�x�0@<
a����q�^�1Y���4��$�<�3�i���'t�)�"�x�2�,Z�A�Pyf��=w�fj��\-��'���1s�v��Ԇ�&���сL�$['M�8�BpX5�N0#��E��	�1{W����9�B�YDì�$��O�({!�x����}Шj��޺[���:�n�$Z�B�����Q�1OLɲ�''�#|"�@��E�*Ҥ想bJ})���e�<����v#�5JB��	��M	c��hX�`�O����S	w�H�Y�D�!h�X��*�FG%�M���?�-�n�@�'�O���bbR��ì�NEh��ڽB�\oZb%�ᙵQ�;�V�D\l, y��Lc>
��Øg�݊1�]�b.�d�� �ܭ.��Ia�a���և�C�Oc�\0W�еg��T�!e��T���1�'"]K�_Aɧ��J��w�FTl���Vb��h\x�j�6D���E�ǲ�M
� c�v1RO5�U�?��qo�;'zY*R,	#o8�5hǯ�M���?�V蜎R������?����?���j����Q����* ��%�ǃ/� 8�TbP�Z��Q)+q�x����}D�3��J���#�v K�'�)J���n��TC���Y�Q��A���7h i*��K�:Z~�;B[�=�剢-�����y����ab֍O�<���"J*�b���/ D��r���9p���臿5�X3�{�*�Gz�O�'������=	������+G*�[�N�}�5
��'(b�'P�G~���ȟXͧ&.u�'���R�N!��.	&5�i�lKd���Z@�'��E� ڡD�DXp�G>F�Y�����9s��D2��{+�3�?ag��)��Rb�F�p�!¯O!)6!��E?k7��vl�8f�03��4!��W����b@
�~qK��Ǒd�����M#H>��+�'���ԟ���v6�@	Ń�oal����ƻ=�o��b`���X��Z���b+��0�jP �@A�X�O˪��%oU�r\���H1i�z����D��yZ�l�@�T� S�W�d�z��o����ǃ4�,Q�Y�)(��=Iv�����	ܧ3�ݓ�O�S�Ԍ"UD����'k��'`=��S!��8���<ي �w��I�ː�BU'�D����Ő�v��2v���iYR�'���#��P�����B��D��Հ�T�5�b���+F��MC�X'-|z:Р[Ej�E(�K̔��Z̧D���b!�ol��:C���u�}B��os���̴ "���AܳC�,_w6`%��󉑯;�lqHX�yh���.^2����	��''�)�I�O<�	�/�e��D5�ޑ(��	(��C�	�-P ���:Wj�rs�Ǟ#��"=�����&�J��+Y�����ˑ��ڴ�?���O��耥Σ�?���?9�� &�.�Oz%�խ^8zx!Ad��<����j�
j�J9b�۝u38h�P�V )�xp�O��YU#OC�E����/j,R�x��Ee,|�#"�,!�L�7�	�Жʧ�O6P�E� �t�!�E;'d�)eV��*�m�O���O�㟴�'h7�ёW��^b�I�I�c�ń�`SZ\�q��\�&u�WLMp̶�o�4�HO���O��}`�a�����P���	I
phR�@������?����?a���*���O��85y����+@�x����"FG09�#èx\���	9O0(�I�FJ�p���#H"tAE�,R������-R���5[*��i����'n�q`g#�F�C�I�@���!���F��X$cJ:�vB䉕[�,YaN�����ȇ;u��w��&�| �:�7�On�d�?�ôg�E� =��J-	�m�mwӎ}q��O`���O���Doԇ&� �{�Z�l{���@7L�f�ҤE%��	S�
w�$���%��#Q�t�$I%5�be�CFA�� �����!B����$JD�R���!G�D��ʤA�$Q�СA��OB�D��ˎc������s���#�B]�y".�hGl�,�`d�CǁX��K
�|���3Z���",��Q7�ITV�N{�h��iir�'�ӫΡ������.�.	�JCj�,$�4�Q��MSUe�oi����B��pS�rq"nwĤy`Y٘O�	h�
R?r;05�'�),� X��'��E��^+H��@��D@�*��ٖ�'HR��}b�	 �1��M�B�ަm������Y��?!��_՟L@N>E�4�,(J�	ȓ&H�/�riXR�G�!��o�����,�)� ����Hّ��1����=D�qq���ai��v�Y� �)o���0��;k�i����$�I���	��u���5fET�Y.عr��ܜe�6a3�No3�)8f�6F�֍5�Z&_���`-���Rta���h|��K��e��A`��ݞ�Aކ����*ߢqaʛw���W���%����I�C���F-$5$��!(f0˓6����I�0=� � UA�"E܌b�`]� )>�T"O��j�AB$k$��zF�Z
E Qѳ�i��#=ͧ������a /����b�B�Q�҅)ᯊ�{��Ă��?���?YaR?��I����u"�!#ީag��}��Ɉ����Na��r�S�TB��Ĭ���|�g��X�ƍ���٭>�tT�Ŷ3e������fO�i��@w<��" ���i�,�h�C��/LqOD0�q�'�f��SɅ;)U�<�PlU�-�t9Qƭ`��lZԟ$�'���4���$�[�|@�x"Q� #��}�HA�<��JU�j���O�(¬��~}�+jӦ�nGyr��(m��6-�O��d�?E���ض-�P(!+�7\=\���}�f�
e�Op���O2��G㚬gvL9Q�ۺU�p��7
��X�m[��X:;��`1eNI�;c'�62�Q�tZ�jT:��!a�s~&2  _-�f��
�*6�DS���$e�+�(S�<��+`�'扮>�����u�OpJ�˴��0B1*"�	�k�j�<Q4�A���L�" ��6�J\X��8�O���Q��nR���ɻuq�Lj5V�p���^��a`Z����)�E&�e���3v�A5>\�E�	�M�8��{�l�*t���=���'��&�%�.D�tB��T�*���XV�
�� 9�r�*D�<2��Go��T�W%DN��%�"6D��֡\�s#@��'��v���J�4D������;�0�â� B`�"�)7D��Cs���ys��[���q�����yb(��5�y�C?=d����(�y��H�"�ȸI����3�d���&� �yR+�d�E
G�"(�L`q�C�,�y����"$ ��GYd��)�(�y"��15!0£� 1P���av�>�y2�A�Re�0Bs��_�\M�!(��y�∣1�>���ت<ؑ��˛�y2C���<u f�=6u��I@NN�y2GT�X��&.2�V ��]��y�∘:��qQ�# ZU>�т-P.�y"jW�|��]�k�1X�r(�Ό�yJ"D�Y��
 S�4� ��K��y�`�NG�x0�CP��v[��T��l�����2 r��	D���P���a�D"D�����ǜt�@X�*���p��zL p8u�Y���>��(܍*ENu��l���Nt��/!<ONt��d��GNu��'q�p��:׬`�go6;z��,D��j�;_d2�F�1x��X�7�D�P���Z�� + �#~�F�S������g-7ED�y2��W.~��t$P/���{��\� �s��W:���_�g	ʤ	��L>�Ӡ$N���eؔ8�zP
�`(<i�B 3�XqP��-	��3�c�	-cb4K�5G�`ؖH��=����*�p(A uA�[F�V��ax¦��	���5�=�0g�ڜ�cG�"'����v��E��U��"O�0����";�T��]����b��P��O�X����͐<fx�F���G�'���[���F�Q:��:�y�KU5��tQ&nNg������X>TT��bZ7�?q�#˭z��I~�=1�`@�N0A��X-%@�hG�F��`2�hPup�5�q
�;��5+2k�h��P�OX'��`-�Oz����4fYȐs�A�?�hi��I�WR�d#G��'��1ʦ]?����N�q�N)IvꂬY�B���"D��r&�NI"�9�e��?��H��<��@�F��Yߒ�K ��W�>�"|��+]�fM���#����p��gg�<��#
�$�|`0�`�_�!cUKՃ	��K��&s�Va���5T<&?a�<��4�� ,�9@,`$���~<��/Tq��0o��vT�K@�ő>�)A/�-spFii�I՟Dd^��d��ϦTc�͒/a���B�� *ax2�
�.|��g�5j|�R�CA�g��y�1j��r|Ua�˚�^M���'��%�'0Ϩ��q��(x  �K�P!C댡G��AROǚ���E��4;��{U��	.j���?�y�mɓ!7�@1@�_(	
PY���K�\�=v�4C�����z�ŉ��L>�� �(
<\<�u-�%o�PTC#��Rh<�bK�
琁z�=�48	c([*�u�t	�7�i��S�? i��'�ej�y����B��	�&�'Y<�K�NQ�|�'���X��4*)�@*�@�$J��<��'�,pc X�P"}k��)GR�P�{⇄�)`�ia��<��S;E��9����vV81� ���M����pɄ;>��5��{�<���7�UAd�ϻ5�"!�3��=_�
P�q�Ud�z�Zq)2����à�M�|��w�)�a�KW��X�Ɛ|v�M`
�'@�`�lֽ}� !�e��1T��x 6����5�i���2��#��'`qO��@(�8sĄ���c䠉�`�'b�`rf�>�"��T%ىN��,��hW7琬�!+ںh��fL�2M�����Pyіi��[�!t\�c�U*4�Q��i�08EpE��ܥCq�xӢ�hԠՉEpl���Ȃ$G���Kc?D���C�;js�!��- 6@~�M��l��P��AMA0�qk��FKJi�#�u�Q>Q��'ħF� �K�Q�RuS��X�<��_�W^��@�J7��h�Db�z�y�A��M�ĤPm�Ȍ�J?��{2ٗ�v!��l)Hhr���g��p?��E�0D~͹V��<��jDG�?S�Te-��Ku
��Q�ٻf4��2w�'5�t���ۖtq
<��:;+ ���A�X�<mH�ȓH`���&"ou���:x�"��C�[-����ƌk�!��,h�d�U��
�X��ɯv��$��b�|U��n��<�����^3���ɇ�:�ę�%o�?<�U�$(ֆ�!��X��8��_42�b�k!�6w�N`�a��
|7�X�Pm�P���?��$�ɇ5�m�F��D�B��6D�����=_Vl4 JS|�m���V@a��BqC"�1ǣІJ��e�i������	Y�� c�����&�K����7M "fn��C�б!��mZx��h��^$����%S-���ȓ{����`ԛ8� �y�@�t����&�^��M�3'�ܠB7A�-p�Hl:ʧ0�rh
��ׅg�XL:'�9�H�ȓOq�m�E\g�x� ��s_H���Ʀ6�q�ADǩd��O������+�'�M�$��'�2���)7�O$|�w��*�R����~��i�%Oڔ<��!�F�9ukx�e���x�$M��I��h ���+���D��8C��>����&��ə�F�(m4L��1�QΦAÀ�XK���P�!C� �h�)�$�ȓ(]V3pk�%z���'�*:�e��{+��t��/�PP�3*S��m:�'e	Z��	¯)��E�ő[�$��f�PA;NFP߮eCmZ;v�0bD�C��ߴ,#(Mj�j6��ӧ˸'I���&ś[����Tb�J�v@p��=P�%�AH�25��*�mZ�]��I��Q
Y Q���r�&��g���N~�zb�
8z�xuE�3a�m��%W���O�Q��O�wt�1BצO�`�i*�	b�jA�,�H2U��! �`�T"O�m3@�[K�<��E��k$f��6�OL�[0����]"3'W��6����(��5��0 �M&dY8Zh�@�"OP�!�!خ5���h�芩y~�""O,��V`�XG��0�)CtSu"O�P�2�ǐZ<M�� C9;R<��"O(��aM� Ί%��Gޏj#�!���'UF�A0�O�d�4E��:	Τ6�Z��i(�"Ot���{�h�G_�@ɵ�	�b9v�3,?�J~�M����TY�� 3bE�ȓ
���QW�Vn��Ț�J���$c	<5e`�&�,:��Y��q�F¥�r��@�Ԭo�[V�&D�`����"���#��Y�u��Mc����G,��q����I�D��M0�CF�6���)ƀ����$B�8��aDd��~"�'`�,y�r�_(��Q�@"�y��;V�~=��N�.����U/H�̸'I���,F�$�آ~��*�� ��q�� H�RsJ�<�d�R�ݮ�d*Eخ>�z-��f���?���MƟ����<�8�
O�'����Hh<�V$�@�����
�0��@��.B�EB�����{ެ�n�1(��D��It��)���	2?���b�6	S>���)r����f�I�>Bs��`��!Z�b�?�~��`��#9*Q	�
O�I����/�&�C7-�}y�%�x�fJ0r{��C@Iu\x����2hq��liSěR�v٪�L�(v�v��"O�� "�^0c��8����X�~�j��-b��1����H���e��v��b�'�je92�=Q��yQ@֣����
�'َ� ڜ�D5d����ʀ.7��p��)Q@UA�C�)*�p���*�p<�f�'?VX�F+�G�Zء��Q_X���@�FHĴ�G#��~SY�gOY���BM�8�$c�bW9�������FI�.>�¥b�I5<U%����j�	�<T{E�ެ\�����	��,*���u��S���2��;(F!�D�I 6|� �HF����M�76$p� j�JR�ec�ϛ_���zg��>Y3�H8G���"$�"|O�,�Ā�`�<��L�$��x:�DV��D۰�=n��5J����s�4�cB_���<�ҋ�/J(&��ӫ@�x���"U��s����Q�LNl�(Pǉ��~���N�b�� �q�͂Dݪ=��Ih<���� f�H1cP-���8tNG�h���)ND�~���	J�0Ւ�Qe*�Z�P5���۲d!��	j|9���n����g��4^fJ���зC
~�*Ox�G��O:1;tO��[f���fI��\�X�"O$�$Y�#�+rA��f��7O�$;��Αb�t���2�j��^�6͊�hѲNa}���%�d�:l�Ie�y�m�W��$r!��M�&���Ө j(�"��	v!���d�`b7h�ca�R��Y
!�$J>�t#2Z(^~"	�t��{m!�E�}����$Ɩ<����֐\!�$+cLl��j��Z��	�Q�W�!�@�Ĕ\�V�p�xQ�O�S�!�ՂUE���eԺ3��h#e\��!��2ᡡI�)/<��(k�8$�!��JVԹ��U�e8�����!�D��r�^��&�6MP���ĕ�Z!��%���EC�,pNY�Ӫ/P!���	n6t�EP5��I��(�*)|!�Đ�`�����(�k��D��b3�!�D�5y���e&V ��Q�e/E�w3!��+��)��Q�p��� Μ�5 !��w�֭۶T76�*@�$��.!�ך7�4鱇�5iYl�Au�т'!��]f����
@"Iv�atAٻ>!�D�x�L!���xQN���Q�Z|!�$��}��+P�3!�(�F��Jv!��{ժ�V���J�yv!�dE�!.�R�� l�j�����|W!�d�m����ӕ{�HqZᆄ�r!�DC��q�3�7s8�9��k�fT!�$��TA�UР"{nр���%D!�D^]��X2׬S�`��Q� 
3;�!�<�B��G��  ��H�GD��!�D	�M�N`�B�1_��զQ5!�䍬H� =ۂ �z�����N��!�$��):�1`$OI�&e@�H�
�!�	7��hӡ�� T��[6�&u{!�dޥZZ��!���r�d���aR--t!�dA�+^i�r	' �y+w�(P�!�0�V�f��P6�ܣD(�KP"Oʸ�ª�*�,0�"#�����V"Oм)��pP*��oY }�h�Q"ODMY�(܂*J��=f���"O|���֜a����p| ^.tB��7C�� �E9�,��Ht�B�ɼt���@���*����	�C�I���Eٲ	��R॑�A<r$It"O�@v�Uga�U`�E��س�"OH�ǅ�9�\��>/�Bd[�"O�d�Չ�#z�BDa7"̀K+la�F"O a���G���R �&�Lۢ"O�d�7`��F��U����#"�vuS"O*`���R� HT�˶y_-:�"O� ��{6��#t�p���|NNm`�*O*��&�4d�ftSW��#W���I
�'��D��H�0K�\����'7�6ix�'�����I1�<��$�Bt��'@�&�`Y#�"��q�Ek	�'�ZU� MF�Fs���7&]�\���'�2�kf�ͨ*筁�B���y��/��D[B@"D�e���y�,��L�⡸0_
|@�|jP���y�K[ -�$�V��n�Ԥq&	��y�D�;k����KŹ���ҡ����yO;�TqRd&S��
vo���y�A�@b�ˤ�P-Ҕ���yͼ6�@J�ʚ�8ady���y�K3v��y( "����` �#�yDF&1��#��/kj�j����y�ӰƢ��S?!�jp�U���y�焲75���D�o+V�B�g<���Ϩeb}Z���3`��qFы:C��\@�L��	Ȥ�4��)�P� D�ص�φ"�Q�B�&,�mB��=D��q6�(7���@��Ǫz*R�2g�=D��j��x��6fA�2T�{ �;D��p�jA��j��ڬ)������.D�P(��Y�l�9B��09΀pg�*D�x2)ێ����#k'�0�'�-D��i��Ņ&��%Av��/r�(*?D��CQg��@^����	 �>D����!�� ���L}���0D�Ba�j��bV��%23��jU�0D��y a��.��YǣJj����D/D��3�σ�q3����D�V�(��F�'D�<S���iF���VH�zPqK1A;D� ���P���Hp��("6PA�&i;D�Ȫ3"�<H��-&�$qI�&D��ّ���}��
H�S`"I�ŏ$D�I��Y�:~��D�D�d,�XI��<D��X��uB2Q���A�E|��;D���"��/��������t}&��q�&D�h���-�FQ!U�)��k�!D�(Y�`�C]:��Pc�h��`�R D���F��l�9AT�^�'��Q�!=D���e���8y	�[����;PL9D���F�)^u�����^���SQ6D�ܪ���
9!F��*� �S(6D����w�:hk���v��	5D��ju�$c����K)=$P@�>D�@Ӣ�[D��D���_� ��<D�|!'d�+\� y(��Dr���2�0D��J# �`1�����e)�](.-D�p+�I�K�����+V�ܡ��>D����%�3`���K��	[^ڭ�3,;D�4I!EE'Z^q�W�
3l@fd��A7D����]45?�C�����X8�!;D�����O_N-bꆚ���,.D�ĉ��������34��8@%2D��IbK�t"ز6�NWc�y 1D�d!��$N1�8�c��$+� p�a0D�hr�M��tUdq an�!s�
x� �1D����!N���c� �z���*��.D�P	� _:�������H�t�"+ D� :7�Q%`3h-��F�?@E�U*O\�g�)}^z-�g�"sc���'"O6M��o ����2(�.�P�"O@ՙ��GN��Q:�� Uֶ���"O� T�C.�x�L���E�`lp�d"O�А#��2�]0�.��>>�#a"Ohp�NϽ4�]`� sX��r"Ob�`D��2R�~�w�)���qF"OJ}�"�_�pB:�%❽Y�Ơ��"O�����?I�>KBE.��(�d"O���	P�IЩ�b���T��58�"O��&�4��|k��i�"O4�+���:%���z�NA�Gc,|Pd"Oh��a�dz*����/3T�9f"Ol,��CH�96a�6!mR.�a"Ot�$�M$U�e��m��U�P�*"O���7#���&T��F-e~�"Q"O�y�i�'t?`�a��Q2v�A�"OZ�3��ʠ,^���/�z��D2c"O!�Q�}�J����Y�%��Xs`"O����K�)G�|!��B*M����"O���a�*��q$c"-�`CR"O�|s�aE�{�U���ߟQ�.��"O"�:��rBM��#�l۳"O� �#L >M�&���I�h?�i�"O�B�iф4>B ��	;'պ݉g"OPQ���I���zB�ˢL�xT��"O�ܘ�h�pK*���,��!��Y(G"ObsR
�=
������ѡ*v�`��"O�)v�U�	F�*�"]kp�3�"Or�9U�����u�3:4�f�'�!�$<^K��7����qag-]�a|2�|���:�PȀ�_�70p���Ĉ�y"��|X�I2���nHQc�*C��O��=�O.j�d��9p�6\��]1++n�i�'L����HP(Xwiϻ(b����)��<��nJ�*1�ǂ�J�$�8�MHu�<I�M��B��I1M�D��L�o�<�aA�#2�̸�6��2v*ă3A�e�<�$E׸&�(L�dA�F7���C�b�<�΋�Y�p �P��A�"��[�<)g��<$s �$M�(�p���q�<9�&�m�����C\s��dH`Hq�<Ap��2,�Mk&R�R�+���A�<�E�_N���V��$ɞT`��{�<ѥ��c�v��$-�79͹2��v�<��o9|dB�3^b�1���J�x~C�
:��Ro	��lA��H#0�LC䉃 (�"H�N��64f4C�	�x$�HB�EF�����6�B�I<@:��!�	%��lO:"�B�	�[��0	��
����CO��B�	(g܁i�!�v���KFC�:��%7EV?����р��`ÔC�ɤaz�I�f��Q��	KŜR!^C�	�)��<H���4)������݄C�I�.�`�HZw;�H-[,�fC�	:�ȡ@��/U�%�UZC�I1>�yӲ��HL��6哟K�C��.H�rԛ�E�5�Te����>��B�	>9B 	�� ��	����TIY��B�I,q^���W#�3P�^�GJ̨X��B�I=�0< �(�.C�D�Sk�5&)�B�	�!ݞq !j?r��5��H�g��B�IZ@P������(0��n~C�I>(���*v��T9����ϙ�2B䉅V�<t:�$M�[	Xm��O�\� B�I�'�X1B�#Tq":�Hv�N*�B�)� �yy`O�1iO�� H�kvB�c��I���I��|T��BFI��o]FрQ�H�Q�!��a~��R��N���H�$����0l����=�g}�'#���X�a�NɄ�#f�� �y2o�00�tas��3��P�n��M��R8l=����d���	�:�tXq�V�j��z`�<�.O�P3C�F��B��aN�=�
=�'�lHH�IC�_�e�"[��L��{���r��b�����@�OR�
�J`�K�H��@s�"Oh�:V�'��*M5��e*�Oر�M�J>��1�gyBO�?d<t��H� �zT�\(�yB�2���Rd�@(G��0)��A~�n)�
�'�~���A�C�6]D.�*5&H��ո'��(��b��jU�c�ٗ&J���'��	dJ�6n�����J����'^�	��$�X�a�E�s����'���6kA�d�6�34��pq��'���%�*j@]��ӛz�x�
�'�&|3�� {3���fc`B��
�'�^�"V�q�6����H�]�-�'Gr���Z4�b�����[��,��`�L2s��l��z��'~{l�ȓ0e�x�E%ƃf���
��5�~��ȓS�����[+D�	��ؠ R�مȓ�\S@�Q��Xݠ7b�%�2x�ȓl,аf!L�0�(��웙92��ȓ\�9�@G< ��3!��	f�(�����p�K��&��5�9]3Y�ȓҒAz��S�5�P҅,�5$,�ńȓ-�� ;g��B4���O0���'�J�K��^4S9���)��A��.rTŁ�^(r��w)X#zmhx�ȓ�+� ޹2ĕ�3��,R�͇�Uę3��	�
����L0�i��t���0�)!
*:��������ȓ4f�u�C,5��`�F�;.(��9t\��&J��P�H�FD��ȓqC�9{��R)�4}�
�<e�29�ȓk��8p0�ӵOy2�k���l
���ȓ9��M���;Fł!���~��0�ȓe��օK6�P+#�S�/�-��9J��bP��k��J�䩆ȓe$�(;r�S�[���h�a�ȓe��TIg�5;[V��U��z���ȓfPj��*r��@�D�],n���,���"�Q37+��q�+�<��ȓ)�Z��e���F�=vr�؄�SjZ�)�.�<i��A)�Θ�_�Va�ȓK��mb5ν;V��{b�/^|a�ȓ0���3�J\�>aX��EU�t���ȓ:����4 gͼ%+q�H�de�8�ȓpB�i��"����ʤj�@��wl��'	?{~-x�g�h�̉��c����ɟ�=w.��4G�bd9�ȓZ 9���e�L���2�"E��PI*� $��nŲ=���Oc���-��13�v�zfc�:<�ȓ?8R��0�.]b���� �%V^\�ȓ5D�)2�2C�$�3�0}߮���g�L���'����}XDO�. iF �ȓ<V2��dɭ5��#��*޼�ȓn���`vo;NjXBB�-��-��9*�2&#Z9���ժ�4��0�ȓ>�h��F/;TI��22�`���S�? <�!�+@�^���q���>�zy�"O�qA�U;5���Ja��1W���� "O�"egŗX�l���n��bZ<�т"O+�L�@!p���K�P��"O�DA0 �� ���zQ��'٦�Z""O��%�,dj��Ώ�QҦ�u"Od�I
���Zmd��&1�� �"O�ta���yh��fėt��E!f"OL��@��*��L�U�F2m�v]e"O8�`H�p��B�>W�P�3"O�P��OԆ��wK*rX 2�"O���OѿAgEDА*p�y�q"O\ a��_k�=��c��0\�A��"O���J�u�<%�@�1Y3
�2&"O^�ӆ͐���	Kd�[�f�K"O�k')�-X�e��,л3�N�2c"O�#R��rhR�eL��"��"O�y3�*T�O������G��T(�"O�T06�\��qf�;�Tl��"O6�8 �Bat���$�(j{�@yT"O`�#��ZcTv-"�ͩ	�8l9"Ob\��L�9"z�
��A�(٨�"O.���  �   ?   Ĵ���	��Z�wH��:X���C���NNT�D��e�2Tx��ƕ	#��4"�V���ą�aV�mZ!�����2L��Qa��u����45�����lۤ�M�a�!<3�NZ�Y��@k�m�5����I͟���.I$?��T�r�N#'R�q��N�a�P*R\��jeR*2��KJ�(p�L�9��e�E�#h��f�
0?F85a��H3<�IePn�Qt�F.;�ʓg�y`����:��'L��۱��%�����PM�\��$׍h|ɋ��.}"�N�s�X#m=}�&��0$R�Θ�;ۊ{��	 x�&M�E��	d	&�ְ��&�V��MQ���ۓM^�]���- i8P&��~B��E�xY���*}��e�A�JEy�L�h���g�.|��@!�2L����@8b�(�J�p��M\xl���S��\����j,�J�[��1��N<^�d4�`Qp��
�h�ƹ���b���.��������yr�����j�$R����)���?����
f�l9&��jq��n�V�O��k�(
4Rf xd��;L�� ���G�l�0�a &}Āg��=��'.���;B��.KO�H`!B=Z�"��T.�L�x}3@`Ĝ��$S��+&�����������K8��߂�� �&fQ�do�>���2�-3t	a"��<���#�B�(3�O�	o�1�&̡g��q�����{Q�)�R�h�<Iƙ9I�6�s�>���̊V�D̓t�a� G�.���X&eOk!T��',�Ahk�4��6^�bj�r��!<�:��� Yj(<���@�2Wll�D#Či�'�6U+Q#Ɗ��A��ZV"�g~��C̜�}�,T�Q��4~���[��@�4�sG/C�8�);��I��́>� D���{���C޴�x���!�x4���0��'����!H����D���o�2T��Ч��p�ȴa��y����giFu��O(��2�H�R�y�N�[UEb��I/Aw����$�<u� �g"O���
�  �X�3��O���O����غ����?��O����D�I+G\,A�,	�\!���&#E}��{�f��Xx�V%�<WW�d�G!Ec�'S������H^��d�F�-�v��syh`���| ,��#�ܒWҖ�a�6'�1��yr��?�T��	�SWD 9�Nڔj�Z���.��~"��@����¯H���a F���yb�^�&'S�N�$�T�����7ϸ'U�6�5��X=C�4mZ�o�6���Z`��7#E@q�$ۃ0�)p���?�Cے�?Y���a�,O1l�Y�"��©��A�_=�UA�!Ǌn�����*"�����+Gr�R5E�\�T�PőW���9ۛq�PԲ�P@!��⇮�G�'hέs�"�LF�[&#���&�J3�"<zd��s�����{�:IzC�x��\��s p����/Z�D�C�T�T=�T������zf\�!��iu��'j�ӻf�z�m�bk�,VΔ5B�-kW%ɓr��az���?�T�ݩDUN�Yt4U
x�k&���~b��?("���ƃ�9�8\��jP^�I�\"q��X�,�^�p��}�Oڜ�ʶm��|x40v�В��M�M<Q �
��DH>�~� 0��暇l�hYxWiG�,�Z�"Ou����|�:�Tg���y�6�'��<ɇ�w8}9'(V�hd��ʃ�k�B7M�Ov���Oz\Ж��6�f��O
���O��G}{JŻ�P���`kG?P���L<)fGۗ~�t��|&�\�&ԟ7�����<�l��۽��P^��ʒfK����ēUZ��U��+'?6��Þ����Z5�7�$�����L<��¼Qhf���+�19�>��Lg�<A��8.���H�jI|�)�B�w���o�����x�O�Y��8�L�|�
���+�i��@�c�^���D�O����O򘬻�?�����4�V��%����6C�H���LD�,4�+PX/�<J�J�7�$4I7�I:q� ��d
�I�h����Fu�1r���mox���!B�k����x�'��ɢ-X39(9�&OA.y�At���?Q��?������1D���)㏋+ҬI�װ-{!�$�&Sg��ȇ&�bX�e�
?hCqORmZ�� �'!B��~
ݴ1��R��\�"��PUc�\a��h��'��dœS9��'󉖃"��8t��vZdi��ҰP����"�T�T�b�(l�u�����"�z>�����0�hx�^.<�Ԙ��U�J�(8i#��E�����Ñ�MK��֙�O��:��'&"[������z�� �Q7Z�%�v*"�I�X��+@�T�c��V�!�0�A�C\%:oB����l��[��h}��e4������'kbZ@@R{������K;KR,7�RY�1ZZ� 
�(BB��>Ъ��	���C3��H�q� /��i7��"3����i�~�R�&1Y\ŀ�L�9�}˛h�I
 N�p��.A��'$A�!dXY�}J3�D�	�R� �I�f�����_�I/$����Ov�}2�4]�ő������8c�#a��a��O���u�L>p�\I㏓�e!��2��'>�<�1�Ɖ%[ �8�,_xTPrg��_j6-�O����O�|+���.F����O~���O7I̆ua�j� )�0$i
<�&b�,r��&,OR� E�@,3�"�!4�S'g�<����$�99ay�(���4�Z�j���&��	r��%��&L�Oq��'�H����M"E��q$_�f�����'�!�sȈ�&3Ȍ6��mzI�x؊�4��O��b�.�
[��FU�(g�;}��KA����ʟ��	��u��'}�4��H����>tŌ@�Ч�1q�^�@ D0/��3�
�+(�Z�I�>4~�����%�(O��K��4Ew���(�=s��h�S�rA.A#�� U�hz�)�� ö�(T��/�(O��26&ҩ'�h�X���$;6��Pf�	ce2�$�O&8QGŏ&a�P���L:_�:�"O(8W�P?tt��a�Xޤ5z����Ӧ1&� #)�&�M3���M���m��i��j�����5�).
�'^��'��6���d�
R9��*ò�,�g
�-X��b+ˋj6��ΝC��X1����(O��"-ːzY�Y�#�w�4X��%
�%���b�
_�@-&��%+hhQ�Hb=�<���$�l���~d }�ҟf.A��$$b!��D~0���#T��Ѩ�#ς#���d�?ʂ(R�Ĝ5Z!nd��K� �p`0�(�ރC�n`n�ҟ|��]�D��cK��CZ>
+$E[ )��}����$8��D�O��$��=r�Yh��բ8E*�#���J�:|r�*�~��b�i�h��<Ld��!cC�r�ɪO� ��@$J�\ZZtCB�S��$�B�
l�Ei���1��P�b�`@�N x��\�P5�d��@���&���/h����Uq�I�7%��!�Y`X	`��H�D8)@C���x�o&ʓh�r�ACc^�R���O�X�d�>)��?��M4�6����?����?��tV��'c-.9�<%�������O�}^NQ��eŨe�U9��
,���D�z�Or�(�hҐ9���`%�x�hU���Z�B�©��	C1;5XPV��)O�m!�<�4�ֶ36��}:F���������P�(��&��M��i��	+JM��,O�6M�e�~��� ь1�6�aj�!
V�E{��I�i3J��v�tPq�SHq��'&6Mߦ	$� ���?��'t5x0�X�w|�a���/͒��f�<���g�O��D�ON�$⺃���?Q�O.�`�K�R�5ҕ�,�IQ^ц�X'ڷo��P�#��~��uA���Q�'��\��Aѧ,:d9���Ug~|�C�>rtE�!c��K1��y���P��ԁ�/\$q��y��Fm
D8q��i��=��O$R.A��Q�~�ŐĎ�
�@Ո*ӆ��cNW�yB!&x�1)BGצ-�P�b����'פ6�!�d�&-��T>�H��_�Viە���4`l9�.'�	Z؞$p��?-~Š� ?e�	��*%D���$�K�6�0����tIXI�'-8D��r�ˏ�[Y��2���WN��%�2D�� ڭ��XF�
`�p���JC`�P�"O4�z���/PW�R�E��)�@eå"Od�)�hN@���w�ԬfӢ��q"O�U),X�dZ� �J�i�����"O�\ئM�!v ����9��Ę�"O��aE�V=���K��̅-\2��"O��Ӡ��׸��UC�K����"O��B`��~ȁ�0e�T��(+�"O(��$ѻl��͊�c�����&"OP�ԧ��9:d�P+u�u[#"O(A�C�Ǎ\�)�@� 7�@�"O�|@�ꇇzU��@ĖP=(�p�"O0��C,8�Ąp��G-U�b}i�"O4UQc�FhA��Swz8�"O.�ѢԻ��1b-��zX��P"O��YPK�%ג���+F.�,"OzEag!��=^�2��:�9"O|��W��̤J5�Uv�Ѻ�"O6��7I΋����W	ݛs�4ً"O�1�(��'g�M���@�炡p�"O�T#∓*L��law���!���؁"O���a��4=���<|�`��"On�z��ZPyC��\/9�2"O�1���t���s㈼fXH��"O����F������N�q'؜*�"O.�w���.;�u�S�ȧ`�M�"O�`I��I&�Q�]���:!"OJ���×(z�[��͖b�����"OΩ�,[��B3͌^~��z@.TR�<�%K��8�ˌ�N�&4{NNe�<a��0����FF��uz�fa�<!��wnyf��u��8VƂZ�<���47�"m�`N� 0�ȃ*�k�<AQ_�,F4�JW�]������A�<��@C�u�����
) �0! \h�<��ʢxV�y�U�E��-�q��e�<�L�7g蠻��H�+sbDѵ��Z�<���#{�
hٴ�c�n�3��X�<.�q	
� $k �^V=C��\�<��̥A�����
xx�Aԍ�_�<	�FC7d�Ys0�vQ!X�<1� (v"����{�ДkB�@V�<)��ЯHVz��T��x�x��CO�<�C�56]��`1@�^����7IH�<��ڗf8�A�oWm+�,г��_�<y���/}���ȍ
�(��R͋w�<��(|�,�����Q`�����r�<ac�=`.Tuz�A5�`a��k�b�<�g&�"�bX�w�^y��!�W�<C*\:E?@�pSNJ�*��a"V)�J�<y�掟Q7~��-� Z�fm�A�ZH�<C	S VG�(cj;uL4d@��C�<�Q#�?Z#��;6��1Xhts�'�@�<q��+`T,H�i);?�4�Uz�<��FM�-"Y�P�L��jyf�V\�<�� t{*�"-�:Ӹ$�K�V�<q��ޛW<F�ڕe?�Z9�Q��l�<	��I{�b =Lv�uÈo�<�Rʈ'T䁷�݄<�ݳcjQm�<9��@��̐bO��V�C��t�<�HޔnB��`K7]@͊�N�h�<q�& 0�X��L�0he�QJRH�h�<1��@$����J�|b��z�I�~�<�Q��-�&r#ï3�DL��k�z�<� �0QG�ޫ]���j'�C�*n�=�"O<��o�#�D����`G�M�s"O��Pb�_�V��[7g�&G�tcp"O�C�M�['�H椉�!C�	�"O�P�+��wO��{ ��Y[h��`"O�ԂG���WN��˓h1g��@�"O��q4�d�J���r��ڑ"O~��c�Q�j�!zR%�+^n�y$"O�����ISZQ�#�X����"O&ɈG�T�60y�W�!r���c�"O��'�|+x́Q���4�n(��"O���g��3L�A������s�"O���2�����)�͉�?��ib�"O��Z6L 8	���g����"O����d��2 $�r��ܝ%�~x:G"O���3�h��]����j��U��"O�5SĎ�*�Vi����z���"O\�lʔoD���k[0��S�"O8<c@Uzq�D:�Iӫ����"O"��á-� V�P.��ػv"O��3�h�/Ux��Ԥ-�p�)t"O.{�M]?PU,``D���}���r"Oh� Q��)�2�;��ډX�:y�W"OF@�$/���lH�-ȶ�(�v"O� �5nK�'���;�ˈ#�"���"OL��R'�E�"$�Ǌ�9�Ty�"O���"���(B�aBk� =���#�"O&L���_�"�(��q��$ywFM��"O�!b�c	4 3P8PuI��Yu���"O89�n��P�.�,\�)�"O�}Z#���W �E���cY�S"O\��*�̰�O	'K3��*q"O=bJ]>�Yi���$P����%"O�L�⓷0h�e;�U<^�&="�"Op��撪%!���S��,(
���"O(3�T�n�0QGL{؍`e"OЩQd��J�&{�c�Lg�Q��"O0K A�<t���|b�TÇ"OF�)v��;0�� ���/M=8E;R"O�yD]�g���C���l�
��"O$�j�)ݛ���F�A�6 ����"O��A��,e�>�beeN�nk�(�"O� +��O&��#�5If�K""O$% 4�ѡ9�d PBB�:b���d"O(���Q�9f�p�l�,���"O��ĪP#+�����pt�LC"O!�v��/�L��#�CU�1�r"O�U���t�����y�D���"Odq�I V�7Kׅ\�f,��"O�0�"T$a�Z���_��5"O1�,A.���1�jA"OxY37�� 2� :S`�D�B�r�"On<��枯Z���s���?��mCF"OvT��M�{�	 �"ʅ��b�"O,���!O�C�D*t���!��ɕ"O��H��[�i��1{ǯɘI)��"O@x����%o�٨�P�=	d�CB"O�8��L3y<�&c���4%Z�"O���d�ԿGC��!w�ӧD��\�"O,Eto]�X�T)� Xl�iQ�"O�Y8U��t�=�a���w*�=*P"O���CL@�fD���/^5$�`L�s"O�P��7/ڀR�&Lt���"Oȍ��AM&c�&�HB�ީY����"O� �Lj�J�^����݁;ʜ�"OZ�k$ ^l�,#�S4�;�"O�p薯/)���rM0D肀;�"O̍�f��GO��Q�f��ni����"O�@#�	�I������Y�z2�dHr"O4i�H����C�kϤ.���:�"O�����ݗ6��8���;�v1��"O�� ���<�Z�)��t��	�"O���é�@d	�F/L����"O:�� �5��8C#nJ�1�D��"O�Vk�	G p�cL�l˔��"Oz)�ݲW�I+V�Ĕ5��'�J|k!k�_Ɣi�+щ\�L�p�'�ޤS����*_� #fg��%��'Qd�r�%A��z��ү�T��'�.���@Q�!�h�ab�֧քB�'�-��c
���1��¡��љ�'��0�&�ø�	i�\�(���'�2��"hҍ7�vQ���x�����'1�M��>����̕=oJp�x�'����>���q �� ���
�'܆!
�$<������5�
�'�H�Z��\�M6�u�W�vh,,��'U~�iQ�\kJ¼9`nԘub^���'�0���CTxB�80	�9_�⨨�'��z�V ���'�7L{jI�
�'0�)�� 0T���H�G��B
�'e�M���(5פ�B�ƬCh4�
�'ht� f�'4�Ab�8F0���'���`g�JfY�\��jѱ�L ;�'m��1!��p�Z��D�= [<EA�'
l+p��i#�E��h���u��'WnD0⦃,���k�(i�1��'����Ŝ$tz ia�Eft�!�'�.�X���/n;D��� ���i�
�'a0 (�菌"�@�a� X&W�0l+�'>Y@ ���ԬS�ɖ�b����'��ɋWP5���l�>]����'cR��!�HuJ�Ap�G��,�
�'������u��ƴ;��r�'�j�P���&膜��E�-V��h
�'�lX��`��2	D5g�Z�2O�T��'�iҖ��pU�t�E�)X��
�'�J�Q�gH�n�z����4�!
�'��Yy!L��y)T�j���\�R}�
�'Z��У�/C��x
ԅ�Y��a
�'��E�������M �*7�'D�X����W��BG��/:3@���$D����#	�R�	T81��Ɋ�o�C!�D+L~4@3���#&���/��!�$Ǳ/���q��\�J\��̈/�!�A�8V�d���N	K�%D�!�$_� �|��=�@!��E8�!��&x,���C�`����T.!��+-�� Y�G�8t���0$J\�<!�d�_`J�d	�?48�n 8!�\�t��+��\+a8~d!]?D!��ҥcM-�PA$3�.��C��ȓ7��q�ڝo����,�nq|\�ȓX ֕���M!v�>�y�ş�^��6"�yqB�%.�� �Ud��|�ȓFf,y6����}��Lڨ~����ȓ_/~ ��F�{u������4u����q24Q�g�I��6�*kZ$�y��S�? -3��>V �yPd40U�L��"O�C�\7���ND��~ CB�'D���ȧ?�k��/>XŻ�V�,_�y"B�ˡOR���SpL;��շ:�|I��ڣld$��e.�CѬȟ(�Z��P�	Ա��S�Xik�fД��P�O�V��ȓ_)�\Y6�۹SX�����/�ć�
��y��$���ԧ/ww1���l�� ȓ:�ɐ�Y P�ȓg����*9aN�L�V��������9��FԞ'l M�@���l��UY�+7�ħ|�J����I7vW�̄ʓ9"`kEd�C�2�	F' \`B��Z=�6C�w�д+@��U�C䉷Z
��H,}\��S�Kݻ(���D�:V�Zp��>H���� �U.�!�$Q�_ �$b�5��p�!���#z.(��p�.WL����I�/�!�d�g�L�iU�èYOD$8&��7�!�D�ZQ""�!,�	{C%���!�$��U�D��7�K�V~]�k�6,�!�D�<j�~�:臑w���Т镂S���P	�c�Y�O���J�K  X�$/�|.��	�'�(��X�%�R�� �B�=X��+�'x��XV&E�M�ɧ�� DpQh�:9��V ��(e���"O��h��q�({���V^5{0Z�p�GLɓ�� ���c8���p!H���KA�0��+c�7�O|�YS��\�6�� Vo�Q!�� �Ãm�,p�`B�ɽfiԡ(Vl�5��4�/ȹ �\#<9��;MҩAU��i��kN~J�h�_�1��t�,9 �|�<-�H���/վg��q�.�\;��/�H���'Ş'�s�&�5�?E��'���炞`	|]��
ھ+�ґ��'��XRO�/{dp&�٘4T�BS�iJ���m�,C�8�����ʣ?��'��^��9!zg�í^}����	�7�:���Z������O�4���
!c.TS��Z�j+p��O�~�K��? M0���"��Un��>�'b��<���&I/~ 5È�\9�����
I�J�aC�ev�C�f�FASd��D ��*x��t@��)#�(0��Z$ K���`�>�Ov���Řg!�����8�Y�ȓ![�Mh��x�X��͎}ܒ�l��i� L:D(X�Ե۵�'W���֋�� ?2�`DPW�!ۓYH��bD��)3��zadџ)������C�%8�^X [��{Vd�CN˵�p%�����P�>)$R�j�DZ�imWf���������p�{�ń}�8�	�HˌR��C�Ɉe(�H��
A�=ԌS���r�Z�J�4|.���K�e�!�%g>�g?����>T� �9��W��˃OR�<A��6��J��+d��¦�G0$��p�e�Z�d�,�@��^,
z�3�@T���&��k7R���XBLz݆�LD2`��F N�V��cH܍%�T<#,A".��4P7�T�{�܆�Ɇ;B�ڄ@V�Ca�92lF�QB@#<�0B�M�v�����lqJ~j�ǈ�#r�{�eK0�j�� +:T��B��ڹ`#���w�h�0��#x|���ڙ ����f7-��)��͸�Ø�q��0 ���g�J|00$,D�T�č�*#�
Y���ML@�1�<)`a̋g�40��p8�� G+�8�rѹ"��^�B�gC9�Oԉ��$A"d��O�uM�\�C`6+΀`��-Z&�|�Y���D�`�� �i�"eG~��:	&#5d�[�FQ)ԉ����O�H�4����5�B�nd�4[V �
�����Ǔ6;L��T"P�/��`��.*�aҭ�?�LLsW�2#���`��S,'��a��[<b����a��$W�!2�t�8J|b(9���W�L�W�ۏ0��C�.�Ƙ�q��nl��ե�|鳢n��=7����
z�7��OP��FS !+��4h�̠�B�Z2H������:,"Q�P�����N_,�AnZ�ed�K��	�x��h���&hz�#?���޾R*l�0J6�~XgGs��x'��Q,�����<<�v� *�Doǃ"�-3�O�5��Ŋ���(a��<���!x��S�+��p��S�
d��c���Q �D���O�!U���)�oӉO,�u���	�p�,�#����Bk ��	�'(ZԺ7��.&�h�I`�Q�O6<!���M�[���cP��$�����4DP>��O��2 L�>!����$`�,5�=H�"O��&d]L0�ERC����q�i��
�ή(�h#�ը΀}8����/� ��i?�M��KF1l az2���?��U�'�&0�0}�j/Z����*B��6=F-���S�#�O2���-P|F�ҕ��L2��
����lr.��$K����@�c?}I�N|Z`e��S-|��!��[�����^�<�#�q@t��*��#b�j�%�2pMeL�b�; �V���"��QF}BO@?1w��*P�J��|{�. ��y2��Q���k�7`#$L�Fn��M�3�X���m�h��	�H��Tk�w�'�`�Y@�݃b��+@k�1j�|��~����<�ă/ĒJ�1+��Z�&��D��O@lq�(����r�a�H�y�xp�CO1���D.[���'��F*S��9p��g{t$�t��bf��a�ڰG�=)ǆ�1 &�B䉣L�f� ��H+`,��.ߴr�*8�Vl2���΢8�r7-PU�O�J�l��!JQ(X��u�A�Y�Hp ��7X$��O(�����!=�Fmn��v��%�?t�2�#۸m^�"?��M�#= &kf~"���BM��4���QMY`�ζN�ؔd�52�����E� ,L@��@�m	�X"	�cT}a�E'?��R��<7��!�<Q��,� !�2B�&��t������ �F�{��ŨC	�y��|��"O���Bb-x��E�CfV�"��ѢW��d�у��V�$�U*P�i�
"|�D_���ud�,<!��B�!K���i�� D�
@�Ka*�����!9X���p�{��}H H�%U��9&�Q[np
��9M%��Ԭ�=d���
�+p���Ė'f�R��({�Li+c@A�.�(X�MH�9r8�KUTY�D�n�R؟h᧌�#Z�b<x�"$z�d��#D����D�6���s�	:���&�<D���r�<,z,�y��2{��RP�6D�D ��;XX��g�Tܵ �4D��Q�f9/��tgc��4�d�i��&�I:>2굆剴=J��vnԑ^�R����N��䔔}��U���K�� JV�$�dU{��N�j����i��Y���		���"w�\�TQ�`�� ���������z�h��g�t&ق�F	�yB��y�p�K�b�A#��s�`��~��L�W[6	��-��Sg��8��K=q�iY�٢B�2C�IJ�6`Itg�7cl�ӳ�¸=�˓�ލ��G�2Jc���D��l�z�kA�҂bN�IJ͜|�a~�n^�9��d�G�\ �A�
�_��؃s%˦u;C�	5s�\���*#��py���_�#>�bF��}��@a�'o�Z.�"��'��q�H�#�D�E��)ҥ"O�s�@X<U��s&Bľ3�� ��in���>0ND��۴o� $x���i`���$KJ�6��˅)u�F5��'�r`�U��(&���֮>�p�B!&E�i�j�~h��C��鉿j�hs���2)�0�����PT�����7?�BPC�J%}4� P�C�p|̹Ì�7t�ޑ�F� �����7�O��cナ
btò̏Qֆ��F��,.T��g듪J�t��ğ0V���O�D%���\3����E�e�z�4D���Q�Z��1�U���58c�l�]����e���HiY��QFN��ҍ��w�b�;q���w]
�X�+�%3����'%��+�k���E����5��cRj��=� Y�&O��.�SG���4�I�n�D���J'3#Be�cG��C� ��Ğ!�@��%�� L�r/!ya�L���dE \x�kwr��@SL����C�Ji�4�G"f,,Dzbi�i�Hu`�)�"A%�E�Ыq�$�@��!�Ã+�Ьa���y����i|r��V
M�^�-�@�6�?��/G-%�ջ��N�~`1��iZ<�&If�7,�@@y�&�:s^�B��O���sl�J��Lq��֎r;D�i�O�ѩ���4G(h�*�K�|Fy2�@�-0���lM:�q� �ڛ�p?��n�4CA-���,A�`\�$Q1%�>dsW��Y?���S�? �}�D�؎:�t����D*l�]����7
���'FW9JoH�$>�X�.�;'O�d�%*�3�P#f�#D����&�"U�,"���h����k�<���_�pN>E�$�&9� ��g����	GV��y�
n��3��G4g䖜JC�L���'�N�#F�'�Q��a��4���8��/e�ȓ���&d��i�v�� ^T<�ȓ+8>��C�T
5�t�".�*����ȓY �j'L�.�� cF�>�̈����I�b�%0r�9�邰1��d��D�Ĉ��mK	�� 	�hOJf���<z]�"�÷^���ṙ�O�0ͅȓa�LY��HS<к�(Ȃu/y��]���Ɍ�! ~ˢ�ӟ}Ʉȓa ⱊ�Oy�@P�J�6����h5̱JFBO��i��
�*�0��ȓi���z5�ě,���)I�<A�p���V��S��Ԃ!H���"E��%�ȓiD�SP	�1��	Y�G)9lԜ��b���Xw<��@
�/2�`���7s�tY�ǅ�"�x�ң³ �tX��F��ْ����,��W�Ë+Jxd�ȓZ�Pc���{ "@pr���ȓ\<P�P���H�,����ʣb���c�yXW�ѕ��d]�a&"O��F�>pټ�SaKD`�("O�M���9=^=��gG&�N�x0"O,lX�I�1�Zڇ�"_�����"O��2�"�*0Q(	�eX�j��h"O�x� ��{�&U҃D׀)��5c�"OM�v'��vl�ҡ,ґ1�)w"O:A��� ��lÔ��nL�Pv"O(� 5���'�(5��B�q
@�3"O�8� �<?@x���M3~:hE"O��'*ۃ7� 9I�DEF��"O�U�2�% ��Y�����V"O��0!d֫w�V�!K�D��b"O�!�U�)\3V�ۗ`S7҈��"ON�4���{cL��v�!�ȬK�"O؈1��'-Qf@���=��5"O��2TH��&�{5��&T��9&"O�|ȗ<�8��C@�`��@�"O��"��>���`5E�9��"O����m�H<D�qnF<;���"O�h�1<p�tÓ/Q(:�;"OB�!���(-;��Y�n�Q�v"O4A���Y�(��*6���Q��P5"OX�o�{�V��������"OL����I�䰒"Q�Z���R�"O�h��.ͻ�l�P�G�R��5�$"Ovhh�B	��!d�� @7"O̸�cd_6s�8�&Mar P�"O�͑���b�9�c��؆"O��3+L�x��'�|%�"O�hz���Ŋx�wF�1�"O��*�F0bgF������,��ܳ�"O0�6�9%D4���s�=�"O��W�i�֍�r�.F�˔"O m�CoʉE��pX�y��A�"O:`;�jV�&fr� �n@���dx�"O)xu,B�TlLqG�%y���b"O5c�� �����?u4� "O$9;7�Wi��)�I@�Q�T@��"O�T��+ūf0Qa&��5R����"O� 6�f-���UB�<L��r�"Ovt ��ǥnM4�Q��f7���"O�E3��C4]���ױI�̡"O����Z2gLyJ!(����"O������D�B@)�bN@����"O�fV��-��C^ �͸G�'(��UH6gsn����
��\��ӑ[���1r珮fx�ȓK�ڀCV`~!c��V�|��~�<I�"�=���qa�o��Y
ƆCE�<�C��5�T��E�(4�$��\�<q����ƅJ�U�XH���'a�S�<	3�
t$$��$l�s���BkPt�<�@��	u�Q�t���
煈j�<A�GU�N�@���
�$����k�<��Iy��b���<��ԯQd�<����H�p���	��� Mc�<	��B��Jr�O�(>̔B��]�<!�m�P��T� B@V]�<�� ( �����I�&T�I#_C�<�bˊdŪDr)ҝM����l�B�<�$����6K�U��$Q���{�<i�$��o��:�h� D.р%IN\�<ib��m��T7�_���YX�g�X�<��i�9�ε�,���hH7dY�<Ab��#w���� W3Sp޼�S�<yg��pR����P��2!�M�<��N�S q�BU���P��V@�<)qk8cYЈE䓁��X
fF�Q�<��j"5D�-��/)b�D�B�)�J�<q,�:?��Ђ�f1zV�Ƣ�P�<	��0h��u���]�2��Ѳ�
r�< cW@^���ٟ, �bvG�k�<�c\�@V#�Xш`�A�<��bͨ$�x����A�=���F��}�<��lҔn�� %C� �l\ �Ty�<�Q�G*E��I��ȌM���t�<��ω}�Ab�	F�1�b8�k�s�<Q���5dMpCA��j��aj�^s�<!ШN�W6��wIVx���Ae.Yp�<�s�ʞ#W^�P%(�<P��I�Ai�<i�����[@��D@���-�f�<I��]4j�фg�y��`Y�ld�<aᅬk����Q�N�8��r�b�<AŅ��kV�u;�N��V�����k�s�<Aj�>`5b�AL��3�,�#Ҏ�m�<�b�ݺ49��X�&V{��=�D��d�<IR�B 7f�\��a;M� �D�v�<y�Yy������e�Be��g�<�#�Ɍ
���@����2 @w��c�<�2
��� ��vg��j�K%��f�<����?rJ� w��L����a�<Aa+�a�<\i�g��V�BXb`̈́W�<�U�Ύ6��8	�n�y�p�a��[�<O@�y�xm�r!��WD�d,�}�<�M�3p�*aF�-?�
�i�<�� _�^(�AKU��:��})���S�<�#�^1&p�/:PV��0��d�<a�`ێ
"֠�bW����D�^�<��� s���ʧ[&��3�.�`�<yt�%T�=G��	v���u�
W�<�"k�+w�,����+0��H����N�<I���.{�����D��	*WLEs�<a�_/wk<}�%���(}x��U
r�<��ab[s|0�d��S�j(ӑ��q�<� �p2�/��I���J���"O>(����z ;���gc�4�"O�钅��.CO��!�7?��xw"Ol�H$��/�:���%p��Re"Oް�)����s�Ŗ�;�u��"O�ԙ���';�"C��	����@"O4�s������b���X}*}C�"O�Y2��Q�Fr�1��� {(��"ON���cx�(�G�N{va	�"OX�+�i��-4���A�|��CE"O�<����y��ꅤl��D�Q"O�퀤 D� �fɹu*Ӛ{Ҝy�"OXֈ��~�a�	*�NR�"O�T���B�M{3�V�Q�.��"O<EЕʛ�J~8iBD��!p����7"O�}�SÜL7�Uz�5^�*�"O~� #j͇�.A���)[�ȜBF"OȽ�E*��dt(^�S`���"OrT�D����0��럗r;	W"O$uU�O:�6 �6h��l9D"O"�±+'7�8�Se_E�蠥"O$�j1�0X���E͖+�0"O�����V�b\�X�nD���r$"O�U�Ƅk���e�A[�0�"OjX��,�,5��`���zx:�z5"OJ�t��kA��X�}�(P"O��"!�K���c��^�t�4["O��y6��=C,���1��w]>P1t"O(�h���Mm>EH���6MX�"O0C�I�QD�ly!��Y?���"OЁ(���h�E�a @@�53�"O\��A� �}SnX�T��  "օ��"O"paÃխcO�	[��� {��0$"O���HI`p�3r,\�c]��r�"O� #1��%V�|��E�L6~�J�"O~̱%f�B���2�
3 ����"Ohp���5��혖�X�W>i��"O���]Y��c�ރ4�0�"O�`�ѥ
�j�V�
�_)�!�D�*o��l��ڃgp�%낹Y��B�	Ѫ��t헝#�t�!�5Gh�B�	�	�٣�BK#�����'T�[�B䉘A2h!��S�~@t�rEABrjB�	�C��%3�)Y� �d��[�>fB�ID�D)*ũ
*�>��@�9>jB�		"N�G�X�5�����5�B䉢K�� �q��;����ɾ!�hB�ɮ.=���_Yڠ�p�G?Z0B�	n�nU���
(��U��Ē\�B� D-���B!ǕP��DR��D�5� B�	�N+x�۵�J�zX��h��C䉹Hzaq����>H�ӢA%V}�C�ɷ>�5�Co�% r� 0��P`�B��6/Xp��˟�h�� &#��t�B��A����Ӌ?��sBc�8g��C�I�2b��`���C���r�5q��B�Ɍ(��x�a�Ilt� �e��G-�B�	:[�r��*W7?���%��_�NC�I��^�K-({�1����}lB䉂wfq�D܍���K1��3	:B���ۧ��3�Hѐ�h�F8r��#�,D���Rg�=�d�Y�BP3B���� D��3�BI�H:b�jB��i�(���$D�d!歙25xI�����ڢ+ D�� �i�4��!Z����nfN}�#"OιJuk��W��dP�6Up��d"O%!f��;Ӏ�:���u5�p[�"O��Ҳ�Q��<(�bU��ܜB"O>��wG[�.����#C3�`��"O��.N�9�P��ca͟,5��"O�l���ff�9r��M��` a"O^��#�ܧCa|C� �/��{�"O(�C%߃J�f��O�
�|���"O�t�E�Q�9M2E(g/ � �v�p�"O�<YƥN!+
p�c1eKl�܈�B"Oh
��-h?VY���Yæ�:�"O�-cDһG$�L�6.���Z�b�"O�t{WI3R�#�0~��#�"Op�a��_�_�<c6IϽ	~���"O�I�ao�2	�N9�!�U�㸤"O���.Ӫ(�(4Ю�[��#�"O��b`���;e��2��Z0ib�p�"O(��'Ȃ�y$iÖ�T1`\���"O�q�#	�}*�|�u��a-���"O<B�Â"qtM���91t��"O�2e�*M�����d�r�� "O��W@�4�����X����"O�*1
�S.5����+&�b� "OƜ�3�2��*��5<���"O�a�`j�#<U��ue��:�a2�"O�1���S6!���:��B&$�Ҥ�"OnsU
Q�BqNB��E�P�"O��I�B˃|:x����ׇw�p0p&"OjHJt.��o�h�1���;Z~��"OvZ�#�2ײa��̞9K6Y��"O��*ulH%o��X CEU8lh���"O���UӋwN,��SeڭPg\��s"O��[��K/j�H��*�U����"OZ�q�؝\MT�BoHX��Z"Ov-q6 ӡ.O�8��̷C:Z��"O�a�&���kl�P� �i9f��"O�-J��J�z�����	����Av"O�R�-.�
��tNQ�!Oj�E"O�Z4��>=^������s��Ek�"O�����N�@��6��w�����"O��h�hJP�!�J� 4L��""O� �Wo���@�ֈǱ?�p��"O�T#���[OƄi%(�]��K�"O��
��������O�G�ʸ�"Ol����ռ
�D`Q�M�e�T��"O�;F>p�6B "�\�$H�""O`��dE��D�b�a��Z8���"O�8R�&�&��p��~V@A�"O�԰&���n���`��BL�p�'"OZ��'�^����@��ECr �"OT	����%J��2�	�VT�+�"OD8H�]�"sn�ߡ�$	�Q"O��
��Ř^!A��O�z� ��"O����E�XI ��9Gf����"O���!�ԁaF��T�T�6a��H�"O�yjT��w�b�ѠM��!K� b`"OJ�hq��N��]2lE�I�XY�"O����@3L/$\��͑D���"O�9�E�?A]���o۳PXe{�"O��"ʓUL������Z'"O�A9�0�y7��'j�8���"O
��L��Y��`�Vlu �&"O�ɠ�(' �
���(�<��3"O� �y��]%K��IS&�-�~��"Oh��v�6	���J������b"O�Q��̷}b�Z@I�!�B���"OdIY� Q~+2I�BK���"O���&)�_�%���5J͢�3W"O��
��f	���%��<;E3D����-$T�s$D;��yk��5D�P
���QZ��(T�.g���Q�/D�`۲�p���8�'؂$�FG�7D� ���L"g�U�a��dZ!��+T�t�aő�C�����R5j��&"O���L�Q�"%�
%c.<��"O2���f� |3�RN�]�P"O4�I�P<Ri r�A0m�L=ڢ"O(�s2�҉]{ơ��$C�|�J "Ov�� �)Lx���,T�v[�A�7"Od��!��B@����/V$a	�"O�8cH\��$��ƈ۩z-𙲀"OH=2f�V=s��4��rzjq	E"O�M�썦C���C&� �L]�v"OFq�Ĝ�Uq�-���i��օ^�<����/T �`Q4�t�` P�<!���+"���,C/�R%z%�JO�<��+
�e�(J�׃f���i�F�G�<�EHf0�9!$��]W��
%�l�<!�o�9?6��[4/V枭��`�j�<�j٠4&Ystj��D(��_O�<qa$L+}�����3_Tm���DK�<�)ȵ�R�i��C�
 @r�QC�<Q���Pf����	X��3"ϓA�<��#��Kn�dK���'JF�<IQ��E ���D����xcBb	�<�d��NJ�Tyt(��g�x[v)�@�<	����nV�K��J� �hIk���q�<&�T�(��)� +C>v�jqKq�<	e�	^5ꤊr�D&z�HH r�W�<y�'ԁ]�9�Ac�:�00��CR�<����'J��Q���SX�t�ӄ�J�<��ɞ٤9�f�>)i����a�p�<a��%ŮQJ�+��;��4#�"�C�<Yec�6Qj�aDE/7�@����g�<�� �(H{>-a%/�,>@�E�C��|�<!�Kه(9�u�gQ%|g��v�x�<A%l�7T<l��`TC8D�`K�<a��1\g%�a/͐0Y�%�Q��@�<q5�]�;��d���� �]A�"��<ɔ É-��}�.+čH�B�<)(F�� !�5��9$&mhoz�<��K]�7 �g녎	�0 �~�<�G�3��<`rJQy�V�{։�v�<Q!�Bx�z,�@F����R��W�<��(�`�֠���R$�y�<�QJ�.+1LL�"Ow�����AZr�<�bO#*2N*���>c��3�"�k�<��)��,GhР& 3J𜒷h�c�<�M�-4��[��]�0�i���t�<1��9E�x�p�i�^�n�ɖG@f�<��H��E�L}�G��o]z�A�m]�<ٰHH:%R�8��.en��@s�<�C�ɚp��h�	�-n��E��%�k�<q�G��W4hpRMZ�xx�|�waQi�<�Ģ�K\��I�Ϣ~;t���z�<Eaκg�P=��Q-����)�L�<�`f�
��4����o`�#�`�G�<� ��ڐL������^�GԊ�"OD�
�f��z�th#���6�0D9E"O�,15��9Ɗ(R��#�d�XV"Ot����30)"��B��W�Tt�$"O�Y��+�9�,�� Fi ,	�"Oа�+�$i�����ӣ@ �Ȇ"O�lS��G��*2�Ě3��Q"O~����D������e"O�ۦj� ���+be@+�>q0S"O6ء��А>�I!��Z�ff�T�1"O��aO�<>�X [''��-B�s"O��"�)*ݞ)x��^�.-��"O�����!�dٰG�V'`�  �"OZ1sg�8\댬�c!K<j� ���"O6�ر6:>h������U�"O���W1~��-#e-Q����"O<�a�/B�<��e쁳D���"Oƀsg��9p�Rպ�-1DA`�"O�)@�f�0��ы�
��du�U��E{���C=_�$�� Ǜ7I��8Bm΅#0!��%&������z�^ݠr�YV�'�a|�h��>�9�I�@�t�������?a�'&Ra2f�X�|HP�ˤQ�ε��'�@�!��$r[|�" F��h���$4�g��[@X� �=9Ы�����ȓ5�Lh��Ӗ�^`5�
u��l��F�Ѳ��?y���A�IH����Go�87Λ�	`�P���@�#�f �ȓ, ��#M�W�Lq��"�^r(!��\.�Ib�K��D=#�/i�B%�ȓf���PC� ?�<|���-�Ґ��nS��`F��<-l~�&X�!X�чȓn~J��s���F��4��ȓC���E�z�*�"��o�XɄȓ �zm�P�E�s�tBV)� K�مȓt3(�I�K�N?��)6��J�ȓ;޼]�%DA-ONV`Q��BD>���?w��S�}���Hfꓡ5@�(�ȓ��e�Q�Ș�C�!��u�ȓN�,� �a�
��q#�	r����+	r��	$W����V�ޭvOrI���|Z1�U�9��u����&^�$	�ȓ<�BA�M�%6FV�)4N_Q=��ȓZ0�y�ǡH�P���&IW+��l�ȓm��pd����	Ԯ?d4��<��yA��F���V��`6���ȓN�:���%�0�^ 3���}8�]��@��M0e�X�x�u/V�ȓ/�0pQhSiV��b��+v�Pa�ȓ���A�Q�`( q
T�U$Ȅȓ��!+��L�XWXzv���V
�%�ȓay�����ȼ]��Q�� M�Lt�ȓ	�� `�jU3L,:��捝y�I�ȓ]Hd����*T@���I͚p]�5�ȓ{D"�j�.�3j�ܒ�꙯X5���vnJ ����sK�b�X(,1R��ȓ+�b!��ZT'�	�¤]�I�H����<��H�T��`��N�o�p���g�<a���i��M�@�4�N�;�d�'n�]�f��!k�A`eĐ< |�IW⇻#��B�	m��( �ջk�^���E.v���ɷ�h]�6��!x�#e)b�y�����G�C�	2|�]��� ��(D�R�m��� /<�I}��ti���>����G�58ȵ{�@#�O8ib3��� `��.4zjk�CԻ|��s"O�ɚ��/���E"ˌ�m�g�	,dì�8�4��O�(eppi�,�8It���v�F���'���� ��2������ 3�ݺ�'?��Ey���Z�:+\M�?V��U"�@6�!��D?2Rq�@��8`h��@��4�铻�>�eI�=F̊
sW�д��h�<�U Q0.с�
�^�p�Pe�<	�.� 3���P�_0~��Wa�<9a��EO��{1A�r������t�<�&�p���`��%B�]����o�<����8�̅��KD�ZEBd�c��s�<�F�	J��W�6DB%{�!��\y�d y��.)�ⴓ���v�!�Ď/X��zg%�2��I#0O	
<�!���b���H��Ց&����'�� �!�D��!�V��KQ,[�\�:`@^-Y�!�����}�`k�!H��|:�ҥ.C!�dPC�� ��W�e�"1�q�	�e`!���M�09�E֮"|L�0,��Z!��@̙��DQ���0"-�
	K!��>��`C�g�2T!��Q�1!�G��,�P�$y�tѣ��2}!�}�,��$��2\<�VG6_t!�dW(bF�<Q�K�S=HI�f�PCO!����]���99|�Ƅϛ^P!�DY�#��$B�蔚r~i�e!�`L!�K��p�fȔ?b����f  z@!�D��(0�@�Nˆ�4�P6lӡ&:!�$��py�1�ɓ9�tT)p��z!�O"!���@⌣wJ��v�|!�Ĕ�B�&��!L�jcPypb�Ӏ�!�Ӻ,���AhJ<lQU����1l�!��� �H�(C��F`�!�هS!�Ď?q��k#��5p�h�E�:y�!�D�(��2K���]+3��!�d
�'Z�mZ�Õ�a��e	@�AM�!�d�+<��9��%1��=H�)4Ok!��_;|���Q�ϙ��÷&;`L!��"wJ��9��4s#�dZ��Ͳp=!�d�f�xy�<zy�1�
�,!�D�.���r���/ejژ/t}XS"O��F
�0(r�)7�ϋ,��5QA"O��jsmħ���Id�ٟ.`�]�F"O��Y���!v�p����R1;�"5�"O�XrdĭE�52�i�lK`�8�"O��3F��-�cR#�25�;�"OL���H�%�����4?:0=��"Oh�!�#ߜ7�>hZ!��);  ��"O���H�
o�@L���)
����"O�Pǭ8"�t����0I˶�B"O����͇J�T�1Se�g�T{1"O�p�J.7�>ԡ�=Z�`�f"OLY�B@[�Ff}Q��j�$59�"OD�xuI�%�T�p-Z����R "O�����[v��ֆ<J��P�"Op�(��~�~�R��.ldZ���"O�hcGcK9@����`��{x��:D"O�a�ccܪ��ͺ�OI�)VJ�x�"O2	�թ�!%�1��)cB��Qd"Om���� ������P$B���"O�y�Q�2K��TOW6	��h1"O.��S��o���"� \ӈ�s "O�B��)�ؽ`�PXf�U@"O� �Q31oݹ\�&���
'ul,��`"O(�@�W�(*��y�D��:�Z��`"O|�&�ݖ^&����#9>L$"O��*� �(��В��^�h��r�"O��Ă�,�-��#�2D��� "O����Jc��G)�Dl��"O���c�\�9ήЀ�H��F2l��"O��8q�P40��g�#���g"O��X�͙�$p!�G��1L��"O�9�` �.�
ta3�ԳG��$�@"O����H�$Bx�1�Eܦ	���0"OX����L�X���D��nAV��"O�X�sE�'�YcsAk9 ���"O��Se�	�X�q���=" vͺ��'�҉��S6�2t�J���:VH��|�+�Jښg�j���O����O�|0r��O����O~�Rc,��ƚ��F�˝R��I�|�D�&�#�T��d��
�6���Ń�l���G�UR/�X���:A���%��JD�1�#�'����iW⽢dHF�_�͙��s�dY�+^6�M�����D�O���'b%
���(g�:0 �´+��p�ΰ?ٳ	�5i�mB-Wۀ���o�~?��aB���T��XRdB9�u��'��Z?I���Od�Q��ʈ�m���4n��q���?����>�r��� wt�@ň@f�-�C-�,T�AIq��cߠ!�̊������O�'�p%I�	Z�D��녃$�.P��%��J��B3A�tA"�F�,T{�`Vt�'dEs�6��fFi�^��~R�d1n�"�d�4A�����.%fb�4�#=P�L�[�̸�&��/W���4�D8��޴ɛ&�i|z4���:#12	C���[U����'.`�I�]u�W���!�M�K<q���!���c+��H�b<	v�Y�μ+Cj�׀�l��ХʣEޒtrq���?���"ț�HQ(r���cJ�
8�H�r�i ҍ[@!M4��XA��Y!�� ?7:4�u��K��Ɯe
g��$\rUy�n��~6��A�i�Hy���[+��E�<��a��M�HB�1��lBc�G�_�n1ArM��A��'���4�?��O؈� �;�MP �z?ڄ�1�ɩ�M+#�iu�`�>����F��+O
����T���S�
 ]T�r��?��N�4,��h���?���?���x�$tӺ���  \�!S�B�7K��L�afq�d���Ԗ52�Ǔ;|EN�������S���'�$z揁�F�68p�GT�&��fB"U��p�TC�@{�y��ˀ5��)�?jl���@ƶja�	�]�F����;Pr�q�v�o*�����<iO<����?Y�OR��0MK,uT�xs�
gx����,lO� ���&@`q�So	�*=�y�G����M#�i�ɧ���O��ɮ_d�, �]��nEeTJ��O;G6���bY���	���IF��Q�I۟T�	;fDf�@g�P�[��I(�%�O��e�焂;;Jjh#�oיt7���l֋M �h�Pb+�/]|�[�iSDD��R�ށ4VV��bȘ)Uv��a�O�3"���	��/�NI�&ʓ``��ɉ#���p�d��ҩ��Q�Q���f�-�MS�����O��'9|6P��@݃z�!� *����; @�ƍ�v��Ɂ� W�i�^m���'�7-����'ݺ�գӨ���O&�pm
��%I���U�2�4��1
-�*Z��'b�kQ�G��U����o��"�TrfQ��-6��xiBU.�HO�)8Bo�1()Y��)R�M�0�X�ܳ;2��r�L����)�O��n�2��O�*y�r�Y'pxl"tH�3�P��'��{�W�D3�ϝg�����C��P���7�OrLlښ�M#ٴh�P���Lv��Ǆ�:���O���OF�O�b��x�m
   �   @   Ĵ���	��Z��wI�:/���C���NNT�D��e�2Tx��ƕ	#��4"�V����cV�m��g^(X���Q��H��h�:ǮM0TeB�	9���#�)�M3�Gٷ
��n�����Թx�x��	��X�BHM�Qp�Đ7o�x��� �Qf��`��T���!�M��$RK����? XQ�&E�R	#��01�t	z#DF$��	>mPV�c��B�W��r��y�RN� 
֔�'X�P7�ɮG�pd g�E;����3!�8r����0k'}��E�~%�e6}ҡ�r������P�B�Ʌ���%�T�c���.L�V�����R�ē6 �!0�L����*�jq�u��`��*�%��~�˝�h��]Y�6}�(Θx�
�H-}��K�K\���ƽ�������:�8��0V��e�H!� G+5>��S�L�:�Ґ7���i�}�l�҅�!G�bK���tg��mo��M���+I�F�zl��8O��B�)�:7f�[C��F��HQ��'/��I�g�>��E�V���Ƈy�ns<|'OL:(٤a��$�<���
5n0^kĨ�OPm �-��`��D��<� .ЃS��wő��H��6��Z�t�X���E(d�UX�fB^#Kpr�N��`�LǢ����)�ޝ��+j)�I�灰l��a&(��A�V�ٙ5z�$�dR ������?�'�5&g�(}�b�"��J�lF�z�бK��('�&��D݁0t�T��h��# �~Hi2>OZxAr�J�n,�U�0D��-�f]�补�ǷZo��O�#�ǳVw�'��$P��� ��99vJ�!x8� "3+x�|%�D��*C3#`��O����^7#��k3A�M#��k��a�ؚ�+N9N��-:c\>Q�ҙ�pk��o��[��9#��[�LI�Jh��F�' �9C��հ�:�)Q�R�Q/O<A��A J��'�49��FR���8&������k��`��n��=K��Q֧ݥ|�$�,��_�tb�b�Ё��Y���4)�`ּz��#+Ǖ]ڨ��D!  @�?�"O�丗_��R�34+V-I��a*O^��Ϗ=�Xp�%"
��A�'����'��{"X�!E��2�'�0iCA�����Q�� 	H��p��'�����9���:4e� 3��*�'N:0�Eǖ&-���"�nI��1!�'8��&�/�B���o���Ly�'��8	����&��jbLE�� ��'؄�c� P�P����˶q^�Q9�'��kV$I(!e�0��G��o����'�>�����#1���X�䁈V�d ��'�^ ��@ �����2D���	�'󐩑�B�(8�T��?s�Z	�'un`�0d��<��m���@�'a���'�ʨP��E�K��t�Te܎5�n�{�'�T����ǳGd�j�-����'�fE�bB_�^�2�8��ъ-M��`�'�n��/5��YPE`�,��QZ�'1�U��B�	y�d$#�@X�,�8��	�'� ���bY�8w:�zCM�1S��1	�'�����M�*��Lk`�^�t�Ƙ��'�Yz�L���Ʉ暵n�����'��6Ϟ�X�����h�~��'H8I&"��t��#djv�I�'�@Q
��E�Qa& �)pI��'V��Ԅ^Q�=�5&��jd`�' ����A��~f�I�H�������'S�i!���;4C�up�-�����'r�iQ�F�.����n�4 9�a��'���U���u�\pH��U"yx����'.���j�<Y��9� �V=o����'}@qj`�X����(��s����'d�hS���NC�M�P�'\=v�!�'�Iq�#_�)�W̸xb�Q���/�'���T"�V'Y����ݲ�ȓ1��a�-V�i��4��k|��'ў�|�!#q��� �Y%i">���L�<���?3f�sd�_k���1��I�����0>QA��8R����M#��<Y���j��<ϓl�1��a�:a�T�HQ�[�=�ȓW<������1S<�P�o_54�P	��3�����A�%r��p0�GV5/� �ȓ=OpC���P"���S*����ȓL�<��4�$e��qsG�^.cY�\��>�Ah£^�vґ���X�I��8��ފ��wƛr���ӗa,FO��ȓx=����QN��E��9�4�����6ní �8��Ʋ��5�ȓ�Ĺ�rn@�eB��7L��0�ȓG�v��aP�&��Dz�쏌 b<���_�<���6	��Ⱒ�9Nȇ�0���b'@E6h3���H�ed)�ȓE�z�;s�Ơp�T�R��,3��܅�+ݰ�c��J��Qsa�;��ȓ$��%B�ǘ/��=3>��ɇ�b�"acr,�"i�-+1 Ǐ�\ �ȓ�0��m|x	���ċ<��݇ȓHɎQ�&!b�B�Jd�J�0�M��P��9�LY= *(���6�R�����hH �E�����o2Gu�0��%��X���� y2��F�0TͲ�ȓ>\H�%��?B�� �)F���S�? |�$�_5O�������,^��e��"O�%�
=Yb
�H����f�e�"OJ���`La���z�ܻ;o�A�"O�D�F#R:r�8���JPn����"O���Ž
=��0#�,8b�p�6"O��!j�GVvT��	�PB�@�"O��s�ĵr��0:"�*52}#�"O��X�^4fRա��֭')���C"OZ8 �B5xXL+�A�T����"O�ǁ�!�J�X'����� $"OX�G���xv�sE��}�T�|��'>n��#�؋~~x�� ؊Q�"-��sl*�P�4z�`��]�l͌��"M�~��x�ȓN��Qy�N��AY�\�U�;�R]E}�i��h��8�G�.zM8��\����V"O���W�sr��j��������4Oj���bͶV�1O?��2A�B!bWnW�G3<Y�� 5D�Ј�kC*i�B����$.8Q���3?	v�e�j���I�b-H�Ҷ	�f�"c�n�����)]�ƥ��ENj�������)����Oy�cΒZ�>Ms@Iũv�l:��OQ?���ķZ�)�N�}H9q�B)D��`'��%g��@��Px���v���2����Ge��Ac��
Vr���Ǫ"^B�	"G��u�eaܞO;V��ņ&j�B�I?y�����۳n����&�"<��B�I������V5�h�焅#��B�����rq�H�u���`�'jC�	4,�8}S6�Y�cp�)F�C-JC��6!���Ж�O�vE3C@'�(C�*NUJu2�����`!�g�r��B�	49�� ��3?�ᵩƈ:C�B�ɞ4��������>��T��[@�B䉈6H�t��$�$	��Ҳ�ߜ��C�I�b���q�%b 떇�1V�C��RQ4)�$!�uX�q���֒LzrC�	"f\�84�A��v�r����0B��0�.� &��#ˊr�J	ॡ"D��dXX���A�%W�/s]�V�"D�$����_���D
7d��0Tc"D��P#�ÄTH��Rs���X����.?D����̜�0��\r!ED2�z��Մ'D��r�&ׂt�M��*=v���#D���Ä/41�!�n�kitm��-D�����B'Xs�������@19b�,D��B�5W@�H�FJ_�$u㗏?D�DS4�1K:�`��=�����<D���/вU�S�eΫ"���qЬ0D���Ү�2�,*�X��R3a-D��W��MZ`�Б����q%�,D�h�4nQe�\�j�L�z'�u�,=D��:�(ܥYt��u,K!y��+ҫ:D���d
�GM�񣠜�g�4�%9D�$CS$A�e�-r�P�2�S��6D��K�b]�Xt�I�_�DB��3D��!����w͸�) .]�us�
2D�\�gM6>���E5Z�j+�.D����.��A�nɉ�b1zu�P2f�,D�T��C��H�%b�ws4`K�)D�`��l�[���
��z� �a#D�i�Y-g��C i��#�L�4H D��)�Ĕaaj��ɬ#���;�,>D�����d��]�����,�鋡�0D����8�5Hr��}1��4e/D�� BI�!��V�pPe`�_~�9��"O~�ے�nڦ�kA@˝4m6�2"O��4 ;vT��,��j4s�"O�XR�;QZ|@0�T�f۞P��"Or�x�όp����K2!7�0� "O&���)���`�Cꗼ�����"O��ubl�42���i�h-�"OXJ��w�v�����1b�ޭ��"O^����1r= 4�г&|�}��"O�S�m�\MPq�CƯVdɸ�"O­��IY+s�L�RU*��!JF|�"OԵ+�DO�v�
(hBjԡrBL��"OB�����1���b��"Om�蝀���ef[?	rD��E"O�+���v��`�GC�\�as�"O�T۲�Z�\�:�
���@�z�yD"O�9�G�O1�T�;c�R��TY(�"O� 
��+�(0�ۦD9�pH�"O�d�(�rw��e��4*��B "OΜ8rT�i��8sĤ�1_3�1��"O�L�k�*!�6�	$
�G;n�z%"O�@Y���iOʝ�2	M%% ��"O	Y2E��)�z�bT�^"|)�"O��6��LHDEkSF�#c�:�:r"O�D�H7y��![��0�ဢ"O0-j��8>)��kź	�L��"O��!4	ۇi��8:AJPk�y��"OL �P^�L�Dx��N��\ ��"O����j�k�j�k�(�#J�����"O��E@$|l$a2�Ȅ�:wrJ"O,L�W�1F�����1\t�8T"O� u�1{�2�(��G�>N���#IΦ	ܴ_t0 ��'�1=u��'�B�'��֝ߟ����rM�����^�@��g�+Wʌ�	�}�6��T-H�I:���剟FژTIr��a�@͓�)<PD�ahŪ��P���4r�}�F�~����%T�\�%�JI�U��D�� X�I& XB��I1�M�A'�~�'��P�C���=]���vETN��9��ݱ�hO?�$_8\��q���>V������O�yݴ]��Ɵ|�ב||��V��Z$�?X��ٵo^� H)�
r? 3-u��$�O|�D�OR|��g�O����OVܺ�fˊy:&<{�#ݣ3��LRҨ�=���{�$�VP�*	�$��-� M!#Q�{B%	ep��J�5A9�%��[�'�|�C�TIÎ�ڗ�U*��� QG�>MQ��[��OR��g&#(5e��K���*�*fֵn��h�'�b�4��7M `%�b_�=�T��QO�?w!�Z&q�#�� H�h�QO
�=��Dl�pn�ty��Á|$r֝t%>}Av�_yU4i�K�9���2#)�ܟH��G���L�a�i�b ���3\N|��"�oEN�aQR�iє��]|P�"�I5ʓ[��Ŋ�� <� ��Wb�%c��]�ĉ�-H�3�)�%%7`,0^SX���T%�P�c�{b꒏�?��i:j��7��0خ��`���2���&J���`�	�b>E��?�`�
�AX �[��K��p�D�K8����4ћ��iqh5
�i��E0��͟�F��=�'�V��MC���?y���Zᅏ��?a��M+h������Z��<�� �b���I�N�=/;\QZp�]&��)f�M�#�j`��W>����@��[�Nc�Ü[i<��]q�Tr � �m50p`��AXY�F9Y���������L#V�!JZ QQz\2�kZȦqᗉ�O��	Iy�'���fN�<@\�!�T ��/CQ��B��~r�'�ў$�>�ҨgBv��F��;)�x k�]�'M�7��զ�b\w�ؒƈ�2�R�i�J#��(�r��O���A�nzD)k�k�OL���O8��I���M۴�þYJ�Q`���"M`��䕧]X�D2փay�RS�&*;��ۤ�OK��@1��D�,Q������������D$4�KD�_�h��IxQ��[yj�	ׄ^b�䎏�P��`'�@�2L�9Lqt`�P��t��ȨC���?a4g�?	лi�����d�O��Sf�B�����G��B�����EO����>h�ʨA�B	�|RKj�R�o�yR�'}���Os�I�S�E3�������)�#l*����_"��	ퟨ�I���SĆ������;d$���nZ�m�b5����N�E㥆��,*��$��-4����/6|�������\{4�݌K�����'�`\��ddCF�T(^*�c�\�J�c��Z�j���0G~
� F�ꀥM�j	Nu�V뉠.l����>��m2f�*�#ԙZ�MG;c�R���Sn�f�|ӎ�O*���O�O
ёu�  �   "   Ĵ���	��Z��v�D�8@���C���NNT�D��e�2Tx��ƕ	#��4"�V����-	���џ4�$x�s�X�n,��H��>��#��<S@5M��!�'T�uw�-�����n@Cr���Op,���/e��9�bH��,� 6�D�{6	�/Ol�Q�X��A�O&D��鎺=&�݃ꂠP�8�->4��Ѳ"U��[��C�#��S]�3 �E��h\ r*�p4Z4p�I�S����H[:Aʰ�2.݀^�� %�>�-^��>�+q�>	��.�ŉ�' �܈]s��C���RǏH��	#(����%'�Q�	"l��cb��|�h�JXj���J��P��A@��k?�rD�ny���4�>��IY ������>��b����S�5^?��Q�Ω`R�p�.*��~����`�7�����n�I��-/n�(����E+�u�U���K���'��e��A�/�f5�' �9��@\�:_.mΧHcD@Y,�l�'�'j�����OX 2�Ă`�'���E�Ƃ�~��O�|����G��l���])�< )e�o��T�N>Q��9Lڒ&�4�`�X9d�66��V�p�1S�D�7
��vۛz�IV1��F�&�Đ(��X3f�>��Ɵ(I,Xգ2m�B{�)DF�X��q�W=�~��O�5hr�I��ԟj]
5�0���רӈ]�����/�tm�'p��ɺA_�	�[�X���'=�����?Qg*IjY�{�)��%��`#TȐ.z��ă%:�P�O��w)j$�rF�>��;O�t���5Ű"1�@\�J��OR�Љ�F��ē�y2B����b�)6Jݤ�A#�ߟv�$���KD�p�^M�˟1��B��-�l�2Lܨ�qp���r� ���9�p�LN(H��AӴ�ܹ|�ʓ(���L�`�	�G�*� �M3�Ҋ�ppC	%:� �˚�<
(�f)�'ʾQ��`��' ų���}~��ѳn\�5JKj��m!��%{V �  �B��80̤�t(�5T�0!�T�S^+��i��H
�0J��[�53�xhH���k�rL��I���Yɓkb�����4c�TR����.�h4ѱ(2D���u�Ls�h�҄㌊|H�҅=�	�F�uc�BǕ��\��-�<o�����uk<%1�"O����_�%�:��a+��H�*���(�9= ��YF�x��!�g}��\d~m� b�*�VR���yrk@�����ߡx,`,   �
  �  }   $)  �2  ):  �@  �F  VM  1Q   Ĵ���	����Zv)���P%G�AC ���W�H�Ąa���8F�t��$!�~-�S�'ll\�02��0JY.:��1i$i k�(��"OdȚF�3E�ę���Lz���`.m��BS�P�4�j�!��f^�bd�%"a�\�4��X.*Y�gc  UP��FM�<ռ��Ţ�I�e���p<�k�K��l8�<1�+��&�	���2�z#��N]�l�˃��l#�����gp� $mȷ?פ8k烞np��Ǡ�iW��&
�0�?q���?��>����O��)�L�}G:qqV�*�<h���ZLy�!T��p>���&B�EBb��o���[M�pyb���p>YG )$wv�i�F��ΰ�(�@y�'��?�r�'� �ha,�5ЎZ��ޗe�d�i�'�����ܚL�#�ςV�bEx޴+ϑ��Z��)/_f��!([,����<!�v�bu��f��IğX�����]wN��'��i�x�ā8��1Z�JΓ/��4(�g�R���:l��N,�P�H��ي)A��8b瘧[��}g���?���5	�84�0�Z�{�H$i�`�K$!��C}Rj�
��BgiHB���2Y�!�d@�$9�I�!-֘���Ш+��	��M�J>�l�f��'�"џ��i�,�uU*��/��0�\��v�i�x���'��'� @�P�'�1O�)�n���m�g��!B�V��ў���//�'Hײ`��8�f[1�N;)DN�G{Ҏҵ�?���ӌ-ਙ�B�C�R�����	Q�!�C�	�R���F�۠T�E�rub��$Ta~�DӛIo��qJ�M֢8�� E���d�2�hnџ��IJ���+.Er�'&��ˌ818�%���%,w��U�j�P�h��O�b��g�8�Jm3�H�-a��r�f�2_(& �	�4��"<E����z�� V23��@�c	W�B>!�<�?q��|���F�E�c��D���*V�*�xB�	�1�t0`���w�܈��S"=����$>b���I��l�L�rՋF#:渊ߴ�?�X4ƹ����?q��?��`9�s�%3r� �UW� 9�GȂI�x��*#%�$r���dL�@�+�ם�?U����-0�xt�@�N�c�a�Dۊ��ݚ!�
�8>���׀k^�a� \>�� h��^pF���R�L�c��CW�@B�ί�$�7mu���d��H���
��x���ĺ��' ,�t������z8�Ty�4�?1���?�J>�O�Ӝ'�<a��/�r���PcGAK�E���b� 8�'0����\�� �'����|�b�ab�U�q�x�S�On/�h�G�'���'�2�e�=�I�ΧO`����Xp�4HRe_-oT��A B�"./N`a	�@���z�X�cf�ԝ5a��Bc("�Ȇ��) ����;N�&dy$@ '�BUr'mI�Q�4�ȓ@�x��hD����ڴc�"i�ȓ5&Dj�Q1HQ�鉴ʲud��'pt6�?��(}����O��Į?��%��/v~�+v�4�d=:��}�|,+��O����O2��M�O�b��2>	�Q["J�?i�H{BH����=�t
B[�O��Q��b[;f��Hi�+Ls�+��DD={�R�;§Up�-���ĭ���7��r����~���S��$)����R�>�؇�	����N$V��	����R�8��������%pȩܴ�?����)�*s���d�O�A:.��}}@� �^&1Z����C�-�C�x<�5�'FϦҴL
g�(z����|���d��lr�ڢp�ā#Ak�)V����'�b��Ҥ#�8�!�ލ_(�!�tݱRT���@��O�P��BV���ՊФ7�-C��')f���3��֨z����|���ܴ32��1��P�"�����*4���?a��?�)OB�$�O.���&�z蹢lԧ"�k���<aJL#�n��&�$�����)�<A�����W�W�Iڲ%�PN���4���n�ş��	�(u&mh3aٟ���ΟP�ɩ�u��'-�1K�i:q)��;�U���8���<I�i�VƺX����"�0<��.)J��pP@@Q�=�T=y�Ey��w=(�R�aO�Fxax�-я�&1��k�>n�\dx''�򤋮-��?LOH��r��D�|����X�bO�����:4m�M
3D�
���x�nզ幈�4�֓OȌ@TC��,�(��c��h8p,�0UI�)Č�O����Ob�D�������?a�P�����[":@��pa%ů"�@Pz7�N	��`�M��-:�|j.>C� "?��mEY��G�?T����6�+CAP�5K ���5ͥ[sf�l� ���&�'m���9in=��O+r���W&�z03Ǹi�,O��D�O�On���O�Y:W�A�'4$�����0����U��٦�ID����t�9/���'�\��I#��n��DԦ� �4�?Q��O6R�����?���y��;(�-+�K>�<�O�/f���/M-c��'�ҍ��F�@��J�
R	xC�Ӫi��A�S*�0� �`F/v���e@ݤ<���=��'G'u���l��P���Q�;LhL,�� ���B�Y,K�L��!�7‒#�5�~	�=	W�Z��"ߴ$��O&ʑ��f�1N)�[�o���ip4����D!�i>�Dy��R�9��+���,e����F�?�>���i��7M؜E�"`(wo��L(��,�14���ק���������O��'}�����?���(gX���e�"&�  �
F{�v��7,r�ɦ�2��q���Rg,�������,���Xh�aw��b!p("L����9�H fh��05%ڛ�����˕h`� `GG�[R�'���� ��*�<��0���uK�l�����I2�M��i���SMARqI�+H���6a���'���	Qܓ?<Bc��>"tEy��()8�Fz2�u��n�t�	�?!x��!�:D؃�ȬC�d��HC��M;��?�Q�A�_b�]����?����?`�����'�d3v��w����L�T�;���S�l�9'�]�q8�<���a�40�I�gbDE���T1o$��B�I�8�%�X,S�a���V�J #�A�|�J�(֐��B���y��0E^���g_� ��i���A���^�}_"�(LO� ��?Mb] ��ʬa�|��"O8�a "4 \D0R��fi���ƿ�M���i>$��{eiǆ`�h[gG�W�@�i�JN`:��[�a���|��П��I���I�OF�� $?�l҂�T��Q�!L��n����­Q�F��*�4dy�i\v�'����ST�%�䅆�	�4�s��rd�9ؒ&Ծ{~�`�1&���̀Q4�_�'h�1��|����btDN������C L�x��iQ�6��O ��?���������}
Fث���#�>���Մ�y��0tT�5�����B���� �M#��SF�ֵȅ��\���Ν�R��6��O<�d�Ok�M�Krb9���ca0H�j�-������a)��'��Y�O�w�� �ٓ��0 "��ӤS����m����0&�H��=A�o�2\�j�ȳ[^q�p�8p�N�p�]�X:��1�O�T����G)�U��Ex�j!�?�W�%iY���bM4MBţ�y;�B䉦g��p��!N4n(�`��%~��$MH~���.��]��\���@��@�,����G��lZ�(��I���=%���'n�p"�JZfÆ�<sIЌ?���+�
_�^�@�Ҩfti���;�|%iuK�*�1���c��<���܈6�h��g��O�]@#g�(Cȡnm���K�=ì��d��L�����l�f��冻W����10B�'��)�	�O��I�e�TAj"�0�a$��=f�B�	�E�T�u�ţ}����q��4�(#=����!R�yf#�'yv�TL=8
聡ܴ�?���YR N��?����?��{q�N�O�<��&$s���jH���i�d�|y����p>1�)�Q� +�j� %���[� �{yrHQ��p>Q$�^]���Ѭ�'2�8��ly�G��?���'�:x0��М��HiFO�����s
�'��蒢.S���ҖE�g�:��ڴ"����D�0�bВ�l޷����q�Kc�^�FND�W��y��������^w���'���"'!B�2x���-8Ph���Ԝo�6��$�Y����W�6}v�@�`Gv����ָx��}�ָ�?9��"4\)'ΩN��(зÍ;C�!�Č���볠��:���P�]�9�!��<U��,B��]��삃�^=C�����M�M>	��=Qz��'Krܟ��Em,@�2*�+u�P͡F�i@+R�'���'����ԫ2K� ��,X�c� �ԟ��C�瞨1�>��6��6f��9��IY����$���_�dI�!KT�x~�y馹�4�1��B�LI��N�} �pq�	$�b��QT�Oގ�yS�2yK���j/8�"	�'��p�N^ ,��\��jT"1
F��;��	�����+l��T�gc�ꓴ?�U�|�	S���'l��'n��3҅Ү>X�!�I�9�Z���wӞLKFa�=H��7�S2eR�e����>��Q>��SJ�U�� R7e(��i�KR�I	��~}��u�@�4� VH�b!���g\7_@D��l����I�::�0��ǌ¥k$�C�NY]��$�2b�(LoZ֟��O4��?a*V�^?�AŢֻA_�Y��T}r�'��IO�'p�J�Φ�&AG�]������y48�Ռc�0�Ox�d�x��Z���	�?M��
�0G��([�DˉQ�@�0X��M���?aG���5���?Q��?I���Z������dv����!b�h�#z�IQ�(8��>��ѧ���d��8Ӆ�U�Ra@��{�hI `G��j��X¦P�>Uȅ��u0�'u7���"n{�h��'�"�c��L%+�����g1t��(O�h���'�7M�Q��ޟ��	h?�D�8@����Hػ]ǈi1ŊCw��|�'? �I<1���<e	��\8B*�a����]0�4Ct�V�'��6M�OD���Z�'EY$]���Q�(WJ���I����A��J������?���?AA�����O��ӜI[�PSeË)p�)g��2K�Zh9F�Mn(��I@� ���mˏT�2�h��l�(��e�N9: ��1���y@�
}�;$cM��9����0����3a]+w\b���3��O�� 4�p�#�.w�r��A錌G���3�"O�����o�!b�!���Y�"OZ�y�`@7��X9 B�>L�vx2Q��c�4��S��RǼi�' ���8�9�'��<
�t��#b���I�a�2�'�B��KS��i�iD�GR(�ᯄ>RLr�xB
�.��!���	}@�UR��Đ>S(rey3�N�<�t��V�G}6H�[�ڂ2>yx��$`�%�a�Ff�X�I"#ޝp1OV�IB�'��"|R�KTnx���(M
&���0O�n�<1P�R�%��Q	�L�#Ll!�/]hX�d#�OE¶�Bl�mY�!فSz�}�X��qCA��Mk���?�,�n�����O���}��JXxF��0n#?�8�m�tL��*��A4n���\���b>�bG����o׋Qm�1�
�ܟ�	c
R�'ܨ%���.�0q�/	W�O0��c#C!h�4񢀚��9"�'1:D �kɧ��l��)>&2\S�a�(D���'�4D�P��a��rƐ �����(��1�p�?eؖ���9 ��υ�k�H�J%����M����?�����	��X��?y���?y������bT£�Y�d��l��U�-�5	פ?��x�E���YB,�3���k��Z��`c��)!$ĸA��D��C�Z0q)	���C���dI�TL�C��ښ%F�C5�� ��I�ik��X���:`��e��[��;f��HZ� D��i3��s��{�(�V���R6�~� Gz�O�'���BΆ`� D�!��� ����;~�h��'a��'"L���ڟ��'}�6����!4�|�����d�5j� �G�'O
t e/�@����'M��K;6L)5�G�O���d�C�J��{�lь�?�0��  ����ÇD�Ф ��K�o�!�
j�F�o��B���c��JU!��.�ҐbPO� '���$���u��<�M{J>�ժշ>���'T)���ì]�J�����+cP�an
~�A�	ʟT���e˶��f��j����IS�`�H���O,�1�/�g,\x �� M��1���dٓJc�Q�Q�!x�0s7��7Cm�瓻�F�K�i��q+L��1�R'�X�=Y���P��xܧ7����MJE����勃�H��'G"�'�~�S��*��dh�ې	�T����d6�T
���:(�.)���G�_g��U���(`�i|b�'��t����IܟXar�Fe��Y6@,O�Z����M#�� ��^�x��'t\�Q���R��ḨF]&�v��9@�i��H$|�Vi�HT�$b��T�}K$�{�k�1/�p{]w��ͺ��iؐ�* RWË�(%Z$OR
i�&�D� u4r�':�)���O�	�;ft���1CU����QI~B�	
����gB��K��j��Sw�"=�B�"/V��*��P-�ЯK�F���4�?�����X��n���?���?Y���n�O\��"	�9�h���I8f��SAj&]	2< � {N4b�%𸼗O���1c"$UdjeI�&Ԩ�#�#v܉�V@��=�Șa�KF2x��'�O�}7�R�\3De�?&���X��jU��Ol���O�� �'V��P$���V��0q�nf���ȓV���)�]�H�j�I͙
j�mZ�HO�	�O��j�v��F�	�>*�-K��S ���p�DҘ,nd���?)��?i#����$�OJ�Ӈx� AK
B�D�e�1���{��28t`�a��6{�� (�g�'(�B��#��%ӁD�t�ja��-CX�ɐ�*?���u��~� ]#�Q���u�=�Ѩ�ϟt��ߞ]p3Q��4+�	�%��M3���'��>7M6�,���U�1P64�F�X�d�!��˳O��*E.U>{M@BBLP �����M�������7��hlZ����	@�&�_�ĸ�&T	^�rw�Z�1�R�������ӟsd�*(�\��rK�3~X�NJ,V�F�ʱ�^qD�|"��#1� "Џ�e�6�<i��^q(����E��ҡ�/O�W��%YA�7H.��A%���&�L��WWG��<I��O���ۍ�i�ڰp���8��� w/Fw!�܌DZ̝c$G� �2Q�f/��xa}""!?��K;3^ ��k5K��Ӧi]~}�l�;r��7��O���|� �9�?	���C&�\�;����M6JǾ�`��i�J �5f�+m��=��Ԍ(�:h���@"Zs����I��������M��򁘏F���$�	��Ѕ�SzJI!�7�&x����Ovx%�`G�8L�!o��%�t����'~��]�ɧ�� ��P6��w��80d&�2ō(D���e,�n��5ѳ�	ͺ�p7�0�x�?KU'��GF�P�w7zԓ�iͰ�MS���?��Z#����?����?�'����Ơ����$��̋m�H�(�ӥ��a�1	��`�rȂF+�/�=�jE�x��'	���Q�X�T��J��3�$0����d�VX3T��(��(HU+�:W͌	Z�O��1��2B��� #����%X��"#C�Ol-��)� ��ѥL4���'�s�l��"O��!�>Bv����=v��
'�iú#=ͧ��l*`-1"U�;�̄���<��	�v�ɻ �1����?����?�%������Or�����)jB'$��3�d c�} g�O�hAM!%"j�qa!�.7N|��	MFh! ���	\8���"Km�,ð�͌d�;7�"���A�+;Z4h!��I0h�d?Y�Ջg��<c* prfώ�uʭ�ȓ��<0�h(,�v��˔?su���}���V1J�D�@�>oOB��'Ot6m4���3T��lZ�x�	x�EK�;
r\�Իe~��3�LSȦ���̟����(23��MNp��K�3G�.dC�S�҉˷PE��Ń4P�AK�'k~�����
,��I��N#���V���o��%���( 'I�X�}D{��+�?���ӴS�p��tH.�X@��m�0BB�I��n%�䉄�4�0�@"R�_�*��d�[~bg,�R-K# ���rs��-����IK"l�(�	R��N�e���'h���u%{J±�rʜ�MZ�@zU
iӎX9���OLc��g�C�tQ�U'�9^����ڛMs�5�ɤh�"<E�D-PnLP��C
=a�|���%υ��d �?Q�|����>2Q�Xgpd(���
���q�'!�;�.�Pʶ����0��ڋ�d	a�O�N+O�N�l�I�l�#�%���p�4���O� &�y���d�O��$�Oz��;�?�1p�@�qd͐����gȒȺu`��3���`Ӹ�h� .�� l~���(�'�8)ѪЀ�U%.�����'9|C� +d�J��SD�'f�zs�[$x*�=�����Q�,O����'p\��G'w� dS%�ە}�ta���G�!��3�Nra�/�6���۬����&��|zI>A��<ʔP�fr�����!?@�#	m02`��ϟ��Iş`r]wSR�'���A��\�����0`&$��AU�0�(�w�ȱ`4(�CdGN	p�š���K3^�z��ͱaP(=B����.�v%�� �ܲ�J
uH��GG~���;sH�+#jv ��\D�'&�E��:�@��O�gw��Y��I'o��u"O(a�reZ7��)Ӧ1p�Y�"O����^�,�L�0ЩT~	̼�DR���ڴ���l�17��#��%��ějdz�m�*�4�3%ꜪkY�;�V�7��B�I8F�v!q�Y�2a"E��#ة}%�B�	�K��Wś����l�2{VfB䉴;��l����Q��U����Z�C�I�5�AbCЋ13�!���̓d��C��Q�KE��%"��i�0h��cC�	�6+�<r`	��q9�勷�{�0C�	�K���5���`,
4��9u��C�	�,�T�� <"����Ä	'��C�I�2o�4�E=������ymrB�IZ���Js�Q����wC�)7v2B�I�*��Rra�-)�<�����A�C�Ɇmh� itJе 9�/��B�Id�4r��1 ��h"i=�C��/h���F0J�J����0V+�C䉷r} ��ɸO��-0�V#�B�I�}7L��5�B:-����p��:MS�B�	J�b7L&QF R@'���bB�=^|��2�(\�����U��B�I�3�Jr�	1A�]r���uɰ⟐q�&	v>�S�ň$�������ea��>D�H
I�!(��f�^�X�H��N�� ��N>�F;�gyB%Ęd�yZ���{�ش��cѾ��xr)Up䩢o�49H�ҡ�4.���VW�jz�I�'�',��$�Ȩ#'�Ұ-ϐA�\��ϓc�� д%߰\���'Z�t �ݓV�D�;�"D"x�1�'�J��g)J�"d@��L�834�@L�DʄhC� �fi��`I�?|,DG���9W�!�2�P�<~�H�����y����0��x���Z�9p��cF)���'
�����a�f�0��L>i�J�cZ���`°	�ٳ	�'mKN�Vc�p���O���Ţ�&����-h1NH����O�a{�N�)
��K&��&�Ѱ'B2�0<Q�oLqP\"4���}���p��=,��D�9tnȖ'��K@!��S�? �H���N �c0a\���$X��r`�Ѥ]�pP�F삀��hF�D�LKݴP*�㄂>D� �*�$�y�(E�xIȱ��ј��q�gb�ARu����<ytB�9��hH~�=AP�K7��M��׾װ���O�B��(BT�[oG^�Q��Y]9�86���g��D�r�?%��$ӑ�'t`�`N["�0�@'�*F��dh��$�-����0	�|* ��=X�A#�Y�hZ��+X�+,X�K0D�hs��̏r
��2�F�E�j��v��<)$�ڈ[�ĩ!��-bZ`;������� �W�	c�3K�P�"O���ƃ�H�6�sǎ@��
�p�A�>,��ъ`c7��E�P('�1�1O�@4�
rn�{��ڌ�{�O�B0LvɄeh3ˇ�q�d��%'�A���b�DH�v3|YcA֊�p=)a�]�pR���+?�`h����U8�tJ2/�e��m£n�J�oZ5<�P��� p�k����B�5p�����!��`׭��i:��'���AŦK]Ste��	�U��>�GbM*-f��ꇇ�N�^=�M-D���&��4����H�S�6ȩ�)�/2��I�!�<�$�������I�;�, p�BU5u<\���/U��C�ɱ�n���7w2���`=a�����*	�}q#+ �O�z�HP�/��\�v&��Dh+�'W���!��AZ�E �3$-�d�2e������	8Rz�@�fF�PC�Gx�����]!�%�Cⅵ\AR@��]��O����# �	�Jƃ�K���,�����mZFp�,ӳ����ࢗ�&W|ACr�<D�@�B�C��j��٦v�b�ﮟ�y��^�G���qi_7 p ƥj�Q>��M({:R���&َL�����*D�L����5(����W�\.}�JU��ߴk��\�`�Q���ʧ�W�
]R���|�=1�gǰAl�R��A}��ү�i���*a�ԏ=��I1g즄   ͖-WPYX&l�C1!��jB"BPl�ד"sHDb����k�27闗[�*�D}2�L4&��L��"F:S��y�7�J��M���C����SSG�iH� ���y��jIxQ��CX�qUmY��~ROʛ���¦��J�:dI��R��MG�t�P�ep��+3B�	dV����W�y��2��z�P!�Vs��A���!R�L�G��& ۺB�=�ו~V���nE�E�A�it �i���B��~��*j.8��'��h\\D�®�#+������ >�����M��<�@�#\O�܋�@)<�<�I���l+����ɭO���a��4������ � �Z6큪+�ԁ��jްd<��E�3d�C�ɥ����킡R<�%;"C3��ɇMW����*�92B�Z\��6�'o`��b��U�z8��+�3r�nB䉑G4Ҵ!V�	�s$.�Q�xF'E�AP�Eo�2Q�De��$�F�i�W�t��e�ӃX�V�0%�E=h�F�����q�PeÕ�9@���ѥ���h)h$�\�\�-}zH0�Ӌ���p=���*Tx]�5�K������v�'~��Cǅ���i�6�Y(�
l�޴UY���6b���� �\.i����'�R͑�P(�w�(��`��'����D�����i��&�����t�O�x0{���--'Fh��c '�����'mlɰ��L��p��EA�3�8y�;[NDz��i��(p��K	��'<�qO�$���äF{�)�������e�'��Y��z0Tq����ND{84�GI'  c��^`���ǁ2�1��V>ْ�R�-Q��"'a�X`7��9���Ӧo�d�R��S4m��aC�i���
�%D�(s�$Gv��#�
xD ��F��� 8���>���" �&ZM��a�Q>"��M剡�S%e
ax4
!D�@��˻E��ܐ��Ƴo�vYS�#
>0�Z�	�ݦ�y�I�>K������=����#&��1+�MQ�SM�A�jT���[!Rζ`��D+y-�TY2`��t@ ��emT��ՆB�C�J�!5`�q7�,
��
qV�1�QE}RW��P��DV�0���a��M���^�:k�uxB;9P
���E�y��V�b���W(*���RB���y��&f<Sg�\�Y�`�"aV��y���|Iru�%ƒV��yb(�
�y��ds����d�3?�����4�y����DyկS��ZL�s!��$ڋ>���D�`�r���xJ�Ss'SdVa|򅈺{�!���� ����&D��;��K�f��3"O��WB�2���BoK"8B;w��PF�\Sf�Ni�O*α�P.�<L�ft:PbU��@���'���bˉ�E�ĀCI�Ufm��c�<m6�	�L<�D�>qU�['?x*���Ɛ��Ff�<��>wt����BX��I���_*��uOG��.���L�P��wɊ�X�R�d�͞L��z�'��T>�j�/��xyd�U�O�z)� I�(F�F�9D��)�f߉_@X|`���=V�
�kv�:�	��49v�_��?��c�%K�����(Ѐ���oE'�6��ȓ,%.����O�~�pE���@��V�.X��7��X.Hx�� �����*v�h(��&+�:�ց^Y��B�	-N;԰�h��8�fl���5>4�K+/����dֆ_�LX�K1O��i -Q?����S�) ���'��Գ��F%� �Cľ~��$�1Ò8�>�A@�PF���dP�X���d�o5tB'��Uz@P�2k����'+�m�6E�̃����C�������!knX8�e����!���P�H]!��.M���R�E�ta�s����Ѐc�`�P X�D=�
@B��I?}�H�0� �r�!�/�k�o�.�x��zA�r�LoZMZ�R.c'���4h'ȅ��ńe\ �0r�'R ���(�pNE/8����	ϓN��)�tFUx|���U) �(ܺ��ȯ�ӣlV�\�
=;P�2$�`zA��%B�����4�0W	+�ğ+t;1	S�W�px�T*���OK���	R�W�l$��{�(̩a~�B�ɮC~:��������1f�ߟ>7n�8௓a*:Yx�����w�&�g~�`L�'��xP�`[�_I�"FK��y�<C�@\�n�BÌ�i]����1PԵaV�(0Ę��yB��:��P�M�*7���z�.�<��=Y��Ʊ�����;,7��v*S�*v�q�A�48�I�"O�(ٗ��!&�X����$LF0y����1^fu!�lOf|�&OW2b�F`����$۶b�%�ȓvyr���s�=���Zn�i�/�`�P;K>E��'�aq���e��aP����U��'춴���G��Blqg�*.�x1�O�bj+�OR��Ю�N��v��l���%"O~l���q����mO�kT���"ON�@0�_�Tt�q�	t��s$"O��������$����S}:��"OX1#����H��hJb���X�0v"O��� H�MplBM�%�0K�"OZ�����#�bd�D�hS�ih$"Oܠ��V�")���0�r"Ox���C��~8T����u�ؘP"O�Q*��v϶أe'�N�@v"O�\01C(���h�Ɵ�^�J�#"O 4`�X�@c>��g&ޓD�N}��"Oze14�
>)	4�� F@TB�A8�"O����n
!%��Gō�IE�Ѹ"OXA�3�ҭbh��++��8�"O
�k���[W�9��1L�TL�"O�DY��W�+���u- 7J���hE"O�X�B���P�j��-	֪�R"O��iv��N3B��"���3"OrMh���MͰ�2���&@f�7"ON�A!��@�c�� �3T����"OЀؔl�H1�P�E��/R�q�"O�����߁*|�5��E#
U�<b"O�����4T�V��TB�?!R:��"OF�Q��9����`�#EWH��&"O�t $_�^˲0�s �+kR�H0"O�t#��#'�n�c&G�Z�|��"O)�r(ϒ[p`Y�$O�"hҦ"O�@`P��#(�R�`O�*%�a�"O��x���+.��[VmW�(z����"O� d�g��M]T�2qX�vf��Y�"O�����.z|�ۄ��?�dӆ"O��8$؆�IE�X�7�b��"O�dP �]p�0��×�2ް�e"O�`��P�=`a�tL�OxPȄ"OZQ��"B�,Մ�pă]�H ��"O\1 mP.��K�BM��'��yr)F$6=����ꋢ9.M� 'C��y҇�PE�% �eI50k&� ���y���X��m����q���@�FB��y�#\/Xvpt��ɀkw��
����y	�I#�(	�i֪W�� @� �?�y����(�naqE�U�IŘ�6,�%�y��ɟ -<!1�a�E� ��݉�y�H Gvm
a䉲S��S�J�)�y"��.��p�#��5A "0�y��/^h�I�Nշ]܆�!Q,�yR�	�F�P�@Fh�~, ���+�yr ��_P6ʣ��dbڬ����y�%��&�n��!���0�"�]��yҠĭ"f(qQ�� ����%I�y�b�^r8AWh�������yH��~����� =��Y󊇥�yى>�|��V��!D�:�o>�y��C¦�S�"�0w��Y�Q���yr��*p�b�g�Զk\M��)�yҡ��9@��;d �6o����S픬�y�.1�0H�fP�p ��"���ybG�36�h�3&�l8�)�C� �y��.7LA��f'	0Z����yb�U�,0U��ΰb���怙��y2���Y���;��V%;�m����y�.��mZ��^�?䈍8�k�/�y��s�0*6��+5衠�ޑ�yEY�2��%ZSN]�'s�<�����O��(f)يR��<����d����i����D�_��5i��F�a�1r�'@�;�G'�xY9GK��T	�'2*D�(�4�1�VK�A:��'wa`a��)�EN����@	�'�j�j0��;sq���`�����'�}��dܞ4�V�;`q�L �'�`�;�/��I�� �E�f��']��ո'\J��A �]3�\��'�zT�ĕ�z��8+�صV]�=�
�'U�@�`ϝqFpE��C�;�n`s
�'xbT1���*����2p�M��'�h<�2�0:0i'�2$'���'Ǟ����]�)���C����,R�4�	�'��U�q!H�[�V����'�		�'B�<{7�*=�aI�.�Iw��9	�'��y��n��B7���d�kc�@��'7��@�(H���d�ǣ\Y@�Z	�'���3�"ݣ����\�Y'��b�'�ظ�2��t�<���.�5a$h
	�'��YkS��>�L�W�[r���Q	�'����rM�x�`'C۞x��<Q	�'I���v+� ��p�K�|���X�'�:���+);�Z�c͕q�� ��'�������1��U!�%>���0�'�LY�
'���1�S('����'����DYYV6U �aC S�(���'nBȃB�^�J(���iAw~0�
�'�Z��L��I��o�LK L��'�P���å}�"�2�����8a��� ^�kT� ���g�[�
�H;�"O��PO<v���8�#9����$"O�l�5�`�d<ɦ��<�ZMJ�"O������"}j��GlbF��T"O�X�"�F�1����M�Gj�G"O�(:��ZF�N�j"	Td9Lk�"O�]R��Wu���B���RL �"O�$�s�J�(Z�-H�����"OM����ZtBMy�j+h� $"OX�@�m��V�����i��!����"Oڜ���ĉ4j��0�)X�E���"O�e��hK Sm���!+�U&$qB"O�|�%j�E�j���ʒ�U����"Oҁ��\ /�}� �X�N?%�2"O�t� #�+�F�#���;.�#�"O8�!�=(7��X�G�*�٦"O��Q���r"n]��BL� ��"OH!9��K�0���{b���x��r"O�2�ƚ.�.y�p"�&n>]�"OzY� L	��H�`�B%B��7"OY��-i���j�+ �Z��d"O�Q��5[H2m�Y&z� ���"O(��!,Č/�YIk;�nP��"O�D �M�N[���� ���#�"O �УeRQ�h��sfs��a�"O	S�� GB��d��.5�$e�q"O*�E��Wt ������"O|�pE��:�& ( (�$��+G"O�0!���f J�mT�H���"O
0�҉Q.��I���<�<{�"O��Qψ�D҇i[sd��%"O(�4�� K����C6Uw.�X�"O�Ai����,�nl�(;v����"O0`�*@;,��aTD���V"O^�x2N�7A����.�04�Q�F"O\�+q�D�s���2�Ζ�zP�� "O�(�Ǖ,:f��ïјiP聑�"O�`q#��W�X3e@�?}]�툳"Oȡ��e_�#\�I�MF�s#��1"O\m3���-5��rR�T�C���P"O���Q�<8�$�3#�b��`QP"Op��Q�b^ms�+Q!&�8���"O�@ӯ0�L!�c��5����a"OTz�(GNkZ��JqU t2��{�8��F�{o�Щ3��QC��QJ&D�̈���*������A��j�g�\����eN���'�?���f均A`������ � ��!^􌉖 �:OZ��p*T�!g&�a��e�_��Dx��)�!DB34xE��fې<�� S�fQE�<!v"��]���J���=<x�
�'B�<�+��o�H(+��3����'�d�<1���V�`L��).�������t�<ɡ�N ?�Nͻ��~���*�$�s�<iS�+zPɳ�ÒuZpb�j�S�<�-��,�D�/jh��cS�<	�iΘd��9$bU�=N\ �D�M�<�U�^%;m|Q�$�|P�|��I�<��`��}�>�kEC'j�p}��B�<��$�s�NepCMX�q
&�yG��v�<�7j���V�Q'�
a�n����}�<��f����Ӊ��U�ܽ�V��y�<1g�p}~���Ƙ�>�XA�-�K�<�h�K�(d�׍P
%�tX��r�<� "#�-C�6\��S���_H<I"O���CP�ZX�N�*V�ˢ"O����׻
��9zWؾ\���"O�����d�
أF�J��t��"O�H�1 ɝ8g��N�|�aP"O�DB�nS�0E�p����,QG"O���G��XDԲp��(����"O�\hđ	�IR!� �ؑ"O����C_�E;T�oW�CH4"O@��C�'�ȵk	1$��I'"O��`��M�8��U�vꉕa,�!�T"O�0�����Mږ����*�""O�AÇE��VQ�TJ����*)JV"O��c�E9�z��& l�>�rf"O�x����-{4��$�
\E�	�"O��	�ֆ`ق	���3�{%"O�uP�d�!p�b���Y.��2�"O�u¥��;$Z�EG2 �{`�'f�'���6�Ǿ���`A�\�fҔIb�'@%���4)��3�A^�- �}�f�6CV�O�OG�0b��U�N`����"�UO��	�'�T��D���8�Bq숑\dt�->�A
�>�>�n@q$gM��i�I�d���� ƛ��_�=V����+R�(�v=*��.Y5���s�'��1�bD�*�4Q7��+`��;�87�Q~"b (��	 ֎ $ ��Q1��-�y��]�b����ŊF�.��؃G�L��'>��(��?��A~��'�0P���P@�&{ҔC�	WB���_++x܅�6�B5��<�G#7OB� �h�"0��	��mʀ"Ot@b���7���YC�,�NX�d�i1�C�I;J!�V�D�\���q��: 6�B�I&m���"��4��}F	�"W��B��Zp��T�"m�)k�,�pdB�I�.$�S�`�梱�Ԑ<�(B�	�k��8�h��d1�ģ#K��C�IO>��#B�s����HH2�B�I"��q�" vt�D�.y4B��%N�%"a͍S~Pr�,�FPC�I�Z����=v21�F"�1݂C�	��ԥ�O'K�q3�JF(B"RC䉪 ȅ���E�|Q䔈1/n��C�	�$�F���ީL��#�����C�I�_��Ǯ�������?\��C�	�8������;Z j%Ђ�D[�B�I�(ΌI90��DŐ^(y��B�3����n�{Cd�b�(�10�nB�	�?>=1�Ñ)�V�k'��7jZJB�r���桙8�����ɻL�B�$+��i�慈U3�ՂW&
ΚB�ɪ�R��ak��������B��B�	�d����3�nؖ�O==�B�ɻ�a� �Ͱ�nEx��3l҈B�	�w�<I1��4*��$�B�I8g P�+ѪW�E��=�H�� e�C�I�	�҅Z�[:psZ�XR'J3�\C䉣]\2tyU���&��<��B�I
H>�B�.Fds^1�c��x��C�I�KM�� ӎ <2%c��G�j�4B�I�#k6����vm�@��IE6+�@C�ɦl��:BшU^��7
ؠ*�B����z���=���WoT�H�pB�IhL�-PT�"c���jѡOuHB�I 3�be�7��1�O7�&B�)� �e*@J@%5�^�Z�\["���"O`�� l�P�A0E��&��#"Oԙ�V F�=� ��=q͒�"O�+���	U���"��v��#"O$�I�)4�u)�Kȑe��]��"O�,z�H�":t���
u��=3�"O�i�X/S��b\7���rC"Ozy����~(1�ꁟ��4��"OD9RO�0:��#h��	�"O>q(��ǧ[�"e�7ⓖ2t���"O�����q5�̣�@�8bf��K!"O��ە�E?T*.�*�MZ[�H�"O$1
Hݔ%��q��w;���b"O0�{���D�(��R���G4��"O��b#允QC"9jBl�2uz��v"O��B0	�1�v��WJ,Y��Y ""OP2�@ԓB�>��rb�?�	r"O �;F����� A�`)�a�"O�-
��C;ج�cOS6q���"Oش�E�R���GH�h��N7p!��P6���I��h#2�J0{R!����D8r�z���'�,I`���5�@� &Q�|q�y���&\��x�ȓOG`��!�!y�ѫ�/S�C�ȓ���B.R25����Q	�'Z��M��!oR�h����s�1��O�(F�>�ȓҬ���m��	H$�9�D��Q�L�ȓQl*d��`��7�j�H��ϯT����ȓ#��! 7cY|���̄9�pL�ȓ0����q#�!�͚B�T9�x��=5"���V�5�t$�0%K�z�<�ȓl��	�`D��i+�)��P&q�ȓN�>{��Z�m��i�"
��V��H�ȓ.���OT����u�� /:Z���2�X$zp1>�� ���(�ȓM��H����w��D�-F�Av����b����A�2#dM*����&�B����i��͒!"k�9��˿�b��ȓyж⁜�o��YE�X�Y�L�ȓ%�@�� @�?      Ĵ���	��Z��w	�;V���C���NNT�D��e�2Tx��ƕ	#��4"�V������m�� ���ߋN<�+C�f� ɲ���k��%Y䇃��M�"Z��.B5m���A�c2�	����X�z�Z�������ճeF���J�\�@ �l��}�*\:N��_;l`�X�t\�v��E�R����iH�*ǛHC剭L�$2%^*ur�^�|a	�y���'G���w`O�9a���2>���Q���t�dH'F,}��5����.,}�[�XI�e��'JF��}��呱�l���F�O�*���ލ��G�D�Ƀ���ĉ�>!��Zf��M���;�J��~$8�4��?}2A�G�5�ta9}d�5Tq~��A+;��8���B�XqR�Õ'�(Pd�M��ʆ*o?��<O�<H�F��yhݠ�U%΄�B�\�FJq�R�6}��ޱK4�+�2}B�Xa� -O�,�V�0z�l���66h��xS�'��Q�E�Ɂ��I-8xxFd�F�I%g��p���"/���*��ɂvebT1���c��'��Dˀ�@���H�;�BӦ�#qnS8B=��ĦGS���W#$?��V�68�|%���$Շ>%��'�,}�'� D��E��l^6�p�( h�	yPI���H7p=BL>!�b^;~����L�|hx'E��K� E�bB$���;r��|bA�,C6e��'.+t�U�b���0��<hNa��OF��ʋ�O�'�r�H�ʉ���P��TJ��:g�!#���n�7�p�O"��E�;��'�Q`��ΐ::I�E��
��I���~=b� �nW�A�@���|�Qa�3&��V���i1 E�Y5P����>G��eF�v�@�B.�w�F(�'����mI>��uc�m���
y�ɏB*��`vG/c܊%���/L`~z��nj�O�mZ��ۗ`w1O~�P�Ι/�40�$�-�r�b@I�4�8C�ɦi� �  �/@�@�$$��VH1B�"Ov��%���z�4(ߛ/�nX�ebG!�r��#�׀�p>�Ŏ<G^0 �3,C{��8���Uo��ɔ�N�r���q�{r68f�^"x-^`����%c�Q� e�SH<9G�(IΤC4b�D5�9)�i�y�!D��8+�a��3t�7-ٹ4Fc?�b�R�4!C�
�{���d�8D�1sDP�UR&F�a�v���1s�t"�	J�a�b�g:�0�?�'�4��K��9�5��0y�'�bшB 6u���j�!�P�(90��h�BaQ3����2q	���#s��xb�ͦ��[&FP(B��j��K���<��D���0���j�,�����!8��d���0�����D�5|�2�'C��կ�/S&��5�Vk�N<ٓc�F,�(peX1�� �mڄ��OE�Y��Ϙ1/��!{��"Sb:�b�'��RC�9V�LxÎ�6"�q)�ёi���aq&ѤwlXh�$*���OZ�> �ر�h4(��I�o�>+����{X�- g��he���v.gl*��"0f|q�R��-��1�v.0,OX�b��+�R��d��w=�=q�'fRl��7��<u�q���R��Z/� ��P<[��[G�MH<�7��.x\4a�V$m3(���$�E�-�(���,�%8�<���U3��O�N��,O/O�B|r���w�~Ey�'���#���X������97�X�ʣ�r�~!�ѧY�������	���+��I�e��s���=|�B�I�����ˑ4܀3�lW�?xn7mS0v8��Γ;0����dU7l���!�D��N��(B�/�a{2*�)A�D*�mʊ.���DmY�Ij2-rR� �'zH푂�8D��ۣ�T!9!|����u�ib��p�'�l4�g�2�>���4��*��h`��	֎$D���A����@�f�-%�^�YFjd�<�1'�'�)������	V�tM�?5G�`�4D��H���L�@S��"���s�2D�̊�옕�b����[4.M~���d2D�d��R����IgM[�DA:�K#l0D�ʕ[�&�"����#�&%��d9D����ޣ	ბ(�7m��1�&D��[�� �D�楑�-�(p�&D��j犘�e�8d�q��V���W�$D��{�N6��e�r�3�x��e$D���S��6��Ғ�@���3�?D����߫Y0ܘ�􄇳�z�	��0D���GA���-r�(�Hq�5B+D���qi�={� re�:Wڔy�c&D�`#��F)����fֱ�@���8D�T{7`��u`h�"0@
u���cdO+D�$�S$Q�^�|��bĉ�l�H0X��7D�T�&'Q�q�z����H��Е�2D�� �ƈ���
�(ֽ(��u��?D��ۤB�Z$I�D���LA��z�?D�����	�"�H���$�rN��kp�;D�0E�%;�1�v��' ��Q��k:D����#$�b�:�.[�
��°�#D�D��e[�bM�tJG�3W�w�#D��5�.�����D	$C��ۦA4D��y��
�1U ��4y3���Տ3D��գ;k�bŲ��SU��;a�2D��{��xji�#�S,r�p�p$�<D�h�� �Ob"�p�W�f�r/9D��Ғ �3&���;��S�'w�b��2D���ǧ�7&�J��#��l=@�3�
0D�܊�+�tݲM�f�BH�.��qN)D�@"�m2��4s�n��Nf���k7D��$��\+ȈIe��&P�Q�E�?D� �ѧ�_����ů
�?9�aJ3�)D�d+ѭ)e�.y+�G(���3�(D�����e�xtY F���p�,D�� nu�0�z��V̇M<"y*#"O@��+K6t��Cc�_!s���"O2|��2` �����l�\H�D"ON1( ��;5���&.F/f��v"O^a���FL]T��
e4�` "OL�8�a�8\��,����s"O����L��T�D&/g��#u"O4<��k y8�b"�O<]�~M�"OT�*�Očb�Ƒ1���<�L�d"OX� ���d��f�2d�~��g"O�횱k^�C��LZ�ܠla�mi�"O8L!��iJ��Ʈ�W�0	�"O  G���s��� F�F�R� "OVt	5l��QqP��e	V �d�Ѳ"O\�� ��
?x���)`�L���"O��+ЏЖ h�RIO��.x�0"O��J�-U<.@�)�$U��2"O�Q�֩Bh��a��勂_"���"O�P�B�?r��0eƳz|��"O�#�)Ύ;
�-���^�_r
�	0"Ox����6&��H�
�c^��"O�����%s3�U,E�htY�"O��Rr��_���G�Ę"��y�1"O��P-ܧA������zljy�U"O�ͩ���L��8����gX��Z"O*}��D�3FQ�9D��=uw2�	�"O|�1�ְ27�A��EԌfT֬з"O��&J:g<I�$]�OJv\�D"O4}q��'A�F����N2ؐ��'�i���E�0���C\ yH�sc�ȥo �B䉏K�.�d'D�)5ıh2n�$�B��*I�Q��=���AW�;o��B�I�BN�Z$h�	+P6h�b�B���C�	�H�RX���^�P| ���+j C�I7*���e�*4��`��#�B�I�F�B�x��Ǜ2�p5��+I���B�I2Vvv�sO� ?��Y&M�.B䉂{���XҐ@�a��^��C䉸*����&e�9������j^�C䉔erNX�LA�U�!ЯV}�C�	�}DX	�4B�4\ie�G�Z��C�I
+�V$�WfυP�0�􀍏�^C�	lc;�쎁`�0c��18>LC�	O�q�i�.hh�rb��]0C�	� t��C@�A��8F��4��C䉥.�����E�Q-,��W��5d��C�ɐP�8�㢆�8ֲ�R����DC�	����S��L��hq�p�&2v>C�I\��e��6�@���1�C�	-~�e��#��\B:M��!$�C��/8$Q��LD;#��M���Q�)5�B�	�H�,Y"u� K�}(��[;N#�B�I�^�@tå���*���X��ՔJc�C�	�ז���t8�Yzs���~��C䉍yPΰIcM�A��e�c�C��(T��e��3s��@'I��[�|C�4e�����ԝ�R!�iI{�fC䉳N�L�Q%��rb��u����B�	9�������7�Y-nC��~��0+����P��Xlq�B�	(D*�2i�={�l��!��7Yw�B�Ƀ<@�Y��DS�b�:DΎ��NB䉧b)�h��̑r��M�����Z�>B�ɅL����e���j��%��@�q��B�)� �<˷�*���rA@t��1"O�����3I������{ ��""O��ԍ��'��XCn]�W�@H��"O�	�Yt���窘oP�0R$"O@�QM�y�B-s3�ߊRa�*�"O\���B�>��J���~\��+"Od����}���f����P���"O�욣#�&M�>p��L��va)#"O2��%���z�Rw��z�Aw"OH`�N)7txCM��hcRl�"O�}ȣ�.���
�17F<}��"O�����*Ǿu��cJ2'���1"O�m�"W�eV�M�R�M�n-�s"O&�)7m $Np�,�tN�#�xYÅ"O�5˰(E=H Q�B#��]� "O����o�W#�kUjH1u�f�`�*O! N/x��T�4M4*�$4�	�'5r�⡇�U���c�kD$r* ��'�5x�Ú<
z������k�=��'#��B��4R6q{��4Kp����'8��SI#�zU�6��@l���'��<��`�|e�4���3[Z	��'��}$�H�w鑅��7����'1���C��27N�b}�,5�
�'>t� 5@�I6�%%��x�8�x
�'V>����!p6���>���A
�',���nU�c*��t�[�>��TA�':|ї�D]F�H���
g��0�
�'n0i�e�	]��%
!i^�_xX9��'1`pBG��z�ʸ��'D���;�'��9J9��aAlO�A֩��'z)(5*�2|�phS��3M�(`@�'�,��Пs+PM�#LբI��	��'�(�@N�=lD����R�,Lyj�'�J��2C���<�9$� (*μ��'��1م)�,`W�LQ#G�'T:5�
�'��9�UC@1R��XQ
�U��Y��'�6-)v靮DD��ᣋT���B.�S�����x��B�F 5R�t��F�:L@!���۲ ҴX�PȢF�ޣ=E��'P��X	D�J��ç�9#�<�'8l!�$� 2����&X��ش#(�����o\X��ՊM-"Q�PA�cJ�Wa|r�|2)�6
O�`M�|����-�?]rB�tč`�쉨c�x�n��2R"C�ɿ:��1�a�٫u�(B��M�Z��B�I�x�Y!�F�
%DU��F�nzB�ɴY��x GF��YH�B�^�x�vB�	�	yЀ���/'G������5�C�T�,x��D�U�A e���qQ�B�I���\��V�_�)B�� �{��B�	9?B�qY�k?���r�h�8MMC�	�qiX�P��E=����"G-VC�3��{��t(�HR�d5qTC䉼.��\�5:�D��pΆ?~4C�	$%n$�c�\<Dyyu��0�(C�ɥJ2fa )P`0@�λJc2C�I^��2�O��`�vKZ
~��B�	#�E�gK�9f��QC�I�bB�	:(�d�"r���:|�t+�I*E�pC�	!L�Ni��͑�U��^[�%"OVE#Վ��'��2T�9���+1"O�|����]T���D	 ���p"O,#���X��S���W�8�В"O� �P�$�<��Q�	V�0��"O>�I��Th��rՃE��HT�d"Of�Za�1B:=`�AB��:�`t"OH���N�YO,����	��HR"O��!QFH7v<��#%<�Z�Q�"O��Y3/*|���I�hr�"OT����$[�tI��K/��"On����_;2r�0�NG��H��"O��&��,X�] �ָz�@�P"Or�A��K%P�2p��*Ο���h�"O�;T�ۼ�� W(K���X�""O����	�9N��!$B�
�:��!"Oj�P�O#;Έ)����6�<��0O@���\�����X�yD�a�'Z�&a{��371�VUxQa�%�qw�B�M?Fk͇ȓvE�S&E�' Ǟ������2w2��>і� K��ħ'��pT�<Hj���@T2S�쌅ȓ�֠"��P�0@L��A�ZF���m�'4�G�,O:Rb�0v��M+6�	v/D�
�"O�!��`��(�
�h�mݵS�h��4mY4k���=�Od8���ߏ+���[�l��L��|��'�b�nZ8cl��DIP�!��3p�ZRBL(�ȓ6�����L
�O�b*P�D�}ن�=Qvb1�S�S D�]R��F%|��4@sH4D�B�ɯ^�p7搤 Bt0�c_�0�6#=Y6�'�v�ҁ��%�5���^:j�N���'������M�����dղ^ǜ��ȓCM(*���']q�A�O.z>���ȓ%ԁ��io�L�zb��+�B���w���B�u>R���&z��q�ȓ��i���
�
q�H駠M̒�B7D��@��/9-Ą"KF3j�>��)7D��HUE�|��R���R����!)D�� �
�#s�ThA#M�J�2-P��%D�L����?[��i���<C���� D6D�d�g�ڔR]�(�gM�=�,z�N4D��bD�ϻwb�x��:'t�+�G?D����ES�M<v��d�4,��Y��?D����-N4u�:�x�*ރA1�?D��W�q)��@ͫZ��8��[�`�!�	E���˥"���=P��\5?!�$ۙ"�~�OA�!i�UC���j$!��%uD�`��3W�L��LJG"!��,�������[�z���H� R�!�Dc<���N^�w;�Y��B�<@�!�Db�&�jP(K�l��Mw�� Y!�d߇Ek~xs���3V�@��Qcõ/W!�×ax Q������� *!��͆u�HYӄ+X�]���)�o�)!�D�4q��h�3�H����I���h!���B�؈	�Ώx�P#P,!�dJ�l+�c�F�\�D����!�D�!;9�\�w�L��Tb`���g�!�D�,�0Ap �Ej��pH^g�!�$��am��H��ߋZ7�y��)`.!�D�@�u�،M̬fḦ́l !������ß> ^l�yb )3�!��N	�6\P�1kl�����!��3&�	q��d�e��h��a�!�d�&��ȁ!,3x��S��*k�!�$Գ�8�@�l	F�Th�f�ϬK�!�A cJ*Ѓf�	����"INV�!��	I@���d�"`�lىcȒ�*�!�DB�H�Z"˭~�ޱ��M#T�!�� ,���F�o�����#Sʬ��"O�}����W"�3��T�O�(�`"O�|y�Y�j~��F��Q�`C4"O�a*W�3}���2�L
&J ���"O4�a��,A��F B��[�"O�܊g��#R���y"��r���"O�H��!B��@���
ن>��"�"O�Z�h_�i-��Y�	�Iܠ���"O@���$3�\j��J�Up�c0"Odi��_!Sp6��Ӎ
j�Iz�"O8Q�		'C]�$�W�ę1�j�"O:D�E��:4���H�=r���P�"Or`��ܛP����&�!	,�"O�(Y�"'Z֠Zw��'���"O��{�ЏOV`�c�E�
�"OjXpL�1#��U3i�z���"O�Y�Cޭo#ܰ�焫-�(�"O��)��BN	L �=*�z�z�"Or,Q"ff��Ȗ-�<T�&ѳ4"On$�ֺ37��0,UBv��@"O(u10�D?�4��R%	(� "O�+w��wX��l�3�>P;�"O��Vכxk�eI lVC$� "O��X���\[��E�!�BG"Oʘ"D�	#�Թm�<!��"O�ȅ�[4c��Y 6N#( l��"O$аK�)V�M���Z<*��I"O�L�$kL2qŔ��E@�<U��Ż'"O�lpQ��a�~��/M����	�"O�U0�O͓L)5[X�UAA�"O��S��6�UQFP�1�{u"O���C�>Q�\k��ܘK�=a�"O�ͫP!�90�<3��Ë`�|�"O�A V�  �   +   Ĵ���	��Z��v)��;^���C���NNT�D��e�2Tx��ƕ	#��4"�V����ư/̭m�#5#Jġg$��F(��wMޔI�j��B��^C�aٔ"���M���^z#뎚/&ͶTB����T�Fl�IɟD��!V(7T�SW+[#0��ua7A�3d���V��P&ֹ@X.]�M�@Ѳ ʭ�Q�ˌ�^ly�#gռp90��"M�w�I�.ef�H4�E�I�2�J�@�:��1�'*ܥS!�C
#θ�����O�;�bG1����+}b~\dB��9}�S���e��x�:�$� !����_E�tQ�������ē?H�<�DZ������V
$T����4�U�1�_*�~��l9���_�i������?��W�����T�L��L	�[�\8���9,:\���b��DD���)O������Q���]��	0uiӵ� �"�#�6P^�'CҘ+��!�~�'`�٩��� B@]�'xz��p�I��Ń!-İ�8	���:h��@a8���x.��:��|b.���Apgŝ�d�:Q1��d����P�ɨ32$(!��7�$��R`h���i����C�����mB�H?���Or-��!:���<q6G�,��6c�ķb�RDPwEZ,��:�׆jqJD��ē�����*�?	W�ҫTQ�	j�"J�������"Zf6x !1ju`�%�>q��O����n ����Ǜ�?q�Y�s��ɤ
0���q��<`d����G9.�P4b�'b2�0�$
N}�ar�<.p��U�@C�'�� ��o߯��8���7L�����'~1Gx� P�	��~�R+z�^�@#`A�A4F���	�79(�B`j=>�c�C�2��`x���(�l��B0�xq���;2�j��'�������D;��"L_���G�|�l��G9��#O<���8yu��hTe��y�� �Ϛ,�j��WF�I�ɐ4@�r�G?�,Y����� �3ft CA��$B���"_f�<q৞, 2  ����&l���
�'�0�qޚ��Ri�)2^d�
�'��6K�1M��ؑ�)Ƕ/9\E!��D#�S��oʢjP���'"���������p>��K<�n�����Nَ��I�@�<��h��q�Ľ(�M��8J�pҥ�~�'�ynO�:�u��7I�}���	ިO�"w���y�L)7jX�N���g��$�pigoB�m���`7)���Bx��g7D�d:[9�(D���\00��0�E��y��ڭbϐ �/� -��	�Ճ�4�M���s����".��� F!YDJ�9OB�=E�$AA�l�u�E(D�,���)��?��'��u��n˓7;IP�(۽>�̩��'Ř-�
'L%���֋�6��	�'8D�3 �N?ZАf�#cr6�*�'OvyYd턒��P�u�]�)�2���� &|� ۧ��3�K+�i�"Ov������E�>���i��	�5 �"O:<pw�аZg+&��}Jg"O2�J��L��!�*V	+�Zi�<9slɓ~@fdREY"W�����Ap�<��.O�υS;3+���d�"��Ćȓ2E e9�'��"�$��kҳD��x��w/�,��2�8M�C�4N�4���s��򤛝4疉�BOӱ+S��ȓ2�$xѮ�1�5��'P0(ɤ���`rܠ���0��$��mB2	����?6|a�T!��h�歟�F8���ȓ[�n�1!Ij��m��A�h��zCf$bM5_�D�[!j��F\25��9�`4Q6�\�6e�⣞1uJ͇�(�
���xu��AC���C�	1��a�`J'�;sEΎ�B�ɒ]v���b�ԐT���7�V;O�B��
����2⋞��`�@+�uQpB��#�[v�"I\:�0'u}�	�'�s�2A���G�3G`�H�	�'��x�Ί.o�.$;'�����5�	�'�Ш��؈0�6�0.�� 	�'��`ƕ�t`��+<2,�	�'z���&��^]L��D�Ʋ�f���'��0	�7�:���G����'�ZS'c
-3��52���>@d$`�'	re(֣�gؤZ�fB0�,q�'؈����.lh��)0 ^���'�D��'�R�\��	jb`ۦ_�潓�'$�<8�-�!�����ԉ$�����'t�Z­Gzq���&�1��#
�'�B�:�	 I��H�%㊆qdl)�'��<�-O�^=�T`g��\�B����o�2:R-W/V�H1�m��	!�� 'z)<�q��\*����]^.!�&f ℉���<��iba�I!�T�L%`��&��^���PGH�=u!���ZȾ�ѷ�׋�V ���!���8�&P�}{@��b��
f!��Rm���El��|�	�s�\�!�͋���s���L��썁F�!�d8:O���o{,<pal��Uq!��?4	X�Q��8F2`ɶ�A�b!��H�H�2��%E�t �S�^j!�$��9.��[�H.�r�{���,FE!�d;`�H\:H(e�Z���(�Py�I hDșp/�pX�)�y�$�+�>�0�%Bse@���N��y�l�5:�Y�����;���Q����y�h�8E��,��"٣g7L�{���y2���k�=�wbB�X)\;d�A7�y�
�Z_,H��)	���҄Z7�y�J�6��5���.���D��y"��*=���Gϣ"x&���Ȫ�y�/�[�b��*�AmH`a㕝�y� ܍/��Y�s.[�Rr��3�O7�y�!L� �!�$�B	߁7~B�+
�'�b )ń�
;�ݺR�/�m�
�'�v�[&�ێ@C�|�
K4�
�'?8Ia���R!	HA��2bI�!R�'� �6��;�p����y�S�'�l��8%3����@�4��9 �'��țЯ¼:��C0J?,v��+�'�:X����4wjlS��B��b��� �̑vo�� �R���5�q�E"O�l���9$x��Ӥ��@8�|z"O�YiT��lcx�AÊ�@�eyg"O���֫�?��x6Á�[
��S�"O�qJc� S
 t.Y�Y���U
�y�K�" ���Y *�m���0����y�HT�QA]�Z8@������
�yOѧ$�8�ybI�:b|��w-@��y�g[�#|�s��ޠgt1W[�y�}0�TP���>j$D�
����<Y��+` !���Qx�H���	�!�����3 AŴK��[�j�[�'Jў�>��sl��(��r��	NF<�P�'!D�ܺd���N�C��B�7xAѓ�?��a��,��kN�c��I�q�0b7�|�d:4��9% 
���C�Y�5.�(�"F�v�<�eF69y�C �:m��A��ITx�|Ex���8�FM��OбjJP��l��yB���AII	;�H��q�"�䓻hOq����'LEgr��w��=����"O�ˠ��0a�V!��%��-a��"LO(�y4� w���f�W d�"O�����$��mK4�L5/�VB�"O�Ѱ�"KG���)��	��#�"O���kD�9��}�@�D�Z��"O�= ��8?͔x#A�U0����"OER�+M+T�04�$��4K)��AB"O�I1��[Z��K�|d��ӆ"O�2��<rZB�㑢�J�B�"O(���j[-"�a�!`ԡln���"O��8�l*.:k`M�X[0��"O�=�B�����@�2Q\Lda�"OZ!��K�:��	y挐"&D�\�"O,�ɰ�L%Yu$ 芀S6v�q�"OؼRD�`|ш�m�o-�,�"O.�ٗ��}�T�S�j��a�,0�"OP����$� �H$i�B�V�i�"OFU�'c���]{f
�>w�<xYR"O����A�M��B���`K~��"O��i2�ιpW!��|n
�A�"O����,�)R,3�
	=k�$�yf"O�:���9k�ʃ7��@�"O�!�&���{&�7B�P�9�"O���+P�(��֦�E~��Y�"O�+��#�x��;Y��1�"Of�xr�ͭ�080a�MB���"O&c�#J�$�d|���κ{%@ �"O ���c��A"��8t|�`�"OΔ���S� �u��!�Z�a�C"O���l�(1���ӄ�+%l\�#C"O0J� S�|�h������;�"O"�6�Ɖ'Ҭm��'xeE���@�<���ݽ/��Ԡr��"���Q�� I�<�D���dV�Ȃ�̦zmXDQ����<�1LP4�DH¹J��!Ny�<�F�I��ຐ���(1�A���	v�<�G��5�M���(Ӝ=*"f�r�<	g�)o��aC�	M��|��+�n�<)�J��� ڲ{>�ꥥNW�<��L zM�r󌅨r�-����Ga�U���Q�x�
qjDk]V�b���H(�R@C2&쬡f�
�M�<Ԅȓ������W� i��COԻ2�����$�vm0D��/��p��M
DO,���S�? ��D�,aB9r���/�(�"O`�W͖?�H�ð�FU����Q"O�25KQ����aB[y9��"O��(��cʤ��Oc��Q"O�l���4.��V�.t w"Oh�S��A�^ɠ���K���"O&�J�j�)A�� k� v@ }��"O�r僐-�nQ�#JK�{�1��"O��1�aNz�v͚2�Ϣq�X��"O61S�cҨ����6���E"O�Mb�Ɠ�i�f=��f���"O }Q�H��1p��#�|<� {r"O� � Hk�L�`!��c�Xh"OzX1lE�f�NX��T'O�TJ�>�te��O��m�L>��5���:�r��P� 0nRT$�o�o�<YEi�u����P�M�|���j�<!�
<k��裃�cnA��e<)�*��:�&A�/��#B�!!��'Z���/�E�P2
�/�,diw Odpz��4�F~r˻��t��3!:(��WП���Ǫ	.�&}�`G�F�F�84"Ol��3-��b�d���D�es]�F�O����%��=��h��3�b����i��8�����U�>0ļ�ǦV6Kl!��ɔ�����DǵO ��	5��?C�\�P(�.|NtT�4�J�RGr�c�?��?����s�(DJ5&�H�(0�Dt؞L�����S���ءp�{a~9�T�l�L	&�	��T�WfG�R|B��D[�A`���"�&�<�t��B��O.��,l~��H�3]�`
��0 ���Gӊy;2���T�����F& �z���4���@#�l��X�(.r!�B&:bM$�K[E�����׳>&j|���V%C&�|�5��?)�C�'���
/��W�4zvə��\�5b&$�"O
m�!�%��,C�T�������$O>�`���g^�h�/ݞu�\w9�����צ���� �4e�@�Z$<a2=k�,�O]���4��p=A��}1<ݓ�A� n�’�.��4Y��q�C�E��!�t�Ø(��:SŌ$V0$Aĩ[K�2��r�#0QQ� �q 2g�e!Sɔ�N�X�1@�<�ɧy������ ��q�n��O��]�G*L I�� 0��4���p�T�(v�ۗiA8���`�)ȈrJX	�
�FN���u�K1Ųyą��-Dt�`�ď�]q��P�l�BW^���dƈBI���5�ˈ1Ŵ)t�E	.Cv���r��Y�Q:NE��Ň�/}4�B�;�:e��f�b�sj�5_������,V%�{�J�=b�>E��k��u����xŖ��A��*L�d��㇎G�ƀ����C�n�P lF7T���[דZ  �����g���K��tSli����)`� (Ō�Zb�PpW�V����r&�PU� ����r^vY�q��.&R j��ȅ�*b͌*0~��8�f�=jz-a"ѱ K4,����mlF�Ƀ�W�*�	3��Ѫ;�`��Ǯ��p2��0����O׉�p>q'�\97Bx��F�l�&Ժ��	v�q�Ä%LaL����.=�:�8�A�:2Jt�\w��� �!
&�^�f���
Wf>b1��ޢQ5!��Gg�x��DJB^	�	pV�x�d�	�I�$\�%��bI$��G�G�f�|�����]��	�~�mZ<': ���Gc���G�I�lFr���Q3}�H��[�X��|�PN}���$gM�S�J�Y`O��J�� �ǁ͟Ky�d���yR.Дi��sㄑU�f�P�כŸ'����k�#p���cmџ+�����_��0W�
?5w���w��a~�[���(cg"t@�'uf��4U<���^�=���B'	?l\kE\#zP�ɺ��/*~r��S��4T=�S�YX�.իg�p�Ȕ�m�d�&6z%!��&�x�b.&(���kEE�:VB���+�d��:R^P�3E���Q��8���O>�eԤM08��U�fyzh8�KD؞�J�lϏvm���*Mb���p��J����U��>�0h*���,
��=�iZ�\�����'bD�9�OS1Q@��fI�$[�+��D9fL�	���0UP���	� S�a&�Vt ��N�w�$�3�A�$.h�Q�'��\��D����{Gb�3Hx�)JjM�`��J?t#�{d�[��H�����ϿsP�[jl�����kX��8W�e�<鴯��)Q0�CEl�pl���O�*T:��E�n�� c!Fj����.qOVqCl�"S�X�%�++ �� �'*��@�U63�Ȉ��J��舳�[.6�)%B	?�P�A	�9����	�5���f�5e�*���a(f��#>��FZ8ǄГ��$p4�����B��Q.ID�#eB�V�����x�<ɵ�
Lr��Rdߟ_��i��w?�C�!���T�˵jc���s%+�r��i���j|��BD@�8�����S�? tl:��ƺŊ؛Q��R0����$�R]h���4z�95��JJ���'���S�V�k��X!���Ԓ4��' ���#.���@2
��%���@�:�FIy��$��}���qt̒�%],	�Z��N���y�ډBL2A�A��!<d"��6�� �y	�}���U�W���@��Ũ�y�D�	Y���c5� ����-��y̉
I�,<��L�s�&��m�7�y2N	l��UJ��@S&�qH�yBd�%X��Y�+��C4�p����yr�I�$^>��'�[0��R���y2HےGS���q�ƛ-,"uspƒ#�y���	;��ڴ`H���W�ِ�y�T%q0���7��3	�p�F`[�y���q
���oӞZ:6�0����y/޲�*RW.Q,:���oF �y�fH�z�~�zva�":2E���\��y�/�/r֨��a�,O��<�@
�,�yb� ���h�"�	�� 9��ٲ�y�T�rD�e�
<�
Ia��F�y��B��aJA�ш|�����Q��yے�L�f��f��C���yB	"�� ��j֪؂B��y��aƸE��%�H8�hR���ybf.�h�7��+K�.}��.�%�y"ܑ^���t�9�t�8�Э�y�H�7
	<ԉ'���0�BuB#��y��Y8@D|��$NV�#^��ۑ��y�Ō�gSj����'�b��Pj
�y�KT nQD��a�:$Q�m�L��y��=�>0j�/á$E�h
� �5�y�D�)N�BI"�O�m^�"�X�y�"O51����*��}�)"��6�y�#�?Ux��T�ϡ0!"uq"����y��H/T��pi�!��JB��y�`+��iن�7v�n�@���y=O-��sn��a9|L20o^��y�ϗ�h�3���N�������y�%��u�>�[����S��	�6��yrFĺo�D�K�L`�)8���yri
ml�(�$%ң;+�%dU��y2n� �` �ŀ=<����,���yb��/Dt�mÐfG�g� ^��y�h[(F'�atMG�m�T��F ��y�mZ?;���n�f�ԄrJЍ�y2F#}�Rtk���Y~^����R
�yR'�Eшaɠ(��9x��J�E��yr(�=>�|�����2qz��fB<�yҮ�nw���a+ ���Bj]��yҪW|�.��+H
$�l(;��P��y����6�"�AV".N���E�J0�y��[� !�)��6%.�xp.+�yB�IL2$��GV�;M�hg�X��y�);����Y���SKҀ�yB#�[���6��r	<�J�����y2eEb�L�QC�;rL��/��yRB4aú���	(Y��`��Ƶ�y���#����ѺB�(I � .�y��U+x��k%�D ;��R܀��	�'�@pa�Ǟ�S��ंk�|���'�4���� �T-�Ӆ��b�p���'V��%C�7� ��BiO�_���'�d��&�ϯA��I8�+�+Ubnx�'�$IP�j�;mO�"�&K�PƨI���� ��{'��+ AqE*�,�"O8I��OM$}�D@����u��h�"O�F�+q�qq��XR"O*����Ŧ�Rxq���q�3"O,�!�kM���a�3+� ���"O"%�傈|�:T	��¦w��Д"OʡY�
��w�����_7����6"O���6�T�;���9� �).L����"O�����W��qu��1&��"O��JB�^�!��Iҳ��$��"OL�	�̅x����d�5^���"O*Y3t&�?{�1�jʀ��Q�"O���ũM�ʀ#�oӠ��(�"O���%\<I�b���5�� "O�$X6�F}	 |�%�.��Y0q"Or����<{6MH"�
s�� @!"O�EK7ΆlY���r���&���)�"Oz���O%8T�귋�>A���!�"O�X���=c�����Q�޼�u"O4a)��1�`��Y�V�l(�t"O<АR!��i���:S/A�ez���"O4 P��
�n}:���QlN�qP"O^�RE�"��85HEZ�
�H�"O�kń*�h�i�b)��`�"O���b� Uci���E���1"O�1àʧP����f��~Hr��$"O�*'&ιD �0K��O�$6XP�"O�XB�O	Cr�x[E&� d"OL"�F�Q&4�	�$C�[X����"O�LY�%\�G �X; ��� 1$�Q"O,Hi�=�X�0P�]"��(�"OpHp��,"���Uf9@L(Y"O�� ��V�/�F�#1c�:jM����"O��z��P�L��;S:D�HU"O��1 .ڦF�^�0�`M<12((�"Ox����6Ng�9:nǵ''�tç"OҰ�2��[�T#t��>�,BV"OLy���M!P%�q��Q�@0"O\BEnԉ,
.[�A�(z�\V"O�(�����D;fi��/��A� "ON|�����Z�A(U�p��1W"O����F�%�<���K�1~�0�Q"O��:2�Wk�;T�B|�¥"O����$*|��H�+�E8��"OHeH:x����CI$�"O���b◄E�yb�GL6P���"O4ɓ� �i�e�L0'#~�Sj�<�t�CW��gH4K�=���WI�<I�B�h`d,1bL�5U ���&��<	�Q9h\�)T1o�M�ס�a�<�1F�)��$5�ES��b�<9�"�$,bfb���Ҙa��Z�<�C8}��Q��o�xؖ���[�<�f�Ee�-��Y,�H�F��Q�<y�%��:�|���%	�m���lA�<QpE̫'	F@��Nf.��vE[|�<�����9��M�JU�8R�"e�<aFւYa�Y���
ci���LH�<���D���Aėt��)GE�<)!`�&�U0"H?c���
 @�<Ĕ0u��l��A ;?-����BA�<a��Pe|��7��*(֦���}�<�h�]��B�E	�C���� G
{�<i���u�>)��!��4��S�~�<� ��cѯ9~d\�w��3,�,��!"O5��,5Ό��'�����"OܤӧGV28�\p1��'s��p�"O<uڅōT�����@+&���X�"O2�Y�

�j����;%���#"O��%�d� ]2�f�:pG 4hT"O+���}���/JD�B����Vq�<���(
P��*�V�18!-�e�<��哤)i��1*��!",Ap�c�<I �A��am���k^_�<� �0�D��G�.tծR_�<��l�9��Ჰ
��U�
�s�<�4�	i+d���&M�i����̊a�<�b����a:/�=@�J�A�]_�<1d(ҟK�X)ˣ�
95�$Q����X�<����-�����KISN���F�U�<��N�nh��
$�Z�"��'�L�<I�7A;�ـׯ�*a׮���!�C�<�"�ȯI\0��[�n]�;��V�<q$�_ ���
��"��ѳb�V�<��d[�0\l	��!Z�Z��AcF_P�<I&N������Z�0S��E�<	CCU�+�
$�d���]&��IN�<I(O�k����"o`đ��P�<���H7F����7���yFd�T�<Y���0-�\�猔�6 2i�V�<�P˔�Vy�Ԡ��V�F�9A���Q�<�)Ar��a��#	8�&}�"�MN�<	���Y�HAB!�@ 9$����g�<�U�UMP�@��J�e����I�c�<)�b�`��EZ�?p(�TJ�[?I0+T���>Q��	U�t��	�	��-�W�ZQ��H��L~���	�9 ���c��|B��z��� ;o�C�I7 ���	�ː�Y��ҥ*�#|�c��"W%��h׎(G������^�js�݀���J���yR۸SLZ��p?}�|$Ⴋ	!_��CuDEk�ɉ�H��	�3�N8(��E������� �PB�!�BYkâB�X���x�I�<,6-��nbNxXf�7�Ox��c���$Kbk�t0<0JW�'Jb�7�F�D�����(,\��/ңH4� {�D�0�!�KuT � �Ӻ0�xd(Xy�Oqa�{w*�~J�UC��EA7�[8) �+��@^�<�`N�(ͪ�Pd�@9D�5kS�U0��XӢ,:�ĕq���D�cؑ��ۿ81�lCĊU6�!��Q��yK��U�L�8hih�7���R�lâ�R��'�8��3L� zl����=A�i��~���+��F?!��X�B�pJ�a�=ظ�!��Ij�<�6 �&��0���,�`�Y�EK_�'X������ݜ��d�`�jY[��΅	2pB�	cA�Ls���;vaF�%-�z�tB�I�R�BS��/L�@irß�UzB�I�\nT� ��i���#�\"g�rC�I�n�����!<K�!"oڡf"XC�I�|_�$`���`�j��Z	�~B�Ig:\ب�H�<�|$DNL�WM�C�I�9Шa�gG�
�&,�4囬P�!��K�N�<d*��p]I�';D�!��\;�J�CӤ$n5t��Gѣ-�!�/Q2Px���)U/��#�FI3�!�D��2�=Z�"9M���`�b��O�!�<���cD+�-�n��#Ӄ�!�DG ����Ł�qC-ᓢ��!�;?�����D۲�&�!�-��"t�,�,��H+�!�� b0ce�Fp�5�6���j�#�"OX�Z�kĊ&��d��B�X.jq؃"O.|�m�а�l��P�r9��"O�H��┷},�I
�+��S��"O����N�>V�1�$jC�"��q�P"O*<xwm�+i�����^��P��"O�9z -)� $����0K�̼(G"O�QpD��1�����\,�>�m*D���DGS&��	J�F�t]Sp�!D���`��m�r`jv/�q��E�� 3D�H�cN	XD=p�-�*�m0 .D���Ҩ"+zٛw� 8�N���-D�l�ޞ7p���k-\Dy�v((D������V
"m�/h�v��S�)D��r��ҫL�p�y�I�+��6'%D�x7.¶H�(əU�ǫ2�B!D�(;Wa��p-��h�E#�t�/?D��aҬ^����	�T"�퉧/<D����P0qU�(1��1�:D����-�VL ��"?4�ע;D�	�!�7c�~�i�J� ���#�**D��#����,+j@0��F�3ڈ�$c*D���w%ʤ6������g~���C�-D���TiJ$���`N�!�� ��<D��{�j�B��R��ߡT���i;D�0�g�@: ���� ^���1b$D�8c����}^���Qaѕ#%b�"�/"D�ЖÑ�/�����HX�1N7D��*`%J�;+��pbj��(���4D�(��B%$�^�q �G��};Ќ5D�|����~�f	YQE��8Y�eh0D��Y�$R�!Nn�jA$ЈV�q��0D��h�A$/���E��D����7�,D�Ly�K?#�<%@"N)X��_a!�d�H�b�RB�8!(�i(b�;$I!�d΢^0M0���W���x%�
5!�D�)��<���»W� �;��\���$ʠ>��1��kp(��G��y2��F�FY�墓_�@ࠤ)Ď�y�W�&�L��'�Y P���W�yB픣'�(2�8[*<���Y��yiS�&�ָcPe�<&��±U �MC����w��	a�rhKݴwV���m	"*x	�c	�{�8�pw�Ig8�,��f��m	*�Q!�N�D6�0�&h$D���
5)zU���?/����)�y�^,NŘ�2/<�tz��=�y�n?��p�="�"<���y�h�9H�dX�n^��<��@��/��O���OO�Ep@�δ��0� f�������3ʓ�����@c��C�<�pWŃUrO*y���ɐ�}8����E�n�4��������8\-Q�"}���v����%�Z�vU���O��Ѯ6�S�OӬu���K� %��2�EJ�B.]�'�:��%�a�$	�S�@4⒅��Vuj��p엽�?9u*�.X�lbE�O�ћ�B���?��F ��Xٺ�(T�R�rjl�Mw��^%V� ��?��t�N1$l�b��Vڡ+g��$a�@;�S�O�	���\#YF�L���am��0۴a���<E�tgP�jܤ�����%*��-vQ�\�
ç;^��P�j�������U�F<�>y�1���ɣs����F�HJ��� � ��O.Ọ}�I��0���E=HK~�;!G�3=RC�	q>��	U��Tr��DG�w�dB�I�o�>h�V�:{�x�kfƏ�.�B䉆,p�pUEU�#m
9jo�`�B�5�.�*Rƚ�^�+eEL��R��d=�� �ڷ�ǐGr�j!ݶX�l�C	_*}Z~��V�i���v�*��I�����
���"H1`�R�KR�y��Z(v*P�x��� t�T Y����y҅�
d�(�i��ޛj�����0�y�$�R���1aY,q��ر�h�#�y"�[%3�Q��d�2j��P�#��yR�Ʌo%rm@eECe 쨻�D�y�*�-hAz$��0a>`-�D��y"��$ft���dO�L�jŹ�&�$�y��N�*��}d�^�?�h1�V���y�I\�%^�y���8�L��%�!�y⏏.r��tgA�nHäKN��yB+��w��ͮp�4ف�h٥(xy�ȓU/
��tl�%T8;T�ݡA�$��ȓ:D��CnS4����	?�6}�ȓGt�|S�e���5�[�O8���{!�t1��Ǵ*� �ҧ�� 7`���^f��G�KBiʗ Om�(�ȓ��=��R�-�E
�H�MWޱ��py�E���Z�t���#�A��8	�ݨ�恡1΀�Ɗ�
n!֜��?�d�83��8v�l��W->#�VT�ȓQ�Ls&��/&�\��@�Y�&�ȓ=�\���J
�j��FX�=�ȓMip�6)��\�bu�[�q�ȓW(#S͛�삱��?J�.P��4��|�e�՘&���ԇ=~�f��ȓ/D� %M�J��q���@7s���ȓ.�!#$��,NA�@��
pȅȓ}��xS��8\���Y�	�p�ȓy��<�gD�.�ҡ�1�Ǽ	x���~y�{FB�:���!b�:t�݄ȓ'����A�$%	�K���ff|�ȓ/��iVU�3؄r��;E��Y��_z���!��R~���r�C�\���zN��u/BTd0��)2��R�$��k�-L~�z�ƁE|็�H��Y�r�G:��kU�:/�������JEa  !�	P!
�E��a���5Z�e� j�hD6wZ��`ڤ�����H����e�nu䡆ȓR��)bא���-(S}�0���A�H�/P��(�R�$_�܅ȓZ�h����8��\2�E�Z$�H��>����� ؚHb�V�G$m�ȓ+F�� ���.P��`r��.;��R�2�a��7dkD"C�ʢ�T���F��9J�KT�i���9��˸<�C�/��p#�Ĕ(Ӭ4��:s��B��:Q��C9W�M؂�]0XG�B�I�*g2E̙�%:1=��MqPG,D��k����G�F��DmMcR�H��+D���Ti��X�V4�ą%)��D�+D��Sp$��p��5���ӹY��*�+5D�t�pbAL��[�g�����1D�x�b�W�KN� L���x,J��+D�칖���3UH��4���L�e���+D���q�K�>Z���
��
y���+D�����w�1hBi�ZT����%D�L����jh�8;�剃E��l�ì%D�p��Js� Kg�	�%�Ģs!�$\�%c���H�} 0�XBNO�Y!�
�$0��cת�{ᖍ�/K!�DܫZ�E"4C�y|m2 �Љ|O!�� �*R/?,�8�.�W��p��"O��QW�C�	�xd���c��yP5"O��� L��dQX��1��Ic"O��:ƨ	�zq�h�!�$M'h�<���[�p50�U��C(�<)�ت)n(�E��2�w�<�F*/�T��S���0j|���q�<�%�B�0TaEI��M�����p�<��o��]�����D�I��1���C�<���\6��@�����'�HV�<�aBq,}��)c�R��&K�<1��M~4���SAZ�j_���s!�K�<i��ɗ(�:ٳfu��@1��C�<-��Ũ7�KF�t��u�1�*��ȓN@�;��I��`���(�9��H�0Q�`�\� �H!�^s<��ȓ{+��:���_v��P��|[0��	��Eh�i3m��y7ǜ��8��X��!�`%Ob���Qf�m����j��[�a �a����w�T0���t��\S��% 4[ ���'��8�ȓP���,�	��d���Q�����}2���U?[��7fW�����ȓ6̋�l��J_ t1#mJ�~�X�ȓ	G�ɓģK��u�B8 6����j0���K!-#���o�$�ȓO[8��U �{8��a�
pr���ȓ"�,���E� ���î���g���GM`�&��í@(F�h�ȓ0�l �q�[�7�P
%� s����\�<E[��M�8�^P�Sd�~��P��H��h;��G�!�x� ,@B�~��IC��O�+��|��%�Aw�u�ȓ^�Wd�3}S�@�e����u�<	���g���"�= v�12!�d^����J!�k�*,�L܊{�!�L�y!�L�c�Z�p���f�[�8�!� (���LIF2b�C&��!�;%7rY+�g� �-9F�ޟ�!��19T��
,i��&k�:z�!�ɣX��A*�)�.0����#�W|!��9��-z�ã	�
���޹h}!�D�:
���FJ�.�~L{��^a!�G��"�ABIHuN�c�LO!�$E�@ց�uV��iK��DC!�D�?y�"m��E�Ef�`���^
2!�D��^E��:����p|t���M*E!�D̓cu����I/%�ɸ
P R!�Q������%���`6I��5W!�d	%'zBhz�G\-z��`�� PP!�d�b�F�x�h�C-����)m!��R��=Yr�Y6�yv��.R!�D	Q�ph(� G�X�B}��$�!�$�*%�8b3j�}r䝒�*�`�!���0Mu�`�z
z��F�0 �!��&Y��TML�@��e�A~V!����hp��!Z� 1'�� Q!�D��p��ԃ�&W<4�,�!�#Y0!���&y�(�a��5�1�LR<!򄏕��A��@	�T�@�ppe��
;!�d�	G��$��������B)!��<�&�Af�
b��:��!�dǮBZ�Tp���'O�j|�$H�!�$G�t�ڸ襪��8��rh*7!!��  �@uE�(��aS
3\�x��W"OsK�)X�`T�!!�(��"O�p3#l`-F�I�Rr���"O�t����$��L�b�n
j��4"O���D 3�����>o
X�v"OT��pL"{�d����$Z�l"Opa2��;�ڔ'A��uR Y�"OM�3�+<�dy� #�48D�8��"O�u��DѸKr�z��р%��""O�Hq-шe�
�D.�&@r�I��"O <��M��,H�<q��H��$/�SⓂ�r��5�I��4ْ.=JgC䉧��9�F��O�  t�C���B��z�
}x�ɗD����NC�+�nB� E!�	�7�����d��@ 5��C䉵!�6����L (��0��_;PHC�7ql��C�R8Ȩ; � LnC�1���pwm�!��\:��Z�m��C�9��� �T�tyǚ%<\|C䉶bj�&��&|�a�Pb�"˜B�I�:*`�3��)�����B��B�	�]��� +G�B�ܐ�lۤQ� C�I�)��Yhpɛ�G���d��>|:.C�	!XeV����5h��Q��n~C�	�3D&!Z�$ԲYw�Ic�G�r��B�ɮSkx��nŲ7�|h�E˂�rB�I��v�[��Өg(�;���9hC�I�0M"��������\<j�B��X8�ۏ"�H�{�.���ZB��\�&D˷�3:t������C�	�a�ڕQ�${��)�#ܒKB�C��4'�H���k�;}=�ɨ�[�.`�C���V9)!#S�P?���aN�P�B�	�v
�,��G�R��yd
=PB䉁��u�S��U���"J�4m��C�Ida����R�=_��9#`�c�B�I$
JxPT�EVN��ׂʺ0�dB�ɜ����v�G7T2���kS�,�8B�ɎƔ�H#DΉk[�l�r��6y�B�	�2r��c! (@�h��ѾkB�	�<��0J��e�N�K���%��C䉣x�X!�FM�:>Z�`����+H�B䉶`��sԍ<�vX8�f�hB�	�/��� MC
�8���D�v�RB�I4�<8��ǈ>�0�"JC�/&B�	�s��%�Ц�n?b�(F/�38F�C�ɜNI@5�A<{�͕h�nC�I�v���sp�ۢ���q6ʓ�KB�,'��ı�D"�`y꒸"C䉖 �"��*2~ ��d�O��^C�I*~R����	[�"�PՄL�Cq&C䉓4"|� .m��(�Fo��p�C䉤,_��ك�����QfR�^C��6k=��P�BΗw�~u�B�ϯ9�FB�	.�0л�B�=@�["��$B<B�		dR�:�!D/T���[@!$_)�C�ɹs2� �?(�x�Bb�_5�C�"\�"�h K��/�~pC�Ģ?��C�	8F.0��I�V�x����;��C䉚�ZlpB� M2�m�$`�C�I"Q�T��+��4Hէ^%�C��'���#K�(�J����C�I��t�� 暡;ΰ$sr�!O��C䉅w�LcЫمj�t��l���C�)� �����|��@h#h�-y�.[@"O��4�ωv�,��cML�x�@�3"O؍yUȐu8�Y�->l�$��"O �0���tbH�ˉ<f��}ɢ"Ofh�hZ5$8�Y3g��@āX�"O�b�.M^H�p'�
<
�P�d"O���w   ��   X  Q  �  3   c,  8  tC  �M  pW  �a  Yk  8u  �~  ·  [�  �  T�  ׭  X�  �  &�  g�  ��  ��  2�  s�  ��  ��  H�  ��  ��  * � l  �  @) �1 �7 m@ WG �N �T 5[ �`  Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�� |d��"O
`�(�;���8���-0��1%"Oj4��ND^[��"3/9�0|H�"OB���H��*�ʞRy=a"O�味V�!X��!&F�:J�$���"O,��a
���C�Ą�M�"O,$3%o�-���p���+Ն�:1"O��ݢ1����`���y14]2��i�<�6��{_���c�H�`�fX�$Kn�<��A̼VI�xR[�)�Ć�pඤ�ȓA5��('nߡ4�� �)˩%� ���,��r�؊b#`T�eT09���ȓ!�b��g��}�8�F��-? �ȓ
K|m�ș�VṔ���2�%�ȓ"R�X�j�4JN�1�˘X�i����̹	_�jZ��1!g��zܶ��ȓgil,*�J�
j�Ne��i�J%b���f	�(U��:���G��$Y^م�~r�� S�%T"���k\�jx�ȓ|4�1�îJb��@ӵ�ݩn�V��/[`�"�v4�R�!ʎ<��M�ȓ`:��z�ؚh�J�Z��$HY:	��H��p�m�C1��!��B:��0��EnjZA V;9����J[
2���	��4'J�EA�IVW&��~�(aZ��ӹ�>� o�Y�|�ȓ�f�A�
Ο7�H��M�$�����mޠP����/���ANXo*�ȓTv�����{ ��-7�*h��I��sB�8�8���3����ȓNe*M�悡;������X�o��!�ȓ'lj�#F�m�+R&;�|��2)n�C��0S4���T:
b���:�0!��e֊��)��ͷV��,�ȓ0�&�8#���� ع�L�����;�P�AFdD��,w�6d&�ԅ�I#P�����L]D9  i^�D d�����<��Ë�n%N��%�_0��hK1M����<�S�O���˂W
�0�.�B������h��iX�ܥ	$�t�F(ȿ/a�5�$��<��)6�O�I�!�$dhJS���J�dݡ��'}���[P@�K� ��a��4*ue���yb`�?R�@R�T4D\��*���ĕ RpX���"�Y8�A�؀c<�&��HC�+x�ő���w[0I���]�]�B䉽��ḇ��~F�@ Ϝ�{�*�>Y����./Y�L)∗�.�+NX�b!�$R�A!�ݐ�A�Ao��a1,�!�D�  u�A��7Dعc��!�Ď��ͻtʇ�&8��kߩr�����h��Ė+1���&A0�"�C�R?=j��e������]	<?���O��zd�aE0��W؞x8Ѐ�L|I�Q�M'?�+�X��ϓ&YȢ&�]�d/&��`��W�Dz��7O�`xVH$��"�M��Tҩ�"OxhPQ�^�1�hI�ᯍ�~嶼�W�G�I7��=�6i�QĴS��3K˞�Fʛ�HE{*�2����<��1ib1��E�&!h#�0v�4�ȓhK�B�4�"����{9J⯓���OPdF���En�lZ�mHQ�t8�X���>�OL�9c�W�7@N���:���!G��P8����P�*���WN�=���3o;�Ho:� "��� �};� !*L;��ܘW"O�U
�g�{'�9��ޙ=�T�Y��5�S��yR�Υ[��a  M�8x���G��y¥�

Rd�(k�d�� ��y��	T�'l�����g>��=0�4���'���А�ԫTp4(+r	E.H��'�vUc��DkT��D�06j>���'.��R�G�W�j���6�$�K�H��	�����R��h,���`�|�����<i�'��$Q%)�X�j�g�?���yd%OA;ɄēZ߰I�Տ0�|��F|��Dx��)Ҁ$�:<J��h�*V�Dq�L�'CQ?ͩ3`)h�j��Lz0r#-%D��Q����Qi����o�L1�J#D���v��;:�
�)7JO�~-��U=D��{��fĀiiJbɰ�R�e8�DΔ��=��O?i lP�۩eM.�Si�F�<AG�m���Ȃ��	QZ� �=��>1+O��H�����RG$ƫ[�(j�"O�kD�X� @��"4Ƃ�t����I�����]jǠ��B�V`b"�%Y�2lԘx�>O.��=�~5�GB9�!�f*�)H)�3�Yt?���)�'5�z�{&)8`��L�% ^-P)�>���)�T�A
�n�)��UW�r(�¯���y��'?�}R�R�g�t���Y& 6Y[*35�2��5�g?Qd��$� ���ގt�l���g���hN>ف��(X�1��E�P�L�a�D&[�6�d�n���+e	#Hh�42d��|�Y�ďa�<���J�uT8�@���&攭�p���E{���])jq6�Q�V�4	ip���<��}����W9"i�c"K>�"�6�K��y�'� h����?�����d�3c9d�S�'���p=�`$��9�|$1w�ͤ8�F�2`�iH<a7ǓnJ0���3��P�C	.R�����ç�����2��.��<���Ʉژ'0�)�w�,��@M��B9���Ŭ�M���Q�'&X��oE�.����#�`ji۴�Px�GK��*5h��y~�����T���d@A�'U1Oظ�c��>N�X�����	U�Q�w"Od��3�=|[�lp"�k�&|"2"O0��I��X�R�3^0@��W��J�������4�|S���,�4�͓
|!�ߦ{:�eI��ֶeWʑX��Exa�D<�S�O������>~|�8�e �a�$���'cs�g�����;X��lZ�'%|գ`A��a��{d$[�e���
���ZB�0@�/_�nq����%�l���iѰ\ud��j,$Ȁ¨� `�p,�' �IQ�)�'x�N�Y�M��5�4 ��QIƀ=��}��PD׊b�y�5�
�g'x�ȓU4.� �E	XIb�%�3���ȓU2�x'K��^��ehwB�mU&��Ɠ{��Ѱ�<q^HpA��(&���s�'붵 ��&:���E��R�p��'�h�`�i�w�<l�%g�;ED����'�B]{�蜋d�Łլ�?Q�=J
���?f5!3!�(3x�� �-T���ȓ2�>�����1v�Z� 	+J[nh��hO�>��J.=Q���t�]�5��G&2D������N��Us�j���i��%�=�O mI6��3ɴiP� ה���k0"O���D�?i�Uc���Y1�]��"O�3�)j���K4�ɱ3�!{W���Is~r������!ɝ	�NY3�"Ȩ2�>�0�*D�� 81�ɥt�<%
C��3�ap �'�ў"~%&B�z� �%�
~�d�0*р�p?Y�O\���ԓR�0��M:*�h��"O丰�a��E�ǁHXѢ"O�qw��f5�p��J�8e�Pj�"O>��e�q�M�+����m�f�'x�?m�OT�r($�1�T0����L3D���EF>��a���r`��
І+D�T� Z���*PS ����-D���t'�)���Ӏ�5��x�g-,D����m}�������v�%+��y"퓊'q�}���B?g�كœe^�C�	���a{�'T�
W+�(U��x��	�<)���H�	�f=�5�[�3^�Uhq��!��C�t��!5�)��Y��eT%�<����eڑ>�AX�\�!��-���8��D�:4(Յ�["��u���:X(��	+�l���?�q��tыeHZ�9�lݙ"" T�'�?A�� �o&.ժ��'y|Q�)D�(���q���G��l��15�'D��!S�W�Sy0��sˉ 7	����g0D�������!j���h&�ʣ�8��ȟPq3aIHL�b�"ԫp���`"Ob-���סvG�i4+�
R����"O�qb�t�L쨒䁯-��}�6"O����K���G���1���[���|���(s4���IA�yr��4ø�p=a�O��I6ZR8Xv�8s�|@�c��=�B��1R�n�rE[�vך��l�S�^">��j�>!�d�]�?�
%��W6h=�EH��"D�x�����	\��ř�e1�&?D�4��M�?)�9�g����Q��!D��E&����h��u4�P8GM$D�<3$f��?����*	x@����!D��ҁ�E7�J�@��������>D�hP��ŇGp�	qCe�Ib17D��i�E3*�V*���$�^���7D���w㜰v{D�( m��;3�1�%�5D�P�tM��=J��Jp�r�x�;qk4D���u���(����%̛IYre�aH2D��Ɂ�_-K�Y��
�(2��S$+D������TbtH8B͑(� `P$D�th�'�Y���1�C �f���j$e7D�ܨ�P$-�E@���$B\���ҍ/D����t|������_�x) c.D�����D��-s&�`����K2D��9#�--J���5�>��`��3D�,ZF���W�Pu�W@�1NT��H2D�,$L�?\���b)�N58G�/D�X�3&d���Ç�X����B&-D������"9�(���1�
}C�
,D��� �L��m���S-2����-D�P��_�{̭9�P�Y�	g�8D�$2�f1������϶���Kq�7D�T�To��-�����Ȧ���c�6D�XS�䎓�t���-;�%ʳ�3D�<�r��4�iA��̲	J1�6D�\�&≊=ӆ����3$bf���4D�p��7gr��PT��1�(#f�0D��` ׊e:��tH�N�TH�t*"D�Dy������d��0n�4�2.D��V"��x�
D�0U*ȩ�4!*D�xy@Ɏ�VP��Jr��vp��`�
(D���R��@	��q H�}N-:$$D�� ��hB�F.'��%H�)���CA"Ov�8�!I�@�H+�m�(r��$@T"O�<��.�T��$�6e"ԣ�"On V�05T�����?M�KB"O*d+�O�}J�Չ�莓G6ⴋ�'�2�'�B�'���'���'xr�'�d��c�j)|�sp���xz�au�'B2�'���'���'���'���'U�(fl�e���C�\�w"0a!�'
��'��'��'K�'�B�'��4��j��~���8&��P3�'���'��'���'�Zƛ�'-��N�#��)��(o��4�)�F��'���'���'���'���'6���;jV�Z��_�h��|(�-,��'�R�'o��'V"�'G��'���B,��%9㦉�N`��B�΍#iC��'�2�'���'�b�' b�'mB�ߡr�R��
�4)���hG�]��'�r�'��'�"�'��'��
G'�p�BV��.`L�r��J3��'�r�'���'���'��5�4<h<)U1 ƑÒD1k�B�A��?9��?���?-�M��?����?1U�CI�eJ�=OD��Ǆ��?1��?����?1���?!��?!���?�T �i$F$8&��:1Z��x���:�?)���?���?����?��?����?Aw�|��� U1�� CL9�?y��?����?���?���n���'=�
�"c�b)P�Qw�9�pɃ9<�˓�?	.O1��I,�M�c�G�t	�|a'�֜^����T�߲#V���'Ղ7�3�i>�ɡ�M�0��@F�  �Mp��")FoқF�'x�iQ��/#"j�� E';=�&�9`�g����e�V&�L��<�����%�'v�E�c��e��k�#Km�Xku�iF́y����Ԧ��:-Nl�ס�3ܪ�X�ɐ�����ڴm��f5O��Ş���4�y�
?���s¨�<�N�;�L���yjɕ ��#�+D�C�ў��D	���#:$��Hc��8�$�i���'0�' 6- D1O�4��m�vsB�#D�ٜj�4�c�!/��<��d_ʦ���4�y�\�H�
�r$dy�S2`s���<?�ͥCc�y0�#�@̧i��\w&�d�3|��$s���g���0��������O?�ɥt���� ���"�>�+��D�4���	.�M�QWg~��z�r��S�����s �9�l�Ϡ�	��M�w�i}�$��wg�F��\9���P]
0(�0��8B@^�Ĝ�O�%Y��-%�����\�M#���?q���?�"!{���2�ݒ{±rq`ʫ���֦��5i˟�������M��'�@�ґ+�3!��->]D�U�ʳ>�¹i�6H~�i>����?5� m˧;UJ4qG���ZL(��#�61��=���Cy��ZD�xZ��N`L�'A剙*c2(�`�j�^�t ӑ_����ǟ���͟|�i>�'w�7m�c���d�.a|�`- >�-�)��Q_�L�U�?A�Y�0�޴<��v"g�@��IA��y@"�[1�9q��˨c�
U�D:OD��)_vTQQʒ�}AF˓���N�Ha�9x����T�lEpp���?Q4�H8v��|���նn�D ��I,��D�O*�n%<9j�'ou�ƙ|/U?e��E�V��^vْ��� N�VOl-n��Mϧ�8�*��EV~"-U=l6@����L�@%��EWJ�`X�h�P�|Z�P�IƟ��I��0���ң4�Tqdc^�(�>��:�,�D�O�^���ɞM�b�'��_>8D&B �*1�����n4PCPb'?!R�P��4`��E �4�J�)�<u��hT���-E|� �X8?�ͳԀ�#�"����<��M଺`o���I�M�!� �|'�����7s�A���i��V&Ă*�f�⢦@)4����K�HUB\�R�'k�n�n�\p�O*�lڢ&=HlQ���3\V�a�$܍9b�`8ڴ&ɛ��/Z4!�'K�'"^T\�G��p{��{?�)s��9���rfj�K��sy�'�@ �&�m��8B��բiӤԛB�iӲ�;���OV���O~�?�b���6O�.!k�њ��C+jm[��_��&Hl�b�'��S�?���R 8���u��H���c $U��m6d�J���N|��8.Г���H�X�O�ʓ�?9�b���;��ä;X�����#�R[���?���?�+Odlm'y�B���ݟ �ɸV���b���$���#|�j��?!g\���4I:��+�K�?F(
��F	*\�eI@@و+�$�Of��⤒	c����<��'4ȹY$��3�?A��#S��P5c�3�]��?���?���?ٍ���O��X�'��Xpp�)x;�h���O l� �0-�'�6 �iމ3��gؖ�"�ЉT}f|b��~�B޴&�fgu��m�3݁>��D�O��"��\��@�Kig\ ��hPr��4(1
��O�˓�?���?!��?��Dl8�W�Ԣ{�>��'�#i�@�.Ol�o$11�������	|�s����� v"2��@��3@�|���V'����Ʀ9`ش׉��t�OL�t�F�{���l�w����W��5l,��E߄k��ə
R��#`E�~F�5'��'A�t�u�'�n�Aw�@�a�4ّG�'�B�'�����Y�L�4���� άA@�	:�R��e��03��6z��'��'��=`�f
`�lڮk�d�Cs��re� f���%��4����̟PiL�b��s#�syb�O�� X�*� >@�P�(p%0c�v20<O����O����O����O��?q�qi�:���aT"-~=�3�����؟شe��d�.O�nS�	7 )���0I�1XX1 b$���`H<a��i�$6����}qV�[,,l���O���E��m��*�����"�@�bf�j�N*V�~�Ob���'�b8CGo��k�d`�]�=��+���������}y��'���!@����C����,�,8(N�j)��<�M;f�i�O���N��$M�?����L���O�-H�`4)�ԟ����:��=Qy�x�I>	fk�$eB49Zf%�E��@1.���oZ�`��埜�)�wy~�`�à�O�Y�N���;P!2,#gH�6�����OHoG�7��	 �MSB�\�^TЭ���\���������s���j��i*�`��p��D�O,Y!�K�7b-v��c�<	�- �vq���6( �0��	�<�)Of�D�Op�d�O����O�˧/��! T"
���W�[��0�кi`�I3d�'���'[��y��s���[�����ҠVR�hcb*�+Hq�Dm� �M��x�O���O�j@�e�$�y��-,�p관ق..~1Q��%�y�`8D���(�"W	�'��IƟl�ɞ4��E�U�
�h0R�E}gT��	��(������'��7M�/l;����O~��ǁ^��ܸ`�4��99�ԧt� �Of�lZ7�M�ǔx�HYv�C):Vq�gM��y��'�0�2�Eƥ>4��B�X�l��3�
�PS��,�P+��0���u��M�]`�	�����ߟ�Iq�O���M�:�l�-M����w�B��rh� ��Ol��Ԧ��?�;J P�#���p���5{^d�\<��#tӆll��4���Y!~���I�؈��� �&J(\؅�J�A���jBP�%4�mj�E�	iyR�'8R�'�B�'@2jM�A{�`F�( ��5L�01��	ҢŖ�L�����OJ��!���Odh�%`#~�p��7~E�JY}��d��YoZ����|��������\p�)��"�TA�@����S�8��d�b^u�g�� W�ޓO\�;t��hR��P�朐� ��?���?���|�(O~�lZe��	7%H�jC�aD�P"MY�/Ԣy����M�Z��	��M�b�i֐6��6���	�E��/1���4S103���P��d�OLS5�
'���ٗ�<A��׿kuIR(^=�J��}9Z��W@�<����?��?����?���\��mH~�Ƞ�b�x�S���?���>n��aH�	��M�K>���F<\M*��'њf8�r!��-j�'6-�զ��F;΄���q���	4?Ʃ���)C�� �/	;��ȥG�	�Pd�'�¹�zL!𫀚k�\: �G1s���)��Rx7Bʪ� Ԑ��(W�]���E#~�:xҒ�HO� 1֚!s��Ct,�<�P4Qt
�q�c�2]��tÀ��P�`ȣ$��n`�G$�[[�`���<KQP����GyO���E�K�!��T��V0�%H�Jx������6_y M"a��:��$���� :dh@�?$�B|BS�C�$��ċ�7H����� :�����
b����50�c#
j �KFG,b����C��*�e1��\�_"� ���3� k��'jb�'�B�Ò�(��;X��Š�!�9GF�p�&���O��£
���'!o@P�6D%� @��m�?i�QoZHy�`O�i��'%R�'��4^�֘	Z:�٤o��4��h���k\6m�O���\���b?A�1D�!�&���ʑa�cӞ� ���O��D�O��d��Z˓�?9�9B\8�jʹ�F��J�>&�&��t�i�\P�7����A��N�!�����"��Fb4#!�W.�M����?y��8Ob͊�P��'�"�Ov�(&��R���C�K"O!�Z��iM�'��C5 !�)�O����O���0���NVb��slΉ*�tI+VO����I��A�'�B�'�|Zc�� !�d�V�i�q��-x)�`�OT��T�;��O���On�:/H����T����	(d霈CR�؍���O��$�OB�O���ON����>9�+��p^��A�p0��O��d�O��D�<)�a�9����M�����B��LA�$��@	�M���?9���䓜?1���W��`�vG_�:ء�C��Q킑1N�>Q��?I������E{N�'�?����pA��yhB��w|��'B�'��':���'!�/$���W+^+nT��m�/ƪ�m����My�%B	��̟8�I�?ɲ��&K�����(:� ��b�N��ē�?���X0�`ʌ��,��5	)M�$A�f�qP���i�剖�8���ӟ���矘�`yZc2NUHT#�7p~"e(�F�x�����4�?���?�PY���d�*U"$�K���S��X�Ę�M�ҀI'J��'!��'���.)�4�kl��p�2� k��,���2$\t����Ȉj/"�'R��'��4P>�Q���SLڱ%�DQ�f',u��q��ib��'��%�8>0O���O�dL1I�^PKt�ږm���F�!ȼmn��P���<�'.����9O���O�{�\P�q�'n�i�ǈI�j�%z���ئ��Ɍ~���O<�'�?1����$��6*e� �
hp��˳�
�z9m�x �j�� &�`�I�$�'a|m!C�,=.�z��?xZ͢%JJ�5ܨO��d�O���<���?�6dE�J����	�����G�<:Iޙ����D�OL��O�ʓ3f��4��d�� E�e�8�������qp7Q� �	ߟ$��{y��'}"�ϛ�B�=���c5E�j��)�iT�T��?����?i.OL5� @�Y�ӯ;��͊�eۇ�]QR�ƶoL��4�?�����O�������ľ|�� ������=4�� ���i���'��ɡ\#H��K|"����1W��[r�A3>��yrc&ֈ)�,�'��'�xH��' �O��ժ#򝐷I)=��ձ�"!A�fT�<*�J�M[T?����?A��O�9��${+8�iؔf>��òi�r�'w�) �'WX��?�'��i�"���+Y{�(-I��3��ش/�����?��?����?���ɟ�1��%�@eھ� Ex�ɀ��M[�LW:[�V��<E��d��xL9wF� @�f�X����t��7�O����OL1!fζ<�O��0��uH�2����DE���r1O�i���}짒?a�'�ȝ8Q	Q�y�����+Y��4�?I� 8���e����ĉ����0e
�=�t��@AҐ/���'��zV�����'�R_�H�	 L���"�
>bMsw������ŉ�ky��'r���OL��E3Xlɶ�Q�Z�@Ӆf�6�Hd�0`)$1O��$�<1���P*�O����|�jQ��J"pj9jܴ�?�����'\B�'����GN�M�ff�^�e{�	U��e��  c}b�'���'�	?� ��K|:E`U r>��q�ٵ"x�����;��V�'6BT���	i���'V�)���,$
Iw-�A�-�#�M����?i.O� 6-�p�S�H�s��[G!#|�X��7xZ`�郧1�$�<����?qH~�Ӻ�v�6 z��ʠ&
; ����a�TŦ��'����G
v��U�OC�OLf�%lD83$��>��ACb�P���o�ȟP�I����1���<Q)���)�0eʐ��G(�*��CF��M�ц�1<��v�' ��'��i3�4��)��$tBKcA�]'$�m����k���ß���$���?���y��'�.�@���XY6 �~��=2�|Ӱ���O ��E�p	��'��۟L�Ir�tɂ�X�u�TEb��!I$���4�?!��?��&L�i��3?q��?�YP� ���+K�	H�(��1?�6�' >�0WN!�4�����OH˓P���Y�ρ�Fn���U�NV0�=;6�i	���rX���	��x����ɝ�Hhj��G�l�l��0%�ݺPo��M���?Q��?��\?E�'�2��2�Tٰ%�^�`���F%�/K���ʛ';��'��'��S>)a�-S	�M��
R�-���Ƥ��K�t1t� yn���'�b�'�2�'R�����!�d>�X�}4��φv�t���E�:5B�6��O����O6�d�U�$n��qSr7��O����&U����*˒E�<2'�v���l�۟$�	џX�'n�����>5`	�}�,3ܕP܉�2.�����Iɟ�����ܹь���M��?!����L�!9M�G�#Z�|tj�Dȑ8�&�'��	˟\�Wi`>)��my��MS倏Zf��FJفd����p������'gd�R��f�\���O�d�H�ԧu�♸E�ƹ�҃�4qI"!J��ӧ�M���?���<����?��Ov'�[{_ZU���	�Ddr޴VW�A�V�ig�'���O"�����8u��[sߟM�2�eɬ_to�������(�'��|��V=���0�_����νV��D�UdӘ���O��䊳8�Z��'��͟��'p|�Y�(�l�4�q,D�	�v|�>���a̓�?)���?�!gY*6���˴�ؒe<�
�K�2a����'m\�"2�>Q.O��<Y��[p/ܱc���cqc�bS��R�Z}�ܒ�yr�'���'e��'v�S'�Z`�U�=�f\c�)ǆILm)cJ��Mc��?���?�5Y?u�';2�ɩi,:����=�I� I�wȔL�'�2�'���'9^>����Mk�IR�@B2�V
O&N����E��)J�F�'���'�"�'��	��T��x>7�.}��vE߿l��ܺV��
0���'���'���~�"N���f�'5R���uj��(��3�N��SřKA�7m�O����Ot��?����|���~bo�_�.й&�%E�H+�%X��M����?����?�&�W��V�'���' �dŗ�b�:HZI�g��xQƊB0!�6��O�ʓ�?)SH�|R���4��f됼O,t�vlI�0;z�����M����?�Fm�,~ ���'���' �D�O���S9Z�(��~����ԹQP��?�D���?�����4���O��ǡF3|{��!��S^��شU�谳�i2��'r��O��4�'���'��xW�R\�Y�(ƥSM\lX5*l� �ש�O
���<ͧ��'�?ɇ�E����bB#K���E��l�R*��'M��'2H��%%��O�������F!��3�@��@�P n �A�Hb�.�O����D�Sܟ��I�Tȧ��[�!D��>��<��!��Mk�Bi�`���x��'��|Zc(D(b'ڟ9�dU�S�f�`P�Ob@ꡈ�O&˓�?����?�,OL`aϚtkn]!��3QY�$�%R"!�\�%���	���$���I�|`��!6J�5�֥��.�x�rBA֭�.�IRyB�'���'H�I'Szz}�O������M^H�j �J��I�O��$�O̒O���O��#���Oxl�B�x���������� �@}R�'���'�	�H~F�L|���8� 8��$<{�5Pd'(9��'��'s�'%����'��S���4��?�$�g�Nk��oڟ\��Xy�2o�������ʸ����-0��=�"������@Ks�	ݟ<��*B�X�	|�~�5D �7���qb[�@���ංM˦�'�4��e�gӦ��Ox��O�|�Q�ƴõ��P �R�D�b��Hl�؟\��"J*��?�~� J������( ��GA��&/Z�°i�t�j��b�v���O��d���T$����D�!��3�p5�5���&��q��4oUĭ͓��S�O�R��2�������	���
�c�0DF�7m�O���Ot��u��{쓭?y�'�H���kW�-C��0�)J<wѐ��޴��l��|K����'��'9�̻5Ɵ99b ��l�1��{������[N��&���	ן�'��X7A��H�'PG�"�z%�ҧ����P�ϓ���OF��>�IZ�M�h���BP�zT��'�
T{!�A��?�I>)���?��^#\�止�ႭIڍ��Ǒ��<�����D�O���3�)�3r]�qϧdx�1+�o��0"�;�!֕J:���'V��'��'W��'�Qcp�'����ׇ�]�h��@\GtH�4�>a��?������-8�ą'>�!bk�Ѥ�9ףSdTH�X�B��M�����?��-kZ�2����I$��Y��J�h�� �m �o�L6��O��d�<�pi_���O���O�}�EA
�T�:���*V	$��Q�%#���O���-�*��>��?���M.	��=3AT�
�̽��@lӰ˓`�iPQ�i���?	�'a��I�3�0`cY�5��� )ښk����?�奜�?E�Oo*l�V������`�Z�_�X�1۴4d!����?A���?I���?Q���	�7G2F�J�l�A����7���H&,oZ�,~#<��D�'ox�7��=����k"H)� y�Z�D�O��䍙�<���O �'�?i�'�:���.�̹��˖+���`�}Rʙ՘'J��'kz��Ƀ'] *����A�\��6��Oq)�@�Ԧy��ߟt�I������I=L� �����fN\��4�8f���R���'��'���'B�ӭl�b�Z��D�w\"���#Y�¸	V���M���?����?��Z?��'"l	Th��w+�8�"����_�t�r�p�'��I��t��H���',�$2�@w����$�]y
�!F� �	�mM릝�	���I����	Fy"�'�2l��O��@
ƻa��ek�/��K+H H�Mu�J���O����O���O�H�Aj�T���O^�Hv/�}���S�߶(�����a�I����	~y��'{�s�O���O�[��ɼ	�N4����osS��'5r�'Jq��6M�O��$�Ox�iOJp8��,ƺe�$(�QjZ9cPmZΟ8�'�R����Ԝ|��Mkwo�8d��l�Am#)}�������Iԟ��!CN��Ms��?�������?a�4�.�K��Ϥg�0d��a����?$��/�?y���4�t�Oi���P��7P8�p�Dў+ђ�޴9���a0�i�'2��O����'���'0������t�4�_��pDf&m�ĝ1A�O����<�'�䧯?d�/9�d�2qC��y��(�"�Q�F�'.��'�n�)@OjӪ��O��d�O�������,�ʼ�@�Q�T��7�i�bR�X�*}��'�?Y�����D�T ��J��1HR���M�����M����?a�X?���p�I�6�Xb̮�x��LȰqp� �O>(�C ԙ���ƟX����'1TIrS�!�za�bOLv*�`*�,�0�^OP�d�O��6��"K^�u۬"LD	S-B4���V(,�	ȟ���������4�GM^R�HK� s�(A��UZ"�����Ǧy�Iߟ��I`�	ߟ���,|�@W!n�p�.�+Oy(�$,2,���R�x�	��IWy�	�?Xj��v�#��xk �����6N�8 �c�Ǧ��	@�؟��ɸBNc�����.+�Q�!�X�w������m�:���O&ʓE���)���D�'����D�4E"  Q�h``v��-�^O4���O��#��~��#C�M�����ID�u�P��ZĦa�'f���#�j��E�O]"�O��)��,�.w���j(�[�.�nޟ����S��#<�~!�� &�H�D�*W�T�H�cJɦ�g⃝�M���?����rD�x"�'D�x0�F&Z�����Նu��tLgӖi{7�)§�?Qcܠp�-�!�K0e��S6@�9��'2��'�䡚N'�d�O��$��L`C��M�>,��R[�$K$��>�zb��IΟ �	qZ��xw%�k�1D'�.,��I�ش�?Qr�#F��'?��'�ɧ5VJ����ę�Z�;�8�b�;���@%[�1O<���O���<�F,D9g(��#ȰcC�Ȑ�A�<>,��F�x�'"�|�'��ʘD�����M�6~XjӃ�Tg���y��'-b�'��I�r,N=R�OS�H�$n]�	D���� �,0s�pj�O��$�OD�O���O�*S� �Wi�
4=�l��Ғ{|��:��>����?����$ǩ\&>Y�YX�� �'I���ba��c��7-�O"�O���O���DG�'?J��f�ry��:�慴��'�R^��� ��)��'�?��/?�p:f��o��x���>��]b$�x��'}��$�O�S�^@Z��'ȴ��"�R6!n�6�<a��@=��FD�~���d��8�E�њ}��îYo2Aal�J���ONiP�)��sp�|B5ʂ�_,��al7���z�2Tl������؟@�S8���?�1fY�Eζ���K�8�J����]�0���J��O>��	2g!�1�n�=VV�A���O?l���4�?�/O��A��<�/O �䤟���Ʉ=B�$qp���<�^,���L ��'+���v`3��O����O4�� 䥣rN��S�h�+rh�fARy	òiU2-��y�O�i�OZ��9}�`K]���F^@���ئ����d]1t�1O(��O����OR�$Ǆ/�ZM0�X�Q���]��h��<y���?i�����?a��%��؉�@�(�y�q��)55�mKtb�g�y�'cr�'��'4b��%j��l��L�h1�"b�mT�U��;5Y6m�O@���O֓OB���O&����df�f��9
���4!W�]3x<���Y)����O��D�OH˓z-��
�[?���9
�t��M�3�^�Z5e�S �Qߴ�?i���'�V�k��$��^9����$��`��Л�'���'B'ϒ{3b�'8��'x��ҝC@j��FLH�ȅ��}�lO$���OX�엲n$1O��.wf�8�޶q�qi�l8�T���{�<�zd痹�8%�#@9G8ډ�6-U�]J� m��1.�#բ�0��]�Eٳ?�-8qlQyFȉ9����}�9�qc����QP��U�')�EsE�W,0���UlӎE�0�&B7PK^1Q2b�9V���$��d6��ctf?�h��nքQ6��(�a�cZ��z�c�3(�d"�V�vȚb3M������$(Z`�5n�)o2��ub��4�bc��B�(j�a=QnDy���,�b���xˊ��4�	�*��E�"AR�/M��'iB�'R�i�)�Iޟ�R��� ��d�cG��!��Bv
��@`4 �jj�ȷ�)�p<����Q�
S���aݰ�cT���)wX�vɑ%J�la���vk���'��#<a'KǥG����]�$�~Lj���n?I�P����In�'��29Z��d)R=v ����GFYG�B�I�h� (+U@׸;���07�Ÿ#5ths��4���D�<i���Л&L\�@�~=�e�ބF�h�� ����'W��'���	�O�r3��!ڒN�)��*�`Uz<�Eh3DJ�����p>9��er��e�مa�(!�媒*Q�^��w��<p*|��ğ	N��/x���f�T�*p���aU�5B���ͦ��I`y��'_�O�Sj����&��/R=JAX��5x%bC�ɝU1f-�́)S�10E�fc��	����<Y��R'8����'K�V>��'��C
Ȫ��T�g���CV%���	�����G:���I[�S�D�~ �L	B�:��vD8�(Oj<�Q�ӻNa��I�����〈2o)1X~�<)�����|A����EG\��OR�5W8٫!���F�q���YY@ �pK�{�a|��7�D�rdp���`�LC&���̄7%��dωE0��'p�W>�T����������j4*W8x."�{d�E$@]1�m̮n̚!�$֥t&�`i�$Y��?�O�1��Ɗ)2�����z�̠׎�|�9Q�N�J�FY����N�F���O�Qi5S�<	(,��ʋ6e�L�0��WCp���O��S�SW�I�1��H���.t�� P�NM�pK�C�I3X6�\��c_���u�]�`N#<Q��i>1�	?a��9��Z/ql^$��V��9��ǟ��ԍ�,]rA������Iڟ<�_w[B�'}T���/֊a?�Q�Y�:p`�'����
�I�� ��A�y���dGH5P/���`�]��ɛ;f�j�oھ�J
��J����~����.|O$�JB�ަA����I,X�>��"O"��s��7Xt�]�w�Z#L��06�MP���RU�7��Ϧ!��.�]���Q�#����#R
���p�	џ(�ɘs�j=�I���̧/�t	`�L�I���Ed=���S��ýHa�\q��cd�����'�8�Q�?g�Xx���.g	Z��WF��l���s5i�=��U&;,O6s��'SR��>�� �$��=?�-:4a/�'<b�'�O���Ʃ�3ă�R� �gD��`��C�	�t�9XV�;A������m��I<�Mk����M���n���X�ID���&��A;���2�H��OʹCF��"�'���u"R�T>�Jg��V�fψ$b>!� �,�/�dG��8B��<����,Pߘ��\��(O�%���'
�"}b�K�
yɌ��bĔ�gu�;/�b�<�押W�`YIC��f���JD)�d�ȀJ<AW�բU3�<�R�!����F�]�<���]ٛ��'��[>��ҟh�	⟀�u�Z�i���p�@6i�:m�K�{�r���i�S������j����Am�@� e	��4��c�'*�S��?�����-v�\H�QmQ%�R�y�����jO>E��V���
�⁠V�����)��|��Ʌȓ�Rة�DֳL3��ٴ���|�Ex"�)�S�$���'�Zlyc���;G��+p���^N"�'��Y��)���'���'A��]���]�8.b�9X�h�0�ʹ0�^�Ɂ|Q �z$FG
B��	�"sh����	U�4�O=\=�)b+%����_BhR��?� ��DL�%'���G��}V�h�($��ݥ8�"a+lOV��S
��J��\w͍�F^hH��"O� ����oʆ򱓐��1f>D2��g���$�|���?Q�7M �kѸ|Y����+�)���K�Z�d�OX�D�O��s�O���y>5�� 
;�#��ӶL�������kEB�UL�����D�(vX��D�0$pA������X.>�z����8Ү��C�X�LOJez��0^���� ��5	Vj�O��`�'sh7�.lI6��B�%i �14��.!�#r�Ƙ���҅<���G�1�ax�퉨L�����O? ѾUs���H�牳�M�O>Aҏ2d��f�'��S>5B�k�	H�(�U���\��Z�6᜴�	����ɡC�pUoZ"mZ  '+�<sx)p窿?��!����Z�9}����%�;�xd1lڳ_�܂�̃A�½���+^:Z�	�RPT��u(H�
����׋uvdR�|�g׋�?��yʟ�ɣ�9����2)��"��y��'|��a�.�,�P���"����k �'	Шq�'��QBP�`�`���	��'~�1aG$u����O��'?����?I��"�yu�H�17��)3-J�z���Q�<bGdtY e�D�T>��|�Ʉh�Z	�$B�'e�@{5#_� U�L�4(�LMX���<nX EC��]��?)�oM B:t�-�;:%&��H�r��� ��������-2�������#Ӏ'W�Q��@J�z01$JH��d��H�t!Gx��#��|
��+�4��5	�hHђ����p���?	�M]0�Rٸ���?����?Ⴗ�8�4�
Ѣc�v�H�����rK����O�d�f@r	%,Ozp`Pn��^@�'�Զ��V�O�Y��J$:�0��#8,Ohm2��	��V	�7�aF��P��O�50��'1����Қ��U"����-i�*+9!��Oꅑg�H1R<��)��K��i�B�g���d�|B����7-�rH�uB�-�%-�ȉ
7G�;u`�D�O����OL��5`�O��Dq>�s�A�Ot��S�:T��9����f�N�|B'����C�Y}�t�S�߃W��<���ƕ2��|� ��?9ưi�|`r�D��0��	�
>Ut���'*j�ЀU9$o��b�^�<U�,��'����¨<��� ���9�4�'^�c��@U�	��Mc��?�,�,1��� h0kE挟qT�cCU25|�D�O�DǠZ���1�|��Ȑ g��h�U�^�/��Exd�P�'a�E���	� &�L��r��#V�!t�H )Q��2��O��F�,ђ#��P�����(��S�S��y"(�H햌�#�؃ F�8 tC ��0>�U�x��Хv��<���:�p=�"��y	�3W��6��O0�d�|�����?����?�R�f8a�sh�
���ȭ	=���������	�7/б���3m:L�$.(�2�@�R�������;�X�q�ΌR��aAvk��s�'�1O?����:�Q¦�#M��rǔ7�!�d��M�,��`�m$e������,+���?��q.G;,�F�"�f�i������ɱ=�֠qbD�֟��I�\�	��u��y��|��p(ț�/�t`ci\2�~�`Nr����DD<04��ԄK "DU�Ѕ�u��D�8bȅ�I�Ax�EQ1A[�!��d���O��~�₶�?a��'��I�C�����A,x�
�'�ɩ@�O!D��b�	Î)��5�p�%�S�O�Ƙ*�`jӀ%��,��%Xx:�Ս:1��X�&�OR�$�O~�Dؼ+e��d�O��]L��Q�ԫ�H�脄�t�� �t%�<�d�b��z��P���!��ܪD�آ�E�q�H,�wc��w�Z�a���P���x"a�O��m�&i�~[ e�%�2�EZ>P*�B�I�J��q���g�8����W�R��B䉥Tp�K���@m�Lc�J�{�����'ϢX���~�H�$�Ojʧ,�|���oZ�U��U1"�8S]R})sC��?	��?���، 7	��i`��S��䟙S�������&U�
b��#�(O"�C���C�|��J�'|5f1��#̤>�\� P�ņTjEGyB!V4�?٦��!��Ue_�8�p���@���B�	�g j K�ɟp�zаd#��l��dYZ�Ih?��������N^�q��I�"�xՈܴ�?������A�!AD���O*���1�T;r�Ѓ@*��Uǒo�J�I�7Хy` ̥iU���5�R���t��wu�=�%A�$}-4�Aq�N�2u2�@P��lv���&�7�6�(҃_2�D��;s��X�w-�<9���I�#+F��l3�ώ�?���|���'&�CV���XH�	S���Q,yr�'�T�*$-|UK�+��O2��Y��g���� ` ��LW�j$�T9�����O����}�4Ep���Ot�D�OL����;�Ӽ;�k��).�L�a���C�:�9rJ��t���į,��YB��	��,�g�'4� �ĪQ.	,B� d�@�x��0��%�O�YoH(,�KR�\�*����hO|u(����.����9�P�s��O�lp��'"���$	�*A>��si�'j����B��V!�Y�4�����_mj���͛�'d�Dz���̈́b�mڱ;
�L �E�
�^�օX���	̟t����4A�mA���I�|�$U
d���*��� E�ʜ���"9�H@H3��(�����L���B�NJ�.�c����TY��d!I��Ƣ"w�8!� �,2��ً���!YL��'3P�r5�:cf��0�8T ��k	�'���g	/G�����$S'�pH	�'���3vb�(4��h �ՑXlȝ'��b�XK���M+���?�*���
�^�e��@��S� ?���D�O ��ɲ��+�|2�nP��b���kyv��wkDc�'���)
.�!Ģ�)9h���ӪEUQ��zT��OșE�4ȋ�?qTa�퐭 H�P)B�ė�y��*iܬ��eV�Q@Q��0>�D�x�y(����s�2i§���y��ܱ�"�'-"T>��I����Iğ�PL�8�#���sV��H�^�X �$�,2�011���$�"��O���y�IU0:�x%��Ԯq��hC$B�t�đ���X�P��mb�K�+pGt�D�Y0 Բ�q4k�w���epU �K����c�rz¼��چW.�����qٴ�?����'� �F�N
�pM A慧$Ö�Z�'gB�'\�O��8����Np���FK�,�X��)�����v�V����)�	�U���œ�T�`I��>X�v�'z�����O<��s(Í[�p�d�O����O:\�;�?1�/�Ҥ���	 7R%��f��"̓�-M�h�x�� C�H6\�Bd\`�īʛ-��b�H{�OS0-��b���
3��`e*/@���2�F/���3��e��S�H0��V�F�@� h�� Y| h�+E�R���-�B�'[���|:��L'O>.ԉFL�{�Dc�&A~�<Y$�P�mB7�V���IҖ�:ݑ�,��Oh�#̚H4�i@v��R��8!Hp��no� �C��'J��'��B��Er�'��V�^I�+�����`y����]B��x���2BXm����/Y�=�Ǔ��`Uc)\��x���~J��C);��x%j�/&,`�S"!)O.0�R�'w�"��ba�dCE2E��xB���w��'>����?�O�
e�'M�.8BVՌ\|r�+;D��[ ��}^H+��!R��'y�|��O&�2�j�AT�i���'�哭s��T��EQn�z��Oɮ(�ʊ���I��(�fj�;�f��N>�O���b��)<T61�&0~tЊ�����K�ϩ&���uj�Y��I��O~��C�L�QLRɉ�a�n�����zR�,�';qR� ���/x"*%
�LUf&|��j�Ő2�
Yڑ�W��ji�P���ēW�V��#��v�p��O7:��]�,���p�i�b�'��S�Y���ߟ<�I�u��x  ��j䰙zG`�4!@tc��� >@��E�ѰAa������i0��Oux`A��3�����ʖ�!2��p&�0z�Y��<���1!�^26gQ?�ڣn�ذ��ض\�Z�#�@DS�!����O�i'�"~�ɵx8vOKU�t�{��WT�C��(-�|	�,X�2�D�d	Lld�#<1v�)*uH�*�	ڱE�ɔH�Ѩ��?���y�Ҍ����?y��?���N�O��ɴ?e�8�$�O�n\`r��M_�$	<'���������j]��!�X��0 �O���b�!�Oj��aa�2L���{���`jك�O�q�u�'�r��DU��̙u�8m�4]p�!��!9!��I)E�Ph��-\)V��t�E� i`iEz��).��n�]�B�N�y) �qq�Z	|�|(������؟d�ahFПt�	�|J�AW����@�4b�x=x��@`��d�h�P���I��j�C���1	&��	�h��ЋQ�g�Ba�<�O��
%�'��7��]=�FHڲ��'��K�C�	T$j(����K;V�[s�R>z��B�	�k�Ƞ��䚫z�
��r�|���ɥ��'b^��	y�J���O�ʧ]X����FЦ^��@Z��Ѧ?ײ�9�i֎�?����?y�Ɔq��m�@�3i�V�#�C��ӄy�d�aO�sCNAZ�b��\���<�'�Ɲy{����E&��˕�~d�U�_�Yxh��z
Em�0a@Q�3��O��G����&t�Tٚ3��3B92�+@+�y�^+e��|��Ӱ@j<p�UѦ�0>��x�'���d!@��6y���nR!�y����/<�7�O��d�|�C�?a��?� b�y%J�+�:���e��i1�"�g��4og�S���dL�e��sH����(�j�Ƙr��g�S��?��*�)Dߤ`��hZ B!\ᩕ*���Z���?q��?���'0��oƹ`}$<r2���8�\M��'��'o��D>;��-jbbC�Dx�p��d�p�'U�S4,�hL ѡ��%����q@X6����ϟ��Ǒz[�a�	������Yw�b�'��cQ��+#�]a@ 	6Y*2(�';��h�.�0	�	�5ܸ�d�O�v��\�ng8���|,Ȕ(��
f���bpE���'�Ų��oa{rcڿ:�8�-��\MA2C&�yRɍ:Ψ#�g����4��)j"#=E�@T��6-T41��%�Dƌ��c �N�O>@��O6�$�O�`6c�O��do>����W���Zq#��zf�
�j�t����8.x�X��9Sz@K2��^�'=� ��NDơȵCЕN�Q ᬞ&,�L����E�LHҹ�D��$�6ͳq�	4Q,��dCҦs @�2f��$LP#M}n�E`(D���sG�_E�|Y$f��`S<EԬ$D�,���x�U �	�	y�5�(a�Lz�}��/l�6��O�d�|j�`�>+�|C"#�*�	���½x�~؛��?���W��l�������Χxx�(�D�!q`�H�B��HO|��$�Ӡ#l�8���b�,�1�F"��<i�/�ៈڊ��ѠitYsf͍�~a�HA�#�	s!��I1K�p�b��A�W~ܡa���1]a|1���%&��+2��|9lU����1\�D�30,m����	M��	%�2�'N��-N1��Ö�l���k�'T:��G�,}��J��'���?1Vͅ�����B2C:)�cf�
c��\c�AV7��O?��Z.#�te3`�J0 �&��!n4��:B��Oh�D�O@�D:���@�!~�0B�/�O������(�	fx�<��C�47>(��&,w�zȑ�N0F푞��O��-��)X;Hr;n(��1a6�'�bNK!b30�1�'9��'�rNn�=�	͟�:C�@�fM(�,����խKW󄔧���ɗ2^)azb�^�sh�y
gf�%��i0s�Y�
E:� �"y J�#�-�R�]�O��FxB�ƨ/��hQ�&޻��`H�C(f�.�U�no��ml�?��Z/Ov\��+Z�Wa� ��o�/e��v"O�`#��?_�(4*v锬 ^T���R��A��4��S�dX�L pF��M�	��"_2jĠN0&aɵٖ�?���?i��B(YQ��?ўOw���!��E�j��#g�)u�`�ؑF����Ä�,US�M�*џL���7v��٧�Hr��A!i�@7&�	1K1sld�oW� �f��wA�&� "<	��şT�ڴ.J�a �/�,}p�b���r���76XɪdA��|�z�Jfd؆%B���y*�hh6&�1l�4�A$�cj:����OF���F禡�	|�O/D�q!ǟe@Z���A/}��A�O?��'�b���<t��'��R+�Q��<O�ӟxȼDSO�Vx�L�Ge�r��<�b`E�K�b�R���d
�g�{e�a����ݐ���:��<z7��#T����pm��)�1O�����'�h6M�O.���|z�)C���h�P�լ��P2�M�?�?9���?A���?�'�hOVEY��#Es�8�"i�B�@:!�'l�O|���2(ʽڃ�A�Se�\.4�D�7x#��n��D��I���ωBB�'^B�ѷA���d͓<��ݒ��_����zw�'L1O�3�H�4�A��	�+�>��C`�>@Z��K� 0Dx���'ڎ���IO�O���r�D�,?͜`z�8�2�/���O=�� �6V.�a�@
חwhb�Z�"O�<z1��9)]hѐs�̰:I�]A��	�HO���)Q>m�0a	Q�̐P�kH~|��IџT�ud�w��0�	˟��I���XYw�wF�80��>V)��MB�t��'�(I��o �-{�)��)���	i��-�nn܄��H�2}�R$1���S�C���I� ����j؞,:#-/���a���?G�)�"�*D�P%U�%�Dq�E��,�E�FHhFz���;}A�o�k�`��Ę�@�	P��!������x��ܟ �̟����|�*�J�hE�d�ˡnt,E��+׎>`%p�
t<�{ߓ��G2w�m�g.
I�����m�=%$1���=Iq����I(~�4J^J*�X	 f�T�%���	͟��?�O�����ǜgh��b�V3N�	�	�'�t�`jY�3��u��狞t`楚�'Yh���D@�?��l�����_���,%e�|hGD΃n��8�n�0fs��;��'I��'��J�'h1O�3� �x�b=����!��3�~��E�əea��%U�n�ZČ�y?����
�(O�T1��'�6�A���	s�$���N*8��b�	n+L�`�#������s�P�C t�D�H��Y���0P��?�OT)'�ܣ��ӯ�8��⮀[a�Y��y�b_�P�7�Ol���|zWdT��?���?��)ػslIr��1K4 qm=1�\�������	N�$���GMzeT��!7� ؖɟH�����I�%4�A��.]�B��F0�z8P�'��O?��� �0 ��M���8�``�#!�ܮE�%�C1nj��BOU"��T����?M(�%��:P�e1'�[8&���˟���8(͊M���_��x�����Ʌ�u���y�C=����[I7r�T�F2/W:��f��@�oc�����?�=a`�
��@qp@ܯ��E�S1�J��0k}"m^0J����g�'���C��3!��`൧/_Z���'Ϛ	����?9����'���1�xa�"�#20��	Rn�,8;B�Y7����	Ѡ �f���(��+��j��D�����xyr��Df7�r&��6L@B�.<���;o����O����O�R!��Ox��d>!as��O��$˝L���J&�8q���3��'{ˍvy�a�6F������f��%�#�ۏ�p>��`��(P۴:Ȁt���ȑ/������|ܮ���@!���	�f���u`Rd$q��5_��[w�^gd@�,�m���`�P@�}"�݌]�7��O(�$�|R���9hw��7�@x#�D�7W�����?q� ��HpG�7��V	V?�O���� l�bˋ_e��Ɋ��E�����Ń:$�в��$�՛6tK�i�8TN`8���δ�(O�H[S�'�06-�=�Ia��L�]��T���Qz�e���$�b��s���C �<r�X]{�HǣM�l��&�O��%�� d��H^���� B\���i�|KF��-<C��	�ĔO��}@��'���'mXpZ6ǝ.$d}ȵd�^�X�C��M�_}CC��\*��k�O�SY��t"w��;T"�$��KV(�$q��@P'Sf�m"v�v�dbI���?E���q��x��c��Q�&x����6K�\)�����?���i�X6��O�#~���i%Z� 7Z*�([���͟0��	�V��AC�L��u�.D���:Ր#<���I�?e�ɮS@�<0�l��s�"2�,���� �4��&]۪)�	̟��	����[w���'/����O�2�rS�!	 ^qcD�O�)ôU�ț#������D$	��P4/!{��±%�ݓ@,F�D�J�4�;&:����ߟ��GyB	�`�
�)��V�=��;� ��~"�N��?���'�ڥp�`�L�f�([�p\��t�<��o�cv9�f�^N��P�$��T��"|��hF)���&�0���bD��+j�EQ��Ã3l��'���'��MQs�'�B>�Z�03�'f2C�/p���B�,P(��p>	@�MxyBm	eo���=f세E�Ҹ:��$��ɰI�������B#p5�4���;���H�C(D��'��r�JQ�nŇ~9āS֩%D���Ɨm��x���&6Ȕaɑ�v��"�}"���J6m�O���|"�#]���WlC.Nƾ� ��������?���F��㊛�h�ɧ�IƻWy��	A��Z��A�ת�/Q�����ʻG:&-D��-(���qб'�0�ԥ�(OD�@��']�>Us�⌷J��05ŉ[AD%37�!D� ��Ǎ�<-�AX�A6���C=�O,M&�hi6�����M��N��>�@B��{�\�k]���$�O�ʧk������?��.���r��A���]�7&̧��c����@%Ĕ��o۱J$؋����?��Ot(� �o�uS ��0��1��JGP�ސ����.�xU�`��ʟ"~�ɑr�V�H��Q�?و�ȲEN�H�>Wjȟ���y~J~��M/OF��ӫ�G� �cQ$"y�X��"O �!��J3��qNw������HO���'������&O�>h0Q�\���`0�'�c�	',���'s��'!2�~�q��ߟHs���Rn�!N��%��Qb�B�T
���� O'���j��6\V��}�'�*%b��	)I�Ѐ[$EC&x�^i�CH^"Ly�'� �U=��e�Y�����	~��"����_����G�ܨ�'��Q���?!���'1�>9HM8�EI��b����)�B�I��h�&�G�*�<,� A��tȌH���I}�P�rB���M��.�]��MK��].c"	AoW��?���?a������?q�O!��0s,�Z���K�:6N����߿y� 	g��v����5,Ob�x���̴�� ^��Q��G;�y��� r��YDɵ*i��˓C�}��(�M#�F��?������H�m
��ҵ�Zm����U[��y�!Y<{)ʕ0��Ҹk;��;�yC\/����]k�d��5�]�y��>�,O�@��榁�I�O!���M���h��'^Rx�W
�z�b�' O�M����T�A��0�	��'���*a��$MM�p3���7$�<��Ҝ+�������]���2�%Y�$.́sޭULP\
���b�092��r��]J�"Iy̓s����I;�M�E�i�"U>�3*D�H���/R�#W�Q������M���/��gyBbT##��	 W��U�ր���0>��i)�6��OXSCX�k�~��C�r��,��զiⵏ��M���?i���2&^�?����?�A��K�Tp�r�����!����������<��5���MN8P�X?e�|����j-� � �N$�Q-El1���3K�aalAIR�H9(����5�Ô�h�iۦy\��q�	�v� <�$��)��a���'�6�DyJ~B����䐆"|t#%E1O�6p�%_0A!�d]3ph� 2R��~E�%Q�A]T�tx��Dd}2�� C�$�@��2��'N�1���'�Z1I� �&WxB�'#��'0���ܟ8�I�F�D�w�29>y�afX�K�@�G�Z�m��ba%��?D����?�Fz�(K�?f!z���;Ĥ\��h�]�l[p�Թ!��U�@N�<�$p��Oȑ��)u���uDe��H��Q�$,��+��8�#��O����It&�� ��#`ɔ��nūCifC䉶+Į,�V(���d�+�k¯^1n�@����ʒu�ڴR(�!��kГY���Ҥ�W>ʸ�!���?A��?��  ��?Y����@Z%�?q��P�I��L�%�!b�$7*�vQ��	�`,�&�' f|a ��K�:}�aƝ�i��="1mB-!a��*˓"צ�����1�7 �h:� ��/�*(�*D���m��(��[1.ȡo$���6D���W��)�`�@2�~�Ѫ��g�`�}"�� v Z7�OZ���|U�Ѩ3�%R���U#����bܱO ��b��?Q��Wo����������2i2���L�4�hw�^��Q�(��j6��
Ȧ��Fʙ�T �OƯ{F�Fy�ᄫ�?�V�ӝzJ\Y�Q)J�p��Z�D��z	>C�I�t�l����y��4��ꊊUe>��Da�I%K$�PvÌ�ftZ�m	=1 �ɔ-R�b�4�?1����О' �$�O�����0��H�c&�� �$���͒2D�X�r@사�ik�Oƈ+��T>��|��.^IT����4qh<%��l׍���g�X�
���D`_����)��0`�+"l�e�cJ
6hEj��R�a�I��M�v�i����O��cF�֖4����	�8?��e��<ON��9�O�e�ʻ"���&L� ଙ��I��HO����'���hp�BR�D,<��&��>hb�'�^HL�/vh��''b�'�>��؟����zGm�����đcgی5�0��z)������b�F���9 J��T&A��䐝Q4�}�C'3fq��ˉ 6�[��Z:�~B[��?���'��r�/�>��P��*�4Ud^MY�'��Zv�)_�6��A�*C�6E`�3�S�O`��lӼu�b�P�t�QeER� ��R��OV�d�O��Ś���$�O��e�����O���#B�V=�%p�	C�`	���'c�e�.O0�F�Ās��Q`�ء&Fr�pg�'����E����*�l`�H=>b<�M�y�G�%^c�@�+�cEU�S/E��yb.��ZMa�f�/[��-��!��y�F*��q���ڴ�?�����鍟�d�
�� ���[��d:��ʳ/�O����O�,9e��Opb��'Z�&�3�Ğ�[f���f@�\*9Dy�E���ʅ�ǫN8B�PH��Lݽn��Abs��%4��Dx�O�.y3�Ê�S��|�H�`Cl̐
�'zZ��IDg/����B�Ex�Ȑ�i�'AVHK��֗
G����G� <��#�'���J"�z���$�Oʧ=h}����?	��i���/к0��O[�LzH�+��?��y*���XeA� M��a���7_��\��Vvy��Gx���'�0���>g(+b�L.ly�!��K���2���O�L�m�s̎t�e��6�Ψ �"O�݉�-גf&��^X+�X�O(�Dzʟpar�憰#��	��^#Bm4���O����T$�%�f�Od���O0�$㺃�Ӽ�2a_ A��ꂪf����Ʈ�?�&Wx��a�C8k (U�W���3 �э�~�	���>� ���Ñ�'��誵�\ Y�tbA�O*-٥�'  ��䇏R�t�b4+�v�t�7���j�!��Z2@�!�������I@���Q�P�Dz���R�@��!o� $`h� �O�[������ß������b�
���|b䄛�$�������6����X9-�/#�F����~�剽v6�:��Q1���K��O� ���-uzr�'C��0��S� �u��?e�ԃ�'�"�ض�P�M��pUC��7�����'tR���$m)s�mG��Pp��'@�c�\�t����M{��?!.����HL�FHr���.C�З@�b�<���O��Ă�M{*l ��I�|RS�	n��Yw(ֻ�h� $)�}�'�pj �RR��>�ʆ�(4�����OjNQ�'k>ʓz������M[�i`BP>5+3��!	z����`J:��!�����?E��'Wr��qb�*]v��/�9����V�'ɖ���d͆f��A0#,�6-pƜQ�']��EN~Ӓ�d�O0�'n6��A���?I��^΂��V*Ɖ"�^<�c� �A;�-i�ȕ��?!�y*��0�����q��ýr��y`r"ȑ`���)��x`4/��[}ucٲmW(��i��E��I���S��?��C�<d҄�smQ	4|-*�CL�<Aԭ��[�F�[��E~|
�MG�'��#=�Oe
hI��6!*M��A�H�*����'@rbZ�|$,���'o��'7�aj�M�i�q�v
O�S�(���&��g�v�p&�٣Y�:� T
�{�eHu��P���x�'��L�uO̡2����1%J�FX`���>l���C�N4H���p����T]M�l�q#�Z~2g����(�7=D���*�~�L\�?a6�'0qC�n@��H�
�?0d�$z�'��#��!8��1qaBϛt���Ơ%��|�J>�dBҪzӛ�]�]��5�� ״@��	��A�+�2�'!�'�%Ӣ�'�4��<�%GP)=�E�g��=&��M��K��F&�d{6Ŕ?�~"A1<OD���C�$
岑#V�A%��pd���.����˓"]��[W� <O ����'��7�8e[<$�$�Y1BH��@8?�x�o�F��>�r$��(�,,y�\zBB*"y�B䉟r�ʁ�'��Tx$�� k$��ɇ�MK�����"�2l������q�dJ q�eS�l���Sk̩6��pY��'��'�H ��'{1O��e(�Kȑ�Wap̸vO��cq�<���T�O:X���	%X��=�Mdf�(���b ��)ҧJ&T��ѥ7� 9 tHU0J�Ā��	�� r��#SS�$���/VD ����@άa�A�T6y������D��7D�Xu�i��'��S�y�&���ȟ��ɜ0:��#��>mP�5�c�͑o����%ğ��<��O^غ�!�?[S��`�L(2��*W�E<\u
#<E��3�*q����I��@�%��&>0t3c-��?镟|���'�����ҍ�`��4iûL	��	�'�2�˔⊶_�P\)TM�Hs�Qp���N���i� R��ɰ�Ŵ3rn��Ԙ]$����O�Ձ��A�F�X���O:���Of��;�?�;4�00 �֒:\����J�!�<���y�H�	�KC���a:Y�e1��R�}�/���{^M���H����ɂ�&�Y��\�n��	̟&���	ʟ��'?�%dn�Y�r���ON���
�'��=C#��M@Yg�ʭEx���b!�S��W�������M�B���\\[	�4�ӡ���?����?��"�rm���?��O]���Z
��l�6m���P��0w��(�-�.j�8��'��%	�-]5Y�Μ!�F�	B�V<j�O2eh�X1���1�`�jūB�2���IX#^������r%*��-��Lg�h�	ǂ%D���2��?-�A1'BD8-�>!c��!D�X����(r� ��P!7!{��*�$��L)�Ȍw>����эI�|�ȓz`��� `k����nޅ�&��ȓ΂���$gXΑa��3R�p��l�H�2$-N�vy��L�&� ��ȓu>�%��Bŷ� ��'θj㸱�ȓ/��l%��
H\�q��~��E��}<\A8w)>E�&�X��Z-M�2��ȓ.J���Mp�I���h� �ȓS�V� MV\���	�'g#&���S�? �̂�#J�9�� ap$�2�*�Q�"O�E��4q�M�6DB�$u��k1"O�Lq�
�+ .����L^A��R�"Ox,!��<�����L-�M��"OI�R]>��'@޽K>Af"O�<24IZ,j�f�d�ٰ�5ڡ"O�ș��75S�܊d����1 �"O�-�.[��'��(ߎE�C"O�e�Z�$��D�d*X�qj,�h"O&�+3��:��R+��{��	�P"Oh|�L �8�H���cO�3=fD�A"O��2(�:9���S�ǰgK���"O�`��:psf�c@HĤ~-��"O���Љ�:)�D��b�-�̪"O���%��^)`,:���@񞽡�"O��xg��d( Բ��L�*���S"OP�&e�r|]���ń:�|� "O�Ę�Ș�k�,���Z��Y�"O��2ǃ�Q�ƥ��l�L���Ox+���� ���5���d��b;��	�\L�����7g��^��?����U��M�r��q�ʡl5,O<�ٴ�	��m�Ҙ3���3�tD�#�� ����� �3���I>9]y�3�/�3扽TJ:��$�B� �q���} O�(��/09��Ke�ȟ�P����'S�xv�oRj�S���v��'��	�M���Ɂk��g?91-V�Bc|��Ѩ¸%M���dBڻW��I�1˚E��ɕ���T`��P����$��`��u�'A�{Th�/H3E����r$�s�Z m����I�R���3"(K�1R��j��Ъ�o����s��3�2��F���EA<E��'9�h)a��ծV�x��ܭv�]ᡌ�:;Z���KA��0���F�5�DP��i׼o����'q��E��G�Ӻ��s� �ƪSL4 T�`o^8K$�9q�B;Bܘ)$�xr�S�2�3W@�j���)o��w�.UjC��{y"�a�8y�� w�.T�����	8@nD��4E"|����'M~�g}�#��4]@�Y1��w�NUBT���q�K���UC��sC�D%@}XX��	#Kk�Ra<�e�H��a O8ʛF"��g<� ������	�4�(5���I
oRe��$ګ ,n$�ċS�J&Q���2)%�ɵN#H���L5!�.�9W �"�J��dͻ.�<|�w�P�mĂ���a)K���pɁ�><ʁ� X9h�D&��遘|r���~���H(��E�%�:b��f㉩^�q9Db�Z��'�ԡ���<`=� XCd
�<Pl=3�SnH�CVS�����#�����_Wj�KS�6������A�J:D��i���W(~O>ӂfΘF�\��U�g��A��䲟4x��J�.�<[�#�2o<��mh�U��3%Fx���	S��M��izb�`���8�=!ebE�i�џ��qH��h�09R�+��TR�Q0����u�����r�x�?���O�qO*�jpD��=�!�/�r�R���O�yz��U.SX�d����f�Ńx���Ϙ�3�fA�Df�D�]�f̀�	�H�|�x�y��:[l�z��I�L���XC�R�+H8�VE@��o�X��Ea�$ˀ�	�u�.$�F��#(���y�.T2�*	oi�ĺQN߹oA�\���B'����O�ɻ��å
�V$��%]����9�>���{D��8�C˻}V��D��Z��䏫3���I�oň̘��';��O���h�>���[��Ã_��p�ըu�����Y�Q#(��	�1N7Z���I	���R�	:��`yP�B�zP�0����Zwp�ٱ�@� �'$l|xq��V.P�6%�9��AD��g�'�X�
Dmʴ��q����^E�����O���َt{�iz�n }�������t܂,=
�d���ã��A�j5:!�S6BY "����b�"�s�hƿ�ē}EPD����?�Du�B � ����ձi�!���L�s�z<�T��-%qR�� _6���'�Z� @RD6|��wfC�'* O��'K�=��h�pO��[��bS� 92d��A�6Iw�9�)O�dG0�i��zJ�0G�:�;cI:Q|��Ɖ��s(t,10���wԡ���(8�?ѵlI,<U�Vb���v���H�$���C5/�v����,o���G��8M"�䕺Q&Ez�苐nT�yu@�W�^�i���قoºPC�I�!9�\h�]�]�`�V��u|t[��0y��i 6m���T��EϠ��'Z�i>����	������W
�h##�JR��aT�0�D\�Z$f,�ǠS��H�hJ"-�J~���Ձ(��T �Fիk?�i�*yy҉�� Ѱ)D$2�@�x�mI��کxq�r��Fc�Ε�F���G����hB0$�h�3"�L�+��x0G�ПA��?usq`��%qL
��rN����LI}|,Ւ�ʙyŨ�
��
+G�5�C�C ���S���pџ�@/n���v�@<_�!�q)S]T�P�[�-��A	��"���H/f����A>[���������;)g`�#�UT��X"b�N	�ax��.(z��B�1k�J�X7�4�;#���vI�bkG�Q�bȰCB�w�`H;Db��n>fEYa"��L�$�{���A���� ��5*�*t��w�I�kn
�j&�x��̳|W���D�A=FDP��R��?%?�ɢ`�j>j�H�e�+j�bM#`��h�<�b�G�0І��2'Ǧt����-3�e/}g9hb��P��_�x*�!l�����O����'�`�~� D�C��b���n�V�@�)(�`A��(wH�=��b�* �C���\��0��D�dlPc����x�C4�� 5�ժ^�fJ��E�G3z�Ä@3-�j���h�����U�_�b�J�qMA)^
2Dʦi�:p�`���N�T_��(3��7��!��1k�T1��O.zR���+�H�a��՝.UZ8 /܎VB�?U��0tN�]-��um	�{lh��W�[��O��]
EN�
z�b�C���Y�'d���� V�HE�%q�\�S�O�b�ơٳ0 �C�n�ZL�%�!,��<	W	B f�����,� �'������]�{�ˎ~�#懟�m�@h���0��z�Y������'�f59�� �d�츸�+�(	H>0K��#�
QI�Þ�{9�����$-f4�=ͧR��<�3�D�G�~��fk�>��c�P�8�X�8D�֛l�a}�fU?6�x�a��5.��1��KH�V�a��{��|�F��0��2��#y�A�j��t��IAp��|[�c��0� �ODa�4��QJ�C��^<�ȫ!�ּJ����R�l������^
z����-nM�q�Kw�ȩ%�Ɯ
7���V���M[�oI.Z�f����A�Y~4�#�Q�'Ė�Y����Y�b�z-W�_����'bp)�5O+=q���nQ�_2�����]{�П'��Hu-8h�p(�1G!ғ
�2��`  c&�#uŏ��$����,�V 4n���)X%F��Jz2��Sy��B��D7+��P��0� yrm� B\Uq4*����>i*Rky�P�a�o�^�+��6 "$���/�i>y�s�aYځ�Z�S��H�;Od��b�\���{���x�dk��'��ei�"Qh�>�	 N�"�!��a��
��x242OT��%
 ��p�%G�.�6O�  i��Jo�y00���)���J��EA���'x���C%%ړT����VH�1��c��>|7�Q��.O�q�R؝0MݠT���r�N3����'��-Af��n��s �I[kGq	�T�`����b�ߟ�'��D�*T�q�o����dC2�i>E���>{�=�E��I�6��`�[�w�⬢7��!<�]��O����f��Mתu�B-�|��0���擧2�lM�֭�n)x�Nh��Ƨ�	�d9g�3+40���3�O0���C�!�J4��%J�6@`$h&Ð	k�A�e��jV�"���։�%L��-z�$j"ˀ)+@�U#�Mc��!�6��1�P'th`tb5��b�'Xy�b��l3�:XXL:�'��D���D�n]��Y��{̮�(�O�~QZ��'��q�C��&H�E���4�<�9�����EB��a�X�M�^!���/�-Y�(ĉ_F���0�2O����ЌI���2?�@Jb-�?F;�xP�C�@����/���>��-�� 9*T1uD_ \C���x_"���2�i>%�ѡ��gr�X��d���2`�� 9�았Rq*$)��D�����b�,�b�v-�Q�Ba�-C��8!�k-n��	5n���0�Ɵ3;����6��">A7��.�jA��	�d���5+���p��q? H����,A3��(N�@���H��1#��(�"�/;3m���d��A�k��i� ��7��O�ʓ��i��`�H�!���}��M�%νb-\1[�`�f�$�Ẽ?AJ���u��<b�EҰD<��,ޝ����xx�p�N�}�9
m�&i@�b�D��M l����������t�t+0 �|XBB��s�IKֺd7r tE�S�����Qf0�����5I��,q��h�iA�in� )�JZ�w~j�%*Н6ؖd��¢�����BJ����#&&� ��	&␨�  ��Xw�0��L%@	��-0ـ�=�Zs�	�eJL���U�X�lZ�A>L���A��"�Ks�A4�%��Ӥj�%;'�t���9���q'I�u�JmR��@O�-�g��:��DEC� d��(�EM#�y�H��_�6kƠ?�f J����(ɲ�9⒟��fS�0=i�h�D� g�L xE� ��4@;�@~���D��I�����!#�L���I<�P.��ٖƉ�6�`	 �霬�ZUx7M1,O���������n��z[�9#5jϤ1%T4˲g�)^��Y�.r�vl[�FL�;F�@�M��ELh�OM��O���o� %��ؑ���F\,�W	t�O�Z�lh�}��;{�`�Ր|��i�~e�B�
��YӶY�D�B����G1��H�	��O Y+�M!�I:t�ŸqD�/e��)��蝔��A�(H��$�P������O�n��G��
,0;�!��g)P,&'�8j=������n��OA���	�a{"�
��p�'�d0�i�ڣh����|1� ��G�h��Eڄ�L����c��5�p�A�-�ق2�A� e� �ϖ6�q�B&W4�ay*�[�lm�\�h~�8���W�"�ZE,G�	�Z�ل5\� �x�*��u��F���x�Q��j"�XA$W�?c��� U�xWz��u	�L�v1rc6��(u"�`����Z/13�i>En��S��qSd$6tt���D�	90�;�.W�FAaEK� zzH��dب3]�����e�2�%�&i-��8׭+��0S2&�xyJ?)�m�8)�Ij3`̩N�ȗ�J�H�+���H!��)v����Px�k�1Kjz��R�˸1��%�ݝs���I�J�ƌ�D�Q�n|�YS��W�*F���6�θ8sĂ�R��RTk�J�d�{#�BFY��VLȪ�N�|�>���C�
����&�h�V�x2h
c���tMR�z+2l��k�GC��	�R��X�m?��g}N=DR��� �8�Q9wŋ���|�p	�v�7e�����@ځU���u�4�M� THt��+<k(�AtN�'D�<��A��ʼ���
-$'dyA��#<O�	�	Νʵ��/Z����悈�Q���t�̉+���'[������Mno� Fn�}���5��l O����wB��E!�rzX�eѺAL�{�;O���=�G��>��Ă��l��d�̛�N�Ԏ^1K�Jm�\�aT�X�S�L���<��-�XC������^���)b�P"m
��s`�O�v�@h�O�\X�&@>��k3��nz�Á�@ )���1�g�J#z�q��Y�P��W&czv�'�@� fW�F��CaT�\���[&�6jfՈ\��d.�J�ؖ�ѿvr )ˡ�Ʒd�V��&�D�-Y�i#"|OX�G�;M<��Gd�W<\�y��1����+��:Ħl2E�ԙs��|2Y>��Z��haaZ�RUU0Fk��!�$�h���)�^�����#�
mOp����OO��r�OV8$.����+�*-�`8�5�ֻud�P`qkT�A�1�Tf�Pz����Ɉ6<�a ��!�+��5Jf���CA�V���ȔlO0���I�h	�!ɾ �&��u�\�f�b	�S �I�Fq���� U �F0JĪ��)?�O��b��EG�~1�� ^9x�(�h�*HT1���!��7+7��Fg�v�l�a��:r��}��#,�6�"�Q^�084�:b��!ȃX�K�H����$d!BɣM���M CZ�'VkL՚@��d� �(p���,x@!�$��S��೧��`�xXB�/V5U�Z�z�L<��6�/��Ĩ���0F'(�S��	 ��L
��a�}{ӎ�?_jv-[b�$,O����9?>��X*O�Pks/�zM΀�p�J8L$�@��vw����4P��Y���B�(�]�Q��)�5�I6,��Q����N�$�cE��hW��O%�gM��(׾�?I���˗,�N�i`��";�m����m�n���ԉFv��+6�δ[TjY�V�'�(�Q&jƭ#��!r0:MlM����1v�؅0��r��O_��Ǻ{T���\��H�DكqRh���J�<�r!yrHP��8R�D�G�I!y�9�?�}���
Gb8�`n� f���DTF�<�!��͑�"`Lh�a� RC�ɾ	����@��A��Q��5PbB�Ʌgo�ȳe�{m�x���x�rC�I�5�r�yU��pt��b���z�@C�	�q�h�sG�.m���V�N(tC�(o� W��j!ڱp�ʟ7.�TC�f�h����؁x��	H��p?nC�I5E,�Y��8�>�>��ѡ D��@3��͚�S�\2Ę��>D�A@N�(�~-9��v�-h�
1D�ĸ�C�����j7�O%�7�a�<	dG_=,y8��b�F�}Qf8I�DYB�<�vn�5k�&4>�؈s�@�<�w&�d=�d���y$�U+�C�<����&�&���aS%ߎ��P�}�<���4�dq�V�ND7��bWF�S�<Q��ݑ<kẓU)ј�4`�[�<1���$%�(-*��C���]�1�GU�<y6JS�?>\�z��P1��Ja��I�<Y�/_T�UGHI�3�S6�H�<��`��zk8�a��@3j���0	�@�<A�������B�U	|,P� D����Ǐ.K}�ๅ�R64�H�4D����:^�q�MҵQ� C�o3D���W� )f��Y��N%�X�#1D�P�P�7r\�u��b�)�F�Ѱ�9D��[�A�,�&����=4�"��G�5D������Zo2u��
ͣ��˃�2D�*b��Y��9��Ce�t4���$D�|@ï���ĕ�ů�)-F �a��"D����dףK��E�ňE�n�Ԍ."D��1�䎠c�.���!ǀv�����?D��ĭ����8��@ F�Δ���=D�������Xĺ��a�bТ��<D��A���B$(��E�ni���.D�\(�(G)�(d	@"
l�L��s�"D�X"B&��c!��%@�[{ά�"D��1���(^j [2 ��DP�g!D�� �Y�$�ʴLo�P+�,E�=��"O���ء,ui���	��`"O���bLË��Y�u��)��Cw"Or�s D�7�Pr�AN�i�����"OX�X�=B2�� ���Hm4��0"O*����S��yPmٌTvHyb"O�p�q���ym�Mq��L/Z�$�E"O��E�Me��u���&���y�`��n2�7�M��X9�DL�m�!�Zo�<��  B^x�0,!�Ę��Z|H��X>�x�P����9eD*O��(��D�/�yB��;���ہ���%pv)�R����y���&P�1��Z�M��sbC� �y�+#$L�t�����(h�I�yR�o*��K�9�8�`T��y�k�8Z��A/s��cc�ə�yB!p� ���j_%����7O��y��)��S2G�a<����_��ybI�≠P(�����	XС��y��	/2Q*�3Yp4adJ�=�y�fˣ#��4b���	w��K%_��yR/�`�ؽ����gt�X�rB�	�y��,'p������8R[��ZSϗ��y�n��}��0j�N2Н�� �y�#��dR���e�A�H�X8!�C��yBh��{Wv�K	[��ՙ�F��y�X�J���[$Ȭ���E�y��I�6��bF�_$�H"�����y��1`hx����2I���@�.�y�ٲ]���֯ڝ|D1�m	�y"�,m�<ҴI�|i(���]��y��
t��0��e����wŞ��y"h\�	h��aҋo�f�YwO��y�Q�+Kш�K�b��X$mP1�y�1�����A�Zo�d�3���<I(O^�qM�$2w%��r�#Z���ȓ�����1[!u�2EN�u��IG{��OƵ�e"��C\<��V���'�d��� ��9�Doٹ|����4�hO?7�	D8� ��7/� k�P̠��d1�	~����ơT?U��i`�DD3�pC�7I<m{�b�j%���¨E�#=Y
Ǔ$����f�X7��
%�7xh��>	דi���G'�|v|��IW� 8�ȓZ�n�f�G�R�T�9�I]6�!�ȓ1���a�K_�+V�m�r#J�[����C<��S!�萅��Ol�1��K]tX�D�O\8��Ɨ?Л�Fي6��p���|��IM�x���w�$T��'�H�i������9�ߴj��c�i�9[����M�����ȓ �J�h>]���9�e�X�Q����ϓ�ē9�!�&�9"�a���Җ3?�ȓSf�E�pI*>�� U, t1�'�ў�|� /�MB9:��O~	�M��A�<��	ȶ<�p��e����"0��Nz�Y���$�O�p�ŋG��ˣ�O�(Fa}Ғ>��C�P��0xc/�^���3-M�<�7�Kߤ�P�]=oKd hQF�<����oA�쐇hā8i���ǌ^w�<1�g��d0ES3lJ�cźU)Å�W�'�x҉��)����q��a�P5�yrlP!7�m�p�Y�¼b��P�'q��*W�pA���+XYn�(�P2�y
� �Ĺ�(G�3�z����G
�j�k�'�!𤋳i �%韢���N�<+TaxT�p����V�!�DQ`���@�Se�M�*�!�$�k�j���@=u��x�p��k�!�D�r]tI��1`�QNŴ,!����q���J�� J�o�@�!�.,Ɯ��N�D @!��G�O�!�D'j�F�wƱ2�E��@K�"M�D'�O���gD�B*-�%@�� �P�zd"O���#���2~B�i���1���0��'��I������]�r���衄P-��C�I5ey�����L���2��/W^C䉎hX��`N�!���@�v�C�ɤS
8���L+k��[S�]��B�ɔA��qY3�	�3r��!�W��B䉼'�8y��P{`��(�6-5�B�	�,�~��p�)^��;�M+rtB�	x8�P�
����y��)�kC.O������
;�(�� ~�E�R�!�22��3U��	&R��c�Z. �!��^'*$�ٸ�I�� ����<-�ax�;OPb��h�fǟ0��T+�FѰx7��q�-9��d�����X|V��2��M:"l񁱦<D�D�2͓�u��|�������/;D�D9�.	,����*�$ܐI�u�#D�� լ��ܐ2C~dD<�D�4D����T�bu�i��#7�(b�A3D�0p����g��,�p��$ ���%�1D��B0E��,#�;��,q�1D�L�,o��yK���8vC�91e5D�@��ͺa�����.��.}@�-�iQ?��Cj�2!��-�^�l��h���xt�Iz�'n�D9�i� =w��5aBg^V�
�'m��saW?X��C���ZW�M@
�'��0@%j�S��x�V��V���	�'A�dI1��&x�;�O��O	0J	�'��X	G��#>sL��#�<*5��'6�u`L�b ����AQ4�~b�'�|ȡ	�8r�. ��jӊ(����˓�(O�qˑ�� }A���$� 5�\��"O�87���A�����Y�~'�`"O���4i9�8��-ۏ%ZMx�"OH ��m	�g�	�&"L.Y���"O���$��=�2}JU#� :F��Z�"O����*,�����	�xR����'���+�����/���x5�H���B�	O�J��s$_�?.�l��쉞HvB�ɫuYN��#�"�ZS�a"<�LB�I�3��c@�HV �D��9r�$B�I�Td$m�-�����`���/��C�	}IFY�A�0��d�2��Si�C�	��|$�s���~ �$IE�ts�C�	�Pt\��aH�Z/h|���)y�d�O��$� N
%�s�#�$���!�䌉1fޤ� �,�ft�ìwU!�D����a����Bf8h��ErC2�)�X�X�3��H�xAs!	>^\�5x	�'�X����9pN�="���C�8���'5�x�a��Ds���E
Mlt4�����3]�R��ro[�+V* (�$`VB�I�zR�d��'l(�I�&N	4���*���`��`�Î�Q'Cƣ�Py�ɉ?w����ԈĲvo�����HO���$_�$V������5��P�a
ҷD�!�� H���(G�P�$G!�j�p0"O�AK�5f�nQ��D��H|��"O:E�,�!{6��b��e}z0�s"ONzDҾh2��vjT$`L�""OȬ�NZI�\Q3!�ǿK�PAu"O��â���iܼji�I-J�[���*�S��ԬyL�X:b$>��5hgd@�*d!�d�D�"�� ,Upd4�q��yxC�I*l���ХH�Sx� 3QlCQW�C�I�B�a�a��LlRD�6uZ7�Z���?�
3($��)*^�NY���a����%�i�	�1	>I�U�A0C�����eP9��B�ɛ"���!t-A���UQ�k��D�>��4��)�'a$t��|�t��A���<q����AӢ�4J@H�3o=+�$�Ca�ie1O4���ψO�	�'�"[�n!�����r9�����'1O��JS�"#��9�B֯&�P;Т�4�PxB$��.�>D��D��W�(��/���p=	�A~�8>|��e���p�\�p�ͅ)h�C��"������.Oat�ks`��U�Rb��a�)�	�?HHP�BMO�|:��*R9w#!�D�,ds�,8��Y�o^��2VOJ>�1O���E�ŞvۊuIą	B�.a�&K�ag�Ʉȓi,����)� 9⢂J�$D��>��'�>�ɼM{z��A-¥]�����Њ(�BB�	w� 9�&CT}Ŷ�"F���4� 
#"�1zݨͱQ��t�´pŅ6D��kP(ݢ.��}��՚j����$�2D�qv�@�3Ǵ()�Ն%���k�0D�Xqf�8c7�x
��85��p��#D�BtԈS�^P��%ġEpdM��� D���J] 3fm�ƌ�3 ����?D��C�JR0B^��ې
c��L+)D����d�"$	�E¦d�AX��"D�<����L?5kD$n�����
?D���"��`�b$yӇ��J�>[��2D��
KճU��U�-TAÂ3D��ړcӏ�6Y�B���;@%�0%D��� �A=b?ZA���:wf����!T��`���|�RNܬy$�p"O^eKL�F$0xp��+a7ށۧ*O��ÆќG�Iې,�'h^�	�'�Ҥ���]�X���rp��90���'�F��!��@�x��l�<���
�'���:E@\$3���*w#�0���3	�'���7I�;4NTu��� (.�pJ�'rʙ���ͦž(ۆ.�M�M!�'��m����Qx0)c���*��� �'��P��c\4O�y2�w;0��'�f5���']��!mKg*��
�'򅢦ᕏ�M�@�^uS`z
�'m>{wJ��'�VA+ҟ"�!
�'�R���nU�����P&�Ӏ(��'�^<9��G�j1��[Y*�
�'�LT�B��~�HM��G��P����
�'��Y�b�)%,�q��@=B ��'k�(�C�ݤsJ�X3���+�'p8�pd��U4�Mk'�N>M�nyK
�'�8h�W.K�]��QVꊀH��
�'�B���m 5ج��%��Ev�1
�'=��D5'��d`�J�=l*8�
�'o���A�� 8'^D�$G�==:�
�'����J�����:Q�''�R
�'�tyH���o���a�d�)7�	��� <P�B��J��l���#t4�\��"O0��$K�][dt�G�T��F"O�1�g�%InkʫGha�a"Oxq�W��uҸs׋��
�DPj`"O�M)��T�\4+%j���h�"O^��S�U����)�3��E"OȽ��c/ebV�)th�S�2��"O��[W�+lZE���%��AU"Oօ���78v�he䌍��u"Ou�Ah�a$�@DR�R"����"O�h�'R���X� �L�i�=`3"O� S���}�0Py�HAq��
�"O���cO��(�X �N
[�*�"O�	�cә@����`@V�>�P��g"OX諄F
+\SL,aԅ��$4�3�"O��Ԩۼ *���Ȋf" �F"O�	"��(���#�;3��)B�"O�L�tk��MX0��D�۷}�.�+"O�Crb�? �J��Vc_q�9�s"O���.P��>	�@�K�fg�0@"O.�X�#�*W�q�!NR��"O��RhS�G�P� &�T}"E*�"Ot�Z��8w-`�Rǫ�3ڂ9x!"O�eP�ٻs�B$�7k� -���PV"O�+¥��И�3Q�8(� �"O�����?Z�	4��+~�yQ"O�xp��& �P°�B�+��%�"O��{�� +3�I���� �VmR1"O���Ԁ�"T�l,0�é{!ڐ�@"O�Z�nԑ	�0g�4,p�Ń"O����i�Ld�$D�|m��I�"O��`#A��~��fe�I�f�+""O�Y�L��3�p�q��A��d�"OΰR�B��=�2`�'A̽D��tq&"OV��v�~��0�m�"r�T���"O4�c�f�5EZ�0��ͅ>�f��%"O m�!CH$s2�����ZxD�{�"O���
��he����	�Uc@Ȫg"O��c�h���$��i�)CX��1"O��r��g�pt����0�d�&"O�Ѐ���a���I���E��"Ot����S�!_�$����/g�ԑ%"O0�@P��,"������A��"Ox U���Ciy�Ђ�A��PZ�"Oz x�K��|�@4�3�H���""O$�qB��$>D���v�Ef"��#"O�92�ͅ/�$U�r�_e�X��"Of� ���BBx���ԌL��"O��k�G��D�^����ܰ?δh""O��!aʲMj��r��4S&r���"O@��/��@�`I��cО*��#"O�%�2�ѧ.v�ZQ�W�V��"Of�!��C��� �"D�G�"O�X@EȔ0V���bW(�6Ј�*O4y���>�&�����z*=9�'Φa��)݈7S�AC�"^�4��'���'c�,-tȩ����_�d�
�'4XE��*\�����gR6�Jj
�'kBH�@��`�x4�m�|��p��'��9���1�b��w�J8A/ʝ��'V(�{�N&G ���g��6��p�'�N٣�I��L�J����/<tE+
�'2�1��<V�\��#P�)�	�'kN��CC� b̨H��M$H��H	��� �7� ss,���-7`
9ȶ"O8H�h͒8�N9�U�R�`ef�p"OT�w���Ĺ�aFJf`��g"O���7`Ԣ>D�� �{Nz��"O>ՒN�Au�q�J�?>�(�s�"O^4��gE��dl�j����`1Q"OII��	�εi� 6���Cw"Ord���]N�����H�����"O�HC��οB$bxi�o7	�5Sg"O�P������z�bG�1}�]rr"O^L�@`��W��"&�úN?�<�$"O�y5G���-[䌉{56�2�"OBL)FQ\���.>�Yq"O8��$��r}���L��PL:�v"O�h�,E�?TT�)W,f��t!"O4�YT�F6s�2�S .E��p@�"O!��f�>DE(42S�B�Ř�y�.#^L���GN(hbR��wNU��yR�R�0"��*�̸/������G�yrf	!I�y��H�t�
���
�y��@�(��@Q$�u��ň*��yR�_/|H�HQ�@�(xE�1H׋�y�-��XC�p���6"�$qp &�(�yr��8��1�(��p��Wa]��y��/.�l�ā�H�аRw�*�y"]�D�`���6�b�ѣ��?�y��	�A�����,+I yS���yB���K�$��e�o�"��!�B��yR�-D�X%� �X �)�)ٶ�y	�Z-T���(�'J.�Q�s ��yҁ��W�8����Îp�t�o���y�eE�l������4s����N��yb@J�w��衉��Rx�C�N��yB@۴�����1�K���y��D���q㦓�o��q��ʔ�yRX��UY#C��o/��A�b}C��6Q��U;��;h�������B�	�F� ��aF�ZCz	8�ꃚh�B��!�b��#%�B�T��B0ȮB��<Udx$���	,}�Lyb0c��N�B�	�z�p5Ba�(e�+�#G�L{�C�A��%��ۙlA�+��ǽ[�C�I!,�~�*֓e.��J��;HC�Ɋ�T��F$~�BAY��]�C��31Td0HMN�,pt�����<E�C�	�O�R4�'�#u]D)Kq�=C1�C�I�f%j��'��u��ǯr��C�I7�%X&�e�
%�CEóu<vC�	&R���Ba>gG�X�q��hٜC�	0c��)2������A�e�C�ɟx���RC%Q/t �@S� �3
bC�I�[�"6���[9�\�pH�."*`C��,Q[04��E�`�h���RM�C�	/f���Is͞ 9����� gE�C䉖v-(9�9��Hu���B��B�I����E�G`z�lSR.�+h�B�� /�Lx ������$C�m��C�I�J�<u8��Àon���%r��B�	&h͉��@�@��7�M�<�B䉹x�(ْǩD�Ry��OM�LM�B�98�P�y��-������C�6����'_�UD��
,�C�I�W?�ɚG@�-�!ig��6W�C�	+x��V����D��n�����"O� v��SX,,L&(W�>V�h���"O�p 2��/��\�R��|j���"O^�0"��)aϦ��&��oQ��b "O֔�G$E�� �����
Nhpr�"O,��5�yq�d ��bD����"Oh�+����E,�9��%ˍ>�,=16"OR�`�K�~i,z�=��56"Oڐ3�]uy:��L�|�0'"O<�A��C�S���jv�Q�O��m@�"Ob���^
5���#j $��m)�"O ��F��G���@U
݊S(�(�"O�t��FG�V��(��)�����"O��q�B*h��z��R�B(��"O��A��\!�0�Ղ�5+�zU"�"O��"��$�JXj��<��q�g"O�t`G��Q����p�=4��P!�"O~)"3 Yw�T3.;%�h��"O�BS�8>�@"C�R�Rz&	�G"O@}�RN�.
t��(���E��"O,��b������P(;��$�5"O��c7�Ϻ1������z�T%Ò"O����Q�ƙ(ԧ�15*][b"Oƍpȉ�gǜ�Y�g1���xP"O^�0���!x�	B��&���"O`@
�G��)�6�h�fO�'��<3U"Oh!�P��$qtY�C�6%4킰"OLYXe�f4 3ek.\���"O�Pa��J"xp=4�˃B�hr"Ov���-�I�I-.���"O�ʍ0h��=9u��Td\�b"O�Р��ۉ1\�0Yc:25�t"Ot�bmۊ�2�Xd��,%9f͈c"OF����(LI6<XSI�>aN�Q��"O�c��)���ZB�u\J�"O�d�1	F�j܍��j
�$,�3�"O.-�e��=�D|� �w���q�"O�I�� �jY�����<�,�t"OV�CЭZ�q��� A�b��a"Ox,J�S�b)�X�(x���ɴ"O��SGP �%�4HJ�q�x��"O�h���%(vЄ3��pl�͡a"O�Tî_Fʁ�7�MYN���v"O���@ͽdY�m�
ɕa��x�"Oz��Q�7�.��hV9DHf$1&"OhA#e��-psRp*�N%b349!"O|°E�Gڙ���X&@�ix�"O*�{��?(� �qF4!���P"O�,�m*a��\�.&S����"O�F�\%`��w�B5%�H詡"O��a��
w(�g˭�p�8u"OT���N�9u按e(
1*���Q�"O
�	%&�5I%�!aH�g���"O�m��d	��0��D��("Of@��Z(=ДlDW ��PiP"O��X�*�B%��
]�TfD�AF"O���D�L�=<LSA�5`Kx,P"O4� �"C�vԢ�C_ ?7x��"Oj����'	;�X� "V(b,�8+�"Or��㑮i}�bP��8O���Ȳ"OV��c+F+e.<���&>��
�"O�(�DE%X�`�Y��Y*(���"On,je�J+^��<�b�̗/��d��"O���ޜ-�V����I��@&"O��R���e�X����4�@p"O� .�b�k��g�̽kUE�1Y\]�"O�Ы�F��JE�D[��L�
-���D"OV`�!l�M3ţ	"k��F"OZEJ�k��f��X",^�]J@"OF9&��*U�Yb a�*��*g"O��8�m�r3L����>�.L�T"O�X��f��}�z�+��ے?��5r�"O���!�U��(�	�oʎ��S"O��$
�.���αeL�c�"O��떏F�d�`I��D.1�Z�i�"O�����:k�\H���9 �Y��"OjB�hO�K���IL�.WX	C�"O�(���z~�I�@!Ӿ:ߐ�#"O��'.1��[g�N)1ݔ�*5"OQ�(�O¦��Fa[�����"O�L��+@+4�1�oӗhtx��"O<ܙ!���Ua"���L�Dfڕ�G"O�&���6��vN�|_ ��"O��@á�!I���g�HZb���"O�8����C�0Is�
�#sG��Q"OF�"g�e"�M� h٣4�I� "O�@�5�B��S$f���0`�"O�ݨ��кp�ň�D�R�""O4��V`D)~g�z��ߠb��t��"O��JQ:2���b&P96Q��"OD�[7��#o�F���j�4���"O���C�W���	O)*+�"O��F�Ԯ
b��0-ço"��C�"O�	�� ˶Nx���Mߤ"m�qRR"O
i�3l��UږX���4QL*Q"O��Yg-�!�P�R+B�9��y�v"O��;��RC�N�iG�^ w�`�#�"Op�l��t�,�b���mұ"Od���l]	e�mA���T�01�"O,��Ǉ�-�(X��+��i�"ObK@�h�xB�J����؇"O,��#�#؅RSA�,����"O2��M�c�>�;a-P��@�ه"O@{���T��x�,�7�e(f"O\��#�Ǘl����B	�,�|��"O� �0'ß
�ɘU�1drmi2"OF-P���{��8Ȕj9���"On��q�ӵ�Di�T�˛����"O\=Z4A	����OC7J�����"O:)aeC& ��@2�l�)R���ʂ"O�Y)�g{�Dђe��DVdhá"O�d����5sT0�7+ :Uq��g"O0`BoO9N��I��,d�Zu"O��`��1���G�[D��1"OD���aJE��XF�G�NTn* "O�H��#�I�8e�#/�Z��z2"O�(�3���'�zx�rH�?+5���F"O��*��8Gh�r��)'>b6"O�Q*� ^`8	1jO�G&��Q�"O�<�$�9l>eCV����`c�"O�pӱgG 3��<�RFP-��d"O� ��� ��j��!eS.1.���c"O*��i�
 _���#K�0��c!"O���$]91���C�h�/Ipy�"O �S�ȶ| Ҩ+�gĕjD�R�"ONE�1AN=V�B��Sh�G"O佘 �>�I&�ҨF6�!�"O�r�ѠK8���υ|=b "OP��S�˘+Q��UE�X C"O� � ��1I@��U�]�I�zJ"O�}�O�$�h���Z�w؞) �"O�x�(^���\`f�
(D�*�"O����*��%ʜ1d�h""O�H��ҿ,w��HaF]�<$r���"O�\���C����*_�}�:xYu"O.lӉ�%;s����DǑp��t"O�PѲ�E
n��m�4��:5�6i��"O��8���^&칁"^�&���h�"Od��Gb7�!��/�aP�"O��0���nA{^�� �%�yrOˈ.` �6��o��ӧ�yB��-zX�`�M.\�Ap�Ϊ�ya	
I-r��.��L�vq:��-�yo���'	��C��U���yr�#b���r*l����c(�yB�[nܬ���
tU��#�_3�y�'=DM ]�Ȝ�X��L����yB/�o��f��y
2{�
Y��y���JV�����':����"�y2o�C�آ��ڥB��%!��>�y��P�w'�$� �Q�,��o!�'�Dy�cK�v�td`4�Ӵv&Pe��'MT�s��S��9�c��;�ܱ�
�'Ť����^�O��L�B�9�|���'#
D#@:HM����QC~���'V�j'�͘Mf�u"�Ǫz��`�'��!�M��r�^̉�AA	z����
�'���q��̵k�>��)C�P�'D����j�BDάi��
|	�'�ZQHu͂�>�.� k�	n0,5�	�'�z�PR�Q�.QG���a��e�	�'͖��1�M&W�^��Ƥҩ\,0H�',(����(4�ԁ��aa�4�'p�U"v�K�	p��qd� '`�����'	
Y���"���C���T�*���'���06�n��	J��Z�X�xr�'qډ�5�Y/�ܰ�WM�d��h�'`��"�&��xw�����U��'��x�j�E"�|1V D�vE~���'4,)(�E�T(�0�Ԋ?�d)�'�fR��F�}u�9q�`�2\4m��'ƌxj#a2#�b]�%W��!�'аyu�U<U�5ɵ草$$�R�'�A����&�R�II%N\�L�'��p�aυ>
�5�׬A0H�{�'��!�&_0����,�=�	�'D�+n+�@Xס&�
u��';:e�K{��p#G��=��+�'3��g&P�}e��r�3�T�)	�'>X�Ѷ�M��6���0�ND��'ŘAM�<G!�d(�9
�'���av��4#��;�F0q��|P
�'�Z=鳎�z��0S&�`W�y�	�'����A��{ҡ�Ix�)�	�'e��b�$\s;x��֋M<=3 
�'�BБ�蟨#;���
�&4����'\�I �k�6�tz��� =\pP�'�f4���[;�������>9�'_����Օ+Aҥ���T?�ҵ�	�'�j 6��3|<~D�E�I2�&�Z
�''�œDB�ЁB��/��-3
�'1�L�5�z�]�q#�,���S	�'@�*��ԙ~t�����~ѩ��� �P1K��7n� ��ŘD��[e"O~����]�&�
_�H\���"O��H#)�z��t)a���3[��K�"O�đ�*�&̤,Y���+C�]�"O⍛&,�"����h]b���"O��+C)M#\;�����^�mF��"Op@�W��c�b|r��%'.����"O@8���Άw`�{�M2���F"O���[�R��ر7a�nQ��!w"O�XE�3s�L}�BI!O��`0�"O�͠�Gי��$�gB	�J@�0"O�QuO];��hb�P���"O.q��@ܐmT�� P� ��9a�'�z�Ӧ.�>}>���&��jx��'nH{�p�z�x&g���[�'ApPA����f�6�~��'���9�$3 ,��q�!��< S�'�m� E�<��U�1�@����j�'�b�!E�87\�v����'gfm�_R譣�샲/�����w�<�uş8�h�ת#vꊡ�@u�<��t���z��	`�Dp i�i�<q�'��1�\K�o��A����VRb�<��$>@2Tx8��?}�T��[�<їfĬg����q2��# q�<��\\%�}:cH�'� ��He�<�aN) I�x�Q��"�X�f�a�<ITIڤ3��a2@Y�UcԹ6AHW�<�$�>/^>��p� e��XQs�D}�<�5�¿A5x�K�A��b�Y����P�<�B@_�C<�x�T^������L�<����CK��(]�E[0���`�<A�#�NB,=@�*�8�j��S�E�<nB0E�%�B@C�낣�G�<q%���PU Q��x%���©�L�<�Ŏ�&1�]��-�c}n5K�G�H�<9�Lq�zX[g��T�(g�YG�<i7N���b8�@J� c��Ѭ�A�<iC㋔_��|��X�{�:tb"�e�<�4���W-Z��R�.b��\RZ^�B�=�E��"�f@��e�O!�C�ɒv�R�GR��<�S�(�B�I��������b����H��B�		e�z� R�l� xVAJ�|�TC�>h�%��F��B` 
�<$C�ɾ=֢�	��/n+pE�7�F�$W�B�ɛ\�<S�)x�%8��htC�I
RM^���`W0M������_�>C�5'�ة�� ��m�Z���2k�C䉢�6-��)	��TP��*:8�C�I0[{0%�G�M�?��-Z���W]�C�ɑr����
=~)�EjDcJ7[��C�I!;j�h���ï~�:M��d��?�B�I���$ P��(9�5�΃N@�C�ɾ}䁂#]�	?�J&��68��C�I��$C�HCh���Td��5�!�^�=S����0Abn,#qhT�W=!�Z.iHjei�ӺKg�T�F�A�!�dMc���!Q�gX����$� P�!��G/sD�ʗ�;'9��dř!�$šKD$t��!�?u7иXuS;<!��Џ(vp�ej�� ��!6��7�!����}Y]#o@��檀8�!�䁨?�4�x�ݧQ�Mےj���!�� x,�����L[&��p�|p��"OXԈ�� ���`*;l�C"O P�7��d��B[!�(��"O�|�F�M$�0� �4�����"O�����2�P�+��O��N̳�"O��+ULظ.y�<��.�N-FD�"O^-3'�SԶIk�l�W���'"O\I��|��y��!���b��d"O@��4儆@�j�+����L�b\��"O���S���U/�`g,�6,����C"O���33��<;�a��G�`<��"O��rÌO�EcB�Ҁ+�����r"O����K^�!� �$��B�t��3"OX(;c��@���
+��`�"Oh�@ƕ�!���Ԋ;����"O�Q ���d�\���	� r�n���"O�Qꄌ.TZ�J�ozȤ�"O|��`O�k8�`HUǕ�R�"O��h��m���� ���<��"O"�8�gЪ\�D�qb�84��"O����R/6�6ѳ�d�?��TCD"O�V�`,� `���-�fL�<���@�|��izb�
�h�,}ٗ 	~�<!ӥ��(�%��B��tx��IYx�<q@�GVs�( ����쳇�Oq�<�P˛�B�b�H�*�(شt�W�Ej�<	3�^m����cǋb}&��+Xe�<�F/_G��T S��1��]�<iR��g־�Q �Yp�݁�P�<�Ls��Ż&�O�e�8x�ԫ�C�<�UcL�	ؖ�ؤ�ҟD/��)�V�<!��Ը5�T��B��l���rF(T�<��g_ *�tp쁽8:уfb�t�<��DY�^��a�57re�Gkq�<q���/�p��+ԭE<�)�5�T�<�!���W�r����-u&�; �[�<�'-��̸�P4H�nkb�X�<1�ʫU�&10ф[It�:�&�l�<���P�dXS���7�����'�g�<A��F<g� ���Q�G�p5ƅ`�<���ߐ;�P��7&���
��"�Ld�<A�X�}wth�`P�>��q��h�<iʀ�]�(%EM/aJa{TBc�<����K����KM)thb2*Is�<!��T�p�1�pj,oNy	%F�X�<aQ��g���K���U�F��`�J�<�o�R�����˱y|\i ��GQ�<��ۜ@��]�#�A�y`�E0�O�<�Ƈ��|=��]�J��,xƀ�S�<!�*]5M��A;�.ƄsTH�ҀX�<a�	�4� ���I��Ꜻ���!�$
2W��I�EaD�V�5��+ӥ!c!�	3^��)wԲ#��j�<q!���Y�ԴcgAD�o�D�Z3o�1=j!��ʆ`���6
��oȢ�s�Ӥ-3!���@>�,i@j+}��쀥k���!��� w�����@�9�N��e��l�!�$�.�"0�@�]�S��d�eϺc�!�$O�]B���`�8c�6���$�$D�!�O�'�m�ÍT�G�d8�q�N�
�!��I�4{�F���� �	��<�!�$# ��P�+OUԼ�H�4�!��V�$��1�Œ�y�|���#G�!�ă8#��a��L:]��јt+p!�� $��j�G�N,j��X��=�"O��J�Q#0|�Qm�x�����"O�T$��zL��y�+J��N�#"O&P���Nv�ia")G�x�@�u"OZ`+�o@�$v��'���P9�"OVx�$�A	M|v����K9��|I�"O� n#�}/h��b��!U��0��"O��sv�ƳYiN�XtD
3�^4��"O.0�Ξ�`5��'�'��-�"O�ibpDI�al��ba��U���q"Oda˅�K�0�P��X�4��xC�"O�țCȀ$����3/�$���)�"Oy(����n6�1bCQ�>��F"O&���L*�XSM�~
t���"O��Z2m�:Q�
(U���J��Q�"O�բ�l�inZ��1�M8���"O�q�dϏꨵ˵*S�| �`�"O��z�
@�M��ȧ^ՠ "OMW��, >@rs�<ZP"O(�F�5{*��$�Uq���&"O��S �YdQJ���d�.n�$���"O�ps��MW�Xyd��<�p<��"O!�%�\J��p"��4c'�qE"O*т�I��l��rg� � dT�U"Ox�T ��m%|�����TXl��"Ofm*��Ҳr$F$��TW�F�Z""O�h�5��%IG�h{Ӂ�/@�� "O0��aδL���ؙmZ�8""O�=���H6j����1��z��pg"Otd�		)�%k��$��Pa"O�ph�'�As����̆�` R"OD���%�jπ�Z�e�/=L>Q�B"O�E#v�O-��P�5n�>_��bG"O�|YS�)�J�AL���p$'"OZt ת�D)�p�<6��ud"O���C�� �i#�D�jv^�J�"O�8!0!"F��g�,n@�e"O�s���,Pߜe����*  F��3"O�jWI��P(�@�@�YR��u"Obq
4nS�*-�H*��U,r�aq"O� �p�R&�ڲ��-yF��AbLm�<)�	���[T(V�~r|d8���e�<٠BG=>��ɺB�_�y������[�<�A.��0'| "�G�0�ft)��_Y�<��Í�Eu��a�
8L8i�Cz�<C�˸4�v�1�bP�g��(��L_�<٧$B|���B��D�>)�Do�Y�<9�����.R���w
���T�<A#*gF�LQ�`%%F٨��JM�<���"��%P�E#65h�H�D@�<yV�B�c���R�[*Z����A@�<�$��b��x؂��!]�������<9���;n���遜h�b@�BV}�<��u�d0󮋛F�fIR��|�<���ݬެ�qCbǖ��1�B�z�<9�,T�Y�P�ԭP�y����@Kt�<�2�ב`�
T���+=.�a �[�<���d0��R��Q %�����a�Y�<I��β�8��"��N� �O�<	��+U
��
�J��2d�+��HC�<� ��=x��Ƀ�M�'cH�[ЌFe�<����=��0�o@"�ҹ��"�h�<���	�;7���� >�<SP�g�<��/*!v5s�����+.T�� >ԙ�N��k�za��F�2>�n���"On���Y�U�L�j�K+��cf"Od�9���=��ܹ��Ц.{�P�"O��� cRoU�t��%��PyL�"O�DRtBK�< S�D��O�8S"O�{�KՏR����6��NF�9�"O�U* b	��� ��C���2"O�����H�`BސxT��~�a"O)c�/7���vꆨe�V��"O0�-Mz�K�e\�9EVб��Ŏ�y�i݈hm�͠�V�@>Ha�d�[��y�E޾>�(Թ�KQ4t)ɗ�y��X�R�pXRE�'[�l�#厡�y¦�-r:���r�P���Y��yR�v,�H�/6Or��AD�O�y�+��y"�r�8��� ��!�y2nO�X��h j�$)����+�y��B�M
l�KT(�=xʘ�+��Ƕ�yb�"-#¬��+¹_��DiA-đ�yr)Z�U~��c�ΈX0���G��y�c�n�<Аf��J����ƨ��y�hA�.���ʇ?������y���)�Z��6��e�����yb�R
9����E�,�\Q����yr낰F+�xX���"ݘ#N�y���u��tW�Q� ��l�]��yR$��[���n�)Fb�@�&�6�y2 U<'�����I�Q��5�+�yR�NC��9ElGv�BQ�d�A��y��/|&`��-���lK�P�yB�N@5 	�ce�d�f{.�yr�	+LD "���/Q����$՚�yr �bEH�<O�(�m �yr#�6=��,	�'ԫ9
�ڦ�!�y"�M;o ,�����+�^x�a#��y"(�/@U:W@��0�t�; �L��yb
�L�,Sf�?^6���KC�yb�G� Vr�i�Ve��g���>�O��S�Ά)����"�:Y���b�"Ol(�$�4g��QՄ
�t��)Aq"O,h���/PFȑ�DN$f�h��Q"O�a��4O�"ѤJ_d(��"O�0W�0�,�`1�Yk����"O�uy#�I��|B����b�P@�"Ox��n�L�+�ZV� �Ae�'��')�H�3�h���T`��AA��� u}!�CK��� e�M$~�Ji��®P!�F�@`ZUB��('�ڰ�hB-)�!��3��8�.!T�X�`���X/!��W�^�T�qm�,t��ȊRfۜ!�[x�0���N�P��#%�ٱS{!��X�K��+C��j���D%�#d�7O�X�s�\x�*pI&%��G����"Oz4÷&Лj����cE-���K�"O�5*�j��JW�,q�l�[�"O����a͡%6�� ٹ7#2��"O��!��>�`2�*3��@"Oʉ��Ԯ: 8q oZ�w&mѶ"O�Tƅ��;P�E�Bk�)[(�x`"O� 0�j�b�l�Kk����"Od0�HG�iJL��
��&]�Q�5"O���e'
10��՚��S�[2h�"O+򏉴*3�@��#O:C�Q%"OZ��mE�`#@��q��|��f"O� u��svH��a}��j&"O��kT3����wJ�y8� �"O ,�ŝ�U�,���ʌ�PqJ�f"O�Ec��<f��q`ꇕ?��a�"O�9���լQ��d`c��]��pzf"O�mä��1�P�"ӟD�n���"O2�ٖ�P�O�P�A� H*K� �I"O�p����.�����I��$�r �"O�)�v�]1��tj@g'7�:�� ��S�O1nL0B�]�m��u�U#ɲS�.���'&�Sa݀
�(�#�I9a�"5�'��T!���5Wu^� �c�']�P5s�'�h��!���z���tk^0b�V���'-z���g�A� 8u�M�ctTL��'p={������s�Egr��'�bQ�d�C,+�5�S�ޑ\�<��	�'7���d]%�$�ˀC,�Qh
�'�<,:�ȉ�l=L=�Ӭ�,|�|�'ऑ{el�'vG��R3j^�n���'��h7E�
|k�� c~H=B�',�8	�N��DҬ�{����X��M��'wt!ja��vޝ` ��I3D�)�'��43�Vw�L)�F�!�\�'%D$�7�M=�,�����F�Z�'���!�d���F!/x8��'N���dB¹���c�k�(Zd��')����C�����iB�r\���'"�+���Zތ��!�R�ĩB�'���zvN��5T��e�ӏNw�=:�'���ӆ�3�шt��C�ހ�'��̢�_�TW�Kt(@�>]�ģ
�'mTM���I�G"0��1��'�P#RLw	L܂�g�{���#�'�,kBDׄF��)�BG�%cD�q�	�'�6�����st����q� 3	�'��\�wD�W`��A �Ǆi��	��'#���̃PY�ڢ�(s��HX�'ڦ,�P!+Zi�u�e�Ěe<����'�NE�U��4 M�CD�+^�
D�'��
#@\�v+��p`L\|&Q!�'SPe�J�~�j}�g �l�����'�nm�6��K,����C	4a'p�'�6e�bL�C(@t��g�%J��0�'��p�'�<L@�e���� A*O��=E��bW�Nࡐ& �*`�\e�u�<ٗ�S��<�#��"2�U ���|�<h?=-�lk'f�5�a2&�y�<Q��A�j����W⛑	�X�@Q�^�<I�`9���!�����d����\�<%D>`�ؕ����
o�� �D�V�<�������1Jى8V�hX��ʟ��	e�S�O�$�p �@7;�a��a!!���#2��� AI��0`L����k!򄗐^�``�	6� �ɬP!�D͏.�, `e�=
�L`�*�hT!�dë*�f�����8_^ٸr�ݷnQ!򤊽�z�{�C�/$�@:�h3N!�֟�<��� (�LS�)2�I��<�?E���
=*9B�P��'v����f���!� /1����y�@�S���!���
$Xkd�^O(fm��R�!�D^�M:,�qg��(����qL�S+!��0; ̒智t�x�����=w!�d��!`��ŗb?�����
�!�� �1RuD׻J�(�ȕ��X<��1s�'�󄖮{�dy�2iO
~'!r@HG�b!�Dc-DpR1gׄHlLp0���F�!�$O�hj�iq���(�6mp"A 2.�!�ĕ�Y%�ɹ��6�D	�O^�!�d.l}F�b�f�2�vU���4�!�$�Hf���B�������c��7�!�#]��EV��u�J������6�!��2u$���'oQ9������]8?�!��Z��`���U�M�
��O�!�3d�Z�`^=k��4A���!�DB�~� �p�;-�P�R�,�n!���9j������ >8�r%�����~
!�- )�]�#��^(8|���32�!�$�~��u���o�)��^!����h8��E�G4"5���N�z�!�<L1>|ZS��8���)V
I�i�!��3 �' (p�Ai��]��C�"O�s�I�RJ�#�'P� ��"O ��&LJH|Ȫ�G�Eg0��c"O���φ�h���P���a�s�"O2H�oI�&�XC��c`F0ʷ"OV8��	�9 ,ȐD�: ��,��"Ov]I�C0~���!b-���t"O`��n�0Y/��)��)':.�Q"O��q˰~�@\���[�h�h�r"O�E�
�2����S�9�~�"O�kf�ȋ"4�DjXhmC1�	�!��.$>�!�� �xV`������a�!�d�z��IBq�R�O�8*Ө��!�$�G2�I�o�9@�ر)Q��!�	�x�Z$�&&���'Q$�!�DӖ'΢l��k����9t��(!��Բ �i��ͅ:���`�j�=V !�D:^p��ĝ�V���[`=8E!�ѪS�9�/=��E��ɚX6!�$�+�8���נm�2��1�Ջ3!�$�1])��h�I��nL��H��N�!�ٜy�3ǂ"U�F!�4��W�!�ʌO3ZP��%�[z%�¯ �4�!�DK�J��PmP9
_ޕ��I���!��M��;QJ�TSHD�ȍt�!��أ4�.y�CK���-��ũh+!�D��Y��(�A2�~�i�%ȅh!��1v��D�D���[R��!�di(*�q�ҿq�<����\!��:
u��[ah��K׸x{�^�E�!�	(5��(6��=v������]�!��޻������7�l��F#V�!�?w�$D@!��*��d�r�W"J�!�Y3ju�Mꠢ�/ސ���(�4B�!�G�AV�X�&���b�l���6V�!�d׃$�
�KdFE43��6�ұRz!�F�	�b=9��ũn� G�Q�X!�$�;gю����D�|&�
uĕ�v!�d��@��Dۘ[�$Q	���_!�����Fآ-*�P���:�!�DүHx�z�C�<
�cQ�!�$��0ژ:5)�t�SPc� \�!�$�Yz�Cƃ�C�n�Y�!m�!�dD&fDz�2�˓4o�]ö�G�lD!�HDvnx3��Аt�����Ҹw	!��ߺt �"�u��aB��R!�ą�<�tɐ����.��[!�� ���56ܴ 7�M�
����"O�%���|�앋f��/�)��"O�T��(02���p�J�|��e�r"O�YђD�:_!8y+�n��M�,��"O�*,*�R�h!-D=G�� �"O��V��2�������0v�p"O�Q�L�)8�}Y7a�?hv�p�0"O�Ѹ�D�m ����ɨcȆ	�4"O��8���2 "��'N�ra�e
�"O����C״�A0M͟a��(�c"O 8ČR�����卤�4���*Oh��W�C*y
��Be@��'$v�*Ƈ��bbrC��/](V�3�'q� h��(0����C/İTߪ���'�*��N2
xzF�^�aH�Ѳ�'� I�HO�#$H�!F�5) ^i��'�1�E�>JP�6h��&��Ԓ	�'�����̐�
����)J,M�H:�'W�i_
�ɸ�BFѠ��ug/D�@��MO�/!+�ތ0j9`�D!�y�@�S�D��P�<,ƌ����y"����c����AP�&�yr�P�JEhd�Xu�aҕ�Y
�y��L�}�D��`ߖ����/��yҭJ7:��� W�Ό}.��v�[��y���c�(��@

�d)a1��y"�ĤIx�3����C�o��y��O�'W��*�G��R��L ��=�yh�$��Y�I�<{� �� ���yO�DL�8�+_�u�F���b��y�	"�ޭ�pO�6tζLPǈ�1�yB��	C��T�F�cw���k��y��V.s0��@` ����,�U�� �yB��,���e���$����̾�y��6.V8���ҷ C�A�+�,�yrCz^!KTǣt��Q�̞��yBO���u`p�^7qbl��&��y'��-�
a�s�O�]�6A�vo��y��?Y.A�P�[� v�5�'��y�"	P8H�í�(;�a�$�L��y
�kD�lbQM�� ���������yr��k�
�B�Zd�#�o֧�y�k�4+��0�D� �`�6�1�yR�K�P-�������H�ԧ��yB����Q�#�=���i���yb�D:W�@d�7I8x��L���"�y��<O<��;�i�[�(��E���y򆝰N�b8�`�+J.Hl��R�y�ߊ`� ���	k�4�6�Z�y�ړn���g�a$$��J��yҍ�/I�D#�ǈI��B"�Z�y��
H�4�.�2����##�y2JY�@7.�C��'x���K��y�W&n+NX��*A�k�P[�lں�yr-�*$MhG��k�&�.��y2�A*��@�`i��Y�C Ǎ�y���U��0���Y�a�8�{3k��y�IF����1�(X���n߾�y�ʜ�v?�}���ٸT�"��u��"�yB�WGfܻ�T��a��Б�y�&&zC&��2(�%�[�M���B�s���{iEz�nؼ&�,X��5�"l��;��yq�E<4�9��F]�wd�
�P��.H81��`��S�? �i�M_�7������ܶw��y�`"Odm���7˜�$�@�e��U�0"O��Ӡ��J��1!�)�bT��"OB<�S(+G��4��_�ڐ"O���g��/����Z��I9"O�Lb#��=���Ӆ��-O	�T�0"Ot�{��,9��Ї��U�š�"OءVn�9���ও�Gf9i�"O����7](\bc�
�/p j�"O��j`F��e�U��$�2�N�9�"O���я%`�����W�L��A�E"O����� �G)J��f��.G�"غC"O,t˂�J�7��r��1ڌ���"O(��VHP�{��@@YQ�x�b�"O�X8qCۙ!��;�ɘ�N����"O`Q�#jܚu�}zP�р{S`���"O�h1R�@"fT5�u��
/ȹ��"OZ��W䆳Mdh�f�1��	�"OR��6oؚv`� �']�G�n(�"O~
�邌`(v%ǜ{�6���"O���	�,��܈pJ�0�ґ@ "O:}HҦKo8�T�3K��Q r"O<ݣB��DB0|r	ܚ^x�`"O���+<rnV4�pG\9@���v"O4 q���%0m�K�͗K\��a�"O\�3�U�N���h�tC8hyQ"O���S��6n��a�5�b�"OZu�&�F�i+��W"3y��D"O�Y���:Mm�SB/k�`�:�"O�cE�EG��Q���_�D�3"O(Љw��6^A`0�7B�6���"O��)�'@3Cj�t�EcG�9��\��"O4)H��9P��Y���=����"O��j�+����v��
�*8��"O��a���*	���CA8� :�"O���ţ��e�&ݚ��=/ڢ���"O  �fƏ�f�8�����%+�"O��Q��'W�n�����#I���Q�"O�
�L��ZE��`U�'����W"O��̋��j��Tk{ޑҶ"O�5�3Q�^�d@�AD�wf�y�a"O�LBEi@�U���Ec�sQh	�"O�؉�F��d��
�,�1�%"O�Hg
;i���Pb�P1gt�A�D"O��5��Qm@@�A@�=�ҁ��"O��5-*9�$�s�hg�:%��"OH�@��d\��H兓=m�^�q"Ox\B3Ć�(v�X��#ǯ'8��k"ORe9�J�63hA{��^[,����	MX��P@ �6^j����@�1�8�:b�;D��\6�Tb0lY3�ҩ�0�� |!�$�/� 0�@\(��-("���co!��͑U�r���^6<3�_>v̺
��Q���D�2p > 2@��=[�M2J%D�����\5Vg~�{Ѫ˯Bҝ`�ˤ>�4�O�>��F��o�&�h���'p�튖�Cg�����DG�F��P���׬t̒Xa0f7\��\�Hb�'�֬`� M&e���eʢ(�0ez��:�S��i$J�<x�h��U��ٙF)���y+Ե+g��y�ʓJYF���J���O\�	`��u�aʙN��m�&o\֑i�CV�y2E�K' �&�%[<�b��_-�Ie��(�z�*4nI�B I)���c9�����'"��l�=�!u���� ï��C�)� * {���c�&�j`��?J�'��q����K(j�X	�K�;Q&q*�'�!�Qkz�1 UU'J�h˥ҹ%h��u��H��`D��
�Ą��?d�C4"O��h1/�5)@�P�2[M��Å"O�aG��讔0B#乚�"O��0����L<֤�l�"lJ�+�T���IO $bċ-Ts`h��=�6C�I�,m��
Ԩ�i@"� ���6R�B��pg�y�c��
m�բ�N�2\�O֓O*�~�) B�{WoUIU�]RF`�{�<�QϚ�C��)��kUa���s�<!5a� Q��[�労h_N�	ƌXr�<aƦ�2"���F'ip�*�U�<�ףK�!���5�΂~�89�[�'NQ���O�D�{��H0KA^qr��:*oD�9
�'j6aHD�	#iJ^)"'"��x1���DG8��9V�T,J���^Y�Q�3j?D��s�A�&��C���u�&D�>&���'��_�>7MŌ�h�$iH?{��BB����a{�,��G����68u�Cf)�(�挓��?��iv��|
��\=ZhJm0�8���D-/�\�"�OO��TL��X9D9��9Xr}��'��9�f�F�3�|��3�<��(O�6�5P`c��|"@���3�6eC®Y/@�rœa�m�<)%F2hpbus��P!8��	��_Jb�!��s����gܓ0<Dȑ�Qu��j� ���a��v��p ��־Q�r���o�	86Ņ�wn6 �שB:
њ����i�8{�'S�ѻ�mS/"��ZW%�.zxdq���'��)F@Y_]��r�鏳��"�'��i˖�+kհ�w��q�I��'��pIOΌY'��U(J��f�+	�'g�(���\%��(T�
Y�P�	�'�B��o؅���Z��˂)_Lńȓ3u�c@�^<,�)�����|m���ݟP����B�� ���S�k%O��@��k�ah<1r��{���h#F#�FL��
�O�It���Oͨ��wCL�g���{4A�+hY��'"�t��+,���_& ��0i�OZ�I1/�ɧ������<�^�"b傜(�!2�D�{ء���`�-i��)~d�d�H���6�<}��'�=�$͞$$�z�1�m��hH����'��0I�#%:5��W'x�6t�	�'�
�C�K�xv��Ш^ c�\!�'ۂ%°ɟ%K��Ф�\~����'�d����.
޸4�PLM\�0��*O�����9{��,��&G�Z"�/��!�DO!�(8�h�)		
 (� ��!�$�dA�DG˒K	@m/��E!�'Eў�>�s�Q�Y��J���)fQ�$�!D���Pl��l6<�ҫ��4x�9I�3D�D ��V�jDk�Ê�4�&��� =D�貖��K,�(0��G�	Ldԉ��:D�����!PE��ڀ�/t!rd8D�HX����J��;�`О(���P 4D�@q��Ur��i@��̠-S�K�1D����n]�	�Cg��PS�㥪0D�h���J/Y�a��$D,L�h!D���Nʫ;����mZ_j����A D�p�"��/�N�7(��1c�咑�1D�d�M  �Zxb�V�(����E.D��2g�"_Rx��O�"g1�E视�<1�'�a{�G�6֠M#�C�#NF�)EA��O��=�π ��
)7{�	�Ș�D5��"OBK�kݑ�v���62j�s�O(�=E�oɇ8l�\9�b$��\�k���hO"<�/���X�Ȫ
T�j��1&�$��>�����;���i�J��bL�a$�`pay��	�}b��Ă�z��˃[g�B�	&s*Ep6�G�
=��T�:۸O��=�~�%���t�h�b�r4*��QÌy�<�CG\8��Ę2�`ۜ���)T�L��Kȕy��a�"Do�cs�1D�01�e�\"(yeo(x!0X��.p�̅�ɺ	i:�A�	J
*�L�! �f�����9U�'���a��K-�l�¦
r��:
�'�`X&�S�#S5�n[q����4ȸ'���s�Z�9�B�:"����@O�#����a"O�=zU�K1b9,@����
�9#�X����ɧ}�$�#�FB�$�~Dѡ��7gU"�<��T>}"��
�?@�1-P!.����-D� cG�T,�6m�5=D���-D�X��g�	2���ЌN�~?�M��,��'�O89 R A��l�ʧ��%VO��K&"O���v(:���K@C@�AY��"O��������T�%4aY$1F�O̢=E�o�&m���.Z�x������y�&���"vG�'$=��q��yE�]��m��$B�XE���yr��i�uY͊@%r `���yR��6���h&�ɔ;6�y`h�����<i�u��� �-��s'��i
�	a��I�G( ���45>Ͱ���%�ȓ9�DPp�:=�@4��f��52Մ��?�OI!�<�R��.�F���SE�<�ԃI8�А1#�Z�m�H�X楄A�<�c!+��R"��{6 ��|�<�F%��$�2�2�և6�l�r��v�<Q1鄌;3f]�t@�+ݴ,�R�o�<�jB3��Mp���b��5�ŦT�� ��)��eE+26{�భ�2�,Qae2�hO��7���UiͿ6^�!Run��cFC�ɪ �*��ߠ#6!���_"_[�G~���) a=�!�F�h%K��͒�C�Ƀ$\ѐw.ؑz���a���C�I�:3�e �E�+.U�uru�̛[l�Ɠ/���
�g�?;"$Y�OܔJV�ډ��?-�?q"NǱ[����.a�*e[Wkf�<D�/�"-�d�X�L��)�`F_�<1f��zh�	���w�|���
�B�<'O &s�űA��Z�F|"��YW�<v�M<0>�2��̈;�j�k+z�<)�GƪٛҢ
tT�h����`�<)��rI�.�� ��S��]��vD�EIV"j�:�[�A�w���ȓ<�HQH��]{�#��bP��� ���Qр3������҆3`����$E~y�@b҄X��)�t*׻m�$h�ȓs�.�B��H�Ӻ��$�Վ2���ȓV|<q$)J,G=���ԍi	j=�ȓ�������3:W�pWBE�Jن�b*܅J�o�J��|(Vρ�+�I�ȓ>�tQ�b�> =j���.khؐ��3������ .7�c��V�	�^���©��#[#5VJI��S�H� %��*ZX	��f+J�Lm��/�q��ȓ=�n�YRlӟ"���8�'�1R���S�? ��i"���%1�J t�B���"O�����j9�\x��Xc��5�b"O�Y"��Fn@�B�����"OH��B�K|D�QV/L"P�+c"OU(V�	$i(@�̓WLe�7"O<���R4'60k��Ѻl�伓�"Oj��c��i.0[s懯C8�Պ�"Oz�2����bǚi���\�h�<sS"OX͙�FA'Sa�U��g�%:0C"O��X/�N�֘�6�(B$S�"O
%����0�2 ҕ�����D).D��e�)-}z�3�	��h�L��*D�,�f�Po�y��N)q<  �'D��T��u'|D瀠#i8b�F$D��R�ɗ5��qm�@?[gd�8�� D��)0���_:.�+F�Y�|���H��?D��C'��+�RE�D�˲G�E�ce!D�s��(ej>Dsě��H=��`>D�Dq�H��� $-�~$X��:�/a`)��!d��T%Dllϓg8L�
�MلmR��jq!ԣU�̱�ȓ\�.��s��3��T�Ƌ�{�2e������/X�P��!��#���чȓk<8����7���y��K�h�}�ȓx���`t�Y�Z�4So�/����v���K�G�X�,}be�f$"���R�" �C�B���Q�D�%I�T����x�hJ� �����a�$L��Tʣ��c$}Y�O�霕��2�4R�)���E��� �(݆ȓm��	�gք*%.ٙJ�t��І�=�5 5�@�K�x����>a�y�ȓOX�Y%a�4_ � ����5i�6���>,\I����	�d�ɬF��؄���p�B��<EpT�r���S���+6L| 'I=X+@��©��o����R�qB/E=1~yx���?n0e��\�̬�b��N����6+��ȓp�
�CO�8*���T1G����ȓ ��R�-L�+^�|��n�.۾х�:N��J7�Ө*�>�a��l�荅�h��� �)o9�"�K��ل�C��`!Ƨ�]�rb�� �ȓF#TQ	�Cá��Ųt,��tr���1��5�#�0v��܊�aЊ_���ȓ^"@���R�rLh	�.؋#	V��ȓ���#w��S�6!�!�݁.���ȓGi�4��� "I�c� �~�bфȓ7:rx��$YD�裏��6""L�ȓ!,h��4u�1���Z(;Nx�I#"ORӍ�b�ҁ0fI�b��|x1"O�9#	����c��5e����`"O�U��G����!��$he"O���tȚ)����0�	39e-(3�'�����Ć=$�tU�� �6~&�P��f֔|!��	>l<Y)�#��8����ě�wV�'sjYq��	w�S�Q`8%�b)Øǌ�Aa�O	6�D̄ȓ$,=���m-�	Q��V�1 F8R�{b�Q�)c?O���a�C-02��BǴSya��O~�P����4��i�a5
��M� �.�k���������HY!Ui��E��	�/)��r�|�+3�~u���;%]�,;��;�y2�ǅ_[�-�Щ�7����'*���j��4�)��%6\�!�M�/Y%��i�hN&H��B�ɭF��8�snW�1���c�&�⟨ᡯDU�� ���ٓY�8�'E�
m ��"O:a��M
3�=��.���h��"O��Bd�,v�R#��0��"O�{A���c�L�X5× |q� ��"O([�mǸ-�8�Z��A:`ت�"Oh�3��M�;�"m���'V�$|c�"OJ���īXîp�G'��s�r�+""O���hý-1l�)V&O�c�b}Q!"O ���ȅ	X,�x�����Aa.9#"O�j%��;�u�T��T��e"O,=!�'F�[��H%� U�� ��"O��#4�Ƅ@TI����.��+�"O�T�qm���x4���D��˥"O�<{�� !�T'mJ����I"O&p�FK�8�0A
>��sD"O��#c�+��<`��� l��5��`�I�n����|��x�i�L�ܡ�w*�7�0?15��}m��c�¸��{�,�#+�t��i���*���,�O��Y����WH��k��i�	��Ik���s"Փg��%�-�z����u\�SH?N�~�R�Β9�y2��jYȣ�M8b����(߯�M�Ӏ¬~��i��Z� ��5�s�f��f��:D\N�΁�a"O2E¶BJ�V��Y�d�޹<��5�$a��n)��
X=���{7Ӱ@�<�g�'��<�<N��m�D�ղ;n���dr�XQoқb6����`��KV�z6�n��pv�9{�D���'��8q��S*l�<U#�ĕi	�<����5dw���vi5T���sBJt�t
��)j�X)��n��U���B䉪YŒ��b ��<���+�({n7��~�B<��c�ZxdXoCm��M��F���1���Fھ�su�C�<�sbʻU�u��T��H�r<>"��o6L^*�ҴA��JY༸�����;CG�_o�a���0uL�㧄3�O��g�$v�n��5M>��Qʠ�+)��5����5\�~������
��R�ړ+KXY�ተ��r��Մ.��dp%��*ʚ#=A��؍B�H�*QK8�2��gȎ�X$�+N;Fǅ9z�;u��=_�đ�$�O�U�����9l�P����I�ֱi`�Dg��6��U��*�4���ၶHu���?�@��5�F��L��('ԾyҠ�	�y@���F������"����qP4��m�dm�hX( ߆`h�Z?A3�k��A�R�f��ü3�A�1�fIʦ�Y����S�
Uu���X����t	ܧd`����n��$@�?A��E�����m�A��F��+ԉݤ�HO�uz���#Y�4�c��*������'[�(��M�/����7�]�b��[q���U1 �+4"�^5Z�[�}�u��xX���0(�.?b�1e�*��ə��:�$��)����h���J!�R�WUZ����ܝ����3h���0�J�< ��Bۚ-�!�dJ�H�6Y�fj�4�qeᏤ����*'K`�y��R�`
q��m�'
{(���wHec�˓h��ݡ��'I{E{�'c8CHӲ ��U�c(k��{(��5�09;+�$?�<��V���r�3�s�'�=aA#J*��F�E+x��ӓK�\���Ȕ>ۂxǈ�H�Z�&�^C�;̆(�M�T��#Ubb���'�]0�jM�dȢ�����E�P��{b�[�#W�h`0��Tl~f�Mp��8BU?��F���\��u�v%�=!:�(��,D���v�3m�䁡�jZ�_e�b�.?�5W��<ȕ�����z�nޢ&ϐ�:���	n�}`�"OR)9��D�Bi�� �;JF� �`�r��v���)!*!�3�� z4(�π�knPm1�#ʣk�!�DW[��3��50W�Y�W���!�D�0MK)�����U�yH��	7�!�E�R��0�T-,�X���-�!�d�1Z��D�@�D6p@�e�b�!�Y�&������J�����.�:|h!�A�Y�n����	���)TmЯ[!���;b(iQ-I�g��EB�[�PA����0�>q���b9ft"��) ����C)D���d�r�\��`Ќi�@7�ա:M�m2�@O�{�S��y�T(h �!H�0=y�AS"��y
� v�k!LČ;R�J3�7"�i,���AgC+^m����dx� �o��m@<�`�'suԩ��+5\O~$ �I�w��bU$�>hHF-AuJ��2Sc(+R=+ �G+%�!�I��4��� .-�Na0$
(�qO22E���HO̙h`	�6rc?]�%��_%��C��Q�g��x��7D���Ш�6|���@�Q�����2���o6Z����Z�Z�"|�'o�A`���9n��M�b(�3
����'����,;�B� 򥟿M�5�7hN�-����jU�&W�����C8���s �5�Z�87�"?s&eӥ#=<OX� g+�#;z2I�c\:9 ��XgaB�jA���K:O{l��F�t$B��">�:��@��B���z�&���O��ZW&��"����˒�(�ď;�Ө���FJ̯9�Τ������tC�Ieu� y7�س!	��A� ��8��5 �'J�p��K@J&b��H8�L~2�_�5l�q�>��-(P�W��x�!^^&J�
�j�"pʀ��J�
��e���-5�*�Z�Ǎ*eܦ����'۔T��EO�!2vHAo�DTHϓL�5
��i�X`(H7z��d+F�J��AA�ǭ,K������x����z1�$Ud
zt
'��<��d	r`:������'@�MgXIH���G�	7-P�rJ�!,svm�.�y�&Y	;�<$@J=)��+s�K�o����	1E�ȣ��ϰ2�Pɏ�D��Tc�وi�`�d�G���G<D��(G��J�0��6	�=���]s����,�:d��H+��ےx��x"lZ�cd4Y��6�f!x��N1�0=I�n�q��񧙰b�h�;4<T��.L�s�*� ���'��\Z��\$n�2P�mJ�Nm���D��Li�Y�e��6o�U�&3��
r'��	e뙐/s�	`Q��37(C�	T�H$a'�6_��I�E��
-`�*�dtyӅ+4�?� 1�gy�&����H�rNQ;rB��!�
K=�yB��}V�7�ӽ%jt�3�^��M���
�`��$MvD��$�
O�r�
7
]'o��p�4���!a|�C%x� y0.�'J	��#��A�/Xt��ƣ�9x�P
�'��ܑ��Mp��%)���n������mU2T���3%7ڧ-;�ѐ�)	�#���� U�*IP�ȓ	��)t��I�$�2��43��8�`�@°ؑL����Y�P�p�W�J���CRh �����"D�(�wF�=Z����l��u�ތTF�"e.ě���	�L�P�h�m�4'�f�Yh��h���Iw����G$^��Ql�>]��Z6�в!�|���Ͻ��B�I"O��(��\L��i
��@�uʂ�H��9cM� )2��q�O@��P+J��5����qT��'i��귫Jd�B}@���r�JB5��x���y�o�<9a�5�gy�)\+F��Ͳ�	�=h�.��v�
�yrK�)Ar1R�U�_�ꕋ%��G���*t��%�@]���>lOVP��U�tj�!pu�IW��rR�'
T�92��'G��{a�i�	�T��,>c�]ZZ(��Ȃ�y�,^K���(��T�n�4�p/��׸'�`�g�*d�vL���S�I����W�ٓlz�}�r�Ó6PC��3��Ph�o7!��ex�m��ME&,#�MD��u�O�DD��O|�c�c��tK����m��/�>\�Q"OHTk��̈c �k�Σl��Ѳ!�'}Ȅ(&"@��a|��>��y`Ʌ^�@]B4`C��y� M�e���,�L&ba;�$ٚ�y��
6_ϖ��!�J� ��У���yb��4�,!��һ��Ex"c��y�$�"(�Qd��h�8��5�y�lA�B9H���wd�/�y�� 
����x�n�a�m��yr�F�j�� H�Es�t�S��$1��gSv�Z �H���@�<�T��ȓN
nѠ���	+�`�=s8��ȓ	e��&��?��@�fA�4"�z@�ȓGfu�@�8N�RV+J.�Fp�ȓ%25���$�2B�� ��ȓ 8��'�)���R%�Y�GT%��S�? �](�F�*���4���c*��"O�h��`��N�Ȇ>[Z� jR"O��{6��-�`-���o��*�"O����(�E(�iP(lVRH�"O�Y�mJ�m�䍡���Q�l�I"O�MZ`��mG����J%Z�V�`"O| S�A
RE[V雐 ����"O(���K�C疵���ڢ7h,���"O�$�!�O*:@��1��>m�=��"OD���J1DT��	x�
��g"O!�QM�4��̠�Ń�B�p�"O (3��M-56���Mˍ�F�C�"O�u�#�\�R�P�@1���}����"O:Yav�ߘzXv͑�fӗj���9�"O�]Ia�%~����O\�5Ǿ��\�<��Hws�`H�E�07h�
�_]�<IR,�6w~V|�����N�&�3H�W�<�	�
b��4��l_�ԡ
�R�<I�mսg,�|��j8�`bA'�S�<�ר�(6���������e�UH�<�7K@
��D@�=+_���i]B�<9"Ԩ{|�8�;.�ި��Ly�<�'jm��-h�d�5'�����
{�<!�+��|+3A�e��kt��s�<�!hJ:]��"�-~�#Ko�<wbK�Q`~��ņU�<�z�
���k�<a0��R�AZ2mJ��țy�<��$�(V�X8�m��l3Ўu�<��eηBD�x;�K&*��a��SX�<I� к@�NDȲ����Ba�W�<q7`�?>��E���6��i��X�<�c	H�1�j(�V�y�čz���yB%���)A) ����7e���y"e9_�p�2�	
�LYSWi�<�y�b�F7l�b��V�Z��퓩�y��:'��Y�E�Wfެ!6���y(C嘽��M	�[�l�kV��	�y"� �vy�P;�@B/<PYf�G�y�φ2���`�u	�xJh��yg@�`*	0��ل2�P������y#��G�y�g �E�Fqb@J��y�9QYdI���������y�j�J�|K/F�}�4�C�_��y�+�Za�C��tx��!2�¢�y�A�  �t���`ͼEh���D�_��y"��]r@}���܉/J�У넊�yR(��i�4���+�I��+
�y��[ٞl:�KK��	#�J�y�@�\n"�1�:j��hୌ��yr#�"c ��ф۹�d)q@$P��y�n���&X"���� ��w���y2�^�D�c���B�*O���'�޴�qģ�n�Ag�'P[h�I�'B��P`�"��B�P6*!z�'%�����O����Tb���'��K����0 �!�a��!*}c�'xv�S�/�77d � �~���'� 	��+ ��퉂�O!xL
�'_	r���<dw��#�%ܝ3�@� 
�'��p*B&G#o�~�ё�հ �.D�'j�1��V�k&`���J�p�l��'��ԩ���9dH��� ]�Ld:�'K&1��m��)]�.���q�',�e���������x��� \��$����b�!ܐbx���"O
D��[;,�k���]F��"O|�뇥�=WF��PN�%MXpr�"O��%L�]P���Ā|5hi0"O��.�`	:��p	^�~'4�8"O��h�J�(�ahR(R�+����"O�ԙ o	��Ҥx2H!9G���"O��)�.ƥ|��-��\��c��U2!��!��z�e@�z�]���4$�!�Dҳ%z�uZB��>��Ko�R�!��5s*�Q����8���ad/��s!򄏵R0���S�b�͎�!!򤅒g�>M�1������"#m�:J�!�D���1�$�JYQ�木�!�@>��+��H����AC�,nq!��rL�벦�>t�B���C��i!�D-S����$M�eh�Z���Z!�^�Z�D�_"��Pn�'�!��+X���4��P��4)�l�'�!�>xxA1a�S8@;�-Z�B�&p�'�(J#�'rq��'Zr�{���ø�P��4��[�Bs�����:X˺X�s�Ղh��i�f�"�T��ˤ9�^��$��E�%�`d�Zx�M�v2ў����rL4!�f���u�O�vqy�a���*V��L�J0"
�'�r���m���ڐ�_Dhxz�4������P�WF��!��MM�?7�]���҇ B�@g�D�2� �!�d�'o�L���'L��B�C��m~�a���i���5#֪zB�p�qM�~Fz�C�M��+���;H��Y�d�I��>��)��8�HX���.R���Z�
�thb�����Z᥏�C�a~b%�8t'�(��j��(��s�Ǘ�HO���2�ݹq �u	׎G����O��@�%�D�uyƅ�a���6U���'̭B�Վ	 �`� �$�&��޴4G���ѣ��d�8�3DW5ԑ?7��?f�h}Kv%�3M����#�%�!��3#}v�1���\��qi��ۜ>��$#·i0�HA�8+�<a��g�~Fzb�
f"���! V4	�cM��>�'01Ҕ�{��s�����N�3:t|sR#F.$������)�G7&7f�R��'�ԁ�B�5V����`2H�!��$�k�T�P��Λ)�ѩ!	�!����T	�rdsB��X��9`瘺T9����Ƕ��?�e�H>)r0�V&ә\҈���Φ�w�΀��p*��r{��!+�U�l��ObvA3"^?ט#a���^z�L�cc�	)P�B�I�qr%k��� )T��!jF�O;�|K�aְ#�(�G�Ĺ�n@�t�u�T �>/�� �Z�^���.�c�]"n �+C	�	9a~�����p)�H�L�(i@� �M��y#�G���t�d-���8Ċ�1�`�A+ȦJ�0#=Ab��zTh鴌205PW�_x�`����5$(���#J~q��˒b��8ã�2�㲊�|�8ap�K	2>xa}�{d�Ğ �\��d��Xi@N>�4c@A �'N�GZT�i�LD�J:p ����~�EP4^����ѣpC�`�f�<�jO�0,���e�3�6 2 �$5��Yc��TTV�i#-҃%	�x*��i �q2�ڀu:��dH��ʵ����B�I�?J�x��P�d�~Q��I:|�ԙ��!�V>�sf.ה}������>F�@��ɧ&~���h��o?�Y*4w� ��dW��!ţں}4q�CDP�!pp�	*Fv���Ï�1N�A�.� a�����I����#܃&�4�7�I�������\T
�@��&�� �@�:I�9�O!fP��+�EJ��CFa��$8�'���ȳF�0A���yRN�2-�^A��yB��/�TQ�c�6 xmiG�L%<�
��ǂ��1��B�I�|����RCZf"y���ׯފ�٧�9�	nGQ>˓pH��Y6옛����$
��M����ySLy�&��0~��)��I��ȓ=��A��2,��u��$�ܹ��V�r��fܞl�t� p)�d�>���.\�u�V�F�H�P3�eNp|���;�aɥ�̖u{�����>z��ȓTK�x�J�5t�2m0�iվN8d���S�? ��[�LعJ�J�I%ϓ!U�4A"Ox�.�d+ /�&2���"O�0�C�@�n�N�aS]&�ڀ�'"O��`*_�V²�r�#�3Hwz��"O�����}����-��QӇ"O�l��,M0|`�R�&�w��D"O<�"��N�B:9b�%[�)��M��"O1��WJC���xtr�"O�1�w�]�=VĈ���MO���1"O����HW�C��:n�%?2X�T"OҸ��� 85�,l۳S�Z�X"OZlxf�Z$hf4��b
�ik��@�"O��ѵ
�-U��K4 _rr�9Q�"OB!p6��0s!��X�!Y��[�"O %��i]�7���2&ZE���"O\3v*�� ���EI "6ik2"Ol�P�4l=�+�evDI�"OT91�C1���u��&	kh���"O<�C0��VN��!!���oT���"Od���O
���zA�H20�}�3"OҠP鎟a��e�d���b� �"O��Z`ɑ$`�<!�TDط��@h"O@̀W��=P��)�c��(&����P"OH�(T��T����a^�(�"O�@	H�hvh�P��F{��Sv"Ot��A(�P��U��Y=h*���"O"��gŇ=Qj<ۢ���f���0"O�i^^in��$Zm��@��"O��3��E�,\HR�?��#�"O(�r�
$�Fۡ'��Ż�"O\)bQJ(R0�}b��J�&���JQ"O�I8�^ �p�� S/.n�x�f"O�)�W�/,��R`.�bZ��1S"O�j�B��щ�-^Z��Z�"OV옠��8xTˁ
��CU"O�u��L��>���6@E4�j��t�$ԍ�*��`�9�'�xp{���,,m��C��ܫ����ȓmL���&Џ��p��$#bXh����A�_j
��H��`��Y��Q6�ټ`��e/ÏlP^5Чb4D�h���j�p9C�\O9&��%�6>��8�V��0rĽ�ۓh�W���wCh@�1@�%��t��I�z$��I�::�ql����%��>L��q2`�N2�@C�	�v�)�V�Xճ5NO=yp��2�矿4 �����Q�Ot��N	7Hp��8�P�0
�'l�-R�HM*m��<����?�ҵ�a�P2�̨n��ʓuhp�|�'J�x���Kb!���c�<)��i	�'y��j���v���P�A��:NP���G�-%u���ތV����?o{��àdV�j���P��yo�z2+��t8����G_�u����+/�	����'�	�S�3�y�'	�N��I��������'q`����A�<Nh`R�,�NH��후*�j��e�#��C�ɒiz4��eM��1/U7��=����H\r��O��G��O�tr ���\���KV�J���3�"Oz�H�$�&I��8�d���lP0A��'M�`�tl�N�a|2f̛c�Ɂ4� �>����K	�yKY�z��Ԩ
�: 
�K7���yBő(J�%b��o��\p�h^��y�#^�l%|����ҔXv ��A��yZؼ���.y���B��K6&����'�L�a��YM�D ��O�$I�)�	�'�ְ要M�W��p��O�&F�~���'�@�w��3u���:�EI7CHX�'Y4�sd\�xq�ǈЃV�ިb�'�p��*���� ɽK��,���� h��J EL% ��'B���"OB�	���|� ���l�c@��"OF�;��W�Kۀ��+G�9:��ٕ"O�q��λg��ȰUʢM��u�"O~
e,V�匠�e��kC�8(�"O���6"Jsc�!��mAA�pɔ"Oh��E�p�`��,Y�oy�y�"Ol�P,.k:x��$eS�l��"O+C���E��xF���� c�<%ĎfF�EJ Ǜp�t�c�d_�<Y�M� Y[H��NAx+,ј��n�<��(�:X��ձ%�E��^M(��j�<��1�t� �(�+���s�n�<9��\;((8 KU��"P�["�C]�<�*�!Y�1��j8؁�iC��y����3��@s"\=�A9�)��y2�^=�\Y�� �'�Z��
1�y�쑸�r`[�ڢ_�Ys��+�y2��~*��#�F �K�Ơ���X(�y���1Č�0�X�Mr*٪�@��yr��bfl�;�n׻�	����yR��>"R�� ��M2+<�"ǭ�y�)YsR&�+V�5rg��ٶAK$�yҨ�:XY�dBl,����y���3*���c��ܽ�5�S��y�� m(���2'˒81ڼ��ˬ�y�^%a�PT�@9ؔA��@8��O ���LV��!X���5�()x�/������$D�'��4L����r����MK�>A0����y���){�d�ґ���Q�B0� ��"��'�|�h�'E�#}�'sB}���&8`p<�@ɝ���'�2�	��)�'�н��ę�7b.) _�8H	�Lt�ҹ���OO�?�A ]�P�`�e�<k�h���#���O|������/[�Y�#��ottb���q�;�S�:p�Ͳ�+I�T��m���8�dO���2�	T�q�R$Q����*lQ��O̵R4�'������F�S�?i�j��=��WEg�h}�P�ԗ�����������0|Z֫���]TB6�^��u@�K�<���N�2
T�y�,<��A��.Q<���N�&������v�
��ַ�
�Gx��a����Ơ��Q{�J�:� b��R;1O�	
�5����B�F6М���O0}��u�ȓZmtT*�,�
i0�m8$#Z!�V��^ZIY��с"a��IЯ�8�P��I�����J��� /B�$��  m�#��U��'� � �>��ӊ|� ����u����d:S���$	K?r�Y/ON�"��{�OD���L�g���u��_($<��`
M�&�|���$:���{�I�9�|���[7i�� ;���xyf�oܦ}b��k>�Ǝ��SbA$c�Z@���1ȱ���+��*�
�O?����*]`�D�B 0�]Y5�^�l<��%
A�, ����~��O;ʑ���A�t���RG�ls�xa@H�R_�<���Q^?!Ƿi��)��O�ݎj
���e[��t	��}�逰� _���I>�g�Ӻ�Z0aņ�y�E[�ǒ([e �ȓF�.(�b	��^��!l�%��хȓb�(�T��>#��"H�@��ȓ7*�Sb�[�B���í��>�<�ȓt�Hy�c@��5���v�P�%3`ą�4������=`�b��&�i�ȓj�Dp�S�B=m��#g��:M:�|��A�Ly�mIms��y�&}�ȓ,�zPA�eL1#v�C�Wt0��'�d�	#ʿ]Uԙ�I�Y�(��=�|�#��x�xzC(�g�>��ȓ:�\s�aG�&�N�Q�!��s�d��0������\h�L�2Qg�7�d��S�? Z�@��	�vQ����i��2"O�H�CdP6L�@k ��nd�,K�"O�0#C P9yvf�hF�J*��q��"O"�1��Y
*u\�a��"AT��v"O�T������v|�b^�X�u�3"OL�P�/{B�M���8(Ȫaq&"O�=Ѵn�	:�� շ.��H��"O��"'�|�� �Kr��{�"O")���Ҥ6��9���d���"O ��B$_�ሓ�M�r�"O��81�ŦEDJJ�h��:pp|:�"O��*D�.Sц�:d�d�$"O��K@HU.��u�&FDK�"O`T��B
6��S��6�N�h�"ON�����<�j�� �-4}�c"O�(�r��;$�e�dÑ�m�,a�"O������.�Jh�6��6-�	��"O|�C��`0���),(���"O�l+�N*j�~�5�R%>&���"O�����R�Y7�|j^E$䑣"Ox��!�U�J���)q� h��"O�����$M6apDȣ'�jP:�"O����&��G��`�e�2l�` ��"O��!FC��`�X�x���qL���"O���)K+=	��XÜb��G"O�@���+���NKMxj�Ju"O�y�E@��s�Y$f��_.�"Ol�2O�9^qD�i��F3V�.��"OBT�%g�&)]���*p0t�@"O꥙��J6,�8�T)Ѐ6mDm	"O��V�G"Jᄤ�e5F�IZ�"O=fo �ɷn>3?XX"�F[!��@�;_���$+�B4��s夁�:b!�d��x��-�C�ѫH�8XwŅ/	:!���6F}����5
`D���2\9!��I�n��SƇ�g�� Dˌ)!�$��8Fn�T�޾Zx��ѵ#�5+!�d5o>,u�0p� P��d!�dU<p�,=)��АP
܁�Y8u!�?K��p� i@�h��4h��۱"�!�D�hj�a �_?D�	c�A_��!�܅i� 
DD')��|���6I�!�\"-s,�P�ǈ(�
�p���b�!�dæo��	Qd�;9Kf��T��hD!��Q�r�Z�,Ć^b���#��P8!�J8
Jt���E%JF^��ň|�!��s�RѳbǢ=�q�1昳�!���;@��H�gB�t��@gN��\�!�G����H�)B#��ⳬT \�!�Dۜ&�h̰�z� �C�k׆!!�d�1Jѐ ���ٳY�"�8q�E�1�!�$��h��(:Dʞ� t�̻�!�䘺t��0�E�<�M`�%̦]�!�$_#��T�$bį'�2����`�!�d��6�(��H˱P���ٳ�͏w�!�	�o;��y��D�!e,�_6�	�
�'��hPaO��6X䪃�B�^�>pP
�'��$p�L8o���K"��3*�ʔ��'���#T�H�C?��!�UfJ���'E`��&�@�X�
r�WD|p��'Ph�*`A�$Z�ځ�ЗS�^��'��YCI@�f<ZT���O�apl1h�'�X�+���_ ����π�Z���	�'�TP:A Y�j�|,2��Ġ ��y*��� "�)q���+�+�i���͊"O�-��H3ܶ���� �Pq!"OZ�����,*5���H�l%��"Oޕ �@y�
���<�`"O�1�� ��(v�+`�^xv���"O�`3��$�X[V��:2J�ip"O�5K�g�F��!"дr0��3F"O�1��$Iu�iB��%y-^�W"OR ��C:Fɪ(@`��*�U�6"O��(5�
V�^�tNŗ1�����"O�A�B䑝C��a	�m�/ɤPJ�"O���I�Z��9k0��+�^!	1"O�L۳HL�6'���ϕ5�:ɑ�"O2�zU�B�CĦ5j6aw�Α�E"O�Ի� �V@�����*iqԭ�d"O�-��c��9߮cu�;��S�"O� �&�Z�������<4�6"O`��n\�*!��	��ѻ�j�I�<���Z2g�.E*5�Q�K��Eڒ��E�<��g��s�1�a�R N���Gl�<1�!ē}Fj��pe� yV��H�k�<y�)@�N�dԳFe_(k�\�hC�Xh�<Q�o��a����]�r<�`�e{�<y�N�5�����	R:�S%�t�<с�զG���:U*�-O�"u�Ir�<I� ��1oʔ� n�)z�D1k&'�p�<q�c�U�ms2����0��^l�<Y����lȊD�I�(��.�]�<1��J{������E�Y(�t���^�<��	ǌt����fF�`�a�U�<A7@ 8T%��jE�Ċ~kt���	T�<qUɋ*0R���VbA7����m@w�<��ʍ��D��r�Q�7�F]��CVH�<��f�Z_Z������P��M�I�<����
��@U��@@4$�@e]z�<��(����4�сX�
D���N�<Q6�Ms� ��HԹQ}�У��P�<�SoO7��)3�ġP���P�QS�<���Y��n�:�&�f�6RsO�<�C�>�hE�F�-0��t٣,�p�<񑫋?5�h�z��*��P���W�<a�&A�X��VL�*@�e�R�<yv!!7�`i��bM q@�СY�<a7,�'6|!CO'R8z��)�T�<1d��63�5�-${JHY�GFQ�<Q���r�H�R�J�f����l�G�<	q�H
Y^(�àC�4@Hq@��h�<���� 7���m��tM����̚h�<�dF�-76�8@AhF��I��c�<�&c��F<8rF����UI&����ps�
 mj:��j'�汇ȓoE��`�R9>�@{V!���ȓ7Y ���o  r�r���H�A�ȓ�l�Z.�R��=��Éyr�|��r�H'dX �<ؓvK�VL�t�ȓ^MPa��)M�F<�I�ֈ\�H�:A�ȓX�(9u�1�~���	\U���P�y�3��>64~!�6�ݘ/]�݄�`<)�6kڋc/v!�b�=��h��Z�̘qCɉc�*��rČQ�2���O��,@P�ґFU��ՌL�b�D<�ȓbc���Fa�, fj8��=�j$�ȓm�����LWt�؂�D�":�d��{�̐3��^�7� bT��*����S�? 6̣��B""���(�G?FcƑ�"O�%ـ
�B6>��`�٭@*�|c"O�x`p�ԣV���E�Q�N	y�"O�-)��ˮI+(�r�d�O��Y�#"O�u���.F	ٴ�Ϻg�<
�"O�0���]p���۵7����#"O��x4h��Pm�!���H2k�@�""OX����`�5���Ń0����"O�ݪ����4� 2G��<\�9P"OR%8���9��@"I�JDYrw"Oj=�	(W�pŨ$ᗮL� W"O�ؑ�	UJܱ������<5�"O�%�%-F�V]�`�@�U�v���"O�X�V�R/n|5:��G b��T�"O��jg��p�6�"�.��:�*	��"O(DuĒ�pgn�+�M$l��@�b"OB$����"{�E�h���SC"O�5�WS�
̈́(0�g˹} �2V"Ov���@Q�L��i� ,S�)@T"Od��7#��~�f�*vo�.k0�x&"O�����A7|��"�@2�b"O�Y��lƒ���P�`
�ͼtBV"O.���)l<H1*T#Il�8�&"O⠁E��l@`y����KgT	�@"O�d�$������c)X�`R�R "Ō��i�> �f����˸EpQ��"O����֘>͚|��%�-`�X�Ӧ"OH�{PΑ�(�v�z�
�y���"O�lb��.�VM8$�E��� �"O.}P��܌���z�2q�|a�t"O�9��DԥG�,i!�f(�k "O�̀rꋍWh	 W �='���T"O�`���q˚E�N��4q"(��"O�����J9'� �WCV���"O8$�V��vP�d�DQ2�La�"Ot@h�ꃪ^��\�N.&TA"O05H2錢3/�Lېƀ�U,�H��"O���Y�� 0bƄڶn(<u"O!���˖%eA2�~�f�$"O���S��v�m`D.�쬹C"O&AP7�0|��$bc���V5��"O�@%Ǜ�Tͱ!݁EYq�f"O���$�o��E��d��Tԭ�"O��'�'x�	���C�i�"Oz%k��5���V)ȵ�D�A6"O�H&J��N���1	�r8ݩg"O�UhɊ[����AD�L��c"Oj��f�"���K"&Ӑ*Q&!!�"O���e��C�L�s��1U7h��"O°aGKQ47LX��B#w78�z�"O�$��+��.�9"G�P�>�ȭ��"O�H�Pm�P�g�5Q��u"O 軅̃�5�4�yC�G5f9by0�"O*�@lE;FX�(���v7��s"O����ݲO��Т GX�sFFY �"O�5jpgV�0�D��a)+l���y2��#^ P  ��     �  3  �  !,  f6  WA  �K   V  �^  �j  }r  �x  n  ͅ  �  Q�  ��  מ  �  ^�  ��  ߷  !�  c�  ��  ��  ,�  ��  5�  ��  l�  � � � 7 & Q, �2 c8  Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�� |d��"O
`�(�;���8���-0��1%"Oj4��ND^[��"3/9�0|H�"OB���H��*�ʞRy=a"O�味V�!X��!&F�:J�$���"O,��a
���C�Ą�M�"O,$3%o�-���p���+Ն�:1"O��ݢ1����`���y14]2��i�<�6��{_���c�H�`�fX�$Kn�<��A̼VI�xR[�)�Ć�pඤ�ȓA5��('nߡ4�� �)˩%� ���,��r�؊b#`T�eT09���ȓ!�b��g��}�8�F��-? �ȓ
K|m�ș�VṔ���2�%�ȓ"R�X�j�4JN�1�˘X�i����̹	_�jZ��1!g��zܶ��ȓgil,*�J�
j�Ne��i�J%b���f	�(U��:���G��$Y^م�~r�� S�%T"���k\�jx�ȓ|4�1�îJb��@ӵ�ݩn�V��/[`�"�v4�R�!ʎ<��M�ȓ`:��z�ؚh�J�Z��$HY:	��H��p�m�C1��!��B:��0��EnjZA V;9����J[
2���	��4'J�EA�IVW&��~�(aZ��ӹ�>� o�Y�|�ȓ�f�A�
Ο7�H��M�$�����mޠP����/���ANXo*�ȓTv�����{ ��-7�*h��I��sB�8�8���3����ȓNe*M�悡;������X�o��!�ȓ'lj�#F�m�+R&;�|��2)n�C��0S4���T:
b���:�0!��e֊��)��ͷV��,�ȓ0�&�8#���� ع�L�����;�P�AFd���,w�6d��r�EQ�( �gVlɦ�M,H��,DP���|�I	$G#\���ȓ"�)���E�B	yt&B�^�LɅ�4�� ��eëF�ڙ��n��R�p�ȓp`@}bŇ�=�$�AUN��P����L��p���_�a�)�Y�!��-��u�5���o}�`iF�@A�p ��F�\�0��[���IF/5���k>bTؖ�;K'DT`�^��@��fnV���Y�b�lI��	����ȓ,nٛ��Ć3���kC��8�m�ȓ'� I ���x<=���޳{��	���`�'$$t��l��-�U!3eL�X���/D�"�ʼL9�ɻ2O�/C�����,��~��$j;��H��GS��DC���2 h�B�	 

��VD�-"(���"��I���OR�=�}"�E�0$\��2�#���89VoWuX���O�IA@�Рg6�5#3�V;	�Fx2"OBj��ÒO"$�;�ɄS��h���I^�����5�82���jW.ဢjX.+!�d�!$bx��iS0:���w	;.
!��N�b�1X �05�J9SF(�?+a~�T�p�2�W�1=���/�>���f�2D���'�K7i3ּ砀< ��� ��,�����O���Ȃ�Y0j��禃T�����)��<�s�Y;=$橛� X=V�|D�ŋ��<�۴�O?� �]a���tu&|a�܊�8G"O�вR�Ͻ$E��↖tc��������	&g�dС��7�����H�7���$�<	��@�ȥ�7G�P�Ҁ�w�IR�<yOD�K�K,�(�vd�.^�C�	���r�U�y�P�s���L�bC�ɀ�b��'��		���%
���c�"O�EJ�)˸R�\��B�Cl$xɇ"O�8	���yO捚��ߡ|L�i"Of�bIǷ0�pY�$"��u3&���"O(����P.PfM����x�8�Ҳ"O�E0@Eдp�A!3�v�"Or]����*{��T�` �<[H���S������$�U%��/��񃶂�J!6�8s��b>���#�L��06�mZ��|���<�7䜟b�ޙ�w���T���$Z��P!J ��!J%
L�8ž����	$x���7�����L)=�)���*�y�Ӹo{�Ѥ�V�]O�%������O��D�$�߱&�Dp��X�#n�10�����HO���
4"(����A�M=��Ȇb��o��I*�HOQ>Ŋ�Ą.92|�*��R�˦)Y,)L�C��<g?N��%E�8����lj���p���>��K��<��� �ۖ��f�(<�شX���D���@ڀm�Ìj�t%�?r�)��Eͨ��Ġ����FX�"`ۧ�yB��!Q��&�#^n}���y�e�U�e8&Ŕ<Uf�u��hH��IQ~��x����iT���ժL�$.���E)ϼS�nTbD%=$������8@b�$�A��0F���,+<O&#<�S,
+�����hB�+ j�_I�<�2��)sa���El�"@�1�]���(O�<��4K *5��j@��{��E� "O��(r#�����J6��Ph� O�<iW����(ZfkE|�2��&�H����K>�dl��	w�੒��P�JhC�A�	z���r�R2K�h���?T�tu�=��W���S�-U��Gֆ\B�a�;��C䉅	F���K�M���A ^��B�I*\��!�R�|�F��p��0	�nB�I��l-�7!�@�yp"�
����~�b#<�����v2Hԙń�#.��A�%6!��"�Ҭ�@�6�ѐ����]���D;LOV�C�� "��<c�(Ԑ �Z1[�"O v�\�]��`ͲGŬ��V"O��ra�٧@��1�b�gYPa��"On��"���|��u�L�W�8�"O���p��"�)�u(E_
��"O�CGK˹w�v,*�G�0wQp)��'o�O~8B�G2��1�fa�d�"O��[@ŽA�t4˵�CQ�\0�!"Oh$�竈�H���*���QW %���bH<���%j�����N�o3rI�ə_�'X��G�D�ɳ9������ .�&�� �
�y2�� ��7�Y�,;ll�g����$��(O>��DLX�Ic�I3J�nȒI�.,4�� �*RuX��O6l>:L�Q+�V�'�ay��!h���F+YY����́��'�a|��W� �8�#��px�"���!���3c���a4͈�RA��Z3��#+:!�D˹>���i��S.�	���h�!�dL 8ʈ㚙5#pb��҇M�!�DI�wA2��"�ô-�*�R ��a{��d�/9���≪q���H$ �rT!�� <�[E��r��Ȕ��l��%P3"OZM��h'�PUc��ϴ+Ѧ��a"O���p�P;
����fk��֨��"O�dׯQ�^~����?a�m��"O�Ta��N9^��"�
�@c�A�r"Oڠ���S=������LO��'"OHp+�鄋Q�Y�Va:+L�S�"OE���M|�YԥJ�u1�p�"O���a-N� N ��E�;j��S"O����k�=����o��؇���G{��i�8/�j��сNÎ�x�jԫP�!��OJ�����d,��,ȶA��DX����<Q�_^(˔��
m�n �JS%݈�቞l�DTp�mM����%0Q�� �!^&sq�B䉑7{���BL��0�ӆLPi��a����O�{��4*4��p!GN<�<*`O�tYê���hEq%e�Hvu���q�<qG�� @��!��1��mQ��Pm�<g˟i�NM���,�jy���e�<馄��Yn�%eF~g��h oLc�<��\'	;b��q .�<�PJ�[�<�ե	�B�.=ST�H�`g��jZX�<y��$C<\�Z���(�z�̈U�<1q�V ��؋@�Ϩr3�!�J�{�<��Uk�ɂ�K�[��X��n�<���Y(4�b����<B���bE	d�<�q/��%@<@03"[	I`@���#	j�<ѣ��!e�֜C�[�������|�<A���"�D�Y�OB8m:l���x�<I�`B0e���=y��{Dv�<	 Z�9�� �L�r��C�-�q�<���s4�7dO7l�\ׅ&�y��R�6�b �a
d�=�F��yMV�Z��p��N��] $ɸÃ���y"CL�nr��Ѥ"�D��ț�y�m!7��0$,
��>M�����y�k�,6�<aQ�/�'%�FŰ��;�y��W�i��k��� QP!��
"�yҀȦ>��A����~i�,��[ �y2�ܜw�$�G�نq�
Lx�(�3�y"$�'$�r�yW�P�5?j$�A��y2���F��E����'���2oХ�y��6@%����s�c����y�iξ	�$	S˒��:��'n>�yRB�u.Z<�hU�icbh ����y2�@�"+6��K	R�0�&����y�Bt�b��9��� ��y��YG0Xԑ`$��:Q��]�y�+\�(��jg�ڢ�:�#P�I��y"n�'7&��A�J�v�HI�N�2�yb�#k���	;?�F<�r$G(�yR�ɂ?ɀ�`H�8��P����y"��Y11,��g�"�҃�5�y��#_���+�.E�3)���o�=�y�L�J�&�s���e8� ���y���2AvB��!�z9�2�yR.�!%Zઆ��Ԋ}�#�
$�y�ρ�@E"AH�7�qx3#�y�ņ38�@I���6)�5����y�$ñU�x`;U�D�D��MY�D���y��F.aL��beT�<3�������y"BN�4Ƭ����%� ErQI��yO��a��t`��J���	�Iз�yR������C�ȟS���F}���S�? ��@b@���Xy ���V���6"O.E	��]"e����d�;U{�H�"O�%x��LY�t��`ߎWZ��"O���3�T�c��µ�߿H�|{�"O��"ܱ?��H���.NCu���'.�'��'BR�'���'j��'N(���$F�45����7�AP��'�"�'���'i�'��']��'�X4��E?/.�ٚ���9e&X,��'7"�'�"�'���'A�'6��'Ф���/��@� �b�x����'���'i��'���'�"�'�"�'��⴬) ��Q��̇D���h@�'���'��'�"���7�Ov�$�O�����ܘe��y� K���x���O~���O���O>�d�O��$�O0��OP풑��FYQ�O�%��a�OV���O���O����O*�D�O��D�OJ5򡊡���B�̯3��U��O��d�O��d�O4���O��D�O���O�����V�yH���:l���$��O��D�O��$�Ob���Ob���O����O�\H���(��xӷ��&/[�0ʱ�O���O����O���O��D�O��D�O�!�M1a���cH�%@ʭ�M�O��d�O���O���O����O���O�A��"�5t
��3�%��O��D�O�����J���?���?Q��?�'$�A[^�*Ť޻'�X��dF�?���?����?���?��xқ��'��"Fl�A
ӀEV���ٔ$��(ʓ�?�/O1��I��Mۑ��;�n��ϳyJH�$mU1�`��'�6m�O�O�9O�!o�� 5@$�����AM��Jd���^jl�ڴ�?����)�MS�'�b�m�����-��d7_�t�S���
���a& U
1O���<ى��]�Mn,��ɝ�+y�
� B ��n��C�6c���
%��y�K��re�Wc	�5iXp�f��P~�6-
����ə�m�:6�d���,�"jh���	�"jch���u��������0�&�o���d�'[�5j�[�|���'F��T˃�<�.OƒO��o9<��c���ՁY���<�,�3�"b �K��bN�I�M{�i*�>Q�<J+�A:C��4O��X!�~҄**���R��3��O����s�����	��	��6܎�˥��	5��'��IƟ"~ΓK�:I�e�r(^=	"�ؔΦ�͓P��V����Z⦁�?�'P�.�r ��)S�D�(�(Ŭ�P$�gQ�f�uӠ��Dݚ6�$?��(�2�D�2����<e�SȐ�2M,ջqG  p�m]���9R0b_&.�XT�0� %����m�(���B*W���;B��K�K���2������,��Լ����Y#`m�ڈxA �(/�A�1��$�P`*���<�3j9���b�o��h��#�&Y���8 �L�0��G<���riT=3?�0bLY)�T�p
�)m�neS2.��up#�B6��(��jS�\a�Lq��Ī!i�|�w��=E��cvaŊ+�\/�����L����ʟp�	�?5��O0����P���#6Fxd:��i}B�'�

�X��͟D�b��K!X���.8p=2x��œ%'���A�9��7��O8���O:�Ɉ{�i>u�"qld"wH�D��aR+B�M˓�_L~"V��$?�П��o�K�&��#�j��Q(Ѿ�M����?���y1����x�O��'7.���FK�z�JNb���0�>y���?Q�O��?���?Y���:c=^"WV[4�rp�9(j�V�'`\h#��&�4�B���Oʓc=Υ��g�5��D�*9B��ųi}b�M���'5��'�2W��
�!T�q��Pz5�M�>)k���tX�O<I���?Y�����O��#d���3�#ύ`=��X1� �"�0��$�OP���O��G�T˗2�^�1�FI#/|*��ʋW<�1Q���	ٟ��Ivy��'e�jL���)� 01����ǂX�#��W���ڟ��Iٟ��'��݉Ќ8�iL�Bl�"e�]NF�j�%C�L�f�m���$��Hy"�'��U���O{
D�E@��-+�=R���
/LoZџp������I[)촓ش�?���?���
�|bD�$%\�p�"�?m���q�i�R[�l��?��SoyBB�	���4p�X��6���m�8I�)��iW�'�����Mi�b���O2���B�	�ORY��F�IV�PC�+�Q�1+�)�L}2�'��Z2�'82X���x�IړD)�����T
���M
���F��s2�6��O����O��I��:���Ox�$V
S� �&��,9G��f��J>�mh}����֟���D��T�'�y�@�T��-�!�\�k���iP�g�f���O�P�
 �l��$������Iǟ֝+�4�#'N�ڜ����`G$7=���'@��?��Iӟ��I�*ٶ\1�K�;;�qF+OW�8�۴�?QN7_͛��'Ob�'�⪹~��'�� r+[�,r��+ƀ��9��� �O���`������� �I��Iɟ�"1�ͧ;N͈�E3�RQ���)��4�?���?)��;t��qyB�'<�`�Fm��͐�P'��+�n���ì�y�\���I�d�I���<����شj"����b����N+��Ђ�il��'�b�'�2Y�l�	�f�瓤'���x���+���rf��,:��T�ٴ�?i���?���?q�Xp��Ҽi���'&�D���v�v ���ˣvtd�
e�����OP�$�<���8�'�?�'�����i�0r�b��B/Ϝ��,�ٴ�?i��?�� �6�i�b�'z"�O.`T��+�6q�"c�k�E�f�e�`�į<���r��'�?���q\���� `%sRJʥ�*���2d,��h��iO剷͊yx�4�?9��?��'s,�i�ʡ�ȷ^f���7.���CBbӖ���OD3�1OLH��y���NW�܈�H.@#�X5���p(��
�7��OF��O���b}�Z����DSU���˜�w����2�ԥ�MS �t~2Z�X�r�$�� ��nC=�@���U�ob��iU"�':rɶp������O��I4W� ��wBE�"���Eƒ_��6�OLʓ|2h��S���'�B�'� ���HS9e.��j� c��88��|��DEj dm�'p��ҟ��'qZc) �H0����0!x���=�ʨY�OԼx�=O���O*���OD���<A�b8^!.lѧGF�Eq�ebt@�55��#"R��'
rU��I�,���r�"2�eO0�pV�K
z� (�aAg��'b�'�r\��ԩ������dV�8�(��Y��} w�� �M�.O~���<����?���f��(�'�v<��D	�vK ��`��6\��4�?���?��� e!��ߴ�?���?�l;C
�U�� �.��)+,a��i��'a�Z��	�<��8�	�-�4<ATc����|ք��ң�ԟ$��ȟ��I=WНZܴ�?Q���?	��/�5Z�eP�|閑s�o�CߘL���i�bP��I+B����OX��|n�M̑!��#m@�%C�N�C�7m�O���C�QE8oZܟl�	�d��?��I;s,D����eݴ@�6L��-R�p`�O���ǋ�����O��D���9��僖vz�e���Xy��˒�[�M;�²���'���'���O 2�'D"�]��(X�g�K�h�`	4
Iu�7-W+4����:�4��������w�~�x!	U�q`�<��kƄq3 n�⟀��ܟܠ����M[��?���?��Ӻd쇏W�����@�B����R��Ԧ���[yB��yʟr���O@�ć�:�b!�t��(x֥C�')db�mZ�飣��M����?���?�^?���n��@y���3���/yP��'��Is�'���'S��'���'�����.}0��)��i���(���5I1�Rhs�"���O���O*m�O��Iʟ����
�*��*r��s��:�0��� �	��<�	���I�$��-<�M�t"���MR�R3�^Qc�߽n6���'R�'|��' �	џ��D.z>0iˋrP�U`s
�%--D�i�iе���O��d�O�˓0ќu������.#�l`rk�:vB��i�Q��6M�ON�O�d�O�5���O2�'����O�U�R-�%��2��`�Ԧ���՟(�'��2��>�)�O��	Խh��t,"'^MC�l�RX��%������`:�(�\�S��K��l���򥝣[P�dk�%�2�M�(O�)��æ�3����d���5�'�䭪$MH3E�:����Ò~?R��4�?a��"��P���䓿�O�VCG�
�[m���� S}�,xh�4YU�hiF�ij��'b�O5nO>���x���"C��!�uX�m�jn��s�)�'�?�A�N�JW��u?V��W����'���'�ػ��<�d�O�D�� i1�J�B��B���Y����-�	�Pc����������+�n@Ѭ1<\
�h�Aݲ�(J�4�?�V��mN�'�'�ɧ5V� wn����nI�$�G�3��$Zp=��Ĺ<)��?I����ޔB�T1�h+e�T�G�p��da�K�U�	����x�I�����)hA�ǆ�YX~�0n�}�|��T-_ԟ��'x"�'rR��AQm����¼y�<�[�+�
��a�%����ON�d4���OL�DQ�o_�޼C1���f������E�Ӿc3��'���'�BW�Ģ�F��'+�T�˱�=~x���M�hY���iX|��'Yr��r5R�>�oN�R�F��)�0�
�C )K�����ܟ��'[n��I.��O~�iLS��̋���z���e�0"�%�����Z��p��%�@��l-f��d��=JR�8�1��J�Dm�Ly�$g�26�ET�4�'	��B#?��GՇ3Ҧm�B�81��I�禭����`;g��g�S�'W���$3)Z�y!�?<#Z�nZt�8{�4�?)���?I�'̉',��9*^�i��>I�l�s'A�7|>7�R�?D��7��џ�9�O1�~��%�����0#��M{���?����!��i��'��'�Zw@U�Ȃ3���8!,�� ���9�4������S�$�'7r�'�l�`����"�(A�g/�"�AfӺ�D��w��(l�˟�����l�������0��J��Tl�k��ĸ���!��>�!F�<!-O(�D�O�˧�?�DIJ�<x6���o/0�����^Ô�P��i���'J��'z�����O�E���M��A)��~D鷤��O8��O��D�+�"�D�O��D�OX-C��Z��#���������I~��p���M���?!��?�����O2��=��f��N<$�`�H5M�4��M��g&�p��d����딓Z�1�SY���N���1t̗%�XI�⦂�;��Pr7�V��1萉�a؟xt�Ƕj��b�	�Gʤ�����Y��Lv��ņ�1N|2�ي?]PQ �fޤkLD�y"F�*iQqrO�.jJ�LQ����>
�P�g-�\Y�e��	O|�(
 '�o
ޱ��H��P2T�Fȧ
fڙ�gT �*)9D�	\������$T�@%��I0 ��5	�%�И�iԯ<.��p��k�2�+�Ob�D�O��� �+^�I�JʪCP��5��=>ަ�����4�n(['��]j�T�3mX�i�c>�)9�-�ҏB�7��QH��1{_0���Բ��,yrlQ�B����gS0�j��1��w�|��T �!���H��~�~�k�+�O��:���O� 2��r��4j5�8��d�2O�61�p"O�8�f�ҧT� �Am�t��;�ɪ�HO�	�O�� �X�xE���s!^<n��jd��O��G�to,��b)�O0���OP�D_ܺ�Ӽ�)S)k!�i��	^7�������;&����<�K��,=Ȣ�g�'��aȅh�.Z|��6�yb]rp��O��H1#�"zL���ھ����D]�����nL+Q��iYŀ�+`���uCR�'UўX�'��5�9"HTh"PdX��]Q��*D�L�e�M?�APt�x�ʭ�D%��HO��OʓM$B� p�i�-�#���j�� ı�rm��'%b�'�򧙄[��'6���!��Dg�:9R�Ҕ�����aW��c�H@�Y�yG�1�ROF�'r���S�������I�:>����Q���a�B�
@ ���S�Oo06-�f�aw�/�ĞB�o��h�LNn�nICb��U����"O8Qj_{�Jh��A��v�����'�ў�؄�ܨ'�	Ad�!���R�
b�p�ݴ��dr\��S?��g��� �U�0% D��wO2!�a���25�'��'�������;C���@�>CA��T>�IA-E�����&iP�0��)�+"th0��T6v�r��Ñ4��'j>��,�?f�1���
BO=Ey��q���?����ܤc2�$��f7d��sGǟ0�y�'s�l�Ď	�7���	{Cl| '�'fNOE��o��~aq �S<0�0{�2O������}��ڟĖO�jj��'H��'J���&�6�Z��·k1��q���v,hj�o�27�<�m�ɟʧɘ�?�d�������	��y�`3�If����� m�d-j�H���O�1 `��k-�9�� ,J���[�Aقƒ���Ot�S�c�	�*`riS���F���Ł�9-�C��;'er��悒}.�q�'%�*WV#<��i>��	�*� R.��)B��ͨbgd��I��,-@��$)L���	ԟl����uW�'�Rn�����j^�|㐡�"��~��7��>�� �.i��a�g��(?�<1TILS?�Cxx�,R�� �.�l�� �&�z��㦟���2�'��'�2�'��	�7���m׹-Y�`�Š�L,<B�0W��PU
�0O��z"�E��z�h��d�|�/OH��6��̦5	�Oq�\�3����!c��ӟ������	<Ő��ݟ�'1�>A�SЈv��-[`�!C8�X�(�R:����☯3z <�"N�R葟���ȴ"�<������ꞝ"p�D_k�1tM��b٢ك���46B
8P� �C�<����� R2�~�<��U��{�>�pu�����IR"O@�,�}9�22�bv��$"OP��GI�	pD��KG�N�s<>=(�5O�`oT�I2"-dm��4�?�����)��s�h|�d��a�`�����,�j�p���O���OE��,�
'����gh�W�0�����tiP�'8#��A�SS��zW��!�(O@�37o��8��R�ā�`s8uST�Ҽu��U�1�^�;�ְ��d@�_�t�iI�>�.-!�{�$P��?���J�`f�ہu`J�C�^��B�O��y!Ѣ��C�(���Y�h x����_�I�$ˢ���!�,w��L����kf�I/&Od�zߴ�?�����遦p0�D�O��V!9�,A0�	u���f��gC@	�p��(IS��Y���p�"ٺ����w	�Iq�*!{�b�R�;^�p8�`�"s�1Ӡ�4&;�9�p��ߺ�4I^�b<h��'���D�T ��>	�\������%J����?�W�|���'eLK��A���df�5E�����']�혥�-m$���ʊ2
*�ڋ�$�z�����'���1��˔$��������b�'8���x�1��'���'OB�u���i�� A��P.�	�!�4qt+gb���C�G"�O�ɣ�g�*��U*��a���7�Oڅ�&�'�B�񓧕�0�|" A�-^����'��A�n	a{�ںAh ����J���$�󇁬�y¦۱t�(R�A҇T�H�3#J��i�D"=E�$N_#Lx�7��s˞HBbhI�uk!	����i����O4�d�O���O�Do>=pA�������.-|U�P���̄fd
�q�U�7H8@�cK�4�Q��DD�#�J�!�֯/�N|�N�ki�a;�Ƈ3&_v����;x�(�"���)1���%=8$�4�b�Ol�q�8��E	��c~�<�G��vB��E*��B�ʈ֊��!��!V�d��1�kNYk��X�,e&�0�Z�n�:��t���|r���v!�6M�O���|�g�lF}!��"2��f�V3T����?)��e!��2�@Q[~�}�Ǫ��6W�� �?5�G���PF�_!�f���8�]`P���.�F����5�f�s��ԏE��ĉ4nO�!�t!ڢ�����VxQJ�`I+�OPxG�da#1�`�J!LN|R�y1k���y
� #e�1%��0��'�}R�'��O���E �3s�����m�e(!V7OڠU�Zߦ���П��O{ظ�'	��'��]��l��ː���I�G$�{�I��	k�T��B�����6��'�Ͽ�&+F#����`L�+Ў����ϐn���(8�m3S�ܒ���,��Xs
w��w��І��F�r%(�
�!r&-kQ�ml�7���O�ٺF��Pű��)�\�
e"Ot�d�G�f�N� 	A�"�Mzb�I�HO�	�O(3�oe��Y�\�R��A(�OH�dFo"�$��	�O�d�OF��\ߺ�Ӽ�g��&�b �siU�4a��h?i��Kق,P��N�ǰ<�g�I�n��w�ւ����G�;sXp-���L'���CI�m|��'qXQ��Q���r�:�����s���4A�������Oܘ��I�L�)�voL�r@�����]��B�	
]x�2�e?@s�H�A2RN\+��4�d�O�m��e���8�#��X��&F$0Nb<����͟��I���raP��	ȟ�ϧ!�\ dG]��27��Q����c��y-�b0s��3vn�Z[������I�&9�3HD%A��	��[X}t��FU�I�B|�K� {X���Y�vT�9G�I|�t\������azMH5QK@ ]��D�2D��c��
�V(鷃�7sr&��.D�\(&��h����'=2�Y1�b�\q�4��vT�i���'P哪z~�U&��jv�=���6�RXto���h��럘Xa���@���u��5Zb��Ԋ���)?(&<p�E�@�� �9"�Q��Z��? J��1�P��X�'Q!�" �1�W�u"�@4\� �M�/؀���*�K�ɕ-؈�#�|�S��V&my����T�2��V��z�<��j��%���ɗZa�5��m�(�L<�櫙�|�ny;�,PJ�0�ѣ��<1Ī�y���'R^>-+@����	�\����#P+n(�$��5��鳕K� l�3� K���� ��&l�ܹ��֟�b>�NЃ-�Z�h�jC( pq���T/Mqy�hY�V���P%��{��Mc���-��ai�� S����1,G��S@B<ns��`榅b -�	��M���?�K~2���?y��"Y��Y%D�.}��@�uM�f]���?��2��(�F�] n���9���Dx��!ғ9̛V�'u���!�Մ.@,8����]��D�p�'��'��3����'�"�'m��m�������K4 ��+�!���0m.X!c�!pf��"�AV	Q;���7�	�����(O�Q���<;
����W�-�D+T�m%���3���vL�/Z��	��9�dq�c̸L��� ��V��e�0h
P		�
`�K��j���k��:��6�''r�'e��'9�w�b�R��YV�.y���T���X��'�m��	�X-Z�ye�t�d/ғ_����'b�	�f^h�*�4H쐘P���̰����45,t����?1��?��eF2�?�����N�/YX�����GNhn@U��)^������0�&�r��'�B��휦N,���d1h{�l�f�����bD�>�����J~#?�H�ٴ6����P�(����"�ȑf�y��y�6�p�!}.��Qe&�
\��C[4�D�GxF����%��=ϓ1����|�H�7|p���?�+������5y��p�����^x��`6n�(�T���O����_��	�#��.@����V�� nHY�Od\�JWa���݃W&^�-(�a���䔚h�8�%�<�L]#ԀR)\�9FF�1F�x���{�P���e��6Wx�Q���>V�O|�Qt�'�@7m��]��P��";w��	���:o�fݙA�A�ri2��s��b�KG�	�.�.j 4+w�.�O��&��1a�s���2��e%��h��l���g��M��?q)����S(�O��d�Oܹ��jϝUg�G(T+<}�_:\�>�YD㌥B����!<.��O1�Wvy0茨����W��*E^<#ᑚ�,#�,�7L��)�b�>��i3�5$�6��ߕkA/I�Z8��b��t���W�E9�d�ɱ��S��?Ye�Ku5d�j��Ȅc�D��Gk�G�<����GX�Br�>,�$�B�A�'ľ#=ͧ�?���� ���L_S]=�D=�?��fe�(q���?���?��Y\��O��T(n���4���Y�-B��N7S�L��fV�O���Nݿ6�p�z&ޟV�Gyr!�)%��Е�>V�Z�*�I ��!��ֆ+UI�(r���OɸX�t�Zٮ�GX��iw��3�P�JE���('���a`��O*-���.��"��#��#���C�I/*�T �N�V�8��5���.���4�(�O���'U˦�hg�ǹ'�XI�`k.+��pSd@˟��ȟ���%�����ͧxt�����D��Ę�ˀ~��Խ�x�c�7yf�H��c@$d���Ӎ�$-ҸIK0B&}nu�i�f�Z]hr�\+��AdFT�+��0a&K��C(����t��O(��'0�7�L�1D|9 �װ+��Ejf�\�	�!�Dʅ`0^	�s�Ƀ`�b���Ύ�"lax2�)� ���3	��q�ȍqm�p��?O���>!�!�!#2���'E�P>ŪR�I�_�2���Ŋ���#@��X�	ܟ8��4�ؤ	�l��i��c�b��U��?�p�Z�V�d` ̇��,Iç?�"��p��4;���&��#�~,�a�<'Hy�Sk�'v����T
����6����d;���O�<E��g�����H�<x�^p�!�٢�yZ��4%��EZ���ÂE�{��B�iӉ'�(����8���P3���Ԁў'�$���Mo���D�O��':|�A���?)��_�fd��F��~��[�bu��zU�K�?�y*����`X;ؒ�ˆQH\C��*Bd^%Dx���'"ֈ���X.�Jpsa	� !h��$���jZ��$���OȬR��	�:�@Ȱ �T�N�y�T"O���0 P��XE���$

���HO��O�B�iR�2L��,ڄc�J�YRl�O��Y�Q���qҌ�O�d�O���ĺ{�Ӽ˵��3�̑��MBn�r��R�xZ����"|J
��5��@m,�'{�Q�$�q�%��p�"ɼFްyf� <��)q�-
g��c���Q���si�i&*�ju���3��kw�AI�A�0jC��d¸�D���O,U��<:�f|B�l��r�B<3ׯ�'o�\C�I��:�ⱆ
:3�4F�	�P���4�l�O~�ҋ�æ�?t=���3�B�%9���u�����	��d�I$c�5����p�'VX�3HܘH�q0���&Q�8*p��A���D���7���P	�b�j����P��*��R#�'G�j�R�㖄R��A��Q�Y��K�Q��Q��$�MK��N����H��Y&.�����D�<a��1~cjA	���e`�� �~�<���j��l���J�t���l��<Y!�i��'a�0X�c`�����Ol˧Y��b)�d<�@�ʗi���բ���?��?��ԣh-�8�/�[jּ���U\�FD4�����g�G�2p����6�TGy�G.�H(��a�}������ݐilT�0��N��y���(b��J#�]�&��Ey�ޙ�?9���
<Dȓ�M�8�2i@��bC�ɓ<�B���+^+`�0=�'Mޣ\����C�I�:���Y@�#`@�c�� {�ё�4�?i���۱C���D�O
�dNw.���V9#��i��_m�ƨ��aN�v�2C�-Jx,���|����0D�v(�*���j�&�e��7mJ�W�Z�޹z�
 #S
��	�� ���w��}��3$��S%R�/���س��&�r�<���O�x���2vnPl���F�N��.0D�y��Wqld-0bـ�nh	�.-R����џ����,�\AvĊ� ��4Ag'W��ɐ
�*`��c�ҟ�����L�	=�ug��y'¨>�(]Br-�i�~��c��f<�B���#��QJ�,K�:C� �O���3+ѾӘ'h��҂���I �̅���qy������Y�"�d�CNV����g�d��<1D��4T�����փQ  K1��?	c%��?9�ܛ�����OlʓY�^��2�0s�j4HwHL�2'��<�ߓND��EU2*f�{��ζD�(8ඵi��6m,�4���<Y�DIO�Vo��qv�j�y�2q+�F[��R�'VB�'�\B��'Ob3���J ˕:��X��)zd�H���B�#�6I��F�>
�L �`�>@�F~­��z(ш]5$H!�G�ʹiq�3k��}kYM��ܚ& �$j�6QSLkܓb����I�M��`V!�:${�ꂞVF"i�j�`�<)���/+���6��B(z9���Y�<qcH�$Nu��I���l�v\����<��i��'e�<2fgq����O�˧3����%���~(0�޿[H��jO#�?	��?9�@���?��y*�xzf�Y8C�\y둎���tC@剦38Ģbg�Ӓ,��A�a�;1]�vΔy�'�D�C��9��>I��(W�uF��� W�b#��(�:D�@+Ƭ6��+6��'Jڡ{�#<�O¬%��6GG�m5�=�6E�@[����z�������MC���?+�f���/�Ot�$�O��K��Z)V�D��n��3��+Uo�.%b�b�ؐy��xY�hG!��'ɡ?��|�1A٨A�'`A"h�uӴ�2Y��+f�}n�Ta�@,]� �36��x�j�C$ O�Z�Ͽ�.C*�����5r��b��~�:��v�ɧ��c�%�^Pc��V�sO*�s�����yb�Bt��#1A��hh�J�j���O��Gz�O'"Y�j=ClL%YH|ES�+əg�B�'�@�uN��S�"�'���'�~���ݵ$��4R��Է)��ISk�.=b]c�9a����߇�lm�`&�?i1��D[�&P�rF^�p�`��@�. ~��S%�.69;'��+"B�JП��l��G�1d
u}�**0A�QرIƏdf5x!�O�~����?���hO`˓I'�B.�d��$8�隀*�x�����?�!��	~���q� ��8�(
�e�ğ��'��\0&"b�� ���/�'� a��ԘR�`Z��O~�D�Oj�W�0l��D�OT�;"�e�� �;�l��B&@�6�(�0�	�������S���r�SNn�	0�6}��XxB�g�<9�ǥT���t)�sRYP���Y(E���'����毝�'vN��Tk�P��|B�'����?i�m l��xWnгF^L� �/D�P���o�f��ŌG�@��3Fo��
ٴ�?!(Ol�JB�H}2�'��1+@`����96�B<Hh�&��L��ɟ��"L[˄��<�O�1�GP�f��@��ou�H���d�<>`V�HP�$�"�@�&p����[$K��<��M˟��	؟��If�t�]W��KN�I�Ĩ�&ˇg�b��s�,�4���LP���K�FPx��*�OT�'�d�A�s�F)���<� Jh��' �3�M+��?�*����@��O��$�O�x��V�&C��2�	ߕG��'	�5�ej����5���̙'J�B�A�O�1��E­A���t�̵M�2f��'�Eۛ�6���B�=z�؁2��^�?a���!��qJ����G��a��l�$��F�<���I�;}�	F�'�N�O?���67�rq:@%�J�D ����0�!�V ������w���_���Ћ�4�b���>�� �B���k�5��#�(�$�O8���$�6.SX���O ���O�1���?�;gt����B�O�<��g�KX�; �	-1w��6K��ɖfZc�1.
���G�G�Ƶ��ɏԽBѧ��~zfY�Dϔ8K���0�ư?I�شs��	+�m����d�8�t��unĬP�)[��Xt�$ܯs<� {�"Ez�Q�@�L6k�8�j�Ny��I��x��'�8:e K�e�l���^�j���e,��|:���dY &�bun� ,��re�D�,��PN�,j���	ן,�	Ο< ��X���|Ң��Ph��ahڽ�B�#E�ڶ�fE9� ��	z)@�`�vɚ��	�1��-��NԎ|d�8�C/q��e�J�� 
Æ���pl�=a�N�k�*O�	qO�%x��'��6m�/ .��C�ܟXXTk���!�	�X��Ńԝ��x�B��B!��"g��H����f�j�XBU����P˦�&�ܑ'$�Mk��?	/�\Hb�Ga���a��j�(��SN��2q��d�O��� �	��+"P�S���s�c�Z��T��O��X���> �D���>rh����d�!_�ʈ
��ƤH�h��K��l�A�'��!"��>���G4O �j5��6 ��O.�ju�'_�#}R��A�!�,!Qj4y���@*`�<!�O��Z,��0]YY'�@��O<�dA�a��#̔.9�r,9���<�UmT�1��Iڟ\�O�,����'*��'��ر��L2�V\�DkE=TWy�D膇,$�c�H9���S���'�l��tA�2x�y��N�"':����ze��Sdʇe
D(2��-z��AG��;<�� 8Blg�DxB��E�P������?���?�����B@�h%؁�QdM0B��i[����y��']�}��$���!bmS8:P9��G��O�Gz��OQRh͖-a\T� !����r��Bm���'`�P1��!���'�'��֝������Ґk��rs�����ӻY ��YF�����2\�=C�#��|*�&ʓFr��	V"Ҫ`�S�0��'��\U�Ҭ��3�8!�íT���ܔ\un��.�����Z7�yzSFՁ?���9G=iH��S�28��'��O~���O �h��[BK�y6\b��\
�E}2��)�(����jA9̋�*iZLb�4�F�|�O���T���u��M�%j|� �F����f�E��H��I���	���$E�@�I�|r��I:`�@[f螆1ݪ@0�ӡ`������ y9&��3��{%��2^t�x� ĂjEh��� ��ʔ��YpMK%�]��&Ȱ�	E�LH�=�E���mqqOŢS�'���.p�����r#�D�F*�'��'2�O�Ӄ�V�[�j֠bw
���C�?!��B䉊0买�V���Ks�ЉK����'�M�����M9E$�o�矤�	Y��Bj1،�OF�6�бp��*$��4ʦ�'�r�'n�#!�';1O�}p}!T��1�� PE�hP��<��T�O$�2�
E9Af���Y�z�80��$�3,%ҧ2p	�����ۣ@��/�@-����Yb
��a$Π�����Ā���(��x���9���M?�r9��Jq@��l�
@�FxkpҀYB��ȓ@�&�9ff<ĠPS�'X(.Wl���쩲�7B0�ԺP�0J��<�ȓ OԨ�RD>�&��3�	a+ 4�ȓ}�J카����X`�O7�V���,���J[�*!�#A��_W\���S�? �aR��þ?W��`��=J���D"O�Y��"H=���V��";�D��F"O|0��ϗL���0�eϏx�\�y�"O^�I��7�<dhsN�0؂��"OJ��#O+N�>hW��U��B"O�,��N)�`Ba�M�p�sT"O�ّb��`6�5�*��P�"On$yA�Z�_4�������{<�r"OD��7"�p��P��`�"O�lE��r�д:R��B���"O�xH#ɟ�6e
�ʁ��Ŕ�yB���!��r�/�xk�=��OQ�y�	�358����N?v��;#���y"Ox��b���ag�UJG���yr�փn��+#T�*$I��5�yB��+
vpQ��K�T�	��y�BP:	���'���0�饇�1�y�NDI�6��`M߷~;8qC�l��ybC	�A:�{� T��Yr���y�D�f�Z(��
7�2��B�V��y���6���ؓ
��8��"Z�y�MQ$s>�(d�E|�R�-]�y��5� �*r6 +�x�kы�y����LJr=�����w�ђ�hІ�y�hN#U�Q��պk;�p7(A�yb��%�|�AG�_3b��E�]�hOp��i>أ|���<Y��	�lX`%�qڵ/N�<i�KP�'D��+2Jd <<
�ͦ	���X=�FȁN<E��4r��²�'0��T�,�!��I�y�H��}�@��ăL�e��h�,����a��Oj,�'z�O�D0m�d$����-��F��h ��y�L c��n��|R��O�I9�M��`�
N�Ip���lk��G~�� �a�b���-,O���@��y�\@3a�ڢ:np�8��;���S�S��d�	���~�'�$���D\&����EI�+m+c���x"��874<!�
[�H'6�;�f� K�x�q�ONm�s4Od�X�D�O7�:2�B�@�_x�%qя�3�0>�w$��>ԞH�
�C1"|Rp�[�
6b�钤N�K��9+2�$Y�
��mz�}Pt�K�J�b��N>qf�:���6�5����#f�'at%���& �$ف�eJ*���O����͎/d�5(&�S�?�|�"暞x]���FNO�"28D��K�wX���e,�~��Y��YH��@�c�N�0B<�v�.[x,���ɔ'�c���bh��AR�_�A�L�O�F�w�<f2�3n�4�PY��'����B(
�a+0���F���Q�"��:�\�Ʉ@*x����DL%e�����&p��w�ƞJ|��)�h,K潫Dn�"�<$�>�u�X
O�*�㲮��-��Y≅Y��Ab�ݱ:�ЫDϐ|�*c�ЩL߰<-*X�!�a��)�k;�; H�b@^�<��%9�!�10|���Aa��ɇAN��2˓M�ڄ2fC�T�#��ݾIa����]#�0�{D�OR���d�O,�z��ES�B��7���le�����BJ<y�Ǜ	K�X(*&F��!^�m)�G�}�ax�:O��Vf[	>�����Ŕ[*�
���?W]��F���#7�AX��q�-X�(tJ	;vK+B�*���xSN=0�� ��~� EF6���!�M���i�����i'�شZq�F��<A �>I�#�!B����c�C�I�+�IגG���#!J��c����A	�x�D��&u����m�"8*eh�R�	rӬ^�v0����	eX����Nж���K���\@R�H��}� e���=qS��%H�p�AE�9;�q�խ�'w��S��5F#�&����uj�<������>y`��heA�lB�#Le�gBşnY����B -&,ayRǔ�]�;g� �XM�p�щl���Xv̆�?,�i�p!q�2#=���T�l-9b��?VO4e��X}�@ %�h#��H��������p3�	�[�� �,R�A�d����kx�i!a��R���L,h>(�����V�fqɅ"�?^N�����B�'���c�'=)+�5KP��5������6��Б�*J�D�ӺGzZw�F	s�̀:s��JP�Ue��1Te�G]�}�w��u�
bb�K�&�-#�!/O�@Fz*�n��=R��@ ֢d�h���  1�H#f�OP�$)A�M�Fq ��^��X� �aR�'E��}KR�۵8�����ɿx0�Z��a�$+���(\C��^��%@�9��fJʵ=�m�O0��ń�+� I�,O�X����9Ox<В݄ qlɃf���1�<�+T�+��(�9P,�4�'8ꠣq ���O�P�6+3bC5X��/S�4%��*3�'ߦYkB|��bBdX�F˼���gy�,	%\��y�s傲X�xf���?���/�Op���T�t���"@�q��s��P�L�ğm�$��B����}Ӻ�禓�B$x) �r֭�hA�02�(C��'�֬�`Q�p�������F:$����wN�e�t9{ݴ|ܩB��4WsΈ`3��M;��0�
2KN�p���O��'��]�q(H;bF(|��x"�@�6D�Q��ǉ�~�G�E��O��K���>�
�w�>";zU�Mҏp����Л0��!��'�4�J�ɍ9~S�� )��/?����[��
u��b���7��a�������\yJ?=r2��1���tfB�[��(F�;'+�[�!��a|B�Ȫf���H�~�Q ����h*O �BY�'�n�Yɟr�� �ˈx+��p�5!����Ҁ�KX�!�*�v8�	W�Dt���7
����!3�y!����M�B�ARy�΂
�4�bq����Jc<��h�,�FN	��L�XP��y$��kD ���9���i@(�$=d��e�ĪEU\�3}&Y'q4��$��9�ܽ�WIT�~��t�����
"2������hO�]`ꀚo�:��bǒ;o��+Bɥ@&���S	k�,���F���'^��M��mR��{�^pIRF8�	�p@�������5|Ok�܍p��e��`X�.'���w�P���FxB#�'�
�B�.RV�T)� ��0���A�C�ay¡B.~�bhc���<,��M�>p@�Uc��*�R(���8.�7� Q����,ղ�R�1�\�Yǿ�ʑ�'��l�Z��5̌(L8j��xRc�9pՀ��O2qd�Ö��|�O����E?Oh��� �[	+����@��$��	��R�:h�щ�2x�����=�<D��H�mJ4�P)��ǨJq��G�O�]�eC��*[O.�S��NO�2�Э�w�P+��J5�M�+k�%*� �=G
�@ߓ2�Ȑ�1��*h�������4r�FXDx�g��$���g�*:'�Q*}*�|��a�(��z�B�:X߸x��-�V��СS�ݰ��X@Dk�R��Q4C�}b�i4�O"�0c	�1�H��RO�,�Us3�!&���G�ϺX��I��,�I��'����6�ARS��!B̔�\y��[�	I;�D!7�	�L�Ȇ�ɐP�\�)Ć8t���2?W�-1�(�
7(ۅYYP5�K�'T\��p헎N!\�8��S;J���A��?m����E�I<����?�\��t�n�'�R���]��R�YC���I�L�Kv&U-~���ZT"���=�E�OrR�(��JI	"@�� S�[8jt`%���l�!�דZ�XH��HF�vV ���Ȟ6O5�`"AkX� 0͈^�)��\�rȪ�E] }�J��Vo�{[�c�`��0<	RBՖ:l��F��DS�1�&�$ܵs#�Z�DU
uL�l�'�����\ή�3�Ț�6�Y��(��
!N����3�,�i3o�8�n���W�~����S����H�z��5�r��l���6���h��_�=	f̲��P�?r��pb�Ź&<|�ٕh�[���'�{ӌ�9Հ�������u�2 ����h_6 c��i��?�� �AH�_
����],�&T*f96 ���þ1<���Ԕj�Bl!ۓ7�0�X��޻�ɑs&��i�r���D�m���;�Fh�r���Lэu����.���� *K���n��0<����X�PXȴ�5�F���n����� ̎/U���-���Q�<��%�񦅡0�
�U��D�yɧ>1Ǳ[�@�B4��I� }��Fx�Sћ��'A+�/^GnE�(cU��#w�T�{$�Q��жX0R-�?�C�iq� $����4;�'ߪa(�iŪybZ��@�߅3����
�V��#��0>�S+?���Pb�;P�8R�H�U?A�'��➠�>�W	� 7��y�L�K��Ȱ�J�"e���+�e���"����e2
p~-�&i�8R���؀�#OD���K<i�H,Z���&��P���W5�%҃'���V��t�1O��R��4 zQ�Ia�Xqpu��%�p�:��R%���)��[\��Ʌ
����WD͗f8����L.g4"<�uE��S�P�CW$2�p��=�Ĉ;�U4en+E*�]���;f*J�z���(�7���+�#&�E�c�iE ��	�21xa�Am3\� ��+J>Bخ�'��#=��O�6�
�r�x$X���;`7+p�����i�&LO�:`�K���5�+�*.u:����-�������[�i�ҢR�}Q��'��iZ�JI�D+�Kx5~`�f䆙����$B��!�j���9�nG�P�t��<9�fW�it�K&��,Q"jP�2G�7g�ɻY�0]B��C)Tyd亣�:R�)���>�@��i�ԑBCb�% p��g�'ɲQ;0///N�B�J͛ 8є$�Csq���d$ĝk�!?ᚧ�D	�3�y7��G8��foʿG|���.���y����.v����	4r%��ҥA�A{�%`��#H�`a�}rC�r�Ȕ��C�&Q��L��I�;1�D��	[#���sB�?u����_:8�N	�F��j�bI;1����!�seZ��Z�A�@�K �#"xצ�YL<�M�`h!"	@^-�� �<��]�=\(�kg��9��\���D��gW��*�l�6��q�䧌fn��Ӧ-2�'@��6@q6jIV��<��OXM��b���
���䐋J6,X�
�x�9g-���phӢ5*�p�5���ƣ=�K������ҩ�z1�T X�j�0eN\|*����S������T���`�2�V�B��6�$0}bO�h�P�'+R��a3Oj����cN�[v�X5|5 �!g�'��,�e�
�Z�7���z��h���*�ʜ8� �w?���8OP���y����[<B�ܩC��r�ȟ�~r�</Ď0	��D�5��b�,���'�N0kCKϛF�� 	J�Y'�>��ӧzT~�ed�1A��1KW�-2��ת�?�$�;1t��&Ç:��h���_S��1uO�~_��*�&>���3�4f#�y��!��I�����_Ͼa��^m�����	z`����1 h��	�l����;-"���U#���'�D��O�Ex��n���s @4H�ŰS@ݴpn�A��W~���+�fJwI aqش}� EI��V/Vp(��#��[� ��n��<a)OlP�'4z��G�?1�7{h�K�iDjaCT"C�.�b�Eh
G�H���yB`>dH��A<O2%lZ,!<L�'5� ��4j��m��!R
?�<9:%d^F}re4LR����'s2�qB
��HO�Y��C�=���"�ۓ �~�!c ��;�1O~��'
�<�,�4�����ǁD5��B��2�R���Fئ9r��V�2�(����,XP�N֥R ��d�|+����4�M�q��4Al��|�$m��ɳ���Q�c����Mºe�m�0~E��$��(Ä��'{D������Hx��ȱآ��O<��{],����}�1O�,�O�H�Q$Y6_�t���_"6�0�ӈ��Mw�>7�:uC�ȇ��]�h|p&'�+*$�j3�iy�c��G��'��{�,��\A��Hَ��qc�'}<�Y��R���P狠/��@B	�'R�t��	/WB��!M޿&U�$
�'��	ᐣ>���� W
q�H�C�'3�Q��#T�2��Q�7h���!�'���KD_�q��0TH�vR@A��'���e@�m�� *7d�'i$�i�'.8����^+�
!+�,8+��4��'*@�h@�T\|��s�T�h�1�'�x��d�[�� ���&�&��Y��'g�;w��PU� ئ(
�r0�'xl�0�B#E �X��B�wk��	�'���rrㄛ��� /�vUhq	�'t\R���#Y� �5�>B,lS	�'�L��#��$G���C�4�"}X�'�ޑC7m�9����a��u�XDz
�'�(�+�NX�3a Ux�
�'�z�i`�2���zЬO#dj ��
�'�d�&� �ε�G��4_X:��'u�B �˝ �8���b6_�Ɓy�'���ԇʢ1����1��Q�DI��' t�8!�IBI��y�JE�Yt�]��'�4�pT���]S,Șyw�b�'rA`���(���@B �-����'K��)1Bω^h�۱�L�z��Q�'L��R��e�ȴ��Ԩh�Ҥ8
�'���`!�9.�m��ehܭ��'4�щ��-l��h���<L���1�'�ЭʶM�=,����Y�H�̅��'N�Y�&��&^8ʅD��1�,U��'���	aj[,���(`ǖ���'�lq�ŁV9c.����āZ��w�<��
�}#��j&m�>&�>��s�Nr�<�W�
!��Mף m^I�2�m�<��h�'3O���PɧK�8%���ȓ`�lh��N� 6����5�Ju�V�ȓwet��6�Z �� ) E��>ه�W�T��7�;
�ƈ��RvFl�ȓr�p�n˰BG��`cn�;�e�����R�LQ�B�`�j�68��,��]��Ze�^�GX��I��6[�����S�? ���ԓ>�,Uc4f�Y4�yY�"O��5#�l�%	�LDb �!"O���"���~ϘH0Hm�j��"Ox�pU�D!,�f������Y�"OV]�M0e�8,��	�0*���"O�;ac��a�4��@�@�}]�""Od��0aNT�� �<K�  �"O�႓ ��=x93"�\@"X�"O�dj�D����jF�x%�@�1"O�4
�"7/��lP��-��"O� ��#~�i@� �*|�t�1�"O���H�'w�h6 �<�-��"OV�t)�h�Ш"2A��p�Dڥ"O�	��I�fj�jW��.]]\ �"O�iQ���T�F�E��?pH�@� "O�)3j@�1X���M�~��E"O��[p��KD�9 C��r���"O�dZ���.��,��VgX�d�"O���+)��a@
�sN�(�5"OD�"x���,G#$��q�I��y�ܱnL���!�ǇF6���.X�y�]�uO�w�M��`���-�y�!m�慁@4<��)������y"�[�O�ض �<������y2&�INM��kA0ڍ�G�͡�y��G��چ�N�^�
=�ά�y��� 	�i�] @t� R�����y�\M8mx��ۢf�f���L��y򇛿\B| ���1����ц�yr�3Z0����8"W:@(��/�yR�Φ
N��&ʪ�:T�3����yf@�:NT|���"��!���H��y	F�I4&}����&_-Ҡ�a �&�yR�\�e��k�#��^�L�Q
��y�^�]i�a�,g=�䙠�yRDL�q�$�ԡI:Y�d�G���y�N�N.�Yr��S�� kG���y�@��4���S;k6�iG��y�h�B5|��l�j�r�9 lK�Ř'��{�cH�F� ��eOءU�$�s$AF��y�׺B�~4�P��	N�!b$Eט�y�X,J�x +���D�4U���y��;q�4ݳ�$_AT:��AJ�<�y2�QY,�<�q��(CF� ��� �y���=V�aB���A�*����@)�y"�oa�U8 �P-F>ݸL��(OT�=�O��
E��G30L#'h[�R��b�'V��a��2bh��F�G�l���'E: �D�MvNb"�D.;=`���N��r��
��AU��]��M�ȓ42r���ԕ �|� �k@�����<�H���5B�9�"@B�$rsDT�p(�A�<1�eؚ*��A�JS&BhZ)+�B�Uܓ��=A%��6/�T��CJ�=�<�:���f�<��36�h	��X�V����`�<9e��p�<��DC�JТ��o�_�<�q���s���FOچG�*�ґ�\�<�e�*+���&��hQ����[}��)ҧe�uKv�ʩ;bV��HY�(�����dM��Y��`l���١ ���ȓ���L�;T�&T��!W$
6읆�	s��d�l9H��0�a��"�:a���� ���9r$��%��
f�8	"8��r�Ry`1NVu��Y�L+x�	��S�? �i;���A ��['Cҹb@��p�"Oֈ(�`��? n��#iA�X֤	�"O�����]��j'� jX�p��"O(eʀ��A<L}0s��[S��$"O4 8  �.�ބ�\"<Ѱ��y�G��m��/;ṋ�bƗ�y�-A�R�<�@�@\{d��A�y���8x����2�ո["%�ׂ"�y2*!&:XQ�C!��o����gl��y"h�Oю�H��.`����i��y�.�58����I��դ�y���=t���a��4�Zg��y�,|0(T�ǊuN^T�Cʧ�(Oh�=�Op�qa�Ӽx�Z�ɧLZ�8e޼@�yr�'R�I��i8Yb Ɔ"�����d(O,L0n;?��8s7��h��(��"O�8���G�d����P*Ԝ����	X���	�,TL\0p��ʥ=��2�
!�d��p���l�0v��D���K��!�D�?/a~�2�ײD�ˡ/n�!�$ÿb��4�)�}�d��Ts��'�R9
ۓ!i~��,G�@D�yZ�N׳z}�B�I�h��9T�	��PL����m��B�I��T
F��+C0	��ع,�"<����?��A)ĜL�Ɛ(�
�.;(ը�!D��:���*�=�C$�(1��d}�,6�%�S��MsD̀'.,����EGБ�c�u�<��"bp QiN�$��"H�m}��'�d����9w����2Ņ�W(����Mk�'Pz�`"D��9I��L���i�'�~I�,�b�$�A!N�B�PL��6�: �@d��}���t �%l�V]�p"O����e�tV��鵮�2���+W"O��`%G�l� SR��]�F���
O�6�&7{4d��+U�]Xbu�� i�!��#D���)RIB8Z��0a"�!_�џ@G���\OLh�3��4oo�{@���?�'��Ѳ@�	��C٬�� Y�$Z�O�� '��?��K� !U.�X�"O���ٚc���A&͆-EQc"OVPe��172͐cB��'O��R"O©(Ї]��j����H ����3�S��yB-�?_a<1S� 	{`h����9�y��̚����vI�-�,�%�R��yR-M�9d�L+P���w�`e� #��$/�S�OW��	E��8�t)T�V�O-@�'iL��?+�쩐��F�N�q��/�'H�J��2�#�,DH������[������۝I1�Ɇ��(DZ���Id���D��^��بFKR0�V�6m�'r�!�� ��XR5��p7�e#p���5x!�$�-0���!�
�23�`��si��G�� K/z�b�-M�Q�(���G�y��J��ԍ���0
��������O�~�Κ�SW��aH�$+,��v��R�<Q0�	)ny��� &|"Xrf�Q�<i�nӴ�4��V,�%xv�)*Ӧ[L�<���*G�D���H!za$A24��I�<���͟� !�I���m[�%�}?����ӦR��u�B D�19�,x��C�	�>�z�p�Jƍ��d�?�B�	��]�e�6O�R,bE�]�-LB�IR�ޭ9d�P\�r�(Z�$��C�Ʉ�܄�G�Q;�()�W�]��C�)� >�3��
5�,����T�
%��"Or�H��#��� �q�x��'|L�e����K�dX lZ���HX^��ȓ*�9�E!χ��Dj'���+2t�ȓ^DP�cga��x�"�C�7_0x��ȓM��R��N
�R�b@5%|����?�FjP�j�h���E_�Ipd,��oq�<��{C�$0���
Ou��(��q�<���
|:0RS'��P��T�Pp}b�)ҧ{K�L�4hݷ4`��H`��2�`��#�z�Xw��0����׍Xbb��ɔ����/�0=i!�f��� #�ɋ8�!�,B���<� �8�(�0�CF� �lm�,ZX�<����8�������;5ڒ)	r�L�hO?�I?UL~��r� �(搪���\B�� P�V�:u��+�ސ{�OѮ[z\B�	(~�da��SƠ(���t�B�I�G�D�Gk\iJ�F�� VnC�	�_j���@W���9��My�0C�	7AV��g�ӱ���jI&�:C�ɟ9�x}���
�h%ּ���<��C�	:Z���J�A7	���Ν��C�	�J�!�#k)`���aqI��x"8B�I�8�,��ˎ?��H�2H��fC�I�p�X�pa��9&�B�H��� [tJC�IS `�c�#2CJ"tɂn	�O,C�I=V��K�爺W����L81	 C��AbH}krI[�#�
\�D,W$j��B�0Жx�5�\�ZQ�Q nS�c��B�� #�ZP�i�Sd����� �B�	(V ��W)�,rt9�P,@�]�B��z�U�')�
X�˂�[�>�zB�	�}r�x��[�M��L@Q(P!DB��O H�`��1�D���8lfB�	�(�2��̞�L���
�S�T�jC�	�~gx�!1�,2��𺣢�)v��B��1N��Ia 
���w�9@�B�I�X-��3�ǹn|Ƙ"��1R��C�Ii��2u�	1T��dE�.��C� )%,���ûj:&@S�"��K��C�I�SXm���W�v��s�F�(s�C��!1�虫�D:a����jR�Ze�C�&{��I�c�$A�I0D�\�_^�B�IJ�`6#��5J��[�˙*C��B�	�<���ҧi����*2�K7TfrC�� 6��	�fT;Wa��C֬I5�0B�I�n�� $�>GXE����P�6C��'7Q���I�HG. rk�5R��B�	#7��(^�T|mR��J�|�>C��A�u�e�|�(<�g-�Z�pB�ɠ`}LV�I&A�"h�	"y�PB�	e�0���T�"\|�4#�w�B��-V8,;���2�Lxq�R<=��C䉣L�x`�cm*aT`�A��Q=/��B�ɟr��a��^��^�$i� 
�B�	3���#�7L=���u��*<�B���4؉#��Z��2iύz�B�^�~�[�B^*�4���,��X�C��p�2E�%�S$��Bd2�C�	.(YQgf1
�D�{E��-;��C�	�j��H��LL飓f�>B��C�	>l�0bƜ%L��S���C�	�/��e�Ήf<d b�<<�C�I�&O��UF	<1�"�!t��DC�)� �a1���z��җ!ٞR$��"O���VKC�#����ڭ#�d�S"ORԱ�ǒ/Lڭ�*Y��%"Op�)�u���V��8A8P�'"Oʬ0���.�L�D�&M3ؑS"O��������3�#���e"O8��'"��M�A��\"4�$�iC"O>5jD�
PB�|�3MS��R��"O\�b3k�7R�jTiW�xԐ�P��y���$M���ȓC����[��y�@�/pHY��-39���o��y�k�/J�8���'�Zq�����y�^Q��@��2�ԉ��	��y�g\.����D���3�\ʰM�y��3��c'��'ˊ���Ǐ �y��N��t@(��J���{%?�y��
#R8�1�����A���y2�̜]�> ���R-�i��K�y��7J�\�R�d�3�t�#�&�>�y��£"�*��"@͛:3(٘3B�y��_y�ۦ�ڸ2�fa���y��8u鸘���,qV�b�	G��y��<�h#�A�*#Tp��B��y�a�l��E
���lA^#�o��yJ�=0��	��\3M )q4�C�y�(š3vV��6H�/?]j�q���4�yr��9w>��r�:�$��B��y�"��n=H(���]6$P;�e��y�͏`Gf80c��0.��-��/��y��[o��rC��?!�������y"�E+��t�. ݆lAs(���y"b���%�� ,~0��N��ym�"�^-��Cˊv��"b*��y2���|�C��_�!e�웆�O��y�N
�sfh��B��7.��uJUi���yb�K�|?L��p�Y�9�-K�!Ȯ�y�k�-X>f �C36�)��ĵ�ybd^�Y0d��f�%(���0��P�y�B� b�a�8V�>5#2a�3�y��.���@5�A?����1�:�yB�\	x�lu�)��: �%C���y�e�QX�1�ʂ$-���@Ʉ��Py�-�� � !�2*G�B�ڸѧ(�x�<�IV�b+�y�	�F�,Q��ow�<���:b����r�ǥU ��r�a�o�<�$�	�c�x�&n��IPd��d�<Yu#̵ 4ވ� B�6�T JDb�<����&S�2�3��h�=��_�<i�6]b����"R��r�<9��N=��| !�7[[��	�s�<Q�Ć�C�zp��CO0X:��T"]n�<Y�j��9��X*w�V-<.~���/��<�VF�l8�v�E�eA���M��<i(��)iy34�L�F4��h
O{�<QE�ؐ;ӄl+��А[1tTx �l�<Y��C�bE�4�D7N�%HV�d�<!��K��3�f��N.x���c�!���`�*�B�&F�w��U���ݎ�!�d_c���W�ă'^ƴ����w�!���&��m���ˬF���Q�$ؕL/!��N!�l��"-O�W�|�d�i�!��D� �&qH�&��FF� ˃^�!�DٲJ� �s#ѕi)t!�ҏ�<u�!�ă�A���1�)	�����17�!�� nd�A�.}�\a	Ď�h��"O�����lS�UQ/Q�=8�"O�M��.R�|�|Iw/��)�l��b"O~08�cɇ��<�e�W�\��]�"O��e��>P�hؑ@Fʭ����S"O*��tM�Vi��� �f�P7"O�e�񩀦_�u���"7�%�"O��J�Q0֙�ɶr��aB�"O�u:S�K�d�p��Ae�&@"U"O���C=^�&�K��� ����"O��G��!�kQJ��5I
�q"O,�"vEE�{ \�	��-G.t�"O���kN�,����:Mq�A�"O�-2��1�ޑ��ğ<^疹��E(D�L��Ҍsr����5n�q!!%D��Ȃ�-s���$؊�BUz�&"D� ��$ݿ��h���,t���D>D���ի��N}��gȥy7�0�	;D�<��D3V�&����]V�|�� 6D�KQ ��:D"��d�E�^L�f�.D��;��34��:����Z��5H)D�l����p��ƆC�*FdQ�9D��[5��+7��"�K�;����"8D����cK6.I%膊]56P	)�i2D��"�S"p�
\cpŎZ�r82`*&D�����S�f�Wm;��x�H%D� X%J�'"��֮G|��XSG*7D�X�S� :$d���@�!�\�#�6D�ԉ� d,X�{0���e�����.D��"%m9f�$��bb�l��#e-D�,�wl��EJ�!�.�RdـE+D�|�G�u�D(R�nAct �E*D�$�ņ�>.��@��YON����%D�(�f�P�n�<���YX����k$D��ag&�~���-�?\=�����/D��B4 �<}��2"�4Ҡ��a(D���B�V �ą��^(A�p�&D��m:o��ٸU�'�*�a�)/D��rt���Q��l�Ѯ[4AS�/D�D��ޜ"b��C�^<�J5-D���'M�s�"5rGe�2WƜ�f�,D��i"jߌ-�B�_2?�t��(D�@����H=���u��ؐj:D����9u&Ԩ2�P�p�&�7D��R ��i^|-2mE�Bwh�9�4D������ �:�K�jɃ_2y W/>D�Hb�͞�.�Ha��nƓ2t���/=D���e����LTB�&���$��&8D��3��G�>����Nb�J�kg*O0$XU�Q�+N����ѕ#�Z=��"Oԥ��D{ۈY᢯V�R���)�"O��y�^�Xf�T�_8�\�r"O5�lK�=�^(�����U��"O�سg�?��uSp$M=�`�11"O�2I�4\��"�Bǿ9�`2q"O�|s��7=hTl��J65jT{�"O�ѣ��|ߎ0���0"O8�TJ.:���
�/@E $"�"O��$#
�g���2P,��2�Qs "O�@Ȧ]/lh��[#t�|�"O��Y�@ W� ���ʘ
�mbd"O�v��GL8%YS
Y2OV��9�"O> �&�U���P)�9p�P�"O�a��G�5�~�HdgIGZ�r�"O� �92�ވpB���]K�Q�"O`-�-�(P� �&�P�Y<8��"On�rp�R�^��p##6j��"O���֨H ǈ��ǅ�[!�Tʴ"O薶TB
LX��� @� �y�� <@���!L8�rѧ�	�y��Q�]��`��	=Q,5�1�+�y�U�*yl�"�	�#HI�J��y2j�\UԥH�i] $�r�0`nY*�y�h��ZHN�`  ��l"՛"E��yr/�)�J�r���UH�q!e�/�y�C�%��]�u�1H�aҳ�Ϻ�yn�0g�m(6�֐&Y�yZ�y�Q4i�@�+']!
��dC��y�>?eܡ���H�c@��n�2�y��V�(r"�a���	z����ǘ��y��'B� ��/d�aB*��yB�I2Dn �ҪT��@B��%�yB��*DjP�u&���0pQ�Z$�yBLI>t��]��c�}1��b����ybbMhzb=AC�P�ua�܂����y���i$	�F U�w)BX9c���y2�B
h?2�
� :n���-
��y2�4#0(򇍄p��-i��T��yB�,@��q�nG�����(��y"I] =�lzQ��H~h� �m���y"gOT���;$Dښl'�m�!X��y��Vh���Wϫ\�h9P�횴�yo�'�x��7H��VNf���%D��y��*[X�ab_�U��q�ȇ��y�Ŋ�w+ � bWOzl���!���yR�B��B���-��P�a��F�y�$�/��R	!W���AA�yˀ
T*J��O�{8�qRJݚ�y���_K���@"}�ѧ��y�a�s���I�N�?�K�439�!��X4R`��U�y�2���e�7}��I�ȓF�L��3.�V%SÄͫZ������E�B�s��	[�g����j��ɀw�2 %�$e\�H!����"O2đr�ʟ2d~��Wě~��w"OB��$�9\��!	cc�]�}�"O�<BfݱM�� "�`B&��� �"O���$$�|��/]�'�Z%��"O�H���̤�F� d�^�R���"O�(�Ro@)JX2�!���l�Ҡ@"O"mc�%�C�0P�qN��a���"O`�@+�)�ƠеW��<�a"O4��`�M�Ƽ���{�!"O6-��F\�\�
6�P�]4m��"O��%Ÿ����h�Z�,ɂ"O"���
��D���Lިx�Tt��"O�2�bT�+MB,�SKX�h�,�P�"O8�j�F� ~
<���zy�;�"O����J�Y�@R��S�p��"OMٲ��s.������< �"O�qᶫ� wX��C/w��`"O�qc'��U�>yg��t�"�x�"O�u`f�7'X���C�w�|�V"O�c�� %�H뗬�Yd|*�"O~)C�퉢5G��c��?_^j�"O�9h��j)�x�j%"_&eC&"O�XT�S�#y�h��(R wN�`!"O��s�j��ʡh�wO>s�"O� �6 ɱ,y:��H߶J�ݣ�"O]P ͎=7 �A�5e�}���`�"O�}�T�^�3��kdNVl�̩�"O�e	�-�0R��G��
���J�"O��T�ߏfMz��᧛'MĘ�"Ot��B��0C�t��'�>a@��f"O����lR�_ �z�%R 9�Pw"O���@S�&����kL�t#�(H�"O�lHs�뾁�`��0B��xU"O0d�aɏ{$���6�g��y3"O�!��'���2�_M
�BT"Oih�\K4"Z���,��"O�Y��L��!��,P�b�N����"O���ӧz�L݀qk���"2"On9hSCJw�|��J�>���"O�E(ׅL�5T��{��.V���d"O~u�f��&��� ��/4���"O��A�Ĕ#�BM@�GQ����2"O���S�
. 3�|ф�?�@% q"O�勑��p�B�E2����@"O䥣Q#G:|H�1z�@�)b��P"O<U8�bn�!�1�ǌ��eI"On��Ȗ�:1�4��ߎ,�|l�$"O��Ұ�I�8���@��h{dDi"On���%0��p��ToJ�[�"O�
%͝�iFd����]�����q"Oh��uO
'0�tl�Qi!�dњ�"O�}�®_�&�Pa�V��:ؘ�J"O"��m�	�����6LqZ�0�"O���B�z�j��g-T�}�`C"O�XJF�˷�|Ä�b�� 6"Od��L6O�}����dI4@��"O��PGW�F�t ��J�	LMJ��"O����E�Zq,�p�$�g?��J�"O�1+ƿ/�H�R���0�l�e"O�� ��<J����^9����"O��R!�S�
���S�y�\�Q�"OംPGD2�1�&L�YcV$�w"O�<�ce�iV�q0u*L�^�0�"O��SwmJ>�8#�M(,�TГ�"O�P�"OҞ%(m��¬��v"OHA��B���B�xЯT���"O`�tm@;��	k�(I�x&<ca"Oꉃ7�A�8�z��Ǉ+<�Q�a"O��Q���A�*``F�)+X0��"O��:T�C$JrRE�R��;]%��d"O��Q� ��C�Hr��	XLd"O�d�r���X�^��5!���T"O�ct��B�x��n��3�v�#�"O�|�Ф�|���Nd� �#S"Ot<V(�8�
5��됉E��k�"O��H �Q�|�BI�2�'*��u��"O(�ȶ�V�>���륇ӘV 6��v"OV|�f+>��	A�Y���"O��!�c�v�.ya�ƻ���g"O�X��D0����T
�y�e"O�a���� g��E{Уc(���"OvZ��$0%������"O�:��ڰ���Ku׭2��"T"OdA�s!זhr|��CHw爸�T"O�!@B'T��=a�95�pU؄"O�a���٣?5XX��D�"O�l�gg�:'9�����Pc 9�"O�¦Lđ17������fn(���"O� ��*DM��,�k�cFve�4��"O�a�e"�,T���
ЂH4$u���v"O�h��$)�aًj0@'"O�y�ΙM�2��iO/W���"Ozp�r��	9ؠAi������"O��9֣	�j�Ib��L���C�"Oz��p��.WI[�)��QD"Ol=�d�L�A&	���A>A "O��B'�/"���צƦv���V"O4���^g�"����1s�@J1"O�Y1�aK>66�m��&��P���#"OD��tKV$+�.��e&�%�ZCr"O~��c�������H2g���V"O�l�S��3[Q�(�c�m���#"O�)!6k�;V�:�S#"����"Oxx�e ���$�q@����Cw"O:�(���KH�d:�I[+E��`��"Oؘ	fDZ�VN�{�(Z�m�*	��"O��PT�![��K᭖ %�{"Oډ�� �.[�|<P#m�0�$��&"OZ(��X���%�"�_2�E[�"O�`��O�Y�$�k���l�Y
�"ODa� �I��y�8i�n#"Om�'&TP��Iy��_"a�<h[r"O�h��
��5b�i �����ᛴ"Oj 
$#d� ����b�hԋ�"O�<�5&ɴ\ք��udK2!�]�0"O$m����Tiz����<Y��"O�!J� ۞PH�(DMCm��Ӑ"O���k�? ���lH�!/�$��"O��A�D_�?\H�Q2MA8)&���"O�lP6&\�]nZm�?=��i�"O|�;��S� HD%��
!�6�R�"O�0pq��CfdY:�n�h�%��Q]!�UbФ�2��o�,옣�S>!�h�ZQ�K�D������ͭ~L!���>�,AZ�%�~�T�S�D!�M	\H᢮L�Lzt$[��@�9U!�V�BL���C���`�x��ȇ�8!�ݸVcd=�g�# �"E�dʎ�1H!�$�'��X���:�b)�vC&4!��"GR�h�h�8fl-��B�H!�$�uB0���X�XS�T�aO>8,!�R� a�7+>:2��2M�~q!�d�;"xJ�G��5.I d)>!� HN�S'I�#s�:���<P !��Ě@��yhR�K��1R�jƥ.!��-w^D�2�l�7W��H���̑x�!����e���!E��? x���Q��	f�!�D�Nl�� ِ2w�zdb���!�$®"�M+��x-�6���!��M1��HPw��-%��t	��O) �!���:k�@"dO� C�$��.]�Q^!�H�l�p��$�6Ң�!�.��<!�$�={m���Jսh��)�F�2c3!�C�Eb�#�NM��|�v@C!�I��A3�M*@�<W`S80�!�dO�S�#L�)&خ�;���h�!��+:I\�����+�j�����!��ݕ}�`fE��:UX��ȉ.�!��,k�F\���tK���!d��s!�Y
B@�9�%	�2�	+3"�$:!�D�:Z��j$IT("���![�U!��P��t���I��MA���!�� � �K� ���%-1h����"O�HǊ��Ș1wk�P�u�b"O�P�@�
��Y:S �� �v(�"O`KW䏷-�LъV.�6u�1�"O��@��1'~�Y㌟.����W"O�I�&���}��}[�$\���U"Oր���؉5�� C�iC�O�J<j�"O���^�@-(M��-ֆ*�>�!�"O�8㒭�8p*�'ĳ;���r"O�p6O�/M� �%EQ"J����"Od}JG-�)@tʤi��@���q1�"O��P��
���hf�@%�BP@"O8��c)�^X*3CՀB��`i�"O�������N��G �?M��:E"O�i1%�P�O@J�@fn�x�VM�"Oʁ0r��^<��coE3��Dˁ"O2�Ps�����#"/�
 ��&"O>Ȋ7�!g\ �.ϫq	�У"OIi� ��66	�LM�4�\85"O���A��^(��b�R.#<k�"O�}fg�W#��)�j�}
Yp�"O&�r��/��	4)�;87�9T"O����査w6��Pˮ �6,��"O0�L ylD���]�H ~��u"O�U����&F8��i�2J���"On�Z�(@�)����a�3+	��"O640b`Y�w�h�u��2�"On��a�ΔZ&�a��� �{l��qD"O4��c��)e��eu$ª|��"Ob 2����YG��0#�ɘ�"O��P�ѱ	�1��"X˴�j6"O��n�vJ��1�*!,}��"O������)+E�՗D��́2"O�32�/"��u�s�Z�B�Li��"O�� �ER�0d���h���!ҧ"O�L��b������͏@r�mp�"O�|�#�L�%�\�:$hV��P��"O<h1U�O��@;���S�"M�""O�K� ��_a��P�p�8s"O����+�����.���Ss"OvI�Ԋ��#��UڤKVd��00"O-� ŗ�nn����*I6м��#"O�p8�^�3B���+�<��`5"O�M���ɩ^�N"��	-M�aS�"O����\Z�*p����*H���"O����8�L�5��%��a�"OB�嬛�!ˬ[�A�T�^"Of��LF��#+F�%��e�f�'D�����E�ց'c�=#��$D�Hjbဗ:����e-�a$D��)�߀�Da��x�Rm5,"D�d��s��`R�\+!H6y{j:D��9�JV�%�tԣ�)ܟj����A�6D��P�$H�f4'�Gr�Q�b3D��8U��Vn�u��*�.��(3!�<D�l@Eg��=������"����<D�HC��en$"��խs@��7�/D�4FAV�D����Y�4�����L/D����f�=9���Δ��f�� K-D�v왅�j����=��2�+D�d�"�<� B�\�L�ʠ�*D��8�� ��UY�aƬC��j�-D�0��˛M
�3���E��X�!>D��q� ]��y��#<�v�[�e>D�� 8a*&c	'K�j=󑉍�2;��3"O�8�wL� 9��µ���$S��"O�a��T�!L��C�$(J���"O�,;4�ۃL|��9&��)�޵�"O����jmk�\+"ެB���S"O�4��+�P�j4CFT. 	
�"O�T+V� 5�b���ծ)�1�4"OLqP^�qj#�P�$ *�"Ot!�!H�gS� i�K��{�b���"O^�㠪�W�8���)�S�V�{�"Oȉ��+�)_�$�3��1�y�B"O� ��,��W�Pi�!)��2"O����)j���� �JY0�"O�M:�؍).���V�6�T��"O@��HT�5����k��X��a�"OJI�Ǌ|�����]�J"�H�7"O䨓�M�6`��9�5c�N|F���"O���͛z��q�w�˻	uHPB�"O>���7R���/�?FnY`b"O �ہ��B)R�[�.�^(���"O��S��J��Lx���j���"O�ar�O�:���P���XR�(�B"O��#��Y��`�ƚ@-PP�"O�|0u�<@����ͨ^�B"O�ԋW��:�P�5m��2^�}��"On5{��n�
���˒	'T�<r"O��IB�I�=�B\�ThI�D��A"Ox��s��"|�<�bP���2)Z��"O�5�g&�� �&�9g�XXl�"O��`��ë:1�h8�ǐ���) �"O���sh4u[:��Ag�6(��"O�	����
^�a���@�#��V"O�8ab���AvAa���"O��Au�Av���u/��T}�P	�"Or|����13,��؁0yz�0�"O����`�� ��S��Q"Cq6U��"O4�8��c�@hP�I2#nj<�4"O\�p-={z�dY7�	C`���"Oz�����Px()�2D��"��t"O0i� A����C�^4bE!��(D�dxc.B��(iv&&)���4�*D���ƫ�\TL���6@=���d�)D���3H�|M�����21���fa(D�8��N��B(%d�.$h�J�#D���*���)qD��V=(��uh=D�P������4���V�,$�d�5D�|R�B�[���"���`���l)D����͌�U����j�w�L��bK+D�T�Ɣ�b@b�QC�W�m� K��(D�x�V���c�x U�Q����S��1D��b�EG`�@@ˢo,4$�@���3D��!���3C��(�
I.��!�5D�D:w��W�0HɘU*R!��3D�X�Di�8m消���3<��U�4D������*+W
���GH��p�v� D�P@f/�
��PF�9=�����0D��B( `(�8ސD�6����_v�<	TD١v��j!��HTX*r"�t�<�Z����� �@�@�\��'%Jq�<�Rf��ȭ`�!�&(�2A�%Ih�<񡀈�����J�d� ��u��a�<�`V)�Ɖi��J�>.����f[d�<����72p\�8@V�V�En�V�<1"�>p������u�]Z��� ��/1Y�#��w4��+5"O,�cv�]߈D����!%��2#"O2���*T=iVeb% �
��J�'5��@�%ntY�'W-Y�ڵ��'�dA��l�#U2��j �X=?�*�@�'�~�á�~���'B��!AH]��'g�=��N�a�`(�g8&_��Q�'��|B4��,�*��++H�$�`�'%ڴ1mЋ�(��1��K����'�x��ԫ�Q���:���(?{���'���
�"S���U$�, ���s
�'�.�ZC��eͼ؃E��#e�(��	�'�f(
!/EZN�9��^��q!	�'l��Yo�pv���!�4+C4�	�'�P;�aѲ@��`�Q�H�%;R��'�]�� ��c��� i�6o����'CX�H�99�(���f�h��'(�!5�3DT���#]�}h�
�',8ͱ�
+9���
P#}$Q�'y*Q(��H�����a�xA:�K�'�t�8����N2���+�>]��	�'WL YD�Z�nH	k0�[%�C�'f���g�T*1�E�[��y�K�1g�zĠG�I�N�*�*%e���y�C��5�ne@VJ��I��q�D�_��yR�M�Yۤ�i� �At�Q��y�iZ�	W�,q@.���@��R�yO�%/`p!���;���ks�	�y��֡"IҊ�;:�^pc���y�E�gV=0��01���� �y�ZJ=r�-ŝ{_�� 6,�yk��C�>�����s���FO�y�M�J)���Y~%K$�ړP�r0�ȓ�I5�>�v �H��X��ȓq��A`�'��oMN���	Պ�p�ȓ-�|Zb�[1kђ��w,	>u�ް�ȓQS�$j�o�3R�$b%	#�h5�ȓF�nQ��璷0$��ԏ �z4�ȓTf�8@L��Fx����?�8e��?�	�	WD���Д��e���ȓ56�ۧL�8�D��!�]锱�ȓ4LP�՘d^X`I��>E�ȓ=O���r�?`�4���P�r�x���M�d�U���E����[�������K4�ܪ�|��mOn�x��p��c�N�sB�]��O]
d�ʱ�ȓ������C���Lz��uv�4�ȓ#r=Q��	�*d2:��έ[��8��HŦh�JV�P)�V���l����d� d�<v�Iytb
K*�݆�]1,P�Eƒ]�������Q�I�ȓ'$��3 ��4�Ց��K2*ڊɅȓi�]�T-Z�ݐ��CG� �Ҭ��_A<��Ѭ�޵�a�S?����ȓ�*Ieɛ�D�4��A�(q��2/<��6͜�+�.q,�P/I�<$�-\���#Z9�)��AG�<����-Ŋ\�dÝ�:�Rus���B�<�楆�hC2���*��	���t�<���$|,��A��).�Z�Ko�<��ƮF|��ɳʃ�}��}ʓDh�<A��8Dx��o�*l� �`�<��FQ���.�Y^��ɥ�,.�(C�FA�3�,�!$�r)�ժӴ
Z2B�)� Ҹ�����UЉZwh���Jy��"O�e� ��6W��X�'�(@;�"O0@�ɔ�U͎�"�^���+�"O*(r6��"6��0[ƍ�	V���Y�"O�ݻ �2J!����
�2r��"O�$%�)�\��Z-9#�E�"OB-�q�Ȝ=�Ё��/G��1�"O^x��c�3
t��K�*�D�%"O� ;Ū�6w� 0�M1n�B�g"Ox��q�W�o�������["Oj��0�N�X��4�u�ɋ�иK�"O��è\�H���R�@�5n�y�t"Ozh�5郷~��BǪ�fxQ��"OP�H��ͭdn�x�D��;� 9��"O$�K��_�u�Cʆu��|��"O�Xg���g��q���Z��Y�"O��qc�<z��a��E
�6�BI�"O� ��@1b�܈D3{�%yg"O�q�D�U���*��T=zq�ap"O��ᗠ��<yt���tQJ�#r"OĐF�;p8z�sGa�f�"��2"O�7���"Fze�%H�q�\�Z��.D����Ί>_�3���=�*�2�/D�P��0�����Ų_��C�*D����l�+2� �*a`īp�8:2�(D���Wf�(m>$�PDဧm�	8��!D�H9� �@<����!6���1�!D�����3�`�	�A�))q� D��Yg�#"��B�3~Є� �;D�@��!��U��j��M���q :D�����(N��M��	�� �N��-$D������E�4͡Vk^W�� ɠ
/D�D���R�$�����(g������,D�ȳ5֒M뺌*�!N�B��"�+D�(b�	��0T�w����#��(D��2!Y�S���q��r果� .1D�ȩU���"� �r �<o���C!0D�D�d�7@�H�I1U�⦫,D�4��/7O"�4@��)nfB�ɵ�I{�� H\�ab
4:VB�I3�\;R生/M�%�����O�<B�	#��i�$�^���;�OL�dB�I�^R ۳�	,��(C�
�@�C�ɏz�����L\fސq�M����B�	�Df�;����d���Q�C?B/�C�;gv��`�7$���ڥ�V�B��$F��(q"���zg�)#PNA*�fB�I�q@5�� ��8��:���p�6B��)\�����ȩ'Ψ2ee�]RB�I� d� wǉ�A��܈rcۗ}�C�	�i�*�R�@��v�;f샱�zC�	����)��/��1�׼2dC�j�ī��
)���z�ǟ=y3�C�	@`��/[��V�����o��C�I(*`�u�S�N�6���+W�*|C��0D�.���-B�c�d�X ���t=4C�	���$LS�s8�K󭝉*m2C��.uݰ5�S�S��1sfێ	��B�I�<��M�oR?p��(�(�5@�B�I�
��Ke(̌M����n�#Cu�B�	!G�<�9�'��+����n��B�	��Q�єGn�U�" �%)Mh`�
�'��p��<_J�R�
�%��,�	�'i̘2�^&_��+�+ϯ+�dX���� ��1C����LT9Z� @�!��"O��F�P;��A��G���u�r"Oԥ�OQ�$�S5-݈�zDCg"OZ�s@		l�,�u�}Q���"O�DN�2m�m��̂��<���"O II'g�<d�$薅iž*�"O��f�*�����Q��=��"O��K$��#�L���P8���Q"O�i"�� M���Z2�\E"Ov8� Ĕ�o6�pP�-K�ށ�"Of��� \��:sǓ.w��S�"O,t(��^�2q~�����H�#�"Om�2㏐)��9�G��M��"O�0�"�_e���	����p�"OhXЂ��(=��h`.���pIu"OZ�cէC�v�n��$��"OB)HF��U�倱�^ 1\Mr"O��3�M�\f�(�D��&+�Q�"OB��BϘ�hl	#J�=]���#"O|�k oQd��h���*T�
�3"Oj�$-�,\��43���;>��\X�"O��
���HԞ�)�A8 ��*�'�b��S����= ��`�*%�	�'d�\{�#yH "�E�]�h1i	�'>y��޲G&2b�ۻN�����'��9�`��d�ۛ6�l@�'�(�k̙`x����E+()P���'��YW�OZ��r���%?�H
�'���"n[7o,��u��71�0�	�'��a��0�\�
 �,Z��`��'fp�HQ� i�ΐ1����^��@Z�'g�hSE�\�~<����\�j��IP�'y�y-��}� ȩ`MeL����'����񣊺v�2��FV;/Z�+�'æ����^���OT,��@�'b�e��f�7ݮh�ձ!&��'�y��+��� H��&pZ�'��[�n�v�9�Ӫծ}����'�U��cр2�
hQ��ӭ}HT��'�rxbDnЗy}n�r`�p�'l�,�&�$���#�e�d�p8s	�'��+d�W#5�% �F�.b.��'8�Xc���38��r �)��-��'��APb�c]z��re�p����'������
���u;�(B�g/����'y��If�� ��i�&��i|(���'�6����g��f�[�i�n�
�'@|I`3ÛD�r�#V�^�aЂ��'V:6�� �^���O��bx�'��-*�j�D�zq9��Z Ph�H�'D���6��'"<��j�6t���
�'��=EN�p'&X�!aV;n��)
�'Ƹ��	�E����N�ߨ��	�'GDI�a��F�5@�h�.=0�i�'@�ͫ�b���Eڤ+^�:P��'
\Is3 įm�� R�Ʋ5����'�z�"c��@c�t�c���ʑ��'���Ⱪ�/V�yp�)Y0dۈi��'����(�,'X8�s$*M��)C�'��`�qi6T��pC��#3��Y��'�%S1�ɻx�F�볤Ѵ2a|l�'V�\#S�s�H���+(ΝZ�'(���HD9\��"��ν"M\Ih�'���	ә������C�FY���� �22�?|�
����=J����E"O,��c�8`D�U+P%uX�x�"OFŹC��$O�X0���(*:�4�"Obs�˖�.��1���6Q�����"O��C��S >�h9�d���Y�L`h�"O�!��?���o'I�:8�"O�$ڧ��9*�v����=�~s�"O�A�F�F�u{�F,+,0��"O�yq.G͸ �cm�y��!�"O����%E3q�|�k�,�\�bQ��"O������1a��9u���L�,s%"Oa#��.��	��[~���v"O�da��,۬�Z7c���ɱ�"O�ݰ�l]h���B��")�`��"Ol�j�@�oZ���F�c*B�A�"O�$��O$�B�'G�)�l�"O��"`�O�
1� ��9F�K 	�yB���'��(ŏ�6"ٲU�[���8�}�Q�.զI�GbR��)��$k(ih`��2|���A�W�j���ȓs���`��*X�AH�[�M��(�ȓ\�����EN�;8���ǨE��M�ȓL{����@�{ds�%4d��ȓp���S�h�#�j��UoՅIDH��I�<�i�lƕj�*�b	zЄ�6ԁt�Ȥn�X(ri�G�,���%s:"*� k��)�FX���܄ȓS_T���J��f�����-O ���ȓ ߀��"j�i8U�2 ��_!�u�ȓ`�̼� k��J���`��G>#Ő��ȓ6jP�Q��P���	�7�G�uc����"Y��0t��8W�Y� o�D�ȓC�>{�_�gܼ+#+�*A�p�ȓVAjɻ���K@��	F��ȓӞ�i3KN� ��]k��&1����^��X��L3L50��#�z�ȓ1�\�I���)P��t�rJ@P���ȓ~v����4*�M�Iԑ-���	�I�E�"�J�̅�zՄ�UT��$��8]�~d"�	Q^.��ȓ� ���c=��q�f�ЅȓR�����#�4a޼t�W��!�8�ȓ
B�r�/�5���ƪ�[:��ȓp=nŪ&Ά�sm���,"8 q��X@���W?�,�8$h��W4j���7��(�&�D0q��dΤ.ކ�ȓIG��j����"�Rl�v�Eh�8��k�l0H�D\�O=6PxĬJ!���������k	[v�;��K6-�̄�[�~й�h����M; �V�,_꜄�"M0��d� 
�jt�)/��\�ȓf���gb�:�Bpbԇ�$g�`��ȓv�P��Ca$\���0L��C�Ix�Xa��ğ*c0�:'K5;ԴB�	�[J,`�e�9\���C(H�};�C䉱��]��S:y�#b�0%�C�I�92�-b�)I6�Д��l	d��B䉃p��X�/�"�^�p�NM�5UvB��(e��}��F�'Dq�VA�<Pt:B���Vd�EN  �6qؤ��]?PB�
�*1y`%R+ ��$�f̏�d�C�	s���U�3���pr㍝9�C�D�}�+�#�|l�שM	?�C䉃OiB���ɞ	@���Ӯ��xDC�)� �p�EMR �t`�(S\~�9 "Ox�[%�#_,���� 
,H�S�"O�2�)bl�E+y5�yb"OM3�M �h�hl���k3"O6a�R�ȶ��ɑ�w�d��"O��J�͍I(l�d�����"O��аᄖq )K�n͓�Z�a!"O,ɢUlY;r��Dѣ��!#��b"O¬�w�Ŭ$�Z�Z���=:B�C "O~pB*�M��<��l֓�
�0�"O�It�S�e�`���Z�Q�B��g"OJ|K#,B�'Y�}3�j���"Oұ�c�L٠p�����B%"O��P�ǡWe�qXg�	���)d"OX�g�^4(fDSE�#��t�%"O~�"�CQ[��]k��;S4s"O �뤮���Y� O��}��)"O�S��,hJf	5-�u����T"OD[Rj�9��̓An�B�p�"On�ґ�߯>������!N�J��"ONiQ�`�78�e���L�F.$�C�"Ox#ֈ�&T�B(H�G���,�[�"Ojc�U�C��9h�ǈ �rax�"O�0���,y�{c�D�qnd�"OցQ�b�,3�8�;g̝%��mK7"OZM1S�܈0njBAW�{���Cs"O�ĩT��\��w@�z��Yk"O��S�=[PyYv�%O����"O�����:s}|p+�+����"O�%!�cW�[^��%�S6#ޝ�s"Ol�z/Z�t�h1�PgW8v���#f"O��W�ZJ�
4�U�@�&B܄�#"Olm��/'����)F��"OL�(��);1i3*�5b�!��"O�\ ���F-X WaM�E��y�M͇48��kT,1:�|�ph�y2�B;c��j%���=�J=�#��y�h���L{�k�h��Q��y����Y��C%}�&} �N�#�yB�gZ� �g�Q,zg8t����y�_7\�WΏ�r{��@���y�� �/�� �7d! ��2��Ź�y��ϫ�aJ�N���| J���y�(�?���P���z|�5���y�W�5�����.�b�	�y��@7N�W���H����y��ҏ"C��Kc��5!��B��(�y����_��T#��};¥�.��y��P�^�����A*-�����=�y�I�A�b�z$AU ���4���y2�"kXap3J�B"�ɚ!	���y��t@��PP8>?h�;q���y���(Ш�0(��;PF	;A���y���&+�����&B� M��yb�έu� �dZ�o�,�H` ��y�f%�8�k�qր���"���yr�_�YC��a6��i�~hw`R�y��2�v�R�P W`Z�#�!���yB��udB�/I�~h�Swc���y��A4�!�H� �v9P$I��y�K�.hD��V	�h����O!�y"���c6���\�X��!�y�J��bӀ���և9��JcLG��y�,� ������0ؚ��F
�y
� �<C.	�%8"3&D��lS��#"O�}��D���뱨.?�!sP"O<|���O?~�lH:���<�Q{`"O�%Qѯ�	���Zs���z2��)0"O2p��	W~�V�G�D�gu �"OP�B`��"r�nm�)��І&D��!G"��o�>�#��$T�K��y2�Zy���	ƚ^>xb�.��y��_�ⰀǂU�<���0�y�H��H0�D�B�xH����y�FX�P�U�D��]ZG%T$�y!�"1�
���8@۾8�V�3�y2Jݻ%(�`�'�8>��%�Q$��yr�37WbI��n�1����'�ӈ�yB���I����m�� ����eE���y����B#H �����o��y��C�S|��M�1D	�IY��y��K�WN\:c�ߧ7�b	�S
ƍ�y��$��� ̪{a�2�"̥�y�U�	��[a(]�(,h��	��yRO7{W���w�����0�"ˋ�yb���;{�8B ��$\鶽A�Mƛ�y2��&G!|��%J�8k�R�'�y�1)$8h�nQ+vְ���ۇ�y2�&~0��(M�v�*�A��!�y��H�x�%��g�*��A.�1�y2.1#~��&��1`�(�3Q��yB�Q�~{Td�c蝇XClXAlR�y�J"l����!�X�?����Ө�6�y"悟����ޫ4�<�S4�ѣ�y��,\�r��?Zv�[s��:�y�ȏ&�x����,��5i�F���yB�˲R�"�y�-�d݁�匆�yHO7nvX�I���(��$!�y⧞�0�@���D|�f�������y�mΒ	Nhe�(	�+丕j��ȓ�yR��8
���Хl���$̐�y���#M>V�ku'�f�D8{ԁ4�yr���G��ݓeě� ٶ���yRB�;�x���I1M�yya��yr*K$��=@ׅ�p�Vܳ���y����7�%p�Ag��`�e��yb�À3ޔʒ�˂�T��b�ѝ�y�i�X��8��A���`rg��yΎ�5�ej�/R�t��laQ	J��yb�G5��a�m�p�(	f�ȳ�y�AŻv^$x��)_����u����y��L�l�8����3ἩQ�!��yR�G�ԬA8�튝2�a!�A��yR����qk�� &��q���y��D�<.)�'��k�ʉq2B��y���2Vjb�s�`��g^ĕ��/�y�ělz 	����H�&!ӡ�߄�yn�@ d���)@:�x�qH�2�yb� ;/p����B3x�8q�ծ�y��ސ@V�H��%A�Zճ��J��y�c�4jf%Y1�,=%��kB�	�y"�=���"�E�;��!�&NR�<#	]�$yPC�6�B�n�<��`Hfr|J �P�+Q(4�Ӌ@k����;VH�#"��|�z�`�j0a��m�ȓ*rI�@AoβX B+QrB�ɉQ�Di���� ��Ċ� 1ZC��/%c��h�+�fq�q�O��F�\B�)� ���*@�$�����.SA6(�"O�H��E�&KZ����o7F�)�"O��H���7nP�!Ԣ�?����"Oʕap�O��9����^`�)I�"O�9H ��~
xK����nj��2"OB�"��@�r�(��(Of�P�2"O���$�7�� �>XҵCT"O�L@� ��:p@�AA�; ?����"O�"!˕%]�"qE�8�@��"O�p�3 (vZ� z��X�[Μ#A"O�0a��B�yd�=�e"c�:,s"Od���!X�Q,VV�2�)b�¶�x"�'����f҆%_�Z�aL��2���'%�9`T#�7&�X�C��f���'g�ꄢ�(-�8��Ò
����	�'�)8c���Y;w�փ�����7��T��"nɷE��};��_����ȓ*<���� j�.�P��]x(���vxT��͓�
�R5��W�ҭ�<Y����)��UތG�rGe�?Q�!��M�2n���7��p���Cc�7!|!���i�*x��F|���E�x��ȓ �����DA�	}���[��d��`񶼫�J^��@ +��۶\Q��ȓI`FiJG�E< �ڠ2�)��XW"�ȓ 8I1�Z�uO��R�8I{��Gx��"�S�d �������O�hV	ߜ�y"@�aq&0���I�� ��e4k�Ez���'4T�[�%!���S@�!��	�'F����g�RPp6�׌��P��'�g���>�"2�_��|(*�'7Nlٷ�Նs���o���ԕ��'s�Q'RC̰���&A�PIj��'��1��r�6�qF�8E�x��'���#D��N��p1�c�?=�a�	��ēM5���,@�blfL ᆘT��4�ȓ�r��G%1X8�ks���Nx1��Ii�'�� 5nپ$�6���%� �ԡ	���'�r1��hK>@��[���exR	�'}@�[qƎ
R�@��7�ܥg�.�a���?�S�DNW�
D<pj�#�!5y��c«�y��BaB��$�Q�F��	�0gL��M���s���3l��i��x�%X�s�Tٰ"O��;R��Du1�'�3԰u��^���	�o1I��i�ey�;sb�2޴�����d�<���Ĵ@�B??���Bh��*�O���NT�\0)7�Q(W�N�J��dq���O(���X=a���� �3A,�$��O�����'��ayd�������	�?�����X��~�A��P>�E�x����6��y"E�	��PK����m�^\q/��y(�9��\�u+��f31�̽�y���
Ƅh�sO��b���Cь�y���1Z�e�g��V�܈��"��y�F��nh&=
���d5�8�J�,�HO�����#J���B�s�B�$�J ���G{���'߄x$��P�:�Z�e;����'�T$���ԩ�A�+_�lƥ)�"O�<�)ݲ:[&M��JPZ����"Oh����W��@�BJ�!L��Q�"O$�(w֠18�릢ƧKE(�0�"Ohe� ->���H�\l�"O*yC��ɜ'�R�P0$��,�� B�"O��9���L��4kE���i`\��"O� |�qs#����Xd�O�u���"OΔ C�]\-�u���(�^��1"O�@��$e��6fH�e�2"O�E���\�^��˩;Rh	�"Of���E-��=C�%ǂ68ve�"O�@{�G�LI���~ņ�0g6D�x(w	�.�4a7b�2:�X��f�4D� 	��bY���i�)$`��k1D���K\�7��)���Ĥ*Pd��	/D�`���-i4����ؘf���Є�7D�0�# @i QI��3n��H�4�hO�,GX�-�?7O��s�aK� ~�C䉷2�~؛�k�e���$d	�ƅ2D��@̏
k��9�F]>S&,[2� D�H{V'�.����U��&;Đ*��?D�\y��A2]�+7�ЙL���&h3D�,�PJ;B9
���o�"}�	0�0D�軃���=Ǿ<!s���C���;�:D�����q��5�2��(���j�+#D�D�JG;�yQAǜ��T�E@!�	��Q��O�>��%��8i�H�R�ʲ	A*��/O
���,G��5f^,:&�D���,�"�=E��'�Z}�RIM�a�����(K�jT��'� xZ ��'W%4�ҷo�8���K�'��b��E֘Jc)?%@��M�yR�t�A'�Ɵ9u 0f�	 �yB�CM��R�D?{�~A��ε:�~M�d+<�Ox�Oj�Z'�� �Ua�ݝ*�ă"Oz|ӡ*�]���H��� �5'(�S��y ^�NP2r��5� 	8V��$��>��O�i�F���*�p}���]��B1ps"ON���4����+���%������mr����Kx1�r��[�!��C0R芁�^<BP^1�f�W-!�  A�E���'X9�)��eɧG/�6�O�Q��
C{�ޜ��AC���u1O�b�(��)4�x�Bҷ_*t�V��a�$B�	��� 蓻+LA`��c6Ԣ<��R�FM`A�ʘ����:y���ȓ}P%S`O>z�l�S�կI8	���s�d�@ �DBl)"��-Q �X(r(D��a%jQ�~Q�(�2�bG�]��y�A��^�j���4F��1��͊��y�bE&-'���d_Dd0 p%j��y�L �^�Ӆ76�{�eп�y�`K��y؄ë/0��ғ�	5�y�.QT��]���E�"��![�W,�y�l]�v�X�I����QS)B,�y�U~�БJ@�td��i���y�jW56��xqj�-N��b����y���1t�lp{q�MN��R���yB�OY�bI��(��xq1� ���y���%�n���H:w"*�	�ڞ�y��c�2���HF6q(t��
-d!�d�c�\Ka�_�$���oS( 5!�O'аX��|P��Ή�H !��
�K�'Y#	,e�7��5t!�\q��e��iLX�X2��^4s!�܍&xF�Y%��&;�I�;SX!���??�f�"Ei������'AC5:�!�ϭcY�(�WS�V�Z��7"�!�Ѹf��T@�q���WAm$!�L�,2,���%<YA`�o�<�!�D[�s]��I�d�=.�,�j��T�{!�� ^9�҉�,�P	k��8��(	�"OD�@�J�%��A)�����"O��2EG��N��SҧH(�VQ9�"Ori���ȑ�@�B'�y#�"O���G�.��D�F���
�T��"Ojt��E�)���k�2��a�1"OR%��DY��v�B5�>��Q@G"O.��"�I>D!�3�%=��{F"O$Ff��f���.1�W�4r+!�B�=������# ��\�|!���P��z��� W	Xec�O��k�!�䚢Bڦ�2n�+��:�-�/!��æ�h`Su�X�Qe�J�� n-!�T3������V��e�8+!���3"c$8�GR�G�@��8w!���1{�(��B���(+�P֢.�!�D�*0X��&g�+������L�K@!� }�je!���|4f�	�c�!/!��]�(��1"L�h���X�a��T!�D��i�� �DQr�t�p�m�B�'��[���S��#TJ�0���'a�(��n�����z_���'a���,�=
nN���&n������`�4�Q�/Ha�Z��"�R@�!�[}����Ѝe�ޙɀ�J<FC!��w4I`j�2��,��D_;�!�ѵyL����Δkˢ�`̥aq!򤎟���p.�]� �ia"�}t!�r�ЕҐ�ȋC�j�2otd!�$
�=��M1�aЁ$�>A�a��h
!��1+��@Qk�pA7��p�!���P���Ң�Q|d����L�K!��o$p�ɖ	�9iEA0!���+8��!sO�0b�,<[A�%!�§De����W�4�1��� v!�d
�Q��Xe�ם-���Ćrw!򤋭 � ���� $L�D3t��En!�dj` �kRC��u	R�
��%Y]!�
W��2d��.�h4J!G�S^!�d�W�>t�+J�b)r�S��vK!�dy� a�q�]5%g��BS&A>!�d��SD�TGP�y O�*/�!�%"��[�i�6M���r/�7B�!�������
�)28B�;�X�M͡��7H�,u���ޗ���ɢ�yo��V;�h0�kإ%���R��8�yb��f� �!E@(�A�D!��y�!Y.4v���f_�o���2ģ���y�++xbm���'�*��τ�Py��TY�b�SP�Н~_�l���B�<!�	�-.޼S�	E�����R�<��m^�E�����q\��Q�f�H�<�%@7f6����E]�ڹ1�+�KܓX���5���sQ?����	��Y�-F�'wޤ��G!D���"�ƻ$Ŷ1��� ��L���;+�b�Sb,;?����~�����!�"d�nG�.��Vc
�_���-C}�����E��&��G(����gX�h�T�0/R�<�bmM-@z�	�H(�� <�
H8r㚤A%h�hwKĶ1'�����'�L���V	nd@h��%��M���	�o)��`�f�1O&��"�B�?����B�<R�Lʦ�S7fn hsF�&AL��'�"��")W�V��L�%� 6:V.x3M���Ћ@ h}�x���Z5P,���*����&Jl��]X3%]!C���#�#2����V�z��"T�[�3t�)�
���f��篝a�'�-��1Ǩ�д�Ҝs������*8[�OO �Ag�}�1�`�Ap}"�Ί9���(OҀZ�Kt&{�fΖ�r�ʔ�)�a}��A�}l�	�#�(䦌ktU6�Iҗ��;��Za^��(֩���D
;F�$�i�%~z�0ƔO�	#�G>@�]�U��]8�4IG��
�<�����G|�	U� �x�2t�B��Ă��l��� J�B%K/O0��чN+P�S%L"Uq��@B/x� �a2~�0�͒�=E�x�f���;���O�t����0hd!���,��}z �	�ߛ�C��-&�Ě#1���y�0A	���D��1/�z�O[��5{D�ʘM -�`�ۡ5����H�y`J83!U�7�p�c���;x�����E��FY2�F>'X����O����p�'mԗa��Q�W�)����1�v�(iKQ8��Á�ٍ��$я�,���:1�������R?Y �>!CC~?Q�"�=��3�fҲ��.��*�*I�FE	2��;��/O�<�D!_�.Д��49�Z���	l`��ʴ�.����;��$צ|jr����5as�U�tkǵ7jhY�w��K�ju+Vg��<�Ag���	�%�Ťx�U���E�	H���)ȓ=��[P��f�ڄ��/�;M��,�����a�u)<L�d%40#9�_�	�)g"��L]m[�"���9��䘏�:yI�/�Dx�I��gV�+���!HR3�M1t'Y�8s~���Y��F&~�,�0'N/0]�9���P�7��h�RϠ��`�<
��1c7""8��� ,	�a�[9X��CG��� �I���ԛ&+~�Xqc!><db�[�v���CVn۶<`=�C�B�4x�	���]X��"L�@����rDH�V���V�ԑf�A1�T�itb��$J���c�U��̅�D- $�[�<4��8�/ ��N�	���#"G�!�s��>�eC�,L6$�0�A	_K°���I�%b�h�E��`L9A�\\��挥)���㙍<8�Y6H��T'�l���"0<:7�mh�hEW �p�Ѕ� 4bɳ��D�3f�l@ԫ��U*	C0i'jx0q�&��@��MU�Ӳ �TP��`��7o�X8$KZ%R0%@�Ħh| !C&V:&��Hz�-�%6����4�B�=�f�k�O�홳Ã�2��iW�цHG�;?:)#a�8%�f�ۑ-Y�s����#�1��+b��>ֈ	p7������L��G��\�i������
�T���31�ϯK�\Q�������4��>1�L� �y��i�!�	HQ0��s��6n�����Z�y���TE��'4�!�jӘR�x ゞ�5ZFY����J�4xBNէ3�%�@F�wm�����¥1��u�a�Y."�ApEC�­��%����]ؕ�B�p>��)��z�A��'Ö��VI
N�0К�'P.�k,ɻh��,ٴ��/v�j�!Q�!Ȅ��	
Ӽ렪E q}��Kt+7�|�S (GE�<�  ��Pdf	C6.T�)���Ba�e�&HP"��T��� =��'u ����b1s�)\�F�HW�Y"K!�D%r4z݁��-pn�PW�mRpw��-q��ZWƋ�q<8(,M (����V�'���1-� i�]+p��g(`��C���@�U��*gcE&-�@A{sDH���gB�ssp�Ȕ54A���'0����S�A���=�����졀ԍ�a͈0H�y��jXP�g��1*����O&m����D:1d�S�L��@K�;�bp�_���ܨI"�t��-!�Ohae��L~�}�A��a!�l��m��S�<�G���ʝ+VB����t� Mz�e�!L��b$�f�{޽�t��s?��r��B#ft�5*O0y	�,͡l�X@/�;�0OS"��8�1�ϧ����3�<a1Ҽi2����`��Cz:��&.E�Eڴ��%m3��2�a�AS��<\O� �6�~ێ�C牒���t`��U~���AsD8X��`�,PC%���I��ǤRa��l@�?�zb���udK�m;����Q8,�x(��=�I�q8� P��/%VQ��7����	�T�2Ņ;̬���Ǎ�Qb!�
7H��p�[;+�n���`�%�p=���� EFޥ"P���(E�U���<ݤ(Ԅ�:���"dY~�����mJ!AÓz��?.H�y��_�߬ �&�6y��A�ɍ;?9���RK�q�<qcG�K;t�p`�3i��K�i)5r̴��c�`!����W���:��I9p� �aװn�����ߥQ7��������)F���X��i�$�S�
E��{�'G���`fd��r<2DP��N� Wb1��o� l*�$��@6� r��� ~�d8�v�{J<�@΢#Qn)�����i&�'�n8�B!REJ��q� $5z��ȁ�&}򀑀Ii��;ѣ��"Z6xBh�:���=2���e�'p@|,h`LY�p����GK�5XAz�$ ͂ISWm?u� G{�L��W��-y!�R�P��=qp8Rr`�Bc�4(Q(E
ݐ ���kUG.=�u�#ӆT��mڕw���%�=L ~\� 	Ŭ(���y��q�R�[z�T"=���IS¨���9��.��)s	�d�n���,n_�xЭ_�"��51fn���J��� ���i�e�h$�aůhT�(`=��IZw�5X���E�;f����C<OT���N/VZ�S�jʼ=��c>�C�*�?:��u2��'��(:�O��pdZVI$$�xA���r����P
�%b��m��O�"��Rg�ڟ�hP&��w��9a �00$NTj�ЙB1cs�H�⏃B�NM���+?$�X�J�f-�p�Nn�ޅzAc�w�Pu	CE�s���x�/S�!��,"�5?Jh@�
�@�*�R��#�(O�02r�16^��$���0OԀ��(��qH������I�$rd�H���{WĚ�8� ��Dh"5E¸�4�M<vG�7-Y�EXNY3:��⠀!ԴEq�)�6���¶�3/nft3u!��,J�q��nl� aO/Y�8�):H��b��	�؉B �'o����DHѦ]���9W�$�1$̔T{�$I�e���y���N|�q2��(O���"`Dđ�M+�	8M�$pX%��Y����˵��'/�Y�Dܕm�$9�"	ȹ�<�Hġьr�� ��")�����kÏ@�Pg�A�W�J���	:�"�04AO�	�@�U�Ս�$c�e�7	D�=O�I�[_ݾXiB�ܴz�Z��s��D�a�5� k�q�I�<L�q��%iQ
���dϋcǰ���fA	Xa�dʦ�AD�p���Ho�Dy�f�Zf�L�f% �]�f [��D5j��C`�7d��m��G�eP(!CF[���M;f�]�ncF�2g��{߶g��u��J,%Q�B{�5�$��if�i��dS0ZO�xY��>��W� �����O�\��S��
~�f@� �ZE�Y�%)D�:���7o� $�5�ۇ]�P����
|�h0p��]J�e��� X\Z�/�}��H��ꙂU��0cF�i�����Xl�B3 j�bʂ������J�e˚��D��+i�����ܙ�p)���<Nh�� ���N�ЭQA�V�����1�W�	f���Ti��'#$�ySI5��-x%g�I�<TK���5���Aè\TzԘ��7Q'(�1���2��(U�L�K�4@{Ţ�0�Ѷn\n�ڱ��`�:V�
U���h��=�&蝋��ܡ�
�)	v�l۔�T�+m�<��������B\�H�ZA��ˠ]ќt��  �y��O��/d��UI	����"�A���@N$�FK��E ҄�s�-ړ7h@�ϐ���*�5���'O�ܵz2+�-_�=�b˞U�" �t+�( ���E�Q�+��QՌ���V�}�h����(e���܍]���'��8��Kg����*�	b��mZ�Ȣ�r,�b��&clcf��C�@]��׬?�q�CH�a	�!i���/�d���ڕZ;��X���hO��"eC��VW�ȁ��K��a��S4��
�i���.�����:%��UQ��٦j�N�$��ˍ.T=�%{�W>^������:����P�0Xt��u.LOvx��o�.K�����"a2HB���<
�N���$O�:��0"��%F��J�Y@��K�'i<Tz�a <����;.�B��<bB|�&��7�џ�� j���B������8V��T"�D�5j�$� 3NN�-D�-b#!�)��AJ��"�=����d�EO�-	D��2E�ӿq���V�!}r��'���=�~R�ŜW�@!B.�V-�0��.teV�9�nՠ1�00UB�z�:�Yg&%�r��9��07�B\"�Ǌ�e��I�6�N@b��:	l =7+ނ[�r}[v�s�rU�_]�Ex&��,g��)��	P��%�1�̑S�gV���b��Kק�;��<Yp�޻2\T� �����+/S��3�/�a�ȬP�F�4�y���g��(�W���[�:�i�.G��%AF��z�ĳ?Ov�a��Y��heN�i��4��#����#D�<��+*m,Y�D�[����x��~�P,h%�$)� y���'�<�07��Ir�a���$���1�\�θ[�+�s�r��ZJ���	�H*�uH���'�yB�����CfX ;�x�Ȧ/B�y򤘩P�Hm
�D��5o�w!��y�씜P��#뎙x����n�*�yBDU�c�ٰSb�c��j�?�y�K���d��Ć�
A\bc(��y�`
Ov����G�B�=�c���y��ټPUx���h�'k�>@�v���y�h	jܮ�q��0kuJM3Uߘ�y(O4{�y@���gr��&��y2�	l���s�K�\�x��7G��yA�Ǌ�1�
�6(� ���aD�C�����bT�@7�� ��\rLZC��}�ڐ�则\<P�J���C��^V.�� �9�dاKX�+FB�
P��T�ǁ��>����s��o�HB�	9�
<�ҋA��B-��FI9]'B�I�\C�#���4X���r��u��C�����
C�W:�q�Wl�%��B�I�/|x"v�_���$�P��B�I�"w�9'* 	�N��ҙc�B��<%g,��tjI�!-t��P*,�^B�	� �������a|4��(��ED2B�	�*�l�1�,�#�z�	��I�B�I	�tʰÙ�d�C�Ov�B��UM�y�h��Q"�@(��ҊF��C�I�[�TT�ҁɉf4�����g��C�I��F*�Iy�����M�J��C䉪QS���C#����Qs��5r0�C�I!`�j��"�B�VgxX��GԐC��'8AZ�(@%��B�ĕ@��C�I$� �pL�]�H�Q��A�BC�I�8�p��G�H�vn�
fB�	�r�2-���K�\)�`J�O�C�ɣ!����D/m4�0��I1*�B�ɪgm I�Z/1�B�¦'��*��B�I�:�V\k�l�V@�fO�+y C��#�!���J??{ |ڕ޷�dB��_�8�8cFC��Q�^(p�!�D�#=A��A���5C���3hM�A�!�� 25�3�ݱD�D�sSj�'f.����"On�a�Y�X����2 �d��"Ox���JQ�q�΄jrȈ3|�`�{�"O���t�m�����'#.�5�"O,I�ϙ�6Hҥ�~���"Of��@P�htԀ�ŕ*_���*d"O@����Ճy�8�H$�T�)s�*O��s�.�
AD5ʥC������'JE)u�O�@�Xe �l\�O��S�'p����D6�|�gn;T����'�`�s!��-Ψ�9 �d�zЉ
�'\�E�TG
>L�d���]���� 
�'V�T����lDʩ���ķx�]��'|��@E�?��;4$U�i)�'/�@�eȁV�F��t�U@h<��'��i֡h-d������'�1Bà��BASD�#f�t�'�< �3+��B�â�i�ք9�'-�y�+��8;w��<\��9��'i�E��$��&�
��fQ�8MBM��'>��!�۾?qrM16�U*�:-��'cn��K�JM�i���Lw0�t��'�ZԘ7�zk �aRR,ŷh���'�$��`A�Aa�!�A��o�
���'���s�B Wnb�����] ��'���{2L\XT�sg�]��Z4#�'�N ���I:��;	/ ��
�'��đ��G�G�ڈ ���	��i�'�ū!�:lh\���h�pa�To�<у��B6@�#U W�n pf'�i�<y�Kߺyc���U)֬̤EӴ��~�<!g�K�:�b����ˮZ��L�׃Lv�<ᄦ�&��P���W�E4�m�@IYZ�<Qr���Aõ�����*��n�<yGڢ=:�bv�N'i���3�k�<�W	Q�\��%n�"Ġe�h�<r�A���sÎщzz�����&D�T�U�ݓV���Ӎ�q��9!7"D�HjU��13��#�h�[��[�j D�(ڕC����Y��:a`0�(�g>D�\����>�r�q`���@���+D�T �"^�
`���B$]���v-4D�@��C՜Q�c�%�+_�5�t�9D��C5a�-pQ��	r�Z�7�.�HF�4D�p�ötV�$�� .9��h&h3D����؍q�`����77s���B
"D��������aBW�U>y��a�,.D���է������QdJ��5�/D����OB/�Ba���&������9D��K�K��.�`��#lΞ	o��"�F:D��{V
�G���sCL���cq�'D��2�ǏG��BRF����1�k$D����H�J��4�3(;`�0j#�#D�<@�c\�3}&��`�	 e2A`�:D�(Ӏ�0*j0؂2�1
��s1�.D��9ǅ�%�J����Q�hX M9�	4�$��������d<�snT�fh4�Rgտ
y�eX"Orl�A*&�`� �_e,��ǧ��mJa��Px�8�g~R P��
3��GPBP�Q����x"�M�R��x7����Q����1�ؠu,��r'�-�C��
��$@4��)�b@�y+�/�
8a��@��G6�y;	˓s�|�qa�9�b��6b������@�FX���N<z���f"»Q���T���{��鍎"$}�"�?}R�XX-��#�6P#���!�����ODl���C�=&*Ak����f�r��&*��:�:���B�7��rfT��h���%c7t�
�/S���P%
�7�TI�G��>�j m0�S�? bab���.E[��s��,�vm9NפS���ĥ�9#ؚQW5�l}Z�)����{���<��c6oS n��iP���]�Z���o�<d�2��$ߡz��p�dIr�Z퐣�ǛE�P�#��J�5K����<InE,(剎>;~�a��:���	-R�H;5b
+�l=�J��p<qb-	q#������,Y�y2k4�x�z�!]�@�@B^/*{�A+ �(f;�	x���)w���]�����(ְU<��Wk
�y�4@��\8��ݱV,
�!7��1��	�:[� M:#��U��"{KK��s�H�l:!��q�ţ��N� � ��$�!{���a����.��a�"ME�)���ۘu��G|"�M,�,�yCF�k)*mB�x��
�(�2_v�&��'�d1���>�O�0��H~�d*�lrPř�[��#'@�%$�d��`7�O�����&g� 4���Z�Z�nP�SI��[ҒtB�K���fS�@[�I��P;��.r0ݻ��H�<h�e�tCd��d+#wF5��'o���b�/q��q`%�эU�D�hI)6��:��yz�Fc�L}��W)n'*�[�]��~�8D�@�F`���C�0�)�A�g��r� ��\t)ƭ�e��Uk�8�ě$�Jm�fHϲP���a`
)ʦiB�7m��$�I�Q��)bT�����u��S��K���A�$A;T�<�iu.3W��F|���1tb����	�9#_!x5+'�G/W��a@^0�v�eBW��M��2O���WC�@�z.�,g/��)�m=Ut�y��\�f�0�2��C�a~�X�/��В�(�%��aL`���UU`Al%�yB��1��ª.��y�����0��X�,�r�K�L#r�E8` �����	�G�H��B>4�|0���D�$��p�@^�Y+��D�_�{�@{-� u���b�L��ѷ�7"��,'�<_&�)��	����� �fNC�˨�i�o)$qO��G����)��	�vh �-��y(^�l9v�{�ĉ#� m�Q��p�y#��=C��yb�'B�I � ��c�h�?���^;paG�e�~؛#��b':7LF�H�$X2��z���,�E�lܺ�nɃ&ǔوW���f�F\DG�+4U�D��(�1i��{�Iv �J�'�R�㦢݃'�u�Uj�i �
��E8l)�=h��_�X����Ɓ��P�Z���" �i�%�O�j�2]c�I��*�4�d�I�Ҳ*�\�2T'/|O$!�r.@s�P����}+|AJV��,N����l��]�G�wD�+�
W�"����Z�e����e�٤Q��O�E��2Yvr((��;~[��U�"2�X� Of���p��u��8
�A6�b����A�j@!�y��|�wJ��}��I��Q��|����n<�4�X4<"<L��"M�U���y��F3L�M��C�(ޘ`��\�v��N�:.*h���͈�yg%ŲD"r}1�ޚ)Z�5����y�h�8��2���?_�I{�ϊ1!���ɣHO�g��\�C�\62�4��^�+Ō��qq�`K	)�� ��(B䉩��r�ʊ#D�!dB �ʽ�Џ������G/�HB��)��2P�ɛq ��a�E2>@� i��ټy�N����,G��_#Uc�%0g�F)c��y�-\#rHٱ�  Rd��������ɥ7�
 CT��hOT��LT;nA�V�;;J�T�nn�$L&��V�ez��2wmI�m���y�����LT�4A�"Z;M:�:�
x�b�ae��*������熀�p��K�t��t��'<ȴ2��ɫ���ش(�L0-x�쟄��@.�H�x�� s�t��;h.@�!lΐNb؊��.z(��C��F�J1\{<�:)�<�̭!X�jM�(�%���'����@��lڗd��D��� q.�{c(\�I0��A,:�X�%b�P[$�8
�(Ur��D�O<��p*-p ����	N��u:���^���r�"J�]k֕�TI�064��ŉ[�s&���'��'x�<Aal�=lm tKw��L����{��@�S�m��GH�d��M#s`[��u �?t��x���o��q��"N:m�l��ՠ,T�����[*�+�*\O��`+�8�y[�l�/d�*@q�ǁ�������Z4C�T�r��W|��+��<�I3D̕,b�8\Q�����=@��Js/:\���:�tx "O�ˆ,P�>Lĸ�v)��p��i��Q�n���3�h�j�'��#%��֬о?HМҦ�Wv��Y��wʸɈF�Q�Z���g�])yX���'�L�ð����zp{�������(�2�ǐ��!A+Ȝ]������r5n@����e��8OB��f��v���&� R�pc�3�L�jM�}���V�N�Q�l)�O.i���DBT��n�Ava���M�D.ΝF+Ziяםa����TX�DICQ#^9�C� �'�uK�OF�e5�	�BT >��@��50�v`�c��,@7mق@2��F��-�l0����-X�m:$�ǿkj�E���k!�Y��XZ�����I �k�r���b�-�'Ba6	 �0��w�)�tBĆ���uhCK�w��M��PH�Oƛ��8{F�2��|�l��'>�d�	�<���
4-֯*?b��BcK�.Ea�ʯA�f���cW,(;�xف��ɲ�b䍗,,2xݢ��xB��R�b�XETt�{u���<!1�ϐ>wP��efA�_n��-Ƙ��$�3G�" �z���-ƈJ9*����tt�Zb	���|��D#S
��AP˓PPȲ&d]4Y"
=Fk/Zyr-	U��hK�q��� g�,��e�WN������_)	j�������Ë[�0:�効���DKQ�@<rm�A-3$��{���?���7	P0[�L����90T����P}��կdӲ� '���sz�1�CS#g��P��μ��&��yY�m`fK�VG0�;�G8��DH"'<�q��V!L{>�bl������6!7b��g�-�H�z!Aџ|��@C�C�Kt 0���E-�O�t� փ}8�<�"��($Ԡ4��H�P� � z7���CM�/:���!��)� ztz�b�,\�؃e�[�m��(Q	�%r!D	�R�ο\���f�-<O�Y	��n�H� M^/
#�p�D)��d�&��'�����b�M��eqI�?i�|�m��	$�l�4���Q�0�2B�HгEf�D�22"Or-{� Ӟh��#sE�OAP �7�1P,�)1�N�1QL�T�}Z~5KŠSl��c�%U2HNN<��5�T��t� *Ӓ!x6�
 &6șP�'BJ|�C�U��P`Zԡ@�K�R����
c4񯕧A���
w� L������L]"$A�L�L�`�}R� L9���gM?�vq��"J!�hO@��T ��o�2�1o�8ZS�𢨅�K.u��at&���C�t� ��|��yBZ�
I2 ��>U�1��S6svT4�M�!�"��أL,Mkׇ��D���a�C�Z��D ��t{p(T(�X�D�PVO����h��G]=g����'��Z�g����|jf@�\?0|��
-rt5���c����Â4y��kc2)� ,��ϻ���Q����t��,Q�����	(AA�9XU�X�>]C"$�(!N�l_�= ��Q�"M,�jB ���I��A��:qG{�d�Q`�foI 2���@��Or�;5�Ƹc�$j#Ox:�P�8T�2����M�7�$а�O��u|�a�P
��m�db3�'���S,��"Ua��qw^ȮO��h0`����[{��Ǚ$8 �5j·F��S:��|�cH���$�Z���1�C�I�dt�8��]�5D0�	����B|�)+��ɠm��$R�rti��8�)��q~y��O|��h:�u�b!Ղ�b�"O"��NL(Xx�!፷(;�y
��"�Ԭ�5�V�X����r^Ȭ1����>T�'��;SX� u��*Tn�y2��:P_�8h�튨Pf�@���unPU���fO�I[��>IA�&5�O�qd���0�BZ8�ճ��ĂX>�ɋ�JњD�l����{� r�I�B�8��p CC�}�H����@fC �5$`4x��)Cjּ��*Xg0dzsB�y��j�����>^B9�� c��Q�q? !��_�`��h�ha�\�����5z�6��/�]b�X+��=���Z85�D٨@��2$Ɛ�X��PL��(KBL������F���S��vu~t@���I/�x�ȓd۪%Å���I��Usqn��l�~A��-�,��V"ڽPWbѢ�j\4\�����n��ݻ���^��z���ԅȓ	}�)E�8x���b�(֩^G�d�ȓ>�Ь@h��(�����J�af*(��b�����$GR��DL"?=@݆�z
b��Qvr����t�ه�\���6"^&jMV�u�ߧn���M��Q�e�N���@��S�j5��1�Hp���&�&��ue�5�U��1#�hJ3nS�0�t)�v��2[�B��~r<�HJ�9�ؐ��l�0^�`�ȓ��Aф�,<��aYW�'x���ZT��pTȆ(o��Y�fl��0��]�� S���#�	%L �g���HVH���
�BT�Q%��!I�u��LZ�X���ȓ&�ļ��ʥPʰ�`��<D��ȓj�	���,4����F��00d1�ȓmѦ,ɳ�ɻ+�Ѱ���Bj���e������3,Q���"�<C����7�<\��mAd��P�T46�<m��c�1�ԯ�"���2 �����*z<����6t����Q/I�Q�ȓ�(��R�c�����F	�j���08ʌ:���`y�ȁ��V�dT@-��! i��M!�$��aM�6K+��ȓQߒ��T�#+*P�`R.I#,}�ȓ@fҐі�Ⱦm�HQ�AY3:r��ȓp��Ż�b58!��'�ҒM����U�8eƎ�vz��F�ԻD���ȓ[a`H�Ӣ�Q��2��Z�#���ȓ��}���!x`�4���$)���ȓb��miԬ7�U{�'\�<��ȓZ\�`6�H�aJ�Cp��"����E��d�`i� ��АR#,fJ�Q��S�? �<r����0�FHNE��5"Oa���ȸ0��A;�g�.�EZR"O(Y�$O�l'��kE�Y���a"O:�a5��u;���喕I��A�4"O�-����h�V���Í�rs>��u"OT����6Xkr8�v��>V��*�"Or�C�/���5�p���r"O�a�$EX}980PA�]<�Y�"O|(
3eT�\�| ��anTS�"OZ`;����x�n
�D
A��c"OJ�"$���h�)��^�y�A�"O&�j$�� q� �����#�&T�w"O��b<{��u�T��@�+2"Ofm���57�����#�h��"OV����?.Uzu��� u��Y�"Oxp B�Y$+WZ�2`�?z:Q�"O�Q'�۝U`Jd��ѕ+b6�4"O�q(��]�T}ސ�d`R�DD��З"O�@@��Ԏ3��=��m��'��""O�a �и !t������j�(��V"O�@���&��$��K�k2!�X�P�|X�KՎ��mP1.	!��J1���p�=��U���x!�Ք3�N4`C���i����-K^�!�$ɕ 7=���h�Ւ�l3!�AN%z�� Q]X�SK��%'!��F��]!`��bn�=�'�ݛ*c!�dH�S�����Ckb^�x AC<Da!�� r� �x�'Y�hi���f̗#T!�D�� d2��&��S��H�qO��R�i��,q���8u�Hk��'k�O�i��ɚz�
��֧�r��I�@�4zlf��ɞ�M+@N�񟬑V���������CH|��/�+1U�@6	��a%��4l� �yB%H�`�r}F�J�A�	D��ODԱ2�w!��̠)�@E8�l;E�Dй"�� h��(Dy����;cإ`�芗2�Fj��.~�x��'��v��|�'��	�ᓯ&��R��� ��8��	T�J����p�X����S(�r�~�L?�31`ي7i��*�-N�\�������	:	Խ'#I���Sܧ/�0�G�*��aI��E�m�Ֆ'�",*�YD�O�O���@
�5�ТP&gW���׍2#��=	��,azf利�����}�q��֝�˴s �+��%�+K�|J���l0�t����83X���j #D(�0�T�(1��;[h�b���'=(��0dsad�H+B�,x��=)�'�.p-�vܧ�ħo���c�&��s��H��=��'��1�
�7{!l�'�b?��%�ǋ?@4`�!�uQrPa�>I�A��z��J>E���U����&!�l��%C��M#砑�\�&@yI>E����z��C��FIp$��B���W��y�	�0|`lO�>m��k�C�,���@#R����O��P�?�D�T���5 �i�!C���u�A%��!�(�o��t'�b?-����5r ����I"�����P��!&�5�>�Od#�d����OD/3��2wGC.��=B������CF�X��h ӕ�"��LQ��cdB9>D�l��m�y�v��a8}"o��0|R�l�V0x� Rh��J]��:&��ʴO��el����a�|�hՌM�����ɪ|^���fm�l�>\`�����Oz��� ��.��BA�o��)�E L&C�������)*��^�S��b	�/`|�%`�#� 	Y���y2�Ŭ0:�Š�D]n���X�yrI�|��KDoB�S��m�c���y�ɉ�X7~|yg�ρ|i޹��i�#�yB�!R�I�5��D�Ir*���y)I6}*����FХ7����aj�y�gB�lB��'Ƃ�.�r	ފ�y�k$D9nDr��U4�Y�B��y��O)q�h갫4XU@�I�'��y�C�h>D��`��U�TQB���y2E��w$��
ɚ~�x�����y
� ꀐ��*7*	��6,�ĔG"O�pI��ňa���DnR"c����"O�%��e�>FFrV�4F���2"O2 �����А��H�2q��i�"O�#�T�zy�F�@�d��D"OJ�3VƬN�ܐ�+��!~�AC"Ob��$�?yo��kgKE/���R*O������DZ�9z���	O���'U���0,H%N/tl���Y�KZ 0	�'фe�ɒ#S�jxi��#R��� �'���h��AdA`��E�n��'�����8R��âm��<^��'xc�B�s��=�jA�1�>��'�5	Ť�Eo D��.:Ƞ��	�'�&=9��Ѽy���H��P3�H���'��@���6 �BI�f��:}�f|r�'N�E@sf�6��t�To���'�< 8�$X@t"Lǔ�Xf��'; (���Ӽ>TB}��圔W���'������F�/!x� p���t��'���Ã��1.�xQ��������'^:H��QM"ʈ���O� X~���'�A�&�Դ�$J	�g=�̫�'ߤ���,�g�:E�kD�\4L�']�y�',؃%80�"h�&Rj4I��'���Zs� >�|SQ���3�$q��'m4X�١!�j #�J��T����'b~� k��l�@���״EE�9��'��t2r�U5qQ�T��Lͯj�L��'ՊY �9L��jb(�e��Щ�'�P�n��_�tP��ù_�t���'Ej5h�� ���_���0�'`r��͒�0�����#[��`�'��H@5�\�7(`�R��(Q���	�'�~` �X�Z:�I�s�`�s�'�h��U��2�bH#�h�(��	�'��=���QIZ���F�	����'@F��#��v��8�Q�ڦ�$�b�'�Qau$��*�<\�p��"x�����'~��6�Ýxt����v��@�'��Cub]W����A��P��'WN�*��g��`���`}3�'gYX!���UPղ�*�6�F}��',4��TAȕ#��47Iʮ.��t�ȓ�J�Yb�N�w*l�$:�Z@�ȓ(���&+��Q�LP��m�7F㐽�ȓ�~� n:o���AUn��q��n� �b�q�L�S��~\D��,����c� 7N���*B.d�y��|	6�7@ ��[ ��)�\����E����;y.���Ӧ2�<����|DHe�<90i���Q�p\��n�$Ղ����P�s����xn�9����Pap��S(�x�6�J���؆ȓC%F�3Ǫ˂>>.L��ęO�X�ȓ3��r�*�������GL�^w����E�h�Y�(���`@�N�vXr��(@ �BR�����i h��ȓ`��<��aޯN]�k�����ȓ3x�q�g�%W� n�p�ȓ)�xc�GM$of>Ac��P'lX�݆�"�]����S3����� hr�y�ȓK��=�`��;���R	�iav��ȓCiԄ��$ŷ"�8,���^�r����S�? R�hv+֑i3��6A rl�jQ"O���3e^�;��)��	��i��"O��H���N�d0Q �	>�L(�"O(q6�<{�J�t���H��� �"Od�է���	㆘�{��Eؒ"OT(�׃��#\l12�f]'pjY�"O(�fe_:(��K1H	RB9�"O��r`f�4)r�f�4/��h��"Ox�9B*�����䄚�<�9`"Oz�*� ?dV��rv��	�0 ��"O�(x�l��m(l���S@�N��"O�g��C�,a����3X̊�R"O��`W�[	j��� �M�R��)��"OR�2Bٮu�<|A�KA I�FP:a"O��3 �W�
���Ӆ������#"O�<ac��3Imz���	6�&D"�"O~�ӳ�
�a���@	�	.��`��"O��y⌟�TR����F�Ex���"O�ҋ� =�� ���ap�)V"O�d�#�n>�����5MN� $"O�8��NW92��5��ܶQlF\3P"Obpb�NB;)�Pk�F[�K��g"O���-n{�I��k^�X(Ȁ"OnX`��^:s���q���a""O*E)��Il�a$K99� �1"O x�՘H�2t�b��*'@E�"O��8ᮏ�#�Z��f!�/t��k%"O��#3(�/^��-:�ύ� l���"O�h@i_)2�Hm�a
0��S"O�m@0���]F.�y�Mׅ)�z0I�"O5�6CR�U�Y��\1!���C"Oހ+�J���5���n��P"O��)D"Z����K�g/v$	v"OX ���?~]�p॑� �`�b"O^�8B�q�D��U�,�ڵPu"O*��cT:oC��xG5�n�J�"O4� ǎ0fUZQ�5SĞde"OMAF́ x�@#�A_��Iy "O��*�/ܤL��(#`��iXԹf"Ov�Ȱ���Tɢ�0�kPNB 谣"O���ㅎrS~p��ɄA2,1�"O�p��PA�\l�.h���E"Ov�VG�+~!
�j#l�1)�c6"O<8�"Q�
�t�R�K�3T�Ar"O��3��9��Q�<!<2-��"O"p3���|\4p3T�. h���"O&h�V��)*7��҄�F�Q|�b�"O8T�T�;�@�q'��wd`�'"Oz �t��"@�j��%F؂��X��"O��6*�9��|�u�� ����"O�l��,��Wx�|9�Ǝ������"OԘS�͐&�ty
��ҋ@��	P�"Ox8�aO�Eh"Ŋ��^�g�8�r"O�tÀ�ðn
���e瀏�����"O�	�Fϋ+кݻ�F�2I�R�zS"O85ѧc�a��R�L��5k�"O�%�����l�TQ��o��Q�4U@%"O�Pr	�6&��q���
`�VɄ"O̅��ٖ���k���.	�ؐ@q"O�����o$��G˖>���AG"OԖAz}�^�3��-J岼�'�Ĉj��<P�ʁ�!�2m���
�'��,�N�"��H�ӯA�1����
�'d<\���80�ҽ��^�'x|�

��� ���!� �5eN)z&���cM`��"O@x;��X�jJ<���*F:v"O0��A� ���1� I���"O��àB�f@2�0SO]�8g$4��"O���aҸ+��r��Mm�""O��X��vc�03��O"m�}�G"O(57cچ}��I ��!N�}��"O����X|�1�
�`E�I@�"O��г�z�8GjK�t<�4"O��KR�Ĳ/����aIB@����"O ���H@�%0�d��ʰX�f���"Oji��)�����^�c�>���"O8婦�J�;R zw�52�n��5"O
AW�!���[�`�%�x�5"O$r�lvJ����.i��\�O�<9a⒫j������R����M�M�<��_�&1����ȓF���x��G�<�&�ʪ/B2�c�oT���b�MA�<9���2�X��F�_�YP��ʣ�}�<�uEI�\�4L����J�ʠ�$Oe�<�FH2z��B��
	�6	�G�X�<I�l��P�P��J�dG��2�)�M�<�Ą�����`��Lv��iB�@�<��	*T}:������d�JV�<ё
 lv 0������ ���l�<QD�;��j��.���!��]�>	�aZ���' )��L�!�$��,�FY��.���4nF�T7!��]�+�د+q�]�A/��V�!�ֶL��)㥑�-�htA� ��!�d�>�,bR�#@u��A�)?a�!��U$ ��P�q�	�J�4�GI�Q�!�$�5 �Ќ1�)'7���b��e�!�$��/="��t�_�M�� 7��/�!�ċ�:�F�
U���č�2H��t�!�d˯j�H�{"����RsUg	�~�!� ����4F�����GT7�!��9\�B���Q+Z �!h�0K�!�͏bX���=@K2�O�e\!򤏲AF$���N�06Dm�g�^�fW!�Ć�_mf��d�X�U��5�>"!�+O���9��87 �KD W5z�!�D�=�N��@�A4n!��1��W4!�d�T�8����.徴{�Ν;l!��K��#,�K��z.a�!�dP�j��l��M�p�$r.ߕ8�!�̤���R�m�tc4x!���]�!��)'.(ia�
@���1��T�su!��O1W�F�9�&F%o��)��$��s!�)М�`�܂�0�CƐ`N!�Dm6�$YV&���+�ϥ5!�ޗGKT@�2'W�k�2lҢ��9F!�$��NU��1��F�%�2��c@�F�!򄄠�Vh
C�!q��-��Ď��!������j�0��,핚xU!��J�r�L��5�
��̔XuM�l^!�D�'ʹȲ����������HA!�D�(ۀ�ȩ��Ȣ3ˇ�$�!�Ě�]�	��
�>����	Q�
�!�6h `  ��     �    �  �+  �6  AA  �K  U  �_  Wk  �q  \x  �~  �  ]�  ��  ݗ  !�  d�  ��  �  +�  n�  ��  ��  2�  ��  �  ��  r�  >�  �  s	 $  �% �+ ;2 z6  Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�� |d��"O
`�(�;���8���-0��1%"Oj4��ND^[��"3/9�0|H�"OB���H��*�ʞRy=a"O�味V�!X��!&F�:J�$���"O,��a
���C�Ą�M�"O,$3%o�-���p���+Ն�:1"O��ݢ1����`���y14]2��i�<�6��{_���c�H�`�fX�$Kn�<��A̼VI�xR[�)�Ć�pඤ�ȓA5��('nߡ4�� �)˩%� ���,��r�؊b#`T�eT09���ȓ!�b��g��}�8�F��-? �ȓ
K|m�ș�VṔ���2�%�ȓ"R�X�j�4JN�1�˘X�i����̹	_�jZ��1!g��zܶ��ȓgil,*�J�
j�Ne��i�J%b���f	�(U��:���G��$Y^م�~r�� S�%T"���k\�jx�ȓ|4�1�îJb��@ӵ�ݩn�V��/[`�"�v4�R�!ʎ<��M�ȓ`:��z�ؚh�J�Z��$HY:	��H��p�m�C1��!��B:��0��EnjZA V;9����J[
2���	��4'J�EA�IVW&��~�(aZ��ӹ�>� o�Y�|�ȓ�f�A�
Ο7�H��M�$�����mޠP����/���ANXo*�ȓTv�����{ ��-7�*h��I��sB�8�8���3����ȓNe*M�悡;������X�o��!�ȓ'lj�#F�m�+R&;�|��2)n�C��0S4���T:
b���:�0!��e֊��)��ͷV��,�ȓ0�&�8#���� ع�L�����;�P�AFd���,w�6d��r�EQ�( �gVlɦ�M,H��,DP���|�I	$G#\���ȓ"�)���E�B	yt&B�^�LɅ�4�� ��eëF�ڙ��n��RbpEz"�'a$aѴ-?�@@�A� ���
�'_䱡f)
L{PԒA�\35�l��OH��՚EK�m�6&Q�/�ؑ���5ўD��S,y�E@���y�H�v�B��Jr !2��dar)��c�*�BV$D��� X��řu�ݶap@{1n,D�� dk��#��a�V#[;���+D�dBsʀ���i�u��!;�-�0
>D����	�BL2)� V�bx���D'D���^
a��{qB(X����A#��h�����E[NyC���3/��'�-D�`���Ӹ3��W��{3dm2�
V0�yR��K��b���w�� �i۠��<A���:p-�����u�R5�A½R�!��X���䍏�<��4�g�şP�!�D֑sD�s!��Yh�,A���4�!�$I2p��mЛnr�G��u�!�Ċ�>H���J�Bkr�s� ���$u�PXv'=�q�ӊ��3|=Hb"O�ّ%�4;���1�*�5��*c�'m�O.�lگ"̩�K�"�1!.G#�.�'!ў�?��s"W�М�b��N3]e�u�d�<Q��*�g�? "���(��M80F�)��h��0|O�#���Z�VIBĚ�#ͺH�'�>����I2i�&|zΘ�{�\,3t"��@7C�	,;j��f4�z�K��U�<��"?Q�}90��1f�.d֊t�7��pB�I�L��4�ҔY�]'�(V���hO�>���Å$A�P����e���S�4D�0�`d\�v�r�b$1L�F|��=D�(Y�NĐxPP)�R�Y�t��U:�Obʓ�9����q6 uy��8,J$(��R�=�£X�}��p���^8�!�'a�~�ꋻ,�lx����`���y��߮2��YZ�KM�!`>x+p�67o����,8���'�X9�EO�{�az��iq1OF;D�'avI�ŭQ' ۢ�⷟|��'�,���/D�i�|a#� rOJ|���$(�S��`I�~�"	zШ�eR$�� L�y¢.+<�R2�Z�8����Х�ē�p>I(G�x�" !Y\;�[�kS�<q���FL�#E$]2>j�9�ef�e�<��iG$��-quJ#0��*&�\{�<9�΍�B�9��M�9����v�<�`��&��X��
	U�(��"Mt�'�*��i��n���S�� N~�P�Hؘf!�D�-"�h$a�
]M�����&7�d6�S�O�80 P$·-iZT��Ɋ�0�p���'�z�����05��)9aÊ2$ۈ��
�'���dH��(	�,{0�O�G��4듗�I�S.D���?y#�#� C/��B�	�B皬s��U+$]��5H�.0��a?q��T?=�go��=��A0g�ܸ<o�ݓ j9�O����IH�-m� {F�6.�k"O��A _'�R�rBZ
�� �B�I����ʁ�4�L48�|8Gǆ�f��"Oԉ�$�X�ĭ	&�]��`�2\�p��)�I�<�I�4���(E�B���I��d�<�QfF�Q�Di��ƈ�%�pI$�a�<��͂�rU)� >&���B�u(<��4cb�lR�_�+�.i�U&C3!|M�ȓiL���i
I�z\��D#[�H���	F�'n�����fr����ǡk�T$�N<� bÏ�p=񂁆�q2e�]-v
|���EM}��)ҧ@e�5�øIlz`¶���>���ȓ	�HҒGX��"���\T�G�SW�*4� K-=Ў`�%��3��C��^
�b�l8&hT[b�N�zC��*�����B�0�@��� �%V�rC�I8mt}��^8XJ����eB=z��B�2�Pl9��af�����K4�B�2�H�O�q�ē�#��a;VB�I�[& A8�aI����"�	��jB�I�
fy��C��B/�D�UM�/g~B�I�q&��(��lx�c�K\=e�C�	*T�N�9�GU�HM�tN��XC�I�Wq���S�4�HE���8�B�ɳi% �h�)͊CQ!�c�ԮD�nB�Ij&8� C�^��DK1�̈́M\B䉹	.a�I�q�n�vE 
?�X�<�˓ @��N�>v�q``�Q��m�ȓ+� c$+�8��|�7�C�L���&@�m�G܀S���р��|�pd�ȓx��0�@�ݿi� rT�L��H�ȓ^��P`��-Nb�!�Ô(,����hO�>A@=kri�'�͝���X�<D�� `l��BEԻ:�@�I��'n�	7%K֤j%aX!b�|���)�=��C�Ɇ;�Y�2���r~QcN�9��#>�5��k�r8 ��,	Ю��4WNpC䉍6�z��0�F2P�4{��@�Z�:C�I���)ʢ���1�v�`��q_TC�I=`�b����h�Dl�� 7T�~B�ɊK��C#U�Gi<�zǠ�,E�hB䉦o�va��V�LI�`�YQ�2B��%j��yi5�I9|	cB�!E`B�j}J0CA&x!A�F&B�ɑv�`�bG�H��?(�Q�ȓ-��Ͳ!���5PDS�b��х�\�'�ظ�ńR6a�2�!�A��oJF���'̸`9�N��X�`�p�H�0m������'��H���*6����J�f/���'1���1�Q	G��x{S-��N(�i8�'�� x"�
�b2����Y�X n�`�'H�)�b��	E����
K�Z���'��Ԃ�P	F�2ac�I�HEv��'�	�W� L!�0��S����'�h ÅCY���u�\Zrl�'C|Ջ$ˉR��M���H�O�dh��'�Z� �E
0��G�Gw�UA�'* 5���	p7��+t���G�d �
�'�P�g����x�VMS9\�
�'I,�!�n�%=�%��\���'1�1Y�/J<��Ù�[���S
�'�� q����R�̉�C&P�R�"��	�'3��B5j�|�ac���U�f���'&mY�*��,�H0B�n�N�Z��'XH��	e�E��˘�u�X�	�'�d*�,4��!��셾^d��'cօ3�	\8%)���Y��P�'����ʏ�[t�Y �Y,Q�T)�'�xez�㒐0�� �Ğx�4�+
�'�z�Hd`F�[Lձ� (��-
�'ML%�w�ѯW�tȘ�͙6ђ��'�x0$�L� �QH#��/�Nщ�'��|B�aq��Y��C�)||h
�'��i���Ӌn~Q��cK6&����'j����)O��l�r�&q�|�'
6�;���R�H�����/ �� �'{4��D�B4u��D�.j��'
�J�����`ta3B�4G�yO
/}�F81CŌ�|�J�!�*���yr�	bPN�.N�v�r��H�y�ܽS0��S ��8tR�J�%T��yb�A$�ER��ȑm���1 L#�yB�ͭ/�PS�i >i���kY�y҅J�<Ø��1h��X2L�$���y�z���e�M�,��\7F��B䉡4	j�0�&SfXP�G�4svC䉰,�̝Zfj�/��Q� 2�LC�	�KNf��� S$D��c��J�2C�I-�^YR-�7����D˂_�B�I�ra<pA����5�X�UN�/�C䉼v>)�UH��5��%�-V��C�	,!0<����JӠ��	��Vy~C�ɥQӢ�)��؎^{��ڥ
P�C�� D�*G�F3�pYr���,3�B�	p�R�c�I�$;�:e�c P9;��C䉠4%l���?��B�	2v��C�I,s��I�E�W7S[��YÌ��>KHC�)� �X8�� rc��ca�>qҬ��6"O^��L�q�j�YCnT�_-pA�"O|K'�q�X�I��T7&.)C�"O(U�p+�)��$��lP�L{����"O���ۑ!��H��A�1G��6�'�r�'���'�r�'�R�'`r�'�NE��`�=k9�@P�_�0u�[��'��'�"�')R�'v��'3��'Z��%�ɹ �<ܠ��S���Ғ�'#r�'���'J"�'�2�'��'* \�^&m?�Aj�_�8��Ѧ�'�2�'���'N��'L��'�b�'�lX��=O�H��/O6jV&a�V�'���'���'���'���'h2�'�慩���"F����K�J ���')r�'�"�'��'.b�':��'g�}��1�+�9v����C<j"�'���'>��'���'��'`©V�R���
�n˛ZF�X�C:)b�'��':��'���'LR�'#�	5��{eO[�
�(�`,�0&%2�'��'�"�'�'u��'/���7�֝!F&�u^`�b6*@��y��'yR�'���'�"�'H��'m�3C��Q�W�qY�!�I���'�"�'���';2�'o��'�#%pf���QB\6�!�Da�����?���?i���?����?)��?���;�D��S�!	���HJ�]�����?���?���?!��?�i{"�'�~��W;0�-�p���\jh�ç<�����ش�D;�
L[^�mJ�*�+�hհ���q~�oӮ��"�4���Z��e�����DP���ђA]̥ ��$�M������!��<���-.�`��޽&���'���Rf�Q1*�]���k�V�;�y��'���e�Ol��U�9����E*"���Ee�j]H��-���Mϻ+4�]��Ȍ/UQP�*��ܷ?��T�i�7�w��֧�O�015!�y�	F�a��DjwW�]� �8�GI�yR,MqOd���Ҝczў���T�ؓ'*iR6��;i�zp���8�'��'rx6M�2�1OD�+�O�xC09P٣d�I"n$�ɾ���	kڴ�yrQ� c���1~\�9B��8�����:?!��	�z9���D͑ŗF3��$훲�?�4l�:T����	W��X%��ɂ����<��S��y�b^�WB��hS�Tc�������y�j�
�r ��x)�4����tGݦ6/��r��;);�ܒ��y��mӎ�l�˟�h�]�u���d.� ȁ�8씵�7O�N��X��e�+�AǱ@�Գ�Ñ2o@���ӻlLl�.C8-D����$MDMkWC»\�k,۽OB�l(���]'��*��I?+�!�dN��0|�2�O�&��ť�:i��,`��B�-s�����$S@r�s����r��sd�C���D��0}Ƅ̠-A�E�V9h�MR�S(�)և��iq�t�뛞|���Yƃ��ka�xV&L�q��Y�fHY� ��ZW�����S�g��6̉0�B���p�>l�,1[�n�Z��ہh,U���i�r�'mR�O�~�
7:�H��Te�`+(t��dn���ɽ16���x��Ο��i�iŘ%Tr����,��	��"�!]����r@��'�R�'|�$�'"Y>u�R�p���V��P�T�XU�<�Ms�`H>&T�<E�t�'�2�fT�_uz@�1aВNl�H��e�x��O,�D��!����i�O��ɬi�n�jv�Ή9 	[��%
	�1a�y�	Ѫ�L�����ON�$�-G5P����XJ�8�ɶn��a�-�'�:����'2�]����g�I
Wi�е���\P켑Bo��c�1
�O�Y��R���ڟ��I�L�I�d��, 8�۔�L&����`�C&���'��	���&���I��8c��ǧ�$ɢj�{ء���#A���1�??���?���?	�F��k�O�`��`�%������uvظ۴�?����?�L>���?�Dk�d�*<oZ>$���i�'�XN �XĥU�j��ꓕ?����?����?���/�?����?է�Q�qg�&e�tqQV)��&U�6�'#�'L"�'��53T�C��ē�����Sc&�a�I"
?�m�����zy2�	b�����kl�?w�be
b�e��i0���K���^�(�	ßp�1�4�ßT�s�p4���L��b1" U�h%ļ��i^剨4�`�0ٴ�ǟ8�ӳ���W�2���"V�ͨM8A��[+^t�F�'��&U�i>�I�?O[�R�}�څa�T�#P��i���㐣x�^���O��$���'��S$v�	Z��	b�]��JJ9��iݴ2����'��I`�s�l�I�U��Y�o>����Q	q\�2ݴ�?A���?�ud�-����'�"�'����u���oF��t+S�qi��S.�1��$�<1�cBu~�O"�'����!��0�]��P)�c�($7m�O�Tkp+Iڦ�����H��ϟdI��Z�	
��P�n�?���3�M�n���s8����?����?��?�.���3v�ߘv�h@�-]��<���YVj�mZ͟p�	ş�����i�<A��צhÀ�C�΄0ׯW*n�:h�'R�<����?1���?�����		�;� �nZ,��:d��{�|0�'�B44f`��ܴ�?����?	���?�-O��D��O��)�!~^سW%шW��i NA-Ln�˟<�f������I_"V��m���	{JޡR� �4�$�ӏA�nBBݪش�?����?1(O��d�*B� }Bl��'�Y�㎖4��	���M����?�*O��s�ĐN�4�'Cr�O~rQF�ߓu�D�Ap�ʹ
�����>���?Y���4@ϓ��N��3� F���� .��0B+_�i�F<�F�i��ɼp�8�ܴ�?����?��'h��i��ѳ���X��W�	�D���s�t�d�O.ԣ�4OR�O,�>Q�U�Wm����N�j�*#'vӀ5�1*��Y�	ğ��	�?�I�O0ʓ&XJ*��R�6���G<4�����i�r���'��'���d�!#������ �}��g=�m۟��I��
@
���Mk��?����?�Ӻ�q�������w�C�R�p�*�˦$�0���f��'�?������V b},qHa̗$����-�MS�t�X�r��i-"�' ��'����~�f�Z���5%X�����	�?��d�+)��d�O��D�OZ��O�˧k��Ȑ&D!9j���o3�0� G�pj�6�'-��'#O�~�.OD��B�B�ʙ;��P�n�!��u��=I�;O�$�O\���Oj�D�O��d��@�00m9sL�۵a��e������K18���4�?y��?i��?�/O��c����.t����#M��`��f�W���'���'���'�b&Z�J�F6��O ���R�5)sI�&�ΡrG��0�6!n������|�'�Rʬm��f?I���+q�����#?�PI���Ŧ1����x�I�(2f!�M#��?	����
	%X;�=+`�[�p��с!��)���'��I̟T;$s>�'��s��h�p�ԺE��g���)�\X�ķi��'V�yz��tӠ���O(�D����)�Oҝ��+F<]$QrA��\�*�¥u}2�'
mKD�'^S��e�酐En$(˖�ްVd�P���k��c�ct6M�O����O��	������O��d�kl�-�T�#�~y5�Z%Wf�1o�4���My�cF���t����O疥ӵ���o���P��>�q��x����O:���7;��oßd�	ş8�I֟��K�8y%��3x̪%p���<c�6��O`˓��S�T�'^�'�P�%N4[��*6AN/>��`�vӦ�DKb���m�˟@��֟��ɾ��齟HkT.�?(�$�Jp)u&"�2�>�Ac��<)��?����?)���)�K�lxec�%�v�
6)�b��q�c$Ʀ���ӟ������¨�b˓�?��B4g_�EYUH4�6�@#&J)�h�Γ�?�W�\ii���?���?ـ��q����˭%2�T�Й��Cv
��Z	~6-�O8�d�On��O<��?����|ʐ��%��|�a/�;
h�ASB솧/���'
��'�S��*3O���i�OkL2�����GH���P

B%�v�'�Iǟ��ݟ q�'f�d�O�[�d� q>��!$
 ��Y��i�b�'?創N���`��h�$�OD�i��<( ��0ka��#u/>L�'���'%�ȓ��i�<��O]���6���5��J�9���ݴ��$8]��m؟���ϟt�ӧ�����A��ףwDH�+�D	xS)�'�i���'��DȚ'����<1���Դk�i���h�6l�2��M�Cd� :����'P��'����O�R�'���1e6L{tK�	$�)"e�V6O�>�l��O���|�M~2��^X���:~q�$rs�� D&=���i�B�'fBFI>+6M�O���O
�d�O��OR�����'R���hS�*�֙|r��yʟ.�D�O���f����
Ū%T�(�B^��.�oZ�p�"���M���?y���?�qP?u��#@��B"��Vo�dʅj5ע1�'R�X[�'����\��П��	��<���Һi�b�y ��>q�ɱ1�\#12M�޴�?Q���?a����SMy��'s��7 ���v�᲻�²��RyX��'���'�B�'3Y��#�U���ԯ �]�^]�TiՇL�F�0�	���D�O��$&�d�O����u����.!�9Sc�r�\����@�I m�'5B�')Y�p�����ħu��rA�Ս`�hP�%�r�&�b�iO�|b�'N�b�y�>�5Ä> 0���l$����"�����I韨�'Ȉ}��,?���O�Ɇ>B$�	;!nƕG�.i�&�!��'�X�	P30i��$��u�]�Bm�21�������;b�o�`y�*�6�|���'2�D�)?ѥ)Z>Y���n2st��x�b	ЦA��T
�
E՟(%�b?]��G*51
1#g�M�t!3F`�n�v������������?�(L<�8D�ȕ� {$@�6�Y�>�D ��i��r�'�ɧ�@�DR�WS�P��kP�9�>�Y�n�&z�l�ݟ�	ǟ|���N ���?����~�h�������?*�d��ULŝ�M;(O��d�-H!�\$>���ǟ��I���aJ&GR�"y��U N�Dv�ݴ�?�7	B3��O ��=������G�ZԴC� پ(�y`W_����AZʟ�'y��'5�S�C��׉Y"���7h~��;ȇx@f}�M<I���?yN>A��?�ɐXp�c �׏{��<� �9+O��������O��D�O��ҭ��4���fh܇H�褠!k ���Y�X�I՟�$�\�	՟�gjL��3l!r�t*��\�M3�!k�j���D�O|���Oʓ l�����$G�#bx:ɂ��ؙ�J%�'I�s�H7-�O��O���O�$�&#�O*�'��j������$ㆍv"XRٴ�?I���Ě�A���%>����?�j�$��x���rBߓMdl�`&DȻ�����?K���'�Q�/֎|I*̻��6%�oryB�[7z��7�}�4�'(�;?q@ɶ/}p��_�$��,S��J�%�'��m����i��6@h�W����(Sg,��EכG��kU7��O��$�O��Ua�⟰��k��Js��Y�l��C��-�F����M+nDU��(�P%;��=� �P��Uc6!iG`K�|�L���S
?jJI��dטq2�X`��I�)��5退��7�����S�I
z6)���4 ��\��䞆h����P�3*\���j �� @�>M 1t A"Ք� V��3g"h�K��];z���v9Pl�fE�*eT�q�"J�$��T*G�7hxQ2,�S��}	�Y�Q�Z4ۣ�3�Z`��ۘ^Lι��(@�(6���/�G���I�dO{��A*�P-tPvB"h�� ����݈p���'�2�'�D�b�'yB=��$A��1f��UũKQDT9��(p��,���9u�x�Y��,<Op�P@#�"e��D ��H ,:Ei^�QV�� I�na ���d̢k��#�����2�'��x��,��i�!Х��}��Q c�Iu�'z�@Q��]���m��'���MP�<�vF���Z���aJ$L���GS�<�G�i�X��@&^��M����?�/���J��9�����f@�O�0ȁ��3 f��D�O��d�+D <�@�?�� @��O����O�D4 ���!?_r��"���Jj����$@
N�D�x���>�U�1m�8xj��,J�y2ڵ�F��]�N�*����P;g��'ָ'j�����>�O�P�Z`�/w���9D�4R�"�O㌁X5�\8X\���n9�O<<%�����d��T��$fM���I'�ڐ��4�?q���	A��>���O��$ʐ&�H�aV�J���$)�"�o?� ѩf�z��2*C�d	�h�5E��T��wf��cDu���V'ڿ=�����Δ	' Qv
�^j}��I�(�4a c�	B� ܁��|�]���*���(���� ��6@�Z��OZ˟(�	E~�'���n,��TP!�5*��b �6�y��' �}ÊGx%��ą%H��!%�OZyGz�Oa�
ٝBd1°��Fy�`k����y��'5�����Q  B�'vR�'u��]ğP�Ik��
#�7H�zB�O� �|����4�`�ܻ4j0Q�?�=QB"ޤ6�0��!��>
��1`)�CB��s^���f�1�z��g�'��g"U� ��{��t~D��'��H���?)��Ĩ<I���7�h�#�TQ�e %�XX�<YG��	{��=�5��;!L��� F�;
ۑ�������'�6Y�'�d�j�{&�L�~Lp�C��7"��uZA��O���O��M:Q�~���O�����c�,J�w�dЯR�k�-��%�l������=�M�ϓ.�����.݀HB`�8���e��34�4|���g���tJ���'��́��?Y3�	�&v^����	Iک�D,T���T(\�ea#��S�̬�`C1D��Z@� 8�d��2� �F���o��yܴ��U��8�i�"�'��g�z�X2�Z�4Iʓ%�Р��Fʟ��I˟XhЋ ��<�O�xx���Jg���0�שHX�	ъ�$S��?�h�ㅋ>�����F�cuM=ʓU�����/�H��trV酇o�e�
%'�uHp"O0� �#����*��F�zw�a�W�'��O$咐�h�Ե��ΟS\��=On��Nۦ���T�OV2D1G�'$"�'��	�d��	$�1��Eۿ����Wz�N`�U�+lMڑeM�.�,������yW�֕UJ�Ļp(�F@��/ [���x����m�&vb)�Rƒ�a6��"h��ID��߅��Iˮ����!D8.���#�dJ(;����	���S��?��EJ��:��iǮk��Az�<�����ʬ�)ݛ^#���y�'�d"=ͧ�?1�]*n�@�I�,ϲ���nӵ�?1� ؜+$,L��?a��?������O��}���礝�!�x�X����r�z��$	Ǻ}"�aQ
�\� �ܟ
qFybI�AR6wf\x�2�ؖ�ʋsV`��c��G.=�g���j�|y�O\P6m܉L��8���>�d/�Y����g�!qz GYY?�ҥ�ԟtۓ_��b&e�{��)���&k�Zy����?	���C9���	��Ljw��+O����a�I 	��A�4^��`�$�2O7���ì�zZ}����?!���?I䀄$�?����H�vh�&	6(V¥�6T�Ԭ���C�j�)��Q�Oւu���!��ЍۦC'��h�4� 0�m1�$�	�����f�>vL�+2�ߞ:;PPy��"�� q���Oиo�	=�X�υ)[��]�j̷mT`C�ɻc�X!&���G�$�1r$��1�DC�I���� 2i<b�JW�IeV�ɶ�M�O>�"�Wa����'��Q>�Qw�2:`\ �㋃$>l�)#�S7O~0���8�I���� �)\�� ���_�XPܟ����t"�\��.-*�1�I/�ɣ�@�dVȱp�P5z�$�!NR PZ$�p���~�* 7�E�h"�`��.bqOt�#�'�n#}2�(�uP 7�
6F,��M�X�<	���w�p�䥜5H�F���V��IK<ϑ6�NA��54�
��+��<�B#�lh�&�'bW>���)�؟���ȟxQG�4�Rܺd��HՎ�J�a��&,�A�H�7c�m���?v~n� cџlc>�.طBij	��[>a�N)�,]�h��aRW ��!EZUo�q��uM�{����["[����Ͽ� DiڃdS��p5���šIê���IT�?H>��S�)�矔�!+�6�L�`Ā�#vf�hT�3D�lk�Q�F�t��,f�.m8��$�rؑ�����RQc�P�͈∘�C��ţ����x��"Z�v��D�����	ğl���u7��y�U���� �U��1�-U�k��Rl�vo��(V�_s��a��O���<�Gf\8y�ҥ֪K�A� m��5L�I2t��R���)����'s���j��=q�v81�O�ճA8C^>�!��X	v����O��;�%�Ox�d�O�Y���	Hy"�[���%��捳]��	y�Ŝ�y-\
G��#a�
�P��ЩB�G.<"=A�#�?�,OxL[g/���c(~�,���lł ����CaC��?����?��b`$����?��O�rFօ���k�eq���F3�p�S���I���� �}Ϡ"?�v%�}t2Ѓ�L� #l�,� ��	��BqE�#*B	J�D�89ņ����� 8x���Y���#<x����M3�F�lv�;�!	�Ecށ dƞj�<��e ?CfiC�,I-:h����b�<��匿1��;��N&]�%�<ᴳiF�'u��CUHgӘ���O:˧!��щ�DE�1Ìx�sT�\�$q�W�H�?I��?I5��M�Ψ��I��T��"%X`���S�Hjd!BC1j(e�-=�<���E�H|*(`��O*.J���kҝ
�d�wf�1��Atf�D��|R���׿��xR�	H�S�L�)*�p!�KށL��a����y��X��ip�e&6x�!KӧP��0>9�xr˟�	��	�O]65�Jc@��y"H�	7��7��O:���|j�	R�?a���?i��
#v6U���[P(a�� �^�t�CԠ^>�.���O*�&b>��ǌ&��ըg�H�<.~��u�G�Y�x�!	V�M�V��bF[0oΤ��)���#�c1�Dkc�d����!�!4����*��S��?9pEJ6"&�aI��63�:���&I�<�F��`D&h)!�I�R�ĩ�aXM�'��#=ͧ�?�FoWH	�M{Z(a���"g�$����?�Bz�z���?����?����4Ö$H�=��P���@�1I��!�&J�\%P��cL�'��1��C��IE�'�hq@[>q��#�m�5!"*I��-Z�(s��+Qañf�8������ɒ�
o^���N��&���%TL2�Ȟ�R�`!�߼@A��I E�4��P��	)=���Ё��KK�,��쇍d�C���p�Ê-����Q pRA
��4���O��'��Ϧ�8�x����K�fp�yE��͟��	��4��8kMv��	ɟ��'Ev���K*�rF�Ǫo=n)q/�*���
�n�3��=�`��� �X�RtG��%z���H_
�X��R��`��k�G��Q2�	�h%���
��A����I5�����A�t��0�"D�Dx�lţ'� �aR��"-t�5C?D�P�&h8Zц��3�ωI7�U ��q�|Xڴ��q�6�8��i���'6�S9P���5G��\��bѴw�e��&�ß���ßC%�\ϟ<�<�Oֲ���Q-%�:�Z��2?G8���d[G��?%���ۤE���{PH��"E~��9ʓN��5�I�H��a�v��#H�ҝ3��N�e���`�"O����Z�V�!AÕa>V���'�PO�h��b�:�R�`�48�|+�1OxH�׃����ٟ �O��*��'_��'B=H�ф *��a���">$ji�'��"�	A��R	|���D�K;ȡ����ϿC�D�1zc���D�4.|�	B�8Tj��4��"{'l��ĂpB���)C�ekh��wP���NM�s�e��藖$Ph��"�>���O� �!�+TE�B�C,Veƙs1"O�y�B�S
xÎ�3�O�'m���>�HO�i�O�1�<L1�`�A,bE(��F|@��IꟘ(�d"e�Ȥ������͟�Y\w��wt��%o6��d� �7߶AI���l���Y�O��=d��������#"�Ou��z��Q!�r`xc��$�8$�g��1% ��h �2�`���~R�i���	�E���$~1��֨���2� Ķdw�I�&�B���O��OF�d�O��/�|1�����,�h�k�!���?y�+Rq"�N8Qj� ��*� Ez�O�V�@�����McB�#v[>�ʴ�PI�J$����?����?��*�q���?i��I���"����1����&�����/O�4���@D��N�H� `*�k�<"?"K�l.��g�ʝy�ܙ�����k�� ү�S�J �g�Ӄ5��!��鐖��2�*�I~B�K��A����&�u�f5 ��Ag
�M#������O2���O���HÕS����ԧ�K�x}�ʓ��YHr�ɩjw������V�ԩ�(ΜB��i��I�#��t�Xw���'�哑` �����?P�y&��rw6諕��ߟT�I��ᎧZ��m���4SQ5�ƄE���=B�y`@��&1%$Q�����=x���a�� t윀v��g�"�N. �<K���0����:F �5q1��" �"�9�g�? ������v���Ab��})J�A"O�Ȃ�Հ ��F�Aj�����'�O���,�"�b���/β9���b;Oze:�����	ٟ|�O����'PR�'��f��n�>��g�J1H.��� �S'q��O�?MTd꓆��0�9O@�8�LH�klԬZ�dm��`��T�.�`���B��5$�1`E�Ǎsڬu2
&��ߥ�$h��?���&C�x�~XF*L��e�� �M#5�ir��O��`fn۾D
�,�"�X+��4PA1O��D�<+O��O���s�d)`����^���5'�/u"<Ia�i��7�O��n�������?��H��xq���m�T��&��d�	,1�ys���8�Iџ����uW�'��lӘRi����/2rltX�ac�t��	H ���`B��ɬ{$e)�O���<Qʒ�Z�0x𶡛�	i<%�co\<a�l�@ ]oʽ���6���pw����H���Rx��O�i���T�@��.�`�h�"�Oh���'ڈ����YL~X[Pb��(�ج
��s_!�D�S\�c!�6 򦈐���Z]J�Dz�O/�'\�E��$zӄX
�h�"uu�q �ɢq��Qe�O@���O��d�_X��D�O��38ف���@�K���J�}�`�R�	m����
�Rsf�`�V���O4�	�k̏F���!�ɸ!�Tx�*3^� ZC�]H8�<R���k�����b��>��w�%���� ��e�ح�t�%%	D�s���������y��;#���١���$��P����y���"�f
1��A&��$����y�iӤ�Or,Z� GӦa�	۟(�O�r��W�]�&�hRC ��L^P܀p�I�zR�'d��>#�;���0XhR¢˦z'�@�'mh���[�X��E� ��FlB�� =2��p�p	D+I�~yFP�bH��3����!���|v��f!ɦ!�p�;dc��)�� �1��O�tD�DCN7-�\K3�ЭjҚ����!�y"�C1�8Ys�_�J �T�^�0>���xBk³w˜�1��?2�`Tf���y���>�Z6�OR�d�|���ڜ�?y��?	� 21%li�`�$,!�ʂ`ǲXM|�2�������I��|�`S-��AmX���K΄~U��KJR����&[�1�Ȍ�׆1Jn�#nV�H`����'�O?��~G����ŀ��ĨS�ĉ�}�!���q!dOʅ�2h@�ɛ#��̂���?��r!C�a���϶{� c'ٟ�I�f��IO����	ß���0�u��yG"U.r�{S` i���W)�%�~�@Հ��>YrdWKߎ�� ҇4`P��h�{?���vx� �.@t�
H��%B<�n�������T��Ov���I;|8����?5b@���Ӊx88B�(U�L�b�`�0�As���P�6t����S Z�p�Zݴ2z��[DS�~@M�A��"���#���?����?adlʿ�?	����4D�9t���Z`�E�3�|���9�fp��,՝,b�� �̿8i8��`�*�D�6�a��L&���փGf�,Ѵk\�QU> ��#ӂ����� Śt��V��{L��\���O&�lZ�^�`��V�T�� ��ʹ[� B�ɲ4#��b��L���A�:\�C�	:+n~1�0�ѻ.5��s�IE�W�����MsO>�s
��F�'�rZ>�⩋�d���g�Dy����T������Id������,k$��rL�U�Ġwٟ�aԬސZ�PI�+�"�"��I�ޤ�Fj�J����֌�3Q8SXwȡJr�݅]�(�a)  D��ϰ4�6�I֗|ϰ�?	��S5�����?��8�)O<��C�6,l�l��'��-� )D��/����hO��^�	.)q��kD\�gaP`§�`C�v�\� U.�M����?�,�"�BWb�O���O
�	 aҩ""$�`�@D-Xu2�����7|�*��� �d�V%Z _�M0�O1��h�j����r��
U��r��Ч1����5͋b1�S�6u����
șZ�Z�I1�������V�Ab���/J�u}t=c�0o%�?�)���z��DV��p��\;B�D��E#D�p�6HH4�*#�����uC�?�w���Sן�5�0��fC���(�����8�Z���,�� �	�x�	��u���y�j[ F� )���,ʬ�.G"(�|��,��:8 �c'�*�����O�ʣ<��*�c5�̈��}Y��!t(�Y����5!�*u����
�L�B��'9�T	PkȦ ���O�p*q��P���ޱ"&$U%�Oh���'݌���Z�k��1��N���,����'"�y�Fݖ2����fN3�v����-��|BK>�����V⎝Y��h�W.?*�6oޥ[$2�'E��'Oy���'�R2��Q��oH�&4U�B� ��!'�}Z��]�I�����Cܵ�5�ؠnM�A:��?;��0�OC�m[�5+%"�S�޴
P��S�'
m����V # b����!

D��?�y
� n  �)�N.��3�֩Pה�"ODa1�Fg��yI�$ݘsxk$9O��nZ�ɠ�|q�4�?a�����lI��cTcN�N ����S3&�I�Bd�O��$�Oy�A�9+H{���y ��� ߨ�����;���F@v �ѓ��ZfQ��
v@��+vL!��fYA Du�$�� n6�pG�?� e�B���0쵡@�8�QY���M�	98�~��_Ȧ��	���O�T$¥\�-gX�@�F<�
 3��'|��'u�����"Jv�ٖ$	�X��5��,1����D�K≣7�� �d��B��m
�n�
�J�I�@I��ݴ�?������ű,� ���O��ğ�|ktI�E�N�d��7��(��%�t��IE�T�'�ߧJ�x����8�����w�p�C�����DЙ�I>e��Y��"2�*����J�I�a��]|��Tڣ*�/�� ��.�|��.&Lb�/d�p# 1y[�Г�b����J>E��?�6����۱pn�iH J�/Gpه�+ �` H�U��@0��!�XEx��=��|��#|��Np��2W��2\$:�
��?�-h9�Ř�,��͟ ��/�u���y��G��l���"n�yUK�yr��^:�q���`��y��޻i��|�@BK���%c��}Lh"��qa�`���@�ZHK�O2|�<�TM�%!���Sgj�%|��
h !�?a��N��?q��iu6ݟ����$�I�� �B�W�:�Nl2��:<92%1��/D�<�P�K<}��7��hk�@y�BN�M2�i*�'b*��B�O��ɓT�\�Xw����7咲-�`t���4e2�8�c�'n"�'o�h�9�B�'��)�/S����~��K#@ʱ�\0��c��8Q��̠$Jn��b�J�'���
��MWD��2AԔ8&+Ƣ�.;g�rF$�	p���p�O�U_:l#@!�0]%VQ�=�Ph���4ZE�2�.�H��Å���tR���+6A ��Du�d��3+��
���Mٸ5iD��!O��qkg`O�?�Z��ݴ��:�ֵQ��i�B�'F�S�yD��7D�Y�8"�Y�r�����ʟP����eLD�-��4�Mc~0����E��	D�7&ܘ+&O�� �0�i(o@Q���łH� *Gj�10c6�RI�3�u���&�B�5E��  �E�"c�ر`s�
&a��'�б@�����I�6d2�i�\40h��l!�D�5M��5s͂��,9��X�sb��G����&>��q�P`��zָa���E���To�����I^��m�"�'H2��&e��4`�	T�^F ԋ�g�	%��3��N�O�1�&@�0�1�OEҌ��;1�f� �ܔc$/W��F�R�Ŕ�J\��T�P�r���ao	�E(�15K�xuLEjH9��;2`����S'd�9�D�
�H���aQ�F�?QV�|���'���35��+g'�`!���V���'��]8���u��l��y� �0��D����D�'ʭ��
ۼ5�(�!U�ϊjؐ��q�'���\m��'��'��o�I�i��h�D�N���u�^ڎ=�t�d*ll�U�3XG|��s�.z���6�(O�dr�.R�u�fAGm��o׶D�"�F�bu���C��](l�:{E����9$k��[��	~Xd��g'P�/P�Z'h�9=�I?9�r�DTz؞��6	g�l}ҒN�v�����-D�D�Tl�;:�P1��2 ��P�b���HO�i#ړr<x �Wm>H)�'K�$���ȓ8�H��ݱ^V���`�\/Y�ȓP��M�aJ�]!�8Q��+�@���b0��b�֊>�b�s�C\3bz�ȓ����&WD"\���^8Qrbt�ȓy��dB�{���(���oO����_(T��mI�8�� j��_�>��t��L�� ��	S�
||���A	��$Y����(���{X��Y�m�g/ȓB
�
UK��<�����#�x�ȓd�<I��@��c��l?P��ȓ*�l`��&�9�Z1 �E3����tE����T�Dh:ؓ5$�2]�l���gYN�:A�J�'��X�Ƈ�|����/z���%HB=.pP�Jt��P�~��ȓ3K&��1j��?��-Ze��vq��
����E�08)��L4x)\U����Upu(S�0A�u��%�1l������Q1����{���<p�r	�ȓ'�`ja�KoNd�'d�,$��� ��(�*t�x�1a�y���ȓ,I|�r���a`ډS$�UHa���S�? ́�� hq��F�D�4�#�"O����O3v�[R��&|���"O�RJ�P/f� Pτ�K�"I�5"O���ƧŖc��;!�\8��e"On��\�위Sv�,�"O��ۤ�ʿ4;�2VjL�T���i�"ODAab:/&�����'#��=z"O���2`�).� z�D�.^���"Of�r��|��Ԣt���3bZ�1B"Oĥ���k�"䇭6
�)aE�|!�䏆~��lK��>L ���Dp!��~��`�Ӂ�=�()p����MW!�$M���A�'�7&vVP�@��2.�!�Ă�8�@e3a��&y��Rk)��|BhZ�$,7M]<8���rR��+h�nE`B]�KD���Eg��<���'*��q&\�t��2�]l�Z����@+?AT�#�\�h��)��'X���n�)����H,%
s/ѳ����"O�l1$I��+��U�_�|M��b�)Ѷ����u~���>ӛ�O�T�������w2h����4�&�6���Mt �I�S���F�3w䍹�E�V����"�� Gθ[�TBteE/<�P��%��H��3�� c���s�P�ƍɦ\"��&��	93f-\���&r���'�ؐa��\�x�楃UEH=!�M�f�9f)Ȥ��a.lOǌ2pp4�\%@�%+�_���>钤�?<�Z����%$�"-F<6Nq��&$�ĥ���0)��`�u��?�0 !&&R��@1��q��8�H��H}���S`@/TsJ-� Ј'��Iz�˧��!Pt$B����i���$mاK��E��R'�.5��O��2/\�X�H\h���!��p���L�T*��S�	����XY�d����Bj8��ԉޚM��0��^�M�����HO��c�^:oz���;�4uya�N>q���OA	.j�v���?�B�O'�����Q8~�����(K�����#um��a���j(�q���ߍ`@I�iI ��AJ+0������(F��`�`%��'Ѻ� $Ķ ��1d
�;/��y�(�;����D3O�zV����1 2�B3����`�aM�2!,M��:A�E�������t��'��6]>����&G�j����M3��	 1 �`�H��������Z~"H�"�8��'[�u�44 5�M�g�I4 ��P���2ӆ<j�E�ܴ@#�T�B�����O�|F|�MC$o�ވ��
� psp��O]4E�2�8<�P���Gɧ�'��H�`�<
�񱅮@3�<"f�Ry�0�çH	?��>��	��� ��}r�eH.aޠ@qL<���۰�y�2����O9�x��Q! _�X�P/U4*�p	ȀI��nM6�*���R�Q���!(�4����7s�*%����(�x�jџ�|�6�TR?F��$T���K�1'��S�	_4%<
m ��_(6���'����7�2�x�O�I�|l�O�����?҆I`�kS�F���I<g��R����'Ѩ�а�]�*�p�#Nɦ�q�(�]�f��IK�����1����9�6CI��ص�P-xH@TA
�S�h1��i>=�'b����+����'f��\�l�$(d�����?�6�ʱ�'���:}�,�WC�����Ԕ�'�}#d)�OFaY�k�EܧPc0��3��0xÌa����L�\^��P���#�l��
�D%�q�2ΐ"&
I����1?�8�Zrf=�6���HN��O�l�I	Q��;��έb���3�4Umj��3+,�����g��u�~p�'�aC����}[��A�&��`�o&}❟���GVI�h�h�=aSڙk�-`�p���",-��L�!`Z3���5��z�=1q�Ċr�X��&�F�]a��ò	�?S�H�*���-⛶�ik�m ��xR+k�aZ�a�_�.7M%q��a�� ҀWD�-z���UdTP�e\� ��d����!���{P��$�4�֡�?0�$��+�J:��} f�2�S7����yvZI��MZ�*�h�H�����O4ɱ�JJ?.R�Ts@�T�7x����i1�}ÃKW�MB�q�$'3�^�;���%��u�&�6?)���á��at8�@��92��=���i�P ��CE	��
5�C�_rb�)O$*�#�$O-~ȋ�T�@m��i�O�ͺ���q���
`�`��x!�i?���"O!=��@��1o�|ՙ񫎡�HO<��Ѯ��>-�yB�Ԡ,���g��^m�)�ת�����%��N��E���.;�N�h��H��X��@�,C�6$s�UL�����&�j����$Ƽ��	7�v�9�l¸P;��Bt��G�"! =+��^����|j��F g\�T ��X�D Ҥ+Ә& �,�v�I(@�F��#
��5�lѕĪ6M�4_�H������!�	��'���oq6��O��l��!�D�SBFD�PI�Hp�p�	�ڴ5�h��DۊU�2Qrvi&K��X�'ZV������[0X���ºJ�4]Z����;*P0��!R��X�voS%
&�჆�$�� ��0�����F`�Ad���y&t��e/ק>�e�>|Gz���\?���O��?��#�4O:ʤ�$(��<!ƀ�I��H�\��azB�}�� m�%����B�d)H7O�;F�|b�>ٴOXc�"G�زC�a� �B�� x; a!WO���"?Y �h����Z��=���ЦqZ�F�=A��XIT,��3��11ﻟ��{�aM:%v��f-A�D�Y�C�Ԝ�yr�� ஐ�4�jp
uڷ����d¨3¨�+�a�
^�V��+�k�1OV�I�h�����!ƫ �����ҋ Q(�oZ]<:�z�W�T�Px(zӢ�D}��F�kS��$$�E �$���Z	�l��2��)��Y�Ӽ�@o�>8y�	ݛl/,�/ W(<�������we��$Z~$3~���d��kC�%��+0` ��q$T�F��Y�2O�wU�5R�k�i�������%kC�uzS-O%?p����/���҄#���z5$C9��я�0,��IZr�2��!�f@�tL�/�#<I4ϗ�.H��&H�"�h�@OY�<��Ī.�(��Ot��I0ǇQ�'�|0Gh����t��,�7����G!3f(K�&]��0>Y�#�&<iR�۵JL,�IBܖE���"d��sx��`�Wn�v}��`Q�2g�p�a�r؟�S�
ڏlW2(k���|`b�X�}x���
ӓ=�0�$�|I�m��II#�u��l@<&Ǵ�b��0C�.qG~��7&��0;��Vτ(q�!�M��CF�[WBQ3s�2l�W�y�'�Ȍ	� �M#Ԭ)����6���)�O�ѱ���a9�bǁAِ�bX����۹W�Ȃ� w�Y�f�6����0A�db؁�n]�xb|��'K+SH�C�(�=i�D��/�g�ĩvG�5;�M��@3�0�SAI@�*��lR�K�4�yb#�S�=/����*2^�K��)ul���v�''԰{��)R8��aG�M�+��2mDy�<)�O<M�<Eb�b�N4�����ʥR�8SѪ=:Dy��	!w6�Y�P�� '�ZԢ�G�O��$^@�VAҕ'�6'#@���
�5�� �J�	�+�t�i�':���l�TV�B�44.T2h�&D�).}�hHv �Q?)�ICa�Np�CNS�Cx�0���>�S��
��ps�A?ldX�)>_�~���W�4�1�NF�e2���'O�������kZȝ�T!��{Lmk�k�+؊ٹ��ܹ�I���=��~�Ȝ���2����.��@P�3'	�2Z�<�!�`+Ry O d�(
�%��H�-�.P�&�'��I;�M���a�@��iJ�j� �?�DI��|�7ɘ�	c��;B���uV�����t��HZc-غI�PM�3��@�h	���K.*�v�"��G�������m^�7�Ȏ�~�"�/ Mhʧ]1�s�8��3`U���X�o���s'9��;d���K�ҋzN�TK2H؎#�������ńsٴ��d�E.lRje��Ԑl\M:�M�+�Z��"�F6�Mҟў���� �
9�F%��_��P���N�!ϨP%���*Ԣ���F���9���O��'%�L `�Ȓ�=L��`b٠:��S� ,؆�����u�ݷ���p֊P��9ÃFל�|�$�M-�`�
qAn��鬻è�4Zc�bxa�SKʐN�>����'~��7 �҆u��I��3�	@�1qtMSp �=O�1C7L�,S $O�E��� 4C4�0��sӔ��e%G(r�X;i����u�x���6R�k�〒��� �%��O��ٗ��F��P�CV� ��xv���M��˘�]jv�h�<BO�3ғ~T�0���]�l��2�_"{z���I�.S΀x�����n��$ ��N>9	^3>|l���A7 J�`��ʃ�p`��3��7�Ok̟!Az�� �E�^\�A3ԦQ�y���/ɾJ�^E���������]C��֖'?��)w�VbІ���GJ3�p<�2�̹و@6�>iM������P�Z����R�|����@�LF�!KѢ�*;�,����i����4$�Z�Pa�����<a�aV=i�Ȱ�B.�bs��a��i~2�L8|E�e��d�+�8ͨ#�9�ؤ��lo��'S�|qj0aY;�\UY�61��1����������OZa'PzF{"�Z�9'쒓��%�:�2���2B���w��y9�Y欒-7Up�Iy}�''|��^w��I$X��tpV+P<Ӳy��NF��D@�%E^''5a|Zc0��p���%*tT��"�֒u�ʤn6@��<Is�چ*����;4�6AK�"�"�qh)�3&��m1d�'��S��S�ќ0C�g{�6@I�*��i�t]�����*Ƙ)���&$�)�VM�g�RIl�"��u%��R5�\�G5����$z��[�� �6g=�5�'���	�-NzMi�8O2x��{�c[�><��G^j.�\pA�8e��p�o�䄣���%���Q"��~��D|B�΄R�\l[d�=���cE���<���)D��z�J�p�e�I���iʆ�T��DY0�	�0Y�h�塏�,H4"�Ӽ��˪m�y�po�j����:��D��HwF	���p�rx[92�(�LW�`�����0<��N��$::�b4X���eT!��=K�$�T6u:eHȭ}iF"?Is�Ig	`d����	�n�I7*���Y��;L-|H1��*8 ��W�4?	�jP���@uW�`h�xR��E���3E&� x��Y4�[�|,��0�ġ���B݂9]2�a���!f��� m ����4ީg�N!�兌�R|�� ���@�����s��x�7O����t�����XEB	�Hn8L Q,�!7Z�Z�H�Z�{�K�;��`9a I?##} aH�<�'�S������Ӻo��Q>�2�
�l�� ��h��߶6��A�Æ�Y�0�VO��j�
F�%�:�E�/cK�4���E`e%��kk�9Y��7mY��h�9���r̓P���T�H�N'��@�
 |�̆�Ib	:�"�4"ԛƏٌ�McSMI0�^XyeF]Uy���YU�Eϓ��4n<�p=���sGp!���ɤxyK0	Yi�<ٗc�:}�%c'H���pS�G�e�<V�W'$�y��"dzYC��M�<	���w���P׭]�N��#��"T�l�$��c��qh���2�:���!/D��$m
A��S �,R�*0���)D�<��Y-�d�`!��3C�Uc�(D� �7%-?P�L��Đ-5�"���%D���1�zVlP'�T���dg.D��*dnY��`#nJ�
����)D�L��ԑ	Xzar%�Tr�$�J��,D�| �a�:_|���B2m�V=P�*Oz=��^�`6nTA1�4+�0�pc"O8}��M�Nˌ1�ǉ�z�zTX�"O��$��A�1Sg�͡FD��@�"O���C��8�񒎜r����"O]y�*�/@��}��9��y��"O��a�X�O,r��
�R|���"OK	�~�d}��&;5\u�b'8�y"�Y�1~�i���V ,��$�d��y�i�8v�HP���� ��Q����3�yr�F�R]��Y�J�8�qb���y"lՋ#t��cM�3��	ub��y�*G>G舤���@�����yO8	�8��&��>���� ��y�@՟5�LM��Ē!}��ȃ���y�Η�v�PЪ������p��yb�M=$�fܚ��̢%�bp��!�y�%�(O0�B&)��T}����yR�t�a�@��|�꨸0���yB�ԁJ-j�-�qR8�dX7�yBc�?�B�j5��Lh����y$��<=q-�"E��xgR+�y� 
�vuF��%jgZ�x#��հ�y�>#�s��$[v��X�,U �y���g�4q"D�,K��ٲ��;�yk�)9�`��H+E�@Z�7�y2��4}������5D;���y�e�0cS�Q�E�7�t-�4%X�y ��6k�!hb�E�#?Q��R&�y"�]�x�,�(�$V� ���I߶�y�
&=+�� M�u`��3���Py��!M��Y�&�ˉj�
$�7�I�<ǠLhҍiQ@W �pP2'c�F�<�bM�`/\��:Z,H�SL�<y��'Kv��Q�з����M�G�<yS�iV�:�c�7P.�b���D�<�fƂ:%�0�ȱ 7v�K��a��C�I�OW()/�&��*�ͥ=�B䉌|'m{�%�RY��̌ |�ZB�	h��� K
�<>��&eJ0
RB�	�\�NL�c
ʚD8����Ȧr�8B��7'��]8d�Z�i���aVGĂYu0B��d^�[1�ƭ��j I�t�B�ɾ^��HPE��$������=;�B䉔KÄ�
&��<0~|���/8^B�ɾOԸ�!D,"v4��D�?4�C��o������ztܹ�JŢh�C�ɴ;?�Ȉ�IU�4x�"�&�B��22��T���3h���O�8J8B�)� ��h��S�K�P�0���Z��D0�"OF��
r��=
�/H)K���au"O�D�cO��� #e�_����6"Opغ!	��E��'�f!�0"Of��%b�
��H�%i�,;�"OHh�E�,�����I�h�X�"Oށ��,������h�/	�:� "O`=0Eŏ(np���1g̬9�(��"O�lxF�5!P6�鵆�'��ʅ"O6�9��ȵ�X�'OV)gP�i�"O� ;D%�5���6� fPѡU"O�Yc���*��s��I�BSPya"O(�T�[�<@��]�Q4��2"OZ(q�)#�D�LO��0�	7"O���BM^�5P��4]��]Q�"O��B�Ϗ��02�k�G�>�!�"Oz#Phǋ���	�j����!��"OxEI��{������a�ft:�"Oȥˇ�Y�g�Dq3�T�<�
q�U"O�`�c���z24A �xl���"Oz��#��tk.�p���<�!�"O4��ou���a�u��"O���U�*N�©!F#O!>��	�"O�T�G�	!k�@l�AaS"QqCD"O�|�p�W��
����m<����'��I:;������T�%>����X n7M?�\�!@�a0��	��<E@��4D�L��$�$�ʨ+��ę^�H���2���I"z���вg[(�r�$��~�C䉥-�8R1oM;�hkg��%N�<i��T>���J�S� 1��Gʸpm<�ba8D�$I����J��G�K�\�yP�5D�0��H�;Q0����E�b� S�(D�px�M�f� �	Ł
��5�0D��x4��L_�+�bO*\5h#.D�d�L�q'�u
 ���s�҉,D���� 9}(X�%ȝ��8��,D�|�AC��M�@�6Hٶ7�T9�Wj.��}����<�<e��	�=&�E�&��y2j�R�}+ə�"���qf�!�y��� y(�Q�'��/��ȕOX5�y�.����7��]r�#��֡�y�)I�~ɚ���ܿK+��sz�B�	�� �hȮ �n�8���1��(Dy���TȆ1#�~|c��
��q��'\V���!���L�6�V�c���$�p�>���~"�	�1+��zW+�Mh�5���:�yB��',�1��/���2B
شG��=E��9-(�K�J.+#�����X��ͅ�	Lܓ��@��j�<Hz6�� و��Oxy�����u�lz�]�xb��C,��er!�d�
JNP���sv>�{�k���j�=E��'l�<BBKN#7ˤ�0C��c�E��'��QR�?o�2m]^��li�':6��cU�\��i�h�OU���
�'>22��=`�ݩ$�ޗL��dS
�'��0 tfӖNk�j��ǜI"�3�{��)�	�U�&�A��x�TIS���0I!�D �~��p�%-���A&�ۛ6!��E�C�I�1�M�)bx�hS�&aaz2�DȦ!�8�3�LR�Bb�ᏑCQ�v
O()G@�5S,������1fH���T�dG{��i3`�:��"��"�d��H.!���O�I��E� hY`��VMF<Iu"O� ���O0=������=k�"O6�:��D*p�Zl���:��h"O���l�2,�R����H�= �"O�I�	�\�� ��3`��"OH�Q���<�xZ!Ɛ1Q|��b�x��)�ӷ$�P�(E�5E���R%�w":C�ɧV��ʐ(�`{�8�'G�|%C�I�zhWH=D �QdX�]-��C"Op�z1c��-֢h��&#��"O�PrVF쩳�޵n"X��$3�	Y�O�4��Z�|�lD�E�s
5�'�H��Gӫ:C���2a�*$���'�a�A�~56@����?�hp���y�ED0*�S�e�"�6)Åe����'����""�eɦ��� ^A��+��IZ!��(?�.�æ^�g}���?�!�D$*Ĩ�s��-��0��KQ�؄剃!�b,� �؋H�&d�PF��^�B�	�]�s̫r������X��F{J~�F��c��Dӧ<+����sX�8��O<�c�!����	��T�j��|��IMX�$�6��WnRҷ[�`3}P�'D���R	E*Ű2HN�#�����0D����n�)OSԩ���M� ��e�'��x�1F��%c2�Q�o�������d �L��D���Iǁ�E$,@��xS��	SoGX�@q�6HW>�� �ȓ�Z�h��
,u	>I4� � ��ȓ=�j=��I#	� ��%p4ՅȓpR,iH$�ɂ/qĜH��<&d�ȓ��h�1��g z%���$3�vD�ȓV�Ċ�@0�4� ��&<r`%��fj���k'{���V�.)�l��ȓ+��1��8�s$D
+a�ẊȓT�	����]bhؓW�;Ʀ�ȓ6
8� Ѝ�.��[A-�	z@���U����i� 1�T�ކ=^̡��G��8�b.S-M
�"�-�:�hІȓ<��IX���
=�pҁJ]�6��� 8Dub�I۱ s������uXj��ȓN�\�$�2-�<�iv���I������;T+ճ|���1UcLi�8�ȓ��I� N�4��IY'�Ra�y�>yK<���i��(�V��CU�F|ꢅ�m�!�DZ�O�H�i��I�0�p�C���k��'ўb?q�W䚇���D�
c?H��`=D����Ǚ�u�l1�	�-(�j��>D�@���X�KC���fH��h �k>D��Ҋ��N�r�k��R�l2��y��;D�Ш1 �?h e7
PM<��a$9D�\��,�U�'�O7ZI2���"D�ID-@�V��&h4Y,=1ti;D�0x6�Ӷc�1�· )��@�g:D���L![�tT	���51P�Q�#D�YC$ڗ\u,�+��ʶUK��a�"D�T`3��2f��h2�\\���(;D����Ȟ�W\�p�B��.�G�7D��P`�T�l��A`]�q�0%�2D�x0gdG�k�}`2F�8bvL��L&��Q������ܭ��/"`�	b�V�\B����13 GC�@P���;|,"=)��T?]"�iѨ>��H0�ۯ+�E�&&D� ��G^hX:g���H��K6D����^u�r,[���.f��|���4D�� � �$-AZJ�V㋇�4�	"ORX��
��Ly2�7�P��D"Oޕ3 � I�Q蓦Z����Zc"O0�B��_W�tI0��ynTS1"O��$ɑ3g��{�CR�@��g"O�p����5y�����b�M�@�JgH<��Eܳ*i#�"� a����GM`�<��H�=9l�s!��	��$vA_�<1�,�[�>�I#i�6�J�B#nZ�<����6~�*�"�k\1l��:�-�@�<�S� cd�b -�#�����Hy�<�G 9q�>}��"� �t�<y��Y2k�Yb�?Ȃ�zI_X�<ɱ��wom�ӎ^�[�8��T�<Y�f����@He��$n1�%"��N�<�u!� )J�*�㇡���&�M�<Q��K�Aτh���F#x��0��+�_�<�����?��wA�qh��X�<�3%׷54�J��E��Px��X�<	�b��}#`�L�t�ࣃ��I�<A�Q�`Z$����.��(Ȇ��B�<Ѵ��<�<���1y0��k�`�T�<�p
ؘ6֘��vbӯZ�"9YU��S�<ɲ&%e�0�c󩟁'�ڴz3��y�<y�  9��h6GO>;���jD%�[�<��Ü/oj�q�&d��G
X]JD�[U�<a�M�L��!@$�i�R��� O�<��EM�X�x
�G�a0��'��r�<i�I�`�����IT�GV����T�<�����u\�z���>:gb�0a��X�<�1��m&��"�&%0%�⫚Q�<9��������
e'L,c���K�<�c��-����:������S�<����9��4�W��� ,DBpcQ�<I(Ϳ<r��EN�}�� ���Dg�<��ń&��T�pd�21u����l�z�<�֪]�!���r%�]�T� 𰄃�M�<i�j>!BZt�1aǭEӺi�veH�<�E�uHtm2%)�.[Xp��\C�<W���j�����)����д"IK�<q�N�8�v�pJ��D�9�EME�<1�i�A�L �g@�;r��Ay�<��T�l��bI�k��1T�Ox�<qS,V<����g��&cB�i�n�o�<9PM�2�����a>��l	e�j�<�t�
��B0�r��
���b�<g�S�6aH��*3�(��^�<Y��(4�ʽQ�J'I�����\�<�bީsц�`a*êW�F�C���V�<�Gʞ$h�
5�&`�?#
��s�S�<Q�T�]�X ��+s��ӐK�T�<�U��i��8!DD�?�1�P�<!�Ë�;�@��Ā���c��x�<���+��<JdX7=��5�wÏq�<镂ڲT�a�$��*���H,PD�<�FGaS��X�
ZtЉ#dA�<�wb��WNI;�?�&��}�<A�*^{��:t�ٷA�AY���w�<qo�p
���dʎ;�H���Mt�<��J�1���/V�	�D�Ӱ#�s�<�2O��KCF��F� 4��4�iF�<�%G�3���B�V��\Hpk@I�<I��1.ƈJS�X�:�D,���Vi�<��%�z���A0�r�N�o�O�<� ����1R�L$��N��q"O�|a�o@�P�y0��.1l�%Z3"O�P�3٘B C��+{
��#"O������*,)%`*��)�G"Oҹ�0
$�����H��"O��xq�M�h'z�3�hz<�� �"O2�v�	����I�~7<E!7"O���3�)T�j��nG� �&9��"O�Jc:I���S���l�~p�"O�-�0@��k`�s�� ��q:�"O��z�i���a00�ϲJ���"O���S���lM�KL�N l�H�'*V-�V��_=-�U�D��8)8�'i�ظ��՜(q�A;e�wzD���'�tl0�bR�pWft"5I�{ 0��'�Z��������k�x�)	�'���Pj��m�h�D�E	p���q�'��8��Ŝ�L�>���ԹPF��'��[��@���=���O"9��`�'"13ǐ"[����ga��{�p 	�'��,�]�b��hK,�>t�FA8�'���{�Qa�x8ƀǸp���	�'��b5I�&n��]˕�m�	�	�'�34j�R6�:5��XH"-8�'S4t�1$�C&tT0�Ҝ�H��'��M�!.�b��1�boM�o[���'$�]�4��#�ʑaX4��p
�'جX�W���s�⍯$΀�x�'��:T�܌H,���W(p$!�'������ܗd���9M
��f�B�'.���_(�u1�Oҍ|c| ��'Z0)�ۖ��j��=A.��	�'vB���w9�0��:�V`p	�'�P͋�`L�'�2�Ж#�$h�B��	�'��Y�@o�sܲ\�f/j�B|Q
�']��8��X;j�tx���j晸	�'ڤ�� oX*4�rIr��8_`���'���A@��3BO��ƧQ��a�'��zPAD9'��9uB �wh��'��1!��]�M���Q,U{���9�'	0p��®l	�A�%�H�8R�'��t�u�~��1�ȷ�U[�'�QX����"��E�G�H)?�b���*�4Aa2b���@��O�<E$l�ȓЇ��'Z�����\k3���ȓ]4��6L��;X|kRIE�4����9l���ᕌD-@S`�Aw�ą�
a�1�'n�(�t�BS�M�e�T��6�X�i�*y3�B+��D��u��x���	;G��x��kJ�(��o���c7��2\	`�v��6[�~���xv�2�D]6uiJ`�Mt���ȓ,�с�CB�X-Lԑ'n����ȓu�l����ci����φS�܆���0l�D�H��Df��
\T�ȓL@p�)�RHEC��||n�ȓtR��΃�M��$ Աgg&,��5ȡ�q,�.�x9�eG�@�����`�F�i���P�X��&$xҘ��Ek���Y���d�I�=C��ȓg���0lB�FPR���*d��ل�'�H��w�Q_՘�90'T%6��=�ȓq�	8�G���qg� 5t�����}���h&�� r���y����S�? ����`H�u͸���J8;kz�2�"O$n7(�Tx����ZdZ�s"O�j�O��dBAX�Z.���"O|}�FN@� Z|�7�ԣTu���$"Ol�C��|k�e����t�}��"O�A�F���G��dB�\�K}X�2"Oū ��&4uʹS��.uމ�2"O(зȖ8���H���0IU|�;g"O0� d�6$��cs>uHX�"OL�BG�BYJt�t]��%C�"O��[��̺"34���F���"O9�w�ėV��p	e#��,iV��"O�y+��L�\Ppc��P��B"Ov�P6���/���
�GNED��"O���$���%v��T�Ĉ,�0�K"O��
EGS!g6���`D_ �* �"O$�I_86HfZׂ�'�(,��"O��R�+]�+�Xѳ�c+�##"O�ɨ�%&9&��2��&�x"O.9���$=�҉�A�E"y"� *"O���2� 7��kF/Շ!o"O��x� ͷcF.�Y�-���P��|�<��d�<T�\Q`��4Zh��"�G�<a���'^( H��V�tr���k�z�<Qca��h������#~��1)Ǐu�<�C�r[�(��')',��W��\�<1�M(Ya
95菦Xyh5nEM�<!t.T  dl:Ŋ��>�9��HK�<����OV��$D�q����-�_�<)��Q�f��"Ug�=}N��VS�<��Qi�0%�)Q�?=��fěL�<�t��/��I`��9`J�S��F�<�u�Q,]���Q%ª5
�'�{�<9$���� ��L$Xi���/Co�<�ˏ48������נp�~���C�Q�<���ذdk@�B���a�`<���J�<I磒����{ aɅw���x��q�<�+�l�����H���h�i�<	qKF���%�"I(cI3D����*��<x�����������k�<�q����%���������k�<���йh�($k�C d���
�o�c�<�����[-�<i�K�/WD�<93#ءzSDP2D�� D�a��%\g�<i֮M�)�@���X�2ܴV��!�d_-p� �h�N�-���b���Is!�Ɖ#b� �*P�ԣ�Ǎ�Cf!�$
��4@3��=�Ѐ�a\��!��?�|0�L�6��S���k�!�D�	>e�}`C�K�>t�;� �z�!򄏹b̴�b Ę��&ݱ�&'�!�Ƨ^{~�H�bP:���""U!��{`�m[)U��u��e!���j�mX"@{\1w��H!��LI�x�2%�P�]`j0Ԁۦ!!�DE?���P�i�5�6`4�!�	��t�b�P`�殅�!���ŒM�����>�j����,�!�d��e�f�rd��P��`�֬�J�!��G+�dq� �X�P�L!sY<e��'�n������1X��z�Ç�L�uZ�'X
sg�Z�#����d��=>�J�c�'�4�h��o"��$�׼c�^�`�'��@&3~��h�WR������ �(9��T
��ZO�^�n@ �"O���M,p���?&耀�"O�9��l�%x�1�2)͏ VT�!"O�|�J�9{��Ee'��w�R}(S"O01��_4p,b�:DU0!�E"O8�1u�֙~:���Ī_�t�B�r"O�����U�8,A�(^#N�e�q"Oh�����R���x"'S0"b�"OFQ�
�u�R���/jR1P$"O��1��^�.�+�o�B��{�"O���6g��]k$�4�E�Q׸���"O���B��)��J��Nq�����"O$4d�A7&���ӳg��+��#V"O��20ԵgJ@G[�-���'"OM�tȜ�k�h5���Z+ yP�xW"OV�æØ?J��<`�a\q�	��"O�0QA�}F�p��"�DaԈ+`"O����î(:	J��/Z�y�6"O�e�C��TR�A��5e��0`"O�R#�C�g�D�i�(OK���c"O�%�R���W|����0,b��"O�Ez����D��=���r\EJg"O�A��o��GG@<�	Z�<铢�-p�Z�b3*܆-U� p@�{�<)Qf������?Z�\L��)Qu�<!�T�����U�A#W�N90e�u�<1A.L�7����(��I�6�[�˔q�<�P�]:�
� ��D�H�(=���Xl�<q@�Ӭ1�Ph�E"P+vrȋ@$V@�<1w��7�,)aa��z	z4�l�q�<1��\-~2�m)��>4ih`��q�<����&;�mZ7o�/P|�U�G�<��k
�VV� 32�^�=�rhq�(�@�<Y@��$�HR����J��Ul|�<�B�Z�:�TA)��� 2�\��W�u�<	���!�y�Ŏ�:v_�@���K�<مl�$U4
�B�5Wx TAEAE�<i`EKU����#X�3x���Ǫ�B�<9��e�I��	'@! ���UZ�<Q���rТ��g��@�4)��^V�<i����:`��>� Q�P~�<�Y �Xs�:J�� hHu�<Y5C=uH�y�ɕ5��34K�o�<9���Y�E��9�"�cp��e�<�bjH���QH$Oߗ{���^�<�	��%h��P�1Z�5VnCtW!��-3P͚Чsg1(d̈�S=!�DO�m��E@u琻����aU>!�DU���\PT�6�l]砊{�!�DbKƕ*s��2;�.Ew@�`�!�^�s�$�@ B��3#n4�"�:eѡ����(9��@������yR/�FϠ�bu韨���Js���y��_�`�q���-�ʁ����yb���{���i�/��oq\ɑ2&,�yB+cS,�����U��B�'J��yB-C�C�,���E8O`<	�%Y�y�K��j�(i��WtH��t�<�y� T6�����ꊳ|f�\�S�5�yB���-�$�F�tW��R�<�y��V;� ԙc#^�g�"]c�ύ��y��V�kX6��4�P!]?0�I�(B�y�MN';� �����J48����ۡ�y�Ávb���'�&Ho֩"�%�.�y
� �=�3?�dYá��tWL�z�"O�,B5(ݡY��"�Γ�\P���"O�1a��+;!&� ���
!f�p"O�Pȅ�N�`r9�+��d���"O�S��\����z4ᖻ#hb���"O�#�Hɦ8����@O�����e"ORdJB�˳QG�����>S���"O*���� ���*֮^B�~u"O�҇$NɾQ�׌�4i��iy�"Oⴺ��1&*Ap���W4��Z�"O�����	�S�&(�BI&l�%"O,��`k�rWƙ�S��-��"O�m�!W�L�A�%�F�L�H"O��g�'�@4�*�T%�)�v"O��F���zݳ�+I"�0
$"O��ŉ�r.��TЂ!F���"Ol���.bؔ��!!�F��"O�*3,�}*�x�<WX�h"OvI�E��[�u�tK�FP!"O����ꉘISڽҵ�;�Ѐ�$"O�ų&)��3xn!�-J2k��a[�"OJu���[�4Y�'��|�m�"Oذ��܄EPm��%ʚ����"O�% ��2 2�y��ÿv0�R�"O��a��'+�A��2�|�+U"OF�	�A��e�^�b�N����+�"Od`S��t%�|���w�`)2"O�d�'d����'gk�ة5"O��0A�L�`���P��ur�ؐs"O쭲&_*j�T��ߖM�8��"On�6�J_��S��"J�xDQ�"O���5gP�5������	�:܀A"O\�*M�YDlB ͉J��mq�"O(��&���d� ������D"O�a�0>�����5���"O��g��gB4 ��	Ӯ2��`��"O�$�'қo;�A�B�WI���"O�-ꖁ�+<"�b@h�:�h�"OzMR&��9 �pِL|ب�"On�#S�?k�	�'FОW`%)�"Oxih$j�/�B���A��,t)2"O&���+�.=M B��<.ۘ�x�"Oz��o�kT<Q��M�	�y��"Oġ�5M�4A	1���N�� h�"O�e���/T��M����C:��9�"O(��c<v��W��4%}V���"O$k7� (�m�,W/,��E"Oh�:��S$�da��B��R��"O���]"/!��8��P��m��"O���N��G�	Hw�=_��
�"O�Uq��98$eF�=���V"O^pQ�!Cv�f�$.�� ��	��"O�Ge�LY�k�&�~�)�"O��h�	�#u\v5[�	A�=�:�	"O�P�t-��#����H��׈��u"ONy8��u�tQ�s��i�:mb�"O4�����iMt�� hQ�t�`��"O,`�3&L)�!2��v���D"O@��%x�M����Wh���A��v�<�!!�+_��8cDR�UI��*���j�<	`��c�abp*Y�$5�Q����O�<A�
K��	&LS	k��0�ɒM�<�g]�NΚ��K	#�hQ�D-Lq�<鱥��V݊�ф7k�4,�n�<� ���4-��7?8��">(�6@��"O~}��E�F�*�� �,*��ě�"O�0`ǆ�)��ZBO��"O�3%�H!}�}�`�L�q��@Ѐ"O�d��,T.c(�b� Ԁ��و"O<T8P��Y��\�AZ��b���"O�j5�"����s![���e+�"O�rW�_�����&��$1"O�a�LT��sr�E)�"O�@��G�[2yX�m�CP��"O��P',�%��H�Tk�H��1�"O����TZ���CW+�,mjP"O,tp�I��r��[���8iu�!HV"O��)uB [�����.(_���"OU�dI�	)	�g�R�<b�܈�"O>|KT�T�7Qx�5Dռ%=^�5"O�͊��Q 1� ��eb� Թ�"Otq2�@F��|uJՑ�%R�"O�����)�6�+��u����0"O ���E��2~����Q�>著"O:�R�D�4�,Bu�G$�Btr�"O��9�HZ$
N	���
kD���W"O�A�A���!��(�L_�<X�\�"OH��'E"oTN��a�D^>X!��"Of2���r����ta�7�HJ�"O*[�ǉ4%�6�_/!�2 P�"On��U Γ Y D{�	/Q�}�1"O�P�7oэg��s��XH�L$z�"Ox�FF�"��Za��j��3"O�p�ӣ�4�0�5�OA7p��a"O&��ЃJ RmY��ӳH�����"OR���n�L)!Q��L�6(k�"Oҵp�f��_*f���C�d����"O�E���VX�P`�oZ:w��$"�"Ot]7L�׶���\�z͐�y�"OnH��"
��P0�c�
N||#�"O�PI���BE��*��;:f�a "O~�(Ŋ�C5��!3aʏ=*���'���@s���yp���L
�
�'�� ��9@��g!�4���k
�'�`E�3/�pO�a�疈%�+
�'^ y���_p��U�шٌ$����	�'X1C1hD�K�J�(�����&$D������E��E  ����6D��Wfʱ�>e�V$�)d�@T�a�4D�4���3p(�ҎV�w� 1T�$D��"�	�$�bw����D�!D���&"^�nޘ����2��p��!D� +�l�4U$Ȁ�#��=�<��v. D��X� �.I*`�*�%�
�";D�p�vcVB\r!ԅ,��1��8D�|����CJ���^�;���7D�Z�n,dN� ��?S� !�1D�4	��Ei�j��G\����`.D�1gT=Yz���lT(CV�*�h*D� ófPV�Լ�A��i}��Bc*D��S��ȼ]o���7T�&���va5D�ܒWG֛NVh�"�L� 0<�kŌ(D��c�l΍C��@p���<:]��M%D��cڎh��S�(Ĩy-
��I"D�,A�f�Mt�«�p$�H��" D����
�=v��X�{�� (��=D���GDE8p��G�وpo�s �<D�3
թ1j,K���9�2�7D�� VL�r@ɖ>p��C.�*y_ Q�"O�e��H^�R��1�rl�<4A��"O��A4'�T����Ф
'p�	�"O@s1MJ�*�XJa��j��cb"O|%�6I
*Z p3)4%�B�h3"O�D���T�㴇�ej��""O���BlI�5���yƎ:y�jĈ�"O`2��'$��ayK��:<�$"O�E�*�>+���)�i��rl�|��"O�A���%4l4mB��ړPdT��"O�d����O+�!�C�CjђD"Oj!cQJ\�<�T�h�b��=��iS�"O��C���G�V�pJ�p��-D"O�,pp�)�T�pW�+g� P�"O�x[� ��^�U�E�
��m"O4$ ���;JH��*GN��,�(���"Oҵ0@03NaXwm��t����"O������<��@ٶ�X�WH��83"O\�*����uk�	�%?�Sq"O�NO������H8�C "O�1�e��?��t"$��
"��8`"OƜq�d�(	zɈ�kR�Ue����"O�]�D͌Q���WJփ[����2"O2�r�(A����Y�30��"O���MD�j(��«�� ��"O�}�L�*8�Q�U+�"F�l �"O���G�^Yn`6���=C�tC"O�$ps�L�3!l��Q.Q�k�L��"O$s�A���t�E#�2<K!"O�ԉgӯ#8n�(D�ν�
�zE"OX��1i#3�lY7BR!�^8��"Ol]c�OF0�T�@ٮ6���"O�� ��A��up��ۮ�zS"O���d�X��]���(Ѭ�#"O>i�fEۦcJl������"OD����z�xY�,�6�p��7"OV�:SKK�hZ�� ��q�\�#f"Op���
M=����i�0A�<D�܁ ňXJ��0���/&5+D�;D�Xٓ�����b��>*
�!'&D����`�,;�i��. 2r�<98��#D����ȗ� B��)���z�ʡP�"D�P�*�%B��ʂ��J]�� ��4D�|˶ �.�fLs&��	R��aȅj.D�T�a�RLk,ܲ�e?,v�8�r�.D�T+�ȌsR��t'>�n+�"0D�tks�M�K0�$� cb���3D�$㱥E�Y�ʴ&HQ�1@dQ;�*0D�H10.��y�=j�	�{�Mrw�#D��P�j�C���S�u򬤢�c?D�0�+͂1�B���mMg���+�>D���f��{a�� ЯL':�¹�tl=D��r��S�?�����Q�R��1>D���D`�	&���U�W�I�dG;D� �3+ϵF��Ă$�r(�Q�'H.D��J�� �LlB�s�ˆS^j0��,D����������ԆEXi� ETR�<�@//p1AVG�k7� Z ,RW�<q��`�(ᢆ�c|r2��R�<�$@#H�T��P���`���AS�<iAM9z��GkՄ0�^��bkSx�<�T)E	Q�q9��S�'�:P��k�O�<�a@�s�tR � ?_��x��K�<ك)ɍ0Z&yaCf��eqm�E�<� tɪ"Ǿvd�ydϑ�e�F�(D"O��s� �}Z��W�ͪX�"OX<��ߟcu<�b��QTAF"OX�s�"��;�x���j�[::��3"Od��ĝ,r�n��1*�����"O�|��Ǫ'��Aa�'m���9�"O�F���z�)�$ņ\i��+�"OvH�wnڏ$f��Vc�҅�S"O��S`�F�<hy!*:�N���"O`�@�	odtٶ`��b	P�q�"O�R�d	�5�>�@�����"O��{Ǳ`F�,�TNL�V�@8I�"Of��F(Ҫ'�Fa��� V<����"O��J�(ˑ*Ϭ�`�%���"O�I0�Ŋ;���/�*t\\â"ORP��K*����@
�a���G"OL�VE�^�f,c���^^��t"O<es��*6�d�$G��W���Z�"O���!hCp�T@��=j�<i�a"O(��Q�׊4��ˢ��C��"O�A�� 04 �:�n�hOF%�S"O��'E���˂�6LF�"O0�ǅ\-z��
��ȘfE��"OJ�X��>#UN\�!/Y�7̛�"O��KE+�AT���n�,���3"O�h���5o(A�s��� �0�f"O����������E߱~� +�'I�pr�앭,/��(Bh	%>#
 J�'��%CD�X]�J��ѩH�7?\2�',�TR�CQ�m�*@�4�P�3|R��
�'�6Y���Ԋ9B�=P����-�,!
�'_N��"�W�nT{ D¿#׊��	�',X �&I5׾�3G�@*C�$�
�'��p�1�@,.vnٹ��ǅM�셐	�'O`�	�� �iUN�C̘.�b���'ٮX�! 7[#ꠘb�ֆ,�c	�'M���3�����!�\�|�p�
�'tF�(_��2E�#��tgK�K�<Q� y$ �`GP]b�x׊�K�<Ag,޺u��$xp.H����W([o�<�T�#lRuzr�GF�L�wE�n�<9�H�0q����S��MR@#�D�<�d
� O_�a��Z@/���FaV}�<A�X�"7¸���C�Jd�q1�
y�<���B�IrA�c�ܑg��|!�Es�<�'IU�>X�S�~g@�Qc�p�<��	`���#4��3m���#Nk�<Au��D 2���0?����j�<��D���#��N-T�H��Um�<�C�ˠ$��u��+13�=� �g�<���@�s^�E���O�a��\�a�a�<���*9P�=;NE7X�L�s� �F�<a1���`��c0�C2*�Tī��F�<�cc�sw^DZ1M��)R#�k!�d4�kTĎ!x�
u�K�!�DN�g�XB��T�l�.��Fd_�!�D�eeH��"���X�EDF�&�!򤂜Qb�	�'Hz�|��
z�!��>v��e�&	
.vQ4[�˔e�!��]�z�����+
�v�0��!�D�21w
Qd���"���7�ΰ6�!���4(ۺ�F�S�|�	�c'���!�D�K��M�g��T�\����l�!�d�$p3���6�Ъ5ۼ��&k�7�!�� @HAo �N��=Z�!�R-i�"O�x��P�KlVb�`W(��tz�"Ot�#��$P4�5����C�he+"O�����B3A�*���C4�ܕST"O(����V�8��Y ��)��"O�t �-I�]֌P�5X�5�vq��"O�hѯ��+p����%5��q�"O��r�I�i���M�Bw�q;�"O�����xU<��$��Uk�BB"O�@ªN8=t�|bc�Թk�9C�"O��`��>������|[���"O4,#b�]��P2��YN�p��"O�4���K*U���˂�J5?;P�;3"O��sr�^|Έ�����K0d`8�"OP�aɎ�,����6B~&tH�"O��Y�AƑk���"��6Cv���g"O����@��(X�V��0���D"O�����~�L��qdؠz��)�0"Ohya�'	`�x7��hyr��"O��k�hR�[',(1��;l�� "O���R���8�d��K�+6(
�"Ox���ƕ�r�R������T�Ra0"O�$�`��1p�>]� 䒀nsPW"O��*���.]��b6-��?`����"O���7�m���fL�B$��"O��0� Tj�4�)3�F�U9p�Rs"O��Q-٪D��:��Y`��}i"O �"p�Lj��( #(]$�Ó"O$���+	9;�Vhk��WiTu�"O��["���S6��>(U�ѓ�"O�E���L�������.l�"1"OD�[ֈP '�����,O5_i���"O�![��C%{�zU"�)�]�"��"O�a�U?n���0�j]�3y`e	W"O���"Q�c�(�з&'X`� ��"O(A�/Rk�!2�f&DX��"Oq�@GW��i�����xk0"Oh�#"cׂڢ�z!ч`�b��%"O|t���?V�:��%Y�Z�ƹ@�"O,\�p��^[Z���$�����1G"OFi��
D�V��%�M��Ɏ�z�'UЕY7����\��fM�i��]��'�N �I	#@�fە\��)s�'�
)2�M;(�C�J@�*4R��	�'�4����G�j�n0��Ă�$$��'o�ݰv�R�8z�-)D�8"�	!�'��̣�.�kB$�!�;i����'������E
h�,{2��9ݠA��'M^`ǥɣ^C.� ��$.�J��'d8
�I�U�V-ӣ��,���'���`�*��\�L`�M� %�6�q�'���Q&o�8�XX@Q��EΦ�b�'ڪ0��S�ՙ��H21pC�'D2�҄�LH�5+4�!�x�'�	��Ў|7��ɲ�)m�|P��'40fB@�)��噃�ހh��	�'|d��"@�$������>V�~h �'��!b!ɉ�,�( ����OY�<�'�F�	U��Q+,���E�.��'���K���<��p�V�U#N�x����|R�ě8�"�c^�d:�\��^�4�qӁV u6�`b�qE.��ȓK�ptR�	7:\���K����ȓ&꤫�,��eX�p��FRb����S�? V|�"���[��]YUa��1&�p`�"O��ˇ�V1�����<J5
A�"Op$���X���h�e@�����$"O^�#rOU�%���{�.Ϻ%�.��"O ��K��$��sNyL~T��"O)Kt��E, �0̄�DI�"""OZ��V?ZN�f��$��XHC"Op���J,Y+���
t�,�(�"O��Pס֍���Ɗ�ln$)#"O�l�g�L�#���b`�V�/���"O�܂�B�H摓&O��G6l�!"O d�L�*�%(��X�� F"O�(�g
̩^���0G�u���"O���6�Z�i�IHթV�Rv}Zg"Ob�#@O¼�I�H���U�"O�!H�@��LNp��g�q
��"O�A�2��Q�d���L,�6T9�"O((d�L�^;�T�e���g���"O4q֫�.��1��ow ,��"O�mS��;y=V�P�bj�. �"O��� �̤I>ٲ��.8A�"O�I���Ez��r"�0x�����"O<��W�.#��Sr!]1��H�"O�(��ڐ<����b�L��qs�"O��­A� $��k ��3�����"O6ȻB�޽~��`Q
X��"On��Ufܚ_M
� '�k{�ڐc�"O:�IF�
��EG�I"ex�"O�<�u�4"��,�Pc�if|�p"OPl����l�t�R-N�`�A"O�,���A�J�Y���:��"OJY`B�0f�yKᬟ�
���"O`ٱ�6���p��7+�hL`$"O�q9WE[�@��w��&#�0k3"O��@&��I[O)��Ѩ�"Oڜ@�+լs|��$GT$���#"OtpH6FA���r��1Ҕ�x�"OL5�
�8^�����3;h�"OЀ㰉�CrM�a�J=2bZȑ�"O:�
�&@ �/�'\&���"O�Y� �?v|N9KR�ǗO\89�"O6�qo��#]ఓ��I�b�4�f"O��
Q���p��e�%�'Ic��"O.���2�r5�'�^�\O�}'"O��:���#Xu(�qЃ�?z>���"O�\�7�U�����LSY)44��"O(�R���It!�A��u�&���"O�=J���j҅j~��"O24#��W�A�51-*ĳ "O�A�`G�l b��"`��B�"O��U$ץM&�B�l�@-<�@"O�D��c��]��@8nQ�|�	�"Oz8����@y����&���"O��ْ@ةE�0��B��,��1"O�M�daԆe`��K�nlaA�"O>�I��S/TAL����L6dR\W"O��g���`A����E$A���"O:�2�E�1v#�!撽!~MI�"O�x#EQ�>y�a��n�)Y�"Oڭ�B@!�00{2b̆p�ʰ�`"O���k\3k�R �3�4����"O+�ǆ|�=�R�Du>�)���Y�<�G�86C�f�41P��T�<1cE�w�j�JC�Y2܈�F�N�<� L�q��"԰@���p�:�"O0�9sEB����O
0�hy0"O��;ӄ��aS��s�be�"O:�� ��v�<:f��S�f��r"O쐻w�f?��0�6�d�Ɂ"O�(�D��g@��@�,��س�"O�$*��
�x����oE(gƤ�S"OFԻCC2_�f�zgOW���9��"OdQ��j�[�RLYQ���o��s"O�1��_�E�T�Dΐ:�+"O�$��,6��y���e���0"ON��w�B=z�Ҕkw�b xh1"O�a����X�����	羄�U"O4}��f1{xh�']�݄e�"O�y L�U� �[qm�]9U+�"O!��c��
5٩��Z1�t�%"O���C�2`r��x �I->*�1�"Oj�(%L�͠��e�U�=i
�'�|[򆏍@ ��P!��z��/D��Q ��;c^��D��m� ��b+D��p!�X��%���^ĺ<��-D�����*1�(��iLZh)8a�6D�Dh�á7:F}��u�D�2�9D�$a��=0�a���-4�P�t�2D�ܱ7��L����I\|I��a&D�2�/�J¤<���@�� �t�0D�ҫ�Y:6U�v�ɱm�fl{�.D�\�c̾�ĝ��I�PLd\	�)D�Hq5��(_ T��.�X �dJ4D�؉W44����6	�Pt�`*O��0���KJ����4p�L��"O�8+Rm�-k ��R%�D���7"O�	B�B�`]�х�7J�H�a"O�MA��˯(�ZIu��,�����"O���$B��	u*�Ao޹�$]3W"O� �.[Tm� ˣ�5EB��xQ"OI�D(�	PĄ����I�V"O�T��NJ�x��n�u�G�8�!��۫@���8�����pK�JܔX�!�\�ξ��t,X�R�<���)Ľj�!��??l�U�ߪE~�@j��Y�\�!�
�0�ʨ;��be�y��ޢ~�!�O0� 2�#6��S���j�!�$�n�X(1"��Co>�Р�n!��+)�1�vE��l]���t@��n�!򤁌z-!�#��{>��w�.F!��z�Ⴑh��4>нJ�,�%N!�d��`, ��e֮gRX}��JO�pG!�dبP�`tyī�"?�����"Fs9!�ğ4x{䠨ԁ�W�<��@�D.!�d�.C�,q�ec�.���"F��n!��/RQ����mˣ+�rM1�`�'g!�Ć+!�S.�l��̡g`&V!��7!���ƈ��:�60CBA� r!�DR�Gl^��3���4�(֯���!�dX욈��	�%��X��O�#!��1#��j���?z�D�����ss!��ΥX�p`{���3r0����!�*��y��L&]\2�9z!�[�&�6��` %;UH
�i��t!��<)ʄ 3��& ��g��\i!�i�ڰH�k��b:5�զW�6|!�d�>��hcge͇)�6���4
�!�	t����D^f�F-�T�>�!�� ����W�]�̺b�ȭP3B�9�"Ov��h������,V�e0v�Y�"O��w�
�Y�6�:P�C�f���"O |Pd�q�����	�y6��"O$�EM�=#��$�I$�"a "O��[S)וP2�J�fùD�H�6"O�q�1j��1$D�{~�!q"O��������b�@i�@��"O�ñ
^|�Q ��>a� ��"O:aye�~-��Cr/�9a��x�"ODmaU� H0͢�)d8ؓ5"On��k̰_���YC�B�tJ�"O�XA.�%"Vl#�M�$,��!"Oz0�����q�P5�`�@�}&�r�"O�(�M_�M>��s'���B�>�PS"O���3��0�Z��N�y��a�"O���@���BV�����bp"O��yu'�/fQ��#&kƋV%<=Bb"O�i�q�_�A'��hĀ�ĥѓ"Ox�vJB�>RP����*���"O���u�V()�U��1����"O�!ʲ�΅�|E��N��T�jv"O�M�D�Ԉ� c獏&��h�"O�ظ��>@��I��
 �,~칁�"OH�HT�P wS��B��(d� 8�"O�\�B�w"�� bܿ^`����"OV��`��
G�)�r#P�ZP��Ұ"O^��p���>):Q��5MOr�K"O�����V;_&�� J�%rB�%0�"O� ĬҀ4(�k�I�t1d��"OX���	F�
 y`
�&��yh�"O�:��Q�?��]I%i�S��|2�"O�qIuj��|ܠp�ۢ�"	Cq"O��ÐǇ��B�+�dD�T�X�R�"Oֵ1cÔI%l�iqㇻR��E�"O���Q�R��`��)<v��s�"O��@��=5Z�� q��	U��9��"O|1���J�4�X�D�0M�.� �"O.i����R�F�5ϣ{� pr�"Od�×Dާy�"q��5��yo"O�}���]j���!�l��J"O�Q@��ưK��cQA��,IKW"O:-
��I4�j�o��'���X�"O�3ELU�b�\�E.��t��C"Oj�+�`ͱ4�P��]�����"O����H�71
�����4"�V�+T"Ob,��;)L288�ŗ�-���34"OD�7�_�:�@��я�F�Ac"O,�1�B�v`����I��dx0��"O2!kE�[������HA%7�^a"w"O,m�����|ٶ��0S��}�#"O̔C����Ѹ�đIc��z�"O���6��*NR�z�FӣWf���"OH}��C\78f���P&��n^Li"O�1QǮrJ�P�ɫ1V�5۴"O����AWP��2.�f��q�"O8�� �-_�bx����}.��"OP��fB��+
\�i�h�^�#q"O��c�F�N�ұV}��<��"O���`��S������T9!�V���"O| k�M�a���f�~��!��"O���,-��4�%ݢb��Hh�"OF��p)��^�!2!A!9��8�"O�S,��*�8DP�6�P�x�"O� �ի��Y�c�Z��s蔒B�J�!�"O��0��àWD\� ҥ\�H��W"OTyJ�.�L䂀����)�\)�"O����~d���BX"��c4"O����J^�	�tM�w��e� �"O0@���U����	Ԥ�)e\N\�V"OR��4H
H�&�C<*���0�'�i2��E J?���P`�w�t"�'��sुAddlS�[�9�n���'��К���6�~���IX�7NL�
�'��I %B�e�*�)��ʰ�)D��x��C�*��=y�M;�4��:D���C��?MP��S"Ջ Q����`7D��h����T�xf��qe5D��Y'����Qca9a���'+!D����L��+�Ĭ3p�ѕ!��Uj��=D���7��budQْF7"]\H�q/D�4(��zoB(�,�n&��R�.D��H�mٹ��S��K�?�a��M-D�Ȃ�e�>,@<<�ҩD���ř�-0D����ֹ.�H����H�d�b��/D�<��pFp����F6�@)0.D�`��[�O�!��oӋ X\x{�a'D����(F�|�L���j��`*6�ذ�!D��GhF4^�����:P��
��-D�{W�U�1`���VK�j,��xQ�.D���"�����ЍJ��H$�.D��*�'؝>l�Kr�ϔ� �
�j.D��A��S?N��ء�L �A�N+D�\�p�͡:�4��"�I�;�ꜣ�*D�`�2l'I�������g�&D���cg�J*Y�CD�]����'&D����ɞ���Uh��KjNM���#D����瑅f�e�D/�V�虳3�=D��;��T7̹:�F23��iW�.D�`
�N�y"R��$�&��8�H D�Xb�c�K�H����M�J�b�	V$?D��r��"z���x�b�7M����>D����DDV�[7DۭL�����7D�lH��S�Y��#$%ژ2�~\��:D����/��Ȥ�����D��"�8D� I&�҇ :���#(Q6 �Z�,D�l��#M+&r�L�
����%e)D�X*�Y�:�ǩ��Q���&D����d�99�Dls$iHk?���$#D��� �ɀF�$�8kCjѶ��d@5D����tlؐҐ��#��Y�!�d��$�ج��3� �ۃ�ދbp!���,[�&�b5iG+&�N)����1h!�ůzp6��
>B�歊 �Q T!򄛑[��6h�$�X hA��3/C!�DhA����)#��4c'�B$!��̈́rԙ
��G�v 
U���Py�G5P���C��>o<�s�E7�y��\7Z.����"UL�E����y�"�+z�8mؒo�!Ph!q&�(�y2�M�.��-���Iм}������y����t��!�k�zq+P��$�y�*_+���)�e�*���Xt�E�y�-N� +���穋�& ��.��y2 ɫ ����oI�|��!����y�f^-M��Q�C�^����!��y2Dҍg��E��XO8�����y�oĀۤݺ5�5?H��{c�+�y
� VĲ'���|�d��mz���"O�E�el�&lu��2%sx`|cQ"O��ըJ�F8TYR���	�; "O�C���j��H0�&9�"O��8�ϷsL(l�S4�p��d"OV����[�<Y���v�B�ve�G"O4�!S�� |(Z��%:��a"O\TA�-Ɓ-�(��%k�e�"OUJ���t�8�!,]�x�a�p"O���f�F3ĺ��TJ��}P�i�s"O��k�&�Zj�Y�OG81�\�"OlQ[��:� |b�׽O��I��"Od���aC3j���`�h	*(�y�r"O�Y:���>.mA�h���ź"O�|� F˚g�Zl@�Ƈ5~r|�C"O@���X�G��@�e�Ŧ�R�"O�0���C oV!�BȦ=�$ ��"OH�킫0����'F9|� XH#"OxI13%F�tdy4'{�,۱"OHĪc'J�9|����HAl��d"p"O�2��u�|�V��/|�1�"O�KI�>@� �ƪ6k�4�a"O�e�5�M$�8�w�ګŚ��!"Od�8	�3�z��g�EbxXA�"Of|�@ŕ�[b�J7Ÿ@3��"O��;i�bj��煗 Q�"O���P�ٰ,�`��rII>��Q�"O�� ���kn,2@�ďT���1"O��8a*�I�]8p�X J�9��"O� ����B�G�-v�D��-
�!�� \A���U��#��#a�	^�!��U���F�]�_�T�gA�;u�!�F2u���N\�3 �t�!��L.n0CƑ�yg�0���YT�!�d
+�~��eI9HM8��֯ذx�!�$ �.��!i��;MJp��O�'{!��(N���I�`D���H�^}a!�DѺYrf]����8����q� к��1��V-�;����X�g8���,��l���K�l+�i�t�3Ĩ�ȓ]}~L�1��c��j�o�.�(�ȓZ��zB�x:�A�p<��&�LF{���IP�L����0F{�Y#gP&�yr�In���Q��J�A�fU�C����'��z��K�{V�dK9o\|��.��Px�i,��H�Ȗj�����4U�x�'�%�'F�a 	2R�.X16��Ǔ�y���]"\l �jr�$hC��'OC4c�!�D -,ϖ�{ dH1��uڲ�:�!�DѫA[h�sw�0#���c����!�$��X͢1���[	K�N��F�&�!���9 �G�/������Y���)��� �#��%�q���q	�t: ";D��nF�u$r4��P2p�*�*rX��Eyb�|_�Avg�XjU��� ��y�� ^!\�y�oCGҍ&A�y����_Ȯ�;2��O�b�ە����y�҇H!BI��.�.1�`I�U
���'�zBF�!�P��*E,3�D!�G,���y2$4t��h*��W�7��|�6eP"�y"-�gq��2t-�6 �����y��ۭ)�.H�F�Ús����ѫ?�y�B['^���'kc� y�	��ē�hO���H��jTY�M�|�!a�'_��� LVI9C�\d�"��% 1�E{�"O���������ЇaN�DrU���$�S�	A�A�yU���X�~��cc~!���Mx����)�8��A�_ayR�2��� �}���u�@�"��C�I�Mn����	<n� %)�&�C�*>�d9JgO� B��cc�Z�`�lC�I/%A���% ,0X�wU=
{�C�	-�~�5�R�W�X��)�JA�C�ɰR�J��P�>�B�9�[&Bq�C�I�V|
`'.�2���;!ْ9
�B�	� 7�!+��,e��`p*�-�RB�	0=\![�S�EԬ��u�R>+(B�I�aϬdbE�Ƙ�p2&$��g��C��.�\�J�_q�l��/�[Y
B�ɶ�:�p)�K�p�����	m��
䑞"|��3ʾ�1wCV�LXµ/>i�C��?�D(aeZ4]4`�����`c��	�.�҅���Kzf�`g��T��	F��?a�
2��E� ��4,���2Sy�<��E�)k�~8C&�6�Ձԃ�v�<����F������bD�Uu�'��x�I�&C�5���m�Y˶�q*�=E���K�����f�i˦�w�˵nf��ȓWB⽙�L��}XzӠ)����|r2�S�W�B�����Vꄴ��v��&��7�A��&@�,�⤅�?G�i���o�`쑂�����ȓ_��,� ��'k��h!t�X�U�
|�ȓj�dk�@��LyV��g->!%�D{���AVm���N4��RE�7�y���4.x�My�������G����y��[1N�pA�v��&x���c@�]
�yBl֗wd���2eXЊbǟ��yL_T�nhTJ
�|������@���?�S�O5�Q례

O#`It�׆�~e9�'��T:��Ӫ0*���a�
���\���=a��Y�)7t$*����t<)7 \�<�q��YG\���@5 ���Pd@VV�<A�
�%;��{ec۰kF�X0g�<�t홙N/��ʧ�0Fb���L`�<10I�yT�KT	�*�*Q8�C^a�'�ў�'A�EQ&��/!���ˈN@D�ȓZ��0GH�i��]�H͉U:�-��4��U�Do�.�ޝ��mBK�N����L�w��Z���@�V_̄��3;�0�������a�L4
�HI�ȓg;�솕$.L�!"4@l�P��\�$%���8[Ej$0A̓������k��8�pOU�M_��;���> j���B�(��)c�eR���C��Ɇȓ�F�pT+͟^?<��W������M~@��g\� �LA����lH��=jg+Q�b��YQFS!RTM��6����2��y�uOv�\]�ȓ-��mK1�ٗu�&�p���G�X��	Y�� �X�0���9/�#�Ԇȓ*T��e�z���)�I+p�)��k,��x%��'Ղ��"��fA�Ԇ�;iI0Q�7�V�B+I,-�<!��fHܴ��F�,mZВ��1&���ɂ����9�V"b�G M����̓�(�!��E1@u�|p�d�
$>H,��Ȏg��)f��A�jQ�����������b�J�F{��9O� �Y��D�O�D`�'b�n���:D�>Y���)ʏ,�Z��3D�%$|]K�)��!�$L�{bZ|2T&��2l���㏜K�D/�O���d�,D���vؿ^֕q�"O�k��=��ez��	>��"OT؁��V�$�X�0�(PG��ţP"O(\�b�5t�A�Hϫ'}�4@�"OL`iҨB�S��pq"�F90��Ż�"O��*D��!Jv���V�N�B0��"O�HMS�F6 EBV犈��,�"OR��P�F�J��e ���z�*u� "O&u��mֺwz$}����qJ�J�"O�0a�,^L]-�iA�Pr�B"Oz$�����d�� �5�W&�
�"O2H5AK-E 8D�#ī&Zj�'�@�'�Xi����k����ʖYjX��'-��A�ˤ�������>�<��O�ٮO赧O>�yGn��62�%�"(Y'j��3:D���"-h� �C�;f����N2�J0w-���>�A�Юm�B�^�4M���35s���'�*�"�-�-r���"h�J"�B5�$�|x�<�ҤK�,<���%O5�PX2��7D���±!2��STnр~N<JWLTh<1�I$�0$���Q(*�Ĕ�B��BX��EyL�F̻�ؑJ�Y[�@!�y�,��J8�� ��F�(`g&��yG�K3� �� �>�¬@���y��ƒd���ۥf�<K�<3$���y2/R�#��r��?B瀙�ڨ�y�&�=U�AZ�B[�B��������y�'��j��P�R&o�:@�ҍ���y�Ȉ�-�D������S��0¢S��y"lفb>��cW �3�)R�!�yҡ�cZ�t�0a\$��9
�y��X�L�hL�W6Wl����A��y"*�B�S@����8�����y�4����w&��	����dJ�6�y����JV���\n�ZX:ԋ�&�y2Ҝ>_
ђ�A�k�(��s�#�y򤉺r"��@�f���CDE!�y�gJ�nnx���΄Y�>�*�&U��y�
��p@(�C��F�� ���y�͑)�\�@�o�AXCM��y��ԬӨ�BaF�}�vx��K��yK�g�*��
�{ee9E�X%�y�(	�0�Dy���k<2�Q�e �y�a��;�  R�f�"� 4���y�+�:��� Ne~�ȸ�/ɰ�yR�F�~�jˢm��]	�`�����yҍ�4~�5ȃ$JTm�iAAd���yR��7ЅH#CH���Ѡ��y�b�='J�Bue�@(y¡��y�E�skX�s#*�;��jrI���yb�
��DK��J	5y����B�yB&ղ|{�)K#��`ǒ�y"�V�k�r�BU/Ŷ��lҦ��4�y�gH��́ԏ���y��*�y
i+�A�Y�X���% �y$]�$Ej)*S�@:L>V8b�̞�y��ږ.bh�%͉�>����ئ�y�ǶR����� .0�tА!��y�i):��;�����{�a�G�!��aC��Hg��CI"�Hb�(�!�D�=�\`sc���I�Ĩ��-�!�� 4��A�Y:Tk�b��b���5"O 1%W�!)�2�!ը	B���"ObIp#��4.�p����>uT��ȵ"O�T ��_�c���r�n�
Ns"OD,
�H

½�1��t< ]�"O�:燊�2�3҄��IJ�	T�'*�8Ҕ��8Vک����{�Z�1��	uB��'�� ��	y��u�� �
i�a��'+�@�lF�
i�v�O�oZ��y	�'��M��oӚn�V�Ň�n���yB��7Ĥh����H����؀�yr
�u�8�#�ڛL���>�y��ˣx*p�j�ば<�*U�$:�yb���m���Ц��0N��q�@���y�ב)��D�i��))F�����y�@2:m�|�'�ك;��r#m�,�y�M�y�2U 6�MO4:��'I]�y��3�x�W��D0.q�V�׉�yRa��s� i&�����U�7�y�/^�9�	�&��;QZ5�X��ybn�6O�!��������ĉH�yr�?`��;��4jQ�EKNS��y�͐���ж�^�pnᘧ@��yR�Y��#�g	��ʗf�
�y�a��1�,���D�U�42����yR��4�Ve�W�I= � l��yB�N��B�ZF+D�rL�ɑ ����y��"A#�hЗ��}��a1A���y�חq����.��Jq;�Z��y�%�����[�"f���
��y¡ֹkڞAbW��?��*��A��yr�@�6un]
�m�[l�Y�G-�y"��4	�{���j�J��p?#��:��d��2�h����J�;��,��$Zh<ـ�E>�����B�a���ȅB]Q�'V��g#Q":b?q(ʇ)	pͻ�腁:5<����'D�<�F��|�&�`a�g� }�U8O�뷬�	 �Qh��"~z�O�
y�����wF�t�D+Y��yb��Y<��)l���������$ą:;F};D�W%NM��ɼ>, ��[��jdƀ�
v�'�t���́ݘ����� ^(���@Åb�:K�'�V�,,�@�)$Ȍ}V-�1��?��g��$��@r�eX6o�@*�畻J{�'n��4Lϫu���!d�M&����'��j�wd���԰M�e��LO&��th
��'l��b�İ�d}��F�O8%b��&n3J[a�G5p��ad�#	��F�b,����'���D6"�c!Ѳ{h����d�86#���a!ܢ����OaV) ��H�`prd��y}����M�j�L�v\[�ࣣoı��O�����7!69i �W��t8W�O���)I�Q���'f�8KB���Ʀ���0 �%H*{n"����I=iP�7gP�-n3/�3;��m�� �${q���ӨYF�`�6*���3�F*9�6���儯Zl=a�X�9,v��++VX�ҕ�V6/������(�y7���d��x�!(����C�R��p?��$	�>A�Yr�'�a�zł�.�)_�t]8�CŧRvV�@���ؤ�%�A;RlG��b�vݲ��(\�xE�'�XxgK�(B�A�e��848��$��t��a�҄Y_�V�[0�@��D@�c�%L��E� �B����;�D��YU�
!x@��;t �J��� ul@��БG��I৚�P���t��r�Ȏ�9ޖ��+���r��&�σ<ܒ��u�Q�3� 9㖤O+�dh��D$g#ԩdQ�lJ�����3[3���'L�
,^,T�wF	V���^)~�B��2E���t�PA���\<�7�(Y�@�tO�-���.�t��S��7>y��b�κ&�h����;�$�CN*~�Ae��o��i򡍋�'8���� G��M;��U�H7�]y��GR?�0]F,��f�ݥ��ɝ#�� �b�H�oȊ�3�Qf��>)�h�*����vLٿ�Ɉ��$��@�ӧ�"Ch���U�<4�pq�Gŗ<tD4RA��SBi��cL�ty\tER+�&9R$���#.4X!��o���~!_7�f=�1�y���e�R�.�Q��)V�Ѡg,ȦY�����W#,p��ۅ���S\@cUH��4��	��`�{Ǧ��g;Ѝt0i������<qgءj�c*D_<��`h����͹S�`�s������@� ���7R6��q�AJ��c�O� )�dH�$o��Z�"��	H!P J��I↹i	R\"r?�,:0)ѽO�.�	E@��!1h�K �b�0Sț0����Վα^4��@!�3V��1��	�Y�� #�R�/
$H��I�t�	�c��	g��ۖl��ʝ�n��9!8�����?k���.	q�����>s���.F�br:�م��T��	-u5��c�;��
��>�X�2��	�:����/aӺ�ۑ'X��@u#W>[h�y#�::o�yc!�T�2t��'Qn�Ss�� [�i%ʝ;;�t���Eǹ2H�1�UnP%W�Ɓ�C��*Z���_�}"5�;=�j���w�,4-�(�ĉ�$���3� aI
�$�0Bd�� �:�G��=�����V�%�rq�'6�5�SI2pv�Q�j׷� !۷C�:��9�q�&�~mS��O=,�@p��6@�9�`O����Oz� d���6�,96`þ#�<Ձ�/Ƌhq���@� +0��!9��'Q
���in0(�fW�"L���TJ������aƃSm�O��P&[�i8��NF<7=0�:��'d��6��R�j�KSCB(&���p�ƚ3o
.�A��ƽ44&�B��b��"�Č<	���u�)>(��"j��6G��`Y\�>��퉘k`݀S�x؀,�d��� �>�衙!��\X6�Ɉe��hS�K�o��Ԩ4Cc��P+L5�� I�f�
�.`���=P�.%9��'�Fɓ�$\�-F���{>��9�D#���'ɍ�a�X��GCI�`N�] �J��~���pF�řz:��aV�؇$�ȈW	��c�V����� .A�u&�4=�}�@�l�'�ث%���2R��kL9.lvt�Z�����
R��xi@�ڨX~��BI��/�dQ�AkJ�Z���'�������W���hI �*]s�➤����c�-Җ?'KP9D�T�p�uG�����K�ɂ�{N��c9.�pWDيo���yQ�	�C�H���T�
~�8D(�
un>P�0iS�}�ZY(@ ։E�F�h�f��p=���F:��|��L�-a��Eԙ({`��쏦�Zl�bQ�HS^���=��p��E�+ e�4ET�)~l��`O_���Y�C��X' i�TY�����AC�R�ѰϞ<Y����;�)�����?�ym��t[�����4FR�d����{��Q�� �o��Ȱ��jW�@�W��h��Y�A��\�1��\<I�O���w�5�hY�&�߅��Z�+	:|)��q�mV6�d�S�V-���`���"cnTk ̀69�~��Bh����q���7�H����*��b�`y��2-�r��F>/���2a�$ƌ�r�_� WvЛ�"+>|Ab�.�:Eg�>�s䅃�+@���E&��p�b���T4b@�C&T�ZN�1�L5.�*�r%�ƴ��<ɴ@���`�.�U伨I�(�>H��QMͥ/�&i%Nڦ��g�@�\4���D�'��iq��?}�<�U(��ir���jN�yԘXӗ�	?v�a{"�Z�h�f�n���$tw �rHѣ�X��p �i� �.�~��-Kab�&�@�>���'ɟ1-�=���Ii�|x�/]�E�� 2��%hB�xa"�	�% \�`�^90���y�@�O׊��`"�Gꉳ�A�n<�A"@��:u���!���y,�l2J��wnX<>� ��яB��f��`�,r��'e*��J�+"ϐ�a�']9)*H�qqƂJ��zBl� q̡�2���l8��djN)$����.%V�	�FÍO)���#O�:Z�4��d��6V��rE��:(4��S� KG�PHC�'��M��j���}q*U0,� ����_���Q�E�^�ڴ?��!�K�=a0b�i��I�J���a��L�|�Df/s���A�Y����FV�q�ܜ0%��3O�D1
�m�70�$�FA�Mk�)(Gú�&��q ����0]Bu(��&��(����H$lR<����%n�����$���=�#��'jr`�3��Ÿs�&x90�H�:�NP�6!��rĔa��5gj�� �#v�9ߴ3h,�fl��\
�h���<��Q3�� l��X��M��~�O�6k<^��B$�"V�ъbb	�y�=+CP
u��./)�hW��l3@�������k��0v��Dj5��Iۈ()N0B��Q
e�]$A�{�����"7M�H��d���%���ax�:�%�=��� ��J.X@\a�O�_�6-_��Tm���y��D �P쫖CX(�Iqb%��iL`ƭ�j|��3'�Q�$Q^����'g��+F苐*dfpcV�x�����S .:e�"� 5�h%��+�>y��[0� �v��<]�|q2I��yy����?��L�7�'FNi9U+�'��>�+L5y�^�9���W��\���+;�ش�D�]��mQ�f�	z� K�Lx�,l��kU���y'�,�PsvSyl��G�Hr)�m���e$27�T1t�ī�� ����t��[�ɵe�,��'8��(�"J؎9M�I{v�Xd�@ҳk� *�����e��z۸8�� �Y�
�CY&0X����Ji<��E *66�Qb3� 	yܪ"=)��.0�(e%�++�셀k��Ϝ�ra��RP^����_��S`��?�R�iRJ�S�� �y�P<��-�LTW�4��gEQf�y��K3�@����q�H�E$�B�iE��q�R	�+�_M��yD��R;�]
N�W��d��T���1.8p)���e�B- Th�%˅7B����bln�Ǔ�]�&�� ����Xj���I�G3�!�DΕ�D)x�µ����PTc�>A���-}�^Q�Ĭ�!֊mJ7j��~��h�Ŧ��Re�c��-BJɌLHYy��/\O��zB#�W]Ȁ��F��|ǼcP��UQ�@2b�չxB�+S,
0��`	�ɦ&�J��gA87ϲK �-ғ*;�!sd�	&,i0��"�#.��=�w��p��-ء7G }yÁ�z�
����O2�#"I�SJ���a��`���2:+��	�d]X����ʎ9'���!ȌC��X#0��.I(j<H
�C��� �)"#��b�Y�#:︩����g@v$��M-!��� �"O�-Ӏ��� Ѳan؏%�1�p۳|�ah�O�Z������ �!Y0���D]�'
牔x DTCv�R��5��/�N������h16�J=!�AC�a��D�� #*}A��פ..�ES�!\E��0c��� yt]ʢ�4��O<A˵�>c�$̢�NTf1���I�8IەÐ>b�&�	�Vb9��'+����iŝ_:z�h��F�!�N���y�T���V-H�Q�P��$���9��8�!�� ���������G�(��Ub#"O�`iCLDK�P��eL��z�hE"O�DX#���M����@���p�L!x"Od�����45�!Xb�1P��dQp"O�R�BT#/��<2TgQ�z"O֜�J�n���I�F� ��"O8�s���|����fF���j���"O8e�'���4U��R�	#��5"O8RGL�1��W�ߏB`��d"OVPCAJ�k�`�7�W�n��1"Oؙz� #O��#���!��H&"O�z4��a���(�	з���Ӏ"O�*�L:�:�ԋ�h�v9su"O�0�� s�و�T9��]n.D�Pb�F�?���� 3�f�s�b:D�p���;�ޤrc#��[F1���<�( ��r�QP�	��i�j�*���(aS�t��I�=�JUx��"~�r��EI�md&Uz��]�ZŦ)��G<p�S�`��36�A4�Ϣ&��F|�(ǯwA  �&@f�'{nv}����!��z�e���ȓ>�<h�7�G�rځZ�����%Γ|dl(��GܪPH�ҧ��Q�N
��^�yW,�<F8X�8�"O|#�&��g�Vu��ʒ$ꤒ񖟼Ҡ � V�qe�'�,�@$*\#Wʐ��t��?��
�O�H��!A�r]sdNV�T����}��Ht�7���J�b�`�Sq��)>��t��"&�Y_�u�'�؎}-h�>Ap��Z��bTF��Ӱ��"D� �ЪJ��B�#��\ <ǔ��
z����Ĺp���S�>E�iY,)�������0S6:�H��O9�yFL�C�Й��*�,�V��ɤT@�͚~X����K�3���OʋV�$	p�/D�\�1m�(Դ��u�O�%;8)��-D�  T�Ed�s�c�q��@�k*D���&#ŏ#�氡�J��H�����+D�쫤���|�0Z�l�:|o�M�U�/D�,J�g�z֊��k�?+�P��T�#D��uG�Y�Jh�H��w^����5D��+U��#%����"GW�y��0D�Ț�`�63����-^z�˷�1D���p�]�e��aƅ_�g��s "D������+m(�������l��ˀ�#D�x�D�D����a�^ #���ѩ"D�����A�l:��G�(`n�ъ�*O�� .T�6¤�*�P0'�t+�"O<qY�*V E�u�҄=Q��%�"Ohi(u�L6P�Vْ�׉K����@"O�0��F�.��غ6�X	gغ��"O`q"�:J��2���>�X%��"O�`�����0��ㄜ�W���""O)��C�mxMc����("O1�DhY~��B׫ڵ����"O\A�'ZFL�j�@Z��-��"O����D�a��A3��C�$h���"O�<�e�ؕ/%3D��G�ִr"O�xK`�=*v��V�'�4�a"O�
Ꮛt�rxB#	����1"O���$|���V��d$k�"O�y�BD��Z�B�<�ji#�"O�5Xt�X0��TzAB�b9LXA"O���#�!3�%�Q`�A9LYx�"O��!s�A�_x*� "):�g"Oy�	J�nR�"3���- �cd"O�Y*�Ô-6M8
�2"�9�"O
��l�=6pH"@^�vQt0HU"O� 8�cL�"��hJ�H'+�t!c "O:�f�Jk�]��Ʉ�V�rh�"O8�r�
ԷS���H��"��c"O��I�0j��}�Wf_i��Uy�"O�@QA,�9��V��@��"O8U�l�^f���IS0��0"O�aBBLߏLva���A���D"O�4v��|���!"�_E%S"O�Iv�P`<��b4l��"O4U��ׄ=	b���Ʃ!0�R"O
���aϒ�p�ـC��3�q$"O~��m��%�Hl�6�Q�^��Ѫ�"OV5+s�wz�a�3I� Ҥ��"O>H(Ҁ�A�z�pi�'jl���"O(`�dF��ȸR�L�+$�T3W"Ove#��,ٲ#�G$Yd"O(�kE-�l���9�M��"ZܩZQ"O�P���dɓkK
CE©I�"O/P���Ǒ�)N6��0#��p3!�d�M�H���kD<r-b$�%�� #!�ĉ�)z�b$�N3	�z�#�)i�!�Ā�	������ίJ�,�7D&�!���dڸ�ђ`�-c�N` Rf3;�!�[�rI6������|u�$G�T�!�N�-{`�i�o�#��1p��@�	�!�$ǿ'���pS���z6���@ 	!�!��%ʌՃ����OpT�J��-3�!�D�f� �Q�H�&Rg�L�ѢY�$�!���P$T�1U.R�jPJ�! ���w!�dނ]�ЁQ.2]'���X<^!��}.�)u��4s&�e�m�!���*IB1�p�t밽2b+ڌd�!�d��P^����8�
�����[#!��Y:���2�G5Y�����h��++!�D}�Lɣ�D7^8��,>!�Dڔ��a�,�,S)�-�P�,;!�$/_&�љ�f�9/� ����P�~�"T��x���?:��3����yy���Q��x��͎_p9rC���<s&��5��O>���b� Dh��~Zu�Y�l!�����(���Q�<1BI4*��A"�O�?M��y��	���H����%Q�x��Ԯ>?E��C�"f��8�gւo�b��3�$�!���"I�@�kƎʄ6�d ��֎-{�ɳwP*�aV���C�~`��{1L�G-�,�29+6�ʞ'�䅥O8abv,�=N1O�)ҕ?I��C��+G���nƱL��u��59}����^p���>k�0e���3y{���3#	�}LO�$17��>�2����$I�DP�On4��?��(�Ed �����S�G��<���'��8�%��)�|���� m�X0 ���.�`y�"L+j��5����Q��7m�,-U��(���O�hJG�Ӎd� �.�:�xP���ɺ{�b8[v��<v?��̟�!���\'l�8
�V,^�~�Z7I{�ޑ��̕B����+�-^�.aG����[����/	�]��$�1)V�~�e�{N(�
&PJ�2�q�[-[\te���S.f}���`��j�B���T�s�V����W-QR,x��	��w��eʣ ��IѶ�s�	m-,�8�(Z�>H�D�� ?,(��B�r��Y�S�U2M׼���ҋh&:��;0��'d܊(���A�A�F���	�/���.O,t
Y w��dD���6OC��`��v�x%�D΋o�<�ѡ�/	Eh��gB���V��<	�oR&��l�%df�+�Mu�'�.�X"�ڒ)�|q:1��?1ݺM3ď�31|�R�f��.��JϽ(�"c�.Wh����	#;����2����O�P�� .o|"�H5L3�4���Oti�c��(7o�E�6��6Z:xI� ֵ:�Z�*Cfنop���X���'Y��=�����w׌1��@̈́)����@�}��Q��
$����!l�́k�7D$�\(�hɻ��6-�z�����M9ǣߣ ��:��-r�W�"@�P,;m��~���i���n�G��(��Z>ee�����3;�� A�hJ�E���M9Y;.�Aǜ�$� q1CH7z�Ќ��S������:���R�'|Y�ppc7�[z��SJ��&
�E�'�H� 8h��G���fM�p+W"_����Ƞ.:�2��V5�`	��m�}�(� �n��� RQ����<X������#\�����O��B���;��!�r��:�6M �߯@�nT�J�*�@�۴(21�iC�Y:��(R�lf09�� �2#�2��$Zd̂�.ϱ@���#g��,sU����_��(SM];sm
�r7E@�]�֫a���3�N� _��]�>�x)*��޼y��A�느~�p����:�D��@ٝU-�������9$C�ț  ؟S%��4�dr7�I�}��� C�@��j�!tG��"�H�����1��j������DG}r��:	I�)O"!p%��+��%�V�!��ȐA�4�H��؞;�`�*��֜)d�SAW���aC��b��K��dʹ_�huJ3(ӢhQ����Cm��@�YÒG^<a� �,Q�$�aD	6+t��CQ�jӼ��uj؊V�T|K�gIh�dg(Y�?P��@o%�O$�a�؅;'���ƃ��	#�hg�Üa��a����o1����"�s22��?/����#>
*�( �3�����i�)+���h�dI�]���'+���D�:��h��*S-2�Y���d&<�c?O6�B��[79��m V�B�?��\�4ʒ�=�e�C����􄁆�ʽJ�8f��59�e#��N�w.�耙�D]
/$		0��_̚]
`��>���C�G�<��yȥl$
\��ڽw{�Ň�ɿ)lvЁ��ߔ#R��H[;[���DG98�E!b%̀B������=/ch��s��&Z� �h��]����R�G9)�^ Y2 ��]ݎ�Yc�ٟL5(��
O&y!p�ІL�rU)�χk����5gӕ�Y�4��@�L�VJٻY}0MY�LI�xU�$φi����E7�,ys$��F�b����$L��4�'� a�"RHؐ��@ؘ�L��phMo�09Kc�M���qυ��ڤ��(������X�B�᠈��h�*+O��ar�.�Zi��	
�|����	�=�eK�Л;ZN�(��-�ըmP�0A�9�
��A����ӆ5��	s���!��)�-� Y c*Z�4������
N�f����V�W�!a<Q��e_�Ii�?h�t�"��RP�q�%^����Ƭ-&o m`1�A��YSWl��2�$�h3$�5+P��N[5�K�3�&���] 6Lt�*��N�zHˑ�W6?ԝ8��X����$뇷�bY{0��'8PL�%
�O�ft�qN�� ;ލ r��/��X`/�?��5pG�\��{R�؂t��٩uLJ�)dTCUd[�Y�j��@�sf���i��D󷋘,!�T ��O/���v
	6x���zb�@�W6��B�n����X�E�O��<�:(S���Նf#�]zs��T�zd*U~DQ6�٤4�F�[�d�:K�n���酽8�"�8p`D=CC������,O�@��S� H�DH�N�p�����RE@F������6��i���J�c[��Q��i�"���`� �\Yx6L=��&�ݥV�
�ۃ���f�Q�ˀ�;s��"��/5�,��qA�Q�l�ڠ(6����*(���b���]��[',�:�.���* +�����L�v��6�ӄR_F)��ۂ��)��Xp6Yu%���|15�7�`e1 [k��8	�,�x��m�"(蝁R$�Y����3�:c�Ț��M3"C�/�z�FQ$bII���ȶ��4K�#PaizVDз<��XK�bU!T�АA���?@�!2�*S��O\i*���(F���IS�\::s�L{�'#*�j$�_?E��H�X.~kl��TE7t�s�/n�f�EOL�9��܁� �{����`��3[���K>��G�X�z�*��RQ�)�d��{brl����+gZ�Q�Y�H��㇆5\�l�B�E�O���J�1}n`@�v�I�e}��-Z1P�0�����(h��0"&�M�=Ҹ9K�S��<1g]4 ��$)��C���E���Vz�y�ѩN�h�Q�	ڦ=s��9g60�I��Mk�O�촋@���XP��l�{�A�>�������GE�9,��a��rwi׍���mZ�61(�)��®C�*��4)o����7ol����&[:��"��b�ś'"�&���ӭ�<_(D�&�	�u�쑰��Ȅ8a�HS�/�ަ�;�_.&xl1�OY(�D0�?r+���B�G֦!�c��l
����D�}SR̠��^1=_�}�ƀ�x�H|�Ip���
u_��5��3 ��]�o���ig�2_��{���N�(��+˛rP�)'�0A��C�VL��v	��*j�ybNX~�*d���Em�.��2f�%"�M�7.�&��O��#p͆c��D{D�S�(/X�Vͽj�XP�h�7CO*��i���� mӖ9�J��p��� 7��i������vĞ=C�쳇�G�/�e�A��)�0=�����$|Yd�,?^�e��F�=�a;��ʗF��ң��7:h��!P�<����,��i����K��5�Ѕ
��ʨy�e�j��%h��P~hu��6[�$�&) e���CuG��U�،1c� 	���2�!fud�"�H�0����qQ�7�Y[� B��%�6,z�΋�G����U�I'�HJ��ib�J�fÝx xh��$}YP<��O��#�Àt�(���ѝ6D9y���;)w�=+' �	���+�XRƈ�=$�u�DfX ��H�҉U�d���;Ҁ��Kk�1�M�/�VjV�	7/F���7e�+FϾ!�fH�&1��h����zU�R�l[#m�6PjӋɴ(I�������McTQ�Ikr9͓\Y8�K�q~�:V�΅7��l����fѾ��1�'����4�0�hp�3$8���]�a��JZx`C�ؑG�å`P2����'ǂ�H��ݮ �ЬŅ;wi$䂥Z�h)�"r��
����$�6i禭PD�H%c!,�
��D0�;Di�1-�:����^�<�dR�F��۪O��"7��!������H��Lidͭw
�0��i�p!�C�43K.��qg�C��(�;r��%��G(i2pő#?��1�r�ʣ^�$����T:�(1�c*�-}��,��|�Z��s铡<��-Њ�K%<��`;A�E!��dZ�F�1pqO0�zCo͚<U8Ł4'�^(��W��(1�ʨ�f��Q6瓓l�(붦���)v��at2)���'�v���*|Ce���,nX�� ��N �`  �WP�ѢFE�xO�,���.ç_��"*�Z����d�!�DΘ?G��16�����%X�䆧���3�͝��D��L"����8Êb��R�M���B|���V�J�Qf zC��*1�qaq�;�O�\���Q�|e�s� ��Ra��k�U�aDJ�"�z(��,����FY$B��
�.��CY��R���|�L���"j��D7pdQ�tg��}�D�#b����7�~��I7HH�8a!
2�F�p7l��-Ϙ|��D/�O�aS W���Yc��ru�l1�"O���Y7d� �p�	�.T�-�1"O8���c �Q������+M8��"O �Ä�(dLNe3ХȨE����"O���$_)V *R��\�Hq�"Oh����%_���tCP�K�J�u"O�� J�HS�-�p�{$Ԁ�"OQ��C���hA��Cȕx�"O�a�m�zVaI%��%#6���"OH­%O�<�CT�E�Tt��"O��8��F'T�i�J58��(P"O��s�@��y0l5 t� f��hj "O���1M0Y�l���Ιx�� a�"OP��u(ϰE`]H����3*S�"O�4ZՈ'1n�h�d�_���g"O�D���ڢS���q��xK[3"O�䓓����9}� x���x@��s��	��	�#���!P72F^�@�<Y���D�-s�DpA?x���N܀5�\�,��B�Y"�m�AҫC�����Y=<F">�q�>(6�hB%5�S�0�8iAD�.���r&Z�rf:B�/y���5F�Z�r`X"@[�F���	Xib ��J�&�S�O�b���#Y�:��@ �)g�Xh+�'��҂���H,�C"R�t���O� a�A���xǓ [��R��>����7-�&x�����	=DSN)�r�#]@�c�`\���𩌴$���
OT�Ґ"Ӎ@�&M3iR8Ff<T�I
RDL���_&jEq�~q�j��e9�!+r'I�V����"O��kփ&R|h�Q&�s6�)@E:Ob)PR%�b��!O�"~�`��97�,i1�ee:$��l�h�<)bn��%R)C&��M�P��w��O�Č:5�ƭ'�",O�+�`e���!f�*��b"O��X%��F���K����j�d���"O��aD�8$���8�R� h$"O���V��n�J��%�-H}�"Ot��Oջ#@�G+XaY�$@ "Oh-���L�4��Պ�iƆu5pT5"O��cs
��U*�����-@<��"O8��$�
m�}@c���FHtq"O�!�p.�2}V܄2��ؒ@X��"O�� C��bQJ��)
/���&"O�q�W���#A�Ȉ���$F�0q�"O��sQhf��j��#4ԼX��O'!�$#"�b�Q �܌yI��d�!��*�|���x�����%يc�!�D�!Ǥ�"`Ŏ^��R㖾.�!�+B����(�3w1je��1�!�V�6�fL��N�<�*�ZD��14�!����(�������-'��=�E�	_�!�$ſ1T��u�R	y��i�E�-�!��ѮV�J$+�ʜI�$�1g̍	�!�D�(#6	3�܃y�6�X#k��;U!�~���H�,X�hb
}��kU�\H!��U>�:Qn��n��03�# bQ!���+lBa-T�%*�,�W'r%�"O�r�I�[�qq˚�`�l�5"OV�񠆁�5��$�#�\�*e�"OF�Z%���t20pX4���^%q�"O|�BR���Y_>`7�0AZΙI�"O.0��ǹb���[@
9l:�(A��r<Ȫ&�I�`g�\j؊w�꼄�S�? �Mj�η18$ŐѨĘA52H�c"Ox8
T*�n�V�s��l���"O`�0e�	�/�x���F�^���"O���2
�Đ:�Ã�w�"�[P"O
�q�?(.m��a�*_̬�z""O~9`vJ�	�$ANɯK�%@�"Oʁ�h֞ip��Yld��lx"O��`W��[\VآD
> ,�`1"O���FGТ%���N�#�"OL�`��jA�h򮝯/��=A#"O��4��+9�����*R�*ِ$!�"O�SB�U���ȓi���!"O�����.ܬl
�.�^����t"O^IP���+��HH0�	����'�l0p�C1X�*�a��}"L����7U/�d�
��V����˦
aF�XEm��]��P#.�2Rz�\���mӪ�Z�K|�ƌá��6VjyqÒ?7-'?ͧV��`4$G�U�`�#��?��`U�� FB1O���.5�E��)�J��jB7r�b���y�J�r�`�~�	 %S܍��"J�V���Do��� Ot���f�	T��U��@M�SJ��a��ۨ	^$A#p`k�@3����fk��&�"~�#&L#y~� �,���-Z��X=c�0���N0�����	�eȟ'�����m�Dp��@B�}PqOdh(	çۈ��C��^��$	�D�<�=��$ "t��	,�v�W���o^TyQ�N�(��޾����=�)�?�>��UB/����4�ڲ�N�	-x혥?�)�'�@��W�U*U� A���3+�4�`-zD^��'��]�A?���XƎ^A~t0%ㆺ<�����Oe�����p�V�ZV��̺�K?�����/2���ꎆD����Q4���D��A'4�b��+"V9�lE���8��տq�B�e*�5�u�?����'✁Γ��bg8l`q��U�:� ���'w�o�,/Դ�'h�S��a�	v�	8]%l�ȜsFX�8Gd��E�i�b�xJ?�O���N_P�)�K��s�������� 1�`�h���LS���<6�eȒFI�ɍ9yn(À-⧘?A���|l�q)��@|pXp�M^R~���5����|���E��]����T�3Wx��W�8x+�ɏL�4ka��>Q	çk�>!�Gf�~ղ|� �ߚ<`�V�S�{eD�G�O��m���"�������`�2Ⴑ h�L�1k;
ec��@�*,��'�؉�W�@�Bh���#X��9��'A2�cT��A�mX�W1��:�'n��R��=m��K�.E�N�
�'�pPx7n�<g��B��[�I1��
�'�`��ı5�H� �J�!I$|�	�'�  z'�H?��J���Ѻ	�'粬�BT%:3�$�Ӣ���h
�'�4y��矒"�>�@����p�#	�'<�\	󠎺k���[�s�p�	�'�RF+��j
Q��p�r�'�x8��,ۤ~9�5�Df��l��Y��'ʂ�D�L�h�/U�g��t��'4ⱓ6鈟T�J�1���!Z�t�	�'֪ܩ���p������_1IK����'���g�* ұK��-:�t�H�'0��5�%?�`���[�B5���
�'�آ�+Y�y�������v=
�'J�
���4��e����
4��	�'���G��"��Q��1����	�'1�p�1�;8���i�̇�+�R�K	�'�,`�Ң)��{�F,7MR�`�'SXl
FkW�Q��Y1���/� q1�'������9\{ӏ�!"
��'^P�Ҡ�^-YE ���bؐ oC�']T��9u�A ��p�'�.I��ĭS����(�9EĄ�'k%9ъ�p9D��i�$�pq
��� �����&-]�Xɡ&ψ5��E`W"O��+ìW"�Аj�K�~���@"O���J�_<���)QK���c�"O��tB��O ���皚Y���A"O�S��5������(�z�"Op9qꅱ,���y�+��R%cv"O�Aa6D9����F+��D�D�U"O�+`@�B'��1V��z��M�"O����i�s�|���0��9��"OF4	��M &�P�+i؏%�VC�"O�xh��S!�XC��X��8�"OP[�&_1��@��/K�Z���"ODE�m�2c��GӲVp>
�"O�t� !��,f��)MUbN�+�"Ov�R��0��Xy�&˺ �R�b4"OĴ���	�x�$U��C��ԩbf"O�]1�f��퐈RԂ08�N��e"O�*�i��c��e�wBL��0�8$"O8��� �Y��TZ��x��H�"OH��V$,q<-z3�*W��]��"O>�xA��,X��@���]���xE"O����T2/,�9���2$�ly��"Oԉ�Pc'#��U��+&dԪ�"O�%jv.^��d�I"�*�3�"O ��cᘫ0{��2����\��"Op�	V��$����'옵a�rx��"O���æ����"�)g�ntB�"O�|���3A4�I���/����"O��Q0��$�h����Bw4��"O(�	NӁNh|��Ǒ%`�(�0"O  R&K �1� �J�t#@I��"O(��7<�4B�5��9Q"O�͸%�Db��Y��F�8�]��"O81ӤD�w'�5"�ʤT>��"O�-)6mK> Hir�[9B6�*w"O4dp�NC$�FXK\�8e���"O=;e�[�R�������G�|��"O�L;&�R�]ZQ�t&��=A��t"O��*WO/WH��6f�K@j (�"Oxm"N��gn���%��� 2"O ���:
�@�dW nb�:A"O�����xT䩫�$�ek&	q"O�r�D�dpq�s��1@hl0c"Oj3���k ���؄ ~<%��"Oz�x7��d�+p�-uiD��"O6�r�aϔ_m��xr*�Q|�Ų"O�a�Z/C�0t���ƬP]\���"O0�����+8X�9�@"���&"Ot���ꖂ��1��K?u|�'"O���K� 2D q�㋓50R�D��"O�!x ͈Lla�`+�1��`""O���"�	P����jM�T���"OT���3M"����o�#
f�c "O\���K����H��H2g�� d"O�i2E%�%@<Al<y��"OX�;��$��,�̘�H��岥"O���E�S��)b땡Dܦ�'"O��0�D33�,Xq�	I1q̈́+�"OHhK�<��Z���$Fv4��"O���@:��4���Q�b�P�""ODD(�	F�M�<�)��ځo3N�@"O ̣�ꎃ,9��!��
�#-�!��"O�|����PD&�i�ލ��*�"Oxx�R��4�B��B���F� �"O� ��f_�M��5�ӱ5*q�U"O&��f��,1���g���"Or� �g�$&�;���J��p� "O�C$IƪPm2E�6�џ=�(%�"OlmK�b�F}��P��_S���"O�mjg��m;� I�/ir,rt"OV�b��8E�J�J��g&�d"O^,A5�[��B����� Q���%"O�<�b�83/T�#S�3N>a �"O~�!P 4	�l��v�X�}/z��"OD����q�D�F�J�x�T�"Oe�E.�hp��<�*���"O�<*ǥ\1V����Ɉ0!��%J�"O�,c��\�RH�§K���p�"OV$��	�8유�h�+�Щ�"O��[-C2��욠��!g��-r�"O^���)�I�ܡ�7����NLJ"O�8�q�P1Pd� �<<��(1@"On��t��}C�`��Z�n�|�Hq"O$��� -NNT���5}��"O�8���_�,u���y�Qt"O�E��N�#�1s���)m�Ts�"O�l�6�/#�J3�3nY(�"Of!�p%� ��]���X�Ax�x�$"O@��Y\��+)��Vvd���"O��v)�{g�嚦Ȑ;[\���"O�8���Ҧ&�l��t�̊;W2$��"O�KƁCxH(��ޒ/\�-2b"O�tAZ�X��ݘ���"����"Ol����$���j�ž|����#"O0�S���1Q��I�F�j�\��E"OT:Da��p���],�c "O�Aq�P�,�b̢b&]3/�Y#�"Oɒ�/q5<m8�N�`Ԧ4��"O2��H!Efɋ$�̣Q(�lc�"Ob����Sz�dr���6&�(� �"O$Mp2J[�D��yi歒�k�ȫ�"OV�ٲ���Y[�}�"m	�XN����"O���u w=Y�큡I�j�"O�qお[:������P�d`���a"O�UQi��l1����BSB.�` "O&��%�T�%7�I�%����"Ov�ynĪ��Ij�CZ81�Z�"O��#p��;�"�����<
�8Xå"O�K�GǾ	�6e�fC�&����R"O����c��WPPDB9T�h�BA"O�1
A�2<��D#s�Z�^�j�l.D��1b�7j�H��@ύ�Wd�볎9D�<��/Y�4��aV/F+09�#D���#�L-�	���7��� � D��Q�	F+F�Tl�A���n,���է=D�x�Pf\-RC�mp��Y�$��$��+<D����E��������7�l��A6D�`R*M�6��|��n�V�J�+��.D���Fg�
�~\�$j��@b�@�,D�`y��T,�Ii�.X<��ru((D���!̔?.��[�V'}�Ԅs$�'D�0@���Hp��zKP#y_�|�*9D�Ĩ�jاNZ��׎ey�E�'6D���V
Ֆx5R}�M�,�����&D���q�LM6���ƩI7J~�{��&D��
�-$�V� �:xS�xp)$D�@{��N�/���F��m��� D��Y�lӭZ�v�����v�d"�F9D�� �kى`x�@�ᨊ$*���ZR"O���M)B����ʑ�z��P"O$4
��[CD6��C�W�q��\��"O�i���	%�Ȉ��QU���"O��
A�ު@�ƅwlY�"O$0S��w�4@óO����c"O�Q�s�l� �SbH���}��"Of��g$^�y�,9d�u+�(H��"O�� g��r����@|d��"Oȅ�fJ�~���
� H���"O�Y�(�2Q�����`��k�~��'"O�mrj�%^P�Z������U�V"O�I(�[��+!	)s\��#k�|�<���p��8��!9H����Er�<1#�I�WF�����#G䘜+�/Gu�<�v��-�"Q;��"�������r�<�4 �R�	�
��匠P �Wk�<�Q�	42�(���DE_�Dx���N�<�S���.��1���ٮeĠNO�<ATʽk��y�&�FR�<�ˈC�<��I%F��ո4r�)#bKEE�<�to§�$2$̅6y�N�
�@�u�<a�D� r� �@�i8If�yՍn�<q1E�1/p&���%�?[��T0�k�<���\�T��=ñF���-��`�R�<AN�j$Z���45۞4(���L�<A��B(YC�l3%�єn���!
�_�<	�h�]��Dɓ�Ҫt���D�<���Z�K��G�X���j��A�<iGH%%��y�ſn��밂�~�<���[)'4ɠÆ��L�:�*2�_y�<��E�7 ђ@����8E!*���O@�<	u�� 4D5��=1�$�� �Vy�<�I�3pC�����CD`���@�u�<�C�=4X�"���r��!��C�n�<���[.srHC�)ձ&�f�13o�n�<�W�G b��-�R�-�����AU�<���7�����V>zZls�"�P�<�$-G�j�(@�`Ď2s������r�<��CQ�E҄�@M-sS�кr��k�<�m�>��t�Se��<���V�A�<�
��i�`� ���"d�O|�<1��O�'@lCw�	�pUp$��@�<�� 8  ���^b!�=ry���w�2
�Paأ�ۡ!N!��έ?��q�Z�4�Ȅ"��-��G{ʟRt��Z�Ut����y�T�!%"OllS� =+��Dѓ�]�����"O��*���3���s�f�8y���"O��lQ�(���EA�"d���"OxĚ��ԺM�����=j� ���"O.`G띥��y��탢H�8xAC"O,��T�W�J��	@l�>�(� "OD��i] /m�E:�職´���"O�C�h_�V�TPh�XKP�p"O�e!F��Gf���eA���IR"O���iսXFl��aJ�w�L� "O�Ã��:ep	��l�"O����k!T������P��H3U"O�Y{�Aӧ���3�ti��'�qO�ɠ��p�V����k���3�"O�,�ѣ׬|z�����P�8���"O
� 0dQ�_w&�K�oO�;��;�"O��kV'��^������L9k����e�'�R�����*m4�$�6)G�?��݄�,������@��r�B�]Ԕ�ȓq&4�J��}p`TO�'A��a�ȓ�9ۤ�Z�BֲMxT� }�J���^��C��
�]�D�y��M�P���ȓ�&�)��u� )`A\�{�D���o�6e%_*o�!�SRA.��ȓU�fdB僃 ���Gт����_4ĕ3�Yl�Yx�ּI�vh��>��x��

����Nߑl��I��Iay�.��2�@L 2�ր���F�O��C�	�L.�"d�1�μ�ҡ,��C�ɞ���;E��i˨�eV�ADB�I�E�L� �e߀+e�D��MR6HB�ɹ��C%�ǘ%x"t��ᏫU�4B�)5D�,jKU2NX�sT�͆e�pB䉎xT�H��]5U�* H ���|�4B�Il`L;$G�_Z* 2�#���(B䉮4\���պ`�6��w��!� B�	#|����@ɴL[F0���,S�B�ɯl�4@�����
D:u͢B�>�<Q�2�M�C�����H��>��O��>9s0E��h]�y�FR�RP�AW�,D��Bt%�.c(��i��e���#Q-+D����o��,��0-�7���x1D.D��#R�̕B~�}����J�`�H6D�ȋeew趗�EG�u�p�۫K�!�d�2*�x��d홥w'T��j�]�!�� L�Ā�oɛ��@�H�!�G�l�쀛ᇑ�n�<��P/U�Qz!�Q�crPɣi��=�r��	@oaz2$0�D�O���&�c�Yx�쓞 n���L�\�<���@��t�h�h%���1M�Y̓SP�lFx��� �� _�TKH<{��G	܂("O������<:�z��G���G��h�"O,D�'J�*D�x2/\�vԄ�0"O(ۤ.�$1r���d��WaV|�V"Of�@���#c��0�B���4���'�&�~�k��5�!�&��|��C�I�8}�f��0�"���H_5:,|B�	�e��ɅD�(L������7+��B�i����c��B>L��NO�7�~B䉠ՠP2��O
��ص�L�k� B�	� >��E%K)c���t�lؐB�I�j���kä
�@��1��`��d��Ī>�c敻#A� ��GW�
�*Iâ��G�<q�,��h�tqI��F)px��3ŤVY�'ax����{ ��2g�_��-���ܙ�y�	�}/ܙ($hǲO���Ar���y��	7~�e�աK�>��Dl��HO��=���?9 �=�!C���6L��kdg�<��Q:eɮ��b"�((�.��)�`�<Ac˄K:>L�cg�<o��@��u�<�"9��)�ק:{M���L�<��͒lXn���FO��jI�E�<��Ζ�tKU��g�xfj�(�]�<qU)R�n���oGll�I�)�t�'?A���	y�EZr"��$fMAV�:D���tʏ�~��h� A�$�V�Gg3D��hDO5[a���#�%@"C�4D��X�KN��%G�5>LJ%ȐH	 H�!��\�dM����h���vG�3/���"N�H R�ܔzT�8�B���y	ݦ_����r�f��K7�y�)�'����*�,Ը�'[%QtT�ȓN��p0AB� w�Z�O�rѢ��ȓ!�Z� Ԟ|�2 �4hŞ)�x��=����ӭK���w%l8�ȓ/�X�$�.�(-��m�&~�)G|R�S��D��'�N5Z4��qzC�	�}�Z�������� ��+F^$>C�I��n�P!�Ľ�hJv��cvB�I+x���d�B�Vݰ遴�1*�x�IB�����.ɫ.֚	�G��c�$w":D���u/�������[����rk7D���3�B-)��Xxr��6$D]��i)D��M�!i2\{�ŏE�J���()D�,P3˾ p��q�[�h5���9D��J�n��p�9�Ŧ��F/�l�D8D�`�3�04AV��ң�,|�"J7D�tY"d.Z�64�U�UZ-�wD(D��g�߄[��p7怈 aZ��#D��9�L��|�a���СZ�`!�"�;D��1O�"U��8'�6+Uj�"6�6D���Ɨ�S�41��&,[�� D�,�c&��԰�Ϝ03���+$D��c�'Ɣk$6�1�L�/��}�bG#D�8����_Z&�r䭚�e�v�;�.D�Xgϋ7�py���T7^�U�-D�8(%
#	Ѩ�"� Q�`}�D��C*D�iT
)Fv�P32j1fH��Ҭ-D�ġ�OH�M~�!��i_�l�(#��+D�X�ЉG:#i:�sC��"/�]j� +D�����נk����F��<F�p�a�)D��x���8 �PuN^�a������2D�8SGw�e���\*h�q�*D�(1@*&������El�
u�u�$D��  ��m��`�.��1��  u𥹐"O�q@��PI�lce/�z[����"O�\Ǥ^�nx*r��eRf��W"O���%ԧS�A���@�-�&"O|9�pIQ){��xJЈ��X�!V"O<Phd����eZ3�%!�Bu��"O�1Da��+,��q6'>".�k�"Oh���+�#F��1��%�<W
hL3�"O�ຕ�<iĪ-�e_/���"O���Q
�nlj|c�Â(J��P�"O��*��Ȏ�SA�/�fq��"OYCUGw��Mq����u>93"OT`��Ҟy2��T�-U��85"Ol��7� � ܩ��A*2BĲv"Oxh��χ2v����$҃M�d�j�"O��R��7}�����Q�.љt"O@�5a)�B�3�
���A"O2!p�T'��ذ��|X񓋎�yb&Ƭ4w*5t3Gj���n�$�y
�5U�����b>A2$xS����y�ᛶn���cU�7:�[�
#�y�jD 4.�TI@���y�����yrKZ<�S�oX�n���T��y2)��>��c�IY!z����b	��y"�ڴ��� `��n�(L��K^�yB���Q,b�g��hǈ��D�y∋'6�J��sC�n��m �h2�y�`ǘ���C���~�����1�y� 	� `��%�<@�d2��>�yB,� vN8�`�n	�P��&خ�y"�.'�Us��6e?� �!����yB��2��E��@eس!)U?�y�b,�콻�I$w_~���J�y����,��4bbI�%o)`����'�y_�l��)KW/�B�ř7��0�y�@����h���<0C��
�y%�@0A�R��E������;�y��2]^ţ�$=/�%� fA��y�_�wL!�'ؽ:�nXYe"[��y�E��j�RI�UOР7���qJ���y�hӚv^��E��6g~{�l_;�yRf�@I\�(���(�hq����'�v𩒁�z�OŞ�HFW5C�X��l�w�|���'V␘���n�B�����i��TE�	z.��N�H7�<�U�Ҍ�^�xV�U�>(åc�bh<��ΜkDB�ʁM�S_���E�4n!������Rp!�(lO~p�r%0���#�)U�
��b��'1r!��+Z0-��]��م�N�>Zn;�Ӛǲ90��9D�h�X�J��`�"��U3,�a�;�d�m�l@j�D�7$�kc	8�'?�R���5�Ψ�p�C�fd݆�!��zE#�]��h�c�C!�\���[�S3u�ŏΖ:�:2|�g�ɶrZU����9��陕��i�&B�ɹ�vd��k��f�.�`�#xG� �b����8�S���-�W�'��%�u)U>MŜ�c��#��I
�K��}���v#r0��N��i��RQ�=�c�D�Y�j��3g����x�o)\��ɫ)ǲ)�H�3�ˋ��$��g$^d���[��j��<{6"�?Qa�)ܠf��u)O�g�p�1�5D����ͫ@cj�C��ȗaC����>�R����v͎|v��0J�c>y%�Tb�"F�x��6��0'e�4��K,�Pz��F[c��x�Ɵ�(���O�9�&�b��9�I#{]�p��I`�V%�! !DXsb� !.����$��(� !X�B�]��K��p��,�� ��Ua�ޢ}sR(7�q�����ji�0��<B���yL%p�/��4��'�2�b�$&p�[�&؛C����#�IٙF��0�'P6ҁ	�hҨ���#JRz́Q��C�,��=���� hX���r��;���36�2%��Aa�)>���_=gj�ɘ����2A�8���c�'Z:�`���ZF��B,9=TP!�yҢ��<7Z\E~���?���%��dS�CPA�'Pi��I�#Y���eO��P��?��4�I�`[�k!K�|�) V�p	)������Z���8U�7�m��hT��H�ڼ����(k��h���؉Po�<�dY'>�~p���A����8�fJ�JC�e�S�6	:�	Se���D	�_X��a���U�>���^=F��'��m�Ö<y�1��^4�O�5b��Vk��HT0��	�(ʒv[<��!fʲK�V�PSAZ�B��➠�P͍��ħ`Ҁl���c8@q�`
\�h!v���x$�#�#�O��Վȗaшt����>f3V))G P�X冖��56�	�� E����`�[�bѪи'2�=a��'7ҩ�� �(�l�2��N9b�j�:���	��&�H��D�)`Eƅ�� �+�`�1b-ը�����Z�0L�ѣ�s늹!@��r����w�� �J>��ʦ�.�l|��Rr�,h�+�D����]} I7��S��3DP>��$�DI�G	..:V��@4T��';P�+r��P�����|��'Q��R��M�M̺|�pE?2����E0��I1L
�X���A B.�����ôh!Ȕ��'�DH2�ȡ(�(`a�� I㊝b@mӤdŗ�j.(�*`ɜ�WT��@�˓EQti�^c�D��נ�4_�8�k��T��ĭ��'�
�� ��}h�(�� ?L�d�/�ƙ��Ǝ��X ��2hH����\{e�b0!;H �6$@/�^��,d�>�e���H'~��R�'�6�!���O(`���͔ �<�˥�R �~�bt/$p0�a9Zw4) ��E��D8�F4���GR�v��>AV쓱�hI
�"@�3�����l�ɟ1��ݰR�D�c�$5#@I�C,�	h�-^��R�oQ��P���kiP�QU�0y�Ւ�eK�q������=�g�Ϡ$<���B��a䶐0�\+|J�822ß*�t�)6�K� �΍�$�"!1�ɑ�V�e㺀h��3(B71^�ڶ-��N�4�9��Qqh<�戙=@��р�Ś�q*>q0LO.V�����Z]�19�"2���
�H�<D���e%�t#,Ux�l�R���C� O�d�y�V��i	�a��$�4��<�fl�j�M�wę�S�x毘�����,L��!�I��{��͒A��>K��t��%���'�e�^{�'�Pq��F�l��Q �-!3�!�N>a�Y�";��f�Ԓq�pt�&���r�c]!n�J%	g�	�]|!��-�: �8hcb'@/\����A%�#l��}�6�v�Z�NZ�/5�
�g;8	Ë�+R�ᐢ�ЬG��Y�Ð�yr�[*<�"���y��ǡ�@�Y͔+u-�T
�	!��x��B�R����пj�n,�G�	F�:0�1�E�K�ƃM|J�0i�D�� <m�p�d��A�$�D[�Y��#����t����`��yC�ɀ@�'�f��)�u��#,FAc�ץ[+"L(��@�N�� շ`da�E�uW豄.
�*X�=a�@�IV5F�Ќ=x���ʔv�I�?v��A*U�N�Ya��0g;���!F����:[l���G�+��y����g$��cEW�v��
�c�]�P@�[�h�K�A��?'�)h�@��

~�5->�E���߃e�G�\�r����<!��;9��d�ن}�j���j\���^�f1
��?9Q<�p�MY�Eni��(�!bL���Iuڒu*�W�o�l-J�ٽ?^"�(W�$Ht]�6�'����ǹ�H�"6�[:M�r����@�����K�l����"H��Ɂ��e�څP��űK��t�����!�J��B ô�U��q퉙w�	 �a�{0�lRee�E��b�dJ%�N�A���уvH���#�RY��)�n�d1Zt��*�18f%�G�@�A�mB��2����>	��Nz���B߉k�4ВS�,������9o.���®?��r �ަ9 ߴ{,��� K�2��nW;ks��A�W�-���d
H�n���D�p��U��T
'{@T@!,�+2f�PW��/D7-�Ȧ���\1�)Z�%�V&��i��D3?��h�5�'Hf�G`Fa7<Là�ֵ"�� �ϓa46P� �7$��<�t��xN���o�#NV�(��]���������4�H�Y��e�I��h˘OA��is�I�%e�+3�_�!ԅ+�b��|��OЕ�BD�q� �&_95��Q࢜;5'L$�0�}�T�B�<>,� �Y�W����K��I$�=��CNx��j0]%}�$A
��y`w�L. �i��@2J:|�@i_�r����'6�C�:�à�ۼ��Ƃ�UZ�3h�m�����x�R$ ˖�ȳ��_.�����\�6aB����<�Ųi�0���K�#a�ژ:�F���aЏ�Q�	�ƽ�1dE�&l�k*Pj���ܘ���[�N�:���`�!(w-Αk�,�H�l=�0�f �q�[�L;��@�����=)v@6�hO�Ԃ����^f�ba� �T��٢�|r�@9W���r����@���3ua	*%��a$9q� J�%�q��($ڏI�XtʣG"WXń���*�x�g�9Z(�a��s�PH9�
�`t<�1AD�(��cwHĕ�47��u%*�h��C2r��̻
s��!�.��t�O�k�0I��c��/H�%�wS �Z�Ӄe��,���Ҧ��@��!Q��Q@L`*�#R_��8*E��%�y��S6�V!g�[j�H�KP���p=��@�V�h�7� �H�F�(��;i����ԃ> @E���RG����i�K2&��ӠU�L2 �P�	<�f�ҲȝVu0͹w%$4�Z�ԛ��Re �����WzO���s�?.�6�q&�i�p�����)U�ˑ�%�D��(F��̃��'�+��x��B�D�K `�`쁲4����7n���^��� 8�0C۴?���� ��u'#]��� $RdlP5��Vo���&T@"OjUQ�K�;m�L�"o(_v�y��`��m��'�����@�jQI���>f�`�ЪZh��'���0 ��V�A������:�u�f�ڥ���u�ܡ[fk<+���X�.�,$sLy���ʾIPb���J	@�<�
��յ ��DE��'S��;@��o��\�T��!� �X�}�
H94XP���X��j�E�)���;�O�����6@0x�zGA8(J҈9FY��!�\���匲({�0�&B�Laƕh`oٰ8[��rg_�Ua:x�D��	�y�eL���ilށ#�l��4�䀇��(��TsB�8D�(��I $��aJ����f��C�[�k��x�8O��9f`̽5�瓀%��qj� H���_.����##��񠰏�sΦ��J^�1����Ol�@�D�cQz�`"�ƈ:T���elL�L� v%G' h��S�/<ON��X�V����ү�Qja��	/�������}�v�r�H�~��d�/Sp�P{TH�[i��Ҵi�h�<�"� 8~����]�;��9��L�qy��Vu�⨻��S2�����6U)�����4�	�B�l�<Q��K�w�8�;%�������A7����'7@)9�����Ϙ'�a7�C(z��{E��`�
�'в�+������E�R�S#
cp�tM͟sy�p�!/=�Ou���=�d@)��^�T֔�Y"O:�C�[7�{B��l{�]�"O���tC�s����&�k�%Y�"O@A���s%Fdh�tY��؂"Oy �b/�Y���^�4ễ"O�,b�B�$v����cޏb�敻S"O�����>��-�#N����"OTI�ă�F\r���3�.)"�"O<8���>���y��7HŘ�q�"O�E�@ӜKH����')[�a`"OX@A�,pp<Xe��]�"8H"Oę0OT��=+��@��=K�"O��KF�b��|S�ӭ�I1�"O>�B�k��X���%߀C'T4B�"OT�h�@T2��cdoɑf4���"O���q& �r�P��X-n��ja"Of8�N�a0I���ōb��8 v"O>HY�b�0>�-H���2R.�z�"O��z��I�2ϐ���^ 5�ʡ��"O<�"ᯋ�4+� ��!�
���["O���Wo�=W�T�֯B��D�"O~�`�j�b��4Rr�]��$	i�"O6�R$hLǜȸ��F���Ԫd"O���D���fMK5����P#[�<�S(�QcLvd�.q ŀ��i�<QG+C?J���s�쁲B���Xs�<YQ�;NҊ`� ��^U0���"LA�<Yg�b⤣�V-yD>,�CA�<�ìX>��7�[�"f<=7��B�<9�$�,d4\��E:��UDm�<i�F����Ga�7E�R�S��v�< AETt�^(E������p�<�`ѣR�`PLгf����o�<���XH*f[.hC���tn�@�<��̛�b�,��b���0��8i��T�<�!oF�f�t=RҬ�?Z�d��XN�<�G �<.����^VR��3r$�J�<yD!ȡk��H � $~е��fLD�<Y���:_m�U�äƂe�t��]C�<a'H���l��D>;�Zgi
}�<y�@>`�����5B���h��y�<�EA�'��Qq1`ÿ=��(��u�<实�Jo2,A`���@��1tl�p�<ٵ�ȭ�^0 ֟Z[�%����W�<a��R�7,��ڙ^��;7i
v�<AĈ��.m�LY�iW-/�nQ�$Pz�<� P��b�5�2X#j_6p�9�"O�<�@	3f�С��U=:�䓅"Of��!i��o��%�݊t�FU��"Oȁ@7�%U(� �+ɤuf�is"O.Aɦi�)w�.y�3J�%w�4�"O u� f�3p8��P��K<��@d"O*=Z%��j@�̙ը
�T��Pq"O<$��K�G��5y�ƌ�yA�"O��T%�]��0sc�Q�`�ĩ�E"O���uI]�D��!�qeӫy=�"O�����&����2f,H���S�<	&��-:V��eR�0�\8�$-�E�<!��сet��Q�P6<0l�㲨GC�<y�ΓCl�rצ�'����G�<�b���FX�=�HD���PG�<!b#7�����*[p��t����B�<Ag�ۊ �&�85�*`_n���A�<����D��@�q,�/9���7��P�<-�(q�e�z;����F�J{f��=�Y�pF<^Fs�
�9��Ɇ�#��Ǫ�w�����+'N&(�� ��(��
�U��P�#GI0 ��h 6A�V�B�ȳ��J�\^�T�ȓ��h2"�0&\�C���
Gک�ȓC��A�bE�8��m��#Y)t�ȓ@�$��vDK�
��,��� $o���ȓ[S��l��lr��P����D��VR� 7
6��m������ȓ~��,SN�򨊁DCJ5`)��_u�yf�?���i�@��j�"Ot��qA��p�X�R�I@Ct���"O`#�6<�8�U�?F���"OHwI�N|!kwhۦ�F=Y$"OԜ"bO��Z$ ��aK����A�"O��0�B�T��B��E�U^��@"OF<�$�:P�0I�s'��ER�"O�HI5�J�^�:]��!&#�=�Q"OJظ�������4-AH�"OZ�8�H�

��O �6�N�9�"Od}2s`�A}%�Ύ�k�͛�"O�R��N�8!h8
f�3<|�Tkp"O�s�i����IwlS�T��
S"O����F�-j�9�
[�M@q�"O����Z�>
���HT���8�7"O��XBe�9�oҵ]1ΐy5#D�|�RKJ��T�Dν4.��7a5D���W��((��!��M	������#1D�����Y'B'Xm(�(ĥ��LP�,D��s��AT%�e�D3yIȤ3@�(D����@E�"�!��c� ���3`3D�$˓��O�̸)���<c��r�'/D���
*x�xHzL��q$1D���'��kֺ�S��J9NM�҃1D���C�F$x#�o�T�Lq�֬,D����[c 1qτ��� 
#�yo�u�F9���\�vb}(2Ǎ��yrO1�pWi]4J$�����y��	3i��Z���#кM���]��y,C1$�ɷ���>���カ�y"�[���B"�)\�A���y�iO O�����ν/
|R&�%�y2�ܔo�ړ䛾� C��["�y�Ε�W�RpQ�B�

vֈX#��<�y¤�'|��ZщգxĜLc`�M��y
� t���*F�BK�Dk��T�B�֥��"O�@�BG_"8�C1�2_��a�"Od1H���!����U��"y�dڧ
O ���
�ڄB��\�]��5�2��#��P���(%
���d��.�u���ҲN��cb	@�ax�'D��%P�.��N�&X [��Z2J	\����B�7c�Q�ȓ��a��Y� �`�✛*~��'�`���C��ph���GA>i?}	C�F#t�JU�֫X/6����#D��#b�39����+6S��8'O�.9%!�͟X�V�RC�	p����Oh{�O6`��`��`�dY����,J��$�� �~�'J��4�v ^�m��t
W.
a=
bJS�UG����a��D�bŚpF#��=A�dqƽ�f�)�P�QQ�H>@ Q�;Po���*�|�0"O:r��@����(< Z4���i�9:!GT�C�y��ڵ	:��%D�t!T�Y�K=��P�Fy�cAC��]���X��a��Q1Xy��I;��0E��D�S����yG@Β�`��`�I�<6�(��Ik4�h�D��QT��4@��A<V#Эґ���#O����n��C��+E�����cB>I��ʧt�~b�|��7&��!7�q��p�+)�$w��8r��%�mS`�]��g�\@�9��/V�F:P�c�!75`��$A(H=|y�A�69;^4J3ÀF؞H9'���;-
e��f�*3H��E�v���c�Q$8hPlZ	2��Y���RzD(����X|�xs��+�k���t�
���B�%�6�
ǨN$Y��D�~Zn@[�& ��Q��M�,�����Ƿpf
����Z �ʨA:�iف�\�\���-�5��Bc_y�]H�G��d%��፜(;x!Cϓe!��Q-]�/4f'X�2��(�1I3���ו �A�1��|�4�D�P�}�daqb�
:�ר�0K7c�4��/� �,� ���	KnL��"���
L|`rg��(�)��!��5��$F�rx:�"��;^P ����ՔP�p��T�AZ�N���e)[�TQ9%o�{��x(0�� ^�dM���'R|܍a�B��5�u,�/F�a�g�v�6d@�Y�X�zq���QzԉqW�c��A`.�~m���1 ֱ���44�`SAH��Xr�C�ӸT�]���O�xl��8&<�{�,Q� ��P!膔]y�س":P�y�q���jH�e�)<�ɩ�GV�8bbd;B�gx�̱����<ktPC�åUW��Ҵ���2$�T�N�8�T	3��
Lg����M��IN�8�3�T�tT����ޑ�L�,ё-�&`h�⒠,,p:D%��R�.*Pr���h�)���C`#4=�A$E�Jx����=odM�!cR�e�������6 �&4.=��	�/$��t�Zy˲t��A��=G�h���øNض�g���踉ӄ�'(	:�	�ǤP����?@���{�@�Z%(�dȅ�2�Q4�
C㉈sn�i21J��E� <{H^x��awf�'���͓F�(��
qh�Mj���B� ��C�Yw����a��x�H0(�p�@��W��ч��0*�~,��CJ�P���cցZ���5�4�<YX$�*@��2�P/ۀM\D��u�.e� �!L3	�Ќ��,�"�AuCC+{���I&
S"C��'���q�j�D�����̃�S8*����b�.Γ�p��B"�u֬�(f�X�v�`]A�>(/�<j'�:�Ol��C(J��� �X�)�,�R��ǝ-� ��ԫ݊v��«C-0�v�͓M�ޥhG,��*� �j>�̻�'��ܴk�*\10x��SO�ܒ� _�|)�b�*�.L����.Lk���'-�y��*}lٺd恛T�@Q&\,�4x�gA����·qrP�ظ.%���1<Opp�G�:*.��hо^R� a׋�&���+��<N����r�\z1�=%F@��DI�)�('k@e�'�XP��p^��h���GF�i�� �'@Q6�a�
ʻ(B��7yuȺS�b�2�1R+ٗ#�v�k�a�_@�\Yc
�$��Qq������>�e��i�Xљ�7s�Z��!��_Ϩ��f*TnLKI��>�(���馍�۴��aZ��F0E�nܜ8 ����(~�f�S�$��B\��$�.��0��-4' ��SKGMO>�[@?�7��Ħ��B�J6�P�f��`�Ψ�k��"*�D�'ΖxE��,=Z:D�.��K���<ٓ���tDR��+@��Dze'�{��k0�)-�����kD4pby`�N; r���	:m�Xp+���tў��!'�(�B	'ƑR�����!�dƐQ����3(@�}\����W| Qk�(8��I�VS�4���
/"|��!W���y��H(����I���9����6W$��YPLɇ���`I]�m"�Q�"
ʎP�@��?�y|�RT��`�VM�;{�<�D'b����l�P�A�ƓF^��j����e�\�!��H)�)TeݮU��I�M�W� 8����Ej >����A��L��H�O�H7���4hC��	�A����<�p�����=x��.�l�c��-��-��cT�A	R�8Ab�Qȩ�*�-6X�bd�
)LCa�*�ў��Uc\2?���e�
��ػ�N>�D�>����0��X8ܙY��-_��� �N>��7M;�eN�%�^���^�\p�PccLZ�v���c��Kx���.�BP��)]� l��h��{�h��9�̙����%M��-��yӚ��cR8W;(�T��;'�^4"ɔ��bm�����o�<9�,Kz��@P�FC	(�F�!e�+EǠ@�犎Ħa8!�Y�>�z�
UY�-�F��P��_��ҳ*W��yh��G=
8[��J�p�B �g���p=��6��e����# � �8�֝m�����탋�wn@%np�v�*� �� n�x�
�@�����8 �Oҏ0�JMzcm�_�qO"��F�O-uW(X�%�z�`�9�
nH��B�4fYecޞr; 5
 (�Fyx�U1��!�YW���Ь5�p�!����8���e�)
� d� ��UTb��q/B�\[��nZ�o���
�Ϻ㇁e�u#�Y��
!��$=̰m���,D�H����' �\��!����XX@c�	��L�=O D���;HȀN&�J�YRAA6
��d �O��GJDuI�z2�)O	N ��'��
2� � c]��&H��KǾ=��tUbM��0<��C'=�f��%U,Ĕ��3��O�q)u�+P�x2��8a�X�d�ظ(�0Œ�E�	�NtQ)=5閝�Y�p+��)�z1ܾ��	��`�nC�ɼC�,�!T`Ь�����͖�4�I�N�I�M�:c��c@�I�@ �T�a��SҼ�EcȎ�b��w ��}p6/r�<���&�Z���3�B�sG	�/�`�PLu���lE�ro�ͧ'�\1�lG.0ȉ'"h`ò�6Y愍0���vF�y�	�~�a�!�Тx���O�7�0��t���@���:#���� 8��J��d����Ē�8�� ��.P�`��HKRL��cf���aTę.t�\[%�ړ`q�u\q;ІͭE5*��2.J����O�Z�����fw4��I�2�0<�'Ҝ��(�'6�|����3��$.*�Aa�92�	Rw�)^�0��ȓ|��A`ɕ9M&\[0I"I�\��'ZX~� R F>�H����y�nO7�3`bďfL�	�"��Px��9$��qa�Uʌ:��+2F�8�,T���Y�^%��HEP�N�څ�&�M�~�!�D[�f�,�gT�M�Bı�(	6�!�$_8y����E�Zz��6��a�!�E1Q��%31�H/^u���©��V!�Dܧd�L9�HؙV���Z�BeY�'�0�{E��=Pk`�XB� ���0��'����F|aE�ف%�P�xu,X��yRf�AR��h��8'��� G�S��y��C:'X���c 8M|�Yx#���yR�_9=�����8����p�X��y"��+L��&Q%�DВ�*�ybiL�/kz��4* ����sG���y���l5�Si��{��tX�i��y��$8�Ah�Ό�g��i���y2.G�Y�h�Fk�f!�]��IZ��y����}[Rء��Ѿ
��X@�&�y��E�:��Q�nєt�T��/�?�y��8d��D�EBb_�]�T ���yB��\��[g.L�f_$ɪ�f��y���=|�`���K傔�Ʃǫ�y"�\�N�ڴ�6 �W<IW'�!�yr͋�!�nH)w	PL�~�a�J�yR�K�(��%��ÆO��1A�0�yR�A�����X�.��!��yR�MMR�P�g��Ԣ�J [��yrI��i@�PS!#�[X��AX��y�ܢ59�({G���H��J�����yBK_�=PTM��mߐr����_��y�°i�da��Ibq�᷀��y�ަdGf�򒈅�v���1ĂT�yRL�!�P �V�?�J��.^��yb��(�L٢3^1 ���g̹�y2d���\-:��4dmxUP3���y���pXU8T��Q r8Jb�9�y��Dz�iѣ�Q׼$���y�M��D���q2��%�y�q��6�y"�\0E�$�ǌ�5+[8,3A��0�y2�=f0��xP�V'0�X��$��yBIO�2Qi7$�zA���y��ׂ8�)�4m,bi��z��!�y�
ܱcH$��â�,�����
��ybC�����ɨ
��0�C�y
� ��S�
S��(@c4 ܾb����"O��
��9�lt�'�Z����B�"O�DI�Ռr��X�p�2Y�6x@�"O�#�%P��@$y�횽�9�"O(�sc�8���%Iæ�(T��"O�e����?.��0���O�BuJq"O|��s�ȥ0�.����7���*O<�`%�}#��8�?K-:�' Ը�B^�E3 �
�� �(��
�'鶀p�-9X�>�IQ`Η j�L�'ir��Ëp�#��
���l��'r�g-�*,�(˖�Q��.�		�'&88��Yf���;#B�Ie��I�'DRp$Z�� �҇�0F�|�k�'.���J��;R��j[v�!�'^@�A�, 4N��@Tr2�ȃ
�'gu�q��Za�ek�+�kq<�	�'��!2 iЃZ뜝�ҏ���q
�'�>|���HVX����
#�|�;	�'g����`Y�d��Ђpm۩�x�x	�'x~t��jB�A�4����y�J,�'vt(WKr\v���ٗ��yRG��s�^q�U-6@R �Q���%�y��WF��$�8n*X�H��yb�T"��5�Bn�E=d�@�i��yBL����(GBڢETR���k�yҤ�6�@؋��SjL�;U�Q��y�O9:`{׏ˤz��4E�y2B"y0�DaD�L0E���Z�y��T�\�0IRE[�	FH��`���y���8GBl*��=Ux4�Em�;,|\ȉc�f?�҃q��Ê�4�OY�i]� x��G�U<4;,L�R8zX�х�<Y��00�H��I>��SM�jI�dp� F{|�@�G[M?A�ó1��S�x����O��ۡCK���	X�B-z�J� �;;��"k� e�*�S��|Zw�$�W!�3����Bt"��Ip��`b��A��ا�	�4'���0UM4'�5eG�:�O@]����{>)�t�{y���ɔL`v�{�N/�$ҩ'���z疟�A�*�ӳ]�,�jB��2Y� %aT�ԷU���	�:���	Ic�)ڧ*
AZ֦�+o7 j4�(>2�m�H��6�M�S�OڸxXv˱H� (񓁝B�Y[���Ǧe�<���OʱO��&r��}�g .��S��#��6�X>��	�:ٌʊ���uW��T���eA�4Y6����۶mt�1i�h�ߴ�ēK��d�"�Η-6T*q3u`��}I2�!1<O~�jS�R��M�K<E��C3(8@1��u����@�a?ƅ8��C�c?:(X�Oa����#]��Y[�b��i��MQ�JL�<�%,?�Dժ�>��O�P���$���K�n����D(%�ɍ�����������CӠ�°O�j���1�I���ɞ%��i�C�S≾��O���� �?R�cvG C���ٴb{>h�G�s��L�ȟr�{ta��UQ3�͂y%��rv�9Gt7@>*k"�dӞY%>�D�<��	K�H���ئ���&��	:�6�5��S�~y&��X���4�ħ$8����ǜS`��HW��Cze@��޾P�~�1�t��Գ ���,Y#c��,Y��#��"�m���53�l��%X�r)�h("��6o>1�O� �:@(E��� a �L1V�`}Q�-)�Pp�IP}ˋZ�L�ʧ�Δ!t �e⠩�g���<ņȓs����Ƚ��H���ԊE�E���ڭٲ������'���0�|��ȓ�0�g��TN�Xa�C�+���ȓ2�(Kqe�F���!�KF)m��I��v.�e9��,���8"���z��ȓU0�H�ׄ�$@�� �,htm��*&�!�9�0
@�?려���� 6�K	,�R�^�����*�� �S���w^�9$ǀ\1⤇ȓv�*��Ec�~j���^R�E��S�? �U �CC�i������<{8�"O`���bW�7��u���&O�E�p"O���� �j�0<� ��g=fPi�"O�8f,ڌz�J԰�8c7n��u"O$5j�����Ph��	�'&h���"O� H�a�w��|9��.&�q�"OP��4�^�z����!�����zQ"O "N��rl� g
Dl��Mc�"O�L!�땑 �N�9�RBu̽�"O|��+�tr�Ň�=�$[�"O��`c�7Y���ȁG�KT�y�$"O||�Cj��_�vX�T�M4k5V��"OV����Q�j�֡v@�,AP���"O�i��h��n�4�j�PZ�V�:&"Of����
>T� H��O� 7�2l@�"O�d-ı)Q��ʔ �kV֔ku"O
�+�B9%`<Uq��Q[V��"Ot�q��JBH�:��*uV�� "O��rC�3ep���cC ���"O��P�
��508��F@��X�"O$щ��P R�k2�UF��B`"O-:��Z�5�֐�B�cҜ��"O,�ۅ�	8P�i�W� !w����"O��r#L53�>En�8D�А�w"O�(C��k�Z`�٪:�j�[�"O��q-ɔd���K��C�2q#�"O��t��<��`�ˀP��z""O��rF,S�Hthk0����yɱ"O�B��f&HdK��5�f���"O��vg�<BДZ�䞬l��ՙ�"O�e�#eIu���4/�8C"Oj���ț5T�xU%�(
��u��"OJ�ǩD'a���:�I[q��h8�"O�,�3⍖Y�=�Į� ���j$*O�L9R/�a��[-aL&iB�'w�io�4Q�n���B�	���k�'�Z��D_d���E����#�'`i�g,�~S�
Vf�l�}��'���f%Dz׌���N�2E`�'ܸ0�7N�6t�fiةH�6HR�'�TP��^(���fԒF�����'�\�Ӏ�pkn�����-�HT�
�'���:E��Y-:�dFU�,��m�
�'g�����P-jTD�أ*(U�t��'��P�K�ar�b�gI�K�Fl��'������`��J��@+�'����î��y��� �MۀNܐ���'L^ ��`P�Йv(_+Ka�tC�'|&i㤂�"n�,��j��5)���'e�d�Q� l�$+
'�,]��'3��۱e\'N�xX������ܱ�'f�\@Wn�<=����7�׋����'���ZS�M'W���aT���ra��' �J����FCx��fa��f�~DC�'ά��+֧[{���
�t%��'LZd����;p��I �&I�'&%@`�>Y3��doB0���y�'����׫�*'��%q��]�xv��'�	�T!��L~�D�,�1j��T9�'!J���/��0������{n`�'
���a�w����r( ZG�ظ�',Vt�!!f�L��С�a��!��'["DBQ��&���i��#C����'���R�ÐZ\-[SH5��![��� ��*��ʸi���b%��L�\��"O|Y��� R��Uj�"V��� ��"OD�	�'�&,�S�	�K.��q�"O����(�8J3�޷!j��"O:�ʐ����`!�u�ްBzr<��"O���צ�8(hݺDaS:K}:x�@"O��1�9�D@�n	|T�mCp"OF���9F6FU�"CO7cq�Ġ"O�� k5���!Z�m f"O ����ۂOR�l���-!O�`
�"Orlw���ؔ.�yP���&"OX��"�
�hTR�f�C�
��W"Ot�Sfǖ.F0������5hl.�S"O����	n|��X��>��a�"O$�c�%ϣ%�3c�ݒE�8�3"O �{��X����E_�f��x��"Ol9�u�>/��PQ$*]�+����D"O*�Ɣ�b�����Q�u�m�a"O�����JD��&m[`�{"O���L��;�Z��$MQ�E��u�"O��S!R�ސ�Cؒ&���a�"O�O����ɍ�
�T�z�"Oh$���K*�8�I�Ar�P�w"OPT�b���Dx���}3x��"O�A�2�_,r�b�����E&=R"O6y�*��Hf-#2��?u�H!�"Oa�uO��z���{@�={�B���"O(�xf!�/���+TcbxkQ"O�T�XN<�8���,��9f"O�� T/ƪ.AZ𰈖-�V�"O�8ڧ�ќ9�8X�p�ُ���I�"O��"�$ЅSjЍ�V�S!6��=ˤ"O6(��1���㰇��t�^�"O�T�T��?���j%��	h�"OP�rã/vb�{W,P�M���"O�d���6#N�P%j9D��K�"O �[�%�<\e�t#�.ƌ�����"O L�2��J�-�%EJ鰀i�"Oz�`$���&��Ч�I��s"O���kͶ��pa��O�c��P�"OQ6ԃ����֌,�	�"O���稇�^6��{�G�r��L��"OZ��`��wh�mB�P?�"�"O(�H!D�?�L��n�$����"O� � 9g�
4o�5_�=�c"O�l��	B�aq��t(��b"O�T(V̓���Ѝ_6.i�q"O�Đa�|V�Z0��pu"Od=J�%�3�Ԥ��+S<+$� ��"O���2�ʨ�:�B�̟6e7��"OL�3�h��Q���uˆ�~�D�{�"O�m����@�� ���u�8�r5"O��� �S��T�	fq<8s�"O�a Ō(���8���F� �{�"Ov�2b%Ĉ	JL�Z&I�0(_��(�"Od� s� �j�㩄'f\� F"O�MZv��qQ<���{�H��"OtYk&��FM��@�1>x`�) "O�� �̈}H��#���P���y�"O�ɀ��a&�(8��H�&WQ����#�y��̛�?�������DE�<�rM��\��̚�a�&`���Unk�<�T�] 1-| ��F�,M��Ջg�<a⯒�td���'�  ���`�<� ������c�A
[4q�"O���6�.x���c�1�ޅ��"Oh�rB�E��<06�H�z
�yw"O �3A��i�����̪5�:S"O:���8����U��'�"�b�"O$��W�K!^T�¤Rh�*�z�"On !Iܪ=E���!���W"O��a���0w�(t�0�F=20@�D"Ov�Z� E?2�K���P���7"O���#+g����ҿA�TQ�"O� �w��3J�H��l����y��A'L��`�`a՟���� i��y�8a��w/��0J|Ys� �yr� E`vš�-��-��C�E��yr"���pSrm��)��1�Q���y2�X27�>e�����)�|�����y�J�5$c��K@!����B�y"�86�ٳd��+k�F�H����y��C�J䬭I���sjz1�p�U-�yR��D)�F	�T�*qk�Mǯ�y����X@I���Q���w�̷�y�#��H���Æ�S<|gz�wAƑ�y�;0�A�� x��U������y�#��T�������1���H3�y�GJ	,�u9P����+�:�y��\� ��f�]?Ij��� ��yrLБQ*�qɴk�qf�y�ǖ=�y¡?w�x���ey�t&���y"!��6���Y�)�4Y7��i��#�y��ش|ft�ȇ�ר��1����yB˞�oDL1r��D.c@b�Awꞇ�y�-[^F`�"�O� �!�N�<�yB�P�[����G�H�0� ��+�yK�p&d����Kj$�������y" �I������qf�I6DF�y2R�i4t
шM~/(�P�����y�]>:�^(� Ji�X��,�y2�[ :�><"�� c�vL8��;�y�B�;�v-j%LE�G^��͋��y���EzU��ʌx_���$�C��yR�^��D�UbY(s�D���
��y��G�m��
��5t�$y���y�i��<���cc
4\LZy��)G>�y��R����"���
��e �	_��yr@���|��؟3&������y�!����\��I�71iv����5�y�B��
�Dz����퓶�y��,r�nS ��֙x��ս�y�ߑlk(����܆Fy����y"̇ ��W�v�R�Rۛr�C�IJBԐ���=N+ĳ+�P�Kt"O,� �ɖ+>_�4�2>.��	��"O�,�w�
\���#�N�N��"O�$�J�I���W�Ge��{G"O�����S��8�p�O����0"OڔH"�R����PAHW"o<U�"O:��P�̙ZJH�ҧ�"�,u*5"O�!�����ĸ�G�@���	�"O�=��O�1s/� �Ɠ�J�� @q"O�X˥   ��     �  9  �  �+  �6  �@  �K  �V  �_  �i  Ku  \|  Ԃ  i�  ��  ��  :�  |�  ��   �  B�  ��  ��  
�  N�  ��  ��  >�  ��  %�  *�  � � V � ( �/ 16 u< �@  Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�� |d��"O
`�(�;���8���-0��1%"Oj4��ND^[��"3/9�0|H�"OB���H��*�ʞRy=a"O�味V�!X��!&F�:J�$���"O,��a
���C�Ą�M�"O,$3%o�-���p���+Ն�:1"O��ݢ1����`���y14]2��i�<�6��{_���c�H�`�fX�$Kn�<��A̼VI�xR[�)�Ć�pඤ�ȓA5��('nߡ4�� �)˩%� ���,��r�؊b#`T�eT09���ȓ!�b��g��}�8�F��-? �ȓ
K|m�ș�VṔ���2�%�ȓ"R�X�j�4JN�1�˘X�i����̹	_�jZ��1!g��zܶ��ȓgil,*�J�
j�Ne��i�J%b���f	�(U��:���G��$Y^م�~r�� S�%T"���k\�jx�ȓ|4�1�îJb��@ӵ�ݩn�V��/[`�"�v4�R�!ʎ<��M�ȓ`:��z�ؚh�J�Z��$HY:	��H��p�m�C1��!��B:��0��EnjZA V;9����J[
2���	��4'J�EA�IVW&��~�(aZ��ӹ�>� o�Y�|�ȓ�f�A�
Ο7�H��M�$�����mޠP����/���ANXo*�ȓTv�����{ ��-7�*h��I��sB�8�8���3����ȓNe*M�悡;������X�o��!�ȓ'lj�#F�m�+R&;�|��2)n�C��0S4���T:
b���:�0!��e֊��)��ͷV��,�ȓ0�&�8#���� ع�L�����;�P�AFd���,w�6d��r�EQ�( �gVlɦ�M,H��,DP���|�I	$G#\���ȓ"�)���E�B	yt&B�^�LɅ�4�� ��eëF�ڙ��n��R�p�ȓp`@}bŇ�=�$�AUN��P�����xyB�1&0��5������yr+L1�����L�?�H�[ǃ�(O�=�O��<��hçc��xH2,S(�\D��'�X�+UʜP�> @Re��'�Iw�8h�E�R�*�Z#MT�r���"�7<On�J�}"F��^)��5��M8���5+D��yR��[�H�9�//x^u�ċ���=яy2��{T�(^DF8@��U�x��B䉪3�`a;�-��j�́q`MS�U��=��''�����Ț�f��[%FC�8���!n6���H���r���7� ���N�6��E�+��F݈js�}��%����c�Q���=�#Y�Q���4xQ�҄o��=��!��ل�3��l��j�B��]�kW�L����*��� ��O�o/$�rrKү@���Z 8���O�|j��C���=��a���X��!>�6)�䆉(J=dC�I�MT�����"�nh�'�U��B����,w
C�O�Far!���l�O���	
5�Q�ƣ~nd�1���L��䭟� <��Ȅ4f���i�aM3~�ea�"O64�(P,
�jعj�7�^%r�"O舳V@N�n�h� �n�a��<(�"O�т�����,�TG�-U^�xR��	æ%���JdH�4�8�T�+U�hC�I72Ԥt�b��n5�@CK�G�.�F{��9O���ުڈ�SQ��G+���"O
;��ǿШ�ԧ׺w'塢=Ov��D«)�Qb�6mf���џ��Ih�O>��pUB��jZԜ�"�ܟi��C�'y�	�bBX��I���:��'N@�i���X��A����'S24�
�'�pZ�-��Pp`��H�$2�p�<y�n�k܌T��eV���z�Jn�DQK�O�̒o��v��\�b h�e�	�'��Q1E"��*���� B�U/��{A� �S��?IL%Kv`q+w�J����I�<y.U7����֫ƗR�}Pq/�I�<�%A�
~��Ǒ�F1CH�<�FFF?XQXq1��@�)!$q�#j�<9#-Z�X#�㌷W�LɃ��h�<qt#=n����H�0%%��� �e�<	�GڀD)"Ma�`X�]Z���n	a�<)��6�j�SEk�(���a�SV�<96��u<E�@1m���e�k�<y!�1_����i��@T -��aTa�<A���q,�Q�{��	1cS�<	 M���� b��=��=Wj�P�<���S'�,�S���/��PP�<1P�	g� `dD�3�"tP�U�<i�F
;=�
7C��9"SS�<�%.(�H�Z恆�L~�H�r�LN�<�`�<Jȸ���D�ug���vLK�<��ʚ�T�pK@���s�\�<����n�i ���%�~�S���TX�(� ���	�Y�v'��D��NV6\?!��9S�Ē��Ξ3��b`�יL<�z������{��)%h2��(
�3�!�Db�B�C�X�H�&J:�!�&J��Ӓ1FRᩑˆ�0H�}���\[5�ޙG��$���&qr�S��%D���p� N_6�k���&���i�%%D���d��<C��C��{���>D�Lp6�ܯ]$���n�A�F�c3'�-�S�[|JyQ%hŧo��`y�$�*����ȓ17���6�>;L!�r��_^^h�'�B듌�$8ړQ�Y�4����a�fh��S����'��PI��*�X"�Ɋ�>�����)��<�@��<�v���"�7�́�ևA\�<��!��c��8��e�@b@��d�<aP
T��2�� V=z�didJ�v�<�'73����h��?��C�"L�<��Ɩ�{�8�+�bwC�<ӐJ=�!��	G�,ĲQ��	:�|�hKN(a{S��o���M	�+��~l֨K�g�*g��Cqc.�D�<�O>���D׀(Sꝑ2���o����iРZv��ܤ;J����GY��� ��B�}�Xh�'��P9��8f咡g�08��'�z$!s�ğ-~|x�E<x�0!�':��E�HN��|:%o�?�0��˓�(O���R@��;�hKH>%���'趘'�Ċ��5�|��S��@��6��p<�S _?i���ޥ�4�ˠ)�O�'}ў�'u���'ŦQ������4D!��PgO� �����O,W�A5�`�A��'��'װ%yf��)s��LQg�\�����'`n���ø_�`�!2�S�Ѻ�'��'�d>��?��G��0���C��E3�ܡ��):D�T�҆;���Y0��(e���	q̢��zH>g�>��O�BY��1d��A��5Sw��J�')(�A-+�GѺ ��'WV��0�72� ��	��hA��>�O^��u���y vL�@䊓l���*a��y����	"�pܐ�.O�b���'EM��y��N�]ڈ0�B�a4KƯ�.����d?��4��S�Oߔ�y7.�$�X%)Z�W'0�	�'ۂ)V&U�f�x��H%�B���5Oԕ�+�5�V����=o�E"O�dhv�C=xp���,�hj4ٖ"O�EY�Xwj�����<DVf
��'u��<Qf����"Gm�9�!ʷ�C䉵#���g�X �Q���Ճ+�B�	@����Y5U��PE��-�VB�:_Ďh�E��,Q�H��U u�*B�	6}�hu ٽR�؝�����^B�I�O�ա6�W*S��Ċ��;+/�����"�D
49�:ȹ��س1������j~BMD(Q�*�#���2��-@�ǝ��y�"��e�>%�"�K'U\Ψ�5o��y�Պ,&�U��ɟ
SP�DR5'J��y�����8�MP�L;��A	��?	���s�J�ul?3ܺ�(�@�){Ў���'�\�a�Ѱ<eOP$�,	3�'@ar��]�$��t���y���gbF��y�	�oT>y��i�#\t���k)�yReݨOx)r�OPo�^-�V�R��y"d�7¬��肝7'N�j����y"��pMҹ	q-L�_�,0TB
�ybſHX�-2���Ss�Ah�+��y�$(=�+�'�&z��4�2H��yb��?:P+d�O�}�Ԕ�\7�y��	%c1���c�s��T�$�y��;!�̫� Js�0!�f/ת�y��1p�����*o����DC��yB� l<nX0�p�-����y2��C�Ma��_hg(�pm�y�"J�0��<Q�f
gt�12nE��y���t*�L� �P�1.����<�y���&���\�#���C�&4�yr�4�$�R�)����� Γ�y�/��&��M���
��5эS��y�M�=j�:�"6�ң0٘@�ޏ�yr�96@~mX�	�0}jZ`����yR��.N��]3W�U�&�(�bi	�y����U���g�q���s�ά�y�Z�p��9�I�z����@#��y�@';���g�@9C�t���!�y�%�A�\�(����6���@B�>�yRN�p;��	�Rh��UkT��yb@��Dh�@ᘞY6���*
�yr�V1�d� F���������y↑$��FK^�r*��I�n�K�<Y�`�;K�� Xg7�``��JB]�<ٕ�=I��#�A24��]��.�a�<A�=�"بP#�D��0+
V�<A�_o"ĔH�D^�	F����"�F�<i�O	�
������u�@x����w�<Q���4SE;$��9�R�#Ӣ�r�<���ݻf���i���& '�(p!(�I�<� F�J���;���AӇ\J�5ʒ"O����F�/X�ȸ���Uq�8Ԉ"O@(lF�30���l��\��̚�"O D��U!��Ϻ\Z�9{�C���y"BW'%�*=8�ʬF֦���m1�?a���?����?����?	���?���?����Q��H��Y&KlT���T'�?����?����?���?1��?���?	$m� 2h�l@2J�(�����?i���?����?����?	��?����?��A�%o��A�U�b}��p�	=�?���?I��?���?9���?���?�gE
1�����Ԃ#v�,�#���?���?��?q���?��?!��?Y�T�D2���.؋X�V�iB�Y�?���?!��?)��?����?��?�d&�\��
慖�xqo���?���?)��?i��?����?��?	to�.jz$��,�"�$���C5�?Y���?����?���?A���?���?)�)V�QX|�Q$ha�iӊ,� ����?����?����?����?1���?��)-j40r�ʓ�L{ĬK�<�6�y���?��?���?����?����?)��+���$�U�B#��zp�Ͷ�
(x���?���?1��?Q���?����?)��P[���Ŷ�ҕ�a�`�T�y���?!��?!��?Q���?I���?)��p�L�Ȁ�B��� �&�;�\�x��?a��?���?���?3�i���'��u�4ـj��L��������%�<)����󙟘�޴JN��K�T�5ƌ�G&L?� �$L~~e�2��4�4���iӀ89E߈M7t�ya��j� �p�Ӧ��ɦ	�*m�Y~Bo�o�$!rKM�)�t��-bS�[(.59u�ο"�1O��<���	�*�K0 V�QB���Nܨa���m� 
b��r��y�
�+�r�pa㙍�Nģv#�0>Ψ�w�F�IIyJ~��bK��M��'�,�������A
�I>�!���m�������b`��`^B���D�'n�1!FT�	��}�7��mJ�ʝ'c�|�I��Ms��̓3�,�b1��S�P�!\�R�2�BG�<���M�'��Ɇ|z��Q$�1*vPb��s�^�}c��І̀�"��|z�ȍ��u7J�O�sE��v�Iɕ�%MF�����<!/O���s���&�W�n�6��⏆�FT����p���ܴi]���'%<7�/��?�Q��J�u� ���a�W��q�c�O �$~�l��6G�7�"?i��ϪQ�����'�CB�A���"�Bi�d$X�$�كGc�3
�SA��xR�E��a�:r n���!�3��	a�&]�0-�yCưƦxbq!E:&� S��?(��"O�<��$yp�'�̘Z��|:�"J�@���g e�Y0�N�sYm�Q$� 6`�D��A�O�t����	iz��Ӈ�/J���IE�Q	2�Ц��7P%L��4�ա�c��S��5f]8�b�LN�E!b=�'+9 ��vG �{ۦ�G�4or��@D���z$*E 6����`	��M+���?��"����!'X6?
F�C�aĞmM�a���d�OXб���O�e���$�O8�	)�ԧ��+0�0qF���#
��M�!�H��?�������ʓ���J�R��$�'X|t(����;�*�l�%��8X�4�)�'�?�D�O�-|]x"BT6���c�w(���'J��'gr1���'�T>�	{?!��Q>�舑� p�h�C�m�1O A��K��|�������F	�z���I����D&���M��-Z��J(O���O:��|B�'C�����c[��ٱ�D�2��f�t��� Qb~��'�R�'OB�'b����d��tw00�A�) E(k@m[b�'���'���|��'���ۙ.�H�♈)�������U���V�����O��d�OB���O����O�ق`�\5 �,�
r�� ԰;�b�O��d�O�D/�D�O��W�%y��i���C6&z	����bA�Zj}r�'���'�B�'��GX>E��N�����l�T�el߆�n '�p�I�SQ��%UBrO����S;P��߉����Ѳib�'��ɑ5��u�N|�����$`�M)�皭XD�ŠR�I�l�4�o�uyb�'ObBͥ��0��iZ|Q���:
�,ZpkJ84k�zӼ�zM�uq��iʨ�'�?�'ch�ɽSUP ��ݔR�F�!&3�7��O��ʿ����|B���&��D��j%zhP�O�*�܌ bny�|�R�M�Ϧ������?)�I<ͧ��9�t��{ꐘ�$�R�y
p�i7���c_�p����d�3�ҟ��SC�W��`G�*2f	S7��MK��?��[�V�QՕx�O���'�^�CG,�-Ҁ(�Uh�$ir�V��>����?�Q	�a��?����?)��BlE�����X�D@�(��?)���' |��e9�4���D�O�˓lE��@�H#U�l����	u�Aᖰi�҉ֳ�'���'�"�'��G�R�I2�LϣxUB	��v�μ;�
|Ӛ�d�O:���Ot��O\������0������"�����Y�$��AR2�0?����?���?Y/���WOҦ�ۖB`߀5"�a`k��@�d��f��d�O����O��$�<��$p��'~�Xc�������8�m!0�8�S���������џ4��2n��޴�?q��b����ՁRM3~�U���LԢ��i���'��_�x�ɹv�$�S��T�Iq.|����\;���u�@��l1�-� �IΟ��I(F��$�޴�?���?���X�l�@�.}Pȗȇ0<&$Q��iRP���	����S�������t�? ��{p���Mu�@`��	*隂�i��'A��Kob�"���O$�����	�O���U��
<��Ze�شd�$t %�W}��'"���7�'�ɧ�4�~z�h�6H��#h�0_����r�ϦyYr. �MK��?�����'�?��?Y��y�J\��cZ,�j��BJO�&�fa'��'X".ۗ��d��D�O�u�q�6>��h���O1X,���b�D���O����!m�2Yl�� ����4�I��]#=����NR>�	�D#F�V� b����1�I��	���Y�ժ-��	[�Z �8X{�4�?��:���' r�'~��~��'ׄ�{��@u�eA"~��O��5<O����O����O��d�|"���q��Db⨏�EfX��/��Z�(ذ�iM��'{B�'��'���O�uQǋ��Eܦ���Iԙ\�9�G�>��D�<i��2�?9���?�P`�{��i5,��1�W�D���ZB"tFn��Ž�pT����T��՟t��ZyB�������4+�:�+P�3��ݫ�	��x�n��D�����Iϟx�	�vM�ߴ�?��K�d�!w �z���p0�L`��}�!�i�R�'�S��ɉ;���Ο���\�@�"цB��Q���͟tj�eo�؟x�����$�!;ش�?���?��'���si��b��+G�6J�-r��it�S�t��	L��Ο�����4�* !��7F<lAҴ'�$	��dnş��ɖ �갋�4�?���?y�'���u��j�n�q�,�a��+պ\P^���I��FX�	A�i>Y���쓠�Ą��!:À+c��zq�i�vM���u�����ON�d���I�Op���OT�`&-I�uI̉��;!#��h��C�����D���	���0�e>$?��Ӛ2pA	� �IX��ғ�5���4�?���?�J�]���'�R�'���u��=e�8����$3�2��E�I��M������Nc�?���˟��I=e4���6��/����NZ2pJ��4�?��˰_���'R�'���~�'�L��y	�T��F٩�c}��V"�yrZ�������D�Io2���NT�f0��ɀ	�!K,��˃��M��?a���?q�]?��'���,����DΒ�j� 8�%�N7t�'���'��'�'���'��H�}�6M9(C�S�L�%+�)(��o��`��џ$�	��'F�%Ԏ��T` 
��Y-Ԏ+tKĬ�`� ��l���O����O���O&X���KȦu�I����ǔ4.�����F�j�/�M���?	����d�OHq�D0�v�䷟lH���=.�XhL��
��TIp���D�O���O�4as�Z������L���?�0�
=��x�&X[�Ɛr6&��M������O(���7�����<��e��!R��pcq��hd�yj�	n��i�����oȖ7M�O,�D�O��	柶�\�@��йT�R�eL�}1O��3���'��� �Ek�'^�i>����=Ad��oȐ��D
1
��ܨYN����
Μ�M;��?����Z�'�?Q��?�e�בYF�8ڸdL^\(Ճ�!ZЛ^@  "�'�rZ��h�S��3�lV�JPx,�(�S
(�{�ڕ�M����?�+~�y{�iR�'
r�'�Zw/d�A���N���dտG�����4�?y+OV	��;O�S����֟�Q.ڹ�pr�\+]/��C��5�M#��Bi`����xb�'�R�|Zc�lը�,L�n\p��Ͽ.Ѐ�'+�%� �'��	̟$�Iq�S4I�T�0�iƪu�^�h'��~��=s������?q��䓨?y�[�&�)���'03Dh�"/ޯ}������?9+O��D�O�Ĭ<��I��n���6\�@撺]�t�P�L@�w��I��h��f�	��l����.'���P'^<R��T���J�]��쉬O���O��D�<�0X�^��O14��s�� }��J�E�N:h{��p���$7�d�O��D§Xh�$'}R��� F���fF� ��P.��M+���?I+O�u����@�SΟ(�ӥ �]+����d~4y�����i�I<����?�D���<!L>�OF��@ ��kfЛ�>⼴;ܴ���.�\lھ����O"��A~���2$Jd�Ѐz&B��Mk��?i�n��?I>�~�!�Nt�A�w��� X���UĦU��F��M����?A�����x��'pjXj�}���En�wE`��q�sӖc11O̓O>I���=L�%Q�� :X�0���բv�Hm�4�?	���?y�����'��'3���rxh$vlK�tޢ|���V�6s�6�|��l����$�O����	J�ze�'p����--f5ڌm�ȟ��uɟ���?Q����[���-�(����sQ�bG�K}���hW�X���	���cy�ew�M�IV�:��lb@)_#�*�(9�d�O���3�D�O����1�j\�u�N�]��)�gF�G
� 0 ��O�ʓ�?���?�+O��G ��|�b�[_h8*NPP˖p���{}2�'���|"�'��e�9&��IaG��S��B^�R'\k����?��?�-OT,�Bk�-����a�-c ��D+T�5���ڴ�?�J>!��?I6j��<�N�\Ss%�?p �����&%� `v�d�����O�Z|@��%��d�'@�t$�)tp�T��o��^���ڐ�HP�fOV��O~ Ȓ=O��O�ӻ$�x3U(:�#�"H36��<I�-��xB�&�~����J��,s�F�V\��d�Ulv�F`�����O
�0���O֒O����ŀ�v���J�}R>uC��i�����r��D�O����(\&���	-P�"%eA/�qa`�N�^x�+�4m���̓��S�O������;� ۔�S�dp���UIY��(�G�7v��3��H$[����0l��hML��9]4(���T�&��(��N/v�����;/,�ӀmMz�q�U�'Wh�w(��rr�pc��	sJu��jÙ%�b=�g�2g�)�X:�9�tb˝k��4S��9�<�Ҩ�C3��ٕ�B(% Q)Q
U->���MYq��I����xm���.$������M�~�t���	Ңc�1��o\ Y�� ��6��}1K�PO�}��N�N�6������|����ɢh��U�I埘�'m��ٮ#�������<�h�Ij�=�@Q��.���� �J���O�H�@CխOst�����aCf�5iJ��C��el4I����T&�7m�p P3��$
9�bs�|#bR�O�F�JB&ZgO@���"Oy�T�F���k��B!a�Ȼ�"O*��BV8t��H�V�$�Dh�7O�xlP�L��a��4�?�����II$ˈ��sQ2v��i�em[�/l����O���O�I��F�m�BM�2��/A��`&JUn��'5�\�"C��|Hт�7�(O~�´!.����DJ��p���~a�ϽY��W#��(yL�
�ɑC�'�9 ��h�2ʄ��>@9P�$�+;��Ȅ"OL���������у�&d��'fO�9����fW0��B�2Q�b�	�9O8d��æ�����4�O.R(A1�'!��'Z\]�FM#��AӇ�@d� �y���S��x0�<Y��4	5�N#%��'ǘϿې�7��2�H:X xv�	���3P�]�t�ʄ�ʪVМt�s�����6�U�"6������mK t	T�m��$�O��S��w�I3�-"�. )��we�U=�B�	�Q$ޡ�!&շ~=�x�BK�0an#<���)B�J��a��
ՏA�Q	��j	�?��^��iQ���?����?a�[�N�O��D�*5�L������4���d�4�	�[1!Y��@�Q�Ѝ(eџў\��fI.W���ÁN5L�1�X>�?邃�98�p��W�8)�^�3ړ"Z�: $�jm�q�#�ח �,���"��E�	���=�#̓������
�^�\ͩ0�_Q�<�P�:o��L�~��ѧ�_5uJ��"|"���6 ��F�ؓD�H�	�(c� rR	�I��'�2�'irQ���'3r;�,�� �[`D�I��I#?�2�hV�'�,��a)C-KD^���i<<O�	�"/C6[+�x����9���vK�"D�+J8\���РG�^��@(�&���`Lj�{bM_��?YS�i�e�P�:�8��1FJ�Z�@�(�'�E�ԭ��b���4$^>a���2�'��t�glǲ#6PAį�#�(�J�'9�7� �˼s�\o�ßd�Ih�t���ҹ2�m�71p����O�;�`�'��'v��%#�"-3K*?��T>�XFC
r�1�b"�)Tϔ��!�N�(Y&�J�ȡ�b@ֵf�\@�W��A /\!\��]�Wk��r	fAbd�M�'E�L���P��>=:#F[��,�(�<[j`H�k2D��Bg���b��؈h"���͌E���N<1թyV��i� �2 B����<!B�ѐ*	�v�'�X>���K�ß�����Cҡ�2t�`,��F�%���Ж�9r�Ҵo�8	l�Y��Ɩ^��Ij1�ӯ@��(�|��(X.�80m».��U�E

�W5��"�̗:���lS�_�rX@VCǨle�d3��;��Ͽ���A�B�Q�%x"�����:�x�1�Y�&
�<��e��?Q�)2@b� Tm�5/�f`@���<����>d"Õpd��cH�0�l��l�H�'Mh"=q���?����hq"8��a��2�c�c_;�?��P|ʀy����?���?���	����O��ċ�^�J��4�C�=���3�P&(�`d�k��O~��E�	��e�ݟ����'K��'�zUYE �
��T�a(�+g��GI[g|��1�C�2�6G@���t��xx�q�o�h~R�Y����
�$&$�(��@>�~�Ն�?��,�f|Y�aޤ���О<���ȓOْ�2� P�V�|���#ݟ��Ec�i>�%��2���!�M�T,��f���D�|&�A����?Y���?A�Z�=����?��OS�(��4P��%Î-hu�W)|Ș���	:�p>���˦�j�|[D��ń(4����&�%�����I�@����֦�#��X,�pŅ�,eNH1�'D����Ō�GN��a��@�eF�+�.&D�TX�Y�{rT�qa��;��}{�Ff�hAش��T�p���iqb�'��S>@���"��X��9MW�F�NԪ�������ɟdPfiI�Z˺i���@�X�6��|zf�p�v%�ƛ�l���YB�'yD�Ye��X���:��Vn�'#(�1(0�̋ ��u2W�8�:Dy�,��?�����BL�bh�^�.����J��!�!.A8@��B�5Z��0���@�a|i&��Yb��X-T.Xj� ��2����)�r1m���	l�ԅШ.���'�R����L��ϑ9��m��$� #�4���'�1O�3$z@��vҸ�Z��c�<�K�j��O?�� ��� #�7s���RɈ%)��4K�-J�2��dm�)�� �0ő#�����PN�z�X�,:D�X!�j�1C왚���D�0��À5����'^׀p���Bjڍ�+W�l�l8R���?a�����r�����?��?)����4�,U[�SB^�[�`_:<`�&��d8BٹuB<�@�
1W���ɧv���	�=0�����>n�J�Z�!�$~��-�E�tY��h�?=ʷ+G�(a�x▜���,Nv�2Yp��V��ԊٟThG+S˟p��ޟ��<����$����,�C�Dظ��A	��S'!�P9�Ҩ�I�2�z�A���%1�HGzB�Oh�R�t�5�'�MkUJ�
9@v�P���3gG���G��?q���?�����9��?y�O qxӮB�d�T��%��4�PaX��0ѮU9g�C"b2�;��X�%��#?��+� t��r�L16�T�c䍖�2�(Q'E��`��O�v��y�b,Ӕ�yҫ��������� Z�o� U�T��S�S|\��P'#D�p��
�R��w�S�^�B<q�+D�)�,��!�9(�G�^����`�s�T�ݴ��}�LԻi��'�ӸH@�ճÍ̞}	x�҄հO��|������I؟Læ��,њA��O�Ke8��1�ٴx��ɘ�<��5YP�T�@H�����(@Q����B������/w,L��4fq���a��%�>4���!l�R̂B�Q�3�P�á����0�P��	��H��A��JJ.ԠaphԿ��lA�"O�,�ǁj�L,����c��"��'�NO2��T�Ď/9��16�P��N�=O@}��!�٦9�	ǟ��O�^���'-��'�h ��N�cf.� ��>K��RCnΫFo�9&`Re�X�W*�O��Y��P&DǟL�vx�����$ɛ�C-�l�DjC2-��sBL�%YW��]w�AC�b�����*��j�y�J1Ѕ���;m��@���L���WC�)��$�g���h��e�g̿#��C�!��dʡ�ı_ݬ�`w�N�#<7�i>�I,�@P�� ��+�)��C�
-�I��Ps'e��eX����	�H#^w�w��h�c ��1x�(P�O���q� ���oR)x�A�41�X���>��t�-ʓT3@��ƛ\��Yul�e|.iI�%X#b)��eO�'r����OJ� 7{����#��drPap�*P�Z��֯R1�䃂~���'� �S-K8fT R�A`/<Ar
�'�B�Y�Z�ț7S�a�FjT�i��#=�'��)5�b�i��q�Eߍ>f��P��`����'aB�'u��ّb���'�		VmR�'o�a`PN�+��u��l)l�\с�f�h�'�����!�>�ơ	ק��4S�H�6�\��/�M���	9�ޕ�F��;gnt�P2�O`�<��&�P7+ɬl(�u �)�Q�<1iˡw�
����?A��z��Q�<�P�iw�'���w�h���D�O�ʧGڰ�&�A�w�NQ1U�L�~)���HR��?)��?i�֔�?��y*�be�d��?V�^���.4i�4�	�w����Eڬj�>���jO;��MSi�'�<�"��h��p�O޽IkrQf����h��"O�dEĝ�X\1���$!�<��2�'��O Ha@![�=疥���J���%��>O�I�����y�	����O7@�s��'��'/�]c��L����� �|���.ul1:!� �*�8C�.�;VV�bR�ۣ4M1�'5[)�xٕ��Vl�D�zb����ď�MF��(BOɍ~.������?�x����g�L����������f�ǝE�h{�KĚ�?���|���'��w���|��	;�T��'����6q:�B�O-7��H���Ln�����'�zt�'��=���ɑς45[�j1�'��a����x��'�"�'��b�E�i�i�Q�+7FM)�jF��V-مk������&�O| ����:| 	T �6^�>���O�i���'�D%#Fd�� 
(1��oP)��P�'l�p����=�2��=}��R��?	�f�S�V�<!��Fۀ�9�SwH��&ɻ�Sc�	 �q�شj�!�{"!V�/z�����?	��?A�-ι�?�����$B46�>���T�t3��у�0_p�b�K�aM`��@$9X���#L�fDy��˛SM�����5e��QlS�_��1���&!�h�@�,��K��TBR���Fzܓ*���I��:ʊ.!M|d���l�Ỡ� D���U^B��� �$�^��#+D�\���U R/.0����dDy�Q*h���ڴ��M��3��i���'M�Sg[�)p�+��>��a��+S�,V�;@J[���	��3�H����A��\�װջ%_���I��lܬX��E52�+T�m��ԃ��&N6���ޅ�p!�G�]����^뇫J3x����%k���[�BI-N�L➰h�$�O��}� �Lu�]�%��H��R4{���T"O�����q#��J��
�'�.O�@���lHa�����n���g9Oڑ���W֦}��ٟx�OX"�P��'V�'���#%�i�V)�#k�)J��
D�V'di�g���פ(�L�v�<U���Ͽ䱵�|�#s�Â4���q�@Y��{�ڷ!~aЎ� >�(�!%7��i"Bc�����#fE�9t����ܭ]_�����;`V<��Dy�)��$IT΀�%:H�u@��q�ޝ�E&D��� Ki���p��(j�ޡ���6�	�\��4�T�dU��`ӣ�V���e��2u����O�u!�m�'\�,���O,�$�O��;�?�;Ix��mP��D�z� ��MPJ��B͏.��҄,7cm�	��#��|�RI=�8�,�4�ȡ<2,)�d�G�����+ߌ{H`:C�X�h,���DH�b�C�� ���������$��$MpMHT�Ԕ[ɚ��c&�3<�D¢z�ҥf�N�'�X�	ԟ<�'�����Q,$��Kڥ'�I��O��=��R.O�$�A���.������9\66m�y���M������'���D5�$l����܋�!�*�t�sJ��Q����	���Iß�I�x>����|⁌�T�n+b��('����2'��#R[X(���6[F ,�L�.|e�N��A����K�wv̤��q>�)�I��M[��D�4����dl����Z����'9���t�?�OS�E�g��7�8qC�)hN&�2�'Yhq5 S0�^D���¼t�T'��L�����b�֝�;�?�����D6���0�'Zx�Ъ��)B�AW��O��D�OJ�����a�RDY��E?l�L��|�3"A&T��Q�%+�]�*�r5̂M�'��h�0�8D�>��&�FM��lsK�P�[$h�$M�J�)�=7�@�3jZ����=!u-����`����M��tC�H��ZR$��
�(m!��/��jacZ_��5�̔	va|�A6�
�/�������0��3!*��Ě�5>�l���	A��ϝ�x���'0b�^X�)�S�*B$8-●��bi���:�"#�߹J���T>Q�|�Ʉ8l�E[��ð7L�4[�)��T�tL�1�Q�U���Q"���I�v���¦��->�ϿTW�����b @�q#$#�@rxeX�-ɧ����O	�Bic�_�4���{v*N��yB�������K�*T`�V���O��Gz�O!��T;[h(B��ŝ,��5�������'V��r�A�i��';b�'�����$u�$e�R�/u���T#�,<*&Az���0
8�$P�q�u{�¾?=h��$�2t	�T���j���]�
�����T�>a�D���Ų�,����d�W=Z~�Y���_��Ɉg�0e����Y��]R���h��I�n�8�ɒ�M�Բ��,O��d�<a�k\?Ag̔�WA7O�d����l<!�'�-�Bđ�5?��i��G�%L��3�I(��l��~y���C�:�ݿ2p`$�� ]���a!�I?nh�������ٟ�piO�� �I�|Z�(D�
��l �+	�|C�96�$`�(��#�4��K���<Y���#s���Ъm��P���Z�`t�Ы��L��	�%n�?M"�hH9� DDxR���?QF�i;4���hO�E��{1C�p5I�'�:����w�pz�,�l%���'���G�\�	� ��?[�X�@�';06!�D۲,�\dl����Io�t��xz��a ^�[��x5茌��q��'��'�@t���٣N�)�R:U8�T>��$�&3�)xc���}�,5x$�?�d= eD��6`t�Q�G�9I���yd�ߣyM��ق���`fT��
�B�8�o�J�㞀�7o�O�G�� ��L�ޡ�EY�4�Ah���y��Ú3�hl�n�OEB ������0>��x��3	����&��
CF aٕ�ű�y"�݌SJ�6��O����|rիڠ�?���?1���M�N4s!!�7or�n�K��X��N('f���� 
�`�*�^b>��ë:� �K�O�2�d�P��;Q1<��P�^�l��Q0-ƿ�Z($D��� 
�IѴ�X��Ͽ������'BM��<[P2",�|�� �Ovb�"~�	���M�5��/:%�E���V:~C�I�]�>lС뎦s�tM�f�T�E�"<qB�i>��ɱ1A`t)U��S����O���Iٟ����:\��p�I�����X�[wW�w��9�����%��l� X��|8+/�x�d:��M�qcNu�cK�����鉸F�L()�\:Z=.F�	<4�bg�H��;6�اc��E��e�?�oZ#ZSn�3E2?!4k����Xŀ�,>�q�G�Ak?1&��럠��I3���G�Ýu�QBqBW�<%NC��������=$�l�����T� ���4�J�O����æ5����2Mcp�� ��������L�I��z,�	㟬ϧ7��h��Ϻ�l��6�ӻ>��ƣ_?"_�4b��[x���l����O.Р��  ��}���U내��֚v�N�A1)I�O;RYd
� ,0�7��5[Ρ���J�-�"�'+J�23&�ga:�wm�o-���!�|B�'+b��?� "<��n�3s9&j��	-m��D��"O�A*�(�XqR��&�X�1�^J�5OLnʟܗ'������~�����iD�v�3�F�U�J�0e�C�5Q~�J���O>���O�B0��2(�,2��^�g�$lQ���f�td�� �
@��DDd���0�(O�ҁ➸0���1F�
T3�9��u��@�H�n�.@`�,�!m�<EK�.W@���,�I�!U�PӦY؎��l'�6��%IM�C�*镨���y��'��}��W:p�D��∘jL
I�E���0>���x�Ku}jE!�MW�[}�R��	�y�GI3N�T7��O*��|:!ƈ,�?���?W�Et@dçN�U_��z$�TyB���C�I>K��6#R#as���wW?��|��>�|��k�#�*Tj>`��a��k�ր�dY�t���%
��u׆�/�>Q�O?���Q�Y���˪w���*�6{��e�Oc�"~���d:���O��g-���&�0`6�C�ɪ1i�-xҥ�	�ti���##�#<���i>��ɕ�d���B#ъA ��X"e�v��I��*٢p�5��֟����(Yw��w�����(�hl0�C]0�<��h�.�������3k��`�×����I�t�ȸ��՟^�=��%?���C���C�����֪y>��ӊ�?�o�(*�}�=?!%bܢ��X�TK�� �$p4ɞ~?	TĂşīߴ8��'��'!� [�H�:c�*6@�����$s��C䉛){�c�h�u^�y�U3S�Eb��������<��ع<R�V��Fƀ[�	�t��O�>[��'���' F���'k�;��Ȼ@fęI�`H��Q�r1�RR+©c��/Q ��Ө�/��y���
 �DR�> 6$����	|�z��Ɔ"w&�+c�D6��A����>�n��a!\c�L3���I��M�B��
Ew6����P�-���\�<���=�`|Ac���z��0k[n�\E{���>>t(�F	�)t��nW��y�x�*�O�3u�q���'��Bd6��CC�5J%��Q���$��(�B����l�	Ɵ��`-B�z�@�ĭzVa��战����0	>�IC�$�.W��a�`�	\�Q���-�+?D�B��Ѷn�|�fպ#KB�5�B�	Taӓu��sa������j�Dܓ~Knx�I�M�P�	K�^r�{Q�K{����팁;T���O���X?�n�  j��3~z0�	Ca|�/�K/�P����T�t�AG��$�d�|%m���(��Y��%��b�'8R)�Tl����7S�` ��-I��� � �o4���!�B`�Wh�~ڊ���~5:-�kr_D�Z��L��,�'Gޙ�:qX�C�<�A��n��~G����yO ��f�~���HԺ��H y�i��)�&l�N؀��@쟼�<E��~̂��Dα�x z� �����ȓ���� �(F��2�#����Gx"%��|��N;B(�%�<[�(�x!n��[�J����?ag*R�ɖ!����?���?�1^?�:?�
�/a��5Y���C��� �R�uTm;�I^
v[��&�?�����s�Gՠ P�����J%QE� ��*P��PÁ�=^�*ҟP�����(.�=�!!�>٧��u��|����|6>ps�M(�?q7�˷�?)��?�gy��'��ɔM�d<#TN��"WX��ƍ��C��֟��)O�T ����&o�`,;���HO���Or�t�$E{�ir]�����(�\yƔJ �3�'�b�'Ab+� ;x��'f���8Ҳ��b��j�H���}M�A	�Ǉ�9Yj�`ř{ܐ�{D╏������8u�k�ɑR��� )ԐC�T8�0�I� e��ذ���x&b�"�6�2��-ʓ�ބ��՟����2�88�0
ær����
?D��a���-Y��	x`d��Qz�$�G>D��P���9�cS��4O��pr�@��4��Ajh@D_�����ĠD�M���S�#�uٖe�FJąJ���'7��'����gM	g�&rvc_�N�J�!խI�Jd̨�w��4�� �6;+�R5]�(OT-�e;�l�3�`�+ N,(���mS��:��N]I%�V,�*b_�;5/�(O���1�'�7m���m��{�4#��3"�YP���]x��(�O!��s�8��>�Qci��>����g=�Ob&��jf��)�X���,)�X[ы{�\3r$L��M����?�,�̵b��OD���Oh�p�
��Fer���M=�x�W�ě'Lb��iX;��9���@,�M�O�1�R���r����f�$���W�m%�� �/��B��H�LF&���؎��'�H��T�DF �p`�����Ň_ �
�B�F�<�|��?i�Ԗ<f�P(��@�WeC�<	���>Q�� 
�Z�@"M�u>��˃DN�'�n#=ͧ�?	�C�C���r���s�,�[�c��?!��2��`�'M=�?����?��x��.�O:�DПe��9�� ,�D��T�u�A�U�V9/��@��m͍:��Y+4ҟ#=YaHҞ5���҄�U�m�ڂj�=��=P - 4ȂU#�`4���'�HOX�%C�6}��(rEKS B�B�	a�O���f�'V�{2��&vJ �	ԥ:e�ڦA޳�y
� �
��oEjM�@��h�@�)T%W_���t�|���!9^7-Q�`�����!1�<�!	ȡfQ �d�Ol�D�Ox9�Ae�O2��j>!��� 0T���/��1X�m�:+��M[ �D�>>�h#��ư<�D�]�|]����V,'����ʚ�c��(����v�fPs��
	�|�;�kC�hO2���'��6m�e9���!�/c� �)�,1!򤛇[�^���Y-7ެt���V #!�d*;�N���
&��I�\�N���&�1������OB�'MJp�tL�n�����.�?�^@0t����?����?q���zS
$�
4h�di4h����S�nz����p�|5s D��<���֥TZe��	�K�<u
&�N5DV�K%!J�eH�M�^e�HB��	����
����̟4����<�O�����*��r�6Q1��@茡1��'��O?�I $�\}��ʙKe��R��b�
��d�i�	�L�lZ0�P+Ap����R=y��I
M���4�?����iD8�z�D�Oh���R�AIf��4��@��ʹq�:]`��RFDyI����f�F8�\M*�Ss���M)�n^9|��1����v*��Y���)���*�|�Y�%!Zr�X���w�.1H���<�̍�S��-JvS�
҃<��|�Z}���'�*O
��5'G�u[̊���MFfi��"OR3�#�Q�LJ���SL���ቪ�HO��oʟ��r,˭*
e�	��.'8a��������$f� �qBџ�������+�u��'��͞�̤sW!Ы6ƀc��,�~R�ӣ9�	�3��?����ĝ�fhH�T��%Vm�i�4�1��$�8Z
�1�KG�>�(��ɯK��d�!<N.����@����I$@�,��'�M)O���O$���O��[���"�	Xo f��Bl��Y�!�$�?=H6�p��(PT4i�0L�$�Dz��>a,O�|y�����a���Ѐ��j.�*����a�՟������	g��m��ɟ�ϧ*�,%얈�M��n�Y��'����ݘ\���D�,F�=�4jqӆA�����p�T|c֩պ8.>��B�'��x���?��ߑ/�8p�eB�_�@X�f�?����$�O���'a��)���$ p��Яɀx��p�ȓrP�Ǩ;E��r�Ѓ��Eϓs��Jyb�48�6-�O��$�|�⧝�S�Fl��i� ��;d.��S�$l`��?	��K�����֘���� 6�q �X �.%��]dQ�H9�@7�')|(`fN�d��qHL	:�)EyBo��?r��&,�P q�B�b%2��WP�zB�c����Ac�:|a�98"�R P���$n� (�r! w14�v��e���g���	8�lp���H�	r�B��r�'��,�j�pL�_�� QT�ϪO�J���� C�²V�|�O1��yB�%u�քP�h�c�i�j�)L$�����u��E!b 2�J�R'�=O�<�~��F��JÚn`�+�G����Pjq��ݟ���4I��6�'�?����@��[`��Z���Ѷ�J�zT���O��d8�S�'E��m!�mZ�h�KX9��̢U�'�&���MyӜ�O<�*�c���Bu�6�
'��^��B24��	��� �^��#��qc�L�g�%D�䣳��, X`9�`f�j!v�>D�@YSBYs z��@��$��x�� ;D�|�G��2�"i�R��Fg�\�66D���D�3�����׷e�\�
0D�����&����TI�)�<Hӣe,D��as�J�M�T`kgJ�l��Mb�F,D��`�V�OE�|p��,��}�S`+D�̰Q�Q4"9*�N�w"�ō>D� �똸&rA�.A�^)��=D�XR�	�*��K��6�P(x�=D���e߽lO��볬�";�D��f�:D���b�56_�%��-��<�&ث �8D�t�!);�j�§�Z�WB! 1.;D��@�
z�
�	�sjId�7D�H倠Q&r$Q��F�0FZ]Y%*D�p��R��`ˀ?�Da�6A(D�ԫ�)&I��$�Q��,��
��!D���o� ��qf��A�P���)D����ث�l�b/^��8D�+D��y��̀4�RGE�W���Y��5D��7��.\��I��3F�܁��2D�� ��in�=`�̄��
�6:jn	jb"O6!YC�^s��ITjߌkQ�M��"O`�S�_��p��fʤ+R����"Oz�B��F�p):��H2ZjJ-B "O��k���.n�*5ᗨW�/[�(r�"O�}����X����`Z�;�"O��Y�� /�%h��9PD��d"O����f�xI�Eܙ��f"O���ڨ.��1�2d���a"O��{cCD�9X}{e#�Tz����>���V�i(�]�7�iy�7-�|}J~Rf�4�Hj�m?�`9�HJh�<!Ra�� �H���K�K�Ib�����T�{�,ݲ�'�8c>Y(�LH����2a�d̩�όUBD����*T�!��!=�!�K�E��%hu�B�8��(g�i�|(ⱠB�D-nT�w
W[e�z���޾l����*α=�����Ꙣ��x���xG��Bn�'
�'ˠP��D�P�pe�X�&�%b�%�!a<a�
83�lI2E�vpm�&kL@�	�vm��EǺDLP@cn�	�����&yӵ&a>-a�E	�D1ĭx�ş�A�,"��14���
T�0�jT���ƶ�,�k�/�P���V��nm�0O�1�Uiⓥ<m��~�&��f��;)��x�)��6�h��=�0O��i2!֦��*��M�׎M?�"@I�$0�3j@� �8��IS��)�W�$f�Fjh�b�8h�"M0�_\6MN������n�tjd�n��BA��K�*��~�,Ù'>�'#���(CGP�=/��s�"ч	� �
ҪE�r�����!R�����Y؀�%��?`���?�Mָ'����.�a�������[%�l��#Ee�#U��HX�h��
ʁ9B�@#Q>�8��.�;(��ɇ~��f�� �(O�p�&�+{�(����<>���b��>q��J��QsE�+���.�o�䚘I�Z��L�.��q�H|��O�A�'ӨL+(h�c�0:��Y���i#�e�a%�L�B��T၎��
,/�(]@�!J�e���0W�ن\
������%T��Z��'�<���!V=7��4)�.!1��x��Ӟ/��}�wo&�A��[�WhzH��` ѐ�6��u���w��ñ��w��T�3ˊ�2��z�TP8� �VI�kN�� ��I8�p-9@DS��&��� =b�hܛ$a�	��:ei��6��L�E�0:D�к3A2?�H��[m̬؃��).��!�f��\U�GD��nZ;s��!�=Q7�S�g��0��<����#08$z"A�9��!cċ��ky�1 �g�ݪ�؞���Y�(�>�HIq������[� ʹ5a{�U����kէK�7���-�\�Zd����B�V2aN�s7-�:W��1�+TH�����!BU�u�\���cClI�ih�L�f'��,|��dY�)�M�b/��B�|��\<3�ْ�oXu�� ĺ_ud���$Ԛ�d�5��mi���E79��cu�� �.-�	+B�#%�^�'�)F�eD^�9R�.Pn�����O랟���Ŏ(ag�@$Gc�����+I��Y��B16�Ep0N]>qK�x�]�>됌�cA�3�ƭ�v�\�v�4�ٸy�49eb̪��?�sB���G�L�50���A�6�9#�Z<I�}�x�Y6/p���u�\8��it
�8����i$)��@�m�;�(�)�h�az2O��5�� �o6K �J���2I8Z�@Z�sl���H<�HO��ICK�\-J!�%˯y6J�	W\���%�I')o��K�s}v��Ў,�	63�v��Ԇu���ܦ��<��F'nb
)P"K0����jM��I��E\E�B��eV?\Z��=�I]�(8���v�
��6Ĉ\�d��Ѝ��3�h���,�@�Fz�>��W�p���0��<6B`���Klp��y�"�	5%�d�,��$ �8�i��$�~���O��ˍ����L�$8�"�NT)6��Td�y���Q��&~C0�p�ϲsZ�g���T|���#;�\��U�����>����;0f������P:���U}��ݍ*@�c+M�?���!��HO��[��֣G��ճ�.տ"���V��{��7�x�BF/8���(z��]��/H��A�UPDY��I���ɚ��FBδ+�� 
!k��䈌	���b �\�"����\�A��F{B�V?��9� �+x� ��R�]�4h�&.�O�M���4h]�@sцȽ5� c$�$/pM��-T���	�@���ݼEV^�8���1�ҥj�E�V����$�*f-" ����@?6��d�"{~T�V�m^��`��$[@}��&�F�ؾ_��F�-�^ �����&lQ�/�Vՙ0��!�0$Fz�)�+6n|i� շ+�M���0�M�������&���3o�'Ę�g��O~|bN<9ǈ�`��>�j��&���+'�, /�d�r���MQ���>e�Ճ��,�.���M��?�S�\� ^u8$�E�.� !P��>TX��E��X���'`,)(0��P�&�q��ΆN�*x΂�BJ�dr�l��� ��L>aVY���o8J,�v@ĕl7 �J0�:�O �l���?���V�]����#1*=�������h֫ہ��'x>�q<�<���3O�l�[� ��r�-�K]�zy['6ړ�~r�A �p����^=�R7��P��,�.w(��'a��{L"�p�R�P�q�B̈O�S�G�j,
��V��(s�:q�i�*��I!tP�0a�CN#b�O���A	ER�Lh­Ĥ;��,a�KI�V��R �ۤ�p?q"�!k��� �N�"��C@�gr,�B�i�EzZw�8��@K!I��N�~lPJN�?ݎ��S7a}���L�,ɘ��߀]̪��i[$i�Ȑ��O*Mbb�����b���
�o�D���|��Q�R����"�x�F�*C;�^�@�E3�n��zc#x�����/Z!nz�7-��qb�(�A�tc����3�	�K�Ќ;'d*O`�ge�8x
n�<!#k]:=������M*5jd�Cߦ�Iè�{?4�²�R�Lx�GNf���I 2��h:�`����QCnUpF& ����s���a9|O�X�3�K���9�׮��~��E��xC�~�;o�b�e���%��(ۆ�FU�ϓe�(ق���G!F ��fc](~Y�p� WG0��޴��D`�$�[kB��Ǝs�rdrtë+,�Ҍ�v��@%�xy�R���9G`�&���m��(�wƊ&�P�-��v��Z�	�v�FEۗm������@�e��jZ�m���O",�d��$�h#=�eL�c��2Ղ��I�L��CG��ƕ8�C��H����5,@�K��1���B	������I3^@����,���R�HMFHc`a�|zr�p#
�} �K��<�}/B�Q}���� =��a/޵J� m1
ӓH�ై�J� ��O�Jt����
�?�*Eڀ�Z��($�T��y"OE5���&$T��TLQ�B�V�i拈�\�Bl�b�D'}|�p�R.��T=��q�V��&>�I�1&�6o&qOa��S
��bU.��������s��L$#��H �L�u�F�)�Ig8�e�_)t5-D�X�(��p��f�t��JG3!Qa{�kJ�d&��W.M�l�B|A��G>��H�iB<eҕ�
�,a���Ǔ�G�J��Ǌ����'%��jM�q����FE%D�ɗÆ6�{RJ��<i0mjWi]�1+x�)t�DG�ԋ��[�\`�����$$��T1SՉ��K�����ǀǽ�0����M�bP�b���z}J�`B�I�Z̨a��'XFĢ"��1u��6&\��R�_%>�Ay���Bdb�'����hٝ�M�u��)Wb���S�I'
$��;Ԡ�qy�y=�pQY�%RF�hT֘|Y�\QpP[�#�2NZ��o�> �� ��W�(*�nZ����[��P8�����61͐$Q�B�$ �Ɲ�Ʌ�^��`�Y2�c��]r�)���El�GT1:��؜ZCf�h���X�̀Ն́?9��3G���hځY��c!ˡ���SL��;'�R���	)/��q�?i��Næ�;3�� �0�WjU,q(��	0�;�dE�"�
0΋�sc��	�C0?%V�������YV�0�˘�i��$�2hY���M��'F�M��.���5���ȴ�V�2��	�A��MѮ�'��D9&�<	����Qm�y ��X�'�����M�g�'�.TK$��,�I���Z���@E�R�r�0�F�'>u&��=�����G�D�ypS�H��80�aKcӺ����)�q,A+%��� �2���	1*��N"��#��N���$!W�1��u51|Xvu�d�ЙR��يt�`��j�	٠c���b�韜+a��q��Jc�?��5OhӃ�!|?H�:$G}ʰ��֓��*�@�v:`�4ZF��E �/-H��J�l ��ΧK����eO
u	x(���Թ6�� ���*���R����?L�i'��K4�D|��	R$�2kƤm��Y%�J�B�"Ml3fM�I
�q�,�(��X�?���р)�l�d�Փ�$�س�Q :�f��_X��n�Nd^���Gn�����]����F��. ��s��O��'��S8M�츱_RR���Ӆ��^� �����*#�)	Ón���� �߅gu�6�K�RҪ���:%�2����+���Ґ����'t����4En��[�C�p�=�d=��t�'�D���V*\&�څb � Hk�O�M��2 �@�֎���>�HA�OPU������W�T��T�^4c%U�HJ�M�􃚻z �݉b���*!Hˆ��O�'����㞩�0�2!�O��p������8e C�~�o4w���M3!�|҂M,a4�Y��H"4r�1�wbr���Bާy'�ˁ:��!g	I"ftzJ�bA7�M;R��O, K��^ �^-&��Y�t�&�۱Z�||�@��)��a��E��.	�JW^I�3S4Nb���q�X���uR��l��ic���R�֕9T�,5��F%&�)�O
@���F	(����c�&o:\ى��֊hn-c�؂��dۍU���X��E'|���E�{�����I��bG}�#O�}th R��3E��+r�i������"M���q���~Fz����Mb=07F�G+`�B�t�i� .�#3�4�{H<%>��E�~z'�|VЁKuZ�I�|"&���7��P�c��a{��� ��Sf�3P��P���{<�^����J���!�����H����#��Z�ˋ<z�	B�nM�&�\�h
�orH�#" �ua�p��"VtS�+��Y��;U�����A%�P�	��ܨ���Ǝn��i.\�c�I�0f0v<j��Y�[ 0�hP"�9{��Z7 a8ըT63v��֮��8���)�8
�*���C�- O�C�^-jnB����B����Y��(ЩA�=Fx�f�1#Y���Lέ]2�
7FL�_�1�MI O���L<%>u˴"����p�'�%q�I�1hq��1:Y�EFJ27����Ӽ�B�S /��PBӇG	O�V��NG`}����y�JO=6:H#�!�7�?�ë4�	�/XcT��&/���3r�`��A)k�er��9 ��	�|MJP�ꎔ���1��l�1fS��~rOZ�<)�)��r"�D�X�t�)����!�ē�04r9�%�4|�	�^.�!�$J�z�d�h񲰻"��?�XU�"Oz�
@G��qM��r�Ǟ :��P�"OdX�b�I ,yhgi� 9�p�"OP�;�/�C��A�g��@Hw"O �E�C�.� �s��ѫ����b"O�<�5��68��`[�6в�I�"OL ��F���+ �I*V�|�"O�"'�X�}2�j�-�"�҄�w"O�[q�y���я@�aܨyi7"O� �	��4�C�W<'��]�e"O����5/9�	q�'=�&��"O$�U �� ��L�E��S�"O��I$����Psq%�Ѧ��T"O�������Ij�mx�c�}܎��A"O|�@�	�x
}���`� ��"O�+�5{�B��J"=f�{�"O�Xu;Y��R�+ �H/���R"O��E�Eҝ2��Z�-.��"O\E౬��c�hʆi1|(�#"O(� c/�>EWx��hU7p֬��"OF,��%'`�[��\���D"O j4@��x��'	�~�h��"O�d�ϘG�Щ�R�6J$Q"OX����V��x�B�o��욶"OR�YUBP6.ۦ�R�*zPA"OvtZA��2+x�pp��9'Kl<2�*O 8�1AV�sA�uCB'� t��b�'�:Y(�̉��j��6�V�� �z�'���k�dØx�4��$��@��'vp�`�/ryX��Şr45��'7�|kW�N�)�v2g���`��'��phQ-0fkjEyq�0�1��'�f� �a�7&������Z����	�'��#�d.FS6P'嗛[���	�'�F1�\�le(���	�T�̜i�'g2�21LH�{��4u�ϦZ����'�f$���ؠ�ty�tM�5a*HT�'���(�.O��$� ��
$�eH
�''(�2���c�t��3��}�jDB�'�ŃC��9"DH��h]{S��Q
�'?^�z��10�+�=l���
�'\RL���P!0��8S%H'h��MB�'��H	�@�6@.:q��D��\x`e��'(ؔa�AʄR;,U��6U^8��'�(��g�wl`p��˶I�Vh�'����`�na�p�X&FB�5��'�� �����-sc���H:�
�'0�d�b�G�M�1p�bH	tW�U�
�'�ʘaGð3':���GU�t�t`�'4��i6h�5|��ㅌV�zs���'����D%F*)#b��s�H�	�'��0z�I�~�J4�1���vl ��� F!�ϩT���'ѦBA���"O��QD����r	�>&$Q��.P�ԩO�gb�ir1�6Z�p�ȓ;���[��l�r�q�f�$��ȓ�c���,\����`�꼇ȓ@�	�Ov9��b��yJ$H�ȓ<���c4ͅ55�L2'��(!�9�ȓL?8�R���8Uk��3,�x���0� }jb�\�/Ĺ`L�/$M����-�q(lcD�mi�m�%f?���ȓwT�$J�JF���S�ZG3$���BuIa��e�HA�d�&J��1��,l900i\ z���HA��C'��ȓn�����_�<O@)�dgK��
 �ȓ����+U�]Vp���"X�ݲ��ȓ[�����^$H1�� ��*��>Y�WK
D�0�G�b!���DJ��89
���͜l�Q��2aPQ�v��1��ȓB��%С�	D��1����n����?���I����&(ʝ�SJ5l	����1�Z$AۡM�@i�#��ڙ�?���~�d��a��L��4��ɂ�O�<	��/��hAե��;�|1F�I�<a�m�0a�~ �a�8[�|ի��GG�<�TG�6��R0MD3)�L���F�<��O,n�i3Zib��ȅM��~+!򤌈��y�mÓ�x��^!X�!�X��@�RoE@�,4iC+�'�!�D·-i�hB�V���IrC
�r7!�ḓP��1�w�O��<m�fE�s+!��>aN ���0BĤ��R���=���G�4��:L��H!��I� T�S,��y�EؒQ�j�q�#ʹvv�ys"�C?�y҈�W��僢��?�hHQ�G"�yr�O��J��Ш:$$�$���y�)Z�	o��1�.�3� )�t/Ǯ�y� T$ؙ��*�4Sܚ@�Nܛ�y"�խA��蓄C�:$���?�yB�P� $X��ʨ��_�� �6O$]�t�nct��DJ?�ؑe"O@1�K�@���(�i�?h�ĭ �"OL�1�
6-��X�T��2����+�S��y�c3P�ʕr�OҀoOVY	�K��y�k�0���˲�O?faiauÚ �hO���� H�zq�2�K6h^�9��C�azB����0������	�^]����Nul� �x�I��}9T�f��%XH��!����<	��ITPU���<1�lIE���:ЮC䉢z�����D�;8�[ l)[�B��4I
❲q�+��$mĕP4�B�Ɇi��H��ձS�eL�l��U�Т<E���X�;�~ p���h����4�K�y�_�#����d;B1����)�yb�Q6B\��fOD�Y�,���b³�0?9*O�u��CN7{���eI\<��,P"Ob�)cc^<~��X��1Z��M����OX��&DYoNe���2p(�7 ���p�'8��	�b���&x�4!@�|`B�ɢy�����s�ٹ���q�����/�/���qr͉	JŖT��Z Ms��ȓU����je���-M&�t��C�J�x�A�z"T�cI�*�.��ȓ_�؝�_$'��)sh�$o[Z؆�(�$�1DW��h=��D!ˤ���S�? �����?���2jD�,�8���8O����ٕo�PB��[��
�G�,�!�Ą�H���ؔm��6\!D%�
Z�!��	�H�$9
�M�ss�0�tj��/�!�$��
�p���#��=�����;,!�d��l�AㅒZ��-����'!�#1B�1k�]������e�!��
{NX0��hٲx��D�w�*+!�;�&�Q@"\#4�\L0��:p�!��qi��K�"ϛ|�
�3b�r�!��4kz�\R��ܤ=+�`��c�(+�!�DI�Ĭݑu
@���� =�!�$Wm���Ã�+ �,cSFX�p�r�	4�5�S��?��E�u���'�M��pE�1��c�<����KF�`�2�V0l�E��)�v~��'��Ձ0A��&��u*��kk\i��O�ʓw;���`�#���5F����,��q(D�͌2�p�H�OӲ#���Ez"�e��m)9w���6H˽A��[��y"-T�|ؙ��R�:�
��Ύ�y�4J/�����\u�.ӭ�y�@�[y�Lc�ϛ ^�X�B��y��S	���w-��tC�C�c� �yD���,x�hn^���M	+�y�O�j�~H��F�jE��#ŗ�y���K�
�����i����:�y��» ��]�"\�_V� &����'Zazr�EUo\�	��-	Tj�2B�7��x�C՘��;PG�R�B�j�K\�aꓑp?q@NF=A�|�e�ɺ$.t8S�+U~�<��L�	�*Y3C%�7.����"�N�<94b)����RHƗĸ���@c�<a�6h&�
�E�[�mb"*Zv�<��,�/�t�YDN����Bͅt�<yq�K�3���z�N~;p��B)l�<�Sf@�4��t{�Ĕ1kض$�)Jo}�'��|2-�U�ȁc,U�#tڽ[�e�۰=�{�j�4=���`CȎ4 �QG靖��' �z�*�_�\����Q�2�`A��L��~��)���>��$[.�pe!��W�I����J�<�&M�������
�L�ީ `I�J���=y�r覹Cw ̿J�$�Q�a�<���D0xN #`���S��;�#�`?q���ӹ]��
"l	�Tʽ����$�ܢ?u�S�T�\$�R������3���s�B�5REKI�Y3�ā�(�[���'��If]�����<	j�N�F/�B�	�AL��"��r�4�-��zU���B�ɱ����O����]�1�'o�%;�4,�c"O��ۓȁR���7D�%n� ���"Oh;��wZ��D���%�Y��y���!;������4_ �j�eM�y2i^�h�.t���82�J|9B�� �y���\n�e'Ȥ%'��a��8�y�"ߠg��5Y �̅!D>�j���'Ǡ�=%>��RF�%FR�����D�tL�4m?D�1c��R�5�S�Ϛog���9D��q�f?1v�EM��z�sӄ7D��S����-�dD��S�\+�@!�$/�O*��u���F�������>13�"O �L�x�湲׋�5��Be"O�kŎ�T��ݸ1� �� &"O�z��	�2����*ͩ}��Qh�"Ot� 3�֦F>���1i�C�ār�"O� �ui2iB�a�Rd�E'	�`��ّ""O�����A;r��Hׅ��> 	��d#\O�\+5�U%w���n�;1�	��"OR:6�NPLkv̝::��)�"O�e���qY>�����O���B��'<��"w/P�G_��*��ǂ�2iCү)D����G�|3���S����'�D*�S�'w>��w�\�g�����\�R��̈́�>L�]��N����0��@^(�ń�|�z�� ��� б4�ڎP�M�ȓVD�لč�DkP�Y ͦM��7@��Ҥ\9L�LiP ��9�.X�ȓ��bC�Ve]M3]K�`��i$v(��I/�'�^�ɶ�ȓVA�<R��	�h�V�9��/�� ��;�d��U�V
�Y���+����H�p�bo�M/�(x���5'�ȓd86Q���,��`3$�?NP��ȓ$Q�t��$eT�+QȌ:n�E��_��e#��`a�h�I��#>�1�/�.�`G���=+q��
�la� ¬Z�J�@��'����ȓa�����J��\ؐ=:�AH����O0r ;B*� ����4n���ȓMĜi���f��T�`�ʰI������^���LӉa���1C'>��̅�a0�+�eM�S�b���&(6���w��ę�G��_i~U�
W��ȓw���It㟫>������J�Fԇ�P��Y�!^�c��C�?n�ćȓ4'<`B7����¨
�E�"Q��X��tY ���:u�D+d�ǒfR]��UN$�CID�;W��)��]��D���7'@��4
T$��� �����=�;/�@���O P�<�$B:#\鰔%��I��)���N�<!���.%���I&R)a�]Q�<�-	~n�[�$�Hz�Qc%�O�<��^�m\A	���Y@�b(AM�<IU&|g�d0A�PE�b��`L�<q ���O�XamT>JF�sS��M�<	V-��q<�u ��2�04��K�<	�!͛��`�	�U��86*�E�<ѷ�ɢ!��lS�DC�Gmf���N�C�<i�M��H����Ȇ#�	��I
}�<qu��('/�XHT�k �N�v�<���K�|��$��mI~О|	 �t�<�5n�/�8���܂ ��4�Bo�<Y�̋c���&̤t�p YF�Xk�<��bӒ,[re��+V䀒�@�<�hS�}�|���V�%|\x��	}�<�@`ǘi��H�B�`�neh!c�u�<ц�\�fT�ˑ E#V#����C�p�<	T�ލ]��Pp�a\/��B�<a �P)=��[��D�1d\�3d+B{�<iw$��T���oF�:��S6Ow�< �.;<����*����"OZ(��WW�z�����%<B�+#"O>�:�
�+3Fi��!�}\S�"O�����6 hژ34�F�f���"OZ���D�*1xlS�S�FF��"O\(󲎝�I�\����xE����"OJf���L�%JL֦.��"OX�3Q�F)pj9P䚂/8m��"O� �,�oI:��!�e	����Cu"O)����u�򝰒g^�I ���"O�ʧ��I���w��"���ȓ;Ǻ�*�U�0�Ѐa`�A2T�����{f>��dGB�F�y�◔�4�ȓP��u8�ƕ97(Q�v@j�
���M���hag���$E3%$�$v~���X���0UdL�dzT�ڱdN��^̈́ȓ�.8`'c9&�� �3"�9d�m�ȓ_.@���F�;/t���cj��H0�ȓ�x�K��ˊ%�ى��
�A8%��g-l��Є�,8U!aJY�^��ȓY�a�hIO�d�l��>	L}c�'��P�a ��U~5�Тٔ7y�1�
�'xL��ei�4���Y���6䮡s
�'��9酣��F49P�&(�dђ�'D�h��/gt�x�w��+#��k	�'�t`:EM�)[�����J=	�T(z�'����#"�%u�*�2�k�: �q�'ad��u^r%2��]�n��y��'��r��_^)�Ds�nߋSu��Q�'?�ݢ��l�.9hE 	�z}����'�����,{��5�U��ts��Z�<c��2C\Rq��"_�%�PE�IJ�<i�O�mÐu#t`  ���[B�<��E����,��hډT=xICD�C�<��!��^u�����u��I��#k�<��M�[�n��F*A�
�)��c�<I��R�6	�!�oOH9��\^�<Iw���^��` �A�x�pɸ��u�<��ꁍ ���� �l��e�4�Xl�<A&)�7V���J���^��@��Om�<��A	V+bdk��E&Rb�pc�aDC�<i3I�5�d-s��+�	����}�<Y�H��a�p����>6�R��|�<�SjC8;U��ӄ�r�H	����s�<Yc�I�D�v�a���^���'��s�<�.�Bq�}Rf��:h,\kG�v�<QeDۂu�pp��<VFUSď�s�<�d��5�(��:d�,�ᶪ�e�<q��Ѡz���&BY2nt��dXm�<i�C�j�BA�P�D��0	1+�k�<y`eȝ	��iybK�6>��0�"\R�<�Bd]=g`jH��$�x˰�if��F�<yw(�"b�����$�\�y�B�~�<9�A�A��bK/:K�����}�<�rIӧ2�Xaw�ǢD��I���P�<!0��Y���@�"�}�	B��I�<飉S �ĩ�	L6.=X#ĀN�<(�&+t�L��d�+=���Cv�<тL�Z�ƨ���w�� ��v�<�&���X�|A{�GB��2��ab�s�<�g�@��~8�f-�+L�6���R{�<YQ)X����A�F%sk�P4B�t�<b��z�ʑ��	�y�EC^�\B䉠MG����ſ2�hb��2*F2B�I�,��h�L�(�d)���A.B�)�H#�>T}P}A���	c4B䉕6ڨ�6o�#p~@�����BqbB�I����� �_@�Ga�W�B�I~�E�B'i�R��cU�@�B䉳t˖�� �6yPzr4��D�C����[1�$S�68��1u��B�It�؉	�ŋ^}""��.	�B�)� ���.�o��y��L�M�R"O����.�0��e��; �y�T"OtzD�Sqx��G�4I��x�"O����p�iPmN�:��� "O�\�f�?/�������Liq"O*dapS��1�Cg�*a�r �c"ON�x�nM!yY�0!L!Tܘ�"O��z��A�v�<�V��
�P��"O��ȃAȉ3�Y�cG�k�!:"O�p��K;8�a�9ڞ\��"Oh R3&�*I��b�5���r%"O��*хϧx�(�@"��Z�R1��"ObɛQ��&;��p@�Y�ӜI�"O��y���)x�	� �k&�0	�"O����ұ|B�<㲡9�UT"OԨ��#4>Et�˷%ݱa��i�<���� �+�>q�lP&��]�<�s�	4h\ۂ�Ih�! ���Z�<����#8M�8f�S}6�����X�<��.R}�nM��C�:&��`�}�<�DL`@0�ɔ�{���@�A�<IO �r�� )ӄ{�2����U�<Qh�i�|0B��0J����VF�<��I�u�YYT���0�,��-�C�<I#��t
��k�aUEjZh+�͐d�<�V�Ћe��ۤ����千b�<�X�$�^)P��2"5r�Sd�^�<�Gf� $�T� 吵C�,{��r�<�r�O�!��F# �|l^+c�n�<i��5SUм���
܌q͍j�<q�����̃q�H�b�:�z�m�<C*I4
���i�W&4�^�O~�<i�@Y�<jI"���7$U,�0�d�D�<Y�����P�2EN�c=(��'�C�<��5~R䱪�$ˇ]<���API�<�&c_� ����g�Ӽ�%cIG�<��>D׎Q1̌7::�y���A�<q��E�T�օ�� �e:��:c��A�<���ƴ�8I��D؍k1�( ��@A�<���=w��p��Bɇf_��Sh~�<���11l��B�N>���V"Zq�<��!?V��Ū�vUZ��%�l�<��ʁ !ܨx����j$J�0'%La�<!s��ub)�V�_*B� 3B��x�<�e�J�!$�(�+R�Q�&8�R�x�<I`�D��4�H�n�:����MAs�<YV(Tj��KC��N���Ky�<�rcF�~qK�ۚ�P`Ȕ��v�<���8{�ґH'fٙ��I�5nCY�<iSI5E8����Ǫu0*tK��V�<1�N��Ǧ��B�ſ,��&��y�<	���\	Ȉ���8�N��A�L�<9�K3���GC܏f�H-(`F�<�F[z�>͐v(�>�l�s!PM�<q揇40�@�Ѡ`�=�$�6&E�<��ɕ,��y�JΛ}�N�d��C�<�Ш
�hѨ�#b�B#g�sb��Y�<�IL�V�����n�m�D��h�|�<���X�D9�0M3�L=#��c�<�R%��H�\�������P��a_\�<���Z0p/.�����H֩�@(�|�<!6��e��ыY�P��{ӭ�L�<92b�?��ѓ��Tf��+��S�<�V
:�D)t�ńJ��䉤��Q�<� N�b�+
�=KJ���L�[�4�P!"O�e��4P�d��"WV��2"O�Zsm
�M�j@�
�Z	�"O�x�e�)f���$8�0��"O>p���L-M�N���*�>��y+�"O�!��b��y�,�4d͹F��uے"O�`ۖ��G R�1WeZ�K���AE"OZ@�` ��|�zw$*K�^!a"O"�!����:�|҂�H�<���"O
9JCK�8����`@;M�1��"O2m���P�00!o=f4�`)"O� (���[��"�T8y2j(�"O8t�K�_�B�BI�q1*�p"O
ȃQD�$1Pn��!ǒ�DB5G"O��
����h���D��$Z�ʰYG"O���QS@-���ӈ|8v=�"O�9'(̦9f�eH�kI�j}0�sr"Of��iZ,
��l*c���4oH�q "O|pCsD>���F�-�Q"O���AJ�2>IH!�3�� N�����"O�X�g�ۻ/�6,ȡ��?r�"�
�"O��
��R$<�� d�;��] �"Ot�X�o@�������`���"O���(��"h�eA�KFlm�D"O&�1�k#Jԥ�!@�@z]�"O#A�T�P`� ^$l/�{"O�1�S�$���Z�M�'3D +�"O�!#�/� h�2��ʫC�V��V"OtQp%L.�Ш�V'�����r"O �H�DإW_4��ù9�H���"O@M�g����&����X�f8�9r"O�-���ъr��h�4�߂G�~%��"O��rP,@��=���ߩh�.4r�"OX�E�Ƭu���Q֮.�>!�"O��`����73$1��K.{hr<-�!򤀋�.E�`�ƍw��� ����!�D[�g�"ؙ�O�;�jdI�d�/Q!�D0_l��&�]+�����=�!�J�*�YJ�h��A�l��F��7�!��*X��<U���u��Ѫ!�ƍC\!�D��6�	���
G��]h @��Q]!�$��n�PYr��Z-�iY�!i>!�$K�N��$@A9
?,�����(`!�d�e(� �Ǐ�<I�Y�ņ?!�$	��j�a G�+���g<d!�d�+	��r�`Ï;#�A+�#�
!���c/ԄBs���-.��S�%K�!��+�ٹ�� &�(� 6/�!�I�~Y Äī"¥�w�t�!��/
̱�A�Q=(Q|�k�E�6o�!�T�T���C�̇|��rk�5k!�Ĉ��"�qq�� t��a��55^!�FL<S2���X
"U�s�ܠWI!�Đ�t�����X�A���P��T;M6!�ā�i�0M�)�o�X
��Y��!��ɪlȀ��j>>���S���]!���#sG��( �~�HBsn�jW����U�r)�SK-h���(��.�j��ȓ~TQcɲy�����OB�ȓ��p0��'���2��Э����������e	Jz����*Tв�ȓ	hx�)��1q��J����9�u�ȓG$��K�NZDF�M�� +[�p��ȓvXT����o>X����_$JI>H��S�? j��AI��&���q�"��\�p"O�E�/h�:u�G�9�|�
�"On bࠀ*��(���}����"OLY�$J
i�Q���\k�"O�ݫ����>��Eb"��lvp�[%"O�T���,h�Q�ul�9!b~0"�"O  ����sJ9�aI,��]#�"OԘ� �e[���#�I8A�ڴ��"OR*�e��X/^M��݋X�T@��"O�и��>0����Ȳq�R�"O��:jͶM����tF3?���z%"OH���*����	q�[�$$�1"O@�Q��	$)"j,;,"	T���"O����C�&(K����Jl��B7D��q�&v���# H*+V�ܙ �(D���ڼ�����n»^@D�X��%D���ǌ	A/f*���]�Z0��k0D�0ᵂ df��� �r�G�!D�$�!(\�V�OZ]���PFe5D�|B7j�,\�lպ#��>ٳu*3D�T� �jhtr�։s�&i
#O>D�lA�S5A	���t�rp<D�,��h��>\�����&���b�m'D���#����0X�p,d��d��#D���N��w�����	�0��u�"D�@X&�jas-��f���; �7	��C�	�$ ��j_0�~a�e@٪C�.B�ɱ~���b�	�[�^��׫�b)�C��$킍�Pf�)2�B�f�s��C�.D�t�����G�q�p�i��C��
���dM�a#��!~�B�I�
Z�Y��EMH܌Ѱi^(��B䉨����EФ������0��B�ɟ;�����ؽc�FE�B�	���h��%�ڸ��FL�T��B�I;|)�L�h�d��A�	��o��B��	��@g���k%����D� :}NB�	ff�q��)�A�6uzu��6Y�dC��E�<����?i	QY�)đR:C�	3V ۄ��B}��CVF,� C�I�m�ε+�͎`��E!�a��'�C�	,
ʨ@S��&6��LL�.\C䉨 +�tR2��+��UR�n̈KT�B�IS�d"��P����/0�B�	�,��隁ˊ�&zقf� <uh�B�ɥ�֥���*���A��Q�lB��RD� z4�C,]���RO�!��B�Fie�׍�%�p Ӂ&C��B�	|Z� sq�҃p�2c)�-@�B�I��L�'�O�54�B��8|�BC�I�S|2y��`�{Y<RDM^yC�Ii��-�%Ǔ	�@�؆�2�B剮nXX���AB�?����N��Zh!�%��9�䑎]�0L��!ST!�d�y��lirn��<�Z�*���o�!�Ę@�b4��ܟ��t�7���!�� 3��|���	;/�������!�O9G (�)��q��%Z�iяL#!��>KV$�vj��ʘ�h�1Z-!�I�4[R}�L*�ڑK���6Gx!�d�;n�fɃ��؝����x����ȓ�0�G�9L4d���׉VB͆ȓi��*D
�j��)��#$�%��\+f�IU�6�,�%�WS<p��S�? �Q P��@��[P �.{�4��"O�r��ժ|�Д{�!Т"U�l�!"O�c�E2J�qu�_?#C�#"O,�{�L/aB�#�II�/8� �"O�)P�
�� ��0�Œ�%��J"OVVː�V�>�ʓgͥ:�4��T"O��  �I-B�@L�@��3b�UH�"O��c0
R)|�t�&�ڪ3$j� "O��b���k?,���;L���"OX�Za�߱$*�T�K:| 8A"O� ů�{`�{��M�+Ds�"O8�G�J (�(�X�JN�Ԓ"O&���m��y���¢i�	ai��;"Ob�@� � p �"j
�\�*q�&"OtD���!h_�(�2k��~�X�2`"O@��ݝV5Z�@�j�>���"O��2h\�A�J���)%@��Ha"O>)�$�T�=�d�N&H���l"O�����00�D)��Y}ⅳ�"O�,B���
�,��煨Tvd+�"O�pÅ�J�`2��R��ֿK|@$�d"O������ Z�\W'�*ht�Y@"O�5	@Eڔ7�,d!�dZ#fPjH�"O �s�O�2����d>|?�9�c"O���MS���� eN:���"O `��#�R�P]�#�V"tL��r�"O�-*��8g���"mťX?D�"O������޴;D�߉
1:�"O|1Z mװ�va��%bE��qB"OD��B@&d",�Y�.yP��S"O� 2-޳��s�K�_M���"Op�Ԡ�#Y��iU+@�?7��c�"O���娔�"� �8R�#2�|cP"O^y� �̾,|�xض��1.%P�"O`T��V�k�6� G_�,�F"O�|�,�����{G��i�Fl�"O�����x#�AA�̎��h���"OlH�n�	�l �LT%���5"O@�����O��+�P
��"Ox����L�*-�\ T��\k�c�"O A�DU�k�<Q(���g8��"O8u[�JF�U�D��7>o�L:�"O`�ɴ�Fy
����(�=2k\��"OT�;��D�0�%�a�`@�z�"O�����q�:��G�LZ���"O,�u���%r֥I��Q�FV8��d"O�5S�+����� �)B�p���"O���&�%Y�1j���Q��#"O����`[���)3Цʍa��"OxBe�X�"�X�K_<[ӈ�8�"Oܕ�w�Vi������+�:-�"O,��mʪWlj�����D�n���"Ot�cB8d����Ţ_sJ}��"O�TZa�X�s�V����Hd���!"OvH��'AH�c�;� ѐ�"O~�i��hMFuȡ#�^�lP�"OF� �PCļ{Џ�7��@#�"O�$���o�J��@�F�^@��"O:�Aυ�\�:T�#��0&�0yi0"O��i�/A9zkx�p3E��B�Nqt"Or�KѦ�*P܆����U50"Obe�����
u�
P82l��"O�UAWcݜLՆ���2N+"O��nЫo��8聉5ܰd�6"O� <,�͚�t��)!)']V�b�"OVڇ�A�Zndъ0I�a���B"OVh��K�-��C��W�oF�ыv"Ozi���q! $h���:갱�"O4Å�ݫr9�ыp"׀���E"O޵�6kB9/�i��T�dY��"Ob12%٨?���f:z���"OT9{F�rp5�f�ƾ
Ը��"OX��U6�4��q(�jW�9�T"O��R��9ߌ=�!ɻJm���yR�I�Fcx�	�D���	���y�e�@�v�z�E�
S[�|����y2���0H��堙�`�ȕ3�g�yR�b}`B�i�;[98ŀ���y�L�h�z�s5*��d�T����3�y"ET�N&�@�ņ8�=9!D�5�yR��p�veJe�4pX�p�B
�y��.Jt�Dƽk&(��F��4�y�&�Z�"�{5��c h�0�C	��y��r�yf��U�xp�C�yrk_*�b9b��K����y�Xıb�q��UjW��$�y"
�u���hSm��:���!n��yR�A1X	T �H+G
ܽ���R��y2+U��
���.đ?��jҡ�y�("<�0�����[aȜ;�y2�������ߴm�X������y��T2XY��&��b�rТ `O��yr����}�f��]���!s�y(T2���� �^= Y�<9ҍY�y�GE1|�|QS*�NFxm8rb���yª�%N��]�B�Y�Y"5���#�yb+	�5�X��s�[9�6`�E���y2nݰ>dZH�t�H ֪"@�$�y�T�0ܶ1Z1Bϼj_0]R�R��yrd�+����!�^�Z ��D��y�H�n9�k�"[���b�	�y��D�0/�q��jǣ��0���̵�y2 �zn΄��+@�*Cc��yr�F�f��l+����y���c�+�y�풷:��$:áܿFХ��J;�y�K��2$X��C\#��qq�,���y���KмX`$D�'��r�'��y�ܕM��5[�m�V�����yb��;���жdT	@�x�L��y2䈟�D��R �*�PC	N�y�J�=a���g.	r8��!����yR��3;I9��\�ql���`�ڠ�yB�-*�yC���ذwaD��y")_�P�T�ە���*V0���y脎r��\:��<��eصlF�yR�U�JaE��ؔ9��@ⴭ��y�b?Ф���1c�Ũu���y"��s�,՚eŇ�V�0�S�$Y6�y�	��(�6�1�I�"��<��G�y�
M�4,2���N�-��L:�y��T�l~��P/��`QK�V%�ybD��}v�0�b�V0���g���y���6u6!�%ER�f�yb�_$?H��v���hZ%���ݲ�y���;v��B#c\<	���x���?�y"�ͱO�nT�\i���1��H.$v C��(TD�Ӥ��)bK���D!F�w��B�ɟG�r(2�"��`�����B�)� �hj&��=b�b!!GD�2��[�"O*�K�.�vN�1H��B��rXq"OT���JO��"�d�-n؁�"Oz�,�F�z��E�l]$���"O���G.Q�& ��E�f!h9z"OM��mM�RnL E � N��"O:Y���zX�E��N�
#�ư�"O@lٓ����U��L5/�v��R"OD�R&�	
/`�����MJU"OL�A��!d�xD`'���e�!��"O��W���Q)n) P�>6�6��"ON�A抍8D��4Ð�q�Ρ+T"O� ����IT 赢	n��(��"Ob(a��BQJЖ�@�U�p̑�"ORY!�ɫ`v��`Σ(�LP@�"Or8�U!TeM�=�
O	O���`�"On���NW��`�d�.\�x��"OEh��� ZJ��4 5! |��g"O�5A�FY���M���$�B"O��	`N�)Z��-���vDr�"O�A P\�X,rp�r̟% �.@xf"O�hj�)ٛ_ժ�!���=岠��"O�$ ���	|��q���T�1����"O�(0��:#������&�n�;"O6�!�j)�W�.�"�"OM �A
Y:�b��n�:�XU"OJ����X�<"��䕜2f�h��"O�
��ܠN�|��rd��s5;	�'���&ϙ�4�f���Ɉ*Ϯ��'���`�_�K9XU�7��́�'�^}r�F�*N��!�Ȍ�j��(�'���SΔ,�m!`����3�'���ұ�ĚcG^L�g��yGv)��'DBɈSS6a2�#P�
�n�>��	�'�(C�� $B*�|� �b�{	�'�&�1�a�lYd���*�=\JR���'���xr2�,�P��X0 _��8�'/
Q�u�Ԓ<��ݕb���'��t�ܖO;�I"'ԠNI,�Q	�'�}���@#�r,#�FX�JP-��'e ]�Ů�,�`az���o+���	�'>����ٰV�.1Q�E��tލ	�'�.ȋg��@!�sID�q���'���	̮g��c�L�}	D��' ��6ݤ"ZYP�_�a�h��
�'n֭X7m�")� h��ݨ]/����'f�SSH۬a�@#�`X�[�͠�'�Y��B!�8Б�f
;!�2E@�'�DI����u(�ٟ"�T��'1�x;�K\!?t1���I��4��'1���'@0�W��?��l��'��`7"�4N2x��U�=X9�'�8�B$���j��%`a�������IA��|�yTNQ!=хȓ>b(U�GhX�i[M�2Fߊ$Z����u�D)��
������1x��#��u(@ʑ� �D�ze�U�ڝ��G�2\2!*45�Z���<	d8,��u���vhE
|M��٠�Bq����N�"�jN��c�N�Z"��6�J���^��t���L*�"�/��e�A��JVj��wd���X�b�@��k�؄ȓ/�������G�2�z5�ly�ȓb��5�oS�W��@�a�x���S�? $q�m�8�āO��G Z�P"O���d�4tf�m�GN�<��9�"OƵBg�X3#⽓�G	S��� "Oy�V$[�<8�uz� �f���!"OJ�jU�W
H1���Teq"O�� �1v��r�Z�_���@G"O� !��ޒ9p���-���i7"O�!�g�.��kQ8f�BT"O�|Rb���H��ʁ�l�N<4"O�Px��+~�n0c��P>^��IH'"O������Z�x��(�&&�p48�"Ob9ϛd��P�w�^%u����"O�8�1��+V
�� '�	�~���"O�DP�D݌k8i�f%m��{F"O䜑� ��1`gÍ�`dꍩ�"O��BW
E=�ȜX��
l3H�[B"O��*T�%G7Ƽ�q�i�lq'"OH�����~|Mx��}�1��"Oֱ��/ϕu�\`FJ�g��18�"Of��D5wÔ���ܫv��4�"OHWk���,L`��V���!����{)�|J�-jt�8�7P��B�I6���W�B�i�J� u�B!�rB�	�)r&rg�@�<z�+`�<aPB�I�e'�Y�0M �o�)����'85jC�Ɇb2����M<:�2y��!�)�:C�ɠmI&�H�1H\�2G%^2�B�&H�d	0�ʜ&�R�i��"`�B�I'y�(,���($����&O�&X6C�	�4�N�����I�haE��&#�(C�	��x��$_�NG&eJ��O4C�	�o���4ES&$)x׎O4r) C��Q�ؤ�V.�p��{&�ϔ*��B�I�%���S�#�0���!D��B�I�Q���x��J�T�)��ܻS�B�I)@|⹲�
��C(��
U B�<B�	Y�RE�6A����d2B�WF��H��F,46��@�"��C�I�	�i�蓉Y��z��٧-L�C䉫#�*�se�"��#�c�!�C�(=��x��A��D�a>O�dB䉨/:�{��JWU(P2qT5<2B�(C�"�I炈%�TTpc�5�B�I�k�HHz6aO�H3v���&��q�B�	��lYӦ��	fx����m�TB�	�%�<Y�M�"[�^�9�h͎0lC�I�XMΈ��$�%<脸�b���2C�I�T�c�HÎ_ ^�q��á��B�I��@������`CT�I��B�ɢZ�6�( �Mm�4i�9��B�I$H^��8�G%I*,=�����$��B�	�|s��i�'L"�&�b���P�@B�	�L������P2	3AK�/.�rB䉷/:h�Cp*��J�� ���5O�rB�0^p�%�s��V(VIᷤ��nETB��yz��z���Z�H�!�z��C�	 m��Iq0��e�.���;ȢC�ɝ�L���;����΋�b�B�	�6�<�0B��07�@"�(L�B��Z����Ć�%ϼ4I��XƬB�ɲu١2�(3���2�Η�;��B�IR�|���J>�hP�
Խq�bB�ɊH����*ś����Q��f�8B�I�c&
�hA�O)��	 �-�DB�)� ��C6�V~8���F���9C@"OVT�T� ���D��&��QBU"O�@i���4�v|RN�	Bt�p�w"O�h�A�@�.�8�aAφ�[d��w"O�\�R�[8 t|�Ь�jo�U¥"O
(H"��HV�j�DFP��+�"O�݀c	Zw�ʪ?4X��b"O<����@�l�|;���G.��R"O,���l���^0Cs�Y.1�a "O��fAݫ*��5)T�{�Js"O�����Ǥ*��`��ߕR�`�Jb"O�8�r(&D�Ii�a���V"OԬz7���B6�
�Qo��{�"O����� d¦��(� wz(�C�"O|�q3g�n���]rٸW"O��J��@��х�z�n��"OJm�v��9�=��#q��-��"O�x#�.��h�vIʫI���Q�"OTŨq�1i�3Ȗ�*ɰԚ"O�ɐ�!�8�9z�d�F��5A"O�[�# %<Xyy4��ms�Q�"O����[��&�{c��`�0��"O~�����B�B�*���J�x|!�D\�q����ЬJ
x�$��'.!�D��`�Rg�@�V�C`B��!�D۫_��P�`�)&���%Z"aW!��\+�,�C';t�Y8 ��:LQ!�\�-9v{����}�����W�*C!�	61��P8�
$(ׄ�ǅ��)�!�O��=2�g���@�Ǣ��-�!�dе5F���*\6S2n��&Y!�DC=w2���+1ڌ2Ҋɣyb!�$�9[���TI�18K"xPW	A !�dJ�ux$yk���#�n�8rNľ�!��?Cn�Siϯ	TF�f�N�,�!�$5`��!C�6b8�a���Zn�!��J��H�c�KQ�-�5�Ik�!�䚐$��p���i4"��E!2�!�D�watЁ��r6�D)�B���!�d�.$��x2�E0d&"ȄbQ��!�D�x�t�م���+ V��&/�!�� �����5$ita"fd�!�D�B���"��+f��)4k��*2!�"\k��Cf��)X$l��A*}�!���3`r��f�e;2$� %ɳw�!�䜖L۪P�d�+��
��z\!��x��h �ɏ��p���Ԑd!�@<�,T��HGr�\Y!b�V�x�!�D̴q�����	�@V�,�2 0!��݈pQ�q`���;=䱰7E�G^!�D#;8�1��Y<�����	M!�$*~�xj�I��U��X��?~H!�D
�_{&���.�1m|`݊d�,}F!�ӄ)R򑐁��q^.�g�S�<!�D�~�0�����0⦄��2Y!�$��Z� ��j��2t��!�jBD!�$�--�(A�o]!M_t}�*U�!�d��t(㴮E�qi��X4��,�!�I�=�r��R"9POnc(u!�dG1H��7�W�'�xl0ŦC�E	�B�	�e+��p��ҳH�\,�ާ|۔B�I�*�L ꃻF]�}!'���ZB䉹<U�X�Ś�f�.͈���I�2B�	�1˦	�B��}��Q�	-*�6B�)� 6��'Q�.��@�0�è`=y�"O*85�O�4�&�r�u��YYR"O���Ĭ�%(,Vi ��U�;�-��"Od�Y D�x�CR������T"O�!x��UQ�}�C �Lօ��"Oġ��.�i�9r�P\�g"Op��3l���J$�pl�E?�=A�"O��B�*9�p���mQA��-j"O���OƵ17AtL����@v"O4��V�Z7q�\kw� -x�@��g"On���]'_��� �	Y�CA���"Ox�����ca�ű'IӀr,���"Od\���Ht4�{!�8i|���"O�xk�o[,l�&LH�E�"�����"O����Do��FFӳR���p"O�%� Efp� ��;�d�pR"O�c���!?��Lb�U�X���W"O���D��V�X�;���q"O �Kv�,v@�@B��z���"O��̐+>H��á*�:Z����"O$���N0l~�\P�ɘ(@�-!�"O2"�MT3P��r
��}%�9�"O��aF�P-�Q�ֈ��>n�Mz"OJ{Gt�"��`��
`B��"O�I�aF�A�\���ٻF"lp��"OBѲ7,� q���$D�@���g"O��%���X��A _���1�"O�5���O�a�ځ����P�æ"O �I֜q��7oV�!�Z��"Ot���E��8ޒ��1�ۉKǰ4��"O�����j�p$�"��G��3"O�X2t℔1�8�"畲Q��w"O��P��k���JTF�|gH�"O�	�')W�4�f�1�(����"O�	��?kb�(�⛢��� "OR)Y��9�*I1�gߢ#�Ā+�"O�p�s�P �t'�r�.iZ"O�%Wf3|s��QA�L�r�:|4"O8	���٣�\)���HG"O*��k T�����1{H�"O<�2���']�<(�
�u�|TC�"OHAa��X��(� ^�t!�dP�"O� ��	�-���;�>\��"OR�R%�9b| �{��j�Ej�"OL)jŉ�mWf�7L؆W�!R�"O��+GFϻz��Fh�'D���"O����/z����!<U���w"O�40�-�l��9G&��㔭st"O���D �L8ތc��M�*��=��"O��[����\����G��&i�|l��"O��)�H��/Q:8�ǋ/H����"O�<��'T&U�ʌ��!W�~]��"OF����`̴p"!7lҜcc"O:	r�JѶm � �4i��@B"OBT��aM�~O��eK�s�恙""O �BjF%*DX,�I�fQ(�r�"OP�t�ơ8��d`�ǒC��s�"O�Xp�i�F�blH��m&fI�e"O��z5銯�N�bA��1}"E9A"O�j�U?�:����5` 1�"O�Q���KH}����:G���&"OY�&)(�����Ғo/��*�"O����R�9d�s�'W@��B"O@i{��
i}@,(ڻ f-"O� �=HÊј}�*,rB�3���bE"O�X�A�	]Dv�%�6l��cA"OL�X$�C4E4�EKZ��&�8�"O��ᢎ�0Ud�0(�?'v$��"O�p��	\X!���<r�%��"OH�:���ek@��Hɗ>hl�"O�5��bE/d�~��
>
Df"O�hw���@-���M�i]xM�U"O�!���Wm8�@�M����R�"O\���,}�. �'��v�&�pC"O��c�?D��Ie$J�v|;U"O1���?|��`����Is"OHa�BG�F�I�l��H��A
�"Oʭ��^�F@H*��J1=�n��"O}"p.R�s��l{!ϕ�J�|��"O���j��H�gL�6�x%[�"O�(b���Z�v����),��q��"O���8��	0&T�V!v��"Oda�ԂI*�b�1�'=Ҭ�F"O���3�[�uNp �ţ��%�-��"O  p���v��# G�Zs"OpH�!�sF4rᡅ)sJ���'"OĘ�7@�0��)
@�E9�LZ�"O~0��
1��0�f���:-��R"Oj��ˁ�]�+���>j]��"OB틧�$)o�����}�&)�f"O��*Ĩ=<��)caP6#쐽
�"O���!k�Y%��"烪�����"O:�����A���1E�dX� â"O
ܛ�1B��ɸu��`��(U"O��ƣ,9|�Ja��W� a�e"O^�*Q�O��8p����y�>��g"O�L�cTM�%�r]�z!�Aڂ"O������&=�m�bƎ#P@��'"OY`S�\7w~�YR�"A�h��"O�5;"n�Q��i�4��&�F�Ɂ"O i;a�˾D��z!K[0d��t"OF`��������阗*�r�*�"Op���K2u��������-{v"O��{���'D@9����:5U"O*�ZC�4*H$��5o�FD~ԁ�"OƐX�'՟WU���'��:;$@�"O<U@�!��^�0���}�.�{$"O��K1)�~HX�s�5D�$��"O�
�Ù3�x���8wR(re"O��2d���� 2�@H�v���e"O.ݳ�g̠y���i�Y- ��I�"O�L���F��>%rb�E}&&��'"OV��lY*b�D���^:fz�ȃ4"O<Q�rl���A��F 0m"OV��Ro��$S�DD�_�T���g"O܅���/a�,�w�� [�s�"O�ȴb\ .�(�_�}��C�"O��QQ��0QHX� O�ܺ��"O ��6��?��ѻ�K�r0���"OBcK�DJ�hXf���$:�"O9���)�t�ٴ�E:Y����"O�&�^>p��ţ�	����� �b�<�p�
P�,���RD����+�j�<�� ,~$�5��=y��{��\M�<Dß�xdM��/Ģr�ڌ�T#�E�<��o��Y3��Q�D��:\���H�<y�"��x���`ۂ�-OV؇ȓ~=�+!E�+!b�����\��S�? P��.0lu����N/��C�"O��� FȈ3�t̑B
g ��2"O���t�Ƨ7�t�00
I=�Q"Od�Rm�'_��h�oܹ�N�K�"O� �D��0Qh���/7LBP��"O��y���R�ԓI	*y4>��"O�=���S�1*�:�BN�t����"OP%��M��{6:�"�l�d_>��"O�!pG�A�H��lA(;Y��Z�"O|�2 jߩ3�d,�Eѭo�e8�"ObU�G�I4x����f��{lZ�k�"O��ڗ�-z��[�b�?UX�A"O�\"E��;
PZ<0'���/F�U	"O����)�ԩ{���8��87"ORĂcE���T�*���6y:�"O��@��Ĩge<�@���/$ �a�f"O(QHoF��|�qD#.�� ��"O\���6%~`�yp��;�6��"OxW��"��Р���+3.vĉP"O<�*�@
,i�di��z�^�J"O���A4P���c�ħ��h��"O�bU�R8�f��)�3�$hS�"O ہ��5W�����K�r5�P"O&�� Ո9�P�c�U&&��T��"OeIG��+ʈ��V@)>�<��q"O6��
ב[�}��$I-#��2"O����%B�,z��`�y�F�qV"Oa:�R6zy�H��O�L��@"O �Sp�9R ��5O�m$"��V"O�<�rHH�jy�Y#%R�.*@@1"OX`�s���f4��p�DIR��Uʂ"O��)P<w���3B���P�"O���'TU��9��.7ޤr'"O�Ȳ읡a�xu��w~u�7"O�rp�2�ф�U�l�J�"OԪ��K�&�>IIu����C"O�`[��R��*�ȓyDX*F"O�uRƓ�f���#@�L�9ܠ�2"O�4�N�jdn[7c۞7U8 x7"O���e�ͯF��@4�5X`^���"O���bƒ�� i��C�Z����"O�Ms)
�h���TO)J�B8I`"OV�q�,-^$p��E����"O�5�'HK�
��q��.� S"O�A�S�\�rqXI��P�e��(��"O̥���K�0ɨ��0Ɲ�!��%!�"O�����M8��x*�EC�N��\b�"O�	�f� r�Dh����)l�@�"O�h�AK�6c��d� H� �ڥ"O.�V�S ����f!��Xk.8ZV"O%�k��Bz�IpG��5=Ľ�d"O$�UD�f�F`J���W��1ze"O�Q9��ѿԞ`e�Ү$I�M��"O\� بA��IUm�$=�L�"OY�dZ�@��4+�	ӳ#��� "O <{4�U+�t�S7)�v��!�"O��P�OG9U�P7�O&;t���&"O�Uj̚rZ6�Gnl�Hb"O���Rf���Vy-D�i��M�<��o]�5�^�ጻn���y d�I�<��"ĩ3�,E�G�6-�,X���YJ�<Y5�;U6X9����@���@n�<I��p�j��A��O�E
�Q�<����x��q{Ԭ�-��@2`�O�<�   �ǷIb&��`�*Ln��zU"Od����ױr�"@��j��m^��"O,����A5��t��H�[���b"Oؽ�NQ!tv�شHBC� �{"O,U*Q���� � 0���2!�L�<I��OA %�����D,]�<�(ǐa�I����gO`�P��Y�<Q���/(8���Ι7UVMP%�CR�<�$)h<t)��G'a�u���Q�<1��?\�b�k	'2�%�N�<	b!	?p��3Z �Nh���p�<��f�fo|��j��&��	2� �S�<a�Ύ?���V��$�(��*_N�<�r&Y�l����W����`b�<!��I!<��t	s��5Y��R�<�u�� t$V��K�F�Ĥ[�&P�<qFF�E[@�أ�_E�^T�ER�<Q��T9"~"�*�Đ.6�|�0-U�<I��\Qq �	?ll\��A�N�<!�0ɺuC��
�84����SH�<��,S^9dl����9zcdu��Yx�<y�N��[�I��X�R p�Z��t�<Y��\�3�^E��Y�G���Qb�D�<2D�
<yr���K�&)�
�\w�<1e@_�8���*��@�l�V�t�<)��_(�� Y�\_�(4jj�k�<q�G�%���"U.�Wb�A�!Wg�<�4�^�b�
|�eN��e�����n�<14��릐[1&��C�&�K-h�<a� �9W܌p��Ε"4�騆�\k�<�QjJ�FyC��	'�B�Q�j�<����>D���0M ��(����J�<���+�9�:Q|�ƅ\�<A��\ԵhU[29�J5`q�l�<��� �i�SJ\�$�`a��]�<)��Э,	|��܌V:@�Y��Y��0=��B�L����D��rL�g�XH<��Ƃ�=��X��@����Hfo�F[!�d> ia���`��tJ�NQ�b��yR�do�,Y�U!l\�dcq��zB#"O�(H��0;�]2q�Q�m�NDX���_?�4�H��:�L�i{f��a!�G�X*�"OyQ�۴[�U����+��%S��Or�=E��M��~]��)�,
��
��^��yR�mZ����,�L��m�5d��y�'m"��B�H���r���$�yrL
V��xp픩+fpK@J���yb$�q8R+ֳ9ŰcGnW��yb�� Z�Iy�"Z406�@g�3�yb$��y����%�
`[C ���y�N^�wDj �&iٺ"�ΙZ��]�yr攅�R�3c��k���DV��yBO�Q�0��L5'���r���$u�h�>E�o�mj��aq���"��C�͌�yrnJ=NlЬ@��8b0��%f��y2�]U^@ySm�
�@�`����yB&�>����4��qyCG��y�M���m*l�5}��D �����xr�0'�u�K��V�A{�
���hU�ē5�y����e�&�h�>��P���L�ᧉI�Jc�S�<K�̈́ȓ<��U�-U�v�^|����D]Ф��\.��QEVxm��J'�p���&�������x"�EF��	аgY<� �Qi��n����0��0�	M�O��I���r���R@3o�J݃"O����h2T�2�`����f�d$*!"O�8��F�+�ݸ3*^�/���q"O����P�J�̲�i��YԨ��B"O�,�ŋ�	r�a)�hݑrV���"OH9�����hʛ?���"O�衢�K�:���&��&��"OƘ���1ir���k�(uC.���"OZ�k�I�#b��9q�C.d����p"O�!pł�4A���j۸�d9��"O����@
.lJ�:�`�"�Q� "O��T��o4~!8��O8_�(���"O`�@e��F���`M�P�����$LOBِ��]9>i����f2N��s�'A����`c��г��)��ҕD%D�X�s�G(���3��
�H$�E�.D�8����l��F�F�qGRH�c.D����ِS��<�h��r:��Pr*&D����;[Sda1NTb����B)D�xk��)4e�rG]6O�tmcD���ԅ�I�K�J�ӱ��N_�ai#���B�I�7��sb$�D����Sk��NB�I5 �h 3��ĕF�h$ϗ!�hC䉃*(�Y)&#K��1 n�8G�C䉒*�1A���*4 8L8b�Wq*BB�	�l���i��� p#:E8����nB�I��Y��DO�_,�RTJ��hB�	<p\�S�a��s��
ƣ e�C�	 ���#@A1�����/d'pC�I X&1!�)؀��ls/V�F�fC�	;Ǌ�1@.ӍDI^P�AA�h�C�ɪd�8O�_� �õ�3i�C�%Y�d ��;���ޒ0�B�?2�\ �~bb�j� Y�P�x�If؟|�Ҧ@�rm�5dN%=�����%�ON�Q6j�Z���"N�,�U��6���ȓe�`8�V%�R��c��N�dF ��'�ў"}�E���b���e�
��@��
e�<A�P&}\@,��c�j��\H#_�'�Q?��Ν!^CPe�I�kD��[��2D����Ɇ"��e�5셛
��ъ�O2D�4"1��*f���5z�����ɵd\!�d�IޤxہU�J` ��T�fS!�$��[Ԥ�KJݏyJ�e��/K,n�!�6�^�����w� ��Α�,�!��R��`PdY��8��nպ9�'���E8�D�s��O�|P�)�!:Bڐb�'w�D�3SBT2R����b���N�!��S�` ��A��n�$="un��!���\�����d������<>!��Z0���W�3�,��D<ONa{��z�	 k��b@�8}��qG!�>B�I�o����� 6&ʨ���� �2➘x���Ny铠X�i˱�:f�����B3r�
��$^~��3'b��`n�"�t5�eg�F>������O>˓ӰQЗ��2��e0�J�lDyB� �S� H��;���\iE����$b��z�D��]�ꌚAm��3b��'���';ўb?�sߴ#�tq���&2������B(W%�i��{B�pӧ3*as,�t^����V�r��#o��:����T�GB(�ȓ+�(�j ���H�0�󃜝\V@��ȓ	P�lQ��
� ��u�g٘���S�? ~	c&�Cy(ΐY�閿(�T��"Ov�"�
ц �zˇ�����"O�M�c(4R0��rJ�H\���"O❚�g�o@��&�|J��[D"Od�t�Ϩ!u��a�ȏv ��"Od8�"��mw���!�E�b�E�T"O<dbQ ��9��4�	�I/T(��"Oԅ�BAU�VȂD� ���U�$�"O�q�d�--
��''@�1L&�Q�"O��*���J_T��cY7H-9q"Ob��F!�8".��ցٴ*����"O��b��W�#�!
��9m�1w"O(l���H�ab�yү_�X/��"OL�
���.P���HM�$*"�au"O�	 A4
d��;UEܒ5���"O�J�L�z�|B��,
��w"O��K��A����c��|Z�S�"OڐXe*��$������'a*��e"O�-��CӛZ?��lʷc](���'�Q����G�&��W�����(� 9}�)��8	`u;�L���`Bc��:dB��V�Wb�0�A�/_w�㞸��	E�Ez��/��q��
S��C�	)Ek�pC
˗:��2���2����'S�8��*R���l�5i�&*0��H>y�A��97f^,,�Z�,��["�̈́� ���aE�f]~�J�B�J)��Zn�k���*4��d
%싚r�쬆�� cDX��>���T�<����.;�u���]�x#�BO�f,2<��):���f�	�PHc%���es��ȓ�.�t�ޓ+���wɰWg+D���NS��P0�0/�D���`<D�4#q+��k7��WO�*��#q�9D�PP�2F�ᢩK>14�`�t/%D�Pf(��촋��լz�����*"D���%L�"�x�L��)l���h%D���p!֨7 ���E/���`&*!D�x�ᏑA�,DZ���"�~8h?D�� O^x� P%���y]�&�=D�D�5�ژ���f�� ns��:�n!D�� �B�l]��׬�#�*+ĥ D�DC���0�� � 0v=��zGd$D�h��&��%��C)N���M"D����*��R����2@����
6D��2G�u��S�J��r,��	1D������%��re��iAL\���"D���JF:	�L�d���2�;D��3�e��3n��+PMI���ՙ��&D�x�蒐T� �;���X�V�X�G%D��wk2V)���b�ł!��i��8D�@�v�V�Gt� ��_�Aq� C�9D�hF#.P�0��$
���N*D�|����:>�`�[c��(\�d 5G)D���um��D,���m�����Rn9D�� i�.W�FJO��2w���aN8D���Y�"!� ��.b�(`���8�y�@�:J�R�2� x�ı�%o!�$12Q:���9�L�{r�	�&�!�$ԫM��0`���-n��AV����!�$��FG��٦��?�A��`N�(�!�Dފo�
�k#�V�½@GOBs�!�Z�%J��Į	Xi�Q+K'5�!�D]1I3��1�.ßM�)bϋ4,m!�� B�[eM�t�����.�t�!a"O.Y�L�yONa�C�+6^d��"On�2ƩV�	°���h_>ގ�y�"O4�PC�8?��ȩq��^�:{�"O���Ǯ��)(�|x")N�!��KE"O@Y1%� :�(���� x�����U�T}�a�w���3�@'z%�a�LN����f$D�l$�$<�F�p#�t��-Q��%D���QF[�x�X���^*+6�}J� D����u'ba8�́�JS�ڢ!"D�X
�G �`	X]�R��s�Q�K"D�����${�j�S��C�(j��"D��R5!��Q��\�4I�~���y��5D�PQ��W>fBd�� &�#�"6D�@���י'�E��.��l�T��	2D���օ�)r�B8�ů��� �4--D�lK�d�t��(�*�2r�b���M(D� �d�<WK2�
�J�?�|�	G$$D�9��BX���W쀳��U�1D�p�!Dɡ�,i�2i^� �,�&'/D���a�؊mՄ"a��:�|ႂE+D�(*�J�˒�Xv̛�ږ��a�/D����Q��|z�LU'SU�q$,D�00C�	#X(�AӬ3��!��+4D�P��G�-�@����
I�M�d�.D�p'^�ʦ H��ف��� ��:D�@ i�zuI��"Dn|�C-D��Q��5)�]

T:_�eP�H=D��8f�9=�%�elXc�^ `!;D��J�n:R���闤W5ie:y�%�8D����e[�$��Iѿ^�"��Ħ+D�8��Z�dq[%c�#�.$;�k(D�$)�G�22��Q��GL*>�`��'D���S��$�P������%%D��&�_�?�PY��n��]��	��G?D��Ӵ�F�"m��n�5p^��AT{���DM\�D�t�'���S�ڏ#m�`
���3�=��'_R�C@"�7'�I�9
�P;�y�m�9�X�E�<���������Zr�n�m=���&"O6�j�f�l�ȂK ,;`Y��ӯum*,�昀-�6-�,I;�?�'
%���;ô�Q���E�x��'�F��b�*6G�1!�M� s�$�S� L�-�P�ZDےA�g)�<԰<�5�I9(��&�̀&3��V��s8�X�3Z7
��X�@[/d�h�HnG7)Ҙ5��,I6,M��Ff�~x�
�'1���k��9n�(�.W���H�0Z�] %�,Y#Aw�p�CM��1��:O��y�6�	Q�G����"O
ac�႓��i��l��X�2 �WQ�P6��H��x��5�C�xyq��Ԃ�Q�8�"B�B��qC��&݂�Z�`*�L1g�޾@-�E{E��q\
��B`��S��7P���G'%��=4f>���A��v̬ jqlJ-g;����I�`���H2.��وcF�cNj(7&%R�8�#G�#���`���qg���M+v�Bm�w�ȣhjj���
I�	U��F��ȸӁ�Q��5�+
��5At��M�b��d��	J�h*`O�(ojB�I�[�-q���s1�t�c͌]��91A��@���Bǃʅ0>���
>��38��'��%�p�F�*�!6(6 ���|��H��بr&���Ůڅr��l	��0b&��B��M,^�aP'��5�F�I��6�0����a�'��<�?���"g�
8(�d�1 �d�@?H������܎8ԍ�0���
(9�"�L�/��5�&�!E�xh������!'�a��@@,,F�I���p �-z�4��'u����V \F(&�	A'_�l�(�ȓB��s4�
7�`��b�;d��Dɿ@,"ӀIy v����W^�}(x�������XU�Vf��csJ_�^�����/�O��h%(�����3GZ������Խ��p`q	�-9|�9qQ�		L�X�k �L��Q��!��f�� "J��n6=��h?��>�S3(ݫI�i�l zkV��� ^���Z�aO�mp��	i�؁l�eK�%	�t؊���ܭ�8E��%���x�'�^ڄA��<$P��5%���A�˄�J�yYH?q�PÎ�@q\}��=	�R�M"D��&�ŬQ
�u � �=���1��l}F�bU ��'��@�M�4v:��ԛ�k͟6t�Ę�gA��S+{�j��B���ү��d�mS�L_2�B	��Q~0 Ѱ���q��qX�ͅv�ס	��I��ÀQT %A�,J�8�h����=�ax"I	�dV��`�Ҍpq�M�5��-�&A&��R����$.�Q�$�S&b0��	j�� ��"�.�"1��R�[���'_,UR��L&����m_�e~J��`��%%[�H�O���[�-L�s!� T�ҰD��=S�'�$�� ��8~
���o�;Ey�&*S�{��S�/�@`�cDQ'm�q���	�(S���./K&tU@�B�7�0�I�A�ph<�5(�d&��C	�'t�@Sb��9e�D�R� �1�D0�Ϸ"�̵��-g4"=�bV-hS��W����v��o�����L�HWrl�Ŗ��ty�`�H�Q�d��ѷ��u���Ӥ���XuMA�O�|���TO]s�`�*��i�0�����'�2p� �A!U@~�"2[� �zhqL��9^y*<j�AرS������,�C�	�}o��ᆪɲ9/�܉�a�2���f^m�� ���acࡃ�l�c?]Иw'%�%�3Al�Ɩ5e��,�
�'�,��p�[0����F`�  ��ÿ!�y�e#�D�He��σ��`�Z4�O��!��OAi�P�BS�+�j��u�'�l���i؟WԦ�q��/}�t=H� �rg�e��84՚'I�'����	�z�P��aC�@y���Sl@M�=��$ެ�f��4���'`�8 ��8K��1\�YI����
\�EK�@��C䉪N"Q�K[�}����`�&a���I��������I�]z�kX(J.A��	�7��b��ܮL pA�,G�m�!򤌗 ��щ��*g�j���ə���Dq�	]KvR�j�mF(?��ݓ@�~J�}�
R�)��i��R,n_�DYda���?�Õ%+Z�,S�`��&vp0!� �ƴ�4���b4�g�İ��&<]�LYUΛ5�X�`�4IV�?�r���ku�p�l��c�6ih�Io��B�*&z6��8���0R��C�@<\O�d�̔�#��	�OyZl�7	T�3�>���-�;PG��Q!��Ģ�5�^)	���#}�V)yUJ5�I�M:%q"��I̓
N<5QbA	i��?�:k��"����4Y�'��-E���(��*���؀nR'� ��qOȼi�"^o]T\ss,ՏDlp$: @L�-���E56�V�X�&�# �b?���H@�3j��$*�]S�1)��+;�,�z��M�T탅E��f]佢�T���i�%
lrĘ��ɘ/k�\���_z��V��_����J9Ch��QХ׊lrج�i٬m�Z��f{Ӹh�C	�?�:�"S�9g'褫��+O��ʐjL32펹��n�,�
�`ce��Y���C�Z
n��$�56��a��y�<�� ��)Lܠi#O�y���_�'D�$���fM(L ��bG��p' E�OB,c��Ǔm�Xl�R�2Pڰ1���3W�f�vnĤ��t�vw�mʰ�M��U�f*�+���I7'Yf}͊�Qo�D�}&�0���i�`鵦��+���3a!H�j��T�f�LZb�����;�,�F�MG�TP6s/:4�1im��v���P�+�Ǘw�x��fB_ l��(E�Ap؞�ĭ�i;`�:F卹����u� 8���֬g\ΰ�P��=�v�	kC�m0z�B��;
����M[yBi��=�i�� M���D)U��O�hz��K06j��R&Rt�d�q�Ρ|�^�8�%�l�&AdS�-�(��I�EUĤ��q��H�#H�<<�Je.2DY��ǲ<���U ��x��ÜL�p����L%�q���T_*�4�O��cŨ
?z� C� Pm�'�e��H���l��ӰD,��.�%+�ʤ0i	�a,-��ҺR�}��X?yp���'�̹�;]V�$Q�سD�ڔ1���	d*0���#_P�Ӳ��t*��=D.��(dB�.
:$<��(Ȧ&��+4b��E-���p�0��HR2����@���5��� IR�D%Y_�z����0Xџph�R5-zA)��5D}�P��S�k���,[�lA �K̚Uߔ�����7x�|V�T�2��e&mӐ���(�{�x">�7E�5NvX4&��#���*�e�Syb�Q__����Q
A�a���L���	><�m�$�r^ɨ���7!҈ZSʇk�,x��f�!@CbM�7�x����!Chp� ũD&�@�˥�+/��(Jt���V�T("iոX�v��� @lt��酃!�V��E*�)+���14A�|�$�P���퍍q�pX��	;���cvJ|�V�J�Jz�S bF�HXp�DW�e���$�Q<'�A���tOh�k�@�Mu
�+ЂߘA�VdW��#.�e8��I�}�$���0|ў�����F@T���k�(uP��͜��Pb��y�m����'��y���C�#�Kˋ>�ؚ4MSL�2ЈFA�|�֠��J���'� ���O�Jj8%�
ch)��4\��E�%�	�$�0qy �#T�u�%i^�Y������b�%$]�X� &ĬA�����P1���R��-gV�Jm������		l.�c���o�9%�ݸX)R��p����U����1U���B�
i(�c�jY�n�
=��w�~�8b�I�@.�(B����EO1C��)VH"�Oy{ ؠ
�0�K� �haU���%�6�r�f�:y����`�Qjƥ0rjB�2gډ�A�n�xy��!�$6��;s�6$C� �.�ļ��L\6Mr@u�B����p�qk ʓ����L4HxTQ�2FH���l��	�ک�(W�Ůy���gP�h�E�˹I�h���[�/يԄ��US�U����Ќ8���Q�x��@��4x��#��	~��G\�V[�y�W �> ߒ�'�P"}���ݱe3�9�2e�Y�)iF�ث �C䉧 ���#���du��I�� a���-*�5bs�YC٠��)J�7��Ԣ�2��Hd�˻O��!�w���X,�*��"�:yh!��*����K�rrn�����1]84��2Kp�)ї`P1�^Eh�Ń�")���'ޑ{)�QM�2X088���M>A�i 
�v���qr���O��c��˙/w��3�մ<���kӄ�W����r��<@A����#�Vü]�t��'��{���k7P�Qu�;|Odlz�n����$_) Ĥ��j�u�ȩ ��˟yM���i�b|J�n݊�����Ğ�ָ��*F�#u͙����b���+\VuR�b�<I^�92�"I����ꆆ*N��y�n��M[4	8�N��e	�>�7BljD��9�X���H=�y�*��|`�t�"غ'y���p��0>�CL��@�%)�<Z/���4B@�S�z7k��n��m���	�O,�ů!u�j���˟_&���d"�=S��0x�(m՜�����_����"�y($H�(Th߈���$�]���	V-z��@�>���!�`C4�̅"TI7Y�Ӌ؟t  y�L�h��lg	
�7���I���fx�����6p���PC+˙P3|qR�'�+0*^�)J�6���c�&aw��B"E�r��(r!���h��8�/�*<ɘIQb�"D��DB�/XZ���ן򄨣�   L%��� >x���ɸ$�ԢH��4:t��P�;� ��`;��D)+M�Mb�Fğ�����>\I+�!�f#����gL>E<��@*����;�b��nt��c�#`�L�����w�L0	�X�L>��'r�}�֦�s���2��Yv�'؂���I��b���1&�\k��f&�t���S;܅ЗG�;

y;�� WF��R�	~}����Q
ZQ-B@�~�h��
�^����k�����I!�,�Y�V 2�ܣ%Q~
8K2��'��9��:@,����{�<�F�V�<A�p� +R"Қ�kUM�\�DV%9B��7j�<�����GH�|�Sd���'Y�m�"B^�< q2���o��)��^JD�6��gV�L��ʃ�`��U�E�e���PV%m�Zi`R������f���VG�� ����EJ�����|F�����%8 ��%�N
 �Ah�;_3 l��@P���
��=Y��1tْ�KW�Qh � ��M8�lk�3&_Z���¹2�$�*��q����H HT=D�!�$�%�@��� 虚f֗:��A.�{��/(x$����h�O���E�H�6�.H���M���|��'�D�Pˈr=�����C��H �ս��0�3O8�!�+O�����84�u"S�Z[� �Vʸ+�^]���~��F$���!� 5��]X$�TUxp:�/˝� h��Y���"g���"�a�3~�&��\�82���E�h��y���'�fɫtE��w���)�Ιd�5s�'.�4���U/q�XX���r�@�J����"f촥��%Ř$Q�}j��Ć5`�\���iN�e�œU�<iU�^7Ͼ����:��|� �U��@��K}2��-'�b?O(��N�i����!դL�0� UO�L�"� 5.P��#�3\Q�� ').� H�b�X���|Z){�d�#�.��4�Y�Uw���AB��p:��Jj}R����H@
ǃ"E����S��y�*��;��%G��I4�ɹ�h����'���H��<H·+��D���R#�0�9��"ONTqG��>�4�T���=���"O�D��[c�)`��>���Q�"On����%4�^� ���b�؀�""O,@B�O�#q�H��f�Z�m��A�p"OnT��⚳O9����A��ZGB�{�"O���sMW ,6�"��#k��<s"O
Ib��0�\�!nĴS+n[�"O�]�#�K���ȍ�y�"O����U =�hA�FOq�Na�"O8��B�$ �f]��Ӻi2l""OfeА������!`���L��"O���Ă0u¸���p�u/^�2�!�ĕ=U��a�P��|�f.]�`�!�}v\��7�X� w��E"ƭa�!򤉃]G.����\�cl�ФO��C�!�� ���k�7hr�b#D�|�z��'"O������k�,���5h��t��"OLd�IR�1Z@#��Ƃ&��A)�"O��8��4Y��ҁܡJ��� a"O`@�g�؋tU����4su�ً"O�Au	@Z+.��F�E'	�d��"O~�1��$�Qqs�C
4��b"O�L��)�4�U�7��3F�%8�"OL��.D���9!v�H&rqč٦"O�HȔ�å'N|�r���0p���"O����KGJ9��Z�����PX�"O�²e�} ��s2�_�;�
-��"Ox�XG��5i�VT�Y�`�H9*�"O�q� �үV:���3F["S�^|�s"O"��-88䭠R��6XҐ(�"O��P��~�Fe�%��`�J�a�"O8p���.!㤘��	<z�|�"O���?h&�D�$	�j�İ�0"O�,zRB�*���QЂ��;���A5"O���O8�F���+P �X(ҵ"O> BL�~�I�7�1Pa��Ɇ"O�*b�A6P�䡲�dN�0x9{�"O �)�nb���8޼��"O��C��J�$n�z�Ȉ��=A$"Of]�Ao��s�PD�`�U���*�"O���q`W�M��Z�C�/2�le�b"O��h�	�4�,����PP�Q!"Ob5+\�h2g��e>}##�r!�D�>��,W�=Q@��Q�կZ!�D� m@x�zǅ�+Kތ0��)<!�Z��|H3��B1
�L�+�
!�V�3�2��V�4nŦ92$^;�!��9��Ju�����qBNݨq)!�d��=��墤�q��LQ6-Y�t!��xC�M:������@g�S�H!���>OZh��F)L��LjG\9'�!�8/���F,a��A�`J�|�!�!_�lX!eS�T���#/��>�!�־s��	��
]�Q�O�!��IG�ݛ֮Ȝ=��y��)k�z"G�v�*�RPj��Lr�-�d>���k$���)��9D�q��< ���l/)q%�4扯 *ʕQe!ԑ&��#~��� h���ĥ@9*���S0��o�<a[��NKr��9��sbΑ� ����iD�%�E�۴sM�-"��L����M�o�Љ(҃�kd�ϐx�-���pȘ���1LL=[�,�5:BN(�a�G
���)�DԲW�$T�˓�K6�ܨXv��ٲJ߄��؆�r�n�Y�G��y|��+�E�X�(����E�.iS��ʛ?��K3	���Px��U:4҆Mۥ'�c�Jl�w�K#��	�7�6��&��C���
��1j���{S�؞r^����C�\����V���b�!�X5� DO3T|��VD8�R�#��D��u!��l�L�����\�a'剕�4y�T�UHP��ʻ��C�I�N�-����j?t-��`�(i��QM��a�<��0���2&��W��?�*Z��4-��Inx�-�ƥRr8�0���6#��IG [L�p���%�m�xC��U�����`ڑN�@u��!�Op��C�B�}rf�٦9� �ҙ� �2Ix�=�D�0/bT��� L�$4'?���! 5NI��!G@#��ܨT'/D��qS/�?02�r�ª:=�8��Қ0���{�� � �>���C�$2��(���ÏayB�ȑ� )�u*ͻ)�������?�rj�(�k��6c�x��RE�#T�:����?@?dUKfl�)ZzEK�"џ�J���JO&A91��(Ɓ/��J&!Ѵe�YE>r�Bل9��p�'�k`�p#SB�?]Є �̀#+�1�&�'�Đ�ө��b"X�S���b_�M�,O��P�o@���A����6+�H�w�يU���H|R�JJ�[�0ՈP�=��V��J�<� �C�IO�F�r����k��4;�K�c����V���X�F�ΰ�O��x�&0�~�@��57�`����m9��i&��2��?��Z112��ЧS�-	@v-0I\T<���B,	r$١!"P�c؜5�tıO:(�F}��?g�I��Z�S|ƈZ1�D��O�5kT�޽nRP�aӊ;Z��0oX3[,"erTaR,�@ ���{���U��'E�~��8:�����m0$���S!�����6ǂ$02/�;�	C�nO�2�E��	'����C�扥q��$15Ƒ/�ʥ�ȓa��P�,O��Q9��O+}�8a&�у
*N��H��Dw戲G�S�SB|���겟h�v��$ݪ�+�!$sR�w%�ORd�jø&GŇ�wX=Y�^��b� "w[b�_���s"ϭl�����J�I����� �m|�Ta!A+y�ax2�%>XE��ˈuF�K�'8��M6j�=���"�02�C���c�~$��	�]�Vл�j��K=ĸ3���O��'�|�A�@�M��)`+��Bq���Ft"8�O�\�����)J+�l3`�	�'�b�� ܗ=����d�/G4�7H�+{�Q���G ��BD��}�q��t�A��S����,�e�|(`H�P��C�I
6Tnh�g����0�O�k��9s�Fx]NNO1j��LҦ�@�7Pbt���� @�+	6g�Ȳ��S����Dۃ1mj�C�ɉ��4y��$�<;T/�2]:��p�S�4�+�j�1@�J�"�|�֠��C�t�R}�t! c�m�=� �ΰx�:���&�M��[E�
�	��G؟Zi�b�! d�Ѓ89b�h��"O��'�iKP��D�k�(���[!m}���&dĊL�P��J ?�����N��{�(�U�4$�x����Z�<�L#zD�٥�1U��B������,r�Ĝ^�4������x@������wD��C`\ Q�L]�gdJ���>�WĊ�0)qEL4�6�R#*�M�AM�gE�iӠ$� i�8��b�f\�ۓ �5��N�[7j��DG^Y�J9D{�@@uJ0��"f�+2�ɧ�9Q`�;)C�5��ȋ;�l ���p���Bv�p�C��rx�/�	*?���=GU�1lFb�|��"��G�h�c�0Q�z�u��L=��k�b �`J>C�I�3F���b2pn$*4b��3G>�B��.Z0wa�#A+��P�2�$���=��YaT�� ��҅�v}a��@|�	8�L]�wN��#�_�x�,AT!KU��9�A��:�%�ۓ�X ���G�d��Ă�3��G��˅q��QNӈ<$�H&.��Ӓ�۝o��=B�N5�h�Q��u���m�;[3D�H4��s��o�Hu��瑲NJ�'X��EM�@�A�L�z�ZEE��DB�>xt�D��0o����U#��'������O "zuG�,/��]rj�@�~��gI�Qz|Ẳ�ݤv���(d	�)y�n�%?� k5J)Z�͋�l��N�6!
�ʐ�U�N�ڀ�X�����doS���~ʴ���@�P�R�MG�r��dL�+�RL��KP8u�b8�A@ƹL�ʨ�@�'n̐�FM�,J$��@)�@�����8j��BAĳr�4�2�T�z��ݠ�M -Jcw�/�X���.�ͦ�����nt��f
<&���׎�o8�(����-�^� fJ�:}��<r�A�u�H�S�&򰸡a(F��kGM�9FT�@YB�K��l�X�K�1w��˔��OI|�u�>T�tYK�e�$=�ՓL���n�
Lq2�)H�#�����\�h�ԇ�2{���S�����N�'c�0 ���!a*0���*��DX�?c��L>�2�_�X�V5+m0����ԅ,�yh ���hazq�b��]�JM�R@������=���Xc�,����ԡC�ty�l����� Ŏ_�F4(W'��=���])b0jqB��Jy*c/`�@&�֦7�Ha�A�U%G6-iFbW�a9|E:-��X]b�!���$�6A�l�C5r��ą.�џ���_�f�	7O���Hcw�ѽt��0��mǦss����FG���!�jI j�n@rG����=�S 9K�xf�P8�>pKg�hyb�ٰ@�  ��\�H��Q��@8�%K� 1	��E�D����c`�џj�I���K�\���2"Ol#�[+d<=�� �����(7*W�e���:� �?��!��r�~�H�~b���^�v�s�w�(q`�:vQ.d�R��3IT��#�C�49���U�#e�����Ϩu��<s�
�4d�� �Q��z��2�j�Q��Us�j�O�]�W+�~�K���q5��"JА�d�;��O(�s4��N}�PP���<�8�z�'C?"�D�Ԅ'0�46͟�	��pT���LI\i@b��Ӧ�[Eaң�`xF|�\+CC��� ��60P�1��L5����]�b�(�&ݽ5�tqgj"+*��U�Əj��3��r��qC�@ 斞4"�����"m����Ңv���d�~��=(gAJ�.��Ya��34\��7/� t�H��aM����+Cř}��=0k�hX��:&���̻�<881� Q+��)����D��Ʉ
�2�@%���� hYCv֑8���
VfLQQ���Ed�]�1��m�������Ј��Dyȭ@-��?Q�j݃00ё���zLh��|�'���'�VX�A�A��ʕ" F!O��鈖OՒB7�U1`<M�j�$h[n�F14�[�����χ�H���=� ���E��F�\�p$��� CS�|r Ó7�j��M&3Ai�LP$�$(!���g"����=2�Th���G����O�M�������S#J�h�cǊ�q��Q>~B�a��,��b�h��Y�rw
ћ���M���2� �g���yǇ�}E�q���g�)̻S�(l�@�%Nl��e��j����R� t���q����S��w9j�kF%�jčb�JH�:ب#ǿa]���faݪu�����4t�h��,K�yr�9ټ���*ӄw�B g�S,�p<�fj׫O�92q�\<J��%}Te��F�!rf��	�FF��-Q��\`4j��Blf���=a�,B���lS #lKp�'۠ Ƙ��� ���C�K�7k\8x�l��r|���'��4Rэ�K� �*^m!�D ���֋Y�u0�)2��ڹ1TN�!r��b���!��Y�$���kå�#���pU+�j��[2 �5Ĵ�ºB�V��%(D�����ʞK��]��EŖ}<�"�EF�mB�̑��]OZF@��ЪDVz�Ɋ�J��M�?!���?$b�*r��L�
�YIx���Y'f(�K �>>v�֫@'>�YX��m����V�h�T`
ߓg�<}�b�_R?��*g�w#�uD{Y(Lآ|�G�Ռ:��e�u��w���;3x�xc�&���2�Q 1>]�ȓ\�jI��=9����@� D[��ϓuk�)��ܟ�98De�=X�d	i��?�'�ֹ&aսC�=�Um^A��ȓ	2aHAl��$�	�P!?C?ެ�a����bZ�A�pn�#dL�O�㞼v��'g�&����ÎKʞ9��l.�O��asl�*oH�3��H�h5�M�*'��]`�E�dD�`����*Հ��d^�4�8 ���%.Hɦ��$�џ(�D�a�
D���Z�<`�l�WfͲ6�l�&lF��T5��D����ȓ[�� (C�Pe���]�qؤO�\�5�928�ȡ�P�c F�Ħ�K̢@�`+Q_����iS%�y`X!沀��E��Q2B���)��NJ�-4�l��8LH����|�T�sM)3�&:4E�uXQ�ӎ�Px"�Z��iZ�@� �A@��9qD	j�.1���U�"| ��'r�pBA��tM8�)�K�`�	�@V�)����'3�4!ۥ�D�.� D��:��1
�L�
�ʤ��$ D��[4놃n�z���/Q'/h�E�?}B��#MW�,s�*��|�v�X�>�'Q�2<xbB
t95z�,���ȓ>n�)
p��8��e
O�#����Y o֔��o~��B��Y����g�N �GH-����/+9��`�@#�� חdO(�� C-�lQ���0NhA1&�/4�"	ۓ3	��9b��C�0� �I�_2\��	=ld(���; �\`�0��Ot�3@O�"C�2�ɔ�>�ѩs"O� �anW	%s�K樋eST8���>��������	ڑc6��F�DM�ds�H�HGC/�)2�٥�y��V��QYT뙗=S�y:���\�b89u��G�󤟦������L>��L��	}�Ԅ���� �v(<q�[TM��
=j�t��ǤP�^\� Ŕ�S����a�g��0;���~�P0s�мU�0�A�L"O��30�MF�@�������2W�Nu�p/�1A� ��M+�yb��9hB):s�C�;P��y�/(��s�4�c �T��L0'-�'��<y�C�)2ܽA���8�T��ȓ �Ա�j�F\�5L�y3����P��'�q� /;�3��#,�
]�'%�G0^���c	*z{��$/�X8!�J<y|�`ŋw���җH��Ћ7�'�5��� �q( �0h$S7
5�
ӓ9U8t�R)���>߶�З�d��MU�S)�0C�'bq�(jR�	r	�]sC �-L㞼)����>�*U�0]�`� ᫃�)`�q�v�H\�<A��]�")�̕>�v}[���[�<�K�.(v�Xs���
5�Z�@�\�<�e��C�V�b��H���7g�Y�<���E��r����A-�X2w�EU�<��I�Xf0�)r ��~G�As��t�<Q�`���8 ��)�E91TM�<!��W��­K���r�va���O�<q�,6q� 9)b��`��*�jJ�<ԩ4/zY�S $p�d�`@ Qx�<�+�R<>e�ƨ�˚�8�$X�<�vȚ2KΜ������Lȶ�_�<� ��0D�ܞg� �y��,P�	�"OhҠ�K/C�@!��G�Hq8"O΍�"��Ak�}eGʛ;�( �"O��
W���.�Z��Ӟ�Vd2%"O��c� +垭��Cx�@���"O������E�ƹ��A�H��tR�"O��{�I�;�H��@�I� ;�"OT��� ��]���9 [��h��"Olȃd#��#�|\x"�>N���"O���BÊ" ��׋Q�#��-�'"O��!�¨:�9�ㅉX����"O�ي����:h ���6���q�"O�%K #�.r;@�c#�L�h�p�"O����V�"�~�1�2|�T,
q�N�j�t=X"̇��%�Gh�by�@�p�O�r� @/L�|��V1p��d�1Ǌb��ʔ�>~Zb��ȟp�����-��K��8�b"W��M��'������*'�>�}""�٬	��9xĚj���J�D�Hy��]�j����5���Sӈ0�0��9��_Б���O�4� �����O��}�V�Y�@�&	�SGŢW�>����q�M�:tV(�'��\�>YH�#�aHnh)��Û@Fx���T;��T��Oț�0|�DNJ"U6�=[��� cg�0N��z�:M�掠�0|��nب[꒺r-�}��%�qy�NI(K�ȱ �!�$�?Mٴn�T=��BܧkG"|ǆ:"��)��3|,�y�f��qm��+��O�Ḑg>P`���chj�:�DR�oNЙ��@�v�Q1���M֧0|�O�u8V��uD��:�V�wB��8��R�C�_F��=KF�����"|b�ĝ�c��ؓA6�&ԳB�Ú&M�]2�_��@�J�j�|J~�E,k�D���:v�JE`'̚T�I�u�T���n8�)�<L��E�Rl��0��}R`�@�,��	b�����B�)�'�r�`r"�&�d�Y�	Խ~�,o�ML�
�D6�)�uF1�Ɋ�\� �"�?y�� �vN��|�u�J2@/`��'><��铏sG�Q[e�eY!B�4{|���|2b���M��~����J��᠂I�C�3qm~�dE*&�`v�:�#�'�E�����zrjP��!�C;����'�(��7��Mɧh��p`gls0D(0�Ϸ #���\�6p4t��4�ē�0|�����rJZ�lL!�c����ܐRƇ�Z �Tb�|b#�Ǖ2�ui<k+����)6#|OT(��?O�?Y���(o`h*F�p�\l W�_a?	��i�`0�'�ms[r��&���>Q�J��h�:�r���A�f p PQ�<�ceϿj�JI9qF�u%�l���c�<I��ٴ-��%02�|ƺA��Jy�<Q��z.H�ۥ��<V)�A1w�x�<	eA��#��8Xbe�K@,iy�"�w�<i�ʐ�0T ⪃5;�D��n�|�<��)��n����l�0`�<����x�<���HVH��.�)uTy����t�<�%%�ri�3f��0欢E��e�<15�S������ɉ���beɒl�<af���9�7C��#P1S��~�<����n�%R�	m9��E��_�<ѴkOpĠ%�R�L�F��l�� �U�<�S�ƨj�" ����j�i�"�)D����u��e,H9R�U���(D��C�IC>+��dB%�?T�D��am,D���5H��YE�%/I6}�c�*D��
V303P$���� *���	w�+D�X7)��~ �d![(8B�)G�(D�\�����g^^��Z~�i-&D��3�@IR6yjwc�=p�p�c��9D�( w���_��h�uY����g4D��kp��!4�J05j �\0�AsW�&D�8ڃ�ڑ~Vh��[���xE�/D��"��$ ���l�Jn��#3D������=|MZ�1B��%�2ᒁ>D��"	Ŭ���q��0 �H�8�H<D�� �u��	�* +�����*���"O��K1�S"���suǀ�X��qiE"Ozd�nVv� ���k��H��"OP�2��_�E���f�]��`��F"O��w��;8>8�P�����zb"Ob�sWm�$b�L�3���<���"�"OXA��V�Ih&���h�!
���"O@%���2S3��h��_zL1�"O�Er%F]�d����f��%��"Ox���+G/
�tEE0{@\S�"O�9۶�
@���T�U�|`^\hT"Onq�t,B+hyh��V#�`{r���"O�9�B�M�6�p!@@LV��"O��9%��$+��X� �^	G`�q�"O�!�猐2�����ߓ`B"1x"O��˱/�#*��2���;!X��f"O�܁���*�y�fO�y��"O���ҪP�"��&�
e�s"O���+�1�0SJ\"r<<D�"O�tSr���7�$҉ҍ�4�	�"O�M�!�ٻ��x�3B�%
9p"O.�2%J�kHj0�'�5,��"O��{�׈d�p��V�R�*$"Ot1A�m835��J#�Ub؆e�e"O�]0�✱&
�3s�[�Q��,s�"O��Pw���a�(CK!o�T�v"O�  t[8���qM%o� Ȃb"O&��r�Ý .�cu
;_z�H�a"O̜ҡ�~�u�b�Oy�$��"OLp�$F'W�ڌ���=����"OVL���Ar�(���B�80P�5"O���r��r� 2c��*u`�3B"O�xk@��vq� �&q��@"OV,��L�D�H��¬i����"O"8�L�|iT5�P.P��>�ç"O6 :�$D<z�8�k�&:$���W"O�a*
�{��h�`�D.y�*@[�"O�[���|�
P���Ŧ }-h�"O��a�eU����j�$@�N�g"Oh1��88��}sE
�#z��"ONіoV�j�X��T�v]�Qk�"O��r*�/k����cM�b<Ij�"Oġ��oí�� R�C/!LP�9�"O��4 
�E,���zg|%V"OP	P��k�04V�K�&M��A"O�����P2_eɨbj�2vI�d��"O���IC)?�� �&�71��q�p"O���!��k>���ʞ,�\`U"O�r(ڞ)�8�$�B:
�I�"Oz�X�E����Iۗ@�9�"O�����!.�*4!��Bo�8�˳"O�mÂ�'���2* ��>�q"O�K4l��tU.����._ ���%"O&���*
���
���"OP�����RO|t! �X|� "O��� O$j Q�%�v�HQ�"Oa1�cZ>L��Y�V�� ��R"O��_����E%R�HA�'qށANw	 \�靾r����'�����,Cm���@�c��9Z�'7ؽh�K��a�8Q�DX2�k�'g���d��Y����3nѷ�pP#�'��U�D�
�G$pڑ�[�H�J�'�bp��U�w��5��-��1Nz�C
��� t ��F�#3��IL]�Z]bU"Oʁ�@����� �@@�Cg"O`E��,٣b4�,��A	�/��ɫ"O,�A�H!i���w�-A����"O~��PJ��A�؀��`�5l��5��"O�I�ס�.M�� �/��*��v"O��A���2Ą%	����(q��x2"O���^%c���ۋ)o^��"O�qae��k'�s2O\�,`��F"O���Q��V��$EkP5��"O��)d��N*���'�L�wK6� r"O�5����F	��sC�~M����"O@ ��)�� ��seH
F@�3�"O���3G�!���
P�S1Ux0"Ov��g�+D7t�#���0���"O�隡�&mx���7i��(�"O����!��m�d�u�[�W��"ONX(4N�h��y��͍�u��H�"O���5<��kM�!���8""OĹZ��Ӗx%�%�!N��r��%��"O��;�B��d�0X0��^���Q�"O~刷L]9,nt���M�XTѡe"O��s�ς!��]y��m��(y�"Ox���6v/�kgaC>0ځ�F"O�4�
��b�Ȃ	^
�P��"O�)���OG�m�U
O�g�^�9G"O��*F'0L�8�2
�h�X�6"O����R�����cAf��d��"O>������F�a3bH�5�8�g"Ot�a��'��<��ٗu�j�e"OJ|�FB�5;3��rs#Շp��·"Od����KL����{w��+v"O
H���1G\�@E�0Y��hE"O�\�d��tw�0S����5j�"O��R��Μ*�.�Y���z{ة�Q"Oz`@��<p��t`'�$bvM{`"O��W��G�ta4���.�,��"OJ�*Q�J���� ^�G�H�C�"O>e�1�Ii��3���T����"O�IQ˘�--�g��4j#"O��W�¢0 �2��
i�:��R"O��� J(e8b� |X-�p"O��7�]��0�H�~���*�"O������?�.�1e�0���"O�q�#Jސt=���C ;��@��"O���l�%q30!�sdLD���+�"O,�z�$�$]�\`z�ȃ|�n܉�"O�P�i!`RZPu�I�n�nP�U"O�����ЏJp�@���o�Z�Q�"O�r��^�VCP��u�W"|��4"O-�%,�]�J؃�%K�	�:�"OpV��xH`���Lra��jS�@�<�D�f��� F�?�B�z�JR�<�����-�0�v]�=��'�V�<1����u��|�,�E�T��J�<��0h\�c�+P��ŉ�C�<��$�WD	B��ET��w��W�<9Q�!ȼ�U��$gc�Cqg]y�<�h��:]h)�B)$"���#�%�x�<���P����K��P�Bi�<90Ȉ�"kDI�ŢOC��y��B�<��c U̚tqD� �0�M��N�y�<��ANq�����9 (Y\�<9@�ǚ0�6a;�耰T�|�@t#BC�<� ����� &� ���#X�(�"Oڬz��>��U��J<R�NTPp"O�Lس���@B�8� �2g��ճ�"Ov�K���`_|�@U/�e���$"O�0"3ꋹc�4,�Ʈ�(m�t��"Ot+�i���R�q0N��D�"O^1���'LV�j�̙�N�t�0"O�9J�n@8�F(;b�ڑ/|��"OrX*5�Z�v���_���i: "O�8�\~�t�d�NҠH��"O�yq�C�azr�1���2��	��"OL���J�Z��1hd�	E�� x�"O��*�eC�S.�8f�^1��b�"O^eo�8e�f���O�#�C"O q�� cR0�o�,YCE"O��q��U=Fg�y!B�W�]"9��"O~�c�H�Z��(�WMƹq+�Lja"O�=�w�+���`�l�]4�
�"O�g�b2�C�hXU,~H��"O9�5�X� `BaQ< �My�'qf�BT�A�A7��B�Ϋ	�
�'��Z���FѾ����R�Fѹ
�'-� �v�­u]��䎜&y�<��'��bcD�= ��	�y��:�'�`D���A�X����%=���' R\!��454�jq���;��%A
�'q���ʂA-�`��H.(�yR	�'.��$�JX8�Q�g�Y�6>���'=7'Ր)U峑�χ>O�L��'0� W�<�ư[��`H�]x�<�%mA[��؇�Yi�1�w@�i�<I"��1X�M�SB��w�Np�<Q��2o���r,��LE0̱���C�<� 7zQ���ȇ��q��}�<�sRYl �+
.��a��D�y�<&���nL\��pDEC$by�G%�q�<鱉L:��(W怍����0FFf�<��ş �lH�����5��H�<�%$�6���3v*ӭP<-c�JH�<�7���@]�`��,m"�9``	�D�<��\�I6���
ν��a!��}�<ٕ�Њ%�1�O�X��4�D�Bx�<����<�~�:@��VL�'�x�<)%C�    ��     U  �  :   �+  7  �@  �K  |V  a  ]i  ct  �  ��  z�   �  a�  ��  �  )�  j�  ��  �  :�  ��  ��  �  ]�  ��  ��  4�  ~�  ��  ?  ] � =! )( j. �4 �6  Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�� |d��"O
`�(�;���8���-0��1%"Oj4��ND^[��"3/9�0|H�"OB���H��*�ʞRy=a"O�味V�!X��!&F�:J�$���"O,��a
���C�Ą�M�"O,$3%o�-���p���+Ն�:1"O��ݢ1����`���y14]2��i�<�6��{_���c�H�`�fX�$Kn�<��A̼VI�xR[�)�Ć�pඤ�ȓA5��('nߡ4�� �)˩%� ���,��r�؊b#`T�eT09���ȓ!�b��g��}�8�F��-? �ȓ
K|m�ș�VṔ���2�%�ȓ"R�X�j�4JN�1�˘X�i����̹	_�jZ��1!g��zܶ��ȓgil,*�J�
j�Ne��i�J%b���f	�(U��:���G��$Y^م�~r�� S�%T"���k\�jx�ȓ|4�1�îJb��@ӵ�ݩn�V��/[`�"�v4�R�!ʎ<��M�ȓ`:��z�ؚh�J�Z��$HY:	��H��p�m�C1��!��B:��0��EnjZA V;9����J[
2���	��4'J�EA�IVW&��~�(aZ��ӹ�>� o�Y�|�ȓ�f�A�
Ο7�H��M�$�����mޠP����/���ANXo*�ȓTv�����{ ��-7�*h��I��sB�8�8���3����ȓNe*M�悡;������X�o��!�ȓ'lj�#F�m�+R&;�|��2)n�C��0S4���T:
b���:�0!��e֊��)��ͷV��,�ȓ0�&�8#���� ع�L�����;�P�AFd���,w�6d��r�EQ�( �gVlɦ�M,H��,DP���|�I	$G#\���ȓ"�)���E�B	yt&B�^�LɅ��wyr*\(u�@ UV$ED02�-Ə�M���sӀŃ��L%'�r|�f��52���5"O���BO�876A�%x�`J&"O��@��~�nW�8\0H�teE�<A/�6r^�=��OA1 D�k#AX�<�A6I�P�j��B�0�SJ]�<�t"�>{D$1�dȫK���b���bh<����d�n4�s�C6P�NT�T�E��y"�')��m�):T$X��䔗:,.mi��${��E��$�@�Xe��_�F�:#�_�yB"�	s�9�1䗿E����A���y�	Ǌ"�
!�حNn:tbqa��yr��ZCpܪ��Csld���W���=!�yb%�.��m����=1���*��yb�խD?fd	$HZ���h�E�a�\QEy��9O6y�D� CqX8!��A=	z�!#"O4l���	�/��]����n��DI�"O@��B^XX��V�m(=h��$�yҹi)�c���SJ�ODIi���.h�xsQ��E��B��~B�@���!���D4a��������(�xźgȒ�i�2I��cD,cĸiQ"Oиc`�A�*HV!���A7VԌ	��|��'K��*ͦ���"����� �m��	�վ��1EʓH�̒Q:O���d�w��� �D��(4z1ڴM��IZ8��$��Q&�,��P�$F-@�h(��j,D��Q�nE 7���F!Q�	�Z<���<�'/�{r� "�li4��*:��$�����p<aM<灵��Y2��
�d ըP[KF� �hO�S4U���a���?��;���P�C�;��$�RI�&"i�<�g��E��C�I!f���"��5I�d�ɋ `���hOQ>��I�}L�� Q���ը�O�B�I�E��+��I3|�b�nJ�1�P����p?����<8j�y�Hύp���Ɏg�<Q��KX�� 4/�$H��-�4.�a�<9��\�\�� S	�
t���`�Z�<qg��Z�����-<�@��Sܓ��=��$�FHUPơ�'Fa4-r��N��4oZ~)�f�΀.ל�rመ�wt��Ө����>��OH��<��L��Z<Pv�@���i���	
�a�m ���0	�xⶃaA!�dV=�=zv�ܼ(\a`�ۄ
,�	��HOQ>�PQ@Ъ��83Ff���*��$�IQ���'DŚagjP�a��:5���e��-�ȓC9�=a��ˈ.~��j�/��l�& ��Q9�-���
���Ĕ�T�l�ȓb�zT U�R�h�>X��O!\P��@���@����t��l`)ϨV߼����6�H�'t�i�#L�(���I�4C�^��.��S�O6�=a���6�`������?O��=���OyBK
/���@��$��t���O�x�3�'��v�i��x���<&æ�B�O'<����en�����؟��.�S��mܲ1�Y��悽9&�H#@��,+���Л#Ы�,֛F��"7�J;�!�آ@Ӕa�q��@L�K��P�!�d�Ȁ�[p�[�X�4����B��I��0?Q���rA�u�u`K�L��ܣ�m�h����'
j �S��}
 ���ć<sʞQH�'{�m��ꁨ%�v@i�m�Z,b��$ғ��)�O���?Bl	�p4�)x��2M1�tєǙmy��')����h0aCx����4.���Ì�dؖ�?����'�)!��T�n���N4(�2�럴�'S�OTi�礂�p,&0�	��	4����'����'�t�`����{�O7|~��;�O,�=E�T�I5O�r�2�H�r\�Pր26X�'���0,Or��e�_�<�����M�6���O��Ig�Ӻs���2��q �%�m��� 4�D&"9 -��P��\y�郂]�$:iY&1M���	f�T�d�����+�X�i�G�k)xyD}���)1���0�6{ؤ���(B��4%n0mS`��y�*��+"�D{J?�YU�Q M��yB.�a�*,��?D��`�2��ti�n� f�T�cq�>�y��O�f�ehG�~�q���=x���z��6-Bg��r�eܲ�r��E���r�ў���ɂ9,����0Bl�{uf8$��=�N<����8}���i��$M��٥���y" ��nD.���/��@��u��Ѧ��<��o�>+OV9��O�"�(���Aļ �v]��"O�̱6
H�W��)Q� �<9i�4Se"Ozl�1L"e�0�ڀKVj=`�'��d��d'8�!�3�!9�c@�(�}♟\��� 'pn���M�)'�<��W�/ړ��'���rB��b�F�ج
r'+,I��'�a}g��1�ŏ��(�&Ya�K;�?щ�4�8��'?��j'ҸP�ƻ�f4�Q�� iX�#=��S�? �PХEׅK�|�A��ԊQnm�Л|��)�ӨZ`>���ܽ|��U��_�C�I2�F1�$�ʤR��%�s/6�<u1
�'&�Ј���#�>d��g� _�D����O����S�Q��)e�9x�h���"O@�ц�Y��b�
�.�0u*��'UV��R�#���L�6L@��n5��"$D�`ZB+��N<Uk�)�VYc�<�ٴ�p>ѷn�@684��]c뒡���$��d9b�Q+Z ذ����,u���/i����򄏄���-�'�x,�KӈF��\�c��bӬ��	���:�:�	Y|�XP�n���Ę⁅(XN���'0	�!� X�H9C��.5��=�I��F{r�x̓!��-Z��Q ���DJ�X�̉�ȓk������$0�.	2�ŏ���u�'oB�i�1O��g�ɫi�,�7�E�E����&�������O��	T�� ����G)VR��碇;�M��'>�E�tK�1_�̹��W"
��F
��<��4ø'�V��AFH9�F�	�CsD�@r�y��'�X�
��6|M~���`N�c�T����4�S��m�=�,�qrڣ:F��uÕ�y�I�'�	iZ�������eKI��D{��$��9��DU*M�g�Y��*���yr�� 2�x�&���6��s� ���f��a��_��3�h��5kL�ȓ RdA���(��HAqB�֘��ȓT|�[ !��#�xiuݏ"J!�ȓWٸѰ ��X�����1����'�~}˕�%zeI����)�͇�=���� N �����pt�9�ȓrV2�`!͵M^6��ckݦƶ��ȓ��Jd�=oA�В��RU���'kP SMȸrւ���S�F�����>���-	�H�K�r��ąȓ�@h	�ŊC6�xSՇ�/�佅�*���*W����)��F���ȓt�ta���P�d�t�iŪ�\zH���{ FH	Q7�8yr�҇@�����XqF��<A���б����8�ȓ}T��e��
 *�����	LpdՅȓȈh���I'����L�=?�����*"�%��=.I*��?��9	�
�<��Lö���y }��w�L��1��8,�Yb�� e@U��9�@X�䚫Y��9Z�hO�i�j���*m�!�1�ͯp����W��F܈�ȓ_�\���ݤba��H���3r���n�X��6Jڽ�� 
�L0����5�hG�L}s������i\�Q�ȓ$zD���'�7ae�L�b��S��e�ȓ.�	��c��d�x� )���i��_c�*� �=���E�ŗf܄�4Ԕ����[�(��2��%nT=�ȓ���P����x_�!�	Mr��ȓ,�uc4�]�#֌��E�Ȟ+���ȓ92�I[�D�X�i��%t��L��K)n5
�)T(|SJ�r�J� n�rͅ�k3t��&և!�l�J�E�vi��ȓ)�~1��?Sq<�Z0�֘~7�p��;�}�Vi�<TW�6�LXo^��ȓ:̽1�Aϋe%�aQ��y`�ȓB)���g�<G`� eͼe����3�xtS�	�5Vd�]Ф��-�"q�����p����0����)�+|�$d��S�? �Mqg�;7�r����K8%����4"O��%&4�0����h����"OXLjgk :"��sJ��Z�v�a�"OD,��'S�#ԴT�Čc�Ό��"OLٹw!�r��� LVoӒ�:��'5�X�X��������I������&��;Ej>��E�Cx���	���	�������X����h�Iן���4<h.v2����,i���5@S�����͟��IΟ`�I�����������$J�ٱec4� dC�%q���ɟL���l�	��������	���I̟\�Ǡ�kC(t���A&���X�u������ğ���� �	՟\��ܟh���L���2�/�%��*��V &�2����0����x��ʟ��Iß��I��X�	,�x(�Vd ����ZZJh�I����	�����ڟ���ڟ8������ɶG�њ��_9{C�@� ��F~�u���`��@��˟���ß��	ß��	c���z@���.�	���I,>YBP��˟���՟��Iş��I�(��˟|�I)46��"�	t�Q��!	�B���ԟl�IƟ��I՟D��ş��ß��	*r��|j�O��8�D����H��͟��	˟����ҟ��Iɟ���RN���!&Ϟ,4\$��KLr���ʟ�	��d�I������ҟt�I/c���*Ԃ�4^ͻ�H�D�8�	ڟ��	�@�I����0�ڴ�?y�Uf�ܚ�?n���Q�ӗ'���wV���	ay���O�Ll��#�'�o���0C��q��=I�E1?�R�i��|��~��i�8 ��̅�l}�/��0���cӲ��Xb��5r$��sa
Y��kԛ~r$KX3�)$���vl�y�`�k��?q)O΢}b�gĿ:|P����0U]�uAEb��,>�VA���'m񟮝nzީHg-�"��9��OU0{���0ҁ�
�?!ڴ�yB_���I�b����F�:h0Ő0�0Z�<2��Ƽ��dPa4P�����z8j�=ͧ�?�G�	ce�)3Ѡ�� )
F�<9.O�O�l����c�p
 L9��0
��Z;:i�eBg��2���ܟtl��<��O:��F&ֱc��a���1"1�ŕ��S�#��0��b�(!�Ӕ3�PB�+ǟH;5͉�[��(㄄?b�{���ty�\���)��<����dR(���DM ,&�۶ ��<�W�i�H��ON�lZ��|R�a�F�f�0�eɹi�`h�z?����M3��h�p�a�H~�#�`F���*;�%��ѡi�)p懆�]�V�&�i>�'�O���ie	24R�q�� �<��O��n��rb�L�SG��/^��Sn��
"}�̓10U���<���M��'߉O}���'�4y0�� %:;���c��G�8�p�Ow
�
�O�=����i�,��R�hO�����$r��*��؈@Vyb�A�O����d!�$٦m�DOc�h���
�����"�ę��G���4�?IL>�g?���M{��#E\|C�f~�p1�� 1#ڑ;�K�=�<d̓� ���8	AP(2��?���ں+w�h�e��i�U����'��AD���c{�4��HyrS�"~2�#΢d�<��F��J���ŭ�|̓ �ƈ[��D��$�w/�1 Ϩ�˷�F;~�(�'�Q�<(O�7m��������H��l�胧��7q'��ԥOcn(pǣz����\��#amޤMPn,$�����U�����G�����
����C��&���	M�ɂ�M��(�]̓��	\|?��8�i�-nOj���J A��	���O6�x��$>�� �1�*�0�u��]�
�d	�ۭ7� #B2?�'qi$t�A&�$��x	�y��)6�A�����_�2(�/O���<�|�'Ĝ6��,��2�'�LzIr�&2�X�����;޴�����'1�v�e�&a4�I��}zJ��q�.6��O���׿O����O�M��� ��c��� #5H�xT���b�%\b�0V�|�(�'ZR�'���'��Q��S;�����
��,�+����-~��ٴ>�H͓�?������<I���yǆۖZ�x����8����4@æ��7���!����4����������MJ��YV~�&��L�.UXUi](eh�DҀ9���qElR�L� �=	���?��Ο/lE�)��@�
P�Qf���<�.O*�O�	l��<b�<�fF�,!S< �`eB�J��`s��ß�&��j,O���b���c}Ri�cǔI���P����S*���y��'���:%�K�p��O|���_�x��O��*�mW-�6��"ج}X��R��<�,O���s�tԮ�
x���dOB�b�+@�VI����1���"?�iҘ|��m��EJ.l�6`�רՔ}�����'Q��Jcӆ���?dz�>O��dP�A��!Y��I&�~i���%�:���n�@�H��7�D�<�'�?���?����?���TQ`t�]3�xs���7|˓G�v>u�7��OJ�$�����G2Ob���41� ���J�*0�v]�ƠŰl�D�'":7mCȦ� �S�S�?����#��5�C���$Od)CC,؅����s�%>�b��':�؇JJ�t��P�1�|�Z�<#Vo�"W�h�FCռ+�`�ʍ��<��ԟ���۟��qy�bӾ��6O يa��W#1㍷�PP�U��O�ylZc�i>I�O��o"�M�T�i�D��̈́�u>���7�EE-���w%�#,D��'��dK#naH�;�M�uT�I�?�2X� �]y@"� B6��!��^��:B;O*�$�O����Oh���O�c>������
�v�B�?��8���,y�^Y�'",m�z��w:O�d�ͦ'����m�:$p�Gɯ
m�*�7�M[�]�|�4;��OUN��E՟�yB�'�:���W#7�|Y���/e�m��ԛC"8�ڱnI�U2ў��	Yy2�'�A.�;�*X-�Xr���y2�|"Nx�||Cg�����I
�M<�B��-S���cF�2.o�	��D�Oj7s��&>9���W��!Z(H�f=�T�V5�\z%�A�����<?a�'#:�D)�9��X�5�ߓ<j��8��ɫ^65�(O��Ĵ<�|�',p6�շ7�^-��@Y�-����霑1�8}����4�?�L>�g?�޴5� �eJ��zD�[������A�i��A�x/>q�'�˔�$N������;��$GjjR���:��I
Ԁ�	1O����<A����%i�Tp+0��G�jC�%P0Do�n}�c����J�S��M�;<�R)�fgT3sU��  �GQ (���'w�6?O���?��S�
���!���,d���9$(37H�$�؋"o�牙CR|eB�D�0Bь�D{�O����S��񐥈��8��vc�)�y�]��'���4]t� �<�@J\5 �� �G��4�m���?	J>��U�@�Iئm�����'"ءD	Xh�Y��֤3?��O�� ��	K�(M�������jA�tFMߟ�g�[K��B�� wv�h��͟|�Iݟ��؟��|��h>��?����N����"��:/P<���/䛆kI�y��'s�6m+�4��Ή�!e09z"��<L�Tvj/������4
֛��];p����'-R��DN�I��_�2�\�(e�\ 
{,ͪD V�>r�񡖝|RP�`�	۟���ӟ����pd�9/�Xd!�K���8� �XQy�fhӒ9�7O���O�����d��'�h)S��:^���r�߻Y����'�7�_Ӧ�c����'���'S���W��!:M�|�UE7^�><�� Y��I�(O"m�&F��l�+&�.�'� �0gA�q�v���퍓\*�x����ħ<qJ>Y��i=��[�'e�0�5��ΆM�� yb�U�3O�m���$�泟D�	�����_{l����t!�ˋ?'����½ J���~�����1",��g�OJ���л�0y)���
��C%Z�B���:O����O.���O��$�O��?�A�ݤG��˄m<��ۅ%q�\�Iݟ���4T�V�'�6�$��Ơ���6O�JA���tn�)�Z nZ���ӧsY�� d�OqZ- &�[%�y2�'�(K��%�r�A���J����a@��?���� dVў\��gy�'���I�Q�Z҈4�H��Z(ɚ'��'#�6-���1O.�'u�l��s�ѵ7����MF�.�'�ʓ�?�4�y��d�OP�u0�˨j����`y=I�WDF|�
�q��:>Ĕ��r��8vx�)H>��� 4�B��媅�i� �����?�?���?����?�|�,Oڸn�:e���	�X�<�c��{������<?���i��O�1�'�\6��<X��6�?v��E��12ք�l���M�&gܐdF���?�w N�.x���B&���fi�Ѣ\	r:���˅3��D�<����?���?	��?�(����ņ��D@���֐1�8�ڦ9z�`u����ß(&?��I��Mϻ)ʹA�P4g�b�k��X�=�<�7�i��6��,ק�t�O��t4<(�y��'��LWi��jLfxH������a�'���(
nv�k�|X���	����dhF��e��(G�#�3k����I�t��ryBOퟰ��'�r�'(F��$nn�|;Q`�r������c}�`Ӝm�?a�Oĩ
WK��T)p�b�Ҫz��&<O��D?q��ڷ�K�w�˓��4���-��]2���Đ�� n����҇.�X9���?���?����h�d���B��(��I�j���WO�Qnd��MӦ�k��b���ɂ�MKK>�缫�@[z����bN��l���#��<���i��7���ICeJ��H�	��$�ei���~Dz�.2.a�p��Ɋ/s*P�&g�npƌ&�T�'�r�'`��'t��'; Y*�ț(*�|���oN�+"W��X�458�pR�ip2�'���#�y��'flȺ���^��v�<v��⃦>�U�i�07����$>����?��کH~�I�E�S�z��oU{\x��G�FyR���5٣aupўĉ��0jڊ��q�.hGB@�s�ܟ�'��I\�	��M!��<�IƁd��� wᄨky`X��	�<���i�b�|��~��'���'�	Q�J���b؈'��wk0-yG)�-^�	�'���&tA����P���d�(p��Z>�P˦C�
n�24�%�t|���?�.O��S�O6�y3DS�k��`��,*~�y"or�6��Ɠ��
ܴ�?�(O:��4�S�E����p'\\��a�̖'^���z�R���x��3O\�� '�n���;�*���H]�E�u�1A9M�FY(R�"��|Z/O��	�cK�X+CŊVo���� Dk���(���ǦM"��)�	H����2�Py�f/;Rhщ@�����Dy��'���=O$�`��AO�Q�0���`54�G`��!���Ͷ+ �ّ��d���Q,R���$�Z�����R�hB�D��L�!�ϥ���J�i� u#���%�&\�џ\�"K&ڭ�6�]�nqjS�Kxz����R-{�B��僇L�>[E$��"�De��;J(�l��_P*�Ia�Y;W��qQ`㎝x����#�Y�? 
U���q�=�b�_lC�Dڱ*W?)H��vո8�`��L��Z�IP$�N��E*a��]':��2ڀL�ͪו>�����j��&��3,T�&��'4��']�'5��'m�D����88��1��R=08�Rm����'\2�'���'?��'�����{Ӷq�'�>h�D�u�(aŲ�����t}�'>��|�'?B!Ι}q2 ~H���E�`����7,PY��7M�O��d�O��d�O���_�|���|z���'6!k%j�69�nQ3�Z���Ig������I&=,m�	���	�O�l�y��V�YX�,�VV(h�޴�?y��?�j�@�Ĕ��'8���I�U���"�</�dt�B�W�/$RO����O:0�j�O~���O��O�����)HGǐ��b��h~(W0f�s�	8U�>��qDP81�:�v@�0a�P��{l��k�;z+lPC���R0f�H��Ѿ/�y�i�'w�C�	 !���5#GH݂�yQ�^&;J,r"K	�T"V��������"�'1�̐�d���9Т[,:̲�H�-d��z�ȅ�R���u�H�:c�za��a�H�U�H�S˶x���>��'͎�F��h��&t�P��bq�����2?P�1� -�j8ДhE�?���j���3����˟����H�_w-2�'&H����ͲW�`��(�|��4�g��2c���ꖉ�p��S��Ƙ����I�d�P8��m��9T����E�qX�R�IK?s��%�s%�6j.�g�?�������'c}2���,��O�/���҃�~I.�?)%�iN6m7�I���	XG$�Pq��a
�!�.T�G�!��Ob-b�KX&F^	���=+��)y��	]�'�T7m�O�˓c6��{��i˸��K�Abz@c\K�<t��'���' ��8�2�'�}�1��JW�u���gB]��h�Q=d��;H� �@���ci�"?Y�� =!���C}}^5��L�*���rV��b�F����(J���,W�S��%LY���P���럨�A�֐wR�QoU�d��X��*D������#�H#S����I��)Ọ=��̍�g��L	D-�,Tܩ�׫��<�!�i��'����bj��d�O��'�։++V�Y�b�,��j6\��a��?���?)&��8p�;t-�*7��S�T�³AO��^$ V��� P4�(O��B�ϳQ �u���|�'v���&�Yw@�3D��M/UDy�bQ��?����'�?)��H"�D��U�'��(pI�>�?����9O^-	+��-�
�8��E�rv�)0�'ҤO4k�ʙw���7k�9XkZ��=O"	�G����E����̔O��1��'�b�'r���B�4%�r�i��0t���2bA���/5�m�G�t�v�T>��|�	�*�L��л��6��~�쐐�H�-�H���N
Q>t٤H Ɯl١.\ '����Ͽk��]@"��oQh� �-��&������ɧ��r&�-j�ޝ8�IF�}��1
A)�y��]<?td(_I�
|�Dķ\"<a�)�Q�X!x�E���D�`�lu�ի�?�?����L�&	�?���?)��o��n�O��+6&�0ud�:��5��Շi�
��44�V�҃Cҡ<)8p�!ɼ?�=&�-TV����3"z"Ѓ/W�d6m�f�PIU�A>2p�s��hO��b�ЂyÀ���]� TY�O�F�'iX���͒���(�aV)E�$ہ��)�!�84I�E�k�,�Ly�M��:C�|Dz��� XGL�oZ=��<isԞW�T₦=>p���۟��I� h��������|�p  ۟��ɺn�n�Ӡ(�(Pi��xrd�;�.���O��I=8;�%
Ù�Z��]KSH޲*����M y��Nn�N�� "
8Z�Jp)�/��/�y� "O���%�\T�x�Pd�ņ[ϼ\CT"OlmpJ�w�`E2�O27&l��b1Oz��>I�hϢQv���'e�Y>�P&��5Th���� �*`qG@�͂U�	����	�ܴ�.Q9h$q�J��?�O����^���B0�Ȼ1d\tY��$��3�A���*��s3A�!D��P�/Uv�T���@�Q
 �Q �#����'����G�td�:n��Xs�1t�L�鰦F9�y"��;�����hL&q�h����0>r�x���$0���m����V�y" �?E�.6�OP���|�����?����?I��S�fж ��	9l�i:t%��\�eI��8� i9 ��.e6~=�b�?y�|�݋' $�{2"�`��22+�<b$�@�<ar��jF��V�B��MqDҢ'K�����B����w:�=��E�q7$}�W�o��0�CۂLY�d2���O\�S���;V ����H3D+��D"O�S��ϥB�dP����y�&��	��HO��O����1�6�B���u��0)S��OL�n^٠�N�O��O�d����Ӽ��A<CL8x�����;�0pN���`�<j�PH����%����g�'���#m�CR���ޗ0 �q�ׂ�TPG��h��50����D�i6eҟ���Ϛ3$*����۴�|���:-���M�>���'戁ȥ�@�){q�sJ> Sف�'�X��5� Z@��Qā�#b�jE�f`*��|J>iĪֳs��� ֥�©J�8��I�b��p�J�O~�D�O���R�?�����OD�1U��U���i�<QP�	+Q,\�c�]1_�k�h�F�P$䈂��OE�4��p����6�OK
,!��#�h����Ř�.0ط$�
H�\\0�F =�\�b�,�dF!=�lӰ������< X`�S�Z��D0�"O�E��͔������J2Hڈ����'�ў��Lۻ6���'��~ݎy�� a�@��4��"Z�s0�i|�'�哛FT�ɲ�ı:�p���;GW�I"�
^�4�	��K������<�O� Ȉe�V+0���g A�~�hLÎ�d/Z��?�"��
�f�0�ƐN&�@c?ʓ7������H���
�D�%sh��e�+!���"O؜2��=ظ$�`n�����'�XOx�k#X������:"�����=O� ��	R����͟ �Orz��V�'z��'TV���	�u�6�� N�Q�[A��}���E�^o"�QV��O�Sl�矀��ß0�\��t���b-|T$�b��0mB�d0`Jݨ�8a���?��X�W�/��;wM��hf/K>es��LQ0ls��ʌ�?Y��|���'{�E�(�0l�rt{�D�rZ����'GҤ�R���2�"�s�>��� X���d�'غH�Ę%o�x��m�gI��v�'x���e?�PZ��'���'J2Lt��iޝ#%ǳU`��jT,.<�11R�������/�O�|��O$T��E ֊K�X0���O�C��'#Z" �]��E�aD�=41���'�P��1�a{rJ�  ��Րs��Pʩ�@���y�NW:�j�!��]�<)��0���m�"=ͧ��Tr����i�&��呠8 �
ӡ�-hJ���F�'r�'b5l���''�I6^���'\9�f�Q 
<t�j��T*O�U��p��M�'�j�;צR=5f9rBԐC�T9�RG}�	��M��ʏ�0��F�	��4[u*W�<#���VX���Y�&h]�B��Q�<� ��b�ҴKp ˈHl~��!��<�A�i�'T&!)P�b����O4�'
�0@�l�SΌ�P���hFi0�T��?i��?Ƅ��?�y*�PW�$Hw^�q�P�� �Z�'J|`��)���a#G�;͠L�F[.dQ���@��O�eE��T����T�ҏ2�6�Cb�[��y��h?dT+p�B#�}�H��0>�g�x2�3�P�9�@B�u@��2 ��y2���&6��O@�d�|2vD��?a���?u�{�K����|��@X����G��tFO�b��8�h�/O�(����4� �1��
����&ĊZ����R�GO:"Y�@�H�sD(Fq�x���'� 7�
ky����Ү�Vh��i	��3	nJ����y2�'��}��xX4�qBOG-��-����O@�Dz��O�L� )ZI�ۮmZJ��̛�/���'�´����Y�"�'b�'DH��<�ɶ"��	�뒰u,�=��O5y�p��x��j��R�z�d�
$��v�'7h��b\Yh��� J9�A�5O`���C�9w0L��U-7џqK��0o����Q�Q%2���џ��f����ش�?I��?q���?)�Ӽ{�C?U����I�|�$��
U�<qa��nt�p7�ϴT h̐v'��8��4�?�+O���EZĦA�)���:�:�)X4�
p�f�@ԟ��	����	9h��͟ Χ����֟�3��;8d��3��}В Q��1�Ox�*�R�LK��ip��B /7��Hء�0�OJ�b�'?2 [���������R.��{����ya��.T��25�x�R�-���yr����j���#y�q��+#�y��n���OxP�Ċݦ����T�Oؠxa#�����E,ʕ0��5=��'8�A�u�J�R0��Xt�e�,6v-1T�."$��paB��K�as�����@�Hq��!�L��Iu^<��-x����P���
G`�9B�R�q����'|B�0ҧ@H��#peG�rᐔ��/�Q�̄�$K,-�U�_�kN��b����,d��ɪ��}9���g&�1:48@1-�� ֞����SS�i,��'���~㪴��ҟh�	�.�h,��D�#P,,m��.kI��`�+'ą3� �����5�Ǫ��a��c���h�A�c��rt�ēm?fi;gO�Uv�:ƨM7tW��5e"A�.�Atg )W�F�zW�*��;���"�C�!BN���mV?w��q�h�/�?�6�|���'���oӐG�!�N{���'m�HrDm�rЁQ��qQ:���ĕX�����'>(�3V�r�u��IT�\���'&���%� �k��'4R�'*"i��i�� �HƯ����tpc̙���q4�O�!g�'� ��Ȋ�.���i��^�S��]�%,�ܦE�X!
��\����9�r���a�N�,�A&�)�	���N؞x�*ۖ@�0��2�$_X�b��-���I]�4-[6Ȁ�p�ȉ���3
+��4���O4t����a[W�h���p�왼g�i#k�����	ܟ����kM�i��ڟ@�';VI����+G�y�"��'�F4�"3&=��
^,b0�p1LH���OJ����LŒ� �g�P2�"W:P��h���ΡVo�lqW%��C)�7��Q���$ÆU	r�m�$!���.\\���ꚵ��}c���Ҧ1�ITy��'q�O��L�v�k�'�/v�"���S5-�LC�I�T_�P`G�CiR� 3#C�p�扼	>p�IQyR�_
�$֝ş���Z�T�A�y����v,�=b�X8�O�i�9���'���'���
Ӏ(k�R]B�j� Y����v���Z���h_&}�8��4���%��� ��(O~��n�=m�� f�б6@z�zr�R�$٣$
�z�p�(���W֐�`aaUx� ��*��Ux���*�'1U0pR� ��)�h�� L��-�ȓ���A�"[I�`�ѠA;l{\p�'�ў�0�ē��xcT.��T�V�Q�Ȑ���Yϓ(_�����i��'�S�#����Ο��4��)b%[�d����N"cܹy�M�;V>�-{bI�K������4���^qp���/\,���m�.yT��'�ՖpǢ���'O�O�����L0K�^���#��#�Yk��w�&��e��z\F�v�Y�9z��P�R\�B4���O���C��4s�P�����6"Od01���*�yzI�&�2�	;�HO�i�OB���&E�Xѷh�!� ���OZ����	�"@��/�OV���O���]���Ӽ3e�!F.b����	6� �Eǖ{�t�kW�� -oF��G�n�	���HO4
��K�Nd&�ȠlY�s�a@Ю��	x���@���!9c3���a��訣�Ԏ	'4��'r�ȧ�"CGlH�F�"�����cdh�O���I!k���'mG��M{���3BC��PłQ����!�`)��`Ǽjdq���4�*�O,$3f�O�ш�C!,2H�*D"�-��b��N͟4��������B������xΧ.���(�M
�k�$(�(�d��Ga
	��!�%�Gn�d��ʈLzfp��(3��� 2#܀tNx��R��;30 �2�Ň "�F�Ԍ/@r(B���D�X�AӄX��q�I>y��џ$��4G� 9 ���`�K�{z�U�ȓM�yw%�2�P�eoÐC~�����y�'�6�B�ٯ@8�<XpK�4m�*ܘ�'[`6-'����WK��l�̟��	t��� �2%[���8|4m#vD�)} 6�#�'�B�'Wj%�D�'�1O��1�� s�A�6+�YӤ�Ժ�~�<�j�h�O��`KA�c��bA.�:����D
���S�^��9���1@�8�W@ĔS�:B�I�eMX��AC�S6b��!�C:0Tt��$�q�ɯ4���y%3-/0��遈do~�	�;�I�ڴ�?�����	�$hl��O���gp|�R'��Y���j�
��A�,C����Te��9�����S�d��w��1a.m����v��-�:���gD%��q�'M2G�e�J��f�}�]�c����b�Ŧ@�Q����8�pU��ߟ�RH>E��k຤�c�b��JI�&%��2��L��oo�}�Q.�bhT8Fx��2��|*�~�,-�҆�"{� f�@-K�&�x��?9�g������?����?�v��8�4���3�T8>8x�yQ���?��4����NQ�@K� %d �R�!v��4ғU�|�x'��*b|��p`ۘkΖ3g	
�wwV��@��
�Y%�y*�4P|Tu	_I~bk��2�[�J��l(8���%�~R�ݒ�?yG�'�\��U��`	���fSo����'�j��A��Nޜٗ�ȩ%�	2�E)��|�K>� !��]���ǜ�tx��J�{v.(��QMzb�'�b�'�x��'��?�������_�L�.�x��p�m$Ob����6�
�FlP�'�¢?�7�S
P���Œ&�ֽ��	���
d �+�).kf�3�k�Z�X�۴5�pI��#P�h��]����M{�hٶl"=sqdD=_��ex@b]K�<�Bo�����;�6-��M�&-D�<	���$��#�C5gd�����<�F�i}�'-v�x��l�����O��'7=�7�U�^�"a����DFH�D�?���?�`	{�`����C�T>9V
KZ]��/^�]��[b�"����	�L^[S����/w	P�T����i�V�v���(�;�*�3���(O�Qy��'t#}�f(]�@u;���2���Ѡ	S@�<1�&�%_�<D�	�C����'V��I<As�ԸT��u�5�D�iU"��<)El�Q2�6�'�RR>����̟��	���S�3�����h��M���a��)F�9��ʶ����g͉v�Q9��hc>�� �)��"U�Dv�� +AJ�j5�\�KC�U:g�ڤ<G:��]�a�᭻m��yFi�\��w�l�* !ǚB���0-�8%�/��"':���O� i��:{.����q� �*�"O�	xG�M��"4I�� ,Aa��;�HO��OX����JU���� ��<>���T��O2�D��as��1���OL���O�������Ӽ�%D;S��u;��]�D�g�y#52��T�����H@�{���'�HO���%�+����/-4j�BBI�0z<�h*�g�&.LV�B X2��	}�R����6=r�I<h��E��]+82�
"�
�e��I.
�R�P؞\�e(\�,�����ɊBh��y��Q�,���S3��	<�F�V�ʏtV�"=�'��:~���i�^x��ɑ�m��1
f�<cIT���'�b�'FRK�*}���'��	M'Uфӆ/��I�ԉ��}�\q���Z��Ȑ#>\P�t�;��=h�����;p�t�[!��:��D��:Ix��Ґ��#^z�҆��M�ϩo{�=1�����p1ڴQtx�ஔ/�\��s͓�C��=�ȓ�5�`/�4����FAX�&��ȓm�<����'P��i��Q;I�(�͓g���|Rf�&�~7m�O����|:7o�)Y��u��?d�fo�:�����?i�b����CU%?��^u�@x�F�a���:�r@���5@yt�Gc��(O�dq�P*���p�i�.P4�̃D#l����� �sf�E��/�� %̄"g�G�&1D�6�����m�O�T,����Z��J��L!.�mQ�'t� G��*=���C�A�0Ů}���'LP0���L�L:�e	wӀ�P�'�摃��tӢ�$�O�'o�����?a�2���{7"��&ָ�����j�.Fq�%��[�#7:���}����åJ6M�I�֣�	��مǕ3r��TG[/Y��m�ɈXw��mHd������i����sr�җ�^=�L�iZ'I8T���h�)�� ;�.Z�� v��&�Dc��3D�|����$Z�4m��F��G#<qV�i>y�����u1s&��w�V�:%�
�f�����ğ8�V �7��4�	ݟ���ן�2]w�w_1SBڠmI�'���U9���$����ʱK���o�Ij��Ҕ��t�	��ty��Qf�CRM�p�ne�j{)�nKR�=9t'\#s���s�R�@b��z��6pa�c��A[2�0�@�M}��ɂ�����Y؞d��Q�	�4U�a� (�D+D�����[<j5 pG!x-������HO�),���z;��nZ"0���F�Ē�p����(K�!�	ҟ�����|��.����I�|��c��/�ҵsaB2��P`f��C��x��+p��bb,H�fTX����	�86�T�;�JϨX#ReB���f��Ϛ��ۮHn��K��p�(����-h8qO�܁��'�(6���"�*��g�o(����oϟ%!��H�1���gF�w6n��1�!!�Ud��  �k&{E�T�l�Y��$� @���4�M[���?�/����F�8ifHaBJ�rk�I� ��*!��$�OT��[�9�ШB�S!/�� A�E
���O�`���"B�;�2��O��DԸ�򤌖M�`m��N�����k�(����au�D����&5��|�a�J�2�{ѭ\�
�z㞠�V.�OL�E��*�cc��C�Ն8�V�j�Ú�y�&��[�����"Ե-ܩK��S��0>��x"D�S/6C���<|�;3١�y�f��\�7��O0�į|
p�A��?I��?)G��:���0H�L �	��!��z�� �:<�"��F�֙{x ��c�?q�|���"l^�Q��"G5�-�㝸���0`e�İKe��#	V����"^$Pm�~A:�*(��MϮ��I���Q�?�8�@�������'��O?�����lx�A�9\6u"���2!��)1�`��4�Cx�I�Dǭ�1Oh��R�����'ު�'����}��(S�-Ą g�'lrO_��d5��'�"�'�	�~�;pY��`�/�@�AQ+��=Bt�*t㐳5��<3�G�uH`B�w"��lR.b��w��IK�E{���S��4ȗK�FF���E�Q�S�.9��J��N�x�4�J9�����9��փ�:����.�$BT���ڼ`=:��ݦe��t�'�R^��j@��$�5D��n8	@+(D������u���R�j*@�B���$�HO��)�O��q<�=�c�i[:��gm����A��*0�����'���'.�KQ��'���H1+����c�W��A����N�T��aN���>����S�H����ڊ򄘵�>�7/_+`�I ��H���� 
�0"���V��Iմ� �n�4Բ�R���*���p��A�G�<.Z�qy� ��&���:�"O�hc `ٟ"�e����j7a�&"O�� ��@�
q
�@�K�!�d3O�	ma�	`��4�?����)�Z��+��84F����bQ���O��d�O|S�&]��4*���&=QbX��@�Uf�(q�V��-��9}��1v&�4<�Q�T��LZ�;�ڵ�B'8\��!�-ÄASc� "��@�F!�4(��+@`�i�P�I��*��@K�O��qqVjG~����l�8-�}��'�[���%�ha��)�Y�伹	�3.�'��ء�H$JG
�*��JM�%��'/v�0��`����O*˧]̤ Y���?�� ���(4e�0� £>�j�p��� 20���$|��jA�س:l�SZ����B���-�N�d��Y�с���G�f@�2�o`^%"��o��E#���w����	L�@뷤c�B��w�N�L�B�*���O�Ӧ�/1�Z� �o_+C^�/�y�G\0������)E��7���O��Gz�Oz���=C��B%."?�tͲ����e�2�'M�D��C�y�"�'���'�vם���	���qc��4TB���(J.D=R51�i)r����D�E��XƮ�qF{��R!�2�򂮉�dP�ʂ�ؤ9��P1�_�.�FH# ������Oސ�`���R���} �F�2oе($�,4�04��'��}��O�r�l��JW�5s�g�~�<�Wh�A=�l��b8�D1�똷z���`�I�O|l�#ܴ,,`��'H�C���H�)�g������?���?K�?���?A��@�b�D]���ΚaB�u�1d_�_�<���''�V��w�X$���?��#ҹ9���5(�v��F�!�$(��
�2ݢ�"��Ϫ`b�	s�,�覭Qf��F�zx�&�|B���?�&�i��	� OoNE(��M�
bp(�"��O��d�Oz���O��� �D�=y��Mp��8u[vx�o�3�1OB��$R�^��`i3�IdVB �r�?dC�čᦵ�ٴ����4y���n�ٟ4�IG�DB�����P-�:ym*I�ׁ� �6c��'���'&�k�kC+�����Mc�Ir�'�=���ƒ|�^�{��J���EX�U%�(O��C��Ɖl��h;��F	<�E�ԣپ"+����M�ҜA��ӹ ���
�&�ؒu�>��n��E�4A�"b�Y ��:zQV�8���'�rmCW.WD�<j���P��P�
�z��'������)И���H4Oè�{�'�:��y��D�O��'�A���?���\h~{S͊�p	tK�ES��EK�ګ����Ķi,r�#�&�O�x���y6	��hsDmA�!�E���F�D�؊ `v�p���8yvP(Qs��H�F/���]["أd`�)'\Z`�5ʂr��ť�=�?qו|���'�D�;�F�5�T�K�
����'X� ���-2���U��;O2E��y��'��"=�'�?�D��=lX��f-�6l�<����?��?P�Y��!���?���?q�c���O��(~�����(�LP�t ��5
�D�/p��}�S��N(�dL�P���y�!��~��<��>��	".�j% [�Z`I��	�����X	���4|O���$��B�(�!#�^�~m�"O:��S��k��!34�>�AqA�d�����|��2�6��� ���([ ��Drd�D
Q�D�O����O t�2@�O~��r>]ۧ�M�
f�h�F��2{B��O�4Ѷ!2a�(��$`�!�t�*�:�U�$�Q���AK�^�aP��N�����/��)2ՊD�U��-�W-�=}Pn���+׸d�Q��[6��O\��E��ZYE��X�X��P.	��OT�d�O���0� �GmA'
�� Y�M�=46���Bz��Q �1�|���U`+��Γs��&�'��I�\�Hi��4�?�����)W�3��*S G�I�ZPl�d����D�Of��Ov�0�,�e� 9KfF�Ih����|R5�E/�D��&D:6) ̺�$l�'�qs6�K
rF䃵�I#6@�|�ä,l�l����>#^�C� � 
�@��#!�)d��-�=�����	��	�k2<�����?�(�c`�z�!�$��Uu6\	D�<���B��{@a|�@"�L�x���J��)0� @�E	3��	,
R���4�?a���iT�gq�D�O
�$��;rT)�� +} 1R�B��oJ�� �K�$򐱓��>BDeh��b�d��w�,���>p|I 
��@�lP%*�F
*���˟.ͮ��)�	k���3���B/��;@��A{c�<K�,��7�N#8(d��?�d�|���'����썪�F����*na���'�����BE>e��Rp �h�������l���4�'���c�NR9y��\�tc��^n�y��'��S�I�u�'���'��B}ݭ�i�Q	!�8w���(�	\"
��ãf
dЉ��ʕ�d�\IA�G�`�S/`�����$Cf$�ᧀ�`�`�vA�-h)8�7��Fc�P6	=kz��ԟh6�P�Rݛ&�������i6�6��5';��T��Q%���Ca�`�D�O>�ԟ��ǟ,�'�Z��)�4C�8���O +��
�'�R*E+\��k�?J�8�֨+Z�#=����?�)O�Dcʦ� ��E�X<���Pf#RtsE�I럸����$�I�3���	��ΧEL����h�"�F�T���FT U2F�3R�;�O�uyX�8sD�X,�x)f�ЁU�L���-�OXY2A�'W7� ��R@矔1�"�y��N�=����"Op�����<;�m�1�ؒ�"Ofe��F�$D�����s���g2OJ��>`��]m��'��V>�`�@�3X����F�< �X�öR���	㟼�����*��*k�|�p@��n���~<Ҕ�_�A��A���Q3��r�	�@}�<��K҃Q�t�� QfR�U��&�4�2e�,�nIY��:Ke�F��22E�=�#�̟�i���~���s'0*�bp�.؅�PyB�46>b<a��/v�"�"�E\.�0>���x"��R��8*�˗fl�P��L�y��ݦi0���?�,�d����O��D�O�A���\C�X�)�"���y`�ۀ��7���A�ȝ@A���1��'���<	b�LS �rR���b��W� ��GgΥRP��9V뤭1�HL!���A�@��w?V���8+�~)��$1d����C�L&��'��6-�Op"~�I�vX�q�d��+@��뷣�$nv�Iԟ���ߟ|'���?�lK�|,�����rP�lI�\�'�6M[�U���M�a6���'$���fC'}���`g"P+!��?ig"���	��?���?�w��T���O�(�f'5�Tp�b�6ng���CC��l+@ϙ�.Y���uF((W��	�3�&�mK�#���P��Þ�@�Nʬ<�A���.��s�?M�u��zVl�0�����gn��.1얁/FJ<�%/<DK�DK;*��)lOF}rwIӅ~t���i��A��"O�!%��0?y�<��B
�!�b��1��a���d퉨+�����lX�R�"�@��Z�[LC�I2>��I��9�0H�5oT��@C�Ip��"��k0h1�c^��"C�I>w8�逄/[/A�\���	���C�
{�uC�-[%��ǅ\-�C�5"�xAH7�-�����5d~C�+%�z!���1Q�XZ��  �B�ɲ���B�b⺈YU�K.t�FB�I�%^��pq��/c���� E!(B�ɠ5��!�f/�O�l�	#�Z�n��C�� Br��4�X�7T5	RBӫ-5�B䉾u��	9��
^_���p�.��B�	���0S�#몡�VĕC(�B�	�!��0�	�iA��̔�DO�B�I�R���6�Q	 �1
v���R�0C�I�u��Q�	�r��HA�#̔j��B�I���@�8@g�,� �	 ib�B�I���K5��C�`��v���~B�I�j�:㋞�&.|	 �.I�nB�IO�l��,�l8ԵQb�A�{�B�Ie.���!R^��p�wb@8�bB�	8oD
A[�͘�i��p㇃�RB䉓F��`�u���Di��� /��sxxC�Id���:Q*ܝhC�D��$Z�C�I�\8�BߚC���#Ő�S4�C��2Q&���IuJҤ�#'�2V�pC�	0�,=�3���k8�$%P+3C�I�,�qҲfV:=o�����n�C䉛FI��ڠ_�O|�;RK>U��B��&H~\��7��(�ӆm�k^�C��)q�����1,�S���!�8C䉕L��@��!�?;��%ۀA�X�C�ɠ�lɋ`mOg�(�i ͅ
J�B�	�A�8�N�;,�:p �N� =��B�I�-ۨ� %�mY�z� E�g�C䉍K
�[�.![�,K#oA�!`����Ei����ْtr�S�Ol]`T�Q�|5�� P��}!�D�R��1;oD�S[-@Ua~Ҩ�:7���!@�w>��R�FL.o���O���%凲t�rx�;V�n$?�i�59Rg�V�3$��jK�� ��=�O���f�J� �u,�Y�#V�I�>�ZaGH�`�X���x�`D�p�C�U�Ա��H�|ɸ���f�(RD�������>d]q��/s�
+�����%Xw(���DКS��|@�!
���Y�q�O֝A��O���&>c�8�ǫЫci�p1B AA�̱C�H��9<
�8�N7c��@�'��(��Wu݄���.��Z��R��B*x�R�E�9hm�9���� ¥ju$܏K���'��3�t"OPzuI.~J�4b�	�T�"�3B�1O�(K׀EdLR ����^\��ףy�b���"�#訝�DȞf���J�@*�0��A�����W#����X%`�Ś�{`�x�BШE��4����Q{j:��L ��'iNʄi�+x���`
�/"��%Ќ{��TiHw�@#\�yB�%��!�2�k�lP53�	��B�j�6�%ÜO�R7���i�a{B�ݐ �j,@�� �tn��y�G��&��"��K�.��7��xZciX�s�QcG�Yx�m�n�J���E�}��3r���W_68��~�	�f��E��.!M��jfL��p<�m�x8�5����Q��E ��ќmњ}�%��
\/.�� ğ�����N����
ǫK�2	��$���D��`��:�� X'��rNY�-XE�	Gd<���GK�J��SU�<@kDc���!`,d��Z��MZ�h8��>}��'4&�r K5����k��N>��ϸWI�İ�kк@y���g���{��y�L_,;�	���E}R"	"`�0Hs��V	���B���#"��!  �7	j���$TJ�xZc���1�A4�����b� 8M����@�O^������;�f�ا�L�:�L���'��U��j��s��6���=�b��0��l#&q�g)��#��q���`�O�P�9�d�BE�,���Iu�&y�%@�$`:�0��oH�H�����&Yx�ɰ6�����]�04� D8F>��h85�ƪF��Dx�	ǿ�|�I� ��kx�h��'��'�D^�g�p��M>I�g[(�3��^��ң�
Q�s��#0h<�1��<���N?C`ߍW��]S��F�P������Ҙ&��z���M��ô2s����~)�T�\�m��)�1�r�z�s��|��v��D��䥟�8��w�F�k@/վPT~�[���:�>�zǓ{BP��g�R����0�]�c,-��a�?H�̄�U�GA��u�!�O��I���:V��K��S��|���H�Z�,,��	ڲ8�d��k�-�� ��� r�'����ɓv��AY/�uv�9�}2��=*5<D��&R!*l^Pk�@�'�~��'�J�GB<0C��Z���C� 5��QZ�@�/�{�R؊@��/
�Ѩ)d{���#��Hdџ��v�=�ƨޘXWa�@�F}�d�3(ꌋqmQ0V~����5��@"���1��/����#B���O%̓��X����b�{�m/u��:��Z
�x2��=���{��6|�h(j��H0,�i�T���	�]20�NQg���F?�r��`�O�7�� {�D�+ۿ:�5�T;2,h�*�ΣE6*�L<�Q��lU2���7��hC�m��$t١	�r#P�:�S�q.8���?�@�DT	I�v)@F��8ΓO���֍�<�B�1�D�Ƭ`�ꏪ*]8�ɗ!�8C�<�D�Z�@JqeA�D���{�X�N| @��T��H�A�W{�Ĺ��g8��ئM�6uyU'!���p5-@|�ڢ>و�W?�!Ny �CC�=��0�D��}8�pr��-)L����`5.vF�сF>=�8�z0����,�����~���|:���d��h$�Xy�U�4�h�Z`k��HSĚ$�TO%�ӱj&�4K���*����F+,ͱOVHq���M��`A��իx��a(��O�ml����#D�*VIs��{�&`Â(�K�I�y�L�A�!�5R�HI����^ԚS��9�rX!AH����OP	��Z(���<EsEфg�<�ա��^pj�m��(.�!����5� ��
aT�$,Z�+�4����_���O�N��B���G
��'	�r���c�
8����|�\���Pf�d)���_��q�J$y0q�R�Z��ē�d (srl�[Q�'q�,<[nV����Z�E�����A�N�D�gJ�83d4%� �VǄ1�
�j�`4_:)�!*�I�z�A���5zk�E.�_�t㞌 �ڏ::���$&.��Y ����2� ���3AF*h����N��*%˞(۞<`��f؞2e�]�� �W)g���`�]V8A�aA(a~�p��@8��غjd}A桞�Lw��E�I_�B䉲���%ϒ�>�<#֭Ħf�)��;��4zB�K��̅Qvh6>��X�²$�,q��LY�0�؅�I2	8tr�$U"X���򵧖�_)0�Y�N\� �p�ݨEr���D?Ra�窜;FyVDK��޵r����h�88.ʸa��,^.���?�VU+�F�=]�����ºA����fE��T������@�i�ʌP'�%ч�*7(8xk%�VΨ�
qJM2=�ayZc�)cT7\�I�%��Dz3�'L�����ϟ���y��ϳ�.����'�"e��َ~O��0�o��@0��?F���IC��	Ag �ѥG \O�QruJ�9�t���?���RDn��S��I�g��~?�]�K>�c��>��\ѧ�d�	:��tܓY"�(D+	_���a%��*�~a�=��EH5?0���W�@�����h�ɼ ˀ he��K��P��.	�	���	���������=�F��QF�I������=�cOЦ	�}a��o�]�D��p<��>�d+�%@4^�x9�F!��)u�l�'��)����3� �U���L؆�kaC�%wf����-Oda2��-yܘ�Cߺw�v1�"�R�u�w�E3.x�EeDq��ԛ&�\�"��ĻH��]�Ҩ"�DYH��	�B�p0
��P'���i����;!N�#���%��=�R��0N@@��L](����"�:���p������ƭW�֐�iY�ncH�I-5�n�p��̰Kr�$K��@��&��	&T�RT�c 
�ܝ:P*+��a@$U5|�������I?��� �*�2	T��~����|"�@�Wg4}����=MY8�;���2�T�z���<�ѐ����p<�1��|ن��\;`���o��EoZ���r�oL2�"���O2��N?e�CV?��6� �#"�8�����F�I�.��㉨@cL��B;=�&���n��m,��B0d]� �%y�HD��Q`�&r��0Y�W��T0�����'H�p"���=��a�"sXv�8�ĚNѼ8 �BK8`/�y%�xs,��0@^a�fێ_�@�Z�!j�h
�O&0��'NY=���go�<y��rR�F�s�D`�קE\}B䅳���!
��~���3A���L���iE�_7JR�܋��� �T��0����t� �ڝX
�䘺PX���Ն֏T$]�O	m�	�m�8�,�2�࠻�a@�^0�Ң��YA�#��K����D�0�"�<[�{5�����3gF3n�ɲg��w�ȹJK(Sf��CN��Eʽ?�̓XAJ �S�X�N��ܘ1�Ahl��	Ǔ"�:ܩwk�F٠����R���OM�^[�����d�zrI�I�Td���!|�3sLN�����O批#��<�" ���<�"�]K伔�v�D�o�=�I<)��Z_%yԋ��?�e�������!X�g�H�zi@�T�@�r@�1Zma[�ʑ"T�tI'܁G�k���4�[!`}:&��v�'=\8`@Dx�,hу���|p�(�˕#&�DՂĒ6}h��j���"��9cL\=�i҅������Ƙ��V�"���#���LMR�ɼ.U|�"�![=qb�B�$Okɗf�~Y!�ǟ%jр-;�ǪVϛ֨�?x��F)�E���Y��1���)g"؁������>���3C~8���gBc���A��,mxʘ
�"z3H5����;Exθ���Cq�(�I�zNL�R��+Px�0:��bʅ\�\��W���X��YP��0A䀉(�'#�V�(��MF�I*���U
�L��" �<p� �I�r8Xe[V�܀�z���ϙ�l"Z��pcۏ>��9���7MT+8nm��o�~����kY��|R�*&�L p�`�29��Q���H�,��`�� G�v-�WCh���P�F9�s�l�Yu��X���4��39<�ҷ�8lvNqAvl,-C�8���'����b�7$G�xZc���L���Q"��K�U�@���4X��p�'�+j��yh�N؟��ӕ~��f�~��b޶�j��	w*��!Ȱ)�H*
Ǔan&ݫ KS�`C.�"&���m|��q���"�Vd��N6vy� �[��Z�%�&�X�ȵ���$[��2�ȕc�?��9��F)X��&�	WXP2%͖,��j����`B��Љ �j�9X�=�3���Jw�!�π�Kݔ�5.�
G���2��Ij��!#
$��rs���c2ƒO�;�*
'p�1�g��/?�ڭ U`N�,�s	<����'���D�,LɧjT�@�T�p0�;U�tR��ÜU�K� @���T�_�p<�1 �EJ7߫_|ĕ�ϒ�&����'���U��Q�\b���0����l_�(�"8��� �hS�=�]�1���>�ĥ��CW�	@��`:\O~��bR�D��(�b�[8Z��aH��F0*�l}�M�<tdQ�J<�@�B��ɠBM�Li�
B͂M�\D�,�.��V���/�sk\��=�F��u.�� �nA4�-��
Ev�}	,�CPKW?1�(�k��O�(ړ�RD5t����"߰=��J��t�F�a��3�
�m.��Hb�>[6��;'���p<��w��$��۩ �h4yV���f���ޜȀ��-[�DZ�+��["���6����GW7D#%�лS���"c������i� bzR  ӓ���ɰH}�����D|����}t���(�Gz"�L~sv�ħ~��c>���K=qΒD��ЅB�xY��M�[����' .���R�/��ϸ'	RU����	�� GO��Ybߴ
�4�3�N�Td(��g��"|��&Qʺ�f͉[�	[���=%��(�c3-�Н�aɎ���>�wjYA2(�7c��z�`ã�~BI �Yթt� {��ݒFd����:&�w� ɑF��?��xj��'8�yhՉȊ#r�A@i�';:0SB��C����$d��e�|�3�[�n��)�'�@�S2�W w;�Q��$��w�Ԙ��2E�q�4)�� ��Ʊ*�(�ȓj�>T��J�9��0�/)mj9�ȓ�`�be���Z}��rfիT�Ɲ�ȓk�8Rm�"N�CE�e�\����W�0_��"	W-X�١�"Om�7"�]ˮlJ��ɿc����"OREF��d��92��%sZ�سb"O$���G��96&���ǇFPZ�1"O�̒��V�}I<U�ā�N98Mag"Op�F��3a\�˱���,�q �"O���a�7h�@�K/.�hX)�"O�@R`���+�@�Y�難SZ��XF"O� ����B�:R�rQ�CH@>$+R
u"O��ۅ�ޠ/�4��0�q&0	�"O~�p3�T�p8PL���J3v6����"O�5��)Y��r���a|<��*OR�k��t�6���W/j"P)2
�'�vCǌ	5�m�!K���	�'���6��B��y�d�.��'��|Vo'*�Tz���w���(�'���bcܲ[L�pAK^*u��P��'h�\C���#D����%��f�hD��'��QPq�ʎ-.b�6a�J���'�(9	D�:wRhbg#� WaH�'�F��1O�]�I�/[2Z��
�'���@e��UX"�� �1L��L��'U�a8�'=#����U7����'�J���&/�H��o�0
�\��'p�}J�UJ�-zU��3p�)h
�'9�4d$0Z��G"b�H��']P��c�&���ቖ�\}d���'5v��nWz��X�qO�)Uؚة�'��ij�A[�^�A&� ����y�
QG��i��̊�"�L10T�L8�y2lpǖyAAI6� ���6�y"�47��-#����su(���y���UI!d�ф1r �D$�y�D�
���+a�� k�4�8�����yZ��i��d�0��Lx#A��'H���!ܝ	�RQš&o`܁��'nԹ*��P��-!%C�+vt(<"�'0蘹%�~�<�˔OX�W���
�'8,9�DӝIE���Um��F1�(		�'.�uk$%4D�8��fR9k�L`�'�Z�	�M7�Q2�BZ=jB
��'���:�cM��C�S1`����' �,�sN6�\��7O��*5f���'�%�Q�Y�ax�l�r�\�'@���
�'C�4�@ga�D�1��	�F��y�G�^xR�2�M�"W�91�
��y�)�jJp:B")�SU)�yh�!Wu��C�֭`��t�X��y"��:��e��""d������y��V�6���Ӥ�b��YUM��y"ˆ�=f��EʢW9�Y)�b��y"�f�������Mi���)C-�y�&	z*U��C6wr��b���y��� �.,��i�C��聭I#�yE�2}4A�PnK��,p����y��L�J�(Ϣ>m��2����y���,��q�����z �Gm�x�<�M��K�C'��ax�ˢ��H�<�G�G&L(�0�	=��0��D�<	s
��"�J�Y$neѪ�i�<��GQ�u����~r�4S¦�n�<����+��#�m�6��@�i�u�<@��w�>�(�g��"���b�^j�<�֮47$V�� ��joV8�@�c�<Ifg�>��s��H#$��i[U(�`�<�m��@�!��!cw��J��A�<��ˊ=x-z	A��a��xi��GW�<i�h�)>�~�i'�K*�ʉ�g U�<1�.��	�dT�f*A�c��A�MN�<A��Cx�i����)�����E@V�<��œ�,ʙ�
�4+����cLUQ�<��ɮi`:���cҨ��"@�~�!�� T����՞\&�#��C�Z��`�""O����aт�ūd��d��]I�"O���%mV8s� �R%3u��"O��Cp+�O��k�-^�1	���"O" ���33��������b�B%"OVX�`�M�tpQ�4'<i?�9K"O.��OJ�^~�]�b��R�C"O*�ѣJ�!7�$��#�'�!"O��+IF��h����F�I`"O��ʲW�+F$��.ɴv��x�"O��"N{H3N�	q},%�Q"O��!ሞ$ .섉�M�Iu��H1�U8�X#�_hW�u����z�q9�!D����%2hr���V 8�B�$�=D�kTgB�cYp#%�S�S����<D��X��ܓRHb+T)�����ruf�<���ӗ:����0A�{jI��U5��#<!��$�O8��+�kP�����6��&;D� �(�*;x����SI(I��U��hO?�$8/�ZR
�=%���1�!�:"�2x�`i�"�4z�Ɛ�P�!�Ҍ}�����B�؃��s�!�?9��X�s�]�y�"� ��6�Py��Z�}��x[0�	uT�f/ڢ�y�g@�Y7	��J��~�m�vg��y�L�g��r�(.n�.����O�yR��=Po҈��,U�5^2i����y#������Uh]5۠if���yҨ
�`-�����bA Y�Ħ5�yb�3_6ܚ�^�P� �,�y�B�8�\�b���,V�����\,[��➈�S��?��%���b�G�؞R
Q�<�@nM06��1����
M����N�<��#Լ}`4��\�@��q�ªWs��l��Ц-�reV�m�r���3wx4	 �4D����	�nIX��2w�Fh���0D�̹WGҷC�,��M�F=�<�AB0D�lS6�O� "H�@�M.|\! �/D����J�-�$e���(XV� ��.1D� 6��Bb��2슨��ԫ�,#�O��'��BGb�	�p,3�d �y���cӓ��'�.5�k[,P�*xiPo�w␉K>�'qOq�$��u�F�-�h �_&�m0"OF�B��DP�� ��2;���9�"O
���-���t���n �R+.�S!"Ov,ȳg�W&�4�[�".Wb�<� ��:9��Àeت�tYH�aP^�<��/N=8�x�0����iz���<)ցU�i�%� iJ���!��mz�<aB��mf@	+���rQi�Ev<	��n�2�74�`@�����1Ϙ��ȓ��`p�E?eJ�*"(ŪR$r�Gy��'70,��	��2{����N12�z��C��8+�B}�rf�LR*yP�`ψN�\��D#?y�O\E�V,&���Q(�4;�X��"O�ywsOJ9W�ߪi�����"O�`�P�3>¬�R���o�p���"O��e`�2G�g��bx$�"O�r���n�jx�gCA}@���'��F��R/&��d2�оGʴ��g�.Z�!��G� Q��d�H����G8!�8�p�Ar�h
�9�@�j!���6-`��R����<d
̐�O!򄝯d|��%eR�%X�`Q�l�%!�!�� ^3��B�I�\��	4x�6MA�_��o�_�'�Q���d��!#�TMP���t�>�@b�0��O�6�r�(r��I�Qͳ�a^��壔�B�!�$ԝD$eZ�b֨^㬴QW�؁x<�{RX���'>��x�J�r���T��3�F���Io��V�X����{��T��׿K&��ȓv\`�/�"F�=a_9	?�%�ȓ3��={2EWG�傗A@����y������gx�(�,H1>.���5��J�IQ;��;!A߃N���/�PA�E��1'�=QUϨk� ����'�ay�H�'Y��Y� ��$� �S`ڶ�y���0ʤ,��4aA���y�ő4;H�up����C&C���O�#BF-շ%��9����))�TY�	�F�<i" ߿�
���$/��M� d�l�<a��P^�M��'� i��Ej�<YQ�	� �#�eM-^P�HU��i�<�㹊`k���"����-��z��D__��Tc��^���BG�G��̅�	�>b8���H� ���C6���pw`��Rn~j�< �(��c��%8a�&e��yB��8[�����g�$+�qb���yR`�4>Ҟ}����\8��g��tX�蓡a�V��x��&U�ѹ�'6D�`�O��z�Q��o;�(KT�1D��פ�$(!H�����|0��/?�
��P�!�MW�\,&��beP�H����ȓsӈ��&�lH��$Q-����.�ְ r
��|Lt@*V�JX\�ME|� ?�'�Z��tϷyT��!㉸p���2i@�a厓rw�(вG	1D��������Y�H��#�#f@��0ReB�<�h��p�/\O4,�=q3�)X4�-*]�vg
ԋ�o�<�����>���L�
�BQ�ŋ�$s�Gr��hO�Iu�
'�D���p#��G[Z	�@�>�����ba�6��p�7�_."
x�*���s���������a@�4lE�a9D�ܫ �\�^��Pp�#�/�d%�r�7ړ�0|�1j��nb(���>�B�:Ņ�Q���'���0i�E,҅�����P㲀�	�'��Ɂ�Q��b��C<_X| ����Ob�}� '����8�a\72�(kW�GK�<Y�@� �0�ar�7 K��z�Ïq�<� b A���C��m�ޡ� Li�<��M��T�v��p�Z,6�B<�Ea馁E{���i���9���4' A�$�
 :x�Qh�'7�5�AW&
�������:��'���ޱ$���Z���}[:T�	�'�2��a�ɜ3ΰZQA���`��'�*Y���j�F��H��
& ��'��h��a\�j\HA!�	:����'��C�ۊ]�]�Ι
��9��'�>�ⶅ�"z	&
ޤ�B���'�!Z�a�z�$`ՀB�z'4��
�'+�%P�A�s��#M:s�`�'��cLv��do�3r^i�
�'�d�`'��@J2E�4�K�g-��R
�'TMA'l�ʦ�d<^���'����Q��-��\�'� P�t���'���Y�&
�n�H�@B.Gۊ���'��-���
�7���:@ܠpӼ	��'uX�	ӓ~��<�#Q�6�0B�'5��R3�/~}:�	���7F9��k��� �H�a��.��͠ �,Zצ��!"O�����;7�T� ǆM�z��m�P"O ��ˁ<��`U�T����2"O�91���>�J��i�%j@�e�G"OJ�@�j7zua�Ɍ�bD�ؚ�"O�ii �Gm��i��9��9Y5"O��)� T�
������hɀ��6"O�%x�-�;��R�o�k�R�2R"O,�2는<����'��X��̛""O:	�5�L�L�d�6g�!A
j�"O�`��s]�4�U25
�u"O���&�h��:P���_�RQC"O��d�IJQ���"O(%��i�X��b���n]�"OL}�#���ęBL��&���"O��R� ��N%�d�����f"O��P��2���[�ǳ+{�e�"OR���@T	 �Q�f��p�ԃA"Od�cl�~A$ִTJ�
�"OI*f�ڮ?�f�S�HH?�$0�'�ĥ����h�ݲ"
��H�X�'���a�,eˁ�:WԜy�'[ 8s�gL�y:���ƅ�+>N���'���a�p˺��
��y�'2v��ʉ�v�,�b	L&����'D�!"�L����I��-3���!�'��DcD-�4�QRP�^<aΖ|��'����'+&�d����ņN�Y
�'<��׫|&�@2���#H�D��	�'�p "#,�z}4��&�W?I"Xy 
�'� #Ӥ�rB�8�6ď�Is	�':L��瀧0t�e�V7N��8	�'VB�rU��`E�HqO���'v~ѣJ߲�x���L+h���'�b��f�ýfХ#��)��0	�'��		$� �A�㇌��ɣ�'�*.н09h�����3A#����'<����M�K�vZ��\/j�`��'�4
��@�1 ��X���!�<�8d���O).��C�IÊ<N!�O�<W����M˃�ݠC��}!��ݱ6�q��·/����Z~	!�D�,I��fK���Dj#�I�!��cf����0�����*Iq!���o�jx A�
�\������C!�$Y�Oׂ�������0 W��!�$�&Qж!�.�+=Zpె�7l!�$�J8��E�:O>�yu�I	b!��9Z`D�!n�)��(s���]���!5Q`�J��b��Y1$�P�y�D�����1���.�8Phȓ�yB���Z�4` F�|`D����y��X�y�HR�@8G��ݪ��Հ�yČ=r��{ab�D֜`���yb	�m�
�����K��؀�
�y�I�1\��U���J��h�`�'�y"�	"�Фmէ��	�3���y2n>p^m"�hU?c�)�х�yr%�H�H�E�%�4���%�y�cS 6V�d�����0hL�yR�^�v�ň�X�N��w����y�IX���)��		7`�	���y2k�)cv�u薏[�z�N`8d��y�g��d��`Xä�<�dq/��y
� ���Ũ�r���f', P���"O�ap��
�n��j�CH{� (�"O||C���+b���E��&Mb�"O�$0�K
���*ឭE&X�"O�1`g/��eol����<6@<	z�"Ob���5+,�՚�e� X֨U�"Oʜ�r��4϶��u����6��F�<�LH�ad�b��:^�ěU�D�<�p�L�J&ʵ��LS\��V��B�<�ƍ��#��'N����`!�{�<��Né+�0�EK�-]�@T`CB�<��^"��t�\�e\aJ4��|�<�1��<H��B�Uz/6I���UM�<I0k�;1 E2�dЗ Z(Y@�L�O�<��Y9^"B�R�脖D�:}���BS�<��ШF;�P�6IO s�@P�<�`�Es�HQ�E;�IAt�LT�<��`�a��j�X6ؕА��I�<�P���4�USwȋ3O���eMD�<�E� .�\�F��B;� 	B��I�<a��H�Fc����,'L��˕E�<��/����������T�"�"�@�<Ad�ӞVZ؀� X�j�$Qy�<�a(^)i1Nty3KRT�T�D�k�<�5�\= G4+�"L�s�D��#M�n�<�p��]� 	bRa� �<e���g�<�@6e�8��w�h�jq+�F�c�<�Ɵ>}�ԃb�	D�D$GZ�<1O�0�����S�\ŪQ��Q�<a�/޺jZ~�VG�SzNT�CEYv�<���9#�x-�0�&�6��TA�n�<Q�-ʊ^�^�k��o&�����"O�P����x�
ѣ��p�QX"O�$PG�� u\���ʟ�+{�I��"O��"�@-��I��Ϻ#^��҅"O�����#@`M8�A�/H$y"O�P򆅗~K.���ʒ�s+FĪf"O��$�Y�qK� B�+�
>F���P"O&��F�P�,��h0��<4��Y"O�������d]��.e�p��"O��+�<�`�8�='����"O�{6!��/9�Q�+�O�����"O�bo-n$͛3�pm�=�"O>��-G�}����)pW��r�"O����pO�y��
L�8�"Oz`Aէ�:Ijz�'�O-@D�r"O���KE�*�0y�p�W�z^a��"O�p��(5��Zw�:WT(["Oꍡ�&�
���\B��"Od����n������Pvt�ɒ"Op�!�,�+)F<k�fwzH�j"O����ǆ#v��7k��]��dy5/-D�x9E�ڊQ���UO��ㄜ0r�)D����%V�Aް$b��F>pƈu{�&D��`�C%r�8��È6'Rݹ�`&D���g�%>ܞ9Y0�[��E�q�?D��t � j��{3˃�Vn�]K�&?D���@@��b l������|����"D��r�p���V�����b,D�Hz��Y�J�P3&,�����M6D����^*g����hB$T��a6�)D��JTE�.|D��#�� �#h`� �%D��30) J���A�G�0�\�Q��8D�`�U�]�m4�����RX̀�`"D�� ��wÞ8Co,+p��tKhDZ6"O6-�q
�9����G�̱`J<+�"O|�a�̀>Tn��j�Ҫ9()�5"Oҝ!"œ8&�*M#�"��+0	��"O0��_�qM,����ۺi����"Ov�X�Dߦ͞�ɗ �����xt"O �b����P�R ��RS�"O����.���GN�5���6"OV��eaR�a�4uy��BI��$��"O�@ꁭ�68n,��R�3u�0��"O8��C(  ��}cA�\�?�I�"O8Ļ��^�zqC�
�]&�W"O�|kO϶a�
�j7e�-\�0�"OB���g�kH�X2DE�P�"O<D��Ļ]���A�X%z�Ht��"O�
�kſv��y{��[p�V���"OLPQ�=a|�kG�ĥ*ٸ���"O6$��Ks
6���H Wil�"O�R�	2qxr�6葍-J����"O�����6��DA"�J(^�`�� "OQs��ʲ$�5igC�s�Rd;"Op]S��m!z�ӣ��"c�x�"O��)�O#@�l�Z�/d�xE�"O6�:�X�~�:�ra�B<~6��P"O�ݩB�I�>�N(���ȠT{ �!�"O<�1�J�h�P8a���gw*�v"O���b�N;)��"�"�jf:]�"O�m�'�>"-q�"ʡdt
��"O�tx�"��2�n!'���N�i�"O�A�M:r[V(I��V2�@e"O~Tb�U>����LV���"�"OʙB���h%�XI���<�v��@"OKݶT������B�P�@5c�
�ybm܎!ʜ�p�/F[�L��lʐ�yD�9#~Ȓ�N?-TxA�VE6�yB��?}h�5A%�F3k�p�F��y_�g]0��%I�<"�Ր�OW�y%P�E�X]�r �%h^!cP� ,�yiD���a1@]�� p����y�&ʓc�� �᜛�p-�gjО�y��O�cJҽI"��+,P�C�@��y�)�12�n��񌈅GLqr��y",�Vz�1�֋@	�� Zsl�;�y"�O�G3|Tb�b�2iqb�8�	Q�y�kY��<�z��=ƨB���y�JE� �1[��¿W�m��g�4�yb灨q��e�e`G���)C8�yE��bK�D	��ƣ@�ּ� ̗#�y�!�U��"u.�%����9�y�韸�T�PE��&+�	���y�#G. ����H�l,`��2�y2@�^V�,ۗ�π==�ᡶ����yB͜�U6,��ėC%���%/�y��޲U� ���	�;5��Y��g6�y�?(b�ݪe
<&`k�b���y� �:��,(D ���(U4�y��m8�Z3-O��(���+�yrF�I!�$X4h;�l��	�yb�ڀ&�R-���\�f����/�y��է!�d��#�)�J\j�'��y2m�J�،B��C� ����y��Η	S �`��HԀ�F��yB� {� @�]���YdEܙ�yR�b�m����F��PQ7 V#�y
� ��%�,�"����	րZ�"O��'l�eZ\ ��Z���@�"O�qC���8-ɃJǟ,
�0"O�pxf�_�>o �z1��G�t"OJ�Z�CZ�4�V��c�&�ac"O� z�

$0�jTؗ�D���"O���`HS�Ob JQ	�$�R�1"O�AYD�C=Aa�碘�"�ReY6"O�����%�H�bկԥV[z|�`"O2 y�*mi��F��*��;7"O���B�G)I�tY��ǠB�M�#"OBU��%͜~�h�4nΏit��"Oسg+�#*M�})�fϣ)�Vq��"OJ�
����8~�X �� �~�9�"Ola��d��!kç5k�1�"O� ���	3��UZ��d�fI�P"OX���d�"��p��[ämZ%"O!�%M��>�m:�9��C�"ODA*#H�-P�l�3��6v����"O(ɸ3(�<c��x���E'[�Aw"O�����[-?VB����NG���"O@��gMW�th�� wO�
�"O4�`�+�I�X��p�C4><���R"O���.\�
��d�A�95��"O�8I���Z'~e��0h9  �"O U�AdD�6�fe
�ט5��k�'J�{��K�P*����}x
�'��TCטV�j�)�YF�	�'�zفv#��b�fHRĉ�g�$��'`�l���F5I�-�D*̶���)�'�Ū�&�0Y��Z�Z�m�-��'rJ%M1t�^�T/εZ����'�ҡ�Q���5r$���Z���'�\�Iĥ##l�� ��V�Y��'"�T�G�ܛK��DX�[�w��k�'0�бc�Q����c�5�'mbh�G5�ɚ���8a'����'"���@I���+��%�$T��'5� `�.C�J�W�M;�`�Z�'�C��@�Q	tlc��� z����'z=
�c� ?���Ń��eMF��'������ �N��!�3Ұ�'���4Iɲ2�8���BI�B���k�'0�JV�
�b-7��e��!�
�'| -���K���kV�
� P�'���pŀѣ^XZ���?2|jH��'���$��)�jE�TH\-���:�'z@�ز�N:
�������
:|�ة	�'�������7�� Ą]�B��@�'$T�b"Q�
�:�(S�Ϧ�����'�"P��M�xn.)��˂K��i�'��,�k���a��(H�F�%��'cv!rH�4� je�K�r��i�'��AR��/�J�5�(dpd`8�'�`�h��u^P�D��k�.�k�'��j#f��7��MH���,a����
�'lfٱ姅fp��bf\�-�*5I	�'��%S�ņ2U��¯����L��'�6�D�ɵUDJhIVJY�(��'��i"gC$s���ť�(�Ę�'�`<�4*�2i�M�5&T��
��
�'�,�i�����TJ^p�&H�	�'Sr�r�����UD�%e����a:%��i��g��z0��5��8��S�? �C�蒄e�j�z��4)��0"Ot�{&M�; ܞ��+�,�@9�"O29�G���i'Ef�l�#�"OV�{P��������NZ��}{�"O,��tjM���Q�b�)C��a�c"O�  ظ\p~s��Ǚi�
dRP"O>�.D�́�!mM�UnH�R"Oz�F%ą]�lT����%z 戲�"Ox�"r≈G�� ����v�(��"Ov�SJ_%V��qB1d̊"���y�"O�y:4E�6�d��aC�#M�(0��"OliyC��
���z�
,2�UU"O��2�O�k�0 @Ԕ!�,4��*O�9��ޭ{8Ba�6<s��(`
�'�J`RAg[�p��6!�'7��)
�'Y �q[�gMv-�� j�9
�'���P��C�R��s�#��X�	�'���X'��D��E<
�qH	�'*�`SMGz�֘y��ڌm��	�'5�Q0�
��R5��8|�,��'R ��ܞ2�F�q�̀f���':8��;+P�hw
GI�d��'��i��F)n������?[ո�'�E��nd�H�2	�18�쑢�'
������5����I��}7�%s�'���խC�(,s�#ԍoB����'�"�{����վ3����A�y��3=g|(Y3��[�PtA/�y�I�n��Ӵ��Q������y�HIj�[��M�Ic��#���y��(�B�;uG%?�UJfI:�y��Rz�و2O�$A��pF@��y�MȚ\�X�*�@�p@ᒭ��y�d�;X�� q�\�?����n��y"'�?K̴�Z�AW�c��Y%h^��y�E�N}hSeU#e��@A��=�yC�Y<&-�@h��E�G�y[9S��m�(�V:�E+�Ꮸ�y�*�	/�D�b�̉�J�0�"w)�'�y2�L�|��ؾY �ٶj�y�K�sJN	�#�#_���K���yr	S_��5B`��[�z@A&P�yEK�VN�9W�6	��h��_=�y�"K��f�3dD��gD�ybcH�1s*Uȱ���5�吴�P�yǓ�^����,W��*1�"��y�c�k|B�
FHW�}�h0cB�y��V�v��/	zwxe�@���ybgٳ'�H|�aDR)<���^�<�F�q��I�1��ve~��(�e�<�`�܎;�����F�C��	��/^�<��&շj[��q��2��љ��M[�<�2��(��E��z���.
Y�<9�fʬ\��S�'�����q�L�<��U�
Ҟ��d(��5�.�؁��J�<��-0Xb�p����|�2�x�-FD�<�_Lak5D*6G���a�Sh�<����y^��ˉW��b1'�d�<a�唕���Nಝ��^�<���
K��z��ܞxܘ��BF�`�<��`��8�K�@�y�X���H Y�<!A��v�&Ѳ �՗��
��W�<-|�UK���@O���b�ԎD���o�4c���
��n	>�l͆�S�? ܩ�J�;5Δ۲��:.<��u"O�mٳ�W< �mrs��[-�a"Or���wN)�BJT'|�D��"O`�h��J81�B���c	,x2@@"O�1Z2��?��A#s��:0�y�"O2Q��)�������kF"O��S�"MB"0$�$m�P<�Ybc"O.�(��o��LS�U:0f�"O(|	p��?Pӊ����	V����"O�� ( �V��W*�z���"Ot:�?W���r]��9u"O���}�l�ʢ��1TJl\��"O� �!��8a��4Z�M�i:�,�"Oޙ��J=���䋃�{�b�cc"O\TAw@]	̼P�c�>!C���a"O�h�5RL�a.�?A-�9�"O�͛#H� �!8�#0{2���"O4���JŐOz�$�p�ʨa��d"O�����,k.�=���Q��D��"ON���4
�����-U�o�^ s�"O���P�[�P�0�(�_8(��"O��Y���z�Eb�U�@u�}�"O���c�r0^���ЋIr�'"O��)���q¤L�D��0zh���"OBW���,�p�D.̎M �| �"O��	�)Nq��q���zp"O�;A�X|���bK��y�R�c"O<�3���:*�謲�HWd��h�Q"Of$x���Rά�3!�������"O�qU�F�RPh�q�j���,��"O�hhdV%h-�S@g�� ��"O�w��5F�s��4^�@�J�"O�]�T�DJm�m���`��p��"O��ل��#�<�h3`�s��[�"OF3B+�pLh�	mb�M�1"Ot ho�"��P�r��5=n�"O�:4�R�"�#c����b%���yR $��jTBȌM4�h@R��y�ܰ*��xڵK�5u}Ba3r���y�@�(DX�C�8kr�	A�̑��y��V�hy�AH�U�|J�#��y�
I-/�b%瓂>p����o ,�y""N;*�@@�Î5��H!3� 7�y���XD��{v��/<���a�i��y�DL'3qV%ц���8o2�(���y���:�ޜn88�>��Q�0�y��S2�j��՗7��p ���y�	�Y�䬫&�˱3&������y�OE���(x�k�3�Z�XWoH��y£���	��j8>��+֨�y,�2��Y�D�%���æ/��y�hگ���hb"�;}�\|�J
��yb��#ԉR��ɾak�<�m��y���	Q���bQ��x���F�*D�����0<r��լXGt}��,D���#�Hu����$���z&Dܱ�*D���� _�W��)� J79��H0�-D���T)EJ��I�%��	��(D��B'�4R���.��,w�U��'D������ra�W��(p�`�� (D��)b�Q�8����ˣ7KZ��J D��X��<]�(x�nE�F�k�#D�D���A�}�2��WH4U�0M��)&D��:K
�p�+�`�yc����$D�� ��'�ҍzJ\��D���t:�"O�9F�����K��	�7��R�"O�x��2���$n�?q��
�"O�@�'��+8X�%r�/�5���A�"O$|�b�SI��M���#!u��ӧ"O�0M\)Rg$d(B��+~��M1%"OD�8d��tZ�i�IH���D��"O�8��\-^�`��T�\� ܺg"O����ֻjS�4�#�6�,�QA"OPM�G�k���R���E�����"O�9�&-W$!���zp�C8cb(�b"OrDr�BO<TU��b��.�8�y�b*p��1	�
��,�c�E �ykWI�����c�n��MY�N��y2�/;���Q��ʁg��H�' ��y��3j��������^$k���8�ybΊ2#�� 4��9�xq����,�y�⎎7L���!�"4�	�[��y�O^�RcT� 5�՚) ތ�g-���y��<-������~xZ�dX<�yNՐ}�����I���!�7�yaQ�-�Z����4�fY ���yr�	/Tf�5��vb���Α�y�hۍ|F�a���G!I���֕�y��D^L�4����`X�:�y�h�?�l��fB�θ�S̖��y2��s�P¦��u�[�H���y���]#���F6>' (;"#M��y"!�,/	P����,*:Ъ�#[)�y"&�s���9$'vE.�D*��y�֑~����.XK`x�&EV��y��D�^،Ԙ�(�?kvm�w,�>�y�%��M�������y	���v��y"�T"w� ��Ԣ�r�"�	���ybi�Q*\њ!��^��a!E`O��yOG�t�D��Ћ�W�l�{�'���yr.��_�H	���:�٣`+��y��.i�n�b��%��1�'��y��*;.5����` Q�N]��y���7oI=sq�-bN�h�v퉉�y���Irl��!��!��dp��4�yBlD-� �*G2Ϥ1��.C:�yB �&~)���c��oL�����!�y�k�9"�R��a�i�伒�cx��'K�bW�x��S�-);�*��a�%D����K;~�d�	aIV�*&��@%D��
w*R�pP. Y�`A/h�9:@!D���Hʱ�rw�^�r7�mc�� D�`���@�I7�T�Fi��
~)��f+D��G�K�0�Ж@[+[-���&D�T�%o�8�qa�ձ+��eT�(D��[Em�Hd<���:!����f�9D��j��71�I�#�R�Mf�He�7D�T����0��X�M#t�^iZ2o:D��� nCy̨}��L�W �h2A;D����٪n<$ͨ��C�M����6*O�՛&N9
0꘹a��6F4�F"O�p��*��m�`�K�==�1"OƵi�oLx�0X:�c�;{0ɋ"O��S��˩�2Ѹ��x���kE"O�k�(޲(����(���sg"O<X9 ���T+��za�E Mk�5@""O��:ԅVf>,,�@�����sF"O@M�p�ކm���cTiDZU�xi�"O� "�X�cB�"MP43�IR�5O~XcG"O��ۗeYZERQ��Gŭ38VI��"OPE�c�^�#��TP�&��W|���"O�8H���"Iب��B�cc��`B"O<!	1��.��D�C�)����F"O]J�Ǝ�,��i 7ȅ4�0%Ra"O��1q�[p�p��U}�fPB"O�ЁgԿr}@��C�� w� �	"O�abfԔm�KubCZ��	��"O��@F���B�qq��Q	.I9I�"O�إ�֙y�t}���?sG~��G"O\2�(P�H)�r������"O���e� �C�@�����!hN�T��"O���e&=��3��8D��Q"O>��$B��a���3b-נ�y��H,"���(0!Rq��ɇ��y$��N�L�j��Q�ڼ�򦒨�y��+�5�&
�>��HUK ��y�)ߊ;1��薃r��S4���y҅O8xJ	eA�h/�:Q-S��y��A:B�<���LK�*�0!�� �ybcA�D؜0��$M~�|rQ-Q��y�	 |yb����E/{켝 Q(��y��A�2�5�FL�"m�j<�G�;�yR��e�B�k%,	9���q���y�'�(&;��`QO.4?��	����yB`�]Z������=%�,�CE�B5�yBm�i�pC��Ô�^�"�L��yb�� �����.M�f9�yBo;}�`=@0������H���y2"���QY��D�{�VAbGH���yB�F��(��Ώ!��҆G��y��ՍO2 �cM�Qh�R&��y2X=_�н�7C���n�Е-X7�yb�wPQZqƞ�G`��#Ή�yB���QK da&��E��԰',V��y2��0:�Tq��G�%�HT�V	��yB�F�NDl�����!��[�&�y��zI��pǫP/M �pV-�y(���X4x�l���t�i�"P��yb��B�l�A����t�6J���y�)N��8��Ѣ}���0sM�-�y©�� �ti�K�(}��i�ыZ�y���55��C�W*xҨ-A��+�yB�Ό(��T)�D�̭���=�y2�A%220P�aŖ)�"=��!�y���r*�sr��wU&��u�Į�y"cͬ��*"��&"���) �L��yR�P	��`!�M�k�ǨI+�yſ 1 nL�{��R@+A��y�BvR�` o��z0�Ӓ`���y�lJ7f����p&�����Q��y� Eze,,4�B�lD�1��[#�y�O�Q-(�a"K�]�LiS��Y"�y���/mɖ �dL�dz�H��yҨ]'a��9B�O%y��x��ٸ�y�L��{�@���I��Hx�uP��̚�y�&"Tb��-C���a��ٞ�y��ƿ6!��5��d�����&ԟ�yR�S�<]��x�j=X��,�"� ��yBǟ7&~�Ee�F�Zɔ|�������$�<����h��ĝi\��ydG�"�)Q�+%'�!�dI/DT��3C˙I�>D+��ĄL^!���NqT�4��!o&��R�ˡm@!�� &��wE�9�̔�b/B�T��Z�"O>��U��g�|P�n��D�z�"O���a%�#�:���
�ND��"O�M�C;*iC��T�]~fP�"Oj�"�g��i*N�B+Ŧ!�����"Ob)y���{x���n� �I�"Od*`�\�o�а��Ix[�\y�"O���M�Rq�Q�W��>,D�bv"O����Βm2 �O��'% x�"O��B����=R��!D���D"O4Y��OU4\��	�s���h�^�P%��F��'̈ˠ�� �ܑT��\�x�8
�'\�%�#(x74�I!�L�	`�'6`�"Չ ��Iu�iI��	JH�<)pc�?s�
�'�Q�h�R�WG�<��n�2�fx��H�-sb�1@a�G�<�T��i�p�:����kz=9u��j�<qA��<f��u�V͛� �P��*Qyb[� $��|�5"����sŎ ,y<!֏�t�<��#�a�LВ�ܳ?��0����z�<�����D�F#@�=��=�hZt�<qa�-�1���.(���)��s�<q�J4j{B�b�
�+�� "rJJ�<�����g�Lpsb��#xo�4p�GZM�<1�M�6�"(�n�8Z��5�MIpy2�|�X��Fxң�*AϤ�3���Zy
"�II��y"��b��)CF�}Q��#���yBO
<�$@"F�ȴIlnW��HURB�	7v��T! 
��=� 85a>'`B�4ej�Z�ەaB�I�@+B��2B�I�$@�K$$�H�@yYXB�I/j.~6		� �G�� !�$
�h\�:1�ƟNƊ���I[�!�W42����&���T\�Ү�l�!���P��a�n��>�	n�+v�!�Ds^�`�52�vP5���[�!�D�'D�yC���%>V<1��J�0�!�']���[�;&a���.7�!��T�x�����!�1KT
uH�I�_�!�D�6
��p�V�L4[P3&�!�d�]�D����Ú�%J�T��'��� ��7N٨p:���=S�d	�'@�e�w���=U�ę�i�N*���'��%���T�rM���!D�	K���'��sB,,�t���^6
���'�4�����#e��!�(�/�ޤ�R�'�a�t#ԋt�q��'��.����կ��y)ԙ+������
-Se)���y§�#B�H��p��/z�0�XdDG�yR��+o1��Q�Z�~������J��y��K'��#"G�t�4Y
�B�y�$� �X�0��M<g"Vx����ybU�c���cq!�%M�$� ��ա�y�m͊gqFY"#ݜGx�S&%Ś�yb	��Z��	�1���z����y J3X`q(��Y|�5�ӯJ��y��ݑޚ�	@���N��`��-^��y��Q�%j�11�뜈e
� p!�$�o�h����TJLA��~�!�¯x
B������Rsl	q+�7h!�WX���p �YWڀ�U
0 �!���Ay\�8�BB�}�� ʦ��L�!�Z���"����4��2�A�#~'!��ۖM�������J��H#rl!�� d��G���B�R"�{�^���"O��V�����Z���=����"O\�C���2�3t.��l�T�b"ON]�O��38�Pm9}�DQ�"OmP,�+9��Њ!�Z n��t�"O�p�gbߚ{�N��2�LL_�"O9��언�L�ەQDC� T"O���C�_��H��!�7:΅��"O���tbٷ�P`v͜w�i{f"Or�IA� ю��4��H�d;�"O�ԃ s�tY��C�^���+4"O���E ��%�g�95 X  �"O�����ư&�.!7��=<�֩��"O�pHBń�M+D����-~F�� "O��X���?nT�!��	�H���e"O<Q�AIHDʔg�5GPE�"O�3	�tD���剀=j�|aX�"O<�G�R=0ɮh�Q��P "O �e�Fp��ȂFI:ݬ�f"O�d{��9R��x ��$�6(*5"O�q"�͙�Fǀ�l�0'�ܛ�"O8�B��;s :'쇃|�0Y�"O^1`իQ7ty��YgKHnd�q��"O�|@���[?����q���"O��ao٠PHLQ*���#_O^��"O����62�zɣ�c'��"O<M�%��
-�(d�ѢT8I�M1"O$M2�勳~�J�z�a�5����"O�ax�S�T�RFK�!3��$SW"OF(򧚸'���1�W;��(��"O�0�G�F�5�V���'�"\"�`B"OƝS�5(MzV��E�ۡ"O��!"�=hՠ\ C�?;���"Oj�W�Ŝ�B��	Pu�"OB9��!�= /vY��F%B69�"O�ԙ"��BP,,aÆ�Y1�q�"O�(p�
���&!� ,lt��"O�T��i�2~�:��2凄jr$��"O��C�Z=H��#�C����t"O�e�7չT����c �:_�0�i"Oz�S� �q�l\
v��&�^��5"O�(��@�<^��P0.�<lp�ؔ"Op}X���=���c�4����"O�0c��-{-���c2Vp�b�"O�)�)�/^�8��c��9��-��"O2�Q��Q+j�Z<�B�A�/�
	�"O�8 Sb�0j}r� +E��Cd"O
DC��|`PꐧGÊ-:q"O�c�%��0e~$h���P�*�0%"O$%B�9>�0�q��Eq��@e"O6�Æ���\1��9�Z�]����"O�P `�_j�^�˔'�]�4u;�"O0e�@OO]l�LYBe:Ax0pd"O,@��$A(F�QK���+J�cw"O�LC�DaQ<Iڀ�M���)�6"Of01���*�xP�aQ:L/b}�"O��G^q]�tBt`��$}�!"O�EX �Q�Kwpd�Do�;��p�"O�=bW�%k#�tmȲn��EY3"OB�u%��<���8�K�=pz����"O$x�6�Z�>�Ɖ�]k̘!B"Ot`�/�T�h�[��v�A"O��8��OkX� a��1?�D�S"O���r&�6^-rM����h���"O� ��xD�	{��A: �T0L�"O�#�Ŋ>b�vM@S.�ZΠ��"O�=�N�J�`	j�l�?sYb�@"O�Q�ns,�w�
2&\���p�ȓ�x%��J�;(d�"�6|�����%�a��N(bZ�0J爓���0�ȓH��#R�,K�Y���W�r��ȓzN����F�+'�T�k� dn���x��Ҥ�*��pcE��Ն�g`btQ�E,|�p���ԋY�)�ȓcyl �(:�H� 4BZ;����{~ez�-�-B4���?@[�I�ȓBD�����$:?����E�0`?�ȓc��P�E)J!��b�遳�݆ȓj�*�(��P,J�L�bgN_2wRĆȓ������P m�R!���_�आȓy|�PWl�s�ʜA�㖒/Rd̅ȓSŎ	"�wB��$J�p�ȓ>���v_r�,���]�1������M�Ňɋ]���"���B/���ȓ
Ւ���Z�Z�A�n��
����ȓV��H[ ��J��1SN��:慇ȓ?��`ۇ�Ϝ_k4�1�1$�b5��k�vpx�$D<Y����h�d5�ȓ�h��RM(�X��_�*���ȓdf��ӡ�Y�NH�e�2��p�ȓ{�0"T!}zmд�_�:��K�r��ͬ>@t�w@>"RQ��k��$�fI�)7���A�h0���7lpA
r��H�,��.*����ȓ\t�9ʠ-�<P��ab�ٜS�����G�TT���,S���!��x�6��ȓL��@���M֨�Ъ�B��ȓW���"LW�ʁe��Q��d�ȓ<�ܜQ�K��zH�� D�8
�Q��0S�a���߈3���4�B��Rф�$(��C�P�� �Ƕ}�����V��u8�O�&Vu���4��2}���ȓT{�i�#��@���� �,����󨹘'@םM�� DcF�=8��ȓ*�tas�Aϑ ��4�
�K�ه���k���6*�@��-O'&V��t8ꅩ��E�e��*�D�]�nC�	��f����Jy��GI�'URC��)�h�r�#��{�~�1T�-N�B�	f��RSj��%�FP"A���)˄B�I�BԆ����H�`nh���;I~\B��t�FX��
=SG�l���ekRB�	�X�
Q�̕%��I�k���jC�I�!��)��Q���
�Ú�9�\C䉠T%\ �`�ٟf��챣mX!J�PC�I�����J��n$����<�~C�	;u�麤B<V�;��� C�I.}���!��٠{����A_�|tC�9Z(�t�V�sS���<f��B�I9QX�fN��Y&�:�NQ�\B�	TI"�H�/���v�ȿ�\B�&`����b�ϚR�xL�!2�*B�	%!9�����Җ`�x�v �K��C䉩Mkܔ�d�C�Δx0wdI�;��C�3VsfY�󊉊`�@�jf��=XB䉾U}�{��<B�6IY7�B%E�xC�4I� �q�E��(;ٲti�f�lC�	�WC�pc�%ʍ2`���D��e��B�)� ����C�J��)IdHA�*�v=�%"O���/�p$6j��_�
Y�"O�X��-	F߲-���X�d�@쀆"O^��R�L�G$��Ҧ#�@ԓ�"O(�q4��,0t�3�%�����"Oи�C,ϏGd���z9TG{�<i��R:2���Փ6Q^p"cJQ[�<�#^�]D�t�׎/r��z��a�<��P�"�X�♕L�d��f!�\�<IrjY�-�`�D#�$^j�$�P�<��BU"Ib$xe��pR��DÌO�<	���qw��UO��*�r���`\O�<���[J�xEX&�EH��Y���L�<�6���vT����dZ�ȥʜM�<�օ
}nAҐN�.5Eh��G-NJ�<�&-����Ҭו:`��S�D�<y�cȏWӰ�ca@'[4��g�j�<�UN�u|��b�����b����@h�<���Q�8!l����F[���R�N�<�w� �����R5N#��z�͘_�<�D�Xl�P|�҈0G��q+ϛ\�<�QAE�>�.�A���snt��a��a�<!���/Z`M� l� �pኅEa�<����3|�9�U��G�H��o�u�<� ;r�ji2��H�s�*�K��0T�t�`�Ԅ'�����5[
�9ᆆ9D��s��ë
&��R똩'EP�0V$8D�xj�I��cĂH!L�IRD���3D�dk���.6��%��P�D�*$B&D�H�i�4Y���ҫ/0ޔ�@�7D�t��π)	f`��iһq��]� 6D�()׈����ɐ2K��1W�U���>D�|��ǀ%����Eړ�&����;D�X1a��u3J[ �[(G>��6�:D�<���=g 혗@��
0\�D#D��weI�} D�o�lB+"L)�y��́Pwr��w����S`��yB	�?���h�l���'���y�9.��y�W��
(8P�5a��y2)̠Ow\��e�#t>x���j�0�y�'J������		r���"�y�'��1]�\:�
� g���٣���y­���m�E�_�-���q,��y���d��d8��G� �^��#���y�F+)��q�7n�
H�,݉�?�y�O�Cp�$�ggS�l���y�(��y�iZ0,6�U��)A�a>�ȫH�yRHR�$��Y`�F*X��5�o݉�y�I�T�TQ�R�%�μ��j:�y2B�O�� �͒�J�x����y��@������ l�<ɲ��G0�y�R.L�L�aaʗ�Q��  
B��y�{�����2��yCi���yr ��P��-]�a��8E ��yr�Y%Bg��j�×���*%@�6�yB��3~���Q9����	�2�y��O5���%�R�/��`'G��yBi�7K���#�&$�,i�僋�y��?D�XM#PY<�h43�ܓ�y�Z�. �DJ[]�Ē��Q��y",Ǐl��j��D.�hvÒ5�y���\7�5˖��5+�]�uOZ��y"'�))�Dy�h���&L"����y)Z�qa��"faV;Nth!�߇�y
� dd`�nI0�:��
��3�B�"O��rb# �*aj�7��2�"O\�x�C�^��@� gƊkg��"O�I���6z�����'F��"2"Od�m�9ט��:8N��"O~�:�i��i��b�&)$��j�"O&}�W@̄T�B���S�X0j5�"OBA��W�F7,��Bmĺ('�I!"O��a�A�,�&���%>���"O��K��G]�ր�g�f$z"OR�F�<#z��!�`��lڒD��"O^QZ�Ů;���r���3�0�*�"O��24@.���f�N�A�خH�<a��BN��v�)�:�gWg�<�ɀg�(�Re�#�NB�.�e�<���Ҧ|H�i�\�-�4�+�c�<)"�M@9 m�AI�|�I�o�v�<S���w^�Ce��x�p��CBq�<���.J@�KP �ݡՆSk�<q�¾NV$}ٔ �A�������e�<ir�D�k�# �@i�@R�a�<)�+F���9C��>Y	Ę8e�^�<A��6��҂h��Z�`�"N�U�<����%c�V쑳*�>Hm����P�<�`�ݳ�̜Y�(6*��=�0�AI�<���ցhU�T B�0 p��i�E�<���ȨOVr����J�U'(�
���F�<�cş+��MB���Y�gH�<���o�1)Bϔ6PM�� ԡG�<����.E pY��yI�x 妋@�<a���!�ԳtG�it��v�]r�<�b�*�̥��̇�К��Jv�<��C�)\8�m�3�Ĺd3��C�
�w�<yԎ��\�P�I�+EQA� �]�<Q �]{��٢SgK�P4�V�<!F	�4ClpiA��������R�<�$�R=#��"ƗKk�t��Q�<�bN�u�����)�f����HDI�<9��.y�
����ҕs&$u� h�B�<���&H�!������p�|�<!tiF�]Dʐ��&�/EN�T"y�<ch�"/��Cܭpw��D��}�<1F�Õ9L�2A��'wL��h��}�<� @L�jԢ��)E��w�<10�˹��4�q�ˢ0̢���fUN�<�/Q-52��, "��L@-�Q�<9�)ˍȸ�ڒ Ѐ1O�͒��%D���- x�l�+0k�ULd Ra $D�Ԙ&� Ug~�ڧ�yFZ���i!D���(� )�yǃ��-SV0��4D��F�m�: ����<'����1D����� uf5"g�1V�H�p�<D��j��&"x��c�%R�xp���C�7D�Ȳ"f
$0�D�JA��
T ��!�B4D�`k5�˚<���v��D�����3D� 때X�)N-�`�XN�:2h1D����$��D�
TDL:��/D�:��� Y�����\�P6�3D�`z��g���mo�2�yD*0D�H
v��l� ��)X18�Fd*D�!D�p�$&�a��<�#Ղ)���s�$D����fF/s�:�B����� e�=D� �?[��2Ta��Q��	���9D����(��jr�eS�X����S'6D�� �;CI��C�6��e�׬Z#$��"Ov���T%eN4$i���8���q"OX9�e���YAlIt��0+��;�"O��[�R$PDT�$�PJ7P�Q""O0�r3�G33��da�̈́$g���"Oj�
�	@��<�5\�E$�0 "O�1��+ۺR�,x�jV�kr"O�� `�ɒz̲�zsI��r"O~L�l�6��(C��Q=$8�2"O��BdĚ'4NP�a��)���i�"O^s�[�4�6챒-
7A��E"O,i(�I�����K�A]�9��2�"On�´h��c�^� q��?$��"O\�1�5����e ��_b��3"Oz�
�FF�0����I�2\""O��!-QK��H��oK��l��"O�R JN��r��I�>햤�2"O���m3BB�3U
H>� 9f"O�ƬRl8�1fHŅ2��"O~y:2eQ�V�R��� �:E��"OZ9�>�ܹ)��m	@q�R"OD��e�O�6�V�V�����)�"Ov<
�+�8?��̀�O3��"O~�ð�0֐��G2K3����"O�� �W�8hx'�G�GS��s5"O `��'M�Y̜��^��:�ra"OJ@��y�8
KPɄ9y�"Ox���"j�(�B����"O^C��%�L4Y���	%�pUB'"O��X �޽gZ���J9����"O|]I�L_9vN̅��5	aF��"O��� 0w�(� �H���-zs"O��)�+T.8�IR�/ء��(+�"O�-hs.M9�&qQ���@hh�e"O���u�-}�8E��T�s �Pȷ"Oh�b���2T����b�|�Y�"Oh�x ���S��i:P�X z��DJ�"O����,�TP�	��D�;�޴0�"O�t��0��p FR>Xa���"O�����:�r�D��qOVT�v"O@-�t����������_:.��"O.E��B��K�h�3��0���""O�a��M��5H� L�Ut
t"OJŚFf��I5��ᯄ�

���t"O
����Áq>z�XP;���?�y�
U����L" ��pe��y��
62╲�K�{C��Pǫ�yr��;���O�B(d�L\!��'}ў�Oi���A��2) #O�.U|����HO���	�����7Zj��"Oɫçʍ��djA1YI���"O�a�2cS�0%sI�F^���"O�ؐC�?K�&�їm�
޹�t"O�awkP��Hb�[1R�ؼ�p"O ��A�M'u��t�ԉ*sּ �#"O$�`�DD�.a`t�vF��k�ք�w"O`d�J�']����R@	�2��1�"O�x�� GT)ن���8"t�q"O��	R�Z��5�j}���r�"OJqQ��Ѯ +b����D� A�%�y2�1Bd���JL�δ��iT��y�e�-l��xCa��2?ݸd#��ɣ�yRk�$&�R�1��էF8�zW*ܛ�y�MP��]1���Rz90�焀�y
� �,��#�#M����o9��[�"O2I� � �=8�x##�1����"O�a�C^Kzr�h0�ؠi~ *3"O��q�7I1���Yz�"O�}"diڀoi ��7o�&��"OT���-cp�d��KX�>|��b�"O�I��D���Ij�=�0�u"O<[ք�6���V�2Rj���r"Ova1EN~�L��1'�aPp�8P"O��Sf�<�u"2˔�"���0"Obx�A-t���C�?��E�"Oxe2���,t���V/�r� V"OSQDݵ^���d*�n�Z�@#"OZ�����>R�����
,���Q�"O�<(th��TC숞��p��"O@%����d5�Mb%d�>4��0�"OP�$c�m�ґ鷣6+��@E"O�@�C��ZU@u��7(l@�4"O��a�L�HGTS2B�-S$E�"O�����
a6z0��!��m3"Oڙq�EV'{���ӯ�d�Z\�"OH���nE�'��`�;�ht��"O�Z��	��L r�U,M�&DQ�"O`���*�'��;beߢG��]�R"OB8���M~��bw��j��'��$_W�	�f
��	�̎3w�!��"�1�(�@���g,G o�!�ǄIP���3�.7F,qkJ�z!�
�&�
<��Ț�K")���I�Zr!�DɌ&R�s�"@'�6M���ӼuZ!��7 h�]�F�
"P��@&��98V!�Ռp�́өG.ze�(�W���0T!�DC�;FB�)�A�~n%&��kF!��U�
���1��ȫwj�I���'HM!�d26:l��d�d�`A&�1hS!��2-�ዤ��WQ�T���(7�!�d�5R)�7�� (h���eb{!�DϠ`晙v`�	v�5��K3Nx!�ă�q�:ݰ���YĠ1�A�/?t!�˺^�~4�V"x�����  ~!��
&��u-�d�\�I��C6�!���H,�=)�H��T���BU�(!�Q�n:"�#è��W���@Ё�R^!�䌯LZ���ܘkX ��m&)t!�d�)(�BΎo�V�P.��HO!�ą�*HFU��	D��I%�ɽ`1a��O���A-_4(�������z�"O�̨��a���7�?`H�@"O�L�$ W��Qҁ�<B��"O��p�ET�s�P�s��Y-�h��"O�J`�B�Vs����m��nh(B"OB=��N�C�~]K0�3m����"OzEs/�� 0X����ĵ!��e1�"O�5KWCկ� Ѡ�!�c�S"O�@v̍�ݒ���JT.(��"O�M�FƞKG��ʷg(T�`��"OH2)�	Q�U���W<��2C"O�њ�,��c�:��0P��"O��k��	|�)#���j��"Ol<SW�D�  ��`ŏL�s��$5"O���G�-L���� د+|Z��%"O(0�����E'����(�g�����"O��Z��D0;~\;d(�!Sy $[c"O�X7+�70)0l:Ӥ6 �X��"O� ��J�b��)��d[���̩""O.���`�3{��]�%�9�~�[�"O�
#oC�>	�U�P�3<�|@ؔ"OA�G��:Yg��d�����"O�Q@6)^�MAjt��"�6]�*aq�"O�� Č~��4�a;U���(�"O.|@v�	�U���sBO._��u��"OfHAg�Ԣ0�j8(� �e7~t�"O�p3���3w���c��3F��U*w"O>p"V�O?L,�5p� �*|�hay"O|�� �M�Q���	���<ȡv"OL�(�(P�K��� �(�0]cn�s"OB�J%Y @���@6Aׁ�^]*�"OnE��aQ�Hu.�	��O�B��)��"O����D�_;���VM�0�N�B�"O�0µ�G+MqМ��M>�फ�"OT��ΣS%zS�nH0ێ�P "OxY��M��Zd<xV"O](��T�Ie���������"O\�HbmT�h_���hPv��LY�"OdV�1'���\"aҐ̊�o�B�<F%A&}ϤE�2@B�*�y��S�<I�cݗ	8%�a�4(ж%B!�P�<�5���bI,���#�\�5��$�M�<�c��)�|��!�5`"(�QJU�<Q�a؁?�$u{ŨG)e.,r�.:T�$�f�^�}v�����\�*���"B:D��1��\!u���J�*�Yr�d1��<D��	��� u�̺'ma�pBc0D��c�)Ҡ*���}���:�,D����X� ��軕H�k�^�V�(D�H3�O�,n�a J�8D��S�+D��s���^8r5�S�_����(D����b�?H`d�˒��уS2!�I� ��U쇐mx�ъ���2t�!��	�&���G(��[i�)�!`Fg�!���j�8�X4�X#����'�G|&!��4M2 ��ٔ+��[b�W�'!�J)w�&ҥ���d*�M
0K9!��P� \�t�[�*
-R�I�,!�d/zaʹ���(��)J)M(�!�$��E���a 8�V B�+�!�˖L��0a��]#��#�/�ct!�䔍 ��T�[�c�l=3����Py�
�
H��3@��=��b�iA��y��Y=�N�u��;6<Z'
 �y2bI8;�$�[0ǶF�M�$��y G�6z�h�� T*��8r�P��0?A�� 7\��u�WLXL�NJ�*g�Ik�,HU�<�u�-9�R(`S�S-z�8�Qi�V�<Y@5}�$s7B�|�6TB-�Z�<�FH� OU(�S69^X}["mP�<9�$��-��K̳\*|�` �P�<)��4w����d+q:�����R�<Qe'�&���CA�K :�h�r�N�<���4{e�\��d�l����D�<��F
��� 2�K�3�F)#ea�@�<Q���u�D�R��3C`
R��I�<	�/B��A�!���,j�!I@�<��h��q�ZQ�-C0D�ɠ�Gi�<Q&�wi�d�V�PI*L5�w)J`�<a�.��e��U����Y��`{W'�_�<��/w�=�ƥG�Fbp�B��LS�<I%��U:��p��<i&L-����J�<� Fp�v��
W���w�>:�2䋑"O���kM��H8c�H�N�^��"O~�1�kY5l 0�gJ�"���#T"O0�s�mQ!,�F<��)�%4�H�Q"OZP7\�-˲E:��ͬg����"O8U1!��q�	�W�:/w���"O��c�d�6-V��_e���"O���d?l50���h��B"OF�+������-�I�� G�U
f"O�3�%X�2(0W���2�p �v"O\Ywo��VjH (��[�X5��"O1i�k��Nzh�Fҭ/x�$��"O�l�o2p���"+Uc���E"OzԢ�c[;_&���/v@�(�"OĻ�ˇ*@^<���='��JV"O(}��BS<�D�A"Ɏt���*"O�ܑ���� �4ա���9A���S"O��j`列2�Ό	��ɐ+]bHX�"O2�ۓ��!w.|�4fO%TCT��"O�1h��B<nۖ��%�W�D���"O�Q�]4��jG��-/�`"Oh��DV�OSL�JE�E�Fl\�"OPx�!�Òk�&Uq�� :츥hA"O
	��H�uMr�3��2�t0yS"O~Tba�>]�(��J�7l��ȫF"Ob\[b����ѳ�HF�t���R�"O�y(��C�*�X�'��h�a a"O*��S���}�h��kְ=D��F"OD9jaA�B�ȅӆK(;NP�"O&�Y��ړ:���0(�=Z%�HY�"O�|#h�-2�ВAn��Ipx�q��'3�h"�뒼k���z�A-n�t�N/D�,����0�&
�.������,�*�S�'j ��n݇T@���J-XCɇ�{��ĸ�d@Yh�*��%H�zT�?��05���\3pq��s2`�:�����F��e*�ƳG;�$�ߴ=�ΡQ�'ڹ�ìZj� ��&��'���
�'�P��"��&[��5��HE/b��Y
�'

�K�tY�"f#}*T	�'�1c%j� 욶H'�Pd�'���!�J��TW�rf�J���j�'���4l�v�m���(H��]��'W`��S�7t���8C&J�2�X8��'Wf yG'��P�H�9�*�' �`�"�'�(�r�(��%�d�
!��;�'��z��,C`�꣄�"�r$��'9j��(�j�u[ �O�9!�'���`�dP�l��X���C�	��=��'�������t�FP1/���^�8�'60�� ��yh���i�M����'���7��	��0;h�q�y�)擡8"�Q���>$6	"!�
�#� C�ə.���B�lQ"DO�����2B��B��;
Z�\�$�P�e�pH" lB�I�)��!�"�'��3��C�2l�C䉭p%<8q�F��M)���?k��C�C �h�I�.B��0� ��|9\B䉺-J�ujQ%��>�d��×0tv�B�I&l���I ��*�f�Qw��F�`C�	?R�쑪�AK�r86�ܕ%�JC��\���P��҅AD��"��(��B�Ʉ/ńU�2M�'|݊ �V�2�B�	���DkW#��-)�X���r��C�)� 6�r�.O����d�u��=:�"O@�j��Z�Vf��E�&��e��"O����k��i��J|XI�"OZʑ�5[��|Sq�J�G����"O����J�'!�ܫԭX�flT���"O@� ���1pRZ���l��y��P "O`��� Q�j|���3J�lk6"OJ�j��,A8|d���7�h�"O�S"���K�2e@���(km*���"O���Al]�W���iɡco���"OP��"O6t���"R�,z"Of��	�S�v�!׆׶!%�r�"O� ��o�n�D�ֈ�ZfU��"OȔʗ苨k TX�ƨS6����"O���4k�o0d��ƅ��Hh�3"Ob��'Y�q�:X"�%�J�(h�"O�qu)�&;`�Ke�V��P�"O4�EU����`���]e8�J�"O�M����"&!�8T��QP�I�B�IZ� F�4.O)PpQaA�A�t�%��1�yrJ�em��G�8�~��lL�?Y�fA1	����W���2h)r��j�2`|=aK�?�v�ȓM&���%L_4)8L,+&$Hn",��t�'��M���gE�x���YF{��#$��"ѮY�K��8�����0>�g��\�.h��k~��${��JHa�x�f�,֠�w�̲������ �.�6����:W�@j{�O�8s:�u$�46$\�U�.j��˫ �ֵ�B���/9L�a�n�m�<� N_��]��A8k1\A�S.����9��$	X��Fc=�D���	���i��9~8[�P�J�y�D+I�<Ѷ'��X���ZF%�	�IIo�x�$=�}X$���s��PЦL��&���H���Ѓ\r����ǰ�@�S��/LO������s&�5頧��R0O
<R�P���ɁA�\q 	��+����se�iޚ��|��:S�7w��%¥��b�����$����w��7m�X���-_V(P��؟z�RI��\����F_�P��*�"O\S�(�E�������3���T%@4V�"�tȊ�v>�0-�JUTC՘�D�!HQ���=
�)[�Lk<��V&��iy��d�p�BWLܚT�ar�2*E�t ��v�֍q��$b[����t�r'L=v~�ɸ�o >/�~9�*�?j:x��I>.�v-��ʄ�;`.T1W�_�/�"�HF悚6��]���"��Bgc"�I3k�u�tS�k��OMv1�fM\B���ӓ`$��@����@�5��9���o��Et�;?
B�ӰWj݂��
�%@�QDe���m����ذ;Ѩ�;-$������%U�ժ�Һ�n����ڙi�DqU��-K�Ҡ#��āX,H�󮎆>��%pHɠ?n�A��N
+z���RX�r�JՅl�&��p�� ���a��b�P]��	�dTyrn�@�j��Uo�6��'��r'�)@󩉱6�$`2�K8����I�3�8X��ʎ=�!Y�<���	�ϒvr`I��T�r),��S�S� M0Qg���oZH���ɞ�&P���bH�_�L��䙽"i�'�\ӤY�&`�e���#����!5LJ��3�6� d�Eʞ,&�rw�S�4$������Gx���'<���PMîc�0��*�1�$�c�;�"�Z�A�=�5I�,�n9���H~3̂��y���7��*���m+��"��~r�iرO�42��H6��'mp A���p^�Uqm��ZQ�r��$�tSW�ߗb�����E�*�` BJ�tW��^yr$Sb����næf�>�#H����<�&�'d�0�c�IL$y� �#"����M5S��@�bؽD �PB	=N*�\;�O�=�'�T��BR?b����'^u'����i��%PUqD=*0�s�,�J�HP��|��L���U��jm��P���r�<aǪr�z�+�h�?|��(3��DF|�jw�F:��؋g	��0�Ax$D�j�S�3�Q�;qx������ IW���ʅ�y#�<�ȓiy�Y�'ʪw<,T[S�� � Q����Iv��B��C�1=��@R�i{�I�D�*ʓ����ñp!LM;�'?��,��	�������DR@�gg�6� Xrb�7Pc�U
Z�ʵ�pOM$�T���M�X8�,�I��eN���/�J����b m��aAƴ�T�E%�la�D/�
1�~m�G`�\T�i�O[(�P�ҜF��]k�n		#��k�'Z*�X��6\Zx6D�"N������I�P��I@���dEx5Ҥ��	l��	�-=�'4������k$`�A
�K��q2�h�)=�!�� P�dg_�E�0aJ 'pvl��j>@v�@4!
u�ZR�Ƿ
��t�ɖ#]2e�a�2��1�3y8j����n�����ː,�89ˑHH1Ѩ�yDF�-@��!�S3����Qm�wJٌl�J ��'ףv��Eyb�P
a�G*m�N�ח��*-�i����$���y5�J��yrG��n!^� �IؓJ8Pis����?��40krIG�#l�I7.\�4����Iv麦m�=�ZeA��K�?J
B䉆�J1Ť�n20r��$��C�ɍ(� Ԏ��p��$ۜ&@B�ɿP�(�  ��<<�đ�B�X�C��Y

)�����h0Y��*d̜�
 ��h��?�)�'�}j��`�+L!$W�\9P"Ov�
5F#Z]c����O@�a��.GNH#�I�e���n�B�<��*]6*���臏R�!����yX��Ey¡��X�*�G����cwd��y҇��~�t�j�Dڑ:t�BV��-���hO����ȶ�p���焍_��G"O�@�U�L;�
��R��Mȶ���"O�-J7��9V�u� F\�G�8���"O�(�$ 0��Gް���B4"Ot1��_ HX�M�F�\C��y����lc��?O��r�Q�I�����H��-���!eąeA[[:�d�?U�g@�8�r�@ՈDO~ԑ)�K-D��Xe�&O*$%�6�WB��KT)�<���[ ^G@ i%�0|�!��"`{�4�ō��QlT�#DVX�<i4,��~��mX��O��u#�@Y}�<Q�݅w�����	q��"E~�<����7`i!���Q� �z�&Gy�<1��ޡ=9.�ń�N�s���Q�<CT�n�~�+5'�0��|S��M�<)��U�W
uA�a%3  \)�f�s�<�W)��"R(�R��-X6I&�n�<1'"WPp!CGǒh� ���GMP�<A6�)"����e�"Mz&�0$��t�<Bh׾8�<yB���f'BH���m�<��)?J�h �Ʋ5>�"��Em�<q�����d�F�D�y\)֣o�<Q'n��4�@(΢Z�`��f"�e�<Q�k�!PM��@�,�bEN�g�<�b&�A���� �
hȱZ�LT�<��&D�.�@g
Ǉwd�`��S�<���ԧ~3����S)D렼�BaL�<�Q�F-1�t�ׯ*$G�����J�<��!Lh)*�c�L�DaK�Pw�B�ɛjF� S�o�7{*怋��QE4�B�I;>��� Bƺj��j�"��"�:B�I�[|�mwe
?H��mG5I��C�I�n�ԑ�I9h�����P�(C�	�}n�c�l�.�mq�-�omC��. �ڨ�h��s
�,30�A<C�I3�^���#@�bv`$��� ��B��Pkr�ʕǌ��U8p�P�!�C�>��c�A�%�������C�	�1��`�^*:s\�7�
�\L~C�ɛ-r����O`�)!�@$�C�	}-z���I۰@e�-c�i��S'zC��C@T�@�"�s��	��AȪH4��$&?�Ty@	كB�Fl�ք���!��\�V�sR�ݎ�H,E�ƛ&�!��B���5��$��+} �a�5D�dH��V6�����.�`C2D�8��зW�8aP��Q�>u��-D����]�4Lx�ِo��}A�*D�� �@�b�T��r�`��!~����b"O,h�d�\�_������dh���7"O�M*&/^�ZߤL�v䋸Fl�}��"O9�kA'Yb�ґ�ن�B��S"OL�P�b��=���ȇCDX�x�cB"O����OF�Y)�����{�"O\,1w��H~���U�:}�x�@"OF�)ED+4LX+�U�c��2"O|ل.�CW<��$#\j��"O�q0��{P�&㊐@"��5"O��P)���(x��W�"b�4{Q"O�[�O4h8Yq0�Ɍ@o<���"O6���iR*�a�Vᝃ]x\�$"O���b�;>��9�&L6M<��7"On���	W�p��DW:H��!�"O,��$��6����F+z���"O����s!����[�|�"��'"O������%�V����P,\���"OZ���5�а��k8
F�4+A"O^�	Qm���B�_?,5���p"O��j���+�V�1
��%�y��"OV��h��+����	��Ux�"O�dɧņ��q(9����"OҜk��]�'�@q!���!��U"O@�@j���i�m�3d�
4��"ObQ;�ʔ=���gl�## "��"OpD ���@ ���投�B,&G�!�X�u}bI�EDC��5  H\�kp!�d��E5P��er��2��7�PyƟ&�С�E�թD����y�ʛ6X��=���M�i8 L���Ə�y�_`-X�	���� �l��'����CR�h�H�� ̔#��:�':�q���,1{���ʉ!����
�'�0D�H����٨�g��5�0%0	�'�*�������I��\+3�2m��'�؄��KÿqUt���N!��ɰ�'b�,�o�z�`�/ �����'��b����3�ܤ�'�ļ�,���'�f�kD`��g���i͐�o�H�
�'�@`��FJ���jէ�
p:8u�	�'ۢ�S�Πg�>ʔ��_W��	�'��E81!�=(�0,�C�=d�X�'�u B~\Y��¼�l�+
�'&��01��{��a��0<��!	�'��ŕ)g[q��_�@�a��'NY�q+_�l�:��,(.]8���'�Z��e�z�X�"�з&1�ar�'Lp�p�Q�^���dO=nl}1�'����q�ں�N�2� 6	B�R�'pq�� ��P�V�Qi�J
()��'ϼ)�"$�UR�:���C|li�'h�ZQNϣ%Zz��h��V���ȓ9u��C���&���cK]�-A��ȓLs�B���ԍ{@
هwkvԅȓ-׸���H�c��m۱��n���ȓ3Dq)��`:�u3��$j�͆ȓ,�j��ӈٮ@jŭV���}�ȓ`��寖�{�Huڒ��?�ȅ�{2:,y��W&D��)���X����ȓM]i��V�(s�h4�\�7�
 �ȓ> �����-1���{��%�\��ȓn���3���z�d�El�>>�A��(�� ��7ްx#�K"��S�? 2y�^�EqI��H>Deh�E"O��A��=50�kRo"!�))�"O�����S�ΰ[�n�V9,��g"O���$D�Ik���Ϧ7��y"O�xAKT�oBZ-;1-��[����"O|��$�R�uP�쨵���(��"O�|rfE��c��PQA�O%X�"4Z�"Oz�S�� H���� ��|�L��"O���e�i!B�R �M�sr�}��"OL���˧DB]� �06qʕX"O(����1�6�6���Ju��"O�0K�� AD�Z���Odp�W"O�HI���%Z�
�j���T��"O��9s�g2}����Ol��Q"O.�B2H*pw�\k��ǢBR�:�"OF�n�q��KPIJ�ԃ6"O,�!LS�9��Ԋ��j5@5�u"O��B�9
I�抃�z�Zu�"O�@�ĶcQ�B�o�]6��""O�!��H#���Ã�SO��
�"ON�K7��3�$���4��"O�����[��I�E֡D�"��"O:Ԡ�B��hX��# �O�����"O"��UJP�	^@(���;5���"O�ɷc#/�蝳�bC%:F! b"O� Aa!-.�*�����.��u��"O�I��H�)R �Dq���B��%��"O��8v��)��yya�ɛ+`(��#"Ov<���*<6T�a!�H��B�"O��k�*B�'%2��!�2�~X�"O�M����d�}XBď/q��a�"O���B�T�v����U'�K��i"OHI �-ԅ
��[3�K�`�v���"O�t�_�|�"e�"b� �0�"Ox J��
����b��F(����"Oԕ��KG�G<�=I�hH:�,�Zf"O�-KE ֋xK��@�	ŦK��	�"O�$kc#yɊH�VgU�o{vu�"O�I��WoS� W�F�FH	*O,�
��;j�����Q �
 ��'X̘���_@Rr�	8�!i�'�f����(��D�A�Ϣ�f|p
�'klh;�$Qr�������� 1�'�$�3�O��zH�!��ʁq=���'}��YEO��77ڴ��j�*w^5��'f@#���%"j�H6h������',�s�ǅ=�3�Ǉ(A���'�h�Ӣ%�&�(kefK�d֤�b�'�H(i�FͲ_�( kd��d�pj�'��̱��G� \8@͈�l	�
�'P��e� 7lMe�	Z�
�'�\i@c��	�jT�w�4[Vdp�	�'�y�WoE�Fp����^Yz�'�������H{`p !�1|+0��'��ȱ��(�*Q�##�#r���'������ض)x��S ր~�"���'ή�������Ȩ�� ~b��2	�'�`L��L
�0�zwK�$*�x�'��E��ƞ�g�D�i\5�Z� �'"j��D#��$V�I�G�x����'P��+�h�P��$2�#��d��'a��8D�h�d�cek�"q�dh��'Hh��<t���t(_�v��x�'K蜱�AO����2���I,����� �E�FD۷!y�U��EZ_�Ll""O~X��$z��ҡO̍�0ă`"Ov1ɥ	ʏn�fUj��̛�|س�"O��J�NĐ��G�L?N �!	F"O�������J��'��B-�\h�"Ob��$� 8�� S��p̹��"OXP	�,G� 0��a�K%1tN5"O(x��F�5�"�aN	Lz��s�"O�)��IC%���8a�[�����"O(�;T�S�,���xlUys"Oz$1T��%I/�U��͘�E�2C"O�!`ʈT=p���Ũ3�H���"O`�a!�1i�rqB`Q�D�Ȝ��"Of���"2X�#afyۺ�p"O���!�D_zqD�Z0i����"Oڵ�G`  ����T����� �"O�hpCϵ}���q���4��da�*O��k�	N�ղ�	?{����'prI��M9*�Yx��@\(���'�h��A�8����N��JG0�i�'���� �[Z��a )0����'w�4�ƃ���Za��m̹�Q��'��<����uȖ%(�*����C�'�N��4�E5e���.I�}���"�'�dW�Z%>���1cB�i��{�'�:{`i��&�qȊ�[r:-�'��0FG�/s���6FT.I�T@�'�,��H��^�8Y�=�3�F��y2e�6}�Ƥ�.�\�R(33��y�D9C�~ᘕ囂L��]9�㛈�yN����CآI�'g���y"�
k��f&�(0�4)֏̫�y�l�N9������ $�|��Ь��y��}V:I�k�(펌��Dƾ�yҩ��!�t@+Ԁ֟@4�* /��y2�HV8�)��s�^8���ȴ�y�C�'1���MԺc���o]��yₑQu�={Ή�Pp� �h��y�o�&j}�չG�+U� �Z�ٜ�y��C�;��%0S �r�:����A��y���-Wqȭ��� �l��yR��D��y2+T��HH�PBӤ�ڍZ��נ�y"�L#cҙ!�FίZ�\T�`���y��	6��| C�B�^����7���yb ��[��#͑6V8��'����y�J�V��k&gP�>�B�ذ�@.�y����F��=[
��{<Dh�n��yR.��_8l��iK�ܠ�h��yr��>�+�!kv"�y�y2�v�q��XQNIy�g���y���9D"��\��X�uc'�yR��Y ��RGݳd��%H��yB��'�^��"gN>�E�,�y���bb��KM�8���?�yҋ���z���$-��	�yB��$i0��h�t�~<��N"�0?9��е�:u�bÛ5"����H71������o�'�|Y�����Zh�ɰo�4 �5��oɖ��5��0��	��>q[��OȔӧu�[�S-B���U�|]�P��`ݭO���3�TN�S�O���Ğ�0��S�&��.��l�����I���8E�On�U�G���s���0`n�qQ�@��������'9��ɣ�T=��LR`I�} �L�O𩑴�2�)���<��3
ӎ*q���S�N('����Q�tP�?E�ď�_� �FX =�&������=�u*!�)�g�? \<��el��(�m�	r��S��<@���É8U�|�A��Na6����7qO�Yc�'�)�鋼'�ΌRen�~t��jâH�6�����+���NΝ	���fb�L�5A�'%�~����O�>�2�ț�J9�<�����K�:ir�Y�s���������tL���F;e��qSi�H�܈�?�	6�R���P&$Eh�gH+X��KB�Õ,M�㟒�p��R�*c���W��JG:`��>��H��?�J>���ܠf[�	q	��(Z�0f�"-i�d�K	�㟢}*E�O6Q��e�3�^K'��`@�D�R%�`��O(\��g��n]�B��2��-��$s&`xk�͖u��oL���
_�2��A�p`�<O�F1XwW���'�������H
2@t��GN�{�&��G)�;���N��I�?����\0hR�ԣ`(E�L;�@ـ�CO?�2�^�������$@C�P�)2-����d�_@`X dN�y�p%�O� ���S�~�l���ڇ�	,)��"l�)�~�ζ>Y��xZw��0�51�D�k���U+
2�X����:d:!�_We&!i�ɬ+Q�:ç]�V�!�d�4w���F*�d�t�E��S�!���S��A�6��.D�&
Ȯ;�!�$��l��J֏�z�q�Ҩ��!�D��m�X	�`NY��C'�K.M�!�ѦM��L17��!p�%!��ʊU��T	%&E�0���)7�-h�!��X0A�ݸ�'2���C����!�d�9,o���iQ#s#�	�)j�!��T;;��	 �ͱ�H58��5�!�=S|&�r�M"��,R���-�!򄙓�e��(}���1nݡ�!�䄸ҐȺ�G��*T��NV�{�!�D��t�څ'���uod���n�l�!򄚒ByH��ʎ�uF���%Ծ �!�$ׂm����98��G�q�!�ϟU0ag&��w���֪� 1�!���^�U9�����f��'�!�D��=�KI�5�PC��ƽ!�!�K=4��0���er(!U`.k�!�	=-�hɲq�J�DW��pS�D�1z!��IպDh��ٜC��J��7t!�D1,/0H'
ߗl7�m��Ӷ2^!�$U�i.�b�M�E8
���ʂ�c'!��MlI���ŅI!R4s�'�o6!����H}���P�� ��F.!���Ehle@U�Q�T�HȅC�+9!�](n��8��FH��,���:Z�!�DI�C&�r��(F�`L�$b�3�!�Ĕ
3*��!F���}�p哧��1�!�������?:�8�� �&�!�d�?;��l��ĵ8�~̹���!E�!򤙙M�B� �'X!���s�I�=}�!�d�����h����芷U�!�$G��X���(�btA4�L�g�!�d��6�
�R���&^�Ez%���!��Z9�8�Ts&E�5c�J!�dQ$t��8��	h48:%��Q=!�D_���%��^<�B��1!�D���a���Na���2�̎�!�$�!hx`�A�d�(�z��K�.�!�^�YZ:�#�h����ãt�!�D�']��y�k_Vcf����&G!�$?m��A� ,|LP 2�	�a!�dľ1b���FD2Ja�y���_!�D�#��ŀ��!}�0eC�c��(U!��U�^��e�̃���0��'O!�� R0@eN�+�j�{���0'~݉f"O�cC�Ȟ[�K3ʖ='�,�"OnusuB_(� ��JX #�-{#"O\�����I ����[�w���і"O��#2能(�^���/9)P(+�"O����j�qbR,W�%@T��"O��ӭaz�����V#R�[�"O���Jۧ&L�Ԙ���	/(�YB"O��鱩	#Pc��#���"�9�"Oj�ʇH��$g�yH�i���~\�1"O�1�ҽ���iBy H�3"O�5@�nK-�% ##:T�6�	w"O�A��`)&�Ӣ��.[ళ�"OT����1ng�����I����"O�U���jt�'*�~,Ji#
�'��Xt��5s��{��
��
\!�'`"��T���:(�؊�ƾq��p�'hr�K�ҵ)̝���[&{r6u��A��0q�`L�C8��r&�7a.DY�ȓK�H�fC�H4챕`մ5�E��ltRY��X S��a�V�	�H��@�ȓ|$���64�!&��q����ȓ"!�}*3�� ���g
F�̍�ȓd/����eP�8p�ԠT�ȱ��7�8, wk�#(�fē�\����3�X*�'��k�B|p�*ߗG�xY��@6>���O���{��X�h�m��aR���hQk,����6 j���~��� �T��
�X��+����ȓ[�Nţ�J45̉�F��-y���ȓd�&��#�9}����ѫG&�ԇȓyv	�!� E�n�z1EP'S�f���7��8�B�`Y(a�>2?"��mm2�����QY��C�J/:͇ȓ7��B1A�>�<ĸQ��7t�����O�ȍ�C!��-�T��K8]�A�� �2����_9< � ��+f�Y�ȓ)D��I�E�-�`���U�<K�t�ȓ@ �S$EH&p�b���r�]��g{le�Dϐ�A�ĭ"�E<����ȓJ��b�ȇ$:}��k���:��ȓw��}:P�P�~��l�'�Q�0���6������]�I��H�dJL9N�Z��ȓ/�8��`/H�X�������ȇȓ}#�}{A̅�I^���$�5Y�0�ȓmq:�gH=`�J�Xa��1����ɥ�ܲs��I���3|R�(�h0D������ʀ ; jՉ����Vg!D��ɢ
������ꔚ-��m��3D��Ss��,c9>�1qeR���T`7D��@�ٚd�B0�gI<pbd�2wl!D��.�'e��З��TN�h�a D��rc"N�N��%���v$!w�9D�$X"����R�D�@�2D�(*pF�$u���@���
\��-S�i/D���+�%���Ů�
7�إ��,D�։�"/�`U�w ��c��ѪR-+D���0��WBt�V!��d@ƁIv�*D��;5�*���S �k�zm(D��ó����QCB�T�+lp1I"�$D���_�Ndc!�βgt��� �&D��[R�O�9EnM�P��N�kUK$D���V����(�`�J���&c D�� E�גi�02uK�8DXp�#=D�� �0`G6b����cf�x�l#�"Oh����;^���f�l�F@sp"O�D+f.��d�U �׾-�t`q�"O�i�p Y�lX`����	 ��"O\{V�_��w��	wȞ�ST"O���A�7l�d�;%BI���2"O�بt�7X��a��B�;}�l\��"OD$X`̘v�($��(�$I���v"O�$�M�C������o�rX�3"O4�8�h([G��+c!I+b�H	cR"O������z��a�O�	/t<r�"O�E�W��T��z'%3=a���3"O���@��-e��Á�ңE̐�S"O2�C�"�����z�K)p9Z��
O>7�A>|g,�SBS�"�2Q#ڥf!�I�1y�AWD�*A���b��5�!�$J�r�m
��͹P������ڈ<b!�Dӹs�$��#�$(�I�u��?`!�D\t����勃8Q�	�d�?W!�E&*֘Q��g��Y� �H�Mv�!��Ѕ)�� ��C�_Yn\�talx!���b ��3"Y!D R�9�!��.>-r����l~���O�!�H�k	@љ�� =:� �Oۤ&!�$��N�d��g��N�nhȁ���!���(��P��H�8-�R�d
��'k�|IeĮF��x@R��#J�
�'#��� ѣ4m@\���B8RC����'B8�9ƠK�*Y��� K���1�'SތXR䈷8�ؠ8��A{���
�'m���Όd<����=9���'�b)���<<��1 eM�bꙋ�'��a�r���Bi�HH��z|��'���į`�v�5J�4�Ji��'KFa����'�XPC�8�03�'�B40�K��]y�$���n�e��'�����U�:���D�Id�dA�'�f�T��]
�D�$B50�b��	�'�QY�� 1.,Y���x�|�
�'Snřă�2Xh�"�I�����'�L��rM�w(�y��~t����'�N��V���)3���n�Dљ�'C�-(aW25�8h&�ܨ|Y�u��''�)!Pi
#�����"��G��aP
�'/��	CĞ-nf
@Z�O�4jhz
�'�{���"���%枞_򲰠�'ٸ]bv��z��Y�-��P�}S�'@8��x�p�"�
�<�H���'/d��N��<MR��[�H\�'�����O�%֐p���%-6�H	�'��ajū�?7������@
>�l 	�'Ԍ�3���vP,�	� F�!L���'�Ĥi�"#wJD��%9 �x�'�5�b�<#+���#'đ|�f���'|�`q��Oe���A�
ͩ�'�zYP�D�4*��bA��~� {�'��Z�Kמ9=��H�u�d �'�5�F(��mT�,XeB��<т�'�Q���07��zD��z��8!�'עpI�ϗ�6̽P��̒"O���.�>�����4�����"O��j%G�s��e ��O�\}�"O��1E���E�ؠ2CH�\DέE"O����F/h�"$�/
j@D��"O� �3�Δ
�6|�îIM"�ј�"O�,rb�� ���۔�bd��)�"OzT��D.����L�ZOv���"O�0�b�H�H|���>=da�R"O��Yt�_���+�[��.��"O�p�6E�D���c�^�x��"Of�jW��Ḧe�F`J�+"O����L_��궁�$#��p�"OP�3�n]�=�h���|�W"O�l�6�-@+��r#��5u��$r�"O�Pہ`E�b����h��Q "O��b*��&�0UA4Rt䨽�"O��ãܢz�*�0������"O���k�<861�&�'W� ���"O�p갈Z�� �J�T�.mp'"O>�"eU#LA�};�i���A#w"O�Q�p��'v�<����*Er 4�S"O�Y;��#tHd����'}p��r�"O���+��Q��-�YS�"O�-�PA� s@�#�e�9i�j�"O� 񖱴X�3�ʋ91H�3��
	�y�(X0i p  ��   .  �  �#  �-  �6  �A  �M  MX  _c  �m  �w  ��  	�  v�  ڗ  ܞ  ��  ��  ߻  (�  k�  ��  �  ��  ��  ;�  |�  ��   �  C � �  H �  �& - �3 s: A �G <N �T [ Vb �h �n @u �{ ?� ��  ԗ P�  `� u�	����Zv�B�'ld\�0BHz+��D��g�2T(���OĴ��g���?Y����?�fY$E+���J��"�
ӂ,M�4K�C"I�[�L�pelۦ@�J���.J���[�b���)�8���I��P�82�.s�أF�8g�p!p�̊t�r9�Q�L��Fp{��	��;7b�C���?�3j�L��I�/�=2�q�v��u�V�i3+G%T�b�¨F>�p�
'IFp6��������O��$�O��ܘQf&\8��O(qo�X1� 3����O��n��M*O\�D(8b����O��D8`�ʠ��*$�fd��Bțd����OB���O����O��ە[뎇%i�� د &�!�����*;��0m�b��R[��y���Bw�Dt�'��d�EC�{�a�@��(��rnЙy��I�<яR���	�(�K��dQ��2�Q��C��J�m�^��	c�^��O����O$�	�O�ʧ�y�oK�	Z4�8�e$Q�����'H��?�d�i����O
�	�V�ȶJ�7�g�܂��ݣ?l����Ë/l�JM�GC�<=�ڴFz��6��D���W�~������d��<j<���Ǔ�v�z���'O���#��<[|s�U�~���pӨ l�?�;�OȘ2$�i$JU���ZZ1p�N�k���QR�i�4��D� F�Ł��X+=�H�mZ�M�lq����] �4&����G^�h ܿ0@Fԫ�	�����d�&@���a�IdӪnZ��Ms�e�@�>��\KZJ�!��a�l���lO�Z�eH\�.�ne���T0Zi�1�C X���)�i�7��ڦ���B����Z�F=�H��"Sx諧MƸ.�nsRu s����McS�ԏ]&�rA��v`v�rB�E�?���'��jj��wE�"]�t�s��$�H��i3~���'G��O��F	$����"P2�Ƕt��a�rL��7h�`8PLP<R7�'#(C�'�b�'�j���;E6���}Ӯ��$�Lm��� o�(�5�X9Ll��A�q�D��@'03�
�y��)�[R٤��k*����!I�b�J.�Ɇj��PHX�
���U8�����O��D$�d�O��ģ<��J�hX�%FM�O��I�ئ}Jz�B���?�Rѧ�~��O>i��<ͧ{"r'B��A�e�x*��V���?Y,O*Ѩf�����Ia�'�yw��=^[��eD!�L�Hs�!�?��W樻�+ٔ��5A�$n>[0��/��V����7&�-Q�਀��ט;�~��'�qpc����mA#o��mR��[3�uG&ض!Zy���O����)��xqe�8'�ܘ�ON�""�'�67�}�OJ��["�(9��HR�$��Lc�A3k��D/��G�.�7N�!���S�@'GDnPb���`��o8�MS�fJ�60O�-2�'��Ԛ�斮x���'p�S�T@؟���ϟ$�	ay�'��/'ܕ�7b�� T�ã��2
��"EP"kj�h��R;�~�qrU>���|��'�lu�� �={儬+P�E�to6ăC��{tM�D(ĺ�f�ǃ9�����n9��	�KP��3LeYw��*X�@����1��7m]SyR���?Q�'���|��҇q�@�Ӊ�A���	eB(	)B�'��	՟���OTm#b�0h;���@�u�V��@S�C�4_r��|�O��W�%퉗C
ֱ�6*��j?��K��%�1�O�$�O
ʓ��	}>-��'Ů>������2z-�y9�EԡJ,xK �Wi� ��Ԁ�1�������Z�|�¢���x�1HZ ^ߜ	���Ѳ(��@17�^�X��ak���R8�H�=���(u�Py aR8>`��\0rz��	��M[��Il�uz��J�$��{��Nq���X16�r�'�r�'ex�z��H9���W�P��^`�I>!�i�<7-�<�s��/�Iğ ˖Ɉ�<�Z��Q�~��� !�ڟ���K1���͟,�ɹԆ�%�ޢG��aⷖx�S�H��M���T�X0�db���8L��G~�Lީ=�6Y�Fپ"�l�ٱ"R�o�r�N9P�䤙��.����a�N0#�X�v�F�u,��I��MSB�i<b�\�{o5�bl[�?�ڼ�SAG�i1����,�Iڟ �ᓼW<���Ӫ��� 聱��)�b��E{*��4l�,JNX}ȓe�)[�
�!�8T�(+ݴ��$�4'ā*���Or��|��?a`FM�YD^� �I
v{��Y�f��?���x�v I�ećAn̓�?�/��˧i� q(U# <�����2W���3�O�@���9U�Z���(;<����A�S;�丂��\�ƽ���
D,n�l=*H�I��M�ǟ���iD��$���hO:6yvu��	�*��'d"�|��'Ar����r�ղ���X�I�8�R[��7����͟�n�R��'�&C��C 7��(s���i��[ٴ�?!��?�$+]�B��xJ��?���?	�wˈu�4��>�hE�Q�=�Z�z�+T?i���Z�(}����O0���pLhK<�2m��(�Peh��Br�^\����FU�q�[T�Ĺf͇bEN�	qJ����&n`�5����G�Ι;�����	E�^ͫW�m�xm(�O�(Qt�'Q1���'�ƨD!�r�g ���	$?9��'tb�'K2��>�s�E�h��v/8~"T3��������A��4�?���iV��O�4Y>��f�&�idE%մ�`�T����	�؟��	��	��u��'��6���3�3kY|����Xf�RU{ۖ
}`p҅C	�I�H�e�9<O�̳ƅҦp��x� ��}��-�p)�i��bb�k
x�4�Q�����5�2ړI��@�PB�-���2լW-"<X���/�ϟ���'LI1�@�59f:ЂF���h�ń�n�.� ��4��(����>���'��Cٴ��k�2(Y�i��I�k{�-KW̓`�����'^����=���p� �ʧeR�Lxe�g��I*�=H� �A� �	h��h����Ն���/�
�L<����iY�O��*�Zx���0�&�8��#N0�0J'��d-id�ϔCld1�E�;Ƹ'����ě�"�<�!�����z���氓��z��U��O�y�#ŕl�X2��!L���"�'=�7]�g�h� х /D�Q���_�P�n�iyb%��Q	2d��S��O���1��[s/A/3�JAB!�;+��'�PC��9ȸ��/�!"6p��ʹ��3ʟ��d����m� �P���xQ�0?IR��8ό�	��8e�h(�.?rF�+��![�����"n���b_Th����s�ʴ�'�ְ��k��
*�'����S�0��Jي ��B̟�hO@��iR�U�~���P�P$�'�	=5@ў�I�M�g�i�'��h)3�D�"Ob��Hp��6�m�\�ĺ<1�*ս�z���?�����D��o*n���\-^�rpQ�ݧ#����FHinA��ɚ���3��|*�'��z�)�I?�MT.�ȡ�-	��P��>N��]���.S�XI�q���@yz�jز��iK�B��s�9９S ��Ӗ%���h`��:ƭ{�X�'��Ec���ʟ�'@ȉ�F��A#�u��)B�$`f�j��d+�S�i7B6@�lP�Em ����?(��'��6-Ӧ)%���?a�'@PY�����4���SFT�G0p8E!�}���#��'IR�'�bݽ�I֟ͧH	�"AZ �f���CR�ȸ����*8�1#/L�4�PQF�?�JY��G>�6M1H-/��a2v�|�Ug���hñ�W?VR,���lF��c�,ʓ%~��s�Nҥ��B�n�p[���G������p�'���E��|H��iwa�``���uF>D���V+įX!� �S��S�Y��/�d��)�IJyR,�.J�7��O^��BӦй� ҩ0�p��W��Wq>�d�O�ZW��O����O���4fR \��x�T��aQn���K��77�@`0�
�F�h󍄅5o��A��DH�n#X�5��RE�<� ���)I<5H�Ɣ�$n�1����%U4�it�]D�Yѡ��/�'Ъ��{ś�+�<�3�G�ER(sp��+cq:��Nl�m���O��U�Qꂂ-��l!��ή'���{�8ț�*��~�j@�A�=J�p�$Ws�:6�<A�� ��V�'���R�D�'�|���u�r@�W$w9Ј��'���O?F<օxt	�y���ì��O�����
���S�F���ȧ(L�dt��Uه���F��`d���e�U��HW'��]`u�B�K�!c3%\��pJ\�\����O7�mnH���ʺ?G��r�L D���D�|�"�Ʋ'��y: Ɖ)qpպ�#�S�	���	ӟ$G��OE�>�`��N�2O�����䔉����d�O��'���|R@�)�P�@-҉YY�p�R�
��MK���?��@.��� ��?����?���y'm�s Θ� �Z�<:,Hi�nI�qn�l�	4x�i�!�z����ʋ!	Dq�R�Xqz��� ��M�r c�L�a ��+�O!4|�XH��*G\�K=?q��;@`M�{A�7-�ByrF��?I�'���|򇄇Z�D8�V�("� I����<��O�=��O���L'}��1z��
���S�W���ߴO��'�6��|R�'��	XH)����bڻ(���	���m�}3pEE�H#���O���O���;�?i��?���M��9$!��?"($ � +,.ib���u�}
�N���r�%N����?/.&�Ym�� .��E-E(,�K��.�`D|B��X�89Ɇ!*�
@�qD]�Dir1{��G����?���<񴣎�Bn�]��HN�$<�%��G��y���0��H��d���"S����?�iU�|�jIoZB�d�9 �7�O<��]�t5YK�y8�j�"+��d�<���?1�O�x�g�R�?�c�Ί�j.�]jf�,�p)��K�z��QOH%s��`A�i�'�|c+F�j�6� ڴ<,,R�%��H+�yP0b�%��I�OZ�6N����EU2#��;2l0��2/�p�|<�'�B\�Ҭ�lT4a-N�m���H>���(�G(p�:�� �3!�Ȕ'��Is�����}�B�`eF �OZ0�A�M�5�f)�phئA�'d�6ji����<�.���Āw�|�fIC1<F�큐e_�
����O\��B�<�A� �A�,`��o̪��O^&�	��XQ��|��'W���2�� h�/�21bl]bŃ�$�v�*s��5�(k�G�[!���Mn��
L')E`qzԍ�V�IOR����������i>i v�+W�#�A
�>����*<O�"<��;V�2�0��+A���[���M�'�6���|��B��?�Z	�q��&(�`�i���M���?���A�,�,ԁ�?���?���ywI�(0ѓf�I��i!��� �D!�Q�51r���H�E����T�|rk�AU�qHW��x��� ㇅�0b'b�\����5/��a-�j���[v�L�A4�dX{a��	��ِN=l��rq�'.�I�z����O���6��9.��JSB�>)�\������ȇ�M$��fl�TDʥ�p�ëz=;�OXEz�O�"_�hR$�*/BL�H%�3P��D�W�Ǵ!��ٲڴ�?y���?.OP�'��Aڮh~���5�I�nh���&ʂ>�P���"itz4�Ġ�5o��X*��)����� ��z5�MF��Hh�瞗uSࣗa�/�MS�ɑ0��H��E�2���l���E$�����ˁY�ҹ�q�[0q�PH��M:���$@��mc��D8g�°��fވ1 �1�*����y��Ox�<�<�a�B��b��.{~�0��r�	��M[b�iW�I���tߴ�?y�'�R��C��(IS�Ti����3Ũd������O���v>�d͟�U(�sA(*��!����n+9�G=
��`7A�R����)CQ��c�
$0�8�aFf@�b~j�R���C��Ij�*�$8{<�%��;x@&�K��>QŒ�#�!�I�P���$��]-O��A�>��q&� ��l
՟|���d�)�N�cǘ	_�a��16��=�?)��4�`mڬ+��[���2؈'�ȴsS�ٸ�4��$ˬG��n�͟���]����`'r�B�:l	��		5X4^�jG�D����'�0�"���fʀ��3*O�������h@�,T�?HA�wb�jэMʀ�Bf#?����8,�Խ2G�5E����G�19���B�tݑP �Ӻ�֪�$f��@���V��Bya��E~-�?1�iL�#}:�O׋�M�d�ɱ��i��P��Ǚv�<q��C8�F!fJ�&2�����q�'��}z�,@({i1���UX�!��M��?)��DL:��?���?����yW�SDۥ�;e\N�#�[z�~��
�)o��m5��6}�]ٌ�� ٗ}`���v�$��U�	�8�듮X��cEI>������D����ȺL���R?��n�7o+��*E�RY�%ɀ=H��1�s�O�{��$:?Y���֟���n�'��y�d�߭_[j����&>h!��"O���a��.p�~�:G��]�d Z�P ��4�����<�a΋!,��5����,�X��b�%O��������?��?q�!���O��Dh>�{�Ʉ,Gn�E�z�d�g��d��7���k�T�JVK
Z���ޤ?2P4P���<8�|L0w�Q�eU��0��˅WĜ:�MJw��B��
�P�Qs'�4���O^�Q��'M\%��	�5I�R�b!�Ԓ:�r-4�O�!ȑ�ZqD���	��^�B�"O}� �Υ1Y�\��)�:H(xÑ|B�wӒ�O���,�o�T�'�Zt*V"�h��5[��X�- 8���'5R��cG��'p�IךQ���0�BT�B��BȻXDb�
�/��'�Ĺ�7.�qA��H�;�!�ztr$��;l�x�%MYԪxJ%%�t���Dg�7Fڡ�To[��M�qh΃�O �y �'����i�Tؒ�Ĵ~��!8�D�O���ݙt��&+B3u*4��4�P�!���$�O�0"WAD5l�jQ!c��5�&�s�'�I>!e^���4�?����Ww6�C+P�R�KBlX�M�Z(��D�	~�$�O��N��n�ĝ6g�2�KVe���?�	��ǰ0`䰛�%�r�=	�
!?�O�
O��Jh����a5����OZn1h��Ӟ*��a{GǙ�c�$���OR9���'B�S�(��.��aF�8b�ö4R���b��L�<	��ǃU<���˱p�\���L�'�}w��5�8چ��,<�|�gc����OP��+/��#h�O0�d�Oz�Dj�a�e�̆/����R*N�\��ca �h�V�13DM&<����.�Ē�.��O<y5$�?7�rX
Q�Ŭ{��Q���dcn]J�h�%"����O�,D��M�v���iV�L��1#47�l�+��%n��Y���1���v�'�Z6��O���4��Ovc>˓�?Y5i��f����"A�4�X0�ԋ�����&�S�O�HE�'ėt��rrh�E��D-O.o�1�McL>ͧ��/O2����u�xԋ��M�R_j�6
��<5+���O���O�D��z���O瓇!Ϧ�C�+S�
j��b��B�'#�(3���;&:�0��	�kV���Z��!�,ϣ}��	B mFi����9J�.��牖i�x9VmB�I�̘Q��!ov��*���OB�D*��O�x��L�m��X�G@��r��"O�$PQ�Y�g��PA Z�iѳ�|��e�&�D�<�Bėp.���'M�Z�����K"x�6�_�^O��'Ԉ�Ф�'��2��<���Mj���G��h/��V5}����N -���h�V/lt��F~��K#p���SҤ��3jR�yT�d@���q�V�"��M_̔�UC�$��6��6K��'��;��'��':�Z�X"sܚ��Ģ��Rl"�0�'���@6̈�&&��cA�F���p��xn���&p����l -1�}������2����?�������6C��D4]��x �ƈ_��(qCˉ��$�OJ��/��@P��],k�yyph��h�B���)�p�	>���PV�aG
�X��f~BE�x�T��0�{���E%Xv6E�
�Z�).����y�-�1C�3��	:36��dWR�)�']4X���/�	|��E3�b����ȓa4V ��BW *�\�B�GL=�Er�!ڧ� ��`ƀA�qH/ȷWPV���4�?Q��?��₌`x.����?���?i�w�HH2l�|��Q�%)�#�J�f���X��R�`� ��Rf�2��O����i?�W��}-*��6N*_z���y �T�',ӥ �p�Jt��=T&����"�S�
5���O� 0�k(��zz�1�A#�`���k��Ē`���'���84(P��6�#R�˼Y���'BZ(XS��YQ450�@ʥ(��q-O��Fz�O'�'��Kvc%.�T{  �/Kl(���X�f��"�';��'�r�O���'Y�ɒ�\N�ɁgK�
aI����gD�X$h8�Ahٸ) ��G�7����DKj�'�搂%����&�Y�ƚ_�,�Ӫ ���`bi0�,���	�T#?QM��VL�U'�(H�����N����I��D{Bቄq�������n6�A���8����5�ɱ'�Nxi�K�1zZ]2p(I�D1O��mҟ�'40R-�~���	Q�)H��
*U���*@а���?�B�T��?!����	���u�q�Q�p��Y��rw�͉E�8��Q�����/��k��ȖB˪@�$ܛ�=���P	�����E�j<j�o�(����Lf�!|6��ӟ�'Iv X e����C�$O>'�|RJ>q
�0��,��@�Q[�Q��`��R�n��<���T>U���v����L��U�����ф7�����|y�f�l�6-�O����|�pN��<1��N�@����̛=�P���5�?��/h���ˀM�@}��'�G��&R>їO�|����r��P'LX(,ބx�枟0���թjxb��g�P�_W@�P��+�bc>e�Ac_��顅D�r?��0(?�s�៌�۴|:�>i�'v� ��(GCҶ豗���H0��D�,�� Z"���1���-���H��	��M�e�i91�h�*���cw�ų2��1g�n�Ib�'�R�'���H�9��$C�'�2�'H?��e�T�Z��dpJ�Z0QT�E�EHS.ltq�P��O���#�/I�1�1OL�7�P���H@�J�}^����X��I!�O�{t�V+�1�1O`t�v��tt�Pl�|�;��'�	��P�d�Ob�=���:E�
1Q�%/��J!%���y"k�.Z��� �jW�y D�@�����WU�����'�	�g�&�
�`aL� #�Z�(Հ٫� R)`a<���������
Xw��'�I�~Ō�+#	�������hM�S��H�"����cT?�bQ+E��j�'ĥ�ĈЋ_.��#��v󘗌<�>�S%��QHޱ
�mۨ�d���)�>o��=���d��2�+��W *� ���9�F�
��'$|���˵�>��4)��K���x�Ji!�ď'v������ �HUS�BN�'?�6M%�$�1kMnh�Or��>G1'�	�g�9
B�F*'1r�'�ZAV�'5�����,q�ʹJ��J�?��D��w(��0C�¼ ��M��/]�7Naxba�z>� Fi�M�� ��'c����NZIIf��!�p�F	�	Ót�jL��џL�'���l�/���c�m2���jL>���0=	Ŋٹ�2� �枼v^�kP��]��$��gf���_���ˊfy��_y�b!@b6��O����|R	���?��P�|��]�e�R�50�H��͓.�?��R��𥁬|�|�{n�{�*�,�w�� �S� ���iRI�tW^�'`��  b������w�>Q(
�DM��#�ؙlN���=?	�G�����v�O�����RM_�z�)p͟�f�<�'T|QE$�~s��
���|֌ڏ���n�O�L�Rbٸ����19<�0�M�����I��i�O����O�˓!���9�ǛbڈA��BD+L�<���h�c~YQ��'y�d�g
��Ϙ'x��0��Ö*2�Ղ���U���A]�#��l�Q�'�8&Ƅ���Ϙ'�.��qdU��,��랦@IB�����=M���'9ў�@�!	8yD�P���e���;�E�J�<AE	۪&���Śb�`�s�MCy2((�S��_��Q���4D(�!��+יC�*U�`���Q�`AIܴ�?1���?Y.O1����'��wFL-�T-N1^����뚋A͒!d&Y�_�<Ȓ� 7d�l	E�S�NPjV��c�xea��Ye��P �k	-Q,B�OZQz�YE�I.$�F�����7��9Q�A�x_�|�`��Oh�d�O⟘D���e^��Į�x��h�����yB�Qoa@4T��
_`�a"k΢��u���Vy2$�w�@����s���`����̗�n4Ec�'��I�����џ�*��V�Y������v}�pAO� �Z$��KՏ�H��$�i��D�4oV�<:ӋڛL��1�B��,h�HQ���Qx�@X���(x(	�q� �qADa�	⟔�'�� �`��ZF,��&-e�a�M>��S4^y�6��?�$�VJ ���ن�I�?ie_Z���i$��| T,�ԕ'��r�U����	�O��*��"�@iC�*]	쀘�F��O����� �����z��}K�;������
�tygF�>�̐�a�U~�+��Z� �B�Ǫ�Z92���� ����;���@�p"h]�������O �d.�'�y
� |t@g��b������{�RP"O�) P��Lb�b���r}Q����h���x���h<�a��ۤ���!��'t4uzA�4�Q�L�5�C!V����=��!� D���!��69��:�g��F#�u�$ ?D��Fk��4P�U�ǎ�fX�	:�O=D�����۰	I�&v�Vq�M&D����f�����V���:<J�$D�h����Y8*���h�K .iAg�<Q��\8� �cZ�t��	��@�UTz��$D��p6II�r�|�	aB
�Py0�.D�t�P���z�D���h��l��n.D� I�F�D�R)�!��u\�q��*D��3�	�,���!D�H��UgF.�O���O>�Y L!j�D���!��,�8F"O�� A���4P��O$ �\]�%"O0���K�!��LU�ӑ9��S"O^�Ib+1�pY��#H5
R"O$�3w��j\�@����_����3"O�	jc�E$Z,�<�r�Ve�L��}$�~�2ōF���v*��%��`�r�<�4��kJ
����\*/z�$;r��l�<q�Jۮ!Bdc���I~&{GAT�<���={��ɢ�a@<����&@�h�<!�A�{;@��"P�"���jK�<���}[+�"<z6 ��$N�� ��O?Zw  ;Q�kN\bU���C�g�<����w{N�*�h��z���#�_�<6	�z��� p��Q�� W�<i�	� &��I�W<���C���O�<)@N�/��5s�&\& �=a��Uh<QՌ�!l���4o�D�hy���1 ��*�OnbVK v��yV�Q�VAn��B��.����v̋���J��A��̶R+d��/|c���O�D�<.�|M�4$��ZLz % ��%,"�^�Sf���\%NDy7h�'f�H�#".(�
�j\*��W�o��p�NO��M�TB�K%�bt��^���pJWX��t��d�1tP���G5�d	8c�r�'+1���ӤKߵ`��䁐 ��o�V�q�_����I&!���$'(g(�Б'ϟ4*����`y��S�D5P �1���sKF ��ĝa3�$�O��Ľ|R�X��?��c����6��c����0*���dS�Mx�,�I ,�Yv�|�v$�3��ZF�'YJ�A��&��=D(��U�Ϗ ����C�|���V'm�nh�*ׄjJ.�� 	+��>��&�ƅJ�	����:�w�m�@�D��O���5?%?y�'���ѫ(C����3"JB�`�
�'XN�����J9]&Ř>; =8���i�O�
L
BgY�0[��R���/�v
��'P��'�"���^f���';��'����'l��	RH�R�e�́*j�v(����*�c�T���������#�d�!F�>y�ə/0�x!c�|kyxE��)�NA;�)),�:�X�d$.�O<�s��j�ĝ�S��%S��)NV�K��΍'}�	�R����O��=y�'�P�p�'�8�Dϙ*_�}9
�'�V����Pj��#�Z5N�����qב��蟔�'a������9>3$�^xf����)�k����'���'�b�O�'[�)֮QO�Q�r�$�j���kl���pHЄE��`�
��"��D�e\0 ��5ؖ<ӰJ��k���!�a�%� ��KŨ9���;�U���O��X�'��<s4$]sx���Ed�"C�'rў�E|"�ݚ�*�(��\ _qc���5�yr��o�n)�B��ZfV�ǉ����D����I~ye-;��'�?��O��u�KOF�\��p�&����D$.����?a�R�@��$�y��鳄�?��\�&-?~�D3qZ� �R1��K���1�!G�o�'"�,{��W.�)2G�aX)�t�IAV-�4�q�"��$����
��1�S���	!�MSf��tgҁ����c=E��E"�ظ��$0�OtQ�O�P�����@D�G��X��'��M�x}�SF�' ,0a!�?2j���'@� V�t����O��'f1�4k���?�e�K���+��:V���w�E��?q��#� �mY>K[�Th4�
L�\h�1`��֘O���kʀ,,�ry�����V��H�'�����?o�����F��4�U�4����}j��\�Q�R��~�xRF�<9�Z�|�ߴ.M�)��"� B��N;crX�"�A ��a"O��" Z�Gw���n�.2��i
��ȟ|6-߄paνJ�n	�'V�b	�O�$�O�]�2 ٜn�p�d�O��OJ��?Y����G�ά���BI�M£ᐲu�h�^�If�F�'��]�s��g��
O�.&"ͦO2!��CJ;25���O�,c�(���	kn�0d\�EU����������e�BHX��>�3�$/(ni�COΌ��]������=9�Dk�f�g�	�<��#�%6ȪL�B�<H0Ԩ�fQm�<�q,G�id�+�\!H�� ��ޟ`��4����<�sDʂyd*L�E��'�a�D��M��Y+�����?���?Y��4$��O���x>�*%
��=s�Mj�Ǘ|DV��j� "�8�0B�K�6;�i�D&� [�j�S
ݐ�Q�L0�ʆ�H��Rc��Q��<a�zX%I�-�?s,Xy���*$�<�[�C�Q��(T�O��7∟_�~	��%�c5�
�1����#����cfX�9�}���'pXe�ȓ9��Xb��	X���&�K��>D�'��7-�O�˓?��42ži+��'|�	L0w�� 
O�Pl:����(GGrC0�b�'�r�+AS�]��;g�i>����B¶	ۃ�J`:*9R�(�����N\�V��1
I-f� �p��@|�D��nrB�p�$''����ɉ-�����H�'v�M����fÎ���C�cZ�ч��$����	4Lx86��*�`���	���$� <0�|�q"�	�A��H��Iɟ8�Iǟ��	ޟ��OA�v;���g�8F�{�1ܢ?�v�$8��苕�w���J2X�⟜B6�<��(�?��N]���W8r�t}8�G�j�L
bc�ʦ��	�&��M@n�������SΟ�UR\��V>@d��3�CZ�A�1�4��Ms��^f~���y� -�����k�ԟ�ݏEST�a�g���0���
���P��',���e��Dݑ��Ɵx�S埘ΓR1V$��`��2����ntJ(:FC�ퟤ��:/����	�<�� Uhnz��Ѱ8O���N�kF�e����� 
�0b��O蘣��'/b� %7Z�$n���	ƟL���?̀#��
.@<�r�-²ƈT�gE��?т��ԟ��	�x^n��	��?YF-Mn�;���آI�"L�V	���;BG"]k� �MC�'1Tx:��?)D�@���'��O�0�=+t�!�/�4]>N���e��G��$ڀa��'��]����q�r�8�'�M[b7/�6AB�L�;��y��-/\�tӲ�iC����9 ��'\�Y���~���?I�F*��:we�4O�,�@1�g�F �"����*�6-�ԦE����pz�-I:<�	�9I#��4Ũ��lˤ;���ٴl:������C�?�l����,O�䄍� �H��*T� !�$�C�qL>B�	7����cC�z���1���HV7��O�D�Od���j���'a�[>7�U�en�A\�;^^m��)Jh�f�'�R�'C"�'�2�'#�'����C��J�P�|{�]�p�sݛ��'��	؟������I��x�O��	sƏE�Y�Xs�/_Р�0w�u���D�O���O����O��d�O��'�V���L]*�B$T�X�����O���(}�ҙ ���ZC'�S�� �Dү�M����?)OL˓���~��[�����NIVP	a����O��d�'>)������`�ȃ�̔@��ȓe��uHf-���&E<at��ȓT��Ph���8�yFII a�"p�ȓD�̅�)�ZF�5����V�X�<Yu�B�x�ͨr`бbT�(b�jK�<!��W �8;c�$f���UbMo�'q��' ��'n���j�
�:���-�N�1V1�\7-�O�d�O��D�OF��O����O��DU>��Ȃ�̽B��(ꔪ
CF$mڟ���͟H�Iڟ�	ʟ���ǟ(�I�,��2P�/@�	:����L��4�?A��?����?����?9���?���!^n���ߗD82��N���y��i]��'P��'.��'���'E��'���S�n� �-�:D ��Bbh� �D�O����O"�D�Of��OL�d�O�}R��RЙ���)2����Rɦ���՟���柨��֟ �IƟ8�	�< �#�l4�A�3H;:�6�Bn�4�M{��?)���?Y��?Q���?1��y�l۲�
�ʦ.�"m�EΕA����7.h����O����O��d�O<���O�d�O�QFJ6A��:D��@	@�"O�ͦ��	��������Ο���Ɵ`�	ɟ���n�`>t�IAj�~���I�;�M����?�����I�����֟d�Iǟ@��`J<�ib)J%}���cqd)�>�ݴ�?����?	���?a���?A��?���5M�����,�Y�`T&KPܰX��i^��'�2�'�2�'#�'�R�'$��8W���F_�@��蜪CVp��Ԭ|ӄ��?�)O�"~
DI�y�:��.�1M~�%r��=�MK3��G̓��J~�$�i���M?W�d�HT*��Gl���#Z/�6M�̦��������	�O�T�ŠmӸ扲M��\ �L�����C#T����I/��x�Ԋ-:>0F{�O��D��b�`0���0+atLچ�Z�p�2V��%���4�rQ�<� l�xE�֛-
�	�G+�=��P��@}B�vӔ�oZ�<(��,q�d��x�IPv֒C3"[��3$��}y��;v�5?�'B�朂_w�f�I:s�D��`�t����g���P��'?������<'JYq��O�	bd�鰩�OXeoZ%+���\ޛ��4�ZYjK
@�ݳb /#Fl����O4m��M���]�hE��4���/D,�L�`#$�ug,�(kj��3C�dE�t��Ԩ�hO���<A��T	�zMc��
�St�aC��������]��I;�Is�'�����O{U��g��f+�L2FY�x�۴��=O,#}�u�+��5D��,8�ypf�Ek�"���Ri~B��#'���笜�h�U�O\���w��ݽ����i��k	��SCC��FZLC�ɸA/,�(�E��=�%�sd��R��b��S�/P�֬ST��	$R�	s�Z�2Q8����?O1X%�.<,bQ�R�R�Oe���G�_֐�"�� U����E���4D��h��]�s(�4A�k�@�O VZ)ؑ�Y�=E|p �S��|8@D)��uhs(٘^N9ȑ�Y�8Mh �� ��ͨh�T�[y�Y���9�RP�T��C)��ն���H�")����(�`or��B��r�~�JӋ���D�Q��p@��:1Z�"��BÂ���[&C�Wbpy @���(��S��X�tԚ凔0`�z@@�=U�4��IF�QVK�p����4�d�T��<"a��QǏ�'a�����
C1����[��.:�~��5�="�E)i]�g��#jD�S������%�6��=Զ�V�_')�T bs�����OZ�h�'�5%�����v�a�b(�O����O��d�<I��4;J��'�?�'�����*��'Ұ���-A��z�����?!���?q��>6ƀ��iK��'�O�:���Dh�����ٳ&���C�'n"T���	�~�,��RyЇ����;����3��-�tG�z���'y��8O�b7�OL�$�O���럒��97�8]h���#g+<�����0˓�?����?�L>ͧ��)_�&��a3q�'�ĩcv�#c��H�6�7��O����O������$�O.�$Ҿm���E�5�%���?�
����o��3�	������g�hE+w�P�i�S�IY��M����?�;�hˢY�D�'�4O���E�Y�QbT)�@�/�J��`�'f2V�p`n�M�̟d�	ʟ��G�0^�$��GGvy��PUj�ɟ,�ɸ$]
�zߴ�?���?�R����<�dbT [p4:�(��)�T)�wA�Jy��P��y��'+�'-��'��S=R��rBӭ#H2�pj��.j���� �M����?Y���?� T?)�'
�B�r(�3s��(~D�W�ê*︁Þ'A��'���'5T>%!%Hˁ�MKQ ݨO��)(�oO�5�l+5D@��?I��?Q���?����d�O�u6�"e��#վQ�V�`rI�Ո�pSJ�OV�D�O.��OV�D�O�,*�IWƦ��蟈r�m�+,3(�Y'��8����W�<��ٟ���uy�<�FQ��O�<O|p0�3J�e��ψ�д�'6��'���'^l���o�"�$�O��D��ƨjւ�(*�\d
�S"YX�1�-�O��$�<i��d��'�?��)�2��'>$�Ke酴p)�	1R�]���y��?��A||]�ӻiO�'���O����'V��p�e�$O����,F�F\"Y���*	p�����|���$�?]شkߧ%Fڐ��@�&ǘ]����O|����ɦ�	�����?Y��П��Iݟs�D0Z΁�b�ޅ	ln��w�Q��\ɦA^؟X��ny�Oa�O��.R�^�����O�[c*Yp0�0'/$7��O��d�OޜH�������O����O�����A֑Ii�=|^�,���;�ʓ��$�8,�i>���ܟT��:+� ��� +�&��`ʺ׈���͟�z��C��MS��?����?i�U?��Ö�ñ� �^���[a'F58xQ���cT��A�p�t�I��L������	wy�)�� �q�߅=��
c��5v:P��-��Ot�D!���<)�
�K���P������J�FV)\l��<i���?����Q�M����ӓB,��7`��y�͢���8	sj�O��:�D�<���IZ?1���>�l� �@�<�H��&Uey��'f�'��ɨ1I��K|�2�Z�^��b�%"&���+6�M.�?������фn�qOڹВ�گ&����5��
.ַC�'�R�'2剅M�ġN|���ʕ�I�Y�Vʃf��P�aP�����򄒲j��S���A+'�J!`
g�J����<�sY�[O��^>]�	�?�a*O�PJ'rW&1�f�?1H�$�A�'�剠L"<�}�sJشP�0UL�1W<L�@P��|�歑��M+��?y����c�x��'��aI�\�P���QG�W�v$�9���'��q��������C{�rY�s �;��I�ʕ��Mk���?q��D�Rĕx��'	�:O|�Z�n�c\���n�
?q��������1O����OJ��]5;���I�G�f4(�L�\��d�O��8h�C�	ܟ���v�I�x��XD�W�M&b\{эݑR�f��'�a�y��'�R�'F��d�����J-
?V�S0)X�d����e��#��'��|BS��B�Z����R��ջl�j!˅BN�?#�c��������ny��Y�>1��I޴)s���uV2��s1)�"k�'p2�|bW��@¥��ڦ�@e�ꅇJ�D�sg¬<���?�����C<Jwx%>8ǈ!>�8��#�19p� ����Ir�Iay"����'���Yp�L� �q�ҼE�N0����?1���d ~l��%>!���?�� Vu�!͞!�j0�j�N�h �|"S��K��+�Sꐮ��Lmn�ٶ����Q�Z�(�'M���+q���'�?I��;��	�_-��R���V�8Dٖ�]��D�<i��ZU���O��X�jN�ap2��U=hAUs�tݴH�3�i��'j��O��O���7<E�4]�'uv�� �V������zDx��i�O.�(���0&�����z��jA�Tɦ]������hֱ1I<���?a�'u4�J2CZ3��P)�.�@����(ܘ'a2�'��d�@�á�-!ۚ��`MF��2�'ntj2�)�����$�H@ӏ�)|vе�G�G<�誄��ky"�����'���'d�[��(�&K �D#��/��׋oA�$ۉ}��'��'G剫7��� �E����Y���j�jO&�I��|�Iϟ��'�� @�埾��b�=n����/�88`�p�|��'�'o�I5D��	�V4<�S�C�`��|���n��˓�?����?)/OܸB�kw�Ӈ1����	�%*H�{�bƞ�&�����%���'P���{��Jʠ��� ��xɎ�!cJ���?���?�/OXqs�Or�Sٟ��-9�ճ���##�~0u��O��\$�4�'
����ԟ���aO:T^T(��A؃�����'�!L&\�9�4���O��Ay�i�,֏	"�4�d�V�__���IDy�g_�G��O�>�စ�s-���Y�=����s��P�E`�
�M���?���7�J	T�p�b7��-k�fΝjp���58���3�ɟ0F�ݤR]N���I9g~�X&���M���?1�1��� �xB�'�"�'�V@S��!XԴ�ժN�2H�Q
0��̝<i1Od�$�O���.@LbQe �|!��x`	ϱ
A�d�O�����M�Iȟ��i�	_�0 �F_w^LZ���D���'�^8��y��'���'o�I�m����씱�M(%��kS��	�N.�ē�?�������d�=����2A�rb
���J�.f��aQ���Od���O��C��A��O�t���W_�)"+֏j��X�.OD���O�OFʓWi����U`H�֊ɤ#y��3f)ͷ�p<�'�b�'��\�\� %ۂ�ħ~���V^8l�8��*k�+��?aI>!+O�9 ���'<��0�#{L�j�L	?KR�'A�W�@;c뎝�ħ�?��'_=۔옵���+�M�4[��PI>!*O�2��?U!7��%'��0����3&h!���O:�(�ʜ���i&�ٟP��.��ٔ6kNt��a�T�٠�=�V�HQ5"�S�'D��s��J�pp��#\GJ���z��9��4�?i���?�'#��',2�6f-F�!��ƊO	|��SJ�).K��O>��I�c� h1�W��"���i؃I���!�4�?���?�gH8XǱO��r�D��AA#(�H��cA��0h��B2�ɕ��b����ٟP��8A��h�߭"ɸ�s��ܒ�H��	ɟ,��nJ���'���|R�@P��P�bFT��Ir%U�ɒT�Vb�d�I՟<��IyB�(	��0j��Hi�j�Jwa�:6��/�����%�X�'�,��+׎9|̵�2�L%91��@nS1��'2�'��W�4Y��D�z����b{����IG>3t�I�I�t�Iޟ%��'��'q`�i���9���s�B.��P)O��D�O�d�<q�HIEd�O��!aTi�?תp�V�"���f�'r�|rQ�X��4�I$:���[�똚"&�M{����C���O����<IDHJ!��OR�O�D�ɣ�GX�e���&<�� �|�[���c-�SjS��$��HR�(@%|�xt:c`���X�'��i�a�l�V�'�?��'g�	4<�x
E�R�n�*@�5�Ġ^�H��)���#	�b^���� @fP#t��O,�ER����̟����?i1H<q�5~j	�pꐣ_�z��w����`���?)�
�8�����y��(xD�B!	|�F�'�'sb�P��/�D�O��D���G�N�*鲽I�/�.��e��@>|O����Oz���
uh�����Pd�1� 7.;���Of���E�^�I͟���v�	[@l�;�#�U�L��3HN3W�&F�'?B�'�剣0�U�����jHB�؉Q�x��\�ē�?9��������؀Bu�	'7V��k���h�O>���OH�Ĩ<&O�7vC�t�җ6�����=L���M���d�O0�D4�D7�
hcb�������Y#bV�q�'	r�'��]���M��ħo�����H�9�*�(�c9�ʵ����?���$�Ol�dZ �����"�o*<�ъ�I�d}�7��Or���O*˓U��4�w��D�'��� T4K�k@���l�JD	A��T�p�I���"%.���DĈG�x�:����K� <����/��Y�P�S��M-�8��8��'Y&[�ś�a�2�6�:9�@l���?���LM�����I�
��&�D�UX�Ŋ� b�L�䁫u=�	lZ՟4���������'�� ��qЩJ����Ф���N�I��'�$U����3��`�Dk�15l="�J_E�a�SL�2�M+��?Q�
�U��x��'u22O�0ˠ/(
�x0a�W0`�hB��'��'�A��4�'B��'� }���F�1��t�PhF4`e��j��'R��}`O:���OڒO8#�*��?�,���L�(��"���<i�D�7�?�*O���On����;���fDj�ѱbIF(Vq��$FFa%����ݟ\&����ݟ�3�H3x��c�_�E�l*Ph
�h�.�IYy��'^�'d���CH��2�h�b=[J�ѱgb0DjVU�(��Ɵ�%�,��Ɵ�8'�՟�8'��]К���@)��;��Jhy��'(B�'���4}&j��I|���a l�!�V�cb��z0��#�?���䓙?�nB����DW�$ 2kZ&Lx�3��E����O����<qS�9}��O��wHQFAL�����@���lԚ@�|R�'�B�Ē�y�|R1������+L((jc	� �
�8��'��	�D��|0�4��I�O���\Ay"$�)�/ �&ą@.:%�����?����?)0���<�H>�}��Fמ>�t��'������� �ˍ�M��?����z�x��'|p8"��,t��X�9�b���)�"H63v"�|��)�OD��Ef:;к$b
�.xZ<�8 J��9�	ן����B"^i�M<I���?Q�'�LU�!T�r��44�X�x�����"s���L~2���?A�a�J�I���%1��iTc@%h����?�&�:6�O~��,�$� @��r���z4����G�.˓U����������O2�$�O��>�V����JuM6�3 ��&)8|�0�$��O���.�$�O�����O���u�@&_쩋�jM�`�$[t��O
��?����?!(O����?H�&	n�U
��f/Ҝ��ĺ<!��?�K>)���?Q�#с�?i"���5j�Pf�>5�v��2�Y���O���O~˓3MN�Ԝ��F��C1N1�a�-j�8�3[���'	�'��'��a���'���&-�0�!���?:Ķp� �\�N��6M2&0h�'gؔ
r��2���EH�1�#���sn�	 ���?-�ij���$F0-r��+��n��}�	��$'���O2�o�O����O���dEv}P�Qr&^f�d�!���OF�OX�d�5���T�K����)ȇ$����I�R�Ȩ��'��1�v)�4g\!t���&� �W�$���e'hA�$�0Oje�Eg�3��#�̕>�!)���4��؊�(�U���KY����3ʉ�6���C�Űj��h���ֆW���:�+6�\֊�D�R=��	X�5���s�Ϊ^� ��7�ۘk�D)�,S-6�yr&��Y;�b'�7@��H���,qO��A�#�#jj)�@�K8
�	��#ƇhE�����1*`8!q�ͭt �l#�舉!���:��(2���Т�O��d�O�����F:K� ���Ry*���1,��`��م5?\����ռW4b�( ��˕:���ʷ$At�Oi�`HS�r�IK�LUȩ�}B�S�?���S�u��5;�fK�`�YCp�+y�NB�ɡKƜ�is���yb���7=���Z���D�+�	���X�t��'B�`Y",�SK� !b
ާ@F�f�'�����CI�b�'��i�%�C%�,t��9JQ^�6��)(�S/,"��铫5�u�p�P�����t.�� Sn�=�xDC�	e=nt�@��/E��Ys�-{Z�$i�˞ڔ�F��'6~ദ�l�λ�b�&��r���B�p������'�6M���I89u��F�Y�`�&l[
6 nT��JA����	��?	
�#EB��w�U/;�L��V�9J�zI2B�'�.�Ms%�iA�O[.X���O˛F��]9na�a���3b��d�&@T��d�4��� �O���O���������?�]���`"�W�7ՠ4�e̚���6�z�a�nO9 ��i��	K0W�9#&-�.�M�&�m؟�.��9��k��H��!G��7�12��<�O�z�M�!���8��W
A2�"Ot2g/ŉ5�@Q+ݮ]<q����8��'08�����D�d��;p mS���0G걂�aJ��?a��?i��Q��?������rg�z�gNi���r�D{In�3��+~e�R
��y2`Ж��1�)����]�m@�w��P�Ç�\f�ybg�?Y���M3�� ����V(׌�H�tl�M�'�ay��pe�` ������2�7�y�mL�vg�S�dԗ?HL�p�&�8	l�۟�'�,keh`�����O��'v.�R�iO�9�3M09�>�
�����?���?�α�?�y*��CF8S<�u�E���0�H20ċ���'�ҼЉ���,ҮXN~��T�π+4IwG���'F��1��%�Q?�9U�řC�9rr�H�\,i��&D���OL�N�Ę�A��o�4D�#f%\OĜ�=��Î�@��!G͓^��5�m��R���nzӾ�$�O$�4�������Ox�D�OT6��Zm��p㮑.{�Ȧ͕�gO�i��$��m�q^���2wԟnb>!�'�X�Fׁ@��:��/`z�	�W0=!G![!Cŧ�="��@v���yn�'B0�^
4�Gg��^�� L^�`� ��	
��c��>�S�? ��(t��	*���!d�#y�T<j�"O��!�G.������ȗo�N `��H����P��ydՙ~8�4Z4	ǒ��ț�%���?9b)������?y���?�$��:��OW����h�gS�S�.p�*ݷMY�u+aN�4x�eQ�O^�B��_w��">Y'FʔZ�q7�R�d+��j�Q+G��@P�[�^�$=s6䄧"{�m��
<��i��y�z�O���@T�yؠ�W����qS�i�(�O�|���oz�0P��';ȸeK6'���y)�"̅D#mMt�PI U �A����%��aqe��M+ڴu�#�Lx�.e15��s�l�ˡ�'���'�pqR�'W�9���xƫ>eӴu�reL&P��䂧H��O}� �%�"q+��4�6N��D~�ƴd��	C3��YOn��Շ�2D �D�dÄ(S��q �B�k,C5��uELD##�C�"'�������lZ*�*TH��T�K�T�fV�+�&�������O�⟒�f}�S�ݶbȌ�&N[$"��$�"Oڬ�P��}� ��FC0/Jڹ�f����M����\�9	��o՟��	e��&�?%/
�D�G����`���_T�8B�'.b�'�v���'%1O��OXSbkA���� ��0^�
���DS���N9����!k��P�$�D;Z��TC$�d> ��f+�'���l�{ת �f.�h�X݇ȓh�(���P�W(�4\��
���	*��'�R�x�AC L.�䉱	 !`����g�ϲB l�ן��I��; �FT�Iß��IΦ�[2�ߢWr�y@V�r�*9�a#�[�!=m�5i���i,Z��k�'!���U�v�p�j!a��z��*�%�Dܐ�h�,��2w�����ݠX1�\I���O��ic9���w�q��j�%8�|d{��M8R�(�' 	'�?����$�N>��w{TdHP	�2�^���Q��T����O����ToV��CO�j@4�p�b�.gSqO�EGz�O���i�>�Bt+�!�ν��Ɨ����#���Oy�Am��"ab���O����O�����?���߁�WND�f�B	p�J���U��Ml�Ni�1/R̄�	>n}�����@��d�R@�q��6��K�H���؆L6�����	�dP��NF8N8����
N����IF̟��ܴ?9��''�˟%�|q����HS�psv�ܳi.hB�e����e�U+�Lk�W�*HJ�<Yw[���'�ƽX�vӂ7��VI�LN�m�2ԙ��f�\9�����I�s��5�	���'N��:W��u��r�S-R����3CY>��\��	� B���
&�GT���X`��ga؍�GiZ8Q9p}��b�`x0���TY�_�,xݴ8n=�Ӧ���;j-�I&�~�,5p�R�����>Y��`���Z��y��$��d�L%� b��C���ON#���>/�=�r�R-t��[�"�^��7�%��GI���oɟ���x�$f��Ԑ �lL�x��`���:l�`A�'�b�'�D�Ȑ�'�1O��O�i��Yo�1�$��#>��1�@��r���=�E����,!4a"���K	M��"�Ec��CaD7E�%鲉W_���V9. R2�w!~�(�b��vLd���7��'*:���U>$]QV��Y�Z�K�b���h�o�������S\�|���4�Iæ��1酝s�8�s I�q�E	\ "��0�E�u�	���d�Y�X!1�1x �Us1�N�j�9��(�Ԃ�� ��I�H��		���B7�K�S��8a�h�=C�P��b⛶�<��G��?�1 �V��so��,6r\�$��
X�����?�Gǁ�Ohʌ�Ac�ANY	��]�_X���M��R�-�Jñ��D2�@YtT�m��c�!�)4�'���',"�g���������%�Gʇ�n��(@�&dM�6��� X�U@�z�I�,��x��o^���|	aH�!]�^��L�z���b́�'ᄙR^wun�S��A������Jx��ҁ�9d�h7��cs�H/�Obh��3P03�>_�@mW"OZ��q�ŉ;�,�I�cҮm�j���	!�M#M>��gT�N��6�ia6TS&G:��];҆R�D�j��&�OX��O����.�OH���O�m���K�0�`�`�)e&�@Sꁧ;�+B�3qϺp���4���ˈ��U�e�J5���NhP�G�g�>�bmN�9(l�eF%:`�5	��+�,���I�!R��D�ꦵ��� j��A��M��T�%i银?������O�(��t��7�ܸc`�i�e�
�'��g�U�b� �q`]�^T�`2���%��4��D
�[b�n���`��l�E^&u" {��Z�g��H�ƪΨ:,	��'�B�'�d0��C���6��\��BUMC�p�x�`�����A��̏e�|1R���?i�U)�DݎO��P�7�7	VH��o��j��۸9g�q��I��Lu��-�f�P�}�ɓ���I6h?�p ��@	u���A�"O� E�A&�9���s���q�"�Se�'�➠�'� KNP�;��I���h��E$aq��i&2�'?�O�`L��'���'�&
��� �ɩ:���CX�v�ޙ��ˍ'Zpp ��E�3ONyq�O1��	T��=�@�\�̬�[`��� X8��+8B��y2���3o�@i�m.�g}�Fe��Cfώ�@)Ґ�J6�j�d����(O켥���	7�K�}�!{b�-���sϵR!�$R�J�6-�1��+$'L��`���sDqO��Gzr��>	�4}�^pi�J�!>���KF��PŰeї�'����#b���'��'��ם�����:\8���
�n��'	ͣR�`� �i���8A�Re��5P��'�~�1lU�+wdI�b��u�V��4	X=�#��`/F�
�9��Y 6��7�H�X�����m6	�n�dGi8����h2UA�WEŲoth�`&&�O<�(:ФQI�,�F4m��� �Fyr�}�v�O�9��̇���l�C}��ae��,nx��g^( Xq���?a�^
�*��?	�O?�X�����S0/<�Зb�+o���Xa朶^�a{��$�ē_�dP��@3O+"��"NAj�|Ć퉅]���O?�b��,��|1�����I��̀P�<�'R=z͂�c�j�-�z��ĆP�<���
��9����%?z`%2S \��b�L['?�M#���?A)��L�4�A�*��)���$p���D��o�d�O���˩~��� �|�	#	,� �ta�;����A�� AU�c�����<�SⓁ\� �k"�V=�QH1�ЀJ�Lc��4 �O��G��K� �z ���Ĉ}���sħ��y�M6[d�y�/ԋF�0�q�M_��p=��!+�.ApÉZ�9u�� �Iϙ8ܰ���P��M����?���|b��\��?����?�ܴn0)K�ƭ�(�f녩L����S�'9����<�Eݟ2b>�ʞd3�ӗ��R�"6�^���-@����sM�<As�>���*n����!AT=�D�1�e,�dDp���$�#*}pes�,;M؀�
�s!�䚛e��tZ��E�@E��A� l��?q��i>!�'4�HZ�uf`�7�B?H
P�Ac�Ojm�S�RF�,��O.���OTd���?����Վ	M�Yh�hJ�J��R�e�T� ��' \H
�l�Qk`��/ͼ*5�xP޴jNJ���	1r#�h�"��@@�U�F%F�|�6��T� (�OȨ��;HH���$�S@4x�"O*a��j�(��q@�eP�!<p��Ɉ��'��|��pӶ6MS�Q��SE^�<�zæUS!4����	@����l�	,&T���cC\iU�m�I��m�J�E�t����ϭ(����*<�8�0�eX�:M����2A����D
E����-�P��!kj�z-$m�'��E��,��m��5�Mc���j4���m[�eC��_�r����$�O&㟄���|o�4&������Uh��x�k�b��'� 0�ԃN�*!����ެnW4�hf+�5T=�mm�uy�)Ȅ]�����T�Il�4d�{��@腨כ�b��d�\�,;l@���'�b�'�@�����K����t,,ƨ��-�j�\w� u�&��`���ŀTr5�?!b̃�B��!��-�$h(UG�6��.|�\�2���8B(5) ��\P)Cڔ��O^9�'��~ʄ�X#Cv�(ƏQ�7���	��O�<Y�Z2xwBL`7�ڸr��(i��M?���4����=�#��Væ�� �}��4J1S?�T��Mj�����O��4���F��O��d�OD7��G@��P�ɗ,m�����`|V|{���f���A�G�<4џDb>�O a�7^~di���S��p����*V@��gvE�d�\���D�	v9b�a��7J�1��+!cc���I7�M�U�K?��SP�	�d����ȡQ�Yp�kUwr�B�	�,����&ʍV!v=��R`��'���"�a=��ͦa�4d�L�x��@��E�����*&�?4�.Ge$b���?����?P�����OWa
�I���(+8ThTՁ���M���R;#�����������]��"$
�|���B�D9�7�A�o�����/.��Ju�'�&��D�24�`"��L�U��4��4!P�L�ɸ�M�x�'��x��I�x�����H<NzdG�p?�O�\����5!� �%�< ��I��M�����N�V�i�����k7O�)�9�oX#.�r���'�b�'|����'��=����@@U�8������D&@Z,h�V�$ڨ��d+5C���eΎ_���G~�K?gXL�
D逫�Z���@1��H�-�b�C�`C�޺��EQ'ZYP ړ��&}z�'^V ��9i�6�Y�CN����R`����+I�<,lDy��'�X���ߦb�HB�	@�z�! ��� �\�(GQa�0��ԫ-�����*�Mc�����ڄ_B`un�ӟX��`�� �Eb�4�p�]��q�s�ԩ m1��'��'��!�s��w��R�<�Oo��Ǭk�D����5�^��p�S�>P�O���WH+Ǽ,���0nLf��$蘅S}�ǥK�ZW�ܛ4�����'�$M���O�ƭ{Ӽ��,�i�=Y�v��AJ�
�(���h��(�Fl�?��S���$ѫy���B��6&u.�z��ӒP��zBb6'�J}+S��
�������9�P���c;2�x��?���|�G��	�?����?�ڴ?�2l؃@pI9&�D�s���Q&��`9�tHQ�K�Zf��Iܴ�������O���3M@~��v�ūKЈ3F�X�{~����~ �8+�&� �M�t��W�f���D����yMH�"����-�]G��3+�*�$�צ��)O�U��0�I;���IP���>ip���!򄟭��r���69���"�qO��DzR }��{���5+��0Qt��e�ׄXw�@���ߟ��@ᅽ\LdQ�	��	ϟ��]w2����悋�r�MC�(4�a�@ �ɦ=0�H�SA��ZF�'� p�':B�����"�~]yش-~ @2o�����'<5�Jv薸~�LM�� GB����F�?��i!4OL���O�OzЉs���� �kL�b@p"O =Q��оq�*Yz#�UO�L���	1�Ms�����M�v[�lѦy)�4[����"5A�L�%
��?����?�VÇ��?!�����Y5<4h�L�Ro� (�a�@2l��)��Ό<@s�s��hg��5��8�q&��M�0aE��Ne��/�H���Ä��|Vh["MX�����/�|�➐����O���m�����6c��+f��e�0�ȓWi)d�����%9��̷c�F}R�S�S�\�ag,'}jZ,����"�5���i��'�!�dc���d�O��'rn��!N���z���m�/;V�F����?i���?1�St8	Kb�0�������	eݕ"��`b�hVh�_|�|��4�Ɏ�<�"�LH�CB�)2���zخe�1ˑurMU(mC���Q-�MK�@�jc�0P��ɋը�\qah�Al�� (V.e,��"OP�@m]9��p���Пw(}Ya�'cV�dK5+�cV����l������$�P�-�U�v�i���'��O{D4�S�'���'���� �O��qa�� <!�tp��4�ƐaƯ�@�����7����O�1�*�͓xX�J4lϋF>B�QE�W4��t�ģ��w���eZl�x�a���H*,�wKC����yǃ���Ղ��#c��)w�U&<�l���&�x�Y�0	��?$D1!�c�%J� D�p���^���*��z�z�H�>���HO�	�>���آF&�s�՟Gʔ�N�8J�����-�D��'���'���u�	�	����J�! �\
nMK���%˛e�`� �͏�iG:0h��';N)�2�_�+��"?P����4F8�L� 	�Sq )�ʌ�p<yk(?���B�
�8@8�$S���g�O2m����?�����M{,L���Y-j8d	��T�MQ(���6�2�r���i�Ⅲ4��V_�yFy�a����<�o��\�V�i���ڐ��{�xm�d�U�S�����O����O"t9���O���a>q���N�
~P@ ��C1=��y��دAsX`YĥJ�a��]S�K�*}�\E#���91B�
u(�:�5�I(w�z���(��F��S&��݌$�T���X曖�j�L}�b�|���?	s�O⼀pbw�rq��G�1��u!�"OE�
	�*�* �M�@��h0r�IV�O����������(	�d�XHˡ���e�<���P��M���?�*�XI3��
��L̫MkN�9F�Ͱ�D�O��W�PQ�
�#���J�2}�q �O��Ú"jxxBlD>Y����Κ&'�Ob%�����<R��sŪ(����M�$kr<�Ć(NB�Q���~9` t��'��C:������+z��%>��O�4+
��u�:��'FP�k��4C�%��ߟ"|�'�Jxr�C�7u� ݉�@�ƲY�ד?�qO�E)�R��� �J4%�y��قK���ش�?���?�'bt<y���?����M���)
�b�"�W�!�4 �aP�.ZH�r�0$8� c5O�E�'˘�����&�Vx�@;���2b����vA�1+]�]� RQL��<���>	�.f�L\�7��=��i�'��`L��d�Z1mZ��Y��>���r ��#!�̕HZ��+Յ[�\r��'҂���� $��q����v�z�C�{2m2�l���Ӧ��-_i'���ƀ\�&� P&Nˁ�?�E$�<���?���?!ְ�|�$�O�1n��	�b�׶ma2�!�I�+2]b%��9���r5�'����p� <��#��E�}�&oX�	��x�I�!S_��Xe���u�&�9q�"<q2�ķv��,��E�"*
ZU24��'�Hxk��'�T,�ri|���d�<�����m��t��SF�;Ba\��r���hO�>-#�/ՊTN.p���UU��#�I�22��'�6-�O���O/� 2ˊUݴ�M� ��۵�Ê'\�J�թ(r	;5���<�I��)$���X���|�cJX�xB��B��OLygT�
sTP�5.�RT�$
 �'�Yq��	n�	��.Y2-̦m��R����tWZ����_��'ʛ���&�| Y#��-%2�*!�^J��<������'����5�Zo� ��(����M������	�(�J3�ÔU6����>1-O����@ݦ��	���O� H��O+A�1�dS-S���FK:/���'(2��Y�b�T>��yB4�B�鈯RD���Ƈ��ӱO<M@&�)�	�[�0���	��Q�����(�=*��O�9
"�'qh�~�B�\l��b�">�ܼa�)^\�<1�&
�W��Q���	�lS�HS��X�����{�J�~���A�.�)F�2��o.� $
�ݦ��Iʟ��i>Q ����L����m�X"h�vo�$*U���G ��"�B�O�c��[��hOJ����_$8 ܡa�I
��\�,�f�'7^#}�'��4�� Ġ{�P"�*la��[�U����`��H��I)�r񡱦�R����@�7=�\C�	�8���ᵍ�.7��!eԖh\D�lx������ֳ-^f�i^u�*��φ8�~"���yB�)�i\ :�Lx��e�<A�@�%��rN!��_�L)�1KҿTC��R�)Q��i�1d0�Ofe�% _��\b�#ʹx3�	i"OȂ�잂O�`T�a��>7`D�"O�hr5�٣*��@;���I)
)i"O��`gA����mJ��ޢ0�(�"O�H�C�6��y�k3P��uQ�"O��V)�;����B��]���"O~�
aoX�`��ȃ�dV��+�"Oұ���j�;�圦8N>Q �"O� h�O�73�R���N39P�)�"O|�a� �P�n�X�l0�����"O�Ј&�^&f"�����7����"O~�Z7��$_,�j���;"`�=�6"O񊃪��x� �̫^h��9�"O���^=&`4H�FKC�\�,�u"O�uc���57Z�U3�+^�N5r]�U"O�� ��64�n��@��2F�"O��()A���ҢU$U[TA;�"OF� T$�.b�!��ˆ�q:���#"O$e��N2b �(@�As�N�kS"O|*d�&8Ĭ�����2OT���"O�x*��Q ���Y'a�4�"O�30���D��y�c��r�<�h@"O��k� *>:�!���F-p �b""O2�C��Qb*d1F"V�&xi"O~E�!�)�2@��K�,J����"O1����h����G��w����"O��A N�c���#��5�"�b"O(ܩ3���uj<�D(eL6�B"O����Q����JDJ �
�[ "O�a�U=Mm���� AVn�#"O漒�LD�9j>��B�R�Xi�`�"OBu�r@ٰ&h���a�)
bD0K�"On�q�B2����˾F7��3�"O.�P����!��̓�W�^%8��"O���&�z��Ic�n�1(<U�B"O��'	�4�����l �Y�"O��A5�G62���f!Ø&Jx+"O�8�E'�>K�Pܓf� ~y��"O�a��V��(;�L?�=�"OP1(�`�>�^���K�iK�p��"O�� dʁ9���HD5e�M�6"OD�Z�j3&�l�'� '�@��"O�!	�KB99���@��`�ީ��"O�5J" �=UT�0��'y��S "O� T�𬋝�Ь�Ġ�%80��"OJ�µ� �8W,�Ȑ,LX�8�R�"O8�C�#�/ �ɰ���%�Ph!�"O4�����ci�5p�Lp�����"O����x�f�A2C�>3�N�9�"O8�[��N� �yj����Vp��"O�Ԣv�*P(q��K�57�.�
�"OL�`�S�+
�#�K&{��:�"O���I#�j�(C:y{��S�"O|Б�C�f���1�'W |Q �!�"O�Xd�8p
E���} F)b�"O^��0k�c���)kU:�L�S�"Ofd��L-c{��7K�Ge�)q�"O�ip7��H뮕���-%?��Q�"O�i"K̚2f9�4�F*XD�P"OZ`B[�eS��ѽ 4@��"O��Aפ�x�f��@	�7,� Y�"ORѨ�Aڔ-��ś�);p��@��"O���Q��*;������Pɰ�QC"Oj�#�C� Ԥ��&���Yp"O�����%xI`�#�q��##��M�8➔��Y��c��/o4��ìD:6/nq(Ѕ>D�L3��[�D�d���;RDA���4b��iR�M�]��|�IԈT��)j��ԁB�4q�������<aէ� @�>eڴ��yRe�]Ŷq���ǋ]H��+�y⥐�
#�Y��'Eph!VCݖ�ēN���"LF;.��*vA$ڧW��QY'�� M��L�&�(]�}��*�b�BAc�rπ�x���a���r-ǯ2T1�'%&#�`<�3�d�	*�rФ�6�H,��jՏ���D���E��IY� ?�8�v�ӉRa��C�Y�.��mBp�ɒo8��dƃ8��M�5�Z�b��qy0/
�=[�x"헝he�%C�@>,��x��iCN-���K�R �k5"L<Ch��
�'6T�u&���@���$�(?TJ��r�/ITu.�B���i�ȌE��"	sQ��G�G�h[>)���y2B�+Nb�b@�8~��ݙ�BŠ2.*���f��7��K,D$J��L>)��	;�(��+�o����@�X(<�6l��[s�֋$�Й$��Ph���g��23*~�(1�ʝ��=�j�C�*X�b��AH4��&+�W8�X�0���2@�p���gZ��n���Պ�
6_D�C��2fp.B�	6	q8L�3ꉖh�D)�r�8kV�'�z�z��I
t:�V��t�>)�Ն�(k�d8��#դK�&@D�4D�4(�b	*���R��E=Bi�KR�V V����i?�!��[����'n� :G� ���S�0��b�'+��R�u��p,�	x%ܐ2!C/��i'� e�ƙ��I�e^��nQH���Q���=����DѐI���y�!�����	(W =�0�Ǚ-ʞ%B�F�j9�B�ɻW��m�V�M�5	V�#q�NE��b��3Q���D�´k��S7HX���٬N@	�rJI�r��B�I-w�E��޻�>����	ge�L�R�d�2U�>����Wz��)Æ�|�@��ȓ���#���s @e��e����d���F�H�J�#HUv���J,�b��
�q�Z�q�����q��(�H��2,�*w&��J%��Zr�l��X�����>G��r���(�L���q�t�P)��u8��0k�,���ȓq�v�S���5W�
��w�֠N��]�ȓ6� A9�	��j�v���R03L@��rot)���^1G*���u��'T;�ȓbs�`k��ײmOpTС.�$K����ȓ,����2P�@Dj�ƽl�t(�ȓ\?��S®����� I6O�D	��8���ORd^=
BÔ�Dl책ȓ��@P�b�9���a��[�/XJ}��S�? D�� bLVx�D�/����U"OX%3�Ӽst:�9B�f��(�#"O�Z�E2y](��Rf[�q����"O���T��JY@�+�4�F�p1"O�-{�%R�K��r�Z���I��"O���4LG�TѲ����ǸY���JP"O�	�B��WYD��l�@��M+b"Oj,q�!H�b���K%3r�<�c"O���!Iv��;�{�8uJ�m�<�bl��`�x��W(ڸM����c�n�<!��S(m~:qNޘ��7Oe�<�A�ߧU�X��.�O�:�T �`�<AcǶ��d�Sgt'���d{�<AA�>}���:P`݉3-��
u�<�g ת~]n��&o����!���J�<!�90���̢�1UJ�F�<�!ʏ����4�ӜO-h��T�y�<!�,F�k\�]yp�D'2�d�!e�M�<�Ɣ;>0(��*/J�}XֈE�<����2HyF� +�?6R�����G�<�f∐:T��b��?Z� T�wa�C�<yDM[6Ip�<*�j���MB�	M}�<!�f^o����n��0r��L{�<��Ӽp��l臬�( 
��uK�r�<�a�,���Q�\�E�)�偝q�<iUk��[� �J��� :��92�t�<��/d�� ���^|"��u�<�SM�W�<�ӴE �j�"�d_]�<��䎞�n �BԤ-�<��B��X��%�O�)v
G_f	
�KƗ]p��Zv�'��I)g���#�O��:��,1B�,ThB�	�'�������_V�(�`�'| �>q��鋫�� y���͹�LJ�{��C�	�K"�IwY'4�b��Bɱ$o��	z��h��  ��db��ZE����"O �t�J9T����t�@�d��u��"O*�3�(��Y�Ça�!x�ʐ��"O������J�4uo�j��T��"O�i�0�H$[�JCm��Q��9��"O���S#�<y�vYp�Qp���t"Of\�g� `�r��c&_�/}Ii2"O��0í�Kl%z6�:qe68��"OR-��J������5@����"O�9[�J2G��9�4�- )����"OV� ��._�^�x�ӗI�9���'�����y��	[Ǉ�#f���p��EAj0���2�i
�M��?Fu�q��K�5v�ą�3JxR'/Y4�P!QBb�gŒdEyBl)�S���G'+��2�o@"�B{CCK��y�aݤ>�T:SC]���(z�����M����s�`Hp!��]8PՁ�8��"O`M�S!=*u����\B�"O����ڊ>&�<��蝊 ��9�"O�mu��+�d�3炾��DT"O�X
�l�/q8D�p��� |���*O$�h0*�)f�@5 u.��4Xd��'g��cń��qD���W(����'8xB�M |���(A$$�[�'JTLrsL^���Z�@�o���'pٲda��QR�Ag;Pк
�'O�	
	D�5`p� f A�?El��	�'H���e�k�	C#+�C��D�
�'�]K��~� x��Ύٜ�R�'��Ӳ�W�R'��4�y��QS�<� �����-!��H�u��	#b��"O�(��5<d���%�e�B�i�"O�ٓr��	AU����AW�LC����"O^D�#���*�<5�a�9� X�"ON�)�鋈,�J���jT%�Py�"O��(d�����q���D`>9�W"O�%"�.K�dY��)]�����"OD�s�ߊ��D�Y(�Y��W)�!��ڐxj���EL��Q��S��!��� gZ�H�ڦr[r�a$@̷G"!��jxN�ŋ� �Y���!�䟄-�l����ݩ"��x��_�j�!�Ċ�7<HM����`E!�g� [�!��-y��D�� d�R\/!���"�����ʘo�9ƃ�.D�!�̓\�Ap��2���U��X�!�D�W=��ၭ�R>,ЀYj�!�d�7�8pQCI�8���v`� %<!��HHPա�Of�PIr�S�!�D�*1v$�@�	x?�I��n�+>�!�D��T�Z��&(��,�7�!�D��	��jq�;Y}P��Q�^�Z�!�@����_ ��zr��:6�2C�ɻCx���$�����[�h�!� �Ctx��l���1^��EXq�;>Tr!�7f1D�$J���� ���K�:DA
�N5D�@ ���4Z���(���<_Xtj�/7D�X�DCG�f �!b ��#D��ӳ\ e��C��@�S�3 n"D���p�^�lÜU�J��|�I؅�+D�<`��ёgߖ䡕�I��kp)T��0�?:�;�n^j�e�B"O��c'�)�6�1��#3���*�"O�]p�K�l�.�U�Ѡ_��Zt"O�(�H���qҎ�m�X �!"OhaJ�Ŏg��`� ��kh�!"Ob�VCY����˕�F�q�$�p"O���+��ko� �PM�|��"Ox�V���A�AY�Ċ�2��x��"ON��I��Z"RQ�E)^�� "Oh���F�������IE[���"O��aUBӈ;7��r'�[	&nƠ�"O, `qCM?z��)�Ј��EdP�
"Oz4�eJ��Ҁ�bAHM|����"Of�Є��1nՊ-q�;Rxv�*1"O�a��͗]�@�4j]$�4��6"O�52�E��p��x�fj׌|g����"O�}Pu�� ��I՟&̰�v"Ol��bA�/ks2�0"ǦX�L�*"O@�qT�D�;ڎ�3b��'�\ѡ"OY�c��2�aP��Йi�F�c�"Oh�볇զe�xʁ��~q4��"O8m�5�E�u�Dq' Q13fP=1�"OR������q��b*�(�"Ot!a���	K�=Á�� S�DA0�'�MӁ�;� e17��5Y����!��i����'�� �L������Of��>a�O2a�;$V̚�� (�D}��"#ړLX�=���5A3��3�
����
cI:F��*^����B���ev�($�x���{�SҷĞ7E��� �F��&�[4��4�f��6Kʦ�yRe���K�eF*,3�m8�V��ا�t+�}1�8q�
�?����jw��Or���͎8���b�̉ ���A&�xR��0R�.�Pq���xOx��4ύ�P5|!���h�S�O�"p�.@:W��vbˆJDA��''.a�au�\�+��m��I$��?A��w��yD���v�>���,��>f� /O� �����
W�FtS��J�J�< �[��r�������
A�:�x$ �7h6��S�? ��5�Μ=���hƶ.�@0���d6ʓNfl�	���1�*P��3�Ml����5c�+pi�� �;���â�Y*��� ��
��v���O	c�.��;�(p���ш8�&�� �dT<��x�@�7�4܋B��/l�'z�1�����P֫X�X�`9��;s z`%��)%=�'�ў�鳨���R\�G���'��%�N��~��K�&�59�H��$ɿ0Z�mod��V�Ƶ �,�CU�%��Im���n�J$D�<,c�ep@��?)pqq��&ғ�~$&k�qf29"F��4x����o �!,�2Dv��FH�6#�0�<���a4m1���N���J��bN��''޺wYV��8

"���g��ȋ��M��n����J
�O��4w?N1�ݺK�9�B�9�~=�>1�`^����:�`P$6k.4��li�I
؄x�ǈ]1`�r0k�/D|I�գ�E��9�O�?Mb��� $;�1�'P�������6�B���Qs.y ���
�(O�ĩj�ͯ�Ar�lZ�W�	����ĉ�y�3'��@���<m$��
4k�EA
�<YXwL���I�;#p���"#��-���W�o�
\��G��|�U�?V�a{�K�/0*���Ώ_�:�`�
�� �̊�"�<�
� �O�H�dD�\A�I)� 
�(]�3��OB�c ���ݏbJ�{����7�P��<97���sSP�;�ϭ0��J%��3C�'x�j��Կ:����s���.�U���f
J�%�T�R�WH�'�h�(F��6X��`H��D�"�q��(0L��I2=�B�qAM�;<Q��I8fն�`cd�F@��C�'GE�I ܦm ֋�h�'�8�Jѧ2ώ�ON�PC凸sGHy!/%xr<� ��k�'�N�_b�#��O��z��O��xp-����ȚqN���	���xѵ��$���>��Y��%��m�f=�r��x�{���\q6��$-�?�CH�W����o���8s�!�)A��ɹ ��5c2�ۤ3y^���_�+#�	6�>A�g � ��DMf��L8��*�ē0�u�3�r����]�����؟t�7Ƕ<��g���|�'^�<2Ճ׮.���N�3�a�
��~r�P�4��{C��z��z�hE�f�6�J7�Q���)�`��ĤϦi&0�?��'�m@���~R$��&l6��*Q�U�I��M��ˉ�do��k�n�9(��6eN��6S���p�i�S���𠋕�AN�O$$��I��(�s�4�b�B�R�A
�?"Y�	�tb�
~o@i�$!0�!�M� ,�6�����"lҔ�'B0��޴��T��%
xz]w��,�r�CC�+,qOʠ����5,,P���J�^6a+��|b��U�Z�+ �T
[>ʕz'��xFZ�[�͉���&`7�Y��[q�j"��X�/]��؝�T�O:�z�"�ά{���5�͹
e��<�S�5Ƈ=t���j4DN�I<�L ��T�e}L�B5*tӆ�
3����'Cd����D��wv�j�D��I�����6��Gy��2��Q��#a.�l�U ڏg�}`�iF�@���Z5F��e�E#��u1H<�'�J�����d��n�����g��A�	��E\-M�"t���K�Um"� 8����"%Z�J�<�Y�j��!�~�I"u���[�� �AX�k��L�uP��\c��OT-)��� G�`h�s��
2 "әx"AU�k� ;�.�$��!��M��T�`J��Rhb�4���M��*W�A*��'�l8��m�8u��ɨ��m�X���#I]ֈQS���*�|��R�;��?Y�Ȏ)#N8���� [8�p�m�6>,��1挳�	���s�$��'�O<�0��"a��9���m����Ch�'/�Έ�HT��#�6�YpH�ki�X���-NnIxSJE26�$UY��BI��(OT%aCB�%�*����0��pa �$Y�ӨX�%��/WFp 0D�Q�.���#�IP݄�2�¦5K���1d8H ��_}�\�c��'j�{%�֊U.��}�j�+�D�[vM��>@�q�煔�ē-|z�-�*�����=iS���*ؗGB��"h��В4!T�X�}x�%,�O�iq�աJn��#��
%��|���6`^����~RڨR���w�����w����!Ff�H�ԏ�V$�!ႭY�Z^�da���`��OP���}��cMf�1,ŞD&рa�O�X.��<�Yw��4�aԀt���@�_��� �h�H�/-���p$�܌c�'�~T�P��|Qf֑O� Z~52��D�
��Xp���?�S+�`��t��eW��oyB�'�]டBD�V烰K���پ=kJx3Y�\�'�֕�$nB�(T�}r�Q�#� �K<A5���5aDY��<£@,)�PL3��f=ʓ�yr�����#�α �ME<��,��"��y�\y0��+ [TU�FȒJ��X�#��\���M['���
�r��g�>���/_}��;��I�<��Ĩ?˓�~����;���6��u��B���9.�<�_w�J풎�	Z�M��=�ģ6͐H�F( џD�� �bX��V���A{�z�SLЍE����'��p���W�	�ժ;^@2�C[�엧�􁝕l>`�B���T&����g�	Jy���+p�ΰ������C'��-�'��5B���Ѐ0����G�����N�.P�'��)�3?��E�0W�E*|�P�EB�$ihrA�TL�0�\���&���I����r@�1y�@FE�O&�ƪ��O���W�xz6i�U�Ş�~�Ϛ;6�H3��
ل�fM��n0��<�Zw����&Eܬ~�(ebĊ��D�E���jU������e �AE�'���3\�,�|�6΀b
�-P	� ���e��Nf���^1/���	5�'��(�`��0O���#ݿ�邋���M�d��O7��؄�(��h�i�k�D�f���{�<ܒRj�c��U&�p���56���E�2��7 ���T�^�'���;a,Z�+�z�H�OM��(��$M�SF���ƤתD���Ұa:��?)��w؊�뒴EVЉ ��Os�hK�O��=E���ހq��Ј�7j�<�@�i��<�Zw��D��KP
�ީ{����$�Y���^�$<��2���LC1O��<I���
C�,��0, �T�­2��b��8��Oғo�t0��'S�Q*R��\~$<�"F�<1¬��$�OV����.bxm��eJ��{��D�� l��[�_8;�`��ڶa��'L����qY�!�.�XaAfK�H�@7ʓ�hO��q�<�T�j���"A%}��
!\�.�quFՎ�)Pj�G����6�$lq#��:lи3S���kP�R�V��C��)�'d$X	�D�&�)�f���ȩAB���c!�08�ܘ� �E�v�!�'����&Ȏ�}�����<S���O<9e�����o58y���E�# �fD0U�������b	"	R�n�FQ��L\�#�H�����I]6Q�j���j��A�'F]���O�S�$� 5YD ����>lt��q�x��F6qBC��`�ތ���?khl�c/��ا��Zw�đ��cR5syh;Մ�8,I�bD��&T1�O���� ���"�Ӻ�=�H��I�w:��	��>�\��O���e^x�Sr�y��U( .0���B�J�"���*֬����j�"0Wb�b%�O|��1�O�`Y�����}��iݟ��'� L�ܴ5�F��5��O�<X��/X!܄B�ꔹ�2�W��U���],N��#&�
�~2����D�O���R?mP!�-	���й��i)v,Ж@��X� ࣭�����-����8��x�a��f�V,��@W�?$��`a��?i"f�By�' �yZ���O�5�c�d@h��sK�?���a%.P��DW�������(O�~���&�S����ȓ'%
�r�)�M�g"��O|9+U$}2煓;�Pi&��~B�S�d�-&�^�<a^w��A@Q��4�~�dټ�~?uY\h'LR y��\�V����'��8Ñ|@N��~��>jr�ȃ��~ ($��a(� ���'ڰ��P�20���d�'�AHT?1R��$2F�[��=�i&ng�T�#��@�&b�d9cx�,�gW��ēBF☑��؏	�������Vd��9Y���OVe(`,>�0A6L
t��<�6t��]3V$��O�XJ��K�|l�� ���O��ئ	0���'�<�
�C�A���P �'��x��0�k�
�T�}1ǈ�*R8Ey"��t�K�M�k\VQ���
(��ɒ�N���ܭF���#lO‹Ѡ¢p��aZ�
L��r,8�b�C䖵���i���ɢC�&Q:@fI;;@h𛒇P�L4r�>�@��Ov�H����O�D2ts�e\�����<��'��s�>�%�0����xOP8�v-E�C��#3-����5��?�֝+h��c�Q��刔�����at��3Š@�rD�@(N�<��/�y�����(���ޥ	��Q�k���^��(OQ>Uۦ,�
3�.��"�ΗB�jՒ��]��(O�֝�8��Ḅ��{�
��QC�Z?AĠ� u0"�K���6�"<i��]��(O�i�� ҳ1L�C��ʠ'_�Ͳ �C����C�/`�ʄ�K�:�)��84� �\�g߰��2�ɓoPfH���4'��m;$B͚<T�{�J5��+^��<J�B'��8d�Q�֓O�1�r�9V�|p �I�S�6���
	�i�.�!��%���O.�aQ�'��'�ldҖ��{��ѫE�-�`)���V-I������0<�C���0��)Ǝ�ӂ�7<�=C��a~��5
fh��=ъ�A�,b}���P�@S�}(�C���� h�~�H\�C X�i]>�)��
�v9�*�1Th�l�+U�;���j�]?A�O�<I���f4��B�D�FҜ��R; \,����5.��Pe�'M ����=\���S��+fҝ�SCĘ����	�U��&��|�H�s�דe^�O�D��l�7g�V$@D+���� ��x�ğ:(�i�@�	?���C$�?����J�v�S�O��}��Æ�STpq�2�м�Z�4̗{�l:A7h3
�y��5��?Ộw1F��h��4
ޙ��&ӝi� �i�O�S��4�)�'��C��8h�dk҃�U$l����	��C�b=�⡓��Y/~�V���'A������or���"㌊<�Z�XO<��M�9U��O���V��;&K>}D���'xЊ����;V��I4��|���?+��aaM]=�˓��T?I���0I�DX4�a��육<_��iy���3�}�V��5!&���4�p�K>���I�?�0����/�*�xPϝh�<Qdl�9��ik�H\3��(�f�<����
�Y�G�
�w�8�p��QY�<���*dy� [q
^(Q���SŬLU�<��LM>1��0���-_�ԡ�l�w�<�rJ�$>f$�$�' �EuEY]�<� .��B���d%��A�+��!�G"O.�+AmT�a�\�y�a5Q�FXs�"O@���!�E�d�v@5,�d��V"O�=��E�,��v�Х:�\h �"Olቆ�B�/*�#�OĮ_�(��'44�����t�Q�զ3����'�Z������5���@�b�>7�T��'�|͐�+K%��A�ƍ�b���'��o��($�d����f��X��'A��2�a �*����9jc��P�'rBjQ/%`l�d�;9��hP
�'X�X���ݠJ`>�2��N)aK"�z	�'mX�����,W��
�V�T����'~��!_�.ؒ���e˨��J�'��!��*�JD*����ɿx��� �'���҇?w���P▰;@XP�'<��c�DBjj��ɷ
(,{��	�'��=;��!0�<({�dӓ$�(	�'vdKe�Q��9h�Z��f`�	�'�r鑀�ҰHZ��0�������'2t�CՈ�i�DX�hH$Ct2	�'���෯λK�~�� ��.A?��'O�Ͳd�5�D��`e�0�����'`���B�k����Mqk���'Wy�P�&w2x�s�C-pj�;�'���Ul�*H�r��sF?_
1�'�H9̅�(-n��ּbT�m��'���:��U!Kv�=P�"�J?b���'.>�2���m)	P�L�:�:�'�ΤY%�T�"<����dK�8:D��'���H���*+�P��	H,AF�ų�'<X��݆/8�hצH?a�U�
�'ɐ����ԍ?
�Y���G�2:�r
�'����cS�A,�e$��=�8�	�'�n��#�I��l;�W�8'��K�'f:��D�$H�\�I�o
:,1$H)	�'����I�K����
�u&�Ŋ�'����
� ���R��O>s�j�Q�'��I�f�s��EMC�k�"\#�'ޠY['�']F��)�*�4g):��'���`��K�(��ŭ�0h���H�'�<�� ��#�9��N5Q�Z�'5L���&ʀ�����(1�:4��'��)�D���p|��7�Z�<���k�'b���*�ciN��@b��Z�'�~UC1{��97'��T�@hQ�'�*P�D	��+���U�D����X�'���K)t�,��%T}���'C�)ʣjEv_ܥ�tL����' @b��dŸ���C'iT���'�����oPW.@�S�T9K���'} �q$m�oBT��Ǝsn�x��'��E�q�t�rlN�q~PX�'g� K,�V-`���8e�b5+�'�l��)HY���,Q�.K���Z�<��)ִA�\�`�mF�p��B%Rr�<�2�M��~���<<_�9��ŗk�<у	�D�6����7rW�چ-�i�<��D(mV��J�%E�Y*�I�g�<qA.;m��@��ʗbf�呓��n�<A$еK h1�3����EA�<��#�N.\�󦣒�-&���z�<�E�P$%-pB�cѓ\Ґ�iPQ�<�`�91�p��Ŝ�~/<\��N�<� *l#�mP�-W����O#6<��"Ot��f+I�M�H�(�D�1���T"O8�"� &2󢵀7���Q>�(s"O��H#U�f-��AߎS""D��"O,l+�HV�BJ�xb�Ĳv֭xs"O2|����"3����$궍BC"O�Lx�ƁV�>Y
��«0a�"O����g6ON�u3��H6�����"OЩ����r��͚$F�� �jݙ�"O�z�/��I��q��J�e�In0D��BEOν6�<�C���gr�a�'�8D�8 ��l<0�  �A�TZDk8D�$���3�rR��H�y���2D����BL6l����BB�%|�\��o1D� ��Ɣ�� ���݁y�x!�C%;D���P��`.0	0�E�5� t�%�7D��I�-]��D��M�;*��AQ�)5D�8	��νS��u$B^KȁR%  D����M <@:(&B�Ri���#D�pDмc�iը�-X��Q��a"D���,�/nD,��)J!wr���'�>D�8�[8t�2�#��_���b�;D�8#����?����W<O����&D�<�A�i�D��ł�Z�zF�&D�`�" K�6���) ��8m��l@&�(D�HE |���
_�nPie�<D����اm���B�j���J���o7D� h�b������n�z0�k47D���@��1�~��`_����c4D���?F��Fm��9�\u���'D���π6� ̳�hC�PeXM���#D�(�(�>��ᶨ�J�R��`�%D�d;w/?�:U����<L.��"D�2!F�F0�Q��H-r[��AS?D�`�v%Nf(F���c�3j�a�M=D�d�ūG  ��`��
ƁB�us@�7D�t˔ A�E Z��˃vn�� )1D��6eآ@4��� 8pt �4D�p7�X6>ȘLC �H�7������=D��)]�b p4jQ�Q�.�Z�aP�6D�+p�Y�
m0%L�d�p&�8D�$��l�:VerY ��=s\t�51D�<qQK�	lFl�!$�(I#F�P�#Ó�hO?�C5�Ѕ	�Q��1�F��/�!�/W���!��W�6hÐ �;W!��<v�,(��,��!zFO�l!��,|�ĹJ�+\�RGDG�j!�$���Uy%B��\ݪa�;+�!�d� x5$�퐮P�z����,b�!��0���{u'�o��i��Y/I�!�6	�=뱪�1B�2���m�!�Ӷ�bM�T�<�-Vm�!�K�%��jL�:��X� ���0�!���MȆU���҃��aɥ��F�!���+��CoC7=FxSM�)d�!򤆣<��D׎�U[:E��"�!�D�"L�hR���� e���k�N�!�ӷ?���R�GGKp��"�1a�!�����H:$-�`65��cW�3!��^>t�.��bE�(���r�Úy�!򄕶!kܱx��� 뒰� ���!�$�loh�[�"&D�h�!Gf-�!�E:?��ݢpfF7s�j��<a!򄏹E��$;��_'�ڜ҄���!�� 荰*���T�Θ�a_x���"O慠�@=wkj�P�G����
�"O��P�*c��AC�e��=�"Ot`"�<b�`�E��G�HQU"O�����/���s#�!�B�23"O��g�ӓn��$ 7E��'Ҍ�r�"O��#d�~?��%JP$za�EkP"O@S�Fؘqr<�8C) �wM�-�6"O��˗���6X����*�&laQ"O�};������#��/$����"OZ	�Ԭ �Oʾ@cZ1
V؋tD\q�<�DB���b��Ϣ9A��W�<�!�99�
�)��ߔ>�x�Ș[�<�3�W�v��M�cDI)��0�&T�<Q�c�^T~�r�� �N�<�"�gFL�<A�HڍR�0Y+��ӜQ��L��G@�<��
oL�:��HԀ����w�<�,H�l������I9!\�V&Xv�<)�Ì+"2r(��A)�n!��hGv�<�a���M�Ѻ� |�v���s�<�D�ȂaתӠ�?2&(��u�<�1/C;C��I#R�\ B���I2
�m�<�f�45�-fh�K�ȑ�&�b�<i�N� Ь$�Lɗt����GL[�<� �^
T@T���(�I
���Y�<���T�_�L��p��y��{7/R�<�e%� F ��I�Y*%:%����t�<iC�G�.�*�& %R�Y�%Hz�<��-ݻxCJ�Y�G�a�� &g�k�<I �N,<�1�1��<�|��Ff�<Q�H�$SC�T�fG�7�,�1��M�<�� ��`�P��G&Բ4[��EK�<��Z�D�bm[���},�h��.O�<��fB%Jy�� ��1�X�j�,�t�<���l���K�f8�$�WX�<������`Mƫ`|�;"VU�<ynY�IZ�uI4�ֱz#N�"�P�<���
Y؎L�1��-�)劄v�<���
�ya��χ"}H�班]!򤑾e�x�Q)�|�qæ�&]:!�Dڙ;�츸��)#{
�҄��Z!򄆜+��%��$z�X�"�T�!�C	K �5��gC�� ��a�'4�!�d�;|F�(�� �$9����4O!�$CML>�d���'�N����=!�.W���I*M�$m��e��h!�DB�zI�0��DYR�,�"�bB�pi!�d }�hp02!G%	�H(HS�^>!�$�I����+��J�:m�F�$"!���꒹�V�I2�ҥ�U�g!�ċY�����"@/��$�=dR!�d(u r�C ��#/h��I8!�Ǫ=&������/
Hxqx���' !�d]�0�y���O�,��\��*S�!�d!(��E�fG�J�̹�oϐg!���ʔ{��D:j�0�  IO�R!���(�a@�A1�(ˀB�Gb!���9�<��c�[2
z�����\!��GJ-r�nP;[��a�� <[E!������`bT�5�\��񎐼 �!��"z�v�(~D�!��[?,�!�ٴ�(��5���V0���%�S�<�!�D9�����e*<��#�!�$Q7A~�1*67$�����Y�!�� ��D��Zf�����=U>�[�"OXp5-M�kF����nǪW9��"g"OpTb�m�1"�*@+�m� Hh�i2"O��	(x��@��8`��v"Oj�[�%ɮMIx���5]Ll�"O���$�H�'��CU��3�*��s"Ojpz"^-M�x�@QE�N��"""O���fAN�<dJ��C�2 ���p�"Ob�Rc�Թd�;"��4���"O�h�g�S�FL9v���*�,`"O^4�g�H	K�V�i��s��TCQ"O���5���^�&E��f�1�"O�,���M�A��4�$�+b1�m�"O�p�ݦ���	 #
z���$"Or)�-qE\�sR'���"O�`Ǔ})�@A3gѮP�d�E"O�����Y�-�]B���"O|�e��X���CE�6ox�5"OVq�F$#0PU�B@[/'=2a�#"O�DP��,	�ت�)�$ ���B"OP�CtƜ�J��`��狋Cy"�8"O�0���
�$c��@��Pr��	F"O<Ȫ��/qm��Y#��60$� "O�j4�]PT�j�.:����5"O�mA��#!v�`�bLT���1"O����Y�
]b��AR�H8�w"O +̓iƖ�9c�@��:m��"O|��n\�w'0�V��w*� �"O��&P�HX�9V�Cդ8� "O$8z�⏿T&2�Ha��j��6"O���AcB�o�y�e	8�M��"O��Y���9Y����Υwl���"O�ᦄ�H�4$���ȸ\Otx��"O�܈�5##��Y6O��]1�	x"OЄ"�՝A2�E"@D�9&��bP"Ov�����D�f $n�h��$"OD�B�ʪ�$]	R,P�Hx4"O�B�L7|@�J�mϷQ����"OV�{Q�Հ�T� L�2�t���"OȰ��NT!��,��я^7"�Y�"Oʐ`��U��Y3�`8E0&�{Q"O���Ê�L�hX��DD;/���+"Oz|�Kό.�<rW�޴SU�)��"O>EKw�I.m��pC_�|$Fhh�"O@���F�:6�"�.��)�"O�`�,Ƀ}��х�Ԝr&��k�"O�T������
�b��7z�5� "O����E��
�1"D�"O�}���0=�I�C=O
xqr"O�asU���X�x�x3C��^	29�e"O$���C�vK���"��!�i+�"O��3�P�E�^E&��D��0F"OX�{�� #A�'a�(��i�"ONt	&��s�W/�X��"O�p8f��0@҆����D��4*"O����ry!�h�7V��q"O��%�B'C��AP��/�3"O6dȀ�C<��k��x�z�a�"OX��G�ǪM��9�d� 6�B]qC"O�l��<o����#k[K���k�"O���/l���q$�6A��Hc1"O$I� �F�$R(Q��[w�8�c"O���7�Ζ&�:ب��#TZ�#7"OT�;#/�'$��=��-J�R�(@&"O� �E3!jU�U��e�R^&�EV"O�L�Q�8�8!���O�DM�&*O.��4�ǝiY@0�J�Up��'u��[ �љX*.1 �,Ъ���b
�'�*���iI���k�Dӆ`�(�K�'�`��7��.�8�2W�՘WR(�
�'�lP�G�8E�V�s�F�>&0Ѩ
�'�,��eK��W����V��(
�'��e�ʃ&)���󆁚z�u��'|�J�D��8�$\�R��j��T`�'C2l�Ƈc�ι�\����'�Z�Ӄ�L����*���*=����'����$o�=�Դ[&��4c:iS�'O|8�Fq��ݢ� 92D���
�'����jH`!�Ŋ  !8C
��hOث3��+C�2��/*Y$�j@"O���#&	�R�.[�%ؤ�׀�y¦&%�l��(̋Q]&|� �M��y�iA��ܹfF�?}2��c[�yg�'5���Is-��3�H��ר�yr!��t��B;	�.`A�̟��y"@�U$���ď���Lj��ϣ�0<�����U�zh�#R�
��yG���N�D�O���D{�!��Taޜ#�'�"poZЙ����y���d]~9��Oȵ�m�"/�ybe�<���! ����v��0�ykV�]�p݂�dZ*�@���y2� �9b�*Z+PJP�ٚ�y����DRZ��� ŠQq2�Ĉ��yB��6	ҔD�v�T��z��W9�yRCEW�`�vOW9ڀY���߿�y$G�OU���N�{_L-"J��y�B�&�6$Q ���('��h���y"n�n" P���5`d�(�,�5�y"�ʒ@�L��f�V'�|8���yr�I�k\N ²�a:�[�JR��yB�ȣ]��A4F�P�xI��	>�y� Y�t�t`�cY�'��åF� �y"#U�|]�P���`�U������yrk4yg����M�_h���و�y�(N�-7�����I (���:�y�ۄ�DX���<'�i¦�խ�HO��=�O����� S�.e�"$L_���H�'a�Q���K�y�Q�Y��l�ߴ�(O�~n���� dM_�%bPYG��>��C�Iq�t�3h��]�~�Q�����Y����OD�1��.�d�Ʉ�=qcx&"O�Q�vb� S���g�#��eiћx��'�$@ݺ^!�`�UO�,r\k�'� a��k�7W��c%�V�}��	�':��Qe	�F8,!���H~p1��'��a�Or��is�D=~A��'��U���J�d�9$�
�b�'7���S�ޜT�܅�� Ή"i��'c D���G���@#�P��H�'b$��8S2��ǣ1~5�X
�'4`�э��	�ڄW��&)<$��'rbaW/ڤ)�D�xq�Q��]x�'Z�Q�dF��OE�x�Un׳SR��
�'Ahd�d�^r3rApP��/�P��
�'	��Cv+W�l�u[��[�%��h�	�'�d�E��W$��lX�!�:L�
�'��ЮF s��ڎ�D��
�'`��d.:��ڴ�ʤD݊���� l�0A��vդ����[nLIT"O���	�)|2~9��h�Xr�t"O�� g�߾]���''O)�(f"O ��QOF$h�U'�7�4��"OV����G�~�"0�'���$�z��2�'3�ɗlJ<��$(sʤ�T�٩=��b�P��Ц��Ew(Tw(]�tq�]�r�/D�l�g��9��=��*�7X������/D��q2�7\����M�1X���(�Oh��O$��AF�� �ڈc��Y�h���"O\��S埱"4#�`L!Xdݢ�O��������w*��/4�hA+1va~�Z�,;�O�H�)��`�7�)�	M���O^��P��)�x��%܊����i�<9RhGAjl+��C� 8V�rF�Lp�<�KB�b��%O�,�p9
qb�i�<�EZ�_� ����K�ԩ�\�<�¬M������,#R$���"\��hO�O�r���T�c	č�D+K�,{�E���;$��+��]>}+pة"͏:|ʬ�`�L2���<���hw���6����p����`�<��BߤͱF ϙrh���KH�<�5*H&0�ԁ���*V�;agJC�<Q�.E�|�t�z4B�2Ð�k F?5���)ڧo,��YAȶ��if ŀ'�$�ȓ[&��h"�!&��u{ �W�Q��A�Aq��� S�ɖ�@9�୅�6���I�E�@.�]�p�3U�Q�ȓNq���G�?z\��g�C�:P���ȓ9�(@i��->�\q��B����}�'��ɡ��'(�Fx��	G\<4���'.R����ʣ��M� gٹ"�4i�
�'&�-��gn�PY���ư��'eb�
�!ddX 催���H���.�'��X�'�"mب4'��)�!�ȓ7�<X� ��Y���e�B�����Ij0���N�����ř�tx@@�ȓd��4�]�Y�e�G��'����+�¡/�y���*��}��˓�hO�Sv~�E�t�҅H�,ת'lLpT%�6�y2��,LPt|���0� � Ԇ�y�$A+/4���@�&M]��A��yR�ų�j��f�
t��7��y�`N�B
���,�#y5�az�M����	[���O+N0�ǥ^���q��,pV`$�4�Pxr�]�j�x�/�^rfB�gL;��x-��\=�o�--N��eAO!�dޟqJH�G��TL�h1�T���Ia��+?�I<�O��$�T��dJd
��c��q�����2I�DT[�+Ղ�����-��M��'��T"5픐Eܼ��cH�T�l� ���-��'��q)�d2�"4�ܠAdƭl�4���/�X�Y��$	��IX+/ �ȓ���9�a�3*������۠D�	�ȓ��� �;6�l�:��^�(���'�	H����1�>5��V
6�0��.��}R���'�L�楳�&^�j3b`2:D���%V�,qkfC3��S`�4D��C���;��X`.�@W�0�$�>a�a�P#�<�S�ˀ&lgv���A��Z0��"�<������~����J���ϐU*�r�j�F꘨�ȓ2j`����"<g�
s�]>��%��h���i��l	����3}�H��S�? �p*1��]7�MFfO��0Ҳ"O������^<�L�t��>U��"'"O�Y	�&dȱJ����"O8y.F+'"�,��	�<���"O�сUS�V�"1 ��A ��`�"OR �6��l
`�Ggצ���"O���7	���<!'��>;�1Z�"O�����SF:%��t��r"OR8H�$X��ɒZ�p�a�"O��ȅ'�Y6H#sLژ����"O��õ��##���Re�,Qά  �"O>,�% #;��"�7Y�xi��"O�D{�lB=1�48E(�({<9XC"O�4����f���\���{�"O´;w��*F���S&�gt�-�t"Or�sV.��iʈ�HPm�-	s�ةb"O�}CD�j�I�H�d2mM4U!���;%f�#"�y��!3�L�!�D�9�"-F�*���k"�G�!���"���Zs�X)u�EbЋN�Z�!�Ď85� cR+[�s��[BI�T�!�䆺^N���F�+fB؊�g
:0�!��H�T=B��g��<|�su�<%x!�$�@Ia7�͒ �ݲ%�F
!�$�}���׋�66�pK�=U !�D1F�̓�e��d�t�L� �!��ָM|�If�3O��Ȑ�)��]�!�$V!I^�M�ѮǛ}@�8i�.X�!�:|8HB��"@L�p��]�H�!�D�GX������/��'F+�!�d�5"#,�
BPY�b���&v�!��Hh��Ԡq��#Z!h�!���	���ifmG	E��1�RhS�f]!�č�7 ������m��p�"P?�!�
�l� �x��N�@���'��!�d>h�^X��kԘw����F�OL!򄍐ʎ) VY��a�& 
z�!�ְ)w�4�6��!|�T�!0�5�!��)s��y��%h���I$kE��!�S�Pi~8P@�|�T��d^�y�!�C�Z?��q�枕w،����
:�!�Dɮ Ӱ�Y���`ڊx3�	�)�!���#���X�D[� ��gJ�z�!�D��G��驵��H�.�8��@�!򤔶A��D������-Ƞ-��Py��*o.���DKA�H� �8����yr�Ƭ_��1�$IE�1��8!�C�yI�bpA�F���`������y%4.�nA�r„k�JM[�h_��yrf�\�"x��J� \��Q��5�yb���]3d���F�0N)���`k���y��A�Y���k�e���PjW��y�̚Z�������z<����y2D�@�ji��%P�a�Fl�0()�yҧ��3��*���6Y|�@����y�h gIjC`�M�=��� q���y��^+,v���a�>M��0��S��y��_�P&&�	��[�@��W�umhB�I|��4�f��0W=0�bE-�A��C�+f� �h��x*�j5!A,@ݶC��)�f�0�М8��D8v��8�C��v�&����a�uR�4G�C�I�37p$�b��@end�B.٫5�\C�	*F,&�F��+5@4��I�m�C�)� ��	f� �&g<1!��3�^��&"O�dvb��d�>�K�ٱp����"Om!�:�9��,!
|^x��"O��A��� 7PMH,�LX��[�"O�4��eV�[��s��Y�XMP|�P"OP0R2b$L�N��2��BX�2�"Ou���;CܪD�s�D%1"d�85"O��#��;/��Q���u��;��=D��#D�˙N|��ˑ^��\�Ģ&D�<�v�]� � 
QL[�u-^H:D $D�8�% �-��qbh�et�Q�n"D�D��ȳD��T����
W4�����;D�Ƞs�U��Q��n�nl�[�O:D��a���8N=ۖ��C��t[�8D����ʷI޼P����%n ��BE� D�4�	�7p�����N��h�J'D3D�����c-I�5�(v���K0D��h"�]��c�W�.��3�*D����N�x�$�#�&���o)D��X��^�@I
A9R5�5�(D���$��Y���V�H%"�B���,D�T� MȂ&0l<��j��]s@;�4D�Hi��л����]��A7D����nP-��D*d,P�C{�p�e�6D�ԻPH3i
��1I2n�lH�M6D��F턜'��aIjH?~Ѡ8y�/D�H*J2n5���EtTyZ�)D����*�����@�(N��TJ3d*D�D{bN�Q�r�*G-@���!(D�4��ٶ`��(���"V������3D��`@kNK6210T�B�x�����d2D��A��1�$Y��_$,�R��!6D����Y`��24�^%q���0D�t�eHʴrh[dC	J@��1D�آզ
�<	�	�\�9�: yp�,D���&�ߜ2�8�zv�^��$H���7D�|1�썑^�Xu�am*�`!r��"D�����ܥ "ڙ�E�U,.�⑺��;D�H�P阆7���B�F�9e�����7D���2�C2fj\g	ԶR���{��/D��(FBY�p��*T��u��I�3D�4H eυg�"��G$N�Y[�)0D��x�o�;v4���G%��k�4)�J.D��"�P�Z����#'�����-D�D"��K6y�lt��i[:lz�(D� R�&��DS����;I���'D��@3�1�(�j%i�9$�np���%D�0�fa�:dXA3+�I�f�9�%D�@���A/�DYH�n� 7.�
$D����ƌ-.��X�%��07%手��$D��%���mG���1��3,�~PJ�"D�,1WMN8^&-�����I�8(cQ?D����HU^;jؙ�+F�gd�۵�1D����a�x�fq��%��-6iIr�;D��q���Y������2���n>D���e�B{�M�2��~��vh0D��jf�A,[�:�h�k�4�<
�	,D���% 3]��q�$�g/R���@*D��	���9Rtih��[l pJ��'D�LP�+͸���13��.{Ԉ��$$D��q�e�_�|EH%'a��� qd-D�4��d�P�bU{� �*İ��rL(D�xs��}2QҒ뒶<�Д�`N%D�p85����y��̑�{� e )D�� ��A�_A�f\�A�)yG*�"Of (C�L�Ł4b[=a�0��"Oґ��j+|�H�r7�Սa-�@"O2)��Ē�E����1�A�I>B�"ONa����r�A�[�~��"O� )��Ɩ�AAA,Ĥ�;b"O
�:lŉ=LL�G��}��͑�"O�IS�g��Ja�(�(]$GUd�B"O  ��a��+�a�fB;{�̆�~�
M���Q�o[\�"%%�"i�`���P�<#`�I.T���j����n-.���D���0ۗ{hzYz4 ��~$��!��i#�qN��I0�EM,��-�lDS���3!.��F�ݼe�|̆ȓS�XQ�i#;l��H� G�̄ȓv��
�?#(�����qڎц�n��@�d�������0oɘمȓu�����#[��;$[�/�4��z���K8$98E�sLA"J�ZM�ȓ���@6�<7��T{���%���K��z �����4��D܄�#� i�Jl�� �Q��5��^�ČS�C�U���#`�:����ȓB]����a¸=�pca/ͽ�,ԇȓw�,����U`�E��FȡYCH���}4�=��o�4�p񪲁�\k��ȓ �R4(G�˃y��@�w"D?����ȓ y2���I�{H�����͇WOD����4��f#��Xa��Ŷ`�ȓ%���Sfh�I,�AIu�ai֩��j��YA�捰b��y�@��o��	�ȓ%ҩ[sm��F��3��9:�J��ȓ;l*)c�.�:d��Q��2d���q����Q�,���y0Ŗ�
��������`�F�9هb��F����W�<����]��8���ie/�`��oV�:V�- ���v·�7�p��o��A Q+�H��r-Sc�����4 P�|�ev�(_j0��FJ~xx�ô�&(k�腐rJ�̆�2*NIp!�P�\C���G��J�F���%z��*��M"^�Z���m7V��
Z��K���>�5IG��5ޒl�ȓa���k�&�4oӦ���	@�o�Y�ȓ=��d �b��<_��`��܅y8m��T�C��;!jը�ͷ+�j̆ȓDd('F�#�4��VŜ�E���z����ì�0ep��5�`���Ej�i�f��T�lQ
!��V�R-�ȓY�T}�e�V.:�^؉�[(Z�U��.�p+����i�Q@%�O~8�ȓ+�nD���An�l��o�_J=�ȓ/'����Js�qY���+�-��xSf�c�IJ$t�+�d]���`��Sf�Ś�j�0r簭�ָ)��|3	�'u��#��>P�6�Q�O.����'�X�'���M#H����h��i�'t������^��<p���3QJ�J�'��2T �50<=2eoE~��L��k#�� ��:V[4��V�c���ȓ~�h�Į5`!�P���n�,��ȓS݌ +�FS�+/9y���*�g�<��ɕ9�j��� Ѳ1���2wx�<��<s���q�#ʲW��Y*&Ȓk�<� H�("愊r�:䃐��o��"Opp����XO�	���B?z�4�Q"O`��V`�73@L]�"9��
V"OTP*��+&@�X׭c�$��"O&\�S�؆l=Zh��8�Q
�"O�%*3�
gFt�Q#�;d����"OvY@�N5)��4�ڠ{>.X0�"O�p�2ɐ��6<˃ꘅ6���"OvE��ȃ��9���ܼ"�J|�A"OD�A���n�j��mF�f�x�1"O� ��a*�x(���!>рd�"O@��#��L�Gi�+�`LK�"O �%H�3|R0�u�4>�*�"O>9p5��*F�,P G�8���d"O���_��k�K��M�H��"O�����>0�u[R
 ,7�q�!"O�jFM��~ �T�@+=|�T�"O����Q)]9����O=Sr��R�"O�P�J�e��e!��MY�I��"O֤P��\�8�&pA���DAhxR�"O�R$��d�3q��H��"O�Iӓ	�	 P��qDP;#h8��"Or��4���TEH�c��e�U"O���2�!��Q�L�Ӻd�"O������'2�;b�D��r�b�"O��9l��`�FeBSPU	�"O�D�"�= ���M��PU�.T!��;��1�F�b������!�	L�V�cĪF�3R��u�Y�?�!��%i��93`Ҁ>��8�	�66\!�D�	�r:B�����f�\|�!�d�*�؃g��P�����)�!򤄜Qr�4��\�����V7s^R���S@����m� ?Pؔ+��׳��م�Y�D���-��#��0��?[�`�ȓ5�"YugO�Z�c&L��O*�q�ȓg����N�v��h��'|�&݆ȓNmH��cN�>���@��%v$�	��1��/_�q�� lѸg�؆ȓe���sa�4#���+K�F��8����$�W�|����P���gk:хȓ���m�=C� �J�)J�SD����F�t� ���-`����~_�P�ȓE�����b��@�b$�F��=�ȓv�b�B�`��A����b^�0܄ȓE���.jg���W�]=b��E�ȓ |�h��-óR+���P�r"O0�p�'D�&��h����`"OVu�r��/p�,�@+��yO�Hhf"OUHcA#|yIJ�JG�dZ�YЁ"O^���e�R�(�g���!a�%:$"O�u;%l�0��aVJ�	'���Z�"O�����'
r�T�,ӎtO "OT� /Q �(���R:~<� "O�����W�FAl�DG�-�u8�"OحH6F �i���Y���o �"O^41�a
80�5SԌG�+언 �"OF����79�(t�uk�g��p-�y���h�飅,#^,�"�.�yB	C^@(c��p=�)����yr��#Ir��y$�Ŭ=E"���X�yr�^� �,��: 2i���ԟ�y�/\�P.�M�ȅ�?4䑒�H!�y2�I�c������dE�xAgFD �y
� ���cp�ߋת��A"O���L h#ڍx��;+�R��"O
�ؔ�H���r ȄB�Fz"OT�F&�+(�
�i��@R6n��"O���]_㶭2En!T�9U"Oj�H5���� �!,��H����"O����O�>O�61C�
�
��-ɢ"O��C���+8e@A�F���?�����"O�C�G^�U��TX��K�x��"O�I�Ŧ��2hr��e�Ise�V"Ol��`Q��� ͊]�
]�U"O*AZ7��8�������1Ӻ��r"O�Qx���v��(�c*/F��9��"O�Q�eo�("��6)ѕAj����"O �2�G�PD��M�?'��r"O�d���P�J�͗"fhak"O��A�]�G���e�$a�x�"O�lPr �7��n�RK�r�"O��[����r�0�MR�n>���"O���Gj/c� �q���~�H|@�"O8`�bCV���$�$�ɷ���_�y�Iw�,p ��X RCF��󊆯�yM]5JK�a����=N�V��C��yE]�:�����\ON�A�&�y2�7G=v�� bE����f�=�yrg�-w��I�� !5u� º�yrϞ�NgLA�OU�m������y"��$����5Nq�P�AF�yr+�+3�e�$�5Ј��/\��yb ��fߌ��#SZ�0QJY��y�j
�,��6m��{�� @0���y�a� ���x5�|���P�ygB�m�h<�v%�ev�� D0�yb��9aJ�I��K�%X��0�L�y�A��a��q���M� ��rF@��yR��4y(H��1���� $9v���yb�B4�h�C�� �$�z-�E��yRi�2x�!H]�G����o
�y2�l��A-�J���,��y���#��Jff�pwBT�H�6�y��D�x1()�H�'mm�-:,��y� �y�)	��hƲ�9šώ�y��O�$�𼛆�фnUv9��Ȍ�y��?4-����)[�`ϊ�!��Ł�yR͌F���s��0��|(w�y�G�#�xU�"NW3�l���T��y2��0�EX2+��T�o��yr!ޤtt�%bш9f�qËZ��y"ꛐW�h@c�AÖz�p]���ĺ�y����@Pv�B��p�F���y�O�2��b$)�5e�4���y�V�J���a�杲W�F� RF3�y�� j��D�J%W�����)�5�y"$��F�N�`�3I˖����8�yr�h���`U�,P�Ԍj��U6�yB'ķ5�"T�C�K�En���1*V��y���3O�4�5l����Á��(�ybU>B��}J%�W,���Hr Y��y"��dI����.��� ��Q�0�yB �]��x3�1i�X�C�3�y��i^��`���c��T�-��y����p*�W�6Y��$��I�y���-p䵡�A������I��y")�9�<�<l+��0�'f�*���S�? .�Q󨉩ln�Kd���SHpu"O�=��M��04d)@bn��a"�*"O�=b3��!�2��jA� ���"O�]if��LL��ц���s@"O�⡀G�N�ʽ��M/m��|*"O�,�FN*6UTMs��م��e�4"O�k�� q���FP�q���u"O��� +[�$��0o�J J$"Oy0qLے#�y�� =5�	�"O��C��-��Q�A��T�ji�v"O8�c
�B���;2�ԆO�t�&"Ot�P�������o�	�N��"O�Ek��V?>n�d�����"O� �, ~� c܂ �d8�"O0h�@$��Х�%��;�^Pې"Ov�&�Ӊ�����a�DuYR"O
�s���D��I�"�*c�f�Ȓ"OZܓBFR�X���;
٢�jii�"Ov���G5K�Pŋ'@M(���"ODPVA��1��5��f��H%�H(�"O:ܘ5�̝z/vI�E�#�2i1"OTy#�kʹ���рm�"��(�"O�|����>&����ֳV���1�"ObL�C�M�+Π��s�Ss�L�`@"O��$�����#�+� 1�"O�]���B�r��&Ø�TR���!"O�e�P�
`20١k�0r��2p"O��rCE�$�� ``�V�W��1�"O��y�`��i7�%�pD��^� �g"ORp�OM�LI^\ZSj�2��q�"OP�c̅��q�a�Q�}�����"O���a26*�i*bh�)�@9��"O-x��юU����F�l��p"O��"cᜊW�`=+��A(�	cf"Oޤz5e����b��/7��)�"OD�B�h��v��h��M_6|���"Oy�Q`��m����L�b��D�"O��k'AceMR���.aDZ��p"O6)QC�8=b�ժ�?2C$S�"O�-�skN�@���;�iG�pM��"Oxu��ܩ �>�sv��;*��"O&���	4vR�!7+]��yd"O���œ�+��r��7���"O^��	#2�Aӛh�����"Oh��'i�HR��� �ɧ�r�S�"O��0VE��Q� �[�C�k�J�R"O"�P�G�(�>����R?�^��"Obl�B�ͫ92��IF�ԙnD-�"O&ܡf+@m�Zq�g?i	(|5"O�!*�K���H���� a(���"O�� �ѭ6�����Ĕ[���R"OB��Fc�*I<�@ǲ<90X��"O�9��Aٮ7W������l T(�0"O^\q�e[/�����N;@�v�R�"Or�I��
�W�ya��݉$�f�{*Ov�k��ٿ&`�� �Z(��')^�k3͞���LP�]��v��'8ݑf
s>d\�C��p(��'$�z��΁}&�%%�_��p		�'9]`�6r�N�
�H����'�4E�K_�l�LH�M�c�@�'#,�+�C|lPɄ���Y�>�b�'�p�xDlG�`�lջ�)�=>߆dx�'�TĠ���990�#B��a-�E���� �1�ׁ��Lr8b��
=T"���"Of�p O�!��tm�2sG"Ax�"O4i2��'�x�2�Ʌ�X7��X�"O�M)A)ǎk�.�9b���*�9s"OjD�B�˥v3�H�'��
�e;�"O��CB�r �xŇ}����"O��ؗ�� wf��y���V���"O̭*��Z �P *��G���C�"O���Ek� r
�I�<HԢ��F"O�	 Q�^�T��'��V,�-�d"O�M�å� 7i�E�tQ�r��a"O�t32nق"��(��E(jt��"OL����v�"Q��߫A~�+�"O 9#�
�����)u���TАk�"O(Y�u"F��+\�V�P��O��y"I�r�%�"e��T@")CacC��y��@�|X��� d��N�X]�#O�y��Ѱk��sa��Lrb� w(j��ȓm\����C�}����$�2$��0�ȓ@�]��OD�z�-�A)�+.X��5r�4;�/Ωa&l!z�Fq'|=�ȓB���F��[�l!K�.�$����pK*��MI�T�.|;p�W��ް�ȓ�t�(`ט5!��3W���]z�9`��8b�<��m֊47�a��2�2�BS��F�
XK��]�`$��=7���+$�(Q���u+�;�"O8�G� �a�rd[��Ã���""O��+�̐� 8� ��j�z%�"O��`�c��0�TN��d�4�b"O(钐��(m�2�(w��r�4"Oε8�)�>y�����<{6�Ͱ�"O �YӇ�D�@HC��9��=x�"OD I4aŸHK�c��ӵ
���"OJ$�A��)l�Z�v�P�X����"OL�ɶB�g"@}c����<a�"O�l��<c�N�s1��u����"O�V�/8�Ԅx�K�BD��a Ƅ_�<q+��t�P�ǊY�}��y��X^�<&I��"��E���Dny�����a�<i6&�;j=�З��6e\	�Y�<Y^�����"1�v���BG�?�!�D�	"hӦ�]ym� �#_�!�N�cxr0�Ֆ/z�ٖjI�r!�D�sX�}* �gt��R	ժyk!�d"J\�����K��7n��cT!�D�>�6��� ݙC��0�`��?@!�ė�8bP��'��Ґ0�b R3i!�D��|�����}-�	��̍;!!�$�k��9r&��Iòˀ�y�!򤁰���d�6%�\}23%�71!��L/C�j�C��\>6�$U7�W�`8!��ݧ)����͍�jᨱlSU5!�Q���廣��%��(:���!���%ΈXh4@�:�v)g�դ'�!���y�]d.F&����Z�!5C��R]��a��	p7�X����(�<C��:0��$I1e�J��$��U�C�	-s��q��O#m�4<��LZ�Ol�C�	>i�(�3�
���ŹvC�	���)�	مE��M��!�@C�I9�h��X�X���üD�M�!"O̐yp�B;_}��ˤ��av��"O*�d���' ��9�%Ձ^�d���"O� 6\
$�	
V�ƙhJ�+K��Ԙ�"Ot�:�*�0Va�M�B�ܟx���P�"OzYB�/3d�>屆��"8��"O��H�o�  J�9�Ԭ �@bxI@"O�IC���L��r%�6 ���"O�PA�Ɓ�p,@=`d Y�b��@H�"O�y�T	�>�� ���Yl��""O�LJ��kfdl��m�4���t"Ox���胏k�V@����1��y��'pP``��LA��⑌Q���A�'5�q �.6gp�P#�.Ό�
�'�z��O�%<(��	J�@Pي�'� ���/	�,RXL!�* d�p=��']9�'d�DuxĠEB��`�'��&�	�=��D��2I�4�	�'�<L[F�@�2I �ȹ+�d 	�'�h�����T2���,�P���'ᶕ0� �8�ܕiQF[�IP���'|D�CD��{����3�\��'}b���8�@H��\ Z����
�''~��GeX/���)q
~���8
�'�Ό�F9b�p����u=D�[	�'�0U��䲇.Y�<�*%J	�'�*�@���4nD<�����P�Ɖ�ȓp��!*&聣,\j�*�o�#!Zp$��(X�����,Pb|�7�؇C̰��6�m�&B��ݸ���ºx�ȓ"���䢎�m�u	�̸�,Q���~����D$`�a.C6L����ȓF�|�q�
)�A��g��Sd���4b�p1��Q ^X{,�)bb݅�钱"f�X�@�)��Wol���Cz܊��:i�y"�q\�Ņ�uϴDxa��~��E���Q�|��ȓ�v�Pb؄F�b����"*=,$��\s�L�U�%sԨ�l�&0���B��eg��9G�D.�@��5��=r�)A�p"�SvN�g0��ȓ&��9i��%jAB�C�J6n�ɅȓK,d�s��m�TY�瀇p`���� ޶B *hH�3��7n��ȓn�Y�. +�Z��`tI"v�#D��ZqC�	R<UB"S�*S��Ӄ)%D��"5h�϶LZek�=f� ��"D���NЍ}|�Z֮�n����##D�L�UgV�kBh�q�_��b����,D�0(�f�	�BC2�@�S�x!� �+D�\Т���� J��^7(v!���*D�<I��&WX}�`FX�[LL�qaH)D���e�o�DJc�)w�|\�"�:D�؁4�^2$B�JAj ~�0�K:D��BN��.)�ɟ;x��tc�n5D�h�g(� p:�z�Ϟ�Q�Ca6D�Di��km� K怂($zұ�V3D�����!	�P�S��k���Ԯ&D�\�6�P�!'v��AM��T�|��"D� �u�ֺ v��n����16�>D���B��pdH��Ά<ʢP�%>D�T ��R>,X˰�ȯ^$r�*B�=D�ȳW�O�90�a��/F"x�x �:D��a��B%4&8�@����r�-:D���Pk��\:A�dm@rv]��d=D�`�e�NC��I�0f\(T�I�a� D����F8Z4z@9�ƽ/(�A��"D�� ~�Ʉ`<_Px����y����G"O���-
�x�A��&z�~�X�"OD9j%��C-�(���b���J�"O(1��I�m#4q�����(�"O��j b��(/v|i�(_�u�<�Sw"O��kb��,Svֈsr��W��ia"O�]��#�?s�n�����*!f�X�"OL� E\���
V��!6i`��"Oʥ��C�qF�} sdE� � �H�"O���Т�0Vذ�$ƴ����"O|�� ��8�I ��Z'n^�v"OЄ���bH>��`E\�AtaF"Ov}s"�%/�V����h�<���"O�a˳��2/"�Ш���#}��'"OD�%�f�,i��&;��� �"O�g�ؤI��	��!=�le�"O&A@W`��2������P����"O^�J���w̲����H!܂%Yc"O��A%	X%�@"���%<�f"Onc ��=u� �����?��S"O*�d��)9rj C7Ďm��	�"O�հ�!0&\��s���@2�5(s"O�\`�̵	��}WB1{����'j�DQd��O�F��`��	�%j�'J�q��Ў2�:e�Џݼ+��t	�'2���C8���rh�9~�u�
�'ޜ�zg�5�yi�-�����'3� ���=ya�����K�-[�@�'
�BfпRܦ�� �T,-�Y��'�|�0#���J�]=^ڊĢ�'J���Θ�.F���fU�\#}��'ѾI"��� AA�f�Ӧ%7ꙁ�'��1�s�R 99�A�e�p�J�p�'��!"p���`yp�i���%B�T�<Y��[R���&�7;0p�3n�P�<)�,�Zh 1*��Ň*1�Lp ��f�<�`ү0���'�D�`��,Q\�<q��R)��#����^�1&�ZY�<�u+�
^m�`"֬9�d�)# XR�<�b)n���c�&!Z�qva�J�<���bD���-�56�!�a�_�<������=�	�Q^Pi`�@�<Y���G�L�p�.�O:���F�A�<�FV�6�B�K��S}�bY�Êe�<IE��J���
��+;����	L�<1dd�k�BۏJ
�97�ED�<9ը\>�ni�ƅȤ ^x<��'FX�<�A�	�P��(�n� G|R݈B�Qo�<9�&�^	��0�H�WU<�!��i�<ɀ�-#�V5�uLW!\8�y��a�~�<I���N ��:A��+4��"�!w�<��vԨ��1ia��3!Kq�<��ߜZ�B<�"�@1V�eӡ�g�<��'4����2!�0����c�<9�#�,\x�5�5�P,D�=�gKb�<�&O�Np�Z3@��8��r-F�<��(�={z�h���%�*��w�X�<A�j��h@ �6(�IzDU�CN�x�<1!Gèum�@K��Q�JY�ce�p�<a#`X�+����a�ѿlh�Hq(s�<Y�jҊj;���1���8[f�S�<1���[��diB�ؽ����"��i�<9�-Vvn�k��U�,�Ѕ��f�a�<�Ǐ@�����T�z�����h�<� l��!'ߴo[Zp"	? 引�`"O:�a��]J�H���
G�J���"O�|rń�	����ܫX����"O��#s��9Ē(bBƊ�~޺��"O���lF�z����20ʮH��"O� �h�4�й/u����� H�y�O�k�D�����Ҡ������y2oo��X ��)kLcƄI��y"���G��lK�GS��2�Y�@+�yr�K;}��p����{��q��H�y2cqpdԊ�N�q蘘2(��yb�N��t`�K�&?TN���BT6�y"�1�Ҁ6�E 4�A�d��y��­A���Z��"$*��5J�yI��W�
P� M�MK|P�� �!�y�f�	+�e���H\�Ъ�ƙ��y�I�8vs�I��Q�E+�:����y�
�#{k���EV�kFxx���yb��j�h�V`�l���Ì	�y�{^0�A��X����+A�y"�ɛH(�BWH�O�
ܪ�d�ybÐ�E;b�q��P��|�q]�HJ
�'��]q�Ď�D�8�S�ǏT(��b	�'pҩ*�m(|�Q@-^�^	Ĭ#�'������>a|� �bKT&,�T�	�'�[��2�Xx�K0L�¬
�'����
�+�&��(�$5�	�'ExX0�B�*Y�w��&%��h
�'\�Z�bG�wa����
�8va	
�'�|u��Ζ�E��l��F�F8�	�'$� D(��M�80k��52@b
�'�L�I�4�Ф�nƈ�hM��'W q�&G��u�uJP9yd���'�d	���GQ�y0%B�,(4P�'FZm+���Wm��2Ѡ��%M����'3(��D�,l��J�HԹ)�-J�'ՆEi,G#n��H�脟lP\���'C�<*V�H<C��}(�]:P=��'n|���+�`)珑6?�q��'�zp���3v��F ����'�� bb�S[Ҩ�&?|��l��'0P-�&b�ش���tP�P�'�z੓fV��dH�I�r�.�(	�'0�y���^҈���L�t��A	�'� jb� }�]�(ZM�-
�'�n���!#��!�&�h'����'_�U�c'k�b={6�15:���'�B���i�.)T�S5��>w|P��'�N��'�,<۲!�#��m��dA�'��	�aIы#��
�,Ei�)+�'NN0��@H�i��Zԭ�	2g$<z
�'���gS�z�4��F+�>%9�'Rp�� a��C�����!NY�S�'�j!@��ФR*�e��0G�����'����*5:)�!�L1N"�!��'
�t����L=$#�E>X$�x�'�(���(>;�j�bЧO�a��
�'u��C2"ڻ�Q��
'�ⵛ�'܂$	w&
jD��H�+8 n�pX�'$R	s���*I"9��L� Hl��c�'9��
��S�f�
WfW�Lz( �'ؘ���8U#����$SɆI��'\�#T`C�#R�4)��L)^�H��'KV(h4���<!z� P�
%��Z��� �-�E�
c�l����j���1"O<$�G{Ā�SDb�q���aB"O��n�%�LaF�ɼ[��X�"O����ǭt�l-�w��-j�t�cQ"OP(J�IR/4��Qt�%8�vě�"Oj���7�L=�Cm��=`��cp"O�E��OǛP\n��ĩ�F.���"O�h�6IBBFn�(pg��(6�D0 "O��c�ٗ*����q*(p�"OT�y`G��e��4Q�fp\���"O�L0E����SEĀ�fR�83"OJ!����8P�(h��h.t���"O� ��i�|�q6�Ɵ5���Q"O�8�4+�r�xBZ��T�"Oʥ��)�4�R��b+G�����"O�a�f�ǐv֢��I�z�L[v"O�s�>a�<Q�	V�Zl���"OH���c�~��aا��=QvL�"O�4c5 L�>�mB�NB!(��"Oi�C!����4T/���"Onp�!+�V�N�;tIW*y��A�"Opi�V)�g��h`WE�b��k�"O��[u� 

����ϒ[k�y�"O��1�Km<�# &A>5`��"Oh��f��p��ys�ӅkE�S�"O YrCA�P��4JУ̯Y;z��"OF9���Q�j�q�M�I5>0[�"OR�猁�;�9�t,	�Q�$*�"O�¦��"
?�e��j	�nAR"O�ź!��Q^��BI�>r� �"O�T��N%Z��=Kb�ˆ2u"O����Δ^\5��ۇI�
�x�"O.`0���Q��q0)Rw�lY�!"O��󗨆4[x��H,2�t� �"O��Pȗ	T��p1���e�"O����+�N}b2��֢\F�j�"O�Dh *����* DWe¼[c"Oй�m1P��!�`�N�Dt "O:i;D�ƅnEI�o\�M3�9jr"O��$U>
X��`.��	D�  d"O̡i�o1�b���,^���I�"O�=���@�X$�k7��o���Ӥ"Ot,�� �<�j�b��/���0�"O�ȃ���,N�!��I� 2��H�"Or��� ʄv���ǒ s'��R"O2Eӡ�#Z��'�f	y�3"OR�#!m�8O$F�{q%Ҋ�`��"Ozeq���H�\X���H2�R���"O��j6h�$Z��Y����$J�ʝRv"O�[��H9����!�3ĐS"O$	�EfΜ6,�"��"tTH��"O,�@QM����)�
��}��h�d"O�4e�Y�{�с�h��}���Z"O�X�h�$D��t�`'M�j<�aA"O������Ӯ�b���5)y��"O�1I��_����V�Ԕ%k&��%"O� � �B� ��9$��#�:	�T"O���D��]#  �I��n�Za��"O�4!!�{%iX"�Y2{v���"OL}S�C��<�hQ�*tp��"On��0b�>9<0a��גDu(�sS"O ٩!*PO���&큩a����"OD�2�[7`'6�a��ɾR!-�v"Oaа��yh��Y2�ܦ.����"O� ��S+�Pcd,�jзQ�Щ�"Oh�[��G�i�6X���Y��a"O0e����,r�,�ʳ"Ҟ%��Z�"OV	S�fA�M\<�ȧ[�`�k"ON�he�O�;��p�0�Ch����G"Ov�B���5}�L��q�����=�3"O$Y�/��w5�CfZ�M����"O�)" C(FƚL+� Q'N��E"OhЎ��r�$b6֜3	�\��"OHy�f�o��$ q(�X��y�"O�����
<����"f�2_�6�"O|�"P.D�[��Ԁ�d��K�:�X"O� !�&��|��	G����X""O�9��1C��;�	�<��̲w"O�H��朖z����Qʂ?|fZ�2�"O4K���C�MB���e�ލS"Ox}Q�,QD&}Y�hċAT�Q�"O��yGK9z��ǘu.���f"Orqu$b)R
�MZ2F�r "OI��]d���Z3t��A"O:�XS����JA�r��6k�#�"O�i�r ��n^��� ���"Oi���B4]X�ԋ7�¤Q8fY`�'�\jd��(�عp�ʏ
�p[�'�z���+�>v��A �z�d$y�'�F�S�#61��P G�~
XjՏ7D��#M�2��d@�P��ц�3D� ��@��l�r�׉\�ȵ�/4D���A@+`�� ���T1O��w 2D�8�@k\9k��݈R
D�eA1�;D����R�KC磞�X<��Z��7D������AWj�7�7h>t�!3�4D�(!T��|A8pQ�OM8��"=D�|��镁������.ْ$.D���2�ڝ�q�0�� i�`��@c-D�D��㑬_e�i�dY�Qf�0��)D����J�J
|C$X� H~�J�)D���}l�
��b�
@�C1D�0�CJ� o�iB��
%4غg :D���P���E��X���^���Xo,D�$*E@��h���SA���H�o>D��P�̗e04�1��f�|�Ha�>D�a���T�T�[D��mnԒqK=D���%+�L�$� ��5�ja��9D�PF�]"T�La23A��PO9���*D�4�'�W�24���L�����H=D�|��B^>u$�h1s�˥-@�y���:D����x�xJq�^ (�h����7D� x*����Ʀܽ<�b�05I1D���`�E�{��b�/�	`����9D�RW�߷D��k@�I�fo�Ű�)D��R&���O0��a��5T��R�L"D�0����D�<�D������g�*D����Y	'��E��~��h�m4D��1�@ܟ�l�u�
�Cɂ9l/D�|ԧX�U^:! wlJ2G��r
-D�l+�h� _����Ԏv��\r�*D�$s�AR�F�T�T��7|�W.D�P*s�99$���dPJ�T�N+D�h�C,ڂc*F�)!�[�2��T`(5D��y#�C`��`FǍ�M!ц�4D�P���X�b���ϭO�����2D��qt��m%�V�̲b�˧�:D�|�W�����ī@M^)u��<v:D�� |q�����9:M�qG#h,=�"O�D���Q�SD�%z�e�+{:���"O��j�KL;5:0�
��RY�xU+v"O�АԌ�%F�ba���C8F�*m�"O�Q��k%yЬ�� J1��"OH��D��-G�^��N0g���"O�(REğ&��{լ�	b߆i��"O�$����bb�9C��$��I�"OP��AN\r:��SҠ|���0�"O��#�˙�Y��`�e�dҪ�I�"O�-���,Q����Gf����@�"O>X��<��Ia�d)��|��"O�л�G�#��h���O�(h��"O�DK��Oh� �đp2���"O���9mF ��G�O�|!�6"Opp�$�&n�V���oVJ�#"O�]`���^@�*F��qO��g"Ol��~�b��3��;.;D��"O�<!g昳	8��`�F�/&��1"O��U�:
m�fF~"�z5"O��(Do |c���E`��9ؐ"O���Ν�S�d�jԋ�	2<!�"O�9K��ħl�T��kт:��iV"O���N�r����W�-޶��0"Oa@��J,!/�̈�	B�컕"O�ĘVIY't�}�F4t!���� x�*G�Q8�EO�	�!��;K���o�ި�)�c�'UN	�5��	G<:��5J��d���#�'6���-V#G���T@ŤZ�����'��L8v-\�G3*$2t(��Mb��y�'��|�\�W!x����u��Y�'%N�6���]xIzt�̶r�Ƹ��'�H���)�����v��
i���C�'��A1���,4yS��`R�ȑ	�'th�x3G��v_���b��f����'&�8���+qW^�X�&u��S�'�^�`�ڭX�$X����j��8�	�'D�#tN��PC$�ZSo]'O��Ȋ	�'�t$��ʈt����ņ��G;И0	�'��yY�Э5<�,�Ԣ�(s>���'x�uBƃJ<5fI�#�]�,H,��'-|�R��=;@Ё9�i�\�.��'�rLh'���w� i�Η'�:���'v���H.n�A���$6���
�'�R���I��d������'!44�E)�fѸ�IM�%���'���Ae�P�B:��[�~qL��'fvY�LC4A3D 1Gݘp_@�*�'��)���3Meu�qǟ�a�v�z�'bf����Ms�`!b�,,�5x�'}��q&#�K�JH�E^���s�'��`�K=~�S��T&��	�'��8�Sd���)��U����	�'O�!a�U��}X�)�RwT�Z�'RT�$��"u�҈��d�F�����'XR�)�˙��e#�/�(D(� ��'8��![�H"�� ��?J���'m�����"��C�f��7�)��'�(ЂC$�8��2��U��'Rh��$-�rx�t �)0��A�'�u��EɃ֤`q4n�-%�Zə�'*�!-��Zɮ�[�b��2��H�'�:�9p�j�^e��?̨,;��� 2	�(J)B9�Uz�U�{y��Г"O�Yx������O.E]̙�b"O�Pc- 36}&9�c��$fԁ�2"OQ��:er�ɋNM*w~X*""O�Q0�IZ���1lܩ*9V��'_~��C`��@["%P���l�
�'�� �d��J��g�*40�'�<�rNH5�Bh[⇈w;���'�*��P��'-�ahƩKᒄ�'d�Uug.��37�K�.t)(�'(�%a�(44��&�
,}�F�H�' ���`,�[]}S��Nt��;�''x12����z��������lB �'\�љS%Or�*A�JK�NQn8�'W�հV�BP���;e@BBR2�'��Y�"�,�j!s�E
m;����'uf��0Q�$�NL�sU�n�f���'Rb��aa��S��6��;�'us�i
>L3ȕSd"�,�}��'��J���2�z!i�jT$�y	�'Ű8�SH�ӎԏj2L���''����cD"M2�i�cʈ�m����'Y�$�PE��~t.�rc�O)(���'вI�C���B 0����Jސ�y"A�\Jp�C�� ͸!�T�֌�y��̷ai"�+\�B�ϕ+�y�
�$:*�م#!D1���U�>r����B%�CéR��j�SY0~g�|�x�l�W��*�"��hxHRu��y��9Q��� �h� �@�*2�y�"O�Y��@�eK
Z}(]��&I��yRI��n�)���L�~�j�(�yR�F�{���ٗ'Z�BS��	�K��y���PX┃6��8��V����yB G����/3!�����K��p<Q�'�qO�� t��-jL���SMb<��"O�h�dQ�S����+Ԯ:5:bg�x��)�S�v�D��vY�cB9�Ǯ��@��C�	�1E���`É�f�(��4`	9�c����>����&��6���:"
;p��C�	)<��Cu��4���e�M�V�C�	�I8�R L+h=^��#X�����Ĕx�'�Fh�bNovh ��U�Ԫ*O>c�8G{�O�=g(#|U8�!a�	5 �L�O,�DzJ|�' u˗�.]ށ��t'z(	�'B$ya�Ÿ&R��@�Ӻr�H(�'q2�b]�a��!�@kP�g��R�'�إ� �%|��щg�X�Z��A��'}J-��L6N�BE��Ȗ�W{z���'�2@�f��Be�It^i�T�W��� �O������uV�b�Ǌp��9*5"O�|Y��J�{��U�t���R���"O���4���p�5+�'�X�
s"O�|�0��p���ߌZ&$�"OΘ[��^Xͻ�@�$wΕ��"OBl0Th��9'�0� �F��~���"On��%ɛC�D�J�O�
a�a"OT9�����2$D2U򌹙�"O�����F9�}��G�5=h]�r"O�,AЎF$Y��"� �b��p�W�'���&	�,���ŷ�@��a&�"+��C�I:r�$�VGo*�$)��R�g�#=)��T?I��E������iђ0*�!� 1D�x�EI�V��h��A�z����7A�O0�=E��� X���$��s��؂��Z8FL&ؒ��'��O2A�g
ޱ!��$*d��7�`y��iLI��W�S�O\�urW>����qſ[V�0��E%�S�'��ɵGe���5�<}0��m�����<�
�A\JQ�!f�$�:t�։ȮY�m��T>�Ex�
��\i����\-�����d\��y���]�QSъ�v'�hf]��0<���D	9_;(��CT�%��X �̇s'�|R�xb�����C��:<S�E��;��d�]���n���.G�Sm�`��xV�t�e�>��>r�3����H� Y1���`(0����Xy"���_�x	h��"W�r�JO�)�y�MOo*���,���[§3��O�jƋϹL6p!0�^4L�era�_�<���*:
Zl�@Dq��0B���v�<����+A������<EJI�u�<Ʉ#V�}ӈ��V�'Ix�U%�t�<���x��u�ՍC�� �W+q�<)@�2X8l�w��10V�1���e<1�Sf��f	O�T@x�&��U�0F|B�ӍW�:7��x�;��3[\�B�a!(�`'�D�)<<H���ͧv�B��1T���H$!�;*���2��ͤ`_���hO>��T���EPV�>spn�з=D��&%$6X�Ȃ�(8@\���;�O��aa&p��C�	-
8ӷ�3Br]��p#��ɖ��&HK�^S��`L���Op����UJ�x�!(0IOH�[f�M�<��(�8�P�1�(06:	1��F�%�c�g���R��F�%g�z�C5D��͖���t{q�"^�a�O1��9�O��`$�E�P�Fu*be��3�'�����n�R,@-��#��H��~b&(?�V��<�|�r�$sLF�kb�Җ9���5j�A�<�v�Y�~m�t�ׁ؎H$B���G~�<1��C�t����Rȶ�R�m@f��Q���O1�U��f�'^Y)A�\���q�O�0(�O�O��0:�˃�P1ɖlA��0Y[�;�O~���;B1c-�s��@���c����)&�
��V�_Z�Y�1��
J$����;�D~�,
6��3�|���6>�R�K"D�DY"�L5w�(�Pɗ�ߢ��c,���~۲m"�`)i�@+_�P�0"OP�v C�*�\E�)G\��E�!"O��'�]�,�r��J�hl�`�'L��N?���0C,e�7'�5X���I��^R�<�A��{b��-�/%�&���Q���d5�3�`!z�����br%Ϙ)����ȓ�fM ��	D >�BpbEA�	��qx�h3��ys���ekŴp*a�ȓl� ����/u|��W*F�+枬�ȓ\jrW��L9�!�-X���'��O\�v&]� �\���3B\Mr"O]���6)tP,R0�ΒSmI �B���O�.��Ah��Tl#��
��}2
�'��!7$G4�F��&I�VP��'!4듆?�(O�3�	u�F����S�q�`h՘��B�	Q#�IQR�@$%d�r���p�5�`"O.�'�������i�	#⼼���	Y�O�����
�x*����b�k܉j�'�p��aɷ1>(@�/��\�D�y��$0���L�PIŰI�U���{�ч�zM�T�Ś?HC���B �\�ܱ��y���0}A9�X&z�f1�bH)/�C�)� �x�G�O�GQ8acD�_�T�X����O:c��Dx�NGB�#N�#�~�ӕ�]���'=�OR�	vyr�V�Y�4�� �ɚ2�����P!�dֈUӦ���*J
s��")��2Pf̓X.�'��g��~��T�T͸�ȃ���N#b����Q�IF�6��"��,�E7A(@6�n�I>n�Q��Od�`�󂟖��}�B&� ��!�	ߓ��'���g懤@�� a1�߉N��"�'�"������=V�0~�k�/]�E��b�t�)��.Γ+���yƈA7,��M�s)� l@h�ȓ` ��ʖ��9�~��@�~��I�X?au�x�KCp�'STE����D)�� �
�W^5��'���a߲9ǀ]hK�QZ��ش/U�O��)��>�fɜD��D�)Υ}��M꠯GE�<ɢ��;�&M��&t�Xi���<��x"�q�Q��&aj�[����y2 �sl4T��Gȇ��HP3�͏�yhűp,�2lZ�����y� R1;�u��dR�Q&����]�yr�K�j���96A}��RC×%�y��L�h���c*{��1Sm��y�~1�w�fh !��b��y���de�Ո&f�e�~�h��7�y�	�U���Č��Z����p���y�C�H���e-�)��!G���yb�úܔZE�/ ���-�%�PyR"ָ-:�T
��#��x`'c�<96��8>�$DJ%k6�c��E�<a��Y,e�t�0U�W�K���$�B�<Y���[����C b\  ���|�<��̓�jrz����P�e
��y�<���͚+�V�`P�ܼdߎ)�4A@r�<q��Q#~d��!ʈ�^#l��R#�q�<y���:1mBX��m�a�@=���Wo�<I �"�*���J���0�Aa]`�<�/|��J�A7K/X���Y�<1'��/B�@R��!&R��'ϋW�<iց�#6��|�&�	Rv�Ѡ.S�<'��-nވ�,O�HJ�\�LR�<�u�L(P�x��)٤fGܸ0��E�<Q!#̗>��e��n�����KŋM�<y����mv��ٝj��p�~�<9�#�+3����,��~@L�R�dQ�<I򢅔��efK�,`
���DJ�<���\ӄHR#ņ=r���[$C��<A��^#���2G�B�fJ��k6��x�<���̺b,�e	�1nRd�ȰH�o�<!1o�{Y�L�F�BK̏~ټ��ȓ@�,�PƃM�tT8\1.ځE�楄ȓڠ=�g%R�;��<�עP�� ��{:�2�Dޫ/���0wm��gLr�ȓ|��R*�J$�0@'ظo����ȓN�<��(lɪͨ�8d66T��d� �z4oΡq����_�1F�݅ȓjF`b	���0ի�-.W1�ȓ��=i�d�'^�t8�c�z_���ȓ0(�;�K�W7̠Q�իR��E�ȓu���M��b�8�9&̿~_Υ�ȓ=�ީ8�X+l�ɳ�f��	�fi��13t!1$��m�l���"G���|�ȓ�n��am� `0>�1��g�r����̙�T��']��A��e,ȩ��v��!�%���p���i�T��}
��� ��!G�������=�T��S�? ���2���B�D���!,bI��"OL������M�&�qm�J&"O<!2W�H d��%+���NS6���"ON �%ו4�J�J��B
���)�"O��pa3e���S�f�ri"O�:��V�Q���'��=�8I "O�8����i��4z"�
��ti�"O�Ǩ�T�0���NGa�fHI�"O�y�֪٭zu�)�0���~���a�"O6 
�8`��A�ڞ��|��"O�t����j8!��h�6\��"O��0�`ްf}��zc��� �)G"O�u�����'�,� ��#�!��62* 	d/S���K����!�ȅAC���&J���8g�!�ĉPMȤY��E�=��O�)�!��#T��)C?7�:��-�~�!��ʟ}�d��ۣSٶ��)�!�d�T;�R"�̑Xi�Pv��Py���3bpXY ��� ;�j`�%_��y"�VL{
m�/�,�uңn�$�y�4r�x��^B�0+C��ybѠ1@���20>���I���y�?%�ҥ��	�y� QD�6��'Vaz��K��P�1"b[(&ۆ\Є���yb.�&E�}Xi�	!��	*B'�y�J��D��0�	����)c��8�HO&��'?�яp<��kK����,���<��M�`k@�C�,�>@C���V��U�'ka�d!�+a���Y#DICV���B��ē�p>����a��!���G4b��L��!NJ�<�%��v
~d���E.G�`�EE�<Ѣ!�~L��q�L��r��U"�gMj�<Y�'�;l��5�ίN'Z�!# �Q�a���O:�*�*��~�r�aU)֙2��b
�'e`�jq�@�� �Eh�-@24�!��),Oxh��,m�he���P1_����a�'��D::�� �Fܧ?s��вA�4[�!�lޢ┮�ZI�%`v @�e�!��i����	�@�~q{�G���2O&1O("ŉQy�ذ�d���!��}�<�A��4ڹ0��`I�1���Tq�	T8��9�(O"{�eb��ޖ=�gw���'W���O	���1G|��4Gש�R�g�2@sVC䉲Wqr���d��C�XeX���-L�Zꓐ��0?QH<%?�	�'͝p���U�D�٪U"D��ɤg�+$`��s�><T��<a���S�X�T���Q;G�-[ ����C�	�:�1%B֬lf�@�FI�2��˓�0?���  d��0P���@�z]���V�<6�ȓ9�5ۣ�'��l��-�U�<���	O�8Y�[�3��XGfxy"a�m��6�,O˓�j�ņ��� �#�̰^�����f}����ݬ;�L�p�o^71�|�Fz��'Ťpz��@�F�DX�����\%C��$5������P�Ȳj(&�h���2����ȓ&�Va���js�EH�g
�R$��ȓL�=�6�� UȘ �/�{s���ȓ �����-�}��@��lZ.܊y�ȓW:l���)��� 3*���9��zx��e���#��/�m �Ň�ij|�ZGl y6��7n����>#K��L�h���B�͙�a��4��h<yee��a<���/!���vEl�<� 2��g@
����F<d���;4"O�D������q��r�(��c"O؍µ��5S���	��)`��Ц"O�UZ��!{��� �&�.��"O$0��-cV��{��� �R�r�'�Vq�qۗ�D͖X35a̕W%:0��h|z��Cb¬y�����Β�6l���ȓ`(��9��K#3�A����&	�ȓ9����g��_�� J�*�%�	O}��'��̨�y*��6F6�;�LI|6��pF	��~B�	%"�ͳQF�,K,�;�ǯ.�JB�	n)`��q��:h���� FB�	'����H>�����h�[�'�)��kU&L�.�:�l��
l��'������!��[��sD,�a�'�0iբDs����딅g	��!�)��<2*�<6�Ô�M�d J���I�<��&��A��ːN� ���2���L�<���qސ%	C�E�^�R��Ԣ��<Q���6�����Fʏr$�Ջ�B䉚@rn����N)9f�5��N��6a�B�ɶ\�V��c�ŧC5r��QK�ݦB�ɛ*����!1�L�WB����B�I��`E�DF�!�ιѣc�8�.B�I: �!r6��s�h91'�]�hNC�	$�d5:uX=M}a��%�+�����9���Iy�"
`!T�r�6{;%�O���d�;F�4���@�#� �C[�E�!��[�h62�Xg�W-�} dlȄh�!��҇q�@�EI�&<t��z��[~4qO��������q�
��l,��.�-��ȓ7d�U(�H+W��}2@��*� ��O�@���r{PE��(��!�������v̤�f������H�<Y��.u���׊U(q��E{��Od���㮗VG^��*dK�̊�'w��bl��|��@��Z|���'U촨tj��.��)Q���XK��'�p,��B��#j"�p��a�����'���Q�^�-v���t옗\�d���$7�'P6
,�*�(s��=��,>����"O�1��. 4bz`�;�j�x�|R�z����_��ّ&�i:�����N	o���(Sh%D��s���d樫fZ��b��A !��<�TK���j��E*��5�U�Hi�<�7�ʘ
��9b��)u�@V�
iy��)ʧlE*p�0�	���&g�&|���a9hy����dT��/x)��ȓNp͒V�A;k�1B��	�x�ȓK�b�2�	ް�8l�1��1Ҥ��ȓ9��]���B8�]�iE�cf�la��(���I�_�,ٔC�za�5R%��C���u�ҫ��32И03-T&�p42u=D��y剃`p��N��@�:�J�*z�xE{���Q:q��HC�'g���"A�Z�!�$<"ٲ�G�D��'M~�!� I�����TN(��%�2U�!��
�:��ǉ�%R"���!�D.#QXp��d�G�ވ1!�R�5��іF�+N.�	`�EY�O���\E�ĉ )㪼��M��<�LLs�l��0<!����T�4�t��
K�R%C0ː!$q!��}č�f�L#�,����@VqO�󓾨���#$� � �<�b҅M�D�`�d�|Ƨ� R�8Q [	����Rm͡�X\	�"O��KO/uvX��-ǪQ�$�0�O���2#_"b��s�M٩^���4ړ�0<� k��U� -x�i֤���IBM��'�Q?���o��6��(��iR(w��X��n1D�ԑ�" 3GBD҆�2T�!�Hn�8�'Sɧ��"�D�Z�-�cG*U{�	��ʗ�O
B�	�F�u᳍۪p��#&L(��C��l�T��0l�st�!
�*��d�B�I�;4d�dk�z4�E8B��,�xL��#p�t僧(�k���=[.̈́�O�Ъ�DP6UL��ȧc��Fz��'��`��MϯW�|���&V�Nd���D1�*��F�S�+�x|� �	�d�x�"ODT�jI;��	�菋H@蝑a�x"�)�FZ襚�/S�m�H�x��C��'�� �'�8����QiHC�Ʉ<�$ "d��X;��͊yhC�ɫ]R���Pe[_'�%2+зp�
C�Ik��}�Q�AU�������Т=ɉ���OF0h���&#*d���P�v����d"O���PNUWaN4b�aQ�u�:�Ar"O���ܑɮ�x5C�D%�)R�"O�ո�/ܐdJ�$>,t�ت"Oج*�(�3�H-�߃j|�"O��z�gI�1j�U���2X.i`"O�[f%�{p�'ۓGSL\�'"Ox��֊;�4'�>tJ���W"O��P�΂"7�4ؒ!>f"̉�"O�C�7��q3���o5��J"OD5r�+�1:�%!D�x)4{�"O�\{փ7�\�R�@�( v�z�"OF(ڒ�V2r��8��5/����"Oi���gMb�jZH�ꄎN�x\!��Ϙl��
�ǒ�+	�t�C�D�"�!��//x]���W�u�n�*�㚥�!�$�=0�΀;"���}�SE-k!��F3e%p97�0iB��g�~!�ē�[Hd�{7�H=�vi�D��B!�D�;���@�M�����	ÆG!���&��pD܉jv�3�eͤ)!���(���ǅ�P҄/Q�!�dM�8����6!MCS�١�#�j�!򤔛E��`�4"F0o��eyabY	q�!��yՀ�[�;v�r�r��;b!�䇅/;XmhC�
~��ՐE�P� c!��	Rrb`�/ݼZ�z���A6W!�d	3E�� ��R�=҆p;� �Py�N\#Dʶ���a�[�P�T^�y�T���Q"��(G���3�yR�^��
�R1Ƣ%���.^��y���>vlJ�e%:z��6���y�N�5O�	b�-�
^��sf�y�L�f�Lź%'����i���y�i�W&��8cQ�#:j��A��y�hA���!�j��i�g&�yrH��$����j1�iY�'�
�yZ5rs,(F@Z+cgz�0%�Ӊ�yR�C�B��u�q��	�NK�yˌ�m#h����7Y,e�CO	�"��t���'����G
=�@J�d�0'N	)�'��6kQ�y!lK1� )�~u��'!��c��I?P���{�86	��b�'�ra���	JmA�k�8#,����� ��cKC ='������	*9��hd"O65�0*�9#,P1@
^m�(F"O~��(��d�jy�s�R�`�j�Y�"O:��b}ɰ2��_�", �"O�����	��`w�
�2��g"O��Y"EȚ�%���д����"O��H%��+Y����RO�b�I6"O~u�rn�-9oX����	;g�f�"�"O���w�|��#���{n�pÖ"O�� ���"L��f�XM���"O��J� B;H|"@�g'M�m��"O��Ŏ*�v��7+;Z�+U"O�p2p��LǦ`��k@���)��"Ol
ō�.v��I�$��D�ܑ��"O�њ�9T�0С�����1G"O5��H�	I����uc��vq���F"O��0��3ag��pv@�Zb�!�"O�Je-^6V�5id�@6hpj�"Ol�1CP�>*������@)<���"OX4jS뎱k{p� O	(�^�h�"O��;a�E�k�\�C�@�q`�q��"O<D�ǅ\&z�޸�FꗋTYf�г"Or83��&s���z���M��
d"O:�#e�A IW��Jݻ~�r�"U"O�� �f�T��ŉ��{��])E"O*�1�F��y>�3b�YX�0�"O�\QsH4lh a��6^���"O�,2�$N<5�2�"'c�/2FH`�"O���iZ��a��=<��"O���TCW*l��Cԃ�k�t�s�"OjuhU�I+W��&��2�B]R�"O�E��	p�v,p�\��)b"O��#�&��0�;��G-{Rhx�"O���2l�%#� Y@���SaR���"Od$��!!rc�����*0A����"O``fm˼��xQ�nʍiN�T��"O�9#�L�ŀ�8��%>�u5"O��W�/v�Ip�D,p� �"O�U��	��8���o&�`�F"O�t9w�TC#���M��%T�<�����'!�����X2oL�g�l�<1�D@"7��ʄ���{�&��� �o�<)�nJ�4J�oW��4偣�a�<��@��0����g�9��I0-T�<i��9H��Uq���/��MY�"�k�<�L?x^�A`�$=�H���
\�<)拗�qy���Ae�$b��a17CX�<)�m˞0ʶؚi8tWd�PD��Y�<��)+m]D�	BI�2�zu���Q�<q�@��s�[ ��t�d [��O�<�u��|�Ir"m�9��\��D�O�<Q�H� 訨�O,R4��aa�I�<i��?8�b�C%U�}��2�!TL�<at�+<��Ҋ�-9ؙj&�g�<�c�œTfp��w�2q��`�"�f�<�ԯD�Q��-�4��Uiqj�<)��[�ip�(���-�$}�#�N�<	b:���㥀��CSh)�œN�<Y����'�!�3mYf�hY�BF�O�<�C�;O�h)IW%��l��Os�<�C��|��PIw��+�,�K��Ʌ86l�ȏ{��"�g}�%�N)���)٩g$M�����yJ�A��e5�^1 ۦU1�_�@� ț&P����	� �tɐ���n��5�Ŋ3���$Aj��e*�2��)� ���Lv��E~��Х"OFM��ޘ7�ذ��/��Ѻ�xr'�\)���Ŋ�f�G����fݘ�z�G��gB�I0�A���y��ÂV~�� .��@��1�bG�2 .x%�����Y9첰�~&�L�w��Gg�8��E�\М@�
*��+6�ǘi"^��"��#A���Q��mZp�ٶ�Ԭ+�$:D�{؞� �7�Nk2`�*s����D)O�����l���r֣Γ'.�7��=wx�D�
X�ia�z�+!�dW5;f�Y�(1Y_�����P�DX�c���A�"4����g�8�H�b�������*1$�����"O��cs�/������L���"L�0�^Њai\͟$��聹D q��':p�t�� �N�I���A���q(<��	R�J�|�D���BKh���,B�M	���dh��LY��k�$)�=�E/ٌx�$���I����D,�L8�ċ��߬ V2qJ��K7x�o�� qhUɖ�-V���Q�[�^�VB�I.A�Dl��Gьr)�4;��]�^�'�V A$�(����U螉L7�>eJ�����Ԙ��.�:q�1D�0�֫�-	�I���9;�=�!�m�J�r��t?��nɴI���'�P5����Sq�x`E�v 0�r	�'����#Q�I��PEbۈJ�%�7l½,?����I$R'����I�u!#���Tx�=���"���=U|�)�� ��y����á�5T"�c�-Րz��B�I`���3J["nJ:�dG�ul�b�� D'�to���S80x����I�Є#t�J�e�B�	\ۂ�ATG��&7�0BT���M}<xѕ]�>�>�,��E����0XY������hpx�ȓN
ʹkb��"�<j���YQ������DPdV����lU&VQ��>�;e�M�|S�I�q�S5@��Ćȓ����o�2ND<�$��C��=�ȓ~¶0ȥ@ʃ1��qF�U`�!��s�s ��F�!Cwʚ����ȓcr�-��,	9 �9�$#�R]�ȓ#�Ĺ�ȉx(4ӕ}?����|K�|����R ��,U{R>B�ɅX�sN��Q��R"PO�B�?sti��\���D����!DB䉇X�ra�*��JE�q�M1��C����)�R�
Y���ͱnC�3glZUɢ Y�1�0\�Ȟ*-$*C�	�ļ�J�!X�L/N�ie��Y��C�IJ��Z��҈8�v�����=F�C�	�|򪕛���*�*�j�  )ޜC�/~�D렆�/_eF��p⃅N�`C��(��#�-ɨ��I��SB�	�=
z$��c�E��,�̂�a��C�� p��=��m�,~��TH'k���C�I�)��ZҎ$0���%n��>w�C�	 !D�##�
�Jz��3`\
hC���RW/Ӫr�,��n	�-{�C䉽k��������yAW��,q�C�I�y#DK�Z�i�u��3,�VB�	&l�)J@��-~B,X4oB�hC�	8~bi�0�ӝyt�!�j� C�IhR��kE&��;���J��4/P"C��<S|��s푱<�5*��(2�C�0h�N���K�"� P��>m��B�	� (��fM��屐I�9��B�	 6+��EK�P����GǴk"�B�ɁgR|��_}|܄Bʅ
;tC�	/�&(ۡ㓛.������B  C�	iK����j���ᮞ7=S�C�I�VـX;�D�t���sF^�{(�C�I���t�#k�6T����4h�!@ªC�)� 9hsoџY�� �פ�.�1��"O��4�	�{ePa�SlG�Bd
G"O6� RHܻ-�0�w�	��!!�"OB@�5�X:W#��Jr�["�n�б"O&����L	.��:&��:_�t4[`�>�7{Nܨ1c�"K��J���#R�ؔ��	~}2*� @~�� �\*$|���ӊ��y�]�
O�#N�ot�i�S�M(��O�#r��2 x�A��Q7���:���D�<a�!� 4`�p���-iհ$Sm�|?���SfR������Hó+��C�.��"O,����q�4��	�<Y�DŹ�"OH��$���N�]�f�)�U�"OX g[:zdԅ�r�@�r:,I"O�d�S�Bl�}P 'Ms�[W"O��WD->��lq�� k]%("O�� ��0'	v ����kD̉"O"(�k�U(�x�����(���"OZ���.g���'��a%\�
"O���c�%D����C�n�cD"Oh�ȡ�Ŵ+~��+AD;�PI9��'+ZD�
��;~��[(�dd�� T�G�f0^���I�>�p}��Q"ǱR��):���Qh�Նȓf�����%'l��D�!nY� ,1EyR�2�S��S�~��HD5}y�yq0�X�y� ��Vx�MdFHzO�S�I��M���s�Z �0dN�`F�ۥ��@ b�"O@���B�d��{��*��ȵ"O���%��p6� �&BE�m�x�Q""O���Aj�Oڍ�s�����r"Op��'C�k庵�!A�s&�Q�"OH�A^�,��rD��cB����"O�l-��?�2�i�%C.��"O�Bg�F�tHzdO�'����"O�Ĭ�mp����<�s3"O�ܰ4Hѱ�"��m�.�ƍȥ"O�I��X�>�^�p��	�+�R\ F"O�@w+��D�����dX�"OrayS����hń]L��Dd"O��	0-/1ԭ��)C'�
zR"O �t�H� خ1� �Rڜ%�w"OP�袀G�A���(AL�-�0!�"O�]����:|�9+ŇFjr�rR"O��j3�]$����po�)^5@"O��˅MA%�4+T֕|�l���"O|k�JI�!�UYЎ�$Dz�y�"Ob�Yc�MqdP�COţ,f�J�"Oj�PF�V@�L	�W �#O<�
�"O��B��^�>ㄹ�W��6 D�õ"O��`���{z�� � �H!p"OB}Y�.ļA$@�t�U�!븐�"O��"u�G!!/�!���'6Ē}�"O��!�'߇C���w�)Eo�X��"O�E8PG��P�
UX�!� [䑫!"O�x!�+B�r1��� TM:�"O�
l�*TH���x�@u��"O8͠"���"ՑG�ݎvw�X��"OVm���
�R��͈ёShj��"O���
�O�>4�(�z���@�"O,�9���+ ��%�q�"�2�Y�"O�1Pǡ�)����H�<*�"O(0)�D p�b�`f�o�Ɲc�"OX�2��EAru���ֹ1���"O�Hs�ɍe�ܽ���Q0b*��"O� f][1o�D��J�E-X��s�"O<�J�+�K СCdE��U�V"O���9gs�h�KK�b	�"O�dZQ*�1<�	Ye���N�{v"O��$3ru����Sܾ�"O�!�C@�S*h�y����a�|��'"O���v�H�k�&��E,�!/Tk"O0u��M�w�L�q�l�m��1u"O��zcH�C?d�+�X)7��H��"O��H�zQb���+�29����w"O�\3��	:y\h���SqD"O�e�㯑�WѸ�
��B�@!t,�"O�Ƀ��-,r�J�	�((�(�۲"O �Ǒ&PA����=�ڸq�"O���㚹`�0De
:O��@�s"O�Dt�C�
�ĲR�X m�.�`u"O���`�K�"��L�N�J��ܰg"OTh� #ݚ-$&y;w⍺YH�]3B"O�UP�j�kz%� �#O&�ّu"Oz���$]Km��RsZ3C�ⱒ�"O�i���Χc`x��HD&&��0CF"On� ���*�!�"^�#��,2"Op�P��ƾ|22�0cb��e��$H2"O�ɻ�V�{,|1���ʏ�T́"O����d@�XZJ:R ���,�b"O�����i[D�+�&K:J��0Kr"O��1���
���Ś�w��""O@I�iƥ���"��AU�-"O�tBU!� =��=�R�B�%_���U"O���5d�>�:֭ڱ���� D��c &Y�.�����[�,�l!��?D�� �ɻq�l}Cp%��v������6D��u��+$6 bk f���`#D����L�j?
��` 2�@�M D�xФ㖣3>�6N�g����a)<D��z�
F�0 %��8h98q�I=D���6�Ȉn��`��Z��c�'D�@Ҡ�D�;ax	;s�O�B9�-��+D�,�QG��#_�-{�C+ޙ��k&D�p���94I�A8U�ͣ{�ڕ�r&+D����BV���ՋH95�5K�(D����,3SR�ABf�<7�H�3��)D���.F�=�*��Oǩ%(2P��&D����I�*]ֈJeF.�N`�$D�\P��z-�؁�P�} �j�F1D��W��#a����1�/"C�]S�J0D�p��<_�^�r�͏�ǂUUf0D�P�g�)%�=JB�;Z�z��tB(D�P���7b�\ �aG#�|I�rB+D�x:���i��#T⏉|n�M��h%D�ģ1*@�*��H�mЅl���'#D���1�h�|2�O�WھŘ�>D�x�턷-Y��@Љ
4}b�CQ,?D��(��5BB���e*T#*H��Z�j#D��oB�6L11$�aEr�a� D�,��ֲ!�h�Dɟ/r�H9r�L?D���%HiӞ�H���%�|4�#D���!m�"{��|�P�ǭQ�h�ypA$D�i%m�.Q�	�B(I>U���Z��&D�p)��0Ql��AbS8!�4:�N$D�ػ��&�։��bN�:fx� �h#D��`�$�gK2 &P��\����>D�|A�Ò���!��P H�С	�$9D��W%�Kά����v���7D�� ]�#��73PP58��ŷN���P�"O�\0�M+��iÈ��e��$)�"Ovu(C��%2�d�S�K�=B8h0"O8�����3p���#.N,Ё�"O\�zǣػ�v�� �X����"O !���|�XAm�:.�����"O<�9�)Hb���X�I�|c�"O��q�ႊOP��*��$o���*�"O���B�@s�c��={�"O���E
��uە�϶�. u"OҴ�@ݏo"��c�e4=�r"OD|�v/��"���������<i�"O��"2�$��D�8<���)�"O���f��l�!O��ɛ�"O���&�M�}��,(` D�2��9�"O�53 �I� z�ܩ/)G�,"O���Ľp]Q0��p昑�Ǉ�P�<1�)�`�d@�'�X񺶭�V�<)��+q������$�@'T�Գ�+�-�p�5"�;F1�9J�a-D��Qf�����(ˁ$�5�7�-D��i�IW X��Y&K#\�`��)D�8k�I\�9��YM!��g�'D���$Ǘq% �cP �5H���c!D�X�t*�SEy#�R8�����@=D�|�«��?clg�К 9��g)9D��	�)B��BG���6}��#��5D��k���V��t�*Bʩ�
7D�T����&-L80�6��7��]A4D��J@��&9��� r N���l2D���5�	_Q���O;9="����3D��PSj[fȁ��H\b蹫T�<D�`K0�L���Ar�b�Z�tS��=D�lHG	P65(|�`g�v��y'�6D�,y�i��~dِ�4��Yy��9D�Њ� R�r�*��H���7D�@�+ &"�v�8���3F0A�� >D�(���7(i���A�=i5}�?D�t!�F�=v��bSІAo��p�;D����ݦg�5����1䨨ǋ%D���@Ҝ\�uz�I]l�D²� D����fL/QW�����.p��q
%D���#J_����6�G\"��L D�h��E�3O���N�T�.�X7M*D�d�5j�}����6k̩]N���&D��͟�P�����15��p�#&D�P2IRF�8�i�']s�H�C�;D�\��#�$
�� 	��Ks�T���%D�H�O�t�ܝ�c�A�+$�D�4##D��(eE�
.$�X�!�'@h۷+<D��ćJ��������:'0�yU'<D�(3�N�MLkF�D ��P��&<D��)�2QYL����1䌈�v�0D��j�+��9$n�4�
|��a1D����J�����[/X�	�Ǝ-D�Ȃ!�آdG�ؐ��4՘����>D�� f��o�:$�U�	j�n���*O����m�|��o��T@��K�"O>���Z=L�LEq�@��cG�-�"O����l̓zϰ���m�J ~z"OR�R� �|�(4���L�^�EH�"O�|��B�Sa��r�F@k���"O�-�ՊL<vQ����@�.�x���"OB�R�)Ӌfj	
v`
�
<�"O� �� i��d�Qx� �J��U��"O���p-Q�1�"�	g���j|-˦"O����iUcP8�N��]"< �"O4�s�!�3C�v|�GL��^$��Ц"ON����:�,��+�a�C"OpQ�TmZ&:���Z�ȑ�6kf�%"O
AP�!^'����"a��2�e"O��0"OR�Q��0Q��b��� "O�i�G�_,wn���$! �b"t�8�"OJ\{�� @�T���À/H4�R"O�1�c,�� ��q��*�<�"O�Ր�F�q�`IU`ɭN��H�"O���2+V7Qn��b ɋo@)�t"O�l�	A[��d�3�;�mj�"O	��KL5�< �EY�\���3*O�JǧE%(}�m�r��
� ti	�'
`ݡsD��sxt�I��� �Xe��'�ƁЃ�E&&� PH�a��vWT|��'~�j�a��26�@��C;|΄�'��U⁄D�<���{�[�$Ef��'��TO��*}-���H4� �'ά�1�(R6��yy��҇��}��'�^�
5;�DAʗ��
H�=2�'ȪA:�Ŝ�θ`1'��xV���5|R a�I9_YHԑ�g:.��هȓm̄��N ^��A�%�&���S>�(�-W� ���4�I�a����ȓz�塥!��l���Q���G>�t�ȓ	���`�.I�M� )	�|$��<���(D�
G�j��u����ȓ�lil�=㌀��$Ì#Ө�ȓH�\���:p��C1$R�:HL��ȓ�E2d'V�4D�|㖪�u�؅�RP>���lԤ/L��
���%�����Y7���BQ�2�2soE��I��&���)�A���apǉ%��ȓh�8���ج_b����Z�~� �ȓ����/͕޺��N�:����ȓ�`Ѐl,*��
؉>��ȓC��RR	�V|���k����l� (��E�-݀@��C�q�(Y�ȓr�֭�G�-X~0$��gY�j�1�ȓ6�8D	�)�4E)
� ��B�%a蕆ȓ<��1s��wJD��b��}|�-�����
��M|i�Y��<�N���'@�m�ϓ(p��B��p_j4C�'�&�)7��@� �*M+!�ک	�'�@���� �
m��I��v���'��@h��[5Tx��U�8м��'uJ)t$��(~�s�%����'K^*��S,~py�Goǋ��M�'���� IKD���g%E-P�0
�'�BY�&䊚~*�z@�;�0d�'8�9$.
��&e�׬��A6�ea�'�-ӓB�
R���hZ,4R�1�'/�����N 8�#Ʉ�s�T���'`��c�g'Ye���@��3ab
�{�'�|}BP��-a����P�P��1
�'O^�r�G �^�	EG�%�
�'x�0�f%�o��-�-=�F�
�'� @��Q�
��3��U�X)*Q
�'Дz��}�2%���P�+|��8�';N5�%�6Q6����''����'ܰy����X�|��	���z���� 8��� ݉^�ȍ�E��1p ��"O�D`��-1�AH�B|z�B�"O���F�6j���ON�h\Hq�G"O!�N�@�8a*3.�>�����`�!	��������㝿b��҄�zS�#>������,U����,�|@!�����6�S�4����~�X�-
�hr�lP���'sўb>ez��ľ�4����(R.���+7?a����)�.Y� ҭ<�~Ti��1��Q����*�$[+7r�Hc�GP�D'�e��H�˓�?Q.Oa�T��=�r�� �;z�l1�2����y�֚pn�X��BR}�㰌�6��'�ўb>u�b�
"ݰ��!#]�	�.�Ð#,?����9��T�T�X�|���Ô0�v�	E�����L�fg
K���
	+[4T��+4��mם5���GQ�d�k �%D�<I7�V�nr �/ۡk>��{A�$�a���Od�-s�W�L�j���"H��O&�=E�4��g�2�'!�%XUr�TE\��y��)�'Yw괺�h>5H�� �z�ԉ��''�ɶ��$#�ĥb�D9������ŏ?�q�D�
:� �6I�\�D�<�(O?�	>��\:I�6}�v �˸�hO>=��OD��9%K� �YdIg��D{���Ś���$LI�	�
E��(&X�=�� ]�����T~�2C�VZT#<����?�)���vn�ex�kנN��uRD/�O8O��Q� �1<m���� �r����|���� �p������5 ��I�SK̭�'��6W�69&��7:B�Irur��w@�@<<Yi2�]�0B�ɑ/d�=(���>6L���a�K�B��!�"O�~�P�i�fЋ *�C䉔IT�!��2o2��-��E�C�I8t��I&��#_�@���މ`^�C�	6}�*Hd�\��Z4�!,�lC�t�l�C�005�q��)2!ZC��k�nm!�N�� p�"8&C�	�-�����3k�
� �"sV C�	&*ŊL���׋ry,�@4/�;]j*B�	�<�v��	ѹ2\�j�E
aB�I�0�+7h̊A��)r�֌)U�C�ɺ�r@���+v[�]��k� h��B�+^q��+Y���BVb_%jӚB�I [i輢wf��R� 
ߢEfB�ɼ[����+W�A�D�Jv��}<*B�	�hn�5�ݟkXD�xg��5��C�4�t;�!�Z���A�eIT�&B�I,��c�E/Mr���#�!30�B�	)E����.F�v�y�E	�{��C��"[��1�-ܕHJ��K[�t�C��
;e�9+�C�;�H80(W�o��C�I
U��*ȝ?2����&���}ۘC䉦Y����gco�!�"�� }dC�I������?z��P@Z� G&C�I'Xr]�kP5AN�(�9��B�|�V�� e��M�L��#vB䉐���r�Iڗ ��
�pU�C�	(� %sǊ�xK�UiJS~�B�I(J������
���Y��.z�B�	�x���d!�3��� �̩-�zB�>i�jȸ6`M�G퀘��ꄠO�B�	��e�`�Y�x)D��"ZB�	yP��J��]�u��0
�jB�ɛj4�0��޶ᠡ�te�6�RB�)� ~������<��i 7�G�}��Hh�"O���w�U;1�P��u�_�)J�K�"O�y�&��;f_6���D��.T�˲"O޼��J�
��7m[�;�%]��yB��@�,�a�Ȧ����j�=�yr߶1�Ѱfdֶ;����S���y�G(A�E��B1�+T�3D(��N
��&"_���Q�ǈ�7g-���ܝ���d<���e5U�\ ��'��a�SD]���T4ZP<��r�p���]�(k��T.{_2L�ȓ<sȨ���Q(tƪeC�$�4ov�0��R�iz��݄8�2��o�2ćȓB����Al��:������Tی]�ȓ��|㳄R,N�V�27��\ԾՅȓD��U�&FP!a��a��+������<�#�vs� ���-N�^���]�кE��a �R�O�%n?�ІȓNK�$�P�< d��R�J�"W���ȓ��{���P`�E�,i�̄�{�L]���ϕ.p��dUTe2��ȓ;���	@��*>FT(	��s�z��J�.�!Ԍ�r���@�V|��M�ȓX�~�%��"���е�L_S���ȓB�L�3�v��(�Uk�>5<p��K�,UjE�۷W8%q�J�2#ڄ��F�r}r̢4)J!i2O�x=~Q��3H���C�T.B *�adK�A�:���t�d����=h��LICH܄P8,x������;��iY���!T�0D�X#Uj� N˼�S�b�IP�q�+2D���LN&b��i 7$k�n�0U�<D���e�
#+�!�U'��&t��P��$D��Rb�ʯt٢�Pu�b�h�v�.D��R�K9$���qe��.-�ġ��!D�,�o�E%�a�3��� �:D��ӁD�pv:ى�Q5wߐC�%D������<�B)z���k*bd���!D���gЋx�JE��*��=9R�K,D�,���'���Z`�`�`��(D�$��OH%Ra��aC��|��P;`�!D�T�D���E(��Rl_@���4�$D�\��&�2��u�qF-=z��fK5D�di�j�V@�ת �t�l 4H3D�(S4�J-k ��c��qKt9U%?D�Tz��I.(�.Uh@܏\���H�i;D�x#�)Q�(�j�:�@�'�1s;D�@c! ��"� ���;W�E�"�.D����QP�I:f��rf$�ZG,D�h�e�>r�\+��ŭl*�R�%D�����,*	��c�bŵ$��y�+$D��R�8Q#���GP�E�-��` D��h�e��Bz����
c��aє'1D��R��ޫ��)����9!bt![^!��Ȩ \� ���� �ʬ`�'D0t!�[>y:^��Kڝ$�XQ	�(�E^!���ta^�*��'�P=a�'K|N!�ѝ7"4��w"��a�(�# �EL�!�=7 >�[&�R'0���G���!�$���!ڤe8�l��$)9S]!��M�S1���O��B�pqS'�/}�!�Ĕ�CܘH�rB�$h��y����T�!�D_5P5f�E�/cz��0j�!�ɶy��郶�խTR��r!�؜h�!�� <m��+�~=BU�M�`H.(��"O��@���w�^��׏���y�e"O�Q�PO�m�4< A�Ag�\�g"O�i�w/��I�6T�b�ÄIl|0R"O&��'��&:bT���2V7@�D"O�$��֫TG�A� ��8Y0xAr"O��Cѫ�h�&�Ц+��""Z�c"ORXbC�¢B��08�8
��A�"O��v�"eӇ*ŵm�
 �"OH��'[�y��H�u,ڡ ����"O$y��Ĝ�)��jS��;�>0s"O>u�� �N�� �-i�Hb�"O���s��Za�ũ��@["O<���!�
����A�'\,��&"O�]�&̷>����ƈl�z@:"O��9�CS'E��	TC�1�2"O�q0N̍4[ڼ�U��7-;�T:�"Of:�j�8ar�� �D85"O>i����/5��b�4~E섒"Ohi��έ}oܨ�'����L��0"O�= Pd��o��`�R<^<�B"O��A�ظ�V���d�.`�m��"O.)ؠ蛺9�(�"�=�t4p�"OP̒G,B�yS4Ea�LD m���� "Oh��C�~}�͑ƥO�:{ Lc�"O,T9a���Whjd�΢l�i�"O~L�3#.eH�I�J��d�=�"O�x�QK~	]�p���e�MI�"O(�Iv�L'4,�`'� ���x�"O� Æ��<>�I�ǙXȰ��1"O"%���%n�`�CdZ ��@!�"O��� �J5y ��Dg ��� "O$��&\�t���K5%E�6p0Y�p"O�����_�\e2�	:;l�ɡe"O��;�Xx	r�J�M��z�q��X�<Y����
�l���dY�s��j�<	'�ԧ7��lK�ێF�p�� `�<�4�V7Q��i���z��q8��QB�<�����ք�dO�S��]8"ȟD�<)�뎒p�*��t��:��Z4L�L�<鱠� ��z"
B��i@�p�<��M�R^<[0X���vj�o�<�c��0=S��[�o����t"U#n�<q�H��R�B.X�6��cF_�<a`�Ȟ6aKt�Ĵx��y��TX�<�c��Gʠ�qf)�-Z���7gC_�<�`\#Hڔi��9T�%�T�<Q5˟� @�`d-Ⱥg\�X�fN�<q6n��5T�1�dML ��a�c�<	��l�*���`�%T �kpI]�<�P��%V���j@�[=Z���Q�V�<�����H{��w~b��p��x�<���=R������!8�)�q�<�W�����2G�Ba � 6̏p�<9�PO�+'Е<hX<?Z�P�"O����(-Y �A�%ŢZ.Vu+@*O�1fM�p&XHam- ��p�
�'�� �Q��i}p�9�K��u�'�:��`L>Lc����K5�~� �'2��ab��%'��iA %��	O��'�Vi�0��Eڭ['[� p���'H"���j�� iND;GG�"%j���'δ���zQ�$�&$���J�p�'7���(A�p(�ö��������� v0QH�s�$�9�59�r�C�"O���C)�bw��H#b��xNM0"O����)�<vv�(G�X|=�-�"O���V��R}�ܑ@*U.t5�y "ON��P&��U���x�V�63��r"O�p�"�T�7�&��(�'I� ؅"Or�� ��/#�Lu�sG������"O lA"N�? �.ei��-���!A"O~ ��V&CF�Ã�)�X��"O��Rw�$=�� DFE" ɨ���"OD$h��.���B�+��9�R"OV���\�G�lL����4[�XD�V"O�-CE�N��渻2�-���"O4�* �(a�l�)�HI P��Q�"OT`��)~դxʱ⟈|�L@ �"O�
�ѐz̠��P�U�7Z�`b"O܉(�iC3}�:|���
[E���"OhA&�*,U������h�HSW"OR�"W��.�P���<q��1�"O��31�ӮZ�����HQNE8B"O��jRb�%E+r(۠2�)�"O�+deG�Ф#�g�*�59�'c�	�4գ0��@Щd���yf_�V��$8&�C)d~فt�(�yB��+/,��t*hyD
���y�(D7B%�xGhY�!,����y���)0�t9� 4t�ȑ3�� �y"aP�A:�p"G��yāѲ�/�y2���5l�A�&G[Y0Mb�T��y��ԗ<�*���ױx��B�2�yrJ�bVe�߈Z޴D�	�y�덧[��AnX�"|�w�y/�x�	��y� ) M��m���?Y�O��~�m��O�,C׆ �2߸�b�݉^�*Qp�i���"��wn�<�K��:G��S�?
P��l��˓G�
A�`����\Rs�D�Mޙ2��-�(Ѹ@�̢	�lP#��)���r�M�֤���y� 
�q�옲�.s,��R���0^v�'�ȱ��� �x�b�'}Ҷi�:�� L^t�Y�aG�H̨Í��*�S�$$
\���b A5jK<8p��Ķ�~2�p���oZG��?!��Wyr���<s�����<A��ɸGCd`R�h�$��d�O�̩Q#�]��D�e�60c�
�bؑL�z�^�0��*tz<YES#Q�8�'@�@5���+R�s"�
���%R��(b�g��Q���y��ަz��SV�;�f�$݃
��v([|H� .UN�x�ǯN,|n�;�&jӂDz��Dn�~a�u �7j� @`��$�@�u�	HX����Gz���#];Z�ҔxA,J	q��F�'�Z6mX���i>%;����M��?��4-��Ya���09[_�~�@т�'��ɛ��'K��'��U(�,^)I�p1"��'{�;	��h6	���ꢇ��_�VE~��Y����#"�T2d��EuN��&!"@}��n#y��� �p�����M#4�i4��u!O�t��b�s	�ś��O��$*�)�x}���7Pt�F�q�QAC̞%�p?I�i z��G�υ<�д3d��3%]���	"~r剕&R<Xxt�K��(�	s�D��(�2�i�����D��a�$��R\��j�H�O��Y�	"i���`v���䘍���ՓV��T���|�]w�"y�/Ȍ`�	�㢇�R��}��O�P� ��N"]S�+q����	��)�J~���DR�������uW	Y}2�ܔ�?���i��7-�O�"}"͒0'R>��R��>�!�1�	A��O��=�N<Q ��}F��r�߮gDn<;�%y�'m6���A%�0�f#AN�Ƀ���;@��L��Ej��	_yB◙#�7�1�X���6���a ��Jt 
37rhoZ(�xMsr�;S�4X��
��$�O!!C�����$Ⱦ^����E)�\I/����ťN�� )�l��9�bU+�^�?�H�O �%Ε�& �i�FP!�E�a���Ҍ*OF�P7X�Pԇ�O��K|�	Ο,�I��m���j.�X���R&1�@	��a���	@���HO��U��]���1��ÑC�0�&�O��nڍ�MS���?����+��+A
w�¼�S��(]��s*�$�9Si�O����O ��ʺ���?y��2L$��ęuaR��#�u
���8R��D � A`�]#��u���R�'|����	�m���㌋�za����.p�x� ų
W �`��
(vm�DG|�'vV���t�? ؐ��H�2S��,���e�3�MC�i�bT����n��?�iq*ͻc�v�"�w��f�!D�lY/�+r��#wi]�Z����̻�`�I
�M���i��O*�D�>��.�< 2  ��     �  �  �   <+  )6  R@  �J  .U  H]  [i  �t  6{  ��  @�  ��  Ȕ  �  K�  ��  ҭ  �  X�  ��  ��  �  ^�  ��  ;�  ��  W�  ��  �  i � � 3 � :! }' �*  Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�� |d��"O
`�(�;���8���-0��1%"Oj4��ND^[��"3/9�0|H�"OB���H��*�ʞRy=a"O�味V�!X��!&F�:J�$���"O,��a
���C�Ą�M�"O,$3%o�-���p���+Ն�:1"O��ݢ1����`���y14]2��i�<�6��{_���c�H�`�fX�$Kn�<��A̼VI�xR[�)�Ć�pඤ�ȓA5��('nߡ4�� �)˩%� ���,��r�؊b#`T�eT09���ȓ!�b��g��}�8�F��-? �ȓ
K|m�ș�VṔ���2�%�ȓ"R�X�j�4JN�1�˘X�i����̹	_�jZ��1!g��zܶ��ȓgil,*�J�
j�Ne��i�J%b���f	�(U��:���G��$Y^م�~r�� S�%T"���k\�jx�ȓ|4�1�îJb��@ӵ�ݩn�V��/[`�"�v4�R�!ʎ<��M�ȓ`:��z�ؚh�J�Z��$HY:	��H��p�m�C1��!��B:��0��EnjZA V;9����J[
2���	��4'J�EA�IVW&��~�(aZ��ӹ�>� o�Y�|�ȓ�f�A�
Ο7�H��M�$�����mޠP����/���ANXo*�ȓTv�����{ ��-7�*h��I��sB�8�8���3����ȓNe*M�悡;������X�o��!�ȓ'lj�#F�m�+R&;�|��2)n�C��0S4���T:
b���:�0!��e֊��)��ͷV��,�ȓ0�&�8#���� ع�L�����;�P�AFd���,w�6d��r�EQ�( �gVlɦ�M,H��I�<��!�]*A2'-l�ĵ���@G�<���%.H]�CV�+J��Hg��A��X�?9Q��;� i�;CO"���	YE�<��)�2tN�P3"��Gp�I���h�<��DD�T�rĮ��w����JN�<ف*'1:j�Q�^;x7��E%D��1MM�)<M9$fǭRu�1�`�!D��SwaT:ir��j'[����2 <D�4Bf@��&��-��I��rޔ 2A"6��y��>�ꅁ�dC�l����F��B�	�7&��)q�ΤW���YC��� ��a��h��H���74���9��<��"O���C�x�P3���b�e�7_���I�}[z��Ì��S�.�@�AiC䉋(K � N�AS@Y�3ϗ??��B�I�:JvԂtc�d�*�� �}DԢ>������zp0�CY:XVƜ� �]
9��6�0�c���S�?񄡢�*�o܊ �N�'Df �$�B���'��dEx���ṃ>����h@��Vɇ�Q3�բ�*�a��fË�x�����*�X9if�_�?�����	VBa��G����ME�c��(q�H��h���Z3��
�͇+M�� ���jч�9���p���;���"צGSx.���f<� �ah�� �D(RR�d�b��`�<� )���׊T�@��t�_�SH��"Oz��1D:z����Z�5+����"OVx{"�x�A%_/!`d8�"O��B�%O~&�q�J�.n���"O��+�H
���%�ѽ8G��`�"O�}�'�M�Ĵz���4G�5"O��i@�]ɐ%���T� ��"O��J��ɓ:]Ss��4��Ԋ�"O�e�f*�E���rWf-q�m��'�qO0 �H��^��(@U�gCx�I�<D��1#*	Rp�y�T ɚ#�h�R&,�Iy���'X�� �gE��l��c�:��m��Eֺ��6��g
���7��{%
Ezr�'�=%��*$�C��1:�ԋ	Ó�O�6��?�0%��jP�T]�E�O�z����$�g?q��V&�&l�voȤXW��{%�l�'L1O�b���A�	.0�(Ȉ��V�<�3E��7�y��'P�Q�"�N�	���@�H3��ܸ��Y��G{Zw|F����}�5�oE�z��9��'Ȑ f��6���˔}QfLш�'�xp�hY<l��Qo	f�6��S�'��O�%�mء,��5i�|��x�'�#=E���CR|$i` V�Af�9��AY`�d,�OP��>�:� T � P�aR��'�1O�d�T�F�ct읓O�h3d"O�4*�ҏ�,���k��E������$�S�IۖHn��$�D?���i�l��+!�ߌ5͞�rPI�oӨ!�KZ�p!�d�{��8�ʞ�@ ���f\!���rZp�f�
<f���I��O�!���A���E,��C���E�H�!�D �#J\�3C+�5,(�YaDL�x��}R��83F$�*�i�@�(WhH{n3��e���S�0��p�i�����䂼j8C�.���8��T�Q�10�C��A셭�8������+B�PZ��hO?٣��=Ql���A�$.m��q�UE�<�v�D�kȾ�AsEϋd��u%H�~��4�<�gҪ%�H�cI��p��٫�)�wx�P�)O�����Xi�l1a MPrl���d>�S�i��l=*�j��[��\ʦ�O��Py�:�fM�� F�t�GIM���<���$��C���p��-���0����x�!��8���R�jĞa\l�vo�:}�Ib����j��n1~(���
%_��!V�-�O��O�	� ̻{+R����	=�l�fo�O?A�����T]��|ZgEŷi-cF눇��$�2�Mc�<i0��qc��P��E��m1A�T^�<Q#+W�k��P����6D}R��$�
s?������� [��Q�i����09��d���d,�$(�9H9�G����t����Ci ���Iߟ��u���:!@q�ȅzf镉$�6��'ra~��dv�����ΌO|ty鱈^���OTO��O����pN��7�u��戏Ģh�
�'>�$-G'U
9�1.U!��و��)�t�ʭx?Lj��]�Vd
��E2�yB��,~0��XQ�?��5���y���2M'���A-C�Ԑ�36�p<�.O�O���B���1�z|b]�w�(��"O,yz�b�(!#��J�&�0������'ω���4TlC[�R`	���8t��"O$��!��A����`(S�/�ppx "O"L��^L���!Dn�Y��"O`��#jM%��p�_3>���I�"O� 2��� ��Y�`�#�:a�p����J�O�y��Jވ�B�C(מRqN]��'<:� ��)V=��#!i	Ϥ�-O��Ez���pp�4� *W��.�!�$�
:@�:wE��x#f��w�_�5����?+OEGb�Z�X��9��$���ҊU��0?y�X��L]�zٚ��AV��0��%D����
D�r$�wn�\��Ţb�"��hO�� N�,@����!|m`��1�U3w�B䉁S�0Bd�_0��6T�G5��F{J?���I'C��K�Mߐ\}J�#P	6D��9D�@62�H�)W�
��W���<�}��9O
��oGq�P�E�o`٩�"O��q$�׵B b��6i�+~d���ī����8�	{�'"�Q�`_�T�l��O�
6,��O`㟼����$��t1����5�LT`ӣ�G�����)D��:ť��b9b<�4�1�^9�$�+މ'U����E�	����
҂��m<�����n��:�D@fdj�*�-�DM�%�:���x�	�h���O���z��Z��F1c!>4�@�r��(Oj�[�G��UZ�jI�0Ȫ|�����x��P�NܰǪ�>:t�fD[���?�Q�>�˟�aX>�յc�D�H�A�y� �ȓG^�b�-����W�+,rP�{A�-��ګ�0=ْCR�_1XQ���K"pX<Ta!��m(<�شan��R�� ���	�X۔��=ѝ'��x���P@� !@_3$8��r�+"��?�'��a�4���pL��8"���||:8c�'��1�H �hO�����m
���'�
�27(�D��aGb��g_ A
�'B��{���(��E�g�Y:\~�9��'�4�¢��S˂@4���M�X	�'��pҗ �{�˂�1&F ��'�^�*�#��C��L �D�#U#|�Y�'�޹z��͇˥?�δ
��x�<��"V4�ܔ��<9}���c��s�<��G5*�0  a�NBG���dMXY�<y�G�{���*Gobi�tb�^�<����(��@K���" M��P�CE�<�sÖgdPI���Y��.���[�<�P��>�Iw��64He8��X�<�ce�V[2��!�WK�ۣ#p�<a7��l�Y����L���"o`�<�F3} �X�r@ݺ4��	)AdRG�<�X�9�r�Z#��33�0��'_�<!����E S��UB�ДF�Y�<a�M$O�lA�e� B�YP͉W�<I���0�ZG�7ݔ�;!�AW�<�sl�>O(Ii�C=e��Y�m�O�<�`2/
N�KMŲ^��x��w�<�pG��E�2l�PoG�t��p� ��H�<7�߬)��I�'��P`��
��FA�<�mܪG�~�h�B��~p``�I|�<��I�5?����ݺs�j$ꅏ
u�<��i/H��,Z2JR�#L�P��G�<)�#�obaq+[�M{�����{�<y���:}����S��+�H�O�<����r�>`b�)GHP����o�<�NSs��Q��焏��(Q@��Q�<1�V)5�}굃�`��	1���d�<!���WP��(�T����%oY�<��̀![�����mv� ��R�<ǌ:crJ��̚� ���\M�<�5�C�wO��%d  9�ɐ�q�<� 
`OP({�NT*���G� (�4"OƜ:�"B�a�@�@�'���U"OU����^�9�B��7�P��F"OR����!zѲX�FV�|���"O칫���Ί9Z���8����G�'�r�'�B�'���'�r�'���'�l"�j�8f*� "�ᜳ`�g�'���'8"�'���'i�'Hb�'��`0��Az3�$Ce�T�ij��'�"�'\��'���'�R�'p"�'��|`gJtEp�J�iŪ,ˢ��f�'U��'��'���'B�'���'1�����TVZ�H,�>'�n=[�'���'���'�2�'O��'�R�'���z0�+%�JcP�7�"E���'��'�b�'���'���'��'Ƭ]��e8�~� c���+C�+��'R�'b��'���'�R�'���'u|�k��#�	
w%2���`�'c2�'z��'���'���'r�' {7E^�E����$���8�Br�'}b�'`R�'���'�b�'��'��:@		/h��@7��7m��A7�'���'���'���'R�'���'�UA���<-�:6� w�P���'��'�"�'���'R�'}�'��	�䂨L`P��C��}��;w�'_��'O��'��'v"�'��'QB5��L��)��$J�<�U�7�'�2�';"�'�'P�jӮ�D�O�p�q�e�pQic�^�r}�UӏZGyR�'��)�3?�ѱi�쭣!��c��u��&+��H���^$���榭�Is�i>�I��McR�g�Ԭ[�H�9!+� Qh�cd���'M�Qĵi(��O�RFn�!�������HЧ��� 1z
���EwLd��N9�Iݟ`�'k�>�ñ˻��=�-U*(�$���ٳ�M����y���O�H6=�"�q���%D��0�7�]4wN%�v*ئy�ܴ�y2]�b>9�d�M���\ܣ�%��'� ���DE7(V���^25��OÆIH�t���4�
���MY�l�����]
�L�ʂ���d�<YK>�C�i�C�yB���P���c��,��[įϗH��O��'��7���̓��D�p�<�0)��v\����S��:M����e��b>Q�3e�ٺ���'� :u�C�#r,L�R�ؚ7���2[�̕'���9O�|�P�U%'�\*�I�YL���2O�nZ�K_��c�v�4�Rm�'A�$c}�ŉ'��I��"�1O$Ln�	�MS�N\@�4����&-rv�U7V�țSjǵ_��ɂ�ʞ���TG!ѐ�r��
Tx�鑉�'Ei@�P�L"q�Tp  �� �����E/��ġ�$s�����D}�)�� Jv�`J�(y���rPm��\�t�bu�ɵ �t��B(������և{y[@��/�2,�!Ϝ�G�XX7����4}�s�ſ ƴI�eӍo7f����Q5��y�p��aWhd��M�d�p���n��3�p�D�e��Y��E�[��M8ĻGO�p� DqmR^���djW����#�Qyx�0Q�I�r܎��c'��7�7��O$���O���矬����$X8�{�Q;~)���@#)x&h�'q�D�sb�'�i>��H�R��h
�)@�ވYuH��$�i��5�R a�Z�d�O<�D�����O����O���mݩy�Q�S��#���Zf� ͦ-9f�㟰�'���1�O��O?��T�2�p�T	�+W���uC�%^��6�O:���OV-�5��ߦ���ڟX�����i�	�bB3��]	C��5,�\�iWm�J�O䀩W9O�Sߟ,�I���P#R�}��%���#[�F)ڂ���M���*��@�S�i�"�'�B�'dj��~�jU1w>��S��MJ�ʧ�Ŵ��D�5=�1O����ON�$�<��ɲp*�1�d�,~x���֥��ːR�D�'N�P�@����<��'p�i�)3M����̚'��z���Iܟ��I��t�	i��k����6MH;�`���M4v�.����$0	o�џ���ݟ|�I��'w������+�S��R�-٬&踬�+�yG7M�O����OJ���c�$�&! �6-�O��dK�B�8�d��&Z��S�F��kf�oZ�����ßt�'��������'���̃=&1�r�F�(�d�c�X�YΛ��'F�'cb�� �(6M�O��d�O��i�2�)�P��x�Y��%T$!J¥m�,�'�2�������'��i>7�W}�3w�!������[����'��/��5q�6M�O����O��)�V���S�.�Y���ŀxZ .W�378�'��Zl���'�i>ᦟ�h�fd �H�NQ8�J��x�F��u�i���Cu�z�$�Ol������O���O�Ir�U?u@RlC'v�=�v������Lʟ����h�go>�$?q�s�a��\��P�$r�tH	&K����	ǟ`��3|I�t�ߴ�?Q���?y���?�;k�يE��5s7�)H@0n��Д'3�@Ҙ��I�O0�D�O����O�5ܱ�sD�8@ �A�D������JT�h ߴ�?����?����K?� hۻ0���
}�����z}�h���y��'�"�'�ґ�t��9g�@���V<<�H��4��*<�9dd�|��O���O���O��	ן��wˋ�U�j�w��3.��Į�p����?Y��?9��?��&��� �i'Vq��/�LV�*�B�d ��af{����O���O����<���VH�'~�^,�3�I?q�d��C�Ós`�Q��ir�cCcSR�'��I�6d�E�O|�3�Hf��Q��a��(�pt+�� � ԛ��'��'@�I/l�Lb��r�-������6f� �B�d�����O��R(��!����'���/�!f:шH�(���A[1a�RO�pd�yDx��� ����~o���R�G8,����i�剆S�� ��4#(����� ��d�-k.I�����p���kŃO
�v]���d/$�S�'v�40!��7N�X�[�.$��o͂��4�?I��?���e߉'�	6E0�)���u���rÖ9D`�7-�6Z�"|"���<c���a��a�R킥>�HM;��i2"�'_�	T#npc�d��K?�p/Z�BL�7E�.UNRm��"�i�n%�)�<��?Y�h%,��)��R�$ݠRkI�>���p��iX$�.�lO��$�Ox�Ok�ѐ$U>�iB͠J��q;u�^�tz���2itc���I����iy�b�ET�E�?z��=�2h�?�(\(t-%��O���>�$�<��EחI1㔀\�N�3,J��,)�<9��?�����@-<��e�'6����uN̡X֝ۢL�|��8�'a��':�'`��2C\����j��0<Ֆ����ʚp(z�'�B�'d�S�L�Eۨ��'r�P�J��$��H�JF����i���|�Q�����7����v� �$�#L�a���mo�6�O���<yAc�5��O��O�v��1�Ζ><�)��W'e� �Ң$�d�<Y��L����[1Rt���U�j���0�Ĭ65�VZ�X��/�!�M�RS?����?9��O�hY��I�Q2�ɛ��i�p�i��I��"<�~J��H;,��@�@)=�L��c�����1����M����?q���7�x��'
 u#�/0�$L�2Jэ@��S��~�%L�"|J��l*0�Ѩ�4��h�g�O2���i~��'����Z�O�D�O����3GBm:�H�z���x� G>~��c�|�t0�I��$���	��Rt��a�I
O��)	Ԇû�M�pK~	יxr�'`�|Zcu>��&��V�p��E�m�xa��OP,"3��Ov�$�O���f�!&�c����%�B�a�E�2ya�'"�'��'�I6 -�����&v���E�S�"D����@6�I��(��̟d�'�f�ѶEg>�SJ W<D���ߞP�`C�A$�d�O��O��@�	�'�F�dX�MiZ	݌��$"�O��D�O���<I��W�O��s��NV���%��:����Fi�8�>���<��j�q�_X�ʂ(��4�vI��o}��l�ß���ny�n�(�z�l�$���
�M�n˘Q$��&b_:���d�r�Uy��1�O�Ӧ	������b�.��7٧o�6-�<!ӌ�*˛�-�~r��ꄜ�4+�Y7���+P P�P��oӒ˓��aFx�����sL�܃��0�D�s���MK׫̔3���'��'���&�I�s:�J��/�T1�2$��FM�Ip�4XלGx����O�G�H�7�����5���BOڦE�I������=�^�RK<!��?��(���AfY�>�\��SBx���"�d��j�<q���?���d2�	3U�X����Ԑu"��i`R��3��c����򟠔�5f%X5M������{	�qv����-�1O����O����<�L�H@�臤�K=P� �
��+�V��2�x"�'���'���pyR���q�=HHR(l`L����Y��L[�y2�'���'��	�~�x�ЛO��u�a$��p� ��Ɯ)8|�(:�OZ��O�OX� �t,�'~@�1+�0f�TP��
|�&��O���O:���<9b	F�~��On��+B�K%���	#��eD�]r�.}�(�1�$�<��DZ�j0���g��Ir�;�d�l����Ity���a^�8����R� 7g��O�`0�ܞ>%�q�v�q�yyBHŵ�O�өm�P��`�<SK��:�Fc��6��<��>5�6-�~r���e��hs������BR�m�@��e�V˓|�vFx����2.�t��`N�$SvЖ0}?8Ml�j��4�?����?��'G�'�B�K�H�T$��~��cv�^��7m�1M��"|*��h �Q�I�Bf}�A����Z��i%��'>���WrOv�$�OF��-+3�p@�b
���`_�:I�c�����/��ɟ@��ڟ��M��m)����/	��09V$Π�M���?����x��'�r�|Zc|2͈Ǭ��ds^Y��I�*$�`Գ�O��" �D�O�D�OV˓'�,�1Pd"UO@Ӡ�=��j�FgF�O���=�d�<	�&_�3	sbE�:W������ۚ�ll�<���?y����>}d��'�J0��!|���FK�8���%����F�IHyr#]���dC�=�ޖ��aԮ�I �H�O�D�O���<�6A N��OzDYi#�ŚSV,�Sh�O��ܢ�o���d.��<If�X�Spf��0��Y����ҕ���mZ�����by�(O�?���(���&��C肭d�`��fD�U�4��Z�DyR�P*�O��"w��J��&"gl����<�7M�<�a��\�VM�~����:���X��n϶	V�V�Y�u��<�D�`���B�VUFx��$�X�^B�rb:Y�x����M[� ��;M�f�'���'����)���O�l�^�4ـQ��a�N(����ɪ�n2�S�O�b,� R�����;���VMO�J��}(v�i�r�'���Y5�O��$�OZ��"k��%r3�R�n�H�:R�WPl*����O��d�O�}GB;^���rC
r��I��N�M��Hwph�I<����?�M>�1/~���
̙k� �IU�`�eF~2�'6��'��	TIf8A�*|��UC��\"R�񆇡�ē�?9�����IR(r\{�&�,�T�;��S> {�c�4�Iџ��IZy")ѷ'���S�����d����4���O�kݢ듡?������(O>��)��81�H �R~�(X��[�H��ʟ���VyҀ�(��Fd�4������uNԯP��
}b�nZ��%����	-�u f",vHe���q%7��O��<ѣIR�vىO�b�O%��p��N��@�o��>�D���3�d?�O̐�k�N2H��sB��n���_�,Q�]��Mcd[?a���?%!�O�u��AUgp�Q�U3���R�i���'��}�W�4��'�*qS��>@jhH�2i� ��޴}���1�i��'u��O� O��ē����ވ$�@!
ܕLu�k�4 ��D���Ϙ'��`���R�PU)T�z�)2���h6��O(���O.�1��M�����	ϟ�JA��Gvj��`޺&Lx�cq�ԭ��'�%�y��'2b�'V��3H��`S�qƮǿr>�r�����U54�(��>y�����K���7R%b�a3���%�`.}}�����'��'f�X��ҥ��+gh�2�H$�081��'=a2]�I<a���?9J>i��?��K�� +ʉ)���Ԫ=��	9w����$�O��D�O��\��|�D7�dDp�*�)h��5��,�f�j�X�[�\���p'�X���� ��ҟ�c� K/�y���O�\JD�3@�)��d�O���OJ�94lĭF�S/%��2h�'.����mt}Hݴ�?yL>���?��Ʌ�<9K��u�7+��a�A�PK����q�J�D�Ojʓ�^��ו���'��t����<ժ�GKn%H)�E�A9"DOH���O6�	C��O��O�;">lBt�"�D]8u�$��V�i�I�c<Pͺ�4L��S�����$��n�F0sE�o�"Y��S����'g�/ҡ�yZ�"}��삅}צݨ@��8þ��Fݦ����M����o̟��ӻ�ē�?�`a�"	��
Ѥ�(�0�(�^�����y�|��i�OJ4����'x��g�%2B�Y�Rgڦ��I��x�	�?s�[K<����?��':mz'f� <�<9$& hd���ݴ��nm�]�S���'���'������@XG��|���hӺ���P�}%�h�I��p'��،$�4+�c�Rj����}���Ghi�����O8�d�Or�M�$�-)X��ǨE�7�0��C�=#�ļ�I<Y���?�M>Q��?Y.D��'#T�;� �a��;T�Q����d�O��D�O�˓4�T}�t5���JSc�-x������M^D�x�x��'��'���'u��S��'kj�2ve��K�ʨx�IT�N��0%�>	��?Y����d� ��&>QY�@��X�0lU�K�z�S  .�MC����?I�le�Q�����<YQD�I�/ĭ}�L=���'O[ 7m�O��$�<���Z�\��O���OAD�a�K h��3pf�&ꢈ;d�1���O���������7�T?}R�*�/��(�S�T���Au/o�T�#��h�i���'�?����Ɍ,��u%��o�`y��eX$�6��O��$�M��D$��i��s֮�T�ry���W�I���҆-͔@��ȁ'gX
m%�l��C��q�������I:%)d�G�$gk��,4P�5)s�2a���e�:*�)��C��C��f ���-ӞM�Q���28��H!��� �jP�pnߙ9B����^PhkQ. ���Т�� P�;u�,Fz���.˚k�H���Y.�2%�s��lQ񥗒)	 @S��8~
}QF��CFYy1RK�a���T��i�֏�����JF|u�A���?����?)��F���Of��(D�ޖ"�n��GA9̞�� �E�C֠�L,9�����'u����jޭu��А�
�?9���Q!ϥ>�@s�I!|O�L꓃��*��W����M��N�=ro.�O��X$�J���ś �˥Mn~��P�'X�'=(��M���E��
23y��yB"}�d�OvU�����Iٟ  A��3����1̉�w��@����֟`�I�/��x�Iǟ��I"��Y�)��M����eQ4��gUD����6X�$�U�D���O��kեV) ����K$.�@hƫٟ`�04��E$?_�`�%R��BY0���8k6zAj�{�F���?��i�v7��O��Ƀ��?c1�܋�ᚌb*����<�۴��O���I�P:����<��aɌ�1�az��'r�I��M3F�K�syL�����=?q����C+��V��(F�)N�p5���@�O �=���'����%&ZR���ض,��Q���'"ƃYUB�T>�aJ�h�t�	~F�Ps�NDI�O�0��)��9y�4���J�k䠋�Hn��':���z�ɧ�O�(@�)�E�~��c� �j@��	�'ה���F�pP�9��ȏ)*4d�	ÓHU��� p�6!Ԝe���P-g@Xӷ��`}��'��(3\Ԙ�r��'�r�'��w�$�K���
�d���F8!Oйi���� 8����O�<�a��V�1��'��q����&m{r�s��6}�t�"a��|�lݛU��O��r���7����P�ڴ���L
)�p}��"�"&�p͛����ą El�O�ў���n8]�x�'ŉJ�ش�%�>D�Ļe陋y#R��� C $zK�=8��Ƀ�HO�	�OR˓4�����A4j񒕰1�T���&B�
�p���?!���?Iŷ���O��?���܂x�z�3u` �GO0�!��4���oϒ,�䜰�G#�%A�Ĝ�Q�>B�	�.�8��C^�m�`=HB�A A9�u��
�OPl��	�d�X����{���'��&C�ɖ7!{q�W�7sNi�"�ޏ{�Xb��K�}��4|�P7��O����e݆�@ë��`�z�qd���` �d�O�iە��O���|>�9 ���MѤ)gO��V X�Y��%7�%��@�7tZy�7O���A`���	0��h�Ț�O�����)��p�1b�LH-I�qd���
�_�<�U����'�݊�zK�'Fx &�T 	X�x!n	ϺaP�'�d�3��������	�2���'*�7�6v��1A�I�)��jAL#���Od!�1D�]����ДO��i�d�'iڄ�����R�Ȇ	߉M�
	{4�'9"��Z��M٤*ݫG4�'ד++
�����IR��t�ӆ���g������s��<�D9�W��-���#���7N��mi���C��ZPI>]��늨ZajQ���� @��@�
,}2ï�?���|���ބ	3V=���þQ)�T@S'Q!�y�EC1SF�"�G��M�X���	�0<��I5:I:ic�أ\"�&��t�"4��4�?i���?a���f@x��?1��?ͻ+($BEW�o���AA�܆6��1�r$�:T����tԁ 	��1�I+��Og(�'���;V�� ]8�u��@�@�QH�R�L��E��)(D)����>=�M?E�AfE-8B�.γ|�v���Ge�U3�*�. �D�O��d�3����Y������&�9GJ��o����E�O��Ɠ�h�{C��*N�[��~|D��'��#=��'�?�+ORu{,N&e���m`D�8�g7��ᰁF�O��d�O��Ӻ��?�O�� 㒭H6F�4��!�ϋ~j�Y�ԣ��x�IE-S*��;��H� .`�H�,�z8���'-��3CN1���X�h̤U��P���9�?9��'��E0�J��:������1>$��'F�G�Ul"�;s�U(|�Xy�N*�ɝ<�����4�?���g3�캗ʇN2��&#��Ko�����?I3���?������ s���兕�wz����5~���X���"t92o&S����0�)�0Rׇę]�H��s&P-]�\Jc�I۴TSڕ�(Z���-�Zl�-E�53F��ɖ"�O��d�<�(�J�@��"<a�C#��<����?����Ӻ3쒅B톷~�e��ֲe$!�Ŧ��@	c���bTI!+���C�H�'�����*h�|���O�˧|VM��*=�H��c�l|��P��^;FۀY���?A�C��&5c6�4�T>5�O������/Bب�����n��sH�X�F&ל6���"� `�O�NC�(S��C/Cy 
M���'&�OJUl��M����O�xQR�ǐ�,)��M� ���b�y��'��y�Dݗj��LI��]�!5Υ+P+��0<�I/YN���5v(�u��<�Θ��4�?q��?�`ML bF�J��?Q���?��;1�� y� ��q`v��
�jX9�Ju��� �	�R�z��I����O��'h�0aDL�	��Y(���:�f��b`�q�4 c��k	H]�0*Hn�hg+�|Z��i3T�̻g��K @A�ezP�N�+D��b�|���+�?�}&��S�HL:!ԹRĆ�%�*��6�"D�X:��^"�p�H]:w�ܴ8p!b�d����HO�	=�D
0AK��!KA�6���Ԇ�`B0,����O ���O�Ю;�?q�����!k���v+�=��0��9y��3	�',"\���5_� ��Q��zW���x�h�� ��X#�!F�X����J#j���*��1saʐ�`U���2M�
MNLI񯇅�y�lY�T��@	 �:����^̘'/b�hyTč�M���?�c"���b1�2-�u1&NW,�?��l�����?!�O�Yc��T�;W6� Y��p���d�}�ҭ��J�QI4O�J���oиB"�>�3O�kyr�0�ѡ �( b�a8���"�OZn���dq�r���O�>|���IL��O���3�)�'K�zI��-�hg��� ںn߬	���4<�&`��z�hiâ��/Z��a��?�yR^���3	��MK���?�-�4e!4�O� L��Z8,)���K�M�֏�Ol��S�j36!��dP�{��Ŕ��I�|2��N1z��q�bf�P�e
R��).�̅�!�Y-��e� F�k���"*0�	��_��t��	�?"�.����[,��|@�M�	���S��a7p�� n�T�J�0�:w�8��.Ud��d^[��|իE�r0�ቷ�HOu �#\�*:Z+B.ђX��J�$Ǧ����|�ɕ����mF����I���iޱ���2e���4�-9�����AƜµ끚��p��H��h���%?�.���8c���iB��MJ� GX1�~@2׌���(�5�JVoZ�q�oḑaZ-X�Oi�=���ԩj��1�$�"�P!k���(�M��]�� ���Oq���'�	T<E�,���T��B+u���v��'��{2F+zL�1�(�u�d!�s�ǃ�����e��4���|��'���J,l@vݚCƛ�Y8���kW>=��4xÃ�i����O�d�ODٮ;�?������H�aX�ݢu��&(l�9�/|f���~�����B�2�,R�2(Naat�ɇq�n�hFA��R���G�0E����DfZ�q+�œ�+αZ'�*k��E�ɎS4x�d$�1�@u0g �.ypd(,%��#�Op����:�fEIm�3^eˢ"O�E@R&A�k¨@���,<VX����DӦ�$�Ȉ�i������O����Ǧ2J\���?.D�a���OP�Dޟ�@�$�O�28:MX��&>�x�ݲg��}CI	�,,��"�ʔ�Yb�]BW�5O���r�D��M��"*�La�LV-+U��(�o�L���B"�V��ax�D1�?	��i�`�:�P�N��NP���b���+��<	����<�PN�A4���� �b�c"Ne<A��i�l-�d�\�0���Q�h	r]B�9�'��	�0���޴�?����)(�0�<�p�b���
#��C����O�l���/���w�Gy*�X�'/5j,ڱ)�)�8!!�].Ӡ9�O��#ED��o( �Z�#+����:V����oI�39䕤O��E�'�p�O�mc�H$�D0a��q�NQ#�"O�,�wl��"-ȥ
R,��$��L+q�.��|�鉉V^�e�&ꅔ0�04 A 90���`ݴ�?���?AVc@?M�H����?i��?�;:\$R�@��J}�D #�ȰXdYi�yRū��<��ß�\����=l�g�\�,Y.��+:�4��փ P��J7 �˨̱K>qw ɟ�>�OpmF#O�N	N�RT,��d�[0"O-"S$�$\Zt90"� w��V������S9^�~�j&�����v!/�^̸��U \( �I�����ȟ�b^w2�'��	B!ab�U�� `G�}��l�<wN|4�aO�YЖ�7N����ڑ ���)�!�D6N R��ЊI��$��˚�i�l�E�']���DѰ=# �� -\(bO:1���@!�Ċ4!��)�d& *VF	x�`��1O���>QA�Ȃ"����'Z_����b�2�ޞD��1�	ϟ|���ß��	�|2��>X�� C�����TN�@��.
�j�)f�̂0��x���&��0�4"�8g�I�Kr�h	4�ȴt�6 v)·CA^��J�\�	��ē�h���ȪH���sDX^>��+M������=��ũp�EʡFx��i>��ݴ2�0�h�F֎ >1���Z�"K>!Ҩیڛ��'HRV>izuM�۟h�����E�PE�'e�8%��*���Ʌv>l��	B�S��OZp� ��a��q��,�^�*��>)D�l���Obvt+�!��E9���n�,oݬ�J�<I!j�O�\%��?-J�&t��$�7l�|H��ҶI$D����^�⃎+M�fI�m!O>�Gz��f�X������X�� s�7��O��d�O�D	�o8��D�O����O�N˜�8��G��:K�9��ʹnt��+O1^;�$X��8��Ge+��DV�����Dn#K6�d`��*A�Bs	�~��0�ggעBv�: �f�ӿvq64�6��Qx��ŷ:{{�o͏}��Z�J�Ŧqiܴ�?a�C�?�}�'��@Z*�B<�S��c<vqg�$[(��',��˟���'ߜ�� 5)�.��\�t�2�r�O�0l�M+N>t��?�'��%�3�̈́*�TK��$�L8puԕ>w4����'�'���mݍ�	ǟ�Χs8"4��F��jP6���
 =�� �e	R:J�ɓ7b��i�d �0NC:o�L��Y�b%��^��� �&P�ܹ�iQ�>�H��QK�O��I�a�ލ��4)K��OН�	I+M
���L�4պX�B&ۃ:���-�O6雰nջT�љC&L69�X��'i�'���� ̦%L}����+[V�C�yrG}Ӵ�O`�a���z���'&��`dG�T�0`cV ��d����'f�'ը`	b�'�	�c1;��ԇ!Ĭ0�f��� ����d"�1��ڹ�%�')N��w%A�s;���� ��?q6�]U�2@��'3��,[R8���T��O��lZ��ě�d�����y��lz@ŉ~01O��d(<O��C���% L�dp����&�0	"��g����`���wŏ�c $y�A�%wy��$=O"ʓ0�z��p�i���'T�#�-��V����(J��Q�͔V*����ҟ�0^WT�I�#�
X�{G2O�T��Jݑ@Ġ���o8��n���I%;���p��r��9r��%�'�RI�� ۃq���gG�8""ɦO��1�'�
6MPu�z�S>��ƦT�u6�ضiY��c�@��Cx�LSa!ā5��pXTI�S�`�ƅDu�����2�gy�11 !�	0��P�v���*�8	y��i��'���[�L	r�'N��'�r�w�xU�q��C� �@�Z!G���M[�=&��#ׯ 7}�9:�� �1� ��O$$
��֪R*��q)W< ��9�p�ϻ`@�1c�dе�U�r)�$�d�Ħv�D��L���ϻJ���b􄘛B�l�i�2X�8���i�ʓG��I�i>���J��`�-P��%:	0�����ԡs&n�R�����ڵ�'[�"=ͧ�?�*O�ȑ�˗ 8S�CGB{�`%� +��J��S�E�O����O�����3���?�O��+ti�;>��4,Nj���V-ʂz�PB �Ϋw��{��غUM���c�]�ʜ��Ϛ�1�� �&b��*\�1��� 9�f9:�
��1���4\٨ro�0]�J��#M��hP�47W��'��Ο�?�S��
��˦
L��XЬ�O�<Q0�;+�z8 O��6��aY��M̓EJ�aQ����~�-�OZ,U#f���ȳ���v!�h�O��I���'�����'��>�D-�@��Cf�1��&y��ʙ� �v(ͼ��4bG/:Ѧ���2��O�`U#ۼ"����pɛ�8�����Wx�Ub�lŬd} t!P�F�Yjd����,5��et�6�')�kU�[=�6�b��*WJ���yr�'�y�bQ	���b �BJ�YY���'�xB�n����,�F>�ȳߨ^6Msw*�O~�k������i�"�'� w�T�� *��K[�	��#��>�~5���乲"�O�X� h:}*�6�'pFdI௚�wȡ��D0��OHP"4� Ţ��'�thR��ש,gNq��чY�P�OȔ���'�7��d�SR�E���xrk��13>�;AR|(b�t�	Kx������t���u.�-:��+&OrYDz���z�p�7��`sJ���* 

7��O �$�O�0@p�<��d�O&���O$���	M�<�g�+C��(*V�U� c�$AרJ(J��{�mG*Uٖe�'�Ss�I
!-\dq%�-ˀ��4��N]� �a�i�b�"CT�)�8a�Nś.#�t���q ᣓ
�yǧ�B~�0�ȑ���ܓ �O�=w(�O�̓`���D��¶7K�I����r�d��Or��gO	|`�`���u��u��?9��i>&����f�?��9�ʊ�m��8gɌ(���[��Qޟ���ڟ�����u'�'��0��h�ЏȎP���DV�.:�9�I��4������j ����A?<Oȑ��.c��(���"t�i��R9HmJ�(���� iA/U�Q�҄9ړe�R(E&<:�z�Z��X8t�����<�� �0��G
20�@C�#Y��:��ȓP0�V�@��AH�u���<ᶷi(�'s��ULo�D�D�O<���!�
xaL���G\���%�Or�Dý%�L���O��O��àu\ ��'	�Iq�h���AW�����5nέ0&����O�ۡ	ߤs��`(�(�`�Ӯ�(��D��ڵP�
����P�����F$p:j���{"�8�?�C�x�Jno<`�WEV�jx�Y)�.J&�y�J�V�`A+ʓ:0hn|H�f(�x�#uӮ��BDw�lU��W���y�*�䊏G���m�ןD��b�DN�~Z�k��\k�'	�d�F@H��I�q���'k�a%��|fZ43d�]�>�T>)�O+�1
W�����FP��XN�p�gޔ ���x�j�9+"Z=E�dG8O��1�
%-�-��ڭ���KZ��$��y�J|RI~�"lK?`�e�W͌D�P*�ʂc̓�?�ϓDБ@ ����zh���F%��ɽ�HO����z�dQ� D�6�@�E�ئ��Iş���[#������� �IП<����%��.��	狊�+9�d;t�l�^%Z3��
KǨ��B�C�p!�|�`�>ـ U�|&�7LʑjЄ�! A�:n}�$�#E�V�oH0f��ر��EU�ӥ�M� �h�-{W �/�.�A��Z^j�]�A<��]n�M�)�3�D�H~ε�d�̪P�.����1H�!��̫=�jq!��הY־I�a�E��O��Fz�O��'��E`sEO�?�mQ&GۀN�����Y=(��\���'jb�'��do��Iٟ�ΧN�|�r�c�ʔ��S��xVص���5q$���L]��@�tm��p��� <"�۟z�aC�	���S�.��3V(�Y�&ɕF��q� ��{0�քv�$��k0ܞ�h9�� ?_L8�!$��s���D_֦�H<����?��"�&y�<�2UN	&OjA9�GJ �y2"��M�A
E)� �����=��'YH7-�O:�g+ȥ�R�ir�'-,K%�0%�;1�'��@s�'A(�&��'�Iޗ���B���Ha �'	��wN	1\p\A�`c��(�v��
Ǔ��	�o˕;z����ߟ�0H^�=�"�3w�B������(O�D�@�'c6m�䦵�I�au�ђ�cϔ(�(�
Sg�, |ؖ'A���,�h�uTJ�@���HFDB�I��M�s�G	f�*�+�Ea��Y�uh��<*ODѢɗ������O6˧)7�؋���^4	��Q��摱C�@
��I����?��kP�A���M|~rQ>U�O/��"���,@ʡ���g
}sI�h��d�h��� H;5\`8�ǖyUJmPJ?9	1�m¬X��ٛo�X�P�"}�䝳�?���io���'�'��Dś�t�- ����uۜ�[��ϸ��'����?�$G�%t����� [�x-�2#͙P�axRp�0l�����4�?��hL~��e �r���CTOF=*���'�'��=�O�*�r�'�"�'L� �?
w��U��'6��.�k|~5�K� a�iR1d�b>�Op�Ca�.������ѵ-I��Ѱ�<p�B3L�2�;�3�$	1ben:D�� <���֠8C�b���O�d�=l���Y��I����@��=t�r���ʕːE�Ɠ`���C���8mT]�7d�%l^���'�$#=+�T�ʆeB��ޑ3c�+�"ݠ(s��:�4g�)1���?����?������$�O&�ӉC������v��te,Pr�@���=��T�L~���,�� ���(bF���C�ɍNt4Q�鎗�ƭw��#�4�e��O p���#x�����Rwh����?T,�C��}ߢP3vk�6�"���Q/.ئc��P�}���, &�7��O��Y 7�c3g+�Ȃ�� �$�On�`� �O<�~>�a�O�O�����)
��r\�ep�ˑ�'4z�����D�2�P6A_�y�	Ɓ��p<�C�ş�N<i��\�n�)���T�Z��uQ$K�<Y�j��q�Lz��(F�l1��\K<�G�i=���FlX�E%��bP�1I
�'g*�a��_;�%Ȁ�	/�"
�'4 ˶fYo#��Y!h�--jV�h�'��pA�6v��bE� ���j�'����㚟����>i����'�	Ѵ�T�Uuv��Z�LA�'�>����)�d�Ɂ�Ň�&�
�'�XY��\9dT����f��1
�'�����=$��"�OC�܌�	�'~�L
�l�0 *d� ���r��'E��
��ԲC�+���H��'Vm�M�l�^���A�'?P)b�'{��xs&	�yp�(�AX&4��1	�'SP8�Q���wҐգF�W{�8�ʓU����a�?
��Q��0�
%�ȓ{�Jy���%z,�1
7I@��j��ȓmM�Taf��%���@K�* ���F�q	E�}��8�)�#"^
���{����

oO���"V�C <�ȓb�(�ED�z�Z��%Ϝ}��Ȅȓ+�b�i�e1f*�@�� �M9`̄ȓ
�-�V��Pt(% r��u'���ȓ�81����!e���f�T(d���&t
`�3A�N��I�	r۔��ȓ¢�6c�A�|p3���
L���ȓ'�� F���w/80{B� '�p����&�2�@�K�j��&ǔ(}&e��,���Q��gbb���C�$z����(��xDm�>$�Ő"r�bم�*�����eP=��%"0�H����<4��dI�Wh�9�A�P�����d��r�E2	!&u�@#C0
T��S�? $�C�%�-A�fE�H��Y�A�T�2�0bF$x��d"t"O�%���`}�����3���gn��}G��r�!��JʓA���É�HT"(���Ex��y8ƩN��P�KE7; q�>Q��~���'�x!A &~Հ����� J`D�łW0R�`a�SȊ�HO��	���w�N�F��F�J9H�b�.��0��0.DL⟢�D5AB���$e�p�L#�A�GS��AH[01T�2��M�%�̉P�֬/V�{b�^�L(Dxc1黟|���s�S�U�GT�����e^�7�ɋ������r -C���i%.��(�^��t\GR2�sU��~���'�����C�4��Rh
?/�U8N�h��4>�^a�t$�>��A{f@.��?c�,xt#�57а����)r�1��IN������_M ̓�I1j�ݘFkY�"`j)���	�1���nM���J����wF�$FѼ=���`���E{��I[�xJ�[2B��$�$	S%�%mTZ�s�I	4�F�җ̏a�峠�Z��牧8����NŕKh�����#2�����!���
�.��*.ȹ��s���̹P,�a�EH͊&m��:�i]��	�J�ԭj�N=�����b�葮D�	J��s�U%-��I�H�6�����
�@���A�V��"<y�٫���K�7�N�[��oң<A��ԟ��e�4t�~(��
e(�u�u�Z�PMAc�G�2���<��*%��t�q1ﺁ��ϸLQ6� ��[�6�\���i�"�Gy��	d�����EF\�gF�t⡂eH-���8(`Pw��
�s%LԿY��OPj��B���k�)��<TM�Q�O���.��?���@>j��*�*@+f<	�$�5��1
�a<Y�J�g΃LQ!5��p�f��A�4,O�e�U�\�4|�LI�*:K~QcƟ>��fE:4�����L<�ɔ��p��s�lMx���;.��W�ő |59�Obx�̊J����k�&qД�R,�L�̭�p��j:F�<��1P��V4�F��o۪N��z��2۾Jql4ғg�pԚߴ��O�z���L"w.\,@�D��#. �2k�I�Dȸ��rJ�r	���6O�\O#E�"UCT��\�:�R�j�	Pr-S7@��h�Q��N��� (��OT��e
�!W�|Ɂ��1o��I��F�D�x���L�\.!��	��~�+����u�*%�I<A��x���СR��a!��\yBG�J�	�yH~���	�<zz�O�	���\<E�\�4EW*t�"��eV��O*u�&�4�m*Z�fE��7)f( ��Z�	��x#�n��v0��4E�<X�5�
;/Ң<��:Gm:-b-�O����圼+��m#1��3i�8�/-�p�<�.*��\��g+�	n�(���Ļ
�`�W���^� �}B���  ��Vh?���\}yB�i�v�x@lU�U䲥	T��64i3�'+�� �-]�2&�P��s�@iG��C&v�z���X�4����C��b���	zx��FC�?��D �O�柸u�-�Iψ��q$f�����j�67�'�BUQ�'��ۈB �p n*��*j��q��i����0�԰sZZ��B
'X؛��'��rN[K�����52p�qq�j�"C�|�Hm_��L�{׳iR�R` ��\���EzZw��0��M/=�k,7"��Bo�,��y	��S���p!V�N�	�Fˠ�>ͧ�qO���@$Z���� �k�A��81�O�D�6F\'Bh�(r�'B�,;E�K#Du#�iPP�e������m~%+ற����*\�SSʜq�r��**7���	@;|�
�DdV"&@�,p@E�h ��C���f$`��2't��X����$��y��<Q&�\
�܈EMZ)��	(9�����X��37g�gJ�㟼���?4��p�P鑳� e��}Κ�BQ��/��		�>*�Fw�h�7mΨp����Jt�L�C�0S�CBK���<�S>4UL�A<�X%��F%.W|S�&@�i�1��U"Lq�U�p�!e*�ԛ4T�`�W�Iº�	J�6dpS,"�r\���Ga�\����U@\�(Lؔ�U��E���C8zEDq���ŷW+�))3p�
-
�[�$����(O�����	�/�B��N2�X��Sz�\̓� ��`k��#Ak<����X���(Fހ&�jS6�J#=�̀��'t`i���~Z�Ɲ>g�Y�&�T00�hyp��`�D� �����b� +�Ѻ��+^�O�}k6��cD�s�� ;4�s"ĠB{n�Y2B/Z��yb��}�	�Ot�w"H�I+&���m
�u���`iP'?�����jH����e�5S��9N�z�KX�(��]	j� F��s���S�,L*��}h�R��Ey"Kڹzl��`��C*u��u�ҋ��]�>��*U!W갻���"N)T��M��.��Qp�����҆�W�0�B1q��.jH�<0g[�DEy�*\���,���
2~���XFB�Q��0���2�d��F�H����h�.�!+W$Q�+�4щ҅C�1��3��>a������{%zY"�(R�M@6Ԁ�H7	 �^�m�ˁ.� }�s�T$D�?���]
ExE��bTq�3Č�A:>`�G�X�w\�a���OD��	��6��;|Y�f��6�#�τ<$�(�#�ˇ-�lp�e+1��?�!�ǔ<dX��&4,�}��b�D�
C���?�l@��'1{H` �Lܺ��d
6�>ʓ5!�E�`̺a�IgNe#T�T�'�м�>!Q�t/|�5㖱g�h�;��H��zD՛%��+���Q%��q1A ��~b �
Q��	`y�O�\	���@�~�H�H��!�V�0�� 6k`��b�|��aU��b�w@-��l�1����eR���`� �piU� 8�G�% �8zVBPmyB�?9˔ ���I�9��"�%=��O&Q���ԭYyb<��nW��&1Qt�i����1#_lx�4C��3CL�������Y)Ȧ>ao����<�Ӭ(�7�V�LPݘ(n�M�+g��{C`W�*���N��8��O��<)O�� \:4{~��A�R*Mx8�d���'� ��ǈߣpi���F�
٨5�-O�6-��!lSB.E�$�^��򊋤}����22�B���ԟ�y���n�x��`�	�X5�V�߯ �~M��&��*ɚD�E�+���4�ǔ��g����<%?�ʀ�K� ��aؑeI�S�����DG���dW�eMN��6�3]!2a��"P�-��OXQ����LJ^(K4$<?�!C�Uy�T�#G�~��)�JD��#��<"\-r0MI�C�2QX�LԪx����'�%��?-p4EY�&�N�8��5p�&��pR]��3%��*Y��h���]�y�l�d�9���sS$ߜ7Lc��3�&�\:����:��鹧�=���*P,9�aj$ ��!�G��
A�I�'Np��� #��S&�R0O+dA�a�rgV�1�䖰���ѣ^�� +sn�<� q�Ef�[�Q���'�J��Tb�?|��X��E��@)L� ���;b
���V�A	RJ��$��%&`ʷC�?S���5�O�o��\`���?�S2�+H=�)X���;�Ū�^��,��^P�[��r��.�����-o�5���Cn!n�0q:%�^�(�D�O>�=E�$Gç$�08�K��0�����e�*�� �>��BVg@�I�0���eRG�w�ɹ9������L�U��D����@ʓ�(O��;eqQ��x��'Pg����=z�1Ê�7_�E�k�+}�a٧��P���x�-O�y1�#<��<YQ �
�|
W��!Q7��m�C��̅"n�$�G�
�YE���a�O��0p�6S�����/+"0ۓ.l�&����	�&F��<�4�S}1���Ʀ��Tpi`�cߣ:��k-��?��®��X��Ĩx6���f�Z4�lm��'���@��c�]�S�O�:r��, � �!7O��t�� ����B��t
�
��@XGf���	1�L���SOV��jq/�_K��I,}jy�?�'k�t�� ՏeQ�h���b�8R��$�l1�$�>� a�\+�d��4����Ë�N���g}D�Oo�4�N L�ػ�.͐���Y0D�g�F�t�F�B�ûa0"<� �K�:��@�<>�����K��Hp�	�8 ��.	��;���?7-[9}'D|�����z��;f"X�.�p7픨oU��SU�ǡ�(O�t�T�F�z�(�9�ٹ6���'e[�H�b0�ס� Q��O:�	ғ3�l�D:��-aL
�1䢅�&!���̇8e�O� �%F�"O4�0+�'�Bu�/Oh7mE"qYD���L��%��a��ؗ{��%%��,ۀ�O��SΓ��|Y�oU1����A��*Fy"��t��k�t�b�O�X�N�`�/��X���;�dL�C�$O���^C�U�'I"_�έ�Q�>�R!^r?�Ua��J�hp�1l/�	�b��8��m΅"��A�$[�?�$a*J>A�,K���O�I���O�K��xT� ,k��0���܀�M+s�S
�a�#��?c&C�A�0�D��	���)"C�l�<l�`bٙkD�G2�\�L��'n&����|o&���N՛7���Jv��w�21�\��%(n�����w�0O�rJN�cJ���Ӻ�I��>����(G����X��K�⑐h'�-I��$!A���-�<}2=�W	˲T��@�O |^���/�c쓄�@���"�F�+TH��V�E>����O�1����<�l,S �7$�Iq��dʹg*ɨ�ݏnܱz�����M�ēkh4s���O�](M�ʽ��VW0)�,˥�(O�牼Wʼ�;k0��b��BcV6,ps'��CT5��X{F�kwf4�9	rc_���0�8�I���	���"^�,p��>p>$�'���$�<����ʚ��6�x�'��᳐�ԟ��[aEN��t=�1�D�g�,0')D?	���3�o�[5�L�u��"3B��DB�y��Q���I	T �¶�DIh�����d.�'�v�݇{H�]*�bX֜ʏ�LƯ�Xq6�J�F\Hڄ�� Id�<��ԟ`�����=."� Q`�%z�(�Ɗ?hm��*(R��#=��y�J�U,�բe��{w��rA��"�;���O^����
���'/�Ԡa�Uo.��3@ě>���&�~d�#>���U3;��y�ƯL8P^�řE�\�<IM�J$<�`�C6zn�!v��}y��|r'I-�(�򀃝.]X��%�ȍ�~򅗵J��[�W�pA��,v:2y���J��-����q�Y�]��{��������,(�5q Ԣ�����ʲ��D���<Piߵ%a�}�-��f�����a�!h�y�wG)>����"eY
^�=r�O��%)h�}����`is�W�y�
�3��2SN���v�|D���Q���7��ΐ�%{�Z�����>�ڹ[�hĉ,��7ML�Pp"9@���O��M~��a�[;c��{�/�C$rb��I�� �\�48���/m|���!�D�>������	@T��/�?_��dLu�N���(`�B�ȓ���&���Dt�a��Ӵ1�4%@e��;3�l�@@�	6P�>L�DC"޽1�J~��#-1����O![����T�ď*n¶��!��i0v%�!n �=7�O� �ݓ BѺ2��h)2E6j��hQ��]�m��םd�O�ځz�Dݣp�Ja2�C�?�䔪E��W��<S�6aS�����R�+Q3�8%*d'��|L]�Tb
m�(8p�S��"��9OV���'�)�|�J?�Y�H�i�$��E��H��2D�d:�$Ng7�I� �,��x�B�$D��"���x�:���3�(c� D� 1���c�DQ	�b�Jnԙ�3D� ���҅{�t����2R"8@*P�;D�0�1nP�X��QJ�C=��`��&D�����QHZq�0��	3Ϛ8�':D�H"�!�$K�>eev���U&+�!򤞒W�@����T$y)d(ܵ<�!�F:!a�i��D�9�`�s��p�!�RCP��A�ԖU��AKSǕ��!�D4V�`�Kbcڥ�ڰ� m�A�!�d��l������4J\R��B�'�>E�#�ɯDxDi��p�
���'�6-ҒB�F�БY0��X����'D0PQ��M�B�����cx�]#�'��@��/ wD�X��+qT�Q
�'V�Q�B��Q��� �,X2�	�'�N��F��r��4!����'�kG�
?i�`�3F� �02�'�u�'�Kj������b��)�'���5��++�e�b"��U���!�'��� ��Ko?nt�ҌƶY5�$��'Ђ����C��YQ&\�T_0���'�C �^�F��*&��^���'�T��q�8���;��;+O�c�'�@|y��n�Ρ(3MʮV�~�k�';�`@���_��y�B'<n4��'X9��ʃ�5���q"_�a��z�'��a�(�=+�䙐��$���'x<��a�e���Ӱ��?7f5��'K��S�bEq��S�*�E��'� ��@�dܭjЁʫ�*[�'�(D;��_��7�K�J}q�'�� �O�D5�	&ԋ2�]z	�'Zp�o��;�p��̿s֔�9
�'j�E���׿R�&��1aU�w`�B	�'��p��Lϸ[�
��7pi,j�'�,�@�Г_��Q@	R�;��s�'պ�)�Ɵ�'��i�1�4���'�4a*f�ؖcN��@��
�0���']V��cM����m��L�
$U��'��nQ'y�H�.J����'W>)�C���2��SF���Ф,i�'���	 H> �:�"Q��.���'e|��m
��A�W".<��'bX,� �ՃkT�,���O����'��@�!bG,Z��ʡF�*A޵B�'����B�1��|��Ǘ=#@<��'�@�k�M�-]�U�v��$ ;�'���k��_5��Х��l�
�'u��KL8n�.x9s.2DS	�'���pbC�3x�p)���+���'�J豗���p�`�*IRϪ�c�'w�i��Ă`h��J!E(�4`
�'��=���\�L ��G��KRԜ��'��["�	�z 8ԉ�!�/�����'K�XC�#�2!N�24JW5&����'�j�	�\.{�%��@�o��|��'i�p�$_(@�Y[w�>z��a��'�D�Pf�u?�w�_	�<�;��� �P`p�K�g -���x���"O
1����$O\�ȨVf p���"O8�cV�aB,�0�h�X�"O,�)pÂ�P�8pr�Տ9�|1�a"O�T@B��с�OAϨ���"Ony�v�O���T+�#�)�"O�9V��(-2��J��J7 ��t��"O�)З�Ga��9���ď��Q�"O��6G�e>�[�/��@�����"Of�����r�ӷ�τZOf�p�"O��# &L�,��l�īA
D4j"O�E�i�'6���_)gR�Xy�"O89��)BW0\҈I$a�(�"O&-`��['�Zi���K���"Ov!׫Lu��� 3댺=3x�C"ON�#�
�e
5˄
CL�TQ��"O�t���\�G���EHK�+�P�2�"ON�Q7�ڬj�ʅ��-�JӨHhA"O�������
�V����Њ���"O,D�do�$U�j=����{Ǡܢ3"O m�#��LF���#1#��PS�t��	d�v��o�`���JBk��a�ZB䉁o؈�%�(?��e��'(aB�I(�m�QH�Zp�p$J����C�SEzd�W�5	�LQ�`[�
-�C�	�m�B��.z��t�%KF�=�C�ɊU(z� @�2��k�*+v�C�I�3$�j�b�$dX�HGE�2x�L����;��|�'����b�<odX0��+Y��ȓIΘ����ޛKF\�UF�O8-���"���	�=��e*��HO����ȓ:�؊�`ػ&F�ʷcߎ&qL-�ȓ�(\�c�M�~����mͥrl���U����r�ؘn��e�f� 8Bٰ�ȓQ�����ſ0.������ȓr���Q��@��a�T���1'P��ȓB�-A��ZgN諐�Ȇ3�^<��M��hށ/�\��nD)��=�ȓjCV��1���D�l)�'���D��U�ȓsT���aN��i�����>i��M�ȓT=�8	�lS�&Q)�W�_o��Y�ȓ�  A���m�@pq%�Y�;��$��C�V�
�	J�X�� ����	��T��x��PB��8`�l���&��Ԇȓ>~��
F1�)KԃN�e���ȓ]z�{�B�!K&���+������d�	v/8�4����cf|݄�xI@0�D�B3��Q��/�T���O��Jx�eٳg\�Rp�`��'9�Op	8�,��9��9*p�L�TV�)"�'�!�d��3�<%qFN� V�M�az���]	\��,�4�@�|H��Y���9!�D��:7���d�RP��H�PQ��G{*��4(v'ڣ"�ޭ ����(�rG"O6I�w PO\���K
hs����"Ob���B6sm�["��{r��P�"Oj|��jұgk�lH�KU6zI�,�b"O�aCf�P'Dr�d�F�� �"O�%������4�7j 1�u�"O4 
qM�>�x�"j�:'� �jP"O,��bJ��غ��SU���"O�XI�K���`c�*�A�6��R"Op�K�m��B�"�`��M-k�b�`�"O��V���&P,(��.UҤ���"O� Z�1F�L�@UJ�]!#*h8)�"OJ=%��k�
%(`Νfe��"O:e ���,|� � �o�l��F"O�ݰ�̄\x*T���y��}1�"O��)���V���"?�H��"O� 䈃n�y��(sS�uYP"O�"2��!��KXwHL=��"O��ZS��l��G(C,=2zQ�"O����G�p8���Ѧ��)��KG"O�Š�!B�[߼�ۢgL�F�6$� "O��a�:x@��j�f͙R���!�"ғǈ�� c2�i�J��@ -����D6�S�O ����˂J]�mA���5�x�'7�u��n��B�J��u��u�ع�'�y�6��)HPE��l�5j�����^X�\R6/	�F�^�����Tp"�1D�l������)�$M�8P�w.�O��=E��K"x�V�a�-_�����r� �ў�F}½ih�ЁaEƌJs�� T��9u��)Ȏ{��'�r�Cg�N�B�RHRC!^�z�����'V4���؊j$a���&v���S�'n��g푣(�u��[� �k�'��$З�JW�r��U鄚}9ƥ��'?�&� �AQ$i����i	wK����=�S�O&�L�	�b�᫡.�g���	��hO�=#�i�2]b���=�.l��"O6 '��R��Dq��F��]C�"O�$H��*j��2g�ՒB+�x�%"O��#��)z�i��K�(T�����F{�O��'2���s/F��6�H4)����ʓ	�\�gˎ".��y!��,}2���iʞ�0B�;�ʄ��ҼQ����R�̵��mK��ĥ�$	 h��O��D����%��q��F����G�}�/\=�%!U�*!.X���MX����ňxQ���!�+y&8�'Xa~rO�W�'�	�"_
t
󢁨�yB��
pM��Oš LA�2���yRk�?]&h���#
�z�������y��J���q�N�7( �}괪̙�?9�'�n9�n�j�@Mx���}�(�	�'"�����~�U:�cpl ��'W���+�-U�<P�aW���X��D"�S���B�D�xM��j��(� �C��>�M�QVN�/T��,rΊ/-� ��u$9ғ�p<������%�1n�s��Rr�<�d��֐!�/�"��-u��v�<٣���R#�չ#@'^
h�hţ�J�<ylL�4|BI25L	�E5�Y8��G��H�'-��;DH*2�b|j3�
����H�E{���(U:B�ݰ���3���RÁ]��yBcF!D�d|[�1�4�*�O�����6�S�O�tQ��J$$> XagHZ�=�0���)���=j�z����ԏv9�)I��	a�&��p>y�bܮTA�1�7���F+{����>������<KF(����;8W���6`V2pt��$ƂZQ8���	'|o|�K�*u0�,���'8�h��Dr0M�	L�Pt���	�'2�T��&�q�t����F��Lb�'�r��!1"1�"�!?C���b�)
3,�"	4:�&(΍*��z����y�MO�kf̉�d�.P4ٸ���*�HO����b+v�Ñ�39�ls�H�f"!�DD� s>�#��3?Dl�W	B/tqO�=%?� P��@�2U\U:��)�Pqg"O��@��';4�$�ܣ.y�x��"O|�X��X�6T"���3_��"O�Ī��]Z�r(1��Ȱ_Z̓"O�Y3��Y<7�8�@�	"UQp���"OJ��$L�u;nq�IaA��yRM��]��x&I�)<ܕ�G#M�y�.T�.�6�*C�-6�h���g��y�(=1��"@޴zjti�c����yb�	yVza�BΑ�z>r� �I<�y"�׶0�Π3*�\��,z����y�/�"t@]c�D�"R��Lf���yB��g�V1�6GM&Jn�U�%�� �y�A���y � �B�\8��\ �y�	�?�̴kӃY�@��(�.S;�yюX&L�a�S��Р�3)C��yb&�}&u)wW���{D/�/�y��er0}�!��n�5T��y�,{�x@Q'J�6���Z��ħ�y2Ι2[�$��"+Z����W�y��ë=���h���'��iK���yN_�k�B�J�aQ�����B��y�ʔWkQB�3��i���<�y�gM+s��X��Q���IR�U"�y$�1i�L��c��NXP	���+�y�ʐ+py2���hI'vU���3���y�+�m$�� *߻g��ÇO)�y��թm�x�*"�,[���s
��y"*�e4�-"dI@[=⬘���4�yb+O�5Dj4����bD�R-�9�y�gG:;{|���T�t�������y�ώ)n�����Q؞ɀ��&�yb.�|%����ҞK��UJ�����y�	sx^ysUf <��x/��y�(D
&�=��Oۏ0;����
���y�"a�P�T�4q#���&�?�y�n_�/xt)Y�L�p(���N��y2Ȅ�����g�1j���M�y��T�N�(H��V�g�v(#���y2`�H�����Kæ]���'��,�y"(
"Ԩ��
m���b**�yrhĺd:���Z��@�'���y��G�l�.ت��̳N�Խ۶��yr�t�H�*����A��'��yF��~czL" ␰	e��c&�ұ�y�nI�1����J
�z��1ǋ��y�72B���I='P�k�����y�I/+R������||�l�`G
�y�gB��LE8J�yV�]R�D��y���+�Z���{n�����H	�y2&_|��B��_uĊQb�dY�y" ��zE4�;f�rf� p`�7�y�1[
��f#(W�4�b�8�y��J2\�1pׯ�<�p���Q�yb�ޘwPM�e�\	�(�#���y�Eخ!԰�Q�79��R�HR�y���,�Z!�a�@����4냛�y��++�b�r��¾����yb(DV~f�����s]�,��ݝ�yr��B��Pn
<s'��HL��y2��x,�a�C����mH+�y�$<\;�8��h��^�D�hA�+�y2�F��xv��W�XԨ�Z��y"�ұ^�LM�g�3V� ��b��y
� �qa�M���0��^�a�t�"O��Q��߫&���`�"�7ad�e��"O���G e��liG� F���T"Od�1pI�m-�0�UJz��AC"OhiPb�ˏS�<Q�&=�bJ�"OD�`�-R)h��LjŘ�x�PE�r"OiF�	YM�t�dA�l�ޤ{�"Ou��A(|��0�N�$Cd�"O�C���
)�mY��V�[b�T37"O�h��6���cu�� K���"O����ۼw�sF�L7x�#"O �� �����Ť�14F<�Xb"Or���]�~,�����H0��"O��"�BL�}95��qEL�;2"OV��%�V�m��2qVMB"OvP �Q��a���$�q"Oȑ�ӧ̗cƅ��Ⱥ ���Y�"O��3q$��{��8���J�U���	"O�m�C(6�L@�fE"�"O�}4h�i���h�X1;����Q"O I���&�fU���N�g�*��"O�I
Gc��8�P,ㄥ�fi���g"Ojy�� �:3��R�N6]�,(��"O��dKPZK��ӌ�?��Q1"Ob��O2p�RUY�LF�;"OFLXЀC&K~>u
�	�3?�
!	"OF����FZ�L9�cF��d�1J�"O�����'d�d��ǆ_fh�%"O�QB���V����[�����"O*!��@:�fZ@AQ)d��PB�"O�k�D��5Sb�EW�4����"O�07�AQ��� j��s`��r"O)Ѯ�5i=�5�r�Ǆ*]>X� "O��!��6Uy �^��T�7"OrqY樑:`��=b��P������"O���k�G6��B҃��d��U"O�=��5�>`�LV�Ń"O
�{��ɱk���ڃ��
��*�"O��˔o�x		"���~��4"O��P�m$�J��8u���"O�A��d��S'Tm�A�V�IO*	��"O����C�Bx���?$f�@�"Or���cˁG�T S�3�>
U"Ob`d@C�|�����/V�7VE�&"O��3E�*�����;"����B"O�1�׶-���TdΕ	 ��ң"O:�pѫ�#���Z��M%P`��!"OB8�#�Z2��@CeV�N�L=ѐ"O4`��������E�Z����"O
@�6,��t�S��� ;��}�"O<�R@ζ�����ϊix^��"O�ԡ���	 �)wnJ���5��"O�i��`�-aB�:NIb� �"O�r�O�b�	Ƃ[������"O܄P��ZR:�&�I�w��T(�"O.�3%c�rN�-rFAG�6�2ЊC"O��C����2*�jŪ	�����"O��S����|�k��:j*4�%"O�-��)�6'59��ѿj���"O�����&l�ksH^@���"O�h��vhP�����/\�,���"O���1m�<��IP��9Z�f(x�"O�C�K�-��� �N!�<<�4"O8(8����`������8�c"O� @Hڕ�5By�l��	�k��"O:���$U*}�Jc�)��Yg�� "O8�k#��6x
5 dHQ8A=���U"O�]��EDvV��C1kR�p�W"O����C$~�] �e�O�d�q5"O<�I����8���9RD�(x"px6"O$�XcbкLa0����M�e��z""O>\�I�~��c5C�X��)�"O��wLR[�~�أ�T�A��0"Of�2)Ɵ���d��Bq�0�3"O��RD�cu�|��P6iY��"O�i;�~�@0e�uSL�2"O�@@`��5]�� ��k�
��"Oʘ[BEN��5:�t�D�rC"O\�� b�,�8-�6'08dT$c�"OT1Tϊ.p��z�/d���B"O$�!q�A�-�@��b��wIHr"O�����.M��'hLx�
6"O��Zc�s�59TFؼt8 ��"O|D���<� �I��-!^:�"O\Q�O�1o���A�2"�!B"O�ٖ�'=�>rÔ�o�R V"O�,�rn��[�Buy��\�vj�"O�PV��7w�*L�㪟�(����"OV��&W�X�:y)vD0y�ވ
"O줁D�j鑖"�#q�r��"Oj�r��Y�EX��($��2p��%"O2�Y�.ѿ`JZ���ݱS��h%"O��,@5tM*��H��e��"O^��3�Ξ|�K���t��"O��"�S!�ZT���@��8��"O�h��[�"/��*�
�9��Â"O��X��"��d�p	�5�|�qR"O|m��#�>\��pPH@ �6��"OD�:�.��p3z����M�04"O�1����MX�(p���-�죓"Ozx��R�-T�*�ƅ!w-r}P5"O��p1 ����i%;$:B}*"O����$����d 7S18P�"O�͠��e��̒a ��X1Z���"O��h�m�442$���O�hC��["Ol���<,�2��% aQ�u"OBbA�
7Q� ���K�kYV�� "O�A���23���K��-IK����"OX��[QN�L����0.,U��"O�4�DX�zmD ���>�a"O��S_��`	c�.W'v�8t��"Oج*v�a�%�d��}�J���"O�١g�U�"{1��l���c�"O$�*ӆǡ_�D:5kˁ%���t"O 0#���*JOH�*�
��
7"Of����'P�> y�+H&D�"O � ���t*��RF��(.�!z1"O����%ִwʦ���˻DƚH�"O`aX¨�?���9���^��T*�"O	Q�EG'u��$�����"Ob�sg�Z'D�[C���]�Z���"O���#l�Zq!!I**��p"O���!�7A��:a�?����7"O@�6흏'���um�~��[�"OB�F/��M�.���n�$���"OX1y��T�؂ ��D& ���T"O\��REW�9$  ʣ�-sZ�8�"OZ-�0)״XC�u�ӣ3dt���"O� &�)����6#���-N�TpE"Oi���9V��A�C�1=J��+G"O�!p�j�*P��������Ҵ8�"O~�B��~8:U���݃D�֭��"O���� �3T��:��8�Å�"OT8R���8� 85"'�d��2"O�I "�Q,�l���B7	�h��w"Ov�
������KsR�s"OP8�bI�>�0VC�Fi:�h6"O"�A�X�o34�S)hTB�"Ox���(M� �dNL�u��4[�"O����(ߺf�<�(Ս¼5!�Ph�"O��ڰ�B�BZju��+��h�ܣ�"ORY��Ϲkvn���ٞv�D��5"OF��Be_�T���F�X � %"O��;B�'1E�E� @��J�cv"O�D�d@��<�T��Ѯ��D�P�"O\y��&��l:�^
=ɂ�!#"O� ��MЃrF&PSP�F.���"O*�T��:G��jj+]����5"O��j#$T�6��!�V�+�"O
y�V�ظ(f�ysfBM���pU"Or��D�@.k�)�cc�
Q�2"O]Z��נK���D"P��n	Ɇ"O���ƪ%a.d)g��2���@�"O:5+j;��x&�y;���B"OB�$T[ԾP�G��:y�hA9Q"O~l+�E_0/Q��bC.�1{,�d"O�,�Fۣ���(���^o��9'"O�M�bh��,��9�pŃ�2z8�U*Or� @��j  ,�񪍵ۚ�S�'��1!��v��E#� Y��p��"O踁��.�r�C�i���R��'D��aG�]� �4�0���ZmX嫷�2D���ԧP�bV����0hd���F1D� ��O8�$c"��4�B���-D�p�VBWQ�l9�̈  ��e�+D���'�Q�@��{�郯=���+D����새7fN�R5H0��L:3e*D�0��#$��X�� �`N4�Zd�(D�xH"�5]�j,�#�	P�6�A��;D� Y���x:��I��xB!%D�$Y$�
��R��U�(��E#&D��!�g_26��3J.Wڜ�"	&D�("5,o)#FiK6��c�eB_ơ�d��9h����.�
M��P��y2�G(`n��L)z�p��7�T"�y���+<z�`���p��i2GJ�<�y��ۖ:SNdB�元��;�W��y�M�/R��1����7�`%iL�y2���Wo�q��	��J��Pb&�y��Jk�V`�uaWx�l��n��y��z	"�(�,,$o��pE�
�y�B��8H���ͮy:�R��3�y�*C")I0��M�1.�B4�$ ���yrB��Z�x����&w�:������y�燀:gx$�ek��|(N����yrHξG�ɚ�MN�qaV="�ɴ�yb�[����ޕ^�V��b�yb��^f�(*5Ä#S��"�,��y�jѬ^�dx�1�%+:��A薫�y�P�uU�ݠ��5.<�VK��yҊ�5�l��׬쨵ؖ�?�y"gQ	��Y���΃z'�hv���y
� ���ӊ�2j��$Kdg-y��h��"O��@4��l��3'`�KWlL��"O��8��,T~5���9-�"O��'u�N����9H2���"O�$�7ł������C�[L"Q��"O�B�G��o��Xz'A�.V�<q�"OpL�M�G�E��a��>^|T	�"O��*DE/'����f�.TP��0"Oz%[P�ӮR�
%��g��̅�"O| ���B��Z�k$�-+���"O~X���թff�3��5��"O䑓 �1(. ��s+G�<��-1�"O:��(�U�u��U+Xz�y�"O�l�TF�qTͱ��T0j�<�'"O�`��,�Iש�jsVxR�"O�PSv+��\��a�T��"\đ�"O*����?)�@	ؠY��9�"O�5�ե��oJ^I9�	֥ul��(�"O���@�`�*�ƿjH��"O$�1 ��g�p���I�<����"O�!����@FHH;�E����"O� 2Ѧ�=:�&8�d��.�PH�"O*XC��F�>�"�p#)I��k"ON���k��q��Bra/3V�yhd"O�:V��*qu<��t	O���A&"Oġ�!k��hmjwG�x�v虐"O�Āe�6o���M_����"�"O`钢�EgJj8H �V��ؙq "O��YV$��>:�qxpLW,5R`��"OpUX�g��X���XP��ũ`"O��X�G�h2�Y�s�ۘ=ݔYI"O@����*U��Mz��$P3"	�Q"OT8!K�g~ٱ��	G�Ј�"O>T��C��0l�h���F�Rl�9e"O�XS�߃= �yu+�1}�A"O4y3�O9ǀ`��Ț(%2�V"O:���C =CA�(@5I)	��Ɂ"O.U�#EuP�j5"�&s�L��R"O���`o�-��b{�̉#�"O����@̀x��i�w��g=��1 "O�Lq��0��ƀ�
sG����"O�CQ�0隈���D1�F"O���䂕�c1�R�
�Q��"O��y�l@aŖ�B��"Heޅ�C"O���T+1�f�RΔd(J�y�"O��y5�*X"�B4:�"Oz�ۣ#D_HT�a�H�! �q"O�`"� ޘgVI`�@��i�0�"O�����_:�ֹ���\���Ͱ�"OKR� ��,��[�Q2B��"O�a� h	�6�L}��D�"6�"O���7�+�����S�����"OX��#ʱ^��eJ�L7p��"Ol�ӵ�/C:��*b�ȣjY�Q"O������y�,���J���"O�)k���=W��X�&�ډ)=���S"O�A�c͝8����cL�N��#"O�A�D���PB��A�LϸCL`�"OU�%DS; �D��?fƾ$Hs"O>ԡh��3���R���X�p��"O����/"!� ���GL���"OY���4]��aw�W=ȑ�"O��uI�,L�b(+���&�0B�"O���X	A��p��N�5n�S�"O� ,y"�I@�v߲H�c�Ծ]�6�Y'"O�%+��[�a��x�'�ܡ�~��"O���c&��C;4��wꕆ�b���"O`���'l�VȺ��ޠ��|;A"Op"�L��G��ܺ`gG��|�"O���.�8^6I���Q1F�X�BA"O"�إ��=0�8�ӦC[4JA"�"O��Z�͑�t�a�A7Z0�k�"O����oU*="`�c�Ś##b8�"O�()d�P�t��\��@�	[����"O�!A�슀�@	��	GB�X��g"Ov�A��B�q�2x�"�V���a�"Op���˓�)P�4�Bhy>��"O���wH��h�p9�#�B�fẍ�3"Ol�#�˙�&X[ƤQ'e�,�w"O|�3D��&��pn��]��$3�"Ol�:F��%7u��1WM��Ui\���"O���d�eg:y�u�d���T"Oj�ʥ	6_�f|J��ߑa�HC�"O$1��h�y>jL�E�VL�E�@"O:Ekq/��Kᖨ��C�}X��G�<��D��a`�� �:�Vi�2(_T�<ac� �&԰��ө�%C$Xh@o�D�<!�a��W�(��&֗���K�l�U�<)�i�$�+�(�H_�H�E�FS�<c";DN ��EX'�� u�'T�ؙf�0F�Q b� 8#�i$D�X��d 
9��A�D=g"��á D���P3�
	#r��{����-?D��`�C<�X�;�gL�� � 8D�l��\�Tv�4�����'dx�p"D�$vj,ΔTy'�D�W[H�:�$D��Ӯ�3�`������n�� D��acKNq{���[�`�H��WG<D������n��F��+>I��>D���U���R�(����3�����>D�8��5u�ѡ���8�d���9D�|`��ɜE����b�b��F2D���28a��9y�:B���hV�.D�@B6	�	vl }Af��6x���*D�<�� L!h$3�JT	?�\��wi*D�d���Q�24���L_2���t�;D��g�N*�V�-���$�8D���6��a��)�!�$7D�ؠ1��H�z�9�(C�.�D5�4D�����V�R+!/�F>}c J/D�0���W'T��a�ą9�%;D�xW{���{��95�M�9D�4 ��Ėw|�L���F {h|Cь#D�<���۞g���*��,R�*8�6�4D������!\b�	CJ�(���=D�@[c� �<���T :j@պp;D���dH��D�C�^PB���:D��C���vc�ma����=D�H�1��y�t��Â��Q�d9�V�6D�L`a�TY[&E�54ah�3D���+˨{�,��� (��@�k,D�����R(���*�?L���q�+D�@1f�-� j��U3#�x��'D����'9�e�V�����ү2D�X���Y�|��f'�Ak��1�/D��Bda(\|�H5�4v7����"D�hY'�->�"%!̖6�.p��>D�@8���rNb�Ƣ-@2��ag;D�� �$2��ມ[�Q�����S"O I�P� !f�(�*`/X�j�ʜq�"O�\Z�=qpXS�'�H����t"OD�Ƥ�`Z�����T>��xP"O$�ĒT�j�k��)�\"O>�Ӕ��>����_�M�X#�"O @ ����X���$����"O��#�ː�?c�yaփ�F�XP�!"O�tÄ�#g�6@��\�:`(&"O�<"�/1	b���1�F:x���"O�a2�+Z��$���b	�a��i��"Oj<�S�^�F`��Ƃ�t�"O�=s�)G-ݜ�g�ܕUK>���"Oj��s$��l��eDYX�"O��Y�������ǿP�i�"Oz���E�m�D��e,��lo�峐"O�)K�?Y6|�TK'{��'"O��Qn@A���ǩ۽Mt�y#�"O<�X�F��<�ZlC2銉sZ����"Or�VO�.@��0f)A�UF�j�"OQI�G _��आ^�#;��B"OH�SQ�G�����ԍw��9�"O��7��� ɑ�C��SfE�T"O�jW`B�l�4�0�#�0t�գ�"O�}�l��r��, �O��u!ƕ8S"O�b���I��UAuV<��"O�9c�+�(%5~pB��y�s"OJ�r�aH*S`�lH#C��W�5�S"O`j��׷�,�1�@��~�s�"O4h���#4&�<�wBL�d�T��r"O�Y��^�kw��"�ì<҈̹�"Oz���?v9�HX���vk��
�"OX��5jnM��X+/L�|y$"Om��Em!2����I;mҬ&"O���G)�:M��dˈE	�`�c"O�ũÜ�G�,�	7��?1��X�"OX��N�@}�Cː"��u�5"O�	0)K��@���F2�|��"O�Ah�%M�uRb�ˑ�A���0�"O,@��n�	JД��t�EL�e�!"Ou�# �{�V��c�6,�h`"O����M�Kv�����U�I���;�"OB���,�f��D�A-��u"O\�[f�: *���ׅŘ0�0Xkv"OBI�� �9(�$Q�t�Q� �Dh�"O�:3�^8cՊ��V���&ͻ�"O��"��#}��Ad%A� �x�C�"O,|�gmۦzC�1�Å,��e�(D�ds�����:`�f��:t
��j!D�<��)��)P�(7�ݥ���qU?D���0k (�,pa�i��{T����=D�THf�!);2P��� @�L���:D���Bm<(�H��Y����y.%D��Q�G/OF��f`�sg��-D���UF�q�����ԟ�|-
g�%D��3�n�!M�<���B�n����'D�����Ø;rї)928���'"D�,P���3�,�"�*ה!P���?D�d)֯�SY��Q���$p[��>D���"�/���`��1,ڐܛ"�'D����$H�X(
���'T+C?����/!D������r�.T�3�� ��(s�  D��a�2��`{3�S�D��-k5�<D��SV"�4U8���bnАfͰ��A�9D�� $�͇R�8L�4�ںHȆ�h6"O���d%z���� Q��9z�"O���cR6��4��$�*9��lbC"O�E�W�L�rT�&��!��-b"O��1��Q:5�x��`T�x�	q"Oa�C Y,�Eϋ�L<�PX"OL(���s��� � jݺb"O´B �,�P6����,Pa"O~8��Q1y�Hs��3�
\�A"O$Pi�➤M��PD�I�2p��"O� )���Gi��ĕ-�����"O�iX��̭:W\A�ǠO*�J�""O��X�	��j�]:g�_�[���!s"O����>� -����?a�:%�G"O	r�L �
��7f�$5�,M�E"O�Ⲃ\�w$�<��K�,��p#"O��C�KW��HRj��Z��Ց0"O�x��^��6	�-jqu�%"O8�C3���0p��g	�f-��"O�!qf�)'�v%��A4�"O��Y��_�_ ���P�^��@ W"O�����C!}�䩊�X��"O�lۂ��^���c�I�1� ժ�"O��CdM;nz4� �ܑQ��hY"O�3V����ICjJ�`��%��"O�q�ڂhx6�"�U}�\�J2"O �`j͹�D1Ch��S�P��"OZ��C	�_�ڥz��2$��q�"OP�G�D<o*��j!ݐ6���"O�釐,I��CA�Oj�q�s"O|���$�$�!��8��1A"O����c3 ��#�)pc�kק/D��X�K&)9) g�y��i��o#D����A�!t�(JU�ƚF���F�"D�|0'�̮i������E������
?D��Ҏ�6?����aD�oV�]�e�/D�d��)�c����*C�Fd|�B�-D�4��_�|�4��u�35W�8�+D�8�c�ӚtIJUAC�>�d��(D���ğ7*��h7�ϸ=��XP�;D� �M
5�x���j�|țs�;D�䘕	Z�(�
6���*�t�p@�5D��C� #!ޜѲ*D�)��z�.D�|4Eԃ�A�a$���F=��`8D�
G.��H�ʶO���̨�.!D�<���	q�D��ϔ7�p���1D��P)�T�&�&iv���W�"D�X��W!$��Y���;,r`��R�-D���U�),[0�	1�Z���0D�@R��W�����N��Y�dq�<D�|�V�!|nbı��[������&D��sm�yNJdKw*٢��9�W8D�k#���H"�(�	�J�F��5D������dqZ�I��x$x�2D�,@ ��5IW��x"�C�+
H����.D��8F*LB� 4���S��j�u*O
�V��e�'*��>�B�"O�9j��d?L	��NH)z� �F"Of�9�~�px�M�5D�tI0"Oz) c0���+ďM�(�*W"O���X�j����g��z���"O,��GI=>�J1A�GױY�,��Q"Oڜ��DD��D0���_��\۰"O|�	���)��0"�J4,�(�p�"O� l��Owj�؁���&�6D�3"O��0�F�=�z��@�FB���"OF��wgzYx��}=R��"O�p�9��T���M&/J8��"OFL� ��-����4��4O2��"Oxd���ÿ%34ڧ���+��@�"O`U���+f����Y3���"O�@�fQ�/!(�6�A�GR��1"O\т_��p�*�+x̱8B�ş�y2�,��˒�S��n<r��8�y"��4�I'�1a=Θ:��X��yb�R���Ɩ(%�d|�,ȓ�yB�ƛax�� �l0R,K�P>�yb�8>��EA5bCDMأNê�y�^�6����J�"ٌ���HH�<A���?�d���-N�4�(SX�<aE��;_T �u�ғ}Ֆia��LU�<�DkJ�f׌eڣ��s_n-I�dQ�<Q�,F�[L>)���X���`2�J�<�Sl��-��Sw��I� � D�<I�@=5I�qJ�A_47J�I���@�<��G؎|���Q�mV�lʪU��d�p�<1���@�����1D�����d�<4C�x�l�g�Ѫ(�4}3�LUd�<��H��lp�q�7D�7b���WW�<��bG�{�F}�*��=���EH�<1���5a�'�JT�i�OC�<�b �6X��� rLI�"��U�g#AB�<��d�58����4���_��Hs	~�<���Gv<M�K�F�z<�!�
O�<i���,JE!�n0P�y�dJ�<q���,"`�`%�x`��H�G�`�<�ՌK���#ѣw䚘бN\^�<y�%���8А"h4}�N\��h�\�<)`%�='�c e��MDIh@�p�<�g"R6(ؐ6�ަ&E|��&�e�<��b�Elp���L��6�V]k��L^�<��I5r
MS�
ɭwV�y�G@�<���@�\bFyWJK*'iܐ��aYr�<����k.��s@B��b=X�s框t�<a�O�@V P���̲6��Q��f�<�R��[M
�a�C�?���gD�_�<EI��k;��J6P��Hb��g�<��JՐw��넍R)G�d8��l�<�e��9��n�&d���9�e�<���5z#���'A� r_piY�FJ]�<)�L�(n��\��oJ"m<t�����N�<ar��0g���S���oZ����FHI�<mo�$�r[:�2�� !�D��v<�Yʡ�ۂW��Y���քQ�!�ē:zL,���J7t�"$Sb	��`v!��>sǲ�Q�̋�|����&(�=\!�$I�z|
�hE��(��K^y6���ȓ1F�%����r��z&�J[���Xu~a�s#YSK(����,K(,�ȓ `
���U������EC�t }��v�������@�2�� �"��`�ȓP3�8�2�0j8$�%C�合���^��'���ɘҪX03\�-��7sd��*D�3v�%j�Y8��ȓT� P9S^)�xD��*�%N|�ȓY*:�	$�N�
`��Du�<��ȓ�,1[�I��l<r��K�#,:��|<�ag�V`&J0�C��(YS(���S�? �A�]�d��m1��H/w�6�p"Op�s��Xai|X�`-�W͆���"O��z惥oYnl���ݻd]�K�"O��z�o��9�~]��+jl(@ �"Ot؃q�G�P��A���
T��A�"OHt,�>0�RX��4JJ�-�B"O���0j� 3!@��1-ޕO��H5"O099��L2,`ۅʞM��Q��'��I�3��64H #�i�5/�d��'��tF�a0U��\�񠑀�'d
h�d��=�}��lA�R�չ�'�D� �G2`𑍇$U��)�'��Mi���6ͤ0�1'[�	�*
�'>�E6���7$�i�/�!�\��'�V�����M��x��Ő7r��b�'����s�M�Z�D�U��)w��9`�'&�e���Tp����ԨANe��'+ƍȅi�Mz�ȳ��<8�����'����Tm
s��!���+��e��'^�(�j�[�^�ɣ.�0����	�'>�-�t��=>������3Zv���'����(֡|;04�
Q*�b�2���j� ��	�K��l�FE�s�<�'DWA�qR�� 4% �A�Ff�<��
?W�dAc�9���e�<AǦ4;J Ȱ�JYlL�����`�<����-��M�b�-��ȳ�(�s�<A�.;��aKf	�5d��S��D�<!cϜ�zy���� �2ծ�'}�<�U�іI�pa�6��M��5���u�<�DI���1E@ \��&��[�<i�Ϣm{�M���ar���#	\�<� ��6HV��'K�TH��[�<AFlK�
G ={C�7�ZQ�7�
Z�<a���/j���K���%TLy��)�W�<�c@1<��1$5D�r)j�C�n�<�W��
���Q$��\B�i�<�'�J�0I��.M��Hr��h�<�#Ǚt��`!��'N��e�נ�K�<��G�z!P�bT��-)��P��"�J�<iFҚ'��{f�ʧC��c'ƈ{�<�oT�E:�q�5�
ENF�s�!�n�<���*0|0���)�*Z�hXs��h�<)�(�C�޵C�L�(X����d�<!�.��q{��n@E$����UZ�<��� ~؜[�L�s������P�<�$&O�ʩI#MS~Zz=�K�<ٰ���4�D�o ��	D�<I�����z��'x �r $���yR�A1ۦ �F��L�n@a�-���y�(Xv��xu�D��Q�I
�y�@�{� Q[d!;��B����y�� 4F\��A�D�J�a�t��
�y��
nn��%��@u��+!&���y����6E�4g�$BЉP�!ϣ�y���0��Ed�n
5��,��y2��+�i;N����1��;�y�����lK7IF���JcI2�y�䈇t��@'`�U2�(���7�y"FO�y�8��B� I2�zbB��y©֖��T P�'��x����1�y2���2��ma�="1����*(�y���5�u����HY�׍̍�y2�3YF�8� �p���y
� 2�����86<�-�����J
l�8f"O����OR2�ܕH�Z(8�ܜyB"O����֦ �����;B�4ɩs"O�(��d�R��BF�Hx�u07"O�$�`�!{�5�2��&��R"ODd2�9K�EŊ�J����"Ob�������Y֎m��"Ox0HA�OK������I�Z�@A"O�X���A�d��n���&D��"O��@w��9L��\QD�c8��'�||`��<� �Tɢ���1�'H�0�B�$�;4ʛ���"�'�*���F�	 8ݰ��vƼ�Q�'_�TG���3~�؃D����
�'�*h0��Y��z���&,>@I�	�'����`_{�x<���D�n�J �	�'���t��!�~hi�3�|��
�'n�,ڑ�v<�e� �&E��'��D1(��>\"�gI�g(����'�xxRc��kVhY���P�_6H<�
�'8�ء�f
�2��(yf)a
�'#ڥK& ń����l��D�q	�'�\�P7
eN�E�D!�z� �'��,KϘ:l�LKc71.@i�'gV͢`�DN�R8 '��,���	�'Ȓ!�EI�P�>�8�L�4�����'��R� �F�)피-xbPp�'%�9�H�;3��
��@�{䌜
�'<F�� X�gR4)*1���u����'��|�n�9K��8 M�{�h�j�'�p��4.��K��L@҂�a�BD�'��pR�ˆomP�qhݠ0<xi�'�(��(�ji�C �%,&���'���[�&�^� =� ���g��d��'�u��)�*r������Ya��8�'t�$S�K� �T��վ>���'�,��� -|��%�� :IO��'"���5�z TY#Q&��j�Ҥh�'�,@(�n$:��b 	^�8bD��'2V��1푴��T" �H�\T�P�'Py�(�*z�"�E#(��5�
�'��)�կ�*8,��Ѹ��=s�'%a��ˋ? �i��lՑm`A�
�'��!C��Ml�aYЫ��^0<�
�'4����-ؕeN��;�S�XF8�Y
�'��-�ѩO2��zgj��kv��
�'��h�
({��mivF�w��
�'VJxiմ�*i!V��}���	�'�*In-P] ��̞f�5��'�,���&nFq�ĕah�6"O$�sgU99VU��l���!"O�� ��  6�D�l� ��z "OLyA���=���0��`��+u"O�yrT�V~������A{Q"O�� ��]��ѩPgS�!�]_�<�@�PЀ��7�G'k�����!�@�/2:d9TaM�?�|���!�D�:J�T�aG*�w0Q�°!�!��G�z��̙ ��)8hp�Rr�־y�!��*w�J����5�`]Q䤜�/�!�dT3G^�M�S�VP�^���1`e!��v�N0r�L�o�zi �DR!�d�`~����Ōp�ʴic��� �!�d�+7D5��K�r�tU)F�7h�!�� ���f"�_���`�JF)-�iYC"O�T�k��=������&�h]��"Ovh�g.�����˚=��v"O�����[�'A�	� � �(��"O���T�&	b�u�Ǉ�;BŤ�S'"O8e���	C<�S-�>����"O�I���E�eYP��l�2`���	�"O�٨To�k�A�AD48��qQ"O�ljRk�^ݢ�Y�v�B!q�"O�e����6l�V�!�P�i(NXT"O�m+Ι�f8N���	�R�X1��"O�=J�iY��T��g��+~�v�ٷ"O��fҹ:yD!ӳ��>	���
"O*�`0A� [�m9nZ��!"O�)j��^�?��ԂU����f���"Oj�V���C���B�ꖻ_><C"O��a�"K"Uh<Ф�2)<("�"OА e�����3���~�er "O��[f��,,��R%��6�d��"O��1V�=T�$�_�uŴ��"O6p��6*���ЫJQN�Ӕ"O��N�-=n���5���c"!�s"O�4z�e�,ef0�@���+��!p"O��Y��P@�u��D֟@��@�t"OBt*֬�(j���rdM�R~�@h1"O�"A�:$I�B)͜���"O��n�u��2%�V1�ּ��"O^x�p+�G�\\��V�%ߐ�4"O1���I�d��,4[�|�N�s3"Ot�bL�-'<�s�֧U�^5��"OZ����ݛ�fF�:��Jv"O�Ls���|O���=m|M��"O�k�B�*�Ārw��aN�x�"O�|��!ߖ1��)��-D�x�vUb "O�q32ޑU���͂"h����""O(�C��gҌ:����?ID�W"O�R��eh8B Ç:X�0� "ONu��Fʖ	&$��o��� �""O�%�@�R�	������֐_��x[$"Of���ίS�$0e��H�\��"O�P'�Z���0'�Iǎ�P"OP�8��B�#�)2e�.���"Or�h �N*"�I8e^�A�H0��"ON�("��$JD*a³��=-�&S"O�if P�F�*�Č���L-�yr��`!X�!���8N<!��oL��yb��8}�j�Y��G�D�LXר�y�[!5v�)��A6���`��yR�G'\��IB���e W��y"��"��=�E�|�Nj�cM �y��Q�U^�� ��?t��ْ�ʃ��y"�J4(�Uq)ُn�Ԑ�TJ��y�&�!Kt�!E�h�"��,5�yrc�Jcb�g�[6�m�Ĉ��y�hތdq8��W�N 4��ȴ�8�y�ݙ')��#A�A)Jv�`���y�$:%�hěT�NF/�i�mH��y��B<)�ʤ��E�8\��C�Ɗ�Py��<hT��;w�Ĳ	G�@��-N`�<ac��mk2ES��̨#l���.\�<��'#�0� rA�#sV>U���\\�<IB�Z�1��e��K�r�GVA�<)0a�+~#�Y�兜[c$\� �{�<i�E�/�>DP��I ]㊼��dJp�<� @}�"kV�4��͘g���p�pq�"O*@3F��yz��Z��;m�eɰ"Oy�����[�zeء!x�Q��"O�`�5#��G�W85��%F�ϱ�y�G�{�@��w"�(kD̪��.�y�Y8��S�n�1Wt� �yR��Df|1E��)D���7�=�y��-@]� I�DN�&'�S�����yR QBnB�T� �u���fG)�y�+��bwp�XqM�]�&8ˠ�!�y���2�n �Eą@���$���y�õ��۷�'��y{ԍ�y�N 1�F]�UC\�W$�c�O�yφ4.����F+.zt�SF�ybǉ�+Uty�0�B� �lRc�Ⱥ�y��G�t�r@�/^
#(B��2�y�CK5\�$�4�~�X1�'B��yr��-������3w�N�C�&���y� I&HN�yQmL�g4�,�6LB��yR�Q�.BPL����� �{����y2˄�I!�y��/D�u> Qf���y���+:x���.��Z��0�)�2�y2�	&*%�����c�Rd���N4�yr�8N7��qTK�b�L�`��ܠ�y��Y�O��#	���U���7�y��]�Tc�Q�r&мD��!���y�d��1Ʉa���a����M�y2��N�\T����-~4 `�&�S7�yr#O�q�b��)ZẍuÖkR��y���;�R��دY�TA��3�y���0c^� ��9P��AZ��Û�y�"صdon`��G���{��$�y�D@k|��B?��0�@�-�y҄�e0`�[E�
t<��g/���y�%͑q�j�!#e[�V�	2G�^�y�m�V�Ztz���H��T��G���y� L	;�T+�
X$EK��q�K�#�yC�)�<�RRI؝o�li#,�y���LE^�D �*bF�!�ՃR��y��0Q��1����Y���R@��yR�ǜJ�y�i)��2���'�y�aW	P��頧��Di;�O��ybL̨7]D��'��c�A��y�!N� ƘѤl�9~ap��!H��y£�rv�mH�L��_��\!!)��yҧ�
9�Pe�S(��h��=�y���8<ݐH�!�ш0������y"��T.-�Q"0.q���v�S��y��5�H��1�T�<��c�O�<1 b�"\*��W��z!��8&HK�<! �V0u�vTj��%��їK^�<�cb�X�DDpR-Z�k�и��Ir�<!s!6,�\$�CGE0����#$�k�<Ih"B�^\J!���f���7�yB 'oo�P�@��U��.�y��BBqܡ���֨.�٩ӡ��yB�$�D܈ħS"��s�P�y"/D�i�\���lR9+��˂i��y�[�h�!2�j#�HY�ś��y���G��jӪ����IB���y"C�7:'�thd�&N4�x��Ֆ�y�`�e���a� ��IBWCZ��y�OKW?>�(тA�:�i�-�y�FI�(GTĸa��{7F�QW돍�y
� �)Ę�^0f�a�h��.tZ��B"O^Ȋ���KB��rc�ȋM�c"Orq L�!�b�EG�fH�"O.�s��):��� �ǭu��Ȁ�"O�ۄ�]N�v��WgҘG����"O�uA�H�7v+f�[`��;Jv����"O��z�I%Q�N�9󌂇7N|Y�"O.��S��-r \)@#kWPA�؂�"O�	qpѡ4��	�R0+
��1"O��#E�U ���F�J�z��"OF� ��?��%��X�4:�X�"O�9	2��7T��A����; ��U"ORy)A� %�4ِm�>�h�"O��"��F�\�z�Í�>r���"O�(�a���\�Mm>�"O��B #��V���$P�H�"���"O�Tbtf/4���QK������"O���ƈ�w�1���I�^�2�zF"OT�����'5p�i[1~���2�"Of��F��U8Wk�;�`���"O��)�ķ}Tӓ��<w�Q{�"O�C����6�&����"dH�Cb"Ozuh�B���i��I��K��)��*O��&  3.�D�cB�!`ڡZ�'�zH#���Uβ�02M���2�ۉ�4�	XV(XwO)�@9c�┉���ȓ\	jL�W&�q��M��_A@U�ȓ.2��* ,�,ie~E �A�n���e/8kJ9_�X���&��Q��d"?����"W*e��$O54a�(W��0fv!�$��V�<�6B�
>ʴ�5�Z56?��d1�S�d�38��(�ǚ�/| ;�
X��yB-�
ȴ��Т�COdY�@'���y"�V<���9s�6 � %���yr�A�m10yJ��ճW�-R����?Q�'�r��㇛�+�P�1e)�Mr��	�'�hd��ն���!S).�b�	��hO2�!QdZ�f��1�5,�.[V�Y[3"O�A*���MI�JZ���`�i�ў"~n�7��Hq��!�F�2U%[���B�Ifƴ�!�RwDݘ�(M�6�j���������
�� �f�,h�D����3	@� �O��"D owƐۓJ��;����g���vN��HD�.�bu�ӮٳD��{����I�+q��J����!A ��!\ +�l�s��)�矘Se���>��$��b_0E ���d5�	y���)�O��"t��-ڄ4�՚w�P�`��O����6W<�: H��[�`:��R(Gga}��>I6�n��Y�F6U!*�[�#�\�<%��r�"y�U2E� �
A�KP��hO�O
e#���	l��գ��Q����'�����Q��y�P��K�q8�'�L��懬-�~D`�NE�B ����/}r^������Ц��5=b�Dܭ9�v�B����#Tu�&Q�Ne�p$>O�"=�w"�:�2P����&k��\Q��N�<9!�Z4DiNA�X+2|<y������;��i�a���>�ص�I�W�����8�A��Q'y����n�#	���ȓ5-�[��V(l�e@Ԍ��1����ȓP6ˠ�@*T:��s	g	�rm#D���2���v#�ps��"b	���+D��bP��~�d��� �l�.�;�,>D�܀�*�78���Ch��$;,����<�<�S�g�? ��٥� ��)x�G��X�TI�"O�H��V4�zq@� ك�(IH�"OT� #��"<BJ	xS/K}�tK"O�|���� su^q�5RaVHSu"Oz��=Q���UB�q��K�"O\��4.M�
����gԗ��D"O���&H�"u"�0���F1:������_X��+#�69�|u��%�<���xu�3D���d���h�`��c2��:@&D�h�Kկ
�� 0��^yt�2��$�$2�	`̧�?�K�Nd:��n@�5-t��g��:i�B�I!d�H]0�c���>��6�\�(+B�	P����p"C�OA����U��C�ɴ[!t�$��3<H΅Y1�� P���?�HO�>apGnɗS�\�� N�76���,0D��r0�M�}i��7�-lu֐ �A.D�p���E��<�� E[c�|˵�(<O�"<A���
��(�vˊ���Ș��t�<Q�&MⰩ�gY.D�Z��gHs�<yG��e|����)m�n�#KKm��<�<�t�6D@��S�@]�N���E�Tl�<���N�oӚ�+q�T";;�x�#
T�<����N�d\��]&dMhY���R�<��K�oYP���I�\��i0D�L�<u�ЧDb`�P�F#K���ȓG`�Y��M�h�ðj�(�^<�ȓ@��xȥ L�f���d�j�ɇȓ4�x%JG͚�eW�Ѩ�hQ:���'���D�����7I����##�	W%��Q��&es!���P��p�Rn��W9����']!�d)e�4("D�=m��e���L���D�$+U?#F�q@�нt5�`�����y�oܛ�> ��a�!�ݙ�����y�kg�<:3�J����T/N+�yRĜ>ĴL!	٠ZX�5�A��PyBb�c_`E��H[�D�����D�<���9<�0$aC�>OT��.������z�"�Yр,a/v��p������:f~	����7�A��%D�Mf����[�"	�`��x�d-�$�A;a�X��ȓ[�phU虓N�j���A�� �Zh�ȓ8>����U7CQ�)ґ	�$Zp(����
'ў�}
AeΒs�$ل��K��c�D�g؟$KW�'�@��D�A�����:'R.�ˏ��6O�)��ςyɾ��N�M=:(�q�	u�Oi�b��#��%8r��j=Z1�'T@���
�"T�@A�3XCP�*���If����H�4��ʑ�� DB�	1\=��bB�J�m"d0�j 0".B�	?N�H	�p�ej&�x��C���C�ɳo�P��bnތ	�"��FA?Q��C�I�gצ\�'$5{D�Ёe�K�m����4�ɦR9Zq�\\��[��;�6�,�S��M���
�]K�Ч�
��P�KR�<���z����D�/N�D�Bqˁ�E����(�ɦ*F�BgD��p*�#T�[ ��C�5N���+�/��d!�&jא}�B�	�x���.�ԐG��C}�B�Ʌ���'�Ԁp� �Wl��.L�C�I9�����DmTC�'��Iq"OH!	�8"r�X��1р�"O0�a�N�)��eV*V&J����O���W�rD��"@ӑm�`�rFe�t�IQ����Հ�8�QjT�Di�x�8S@.���)� ���D��T���hc@�;��f�O�b�PF{�������0z�R� �ѽm,`zg"O��(��(8Z��Ε�h).|Qg"O��r��>B�| ���(B�;T�$G{�剂"/aZg�ߪ��H$�
��B�	�[��R"�u��P��I�m�2��^؟�YuoT u�n�bK� �F ��� ړ����Dh�h#�Zs�"uy���As<)��<1��哝	6Fi(��T��Ih�O�
lB�I6A��Qc��
!���C+mƞB�	"{}vI�cC�@"�(��ܷ3�h��hOQ>��pdԥ{��)D�_�^r0��#D�dz��U=�@yS+���ͫgj�E8��Ez���0�")"�/�$��Q	��
�y2@�:_n����G��c���M��'�̠3ת�n���P�D�QM�H	�����Gv!��J=�I�
րvB!���,i읺�m�8�șa�ɀ�E:!�D�?�*p� m� �h��c��8*!��:q�L	[$���.���&�Z�6!�DV�o5TaR�.C�{��<"�CM!���4�T)3�E��H��)�v�Ҿ����7�S�O����㟩��DDG$*'،#�"O�A�`n���~p�'��*vig"O��&�;MV橸��G�%=l�ۖ"O
���X3���`�OIW�N,c�"O(��^,`~��c�DϮhhz�Z6"O��؜��� g�ʇn_�}B""Ofh�@�»},DB1]WJe��"Oj��g$^H�ڣ�פ9:Ir1"O������Z��Pcq@�%M�΁K�"O| ZQC32���(�R5�1�s"O0p�EEAg��˗�`���x""O��:�DS
n��:@aW�P��sB"O6Se�h���oR�o�v��R"O�Hȓ#��f$��F�I�S��@ڔ"O�PB0#=R�Pq�CޖF;$Uz "Ob����[�V�Li��6A2�qs�"O�K�������v&�(yv"O�� �XGʕ���T����"O���w�ƅ�����5���"O��)W�D��5��'
d�ȓW=L��b�I�L����[B,�,��r8�	��.�B�`�;��ȓO
��t��d�5y��N�U��=��qo.���@�P�8�̅�eu�ąȓ&} ���N� ���ʀ�D�ȓ¶�	�ޗL3xA��KGl��a���ヅ��A�tꙃ@2D�ȓBt���s�Z�\��p;#*�-Ƞ��ȓl�:E�F�[P�mk󯐪jn�ȓ[�h�IB�+?UXY�v�')s�ć�/��U�e�	��-�!2�й�ȓK�tQ;�	&;ʅRE��$8^��ȓ:D�a����J���p�C�PP�h�ȓ��ɓtE���� �$�x��4�5H�`�nE�IZ��O��!��2+tUb�f�Sn��ȓjV���	ə3h�dPf刿ފ���DTT	�����<v��4, �ȓB�*`�a&��
�L�t!�d͔E�<����	cyS�Låi|��`�g�D����5�ўUF��i���,�Q�ȓY�����Un��I�V�&Q�Lȅȓ(R�HJr�[;6���rV�����S�? �t2�I�\Q�G�E�0���"O��Xb�	8\�l�âU�Q�dj�"O�rG)_�Uc�Œ#!�K0�ՑB"O�uZ���?Z��@�k�.$��"O�}8�O�J�ʬ`�
O(j:r�`!"O^A)��]��D�f�҆`-Ԉ�"O*�ѳ+��3/��1�]"1zy�e"O�qhG��&z>�pD���␉#"Oܰ1c��m=�`�E�!<�i�"OB ���¬���E� ,w
�;�"O��:�ßMa�!	1�1R|Te�"OD(#�[�^�(4�d��;2�"%f"O�$T4z���JsB̕�ex�"Oܜ���,NR�p���tȜ�QR"O��C�ʂ_*H�灋8U^	�S"O��(Q��,^<p��1x���"O���u�ۭ�8@�w!�"O��D�4"Oh��̎�k!����Rh㐔[S"Oj-�Ud��xQ�φ�R�b���"O�PZR)�;'JhIs�HAS���z�"ORpqb�]'��Py&홱d>�R�"O��s)G)~05A�mK*te��A�"O*}bA�Ϻn���2`%Ä^Z`Z�"O�6�J�9.P5q�/^�4rh�d"O�tSB�771LM@E�-%>�V"Oh����9g�B�AG�^�tI�m�"O�0avE��]� ���r	I� "O<#C�ܯh����%�%6����"O�Iӡaù#����� #&~t�"O��Hĉ��H��F�H�ur�"O:	9�E'0V�2�cCt���"O������-D���A3(���"O�)��# H���)��q�����"O�P���*B�,�+rmԯ*|l�{�"O�x�+�;	��\��È�[���s"O�!���=f��u�B\n_���"O$@�����AR�@)��R"O��d��7|^�s��*h�H�"O")�u�+J^8Z�N��y���x4"O@�D석#�ZB�="Kdh�"O.ѡcA�p3P0SGd�3o�P�"O�� �"�1H�A�3%���S "O��V���flze���}_X��"O�02�'"t��E!� ʹ�ۢ"ONa�U)	�"g�؞}rҭ��"O(P�#.[��M`���<����"Ox�0�b�~��""V�:˸�q�"Ob�3��Gs��TC�l֑%���3"On����M�Q���G#r���"O��xw�;kЕ�!\�|�E��"O���t�p/��CG�'[:��"OF|���G2�8:�c�4ml̸��"O6e X�x�Q�VA�%[j�I�"O����K+B�\ٓv�H�(8R�I�"O����V�XMvl�"�٥R��*�"O4���o[5f��k��B�:P2�"�"O�\Q��W3+P��؅��0yQ�͈#"O�Š��^)Q��u��&Ј(vD`x�"O�\�7�D?ha#V�Z2A0�p�"O��SfI�#����̖D�Xdp�"O�YY��)Q���Bg\�NR�ar"O����I]3���ש��Go>�"O`}�#�>E"�X&�P0|&Ta)q"O�(9����p>�
�'9s6�	�"O� $�*ELC+\U�G�0�"P�v"O�����G3\�n�0�Ӊ%_�Q�k���|<˵���O���u�]y�e�v#�8d�19"O��c@�ĀlQ5!^�"N"���'uH��P�T����?=����ڎ\a*l%(�)y&�{�6S����7"?<�X��u�\�k�J �@R��k#D�,���Ѽ���޹eu�QPS�>;� �6����̘��Ӯ8�P*7�+|��=c�̀Zt�C�I/"����C�HQ�%� ���غ�B��UX6�$e���ؖ�<��b�ZꦘhUGU9]�h0i%M�O�<�ց(9��`aDN2s�Z9�c,ҽl���Sj�#J�w-��<��Mc	��:�����L$Ӧ`�x��хւo,�Y�i��fj�t��e�2!�BOƈdE2a���wh<	����q� �s�dD�Ci�r�nX� d*65�U����O�P���舩��td����'� &��@����j�#v����$a�g]�QZT_�ϝ�����6J.�	: j֧m6�q�f�w�.C�ɻS&#4'T�r�\5C��ßJ3��`�B2GxXaB'�T�G�>�特da��ڗ�ƂA
r|iÃk���D�?����0P�=#C�M��""ƒ�K K��Af�	�O��P�)֖a|���Z0ްq0e��0۾Qx� ڋA�ly9F !�S�h���1fE1q�]2���h�B䉕,#���� �Q�*Ԝ��@�b�uS�e�AA��T4�<q�B��{�
Ī1�'gs�U��(I\�<qUcZ� ��]��c�!r{�1���X#W4�))�)�I8��'\c�����a�dT	cFѺ6��D
E!2lO� B���J�"T��#Äf�A" '��kj8*���iG��)�A[C$��P�NT{�eϑK���?1R� �3Q4L���(�'��5���B�v�8�"f �r����ȓ�n�[��(�p�9v�\j=����V�D���=E�����[�B�&m��S�%�:D�<�T͌�5N�C�ĭ��,�d�;D��A`�=���z����Y� 6D�tP1��A��=Kƃ�]��r�c;D���-Q�v���sELݟ8� i�a;D�awo%m��iUD�I�QX�b,D�����0���S�+K,tD��s�,D�ܨ�lz����-�<�|����1D�`���ߩ{Vrt��E�,]sD�-D��q�Y�Y���Lϱ*$ �%*D����T�Jq�R�*/,���)D�����$��)�I����c�3D���!��xQi��Z��ʅz��.D���VN��N��� �O׼nv����,D�@��ǆ3(}t��P�\&\���%9D���ǚ4�U��g�-}�X:F/9D���E@7"L4hC!£aˤ���*D��0����P�i��J\Z��)D�S�D�rԘ���z�vip1�-D�$���
).u<����,ِ8T�'D��{�k�9߀ٲM�)�| cf�$D���4�\,{�u�pk׃�@\
"�#D�K�j���m��Ò�jU�>D�`�W	\�Rl�PPl��%K�)�E�+D���"농:)N� WlO�ԹA�N(D�,Y���[f��f���p\0g�(D��p�"بO�~�#�K J�t�G�8D��87O�0"b��X�`4�&��	7D���&��TrD��Uև�����&D�$kE��|����a��	{��ւ&D��D�ǒi�@��щ���}PM$D��qkԝ#��]K��]0�}9�m9D�tE�}�q�G�֠n>pIɐ�9D�\��R��:L�艣��:D�� �N@���@�k�8
��"�"O� Z�Ŕr�왕C<��-y$"O�$�)�X��z �UA���K�"O~-+q���:u37�@*F�ի�"Of�jwmwb��ㄐ���` "O ��ET�z(���A�a(Q�|���ɓ]`Sq��=�$�A� �!�$[����JSԓ<������^	Ӱ�=E��'괰�2�9�4I3�Y 6x�z�'Ls��	B�2|J7eٶ�'��j
�N�����߱h����P���0>iL>����%E�d	��Q64r>x@B�D�<�s�8uz[t��$�0׌TC�<�elY2	T,T8r)�+4�0�/ E�<�`IߖO�b�apH�;[�DR4�GN�<�C��pX��Μ$��͘�,�I�<��I�7?�4�'#����t*�	I�<�cCRi�@�`&�>A�r8Z`�y�<AA'��HZYV`V56�y���w�<q�jӃ|r^Ly�IP��|��Aes�<���J;G�=���:�}���s�<	�H�21S�W.+���2�[j�	�]T"#<�~�S ��x?�(`���7�'B$C�I?�v0i�N��E$�X�&ŎEf�㟠ȑ�'Z���&B%`>q���I&	�5;�'ZZI"��7	����O2p�Y�O�����^��-��H#_R�� �'
�O��a��)tt@�b�5 	�"Obd�%	�%Dڽ�'�P�
c�K�y�?~�^	�@ǔ�^���pG0�y©C(_�^����M=Nu���/�y��ҏs>ȭT*Q=����GD�&�ybbR0jdvL�3�	aW�@����y�Y�+j�4�K�g�<9�G
�y�MY%��٥eYS�ڴP�%'�y��A�J��i�$(ڐN�ha�bF���y�d){ʬ�Г�+w�ֱQ��
�y�B��}��d�;x�6tqD"��y��0M���R�����l��ӯȿ�y2���T�n�8#�	
���Z���y�Iߒ�
���J��x����R�F �y��B<A�<�6eA�{�Hh�����y��-U��"�	�|��)�(��Py(�9y�P(�%ț>P&f�Bl�X�<��
5/sZ@3񄔖5�H��C�<1�F�L&�00������tM�{�<)�Oפ`�rѻ�O�+�H��J�<1�%��t��#h�����{�<y���ઑq���z�� �%�[�<I`A
T�d��C č!‹���M�<1ꆁx��� �����$���!I�<�� �\���j��*O���I�J�<	¥���q%	֜;VPɊs�@�<1�+��`�oF�Xvv�W�k�<�'�^�}4�p��0�I�0�]�<)�k^�����@c�k6T�)&��_�<�CjW����R"
���#�S�<��ꅹxB���Á�&�MP �r�<� �Y�nK@��g�H������Z�<Y���3z�a���ђ�̡KB�W�<�PI �H�ɥ�Vo��5Sp�J�<��O�|�9ʓKF�bv1;�IA�<�d��@��P��8��,�RMX}�<ɲ��w�<�K��̕'��t�*Cu�<� �D�(�hH U�G��RP��"O�1�6��.�j�{s)܆b<F�"�"O�i��\�I�"P8u�Õ4h��"O^��vf�9MU�5Q�Nb�LX"O���c�6*��ˡ!��6p ��"O4͘�l��v�P�Z2V�"O���צ�-]=�bKҳ)�aI6"O�J��d �	�B��8)pp�Q�"OX�5�C!�Q��+��q"O|Hs�K��*0G#^�֜�"Of� �j�QKP�2����"�  C"O�Q��铯|f�F��.Q�\�7"O
�%�x��jC��2gT*���"O$��L�@!�X &�ɊF10�"Ov��K��c�xjfeQ�pL��`"O�mZ�;�Zbcߛ]R��"O����S]�Pq2`ւm��H�"O��+EI�4|zi��E��.X�W"O~��D!_*� ��d�<���	�"O���I�d������]�lB��"O�����8f��r ��$���"O���5*́c`����Z�cs���0"O��"F�u��Г�+#�D� �"O ��e�	0��Q3Nek2��"Ov`Oۿ����EkZ�vT����"O�����0[�`W�Ѐ	[���"O*=�Rg��<��5i�X%�e��"O�0Z�fS�1�d��шP�:�6yF"O�PHw�8�j�e��$�����"O0����;��1�v�I'^�v�$"O�H��N�+01L(5h�pTB���"OXt0�.я2���BGN+&@�$0"O.mb �I�w��x������"Ol����I�RdI�T��D��8s�"O�Ԑb	�]*Ȋs���9��!�"O��S��.:�T��ȵD�$az"OL,+�c�����Á��@����"O\���E�j�� j�4��]�"O�uqN5<+j��T<{rx��"O�e�V�r|Bf�ѬS���%"O�p�a��h���ƨƲ�Ε w"O�IS&cV(M�Zi���G�8h���"Oґ����IBL��ϐ�vn�� a"O��;��ja�/�'\��)�6��)�!�DX�o�����
ɂ`٨�����,z!���p��������`]�.ԶYs!�D@�n�:ؚ��\�[�txH'��[!�İ bh(�A��|<�1P���:H�!�DG�	|�Y#pJ�/*�HU�H��!��%J�>L�V�1�d�O 5�!�8{툑�ե��W�����}�!��;E���3``�,qf�i���k�!�dr��a��f�7a(���KF�!����q���O�k�t� U
��!�D� *�Y2��Cx�	R jM,<�!�WNJ�����֜\6�\����(!�$�|��UXU��,Ҡ���1!�E$�V��1Q��L3!�	F>`$r�fQ�[㞙!�e�3�!��*)�h9�� c�f`ʗ� ��!�D��Z� �h7l�5�,��eϮ�!�҃F�ڄ�%��(��C׈ �S!��ʋ �pI��3|�6Pˆ钅^/!��v����)�z��§��m!�� "9�p&S�FE�����ȯgix�2w"O�ɱ��;Xj���T�]N "�"O@��"��l����	�`"O*�p�拱H�F���L}����"OpL@ ]�[o�%!��چXP��"O�ERf�U+&��uaJ�,��L��"O°Q%�G�jmҨ��I��t���"O��P穖�V�,p�b�N�p�"ODu���^�Ҕ�W<���%"Ot�0A���8�.�;1ٴ}��"O�P���8��킳���'"O��Еh�k|� �.7�F���"O$@ �ED�U���j7�<S"O�� R�;��Z�j��qL��HT"Od��fG�;Ls `�i̇%@�a�"O~��ŉA=���Q�hT�ސ�6"O ��O����X6D�`�"O���E�lߖ�$$ !$%D��"O�uxCk=L{�����'`�I`w"OD��G�.9��-���ԭ(��G"O"�E�<�HY����0��<u"O�T �'5�|`Di��H�"OhTSBL$d�eh]�A�v �"O$� b�oǂ���lO�d��� "O 	�&�4M�@�Y@�D!Wp�L�r"O�$��Fݜt�"!�R	ۭ*��]"O,ջR����Yk�ȭ8��4�@"O�y�@�8}��U�xrb���"Op|d�P�w�hH裬Z�qa5b'"O����ɬ���[�Y�qX�"O$5Y�ϔ�����
F%}�q"O��"/7��Qgʁa�H	:�"O<[F��RH�u��IB���W�yҡԛ�f@��O��:�
$:���yr�H)g�B�2��ߋ>�I�teU�y�G�V
���͉�,Fh��`I�y���84st4��œ)��e�$ᙈ�yB�1E�t! �F�)�0:�h���yB�A9�օH3(-/�9��H��yb�p%>aUH�"&��i�AK���y�@�C|��˵�+^��R!����y��Eh�ȉx�e���Z�L�/�y�Y�m=Nps�
���c%��yg� ��H(B%���f �y�
��� �ɸr0�dr�hC�y��ǻK���3���hx^�W(�=�y*�+h�hRw)��a
@�V ٱ�y2�ցGf6����U�5FnP��� �yR�F�D��\ �cϦ6�N�c�i[��y2̅�vq�!�ц0<��1�J�yB�]=<@E����;�4�؀���yB#��4w"��%��x���	�-�yB�Ò.�<����n؊��0�Ͼ�y�"U��*�j��a�T�者Y��y"�\�l(�Hb%��c
��'����y��Z.0¦�p0�
5\X�HJ�$K��y�o@3T��zwmY	P� I*UM��yR��.1��ǅ�K�uP�n�	�y�� kF������"A�M۰����yR�ٟr�D�W�=9�bp� �'�r�Q��שLU\��ȇ}����
�'�
�hgm!~�>HZ���m����	�'�ށ�D��Y�8����H�\�|�I�'�Ь��!�/	���+$���h��� �a���?*r	!T�өDK��V"O�%�&�P�����M�6#M���4"O�4��a$���8��9t�9�d"O6����,b	+���+O��U�c"Or����QbHZA���58��@B"OD��I�-b��tCHQ$đ{�"O|e����iv������
���r�"O
@�3�B=] pQZ��ތԜ�!1"O.�C�MP!gr��#�D� �t�"Od��ۈ"���y�xƒ��B"Oh0��ي#�`�BU�.�^���"O�tYCm	�$�hi����0H,�"O%p�[�i�j=�T�� a8�bw"O�� ���<�& �U��
��)�'!����2$0�͈�7?��a�'�|	��MҪ'�(iP�e	pwB�k�'�H5#����l�jY�&�LjE��b�'��y�oɛ7��z�NڮY4q��'��+TK�����������'��$���֘/ލbS��/����'Z���E �7Zr�}q#�[�$�r��
�'�PD8������@I
�'-jH���[�4͔�2�T��j�Q�'��9����?[dD�f��s�d�)�'�����ꚦs�n9��u�,�z�'b�(�奊Ȇec2D-3�$���'V�=d,ʫnr-A�P-0`���'��M�Q�����s���yʬX#	�'�M�4��0Z{,���mNi�'_�P�WBՓXe股ӵTO D�
�'Ʈ�;��U#M�v��$��7W����'��ѩe�' ��`&�,@��#�'v)Rf �=!]��pEӤ$�H3�'ΘBT�ɩ$>ɠd�߀$0�Y�	�'�(�X���>��U��`9�&��'XRE���N,(#Jl�u�_4p��,8�'������ �d�Eg�{:V���'¬]��ס�K%�[�i�@<��'�b�O�l�>%k�jV(`u|�	�'Ѫ���X!;��P�OU,s*��x	�'����N3!#�I��Fh ̀�'�Ģ7%��)NѨ`�ɵm�J!��'�\��Z$n�e�֊ݝf����'?�L��'���@VY"!H�'X-2 h��z�J���o����A�'Sp [���9K��x2�X�'��DA��:#T��$.�	�ͳ�'���K��نs�DP�hސ��#�'O*x�u�K1,m��Cژv(Y�'�0��
ZV�F �㌵]t���'9 mH��3I���+r�j\uB�'&Y��K9�`$��IF�\���'��)סV(V�. 8��h2(��'^ԉjf�h�y[�H��X3�'�Ni�e�f�Pp�H�<͓
�'��iw���eT ��gꒄ6f<!
�'0H���<[R�*�"�<&����	�'wx@��B��;���hŬL )Y�t
�'2�9E�ݨ^�N
�˝�+� �Z
�'h� �d�;X>@���ۗ"5��!	�'^�Q"K;6¦��#�A1w9քP�'d�m��d��H6Y�)�,i�L��
�'浩�Đ�4<p�0��e����	�'H�r���4�L"�o�8PA�4���� �ᚦiC�X�X}�O�H��YЅ"O��
�F
��Di�đ.��b�"Ob|0X �SDfY�%��vh�V�<IC�́9�dX'-د�j�1���P�<)Cf³��9S"ب�P��_Y̓�h��ޚ5j:+Q�_�4+���<�E�ܱW��!V�]�!������T}B�'�Ѳ���"�H� Ǽ@� �����hOQ?���B�+8�.��� ��Ѐ�>ړ�0|���B�:.��ª>F1
����z���hO�'���c��D�5�䴻�"�Y&x'��G{��DE]�
���iU��
s�z :�����<1��0|ڰOK!|�9Sm�N�Бq�L�&�ԅ�	�Px�"S-ޚ[ *б�K�O���Dl�$
��xN���Fȁ=_�~� ah>��O����9YM����L� �t�HOcΓO�=�}2`"]�uI�GY�N6�����Oy��)�':@h�+@$,H�`x�pŅVN �ȓ;Z}82��)'�Q�,ՋDàM����<1��H2a��H;SlJ2~�dy��m��hO�'n��M�������⎕���/��<�S�'u!�a��f wA�sO#�`U�'�ў�|��QF�1ۢмc�� �B�Q�<Q��Y�l!��鈮n���tPcy��'��	c>�"�@N/]q<�2��$0�C��<�(O�=���9���Ӣ@�p�5C=�ʴ@Н|"�)�'Q�E���Z/)b4�V^�U����hOQ>����M��� �mCM��P��Oޢ=E���ۦ")�	P2�2���'E �hO���D�6 p⵬A�>-US�i�Q5Q�\D|2�ƶ*l����4Q�����
}��p�'(D�l����#r��pyW��7&!X��&D���j�L��`�MZ��<ȵ%D��Z� I��rO�{��8�O$D���r��QҜ�B�AD�.Xn�s�&D���	�+?mvE�`�D~�*�;C�#D��1ac@�T�e���3��x(#D�+���V�8���,7?���'�6D�ı�D݇& ��r�PL�`� ��>D���R q��M�p�Q$.� ���8D�H8 b2w��,BBS�!��%��8D������!���DcѮ���32&2D��A�%�-qv�۔AO-��Bq�1D�@آ�ݮ�`�(�
�yc7�0D���!��l^�U�i3����,D����� %	PP��F2�5�1&-D���s�S�^�i*����w��z��,D���FV���B� 80�ܠ�-D�P[�`��|]�=��hY�	[p!�*D��i�.l��6����(D����),@k��&F�->nhT��f&D�l�#/�5�+!���1�TtR#D�$!�^훤�ښv��# D�TA ��R��s�m�	�tQ���>D����`V
]$���#��1C�<D���A@}:�{VBY6�`aZb7D� ����^��qH��$8���A4D����D��4����s�<�$$?D�,s ��9�����Ɂk�r�x��1D�h�0�^8D���!%��h�i3�+D�<���L�l(�� EG��+d$D��#E� ,>���#w��a�4/.D��Q��٧
�F�if�!�'m*D�l�w���Yh�UI�Jp�s*$D��J�!�	7�\1b�H��<lY@%D�� �y�g�Y�xx(��ԐR�"O^����ϕ4\v��G�=[�0@"O��r��9�>iYr��8�x��"O�}y�����@ש���� V"OP�nC�L_Tq�	[��hXٳ"O�Q��H�2.��(ۇ0���"Ob��,^�{d�	�3*�E����"O�up@'X�l��Q�
�?ItM`�"O6����"+����ᩎ�W�İ�"Ojh�$*5Ȫx;�'�&�I�f"O ��*N�����e������"O�� /��zԞS����;&|�"Oz�� H�v���g��,x�V�r�"O��ʰ!Q�j�
��S�
ٸ�"O�x�A�H�0e�����>R�)C"O@ER7�Ӵ��Oĕ��"O��A!��.6��t��%}Jl���"O�a��Iׂq��ɀ.ɘ/́3�"O𨻇��&2���M_+%�A��"O>]�0Ć�9�����'T�r�"O�M�  �^a�MC��Y��$�"O���n��v-�RJ�
"�L�"O`a@���=8����6��h�}��"O,A��ŗ �"Y *зa��c"O��h%IY�C�pP�*G/dh��`"O�L����k.|A�ת�Y�U�"O��4+οK�`8g�F,�����"O�x�ע�>	N���=1k����"O�E�D	�Wj�h�̈SWRٙ"O�\˔��n�����+����s6"O���"�6a�r�h�=���ѣ*O�(` �W�2��DٓHJ=H���'u���'bW�~x�C��2	����'K�(����1b�Dj��	;^�%��'�����̄�����(,�Dec�'��l5�A�X�$�Q@�&����'�&��@A"42��(%�U0���z�'�l��tLC2$�$;8�t8	�'�aY��>1" a]h.���'�U17��63`�$��d�<���;�'��Y{�P�$��t�H�}> ��'����Iҏ(�"#CI,,*<@�'A4�Pb ��/���z�h�'��t��!~8��c�C��L9s�'6Z�����SǺ�a��:r�4�R�'
V$�@MH�.H�A� ɚ5k>���
�'�Ή��̯>������VX�0P2
�'���G,S�ݸ��!�Z���'����
ér��Q��eL(!Q�X��'�~١�],z�9��ƆD����'����%��|j*;�+���'m�E�"l�4zŮ�{hZ�]�i�
�'E@��w��Y}l�����}����'�4�1�×}��q���sۘѻ�'DB��"Ƞ$�zD��:{�*J	�'�	������.�F��L��'Z��P��Q��r��۪9Ȕ�z�'g�m8�T5Z���B��j(��'G�e�C��gV|��B�%?T��'�P|R� +7��iqfC�����Py�d,ͨ|�fBP�&�8��D�e�<����Y��8u��s1��g��f�<�ǡ�1�&ĚҩxWZ`�@�We�<����2|ّe
�8HC&)ef�\�<� ��J�gԉQ��j�cOi����"O�u�t��4QD���"��z�B(�A"O̸zvf������RE�K�����"O����˹+x�
2���T�"Ov�m@Se*�j3 	�hת8�P"O�q	�MB�u2R����ܿ6�T��"Oi��)E�
έ�V��7j��e#&*O*:� 
�w����G:�� �'ºЩRJЩB�\i����?/���*�'7�)�̚(�nlQ���.ZZl:�'�TEJ*oUڱ��aƧq#訳�'�Z��h���Ă�6��;�'�,E�g�(�传r��).��a��'� S>�U�EH�,B^��'�ҍ$��!=��
ɽQ�(��'��IIs+_��fYP%O�N���
�'тW��YkT�p1"��iY`��WJ)D����Ėmk��Cb��*
X���:D�(0�܆6-"T�c�ɜMU�H���7D������1)�B�`� �\����4D��`p��8˴y��*Da6�c�3D�Y�l�=����P���a�$#<D��z���f��lJ^)Rx)B`:D��x 	��_�`h���c���ą6D��97���fƸ�q)��cꨕ�&� D��BG׏ĺ���#kn@��>D����Odn*�BV���XЂF)D��+�ʇ�;>� ��
�83�C�B;D�,����$����G�{�.-���7D���f��[�x��En�9��2�5D��x��Ĉ"���!E$�

����L!D��B���R�(���,ŲH{,����,D�p�׍�O�2ii4�B�)�L]��?D��!B猑�\xjW垤C�>��b�>D����݅3�!qV"]��<���<D�y �νp��=8��M���5�:D�la�U�U
lIh j	� �F���8D�*��˰BѮ8wŜFR,a)d7D����k�$ ������.�愈�/D�|�RE�&�2([���
$�CD/D�<��薁!2B�h��ˣS�4�tC,D��"D��<�9t)ɢ2!����?D��D��n��e�e@Ɇ�.m��(D��
��0	�1�W!ǙN��\�T $D���#MC�?-(x�b�R�'q8E�5	$D�X(�f�	�����Q�6&}b�&-D���fd��G�AA%��9�!K�+%D��&��&�����I�dWp�`$D��$[;s,�TH��P�d�� D����S�["�q�&�Q�5c D���T����;�h*B�X퀑,=D��;`ák5Lp� v���R�(D��c2�}���jŹT�@!�H&D��Z6aS�-9l��+H�0D�*��#D���P�� !�E��҅U<F�c� D��1�h	60��I�CI�'�
��f�<D����˓l�Nx17'M0�P�d6D��#�.�4n.R%�@�I��'D��h�胟g�\{�c��7�(���"D����&�� ,T4Kg�x�*���&D��C��
W�>X��眅2b`��1D�ذ��G����y��Z�S!�8s�O/D��)�j�.K;�A�q��V��@S�0D�#�]W�>��A�ۂ�\a�TJ9D�� 89�&�_�#��pJ&,�/sC|t"OB�W��8M�������LX�"O6dk���:.t�hg��F��bW"O��IO���1��]&HۀC�"O��9ŀ��g ���Y�)�n5��"O�وA/39o�@�����y5"O��(�*_#� j�HC��P��"O\8� ��U�$51nL�}�H "Oz!�!O��88T�އ��� "O�x�r$%+o��R��@���D"O�P�_??`�X��'uJ���"OօR���J�[��ɧ_�d�"O�PB����s���P��:Cj���""O�	ɖ	ԥMlX��A0/n���F"O4uZcg�8��0_NX�Q"OA���@�\�b�E��F$��"OlA����Lb %04+�k��0�"Oظ�6΍�*2e񧊜�6,�b�"O�Q@�A�6�AQpK��`�)�"Ofm�@�E[Q"�,�YL�ٲ�"O��3儂�?A��`3i۲\P8�B"O2% 1\�`��ai����z1��"O�h��;���(���P^�S�"Oh��0��-c�Y@�d��mZ���"O*��i�u��A��b�1?����"O~���H�&L"u3w��5%Ȩ�:"Ofa��^�,�����L� X[g"O�Y ���h|�#�L�#�p	�""O�%�t�����e���z\ �"ON�P5�եz�L�'J��մ� �"O�	��.��>���G�3f�HP"OЭ+ӆQ0.�n█�/N��{!"O�s���@X������x!���"Oޱx'�ۗZ�����S�(i"5��"O~L�    �D�h#�3����J�D�,��j��(�NI~"W��>˓]�&X9C�&���K�ܹ��3J&5�$�6�!����/pd93�T���Q��o��D���O�JP��+x�25�5\O�'pj���kX"����D��\;��U�;nDi��`��t� �FC"��deذ\�Z��=��O��"�	3�'B� �/C�1y��R4�ĲHB���I�4����7n4�Zu�ȩ=s��Γ}�d�H�O��S�gyr��T��(���Ű�2d�@��yr��rO�����Y�p�>�����GW���ʔS�#Ҵ a�G9o��Y�a������>	���?Q�7X��PP�*���)ƋW�<�ªI�8N��zc��,m�1�n�v�'R\9iD�S~���b}��c��ĸ9Q�C�	�-���h��ֻ���G+Q�2牊w�j��?E��!�
�	�B2zR@����yJg�K� �y����Ei ��	$�6��dʦ7.�[���|��Ւ��-zj�~r��?�(^X�8�!��ވ�p	s�<��
����MI��P���(3D�k�'��(��I�/K��`�儜t��8�2j�*~�!��f�(�PR�?A��i+�	�2P�	51�#<E�LVg�.)-�<jmr�0�&���y��B2"C�ыK	b5�Q�aC2��'4� ��I"4�X�����+�������B�IA,��bj[����E��VRp�"O�m���O$�n1��H�YJ8�A6�'IQ�0�jQ�rN�kVO�",RԁF.!D�[D��W���Q�<�ĝ��?D��"�#н$�ґ���{3��Ɇ=D��z@H�r֊�t&��,�c'�!D��ӮQ\�Vn�U�2(�<D� R2��hq��!�]Fw�/9D��!���OM�q�"Yi	^�xV!4D��p�V�S¬e��J�Srĉ@�6D�dh�AD�0|v8vlߜv͔�Z�G6D�� 4�!��.c�4́�c��uЭr�"O�Hp��3Q��8���Y�� �"O�P�'/AD�I{GϴV�����"OD(qr� '�luCë(��h�"Op�K�7MXP�آ$[�n{p@H�"OP�a�@ٷ!1�e0p�/u��KQ"O\����%���R2 S!Jđ�R"O�T���Ҟm��$OXO%�ԩ�"O�P�D&��Fct���I�,<��b"O� ���0_jE�A�`��`�"O��J���;5�Dճ��B X�2(:�"O*�p�
7=KT�QIC"�谋�"O��q&�;T9X��t��6L�8�I�"O~ف� �)}�E�דe����'"Ox��[�"�v�����$c�lv"Op,Z৉�cP(aHg̖�DH�v"O��G��N^��j��J�|�h
�'���SD�]h���(� c�bb�'6�5�wS�(��E��@�.;�4�'w�كen��0��7 �$�6T�'�aW闶\or�i������lJ�'�^�Y�/��Uj�i���zΩZ�'y�b���0�Pi`����X�''.Dh�Đ7gsh�R��|0����'Tx!��ϫh/V�Z���p��ؠ�'Ξ��Wi���|d�TE�*k��E��'����*�-�ԑ;dC�f���'zңL	�z=�3�gU6���'����ł
0�K@�ۋYVH9��'�T�$Q�d�.���+TrL} �'��$Z��7#n�����1ɕ��,D����ǀ�Db4����6���J�A6D�����X�s���:��A:��@W#D�8[�b6YD�)�Q#mz}�>D�0�,ʩD��X#% {f	8cF#D�D���
j��Ѫ�O�9B�Z=��M?D�(J�HB�5��`P��1�����?D�d�d���Y�L�&/L��!�e:D���W�>%F�ɔB��h�
5 S*O�<0ckގJ�"�'�ҡ����"O
���LӋN���Bl;.c���"O�I�gD=�h�1q�5\ДQ�"O�� 2�ɂ~��-z��N)@�4�Ȅ"O�	�� зi�嚢cֲBa$��"O�P�'O4m�(��B�Vj`\�d"O4xK��9��2�פn� �"O�dȂ˟ (Z0�@��9_�0��"O�x����>%��zA�cOZ8 �"O��P���I�-ji#X ��z�"O���CЧP]��IfI��u�#"O��җ��
0*��$�K�b�ж"O6�8����8V�}�t�8;�T�#�"Oݳ�fz	$��`�ȫ� ��"O�-r�UӼ��5�͔����w"O���]�8�(�HD%/����"O0��&��
IQ�����-R���"Oj%ST�J�]��܁�1h�m�B�+D�dC��O�Oz�a��E�5�,����4D��1��_�KV!)�� 2�`�	5D�x����_kD)(E�P����y�g0D����FZ�N�� N�5B����o-D��Z3#B�\�a�J�$��Q
��*D��	E��I}P��D�.�}�$(D�� iT�Ov� ��`�`͡�B"D�� $���(�� �@�H�#��v�n,�"O�����2J1z5��C2aq����"O��
4d]�B#.p�ƆG`�A��"O*���W�$�n�RS��ac�\�w"O�$x#��&,�6� G&2o��� "O��
pf֝�� {F�]]�=��"OZ\AR��pi��k�f]�J��)�"O��Z"�B� =����r��D��"O�%��
%qK�X@�)l��#�"O�<��Ȝ�?�>�CE�̈́eb�f"O�}�&����1*D5�TH1"O�)񅀊
�.�����7V%�yR�
�a�)�I��A�5�ݳ�y��^,�F�zᇉ5Q��`U�y"d�6��Y�Gn��E�EF���ybLF�>���C�� ):m�q�P��y2×�o���iǟ&�0  �����y���� �H!�񢀁H9�y�nD!V�ʉ{��
Ji����a�y��Y;xa���%KR3��:�%0�yR,�M�:u���>���D�]�y��Mh$P+aL1�.hB�ŗ�ybg�6�������G��5����y2�4?�t��d�`Q�u��#�yB�S��4M{� ��P0���u���y�&�YáX
aN��E@�8�y��	']��IVmDZ��y��#��yB�C�bY���0!�SӤ�p4�ۭ�y��{$���@�ީT��a��U��y� GE�=IUL��f��򠝊�yr�I�J�Ƶ��P��qn��y"/��_D6%���1ޑ���Z�y���&��=91@F�J�JL���G*�y��1��z�@�J+�x`��8�ym��oP8��TK�8~��7j�9�ybjWGj��!���ޤ!w*��yR�$��9�B�$͘�'�0�y2��ny �2 ��f0*hs�B�yrEI�P�J|��QH���b&�҈�y��7pD�(.�/{��I"��Y	�y�'	�&������#j;�A��A��y�Ppt�Іu�B8��R��y�spd��#�4+���y��_�9����JY�-���H��y�N7���p���(�
\�����y��R�<�ٶ 2wx��W����yb�ϵ4�V�)$���n���	B0�y�f^�[��	�a�!Y����F*^��y���;���DC�]L��f
N��yb��*����H�n�f�
d;�y,�=�8@G�2X|Q�qb�*�y2�PrR��Ro��Q$p�z�BI��y��?;��xQ�습H�Zl�@FЬ�y��[f�"W���Ch��I e��y2͊?	�]� K%cXs7��:�y��L7��p���#r5�!�ƤT��y2�C�'*.9��'a\^Y�-ݵ�y�(/=��R+F$X�>����(�y�B�(�`X���]���a@�%�y��!�wfO��U��ML$�yFT�I���傂i9��k��Δ�yCߔ�RQ*��ڐq~����	S"�y�ğ�	z������')��d���y��7��AKl�#TL�"�˱�y
� ���SD[�Vu�U��$ $F����"OXص�Ҋhl����CZ��}+�"O}Yr��0j瞄HJ;"��Z�"Ork�@T�&`�Gn��"� �#�"O��4
%*ǒ��PO>H�"O����䍍
qXU����R���S"Oh�L��qC��`!�^�u��0i�"O�lc&8S�� �C�7dgޤ�p"O(��L�D(�F�M�Un<]z"O�`Ju�<q���P��8Jp$;e"O�\�G�/{U4�!Ђ�?3:�I�"O
�xR�P)��S��ަxw�	f"Ox!!¤+^��9�C!����a�"Ovh�uEY#�p�f�<t���R"O4,���/���3@�~w��Y3"O�jG�ֆn�@H��S<Bih�&"O>���
[<��� \��;�"O�<�f�Z�A2\9�GCRb,{�"O`�quG�	 0��L��8H��Pe"O�;��S\"$ҵ"��#�(�"O��.�̴20��$(J��!��,o�!�D �0
�3��R
�I��lʩK�!�d^�?�T��`O�l�������B�!��у.m0!RU@<f\"5ёJ(!�D��.���)��3	>Jx�GHE� !�
SŔ�I4�5Q)hh� a�wy!�d.uV"8����(<�>0(%M�D�!��d"� �&Ü���<0Ӈ �!�đV7x!iT��nτ���.Sg!�d�de�Hv�E�T�)�!���yt!�X��<ヅ��{��9���έW�!�ğ��n�S5&�v�ġ5�SNd!���
b�[afX�|x��BD�}p!�DK<P봍�A�A)i��10F�7�!��I?�,mp��>_��1��E�
u!�?e��\Hp��+?�,��m�!�$���d
���72y�O��!�d�FZ�ɻ�E�5�^��!W:?u!�[8F�� 	��&xє�y�@_�+Y!��O2���3ҡ�/�J�['��v�!�d�5s�dP���fÊ���H��l�!�d\+=#��w��*w��-���O�I�!�X� ��Չ�*�R�xS�gO�g�!�d^1Y�8�����X�%���)�!�$�!5"A�e-��!���7I�!�$܅�X�Ꝍߢ9� 
C�'0!���=@ �ی~�Rl�C	�� 5!�M!"*���WmY8��̠UC J&!�'_���D/�;@; ��,?9!��I����'W<^��X��܈b�!�d�	)|��B�F:|x��W�O�$�!�V�nZ�`󒎂���z�aڑ�!���&tD1���� �p�j/��{�!�B�ۤp��!��Ըsn��T�!���g)���_�1��Q�N�R�!��ӧ�,p��j[0<�>< ��lG!�d�.s(T����@=��b�lN|X!�M�\K��C�J��V��v��4!�Ā�e��f҇1m��#�eܭR+!��&_0�)2�Z8BP��j���3{!��"O
��Sj]R��4/Ǫ8�!���<Fg��0O��a@��*�nIwk!�Ǒ'��P�ԍ
sO�EÑ&�4W!�Ė	�̥�ƌ_�7vQ�r�ֲtE!�� �pZ����, �iX��6�^���"O����(�r���ˊ�w�e��"OI0%��#:�{G�Ɔl�<=�a"OX�S��)�`a"5e�P���b"O�Ԣ��~*lPPdDO�y]@�"O���&!O����G�� N�@xe"OWL\$"����9/�-���T�<� $^�
%>�HSD2`��#7�AS�<�+�('Q��ިN~�e�C�^q�<��'��A��<kRfI�n������f�<)���d��|��K������a�<�7n	Xxi۔A=0�z5]�<���4h"<���" �f-pЍT�<�BH `g�(�"i)2M� ��R�<!��W�r5��F>j��SŌr�<�OÃ2@�a����h�<���I�h�<y�e�%lJ(8���G� ��l@U��k�<��*َI�0Ի��3Pm����a�<��\?Z.P�����OuVd`'�\�<q�M�\�(�sk�%� ����NX�<��@M
�
AJ�,�"ad9���b�<���9`8P��Y#������P�<14�D/d�Ѐ�����ܵA���e�<��"·fF�E��B��x/DPI�LU�<�"+"���BLB���I��
J�<7�Q;9��U��	_4?� �0L�m�<��D���iŪ��%�be�"�i�<I"�%,z8A!D든/�^��%�}�<�a���0�$ k�䗋k�
`S�/z�<�Β�訒��Xi�.�R�<1�dI�����擐�zђ���H�<y�`ԎKh�Y���dx9�c�SK�<i�J�
#��Z�K��t�ƜK�d�4���L��N�)�dX�V��O�8���łBq�!W0G�K� �y2"A�U}P BF�Y��ㅃ�9�yb$X��)Q�M�s�6��%
�yRdՁ�萉�)�1j�@9kԬŧ�y��̥�$��DmB�\8R�3�P�y�"дI�4@37�Y�(Y����y�*2u�h�/צM�"�U�ԗ���n�&ڄ�I=��0�:�u�K4ꢘo�,Vy�1kF'��}��F�s���j��i�~������0@<( K� G-�`"�A�^(�U�!��F	z�BI�B���&���K���Y���Y��l����0�f8H@���5���)n:���A��t�9��ێ=�:��/��)�T�Qg�#
ز��3�#��|CA)��m��͠&��z����O�i�WLF�Y]z���`_��y�Ӭ0@}���m(���նOJ���y�t�Ơ�+�R�)��UZ~��C�$Oc�U�����"P]S�Ň�+<6M�$f���#1"�u�O;��ig$�= �0�yS� X�Bǜ|B-��Z��=�}B�n��2i��/O��Pi���<��4 -�1��)�]�$�Eܧ�yr�A?}�-�CHG0S0܃�RJ����hO>Uj���5Bf��b]�7D���p���IxyU�"~Z'���F�U!ԏ��*�^}jb���<a,O��=�|�P���6Ɋ5��2k�� a�U~�)§P���`oT��M��h�0�͓�hO?���G�T��-�fW�P�{�@q��0|Z��)?r�M�D��h|�y;��q�'&�yrᅡq�dP�$#->��K�����'���hB��$.��!�A�9"Z��RaF�(N}(�Έa�<�%��t)��Y��`�r��J\�<FJ�2��Y�DХL��0rAA~�<!��N� 0�(�̥�0���e�}�<yE&c�4Rf�$^z���ǖB�<AC"I%{�H��
��	TrP�@N@�<����������5+ၛ|�<� V�Y�A�+ھ`�F�p�9;F"O�ң��=�z	�&ʟ2�t;F"Ot����D8$��{�)��8X$�2"OR�
��|��`Q�
[Q"(��"O�؋RM����)�(�)G��`6"O<��Ѯ�\�hpr!EH��!"O�X��o(+���FH�XD̡��"Ol�"&��D�!��Þ��qP"O����"�	uVx���j� h	"O� 31�?/�00p� 3q��=��"OKƥ�5�1���� �f�;$"O��8!HE�pZ����|���j�,3D�l�V�J�}a���6HF� ��yA��1D��
�L
4�@��f�	)�P��d"D��*�I�h�8����ߟ��X2ӈ=D�`@q%G�S���(�n6U���h�<D���AB�5��ݡ&h�qv��5D��[�a�j!���B�8����cd6D��
�7}�Y�qM�I�,�#p@5D�qi�|Ю�4tF��1-RC�	�5,~ɲ�"�|����oC�F!JB�Ɂ[ʬT�箕���);��$�B䉄S.��V��0�\���I�qaB�I#1*(��t I����ꌒZ	�C�4)��MԄ�mB��჌���C��C'^��� D�-���WU6��C�ɞT�`�HS�'-����$�,�C�	4چ��S�7�T)k�`>D��B�	9~�����siA�	T�B�ɀ6.u"��$"����b�9��C�	g6����%��h�!5��C�	�F �h�v&ƚo6ց�@�::tC�ɑy��h9Gjϐ,R�=pğ�FC�	�+���Ï�ra��E�K�[ddB�	�~�
ݛ�hR�A�IsF��5#�NB����Hg��� �l�����\C�I*5p2��2�y~8�����X��B�	�)	�Н6\
�b�^N?�C��Վd��,$�	� hO
`:C��j?�xCW(��P6� {��K(L�B�+�()�t�D�*�����\��<C䉍��9�B�f���0
@�C�I�RK�cpB�-O���CH:��C�IG��,"��Q�FR28��&����C�)��x�g�y�L��NA\)�C�I�[���WB��"UɕHL�ޜC䉿��4�!%^�5 ��N��V�B�ɪ5����	�W��{ӥ�35��C�	��T��M��?$y���� ̘C䉄R`l�K6ğ�X��x ��-�bC�IW��	z��]�SC��0	A{PC�{��Bw�]�,&d1(�&�\�JC�8'�l��v�ȩ"�,]K"B�'[�.C��Z�|���ǝ�a�&Es �^�C�ɂ���Hi\T;$�(Q�L=1�B�ɡ`s�	أG�@�(�/U=Pp�C�w��R����4�@j}�C�	�q}t�p��rX(K�ԄB�ɇY 6�(�� M[���VƜ�:�C�I�9��(���u8�x�^�j՜C�	en��Wǌ4�ja�Fj�Uv�B�3z�@5�p�F�`��a�6�}&�C䉩L�IC�z�E�M	�C�I�� q2�H�l��oS�a?�C�)� F��b�Ѱ|Htp��,Y8#�ȷ"O�	ƦF(.�@]A���7�]�"OnI���F�^�J�j�踱�"OZxxc��8��ذ	ވU�0���"OⅈEFՙk��H�Ɣ�r�4��"O  �H�D�>=��kȄo���"Oإ��Y�rd�a�ɒ&	���)�"O*,���Q�upb��WB��(�"O�Xd�"\8���@�j�� �"O8ik�	�, ���ϋ�Zzh��"O�XW.P:'rd�����Tu�j�"Oȑ�J��p�8�Wm�69_6�14"O��QgM�2vxxc�U�5b����"O$��ও+LN�h�g�L����"O�U��m�##�QpGR!]h@̺�"O�*�/�8/�t�e���%���y"O�|���?�L�R�P)G���P"O������7ip�P��� �8�(""O�$N�f���N~��,��"O �3�AX�-�����CX�F��PK�"OB�Yc�ܵ"�Z�kʞh�r9Q�"O������'�~Q�"����0�"O��4�ޓ��[�Ǜ��9"Ol0��n_�U��*Ư۴	=��q"O.HpU���s�����ǌl5�<hW"O�qq�΅?��P�%d�&
(5��"O$i�G�;D�t����D�bAC"O$��a�%��A�o]{��Ѱ"O�M"��?nf���.�=�Z���"O��Bs�W���u;��0T�@œ%"Op%)��Y�!�Hx�@�=�h���"O`�Ƌ�(�>A���2!I �3r"OH����H5��8 9�a1�"O�ܫ#�F�f�,2GڇM'��B2"O�	;D��(־؅�4v<\�{�"Od����=r7����Z�W����7"O�!ڰI*9���I��I�f"Of���-Ɓ@�潲�a�/���+"OZTxO3�<��4]!�M�'"O�X��\��l���*& �m�"O�8:��Ǳ*R�D�vA	O�Uz�"O��QG�-G
�c�϶Z�"O�T��GU'\^	��-I�`���"O����G�DK�i�L2��Ҁ"O,� ���@DZf��!	&"O�q���#[Z���d�}����"O�lA H�%mp8X;W�J�z�:�"O�\�U��`��(� �5u%��"OP�S�P5D�dY;�`��&��"O��z�mDa4@���,�u\���"O�PxB�KI�T9���VUbʁ��"O�Yj�$N��1��P���ݡ"O�M�ei�(B*��¿*�����"OX�a���#{]�
��N���A�"O΀Yᩜ�((P!�Y�rm���"O.�ඪ��sӪ�ᅋ�)VV�Q�F"OT�Q5ꗫe\��d_�;c��	r"On�wER��Ub�D*黀*OF±K$A5'6����'
�+BF����Y�l�A�]��'��<H��O!l������ I14��'��,�&��,�h¥�Z�IN�Y�'}`9B�[|� b�L$v�� �'�P�÷�Y$�8	��F�`C�"O� ���3$Ը�A���ױam\I��"OƸa��*�(%b���>P�P�"O����%f���P  Cv���"OB5���"1��u���H<E��C�"O4b3$�(/p����0AE��S"O�)&9�"���f�:Q��ySr"O�5�Ua�4&Z����R��<rS"OF$)���3qcX���_Ot��A6"OH%�qgS�L����	O�RZ� �"O�e�e��L������GAX9[�"O�]Q���M�� �����@XT��"O�+S�E���Pz󥎧˔�s�"O`́r@<*p���1���C�Z�"ORD�jS�ȼ��sɎ8r��B�"O��Z2`�4o���L&��QQ"OMyR�/r(��&��S���2�"OzY���ܽ�V�	`gO�b&��V"ON����p?�T���1���"Oȓt��[��s�㑸A�*L��"O�D�Ū�	m����t�:�
"O,��aP�T�YT�۲c~�9;t"O6����kyJ�s$'L�id\�)�"O�m�g,
�aW�eDP�n����#"O�DH�ȗ�.�vlp�!ن-D`��R"O`� �����s!��^\�2u"OX���"x���c��-ژ1��'����n׺����ЈW�<��'���R��F�|<�ii���O�(��'_�8jP-ץK	�Mx�PT\:�'5���&�S�O�����\�F��A�'G,���nِ�d���	��?m���'�����
�8e�2��E��&=�: �
�'>-��D= �J���Z~��Y�'ㆥ�a�j��+�LыJ��X��'�Z�c�W-0I���$֔
^L�	�'�`�pƏR�`��Ă5��	�'[̕�Ҭ�7���� a�3-�f�	�'H��Q���?s�q 'H՞+UFu��'` �B�+�(a�G�S�07\�s�'�2�i����1�d��#N���'�R�P&T*=��3��h|�]�	�':�QXD�H#�u I�KGX��
�'X�cS���	�4��0��'�n����ܳ%�\00�_'U�����'UnٲDN�'7�tJ󣈍C ���'����E���f�P	��590h�a�'"253&CRKuh��2Υ$�1X
�'�2�zgG݅3�X|hr��f8f��'7�s��U3SI�i[,C�O&��
�'Ĝ9��ȃd����%����	�'���V��� �,ذl���'"ܹK"��FU�����|H����',v����>cϪ�Q�!0>y���'�00���P)\
V���-=l��'4����
?Ont ���	�P��'V���f!��G#�:�&� �'���j;5��P�V&�#20����'��UQs8 �np���]�� I��'���0@fG�7�*PSAF5U?����'�r���cI�:o A
��Q3R���'oR4�%�
�Rv����A�ɋ�'��h�dV9w�� �I�n( !�y��'Kx�:2�Ԧ�F�T���w�f� �ȜVI��� ���	џ@�#M��P�17�i���[A�UC�$(1���?�Js�Ӧh�:��L�>,����D4��,=I���-��z��Հ^(k�b|2cJ
Q���� d�jцP) �t!��.�0l���*��m���Kɦ=3J|b����$��"Cj�	D���yݬ��eo���?E��'���b>��xW��8+b�a�b��p=���iǠ6�>�F��>�NѻQ�U*Ԥ����L�,(Q�uӲ�D�<ͧ���}�&K=e��s���)��_�sj�pP�%1)^�1#�Un� = צ�
�S�?��8���Wf�`&��sD��<��p���Q8Oƍh5�%}���B��:7�����$����ͻRQ@����_�r6P�r�9e���*��'�7��dyB7���?���Q�b�	73���1�כSTP�@��{����� �J{�=X���6iD�%�Pܓ&�r��d���ɖO��t�i?X��/Za���UC�+%쐛�#�O�$b���x"���O����O���;�?q���M[����=�@���OT�H�l�eڀ$���
Q|)�7�'�&3A+��j[w��� 4@ ���$Ò-��m�*FH,�X�ƞ�uG�IP=N	P.K�n.�ɑ�(��b��tq�Ô0�?i��iD�7��O@˓�?�K<��-'�@�%ʂ�Z޼@qiM�'�ay����԰�I#Qd.}{�
��fDmZ[�Ow0���~yr��iq.ם����ȗ#���7
ғe�V�B��?���?)�% ��?���?��[+BXaL5�
1Ōz��r -]u������t�4=��Ey�/erdy:&K�*n~䲃�Y�_D�v�%~�H��Ǭ_� �@����XR̵Gy�\��?��i��r�mz��1*�#ܱ6n(�&�%��[�l��c��|��Om�W������6钺u�L`b"ONI!�jE�m��Uɀ��6J�`�ԬH�Vp��4����?$�fe���?�J~j�*i�d8,���2���v�h���3}r�'6j�إϘ�r�Xym��]���(#�K����g�O��|J���j}0҃�F��H�}B��MJʡ:"]�Ph�ت�慖I|���ܨ3��9��D��1vCƠMn���Z�5De�	��M�՚�$R?����	�7��0Hh�F.|	g�����?��S��]>�99X�s#� :G��m�GÄ���Є�I��M�S�i��G�1��1j#�G�)/>p��OU>o(��cI�7bn6��O����Of�	>^|�d�O��dtӘ�*�%2iG���֭�A�H#`D�0z�ĺu�#Z�JU8��O�Z cS�Lr�t�O����;m�c6Lղ&�`�Uo�:x��գ� v���*�˶[���t�S�]i�-����k�و�����d�Á�=*=��sS���?�'�i��6��O��F��O���d�/2$hy4Ù'r�l�iM[�8���1��������B��r!BP�'/�e�Hl�[��?����uSVK����	���N�I��T@1}��'`5�@ ��yX��,R~i���:}��'�n
@ ��� .K08ₛ�X�<��)	5^����M4|o0�yqDV�����fN�n�%J�T��MZG!��|:�<�G����Q޴b5���'�$qF��@PL�,����5,��a�D�O㟢}2���.lö����@�@�⥺��~8���?�MۡCW5:�����C�1����/5�UÏ��'x�'e�'�h@ ���:?Ȥ�B�/�;6�2�y�F�D���>1��яA�:��4m�' 4�"C�7M;����i�<	�nJ`4��hӞ��p�ǥS��kS�]�=m ��'���E�F��t�'UĦ�YT�	^��Ma��%<\��E�� �@��5(q�h�� �I+;[�$r2B�.0�����L�0�9�O;�X�Q�z����N�C�*�0�4 �qO
l6�'z�6��-;xF �"K֔��� �L�~�AO�x��� &���~�A�Ae>�����e�z��ŋaO!�Y���$�!�� 9���a ���ՠشg>���'*l6���e�jpl�x�	ߟ��ӱ-.:	"ȓ
�P(�"��_�n�c
�����Iݟ<��
[$���2!�!z֘ D�m��Z�̟����&���iD-S�C��:���N��1A�EN'RaH��$�ѩxHҐC�GTx��Э*��ɩa'�C�U�'�B�O���'_�6M�¦��I@��{y�2$
�y?B���G�X(�r���	CԀ����	����%.3��T�'U��x�hLm�k}���;xb��Qu
�(�~q��j�(��I���$��GzRhK5 4  ��ip�@�����@��N�6���'��Ո@-f�����n�pEA�
bZ�$ե
�n %i��Y��:�V�e1��D@��2���[� ����?9Ɇ![��8G�C�yxꡯR@�.�KA�vtx)P�E�-�ơ��2��i��) ��O,�3�DF'%�0�� D�b�`-C��ie��0��B�V�6�D�Od�D"��FLȈԨK�R&�Ա�황|��?��S�? �����=2�t�a�!"O�p-H�F	��M�������'�7�矒˧V� 隀�i=��%ә]c�*�f4X�yJ���a^@���O���B4 �n��OH�D�7��Cəa�-����8W�a�e�Ӵ@	��$YW���#"U�o���rw��>K䨐'D�n�J��P�ǕN_���B*0P��%��.B�LŘ��D��z���*g���$���1@�'Y�i�cށ7bֵj�E<`��\��Cy��'��O�O0N�����t[��S�$X����'�����"�Z��/<�Z�q��ʖ0:��l��M��'��'z�vEU�> T  ��:A��`AĦ�C�ʝHox<�e�;*t�`��p@���
8w\���@�	<-Ȥ���]�5Ш���T�e��!�F5z�]�\I�\;4Oԟt�v��"kS�D9�U�=��)��� ��4[�DqHF� �.[\�ӧ����`B+}B�'>B�|B���;$�� '#��a�F`B�� �8�������e*\�|��� @U��S��l�@-l�۟��ڴ;2!H�i���'z"�O;R�P�$P�Ό��e�97Nm���ԵsX��';b�\
n��3�\�-<��ƃ>Q�հ���DY��K�#�Z�s (�j�r��6�7S��O(-��/�?�L�*�̹;z��&�Z�l��U��'4~�;f�	H.�1�E�*�H�>AgF��Xb�4Kr�f�'E�O����1Q�F�rca@1-�l̋�/,�	��"|�'(�Q�՟e6���#dO1+Q�hǓ�?���i۔7M�>�w�0>`l�C&�!*azA���}�d�OO�"=g�?   �����O*�;�?q���?yq,:�4��"�	1�$�c^��ٴ�O"'��� GCW^2!���\�w�"�Gy2+� HV��+ДVn����'[~)��X3O��� �
� �b4H�%�pP�Fy"'ը�M�c�+���G'L�y�Z��&]ذ7m�����ay��'��O����'w\e!��ݔq�l���F�3�y�&�f6��h��U0�� @��~b�'b�7-�ϦQ�?A����5� �  ���KZ�i���:�'M¥d��Xm�x��?�Oĸ���  �A�%xִj�j�#)f��'�(���$O���o��-�SŅ@(^m��h�LԯM��@P!��0��Ο��'��3����BA��TT��aƈ҄y]�K��ɬ�M{��i}�ӌ�du�1eˆ��D0�M�glhـG̐�?���?I��t?�9���?����?) Gl�*獟$*�8̓��՜tG2�YҢ\1H�{T�g��Y}�)��e���T�O��u�hD���Sb�B"�I-~�d=�ǌ�l��qa�'V3{@H���sP��5����صQ8�'���J��Ώ5�b4؀����^AF�����I�p��1#ȉ���O�6M�7l��\K�
1, �hV�M��!�d�L��	���l���'K�vKVI�	.�M#a�ig�i>��S�?�'���R�1�H�q+Ng�ԙ��F(��x�$�V   ��M�/�e8�34��i���C�B�b�zy2�ܻGg%hW�73��$[%���{Bw�_B�t�ӯ�3Q\��RK|��SS�dʓ�����'��0 �
Q�Lz���Bm������J���/��gyb�'����!]�y[��o����9�y)ܪ
ÆP)5�L7�����< ����Wۦ��4��4����쟀O��5Ϝ�+	N�xCD�,`5��E �BH<���   �1'�J>'ޙlZ
^kB�X��N��,��#�ɛ{�lRB��9R�R�ڡ�_IyP����B��3���%*�=����{���"�퐪b�qOJ醾i��Њs)U�M�F�`w�&n��Z���a�J<����?yM>y��~P@��	�h�T}Sb+4p�d �D�>q��<t�@4T�j`B�!O�p��T�b�v��˦q�۴�?ͧBB��D�i_R�'��V����z�	d)ֶI��H����-�z�$

�@���OJ���/�`0A�-��I�$���Ϟ��}�e�@��<+�싑I�R�C>�,y剂K�����	py�k�#�'P ,	��M|�	�� �J�C�#��ZB��'�	z��কr޴�?�Yw�\�e�Ǉs��a�!�_%ri����'b���0r�(�'��\����(U������O��nZ�>bU�� 9��3A�-�$؁e&Vv���?�J>!K<a2�V" "  �f��`�ɽ33*�(�}s����9!x� � ˲K�\�ӍN*lq�0Za!�`X�§�	�|�����5���G/`��!yR�m��D:�ЍU�x��	Wy2�'�O�O��@��ܰ����� 8-�@���'^�&dG�&�&!�S�j�X8!r�Q7B�qo���M��2�'��'ě��ƴ[ T  �[��y�'P��p�7)еj�H��C�Ƌ�4�E}�OmӨ	n�����ٴ�?9_w
L�dOi^D8K���8�B��U��O8���O�� 0h��(���O��d�O~���wd��2�̼��Z�U�TH���H�g�����)O�A"7O���d�OgZ�#c+ߢ��dG�~t��,�a�*����2Z��0��A� E�^��+:��6��$�<Ұ�'�}�Ŝ�\��a�@	O5[EpE� i@覹�	2M(��	)���D�Ob7-B)j��i�U邩%�>)�&JH�r�!���(M��	Ԙ\�#�8R&���	��Mf�i�i>����?&�� X%�D�8g^�"1,H�2qf�'��nH<�"�   �á@,@�87G��X}b���W��n��	��Mc�i{����h�$L�𦧂�M%�6k��b��)�gyr��>ktR����A��5�M��p<9��˛FFp�\�D2��@E �%{�ᙥ�ŸN�M�O��D#��,�+�*�� @�?AW��̌q�e�-N��ٕCa���?E�,O�uY0iW(������!���'��em�LTl�m}B��<��k�޾nr�a�bA܆������%�<Ez򂍼 4  ��@ӥ�O�il��M����H��iT��=�@��G9�-���>�����*��?)�#���ه���+�T�0�G+�vy���O�ȠUnǑi�]J�"��`S�K�'�r�D�OB�ۦ��d��N�O����O����%�y7�R��"�$1���&㈓50 1���.'<�x!�.�:GL���O	��b�D��+O�Q����)��	�A���A�V1(��SNҘy�ڼ�P�-6�O��}`F�DXy��~���n)t��W�=��lm3���ן����,O&�mӪa&i��Uqf�J!-LVUvy�d�sX�t��(��@(��V�^��,R������ܴBƛ��|A��4S�T��JJ�^��2��Q�Tӓ��9���!�4��<���>0ʅP�d��j��1Ae���]���-z䠵j|�j|�uŎ�qq��񢄈��(O.���ۣU�r�R�̊<J�4j H�$�� EJ�)S��T�&9Eod$�1�i���{RH���M�W���U���D����p�!�)@�{ǐ7�@������a���$�-$�2Y8停�qe��KBÚ��I}X��F��+L~z1y��wRtX8"f� K:���'��6UԦ��i>����ɽ�M[���?ܴt����V�
,�J5;q�ˌy��I��'	�����'�2�'�T���V 
��5#NƗi�����D��ɑ(;:�>���hm��(yS*S�(O���ʗ"*�����m�l� ,����菗i��!瑳:��M���?� �Dyr.�=��iq�VqӤ��c��Jf'v�`C#�1"����&긟���F�S�O��$(���_$d�K�Ϩ-�;��?9Խi��1�b =��\N�r�!�4nL��?������ē8�P  @�?d�3����!�h�<B##���	G���)��)���g�<�`L.Lv�gE�+������g�<��T�=� DH(?��b��RM�<QF�-$	�!a����z�Z#ȁE�<�5G
�gwfDᕧ۶t!��Mw�<	塎/Xp4P��S�!W1ow�<��
E�Pwm�!uQ��h�<���.�ҙ0U��b�����c�<�3 ��U@x:���)C0�5�Uw�<a�nB&~�p��H�	��p:a�Dy�<�ׅ�Q�(`�C�6#*PR7l�<�,�iz:���K�u���0t�OA�<��7gh)����^]�E��Oc�<�,��{�5y�#��mbޘ��\�<���/���I�K
mݒ���C�<Q�oY�7� $Y���1:
���c A�<����J����.E��P�{�<a�o��%z.H�YN��3m�v�<QFJT+�*�!A�>Z��f��t�<����9,��JCHѳW�Yw�<Y��Z����ڰ揆a�:h�P��v�<����Jg�� �G�Z0���Iu�<I�)O��8�'��~ 9�`�L�<�7�E!ih��ᵪ/E�����EE�<YanV��������S��l�v��<YSÀ8��EX�]|�Y��{�<	5K�>"p�Z�:f2��g�^v�<����E&� �jί�
8p��IM�<)����0��|1�Í*�U!��o�<���. |p@�V��u8B�Yb�<���	)\M(E��IR=1ilM��Xt�<��� o�\�BV<K���k���v�<q3
ǣ�<9Q�5?��s!�K�<�u�۵D����G|M*ɺ�$�E�<Ѧ�O�iW��(��X�H�Q��F�<��	.*��iG(&بE���XA�<��� �  @�?�s�o��p
�a>�J�!��O&8>}�v�	&Aax����`A��@��v[\$r4���HO�<X!�\�*`@@���)' R�l�@�,0����>䘲�Dr@���;n�BቁS}B�He���4�.3/����UԺ@�aOO3�N,k�BZ PzL�h%�K��O�l *�(�@��<z�3u�L�"O��҂�k�4�z��Mޘ1a�K�(+d���S�V����͙�w�q��'N�E�o� ��E
4$��X��+�'Ҡ�:�8Sq�a�ïMm�)�ݴ[��1;'�4Nx����	�L����ύ+SV�P ��1j�����L��mN�Xp�Z�)��� (�(}�(�1vj.D�L�A�РR"�l�HF�uc8�@�K D��!$O��J��1Ǜ�~mD[�h D���#�^�A1����fL�D�?D�$2��/45d���)���Ɇ$<D��C���U�ͻ�a˦{�D�#�<D�����(&�V=H��K<H�+�:D�L!J��,
���P�p�P�7D���7��#e�j�PL�/&�@�@'D��dk�;^�,�KC/ډ|��9��$D���AbI�(=~���75S����a>D����F�2�&}K���Eb�Z�h9D�|�����-XA���=��d�u$7D�,#v��']�8�r�@�: ��0Y��8D�83��Z�2�|�%��X���u!4D�)�*ʱ	�%�0E��  ���3D�x[�MW�U���)})�չ6..D��YE⎡��`�k1}����/D�� Fk�$rx�3�F�|ڡCN#D������J^�M��%��U��<D��smB&>�΀�`�Ҥؚ��fd<D�� �b�,�h��*Q,?��2�"O���iѫ�֔�j��*�i7"OP8R@�$mV��eI��"�"Ox�Df�6f�`��g-SϒR"O�j�C۲f�R�+t��uˢ"O��0U"Ϭ{�2x��j��L����"OrZsCY�@?D�pQ�Ɓit�)��"OH�s��ݔ+)T��K�Kmȕ"O������h����)UT@��"O d�X>'g��I��)@��`"O�\ʕ`��Yy���rn�jj�m(�"O�ъ�l� ���#G Ge.53�"OT�DļR���mâQ�!�r"O"���GK"�\���
J���"O�p!DI��j��v��p��Q�"O&��"IJ(���ʓ��_�  ��"O��W��*D*b����,b�J���"Ob�؃'�^AH ���
NV$��0"O����NVB��0Q2fEpQ��"O�m�#`3�����$��!�"O�d��AX2�院E����"O2�3s.�)V.5�1�޵$z(xt"ON�ģ^�U�J��u��-V��"O ��E��O��ȱ�(b��s"O����ȭ9���G�B�F�H���"O�16.;5}r�fY���s"O���ZJDk��:yvf��w�D:�y2�,:��1��җlzL	B�ݗ�y"��#&l���'k��W�x�%dU�yr����)�!�O��إ*��yB(ɱ]��L���1ld�Z%�[=�y��@5*:����FHZͻ�CU��y��	&���jR��)�~e��_#�y2R�Dݨm�3�A�H�g�r�<!��/�x'A|U��E��M�<�PKK%W�T��
\>eF�� �A_E�<��,
�p�������C60�� ,�B�<���ɩ�9�*�Ji��;F�g�<�n%�^LJ̽ZGh���i�a�<Q���P8����8rj����f�<�1��#;��<�7I�jf��Ѝ�`�<q �$?W"]qGI�HR諠��^�<iƌ�d)4�q��A�&���[��C�<�׫���|�[��ԡ!�ɹ��f�<!���F� �1-��R���
GE�<��E�}$m��A���Y�"�N�< ��P$�S�Zv|>!�0�HF�<yWgN�@QN�8�V�+=����ZI�<����c����@�"�4�p%H�h�<If�V!WٞTZ1h�v���@4�g�<Y���"H8��!cٛ�j q��e�<��>}v<J�MG��A��\�<�P��ys�E�4���`��X�<��ǹbS�} 2��/�aC�XW�<�ʋ�I�Lu*P��R��(f�J�<q�e��9�@��ϟZM0,��cO�<��W�J���`�jb���ԇDm�<)T$N'
�y�!,V	�D�%�i�<1�/�"h��D��
éZ7|q���S_�<��ˇ�+���L],뒈�W�KX�<�D��!<��y5�˰�:��f��Y�<�!
Q�L�F����-�:�S��c�<�f�>	F�`� F�`z��s@�Gu�<�蝒M��a%#x�� 3 ��J�<� d��#&�j�X�1	R�3��p"O���jO�!K�P�r�J�n��j�"OV��DM�?)�.M����1:���a"O R�}��`���f���"Orݲ�Y�r�e�'#F)&���1u"O���3�2�yU�
M��+"O�	��F:KA��&c�4:�Թ�S"O��V��*���v�3h<����"O|-�f ۮG&-�����!1�"O�m� �ݝHc̍��,�@��P��"O2���/3*ܾ ����>� q"O����.,֩��a_8*w$E�B"O6I�Ζ
�D���@Ȩv��d"O�0 �O�(w<CШH�PPS"O�H�!���K�.�b���<WK\e�u"OQ�M�(R����F�Ք%K ���"O^젓 Q���$.77&��#"O�����!3�T|��Ɓ&8D�J�"OE�� �{cVܩw��/�izd"OА�BC*s/�4�&aM�#��q�T�I��^l@u΅F�&�Ad�Լ.���Ɂ ߒ���X�J,"�*w ���$|q9��R����=?E��K��8מ)���ѡz��F'L[�V��c�����������|:ec�y��Q�����,S7T\9��_�U!���?ib�O!��R��D˕�˘ő��F�}�ޥ�
L����b�C�)4�	5�ӱD���6'�P��NV�W�Z�A�JE/кYM\�cM|���)��Be녧�;��t�a+����v}��S�[��)�<�&�Z�9[hI���"OD��J5��Eê��ɤ �)�,O�Sm�O?��t�ҽ
"���jH=NUx�#�H�,٣(O"�0E�-I~���
|��Y��E�y��b�G[�n��t��]E�Z�� 
�6{�1�FNW�$�	IL�,�<a�J�IrN,y�'	�N���S6A���4Ǆ7{�I��}����;h �$���T�i�CB~RiB��8�{���Wc'j����?����)Һ�~BK%y�xl�}�)�L<�A�]X�90��W�q�F�
�E�!ّ��C�S�t�i�ē�. �w)E�+�6A�W	Y�L�9���z�P��2L|��d�!�~�����x|�q�焘/L� P�L5��Q}r�G ���	Ěl�rCM�P���0�j�'yT�a{&������4�M���٬kF��D��'���
B h"]!�"��Ř�'!�6�"*��O�]>�'o* jE���6�晸�c��2E�49�B V5j�c3I�	���Oszx(a�|����[��rd�B/9<>��X�NO.�F�tџ2m	w������Y����u��'����e�OM� ���Fk��x ��D��`M>0�Y:D��h����Oʨ1���1>�"L�MW�(�%h �l����)��������YsO��M�g�I�::Y)�J�A���R�[E��B�I'|�Rm�WIG�@T�a�ق��B䉪�Z�Y�'�2 �X����~B䉞Fe�¢U>�JU� �1O�zB�I�%�(� �7,�0Y��� #�vB�I�&bR
����2��!{vbB��3+#
���c�;%����F�D#T4B��hn����Y& as�EbtHC��&T��)2�m�:�@(��mGdB�	�~ ����lʄ1��.Jo�2B�ɽ9�>�c�,�%S�XQ��O�l\C�	3J��m�A �
q�VA���T8C�4p�tQkr�5c�t��.�a�C�I4Vjh	#hܪƞ0�d�9p��B�I;YꙢ�`���H��E�\�B�	�?��Jp/I�[f�tE�G	X��B�	(n]&�8�IG&W�t	�dY	KlB�	�Z/ޝC�
�'��0�֬\n@B��+H]��)T�"�M���R.�B�I>H���#�˓:��' Q6��C�	�Ymd����93���"e�(;�tB�I�"0i���.5�KZ�i�P(T"O� �@��l	MÖ9�L�5Dr���"O�!ص��<�,BFƝ�]���p"O^<!��64^ ajWO�b�1R0"O�l�&S b�.�1�&�Bq"O����2���2t$�3v�L��v"OL���$At8i *
'h�Lu��"Ol���펩�k��,b%"Oڱ�����9Gj�X�ZP��"O�`2�ޑ%ŤTG�%r���"O��1m�$3��3f((^�U�%"O��a�.L�C@�I�D!�����"O�e`���&d�j @7��}��"Ox�{�+?gt�S�E�;tC"O�)X�e�5nZ<��C���E��"OP#�B��)���`%��#4�r�"O�p0�0�
���@�6$��r"O��S��)m��Iס��s���F"OF�ɣf��E��i��M��H<D�hic/�;^�
��"��`��D�#<D�t A��7a����-t�j� ;D�@�2��	O�$<:�KS"L���o&D�T(TɎ1.�N�Z���,@�F�P!�6D��kp��)���H`HG��FA�vd/D�DЗ�\>2Ш�W/��Ny}IWn-D��Y��'OL��ӔMؒd�yC��7D�\�Bŋ�\Hr���R�C��<��3D�x��0�(Vi݂[���z�+1D�t���%sdp
f$@95��,@��0D���@�w3:l�*˾N���j#D��'m��\ݐ���)V ����$D���%�⎁���	�U��=S���y�B1��lK`���62VAc�>�y�&Q�%�hit��E�ĵ�R�B�yra��)D���Qe\�5�*`#���y�H��E���S+.F|)����y"H̸t���d�Λ;�x��1�y��;k�-����+�Hx����y�>��|z�ԙ20�q�@(���y҅S<I�@T �i�0���z ����y"�5G�~��7Ň�u�0�W����y��@5d�tsf�H�q�L� ׄ���yBj�"��"�E
�p.(x)�d �yRE\>T�PH�Sƀ�~?�]�Bٝ�yrJ�%6���
�'�*.�Ψ��9�y � 5WH�,?*@i�f(���y���rz.�Ȃ��0P�����ܥ�y��x�0��g��]����hTjB�I�B�^��)G��ɉq#ֈO�,B��9\�Ω;��T�}����!H'+<4C�	!a� ,�D��%�)��nєcYC�ɖv&�:� ��� ��/� (ЮC�ɉA&5���;&Dt���(�!���p�r����;|n=�Al�&v�!�<��Ec�D��h��E��(�5:�!�䗌P�<�� �O��%[��22|!�$5 �<�aR�{�����N5D�!򄄹��Q���6m"�5�g!�D� JR]0� Βu6���l���!��;g�a%�� %�ź�H�@�!�$�r��x��
YY0��� H!��T; �,�!���WrD���ɠi;!�D�Y�jI(�웪6rj`����u!��P�B%�h�r�yt���h�u�!�@8\�ؕZd�C�c_���᠐��!�� d�*�d�`0���0�0uc!"OB�fjK�qU\��g��4u�f�"O��Q I�����5)�s�8P��"O�,(��/q�1B	B� �	3�"OrܪbB�V�Eb��oX��S�"OH�P��C�Nm��a]lJ���"O�P�Ί/X���e	�<��`b"O�1P��X�Y�B�c���~�e��"Oh��")�+�C#G�X�m�R"O2�xd��'p��Ъ��+�X��!"O� ��Ξ�|P� k5eGN�Xz�"Oꠠ�	[�b�dp����0E"OF��F]�9Ͱp"!��;XN�XÀ"O�jv%*+���I��d/�s�"O$����XɞA��Hw@�p�"O��w�҄N/|5X�&�jb�{W"O��R�Ղ/�h��G�+�h�A�"O"��cL?]���	D_�@��!K�"O����T�9��9s�]�.��5"O壑B�!'��0�UK�0n�@p�"O��3q��%?J~	듪H8\ʄh9�"OQ�0g�D�)�e
ٯP�2�b7"O a�g�S>
2���DXVu"O�y���2�����)MH�;�"O��V��
]���"tK.?΍Q"O �����VE�e�D7�X��"OMrtr�!�IE�:�9�w"OJ�t.6bF��VI�	%bPAP"O������dNj�s��J�>��p"ON)���I�th��� "/XD|�"OV����6"h�=���=9t�I�"O���$_�\�$R��-�yr�"Of�3�I6	gp%Z�� +f+*e��"O�i����9�(h{d�0$T٩�"OV��ɷ'<nh ��v��i0"Or%���Z7w
���)ؽX�"OX�{��F�Ne��1`�\(RN���"OZ ���3Sy�	�,�S<�4A�"O��R�9�6�B��E$�̨"O2PrD�_ި���h�*�0-�F"O^}�0$N�3`������ z����"O(-�ǃ�,v�~���?�V���"O�a���1鮼�B�޷rDq��"O��G�&0�^�0�o�&d��`%D���c�N�j�Z7IZ�����>D�8SN���~�P��\�4qT�1D��@�h�?1�n�&DN�"߀���j1D�T2B��/+t~�d��<��%.D���CD:�N�x�oI�0�3��(D�8��2̔��9��9�L*D��:���:6:
��3-�`\�q��=D�P�u�I�p�zX� ���C�c0D��y����FC�Λ3 ���'�-D�#W*�r)��Y�DO�2�X��+D� c�LD�n�T (�`BK/�lp�")D�@��cD���j$�2N��XR�e3D��q�V5>��if�W⌘�ס1D� ���ڴ?�`a�7	��j.EhC�1D�tP$�Mqx�I�ކA4�X.D���gh���\ F�Z`�Q� .D��"�]~��$�m\�&�P�2E�)D���p#N�>��0�����T*L���i&D��0�_17��T����D�"YF`&D��(�B��&�|$qQL��M����j(D�� ���$�N�@$|��D��l{� H�"O|�����C'*�i�Л*H�"O�����j�x�1�Y�Z�I�"OT��T�A�M�e���P8u,�}�S"Oq" ���b�<�҂a����qV"Ob����� Z���$�܁vfHL�s"O�uA��WJʩ�P�ZK�`�"OP����^�f�Ց�7g��ɕ"O�a1gHD��,� ̚�`x�p!"O�u!226���M��y[h�V"O��S"._/n��Ȳ�)��c[��"O�EIG�'Tq0���#o �]K�"O�D3���	q��H�A�8sz����"Od��獌�zd~�ibō2y���"O@5Y�D�R9�1�ń2�����"OR����w�A��֞.gQ02"O���U�[/;:�ѐdפM�
s"Oi��bX�l̚-�S�A�=��	�"O
(g��,�j���RH��A��"O��+��B2{�v�)o�d�^�#�"O�,e�o<�NI�[�<�P"O����&ie2Ѳ��Z6���ʁ"O����K�k78����؟B��q"O�����P���\2���;L��d��"O6��U���j����k'���Q�"O����ӵe��� t���R����s"O��
�Ɏ�^��s�H�""O�`���[�"�pH����F�*�x@"O�����y�����EzFv��W"O(p�`��![�	-J/SI�Z&"Oh�:�%�~ x�!M�	(��"O0�4߲n�Ȅ��邹_
ts�"O&P
�$ֆL�x�rʛ��t`G"O�l0�а&���("� ����"O$HqG��*+�T���LG1H�d�F"OHʦ)���(5�E
ˀ�ɷ"OT��ua[<�̊�,әVz$S�"O�١�)��D<-���,=�9k"O��ee�&;Z ͓f,�*����"OYЀ�V�b�����
#'>��"O$]Ц�[�}�^e�R�Յ`�"�["O80ڇi�>m�&|�$W���(�"O��˴�[�1$*���cƶ:�0�"O��;a꟨$lM*� �T�L�u"O�"T�Ç�0-`�.-���[�"O��93��g��K���8e�`��"OB}H�m3��ap7g�v�m;S"OZu��� J"�([�W���K"O�x!   ��   m  �  v#  �-  �6  A  �L  iY  �d  Gp  �{  �  G�  ��  ��  Ϭ  ��  m�  ��  ��  ��  ��  ��  �  _�  ��  � �
  X � �# * �0 �6 = ]C �I �O &V �\ �c j �p ew �} � � Җ [� � :� g� �� �� �� ��  `� u�	����Zv�C�'ln\�0�Jz+��D�/u�2T����OĴ1ED�2�?Y����?�fY$E+���_(z����Ĕ1jbd�J&�M�?9�����[pZ�PgCG�
6�΂�G.��	_Q��i�tk<��Ya�M�E�A3w��I`#�-�:l�P),,^B�{�+͎<^Ȭ;ewL0�����戽d՚-����WFf�d�D�H��D�|'��D�>��|KW�7;"�oZ�FPr��	؟���������\/z�P�c��8G��sF�L�X0M��:�8t��4`���'��4�O��H��O)�wБ�%�9Ivxp��ǿj!X��R�'6��'�R�'�'����Yw�@�b u$j��q�C/�z4��
(~5*��B>:������y:"�<�@$C_+�'=b�p�[��k+Q��Dg���?y��R��Z$�y���7�pY��یy��8	�F��?�`�iQB�'�B�'�$�'���ּc%�Z�m�P@!QO�+Z����Q�O��(c�4Hy�du���mٟ4��4�Ę��is�x�C�U=s �!�/�7��!��R:�4��L�>i!+ӾRb,t���`ےd���*��|�X�'T������m��(�gf^Y��BՈ�.^��Y���N1~����ݴN����wӸ��
�|� ���M��
4g��h�L��S �� ��M#�FƟF�<�s�$�Z$ �x���Ӌ�;u�,6M��1��4^R6̢���>zZ��3`PH�;&�/�z��=��j�4R��j��3�����HN��D���e��Ae�U���ț�Xva"�\�U�9��O<=��w��m���M��D?G�D�s�X�A:ȳI�N��
�.�8)���T�nHܑ��i���s'h8Fj����#=���s�'��O
)��Fk������ڞ M�P�n��[c�Ё�H�O���O��I�jX�`ќS@P��n�O4�{��F,7,� FJ��l�����OL��?����d�CvHȱ���=T�8����с/�f]z0-N�
a		����h��͒Lԑ� ���]0}1�ձ�
H�ִ�%�$8�r���׶V���j��ȓEZ6�#@jY�]���F��ʎ.��v�D�']>]z��Pt���)-@ę���?������?Y��?������	�!� ��gPS�~A��AI>��?�G�i�*�HUcӶ�
��Y�ZhP�U�r�p�dF���Ş�M�����D����)�Ou���<K��]0R藶Ξ ��	�O���^��iC"j��J刔�N�{�:�	��t��bB��@����� �$	���	�8V��c� �xZ�As�(-��A�[w��x����\-�t�YiV�i@ve� �p��Ð<��D
LM��g��F�4:�8Aʧ偎U���f:F"�'M�O ����>g"����H4]�qr�BӒ�hO.��¦:ش�?a�i��T�r�>�9�A���+e�J.T!��'#�I�?�j��I����I���'�h��QȣG��1s�O��/�i��K�X�{�Q+�|��qh��-=�S�?�b�x����Jl@�	@"e(W��]�,U+�OɟP�(����xF��z��p�I�;�j<�9�T�
ve@�|,�	.�h!u�NA�'Mv)����rʟ�'W�8h%�ڭ'�ibv��^M�V�' �P�P��}�g�$��p��q�����3I�4-@uP�`;ܴ��&�|�O���V� �&�,s��5�P0v�RśJ_9!�ȪO��$�O����	~>�aR��3^H�#t�Z�m�]�Ҁѵw�����%��t7D����,a��B��������� ʂ�}�����DT�6M��gȲ#�"@�7l���LhF�y`,����Ǹ'6����V��Q�"N!:�����?��i�"=9�2�M)/����E4� qB#��	��'���'�dk�b�.8~���!FåOWEPL>)��i&6��<��N�;nx���(�ɜ?�� 1c�� t�@kÆ�Ɵ�	3(*T=�I������t���ř�]���Jش�y�ƅ�S�>=�&I,�|!	�+Q;�0<)��=t�`�f��1@�'2q�R����݇3���
$!����g�L�D��I�4�?�e
P�ɸ�JdhE2E5D鲶��-��$�Ol�d�O\���K:%V4+�bI�"Ͱ!��K���ht�Ƹz��S&b�Ψ�ŀX2��Zu����'�E�]�7M�Ox��|z���?YD%7��eDSCsʽq$���?���S�i��s+ ��D�	RPy���?=�Op�3�͘U�D�C�̀I��\B1���g�\�;��Q���+s��4�,Y�q�1`ӏ�qA���$��R��n����`��1J��H�I��Ms���d�	�I�ܕʷ K1f1���Ș1�'0��$ 扲u�0�妛�X�"H��A*v�`��$���$�Ȧ� �4�?)��i:BB�6���C�����jg�X�K/7��O�˓S�
`����?Y��?�-O�YB$�!x��Ţ��*��9p�Ȃ�vR ���o�ZV�A;ro���ʧ���$�DG��x���(L�e��a�� �O���J�54�D���ۗ!��P�4*I>���'^-`�o�༳2N

}��#%�Y T6\�3�؅�M� �>9`eC���|�	�����r��`�G�+kN�ꂞm�m��䟐��ܟ��It�g�d�A�������;���e�H�x��	��M�6�iB!|Ӻ�D��(�	�|�t�ɳ?��	���*+H�5����J���2��?����?)��>��O�d>�:P�B�j�\��i;�\�q�HZes�iإDiۼ �L�7�v�h��D	5'I҄�Bq	�I����Y/�`b���lO�<)�g��@��f$�S�'dc�Aɐ_�xzP"�~��p���ԡ�?I���hO2#<1����_6����M�7q���h�<�!$��JBU+-&I(!k�ȉ���'��6m�O�r(�Q��i���5:���NJ6.>p]�T��fyt���<���?ٞO������m7�QSv�YD��Q� (H�'��q�`���T-j�\��-�I�n�j�򤜴q� 4(��4S�� H�˃�I�ڹq%��h�<Q�D�.L�]E�g6�1�.Ύe���O�=���'D�6��nyR�Z G ��`n�+T��`���!����On�s��p��&>e�q�E#AU���?y��4�&�oa!��R�O�cf��Ћ��AW� �4��2rl0-nZӟ��'��ӟ���XД:� 
�	*C�ȟ��	�*��L RƔ9Bԙ���ҍ/9pK����E���B��=`Ҩ�s���\�58P�!��y\�5˗^�h�ʂ`B/D6�>n��D�?D�,XCĈ1��I9�FӉ���F�o�,m�^eG��:���p!�V�V��B���7(�����#�S��P�y��0�C�YUA \	wB	C�ў��	��MǽiF�'�i�0��%"�� ���3RT�t��'�'*`a�܊ �'���'�R6�r݈��U":*j���A""������>���o���x1V8d6�b>c�0P�>����s`�.ﰑ�墕�x	��4�?QfS�E��|�<����8(��3�*X9Yr��7�ȟ �'9����?���D^	�d��d�O��=#c�P\�C�	,�<�8�E�K`�Mr�L
6�˓h6���S�,�'�,A�J��*�2T�� b,
)r5C���6M�O���OD�S�'�nı�ɍG�űw#;(�h����	'֘��ڍA[�1 �����k�E�'Y1�ٌ�|����̻]KB9a_(���KM$�<K�bپ
u*A �G�?�<�S3�|�'Ԅ/b�YTČ���c��A87J��iG��&!ғ�O����)+��P��!I��.١d�'01O����9!V��`��A�}��H��|b~����<y�G �v�?��A�ј}�0T��ÿf%(�`��O:��?�����C��?�<����0R@�Q��K�}YN���B+��=ᖮ?
4h��#YDGyr��,.�0�ȕ�M%=S��e	,�>�[s��Z�M{���#rlK�(N��٫uɗ�^Z�'�����*Y��d�<��o�&� �A���W�\�[�f�A��c���a��jNpb�fݛI2�e��Oh�O��=ͧ˛���
�>�(wk�,_w�8:G��n�6�<i�N�m���'��]��'�� j2,�T���Q��ĒKsy���'��*PbnH��š��o9�k��n�l)X֧	���i�RB��gDRp�@� �!����!�$̇0(���@JL�q�f���H�q�ĩ����ׯU���1�R*\�Vp�B��S�*���M���ik>�ڰ�
�p"J�P�]�o�5�sa�O��=E�Te�-"\Q�� ���`��@ў�͓�M�"�i�1O��p�!8�<:���K��	2&�qӬ���<)�+7�����?y����Z:��(�dHG�J�x4��*6�L<BQ���j"� l�G��j.)��p���O���4(E?���s�5i�.�`��l����l�6��X;�*�Q>&Q�O�|�˔6|U���; ��T��$�Պ��ΐ&=�)ڴFT�	!t�v�D����g�I�X� ��*��0
��#)d�P�ȓw��-��[�b�8�#lM�gv|4��ɟxщ�4���d�<)�dE�*۾X2b
e��H㓮_��?邽i'��'bZ���O}Bk��$Fpp�(�4/�<�sQ��vw,@���� ��A��M�?�`��]���y���/�P��K&s�]ҕ�1�X "�o�I�r�2w �%M�(�/��"��1�wM��CuT�O�=�W�:BȠ�2�OSx:������"�
#<����'�f�@ŁD�U�Į��@�|����ԟp��{�ITy��dVލ"��_8�~e�V�޿���O��m�����'��p�VLlӾ��m��5I(2�^��g�53�F���C�O���?����4��,dm 2E�D(fN<a��d�����9�èSWy� ���E�E�q@�	4�Ey�e8����M��F�6e|h㵃�b�P�c'ؑum�3�e�nOJ�Y�`
d�O@�Y�'�b7m�uyb�ə=��Q���J{�a��%����0>!g�W��V����*0�0���JyRU�8E{�O"66m��-���ɕL�Up@���OCi0n�Sy��
�t
�6��O�˓���O��9�V���t����&�VE���O���΃ֆl`�Y�m AX�7-�8̈��m
0���fcPB�L�rf�ƶz�	�5�UQ��Y��Lya ۋ+�,�kS�S�R��PIe؟����k�n����HG�8y�6���6��O�}nZ�H���S;x<
T@�	�
@RPѻAa�!Rhv��d(� ���ԗb���:��Ӝ?��D�mӲ=o�h�'-�����.A>$�HH�"P;;{�D�Iٟ���蟠Y�oB�M����	ܟ��	ޟTϻp���d�]�r2���D$��J�R�:���xwܭ��b+�з*Ar�g�D�f�iŧDQ� v�J�f�qG�O�a��x�J�D�xbjBG�g̓q�j�3Ǐ�8/xl�{�ŷ\����Ir~�B��?���hO�iB��%y
���-ےc�r��(D�3�.%��+�C�� �����Ⱥ<!A�i>�	xy��.#�֨J���'q�hAA��1\���Ҁ��1���'�2�'���]���I�|rA�M1t����a�C�MA�	E���`��r�J$-ְ���b^��R�`�CŨ�<��
D~�? 4A��k�
��A�]�dMIq�S4W��a�Ć\�pЌp�Z$�����D^/`�P<ӳ"�t���2�^#�
�H��'sV7�Zq�'����� $	�#^/&ޭ���5D�����%��ہ-ĘB���!A`4��禙�I|y"a�c\:�'�?9�mB�PV�yg��d2�� яI��?���u�X�(���?I�O(h �؀UT���HD�l��� |^Q``H��	S�e9�.Û4�џaff�:*��H� I�;Or,:@/���ܲ�OG7{98AC�A(j�<D���?y�����M��M����:7�L��E��11�'�2�'��T�V�O�_���CWO*5h����yB�|Rt�'e��$>9Diz�ܪ)(�#����@�8Ȕ�lB�[��'���k��\�M�l�K�*8NE���'~2�'.D�b��X&&�k�b�2w��}BB�����ϙ̺�k�X_�4�pnI�^��O�T�@!��+R���W.A������	y-����#-�N�R�!2eFK��P5�b~"ʶ�?a�in"}��O^̼K��>����s`f�j*�r�)�#P|���S�83���!c�ߨ�hO*�� ��M+�4��|y6h�gF�:@���.ߛx��C��i"�'1BL�l�pٹD�'��'T�8��i� ���t��P�4�֙Sh}Bċ�.*�LJ�B�~/ !h�c[<T�1�ȓO�Q�:zR���bZ�I�m���T�3.6,R�"�^BΩ� %[P�F��J?R���N�2�5ZC`+k��@�1@Ź=��7?�2c@ß��	b�'����ȓ�� 	2���9�
��p"O"��K��5��I�� �"P`@��A�����'���>GD�I�*��s������#E����bM7/���������dA���D�OFMR�9 �Z���-:ȠY*c斎P���RO�|AiÀ�<
�Q1��$�C6"�[q��"FWl�m�B���as․? ��B�C�/ ��� ��G�U�Hb@����'u&1@���s���-}�V�r�HJ28�I��M²i�2\�D�Iڟh��|��CS�Fʹ�S��ũ7/��%���y"'�#&�H-3�@R�6{��R�aN���;�����i?��)��)\w�B�'z�x�DCD:���e�A(p�*��'Yb��[W�'	�I�
~�6䰔cM�y+C�IzI{2/�{�@��"%�2[.��-:��c�{��N�k븸��a$X�\����*z��2��̑ s8ia�M;��O6����?��OnM�`�T��0U�a�Y�5�У��|�'��k�(B����$2?TЉ�b(�Ox����CB`�!"N2!猼óF�f(��<��n�w�V�'g�U>Y�!fM���ȃ�ZP�a�c)L��  �� �	.��}Iu�@7<"~��@Tj>��O��ӹd���h���\�,�D���*�q�(�iÏ��".��[T�]�/��|�� �C�(�"V&B	�0��&�h~2̬�T�IM�O���0^�@���%���Vx��B�!�W�G���@چ
�f Q6��E�џPȍ��Z�IT�p�◻w���_>g��6��O��$�OJ�K�Lx�����O ���O\�]�U�px�F5|�4��e�4�mY��M���·�C	j7�M���2��ēu��蓑c��S%��썮z�k�ç)U�V�»<���dG�x�'�x�7!T�<.�fHcԁ�[5��{�A5��X1���I_�g��>�I��.�\E3q���~F"I��u_l�Ѱ��<��XhE��x�'�#=ͧ��
¤��B������S6qDv		EP���%���?����?��'�?i���?סݳza�8ZBI�!fF�ӀA�Wr]x��G�5���	�"]9H�g˫�V] R*��p��I����dz<zr��2�����+1O�]�����ҝ�u��t��2J
P2}�~-l�����'�r�d�M�x�nʦ~F���D�ӍT.�O���D̈<��QJҦH\PL�s#�,U��'�b6�Uަ��'�>�v�'�B�'����# n��)��|��R�' B�N�?�b�'���\M2�"�'8ǠL�'v)�%�POR]�N�	D�r$�A�����^,G�֤k�%�+;�ppK����oZr�k�m�i(ʄ��Ƣ>��%�H�	n~BJ�/~�"��%)B�~� $����0>�'�ٴ'��D��;q��3u�[��Db�1���z"�0|�0H%\�D..��hy���K�7��O0���|�4n���?Y�B��3bkP�*)�p�'�?��+�ؕ�ad��>a�4��*1����?=�O梅q��Mb�P��̗�VjD<��O�0 ŏ4g�H�JQ� ��8��j�F������@φn3���TJ��~
�B'��C%��O8��6�'�yro%`��xb'�O�@��	��yZ�6<C��^�L��1F&�Qu��E�6ڧ4X�R��/u�RDh�Aђi7��B�4�?A���?a0�Y�)jl���?���?y�w��a钉;�A�g�P;����GƐ
��DԹ�EX�ϨO�1A6H��mq��1'-�Xt� ���
S�`�E æ��a,�2c>c�� x��5� ?��Ƞq��eP4�1��D[�e.az�&J/�$�)f">y�:Pk��C��y�b֥d���b@^�mB�8���d�r�����'��ɢ�,���ㄮ{?���&��.]�yˀ/�ERT��������\w���'�i�%+I@�^X��E�Y�4��GT�jl ]�eH�
].J��[�H`ax"��v:&x�sÄ�(��m�����U����(t�����o���)
Óp$��W�%DQs�폮)�$����ܟt@�4��F��Gc��cxY�gF�e~�R#�C7C{R͇ȓl-*=��nU�a\��:�в=Ɲ'�a�O�����S���ɏ8ʸ�1E,��lu�@Q@Gþ[�ʘ��ٟ��MП����|�����;v��`C�j��+���O.p����+�d�	%⅟�.�`&�'�"��֍A�&I��)��
3.p� ��h���?R�1FIZ��0<	�HDџH�	}~¨ҋa:���A�R������6���0>Y��<%�b�إ��Q;��ZGeIZ��X��b��*���@X��O� l�
1��hyr�^l�7��O�D�|:�c"�?���Α�y���@�d #�o��?�����tx��8�V	Y�-Ùgg&��2ʁz�*˟z���e�h�W�h^��A����ȳ��v�b���͖v�`���Ds��~�5�%/���r��1?��!�KZ~��F��?����h���dR2c���f�7g����F==B�I�W��1 mZ�X���P��#<�ODFzo�80�JmC�ݘr����U�7m�O���O~-�1c�Gm��$�O����O��]:v�`�	�h��;��a�n1(��<b�웆'���)����w�����&擏w�8��Q�O����n
+MV-��O[,�����"�H�e`\�P���Y���*1��Q��V1�~LϮ!�R K��x����0�?Y�O<�9�'�b�'��O�X�H�q�����.����$F D� �䙊s��|Z���t
�p��_B}2
,��|J���d��q����U�v����c,_Q�U��1:"f���O��D�O��;�?i���$�,@�2��q�B
j� �`�>1\Dȷ��.l��5�Cgn�l��(�N�H���H6�P(�A�߷%���Q"��f�*DQ �;-�,�b�ׁ'Kb�ʌH�'�J�1A��f�^���@�3<�Rtc�F��?���';x)ĊR�]�ʉ�S��j��l+�'8�1x��F�g\�ad��c��u�H>���i��'��Q��~��J�f<��@މu��d0s�`\K��?y��?i�����%R@�� �Tl��:4�'E�$�
*�����$c�b!�	Ói3,�����,�����-L�?��nH�'Ȭ��ɑ0|U�2IQq� 	@F�O��D>?�v/Fl��U�s+Dn�2�+Y�	ȟ���I�'b�\�`�le�F��%~�����ȟ��q��3L\���Ej��-��O�Or˓~���i���'�哪Um�����\T~�
F�gi\��u��)S��Q�����d@�0l)$��T,l8��2�S�d�?�� D+��h�*֌9�D���"7?�#�6.d5� ��ksVp;����6Xy!W�ʀw�������� ��� �H���O2�}B�'��H�S���7���)��2����'���y��ډI���1Q�݌L�S��h�Ot��#�:m�v���O/q}�m�V�iarY�؁q�]�?�������Yy&� F�X&��l�@Djv�^&���r�͔e� ���\^ƨ����d�5ˠ-��^#OD��"ɔ_j�9�ʗi�"�DNEL�H ��$���
�m� @�X�a�O�DO2��ĩ�#�O���6ړX��-#��	�%�؉pe�0�]Z�<���QJq�7��P�`�cU�Ly2N �S��_���pNϨ'��Ys��@O< �@����p�4�?���?a/O1��	���	�gz][���3D��٬,2L�kj�i�� @��\�FY�����<`Dz��C��mb� Ѥ��y� t�e��$Є�g��z��T/N\�' 2�Hs.��,����u�by�b��?9��?a��S�`�v*�۸.pԽ�Ѕ�"hZC���`�Y�؟>���"�Z4H��Ox1�'�剁_��bL~*!)�P�`!Q�V(qa8���L�'���'��oϏ1���P*�"uhpK��
���")����(86��*���`��#��d}�X�A��m������5<h^�+cjH�	��H5L�0r�����O(|��'L���p�V�L5t]�0J�⛤� �i��(��;�O�}zi�%5oƵJG�ģ��`�#�'� ���8���i�-�)��{��ڃ'�^��H���fyʟP�'�?�Gf�#������ǻw��ј�����O�x����z����jA�'w�̃@�H�'������I�q�P��&\�gQ�'�����@0��	q�c�^�`��i1D^���C��`�� ɧ�ٻ��I�(�*��O��}���� $�B&�Y��b�z@M�"�d���*Ox�kb�F�~��Xx`��@T䁎�DVz�O�@$���7x9$��'E}2�$���'��@���(O&��a��.$p�2�֮B~�P�"O�s�G��CǠ2v�4u�@"O��G�ҥx	��:�)+% � 3"O\��&�D�R�V�XnX�&��Q�"O��Ў=,�>��7��a�l���"O��1�#R6ݞ 6횮s�pCY����o'�O�@h�J�q!RHb��ٖg�=�6"O���C�oݮ-�îET��0b"OBؐ��3�TTi�j:O��9!"OZQq0a�,Iw���$�HL@U3�"O̸I�\Ms�$�TJC�7�PB�'�4���'"4��#c�8���wn�+UX�"�''����9�VH(wEZ�L�б(�'�8�-RWVhpbv@�HLd�'輠�%�0.���ȕH�5UH�'����u��s��*�(j�1��'4,衁ϭ1Pir�o�"�*��Dϲ4�Q?yq�!�"����p��q�\���.D���O�66I.�R�8~wT��� D�L���X�7�TQ{"���Q� $�B�=D�P��Q�;L,�qFL�������<D��8�j]�{�m���ʻF��A��n5D���sㅞI�R�3V�6�x��O�bs�)�S)��Á�&m1�ՄǼ6��'�ء���R´q��Ű
߲%��'H�4��-��1#�A�G#B[���'y���G�K�o�2�C%M����
�'�yhRf�3$c�T�5�C�S�\h9
�'U���") �M�lqA�J٤6����i��(l
�X�+��剣�� Y�����
�5�nq���<�Z9��w}�S�].�I+磁.B�%�'��9���'.r�'�D�@�KQP�k����v$�4�6���\��؀�!�.']�4����5�.�s�	
�� �vb��f^���8w�΀�`$T	S�q���K�e�">!���џL��t�'��1�ԇ�N�hQ�M�r�"��'1a~"ȕ�/��P�F�D��oe�����ny�㘘rf�Ճ`D�D1d��/W0���]G�l������u�D.��4���'��l᳍��
������2Fj���'�(���J� 9t4�i1�ʕ>8�T>m�|:6�F4xKH C�h��7�rL��&��<EJ�3�6�I/�p� 5�.N'�>]���R�W�9c�B�c%H(C5�f�X�q��O���"?%?��'Kl(Jc�.y� �r���^a�
�'KNl��E�+�QƁ��~����y�Q�0���4����!,�<�����,�t:�iF��?!��?i5DS�n\ސ����?I���?	�'�?I󄏥(@��:F�<1�&�3�+�,. ��q�O4Qt�Z ��T�r �ɟ��q�ֿB`f �g��$FB��Bjʐ&βa*D���z�,$���7d�l�'�dU�'NLd~bbOBo|��p@�#�D!Ʌ)"��΀g��';ў��ΦY��,G�w����@6'�)��JWҥ����AK���#I��8����HO���O�ʓ-��<{�*_�S��q��A��4@�e&kiJah���?���?Q�'�?������A�.�@ƋӲ]����%�:�E�G�Vz�x���F3m����r��Z�FŲQ���.8�5�d�^�>��	��#(���Ae�}6� �X�U\n�Gx��˭�?��Q�6�(V���D�8�cF��?���2�D߲T���I.��L��IߋN�����j:J��d�R�2VD��W��PAz=�'247��O`ʓ9����i#}�� �aL�
��S�oȲz=���?A���?�­ұg����D��>��`[�R��:�9=�� k��	�y�y���,|�t">�Ua��Wc����.Cx�����E��(��m)�2��c�}��˂a�O���*�%A9���oѺj������+0�ʓ�0?�ժ�- y��2�Nӑ/����Xx��X)OrekQ�,��Yb��@�i�.u�4U�`���DΟ���Sy�X>���ӟT�QB��'����0FBip�3��\ϟx�`�8d���X"5����B���"��)҃6h��S0 �e�������2�D ?j�UQ�i�.��[���� ( F�T�P%w�xe
t��>sZ)+�����y��W&�?�������t��� Ba)w�� c�.%��M��6�)`�"OP�3$�ݸ.ʈ(*%��$t�T��	��ȟ��FB��{d����n�w���Q��O.ʓ_�2�����?���?q-O��IS�TDE�쬘�b#\D�0��8w,(TXS(�?Y�qb�?鑋}��B�){N��6�Pf��ig��P��t����X�����!f0�ΟƬ�>���R1���憦|�@��	�V~B͍�?q���hO���!U����S� �&I����v�pC�	�y�V�0�X�7=v�2Cϊ<,
���w���D�'&��;3�����KU��|��I�/���p�dşD������Iy��t��[} ���QW�(����JK�$[Sb�.J��e@�	ϴ�*��'k�'˪�C�2z�H���'�$���]�c�Ԣ�ЯR֩1�j��#?!�����P4��)+��d��k���F{B�	'!
#3�<>�ҙ�0�	�B�ɍx�ԭ�F/A�A� ��M�ʓRC�v�'��I�M�,���B�g>E"7FP�Y���EHؘ)t4�����O������O��D�O�+Ta�Y�J) ��9?�'Es!�wiN�z�ܢj�XCuG|�M�6��M��[>�Q�-�~�U��T��G"om ���m�'���Z��)�$(S�����	� 4�� �_�!�D�9gp �q�9",�q��+�}�K�<�\�!�����i&� G�Fy�'w��'{��'��ɟX�'Vܔ��W�|�A�%Pk/lY�'����{��cUZ�sd;.��taGo �%q^����1��>�?����4�G1l���J��%F���B���)��0@qP��|X����ʟ��ڟ��]���+vBN�z�����#��ܚ�9� ��M��b~|�����y�����������?�،Q�`��ənA�X*���8�����'�"$�$}�|��������ߟ`ϓ2���2����q"1�����(:�MΟ�iY2ů�O�ɖJ���s���TW?���ט��ɋwG/5)�S���?�(˟(��9i�18��u7�'��O�$���]L8��T�J�]3�G֐Ubx�$�j"��'Ld-1�'������u��j��3��x͐*$ܓs�81H�oz���0F�x���O��	��i�O��D���5��f����D�h3�'ܚ
��R�'c\����?!�����s�C��@�?�o�)��d��M��cl�˅,է2����	�M�&�'�������?��mZ7i���	l�,���	@$thD�./�l�x�4b�\Q1�'�����?����?�'Q��b�O�,�2 �ٟrm|���\�RL�B�i1�Cc�'��I2�"ߴri�W����5_�e �M/�E���Ӌg�`�ȓ>����'���y��(�WWjElП$��y"*�~���?i/���L#Io-0c��������M���?q���?���?�)���OF�-ar�^.H�8pf�+/ +�}�'��O�O򥸥"�,������L��4���?!R��x��ř{g�ٙ��I$,#q:SG3�y� @�ha��[*�aR ��y�k�7'Q��P��"x
 Ʉ��y�N�754±�X� ۊ�r�
� �y2�
�I��8e%R�`,��YC�+�y�ܨYv���w�K�D��01dm@��y"ω._���ɳClE1b��-�yrɌ;"Ө���=��1�I��y��\������ߗe�����L�4��O����O��$�O��D	�k���&�8�����#H�d�Hm���D��؟���ş�~����O��d�O��`#d� ,�ݡ�H��3!*�S��Ϧ�����T�	ğ�	ޟ���Пp�	$��
"���je�˂A���Y��M����?	��?A��?���?i���?�FDG�s]*`
�b��e��$�o ��6�'�R�'�'���'1�'j��,o�&\A�e��z0qo72�7�O`��O��d�O���Ot�$�O����㜱��'&> z����=ZLmڟ����	֟|��ԟp�	ޟ4��)6�&�z��̦#���� �,[ޭ�4�?����?Y��?I���?����?1�,�<�j�o^k���� G�%�X0�Խi�b�'L��'YB�'���'��'�!;�� bxإ���ќ"�V�2��{���$�O���O�D�OX���OL�D�Oz�J�	N	[:�t�d��rDĉbwcI��q���<�������0�	��L���0)�G!��x0�� 2�Ӡ���M���?y���?!���?���?����?���RJ�E�g� [���Ь�.����'���'r�'��'��'"@I3^l��q��@��p��k�7m5?)����+�'!{�X�E�2-������#k	��43cj@�<���d�`�n�It@<S�̛$�2�Ӏ�+m��l�1�M[�'3��`�Jo�|{�B������B[�Q	Ɖ3��
5�Oz�(AŖ�e�(���!��|��'��pQ�Y}4��mE�2 Q����d?�D��i��9�K�? �����>t���(\&�pB3��G}��l�xl�<�(��1*UlȫW���7N���i: T��CCn^2re���,?ͧX�޼�WH��ybG'@���#)*UgƩj.î��<a��h���\�%�(%r���R��G�k�kuӠx���:�4�����I���h�f�#m����"�E_�i�P�n���@SQ��$	��`�������,N��]�I�$�!��̽C���qЇC"�Ң=A����D<�����ɇ ~��<�0$/X˓~_���A���'��N�D��[�n�c�����ʲ�_}r�`�
5o�<���Q<t9yatP;F��eȥd�&:��q�d\�n0�I�M�x��'G�/�`F{h­�H����F(������w�2Q���'��'�7M	���D�F�;W��v�	�fY�t2BIx�h��s���4Pʛv2O�,�T������T�56!2134Ǘ�U��0�'� qc3!�DT�!7,�Znz���D����K3�^�V̛�ڻ8[n�hF]ß@��|yBS��~2��<Z+,e[׍:}�~�93��{�	��M#rƅq~�@uӺ��(?A��[9��S1@Ă`�ҙ�# ��<��O�o �M���1b鈴b@�<180hxE+�$��ЁS��4bxu�.e]�,Ŧ\�VO��|*.Ov�I_~����J��Zh���".%U&��?���ᦍJ3�/�	�?I�';h<�a�H9s�>S�fQ<M$��'7N���6�n���Ii�S�?�C��:x.m@3 ѬkRԹ�%bd?НB���7R��ɭ����o�ӓf�;�ēsߺd�G��6=�ry"�A��D�#6U����ky"���OΈm�\ʶI��.O�^��������u�u*;?q��i�|��y�wӤ�$섦9�X��rd ��� 	�ᦑ�	5t�
�aq�, tIMӺQ��G7O�i�d,@'�*�P�p�V4!���۲p�˓�0>� 
E��|�4)�(?+@���&��Mã�\�?���?���+z���2wTܱp'Q�TMz�
eF(#.oڒ�MS�x���$/"�DI�']���Ū��Hݞi����'O�֡���M��9K0��h�x�N>Q(O��hC���E�
o�m��7U�2�F�eӼP�P�O����OJ��⌔�B="���*����3�I������E��45m�'���@vԤ	��`�Eď&*�!2�X�H�%;K�b�0v-Hp�@��� �(�<I"J�"7���S��6�Tx��^V�<��M� �޸�4���I�D0׉������4O�0-����?A��i��O���\-^�Z�k��8n�ф�\�����]��Ub�46f�ƥ	C�n�'����5~>�(7l�8j���K���.ua��v�nL��yQ����ԟ$�	ʟ����X����z�J��sk�=[_<�K2/�dy��i�V ����O"�$�OT�� ��T+nJM҇K7R��EY�IYr��y�'�f7-�Ϧu�ٴP��O����O"��m�2Yz�����;����]��'���M@E�LpQ�M"X�_�,J.O���u�����b����0��H���O���O��$�O��$�<�W�i	|t ��':��f+�
ۜ�:JN	j���%�'h�6�:�����$Lߦq��4%br A�JP�r���Y�m�B��bg`ɸR���<����M��%��
-0��Q����s�#K�^ۖ�hb�`z6�ĝN������$�Iğ ���@���Obږ6P��h;�	@��ܠ�n_�$����h��4/�8ѳ���?A`�i򕟰P�E��J���BG�VL*���K�>�M���iX��N��"�"��<�� ї�MS��	3X�D�)��6И`���'~�8�����"�O�0�+O���O����O�(I�������`ԛZ���a���O��Į<��i��*��'w��'@������A��A�� �?!���.�	��M���i��O����E�D�7)����pb�F<4�z�`0�NԎu���'��4��7m=Fp �'�6$9��$��7�������_R�����(�I��$��P�vyr�n��	" B̉5���"�زk��9 m� 8/��D�O<(nZ��$�0[�O�<nZs;x��$����+G��G��tZߴM���@���ɞ'���ib�T`E�ظ�`˓V��}0a��O��	��6to������d�O����O`��O2��;�Ch�w��@��&ϡ:���b�T��M����?)��?�����'h��;�����J=+��D�?�:�H'�}�lm������'�2�^�HH8Γ ����2��2����]$f@�0R��\><*t���ߦmNER��~��|y��'Q�X� x�Q�%��&����A-`��'o��'{剃�M���?���?ѡ�W�m�( p�.�p�$��O��?�N>��\�h�4����0�D�L��|KU�"@r�L"���@�V���O�6��b�a���[y��O�*�H�FU ~*��>t=
0�R�LX`ո�dՈ}��'���'w��<��DZ^��A�U�R8A*0|��O�Ɵ��4x�Bl���?!ַit�O,�����@�u��57��#�E�^,��Ҧ��ٴx�F�П({f4��'Er�i�p�`2�H�[�c6N�P��&��4�@HQ >��<���?a���?���?!�X�-	�Ѓ��v�"���)����ɦ1qVF������՟�%?�I�"����GcН7qx\�2cXg���#�On�m��M�Мx�O����OИ��� ��#�dq3+�uP�fQ�0���QT��l��y��d������$��,�����[
P���\���$�O����O����O��ϛ�'֞q��� ��Ƭ�9Z�l� p�l�<�@$�'�7-�O,�O���'V6�æ���j��#�k[�.�8������DÍ�2�x�D}��˰A����-�<y�g�aA?(>��0ƈ�����M������l�I����	qy��$��
+�� �1-��&)C�?���?9 �i�$��2[��
޴��'U��$�M@{"�˖+y>�(e�x�w�h�mZ�?!H��<=4�� n�5-T)i��߃+\��)�.=��������e.=�H>�+O&���O��d�O�aӐM�d-��ސQ���O���<Ѳ�i���1&�'��'j�S�S�R� �S�pI�M��~1�I��M;r�i!RO���4�V���/ �j���5�l��A�i�"���D�9^�x)�'i��'I�t5���|rU; ��t �Gϋ5r������=g"�'E�'�ҕ��T����4Ms&88 ˒xyy�	G&M
��@!�L ��D���I�?��Y����4b��h�6�N�w����m�G�����i�@6mM7Ȗq�5O��d~Ӓ��`mЯm�|(�'��lA�A^�=IAL^�VP$����'r�I��	ş$�I����	Z�4/�2`�Un�(�D.�`޴&�ĈR��?I����*���Rݦm̻pMdB���,T�9FI��`01cߴ#�6d'�៌���@�8�������1�T*�U7FC��JK _��hӖ�X�kG@}$���'r�'x�+�n�i��u[`d��x��V�'�2�'z�R��#۴Q�R���?���h(����ׄTIz�[r�I�c�8c����
���'�MKS�iCO��20�B*"�]S�Z�` ��a���O���z�b%p6�ā?�>E�'��d	[.�0�D=O��5d�+q�`4X��ʏ"� ,Z7�'{��'���'�>�̓UiT]�w�J
�9cj<Ds���	(�M�DɎ�������	d��?�Җ�3[k��0�&�¶q��	��0��4Ri�ca�TS2�ζL���OD6�f�j���qs��#�"��".2,Ƹ'�,�'���'���'Q��'��}���J�͙�T1�Ġ�]�l"۴d�|�����?����?�aě�cf湂$2ir�ع���a�	��M��i�VO���&��]��ba��M�.�$|j�e��
0%"��ח*]V��M[s���9�����|�P��9�Ȇ�j�^9v.Z)i��D��۟,�	ߟt�	�P��}y��}�py���O��Ʀ�p8RV)QZ�yҫ�Of�lZ� &����O��mڒ�M�1�'O^��rZ,�cN�'�.�
��*�X��?��49��d�C�PPo�I�?�̻"YԵ�� ���Q�E
&x��h��'lr�'\�'�RU��>�-�̔����&,�Z����O���OJ�mZ�ɞ�'j7�$�I�U�����Ц�2�#z��&�L��4#����O�dy��f
��yR�'��âTM2�%� ��A��	Z�t*�BQ�'Y��O�ʓ�?q���?���Y���s�Ļv5^�Ȧ+U��: ���?�.Ol�oZ<}�]�'�r�?�K��*�����/�1w����n�<�e_��xߴ5����)�4��I׆z�L�B�:K:V�4�ň'��6���gl24b���{y��Oݲi	�H��.��'Ԅ)
���CA�VIV7R<yiS�'s��'�b�'n�O��ɖ�M�W#��M�I�/K�P%¤��$�+4������?�C�i��OZ��'L6.q�T,c̟�m����F �n�MSa"Еn��ϓ�?9�4ih�=�$M�M��y��-�`�G�b�����Ȃ�5|����`y��'^��'��'��?��7cǡȸh@���	2e�@U$���0���ן��	ӟ���N���'�"6�e���w��! ՘�fD� �zp�G/������4B6�'����O����iF:蛜'�
 9�	4|�@��sb	3IPA���'+���~�4��)�䀍BB4)%i'?�&��&V��@Z���koH�§O�<1��35\�a"�k�NP��#&�R�<����& ���?d�2I��L7?I�=� *@Mȡ#7��Q���+%��`�N`Un˛q� l���S�X�`�h�j�l�^l���ϩP��Eꦍ�\���!�hƁE���jd�X�t�����O�yʅ��TD�R��)7�ԌP@N�X�2e@D��%f�ң���Qj��Q^m�8
�@!'��,H�`л���Sw��c�
�Hc� �d��
$O� ٕ*Ζ:Ԅ�%��?�d�2��G�G���iQ�����@���8q��M�]s����b��	6�L�a��S��԰��Y�#:��: bʃ�H�%NMQ���̡޼�J@#k��s���`��jϐH��T���+" q#��L�.\)4MO�!�� !�p iuoĚ\�0{�*���hM�S�8	��y��(�ɰ��ܹ��`Z��(/Eh�Q�F̦��ԟ��	�?9�b#��Nx(u�^i� ��	�K�I͟$�ɜu���yy��'-�i]$H�X�ǀ�$A�Q�DL�o#��'"@�B��'���'v�t[�d3���]��eQ>T[�L2�@����՟���	�l��c��>���E?Pyģ�ك0��Ƞ ��O�d0�F�O����O��㟐���O�ʧ<�2��vӂ���Xpj.�~����5�N��w�r�S�O��(V�L��عe�C�i���2N�.��'���'�<�i�P�\�O��1Op�q+�[&�R/F9[}�u�5�X �'�D��Đ�$�'���'��0ANZ�*@�r� s�����'��H$�"�'��ǟ�'����d�6w$�Y���~�VnH��'h*3�l�����O~�D�Op���O�!{��$vٮ���)Y)b(<�D�4����O��d�O���8�D�O��d_�P�Zq",�DI�f`,i����j��	��(�Iݟ���蟜�� ��|:���$u�����ҿ9T`K�eߟ\����x�	r����|���D���&ԥVgBTGɔ�Y��lzeD�A�v��'��'lW���!L���'�� ���v��4eH֮\�3�,EpG�'�B�|R�'�¥�ܸ'�8H�ʚ�0�����H���TH���?y���� T�'�?Q���J���j���5��u��#ʼ�O����O$�10j>��?щ�I�g��Ȱ�Gʦx�FP�H�O��W*صb��?I���?����ɫ\Ҭ�4��n����U��eU���O��$��Y��$;��	ĆM���qEP�0�8�)a.H>KX2��=2�'���'��S���I֟x2$b���B�[�̗/th�����Ο����Uz�S�O
bh��n�"X����e\XraP�`"�'+�'[d`�P���I��h�I�<)���84m�G%� G�Pmy��O��|�^A�I>���?!�qQ���A�M*>�lp�Jߍw,2� ���?��c����O~�$�O��O|�xV,Dz�A�	Y>��p�1ϵ<���(�䓈?	��?�+O�m���еs˚��̚�)������#�H˓�?��?!L>���?����|���r����Nь��u�ô��O>A���?����򄎱�L�S�?�����Q1p!l��t҂I��$�O���O`�O���O��3�b�O�]!���)m���R�kF�1<�h��a�<����?����$�;����O���L>KK����j.��y���_���'X�'���'�p�;��ʒztI�WC�J�` �/ȷc���'~B_�g%@^��'���OZ��h�j9F�\%�S�L�>��`�|B�'�n�M��O�IS�;7(�n]�v��-�#ļ�bS��(b�EL��̟��i5֝Jyr#��| 哱�$���l^�tv�'*��N�#��Oq��Ä�SHV�Ar1$T;'(��a�'T^0$�']��'c��O!�Iʟ��I�K8���e�?�X���K��m��t�ɝBT��?E���'�n����	4z��]bQ`[la@���',R�' �bV�!N�	���	럸�'6�0�a��:}��[�Іm�2��?IC����?����?�A'͍s���K���JV��n�.�?1��ZR��Q���'��|rQ��I�J��+a�ܲ�o�'��	(fi��%�������	~y�ɚ�6t9Ш�A@н�qL��ذR�����4��B���0�I= �~�8�(A�^��v(I:��ecM�	̟t��ȟ�'jc�2�����K�����C'<& |�c_�L�Iޟ���}y"�'x������@U����Q
�_`8(���6@��'N�'��	�8\!�H|JFsO8��Q��:$���y�)ҽ�?9���?I*Ol�Ĵ|"������?3ڕ��lI�-!"��4+�3��'�R�D���6�ħ�?�w�t�Ʈ�S��Y� !ˋ"�"����O����O��d1�9O�}"0"(	���2.B�Kl�Q!��O �h�q�i.����@��	��B\B���Gâ�h ���_�J%��'"�'&�P>��'
��zZ�-�F�A�
0�g�	�Y-D��I�K�P�
�4�?���?I��*����������Ƅ�
�|��^�2�\�Nc��'���'���T>ŗO��+����Z(Fɖ���'Ab�'^R� �i�)"�O,�FHQ�p�z�r��P��<�+�'ݠ��'�j�F���Oh�ɇS�b��6f˰uh��`�XZ����On0�W��<1+����H��:�T���	�<B��A�'c�Wy�o�%R�I�O��D�Oz�$�<�oW,`�&�ID�S�̕`��%�@�BA�x��'G��'�����I"2��$p�H�}] 9g���-ޤ�(��Oɟ��'�'��П��tLH�|J%j�&���`�nA��K�H����ΟT�?���?GR�zV��`Si�!-q�A����#��!y��G����?�+O��d��7W�ʧ�?��G�bG<0Swd� ��8����?)���'�"��$�pN�(���~k��A���R霔�׬�O$��<y��d�T�.�L��OJ�]�X���z���
N�����|vʓOL���O)#�Η81O�)N�+�2Y+��ƨ�@4�	@�rY��p� R�M#,�����5�'~h�g,ִO�P�:!��D8hT���?��d�BD ��䧒B,��%� nG�K.H���. :�ٓS�O* `��JϦ�����P�I�?��I<�'u�2O�+)�����m$k�5H%���?���?�����I�| O΅#�͙W�܃�2�B��R#�?����?�reu�+O�Si~��ңH�čX�?HPT�<I@����'�?q��?Q�E`!�d�� ��[�jD� ���?A�N�THxB�i�2�'���'_��'�y�9Q^����%z��ݨ��ґ��$R0���<����?����?��7��X�땠/��k7��!x�I2g��)����'��'�2�~"/O��M( (�)�b��I��P��$��%6O����O��D�O|��|��Ne�VV�s٘���'V	~�̅8�%�wl��'w�'K��'��	��z#�|>E��$Q4qrN�����Z
,TpW�ϟL�	���ϟ�������5��M����?ц�U_ɤ���D�M:�H/ЎQ����?a��?a-O����.j��Or扖m��0v�$�$ॄU%/���O|�d�<�c-�_(��柴�i��b&Ŀ4&ڄ�A�'s�1�ÎFjy�'���'��8I�'"�'���Z�U���%s� 0���N�E��U���d%Ě�M����?y����dW�l� ����K$9���C.	~F��+ �'�2�'�"�k�'��Iğ��|r�I��\��]b��@5(Ʉy��*���휔�M+��?)���R�^�x�'J�CK��e���|\��p�'X�K�'��	͟������}c%HX�F[�]��H�/��� D�i�R�'�2F0|����D�O��I�p��r�?���fG	}W����<!�K
��9K~J���?I��Bc�)y���� !�aP�A9z�Y���?i׊9��Uy��'a�ռCd+�$)�Z���o���q�E\My�ă��y��'4��'w��'Y��%%�0)��6�l��p�_�cRX�z��-����<������O��$�O.�Y��F@F��cZ��Υ��^�D�O����O���|Γe�����O��ɲr��Ip<����D�����Ovʓ�?���?�'g�<�R��K$��:7
ݹLH�p�!�ܵ�?����?��?�-O��w/�R���'�n�)A�Q
n$u9b���hpp�'U�W�t���P�	�y�,�IF�D��,�!b�q�XZ$�H52�'"\��h+C��)�Of����B�H=B�DQV��M��-�Ï�<��?i��S�.����9ON��?�����%2L��cA�$�����O��dʨ1��oZ����ӟ����?��	 16�m��R��	b�:H��}*O0��Ȼe�"���O���|�̟�P��\�&i�	u�ч�'E�l�b�a�����O��$���4�'u�	"N��5�v�S63ь�w��|�Z���v��	a�s�'�?i� S�����&�?p�qc���+/���'���' ���e�O/��'�'��⍨1�h�sf灝,����ުtR�'w�	4[��1$?�����\��,�d�
�gͺ}Pxpr�E�����I�<�9�M����?��?�T?��39�q���),,��G^�5�b�'��@��'��I� �	����Iߟ@��f�	W�B԰U�I/�āj�>tV}k�4�?I��?i��g���Uy��'�p����E�Q�ॱ�D�
8�(t%ژ�y�]���IݟH����,�	63*��޴'�i��L5����b=un����?��?���?�,Ov����I�+*2���*Th@�h���`4p�d�OZ�$�O��$�|�d&���'1"�G
�eO��_�^X����
����,���@�	ty��'�Z��O�b<O���_� ͳC��X�RЛR�'���'b�'��m��tӊ���O����pPƫ�&S(�):S�J�\��AA��O��d�<��}dJΧ�?�����ەId�B�!�*z��S��S�;�b�d�O��dI7)ɺ8l�����ҟ��S�?Y�I��.C�)����G8&t�Ҡ��<���\q����?�(O�i'Z�FO�FC|٤$A,aX
=[`�C៼C��U!�M���?q�������?���?Q���)�
�5ֺ<��q�TO[��?�5D>�����yB�'3�� ���<RĨ=P�01׃n���$�O��-���i�O����O����O��ˌS�X�#�'�bp9q$V*�?�����U󜓟����O���7-�f��e�6����$�#�l�d�ONݳC��ᦁ�	П�����0��~�ɩ0�����kHjq��Լ/{��8����<mn�@�$�OB˓-,<D���R�
xr��s��&@'�Q�6+C t?�'���'��'���'��1�m��S����c� ����ӊ����'�r�'�"^��ӓ�L��JwCÍh9�5���k�y�p.AMy��'/�|��'.N���y�,<���KӉ )�Er�L��2���(�	��̔'�
���:�	�2�l�x��  ��c�.�>DJ���O�OH���O�eY�;Op� �Dt+�*о:�!��&t�T�I���	Qyr�S 5�8�d쟚��D+G"��2�-F?`P� �?��OR��ܛT�p�$>�ԟXXp��F7s��(�`�7V��b�'h�I
�x%9�4���O��)ayb@�z0P	���wd��K���?���?qn$�?�N>�}��J_�]Ƹ�K$/�L���P�e^ܟ�X2���M��?����z��x�'�b5c��M�S֐]�Q'7FYs�'
dt��'tɧ���_"I��(��F@,�"��2�����(n�Ο���D0�A�����?���y�b�)�­ Rg�4�,�&��+��'g�驎y��'$b�'Sx)�K
�PE�{ae�8]J����'�j��@Ob��O|�O`�O�  ��h����@� d�fˤ<A��P�?�(Oh���OV��lx��#RXl��*�5)�J���J)�%����ş�%����ş<#�@3V,f�U��p��SUV0'�h�	ߟ���Ry��L=b�J�I�,Jp����13|y�a�		��۟���I��۟��	�d� �I~�p=�6H����	�$��Cz�ؕ'D��'�rW�鵉���ħd�:A"�mϣ(��1@�������?9H>���?�qbR7�?��O�5��ɭXfZx)�a �60H%�'���'�I<*�T�aJ|�����$.�
�����\����ڗ�䓍?	�d��}�����SJ6a�'$���p"��>VJ���S��x�'�@��@*x�f�'�?��'.��I�pڤ�W���}Ŏ���o�	^��d�O(��!d���D(���͹��a�
0��M�"	}JҦC�g�6��O���O����U�i>����R>!��H�$�T��,ԆD̟i���<����D�D�'�"9Ѓ��Q̸���ܯMDԂ4Mr�B���Ot��A�W�vD&��S~
� R������"��,���,��UP�'D"�'�i���O���'�� ن]$�vGM3*T�+�&�I��'s��#,%�4�d"<��Ù��܂P�̎l6t=�&`���I0KB��Iqy��'���'�R�'*��p.�%L�p��&�3&\�AM���ڟ\�Iܟ�'�X�	ܟ�෭ƞ�ژY@EW�"nŨ�-V�g>P��A2?q��?�����+y�j1�N}��r��A���� �{��ʓ�?����?A��*í��'�#�P�6,�$N��C0F̷���O ���O��d�O��8'��O���Op�Q�B����#ZC� @�O6�d8�$�O4�U�(���Y>�uć�{`h!X�'���d�yנ�ܟ��	ʟ��'�yq!�>��O��IE�8+:Y�놅c�ʰ�'̭p�`�O���O�����?U�Sk+ru����;O[����O�OD˓=�-Y4�i������Z�c�(��G
����&�7D���'}���Oq�t1�p�� hӱOZ��z)"햠	�\9k@A�3�=iQ�7+�����<(x�-ǿlUl��%,	��� ��쩺@�G�\�����ş�I����2�.��?���?��cq��'4�Ԃ�A��aA����?9��?	����#{��3���3Z8i"�K7;�.:F�O���O.���O"�O���O�� *W�a����)�H�)v*��O�����O��K"X�� �A�~��'N��d�O�b(L�C1>�1��� ��Q��$X����|��'�8ڗ�?����-)p^�"o&pJ&I&�@�+M��i-���͂��qon�!��	OˊUpR��9"��h�T��h0�DEd��l�vȈIs�4+DC�8('��T0���WH8as��'?@�U*(<�@�5�XF�9�O.������P���׉�mS��K Ȧq��T��2N<�yx�②
uhĻ4!�~�|;�^6a��Q�d�'H�a`3]E�����]8��Ѳ�&�a�s��4L�^)f$�c�0X�F�麋0H��y4|���V�h�qj��Sz�����O~��O����#ۯ?x�H��I_�&kp���L5��D�	���c΂=�2b���Y����@��L�� �Cf���.�6�T�; �P0��Úv�J����Ox��c����n��L>YB��՟ ���J(ry|p�II��
�	v��8B�!�d�.f��� AK,X�H��G��6L��D ��|r����_�n�����#��� ��cc��C��$�O��4�hճG�O����OP7�MF��$C�!���X��ư.I�<�G�z�3����?ɀҟb>�&r�� Z4�Je"�J�<�
xQQV�nnn�+�j>"�*�$�O����M5�0-�ê���4R�W5_�ޘ��ݟ��	ӟD���>Acj�2(7(A��eB5`Jz-8��O4�r�'@
L��a�#B���!�?}�4!�{� ��|2��M;Ӄ\�b~ �QV�>������μ3
"��j1 ����'e��'Ҡz�Q��۟�]�rXpx�q"�2#ʠ� 
�)��c���H��
��=�*��#��D�D|�ѹ>vRux�KR�oL��\�=����Yt�����V�F����@I�Ь�j�l�bC�;}��.ɀ��I�9�$=��L��MC@����
���d;G}�șP�G�K+��H}� . �~9�g%�.�n��# ,�(O�=mZL�	�<�{�O[����Y67qzuR#k�p�U����Of���O��J�ܟ\���|jV��-h��1���	�� f��&T y@�^�Jy���R�����<��F}�x�Q#Ȉf�� �Ԡ�1	�h1A3j��Ao�8� ����<yjUܟ��	զ!�#�W. �3��+ބ-��  ���<a4a��]ߌAk��3�����[~�<��c�*Bϊ,I�dR�6��KU�:�(7��O��-a��IV�i�"�')��(��H{��	��8��߉n��ܢdM�����۟��d��4Z,��J�&�:�$ `�a��X���� ���Q$�$A�8�r�	�U}�$bP�c����B��w� ����E���p7k�i/���ٺu2�,�3`�^ 91,3L0�O@��'�?�	�Q��@	��<�P�pG?D����lF�k)���ǡɎw�M��<\O��=�EJ��'���r��!����[nB�x�e}�P�D�O�4�8�YAE�O��$�Oh7M�P=���a�׉d2@��FQ5W�,�lZ"h|M[K�8wS8(�f��?�&?˓Qi,��eB2sx���̕��v@�)X9��r�A�S����ODk�OA�牘9b�V�^=A�:��*l^^�	���?q�T�hi%�.���n��z��q�l�6pu���7l��H��Z�	|X��;�F�x�ԯH�<��էO���?ћv�'��y���|�$~ӌ�r�BۑP���D��p*���H矤8��Q(�-����$�IΟ��\wG�����w.�B%&Ȫw)�bnT�GZҦ�v(�O`7b��TL���:c�*�c��f�$�C��'b��SD
2*)d� 
86k�a��40p�x�	Пl$�l�	ӟ$��1����-�<�5�L��A7D&D�܂�R�'��1˶"�N��<z�L2�X0��'v�I;]�B�ٴ�MC�C�7I�>ܘ���=�� p��I4x��'X��!�"�'��IM�H鬈JL���7��*Bf�f�v=�| TA#����DS�up�M�G\�"쬐� P)��˨5Qb�z��^S��H�U5t<{0Np����5��&:�p�d�r?YMY	R� 9[E�_�=,��Ҷ�Y�<��ϑ(#ν�f�>R&���R�<�&m&	���r�ʘ�lnJ���Dh-87-6���,�Htn�쟌��U��@1ar�Y��n�5YAt$H�~��x��'���'W��D
�Sي���<�O�Ǒ"B i�Q�Y~�nx�Cb�m�Ol,��*3@��V�h��p�$���i�2
�*� �e�c�@,�Ǡ��c*�O�5�q�'�,6����Is��E���Cϙ鞐�����@�,�0�r�����j�xH*�lf3�㒡�d_f��ds�;�YZ3!U�	9f�H4R�*><e���Ġ1P����������61<��	�x�	���*��I"�*6OȖR<�р�ٵ�M�C�e����.�?	s��'��O�@�ɩR�x�3�3?��)���?��-�4&6J�`K�
�V�T%Q�k���SgP�"	��'s��-8��	�c�+��|���9+Lс�mx�',D#}�'��U��*�=��Q�bv�8�!	�'Qb�k���_(��CjH\h"��{�K7��|��O\рd�2�����D�ol�������a(K�3�T���ɟ���蟄�^wg���Eys| U�*o���cO��]���4 �f� �$	'\OR͈���U�6p ��+�.��0�ؕq�,A��7�Z�1�Z12�����/��xxv��Z����쉌H���2��?iW�i��7M�O���?YM<i��R�S�%�'��JV*$�G.U�F�ў"~�I�d=�=YEeˏx��EX2g��4��tk�i��'x
,��O&�O�X�!Xw�+P;{���%�D%ae�[�'�9+���$�Oh�dF�q���O擴V	����L ;�N�� ��\�B�G���"J�		P#�佇�I)&(	yS���&�Iχ �}c�dS�d2g���(��牙l���>�P����\s�Z�\��c�-Yq�<y� ��8]��	��V�c���p�<�l_�g����tK��>�F ��C�Q36m2�d;�tl����I}���J�;
6iI���w� �EmVy�C�'���'G�T*�`єl�ial�<�O�˚m�@�����a�T�iʩ/�O����On�+�I+�'}�d3�&V�fQ:��IڄO����>���ʟ�۴v��O��S9(y��S-�^,��HF�ñB@���b����	�H"���B.�n��&�'<���f���TO)� N`�ѧ��=�>�J��̄""x�8DkX�u���'K�����G>#q��'%�iq�p���x�4� ��"_ �(�A�O�b��Q��hO�A�G�,B�vqق ��GEJ$�(M�'��#}�'�><�(�7_��PG��n/,���k�O�4'��ۍ�Y��@EN�Z ��j�%WO�3u�?D����ȸ.<q���\r
�J"+<�Ɇ�HO�O@��s�*[\��j��p \��d�OX�UD۞8���$�O\���O�����?������	U�.�ڕ�'�r�:4��X�x�Reɡ)P�N�8 *?���]��O�h������S��3&7tI9%kА"���8c;v��j�e`��N9eG؋����#'i⤚V�D� ��j�#V�F����M��?A�'��[l�i%4x`��֣��)��';��j��[PlN ����9���ً���-%�4 ����Mڴ�
I3� �4~Hsɑ�a̢=�`�'Q��'���pv�'�3���s�l��U�x���,	(�eoK� �A�H#A.���ѿ�H��υI+�����f��j�EW
Y��9�pa��yZ<l`� 4+��j!��O�����Xh(��2d��$[��R�aў�ȓx��Q`�EZ=E�\!�'Dˁ3$���}~ΰ�&�σt�i��I�'+v�Y�s�f�O�0)�kQ���	ʟ��O�|��L-	�0���M�M�f�)�����R�'���υ[i�Ir�jR4?���|^w�J��˜%d^�i�#e�H\��}"lU�!�~�k�b8�H��-��L�K��X	dfN�0�|
v�L�2�'(�O��Gb��#`ì8��NM���p������	�i��Ux3h��!Zx9���L'���D�wܓ/���C��!�"u�@�H�]�P@�	bюPl�柸��ڟ�Sh3�i����T�	��)�::���Qd"$T����5z�n-�P���($.��2�'���S]�g}"H�
o��0Ul�t�(4Y���쩀u�C�,x �M��U2�Q9��Y�h��gY�>���ɟ�/��?	��|r�(�g}-��|�V�dcD;jk�S�K� �y��W�x���kGH�"fẨ��ĭ��'��#=�'����&/*�p	��"!�L�@b�.����I�+юjȟ����d�ɠ�u��'	��[)�|C�eՎEJ�EH/9���_��[�+T����������I P�����_�B��/e��H�f E �!��O4@)<ā! k�`C�FK��� �d��-��0�����C�z���5�iv��X��?A���'��O��� W��t(�B�&2�H�j	�'��4r(V[HV@��M�0��e�������Ity2��V�7nӄa��cߧZ
�m+u�]$6,��EIXΟT���J�d���I�|�%P�T#v(�F�eP��R��9J�,�s�J�jk����hθ"3���$Ɵ	8v�<�r�J�j�8ʂ�#]hH!��O�^�e;d����Dh�@���e.Ј��\+w)��<I�B�ޟD��'�hL 5�A�RV�0�1ꑉf��́�'D�DҵBU� I�F��e��`�<Q4hϡi��l�#HS~AK	6E|78�A���n����^�$�6<\Xic��C�D5I!�nѼ��q�'��'���Uˋ�(��X����~*�l�]	Z����Ow�©�r��%yM�c����RJCHLPghZ�"�
����p����&7��u�ٌ�^�{���C����#�o�4)�W�����9��A L��݆�`:���R��	��!�v�Y�DlԆ���'��s�삀X� s%
B(i2�"E	�>lZß��Iϟ�ӊc�|1��Ɵ������MN:Kޔp�OН^X\LY�'K�3ڤ�Ғ�ə ��	����Y���F_�
�,2� Z:N����ҷ|h8�(�L�2c|9�TkN5Ld6i�������Q���p�ˮdI�C��ѕzb&,�d�T����%X
���V�	�0�ph@��I�P�!����"|�S$֢+F�`R�H�qO��FzJ~b5�B5-�(Kg�E�n� "(V����\r�ɡ�'�2�'���e�E����.٫`t��B��[eh�����>�f��\{���_���)�BM^8� ����#�H�`�(��9 є$	X6	�B��5�ܣ�Oy=�]}�F�Fy�뒒$���Q.xl|z3 >�Mk�$�����{.�UK@�<W6����ክ,RхȓA8}Z�iܪ{��zU�>��Ey2�!�IWy��x�'hT)C�ߏ�@k�%�3��Å��Ot��Oj���
�O��D{>Yr�B��,���ЪJ�E��dʷPT�c��5!nL$�'� �Ң˅�d F��/T��t�1i�e�VE�rn�&`�@A�B�,�<�ɍ���(W�/lӸ@�`��N��АME�P}�t��.�2fV�|�)�gyB͂5y0v���#�H2ܰ����(�y��Kz���j���*:��8C!^,B�F��'�	
��zݴ�?������T@d���˵?Dl�rDV?}�՚�$�O��D�OD��\�m�,�c�F.�M��S����D����dklљW�\��RL���DϠ"w��A�c��NL)leܧcvz�qG��2|v��	��S3S@`��>���џ���)�=�����4"��e#�d!�䖭�Ұ@E'@?u�����)G8�z" :�2gZ���딫y��dk�@��{|)���O>����'������ϾQ�r�'��i�D�x�@Z�{�&�1SC�~�:�`���.@��������d�ß��4�Y��ڐgFF��} @�˅#�=��.��?y&���1�V�3��	ͼ(��a�r�2�Ry�;Y[ȅ�	߫l͓@i�9g$�x���'��O�hE��OVmJ���$��t�N�U�d���"O:p�w*Q3U*�F^�#�d��e��n���'t�����������i�+}�A��'�P�[�(׍-���'�B�'����埌���~Ts����
�.N ��1�!dJ�$F�p;�(K�s�x���I�-.~�?�FÝ�$��Ւ�LT�sv#C]4R�*���6y��i�V��"g`�����B�h`{k� |�~����m��6H�?ɐ�'@�<�T�יJ�^���Ћ.*
�{�'9��3&�)\���9�@�� nny���IX�"Y��q�iӛ���DfQ�B&(����5sm����O���
�����O^�ӷ�b��2(�,c9z@b�̃�`��5脇P3T��X����n�␫�E��]��	"��Q@-_�)��K�D?v�F*�j��	��'%��#�J��� ��I�5� �	]ڡ#Wӱ�!��� ^�AB�",d��,��r�!� � 3��A�@!Tɘ LCQ�,�}b+3,��7-�O��$�|���M�
����`b�	:Д4a`Δ�:����?�����*r �������'����c�F�O�j<Jj�9���`�}���H2� F�4㒙)�B�k�m�:��j`�֙��'���ygQ?�c�/ʋ,F�i2 hSU .��t�(D�t3�O��H�t@�],E���0R�'\O���=)�쉗$��)f��A��t)���rcV4���m����O��4�0�Z���O���O�7MM5pU�y�C�@i���Qԍ�0.(�W����G��;�>Y��Gu4Us���%�.��R�F�s/~DI�G=�$�P���č�I#�5�f Շz��X�G�*O������K�>�S�? pܹOÿ	��{f&\{U��"O��h�0����aŕ*p��p���t���'j��L�	��0<.�C�z���v�'P�AQ�`
�12�'��'4,םΟd���(,�A�U�܉���LZ�pc i�5$�i�Y�:]�7�? ���Ζ=T�<i��7.(9����ؔ"�A-U�X]YCb^�[q`��胳~��p�;l9(����L���&�$@���Dʖ�II9�?��'$ <y�`ԃ��̣3G�8:�\���'�p�R�.> ������&�P�����e��V��W>�}"�A�yD2��Sm.v�~����'mB�'�l��'�0��=����`��IS�>(MK���;9t�B�옳J�z�Cs��iX���F��1Q��m�C�"a#�5"�]+v���Y���$r�8�1��?��<)�$ğ`;�'q��3���6���q�Ӛf�*8��'L<ڐ��B��lA��"]؈HH�'����l�z�n��1��Q�D��K�n�skTQ�i!�'.�f��u@v&�yX f�n�Ҕ��Yğd��ݟ�y�	� )D�A�
4Y�\@����	b�)�A�<&
��`������@3� ��(yA�)Q�s6�x��L3i1��iƅ�JY���O;Ig�����?���p�F��O��`��%�`��;�c��?KJ�7F����	����I��G~B�_�o ��7��*�p؀�́�p=�����"ȅy�N�;��X�f���]���P��M����?��|����?y���?�4hu�	��&�:��
�R��H��A�X����̜r}2�?��|�'�I!P��G̜h4�+_�}`Ц�5u^pz�����X���dֲQ�`�3ƆѰ�f@P�.K�ef=�ɷ��f�>����0cK�}�ε14)������LI3�J�&c�ڨ��ةv� 1�=	��)���;[� A{UM rQL!a��\�D�*��I	�� �`Uҟ���㟄����u'�'���&\x��rph�@�Y3v�V�ڑc�7(� �ǋ,�^�Jԍ��G~�dΩQ��[���Ut�AXG��k?,�c^��L,�A)��x��ܮ{�'��MX@�_��R`��Sk���4
���	��p>�"E�Dx��eK�5O�@5OD�<�S>]/�@��aB����c�B�'�c���Eƙ��M��4mcjT�U�I5�:$y򯜯|W(���'���'�@����'*�?���q
��S)�q��0� ��)�Ԁ3Յשd�������v*�WZ(! %B��j�g�2+� }����F�Ń2��I�,�F}b���?Yq�Oؐ{���\�R���G���rp�V"O�L�����Ǫ6~<�� ^��yBi��.!*-����Zr�9C�_����>y��25ě��'a"S>A��4��KR*�=$�(:0�ʵV
�`����\��& <v�jE�G�/��U��){ݽ0�o�"�\�U�^�u_~��*?�	��e)�Dź�L��)�����U�A�P!{��+�Ξ�|?V\#���ߎ��
&�Lw�T��`ѭgصkĭˏq�8��}h8��`I֟1:Xp{�iH0@(�P��I��'���� \)�Zu{ASu|�B4�8�L�$�O��$�O��
�@���O���~�Vq��̃�x��i�p�Q}6�(�@�I�|p�d��9�d-����+�Y���#cM#Ey�������}��0�G�
�SE!Űx���$H�:=�$�bd :UJ[ȟ��w�f�RK�6 A��աK(�(\�A��Ov�d¦y��K>�>�O$F���j�
��hʖ�Y����T�'��OX"?���-�B����� ��H���G`ܓa�6hgӘ�O�˧�M`��&�9�q��&+lԁڐn��EI�6P���'�b�'Nɳ~���ߩI�吭Ö�RS��<��5��O�3|�}��15�k��яJ�`֝C�'�D��PΛ]H�ձ��G2���K"LI& ���e�i{"1I槐L(뎟F�8K��D�Wz�8��;e�h	qA,J�hq��y�g������⟈��^y��'��'���vʧXȽ�-�*_���'��� EN�<%��z�	 _F0����ޢ�~bP��;&aO8�uG�ibN}�g

6)Vl����݇1��PQ#F�O���O�i�!��Op�$l>����O��I�hU@^d�рb�4����Iv�Ot���	?���Z���P*� #��'l�P���
�d�A��T����%$F`0����o�!�D�f�d㕥�� 'F�s��8�!�E$9��hY����D:�1"u�Z�A�Z�i�}�G�%5h7-�OZ���|����8Og�؊ŐZ�͢�dؘ%S������?��BX=x1"Z$2\Kgc�z��}�/�(�݇s]�=#��
%'�h�GA�.?�c�L�vM�Py�y�����8`�0񉅬�0�؄d�(#V��2�u��O�\�3�'n<�~J��u����nВP^�D��p�<� ҝ�ckP��"�[Cć"LO>��3�'(㞘�6�ѵ0��}z��ȋTn�(�ba��q���;s�i��'t�O]f�T�'���'̛f��=0q���feθC:�����Q���+P��P;8D�'���S�g}�F�OƊ:��2f ni9�I��R��'��:� �'`�#}�'���ja���Q��`�e&K�/�,��h�OH�&�0���Y���H�U/(��%�'x�8��?D� �Ѡ��.,��ZB�G�%b=J�qO� EzJ~B��=L�N���m_�'���*�E:$��/�l��qb�';��'��M�i��͟��@%0��E��#R���(�����\�Є�뒮>S��Ӣ�L�"����"�A�O�t�!XiP�cd[3([���箚�8RRAp�	&fh�=���H��(��F�{c� ��nZ�(�����ܴ��'� �Od���m�/&�X�֎�!��� �'��%���G,y��H���I(�����P}U�����	�M�޴^y��h񦍼nU.��B4bE���e�'2R�'�0J��'l"5��ysp�
+M8���!Ǟ��4č7)fr���ѠVT�E�퉟f\!�oD�'�� i��99�a�7]�4X@$h_���=��K�ǟ�`�'�@��W�z[*�D��6��i	�'*Y�X):�^�C�D�9� 8
	�'%|�s�<8h�Ə58���P"�^�M��hH��i�r�'0�S_"n\�S`�:���+I�AC�������b�Tɟt�<��?	3��6��6+�9��i#!E�"�ExJ|�PJ��o��P�,&�}��$D�[�=��T�O�ȼk��2W�;%]�*H ���'qv}��#�	�:�����$:���
�1qOȴa ]�m}�,�E�!wJ&�ё������4�?����?ͧB	��?���M���ATg&is�%̻P�����b�D _F{r	ըY�Tz�(Ƽs5��9��B$��#<���>���FF������9(�p �NM2�-��W���d8Bd�A�gգ"5�!�M/�!�.��P�CI����֫B1z�qO*�DzJ~��`��#(&�ct�v=�l��_1;Db�՞P�d�g�'���'f2'b������9/SR���/�4K �·��;����,k4�wM��u��z���?@�:�!,1�N!x(��MsU���{��Ċa2�p=	�m�e3 HC#�WhdLQ�
ᦁQ��O��4�D�O���7�D�WB ��h̸,'d�kWÅ	oh!�dZx��FI��:����wQ�Ps�O�˓$�,����i�&��Q�U�1�ݾ@�m1���7c����O���	>$���O��S*3'~�#3$Z#Y�d9q&�S�	8�11�B�Nq:�x��c��I��	�~���DY�I�s�M=�$�:�<w���	�HC3_^H��k����Oⱳ��'r�iڌ�
$o[SV���F&E$,�fl�J�4��ʟ��?%?��Fą
),(�G��x����%�'D�daQ�T�B!��+�G&�p�@�I?���Qyүյ���'l�]>��w�ݑ+�����V�&�F�>\K�-�Iɟ��	�Y6D��X����.y��OJ�nŬ�&�A�_��9���Z0r4�Ov��U
Q��x���Թn�[%NËZ��Q8b
"C�N���'��+i�]�/M�M�p�{�̉�?���+'���'���)�2Պ,_�T���Y�d�Q6RQ�Ū�O��O\��<�b*�*2���$�1i!�9W%�Q��(�۴N��'�(�D�>&G�#���12�N�"��N}���E~Ӛ���O��꟒�;���O����O�6kwx}����ډ��i�2IP��5�Sz4��%J���O1��I&\*��K���]�V�Q+�x*����$�15�0��婉oو���>h*�-b��Y�)Oͼ��l�l��%�v����pDz�a�m��'��'t�D��O �I��x�*���@��%y�?���+�O*���˅P��Q�`ʗRWR��V�'M��ۦ�qI�) ��p�'.%��i�+I��?�b`�-�D����?q��?Q`�����Og��Y�lۤ=n,��!�V�Mc�m��m�R�!�{���׊|��  �T
"��ulZ�,��Z�+G8�X8u��
Y@x�"܈Hoh�b&dc� )��'�\��$,?���)w��~Ŏ8+���)<�!��;q��s��N�f�c��9�Q�tb�}���x�7mg�&" �,{b��)Ej�2'�Dhah�l��ݟ�[��Ɵ����|�스E%2�(3N��l �z$A�k�
���ȌI�@��e�-p`��ۍ���?W&-36�� C�9 ��)n�K�f;{瘘(�ؠS�x1�`!�>���I��~R!�8	�� A%D��q$�Q��*�y�䉒R�(��G��l4�PI%���y
� ����&H�|Eq+�)_�&�g���'	����et�����O��'6gb�*�� dk~43Si�0kڹX1n�-�?��?1�E��'�~]t��U
��B#o­St������g�F�&$��(�n��M[�x�`PC`R�Jn���㚡Jx�N?���KBz�0ا��U��鐭*���+~2��o�Oo@J1N
�p�܋4�R�W�����'�Z���f �fd�5Q�I�m1ד|�qO�K�Qq"��@)ӫ@��� ���g��8�4�?���?�'gZp����?Y���M���*��-�M!y��q���O�lA��M֊q���ۄm�Oн�'ژ�������E^�}�\��C�6��Y���	5:�ٖ̈  ��}�I��H��ɪ[�q*#��\���My�B������'�J"}�'hr�y0���y+[>��Z�'B��E��oU�y�dF5�(��{R�2�S�= �~h�Oľ�0��d,�Gi��K�=�Y�ՌN��?���?Q������.@�g���ل5`����.��|��֨��3�l"C@«?�5r��9O|�b�R�Iӄ�a��	n�)w�i���so^$c�i����\���Vn��4���<�P;�$]q���(q��ן0��4E�V�'?�	ş $�<kf+J�e�|h� ����m4D���Fĭ:�����ÌO[�	�2�?�	Cy"�8L|6�f�$t�լ��t��Wđ���2H��`�IğH�K�쟠�	�|��B�a�X\;qNƾ`����%�]0R%8�� 5\�"�ð�^b�� ��.w� �Y���O�i1�/��P�³`�'՚�r��0� �
�6nvPXA�7�	7
n~��N?Q�K�,^���R��#��yHbH�R�<ɵ�Ӡ,����b�cHxТc�D�<���l�<B
t�Dj���//"6�!��ܓ-^J@l���T�	a�4��5���I�)N�c?�ԛ��E {�� 0�'���'�Ҹ��� �2Y@��P_$:�I�~�]wh���E'�vĴ���<��%��}�0H	<90��[�n*�D#A� ����%2!g�Ѿ��U���kJ���>Yf�ӟt���)��BnJ�&}� #�	�Y="���"O��"��b����LT�-�Rxi2�'�XX�ꍋD-�|�tKL�Vv��
�%���"~�	�j2�<��G��1�dQ���~��C�I�X(�z��:b�q���nC���5`�+`�~���њ@�N���D�z�'�8�3� �!^I�%�&B�����'`��{6��sT=�i�9w���'�3ѠK-e�����ȇ0��y�
�'�y���j��A�Ae�"P��Aq
�'��XB�H#YP�$G��TrL	�	�'T��Pr*T%\��)T�^MZ!��'S<KW�. |9�+ǻtdJl��'�܉KCfTحY]���
�'�b�)G������$ьE3����'����P � UH��b�1#����'����r��W.���@C�.���'(�`�B�2���Y7b�69j���'��Ђ�FؽZ!����"��
�'���GK�&pO>���Iތ.���	�'S^�áJÙ~`tB���m=���'cV�`nK5�P$h2�ĩ]ޢ���'U\�	�.ԥ{)Hea��F?R��ih�'���`B�Í\�L�'�g��s�'߬}�#a�;T�{�2\����'�ΥHP��5���3�� Z���*�'��g �$ixES�G�(L��'r6����1����t�X�:�����'�d�bg�jD>���^3 �I�'P�
��(���䗟޼��'�p𑗎�2olm�W)�7	�X�3�'��I��m��A��-p�}=p�+�'O��@����*��i�G�Q�I3�'�>�3��J0mȭ����~(����'�><Ӧ��s%��j�l����
�'�����.2Qf��RԳ_���
�'��9�b�-s�,K��ۻLf���	�'��j���8C".�xS��>�l����� J q��0i����D3}M�-ˡ"O�]a�bB�%����*;�`�� "OjXb���r��Ȍ���(�0"O����8!ڥ�FGU*���%"O�� ���e��P� 6@�p���yrGT<+��pE!�6�p0�ף��yb��!T$�ZRxy��ۓqnC��'S�%�s	N01����D/7?C0B�9{�Re:��$4�2a�c�D��ĊD�$�vB�9��C6d"��PBR(�!�D��7������ ���`D�<��O� �g�j�O8x��v,����J�6���'�pf ��
�p�@Q 1Dn�*��d"c��
��Y�<����nh�y(F���|���rH�^��a��)0�PJ�g�>��5s2O�xs ��P�U]�8nڲeG��
r/.\O�9���|�BT;���4�½сf�% 3����̈́4 �#?�u�̍22 	�'���Ȥ�C�p$u�F��1	69��$Ǧ/@�SIC�7���OQ��a'd� '�Z쀔�/��(�}ң
{!DQQ����Q*ԲG�]����CKӐ'��	=P�B���Fߚ_�� 1ç"i&�3�nO�H��bs]�.GVZ<�Y�'����P��~�C� ��a�6�'�4��$'O�2�h�O�,�����)����}b��6Vb��c� ,��Q��y2&Ш?!��ف�BB�'W3wm��[A���cF#Pz�	sj"?�y���]�<tay2F1Au2H��I�'þ��fV�5�V(�Qh�5@
l�'����+ؙl'�� &�~�7�^
WA����ȜK�����Fy2��,,��(�D�X�O�v�[�-\�^�xk"�_�`x��O޴����L4��D��|>���9<]
��GYL�4)闂��r�蠛s��S�ӧ���c^1���j�ª/th�����8��'��đ�ĂE�Z��OD%Y�&:eXIЦU�H���� �O�5�2 �3��X���$�&��\�RFӵx�8�H.U�h�P�+��*`<U�	ϓT�|� �kX�/g:���,0}5��J5���K,���6O��eժx�֓O���Aɿu,�8��#�H�<� �ɡ��ܲ1�	>w.>1s6|JvI�Lz���3�4D�,9�Ȃ�q��l�t�V��EI��q�Up ��O�j�O?7�ܠ8��:�di�vX���wz!��D�D"#F�;]Μ��F�}e!�[�]�4�5O1+��2G�Vf!��NW��i�"f7K�:u"�[(Pk!�@�6�����p(F��5\�!�NF�Pd���C�6��\ ^_!�X�YT�@ A�k����D 2�!��M�?�"x�ËB��ʑ1T�ߗCi!�$O�*�(����<� c� V�!�dU>D���m�
d�<�8$���a~b ��h���0��@�(Đ�i���6H�
��F�/f����{ =��G/c�f:C�K�!t�F{ҋބB����kX��1����97lv\U�S0U,5*�"OnRl 6<���4"��~8� �Ʋi+�0�fz�HX��O^?E�ܴ� �R��� ���!��O-~ʰ�2��ٖ�(��Ix�X�U Y��ܹ��>Qϔ������ϯa�J�$&�	�$�3)�(Lri 8��A��+��8�6��$M�;��q�@�� )�X�H���'f����	�>>t�l����O��������� M���!��^��D��:Q�#=�b� $q��8���������W�8^en��%�I�쩒���L�����{��4oX�d)�A��wq�)����>�M{��E=.ND��5���Fr�)��5q�D�!����TI�7]�� �NԑTNqO�tS��3?"K	Ard�d�3uo�/���y2GAlAwfE��H��D�h�� aG�����`D�&��5��iK�p<���z�Jz��ƶ�o��!�r�(�+G%2���[�n�T��D��_:.O@Ҕ��,r�؃)��R8�0�r�	[ިZ)�[6�'3�
V7�9;��Y*jE���	�&YJ��DS�nL��XѺive�󡎝G�ze��T4y�����:��)�
�6QJZ��S7���	3h}`����a:<Mh��im�#<Y 퍴g���8�W�Ou(�q���	�XPcL�QPz��B6{$ �@k&5�(��)� �yk�
R�:t0\PG儌?���si]7g�(%���tVL����i誔��ǒ�qz8���U.P���� Ͼ�����!B�FB�	Dl��xrD�n*��a+Ѹ6�>6�K�\����#5`-�f���p��$���!KQ8��)��F/ȝ����hC�8�šAb��zrc�1xiP aت����ǠJk����yfF�c0 ?~x��Ƙ�c��Ƀ:������#�5x`X���Ao�i�1�	l�}!aoM1E�w&��h�q��偗&���"�Ʉ4|ΌKŁڞx�dPH�i�p�HL��Ij#��FS�5���c@���*;4L��b`&m h
�N}���#��F�~
��EG�?�S�̶@
D}C��D�0���*B��K�<9e��2��e���YYHF����R�9+1�޴Jd�-�eD��P�mx�Λ���$�T�N5�1���O$Cʪ���ɝ>�����'ˮ�ِ≟;���{$`@�x��}C3.7,�92ba�6:<��֯Z�3�:Y���<���>i�ք�|�' |��1)�1
@�2�*Z0v��J>9�	8d��� ���<��D.r��Ot�+�Ḙ!��Ԩ6�G;� �a۴wಠ�������$���؆ �z�"᪂�@:S�BMz @��jԱ�w�R/+�
�5��d��%YY�!8G��Ꟍ��E�-^�9%�9V�e��+4�%_�F����7i\�쁇Ǘ�s��=����3��H�E	}sz�P�)Y�B4�O��b!�8�Z���t�t�kb@qXp&�Bmx��{R���rL\y�C. Q>�(#�¸s�2�JW�G�t�І-3P$��QG]���I'[c�T���O�)rp�wl����@zF�E�G�ĀxC�e���Z���)gF.�1�����8۞����%�9��'��Ȣ�MI��a|2��-a�Hx��"3����a�kUr���	S��1�l�>2��N|RD��44|(M�Oظ	 �L>�f��7�&>Y:%5"O\=����8%� x��eFܼ=���U39�P�k�	��;S��@ԍ!\bJ��K%}�(�6F��I�'�8��-ށ{bH�#%�l�zb�^P�D{��>V��Z�MZk������2}�P
RF�7׾��&����	�$h�M��'��0CS��(:��2�	C�$U��}r�;K�"mk���E�V�U����S�f�he�~Dٹ�iW��17IS�
�n����M�����ʕ?����qIF*]��tɔM�b}�L�s��h}J~���ԏM>J����OFx�eD�3��A�´>.�B"ON)�Gუ7�������%6崉��;O<<j���9Z�zUz���(�Z	��#}҆<���܎Q 
�I��<H �3�
eX��3w�	�J�z7-*� �qEW��>�I���"0��y����Uv�'aR#}�'0�yA��L�R�g[�^zB�
aL�<	e��=b� `�J\e�J�ß�3F�B�,��1��	�H�z���W2M@�QP�F ?,���27���'��Y@������+��|q��2�^R���M>� �t��۵7��p����a�<!��M{�T��'�3\� 8檅Y�I�1[�<����I�TDZ�	M>uE��R+X�I�}�4[#�'�~�r�B��i�pM���hJ�'�	 Kf*�
@I$#�v�z����N4�i�%�)����,����x��U?%#��Rd�(&[H}�a�^=N�V�+�"�m̓N�\���O�G4��?��B-��6���"[p-�E�?<O0������MO(�Z�hMOZ���3-��h���o�Q�
�9@I��sv�S��M[��\u��p�O�2M��y���Vx�2O��e����I?DǊq�'�N�|0��M��G��	�=�@�%��7o8�yү�09ν2�	A#ShhSFn��&��O�!���	�3q��w��T�%�
�4R�Ѐ5��($MB-P�'/V<�e�D��I"T(N�x�"���V8!+Yx4�
�fM�ě1E>�Jy�D އ�y� R9?��Р"�W8Z��4��M;�ǘ^��:K:}���i��L)�)�!m�H�e�ʃ0�\�s�'Xt�{"�j��$k�$π`��%��O�]��ę�$��!vh\8V)� 
R��B��@Xȅ�ɭA\�9"ǆ�iI����¢O�-�ō�".hH��L4���$��$Bv�j��Y�`�uE|�Ɇ�Z� �D���&��s%GY�A4c��E��y D'UU��	�&AK Yq����y�.�'vyj��àu��h3�c�(�y�K�Xjf(z��4X��mŪJ7�y�J� �R|K���^�2��Õ��y��H�(R�4��H=%��y®\�v�xɆlۺ����i���y
� ,I���59HiVA�.xe~L"5"O�T�󇗪&�����
W8���"O�ic񩉔����4�2��b"O�d`��1UF��k؏�*$�!"Oj��O�8�(��uK+w�����"O�A24��=�s@j�M��-R�"O�%���T��m	g���M�>Y*'"O���V,�.%�8 X�My`<h2"O� �E�ѻ)v�)t	�u��"O�$��� �^aR4�]h�"OЁ��Y��	�v��~M�[q"O<�h�ש �[N�"�� "Op�AC�	����P�S�d��j"O� Z��˼y�n����'@8$[Q"O>�K��J;�h�1�Oj$�0&"O��Je��.)%���B$KI^@�"On̢�&T��=��$�$+&��"O&@�h�_b��;�HF1� +!"O\|�����fV�s��-�C"O�X�Q�2�k�l�}+44b�"OrY!�e�&9�}[뜋)�My�"O���C�L�]�:�B�+ɧJ���
t"O����(L(H-1�׾�0�;r"O�5k�'��,���R3�� W֠L��"Ohm��+߳}@���t�G|&���4"O.��Sfʖ-�t� �H�Mz9S"O�=��GA1?#����7=lx0"�"O���Ժs'��Sঅp�����"OM#�a	�E��#�t�|�`"O�d!�Rz�����- *l��jT"OP�q���	m��%�pJL~�MA�"O�ɕ�ĸ#�>h�r޾~3���"O
�8�ĚJ�%��EF�ZJ@�"O�q���^�H�IPe�"oDl�s"O\A�r�'^B��ɦO�S�tu�c"Oٚ�� ��u��d�S�y�uQ.���p�Ο$mC�@��X�Y��?�6��H2���ׅ0��4�mj�<�� rҤ̑�Iɭ����bMJd�<�𢍜P��E�+R�h�r�^�<��A �"�:tb�bRʐ�J�K\�<�4$ɮ����a��.� Ԓ�GKY�<���D�)zqA�3�ً6��V�<�D��w�P���U�nBX3TH	h�<�-ׇ9a����,��X?�Y��N�n�<)�Ô,jbU{$W%_d8��Q�<Aa�P�3Y�q�� %��F�I�<j��FiY�<6RR��MC�<���>o���)��9t1h��V�C�<�AL��I��0�F��M�YQ2��X�<���ԆKG<��E�M2��`��l�<	�@����s����^.Q�L�f�<�!�ǦV>L	�)�7r#j�����Y�<1u��yɠ vF�.`���2�M�<b��#���A6~����+�T�<��\|
���ŏ47$�#oHP�<��]0�:�4&D._$��m�f�<q�r�&}��֬:H��{�L�<�%ۙ e��cԨ��p��}�e�[F�<����=�MHRG�
@Q��᠅�<��B�"Gv�+
#���M�o�<!D���l�L����2<����dv�<��!P�T&�E�~���G�K�<��A�J���)p�σn�0��RE�<�Q3.����`;\�z��!�[@�'�|1h���K��4� �lz5X,e����b��mr�Ѧކ3�ʓ%�~����?���~ʡT�����F"&ꂝa�A��K��������$`�&�9v��'-n�)�',ޮ�)ڥhL����'*W�!'�d��Ԯ�A��˵]0D���?�'�hcqD�1g�y���F�o|���'��	���d!-���Ӻ�睏:���J%zI�=�Ҏ�0h���-B4:L�U���3km�	�&�OQўD���oZ���pr�D
`|������.!��D�.gWJ��'溅l�F�''xU��.�8Ѷ����]�uc����)U�	�!^�-��xΓ)]�D�y:`���Dσ G��bb@�%���/��O:�Ϝ6S�:,�!F��赡AC�a��ŉ5��L�ް��Z�D\�I���� ��O货O��vV��D-R�r���['(�C3bK�D��OЍ�!]4Hp�abޛ.���$�x'W�6z\��@S�S?�తͼK�r4�e��e�dY��(O���t���eƿJ#�	J�O
NTL��D�:i�f��0j��D|ԡ���O�L��z[�i{g�=H��C�+��Ұ���)��<�CkJ6e�} ��^�y#nd+Qh.y4Q�଻i�ؕ�	Ԧ;�挺��T��~BBߌ	%�\�!oԳ$t\�����yR*�%��O�$���d��"�g�$Z���Z(@�#,f̴�#`TꟀ����z���`e�\�z�F�`�8}B�����s�V����C�z /�3�*Y�<y'�s@*X:gU�~�l2�H��?�'������X� "`D0Iښ�hI�1BKI��t�Od�Ҕc�v��|���j�U��)�1%�fhr�J
@�*���@@�bQ�g֠f������*��;��1;���5����	נDZPɓp/�����t
�e�'k���<�Z�萭��fz)��N.ʓ�u�\ :��i�S�
����OJ`:KA't�rԨ
*b����<O�1�GP�(O�rР
"�����C1x�D 0:�Ā� �>Rf�
��'�p��CP,x�R�!hF� �x�H����"�ny��1X�����^�2`|"�-C��'�`}"�%S�'��Q$�1��4��g��O\oj���Jw^����O�0��u�񮖰8����)ht��?��oZz\潂�ǐSR��a���,<�&Ԣ�m��p;!M=v������dR~T��x��?!J��J�."*���Gk��w̐�Q�Ov�g� ����
�b��ya"�&l�@�I�e�.&��F}b��S��I�������`���" ����ο.���d+#^�,�<O����ɛ_ld`��ơE� e�Ǿ,-���k0<�e{$5F<ʓMH�}1��,\h�'[�s°������[��X�Lچn�0�%k�,�ذg2�	2D,�ڴo�UO�l� � 2� �M<�q�ݶ~�5 �J��rQ�+Ӡ]o�l��	O�	Av�P,N	bDX0�>��O8$�iq�L�3 F/_��`��6�2 ȡJ�z�`�p�^ x���h'!`��[���+�p3�\�96��%#ڢ'��9��<��N��(�с��X�'�D\��c�6��)�㦀#�X�z�� Q޴BDMzgm�QW`��P�Q����]� =$�H��-O�@��*�a0�d	�K�tz����B�yZ��E�Q	sÍ6��'
B��;���E ��U��P>˓5O�F�֜~pY���īD���=�S�E�X�{&'b5�e��"�	�YxfA�r�ќ=Wԑ!uF��ް��o�i'��wMy��D��,CN���Ɇ�<�R�h2+Z$L2�3�L�)l9�G���6�@G�x8��'\��i(B�M����#����L0��m�N��W.�-n��b�n�UJ�x�jO�7������T(��LK�fSdyeH"OX�h�"o3Ұh2M&�I:��&8���`�U j^f���zzҔ#d-�G�\�sj�2}���O�0��%z.��WG_�2�D���dE�V�U$��
��8@�Rݛ֢��
�ļ�S	�]�(=�G�˪�����۠�v\�WhټziH��Ņhɾ($`ץ>�̩��$��?���O�
��E!/��u���oӴ�)�/H�L���I���=Ie��7�TibVB��W�i�@w�â����;?��T��	�
@��x��S�GP���r�X�Aڌ@�'�}�'�=��D��SE�D
�n�a�<�ڴu��Z�,��<H��Eo�X�	Ky"�_i0���S�<o���~, �a2�E�bƠz��U-F02��U�R���+e.j0����0H.�8ԧRB�PO�c��aC� &G���p�L�Xn29�W�8�L�æA�a.�c�"\�I�
��D���ԚE��`��������0F�0kԡY�Ԋ�'��O���I+�?��
2�eyǥ�K��H�B@�!A�zY@��J�3��b�$m�tে%�(O���Z�s�р�H��J^dM�"��K�h�4Z0�sR���i�ĵ��'����s�� �
J�� H�Re�;�Ҁ����+-��<�S�Bw I�Vm�]7ҁ���a�aAS�ȺU-� �çM�̨�E��<U��t� ]��ύ�_�`%�\��ǝ�LaCW��?��%��qy�%c�OצN:8��4hql���%	�=:6t�Łο*
r�"sdL� ��{]̪(�1P=��7$ʖ{JLH(`®>��9'�H*hҎ~�8�K��=âm���4?)@�Y� 8�1�G���m;,�#�΁B��T	��|r�σF��tIK�{<�X�N~�㔺M�,� ,��(ۂOl�N����ЂL@�h��i��m8�u�=��yW���"<���)6o�T���DF�#պ�jB�K/�RA��K�G��O�>������2Eڝ�������."���5�DO7�����iR�e�۴Y�ʓ ���2ň��Th�T�rd׍�lJ�'�H�
�O+Of��`�����k�f��d�ф@��� L��ef�9,G 0P��(
�,�k���憜�v#UOp�����
N3<�)���1�$`d�0A
^U=��*'':k̓O��(#/Y��@ B3T ��Rћ� �j��l?�-�5L�j�R�9�%}�!�b��h7���L[��S��\�#���>�-{��«m2���5~r�)�W���O*��i�����9�~@��C�T�d5����F��"��&�(DKW�l�+ !j���S�8db>�D�+}�A��( aҝCS'�2f�4�����	�|"!҃@��������k�t�(���z4b/W��A��'>�I�p�VbybT3$��"�bU1 6o �4�0�У"���'��m7x�	 B��<(�!�0���r�G{?�w�x�F�Dx0t���ѡL����FK����bΑ#.�و��H<��c��؊��X2�b��Ki���'Z�p ���c�8��J+ 9�툭O�O���!�%T��P{6.��kF�Sm�8�
�AS
Z0F�^�&�����S�E2���!T��jf�^,~1:��?��o�:A�3�/&^L�%D, �!�)�� ���YJ4<�V�@�7�f���?��Jf �b0ߌe;f�"0+�=�8��?1�O�#=���&2�Jy�BQ$'�0qpbn��y⪕%&e2B#�v��L>1F%cnv����1c�H��GB�y��ź�iW��8���$U���	��$̨ċ�6#�֕ӂ%�,����ѹ>k�u��c��"P�b�|�k��b��f%�+!?��NK��AI:v��t��CdVa˒K��qO0eˡJ�5g�i�7�����8b3
�O�|2�(�]p���"�4:f���ɉ�b�����k� �C�k�)[�	)`�����\�M[�(�kB��7+�o-Nxk�턫uFB=��,ݜ{2-�T捥R�θ��C�v�]>7m��t�4�g鋜3��H�pjH0qla�vKþ1�On��7y�T,�Y�H�Pt{"�Oxf65��/R�E�DС�M�G2|u�ab[�{��Y�O�<y �G�?��#J�%y�Ѣ�]c���c�C�1W�D :� N�OPH�I&�tq�B�s��5����Ā�7“j�Q�G�X(F*��9���h��2��K�5���y�h�����(�`�K#JJ��;��?�
Ɠ��s/v�0�q)�Km��xu ��@��',�����LB����-	�l\���9���@h��h	>z��͏4-X�x���V��/��-P�I���4�Z睵=$]X��P	��L١�� TRX�gH�O
���~�O�V閧���u�� R�6
M�r���1��hO�y��TB��@W�L�<���O ���� 4'�*4	�Z� ��>OAq�X���$�<��y� �(TP6��xc�Spٰ��%{���h�A�-�?cɁ-k��Q�Áɮf�4��Ca�T>���)&��q���j,����	�l�DyRk��&��J��֡T����@͙���'z@�RaM�[�<X3�ߜci�MȠ�O��?9��*�),4���˜.R���;�%ϊv�8���Jï<?�� � H��Q��jc�C˼d^�>�8!Ί���Й���B}@�i8��iE�[昘�ɛ�'����W��hO����͆f��@�b�Y!�?-�~��z�t��`�W�� ��?԰<�Eюa.>j#H�?(��`WR�55a�7.�%�X�Q��.Rk9c9�Uʚ[UJQ�I���'�.A�	�rV
��CNGHY+��	DO���R�O�)c� �Z�Ta�}"+Se��U `f��B[D�l�822�S" Kex��.�8QlD�"�4<�v��*��y�V�l�RL�W�ɀ��9�<*�uPSL�$���kV�Șw�����z��Ӥ��qo��#IՑN-d��P&�_H�q�s[UF�������4�������`�������]�<E許6�1[�!9�,�щ'��Av(I���I��=uV����}���-`F�m����f�(��"�[���	�gL�Pz5M�� Ӵ�Ę�M?t�T>�	�Dh�!GW��������� H��
02tp4{T�ɹ۰=ɤN�b�D�R������j�l#D�>���:��<�O[�t�s��	j�v���m�6)��h�'�'Z��Ѧ���|�����^?��8�M���d�6Nla��뻟�@��3V����5�|�Rk 1���o�{Vq���Wm�'�|ԸVcS����g�6F�Vp���|�ť�=���El�������H��jA��b��Dfy	��ȈU�|�<�^�@�FzT5�\���V�kP�	 `Ԁ7@@T�d�%|�n��S�Ͽ��F�`��\Pdˈja��Ӊ
|�$`	�A�%����{��9��%l� �&�ſO}��3��ֱ3I�Y�	�+2X���O�:j�B��?�r�=�9ɱDW�6�`�!aG#�O�݁E��=MC��rF��B�J9\^�p�F�p�buN��B�Z�^�r�F2Q*p�`ɟ���tbC�u���9�`�CFD�(�#�HO:�)ʚ_h4�ԁA�"K�ɡ?��A)��"�<4h����KP ʈ_h+�S�6�H�I�B�Q>˓ �j������ۮ���'��?��q�O�\�Ջ_:9��@��#�P,^����[��B,�waW�&����hظ4�c#�=�v$�鉤:����p�V>d�r���	�JH�W����$��S�v��禝p��/Y8\�̛s^5����܌lrJ�"OHI9c(:���[�ˊ6vp���a�'F�����E:�ia�ܿY�HH;�O��b?���Lzg��P����Ղ�q�5�O�����<Y)B�?��@��Ł(o"<��\�e"%�W��,tN\��.ң.��t&?�@´�	�e����5FuAQ�0�O@���9� �Y��N�:��b�3xZ���-��j�������&8��I*��p�cA+A/t	 ���C8��?Q��%q,��,��/J�RR�z�]B$�G�o>�� ��@4���S9D�8�	�g��#r&�+lg�����<qg�ع/����?D�B}���)ҧo�<� �W�3���bF��p����ȓz���*�Oq�9���?y0t���X�Y*B(��n��Kx�g��0EZ@ρ-��E �#7-���"��qF.�)}�`,y��9;�"7D��y��:,�2��b��3!4\� �:D�DJS.[����.@�nO �`�D3D�`��O10�q`�9�zU�$D�XR��&��̻����g���qҫ/D�L"�-�I�8�����q��%���;D��qEm�4z�*�D�� ����>D�X3R�C�[��;3k^h�h��"A;D�\k���m�N}���>A`R�L.D��r�̻a(x�!��;e��as�&D����ЧV*�����8-�Q��$D����m]�p8@i�1��)*Vh!D�Ă%DʰyTY��	?>*��A&)>D�XR�B�*o��骰�=`N�d�#�9D��
߼p���	�������8D����,A�)z�gf��$5D�X:��ŏd>q�⋍$X�� ��'D�P� �6���غ+�th��&D���GH�b6>P����
	�s@&D�l��M��?�d��@I6k丄�U�0D�X�`R,C�x��ۋ_>���(D�آ�O�Y�^�2�,&^"i�4M%D��� D$F�U3����[�
)�@$D�\�&A�=w�p�"�^�\;���c$'D���ё%������[$BOf� cf&D� ��.��m���d"*�z�H �%D���!�@�SbP;�dY�
>����%'D�HZB���%C���["��9Ш�	�'`���H,^R�9S*'X�,@�'Q
M�B
�v�����J��M>��
�'
� �ŀ�"�PT����IN�1
�'\�} 3hW���<�Ԧ�t�J
�'�R�����
Dx�Y�d�	jiS
�'�*= o��M�p%s���i̴�	�'g�%Y�Ĉ;΄M1DkRn����'�J�Z �3t� ���V%a�j�S�'9�#v,>�8@��ױpP  a
�'��p����F>�X�1��jg��X
�'�	�T'��v�s���j|A
�'�ruy�)ǯ+��Y  �a
�'$-:���w���B�����]��'��I�9��!x5�ʗ1�N���'�aҳ�~�1cD�[�\9	�'�r�xG��A��@2��Q5A�t�'� p2�B<�J���N�4�b�'/���M�PQn���oݱf�c�'���4@�$���%M�0r�Z��'�(���B�5u���ū��mbV�Y�'X �*��� A��	:*¢M��y�'����D��?��85	�>iVl��'l�|���0���d�P.�"�H�'f|q�5��</5^��Q@\>-�h]�'�����A��a̎�ro�!��)�'b�4�F)�=T�ܹ�LUju�#�'�\�;�����3AE@_����	�'*���0���f�D�	�ɋ�^i i��'���`$"|��l�R��`���� ��y���TNz���;���jf"O�1�(�4� ��Q޸a�P"O(�s��ϳT;�ՐB�P�I)��S�"O�E ꉃ7��Ba�#VdBF"O�Ip�oʚ���� ��=�(ju"O��1��[t��+!��]|8�p&"O��� ң�D񩰍��`��ZB"O$LIf���<T��0L��Bez�"O��S��M�8Y��`�w�e�`"O�[Eb�?yrT�BJ�F�� ��"O`�AFs�|���R�S�V�0�"Oܽ@�b(+ƨQa���hur�@"O0 1���z��ݲb��"d2�"O�ـ@� v����,�MRݙ�"O`D�)X�wp<��6�ؘdH|Y�"O؜k%�9�"9H��X�'�����"Ot@�m�H�v]�h*�L��"O ���$�>?��h��ä��)��"O� �'�G�.����ǘ[�vmX�"Or�ەD�&��JVł6CD��أ"O�<c�� ��\P%e#X+hX1"O��B�ȯ��G���w-^H��"O�Uj,wIp��B�0N,�p�V��y��>S0�t��B��� ��@��yb(�^w���DFDE�� �:�y�+��{������Dd*�Ц��,�y��IS�f�c5l�>r�+6�T��y�#�Cq��Ԭ��Eu~Y��MB��y2��F+��Ejɪ8/�|!�m��yBdV$H̸l)H�(/�1�!E���y��%NЂEr�$���
�'�1�yB�������f�	f�\Ea���y�O�l�4�SŒ�OZ�aPa�H��y��+�B�!�Ƃ:y����6�yr�C�W�,����s~��bw�ر�y2�
5U.��*��
��ac�@^�y��цHɃ(^��"|85Ȑ��y�'w�j1zp�!���AŎ��y���Let�;b��^�zds�-L�y�M�#��8�P9^� 1� ��y"��[�,aB�gG$L X��%���yңJ
K�nk%@�J0�@�3�'�yB�B2cM�L�)^;�;@k��y�N�/jJ�� /S�Њ��y�8 8a���0&~�%�sᐜ�y��)[��{��� �� p+\�y�:6���5��(�y����y����l�W��)GzL�V	��yr+�
D$�ݨ��^��̃��Q�y��]�k��th�&[3s������y"��"Rjd���^R8�#	��y��	�����P�L�Q`R$����y��%mc�-y`���^��)�
�y��'W)���t�Ĭ�N� n҇�yB� 
b�����U�)��ʓ�y��C	R��	��E�|���
w��y�� #����X!&�x��ƀR�y��M̎t��B'����T��y�mؔlz2��M��T����c���y���j�"p���#�N��r�3�y�`N+D:D9��Q�@�a2�^#�y�[����g$Y�N l�� hJ)�y�/�L9#�B�@f�ts��Ⱦ�y��Ǯ*��+b%�9@�X�R #�y
� 8��a���z<P9�A���`�L[�"O�I��g�$��]��(?G��u��"Od���!#�����";Bd���'�Yf&�-���rE��l���'�<("�H�q�i���GKE�<Q`�5Y��1��'�H�ab��X�<��Y�"����͈�b�w�L_�<�R������?��x1�E
]{!�D m�)�Ni� 1Ո��md!��
Z}C�OD�Z�+2n��@\!򄉦~V|��BK�R�5B���yF!�۹z���q�Ê9\�*ͫVkɝq7!�X��A�M����7 =5!򤚧�ȑ1��kF4�{�/�) �!� ���¥"�����M_S�!�U#jf��X�O�:/fv��-%E�!�'|����1��68G|�#�V�Z�!���Ag %��H2�5��ʎ�?�!�N�)!^y��bןS%�a�R
v�!��V4��:@_#c����9e�!�#� m�2"��lHܠ�%+���!�D��24	�e��*�H���L�!��Evl�q�̨.
h(T)�/u��D�[��h���Y�̗�@z�%�
�%-���yB�X��hIU�ۧCcp| �KG��yr��8�E3CF#�z�a�O_�y�"����(ҁ���S��T�yrG�?�Ģ������l����
�y�Cޘ'W�I%f��	J�hy��R��yr��{�j1ڤ�Ȼ5S��t	O��yRf�,9��r�D=|'�1��^�y� �	��H7G�pA�A��E�;�y2��.�fI0���l*ʐBU���y��B;<Q}��L�[�B5�D�:�yRE�+m;4��A�F�(r���d�<�y�mW>v�T�A/�2Oͦ���G_&�y�'B�i�� B�0J�V�{�ؓ�yR@�+"����(SY�����α�y�n�Uؘ ` �MG,��0�y��Tz��K���:H�`���yb<>B�����-#�La�Θ��y"'΢	|8-��(�d�:兗��y� PIK���WTq�nW,�y��,`�V�[�#���	 ����yD�;o����/ŋui��yb�y�H\HƆ֌w�xH�t��'�y��o�h�j���s�\��!�3�y��/G����o�\�C	]�yb��)	���iVJ�qm��z�Ç��y��׮>�8�$MĈj�Lxq0�O
�y�Y]|����[�H�Aᄪ�yb��0<W�4�#U�W6]��ˌ�y�+]�5���F��	O���҇m���y��ЇK�`]-�?{����	�y�IP*~}� �f.wغ�!��ώ�y"�F	 �ti�DD��i���!��U��yb�A�W7�5;����`ܴ�Q��y"�ь-�rL��`��x�@���˦�y��\�s��)��P�y��e�����y�d�.9δIH���4fr0X`�"�y��0Q���b�"m�W%�)�yG6+m�y([�c&\˲��'��8��O���K��ȂSή�R�'�2H���&�r�YTf��8) ��� ʥ�P@O�{��������0�T"Oz���	4�f�b�Zw�R��"O^�iA
�!vmaeP=%ق܋�"O��!�D� 4�A� *����"O��Kwa�^N�Yb#��t"F��"O���眝����/���"O (1GKKJ�șH�B�2C pȃ"Oq�mW9d��qcF�K�F�ȅ"O�X!r&Ñ;_��!愂2{� 6"O�$�&��ir�fEO��>lz�"OH1ьS"�P}��dX,8��8�"O��9	��s.�Yz���W����"O�yj��� Lд��	?d�ҝ�F"O�ѠQ�jb��pW)'��d�"OFs��S���ɴ��=�����"O"���@�%|T�����44��)z�"OvxÃ�ق=�� 0��m�lCc"Of�i�����I�
�!�L�Q"O�-`�*Ȯ�V\�)Tt���"O�y(��K�jt* #3뜤M28�+5"O�\�fh�
|�����'��O���p"O �`Q��hqj$	�YP�;�"Oz�*5�1'I:s��)I�m��"O�XV�G�.b 3�燢LB}�"O�E VK�X� �"�$XN<TE�A"OLA�F	�T�s2��-k-x�$"O2A9Q( WGf�K�K�H!e"O�1��i(��J(f��ݛ%"O�ѫB��=�k�,HB�a5"Oj<[�gI&N�.E��,�
܊���"O�ij���Xa�*�_��Q�Q"OE���B�,�Hh�l�����y�Օk'�B���'�@�8ŧ�yr(�+c����ui\=���T��.�y�O�Dvd�4j���c+ܚ�ybCQ�Bı�aV�n���!̔��yr/�=�~�������p�� �yb���ܨ8ny�'��X���C	�'�����ҒI�RuK��Q��(��'�b�:��QI���C��۵&T줅�7�"�s��&Hx� �AɏO�
ԅ�pXUK�E�

J��'
�&���ȓ�P���@?�J5�a�]�L��؇ȓg�H!{�∨�ju( ��2/��Y�ȓWt�x+�D�,(�Ó�X�5�Ҁ��TUV��&��q���J'G
�wW�ԆȓT�&P�˲X�~!q���)BD<�ȓU�����$Ak�M�pf��)�,��� `2
������h��J�t!�ȓ;�z�4EVDRP)�G+ǰ^9���KA��sd�� �"����b�a�ȓ&D��i�o͕0�V�$ɺ�"Oz8�����>���M�*��M�"O(�*Uh���=ȒE��P�A�"Oz1Ќ�?�I3tǇxv��(�"O�IQ�Ρl�" gԨ%d��"O��5��6$���7�5S耩""O"��G��o船�@�I���6"Oqk&��F�
�ڷ"�� �6ukR"O$}���9��z�C�j�"O��Snŀ;����!�����A"O���Å�%�rq��%�E�H��"OJ�J���ԬP�
$s��CV"O��](
�h*�ʓPD�`��"O� <
��X@ivgތu$��y�"O"��v�F��ǝ�\��"O��Sa��b0�a�e�D�޸�"O�E�1*�&bHYUMR� y�mc�"O�MP�G�9P"j�2̘�Gd�� "Oαa� �B�
aJᅌ�7z6���"O�-9��6h�Ȩ����!�Y�P"O�E���N�5e���7$�$%��"O�y���EVTu���\6	
�%��"O�=�Q���m�g�� R=�2"O���4�ʇ���%�	�V"O��b��z�\�2��&I���4D���F�6H��������j@�'D�0�7(�g�mHB�$���F�8�5�S�'}�q��e�z~���C���6Ɇ�N��)6�e�Q�
I������U�`���Z�;�:�X"�Лn�L��ȓj21�G�-5\*���&Tj�U��Gy3䫍*}���B3�E*Qo����	�<�W�S�g��B6L�>�����Ji�<)�	,N�
��� w���Ъm8�pGz���N�8�P0���+�0e�ul�?�y2�H�#f<1�N�#'�A��V���'rўb>�pp�T�m��%S���(%��4h��,�O��'��S�i��^��i�@ѳ(�p��	�'�e ��)\����=J+pѻ���'?@8��Z(��K��Z*=F� ��'��HP�c��	C�!�̾԰����(O��e�,�ж#Xh�X�"��8��I��U�be����8/�y�7/��`��<E{��'����5
Ć0��M�!���b�> �'�(��P�Іp��}3GN�(�#Ul>$��æ�Mn�I��o�cw0!�%�1�O��v�IYT��"@NQ9U��<`��ȓP��Z�`@�T��EP�H;橕'v��z}"��4�@�Rz̨Jp�]��^�Ĭ���y��	% y�t��` *jb�JsJH��hOj��d�1C^l���-��P�S.eɉ'dўb?-��/Nwz�Jg��0�F,�`;D��JE/X�<d4�	�r�R�:�O�O�Y��K4~�HY���]�m9��X�"O`��s+��W��U�!��1݈�"O0�3��ٗsFȱj���rU�İP"Oj��%	�=��!����V�p�3���q����R\��G��>���� 	-D��0SH�����N�&������=D��2�OCs ��U�\�t��Y!0,:D�df��8S/~ Zs@64[��q�7D�8@��dI�m2 ��O�`Ex�5D��Jq�7�
|P#���2~��5�%D�$;T����m���%U�@�GHd��C�H$j��u
�	=	�Li�lB�	@x��*ۨ���tDFc�C�	,"P:9�"�_�^����"��b�F{��4�';�� {"͇O�<�˥�y�,d-���G�G�6��|�2I?��<э�d�:/E29��/�m,�ЀC[:QA!��Gl�,���hY{]�C�"0*!�D��(���s%�hZ���bܛ[��hO��%�#�̤f�	��-H6�T�b�"Op��@ձ2�ր�M��n��T"O����*���# �\�v] �O�9s
ޠyΤ0*� 	77������<A�-dHAeY�XT��`Mx�����X�)� �m��ӪDn]"e+�!���"O�Qz�#ēn�l�銻'��YF���O,�b>�xB�"lD\`R�c���&�:D��)� 9N� �Q�Ϻ��ԡQ�;�ڨ�L�`��J�[a��s1�0re@`�;4��+��E��H0��扑6��o D����?�B�*�霝6Hjؓ�	=\O�c����NZ7;
�y ��\�2��r�9�$l�>�=%?��ɣ�b@�n�}�8��FF9D�PcF��6���p�gوH�(���d7D�d�0mΐsf!r7�Āb6(�J�5D�)�%�<���T�-!�$}Ru/8D����0�A�q4�@�R��ZV���%�D	�7B�QH�I�4Y/�̣ �,]v!��9���J�"Mz�V�rp�\
�0���$�<�D*�'P� �^� @���X	��ƭ D�ఴ#ܞ	�B�S�D�CC�9���(D��p�k�[��g#~�ցB�4D��9���3yV�QQ�cA!7U��-`$C�I%�J�y�)A����C�K&���������CŹ�n\"�c�92�C�	�fz��Sr�!,���fX8J��B�I�Y$,·C��]�|ꗉ@���hO�i3�	�,�X<����P�b��`b4B�I2b����VP�,�Hsh�S#HB���F��ߟB(!�KֳV!J	�ȓW�~��F��bg�X�2bӵ�~��ȓ��ס�.%���tK\�n<L��ȓP��au��qP<p��ĭc�����tU��dJ�pO`8�'/\2� 5�ȓ!?��@�l��k�j-)�e]	p�\��Q����f|�Ym���2�H�#1��cE�[��y�[�};��+T�'*�؀I�ML�y��
.�tc�H��y�@�!���yMɰF��ez��ϒk�V�zK��yr��3TH��r�8K�5`��N�y"� �-�'I1Ʋ)��g��yb��/d�\ٛ�,@�
<���j�y�f[?r����.�r���S��M�ȓz-�1B��}�PXSW×4��L�ȓL^ ��"J*I���"`�ͮ5�̓_e��0F��8Rq���0a�L��K�#[��yB&���Ɯb*:Zj$c��y"�@4!]�� �H�>Л�JS���>�Q^��˵%
7K^���6`Ψ�A%%6D�$	5��-'��|���<r�z���1D�܋�%Bzz��Ej�����1D��Y�-d�ɥcíL���kr玫8%��䅇B .!��+��Ѣ�DĠW[az"��
�/�Z��C�[�|�AJ�"S��!�D[�D?y��������҃"�Q�xE{*�&�����6	��j>Zb,(�"O���C���B0hDcB�=S�l�3�IBx����A�W]٣R�H�>h��6D�����
�m;tb�BB��L�SMuӼC቉<K
8��V�6P�=X��	9� ��D$��qV��'ЧO2���n�3~��B��/B"�Q𡂅s㈤sү��T�(B�I;*�Eb���T6�p���K�B�	�	�"Mه+�>	:��!��C䉘gE�YP+ 7.�5zjB*w�C䉪,�V�����ޠ����2lF�B�I6��X	�/�P�j��&2<�B䉁<��+�E͚:�j�A�rU�O��=�~� ���e����a�a��/ �چ"OrT{�B��EL��G�����"Oj�)R�)Qu�|��c/�1ʃ"O,�1�땧K��8j��g���e"OẕŢͬY�X�Ŏٝ1�:�hF"O���\@`��f�׍�ތ��"Opa�F�֌h�T��eJ�T���E"O��H��ب���]
1�h��a"OШ8��Cs��9�.˵R�����"O𠫶ɤ^N&�@�K� ���"O��P�߹]8����C���"OК�#�ql�)B��	E=���"��*�S�@Uƴ�Gi̷Odлb�{C�I�s��ɓCׂ0O40+Q`)[� C�ɳ{P�Yt�n�\8+V��=XM2C�%g�Ȅ2V�mq|���D�ZB��<jv2Aˇk	���(+��'�XB�I�MY�HM��l�x$�"�C�q�B�I7&��!�e�w ��*����B�	��>Y*��;�ra*7ER�A�HC�I���Ӗ(�!`fM�7��K�B�I:j�&�r�c61OC�b�B�	4v��drV~:.Y4�Bz�2C䉟oPQ�� �> X�Hu����	�'�A� %ǲ|��P�C#>mV<���'����E�9c@|�cOL�[&+�3D�tLBD�;t�̲s�}R4`1D�dy�JY�0I���Ǩ(&҄!�9D���g$M�j���G?��0���8D��F"A�nj�Y�wG2c� �O6D��˧	�,7.�Y
�g���G7D��e��f�|5�$�F�V�5��n8D��pBBH)�]�&�	'c�����*D�D3�-�*s���WL�[�xɠ��*D��� ��*����a�M�7-J���(D��7ˈp�r�u�I �"!Sg&D�8�B���tb5�ՆIx�PHC�&D����dH�4��e��C�h���#D����c˚'Y�a�V��1,�^|��� D�� ��S��8�fN�0�(��6O D�A�	%<���"�j��
�����?D�0����+:�FT�b.�)�Z��R�=D�,A�D�@ik�o؃�<�jWe<D����! 9;�RdSvE��G$�
�l/D�I�ǘ�7n������4^��9�)+D�4R4��5��B�o�Z���xv+D�l�N�*UlQaT��9�(XB�-D��#5����x?.]�)��/D�4���؉7f$ZA��9��Ԥ/D��j�]�	���f� �.d��c�1D��kt�
 @i<��#��]�b��I/D��cS��0�����Ǡ�R�R�.D��-�Zق�(:5,�Z#Hʹ'T�B䉊a��p��*S8ŦT)Ə���%��i�VQ�P&�	y)uAїXf��ȓ�$�� ΁#$d�Ճ0F�h�ȓj0����N��T�s�#���ȓ� ��6K�c(0P��Հ_I�-��?ZVX:���_|�|(�d�=b@4�ȓ\ٺ83�աt�6�;`ӻ3��X�� �d�B����I �B�[�tFB��ȓf�R6c�dEf	�@g���!�ȓ���B��i�`�⢮�5 ����ȓcP�c�G_�P��f�59Hht��S�? 8���> nj�!CY 2���#�"O ��'.F�^`"!��b#"h\�"O�SHK�1�������-L��yC"O�|�HC-&G� ��O�2F��i�"OL��a1l�4�c��QD�9�"O|Eib�"eX)�`F2E  �"O@�I�.� O�N�*�mۓ ��˄"OIr�:�,�D�ͻHoD��"Ob�rf�R�0���<|M�|�"O�Rq�� S��rR��o7JՃs"O�أ��P�wcX�Kb)�kN�c�"O����,	�`=�(�'	W$'��0��"OX镯[>��(��Z�@@B"O<x0��[æ1���u� �E"O�L�K�^�R��ǸE�4��"Ob4 �$ޝ)([QF.(�&�Zd"O�uR�-!�HB%K�*p��i�1"OR�!�&J�(��ͅ<؀�Z�"O@����Q�I�"!�	^�}���{�"O��A�(�0:v�Xh '���R�xs"O6ŋ�ǲ ��`1$g3Zp�m
�"OJQ�4.�(H_�d�TeF 2bP��"O�|�Q��+F|PBEn3Q,mc"ONHa�˛�Ua�a�5N?,@�"Q"O.|��&
!��a�ȱ,D [�"O�e����;P�L��@��
%)d"OXI�#b*%cp����ȋl	|E��"OXI0G��`�
�$���h�z!"O,�b���ڜ��lI|��1Y�"O���➈g�4@�X:��Y"�"O
�#P��Ht2����[�k�,��"O� ��5��y"�2=!p��"O��葉�eB�C	�_��s�"O>���E�o��Y0�	� �pi""OX�����Y��0�$�H��l*"O.�# ީ_�\�"��
Y��� "O����X$!xհ�j�eZx��!"OP��	eɶ�[b��9G0t3a"OR��BN�Zd9H��ԭ��7"OX<yvJ_�c5�(mR���WU�<	��0`"`��2b�.� r�mP�<�®F{��x�f���cd��3`�
N�<�eNåk�8�A7�U���	��P�<��&A��@k&C£!��۔��u�<)�g_^f0򇂀	(eT���n�<!���nMp�� 	����%�p�<�F��<iVd��Ч��[�i�͐o�<YBF��s��=�Fר�%�w#�U�<��o�u喱���!K�Aa_J�<��J5��y[��ƴ<��%RJ�<aWN��&]4����4
*$�U��J�<��$�e2x���4��(9�M�a�<!��=mq>���Z2�B4�%�x�<�m][�)y�N��j�� �v�<�Ѥ��T�A��H�5j���t�<A1�,6>�%�u͂�3 ��a�f�Z�<�b�R7U�	�f���z�6=#F��N�<��\��\��&�WhYP2��J�<Y��^$(R�0��C3n-F�+���}�<��Ȝ�i�v�Be.0Z�4s�}�<	%���|N��(�, fEX��u�<	��\����SY���+�y+7�� �d �Pc8��oD��yB �|ش��.h�02�
��y
� f���@�~@��V[�Nl+�"O ���_����W�^�˚���"Ov�k�)5H�<؂OA�a�)q�"Oޝ�$���b^���Q.��%M&���"OJy�'!Y��-bC�T(2fX��"O��bd�ȎUd�Ջ�ŵ4��8"O2�!�ԁK�h䓥hʎ-@m�e"O��Z"k@�\�s�.��"OZ�+d��P^�9��M�}pt�Ss"O4T�ac�#Oy�s#d�]U�Yx�"O�i��]�i~
�U�I4c�,�B�"O�Y[b�����A!	5h��=��"O�h@�ʀ:*Î����/'�x�YG"O�!����-6�B�!���☑P"O���▫FW�J�O�&mZp�$"O�LZrHS2#����n�0k���"O����
�?O#�츑�̟H�����"O���aK��t��}բ�9D^��"O�-�f@>)yT[UCʢ5��)��"Ot-�D)PF���A],_1�� �"O��q�+	�l�:] �^''�U�s"O����cJ> ���l)fٳ"Oli�%a�*7
���GO��Dt��1"O�}#�F� [
�
!���[f� "OZiSgo�Zk|pCҎ��iU�|�"O$��4C�	6C��X�m �.\�(�"O��K�����NE�F�� "O�Ԩ��!4�h#V�	8L�8�*�"O4Ek��3X{� ����B9(��"O�`[4�N�lE�2�E@q�\�k�"O6��R�H/�B8�ѧ��_$��"OV-Q&A\�<jaq	��L��V"O�pC��E3�����kc4	��"Oh�"���ZN�ay%G_�]�"O�H�u��wZ8�QE)|����T"O���CnD�nMj��ä��L�a"O��Х��'x@y��f�1)Â��"Or\Y6�4p�2l��F���8	�"Oμ��.}2XtȂE�6�\i9�"O���Ƅ�*'�+�bܕQ%�Es6"O&����\�+C��#b�F"I��"O�4p��R[�uKԇՊ`
R9�"O�P��DQ�1�vHa3���1"O��&C��V�\�ڃ*�����u"O�@ؤ���M����hX7\.$ɁE"OVh*�n!PP����268Ī�"O�� F�>F2tH��8<���&"O��[��
4"�{�!�G��)#B"O�(t��nl3���}����P"O�8C��8$/�L�P	^"	BJ$�6"O��q��؝^�%��
<Nv1�S"O�,b'���.���A4�I�E[�ʡ"O�����9	8BiS�N�%B��c�"O���E"G67Ҹ�G��\+8=��"O(T�#(J�`�lrWNI�*T�*�"O@�PƤTg�t�SwG�� ���"O�yC��E7<4��'Uh�)I�"O�A#2e�.^��1��1)�^�33"Oz�;���$+ڐ˗@^5Nm� ò"O�q��Bƻ
��ؤ��"J�J���"ON0S�&��:m�����ޥ L2E��*ON �!�.�����'kp~��'THM��.�c%T4� h��d���k�'
4쓵�Ogڴ��� ��U4�)!��� >l�s� �I�P8�6@ڌ/�@��"Oʁ�"D�X	j@�6��y�jEK"O
�"d�W,<��9��ڏ`�A��"O��g�ɫF"� R>O}xԉ�"O���6$�!�C@^�Dn��b"O�&�� y ��hv"H�a"O"�	�L0 M��![��3R"O�}��	�vV`���ALhOj�"O4�7C� �LI�ƒ�QL�k�"O�9�DFK�Al�aA���*1j�˧"O������f̸5��!�'2t"Od�k00`�
��g�K=N�Z|��"O���#(u��#���1ʭҥ"Oz�*f�ܕn������[B�P��"Ol��Cm(<#80+v!ی|���'"O��1�E��W�u!tGR�z��` "O2duN�8�xix%��Q�&�I�"O�����6�Z���ETT�D�Q"Oz��ND�m��A`�)�	ت�C"OH�`�H�k��li3Y���i"�"O|���M.o��ɑ�U/vި� !"O��LR3iD���]:�l`�"O{�+����I�4$B�7ƾ��7"O^�c.Yb���!TMUAI�P"O2�j1� +
����"��~`*"O�1��)��'�%Q�ڏ���v"O��PKP3V�n��O�>�"O�����$% �� Q����"O.@����/{�ӆ�M�0q "OR���hAu��q�h�3<�h@��"OL5��/C�~��H���Y�"O�9��FN�dC��a���w����"O�T�������ٔ��8R����"O�y�DI�>6e恁i�L�)�"O��&"$"��T�fa�:S���"O�<WE_��)�4 �L��y "O��ʥ���?s���%ϙ_7��"t"O,Y1��]V:P�#��=FV-PG"O�Z���.E�,����
@�}h�"O���Ɖ�X�\e2�f�70I�A"O���"�\�x��-;�&��lN�=2�"O�p�c�Y���B�!ZR��"Oha����VP 8��ɾO9��"O����dQX�( r�E]�; ^9�"Oh{2^&OH����e�N|��s"O i����PG8dx@�ڲ$���e"O��F��+�M�eZ��p�6"O���#�:H��Bɹ{jFM��"O�A�����b5���Q!@@�"t"OX� �n�s?�}�� �pW��b"O�C��I��ɒN�iW�P�"O������.t�L}���3B��r"O�����UZ!��Ņ25�Mq�"O4Q�i�IY�H���=|��"O�}��Ȍ02x4��TXs����"O �mL<H4�C���k���"O�Hd�]$hE�,@^r$�0f"O�4�R��d�!P�י|\��"O� rs�C��l����$U\�Y2�"OԈ������� Rv$�3���P"O|�B�m�#�T��c)@�m�&���"O�l�v(���II�#O��D"O8���,@�|s��9\���"O�#+\�a~r�R��^>n*���"O� ` a�E
�z���BU�ڇCZ��e"O4���n��5,T��G�\����w"Ope!��U8V���W�mh�"�"O���`kX<6�y(�!��&`h��"O���f�Ʀ\��F"��>D�P��"Odċ�FѩLOBŀq!��P=���"O6���V�K�1s Ɣ<{7����"O��8v�@{��I�%S GU`hPs"O^-kQ�7:�|U9��L,J�Ba�f"O���=��5�K��j�Pq"O�|�SoV;	&N�9a�U�Lq�չ"Oĥ�4�Փ5�����/
�YZ!��"Or�2�R0
HL�i���"O|�«=:T���4����b�"O8]���o/�ʗU�E�a "O�K�N�<D
rl2�N��d"OpD��i��V��pC���m�Te��"O�V/Ɠ�8��VAn�z�J�"O�L:�o��4�JVG�|�t���"O�ISj��=s�`SFo� ^�t��"OL�q �Gdx� P��#'�� Cb"O�Q��S �%�G^7/���9�"O���A�,8�,��
ٴl�F�S"O��"��2���N�;�&%`"O��'��cװ!����C0"O:�R�!��<��A�V�(gFU�"O����պ��HQ6&�-[lP3S"OB�������dL�'"r<��"O���0�����a,�=����"Oމ�7��-&���l��i �hx"Ox��t�G�g ���>\����"OH<#��$~�c�� ��ݡ0"O\]�"M07��r���jt�Cu"O4��i�5E�Z����D��Q[�"O��V,��_��m; �߸T���� "O�@�c�kc ��AE�"��R"OF(A&jFJd�8����^�ڔ"O��(��(Z ]�����z�L��f"O�i��%X+��.T%D�����"O
m�  ��n�H���pb�id"O��%h˻���A��Uc��U"Orc���q�x�e��H�*�"OőC)�[�ͫfV��d��"O�Jq���&��("4ʜy�.�I&"ON�I��f��'I�V�8�8W"Op�ktG��u�T������.��"O����?���Dǆ�.�0�k'"OP����
\ͺ�Z�#5�MRS"OpQ��!)'~��"�ˊ� "O�U�t��'3n�˕�R�A�4�(�"O���2��>䁹��I�W���"O�<��n�<W6 �����I�"O����(���HD�=u��H�1"O`<!ŗ�K4 "��/\h��"�"OH������� ���E}J���"O� ���U�W[J�RVKI�/� l�P"O ��W*;����Jܼ��}e"O���%h�f��+_V|�2A"O�8�F�R�`K�9�$�(�P"O�����	l7�"�}���"O)K��]��E���0 (�؁"O��t�����:�:""Ol���
_z���a�(b���F"O�VS����Μ�ogx1�Z�x!e"O� �!SC(N�8b`�M��a�"OJ�+�eWzնX�Λ43��)��"O,Y`WJ@,KB¡h��F#B��]��"O�E���$:P��xׅG1Vv�Ԙ�"O�;�.Z-`����Ҧ�{�fU�2"O�\�'ے~���5�W�u�"O�Ě��և0N��5	Ї@��R"O ����$k�u2�G�:w\�6"O�)�wKʕp40T ��"
��`"O�!�6@P�m�B�炟�
.���"OH�`f�����"�1\�t�@"O #&�:8s��2�aD+"��,�%"O�U��I��z��g�S���`t"Oh=J���$j�h�buMкglE� "Ot �!�
8J��&*���ȵ"O��(�OY;�h�ؤ�'n�Z	��"O��f��>������J.n�z]:R"O����� �1�0%ݔmĜH�w"Od����Wu� h�$X/B�z��"O����D�y�����
c����yRH�7?����ӻ "�p
H�.�y�C�?���p$:qĐ˄*���y���caQ���
T�TKS
�ybgձc���Ȅ�L�S�e�Co��yr��;c3�-��&X�G�h�S� ��y��@������\�Bg�]�
͙�y���z�Z�k2,���l
"G�3�y¦]~
�L���X��D��y��c�$�1rǅ|�J��G��y"/3L��ԫ�Hs6�dC�J���y2�czh$���S5f�,jd�F�y� VT���"+1�������y�B ��� �%G�,{�<�d���y�úHo ɀ���)��-�zTC	�'����!����Є��Nɼ��'�v�J#�ĢM�,x{ ���/-j$p	�'4�)�����3F0r�ȏ',XT��'0B��H ��"@��*����'�<◠J+P�X7�B>
4����'ǺM1f���+�D�)N�}�'Zxec��)-�6p����J�lS�'>@��g��E�$����H����'�v�:�oD�m UD�9Q����'b�9A-��=[�i�4`ɱDEH��'��!a4ꊝ����)�D�&�J�'���ȓ�ۣu��h��!5�2m��'=��EUg��0;�L�|�0\s�'��u�ȗ"(�t1��#��r�dI
�'��d���!]����MA�&� �'
��iT9L X�X��A�b�D}��'��I��FSo9��Ӄ`�ؤZ�'Ŵݣ2FF�]G�7ɋ|����'*ܽ��m�V����_�T�c�"O i@���1�:CMI
���"O`���W#|M`9S�kV'I�VŐ�"O�!�bώ=bS�0!�p;$�H%%7D���$�>���h0���i�;D�x��S�D3Z�z1���@
�i�d:D���щ:�V��`�"�^q:B�5D�Ly@JH(G_2���E�_n�*O��%��'.~.�j���D��"O�}(��G�e�zqc ��C���qq"O|`���*��S����X�6"O��z�?iH�à�5����P"O� �m�J�-CW�u�o�F6|��"O>��f�`�(���^-p�H���"O�9�"�ƟH�A0ULњ i� ��"O�:�h�2 T�ѓ#��3`�e8"O�����6��RH\�%��#"O@�����k���+3�[<�ع�3"OH��P�5!��� �M�Yg"O��ôI؃6�JI#��5��f"O ���ҙ2a��c��j�|�v"O*��A"H�6���9�ĜJ7��HW"O����MB5j��S����A�jl�4"O��ꠌ$i��*�B/G&�Xi�"O�q���ːR$�򓠄��z"OD0�VDP�b��h��D���8�"OX��JȐV��`���#;����U"O�q�煭)� �B��)f"O�\�D��Z1��
R�A���
0"OfL�*F�,m�6�]�8v>��"O�a �m�:Nr|D:�'D�n�-y�"O~\�rʹ?L�`�ȠaUV���"O:T�ǒ�%��Q��F	I��"O��ZE����a���Va,�XBW"O��Z�� ;#��eJ�<}ֽ9&"O�l�)O�S��y
��MLi�I�7"O�l��c� �*L��M)+ �J�"Oxyq�H����i
0JK29�`�"O��'L	�3�.�K�FZ3t��$:�"O�dQ�I�Ϻ�����x}:� �"O�CaB;;����j�(	d��C"OVtʡBϻG~R�H�	ވ
Yq�b"Oޝ�
�t�	�pfI><u�U�"O�
u&�
!`�g�ټxZ*d!"Oԕ�G\#<��+.��`B�"O��Ұ)͞I�>��2E��~���Y�"Or��w��AAt�P��@x�d�X�"OD<I$k�"T/ a����j��$��"O�  �ϡ$i���iN)t��r7"O�8`��>5h�C�)�m��(%"O�5��T�YŇQ�<�"O�%��
�15,d�ӆN2tK�(��"O��z@��IXڜˡǌ�*��ږ"O�8���+I˪������Fr4"O�q�p�9E��IV���"�.���"O�Y�#� ��{�˖'oÔU��"O"5[��W�#�T�$�>�x��A"OD��!�A�2J�z�
�\�xH9a"Oh�+S�F5> \�Q�[�H[�pd"O@�kל2�n(!d̆�S��!�"O
���	�B��"nWtR����"O��s���4���9i��H�"O�9QL�`�*my�uC�@��"OȀ2, a*� ��W�F��&�'���'��Q�#1h��F��	����r�b�'B�'�T	bt�_�8���b����'z^����E(,��D�ulR�*�L�p�'�@�I�F±�lK�a�V'P,)	�'��كP*G�X�宍�\����'.ĕ8���"
i^m��FP"=�����'
8M`��԰��1N#G+JU���?����?�򊒲 ���!ќ.عTd]��?���?�	ߓMnR�a����b�2���X�N�T�ȓm}X�h��l>�ѶaKV]Y�ȓF-H	�F�T�?��9Ԇ=j��ȓ{j�b#��
Q�hA�(C<t���S�? ��Cn��N�$=���-#��s�"O��q)6\���1��(�XȚD�'0�'Qb[0�,RV/6.uy�f� 13>��'�r�'�h�Q%ٴX8�R�U�g��M�'V��q�Ǉ!�Z���ϞfU4�z
�'�R�P��$A|�0��O"eO�t�	�'������µ����'� S'�I�'m�I�JW 5%��N-Q�x%p�'�U(5�V.o�xu#�^�2�p
�'�,��!�䈆�AS!��8
�'�� �[��E�@��8T3�+�'BC��٭]�����m�Y�Ĉ�
�'��H�Ø*E�L�'�HY���
�'~�1%#ܣS����U��--2���N��A��(�sv4�Pb>��|�ȓz�@|p֍��?b���!��X�(�ȓuC�P�r䖉v4d �_#M6h��ȓJ=�[�$ӑ3`�&̢H%�ԆȓL��`4��h��L�ڛH�p��8�X� �T͚9#ӁÎH���ȓX26Eqte�sg���R��)<^�� L�DH��r-��C�y��	��bo��Hn�??�<E�4HŰ;p`Ն�	Uy�N�5za8<Q���r"@��͏�y�e�Yf�B����5�,xp���yrH�9T��qsNߴ*z(Q��� ��y���n^V|`�o��`9"���y���?"��di����Vn5��K��yrD�"�j@,=��K���y�	��`y���$]�W����yrɀ*���JS&�2�8`�N��y��SS:,���I�1Y���+�y"n�(p���C���^��QF%ݮ�y��^�U�~��ゔ ^i�|�f��y�'��5�Yb�_D�b&�ߑ�yB`ʬ6��q3�
FL��ctmT��y�E�b��H�5Kƭ=�Y����y�^�r�zOݪl���hC�٬�y���fh�dɋM�$��L�y���h_�8w��$F�:�����y��"V�YS�jQ*:� ���d���y��>� �1��)Af@�(AD�y�D��#���M�3�&�� ��
�y�%�b@�Te��1'ΰ��-��y��Nu�����lƈ{0
A��H��y"�g'4�"��ŕe��k�)ȷ�y�تG�D+g&�,7v�Jփ�y¢� gH�$��/����B\�y��ZfҍD�_S�H����y�l��.}�����R
��6nM��y���>*��j�jM�w��p�	��y�Ǌ�/_j(s0��:� YƊ��ybBJ���X��ʼ{����j΂�y"�E_�0T"��lz������y�iY:>���)�آv9`qy���y����
�q����ǌ�yB��:K����d(V�fN�ew@<�y¬J+0XM	%VY�t��fJI{�<Y�C�$6�ZTb'k�)	i�@�z�<���E�{� ��f��EX.�B�o{�<y4ɐ'$78��(P|i�6��|�<�a���D����!xM.q����c�<q�-Ϋ?ypy�!�X����c�<i�j���ӄ�� p���f�@Z�<� fȱv��ϒ8�@�N6H~�P�"O����Q�>��||he�"O���I@
�ԁ��ɫ`d�� "On}�P��H��·JJMK&�sv"O�X;�k�/g�hkj(A��""OL��Rg��M��� ��!"����"O��Qu�P�CkV�1e.fc���&"OB,I�ݩCA@X�BJ!=E���$"O��	��,�����4��"O�D��>jtȫ��YV�"O�4%�P?���R�N�7����%"O�c�jˈ?İdׯ����U�""OEZ&jA�V�;��Ŏ$��!��"O�M��QD� ��4go:��B"O@��vː�&!���	]	h�5!s"O�,{��Ҿw�X32�U-	W��)�"O&��CȦ8� ��9�e)�"O��B\�1vN|+橒&H@�"OT���-�:�ja'��,b��"O�8��I�F�y���� Ih��"O`�q�����4xjg��SC$��"O������N��[�1�n]P$"OШR�oI71 ���� �{�Lg"OL}�J[�+�t�
���"O.@�bɔ�(zt�"��I�v�h�r"O�w��-��J^�e��#��f�� �ȓO��Dm���K��͢q����ȓdc� I�EE �9Kd8wd���Rkb(q���/=�m(�d+C�҉�ȓV�åC%Y����/SWHn���[�x�h�%<�4`��	qd��ȓa[FT�+�p�P�e���ua"O���F�B�l�"��1�
��tAa"OJX"Y8�ʑF��cyH��QB�b�!�H[0��U��	P�#ŁٙQ�!�d�:���J��M�[S@#'��q�!�$ו���և���� �Ò�a�!��º��|��f�>-�$ؙ��0q�!�ď�c�U��'?��pQTA	;=�!��
k�&��S��
��U+�AZ�.Q!��'�$Uc#��0���@�BF!��F��Ya�(;L��LR@�x9!��9Rp(��@�)?�&�1�H٥9J!�^'`1���B���
4�U�
�4�!��>������1ۺD���C4K�!�D@XJ����X�£a�7}!�D��9�P+�KP�e�V�*��ŋoe!�$^2^��*�+��^�@��1h!��Z�Li�w#���&htɀ�D�!�d����yàgɭVj�\!V��!�D�l�����a�7&o*X8�!���!�H�t���k�ln
�������!�y����დ��hq �5!�D�3]:�
f��q�����8B�!�D̹/�����e����d�Ȟ	�!��G�
�&5����`�ب���U-D�!򄓇7���'d�h5���Z�x�!�$Q�,p	YQbȍ
��P����$;c!���;Y�ɡ��Z��3��8
X!�$�3H�Y6��O�~����!��þ4;�i��h��aa�Eſj�!�$
&�P5`�6@�R�ʵꓴu�!�$,`5ʵ˄�Y3h�W
�)�!��;`�)���@� �Z�;�ŏ=�!�� �����8r�� �J����}��"OF�����rd�0Ӆ#�9/����"OPq�ը�@G��x#ΡFc|a�F"O�}@S�*<3�aT@\6$x`���"OV���I4nh3�o	{f2�q"O�Xk�bC¤ �tN4)q�"OZ�@�'C0�
4�w֐;��*�"O0t��Α={.\��qb�"7vpZ�"O�i�F	X�`�Li��;���"O �Rũ
O���军�g�t���"O�!(�,ի.����eׁ�Еz�"OTł:c�TYQ�9>zV�HP"O���K�$�^����V�f؂�B"Oq��E�ta �C�����T"Oƨi%$�]��4b�Z�>Y�w"O����+'6��T k��a��"O�r&�C=<�N��!��;���"O�hpʚ*rZ�)��/�9�2t8@"O�YsCvϐ��+��
*,Y�}�ȓMҽ��C
ِ���i�$vct��ȓc�%����%�ЁpK͋zYڔ��(��!#�0�iQ� �!�܇ȓVTxb�l\5���"�K���ȓv�v A$�l�����Jf�����B�s��A/A���N�"@n@�ȓy�� @6� t�:P��?���ȓ	��Yщ��F�<J�
@/�T�ȓ&��a�i�T�)5"ӣ31�ȇ�nꤽXfg_::�]�P��H���	hh�!f�{��-x�*�k��Q�ȓN�p1��M�J|�<1���<'wPd�ȓ��ӑ��+o:��S@Cch��ȓ6�b����"�+�$Aa�݄ȓ>4�ي���%q��� ��$j3�E�ȓw�ŋ%� m�8��)���t�ȓ���䦔=�B!ہ�&a���G�ΕX���n��
��O�B"�}��Q"� ���U�_F��4�W�2WP���;�<��ыC�M�l �f���Ph�ȓk��,j0�G�Ko6d��n=5����7���f�7�՚��]1��ȇ�7<�P ���Dz�Wd��gۜŇȓ��H��F(!-ڈ���Yi�̸�ȓ|L�c��Vڬ8ĝ;��q��IϦ�� W�n\ @�_#@0�ȓ b��c5N:�( 0F�J�j`�ȓk�i;G���lY~��p;@5<(�ȓw�4ԫ�A�N�l�j�̇8]�n�ȓ)J�$�`l�5?�5���Ϸv Y��wԠ��#n�h�l]��G-my��Nf���oN�|���CC�.�L4�ȓXl&8�Sm�[7�sDP$�T��ȓM���z��Z�xG������~���ȓa� �s�J�M�drDF������J�2�@I �.��#¯�J�x�ȓ%Rp��m�v������
J�f���L�L="�N�-$r��J&�l���@��,�w��8#Ăi�
��P
���{j��7�ʨ8猔�$�CQ�؆ȓ&��͢���1l0��)1��w�B1��[�lB2'̠r�,�1nҳ/c����:���*R��tQ �[0J�Ұ�ȓ?8��iX�@6�u��vNe��^�(����w��D����',Y,���S�? Qqo�)�L��\�~��qz�"O� I�81�����d$��9�"O
Q{7J��/��C$�Z3|Lܓ�"O`z�hA��ʩ�uàx�.��0"O�`���� ��	Z&a�,N��`�"O6�	�ř6�fX#g�B#*�`�"O�{A.�/�z�Y�E�4��x�"O �K�@�b#����$�L�!�"O8�����s��}Z'77��}��"O6i�Q,�*|݄��%*q��Ed"O.)���?�
M�s�[.6����#"O乱AT���1P�셄EJ��"OF�괢I##��}{�-�<�#�"O8y�H86�:0�w�J�XzTc "O:y 3�;��L��+�¹�A"O�X��
���<`��n�n��@"O�E��(�$OF�yb��
&H("O*�е*^�-��}j�K�*S��R�"O� (���h��!����(!�"ON�PӂM�CY�xs�4v��}c�"O�]�fM��v������Q�l��"O����L.��|ض$����4"O�b-�=F0��.$=k�"ON�:��<��r�W;)���3"O��z�C�P͆�z#�V�# L�Y�"Ot�2Q��E2\12eӪn��""Oν�"��X�.Q�D�P�i�F`"O��;�V�cz<�f,ItL�T��"O����R`�` �ǡK*Nx�!�"OlM���4 
�c��**��"O�!�FN�sMv,◫3;��F"O@$ya )3ߴ�32K.;�"O���sK�&|LWF��'nl*"O�c���"�t(�4��;C^ ��"Ol����uX���uݱg�xP�"O�i�J^�ܐ�!
�bq�7"O����� fdI2�Y����T"O��doC2F�P�q�/�U��HA"O�Ts���㢑�!����"O,�z�/�A�pDq%̓:k��Hم"O�*�ȋ �2�%�.5F!�"Ob��Xa�LP�.�&)@�"O2͈v���`AnD%E��@u"O�t�Q��!qx��bX0>Bi��"OB��G o����
�{��$�$"O:����;ld����%0��`�"O��k�U�:r�h9�E�S���"O΅����1N �{T�K��V���"Od5�Hݗ%�,��4��u�\,@"O8��Rh�hi���C$	�(a"O<m1!�0b@r���A$¦"Ox
�gްj!f�`�ј�"O6i�7�
�t����BICu��p�"O�i���4T��hI�(���g"Oh�j&_���������	�4"OJ�J��^T�rᚗ ��T�n��"Od1�&��=V�`/�>�{�"O���d��^�^�9��T6�:"O|�
��_�v��9����{۴�r"O8Š�L+Yh���힣j�"t�"OHu`@�I#��E ��M�J��"O0��!N�L���V8��7�8D�0�t�D�[Z�Qr�C�9 �r�2D�lyC��04L���#� s<
%�w�#D�� 2q���O��Jf�ʎx:���"OP1ר��t��1�R�gex�"O�} %��{����ӣ;�ȱSw"O�x�!#_'����K�gJV�@�"O`��C�'�������R*t6"O�ٺ��eP=��̡�j��"O���K$e�(`�֡�5;-�a �"O�l������<bv���+�|Mi "O��΂j�����NR1c�n�p"O�ɁuG�&�,!9�nh�X}��"Ol��'��W3�mA[��x42"O8�I^��2�I�G��e�VQ�"O
ȪG._��HҠS�n��]	3"O�D�1%��]�,є�������"O�B��·�(�3
� �8� �"O ���@�x�0�2ȃ�w�zu)�"Oܠ��½|��!�L�[kh ��"O&����V
c	L誖�4AV0 i�"Oz X@��!I�JQ�	K/
@��U"Oxq�ϒ+�"�X��ȡ)�ѡ�"O�tc1$/K-��y'B�9R"O2�I�F�5_F-�� �FT ��"O
�p6�	@�P�E��ZR�t�"O���\Id%�Kƕ2>0qQ"Op��$GX� ����) 8T8" ��"O�u��k��7��	�q��(�<���"O��F&�0u4��ΔS�:�"&"O�Qx'��Mڼ���	�kx� �V"O��`��,f�h���2:jy8"Oj�ek]�~���p�\+RiC"O�l�v�W%%�P�����%f~�kC"O�	�򥌔lQ���!��	�V"O�X*GDU�#\���HT���+"OZ
 �R�3p��ǀ[�~�x�"OȽx�@���F�@s&��"O�͋�l?6��Gi�\5L�r�"O��P�hP���:���S�|	�"O<Ց�i���R̒t��OCpQ!�$��U�z���J
�̑�g�W/%=��D¼#t�'H��*�SAi
��y䗖BͮY���P6|s J�@+�y"�S� �p@�@�5?3��`���y"i�[M�X�P�H?:d�9��\�yB�<S�)�3ۚ��� ���yb�/o6���6��L���4)7�Ćȓ2��sa�F/E�z���%ޚcZ���~ecE F:`R�	�J��D�ȓy�F��w���(�^8Y�d�Y1�ȓ��a���3,Rl ����#}�
؆ȓG�ƕ���.
�X@Sl̡bs,p��6��Hc��;2�6�;�K����8�ȓF@Y�t�Պ0@���g�U��}�ȓT��Q���]!�p�Ǡ!�h��ȓPp�]�G� 01x؈DoCu�u��O7�p�fcQ��V��>u��N!��� ��=��o��.Ն�w��eRw!�>��R�J�yr�=�ȓD����A�H
}?�9z�&7
u��ȓ��xX�� � �y���2x����i��Pc,J=Z婁D#L���ȓ��D�$.3*��iG��Ѕ�F�~���ӣh�Y��
�|��jrh}��D˲3�H���L8D慅�V+:���� u�,{��׊6��H��S�? ���V�*�5+�+T&*p�&"O$�S  �L�xt�ӊ���XK�"O��!�ˎp�2m�ǊC���C�"O���l��rU��I�jH0�t��"O���!�8v9+��ǋpa�q"Oڠ�`,*�R�tpN�SF"O�l�Wc0F�X�6N�HV��3"O�8 �*�i�4�`փVD���"O�����>t�7n�2L���w"O��!��+1����-t��2�"OfD����P�,��☷IHd���"O��y�꓈D� ���

6|@��c"Ot��w	aP|A�iĭ@̦�9`"O�aE�_G��5�3n�>>� ��"O�`
a��!=n�xpխ�,_(�e"O&Q�C������ÐB�Z[�r�"O�� �޻|��H��A2d��"O�H1�5D2�8�Q�N�g\F�Q�"O҄*J�+F��@V��/UE�˒"O�t�D��D�$*�D(XAR=�D"O�yZ�dF�*��+�ݔP,\�"O��&E5wiI`�K>����"O� ('a�:(��(�lZ�{(vu)q"O�b�+܇E��8r|�b3"O~ @�C�}q@��\tJJ�"O��Ӆ�&:̼�(��G^�`�%"O.5�1O��ȴP`g�vT�I�"Oе��F�b��u�F��*B���"Ot5��޵fаH37���^���"O��3�
Փ7͎�:E @�Ĥ3"O܍A��׭o]�����p�!�g"Or��C!�1M(�y���ڳ$ޘ��"O�0��)]$(e��1,ߵ�2]��"O�$��G��Z�����I(<���"OB���l��(��xE�6Y��xȲ"Oб�Qd�=�=8�E��ؐ:�"O~P�dY�g�(��UӘu��)�"OR��p)��9�����'��Es�"O��*�d�:-�S�א�H���"O�+T�!5ԩ���uh���"O����a��!��GH=FR���"O�%��iH:Y���3(ͯ9�p=�D"O��j��Z��$��tz͸d"Ot��s�͞8���RbCO�"�l��E"OCSL½0�0D���"��a�"O&��ebxFtt�t�J�XW:�pt"O>����7d֞�+"D�8F�(�"O\a���U��L$�a�6I:�]§"O ���2�R�p���
Qm��"O��:1����'��o�LŠg"O�)z(�"zd8ɐa��#�Z@0�"O�KF�
�@�1%���At pY�"O��cF�S�.�3�n8Y!�"OP0�Y)4��Y��D��tGḄ"O�8ӧ�
Y����Gd�>�Dl�"OF�2�N�H"�s�A�" �6Q)�"Onr7�F�d��蠀B:1�9#�"O��Wb��@���qRA�9Ϝ���"Oq� &(0� �@B;�8���"O0���7�9@��l���Ɂ"O����1�R����\%��xD"Oԉ�e�oaV@�.�9���"OƱ{�)�a`|2����B~d��"O��d��|˦�
�l��~b�ڡ"O� ���WI�**��z̟0�(Q'"O �cŐ�Dͤ�@���. ҁ+�"ONIs�qtx�b��������"O���M$�2�R!��O��=AS"O��H�L�u 7o]��E��"O�U������y�K*1�`
�"OQ��JF1(�ܚ�վI	"9��"O������O[X����Y��b)�"O�e�CܱfI�1���87�>��`"Ol��G��= ͞�iU�@s�=�"OИ�ED]�.W8D� �ɜdV��a"O�$i��)ElВ�EZfU�]�"O�0�)�s�0\��ϔhS0�A "OZu �Iߐ�@����Add{�"O��3Bȵ^}��H[�D�3�"O�x���K4{b�(!c��T��,Bp"OppP�G�!;�H�9�&Ր�%�"O(�P�(�:2h$�{���Q3~u�v"O� !$�Ģ�`�[b�԰t�h��"OH��`��:=�AP�Zi�g"O��+e0q��a��ܗ-�T�"O �+���-Y&jT�A��NX)�"Or�p!�,H����� !~�Pd"OFD� c�9S�!�@�K .y^�{"O>��Ś?�
<(�.9>����"OJ��K����l�7)��P�"O(y�`K\1E��t�0�3@Ǿ�'"OP��-�h��(
�+J��<=x�'��,�c�1x�\�3%ņ�V��E�'Q\�Y��� p����M�H�~:	�'���re��DC�,˷C�I��(��'Bp5q��̪b���㟦F��q�'�ec	47�J�gEIa�'�nY@�����٩�oBeyH<��)��j#�"�LF>|z��SA���C��-�0,�0�	"����)���D�鉊n44���f]��|%�S�Z� ��C䉻<{e�V���%C^��6L�D�O �	Vx�D��m	9�&��I�&*��B�$*�O6-z����
$FViy$�ԉ��t1�"O��if��2P.@�� IT� �#��j�O:	�'k�"1�a���Lh���F�O?�c�F�;�h�#!i�%�VL��'�Q� F	´@ �ZR��)�'��Ð����Cg�(G����ԯ4�	ɟ�G~��/|�F���+����o	)�0=��4��'d�z7��U`������?+x�#@��O>�����d��0$V?�(��sA��$㟸��f>���6�Ex�A�
�� ���Nza|�i���00 �EB%s��e��	�Wߖ��Q�ɬW\Q��'��a���%z9,���䚍�^�FxR�b���	����@ ۳3�΁!"(V�!��	)�uڑ�����f�Y,��f�)R�{�� w���r���<��z��B��y"E\4 �B�6	]w�6���'�����O�=�}*�E�&@p��gco.�#BlX����'s�Ɂ��Թ / 0\�a#�����<q˓cb�	cŌ׽3�D���@����<���󉙻,�����aY�Y��=(d/�3zܛ���i���C�B�I������&�:s�,D���O��<1%�4W��U&%D�x��]�x)�[5��&^��!�i%����;*�D0cf�"M$|A�̗?l�C�It�\��h�+_�Bi�r�
Sl�C�)� >M��j��J��ؤH�G�[�"OȬ�1��~�`�q�h&k���a�"O.�9�Lߙ����P�W�`A��p�"O���G�F�;�H��M �S(kA"O��k^�{^ ꁌ�v��L�p"O�u�#�9dv��y劙�v�@�ʷO<���]��4���0�J��X?��_�|��ɴy+�hLߜ~p��cd葈����$ۜJ�$�<Q�G��c�J��*�r0�GoI�<1r�;S�dZ���5�����H�<�%g� H������ �� �DF�]�<��� 5SZTU���>i���\?�N<9�O����D�R��,�B�׾.4��H�bϳ*!��ϦRIh��T�C%4���*�W�B�l��l!�BM�\���n����E{J~����B��X�b��Ŕe��Ur�<��I�ip �Ьݖ�-ʀBLW�'kayB������L�#{Tys�H����xR씽55��C�[}B4��w�ْ*�NU�ēd�Lq�c�}�X���o� �����+Zd&����#�,�B�.0�2iS#O5D�����$k���e���zM7 �I���l�?�|�G�-d@�flM�9yj�c�<!an��
`�1�E��0���7&b�'�ayd��/zJl����7TњHX!b���y"'S)_�EKqa�Hp@�����Mk�'@�"=E����t& LbJ=D��3Q��yb�F���1��Q�S&D�! W5�y��S�Z�q8�/���(�ȓf��-iF$&�0��fEOr�e�ȓ J��$'��)�v�E�ާ*���&�xG{��tBDc�3����|s��TM�#�y�NV1Z��Q{ �P�dq�%@�y�'(��
N>��O���-'mC"m�k�v�1#j�3`'B�ɏv�n�z�"���Ź��@�D�@�>ғ���nt9E�C�m�8�Vh�d�!'<O�9�}B�N6_�Q�D�> ��ʉ���9�S�Oޤ@r�Ί��H�&iҰp�Z�K	�'�u�F�42W��$��\}�<X�'���(�.]�"�R���J�L����'���÷�L�Q��a�G!P�<}*�X��d����b��1M
s�LՃA�P<r��)��"O�]�)fR@$ ��O+���"O|�c�$�;I��5s�k��mhӦ"O�8Y�hE�+Qz� A(T���=
G�4�S�	Z$��GX]��p�f��V!�$
!y�^l�w��$-��`h����p����O�p��"�0&��D;���j���"O�=����� !՘JO�9���i9��$�J6(p��!y|H��dY�R8!�$�'nl1A���q4�Q�fB (�d�(O&�}J&�͏QdHA��nG�EM�8 E�|�'&�yb��&0���!�Y�h�R�H"Cӏ���XX�$�0`JqMZ]h�!L!V��8�Bg8D�lq���X^0Zv��<�hӆ"D�����'�\|��d���=�3U��xR Ȭ.�b<�%��w4pp�j���0=�F�$	{uf��PoS6,��(�H�!�J-;Yb��BM_�#B�h�)F8M!�$�"��m+�灂X :�v��%]A!��$*�l��a��豂!��>�!�$I�	& $�_9mɘ��B��7�!� �w���Bw
Nx�nlڱ��*N�� �HON#<�2���OV`K&�H0%9"���c�<� n�ڀ�Q�I$�@�+Vu���E"O� )�L�B����$?�:�s�"O`�k�KS�����?)����"O��!d��09N� dBU�6���D"O|�X$	ܠ�ˣ W�
l�@�'��O�)Ӷ��!D�a*���b��y�r"OԵ��[�� #	�r���2�Ix����փ��)J�� 	�	����4x�!�2O2Nh��ǛL��C� k0�����I8p�13".ԥ'�����W��C�I0%�^Y�b+�,���c3�
5�k 9��hOf�q�;8˸�3F��&�l�9��'����<A��tcT]9$�<Z�.
Y�<�P(���� PCI�	/�i#�&�R�<�0��E����шz��Ec"��d�<Y�X*b��u��< ���/^<a��[��9�a^�j����BX�6T�=�9Q��\�JԚ�{t�>_����I�HO���-�dY�HJ��/ZD���"O^�K#��$,�jaR�
Q�3��(�>����	�GEٹ �	�4��t�C�Q|!��90�#B�6��3u�U�!�Ą7"^��bލxU#�`��j�!�䏁[��M�PlЩF�Բ҆�z!�D=M��Dbm�(jʔ�Fc[�[�!��|�Xa"�$SȎP3Q�̕W�!�dve��k!G	,��lA��!C�!�䖀�u����X�n�  ��!�$J G����	L2#�p=E�ٗd�!�K-"YtA!���5�������^�!����5PC������w � }�!�	9Ih��;�&W1lв���N@�\�џ4G�$%ժ}�H�.ۯVK2d`"��yB�75�� �5�b�#B��(�y�B]��&0ʶ��8UZ�ΐ�y��N}x�\9���zMh@H�h�yr�8@H���p��raP��D-٦�y��V���(qD�7j���Ǆ	�y�kǽԶ}�M�/[崜��+N��ynG9Nw,p�Qa |��kSb��y")�1\�h��^.%��AB��U��y��4;R`�'M����n��x!��^�G�a���8`Ducnݥ)^!���I�xЈE7��(@�X53E!�$̖`^j�+�f�$b��ٷ��7�!�DR(:mh�
��@�p_���Đl$!�D;]�@�x�玓rN�و")K�e!��!ƈ	�%�_T��	I��$!�D�f���	R�1C�PӃ�9�!�Dƣ���hw'h��6�_�>�!�D�0Q��-#u��oX��WOȀ)�!�B�Ta<�"F�+vZ�S�N��o!�K2r�ȭ#d�͖"]���f.�[!�D���N��t��3�֍pe��.~q!�D
2ZQ�|:� [ h��8(�
�!�$�2%�z`b��KN� �
�?f!�hw�A 3eӄ^���2����>�2�!CcU�1���@e[B��l%4]��m�+�9ٕ�_����G��Q�a�	�̐%%�Pt��T��;&@�(E7|l@�͌x�
$�ȓE�1�!���z�����D�����{\�PY�d]�����_"@���hm�@,1b!�ű#�?����S�? ~���dn�c K-��ۡ"O9Wa�+A�H�A�O�.���A"O6=�D�``��\�f���"OX�a$+��q�ϒ*s�ధ"O�T�����pJ.苒O�5�؀�&"O��C�k;'��9xGO���J�{�"O����$&���X	ym 0X"Ov�P�Ĕ�(�n�"��N�'aR�[�"O3�.�KB��ó ��eN��8�"O��6*O�JOb5�bR=5���"O�%�#eN�f�6<�Jw��HB�"O�����> -;r@G>�,4��"O�M��-�2.�*�⠑I$>a��"OyA��� ��U"�@�H3"OR�! ���L��u\�(\Д"O��#t'U/1�.L"U�����y��N�
�P���=\R ��Q8�yb���Hz�!@�� \�];7.T��yRF()��� �!�< z�"W�E%�y�7o�֍)��.�މ�m�/�y��'<�ƫ�/:�^d(�$Z�y��E�ZG��S�h�5/E`�����y���	e���(s�P#TRLxI�`Ƒ�y�H�7p�F�9����[�d��g���y���{�:�X��'%�ȩh���yb�ĭEȰ-z��M� }(�"�\��y"+!n����J��l9����yB�G7.5�ak4��36���s�Ƅ�y� U$>h&��g��,=Z��"b3�y�"�(�X�����PkR�!р���y���Hv�`����F�A�?�yRG"O�D�"R؁q��˫�yr��s!���b$L�n������yI�'�d,{B��I)���yB,�/*jj�K���^1�D���y"�I#0���(���3R82P�S�y�%�FN��b�� u����.�$�y�EP� n���w�؞k:�Z�k�5�y҅�m@�**G�d��4;s�:��<)�򤑛*�ڱ`��;�nL�w���6�!��Z���	�U�ԓ��zu�
x�!�p���� L��*:��t䄀C�!���4��X7*Nl&���Tꜘp�!�x���i%͖H�\��IΕ�!�$��.�~0��'��-fyHr�,wqOJ��ȟ|(��WR��u�?/H�PP0"O�=�6�ЪI���Cp��eJ�fS!�d_65j�]haO�-oapp�T�!�䄘�l!��$8��Ԃ�H�:D�6
OPM��e���={���fX�x��'cqO$�s�o�2|�D�bh@*BH�
�"O8�/NBR`d�4��I(%�]�<�H>��AH �h�4i*BQH%.�?%-����I���D�]����><�D�W\�Z�!��Gc�fy�R*�)J����W�!�$��xD��O
�n��a��=��	p�������ՓQ|n��1LD�Y�D��b�d;���d��DP�@jI�ya�qh��ùs�1O2��đ�BΉ���$� �Е��3|*X��' �a8t���R�X����;���BǓ�~��Ts[��ǆ�.K��y���X�Q��1w��9'Mb��'�M�8�j�* ��r�!�d�=��C�o��0�^yCt�$����d���"~��J���8Sa���8vq�r��b�<� lAx�J �f%��N�)O�̣��O�6��O���ǰ�vD2�a�SE�����T�-@�'����	f�S�'OK�ա��P�^<\a�dC��_a�|���y�23�D�蓭!��*׶��'����"�DN�L������-TS�\��!�dM8r�cƑ�d>�x����o��؆��%G`f-:�&b�zT���\r�|B��@�ZY`V���M���E�]�BB�4N���q� �D9j�b��_��c���ӓ�P<ZUH VԂ�g�% ԅƓd6� �Ո��YVtlzt�9XL�5�
�'��	z�Mޣ>���BD��8y�j���M�(Ov� ���x����wc^0@«�7Q�<�%�\�ߓ?��}�p��vJ.@���.��aE}�<ObY�<)�'M���a�׿cԽP�H@�EŇȓ�l�#�+SjJq�#e��
hA�Op��>ٍ�	�a��	�T(n��Ć_�\�!�զ	u�!�1k��j���c5�����C�ɿj�@B�a�+aF��[!��$!�*�>���%t���Ic�j�f�av�Y�s�!��ۥQa!���
*9G&�[��3��6?�O<E�D�~�`�@M� �xUp���7�y���6js,`��gC�#(x���N�HO���D��3H��:�L�&$5��	P+ڷL�!��:�(�[���)D��h��j��U؛��	���E�T��	��h�ˉ�)�
ur�L���'�O�-�|���=��J"IیL�r}1�!�Z�<I@dq���8�+��P|�T!{�<���N�@41�J�-7�� xF�t�<	��Y�C���3t�*i�x�!dd��t�'ݱ�(�hd�ƌd�<�W*ڵ�`��"Oʅ���?��M��擵c��Hڔ"O��Ωi�f ��]s���u"O����!C8o���Z��Z�K,�i*�"O�hQ��#{n>qI�·o1�}I�
O�7���J��@�B �A�	E��C3��v���I�A�j<��S��t��iɟ1#=�OF�2�S�|��0E�޽z��q�"�ێP:�C�I<&��l���]�H� ��eE Fk�6�8��9?E�ܴA��+` ]���{4A�g�����((���+��4YD-��)��D{��'�ҥ� ������p`O9��A�'^j�@F�L�T�t�PGl��}|  R���xrA+�� @��H7n�� ;��)�ybK�
�8���X�"���l
��Px"�iU>Us֮X�)p��i�ȣe1B$9�'Y�
�%�|I�Q��Ꮑ8�y򊅈|\>(�f�W<z�� Nˑ�y̛ W�~	�Q� PݻGb�Ű>�M��A�6��dJ�l��^��U맃�<I����xT����B�4-��`�԰Ez"�~*�P�j�ʘ�4
ل�F��RFL����?������} qN��O ܪJ�K�<y� �i�.�	�[
)��}bw��S�<��U�NR�q����Y" �Z�<��Ĵ��̪g��^7x�A��S�<�1i�$I�o>���d��Y�<B얓NT�- w��?;��pC�P�<�0�8IW��bk��zR�=J�DIT�<!��3(�����Ď�Jp��a��k�<Y3���<�ڂ�N;4D����B�i�<��l��X�aA78�R�;懚^�<q%��T�:*����H߯k�ą�K�T��əe�xc�#R-Q�}�Cm��7˓�p=1�O� �LAaH�� pz��ӭ��)�V�K�"ObD�+���1�F�� `�+�"OZTcPF#x��xxkO6ͬ����Ob��$�	c�'��i�"8�vH���F �Y��D&}2�I
���u"r*��k���@�&S�!�D�_���'�U��!��
��-l�@~b�xJ?�HA*M�
��>pD��7�ڥm����ȓ��`�v�S�hd UZd�[��ZL%����	�6�������-�TZ�h�PҼB�I  ���!7CL�:�8;q.�:Ya�B�	6֦pk��>1�RMP�N[��$F{J~zPL��y�ϗ�R��X	��SS�<�!����Y�6@��I���g�'ay�䞄>��'�n��0�D-�y����&A����6��aI�̔�yB���p�y(G�,��@�I��<9��D�0#b�TS4�L<�3B�w!�D�S������&tEt�f��!�Ā�y�r\"�+ܝ(2>�阡�!�dZU$^1#�9$d@ �F�5j�r3O��S!��n4��Y"��"0�7O>�n9Q�N�j&�ǔv�j)��-�N��B䉖L�"�A�Z4�<aJ+�4S��B�If����O(]���*�TB䉸CB�Z��N.I%�p�� ��Z��B�($H�M�t`ZP���1w�-v��B�I�N�^=c�əi	�H���5eE�B�	�=�j V�C�[�14m � �B�	V4H�����3&�>G��-���)D��qW�~�؁�q =Y��Ā(D��ٷd�&��$ �&Qh��DH+D��[䎌�Wp��J")�"�*D���b�N��7$ȐG}���	~�D���"g"�e��x�.9� @M�q���$�%�� �lX�AJ�7kt��`Ζ #�]��/tX�3�A�)��ˆ�T�̅��Ge�Q��@�"
ԃVE+oiX���9��L��C���3g � &�H�ȓi"��� *0S��Yn�P��|��x����/��(|"��m�+���ȓB3�d�p
Z"m��Ҥ��i��ȓ-�0L�eN�Y7�m��ām�@͆ȓs�,�rf/%-^�y�EXQ��m����mi��f���sjT�^�vE�ȓi���A�
a|�ЋRe�T�݅ȓ&�4��o !j�h�cga �FՅȓ�$|�U��>�V�� OY���ȓ8�xhˍD5B�c"c��7Pl���Sf���A��X�T�V;�y��<��òFT�K���kEmP�ȓrD=�0ak���G,1
-��"OI�F�^�C",0��L�N8�iD"O�lQ�@�)3����W#;.0Q�"Od0£�� +����2�J�l����"O���a�Ǳ(��=B� �-
�$�r"O*��E��[\m��� ]��Б"O���K�Qm��8w�æh�4a�V"O���,���M�/X�4�R�(�"OrI�aaԔP.@:����r�F0
A"O�]qԉA�X�BhzG͝=\�t��"O*��w!�j�r�aT�'?F\�"O	hޑD6T�A2۫Ma�!�"O����/W��:��4��j�"O6����@\�\������0"O� ���c��W�<i���Q�.�f(P�"OB}[��ܰ^�<�c�* <8�v"O
$` ����|c���0�t"O�sS�P��[�� �>MS"O�QS��۰��i���O�qm��0�"Ox���H1[��9@lxF�c"O��ڢ�A)�0�+1)D@)��%"OLa�i�z7��p\L���E���D�>Gn�r5%��!(��	I��`!AW�n�*dힲmSC�ɠNF����@�9rd|�v�߬dp�B�	-lrL�hDÌ39����"w�B�I>ir�1BX,]�p�!V�O��B�ɫ(9��R�յq�J81��֊bB�I��r	�p*�LZ�s�.�H)�C�ɘG|�H��f�1;��h�'�$�bC�	�+��1�Ț!�n܁㜫G�JC�ɜx����/O/B�&p�t-�8�RC䉂+���t̏�2�����`�6C�	�[�:�B�!9� ���	��C䉃�nh���Z 7���'q��B䉠@}4�6O�z
4���oB-\9C�I�	�|�ڂ���QQ�P���A�H��B�I,Y�L����)�l�WJ�;6��B�I2f~y��y�j�Z�B[=��B��6�����e�,aDF��̊�#tB�?B�2�1S��0$ӧꗤKJB�ɕ��=�P	�D� ��ΔB�I�]j$rAb�Q��b���S�B�Ih]�{�)�#P¾1��@
.�C䉞
��d��%�\��p U��C䉨*渡��nW�e���+\6sY2C����	���N`��YF��n>
C�I�/8 �%�G�~�$�`!Z�"��B�	J�}0�C�xPV� S@�i�B�	�4j�|�U����Fف!��3;�C�Iz� 9����_��0����:C�0=~�q��E�*Β��,nB�B�I?0ߚ�Ӳ�/o�H5z�c�->�PC��'Kxh|�g�֮�&Y�̇�[hXC�+5���K#��o�L�����WuC�	'Zt`�vo�,I
��F΂�S��B��9BT�� BN��=H ����\�B�IqH����0/�@�@mݾ1�C�v0����������p���7.�B�	���I�ki�X���z'�B�I�n}NѨa�ӂ//����k!�B�	8&�"���߁�P�6χ>?jB�	\]tU�q�3o�R�!�+z��B�I�*����-�q�d\*'��ޤ����H��2M`"lb� ��\&B�aD�F!�dǁ4�̈{w��W8q��C���Ob`�a �N�O����Eʘ�,��"�#��mY�'�R�q�,7�
m�f�߽�Z�a
�T� c��A��Y�,��oռl฼f���4�$�u��Z��#kA���y�g�yؤ��I�*b�9���x9Zto��W�"ye,\O���F�(]�֡�0&A+8�Q�CԽ1t���5�ݻf"?�Ѭ�\���'H�	�DT�-
eN�f(zPp��d �(��q���Ъv0�<�O�̩%���!z�y7Bߔ7��mp�}"EM�bRYX��	V8Wf����`�JL&4�d6����5Lx2�ᘿ%t��'"۾P�t-+M~�$CbC�%)u���-KK�$��ė>���O�I�)�_Enl��FO���=TN�]��I�4}���lأ��g��`w�_���y�
˵E��ϓvE���@�_N���?����)*6�뀀�6r��!�ٶ���� �Һ�}˓l,�գ�aY'v ��!�ܱ{T(���憐&�pqI�o;���Â��1=� 1N?� Pq�� ��5#���\�$k��2uqFM�s@[�>]#�B=C,���Ț�TuvU�>q���A�0��3�ȩ3�a�T�� T`��*D��x�0Q�����.wOL�I�"~�Ɇ=	���I�(WR���@�2��yȃP�TX�� j�t:O|�>S(�%b���P2F�/G�l�Ňp?�D�E4�j��?��a`�D�߰v���1���I��gfX Q�K��?<O��X�&�%Z�S��̢�:�g�V
x>�<�AZ��0<Q�I�>"�V��I>1��ǫ%Xn�x�¥}��U�S��Q�'�2	�m*&_d�D�o��~�R�/�L�v��Ei7�yF��Mr`�9d��CӲh�$�J�M����,?�D�H>E��4K+��`׫�,'*AL"6R���ȓ"׌`������B�q�f���:ϮQP���*1���GC5V�(��i�H1FK�2�D�`O��zq��V�`�C+�h=��K���.a�p �ȓcGdSŮ�#
4nH�'�
?�a�ȓn@&	�!���Vy3s%J�G��ȓl�h3�i��*D��K:/���ȓ!�b1����e6Z�"���r�8�ȓ#��
���, iږH1�U�*�O�:E%C�z�T����+�\���ɮr3|��3��Px��T1s�h�ԮW� �ï�hO��l\8X��˵a#擒I2i�ğ�*��5��\V`C�I�S�aC�GM��}0�ݑw,6-�n����);�*�3꧈���C�>!ѩd	��F_�)�g�;p�D���<A�X4x&n��&��V��U���B�Oj�ɦᇧS��}���8��O��t+�9	�<�b�J]�[������I�L��ϓZ��<��	�O�F�r"��u�L܋�s�N��0�U�$g
�?)oS�?��'��t��I�"��ˎ�2�4������|m��aV$΁K�M�M~�����>IF�	�)@ (�W̓+G[0�*�)�- ����l�r�D�X-fx"6 �w�&��#�_�|�� �����"քD̜������T�t�EjE�"lA�=9�b�A����Ձ,� ��)ހ��1���!jX�I^��-ؠ/�f�<�(��5��I��|���͍5pp�S��A���͉ī
���dE&�dPFǒ�ː-����1��r�(P�%��8t(Ó,~��O<)�E��JhTx"�SP-x���Y�'Ԥ`�B
+�ؼ"��Z'��O�N���C5�J�R'��q����
����E����Θ!!�� ���3I�9�4懽R�)��b��Rm�)*��H`z"|�'\"�g	���:�zR�X[�b��D�A.�H2���]>SgN��O�pX�&���v"&0k�+U1w�@��J��h~0@�'|xj �րy�z�;���/�F$#�G��`�'�G���Ia��4pZ��E�ދb�*���`���h ���B6�G�{!�D:?��LYGᎧ�B=����(�����+�"�ل�(D��(te2quə��OH-���F`����?��Q�˛(\&��$lT��p=��],��T�� N6��C�Y-?��Q�n�K�b�-�1d�Y.8��a�.�D?qРo�{����Q&� uPx�dǎ>>W�L��H;��>?T�XɃ�[aڮh硅�Htq�n����X8?��<��$Y�,��(n���C�<E������N�8��}Pv���dv��YA� �.�V���ɟ�d�X}[&G8���>�@����0�?�� S^KhPs�ȑg�e�Pm�r�<����$�J�S��p�w����Z�M�J8��
\(X����D��=%�ݙ�)Sy����漨�O��0(B._�8��0`�E�?�TDx�8��$P�e�:�Lt%j�!Hи� +�q��ʳ7%ؔd��<�<I�R�����7�b>�.����JAh�@7�BpI$��P_x,��a �xU	�b�5ғ�,3#�Н!��M`2�-mj��	��idn���޺K��L��i�a�#,�h�+
�W�|ف���a<$a�!����Z%	7��'dq��R/�?!P���Qs ��3�r�j�{$ckh<�*�'X��h�I�*ް���4@��h�eo4V����QM�	q.2hC��'Y���PD�&H��r)"������I��T��A�"�'��E�q�U�Q��q��E� v͌�-L&����`��9ll �X�b�̜H2�!}b�¤c?�VQ��:��ڕUO�@��&	�O9֬�<���IL1Ą1��˭q�Eq�DHd�'�B��wi[�w(U�Q���79��I��RǢe��i��@�VŸh@�)R�C%�i���%$�;��� �.!#t߶-���8MBH�?n]�k��[�ܡ����#l?lՋu`���}�ȓ�4�S�Oܴ��ыw�� m���,S��uF�ƴw���R!���ld��)}�7�� >exp��0w�͠���&\�T���'2l�[�A��#Ҵ ��A��&��`������ �5d^v�I"AZ	 Gެ�I��(��w�g}�G%Og
��E�<tE�XX�J ��'R�2B(!�6�	`�C���O�|�d��)7�6�)�ӧGJ�Xٴ���ZfS�9�F��DH�*3�a�֏�4n���@�H�8�rCi��@��ɻ>�H|��	�=&����O��dH^'%���ؘ!��0�"Oʐ��U*UG��[
������?OR�BU��9D��H�h*��{�fJ�����	�Qi,�3��%?�dYV�Մ*�a}��J+	T�e*�4W�xq�#H�y���q�U8)vP[%m�6==�,�O�谎�Y��BF�ّ^��؋:_�Т�"D���� ��b�X�R�]na�T���O���*E�"g����іk&( &��Xp�E� a|���)D�m��c��ϫw�l�:���$͇�I;U2j$�l����!0��;�KZa~��8�=D�p�'����к��56�4�s�!�Dǟ6>� ��{��tJ�cք�B�߶�D�;��P���пl!Ёzד$:PD�P�� j:%�1��fӌms��̲lɢ�?�I֍5&>T@�t���q���A���#��� �qh<yS�ϚS�,�[�ҩ^��yR���d��a�H2�e���Y��R�d���caљ ��k�W7M��9C�'��3��Y��	[`���Ǎ��B��aɷ .66ML�<��BtBC���)���8�̀"IR� �kGJ�p�2�� �DG�I�~�:�{��(��"�ȍ�����'���$��p��f��<q�H�I��H1o��0t�aЕ���'�����4�/`����OH�u��4!�zh�0#M$?3D���8<���iށSYe�&� ��Fz�o�����DO@i��UQP��c"�D�����+q�X�ȓ i�mͪ> XX*�N�+�Il�"+��	u�
Ig�S��M�R��2+~�����YQ�qSS
�G�<q�k��CB噠=N����C}r X)�
�A�`�Nx��G&�8fХ��+��H��� �!�O���PN��sf��
C���H+�̀���&d�P��*D��򶌄F�������z� ���<�Vܒ� ��<�'���A0��!����C��O\����:���KE0i�a�"����2�ȓ5Y��0�o�5Z�-IRo�8\�5�ȓg�r @�J7�\0b�Q�����ȓf��
��Rp ��B\mdA��piH �o�I2 �� �TmZ��ȓkfܼ��79��Y�D�39�"��ȓ�d�[�g�OY���r&�~�p�ȓ;�����#%b� *����u��9��?�nt4�7h#�QQ��i�>���];8��t�R���r֭Ѝ��!��Ɣ��hBcR�	�\|��FrD�����sH�"��D�P����A�l`9R.	�L�
�qq�ƬX��J,ܜ	"�Ò2��H�������ȓ,!���0H��l�t�0b3DZه�A�<��_�Cz����)��5T��ȓa���X���/~�&Y�����ȓ�U��f��<��҂N6,{.�ȓ|��t+�G��~�����F�8
|���+������	�j=�%��8=N؄ȓ[J`9r�E֛w,��ӷ��p���|ڜiS�l1D�8)j6�]<]����C��`� ]�~� C���p��fu��fEN$���"P"!�����^ H+�
�Nd�m�tY�p��ȓb��=�¬�xPF�)C.��70���ȓ>�^ik�nҺ���be��9[�%��dZ��{��T� n��G0E���� ���u�v�Y+�
:|���V"Oh �Ӈ|�p���'U�bL�%"O� �H��L	_CJub%B�
{ԄHH�"O��I��<d]��Â��VMC�"OLx���Ɛ+��ȹ�LV�E���""O:�{U+��Ɯk���H��9��"O�X�&�4E�U	��v��� C"O�4`mI H4-�#艡<�p���"O`�P3�#	P<)���"dq�"O걚�ƈ�I�D1�PF:7�� "O��,m�D��1i��7����Z��yb&�e(.lyRD�$jH8�����yb�R�,Yr�8S��r�T�`�@�yro\6%K�а���F�Tp3M�3�yr$�-]<��o˰;��7啀3Q!�ޮ���g�[L�ʩ3C�2l!��5P���@./R����j!��ӽ<v,{�,�sS���4�"7]!��M�\"���Q UC�Y:�6]!� 
r�񣖃P8��a�L�E!�ǦOٸxcNC�@.:4��ֶ*!�L[�X�iga�<D����i
%h!򤘜</�8��ȭ8�N @���_!��$'�$����Bu�u!uiѹ�!���3XI�B�f`�i
�Q.�!�DS�q��"�m�bq4�Ӷc�	P!�H�PhIQW�0.H��s�ˠ"]!�Ğ}�h�*��2����G�0a?!�]U�E�NW�L�TTSa�
�K�!�$U8z�IS L�:<�0H�%�-4�!��+x�mCsk�s��h�.@�e�!�L?`)j#�Մ5y���CߍZ!��\̑h��DeN�;�ΦJ�!�D�,(=�)��T�d�l�k%��92y!�7Z���!R5q�dp@s�̍>f!���p(�QQ�Ɠ�M����t"f!��:aH`{"���-���w���!��	�#mp-z�'�9!�%��(Y�C�!�I;v,�Q��f�:\,� �(�!�$W�#&(QY���0�<���8�!�dA�G�	 ��.�L��$�~�!��D�&�y'�
�Ȁ����(�!�� oݸ�B'{���`��	�!�d��D/9cI�qfʽ��C
'5�!�C)(�X��%��m^䐙#"Z�b�!�ē4y?�-���3h��P"قq!�PŰ�HP
�w?Nl9���x}!򄃳	�X�y�/� ~�X) �U1/E!�d͹w\�㷂�r���#!�2h@HS0���i����fſ{�!��.&_����IsT��&�6A�!�d[c��%�Z9��œd�Oe!��3?3n9�0➴>�L|��&��t!��`&�-�@�t�Z��I!�U�!0�����(�"�s ��#!�dY�El��ț)�@Q���0<2!�D� GP�PnF#��l ���	�vB䉃L��E���<m��
�� �7L B�=%��R�(^���� �»d�HB�+j^�=B!��`�D���&�`�&�@�!�^'�dc>c�ԫ�K� X����ʕL��[7�6�On݋��O�)�<���گS�d�K��"(�~���OӁ��?���ʂ���!
,<�p|�u��f�'U8�h��R�l���~3�?.xmrɘ.����m^a�<�6��>m��ز&� �F�R�����d}�E4}|J6�Ǧ�&���^�r}Jxse���V%�b���Ǆ�0S�!�=E��� ���W��h#T�@(�(�e�G�(��dC 3�^��We�^�3���p��Y�
�9a���gO�1B��T5�1seߦ��O�<�����)��z7�ǔ"��ŨW��Y�F��B��#t�|���Ȗ5�
�XY��5�G�)o�<��4'֡vY>�z�o\R�'�De�$ᝤ?���ґ~z�dA�NYr)����_�� .T�'�h!S�KS|%F����#�T��٦�����P�����S�"�PG̮��<���D�@��d�6�S�m �
X� jDoŭM�� ��3}���'tP��*�:�yHV8�@yb�!ngV ��,��$�$[3�y��@O$F����&+q��"(
<dz��A���O��4ˆzeF�O���`��N�s#����=��<y����v$��w�Ժ%�Zb@è
���A�
"���B]�'$�?����QgmR�(
����t�Q� bg�Յ=��ܺq�0~��Y*�5s���ќkG�B�ɇ{Ps��Ak(�<[$��6-ϊc͜0HSM%��s�f��5�ΨF[���RM�Xat"O&%�(���HB��_�th�A"O0�Pl̕R���Cb�r(I�"O��*��0d�� ����&YȂȻs"O@QYW��6>\xP F�Y���s"O���2%F�%<�4�V�E�򔺔"O����d��_>Z����4�����"O���Q	�~��CMF28���"OT��	>іt�-�V�,L��"O�:��k����/>r�J�'@�HT>����lЄFX�("��D�-�L8K�#Oz(<!��;H�����
#:���h���~�'�̽���#ൣ�󉛜C���0m�1.b��4��6j�!��J��9+�i��s��e@���)X�V��1d"4��T�MR��S��M[�>���@��qlp�2	�Y�<a�I�x=� Ƅ�sPų�$��~�k�5,��#j7"��0E�a��Uق��4|@�8�&� Ȱ>�!n��$D��O���q6o�*vm�٘�D�(05�h��,�O\�3m�2���Ø8�L]���ɍ)���vFO�MN��A�����%��H[��h��dDԱ�yb�̰uڱ����	ä�I�h��sG���H��K6���s�ܠ��"E�(���2�*,D<;�"O��������З�#Q�%���{�HQ���xC�R�%\�+<��?х�ÃP�ec���9��a�K�I��	���1]�@���0'��ۅ$&�T4�G�K�[ ;#�Z{��LPW��s�B���ㅪG|L9d=(㌌� ��X�BuχĶ��H�R�Y���@�@0"���ȓt�����ڌ7/�4b��2H��mZh״�@�B� T*�)��<�v/͆&w��iC#�=\����-T�<���ɥ(%J̉�)�C���a�B�<�BD�^�
��)/\O�}��A�2sƒ�P`�\�<��e1&�'�(��׬�2�4L����� X�p���w�da�`Ѽ�y�K
9U��B����nt��S���O%A�w��)؍�)�,K\�|��E�Y�"!k���`!�ĒN/+)J7�3AA>F:ŻD!S�8�l[�A.}��9On���K
�=f.	f���H�@��"OP$��6Z�%ȣ�>t-3Q�'�p�e>���.J�ޙ���
~���S�nO,T����Խ|,���*ݐ�?qW&	�iJ����;2�9�mKR�<AG�n�����o��#E�M�F�D`�C7t��}�i�1��P󷤓X�b B.�M�<�s��WD9�Ão����`�:��A�Х����I��H���>S~��6Fɾ!�:��WJ�kB䉓y4�)��ô0�&A� �m|�7͆�3�HL���%��=�e������ �ev����A؞�D�ͭ8?4���''�q�p��2Wm������،C�'�"0���\�ș��hӁf�`4�}R �#G��ˠ,�@�O��#uM!=��\�5lW'RKt�
�'��#1�?RцY�t׻W��qIP�D��3�>1��>aRI3&n��j� �!S��(�V`NI�<� ,�#&N�LQ�\����x-�8�'�!�D̔I�a|���A��)����r�u�S��=��� ��e"� �O.�bL�+Jasa��dа�%"OF8
�c�J�.�z����U�(;��$�0�Z�Ka蘏�h�ƽ[f�W��Y��]��z C�"Oq��?H�P��T�z�� HQA�fp��0}"�0�g}�-�yt`��O�h�9��y��JI���p���h���
A%�M#�ɵSЪB4|O����7$� T:3��pѰ1ʄ�'e���Ю5C�ڤ�	 �3�H�i_(iQ��Fk5lB�	4�n5����&!D��"�żn�(b��IQ��"r����퓻[^ܙ��0=8<�"rͅ�F�2B䉥E ^4��ˀ?"J�ˇo? rMjt�"���O�F��O ���_za���-��H�"O���&)A%{O:+V��:E�-:��'�D��C�ca|bߖ7g���WH�
�㵌U��0>I�(��d���	�$;4��G#�$gԢ���/T�qupB�	>,�ԣ���*5R1I0m��*�fB�I7CK��÷�é=�T�Ò�^B�	/Kn���`=O��I�R�@b��z�j��f	.\Oؕ"gcȇI���6.����]aE�'��MI%](s7r�XP�ʨQ��$kЍ�X�Laڠ"O�"FU6T媝Q�ƈ*�����v�H)��[�s��y󏑮s���)w/�� ��|�"O�5�k^�K	�0�P�L4PИ�c�i;h�K�i@���O?7�H�3�hM�Ն�)*�Z5�V��eP!������q� BC���&�W��	��(j��L���yr�-%�9���6BCTe��$ܰ��>�0ɺg����d�	?�,p ���� ���U�B㉱u�ɋ�+ƽUY��b�&Χ:�"=�� X�p����E�>�S4L��e��!a���=i3����y�	ۓ'��))�9 �I����Mk�d׃1�6�'@ }���i�6u�&)� ,8��`��V3&��,��'L`Ha��ѓ<�,%���S�DMjگO��i���}��-b
�Ys��f�v:L�c�A0o�V���	0n�\��u ���#%�} ��IH3Xn(�ȓ���k��&"��C�Ŭy�̥E|��VxoVDF�t�J�f����B�U͊���/��y�'M4�NYJ�ڱD�	K���y��l��i��S
H��Y��y"���:ȳ��ҷy�@�Y�Y��y2�[�j[�!�c�M;z;�j&�1�y� �9���h(^$�2k���yB%C�G�L�13��wk0U�$�S�yrb�G��Xf�!uG\h��g��y�؉Pj$r6�>���Ö4�yA��a�rP����7�*��6�y��B8t�A 6Q��D��n�yB!R�r� %DI�^4�kL7�yR���
Y	5��<M��!� �ؿ�y2͛�:�=8��a�-FXVB�ɗL�`��A�>f�;s��{��B�I�Ġ�d\�|D2��P	�}�B��/cB����#���8b���:C��_1f�� J��K]�)�G��=@C�Ƀ�D���^�x�+�I
(�^<*�'C�yS���;�U��ѽ'm=K�'��� �MЬEz��zI�'��4�
�'�j�'�54	��c�.N��	�'��"��_Iruz��l���'9RpK� O�L+l����
�' d����5�U��*]9q�hA�
�'P`=�d�6VD0���
n��	�'((�p��Y7d
�����4�$���� ��k��8y����m]
e�0B"O�� �H�<z� �:eٸ �@��"O@�A׋�9n�p�d�Z�N,x{&"O`�p���
�l`0�ʊz���"Ov�j�%�v� b�ZЬ0X�"O8��-�:{�X=h�	��d�Ʊ;�"O@!ʰgL�&�.y:�hȄQX�q&"O�h+s�	�	��*��;U8��"O�0�A��h�����c��4��8�T"O��A0n�
}'�ᶡҍb���H!"O]���}\4u��`�E�,��"O���#�7[��nR�4�ЬYf"O�7(
*w,:Ē [`�� #3"O���� �R����%��;D�s"O��@Bdܝ1\�����=��[�"O�e��ұy��<�d$Ӿk���{��۵�<%�7,0IH.�˦���p���I?ax��ɾ�M�$�'�F��v�� 2��\�0̉�(7����&�S�d
L)=IB�Bs&\�Vw��)KǪ��'vўb>�ӕAM� ߖt!'@ �JPc -?���Ӭs�<9zP-`�tq`��A
���c����̼�C��Lc��@1@�Ra~���匛��'��ç9"l�sC	�jǔ]�#�X�+D���=��4+E��Dxʟt@��ǿp$n��d^�L���ƙ|r/?M�Oq��y0T�[;&\i׫ìi�0D[�:OBq��C�զq$��g�beT�W�U��|���o�"�"���hOQ>��cǏ��Z]Vv�%�C�0t�P	�' �]k���5<���0�CH*LuF��'�xS�H_�g�*�eH�GQĐ��7�S�O���[f��HfY%��@���X�O�Ⱥ�OĢ=�O�PI���J���3���!6�İ(J<	w(��HO�Oh�1ዳ� ���΂mح:#�>)�����o<�:F$X�%Tv����=5!�:t�`��TbE %6B�*��N�_��'Kn�Dy���+@h�+� Z�F�y�¶<���<�|��'�|Q����3y؀�`�Ơ�%��4/K��O$%B�I�A��M/|�xQ��B����L9b���I<��U����S�i��h��	�+� h�G�Z#cit˓T>��q��?Qc,O�H�bE��L�Kp��,bd���'W�=W�j����O0H��=���E�@!RtX��J,S��'�Jm�A@.*�"H!�O�����zTP���T59�����j��<�R�A�.JQ�s��h���L����M�$�*НW
���ȓNDF�3�,[�<��&��0�,��J[�tX�d�K%���8xvɅ�I��gN�ML�`��0g_�Y�ȓKO 	����p��!ĭ(�L�ȓAI�T0 ����#2eʥ}R�h�ȓk�*�s�AI4W��㵥�$YR�D��V�u:Q͌�@�>4J������A�ȓa]�,��hX"u�T�It
��N��S���X#��:j���p���T{��c0jƸN�l���*f�ȓ��e��)��%Z����@��BK���ȓ8Vxq�'�P�D��`㜩A�+"O\PTN�5w�L�k���t.�C0"O��N�yM�R�.Q�/[���"O����߇^�t	�m��G�`�I�"O���ǏׄS68���Kd�0��@"OH��匸b�4xAd@�`؀se"O�������pC�rAƣC4\˕"O8�C�%Z�F�sjZ�;�� �y¬ڑa�x �t�6b���A��S��yBO޶yZ4�'�R%qׄ|�d�y�&֜-/x4���U�gJ���$gT#�y2Ŗ7�&�X�oEf�Jܲ4Lܓ�y
� p�x�6Ө�X�JO$*��<Qt"O|{L���I"uIߠwN��2"O>}���>%O�[d)o� ��"O��J��fR��W�̔jl���"O\����)x]�Zfg�"FZ�D
@"O�-�F W%G8�T�$�	�tGH�R�"O`:��B�@��<���>	��h��"O����?����E�}��S"O�	�C��hS����Gl ���"O��+�9�ZE
�nMt�,�*s"O�|A�,��\ Y�*A@�8q�s"O,k7D�<s2���Iݳxq;�"O������zW�0QgIΜd��$"O<h2�F�����呥+Rq"�"O@H���BP���nǅ+�MY�"O@6��'`�(�1�(U���Q"O�@�eƓ�s����M�G�dmѓ"O�y:�C��$M�l�l���k"O��J��*Zf�b�����V"O��ۇ�ԨJ�2�ʒ�>�~��"O���	>Gr(��!�4	p"O�Ѧ�B&8@Ta0ïH��7"O�x���Z7[F�Q���t_���c"O���f��D ��G��g`��@�"O4=���X�$$ܻD��8`H�H"O��k�%W#e�:-��Kɗr�28y�"O�-!ႄ9�I �dʭ&�x��P"Ory0�
RB��J�MK��g"OvX	2�E��yY��vA��c"O|�0"R���$W[ڬt"OdAej��s�h$��#�
_���"Of���Y99�8��c�A��1�"O��A�S,9bP�81(�UJl�2"ObQ{ %�-;��Xg'ڼTVl%�"O����ia��!Q�F��g�4��"O<5�ǅ>#``�cf� 9W܀0�"O�ڶ�^�6߲5��[�-�U�E"OtB̖�V�1�H�r��ҁ"Ov��
�*��3�[:fe�Q"O���@
ݾb=��0v�ؖ����"O.��c�[H@�H�J⠱��"O�Q�4�21�G��(�(p��"O0*�,_��!p�#�	SH�;d"O<��@�F��y���I0@�c'"O�g$]YF^Ea��V�lmh�"O��.U��isp�Q�
�@Y�3���y"�+����P�ZyK"��1^��Y�ȓ 2n�"�ڐ�8�D��{C�9�ȓ��b��(_�`AmT=n;B�ȓ�2<xu�X,ń���Ӽ6e���
Q�5�w�+]ۺlۣ��bQֽ��/ ��Y���/Fу�,��$��ф�P���yb�BgA.$ɠ�:C���ȓmb�=����"A�<I4J�#�����x�V�Bb���r����o�1c&���i�Y�
CX���(�h�7eBE��H��H@�_Y���bA��p���%�%��Bߔ^ <ݠ�� 	B�h����i0��>+hZp��f���`��lj!�<Q��,��_ld��O������9=r�6nXwDP�
�'^u����1P Aj4d�!��0�
�'�L����3��|���-#T!�'F� ��G��>E k�&�4@0[��� 6ESoJ@����`��j8��"O>M0��LP�̎e
�႑"OP:�`<*{�07*��:�$��"O�}pD������K��+�i۱"OP�J��S0�։qk�R�>Q�"OR}�fn�m��Tk@T�Z��r"Oh\�pD�wp���R�/0\�U"O�(��h�!}e� ��'�t�"O�+R�P�9�*���;P���[p"O$ؐEπJ�;Cn��h*��{�"O�x�p�V�p��tgD!<&�"�"O��6O�*�]u�;'�-b"Oڈ�",ߜm�
DH��H�4 �u"OJl
d�\<*%���i^|@��"O���B F:��s�a�!	]�	�"O���թ��r�BU��AL6N\>y��"O.�d�����|�t��Z �a@"O�\�Q� 1�g�:Ԭ̈")D���Bj��"�Ľ���^i�z�`p�'D��s+�]�ڭ��!Q v4R�+�&D�`a!˰P�@�3A�i�%���$D�HH��Sl� �a7Y��RR�/D�,ZS��,X�h�xal	,\�*�
!D�H2᠊%J�����ӐEe��3�� D�$�3@�U9�ĐM�q��2D�Ԙ��;>� �U��Qn�I�g;D�8A��,��3ϛ�y6DA�Ն-D�xiv�����Ř�H&3���ȗ''D�d�䧓<I��X*W͉#���+C)D��2�䏻c��lSQgܛ"�Ը��$(D���ڏ[2B���DN�Z7~Q c "D�`�e�H!G^zh��bʦ&˨Թ��5D���AET�8���JҨ��k�0p���y"��)q���Co�:GZ�)�l��y�'r�	X��S����6N��y"�Xt8A5�@öj��y"!U�Lk*=��ݝ ���q�/�(�yR�C`��)��X^H:����ylʓQK���!�_6�*��C��yZE�"d�P��=~y�I`@��3RqHB�I�&�j�R�& f@�T��#� C�	�D(�%�ב��,���	k��B��!,$�𹤍Y/Q<ĨSB �.�C�	
&)b'��>}\	r��:I�B�I$�`���(ʕ>ON��'��B䉡C�=T瞎@�11&��e��B��Q�8ВvH�@���Ũj��C�	�c�6�Pc�;�.�$C�&j�����E��Ce Æ`��C��zr����;Ǩ�������*B�Ʌda`��a�A�`�<-���٩Y�B��Fv��wE�WPج��H�3ҠC�	�l�p��J�)c�a���[�(4��&���� �rʴ�X1I������*�>,���'8R6�8P]�}͒m��jm���aַr~l����15���ȓ�59Bm��m����z24цȓ)��y`�j�+R���q�%r"Շ�UA^I��Ȗ6]�=�A��F4�D��0�,���	Rҡ���ǧv@�ȓB4`Jw��!U�}�/�Ne`Q�ȓ9'��2lB�IՒ�	��B+|��ȓM� 1�C��"�m�Ɖ̌�FL�ȓ�v�s�m��(�4�@sB�YL(H��S�? ��S�
8�h"��� v���"OZ�����(1��ŰmS����"O���8I�z�`E�5�0px�"O����R��� �`�@ܲ`�P"O����,2-N�qR`�B �!�U��¤����R� �����>B�!�A�i��-1���Ntn��"�HQ�!���B�T��%�9:�P w��X}!�d߷9�6�2G��?nH��o\#K!��./D���>?��u:�a(]�!�$`��Qc�%^���� �<h�!򤖯\z%��"7l�Xk��4�!��

]�H��!۬�jɸ�gMn}!���(B�����*D*��K��C�bT!�є{�$����0�e���M�!��8n$�bԴ.z��P��V9�!�Ā)?fZ(�g��)k@����/.!���L{��+LS8IA1�V�Q�!�?N�*���`��WK���&H��,�!�j�B��	p�꠺��P�6!�"a�ԩ`��x�a&D,a0!�	+e�`a(�W�.U:e0d�� !�Ā�B%�%#V2%X��㝳!򄕟����»̍���7u�!��>i�>��dR)M�X�
���&�!�$�.`�(K�O.o�"��@>@�!�ΰ<9-{���V���)���!�$�R������çѬL�cn�'0!�$T(Q
m	VE��+��U�fL�#�!�[$l��"1�ΥP�DJfI���!�"t6�H'�ƑTU�	�2���/�!�|�}���xQf�x��L��!�;:j�HFB��kl:T�S�I3�PyR�9M�d=�BB �)����yҫ�=_��\җ����T��E��yr䖇Jvt@bB�C>���&)0�yb�طZ�:���E��"�X�H��yrJ���N4�6��"/��d���yĄ�*�>�B�k�(5`�� C �y�j�-����c@���@�A2熑�y2*�nh\��jI����p ��yB-�
;�qb@k�/�"�鐏-�yb+5G� lq��2���0ϑ�y"ڻ_���D.�[�
=r����y�
߻F4l+
�;RBLi���$�y"�'��(����֧��D��0���|.d�3B�[�V�4���H��V�#W4��ը3b���"���) Y"CЋ}����rL��7.�H*�eX�`�ZL�S^���Rc]���Zր�b^t*2��#6��X1ܫfH�S�ko>Py�5d����mJ��lr�4�	�M��B:�d���fSt@6��I�|U�#�ְ�铲?)J>����'R��)�6x�d#��&l�P��$������4�?�@�i{����U
�A`�9RM�3��e�6h�ӟ�'ܢ�3wdzӄ"?��C�-�� �!I��ȵ��E�O=& �1��'�nd[�Q�Y��t�������2�|u�'�����ƥF:��#�(^��D@�ʀ�^^���'e��`4���&oɗ|��'���j&m����NôC��yp ��7a���f�3x4��)O�E��'&f6M9&��N�!5����@�$,���ab�"sQ��ش�Q>;%_�n
Pք��O<a𨸟�K�4Gu�F�'�H7��|�'���*��m�t䉘T�ч,�5)Ɛ�[e��Ԧ��	؟$q���"��=���@7]�q��	.�k��;a��&F!Y>�HY�<�Fyr���N�  �c�?w0Z���V�t/R�e:����`P&Q#F'D7 �"�����e�K�ؘl�9��9P�鏊B<m��'��xt�i�O�d�O����cG�.dFı�Q�{�TT��YT�����@J�Oμ�㤥��B���#�L����	��M�ii�	�zj޴�?I�O���f�Y�	�,�,T[&�ڳ���E�ϝkk�� e���d7�T㰨�
L��)"O���۴���'W �����X�<y#�Y�#�����o��w�h��&ԟ&�� �!��(@zd⡭Eա�`�Z��p!r+��,Fh��$Φ9iM?}���e��p���z b$�@�>}�:ғ{¸�["��jrM�i��4��'��6��5`a��;?�R�{d���^lCS#�O�<o)*`4h��4�?�-OF�'�����.���po�Z@�U���0���I8'�
:� *j9�)`���%��i$'5�����SP��s��٦EN6 @m�e��>	�!/=~�!��7���	p�����!V?���'1=�]�Ra��U�}Y4oJ#����'�����P��b�}�O���$_�}xգ wߊp�i�
���'�ў�?�c����iD�LAs��glx��'�7�IZ�6 l��b?�@U�ίJ�dA!��$��y��J��?a(O��i�D��F~"�-i�5KE+[!+|�p��iֽ�M���;U���J�C��tI�Tԟ �	�1:��F]�8�rJ�Y!Ը���J"?@5��ˉ�z�te@�:|lX��`��:������ A3u���;-b����X7� Ō'ik|�2e�<y��ʟ$�����?����Mcq#֢CCxB4cB8����7)�^?�����'C����`ɔ� 8I�@
W�VʨĂ�	��l��4,���'�.7��O���$��usSÝ�X��Y�n&J<����{H<aR��   ��   f  U  �  L   �+  }7  �B  �L  'W  ca  Zk  u  �|  ��  t�  ̚  j�  �  I�  ��  ͺ  �  Q�  ��  ��  �  `�  ��  ��  (�  k�    � T � & /& - �5 �< �C �I TP �S  Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�� |d��"O
`�(�;���8���-0��1%"Oj4��ND^[��"3/9�0|H�"OB���H��*�ʞRy=a"O�味V�!X��!&F�:J�$���"O,��a
���C�Ą�M�"O,$3%o�-���p���+Ն�:1"O��ݢ1����`���y14]2��i�<�6��{_���c�H�`�fX�$Kn�<��A̼VI�xR[�)�Ć�pඤ�ȓA5��('nߡ4�� �)˩%� ���,��r�؊b#`T�eT09���ȓ!�b��g��}�8�F��-? �ȓ
K|m�ș�VṔ���2�%�ȓ"R�X�j�4JN�1�˘X�i����̹	_�jZ��1!g��zܶ��ȓgil,*�J�
j�Ne��i�J%b���f	�(U��:���G��$Y^م�~r�� S�%T"���k\�jx�ȓ|4�1�îJb��@ӵ�ݩn�V��/[`�"�v4�R�!ʎ<��M�ȓ`:��z�ؚh�J�Z��$HY:	��H��p�m�C1��!��B:��0��EnjZA V;9����J[
2���	��4'J�EA�IVW&��~�(aZ��ӹ�>� o�Y�|�ȓ�f�A�
Ο7�H��M�$�����mޠP����/���ANXo*�ȓTv�����{ ��-7�*h��I��sB�8�8���3����ȓNe*M�悡;������X�o��!�ȓ'lj�#F�m�+R&;�|��IV�I�[�2lh�-O�()��
^�|OX��D�Ɋ(B"Hږ?*�K��h@a��O�0X���Qȉ�ׂ+5Ӡ5`�"O�x�&E6��LRGؼM�8=��'��e�\���@�hd�נK8I�|�PA�%D��90Gr�� �M�8C,LI���6��M����T�uw,�1�ɛ&*LtQf�E:!�$X�d
�bj�|��ʉ�C�=E{���'�p���C�x�	���#��j�42Ց�"~nZEiޱz'�A��9�ʆ=B��B�	�}fI)lOO������1B����*�	�<iU+W-@of47ꙛ+�h[�H	Ch<���\7-���Ä$Q:�P���fyB�i`qO��iS�	�̀m�2�<:�*ԡ9^���^l���uqkLp���M��'�|�S��?O��Q1��9�,���0-�@`�w�|ҹi<1OP"|R��	�~]�%��[��t[fKr�?�J��d��uy(�#6�[�
%9��A�I��O��*�D��ab�V ybA�� '갅ȓE��ahW	 Rp$J֨ɍEX�Y�[�\D{��e+`�
}��B�5s�%�ä#��=�{���&E �	
r�'x���cS�ē�p>��mԡ:����c�]�0�F�}yRZ���<�}���@iq6�K�_�d]x*�ԇ�h�Nl���[��Z��L�#�)%��=I��:�"\��wm�y~Z��B�],@�d$�ȓNxz�`+�K[$�3��G2���ER�`�C/ݱi����C�u�⠄ȓDv|�G�GB���a^.p&.�G{��OP���&E3�$|�G�a��t�	��� ��9h%z2�y�� ����"O�\��B�	zyR�L߂r�����"O�UQ�@�+y���G�Է
�j���"O�#����(lI�HC�/+$1I"O�0�ׅ�bBM	s(�`�)P�"O��D�Ђ�~�x%�!;���X�"O�}�Cf�&F���X=���r?Y�O��� ��ױT��$��
���#"O���C�߲DyH����8���I3S���Ä�� &�"}�-�>~>�vf�M�n���&�J�<�ɟ*I� �ۗn�'N�Ƞ�� G�<)�B�)^0z䋑ԝ8~����lϓB�����MՐ~�;��b��<��*I�x��h�%X�n�Y�+��|��G��S*S���A2(I�TE��zF�xazB��*�2� sfE;#_��M�v�c���	�zڞ��vH�|wv0�W��:NxC�����Y�+�?p�19ơ�?~d#20D�0���.vU�\,9zd|p�)�i��}�ŅA�rod!���E�>ͱ&�i�<Q��\2X�*�A��5�a���gy�\�6H�OQ>u��e�	p�`ƇQ��xrS'=D����ӯ\�v��Sk:�Q���9��Nd�����V����0�۲M��bb��)�!��O\�"�cY8Ou����)�>9���{W"O0pES�*ih8���9m��@t�'�����"�(@���k����B"�| R�>y��'�`�����m�R�K��J1\�	�'@��9��C�xŠ)$&��W�غ�'8��&��1�X��k�'(���g�Ork�����F]�Uz�'A&8��`ئd��� �]�C t��N�|��I!uL<
5J�,&C�1�3�Ν̘���\�B�6�,K��$I��̈"NRB"F��M�b)r���P�$$������c��9sr�����6�Ԭx!ax��$g�����Os�R��,P=�x��-
 <��#�Ab�	6�H��B�@��0m.��'�z`�'�)ҧeJ�Q�P�V&v��R\)$N4��'�a~R�K�2}��p�d۶8�b��	��yr)��k���{��!��H�=�yR�(7E��+o��tт���A0�y�d~�v�c�@�y@Q)E�5j�{�i@�-���zd��^�O1�	�4��p	�!�p�p��DoC�(Y4B�ɱL|Z��g�"|�eq�� _0��?9��	�Gڲ�J�i�'��Rv��[�!�dJ�����'�
	�|�3Qe�Nj�O�����^��@K�1�ވ��M�t�!�$��#���6��-}k �cF2~K�Gy��'��h�Q��6����m��h6y���HO�\2A���_��"�U�6��9c"O~�X�#Gۈݺ�i��)��賓�'~�p�c�V1d�ԛ��/�JH�u��O���y'�h?�1I`c�:FT�B ���=��|�k!-/�hq0$_+d͊`���C1�y"��oX��RM=(6Z��`$�yb&�n�|�e���#nf��q*��0<i��d�<C�j�HG�X�bV4;�]/#!���[��T $90���Wjԙ�'�z#=E��b���K���.��B�X$�yb��f)�����&��]�0I#�yr-��a�$���N����1�J��y2�� c$�uEH�$�R!���yr�%RG.Å
؋R�L)&���=	�y2MA�_0�D�b	�� �3��C0���6�O� r��&��>dB�!b`�yG���"O�k�FF# ����a�I*���"O��Ǐ�ta�UZ���0	dı�"O8�����
��Թ$�C>�h%*�"Ov��%��O�L�be�)x�T�y�"O���O	@q1�I��37 �I�(F{����)>l�ڥd�� ~�XA�#P5y!�D����TX��?:J*j����2��O���$Hkj�	)e��sE|��d{}��duӖT�Q�%���R#��d.��*"O<��!��~��@*���}���'�iFy�$@�j��Q9�mS��ɠ� �?����S5|���U���d�b˃o�@�'M�8Gy��DG��98��F'o$��
tJ�8#�!�dE�d3��;7dEXxD@���##�!��5)ðš����zXz��}L!�׸	讬���N�.	�q����sIў��� Y3b������q̙��JU�\m~B�I�B"�A �
C�ZXA�ҫJ�d�m������k%�P��\(�Y8A����2D�X鲣�YAx1X���6l�A�F�=?Y�0@<��ޞT�,�b��N����ȓ{�`�&�? B�Y2��M	9�@���0pC�жn<�	Ұ���82r�ȓ~�b�ĝ�&����5i�%)
�X��n�.42b��B� ��D�Ǟ<p��o����4�[�4d�<A���E�v��ȓ}<�G���<0ѨW�Z:�*,�ȓh��|��N������׭�7tv�ȓ�ȝ��&[�0���B@N׼T�.��ȓ@��A	�a�T�!F$%���
�B� �Cʔ���Ҳ�K���ȓ�a�+V�y���.Z�c36Un�I�����한8�$�V�^�C"f�R�(Ȯ�y���9%16�j݃-8�%Z�䏘�yr��I�6�r@束>�=�bU��y��W@a!��!K3d"��u�� �y�B�(��B�]��9��Մ�yR.J)d�R1�b���W$(���C��y���T�rS� {�D����y2�;T:���P%m��U`R�M��ybm��U�zZ�T;��xV���yR/�i>��r�ڞP��Kg��$�yB��m��=����@Ŷ!�����yRg��9��	�u�	1�R�C��;�ybOD�\H���D�*DN�*�iU�yb��\��lʦ��8/7�̫CB���y�aH9	|�[�d�:o5n�)��B)�yB.� `.�@��a��kVD��H�y�FJ	4���Q�XjRȂU�̷�y���b~��C��S:�hq���>�y#\<H˰Uj�a�G�z���L��y��� �Rx��M��N]S ���y����b�9��iBLBC(���yc_�G愡q�-Ņ b��KA���y"!ׁiɦ�����3-�t�Sp�J
�yR ǋ= Aa'��5S��k��&�y�j�9ja�wn�	 6qS0ML�y5
��XaS&���H<�Ю��y�� �G��ܢ���`� �%-�yeF�Z�|�w�F�Fi��(�y�G�T[*PZ����zd�F��y«��s���ʕ@� H����ƫ�y�R�Z��`����:+������)�y
� ��PS)U5!n8�X�bT��v��"Ox�[�a�='r���Ⓑ�@��&"O�u���K��4��X�i���r�"O��Q�N�u'���$�b0��"O��!����$�+�ˌ1$u��0��'B2�'��'r�'���'���'^����H��z!�L-+|�]j��'&��'�R�'��'���'t��' z���5�yP/�C���r�'{��'�b�'MR�'b�'t��'Ӻ������u�#V��X�MQ�'���'PB�'���'�b�'�b�'��m����v��4��o��l�
���'���'B��'��'[�'�"�'�Vy�h} h�䥓G�X����'���'XR�'���'�'���'_z=9$"Ћ�P���@ @;&�2��'���'��'���'�R�'��'�䉠0g\)����&Wf�+'�'���'���'���'��'�"�'�`9R����4Ė�J�(��'?��'w2�'T��'�R�'b��')��c��V�KYD�Sg'y�� ��'���'V��'���'_�'���'W��h�q�l�#JN�:�|���'��'�B�'���'�R�'UR�'ƘD�D.�9������˽g�����'��'�B�'2��'"��'W��'R�i�iYPL����,GlD��'�"�'"�'Xb�'��i����OB8�,_H(IS���2ě���@y��'�)�3?�ѿi` H��dߛn5��k�����1� �����EĦq�?��<��i۠����'�XE��ٷv��8�!j�
���.�24�v���x�H7R[��Q�~�@��@A<J!�"*�l���o[s̓�?�-O�}��R�f
�Ǌ���#&-��֯��'"񟢰lz�E�႟)D�����W�>h�X�M�i��>�|*�%ڋ��D}�\��%Ϯf�C�G�	Vh�Y��u�Dj�d.1w�x�p��X���d�'�&y"W�Y�~�8��F́�<�T�X�'��Iq�ɥ�M{�av̓ ��hfE�X�lC�aJjl���>ip�ip7�o���'c�@�g���\0F�����	�O�5���7C*�UQ���5FR�MٳJ�O:���BQ9<�t!0�E;a��[���<�-O���s�l�b$Ւsn�xנ�� !�T���p����4��<�'86/�i>Ub`�ѽC�պ4M��a<�P�Ua��0ܴ:��6�'�tx*¯����$�0NDX��g��#��5`�
�"�p�S䈖�48�k�9��|�*Oj��Z�u�ѵ	��.L���ī����ݴ(�D�<A��$��
̒�k�i q�D�_���<�*p�B�w���?��	�>>���}���Wߙl`6퀗��S@��g��dCVi��9����`M+}�2?�D�oךu��.�8A?�������?)-O���X�VN,�y���,�Ҧ�� u�U�w���ybHk���7�4��O���ݴ�?iĭ�Q���PQj��)����Gߒy�@�@V��<�)��{��G��R��S�?���$����J�l��	��|!����柄�'M�)�':\�ҢԦ>v�1A5�źT��(�<є�i�^�@�O��l��d�'��9�Q�B�r�͉2y����s9OH�O���h�8�D�i�>!;E0O�a�U1w?@h�j�<rqi'"ݑS�Z�1��C�z	�7�$-?�'��$�Oxp�JW/�T���AŒ���U4Ov�O�mn�^c���S�?�i����	AnLs�Cީb�(?1"X��iܴZ̛67O ���	�!EO��.�b�m���H7-%�Rd�L�d����O�Y)a吠%o�L�D+L1����7h��<��� F��	z��uS��H<��i2��z�H(�H+�C�'9�l��%�̲]�I)�MK�C�>��i
�<*�퐍8��5GX���r�dhӶnZ�+	����#?�G�[� �h�C�Ѝ���p�x�2#�*7�j1�"�	|���<��U��\
d�|�$l#v�
J�RU�d�iQ�@B�_�`��h�� ћ�w����S@��_�x,��G�����M|ӊ�l���Şe�^�����<�2�e���T�J�VA�����<QP&
S���䓂�$�<���Q�'J���%���B�A@���۴yQ
�B*O0�dM)R.J��I�f�����4����b�O�$n�2�M�'�xBK�j�T�Ul�Ɛ�P-�y��'�F�.F"Q���_�p�Ӟ,�L���L�0b)BYH�N�%!��,�R�?h�iHਗ਼�rǌ�����=3��QP�垍��7M�/5����ӌ06	�b���F�\E���R�F��z�u��$ɖ3�NI��]7��S%_+�LZ5��=
t -��C�w`V�C&"]?�h�ԏA���F��)Hڑr�3\�K��c�<2A�vE�,$=�eb$)R�$Р)��\2zAZ-\�J��3�
�(�-��!
��"�+W�0W����Proƹ G�5n���� k�S�@�	!��j�p�4�?�Q(�J"�')R�'�ɧ5�C�HD���J�� �x:1/֭�M��x(����$�OF��O����O�Э-��t���
,�Hc �.�
ҟ�Iğ$��ߟ`%� ��ߟhh�îF���������h`�.>�<���4?���?)���?�������O�|:��0T�yK���Q=����4�?9���?aO>1��?�RB �g�fo� x�Ԑ��� ,a�KҌZc���?����?��?���?����~
� *�چJ.\�(�ɑ�f�t���i�B�|"�'��j�0P.���J<��kA�o`���%z<�C���ۦu���T��ǟ4XdcUB�]���ӆT�D@B!��+'lȹ��i�i�J<����?!EC��7�Z��<�OB^����]�_�D� $G@�c�`�ڴ�?!��=`�H ���?����?y�'��Ƃ9���R�Y�B)g�-�B���i="�'d\C6�������O�4�:��$D��H�A�VK3~D��4|��0���?A��?a�'�?����݁����5@}���0�	sPql�-�0hY�G0�)§�?�K�< �>����� k����a�ĥ$�6�'5R�'UT8�!���Oh�$���T�$9�z):E�R|Є���;�	�d'�b���	ȟX�	�J�� ]2-�.<�G�(a����޴�?)����d�O����O�Ok�z��hQ� 0L�z|$�	�_]�I}�(q&��矐�I`y��rN��8�/��'=,8��b�y6�ȡ�V����ʟ��IS�ʟ���2x�aLڋ:�@���B�ӂlCb`ɟ|�'A2�'�Y��R�,
v�#@��=��bP�<N��ir�ͦ}�����R����	U����hb͙P�V�HW�m�qc6i����'�2�'5�V��!��{���'��J0ݬ>�4(�1���!OB��1�l����>�D�O���J_(��dB���"H,B��Kh
���%n�@�D�O�˓P���,�����O��闓o�tc��U�\Q,ᒦ�l�$�\�	ӟ����\�S�t�; �xuh��И_������Ms/O>����O��D�O0�d�����1��67�du�b�pu� ����u��쟼��/@V�S�?R�tcQ�M/FM�0��"p4hnZ%61
e��П0��ǟd��^y��'��[�+UԨ")�'n����Rx�@7�F�$4��+��S�lPC��: v� �囡m�P]a����M���?9��}b8��X�Ԕ'���O�3�H]�!t�u	��G"N�45�����h�Ob���O����"rb�Sw��3O6&dŉ��6�nߟ �3�Ly��'x�'ɧ5Ƌ����0�6¬�!�V��D�&T!ʒO��$�O��D�<q���e�\LF�҉'gΩ3'A͆K|�I/O��D�O,�$9�d�O.����XVhE�� ���Q��ؕ2�h�'c6���O*���O�ʓ��$�O��,���
oWPD����N��h	�4�?a��?�I>i���?y� �~RDmY<� ��<s�
=��D�O���O��;����+������[a�u�Kѱ��y"R��v�]lZП�&���	П`�4�|�~C��	! 3�E��N�UQ�lZΟH�Ixy�IV�)����?���"nR�n���QN�=S�6�:�e�$G��'�b�'�B�`����?	
 $P�S�F�)W��䴘E�oӆʓW(8���?9��?��'���2�s���%ڸ���O�Fd�$���i���'J4I1���i�?1�	KO����ˠ��	f����6i�7m�O0���OF��]|�i>�X@d5B�!?��;�(�#D��7��J+r��O�D�O����|�'ld���n�8g�* 7����Gw�����O���g*�&��S��\���I�,X��oW�$��9�%͎�	�ԩ�ܴ�?A����Ĉf��'L��'Xr�6	� �P�L�A萭 rG^(�7�O2��3	�r�i>a����ؕ'� L����,�b��	�5��)�
wӖ˓�?�I>Q��?�)O�[ыD X�l���M]0�r� �����	$���	˟8��my��'-�IѦT�����"IKB(r�b�I���'Z�'�ꧭ��X(�)ͧo*dɲ�� ��Ѐv�;b��'*b�'m[����ɟ�`pL��|�]�~1�a.\�SS��1�S��<\�'���'���<s�k�c�D�'��%���$�U �>m��|�`��I̟Rj���OB�/��R�T�?�8�����ޛ��'��I՟(��c�d�T�'Zb��5V+]&g?N)�A
�|�&<��m�(�ē�?q�w�x52V�S�dDѮ	O^XxV�կe>:U0�(K�M�-O$)*�h\����*�����'�����v�D���䋸RpU��4�?����y�?|�SΟ���x�ܴnv|`���҅=߮�%h�&v�@Dm��k	�	�I؟���˟���pyʟ~`hB̛{�J��K�1�$��̦ё����l~�b�"~���Ȓ(�%ȴ�����uo��v�io2�'|b5y��):N��1�i�M��\h�V�=��-�%����'h����*��ן��g��!y�)�6!�ܡR�H��иn�������{y"ǵ~"�I�2���1q��k�xY�iX>@6�([֑�r/m~�'B�'��I;��4;!"˨(�Du�'��3'.�5��O	���?a���?-O����O����C�	"8zg�ڠ+�24A4!�3�h�D�<���?������I"5�'i����@�,X����m�:�'r�'��Y���՟��T��쟤I��riZ���/Y��ؠK�f�Hq�'42�'���`xf$	q���'�����V���E(1�G6}kl�$jpӶ㟌����JAo �`&
O�R���..l�ȅ�Ki��Q��iMR�'�2�'��	�$nmӺ��O����4��'��!y��SQ��J��43�����I_y��'�&�i�Oxɧ��4h�<��Мxtb����/e�n�ٟ�	��@��4�?q��?A�'�*�LO� LeG`�L�S�T�UԼP[�d��+"0��������Đ~b��I�N\�����	R:���
Ц�AP(�(�M���?��������?���?�ӂ�	
d�H@
_�<IR��0	N�n���N���'�i>%&?��	2�z(��K��'�Q���%G@`��4�?���?��0��'�R�'Z��u��X�v��`���
*PY3�N���M#�����E��?��	��,��^5R�8P�QYw���v�B�zL�oꟄh��̪����<����Ok��H�I�����ˀ
?��i%V�<���a�\�'�"�'AbQ�p�1c�"j:rK�	�\�*�{A�V*)�͹�O���?+OKg�����O><r�U�B2�8
�P2.�6A�t��o���<���?�����FZ��'+׌a��$t%v�2ӨܦM��m�sy��'������֟k|���8nV~� q鈇V�x�@��Dbz듎?����?+O�-#�×_���'W~���G�:�)R�
��<"e�ft�:���<���?����0����� n"m +Q#�T(��_�ʴm�Ɵ���Ay)�맇?A��:H�88��31b}~���cS�
N��ɟ�������`x����ybџ�:�^'IF9;�M� �!��i��I*t:��ݴ�?i���?�����i�}0�D�op
 ����^iB@GgӖ���O`�7O����y2�I�GHṣ�R�PI�!�*"5����%4�6M�O����O���B}bU��B�.�4�, r��R -۸��gB��Mc�]�<)����,�S֟dA�ʑ ZZ%3�&�{.tĻ'J��MC��?���J�t�"�P�$�'�r�OhdQ@L��oE�8�	�fF$j��i�]��9Q	{���?I���?Y@�H�W�>@�!�6��s�^*\����'Yn�"B	�>�-Op��<���;CnJ/1��p�tR�tF�x�7�_}¬��y��'_��'�2�']�ӧ�F��g���.�2�0�ԁAX��@�j�5�M���?q���?9�_?-�'L"`���5��#�fhuA3��?M�@�'="�'���'��S�|�&�M)���"�
M��Փ�␹)���1���M)O���<��?1�	 ��������L�_#�A�c>�r]��_���ʟx�	ݟ@�ɜWڀ�ٴ�?��\� Q�ɋ�]̶$ʂ㌗sHDyp�i��'X_�(��F���8�k�Ȍ2we�s4����Ӗ;���l�џ��	��|�	�L1�4�?���?��':��	�­6=da���x*�#��i>"Y����b���e�i>7�Wo��!��	t�����+]	����'���8r7�O����Ob�)���$ľf茛S�H�x�P���B("���'DB�ݻ�|�O�|P��0 �w��,Ci"z߼�mZ�V &��޴�?Y��?��'�"���?��H!\��$��8��(��
	7xw4L��iMn���'�'g��'���?����&r��[�cJ�>���A ��]n�&�'�R�'�I�7�m�����O����O����b�d�I,6>f5Jd�kc褊�oo����<��U�<�O��'���&sM|�GȒ2�>�"h@H��6��OPh @������0�Iҟ�ᬟ��I9c�詃��&r8u�d�˫?z�6��OH\��=O<��O���O>���O���։��l�Q�_i�<�Y�56�ai����������ޟ�®�(ʓ�?Ae�&s�����5+w
���">+g�-��?���?���?�-��%��٦�k�҅1�Ң���	N�y�@)͆�M���?9��?�������OHT�c1��O�wA�Xs� ъ �j�K������O���Ot���O4���i������̟�zW��(G�|s�HyJ}��	�M����?���d�O�e��1�J�Ĥ���)D�)" �c��,L� j��e�`���O��D�O�RM�Ȧ�����H���?)
��^��3d㑏GM�0�2�ځ�M������OhL��&�i>7-Y�q�m��k,m���d�J��&^�$�M��M�U_?��I�?qC�O@�!��U4��
�匑VA("��i���'J��ˋ���ю � �2�E�/>���aVL՛��!_t�6��O��d�OH��QW�I��(ܩ�DU�� 0��$��N��MC�� �<1N>E���'�LI�IE�u1 �%G�˪�H�@u�p��O��䗒��&�d�������Hm� �(��4"vD�0ƚ�Fp|hn�\�ɚo��)����?�O�� @�.������ne�Lٴ�?q�k&Cw�'���'�ɧ5&A	�W(��i���5����C�����������<���?YK~#�H3Zl�� ���(�� Ԁ ��@�x��'`��|��'a����Dl�\Q�+�'�`���� �����'��Iҟ4��ӟ��'� 䋢eh>遷�Tc�Հ3MR�x����"��>!��?�L>)���?aQ���<�d��T´p��(`�kV�(!�	ڟ|�I��'��$�4o%�I��N8�w@-��i`p��S�mmZߟ�$���	ߟ`���9�	9����Ÿ?�*�P��\&�87-�O>�Ļ<I�&u��Ok��O�m�dT�4r����1��M� �+���O�D�W�H�d.�T?=��+�6�Tt�DT�t݁Gch�p�kP(MP��i#��'�?��'��I' �DPzPE@��:���d�X86-�O���Ϸe9��b?Y�jF�r~����丫��c�D���ϦI�I�����?��I<���S3
1r�����*��	�?~	!E�i�2 �`�'�ɧ�F��֋BNF�@u���G'�)�t./w�l���	��ԁь �ē�?���~
� ^ԓ����A�G(Q�kȩ��i��'�x���/2�)�O����O&�H�B/b�D���\�<������M�I��T��K<���?qK>�1@���Z�X�H?���RIg�
��'ʴ���'����������'�bbs�O�E|���r�H�V`N��p�)>��O����O��O����O�5���ϥR7�aQCm�"R�-�a�W� �����<y��?Q���v�8Χ-^��0n��p�H@�p�� cIp(�'yR�	ٟb_C!��S	�(����*"�h�c��tP�6�O��d�O��$�<��
�w̉�5f!K�����"�P�D�P�r����	e�'���
�	kB�'��	�?�r�X'�C�q����5m	>1����'�"^�@�$ǝ��ħ�?���;@�'r��rPQcښp�JE��?!"	��?1��i�("Ѭ|��D[�d_�h���M_�V�'��i�%��'@�'����'Zc?�,I6�����R^ 0���4�?	��Yc���i_�S�'`*(Q�
�.C>�2�G�/31�Ym��9t��ݴ�?Y��?Q��a�����B	�!�{ʷ~�-p2A�fL7�ӺAC ��3��ɟ�RH�o)�12u�P�?�\���^��M����?���a].�;-O�'�?��'�(`���4K>�8�C�lB`�k�e=�	M8D�N|r��?���lx�\9��Y�u���ᬙ�L�����i��݄;˚O���O��OkL3)#�����xɌɻ��2����L�2b�H�	؟D��Uyb�ʭxfJ�@�(�0�xE@�횉t���
��$�D�O*��1�d�O(�DA�U�V�I��ͱU��R�D�1"��!s����.�ɺg���^#8��6W�'԰jA(��u���E���^�8g�˺!v�Ӡ�-L���*�|
~��Q�!;Y�y���n�x��@/=u��ZR&�<�Ǧ�� ���{��o�	�Vb�xܓ� ]�>2|X)�505ɼ�؃�Ұ�𑃃�D�fsk �X��A�#��q�$��>�1�A��S�Ĵ�Q��p޶�J�.X�`�UȎ��0ͩw�YG�jᙐ^R�V)��m9#�Ł�-�e�e��ף) �4�#%Tw������f��ם��j9`��'٦<B҅	������#Q��1�'=".�i]�9BIL��n�k�#E�;� �'���#_.�	 �T�E�N@i�o�wD�?����$J�ZЗ�έdM㒿�H�4�Ѧ�ם}� s��J�zqRq�6% �7n.�'����nɧ�O���a� ��uD��z��I�'���b��KϘ �%�֟or$A$�i>�J����*.3�=�5m 4�daH'�����'[��'��Z����'����y�B�H�z=��V�Y��0p�G�[E���&k�;~Ϧ��Ȑ0 �����|�
#r�)[�m��<C6��b��Bf��3�Ҫu�h��!���+��L>��bO�(�}y��vX��1�3�?i��?A����?�}�'X`2��9IJφ(>�Ctɚ9\���P�zńb�e��y�x9�̇2��	��HO��O"�8ܐ}1-� :��I�V� Hc0�\Y
<����?���?q����$�O6�=D-��d��6$��  㖾:E�-��+�y�P��!H�QTn}��"V���O���y5yKP
�9v��4��k��L19$��.��D�g�F�{�@��7��yZ��ra�(��z^ʁZ��38�`����y��0������}�ёf�!�I��i�?:!ֵ��	T�I'����$��g� �z��_"Q��c� ��4��>Y^�`_?Q�ɺ:	H,Zc��3�CV��u®A���`p������	�|ڑ`J�P0X4rUJ[�B��y��4e�D4tg7MB��3C�� 8�l��iyA5�Ūg	D�qaY�-�v7��n=f:!MB1*�t)�)��9s�x����?A����dȋdYZ�B�!�W��sh�1O�����&���\��\�¨�!�!��P��Ezʜ) %��I�٦7�ҥ�aM
���'�d��Jf�4�d�O�ʧJ�}��;8���.םY�|YwG�1o�4�����?��̌Gw����HG	^�x�$(� a��������K���"&�VN�E�TaD,E��]�D0�&��k�6��%��hCx��	'\���v��x'A@�A����&�Q�*>J��O�A�'�1O�P=SG�!єxq ߰u@�"OP��Z�
	d��.D"L�"#�'p�#=y��N9V�h��c��zm���R��C9���'C��'�|��2�t���'���y7
���a8���4GQ�3��+İ9x�I�26��r�I�C4��-b�1S �']�\�km��Z�`Kec�*s��V�1m���) ���o��ҥ"E�	Ƀ�N��rD��A�~�ĜRy��%�?�}�I�l���Ǧ��(I6Uc������
Ǹ�&�`��	��ۃ��r��e
A ��W�>?��i���'$�6��ON���Oʧo���b-�<I �c7oX���cɛkt������?����?Yr������MӚOmH4�������C�K�` ���3�x"AW>����"I֘�J��B�J,L���'��)!�#ue,��W&�!J�0Q�4���?	�����?i����'�L����/V�D�p�J�_�	��'��ikA�@8a�H ���d��%�y2$Ӱ�d�<� ��%��&�'�
� H���.?j_�`�ۤ��%��O"�D�1x���D�O,�Ӯ]3L��JW�W6�&���>��e/D�^��#Ye昨"ja�'���YjB�k�$�����(�+��>�nu��� ,$���Yir�ɠ��I�� �%,�I%u�|�$H]�ɨT�J1�7�Y�;1���`��svfB��&^����C�7"J��`BE��&!�d٦��q�/B�`TjH�eH	��#�H�I<MF -�ܴ�?����ɜ2,^��A�59n96j�P$d��U�Ҥ< ���O�qy�D#b������ny*�.˧��h��۹���b�0Bz@��Ov���֞T�> 
��m�Rha	����O���bX9!���4�G�[���I��1��O�o�Mc����O���u���Ew�5	7��Y��шyR�'��y�GB�g�����̘X%n߲�0<�7�I[��$y�B&u3jȔ
��>�ȸ�M�П�IΟ �v� �9����ǟ��	��а]wm��Dl�iT���I��U����B��y�v�x≷.��H8��i�b>5�K�����ŏO_\᪠eހ:�c�dH��L��'��;"��v[�R$j�@�����	WT��nkޡ
R��'#��\Z J�Gg�] a�,��Dc�M�)�3扄��\Z���8�tʃ��8X!��Wv�J4�N��b�M6(�I��HO��4�D��^��	���Zr��婣뀚Z�1V�Z�d�����OL��O��;�?	��?��"2]��@��U!E,�`��Y2Y���P�H.y+W�'�.����ߊ=� a�2@��3ޠtC��,(&q�3l\fD�@�
J,�0<Q!�ˬ�`ܨ₆	CP��n�+1V���ɛ�M��i��Z����O�K�T)��
�^( `�X�`-��Ex��'��$��@�~Ա@�D���|�@~B7-�<�G-�Ѻ����?���V#e6,�@�m
$�A�9�?���Ѹ����?�Oq֜(MV(_dJ���9X雖���*�^Y�WB*@�^ġ�D�9�p<A��Ru�@qJ%��h]ݴ|�hз܍V��F)[�.�J ��	#r7R��#��	B�J:�g�?xz�
"$��A�!��I!64ر�T��|`Uꃣ�3+J!�$�ަ�$Ԕa���F�$��9�F\�I
���޴�?�����I�"U��$B3HD�|i�G\+���S�͆H�<��O����IԴ� ܉�lOhy*��ʧ*�ޕ����ik��C���*u?�ؤOr�(�L�e��Йc5�]�< ��J���!C`��Su<��OҽC&�'#�6�{�F�T�����ˇQ�hBF�`b�T�	\x�@q1�R�bp���TbB)HҞ�Z���U����H'�	�����e[��Lᤄ�O����i�B�'���ˮ7�xbS�'���'��w!,�t,�8r���@��[N�� �D8?�yr(��Ft�Lq����r+ʴ׸'+6՘ϓL���$e�/&��*5�	'Lf�:ő|Bg	�?�}&���Ԯ�,)��`w� Cz Ey��'D�p��ĵڦ�#���C��3�k*?I��)�'l�t�r���CB�q�d�@�Q`~��qJ �4��(2���?���?�b���$�O<��6�6iyQ��T0��f��a�h�y�矖!�%!��O�Zt-��˃��O:�Htl<dƎ�c�H�00-�V�=��q
�-�4b�N4A��2T���3j't����R$E@�k�i�&��(ڡ7�"�$�}؟l`a"	�Z����J4|�&�ۗ@0D����GѪ0�|-�t'�)B
Q	.�	��ML>ɗ��P����'L��Տ(X�3s'.�RU��/ݲYb��'KȐ��'�"0��tR��+/��O�!:F��v|�٢��U��1��'���f�/D>T5[�JƟR�hj�G.%��x�T�1|���b�2q�(ˉ�$�o��� ���0k�@�p�ۇjζA!�h�!2�!�D��Q%X��f���YK ���!�G̦�N��?N
�"EU�Ci�]y��q�1nuq�4�?����i@ "����O� ��%�\rarC�5`��O����]?'��􊢇:?�O6�;^P�c�l�(Mz�81e��Q�h�'�6�H1"m�>a��)��<�4P0��G;��`3>��v`���D$?	&?-I` X���($��b� �ag$�蟌��	�?�XL�-�9V�I	�杯�8����z�'��X 5-��j_�$Bt�j���lӲ���O��DP*b'f�R�
�O8���O$�������2�I�,������KZG>����=;Pp�q�D�hٶb�*o�b>�Oਫ�iK���S�ÚUyv��E��
��їo�=9� V�[�o�q��'����茖U�N�qCG�N@�Cv+��G�J��L>�tnZ"y���
E�9�@��%Wm�<��A)C3�EQ�T�B0Xt�j~R�-��|"L>ѐǜ;`ڔ�ǡ�KB-v<yr��w����͟���ן {Xw���'�)Ҁ ��*�ɾ�)d'��HbD���D�tF����F{$��`�7��O$)���>�hi
�L��oD�1�"��yKR��I��x����e�@~��#8�c9����{z��Ku'��A�qS��@��͟��?����<��b�<��-�GH	!�yO+U��yФ`��J<q�I����'9�7�O�ʓ:S�����i���'J�Y�j	e�$�Y���K�8I2�'���J
���'`��S��1�i�a���3cF��`�[�m��w[��YH��4��j���S�JR��(O�yj�C���-��z�f0�����}�e�RGz�8�F��4��"ê<�(O$ѓ&�'�xO�T�q���D�!��||p�B"O��f���E@�5��D��cu���rO�lZ�/
��ǌ� ��$z �A>M�%���ſ�Ms���?�+��}���OF��'�ʮ]D�T�P�Rm��"�/�On�d�9��e�F�;u��i���O�V���ވ"����qe� {�<*1���	�6��= 7d�"Tj�SNh�b󉋸PӀU�V����P
gϥna�D�I����S���r�CvhY�.P(�g��3%8�E�ȓ�����@��xI�����2a��q����HOda���dRr��MX�ZZ�Y�DW֦��I����I?I��8������蟴�i�ѡ.�r�x�˴�[@}�|A�ES�Ę,O�I��u1��':��F�2|.���$7�|���D�3Y���d��qZ�(��O��	�[����N�6�l^#��+�o��f<�'���S�g�I�=�FL�&�߳�]�bΜBB�B�� )�|˱�]��T�0�	�j4�oD��"|� �Wl�0y�c���P�jΖV�hDP��@�?Q��?��{m��O@��i>�҇�=Ry� ���Û`� �������[�`"s:8@�B`x��"u��x�P25#�������4��̀���eZl��2K��~jMI�o�V�'\����S3}k4�Ƞ���f�ީ �O��?���'���'[ kyʝ�d+�0�E��'Xd1Gc�P�z�DAÂ;�呎y��<��!jd��#�O0����#=�a���D/p����Z�k��d�ODta��O���a>-���Ip�r��`� <�[愌:��*�lL!������x��Aǘ��R��'1FШ�&��9xF$MY�D�0VU�A3��%Ʉ�܈O���'ʊ6M�{}R'Y8`g�a�T<6��� �6�'b�'מ$�b��i40h2��*[��*�'(`7M����+�O�=T�8�g��t��d�<ѷ杫 Л�'S�X>�PKԟ�p�S(�0�d��0DBa1g�ʟD�I�p'���"�@V�-�i[*��ʧ#nY�'��<���R�ѿg���O���ԣR�ol�Sa"���iD�T(NO>Z|Ã�yV~}HgB�2��ɐ?���D�)���!ڀ�:bjP�|W��k�a܁v��B�-B����m��E@� A%�,d���D h�'(��$�щ?cH( ��>T�z���o�����O:�Dɠ7�(��@)�O���O��4�,ۀ�Ė�xb�A� �V�B,ź,��l)"B�?Az��y���-�b>�O��e��g��-��hy<�*B���M����i�:ep�Q	ӊl3�;�iɯ
zl���w/L�p��`0�1p��8��\kT�4�$�8���L>�5&ƴK�X!���� FV�4�Mu�<���^-f��<( )�9z��phV�g~��-�S�O����҃L)Rᘦ�5�Ɓ�ס�@�{`�'kR�'��l�5�I؟��']P�L���v�*�id�E+��ԙ��*�dQD	�q�\(��"O&�A�l� �w�
�>��5�sFt����7��8_�v��OV��p<	��Dw�Ш���
��D#w�9'����+��?q�@�(�~�A��L�B��$�r�<�&$F�WyH!(`�S�b�-��Gp�|��O$51U�禭�I����Ɖ�(q�Z�9աG�aE�x�2�T����1A`(�	埤ϧR�����Re~ģa�!U��P�7��E��+hl�l��1O��U��Ol1I��A�~j�B�D-"�Ƙ�ccFYb����^��p<!#n�̟*L<�v�ۤ$F�!�Kڪ����`��f�<q���~��YЧ [�m�țAf<�b�i�\m�C�(�8Eآi$o���ۋy��?A��6-�O �ĸ|2�h��?�QJ�'� ��C�͚O���"C��?!��1��G�!혧򙟴Z��H��)r��'*��iѧ,}" ��}T���=�փW*J,8�@)*X�ٓ��T�Ā;RPri3��	O�(:e"�M���(���_�rD!�ē�/�ҡI�X�Xh��8axR/ғ"����&_3f�<\diO�$�i��i��'��yؤ�q�'�"�'��w,Z���G�nTf4�ċd1f �Ť;�d�RUf����|
� J{g�:h` o��3����$�m�I4�����|�A��u�V�r#�I狚�f��O�I������l���8�m�i� ��� 3�z���7� *AA�7Dn�����Rle�'�v#=E��%�eI3N��DCT�����paB�i!A2���'��'-��]���I�|2 �;@��j0�X	� 0!郩P�"�;�f^�5�jp�F5��8��"�hO����V�4�0�a�D��`;EL8�Q6��!9�����B,@8,<zB�3ړLe��x��A.$"Dq��oVkc>L
��ʟlJ
��h���C�ʜ^ϰ	��ʟ*�Nɇȓ&4Aqd ߀7��-��U/�0�<i�ԱK�րlZΟ��I  ��m�g��,A`*� �k�(&Wp����<:�SΟ����|��LѺ#Pp]��32���c�\Sjh�#1l���D��&ؚ��d�h��9@��%��Z�4D@$��U�jഀ�,Q����9VT��ɳ��}Y�LI`��a�&!��Z�t����ȓk���؅�:}�A(�iW�3*�4��;��d�'%�dUc�6�D�5���'߮��v�|ӎ���O�ʧ;�p� �*�487��#c8T�Q��+,J&Hh���?��*�X���ʞ/O�h1�i��SV�$牲P9&���U��j�"�Ӝ��ɿ8H�MS�B�l �Pg˟�(���1�]� L97�Į+�jt�>	bnן�"ܴ�?A��䧳?��/E7P�4`vo-���2�̌5�?��?�����<�Q�E(u��aA`D��B��E��R��D�P��	"a�O�V�u�d�O"i�m�����������)�@�>�����������)Zw���rBϷK�x9s�](6+����הF(��'��x��C?�����0Q�E���=h<$AO�/I�\��Wj���[��s$<�3�$�5v �+2��35���gLJ)��]'��g��Oq��'�ĵ;��ؖ)	�ӣT�| B�'�2���R��P�!��Q�
���O�Fz��I���x����D�x :�o�/M���.�5'����OF�d�O�|���?��������!?L\{g�1*���f��e�����C�=@�N	�ъ�xA
9p�<%6�� �3_���h�<��X�W!�g��K��Ay�l�dĔ�Ur��p���>�=#@��,D�^J؟��$d3�28��G�p��U���%D�!b@ŴYf =aR�ݜ.5�9C'L#�	#��'�H%�Ehtӊ��O��j�9+�I(��8������O8��ߵ\�l���O��Ө G4]�DiX L��Ikv$1
@J�(o�N�@��r�����2/ǼYB&�/}4@`���Y�P��H��:�Y$���KE$�걮Y���O�y��'��O@̚�d�rh�E1#J�'Nx��"O�q
P��)]�ꀙb�O-2~�lP!Od�mZ�YV��"b %˂�0B-Y�b��"5�M3��?!-�����O��s�B�c��R��1[S��P��O���]�<��Fㄮ2��S�tP>�:�$U\�B)�Ai��7VX�S0}rg�Co�4���Q�T�B<��s�O����-�q���@&�;U���J�8�c�OX%'��?]
��sb���Ee��8��b`�$D�l�@ `RJe�g���ࢥ�$O��Dz"H�; ����ńhgp�j��G4DB�'A��'LF� �=2�'���y�'�9s�n�fե/�|z�
�<>jL"$K�b��=#!j �җ��yR��Z�Դ��+�yD�0���-f�&�C�>Ҡ��#*N �R�W-j��s�f���g�y�'�C%hVX-��� jӒ�t�����4�?1PMZ��?�}�'VriF��8��-6:��%��F��O���$K�]���-i�ܔ���3����M3#�i��'��S@y�k׳[t%{W�	�l�`�g�X�bPb��Q)q�b�'-2�']v��?i�Ob����.F���᧘�3��i�ʂ��h�b�ų$@;�/�9�џ�0�#�AഁR?��� �G�y��U��i�蘫���+AH�蒮sv �Fxb��Y�䜸�l�r��KA�һ�������?a��?A)Oh�&�	�+Z��-�47�n�ђG\?~X�C�	�4#�I;��T�14t�DmA5�c�p�3�O8�:�0h���6���OV@2�хr�TZ3/� �%eH�O0����4���O4�E��d#�$ՑclcB��~�,���OV(h�x�i"��'Ბ��9b_8��3e�k��*ǓY��m��#��q
��+w��<�@i#u�ߜ3U
���N�4�8�lE/�:L{2!��ZԤ���1��o�`�Zܱa�ЗX!�\`��J.ޘ'��Y��j�����6�|�0�\��?I���$'T��7�T<@~�X*�r��'(r��N��D�G�M�z��AЂ�Li��Y��j�[Z�Q�X>t��7��g�>t�OnU#�i�*�(�ᱍD�izh��� �#��9.º9%��$?ZDSD�>2J�ʟăN>���W�����<l��ExT͂Q�<��IW%Z�t�zw��1E���BTO�,�����*$}n���A�+�H��%cV�p�@�nϟ���0*��7���	��	�杵W���!\�ؘ�̀NR�Ȱ*�=w�zP�/O��0a��&�1��'���%�T%(���H�#��Y5ؖmM�˓QT�C�9�3����6G� ���3�T(BҢ5h��M$�4b�"�Oq��'��C`̷B��|�K�*��M��'�j�A����\��p�תzʜE��O��Ez��	N�k�f���e��b��",B��d�0f+�(R<�D�O��D�Ojͯ;�?9���T&U6_�L�R�M-9Р� �(Mf$��,I0��Tp�F9�� 	ÓF&\�S��OwF��$ז?= %�a%�&%D���A�~׸��!�_O�49����,�5�2�\�zƌ��^(5�&��O�8oZ�MÎ��&�ӕ	"�u3�*�1EBPE�����3<�C�)ir��kC�%H���t��3޸c�,��O��h2 �zF�i�2�'�HDsc-�,D��U���U rn�0&�'�"mG"y�B�'���7r�v�
+�����@��L Wm��.ٙ�<W��xB�Q�<2��!Pu~��QӺjfχ3`�9Q�2`P��D�<��$�D�>0v,̒TI�"�؝1�
Ǔ�!��6h�J����A�|���D�H�!�dɦMत�[	��j�@��d@x{��;��r>Xs�4�?����I��2�2��R�b�BQS#L�ɸ��?->�$�O�h#g�O�c��g~�TfZm1�ʀH^�S�� ���6wX"<���a���b�)�B�;X�<Y��aK����w����I�F�2}�""־Q�`��`Ɂ�$!�$Ƈ-P(�shW%l�l���8Iaxr�6�L>e��FB*d�UCvańC��Ѵi82�'��O����'���'��w�L���r
X%��b�;K�Cg� }}�y��8,$�����m������qO^�+G�'R���ĕ3��L{���+f�z�q$+�D�*f���L>فm��>#V�"gÇm6��2��}�<��C�&����[�mzJ�G�|~��,�S�OQz���A%qThJ��@���� �:)�0�ˡ�'.��'�aw����ȟtͧh�vԳ��ļ��իA-:_`@��r&O&_�Lcbʐ���=���:�
xA�*ڴx�0c� I!�(  +���x��
ߓ��`;6�4+�b�Eؠ�8=v��ԟ`��Z�I֟T�I]�w��� �xbɱN��Z��i�ȓHjDCP��)|�d���L$Ra�<3Z���'�:d�CFt�>���Ob(��K��i¸\����(ypQ����O���/����O��Y�fыa&�Q�B˦m��	ߊL���:�%,ґcd�x��O�
�B�	��qGV5���Ӥg�x��.ٴH��9S�k�>���3�-�u˦E�����'ɠʅ�J� ��&�՞A�ڵ��'��'��O>�c F�� *$�5��H���*�(��4!.�1���[�z�I��;�|�̓��d�$ff���O��|Z�L��?���+N&���W
��X���p���?���p�PL�J�.;���'ME�</�<ʧI)�p�!��qt`�A��ƚ@���O`T[��P�%�Q2�	~5�p��(B���Q8@����lPE��
r��''�TI*�逫��I�ON���Oʕn���D�O���+W��	g�Q.�S!D�.f~q&����b>c�0��̦q���Dj�7J`�M{��/O2mo���M���O��F�'��$H�����Xg�?���A"�i�2�D�O��dސZ4x)C�O����O������U����'1�D�DI�-*A"V�@8�uk��O�����]�1��'z8d���ے]R4`�4�F��Ҩ��^]`��dBNZ P����M?�i_x0p 6ﰡ)��q �:OY&.L>@{&�Oj�d�O�a��$�Oq��I����`m���`�:��H
0����ńN^h<іA�I��zt�h!#�L�Y��'p�"=�,�.�u� �fS����І��3Pp!7�� ������?���?���*�D�O���_�"��*jur$�����S�0Qԭ�y� ���9N�U��B���� ��Տ<��Has�]O�줇��M�2<AWg�I��[��J!�r��OVA��I4RZ�[�\ y�i��(�)hRxB�IrQ�H{�K"et�u��%�$ifBb��h�}���\$�7-�O�Dɯ]�����,l�I1oW����O��)���O�d`>�ЎD5~8�`"�M`~@K��ʎQ�D�U�	_4�aT%ml\E" Z�X$������-f�hű�#��;n��`�B���f�H�) г����#����}�)� ��bW�':�[!d�|�� "Oʄ���&����%�������O4yl;1KF$s�n��\����
\�asHc���fX-�M;��?(�x���O@J�L)F�%�sk�><��d��n�O��䜳�N�p��o����a��)2��Og哬km�e	Y. h9���%m��']�`S���,���fKL��,��f�ɛyG4�:҇�x}^Ic���4����������S�'G��I��_�[ZH@P@�<^�4�ȓm"��Z!4�]���C�|���I�HOyI״<�h�f�n5c'�����	��l�	��p������	�� �i�Q���l��`C׻I�NmӦB�{�(���f��?�6h�/mF$T�|&�,�u��JC�e���ג)�=p%L	lW^]�c�-�?ab��W���>�O��#2�$-]t�1-�p��'�Ir����|R��6D:�I�j�n
 K���y�.ͺ6Qҁ:���Z$d����B����l���X�킼���#5,��0�r�RF�6�s��O.��O
���|���'���?I%��;B�
���P��3�2��F�6
SpȪ���g�Z���I=T{�HؠK� �FŸj�us�<c&���z��aj�l;��˓;:J��5QpJ��X�.�K$.�2��t��(�M#4�i��V����m�K"��#`�3#Y�K7_�9N����/�@R6���sc�G�/o^��<ɕV���'�B��	mӨ���O��Xp
џl_���'Y�mǄ�O0��� ���O��[3p  #ǂ>k��j��O��ZR�E	v������ѬQ8��'b�J�J�vp��Ec
�L�R {ө�<h��t��ҌF�5�A��zQ�W���I��y"���?�g�x����QX�%GK��؍['���yr,�`$ֈZփ	� ��f�Ɯ�x��jӈ �1��p�FI����{�&P� �(���_�2Tl�ӟ���e��"��7N��3��0�4��N����v�
��'#��W�3^v�d�b��9 ��Y'�~�*�|��$�)�uq�ƨ�m�T��P�Ȗgc>�듫"���K#\��b?�@nW�.�T�*� �)M��`<}"�A��?!�|������]��2��JE���;'"��yr��	�XY���<���A�Cƻ�0<Q0�I�F>L��tĖ\�d!����$^��`ܴ�?a���?1�G�HĬ����?���?ͻp��,��  ��*1�s�Y �d}�yT;��<	�m�XG|!�́3��X �cK_�s?���ɟ.F�+VEPW:�"�M`�
��J>�b�MƟ�>�O8�XR����:�شʟ�}��HP�"On���`�|�$���	��,����9���ӋtYft�c'�3u���
 ̔;?~*���Y*�=������I�h�[w���'��I�
L��d��e��`�J.�����']��-+�p���@B?�v(9�/ʩ8�@l��D�gd��#���f�lH��'���X�#]�^�޸p������͢qk���?I��'����e`�\��父Pj�	�'J���)˽)b���6�� Gx�1x�y�H2�	=]d�-�ܴ�?Y��\q�����ۄ	�V}�����?y�䞴�?�����j֟�?AH>��	\e� �DW�b�2tZ�Kx8��RA�4�I�J�5]�S
�Y�3 �81���$�1tMRc/��pC,�(P	J6yN-�ፂ -�!�$B��ɰ��Y�L"y��Ǹ4!�����a��Ț�����,�|m���2�I�zbq�IƟp�	U���L��#�a��Dآsh�I@E̤3`��'Z
�4�-"� F��y�U>U�OZP�s�>s�PE��'M��H�J��3��A��1!A�*H�����͸(&H@��-N�o�"�R���(KZ�e��]�I��M���i.R�	���*6@�)f�5Ac�^:bF1O���<1����V0q#$�(p��s�Ϯ6ax§x�0EmR�^|H�J�I�8H�`���/B�(�zX�ݴ�?9��?��@�Vx@����?y���?���iCX1�'J���1n˚e( ��yB�Ɓ��<)�,�WL�}��X����T�g#��牀#�L�`���2�\0���12��1J>���ß�>�OF�`2�H�g@�t�eƬ`���9c"O�t�wF�v\.�X1�@�ڌ� ������S�'�"UxF)�9�<`��)�*%0�����H��I���IƟHp^w���'��)P	lY$5# ���5&�<3�KڟM�ddZ�O��B�B�+Xi(r!\9|Ŭ��T`�qI!��+�4u�Gd�eT�Y��JW��(��'����  �!���9
�q���)��!0"O<)5-ʪB��$�����W���S��DOa�O$���C�i���'Id}�b��$8.�L���'9D�e&�'f"!Ճ(Z��'r�)?v��|�,H�Xd.-�-ɀ7�5Z�F��p<�F��n�Fx�R��Cm+��	�ф㉌r�$�^�9d�2�e ��N��#�G3o�B�ɶ&��y�Oٲ1�|��I_+�C�		�MQ �&����� :w
�c�c�wܓR�r-�ٴ�?)���	�g�P��_`��]:P�b�	�,�"`t���O��z��O�b��g~�㒙!<�Ҧӷp�<�zv+Ÿ��6X�l#<�C���c5z̙��Q�-�C��]��^!r����r�a���`� xJ��Ͼjk!��a4�C�bܜK��X���0axRf#�p]^��� �5^������(6�jT8ǵi�R�'."�+�0͉�'�"�'��w� �d��7J�	���B�&���$ѵt��y�IҘ3ya� J�L;N]s,ߧ��'�p	*�>�}�DːMQ�Ub�b��g�li�y�⃝�?�}&��+�J��
[��ɰ�
��z%A�&D�\�#��$2����CG1�V%`WD1?A4�)�'i�p�B�W���}�WF@�Q��B��۱	,��1���?���?y���Z���O>瓗Y�F(�6���A��:)�P����pŒT���G���Y `֋�]� �' �94�E�A�)����A��s�� �µ)c�`G^��F�O�e���`�de�Ĭ�KV�8�4J��B��)7�"t��#q�J��� �*��b�\j�}�  1�X6-�O,����.*�t�V����8Q��e@
3���d�O����O��f>iʕ��O,�O��&�L&J���20��E�(���'�����"�۬.Αǈїa�@`[��L4�p<f��$������ QC�G��P��$D��jŊ���H`6lɩ{�&lH%I �X�۴��P	��#+�fA�-� %Cd4�ȓG�<I���<@� i37J�1N3X	��v�����3�ub��O����V�|��B���lXPtZ�O�,Yz��ȓ8B$���6[/4-"���<G�� �ȓ5��~���%O�/�$y+3��T�<�!EW�A �*g�F����WKJ\�<�ͼ
���W�����A eG�c�<I�HP3bE�e �O�hȍ`�b�v�<a*N'���u���:ΪH8�$�v�<A#��L�����қZ�xQJ��t�<���P.8���q��.H� R�l�<�WiȈ"��-�S��&�^�����q�<	���=�5@�hԕ	�:�0�x�<�Q�Z�Gp�=���&�����u�<f�ف.�@���A"�����'\s�<y��"l'P�9V�C�5��P���Sr�<і"3D����@� y�����d�<��l���$Y�ɕ=(T�,Xz�<1���|=(ҩ��|4�΋v�<��kѩX~��c�M�I��}0��Co�<#
Uj<����(tw|(�&fCS�<�FAvK���U�[�$�� L��yL� ��T�C�H0r���c�ć�yҌL�Ũ�B�H�d��S��y�)N wP���63Ҫ4��@�y�O�*�T=�5�;k�؝��&�y��O;]D��'f��74d%�D ل�yҊ�~���P��5\8���Q ��=��K������"3�hS�JH��j�Z���+>��$�ʟD�Q����MnZ�q��4$p��o՚��C��\}�����$G?>'��L>aC�O��Y�?z�$y����d2n��ɓ%/��ɫt�ΓO���OIdݨ�!�o�^�]�=�0�����;.c��ajD$�g I򉖡~ʟ.g�<�����/�j٪��D�V���B9���R!.YZf�&Ke�qr���6Q�� �9	�� ,�����h�Zb�� ��s?y��Oh�Ç`yZw��!��xB�XM��_ ,d ���	/Ĉt�@���N��F{ �#Y�n��u�{ޅr��	8#rm;q	+�>���XߞO*|���i�u	���=J�j ST��|~0Xf�+��?B����-P�Kw(X��'4��'��+��D�G}L�He�~�T�J5�Y�'%�3A+��K��PQ#��+���0%b$��'͆�5ʄ��plT*V�;��m���L���}�O��}�,�}\�q��&P�h������9 X�r��1y���c��۝bN�⟘���8/<���&��)�� /�)��I8�Q��>�z��?=�j@���;(��U������7��o���Dy��{��	�Q�s��gN��fu��)&On����'��-U>#?�cF �"�7
�7�S`�Y�c�XbL�� E������IRD1}�!2D�+����8cm�#r��2��O<��өm~Lps�*ʂ� � �C�e�pɰ�A�L(t�&�-}�&�ZBf�L���ČR�*����K�
�����^��� �%L�h��[E��c��'i���f)"����Gq�H`�g�e�]scM�()��X��*�nQ��>�1N>�����[}�%ȔRa�W�ġS:[�:LނM+�H >EHH4��:Y��ywD,M�0��k�
-�΀
r���'I���f�'`�h���Շ1q��hB
Ֆ���*ب{w�O��2��=����V�A(�(UY��>��H�"���,����,L4�%2��3nrQ�<�"���lw���$\!tp�$0�γt2T@G�B����CC\�X��YK�/S%4�@�#@��x�Ĥ�!�-?yÀ��'�l�k �Âݱ�%ݝTh.9�,O8	r�^�4�R�����[`�e���O��ٶ�6L��Gđ{tn�3�ɺ-�Z`!�����D�C�>Y(O�x�??��O�Y.:Ÿ�K��b�4Y��_0	x����C�K=�8(��D�/�$�O
5}�ݛ�@3dV	R���21׊I�O�ʓ%�E|"AL?<w�i�����	Ϧ��p��U��P��Y�m
SJЦ#�nu:N�
[l)`Eۤt��§�$B�si�?gFS��N�'x��C��Q2�.,���� ��NA�[m�Q9t#�&y�����
3k�R�	��2M�c���oq�1�ڴT7�������rN�G=j��a�ʜ��hB#W�򤗡j�~���������A��z"<�Beф[l�5XRa//�˲C��m��ɐ�hY9�<�t��F�:M�a�@��Ԣg7��3�F<j	��b+�CH,xr�Z3�hš
�s���x�,(T��5c�"��(\�I@����$L�	���Î��Ѣ5�Dh��ŦOsV�ц%ӁL)D,1�I�H-z���aΊpZ�e8�!��e& ��;Gh��T�_�EP�`�$�
�q��I e��kUśAVL0B��p��`aD����O(��CU�o��C@�� ����������di$�Vդ��sL�/>AyS�P�?����'J>y� ڻr��{�L�*R`�;��d�G�\إ  _,S���3f�z`Х�Q��	`�U;^�9�g:'�1�w�3�~�Y��U�����Ԗ_��n��S=ڍcR(�������%��G�
9��Ot���ɠG'zM�2ʙ�z��]��JJ�4��lr`-(�)�F8W'ʛK�ZH�NB���ϓL�nl@�)_��Ha &=�di�{2�^f������&T�+�[>XI ��>Y�CV�k@�����L
/aTe�S@�<�,�->̥�NE&{u UZ�KFa��jr���p��xWJU+~��.��f�9	��ؠ7%D���&��>a�yk����^��@sF�T�7�����mW0��q�'Q���D|~2�;5N�f�U	]��p1% R�svxy�,)�\����K���H�4���S���l*Yh�a�;o��h���T���DĄnSh�?�ڤ
����<�âX
A���:&T	�O��(%N%�2�{�U�TR$�q��THS��DUQ�.��,_�5��G��Mpj��nĄ��Ox�]9�M����}+�lJD��
�60����T�MI%b�#;/�i��Z ?;(�E�ʹ�f8�O��5�4dj�`��F2g�R�J��S�_`��	Ohl%mza�څ6?���D�}r�&$�I�r�؉4�|[`IZq��!;q�5+�	;}��N����'{��ğ�'P�0��B �	��c�BŉkTJ4 !��a�$f[�T�<�ө+�J5�;dE8�f��vB:$X��S."քn�J�*��B�<ye"Sc����б8���ٹG��t3@��"<Y$D�#�v��3���b�`~"�A**|�Q����v�,�;�]�O*��B'A�H+7�S���Q��I)3�C�wO�����Pn�ΌZ'�F�_��t���̺$a�p���܈5�n5�#\�^<ȭI�|�#]�Z4؍	��_'ޭ���#
���`+�&�|A@����fR|@B����<���M,V1]�=�V�ͳ ��ɂg�5 �f�QB)�i��v��)�+o��KPM�n���?5���(�Ԑa��ב,l�Q�!GEl�0���E9�~���T>��K���a ��\j���oN\v��@�+�'Vax`�݄���0O���c�4��<��C�B\��pfp+<URn߮��'�<TPfώJ�Da*�mHN�'�>aQ�
V�n���돯l⤣��!@�� �����ؚI>!���[2�٘�.^ZL.@&�_AA&�K#*ݪkZd��cߍ�$lB�t"ҬDy�"Ę/��E�"g֟Z�R0�%�y���!$\�����V���d������F�W�R�B�X�l�=ydÐj�qB�.�J�PCqoa�n��p �c�c�,�� e�D՝M�� �i���q	fiPs�\	zM��6����h�&u�H�É}��,�(��tQb��X��]�s+�;8�����D��=�go��2��>�,P
f�3�<� R�m���
ވ<�p�(�a�	��'��x�s
,���8��O��&����/ծ|�
�����0R����'���O��͋U�I(\��)bg�)��Y�(`cǙ�>b��@#�8A
�Y���L�'j���0�	�`9���ȉ�^���x.O�Ob�M�� %��I�AF2��̇jr�T2r�I@U
��Õ|r�Y0 �
���-��NA|y�"�_�'@����(��!B�y����e���hM�4�T';(� �WQ�\V�Eq�4O�°D\-�5��_�xC҇ǝ`��e�s��v�Q��d�x�"�H6z'�����$ɥs��!�7�f@z��$��E!}y�&�]+@!�4O���&م3!� %>˓P�Ľ)u�D�R����ƬQ�L��Q�}!�T1D|"�]�t٬�3��Ƹ76�)PCMܸ?���S(G`��:�G��ԭ'��8�O�0Q\Ԭ�׆��<�p�c�R��$�& �3OB����7��@(��$�Y��8��P�W�R=�ab�!�uˀώF@D�͉� ��<�H>�ř�`9�=�JK�Lx��c Laܓ^��3(Es3'��VX\�OfQ�bn_.A%��P��e	����Sj!�Յf���<w�h��o�=�1s��wz~`�wϙ>��Ae	�1����t� �7�k�i���t'D1�4 )e�ڻ4�*��"��'�T����?	��e��b��*�E8��;aMl�h�@ZCV�EC�L��'�OV�S���<_j*�X�aT�PP5c�iE%x�O:�'uB��4"Oh���'�>e��iA�h�|Sa`�*y	Ѕ�C�I5h�.���q�{�E��	*�ɐbX}��n���(x$� 
��9-�XS�@�!x�Vۂ/ڬ���ă93O��q���0Pp���'P�I<��O����'����~��_����&D�$�1ᤀ
4�v)����`@ G�:S�
�>A7c��z�́�t9��	@�B
f�X�+���>
|�س�i�X�	]?Q�KԾ=x�S��t�1VӘE�c�]�N��mH#tPH�>� 4R�XLai�=6��$^T�$z-��gI��[oJ5��a݀s�����Jѿ��$�<�'*l�xW�QMk��=�B})�L�T�L�A� �(6����#ķ2K�Hq�<$����[k����0E�rh�f}��I4��6������1�W�^��Ʊ�$�b`G{��_�t�r����?CJ����K�+o��x�v�'�bI���>T7tԢ�ܾky�Q��#��?j�Aq�I
>�칒O��yǧ�8����b�O��1��%|*���lX��]�G��	׆ڕc1����BA��Vc��R�㐅�l�',L;*��&����j�H��@s\h���Ѥ/$���$�ړOVU�B�O�p�q+D��r�Os^�!���!�,̲4�G�F�I�0��>Bx�6���x�h��'� l)��W?Ȝ��d��;$�,�'Y~��T� `�!���G|���^���I«	�:��+"g�	K8��d��56��%��P����!��)�������D�"�*9zt��eS�)��t<�t�Cf�Kϴm��&1�q��@J��Y}��M��D˖{�(���Ew��K��D�@�H��60m ">����3)֘� � )�0������^Yl��`Wˉ�&} �X�Ι�Zg��%v�d����C�~d�y�D\����6�m�FXX���X"O�hUȖ+d�t�� Z]�t�O�3�$	m ����P�&����\#6l�!�*ھ�
�����wa^h���V	/`��Ղ�'@Q~��&ZZh��&���y ��~Yz�4!s卋Mn*y2W�͏O�4����w<�)�����
Cm�31�pK�@G�Zۜ,rrl	F+��2�'�t嫱��gGF�b��O��qI��)�R&D�'7B\z��c�ѿW�`b���g���S`a+hR�n�rq!���O�J\6�Qt�-4c�a� �$"�Н��mS<W �	D8&s��$�3�I(}պ��$�Z�I'n&jr2���/@�+^�Jv��4bV�$#�'T�e�'{ Te�W ������+��Yk�,�HE�9���*�$0�O�ES��ĉ���U��=F+>��4�'IJ��E),�|�a��ӝ��DQ���O$sC��jh���
�)�B���'���@�K��6���4�9-Q� �D6^h�pV��Q����,���݂WN���0�>��S�O�iy$&Ҁ?� ����5�.m���$Lm�E�o ���������/��q�p#сu���RD��x|���'	�y�n�ʘϘ'[�! T��3J~�(�Ӂ
-�H�'�,�S��U(Uj�O��M�&�68��R�� J�N�7&�	�V��d�%������18��|�@�?.�-+��ؕ;�������qOfmz��'j�p��`InF�ݓ�ߟ|��.^���d��*Ec���jD
P04C㉼Z�P�#Eш8����5��=�2��i��)��V=���J&�u��,�禅��hU����;.�t�1K/D��A'	[����u��3ytJm�"d^;4�p���'��<�C�Ķh���g�'K"HK�K�U|`� ��&
�I��I=E���FjY$)��P��)n�D����  3��x�
�@娙���'4�z�"�֞\#&B~N��Q��$�2FN�{��%+Ϯ%���I�0J�|��U�| Z�g���D�!�� \����=:t���i"*ɚ�'�PݡGO@�:}��"���	��?�����V�i*� _�N uX7���<Q���h�b]�$`7��-0"y�<���p6����Ƅ30;XpK��r�<QW��5"0�kщVD�� ��n�<)� ��O��q���Hg��aNTe�<�l��)��t(��g���S( m�<��O�<;H��$I��`�8��i�<��'NM/�Pkc����0���I�<��'����x���T�#��=0f��_�<����	S�ʃ,�f�p��#`�P�<��931�9PŮA�ڥ[4+PK�<���9~@4��m@�*��𐶧�o�<Q��g굑2�J2"(a��Uj�<yE��D��������`+N�<qF�[�I$x��i5_&<�@gE�K�<9�Q�D���Q�

/�I��BE�<�ܨv18���X;m�H�#��G�<��������`�hz	��X�<ɗ�\4f�z�2D�=��4y�SV�<�Ei��**�@0
sS�퀡�U�<��G�'w�
�R(Q�=���a�fW�<��|Hٻ�`_.���t&Cj�<Y�T:��Q�BC,�q ��<�U�'It`#��0��0�
|�<�얻Rd&s�Te�f�3c�CC�<YS�8���͑4� ���XS�<���,�33�Do��!jӊGt�<��΍�x:B��"��v���#D�G�<�2"�'h�p���.�,c�̉�o�C�<i��G�"�p����*P��$ڵ�S�<��HU.%Ȕ
$r���	�d�<���K�F]���g���;��z�.�u�<q��օW< �痤�����o�<�3�;v��̉g�D�/���C!�D�<�t�n!����#�	l�4����C�<&O�yP���o҅g"�x t�B�<a%��K�~�ֆI.,���i�<�4 �?3������>E��]�R�]g�<y��/#�4��V�]��,+(P[�<���8 ����@8��q����q�<��#(i>(`S�ԙB�z�"��l�<ѣ��>.t��ؓ"YM~h����k�<�DD�"�r��&�]|�d9sӌCe�<��c�%a�Eq槂��v�
�O Y�<�fOέ'\X���5
���*�J�<�g�I�s`�����Ӵ���"c

L�<)�NM�5.F�A3���n�걂��E�<	U�ΐ�V�b�0ad��p!Dh�<ɦÄ!EJ0�eh՜7x�Sҩ�H�<q�K�|*]i��]�:H�s�]j�<�b	�+֜�zf��N������<)��eʠT�%D��G |r��RQ�<!f�P�"�J	���Ω!����P�<!"l)�2�J�:X�r��Q��B䉟:[&D��mߦ2+F�R�yB䉏*V�i*r�� o�P�z#o�B��P:N�+�-�!�&�z�o�zB�I�}�j�y�F� "�:eH}�8C䉲>a�8'J�$H%B��L�8�>C�5G�0A���$#9H�R�Ë4�zC�	H���8�7�b���ldC��"�tj燊�1	^̃�&Z.>�XC�ɛ2�E��wd���,hq���S�? RL(�Eb�"��E%O$)���B@"Oz�Рj�"+e���C�!��,;""O�㔤�+	�TZ�!D14� Q�"O�2�t�aSc��N��	�2"Of`��fN�s7	���f�പ���\�O]ʭ.-Q����E��K�łC�<��/�v�Papj	�y���+�!�|�<q��ڛD���xg��*�k3&^�<Qe����Pp�(c��ጂ@�<!0D��c��d�bǤ}�Y0w%BG�<ybO�l�B�k
�!�ļ��Ǚ~}��'�`}8��Uhm*3	F�-��)����α3���2�mj��Z�A!�P
I���3�@Z�q0�L
 џF��)H�
�����|*J�A4,���yeN�u�DI����t��`3.A�}PB�	�F�޸S�#_甉A�cJ�=l����q����o���\�"c�G��l���;D��9��9bT J'BY�1�|�p�:}B�S�Of�]����D�Ր��� ��1�	�':���ʗ�%k!�#(��C�����6��<�S�'=���aS7A�|��gҠ$ϼ��aPʅR��U젓0 �O�&y�<��7�(�i�HC1N"j)��KH��܆�[n4��w�ϸ!o��Z�n�*�X���?Q�'R�d�K'y;bX����s�'P�	_}�|��_�D��*��@���A�υ�y�)X�K� 9��°1�¨S3�ٓ�ē�hO���q�[)��!f\�D��@b���|�O����%��Q;��XM[��		�'����w�� 
_�B����'b,�	�|�*��
X�>�|�O���-ھ㐅� Zj{l��"OLM!$ۜv�
�{� FOD�}��'1R�jFE�e�t��Y�O8��'/�"=E��D�V����^>K/�X�q�O>�y�D@��Mp�% t����K�yF!���U7.� ��`NrqTc�_<!�$	V�����9�ԩ����T!�$�N0h���BQ>/��t�5��&E!򴲘m���
Q��Ui�<䠠�ȓ��ȩԨ��9���(1A�D(T�=ۓ5��$Hde�JsA3֭
�2��l��I;�}��KH<9���2�G&�p@�����+֮�	>��|�i\���E2�Ӭ>�.��!V8e�2�nJ�{n$B�	Idj�w����e��/	�
���$�>���]�Ҟ�p��7x�6�9�+K}�<��bT���f�Tx��z���N�<)��B���"��	:�����K�'��?�
c�����H��)������f?D��h�K�5M� ��Vm@A�?D�L
eٝ>���*�g�^$r�zQ*=D��ro�3% p�V��"X@�*Q-(}��OV����1EߊL b��(II|A�\\1��DP�l�́I`#Zb�4Ii����1T��D+s�¡s	�����T��џ��	r�OP���B�]g�|h�d�
h <Y�',�pA-LQh�j_��	��ēXEp1%Er$��Qg݆fG0e$�\��� L� L��c�,^��c�\�x�B�?,�z���g��ۀ�L26B�	�X��[�rk�bå_tڽJ�ǂ��hO��퉲��%+��Dpi*��6��:�B�)� 6\�P��F[��!�e��%�|�f"O<���I�1�:�����Z�(P�"O�}I���  \�T��%ׯ�3"O�y)U�^�d���"���j�~X�g"Orp�s�\<I����ņ	\K���)4�hֆ̢ �~��䊤8!ZTЕl4}�i���0?a�4�yr��Zy�ꋣ'��q �a��+>��)R�V)�yҤ�a4�x�-��&�$�K��ˋ�y��]�  m��s:d�����>��O�T���9��$���� �.P�s"Ov���l��B�B��E_d�R8OF�O��p/�'a7��Q$�3')�����&�0���JP@d���Y�Ҳ���puB�ɨ:��#<E������ıW=&���F��+��|Jܴ;���B�3�� o���/F�$5�Ob#�	׾h)�
ujK�hԮ��"O,,;AD�iU"�X����1��D��"O����ћY��x��ȣ#�&D:�"O0X;��Q�fɴC=��`"Oj�!���+؀��4��<GV�pXq"OV�eJL+R���d�$/K�Y�"O�h�l��,J�=
%(�<+C�X���d$�S�S?\�\���K���i ����LT�C����Y��
ͩ��� r�Ճ;�vC�ɺI�H��'��11���tG	&t�B�
/�[4�T%ad�8`K�vC�ɵc�����^p�<�U$%`��C�I�Q�(��6%��,�j�$�L��B䉌-/d3s��_Aj(j��ا/^�B�	=c�|�3ƙ���"0���B�I�3ݾug�I%�t|���dz�B䉆r�$�8��ހw�\`�c&%��<X��'���%�ĪKL�z�j!0�r�<�@�6��0r�	Շ��ⶫ�n�<�I8����wl+S��uJ��h�<�dn��w�0��C$"ǄR���Y��'�}���C���q�<��E��'G��X4�I�����0����'#>����,��@Y/T�8ׄe�M>�����i����Z>��;�ğ7ob|��I�<٠ �*m�6�k 
���i �M`�<�D�L�9����HF4WL-� �]���?�����GT�h�c�R�Y��f�~�<Q���$���c� �{f��kU}y��)ʧFLѺ�$K��L�ҫ�� |�ȓ:�R��q�(��d��4]�5�=�ۓG��K���2J�f$��
銵���?	�@A&f��-Qd��"!� b���<�q�T�U`�#a�V�).�]��o��<��)��	��DR�fVy�@, ��|�<ѣ$P31bQQM�"$H��n�<A�\���ҰKUz$!�O�R�<y��_�1|����ѽ8J�``��y�<�7&Z9�M ��;[¬� T�M\�<��	�#s96q�s�M�I��HFA�Y�'�?����Z���+��B�$0B�k+D��� �A� �4S��!��)*D�P�!�9d�R��g$�e��(D��s4�цy�x&B�C	���� +D�,j�#�nY�@��K:Y(D����!��m��;���M#�D%D�P��ҝ,�Q�%/إ+�A���&D�L: ��"��B�b�_�Ȕr �*D�#� 3G�`�:��[�":�P�5D�� LUa2��=_�%q��-� ��"O�t0!'#U>�{��O ��4"%"Ovh("!�\uL�xbC\�C�"1��'cў�j�:*28���D!=�)(!�6D��"#�
���(�0�iD�5D�T�7��!-* ��e�$y����"?D�$;�C!��9U�[�h$�AsI;D��	G�eQ<�t�y��ً�t�<y�-�l�#�'X�x Lʇ��Z�<9���u��-)A���vlv9��ɐj�<��E�="ma�F�,zPX8�Ge�<�4"ߞz��@�6)��x��SJ�<��Ń��Ɋcd®yc�#�k�<���/Fx��6a��=a>�+��p�<q��O��٦�[�MfX�� @p�<9D.Ϙ.��paC�(}ڍ��Hi�<فE�9�\�d���UeDc�<q' ����E�s�ă,���zwQg�<�3�Y�3�<$�TA�5�b��c �c�<��ͭwVm
��2I�P�I�@�j�<�5l#s�T��֌�{�v@"P��h�<�3�I�~m���ƪ�8ږ�[z�<Q�+�*JE��M%�dt�eIx�<IQƐVTXx�꒢-�C4
�n�<��i��O*p@��9�����D�<!�n�:(�D���(^6%������@�<�Q��3�$��Ç�o>�<��+��<y��˱�~�Be�0i����� |�<y�A
#dO��Xӈ�-?�V�H�I{�<�2��" ��\*��B+o�Ț�jZ�<�Q��s �@�Įδ�raa�{�<i��փp�hA�[P&�*��\}�<��֩ �d�@B�I�͉w�<��It�pĸb��86���&�^�<ɣ�(#*�9�FS3����fJ>�yr��?CK,��*^�r�Pc�8�y��ڒt,���Z��4��,R��y�nB�~A$����G��X�ˊ��y��͠W�漪4#� 6A6Ȱ`�4�y��t����E�>.�^�0����yOØlpM@u�� ey �4�y2�ӌl)ܪQD
�-��1�f���y�mѫq�����v^����Е�y�![���B�Fq���y�cЀ�y�d��LA3c
�]�DiQ�%���y�j�1����r�	W	�x��M
$�y"+�,ef� 	J�T�����F��y�l��oʅ�˗D�e�қ�yRG� ���@�
:�lx�.��y�*ȟL�*����M +_4�����y�lGGu�!���%^h�3�y�C��@����J���Д8sč�yb��/Y,`��xࣲaĘ�y¨��zR(8���4��A8�lF��y#U�&0�Ma�� :!J�@�)�y\�]^�9׎�$]��z`�0�yr�Y�[�z��̈Aq �RgW��yi�7\e�1�ԋ�'4�2�[�䁽�y2�.s"&�) #Z$1(�0����y򂘘�8͢�O#T�̀R�l[��yB�TQU�4��M�M"����y"
�"m�N�h�AҶL*�Hc�b4�y�/Jl��|����K��I��H��y�W� �u���n�8� W	D��y
� �����	@���@�͡^Ք�H�"OrLR��C�I���aH�+�f���"Oƕڃ�	8}���l���2"O"([�.*Y���C��#D�v<I�"O|�'BR>��G]x����"O��B�
�$�)�,��4��e��"O
�f�0ZB�T��,��H=��C"O�H�Q��*8[�Q�4L� =����"O�AB�������̞�3���&"O\)@�2 p��%G���I�"O8A�+�3J��93��2B{๺B"O	0��͛"ު0
s�-����"Or}�@#�^
�0����T"O��QJ�b�tP ����w"O �8%J�`8�!��DrP��2"O씰R6Z��  �H	lPЫ�"O�0�@�6�N�b�W>Nz� �"O(I㄃��7�
��B.�	+G�I1"O��fG��W{tMǬ�=-Դ1�"O��p��q�%����<G�B�"O4������2�H���,M)FD.@��"O�Q�F�P�yY�D	@�;2�*W"Or}I풍�t���mO
m��� "O����� �&���܂]�.a�b"O�|a�y�@\AeK�4ʲy�"O�	��E������I��y{�"Oƍ�����}����F�8�:#"O�L�4ER!�h y� @8T���["O:5�1,�@�"��=��k�"O�9�Un�
,F��1�.Lۨ�Qw"O��B�Ĉ$!+"�B��Ҧa��8�"O򉪵�>}��t��C��:퐝�5"O���F��p�41��F2"� l�&"O�ШbȖ�%��d鈩;��"O�Tї��ho���B��@�����"O`|i$c
@U��B��Ix5�"Oz4:��&g e���Z=��@"O�i�`'�)��V��U�c*"�y"cr�4�f
�NBЀt,��y�-�!`0��g �@t�u��ƀ��y"�ԝ\	�M8AM�3��� �B4�y��L���y�d���NH�y�EW3AkP]*�Α�kxl�����y�,4��|�uF:glj�����<�y�"̸/�V�3�3.ո��"�<�y�CW6\�����*��DD�� �y�F�o�܁p0����QHG
��Pyr+\WFJ�ٰBE)4�Y1�N�<i6�F�0�|��
�'N���a(�@�<��k�:�aǤE%xJ�C��s�<���`���T���1��v�<��E �bu����	e�VZ�<��B̬L��x	q��'��Y�6ZU�<q�f�>.�C�ω*�41��*�Q�<��DD�)ȹ�ff;�x��A�C�<Q&	�2���咷M	�X$E�s�<	��A�k�2��*]09"t� 6/t�<A4�Ȱ�[&�O���)bE�Y�<�$hB�������БXc��g� V�<���0�N(��,��T�|�3���Q�<i�bK�0(��w�ξ_��c���E�<�eF�?��8�dJ�,%�=ðg�F�<IO�K�A��a�O�B��p�NB�<y���s�i�R)��%{L�:��|�<� �qkc�[���ݙf%�P�J�"O��rp��m��8x����i��|8�"O�WEI�5A3Ҙ,�"���"OP`�/��V��$�%�1k���"OP�S���7O��q���cP���"O��#ƭ�J�� ��<\؀"OЁ�O@��88�C��!|�mT"O�aWF����1͉4v�Uڱ*OJ�)L�OjDQ��%]&���
�'`���f��P��Uaَ"'��'��mbЩvl���"X3Ѯ��'�
���LZ�����lR �l	�'�f��5�^�&ن��L�'B���'�=3t�¸$��\
QaP�?�8��'��]1�� T���S%6
സ;�'R���§�' 0��/P�z I��'4���A,�LJ����I	o��k�'챩�Dɤe.�U�B!x�����'����1ň'/N7��<&���'_`�cr��4��i;�HW3evٛ�'��`V�ąJ���qsĝ�}R)
�'�z���iR+�`}B?x����'���W'���ע]+EH�8�'5���1���h����B��ܔ0�'&��zgm�;+��rG�
%����'��eK��[�	�>��Ř�dvޱq�'b������9���@���a6��'ŖT#��ޕZ2�*k��Y�X�[�'@�JU!Z�^W��
��ǻ?��dP�'�z������8E���5�P��8Yp�'��j2A�Fr��%FU�FP��'��9���P)m��3�Nɳ83z��'�xe�t�W�c�pAH��,�L���':t���T�b�z�y��T�4�2���'��& {K�2U�`�z�Z�'n�!�­4g׾��Ϟ�[&��X�'i2+��;P��IBdeW�p]��'!��9s��|V
>"�2Ց�B9D�@hG�C�'���YWh��#^T�	��!D�HBb���]Ғl�%�� �N@ E>D�Л��X�A��ɘu�Oi���;D��"��h��x%��(�J�A'�&D��0W�ʘm��1��	�:�:��q�!D��y�-E��=��G�)�u�3D�� ��h�Lɓv͋�{����i2D����Ç!�0 �(2��P�$0D���Ro
�b.���,Z�P �'/D��)��*��"%�ƹ0���i`h,D�4ҁ��x�DU0�MJ��M��+D�XR���u�2]��*.C����B5D��S�e]�U�"�����%Rέ
��2D�8�w �gb\Aa����j��.D�LP5��6���c7�^.����-D���%%�qؒd߈$�VE@�+D��B�+1� ��F&�/.Q�@��4D�ā�AB�j���Y�'��$�¤��=D�6o_�O2芦�
]�6�NR�<��dI7n�HR���[Հ�AVw�<�$#T-_D��B�C�LQ�f]k�<9be�K~J��ҥ��԰!�Se�<�7��.����r� ��҉ �Ag�<�e��\Z�`�\��2��j�<���'�-q�o��W�v����Fh�<���,�08A�%bp�(� �b�<� �ĺ�&p�F�0c��I�0�B$"O9A�%�����F��25�
\��"OF�s�畆{>�!�P��Y-jw"O��z�fK-qv�S����	�
)��"O.�B̝?�����X�;l��"u"O�HW!��(vt�(��ę)W�l�"O��� F�2p�bCT�ڋ@F�)s"O ���Y�_4L�)`�B�0��=b"O*#��Em����Lؚk��<�T"O=R֋]�%΂�8�ˍWr0�PS"OЬ��&� ;��dk��*���	�"O�@S����[[bQ��W=�Ƽ�""O����0�� �sraɣHoL!�d�:yB����
2uȦ(ڒN֔K!�ĝ�{�@RF�ڂ:���	��\ 	;!�ď�I��(���"��z�"X1R!��v*�-$nT��!�!��Ý_A\���N�	�PA��6�!�D��R�h`����]�FZ6r�!�d����2�
)(s�0��ս2�!�$����s�bcԉ8e��-�!�d�yA�9A�LR_�QZ"�sw!�$��J���A�A&n}K�g�!�Q;������{2/8;�!��&���nUzb��I�LT��!�(Ij�
Մ՛og�`w?�!�$���l��m�T�p�鍵J�!�$�ha)v㟾� �3t"�!�D�7<�� 3�.-�����)+�!�ţ*�$	��b�A�� �EG��!�$� |yh�SD��|��M����=L�!���u����	B�|�J5��!�ڐCpl����V�0d�E�_{!�d	@x��5�_�D�̽�u����!�DҫR�8C��Q�u�P0�tMŵq�!�Vn�<�J�n )m%����B"O`7/��t��,˂_�r�>$�V"OnX�c�H�C*�6�p�P"O��� ���B�6|(r�$L��9��"O�ö�A)nΖ���L8g° *O��p��T퀅[&��)V��]+�'�~�R�,�$��a2f���Vaޝ2
�'t� �Wh�)Yoj���P�I�x�	�'#=��#��J�t�S���F)Pp`	�'�R`��nԎK9����-/�LL`�'MLez��I�f�[C��8�"�8�'��,��{����c���X�� B�'�r���*�Qn���@*�:O���p�'��c	��.���r@*�{6Щ�'Sd�Yw��#'R*�y��v>x ��'_ (�1�ۄ	��vc&Z�f�p�'*���A��S;x`VhC�S&Bi�'N�A(P-C"RJ�m�BK�|<ظQ�'|(� 璸Cp�LL��'m�@�va�L��9iR��&<�2�q�'�>$+P��$V~���i��g�ȥ�
�'B�dQ��I �$H�q)Ѡ4�d���'z�<��k�9I��̠Q&C&V�$ ��'�*��w�w�&�����J�$s�'	��S�U��h� �֌;�:�'.�Hɖ�V���Y�389�'��p'Z�����V/U�#�h�'B�h���j���` ^�zd��':�ebֈ��N��80��K0[��� ��� rx���ʼ<�t%�W�õ`�,�h"O�Q���We�D��(��$� �1"O�����X�p4�C�	}�r"O	yGJ� 9p����	t����"O�!�Gس+� ���E7�T���"Oz�8U:x-�)�3�ք1�q��"O�����ŀU�x��TT�t�E"O�ՙF��B�ґQ�A�ED��H%"O
7.�v���5 ¤Dx�["O^�K�j	�u Y��	"/�RA��"Oĳ��.'�����C��]�\�Р"Oެ1���c���1�J��"O<�Z��L3qi��!e|�x��"O��x�C�%&�2�%7�.��e"O����gĵY���!�)'��Bv"O�8�g�H�IK�J�8��"O��0� �n�=Б�D�&�u;�"Op +R&Ro�p�z
8>l�s"OLI���т3�D��P�E�_��)3"O�U�^�M���Ѥ�nS�ݻ�"O`��T�W�~l��ۃ�	5��k"O��*�NNst�@�BɗE�pd�Q"O���$�'Y��)A^ �<���"O^, w!T^��8W�&¤���"O:aj�k�G9xؤ��|Y�@��"OB�D��,H��rf,�I��s "O`�(�0n��yd�N�.��u�B"O��8dX�R��3&�_�L�1��"O�$��F?(����!\���y"ORл���*4?�0Q��
��0@"O$�ň�L��%��<@L��"O�#��9r���3���z,�,9�"O� ��O3C����P4q�܊�"O�u0F�YPo�h�$�J/ID>̙@"O�Ё��6L\�m ���]JbTF"Op�qf%I�N%�y���ׯ;����"O� P4C 0�x���C�
T�*O�uiA^��*��%.����'z�� �g,u0u��U9,�!�'@a�FH��2���CĮýS���J�'� őL@>2�n\3�闩^�X�Z�'Ť�Z���$,��D���Ya���
�'ԚỤG�'#���:�EG�|�0�X�'|TeɅ��S�r����� ���'��q ^3-KZi§�0�"p��'S
�JF��2\��0�A;l#�L��'r�uq�a3m=&��A�5�*u��'c�`�H��V!Q�&!V���'�Ԑ�ȏ�kS��SE`M��,x�'�$�knXn��=���V�����'u�\������Pd��R`V��'���Q���Y?���3i4�n���'���2�Ȯc5���#B�70�j@��'���"��*�sԮ�V��5a�'�QQd��&B�2e�2�U��\)�')����Ə�
�����J40U��'4A`'�O�XJ᱁��*��	�']�a8�&on�{�9��5��'��3�&B�,�t9�51��<��'�Z��ӿY}"��ըڻ!V���'`�ç�_`�������L		�'���Õe7�\x"tA��N*t�	�'&l3��Bʾĩ#�͡X
��t~64��?f����2#ӖQ����S�? Q15��L..�)���Ph�LA�"O�\��jʈr�f1 A�'�v0"O�%z�B�\Ģ���;Ю�zv"O�A�5m,1	�Q۠$1�vh��"O�1��cH3W}����DC�S�D�JG"OB�# �_$Xj���
�]q���"O���D��)_B�ǆ�Q:�<22"O��0g�l�B8�LA�/��W"O�%J:o���Ӳ�ݬJ6v�v"O�a�Tf�86OT�9�#��$�l�"O�1˶΋Hn�`5	]�Ao��C6"OB��Ν.Ē�b(؄p_�]�%"O:M[�-��@��%Y�UJ��%�"O�-S�(�:cX%(�D�5
RL%��"O�q�������g���0���p�"O�tcG)C�# 4��'C�?7��$�"Ojؘ���R��q����?	/z0c�"O�$(w��%�©���LS (��"OrYP �U�h؞!�7֞(�s""O�!�%"E5��\��M��)�N,"O�$��iI	&#CF�8��"O@$I��_=Q�a8��S��q3"O�		B��l��U!A�r�qj�"Oz�C!ՇP�e��	���p;�"Oh��a�821�i�GK�F��5"O�Ԫ����E�YcG�4�m�`"O��bF�{�)�槅.l����R"OP�G	�=f�*W�J�#Έ0�"O���F�3�ص��H�zP��"O���W'�&amhyx�KE�K����5"OZEB��JQᕈkZ��d"O:��ώdz����k:H"OhP�fbRWl��Y0ƍj�ʥ��"O���]���cu�I n�rٳU"Or)� )����2" J�Nu[�"O8����/O�`�I'b�W�Z�ӂ"O]bT�]3�5��X�U'���"O� �+1j��SA�,V��G"O���C�0d��3��Ƈ���"O��R��]�	˰̒RƂ��vl�"O:iб�&,Р��.J�bdr)1�"O ��a�K�4�@�,!2����oB��y�.��T�|5q���
�<C�%Ƴ�y���2���ЇF�T�W�W��yr�	�KPͰ��ЗrQ��h �y]�!��{v!Yb>�SPD��y"�ڲ ;8��nP{6؅�Vk�"�y�& �D�>�S�	ݠqf��V�S7�yҨ\.��8�%i+;2���v)R�yr�JdS�}!��Q� �6���y�Ą�F&�i�4����-Z`�
��y�)�%TP Y���:��T F>�y��z��Q�����8�y"M�j�Z�Wc��JQp��=�y�F�4���dKU��)"ݫ�yj�
�4�94�Ls��ዒ�V��yk�?v���c��H#?vR!Q�&G �y��!�4���Q%5�҉�W��y�,>:Ȍ�+�+	p��@���y��_6ΐ��OƑ,+m#!)Z��y��Z'd|��_Q{�ؒcJ!�yEV-B�*�b�΅R��Q�"��1�y���Vݬ�)��N P0p�q��4�y��R�n�v�ҋ�dR$��y
� b	� Ż3s�i�!}P��"O�X)1H�'z�=�r�ì:����"Or�bq����JT���B���A�"O�d*���h�D�K��(#b2�"O�h:ƈn<h!S�l@�9��I�7"O��!��P���pQ�+�,��"O|t �@�O�0������"O�YG�ˮq�v��"��k���Y�"Ox(Xn��Z��1(� ?}�0k�"O�,a�Y��H����G�D�=8"O��{"d�t����)C�(�w"O~����g��A{a�_><�J	c�"OXq i�+s�ܡ��'�5�H�W"O�Q�P!����b��)צ���"OVA��>PA��t%[�,�B�"O�z#��e�}q� ��@�"O������)Bh䍰���>�F�"OJ�;�Br3B-y�-��*�\i!D"Oz��tcq)���#��2�С��"OTi����x�u�4��Td`"OB��@(Ԋ� ,�%d��"Ozlq�8�򨣅�]"���"Of QEj��#~�(qT�V�;���j�"O��Ȁ-�?+
�	��%O�r��"O\�*&�ثn,�8�ď$g� d�@"Oi(���5&��0���-�3s"O�
�J[�Vr�	a�
>vMnmk@"Oz�"Q웟� �%��E�	�"O����ψ+�	�� �8���d"O��CqJԓ�|��kM z��d��"O�3%�X�15 ����Ps����B"O�=鐍�'UCrB�iaiNPPu"O�e�P	%&��	BON�RO��jD"O�ѻt�չd�2�Y�@�~H.�"O�Y{��	�����=_6�P2"O�Sb�	�āz��6ɔ1��"O�T�*�?|�ZE��)�R,��"O�4#�O�>�uj�*L7e�r�{"O�𠷎"17(C�
�%w���S"O��ЁбV�2���fO	3"��2"O��s��g�����K�5<�U"O�u0Q�	yg�B@k���E"O�ؐȉ�&�Ѝ��A*�vp�F"O�t���X F���Ib_+}ߞ���"O�̳uLC:d����#�ל0۱"O�5�!�AՁ�C�Ҩs�"O.$�OF�6 �@�˗����T"OX��k��?��0�#J���!�"O�}��]	u�Q҈S����2�"O��y���x���;e��+O�p@��"Of(r���6#�X��ƕ����P"OJ�cpfȷ*�l��Tf�2~F�i�"O�xxvd�5n��pr!E��"O\���$�M���K� p+6�"O$؁tN
/
��´Č!U'tթ�"O�]��
.A_����#�c��W"O�4� Ɍr阝�4��::��g!���{`��sdA����X�.O�:>!�̋g��X�c��*�^�(��O)!��4	��H�%��>i����j֑J$!򤛌j&�(�U��"��T�#w!򤘼i�(�/W�h���A�t!��/�^tx� �2O��¤O��%!�\`�,���n@�(9(�@�5z!�� ����
t�.(`�"Ţn���KF"O2�L�8�4���ݣR�h!��"O|Lb�1?2R;��W0'�v%r#"O�X��Nʊ�hE��呪f��iX�"O~��E�K(LZ�$�� 8K����"O\��F�&B��Ѫ�RM{�isB"OR��� ��5MRqK�L�`"YÀ"O�U
��ߨbq�e�*l.��s"O`p(�ٵd��EХon��f"Ol��#�4nO��ڰ�ϡ=7�5�""O:��"KB���i�[WO�M�a"O,�򓄎 �,mj6����L�0"O`)Q`�*r����F���X�"O��O%� 퉵Xl�"�"O�(#j_%	��B�!���J��"O( �ƪG�fY\0i�E�4iI��"Oެ��ރb
|(	�$�s7���"O:cG��(��,
g�e&U��"ODD��ƭP?8qQ��¼��$�y�B�<��ٰF�	�l���NД�y��ھ����l�v���0���y �l���e(J\	%�`��yB�п'�n�[�ƅ#[(�`�o��y���/��i㦘����;!��/�yb�K� �c�H2�v�� J���y���a����ȉT�𳇇0�y��Ay�z�3l��<���Ɗ\-�y"LD�x���c�I-Ѳ%����8�y"�ɶW:.`�sj� %g|9{�Ƒ�y�Ě Gh5[7��J��Dl��y�*��F3�#�)����bU.�y��S�\���	Cރ@�ꈙ����y�m@�3�ԱX��4.g�i�0cɅ�y��� r�Q��$5(.*�k�/�y�&��X?�Y�&)ݽ�p�Jd���y�@�*��,����~|���6$�y2@��L>��Y�(ѧ+9:䱴c���yB�ܢS���ba�Ί"WaуO��ya��W_}��W�d�F�1c�V��yR��;c#�!�`�C�E����@�,�y��Ͻe�,y��ø'c�p2��R&�y����έ� ��'N��r2�A��y��;W� P�OS�O�|,@��O��y�BIS�(� Ջ��Su�t��y�Ge|���K@�Q/�h�@j���y�Y/J�D�z�N�#a��d����=�y2Α������F�]�M�d��y��!�Oԓ 56@"�DN��y�ā
���F�Cmb���,��y��1LZ>��Rɍu���&lE��y�gT)�H�8���4CC�}��큍�yB��y��ѰV��>���2&K��y"��>X@Z�#P�˞�	��f̟�y���h��0�dňy��Hyv��yR-��P@��q"C��#�8�Y�B^��y�E��eK�u1,�0f����
��y"!��>�"�(���(�7���y2	Y� ���k��>0"����U��y"(՘=�|��B[,'��IE�S�y�+C�4����T�v*�DQ��yr⊑f�:D#�žp�2�P�+�y� R�z�����Z�l٦*ʢ�y��ԲB.\�����
Yg�8������y�I�%:�:a����V�E��y
� ���7�׈>vf����
6�,Bu"Op�R���3��9�1���5�Fy��"O���dX7h����MS%��1"O���c�"�\P;d�ۀV�Q P"Obͫ�芰/�Z��;>T�"O�U��$*,��((����)��|�"OfuYC.ܭ}7�pA'`[�R�D���"O���R@U��nd�M��p��S"O�UR����z���XW�
AX�!p"O �b�ټQ/T�è�>m�l��"O�T���!h*���h͔vf�Ei�"Oq���83�t�W�L00��"O����F��	�0I�E?�D�r"O�(����9��ҹUR��(V�!�X8��r��ҠUU�q�i '}�!�%5�Fҳ�	�/[L� �(Un�!�D�^��#�+mD �a4�@:.�!�Dج�F���ɜ8�5"��S��!��+	��5k���f*�qQ'��:�!���R7h�3����[���s&�K�!��~��	r�l!wB̙ń�B!�ċ�B,��GC0A	�ÄU-#!��](T��c���/jCah&F�A!��Hv��AE�q©��;
!��4E�D!�"h �;fA_�!�$<a��k�L6JZȤ����}�!��C&zD�� K3CH�M3���0�!�F8A��QS$�ă1`n��E�/ �!��&Nb�T����oJX)I�-Z�9�!�Ml1��8T�-���OZ#K!���6UVHy����"ai��<f!�Ǌ&B�ê��x��p�薕A!�ݱiv�8�eҊ-�tP�g�Z+5!�U,3����k��ǲ�12GQ$�!�	�$���B���6�<<�G^)_!�d
J+x1sGꜯ�j��-!N!�?B舱�łL��=��o��h4!��ݿ;G�k�Ľ.����u��D!��T�l��Č�k�
�o�H!�䛧Bm�Ɂ���p�a�	
�:`!�T[3�0`c=NYDt�TF=r!�d_i��F@O�RX�A1DC�}f!���5)X	�Ĝ�h�Ř�  J!�%w�>ف���-��=*ʃ�gX!�Ѐk0<UI��8�I��i˺3>!�M!pQCV"![)F���)�<W!�d	qZr��BA:ai�(;f	�!����Y�go�v����!
!��0]�M�cmҀa�n+���hp!�Q2���1�"v�	���/e�!�d����UZ��KQ�V�����!�!��C,+~m��N�>_�~iVl�!j�!���-��	"e$EN��Q��JN�c�!�V+e�(0IR�d��X�%��D�!�DF�	�"�c�cڏf�
dy�.�g�!�d�:uH�qbݸf�T���	��!��o�`�'`h�e&ӵ<u�ȓP��%�HP�r\x��u�'kl괇����pPR�f�T��L#:����ȓc� ��i��8��$�f	�@d�Ć�d;!0v��;OU(x[l��4�"P�ȓ ��0a�ܖƺ���ߙ����ȓ#kz����_�r`yXbE�\��kU�d F��4b��{2n؍p�����S�? Z���M]3���Ze�^�P2���"O�!�g��j��xG�7*�є"O�Aj�`]�l�X���͎"q~���c"O6(���̓zc��E��"G���yU"O���h��2C��d���aV6���"OF�FlˊIE�b�n�1���[�"O�л7�E��3ӮW!0��f"O��ŽM���b��IH~��rw"O��{�j�.)BF�/K|��"O�\�Sl�
 O�a�4�Љ4�A�b"O"3$��8�6�C�KR�y���"O��+�R<��8S��Z�J���&"OJ�BaL/5=�" ��a:�DZ�"OBp�w��|�V����\�΢���"O:�8�ffB�� @j��b$"OXI�&m�B�B������@8�V"O�qw�̄ml��pO�x�&PcS"O��@��Y�0�X)�B�GM ��v"O6�3C�Ȉ�6�� $�>V�EJ "OB����@L��b]$HE����"O����� ��݉�f��U9��##"O�����5�29	�F�G����7"O&�+��նFJuȡg�y��4�"O�%i&�K�D�nq)C�Q�r���B"O���W�E�y���	Q�z	 Qr�"O>� f,�,"6F]A��ܼ�Ѻ�"O�<fK��8��lX�B_͑�"O��S!�		�q��(�^d� �!"O��c��-�ґr����xM�"O(lqV	�o� ��%�E9A·"OJ-s���U�t@�Ƃ�,{Li��"O��KBl�<O��ʄ
Г2q� �"Oz� G�_N�aC���6�
�J�"O`UQ �\2�N�Qr
�q�5�b*O^�ca��� ���В.^�*
(��'>$}
C�L d��˂�u��a��'��%p7�\6"�����S�ii�k�'����3Ȑ?s��%�t!L`��u��'F�0z���"��j僂�S����'����ޣ3�
�I��$Gw
9#�'�݃5��%4T�Km��l�����'A�501� *D%2��R�`�
!��'��a���Ԗ���� D���x�'����!.��HQ�7�ry*�'h�9[�ɵ�|��ga�1F��3
�'�Rɉ��W5��
B� G�>t�	�'qh'�
�(P4�eL��F}"|��']t��É�z>.��C I%1{&x�':ƭ��
���\�SJ5��a��'���A��rkxy�Ҥ�'V(D��'�DA���(���3��i��]��'e�E��H�] �"
C�Z[~��'�4ܙ��_/y��B��}��u�
�'�R�pb+�0��=jT![(FI�I9	�'���
�U��,l�.�*6�Z�	�'>fi�G �	52�G������4D��Rgb�7
���{�pr�ܓRk2D����iR�!�D�uM	-�x��0D�8�RmW�l؅�s�
�
� ����.D�0�ᨋ`���B�I�D��-���1D����S(e�+UQ���B#*D���5�
$E��G�[G�y��o*D��pL
7[<��a�:EM@�'D�\�\f��$����.7�@=�0�#D�� �L�$���(g͎5e=��5"Oz���	Ŧ�$��V��O,�]��"O�,��W&����+�+~����"O���e"ݘV"������LGjU�1"O@�I l�� �,8�ǉ��M41Pt"O<\�e�*�,����8[6>i� "OR���hJ�/|���Ȗ+ű "Oց� Axf<�bGȕ5�T� �"O6L��.�<f�$UiB�Ȓ[�.<�"O�䪲��+�R��V��#�|i��'<8%��l�T,HLH�	�<θ0:
�'dЙ�ŔX<D���[�d��'�9أ�����i�*��~-��@	�'j�Mуm�/9>�ܱQ� A�`-��'����`��w.\ъ�@�6*ڨ��'�&qC��"l��9�J��.�i�'Y(���#X�"3�]:[����'���ж(��{J��b�Pg��Q�'ܼ5�ũ-9=*)�C,N�
I��'�(�����Hjl�5��&^���'
0��ĮVa:B�3�ϙ�(��L1�'=P,�4���g	�u��l�j�p��	�'ӎ�86�W[�����"J��k	�'.��MȆ9�셣�/�04PQ	�'�4��������H9��
�y�	J�j��(jӊ��4 g��y�V�H�Dȋ�����l����yb��3M*� !�-D�����j�(�y�싧d�F�y e�^z�Pc��y�^"?#�=�U#� )��2�+���y��
;3��U�1��=�fH������y2b�Q�"�e�����m��`�2�y��S@^ѹ�!�0 -V,��D��y��NP��_H|X0��Y�԰@�'��mkFOLG�~Yr�-�J7J�'yE���\��9ST*��W�I�	�'�L@��(�E.�`̾}Ux���'�
E���.��x��mڶp��4C�'"�4��v&T��G�3J�x��'�\��Bz�f��7�5%��k�'�����
2�Pڴ�P�"TS�'�
��2)�TF���ǁ+5�ԄK�'/\l��J�`���#�c[�2�
=X�'EN��Uo
�e��%�v!�2�P�'sZ���O$0��Q��X�'=8��4��A`�5��O����2�'��c�nӊy��@-�4P��Y+�'�������{놵�G�	�O)�x��'�L��W���e�R�1���0E;F���'_|�Y� �4Ex��g�߮6����	�'���fb��0g�`6_�*�B�"	�'�q�3i�: :��p�e�&����'���5Έ�<2�a֪G>"rv]Z�'��`��f�7�B��to�:PrX�3�'��L��@�t�|aN�&Q��I�'���7iCa6�����O�"9��'s^��E�ɹT�J9�@��8)����'ָ��O9Zi�,�`k�}*���'+b��-��d��f�L�tH,|S�'}��P��g*�ej�l�0P��'ٶT��d�s���b�ʓ3�N���'��h��L>�d����
2�p��'y��8V��db؄��.  $vnŲ�'.9AlB�e�H���� @��� �����2
LA�so��n����"O(���@��q�7!-2�>	�a"O��@Dg(I�����_BΕCa"Oҵ�f��~�x��b��!6��94"O���L�75�i�щ�7H��E"O�eb4�	+����>|��H#"OVH���3$�\�ӑF�c�� "O�,�Gc��Ak�-��]�_���s�"O6�ڱ�|{�%���"O@I��H��K鄘��C�13�x5�"Oz�0���^��q�4S�{<$9Q"O��B��V�-�j]�w&̼.N�%ٷ"O��H�/�v��$��26��"O����ʙ��T����E5�̩�"OnŀìN%bϢ,؇�E&.�x  "OP��C�Y���r�Ȟkw.�qu"O�C]�6�0)�7uR��s@"Or8t�K(P�B��a�T�T���"O�@�RB�(0�Iݴ���"OL�,�#�XS1M_�N��&"O����ץFT��pe�Q�
y��"O���g�����lZ�A���ؒ�"Ot(��
�'��4q���_�(3�"O���@etʐX�!Ϝ$T69�"O���V���FZ�T�A!�B)n`[�"Of�a��^�G�8�
֯y0��@�"O$t�Ѓ1��	S
/I{rA@�"O��c�ӥ6����
��Ctt)��"O�|��j�UL����ʌ(l�qy"O�(�)��)�r�N˫-� 0�"O֠(��NB騬��͇#;�HI�"O�ʧ瞺4�V�`gǯ)/��w"O�+5��D�@�w#��Hh�I�"O$ѐ�+M
b��0����+
|��"O L10	��b��&&�I�(�"O�  唐1��,�f�
�!	\hS"O�}b�jV/by�W$�`��2�"O�0`5�N���D�S�̿A�r��"O�YC1��O'�kS]"	<���"Ohd�l�<vt��J��̩A~�"�"O^%"�k_3(F��;�ABD t��"O��x!M)p�D�gA�F�$})G"O@���jB5o`��p�-ck�1�u"O>�J�^*[U6})�c�0Qa�1�$"OY@�ެG6�pb�YJ��Y��"O�U����n�������A��"O,�
'�U�k8�����%	w>�H"OX��":efB �vƔ�Z����"O`�! |��"�
[8`�F��"O*(
���â���0�vTbR"ONI0�a�#�@E� ɒ�v��"O���#V�x��x`��;�����"O��KDj�9��kMK�1�����"OVi� lےe��@ mP�d�Ak�"O,��h�Rxᐲ�
 X-C�"OD���>U�E*S�ؽ�>�ٳ"O,-)��%=�����������"OT�z�a�(;:Mc�*̣x����6"O��AT�]/�$�S�^�@�p3�"O������~e���1����f"O�H���0��@�M�)XJ��"Or���C� [2|�QM�4]:���"O�MBec�<��	�Pmɼz0d�w"O�ذ�F���J'-�6z��1�"O� ���%F_#��1��$b简I�"O�!H��:��I�c∬�F=�6"O�U`6B�r|�K� �,G�6�("O(��(�4[M��zQ�A�+��̚V"O��qR-�(u'�!��-�2]`=��"O��`Q��#�H|꣌G�/�h�j3"O0��tb�i�P���*7 x@��a"O�8�f�!tȢ��E/ڥ{k֤��"OFy���Ǽm ��+�kD�3���e"Ob��qIւ|��AX�䐫Oԅ@"O� �	R�h�ۓi�'eﮅ�"O�h*f��C��2�<I��"O6�y�]D�@(Q�%�.�\t!E"O.���ļ�Rٙ�D\"�a"OLBÍޕ9C��#
I�y��"OR�rLY/,骘xDǠ`��0"O�P@F)�S��m�2J]�L���'"O~���ψ�`=�P�h�,w!A"O�t&�N>|hÓ��Xx>��6"OPC��FPVD`pF�X�I��"O����� s�rA1ǟZ���!�"O��2`7=f��х��z�e�V"O|�)�JG�}�HB�اym�ݪ"Oz0��kq$dXj�#R2=�"OhɃ&
=Wn��#(�)�f�˧"Oh�R�#���J���&6i��W"O�us5+֊D��P�Fºh^ti¥"O��;��٨@E+F��j����"O�L�SE�Q�hpB�K:0d�:C"O~�0vA�:m���j���Q�A�a"Ol�k�ɼ/V���*E�Gh�9)�"O�$�DA�=Al!)�B�!^i��: "O��KG)Ď>r��j��ڋTa���"O��F�3Xf�QcA��42���Ie"OΌ���il�4�K{�8�Zf"OH�h6^�hy1)���V!�"O� �A�0U��@;"��)iцYKv"O�����t *�Dh>YXp��"O�E�Bg�*��I��ǀ"b=��r�"Oԕ{�ꑒ�Fѓ���2j��$��"O,I� )��Q�*��Co��`"O�d��cjaT,M�I�NU�4��2!�DU�|hl�(4M�6�0�5�ԸT�!�C�`F��u)�=jk�x0��^�D�!�$W�E���*PO�c{����GB!��otn��S�y��@���!��: :CIL7rp���Tq!���� E�dl��9R�̾An!�D5�$��u�ެHTdq�7�O�B	!���6n�B������T�۳;N!��C�lc��3�5XxV ��*EQ!�䅯dS �	�ۘs��4
�S�!�䅷B٪1�hЌ��@p/ �!�$��M��M���]ͬP�e�J�9�!�ą�*��٣��� '�6�8�p�!��*HT I�1D�cp X���r�'e�IQ�ʙ4�ٕ.�ʴ�'T�@ 6͞�h�Z�f
|�i��'}h��S�_�(��iV,?z��	�'i�=�oU�|�&���׌	bC�'���B�N@�g�f��'�$<�G��e<"�j��ɷz�:��'�AJ'�ǁg�r`f'E�n=Ꙛ
�'A�\`�R����s��3~�h��	��� �T���Ģ���u�B8J��-b"O��ă�Wr^u["Y�Ǹ��w"O���)��6N���,޳��%"OX1��Sٳ�T�H^��"O�E����=���C�y߾M�#"OtIC�ֽ+�*�3�KO�='l!S�"O.�+��� �0��:@�L��"O�P��I�n�>��C��98C-!V"O�8T��e�|��䉔�X2�E��"O؁�K$�])�i�+s!��""O>��v�Z��롨� N5Y�"Oڭ��e�~c���!nJ�*c"O�A��->ڒ0��mA9PRmPD"O@%�f#H?|�f���E�I�t� "O�Ik�e��lP���Ce�h�1F"Ob�����(G\�`���
�y"( pU�-6LY�S�X� ��ɱ�yr
�T$ g%û?(d�����yb
�(b�ySDgJ�2�����(���yB�X%G`��X4V��ucƀ-�y��3B�%��'N�zMN0S%�yG�I2E;GFH�=(�@CGT��yBl�,�҂V?f������y2gM�
���懐0�R�C�G��yoεX��<P�g��*w�a�K��y�ڷ�Y��%,m3R�HM� �p?!�O
ij��G:rri6̂v0���"OFQ9�
l𾕀�k�.�U�"O�=��	�_�)+alH�X �"O��P&���ɉR��9-�,=�#"OP	3�'C@�����(C1����"O�(�$k�"�U�CiU&u���'��Ip��d��اn	�>��V�^�?$�B�I/M&����b�JrXC޿E�DB�!n~cp掽	_DI�@*b>B�I/1�|Us� �<A��F�S�,�����	?i�N֬�
J#0aVS�)��nڶtK�ݳ�H�+��u:�mS���C�ɮd��w�H�93\�aqm�7/8�O��
t�'3qOz�R�D)�|=Z�ҥ;��� "OBP��H�U��$˦Bӻg��и�i>�C�I,P���Fnچ��(2C�I�j�ܸ��Ϻ-���iÇ��f;�=	çsG���'�ܸX��@d��D����hO�>�Bg��& l�ݛ�Q�h'H��W�O��=A������T}�� ΁*Y���tA��\"�'f� ��ɝE�����Avb݋U�L�j(��$���:wOƢ%����U���KT��0>��)}"CQ�@I�C���Z�D��m��C䉞i�6�8�!�����	�~�8a#!Q>-(`m�$_D�)�o��"�0�'D� P��K8�њB��/��|����O~c�pn�H���dϭR��ti%�X�T����N�'Q�8*E�'�>Y Gˬ@ht��-��t/(�P�;D� �dH�V��*�A kr� ���O��2�	e�O���#�*5��Zg�FG��1��'�U�"�v�H󗄕�;IJ�-O�=E��.u�谺�e�uz(���yBC�	���S�ϓW<�����I��ybC�,����Ն�gT ��A��~"�<�S�O��)��� r�bq��A�/U�8��'� �B���̮DZP�T�T��8xK<��&2���L�*,`�9�)��J�d���	����	�c;i�b�+-�ai'O��gi�64�(O��)� �Ms�\2q8�i��Ck�Ă�'j�@?9@���H�(�"��.4����zy�'�6��6F۴~�%�@)Q5J]`��dR쓯�)�}3��P7c��d�i��9i�!��>iW0����B�5���7��7Z��'{a|�A��U�x�!�/��|pه�0>�I>�#��Y׾�B7/[�r1��ْH�E�<�V�к")�m���� 
Z���2���' �I_�Os�1s7(' Y�cs�
>�"�3�'��p��
GB��jw7����N�D{��dm��ZW��r�Y sԬ�(��ب�y�B�)G ��+�E0hj�i����'�����D?�$��q^t5"��-dF* Q!�CX�d�>��Z�+��x����H����0Yi2B�	!|D�%৩AE	��L�3X�VC䉪W��3����d���@h�c�BC��7UXY�BN\<`�8ck��O�|"?Y����NA���Ҟ"<��$��X�$ @"OZ}zAN�wnl ��$#ö��0"O*�r�!�)��ց�"�~�I�"OB@7����0�',0�ђ"O(`@����5���ە/�%p��&"O~�I�n�F����-�
Zj��񓮻<A�O��)Fx"��q�hqc���t�B�'!J,�p=ѮO��d�O,5a���3z&M�#
�Bt*(�"Ot1��G��:�ĠS`4Rt ��d4�-�'��)��>�X��$Z�3L u�ȓ9� �"�o�xAbU�z�%��D{����]r�"���G�4($��ʖ�y��	C5]�Ƥ�j^ⱂrb���'��z�F!U��R�Ӌi��
�삻�y�F�k���F�� ^�������y�bŝ�la��ŏ!K
�cDF����#�O4��p�أ8��Y��
��4��"OF\���>�q��Վ ۞t��"O$Y�e� �#x�!�$�sa�ekg"O҄8Qh��-���&e�, Q�d��&Z�'<�x�� ��Ԝ��#+����W�p=�}��\`N>!�&ut=�Хȵ��?ٛ'9��{f�0l=�B O�#,���p�'yB���U�1ЄF�96���'w�8��I����A�<l���'�x����^���	�:+��S�'.�ElK>r�*�Q@_9v�pa��'��p  ��7x�p�b�l��+�' ����3D��eSc�
�a]A��'1�c �}Ÿ�A��K(W����'X��P��[����	�/>�]�	�'���
�&��� �o�)e[�h �'���X��POw~�1U�[�b�r,��)��<A7 �	iH� ����{�, ;���'��xB�];F��;�"�&w_Ƹ�b�&�yB�'r �fL���[v*�"ؾ)��'��L�Q(��J��L"�N�?1;U�D�O?�	�<�!����)�L����E$u/@��D1}2��E�Y �*[�#<:M:�#:�<C�	�\8���M��6��Vlv.˓�����+0h�F�����XjB�g���GV*�Hz ��o�T6�"�S��M3�/��B�xQc�S�]k�RɇQ�<���90n*u/x���GB�K
�l�ȓ�v�ZUOL�*lF���Y=�����	H�'R�QC���9`� XR�\-% �
�'+ ��	O� W��1B�/'&fMh�OD�=E�� f�Qifd��g6��Y6"O�ً��N�3�4{���$Μ�#�"OfE�fh��� �WK�$4˘a�'��ē���X�V��M����q�7f�!�����a���ol�ꗣ�/+����d'�I��A
~�d}0l�y�	֔DV��)�A)t(�(x %��y�E]�	�b0���I�n�L$@M����$*�O*a�G��?�ͪ��S�\�@W�ę�s��)�%��eSPU �0T��ȓp1���S�d�Z�c��_8����a�\I�0oF3)�  �읻)Z�p�ȓ���6���FPu�ĂN�C����ȓ{nX��`�V��v�s��N6�|��T���Z�*
)� P�fI�<=\(�ȓ-�f�����n��$��RI�ȓa�:���@ڹG�V5��8:�n)��C�Ċ4邜i���ԬJKډ�ȓ��b֨"!�Mpa��w�t�ȓ)P�����GW��R�p~��?��T�8�����:�I:�G�<LZ�1rtlP5L�&8��U%�"<D�����*=���j0�MM���I.D���'㊬&���Q��CS�88�0D����Z`z)�a/H(��1�/D���A
��S� p��U	x��7D��0���u�~k�v�~��"5D�d��̖�G��x�3%\�fyQ-1D�8C�*F�
��O�n8��n.D��"�+A''�ꡂ(��h(T�� .D�,0��ۘf.p��U��7b�@H� �/D��xt
�4M�����n~�¤��:D�0�d�D!=s)�6Rځ	Ch�Z�<	t�W6M:�����'��d�_b�<a�ߘAr�!��JQp��H	D.Jg�<Q�,��89��B��
�)LLU �H�{�<iBBF��^#�Ζ�g�m���N�<�A��38�R��#�<�5�_K�<��\� p��"P�-@�	�C�<Y�cF&y6��� �7M����@�
~�<��?>�&�ʦ���9���+Re�<Y�ޢI�n-JG�35H�xrB�J�<�1C�`w��2�����h�#DF�<1��+A(N԰�n�H��J�<9�G�1b�ՂA��F��QDEl�<iaGѳ6��Q�ǐ�"�Q҉�k�<ya�)Y�*D�`�_�%�B b�<Y!a�(���	"+L���0G�s�<�G�"ː���T�frB@��q�<y%�)����"a~��@QW�p�<!��/*����Dh�q  _�nC䉎i������(�ʝKEп|��C�	�}a��	E�+@���.R(��B䉅$�t��˂M��y
�'<f��B��9C��y�� �r<��(g�BH��B�+0�:����H;X�+4-�N��B�ɔ��T�S��-�}��ɵP�PB�	eq�p ��"b�$q �)��Y�HB� �la
'N2��0�Ęv=�b��HV�q2��x�(�%w=�-�ԣ.�;�v}�K�~��KeIǴ��C��.c4��HTGK8I���@Ő�.B�I3EEr��AO'p@��ؑ���>B�	�N٬d��wѰ1{qj�x�B�	.2���D���n)�W�_	�4C�)� ȡ�qCM����Fh�R��ݠb"O�A���I_8l�U�U sz���"O���& ��$FB�0a�|� "O�$(�Z�⪌Z����P&�pw"O���CZ9�.�{䅞�B��Q�!�$	��`�Y�&Z~l�`�4)��!�_.,�TÄ�_�lV|h.�"U�!��X�,�bl�)@H> �q�V�G�!��<X�`+�AJ�<���C��!�����Da��̲H7��X���3�!��?Y��݊U)͂���qӮO*�!�dݛ]4�l�@K��&݈(@!�d��>P�LX�K�����FmE!򄍖>��r"^�M�$�IO�^F!��E��i�' ��p�^u�t �6$!򄂊iz��@��v���ࣅ֜�!��T�7 ���&��m���b���;�!��M&5��1xf�h40<�Eh$�!�d>0�����Y�a�ɉl�!��~�&`htEǓi���'� �!�U�Ez�Śq!�Y��q*��
�(!��SXh��6S�4��oB�8!��>D�� ��iG�g�BXz��
Aj!���I@$i�$d)*r0��B�P7mm!�$�=e�( "퀟m�I�5�Oy!��W��a@���?9�v����?X!�H���]a��Z�d� �M�+X!�$7s���ւ24�|2,�T_!�G1�R�ӥ+��|</4!��J�g[����%�5�ذ)�o�!�'��Ĳ��'�����^J�!��3����쏥r�h�1k�/F�!�U�^@1j���W�R�Ǎ�46!�$��
�p�kN���M;���:!!�D������Q��bU�d+��$!��[䨙 ,F%A��IQ���&&!�VRL�� 
�h���ď�)hhA�ē��%���+)��r�"O����9TW�=�y�!E�d�%(g��fڌ���yb�&f��p�iS�^����G��|*8��5K7�)�S(K<�� ���sꞵ��n��aЪ���
�nq*�n�+��)�'4����`P�-ľ$�`���K ح�a��0O��ʉ�L>t拋6' HzV,�>����Sq} �2pj.pA���<]�����rJ�9�/
:%���QE �{B���!;LO���B`�"�t\���X|�<9� ��)���[aW�;�QD~2F	 �RY!M>�Cׁ����!K̐Qu�L�'%��PV�������+�����ϟu�f���0�O�� �!�b/
b��i�H���P!<��Ё�ѶZd�Ԩ�K
9(!�s�ފ����Or@��
�?�BQ�ҏS�5����Ǖ��8�O&x9r�1�3}�P�R�蒀'9'h�@���~��W9��	9SEJ�ayb@��p��fƔ�%`0
s�I�3`z�gAkaF�D~"#��fC��A�@
mLܡ�#��^l�ya�	��o�$M���'��Ы2�ҭZ��E���(c�ܙZN �BJ�)�H�Gy��<���x��]�XL��$�P+@Q��YׇZ�I#�����a{  �����pH�IǄx7��j��(�^�/I�%�xP��J�%��������iȁ.Ȃ��`�R()��W��<j��0�2�XY�$L6|�>�b|�h��敤Pp!P�%٠Q�'� ��"Kz�(��ɥ} . t��R	@I�A
��s�P⧀�0B�ؕ��'�U��ǒ?NX�&ǵt�j�V\@�}���'\):�ɯ#�4D�<X��a���
G�١��đ��h���1��!���`ד
N´�=�k�&bR�����ݬI�v1w�ED��i� �%x!�d�u�$ %g�1er��
g�Q4n�!�$���tXsj�J�.��3F�2F�!�� �hj �5!B��Y��-ʸ]��"O^
�dY�	pF����3K��uy�"OV��WL�d>�s�J�52���"O�U1%
�������p�zx��"OV3�'	-��;Ո'N�A�4"OtᨴHV��ڄ��N3#��,��"O´��e�����fH,����&"O�5p���0z�$I�a`���'`>x0����VO� ��	�-������',�@���/C����EJ�0����:0Y6�3���:	}�$@#��kF�Po�^�<�F.�X�j-I�	Kx32���CT�M����q�r�vK)�'��Lɓ�2k\� G�	y��p�'Ծ,r!��S�	�J��bCϻnFp���	�W�T��`�U�(<���f ���z��<9�$*���:�燎*=6��f�e�	(:8��F�'=�ؑ�i &0;��6S�3�C˜J�n0�P���@u����(x>	9��, 5ʸ{Љ\>7�����`��qO��q��A�� Ӹybr��C'��'�����֕�5�ڬ}�@M9!��a�'S,0���q̓ZUj0�t� :-���HB9BY~!;���K����by����U�zЄ��-��?��ଡ଼�_�����M�X�H��Ī<����589fO��$m<l~t�JtJH��~bl�T�,�x�!F�Y��U���w�b%ՉÎRn4��'	�@���h�A��]�U9$��	�)�<QWa�,W��B �@�F7qX(�T�{"�A������<d����Ų[�|p�5��=wX$�3��/,+\0��	G�Y�ax�B�0��� b�,3�~����?6zm9v*�$�:�A��H�c`���H�r dG��#U�Ȅ!M }cr�UϤ���@T-fd����M@������7��i$ 4���B��ēS��:�hY'@^E@��Z*24R��	�2��u*t��5��O��`"�*U�,�l�	Ū?��я�DөT��� �%I!F�a�H>�*D�ϒzkX��a�T<?Lq�3�6E��0���O��1@�B⮓�qO�E �@�$A��YcOF
l3&�O$�q�h� �3]�.J�O2p!�h��R���G$�4P�M���,�r���:yFa}�G���nT[�i��f%(:�QYuR��A(���dKB#�����jPK��J�a*0Bq!����$�V�;Jx���̐2j���v$Nf����)R�_��YtF]6jB�=i�0d��%�se\Ci�U������ls�)�39R�1�$����Ec8��cGΕ{P��2FL��/ >Q��"6D��\X���_�Ҍ)��K麋P�61���P���� �"
��h�OV��Gl��C5��qO�D�/�<u��d�n�P����O�Sר">��D�V�L�2j2��'E>��1��՛r/Sc���5.A<?��T1���*�<y�n��ps��M�S=��2W�Ó<�\�����2C��s�c/s�6(�s�Y�t���R9��j�.��<�J�6I����-D^S��wg��[ dC���V1�w�}PDEcR�N�4Ŵi���(�T���%�6#|�hS̛�hٰb�<�!�lX(�Ĩ�1�̧��J�-Ч)	��A��Pb4u��DԸj�,mq��@�S`����$��=J%��$rQЉ�2�٪B2ĕXJ��;3%S0R�q��'O��	F�+�ٓ&ᛯi~`��O�Ua�h�
�l�s�%X���I��i����ц1+]�x�3�ٌ��J�K�g�
�Y��H�q=������V �5�5�̅s6��I,?
�Xe`�R��Az�v�a�`%?!������< ����� 0�'XN���0���;���'� [$|�vH^�jLءh�n	!_zx��E�n��y���]J���OV<�MS�a���Џخ-1j�K	�o��e�|�pa�Aý�  k�,lf����ڕcTfЪ�	!��'Ub����)�3�,W�� d"U�]�b����W #�'�f�"�K/9BB�E�����4���D�u#"P�.��|��-JP���/�H��	v��3Ph.nD"ɡ�G�
��p����z��@�n��9٤G�>���+I��m�)Ʈ�~���"�f�!�dG�r�X���-�>N����!�+��|�Fa���W�T	L��釥|ta�A�7�"�(�����Py���*z�PǍW�9UTu���H� I�J���2CQ��q��'��2 uh�"�/0����'�P��@�� �|�#�ɘ�@�x6<@Q/IG��xX�m���- ϟk�~��TB*OL06(>z�!��O�}�#D�wltm��ML�=n� �"O�����/BzN�:%�$7�4}���>�U�ʁJi�q�p+�:	�#�����#5�}
D�2"O� ��k̰�0��ȕa�8 É���a�, P��x��$BN4Y��߇HR�EQD����x�	�*q�"�(rpL��nT,F�;��Rg8��s�n�G�? n�R�ݻ3J� ���(=�$�d"O�P�C�!	�p�3G$ź	��*��	��U���I��Y5˂�V�(Yx�k�-�;B"@�u��qܓ�h��d�CL����G"F��B&
�h�I%|4,8	����t���Z��UYrH��{}���ߴk	@q#;�p>�*�	v�����IC�A����FAz��Qk�����MS���y�ֳ�Bp��]1^�2dy�ט�?�-�/c"�Is 8�8hKC�ʁD�U�E�9�I�F� }���2?���B�f�
 Hs��'Q�т7�Ft)�  ���2O(� �L�%6�c�-���K3C�G��',x!F�,OE���i ���F3�.B�W�� o��S�OخM��ׄj�ty���Wl�˄��m�dq�
��0>q0�=M!HL�" ����s)]�� (q�D"dm�@bd7O�� �Ü%)�̸��!��!o��"O�0�6 R��z�!�=DZ�4�R�d#._�Qy�EA�����p��N�j �1�??0�X��"O�)3"�P,��]  l Z���1+\� � ��B�>q�6�gy����2��!��vgz��.ܗ�yr�W�k��aA�(�+iJ$�Q�<�M�T-W�.Mp�e�y���1qn�A�ff�
Jƈ��I�od���4P�ha�%Se��C���{�j�!q*D��dJ[�X��,��J���Q�3,D���הk� ����X�@�4�!(*D��:�$�lT�Ea#L�y��o5D�d��
��+�^I�Ѝ�	j��9D�� g9S�x(��F�,2>@�@�7D�`�/n*fKI�lŨec@8D�����6)zt(��MG�R�ؼq��7D� *R�-}����CȂ v�����3D�(��ٗ�D㆞?)란�#f*D���m��b�2�`\hYl��f�&D�Hː	�;���g$*F�Vl8D���vBݿQ�怑BJ/c,t\�4D��d��mQX���T�n�0��B�3D�`҅�P(�h�u
R5gB|%��,D��Cl��4Vevi�<^����,D���/�qHb�G7b�e�%�(D��[�nǬ)�8ej��G���S�-D�����T�ތ� K¢_��P��'D��X�c�1*�^��eA�8�N��	$D�l"BɤQ~�8���\�	b�j�a#D� A�h��氛c�1(����o!D���'&T�l�\)s��ZH�މR�$1D���ȠLJE��D��JU;��/D��s��dа��K��'6�!E�+D�0���G!pEj��Q�M�f�����&D��JV�3�"���كj�^��h.D�EC\�[��P�R��(�4�pV�,D���d��Gz�p��֜�����+D��B�B�}Ivʖ�R�5��4��-D����%81W>�*�aZ�D>|p���+D�H�@Eu��U�"Lk��L��C'D����.�Rܞ�B�c
G1�i�h'D��r��6{E2��.Q�4��1D���G
��lG,���ǯF����i/D��:���a��Jb�FR��`��A0D�T���&h~��R�ǓY�ҵU�0D����Oh%B�b���Vb!���=D�T�a�^�L���S!�5eaX�O4D�\�v�Z�T�1R���B"٣�'D�T[��Ι�C���Aހi#D�,Z�lSOB������(]���0�%D� �ӌ͎1.�Tʶ�/:�ex� 'D��9���a��=# eߢf*�	���(D�� ֭�@ ŤQp��{dMW-M��Y��"OheK�`�4S�2�FS-p<'"O�����כM).A�G%\� �tK�"O�Y��KɯUZ��b�JZ�~`�W"O<ihR(�:'Yд����G��ڵ"O�|*6�[rP�S��2Ԣ�j$"O�s�kP8��ȗ7B�LhkP"OJ,��P�.�@�уfX�2��۷"O�)��F)�6���k	\�����"O YUcذ ez��0�7'��|A%"OB���۷�2C�"?�45A"O <z�"�*7Y��+�{��H��"O��@��H�},�i�@�F7B,0�"OJLS�C�
���D*��CNJ]�D"On� ����l.��d
���!H&"Oh�2%�ʬW�x�j��jâuq�"O�H�'�әNr��'�-S�>X�"O��sǃ�.��z4��v��yR"O6Ͳ�A�D�A�� -?�Ν "O�9��-A�EeDI��"O 0����(,����E *�h��w"O�hE�D��P��L)(`���"Ol�ـ�ʆJ���@�h=�Dx�"O<x����47@�,4<��ؗ"O�]��,U1 �fI#��Zp���"O�����\�Y����/�T�"O��$g	��"a��U�P�D"O����T#Q�j�"��P�3DL�h�"Oޘ��)��pM���6���Ze"O�!2A�W���r�ܨOl�KP"OD�����:������`,�p"O��bs	ؗ7l���ѭM�OnB�j�"Oz��B(em~�	vJ0b�"O�U(DM9hʎ����34l�"Orzg�N�lT`Yꂢܲ?庑��"O���	�)�0R�ܪ �ք �"O��3� �9@�k3m�&��"O޼�с�c�v/�%@�6��e"O�,@��X��J�pQ/<�$!"Or�������*��U�a���"OX3��C�a���!�/w�:`Y�"O��2	ʊZ�`!D�	F�v��"O���CD�K��īǧS�Li�"O�Y�F��l�2��2�z�S�"O���6%�9��0�C�1y, 
\�&e��8�� ��|��i
8)����j��c�&TɡNV`�^B�'Ԕ���CM
Fn8�s��+nH�hZ$Zs`��	�\���)D*��Q�� �Qp���~��|R��mY��4�Q"���2e�c�H�P� ~�q2O�3�̋�l�Ԉ2"��a���)��ɜ0��4cQ�
�h�܀�~�V�]�f�<�7C�wx�	��Q\���-Q$;��5�����,،�(=3�gJIf9X�K��
ƚ�����~�)��`	NN�*�+eƮ�3�'J���L>!��*�gy�+�,/^]2���@R�z��a����P���x�,$�Z��DDPД�ӕ�J]�@���w@`8�-ؼX�����DB�z� �ÂB�nB�P�C�W;s%t��S)�>��p�-,OL<�ԿKU�I���I/F�t�0Cl̘rn�Ô�Mv>�<�!'C-C�`�`ì̙��O��93� ��\����30�l�y� ��4;�@j��r�O����QA�Wh��ccP�:��y1N�:!H`V�84�S��?!w�GB�!��Y��Li�(W�w�f�)T�;}�j�,���I�7=*���� N��T� CF?ki�_e��0���G;[����rnݯnM�	:�_�c�~�㵨H�)������.���/E+jԓ
�Т蠱嚉l��j�iTz��"-��5vh�ɥ���3��M�ZkC�	t�\4	��� Zm(i�$P���"��e�HE����`�&�!�*#�'3��MXs.�C�8�۠���ԆȓM{�8�k�	vmPa{�V,[,朆ȓ8��̈��@��	 B*Ȇʓ{4�$:R��D!��
�cx�C䉩_�*T;m�rĚ8;�	ߧN�dC�I�4	������:/��*���-ˊB�	��0�Z��]�[݆�sa"@�hB�I'~ePM ��]>�I�PO��{NVB��n�$�I���R���B�����C�	4�f�SuZ�Uj:Y{�&ҘbDB�:���A�)�hio� 9����A,��B��=����	uK,D�(-�0��r؞`���]�4z��iF�A�N����?�29�5H�0 ���'��ģ0���ajV�5l�E�h=j�{���#J�)��ބ� 	G��$R:M�򼫶­\�b�"��/�yBH/D8��C��cr�6[���#�5�dl��'5��F�,O
�`�%��+L�Y*a�)9��Ñ"O �PD�1���i�3|(��u�;B @y�N�@=(,��'�ḷQÔ�4�<j"��"bX�	�+�� UHD��hp�aφ�}ۖ��\_�} ׷�.�Z	�'j0p� eT��ܹ"&BN�j)(�{ ��$ CJ-�ЌD����=u��yBRJ\Q����%ON'�yn��^��4��D>z�5�WI>f��E��!LAx�'���S��d�S/�m/��[b�P�M�<���-4���5/�:_��-E���oC�)�!Z�>���IR5�f��Z�������H�@�2Fʍ>��L��5<OD�Ɗ;��\�����8�Z�ztoG���Z1�A�Dͼ��Q�7D����bI3,�$�[��q����M7��]�{���T��-|.�<ˊ��7;�4D�%��t�a��L�!�b�l��v��*7�,jAb��[�v�p�iy�Ą����?�'GbM"��Vx�h�d��rUzY��'��\3�n�x4 �F�gG�XPUC4V�aЁ.�CX��R��-m9�{�-�#dfJd��M#<O�K`m!anFt�O
�ӏn`�I �8wm¤"O�0k!n���0�Ǘ��b�`3�|�ם�l�Pc�Ns�O`18��٨w�W��XS0CCL�<Y5��[0}�a�-2����o�W��H��G	������5p�ەa
=ľ%2��P E|���8��"���/�P�aSȃ����"�)F�A,��JA(5�OB�K�g�2f��-�b�J�3�z8p��'Ȑ��.7�$�'�P!� �t͎�ђƅ�f�Dk�' ��'-��&,�i�m�+�N9�O�P�bڕ!Z�ZR�O6��9G�ԥ�`�͏.��3�'|�	Paʆ)|��
�w�N��c����I����p���|�ێX�@����!�<%P�NC��Px�͇-6�Mh�.c)�I���<��H0��Їc�
���(Uv����!ˏ���)\5C;l��dC�/7ZL�w����
�W����P�j <	.�z�y	�'��%aX�F�h0��Kׇd�<IH��p&oW/��	h��O�c�/J6l'>T�W�ۘJ�n4I�'����$��a8( �A�_�Z��5��HKJ�	�[��!���L<I�V��p��	�"a�%�3�m(<�@�����`�W�j]|��uJ-%8	)p
t~���X�d �)��Bw�E2th�A�x�T�|��yvIPa~򁀝JLh���++[�A�#����y$?E(ȩ�2*�@ޜy� ��ɰl2��Y3�?�a�Di]
^e��;��̾nȰ"c+!�y��Έ~�|�SN^?13Uí�G���O� �`�Z�-3q��';8�{�b�����;X,�pH�'�Ρbs�C<� �����#Y劵�53"�c�Py����)���:.2骉+���x���Ek���F.�k~Bc[�Xr���ܑ[��Y;4�\��y�ޱJߔ}���D�WO"T�s�S��ɉ%��X��'P��a�� �0�$i nQ<!ņ��R�SD"O�
ъT�^��P��e	+a�0����!��a�8��Q��x��f������Ǚ"��2@���x���
Q���bĊ�q�"A8���$?�� %��|؟�2�(�i\0\�Gc�2	o�9p9D�`��L�Uxxl��%K
8����0D���Ā�JL����mJ4T����"ѪLi��{�� RD��)�`��SG����,D�|�h3��`�"i���
a�� 0��x ����(�:A�2�B�liL�d�&T��z�d�
���I��<�P�ϱt ��C�B�Om�Ja�N�<�.�$���b��b�*E�Wi�OܓI�.����F>s�"~�ե��FklT ���1�e���_�<1 E�\�F��`g�&%��Q�^�����H��^)�(��I���C`�xs��X1w��	�'wPa�f T`���鎣#nJ5ZqGU�L`�= �F���0>� �L��P6���p�xt)E���R���"Z3
A�f1O\xY�E��&��5 T?D!�0�""OU U��AAх�� 'T��DV�"X��'h����Tp;�-ѿD
0��Q�ɜ{@�8c"O�ЛTg�2%���A `�6^��K�A�<Jr�<CB�>��F#�gyRJՈ������N:.�P2�G��yb��>Z4����J�I�:���W�M���'p6QA�}I��xt擘!$�AP��=Kjh��IT��S�T�ܫulL�Tȩs��§�5J�&8D���VjY�Jr,�sd�`�n���n5D��Ӆ�$FI"Q��jJ�;�j'D���d�#2H�rƯǡKo�#*1D��`4��4�p%���D�u���8D�D�ѿ^7f!����&Ke�0)ť0D�Px��Q�4�F��S4YpH:D�DS1!��=�
L ��XQ�Yc;D�l�ҡ�?��lsb��2^3����9D�<�V@�<v�:Q��S�܉�o4D��R2�K�lx��ұ�ѕ��fA'D� �g�X��m\h0�!���f3�B�ɷu<��CE�F�jR\]!v��D�B��5h�m��A3)�*�!4FV?}�$B�ɘG�n���,��/�*!33�/D� !4g����*��0�T՛�g-D�@��dg,���˵{05
��*D�0��0���J!H� �%u�*D��z �X2���5�D+U<����'/D�`���.gX�H&�él�r�2��/D�Ђ6K�x��a�!қ��d��B+D�ЀF��x��Y� �����r�(D�@+�n�*�.ݳ�bեh��	�F5D�H�WƂg��S`�+p�fq	?D�h @�A�3!d��ĉ�^�(�l(D�ȁ�ɯ@��[sEʇ�beb
'D��+�n̎4��L;�K� ~�!�`6D�<�f�I'
��(�dd6i�h�4D�,3��B:F������K�Y1�< $M>D�g��>�f�*��6.�9r�=D�H;�`L�-<r9��6yA�Ti:D�|"�EH�z�{�F�VQ�X�"�/D��eC� H�u�#'[~�Ԥ�q� D��i4aڈ�0��ʩ��0�o3D�0��H��``�I,պpQd�:D��Pw
ٌy%	�k)lڱ';D� ���B>:�6|�f��$a�	zb-#D���Î�>���uǙ�}����4�>D�,�v#��X"�m��O�^X8SƩ(D������JM@�����I�$�p*D�� �,�G��8f�X�W�R;"
H a"O$!s��D;
������O���k�"O`�e��.�v-Ze�O-'�
����d�. ���4��_(����V�RX�&r���NMzTL�a����(��D�c��(�`��4�����&�d�'�ў�~b��3\�$��tO*��$E�h�'�a�d������ �/���+V��"��'�ў�O����G��m��Ð��b��K>ɀ�$�	[��T���q�!�7�v�b�	A-���͓�M��3��~ҍ{ir�hEæN(���ƆƜ�MkR�[-���ȟ0u�")¡XhJ�n�>^�\=�''�/��'�^9�7s�?Ir�G�;Ҟ0��G�,�.�����N�'ў�O/de�!��5h�P䭒���ܤO����e��D���.J���0aW?x2d��҈)D���Mތ?)� �G��E�^=��h)��F���O-� A�73�8d��9S�@p��Od�=E�4F7rTSVm�/u�1ZnV�cFt+�`5�)��Ԑ�k��R��5����jY��)M��0|2� &m�B��R�C^A�f�f�<i�i��5\��D�0r�b�`�H�v�4�Fy��I�n=rwA�!x���b�Cɐf�Q�a�Ot"!�B�3:��!���-)̖���'��5[S�'uKj=�	=_D����	����C��C����xx>7Ao�i��S�'J��B�Ԩ#F����	ڏs�D��'F�Q�a�d/6`�l5
�i�.e�Ȕc�)�M���-��Ħ<E�TH�fK��$�Q9to�J���d�Vec��x���']��X�F0��i��OuH@؅BG6Y�ژ�PG]���D�$}b�L����)K
br����#G� �A�%ɺB�!��>4D$�N�u jq���v�!��Q4�Z�Õ�# ~<1ӊM8#%!�D�?f��5z�Q�D	���v�х �!�DL�Oc��r��$iu �۩&�!�d��}6��3e�g��=��aJ��!�DצT:9b f�������{'!�D�>��i Q1X�|�@ט�!�䛸!��� �ݳ#���#/ 6>!��J�=�$�K�
$f��� %D��4!��;�H��� �'p�`8�
�%!��2DRd�6n@Y��bȴ+!�D�V
�L��Q6/K�������!��h�-aa�^�gG�Qy׭S��!�d����b���Z-��mY!�d��0���8���:nL����0�!�$]�4�JE�p`ώ\<\|��@�*�!�$߻0��X)�%
ƈ�(֏�5!�!�@�k��D��,���H�!�d��ty��k�ş!N����K݁Wm!�DʃoC`:�*�0Ed���ِe!�Է�9g#,
�p�z'��X9!�D];4��:�bG]���`�C;3!��X"O������N��0z��*?!�dN�a̩�t��m���7b!�dJ�mE^l��fMMXA����`!�Ē*5�|`�1�!=3h艢�S+M!�$��q�.ћ�-3#>�|��F45!�uR"h�,O�'�\p���@�9>!�䕯sj�D�Z0�����Kk�!��X2,i��1&DF�w����H�.!�DV2@2��9��}��p*@�tr!�d�xo�� ����-�A��銉l�!�d�7yC�Ku��%���(M�!�$B�)E�	�傠��4GȢ!�E30�����A/�:���/�N�!��W{˨��q�\�Yp�����@�s�!�� T9��+ `0�rS,GW���2"O���0o��BtY�J(#���"OB5�v��*1H���25�|�""OБ��6؆ș֨:N��S"O�T/ r~�HJ��F�_�P��"Op�q�ȄJ*]���F��`5"OP4�bI\+&$���K�A��T"O�8P��)Q�|�aEaJ4Y�
% c"O.�A��?MLH�b"��)�4��"O\p����Bp4�:6�Y�|����"O�@��
X�z�#�H>Z�s6"OH$�d̯|~\�
#�-�]0&"Oشq��	>gÒ��cH�V i��"OV���T��`�(Z]��$��"O�#sC�;H�)7�؄����"Om��ZUyN���N�l��M� "O��	�]%g��Q/;U"F�"O���в���Xg͓�a�pܠ�"O��2F��5K�<2!� &e���"O.�����]���q�L�oe�)�"O�0!N�:| \u��J�ua�9�"O�u��<{����aHޣ-��pKv"O���q%�i�̥�#�ܲ#����"O@Y�F�F�"E�G0��9Y�"O ��Ta�.qJ�'� rA��"Of�`b ��?Ԫ��`!�1Hu����"OJ��uٴ^�9����#6�	��"OB4��L�5��p�$4걙�"O��9� ɞS%�5�d��*����"O�<q�m�5(&!c��ĒG�b;�"OJ��6jK�/�JE�G�m�X�v"O֡zWe�9m��B��E�Glju�"O�a�FO��kLQ�ŮS3#.|��"O��� ė�hzJ�Y6�ƀ�ܸB*O2yV̹E�d��Ŭ�%W �I��'v�y��_2hS�e)L	Oz�@�'ڲ�`��U��X�8��E�o4���'^�u� �M��z���(r@�] �'�5i ��e,8���O����'(T�Y���6!nt"`�������'�~�b�O��D��EO������'?d���`��D�分�H�UB���'O�	8�㝜��h��H�:;�Z�H�'d��� d��?HȲ��@�u��'�(J�㗼 ��y��߱;��%�'�#�i�&7�x<���V27�4C�'�"�~a�˺t� �r@���y�%��,iZ%�O0gi8���"Ϛ�Py�AWBt>�e��!΢��H�<qU@�*m|Pݡ��D(s��5��y�<�tݟO�i��V�Vͮ8�a T������C-0i������I0D�$��EΨz:��*�	n��B�3D�q��	����@BA՞�1��2D���d���1rK R3H8+ҩ2D�� F��@�����1u\p�3D�[��� {4H��w��2�����.D��senٯW���w$ٳS�4���',D�(�d��d.^�KIU.\� �)D�,�Ѫ�x,`O�~P Mrq,4D�l�rHU�@�~�6R
M�&��P&6�T���E��զ~/
�R��=u@�C1���ybO�3v�
=��g��)J&����ƴ�~2�i���}r%�@�?���Yҹ)gڠ���ޗ�y
� 
`,"��J�ANH�г��>yߴ."a{�(�"�`�2!N�|�����=�p?�޴�?�+��)T��x!A�%S;j̀cj�n�<��J؜d�f�@<���H��l�'��V��#
'�1�o�1y��u��H�@.>C�I�Q
 t�%�9[�]PS�S�y��	��Fx��ɂ�	��}��@�DPJ��D��M!�$˗N_�L���
?�Ru�F�aJ1OP��ֺnq8����;�7AO�I~B�	,Z\���)���UC��6KB��[,P�Bd���A�z�p�%�'�HC�	��Z�f��'86��N�sZB�x��Z��"J���b^+w�HB��3i+9X�-�H ���B^�B�Iy�L�r�˔3�`��ڬi:TM�ȓ(("���UZ�@��fry��Q���4H�)�d�y��ȓ	�� `���@�3b͠D.�ͅȓ'r��#�+�8)�iǴ!�Єȓ��,%�	�'��#q]�Ur�#D���$B�0���bNGm��kU�-D�Dy�C9##����A�WR� !�+D��he�њ����:�<�q�*D����b�p*F���
A�le*5D�� a��lѫ� �Y��i %g1D���6 ֱ`�NޯU�t�w�.D����)j��x0�Vp*�
�&D���#�"�`8���)n�@�F�"D�d�w�_�bv[���5&G�){ա$D��y��T�J�j\3�V.-2�)��"D������a��]�-�I^¨ %!D�(@'HG�rs��'�Q�6S���`� D���I�e�"!�τ;�] U�=D�(0���;�(��#O�>�d�Q*:D�@�"��J (驖�' �`b��+D�|XBM� 6�l4����8�lQ+D����Q,D�(����y�Z\ڗ�#D����>�,ЇjG�<08�i&D��pE� >ֈY� 
��zh
�
$D�T!&�62d�ċ��BA��F� D����e?rL@��Μ�5���C�	 D�@kЁ�>Vބ�ǎT�[�!<D��1�cƵv�`�Ys���S�-���:D��O*A�H��f�� �I���8D���w��6�R93���I��R&H8D��hc�S�A�
��v�]�A{�aR�7D�@�D�OBn:��"��Vj!&�4D�d�LA�dP0:�hɯ_��/D�X��
� �Н�R "z����0j#D�����z�� K�G�9Oz,p�?D�(�)0uʾ�
��M��JH�Gc=D���'�ٶ]vlɹ�Ϗ/e�u@@�;D�B�o��V1���3Cv���f*O��¢�'�`%���7Ydh���"Oڥt��(e@���nW)x�}�"O�h�6�%>
���-]�c�4Id"O�H:Bf��q���뢭I?}ڠ���"O&!P�j�A�%B��9ͮ�	`"O^U��Y�!\�����(����"Oԝ�����Y��lڹX���""O��0�咇�� ������1�"O����̵PPS��8�J�B"O^�B!�GK���	��	&k�2h�"O���V�;9頵�F��A|.-��"O� �5��97ް�/�s^Z���"O��{V��4+.���wo4C�)E"O8���%��2H@�n�&d[��K"OaÕ��1>z)��'m��5C�"OlE覃ܗt�,��%և`��i3�"O��[���Nj|��K�(��|�g"O0,�W�ڸ;��1zh�4��A0�"O��'cK0����/+��%��"OV�ss�y���#˞t���a"OF�$eݕhe�(KѴ9�XH�"O|=�c�JQ
>Ԛ'��μ�z3"OUCgG�i�t�9vK�+sl�m�"On��`�n�tث7\�I�DA��"OF%iB	�d"b�k�"�63Q*�yb"ON@�w�؜�B@1#F9pC"mb"O��dG�֒���
�����"O�a�[�Of�Ad�H/|n�Z�"O�1	W�܇!	��0Q��_v��F"OPQs�� �zEb�8qz @�"O�����s�Y��'^����"O�m�ɞ[�y4�ڜ?���"O�ӆ��˚L�D�#=;�غ#"O�5@Z�Ny�T�aڍEЕ�"O9�"C��x�Ҥp���oV���"O~��O^M(�xC�NU%Xd6�z�"O�l���i*LCp�ّ�q�!�DY�B^!@s%�S��I!G+O�V�!�dp���0#�&T�0�! �S�!���954U�G�ZC9��� N�.�!����&�źd�HO�Tr�MN�w�!�$�13�Dy��& �B1��JF�	*)!�#�6A��l���9�C"G�!��ͣz �  ��     �  �#  m/  n:  �E  �Q  P^  �j  �w  N�  �  ͔  ]�  ��  �  �  ��  ��  2�  r�  ��  *�  q�  ��  ��  ;�  ~�  �  ^ � Y �$ + `1 �7 �> +E oK �Q X �^ (g �m �s &z g� Շ � [� �� ��  `� u�	����Zv)A�'ld\�0"Kz+��AI�/@�2T����OĴ�g����?Y����?�fY$E+�)�Lͤ�4��I� `LƝ2��O�7���p
[�U���a]?��΀���iN5I�����}���rϚ�AQ���B�Qb�I���]� Წӥ]�B�95#���$��h,�H���Ei�V����t�B��Wn�ՙfj�2���\�R�$�"��[� ́F�dl�i�"Y��ߟt�	ٟ��I�~K��rK�z[z�I�٘7Ԟ�	П\I@J���M�*O���E�f���	�O��Dɴ(����/C����T��/J��d�O&�n�֟�������	�!y��'\7D}	�,ځxx��*e�x `��{ J�-�~=!<Ol�<�*�22b8���`N�;7�I�k
��d�
"u"�jwiR^}r0O�⟰���ʇ����^�<qTo;~�b��XI�F��(��z���0�D�Ox���O����Od�'�y�iF�"���p`Y[dHH��]�?QÂ�3'J��	i���oZߟ��^w�pQ�Ki�F�_�H����X������rX���^��<Ezr�	�H���S�Ɋ9��d V
F/�u�� |3�(_Ӡ���N�g����3@�5�J1��,d��Jz�l�M��'z���̞ 7����J�;l�%�X��%����7-@)Q���aD[�J���1�B��M#E�X1���aڴO����2�K��ۊX��EZ���$y�
T�&h=Y2̨P�$(UhHnZ��M[c�inVD	�%Ҋ*<&%W��+Ac�%�aˍ/������$� �G �;��� i� �U2Q"`Ә�m���M㥦�x����?^y��Fll4$;�P<z�Ε �,�9��՛ֶi���GB�&��� (�(|�ؘ!v�'D�O����c��2��CB�f��P�lZ�s1�鈔A�O��D�Ob�i�����)�����&l�O��QW�	`�Q���ڮl͆�W��O>�䁂/#����O8���Reƨ�Qd�V�V�mZ缓է�0>~�P���1t�z�x"�g���b刪Sb�����Xyl�;�.�r��Uy� ����0<IU�vy�c�<a��Ę_`d=��fХ߆Y��*ԟ��	͟�&�4�	��0�'_2d��}�[hU�ؽ1e��T`�:2�'�t �T��2�'����Ԍ�O�))�cčYe*�aN�J�N�(��'3�3?v�3ݴ�?��D2��HhUl6��!���S�b�@����'�RjT�}�>yKu���?I:�AV�J �>��}*ՠN�"2M� �e�V ��,�0����9.��I�+U�V�Zx�<p}ܘ��kCJ���g� ���)��� i0�nK�Dr`���Zt~2�ݖ�?� �imT"}B�Oo^��pԮ-� ���J�;�X�����'E�?a`�oΧ}e4Ⱥ�J�>^�9FL_{�'��}Ӑ�m���H�4�y�h��r��'h�8g6������?y����� �����O����O�ʓo�i	Ō�(k��Q�a��_�4��6@�j���$�$*a��JG�������(�O<�bg�#��d[�JߘUIVU[�*�lA��,u��QD�0L�豣A 4��D1Y�w<6��e�'&:��rP�{ �D���i�j�9�����?!���(5�ِ���9�"SR�M� F�@���?+O&��!�3}/ӋwB�LPS%ؾk�Z�Y��O���Ӧ]�ܴ���|��'��䛺��7�N�`�]�|���p'�<��$�O:�ķ<+����<E��S�&��pk�J.]C���= �5��0�0p��B����Oj5�C��@�ɱg�M�op �0U+�  �����x���U!��a�$ �g�P��I�{RoV(`�8�K0'�%���Y �5�|�3��\w��#���'��Uy��S-qz��篔������'���'�a|��ՋC�x�橜�^֪E��7��!͛�Hu���J���\��	0U��x�$G6��4F�>�`���ş��HP̟���Ɵ�l��}!wF�� Hy�l�7|��c�jQ ��Ҕly����s�/I)g���D��j�IS�4'�~H�g^��=3�(&��rB�I�XA(�����i�(�l�՟!dD�$���FJnh���Qy��'	b�'wa�\P��s��'�����$m�D��y��|���i����c� p{r J_���al���Z׺���K�?q����t�$�S��	eg��Qp+T$B���O�0I�m����k����a���Qf�@4�D�a��|�TS�W�6��uݴK�R�����"P��S��;2=�ѫ�h\?Ξ4��_�� -�c�����B��P����Gc�"�]9���XS'�O�n���ħ��O@�A���с���)#��>1�
]�H>�����?�����R+I��E�B��]?3
���U��2�?Y۴�?ф�i�¯Y����F֣'�6@QK�&֨7��O���O�ls�3�T���O���O�]Z�n-�&�_=��aCч�+hЅ�N��X>�A�ӎ<��8@ �|���v��O���vhI�QVZ1[�N�\M��D�}�Z���;<�B�HEc
:�F0�U�|�D�"xλ�X]P�f��}y�d�U+�O�d�#ٴD��X�bY��`�矬�I��4 bεP/pLz�r�p����0�I��d��ǟ��A�g��G�Z-�$z��۹s��d��1u��	�M��iD�b�D�D����|B"�<8"R=0�c�_�p(��AR�|RP@��<i���?��7#�N�O ��OJ!z�N@�G�@�i��(hF����.D��طK�6���5��	}SLQ{��ď�w=|�pp��) �ց��֋���G�R�تR�ݡr��)2�\æy�3F�a4�}&�`�3�˨c�@]��WÎ4����(r������}����8\[LL�U�M�!�.��dI)R#ҵ�	a����$?	�<3��"���v�]L����U! Q򉉳M�V�i���88��x�4�?9�'a�܊aCd#pip�@�e�������O`���Ոur��h��6	��2+� �xaB�-( ��D�{��&�"ᡉ�dX-OZ��o
�A�Z\�ą��A�G�J�	ǐ���!�!d��YItȒx�f��cʄ ��'6��Q�{
��e�<��`˟e��	 �8�Z��$�d��C���O��2�-��*���JɌ��T�'z�6M��Y�J�/G~J�	�՝/��lGyBJ���6��O
����O�y���,vx)�dԧ#@Fy�A�Oj���k/�}���KpX<x�Ȍ5Cl����=.�-W􌻴h��w�	���^�s����'��*�B�L�����E���A���.;*d�E��,%)���Z��^a �wy�|Y�R����;�2�o��)G�3�2!cF��?��H�S.K
8� �3�B>M��R�QiD����[X3��B?��?y�i6�:� [eS��׶R���P$G9SĖn�㟔�'j�Jw�O�B�'�W���Hψ7?� Y��Y	%� �$�~�xX0E�WtIy ��zS��OI�DB�g:�h�'Ď��%�āx��x�Q��
�hrA�R�i�L�5H�:&�D\��!��%�fexZ>bb���ݺ4q����U;Bp���7K8��o�5��$��?H�O��3�D]�`�C嗎JE�4�ľ�H�tD{J?�cF�SAR�yC�]�@���&A�O���䦩H޴���|z����ߩZa�1�����m��%�+}FP�`�fҺ��?���?y�'�?�����g�S��h���"�T!�fD4Vª��ρ�=8�	��kMV
��*�J6�Ua�H0e�^�<&��.V���$(��
BBR>��y�̉';���s�+��V�a�����'�6\KJZ7�.��D*����[���?����hO
"<�5k^� )v���	_n|�� ��J�<a'*]�T�d�*�mŴL���j�G�H�	�M�����KBj�m����	�r:Tyu�	�y�.dH�oP�2�2���󟐪vCCş��	��|��İjd��ٲiP��r4��ح`�>Iyu��R�Ӱ����ix�I??�"p��LZ1�2�y�k̫I��h��w9�`�=O�D���D�`n�i�0Zzj�{�c-�?��i�ʓ5�*9�7�Vˎu�mD�3��%�F{��4��)��h(��^24�H�K�����?!e�i�`ݳ�*�&U$���u�,`�й�ֆu�x�3�P
��i`r�'u�4gU���	�eΨ̺��]t󠥰b!j(����� ѥɗӟ4�'�T>�'�4�υ�*��ת;&�Y;�O��k֩�(El$�#E������ͪbg��P�KP��V����`���� �O�m���H�^���A{F��o0�ݚ��ڭ">�G{J?=�d�K�u߰	��M�R$p�1Wf#��Q �%r�jc>������!���C�"���Ѧ��	ʟ4�Ik���k�M�H�	��t����q+N4�F�ir/΢}S���)�)#�*�ޟ(J���`�9��(O��j����8��A���eu��0�
�F�����L �J��u��J�1�1Oĥ�fGI OF:6�=�L�� $|�P��'�~���z˟�'v*5�B�¶@��xG��8ӤҲ�D8ړ���$zx�� HWy�tT�,Q�_��ɢ�M� �i��&��ʧ��*����״I���`[=eJ�ɆiTzD���`,�O.�d�Of�ĕ��+��?��Q:�H��$������J(��Џ�;N`�� 1�'3*H��a�9�I)�EK�`y�|��Կq}���S�B7x�0AE�L1�����!Tp}Qq�܁&���"��Z�ҔC��'��7-Dc�'8��zy�O�/	*:�s Y�HE*���0j!�D�f. k���}|��V��� B"c��IۦQ�ܴ���A�"���mZ��P�-"�`�F$Ѷ#@aC0X�^d�Iry��'��?��8��ș33�X��Z��~ i�*�rtN���Z[:�Q�HW�G�0)���(O��dh{� ��i�f�0�N(5��(�ʃ;p~��#�#\L�#΅�<t�d��r�ɛ�$��T�}�.O(ŨcaL�\f�}3�LΙM{��@�|"�'L� sfˑ8=�ThhG)R=$`Ls+O���hO���!��ϛ4�Th�� (�r։��M�/O�Q���Zy"X>�����E�pbV���!'��~��	���GE K7@��D]<�������!}v0h�c ��$
�LI4	B���4�`c�[���$�*w�U1��@'RDA���7��ׁߗtc��"��矞�JS@Z�+?��(�# 9�V!W��|YQ��O��nZ�����O�P\jf�$[3�8��(-m��cN>���?q��爟>dq��
�L:h9��nμKQZH��|�^���� ����<ٝO�F �����q�JN,�(!*��?y���?�s�
�\����?����?��w� ,�'h�'�xc�GƵJc ���	D�F�.��3��rGt����� ߘO)�O���Ј��6�rH`7B˧i�����)�`�hr��@J�\J#�R��BU8K?)����.~B�]�yN$q���CIF "�_lWJ�D2?0D�����A�'
2��C�a=���!���Ό���"OnuS4��C�>p�f�>_j��gQ�x ��4���<���[�P���A�]9-!�d��aQ6�\Q#c��?i��?��\��؟��Io�N1SQ?k����RK�C�z s����%8q+�����=���n�? T���m�
E����ՙ=ż "�D�L���iE7>�`��{�'C
d��	U^N�����ը�T|�خ�?�Ҵi�7-�O&��?���?�͟�9�d9;�2�aF4u[�e9f�'�O�m�怍6j��S ^xJԒ|b�hӎ<lZSyr��6m�On�ɃS�<`"d#�>
	��H�I����<!���?q�O����	LE�(�+wA��>j�=J�G�/NQd���KT+n�,˓�*Z�yC���b�'y`���Z�Y�D��0� 6hk:y�d��<![�� ��&LR0T�ǍI�Kc�L�!#B���S�|BCB�?�R�ij&˓>�m�CM+9��)�e��<@�&�@G{��$W��$��@�<�:Y�ԍ�D��O��=ͧ+t��$�W��]���)���i�̔�;��6�<1��Ƨi��6�'��X>�A��� '�9S��T���[.���8S����	�%bY�2MΑ El�����M+(�P�'C/�TxG�Q1SqT��l���Od`�$I>��HR�>�&�}��j��[�8�sD�E�ܼ*���Z~�L��?9b�i#}��O�d�2�3ZB2`{�O@�!��|���O�`��$q�hzb��?1�p%�����M���i�1��,�� K����U��86"tjEab����O����]�P]�O�O����O���`�����D9\AV
U��8�`�iJ�� ��OQм�!o�3Ab>e�2閖/��T�8�� d�
d��$�V�N�r�p�� ,�eO�Q�lQ��ɇ����	3�r}�ыs޽j��Z�L.�E@�6oV,�X2�W�1Z-O�u�r�'��t�?�O��Hea	6it���:v�H�xdc<D���4��|8*��7AϬq�BQb�J�<Q��i>���|y�	J��IR���0X��@QG0~��$ ����'��'����?1��i
��+'8CȤ#F�4d>��s+�V�07�B��K���L#?B�\����b�3������=Ɇ��\�G*$��'?�<аF(:w ���e�"��:v q��OL�6TL ڴ\00��3���;�Ġ�M+���$�ۺS-O�˓iqlU�&*i#~����֎j���OL��P�'"���O�"9OL}C��V�.��g/q��R&X�p�I��M�����Q����?�CE2mv����#Li��V�L��?Q�>�$	���?ٛO&tݪ��(}��nA�]����,�01b��Pn�D�ډـ��~��"?	�-E5���Ԍ�B�8�
v5�}!��P���U�+�p�����/`ĵ��^^��@�F��O��D4?)�i�7~��@TWO��G�o��T��'#J5<�(�s�H,	��Q@9�On��sx�[�1`Erԙ�3?�,�d�<i���)�?���?y+�(  0H�Ousc��\w$�ƴK' {b�O*��C�e���w�_�Gf\�`�ۏlꜨ�O���[Z�0�f	� k�e�2(�X�ZP�S5$�Vp�e7iO� g�P���<[-T\Q%b�?��� ]�7	"�#�J��}�D�6f"?aw"UΟ��Ia�O�$��x�`�s��aq�A�$b!�ā3Z�8�� 䒱/�z| �ķB�џ�����q̘����͞0�J����2w���'=r�'�le 5b�w���'����~�!V>���ӤAЈ�p�{�႖s"-I�.�6i�=���'Sv��A��$�*�ۡn�%kW'�;5�EX�%�%<zv�Z��R�f=�8r�Y�OE��[�W=���)?�n����b��9� ֕Da�Xs�iB"H*x�R��OL�G������F{k��R:�90և�,��ja�	�!��7h�V�@��YȰ1i���)Uz�ɒ�HO�)�O
ʓUr�a��  tPK���/�<xf �{���?����?�������O.��x�F�Ƨ	��`�K�X3�5X�N�W�(0;�]Q��$a�� ;��p�re_Jo���`놠0�� ��/>*y� �1Ĥ�Cp�¹�HO�q6��_x�08�	*8�Z�C�dٗ<��o�~Gzb�;Ұ��� �Y�-ig*�������O ��?�.��d1�	)�~��L8:�	����J�*����	��M�!�i�S�n�Q��4�?I�
�����O�TP2����F�p1���?��B�#�?�����MB,�"��Āw���v�<k]f9#��٩�f��tjǤ	�� �	
V����v(_����3���`��D�r�92;�Ҹ ���F-J.���Ӧ�Z#qO��i��'^b���&B�=�l��R�Ja��6a3���O�����9{��� `Ú�U���"��,�1O��=�Ot����g��B�V=*e�$�B�ۅo�\�hYǃ�*�MK���?	+��j#�O.�!ӁP�~�"@�H��F�x���O���Ÿ5BtP�JP�}�48���I4�� ��롃�.րS��w~��
 (�(p&�TX�p\#���'N^�|�"(�)Z�i�>��k�#0�*T�RIh�	Gl��a�)§@�X�&k�8�b�њ4NU��]��WF;s3
Iڲ-_���D{��'9"=1�� ~�:ԋ�$2�4���㛦�'��'n�㬎
 ��'B�'*�.�&Z�L+@G$I��\"��Y�:tjݣ�iįRI����m��0	vU�Q>�ӭ�'?Ƭ�b���~К5�QJ��4�v��!w8QK��J�Is2�AL��@^"`�� ���O�:��� |��Q�d�yf�� ��J��`�Х�'�� �����?����?�TAnLE�r`���?����?	���?�M~�=y�*�_�v��q�J�Rg
�������Nɦ�2�4�?a�ih�O�\>9:��ɎTq*��h�Eh9��&�S�2�'���'+���'R<�DdS"�
�6p�|�ʂ	H��bU:oVv�k���/��h���0P��9F~�&S;,����gQ 4�m���Vp��� ��r{����I���%H���5C t��a�Q�"����e&k�T�W�͢E2ٱ���8�Ip�'��dJb�G�.<Y�Ώb��\�GF?D���3k�;��Mچʌ/C��T�D=�$SЦa��}y2�_4q����?�0lڇ3�'+
��#��� ���?Q�-�8�?y��?1�U�u���W�݅eԀ��*� R\��4M)�]Q�J�	Ԏ�x������9au'��v���C��#��e�%+܀9�U�(�:*L$yF�Ⱥ_����I�>K���S��	:ش�?ĩ�����GKY�(\�|��F�����O���4�>§w`>Y"`*�'iFd �e(N��<)��T>��ߴX�>%��L�ц���n��$��0�i�J{�H%ɥ�O"���O|�D�i@��O��S�%hTKçH��Qð�O��D�w�����i�,�Zx2 �ف6I��;�O��S�Q�D��J?)��b��-�8�V=�y&�*zʥ����Z���T��i,~̪��?q�kG�~��U{�l)9�X����/?��F����Iz�O}�$۹s�X˒���^>8�Q�Y�xu!���W>:��6�=��x�RH۪e]џ��IO'p?�C�JD�#�( cDάIc���?a��3�)2��\��?����?���~�I����w�U�h��XAK�n�x�ڴ�?!7�\�#J�+�Q�\�B�m�(��b$~��9"�N�-SV��%N�1ܵ����9��b>}�L<�sΎ�-��Z�Ȝ/���21���MC�i��ǋ�.��Y����0,�b�I��έa'�U�<(��ڟL����	�����'�b�In�0�$��'bB6��ЦE'�P��?Ŗ'���d�[$1�	�s"R7Z��q�G�X�)��?��?�����O��S�9�8��e�H� p)��nȕV~t�B4�R%^T�J!���L�`�`J7s��f��.^
���F�˗1h�5���Z�U
%��U�ob\QA�޹$(d�P�G�n���E'F�!:"c���E�F�'%���V�Y�G� 4q����U��d�j��P�"k�9��]��%�x��ę�'D�B��6Pp��`�XƘ���$���5%�HZê ����O�8,������{�\X�v��A�d�O��i�L�OV���O����V���#5h�	w1L�AADR�D���Z@��z�hك�K�����p��$�m�TU{'͚$gc���f�I�t�̰RV��Z��=�����IĽХ�A3RV:�3�,U/��'����;���~�|�DK5hE8���� DN囧�+�d��?���O�1Oؕc�;7�v��Q	¾e/4$Pe�$"�S��,�l�'�V3"@͂d��#-f@�ɳ/ܦ%�'~��>a���
������q:8<yf.�'���"�J#����O�es��ֳfM(p97��B_��p����W>���$�
�$3LB%%��RbV\~r"�)=�T ���$�Rp�癎~b�	�	R(�H��O���Rt Yt���xuD�KPB���O,%!�'y�6�ۦ9�	y�tK	<���U�b۳#���*?��9�Ioy2�'��)�O"�D���
��C%�;˒���J����'^�IΦ	����I�<��TӚ�!BPP�K��ͦ���!�iI�'!�ЧL����'��'a�2����J¬ �Z�d�Old���wmS9���c.8�@�����g�>�A!�)� s������9�R�����q�,�1&�)�����OW���w��>q�	����1���X����Pnʮ�M["_��j�d�O��I-&������ � ��Uj��/�lL�ud�ϟ�'!B�'�?]�#Ɗ�F0�Q�J�%�IJ�lSğ����M��i��v�T�'�Z(�Ш��nt���UdV:�2e�$���P�$��OH���O�d����$�O瓓"������	��˜.&���װ������t��U����4Ӝ�?�R���|����G�N(6��8�b���Tk�|)Wo>}f�kP�&��j��GK��0�D�'�I${XXՀ�	�RLZ�CA�S�hU`�O���'ړ�OЈ��I2]�u�QO�A�Z8%"Oڠ���ӄu��	�#ЗK���aҕ|b�o�����<��l<k~��џ��,G�%!��@�	�Z���C�!ɟ��	3jn�`�	��ͧN��@��i�DJE��m˼�� �>�@�qeY�MZ�H:����OZ�� *tJ��q��D]B%��
���8�� k$��(S>wb@�¨��dR�)�{���	�?i����4y���0C���a|�'��;c�'a|��&BaP�����G��c�!��?���'�� �%[�IpvĻ���U'�Y�����@A�v��OZ���|:0�զ�?�!��v��E�F�*t�뇟#�����O����-�>qP$�1*A�V�ƹ�gD�ԟ?]xT"�F�f�  �ǡp��e���&?��t��m�EC�;�\IÈ�" <�� \fR��ZF¨5�KC�|cQ�N
�,�/����џ�D�T1O� ����
�ixإ���7ot��"O	����F�i�%d`��c�I��h���)�*릴�5c��L�A  �OX���O��I�}���$�O�d�O��}����N�&�
��T��D���4a��i��D
�i�HB��9�ꃴ3xc>}$�D#c���F�a��W	t���ƌ�-by,L��f�xE8t��[�N��$�~�sȒ�/��Mͻ/��|�wFDT�EJf�]8���OZ�g��5�	�pF{��ۚx^�e�3�"R��8���X`�!򤇃_��t�%�Y�|~"�7�ݫ ��I�HO���O��ML(�2'�T�c ��Bt���!�b0���:-v�1S���?���?��'�?�����O1�h��E�
A'0E�����$h��k�E�.>:�9g��L�TH����"�* (T�ȰF�� ����XJȑ�j�u����@�?�"]�)�YW'E�V�qO������(H��@��{o&�裦(#P��'�ў�Fx��S��P�p�$]�0�P0*d���yRC�Hҩ؆�<,_�5���̉��S���'q�	�a��������Q$E�YP5Lv����V>?]d�D�Oѳn�Ot�Dj>)v��&|�
� A�&	4x�S�G*eԜM�&��:�ԩr�gS�"\1G2H�9v�6 +���,R��J�,gQ,���̯%Tb GD�;8�T�R��0�Qc�N�Ue�}�����'����4�T;����N؁g96�K>��.0F@zE*^2v_Biy�B�v�a���)�?���L�YߢA���-)�� ��Gҟ�'l�����'Hr�'��%R`�	4��q�2gCo�2��&�ٿy�4�	ϟ�pĮݲ[\�E�$��3�I�1�O���?�kU'�0��Z��H���o~b�G�.�p=A�HQ�m׺	{�愩B��3b��9��y�'�����#޴ �e���1����'�iA��?A��)w���W&�s	|��D.�~紁���4D�(L�&t @���\-p+8M���-��~��>i*���J���b0���E��.w��'{2�'��б�˟ct��'�R�'g�Κ.cƝ�Q�Xxq{s���8#`�`@Т+;Ё��Ѭn�@���=��P�f����R.Q�S ��@�;d.�+��Ԅ��U�d,�T��$��S"4�	�.h��p`���&�����C�]��T����O��O�(���˟�G{�ŸYS�}��.�!�t}�d�E2E!�dJ"�]p!��e��͈���.��;�HO��O�ʓP�pgj��w��	�Tn�>1�E�^
	Xz��랱J��|��J�2R��`����u�,I�.�2A��8�A.Qh��ʳ�Ղ<J��@G��OJDSn�OD��Ozx���/b�Zt���ڙ
j�iI��
8�u7�ŷ��x¶%_P�8hZԈ���O&Y�%Z_�zd[P]�Е@`�ՒoG
����2�91vC��ey����V��Ex�{gO��?!��ИO9����ԤS�1��gC�1����(Of��$^�:]��`�$��%�b��9��}�A�<	ѯ�-NѠ��re��5�r����dy"��~��'��Z>xu�V�����-nl]H�f��
zl���H3P�ܠ�Ɂ, .M�C�R1J���b��	��9�ПTc>�����qߦ�j��O� "�d�c�J�Q>�1��;D� ��>B�B!kք�:<�'2("�z�-ֲXg���E�j=�$�b��	ܟ���'����6q̄u���'_�JX���I70!��BV�@���-��I�K�cў�C��銵og�!0#!�3v(:�Q��ѧK�B���O,�$��;bliW��O��$�O���@���1%������7h�<UC��L�� yP��xh��f�.sq���5J"z��$$=���4�O��4�B��F2
zZ���M�v����B��]s`l
�?�0��X=n�DI'�O6��R��(.:< �ri5\�6�h���dt��O
��!��y�j�m|i���M��T+`�ϟ�y�@:3�LIX�n�HZL��r��p�I&�HO�I�O˓;0((�S��/<f���ʖMU��:���4��(���?!���?)���?y����VJ✈a���1�jT< x��D�W�%2�\wȄuJca4�e0�#+��M��㒲WI��`UgR�3���11���:Qn	R�bWa&-��*��#�.�Lh���O��
�� �Q�8���5;�
��t��O$�=�����5Tr��Ъ�l7�qE���?G!��#q�Q� �Z�D4YW�A.v�剼�M{���=nĽ�Or=����E�Q(ǰ���� 	p�Y�'�l��'��'�53�D��|�Ul�;X�8�jV��;A`
�p!��):��@j@H�'$��1��A	!HD ��A�^e��A��
�N�|��NH�m��k'iH�v�H�B��
��`�=Y@���4��^�'D!�Aa�oB"&@lX[�C�"��@�'�a~�,Ζ��S��zB������m����+O��	ӧ�	�2��ҏ��H>I`�_�,1��D��������OQ@@��'��[�[j.qcDƖK�D�v%ߪQ���
/�Ը��J"*d��m��'��O��l���Q� %^�jG���.��'[C�$X AB*ИRiOz���S&]�V^I�T�H@�i޲x���%����ӣ8���ھ+|��'��)�I"?� x�N�,&P�z�Ou"�A��"O쨢t��8Kj��Cdm��yFxaW퉮�ȟ��Y�FK<6T�s�Υwcґp7k�O���O�IxV�
8J�\�D�O~�D�O��I�O�@�Q�A1�� ���ĮS��%&�/(e����//�PKƩ�;q�D�'(9�O�`�Ɣ/TK,��B���|�ֽ��( -O"�}#&�� PQ��]?E���� *:͡��[�G����!�dH���:��Rnġ[��ɱ&u���O��=��'�4C�Û�%h"��CH�6otqy�'�F��VLݤePm��P�#T\�A��:���򟬕'� ����|аq�U�2'`-Ц���h1�'���'*��O���'8�	L�%��P ��e{D}��Kp�����=[Flhh���<A�2Uї��C�'o2	{��N�02	+���;�t�f�>l�	[W�=8@�L�qo�UX�Sņ^�OTD�=Ys/;%�NV����D't*b���\͟G{2�I�vjܡS��u!Faxl3u,�B�u�(�u�Q�}Լ�f�*Z|ʓ9����'>�I&�Դ�ߴ�?����TBQ'dHee'��5_eأ���?���?	���?I"�\ K`�0!5���C)�Jȵ1�G%m��}�m�&�����^���Gy��%_�6�h�k[��&��R�)�x�s�Ci݆d��oR%��}*$)�)�<�6K���'.�<��*�񟮹�צߌ@d~�ٖM��v}�YSD"Oqɡ��4h�1�&\1s��� �ާeP��1��t��0& :��m�G�<���?	��?9���i<��[�lor���j} U��Kџ����iU��&T�Wk�� ��9ƌ �\�O��f�xR`ğ4�O�� ��:d�Y���
#+ޖY���~�6���k��扰k ���O:�i�O��ɼ}���$V i<�X�U�)�:y���Ҧ1�Ɂ�|��I�<2k�Snz�AQ�OI�İh�m5bT]`�����C9B���?�ƛ�yr������OX�i�O牿bvu�d��-nQ�`ߛnhh� Ɓ�O���7��Vϟ|�Tc�?7��]��'are�WCJ�¦���\����'�^�a���?��OA2;Or��&���O^�I�T�k� X�)�i
M;(`�sŜҟ���O����9����ោaՉ�?7휒5\�r��ӯ�j�{ �_��;׫�˦e�r���I���sAb<��?�'I��0��͈8~���@æl�tW����yB���?!�}E���O��I��q��ܦ��֎4B�JE�t���/����UCL�-��u3ܴj��Eћ�?��i��	��Y?�Iȟ,3Ĥ�I�p�B�ԧ$>�H�G4�M���*�y������.f�����O6=�	${;�5�S�3�P({.��vRl� j�';d�lZ�g���:ش���#��ߴ\��Y��	�346
��X�:e�Pzv�ۢ2�2�����M�@��+T�RQI��mZ��	Ɵ��	��)�O����|n3H�jR�H6�-�h�%Y��6��O���On���O�d�O����O��SL�
i
��0b- JB�C�V��6M�O��?)���?����?q(�4��ć�(��6	�m��MP[�6M�O����O8��ON���O���;}�H0RT��Z�Μ��%�52.��'��y��>�4��4उY�;��� /��������p�'@��d�^?��C)̬�a�k%�Dc�������xy�R��$����m?�G������?<��u�^x�<aP'��iFq;�F�E�|��OW}�<)���&��4Q��T���`��m�<�Qo
qHw��Bq��
$.�r�<��RVw|�d�Ò ��m��@f�<%n^�H��$b7b���R��Wb�'�r�'`��'
�Ɛ:�Ј��o	�U�zu$@�h�6��O����O����O.�D�O��$�O��d�eT�Lh����;D6"�d�mZџ�������	���������	��I�	�> �r��-�uR&�� �B�A۴�?���?1���?���?9���?A��G\�l�¢�1�0�iѨ�tN蓴iP2�'���'J��'R�'���'lX(8�O
�#Q|�a�R�`�T@��t����O��d�Ob���O���Ov�$�OlIٳĚ:�N�J���ez�����M�I����	�����埬��ş�Iӟ�Sɍ�^X����+�b����V�M���?����?����?���?���?��+� |� �'�"j]E"5�\\���'��'v2�'���'��'VrÂ�Z�ę���z���G�-�6M�O��$�O����O����O����O������~� �'ѧv�4�7�װ(V�-m�ȟX�����	ڟ,��ϟ�IɟD�I��P "���0�[���bκ��ٴ�?Y��?����?����?!���?���>����FX�?�R�+�%��P �g�i��'�b�'���',b�']��'����$�{4�=�6���l�{�a�������M���S�.)��*�X?^l�l�5N��9��oZ�"V\��?��'����O��n�ռwH��b�H@GB�0�`��cC�<�M��i4�d�>-�M��'�?����2{uld�.��i�@�
:|L�O��I"@�c��s	D�``����H��R���<O�P��S!(ɔ��C�6-��A����
�Mkpb�u~R�'� R�ތ>RTm��%W>}D�`�'!��ҟ#�O��o���M�'��H^๚эPSL&UJ�.�?A�<�Wmi��W�c��Q��T�H�l��	��9O�!"�j\�U���#��?�:Z��g�س�j�*3�|��T��=X��O�enھIS��	���!�4�?�/O�)���My�r���Z��B<y�e�a�O04m�&�M��y�@P��Q~�"6;���S��Ǻs!>Ań!S�B�&іQ{2��r��?Q���hO�eP7
G�t��4��,Uk�EQG��<q�i)�d)�Oh�����'�?х������ȸ�bŌϔn��	(�M�7�i��1ҧ,4\�*��8Y���S+H:ыEF�-g䪥�'2��؇�g��Jq�|��'�b�;k�8�ӅMMW8 ���e�:&�r�'���'��'��ɉ�M;��<�־v0D�c�J2>4�ҧ��?�#�i�RP���I<����ަ]��4Y-Fח}����ֵ#Ɔ{���ZB���<�y �Jډ{P�S)O|�	���Qd�,��|�6MD3,�1'��?���?����?���?���)�@Ц4P��~r��!!A_���I��t9�4�8e̓�?9r�iI�'�؝�!h�-�	@��2N�����O��$���a�j�	�'l*�-0��$bwN��`�u�@`���uni ��[�<
v=h'DX�	�$�	؟��I֟$�����!�F�^�r$Kӿr�f���џX�'Ĭ7-�-��$�O|�d=�%LH�U�ԠRshE�i�
l1�T��h��
��d�ۦ�ߴA���i/dN�G���C��
.VL��ˢ"5�u�!��dy��Oy|�ե����'{��� +(2c3�A�(����'���'���'��O�創�M��g]�{�r�R.�P8{!ƚ}����?�U�i;�S�擌��d_Ʀ�h�
Ā�,@C`䆈�P507#ާ�M�"�iͨ�C�Ŷ�y��'=d�H�b�'$V�AuV�p�����Ys��Uk%^������|�	���	؟x��� �Iџ��O�t�W�9H�}�6��@w,h��i�4��'���'��)�~j�V�f=OPA�uխ�H��ã�t�D0�-|�΄o��?��O>�����-<5���6ONT���$6pJ��4��(E�"dؤk�OpHbтʪz�
���-���O�$�Op��ͪy+<���G%�B�E�B�����O��D�O~��2��<���?I��NB��(�㜓qLhLa�D"�?),O����T}R�q�J�mZ��?�*�4Y�5�P�p)����Ϛ� ~��'�R"ٟw�ˣ���E�I�?�s)��9��͓ ϐ`hV�Į ���0��h�0���ҟ��ٟ�	E�OB�dD���� �j@�4��3)�y��0�f0O �DU��%��S�?��$E�� nH�Г��h���G`̟�@�4(3�&OfӢLy��&)��$�O
�@�#S/7�ld��	�#X���d*S7Xu
�VE>�OZ�D�O6���O~�$�O����O
i�aP&sŲy���_'`���a��<׶iv>UR�'��'��OBW�v��t����q���2E̤c	6�__�6�rӔ�m���'���'Jm�צݕ�À '=���ln�%�i�����@�gR���ߧ]��OP��O��Íܬmi8�� ȬF�ƥ���O��d�O��U˦���hy�p�x�0�4OL�P�BT�{
�5@C����m�h�Ox(lZ|�	�����On�l#�M�w�'g҈�uJ�.��qm�6z+b(jS@�>^���ϓ�?	�"�5f'h�J����z���_�0��U�	c�큤K�`�T3���?���?)���?���ɘO�a��ɱ4�]�� P*:��#����\:���'$r#aӊ��b=O��$I����	Qy�F�;}DL�&�y�$YF�47�2��>�A�i�7���^@bh���Oiru�܅qŌ��s�ؕ�R�Z�K^�4>UI�ˈ
�~�O<��O|���OT�d�O0h�e����f���n�)���O��d�<a��i�����'���'���\g� ��O� [�`��.Py����OP@�'�z6�U˦��ħ�js`F�o��8$�Y��$ЄlC�q�@0r ��2G<3*O���Vu�qf�'��V���r���$_�Px��'+v\�d�O����OL��=�I�<��i�1GD�fd��C0 ��>��8���yr�'��7��O��|ڐU�(��4B�<�Ȇ���e�bT�)W˰rùi��7-�O1�I
�?O�y���c�+F�Qm"\"��<����8
�P���� -���ᗬ�?����?���?q���?���?�Οf@�fe�G��6�� P��`Ӝɨ�8O`���O���F��K��͓e��(��fZ2e~���CU�J� q�4Eԛ-y�zM�'\�$�O��\��
W�R��y�,ߙ
�L�v���o�%���TEb�ˤG��@:�QQ&�'�r�''��'o���[�im��1M�H�ꑈ��'qB�'�_�(q�4����'DR&�>=��@�7w�"d�s�B�H��S�$�I5����)��4hBX>i{�ŋ$x�Hɀǅ�.�]ȥ��O,���h,��Z���t��˓�"�.X	0rE��'~���C��*�Kq��g�\����?��?����h��物Y2�]�	�jJ��7L�+;�����E �m�$���MK���4���)�GO2���M�p��Q.�mZ�$��ɒ�4e����="�'�ҡL\�8���߷'!rs�D�/���B#�H�_������|�'���'���'T��'�o�s#���כs���`Dʇo剘�M�5���<I���?i����I�OBq;��@�j����&�;z���#�S}Zt�FqӀ���S���?��S�~6-˒�=t��`�,O|c��
.<�p�'�<ђ�È�v*�dbr�|��',b_�8rdsGE_�iZ�D���)c�'��'�"�'�	��McP��<�� ����^�xR��Jq�r��'pt7m"���O��'��7-VǦ����b'�u�S-S��P�z�B#���b��>դ�&�e�檖�Mx�dK~*A��6�#�	4{z��I�73,�l����O���O����O����Of"|�lXD5�m{6OìG��5�ş����p�ݴt��$̓�?�ҵi��'b\���/��
��MR1*�$?�I[$��O@�1��ov� ���P}ޘ����pe�T�풬p�-�d�1�G�;~����'�
{�$���I˟��ܟ��	���/Dr4�y&���5��M���ҟ��	Oy�nlӄ�Rw2Ov�D�O��ii>��e���k:��V��HB��O>���|}hӼdoZ��?�O|j�'g�"�*�'�>$�x�b���64j�Ju.=2nmKT)����a)1*�$^b��O�˰��5��Iq+��((��i�O��$�O&���Ob����E��FG�]���c��, XyȤB@~��L�'���g�|�O�	k}R�f���P��x�ܒ��#��q �D����ٴgv([��L~�F�\���%�ɸ}��ӌ�T=s�W5H��83�4DL��Or�d�O*���O���Ob��1ʤ���CR��C�L�|I��[����M�a���<����?�����)�O��mü���A�E�В.8~��#�遱�M+ҵi����>1H~z��hy�����)��QE�����+L�p���O�qY��ű#����1i:���O��D�O��d����`&��(��}����e�b��O����O\ʓ}R��cK��y��')B��`t���m�O|}����3!V��ɢ��$���}�ݴ��R>�pv)ս"�������Z�lUXu��<�A���M�iu�/��'o'��a��y�
\Bt�`![�j�,[.��?A��?���?!��)h�8ku��9j��Dbe,��0� ����O$Qo��I���������4�?y.O�9�����6��kk}��m�U.�O�Mn��M۰�i�H��Ď5�yB�'f6芄`�NrJj\�@Y`�I�ݬC�E�Qr��'�Z�M���?���?���?	�IӉJ��i�C��{:L��ʪ��D��y���r�(�I㟔%?e�Ʌ)��M�K��y+3�2Eh�O*�o���MS��'l�>�D�+=���K�Ղ�`iXѮ,�3˔Dy�#�2��y���Sy�'���'x��[�h�ؒ��I�8��,�F���?���?���?����d����hcd�(sgE����U{���d�"%:dnǟЋܴ�?�(O���@}��uӒ�oZ��?Q�M �d�ʵ�Z�bV�	C-H�SF�!b*??��7��@xcd���'K�k��5��k�G�<�|��N��C6�$�O>��O����OV��.§z�pP�Y�B�)��B޿-� �	��d�I��?ђ m�\�ɠ�M�O>!P�D�n풓�ޛ~g�-����.;$�V���4y��F�OB��	�H�=��I	w��Ō��	6pd�W�*}k��b�M��ؑ�ec*���O��D�O��$�O��DV,\��@��?�h��BՓOr��d�O˓I|��lV;�y��'(?��o���eyc�׿2x����@�O���r}��g��oZ��?IN|j��y6b ����?H:���	-�H0Ac#N%Pߦ��֤I���꟢t�u ڒqD�O���僬��VL�b�#Y�j7��'"�'h���TZ���ٴ�&Tɐ��?X��t^�&�<1 �H�<�����|�O���#ٛ��Q(O�����הN����T�I�"��7M�ߦ�	�Ŝ/%�����4�cF|9ʑ�R'RSyo�v$�$������>�"��	&�Z�M����?q���?I��?	���i�%�xT�h�2���bʍV�7-T ���Ot�D3���OH�o��<���^�s�Z��Σwj�ݛš���Mk�i�F���>����B�'|U�d����<ipc^��$��pJ��F7�p��ż�?9aMJ)q�xi�'���?Y���?��8�t�h& �:3"&5J�.�6>�d�h���?����?i)O��lZ$���ʟ���<L"
A�ǫ_�%/:=�i�T@ �&�p�I1��?_�i��K��O!d��ׁ�1�y��	� �t��{Xk`��4Z�؁�w䓓�?a���u���0XB���Dw���$JR�eU�yS��_�4a��n�O^�d�O���O�}��'A>@�F'�[��x�l�;S�ݓ�zG��Ȗ��yR�'��7�O��|R�'p��(@���:�^����܅K�0��t���v�B�o��Bޘ�%x�@�I }-���5�ֿM�R� �nCr���P����Cb�b�����I⟴��埸�I��I�% �X�B-H��2��0cm��'�r6�V�5{�$�O^�4�I�Oj��4�%&���
Ph!^��r��[}� z��l��?qK|
�'�2׭��а���qp�x@բ[����B����d 1Ԟ��&!�,4gO����O���1�"]N�9 O]�uc�.�Od���O��$�O���<Q&�iQڐ3�'s��2��'){��AB�&T��9��'��6��O�˓�?�A]�T�ܴm4����O }C��X�~��VN�*K TD���@�X�ٛ'��BE�d��5��&U7X���?�	\cjh�Pr]�@
B�pSJ=&[��Y��'���'��'��'K1�l��A8&�4\p���)x�`���^�g6��O��$�ݦ��Gly�0�ɽ�MkI>��hÅ$ttzDe��4.���JO^��P��8�4k���O�8ݐ6�ʐ�y�'�mQ��^5��(`��{r��q2.5ql�P`N���'p2�'�R�'�r�'B�9�N�XMl���Β}��胀~Ә�mByb}�0��1������O����3����E�N��Wi�<���'q��jڛ��q�N��	W�S�?�`�r|�BZ�z���Q�d
�I�!C�% �Hp2Ԕ'���CM�<�.����|��^=��we_�k���)��\���'z�'����d]� *޴΀ ܹg�V�hB8��LJ�:!0�����y��'��7�1�4�ƀ�'n�6̀*7<�ܐ`�3"��DS ��m��8o�M��e@��,��?cC����m�s� ���˞vk.���ƕ#��X����|L����Ob�d�O^�D�Oh�D�O���)�@E�V���Ac�]A�c0)˝�M���<����?�J~r��7���4O�T��)-C͚���5�(�@gӺToZ�?!�O��������	^NL]�18O:�A� L�N�R1l�X3t}��$�O����2\�f`�0#:���Oj��O�����c�$�pg[�C�"	�6�1J����O6���Ox�G�6��$�y��'h�D�mG�I�D��Y.TA`c�eDbT�0�	�����ꦑA�4�V>=r��>d���T�~����O��Ć4
@�(W3�|���CJ�\?�I��'�Ե�0�� $������9~�!����?���?1���?�ȟ�@ʀ�o���I�>��i��R0������v����^ʦzP#z�p��'�MO>�'�
wJ#7�(���Nâ*��l���P��?q!�i@N7́��H EO)iG�$�O�ța�7v�����
H�:Y�s�C�Ԥ5*��R��O����O���OX�D�O&��O�p�0#N�`{VH���<@sg�<���'EȀΓ�?����'�?qҨ0D4�I����U(�d�Q�!�I��M[�i����#�������
�xYC�F����!� ��C2�ۖ/�ʓvP�jDHĊo]ּ�I>a���?�1�X�/�����ψg�lݳ1`F>�?���?q�:�f�K|�I5�Mc'�L?���[�<�7�V";��"㟭�?�ֲi��'�҂�>! �i�6�ȟ�xs�_�
� �,�����n�
#|��e6O��$>���)�a�	w��˓�����v����a��b�&ό\|L�У*�O>�$�Ob���O����O@#|�_1��"č�+�6�3�&��(�I柤#۴F~tΓ�?9`�i��'JR0����|�uI�Y�<�1J�ON���A`����I&o^���7O���P
";\$S�C�*�X���:0+�Lk'��"pE�+�*���O����OB�D�O^����8��j�`��ࡵ,:��'I"\�p��4-Tv\�'�2�?]A�C��ʔ ��$<| YQq�O����m}DfӀ�lڶ�?�M|���qׂ�q�p�<�cE>;�*Aas-�^������꟬���d; �p�O��� EYL�D�Lџ$�R|���O���O���O$��P˓�&O��}�*(R�����xP��K�cr���'j�F�Z�O��Z}"�a�&��i��T�P�k�>y"4f��Ѧ�[�4ap��O^�<Q��N����K�>����/OB��E���@��`�F 
3h Hqғ
�O���O����O���Of�D�O��'S�� ���^-'���yq��'zaV���+���ٟ�	�?�Ou��lӈ�b������ʼ��'-{���m���M���'����?a���?�u	��[���=
�6��1&^���᭍�v�D�I{��޽{�t$���I��p��̟h�DH�o�L5��+��l6�j�.�ßl��џ0��{y�}��LPכ�L�Ƀ�԰k��=&��SK�{�t�$���ɷ�����*�4uIrV>9�M�\�YK��N�d?x�����O����$Q��jB<w����2��Y�|]�'�x�� ] (=���ct�����?���?a���OØ�C��Δ�y�� ���@�;@�"i��	��?�@�i�|[�'��,w��O��l1��6��y����A��4��O��mZ��M��i�pq
��y��'P"S�� �5(�؈�a��b~��5�Ķw^��YuC@�$���I�����ԟ`�	֟��	�`��A-Jֆ ��� 5��DB�Ky�b�f�	�����	�?	�O?r#Ϗ-��aԪ�uB��§����6��V�x�����z�S�?5���B����Q����@�� G�`8�a��<\$�ܕ'��xc�
�z�|"|B�'��aLB��D�1J a��|�䃞�m�"�'��'q2�'���*�MUOR�<鄄�0P_V��d��9ކ|jc/�?�Ѽi�R�$�	���$��ܴeI�*� hv�uXa��}���kq)	�>��R��<�����1l�>kp�t*Ob�i[�����6a�b)h�"�q7|��X�?��?a���?���?��	�:e/dܓEM�;XM�c�놪UY��'�"Ff�b���:Ov��
ئ��	ly��<S� ���[�j��K�9e9��$�>�i L6�䟌к�3}�D�Oqt"����Ӗ%	�R.��顉�	;k�;���?YD�O�d�OF�D�O��$�O�9ڃ!ͰH?�`�	�,?疠:�f�O���<���iC���'E��'_�S�
�!U��X����d�E�N:���O|�'o07�ئ�[���ħ����)E����U-����F��VJ���d@�&��y)O"���4-��k�i+���f���C��S�{��	@�����O��$�O���=���<�v�i�0S���B��ycc	�\OF48�H&�y��'��7m+�4�Z,�'�6���V��a��F �pc��?K&�l���M{t �g����?q�j�*b������D�(L���h�;��i�C�8{N�$�O����O���O����O��$$2�KęZ�5��G�r�������M{w�	�<a���?9H~���?ț61O��:�a�_?�@��
�,�&@bg+gӰ�m���?ѪO������IИ]E�@�t2O0�C��%L��E���01�,�r�m�Op\���;�,�1�-�D�O ���O�D��.ʔ1K�/ȡ�ph��E*�f���O���O�ʓZ��6�P�y"�'��I��O��q�f̘)8���uM�p��'R�>!��iD7����ĕO����A���p�$�	Ld�@���?�����F�8����Ƒ9�Ǚ��ɕ`�P��epUS��/�T���O>���O�'�ӊD���bm�� � 3+�@t��#��H�d��+�'�t6��R ���O�m�Е����O��|���?�����l��}L�c5�'��7-�Ǧܴ�h�7��<�ߴ[� �1���*j5�<��+��%X �2 �����-�'0��',��'{B�' ��'F���C-?3^ҡ�� 	-Q��W� ��4-.P�')r�O�ڟ�*����Ę���֚��c�'³���L���4|-b����O���-z��Q0�M_�d� ���Z,!Fԁ�k]�6��	�k�hKr��v�`'�l�	�d;���'np���������H�	ܟ��	�x�Ixy�`�h� ?O�� �`Y�r>.��!�
DnM*�M�O�o�@�I�\��OB�mZ3�M���'3�UV�ܲa~�=�o�=O�&��N� :��̓�?!�n�(s<�06�ֲ����DŬ1c�>��(7X����&_�_�����?����?���?������B�G��l؀�ԏu�p��'�b�'�(7�B$��O�po��\�'�<�c�?z?�$�ȑ..���JR��O\�&��vӮ�I�0�
�I�4O��d�c$��9#���`)���6^�x�aX�
Ir �o;�D�O~�D�O��D�O��d���Yz@�ԯ;KH�IL�2t:�D�O�˓,B�V�O�y�'8b�?噂�L*����`�Ǡ��v/�O��Df}!w�R�l���?�L|���RSZj7kL5M�܈� O�&Y��y0�]7Vq�8��d���d柺�p`�g��W�|��K -�*d9�eVd�v����V��'��'1R1�֙�􅉬���M�Ҡ@;�n9UD�P-�p���?������|�-O��lZy�ށ�pn�{�D�"Tg 7i�ݴc��O� &�A�'!R,�)�lA�bKP�d�I�W:*��v@�PS��SoM�,����ȟ��I��	П���ٟ��IR���U-j,��LP�U�̩4�nC�����y��'�"����'}b>OQx������AC�H�6.`��y��po$�?!�O\���d��:fr1p<O~`:r��'=�:a7�J2=m�Dp���O�|�Q���E��<S��$���6�'"B�'Ud�H���;TdS�����^�3��'��eӦ,�G��<IĿi�V0r1�O�2�'��\�s/÷B0vxKC"R\��[d�|r�'I��-�M�#�i.$7�q�������t�b�
{8�"o[��?	��-(��!%'V�o��z-O���
�m�����z���ߞl��P&��'RRP"Wi�Od�D�O����OX�}�'
���V��" ���d��o4=0�xf��_8�y"�'�07�<�4����>R������۳	�t**g	�����QY�4Jv�K�����'Rˎ|�q���_�[N�8�1�ީ�:�؇� �A����Ӕ|��'���'���'/��'
���6`xa Q�Q�pĊt��ʁ�0剏�Mcr�<���?�H~2�J�V��� S����bIԵR�D-�/O̅oڄ�M�5�'��O���Ox�qI��'5��1`Ç�M,T�ñw��9�\���p䛹.�.���)T���'���'����<_�F��!��~���U�'���'%��'e��j�_�x��43�p�r��}��t1 �S=�0y��G#H��x+��?��O���{�D�Ӻ{������_w�Q	�+�?�еq��
+Oom�C�P�pݔ��'P��	��Y����ȳ46��O\���p���L�>��!� D�_� �Ra��Οd��П��	�������|�S6/�R����?��/�
=t�s���צ��������4I�6�͓�?�Ŀi��'.��T�or���`̺'9r�q�nmӈ��'�R6������09�>��Vkz���	34Ɯ���n�P���a��U2��[`�*��&Ea�	ޟ��	����韌�	���X;��(#�@e�ݝg����I��'L�7m�ik���Oj�d,
�HW�&K���Q'ӏ ��I!b����	����ئ9BشNҔ��O�̑�h�L%��blo�l��/̌']�HQgTJW��?���$J�RI(�$���Eʅ�x�@����:��؂BR��8�I؟���ڟ�&?��'�7͉~�,���L�/O���aa��1$d�PH=O��ߦ�$�擟���AצY�C�42�Ly0j��N9@<`5e���M�w�i<8���S��yB�'����#�I�h6�qW�$K�B�4B�|tRG#M �v8@�%���H���D��џ����L�IFy�O�p-�#��M���poח��)ĺi��Ax�'�'��Ob�'��Q/2.���e��ݥт7M�צ]�ܴ��I�?���?Ͳ�ePw���$�� �h����H:S��4��@�$��,�?M߈@&���	��D���H�w���lsusM��B���@��۟��I埰�	Yy�I}�:��?O��d�O`��A���D�j���r@�����?���O���'
�7M���5[����I_�O�r$įt�TܳcM"A�"�'EB��5@p~aK�Z����<J��Ʌ(I�<�w�	g	�E�G!J9�@5��������	���	ܟ�G��;O� �Q��,��[�¯ �x��[&���jӒp�2O:�$ۦ�%��S�?�	�(�+B���f�*G���s-Gҟ�k޴����q��i����E"��O5*jΌ^A��ږ�R�b���m��w�����# SĒ�A��[��DQ!FQ�ԃ&K&��dJ�^1��[�lϑP��@jg'_&�!��)����� �u��+�O�H��E�2	.A�Π�F̼<\��*Ԫ^�8��0�eo�]�k��H�T�¥)��F�r����o�)\'j�Y�f�&v؄t�T(H���b5#�s.=���M�^�J�!�j�#H:�p��o���aE�ڋՊ�3A�	P}>�&>+�@uʗ:,If���Cd�D ��$xv���GA�t#!�\����Ȕ�G=+[��ׇ�)���AkE�FmD�Srd�{i���c���.d��B7?s�@�V��5��AY���- �@�	 |6@�*q��K�l�¦�;
�p"��ƪ`��p��;4XRIC��*h0����s�̣C� �A(�ǔ�M�
 #u�ΜtG<i��W�M�fɫ��`�����O&�D��f$�@�ɘPK�XR��_2~Y.9!5K$&f��	 IDy�	ҟ��IO��\>U��̟t��'X�$0��ca���~GBxE#��M[��?!�����&�xr�'K<O�U�p��<m��
�C��h��2��'a��'�e�
1���۟��	ޟ��H�e����Xi�Rf�].x���*)�����?���L�$ȫG�Mm	�LRӋȐB�\8����?���&�?����?I���?����?���0\9Pu�W�p;��*䍌w�~5��
 )��'��'B�'��'6*��6lR'a���7�@�m_
-@��@�r���'a�i� ���FƬ�A����e��Pʰo��=��{�F.E����M�i�� �A͸z�P0���O����O���<)%�E�?�����K��d�>!�1��!9������?�����?����?Y�Oh����
3b���96�~8đ|��'��6�b�6-�I��H���?����)G����d9����;���W�\��490r��R}��eȏ�o�b��c��eګs��I2�+�;S�R�f��yb�N�m��=s��-<x���<��ay8� @�"|���	e혿ov���
�&Yb�ݚF��Y��a���i�t�?�#�$� Rވ
�ϛxK�H�RI�-,6J��&g��&�d�!��!$�L�b""�~^ \!�XB`���pW"�v�c��@�\�i�����%�(�ks-I�Z��FG�v	p@���)	���IΦ1���P�0�x�$L�*�b,ae�?�� |�-�.�Q=���m����!�	ֺaN�ҁ�S�i���[e�@�^�I�M�4��U�S3CDs�m�*��>� ��E>��`H
�F�8����>yU�Kܴ/�ޣ|*���M�j�4;ج�ZC�[��e��m�<���U�U�C�N���2���p�'栢}�T+޳r`����͘*`H,`FeI�c���	ǟX�I�N��LX���d�������c��N�&=�漀� ���(����1��]����O*���̓		
b�c����7�	Ly*!T
�s���`AfU�_�@���ٟ�1�+O7��Pe��P��Y&@��K��ۼ�d�ɥ$p��4��2M�� dٮH��G
�p�		i���?����?a޴:�x	)'�<&ˀ`V��w���V��=y�I�g������KaF���3������h�'�Hx�EjK<7�n=��L3R��ѪÎΛAN�-��'M��'��Kk�Q�	П<�'�M��.�ڌ����`�h�;1k�R`"i�����=� ޼ͪ0)�gH$�ڀ�f �H���e;L�C�{Zf�oڱ}�Ha�$L��D'ڹ�4��;b��{p�in�7m�O"˓�?Q���*���h����(R׉�Z$���	m�����g.�R*@���c[	f8��O�}o�ϟ��'���`��{�t���O�7M�1��YSSc���3a *z����mOL ���� �ɏ�\1�"H9��q2a��H��]a��V�:l�O�41��qÏ�p㑟�R��O�I�&G5�8'��%l(�9%%$,p��@v p"H��f�S7��c��U�IS7��$�զ�qڴ�?�_wȔt� �QA���%m�:f2=��'����?�'�� ��}�:��T�NX��-�j1�	n����wӌ� U
�ԄK��?&Y�s�N��&˓G/>]�׾i���'u���9��Ʀ�����Tﺀ�&�/l�\Z%��
�?ɵKƅ-b���kٻgB0,�E��.h�t�Sv�S
n.59zU�b.'�8-J���>i#MDJ������\U:��yk�%�h���h�_���'a��`���x4�@�x)�Pa�>)����1޴ ��Ov���|�C'�3~/ ܲ�雌E��3q�>����=�⊓<d"m�%�^�r�*�q�@�K�'Q�"=�\w��%�i�Mw$���� RqI!J�O���Of4	�c�)�����O��d�OnuI�w���Kg	�D��Y��AKR��(��-�RPtB7mq\p��o����'/E1O(4ۅ��GBt��F)�P��:�a��](|qB�s�\�)!�)+��O��=`E�5hg���)�"�"e�N5P���ӦC]8"B�h �i�R*Sz��eDh�<����M���� Z
*�z�K � P��d�<��Eo� `��J�>4<��SV�U?���.{p���my"�ř\.ސ v�҄&ib�)��T<a�R4��H��f&B�'�r�'0��]˟8���|r#�7�5`����;�&<2d���>ؑ��pf�ِiƱqg$���I���So^�s_��zÅ�j�L��ǀ\�N�$E! :(��ˀs0��ɅhZA3qO��Bt�i�$Z��ӔQ[T�d�0i�x���N�b(<9�N�1��,��.x��u��Ej�<��k�&m9�`�P������~��ɦ�&���v�K��M���?��4֞%�߯���r�ɏE���a�'��p�'���'�툐	12��t�Q�ǏU�8���+�N�z�"�,�6p�l�"��Q�_S�F~�'�*\Ǵ=Zd��d��5S��ڼU^��jq��sO:Г���:�ΡHW�7�M�5�śø'+��O4��7�i	7�y�F��%w�l��0��\>�h�Iş��?E���^�#91��E"��(6		��p?���O���Ϧs�)k������$��ceyr��� �H6m�O��Ļ|R$���?i�4~[P���g�RC�Y���? ����'o�mQvC��ʹ�pE�ns�!�v�[RRO|j�W�~��DCcj1j�m��cP}���CDI�@*�.�r�	���#^FE0�X�R��π R���]�Y�J��"�R�/����]��W�O�ym�M{��H��B+@�yl�ʱ ҺшԒ>����hO(O�UA��ѿS�X�àH�h�*C����M�a�iQ�'A�%��ѐ d��� �\ ���+b�'�D�"7$���'���'Q2��ü�i�QIDB4�^�{`�Q������"���'�,e:�Κ�/@,��O�{��=<nh�蔋��]^�A��]����I4k�L������g�4��9����;�J�z���+[jPJ#xӖ��)_��d���gy��'����7��BT䖤#k�G�	$�y"�+)����F�p���D	��~ҋ)�.� ��Byj�p��������_ri�#��>���'""�'n���?�O��x�B/RbT�ƌ��ev�xbn�:6�p��Cjj�Z��45�f(��[#Xа��rJQ$2���I���7m�ڊlI���%9�j��E#�0~����P�	Hy��'��O���>�2�۵ǉ�"!FE81�@�yB��'�.��È *�dz5�"��	�?C���<�~�n�O�$p�Za#&��4'�|����s�j0J`���Y�nV˟�	��`C�EF���y��s�*�bs'X,UU(�+EnJE1`P��#�6��m{A�I�E=t�2Ŕ�?. �V�#��Y#�U�6�N �"EДP�1@B�P�IhslJ�QqOk�ɟx��4MS�6�'��ɥj���1��\�t����){�$�O�㟢}*���7s�y1�h����J�e��Di�'.4�N�+w�Z%��K�6gJ��j�b�<��a²L�<)����?�*�v�"w��O 6mXRc���˃2 F%�7��Nt����%���	B�S�L>���U�E����A�z3J�q}����O�>-s�%?+��:�o�(�*6��>a1d���QI>E���Q;��YP���a �р;�y��v%�1��ɧ�\ڐ�T0.`�>Y��Ӡ7�`�@W 
�N0J��2�H�P?Xr��?���%O
�Κ#�?)���?���_>��	����F��.P^!)b)F�G���q�)�	k,|c�����C���� &�ɢ[�y�'��;�θ@7����`����O��q�BM�*؉U���b{��"�M��gB$[���dT�\kѼ:�2Q�eF�[��1������.�՟��)�,O��diӚX�!֒n��7n�<q8�V"OR��Ҩ߉[��5-F ��\��%�ʟ`C����P�Ġ<yנ��o����s���+f5��D�5.��ը�F,�?)��?a��`���OP��}>)$E��5ʰ, d��Wt�F���8&�Ǚ��k�0�<�BB�@Q�'RL�srF���-AK�4���f�]�FS\m��[�*�	 �ő}%0q���^��=�
E�!Ä#�$*��#G�x�l��S�	��?�J>����?����;�vl8�ŀ�y��`�I�9�^���t�h�jv���:��P �B�	�Oʭn��ԕ'X,��Ou��D�OV7M��x�9ٖ�ۦ]��؈c���V�y��:_��]��Ο����\��y��^�M�T0����-7<���O%�V- �}�>i�7L{�PE~�V�gd�����~��BD�}A����H_�3�VA����;c(1������P.�hܓ~������MK!�i����ny�f�^-)����Ph5���OJ��5�)�'��=C��ډJN*��舝6	�����=�~�#�d�`Pg�Q)?vt1�|=˓x6�����?i���i�}���`�\D�!U {]��`! SЀ�E�D*��56zB	03'�S�\�+ŧ>L:��-�	N�[B�!T!�/$h��t	4|��5;뢑 Ci�;��x��(Yf�r/>f;���p�D?,I@g*��t �Qʱ������:S@b,r�p����)矪6�3`�H��揋8[���a�/G�-!�d��T�ޡ�]-Jl:�N[0 �IG}��*�'H�dAE��Ac�<+�O�/f��(GKV���'���
�'�ў�)�a�С�lK)�*p{�#֍|�!��v��񃥔�!����1R�tP��P�8WT�a��/|O~�)F�ߞrmbX���5��1�&"O*��j�� 
�S�D��t@��w"OJ�I��J�3��]� ���	wH��""O���v�B�A5)�������"O���f��=������ڷy�~��v"OdQ�E�n��+���p��"OT�"�LA<�y#���Ԡ��"O� �qE'-�� �4�ؽ�$}B�"OL��ʻ)�ph�惨
#��1�"O�Ih2!Q<X4��K� BF:Xf"O����L;OnXH�oC,$`��2"OpC�K�(����1c�.K�ES�"O� ��!h˜z�� R��\-�h&"O�Akw��0U�X;v/K's"U��"O�P�q��X�nhqpe@�{�	"""OҤ��]r����n1�}��"O����B�#@l ���&�����"O�I��DC�.wl��g�/>,PYyv"O�����<pJ���fE�jh$�S"O��j&��^QԸ�	C � q"Ot�#���C\yaύ:�<���"O��0��Y,,�v�x �S"
��(��"O�X��cJ�	 3�$O9<�L�q4�
�H:�*� Rpy"�@���BL�0�RQ
�%i9��HAHHޡ�^��R���6Ra���� �2~&pZ�iE!;�d;%扞m�zB`X`+)���Ұ��e����<	r,��9,�q)SK=�l�4,<m��U@�ЊU�mn!�$�8�8TI�k�18�pRJ�l7�cr��䮔�H�dPF��I��>�U�+v�"�1�n��y$�f�(Z0 Tl�B`[l�6DεQ�O��І��o)1�1Ozƨ�)�L�z���+fH�K��'nZ23۰����,f�ީ{�
�%#i�C�ɞW`�%�
 ���6M��5��#?1�@o�O`D��p�N.^��XvK�5
���b�'!��r��
E�������K�OR ���)ҧ:=�]��N��p�@j�1H�����{�jE��KJ0�ndz������O�����3lO4���@ ��ȉ��)�@�'�<��P�i|yx�'Z5�Ȼ��݊
�'<�1���L�Va�`�",C�8@��d�^n�"}b��P�a�(�����f���;AE Q�'Ea�t�M6l꺤e�]?tњ� ���~�E�)Y��O�>�;� {����ɑP+����O��=E���^�f Ё����i� L8}�3��ۓ�������5`���e�֧:���'��z�	���G�w>(u�׋��o`d����y���M��pK�L�*����)��O�eۇ�.�'�^Y���u�z�SuL�P�Q��AP���,$�����ʉ4B�����n5����)��U-��hdGy�L��U��)!��܅u��,�R ǘ#f!�f�U_�0:N�rۓA����܈:��mp�,̀�����!�In�Lj���b����a��K�V�VC�ɸ>~NYZ�I����2*�Kc���'|������OEV�%�%s� Æ��>GB�9�'*�F"ڇ[6 �DfO<k��Q�CM��~�A�%0~�O�>���ޫz�.] rOV�&�q��&O�#=� jN�,�<�q�l}}9�(��j\�f�Z�;
ۓ9����䈑�I��㦭��_N5�O*�=��L=�s�i�d�z��\+e�sv�jeYO�<���_`�脰`�C�Vրm�I�Dܓ����a��֝�)�<�{��_�]�qj�'Y�W'>B�	�pXy�� �-s�k�#j���Dx��ɀ�L�s�4�]�MN�T�!�>1�i����Ni�!�U�O�1OLa��'O>ի�k���d����k�j��'��ݳ�Mξw!0B'�ʶ Ȑ�fO�z��B��>nh(��`���	��Q�l�L=p���%`@	�<�tǦ��;b�1>�Pl�˘ͦ��I;"�^�<I�K� x�|!�5��a�^��q�PQ�I.a�Z��A�|"��ņx��x�'q�P��i�Hd�D$��@��p�qO�� �bV�_�l����)9v=4�AwC�)��'a��D�,O�i�!A�B�֥�3퓛y*f��B;�	�9�P��L<yQ��(M�&hi�e˳���`�@M�'��hq��h�OHqzCN�����m�8cp��#��%0o�Ą���!S�P��fV8*��Q����{��
��knb��J�$�Onh���I�U�)� ��s��g��5�D�g[��{�"Oj�E��`TՊ�E&l���H%�i��أD�+Xր����W�jEXl�N?��@/�8:�t�yBF�� ��"+\O����M��K�L����=h��"�#T9[�~���nT=$�Y���%;iaxR����);0�Z�)�ةj$����'�R%"�C �F�,��.YA�O��Es$M�? SFA��e;�Xpa	�'F�!� 5A�����̶NE�d��`�wDDc�:)B�M�����~�t)V�<@���	�F�2+v�C�ɮv�n�I!�މVꆌr�B
�#X�r�-F���0N�*D)���mY`�A�"喠aG�K2)|��D�pL���#�ؗ4�d@��B8�)؆��%j*pA+MڙS�B�I�V�n���ҚR���	�*Mo��b����Mj��H ըG��Փ��^��켺���K^�ੀ���P!�D����2aƸ<D)w�.1��s ���fv�C��O4�:c�3?���H�ڥq�Є!	x�D��d�<��-/1���s$�;/�n��E�":�X|��.:Jj���I����<1b�Τ!�ع��~���б&�]����U�=F�r�0����xs ! �Y���� c Yl�Ptq��Bh<���\�<P-�Ud.ir�葆�L̓ix���>���3���OE̬�UGU	!��;�ɉ��L��'�|j�!��0z�{R)'}�e��*��cv�Kӧ˰&�B�Q����I"'[�A �6g`Di���B�	�"<v�:'�~�ə��Vꪠ9��W*p�0��gN�K~j��D\R���#
��D0�Pj�"w��z���$	0����+s2L�ۦ.R����*��i�U0�j�<A�J�T|�riXz��� ���k�w;�9ڧ�]�'VM���I� �$�N�(�]@��R�F�!��5h���퉩�.� v����P��͑� ۚ��O��}�����W(������fĮ\[R4��6)t���ߕT�<��1�&RS����������'�OT����:>�܌*a�ܱ<�P`I�"OJ<8ca�;_*��baU��Th"O�)�*C+Y��
b�z��@��"OV���Qk��˚@��yh"O&�9�$K$j�T�Āիb�hQ�"O�8x1�99-�u1��؋
܂K"O`��c�S�i�*�T�̠X�ڕ"O���N��0�{�T�Ʀ���"O�<BP����Z�x�-�!���F"O�2��<	� I�C�Z���z�"O�������3g�y����*ph���"O`|�1��@���Ax��g"O��J# ��X�"(�nE)%�Z��"O�,yc�P>���hP�&[���Qr*O <Jɼ]�����#e>�*�'��H�	;g0��v@Ȇf�8�'�y��L
F�0agj	�^7����'��ؑ'扈%�������Xu�ȓq.
�q,[�z��m)7�M�q@�ȓ8��Yc���J������W'��|���j�&KĎ��E
�K*
���d��Y��$npz����f��ȓG>�<��gԬu�<y��(�>3"A�ȓY�v�1+&%��<
@��G��	��O#��s�[?Q�*��ʐ�B5��Y������U	�YSa�ZN�-�ȓW�$�I�h�3@gn=� 8A	��ȓp�����z��u��5՘��3%F���Y'> ����,�,Ʌȓm�d\ا�C
/� � ��%g���ȓ(�,;p@G:R�tdX��ܥQ�x������[���dݣS�5��ҁ
��1*�>Jg!�$��fjE(�'��3�\�2��\�]���oӺ�*֩�R���C`�'M�Bq�'"O� ����ޒ_uH)�g��:ɼ1i$"O��S�T6t
� � �� �ؕ�%"O�}�1���-�F�zr�&dF. I�"O�L�h�&U��xx�T�:޸�S"O��2�ţ5u(H�f��q�x@�"O�9���o^�)��ƴv�~�0D"O��+vJ̺��h��kÝS���A"O���РJ�>Ѵ1q��H#+n���"O���.�Y���pI
6a� d`%"O�$��L-��5��!#�,A��"O���� gw�AsP�2H- �"O���ǟl�|�j��U�E����"O((B��
Ok8�{�$�'mY��"O쥁�°\���@B�3��F"O �����$��bP�Q�Z[ʹ�!"O����`Ǜ�$���
ե%�U�A"O��W�+.�L AȜ"1t�S@"O��I0eޭ� }{�"��U����g�]����bn)m�nT  ��q�X��E��y�(��c�����i��l�(��B�׈�yB��X| %�p�ӟ`�vP����y���6*��d`D�"u-l�y2�ڿ�y����\�\A`gk��y�ܡ�Ñ�y��i�l���bӷO-�(i���y�fƽ?����f�;���Zg�\(�yrC§K�b@N�+*�N�B&�P��y�h��P�.��Q��(I}v9��W��y�,[�y��`E�9C�Ѣ�ߒ�y".ç(݌ib��S\P�b�ȟ1�y�"�"0B�c���BZ�Js�>�yb�&�8	�D[7�R ���yr�l��ؐ�&]����#��2�yb�T��.P`��	;qD2')���ybH��r�C��P�n��&L٩�y�&D�$�HH�e	�O�<�SN�y�/��e~�Iz�(��8�(���B=�y�˘C��x�t B%o�^�	����y����__޸)W�X)>DQ`����y"�Y�4���D�:,Ҹ�@�M]
�y�	Ȍ�N�e+4R�Y
Rf���y�n�Pr�T�bh�,Z��X��y�ԫ'�J�z#��6Q����f��
�y�B���a��A�M`��r�gߋ�y�L]�,�D	��Ɗ@�H���Ӝ�y�O)^�a��匩*ݨq/�5�yR
R	�~\0�+F<{�q�0h��y2�*6��L�6Ϊz��I0(@��y�m�/(��йo�|9�IC��y����>�x	��G�X|d��#��y�W�0�B8�F`׷=XZ�L��y�QvT��@P������1�M��y2�U�\(�f� 
��ƽ�y2lBi*��ٷdX(�����K�y���-�|i�J�p����GH���y2m��@��!�^5E\(m�ꏢ�y$Ӳ� ,I���=G�>ف6�ЯRN,�@����T�'-RЛ4�
�>hЍR��R�b�x�)�'ZT�E�Y�v^��l�]�,��'+h\q���>#�@�f�2�����'��Ja���!�`��2� 
x�H�	�'��5N�&J ���E[w�(D��'�����_�'[�̪ѢVn'$��
�'r��! ���}�kp�.^��X��'<@�����8eL4�Ɛ{��� � ��� "Hj��iR��<��3"O�xK�J�(��u��M 	�g"O��:2 ڻ����ꝫ&�:%��"Oj8fG�R1	�P�^��"O�)��	}�d�#u 
"��AE"O^L�fd�#C��Bu�(?��A��"O��[� �?R r%��h���"OLX��A��:Ï�;[(��d"O���3ɐ7#�|�	�=�<pC"O�=�pʞ9Q���#*�.f�F1A�"OLL��=j�s�BƐvU2Yqs"OD "�o� ��ŉ3=��R"O�h:a��?�0���(�6"q�a"Obq��땴%KP�h��5!��iv"OJY9�,�2o�:	93�� 
p�4ٳ"O>T��7sޘ��W0�P�"OD�SI�y��`��]%<+6�##"O2YT��U0HكFgzݒ�"O� �!��#bx���+��,�h��"O\а��I%r(�@�d$�F��1d"O����D�;N�,���1� uC�"OtP�H�:�x"�e�Z��"O�T* ޙ"="I�Deϻ9�&���"O��D���R�v;`E���"!"O�X8��ĉHrg_�H�i�"O����0�Y� �ި��4z�"On<y�
�_k�$!r��� �	�qɈ�b�c�f���]Wk�ݐ��B
z�l�hZ��D�<�R�1ahC� S���(��uyn�G{b��Y��x��vɲ�b����'�Ȱ�j��^�x��%����R�yb��ւ�ʰ/\�JQM^�����e%�L{�}Z�ğx`�r�
�$K���[�̏'X�`�v�|�'����q�2�����g���"�Ԇ~��C�I&o��e(��]�W~�-�_���Q�IQ�'U2A�&�O�񑁥_�ZΊy��4
��%0 n�9Z�Z��Q�4Fx"����>XIdH� *�r�X�
�#�����q�ִ�4��,@��
V��(I�Q���p���1Pֵ�0�� t�R��<qF⒟k^ ���X*��Ê='�.���� ����a�ҿ)����C>i����b�K�X9&�sG����&e���q�#ׄ?n�]ඨ���O ��oHjQ�$h�a�G���C �Px�H��=�@�@���ApEZY.��see,O L�6�5)�d�XZIa�`@#_ J�'S�4����_�`�<PC�m�n�*��`b.mp�ר�0��?�?[���Q��g@�]��(PO��,F?�0���G�4ݻ�*Su����n�_`�	PA҃��a��>y���u^E��b�:L(L�J!�ۗW;ޜSS�E+�V����ԋT���?�1^��q�m�+�~��&��e����Q�DՒ���?�'����4�K�8y�Ahȍ[�,�@F^^�p�i`�'��#|U`'5z05�b˙ )/2����T���pP��'��ʔJ��R9r,)� #A�s_"8f�֔L�0���ǳ���O���ػ1-�e8��D�2FR���r�1�:I0el�E�I&�L���$��C�01�NG�D],p���R�E�>�쐺G�ƭ
��J+@@��ݟTr�&�Z��F�-�HܣT�>���TP&;t�V1l��[�����D#�&9p�4�l��נ;�	�\������"Ǚ�/�����f�E�����Ǧ9Q�͆�8Z��� �3=\��M>�/���g�2l�zyqCE=vL����;�	9"�Z]���(��D��@J-rÄ0���� )�Y�(��Մ�I{�21i��輻 �ҽgx�<�ƃLBsDM��FM\�	y?��N]�K�(�y�o�|1�����KζWʔ1��L&`����?�	�=���i���-���+g,ùL���'����^�$
ޭ��*P�+��L�#�<y��'12-�~D��K2�M��"@�kx��0��T���AZ%��`n���$h	��^%=^ţQ���Of�SF2�;����?��P���%R�̱@1�i�`�B�oRj�Q��43�P�80�ɺ0�3��̍�F�C�Ǹm�.�	��Iv?�K�֘fV}�7�[�<�а�9�,�ci�'�p<Y J��䥰�w%`Y�&���[( �
���v= L<��'i���ҫ4;(�B9_��q����P�!8��H�?! �=I�9C�f5o��0fL�dƱMQ�ɺ�b,�����B�F�f�'Db�'�:�!Zw��G�U���\*�O�hU�]�`o^L����I�\�q�����4
���[+X@�P��9��Ok� H�" ���(�q�G\�}���v�i����{���i�oJ�^S�����4XB�C,[r�p( �(GA��s��,�Z���O�q��5�Me�nik���-;��	��N�Q\��R��&O�݈#�CM�D�ݜU�C��33y��� �	4�SAU 4�6-��`�dH�|�.�`��Q�Ԅ!U��O�rQH3>en�̂ѧ4�I����G��2r䠔n8<J��'��=�1�B�VR��B�fPh����>s�h'd+��I�H8�<�7�Z�6� �A�jH(��a"H; �!0t~�`'��(1��"���C�@ G�G/6®����O?�.���Ha`$�"�@��X)R��aN��m���J�^�\��#U*���B�0�4�ʄ�7CA�&8t��n��f�l)Cw�<�d��F��)Bu�T�Xs�?�XNBpCe���y�c��"n�T� L�p<yV��;����w�2����]A����E��}5���(�	,:X5��l}�U~��H�~����y�d2��\,aюx���ˆ.F�2����O��Z'h@�B��I��M�\��a�>�DA�z/Z�*�㒺=;�xm51�D�������ڱgN�-�"��h5޵aS�i*v�P�	|�LEà��9�<`�����@�c�DLZJ����+��Xӕ�dyb�^o�.(�aI_Ί�Yc2�I�#��@��Q���,0��(�$�*�	8�`��O�·�
q$�����#P}�"��<�~��'}����$a�������8��ӷi��	Σo�,��GM�'�|���W<}S�=���BH؞���g��|���y�p4�E�nJ�)K�jAh�Z@�`�gCڔ꤀�O����M4N��O�V,kj�� �5�lsgCY�*I ��$�M���S/O�%$�O�R �lZ���i* �ą<- y�8t�&e9�	��"��\��F	�7`j�A�`B�cph)&�ܵ\�z��>)c���%�����*A�X�+�ėX�'>ĕ�A�۲	���w�!�Tj�GT);D<�x�"M/L�
�aU�G:��(�t�N�������>�~��u�����{��$�b���E��\��+qM�-/ݛFJ��:޼�Ж�ã"�.H��C�Q�D	��ɛڟ<+Rꊤ޺�_w%�0�M��9 �8tc��S��=�U��a[����eZQ �烔>���᪉�ڪ�Sr�%}��E3Q���:^,8��vv�1��ͪY���Fx2G2��Y(t�9fm�Ia�����$J�-�*b�d�/N�<�'��3���W���q�fE˰�G�#̜-���ٻgyD��'��A�6�$.�^��k�t�t��W�/�~I�� ;�(B�B�k�9{O2ē�Mҋrx$,	�l�%�J�h��i��HxU��e���:��G�V�e���ą�#0~A�HF#=��ł�A�V\�:�y��)��j�3i|F���X��rt�[�J���D
��p<T'W�d�(�w�$@�H��(��ܠs/	�hhN\��tQН���$�^�r5�F�����-�'yZn��0�D�1�漸�bL�V�$)1�/Kr���V��+YCᑊFǼ�Ez��ݪAti)�5O�����@U���$ָE��A�G#M�R�@���
Pb�Y� �:t����H�[�TX%��j(O�Q�.^%%�,R�� +���I�`0mڋ$ �ݒAA6$E^��$�,f�(#?!��˖#�X�wIY�:�ȑra�r(�'����O4e�vI������ �@�7J�Ӑ�u.�xB
#)��*�F�︹[r�ܚd��i��mI�2�V�(�ɕ�eGp�i>mI�Ā�w\�6�Y�ɬ
�V�V14t�ċw�OxP f�~!p�'���"��?˓$T����*�):�*d	�([�N�:<*�OL���'�:���5xv�H���u� �:�&q�"Q�f:�A���J��ac��Ky�J����O.H:�����~Ba@�?7튃��Mp�.�;� I����>qۛV�ÝI.�q#k$	��t�#f�5��O�U���E�+T�:��$tg��BS�'IX%�F�Ϧ����:���@џ��;D	J�a~p��G߶H��	�F,Ϝ��
�=["��#@
�|�"	�*uTFP����/�ڤX)��t`�PCm8���F�j]�,b������@Ơ�/iԅ[���n���8!ץ�=\��Щ��I:UL$��P��\����e��"=)�/�
f�Ń��?��Pp�R}�A3 ۦ4+��R�p�tԻ1��>M�5�eZ�Rl.">����:�&��' <X3�
QID<j'�W%Z1�M��4+f<U%"��m���@#V�	 yF~�NÖ9R��r��/fJ�LBT"���'�
g�QM�Q��� ��AaR̓���(h����.�?ORPx�P�Xe�M�o��JM�s,
y��S�� �h����E��~G�y���(R���-�2�j��,Dr����HH��@r���dR��ɧg�엎Z%��2J�e���$�I=M�><�`�t�(����(��,�秮>�'o�6U�%*�������S��˚?r�hQ��@��ē�M��O�V�C6>��q��i&���%R�(��D�Y@[��"�'�@X !�҈T���-AF{C37��]ض"_�a�ޝ�&MY��?qwaϥm����-R�ԹďSS��'#�	62����$�^�ɖ^,d��a!�h=�p<y�.K&8���qިH8�bT,QB }X�ψ�#���i'X��!Bx����'�$�� ��Θ�c����MX#l�(X�^$k�@�]Z��h�G?�ə_M�陴N�<���NΓQ@L�����/3��9��?��O|���'��=b��0S���c�?N������dE�+���T68_�t#b�.0Ve�6[�P��1shHt��g?��7�~���5V��h�^q���$.*@q��%@uP؊R��
)>��.�%RU5�S�? �]���Xz�E�ЦO�N���G�ε���#4O�u� ��>�3�H�N|��뗖V1��Wf�W�X�P�ԇ>�x�GL�u�\�f=O�b�� d֠I ���\����V�O�!�E"�A@��c��rT�	h��U�s�p�p-޲\��ӷ �UϘ�`��	�&gj0�d�J�%9
 �gQ@��'cQY�q( !91��2q�⟀oZ<s�DK`�ցp ��z���+0H�m򄝠� ��[��q���T����"G�)
�����'-�N��Ua@��{����hR�@�vy��Rn�EC�4�ܜp �/`X��%N�(hb�G~B�^1~q AC�d"@R�����@���T�  �y�'��jra�h f��-�3l��8���сf�&��ɖ<N�� ��ڼ[Q��>+�0��B�H5,���c�p~���O�����Xl��dڐUe.�Ui��b[�e���O/w%�(� ��J�e���X��
E����ٿnJI���@��cҍ"Mh�Xu�^+ܩ���$ɘ'�ܨ���O�&�*֌����Ywj�ɕMh�XKp�^�,�X�%P�6�\ۀ���D������O���+e�<泟��'�lQ����f!�w�,l��%j�0y���(���xC�ҶA�l"?�D��q�p�+�'@i�8Rd̙�D�f*6.TbD�  2
�81����.^B͉c+>�a8�>Rڈ��q(ļ��?�0�:2��\3��ŅE"nXY֭�S�<�uG˯&p� �hL��D�R�<a� s�X�*@RY�x���K�H�<Q��[�Zm2��҅�P�!EE�<�t��<�4X�R�6�$��D�<)��pt���KJg�.����F�<Q7�# h�kPBD����ܖkV�C�I.L�8�֫Ac���Tʎ&�C䉕	�ՙ��_�?Z��A���� E�B�>��pjH��a��]�F�=
�C��f�͸5�~�L		a��	D�B�ɣJ���zB/Q4Yfm��Tz�B�x)�<uM�}l4���H�B��0&?V�B>q����m�8�B�I�Z�(j��K�#1�8��
4��B�ɁB��7 �/ma�L
eK	tfC�	?w���e�$��w*L�hzB�I�j p�
7&L�[�T`���Sn>C��66!���՚*������,"\C�I9'��m�0�(���Q���B���ؘY�&C�'-�Zffqm C�ɅZ[@]Р�.��,�<��B�	�(��GD��<��0¦d��t�B�Ɍ>�i�$�þA�b�A��R��B�I�'�q�5��Ü� �۶>.�C�`Bȩ��]�"1��{�eZ.^~C�ɧ Tj���|��%�jC�	��!�@J^�G�lӒ���IfC�2q���v�T*C)���A&F��B�ɳS��`��S�]y4����ގ0P�B�I<C4�"��O�(}A�e��D��B�5UV����T"s�m���	Ha�B�	�:n�	��ԷG�$��N��B䉼_qr��ś-� ��G�Y�:��B�I(!iH̀P� ���Ӡ��z�B�I�=�5�tB�I7����qQ�B�	5NE��e�"�D��Ü�e@�B䉪Q��a�`���X�]�l[���C�I
a ��qa!i��)��5K��C�	@��!3tk�+c��H�Ɩ�Q`|C�I�~��)#V�2[`�`-��B�	�F�ӕ��.z>�b��E�vB䉵E[&�)E��+O��s&�;RhRB䉄e��Dѧ�]������߉/ZC�	L�	*է>mNhqWJ�Bu.C�I��P���mY:�>ᚥ,A�h1nB�I�U��Lq�A|P�CDɉ�o�<B�I�/�  ��"MNFq��o�07�B�)� �L"$U��B�Z�15tD:�"O�L��F8�d�{�f��n��P*OFm �.W�&�Z���A�VO�!�
�'�� X�bP7Z�Idܯv!*�
�'���%L�K�'��{�r�	�'k�@0!Y<n�I��U�t.�5I	�'h���a��.~�ڢ(Z�!ļ��'�D���B�� �j}�U G� ����'kx����͏w�,��	V��ͨ�'��0�#IK����ɀ)X3�z}��'����1��<[~FD	$��T���'8�qPӤДl*Y
�X{����
�'#��і�^?>�P��ּv�8C	�'��(��o�h[̘0�ݛtG.���'�)�lO')�z��#�[7mt�`��'S,��ڥG8�e;�%ʆ�A�' �C��ơ�>�ӵ� ��D1�'�p� j��3Y�<��&D�~����'��L�P�k�S�aǘ���'ئ��"�=� QB�fHD�b�'�@��@t��Q���:���'ᒔ2c��d��0�
|�d�y�'��X�qb܍6a*���K�np�\�	�'8
t�(XŮ��ǩ�ix$��'��`��-R0w��x�,��H�88�'~$IP.�a��@���Y�+����'|��F�+n���ǩ32.���'	!��+�9T��$� B�j�B@��N� �1b�s�@A�	֕#z�ȓB���i�O�FH��*��2�(P��+P�]��a� ^�����C�����ȓcrX�OM�i*)�U&�6��-�ȓN�F��C�Y�.\��qB�M!��9�ȓU�@<@FNڭ1q���&��10
���\/��hsυ*1v�D�$莾ned%��]>�I�A�:!P(i�j�IWbx��R��pK�c�n38$96g��/�޵�ȓ^@���e�� �  ɿ~虆ȓh�JAg��f8꼰�j��jẍ́ȓw\�:�X,3n`XL-8lh�ȓ�ZLF�Al�h����*p4�ȓ7�LĐ�"҃^��y��'5;p���G*T-:5�lE���L�e��X��T�v�_�d`�L�7�^Ʉ�[��Ac]�o���q@�@�zTH�ȓ>Bޕr��o3X���(H�N��ȓS�$�K�T8 d)!ͽp�Y�ȓ)w��rU.Ĵe�|�i2�P:��=���lK�!��|ѱ͙�:�<؆ȓq�h�#ݲE5ޠ�&�P&<��#��|)%+ںe��qс�.B\C剔`�:4Bb�hT� .I�8B�	4���#��7�4��͛6Q��C�I�LBӀ1?(`  6 {�C�-P{
�0�'#��)�'C�s��C�I"}w`r��f��	,P;S�dC�I�1]tH�q"H�-�������tH.C䉧p��Q"F�3)�M� � [� C�ɱ!'t0C2�W�{I�s��O:C�I�_&�!F$�93��� ��^���C�I�a�\�pf�4~�8��x��C䉀r�*ũ���<:��0;!n�km�C�I0]iBʣK��uL�pBQ��:�xB䉧V�����kW�^��I�wi��KGZB�)� ��1�G�P�8�s���+uA�"O��!҅c�A"5d�*H �]��"Oj�Y�!q�n0�"#_/~nZ��B"Oz(n��\�)��F�eL�Yq"O8̂���D�^,;�J)6�ZTr�"O�a)��O�z��!�����ޢ� q"O̤���,��s G�J��"O�ԙ0�ՂA�Ty�%�x��P�"O.@Kd�]�솀�W�3S܆�"OX����I""���7�Y�;��<�"O��Kr'������[�RԳ�"O`�#!���y�t�-w�(}�"Oup!oc�B�Lr��hg"O�)��_�Ԣ�c��#w��P0V"Or�K���'���m�)3��,@?D�Ѳm�z!� �r).����F�>D�D�b._�q�mqaM+x���1�0D�0����h�yoJ�^�l�$O#D���U�
����҂U˨�q#?D��caIIʲy��jN�k����F<D�$��`J�>*����ᙷ�b�Z��9D���W�O�}5D1�4�҈ma����u� E{��i^*[�:F�-_���g�E#!�ď_<�	̊&���K�N!�D��̰vNʳ�:��⨖6
A!��&L䤝�FbZ�J�#��1!�d�>����2���1 ��r��!�D0w|�Fa�z���6�K�Xx!���*n�H�C��:��P��.v!�d�a�0�墔���(W�W�FC䉀4
��ibC��h���厃�0�C�	,m��JB�P6y�(���(:PC��IM�����a�Q�FjC�	�I�B�G�O�#���a�\5"�HC�I�,l�=��7?p@P ��%f,C�	�K��Պ���E9ȴ�dխr�C�I�"@ �K�"ͼ��Ð(F��B��.&o���%�	�I��@��H
7aj�B�I�n7�4�����cr�(�$��fȾB�ɴ�Cd�B�c lhHvBL�$�B��!Ӧp[b�,G�2��� AW,C�I�7�T1�c���8d��|.fB�I6@��d�ƨ���4j�  :x:B�	�$B<D�Ճ׫a�"� ���
B�Ie��ke��[Z4�
W��T��C䉸O�2y�� da���AP9U�B��7��b��S(x��HLY��B�Ig�F9�Ջ�2�|�*G�#ǎB�ɇd�&P2�cA6K�i���Ŧ�bB�	t�6� �,5{�i9�
%7� C��X��L�2�@�~����f�.B�	�<��tti�,WL��֡�d,�C��9F*�YtǪ
Jl`n��j�,C�Ie4P�����NE�]P��/[��C��d�`����D��m��C=-��C�IT�qAPf;8�JJ�><i�C��B����L<�j�P�bvpB��N7�cw�I�P&Y@��� n2B䉩o�!��K�sqFu �Bg��B�I�i�m�r蠃2cE6O�C�I9���Êe�H�0`Čw� C䉴Rn��^�Z��v�C�oh�B�	*6���aF���(@��.x�B�IO?T�A�Xd����DܲA�\B�)� ve �W�:q\���(�c����"O�$B,�̱;�I�n��L
�'��z���#-���Tn^�]U�a��'�|t��F={�D�Q�Z���'"�f��3L�q!�
WN]`h��'A��;�	ʛ9]��*w(]�z�2)1�'�BdRcjF�6N�6m�o��j�'O�9������@R�%k�N��'r�� ���bd�Q5����'��E�dKK�C� �sK� M���S�'X�2C�N�J��cj��J;<��'�|��V����2	�dHK#�yF��,�<���!ݎ+�%��c�/�y2Aڵ$�*�C�&o"���E\��y�+��M�Q��T)=*�2�����ȓ�� ��EiB�)�I��GHD��G��u�u�=v*�ybR7<�b���;�vp��I,ktԘ҈O3�.i��J�,L�$,�X��ax�N��np�ͅȓ;jj	jC��1$����S�7\Nu�ȓ:t����@J���'�@��� ��{(� �d�X(��Eݟs�,���F���w�����yw������ȓf&2����C�k'v=C�!˨w�@���
���E_��c )ƦA�<(�ȓhQХ��^{X���'e^�brчȓ?l �c�C-��R�#�h�����A��� w�L�sn�a>���ȓig���; �R5e�p�Յ�k4���&�P�QZ ��@D��m䀱����6�@�w��f�^ل�2fݓBB�D|0ɠ���;j*@H�ȓtΪ��@��H�Ƞ� `��d�ȓڪ�S`&V�F����װba�a�ȓbӂ�� ��n���͛0<����V\l��á_�0�H�ۖ(�2P�(�ȓsx�GԪ;
`��O�ks(t�ȓFFu����u���;H�U*`���`�.4�D�j��x����J����m/Le˓/�9)j���C��a/jC�4P���H�w2
��aC�6(C�	�n�Q! U�#:�ADoև9C�	�W$DrLM�:�S�cV�B�	�U�jipL
K�����E�o��B�I���HJ�[�U�@�s2D�+H�B�ɸ�rHW,��Cch�#F�%�B�I:B�f!R�e�UI����G�ef�B�D�pb� 6D��dK�	31�C�I7j+f@�c�P��4A�"J�B�	nܺi5�,:���* �B䉝�&0uK-�J8��Z30dB�ɶg�-�����nP�`X��Է!XBB�	�R,�Q�8���7�vC�ɎC��7M���<�x���R�C�.(�|�2�ݔ����m��x��B��L���1�hE
6��|xq	Z�4�B��2r���P��A�X!�v�Q3�B�����$��(l
�G����B�	�w��	1$���,��d���F'�B�I4-ʂ���JZҜr4$I�&'�B�	�xt�	���'}�D�gd�/Y��B�	���P�Q��o�Ȅi��U4v�^C��{�N\�d�-S�|kÅr׍�y�#1� �7[a�Y������y
� �=�g�[���B��4p=Jq�"O�}�c ����d�\?*<Ԍ�"O:�`����`��/C6�c�"O�)�!�!I�P�rd�p`"��"O
蘶"�VB��yT� �BX$$
�"O��`q�D2xT�*�ǜ,RKl�j�"O �0�!S��i92DX5>��&"Of��&Q� z���ʫM�n��c"O� s6�W�:D�B`b�'2��5{F"O|(�W��3����cBz��#*O���w��v}b̛!�ݝ+� (�'y�d� �7�~����m�����'x^D@��#4ָ]Zqg�#p�d �'k�݋�&��iE��wf�)klؑz�'4��Q��
6�����ޱeMp}	�''8E��T�zb�Q�/E�M~tB�'�޼�%��;ƞ�óΎ�L���`�'��Q�-:E��D�rOW��h�'����7 �$��	��9�T��'�%-L�\CҜ��:#��>�y��:{0��8����e���y�A�F����7�R�~O�����yR��D &�х�7s9����&�
�y�Dd�Խ�$J�8}\��ş��y��T�a�t�� �B9o�P�P$�y�6>a�I�ˉm�`!j���y����T�5A��dQ��B�΄�y��A�������W�U�5R����y�AU�r�0U��M�|hrς:�y�KݭG�d�ɴ��	t�� �ٽ�y�ΖPkq�.�}s����PyB�
++�xj�ɲp�쉗�E�<aWHW��*��#�v��؁�/TA�<��)3P*�Y q8�H�J_C�<q�h�$��s#BS�Q��e3�~�<���]�$n�`ӄN��_0}�6��w�<aq'*�6� g��(�Đo�<yte�?0<�@E?F��(B�`�<�ck�.0n%c��V�Z%P �Vd�<I�n"B��Q�pF?V�hT��.d�<����'{6]Ѓ��"m�i��_�<�a˙q	H�ã�J�O�+��[�<�B"P�d�q��O��2�	�X�<Q�H�1� lꗧ�)9�l
�B�\�<Y��"p%2PB�NQ4V�9�@U�<���L!��S`��=U�Q�EK�<QCJۆx�n�w�T�z����H�<Yс�/5q�x�@Ekel�f�AF�<�V�Y7�v�� �K8@����}�<�vK� d��p8&M�2s�$J7$�v�<Y�@�2v@��j�R�1br���fyB�)ʧ!�"�h� ;Cxdk�d�Ij��8��m�� D#��S�,_
:�%�p��	).�N���޼-�U
G 	����)?� <��2��["$qvM�6��s�<�G��/x4� d�)�ȁjUD�<A����nǎŃ�K@l� �v�<��A���[G�`�xs�s�<ႆƝA�\���Ń:���äE�<�q�N�.�H���<�T�����<Yrb�	u�*1�յYǤ�2Ƀ�<) 
W�a:�R�`�
B�>� ��a�<�E6eJ��-G�Lq����x�' ў�'a��Ru�K��̈�åA�J�J���S�? }b#�V�
E��E�}�B��"Or,qq�܃���z�n��zH "O>,r�c�?�:-!�gڅ!�,G"O�Qs�57{l0��N�u�j�!e�04�+�Ñ�/G�IB�l�r5�W�7D�����O��@+�$H�RE���2D�$�fY�S�^PшK5O�dp�
0D�����Ft� �%����e/D�|�H�Z�\����aܦ�0/"D��2�
+e>0�d��9�`���4D�,)�����ݓQ�H���k5D�T˲�@�0�`����.b�\؛�ct������/+j ��۵_D��f-A,!�C�I+�PL�c@Ew��O89�B�	 mJR�J�ˌ�d�je�s�۷T�C�ɗ#��-���G�X
)��C�9W��t���!(��)��Q�6�C�ɛ6¶-ۂ�@=
���c���cШC�I�7����E�	M�=�fZPn\C�:1�L3���r%�a�<o>C�	�k��4��!�5"C�{7��g�NB�I _����F�"2԰�+�>:�HB�	��iŎ�ec��5e�:�zB�I�|yH���7+��Їi�>\�|B䉙��0C����S\�U`"�X��0C�I�|iAw�^�=����.X~""C�	�8mT᱑ͅ�zC����-U_�C�	J|Yg��c
z	��E�=��=�Ó&�� h��� &�е�qjچL��P��R�Fɡ�E��<9�ŧ?w�JH����?a��ۙ&��9x@I�6T/ȵ�c{�'/ў�;��p�٤1�.�K!�?�J��~�0|��T�t�J0�үEV�ȓҘUB���>oq��e��-G�1�ȓx*�PV��(��N�b����!�|!�ăL�g���o��lN�l���L�B@�8C�/B�$�P�/L�fv�}�ȓ.Bhɗ��'8�`�*�4Ϻ���R�`��1�/�)F��2��Z(yC� �ȓ9+�\*Q��ve�j�IL<Z���'�ў"}�4g
�PN���5?%X��SU�A�<!b$��[�9��e;��9�Ǒr�<�A l�R8#�?H�9�4m�C�<��ùk����תQ�z"*X�&+�X?9����0��埩,�p���P��ލ�ȓ��dS㏙9x�j��P��kȭ��7�p�H�(9lSz5"5O&N�V5��EɺQ(��,K��Y�Y��1�ȓ+���
�`�#a[*Y�C˅V����J'�0�@���"�:�ʇ�_( [(Ʉ�,��PȆC
�Z�rc�	G4|��ȓ:��Vm�(�a�I]�4��ȓ&1���c�.�u��#�e��%��
�
�z��ً$dQ��E�8( <Y��$U"�h1jD?yʄ��n�=�Ʊ��h�v0��&N൛2.��qG$���u"@ ��;L�ا���{�.$����<��2�)y%��"Qჳ�C}���0=!���T�͐�o�:�,B"�Mb�<!eM��@�+�M��"�)Xd�[�<I�bQ0>�)�����P��mU쓇p=i1H��֝0���=������R�<���*%�QnF"����@K�<��̸��9�5@ E�S4��F�<� �t�D�
wt�ۃ�M�j�"�p�"O"�2�)ϯ"�.���Ō�D�x` Q"ONm��cԖZ�0}���`xZ�!"Oޡ`�S�ێ�7g��4Y��ɲ"O��
�h�?~w��y���YV�`�"O	I`U$C4p�4+ζ	XJmA�|��)�S�eV.���nX<D1�co�3�
B��# ��=���
 )��0Q-��f\�B�I�:��� ��s�)Ќ�I��C�I2�@$1��F�A�����R3J��C�ə,7ZЁ1H1S����d�Q�%7�C�	����B�&��!�̴0���QzB�ɓ���[�Eқz���_�M�LB�ɺ`�t��ڧV���†_�d�B��<Z���c��òtQZF���~m*B�ɚj�l��tĂ?m`�YT�QX�B�	��T<9��ۄLaxi��\�aɆB�)i(ź�'\�	d9��螴YI�C�ɤ3���b��/�DÛU��C�		)��Q��^�Y�ҽP��߅0D�@CDf�9`Je���>	�x�s�/D�dВ�72dQx�$��N�&�Q�l-D��م�R�p��5�2Ύ1c��!k'F)D�|kuH�N�\E� ��6u^x3�A<D����P�@�XȐ�A[= � �'D���*�YԘܒ�JI!jx��%D���7��0Ĉס�90,��s�#D����,��;�����+Puxx�%!D� [ *ԃe��� J�
G���Z�	 D�L��`�J�������Y�FL=D�p�r+��s<�pWet[�Yҕ=D���3��#<\��'����.D�P"�J�*&��e��i�>Gp$�!En,D�����Lvl;�	�/ ��]�(+D��0��`�����/k�<���*D�|� Ô�M�xBBC�%�L�d�-D��B�	 �32��3uべN�j��+D�\I���1H�*��5O�4�*��g�+D��� '"� �9榐Fy��:�e>D��8�hW	!q���F�O'�pQ2X�!�$�,��� r��:plt�r+	��!����`�P�;���XQ�t��!�$ǐ}DB(AGk\�1A�»�!�$˷#P4�dʀ�J��)�Q'Y�%�!�$��nH@ɔ��<)�F��u��"2�!��Ճ+�܁���*���9�A�k#!���,A�zP�W���n�����B!��H'g'� �Ü>�ڐ0'���Py�O��g�\��Q�=��|S"E_�y�D�9\�����.�mȆM�y��a���QiZ� 
!r��U3�y���9���Љb�b3�E��y�$i��:C��	�`}�S���y
O9kŶ�k����|hZ/Ǧ�y��7���q�+��]�x�S0LZ"�y�8uA>�[p'XT��!`���yR�C/�LYQD$�RM��� �:�y¦�>Z���0��G����P�y��ةU�rQHt��#8'>�r�i�y�$ص!� �{7��;9�hS�.�y�G�q����ӆ�9���B�a[��yb��)��ܓ�e�hB&�k����yB�͋{�j4�rkG�b��MS�c�;�yb(�!"�ԩ3�� 'X���g��y
� d�+�H�(��0���өAڠ��"O���g僔��D�eÓ�g�@-ɢ"O��8���
		��X�O��N�~I��"O�5rU��[��1����&�R�G"O>
W�ȃ4p��gȑC�
u��"O�I���*<;|A9�fπ>�(�"O�|a�K˳�p�Q��xp(T"O�uX��[m21�`#]%uni�"O��z�DR�T"��(����$?8t�A"O�HYІN *�L-{$*C"Z��� '"OlUk!�^-��kb�uѤ�z�"O��B���>�4��6��j*�(��"O�8S�
A��t�7.<0��8JC"O��	�K�S�f=��)%��b�"O��!ܕc��Mp���T��|�""Oށ��Z��
�q��+f�(�"O�P"�#X�{2Q�6�;�� d"OPѹN��֑:kɍ#MQ!"O���X4�Jy�u  ��h0"O��1Ĩ͹|��겯	6a��,��"O�r4CũbR��;�OV)'��	�r"O4����(N �roI�x���"O4ܪ�*�	vА���-�5�,@�"O����)]��ht
��F�b�DI(a"O��O�^�"Y�h(>\�X�t"O�`+c�(RV!����$@ 5"OF��փ[���`�'B�`���@"O��"�ֵ`[L�P�Ő��B"O�SdH�"�(�#EÊE��""O�H��7>ޭ���.���I�"Oh\Cpc^�N>EA���R�b��!"O��Y0OB �ʔ��]J1���"O�H�t쁉I��C�m��>9$BU"O�i6��=^R���L����� "OdL+S�^�Py1�xZ�a"O@�ao&�@����?ys�l��"O
�q��&$6HH�@ڄS��{�"OĤ�So���)�EӈWؼ�`"O��rዷ�"I&D]7k��px�"O>c�
A�O�̨6�	�|ºt��"OZ�ȗ���v� �td��%`��Y�"O�;ǂֳ=��l���R7vUx"OJћc��#8[��cnN�%$�4[�"O�Qhu�M,q��;�ƭu��A�"O T���l  �@������'"O ��Ѣ��w݊)�M������"O�S`I��>�4;1�8o�8k"O�I��ܜk%x����@Fz�"O��1��R���j����"OF��㯓�'��i���7!��}C"O�!;�C�E���0��a��q�<��*�TV`�W� {�$�P(m�<�F�ǻ(�Rܙ*�u�R��� k�<�A1h� )"� H�]X� ���]�<!s��hR08�K�/?�
Ј��Rq�<� ��?Q�2FID���M���j�<)A� ]_Hu���Ȧ"hz�Mg�<��E[�a�s�!C�du;� Yf�<рW�� "�߅"`{Ć�l�<�s	�o��0��W��c�m�j�<��F�z߄�Jb.^�[)��*� Wg�<����<XK0}����`�g�<i��C��b-I���==�P��n�d�<���#D���p'"�?|�`%X_�<� 8ɡ6iK�s[5�BNV�i;XxJ�"O�$;�l��54t	U $��"O�L�k��n�}"����4U�"O�Y�TK�LM\8���B�t� R"O�ȳ	&6� Y��#��hR�zn!�$м�q�ƍ�,�T��F��d!��нh�40cŖ0qt���WvF!�$�)rD�U	�e9��e�T�ܘ*!�$Oz���� �Z)�Ȱ���+ !��3� �Z�+�L�H�!U�!�DP�)jja���џ7j�	ؖn�l�!�$W�V��Q�X?.�p	PtͬG�!��W�V!֎�:m�� kRD�1W�!��2e��#�1(�����ڶ2�!��ۡU�@4ꐫr��cBX�!�ї|��{����z�8�`�`�f�!�D�?s��T��S!��ZB`�;�!�D��<D���ωn�@V�	�!�˛"甝c�D�'{��9�@�p�!��G7M8ZqB���jV�<q���.o!���;~s����ƃX�D��Ѝ�JA!��3Ks\,�efOd��]�d���@I!�0�6`� ◢�J�iw���}�!�$M"&~�����0���{�$r�!�d�^�,�V#�?R��L�D/._!�$H����W�f���Ѕ�D�!�!�D��'�D|(b��QL� ���z!���nDQ��JYS0���R�v�!�D�1݂\�"�٧!kn���jS/�!򤉩-�R}q�P�dN�$��	!��'!a�QQ���&@<h��*[ hf!�d��L-`��Y6�B����P!�� H�1xU���`�S�	��@/!�$ܦ=���e# �VX��zB�!�d�&�L�IQ	xPx���Q�!�R	+,~!�6�ΓO���b��G�\!�O�SsrE*@��3�����m�9�!�="���H$#!^�����aU��!�d�>F|d�+ ���xݚ��!߶�Py�BE�nK�5k���f��B�	T��y���xS\��e*J�I�X�����y��1d	�����=�(�@��;�yB�C�y@�H㔋Ǥ/��u Sd��yR��a��iwd��'~�A'Q3�y�[���ukŤ�Mv��FY��y�lHV��;�I���	���yB-�rS��2��\��H�� 4�y��ɝjf.x��g��>+�][G���y��؅;64���荟;GN�Ȗ����yN�'~��C�&G]0QVk��y2昙e�:p*�_?_����łC��y2I��e脱�2��`�иE@�*�yB��A�ͪ䏘>D(<�˧�D}�<���l"��˞pH����F�<Q�m�:�~�ZV�ۿ|���w���<	��3]Ⱦ� 3r�]I&��E�<��] ]+n�y�e��0��3�h�<��&R�_�����=/��4�\z�<q��ѫ:�d�U���N>ޅ��Jt�<yn=l&Z���J�5c2��n�<�b\A���x��^����@S�<F�[ �h� Ո�.'��m�/L�<���W2��A @�f���j�m�<a1@.C�P�D��f$˵�g�<� FE;e`�%R�a:r�-�Hۅ"O4����,8�����1a�J(CW"O� #�. ��h�?�*�s"O�S�W�c��bcΎ
�J(�v"O��RF�5$@p!���>����"O\<:�3�^����@>fC�S"O$r"Vgzt�
1��9_�$�j�"O�SԣG����Ƒ s��P�a"O6���J�[��,���o�����"O�{�&ԸK�i�@ĕ0�6-�4"OlAPb��K��!�C���l�>0pR"OZ�0R�L�#�fܲ3��l)��"O,�r��R�:��l���+�U�"O�%��A�6!ڀX��T3A�$���"O"��CjՂQ˴����F<9��#"O���G�^��$[��*8Y%"O�iW�G�,(S���~� ��"O"�`߈O&������νS"OĥIc�ފq�@L�RM=Z�r\;!"O� G�3X��XǩUw����Q"O�QAU/��D^`t"�H:$�<Ӵ"O8=�Pl��:Ҵ0+�A9����V"O�9Y�b܉W3������C@��"OR�Eo�*q����ֈ]B�i��"O�E�`Օ�]��Hc�0��"O���d��/qr��d&M�7ft<Q�"O����(�u9<���N�^�Q�"O�U�r	��z�bvOQ|�
�"Ot��p�(?b�����Ǯ3�2a"O PZ%KFmshQ�4���Sh͘"On����K}�q扚!^�Ԁ�"Oٙ�h���U8�.F�n(�w"O�`Bā����E��:�f]S�"OhثGH�M�����	]9F�v�"Of�2�B;7�Vak�m��&�<,["O�$	��̀P�H�!F��t�f���"O�����{�,{�@�lnp�"O�h��N�%V���S�x���"O�遥`F0EN�À�~elqp"O�����
�~�c솱5cpP(v"O�H��G�ky��%e��`HT�0B"O�<K�'�_��F �r��!"O4�H�a�6d�D��`�-��q"O�6f��LP�f���V s�"O&���m�3/�h� f�%�z��V"O�h���X;v���dм߼ `"OFa��π-�n�n·dȆ](�"O:t
�B$�pi�P�ԕ+�XC�"O*t��#_/��Q�2l\�Z�4q� "O�U�#`��ab��6+�i��0[�"O��
�5wk�}������ 5�7"Of@0%�W�ʩ)���!�%�"O>��j��9�����O�l��"O�)Z���7�����H%-��B�"O$\�D�YpfU 1㏱,:���"O�丰�C�bl��k@�}�j&"O���!�DY��1,ِdf�1"O�k儀:���s�\�M��w"O���m��E����ՍP2��8�"Oh��ł�5e�$�����+|(���"O��tl�W�$����ao�8*�"OZ�D�4)�=q�$_y�x9�"O�-�p���u		Ă�(!��\�<aCM�>0`�ET�6�{A�	Z�<� j%�P�<x�y #�i
B5�&"O��4唹�r):��Z-m��Ɇ"O��PJ9\,B�1�� >����T"O$�A&NěPc���e�%J@�p"OX��a�H����=1�˗"O���K=&h5"8+V(c�"O�<��_8�������(i�� ��"O*4�t��Q��ږ� !�`���"O��cg��"u"���2��`�"O�Y�!$}r\öL�>2�Laj�"OR�Å��,,��#J���$�1"Oj��AD��j�f�Y$�2~��"O؝��*F6���qè�0~pr4�`"O�H8@a�6�rݰ2m�2STtz�"O8�v�b�Z�I��H;hn�x�"Oxt�VgGk���!�֩oZ�Xw"OR�2co�n��|YQm�/O�H0"O�0D۹�,ȖFY,\�x`�"O:����!V�z9��.ۺ�$�'"OL�2�� I����Mŭ~ֲ ��"O�)��M�?|A|U��N�^�T�S"O4����O)m�XT:WmU�	�V�J"O���(ERE(1��ÔX�ʅR�"O�(��J�$r�4�����&W@�{S"O�Q�d�^��:0ۖ�<3�4�;"O�bQ��}@��V%
�T����"O qQF,�-�� "E�"eJ��Ӄ"O
[�
���`� J�*X4�,�"O�y �5 MN��4��B	����"Olq�#�+}h�U�UD�Ar5"O�}"�M-e���0p��U����"O���'�L�d�a`� N��H�4"O�X�!`D�*$��yS�u��"O����W�4QC/��&�q"Ol�١#M����R�L�fc�!8�"O,8���",E�9���Q&qFv��"Obt3ף�)��R��X
Q�"Ox����< �����y:���"O�)׮Z�a�d8��+'	$@�;�"O"�X4�ڦ�б)Ϫc�:4��"O�i���Z)<a"��;W�rF"O����l�3s�h f�C�G=���"OZȣdúK,܌�E�>=DѠ"O�2���}��5㋟^�T��"O9��BO;o$qbqA�),\�""O�YdK�;8@�V@�[2�e��'�jQʅ�SU��́�M�2��i�'<��r���ٰ`_	��
�'�@��[�w���!�L!e�,ȡ	�'_�t[��	+]��Q �۸f �"�'��X�u
��0I�M�������'�䕂�jx	��&��X� R�'��`��n3�B��VJ��(�
�'"�,�a��6Q)x� 6,��
���	�'{�<��PB}�5L�$vQ��	
�'�V}��O�;8�$��S�+i�@	�'��LXoE��X�y���s�0�K�'���{���%E�!��֖k��s	�'2f�bg�;M~0q���T@l80	�'4�����niz90,޾}���'C�9䋦�f W	�[`�X�'�@�)j�>u�f���Q����!
�',y�Ԁ�r��Ei,�xXb5�	�'S�}P���p0ܱ��D�/_)�I	��� jـc�U�����%�b��r"O�e�B�aK\�Hrďz��r@"Od)��e`�-��A�9��\	"On��������D�)��%�6"O>�k�o��2h�8�U U&F	����"O��	�	dq.�:�e�5���"O�x)ȃa���UQ�x�p�"O����hܯ[�PAD���{�Hو�"Oh���W�]�B�Y���]̬T��"OB<�qM�7hn��� ���\`��r"O�¤M!	نy
�AӅwL�y�"O\}ʐ�K�#�"�µ�ӷ1���"OL T��@�d���m��
�DP�"O�(�t�$"ZR�p���R�D"O`��o��`�i�I�mܶ9;R"O`��n&;dȤ�w��c7���f"O4%�*�H���0�s-�h�"O(�"a�0d�aB�@�&�{�"O�A��)G�|��I�,8�V�"Obx:h�q4�%��ٗC�֘ "O@�2�݌BpK�K�Wpb"O>�k7�ѓ:sL4H5�/�>��"O��{u
̥@�z�c�jT�>��"O���"�ωآ��!��M�����"O�-����{�*�z�G��%u�DC�"O{ᇍ<NĵCUI�{���"O��2Gǹ��@ײ5�FpV"Od�A���� uj"J2��A"O��[vB>iI�@ pf ��'"O$�xDJ�^�����N@�0"O*1[Bd,<���Ip��B�lEأ"ON��`FK�[�P1B���1�S%"O*AB�G�vljٳ��7y@>��1"O^����A�%B��z�g���4U"O�9�R��mm2�`'Ʈ%g�}Kb"O�}�e+Lp��J��#.l���"O��c�� �w��b1'� Uy8��"O�u�@ �<���!�f8���"O�Z��NyX�s�a	�k_�9d"O�Ѳ��ՙo���8g��Eص�'"O�Ŏ�4J(;�a� 
6�٢ "O��ʕ@�6U�����=G�$8�q"O~�����/ S&y���=�	�D"O��q��QɎ�[�$G��ƹrf"O���P�Ɂx���%��ġ�"ODU�֤2t�X4�N�`��ہ"ON�V��E:8�V���ݒa"O�K��=�Z��-�����s$"ON��S9P���C�>���
�"O ����B9~��Kgn�/%6>]"O��r��I
%�<����$jp �"OJ]*2�O�H�Ӓ��3L��"O���7�M�MB�q@э�g���"O���Ŏ* �E�C�O�X\*�"O�lYdf�/w���K��ȼO����"O><�"��'�=���ݳ�p<��"O�b�n�؁(F�I�y����P"O
��b4C��Aqo� �<�£"O�S��8'Fȹ�`ы��8+"OԙXG �u� K�e�u����"O�1�BU�b��  �K�C�E
�|�Rc�/8U��(!��C�I8_�t8Ц��6x�yB��@�<B䉈|��ٸ��P�.��@�&�oKB�)� �<�7�^�|G؀{A��o�����"O�AȂ��.d��
7	��*�4H�"O2��q'�5�P�!6��/K-�4"O~�0�fGu�ep�SaΕ�"OFѻtcLD�R��� �0K6�$"OJX�A�F�`S��T��s"O�=�2��T v];V E�'&�E��"O�h&#Ի|�LI��[J�D؂�"O���) [l��NF�v�&!��"OtA��@�&vu�%	��O"ݶ���"O:M�A+�"*(�{@��"u�̽p "O|p ��Ӊ?�){E�|�ޠ�"OV��a��J
F= -�)�$g"Op��u�	�<׆�+f�Z-Bm�"O*�)]:8�tqu�YAV>��"OjU ۚks��jOb��q�b"OHh҃�$,� 	�9_�m�""O�j�ER�,|I	��� �r}�!"O6Ӆ�T Jx"�� ��'�|��"O8��/���b�	�f��"O�ɑT�N?�R���Z�<�ڸ*�"O�=#%A#
զ�i�蜬g||L "O$��0b�'PG��@�Hʌ�{R"O��bPM����g�;{�&�I�"O��0��F#0��(�F��*��J"O�J��Q�Q�B�0s�.���"OR��KQ:hA �bb׽Y�FU�"O>u:�.-�^<:���T����w"O�Q�&	OD^�\s3��8��'=�S1 �ˁ��9wVp��'lXj��B�
aa"�c9��3�'���m�)^�k�M�,W֜*�'�z��0��d�0Q"oTdt�i�'�P�)�$�P��c	��L܈��'xK�V�����K�J���j���'�h�	 /��s��
|@TQ���WB�ɗ>5����Ɓ,��Q ~`�C�	T��}�	�kĨ);!Г!��C�I�I��A�\.@!F�
RLS�6?�C�	�n8հp�O�m��q�ԥ,a4C�ɢ[۠��̓���@�O�qnC�I.>��Q�N�3Q��BQ1XV����<��-=��"vN��@x2�+�bޢ��>CF���B�fI.)@���Ch`���&�)� !O7H �{0G�9ژلȓ+1Xp� �Ԍ/:*�;�a��j�����,cp"Cb*���ծ)��
�� �wʆ�<��8�)
�"�H�ȓ��Y�fͼZ����"��/�Շ��OyR��`���#�Oǝ'y�	0����y�Í.OҨ��_�L�P@"��x��'�5�Z� Y�gԌb���'	�y�@/
\EHP��$;�(��Ù0�y���!�jEA#(K���HEIV��y�<gژY�@q�r`f���y� ��y�@Xkp�X	8&�n��yF�=-��{���q>��慮�yҤ�-O���'������Ƴ�y�N�_���U�ͻ����D��y���X zÅ�)��5���H�y��=�(�s'�5k|��p�K)�y�J���|D�)NU|�52%ˀ�y�
_`�̘1D� I�`�rU�	#�y���I�d#p�@�=[�(�(��y
� ����H��@y �f+TT)A�"O ���B�B������(���#"O~1�v T�RRp�7�7p�l\�e"Of��*I�wuhi�R�Q+4���*s"O�X
�jU�H��#����� ��"O&�Sm�8�h]�1*E#�Vɂ"O"�a���?W��A��3ń(1�"Ob�[E��
WΚd�t�A#H@xt"O�]s�a�� �*sL5a0>I��"O��R�'K����y����%�(A�"O��E�>>�zE@��'��mi�"O����x���H�gV3-�f���"O5ѷ�Ɣ?�h�a�]-2)����"O�U@v
\�EB
`�4�M;6(�qr�"O�pTLעi��A��W�Q�Ȕ�7"O��
�퉱k,UЖ,]�R����"O�R�M� ��Sc�܆b��١�"O
�v�H)� �zpE�F���G"Od��U�U/m��0Z3f\%}"�{�"O���	�~�P�ɟB�\��"O��ǉ���P!#�Я9t��&"OK�(D�p?����5^F�	�"OT���萎We���FaQ�<U(�`���F{����<)��	�7Sq�r���,!�䘋Q{.��&#C�t�$O��!�$��R�d	�i� 9��������K�!�X�z4��k��G���q�ё�!�Ki�)��+%f�ms�L/$b!��@�@�^8���c�����U�Ko!�C�|,�U.sC�j���D��B䉞N�%9�&���Љ�\�p:C��6 �z�
2I�5�����M�*NC䉃Jµ�`�9`�[�%?5C�B���t�0㊷8�V�0���@�C�	��������H)��J�?��B�!G����u�"��f�
�+��B䉯x�#�oS�q`"�%�-C��B�I2 �XU�m>�
F
ϊL&�B��U�� �힋t��	*�H�7Y�B��J��(dJ;?b��F�*(��B�	=8&Nh:�CČSzpab�G��\CTC䉮B_�,�v��U,J�O��oy2C�	�s�f� Po�C.@ꆋҺ_�pB�	6Y�p-^z������� B�	p��{я I
mp� B�5S�vu$�H�[������@��C�If�U�Q�Y�c��q/E�A ��$�>i�*��Ą�2d��Hಀ$>!�d)�DW^�\�^t�3b~��I�<����.�$Јm�H))`�ƹ�=)���0�!�Ĝ�$�84ÄL�$	e�dIp]�z!�D\H������~ !���!�$�=	����[�l�jm�2'�i�!���͖ԠT�O�^)LQ���'!��A���r�^3f ��C��~@!�U�h$0���'�rqs"�]4
!�$C"z��ԈF�3�� S���!�D�(�@æ�Q�,B�L0�A,�!򄝜\���VY�j(���P+�<d�!�ę<s9v)Ro[r- 	�%���!��Ђx���8�GH/_ �p�g��{�!�˻O}�$�4�Qa�0�X�K�"O`��2�H<F�.`�e�F�}��ˆ"O��X��U��@�DK3 g6�!�"O� � ���	V�"]C!$C;��!a�Ob��
�"��-��
PE�v�:����!�D�/�MQ  ~~!�rd^�Py�럮/��х�Ҫ3]"�X`#���y"�ѣ*���q&����J\�7����y�E�Y�]�-�D~���glڀ��'��{��[u."�����,jl��K�yr	؜^��EI9�05�OL�y�ъH��!ɂ��saR1sq�Ӥ�y���,t�51S胁 ���˰%ĵ�y���(jfDP�薑h����
�y��� ���!�$e��թ��A
�x��'�82ŠR<��t�2��A�(����OV�}���T5��'�ś~��m�DD�<
��5�&� ^�t ����<6��ȓ-�ؠ#ѡ���,�t,��f��ȓ2�.���G�%P���v)ŌkWJ��ȓ6x軶HZ�dyq��P)`��ȓv�����0��YUe��boJu�ȓP!|x
��T�b!��X Q�R�^�'��y�JR�]�P8���)L��J�m��y��'er�{fȒ"Di(t���w�p�1�'� h�c�̭���CM n���Y$/D�h�[� �h�腫E,��x6�-D�)�"Z4�B�ȑ(�^Ff�C5!*D�h��3%QZ(����f�f�0��)D�Ĳ��*z��M(bϫ(}2� 'ffyR�|�O�ўT�/Y\s"i�Ƥ��J=�U���o�4��	=à�;3��-m��:&e}��B��s_B`c�A`N�q�UL|B�	?f�{�ˉ� �%���I�}�C�ɮq���,��z���$G�/,XB�ɫZfdp���T��b
�#0�4B�&3J��NX
�xыɌ���$%������AK���`_ԍs�% "�!�ā�t����/�6.v	��ԍX�az��ڝqXt��bG�b�a�@"Ȃ L!�$�)�R�JS�V�}�$E"�'�i�!���"FA�A%cT�V��S��Q�!�D\�����,ς:����KX�!�DL>Q<�a�/D;lb�р@$��3�!�$��
z��bt���$JF�r�B�)h�!�d���	Á$ �\��P�n!�߷Q}�{d�I3^�d���=kw!���H���	Hj\Q2׭ H!�d��Bk��8�a��N^|H2!�%`0!�d4qI�034�݋ D�`@RA. !�ȶe������Q�+��8r��S�!�d�Q!�*�$�F������<�!��)b��hS���1Nf������\�� D����W��	�r@M�R��)Sg��y�HX��`A;y�i�"+ـ�yrI@�b�D���K�'|1D;3��4�yң�i98=#�K�u�� �h�#�y"G
xaX��B�:������D5�O �����5�����kr~��"O��� S�Vj�c����pa�"O^�H3k�hľ`����[r�|�e"O8`:Be��H*YRԤ�'3*ث"OL���)F���uC��p!�5p�"O�f�/.�E�q$�%\(L�ɇ"OI	a�(z�V�jS��(���%�Ş��eKX<y2�?�������
	��J��\�7`�d�}!�� �] Z(G|�]� �'��3� ��dI��Mg��F��K�-�3"O���e�g��,�$g��[b8�x%"O��c�A>A�Y�Ҁ�R%Hv"O��b�NW �tu𢁊^Ӓ�x"O|͈$d�<ɞ���2Ml.�C �OZ���N�'H0�����r|x�G�%'���'Y�&M�]��f�� ��a@�y�)�S�=�.L{T�Z�^][F��ru�B�I�l.V�"���\�d���_�s�B��:kX��Ѳ"�t�4�[T[�t��C�	b'�}�d�	8�e�s��B�C��2ݒ#-R�~R|����3�~�	Dy|��i܃NБ3$����X�.�.}'!�T42^\;G/�� �����!�1O�$!�)��iKf�kE�_"-2��g	3I
h�ȓ��IzfjJ���蒣�]1e\*�ȓi^�)4�+,{Fy2D�Q+h����ȓ0H�ܨb L��أr ��DH9���?!ֈMX"�u"ue�=MD\1�f��<���S3�@�0f�Z�Iܺ��/S�m��IF����:`��<� -�/FPV(��J,?�������q��W	x�����Y;
��gc>D��zd-//4j�o��tv�)T�0D�4���ܼB��=w�:4�ԕ�G�.D��#5/	cW(p�Q�P^��MӅ`1D����M��i����iP�'{���R�2D�X��Ay���C"M�{lx�x�N1D� {���F�I�3d�W+L)�2%1D��Ye`ȋA:~m���M�o���7�1D�s#l&P�B�C���8) ��<D��!�l̾m���ҧO�.<��l�0n%D�HI��M�,VR�̓f�ļ�u�#D��PT�<- �@sa��:[���FB5D�lQ$�ȋn��1ȕ	�31l�	`�(7D�p�A�m~�����Юx^Lvi5D����f����=���(UF�8�f!D�d��5af��eA	(a~2��p�<D�lF�T�0�1�3�u�`�'�-D���wₕ\3�|kՍ�{��x��+D����(��L�p�Y��Cw�Lq�k(�(�	�a�Qc�G�,:�da�� ��+fPB�	�@T���H��PG�<�rC��<� -�s�P�b(��ӥ�;�^C�	23kBAIG��$!<څ!'	��DC�ɚܦ�kaR�#���``NP�& tB�f��� �f�����O�PV�C�In���"�(�?RMt�Ò뉙jc�hG{|�B��Q�f��l��#�mibC���yB�v�8r�H�(�k1ȏ�y��)�'$��UKW�t`@]H�	@�7<ԁ��%|t���J |׸�[��B=a����ȓH5�a�i۳S������ǹX_�Їȓ]�"�fE�?10�����)y��݆����:�p��̒�{|�,�m��<e�T�d|V�$j�S4x��-s�<��'�0cc�h�1k_�Bv
� ����hO?�	2+t�|��A�N	Z��5�C��9&�Fu97KL�4�Q���8(��C�/�-*�sED�_����!�'���1@,U�"O�l��	#� �[�'YP���oI>�ЬX��½D���'���3�Bu����D�aC~ݲ�'�I�i���HAEA >�����'�Dq��
*���1���m��2��� t�X%��8r<i���Z#Q��iIE"O�R�.a3�EYV��(���2�"O���PdB�Y	r�0���qpP�J�"O��!�����3�@�,	��S#"O��`�D�m=���VN�Or`;T"O��Y�*`�UX���i�r���"O�؊蒘d�9 �茀�L@�"OD0�4�Lg� HU��8
�I�"O01��&�/Ej-����X���j$"Ob�x4�U�;fF�#����`^�P�a"O�����v�ye���
X�y�"O�]"ȷ~��X逢�7�V�P�"O���1eD�Q�#��.)v��6O���dۊ/Шiz��E=��Y��n��oI!��
~�����V8�D ��c��9!�DY�g��F%҅4��9�"�=I�!��U(IUt� L>7��B�~!��
8/��$�g��,���I��D�!�$Ŭ_`��kF5a�Mҥ�0�!�d%��m�6g�!w��A�@ W�
Τ�$�<Q
��P z0�&T!�"n�#����"�"�ck�<���R"��&Lt�ȓ
C$K W!Y�x�*���If�I��*���8��k��<9����E/D����#�"�T B 	
*"��k�--D�xkf�^
4�*�I�a[�1:��)�	ן��?�|��eٵ&��sCfɋi��ґ��P�'���S�O=L�)"�ֱ3�z�����a����'���y�t���x���y�}�'�L%�֤@�&�p}��(1���'Z�ԡ�O��E�î&����'7�����ʌ`���B� �	fr!��'K(9!�;G`�늉z([�'4�L�H�RlJ��ˋ�q(�=	�'��p��%K�(s�x�!��7�h�b�'�p�Y�	�=u�P�0��_#���'�BTXo�M���+��O@X�"�'�&�B��!8gn���ɖ�u���'� =���١>Vl|{g#�mW��O��d7�):(O� ���n�~�1u��V�vٺ�=O����0b���Z��N�T�� B��kf!�pf	�)ʉ>İ��䙓';!��#*��� ���$o�<���D L!��:djȻ�� B]�8�c�4i!򤝀;R�����_�m"�!���;`^!�$��d��$�Iq�<yQ�`F{ʟ��` m�?�:q �^I�1��<��};:�c�"D��U�'T����?����I�R��0�@�5݂��L��[�!�
�f���C�Iϰ} w�֢/v!��ޭ̮D���	�[�P��tkƙzg!�p�`�	Û��=�c�ɦTA�8�ȓ �DkOQ8��W�Q=����?Ʉ"G'�,c� Y�]P$��<�
��3t�e��8W*t�i�@&&n(����?�H>E��'�x��� h������!T���'��C'�ڇT��3B�|b�9��'���r'-R9(H�j��z��i��'� �B ��O�~�;��O,}}Dm�'H�u�g��(8~�7��ml�;�' "����/�P,AWmǻYP�' �mѰ�Mw�r�F�5E�h��
�'w��b79uN�#4�֡e���
�'�2a{�����H�0���P8�	��� �K��B�N@��V�S��`�"O�C��ӕa/�T��O�j��Y"O*��p�gP���,�/4�8��"O� (b�I���ô�}|<�F"O����ώm�<ʢ(E�L�L� "O\�g�&q,auMP���pa�"O,R2O ?�X9�ċB	�H��"O ���	��a�J����V�L�2r"O����EO�OtP���\���"O*�X����%9&� ��F�� �"O�
���G��ty%bD�=�h Z�"O��;��`�������0"O5��m@]b�RA!\�B-@���"O����o�N�rB�(�J�"O�l[V�
��N�)ʙ0"O$X�iE�N��@���즀��"Oܸ���ݶR4��X�f�(c��`"O���ʦ�D�{�#�X֎9��"O䵢c��18�`��cC#���y�"O�<I']B�Գ���$R�"-"&"O"�E�ϸBY�K�2�X�"Oz\�0���*g��P�j�Z$"O!��(�5� %C�K��n��"O9�bJݶOF�02F�~JeP"Ox�k�\�H��g�"B��IY�"O��If�CUTR����-q����"O��`�q�j������ ��x�"O�	�.�lU6P[�Fȥ-�i�"O��г��X��8K�D��y�X A�"O�Y�'	̚ O��TJ)w�iт"OLE�¤0jAx�i���#�
e)�'� �����P�AX� .G�:���'��Pإh����*��"G��K�'�\�o�.O#b��1�ϘB�� X�'����V%� K:H(���O��܂�'PV����
i���8�#�"�N�!�'k&0�$��)J3�t�B+ȱ^p� �'�t=�n�Aq\A�!`-�$�
�'�l�˵�N�h��4+�&	�,��1Z
�'���x��-.o<s/�n�FDC�'��R�o�A|�'Eʮl �x�'q��[����,����5)S��I�"O��Bb
���p�J@��4y�A"Of��b�:?"$���)�
/n�	�"O�Hh����-À�,/m2	i�"O^���

�9������o�8���"O��#,�3dX!
��O�	|��"O =�A.G�!wܕ!Tʟ�-�Zՙ�"OT`t���.���7��Tx�� "O�!��i�7y/r4�p'b`��H�"O�S��ɾ7)*�9CW@����"O���a��BƊ�Q��Z#�A�"O�q!�?�UC`%W7|5HKD"O���g�?��(��>.���"O�IQ/�(I[(�C����˃"O�=ӡ'��:�a
�6���"Ox����&Q�~��@"_��"O�$�V�Y�b�t[C�Yr8PPѐ"O|ʇ�̩w���qk�>+���"O�z��5���p��)|��q"O�l3T�ZW
��j���$F�ي�"O�ea2BفL�Y��Y���-��"O�%�� �47־X�b
Jn�H�"On�{��Кv,Ԋ� M'��-�"O� �H�ƪ�9I6䥢u�	�}����"OrI���G RF.�*f�pY1"O0�ٵ�5ZA�Ҍɸ"V��)"O�@N¤}u�,`�,��c: �
b"O��C�%Uv�aPժ�=�"4�`"O����m�Bhv@�HE�tR�"O��I���.0y��ݰ{��&"O����X~�DQ6��f��F"O���`g]�d˴͊�+Q�Y=���"OH]G���>��
�]K.�y`"O(�����8����Q'D�c"O f�Xn0h��d�f   "O�E2��A;l��FT6���"OX�X�f�E������:� 8@"O�5�r��%��P��ǠS� R"O�I3p��`8���(Q�ƺ�i�"O�0��LٰF춥q�HȓP�\�҅"O���%�K��`0�eM<~ž �"Oj�8�%/p��C�����"O��`C�4`M�Z�Y8b��t��"O�9K1��v�`�d���T8�"O~�{׉ �4�tj#��;k��,�0"O2��Τ�������7_̨(Q�"O��@��(/�Y#ᜟ9��ػF"ON�����\�����t��ԺR"O*�q�B��d�h��@�e�Ҩ��"O<��0-�qaQ����|D�+X�y2� ێ1ѱ�T�h���=�y@�m��lȤ{Mp�(��Κ�y���~�eY��֬Y*�3aG�y�$��4=B��c�R�M}��Q	*�y����̻�)���Cad7�y�k�l��ز�
�!N�=�0��)�y�(_�e�k��.'�I��ybB�m�Q@D��eR��3��0�y"b��Dp���g��A阁;֩��y2��nP����F٢��ug��y�N�
��D���	t��|��Z��yb�)N�q#ǆ4>�`�ٲɓ��y"C$ex�4�b(�()�`9,Ġ�y��F8N'P��H�/�F\���ȳ�y��M�����.;���:���4�y�i�.�(�t9nzy�,ȼ�y���|~m(�1�� ��J#�y�S�:͊b`��&v��ӗ���y�^�hʌ��I�H��(� ��y���k0޺3�4�2�Kڊ�y���,���#Q.U�x	r�K��yҡ�֎�ɶ�� �r��n���y���uN��P��:X���V���y"�U�z�5r.R�"_ʬ�E�3�yb-J.y��%A�ݶi��9Ae�D��y"��s��5-N�qj H���y� �q�p �(I�H��3O���y򆞍d$;�Q(��
��ō�y&�5uJ�rD�h�j�BN��y��L� �N%X���\Az`��y�oW�1���S�ϗ&�<=�`oJ��y�,���
��7�Ӕ^Y����yҠ��UwD4#Ջ�����B��y���-	OZ�BE@����A� �y2���W��㩖�ht�5#V!�y"�I�pkfN�;�ll��Ą)�y�)խ}r�[�>.h1�Wj�y
� ����`Цo���zc��T�NM�"O^���KQ1e'la޾t�z�b�"O�� �#K������7����"O����ۀ;��б"B[�j���"O,��w�jV0)ׁ����x!t"O�P!v�[�0�T�����.�G"ON(bC�'^T��@K�u�&u*�"O�{�#?�L�qc�Y�+���xt"O��BA"�>5(���"Z��Y�4"O�A[���g0���'����� �"O�DG&�]m8�� Z	zTH��V"OvI�p�[�W�ND�p	mIs"d��y��A	k-dM����-=A�[�*��y�!��UPr�V�Q�H`0 >�y�G�G*��2c�~u*Q����yB�Шߥ߭w��I�0e��pE���ȓA�q8E�������J]�n(౅ȓRȺE�W�	�<�D1r��E�D�0��|�^�X�1.N����2q�|܇ȓ���$V�9�!.�1S���>��v��M�l8�ڑYq���;�^0��2ľDA��3��(��"@?�)�ȓZMd0殜�RD���T�8����]B���F,G3�b8�B�Y�bD��ȓ���A�E
}V�Dj	��o�$��ȓ3ܦ��c햆�8�Z�DI,ӂ%�ȓB�.��D��ed@(�$�[�uVQ��2�64@�˱�`E�&KH7p���?�pa�Qټ	P�猳 �B��*�B���M$g�arԌ��h0B�I?����Vm���Ec��J o�*B�I)PB��;�O��<��qb�ÞPB�B�I>X��sE���Z�~��`OC��B�.@�z���'�p�3P��w�:C�	9��q
B�XyiԀ�2�C�	�]�Ja�H�vx�@j���6��B�ɴ\���J�C�r��x�ʛ=�*C�Kj
#�`P>4^dz��[8Y(C�Ii�J(�UDD�jh�JF���Y�8C�	$j� ۱8�1�v
�%�lB�	K���b�]�	i�Щ�DܑsT.B�ɱ5_0�"�EG6Y9���L;K�C�	;�6�ٶ��=��` F
R�#��B�I�ut����]&Px�q����l�nB�IS�����FX #|���σX+C�ɔAΎ��i�y ��%G.+�C�I����d�(q�ʹK�Aή#�C��]�����9n0������m�C�0Q� ѡ��Hk �[Gh�:EARC�9i��y���1Je��ã��:m C�I�	�2�b g�@������7�C�	-	6��@��?�,�W� �+�B�I�u�ș�+��_�$�˧��5l�B�	�k*=HWBˋ0���T��-K@B�I�U�Ik�������s��;`B��*&$(��U�l&­�c��o~8B�	�X|�tka�Q�˟�z�B�IR(ؤ �	�Za���
5�C�	_S�T�e],	����l	�=ʰB�&�$��VAߩ9�|j��Ǣ`	�B�	�TSJ�!d�� TC��G
�0�>��8�S�O��D ���<E�RE#У��y��"O����Ʌ0
��Db��g�5�g"O�-��\>���ߨzИ�4�H��(O�π �M `�!oIi��a`n�q��D LOm�d�ŭI�~)pB�V�wበ��<E��y��Z��j����WG\p�<�ďN9?\|���5���#A�'ga�Tlց�Ҕ����$���mB��p<Qf�\��7��%3��@$o�T�� �bjȍ�ȓT�@�R�	t�����e94)�O4�=��T��2�AP
\��YQ��c�<Qs�� �"�)��ˈ<YP��ue�Z�M�a{RIL�N����.�(�au�ߴٰ>)�����U��Nw�@������� ��5�	Z���O��ℎԹX����D��Y�'�B%���Y���C-�'6�ti�'�m�Q�����ab��^�$hs#^�������w�A
bf�8$C�xpD�
�x�!�¡n�"��d��[92t�s��8!�d�j �����f0�APWn��B0a|d2�R9c�8�z��γ8|t�J�!�d��H���� m��I�l�u!�Dݜz��(R�� y�lP8�lG!�$�[]T]�T��6)a�&�0f�!�$A�x���A*Ĺ,��m��©|lQ���C�+�Iс945j���UG�I͓��'�"}�'*�H���U�x\�CAm�V�'�6ɖ:���xe	�B@�}�M���y��8-�رrDɂ$y�a��l>�O��I঑G�4�@�
(�K'"�e�Z��aV��y���dѸ=�Pjƫe(h�'�����>�O�T�Q@F�Xȴ ��/�ޮ��$d9}��;�O��畤9VRDA�A+H�M�`"Ob�c�����Y@�"jFr�0'"O�}q�J_*���$9$��T*��O.����_�
ÕDyR�|͟H!�̸7�=z��A�kip�:�&�9)�	k?و{��IB�L������/u�� ��=�!��6�R4���]Yp�	��ҏ��l���oX��;�
�L5��d��D:�G�#D���L*q��[q�*�R8c6B��xR!S�ȾIX�45"��;v����'�ўb>	��ٛ�཰$�˅d.	+3�=D�` �F�S�h����H�+��Uj$�;��D��ħ���GȜ	a��q2�b֢A ���ȓwK�U�S��jh�Q����i�����~���[R·Ll�qY��9n���1�>KU��,�!ҪF�!Ħ���yy��4�׵|w�M���)U��'�H��4�qO��
�CC�$q�l�k��"1o���'"Ol���ЊA�l��$L2W�*B�nӐ"<���D¥:pD���\�9DXq�b-�x��O��&�[s+�����7ΐ�3�&�`?D�(A�	��n�P�;�dT�r?��!��1�hO�S.Vd��#�}��Q��a�?�C�	#��9Qc%X̪��B A�6+���/�S�O_u���	*yR��#
�W��b"Onp{QmA�	���*���gٺ|:";OP7�|x�(��)J��u2el�,����i�O��=�OD�'�����*/�ԑ���5N���_�' �y�d�N�����a��i�4/֓�y�K�E`��G�+w��Bsi��y�c	��9x7��/�*t#M7��!�d ��X�eG�+c�h�(C�_. E����"O� ��@��sC)y��`K�H�OD��l�IV~J~�9U:S��;oL8L�	A����ȓ<{й�t�ρ+(�PょO�/~��=��S�? f|CP�&=>��PgLG:2\z��"Ot�R6(N����:��42�й�"O>���W7n��*)T 3�,S"O4��ʌ-K}����X'wR=�`�	K���	��i�&h�ujM�wi8���B�5:�T��w�=�S�4dS�j
�}�GL�?$f|�%�E&�yR#�"m�BXxp��+?~&h ɚ��y�b�=1�3�荩:�6h��Ř��O0"~2�Ǆ���p�fa��xV���1&%#�!�Ċt�� CJ>O|D��Gɶn�!�D\���@
��	-rH>THR�0�!�
78sP��O:]��J��m��'�x"=���*nA1�f��I���8&�!���O��0��\1�<��`�?PΨE8��%LOf���* �NpH�`u�rP���Ir�O����D�R|D�t��S��!y
�'�`Ԓ�X3��P���D�e����'T$i�v)<�r�1M�7EЪ�'m�[��b�C�i�h��*�d �O����6 A�h�)QJ�XY3d�x����[�@�N�Z��	&{D����M+t�r�����Raq(���g	�e�zņȓ|�l���S�L��n>U�"ņȓw�"��� �TD��T6�nLFzR_��Fy��]5C�
�A�G�^��$	�y�o�I�D*�N �e�5�ē�hO��$ě��B(-,���
�q�
�`�O`�d�@"��Y�dη��`b�lF��O%��I��$U�×�Qv�}a �j��C�	�s���٭p3�=�+I,82B�n�>��ʅH��vL#G�XB�	'wG���2#9�d���ƕ5*3�B�I0����b��8v	FI�%N�e�c� F{J|j��˱��y�� ͩV[�\`���F�<�U���Zy8!�C+/ f	���QX�<!�E��?J�tq2��~�R-J�I�T�<)��G�D��x�Qꇤ5����e��N�<i��R�glD b��"5�(����N�<Yt%�/A�u�&MJ"uj�NTa�<)E�D'0+�����X`��[�<y�fY<K�4T� ��;V����d�T�<��Cք:V$�3M�90����V�GW�<q�܊|���3��ȰZ�<Y�i�7�����_P�n�� �R�<��(2A@�(A�AH��#��D�<դ�ZDI�-�:t�)k���F�<�V*��
����%GH��ت���J�<��.|y�a�Q�$��d\E�<ß��"����[	|q�ekFH�<`l�-hq��,D�Wqxu�U|�<iDF�l��y���;*���S�<�E�Z�xĒRbU�eW �x�<Y�-ΪPt��r$�3VƩht��y�<���W�!�Jd�4`#���n�K�<��� ��D�cI��~\a�E��]�<��I��!�DW ;�^@��u�<y(M;~��(����U�lQ!���m�<���F�u�Ũ���5>\���l�<�q����hXvԲ��i���So�<�q�^��3dۇ�
i���h�<�Rf��Y�m��BG�iΪM!��L�<1��G.a���۔�ڀr��J�<�G�O"�Bp��ɑA�ĕ�pgD�<�a�Iİc�I�L7ƕ�L�A�<� D���B;1P�+5��:�V݋@"O���WC� G�LеG�|�J-�p"O��Xh��i��2���r�"O�$)�iۓ$\���'_�^���J�"Obx�� �����\1���"Oh��-и{�n衱F�-\bXx�"O.@�GI��\� ��*dH@ S"O4	���*[W�� �ףd6���"O�u�v#�*B$� �V�_1�9×"O�99e�T�E"��� 蝍�&M�"O4]�c�?��THZ��m�%"O��)���%?���@IDz��w"O
����@�\~|�Q�� fX+#"On������ ��(b�eP"O�d�m�D.Y�ŹT�l���"O�p��K��6V(�+�fO�0|ԑ�"O� s�C`E��FEQ$hց� "OJ �RNδSD(5�gEAR*�p�"O��B6�\�Y�x�[�$
[��5��"OJ����KG���^�`�"Qs�"O6���Y�r���H�+�	�!"O��I�"S�M��;5�ˠy�vd"O�����1oZ"I�w-$�����"Ol��!���Tɫ1�D�o�٢�"O�� �ջ}w�,���X*ҨQ��"O9���֛A�b�#T���'���s"O,=���A�7]�����&5���je"O&�����m�\+�Y�o�Ԭ��"OxA�Յp�X����J�"{	ے"O����@�a�8&�O�Tu:�q"O\({A�P�Ѱ�2A��s.|p�"O����F�vP��&lQ"tc@�R�"O��r�P!q��'�ȕ}~�q�"O�j��ڮer}�I�W���@"O��!G�b��ō�j�0c�"OdKĈP�@6�d{B,D�TQ �"Ot�-���P��EЬTS@"OXl�ёy�ԣf#�Wgލӣ"Ot��V�؜;��%Y,�"Q�X�"O(e#V�s76X� ڂzd"T"OJ퉲��o�u��h�M½yC"O(���`E�@ZԠ+'�Gh:v!x"O�<����R��,���H�/H�l!�"O�����7s�Z0���X!"O�E�,G�^+ 2�Ƃ(P�k�"O�8РJ��(- i���"$�)�"O&�ҩA%_M|8��L]0/wn43C"O(}ӡ����!2 lԕpsh�ʀ"Of��tT�y���p���Bm4���"O�����!p{�M	�͖7����"O��ifD8#D���EtН��"O��G��`X��`��d� �T"O"% ����0��Ó��-}Z��� "O�������_��P��9!;h��"O�-Y��D?�� ��[��M�B"Oҡ�b�|u(���nW;�L,��"O(0QL�{Z�D3����]2��0�"ON}HEC�i|�pѬ۰#�X��"ODرdM�81RT)4K��.|`"O@�aiH��\�Q,���Lu�"O�xAw��%rQ��RDi�x� ��U"O�-�4�&cm��1S�'_�d���"O����9V̃��\�a�x98�"O4��O��<ɂ��@�,��"O� �Uɡ��K���Q�j\�2z)�"O��
D�L=OC�;vh2"OH���%F7�\Z7��6.r!�"O��gCǮV�])G�;3B���"O2)K�m������$d�E�!"O*�@E �^�F5�3��0@���!F"O�I0��:zn, ���	��4I�"O!K�oE>uCJQ)K��v�P�"O���u#-����%9r�D�"Oddk����*fnI�����X��d"OJyH��e.��d�t��l�'"Oҵ��S?2P��%ܙ:�`	�"O�	r�׵ �&y��K]���a�"O����剂Rj`E���7E�6ݪ"O��P���]�\��UY�"O>��)b㤅�aaWK��Pqp"O��˒�E%A�.$�D!��1�`��"OP���o�B�9!�+qPQ@b"Ol��1)�16��+��+@�%"O<�Z�'J�'���sɚ>�@d0"O�㵠ҙ\=j��1��2����"Oz� ��[m{\�wfE/n���g"O8u t�û9�����ɧ#� ��W"O��s"Ä�ic���dR3#D��"O��`�X><�����99�"OdM�gMßqt(cf-��^�x�"O��[%�;�A��
Ϗo����'�ɮZn��3�gWM_��ٔ]<L�C�	9G�	��B�lJA*�;u�7�(��剀#	h�`�&(d�8��9D�h��H�!0��v��.�\�ҕ�8D��Ʌ��k8�K�i�c0:M*B� D��'$Z�r��(񬋏�,��G1D�!�c*\�\E���I�~�,�Qc*"D�PJ'�(a �a䊇�{�^9k$+D�CAA;`���BDA� �"M��!(D�LpR��U�Yصl���C %D�|0��	�$n�3Ң�!U�D��(D�\J�B��K�&<8��=/.]+��'D�h�s���l�xY�b���8�ոm#D���G`K�ꆘ*QF@:�@�1�6D�� �+�`jT�\ H4����5D���D?	|n��&��Y-�*b4D�8��.C~D>(p���+,ŋ� 1D��iAȪod���B
�E(�PU�0D�p�*¦ֹ0'�H�=��mKtk)D�<�$�!n�{G�G�!Ѽ����1D��2b-͆MԲC!%G�s@�щ2m.D�$���ŒF���S���v����?D��� N�b�r����F~A�>D��ShV0etإ���65��)���;D�@с!�7��k�dO�Xg�)*�d8D� ��)�P�(qSA�9ru�e�!�8D�8� �L� ��E��W��U���8D��:�@��@(Bd�ϡve`�q#7D��0!�W��-�J�i�4	jФ"D�`aO+ͦ5i�M�E�l���?D���O��U=rt*F�VsuTMZf�>D��*7/H�4Ք`qtE��
G*y� A>D�l�@�ؾN���1��-���2B�?D���
eݐ����n��� D�@!�ks�t�4�QQC?D��ho�"$Nz1��z�ΡpG�2D�"�Ǝ�~�!�!��'y�N웰o0D�� �첂JT�*��1���:@���P�"OZ=�ThA�=9�|�fH(���A�"OP��f��'& �É*?L�Q"O���w	5TtlP���ħ75(�*"O���@­jZ���%:�*$P��d7LO�us$C�%d]���W�H�
�Ȱ"O��#�/aN��!F"{G�A0"O�{G��g��Ia@>cj0"O2�A�FْS��A�dL�La�"O�	H���,Hj|���W�N�0�"Op�R�ͣ
�n ���	!;{ppP"OBx8��S"MV��F35s$�0"O�P(ܙ�<�`�EL�i��b�"O��@%�ڝq�(�ꖀD��L
�"O�E�ٝ��@
4��?[����c"O005��J�Z�ӃBZ!r�p�
�"O �ZW B�"C�\�F�}}X�C�"OƄ�5gZ:k�|w�܋}�`p�f"O���&I��uR(sA��p�1��"O�5���\�1��u:�K�~p<�C�"O�=Zc�.�.�K�
�]T2@ �"OH,��G�Y9�%��)ʝ%C����"O<qs�!ޓi8m�Tɟ�w*tk"O�� ��Ws.�R���K��r�"O��HA��~{�j�MJW��B"O�\�b(��N���%�M�8?�LK3�D(LO�y��`�& ��SQ'\�t(�8�"O=Z��]7x� ��򦒧:+�ċ�"O���3D�7�:�k��!6�8g"O���s�W;f��]�-['o�Й"O0ۤ� $�YY +�0�J��"O&��S�֗��p���4��]�"O0����9B�&LÆ��08����!"OtM�N�]�PԸ�@S�g�L�u"O~(�J�=��� �ʄ2�h�h�"O�Q��HZ�
yT9r0'��D	�S"O@��u�)��Jd�D9Y�"d�$"O.țEΈ{n\��\�&�\|�"O
���'��B�E<�4���"O���	08+W훉7Bn��"O>!)�lʕi�l� B�߲�S"O��H�̞m6D��R�i�Ԝ�g"O�Q��A�Q<YBM��r��5Z�"Op4ȗj�;M7�)'��9Z��p�u"O"�7AE�4��]�!LB�-���"Oz,pd�߶}|&�Q��4f���g"O��( �g]����E�8R���"ObDQ�DW�à�h�����rt"O���P/�"e�=У�2�.��0"O~��%�I���J��%s��1a"O��ò��26f[3�ʌi�"A��"O\T�&��>�����S�4Ku"O��/��D\ !���6� �8"O��yх@*q�Ny�a�����K7"O�l�p�3Ķ�H�A�e��"O��SCư�JGa�(���j1"OA�q&�'G��8�
U˄8	�"O|X��?� <��p�*��"OX���Z�l��ׅ����T+�"O:8�A��S��}a�jL��n<BF"O�,��������E�C^�J���"O)t�Hm��A@Ƀ-wMVI�"O"�z�Y�*�l�I��ӱI-��7"O i*�W�C�J��EC
u�P�B�"O� Y�b�	��ޠ{t@�J���"OH��fk�� I[ ��>f� 5"O�A���Wrl�2 �nV��*U"Od����RKj3� ]�D$�&"O2�(�/L�!5OV<R1�h�a"O��3q蓱n�PH1� �b��4"O�]1�/��0M��P���}�0U��"Ob�A�'Y�[��m��G�@����&"OR(�ө��7��tp$ |�����"O�u�/C����kr�ίoͦ��"O�Ԛ�bΰ@�4₴^�D�@�"O
'�"�<���
7�r���"O���O�,/����'�5\�X��"O0�Kp�P�Q��Y�A�үj�r�"O��f��"P�d4�a��>Ƚp%"O�[Ī"Fnti��	-c:@��"Ov��@��tό	U�Q+,�b��"O 4 ���L�,$ʷ��a���C!"Or�b���z�+&O�E^�]s0"OZ){��S3`��pƇ�f@��07"Of����C?mj�h1�阋m,��"Ob���k��@�k���\�[e"O�H�r�ϫ������'n�U1�"ORY��� 1�tM:BhS�~�a;�"O4C�o�#"���G�%螔S�'V6��Ĕ����ʈ�@�	+	�'jd@�G�!kEY#�i@�0��'�XZ��Ô7�H��ѧL(9Ep� gN&Bf$p�jE+r�{�(Z|/��?al�$[�	���y2�i�j!qg�;-&��[G�
�y2�U�l� ���%-� ��e���yR��$4�����/�(Y�B,�yrÓ��h�1�-V� ��Q�yrh��b� `v-� �|A��Ǟ�yG	Y�`�9�#�z�*�����y�v5.X`�	�	v��m�0�J��y�B6v��)��Ԛ[��)��A��y�'�M<h�@Q\�U�
ɕ�y��A:Lo��	���;/�f�rgn��yR��]0������k�Læ��y��L��bA��a҈{G)Ѫ�y�g�f[��Yn�}�|��-ѳ�yrKA�VR\�������a�F���yB�L���G���i���y"�G;�NMJ��_ @΄CU �y�Gϓ(��yqM��ap�����yRG�0&{�t��-%��Ic5�&�y"dӼ/�L@�TF��\�Qg���yF�}\˒+��H|���:�y�(Ib~��hw8�P��כ�y��ğ\�����`�e����J�.H��u�_>�˓+�8�|�'��ʣ�N,ˎ4���աb�'x�ە�M���h#s�,.�4Ȋ��ȱ\���0q)O�3Ej��
ד+�*�+V�x���C��%�%,O`��),80�k3*�
�b�p�Q!� 8���'
W@�<�g)�qG�y��\�� 3�F~��͹;3Ji!&�ͯ~��?�8��x��(��f�P�rcb�=D����Ƒ��d�;``J�y������+n� �,�G�r�g̓V:���M�~�bT!� ؋��I��ɔT���˓pX�Q�R	$��4�0@���y�뎫l~t� ���`-2 *��O^�p�����*�_kR�;$��hB䉣`�#c)Q�M�l峒D���K�l}Fx��I�b�`}�@����0À/�$�!�� 8ȑcb.j���cT�l� * �>Y5�Ĩ�=A��߀��	S�A�{��;��K����ł�򦍱QBG���R6ʁ2&YJ�4D��a�E^�"|�$�U�z-�%2�f[� ��IŤ"�����Z1[=2
��K��ў����9?���#��3y����G`����	i����?E��G�4;Ę!�A��$�p2��_��?A���S��"P��g�;�j-���O�'�"�O��zb�?lO�5pL@�z'n�P�ĝ���sTT����I�FA�-mڙe1�(���;r г��%|�>B�I���%��i�h�!�^$0S��>�����H��A��i2(���JL�h��X�p"O�6��*���S�/�~Hc��OTX0.8�)ڧ�� ǎI`c@�{ ��#:9��ȓ�B��l��uB�m� ��(?ބ�O���&�*lO��1W�H��;�lڞ3�0���'���Z��i,�)��-�uX��f�H.f ���'���b�N�I�\䂳��+y�T�=�)O��Ӆ�:��
P���\� ��̚ ��3
O6x���Y����]NX���,B��M�e�&㟢}�E�Fc�I�吴_|�"�x8�pDz�bS�I��𩘢3"1������	1De4T��I� _^���_:��0�ڪm�h�'uў�O�l�*�40�P�&�P��Rᠲc��L��y��M�Fأ�J	�FV(X3+�38x�=��ODг��i��a�G,t�U��ޝV�de���,D�D�F�^��2����LYx���<�D���(����a�M�G��%�v�ւ=D�HC"O��I3��.CJ�A�ϋ�d��|9����e�azR*֪;��%���#��"�)�Px+U�o�&�ʶ`D�_9�}���1=?>!�F�"��h#ƕ����I�,��9�2!p!+/,O�ɳ��\̓چ%�fl�6l{S$�T�mnin�p�`����p�Ae�D��*X�8hJ�
@�|�$��1C�}��'iN��|zt�
,�����k�y��<���\�I�^�tQ����ˠDb" `��͕���(6O��͸Z�}�s���D��X�wO>�
����l���:W�4���ēi}� ��B>�e�.W�b�.Fy��Ҡh�F���!d�P̱�ʲ!���)�.T[d5:���]��C&M����&�M�3:]��A[1%bԈ��_(���v�� _*k���&�8��@�x��i��i�����I;D�Bu���9ڦ��Hj�H��{����oB�E�U���	,��'� �ّ�~��Aٌ��c�{�>��Ą�m����C^�Lw8-Q5��d2�x	7�ơD(�� ��L1tz)��Ď/g}p��D��~�9���	F��2P�,�qOn���=Z*H\ؕ�����XD��,[5��9av}"O���7DC�L��I)�ُ����zI ��d(ߕ`H��dO�D>�W��t�rȇ�D�tI:e��>h�؄ȓY���#�JI�!�"@��6Mfԑe��=F��H{�oC&�4d�����P��?;J�83-�SB(���	�$y�ɦ!��'��($H�6��e���˸RD�hr0Œ����� �`D��(2���gE\�r��<�W圇x���CBCЀr����	e
j�ˆf��#��B���yr��>1��aseGþj_�tx�\$oo��{�4R~:����'��Qʎ𙟐�e.��X�n��LY,Z���E8D��� -��(�\�gh�� ��u�d�U
�\y�A��|�R�2���Wx�� �d�qH�٢k� =��S�5LO�`��J�Z�qgJ�!$��X�\!;�pU����"[��Xp'	(4��PV�sx�;Ɔ�z �!�5˘'A�2d�N58<�U����������T�(�`��k�
a��"O��4� Ĳ��Ao094����+O�!Z��K����d+X�>�7B�
��J�K¾䋰H�Ա��t�
 �0e��oؐ�3'g�B-@7� TVy�8pv�x��ɪ$8H��C�Ή�qi̲]�4����,rfjD"Ì��O���� T��� T����2ˇ4c�l�"O�|-�<̅���E�nM��3����y��q���5y�R�|҇匠 ��4���1z�@��t�Lf�<��'�9g� P�c �c�]	3� o~䐋A��d=��h��")���	��g�b`��H!�d�����d���Z�$��i
��\&��|����9%�ˆ�
%(���4L9Pه�=!�ZFnz�}����9���uV��c#ϊc�TI�b;Gw�A�ȓ��A����?R~]�D�j��-��Z �H�`(G.$��ʝ}a^4�� �(A��B�qj�T���`:�L�ȓ;�R|j�(	�xg�MFX�5�d���	�hu�T�D)F���"��"�:���l�^��ǊP�	(t�7��<$E~��ȓc��ux�I�;����e��r��<�ȓB���ڒ��+�$%i��Y�L����WX8p-:cd1��ɟ�!��%��z!4p!��8H@�ՊA�>e�ȓ77���2-hT|с㈟}�Za��W��9��c_�"n�dR�	�>L���Q����De�R0Fǅ�4ORM�ȓ��hzqm",j�i��gZ8Vg.هȓ)��h`���|@;ш��7�䙇�o���ᠨ�{F|!��&}=L��	�� ȑi ���9w�A�jE\�ȓo*F���f�5Uh��2CO�!9�p��ȓK`R����t`���JmPHt�ȓ��!�&#D�!fY�LOh-��NXD8�*�3IN5�,�'L~Ȇ�0_��pjŐ&��-�6.	�1�u��FJ��PB3��$�@�s���ȓCJt���@���-�f���Xe��T�6 S��|DԤ��� ?a}*��JV��#�+n68��#�>����VlZ]��-�3���$J $� ��gغ��e"��$�
#;$�Mz��$d����M�]�`�)>\:�  cg��!��1D�[�e��V%�a@W������Di�$�B͍�|��Xҁ!
(D�Ir""O� p�DH#`��0Oeex��My�<V�]:%�4���9R�T(f�Y�<���;dl��dl@2xd�k��G}�<��Α<(�-Ą-F�R4p�ax�<q��C�9��Qì+`���c��Kz�<����e���ׂ@����Ǵ]�<��f�����`ׇ� l,���S��s�<!pd!ܶz�!��N<CҢi�<a7��w��E�[��ޜч�i�<�g���P.��c"^�3v�� o�e�<��Cӭp�2��BkI��E�f,�D�<��AE���x��r�vHV>_B䉫O�隲ID�F ��2W
��;�:B�	6I�X�	�ǈ;wp�3�'7��C�ɭP7�Dق#چ	Vl��q�U�QB�ɑvD�K��G�l\ ]15�	�C�	*p�d����f�XcO��C�I�����ā'�fhE��,C��u(����O*i���?d�j���M?w|F��"O�X�P0/�0l�P�T��@"O�肂�_Q�V�C�ߏB�p�be"OB-�$�g�z���d6��E��"O���T��o-rTڷ	#�(tɓ"O�P�ê�<8BR��2Ń^��d �"O� p����nj ib&�3E�8�"O���>[)�-+�U�7C,�zU"O��QS�`�C��*u�{$"O����Ѩx�΀q��0SA"O�����
<0�)d��.r��V"O�Y� �U��Y�d�*{Ԃ��"OV���n��ܑ��ed��k�"OD�G�h�} wȲURY��"OViP��]乻�/ԾWP�0R"O�tg�[-��h�vO׆05R���<�'M8@�iS�� fRNt���t�<ɓ�
>r�^�F�A%3�`���Nl�<��B!�N�{eE9�M�d��o�<e� !�Le#�a�#��0Z��S�<���۵H=�Tɐ'� �Q �MI�<u�LOiT[������2!�m�<�O�M LPqE�
X����*�p�<���=U��D
C.��M��,�&Jh�<��A�k�����F
^0�p*��j�<9�M_2HJ�zw�Y�~v�O�e�<1a���U��'Ŀ`�ց���H�<q�2|pT �˵IS�m��B�D�<�ģ�h' Dc��T�\����IC�<)$h�J��Т!A�
����f�<�1%k�^Q�3�T�q������c�<����fQ���4䉎8ކ��f�J_�< K�E��{��=:�"��!a~�<q���r�t��i[yw�uj3f�<I4�V�L2�j�'��x"��p&�Xu�<��G�5 b�$�L>Z3\��3�l�<iB��4w����Dm��8\ ��m�<��%��#�d�(�Kl������V�<9dkM��c�G]�J��8 ��TW�<�� �&Z��	Q
Nd砱c���W�<)�(�p�ʽi�f��ʬ}�SFN�<�TG#0�h -�>W��Ŋ��D�<yd��Q��n�~����Vz�<��K�j��0+�k׵fbj����Hp�<���M lK4�ԛ6EL����m�<��J7J�F�0��bY��c�n�<��!�{U�zgmF	)�h4i fb�<�"��]eE���E�P��^�<y�e�r* ��b�	7�=
֢�8�y���`�l��)
&N��zF����yB�Z��A!c�F�A~`�����y�BB�<�8��PF�C����;�y��ڎ*eV5!���89X[e*܏�y��ʍ1x��`���0�.�A!�P�y�#4��3��D�3���a�L���y�#ת'\u� �	4�Ld��Ň�y�L�)Q���� 8K�]`���yR�Ջ�E�'P� �"!�%���y�l]�� �H5(�"��%��$�yB�'z�rm VM ����i��y2N@�P�<�1���t&b4C�+�1�y��~t���&uq��s�Ъ�y�MQ
�a[�柈�Bd��C�	�y2 ��o"�-;5L���'���y"z�N���[gx��v�ٴ�y���T��p�c/�'��x&��8�y��T*>i��"U+�T�b�_��yr+ڧ"f��
�j�DPɚ��y�`W�+�U���^�u�f��E��y�+�tk�y��U
m��]Z��y
�  ���T�^��b�B��X�"O6m;��rnM걍=���"O|�
�l��ވ������A�Z�2t"OL<⦟�Q:lp�6�9�^%�"O@80q��H��[A�����`"OP�rp��:6 �A�:��Щ"O,�1�^�O��s3���rM
�"O�A�e\./ϲ��CE'W�[��"O.-"�CǛ ��aSM+d�x��"O�4��m.!�K��j�P�#�K��yrE�c�0��G��:���!�y2eD'_2�$'���T?H� ��Y��y+�'xPzp�1H�V~������!�y�Z� �A��E�]|q�3I���yҀ�� �<�c�:_5ش���y�$��+�~�bG�'[K���W�y2.{n`�󄃍Cf����;�y�`^�ecU�\M9\8 ��y"CE����G�νK��u�X'�y¡��Ar0ѪEn2L┠*U%���y��9MR��򬛱B}`Ͱ�'��y����{딌�eDD�Gr�Ԑ��Z��y"!H�Og�k�0"�����y
LHD� �kǥ14��7nH��y2	\5���iJ�/���OO�y2M�%D���#�\��^�p5�J��y�mL�J`x$�� ������y$w��5��m�9k5	&�y��]�[F��hC/�
ax@��!
0�y򋀇S��)��B)�D��+=�y�fۋl�i��	�al����	F��yr�83A)� i�l�7F�y��T�]V&��⃝�h6�թ��1�y�IYU�p��d��5t����m��y���GKPj�D��	� ��u�U�<!���y�r�	tB�.t�x��́`�<��8��=s4�*Z��+�	]_�<�L�`����2*Llw�U#��_�<�+�9t�~��	�p5sA��Z�<�BP�`Ɲ(Ge�_t9c�V�<�J8���3����^��|Z�Y�<���� t��s���xDVlk�BG{�<��Á�� Z7�Y9+�6��%��J�<��O(o\�p���]�dwP�6�UG�<�D lV*�pu+Ǣn�[ACE�<����>��F��>�z����n�<i�Kp�^40��&B���Mh�<��
��]1bH��b�9(vmATg L�<A��_)��h�'��0��$�#e�g�<iA���&���Ѓ-��y��,�u c�<!���$�:�(qMO%J+��!c��d�<����N���
U�ܚP}�P�e&D�\��B�}�&Dy­�.c�D(�@&8D��R%�#-�DA(ת**��CI$D��ۂ��Z�����K�jI��e�$D�����r�0-�J��p����2g<D��QF� zv�`��o���F#.D��7��/䶵��.U�a(Ȑ։8D�p٠k[yz� �lQ!v;���*D��`�I��B��qgI���l&D�ȃ��)5��g��]Ԯ@��.D������T�*Y�wj�>�^Y��h-D��F �1y!�Eɗ��3�a�+D��
 �Q����FS��&�+D�� ����B0��\� ��&��A�"O��E%JW�dL��c�H�@"O�̉�*N4���	�A>瀠�s"O\xe��.�e3V�S�E��$t"O�ȳc	<T��89�N�*X`5ʴ"Op}J[��%����]�R	�	�'9Ll�`�\:(�Ь9d՗w8ȸ�'5�����7V��K�Oݖ��	�'�F0
W_�$Ӣm9���D�z9H�'!�Dxr��$lN��j�7:��l��'�p3Kd�r�*2�'y8bX��')��H �:	D��Z�IZz���	�''�9I�ln\V<I��ҏ~�ꀑ�'@�,��ӫaL���DGړ8�Z͸�'��l����hRaM<
�&ݘs�;D�����#�l�Uȋ�-��	ڦm<D����N4A��24�<W�h�#�)D��s�`�Kz��P��`Jrȃ��+D��jd"%.�L��^8Z�:�n)D��b@әo�*a����ig�+D��U怖-=��;����c6���N+D���'M�ƙq|,�v�7D�<��	wp����:�Yq��5D���o��\0H� .��Ʃ6D���V��!b��� ��))�T���2D��SB$
.9k��:��btZ�<D�ı�
�����k`�$B0<�z�f,D�@�p*�-}��C�h�R{#-<D��KS �-��P�BMi�θ��.4D�8H� �D����BJ�3��ĺ5�/D�hѧU�]z����ۥo��#��*D��3���~�T��eJX��|k`�&D���ˑ�eF�ʥ9C
����B"D��H��������D�䑢ׁ7D�<��X����jBɐ}��+��4T�L��m�P��x�scߩe�:�C"OpQ����S�bɀ��_��9�"O��RSF�x��!�vaN�p���9"O�����s=���Ю���͒�"OV��2B�[g|8�m�r�V�K7"O�MrT����r-(`,�2�����"OT�k�K�L@Lј"뛏���qs"O�q	D��
��q�jX;j� L�"O��C��9��h`�
�Ve!3"OTً�LȲ3=h�q�
���H "O�; 읅I� ��$g@�1�N��S"O� 4�АX��e��P����"O����)�� 4��ec^���!C2D��BY�V"��[vBG�.t�qT�%D�j� �-�p����4TxH9:�'D��#b�t����DaϷS��1D���+
6G��  K)i�Y#�m3D�p��B��1�,�K7<%�E��!3D����+�9wz�-;NɡrStES#�:D����"߽�*�$Zn�z%�Э6D�`s�%��2�&� E��*�e)D��q�ʞ�\�����-����f%D��ؔ��8n�ZӃ�	I�>���I#D�,RDOOm�*}[�,��	G�-�#3D��goP�|��A�5���t����e *D����'�T��3kV�H@��q��(D�\�$D�_��`9j����	�4I0D�P�����pxr]57f����%D��P"�H�:K�@6��*����#D�� (p�P��94��(Uw�Y�"O|��!�mn��)2�'{h�Tʳ"O�]��F=5Ξ��E�8�5r�"O��!a��d����H��T���s�"O�)3U��W�ށ���m�~I�"O����n��EB���Fw�h)z�"O4aA�"�/���k�-[	�.T�b"O�4��˩>~�|��M�"��B"O�	���x�v !�	;3��"O�-� �A<l��Q	�6ɓ�"O�yA��_!6�� T
V}���"Oxd
DOI�[m,E�֣�#[�-��"O�Бg�Ŕa�j\��\�E8f�a�"O&I�"H�C>���0&Xq �"O�����Y��e���$uJ�0�"O�[3�GHZ1��Ȟ["�B�"O�m!�d��2��9�"&�=4�Kb"O�lv�N �����2.�<ۦ"O�E�o��E
��$�����"O4�c0�π�za8�	1.���(�*O�����¦7��Aٳ)�BGJ	�	�'�̓�
<��Y��(d�}��'ń��E`K@��kʴ�p:�'����+L�"�L�6bY�4�S�'��kc�����-��+�P���'w�`Z�����`�ށc���'c�=+po�"P���ĩ��� 	�'3�	p������y���P��'j�#G*�Z�Vm��+ƶT0�$J�'<���kC�S@��mS�����'��X&�_��i�]I�:XJD>D�Lb#Y�u���R�U��&�X�!�$�v�*�/].{��U���A�!��ʴ~dh�`e�-E�j����t!�$��V���A�׌hb�*� �=M!���d�v�6�_�C���y��"P0���)f��\�azR�.h���R�ĝj1�5�H���M�KH�*�Jء�3a��y�4�0|��� *=�p�A��53�d͐��)M<��c/�)��[�H<X�]�o>iȅI� C��U�$����0|
�e��
�1%�N?Tʡ�dBI�r����J|��T�z���z�E�=p�`Yi��
{ �?�~:�j��Is��ĥӕ5��!���N}-��.��O�>}��ޯ.��M���H�2�ܙ(Nb�B���e8�)�'12��qE��avzli%�m�X� #�	��0|��Z����Ł
��;�x�E�� �J|j�3U��	����[O��	 k_{�I#�� �?�'8 �ɳ
��`�8hV3."�'-��q �+`�b)0��Q���!H�fZ TF��i<U1��S7��\+v(W2h��ƶ|'�q����|>�xTϟ�a���<�T�5�:���zF	�?%>Q���_<w�n�R@c�:!�2`HS`U�<y�'5��R�O?Q��㟑7Z���E�j�)Eg]�<H8q�EyӢ,�S͠<I��O�?q��&�2".x�(n�acЯ�ܠSV�<y�-[�<E��lȹI���&k]��鹆n�8y΄��h�t�m��=֛6n�|���)�FKx�k�)D?"H��D�yF���$��44�N ��O��F�d�����0��;�,eo�����\k�F���S%A��Á�C�@�X����.��N��:���|��M�O�'+��q��c�,���K��U w�"���[�`q7^�@H˟��W��%�O�x�'b�0k���B�$>Ғ�S
�'�F��E\-��w⋕�e
�'�r0�'�C<X�p[@J� 4�Y��'@�D���4H�V��J¢Z����'$�<:d�Γ"Mr �dϞ5P���'Yng�ۂ;Ǝ��l�/\zq���� �3����^f8�0�bδ
��a�"O2�2�ʆ |�t8�H����R"O���U�/�N�*%U����"O��h4��+ ���tC��7(h�R�"OP�Я
�z��\�6�zT"Ot(��;'�H�R'+��%
���T"O4��K�,͙�L,��	�"O@�ۖ �(;1��Q�k@�@pl0ZF"OmKW��:s�f9��D��lL4:5"O �@��?"rX��a�KN��P"O�� 	*XU��"O2�֨��"Oh!s�/����(����6K|�a�"O��$�
l))Q��3qH�Q�6"O֨J��jԆ������;"O�p*�犣2��|��`Γ��3"O�y�@:>Β9�`�s�0=9 "OZ$c5�	��Ãi�= �4��"O�a-V�IT�)�*Z�rEK�"O>8����3C���$�Ϗ!˒�x"O��A�S}�
�#I�|��U��"OBՃ�� h�\�qc�/_�R,ؒ"O:�� �<{
8ia�&��~����D"O�A�b��g���ED'�,9)�"O��m�&+N4���b�+웢"Oڥ�
�xS�t�υ�-ȔL�t"ON�ڕ��#�|TA���z�b}�4"O���Rb˳u9V]�f�M2���Ȣ"O>*$*P�yu�([pč�Va;	�'��4n_E��1`ޒh����'#�8�".�!��$��EL�B>���'u��@��M���
u`�'�:T��'"H��jA�\P t�PvȮX�'�ԅY�`O>	�<H�c�
g�
�Z�'�☠�@�Z�s�E4[��{�'�P��ɐ�}h(�Lǉ@W�d��'E��z��P!l$HE�LpDb]�'�U�EF�9
��x��/�1bif�H	�'@�=H�OI6�H(Yg��8_�E`�'d%`���%bUdLj�O*X<X�'B��"b�?a�5���	�d|t��' -6�	�Ê$`rl]������'g�$���͍Lq�i��� |���'AL�0��ۼq�DH�P��)Ddh�'��xdG�}�h]��ۧu%����'
��A���Z�v�����5�,�
�'�x�QC���S1ҕ��II0&7*���'����`S�?.l�9�������'e�)V�!y��QN�.�)�'�d�c��+�� ���2
n�lX�'�(�J�k w&���7O����' �a��k�BH;�-�>;dx��'�͊ k	��@��P."�B�'BxU!��В;�0�1ÃB�R 4��'Ԟ��w�]�eo�<�� D�Ƽ��'���q�ȌB8�`�=$#�'͠M���� h@�`m5Zm��'y��	T,[�e�~hEG�3	 ���'���AT�Öq1��eɗ�8��;�'l�:��:c�ލK��W�^'di��'A���֛ ��}��I�8�(R�'W|��Pφ�Csνh��؟;@�D2�'Ė��VřX��u���>�� �
�'*��e^�h��I#�)8Un�a
�'8��(O��T$�#E@�P�	��� fM��nS&~�d��a��B�J�"O��:1��!,p���b�^�ZY�"OV���%�S�~HӑLJ�j�{"O�|�D�qLҌXdn^��V9Q"O�did�[�"D��,V�d��Ԫ�"Ol�R��hㄈ[@k��ȍ("O�`v�N.1X@ذċ"��l�2"O��%�B�V�(��T�g�d�p"OH�a��;0��b*�/P��U"O�س�W$�	౦Z�e�A��"O�;S��	!vX��JN�td,� �ybI�5�8�f��W;V쓒c�,�y��0Qe��!��F;C즬�� ��y����*ndxcd�U:q�T)!�*�y�䔻a	��#�o�l�,�F�%�y(�zH�@��C��b��E*�1�y�ǁ+Zx 3�HV2���+�!�y�A� 3�����N�}@hA%�T+�y�$Pp�C��(�Ѡ�(ی�yrm�\P+�$�1��Dڂ����y��� _#��1"'�A�jl���?�y����ⶇPm����W�Q�y2��M�@��ؕ��� $oʶ�y2m6L�>���!��6���2�yBH��ĳ4ÍQ���3i ��yr!ݚl�Ɣ��.�KB��	�/���y���"FT�YT��t¤p�"�7�y�o�*;��h��+f/`XR)�1�yb
+���r#�ҨT�Aw��yRj�����↳I0�u0��ʙ�y"ǅ���h�COY#sְ��w��y�Q3U�๣���eΜ�G�Z��yboU��*�st)��X���H�C̏�y)�=75�qjԒUs�A��y�9z胕�ڭMo�|���0�y������3Mwf� &n��y�ʆ�.��E�MI�v��L�y���[=6��0$�	�^E#�f��y�DĶw����2Qv��Q�5�y��Y:{ܞ��1�ȡV���c�J.�yB��'�4��aS�&� 2�B��y�/���bb�70OJ8�!��ybKQ	y�hP�&��,u|P�	-�y�ȮC�%�'m܉+��XѢ���y��^w��A॓/a C���'�y���E�e���W m� �Q�˹�y�6rx`��:~le��#�y¯ca���]��c�\e�!�'Q�C��N&!4��I�$ԁMJ6���'|�Xa�#��g0pP�B�5y~@��'��Q�u
)2DP���c�$U�
�'�:�X3�4'ڨ�+�W	S4F$
�'O�<�����-$K�	nh<�b��C�<�C��-x�IFkԯ.	2]*@A�<�2 �
�C,�?�*�!U��|�<�Ȝ2}n�Y襪ƬL(=�ĦWP�<�r�S�e��I#H,Q���%�D�<Q�g�(��8��^�M&2L���E�<��mH6m�� x�咊$H�Q�1�I]�<��	�'S� �)P��������C�<iW� ��r�q!E���ѠKV�<9P�׶eT
M�*�!k���jGb�S�<�U��) p�S���Hsl1��CV�<�Q��NwQj�B��U
c��V�<� :��\�.h���3��0Fy�A"O���c)��q���RC�́?>lqi�"Oн���	�`R����f&8�8""O��P��
&_F����d�0�6"O�Yh7�1 4�X!KB5x���$"OJ䀔fd�x����0Fhplq�"Oܔ�g�"#�EӲ��$:ڐ"O�q0Pg�F4J��b�ۿF�@4C�"Ol����Q�H��s��P��"O�Hy���(S8�ض��=BOn�RG"O��8%���l/�y��NO��ܲ"O��E��� �||!��R{|a�R"O���Å
�A:� �X�< �"O����ŀ=?� xEԷNA��J"O�I�b#�h��<�F%�<V��B"O��pCG5?D�y���/I.@��"O�P�DS�~��=��C��1�5 a"O|Qy��r���)��"'F0� p"OXI����-���"�Id^��CS"O�`�\�SH�#`�~Jh8y�"O-h"i	*^$q0nR5'��s"OTXK��,GMVU�'�)�"O@���e�.�q�!�Y22|�"O�%��A֨F ���UH�_b!�D���J�[�,��ɘv׿�!�ĉ�%�K�MU#�b������e!�d !��@Ģ 2�.��Ɉ(!��W
7��*���+����c�ܷf!�0@2Qy�o�+�H�hɑ.!��h�X�x����<=���H��!�2'�$��fڎ�4Y���b�!�$9
W�ܣ6Ȟ}}�����)Z!�dB1D��a9!���f�5�$� T!�$�3Ma0�\�D��)��X�0�!���#�J�3�D�8@w�1`cd��A!��&2J������0Y�T���J!�d��w�ơ�ÉA),>@��-G�[C!�5N��2�	γd$��F��!��9�8�a#Va6)n�k�!�dJ+KR����ꑠ)$xKĚ�1o!�

���i�x5�p����!�R���푔�L%;D�X��lC�'�!�$��A�ڬ�𢊧z5>����óA!�Z�wԶ��q,C!e%H�
4fQ4	2!�I�=z�Uadi.
pD	��ڐV�!���q��e��N��zSQ拐f�!��L!�h����:"�q�AJ�>!�W�!�����ٲ9��mc�s!�ϧn4�1�s�ϔ��qD����!�]t��E
.���G�
,�!�q|��f�*s��z��F�>m!��^�d���A�a��+�R��%C�!��a��E! 
Ĩ.����$��A�!���&k��II�Ô=*ڕ�f�ا>�!��Ϡ&�����@��ꡦ4c�!�D�V����`��w0s��ߖG�!�d�$�J)��� �[F���/3�!�d ���i��H�j,�B�O�tq!�&�{���,L�^p��I��P�!�$�D�>e2u�˲yY ���铢�!�D�aQ����OE�W�Шz�'�<ez!��M��r�牅��<�e�Ѩpa!�]�^t�H$�!i� �R�I�B6!���X���S"Ƒ���I��S�B!�� TՈ&�]2Xf�BV(�p|rY�`��&�F]��4�?yڴ_���Ou��S��'}b�'%�ϛ<�����ޜ'nLy23���><q���^���O*��OG�3��#W���F�qe,� ��<�L4���J�f���	(.|�˂x�Od��Y��F�b��Ⱥ�@��3�P�G������M딶i����|�����??p�c@ş�M��;`�RK�H��	uy�)�邷`��c�I��]����J�LqO��m��M�N>)4��zڴ�9�СY��@��,��rV���?�U��2:'�����?����?������O"6�E��&�����C8��r��M��;p�,R��ś�d6g��D�,1��k��1�	�k��)	�O�*����� �$�ly���a �p1Aυ�\����A){�M��#T%�O�M���6�"I��+W/ �����O���	/�M�ճi<2]�D��d�I;!��H��4vZ�aG�l�p�'�a}��@%
/P<�	�BG8`Y�q����Y%�Ě�)I�?}�'�8x[kk��l�D�B���' *x��s#+�;c�����O��� �@��(�ܴjMZ�'&Ծ�dz�#�r�f1BC�X�Mb�IBb�H;sR��<�5Ö�H┱*Q�U�] ��C)�"ň��M��)6��PG�(c��Kn���G�6�I%6N�񦥒v�ӳ%�ʨ1�I�h�4��.3_��?i������O�m�K�
_�@��,��H6V,)W`<$�h���$[C`U���� }V�3I���h�@���ܦq���ފ�M���?����Шt�����{�M e(�P�r����?���Z�v��v-�#1|����O�x�fM6�T�jЬ Yw�|���kAk5�46&�a`��È}B��pp�B��<6fЬԘ2X���N'J.�c�ƴb�X1��
 B�b�"�������l��l��ħ��ɇn�"�6O�1_P��Ո�6|��?A��hOwE�:{�-R��(����s� )�p=�Q�i�J6-�>�q,���AŐ _vl� ���^A���Ӯ�D�O��4���:��O��$�O�7�5�]���^�C�O� %�³��2k�F&ըF���y���:�~Y�O��4@�ռ����
%�&���#/�D8���F�z��4Q3L��B��J�)8�����Ow���n�N1����2�&�(�GV�5�|<��:�F�x�Z��O��H��I�1��Dc�E�,���;fA8Ŋ�߰?�4��H*�AR�WRRX�$	�G�d�OZAl���M{I~����4W�*Ѱ��6�萖b�s�81p5�'���@��o/��'���'��ɟ����U
AD��yDl�a/�7~N�X�E%0��:�J�j�� 9HYT���]���l��md��z�͔���$73��0m�Sz�k�� +0�6���?�W�i��"=�O<��eDI�<�{焛kA�53��_{ў"~���PK�q�u� 4?^ 
���BK%�M�M>�6�i���|�����a$B" :  ���!�?�f�i�7�vӊ���*ƲU;jE�E
	|<
�ط��Hy��'�O1�`6mH�� ��g��+/h� ��e M���p����!Ϝ�{��r�E�|`�
��ߦ��'jƸ!0 W�X���'��S�8xn0"x(af�2~0A��ި\d����?��ޏZ��k���
���a&���hqdS3�����(��!���!y+ܝ�.�/?6�'��d:��P�f��:0���`;�'b1&��O�U:$�k]�,�fj`�I<	$d��l��4C��&�'
��Li���q��DKr#6��$�7�$�Oh�=!�OJ��#�І �ra D,�� ��	��'�6��'�T;!l��Y�j����%���k�ݱ��������DC {�ro�l�'�v��b*P�U���2��Z��EMۦ�Mcv�� TN��"+O>#������[�F/&�U��H�$fT�AD�D9��Ȓi�ʅQ4�zB��%C�t�NP��̜U�*ܤ�t���U��ņD z�T�g�Jm��a���]�@6�My��#�?�}����lm��8|+Ǉ'c$��������(O>��%��C�S�?  �!�� �*�)� �+�	�w�>!ñiHr6��Od�n������?��O��!��B��>�B���U�,Ka��f ��*2��OV���ON�����;���?9�[�~��TnW	o���磊�Sb6��!�?M�M�r�ԾEL`�fa%~�|r�hW_�'Ȓyh���8�݀2�ɠXjf%��gY�8�𤝍"�V�C��Z�zʀ����!a�yBㄐ9rɲ��ڎc�B��R�*6	9��y��x��'���d�?��D��Ωq�`A�ݴI���0�O�k�,�El�t�΁�+�*���O�p�I�MS3�i��	C��Qڴ�?iߴw�����B����E���uIz�{��'@bE�9\���'I��u7�����V,�Lz���n�}J LV^9��,���I7,U�Y���wC8�QON� ���+�N)8D*��m����@0Ec��q̒J�vi��+�4o���`4ʓpF�����M��iۛ�%ɐQ,���%CS��qb��XY���?����d�j��-AW�K��Q шF��p?���E���&��h����$���(�+�M�;=}�[��BOR��M����?�(���".n��b�,U99CJ����ް9�J�7b@���	V�0���}yR�'&�<y�oN�u��>7|h����B�D�4�E�	1!6#�'R�Ђ��t� �0�4��C+|�ɀ)a����Φ�1��	m�y��̂�/�����I�(p���<\O�c�\
��ɽA4 �R�mQ�`F�A� ;O-o���MN<1a��7T��j�aNn(�e��3#R�'��'���H    ��#����{�"O����2�����V��8��M͟��Ix��A�'�h� ��O��D��tU �&�O����O��wYr5;@�'VF\ Z�R%4Ȝ�[�����f�O�0��ɢcl�<27p˧��tMéW�d��(���X�-��F\�aP�(��ܐ������GCӚP*�*P�L^�'(���a�0�P�� �M�˓�����/�yx�l�+�M���y�0���S�gyb�igހ)��^���p�+O�`Zt�+$���#mKFg:u"p��X�Ƞ��Ĳ���>�M� �is�i>���?��';��h��A�*Z��b�Ч$��A�C�X�{q��On��OT�B�s���?I���� B�	C	f��s�G�2�|;Fo��xr�E�H	;"�;�,[R��'��)"m�Sr����k���QLG`�8��������@E���t��4����>�&D6ll�qA�(�Q��2��O�'�ay���zD�e8������#˞�O�o���M�J>1���?�ݫ]���  �S̎1~B�7�X_�&�#��g�D ��dH�@;\��fL�Fo�� �J*M%Q����n�8Ī�K��	_��ڣ.2D�������9S�4�?�-O��?���~3�9��aQ�km���U��C�B�ɔ]�He�E��<X*�[q�#�L�-O��ĜӦMbٴ���V�z��m��nZ27)j4�K^�v��l���B�$[���?�bj���?���?�6n��?Q+OV6�X�i䰦���c����^@ayR		���x�j���$M���]Za牥|�3�`�vay���?YP�in���?U$ 	J-MX��堀͟��@�4��	4+Bu�s</�ę##cH��@@���<�%���-l|I�g�(�n��G`^Ǜ6�|�'!���'*4� ��k��OJ�$�O�Eϛ�v�Μ�s
-a�x��HWh�58P�J�����á�xib���4[Q����㎨ � x@�
�Ki�pH���Z�2��A�Wݞq�2�(}��p�֮ͳ(�Q�4��i�ON|o�1�M۴o�z�`��
�^E:��s�E\�8�6]���Ie�S��b�xq�ejO�l�0�`Ƙ0;� �������)�a�6���إ�Q-}jhK��� G�f�۴��D�>�^n��	|��H�6��汄qJv��>�iA�ե|��T���'b���!�X���E�,O"Ũ"�HE��+��V�n����xbf#'��e0*�?�ȟ����^�
�<�!u�>k4��Q�x� �?$�i��#}"]w�!
5瘗ZĄ]"�[����	ד��'T�R���a"�Ij2�֝a�hc
ǓS�s�nOb�X����Y���RF���<H:U%ğ,�	z�H�'fj�C� ���M�����m��lZt�<d�T����:�������v�.k����BѪah�8���'ߦ=��e���>�Y����O\�&�tʳJ�ON�lڗ�M����O܎��-B#�(C�X��5x�{��'�ayB��rl\��/b�I��8ӨO��$������4�ħ���Sm»/M�)��:2t��hӰ���O��ٙP	�`F��O��d�O��df��xhWr�l��)��vWX5��KS	���O�(6�/,O�![���	�V��W�I�+����O�#���'��@g2�3��N�O��e�q�� 6x�L����%bW��ܴ �	d�6�4� �g��<V|��X�*ŉ����CMi�H�HE{J~�C���E'�Tys�	e�t:ro�e��ܦ�Kش���|��'��D� 	�|��㛆V���hjĖ{~��-�O䄃��  �Dx��ğ\�?E���$�*]a6�7bȗ��S�j���	۟Jݴ����i���O´[��)#gH��[���q�'�\��Ox����Ozʧ.�<-J���?��4i�p(�W(IWb�ѷ�/1wx͒�M͈H�2V����v����3# ��ʑ�/,<jDZ`�	�McD#I�eV�UqC�T~���i�p(p�̮1��0��w�nѸܴG�����M��R����禕���ɍZmd�3cʆ;�=�2�1��ȟ�)��T�_`V��兝�:��$���I��M���is���+���G	Y�zT\3��DرxN>��S�?�\t   �A^���QDV�Ih�1���?a�~;������]$�,+r�J�^/�	�=��h囶Ik���:�Ig�� ��	��W�K!؝�"�M@�0�k���ɉ�(9������Iğ�����u�'���AJ�w Y儇�hְ�����>��$!d ���dч� ��ū�z��G&DK�	�QA�a�5�V����ܓU��.�HI�"���^/��-#?��Dצ�R��D�>qT	��|%Q��:31x������Io��h���Y���G�~�r�P�ܒ={f
�M��izɧ���O��'^��[' |  �r5�EO�ɉSe����$�7X�B���O,�D�O��ʑK�On���O���B�"7زT����K�J�1����� ��ÈIn��D�'f��sR�<ހ��ɭ@<
5�����p� �h�ͳK!tx37�>�'_�I,4�*�P���+���E�ذE`��1��bo�ϟ��'G�T>�j�NT4��0�dAݴ8��|I�n��D��	�u�W�>u��q�  0L���&7����4���-e�:���?����\�|�δ�SY%t�h��O�@����Cϟ��ןX��*�=aPpY�8dɶ���F�r���V�\�i��J�(b�-����-:��<�Q/+k~����`���C	ť��㦦�>x!�tgۥq]��Xc,���(�<��R矘�ܴJ�'��Sag�S���\I�������x�������鉸Imș8cf&%��C�Hճ<�������#�4�Ms�O1W�>cЊ��/��uB�fXN?�".��V�p|����4�f1o�n�It�V�����T�^�:q!ҕ*�ZI�o1[�`�B�kh����U���)�J�?�����A�;/`��c��5�<U�&���M�f���k>���Ğ�:�Ƞ�Ǚ}w�d#���\M���5�HADIk�)�*ᘐȕ��M� �C�8�4RK��l#|n:���˹���@� 3 ��c�П@�I@y��'0�O��N��-��ϗ�?v.�w�>*�,�Dy"�q�,�o�����4�?Q�'�u� Vm��B��M!$x�k�,���yub�d�I�Uڤ��hܟ���՟��I�u�'$�Fk5q#4���ʫ0�j�bdcJ�E��R4�͂_���r��N�t6N,sGK�6��MD�0��'������Z5`����!�=�n�*�4�I�cV*)pLQ��;��i�1-ǀ��`JA���v.���#��x3&��P�E�F�,��~��I�<N<y���?)�O�\b�I>���p����nM䐀�d,lO.�Ö���T<94,���X�"�R��M�v�iHɧ�d�O{�Ɍ*�����<u�V�4P��� �.I0~�z��	����I̟��EFȟ��Iៀ0���kD�`�)�2�t�E��7��a	5�	� A��H�ŃoN��:"�d�@�<ID�'�-A�k,&=H� f^m���7�̅>fe��T/<���	L�L��<��������|U΀hakQ-�I��K�" J�9�4�?�*Or��+��|�%lɻ��@'%^,��!9wEc�<�@�I^��P� �WvZX �/�"i�2�zӈ%l�~y�[s��7-�O����~ڗ!�}k�u���D��Y����}��Y��'r�'�*�$�'a�ݟ��O��)3�*E4h�Ɖ$�<陋�$G�u�r%�`�?i����/�7�jX����ߨM���	�E�h��XۦIC��TM�;Ri�7�U�q�2M��,H�~�'f��c��`���W�$���)$��3w`����Q�i{�4�M�b'I:2W���&X.����eFS|��O���?�D-�	�� �   ���bμ��k��G8!�"yU�}I�0n�"M@j۱&�!򤎛7�~u�5"^��iш�?q�!�� � ���$<�둄�#&���P"OJ|�׏�1C`t�(Ģ��?r��A��ȟ��ӽ��V�'����i��P��J�+eDVIq����ԀS��O�m��O,���O�`�,�>
(��Y�!�OZ��w2B���F.X^�ps����2pQ*������Y�ӡV�s�)��I�*κԩU�Սg�z���_L��	�a�z�'�l<��f��V�t�6�dgݥ� ��n3Ĝ�\�*f4���-����	c�Ş�����w+� `��E��2׎<\��~� t�h�[��r�,i�b���*D+��Jk�ʓ)y�xS&���?���	G9.���d{ӄE���~^~��qg��[�<d��G̟(ye�"W�HM�;Zѧ!W�L0�y����\���X��  D!�T�R��"c����V� ����	�bȊ
��hs�O�_t��8`��th�_��AJ����5��a�G����D�-�RAoӰ�m���G���m�*=�t��%'u��6�K��	�4E{ҕx��z�����R�$������O��nZ�M�L>1d��L+�A�ȅA�!!�T9Vjr����dҋ\�d�mZf�'U萦�Ɋ|1F8�#J�Pܢ�hڴ-�ƈ`���1D�0���"!���D4P�Ǘ@��I]E`!��
���W���D�q�V��b��"bɰY*c� �O\"Dcc��T���݅/Ѷ��f	�
e'$�å�J�Id^\p#Z����n�O�yI|�����	ڦ����>Et��ޮ~6��F)����IP���HO������/��h��΂�8*M1��OrlZ��M�����'����O��{���2��ƛ>8�`JĬ0 m����P4t����<����r_wir�'��ɋ;M� 9�(kT��I�(�	&�ܘ)�j'f �BT�c��<a�m"�����$F�fgܝ�'-C��D��n�>8�)Qg��|����(XĢ5A	'j	���%Z9�q�y��ۥ�M�W���L#��g�\e����2z��$/��O��d!��,�x!�� `����aP��TU�g͂IH<!ǌL>?����iλq���aa�Fs��٦ͨڴ��s���m�`��O47�"��PX1�ؠ�e�Dm͂A�*��	>2ږI�Iҟ��I�xd�O�:*��kIs��)	!� T����+��*��x��	�=�̀���&�	C�l��-�`M	�ɾ	��R��꺇��!ABX{���PM��
��Ǎ�(O~��T�'�D6�S�����a�@�S7�eC0�Q�3�L4!�,]h?)�����h�
e���2����1�<+Z6� ��'�-c�r]�EJ��68A�Ę�S3�����A!�<�#��b�ib�'��=`�	Ŧ�+���f`�� H�Z��`�%��;�?�V$�5�?�-OJ���|&�����>(K԰���
6�zy�e��>A��P'qP�0AE�v~���˚e��8
�*�$T������ڰ��	�U>�d�Ӏ�v���-dҁ���Su����揵�p<q��A�v��d��BO�M�6�`g.Q�Q���شV5����A�<�&ؘ1	�8�,�	 �<1�0��k�IpX���֊  	  ���x1rm
��@�=�����	c6؄ȓy[�œ#J�0U>��P�	L�\D�Q��YĔEP�K�z)�� �v�>��6|ֹ��
����D肉�d��zj���-�jf&���M^�( P�ȓ;�z!8aƄ�#�\3�!�W��P��N�Ҁp�܍��=�G��*��T��w��x�CO��"	{�&�a����ȓ`�x�Z�	!}�򤂷�wW� �ȓy�h<J���/
��a��D^m�ȓ]��4��%P�@���3&���J �iгۙ-�m�&o�rBцȓ,�jh��0K^����M ٜ�F|��'�8��������I�?Yoڡ=��@P�X�6��D�HRRZ�ZA��1��?��=���FC�
"��K���?��@�>L9�G�8�ԉh��@9	�`#?9����֨ɯh����˻k��@!	ߦ�d�g��3� }�����I���$����4�?aYwo|D�N�+3���It��'(���	�>$�E!4:��ہ'ɗrn��6�Ug�����4>
���a!'P�둉H)oT(��q�ҫ�򤓶��q!Bn�O6��|���Y:�?�4	7���KҘk d�0�)�OvN%�`�'��-�%�Hr�:�7�в> �D���^[T�xA�Y>]�;/��<JhM�m@8JA�12Eʀ�')t���]�{�h,wY�`��(:R�)�*��Xm�O����R�K��!��	5x���ʦa۴�?��醮B�x�g�4eu4A(�u��?���,�كk�>Řw�5V���fF�_Q��޴X���|��)������G�0ꦉ��e��&���'b�I;#�> ��4��OFX�U
��c$�@�r�L!�����iߒ�A��\|�4�T�a�&���?E�� ;%�f˓0�쥸e�D�1�ȁ��^)Zi@�̚�h��"0�X�̙����ӭ p"J֬���y��'k����2L/��X"5�}�'�4�������'��i��uJE�#��14�SA���2�'B��"ғ���W+� �n2�@f�@���Y��6�f����������?��s���P�r%r���-؂���hX/dd�[v͏hHr�'�B�';b�]֟��I韔�ǉ�/:qk�T��ִ�ѡ�D[�hZ��@Ո����"u��afL)Q�z�<	I��-���rp��hɸ�$���!@Q`�K5 -�H����Ag, �$�"�PsAdC]̓ �,n�M �)�O�H���c$
�L葚'�'��'��O�$�W�9�б�'$I������,2RC�)� �̃&,O����1I�+�����>!0�i}�6m�<!��7+���'R�iA���nI�(����iY�6��1�ON�f(�O��d�O�;Ș(|� E���U� 9�a`@�Ҹ}]��hN��DHQ�,<Ba �c��n�Q��+�h��=6��Ң��<��I!���Y\d3e�� ]}���,"P��FG�d8Q��B�C�O&mZ�M3��u�EK�pN�x�IF3ϸ\	�P��~��' �O�>�KI-x���'չr����%k7�O��D��%�$���� 6�ս����
��Q���'7�5At�n�����O˧	�5 ��M�d/ɿ{�J��F�0_6�@� M���N�Zs�U�X��j�L>i��3���'�Q�=�z�i�Ka}⌙�o�4T��� ���S�J�.��'T�
��,�����{K��3�e�I��M���)�'�����my���:И���,A|��xB�I�>�L��cCÆU�q�Uh�:`N�>��iJr6-!��4!j4��LH#��	2�*S9&�M������<9%�   ��禑�'���Y4*x�����O,�Wh�3��R����)zD&%y5�3�'�R%�`�"S�|�	U��� �8cd�҆hŽS~6yH�޺�HOPՐ�愇��2��ɇ-sW.!E+c*J�"��X�����C�O@�n��O�>�*�K�6���jB�'�����'C�{T�Tp1L+oЈ}H� ��`Hh`Y��6�O��nڇ�Mc�4�r����	�ʕt��u�Nq�O����O��O�c��   �9j�ΠE�X�"
��L��4F����I��M�d�i}b�s��>�`�(���	@�Q��`���O����-cS��! ��7<�1���x�qO�dW�YH�4��'��]w�4�(D7p@TAթ?X�EYsm�O��"$�^�!P��O�$�O��d������M�4����	�-C�A ��/IB�-׺9�a}�eO��JXjڊ�<�D��ˬ���ڏZ'�Y�& �?ay��& Ø!�&L�� ڊĺ�������	4an�Jv�@�Gz�[��Y��wh|��h������ð�$G{���M�'S&�KW�X�B�����P��t�ݴf�6�|�O����|r�i���{� ���oH����MCw�i������� �5��Vh����C�{ qO�d5,O�Kd/ՏVP�!�c	2/��(����� ��4?�F��DB�
n��@��^��xe�mXQ|�l��4�I��(�'/�z���ߟp��ğ��1dN�\�&��e�J�f,�? '*�@�T���ɱu�\ ���J�zI���2c�$Y��ЍFZ��Ս����]=/�R�~&���J<�^���H��$�<5���Ǳ<i�O��SX�L<�נ҇8r���.2�.U��Iܓ�hO�π �V(9\ⱹ��VϜ]B��>!��iTF7�2�4���ɡ>ل*!ZLxa���3v�(���|?A��O/�	 `  @�?4�A"O�qKU;���&��)0�"O�iQ�g���R�#CaԂ<d�b�"O�m�B�1"�P���3:[��js"O ���Z�H�X�Ѡ�N�TZ`��'"O6��FB�El<���O�/P��j�"O��Ѥ�.�AW�L�,F9P�"O�i5"ݰ_p��0��S�
ik�"ON<�q�ѢK�8�7���Q��ճB"O~��O�/Iu�����tʁ`V"O��7�ƙ~V�{�œucZIH�"O:)�DП:�F�p��C6ID@��"O�m�r)##�"��MK�9>i2b"O����N�Y\@��Dm�,	�&8��"O� a����gHr|����*"��y��"O�l1�W�袵W픁�"Ѻv"O>�10�.Is�Q�R��g��G"O�]规 �"�~�8t&؇}n���"O(9i �]�`�a�2��,��"Oލc��r�f(�#ɓ[��x�"O�-��'F)���R�E�l
""O� α�t$J�� �ufP�x�0ۂ"O�#NN�W�(���B��X1&"O|+�ņy߼��Ţզ]~��P""O�B"�	B�/~����f"O��aN.j��
�ˆK���d"O �3( �y.-b�A-��J6"O��"CN�%^<hRrn��.b"�X�"O ܐ7��X#�p+%��8]"݁"O�T����/S,F�p2=UOHK�"O�"�V�j�%��ĢL?�8Z�"O���Nй~Ŷ�!�#e8���v"O��GL�N��MQ�K$c� ��#"O����j	<)�̐`ê&F���SF"O��wnkoF<�Jҹy6^�F"O:b��ѓQ6b@q�/�k?�)�"O�ˤ��2�4����#n�(�"O�%p�Y2ZM��VT=��)*O�����ڔM��r�GtG^pr"O*�ɑbPw!��oż=a�8�"O�H���(nc84����qeV�)C"Ol�pV#�3H�
A8���2yC����"O���U��d��+ ̟�N(^���"O�T�&�����V�Y>"y�"O8@���8	���3�H�@ "OH����K}��4�1��R��@Q"OZ����I<�l	����7�� �"O���RY� �q��L"g3TȊ"O��X$P9ViA�Ά4z�^Ys$"O@��u  -��ͻ",�&�Pi��"O,��C5�@*2,͙6��-�"OL5R��^;j�N5��*�
�lK6"O�%�q�P�(���p�	0�=�B"Oꈃ���43��Ā�h_�Y�6A�"O@�y�Y�\?�̋ 脫�ԙ��"O`!�����VI�m��F���Z��V"OFdc��Z5e�����%J?��d(A"O�<��ꚞ%��A�吟`a�m��"O� @T`?
!��1{d\�"OV�6�W~����T|�f\�g"O����(6�z����ڣ7��9W"OLq�c���z 2q`���}6�a�"O6\�E��(�jL��b�	}�("�"O���m� @��W�'gޥ�e"Obh
��@0^��1@D�T���"O }Z�΃�q �3�F������"O��VKQr(ę���1�s"O�ahRa��q2ҧP6�E�t"O�5���Y|�Ľ���A�}�h-P%"O�����~,�Jr��Fi�g"O��Z�k�$�}c��� ��"O ��(S�-X��J�)s�RA��"O�(HF�կ}�,y!�J9�M1"O�����6O ����΍��<S"Or �2L2�$�h!�]�o��i�"O����D\�q�����-u��@��"O�-{f�Z�j_�!R��_6�LL��"O��xBo�1%$��!mW�%-He"O4����9)6�@�lI� f"Oh��B�#��E������v"O�����'�F٣)��S�p�w"Oʝ��,�����<�Z�"Ot��f�l4(5*����$���"O��r"����L�<0��Z�"O TZ��/@
���*��t��d
"O� Z�H���	.H�Ñ$+�ea"O�Is�̎�~���C����C{p�"Oʨz#�X��!ጳlx�Sa"O|�sq���g��e�W�ɫHs@T�"Oٰ�f�/_.�s�nܠ^a�ȣ�"Oę
mJ�L���p�&R���s"O���٥S�����9I8���"O*(�筐�mcU��o�NLXEY�"Oޠ �L�� �Rs@o
7
�j��"O��`S������.�8S"O�9���scR�c��ҐR�dA�"O�!�$I�)˲�Ѓ&| `�"O>�Q�-;:�1���G�aKd"O�X��`��� �Q�O�&��*e"On��Ô={�ab�n
�t
�Ԃ5"O�( �V�s�� �Э��r
���t"O0l(��X�7����%I/bѮ}�d"O2�������c�OD'S�P�"O�5�KW�D8�/�V�N�2"Ot�e� v�H9u$'&���"O��JfJ�*�8!��3l�bM0"O����m,[���G��y�lQ�"OjEr�Ú:�����س*���"O�QW�|d�r���M<�� "O��J�bR�@��B7�T�#_�9��"O"U���0qRzY*���;��`��"O\Q�J��_8��ԫ_:W��S!"O�]q�h��4x�h#��I�t�t"OB�cr�߸Qy���-ц�(��'"OV�ـ�� <�EY���*(��<�"O9��\=(y�0��Cm�n`�"OHa"��D�
�� Ͼ+dxq�g"O�o��te9VIT��"�3�"O�	��E184R	��_/��%S�"O\��w
K%�8��'��~���[$"O������_��%a��I�3���� "O�e��9�2�*ԁW�6@Hw"O�$sB����>U14�©0�n��E"O8�Җcֱ)?~q6Ü�A��-�t"O�PQHkl 2voYT��H`"OJ���9!&=���'�H��Q"O�0�E�V�2DHA�nV�(8j�S6"O��Ș���i��,��4�$*%"O��I�������s��&l���"O\�'��*q�,d;�)ҸR�dm�D"O�!�b֑B���)����s�"O�Qi FߤC�����)�x�av"O�����HJ ��ȖD��U�"O�\�c �o��qi��s�z�9�"O&D�w�O5J�t2WǄ%�+1�y�L;L_f���Y'4^r�z�(���y�ǈ�cE�!C$�ڥW�b� �H���y�b_�z��+N�K��\�T�Z%�y�l��|3Ҽ���M�v��L��yrA֟+21��)T�@���zd.D�ybC�[���'!<6���o׍�y�J�!.J��j rs��2�y�/ھ#�4*�N�)@vЉ��G��y�mS�V�|���ݪB>����X�yB�O6jy�ٲu.�?,����,��Py2×���� &c�8�z��r�^�<a��Ր,.*H���#�$��c��Z�<��5�t��>ZSԬ�fbV�<�7�"D<R���f9U���S�UN�<� (���(ʝh�";s��hJl�@�"OH���+�?��ZsO�H�| 2"O^����
S.dc��b���"O�����%)�fms��?�0mi�"O�qb	K�M��5�������p"O��Hg�l���df��!^����"O���o�9 �2U��G�6Cd!t"O`��Tɻ.��$+��+-4���"OBlP�&O�`|���'Td����"O����ê
��I{$T	΂5ۅ"O��Dm
e=��Т�-.P��"O
��n�6!��1�'L�kKЕ�"O�ďV9������ ʕ!�"O�@悋2U�H����ըu"O �т��13��Д!?g )�"O� �֍Lp�Xr��
. hQ�"O���f\�� @��� :�"h%"O���nZ+t�z�:q��K�2�� "O���k[�-�sOΠjo��+7"O�DP�G�?8۞��NU�A��"O���+Y�R�܉E�B.7Z�1�"O�EǍ�s���BI?+@p8�"O�])`N�o�m��̗)(�$�"O�M�K�,t����E�#H���"O��!7���2�cǀ*R�a`@"O�`�S�C�+�NI��X(pFblr�"O$ň0
��rVVE�2N]+!� E��"O���d��9y,{�[v|FY� "O�MHǌ <
 {�͗x��ZR"O���Ø�?^��k�#��kB"O����H�b��pK�6�.��"O�x�D���eh��rh�"O8ҁ�ѐIZV�`0�Cg���+�"O����lӁ0���ZU��X�N%��"O8�G5e$*Ի�����A�"O��P���k?� C�C�"��A��"O�H��Ö U�T2�#�.���"O#�2P���h�'w2��"O2i�@� �O����&�9dV��1"OJU�cү!�L�u��9�13"OF��-J5a$��:e�K�,��L�"O����{| Dx���/R'�P��"OL�*���w�0P�W�G?�	)�"O�5��^�䝩'�I�b3�tB#"OB�2 �<&�*D��K�6F3Z�23"Oj�:Am�1l,�}�QJ��L�:̓"OFA`ɗ/9�X8�&S(.����"O�-H j��/�����Z�r��"Oh`�'(]�]��鰨 Fkj��p"OP�9s��@�ܕ��fic
M�2"O�H{�H!o�H���9nS�,��"Oi��F_�v�
��1{:��� "OdqC�23rdE�5o�7U$v�c�"Oj�!�&T�U^D��Ā12��j"O@]�RMZ-[W�Q�D 2^���a�"O�����W��IA�-Z�6���A%"O�v��D� �[x��	�"O�s�J�R��U�q�´��"O�ejèX�S\�b3NX(��"O ���N�6DJ]hC�B�*q��"O��p�R�\�H�t��;9޸���"O��r�䕅@{�����T'H=@�+d"OJI�4+�f2`PhQ
5��F"O8`Q��?D����A1h.�8"O� ���Ύy����O�3b��8�"O� ��*��
�Q�ѫ� "O0ܹ��y^B�,�zr%;G"O�ݒb��4%ȭ��j')���"O �R���`3���J6#߶�`�"O�Xp+M#_��C`KB�I�T	ڡ"O.l�ae.>�z	3bV�w��h�"O��51y��,� �X��.�3�"O`��D@�&r��§-j-�;!"O��)MX9yB.h��M�2;>vD�6�|��'I,5���L�L�\�(Q�œq,%r�'��m���G M�zA �� 	�H���'�,� �fGm��� gZ�z���'�Q� ��}�)@�R�%��!K
�'/0T��>x���W��ј	�'k$�8��@21p�h���T�� ���D8��0� �]�)�0W�Ŝu���ȓ ����οbU�9�2��#�v��ȓc�(��/�$�Z% TvD܄ȓ>�=����7<]0���u
e�ȓ[��;`�5�X	�%��6_=D�ȓ��]�#��c渡�u�[6y�l�� df�"gaI >%B���zɅ�M� �ԾeXPI�߄Z,|��,�\\J�$ţ2�!���{�FU��y:�t"���wpf���Ŀi���P�8�g�̕~�,hB�B&��T�ȓ-$ �ׅ~!��#a�
#L|Q��,>��2���@Z< C��ܕ D��TB�Z�㏟�5�KQN�Ն�X���� ��>h舕�Mǔ=b�q�ȓu�1����9s~fe��%Vp��ȓG�B	�a���0V2�t�ɓ2�Յ�z���)4"W=�H�q��A�&���Y��xS��,c��%��(Y�[����*����al����������v	2bE�`�:�&�_�>H$E��v{���׹e�l�jw�ďC�@���@<'��~2M�v��� �f�PdOM�<�d�'y�:�s�aM�;΄���n�B�<�Pd�݌�ۤl;A���	Mx�<����-$`C�]3T���)�Tu�<�We�=Q�[P�3sچ��@h�<y�m�2v��\ȧ�߮*��I�<�&��"uth��CE�q.v�RNY�<d� CHh�JA
�$4�Z���\�<Y���>ڠ\�ָBi|��g(�_�<�sM�_��9X"&��#AZ\�l�q�<a�GA:.C,V$3h�@�3�Nv�<�g��c̆m����_�`�3��s�<��C��v�́RȊ�O7��w��w�<1G.�Q���a�,#2�+bŎi�<�2��:M�Ԓu	��T��T@�g�<!d�\:%�|�BІޙ	n։@ ��z�<�ǄN_��9+��:n�E��j�v�<i��!8aQJ�)o
 H� �|�<�u���}�Z�X#��\�V�;ul�O�<�1��D
]0�eM�Ff�p�*�J�<Qg��o��C�>a�i�ʙF�<d�[�[�<\�c��9o&���F�<���.jΌ�Q#ϟ%�h08�W\�<�P��V骥ɧr �%EV�<14H
3�u�)�p\��ŧHG�<q#	�4r���ʶf�9hf�c�b�D�<� H���/82�|4�S�ѐZe"O<e�b��"��ǡ�	����W"O�$8"��\��)��݅5��1c"O�����@��*��Z�c�����"O�0��d��o��""�qb���"Ob��3C�Jh�����wi(��"O~:����%T����=~���E"O�T�v�#���&�Sgp��ؒ"O���&�Jј���ڿe�=��"O�§�3 q�A+��}�t��"O�sE�N�=r8���γV�h�"Of$S˹88�i�((M�8!��"O1SGh�+W��KA�Q*}P]�4"Oz����4yȇD��kaNɫ7"O���.�'o��ܲFN�@�"O�a��P�5Z��8~�]�s"O x"�M8+{�'���,��C"O��7E(��R�X�sX���"O��	b�M:jq �ıTq��h1"O�8!Æ�������C*rR0,y"O@)u"��q2-��.\qa"O	�׃˪��1�&Z�'�^<��"O�ݰD�÷.���F�0s��,�B"O��A�^�P1���]4N�8��a"O��c@��\M�0��/Vv�h�"O"0kQ�Ͷ>�1d V�t�@�q"O�uh�B��� `� G��A)�"OR��d�DJ��`nÜY�4z�"O6�C�Nz����޵d�8<K#�'�R�'�B�'#��E
�-��ix��q���"O��Ƥd��U�0i�H�"O@���m�8Nd+�*?��ŹV"O�2��9w�V4Q�Ʌb�,��"O"�@�����z��A��s����"O����Ƀ{�̡�* �Dhi�"OZyS`HģBL���q%͌�ڤ�'d�W���I�O�^Ո֮S
4�L�A���k0q��lPTm0t��(#��P����r�e�<���7d�j��摞[l���]i�<�1O�Ak�Hq�K AT� ��b�<	Q�	�J�Q�ş�%yi����^�<1B3^ ��c��e(J9Kv�^�<1D�X1��Y�PB�%�X�P��]b�<�C�e7�Ғ昼yN��rK@a�<A��2RX�h`#��;\D"�k�)IX�<Q�\57��p���� �2`��BZ�<��@�'��|2Cؾ�}K��W�<AkʦAO��+�g׸��93!gQQ�<Q��K�����Aԭ�W��R�<���5%�B�%؍7�JD�gz�<I�%| D}�@aH.0�2�2�[�<a�!SO�����S$�\�a� ]�<�qM��"t���t�_�5��*��Y�<�B�^'�2D�J@��>q��/M�<�"��,B蔉�tF3CAN�E��J�<����76�)�hI�#�^
W��D�<Q�d�	��`�ɇ/~[\	BnTC�<�+@�e�x�a�&���L�!��D�<Yt(�+f�	�J'��"B
}�<��˲��g�Jlg����Cm�<p�Q���a��M��mP�R�<Y�cH�c�~Y��jX/=o�Ԙ'�t�<�7��!m�RG�-#�^e��	]W�<�rbJ#+�p��D/ �m�8&g@i��S�? ����#zI�`��k�3��|�&"O�L�֌�3\C��S�hG%�V��"O�$xE�9JdH����#_��"O��2wR.a��fK�<�R$��"O>!�UI��Vˍ/B�P)�"O�ȁd*��(��ɹ'�{Z2�K�"O�)엱����4�� �N�"O2��ìL6Ȗ����6O���rr"OP:�۰���se�@����"O�ZV���|��QRPb� k�.)P�"O��7��>aYze����;�$��"Od��F�:�̐���o����`"O�zc#QJ^V8��`O�ߴ�h"O=2`nI�%|�Y@��Y�.�aP"ON� �k��_rb�� ���y����"OFT ���*V�`<sv ���"O�5
�M����N]��"O�I����5;Ȕ�3*�@:��2"O|���(ՔC.�e�b�hSڵ�v"O�K�G�Q�B�)�K���QW"O&����߁tt�A��
�2� �p"O�Y�P�P�q�ı5AJ낇��
!�E�!�l4���\������-�!��3{�j�I��Ƥ3���:De�!?�!�D�{e\8˶cq���1���z�!�$ �l�d�_n��S#���!���	Cu��3Ǝ�5U[Υ[Gc(�!򄒑�`pOXp����!�'ee!�-N�Ds�G	��|z�g��"'!�� d��<�$�3sX�d�!�$�{p~9�b�?w�E��%��Pybg�	�
�˓�M4q��3E#,�y�'J�%U���!�σ]�I��L��y��8Ca �j�m�1X����c$���y"��5�"�!0�T#p��s�̐�yBl�1����Ae�\t��2����y�F��q����΁!78�1#A���y�I�W�έ�@ķc�= Kˣ�yX!	��dQ'� �XR�M�D���y���P#�k�5VyX�
�L��y����Q؇��E��!�w"5�y�b��5ͨ�;�05�\��w��y�E�=%�*5[��)�<���Ӳ�y���;PϤA�H҅$3V�+�G4�y�c�9E���i�0|lq���-�y�i_"V�Å�@Z��# m_��yr/b؀BP��4C��k��ڜ�y�A�[���[3&h�p��@�.�y�"v�yȵ�� M2��U.���y�n[e���	
ݤݘ�$Υ�y"a	�-/2��1��bg8 i�
�y�N��,�^�����=U:���Я�>�y��$'*�k�e�>In���j_�y"�u�K^<A_�1�0�=}�J�;�'3&]�����c"BUz�B]�b&���'�~Y2�8h����@X#,+$!��'�nDPB��-�ʑ�V���,��P�'�x ��6T�eF�_*8=��C�'vꥩ��ߝ�L�%`[+*{䬑�'����1�z40��FGSwZ���'5��c��#���׉1DK�Ш�'tf<ȑH�
μ,X'�A(D���'��aS�M�x�d��?@���'�0�jEmYV���i2;�&�P
��� �������D��Iv�E��ZF"O~��A�	I��:�`B]<|��7"O]ӧbs���
�&ЙQC�4�'"O*�sQLG�.4��Vk�d)��җ"O�}�t��JHl�a�ϊe�X�Q6"OH(ǫSP�I����g�	b�"OZ!�p�U�j�y۠��	q��"OP�:0a��p���X��r�u�"O<�⡛syl�jT�Ͼ/[��c"O�؊W��3����ͧp�NĂ�"O��� ��9Y��`����%�"O����f5&Mr� !�P�b�*��"O�1��A� z�����Z&Mr�"O�t�G�-8°@:�T7MD��"O���7�)m��l1�Z�]I��`"O&��t)��J�p��d"B�m6����"O^u���D�``:a˖#$�6���"O]�[�sX*�A��Q�����"OX|�J�9J���iTo�$~���A�"Ol��֊j�*��0��+1�X��"O̝a'#�tw���6hŉb��AE"O&]�R����-z�� �F�e"O⍂�(L+O�r�S0�F�k��z"OF	�2B[8ؠ��&҉4��X�"O�K���tn�$@PvL���"O% !`�*.f|UkW�	=9t ��"O^��"^<��Y{p&�6/L�!�"O����l�>~�����E� s9�q��"Od�pϯ3�2�r�Y!. �z`"Orܪ ��;b} ����4�X��"O������>7V|pU��2Jr�q�3"O������;ͤ�[�/IA��x97"O|���Z�`V��
���-|�j��"O�]2�������)�l��F�ȗ"O�$#�A�W����V��8ca���"O�L���
�
2�dk&b�%X��"O:��-D�5��,��U�rU����"O��!᜷!��!"�0,-ҍ�b"Or%kf�({G�<�@Y�j���22"O�d�C(�9!
�m���pҧ<D�<�w�V%>�f��b�C��q�9D�d9��	w^|a���&�Ȩ*E�!D��q���$:���\7o2�`3u�<D����D�:A�x��X�X��\�e�6D����B�?m (G(�/W����0D�H��Mܹ �TаrV�x6b����2D��9c�-s�0�XuȜg�2$�0D��8D�!h����-�8Q��H8�L:D�����RM`r�"�C0vؾ�+V�+D�耳��
�ּH�OԬ@�D���3D�l��l�({��@��J��%=4���2D�;/8H�n-�Vǌ�[Z�|ۅ1D�P��X����$W�ʴ�0D�$�C�ڳRr���6m��%9D�����5	�n�OZ� ��Xc��5D� �d��T.��Q���hՀ�rI'D��ba�]2���7Vc�v��#)D�S���R���a 8&4JH�$�%D��H(�}�z՘��
��*��B�#D���EkJ �@�ˆ�)bHzu�4D�@�%(�9�p4�ZC��Y��1D�|���܅|�0�!ʜz�h��2h2D�`��O+v��@����XnQ���.D����\0�8YfJ��IIM�U)D�� ��S-J<Pi��wky���90"O����cVՄE�v�X�)����a"O<5�2�y��M��ĞL} $B"O�ZF�4y&m��� K>�蒡"O��"	�'G�((�)*m*B�ҧ"O����)ƭUz� X��O�ch�%"O�`��ٟR���aBťv�X �"OFД������b!ĥ6��`��"O�JPμXU�#â��Qn�M�t"OJ�H��ڭ��Ơ׍Ag0�� "O���j
�49r�o�8*@*R"O��P�T�`Q���&
ź�"O�Hڢ/��?�Ʃ�0lLt��x�"O�ek���.+F\!��ꈚ:p@ 	"O�$�A�J9X�X���d��H0"Ot� eI4Z�+V+X'G��9�a"O�M�q��kb@�u�J6X5�k"O���@_�/0 ��W�E,2hs�"Op��ቓCv��S��%O�X:�"ON=i��\�p�b�=1�<��"O�m�0,N�=!0h���MJ�\J�"O֩�%�1'� ��B/M@in�h�"O�����'P}P�v��"\�y2"O>��6�]�v��'� @=����"O����J<I(��0ч�|��"O"a���?b3�uzd�<v�4ʂ"O���pbɄd� ���G���[`"OX��O�8����C���|�l!�"Oz�K+�Z�2-��M0C��A`"O$�A�S�-j�����	�X��1�'�0���ʂu���&�"�(�h�'֚5�a�ѝ,�4iBw@�D.���'Ƽ ' ܾ:��X!�k�(|�\���'�0Y�,�X&��a.�?	w����'���PR"��lW�q���(@�'���NNLJ!P��*MX,��'�(�2�,��~����!�Y[����'��)���3<�	bDK!@|I�'�a���')(��8aă;�DA�'���jУ��.�Z K0a�8!�'�"\�����>��b�ÞQIXm����Q.|������U�����Y��y��O�&�ڢ �J��=����y"�ۭ^��P�.=C\ (�jǦ�y�m��v`p�:�Ƌ0j���20Nȷ�y��Џ%�tñ솟c�xD�7�Κ�y����d#�|���çD0h�C �y2mǗ���vg]�:����(� �y��/(����Cb�*Rƭ����y��'\D���e3&�k%����y�NB�N��ذ��[�  �k� :�y�͋N��8�u�k\b�'�?�y�J�� �h�����k}�@81""�y��M*��4��Lk\];�jB��yb��*.ԬA���<pd�'�y�A(}>�%����dd�H\�y��&D�WAG����3�bM�y2��Z"��dJ�J��4�D���yB�P�d�Q��G�>�J(�&�U��y£D����P g
6o(HyV���yR��2#`Tq∞�|p����y�,�V,K��x�NM�@��yR��3g���&�ׂC\^��b	��yr"^$�l\X"�)�Qg�U6�y
� jq��mG�!��t�u��'~AP�""O4��D��'���C�'v�T��"O�PH#O��hX����9T�L�6"O~U@�@��S�T	1'	F����"O�Q�@��r�� ��	/΀	@�"OvS%�j#�x�5�JQ�"O0� ���h'R呂f#K�J!�"O�Ԏ�i�@�P�X���7"OM�̓7��@nܜ-�Xy5"Ox�P�!ļN�`�e���
�4]q"O���BH�9�Kݳ�����"O*���F� ,#"R�@�<|�F"O�dAI^Ge��.W����"OM�#�	}�J�Z!�4:�`x�"Oj)�`Y%p����S�����"OZ�; �X�46��SDIߎ�a"O�YR 4޸�
�b� zw`��"O��2�	T�^��hp.��"O�l2P�K>�����	ӿ/5�P��"O�|qLթ��T !&ȘvI��"O�rdj����%R;/2�`'"Ot P���|)� 9�!��u�@�W"O�́d����PF�!:���rA"O�� ��Ya�v�y#jڅe뀭	"O���UG�/WxBPz6g��7��Q#"O4�	#$ì@�-4'�����Av"O����(�p�-	G��Y�°2"O`¥C��jm�E�Yi�`0g"O���g٩`�2��D�҄o�L�E"O�`T�J}�|�K�f�,D�x"O�3��.YjAsF��"{�&%q"O�mb�d�llЩ���9@�Zm��"OB���ר3��t#'GP�$�
\��"O�x`��"6-hQcA�	!m.8QA"O.�����__T��P��K�f�q"Oµ�AfR�xrz��d�ş2�t��"O&@[c�O'�tXi�&2�p�2�"O} �5,pթե����h�"O�� b�Äa��8:��=@BDh��"O���	�&6�P�#Z4R/0u"O�2O��Z"�CT�$3%���"O�B���஘�g���xœ�"O����ȳv�T�z�ťY<L�"O5x c׸Gu(��升:9��#"O��Q��8<T�e��F�2#��"O �0�%;��A�G���}
$�c�"O�hҤP�C��(���N�4qY�"O��Q����R�B�2�Lݱ���Ҷ"O����,T��i����Tyj��3"OQ8�n+=�v����Tx��!�"O�}b )U;p���jc�ؙƕ�k�l�<9��������XvU#�H@b�<Au �+q��TC�^ز��X�<!�G�h��: #D�-���B !MU�<ၥKF��ȗ�΁$t�a�֦�i�<I�Е��c���("|$�b��J�<���G<�t�k!��|V<��E$H�<i��=��"��¤b#<y�rH�<Ѣ��.�f����ˣw��ւ|�<�t�=*�dA�҄��e�h�p�b�@�<	C�W�{X�3��J��
t�qČ{�<م�B)X;�8j�Ϛz��]�gy�<!e菳e�V]ʅĒg..I(�FWx�<����h����
�p}�T�^~�<� �A��88~V�s@�������"O�W�˦Z��2�+�>dn��"�"O��d�݈D�������X[0��"O����_�dv�=��f\
,?���V"O�hQR��~���5�]�Hp�-!�D�6d6ĚE��!0P���f,�Mo!�$��\ ���$��'%���a],l!�9�����-kZy��!�p��B�I�m+��¤B��c<�4`���B�	�O�<� ��{U�ܚ!�Xz�B�I�F�J��/��LkP���r�dB�	�b��u&�cW�졓��s�C�I��
)��D%6��z�ʨ?�TC��T})E�S.K@d�t!0V��C�I>r��f��3	�Ԁ�v��/a"B�ɻbl��E�� V��ъ�s]�C�ɯF] �!����ࣦd�O�nB�Iy��7*��'��pb��Q 5�ZB�I#_���Jg�	#dzH��l�pnC�I�V�l[�+?Cv�){Ǣ�I�C�I�"b�������fal}R$L
8��B��,f
��.�*p�ř#l����B�3F�Ys��ͽp&d�za���C�	�Ku��+��C�B���B�	'u[8��dO�	.�����c�6B�	�tlb�d�	���жN�S/�C�	�"�p!҉H�P���� �3_��C�I�_��BWK�,[K6��N)xخC�I�V�n)VOѶe����~�!�R7Z� �� ���?$(p���&�!�P��IlTl�4���'���30��5��X�S�?�f�(�'�b9)�+Q�T�>� E�;=���'.Դ:���M��$��k��D�ƥk�'��]1���N�L�����7�>�	�'�~-3�II�"༙
FCW:���'���t��)�t� �ąH�v��'S��PХK�~�8�)��/>6��'���q����|�h�$���\"�s�'�xzVD�K���r�#�\ZT	�'����ܑ/s��â� (��Q��'5��B�\/>PXp₏<&��;�'�$Yi���#Kڰ8��˚�,�'�6��N��C����Tܱ��'U~̺��U6t�1���F��L�
�'8l4	`���\�E�.;&f��	�'���Y���2Pp"5�V(����'��S��!sQ� ��E� �'��9A"��d�z�д㝿v��	s�'�H��4O�1�0���]71:h)�'��L�5J�=���/�`���
�' ��col[��[T�F+P����	�'}��@�l��^�F�a0gR���!
�'C�A�u�%\:0 �+|�
���'<� ����O��(WFR#v-r��'���	;9��y�f�<p�(\��'�&9��o�8LYbu��n&�8
�'/ P���F���1�.mМ �'��๵ UxB�����R�5�|IA�'h�1�0@��ب�Կv�B�S	�'�LЦ�S�Q"�����:��X8	�'ު�+7g®x6���ʕ1�f�;�'�����&�Q

I�
:�q�'Z<��ŝ�NѶ[w8wԐ��� �(����%�@�Ռ!hXR��"O����;]N4��a)OVN6�A7"O8h��FE�B�,�3E�ǔvH0xk�"O�5�2�Ѷ. Nu���Z� 6|̳!"O:5b1�L<<^���L�-&��"O0ےh� H �ꔌ�,A/Z�Ӣ"O��A�h��'�^� u��%y���"O\��7�Y�d�8�t�[�<`��f"O�uQ��	����
�fA!V��4:�"O>�j	D�"�j�N-3��2"O>M�W^:N`P�yP&��1pe"OXˢK�u`�IP'�і?��=""O��q��D�E�%��%��,p�4Z#"O��@ͣY��qi����!R����"Op�L?}- \�!@*�h�"O�ɺ���(u/zD����]`a�"OTpa� �	p���E%��\���&"O ��q�7ma#Θ	}�����"O��b�.}x�U*��_�x����"O��s��n�⸀��.�\]x�"O��i�c�I^Yj���a:2C"O-�����e\3[z�hڷ��3!�䎐c5ت��0L�֡#tO�l!�Hy�pX��'^7X꒹����]!��C�]� ��℗���0Y� ��!�ӯ�@�����<5�Q�P!�dC�F���G�$A2�y��%+!��}�Lm��ELG 9�2�
�PyR.L�:u�B' \�#�������yl�j4����Ā������y����O��4�5�Y�9�P�ް�yra��:z�D�% ڦyT*�d��yR�M�!OX=49Qn��t�!�dJ/P�ZEFQ�d��4
V�!��ԝI��e(���	4�I�3j�8S4!���& }Ѳ2G���z@r!IʲI!�$ M��P"����M�2g�*�!��v���6�*���(W?<<r��"O ���ʭ�Bp(�2v8��"O�9m�S�jTbqe* �CR"O�BE�P	L|,���L�6[�"O�l�`	D+�CD��AD�F"O���,2
4�Р���60yx�"O
�iA�U��\�#f����b�"O���d��l$;�+W�9�,��"O��8����Z���	��A�6L{�"OĠHp�Q}��PO\�?�\� �"OJ���A_<j��p1 D�6��-�"O"�)�	��+
�ؙgsT�!"O��b�΃��f@�Rm�3bO��0t"O��q�T�F�yB�a��8;�ɪ�"O4p�  ?��C���%/	0X��"Ox����ք?{���r	Vz�J��"O��7��"*Z�a$�=�8�[r"O�dCc�^�RĪ�i�gP�jy�4"O�����(�t�G/*c�Q��"OZ��	�h�d�q�oS�o_��F"Oy�D\�*������ A�*�"O^����I٠��%�۝2�& 0"O�\�g���-����;+ˠ S"O֌��͕�L�zX ���jR��"O����,v\�3�!��tb�B"O�Y��U56���H3��)
�4��"O�)�Э̢_���cfPy}8 *�"O� P��#�EȌQ� W����1"O�xA�Lֺ�֙�ᯄ]� [Q"O�%`\�8�r��֭O8g����"O�H� �q4 1���la��4"Ofw��?mX�UȇSR�@Z�"O��A��P��yb�Ɩ<�x�"O}�A�b�VY���[:Yy<  q"Od8�Mߓ���Ru�ωCt��Y"O<� �f�v�, �D5N���"O`��+>i�rE�5-_�T�M��	s�O:̈s��M�*���M2U[4��'pH�U��0�Eq�iY+ۜ�R�'h��@N�3��,��%�Z�R�'@�\�tF�;��M;�@_Oq�'G�`��bаt����'/ɉ����ߓ��'�Sg�\]�^�wJ �@����xr�F�G�Aѐ/��k������y�ʜE��TDk�,q����ѯ��y��֡D"��r���d1�ݲ�	V�y2蜱:�
�aV�δZY2\�T���y"�I(L�Cfh\�Wg���˞��ybjC3L�8ـ�־Z� Y*$��y�ȝn�w-�C.�= ����yF�41Pam��,J��j"�Y��y���2x��� �	�v����y�K�A�����	�pRf�;A%F��y�۔F�� ��J�|%|�R󭕂�y��� ��+L���Q+�����0>���#:�D�$�,c
V��A�k�<�Lۈ[�$3s-ĩ	�����
\�<YC���ҁ�O��wB(�s˝V�<��Eݜ5ҒI!���|m[c�KL�<�rD�%f00��g�� �+C�<9w��_&	�0ED��9��@{<���,�Z Ɖ0 �և�mN���'jў"|��NH"k$�4��B9�h)�k�G�<�� B 	�d}����d�(���]�<�A��1B.<p@��'����raM[�<)�cҟ;�<iql��L-�$ �]�<�Ad�Ѣp�GM	pU���W[�<i g�� ����1�Ul�[�Y��Hh�i��1c4��g�U�P�WWxrТ*Oޜ!���D�@18�D�b^��p3�׈/Mh��d$�	�vҤ�b4c�vm���tj�
W�FC�I�6(\��U��#p<���T�c;6c���'PP�OZ�X��R*�zr��@�P6� �ё"O�+q��
u d�C�cy!���	l���\G�@�:Q#�v̙H愈
 o!��4}��Cb����8��e�6k!�$�)� �#D$O�s�$�A�
ڋ/!򄍅v�997I��s���C�B]3"o!�DQ�l~�SS�K=s���@WMx_!�C7W����&�.=r�����Pyb�H?N��'��!	�fH�n�6�yR��L������K�<93��Y�y�c���U��NG�@[虁oB��yr��X������S>;Q��ʐl���y��ƍ��h㢯<H(�LJ,���y�N�a�����nT�B�jiؒ���yB��k�\��fS#5�X91A�\�yr�0
�(�O��< r�D�0�yR�
*�ZI@I�4q`�HxG ��y⍓�`�H�[�蓈h�LH+7&H �yrB�U+�0� ��J�xY�`���y
� �	����M.�͸�(�=j$�, w"O�#eɔ� �L[�m�"M,ءe"OD��a
�����6�ϸ0�q�"O��lL�(�F|c�jݟ:�m�P�/D�����J���a���4�ٔ�/D�L3G��nt�m)V�K"j �Ai��+D�����4C�$Ա�m�+`��
7A(D���ơ�"G�R��̈�x�V�'D��B���|-���G�#�d ��&D�D�� (ChT�{'˘��{�$D�<p�k
$i0 {�oʶ2R��%�!D�8��C@"G`&p���A#�}�� #D�А�
Zj�l�+�&=�b���-"D� �m�$%;�q�V�U J|$��n>D��+e��j�.T�Ť`A����$<D� ��J/<)��	G��y���4D��JBH�!Q&$a$�
j�\� s�0D����R���`dH_�(���.D�(��a��/�Q!����p��-D�p6-P�z2�)iZ"E\��t/7D���F��>u`���Ҹ5��SD?D�Lх��d�T$��D�'� %8� D�T���*>,j� 0` ���	3D����N�R��5ۃ ��㎰i�/D�\R��ʠ,6��I�Á�J'nD��,D��q�$ =XX\	�&�1q�2� �,%D�X3�䜄h��Q��
�-��hHs�"D�P��*�?^0�����!D�P0��E[4�)uJ�;{|����=D�D���ʸ&3nu� ġ
�<h��=D�hP���(� ��Af�[���ǀ6D� a�4�Pmk�2�CǍQ��ybAɭQ�c7�\C� �;���$�y"(�h��q ��6fP�e��y2&
*r�u�k04^Ą)�,P�yb*��&�2Pbv�Ĵ%���v*�1�y� \�'nF�[��E�nt�}��냲�y�Z�K�ͩE&ټ`9�P��ត�y�g�q�rD����U~��zt�y��F=~�^x0����"�0㓊K��y��T4M
� �P Y(0[����y�I���t��I�#����Q�y�!#J��p/�G�\�q�`^��yRʌ�x��ѣ� �9Q����#��y�"�-C�2A����:Hh�9�L��yBk���E2� �8�b1U�M��y��Y)�H�N�;f,Y��Ȍ�y2�I"�$�vI��|a1i4)���y��7|��1�T�jC�	h4���y"�ɷ�~h���3P!X�$�;�ycGd�*�;J�J,4��4�yR �1�f��g��xF�#�"�y�	k��𒅮O�x2�ǃW�y��ܙs8��ەC�С��Y��y�kV�$)��d �BxFՒ�к�y�CRDI�x��*Dx�a�'�K�y"OR�J9��c2�=Nf��*�Oӈ�y2)S81( ��e6I�x�3sU�y��ˤOS ,;�ā#`Q��FД�yC�3l��4Hdi�0#
dy�#]0�yBMlԜ�3��'h�#�l���yboٔSr�K5��  T��`�I)�y
:bU�H�AC�)�콛0���y��Y,��ؒ���x��`�GS8�y
� �Ĉ M0A���W��M�Z�H�"O�ЫVV��t@���|4މ
�"O���ٌTcq�Ӫ�+�@z"Ox0�T��:D[���Ѫ4~%�3�"O��[�#�̈ʡI��
<t�`"O��pr�ɛ�d���Gɺz�b�"O��Y5!L�a�<= AH��	/
�!�"OR���j�;~�VHz�-��A�-�"O
B����^S����B"�;IY!��I�@ �M�i1jh#��iF!�$���ؓ���v0����6!�$�:'��H�1$�6�ֵq5��%3R!��Ҷ���b�g@�u��d񱄎<;H!�Z�v�<Y���(JI�4�A�A$�!���iO�(�c+SrHxG�T�!�]>)s~Y�P�sN�P*0�4:�!�$������4��sA~��B�]�_d!��DE"~kS�	(攒Q}X!�˨(g&�ƍS<�)�1WH!�Db���@�a�{-�4	�-X�!�-+vp���w��hd`�6:�!�d-�d��n�/'6���M�Y�!�!3r���2%\�>!��
u�Ή;l!�d�9~�\B��Șp�n�q�u!�dC�FaP������,��s�!���%gݎ�s4H��G���S�A�'�!�D�?w�,C�O�)1�๩S��7-%!�٣'�d�)d�|��IaD�� e�!�Ʊ-�F%yeB&2��ۑЄd�!�$�c��ݐBQ�k*�y7�_V�!�$Cp3�̰w��.l�\��&��R[!�ݥ>��(�c�z����JT���$�זB�~��\�D=�|�3ak�4�ucM>�rU3�Z.Tt��{E�%D���G@�`؄�R	v�Ҁ �"D�<7!guԁY�.F/p��uj D�88Rh��A$�ĺĢ@� 59`d4D��[e%��V�p9��ŋ�Д�Cf!D�T�W��3H*���V�wd�4�`!D�<�!E�.R\0%	����6(�9{B(?D���үE=���9��O�k�ihB� D�|Q5X�z�*3�@��$����6?D���Í]�\r挋�N���.D�P���O�q3$��c���F00��@/;D�$[�g�\J)����$�Ԇ6D�̨��Pz��WG�i*xĪ6D�f�Ke"�u@	D�k�.PS!L>D�0��/uIr$���b�&��E�2D�:�
+�X�G�9mä,*H.D� v��� �X0%�ê?u�h�u�,D��Y���|�: c6�A ���f�,D� z�'F"0�&�hgC	��5C��*D�� ��^'p16C��c�RuPU�)D���@�	rޜP�4D�$K�4e�q:D�`�!�\X��!��f�m��;D����"c�
��J��089@�
=D��"d_�4�v'��=��a2�8D�2W�I�4��ۿ	��(��+D���b �"	)f4��m��XU�E+D�\ٴmڞ8DL�s�ًh�
�C��(D����,�/!�^�a��P�mF&)D� ��k�����D)N,�@���g�!0(_(K��̂Q.Tkx�x�6���k��[��	�q����e"lO8q�2`7�@�-�'jt% ��ާd��J-M�D#�f7��Ѵ�ǖ|aZ�2��Ʃ'Y���E�/-ML���g��_;����w61�� lۡ"�.xnZ���v�j�ѓ"O�@"e$a�.�z��G �~�[To�#V<U:FJB�
xX�뗻D�>��'� �:�J�vA�HkCU��1��'f�����:�����,����B� ���(^�?�4m���ݝ`/��F~"6��i:�A8R���
��<�Tj��r<���Mգ;whY�B*
�֬A��^0rg�AӊH?<�ޱ��,M��p?�fJ�=����Ao_�V�$�K�>�G��x�&Q�"ѵP�b�	P��<~�ػ��2j��H���z�ᗼ>��("��X_�<��͗+DHa�8i��}� ҚF�\�������!,��}b��ۑ����T�<|�$�*��!�b*M�|��B��U�:��B� �p���ɤ|���  �
�,`�K���2J��h�7��
����"�}�'�!1�D��b�����T���X
�'\��G���$�~�"W�En���`���v%Q7�L��T����	q ��aג��>�a!�u�2!z��W�ic�y���s~�,ׯ\���9s,�=b?:*nפ@�x��e��1��Vg:��C�HpR�bR&)%�C�	�Y���F&0I��s��@�$@푆HqtTZ3d��>�|<$ �P�Ӟ:�p(0d@n�M�"#R�0�]�G&ߢ�����h-�D�b��0 ǈ5
 � �8t���k8�@왡�@bQ�X�h��CH1��F{�h'e��4͆�|�(QueB��0<9c��j1�Ԩ�%�)-���a	�h��d 1�\�>TXD`K&-��I�v�����b�I�ӣM���C�!���� �mp�_*)᧎Z��jp��"S����S�{�����,+��d@@E�oS���m����C�({}Z!�c���V��=Ϣ��G��|��oV���L)xqBg��	`���%�>Ȳ��*W�:��5F*J��!
�P������)�D	��'ʔ-X��s�?f�����˕!��賆�!=ݢ��fY�tA�(I?h^�	��MZ=j���0o
���$�;Y����X��z4��+���D�Y�u���g��< ��}qT"L[�U(�+]9"DMse�\8����r!��S��55T����%s�]8'� ]�'x��Qc�v&�@@�1�X[�G7S����H�!�N
� s��	�ř�~(o�	4g�u����??l�$�P�n0�7(�-[�s���ir�Bo��T*�J�
	��ai�u������X�V���P� ̛V�?y�$*�"n���$�<9�5�Ӈ��a��T�
��t���[v�A+u�V����%ǘ5Q?DA���?�H�b�è
&d���Զ�������O<��PB<WR]k���<�D�Z��*/v�V�\��'l��e�s�
��00�����}L/h�0��V�b�up��)������=�xaQ��� v�9�(y��Rf
����X��8��82$lU�+l�������O���$L�dI3�Y�fv��Κ�O�i��A1��Z6�I�c��dܥO�pis�e~�4X��I�ԣ� �.RA(#�(h~p�K?il�
���^�b6�أzО��7�^�:�@�@	�-gA��׭�x*�u�C	Ԯ�D�2���zӈ���"��?�Nͮ1W�aWbOV=r�Q����/Bd�cE�'���X�E	�t�8J�Eac�P�Pn�`X"�w�6lx6
BAA�	##������ �h�/.����5B�8�I�Ui��Bs�Z�خ��m�R�Db�p��"�<O@�ڵ�ۆߤ���ڊP�N y�&I�IAB�A�iU�	�lZ&�B�8ᑕ&�VW�l���6��(:H@D}R��'K�t ��gZ�a���bQ��%
q�d�D�.s��Iƫ���T��&I�|���`���"��I�y�P��eE�:�V�!���JL|��@�XPUF��	E^��s�d���|h�/��U8���T0FK�uI�NG�J��8:��@�+�N);4D���`h���"Q��t�%����NR�BJ�2Ӏ�W�O��=9�ذy"� �T�J����1��K� 4��qWg����2JNB.��`@�<rz] ֋ϭ(�����:�Qg�b���.��؛������!MW�4��p�?a�F�,[
���ȭ4,tų�#Z�cb�����П~.R�v��0-&�+N�/��L�1bԱju�"���������5!D#?�a��1Od�R'B���Ǎ�9��Ƭv%�	�p�=<%~���n�0Lj�
��ځ ���s���a�J-jG
AǦ���;�D�D��ݪ�nZ��rA+
k2L3Ql1"�p���8*<���fC4�6B	�!l_����*
m>P�C0 �vλZ>X�'&}{����$Dp%�Ʌ�ƙ�g'����2K�ɀ���B�4�@RGfM.3�����l�!&D/�$�M�u&�q0���ib��C�Ly��kĈ[���Z�x�:�F{2��R]v����<�&����KUŜ�DM  �ϒV�E�d�[,<��I��@��B�LR$r�`����urbH�B�ZӦ����[S�d���ԒN>�cC����'��<��n��' �q�7k;ޱ1�hX;j��C�I�*$�V��l���b%�0n��e�qz&*�)�'XX���$	Vy�������1�ȓCt�JFԪg���PDk +����<At��+��<فe$i�U��.M�
!*����j�<�c�M�G�1����S8��@��r�<yN�fTɣ�K�7~b�%���@�<نfѦ9|)q%�sj����~�<� �`c-@:v��&�8�0س�"O���F�@/�
�h�K�I,�q��"O����I���A`&�'1�}PQ"O�)�QB^!k� أY�mNH�+1"O0d@���^������r4��F"O�dQC�L0�҄�%j4��"O�,z�h��l<ȔaB�S��z�"O��i҈�,R��#�@Ȁ���z�"O�D
d㘸G����ˠg��P��"O�x����,YoH���ΌC��q"O(D�f%K�T���̅�H�e"O�]������^�f�����/D�!��1="�"�dT 
<�@!�+U!�D��B��r�
6��Q�X�?G!���7���I �P'rA�D>@!�D�<%FJ;v/L �tуg�!��H�!��Y�˝ R�c��F	�!�D '﮸��D�+I:�!�*�f!�d#@Et�x��;L"~@z0',d!���U�p)ؖ�[7>��	�(K�4!�䂸]�,�Cw�����K�Y7!���� ;��V�b8�t��ɞ`�!�d��=-����#�	x'�L����9i�!��K�}�̅SE�M�!�|m�&�%]�!�d�]���⒂��%s@���λ!�d��^��I)�)H�]n�a��!h!�$�\��`�T�M�SD�<�t��x�!��>�ҭҲ�τ)����%�R94�!�S!�,��#E#w�&��I	��!���rq rv�-]�\̨TϚ i!�ԍs�����N��e�~ًt��
-e!���5S^��� ����(�Q�p�!�����7c٣m�p��{�<as�T8Q	|� 5�؟}�UE�H�<! CX���&�s}�db���]�<A�U�E��x1WMR�j��j��X�<!¯��l,��Z�oI�U!E��V�<��N�1B( m��*pA0-�{�<��)�0'B,� d�'f�>|)%��u�<���̩�U�/*�\Y�j	w�<i�/X�6gT$����0nv�����e�<I���!�l{�1i�0 �t�a�<��J1��P��m��	�N��Y�<�cg�=��}�)�>��a�q�V�<���F�ĄÔh�>?���B�K�S�<Aҥ v�e�C�A�?<�P�G��F�<�� ���`��;{��pI�C�<CL�<c,�`ׇ߫j>���SdV~�<!�@E�|a������i2"��v�s�<a7�*9*�a��;4K6mH��j�<ywL��(i��Cv[�b��=���`�<��
�7K�,��b��7:�4�#r��E�<�� |�Z�i�nH�]#�.ܹ)�B��'48��k4KP�*�T�B�!. �C�$W!>�3҂8:Z	��]3w�C�	�eΈ�(����p)�܃d���wE�C�I�j]b�� �
j%��21(̠��C�>c�ebv�M��z�,V9O�C�IF0�J3�ح5�=��l���XB�I-�ع�QLȿ"j���Ո�
_p�B�	�N.
$��*��e�d"v��,^C�I�1&ڼ�#
, 2iY�Ĕ{��B�ɖN5Z���n	Qr�HJ��D>~<�B�+e<V�b�q��)�smQ;|3hB�)� ��ᎀ�)����%o_hX�P�"O`-�e��(9�uQrϝpW̕�"Ob�($A§;��5����#[�`��"OƱ���bz�H� Ѱ9��0�A"On5P����ms�0cwoϸ<r���q"O�UV�߲;J��#�Lgb����"Of<�vE�)m��	
NAby��"Od���U�	^p��"�.?;օ�'"Oةis�wƬX���8���r"O�R�Ӣs��,bСb��4��"O�ؐ�"ϘQ*�醀�-��0#6"O8Pr!F�4+f�C��!��=(b"O��:�*Q2kz=�f�|^r�
"OQ�a@�$x�ع�؛*;��`"O�P(��+��D���Bx��!D��s�/��X��\� Y��;D�|+�N�;qߠ-��I`r�8�8D��
�LR9j`M�$��$fєA�6l D�t���+Mp�[�n>h�	��>D��*��߮z��訴e֫ky���a�<D���#��/mL��;e�#R�z�@�E&D���4�F%')�Q�b��n&TMbģ+D�����H%7��Q�L%Iҽ��#(D��3�џ
��ڴ�T�L{j�Qd!2D����
�r�R��3�t�B��$D�\:�Ț"
g�=�B���Z�.7D�|� �X�J&�|��^�7��ҊM�<��mI�`�������:3��3 ��c�<QQ�Ų��	�
1?XrLW`�<Gɍ +��	�D�8!�- amHE�<�q,�,y"L�f-#�2Qv�_|�<� J��*��(Y����cOz�<!)��=� ��X�
VH��-�~B�	 Z�`���,�T�&,'JyJB�Ɍ`NVlx"��\d��s�Y�^oNB�I�]��yR�K�^<����g�>0^,B��3TE�Ր���8��q��& B�I�S����@54�D�p�?a��C�I�wc�mieg�U��gA �C��5g����
�1��q3jɞ�͆ȓbrF8"֡�y̦�ZGk�a�&��ȓ-j�u�s�C���sf��p5�y�ȓ�L`zE��;v��Rkɀ�>$��3Ff��)�B��D X<RY��G`ԁh�2^q`I��VU��9��<�&,� i�XUhؐEX	��l�ȓL��=JL��j�l\Jd���a���Y�@K`膞]H�	Z�-�tߖ	�ȓŢ	�C�>5���!p�X� ��ąȓ4��XI��wJ&�歏S�ȓO����7M�Q�rQp�߁|�4��ȓ>$xl�������DF��ń����9'��.iY�T³g[ x|��*J�LJ��4��T2!A="���r�̡0�I�O8�@%%B4JU��=Vl��%��Q-`l@�`��$�z�ȓA�m&��5!� M2s�����jC�d�(G:��#�/>���G�*�D4O�җ��K��)�ȓ�LR�o�v��I�D#�Q�ȓ�>�I#�I��lAa��@�T5����rA㐧`�+p�ˈe~���S���8��NR���*�"wm
M���0��M�8'b*KćP�F���S�? �<1�~�,��(�!����"Oƙ�t'A7.'�(�� �E�`��"Ovq��ʃ&6����C�""�t�"O���t�^�q�4����!�=`"O�|p'�G�s����/>K ����"O� ������q�0��)r��"O��IOݶQ��͔�w[:aɅ"O6A�&d�"#��$�'3CFL��"O t2�*�7H�tx��ѭh8��+�"O� ��$�|�d�9��V%u��"Od!��Yg����ƚ��yb�"O����C�6�v%�����nŻv"O~xAdMZ3�0�1ChK8�ܜk"OR���)=��"dh�=U���0$"Ody8 O
,}+��xu�٤P�R\z�"O�\�"%��.3b��EG@�v��L��"O���+��`��j���"O{�ָ ���ӆ��z6�q�"O�A�4�#t�f Q�NQ�|��*%"O6�cad�v���%j��	&��r"O ȰbڣN����ՈśH��0�"OVܙvON�u>��C����6�,٢"O*�qO�t{xU�OC� 9`"O�uyU$є2f��r��
!o�P�B"OK�H>f)�Ȗ ~y���y���|���I���i@Zl`��X$�y2O()��p��ľf"�Y�E���yr�ηqzΙ1�Bڀkh���%܌�y�)Y,)�@}Z�m�1ZJ`ؠc�P��y�M[:�j�`���R�\�S�ʹ�y�i�1A* �(�W6�0x�O �yr'�6kTΙ#�A[�I��{����y����!Q>P2�#��?JсbX�y�,�&tK���	���,��܅ȓ(ˎ��K9'LT-X�O��f:Q��H�T�cFؒ$J����Z�/W�4�ȓZ>�5���T��F	#�� �d̈́ȓ1>P���|,��iĭ�9����"����p���6��)�\��Z!���$w���R��v�|�ȓ�0(�D��8lhp�54�H�ȓ9 �U{⚐>�*�`R��Wݰ\�ȓ6g�)b��N
I��R&��/�6��ȓl��t�BG;�����+�hKT��%��|2-՛=mn���*�����,b@�c!_�U�����%j�Č��Vq�MݸJU��'ɚS��\�ȓ�e����P@H�:�*JY����ȓ5$�����&hm�2��O٘���Q��a����9_W8�,��H"X���qe*��LŎ���yN�7i��ȓQ�l�saE�9|��Q`j�a؞���<p9�"S�}$�}��噡S����ȓU��`�sЀ�sFꋘ{�X�ȓ'�h��-'��{'g�|	PŇ�wN���A�ˆ����	)�PՇ��V�:r��+u�8$��
&����bWT�s�(��sv q��W�XU�ȓ��`�b'�$I���CAC�rd|��$�*�[qd�>P8�̨��!y���ȓR#t�Sfc4ct�)���U��m�ȓL�`�(5�ޏS� ���G����� ��¨Ŷ_��Q9�DW�R�<��Z�I�e�T����C�	��\��S�? x\���	B�Rƀ��3앙"O�����O"8��4Dď:6�z"O��;N�v>��9�C��<<&95"O��1Ƃ��D�W/Y#Ev^���"O���4.ԩjZθ�fH�.NhFaq"O��('J��U�l��s�C���0"Op�Y�Ov�1��<$NE�"O�E���Z�s��(KF��v>����"OTT�q%�M��iA$	�u	�8�"OT���OT�ZxS�	� �F���"Ote��g0PԒ�M� �&	9""O��#��/'���(Mv�=��"O&����_G8
�g�^d���R"O�A���;LĆy����i��T"O�ipQ�
�YX<��#�Ц`wx��"O����Y�b}� ��>�ށi�"O$YU�ќhV��ɴKWy��S@"Oj�3�)P�%\�H���`�ec"O|�;��3h	�D�@=�Z䠂"O�]1b@(��p�v#)g'�1C "O��ςpf
����Kt��"O��bZ�ZF�Չ'�ϗT-��"O�<B�#)�I��ӫ+�!�"O (S��R KH��-�G�Ҵ� "O�PQ*��җ���$��c"O�I�#���6�(��J�W�xMP"OlAㅃ
��0�`$d��|S�"O$���?jB-��CT�@0�`�'"O֝���
6,��N+V9��A�"O�R��ϔ<�`��+�6ܤ'"O��)�	�h|�*#�A�t�i�"O�e��M�� �5��Ѽ}�<��V"O2Փe�́q��=;�
U��$,�D"O��PhԺ8mXI2�����Y�E"O����B��U+W�����$"O�h@�/�R���y�jR��d��"O푇��q]V<@�J��v����"O2�P'C;>��x� ��� ��P�yb��*( b�8�"foC��y�mƩ_j��7j );��t9A���ybC�o㐴���1���30̇!�y"�H�Vv�P���҂7���2�Q0�yB��Y����M^��LA�)�y"c\hY��H�Y:����^��y2��zײ��	U�8Nx��'.�y�@�B������)ֲt��mE�y�j��>qP�W���zf���X��y�蘯y�f��B�L���Q$���yb�� `�(���ʕMJ2@�*Q%�y��C$t�2p�'�v�����͕�yV&���rc%Wn	~�ju
̽�y�) �RҴ0P��iJK$���y$�x�y�+��Ā��
���y�7v��[Qɗ
f��K��y��I�yL�:䈅"��H����3�yd�#�,�!�:�°ju�Ы�y2��=�d ըy�D�d勹�y"eܗ<�ʠ;�	�����@�y�)Q�|.�z)�Qc�!+C�ǯ�yRbĭ ތ��g��bX^m��ϟ�yr�ݳW��․ºd\zL%�yb��3�j���T�a�,��� �y�n�
IT8Lp�@�Y�-����.�y�Ͱor�=�n�[��)����y
� ,#a���9�I)�h�>�r��"O� q�dĮVT���'ʱG|���v"O>�h��l,���ĉ"�ʬa�"O��F��� ���s���vKL<��"ON��4�
#~":�c2<����"O��:���}x��2
&:c� �d"O$;�K�gH��C�ԐC��y�U"Oj�����13�;GE�8#��A�"O�x׉�=\�({�^5h��ě "O,��Ԧ�`b��D�	����Ȑ"O�a��k�*f�V�J@J��cz�e�s"O��b�/n6Mx��Џ3�l�Q�"Oڱ��[O���X�B�K�*P�"O\��<H��-�Q�7`�:��p"OT����"nB�o�/.��!��"O
�
�i��zņ9S��f- "O��zC����!qN��F�r2D"O��#G�2?�`TS�T<�0"O��	�gH[#T�I�OԦI����"O�@�c\�{b"��%h�l2�� �"Oa
��G�Gj��{��L�v���e"Otl�� ǊS���I�7v�T��"Od�%�.%qP�B%+B;l� �H"OL jMI7=��p䊓�W����"O�`��/S��K�'*c,izg"O���'FCG��lq���f}F,�r"OB�{�d@�Z8�T�t&G�m�y�W"O�	��F���B�R"*D8?g�`�d"ODp��&���c�IP>Eo~-�"O�uc�Ic^:	Y�JU�(�>�"ODA��!
��d������d�Q"O��a�Åi"�ĸ�cߝ3�<�{�"O�l��AR']�.�Pl�d�<x�"O�H�Q�!a~���
�?qhI��"O�����4�t�v�**�Zy��"O���ЌP��bqA���e_���g"O�)z�a��7��"��`r9�S"O���S�W�Q֠)Pc��cX��K�"O�5�&�n�̼�ଚ�25*��"O`H6���y4rX#
�Z���w�ɁƸ	��o��mZ�x��J�6�0�I1���Ùj2�Fm^�$�����:⟢~�GȐ�����e�<ps@R��Լ|�]�O�8�@O)��d���Nc?��gK�)�T�����T�r�c׻}�6$���l��,VN=��Ov@�ʠ�E�2,�҄-� 4%�qu'�OZ�!�⛠M�`HC���0|*�ۏ_^N̑���+�˵bĢ2h����ń�)|��!�0\*������|(g���_8p����5p����Ǣq�|�#���R�S{��@��bjyX��b�����n��F�� 6��%���#��K]��8�������M� ���튇a�����i� 9��)Y 5�Y� ��R���D��>y]w?�������cN�@����I�qI�C˹Y[�]1&�I}B�Z>���mǈT9��I#�Œ]W
m`'h �
�t�@�S��BHC�Aa�4dN_�N(�bC�e���S�@�yB��e��/7FS&	ގ8D�����|��G�v��3ĄV.0:|�`I;Iy�xhWP�CMj7-/.�k�'Z�VܹV K�,yT�Ӎ s���J�k�6�*s��rS1������r8�d�р|�\�`�d�C2�3� Ǔ�Px�d�jܜXYDg���������yb�Ò#E �C�R�G��Ip�h�y"��L5��[�p}d�Z0���y�(ΕL'b@Id��n'�X����yB���m=�z�A�S.*�)r.��yd��qD6)ikB*P�<H!�N�y�4�1aW�@�@�8h�A���y��Au6�T��F=�z<�1��4�y�H�zA��4KSidTq*�&�y����@T�_���5q�I�>�y
� ��a��ťJ��a����	�7"Ohh��8I]�;@oݚc ��x"O�� ��_�0 tPk�� ,�h�"O�؉���)<��Ԡ��{lРI�"O��;"��	�D�P��#cf���C"O������L㢬�I!b|esb"O��D��%cO���*ڽ&a� "Ol���*0^��ړ��u�I "O���W�@96t�l�ƀ[yz4�f"O2h{Peօi�&����]�\Z.,�B"ONHJCɡ:j�X�$�bN�IÇ"O��`O�F#���C	<e(RP"O�<A�5,?�D8tQ�T�:�
E"O��PU�Y�-�f��B�n��-"t"O���oX�a&�(�b��"�d�I�"O� ����>1߸�K��K8s�� HU"O�16BK�5통���ZO�!�"O�j�.�/������[�p�p�"O�(3�Ҥc�11� &a�a��"O�1��*��#�<���)qNԨ��"O��v���I�.)r���"O�%صɓ1c�sᄃDC~���"Ol�IS`�x-`9�j�;@��K�"O0��ć�Fe�lBŦv9���"O.�"����`��t%��8�""Od�Y��(#��%�ծ�JL�F"O��`	GD��e�E�6��"O~4J�mJ��,�YDKB-۪�hA"O�Ӱ�K���Hz)VT��k�"O�АC5t���CrHH��fc"O.	�p�ڽz�\��	�[0��ȓ�j�s":'�9:���x���6���
V,��{�dPE푡h�A��Rz��r	--p�u)����	Db��ȓr^�E8a��Aq%�&*�ņ�k�����/75J� ���ȓ{�e�D��h(�+è�5=����U�lu �3\�� )'�	�EI��� X���4�G�YF��ӿ@a����q� ����bX��+���|��|�ȓg����"ԭz�!�B�#\�Նȓ0LʵiS"��H��%��m^.`�ȓV ���b=Vjz�3.��5�d��Pǘ�jF(Q;.f ![�-��ȓ*��B!�;��1넑��i��`���gl." ic	Ή���ȓl#.�pb�_?|�\���"V��ȓ6�>"�Ŋ�\n��W�Z [��9��+�A�K:f�$!j��r��a��(��ID��2Ab��.ӌv����f�~���@��AB�8l�e+*D��5��� ����7>��2j&D��ѣ U3KkHAz�kZ+� ���/D���vn˝,H9"����h�G�,�Ϩ��8��I5P3"��RM�|��'�<�+@�<���:"��+�'�����N:�l�5��7�Ki�<�t��% Z��@�\J�IqSe�<!WI\\�X���eI�9���Ѕ�`�<��0C�q�6ںp��} ��]g�<Y�j&�M(ւ� Ma�%�ci�k�<�UA\��%��S�?�a��	B�<A�m��_:�Ds%bD�g|����+z�<9Q*T�i�� 8��
��~��"��k�<� D���*��J%��)��8�*�"O.A0nU)��=�I^�HfՓ�"O��	q�q��q��?h��p��'��x�[)*�j��ÌP;!��HB	�''��K�O��x6��@�-a�e��'��ƧF=���A׏pr�m�'"N0R�U<6��haj�bdx:�'E�"e�I�D$�p��O�����'��%�}6�Q�@�<H�P��'�iI�-TJ��Y�)`�9��'r���$�/X�*� �BW'O0"L!�'��l�Ui~�^4���>��e!�'BV�3a��7aRl����)���
�'"����[!62$2@I�5-���'I�H�)��}Q6!;���95.�K�'<6T(�@��a�$�eJ�%��]�<!EB5��äm��g�` ��mX�<��d#r��uc���h�0��'�S�<���İ&K����c��N>��E�X�<	��T3�]NK� e�Ls� �R�<�KI�9a� �*i���
Tg�J�<��`��(��g#AG�\�g+�D�<�UÌ��8��S�]*/�N(�`��T�<��Vݲ(��ގ9���҇V�<Q�*��	��=���݇k��}�2�I�<)�)\�f��\��C�.���FC_�<a7��4�����L p��c�X�<��o��1ɀEX�aN�'��PC�]Q�<Q��T�i��-3�H&'�E�<)8ZH�p�*D$��%H�<�FbB�A֍1AJ��~�����H�<a��j���
Q�ש ���CH�<A�A$eP.�С�0,2�4���C�<q���X���IH?NڽR���G�<�T�%_rX���¾3�,�Kv�@�<�����HQ�8��%��D�sCv�<�7���/ ���Cg��]��G�v�<�D���J7>uY��4ѐ9�B@r�<A�L�@��l�G�*)�B��h�j�<)�a��M4��b�'vþd�ՇSi�<��)-K��F��"0��)�l|�<�2�p�Мi��YN��G���<YUER6ՠ�$×:��{���|�<��K�ya�=�դI5T�!�eD�v�<���9
�a�0I�+&��5;W��v�<����&(K�L�&>B�Y�Şf�<�ǤSb�j\+��׶�i�Ǧ�G�<�ՠ�!$�.�B�aų e( 	�B�|�<�qR+��mg �5y6�cD
}�<�!�%=���B�	.����
�T�<�d(��:�����9PԱ8�ĆR�<Yb��<%r������
Cl`h�!�C�<95��'(�f�� �МG��Q�g�<�!�Y�QM(�17����,��KSY�<aG(�?͠��e�!^t({��~�<���NSz���kLV�7��r�<�����.9��$&�b�R7��l�<�O������!)�!x�/@h�<iTBK�'*�(����:.�J���I�Y�<���$�0Q�6"�b5� %]`�<�e�ݣ@�>��p�4�N�dD9T��	�G�9�D$b��1�uG2D����C޺2 ^U�aϜ-�hx���.D�8�b�19�й G	�/v�L��8D�� ��%.Kz�$9�e��y6�B"O�<aC���qh����D��7��hp"Oڌ��DI�M釄G�V�=�"O.e !�Ԣ!��DE� =k>UP�"OM��j^-J�j&E��kJԓq"O��r!�J�wdt�f�-		�8[W"O����̓%D�:�	��h��zd"Op,���7�P��*I�T$tT{'"O���UŇ<u��ɩ%�P90�ؠF"O����ƛ4S*��S�ٵw��u��"OL�h��ЊK����.^7K�����"O�cc�c�ȉ���:�xТf"O���g�,6'*	j�C�xrĈ�`"OP��P)�:�a�c!$_��j�"O^�m��-P��32�7S�ըe"Ov5�flXob����ߺE;���"O̽��F�o(Isş
)��!U"O�$�FH\X�����m��
��	&"O��S�.�)!jp�bE- B��e�!"Or%`.I���4KqWQ��Y�g"O���a�;9f��:����`�P�"O4dP­�'��,0A��A�@tc"O6�$iG<���a�*
!w�dx�p"O�h[�KQ'#�Ĭ������p
"O�X���Y5~=�ڒM��BN(�"O6��'B��\��C��#C�yh`"Oj�A�͔��(�k� ܭ���yf"O~���	;Z��BǦ�?���"O�m� �Ϊzc�y)�d��8�9�"O�ui6cԊsL<��)֧N�6i��"O��d�T4R������=@`#A"O���2 Ηe���K�j�@q�"OԉY%�դ@���d"ŧv��C�"O��Cʡ �8�� �(L�4���"O� v��:f�x%�`��!-����"O�P3�OK�[Y�ab1 �[�x%h�"O�a���Q2 � �jP획7��m�"O�ȴ��N��(�J'H%�q��"O<]��@eR�(A�H�!%HiR"O���2(��Q�7K@�"O�a�Δt�0�+�*P�Mh��j�"O�$�2KV6\rE�E!F_�x��"O !���*n�"�q2�:rQ��R�"O@e#���W�H�dhƽp)�p"O�Ir�K5=��X���7M�(
�"Oh�ꐌE�����ܩO�|�3�"O�p �Ή ���$��'�
��"O�z@K�L���թRϖ��A"O4��"�Q�GӲ!�&K�i��9�"OfqK���NG�T:ӈ�r^��
"O,5i�*�=_��a���XVa�e"O<9���H��-�&�#li
�"O��1%�&��%�Ћ;�!R�"O�{�����q�b!��]�&D�"OP�q4c�U�{���F�Z1k�"O�hkS�Ť-�p�k_j�
�)�"O�� �8Og4SA*ώ5��q3�"O�!3@�`&DA���фE�<�S0"O��"G�Ɗos�j�$Qx%�0"O4��r��(�,�s����#����"O��R��!ʨ����  �4�PB"OJ�"ˈ+~�b7�&mâq�!"O��N�v��ș��>T����A"O�ː��M�$�RK_�U`"O� ��I�� "�H���	F�4��P"O���g��Y���'��?8����"O
u0d��1ɲ�p�
�|�R� �"O�u���Gi�٢��2l� B�"O��`!��pnjMP���mH<w"O�A�6 
  ��y�j�.J$�qr@�E<]پI8a+��y��) a�I�ߘSutHRG��y�&[(9�ٰؔ%Y�;�T�B6@��yR?L2�k���Q5LX�D�ȓ[O*Ђ/�)�@�Ue��f�(�'e��1E^<WE*�膻����x�<&T{�F�kk�)�I���_�<��DA�/5B�)���tOT���A�<�Q$TZyb�'�Z9�X�S�Wt�<	��B�����4��ѻ�u�<q�NK�{�:v�iM��ԇ�l�<��e_��>9SH�X��3NHr�<���U��v��sgW��m{3��n�<�D�:q�`��/�'isFTVC�<Y@��V9�y�R$�gw$��R{�<�Q�c	)��J>���W`�<�S��!�`;�o�L�8pJ�S�<���j�@K�-� [&�|���R�<ଏ$iNRT[�&��kb�#�^Q�<��-�'1� xIc�ķmn2��1��L�<y�i�	C}
��Bm��-���!w��|�<I����6R�xr�ր.݀���M�<y���L�zP�N��OֲD� ��K�<�3쎋tZ���W��~���%�`�<�&� P�٨���9]�5�G�A�<i�d�SZlL�����~m��X��R�<q��X2p[fq�D��_٫F%UP�<��'�/p�l�CăNٚ��'��O�<1���� {��4@D�)SO�U�<��I-��s�3&��*҉v�<�&���H����2>c��S��St�<�u ۚJ�j�C�+��C���r�<q��^f9*!�-������d�<Y�̐&w�Z@
SMI���|�fI^�<�V�3�i"JE�L��a�s�<q��U2�0�1�����T��d�<���Hz�Ę1�̞%Q��B��_�<Yt�&A�&�)��L�pP�7jJ[�<�� �	� R��X
$5xG�\�<I�))ޔ��.����`%UY�<a���jA���町S� ��a�M�<A�P�1�q��+"Q�ր+TÖJ�<�)\^�4	@�F��I�(�K��I�<� \�9�-D1^�X}��(�:V� ๰"O|,�V��F�z�أ��:'��)�G"O2�[��#�q�]�a�61�"O�aug\*���R����)�v"Ov�{���)����u��A��`��"Ouqn��t ��żS�D@!�"O��:�c���`GM�G!�p"OZ6iP��q���  Hڱ"O&쩦e�:��H�M�q�"O^Pxg��m�Ա�)ކI��т"O�p��\�i[��K"�F�(1у"O�H�t�Z�o&����F�B�~��"O�\�1�
�|��x"��!�X��"O��#Q'�<^_�M��'�,�ԍ�U"O� ��m�|��+V�%j���B"O�H ���=\�d����\f�L�q"O�R3o��M�<��Bë" V�D"O,h9r$�&brk���<	�Tx�"O�����a�@�s�Q0 �<A�"O���V�ks�Q�ƥ�.f�B4��"O��Z��&(,�y��@3S�2�"O�q�P��mKaeR#n�� �"O���T3d��DʳB�<8re"OV��#��8����ä�-$�H�Br"O	��$��@Τɂ�ٞ2���"O�������$�L�s���:6��t!�"O�0�#!4�)����G��)�2"O�]����'�h�RAT;U�d�r�"Ob-�d���\�x
$�>/���"O^���*��쌰;F��S�"O~@�PI�%�μ*��ЈJ9��#5"Ob��v��r���QE�Ƽk5"O���0��}�m�P$y�B��d"OR��G+"��c��2|����"O8U�5�Ҽo>�z�BZ>yWP!��"O��(�
C��pM�/���z�"O��!���c�²ىF"Ot��V��=xU��
S�d\ H�"O��j�$1DŞ�B$X�CB�AH""O\e��o�%����UwI@H�U"Oh䢦x�!"�(A:�|�"OZ�zu; �`�q"H�"%���P"OD[ �6Kn��4���bZ����"Oµ�wc�d��(���Q�.]��4"O&��Є�|�Xi��'Ӧ>�x�e"O�qC���q�FϠaG d��"O�y�u�3��q����=r�aa"Ot�⡢
r�ir�s��+A"O~����$7��X����i
�D�g"O4ՠT�x��P�s�'�"���"O"<ZO0@�z�JӠ� o����"O��S�EG�N$bP�@�G逕�"Op�Bэ�9@����u^���R"O����K+R��2a��y�ؼ�4"O�$�T-TB��U�R`L��Yap"Ox�HuǞu������L�,�=Q&"O��pg��3eJ�����$7D|Yb�"Oh�����jh�����,��"O�B�ʓH�~��P��8U<:l��"O�)��ĝN�D(S�]���"O��)�A�=uۖ�`a�
�>��ajT"O�{%K@4)؁%H��u�f"=D����D�v�9�(�Tm�T#��:D��i�_m��E����8D�� (��A�� "��D谁�,R�D+@"O�0�' 9�����5~6��#"O2�l_K������Iy6����"O���p����J䘁``k=�Lk�"OFY)���jX�DaՓ.��*""O�-+�,b	�]��������b"O |�f�]"nI&A�V N�|���"O,1k��,�-��̟c�(X��"O��&F�uH�-��)L��r�"O��ȱ�%y��X��R�_�`qKv"O���B#߆A������'����"O��1�#�2�:4�˺O�>`��"O����7q؊x`�AX�zP#5"O.`"0/Ĕ~��laE��6�Ż�"O�TA�)�Gt��2��#�T8�3"O���ĮM�;�$���z<��"O�1�g@�B$�(�͇;״d�"O6�H �T����{�f��b�P�
�"O�jU���;��X�e@O��1yr"O"a	4k^#������6�F]J"OtŃb�[�!pz�`�H�V��X s"O��ɴ�
�O蕀�AZ�D�n�"�"O�ha`B�D�I�ۆ;�X��3"O4�d٦H��Y�#i��o�����"O�YZ��sV���Ț��1�e"O���%�;��0��/��GEh��T"O�� c�q���;��ҵ@�)I�"Oxp $[..�:m9S���dV��qQ"O�J'G
h\I�N�9�n<��"Ob��b&�Bk:��`M��-�V�1d"OZu���0J� ��K�!@��H{%"O�y�ǁg�F ��jG4Z4G"OV����]���pJ �J:&�
�"O8 :�D[n�	�b��kĈ�"O�t��\�4f��Pu�@)d�y�d"O��z&�߮}� =��`E�eײp�"Or��/a�d
��B���U�5"OH�u��5�"Px&a��S�����"O^(��"�0\3�/e����"O�aB`��`R2@�gOP�6����"O��֎QHd��	���#"O�p���&�����1�2�@"O�![��JsV8;r�$[t��"O�l�E�Y��\�z��K�S�"O��a�;%_�0S��\ ����'��m�V���S��4k�<`F�x�'�"���͊
?Y��N#@��'ܡ��Ņ�[�e��IL� U��i�',֠������Ɛ	�+9��z�'�P`�i�|B�A�ა#訌C�'ՠ4Y =d�`���&Y.{�9��'HhxXЯ� �b��2�\a1�e�ȓ7q�Ѡ���3D,DP�e��9OX�ȓc,(��Q�X�?������3tdq�ȓ��1qQ���2��h�0K�nh�ȓ�"�x@�/�ؤZSf�� �͇�,Vҁ����{�P�s2Kpǲ��i ��{�ćc�H!��P�im@��ȓY�����J;!;Μ�''V��9_�ȳ@E��|�>D����-A�%��G��b��PA>���N->�H�ȓt�Jx!��fn�x`�D�.g@	�ȓb��w�H���Rf^ 6tP��ht�@
d,��*I���)L��S�? Z�:W�_N���2�[��Xf"O� h�ě;z�lU�D��� ��h�t"ON��p 	���8э �nw�l�"OdB�ή	�4�Q��[���c�"Ox�冔4]��{CBאdq�1��"Orz��+˂0��n�#yf:9(B"O��L���L�B�ɒB��(C�"O��sA>ZhP00.Y�q^H�"O �ů��v.���]�j�j7"O���$��<�e�B?V-(AS"O�AiQcKY`D�DK�. �R"O��,�>Gx\�	Ն-"Xq7"O(��@�ZkL�ℊ�;# y�`"O˕�g�2�A1gO!�"١"OZܣ!@�Q,h��uƑ��@C�"O$(���� �Ԙ�3E�R�dA!D"O�s̈́�{H64񡣏�jL�3"O��8�N�wt�qw�7#	0�c"O�Jя��!N�V���J�"O6D��	� ��%L�c���Q�"O��F�<4�t0�Ķ2���u"O@|[�E�~~�Ub�����v"ODPh������D�F�	}"l�u"O,��gC��YȞ���8w| [�"O��u��vD(����Mh2��"Oд���D0�$�r C��e���"O��a��/1d:�ȥU>,�4"O���؈j���q�F ~�`|�S"Od���+JB��u*�y�k�"O��񅋑�hYSO��oa!r�"O��A
:�4��cQZFҡ@�"ORap�'L���K���&��{�"O�EKC���<�C ��j�Z9IU"O@��/�/���A7N4D�,Z�"O,D��G�-��ϖI����f"O�� q�,o��Ph�'�6q"OJcsm͌�$+�q�p���"O�M��(�7sP<�s��8��f"O����"Y�8,Pb���I36�#"O�	+�$���j���]�$8�"O`y3��
���L�3C��Y��B�"O*h�@fF�4�� ���VX��"O��j �L�]�H2-�!V ɫ"O�ph$`ȎV��]�NH�H�dap"O��Q�0�la�Ȏvy��ґ"OB�{�Ö%h6it��'2pll�T"O�����K�2(a�&gQ�����"O�a���F<0��%x��$y�,��"O��a`hZ#�����|r�P��"Otu�eZ�E�`�2�"�i]�� e"Oi�&蘻.2�H����QW2�P"Ol�@�f�"�R��֏�z�zS"Ox ��R�,H�h���(j�\l��"Or�㰭@'pXL5�H2��	"O�i�]���a�B\���"O�;.��)�dt���5e*��w"OHܫ���]��
gm�#D�t��3"O����;~�%sĬ��E�x�B"Om�!HM��Jq��bP�S����"OĴ����.��/��� g�:%!��F*Hn�P�#�Z"�P����7!��ą]<�A��9�ĒW�CX�!���vTXq�X;��0!�"7V�!��G�B�^�&mסO���u�$ �!�� �A�d��/1�mc�ǺS��U"O�P��%B�����M�X��yG"Ol�8�g�0���4.�(v��͚T"OXkE_��L#u��<��c"O�aR����T��2+"b� �"Oj�2��X�+9�p����1
ܙ�"O�P��$�O7f�C0�r �r'�S�<���J;
E��F0ỳ�[� �Q�<���6��@��Z#+�b����O�<$�\��HeL�X����R�<��'A/r�.�z���i�Z���,�V�<�J4.֔0�@�Egٕ�S�<Ie��1~u�g-Y�5���*ǄT�<a�n���t��V�^C��IG�g�<9�M��6�&��b!��+7���c�f�<��E�\����	��`��,�^�<� �5���!�l��q�C�Td�<�"��l�r� �-����Nd�<�IπL��d�2��t����L�^�<�s)O�#n�����:mw�]��m�R�<����o�tE'��3] Q��K�<��J�-9r�B�_2ZUJ�ʦĕE�<�f哛~�@Ⴕ���ܛ��QA�<iwK�gkl���ԛK��!)U�S�<ٰ�L�L�>��d�@3iD��AT�<y�
¹}|�v`F%}8]��AS�<y�K%�~���#�|�3� S�<	W��##R�i %v>�\�4�i�<u'Y�P��(rU��5����c�}�<�CmP<9)0�5G��j)W�`�<᥋��K>d|�#�F�6�KUC�b�<��N��sX􉥫F�/�0�z�_�<��B�x�P��T�9����r�Y�<�f��8=�b���\)n�~i�P@�J�<q����	� /�98��TJb��N�<1�d%^�>!���X�<s�%�P�<q�Ƀ�j��DF�&�h-�! S�<�e%�f| ȕ/J"Q̒��U��Z�<'lX�>��<�0��^�x$NOY�<	�#��`�`#)�jK��M@U�<�'F���
9q!�UZ�<	u��<P<��G�
^' 4��iIT�<�)��l7̡���bƔ.D��"��uP��	|��u�Q���t��l��U 찂ӵJ8|����� ��Ò�{���p� ���E�~�����l���HE�1A� ٓ�R�Ė��ȓ?�8��i�0&=.�x5L>pȄ��)����*�O\�8�%bQ�^����{j�`M����!�Z�<@�ȓL�}Rv���-ٔ��T%�̇ȓbt�E,,uP<y�����}=DS�Ђ1/Z��7��C�}�':qO��~:G샙|���Fn�&Y fm�S��!��c�r�8��W�E��17�YOPɆȓtE��a�{��A��Fي���X?���ҨDH����&@���w#�;	�'�ўb>��D�`&d� -�"��$O�O ˓_d�Db��U̶X
�iۤYS\��ȓ)���ȕ��Gm��h��'$u�]��IΦ�q��FovĠ�9ʬ�J�@�7�pY�=�������aP�����P�	]
�w�ʡf+1O`�=�|��T&.q�EZӀ�(F�}a�G�E?y�N9�O܄q��8���H� m Z����'�a{>� �4r��ɶo�nS �"e%h��"O���6��&a��{�,Ɩ#�LUZ���D>�t�H�ZZT#V
�1��e�>��y��`��!�2��]�3��ZA�a�e*D�ܲ�a�%�r��!�	21��*`j4D��X	�(1�5��}ШQ��<1�*JUHD.� jQ:T�ro�^^P�	�'��O��?)���:7Q~��4�T-b��
a�'="���d�J��*�����M�l����O(�=E�deFs��s��V�')���pI�O>�=%>�а�tԦ��(ݒaVA�%D����E'S�pe(Z�!&({��8D�H�jR�hڒ] ANZ�e�4H�"8D�< %�]�A�`��E�2[������+D���I�:)����� gp��P�<D��cק��2VJ<��]�xa��x1�o�Ԇ�I�
cU��\b�pZ���l��B��5Y����Gʅ�\�Q/Z���C�I*��1"
���p����K��C�Ƀjwjq��B�8�Q�_�ւC�;Q�v� LH�?~@
���9�r�Ov��[�T4����Y��$�@�Y$���ȓurb	B�+F�0�С��@˨.��1�ȓh��|���G���뤁B+ �%G~��	�?��+ĶXcl�Y�LcWn6D�„�4hEc���y:N��U`1D��kd훴e�t�#햣,��x�U�-�OV�g��pI�!�>N�6 ���X�@`%�@E{"�{�"l��/`3�0xg�YJ!�ȓ[h�B�@�N��r�"K�O!�� �	Et	��\B��9P� �j:!��� cL�!!��Xɺ�4�0!��A�(�v��$�/l���g�� �{��T@��c��w&��c�"�,�a}җ>ŀ'4�H��Ir����'Ku��&�@��,��afB���!6�X�:'�+D������8\�H����\�O��`c(D�$Jf�;3��u�q M)��`e%D����� J@a� �4
X��e%"D�x��M�B	@q biɥ8)|y2>�I�b�Q����@Ԏǩt���^��i�**3�!�d��K#z�����H*���2���C�Q�8��	&�4���G�(P� a��zC�I!��|z�� �-�2����_)D �
O��;dևT��1� C6!�舁��'�O��97��&�`��'�O�c�R��%"O$�+��!f�$�����Z���D���'���d��U�2�"�j Np�]R#"OrE���،4�b���N/;��ab �O��=E�� �7r��c�1=��� �C�9�y�H&���r�̗�5�l��J�yL�� �A@%U
Z,& C
�y�+����I����K����z.�ņ� ��@��<:e�B%Nn�ȓI���k�D�=R�1�Q�V�|��8�ȓ/�%�3�P +��XA�G>11%���I]���yD�ͼ��4�pm� ��a�r�%D�H���9�D��׉�g���ks�&�	\�����D�y��Z��Eqʤ�#$f'����p���Ƌ�|�r�'��RD0t�Oj��D� J�iP�L!�=j�
B#�'q�|���H0�P��4(�x9����>!�O����J�Aj��C�Q�*�	�"O�x�C]�<"�MI=�"�ñ"O� �`�P��9Z	m��
ʠ��YJ%"O�H��N� MҐJS�0�2��'<��\�]d�;� �I�҈��l�2�=E�ܴo��|�D��	J��&�_=&#�y%��E{��d�Xu�j=��cH9U��:����yÛ0��1 �Ot�-" CP���'�ı��	6d����s��n*��#��%!,C�66+dd4�KdxM��L��HF�"<��7{�h��] VD�w���W�>Ʌ�	�O]��/b��"�	��gd�UB0�UhUBO��u�R }�4h�A�+YsA ��'ޑ�s�a�M�����ۣJW���p,%�O�I�A�@�#�Ѣ:t�a@u����cy��Oz➠&�xYЍX�\��)U��~/��0�$D�����(&�L�1ۻj�r�A!�t��'�ɧ��U�F+��Qq���bt�C��,�!��#'�X3�HW�fp����'/s��=E��'odm8�@B�u2�Y��)��<(���	�'�\�mD���ʍ=/"2�
�'��rV�ǟ���B�-.p�	�'�*� B�"&�������ss���'hT�5�ȜOt����O�W4�]��'^��s�hQ�U���	�?z�eA�'��]原(+Υ�PD��0��H�'�b �o��O���3��I����'�:��dC�/�B�z��Gِ�Q��?!/O�a��#	!�҉���={#<@U�� LO�����=>�@r��?I �|�&"O4��mJ�o� �zB���5�LÀ"O���RcD9nzQ�׮�8"�ȼ� _��E{J~:�O���a�b)�bf�T�ڰ(��"O��!��}����×�8�������<���)�0W^J���D��a��ab�Y�0����7b:a{2������&<ޙ��m�'!�=*"2�I
!z������V�S����t�G�a�%+��<c�*C�	dњ��A�D4R-v��4eɳ�1D��u�޿S�E�K�"�;D�`�Q��h=�v��~�A�c)<D��4%
)�,uc&��9\J�@��9<Ox#<y�,K�Y��E[��_�B�DqT�Lo8��$����%�B�)��$�z�l���6,O�'���S�f�J�U��X)��@�ls��D#?����Z��`ɓ��<0�~0�r+�<��x��'�����`�>cY�sS�ݼ�y�O0~�!��Ō;_8�bSK���y2bž=v"�G�Yr���R
"�p=A�}"�'"�DDA�+�	�i��	���x"`A�\u8���ZjM��"|�!�d�%ZHڼ�UPo��+s���d�!�$�N�2��EÛ�L�F1y��ߧR�!��+b�U�A�7HF�x�U�յ1��y"�I|h���-� xd� CjB�B�	�Q���ťt8�;���
"d��	��HO�>qB@�_�n-��b�
�DI��%D����̻MF�'
'S3@��7�8D�D)C�X�h�$H�`"B@?U�!�$ǯr�ij^�E)��ǃ/�x5��'�x2V�^*4qk�58��Q�'����ߧA��H�0a�6ޮ�;�'�4(+�BG�,�9s��W�3�`-!�'�
xh�n��L��J+�
�H��'yԺfA�v�4I5 �;0nY[�'5*M��H��iZ�2d�I�1k�'�N��'�*Ij~L��I��$ђ�`��� ����)=�X���'B�0�3"O��3��$;�l"��L�Ju���'"OF�0(�*W���؂�_u�`�K�"O��R�.�������%�)]�f5�r"O���7��,�N���:CL��@"O��(vH?� !����3%O�j'"O�]BW�-l͢=1��]`M$��`"O���E$Y|R!TE�+B.����"O|��6.¢3z\a8����J��Q(�"O䴑T��'n	|�4e�tf\J�"O@�B
^ �b5���!;�d4��"O��qE
;f�`�1F+�N@8�*2"OH�kA*I����m�XC�i��"O|!q�i`�*��T-�GTXH�"O���*E9d9< {�R�0^Ƞ�"OPω�At*���f�(Z��p5"ONL�cG���R��^�*�U��"O���%EW-}�ب)�a�u;D"OP��S��&BDl�[t���M�1"O�i�I��|D<�$�S�7��Г"O�� "K�G�)��L��@�(�@"OF�A�#�>rs���L�$̶���"O�|���]_�x�
���X`@"OV2A�B&����i�,e�w"Oڹ�'�T���E�b�l����3��'�r �Dj��B��@���;�B�S�yRID�g.8d�I���*|�4����y"'�F���C��Zꛮ�y��LKr�-����l,�ʴ��'W`�JEGB��P�(�"ȭ�AH�'���b� 7~l�J0�V�1���
�'<�\�0$�2�l�")��~��]��'<�DS�ف�
ٲVI�����
�'}�	�"ʙ�0 I�oJ�W�T�
�'#�u�5f�ZSf�q#�Ӳ ��'��h+��K*.�q��P3u*h���'��j���F�"q0P�T�B��݅�=�j���P�:��܃�AC71Nv��4FL��P�r���/��`���ȓLp��S�S5i�شk��K�Y�����x�^�K*�-BF��I$�����4��E*�< ]� /@<!A� ��͊Mڔ
�ڠ	eh�UH�|�ȓ9k���}u8�5�.$�rd�ȓCl\��퐥L���hUV�Q�v�ȓ=����!�R�%���+Y����^�©*5Z[��1(A�˧*Q��k�d�q�T�V|� b�k�$�nڌ0�����bQ�nFh�����Fkî_HN��H�5]'$��#�:�y�H˕&�ҙ`����R"ʼ� �H��		WJ�0��<6i���I�mE����_3D��TA�&����d�*M�`ұ
O�oA��E�ֳ@��ʚ6UʈPfl��Q�n5��0K���]��@+��_��>���T�K���Nr~�2�д��� :�%x�ݑ{b���g�)ImB�I�zEJ�Q5��'"�HX��a�f8�I�ĝW�dR.Ĥ>y��>ʧf:��E�01U0!�6x0��W���B��<y޺<�.�%L 8�F���P�؛獋-��h��@�o�f�!���<xܼ,E{bI�v=r�ؒ��LͦE�5j�;��<Ѳ�ھNɬ]�E�M�'���Q'c�X��h�F��_.�Lsu���5�����O�h������|�#@�P,$R *�B�:�'V
�ⓓ9���V:��r���p)0%�O	f8єl�0]0�
�K���|}��'���A�C!wXR�g��>�^݉H��,0:� ��qp�p�#-՝{��	$?m�C���yw��,~KP}S �_�m_�-)�
W�Px�*��!t&�h��?3qV�!�O7x��2Rg
T-��{�'�,��\˷��/ p,�X��*ʓdU��� �J�>�@$ꧪ֤%Ď���I8*���*�H_�^��8c�J�� �� X4��c��}e��%GMD�|H���>�q���p>ic�S�gEn���.�/kv�c0�V~2Iݾ=[���`�)(g�A�1,�.5�������/q ���x+�Uq5 	i�2�v�[:��|��'V6�����X�j ���N�)w��2�E�	a��E+mb�D�B�I)%U2�O����fE�yW�7Yz��SU(�)j*����S;�xB�A7[FZ��t��>,��FeZ�d4��D��:I�ȓ�gZ�q(6 B
ICV����	|�'3ֽ�MQt�|@9U��\LĄ��o�*�����+����$�D��C�܎8�����N$�2�F8>�Ͱc	�.�����SR��7e��{/�M�PAY�;U�I�H�T��t�ðO|�,3���0�� ���D;J 8�Tן�����F�:�}���Ӌ���'"O�%Spb�5f�*�Hu��*�|��6�ݰ +<d��R�8U���n^�)CH?]�%.q۶��?p�F�Ӥ��=��)�cZ�y�nB�I�q�L`����S\��A�փOښ)	��G6|�MrUE9{t	�d��EDnx�w�ݥVWQ��7�T�p�[��U1~I�$#$O�� ���_����1�%/����=w�i5��*R=��C�ɇ����3���T>�*�kt8p2�+��F�Bh�$,�5 J�i�'�ʕ�0��oI����-O�H*f��C�]���Q�6�y�q)�n�|d�@B҃0��	U��v�<a$�C�k�~5A;x��-��¯BX,��lF�WP��w\�9[&�r�#�$�ٹGu�\��wY��+�"��f��2����'X��S�X $�岳�Y�h*�8�"fL�֌	@�"�,>`����)j�8iM��,�#=�h����p��%2K�Q�儌B�X��÷,ǞQ2��."n �Q$AxL=�8Je�ؠ��ɨ%>����!ڴ��� h�0
��I<(�P���G{���'�pH��:��\;7 A/�R�SCI@�"����X>XB�Ւw�j����?HD���6D�t�R��a{�I�j[*`��Hq�҆.�h@Z6�X�@���2�k@� �>��@EY����pd ҭút�,�;S�U=���$�\��;B �DyL��!!>��e�FZ�!�mq�'�m���^n����d�.=��k�/�
�5`CfMfay�"�8:�!B�FL?;���0�@�b%�2�h���� 1�̕ ��ԩW�~"Hܲ`w��IY�J 1R`���N���F��5;gF%��Hp�$�_,8�	R$�_�N�8Ux�*�g{!�D/�N�Z��.�ih���/Fh"�r1LD)WtƁ���]�'��r��Uy�Z��|z�"�/���������y�L�xG�U���,H�Z!�3��8�Wd�5H.PТ�h�!p�9	Ó,=(�(�b�Q��`q���\��4��	�.J��+�K10D�Fl��ǖ�Ad��CR~)i1K$�Px�����M���ѵ�A�2�G��O�� R�Q�> $%�tc;��}�"���m��YC�Ț<��C䉄a�I$	D(�ƭybLç-��EX��E�v���g{�@C�Fڔ%�����*��$=>��K`/�~`���#��p��˓�8��~҇�	�`���`[-Z9RJ�ϰ<11K�+N�jH� h&#ӊ`���$��d�r��*D�|kC�,����˾aE&(�DV�6;�A�@
,��i�)=��x�\1�����Ʒf��Ȅ�g�2풓J��Z�<u�� S�[�|#vO3���2^�P�~&�� g��^��h.t�Y�ק�O��C�I�<!���W�a@yr6c�[ߪI�"��Zp���	�;<�w.ܛPp��RãK��v��d�92��DK��'}ljY"ARn�3c8�+�ύ��y�M^�$��4;gE�^��P��&�����4Y������S��ڈ�g�ƎUST�"Nd �E��9VcA=5r��
6�T�m�&5�� %��?n�2�~&��q��C!j��Ѐ�� Cw��1�D74�|�sh��_	91D!F-p[Ęs
�>��4�� 1�O�4��)���IJ*Mnɔ�A�'�T�Rs�x�Y�'؝�/�O���"o��y�ǉ>sv���b�(C�zHq�F��yr��A7�e�wC�6G@2=�F����y����1�n���oL����LJn
B�I]	:��GA�T��`a#B�R_B�I�Z�S����бx����M��C�I #Ǯ���C�h�HAA5�!ϴC�ɸP����)��u��h�v��''j~C�)� $MQ�D	m�L��c�*��Ah!"O��[Q@��,�Dj"��YJDТT"Oj9�#�Rt=�`!���<X����>�bD�+z��?�U�
�V}�1�,%�Z�O)D��yO��U-��iu ��K�6��g��F��Q�$y��OO�g�_z�YF(�B�3P�+�� ��I^v��a��zr���煸`�-`ϗ�\ꍀggX��xғǛ4$B�5c,@�<pP�9�n�P�X� �v��DP>m��i��U;B��@��
�RQM"D� �������se!��q��LP�n�<�/�r
�r�A����?}�B��tA�-pP�؛���r.1D���! Xo2$(�2����${������'n&�ص�ؐ3��ϸ'�b�a�H�?�<|��%�qK��e�l�p����� g��a,�@�ÐY-\��螁r�}��]s���Q�Lȸ\<h�a�(��O�ɪ0'�j���@F�ԎՃia*|�'H�� ��0�nL��yr��$2h�1p)�7�m��Q���@%V�t�t�@'��F��IΓi����#��
��|��8�y��:Ӽћ�G��y>�9d�wF�$�#]��P��k7�c>c���L\'z<���X�`"yA�l!����>5H�T�׭� Z�NqR�ƿ'�#$˔߸��䑅)�L�'�d���8�C��ax� �,;.�<����Q�ĝ$��Q�H� �J���2Z!�$�#)~��"@�(��,�#�Q7�R��q2ǚ#��S�'rIc���J�(4�f�6LM�͇�EP��…	" �*�­��[�{�֌O��c?Ox�B����5�R��&��9�Q�B"O�,a� [� Z�hH�%V7�@�X�"O�y�B۰QЁ��	�ؼ��"Ob����L���{2��53�H��"OV]��#��Zφ�Z���%'4RW"O:��t���_dT��I�!t>�$I�"Oz�	D	�
�p�h�2"�őT"OJ=�F���r抙bM0�@�"O:f�T?v%f���Ԍq?���"O�ԺS��,G2�a�;m��Hi�"O$9�¹#b���[3O�|�Y"O��vIF*<�`��6��}�C""O��B�gV�k֑��Ѥ6V�2E"O���c&�$4�8��ӡ	88	f"O�DsV�6x�"�;��	'� �"O�M{Rj^^�$AQNOp�j���"OR��Hܡ1�ƈF��9�0�@"O> ��ӤeƝX�VӶ�)p"O@,�Eg��T�di���5�%�3"O"\CR���a��=t������"O6Ta���+|L���GB,$��q"Oȩ ah�]r��F�k
n�T"ON�yG茰1���xqf1	�ڡB"O���P��?>^����c�.��"O�e�d�Y�bM�A35I�<&~�Q"O��$���$� qx���J|`3�"O��3p@L�h�ht��읂
�"S"OX�A́����Ӧ$G��%�E"Oz$� �KǼT�Rb
2F��"O��	C�#nɚ|B�Ո H	��"O�x{ �k����fЩF�ڜ�ȓc��a�26J�DHB�S�|Ղ%�ȓdz��8SM�>�0�H�Zq�����j�{SD�
<�ڵ�D���t�8��/��u	f㊞lp���F�-ror���r-��i���7���A��oyH�ȓ'H����HB?&񋵂C."f�̇ȓ:�P(��RbDb©˥Z괇�S�? \�CO˟n!�)�p��8����"O(��u��2/��zA�<~j��"O��q�ƳSn��9���ZZ=Ka"O�x�W�Z+U������CaԹ��"O>0C�BM;���-��w��l*�"O�P��A�L���"FU �T�A"O�K��#w�`l˄%Xjɦ�2r"O"��P�I�lS.�9�=q�52�"O �����H�
Mڰk�j͊ـ�"O���d�MN*d�I!n����w"O ��Ƌ�(�j|qT��� t�ң"O�i��%A

-�^����7"O�ؐ3I	?ud#�M D:`l"OD���ݶi)�&H�/G��: "Ol�	WC@1G��ԓ�I<�����"O����GE(%$��3�R>Z���B"O|���MO}�d���� ��L�w"O��:p @B�r�KL#xژp�"O�,��C�9ČY	�)�VW�	��"O&�H���^I����"VO���"O�ѩ�(�(A���èG�K֙��"O����_�)�Ĕ�7o�r!�"O�D�&�\�_�B�:�&W'KТQkr"OR����P�r��3*9���"OL�;�˘	!�Ѻխ�	:>tС"O.����,4s�e�@+«Y����"O\�If�"���'j��?�:�B�"Oh���șE�L5Y�M�I�.A+�"O��3G·e�%I�&�vm"O��g�F&L�j��bB�W��+ "O��{�aL�?`�M��̄7_j��D"ON-r�M=+j`8�¬���1C*O��*C랞r�䐥튧r�\��'��	��X�|hM�$�ȠcVZ��'BF��7G2B`����\$C8���'N.D��H����d@�B�1�'+�!��16����Κ�B���{�'h�H2'�	�����'�<���0�'G�����m��!��Q�:�>��
�'I��2U&��58��s
�3̂y	�'L�=@�B\%5���+6�3u�4	�'l�R��'()\���.@e'���	�'W�<k`���3B"\4�Z��'4(�w�t[�xJ��NL
uK�'jÎ��
e��%W�]���
�'���1b�B�ذBF
�H
�'��֮˯y(�3�M/~|.x;	�'����OhKެ���D�p�r�z	�'�pQ+���f"��ȋP���0"O�=�7�ʰ>���G③v�.(�6"O����l��C�����bO�*����"O��XЩĎ|�6�;��= ���j�"OTl����R-�0p�f0��x�"O�$i��2v�d��>^� 8(�"O4�8F��R-�]�ϕ#����"O���d��xjz['��9�|�x�"On ���R�P��g�%��e9@"O�2����S���х�y�"$�3"O���Do(n��c���ET� RP"O�T��'g�dW�B9<<.���"O��ه�TI�R���$�3*,`"O����S2̢���V�
,�0U"O`H�e�+@=6�:�L���*A'!�D�.r�4����U(�J��"l�&!�� ��j���/W����ϐmj��� "OF+���:!��P�ɇFP��C"O]���Gs̴��ȗ9DHQj�"O&P(�ʁ8rY�[��V�3<�}�f"OX��'��:#@�� d��V�{�"OPđ ��"BLڤ���F�j����"OZi	���#8nƸQQ�&H���"OAj3��9�����G��E�!�"O�Y�rD�]�����% �7<4��"O���]+�񀑥��:��r"ObasR"�3r�����ę�ZQp��3"O��0.�3*Ĉ=`FB��RL��j�"O������-�2y�3恁1L�a�"O�ઔþ����C'8yzA"O��
����R"���K㾨#�"O<���K�b�^�!��)<�}�P"O�9{�F�;���b�l��J�x�9"O~�;.¬���nۆ�,�`"O����mC�qAΌ�tnG?(��'"O���T���e�d�7���/�Q�"OrL���ǽgO|�yb#Cc����q"Oݱ�a_H�B����)�"O0�#�EF9A:p��$��{fE��"O��8S�	��z���Ѳ�"O&�� 'j蒝1��H�o���Ё"O0�Pׅ�1�~5��D��"Y�x��"Oظ��+��Ix�A�Vl�y$"O�9��C�x�L�v���@�7�#D�( ��	��[�RH\@��Ү?D��Qǧ�6vҌ�S."�H0&�&D�@��B�u�h$�����q:x�%D��qFD���� � >��4 D�`T䇜I_�,Q�C����#p�4D������G{8��d�ͣf�d���D$D��@�͟e���dG�A#j�k��(D�0k hP+I��<s�i�n�X]��;D�����_����0"g�+c����9D���7jF�;���w ƥ_QY	`F5D���(�m�42D���H	�k2D�TI�N���D��� "�����4D��a��\C¥��Ėww��:3D�0k��Q�:�
�G@&s.��kP�:D���f�ɂe�4�Y���/yǆ�i������'/t�G�,Oᨃ%̴%��M��pn*��O��)Ca�>dݠ�j#Y�}d�t��kP0�k��'�R�µM �@]���ȟ�r��Y�K��0�A�P���	2j���� �א
�e�q.�4��B�	�M0��2���x��%�r�`O>�����<�O����&l)N��:s���e��\5"O���7��>��l0��Y%m��������o�ܘ��x�ϝ?��B�	 T�Q��.�ՐxB��[��&g��^i�T%@
d�!rE��op�~bl+D�P�C6G�O��r`M	��<���9��AH�H�E��U��hw@�D�|�cg1D��+�Ȗ#(^��O�2e|Ր�i"�D�n���Q�3����3}3����ځlܑK�
֜z!��\"K�n��d��GoN���)��9�L>���L���'�(��c�[�<
�8�Á�18`��J�'}�]# �!pm�dI0q��a�Ι��vt�	� ��ɹ��A9�.(9���k�Fa��	0
N��%�����:�,��A�/F;8���K*D�,w���U���k7�����?�y"K�>1��{��W�_>y:��7�y�n� S2�H�`�VCD�BViW��y
� ������M���� ��\ָm�P"O���dƂ�J��T$^�W��e�q"O��x$��U��!�ˑt�����"O^E��ύfMp=��Ǟ'��d�4"OV�AC��++�F���:rHة#"O��J�	��q�ThہD�
�RIh�"O���"��!�n�0d�rY��>ac�]�`�l��?�+k�:������{g,�y�5D�t0u/ڋ-�C��
4�~%�!H�R��j��bF�b�g�
ty2���}d�Mq1J�xA���	xe�B�b96�z@�v%:�sI��+�,�#�o���bgAP	�l��F�P��� �1�@!4L�9BN9��V>�C����0:'"����c�;D�,��銭���ٕ!�`� ��`��<ن�ׄR$�)�4h	�?}#��/oByjF�O�f��i٠k/D�d��픬l&� �0@�x�U�BjL]�D��'`$�gL�To�ϸ'�����0{��0��j#6(�	��q��)c�J75�!�1O[	)P:�r�B�w¸�	�#ߓ��}Ү�+�r�!���/�֐:��H���O8����0� 
3J�r�D��{%`��%��!<\쪦-��y��BN$Q�d���&9;�Q���d�{�f`�$��.C�VqE���� #��Mr� �'	� �RƯ��y��_&^P��a�t��P�Z�2���uR����C�l�b>c��ԅž:�C��2Y0ɐ"4��2��D�p`Ӂ��c<� ��X��<�[�!�4����V�h���ZQ�Ԧt��9a��P�L.ax�M��Y�8��7�IS���y���2J���UH=�!򤛥*��u�%a��P~��IC�I�s��/��PK����S�'5�0zDA�0=F��)�Y����^�%)%�<,��D#N%��H�{g	aN�c?O>���*�!z�59��bO�E��"O���'?�,�K�@�6)�U"O������]ݞ�I�!_��0�"O�e��Yjo�)��'22A��"O��Df�H s  �n���hG"O@J�ğ�C�Xy�M�3\hF��T"O�4�b�6
e&���K��rBF)3V"OF\X�p0�7�ј�|��k'D��R��͇Y�,�c�=u̎��K)D�h��
M�h�JX�˖���� 'D�p�aZF��Xp �?\ jl"�n#D���1�׹4�`d8�
(�V��%�#D��E�A/&%���@�X+^	2��p	!D�P�q�Ȭ&@B�q�T�f�\�yG->D���iS(l��t䀩��k=D�l9t�M`iV�"-�H�0���;D�h8��	
u�T"t���2�;D���G!&����Ճ%��@�9D�\��L=M�D�P�!��T�<�&�%D��	EC�~��(�F�`�)"D�L"`�C(wsf�0���\��c>D�CRX�jWz�s#
:'y��H6�<D���be*%��C'��YG��q?D�P�$��K�mc�J*d���"�0D�����G^� �4n_1!�@��#D����i�zžd��Q=jЦ�A�:D���E$[�R>�R zྌ�U?D��ん�#"u`e\�c�a�A�&D���Pl��L�~�y�� P��Sa)D����A־��ub�;c���U%D�Љ��N�#ɞ�s(I�>�A֌"D��H%�ԦL,�x��+,��(t!D�d�R�Ȗf0U��d�1�&*D�b��Y��p1��T��+��*D�� ��Qǉ�����E� �v"OR��W[@��-Oe�0�W"O&`q䡉��("a�O�F(��"OB�����(��Y���;��'"O�Jg�ò?P�\���U�����"O1 �S�  ����l�~@c"O���hď@��$��`�	JC"O�4"F�\��(�I!ט���"O�ig	�2p�ޡ�2�&N��H�"OPqy"#�d}΄*Ѭڡ1º�ʃ"O~�Àí�8@@��OJ[��3"O&�83F�,��@��'N�� "O��QF�*N����T���j:� i"O���&[mĐu�
A�_��
�"O������m}��!`��+(¡CQ"O�Y�(D�^U@�*���n3���C"O>���?�a1`l���"O�e��hW@@��JB>:*�X��"O�EJ5�K{b�*5υV���y�"OZ ��Ϝu�Hաtg؟W�Z#*Oxd�!X6Y�����*��(�'TL��Q�C&�Ԉ�B�� �0�{�'d	{@��+0M�r������';� B2�ڰ�~�I�$%����'fh�pwOJ)u~��9��ޭ���B�' Nl2�H��  "@�U�*Z4Y�'�q{R䋆Q�.H�'�0�p��'��=Qfc�X�0i�5Ŝ�)BB�)	�'�4�"��aR��D��@8Q	�'���{fD�q�e9%"�����'� qɄs�b��ԎF��)�'Hq�q&��zor�Y� cP�Q�'E.�1",'j�L�)6��u`��
�y���rn��z�$�$�~IҦ.Ee,�'�B{0 �&��(��b�h�O1E{��	�w&�0�"����A�5�%�r�)�'Pqv����\�V�.���n)c�6��0|�cD�-tp�h�*�t����i��hO�4��P�  <e��a��}&�`F{���-�.t��e*Jx�h�7����$W��>?�;�~�O�|�ϲ `r��I �|�"�[VA�;��(�O���鼟�ʒ�ޡ^��q:$C�Y�N��%�7,����![���<ݲҧ�O|�A�1a��-0�y#d�q��5��{"��8�(O�O�ޱra�/6��	#�ܪ=�d��M<Qf:�S�'9���	�mA�o�
2&��'��hDyJ|�(O0��D
�����a����Jոi�JE�'����ȟb��	�>�1C���M�h�ڣ�<a�,�<ѳ�?1��T��	��Eǟ���W@�A�.�£<%>��#��?J�n�Sg���� �."��(O��|qh�)�O����@̀;f�Y0_�|�$�4�S��zy"��KP��_������ �m�*ݩ�D��x%ΗU?��ӡQ#��E���i dg�9l���A�8��'�q����
P�y�C.�(a,=��$
X����;y�>����M��'st�z�|��)�e2�t�E�	ʔ}�5��I����hOQ>���I�e�Q�A�LS�0Ԛ�,�O6�=E�ԏ�<���7��
,�l�p��!�hO���Llǚ��Aj�IR��	!�CбO@6�#��?}8��lư�s�eߠvb��f���l&�q �"Ox�����	�8-I�JQC��ۄ"O�P)��0"� &*ҋ��"Oސ1��ORe:2/A���$��"O�S�Ɛ:l��Ä��h�H�P�"Ob��k�E�M{�H� s���"O&Q�/֫gI%aq_�kCb�qR"O� �u�RK�85�c�9T=T9g"O��p��	�(j-�K�%'<N��"OBe㦫��PJ��1�Y2(7����"OF�QBO^0A�6�QA�T )���"O�9R�޵ A��b��?+(�26"OL�M%��ѡ��׺])�i�"O~}Q@��>���Ge<t��%"O�iK��Ҩ`�L%9BE�3� #&"O�};T��@������x$��"O�4 "�P�F��q�b��))�|H�"O�@iB�Ld���(,��
���a"O~��d��;B ��KD$YU����"O��� *��τ�s��L#D��`9"OHe���3V��k")�=���'"Ov,撔|�l�#0���y4"O��R	+-�tɱ��`�Z���"OVyAw�� ����I��?�+Q"O\���I\PJ�0��0b���$"O$0�UIB�S�rx�)�VW��"O��#�#v�l0k��{D�Հ�"OXQ�eb�w���gɤ.&� p"OP��6eLw��A@�+\VM:�'7�mX��9o܊�
Ƅ~"�'����g�:k*����~�����'���r3}�P�S2p,���'�����+�&5h����EWaJ�Q��'�:q��5.�乲�\�c�!S�'��
FM�w `�&�)H5S�'���i����j���f凶�$Ժ�'��-���W܌��Y�xļ`P�'����b�8S#`4Ѕ��s?����'��ջ���(d߈�1Ώ�X;�(z	�'v�1ʶ=�sJM�p-b
�'�h�B)	3 h�U����=�����'�"�"�MT��"VC�9� ��'o�`Ht�H�>��Q1Vϔ�$�]0�'ܬA9񯓪Y�~8QB�A
&��-"�'Zl�q�F�9���Q�'�1*|�Ř�'�A6l��z��A�(!TЍ��'7�l�@kX1s;Ba��C���c
�'���CC\�`�V�/k�b�@䍍�y"�4!�X�?4v<�)ׄA��y"�_<.	��(�v�jx�'h0�y�m��Dg,�J�f͇ih����T�y���|�pK�OcԎ�O%�y��:)���H=�u�݃���p>Y����~oT���R�r@���{�<�GR�l�@h��-R��X x�<1��ZN�Q��I[�N e�[~�<9b�ʠqe��d�['c�4�{a�_d�<1��D3�X����ߥm��;b[`�<��'�y��y��լ
N�|���Y�<�S��.ku��פ(ߜ8��DV�<�n�IN���.$J��aA���R�<��蟄3 bZ� ",B�-!��ED�<I�������	8�(0;�	V�<�fK�ni�]�ʘ�
^�<��i:�,#�D�I)� �A�e�<�!i�{7����H�j����SǍb�<�Q�L�4�wϏ;PFܡ�W�_�<ƭG J����k"��v �D�<�%�^�Rl`	�j@�Tl��B�;�yG �`+^�4�(D񃎒��ybcH�g#xXp���,������y
� �0#�.�!:�(P#� �♓�"O��f�8l����#�����"OΘib�*{� A�b�h!����"O��qq�G�,�̰ǀN �p "O���=�S��p:�"O,��mX-m\��'��'x�f���"O���t/�i�D��s�ֳC�]�"O20�`�lNb�p��"4����"O^�
�Mʮ9�
\� �χ���2�"O��CwA�4Z�phS��ܵ�v��2"O �k��S�B�c��2�|���"O��tA9#�t�*��b.a
�,*T�r���i��1A��A-Q6<��#+D�)��]��,XSCm��,��c`�+D��YA�:Q���/$�&d�f�,D���a�.���ȑ)&\JD�=D�l���*R��W�6BP8"":D��J�#�sE~Њ�'S�K�8����5D��h���*t���a�@C�P�F1D�`�O�,���if�Luk��GF+D���S�D�J���H������"�B)D�X�TI�2��ڑlI�k�^�Ya&D��"eR,��� �*��@c����-$D��P���mTjT��ꆴW�ę'"D�\�#獎I��͐��;@����"!D��A�g��T�U�N�)ur�$��#D�$j�̮D�~DB2bG ZY��C4D��1� �d~�1;�b1�De�U�3D�<#�L�H�"X�PŁ�t�"��S�4D���%/s�N�����}�1��%5D��s4lU��h	@3NM<5���h��.D�Z�E�n����X� 7�li'H.D��y7͕����5�}\�L��@+D��;�R�j��0ǁ��%m` B��*D��Sp�V�Z��+TgS�;���c2.D����/a�v䨰�R�i��akBf.D� x#aֽVRl8�c8=�\$��O8D��V��U�@y�v��/2�Pp`T)D���ȟ$�����_�T�Z$�(D� �`G,��rLT$h��AW@&D��󂊜�:���E�"Y�~8���#D�0S�A�?h��SH��<`|8�� =D����?\ D��o�%`�hP��%D�бʋ!%.(�	�68|��GO/D�D[0�нI�R����f�`�-D����`�?97 �#`ǁ#GJ!2�*D����ڔ=��bC�3&���g)D���! к[� ���D)߂��um(D� ��hPZ�L�a0D��}�`���0D�tc�Ð -/��w��M��ct"D���Ԁ(I�.��(�X*g�>D�PR��=(o��9���9�ŊW�;D���⊴7`~��$��O�Ɨ�*�!��L+����ܛA�*�v\��!�$X�h����p�ҋ&zb�� f�
l�!�ڄ�  Ȗ�R={Z�Ab�Ɠ�-R!�d�  �F�a��
^@hBUҔp�!�$�]{|dB�HN�+`B41Т�2-�!�d�>N�z�*�͑:EA^43�B^*7�!�$�+2�x0��� $Ah����X�!��.t�XQ��n[X�jT�S�Y�!��%Z��P��Y�!�ŒC�!��3L�TI�'^u+H%"O���v�>?6����
XA:���"O� x��O��+B ��Fk 7�9�"OVɺ`b��]S� R�JG����b"O��B��[���ɗ-E�R�b@"O�-"�nT�A�r� 0)Ih�AZ�"Obsb�Q��*�hڱG���u"OZ��w�&D)�I�)M�^�"O܌��B�Z ��I����"O����	]� (��ŗ<�p�(W"O���FdU,~����� �)�}�t"O���#��?b��P 4��}�v"O�T���B�ʱ�3�Y7f�^5��"O��%!��1
�`r���^� �"O�B  �j�7Ά	���"O(L����7���J0�Ɨpf�\�%"O�Qf"����.q@��"�"O���Rj� 3��Q�£ �P���"Od,�V��6w���6CхބA��"OV�T@	�K#��;�,�b"Or��PDޞ�����
�d�R�B"O"и)�=��Y�J�=�>��"O`���� &(���6��	HM��"O.�k�	B-#�=RҮ�Z�<
�"O��������!���/:��c6"O|�9��l�`LP!WN���"O�pr���qyH=J`lF�u��互"O.(w��.���AŊμx@T`13"O���OT'ER���K�5��"O�%��(l��� U�C�m�<��"OQʇ	�.�V��c�4 ��z"Oj�#��BwTV( b!ڟz���ص"O �	�*�2,�$�aa/mg���Q"O�x�UX�ñ.Q,<��t��"O����aR60���,�F�
�"O\M��l�%:<M���(�L�&"O~-��çH}�MRgkͲ<���iQ"OD��˒�]�	��4ۧ����yr&��`�D���{��e҇H&�yB,:�ެ���B!k�dD�d���y�o7S4���Űjh�@YW�� �y�ߦ����`�]�����yR��0k�콳���djs���<�y�KՕ �>4r���Z�,���O�y��u�
�>>��ǃ�&��B�	�P�F �&M�W*��U'Êb��B�Im��H��P5WfaS@@<��B�	�[��	Pn�3��8�4a�GDnB�	��Ph�t�ɦ=���M	%��B��q!���ƌ˂e�<T4��h��B�5i�H��o�1m,�XF�ǴMfC�IS)X����+�*�33 �?"P^C�ɭQl��tcEk1
8A���!&C�n�|pPN�	O�*��NBD��C�1x9���@�ZW�,r���f��C�	>��YrM��y� �E� �0M�C�	���Mj"��O�N���l4.�\C�	,G�lt��4_S"sGǍr��R�9�|$�V�Q�h�s&��!�Dԣ3�0�@�mܢ�E���!�E0������R�c��=�GΡ|�!�d�8+�BQ���I�'��1�G�>.!���v!����+�!7w��B5�
�8z!��R�7���A���]���`ā%>!�d؏x �  ��B;z����u��f���鏿O~�$�'�т
ϓg"����q�@�q��ш(�|���e�'	6��+�j-)q�C<n�#����/��e%�0<6�I �X�"] R�'��6Q��E�Iyy�'��O&i�Ħ[H�T)[�*��A�2�5D����ԡ"���Q>&�x��1�����
ش��$��"�j��'�RȖ1�=�Ԉ�mY���*V�P��'	Լ�V�'���'0b�ȧF�\:��u��>��f4w	�c�%P��cU �0<y�&���qD �R�С:��T�%ƨЫ&R�W��a��%� gv!�!�	����D�O�m���Ѐ*#�hxxcK<R�&D�t��iyB�'��O��U~RD��I�r��^�lP��#* �˘'Qў�'4R�6B:♫r%��n�Dh�s�Z#|�7-�<�Sę�_՛��'.bP>�� �D۟H(P�%(`PL�1)�J.����ן��ɰ1��%���ֱb���XC��)	�����P�*m0%*�2��X����b �'5ܕ�s��)�V4�DM%$Ζq 2K�}CB*�\bAC���:�������3��b~�յ�?����h��I�]�� D�F�j1"��!35�(C�ɤW
�"�i͓*�FS"��D�ȣ?���ӏ-�e:��)= �مA��H�D�l�����TX�ڪ[7�5��ğH�I���λQˆԫ0�36���h�둘 �]+�@':j������1�Fn��/��(O�5���9f2���ˀ|��ْBR�z�Z<Jc�Z�@�Qgą	1���Ѳ��<� t0�7Ԗ%�p�1A%đB��pf g��'$�����ϟ�'��������daYr*V"	����'NB_�,�IC�g���:sڰ@u���F�L	�-�7f��	��M3!�i�ɧ�t�OJ�	 /����蒭�� �ᐦ&6d��u҅N�4���۟T������Zw�R�'��
~O�8�ݸfsD��UQ�B�l�cގԄ�I�T�F�..�]���G�YQ�
����V�@R�kݕ���F#��pg��&��)B�v����ݎDS�Q�4k>6���g�O�Մ�I4{;�5)!ĕ�9���%S#��C�/�&����P�:/$Z��H�`�O��m�]�I�C�6������D��7��$Q5,݊r��@�OO�|j����O�-K���O��df>iHKЩr�T� �
��KJƤ�`�x�*���i�p�~��6��`��LD�'�;Rd%�"h޵1{^��g�6:�h�aT*A,%F���!�)��S��(�����O��+H�l
K��,��pW���&���	G��\٦ǔ�-b+�ȐC-6傷Ԑ��?���'�@�!+�'j���݂t�������$^�o�� ��s�TF܋]����6T�Nڼd����Q[?S���'�"I��4v_p�&��O���'Gb,���#�>�%�1���ě�����)*��-�*�=p,eq�@�>��c>1���|�XM��/I�_d,
��8?�0�ğd���ħ��O~BY�f��a�d�q�k��A-�IpM>!��hO�-����H�$����n�:}6�E2�e��4m�P�'e;���F�E����sd}M�I�Lx�R���<1�AE��B��?Q����Ċ\���Z�k�0Ox
��b�31�N1Pl3f�d��G�hG�<kpk�|��'BznOf��߾ϵ�&\�&�ѐC�� `jf����ܶ+L$u�3o��n7-�<��Ӈ@�H�$Mt޹�Q���
�P��쟳h�$"0�@���X)O��@3�'���?�On����y����?�`��T�;��0<15�5�^�J�# ��T��mD�x���MS�iɧ���O��ɔSv�)XT�R�x0��j<[g�Y�M����?����|��O�����8���p`^)��k��:[��122��	-c(Q1���$��#?���(<��1%�F�_�0p�\< 5��*`�KYvrdagKM�a�&az��iq��L ���'t���i�;�l;�j	�D� 𴮒 �?�릉Џ�d�<I�OA�am�� R�	V�[p�7X��G2�D�`"0�j��w{�|�V�ߎ?�r����Ҧ9�ߴ��I���z(�'&"�D�o�z�v�v��zĀB�HR�'��7�'B�'����ȓG�	7�>�֋�?Tڌl�$c�( N���g�ř�0<�t�^>-j��pA�2D��F!�1 �VQ��$�T�`���83������	 �Z��O��m�ȟp�R	�q�fYʇ�@$(�&��my��'��O�Sq~��g�a�AiB)>!T]�e�5Ϙ' ўʧ0ț��΃*��z�MF�<��h`���$��6��<1�TW͛��'�BY>c����0���3��e��/uZ��%�C����I�bBd]+Dc\�l����'�?�O�J��pYP_<|��cn�8N��w�\3���4P H����h�2��4GB Lu�B����:q7�����O�$,�'�y�l�Y�p�!��#PBR5A�F��y��h��y�Qd]03)^5�Jʞ��O\�D��+�p��(���*���+�FB�f���':�I�x8�S����I͟��'��=�3㇡j�{�N�6 Lc�қR���&��OtѲ�$M/ )1�1O�)�)�	͚�;u.��s@4�0��
v�>�1���2)E�'fhc>c�ܢ�L���5POPf�rq�O��'�P��蟐G{".��fh����U�Z���ۇ��'8!���@����f��u�N�1'��I%�HO�|y��A�T�R��;.j%B&�&[�r�Ede�����O��$�<�|
�.C�ђ��ڢR�\�J�"��*���ӫ�96��}S6�|By����;c�ܪ�D:W�v8��J�(ՖD��Aڶi:8rt�J.��JEo�'�4��@,�$���Z�v�Ƞ�O���?���?Q����o���U�[��e�b?Z�jC�z `ӱ�"Q��}��#G1�J�O:��'��j�V5 K~����n~.ؠ�DՄ-�@���R��l�'�'���Q�1_v�PĦ�1���woNAj$���f!1;&y��ɟN�Re�C�?���,H���=L��CV炾L+�-x�P�
pX)�E��a̼��'U���O$�a��'�❟��b��>v�e#
Q6X9Z�J��:�d1�O`+u�#��x� Ĩp�}�v�'���Č8pe^u; g�Q�]	�L�N�W�TX�"RDyʟ
ʧ�?!�JZ;_��h��D��5k�N�(�?��(.r!lW;q��+��!X�금!���U��LZ��E�x�P9��mNM���}��OV� �r�#%�وI����˗C,T嫱��7<��T��u~"ѡ�?����h���)� �Y1d*5~�t����:��!s"O�̘&Ƙ�Iƺ�� �L+Sf���I��h��ݢ�T/p������3
9��@��'1����4�Q�`�&-88՛����kA��2D�Xa��ĮArA�@@W�M�tn#D�����
�fh�l��'�#!� D���$��/W����H�<�rh��J9D� (�n�5��(�H�PJL+i6D�PBƮ�h#�<;��1�4����<m8��YU�N�\��xئ��N%0�s�N%D�H�-[�F"����#�&B6 ¢�'D�8a���Smʁ(�fD���Yc�#D��2�U0*��u��8h�M�@J"D�$@��^7<؈tq��x������+�Oh$ 5�O� �*܍:N���Q�v%L��T"O�0y��@"<<�s�ŖF�Ru"O�4�aE�^�v��D$�����C"O H�U�F�V��!���k���Q"O�%�P�Ǆ�A�n���|R�"O<�;�kāE�����NM�&Ԥ����ɸ0p�~�1�N?��mN�F����A�<���`��A�£�+X�Фghb�<)b�
o��d��Al�� zkT�<@�3N��Br�*I��e���S�<�b�Ȩp�9+��۠�6�z���G�<��$�)iS4�b�ρ5M�I�E���di��,�S�O�E
�c�f�D�6���U�LP�B"O���Qc�*k�Ҽ)1�G�J��:u"O4���4a䨊����s����"O8H���ɵL���� �Ƹ)"Oʉ��m��E����H�Z�^�SO�!�d�1I��8��a\ U:N��2L��i��i�ƉkD,Q��1T�ۼZx�x{�랾CET\�XwIw�V;��Hu�;��PLT��r�Rfb�'���?>^  �`3*��P���O�鉀f��)��1zF��IЯ=e�|h��,r]� #�惐I������u�H$|TIb��37�$�@ݨ��Op�$�'^R�	H��ʽ���GH�a��AȶHn�P��4*�/�g�^��@�<�⴪�,?1��T>9�*O��)aAD62H�X����v�4Q��T�� ��������Ɵ̔O�*� w�'\bP=V���>{�0����,9R�b_�s8�P���_�u�j}����iH�Sḩb��-�o�P
֥ɩJKT�̓v�Z��5��S}
�wb�Q����V+�"U����|�r���"�����o�]��lZ$g�<�OIß��Ij~J~��O��Ѡ�uU&��T�_���aK�"O�-Ȧ��h�����]����	��ȟV{����5;�I�i�$�Z��v��O����O��&�¹G����O�$�OV���O:I{T�ܜft��[�
A�wLHM�2$ԬqlQhv C*B���
�fY�=��g�'�b5`�Ne����3=T��Qf�:adV���Z�F|�#cݻ���F�X�DaW��0Hb+B�&B���6bL����3 #?��m�П��	J�'+�d�;[��U�g�ҊN@f�;�Ȝ	
!�*y��|�W��)���Ǧ� 
��5��|"��򤃌EԌy��-5�5 v"�2"����'��Q$t���O��$�O��)�O:��v>��d+R<H	�%�b�d���@bʉ��IBʋh��!�ɃTSl��d��*;��A����6���i���/W\j�8F��~ 4I)A*�r$���6cۗs״$yT�I%����ҙբ����g�q�iRY��<ړ�O ,�����*%�re��P�6,l"D�$�$ʠx����?5	�S!�<�i��^�$#ӫ���OQ�E)恚p���Q@���V$;[�D�I���	(L>�$ C ��PB����-?'��%3e��F<�,\m�T�c`�=�~����PFR9:�z0�|����g��5A]w&�ɣ����BU�����Ke��p��$�7y2�'�1��0l�*(�ܢSm� 6���CP����I�]�����HM�ŀ�k[6Q����F��O��(!�U�Z�se���˓}Zޑ���?	/O\�'�?��3EB�ɲh�:��M�$�SO�,����$�x��0j�<zzmYgIJ � Q�6ҧf�`����E�Zp"�̣GRx]�g0 7��<�F���'0l�}�铀XV8DB ^2,����p牥���O0�S�c~
� ,3WI�%.�����k,���"O��(�#f�x"��vz̨���4�ȟAPEA�kY~��̗!l�X����O.��h����?����?�(O�)ś{�h 1&ͷk���tM�ko��f,J
�\�o�3X��ɀ��?倍}���	xH�;FnQ�JY!f� �`�xa*`����͟�m�>i����*`����^�m����DFJ~�e=�?y���hO~牦�8C��N�m����`�nC䉫&+\�;ӋV�F��a� �XF�$
@���T�'>�I0^�:#�؜V8�	�K�/zL�Ћ&T柌���x�Iyy��T/Pj�p3��цp789�����o�`�J#>D~��8%�������t�'X.�`�ʡ�`��5?`��W$ٚ#�M���k��гq'���E�		x����#f���O�aN�1dO2e����4ړ҈O��A�%Cf��B�`˗l4UÀ"O�(�c���_�n���.^���]��Aڴ�?�/OF�Y�*DҦ��	� �')qQ14�-+] ��_�NQ�]�	6C��@��Ɵ�����7��^6�'��͠+?$	�� VX	�RL�L���w�C?RW�d��bO15�Z�	� s$��27�a63�*��	�Z	�F'�_��u����p[K|"D��qq\R߈L�Q��ڱ�?I��������N��L1�OU9�P����h����CĦ53�49���(��&ZZ@�$�ːt��a-O����Of�$�O����|B�����/E��Y�EcY R�������by�&�2��'�ў��`�8^�Ր�P�i�xp�c0�IN}�O�b>��F$=1W�K�AʌI~����מ�M�c�4H��'�<�"��?����?��'g���!���[`J%�X�� 8�UJD?�f�'�D���'��d��=H���u7@#��W���	q�^�&(2!#!0l[%
�O.��"!AP�I�����?9���?ɘ'f
Y"����j�鈲xۄХ�?Q�M��Ls��y2K�?�����#�O`M���U`��)R1?tJ�b���O�Y�'�r�*�~�'�?q��J�}�r����Ǉ' ��I�n��*��'�jx����?Y��H�?��'% �+��M�;O�N��n�0�)!	I�%Q��T&��L��=O0	)W�'���*��I�O(�����y�6�?�L ���}Qz܀��<n��I)����Opɯ;�?9�'O�I�q�Oś�_��ެ���B0Ѝ�c�9ξu2A�'
�D����'�֘"˟ ��O@�I�l�03/������\����X�� ��X�<�qk�ҟ����?i���<��/K�|��HO�IG+ܵ x��e͜�M+Q	��?�.Ov����I �'���O*aQ�+tm8�DJ�d�t�+D����*� ��,C��7� @�Ik� ��O4�DZ���P�	e�ܴ3�A��HF�3tL��ۀG���l��D�	�H�I�����B��~�0ryPx� �pv��d�\N�<1RH=R��5��MBL��Ӂ��I��?�Ǔ
���z�`?����bƺU�Y��D�p{�.Ֆ(E��RI�7=<5�ȓ�:LQI�7�AʂL(O�0��ȓ-h�;�$��d��ؑ�""���ȓhn*�*��b^���cӷ$px��4T��%� >�!�X7 >����.�����@�Rl���H���܅�3�Y���4W̊U*��í}�l���N�YK�n,��C$�*![�iE~��'ZR�'XB�'Ђ|(e�u�2��`��&)����V�s�f�$�O4���O���O����O���O�Z����7�L�� �YK ��`�Fভ������Iҟ���ɟ�����l�I̟���섘 �DQ{�
F)	ȩ��b�M���?����?����?Y���?Y��?y��6Q�4��&%/�aæh�~ӛ��'b�'���'��'��'�����v�B�N��T����Y��7��O
�D�O����O��D�Od��O��$ݎ3nr���Y�P%�7	��wB�m�̟$�	�t����<�������ٟ��	[�p	)��V�b���E΃y!��ܴ�?���?Q���?����?����?��)��P�V�s�ui�fS�M�;��i"�'���'���'r�'e��'���SQ뀘�.)�.V�5���#w�|���O����O��d�O��$�O(���OH �e�y{�H�$�,F
��*G�Ҧ!��֟X�IܟP�I͟�����(�Iğȸ�Ŀt�����OV~u���M����?���?����?����?���?q�n۶2����n?t}V��iB�U͛��'���'R�'��'���'�BA(�x�32��9!���L6�8?����2�$b�0����-*q@P����)6Ydh�4^�f��<���tn�|��yX���m�=�|�b���m;�Ms�'��	N�6Y�r�mZ@?ec�)~N�	�&[�_����To�ʟ0�箛�u`B}�Ul	_����2Oh#�mЩ0�x��$�9�>dc��'���x��M��K�f�� ����j�13|�͈mU��q���d�p}�Ft�xoZ�<	.���D�ľ�]Z�Ʉ�
����Q���v�qú� "�.?�'蒕`Ywu6才I�X�Q�*��f;L�3��B�#�"�����O �}��{��0g��mS���!@ǀ1Lp)�I	�M���GQ~�m}�H������+� Zc��$9��Ł~I0���	�Mt�i\2,��*�����9�KğzC������=���'F-���@nH;ɠ��C�I��'�1�F��!�ۣ9����a�R7-�$�W����4�`a�<���$	�2]�`PO�i-r���,ݎhqx�ӛ�gӴ�o�OJ֍ɗn�6,��P���A�8�g���
U:)��OJpqO�*m��ݖ����D�u��AH�A�)n:��0� ~)\�d�O��$�O��D�O��k�&�0�B(�ZCK=�B�6��CMb�|�p�OP�lڐ�M"�'/���1����E�'+W�#�v�(�"8���?�i�U=�h�Q"�����|�]�5a*�!���u�: ���>tf���O����O��d�O��/�'>������X�s�A8tz����ڟ��I��MÓNK���D�����I^~"#�$�P������@�fD� ��W0�'A7��Ҧ���:���Ҥz�@�	"��L['>'8�Ѕ!�
��D
���~L��Cr&�W�fy��'2"�'��왡��%�2l�=M����當�"�'�剖�M����?���?�˟`Y۳�D�L2X�YU��9!mtx"W\����OZ�lZ��M�`�x�O���dZ�1
L`�2h/"�]yD%U�.�հ�#[�����W��Өgg������H�I�w�j��	�j�Jcۃ��(�I쟠������D�kyRcy�P ��L	aA�֢'����b��7d��AI�]�0)ڴ��'���w˛�	Ċ5�\�j����.�tCҫj�V6�릥�F��$K4��៤b%�$u]�$��%�[y�(�:�F�2���\��l�̇ ��]�x��������|�	���O��l�C�M("Y�W�רU���B�i�z����'�"�'x�O��{����>wT�I�`6*�y)'�F�zL�o�
�M��xb�O��$�O�3t�L��y��AC��s���x��٨�a�#N���Q^��J�k��JP�'��Iԟ��I&S�!�LِG0���:p4�	ԟ��I��'wb7�#R���O �D
�]���+bMĒ:�e�P��7X�<��OR�o��M˷�x��D����)S���Gv1,�v�"�'�h��$���ތ`y7\��S�I`�`r���<��P[�$}����3'�fh;$�˟@�I���	�D�D3OpE�f]�.��P�kR�����'3�7�̣ig~˓	���d��b@Ñ�S;�����]��l)���OPm��M�!�i6�S*�yB�'6��څ.ɱ�����3&�ai� �6.έ+Edӳ?��'�����Ο<�Iݟ��Ʌ>Z���,Ɋ`R �� ����zUZ�0(ߴ,b���?����/�󄜍%.J,���MY|u`�>���'�7���iqN<�'������б�]5go^M珉!u,ݺ�fу^�rY�,O���Tj�Twv�bg�9�$�<q.��:9(7K�Qexj��2�?���?����?����SЦMZ�����aL� id�L����^�<A���؟xq�4�?�M>q$]�́�4H��&�O�4B�J
�ȅ���7R�$�lM�+�乘'���L3{p�!#�	
���?��;(�R ���̱�x���FXT�X�Iҟt���|�	��L�I}�O�X�9��)R{V��`l6C�Z�����?A���f���	��M�y"��'Qv���-��)!��0'�L �'H6]ݦ�Sj"�P��$f��I.'Ѩ��H#-CL�ţ�`��Z���c~,�b��r��ey��'8�'��K�#�,Y�dL�V�� �߳H)R�'x�I��M���O����Ol���0��g�7%N�����
�F�> �'��D��� `��$���?�Z��5+�n�s�mL�>#^��w���%�0P�BǺt����'��	D!��mC�|�IN*$7hI�n�"�{�H �fB�'�B�'���dP�\�ڴ-+t�����7$�)���=VJjl��B��?y�d֛���r}2KdӠ�u�Ͱ��q�iӠs���K����	޴>-�,�%�\�<���%�Ω���N�p��.Oެ��C�i�V\PB.�n��h�(V����%�������(�靇_���I���A�qC�y�H�"lɿ!%6�CZ+~�؊��7D� �U��H��� �!!\���W�x�kDI�B�q�@ňBd$A��	��\�LAy��=|�Ȅ��C�(Qz�JP't�cС�j�vص��M*�$�AQ4%Ι6mӏ@0�r�N�FYc�#��v�,ɐ�P.gք�fP�Zx�h���.p��EC�U���@o�h)��Zݰ<�e��0�^��Tʀ)d�P�t"�}<�v�N=�������ca�0��T�6��1C胯g[�yY�
�1�(��B�)�V(w���Y���sQ�"����툹H1~4�WJ�-�p4��j�6D�h�bDp��0���B�B��a
<=ȕ�B	f����@-N�&Ѻ�Aq�@'Ϛ���{!�:@

�j��ٶz���bش�?I��?y�$�'���'X�DU�J�5����Y���$�K<�O�D�a�'���O����O4(z5,�'U�ȅ�D��15�zaA�ON��:{��%���I���'�����P�&���­�4��hU��Oy
 �bR���I͟���Iy,�dN�ȣ&�ּx�����_"LK��2f-�D�OT��4�d�OV�D,H[N��t#�?W`��FG<
Rh ���O���?����?Y*O<ܨӅ��?��bW�G�	�v�\�t8hS��Ot�D�Or�D%�d�Op��T�g_V��7� r�P��G��q�	�1@$��'�'�2�'��I��Y۴�?����� "�#eɰ�Q#Qe"ఓ���?�.Oj�d�OH���)5p���O8��E?m��BE�ү	�Hk�*@�8���Ob�D�O��9bH�nZ�0�Iß��f�t�ʦc��= ���@I�/�|��?���?�2�Y�?����?9ϟ"	UK��l���L���\����'�B�'�2�1p�eӂ�'�?Q��o.剙"N�آ�_�O��}A1ϙ?c`J���O����,yԞ��$��8�S���u`t̓_����G�p���䈰v��dlZ���	���S'�ē�?����\���>_��pр�^�?!L2�?�M>��T�'`�z��F�˒mc�����<)�bf�T�D�O~�D$
��$������ϓI^��@��I�w���GP�?H �IJ�7nڎ'?E�I����P#��'��v�V�c�7(H��ӟH�P����M����i�O<ʓ�?"�	4���X�� 3a�	�?���0������?1���?������O�!S�u��H��)I�r9L�z����|LlZߟ��	ʟ\��Kyb�')b�'�P��%��*Ȧ�´��^��t�$NM���'�B�'�Y>Q�	%M�*)��m'���a�փ[�&4� /^� �:���ߟ0�	��$�4�I�<;��^���� X���!�]'-�,�q���\��ȟp�I˟��I埴�4\��ħHR2t��q���֔�"�Z%�?����?�+O^���O����I�O���Z�sW.-{^�q�sÍ�#^N��I��x�'#�&�3��џ��	ؼ�Q��:�L����m��l80�Ml�I՟t��,Wa�&�h�O�mS�A�+p�D⡬M��Z,O��*b���O���O����<Q��\&k�J�r�ѫ��}ZG��?���?� �l���� ��� $�P�X�A��=��4�0�'PT�9�'1��'���O��)� ��0?�4Li�����̃�f�=�?�H�P��h��H20T��2�D�8y�-*��	�R�H���O~���O�h!��<�O�I � )�eGX�� ��Z�2�O��dB�O��\���<d$G�*	���í� e�`��ٟ|�I*�D�'}�z�l�y T�W�Q�:L��)V�q�������?���Wq��?Q��?/O�D�D�Ol
��0��4qԘAE��-}�\%�4�	ٟ<$�0�'=����	�$?.H۵�)¼��k3��|r�'����8���|B���%�"q�VO/s@`��ӟ4�	���?I��?�¤Ϫ�y�ӎk� ����
i��t��3��$�O���O�˓+*�᧖�4M�+�X���>쨵!%�.���'��^�`����@Q�n�🼖O��Y��B��G!*��6.��	ZD��õiV,���D��ցC��ʋ3��#4�Ǉv�r00g�=n0�)��P�ā�P�vp7l�76��c��O��7���O����Ob�O�l����4�������'`l`竩<���?������?����?���1ih�k'D�0j�I�(�'�?a�����?����?a����DY:�Ԩ��/ܷ\�<R�) $B�'����'�z���OR���O�OY@�T�l� ����2YҰ��Ȟ6X�b����V���:G��>V��:R��#<q��
�)�d�P��<��D��VH�<��́�\��I�N;z��@��n#���iE�ß:���7�	�n�>���/��H�V,	��I5f���Kfm7�x�!� 8e�hR](2ja
p�/�$�sgI�(Y�Ղ� �+@�P���M��(�Z&. ���Ǎ;�tpk�E\�JW��� ɵ�N�:D��y�*} ��J�9�'���'S�ם����	�|2&�$KRR܉$�ʹ����F�"��'�z"����'�>0�#��85{~��i�dX��茒��׼�B1�eH y��E}ªN�S�x�ATˑ+K *!��eŶ������?��?�(O$�#�	#,Bz8 �܎���S'B�^�zC�ɍ,�,�@��T�~渼 4(�v{@���۴�?!)OP���dOߦ���Ŧ!��X�(�ȣ��*9aH��$��?��"ﲘ����?i�O��U	񮆡��BQ�!�^h+eM��"L�ܙs �Vu�@�<,O��Xc�i���Y�z�f-��� ���(uFG�E?�:�'�0�ay"j���?1b�>�po�% ��Չ���4u���c�l�<�'�&O��(�G
�@�М��%k(<i"Ӆk����`��.m�n�i6�˕p�B]�N>�GDH�s����'YR_>u��OC��Y0$jP�Y�����	�e��|ff��?��$�^�p��ŏA�Yh�L\�^�*���I�D����J���B�e�j�$�L F�ҿ<�52i3���D���[�/��`Pb�A.N��P�銆��_����I���S�<!�`@�L����g��G�����b�lܨ��M1G(�@��*I$w��)��	9�(Odt)���#7j��+�A�>s$�6�I�M+���?)�]����2�?����?Q�����2m]:�^ [rfK� tSPD6���j3mH� r��*7u�����L<��M�6)���l��`�$@�Q&����O�	O�T���P(��~&��7*�r�h`����;��#g�.�ɧ-��S�g�	�Z;�l���\$�A��&MtB�I��v�8�̓7C��Iz`G�+^��'y�"=�'��S�? ��తM�K��!$��>]K��M�z��ѩ\ԟ��	��P�I:�u�'b>����C�ʳi�6M��F^��N�
Č�|���ߜD1�CoJoX���-����4"@ԣGF`�F���:���:���
�l��JX���	-"��Aq!�P|�ո��JOB�I@��O2,l��HO�b���d�@�tR �!(ڔ��H�v�!D��� ��v��0ɰ"��CD�L�4?�	��M�������n���o�4�����&i;K�!���1��ϟ8��;t4���ޟxͧ{��)nZjc&A�𡟄�F�R�@�=i	�!��A�))$�:,O��S��i[��	T"�z���q%G�{'����M-9i��A��(߰<!�������K�p8G�ˮ���r�O�+j�T���(D�Zc�T�'��`�'�f2��Ydj&�P�B��4�h�#�hB;5QD�i��_�ih$�@4��M���?�.�R�ɒ�b�dyp��?{���@���-z�9!AFҟ|�Ir$dA���QrS���' ��S�d�\7,1�́�lG�(q���ē)\���s�6g�cH�8Rm�c%I~��.���J]'0�����4?��OJd��'��7Mæ���E�ߟ��1D��,q�!D�5���jp���O��Zz?B9i3dݖm�,�(���c��xk�jeoZN��$ʎ`���Ԧn���Jw�S������?����?Q�����T����?I��?٠��U���t��� (B�z����/��Q����z�e		�����L՘O��a���0��
kk ȶD\*&�� p�S=�j��M^'�R�ƛ=ni@K?�26���y�CD+�D��E�Pv4���bр=<��l��򤄮��O��D�ER�0u9���x����$kǬXo!�$���Ե;��٪	p@�"�j֔m��*쑞���Oz�f.X�U���B�c� >��c��`}h@��'q2�'K$~�Q��ޟϧG��|�@FZ�.w�5�I��F ��Pp-�>
z�`֟��=�"��B�0��v�U�%�[�;=��*��Γ{�|鈒jT.hV�+��� O�A��iú��<C���2�	u��O0���	%j(����X>-)v�����E9	�'L8�P��+G�,`�"]�-�{��nӺ�O�x�o�ݦ]��Ȧ��a�C�<�и ʉO-�'N���?I��e$����?I�O�J`yRf}-@��d�O��iA
�#�h0�Ʌ[�>��E�':��c�҈<�b���� AH��t��%̝P�o�a��}ku��~E#?� �럌hN����:P��T
�jI�	n��.T��+g��>
���HZ�;�iU
O"h����4n'ڡA�B��<��iI'O'8�O�t�1�Sئy�I��O��I� �i��}�Ǝ@�3/VAiC�+m~�%�0��Ok�i�8����z�1��Mdp"͇B���􎔛C����F�"Kz����xBi��v�p�rF��G� MssjX/�,�����,]���	�]�{��	 �E"t��cGb#+O:tY��'�6�����x�c�
�h�"O�-��田-���=I��<��@��,hD8
�D�,88�2�.Pd8�\��ă�p��%ڃ��T+����B����4�D�O&��Ϸ:����O�O����O��^8g�l\c��՞<�&�KD�������"DW�d�:[u��8w�x��:y����O]�}kn���]�8A��A�����t`��9�%��L<�)AV�\)�
�;i��h���nd�O�x�����#h@ �aA
TF��b��*8ȩ�ȓGf^m�E�Y���#v �sdv�O�Fz�O�'}x@Ka$p�YK�)�D�b���?%pp�5!�O����O��B����?����$ت��M�1��Yr�;XpL��T$׵\�pـ���{r�F��1S�c�VS�0���S�\�*�{���aP�IB� 3[���PÓG�\L�Ņ |���PI��D�T2����P������gy��'ޱO(��")m�(��g��b�n����䁎��$$�Xqg׾K���CE(	0V8񲯂�	Ɏ�'�6��O&˧�?ɴ�iYºi� �s␀eD���"���^��C��O.�]���D�O�����Q!�ᨲ�T�&��Q�0)b��zTk}.ِtCBBX6�'��ȳp,�q�0���M�/٦p���"MW	���#G�SX�49���O@�m�/�~bئJU�<@��1L]�PDǥ�~r�'�����OzO�=	�n׺X"4��cT� Lِ�T����_�X6���@Y�zc��h�&��&;������C�bT|�mZϟ���ӟ��ӁY-x�l(�B��XN���A2������?	�	�?)�y*��ɘv�fu*�`ϋ~@�;�)@b� Or<�4�)�������%��z����� 4�Or�%�'eR�O��`|�7��*�:���E�`9��"O|0��$ūJ�1��?�,��v�'P��<���e[v�Itn�t�cҭ!E��6�O��D�O$89d�*HƢ���O��D�O� fePS�T>A�-��,��8b�iF����剠q
9�(L�`�\�֥��_�Rc�hP'h;,O��:�	Ų^숄	���Xx���L���Xh�)�3���&G�VŚ"+�9c'~H+;!�ńTJ�-��Ʉ@D
u0IǕ2R�v~���?��UF_�h��b&� �?���˼:���Kg���?A���?)��j���O���v>Ec�͍L���n�$0ؒD���&ܨC �8�+P�'p4]�ah]��)�!@Q�r�"��ڮ.�e��G^�+n�A��I�AJ�T�S���F�4T��c�	(�$�OL��I�)��)Lu�Ҙ��ē��lC�	6Fu�Pk�,�%z��8[�nݼC�:�P��}Rh��K.6��OZ7���6�=��ˋ
c�#`m�0i�(����L��C��$���|��a�hQ��c�*^��D�wun02��#"̳ӬNz0ay��u�������ɿM��4��bW�]�ʌ�smX.ph��ů*��:}�-[�>�b��&=���0!��y�jS�8e�ȂЍ� "�0Q�]��PxBFV�����Yn@;�� i&u�=��L��6����'��T>U�h��ٰ��=E,,���N��)idG��?Q�tg���w-��q���#�>�O��SL��,H�-2Mm��s� B6�OT����H$��9r��D�O��Ղ0xr���s��p����M<i��V���"I>�~�gn�<Z�1�d�� u�*��1O�k�<Q�iO��f�c7c<T¬P��+�\8��a�򄄻ݑ� Z�5����H +m��3�O����O>*CB�=�����OH���Og昝)�ti��M1Q��&FRA�so[���z�'ܯef���a�8�S4����,����q+�n56���ޡF��\��k�/����E�N�+Z:�#w�)GO~�@�w0
�0#�%)���2!LA�.^�nZ���$W	a(�O��3����b6d�K���B�,�!�A� �l�{U���tJ ���JT,+v�X������
���s��:1$�"j¼b���1o]�29�I��4��ߟ��[w��'��I�'�V�#���_�$5�&i�B�(�kc�i�g�<|O،Qѫ;�ᢷ�ԣ1�d�`�L������\7C���#0LB	$1��"�	E��"�e��A˺���9t_�8x�����=<u�0I�"Md��SFN)Zdd9��>�t,{��T~�hfLK�l�*��=�Q��ԆK�x�nZ�do�<J���bn@/)>��z�d�#��c��?q�o�)�?i����M4��R�b�ji��A#�p�� I��_O� DW�y 6���Z!_۞�q�脦*���!g��T��U�D�����f�>�a����L����v�d��R��Q�`�E$_NĈC�I�)8�!�dX/
��8�\�jI`T�iҾ)֡�DQ(:�ebٖ1c �(I�)��B���p��?�Ĝ#2���l����IQ��N����V��0(��0t畵qh��6�4&�����O~Eb4�*^���b�F�k�M14���qn����~��iW}��(�G�/NI�qQD�
R�I#h�ZP��jW4�u��V%*��ƩG����ۥ$�,�8s4�lC�챲�x��&�?u�|����>G���s�H�^�f]�!�B5�y�![z���2!B)[��h��-�p<���	>*i"q,Z��"ʀ>m
ʡ���iF2�'O���| �EYr�'�b�'��;p,"%Q�)�5L�d�@�f!΁2��L��]Q ��O�U��3p-1��'���qCٸ�^l�Ņ��Cՠ��R��0%��ܣ
H�R|��I������_��]V��-�Y���Ed����<���Eǟ�>Of42�I)Yw��h�6���r"O�}�v,�W���f&��fp�,�5�>���)�S;m�T�!��+jd
TeJ o�z��Ri�7h�����?1���?ױ���O��ċ5U^섊CJ@N�`� �9.��}��i9���
�qX��!�T�%j"`%ױ�THpC��(�U� ��b��C2J� �D|BŔ�0"��U�@��P}�B�}�������?��x��'���DړG�TX�@_�-���#� ���d"�O���'+�xݶT��n�e��9�{���M[6�i��	���D�O��`��"�-!fF���bC��y�h3�X��!�H"M��m(��H �p=Yb��%jT�Q�( &[��qW�ݦ+��bT�U�m���<D��*�B��p�Ș�B�/0d��)D���w��
s�\XH���/�>�CW(8D�(K��[�f�����%Y��X 
4D���t�H�I�a���rk��r��'D�� ���%R��Ȅ����?m4 �"O
9;r�&|��X�W��4%8"O��Zd�� �FI��e+^��"O0�s���S��T+v*�@12�y�"O�h�f�Hx���S�ʠr�H�"�"O�<Tcƨt�<�������A"O� �7�I��5J��!tje��`=D���n��ze�)�5� �N��,D��� �3pR1HQ־�ʱAA�,D����BJ	�T�کJF�ߖC��	��I�i�z}�����t�C䉋gH4(�K�/X�PT�6,�&C�	Q'� �w��n@Y��H�Z	�C�I�iV1���A��7�mz�C�I��p#W#ͺ"ߤ��4d��LG�B�ɵJ�L��oN3L��r��>*z0B�ɝ?M��Y�l��E�H���Μ?l��C�	'}`zQ��S>=��Mh:
C��.*inԛ3-U�E�\8�V	Dd��B�I%����Mծu�T��O����B�	����q ?�T�y֧�X��B�	�A�囷���Zz��D;�rB�ɪa�x��F�@o�L86K,X�B�8:���e�^7ovL
��-0*B�I,<���U�Ɇ8��������zB�� @�N�Q�ơlr��q#��Y��C䉯)��4Yu��|A�	p�J-FeBB䉆rX����ݹ(X��Y�CH�mB�I8Ҡ�+&�[F���䇣.��C䉮L@�����P�!�U� À��B�	�n%*��(�8 �5 6��?�@B�I�9q$Ъ�N,:�R�qD�zh�B�I�x�~� ��X��� �M��B�	7B��8�V牛dbrd32i�2O�B䉠s�P�N�	�@|��ǟ;c[�C�	"�F�сa�%�dMs��Q�#q�C�	7� "�) �Q��"@@C䉊ڡ��h^�["��� ���B�	?Әlq1��ij�9���&IW�B�	�iPN(+� 7swN�kOԵ[�C�#��(��т}�t4��LӅ����βM0���'
�1AG�<2��9��-O �`8�'��� V���9TI�B��UʊR��2KZ8�)	A�O0�������f����=!��b�'j�1�v� � ��L��1(�����2o��H�I !�~rnG����1m�.��1&M$�����Vx!�$R:>1/W�0ٓ�Ē�Bz\�iݟ��1�ĩӼJ*�8��'�xh� H� �^�S� �6�
�	�f,�9x�ͅ�uf�Ȇ�^�>Eڀ���?���+���l��P��'����cl֣2�$�J `B2�=�H>A  B�}4���Hʾ=�l-2�o2���M�NA��H�d�X�-	,_�C�I^����K�'G��I��͉> �dȑq�<k��aB�,^�)ޘ�#��&�3}�H�7�H�#@�6�f5�`OR���x���=��CV���fM��';RL��a��`�F�rp �m�Pj��'Z�ӑ	��%�J�'��<���˓GH�PΈ!`C�a
�q?�IZ�-7N�M�ΉduX�\$�Px�ڇD�^�� ���Imt���c���ē{����a�/,�a� (Љ?������,~� �R��E�~q&�	3I�yb���"n����G� HIȒ/P4Cn)Y� ��Jen� �d�-�Ys��4�>��� �2�0�W�%S Y��uH<���0"᦬h#ӴM��u��M;��.� <.y��YX]ظ	Ǔw�4K�ˁ�^%H}�&�La�.���	�`�@������qPe�Nd����mۏ>h�A�J�gL�Z5��(<1v@U�ln �A����]�tE�a����*+zU� �K�F���-B�>�t�}� �qDʢ:��Q��nZ�qR�Eˠ"O,�F�֕9!��	�0��!	ì�k�pq�@�͞���4�q�O���ď�|�b���+A5�<�"
O Qk�F�;�L�Hr�C!N�"i8!���gk
l�sN�#j&8�$�҇Q����]�ɡ�*� ;w��g�;��x2�^*r����7b�N|�<����v�b���mJ�j�6y�t�^�0�q�OιP�/�1��x�� ����>�����?8ԉ�ƈ:��e	�����O ���!Kb�&�� 뜥ip�PZ	�'De�5�Q�f�&!��l�U Q!U^�M"��R#h�d���^���OF�'�V(x�E�?��Q`�'c&~x 	�'*�ʅ�׿G<�up��Қ8���$�]	^p�3dc��2>��3J��N3ay��[�-f��SeR4.y QN��۰<��'��k[�d�l�u�:`���F�D"���n�	Gt���φH�lB�I&u	b�DM�7��M෋�?_q�Oj���ϗ�|��X�@DN�C�����DkV N\�-P�LEg@Ԝ�@�U
�y�6q6����kG<U�~�`)C��j@C�l�|�K����8�É�L<�0i��	;�&H*O�H�8l�I(<�.2JH�h+ri�V6BP8$ؚ5��˴'�P���eR @�K
����լDo^�8��<2��	3a�aYs(�U>�T��,;�D))�h����M��Q�5�IʤHTR�H��Z��$E%���A	Ϝa�{�@�h��9��Qv @�ݾ�Ȕ�A< 푋��b);�X��v�5.��gBg,,���)�Y��8Wm��x�.,l���y�FV!v�H骀��s���6ș`p�n��I��0}��U�_f<�÷| ^ݰ��B�Px�J��$t����[�O�p*`E�0HÅKer$Xp�3G�mJǂ6~�(�[��(m0��<1z̩��շG�RaS�'�r��Q��R�-*5L6N<�f�cX��v���}�b�*��2To �X!�(����Ğ�qB\K�oV; �rt�d۰��v�����O�d ~��h���b��Tȇ�>_,�Ti�d�hU�"	T"�v�ӃE@R����F���rb͞<H�)����P(k��(#P�����l�OVH��Óx� Ĺlt��P�m��]�$��t���s�n�����e��)O�ld��	�Nh臍C1,���O��<.�yb�ی�,�y�E=AL��3�c ��<q���CJ�������U�h����D�Ƈ7�."mܵ�C�	}!� �V�Z�'���y(}sʓO��a$�_�v���G"Βng�#|��)A*2�f͋J)T�W�X�<!���eR2���)4�u�����S��x�@� �����NW�"|�'.�@V�L��/C4]���k�'HH����?iۢ�h���HSmڴ]���4:����,T`U�B�>֜HW���hFa|��:B4V@��R�<X�$�	%����!�4�k�<���_L�@Po��p��1Ũ�}�<ِ�JB$��q/ϥ(H4�Ј�{�<����'w X�Ӏ�\����~�<Өē8�lJ&F��_ߤ-Wb�C�<I�k���J��2�w�*B>#7�C� \� �UJ��8D�����B�-�Z�tΝ:l� �)۩x�B�		z�HQ�Pc
J�N(�PlO�q�C�ɠt�,�a��-;ڞ���,�&(0B�I�E|�K̟$s��1dh���C�I7ݲ%\�d�@���@w�C�O�.��$#�V�,�X��J,O!�C�ɿ7d������?[_ex���IglC��Sc,1�Չ�ȸiS�R�xC䉧K3ց1o$1\��Q MW6+?�C䉔X�H��g�b�
qh�<JvdB�	�1'�� U��?#��,Yg%�62B�	�8���M�+e�@�6�-DBTB�Ɍ?ͪ\�!+��}f�HC5O˽6��B䉐�Z=Ȣ,	\��!�/��C䉜Q:2��ԉF.b]�DrE�T�C䉳H�|x���-^�@�>�B�I�x��������i����2�ñG��C�)� n\�i�l�$�� 	n�s�"O�4xG�]:_�4�i֥�;�T��"O�e!�bJ�h"���
��q�"O��'�B�8z�
�"�~���b"O�TQs�,ZIJ}���t�H�"O�%Ju��*8�D��녊]P�*�"O$i��eS�Z�����W&MY3"OZ�KG��15�)1����(M�"O���q�M63$袗"N;H�.�p�"O�xZ�KL�~Mn8a�"O)�0r�"O�I�v���2��S�w��(��"OԜ ����s�� J�$�3��"O����H�*\b�#"�a�"O��hż��|�
��%$S��y���:A�ra���հ `������y�뜔�ˇ�&	��h���y"   ��Xta�/��l9����ybl��t"�i�K��Q|�t�	��y�:+�q�c��h=c��#�yҤ�|���,#B9k�gޮf�M��g�m���.(d H`C�=�´���h�S��G5���W�B>g� �ȓv�
a��D@9�2B��q�P��ȓip��G j&f� ����YH.�ȓ05Hp�� ���G�ɞ\L�ȓN�&�X���j�,X1�c� d���*I��҇B#�()Ҵ�P�ȓn�����,Ǐ� t��]�[��p�ȓtz��`�Ŝ�B#ȴRqą�(�ȓ|� 1�,��FG�4�U�J N�����f���6 ҶHX��T���XH��3L��u)�R� b��Q�~����bT��qM9;�	N�F������6nX�z��ɬȸ"LQS�<Y�.��(]*EC�J`C6d��r�<�#�I�i�k�a��I'"Pl�<9!� +��؂K �q��Q�HLn�<AW�w����)�Q��MI���o�<�3N�'"�9Q噔[�.8��@�<q�#��P�ID�ս-�8h��@B�<!��/�"̢g�#[Rx��s+�x�<�b0%� �ig�C�~����Q�<���ʇJ�^Pk�E1<�v`�Lj�<�)G�}2�a�4"ě��0�̚`�<����ȗu��@�S^�<ᖫ��
����
�7G���`�RX�<Qs`+q�8�QOZ�H��I��-VH�<1��׬\|AA�(��h�ڈ#Vn|�<�k)�P�gB�k!�0��/�<��o8/�\Y+GM��4)0���<�eA�(D8B��K��2�jQ��z�<1Z
	��n]!�H���		�*�B�ɑ/��]Q�@ �"�$�w���Z'�B�j��ʰ�G.s�� vΆ%*�B��2�61(De�"Z{� xьDFYB䉨"@9b!I@�rv�LC� �B��C�	�Sr$�y����7��q,�<,k�C�I�=��z�ᓡLMX�ӣBΌ<�B䉨Bʌ9#ܻ4��M�IX�C�ɜN2b��b^�G�> jC@ʆ<�rC�)x&h��H�J�Q˖NzC�ɨ)�򭃅�D9d�bԀ��_2xB�I/ʈ � mK�_�@�iRm��J\��ֶWq�hcA@��n[b���|�x�(���T��!��K��y
� ���@�u㆕ȅ���Z*T"O�qS���!B��;�%�=``�b"O��YB�bI.�	�&��\��D"O�x&��21���8�-H�,�"O����&�z�>d�g��Ő�ZP"OFt�q��xhe�JO�"O&a*g�"N�N1j�O�T����"O�Ip-�;of�q���);�J�"O�Qӄ!R��P:�$̜y���"O����:F��gF"h��D"Oty1mYt;����K�=kh(&"O�H��ϐpI���K�:T���"O�#�͑>#[��x��/l4�!��"O�5��%ޱ#�
3�뒩Z�l�Ku"O���a>�U9􀝇1a#�"O`����:8W���b>HA&	 6"OF�pF(1�@pD�H�����"OڤZ򢀎OF�Ҵ)V;)�=h�"OD�WG���ʁ��o%��$"O�8�wd�5d�>}�qN���95"OV�ÔZV"��F��Sh.��"O"]��ڐK2D}@��H;NJ]�"O�9�gi�,~���K��O^��"OYb��0W/h3��@�N�\��"OM��e��4T:�O��bJib�"O���A b
�E"MW�
�L��"O
��`	�9�ʌaEY���6"O��V�ղ3��y�篙%?՞`!�"O2m����6kiZ�*��S�8L�"OJ�(U850�Xj��Ў"�4�9�"Od�5��$<&���kA'��(���'<~,��,:8�*�c�p�,8���ֻE=^�27ƚ8�:B�I4\�qY E�i�$���nTR���j)�`��ۺ@�>ѐ
]b��9�K�S�<���3D����9GT�z���[@
y��@��x�qPH�'�l�	/@�Q>˓�<������=)��
���Z�<\��dV��O.O���c^�,���@n��
yD�� $� .����I(�"=9$"\0� ��2f��?8��� 꼍�c�!!D-��k�6`�P���O2lR�{�̏�y�F(mh �p2��p��*��'Z�ad	�tz@hA��s�Oz,Ia��2#&F9�U��t��2�'��]��O�$��T��`�;9\�5Gf΅aH�uKC_5�~���X���D�_�� P�N�L�!��?bD!�dףOR� �/(�ݨr��|�v=� ��Xqb�&���j�az�B�8�`��U�ҒZЕ�DaH��p=���"4e�P�- 0J%⹘%�#,�
���T�4�J�It.D��Run�$q�f�H�St�H�PG�-�	�$Z�!�
��3+&��0�S��1�E�HO�J��M�%rB䉺&(�qK�Ex'n��r��i��i�� �t X%�sZ�$���Y�L�$%9����U2d���A)D�,؀霝z�i:T-̭	�ܘ8����Ԉ@ˑ
�a|��"nڹⲮ_�]zhQ@�
�p>�I����h�R8S��?z]2ۤ��N�-�O�e8�A	Jx$>c�2��*]�<亃j&
�:� 1*1��?�	�8U
��KI[:�UÆ�� ��bF��єU���HU؟<��,S�Ā��C�?쮘�6��#N!H�1�@4�	�0�`�`"Ԗ_��������J���`���;q��x6��d�<���G��'L��?H~�Xe�D?�i@.A��C���
��d��A9�Q��T+Wsj*��+^I����%�ԍ�0<QW!@�q�7�>���;۴~fT��d@��Hϖ�����5*�P��i	���q�N�A
6�����& {�F�B�umL8��IY��	�Jaִ3��a��ȸ�ЮF���?q�!�`�( i�W!i��9QTl[?�\�p��&�z��I&'W� x�$I0Hn$��Jy2�erv	�g��3�\��Zw��!z�,YP?a����<��X�$aP�GY��c�ۣ9������C$`� @5 aL�Nј�9�����i@"�I�%#!�"����@4�O"��%������:7����5�4;<QأbS�џ��k�dR�e�@i��-�|������D�Q�@�4$b�׊N$U`x�m�����'T��E��V�'ȴ`�'SP��Yg�V�|4,O@�Itn����Լ��j�&_���~b���S��aw�Q+h�$}�ǌ=l :��*�OV9���I�f�>�3G���ۓl��y�i����d_�|zV�|bW��	��{�n-��ڏeV��@B'�Op��̼]ke�� {u��y�*��D8�6m�L��b��1a6�7�]�D7�*6gg�r�2��J0����m�)65���'ւ(�æ� .{|�J���N��U��eHF	
4���U�j	ȣo��~2�OV�'�)A��V��!(���hU���=�٢�D�-l# ��L[){�D�O��DK	;0�8���j����J?�p��i �u�K�*6��Xpr��!k�x��OT����O�����9������D
�r>�:��+R5�L ��1�+&닜S�� Q+ݴ�򤐼2Σ<�(�	i�䍁Tm��I�Ji�A������B�8U�|r�[���T�$��,g��2��Z�'w��7I��e��ɳ{_:��b%ϖ9�^P���j3� auLB2��<���%*��bs@Z\��m���^j����0(,���U��<��O��P�l�57؄@c5����p��i�\��A͏ �ό# �%�O>ǜV��$�i�5\���
�h�I�<e�उ�w��4#$�&��'�D�$\�Y� `�1	�G�qr��ϋ�r1��)�/)$�l�'F�%1��#�;"��F
٦�p=��A��&� �)��Ȉ.�a��*Nk���h�@�R�|���V�<���'�{3�L�֊Q�K�arL�k,�Ē��˭3�lP� �(^�k�^���@� L�t���U	�Ac�h��Z��]!f��=u	�3%�(�,��r�sg�It@�	iŠ0nZ�X�U�C7Sx����[�W&�O����K��&��L5^�4p1I?��)u�*C���h9J%DI�'���\E E�e��e�bB��JE"=�LůL>R1QP��)�r\�dHjAT���+3E�~A�e����D���j�%�.� ��-K�Hbfd˂��f������ʰ=�w�����
*d|��XТ�#$l9�޴3��]C��	?x��j� '��p�4^�(��@�T�|�@��Ҥ�*V�Z�D�c�]�P Q�Z�R+X�h���
?����ٺ[�@�a��-}&&R��O��&6���$@��4x2�C���G�h*��K�k��)��aǕ*�B����2���]ת��+XU����*���(X0h�qC-��(�0��M�{	a�c�F�n$`Ԍ�N^�#VE��@k��V"MH�'��gyb����D�-�HD�p�ͪ��� !G�h
��H	�m3(�$K��z8*z�k�Ns\�Z��idʓK�d�>D��ӺC�a����MyL0�1��M�J4;�(rYџ2���0,�6 �O��E��������ʆz�x2��X��M�+ W��̇#��p���<~]��8��B�^.�ڧGVd��	�K�z�"�b�~�D�iyJ?u+e��EAl���E99���F�Z�ֺIS���j����M���E�,8�C t�ɫ�~B(-?���e�p�S_����._��]p�X2e��!ӑ8D�,�6�P-w�p�̭O��ي6	9�܍�؈�{��t�#|�ڜ[UBF�*<��2c_�y��^*D�%���ޘ524$QG�;��➌�'�l�g�Zj�� �f��i��ɤb���č"u+<�h�F
/�z|���Hq�)P�ʓ���?�G1Wq�`�3��QN4d2pSo����ǉ�H��f����/+�D�!��2qqdC�ɧht��Ѕ��"񐸢p�A�t B�	�<?���l�(]V1K��$R8B�	8% �k�/�>wm<Lb���xJ6B�I�RLI�A�L�{J�W�M.2B�	;@�y�Ȗ�]�zR��^5ycB�I�:��	�-J�$猩�b�'6	�C�I�)�$yY�L�nK �xB)��| C�,Z5��g�܄c�	'�C�I4d�va��d�%ku�2錗��B�	�#A�퉓W�*�*���i
��$C�	�^;�@S7��6�ږ�! �C�	-+���3���z������18��B�	)Zؕ�'� �^֢�e�W_zC� x��4����80@�$3�RC��3�p�pd�ɿZ\@���Q0C�)� ą#�ɘb\N%�Q�]$�TZ%"O�ؚ%��1|<|��.։	��Ź�"ORZ4F��ZO��p nWk>TJ�"O��r���
��P���_�αQ�"Od����"T����p��>?�	ba"OZQ�l�#hG.ٸA�� �t���"O�PW/�&w� �O�P0����"O�Q�$���3BP�3$>=��"O���r"Ɋ�~� �@�u.�Y@5"O�t)3��8dŊA
�*H|��4"O���vCYRX�����l(���Q�<!�c�O�$��VI��yKd�C.*T����#,��8� l�"<�,�Fm%D�TP�AC*v�$r����#th(D���rk��mҴ���BŰf�1[qO3D�<�� ԾNP�KW����ő�0D������.��!O��R��e�*D�p����b�N0�Fē:#��H��)D���p#WP����$�տ���!�&D��2�̺~^��g�(tص�#D�\�p�Jٶ�a!��	H0=�c�!D�lpPB!O��2�P7��#�%D�a�E�>�
��!nN�n����$D��C�&�dB@�A�M�t�ܱѡ#D�\�S�L�|T*� B M�H䪕��`5D�̺p�D+8$���՝_<h�µ�-D���M&�:����2q�FŁ�(D��CEF�d���'��X��@*#D�R�I�*�u;sMۂdΕ�d/!D��z�"ɛl�|]���<_�1p�=D���J
�@d�p7
��S5�59��8D�xi��]s~s�A�Pbj�I7D�t��L��J���BR�'�a��4D� ��͛B|~��M�	�����6D��q�/H��k�W:&l��o2D�d�O��Av�۷�#7�r�H2D���k\�A圼��L�'�l�)0D��RF��;~�D� Æ�.����/D���dꐽSJR	���1l����.,D�h�g�>m�� "��v�xl��
)D��;d��!H�k�L�^�1�&�)D�ks�))�v��'!\p"��s��&D���QE]	_e�hb�G�9;�ز��#D�$
%�z�*�3
ˌu2��i�)$D���C�9�҅���G~���i.D�\��E
,{l颒GG����3!-D����@��=!�	R�JX���8D��0��(�LtڗJF5H� A�$D������PΙ��	�#�V�8m=D�|n�Y22<��H0r��r��u�<S��q�uX����ZY�#��u�<!A%> �M�q#�V��Lh'��o�<��k�=*w�]*B��!;�u���i�<����;ـ�I��ěm�� ra�c�<Q�'�h����kZ�kB���ajt�<)��/p����(u:ph���I�<�s�T�BQj̪ŇD�\#�('UC�<���B�p��lӡQO8�A�Ve�<A�����M)�Q�7@r0'#La�<�g��� H����!I>���nLu�<��Bܕ<?,�Z������B�&z�<���6A���9��g{̄���_y�<!b)˅DE��Phǅ3<B  w�<�hԨ@"���D�y�O�o�<� �8vb�o�^�����l�>؆"OR�B��V�W�f�x� �"S���['"O2�3�߬ƺٱEo�tC���$"O�tpǄ�9� ��f�,
�"O��b��7�0@H�)��WƦ��"OH��ri�e8��%6��M1""O.�*��@��t3�&F�3�B�pw"Ob)��a
���������C"OXd�g�ԉ��X[��V&H���Y�"Oz�ʳ���=��Q�ѐJ=
0�"Oj�J�ĺQ�X8��(26@-{!"OK_�!3إs�+�<P���c���y2�]�|)$�񬚤[~��G�O��yR��vN�yT(�!{6��F�)�y�l��2�Jt�	�wcn
1	�y�薝&�Q����8<���נO��yr/܋J�M#��R�ͣ��y�o0B�&���#̱
 
l��A���y"�#�""L@�6�IDlS��y��ʙ"�����v�քpD'��y�#�D:e�����g.V��@a
��yb��lb��ŉ� w�>ac�Q��y�eZ;3�8lY��2mPHIPd�y����eM��ѤeS�jߠ�qp���yR�@�iC^��6��;]�����yZi����C�V�QrѸ��F7zB�	�6%�Y���^; ^��b%eقC�.+�⩀%L�<'��[ ��5�|C�	��	�F=&ޞ�񄋴{�B䉡^�8��pD�8��p�.�(.�C��bt�`CB������2gB�I>D/�%�FX�C��L!�B��B�	 e����%� 3��4��D D��B�$Nʨ���
2�|�&�]�4��B䉛W~]��g��t��Ƀ��9
|�B䉻3,�B��T(-�~�Ũ�7ܮB�I�>�1���"]8)���A`ϜB��7x���S�1p��x�5n�\�vB��
U���Ύ,�t���\!`B�wzDdZ#��.:����\^ZB�	#q�Vt�����1b\+���5�pB�	�A���Ǭ��:�*�R
�8��B䉯C���h��6$V���̝�1�B��,h?��igm<�h1���y��B�	�]�P�6
�n�T	j���if�B��F�z`���&%�tpB�Q�6>TB�IJ'4�IEb�1?� 	�7lJ�@�TC�	!l,UR���>LA�4f
�`E:C�	�f�6�@����V Ѝ�"EU�A�$C�I&B�4=qԈE�fܢY���*Wg�B�	�a�97g��|}6�ӧd��B��*>
���G�Ȇ;o�u�p.�O|�B䉙	]:Hh�'§D-:,��*��w��B�=H6����
U��qs�Q�t��B䉅z|~�ywe�=|V�E����cݔB�I�kY��dT*XT�Q����$a0C䉧2⡘cTAN m°�C/p$C��;	`�)�����(�j��z:C䉫v�^Y���N#0)"�X�	_�8�.C�ɩM��A��cA�$ڠ'��$m�B�	�Y�24�����I
�G��s�C�ɿ_�x�����]���.w�HC�	�$�2c >|�,��ag<C�	 d ~���ɗ.�x�0E�@C�)� `%2d��VҲ8��_���rr"O�5
V���8xS"aY�!�"\#"OL����d�����*-��)h�2O(�=E�d �=��q����4�)TBZ��y��Q��`ˠ����&dZS�R��ySr��
� 	Z.�i1�O��yR&���a�Lep8rΔ�y��߹]���Ǣ�f(�ύ?�yR���V���Qr��v� �##�yB	_�!
��[s��e2@�A"R:�y�` �j��Pt��3�x�E���yri�t����b
Xz�*@���y��@4;&�{Bc�L�(;�O8�y�,B.�B,��m�;���A����yҡJ�iulq��!�T+8�3Fkض�y�a��i���3f��h����K��y�@L�S���!R!	�� �f�ɬ�y��@�*@	�b[�N�>���'H%�y����gtբ`Ǆ�ɬH��-_��yR��<��d�� 5�d@���yb�
 !��gSt��TP�y�.Av=�)Y��6�^�A�U�y�^(]d��G�F7�%y�,�4�yr-U@�I�	ÍK`����ܖ�yr�,4q�V芢�I��C��yB������范����2�y��B�>��]IQg��|��q�
�y�_� ��4Are+m9@!+�� �y�'�M30붠�c�8�p0�Y��y�D֏un�8���4X�B(���ƕ�y�X�<�"����^�M8����F��y���48�%�@dɔC�0t;"͌�y��Q�;�j��D�4g�����8�yb.��S���
��ӯd�ι�q���y��
�g��Cp͝�`�Q� ���y�NUY �:F�,���QЎ̟�yR*F�76Z���Ǹ3�ޅဝ��yb@�7��|��/>D�����y"`بo�q{�a�M��2�^�y"E"���]2G%�1��j���y2�R�J�\�af��:�b����;�y���-b8��PDп'��<�D���y����UʑSn�.J��\A�ț�y�fڻ]��Q1�)�AX�
g,Ɗ�yr/ۧ��`r��9>܊]�%�?�yr@�4]ޤA�H�=~��� ���y2�\�0�%D��e��j�ו�yBC��`:��0�ϒ8iE�	3m��y��4Q>(�G��k#\�!b�O��yr��[��Z��� W5f�����y2D�v?\٪��Y#�ʓ�×�y���~�h���d��W���`�LC�yRF��I�e �п�����Ӌ�yBEQg�p�i"d�,@:���¤�$�y�*֬~�6u �A�8.w�j��y�mԱ<�!��Y�".b�Yǡ�y��E!]�=�P��=�z�Z��B��y�KԅJX yYE��?Jox%#�ӣ�yҤ\i� �H�l�*qL����yRj�)�(5��c��m8��"E����yRY6Po����g, <�F���y!_�Z��]�j�X�d@R�ʎ��yBG��_� `��(׫X�.88 ��y�CܚV�δ!�톹OQ�4T���y
� ^�8�ˎ1+X\U���V�.��"O�%�䪝9,��i <� ���"O�h�T��s����5��*K��"Oh���9p'�УC��.I��Z#"O"���Ӣ|$�KAK*{�n���"O�=���ɺ&Z���s�ԙՠ�+�"O���D��hƚp@v�P�Y����"O^u��R-%���b�I;n�4U�V"Ou��f��8���H�h�(�ڌI�"O�	���b&�XI%&�J�z��"O0HУ�5i6��#�az�99�"O�� O�������ܜHur ��"O�8���.tt|�uIh�Lja"O,��h�;_�hoM�]S�,�7"OV�ʀ�:h�TxPdG��1S�[Q"O L;��X ���'S�4��a�"O�9뇌�<l(��	�;u�1��"O���e�W�8�0�� ^�!"O`!�D�B	=���1Ǧ�씜z�"O\D�w/N&��$���V���"OāY���6�΀���|��ݠ�"O�c7kЛ��)����:�T��f"O0�B'�4p"�u��S�5��9�7"O��AmX2�h١%�9bF0U�"Oʝ�c�`�&���&O0��#a"Obe���+4�:�k&�Z*\q��"Oȕx�-҅#�⢄X 2�ݣa"O�a�q��J2zА&�
��ؓ"O�|Ӂ��<M��j��^r�n8:w"O^���R4�$�������[A"O$�i%雁4j 	�0�<i�(�)�"O��[���'4; }P��S:�+E"O�Ka2�d3��I�&��:�"OƬ��D�Z'���)�S�05��"O�����Ѳ_о`H�i�&*�"��1"OJ)�@U�`{n1��,BwĄ��"O8��"Ҫ(84m;� ��]L�1�"O$�c�D]��) �Y�䕙"Oz\���;6�d2p�ȝ1���P"O��WEJ�V��@���6��e�"O�Ũ���2K��@�F��� X�"O��Æ�5���#��N�	��"O���%E6uB�mQ�e]$F�]k�"O��V*Ui)z�d&]QP��{�"O����!������,@���"Ol����NWΑ� �;q_�M c"O:���?T�0Rc�ǈ����0"O8�CT�\4L�-S���E��܂f"O��	����z�͟�j����"O���[�o�A�uK�y26=#�"O���@x�p�ѶiA�a�>]��"ON,�c�%F	$5�g�;�h`b"O�XdR
}T���b��!�x�*"Ot��J]�`t�s�\#=�z	�"OdeKc��"ʰ)��/�*ԑ"O��	��sP�8e�Ŝװ��"O��cMXS�l%Q��'K��+�"O��z�4v�-b7���/Ӫ	A�"OxSe��Ô�� @! U�=��"O�E�M��}�C.�ZMh�X�"O&��''�KI���R�G1�%�@"O�y�c�`�<�B�]$-���c"O8�04���>��PH�k���
�"Oȴ@��Y�P���#�)X�x��A"O� |��A��m�|���B��;~�8��"O
�Cbh��|��sBE�x�n]��"O�Ѐ���A���萣��;{tՓ"O�P2r'�6��Y��bҳM�|��E"O�+�A6��8R�a�W����"O�-z�I�0�8\!f���O7���u"O�y��[�a$-��)ܵEA6�*�"O��"1��B�p͐�_1V;J���"O�*��+t�`@C�th\
�"O��#$��4��L`���ǺUhR"O�Y��	D�c��UX&�O�nA
1"OFH�tMٞ �|�HV��/��l��"O�IS�C�E�,�ڱ��&=�vU�v"O #Ẃ�,�.��jƆy���1"O �Ȃg;����w��(��+v"O�H3�CA�@�Pb���2�x��"O���`N>
� ՛6��rʨEj�"O��$ș$�P|���ǚ�X��"OBP�����K�3��x3�"O,�sCɗx��B�I��W��A2"O���DsY^�(q��t��"O�`��֩e�b��q��	r�&�B"O����.�|�F��F,H?Gֺ%�"Oz�`�[�8���pA���)�艨�"O�]s�Q�Z�`E��m�4����"O(���l�@���J}ɤ"O�آ�BLi��"d+߀n���`W"O�UɅ�Æ00�A�g��TS�Y��"O~ ������b�i�G�4
��m�t"O����#Ã��9 � ��?��xQ�"O�iÁ�Όq�H��p��^|�U�5"O%P��x�n( g��9bB0Q��"O�d�NA	Y���׈V|Z��c"OR�dE��g%�}��'=*�x{�"O�(�3G�K��5EfyH��0"O~�� C\�;�e�o����"O>q�fʎ��N�o��\`��"O$��-1>B(��
UvJ��w"O�VL�23�@�qhQ(Q_�p�#"OD�	!�;_0� !s&��\ln�*r"O��9�.�/r���3Wf+rc�d�4"Op�jr�\�zV���lT�"o��y"	(lf��Z��U�:"p��EK-�y⎎1+��8ÂD�"��U�R���y�O�D�Q;dn�=�aw��ybÑ�g��B0���<2&Í=�y2�U�pT�[2GZ<z.�@E�߬�y����D'r�y��τl|�B"�y�B�>q�`C"B�^�	ТȞ��y�OԈ[��$CĬ
M ���c[�R��	h��Ui����ϒ1�|���Z�y�4�@����!��	5�ܝ� �Y!q���iĂқЛf
O�0�'@°d�tzë�� ���"O@���ϱ$Q�PV<w�h��"Oƴ롦bx�qjw-�)��9�"O��*קJ��Z1,%��=	w"O�4���IK4�&K� �`�"Oؑ��ƷLTVp�wI��p�,��u"O�mⅠ�=La849t	N�/�k�"O)uJ !��0J��	8��d���'�I6�jt��;h�<���ŘW�B�	�[6�Hړ~� �����B�Ɂ(x��7'[���H���_]�LB��=NO�uBU�\��y�CH�Rt"?���� FyK=��p��������V"OD�` @@�V�XZC �J�bi9�"OV������
�� B�̭(�<��"OB������^8r���N]�i{J�ɳ"O݃Bc�;@P�@�� J䤚 "O"02�Ү*����wh&1a�"O�L9@i�Q6\Z@&��n�B�"Ov�gNGL��4��_�\l�P+GO:����W�NQ(���.O8��p�w�Pf�<i���*:�c�L=zk�ܑ#@x�<���*Z�Lʕ��8�9�COv�<E*V�-Yv&��A���1�u�<�'�V�/8�fȂm�@E�TJ�|�<tC+5���ؔBK�2	X��$� T�<�@��3�Ir�CSBx���	[k�<)A�ΆtqaL�>p��4#�D\i�<Y���7X~����:LN����y�<qr��,8��Ĳ@�n݊�Vu�<����l�� {Ǝ[/8="(Z�,�e�<`b�f�� ф�Z,{��aS�i�<q�ا$�`t{QLZ�szZ@����b�	\��h��I��m��<*Jm	�%ڴ�6�T��DH<Ag�����ĩ��Xw����eoIu�$9���O����G#Z#����'��-P�@�'��L#��/f�D�b`��먘A	�'�,�[PaPUQ�=0AALY�8Z�'�	:mԭ�~�����I�2��O���� )����f� i
�Kp�\.hK2���>!.O���IU�	X|aH��M׊ �f"OD��!�c9��Caݛ1�z�#"OzM� k�/:XY�c^"�xY�G"O�p�A])M:��dI�u5"�[�"O �	#l��.�4�;��U(P伫v"O�ųŀ�dׄ��&hFSh��f"Ofes�'2P� ���a<�ʓ�'|��yH��zhs�(Q4-��ڐ�7�y�Ƙ��&���σ� r���2�[�7���<Y���~b#�&cg6��.W�l�sw&]�<Q3��8"lۓΔ�?��S���Y�<�d� &�Z-Ri�1Y� �WY�<�����ob\���F_��m:5*�Ѧ�E�'Xz���l^�T�6���FZ�@����'&��8�d,;���q5#��b^ΰ"�'����
n+�	���R"]����*O4�i@.�!1�*�yw-_�W�h�"OJ;��� �	�ƞ�w��Xk"OT�@���"���Iy�@��"O�E֧��W��{U���h@����"O��Qĭ�q�"aa�#=>.(0t"O�)+'�]R�I� *h(,�Б"O8ܨ�g�2����嗦<'�@�"OT��R�ԗ� X��M2�!�!"Op�Uh�
�:�B�L��Cθ��"O(uP�OÎFP���Y�@k~)K"O�hY��;-j��ds3�MA7"O2�``��+m#ع���)xm��"O\��!��=�����c�|%�R�"O�sG�Z�(�[H�B*]��d��"O����D#k�(��F!M)�� "O8�9w�����ЍϨx�bA�"O0a�Y8/�����ǰ_5��"O�X�(12!�S@(�x��"Oȑ`�ɟ2$^�2f T�-D8�A#"O��!�'��)g៷27`�:�"O� ��WN�0#�!���M�A2E�@"O�t���7<� b��=|AМ�f"O^A*��U�~���K]6�Q#u"O֨�"��]������Y5�I`�"Oph��ػ�`��X;$1I"O�Uk������Q�AL�&"PEH�"O�E�		5@p�&��#�.H��"O�d�@�ɐ*����C$فdd��s"O�r��$
J	X��I�GW���"O �,է3@�A��@БZ8~�r"OLT���D73��M���_(�8c7"Ol�	܍:@�j2���[:���"O�!�Ԕ)��EX���<3^u�"Od!����fN�ѣ���a[d+a"O��4��0Iv�򗭌�.�~ps�"O��qW˙>j�Ȉؓ͟�����"O�]��+E� �3��9]�p��"O�x�/o5���ǥ��	J�%"Op%�p���!��Du����"OJ ��b�O����C[�Ip2�b�"Op����-ٺhz�B~��"O�y!DlP�{q�)9- 2Np�(#r"OHMZa��	-Dj��&��Mp�"O�#O�
�x��#�b�ˑ"ON��C`��~ ���*:�<�[`"O��K5�,�4��3�/\�IѲ"O~�� gJ�*W85��&�4@�=�E"O�����.����@�� 5��y�"O~�{��Dv^LȀ��z�}y�"O�pp	^6f#��!�$�v0�٦"O�1�'��
g��m���o���0�"O�˖lU�X��$�F�C0C�����"O�8YG�BW��Q1i
'^�n��"O:Xh�D� g��"Í���a"OJASfȀ�y�r�������Ő�"OА��)�%�i"G��]�pEP�"O4(s�g-,]��h�蚆3�H�0"O�� �!?�}�7Aəc��ػ7"O����@�z ��桟so^X�t"O6)J�J�3D<��"��߈�輙�"O�tېb�u���sTO��%�Z	K�"O�����օWBt��u W+=�d���"O��r�T9Q;e�To%q.	2"O��D�]5��c?5T��"O�D`�e�47$  ���hN��!�"O��[Ǝ�,[����KY	Ur�CQ"O�t`�b8��a�'��V���B"Oh�	d"R�~aEHL(X��`*"O�mK�R�Al��Bhف���Z3"OX��1iV�/�J$Ȍ:x��F"O���.C4F �UJ �Mc�b���"Ob�xw�E�#�� 3��"��ɢ"O6$*p��3F�^���>*<��آ"O�4`0��~��:Ή)31��z�"OvX2q���b<��(�T�`��]9�"O�h��$�>�F��cςA^��v"O��GR��~M�w��K`ʅ"OH���fZ�g�vH0S��1v"T]�"O�h�N�g�N-�WMF+�L�0�"O�a� ������+Z��l�:"O^�	k�R6 1t)َW올�r"O�!{'���&�1L[Ԗ��`"O:{�i��^L�̢��y��� "O��0k*r��DBԆ���<y�"O� ���"�!�̩��{��\��"O�	+�f��9���Cp����e�"O��(怔�5}ʱ�׃�5�$99Q"O�)+�a��er��0�܈��"O�Y�g�@Cg\Q��q+  a�"O|I���Ϗ;����-v���"O ���b��S	v%	��$&ft��"O�-�f��(]���"7���B(0k4"O�D���;�~���	�$]AA"O�a5�I0P��yÐ�ߩ�v2�"O�t�A$�~�Y��Ƙg�"�%"O���D-\��ѤڕD�n�P�"O^�[��L@8����:'�r@ig"O��%�� �|\)˒=섍� "O��T�rV��`�
g�",�4"O m�5D�W��H�	У(x�"O�鑔���6)EI�+h�T���"Or�H�ݰ<�lk��ފ��u"O��kq��L��9h�JEI���#�"O��9�J.�>ܲ��\�C��+ "O8���٘uX�(I>O�*ls�"O�\�6'pLء�T[���;�"OpIh�FB�9�6��E�c���"O���A�)��
Q3i�r���"O|}�sc*M Ыc`�* �"O=�R�͙5�����O )G/�=��"ON�`��<a��s��'g"x�bD"OV���*���L�Fˆ�����"O�1��Ć0L@�`"��5j�JQ��"OޭX�lA��D<�1J��f�聓"O��k𭟋y�����BB2F�"O� ��-`׬+F��),}�"OB� �/W�\lYB�ɓ�T�8Ґ"O�d�rm͔9�d$���G:��ј�"O����� �T"�o�>��e"OƝ;@��3M;�`'`
�5ɠ�ˤ"O�TU�$a&�Z�OS�2��K2"OJ����8u�d�PO�%��$B"Oȼ"GMױi�jL`�.Y;}@L��"O
YJ7M�8f�}��CO�mvً�"O p`�PBX5�߹Z.	��"O e��L��^G!����S�M��"O�Y� �T<*t�
�Cٙ
�\)��"O�8lC":�^���#Q�.a�"O��c6��&���Y@�ʳ"Op��GDR�v�8���wڨ\�u"OX9HAG�/����P�OXb ,��"O.(#cIN9-Ra���UP6�
""OXxq#@�o,��2�4����"O�}�A+I`���ъJ ��@�"Oh���]�U�L�#��́$"On�vK�L�4����#�.=�C"O�4�"��==��)S�;���"OdY�@� +��W��P0����*OD��!��d��]�1l�<=���@�'<���˔-pڀ@H93�,tk
�'�%� �F�����oI9�TI
�'�n��1��n=Ibm@5.�2�"	�'���@�RnpQ��`]&�$��	�'���b�D����y2,׎ɶ81
�' @�Àו&{<�Zu�ZXA��'�
��u(W"�1�Ǒ�@�x��'�Ɛ#�4F�q��).u�f���']| �td�`ib�bA�s�]r��� �]I3f>((��j�Q�IQ�"Od�bW��G��$�H�{�N Z�"O��3#L$x̠��T'4T܂P��"O�A��-�<Xv,���^)-�\Y��"O�I:��S�`���ǗX��T�"O�A��G
\�PY�Aeޠdg�y�"O�3�OK�>
Ujv��I����r"O�)�
ݟa��ʮI���"O8̙�M�%N~ֽ@�ꈃ\sz��5"O���"H�%�Bi��)�=����"O��YU-_������	L����"OΘ
G�E&S��Q���9�B��"O��	G/J�Y����WГ�z�h#"O��9PJG4X���7N|j��q"O�c��˄/}˄-	�W���Ȥ"Oz�3�$��9M���K�x��I�2"O $�!�5m�*@��*�9�� ��"O��rE��|�k�	�)c�Y�c"O�I���łl&xl{F�#X|q�"O��[��zΒ�k2&�7�p,�C"OL	xS��I�޸�����]��"O��i��p\(�2B��>Ӵpb"Ozh��D�L7j����G�y�"Ol<��N�3��0v���=1Va��"O�)�N�)nhX�$4��"O�#�M��X��\�,ޕW�mv"O��!�A�?ȑ2�+R9rЬ2�"O(�8W�ƲHv� u吳"U<$�1"O`+�H�$J4r�A�U�]0�"O��:���{��=���Y�T?�@xF"Ol<��^+�-�w�Ɗ;+(Ղv"OdEc�F92uRM�5�#"�Aqr"OLԈ#@Cd�
�k��:�h���"O�,!��giTe�" �
pڔ� "O DZ�`Ũ4Z��/�&L��9�t"O����A����j�"��q"O�9�t�À~�,���f dE�-��"O�]��B�NH���3*]�\x�d"OvԂ���7�x�#ڍr�nQ�T"O��1� C�9�����@!E"O���e�;H/�e[ǝ��y;�"O�9�[�JH��KǾ1A*A�B"O`Y����R<f}!�J ��� ��"O�)H�4k@���s�0��逥"Op��ր
�L�!c`h�!k�ZQ�"O�Uc��cwzّf�r���"O���MR2vJ����>�p��"On��`H7Q�h�ȗ
�<j��"OZ8yE⇘j�T���_=����A"O�5��=\4���S46�>E��"O��jd��A���R=%��ܸ�"OX��0J
;:����y�$Q0�"Oa�W)N�rؾ��%�|�4���"O�����I�d�q��.�~�(�"O�M�ⅆ3Bs�@0���7��ih"O�,�d ZX��L�*v7��#"O�Pʇ�e�IW�S�a��3"O�Dc��Q9y0���hީ	�~|Z�"O=X������e�$P�҈B�"OvA���Ǟ-�^�0˾9*ra�"Ob5J��S�@�T��ȞF��q�s"OR�q+�t.��x�0&�(�q�"O��%*X
"Hn'&��<�Zm"�"OH��S��6:�9�7نl\��"O� �#�i���"d�4G�y�P"O�����'W���r�\�>�d0�"O��5��5�Z�5#��$�"O����,%��`��ώ� 0Ar"Ot@�X�b�T������^���"O��r7#�6f�|/�*,d\�("O����
+.V�BK��-b�y4"O~,l[�"0�SG �=&U�|C�"O�I�#Hʁ��� �dޑ4hbUB�"O"ѣ��'����Ǭ�.|Gj`x"OV Hk�. � ��؛9�6���"OFh
U�9Ip$��φ�'�ƜbQ"Ov���Y<(L�kѩ���,��"O��a�l������F��58�>�H!"O	�%�������W=t���e"O���-  f����������e
�"O�9���_%;��4��(��x��U	�"O�\�&ŖCZ�-)B�<~��(q"O������\�EV8���Q�"O�a���$h���D�!��	��"O�-����".�4���%�lw��#�"OV�#%��[�2ب2%g`�BF"Oh��A���R�>d
�iR3t��h��"O��E�6[�4���+ߚ��"O���v��.B'd̂R�H�X�k�"OV�Q�ZT�spo�=|b(�1"OءBʆ-I�^�pI��<)��p"OLT��*�D����)�#��,��"O:TyÊF6T��ṓb\+1̂���"O��ؖ�� p���.Y��͐@��y���5��`&�F)��I�蛬�y�`ˢ>^�T#��{\�郒���y�&�4VLࠪ�tb�)�1�y�nӿ7�b���EԟsZ��!�2�y�B	�,���I/�"j��yp�y�o�)e�.@��MP�v��P��ҿ�y�J
�o�>�!��k�R�Q ��yB�50o�Dj'�Z#]�8H�w��7�y�+Qo�䈵�O�䤀���y���-.\���XX��E#Y�y�ݶnt����R�SdX�2�h[:�yB�ƴ]dx��+� �ƄQ�F)�y`E�+��$��@� ,��e`ۧ�y�O^01Le������4�2L$�y~U���m��aF���=+�C�	�rՠ���42ܙ�k�+��C䉾�.X��MĖdDS �4TC�I�6�d)`�?8�4��_C�	�x$��s��Z\X�s�X4MO4C䉶����g O�:W��fؾ7�8B�I*�^<�Â)"W�EY�NX!1#2B�I#R�x�'l��H���B���0h��C�I�y#��KլG��V��%�C�I������ؾ
#rU��alU�C�?.i�M���_I���x�D
�8I�C�	&��Y�]1cV�EC�J:L>�C�"|2�Z��*{�i�tM
0~hC�I�h�
�k ��&z�n���F We*C�u٤��A�g*�8s�F�hdB�	�IBb������X�D�D2�B�I��ؑ�fѫ'���a
B��;��j���[�ր	 G5q�B�I0'?�ܪ��
d�p<@iW3/�C��a<vp�&�tyV0�M�mThC�)� P$¦��G$�(a��g���1"OX%�`�QR�FEa�N�nJ��"O�)�o��W�w��n5�,�"OD��j�Lϔa���Y�` բ�"O���B̓� �۲`�?@���%"O�e"��=ZN<s�J�5I���2�"O
D���O>tq �
hS�����"OԔH��6���)e�!KU-G��yh��o^��0d���`%i$�W�<����\�B�H�&ʊ$B�MKE�<61rjl �k߾�ƅ����<��WK�51S�[)N�x[D�t�<��,ZsNi[���u� ���v�<��IO��z7�
r_�+�Xi�<��HA�'=b)��c�+1���@5go�<�	|��=jE�'a���#Gi�<��m�c�NĠ� C�����V�q�<	�ƚ\�&��1����p��^k�<�� x��0�ש���޵�PJ�o�<�@�.�SgT*	����ā�E�<t��!l򢜚V�Y�v=* ��y�<�ơE�'[�(Y�
 M3 `��Ut�<95�E�:�aE�NP6���)
j�<�dG�V?V�r'Ye��86�l�<9S��'Ob^!�##0g1X��ALM�<q�U8Z���h��өaH���*MG�<����m ��J�z p@#���x�<WM�_�JuK境������H\�<qgƈ/�"ڢ"=�| �I��t�B䉦g:^���I�{��Y��*�?m�VC�	�Ix���s��O�=I�A C�		  ӓKM�C���#��Ӕ^$�C�	�-j����@?0�S��O���C�ɡG�8�S��9tdR�ٴ��%�nC䉵V�Y�� B]��q���$!VC�I7~e���%��3���	���C�	9Y����0eǏYz�p��"بB�	�	~4<j��N�?HXZa��/�B��	t�BPS�,ڠ��9�a�3XfB�ɄZ��հ�.�?��MqT�I7$I(B�ɄpR4�`k@�A�n�dLZ*2��B�I�n��%�!��xMJɀ����ZB�Ʌ;�P�I�]*�]���(�8B�	�P���H�8$�H9𶫋,]�\B�3r���,0�@E���ERB䉄��Pp�:]��� �U�<
:B�96&؍�'N݋h�"��P
<�nB�I?-AA3����>\#A��H8FB䉨'���A�d����p��HYB�A�xl����0[�\ X����i��B�ɻJ��f�	s�X�iBLqt�B�ɻMtʬR�
@�E�\��ǩ�S�zB�,5��@ɀ�
n�ެbE��K�B�I3���!�%b�����O���C�ɤN��I�+))db�#�5m�:C�I�Q�h��+�5PZ���
ʱG�2C�	.tW�y�7�Ӛ7�(��2DF$�C��5vn�
��W�C� �h��Q�|��B�	3�-A�J~2HEK��+�B�I2j6��%�)T��A�H�\�B�Ŷ)�R��Һm�����B�	�q0�k�$̎j�^� �n��7��B�I/Yi�|�a�"�j �$��k�DC�I�EF`�ᱯ�PW
��s`� �8C�)� ��.Ă�A�'@a��] 0"O�I�d툷�"����ߗ�
�R�"O����0��ɀ���	~���"O��b]�*G��@���<V�d1�"O0��S���X"҉���:����""O�x�Ae0<��a���Ɲ(�H�"O�	v�ԯi�81�C�1��rD"Oa��H1}�C1�D�v�j�g"OT���'B!Nʠ ���<�"O���"�c\�AD�K�-���#"O�m9uF<]l�oG���v"O>Ò�رA<MSg�ƍ+���y�F�*X��5���S�����5�y"��y�P�s���4O�Nx6��y��6&�ީa��X%{~�2pŞ�y �4ʨ�P��rZ�x��$��y�"S'v�(\��@�7q��K��6�y�� 9�A���l��� fZ��y��-�&�a� :X7�Đ �[��yBjT�C�:�MD>>tx�[ �B3�y�#c�3�Q�6AeӢA�	�%��'>
��3�<���(߬ ��Y0�'�<Xq2-�=�ưz� �&��d��',�ȱd%ߑ `Y"�(��]Tt�
�'=������������=W&@�	�'��O3 X�t� l��?^ Y�'\�P/�>��� ,B7�p�	�'���z1�_�l�:5�P�Α.�U	�';��I3I�]�9B )	��
�' �@B�U�1��*`�1gvx4��'�Z�ä�ϧ!= a�Q�v��'�^�Q4��;p0���J[C�n��'	a�D�Vv���%D�#�J���'r@|頦>~,�D��c@Yx�'�
h#��
��:�fO� �
�8�'�F	Uj��.����>
dp��'o8�Z�ҝ �*�f�����	�'�Nq�f��'T �	ܨ}��	�'!}Z�c���xi�n�ufR�	�'k��F�"p5,�Q�Q�q]4͚�'�0i���.)�)P��6i%~�H�'|j�ksF����DN2��ܲ	�'�n���D�5�v���I��,��'���ȍ�O�t*Ө�?x+��s�'���������W�o5L=��'~p<f������B�21�a�'�|Iz��(�"t��݂:�H)�	�'�h<�r�#���ef��F��y	�'��\�g�Y�m$}@6�
<<`S	�' ���b��@BU�"���jr~�A	�'L��c��=�&�\a����'���)�!ư��X�&�X�Eo����'+6Ab�	�'�QQ�. 7�Ƽ#�'��$ce�;� ܋�����	�'��&�Fvm�eÑ�CZz��	�'�`E���#)}`�xaF�9�n�!�'\��w��6�t�pKV�X�'����'d˩)��������LI��'���)Qʍ6h):����^,'n(��'A��y��ըF��r�N�*���'2��	���- ��ڰ�ʤ��<��'<vq� ���^��uB`�H2x�����'�� �PC�4N$X�9���oL�!�'�'c��&�nL�� S�$A���� $�`2L�]' 5z��Ҙr���p�"O�]qfث&�rm��%<����"O���e׸bX�����3��� �"O��#��9pT�u3c�5o�0��"O½b�ѹ�@�
"�6e��M��"O"�e�ʡ{��;�
W"gX,�q�"O|����T���<��	���R"O
(p�(8D]��Q��v�|�m<D���F��	���4z�J5���4D���"8�x�
����<� ��?D�����+5��V��7}��}�fL?D���%O����O��Y<D���f�8��C6$�ڮ�8'K:D����FH:M�PT�&g�|\d!��F8D��0V'�p� I�'�\�h�v00��7D�l r�ؒt���y�AY9l�T(�)D�9҇X�]L
�i���Ǩ2D�\�v���(?�3�@6̼�Z�0D�`�AFW�:��+�IU��I0�,D�`7c\dE;"�L4�:�FO,D��k�٪r�2��V���*D�̰0��$G��kU��
�
B	)D���Pn�
�L�W0-���Y�!��l|nLr��߶E\���e?i1!�dK�yzn�`6˅e=Hhs�
�s!�$�f��D�@��<�Y�DU�G!�-`��d	<}@qr�2!��<"��Zc˖� ��Cf�7Be!���0��(�KH�+��f���fG�ON�S�g�R�2�d�ޡ3J��B֨|����T3�Y ̊�1�>!DM��1�ȓ�:�ZV�r46@H�	���ȓ|���{#&�f��;����	�ȓ4`���W�Ӌ?^�ЇВcnX��ql��#O�y�n�3Iѐz5rl�ȓ*��1ؤ�F�{3��kT�"iM1+O����O����|�rK8����>])��{ B��Ra����^�(s �A�W��R�����m���I)��5ohva\e=^d��#�X�b��Tk;*h�0I�s��1��A�hp���C9]�8U�'OͥLiz��z�~�� �[�L:B��v�ڗqy�	��|��d�k\�+�ꏟJ�"� .O��D�O^��I�|Γ-���Q�`�;\x��cT�H1���ȓeL����C��f�[v�˃f�e��LҔXk���:�u+��P�o��t��u3(a���'̰)l"-�2���}KW���r�l˓�ל��x�ȓ�h�HI*��ڧiEn`�=�ȓv��j�ƞ1+|�jCFܕp=YH>�*O1�1O���F��� �"�ZX��S�"Ot,׫[b M�胔2�uɐ"O@�H�Dh�YRA��I�¹;�"Ox���^�C��ڴ���4��Qp"OF��ѮOo��ႂ��"�~��"O�A�#\�%��Vmԡl���jr"OJ��V>..�i��>���ِ"OT�@��Ze��r �S:����"O���aD�I�z��� $	��X`"O�dq�T'p���mѓ}�q)�"O�Tk��L�zv"�JP-�3<ڰ�{"O�M�� ]��T����H]j�"O�!X���.E��� �K�PS�l�*O\����Ze,��鉀y�z���� ~u�Q�,�R8c���Y��u�s"O����(	�����16�^�Y�"O���+���v����:d��h�Q"O�Ɂ��Q1o�RQ�P�T�i�j�6"O��#�eL�(��Џȼ4,�T��"O �(`���r�(�ߜs�*�9�"O�M���	��x���ǵu����"O��yU���:���B�N�p�f��"O��2� ��9�LH��G�n��"OB	X4�n�r���=;.�̛��&D���1�&bD ��5��$X��E��1D�@��p�,xa�%
�v:����-D�L��ԟ?kf�+]�K�^�	S1D��h�*ڈ]N�b�Y> ~�Ő��;D��U�Ň6���
��
|�y0!?D�8S��)Oh�Sӏ*�r��/D�����(�|��4����H/D�H��`z����+{��Ly�g+D�$��E��	�$���T-I�xs4i'D���$m[0)�X����%L�z@Sa9D������+K����BQ�M�F@)U',D����ًk��*�&�,���*D�X���'S !v
\?��yHV�)D�$XgJ�G�`��j'j}�1�'D�����$2�`�e��n��0�� D�D��HK8�8�9C���]��ƀ<D�D�%��"�������I�"� �9D��񇯂19߄����ϡTY�dq��7D��P�&�4�Eɀ�f��У4D��Rw�j� 3NS�Ұ�b�.D���"邱GƬ YEN"[8��� �+D�`Ť��TxP���F�]*���$D���	Q��`s��3c"]���!D��7"U$M&�@ �]�=|�x�F"D�x����z ���h�n �Y�h,D����BL"/6h2N�':��.7D��(���*U�<��7b��*D#1�:D��:d�R,a�h���A� Zd+��-D��k�Z�T��H�S g��]��,D��Z�΃0=d��壓�Tc�i�B�?D���ւ�-_6I�s�O;e����+>D��Gi\	%pԑ�`�Y��q��F)D����ū|�^�{���� 
���'D�4*�KҞ3�r��u)��o���ke!D��qF�J�q��d���T���a�2D�����
ʔW�K� S���)0D�A�/�.+����
թHP���!D�����d��)х�4�	z2G<D�@ ��I:U�d�xW�u��qtg7D����-Qd͓��ޛc'��4�4D��
�MC��(E:�A	G{�@�5&5D���A!R�.�f�z�-��#�0�4D��↫��?�D���i^�Yl�"��8D��r����/h���G�3Z�Lw�,D���`��R|����/��vР��*D��{����tm�&�f�k4�#D�|����Q���Q��ЩL�DpZ�("D� �&��%����1��!p�!D��"��	xV��������ڥ�>D����Y68�t��lG��mj�b!D��`�'���<��T�13���g2D��邎� ��q��aZ*p��:UN5D��Xc�HE�������{�n���C2D���a���H���L���<{��#D�� U(��YZ4܈ᗠE�ܸ@6*O<I(�n�91�t۲n�s�.	�'��� �cּ4��.�pD����'�̜��d�%��5�B���h�~�
�'=��y�[zx�Ñ�]Xd �
�'瞭 �_>S¡�æ�5U=��
�'�2�WgA.%d������T�T]��'p�p� �[�{@�f�N
�mk�'Q�9"䞚Q.L��ւ�3�2-��'��<p�O���T�&@E8*�J]�'��dT+��N��gB��:�!�'�����+6��8a�
Ύ�Y�'�@��v�X�^x��jeB%Jخ}�
�'��A��gY1-�d$��1E س	�' �9�m��$��9B���	�'벬�@�Q�{'vEې���6`�]��'�D�P��\1�d!�-4/r%��'|��Ɂ"��m� xC0֤6��Y�'�4��	0$}p��b�48��2
�'v�К$"�
Z<dav�P2��eR	�'3��s�.Ô�<={�ʈS����' �Ppc\$6��d��u����'�1����+'4�����{�Uh�'.(��F�
R
|�k��@�[��1��'-0gh�f_�	+�Ƙ&MX��J�'9����D���|#��2G�vd�
�'ښaj���p�@��g"5�� �
�'aR��\�st����A�"#&M�'TY봨��w�Bɨ��G�I0a�'����"Fp�ʀ�U�^��q�'��]r��'>�B#��mr�'�Ӆc��5���Z�m^(���'5&��5.���0�z�j�'H�Yg*�2�x�	D��$_�1+�'A"|Q�ڻl����]�[@6-`�'�h�#�a5C�,r�D�"Ւ՘�'hR]�ÏתZ�"�J@�'�(�Y�'A���EFP �pɐWiC=t fu`�'&��šDvSnq�1 �X�eQ�'v�]{��K�����^)�y�A�oX�!��GZ�X=���غ�y�dK ��ǊU�U��4�����y
^�\^�* ƍ�Z���{pb��y��4N(d�2�`ڲf����w�֍�y�Ę�axD���gìrB~�����yr�I"a�.ؒ  �dT��mպ�y�	�Z9g�ޛ�f�1��	��yR%̂4����W� �����ҡ�y�9DѸy�«"sK �j��&�yB�P�e�hd�ʆ&:-3�OS��yRd�.S M��`�  Anl0�GI�y�l˧'��#�CFd�0j'FQ��y"�X�0�<�M�3�8�pe'��y��eV\�����4�b�+���yrY<L��� K�7#�.�1iX��y" N0s�"��VCI�*L��� ��y��ůk4Ԉ8�&#����c�U��y�a͖_
��������jp�Sӌ�y���A�ő���z � 󧆛�y�*�c��P�P��<gl�be)ք�yR+Ю\�\(�!]5w����j�yg�:5��P�K�5I����$��y�C�n�r� ��<�X��#��y��E}!2c�43��]Q��T��y
� ��H�g�+��r�FVE�N�`1"O���P��j6Ir� ��}ж�D"Ovm$ �,Ld������Z���"O�Q&���q�2�0���eg���0"O�4�󢁬H���ȚJp@yF"OV9a��ÅH�J�Iԡ�E]��r"O�M F��R$����@2?��K�"Ov�cV�[�R�kS"�|0��1�"O��3�	�0b�<X1�-S!l (�"O���
E7U�,1pO˷b ���"O���0�Лz�֠z`+B[�L!z�"O�a(�*2f!�i^%����5"O@ES���`y-*E��.t8t(K�"OL�k��q�
Y��@��l|�q�O&D���š��+����!	X�p�P��?D��c��јZ:���ոB�
�sO=D��@䊄�-u�[���2`��5D�Xk���' ʦ�A��؁��l3D�����s������5
"����0D�D��Ì��<R%��P$��.D�8���S#T,��BcC-J����1D�����)PМ��0���q�]Pa!4D�ԃ��@�6�4`���^|���;b&D��u!�|B���\n&� +�H8D��H�D��C�t�rG�{�8�UD7D�4���NI@X*j��;�r��D0D��s�U r:�d+�m�
jL��+.D�ܰ�+'[�Du��'�z�(,�u�9D���`o SҊ,pcG�>X��A�%D�T��e	|���c ��?i<��%9D�|�6ũB�x���ذ$8D�D�u��SULh�A��9�>Ȑ5�5D��)<n��@�B�։T�Uؓ�3D�D��Oƴx�d8���)>�����.2D���׫o��Qe�g��i�#�0D��"fŜz+� 8Gˊ\$M�gn0D��p'F��-�d��
�)iN�P��:D����(ҕ
Ur��%j�8m05ۃ7D�䚳�($l<1��.���:D�D�"1!􍘤�@>"�,��gn8D��[��_1���CTA�!a�����3D������4.2@Z��ߡ-T�11WD3D�����H�#R�U�ïڰ9(�Q�C�=D���@�"iƶ�����5��bcc1D�@U�^;+�\Ht#�$��Ң0D����'�0-0S"� �j��ӫ1D��	p�[� Cҁ�,8���Ѭ-D����u[ąj�	�=���
5m>D���1#ǽj# �s`��JC$���.D�$�&c�%C�>���e]H��We.D��`�G̱}���aN�-\�:P��j,D�y�V�w�`��O��n�3�+D����G��	I��X��)f�b��3�)D�d���DqI��"q���^lS��"D��ХLpjx`��1����V�.D�xB1��)'�t���q7(8��-D��	u�K�h�E�BF !a��"��8D���4J�p��a`��\1:R�9aG7D�T�c@��V^���עD@���7�4D�HA@K&���*��}�TD;��4D� JEE� &U"�c�iD>S �&n/D��`f0��I�mA�~��![�(D�����d��	��j���"�'D�����AŋP
8��E�у9D�� ��D�ʹ^m���ձ�~�#d"OT�q�̛:!���s�h<D��y�5"O����X,\�4]��E L���"O��CK£J_8�⥀(Hb�P�"O���D�)o�!8�$V�/U�h�g"O��!�5-i͉�bL|b⸈f"Ot��(�4V�e���שP��I�"OJD˄M\)GZ�Ɇ%��c��9�t"O�]ySc]� T%J���=����C"O�E����9R���C(V$�!�"O����H_J����H? �-2�"O��!��/9�֩���B��aw"O>0��ֈh���8��I�nj�ܱ$"ODY�:C�i�EC܎DU4q�"O@D3`&[�p`,�H�ǈ
[H�P��"O@t�W'�0cT\IP��, 4ްI�"O4P�o��B��T��"2��av"OX�)��D5�D)p��
�0��"O.�C���3άDB��ܲ�
l��"O*��$"�Y}�%�%��Wr$t�r"O�I��� (-"��H4����"O�̣s+�']�l��k�F 0���"O�tu�[�W�r����0.���"O��x��X�s^ܥ���� "O�ݠ�� �N'� P-
8�8P"O�2���B16-8�+��'�Rt)�"O���&(_�Hq�4�Ww�0C�"O4m�P �A6! ݣ/
Tak�"O��Bf̈�N2��@��2i���C"Ol��K��'���ж�δ-��u1�"O���dX�_�L(P��!s�2s"O��"�iY�}�ฺ,�ZU�x��"O��з�Ժ{~��Q���R�Ez�"OxY%��T��]�R	\W[�0�"O.\C���#DJ"����^�eZN���"O�����*�z������kB.T�"O� �T,�I��(�2�Ά2�6�kd"O8�o�G��#g�ZF�(�س"O�`xw�@�/�����C�P��"O�����2����@�,(z�5��"OFa"�%O8ww<8	fO�W��`"O�űDK���0�n���Q�1"OR9+@�N��H���V�Kڔy�"O�<2 gF�^�&��&	�[ƌĐ�"ORX�	�P>���i@�Z���k1"O�����N]�V���I��,j�*O�D�Ь��L1>u9�ϳeG(��'
�aH�O��->�+ԣd�]��'�>1ɓt ����`{���'�� �,ûm2
���m��ȓ7����w�Q�F�vk׈+�t	�ȓ0�5�!�'!n��ܕ\�ȓ^���Ap��dјY2��шyoJ)�ȓ4� ���&G�z��$Ln�ސ�ȓ"_hP��"
p��y`��F�J��ȓC�^%���҉FШ�k�k������dENt��݋w_�����&���ȓS#��Q�JBx( ���bDD��]�2�Z�"6Y{���eo�&	��@��v�%��6@7>�� M
&c�j���!����1�B8[s�@�SHP�c<lхȓ(#�Ĳ�	�%X��u ���8B��,�M8��V�)Z�9б	ۨi��ȇȓl;Z��O^%�+B��?�x���S�? (@��T	E61 E#S�(�Hق�"O�"��@�z��cGgS�Djt<�a"Ov�4��(��3q�S0?_괺A"O��@ĩ,"xUuc΃%oÂ"O2�����<�:�8��B#~4��"O�C�IQ��X��O�kb��2"O�͢�aۧ}� \9�M��:|���q"O��t+�*�`\3�E.uw�l�v"O<i��C)|
��9#Y�ԩ�"O�9v�S�pG�h�m�5��%"OYS��exfT�RL�x��`�"O� �� 䌵!Cn��4,�i�"O>4��a�0,�����57��xg"O��9%˔�1��;�B�x�6�1�"O�=���x0�1b"a�s���Z�"O�ׂŧ] �� s��-tǼ&"OV���9n��$�@�T��"O��K`A@��8p:v �,t4��K�"O ��E�P�}eJ��oL�e/�L9"O�q��^�uܕ�u�߷|"Of���="�Z鸳FL�I�#3"O(����8(���hR%�M��|�T"O�HXɆ�ɮ���c�r`6 �W"O�Dǂ�5.���b��[�@\�!"O��bWP� ���q��B���X�"O�Ѣ�Χw0�Q���"T�BZ�"O�9��J�|"&���R��H�#"Op	��	�~� ���v�H�"O��r���&���¡����r*d"Od�ku��6���DC��.�(ʇ"O�����߉HP����BJ�\S�"O⼈7"�nXrh���R G�$� �"O�%Z���ly�P��>N4�4"O\�2լ�!������O�|!��"Oz��",P1.��(B_�&��4"O����M�w��q�si�:A�B�:%"Oh�b��RzD����h�l��'6n�����u��`�m�3Y5~���'"h����!�Np��-�IT(��'Z"�ԁ�1^%&H�'�'9�bx��'""!����Ij�0��/��n� ��'Tt�a�mQ[*l�5�E,�ms�'�hy)S�S�&(Pؤ �B�f��'q����)̯����(T!ARbx��'�\`��bL�Av���`4�$��'��5� ��.|X	%��}�Q�']�2� E!{����S�šs�p��'�rH����	u� ;�/�h:U0�'�i��'�g�� 
��ɑi�~�i�'iB�#f�]�E1Z�����(W:��'��LX 9v#��	t���\����'U�<�пXd.��3�.i�L,��'5�ݒGC���Ӑ�޻5׬���'p�����ULY �HФx�:���'��$Q�S9>���3'�~\���'� ���CsHą:�~����	�'��e���}�   ��&`�~]��'�Ѳ��W7�D�F)�]�
�p�'��#��I��tI۶�?!���@�'H�*�ƙ0���(��0����'�����%i(���L� dp��	�'y�h�0��5'�<h6�ыg!hHc	�'�0d���@�T���aB/]Z��C	�'SP�أ,J)�����'	�vT���� � �\
n\��p胣N�,��"O��P��Z .î�Jq�Od�>��C"O��	�*����� &Z�:0�Q"O0�@`�6MA\�Θ�0݈T��"O`��g�G*KM�Y�qæ��<2�"O��i$�Z�eaER1GKx��L��"On����Z�)��#D��4�:���"O`9��]Nh�xDb%&�X���"Op9*���)I�PT�G�GY�z}��"O��@�Zj�ڤE��.u�Kf"O���W�K&% (2%�)5��QA�"O�tsc�_(b`�%cO8)[(8��"O��/P2R`vY�F�ϐP=T�;�"OjԋEE�$Dp}�g�='h��"O$�x��>�L%������"O,sW�Ϫt�,l����K� �'"OB�3�
 +�*��S1z�f�S�"OJm�E��Q�p�q3��	��i��"O�\� eOQ��HⳎ�� ����"Ol(�7A�(�ΈYP-�C�V	CE"OV����ùNɔ��p�V��5:4"O���J�><�5K��t�e `"O��(u�H(~� vhGݚy(S"O
�NO��8H��4j�qQ"O(-`� 5�J2'�<x����"O��k��~4��ő9(�i��"O��P�O�h�8���_)�� "O|
厎0 	�P�a�K-
Ѐ�'"O����Ϟ	����%߹$�Y8b"O�y�3���NƉIP�@�?����"ON!�ը��>
Z��q��g�v�
�"O�0
@#}(��1��Qg�p��G"O��!oD�5d��KG���iW
��C"O�óEQZݲ��'�]O�C"O������g j�����G���"O�#TK6(m΀[��2*
@��"O�0���i^�`  �[����"OD�郥ķOx�6��KD�6"O������Vz 1�%Ȓn���"Oz�[�,�{�آ��m�m��"OV%�`%�'�⢑�RF��%"O*l@�K�5��5GK_&cal)�q"Obm���L)J��`����.(.���"O�t��c]�$�d��0Y��a�"O:��%�	N����3�]�>:�(�"O��U`I]�`R�65z;�"O6%���_�(:��C�Jd�"O�Ш3��gPjA��E���.�p�"O�U9�`��:ʘX������;�"OJ��g��h�6e�G��+��m@Q"O��1nŴe��`[�"0(��;�"O&�A� Im�	(U��+ۀH��"O��I@�LK�p��Ƿ[��m�"Oܕ C��YX<���E�p��p�&"OZ5����̓�U=��X�"O�ɘs��]ȩ�7��=K<�J�"O�����*`���4F����|�2"O���?j��ٳ0 �=��"O�0�D�S�j4z$�$G�*P���5"O�x�Q�O�����&A� PXJ�"Of͐�l�sS !�E܂E��js"O#��w��g�V4q�p"O��ᅌ� W`>u2�!G�'"l�B"O܌ G�`�0���ƛj
�M��"O� �!����n���x�&MBQ"O����}��-a���Rv��"OPx��.��6��颃bڔwo�M �"OfA R1D�~��V0>��ң"O�lq��2��q���V�7(�Dx�"O4d����4�J���E�b:��"�"O�t��F�D��q����z���z#"O�,���\�R<.�#K�"碴�"O��+�c�.���pɀJ�,��"Ol<2�GO�m/P��%jU��]��"O��[�@=]v���8x�C"O~���$O��I�KV�|�r"Opq�ć�&��q�#��8���Z�"O�0J�F�9��%[Î֢G�e�"O��[�iH0� �C#�J��9�"O�A�7�@r(@Pb�μ�-�R�"O��p�HC4s ��3��8�"OH���� 
�(E��M�.��Yp"O��$�B��<��7H� X��z�"OZU��JqX"B]	q�٠e"OAЩK9��,s�`�^�fe��"O>�It����c/֥h��M�D"O�$7!ϰsҼy!���P�<Af"O��ˁl�?	P$(��X�R���K�"OZ�� �ǹx_
�YU��8�T,r�"O8�$E��
Ӑ��s.�@z�"O:�pd�E=]�����(R�@�u"OD����{"�}x�/O�uB*E@�"O��1���u�x�85��U: 8�"O\��&�E*,�t�H����
0���A"O��e-ϬK���B��Pu[�"OH4K�h�@5XO(q����"O0�f��Z���d�"O𶬊�"O0x�/Ϊx��f���,�� "Oܸ���V�ر�ҏxĤ��"O8U�e�S���HC�J�+�"Ot���׬ZCVx��M'R�~�""O��M�G�r��f&�-0�FY��"O�yهK^�^u:؁V�7��lP�"OL(�2��<� �f��}��X� "O��9�j��~.`�R���Y�� 8�"O���� ¥���@CΰT�@Պ"OjM�����X�x��$]�!׌���"O �җ�
�:%J�m�
0¦�"O��㊑F� �6BF�&���"O6��2� �c��-)T<�P��q"OH
ue�9-p����
�ܵ�'"O>��W��/D���*���	�8pЀ"OVd���υ*�(B�^��к�"O�t!W���1����&�3bpQ"Or����60��=A`�V/9`R	�"O����ʴ[��{��@1Th��"ODA�t������A�m����"O��a����"= a�>�򀫕"O����B����
U A��Z��"O`�P⫕�q��c6�԰U��i��"O�HD�)��z�
6��-��"O�M�'C!�����"MV��@�"Ovሐ�M2H�м��+���L]	G"O�Uڡn��O�!!AiHT=��!�"O�)�C��^�D �R'¦=��M�"Op�"t�J�<���y���+/NX��%��!�'����tJ/�����*Y��p��L�a@G#ߪ�`���S�? PUr���:�T�c�����!�"O<��!�d��͋P��U	>���"OD�J� "3���	B#+?�葐a"O�"7�O4�|)����&U��S�'�ў�
�AO !� ,�IWf��2�)D�����@\x]�6� �A����PM<��0<UH�;6x�"�<A����``�M�<����,d���b�lG9�|Tʲ��ɟX��5�&�A�g�8(�<qs���sp���ȓ�6�	-Z��!�OD"�:Ԇ�1��D���_�
j��O�\sX��Iw�'p�Q%��o6�`"��� i@\
�'�nE+�`�7��ɰ��_���0��'J�� B����Q�/N���\��'Sp���E� �`���ލg�-9*O�t��ɦ-0�a��*I7�0�V+VT4|B�	�Hn���.+��U1c��&\?8B䉎@Jz����B2gʅB�Iӻ*��B�	3C�X����X6/������'֦0#�'))�5��=���*E�' 	�y˓�(O:��C�
n�L�
F��T�Tt��"O*�z�HA1M���K�gԙ] ��d�|��)�Ӑ $`͑v��5��A��D�`f�B��
�h��,;E>M�@�A�b��B�ɾy����	b+�xkB� tx��%�I�B���sfk���ȥ�]$t�nC��Rj$�ƥ͘x����wz�c����	LT8�B�V��IS�#�C��3#�� ��ӊ)~T�Sn !M:8��'&�}��DЀX�]�Eö����0?A*Opq�u$R^R�Z��؊J�X�2G"OL�B��A�k�j�Ff��ܘ$x �Df�T���'^X�!P��Sxlh��W��7��{<A�"�4	c�m�N�L��eΓU�'Sax���Y�8ݑ�E�1JIi�]�yB!_"���f	�;	Xu���M$�?Q�O��d@;=v���^$qBٓ�ЂXe!��J�V�
��$`�*;W��q��Y�!�D
�#�P�ۅJQ5*�T���+�>�!��O�p�k�EQ����+jX�|"O�a�r�G�C,
�Ⳣ�;@�]����)��?��'���hp㍪	�%JƏ�u䨛�'�|�8'�H]&�%dT[�b �-O�u����b�g�|#���Z�6���(D�ؓ��H��и")�33�ܝ�7/������OZ��'�ɧ��'�(��cF}��D���
lw��	�'����	7]��^c�P\����O07��p>馡Ŧ-�-rp.E�e�<�#u�@C8� ��ችn|����ܝk��`�z��C�	�'\xc�'F�=��Bގ#^7�3}>E�ܴ+ܪE�L�G�� Ӄ.�(��Dt��zM��K���hJ�r�����$�݃� ��"Y0��C�d���?a�n�4@h��ԁes���$En�<��G�\��e�Le�D�Ţ�f~X��I�>���D��Z]���/b��R��!s�!��Ȑv|A˲�G.U�|���d��1Oz��w�)� ���R.Jlȹ! ��C�0f�@؂��!D2�QA�C2X"#=!ǓkrL��`S8k���t�	��\d�?���~����.����nI*o2��r�>������-9BA�j *�����r��(��"���dEf������Kq�2�m�?�<x#ȋi�(���##�"=)�S�? �����FV�4[��2$)`i�"O�U���3)x$M���ڱ���"O��0d�Ѻ%��H����;` q@5"O�� )`��A�U*z#�mb�"O �zpɈ7���6Q+��H*�"Or�{�oUM�,���ܞ#?��*O�M��|7��z%EЖ�t�Q�'Hx!�j@�H�n�85����1��'�HBR��H�4E��$��'�0��H	� ���5D�� �' ����0M��hb֊-��qK
�'e��2��L�3/`�1���(��A��'{q�����=� ���� �#�rQ��'��t���M3�5ˇ�ۢ��a��'��i�ΐ�q�6��@R��d3�'�权Q)%D�0����R��I�'n5
�-4ܬ�
� ϖd@�'�(��@�ӑ93<���Y�.��<
�'�&��)D(%��(�߯-8�@��',��E��BJ�e�(0�0���'O��"#�2�b񲕁J��e��'t��;s�Q�h�x�BE�
�'��$����N�$Y6mXy�	�'��Qfe�*�L��qO%(�0	�'��1�"I��:��p��@u��3�'���� e�
y�6� �Ź^8��'\���p�XI�Ё,	0Δ�'! � u �)�,�@�$�3}�Y��'1�4��v�0��Ԕ0@�;�'�(1�a
R�4&łf'��{���'�@��0q�NA�b�ުl�NIA�'e�i��ܡ\�>|ɂ̻]J���'Ŧ��L�!��D���Ǣ@5�9�'!H��1':��A"#�!�h��'L��1��#�x�A�h8��'>2��4�3S.�#��;�<��'�(͒�������(��7��1�'^VP��FT+`�����[.cY�'��ѓ����)�,E-u,P�
�'���rP�W�|�L�zŠ������'�qڥB�P�aa�G@$x	��8�'�&)���4Q*��q�A�GO�|�'i�9h�J	�[E�����̵)Ox��'ժ�� �˻8[�ܳ�J*Oʖł�'S�� ��".���P���1��'W��`�ͦP,X��!^8"v�#�'v)���U0��;��[4/� 
�'�����|0Rq�gȉ�)Q�=�	�'
����Rtǘ]Q���'��l0�'����\���`!Pd�>p���'�̘R%���8��J% �~m#
�'�@��HN�fm�����[��~P�	�'3��B'`U��~ah���3'����'4�M�Dn����bh��&��S�'eV4����m}���EXg�輣�'���*�.U�)��R�o�j�	�'
6�B��3���ԛ2����'s$mk�A����0-1����'d�9���� b�R�B>Ev� �'��ia��L�o�x4k�B�"3���'������kjAЅ��?!�ֽ��'�~����xq �DQ��d��'�4*�-De6��a�>�� ��'=���BD7
�� 3 ["3�@AH��� ��R�y�@z�W,y\�the"O��`m�e��X35��*@>$5��"O�UI6��A \��a��.�<Yjg"O���&�{ǐ �P��
:���"O���W��1*�#�Q�'��=1�"O�`z�.V�VA�×�M2M�Z�PQ"O�ī
N���8�CM={��l�U"OR�JOC z/��0��0Fp��q�"Or���g_6O���	ao(1�#"O�yZ$�9d�x����
�Ҍ�&"Oƀ���� >�:e2E���}��Ex�"OHa����!)Zy d��'0t"O�"���/qt@೨�9$�$�2�"O� ��<)�"X� eİq�����"O�-´F���h���I^�)�	s"O4ҋ��Wuf�ׇ�>t�N��"OA���;�����,*��`�"O&���DR��e��r=޹aP"Ol��fDS|!��j��Ge���&"O<����%�qa�%�&	�����"Ob�kAN��U�$�d���r"O)@�L��V%����,��\8�"O�s�lL�$�cw��6��ѳ"O^�1���Hӈ���*_���*"O^�Ѷ�$P}�=�4&�j4j�"O�,"/X *���V�>WV���"O6ȣ�X.�Z���̅�oD�%
F"O���C��\�I�
Br-l�� "O�y����w�X���e�,��"O�聤��hT��ɖƄ� ��hz�"Od��s��\�$K6��&n,��"Oz�H����i��4)rn�whx��"O����?g	���݊e�hX:A"OP
v��%wc\��5+�M놜�E"O�h��VB& �!q�JXz�"O�u���*�F��7���?�&�X�"OD-1B������M�R���g"O�̋�81�$�B��W��B�+@"O�a� /�bE����/�4�"Od�x'�5A�$b5/��&�`i+q"O=9�,�?tBn�r",,����"OvQ � 
K�D��1㕫Zy��"O���0$pOm��$]c�0"Oh��-�=hS�$4��-c@A�"Oh���%h����+*) ��0"OF�Hb��\x(�S��#�0�@�"O��)!ɜ�|4�d�P�M��t���"O4��*:w�M*���4�"O�ܢ���7wg�TɄV9�bʕ"O��Q(�-��2�k�h\t�E"Od�+�*b�:� :.mp�X�"O���#��g�&�z�j�T�x�"O0< ׃�G ��)s�BE&"OZ�p�͔�i���Y4��&��Њ!"O<��rH�G$=�$V$vq��hr"O�v��=��2����Xjd�
�'P t��g<&�L �+�z�9�
�'�N	��&^�iY�Р�B-n�����N�}Y�H�ŏ@E�E������yBl[�Cf��%CV7]��Y�#C�y�AĔV��T;�,߈J;@��C��y��'x%��Kg�C�Fҹ��Cˢ�y�� ~��[��ҫS}�b���y�EU�>"D��l	P�6W�y
� ���S���p��L����a�����"O�5 Ǆ�p�P���G�!?�v0�s"Ol�	� ۜ6���Fޣnx@8"�"OXD[���Ṳt���Ժ_���"O�k��^[����e�<c*]	 "O�Y���#S岵� �P�P���"O�ܢ�/Џw֞l��ܩDVQ;7"OlPˇ,�G�(, ����y����"O�ȡr�'oP<}Y�-��)���0"OT����tU��B�Y����"O|Y�A���t��c�͍@%l��""O�X O��T�$$�p�]?@�r7"Oҙ�A�I�^����-��� ��'��'C�����������V�R�ҹ�B=D�ܑ���?lڌ塲���h����W+9D�8J5���L�|� q�N
 ��a{��$D�;�=kl ����m�u�$D�ġ6�F[��	���V��X���4D�tɲbFq�ܰ&�H�6�<4 U�0D�8�b/��[7UK�Ȥ{�ؐQ�0D����[������">���Iw�;D�`��,�$�B���M��z��4���,D��h�n��:aP�"gϋf��Q�N)D�[�␸D^E�N(l@��!<D��[R�	���E�R���y%=D��@�
�ڽ؄)�	<�X�����>I����D�x] �J���j����.B�ɺ1��K�C؃	s�m����)��<y	�C��55�������^��n���~�'|>x8���sf-Іe�5$Z���'�Pi�g���EC�_�`��8�
�'�J�)�D�|xR�2��וt�'�0��u�  A#R$(j>	����0M�nB䉢W0x��rl�38Z
��^�C�IY0���B�[0@�,��,б<��B䉍}��M�.#z�n�B��2M�<��v���1m	��쇧'׶B��kf��faD�:s�kɌ5���D-�� /�|�+u�S�:+&�(� �??�B䉑0��9��B?m i��X�#��C�%;`<��-�yNR�1pnĜs���*?�W�?L�I��1R��\P�]`�<�'@���T��L$ �~��Mb�<aCm�@B<�a�G�% ^q)���B�<��]�U�
�3�ğgF����oJx� ����Vd�di��K�wi� ����#����ȓT�΀���*�ހ`ViYVb���hd
���7�ny@�e��ݠ-�ȓC�*���BDB�V�ɕF_j�݄�Kv�M���nA�aцF�(vb5`���s����F�Q-��ö�S�8���%D�����^�ݐ\?P��c�Ҫ�yrFO�5�И!rk��:Ī�-^�y�NK4|�& �GXU��CL�yBo�p8�!k��d��`� C�\Fx��)*���%t�Rq[���VR�p��H�b6qO��)�3}�,��z+�Y����<�����`S4�䓋hOq��T��'�$�4�YӦ߇MZ<��"O�B2Bt�|�҂F�-KL䀵�'>�"=���$�9��R����`L<���CQ�~ !���O��keJ�*ti��͌&<Ԛ��IQ8������0xmxXG�Z�I�4��q<D�lH��ѥe��� ��/0NQ�@-5��p<1#����92�A�A�0I���d�<� 6"�A�C����B�X�E�"OH�['����İ0�R
Z�<�D"O8%��_<Gth�j��T���%�p"O���R�f9����n� �`�"ONE��ʄ2O�ι�7@܄
���W"O`زC�ʯ-�6!�C������$"O��z� �� x��(S�u�.	!"O�[t-C�8͡�!S�����XmH<I�@ W�����ZB�\B��J�<�a�����H�1e��L�<���[L{()�S�X��z�� *�P�<����3I�R�`E�ĞT�0x�sB�d�<�	�_[�Ap�؂/
X�HU��b�<I��H/4ʆ}�SF�X���r5�a�<��^P�Pc��#S��p@�+D�Hȕ��X�.2���&�*D�L8a��}v<�J�T�w�����k6D�ȩ%[�]1�):"(ѣRkH%�Ub3D���'�ڮT`��˦	C<?dd�V�#D�8��'	"O�5��
�-�(��P�,D�$��o��@��ۦc;��fM*D��� Jќ
YWk^�/o�\7'Z�<A6��"b,�1BפƩb��-�2@KX�<�!]%M�B���ŋ#Q�����Q�<A�Ñ�G�r����Z���ڃ��M�<	��ܧHIG?y>��� K�<�4m�*�XT�aF0��$B�&l�<a�I7��U�v�I�X1^���}�<i���m���Ё{�&��0��_�<�P"Y8ʐ`�6I?&��t�X^�<��N3s��X#@׆�J�࡛Y�<���,�3�F�'�I��n�W�<yv�y��"�V�n��]�f�g�<�Ң͇^��YRꊒ^��ى �f�<)"��k=��2¦�}�V��k�L�<��G�8%��l���GC�<�������9��͝� �a{ �z�<�U��p)��p��4p��n�n�<�Ek�y{��YPiڶa��l���k�<��H�z�>�A1�H�u�J��k�<A��=s(t#gA�<~a��g�<Qg`I�e{<�8�G20v�y։�N�<a��	DF�����8U%�J­�S�<m���tA#��e8dEҐ����y����W��V�-*�l��ǅ>�y��Է')Z�p	B1 !\��&���y�Ã>	B��A&p�P�C�lO#�y���H,$K��:_�ePi��y����lr�����'^�̀�G�>�y"�'r^�036�N���	b�h��yr-˵T8�	���4-� �� ��yB�&h.X+�b	,P!7Ȅ��y���:4�p��c)�rƁҠ�y��Q�/�ͫ��҇J���E員�yb�M�c��X���D����!�y"�M� 6���o������9z�䥅ȓ*�I�.+����L�V��E��=�aq��$��ʜ#(�\�ȓ���D��?-�n�ɌyP�ȓ-�ж�ɔ>Tr��v"W�|�6܅� ڦ	���X�nǀ����3�x�ȓk������_2p���jD�	1G�X���K�� Ѓ��9�8�
Vo_+$��]�ȓy�Ȝ7!ޖ5I�s<h���S�? 8�%	�T�
q��`��:�)0A"O��� 
� �nm �NY3^]{p"OTP�b�Ԛr�he���	Jێ��f"O|����_�`D���ث3��!�"O��@���O0�����&n�੄"On�{��P�F�x�
����S#�1A"Or�8�N�3nvxI:ǉ�e�@��"OP���!�%{�b4���O�U��u�t"O��:p�AI�\ʄ��{M�ɑ "O��8��=K48ʐ�� ���
�"O���+I#\�t`I�eXz�C�"O�d��뛵"�e���N2c��qR"Oz1�@��1IqHԈm�L�"O�Ub�m�~�`��g�3�~xG"O8��@E y����	"fd��"O|��AK8O#x����# �@xp"O�X�1C4t�8��?*���5"O,4"�oC*tr�X��`ȋ��H"O��8�F�d���&
\�u�b�W"O��b@[�a�D� ��x�DB�"O��� Y"��HS�aŠ��@"OfhP��9ub�����"��-�"O8)�s�Z9b�âF�7jxl�0"O����I� b��p���&
�"` �"O:8"���\R:E�`��D����"O�U���4 c��p䂏���"O~���.��X�4]�eD]40邌1"ORtqO[&�����j�d��7"O��ђ��UFI��v~:�"Ovh�ӫ��W��!#�T�",�"O�Y��n�&( 8%0�kZUU>x��"OL	K�̘�K/���aJևd�ȕ
�"O�Y�E@]�\x(��t���tp�5"O��t�-$���Z&Kl���V"O���O	!,rjhzeR;S�U(7�'�@��� �sԱ�Ïƿ��P3W��`X~X�Ãi2@9�ȓQbP� `]}�5qW΍i�$��m��DB�1eZ�(�D��!��ȓ�bL���h�<� �8T-��s�*5�W���+l\���;!4D�ȓc�����`V�v�p��0P	f�����	7�,G/���B	��؆�JRU(CN��{�=SӎH�9�Jԇ�0�"I�4"�:+�:w�;f�ꁇ�U̠I夛�Q�X����F@p��ȓ7,L9yB	=^j�]��ǀ� �ȓ B !��LG�,�V �͆0�6Ąȓ^���R�MDU*ly����@�ՄȓI�"@҇O�"3p8Q�IG�U�x�� �\��ԥ�~�Ҕ�ՁR� D�1��^���p�O��f�8W��\���ȓy�H�R�JU^�bǁ=:�>���7ۼ�)�@�:約�'�  K=���4���pC�3mu�(�S!6���ȓY�$���ڀd� �!Qm,@x�����Ze�V��LAP�Ӓ[.J��ȓ$˴bP���U\���F�!P�@�ȓ ��t�V��8�P����N��ȓo$Ҩ�S�(hE��� Z�,��2K^pC���m8VukA��3>B��ȓ@�����ȹ�&,���@����ȓi6��@Hd�t��G�P�0#���DWРp�G�G��=�7+Hs��u�ȓl�89�)�U���1*�$��=��S�? ���@G8E�8���h[�3��y�"Ol��F�:F4���S���`N��S"O��A��?O
��zw�����S�"O���f+	��U��ʑ@��Ժ�"O�ja+��:pbc���6"O�\p����&�:gGړE�^�k�"O��i�LQ�!��&J6W�
h��"O�0��"cTͰ�#� �"O��a�k� A����S�"�2��s"On���� :G�r  G��� d�X�"O&��G��%j�t����� !*�"O��a�p;t+F��m���qQ"Of�"dNR?�����+	�܄�"O8x�1	��Ln���E"�}�p`�"OX aD��,-�}�K�/`�q"O�K�J�~�,0�+��L&!@"O��������[��I�3O�\ia�'��8c���<Q�
��(�ZHdwL�x�kYt�<���	B@H8���T�qG��b�q��ZB�48�����"}ڣ&��W�\�+�B#c���7�r�<��/Q�K�FLz�K���c�5.����$F#� �ڨ�|�'�0@�gK�t�زCًKHNx�	�'[2ӳ��c�4�AB;��åe�<���&��&�����'��ePUIV�xŪ��B??��h9�bV��`a_�IE��Jw�C*Z��d�s�C���R�� �����'��9wm@�M
xr)�I�&I�M>	RI��K�(iصNQp�da�� ��.�X|&��4W�����@R�8FC�	?J�J<�r%	�x���ǤE>����E1,^�,���-]t@zt 3�3}�
D4,�Cf�e����j:��x�G��-h0P�"ƫq�`)cO�%]����� �&t�BW)��e��U���'���*�+��BbԚ�f��[;���˓�И��L��n��g]9_�|�ٷ���i�l����M���K�Px��ڂBB��($�X?v��(
��.}�h��j��h;������J0;|�y���#E����y¬֨u���/��w��� #�i�|�*'P����Q�*�� 4x�Ў���>����1(����N�6�x��E/KrH<�G,E9m�����Ԉj� i-r���\�hon���E6~����AWL8�D*FL�6'�E"U�^�]vy�t�1,O�j�?X�� �P�Q!L̈́]��
�4a*��C޼
�f9���N�B�� �|�CvV�!���rjO=' ��'6F C��~D�!� �uϢ�W$�ӘQsH��Y�O��B�̍	=��B��!��)�Ӏ�:]�5�0J��3��H�j��>��o�3��<���>�E�	7K"�F�P�(z]���I�x��C��$�L�����-�&��(J���h�Y��!0���{c2���zX� ��ߖ;��a���">Jb�{v�"O�tB�f����eo���G��"T�{q�� hU3d x�jB�I"?�� ���0����K�<�'@᳁*b`����2��ɖ%*��;4��A���J�#˹m�!��C�|X;�G�	a�*01 ���[4JF�sT�8���2�@���)�ͥ;	>pQ(� ���V��a����R/ڐBAòj�y�$Ѯi²<�b�($ ����SN��+,O�:��D:=�f,�.?�b��s�'x(�p$�\�(t��:a�<C��f(ʰN:(E`\�DMH�GAh<1Ӆ��H̆����̺h��e�Yk≙t�2L1g�W�Rn��B	�}�P�Νix���
eѮ�Y�"OB4�AH
4�jВ�Egˤ��-�t�� �mF,[\t`��گر��'ܮݛLA3]Ѥt��#��ff`	`�'�����gE_�Ёi�=��@��ԽzX��i�3A2��oIe�ay��?v,�B̕�uA�x������p<A��K0Tz�-�"iC�#H��O��	�&�qS�5Nl��Sad��.�v؃��؏z��x���q��t��`� ���QT'$}����!��cϋiO���P�/9���x�S��vgl� �	�PG�-C���6>b��p�"��f�=Q��В �H����b��vd X�c��,	t0���\}���
�P�O�)���V#fo��B��.�r�+C
O�B� �	0t�(c��jӐF�4쪤n_G}|�Z�`_4�.$IB�ȸ'�� �A�~�ně/�����&lmd��Z8�TZG�[����H_a`�3��ϴGd�)@`	���.�8����7��Tc�{�(@�z|�c?�p�����@$=��hs��8;��u�Ox`{�&H�ura���ҕ5�<��'��C� �[3�����ӸhX��e�o�<��I�y�Z���(��~��9��݇0R�%ӷ�9_�,�g�ќc9�m C�8��/"9ŉ'\�Q����0nHi�jN�2m���'oЕ�w�Ԡ5�$<�uɓ�E�L��%���|RBsOñ\�0�z���Xx���@ r�v9"S�Nt�&՘�i,<Ot5@�w�(ɨ��̮����"�>!��J'R�� �?D�Ps�(_?]��-�!f�!��\��E!�D�' ��Hɲ�A�%����u	9�'2T���2"eC��8���|1x��I�L�2�71�]Ȳ(1�j ZФ�(׆LjC��lvc0�g~2&"�z�HfEW:�̽A�h�?�y�F߆[�䚦������`gT��M�P]��ia�0|O���3�G�1��+����a���'��	� � W}�U�uE�QkP@L�q���&
�b�<Q��*�$�a/P�?.�HgP�<y7IP:L��y�T��vT쐂�v�<ѷ�H�PtΑ�j>~	�� w�<��g��f󒁗li�=�N�m�<�M�*I���2/8CcT�B+�d�<�0���~W� ��D�����YG C�	�u����D)V"ʘ� �,�JC䉫e��@��Q���A"��4?�,C�I�h��hfe�r^�T�L�9S_:C�I^��UQ�Ě�T�<I�E�V�wC䉿b$���M�o���#g���0B䉆#j�r�ș��� ���C�!d�I�G*d!���l
�+��C�c�lp�3ˌG�k�(ȹ0̾C�	!M��]r��Ь�`9�B�	�d�XB�I�.��ъ���<�Hs@�"C�C䉠OM��	w���[M*!3���1J�B�	�#�4�d̾86E`���&h��B�Iy�^ 1 �ֆV��5�PeH�UX�B䉧K�<�S��۸}"�Y趍�E�C��s���{񠊣 }P�RkСb��C�ɽ.�hT%�4�M��	�BC�I�p��Q��r��Q��r�ZC�I�^�|����$�����~�>C��,o�(���_�EHz !��K�iY�B�	!]�\pY0�D�ښ�S�KU)?.�B�I�J��1`�D6W��S�f�B䉁N$�ܸ���;�FA��ѷ>��B䉓5Y�ã�
pX�&�.B��#Q{D��r��rZ6uR'���6B��$jHQ0 X��8Q"���Mh�B�	|�m���'�[h��lC�<BvH�T�φo}̀�"�0e�@C�:*���d��!q��	��׭<B�I��h�7��:^C�)�U�I/�C�ɦi��tBu����d|��C��H�C䉤I�Z�0�%�N�$��IS�%��C�
9��B�kѩ)�^�3��ĻGĄC䉷k�5h%���
Yp&(FC��f�D�f�H>��񢦝4(�6C�I2-Cr�Z��*SE��IT-��[�C䉸|�ȉP��R�8i� ��+s��C�+K׺���%J9VB�t���ĲF��C�ɔH��	P	� p����C�,��C�	�9#��ct��_rn��b��UnFC�I�:a4�j6*R�E���KA�u�B�I�EV���I�n��m�S�_�k�B�)� �񣄆 T�80(!�6Ŋ��"O�d��լy��Q(#��OC��"OҨ	T��O�i��K�2-0���@"ON�넫]v��!�UQ>��"Od0��T>.�Bbh�QLx�"OhE5� �U9������4���S�"O�(EG!'2A���p�i��"OP�!η+	 ����1�ʬt"OF��D�]K����oGP:�"O��s�/ّTH�`�W��(o��H�"O�2�nރ$M�A�̑�s���$"O -�oM�tX�� �do���B"O��DEɴ�v�"�nD���"O:�36�{�db��"1��	�"OJ��&D�!�(��G�6O!���"O�yy�D_;X(������0��"O���C��;��!+���\Qp"O�r��B���*,	�WV��9d"O�T�!���V�Вl{X�ڧ"O<L�ю��>)|�Q����Q[�T�U"O, s�!��T].4�C
��3�p
 "OLYX .��W��I�0I¡z7�}��"OD}ygl��o��J�R"���"O0d�� =\$4�@	K+"��"O�H
%�T)R�����ՙf,*�D"O�j��
b� )���O�]��"O�l�un�"8�m{ ��^��#W"Oֹ񃩍�O�����.��<1"O��Yu ȴE��bV��+XJ'"O�4Y��f{��bbbœ����"Oک �ĜR�B���D\0��u�"O(A�Į��E�z�1��5>�zu��"O��Ԇ(5����#�z��r"O�HU�	�Թa�Ag�|��"O����KQx�,4�q
�+7S9zU"Ox���
��e�X����"� A�"O���$fLvؼmЄ$O	2��"Oق�k�8�\���� X 	��"O<�b$����1n�8����""Ou��#$Il�0� E��"O0�����M����� 9�r՛�"O�չ��^�N��c��{d��"O�����\��RI�ӍVvÀ"O0<��B }���#yFD�6"O�����H4���ͱ8�`���"O��f�Lb4��)ʈ`��"O�QYG� K@B�Z''�-��Ń�"Oz|J�$\�B&hl�����wn*D�����A�{�V��3�f`^Lp	:D�Ċ�FS:h1��G%A`P�d�4D�P�r��Z�.y�P�B?@�Md+5D��rB�͋����@��j
�*��6D�����K+:�a����P�N.D��Z���~�(T��.*1��AG;D��(7�>�x�B"f�'2��$�<D�T�cb�?�� p��5b�:a�":D��!�� 5�x��ی^<���E�9D���]�~ȹ��
��S��3D�����=WO�""�׼x�r��3D�l�B�:Z
Xj�-��/
@�{3%:D�Ը�m(r�<xr��[�n1Z��'D���I�
Z����oJ�^��J o&D�p�2�/?ɼ�+p$ܧ���ѯ;D�3"$S�J�`�+&�]	/��R��8D�� (D� Ǌ�T��у��+z6h;�"O��B*D�͐�H2 
�ai 5��"OH,Ӕ��
��|9�@���V"O���&ښt`&=��꜌W�^]�"O4����&p$.�$���<��01�"O�lb�Ċ�oVT�I�FԬxyFl��"O&�#�V�>n����%`�ƀ��"O�x	�.j���X1�m�$�]�!�ƯW�~�(rHŋW:�Ճ� �!�L��s���ZxJ�s1ܘ8-!���c:%AAh
WQ4�)�a�f�!�X�5�R}���6PJ ���8�!�$V0L�Nl���%3�J`Be�aV!�d	 �.Y3ӧ�87��(Q��4�!���s�Z�i�c��2	|`�%F�?ec!� �K��S E�*�N�D'S�!򤊷p����`+�d� �q�!�э(��H�
$6�D9���H�M�!��S�|��Ō�
��(���ǁ2�!��μ^|���>��"R�T�vp!�Ձe�ƉQ�H������ׁ&,!�d�dg@b��@�d�.��t��@�!��C�aZ�c��5x��Pd��!^�!��-@���d�$Oq��C4��5!�
q����Co���%m!��J�Zr���-��SK~�$i�	�!򤆍i�L[ჟ/(4�@ɉ�T�!�Dlmn�����+��ɐ˗?'�!�d��7l(@��ͼc��)��B��!�$�0ALT)�bM�i�4��G�.@}!��ʱrE`�B��
��cņ��m!�d�Bh{s����Y{�F=`!�4y�l�FA�L����ǨZ!��%$��@�!)ZV��B���D!��A�0s�ɍ0'��$`��QHW!�[�"�����[9�$Mʴ\W!�D_�|?�18q��	US�&ojB�I=��9��K�!�C��#:IjB�I1"�f�"�l�N�4���E��%�fB��=��,ȧ�;w�ް�6�	D�B�	��X�BB������Y�`B����`#����``8rkѠkbB�0R��c�\r�~�h`L}�TB�	/V�z�a��$((9�aN�^9(B�I�Jm(Ir����`Hha�/��SHTC�	�Z���B�I$L��!i�OVC䉢�2���I�l��1�ʖa�B䉕8�<�%i�:D<n�)S�ǟx�4C�ɒP�ڥ#��l�f��c'D7P4C�I��\
���M0@Pc���37��B�ɠ\�qp�"|R`)B鎺)fC�IWֱ��H�,t�nH����?�C�ɴID$��CgˑR�<�+��^�t]�B�I-Q��P�lӘ�@Z���#-8�B�In��t
�Q.�40�F�:�FC�I	�����B�Z���AoG��lC�ɦԭ�5̌3Y%�����7h��C��!J2| �m �`E�|1�L:8рC�	�踈�%L-z� U��
�^B�	�� Yႌ
u�(5�S H�L�hC�I7EN\����R�=�.���[�@C�ɗU� �rfϟZH-�*�B�	)!�ڴ룠�'��YRW Ե0O�C�	 �`�G���Vx���s�R�T�C�)� ���5T�f��0Ņ�"l�2 KU"O�xi�Mڬ	��͉%*Ɲz�"OL�s��8y􍡧��D��1"O8�c�Vq3D9 �N�;E�1�p"O$5┈E�2��Ȑ-�

��@2"O�uA�Բ2BVqp���
qG�����&�����X���(6�B�cx�ȓL�Ԡ�
%X�`T�]�H��Y羝����<\�R�pQ(]�~|D���o>��� S�(,��m��jE�ȓ���`Җf���`�K�ڹ�ȓQ���j"o̡Y#L �� 9�ȓ#Y��ߍ^���9���Ʌ�JQ�=���� r��@��fT�a��J�������9�ӎ
�3B�|��{ׄ�9B�]�<�v��n����2}�܋׆C:e�&]�����Y�2��ȓ6�����j�H�B�D�&,��4�������c���a�"q^� ��2�U�"��7�$�� �LAx	������7��� �b�]�&H�ȓ+z�"g��k����Kh�؄ȓN�e@FA1���0AS�<��U�ȓ;h�ّ�06^��DQ��i��| h]�@��<R�L���	+��=��&�:�*����r��ȓ8˨0�O�%��zԬ��J����A:|�a����|�bQDP�v8�ȓ{��#Q�.+DQ����;#Hj%�ȓ#���X���@���14���ȓB%b��@W'��}��A�)�l}�ȓ$$Z�z�)v���cGS�G�����89lAa����+K>P�䉅��t��#�Z��I+����h���ȓm'���Q�дY�����=(����-��\PS���N�b�"�Ͼ{�*T�ȓN�zi�Ĥү2�<`��NwT����4��зH6P����[���ȓN%�q�@�]�h�q��:%�X���Ǟ#!5(��� r	�� ��:D� �1%�9 �Rmi��m㘰 �.;D��X��ˉo6�Y���%5����r�%D�T��+T�(�45�����i�ؐ0c�%D�p��� r�YI�@���kA/D� Q(̄T~�#�BM��x�h,D�X���4!�H)��5`JI�wm(D��!!HK'4��:0%��{���r,'D��rC�Lɪ��6��.
��J�F$D�d��j�>�Q�5��1z8�`�3�$D�T"�g_ *�%�f*�3'���� /D��0C�'|MȀX���\I����-,D���i&q������@0�x�ӥ�+D�pPqC�y���B�a˨\�F1���<D��h�I�����7ȒZ�ĝP�9D�Ts��ǍPӢ9)pG�"��yht�4D���"��#�1�R�bC����&D��2�Ǻd 4Y"��U�P�g%D��pUm�"�HX��� �DDB�  D�����0{D<ZT�Q@�P�G�2D����\L��Uk��R�b�:P�w�2D�DӴ��!�ҡ+S�1](Ne{�A1D� h��ϵL<�}V���RY�*D��3�E
)2��Q��[�_�$����+D���s'w%2��u���M���f�:D�� ��IBN����Y�.׬h��4��"O�q+%#�"~L�49��,�L��"O4,� � �Mڄ��Ǥ3�E��"O��pc΅%v� ����K��-��"O��W���H�I:u�ǟW��E��"OHejTm1}Dj�8�嘖AJ���"O�J���1|��3�k�A2$��"O�<�c�L�?j6
"j�>A-��"O���jH)"�^���]5K�i�"O�8�rŎ � �w�Q�?D��"Oʵ(���|5Py�a�Ǎ!zhZ�"ObHР"���@�[�kG+m)^���"O�����w�8����UMt�3"O$=9�K�x1n�P�M/*���e"O�؀�W��<���FT�@-|<�"OzXr#+�v��Ao�C���"O��h��� '�`dO�h�H�`�"OB�@u�˭4�^�"D��"�ID"O���/*yf���6'���"Oey��O1s�,��o@X����C"O�tie�>���Y����Pj��v"ON��"�eٔ��箆hd���3"O����ʇ�[�\� ,�$~^ĥ�s"Ot\2T���>@�Q�+�'�|�{f"O����oH�X
.��jċ)��X�"O��KJF��JEJ��/A�Z�@ "O��%I�>[���כij&�е"O�m��] )��	n^" V�"O|ei5�T�8����?	IL݁&"Of�㰈́w��`(�ㅉp9*ȊR"O9A"B·W^� ��l�;?ڔ@"O��c�/X 5{��j��Y�2�!��U��У�D�%���B`)C�!�$�Wr<i!LZ�P��J��d�!�d9t��3����0��}��X��!��r�M�5��9���r�mƲ.�!�$52�$�c�� :q�es���!�$1���i���6Bt���ɡ=,!��M�{9Zd����1�Ȓ�I�u?!��ݠQ��C��5U/@ BG�(!���u͆��ɞs�����FF�Oy!�D�Hb@Yɦ�C:/�r=S�E��g!�ġh�P��P��:�jl�3�ΪFk�z2G�#����SjP���]bal1~rL�厘#�
�kE���#��ceG[>)s�(rK���b�9o'�-;pA??��J�r�L�SN>E��"�	:6	��*���;0��"e���� c��ܢ���)�'NWtH@�g�h��l�4{���de�4%}xN>�|�Lʴ{��Χ-�!$e�(g�\t���I19���犯<��O�7�n���I�Ob��[`n��}$�0ҍ�è\TH�8�D��WB�O�4�!��A�a�t�U�%H�m��
���M�XAa@�'Є}	�@a��`y������,���([li���	1M��"Bʪ���r�i��d�Ϫ"��<%>�0H�|(�y�b¢u����0�$�E��3�-"��I�=���k{,Ω�'��8Y��I�XB�kan|�)�4����	ȌE
�$����hoL]�F�y�"��h�DSV�'�"
`�B���-[�}�X��鋸 G.� >O��/��	<�'K֡Iuji�����V�v#�d{�'jrLs��P%���{>�2��ɘ2185���j:i���[ю-��q��ɰ�'Z���O�&T�bi� ���(�aL�,�B1qN>!�A#����O�Z����X��DjR%3�TA�(O|�E�)�Ỏy������ d$��{1h�"O��A�F@�5�^��VB$	0�ś�"O�!rc/Ï8R�y����&9?B��"O�5�ȕ-,���Ҳ[&��v"O\PR�,N(�BU�`�¼��F�'��� A���֌*�T�����/g�����"O��5���>:B�23�T6�^-RT"O�$�X�r�|�jwM˺Pw,��g"O�`��'�e���kɏ�@�u"OLXP㖦P�\�0�)@|fa��"O���"���h���L8bܵ*F"O�"��߈6�V,Pˁ�kT�l�"O��S�:s��:�/	&��a�"Oޙr�&C�dX`!P2�����("O��k�F��lHR��3.ۤQ��%h"Ot�n�� ��®ԉ}�@%�T%D��x��^�'��`�#��Y�$٘��.D�H�d+��H��f�Q����+��(D�H�1�P%(<]I�Q�I]��֎)D�0� �e�h	ck��P�W�"D������}e��u.P%(���D�$D��:�f *�T�C��
 ʲyp�D(D�<���9�� �v�̃1�9;c�"D�(��+Q�$aJ���G�8=\�����>D��gD�:I"L�HÄ��\�l=D�Ԣ��A�Eed�W@İ������<D�|b�ZIZޜ��B��r�� �*?D��J�S	l�Ee(U�z ��Q�?D��C�� (��q�f���D�y�c�;D�\8-�=a�z�RԄNlT1���9D��3�M�#o����	�e���F,7D�t�Wg�x�:�J+=?�d   7D�����	Ÿ́�R���L����Q�3D�;�dK,�}(���v�a�4D��K���?P���d)��cۯ'�!�$Q"p~�I&Q�
���֏�5�!��=�Q����q��M)ю��p�!�ӕ ���%ȭ+� |�0�Q�y!��b2<������~暅�!Չ@�!�$� d���j� O����HN�g�!򤟟\��1U&G�)���c��O�!�D��
W�Ġ�Ȉ�>���2���!�������0�^��Năc�5V�!��F�3�Ơ�x96բ��Տt�!�D1"����F�D�.~ 8SIݶG�!�D^<C�p)�#�"b�2�L�!�ϻ�����F+� T�t��=_!��B�E�IB"�2 �.�J��F!�$կ/i�23�Ҝ���)Jӛ1+!�D/C�p�Q���a��0u�P )|!��L:E���A$N4dѳ��<qg!�_�X՚�
mژ�����OT!�ܴg,�eqէ�b��8�@/B��!�DN�SX 
#ҝJ_\���O�<!��A>�2 ç�KO@��Z��ڒF!�_�4�>��Q�V�QM�p U�L�1�!�E
:a�d ��M`�����J�!��G�N��D&�'#/��Vn�!�DZ�Ky@|��/_�0����� �!���=R�U#�I�2��m�J�(�!�$A�j�ʜP���1�4�b�±b�!�$ވ|PIJ��M4l�̅�
��9�!�׎_�@��NّQj����f�n�!�d��}��i���
Qb����H�!�D��3�xLA�m�
[��u�0�!��!Fh0�T�76���1o��;o!�(6�j��1�H0tI�@�k!�5�>��Cg�(��a��͔9j!�č>��ez�A�|޽�6�-T!�� LԚԆ
c&:�k�)�x���"O���U=a�2ݘ$G��;V�"W"O���G�P�H�f�=utu[�"OR=!���k.4�`�E�3\�I"O<Ȩ� :-� �
U��YfT�4"Ob��B@MN��x���	A�]S�"O���#���44|�D��,Y��"O8��s]*�� _1�F�bэu�<�"M�S�J`��j�
ϼi�­Tq�<�F��jHbd�"C�j<�02T��k�<�!O�,)H��fgπ%d��7�S�<��ۖ?��A����R���1M�Q�<��/�BgJ�Xv��'d0��A�O�<ѓ���N�0���c�xe���ԮMK�<Q�J�0$x�*�l�>P����B��C�<1D�0�j�Co?2%��+2k�W�<y�E I�AJ���N�qh�~�<�5�=��-Ӈ�[�i��Y1��_�<�E.�������IR%b��E�Ld�<i��ЪW��pcR�md�����]�<a3@�8P�%�U�G��p@D�\�<QT��$[��i&�� �\yx���\�<90B��?��q�pۄw\�S��V�<ip/�.���2�l[�;�uc��N�<Iw,��*��U&ٶ"�X�i���Q�<y��+G��ݒ��V
���bPL�<Y��Қj��Q �G�[�.uN�<�b"�'NB�([�"'������I�<�פY˘�a�"�?pE�T��C�<a$��8J����%�����G��j�<�s/��}��˶�	�\1NL�W�
h�<)u��pANx��>])��bjXe�<�f�=	z��7�#6��9�gAa�<�� �)j��Q����9����n�B�I;N��0�A�ȔX����u�B�I�wͶ��vI� r������B�ɐI�e�!R� ,d�	�d��OGB�!ܒ�d472}e��I�B��%x�a
7*g� �����j��C�	u�$�A��(�ȋFN /P@�C�I2$��8��np�����{�B���'�p���JY�_Et�H�ǚppb��'<��R�w��(�6�W�{fv���'/�(�� 
H����M�x,R!��'��h��'ܾ1|�;f��o�d:
�'P"��@B��
k��0�M�_!N�P
�'�De�%D	���@�	!i�RDa�'=�la�݃\<tɢ�����8�'O���v�L;�"�P��\ ^�i��'
�X���O�4u�mK�@[�OtV�C�'@�RV9��h���<�0
�'������5����?0���	�'?�@s�� W�Я��556�a�'���kr��5^�|�ʀ�H�8#�ty�'æ��0j[�Q�lP \�^"	�'��P��i1n�8�w��r}�X	�'m�`q�l�+}o P'�55�u
�'Z��s��!(`�uO\�H!$�#
�'U��0� =~���ǆ)9Ȳa��'� � ��
�6M��"�N�#�(�'��J��R ~�h�ϼM��[�'V$�e�̤ou�9ٖ.Y�qh=J�'���A�`ٰ1β ����
b)K
�'r޸�"ǅ�.��`�v�¦7��#
��� �k�mT&G*���fӨ
�����"O����IQ O��iP�Kʶ#1��ۡ"ON�����?�P8��^�&��"Od��'L�X7:�Պ��9(���"OH(J�%��@Ԋ%C�iPc$��)�"O�t��)�|~$]{TI�8v8�"O!R���>�r��EOV��Y�"OX�1sJԟb�CS$��#��8�$"O|qjW/=��m�RD��r�c�"O���5M�pb&���͛	j	���"O�L�E���g8�	�S,X�]�<��"Or@��h��2ز\R�l�T��"O��YF�
I��4�=uѠu��"O���V��&�H�6��.@�@�"O���7�_�#\`ÓH�7w��"O�$IU>ܜ��������`"O����e��X祟�=M�e�B"O���a�J������=L(�3"O&����;�ޙ���ߑ*N��s"O�eA��*J<bQ.�[ z\�$"O����N�li� Q`f��u����0"Ov��.�Q����R�=w��
`"OV !r�6oX�E�TCV4&V���"O�d�5�F�6��4zQ�Q�MD�d��"O����h��RD��X�6"O�܋G�ĺ��)��nޟT<~�h�"O����hإI�p�PwNѦyS�=��"Oz��_�p����iE�yQ�"O 8���Z;~l0U�2��C`"OabD�\�w�1���^@���v"O~���U1!ҕ!���A�<5�"OLpJfj��\�`t����'{����"Od�i��V��r��W(f���1�"OB\���M�7��S.�tXP�BV"OZ(���#7��J7dH���@Ib"O�� `��$`��l �9��C�"O.���I:Sk�Ѫ�a�%AL��#"O�\��@0m���!1��a/L��"Op�jD���!	������`�"OF�kqg
�D�6��/�ebX�T"O���
C=2� �)n֭U ��C"O�A�0/�� Y6��>FH�a04"O��b4s�>e0���'?B�
�"OZ�:��V�A�l����u �4�1"OF�9��ٱ4��(��W}����"O��3�� ���gE�[�x8b�"Oi�q%O��0�c&��D�5"On���!׾�*����	2�έ �"OD�����P���ZĪ6&�x��w"O�ɺeo�9Bh�T��i��C����"O8�B�_�Z���)�-~�}�d"O�!��,�%x��y��]�is�� "O>u���~A
SHڡP���#B"O�H�E�)q�Ԑ$��&���"O.�G��E'�9Q�*䌔�0"O�,�@i�=8��1@JĸJ� �&"O�(��U ^�3Ǫ5����"O(���<&~X��f�Qp�|�5"Oh!b�)	:C�<�{$J�XN��
�'x&}�B�[�:(�X;w�ƈ��'�Z���̖QA��ǈ��}���S	�'p�ѮΑ;$@R`Cs�ހ��'s�a	 "
'C�r)�0�6q��#�'�ٶ+̦Lp.18�'��n߈ "��� ���A�S�4UvO�o���J"ON|Y7gM)1|�u#r�X�y�`@�4"Op<��D�5G0Q��ޯ%��!b�"O^8Je:"zH��/Ѥ��%[A"Ot����@�NBb�(ə3쨓S"O�	��,�X�	��Ɛ�FI��"O�	�԰� �c�IAdZH��"O*I���ڊ{����GɃ�o~q���'��L6}���$dM�%��y�a��B�^sC� aB���D�O\:m9q��A�N	#è�� ٨x2��; L]9��Q�J�8OyB1�$�"4�Q�h��lR1$�(�xR�0��~�&!8�.�mX^`)���D	W��IH�ŉ�qO"��' d9�%>�1GCY�LE¬	���2o�U�O��d�O��(�O
]Z'g�<Q/��k	��([�ّM�d���`��3��f(,�`F80������ �@m���D��6'�Mc����w	H�a�C�Q���Ć�	�Ё�{r�' L�83��*��8� $XbL��f����iP�J73;
��V��1l%���L]��(O\� oǬ HJ���cù[C�0�QJY�tt�'�'���!sΕ�IN�ko��K30�X�{b�ߥ�?�c�i.�>��v�
/�
!!�_��$g��d"�OB��a"K/^� [��&$$�a��O��n ��Or]mZ�M�۴��Y��(���g�<F�Q�@tӶ(��g ئ��ICy2_>�%�̉��H�G-�Њd�A31:�y�7h�XyL�dJ>x��6mK���m;��Ȋr��p�Ο���w����*	WL<i2�A�D؊�4��Ƀ���kgЍ	�ʐo�zR�땸 �J��W�<�\c�@�{#�Ɔp�d8r��~�b�4tmD����M+�W��I$��ـ���)�汚̇�m�N�⶟���k�'��O� ��������L�	!	&D���ɦ�M�i��'�����bh�B��>0�I�ՠ�h�08D#�FyB�W�n*�7- ,O����jĘO ^mF�Z�%{��R�఺� � m��=�FfW�uh(�h&�Ob���v�@�M>�qO:G�H/S$���Ț��hT���ӹb����e���]ӏ�~:��
�1�*�7J�<ACh�q��S��R��ԜHeD}�:�?��i*B"=��O��I
��oǘ���JE-v{�A��>��d&�I�  F�ڗfQ1��x�4�P��Hh����즱�i>��~��6��T�M�H��P�2��x-���ʞ&O��y"�',BLj��^2{��A��W�'<\�pg�V�>��͑#v��u2�&ϕ7(u`�κ�(OH���U8E�V�+A�\�64���QcN�3��ǎH��k��,'\88�gL:N�TX��{bF��?i��_�=,��s�=u�  ��VP��D���f����d��.XL��,W�� �
]8�!�Ė0���`\�qV0uأoٝ����q:�4��΀	��(oZ�\$>ѳ�`� hI��E�G	o�����8�����K�җ3����i��0��(\�E�P��	}��� %�Si2P��Y��RDy�
�J�!�A eI��铁�(�R���nщ:�X���J�/j�� �i[�X��T�C��fܓ{i�h�I�Ms����i��p�P�A	��xcf΋R����aa�Ob�Oh��I�|��֤a#���(b��`�N�-D����Z��=�ش�M{S`�i��G�Gp��/I�7G�7��O��D�O��O�b����h   ��     �    �  �*  |4  �>  \F  P  QV  �\  %c  gi  �o  �u  0|  r�  ��  ��  ;�  ~�  ¡  �  H�  ��  ͺ  P�  ��  ��  9�  ��  �  `�  ��  ��  �  u � �  Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�� |d��"O
`�(�;���8���-0��1%"Oj4��ND^[��"3/9�0|H�"OB���H��*�ʞRy=a"O�味V�!X��!&F�:J�$���"O,��a
���C�Ą�M�"O,$3%o�-���p���+Ն�:1"O��ݢ1����`���y14]2��i�<�6��{_���c�H�`�fX�$Kn�<��A̼VI�xR[�)�Ć�pඤ�ȓA5��('nߡ4�� �)˩%� ���,��r�؊b#`T�eT09���ȓ!�b��g��}�8�F��-? �ȓ
K|m�ș�VṔ���2�%�ȓ"R�X�j�4JN�1�˘X�i����̹	_�jZ��1!g��zܶ��ȓgil,*�J�
j�Ne��i�J%b���f	�(U��:���G��$Y^م�~r�� S�%T"���k\�jx�ȓ|4�1�îJb��@ӵ�ݩn�V��/[`�"�v4�R�!ʎ<��M�ȓ`:��z�ؚh�J�Z��$HY:	��H��p�m�C1��!��B:��0��EnjZA V;9����J[
2���	��4'J�EA�IVW&��~�(aZ��ӹ�>� o�Y�|�ȓ�f�A�
Ο7�H��M�$�����mޠP����/���ANXo*�ȓTv�����{ ��-7�*h��I��sB�8�8���3����ȓNe*M�悡;������X�o��!�ȓ'lj�#F�m�+R&;�|��2)n�C��0S4���T:
b���:�0!��e֊��)��ͷV��,�ȓ0�&�8#���� ع�L�����;�P�AFd���,w�6d��r�EQ�( �gVlɦ�M,H��,DP���|�I	$G#\���ȓ"�)���E�B	yt&B�^�LɅ�	�<I������t��v��AHZ�<��#I�JF����3Q��j쓣hO�O�D�4�ˇE��	qo���'b�1��h�.eq��p�J�N\�xR��D'O��ZSb
+h��D��	2���["O�L��!A)����TP�"O���D)ƸzM��1��0&�l����'��d��1@�l��bL
�4���ί'�!��xj�9v�Ҳx��Y�A�ˋd!��T�`�g�p�,pS��*D�!�$�5��U���Ϻq�<yD�W>P��4�S��M��耵��)*�� ~j� ���D�<���y��ebP��$H&�c�C�<I�GK:�1��2D��!�FG�<q���{U���� �u��6/�$�O���MwL�`u!WA�(�����ck��nӖ%Z�$��vB�K��#8��86"O�y�@�I#%(d�獊!S����'�Q��p� �~�P$�G�>O�N�i��)D����+R�B���t�>�Ӊ,D�L�5�_�\�<A��<�8�K,D���s+�Z��	�pꅐ%\���%~ӪC�		B*�RQ�Y�9X6PG �O��˓�hOQ>� X � H��h��@���ԼU�����"O&���"Gep��'	�X�}���'�'T�)��xB�P\���҂t��E*�OC�y��&��r�̸r0����V���/�O
��ȦO��`�͎�I�.t #�'1��6}2�S�F�A"���p �SWa
�(O�����;]�E{�ݰ-_��w	Z��"c�HF{J|*���#1�� ��19I.\�a�<1��J7�ht�e$����ؓ�E�^?9�y�k/�g}�M��D�Hq�S:J�b��Պ��y"�_�|�f��'�G���s�ED��y2�4t�T���N�j�6處��y�����`�iŕ^N���Q!���0>�@G���Iʱ>(�=c�a]mx�Ex҇Ų�z���iH�v�"��Ӓ���9�O�<8������
;�d���:O �<���^�{��(���غ'���b����.A&B��9^��A�����Y� �7cCT�$�O���ԟNb?��k�CG�yꢬL7n^fHy�F�^�<ɦ�#1�ahĎS�^Z��@���MS!�8�$�O>�AB)j�,�s)�r���)R�J@���3F)Je9{:�MIu��'_ozlBҨ�u�<�O��@D�9	�m�#'v���j}��	Q~>iJ��'gq�p���T\��qIɞ t稥��	M�D�*w�^�&h�|���  �!�� 	�&AHC�����F/�j�x2O1�s.(��NY7SJ��a��ߐcP'�t��I6F���glݖL��m�1$ðph�O��L��G����49d�UH�A���y"��a��kQeSS�RH0�ڝ��<q��_ܓ`�h[��
`0^���o�� N*D�ȓr��e�@L�*�V�{IH��=�����c؞vG��������TA�@AK���=��{rE�@��is��:M.�� ��O�����d��,E
N���0B�B�T.ڰ�ȓz~L�r  �HE�̰����7�"9�ȓv"D�@�r!q��
%�ZJ��Wp�tzў������T�u��$°�wo���"O�%�cR&�R�fD#qb�"Ojڰ,��C��� ��F�TS�:�"O��c�"˥R�¸�$�K�b�����"O�Ԁ�fŽTϺM�"�[�����a"O*U�i:j5�ʊ�9p6T�"O A�-U>�M؄kB�QU,���"OD�R��5B�D
��̩Cs#"O�%���C�zd���80_���d"O�My@"�i���6
W&UN=0�"O�u��3%�x,�&/�IxA1�"ORAk��Ɣ#�l��N�vF��"Oz� �!�!O��8R�
�>)$��a"O��[�9B+��
�s"Pڒ"O�@g��g�XqG	��6"O؈!�@H`���D�M�L��"O��SBџ{/� ������`h�"O���0vBi"��\^h�h��"O��W	/5J0p"FI�Ra���5"O�t���޼&b*�I�EF)�n���"O�   � ��QK����C�� �"Oj���G/t�:a�@f�,�\ a"O ���Z?5ZQ�1�ɴv/��"O��ɶL�hp ��#���8b�"Op �f�ͤvh��ꡂػm���%"O��q*� L�n@Ѡ L����%"OtipSJ�u�����ɡ)�n��"O� �8H�lz.s�.Ԙs���hw"O�h�!
)k=����@�)�D%�&"Orh�GR�4�	($�>;��a:�"O�p�g]6'V��c+��x��e"O�4`��������	�h�"O��Ѥ�:b�,��
U�>����"O�8�I��[��jQ*�	d�d@`"OTr�S/jµ�u��8NpX,�q"O ��fֲkS.��,�e��e2"O(�3�-�a��} ��F����#�"O��y��tjUJ�	D`���7"O�eP7���J�l��.�A�=�"O(���aB.\���Bā�/�]($"OK���R�F�O�&.H�x!�D�?s2m0E間/Ah2�F��*e!�D �а9%]&2)��$˟a!�D˚[p����1`qŒ4�.�Ą�o'�h������5�A�Ik�I�ȓ\c(8r#��g�L=Q�hƵ	�l��y�8���8y������½y6�m����Eb�)ܚCa��P&NߓBZĆȓ&c�08c�+_$��8 R�\��ȓO�R��q�ЁXv��`�	�F}pA��}��A2���>?0V8�K�b��|��w-�,�Ң�0a�#ə;Aif5�ȓ Q@$�p�o��| ��42�R�ȓ'V�t�3g@�]����4:���
E��Y�f�bWn��+�Sv֜��k���j�ǚGN�\8o�5Ŵ�ȓ>x ���_�7�r��E���xkl4�ȓ>���c��0n��ћ!���i�ȓ8V�UAR��y
�Lq���ȓҔ$�Q�+<!:�(ץ��N2�t��d%��B����H��&́:0�8��H��F�8��N�:��h�ȓNN]����d�1��Y��8���|�D\�Q��2T���	�T�_��� y���!C��3�\G+L�������Gc�������m���Y�lIe��O�ء�M�.<f���ȓ!D�7 �m���NדKT\��ȓEl9�i�ni��z�e��	䎴آ��qg4�`r��y���ȓ`��p9�@��K�P���u�|݅ȓFc`����3Dj:�KԤ���=�ʓ}�͉G���F��Y
A�ϕFrB�I�P��PZD�G�&��u�î�\�lB�I�1����E�$Y�n=�i�B�c����lP�TS�!1��C�	�exL��ef�/v��ڰ���+�B�I�?j�@[�LY2R��
w��C�I�b��=h��\"�Dpf�gK�C�w�lY4�Ȼ:�T��3%Q�g�B�ɷD	HY���?un�a�eP.`N�C�ɥ8��$AQ��-*����C�$\B�	$5�f� ���<���4�FB�IM�%q2�@�2���
�DjB�	�|���a�'�M�%mR(B�ɾ������F9g��â�I�1T�C�	$;t�LAfU'&k�Q�v.��[��C�I�1Y6}�EbՃ�r,
AN�,U�XC䉿m$t���B�>)t��p6�B���Z�zm[�,�^d�eպ.��C䉿Ml�
��E�@������,'�rC�)� ���32(����T>@�a�"O^p�B� S�pqD�G�f=\iф"Oı31�Έ{��T8Gϗ7-p�!�"OJH`���$8&��� E�x�Q"O�\Ȃ@��d�����.k���7�'��')��'�'��'Y��';Z����#`)�Ä�/��Y�$�'�r�'��'��'"�'�B�'�:�	����-����Z��1��'�B�'B�'��'���'1r�'���K&�W	-���֌."L��Y��'��'���'��'�b�'0"�'{Z0B��Ih�][�i
 �f���'@��'���'�"�'~��'�R�'!���dU�[Q�	Y醿�*H���'9��'���'���'"r�'�R�'7D0�Gn$�	p��V����'��'�b�'���'*��'���'�~�"�/��,��#$5(H���'�B�'��'_"�'���'?"�'��2��
&+n� ��ɃkԾ01u�'�2�'E�'p2�'���'���'�>�#wHU'* x'BáV���!��'���'9��'J��'B�'�r�'���e�
2�b���J/8v�0H��')��'�2�'|��'���'|�''́
�OH!~u�S�_�.{��0��'���'���'��'72�'q2�'��Q¦ܥxdA�)ܬ2��'��'��'\b�'��#rӊ�D�O���"�rQ!�E�aР�2+[yR�'��)�3?���i<P�nۮ~�d ���;Q0L�Q��C���dKߦ��?��<y��i m���܎=�i�PM�(Q���p,p�R�$� J6�.?`n�����Fk>��L�� �`��凗\N����°��'O�Z��G�T#_:A���F�,0t�ĀH��i��0�yB�ɕ٦��
�*fMB,T�d@z�a��q�ٴ#ěF:OZ�Şa\l�޴�y�R�$۠�G�U%�n=���y�\L}��/��:�ў��ϟ�:�ڴ8�����Y&o�� on�H�'��'��6�Y�1Oz5÷�:]Y���ɋ�US���7�����G��5"۴�y"Q��
�X2��}�Wo�V��S�'?���
9/�y2��z�'$%�Xw�X�$.k6��I��N�.�q'+�IѰ˓���O?�	��B���+��n^0d�S��j��M��m�F~�a�n��"�2��D�/4�ޡ��RB l��)�M㓶i}�"�z{�Ɣ�\����p���L"��˗��h��8�6��wR���*�5RT�Z�a��B��ߤ ���}&�����
�m�G�!��Ƞ�b8D��!@#T�@��u�ff�3B�,�!� ?ZAyT��gu:l#`%�^ �Ѱ"�Qن��$�9jʌ���*���̀,�ҁ�3�ûF�H�t!I!a����#����F�D�Fˋ:(�b�"��ƱR�M��#N/}��0u$
���BOjD\�*U���&�rY��"YZ	L(��(6��v�'0r�'��D�>?i��]�v��� b��	;�>|�"%���������G��G�S�'v�@�N�2f�)8Tx�zӾl��������IΟ����?�O<��%P4 �K�4i�����L 9��y��iRY�6�'rɧ�R��ï�:��,�{�j��׬ʦN$�9o�����D"�oň���?����~$>9ff�{��1P�X��"�ß�'��b�VC����˟�S��n�y��JO:MXX�a�[�M��M��Չ�Y���I���I@�i����j����M�Q�,��:��i�L��Ţ��D�O��$�O���O�X9�����P� �@*%"�,D��`8��'���'�]�d��ҟ���++�
�۴��3Q۔�H� <]�`�(4����8�I̟��Iɟh�O3�nK�_�7�ߦ*LPɪf�Բ>v,�dL�i"�m֟���ڟ̕'���'jRǛbJV(��eh'EB`��]�%�+8�7m�O����O��$�O���I66��0'>���(�!zk|9Z3H�]4���I��M;����?1��f���{����	~��Aj����  �Ȉ4�bY0�i���'!�	71���O|z��2�F�0��� Lԍ/�����oJ,c2�'^��' R�81�'ɧ�I�B[`��$�,�|���F(�VX� I��;�MS�R?��	�?YH�O5�a�݈5o xxQ�G+����i6��'L��q�'<ɧ�O�y��_$�
����	^>:(��4G�@�S��i]��'D��OR���'���:+
���<'�l�g��)U�:0`�4�6����?A��챟H�$�O����+�5=�}9��O�:��������I�����{ޠ�k�4�?�)�6�����BG��OF����k^l��
��v�J�$�Oh���KH��OE��'��ٟ
uS���n�.@��kŀh�b]�ƹi��ɇ�/�t��?Y��?�M>��uH��� ��ܔ2&�ʯM��mZ��RK�ޟd�I������H�	֟��I@@��!䍍1�q�� �Rq`12�U����?1���?�)O���O�Ԣ0i�[��[�\(4A�I��G7�*���<9��?�)O��d<_'r�SwV$�[a�I;�h 0�b\�	26��O:�d=�	ǟ��	
:���8(����D|�� %��1 ��'� �IKy��'��\Y�[>��	�~��%ѝp+�ᐋJh۴ �ߴ��'�R�'^��y�i*q&��-(n|�`� ̭0䶔oZ��̗'ar�P�������?ט>��*D�W�gadZ�I��O��d�O�YR�`3�3�� �-1�!؆=�aЄiA$1���c�]����5}j<u����p�Iܟh�WyZwL�̱EC
�X���U[�LA�4�?	��ZJ��<)����z]�!��p�H�e�V��M�`�,�?!��?���.O�S&��JwH�3+F<�k&��%c�P۴d{HPsN>���埀Jweˁg�\lYE��N�~,� O���M���?����&5�Ǜx�OF��'5�uC���p��L��΄?l ��ChӀ�$�O���K�+�.�O���ޟ��<}�d�"�{�< �jM�>�l�ן�#p��Gy��~���%ÌL�J��I�5`��0a�(�B6��O��!F��O�d�O˓�8� ��7W�+ �Pm	.1���v��'���'��V�|�	ޟԈ2�Ya�"��CZ���R��G��=��Vy"K�0��8��C��r)�5����rˏ$s,@m��B�'Re8L�t`���5��.r�C��9f��b3���H��G�
}b�� ؃$��3Z��Fv����%P�7\z��c��Tta��$;@�S"�E���-��#%��A�r��</v�C��/�����S�y���J�0�"�R1�����q���9�����;qͶR�}�Hz�`�*Vd0��eֽ}2>@x�g�:tHY�����F�0�9��O�E��&����A��8;�@ ��O���*I{�H���@2l>���O�S_��@=\�╆D��ry�!�����(f�U�G��S�����_�4����4�� �d�.G�:h�-A�\�J������I�����s�S^V�U����5ަup��z��?�
ϓZL�|�uaxZt��r�ƿG������HO0��k��@�x�E��aCqq��ΦQ�I�(���#���������֟��iޡ��e?%aޕ��"��v$��#�EJ��WE:x��Ɇ2��x�SM�S��P����~ӎ�H>�q&@�n�L�>�O�舠�XLvtA��c��@�A�O�L�'/�}��S�����ݟ��ߗE=�[�ą�rd^�1c�|��hO�ӖI����+�O"��v���'3^�/���{Ӑ�O�yr�h��h���y���b�8������R�'IB�'I��� �Iʟz��Aޜ��e@��l�8l ���Hz�)+�/ĠHN�� ��6�ayrkS�A���c�&S�=�:������t8Eɀ&Ur)�Ю�E��x��)�K41C�kX4F �̳��F�"�
�ygA�ڟ�A�4.�6�'-��'{b�'��V>ݩ�	��zdl��E섗~������6���<�c �:(%��d�˜w������)��ss�k�����d	e�iG��'����'�0xM*���fO���9��'n��Hc��'��G�(�y"�|��*��V�I�z�V�J��p<ف�TDdU��(?��ɱ�41��`�}y\���K�d#l�񄞂YT��'^��ߦlR4IԻ90�h3�Ŭ{��=��?����'q��'�R�'�H��ȷIX�����$��P;�'D~6��R< ặ�:;���4�tc��lZiy�a_�1�.6��O���|�֫���?!��^��R�K5�L�)���8@���?���\�0Z��V�4��e���R��6]>�OuFԁg@Ă H`��V
�` 2�aJ��3&�[*#�����
��X���+q����V�jA�t̞�J�K�������Mk���?�*�i���� D#+Sx�j��4D���w�K�v��Ha��)uf�5/O$HGzb��w��� �m��3�v�I�,8�.7m�O��d�O^�DG����d�O���O�D�P͂��C�8*l��`��!(V��K'��JsJ!شv��lZ����f�^���[x;��"�Ru�\#����t�~�@#�i�q��'�<��UK�j���Qs�A�)Z%JF�3�A�)^��L>�����|w�!IP��DV9AA�EH�<��^mjR��g�+A�ظ3�.Jx~��0��|L>�k�m8$��C�I:�R�H�9j<��˷
��?��?!��n�.�O��D�O��مi��
Ѵ��tʓu=^( 7mL�
����h�N��_�c�P�3 [6a������n �xe���.w`��̕7I�&L���g�����嗫�(��@��$#Ӽ��j��mϐ������ܴ�?)(O��o�G�&�H��׺FZb�ʐC�)
�(�ȓr�#w���G����b\(N��=xI>9�aV�9���[�p�B��u'�'R� �Hj��S���lcs�و���'�ֵ���'�R9��|� j�0:�n�j`�T7��$0��2H�h������1#ȍ�|�&�?��
Zv{������� <1�'���zܐu�HZ �Tj�.���-�+u�BEc)/�I;A�����];�OxQ��mP���f�l�B3��f̓�?Qϓ$�6���B�dl|���X�_0���[<��DS�zB<���Dū{T��&�ޕ�y�R��q歕��M���?�+��DZ f�OFD�'��Sh(�:�$�
uդik#%�O.���?d!ʬ���6=�ԗ��i�|�s��- ���q���0���*c�y��(-@u���*@Z(�b�IZ���}z��ΚW4lڃ���H��Tx�䉰.R�/��Ɍ9�l"""P��~y���1|!�� �x�� �1�(P3h�*�V0��'�p"=�q�ǷNVx
2V�*�V�"f��V�v�'~�''p���@i���'5r�y'��)l�~z�G�tr ��gf�D��m�<9�(��1E�L�|&�l��h�Y4r�aL׵c?܁���A-�z��
P���GC1��>�J�@`(\�u)U��LP=j��l
�k<��i��|�)�3�ݠ}'h��T��/d��ڠN� !�!�D��^:8pa�*0~f�+ŊU�7�����HO�I&�$׺!Af@5�§J�ĵ�`�c�f��"N6���OH�d�OjD���?���
��l� I�-B�Ow�IPc�݂5�(���H�^����U�S5C��l.�~*�,P�I�?c�dE�_�jH+���q��(V�G�G>����J(U��Q�m�"YѮ�	O>A�m2�%�T#U� Ǧ�V�H/QU��I��Mk'�i�r[����w�=��%q�&��' �U���*��i�ȓ'^ꜻG�����|�`1?���<	%���?.Oz�xtl������?�c�À1[l\:G �aJ�:�.M!�?���m��H���?��O�����Pf�U�'�E�@!�v�&��(E�T�:��8 ś���.�sW,߆V��lA���K��G;.J�Y���h0��O2t%��� +�?.���� Bn�P��)D�Dh"(F�����<���8��`��w��v��)ZC�U��H�F�+Q�X&TV�'��2�xӪ�$�O<ʧK����P/:{���4%1Fl+vŖ���k���?�"Ɖ�T;,�2�ɝ)dC��V��S>(�bg���ʁ�E�$�����)6}�P�>&8]�Fa�73v�L�ꐃ��O��!%�.H�1C�eM$�:eJ�j�"�O|�d�O���=�C0uq�d��r���H۝G��b����[yB*�,�O,h�#K�]CT�EĲ�jV"��|jfV�Ds�m'?�֩˱d��pTH ����X�m����'���'��Ae�2�'^r��yGÂ~޽�E�D��	WȚ='P�pѣ�f:bD�B�aRQ���yrF^;N	z\��ҫv�lHڠ&%��	�P��D�>?
�0���L>�0�G
h�pqCW.��
�����nD��-�<�4�ԟ`��r���?A��D՘�IB���R\�`�[LH���'-L��&XP�M�c���WA����'��>*O1��ʓ,��X�G��H��3	>({�lp��ăv�L<R���?���?������O�擯$c�={���.2H�d%[�zY2B3� 4�C�t��(�!�"c�Y`(̰+#�B���v�^�	�%�%�F�	�D�aC`�O8����2Q
��)ըæ0��2�JO<O�C�I+i2,2�!~�t���O�z�y��3�ɨ��|��4�?��b����$�%#Tn�0uƗ�ߢ�@��?�i]��?i������>�?aM>at���{�8��!%@�A�vA k8����<��6]��9yT���2`޴*!��1$bh��Q���$�d
�bc����ڂ?W�1��BUD�!�dɲ1)dA�u�Z-D[^��E��8@�!��ͦ�qԊ��	r���a�S&5�<!�	�L5N,ݴ�?�����i�&��dF�ew�1Q�
F�:5ȷo�0E�r�D�O@hА�]�J�:�Re�J%W�T>ɕO�j��#��m�A�#q�,�2M��!Ǐ�q���NZ�`o?Q{��^�:���@�-ޯ
��-P�.}�[��?A7�|��do��4����(�:S����^��yrm����X0M�;��%����,�0<��鉨.N�xv���#��$�P��fgj���4�?���?�C�;O��X��?I��?�;Vuc�ްRq�QI�N6s ^�g�F�"�.j	�\k�g�t���P��c�.�z�X����pt�S�8��	"�R��T��|Bi�4��8Q�ġw����4�X�'{d�O���t�����5�x�	toT�PE@��GD;D������,��:0m��;A*��#<?��)�'O�`Lj�-�feB�h �u����Q�z���j���?����?I������O�瓉p� !���0c뢈��隘WS嘷�}��2W����=yRi�q�����,Zv�d���cNqH��lZ�>YД�'��qhHq����� ��W��a�h�!�?��'�x�RE.$rlY"�a��p"�=��'DRY��C߾#�F% �&��d�
hK�yr�3��:�@��O��� �<_��P�-m��!�d,�G���$�O
���m�O��g>�1�_�b�:���\�s�~�0c �.�j��+�$�i�,� X��(p��d\�|V���֯@�B8�d����!�0���-��^B�<{w�O�
|r���F�'*���om�FO�>QF��1;-b��7Ɔ:9�����M̓��=���O7V�6��e�i�P��k�E<IS�� zuk��ު0	�@`�]5l:�@� 1OB�O�N���i�"�'��S�*L>�������g��6��PiC�!���	Ɵ(kSO���4�቉���T>��OB��I&B�
S�a	P/�<4���O���&RX�x�F(D
��Ĩ���h6�$>a.�$YZ��ި\��H�攎W��R1�`�ɜ��S�'9�����[��� W����v���<����wb��6������*x�8����HO�l2b���)L�kbbD�u�j5򴋏�Q�Iß��	�'��aA�����ПP�i�� ��W�"È�Q��4E�q;0my��S��?)���@=���|&��i`�K�HO�51t�����IL�5�.Ѐ7�ֈp'ƨᱭ�y��>A�M�J7BZ.��<P�g��r���6)��q����)�3��H����4s\$�{�NK'!�Qq�1b ҷ$%@P�"��%5����HO�)$�$ .2
-
�B[g2����f� ��ד>3*��O����O )�;�?�����tLZ�_[P���ьg���� ���w���z%cŢ:h^�	���?�(xsD/	�m[��Gy�aE"m���1*�iPI��W���QfF��wO�8�q�Č1��.�_�Ey� azA�2��s��@����2��B�a���͑�C�\��X�^��y�KF�8
a�lT�_H8�ړ+Ƀʘ'��c�8�5�/�M���?tn@&��Z��J�V����V����?���[�2��?ٜO��1�����C�8�U"Ǳ{��v�X�2���@M�5Ep&����p<�ą@-q��A����/�mY���
��1����,�jJ�M�vj8�D����F�"�|rȑ>5�H)�%��M*D�S�4�yҍ�90����i��E<P2�Z��x"bw�xq�-�;f\����W�,F \�6�G\V�Xm����	v����,O����
DԱ�1�Ӗ,�0eRq�<B�'2��HٴhO�&�̔O&�S.#6Zh1C/"��w�ߝ+���'����(H�?�q��K-�����'r (u�!�S1i��BP�(�E=}�Q��?)���O
�O)&��bD�.�l|��JC�c�^��yr�'�ў$�'�:}(�b�`̤eR�nI��ɉ�k���z�ؓO�#���?oTxk���$��ڇ�������\��>�1����@�	����i��𐤑�O#`�9%]B7���ڕ��aXN��P��N�g�I�3ԝ9��Q(�@HBߨw�^�z�G�W��5��@ *��z�!'���/��%@!8Q��*	� ���y��	��?�}&����kS�*#���x����m[��y��,<�@ؘJԴE�AB�l�1���KW����,jRe�|c����H�H��y�J1:J&�#�f�ON�D�O���Ϻ����?�O�6� Ӈʃ]��i�b��lۢ	���K> }t����5�z�q���K8��2���C#��U�ԏi]�4�S���J7��I��E��ń�w�x«݀`�j$b%ə��4���CϴLl�+��U�a������R�M�� "��R�y��H�b������T��%eL8ǘ'�c���F�J�M���?��߰ �̉0���1�.p���?��-��B��?y�O�9���'�n {!+7P�Ab�%K,,�$�J����#tD	}8�0�sj���l��+܊��X�B��6��j$��2��j�B6���U� -�/0�d�qzt�k�͜m%�H��~�!�S.؝�MȱV���%�N�s�!�D�Ѧ��*F ސ��$�&T��D���3扗*S`\��4�?�����E�0�����ϸ���"}K��#ޕe:���O�=�tA�p"�c��g~BD�#2I�_(�\��$�����/<6ԑ����_�+]zLnE*!A��Cwd��()�WF��ɟ��S��*���cr��;ziPu�j��]�ȓ)��]��)��3�e�L�&�T��ɛ�HO�=(G��v���xF@����1rŘæ�������	'��S�+�ɟ����i�i #��Hr�\��ᒨ6�] Q���rx�Q��F�g�	�-h�d�2�hpF04��[I>Q��)4��>�O�dYV��.j: ���H�5�6�Ȃ�V�7�>���|���=Sp� ��էp]��F'X>�y2l-t	e��̯s14�+��ˢ���Of����ԑ�^;n�X����),���� �	.Y���i�O,�$�O�����{���?	�Okz�0a��xl��C#�4|�d���B�,�����U0� ��/�� 2�ɋ;P�T4��i���8�m�w���&�Qb0M����6�02�i�z	�D{"c�m2��S�S�V�Mb�e_��"����L�6�o�T�d�<����'��$kD�'�� Y�
�l�dĊ�''2M���ؘ>Z�`��
�CLy�y��>�J>���� �0�t&�6#� �y�JȲg�%�"OH)�S/��|Ca�e*V33�R���"O��cU�������zIx��"O�h*Տ��0�t�Sb�1+�r,�4"O9
g'բv�ZH���3�zmz�"OACsl�=S ����Q|P�x�R"Od-Qb��S�~��-S�VJ��Z`"O��a�0|+�CĶ,A��X1"O@\�/��%�r#� c9��h5"O>)�1��JJ��t$�L.�)"OP�#���,X͎���h��"O�+L�AӼ���f��\�rP��"O�m��9X�E�ƅ˞8�V���"O�E@e�܆&g`��ƚ/u�@ĺ�"O@`��E����$�׊MDFѫV"O��1�A�H@ #W�V0 ��"Ot��g��_��;�bT�8#���R"O|��r���~��E��OЖ	;g"O��#'W)u�a8��KX�����"OL�Z�K�n���Z���M��!r
�'�4��@@.]2*l0#�	;��|8�'�0Ȫ����|��=Iֆ�'8g\�
�'�Z�
���JcH�`⦇�/e$���'hB���Y�G���K"�E-(�};�'�Z�;�l
&>$�̪A !��hI�'f`�F��� ���U%0���a�'��� l[!,�� ��  &�`�'����w��A|>�C��"^�d�
�'A�<��j�>���z��� %!@J�'�ˢ/0<�@�Ja%W��(��
�'~�ТÈ�Xm2���ċ��y�	�'�Z���m�$�̬0���v����s��c �͉u���h�4$@ԩ`R)���4���8KA���ȓ�&�+2�_	<�Y0
�8����<Y4
�x
���e��b��|���ٓO�%���OW�j�R�Hj�<!Ө��DY�3���H�*}J���r���H��z���I�$#|�'vj��B �G4y9#�NG-�C�'����'JA�<����|��@۱M� p�L߃Y� ���	�L2�zOhؔ�`!��/���,J�P����7A�e���g=<!�֬z�0	�S��6��q��+�U�O� �Z6��35�0��<Y2��uI0����B�Z�|����fx�Y�$��������H�<1 �~3����*?�(uy�DS?M� �	���0{	^���d�hD��O���O�z:�  �$�k����"O�MYR#P��ek����.+h�£"ʴe���d�L�VJ8��דt�aЬϥR~u1���~M�����%i?�Z�S�f`z��C�{N�aǟT�����.YnB�I��PE��jR��0�r�V�9�b�0�v�F�y����E�x/Q>9���V���1v�@��l��+)D��� ��8��D
 ��P�7lܝL`��a�`]��$ΐ�(��	�~�j\�	�>,?��D;��B�I	e��lqť�fH\Kwƙ2)����6�jXc��'�x�`3�F$~xA�2��7��x	�9վ��#Σ���
#���1�b��
�F� ��2}bn�U���(HE��A���7���u��Qxf���$^S �r��3�?�Hi��'��X�E �$�J@pE�����Ň?�HK���,T�1�A�N �|��C�T�'�R9����<ͻS�8���*R�^���!�"t?�l�ȓM���0ԏ7�̼�2'B��U'���6/R������0��Ԁ�S������t���������ON|q�j�#�Mˣ��7ud7���� hbL�%z@�ґ)Y]i�)�+��y�D
]��ӑ��"1џ ����M',+��k�T�h�o�>9e�H�g'�Y��T�=���B\�4��?˓�n��m���t���a$� ��˭@���d݂J�>�����
r &�]!K��,� �<8	�',�[�O��	� ������ �����]�n��| �A�T��*E�'%� G%	/T92��E�s��<ۤ*��9�L`��J�ckZU9�.���[a
;}�&Γ*⹗'L��1�5'�Q+��M@��ѻ���Ȭ1P�8+�J����1��f~�̋�Ib:�sA��+���*p�W!���� �>�Q�H����?ɃzP�8����m_i�R%�`}�bՉO�m��@�j��C��*��~n�*�p��?�h�ɖ�t|�;�jQ}��8����
�v�x7*�+ �,�8 b��jIzȣcǭ������=a�OzMK' Y7Q����6�Y* �m�E�'�O(���FP�2�ᨒ��&̪�R�L'H�!)S�	�j���۠�I� ފ�� �d���f����a��	���CE���OR���ҧ�&]Z�f.U��1E-U3e,
�d�#�=�,�Y�5O��˟�'�̕���^x(x�(�`{���VB�7)Pl����ke���g%��WhV���!��*TWJ��"�-���>2mD�8 ��@v��rnV�S �����Z+�~��@�b�P�2�G|�'���2C��,K��S$�r�.!9` 1��ߒ$:<��d�  �V	�׈(!I������afe��MX��u�����Ӗ���򁒛	�:M#P�'�6ܡ5iT�/�\L)�m
�bs�R��DR�N)(Q�@��9"����'Ǆ�A�!��<QT��r 0e�/OґSH�;��P/֡�(��o�H}I��X��aEDQ$_�Ą( @��8Qt����-6��D�AT���¢-�iäY�m�!P'�x�D�
lZ2,�2�'[ q�����OTEA���
bZ�j����$�A�F]d�̬"�m�VX,}3�E/�TDC��4ړ[
� ��S8p�"5K��B�*J��J��'4�%�T��$o��8VHJ�+ER7�dL�0MX�-!�D}���� s�C�4OS�$���u��MyՏ5{�@�3O����j»^�(����tY���� a�ي#���+н��A &l�Ov�C�;S��\�b#�,�iB�x��1Bĩ���f��6.F5���-;`��+3iT�J0t=2S�x5Pݱ�ŌRS�ĪO�Oe��/Q1S�������+;&���A�;|11ᐈ]����O� t�&D�u����hL�H�Mk��[?�R�Ȁ>� u�"
4ړ;�PEH���-���K"ćFx6h����M�Q>�	�t�� �5<���"��M�$�;F+E,phQA���7�l�!a��b�1UCD�]�V0�lд904`f��S�D�1��*F���2V�FL̕�e�'����&
�P�yb
�g������E�TnZ��]T�:���&�4��v�nL	�=
�pJE��3��t}�C
J���z4�I���$aq�̊kO��$a���4Ń¯>y�fHIS�d�!�P����Wn�UyJ?7�P
���`rH?�6b�G�'T�B��/�OJ�Z�)ŵW�]
cҍD}:��ĊR]y!��Ey��HB�,OnE"P��I2�;t�`���Y�F�;��1�Ov<X�lʇ�F�SB�=~!�����!I�yJ�g�<��O��>��H,�(OV�B#��
S��Q��SQǖ��1�	:I�U�v��J�dUʦ��fɟ�삇�F�xx9��.���O.��v����OD R�Ųc^�UȂAL1�DmZ�^��ƤR6L�ȦO\-����ƺ�3.���H��pF�L@�af�c`��l˲��֏�!P���$�<��	?�~�,.?�o��x1��!$�H�G�R4aȀ���V4D�(�  ���,�@�_!{s��AI0�Z�v��ɋ{�����
&#Vj��q?�vG���y��~ ��O��@h���6)!qO��b�a�t�g�I�u���x��C�w' �����,\.C��8�>�z0H�k�����љ������ӏG���ߛq�< ���T�exl(P���<���D���'e���a��8w!���W �t^���'�x��7F�3x+��pn��j�U��'F��yT!ٍ4�����.\?6� �'��M�c Z�s��j�(O��ms
�'H���܀uN�mڃ/=M���b
�'�H�
nM�m^ ��I�Bvr9
�'��LȓB\�%��4*Pkʇ>���	�'؞��e�s��@ף��7�����'3�$C�Gݯb���Fk�0��<R	�'ޜ8���:\��)
�(8"pJ	�'jP@�%�	N�
�B!L:����'��i�A�Ϸ\�&���\7Ep�H�'�i7��.[���A��6;���'D ��Z� �=B��Ef��k�'���x'�
A�ƥxe�F0��1��� �$z�
X

'�!�R�Tj�ب "O �!��T�9�����߈�x�%"O؈���%t���0��R�0��	��"O.�P欈�w�2�)C��"2��PD"OL+�eӘ))�p��Ȫ�V,��"O� �C��9E��{����Z~Ѷ"O| # � BNh RM�vh��Jr"O�t�#=9@�-�M%A�Iѵ"Ol%�%(� D���wQ�@�(9�"O��A��Y�:N��� ~:��"Ob �P�E7����oE� lYK�"O�3��U*X��
�cV�t��\2C"O"�9������gy�µ"OR�ò.��&N��遍Cv69�"O��K��
-s��:�g \Wv��"O�@�	M�DaH�a��P�u�v"O��1��L"b���C EaF>l��"O��u�մwQx�AAd�7"��U"O\�;7O���b	� B�7m P�"OV�j�	uT8���A�g\`z�"O�ݢ��^�.�F!F9CE��I�"O��ꖋ��.#����s1@A�E"Oy��F�$s`��&��+ &���"OM���byI6	�rD��"O�M
����qЦ��1jŎ��Ċ�"O�Q�H�=�L)Ci�c�6�3"OHm	�E�?1��)��59���d"O8lkA� 	�X-z`��'GMBU�"OL�Y����8`���6.h"�"O�%����wj��;�ʈ,Bz�"O>���&��8��P*?��{�"Oja�`�̍O��bUO	;V���"O�08�MH���;��)f|���"O>��cʿW��(ȴ�-5h��p�"O��Q����R��Q�AlSc\ة�"O,� ,��@L�<YN2R0"O(�'�U����z�(�4��90"O��ˑ	��.e��1�N3;��La�"O�X{A�@�/�u� F5G��P"O�5��0&���Q��,9����e"O� ��+�:X��`�2�?@ʈB�"O���$�^E;`!���=,  �"O���TA�t^�8��J�R%+"O�|��Aβ	G�=:`�.<�[�"Oz�#����hs�� ���K	z)��"O�`����y�U"!ԁ)\}�d"O:	�VF@�	��T��o�Lx>�	t"OX�ؖeӏ>�e�	9}e���`"O��
���*m't�
�.B�IXp=�%"O�L��M�
�hT��,D�+��x��"O*,�S�N�J��j���
!����y"�:>��4�-&��rDA�y�M����t��7Gۃ���y�(��M��&�:*;J%�#����yB/�u�ڕ±�
	%�|�;L��y҃��p	�f���	���DT��yŕp�n��"����ũ��<�yҤ�H�Ɋ������]=�y"��n!
Ԫޮ3|���+R��yr�Ϲ+�8b�ɥ|��q�����y��I�d@}T&i��<�y"W�4f��c0��L�l8J0擴�y��9-Ă� ��:A��	���0�y���@�a*ݮf��9 jЕ�y
� tm����?�(�Ǯ��=��L"�"O���!<YO2�rP/؎4zB���"OҭgG�?� ^�~���y%"OFp��`2d��Hx�m�X���)�"O���2i)C�^js뉼C�R�؂"OD4��,pn�r *���\h�"O*ݻf.��r3�U�+L�7"�`�'"Or���5Z�֘	��K?g:~��"O�M��,�>��tB���X��#"O����D,.~p�#0EV��&"O��P�c��x@,hU�!e�\q�u"ON� Co�+_9��s Q0-�d�B�"O>�CF^�2qP �1M*he8 1V"O�Q�GH�7M��H �L�1�\�a"O�ձU,2��ÊD�$�"d�"OtU��Dιr@�$�C�-?|� �a"O4S��F�\[`UH�V!?Iԉ�""O��b�F��P!����)]?6}��"O�@�@�9�����O�O�M�7"On���/fx�����i�։��"On���܊o�Fj#�tlaF"OL����&C��ω�: J"O�Uq��߷^1U+ӎ�o��D��"O�	���L��h�V���w��tJ2"OKӓΆ�R�%7o/������yB��:�� ْeʄR�^,#�"7�y�-�;�����O�v@0�Ȅ��yR"] <Prq�cZ <��P0HW��y�%0����,Ө~� H�R��yRGJwލH�I��$�n���JD��yң��/�s$+զ��Jȏ��yү0-���!׀Ӫ8j����y"M�|���BB�yR0!qE*F��y"�ENmle��M[�q���d�U��y��G�e(�Q4}1�qcB��y�MMm�����L��v�����H��y�k͓KtL�Ab�'g2�}0%�ۜ�y
?-��{ŭHf}�I���̓�y���%K-h��j��U-���ި�y�D�*|��C��H�����V7�y2�A)(��:�NزMIGK�"�y��#J���0�����H��C�y���B*q2�f� Q:ƯP��y�(	�\����O8|��10�jѵ�yB�©%�^��ЅVor�$�1ʅ��y�*O�y;`a�G�Z�f08�R(B�	�
���@�$��5'��S����	0Q>�sj4J� â6LNHx�N�h�����\��v��7�rq���?n�|� O�pJ��W*����2��'�ؠ��"O�5b�hS�h�����
����B�"O��c��-@
��񏖆G�5*�"OX��V�Q�K�K���7��y""-WP�)��n�H�Vp���&�yB��oƚ�H�VT�ez�䐫�yr�@�X�@�w,ͯ8�,A&G��y�LT�S	��E�@/dɚ�!����>y�OR@
�,֦��u�T�.f���"OPI)ѬCt�UQ�� �:���Jd"O4a���~�� r����E�Љ�"O����E��\����t�9o�¨��If�O�2����64�mS"�^,R��(�'�r#Y�P�xx�t��*b5�AS�'Y�a!Q�vRDrD��kyX![��� ~}xwd��2��Q�#�V r��Y��"OB�҄�^n�
A@��1'!�Y0"O��
g��n����%��%;���B�"O�B�lȏH
��0c���c�� 8�"O�����{"Z��bkT�&"z���
O�7͜ 
�r��� ��_�h��]>���������8mX��r7��TV|܄�,�8	c�Q�h���Po�>2��E2bp9���T~��;�fޒ���ȓ�v����G�_���9��I#.¼4��<?��Q �[�
��!�_K����h��E�,��_�4Ac�W�Xּ��n,��c�5A����N;!�ȓ=.�yω/"4�j#)�� Ѭ��|ݾuc1.�&eb$	� ����ȓ!��	�6�%}s���-�i�di��=W���8���X��I��ȅ�8:�!��P�@��q�D��1K�%�x�<)����5���r�υ�X�IjPe���L�,�@�kߏo�L�K��Ib���&Dy��FIF[���	�(Dc�"O�I��A ��J����xk�"O$��!�(w�Tj���d.D�����ǀ��YZ@k͞B�l�B/D���)�R��Ԓ�G˭0$$M�
�Op���9��'Hl�rg鉉	�V;t�=���$yyB�i�B�0nB>$��%_'v@���'u���Т:c���!�ɽt�鑎�7}2ᓣD���'�è_N�	4H�?��C�	w����_�r�R��"e��M�'Y�����d� ���wX aK(<��,�!�D�!+����dFu��dô��y��O<�On��Dpp�y8�j{��HF�#ɡ���eN�У*Ço���إf�$�H��y��)�� �WFF)3�@�����0-�$&G!�L�b0��(��R�o�&��!P�/!�dF  @<J��5�$�"g�A
C�!��_�
�k�� _��0)ݤ#�L��%Oj�!��
1Q�ȁe޿+)��%"O:$Kᎁ�2�x0$Ң���T"O,D
��{���c�==� ݙB�O8��	�`��E��.��2<8J�F1D����Kg��3AA�q��E"D���J�G��+G��i o D�p�BL�<D����lW�X;��:W�#D�(6h�
�H�%�nz�i�'"D��Ñ�U�b���p�)�- -��?D�8YJ��h�e�߀w�BŸA�1D�<7ɞ����(�"#lacӊ1D����d"�:�1Z�P��8Q0D�x�@�%Ep�`�`�YlJ��B�/D�A�9��]��I7F����,D��aF�%��-� y�x�?D�`c��ˡ9s�)@H[�7��x��B2D�0򖩉%�t<GF�7�t�'d.D��W���6��Zd �pES-D���G&����a��$�n9�ш*D�32���r�����W��^`WF(D�, �)�5��x��&V�*�*cH*D���$�]Ք404�������+D����ܦ_X�Q�Ȓ5.�I�5�%D�(A��\;D���)sŊ}*'�#D�����L9"_�d(�A�51��c� D�(���\�N�Z�X� 
�>x�d��c3D�� Q��ɺ�L���?G�T]�"O��A5�� �zm���K-j���Q�"O� �O��2���g��8@�t�("O
�8t%L�3:�|��/X|�9�"O�f���������
_X�(�"O����P��w#f!E%Y9UJ!�Ń�6��p��A�D��G.+1!��2I�A�✥k�~qP�L!�Ռ,���)W�.r$ԉ�B�u!�M�X�1���ʝRc$����BR!�$%,���-ر
}69�����!��1Ī�1d΅^�<�Y�oE�Py�a�*^����qF��]-H��V���y��3N�a��.T�� �t�]��y򬕈Ygz|��΅ag�����W��y�D%2��2B�3&���	g� �y��ǒ,@��;�J1% �����ym��:��A�ǈ%Z \�h���y��W&v�^| U�)0δMBUH���y"ėS���3�@��ya@�i�%��y��	2�VJ�"-u��%h�#J��yRK^tI�i��U�j9���uj��y��+j��)I���i�6�"vdy��ȓE�"U��cv<����()Ƹ�ȓX��E�`ӧ)$��� �$��ȓWL�U0r��2`ў�7 N�3�^U�ȓy���(�M�3��钮W��A�ȓÌ�03H>7T�㈁)q�6y��f� P��Ȓ��y�$e�#P@����}8�I�cE9,��Rg+��Z�݅�@�r�ӓ�-ˮ�ǥ�;(�J��ȓs�x���O�'O�rq��4C�"��ȓ4�ʔR2	�K� z�
��u<0�ȓ��pބpy������. �ȓEY�`�u�V2%��ݲ$M�3�$Q�ȓQ�� �l�%0I��	خB�����s�e�ńB�>���&�u����3�t��W��-�X
��^�JI���
U1��Z+*�@��3��Z�4\�ȓ �q�@E�� �����'��d���ȓ(�r|�O�:p{��2�EW~
h���R�lKc'�.��ڦ�[��l�ȓ~�<q�H�L�n�;V(F�)�Ȩ��_

iJ#-#<P�ka��/1�N��ȓ, ��QI!�"t;��4D�X���@  �� ݘ��&�Q�+�F���J�$%(pD���Q��KP�"Y����2���!	�4u���O�nL��ȓ!����g���12 �v�G q>p���=#Z��G	J�+!h��D�i#݇�\y�ۅ.�\!b8
bF[Z�ȓj�rX1��AT���
ȁ� ��ȓw�����#<�u��Z8} 0�ȓIӠ���-�typu���W7u����u$�$T0��,�2 0|�ȸ�ȓG����4�Ȑe :���Σwy���ȓB0���bN*L�5!I*#����,���oM�6��ؐ	F#_X�}��9Jh��I�J���PS�FC�\��ȓ}�F$�GOM�a�"�����09Aд�ȓx��B@�[�.�������$�ȓ �`� �Ȟ'x�+F����	��y����]�03���x�$��{�Hx"2�Y,MS!`
�]��H��S�? �=c�ŐD��İ�,U�B� X��"O�݉"�bv�<@Ц�1T�r\��"O^�� ��>C�;�K�|���"O��K�#�����9�BP��"Oh�:�L?%�x�ےk��n�X�@�"O6,�'&�2�8詒��<�\m "Oؒ��V�>�;�酘�t0 �"O��@'B�q��hٕ7�4��"OjX�4OS�4�� q�CQY�8q"OPI�P�ǯH��]3�_�u=0�%"O�� ��FF����T�0f�"O
}���RaPF��WMʂr0��e"O�5S�`V2tϦe��,E�ri蘚�"O�)SvI�����N�TTR�w"O���sވ+����jRƬ��"O`�C�ʕ"Ay1u*�
[����"O�E�㮋�?dٓ�h�;3S��(e"O(��a#��W��9a ��~B��B�"O��PϨ*
 ,A!AB�v/d<Zf"O��!",�^������ ��"O��A$��\`0@��o�#)f���"OP��H�\��h ��Q�JGl�A"O��@�%� {��� �ya�mY;m?!�#h6U�s��9{.��bc�;�Py�o#i���@��4N0���K��yr��3m � �l��vh�!g�У�y���\ɒPgi��а6&>�y���.(+�h�i�`�A�y�ʾ̼0���k��U8�!_�y�{�����+4�,��S*���yr�V8.���f[�(46�b�I��y"
Կ���)&��-�xY��ݚ�y��&~1�u�v��-��y��y�?0��:ҪƆ���Sb���y��T�r��%�����%���y��6C��8@�֏�X8c���y��ަu�TlcE#Ոy����cR+�yB��
����sJƎl'`	�q(U��yҍZ<]����§jR�ɋ�ʇ�yB�WFX��+s��Aɔ�yRK�%"���&��y��s��y�(�O� �s����05x�)��y�l`h��$$gb���a���y2��.}9�m$�[�
a8����y�cQ�o��1s#N@��r��_��y�)	�=�X�ȓ�2���z��ڮ�y��GYb9[#l[[���Beܙ�y�ŔsB1��JN.G��1�AA�$�y��/���y��ƿ=�V]+����yң�l�@���ӛ0Кz��^�y��P�W��!gM�7
�`�-غ�y"a�,;
j�Xk\�-;N�h��@"�yr�*�e�3�N�����yRn�Qf�l01 �W��3P��(�yI:傉QBFI�N�m��CE�y����L�웴��S��p���yr��lLH�!����R�4���EG��yB����i�d�R����b'���y��L�\�K�@��h�~�IQ���y��"~����%�7Z/r$ Q  �y��U}���С;`��h @蕫�ybh��Ψ�:Jצ-��!*�*�.�yR��< ��e����!�4����=�yB$ܤ
��i��I.����%[?�y
� !���͎:T����V^��@K�"O)@.�5O��#��';�ۂ"O�	y�@��2�h�� S�2e"Ot}����T��aSj�"[�ޠم"O\a1 �aCV�t��I�T�"O�a(��@�	>�a�G}�@([�"O2X�1�|X��Riˣ*$ę"O�1�ɀ�f�1i�Yf��y�"O4!CaM* �t��Ƨ@�[;�Q@�"O
k�+�.��Y� �8x&~�"O�H��Б8wZx#"EL�Cp� ��"O� 2CN�l�����a�3n��2"OD0���KF�� ��j��Q�"O&-u�O��+u��[��� w"O�ur�$׬�<%�qA��+z@"0"O�
GF�g��0ȡ)��t�AE"O��!���l�������"hy�L1g"O�|��hS�#z�`1T!R���Xj�"O��ӗ�Z6>�����eT�_���p�"O@(�#��=�ȹ��e3rJ��"Ox�B�H;y�\���LJ� b�"O��W�_x��A���	�"Ot*�K��KȄ��C���"Ox%x�Gܐ{5��іn+H���"O��[׋R�� ��ĝ"�F��"OR9�&��6sU~1n6���9�"O�9c�Y;)� Ռ�j�$�8�"Ob�dc����A����r$��r�"OD�Z��^/�X�6S�
&�h�"O����j�2.��X�J�!��@��'�軤��$U/(�K���'n`E��'�f�#ïj���%+�N�ڸ��'�f�+�I]wJ(��$cE�9 
82�'@����T�M>QSt���>]v�X
�'��p���4�X��3h��.�0���'-P,⡡�g��Lb�o�:u�y��'���)6�W. }p�x`�U�5�dQ	�'�X9@P�d>�[�@�;g>T��'A�ibt��Ay�1�dd�8�6���'YZS�ǻ~�LQ"C�b�A�'�̌r ��!� 18�SS���'��q]����!��S���(�'L��V(��l��a��'{J���'׊\d�Q	MT[q(x�$��'��![T�ڀ�쥊'fμq��	�'�Bd2vjTwG������ w�H�	�'��,�p��NR��C&�T0u"���'�9�MF�[���x�GN/� �9�'�Z�Y2��t�%(��e�V��'�nu�ݝR{���Ḡ�^4����'AR�;�ɧ ����ك,T2A�'\�T�g�-K�8@&�:.�l��'�$i!эL�@�8����R7hİ�'@�%�o�B��W�K�^���'vd�EEN���%�� Z�(mQ�'wdI.4����a�U��	��I�7�y��?OuP���O���!Yt�4�ybjI	.��XRFK\�4�Á���y�Řti� ��C̵"�L@���ٚ�y2�5���0�'�$�������y���(.f���Ɲ([0���y�Nm�1jrb�mH�T���	��y�i��H\�U�Rm���:��4�
�y�(�tR<y�p"V���H\+�y
� �y�7� 1L�)��v�A��"O iZf$ľg��E*��^���3"O�5�Ulȥz�`�S��,_kj�k'"O���5'�:T8��*H�`�2 "O(�x�!�&� !�J �3�!�@"O* �׉Y�X�P�K�t@��"O�e�SHpֵ���X4�a�2"O�)��R����
d�H0Y����"O(����C�.$PV�ݼ�j�9�"O��[Ԉ�-jN]�d���wIDT�"ObQ9�K%
<D�CG�' ��"OZ�������[fQ&�c�"O�����R��%�4�T���"O����T3�V(�t�2��R"O�j�#�B�r�xQ�J�|Db�"O�L��@ʿl�[�n#��"O�\;�g�~C4�*WH�"g���4"O,�SՉA��p��!qDJ�"Ox��!S��D(��XqkȩrU"Oҡ���I�|���R �ij(	�"OZUA���-n��1A
�f�t�#"OJ��K̄)Z��"i�8C�Mȵ"O:`X�&0��PV0�88ò"Oq�@Ɍ
������$��x�"O�ĸcP�689���s���"Oz��T������D#r`Ma$"O:䐗�Z�j�\eS�)��Z�)�"OI��E�"��'"��Q�]2p"O��:��\�Tܛ�Ç>?�Z4�3"Oj�YeL�������5�\�a"O4�7��
k���PT��F�,1"O�)�!�I-��|{�Ý�V��QQ3"O\�Z� A�^H0���Ke$XcW"O(A��Ł�}4Y���I%P���"O@U)RM�li�E�A�;8�tbf"O�y�����x(6�
]I0"O*4�X�5 BHC���q�;�"O�ݐb%Ȼ~��Hz�O�eڂ�p�"O��y�	qx�/E�D���h̅�yR��y�ēy��C&��y2.��{�.$�cm��x��� Y	�yb�ŀ%}� ��	l��%��'��y�Iٷm*�d��b ���-G�y�Ja�j��m�#U� 9����yR��w{���:7��ZqIH��y�~�^��Kĉ~eЗ% �y/0���1��P�P���y��݈DJ��X�⃩Q���������y��.ߔ}��mG ���f��y�+�[���h2:לx�ph�?�y�!M=� �6��RT�X�V��� ����Ē�����2�P��,�ȓ[� x;W�C&F6��HH�xr9�ȓo�5h�� /}��9��D��,�ȓ2ft`�c01 ��QQ����j��l1q�ʑ\�2Hh��Bm]|�<ip��� h�@+u& i��&�z�<��m�r�Z�����]3PP9d�y�<Y�쏓wKl��
o,(�.�j�<p��q`�y࡜�JQ�'gh�<	�cGQ,���l��v=��� c�`�<�I�'R)Ek6�߆J��h��I`�<�Dʬx)X�j���r�x�R�Q�<A��ώ[�h	*�Ƣ��d�S�<� ��DV)�^!2e�
g9r��"O��!� ��0��T�i�$��"O��WjK��d��`X<8���"O�!J��[+Lʰu���R�
z��)�"O:���jۈh�V�
HP���"O���v�V��*1j���=G*^i9�"O�����)\e��)7.������"O��r�i��5W�|p�V�F�L��"O��P7�Y�N5���ƅ�8��8�"O>��3O��=N�0�f�U�zAR�"O�8J�cJ�d�f �'D�k�^�If"O ��a�Z�yf����${��s�*Ovm�G�E�[6�QW�.�@8h
�'U���u"B�w��C��I�P)�K
�'9���I*JM���&ry�	�'@&Ѐ  �t��h&��>�	�'7,y��������[j�l	q"��y�śE��5#%��)O��Ac ��yr� � �����?6�k���y���az0��C�6zp�0�KӜ�y2g�T���,�rP�cML�y&y��'� ��˝m���r�N�":L�c�'N�y�ҧ��X�.�� ��4Ap��'������I��t�W�ۀ��k	�'� x�����QG�Ɂz,���'C´A`�A(4p@fɀ�p
��S�'�^%v��k5�D�� V��$�
�'�^)8�	ҧ>6i�s��?�B
�'��:�A�^Nx�!@G#;���	�'ޖ(X���3v �b$ϖ	[���'���R���8gڙ���:u��i�	�'��qs�<6�����r�&���'Av�����3H��Q�G�n2�({�'f�m��d��\����ǯ"f�Ma�'E:���P��a�'`�L�'v���#�(8���Q��!f�Ri
�'u����6�zI���^%�0�	�'��Ń�a��)���ui�Vd���	�'�x��C��&9��I�n�����'� �C���#{*�J�O�2���'�P��Q�Wv�R��5Ӯ�q	�'wFL��!)n��I��C g� ��'�p�BЏ)���ةnO��8	�'��L����-<���Gc����'}R9��c�j�����X��)R�'�(���g����fL�~��@�'�j����ΑjH�ջ�+ˆ{�A1
�'���u�ByA��(�� g�e��'|E�$L�T"@�C��b�hyB�'�6�����1�I0iB�P�4��'�8ʧ�Q�&BQR��S>w�NIH�'P�L�Ȁ�7���xS-:io����'f��[�n�/8Gxs�+]v~,j�'�lK�[!`��r�&NF|q�
�']����}C�`����J���A
�'XzL��}�x �KL8U��<
�'��1��;i¬���S�O$r- �'b��p���W�����Uo���'�&��UD��]�t`�!�{��	�'�V-��NR�dk��s�n4��'����E׻��Y��鐿i�u��'(��v��e����n��a�ı�'���;�P�� ���@�^����
�'h��遍ǻt<.1#ӎB]T������ ^��u�#��4is˝��8�C"O�p±��-a��$3�E�, "O�������[��L+G��a�\��"O�U��	-+ܜ��H�2+�!�0"O�� �I��T�	7'D�
G�s�"O�C��
� ��A��$q  P"O�� �jH�r�r���-V{�b��q"O���A�V�>�z�mK�x����"O@А��Q�k֒D�PGI�.?
�XU"Oح(AN��p�#!��Z챢$"OƄ��� ��9�!�3��T�b"O(p#�.ː.��4JG���~�򉺒"Oz�`!�I�K��I���h"O�|
qn�iOp�S4�� x�vӧ"O��ö� T�@�(�m� !��m��"OZa���-6�<�"����D��I�#"O�ـ��ޘ��[7Û,`����"O���fֆ�R�1��;����"OT�1��9ee.�rr�5 �����"O�!�s(zP�D�D�ݺ`>,�*�"O<��dA5rt��rd�e(p@B"O�xS����L�{N�X��J'"O����,T}~�d-��	 B$"O�����X�����԰h�]��"Ot�҇�Od�*Ga��;�TD��"O�U��A)'MD���}����"Ov\�$��!E�H��kn ��"O�8�񬒒`��c�ꎧm�6$i"O���raȗi�� ʇ�	Д�0"O`x�d�f��c�k���X,��"O��*���uPe2�S,��ݑ"Od�$J:��Eq��3���""Oz��V�Q�h��\!0o����a�"O��Q�!����� A��yj�qv"O�|2ç�W�д�ɐ<xŞY�"O0 A!V#L��Q;��7H�){�"O�qRv��Vю|�疙T�R�+0"O$E�5N�^�I�e�\�y�=�"O�C�J1@��H���&e�>��e"O�ܢ��ܭR::!�YR�2-b"O�FO�xY~�Ip��	���#�"OLTi�׭stX��J]����s"Oz���L�n�( ��S����"O~�ك�B�:�\3��ڹy,(� "O ��an��j��fDt�x�3�"O�Ms�K�2\��8�5�pߢ<�Q"Op�ÐQ}��B$V�B�	"O^Q6�B�[7�܀"��;�Z�
s"OPȠ��0f�80��;���4"O�xS	�"K�vԱ�"�<ָb�"O�h�k_���u"A�٩H�yڑ"O��3�K�8#��E�����"OV��s��=i�-:Va޲�腁�"Ox�{5�N7Y���R3T�r9F"Oc"��%�֭̍$�D�d"O<����d���N >�-�"O����M�pY>���CPM;�"O֕�0b�,
�Y)�$����2�"O؉+5 D-pK�D���B6j�T��`"O��� E'=bH�����y���9�"O:]��V2qˢ��%3��Ahu"Orl"bk�W/V��2f�r�8�3"O�P!A��;Pz���S�E��"Orm{g^�&�"5���F�v�K6"O� v� �l�81��1��C�4j���"O� �7kC9ki*A����(J��y�"O$I�s.@(#9���b荹+G(�xw"O�aU.�>x�����
If�R�"O����ϳ ^�aC3��'��H��"O��*u��
APS��x�p�@�"O8���n�o�X%����'=V�`"OD�"
$�x�J'C� -4�xV"O�q�E4.�XH�!Ó>�p�"Ov!��/�% �e�1��(�Xk�"O��(Vn�� ��iB��"Od�6�R"Q���B�e�Taq�"O�#�z;�Ѿ$�D���$�!�dB�y�p����_͐�i$��H�!�D�W�hD�f^2E,]3�-��rY!�d1s�깰���B����3�!򤎕[�PX���1T�!��͑�!��I>T�Q� �:H��E;ԯ^�<�!򤄐�
���J�1s�m� _�!��ܷD���!���u4�Pq�j�"�!򄀘H���xgn��t�,�9Ri�(!��S�Fo���Z9j�I�E01]!���I~�u8�%���\Y��H��P!�Dv$��͝��IҬ�i�!���xJ�Q(�bV8�0�*7E�!��' �(��퓝BODe�A�N9cv!�D�W��3oܫ:I���s�Ax!�U�6L�=���Z�aH�M��B�3!�D^T��!��̜�tU.��t�W�EX!�DO$1��x:��N�Qd��vF$X!�ܶ(
:P:L[
'���蚢V�!�ğJ��!� �8E�5eԅn!�䈺:;��1�D����+�Ç`!�Da��I�#� �u��Q���g!�dGNO�#aBM�ݞ�q&!��V�@X^�����6��!(Ӈ-�!�4�;��1�0��GK+4,!�P�7<��iԊZ�K�Y0�`EC!��[�$��٧I��0�A���^�!�d�s7V��m� f��QJ�(�	tJ!�d؈Z�Z�����`ȧ26!�BY��)�b���<g5!�9e5!�$�0z<>����r{(��b�×�!�=i2�C�!�?E"1�)�!�dڄ��Tq��I�<	�1�tI/!�D���Zu
+{��%����r!�dZ��*f㒋��z�E�!�ډf�b��R�V�p�*��Mڗ^�!�ĊJD�p�P��`����1]�!��8:� 1�EI�;� ���Lս �!�D�{.��DD��V�nt�� s!�D�PN	�G�W�i�P�S�!�+h[!�TWK}s����ta��bC!�d��=y�h�)��t�^��ᮐ�A!�$�*p���0�jT�����!�$U:l��I"G�U�.��"�d�!���k���$�HY']�!��5 l�"2,���R��%A�(�!�Y�,�P-�҆�(3�8e���#j�!��PR�lH�0NK�O&���e�!�č7�~%
W�O *�� ���)v!�ĕ*����B���������Q<lz!�D�MX�#�Cd�dA��T,O!��b(N��`�\!0xz��Q�]�=*!�� I�p��8&��FFJ3dЊ3g"O�Yj0��<=.��cfY3`���4"O5��-I�;��9�1o�SWL	��"Ozj�� "+$�䛒N��[)�E�"O\��홌c�,y�M�3nܙ@�"O�uA�JR(Z�����M
>#|Z ��"Oj��TI�H�8�-�vc0��R*O�%�T �'2�+��r��r�'��I���ƨFzt��e��[N���'�e�#�X�*Jق@�M���
�'_�1)�EZ�P��՝R!���'����6+Ʌ9�4)�ԦOO�K�'� �1�Aq���{J� =�pI
�'v��٦�V�V.8�@�B���S�'ڸqQe�*�bТ9�����'��	/�,�#�O´Y��<�!쎶�y¨�)Kb (A�A�?�v�+ƅ]��y�ʱ�Iӯч.a�����y�a ,��e���N Y;\ȩp.I��yr/WNj�M	d��N	l; `��y��ر1�Vq��z��9�'1�y2��DT�Y��R�hFRH��L	�y��D)�:$�vc]�k�(�q-�)�yB�_%�����z�fY�u% �yb��U�����!�[����!	�y��
S�2�1T#�,U�LC�	޴�y�뇜J� ���=����f��y��6�(���A�	b�蔌O�y�j^kM���W�B!Q�R�u�X��y��!< ����"C�X,�P���y�(��*�W�	*۪�)�����y�j�SW:uPӉő(7����ۛ�yb�ޥ�Ҡ�郗J��e��A�7�yrbL�Y�����%��2I���C�&�y�� !|��6�M ,�2��t��y"A�;[�� �E,�'vh���y��.>��(rN��!�,��e/�y�
I�X�\Ys�/�� 6�y�jǎ_�RЊA�)=����yҁ�?T�l�@MP�%�Pb����y�͜��D��jQ��4��.��y�!�+a܄�@u�H�d�����N=�y���]HN�J"��Vl���c��y����f��0P�@aS��@��y���wM�rD-�[FT���b�=�y�.2a8K%+�@�p�XsM%�y�Jڰ+��B�&�2}�:����yB+Ϗ���r,&%���kQ��yB��$��H�ebG��0c � �y�Xc~��J��Ȫ1���jGd�&�ybm�o�1�M-/�J�@��y��[�f� 5(�u�M�Vl���ybL� bx����� %�@%�E�G�yBA64�`��	R3 �>la�eH��yǜ�\�☚���T�����y��ob��"��#T4��Ç�?�y.���Lk#���-�#+��y�Gb w����v��y� C�(s�=.i����W��,x��x���R�
#G.�ҕၭ4!`u�#�<D���\)�����-.*�����y�ӯ �f�D,0��4P 埐�y�@Y�%�	gm� -������-�yE�\�Z\����J'pYsb���y
�  ��a�2*r)�*K ׺1Cb"O�q%�̹��̸-���c"Oz���!@���3a�:t�ʕЗ"O� ��CE�FE�`�� mc�"O�
4��}X2�c��T>Hs��0"O�X�EV�?����ŏӺe��)%"O�	�d���l8�c'�QRZŹ2"O��q�B�=&�����]V�M��"O��
pʕ�$��P����.GZ�g"O�x�4�N/$#	 ���%A�̙"Of�u	��?q(�J�!	��=�&"OfȻ`-��slȁ� �̥op���"OЭh�$P?�^	Q\�J�����"O`Cq$؇19T؋i��0�"O�0̀4Y��|{B��	����'"OD(�f��!�x��G�ِ\����"O������=,�`�EN.z��Mb�"O�us%I�1V<�j��`춼��"O�qC�o��������:E"O�� ��E*)A�\��K�
i��#"OA���fsD����4%M��"O�m�E�ߧe-���ǣ<6�At"O��"6h��Gch��d�հ��A�S"O^�+�/�n��7�E�[����"O~��qcΚ@f���X���k�"O�(e�L�	S`���&��"O$�"��<|��Ex� B5}o����"O %��BvxR���o��Ea�ԣ"O���x�q�!D6+��r"Ozi!�'�ؠ �枻�����"O���0��LVy �&�l~ yb�"O�Lٴ�?�A�1� +u}0Yp"O8)l��F$���C�gt��!�"O*8��$�0�\�"K�&ְ��"O����O���3���!�A;B"O�x�C	_�L��i���6��"O�bFH0?"=��͕���1�"O���Q���>�U��`���ҽ��"O\I��_;x�3q�L�����"O:��cA]��
M[�D�IRzQ3"OԤ�*�+����m	`e��"O��"V��L�x|��a�0jژta"O���j3=��1 �D}��T�"OZ�"ȫ �L+��y��t��"O�*��R�."�pcK�B�V0�"O��;#*B�|���� �!s��y&"O�eҵ�����ap��,�Fa9�"O�9�*�%��l��8�J)!�"O�x6��~z!kp�5=���Xd"O�(`G��x�D
�@���\[�"O&�q�/�0*/Hi�u�1�Nx�"O��J���&0�P��l��X�$��"O��rK	 D�w�ʿ,���"O��{o��|����)GY�9�"O:���*�\;���p�Jd� "O�|���Ƣ,�4ԣ� �M��82�"O�H�2J�'IG�8b� �8 A�"ON��E�nݰ��i;�%��"O@�#�I y�|ɫ���=/�ࢧ"O�!��J%Gd~`��ώ���mhp"Oz� ��(�F��(�&�p�"Opl���Tb�h�2���:i�D��"O���LR���1'\�OY���"O���7fZ>4r\�(I<�\yQ"O� ��y�f�Sz��[S/��:*
U�F"Oz�8u%U
.���r�Q�a�)i�"OH�ٓND�|+�1��	�{�"OVIx��oP"� �ޮ?X��R�"OLY�F)�|'�0 ϹH�Ш��"O���
@��U�ֆ��-4���"O\8�רե8�֩ �%>(jIcu"O�Q$ B�N8���	!�"Od@ㅩJ�@�VeIU��)9:�ӧ"O0��S����|���*�Y"O�<�r�ͻ9��S�kMӲLH�"O�]�חb�$��dJG� �qa"O`�`�00L�Ӳ�!d��,�"O�����L/��g"D���b"Oʽ��_P�ݘ�S�4�>`@�"O��)�b
<�bPhdF��mo�8�e"O��kf��oh���N7$4�R"O�9��b6EA`����#h�@"OT�j��10b�����ƹP�Eb"O%a�"�Z����Cۜa��E:�"O]suዋpbH�DG��h1�"O���ħȑ!J�U��+�2�YQ"OD
�[s7 ���/�4y~U��"O�	xv�ަ:�&��d�H0Z1"OVI�3���=7 l	��D�~�Lx9�"O L���K
U��i@A�64�9�C"O�����@����W.�'=�T��"O�=�D%'0Ȕ�F��q�.���"O���E���Ts1鈿pj�
�"Oڄ�R��-X���i�`l0�3�"O4d�A��H�%Д��d^��k�"O��YՃ�iI xQC6*jd���"OD��g�X+gB���.݅2a�M��"ON�I��Oj��i���y�e�#"OVDyvl��9���U�:�2�"Of<��dI�x��99'�Z,�n8�`"O�\���|v�6ø��W"O�!�a�ҍp2N��2' 
T�P�"O,! �dU U�d8�q���@a�"O���΄� `��A&a�$��&"O���g�2�����N�
:���2�"Oؘ�U��F�2m�1�|-�0"O�:�&�H���
#ܓy�l�I�"O�ܠ��̜{��(��+�|�P-��"O�q�߽�� ���#��@y�"O�`�e�&AV��2i��m7,��"O~ @b�P�u-l�83F�8�FE��"O����q���ia��6m�,�g"O��#�
L�g��y3O�- O4L1�"O�Q�Wኁ��:���C�L�"O",i�^��H8���5o�`{�"O�� "�Zz´p��G�TT�"O&)�qf^�-al���.��f��"O>�	���+�P��r��#���Q�"O�Tj�+�V~	R�ɞi��Y��"O(�hA�{�BX��8*]q4"Olt�D���K
���� �
̆�yU�:���7��������Y�y�� zM�q�$����T�t	�1�y�➆(�*��qdY�dF�D4h�?�y��E� ဆ�OV٩�A��yr-�9JM��郢��.س���y����a���0/Z5	|�
�j���y"��&z2���N�0Y�|�+���+�y
� $#em ]��`�C�Y��y�"Oҁ����|�i)B&O�Ig��P�"O�(U�f���CuD��=���s�"O�2�O�!`!@�	��+]���"O�YYN�<���7	�.<�h�"O@uh��P@^�)!��>;��J�"O�8[��шG�m�Lʫׂ0�w"O���`ڊz��ĳ�i��M�ޘ�"O���E�Aw� xI��D����4"O��ǊP�T��AY��A���P"O܁��iV1}jƠ�M^�9����"O.B1��;r]�a*E�8$h�В"O�T�D S� cHݍhX�"O��Y&�?���s(	%2	�"Ot�S㌐�{c4	@��:�l��"OP�3k�8n1f`�MݫB{�k�"O�M��C.@.�u�0�N:,�:�"O�\�S���$d�ł�pqz�8�"OZ�(���r�|��q��X����"Ofx���?���Q@�Qj�"O����C�؊aK��2�-��"O�pb���5U>�@���%��:a"O�t���O�n�,�1Ӯ֩s'����"O%:5��7Ը��Ȟ.5��)@"O��*#��Z�ZDXR	��=C���"O��!?'��6���l	&�� "O����^��<������@��"O~��'GH=/:^	j�K%F�*�Q"O��1!�]�Do��׵(�N@bG"ON�[��K$4�<�Tŕ��f���"Ov��"�\?rjx4��^�l]ź�"O��j��V�L^�͍/z�Z�"�"O��AkV1�8�D#�F/P��"O�Y;v�J�8[�%����1p]��"O�%M�ZBѢA*n���X"O�%A].R�
�  @M�7�,�ڃ"O9�%a��"�O��3��B䉣պ�ZB&��i{���烴K��C�?�$�Z��W�WM��p�g��P��C�ə���ۂ����pY3�?�lC䉁
O&�Ёa�4V���QpK[��NC�	�_X��Y�F�/�L� �Y�|B�(l�"��v��3�jd!�V�@�>B�I��j�C&�`(x����H:PB�I�>�ؑۓ�J�?�v����J�z=pB�Icq�y��+(�JE���һ�B�	a��dA�S�.q��N5z:B�	�_xFlyq��� Cs�̼jĲC�I�W���G�8;���d��'IrZB�	����ʕm	�Q$8�sB$ BvrB��5P��E96K��0d����6�B�I�r\m���ϰE��(bOڱTc�C�	�l�ZL{f�فf�Q8H� ZdC�*O�|]
��$F��IQ��aFC�	N�Y9g���l}�a��C�	�mLpب@�ޡYWha!O$ ��B�	m\&�h��C�Pz�󗆍3��B�	8p;ȍ��W5z/|ѨF	�#Kg\B�	�jF+�So �S���'F*B�ɒe�q�QM��,�" �#DH1?ADB��$ެ��PiZ&�|�p�+eg�B䉊M��lV�ȡC�H���F �J"�B䉾0^���ʔ8 B��4��Z��B�ɣR�4;Bkذ(wN ����	2��B�)� �dzC�� �&xUĄ�y�&�0�"O�(��?�(��ՠ.ǂH�"O��8s�\���"��%u���c�"O򰡓c�>^D���G�K�����*O�Yd'ߡ,��XB#;;ĕ�
�'��݃��K  �K�z�p�q
�'�L\��\ vՐ�(���(l� ���'
��;�I	�o��	X�kG�5���'�Vu���
J����#H�}*��';,Y�Ŭ܃����
H�w�d��'�
H��,�L�L�s�D�q!F��';d˧-�B��勌�bJ,mB�'l�Hpp��N}��+�؜.|*���'V|L�b@��k���z�ڼ!{(H��'�(�J҇m���Y��\4eD�z�'?<գ &�W�8�i�FM�v�=A
�'4���J ���d8����9�	�'$!���W�D�1���>Q�	�'�R��陀lR�y���/vR�mh	�'��U2tm�8 o�v��e	�'+(`�wgB"4�X�'�جp�6,��'S&���/�,O18��3<��'q>}����W��$J���'3�a���'o�&|+Gؠz��Z�'�,u��D֥B,q�jͪu"DAQ�'��%xfU2I��a��
p��Ic	�'TrȒ�Iˑ8�T��Rmɉn��r�'�^i�`FZoH䄊芷0����'�
AccW�L�D������>�*���'��SkU�!�*ђbHD�;�ֵ��'���Rtc��h�z��!�5�t���'mXK�-�9
�J�x .[�o{���',D��T��_o���Ǣ�����'����D�@Ų����P;=x�c�'/@�w@��~S,Y��(�!0)�H�'��t4�� j�ܨR�G�&�!��'5���&+��\�b�	G�%>VD��'"6�h��A�N�aZ��=5�t�
�'�eP�oZ�.S�U��+\�\��U*
�'t�eq�m+,
�����V3f��	�'`|�����_��AA�ŘmJ�r�'YL@2p�E;t�j��R�ٗ�����'x&����4)h�5�
w�i��',�pY���9u߆1K"D;v}H���'�]���R��E؆� !B^ �P�'b�x��a��2=^�i��C��ة�'g����D(,R��I�G�&��8�'��Yu�B<7���N��4k��'���Ёj^���L��ʌ3�d݊�'hR����<ά�P������
�'�1��IV=XK�
�vf�h�
�'�(��WM���PB"�>r�|��
�'��m���<>L"@Q@�E��N�
�'���)5 V?gz�w�T��\a�
�'���oI"�\�e��s�,��	�'#��gɝ;C,h����6mٔY 
�'�@,P��ъ.\���f�~�B
�'�Z8�`�wzDK���i�r̓	�'�Z�!���":��%����O���	�'cjMx�+�g�&Hq�N�~��'fN|*�ˇ
�:�� �W�P���9�'�8���EZ0��MI�O�����'�D01J�^2��M_�J8[�'��d*�H�s�2�ζU⾤���� �d��X "�`ݠB�م5�����"ODq�Lɂ>��!" '��7<��"O�-Y��7���[�lӄt5��pV"O���3Jg�9rM�0M�r�`�b3T�Ę冈h
��j�@�h?DtbD$D�cǀJ]Э�r��
�:d��6D�8Z��Т5e�k�1�:��6D��J�M�`y�(�/�<!�2D����L�E�``��My��j�-0D� yL�.ST�y;�,M�T��L1D��[p启G�F%h�.�+V颍�w�<D����&ړV�Xa���	,����Q�$D��Yc�Iv�^9��#��_�	���"D�|	�VC�P4rԪ��@<��4g#D��IC.@9BPX=�T����b�K"D�X��*�2j6���)7 		� D�L��@I�L\d�v��e��0c�@4D�kc��L�`M�0��E���h3D� �F��	V����/{�4����2D��!�&��rc<)�`��"g�ltB$�;D���Z&'�ZD8�ٞy2��֢8D����D�Y��Y�cV8B��@�!D���e`�&u�P��`O�g���å�)D�$p�� be�l�4��e�L��A3D��[�@!=r4�#S�K]�qcР6D��z�"��n\̍�w	VSz�����4D�`/�ZJE�կ6�1s4.>D�r�AKB�Kp��_�j��E�!D�;r�~a4a��S��;��ӫm�2C�&�f@�Nʱe	�x1F�,? :C�	�-v�l�Ėj�ʀ��BK�c�C䉞V�����6J��+毓�e��C�1'D���T�\��Svȑ	l��B�Ɍ�a°/�w�Թ�&ɓ�y�nC䉒UK�}�Ѭ[u ����14�B�əa�tp�)M=��I�`�-q�fB�I�=���S�D��sa250�B�+�h-s�[�miZ�0���2-�B�I�LLP�0�*\D�X�7�B�	�r�`2ad�)OF�e�-Gq�C�ɑNގ�1�G��o��X���&ir�C�1CL1V�^	��I�H9K��C��3xr�i�[ԅ��)��<�C䉠�b�b���DFd���έP�TB�I6d�
��RWR�Z�o��A�C�	�2�rԦ� qjJ�8`�1W�B�I]������i:(1JC��5��B�=�
��dC:��	�#A�OhB�I;�R��N�DBpq���2F�0B�	*0$%JAf�70$80�G �n��C䉧G5f`�6!	�z���1���C�Iq�����^�q��5I�(W�PrTC�I'M,*��F�5��Q	'$-aL"C�I�T� �0S�.T���Pob���"O���3a�&͠(�'C/	T�m*�"Ob(ʴ�3-D�1�� GJ*��"O�a���
и�\�Z�tz"O�ep���d4 ��
�+��;�"O~D�0�M+%�����H�6��5�P"O��7D�LWֹu�Q3R��0b�"O�Yj� �$�2"��fV��� "O
U	(Ȃ~����EB8~H�0)S"Oؠ*D �_�NhK4��'a:�``"OLi�%"_�&��� �"�A$$=�&"O� �r�h� ]���B�������"OT�F,}Z���j@�T����U"O���'G��CRȠx5�Ȫ-�Ҭ:3"O&�A@�/-=�}�7�ͱW{6��"O�U1SJ�cV�TN֨P�"�92"O e��"_�G���a$�7@��)�"O4����"���g��c���1�"O�8ZdbA�.�.��p�U�� ��"O�pQ��հD�Lp�&Ɔi��T��"OH=�J�E
U[d�V�&��P"O���&̃E�h,֛K[έQ�"OV����VST�P�똗YM\�k�"On#��,+��Q˘G^���p"Od���E�?�����zp�r@"Om�2� 2�3#�5R�KF"O��˃�F��t4AS-��`�"O���E�$<iXAh�@чsl��2'"O�D��@�2^��EO�IV�`��"O��{v��AH�lA��CH_J �"OLl(1节X�`la�O�-BRԑB"O���CA��ӭ� J�<�E"O����˗ ݀���[&,��@"O�d�@�p�zl۷��:M� �AU"O��!\xL���o�1��s�"O�%`���K����ْr,�i �"OD$�3դ�2����D�ap�#�"O<��ϕ�M�a�Fϟ(OX�*"O�}(6�S�H����rfL1afEô"O��5艔z~��4��cS�p�D"O����a�y�������l�7"O����49�l�P �oC�ɸ�"O��K4cڋ1ѐԀJȆI%�]+�"Op��Y؈asL�:,���x �z!�D�$t�4҅ES��tx���!�^({ʕc��^Vǈ0b��:H�!����Aa5�!gŚ)�,�4�!�>Q��b�� �(��0��l�8�!���.U�ݺū��h
����H�~!�\=��L�s��	�0+Vɓ�ss!�I�PJ � Ci�/I�@�+���+�!��rȠ�gK3j�d����Bx!�Đ�("��y�.��i\չ���:+a!��ˀ0����kf)ɵ.ڡ]D!�$5aB
q�F�])ZUl��1<!� �"=[�J��~�n%����8D.!�$"��x����]`�����G��!�S�
NU�qn_
b��B�%$S�!�F�@>j�[�FH�PM�À�D�!�JV��Yȃi�,!0 ��r�!�d�V�A�R�
�}kX��gÀ�	!�R:pW�c���#e ����!�܉=�D�ڣ*حP���n��!�� ��z�"�*Z1:8r��T�!�d\�i�L�#瘾<%Űbn�)#l!�dH�u��*S�X�Y�%��LT2`�!��$~�љ��ĄG"]@g��Q�!�$�(K&ap(�,NX�KؔaD!��$?��D�a�۪|�`� �I�:W!�$϶�ZL��-l���pə�4!�߮,�4�m�Op��S��ɜ�!�d!(Ypfy���@�e�<�!�_,jH.��r��?v�$=1E5�!�d�lU(���G�*���Hګj�!�$D?�`���.ב����D@�!�� �Ii���~�0�R���>4�!�$"O�9� և%!V12�nP�6$��1�"O6��6M� h��T�GK�i�G"O~, WE��2�%��E�:P�"O�������U���H%eDN��P�"Oz��쏙�4q3��&*f�5'�'��'z���]w�T�b��#-t����y"��,j�
�"Ń°,����jÓ�y�&�V��ఉ�?V'��B@�Ʉ�yBFݕ*�����k�%&j(J$嚰�y2 �I $҅�M7�P�Y���7�yB�۞��t�@f��|�`lһ�y2�I�[!��(<8���ϭ�yr�F,P����T���ϰ�y&�E��*�B�On^��DE���y�oW3|\��C�� @x>�*d�=�y�N����hԡeL�(s�V��yr�� p��Q��$X�B-z�
ʳ�y�Ò�U�~�"�
F1�ك����~�)ڧ,��Q�B��b=,1yq���6܆�Q���	0���]8D$	R&I?h:�Fx2�'!�<8��B��8Zt+ 3S�\�˓�(O��B�#Eu"��ǃ�x#�:�"O޴bG9�����b�^��!"O��ђˇT�>d�0&K�q�B�'��&^>�a�@�i��sՆ��CR!��˻�2���F��2��U���
]G!�\��H�I�@��mᯒ'!C!�Dמ,�ؘ1t�2YՂ�@�@�'(!��-�����p��� �m!�ď�Ql����ɜ_��R�oZ�b��zr�����e�P,2�<=���Ȋg�!�D�L}BI�G`�_zMd)H�!��$z�j=��/��2�B�'�G�a}��>��	Y�8 LY�v*���Oj�<��*��, �u8�n^�3���ʂJ�<	��U�FZ`���g� �f�B�<y�l�"|����='n�EX�nD~X�����z�Z��P4нK3"�����ȓl����E�[��`�a�J�9j�؆ȓ_`���� SAg�^�����&�99c�0�<X�&B6�P�ȓg�x)�Dn�3}�Y���r���D{b�'�\9{�U�F
\z4�F� �q�'i��x��=���"��.!�5��'~|@����G���Q�@���L��
�'��(A&aܖN[ ��#��@��y��'��E�5@�%,���":�8����)�ԡ�;$��0�e�.QG�C,	.rqOf�)�3��8v�^�s�V�$7@�ӷ�E�>B�''ўb?	y�@'e�4Z�d`��P� �%D��5�؂���Dn��%	.%��ke�|�Fz2��0K՜�����[��Q�V�u/����v���SL�; �慛�W����e�#��<i.�M��,9�>%y���EoB�I#ʢ��w�,>v�)e��5bX¢<A�]�^8I��>O��]ܒ)�Re�ȓ[n�,�w��.Ҡ1R �L�r�ȓ;�,mCr/?����r��)��L�ȓ}C~���[�e�(	"U�k�  ��kh�ٱc��*Q�l�$�p�N���&Āl��č�J�� A����a�� "�lY��D��`��|~P<�ȓv�ص�Y F��P�vj
A���S�? �|"A��:5}S$���oV�eR�+$4� �$`�;sǲMjԣB�s-J���g6D���M�E��y��+lF@�ђJ'D�$���,-�=BBB(@�&D��iׯ	�>�PI%�*fxu!��%D��K�.�.� r닯UExU�7$D��òg�v=y��ʪhT���C$D�P��ҍ8�\�+Si	�8����,D����-�.i�6� ��n�("b>D��R��@�o�
xz�DŚ>��i��&=D� �!ʋ�e`XU�r-�d���R�5D�Lc��]<2~��Rw� 0��Jv�0D�W鎻BZ�с�ۃp��3�,D�dC��YoR�;4�ܒQ�>$��O D�ܢS
N=���tL��k����>D��H5��|/<M �¯Q�ܵ�� D����n�,��A�n��,��UHr"?D�$�D/�.b�4 [��{��|*�9D��ȥ�?A�^82��b�hkAN4D�tJ��)q�h1Zw��O���h>D�����&e�t���Oe'�I4h;D�$�q�8�(P	�9N�j�h��,D���G�#�pT�7!R���E/D���$���p჏%���7�,D��b7�ʘ�=�����Y�&�8D��C	�rҨp�I�15�B�ف8D�l�eіh����
"���� 6D��y�KN����p�l��x�qK%3D�,�O�;�q�a�8"ޠ��2D�h�w���W���"�oR$qXK6D��H��^�Ep�h���8\��5�!D�ph��_�hp�irD��7j���h D��3��:D}���"GԗV���w $D�,���J��!�V�Ӵ� D���cO9C�><�ӈ�[5���O;D�D¡/�"de{C�� -N��a�:D�,h�`��t��"M�"91wL.D��P�ŵ~�D Yv�� ��L(��*D��c�|��]�$��2�lY�(D�Ȓue�*Q��"p�\�DE�5*OB��"��2ߖ$SG"%�m��"O8<���$$�e��g��	c��+�"O�B3�Ν?��P
�h[<}v�"O.Qy�����,[���(b�@W"O0a�Tj,�Ա+���9x�P�S�"Oƀ���&o�&u D	j�pl�"O��9��Պ�Ԉ$e�[�h�8�"O*�����HГ��N��\�"O�Azb��e��*��\��j�"O�e�"��t&%�-�"{�y��"O�[#L�,>��A���gp���"O�0��g�����b�@U;	�P�B"O8�'� �B���
^Հf"O��4��f�l�C�V�\�Zԫd"OEj��|o �3b���[�T��"O���'F@T�y8��2� �PG"O~e����_���I����Lh $"OR��1��)[Xl,�H�9_��!v"OP逷lM�1?���"�T5t�D�˳"O�ifO۸8�� j�R��"O�9Q�)Km4.�C�Ԇ�:e�"O�5Çe�zx[�!A7�hu G"O�17j�2�΅[7A��U�h�#p"ON��S��2`?�!� ��p�j`k"O� .�QE�� q��� H�D�l�2�"Ox��W�
\��(	b��0�j]3�"O(#7��v�r�W'��T�	�""O~Q
Ԩ�#{����ED��s�X���"O�%$���ڳ�Ǜ 	�m2p"O �I砌 &jဒ��-��� �"ON�07��^�Z�� ����Q��"O�Ay�N�:e�1���\�+�F���"O:�Ȁ���.p�4�У�J9#�"O$��A K�Ըq�_�:�X��"Od�+�����LЃ&G:V)�-�"O��Ч�A�����+�}h"O���͔�1Re�e��'���"Oȋ�D�"���'��:��"O,5 o�>+�0��ہg�=�"O���D� �$4BI�),Aa"O��A�ؑ/^��k �J� ƍ��"O\�`�#�� �w���v���q"O}I��)+��a�ɤX���R"OV��6����l�7
)��R"O0�J0�Ҝ>D�ĹR%��R�ڵ��"O0�@P�0c�03ET�H�r#"O�Aj1��Xj���"��Q�� �4"Oj��kF
\����̋���g"O�� ��
�qY#.W(}Y��k�<Y'CA�ni��P95�x�,Y	B�ɼo�d|Q��N?S�4�A�Ş.B��$_>j,�sLɟb����E*G����2K��ћ��T N8Ŋ�� �}8J�X��Q6~��,a�ŕ�!��>^� R�!lʹ�ڑD���!�d�#4��ZE$W9
���J2#�!!��ʜv�JU�kA:�zD�6!�Q!���/x��}:5�U/< �ai��^�!�d�	�69���YO������W>w!���è���
I���xf���R+!�ċ
ʜ������F˝�J !�8 꼰
$�8��ŃG�V#m"!�.r����"�V�&�p��S1t<!��āk��c�ʆp�0e(�M�5.%!�Ċ;/[HXB�'	��bhaU��@6!�D
(͌A�L�:v%�`&�u!��Kt�q��:fB�0��&��!�[ B�IHdE�bg~� ��.!�d��w�8��f(DYO:�8I
&7�!�$G2|����*�{5�ő�!�$M�W|k��@0	��9�g�
JT!򤖩�|���E\>2��)���N(i\!���k~�(y�B��q�fH�(�!�$<H|��&�=�^�y�A�!��p��q8�L8FÄ(
�%�!���KlQ�G����yR �U;L�!��2�6���,�& y�A���&8�!�dө=��l{����Wۄ��!�]�pe!��8x�\)��Ю`Ú4A�b!�>�N�W��xPV<��(s^!�$���t�: ,Ub�
�����L�!��29X�@WZ��q2P$C|!�DFM�J� �K�zp��f��zm!�D�_��%I���j5�IX�FTJ�!��O\��3V�Y����d$���!�d�$(& qh�Y�� X"!�$Q�B���G�C@���]�!�d̀����U�]��	�#�/=q!�dDkF�2t�ſmܨQ*��e!�� ���Ã�
�"囄Eه!�ؠ"O�i����U�^� D-U I
A0F"O��"!-
MY0��&	S(��"�"O�Y@��ЉP�P�3A�C�B$�"O5HaK[*�ڰ�uC��-�:dJ�"Ol�(�o��l
�][3+���0�t"O��rS&V*��!B��Q� )�"O~�v��qN|مm��r����"O؈Sf�ؕ8 ���D}�x�8"O�y����=��	)���6X�b���"O�H�F��I���3��� ^u:A"O��w��Z��MZ$C�;��K&"O~͋Q�\�	d����M���"O��s �\��Ap%I� )��|��"O�(�J��<���@5J�Q� M�q"O�[���	�V9K�J �x�R�#�"O�y��ɍ��1��wؒ1�"O�	���"Y��q��'78,��|b�ŧ79(�=�}��.@+2�C��m܄�G�k�<��H�����p�D�*@���,,5�,O�e!�=7�1�1Op1�K��kzF\Xr��q��]A��'�t9 ��E�M����$ň0�+�)[�Z8��D�?��M���yJ �օC\�h�A���"?Y"Ʌ�,����7���`�O\1��e���s��J���#	�'�0�H󉝞L�h���@��N0�!1+S4������<	H��d�ؑ�6�@��4LHɼ3�F@9Jp���Ԩ��	Ü��`��Rh<!gh�&�D@H��	�~+�8�oH���|�`�d��89��EDD��$�P�L$���b/�	�4L&���P;(/�l*�&C'�^���ΖC�)�.�[��
�D��'n˚Ka<<᥉<��J�N�z기�DF�\����]�p���A��h��\���w���sҔ�r���lꚥQ�֚<�Yi���/���ʶ����d��aC.@@l=(�%S"�a�*(D��0n�D.�)��S�XP�s���Ĩ$�V0(��U��<�4�)`�F,�>YD�Or��À�[�@�HB-��9���Q
%�OR䱃 �?Uf鐓MA�U,�8�1���$��@E��>��R�"2*�<�q,C�]v����/W)�$'��%�̿D���z�˂_P0C`g!�2�=��+j) ��Jx�jSE��@łP�d#��$�fp�P�F�(Y~�b�L��K?�zB��l���G0kHpa���z>"�*#�E����?G�N�ˑi֛&T��g��'�"�;�腾�l�A@E
8�I[R"�#VԻ��U�(�y��H� &���"~�]B�؜B$q����S���H"�_�p��I�$�,2��uhُ'w�}zǮ�@$}��?W���̻:���0��,D �I�(�i����lq�!G�ǽz4�i�̂�F���AR�
0pأ�ޘW�2�i�đ>z>���>|:��1E�CN�O0	I����>M�Р��z͐��e�	<���T	K���3&Ğ� ����c�8("���@�t`�X���-�����^� 	�&A7�h�ZÓ��i	�ĭJ[<H�6�F��`�'$hE�A�7d{vj�gʈY���Ǣ��+�mc�gG vz���ID�8e{OM
*�\lQ�
E�zYt�3����/G�I����`��3=�:��0�N+}�f`ٴO��.��7�ڟ'��ԉP�ò?�*���co����=O�=iT"��M�x��l-�O��ه�ąX�F����1��%���$n��%�-\6B<#H�_<����W�\�R䲵�E�5��1���|~���,~�H���*� }���$��ONhѓ���K}B�ǉ�aG*U�5"D�mD��5��BUP�,k=:��$-*P��,�H���RX��Ó��0<iҁĒ[�4��a� $)�mS2Cc}�i������0��,E�� 	�����Ѧ5�`Y�s��x��ƨ*��mKā�+����$Z��j̗�~!�R�&�.(%<@2BE�3�r��W�ȡ$an�nZIB�P�U� �I�����9�$L�B��pH�>_Ԫ�Zf�'��X�T�ȢZ2`���	�x���eX�Yk� �E��(�T���i���Ak�@�|�P���%��S�O+}R F�K4�d����l
�=�+����O�Q���ۥ1<�P3 �Ȥ\���	 #ܤ�ܡrB+x�d4����=�D�����.�2��'NG1H���Ƀk4ONHsҎ�*���8pK�Q5����P�P�T�F X꒴�q���/�!A�O�O�RN��D^mY�w1(%c/C�c?���6�]��@�"�b(<	��.����o��z*���4M�`�Ⱥ�OJ^�r����M���2���
����o:{.���h�$j��T2�B��%��lYEL�|��ȫ�ϟʈ�ʰ��6S��ꗆ��8��H�L	�u�yxSe�.hJ���o͵͘Ȋ0�چ5V���O>oҮ>I�|�kG#�NE�	D��Qe�]=݈��9bJ&o��t�*��P瑻?�,���`ĩ�<�['��q�ӳJnB���)� �x����iV�, a�Ӭq��"����Ip��&[�D9x���N��4��8�G
A�SJ�p��e�91>��JbĪ,��0)h��O�!��ك.��i�DXj�7��v�-�	����� ��5k�%����	��8d���w�X�RW��:6�2�a��O�(_4�y�'�Hh�1-B�������1R�J��D�&顉~�	?�I��I�RG��
��ؙU˼��Ǟ,VV��D��/0D���OTi�#�S�l��0Y���B@��"O踨�L�6
��r�\�[��Ȱ"O�(���	*�#S�[\��"ON8Y�&�2�NZY��yB�J��y�Ėe<z�鄬]�~.��a�`Қ�y�)F=2dj$�Tg�.H	�f`��y2�O¸���_8l`�&���y��dZ�t�Q̄5=@v-h�@ڃ�y����`:`-yuj�yD"5��o�y�$P-m��8�dlP�qg�  F��yB%�l�s ŷ?oԭ����ybD�v����1�H8�j<%��"�y���/Z�!�iَ$a@l��ǀ�y F-G2��&E l����� �y�'�$�&��G�clap���y���+n<����$B���%B
�ymM�LD+�&��	��qĚ��y���(}��bJPz.|�k�ɘ�y�&Bo`ĕ�S`��^��˰�@!�y��h�p(x�
�N hP���yB�9y���∂vs��[��_��y�d�'=,Jp@Ţ�5Z��K�+�y�g�4.Z�`��ْ]�����h�1�y��ɒO"�}�r+R�f;��K�@ҋ�y⮖3������6[��mr7DB��y�/F`^����#� �J��y�b�)����q�ʉ0+��:gD<�y�'�[���#a�y��d��	�y2ƕ.pb���SOH�� U�� ��y�ϋ0 ��K�9���b�(�0�y��6dq#��;{�~��d�&�y��edD��r	�d��(�ǝ�y�,�*���[�'D3X+<�AuN�*�yBF�q�}S5�PQ��}���[�y��0z���d�݉*���y���\c�����6KJ�Z��3�yr-�]�¥���
P4��S���yr��=��+�dZ
5�A!�l�;�y��ͤg䐩��j�'xx̉1t���yBś=:Ւ�V:F���/��yr!��2�i  �� �҄�' pZB��1İ1��Bɐ-׺�GH�D�B�	�s���r���+M����#N4B�	��4(b���M��$;��	'n��B�:l��]	'A?��|)�.�OU�B��4 |�ݱsD���3M�a|�C�ɞg�Z�x�Y�.�b�)0ŏ��C䉎c'~T*����y�Z,����W�<B�ɫ8f��AJ��+��)H��ޫB�C�	�t��Q�pgܡ;�mǈ�_��C�I�3'V�yj�DI�e
�	JC�	�B�$��F#�N��e�A��`t
C�I�.��X�����-���d�B�*�Y[���9>f�H��j��B^lC����X#�A�[4��
DO�3+DC�I�L�9gVu��SyII�"Or� h��C�i�%i��6�E��"OFm��j !��q��E:bm��"O� ��pu��I�`�8V�o�轒�"ON�����N���hq�_l� �;�"O���vŃ�K����bdD��|�W"Ot����Ƿx����$\��J�j�"O�y[f��:}) q��TNO�d9�"Or Qbb�m�e+F�(5t�`"O�������:�6�H &���p��"OZ��E Kޢ�2u�����3W"O5{ql$s��x�E۱Tr}"O��`"Y�LD�yWb�a\�x"OJ	���T%uH��!��97��ʅ"OH ����7D<^��W���NE��c "O"��l�1`�����B�p¤�qs"O:����������˒=$i($�U"Ol��jǋVk��"G�AJ� ��"O��	Qf��~�PIԞ ;�1"O����nF/�,�Gh�hI�u��"O�U�'@�:1����hܭd*�Q"O��f��%��#�!3Vj�"O��q�@��f�
����MF�H�;"O�р�:2� �` ۜ*�D�+�"O,���=qZ���%@8Gy�X�#"O`ȁr���إ���^��z3�"O~t�`"�wI���Ϙu��ă2"O�Q�Ƣ��\k2�A,%/����"O❉��عZ�xpb+���,0��"O����^+q��ً7�װSTJ]��"O}���E��Z�H�fW��
�"O,�;��&R֡�`FU�WY�,""O �g�D��Pj�E?*z�"O��il��9�);��E�A(~LH#"Ot�Fҕ@Y
���d:0Z5"O@�1�l%]�)����vٜQ�t"O��k�l�>-� ��R�R�I3"O�99���T¢��3��J�x�
�*O�Q�H*dЁ�^XR,c�'0���Hþ�*xQ� /I:`�x�'�ɒ'��p�8�e��C+`�j�'h���e�"2�@A;���<(0	�'d�r`���*+��@�I�y�@�	�'�i�D�	|�"� 	J�,���'n���Ì�<�LCvi��E��,Q
�'ߘ�q�í�.��ɱ?0<0	�'p��4f ѩ����7��Y��'�bBT�O4^nU�!�5$�Xe@�'UM��-M�r��X��(!*آ�'�D�+B��T��O[fN��A�'8�PR*�
y�]��V�n�J�'Tx���̛�T̈��f�n�[�'�H\c���:h~ٛ"b�P�P�
�'N��sÌ�Q���"�N$XP�1	�'�Jx�D�
J^R,��e�	�\���'�\����RQ�ec˅s�"LY�'c�-��
A�>;f�����*�)

�'��0�OB�tfP�����)
�'P�r�#T&]l�a)aA�y����	�'�XQ�F��b���ʐ˜8g�p19�'��q�/U
O�H�Z�HA�O��C	�'��]�/T�/

�f��l[ ��' JL��	[FI��nN�ta�'�H�A�FI�0��4Q�h�	�p��'��i��\h��g�Δ��'a��r�e�� ���e*���a �'a�Q�
	�0�
 D엦}E&tJ��� �[g��'lu�(ʸژd D"Oh�qBF�����}�,�8"O6�P�X�wè,*�Z/��X��"O��d�/_�����Yp5,D�%"O�dn	� �z�r��R(%W��@G"O C�ƅ'r�t�JCY-R�
�؆"Oj���G�?t2�UY4*�f��� "OB�Z�eژ	�J܋f� ��(�"O��J�,�De�@D^�!��t�5"O�����j���qQI	�]�"O\d� ���q�
;�Z!"O�m�7����*"(^1<���"O��FΕuV<lA%��c|�t��"O̅�Qeۑ4$`I�G�#C6����"O���Ɗ=����F�u��!"O�92��,*qKB��Do.`�A"O�q�CD����C9�T�G"OT��7��(S�8e���$R8�	B"O����	�=�*%�ƌ�49rqKp"O�%4
P������Φ}8!�%"Oj����;~b�c�MF;�޼  "O�b�-��m��x��k�Zz��6"O��W�*C@�
�ik^���"O�Ż���Q�^	�媀6`T�xR�"O̭@�M#mȹK�)Y8��j�"OT�(��Ț=�Պ�ûR;���"OF�3�Gɥ\Qx��v�H�T���"O8�G@� �������N�pM2"Oֵ��MB�C��a��_4exbɋd"O����� ~�X�%�ؑBg"O��$�ؚF���PF	��<@�"O��%�ђw5�
&�8^�L��c"O
\K��[s�Z����. 0�5aq"O@�ٱ���NH�hŊ�Z�B�"O�ɁK:Xe�F��̱�"��y"�̱^���� �t(��:�����y2�Z��J�6I�V+²A�"���'sX݂7jW?C�&�����H��]��'�������$v>�C��D����	�'�J��� o -����K4"�9	�'��BԢ�4&6����<i�6���'?��ӵX|)�B	S�6�N8��'l���J���ii��/妠�'��!��%Ӎ9��
��W���a��'	�I#J�d9�<IT�T!XPk�'�x!�L*:�š2��s�>��
�'�j����T�Jz��5�ʻG����
�'x��rE�>D\ �(E�����'�:=�2,�[���"t'ݎ8Zbh��'�u�ר
>ƍ�p���5���j	�'z �iE#��<��ͫ0���%�\T��'J��mB�a�,x���5y�'�&��TJ� lD�XDEMP��M��'MFE��L�:
F�и� זP�Z��
�'������Ol@��`�\�Yߔ�?D�<J5/D�RT����f@&����C5D���BZ��m�"�̔GT�qi��3D� ��Ң{�U���
F����K2D� +%�)f�r@��$��	8A�1D� �S�ыgP�<p��I72�NM�t� D�����G��X���#�e��-D�Ēb�%,|x�Ն�uY��{�+D��ƃ�#�:�"��5F���4�+D��v��8�ЮI�R��g�(D�� P݁��SԠ����8H��Aa�"O��Jiߒ-�P+"����P�"O��x��JB�[UM��Jd$"O��b��ӱTxhA�
�y~�+%"O,4@`��#�����1b��c"O�,+� �)w_ a��,:�!�""O��i%'Ռ
�m��L��	�R"OFP��e��MPp�p���A"O����-�&Aè�R�)��V��jP"O���&gQ�K��32hC*b�t��"Ol ����\v�J�ȑ8���!&"O��IE�S�kC�$R��+hj)��"O<�rWcĖA� ��3���p�P41�"OlL���$Ss2`eC1T���Z"O�,���F�b�` > �$;W"O�a���ĺ�Q����}�N@�"O<̐t�ͻh7��EАn�J��"O� j�cJe(4#2cV'2��l[Q"O�(��CSH8t�JL��a��'"O	#H߈G��z�L־B��3"O�$��I�� OP�b-�$CǶ�$"O��+�DA�+���jLP'��9�e"OY��JJ�\��٠���i�+w"O�ف�AĀp�xDWm }�r��!"Ol|B7$�'$5��BY��Ʉ"O<E��cA�RИ�a�ᘁt\d
�"O �2�ҝv���+5�.���I�"O��Ҥ�n��D!�(��Q-����"O&B"�Q.��yygG�95c��C"O(�K1�ڢ/����`РE7b�Y�"O։pwO�r~����oH�V;h*p"O����k�1=[n����,����"O�����#3	��[����=����"O�H���ن���e
�=Z\��"O�T8p�x�,��vd�!i<,��"O�9ZDS��ҽT�V�&�ԑ^�!�ت!��0#v���g�������`T!�#i�DБsgѠ#0��B�/�LH!�DQ�VQ��k�I��(�@cӬ0h!�M�
���6D�8h&Q���?#k!�ל�r!Ԅ֓]�!r�'2l!�QH�`�Q�ERt7���G�<T!� �d����7d�,��t*#F�(�!�DZ�P: ]
W��u�p�C���h�!�$-X�6U ``�a�س���!��ơ�	��,��g�8�a�g�!�$d�c��*)��h�=6LT��'�F���H1�XAs���;8��[�'�6-��V%�h0��O�?7����'ں<�á�z>ФÑE�[�(T�'���J���6!���o�o�&���'��<	�%��`f����g��f��q�'kT��'�����!a�G(��͙
�'�Εp��<cd2�[q��>+����'����Q��e�z=ѷBN�=i�!��'E��p�%EmR`� ��5G<0��'@�	�����X��(ԃ)�.��'�"�)��W�V�(@�L�"�(��
�'�q�Uɕ<P�h�W����+
�'$�P��ӌfx�+���e7�M�ȓYSڔ"䦞�w[ؼ�LИQ
�ȓaD�,3���d����ȓ<�2���!cK� �N�-�Q�ȓR-�Mk�j�Y߬�/%�2i��S�? ��-V=+t(0@�>���1"O,���˗�0ڤ� KԤB���"O�mABЧEKzm�&�S�m��ź"OXT�U��).5���$N qt�t�U"O���7�\=>�=�ROD����"O�,A�ذ|�D�*A�!}#��P5"O��a�.ˊvԲ�C��&)��B�"O�T�C��Br|@ۤ�Zy� 1"Ol9bbnP`��@��$F��mR"O���!��^ ���6�L����q"ON�
�M'�����ܢU�&H�q"O�}�"���{f@����&޼�÷"OX}R��&�j� o�*u�R`��"O<�� jE,N���d���a�
a�&"OJ��Q	�	Gg�	���@*Q��(�"O��B6�E-��rF �
P���c�"O�p+ǒe�h��`��~�(T�5"OnP �� C�Uꑡ�� M��"OzI�"F�"6pXq@-!5\��"Oh(�PcZ���y�bB��H�(�"Ox��4]��d�Cŭ8Q�q"O�pGU�m�Z�у"Խ)=�x:s"O��Z��0-y�<Z��D�-��`"O�������Ћ!�F������"O)R�
�0O0"�B	>a��K�"OH�6E+F��a�b �;���d"O��a3��&$Ж����>2l��ۓ"OJ���■'��<9�Ε?:P���"O�����)d �+P��]����"O�Y����4/����!\uCf%�W"O��
T�@:&..@0���1�Er�"O�L	��ʨ*DN�h�N�<g8��S#"O��3'�[�,��CάH��(�"O����	ېC�츉U�߈Ғ�Yc"O�YkV�5B ������JÑ"O2�ʳN@�sQ���g�9ȌpÂ�'K�M��$LcH�Y1raםr��E3S�2M���R5,fzE`I>�B,T�,gxAh	�'>T����4�,�P��
X^2 �'҈��c2_+ɧ(���C��8���U���a��c6�'�Rl���[4ɧ��x�H�Ƅ�w��%0�lúm�޹��toNlq��|����L�:m�ܽ��O�"UH�D�{f+	�'����0➳[H
6�L����?�aҟ(����X?�ZH�5JůT�|R�iގ������B堎!�̥��-&K*��\�D�`�K�RT�ˤ�V%��lT�&��$!ua9L;�>��'V+���9^׺H��)�\�I��x��7�˴�p���`�t�,O�O�4, �")���Z���Y�B�N�0���)�S�Ro���X	!Ʊ_��A�칟�x�)ڧZ_�)�č5<�4�jW�ՂQ��m����R���>�`fj���P���X�D�!�>A+O�$��?Aa�fO��Hc��)��UIEj��4s��#,L����RZf/ڧz_ҝ�"�N������ �Va��AB��O���	U韴b���0|"Vƚ>,�K�.��Tz�M�M��<]?0!�?�~��O�O�"��$��V��0rQNKC}�]�1��|��Fjl(AlN�P��T UR�y"gȑ%-�P���_�p'�K��yҪ�/;� �@@.Z�k�����W��y�b�� �A�`��sE)G�yBḡѴ���לc�"Ls����p?��O�y�,)W^�M�p,[/V���r"Od�U�uq���l�
��C�"O8ӣ@�[��d0�KȮ �R@�D"O�$�p��/'n��R `��d9�"O��!���33�t�.	 ��삧"O<�	uEM�m?.�s�γ@@����"O&@Ȇ���ҽ*#�M"'����"O� �
��Ă66��Y��+�Qc"O�	���<*� ��J��[\*8 �"O�5�VF�x=��*��P'}Fx��"O���ç��+�&,�4�=�}p�"O~��CXz�����R[Q%�7"O�Q2g�?oeD��r�#�2,�"O(�aDC��,��ZQDI�$xީ�V"O���w-ų~�4�Fن'B>�3"O�q g
0�R9��31z��u"O���S����,h�%�]�D��&"Or	q���%fI���cّ{����"O�Ҡ�B�������<�P�ȓ6^�HHc�*��H����Z�4���HtN}`ʝ1g��P!�V�M�ȓI#"�I4-ORް��햹�z���*,朁!B�-au���r�\�L�씆�>�xb%OE3/ �{#��"��t�ȓ2*��ᴈ�^�̐+�g��&X���id(I� Ѷ���H������J��DI��SJ.��kz>p���8��W��`:�mQ	j�B剢GY�t�b9�쌑���	,�C�I�;�9jI� !��Q�%4�C�	=;�b�x� "��Q�mB�D�|C�I-ٺD��d0�Pd��2� �P"O6!
�c�rz`�%c�-��@1"O�IQdI�r+`5Z�k<8a�X��"O<�(��@�E����=v/�*�"O���p�z��,c=EftPd"O�Ⱥv S }�Vh���Z�{?�"G"Oث�M�2O,��Y�����`���"OBh���6�z�xQ�ߗ5�� B`"O>�A#�7��	3"�ë1!T���"OdM����Ĝ�@�ڟ#α�"O�tR��T4Ȱ��7�S"O���I�&+TyXv�ϐF$D[q"O�K��ƤqԄ��dQ2g��*#"O=r��T�utN� �K7d���E"O|ȓF��<oj�4s0nȾ`��@H1"O�@%d J�4�C4�\UH&c�"ON�R�L�`�d����(o+��!�"O�)��gA>��f��$��:&"O`��cV�Z�R-�_�2d��"O� ���ĝS
`�"��VCB�C"O� z�����X��JS
/�=��"Oް��FGl.��H�r4\���"O�qh!�9 4va��f��x�༫F"O�I��ڝu�~���eM��"��P"O�ق�U'�x�+D9qQn��P"O�9;��	&bV�sC��1<�\#B"O�+`�
|\��T)��2�Dݺ�"Oz���i�iI\�A��;_���B"O�EI���&L�'ɛ?wS<Q�#"O�Mkdnݘ>���QǊ?aO`(ȡ"O\ajB��v���R#�8Xu�"O��0WL^	-M�&�K=kȰ�"�"O�d�B
Ĭ �1����$U��5"O���(Ȥ[����)�+�|���"O�<���ѪM���pP��#oD��F"O(�'��[��q"�C�+Z�"O��JBID?Gb�ӑ��19��	�"O<%*�IӾ$%���b�� ��5B�"Or݀��ٴ
��t;�T�Ppte�s"O�y� J>:��b����r��U"O� T|�3*Rd�*����u���T"Od�Y2â$����ϗ�]�j��"O8��''�v��Q ��.%�*�"O$�"�ɄB�~��#d)��i�"O򴚓�E�e�@���Q�[&j[F"Oޤ��Γ�@4��ð��-��C�"O
��]k� ���IB"O��9%D/;��݀��ۻF�H�xB�D.�S�$m��m9�'H7D�:�H�AT���B�	�(���E�ɮ%�.�A5J�%d�=IǓN�h�h��ܰ����\nC�f5&����2���XT�\�V�\��T2��/\N���V>����5�O0O�Y	���'�~$�I�5�.MR�"O�L�Ŝrsl	��Q7L�DɅ�v���)
�[R�ͫ(���b�nԽ[�!��^����ZL�]��l�4��)�^بP)0��<r�i���Vb����'V��A��')7*x��/T�^�	�'?P�'%�S�LE
eǇR�h�'!؄��G�8���QD��h��'Ѹ�*���:��8���܁>�<�9
�'ߤ��7��F���E�IfT�Y

�'y�QEA�!�
Ҁĝf��<�	�'z�Zp� �K��P�O��	�y[
�'���r���)s�z�#QE�?<l�z�'�����t	X�r �Z�Uq�'�޸�v��'rC^!�aR"��P�'�>A�wM@��0q�bP˼�B�'v�U�Q�ny�I2R*�>谸�'lH��!�aMd�"�@O�+�`���'�~
�ͱLA�UĂE�!<�Hk�'��$)���F{��3�Β1}\M�	�'�
��!��N.=ɢ�K���ԁ	�'�| D,HD�F�~9����'޶y�D�[� Ӷx �H�t�&�"�'I�YI�Ζ:���z�f�7g���a�'�(2pL��cv�,b�%������'�h�QG��4و���"U<?��,X�'=,�%�Z�N�
5���8e���'wȑ���Q�vu��	�1�R ��'�D�f��+V�*�+rnR�"Bi�
�'��A�\�m�¬Q��T)��1�
�'���RG�:@�5;����"�@�K�'�d0�"R�f�
� cU�M�*���'�y��o]+o��:jY+{z���'�I�weҖH�I#�r���'���ö"�8`ڒ�/�,	Y�'RVUȥK��r����R��� h5��'����ꀱ#*���D)�q��'���P%Ɋh��!"	���~�:�'ܔLB�
]�g`u0�[�t��`�'M,�q�l��^�5���ۙg�<z�'�TT[�E.%�h|�O�_lv�`�'z܉1�m�/]��@6샭\nbp3�'��˂+�
a*P3e��8S��8��'���"^2��+F�I}�	�'�R( C���wAE�Q�t��'\�X�k�%R�N���dY9D�N8��'R�����]�;�A�և= �e �'�2�I&b0�$�!Q�F�*�(��'XB��G���d�5i�ֈ�d9�'�=���X$�����a&�	�'� ��A�� �g�]�:U���� T��h[�	��2'AG�Ċ�"Oh�0�J�~��kAi�"K�hqP"O�(x�
h��ث��2��]�a"O��b5�ZM�T��A�;o�"��d"O���OA�8��+�e����"O��U��e�� �do$��"OR��DgA�T_e+U��l޴qR"O��R��K$p9f��AI��~L��
e"O<�B�o�+m�|<�7�B��jW"O�P��W8`YȀ��E�v\Lq`�"Oa(�*Z� �:�TI]�mQ��* "O"LA��'`<��P�@D �r4"O`���S�Ej�(d�d4�9�"O���,�j�)Z��ִ�b"O�|&ǁ�1*���M�D�M�$"O�@�@�.l@@����>- ��"OȘx��OI��M��c�]
����ybeY6*�D�t-O�L�ʼH�-�?�y��� =h�J�H�$2��2Ūߝ�y"�V��\s�Iڔ3E��H�Ð �y�W8s[ڝ�!�58�#����y����ةXf��!5�Z� Rτ��y��т6�(p�m�5�6ݣ̜�y�M��AlT��EW!��1� M7�y�`�9�
2%��b�Z�cD.��y򧉐�j]���/5\��!�y҄�H0�M
��'�^5������y2��82�q(�k�6��K�JW��y�/ڰ~�PK�-��:�|y�G�͏�yRC�!`�s��C`�H���y��Ւ�~9�F�Z*����^?�yr ��HF|x�")�+N�}#�B䉄 9^��&�D>J&TL��d��7��B�I*%
V��G�C8��A����%g�C�	��ZX:ȅ=g���!AN�ppB䉁
k�h0����� ��R�%CdB�ɐ(+�X��J�;�����*GP�C��=B8h���T(𢘙 �!$�C�I�"���͕�r�Fd2`� �B�q���0��7!2X�fi��$B䉔�t� �"�a0*L�ի�"B�ɏn�hm��	)sN��0����M1�C䉻����P!r䅣���1e��C��k����1��$9���ʆ �2M%�C䉈5NX�I6��Ap�Ab�U.��C�IM�A�BB7p0j���E��B�ɑՀ�J%��&r�义���Q��B�i� �%K�#9y���U�юB�ɽO  �Y2GH��f��Tʓ'~�XB�	>LG��"bf���pP!�ύ�.B�	WK���e� �n=,��vI4B�IK���#��p�ji���ȌE��C�I�+��kt��#IX�H� �'2P~B�	�#�4�YQEW�bݔ�R��kǊB�I[��E[�2<�$�:�C�28�C�O�\8���ӕ7V��럩:��C�j�z�@L�.s|�"�^"�B�I �4��W킊|̀��SݾQ �C�	1TRX�E�O�h�QŜ_�C䉩j�|�"o� E�f��F��u2`C��0�S�Dcd�z6D�Zn�C�Ɍ��!`��uڞ!��!ʹB�	�0�`MC����$?v�>"Q�B䉞^�Ȕ��1(2`�$h��?͒B�)� ��&LX*Z-l�P5C�$����1"OZ\E   ��   T  >  �  �   y,  7  vB  ?M  sW  fa  Wm  �u  3|  ��  ��  A�  ��  ƛ  	�  M�  ��  Ҵ  �  Y�  ��  ��  !�  ��  P�  �  ��  ��  ��   � �  _! �' �-  Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�� |d��"O
`�(�;���8���-0��1%"Oj4��ND^[��"3/9�0|H�"OB���H��*�ʞRy=a"O�味V�!X��!&F�:J�$���"O,��a
���C�Ą�M�"O,$3%o�-���p���+Ն�:1"O��ݢ1����`���y14]2��i�<�6��{_���c�H�`�fX�$Kn�<��A̼VI�xR[�)�Ć�pඤ�ȓA5��('nߡ4�� �)˩%� ���,��r�؊b#`T�eT09���ȓ!�b��g��}�8�F��-? �ȓ
K|m�ș�VṔ���2�%�ȓ"R�X�j�4JN�1�˘X�i����̹	_�jZ��1!g��zܶ��ȓgil,*�J�
j�Ne��i�J%b���f	�(U��:���G��$Y^م�~r�� S�%T"���k\�jx�ȓ|4�1�îJb��@ӵ�ݩn�V��/[`�"�v4�R�!ʎ<��M�ȓ`:��z�ؚh�J�Z��$HY:	��H��p�m�C1��!��B:��0��EnjZA V;9����J[
2���	��4'J�EA�IVW&��~�(aZ��ӹ�>� o�Y�|�ȓ�f�A�
Ο7�H��M�$�����mޠP����/���ANXo*�ȓTv�����{ ��-7�*h��I��sB�8�8���3����ȓNe*M�悡;������X�o��!�ȓ'lj�#F�m�+R&;�|��2)n�C��0S4���T:
b��|�O���;�'t�4,`v�K)�����Nk� ��+:�Zwd�gIv�:�OD��|\�ȓm�@ � Z�n��=�䢜5P^ȕ�>9������C�z!�1��ϫ>��!ҙ�y���pE����J;@<b�Q�A;�y,֕~�詑s�d�� ��'��y�i�6���.�	�I&�A.�Ң=�;�hO��T�W�{�h��/W\}z�6���'�q�"Y�3G-LJ��1��W�|�6()�"O�)23��5�ڄ�p.�3{��[��'����\���0�E�
���V?f%��}< ɓ�d:�r�$�)�8�r&b�'y*"��R�D/v���@^?z
	#� [XC�2m�D��#ޅLؐ��p鎹kR<$ϓ�~��퓟(�	�S�٧qFRC�� �V�IH������W�qJ���h\$]�p4L��'�a}�,�*�a���V��<�tM�<�p?��Osd ��9Dp4�5.�.{�zB��|�'�~�86l(1�,8��Ύk�(���'81O�u�|rL~Za�%�lm�_���/U?p��C�I�Cw�xY"*�GN�qJ�'���˓�hOQ>A�%'%�x�P�K$!{<�9B;D�Dz0l�^�j�4�ڵV^��DW$���"��?�HI�jݍY�����(%���f�<���L_��:p욫,�$�⋈6~�R��0?y��!`p�TZ�g�B"�h��{�<y ��,E�`b�㉙-}F512��k����'�:�Ѡ�6%j`�i��9U^hS�'OqOX��d��_9Xd"Q)��FǖiEL�;&�!�� \��q�W.fk��Z;2��(w"O�Y�t�X��"�!� ^�����'��V�!IG(��I?!�T���j)D��A�H�X���'fG&�.]�
"D���kI
T�v̒ab�K�6�#�O>扔	Z�L��LG-k��a���1X� ��V��h��`�ɡy�!2�N��pxXD0��'J�O t��AG*d}��9���<?�ɻ�"O$�4.Ư�^��^�,*@���'�qO�!sk�:J��qx�O Ud!��V�܇�	YRXjWA�*�\�m1g>`�<a˓�Bx��nH?ŀ�f�5WX�5���F?��	�<!:�Sbb�)y�� �o�[��B≊+�FQ2�R5h��b���4C�	�6�̡:��C/:n�����,cVC䉂iX ��@&U���v��;,(�0>��4%s�`�rB��� � �@!Q���ȓH�hp�A��uL`ȐFY���4��C�4a�"c�V��ٻDN:/�,�ȓ?|�i�E���д� �A�~;\8�<�����01��� N��u�
�
��˳O�qO�����L�O�ԭ@�{������rD���Ѵi�8��	#��lQ3�>o��A��(=XJ�<���;�$�.kpC�`#Y��H�yb�ʿ.���H�b�Hb���oA���+���>}�V̉�>NlJ�	æ����<D�Lr�H�=(��sI^JOHi�CF:��<y.�y*z9Hv������e�<qn��q��T��\)9<��F�L�b��"~�s��YS�C�� G����\	�2��)�����[6`�!@��,�X隷�.D��S��J4ν��`қT���`@���hO?���=3�`�����d��ȃE'�;�!�$U%!0в$��*� ��"$Cd�!�D�Yڮ$ȷNA��X���E�'9�zb�V=���{-�>W��i�6��zL!��],���3� 8��y�&o-�	�<YW��O4�S�4����S�N���&��@��CQ�<!�F�' fU�ll�(#�+*�@X[t��	t������G}� ��h k`��o�~��� �yR��2���`��C(`H��,���y��&	LY�B>�Y��k[��y��\Ψ��੄�{B��������ybJ�2B�p��I$xJE��O� �y����T����̡"��eK��/�y�!9�~�17 ��iv�A�M3Ǔ��'I�R�(M06�1c����%�y��Y6{C8��1-�0"I� 閧��'�ў����j!f�q��O[-	�c&"O Hj��۳Zdz�YQ�Wj� 9Q�O��:�oL��ˆ�&l�D� ��Mnp�Ey��Dܖ��)�]x���S�TS_��c$�ҋ%H�5�O��Q�&� i��1���9���4�IQ���PCΉ�C��Le:%��+a�!�$F�R�~��(~��5ԉ��#�fp�ɖdQ�"~�d@��0�9k���#
�		��4�y
çu�.���+� 3eJ�RE`��y�A��Du�92x`���͈��=1�y�`���a��Zy�b+��y�	�&z\l�r"_vT`8"b�B��hO,`D�4��:��=:��%�����y2!���sHM�t��D�PA2�M���)�禝I��8
v��	�4g��]F*(D�����M�:D}���/8Д���>��S�? �4p�H�We��ys/_�'S��Q�'�1O@���GE= `�:��'1JȕQU"O�	c�����@P�+E��|�>	��I�7o[�\�/ξ\�\5Ȳ��|'!�Ă�e�} M�8xje��d�7U<!�A5ʞp�R��i��t�3$
�9%!�d��s1�4�*nڎ�q��"��;'OxH1�U�蜸E��7)�qҰ�'���:	�!z��P7'�]�h�r(C��RJzУ6���E��2.� *C�ɢ5P��`E��*�9���&��"?���	�!�ѱ�eI|4@ic��Rl!�d��m�d��D��Fŉ����8Q�Ix���佸�T�!|<X���b���v&"���"|�'w���D@�c��};��� .|J>!�^s��aG�'��MQ׉�L��I�բ��Ď#��Jѩ�G0�{�f��!��\�We<��d菞5Q�lЀ��E�|��x�`۪`r��S�xT�qB�ڥ�yB�0��P"0�׹���g��y�D)*�t1S0�.y����#��1�S�O("x�E�1*�|�aQiַQ��01�'��u"��*�� �P��{�"ݡ�'��y�ꘓa�Hi�G yN����'ab!ıY�n�X�jN�j���W*_�p<��O<�'������-q���t�`Êy�����
���@��h9uBރV�E"��O��=E�"�I�h�'�Ȑ|���5hE�^V&l	J�8���]�˦j�uu�����p���OD%�=I��d����샵���"=���@@�	1!��I,DXG݂~!D�2N�Q�F�To��m�ܩS%�\���&O����x���7�X��uK��6vy��L	�K����>��'�2��i�'*Q.e˃=�P))d���!��*=I�cΒ���ȋ�!��Z*A\�@��Y�d���b�U�)�!�"8�Z���fK�N��|��&Ia�!��G$�|��O3�a�0慐\_!���#�؜	��g|@ydG��!�2$�x��a��K�]`g,�t !�
�)i&�Y�� �lB��".�3)�!�Dd$�����ζb@ܥWo�!a�!�$ɀl����-JR���5��r�!�,zԈ
Gܽ�*0퉏n�!����
�t���E�r���-�&�!�D:�l�f?P�HD��,2�!�$�	c~ ���I/
�D5hb	�n�!�Y��`L��o�9v4��D�D�h�!��@�XTR4KKd<�C�Ou!�dΚ��ġ�S#�ɨ�uu!�D�6,���0�[qCN97n!�ǝOR����Gä+�	���z����i�t�c�.���<1�P�ȓ��S��=_fq{4m;R2�i�����cD�_������.Za��]\p���l��3���s$�,:�V��A��h���[��[��߂0�j���Y��06dG�++��%�X�@ *���.�!f-�q��@�%:ir �ȓ=[�0��M�?_�p!Ʈ�2Fô�ȓ�<�Iw�A�d04��Y,/�X�ȓህ�Z�!�<C���%,걄�K�����K�$�ؑ�$T��l�ȓ��8���m��a	!B�8���S�? \E;Ǆ���k'��Ci�	W"O|e`�FJ�b�s�D��Sx2j�"O�lq��U��Y�c�b9fY��"O�(0r	66�����<&��5"O�(@� GN�� EI�4Z<|��'��'��'#b�'�b�'��'P6���Z�*Af�*��E�!�,��'�b�'���'J��'���'*B�'������G9��ؖ�����Q��'��'��'N�'�'���'JB��"�Y0T=�	��h�&Ղ����'$��'y�'?��'J�'���'8N`��C���)�$���dB��'"�'��'e��')r�'���'"Q�@f�9l�P!�� I�.1�U���'v��'��'�"�'�B�'��';�4��ͳ0�@$�3":P�A�'t"�'s��'���'�B�'���'�� ��O�Z�l3��:�5i"�',B�'wR�'[2�'���'A2�'o�`��dH(��p�"H�2ٴ��E�'�B�'��'"�'���'���'� �2�-�H&�I0@�
�]�2���'�"�'���'�2�'�R�'U��'( �
bv֨XJ�JK�Mb@���'��'�r�'���'���'h2�'|�z$��9���Hր TD�b�'��'�R�'���'�r�'
��'����±Z%�� $	T?f�	W�'_��'�2�'���'��"t�L���O:����D���$��D��9�<	��]zy��'��)�3?�ưi،tH�&�\�J����ϻK�2��ș��E����	z�i>�	��M��� �n:�g��H�M�,ޛ��' `-2-���y"�'�$�B�ȇ����O2�*���;D��&�w�u:q��O�˓�h��I��m�O5�d�FNSc��T�1C�&�I{�'қ�w
h��)W�$���B�hʈ]��Y+��fӶ�n��<��O1�����A9k��W�w����#mY:�J��Ȕ� �󤛍n�fm�ChT�5�N�=ͧ�?����Q�rP*�ݛ��D����<-O �O<anZ� ��b�(`'%X�;J���s�F:�K0��B�x��I�M��i5�$�>1���i�4���ǁ��J�Q�hF~B叫,���0����O����S�ц>�r��</"BE�æȒ�t��`F�3��I[y�𧈟�$�����!�U!�� � ŷP��D�٦9@m$?�żi��O�IU�R�̼�eJ�UF��J]�'A�ĔۦM�4�?�V/F=J��'r�#%)N��&�[6�ļ9��aF�u\Iƈ��4r��Vw����n�`�[�H*� M4$�1"T�	G��,���$(��q�w���E��"f�>hB��l�P4Z�� ��}��kP�,@��g�@��h�����(r�L��#&�"�u���0�.;�N�-�İ���^${B�Q�c���I�L���� <�����"�`�{UL�' ��P`�Y����ޢ-�4	�%
�q�����#�DM�{Q͞;M� �����,Z@��մ�i�'�eݲI�  �XuF���	5C�|�v�H��$�ڳDhq���AB�$ ��i���'��O,��gR�bG�Hw�vŚ�LBK���lJy���O��"}�'Ǝa���D�ʥ,�{�M��n�9��F�'�"�'����3���OJ��s�E2R>N�@�U.�}{B�Aʦ�{6C�I��|�<����u%�]���&HR��v��i���'�rl�5d�F�d�'�D�JV�֡�^r���!!˺}�<��jޣ^4�O�"�'�B�B�T<@q�FK!^^���g�5m�06��O�<�#˒�Iϟ���m�i��	0H�@���r�\�N����>�%�e��?���?�/O��B�)K�E�ҩ�R�T�\Ӵ��E�L�"y�>�������<I�z��59e 5H�!=Rn������O�D�O��$�Oh��ĥ�?]yw��t����-�:uB�em�&ʓ�?QI>���?��D��R�PAl�7 ��e��"r�`3�%O�p꓆?1��?Y.O֠��B�\�ӹpaͩ��͸i,(1����!]�F��ش�?N>�/O�]�����x�Q�
�:U�f]��d�)!��'���'^�N���'��I�?�[pN@8B`��ήRs:ы  O	���?��b[`�q��w�S�$�ID�U� �z�����j��FP�Dː����Ms�Q?Y�I�?�B�O�1�!�۵ޤ	��C���e&�i9�ɇ{��#<�~:���/���p��4\((8 W"Q��q
#�����Iğ(�	�?1�'�S�Y�Ԩ�)��B������ߴJJ����^~�S�O�"D��Jt�[%�*�H|+�,� ®7��O�$�ON���D���	ߟ ����iݙ��茌g(�r��� /$����x��z�P��D��<�O2���'��茝�t�iv�ڦ�8@���A9��7��O������Ǧ)��ߟp���|�����6���`�Gؖ(�`X�1��"Z��H�L��'[R�'�B�'��(R����j��`��|gjaW	��M���?���?aV?�'���X�	�x�BF��R��S�f9�����<���?���?�����I�#�p}o� +?.��#
T�}8\|3uEʋhM\�޴�?��?����?q)O~�D�D��	E�h����dC�y�0�uRplZ��	韐�	ʟ0�Ʌg<��ٴ�?�b�R�� L(,Z�
��0Ȁ=��iz��'��\���	�x�������x�H��G�JI�0al�<~�o���������	��1�۴�?Y��?��'Z}F�F	4=P��3H��?|X�a!�i�2]���I�9<��u�i>7� xPI2Ɉ����ƙ�X�÷iHr�'�6��sga�H��O�������OlM����z������j��p��N�[}��'�K�'_�\��P��#g��]�Wʁt�]��!�
���O�7L7�O����O.����r��O*���i������u7�PHV�"�� oZ<3�����̖������'[�����a3��A�h=4���6Nw���d�O �ˌ�6�nܟ4�I����֝�kb�P�Cf��4dD$I�oڦ#�N7��O�ʓM�,�S���'���'c��*�[*=�	1��W��.��t�o�p�$�R��n���D�I̟��I���ɽ���B�-Mn��r0N��N�0�Ҧ�>�t���<q��?����?������a��)���	<���
M�v*�@Ҧu�	�������@H��.ʓ�?	��%$��$��/&[+������@l�HΓ�?��n�m`���?����?Ig�A�4o���:q�bbi:(x+߾d9�7m�O���OB��O(ʓ�?�D���|�P�y�\�����7�z}u���?��'"�'���'�⢗ ��7�O��$�;^$�rU�S82�~ ���M�?� n�ܟ0��ϟH�'r�B�=��T�>� �T"�\�ҵϛ�R`<�iK���-����|��矼	a�O�M{���?�������Z�m��42�ȃ���Y�� ����'��ʟ��v�h>���Ay��Mc����r�45icJS��Y��+�⦕��柼�Z��MC���?��������?�bm��.� �j^:R�$�	V��Iɟ�!�ɘ����	ןh���b>���������!v�uRa`�_�d �"�iZ�K�B}�(���O���������O��D�O��Cu�\!��@�F��4�0}�A���)y��֟���fy�O[�OW���Wޙ�х��{�rе��i�P7��O����O�%Jԭ�ꦕ������T�i��x�i�>t~H�#�أe���(��q�"���O��C�I�M��?-�ٟ��I�UG�II�Xz9Qf�̻+c���4�?)v��,[��	YyB�'��Iٟ��*'`R5� N�Tc�G}�6�?U���G>OF������?)OV�4Y���Vȋ�y	f� 7�\9`��'V�I៌�'W"�'��፰"����"��U)$u�w@�CCЌɚ'"�I�^{�l������	ʟ�[��Ϊ�M��\*2��ȥ��F��H���ߵu���'���'���''�	���y�p>����-�$9�J��a�+I����Oh���O���O�D��Xͦ��	�����79c��0ӭ&�z-3&�X��M���?�����OVU"�=�n����*"�A�?�L�z�
¥O�Sa-p����OZ���O�ݹ�D�æ�I����?	b�K�\�а�%$]N��4�P�_�M+�����O�p�;���O���ZƐH����@0�SIʤ�M���?i���r���'k��'��d�O��	F-W2���Ȑx��͊ HJ�����?a'�ٟ�?�O>ͧ��Ӯ �᳢�!Yz)��Z���7��X��l�Ɵ���`���?i�I̟�I�l����s��\$��Q%!X?a  �4��	������|�J~���rw)���q�ͫ���5[�)��i���'�"�%�T7��O����OF���O�Q�B=<�i4W��%y��;z��	cybd;��4�.�d�O���P�P�0�0L���gA\� ��n�џ�����M���?y��?aW?��Vz���gH�����/`�D��'��}k�',��ݟ0�������ȟ��A��:!R��#u�\��E�C�4�ٴ�?���?!��.:��ayR�'8,|�)|�TTȗ"\Hrt���ȏ��yR[�,����(�	ퟠ��fM>���4N	�����2�y� lU�*IF\#D�iM��'wR�'�"[�����j>��sӰ%�M-��t"�dٵ1���i���'B�'~��' pMb��i<b�'����e	�+CX\�&�����V�g�~�d�O��$�<���o&��ͧ�?!�'u�|�0+HGk hJ+�*(WШ�ٴ�?Y����$V�IUnQ$>��I�?���,O�~
l��Qӧ��kE<����d�}���zI#��
@��L��L0@�moy���0��6MF[�D�'����)?��,�]���!Iܛ1��D@��a�'4��@����C=wY:lʀo�aV���A11��V�ѾJ��7-�O`���O��i~��؟$��C�"��d����'����#���M����W����dYx�Z��ǌM�$�良s:ymş�����S�O��ē�?����~b旍�u��K�=&zD�q�I��Xb�\q�%�����	��ܸƦ
GB�
f�!5��A�Z��M��� �U��x��'��|Zc���rhV2o��b��l����O��"#��O����O��N�A0Ù�l	0x�@D� d K��7d0�OR�=��<9���1:`����Z�#j�Q׎@*M�v@�<���?Q����Zq���Χx�p��D��h\�s��7#X��'2��'��'3剸j�B�qV- Tϋ�wx	���@�'v��'�R��������'W����j�B��* L�[�\�D�i~B�|"Y�x��4�I���a5��W�P03�C�(~�7�O>�ĺ<)�c^7��Og��O���xS*�3�ЃU�Gb6|�6�9�<�W�FV���IHkKb��C*B!U:`��c��&O��v]��rg�ĳ�M��Z?��I�?0�O��!P�n�L�@S#��0����i剫w�"<�~�g�m�d�Z��H?n�<ar�צQ ƃ�8�M����?q��Z�x��'((|Q��c��=b]uk�a@�5�MS�}�����D
|�?  �BNں2�nI�����
�:hk�imB�'����>jFO��$�OJ�ɋl�`
��-3�}�&��iLc��Q�%3�Iş8�I˟ppb�� �
8���}!++ɭ@�7��OzM[�~��˟��	M�i����_�$�腺��[GZ�y��k�>1���s̓�?����?�*O*�0&�۬<Hl�;��۶R$\��2#�,�&���	̟�$���O�= e#F�*��qE�"���)`�D�O>���O��<yd�iW8���Q� ܢ+F�U����<�����V�T��̟`%�PEy�l� ���2��٫R���9t�)��d�O���OJ�A2�;b���Ƶv��e��ęM�$ы׃B�k��7��O��O|��$��ZO$5�1*P4y�|�aE�%ޛ�'q2_�DQp�T��'�?i��JOj%�c�ɕ�jy	5�ܤk��x��x�'>��֮�6��-@�A5b�~p�ݴ��d/fo����I�O^��q~r"Z�u��h�m�3�X�2�#�M�,O���"�)�6|�R��5)�I��\C�!�I�H7mY?@�`�m���t�I�������'�RL��蜢��L
�*�/S�Z�pӄyH@�)�'�?�t�
�
��D��4d�J,���'J}���'���'�p����/��ڟ��#����m˩x���{G��>�N��>y�h�u̓�?	���?�[�\U �텦K�XTI%!Q�dN���'Pt��8�	���%�֘�B���`���)`�f�x�i@��c����<����?����P�+�-}�(�
��D�hh�Y��|쓹?)O>))O��Qe]�	��s`�N#d@j��AE 1OP���OZ�d�<	��a{�I�/���S��G�y@6Bz��'��|�X�,pO�>��Y	#"�,�@$*Tn|��V��h}b�'�2�'�	3N�DXM|bV��~�v�҅L� ;Z���� �����'�2R� �'�f��ϟ��r��pK�"{bRi�&�7��OT��<aA%��qe�O���O+��[��\)?\<!��o�3-9P�`G@n�Xʓ��!C�3?�矤@��4}�0\�V#ًR*�ˤ�i���q;B��شFz����,������kҘ�b�E�S4~�0�ד[w�f]�8YWB�I��|&���.ц�b��c䂀0���a�)��xI�#�̦y�	��p�	�?e�I<��z���00�ݫr
��u.�@۾��i���s���S��L�2��8n��6Bчf��D@�	:�M��?����d��x��'��O��s�J���^mÒ�G�GxD��dA)C�1O��d�O���A*%�(k�D���~�R��$n�؟x
4,�=�ē�?������S ��am�<��鐩@����ãd}�I�'���'��W��x4ƕ�=�P�9�^�"��|�!K�<6�@��K<����?qJ>�*O⢩��_�Rܘ��ܐi� 90(��1O����O&��<���^�LT��kjN��=%EHpƒ05D��̟(�IJ�Ly2�W
��������KO���GB%tu*a9T���I����qy2 ��?N���� ���Q_Z9I�#�9y��e��ͦU�Ic�IGyB	ќ��'�`�r���=3��߃�|�X��n����OR���$�ƚ���'(�ᕲj�|�Kp�?j���qh��U��O��vwjGx��։�e+x���8LۮE��8@��i���4(j��ܴ
������,��DϽ5ڐ#��O'�u+#�����fS���!E2�S�'+M�}	�/�6d�b�Bw���mZ)[����4�?����?	�'v{�O�}���C�D�R��S 
�n�PC�m
�b �S�O3�4{uV�H� �<$�h$ڞM.r7��O���O�PTɜn��?1�'����U�Y%��w
@�3"��}�@�̘'��'g"KW��8IG��t�a �^�X�H7��O���f.�v��?�O>��b�����9	�y����C��u�'���y2�'�2�'��I%Bb�Y�E�@�Z����Sa�P]�5�-���?���䓫�$�W���!�$��J�:�
�l6��z����O���O �!P�`�:�����C� ��cKR�RS�͓�_������&���'z����O�,X
�-dkt-�qJ�PH��rX���Iݟ��IPy�HВ"�H�ж0-J�	2-�i��l����qKI�E�In��Ry�&���']r�*F�9Se�19��Ih�L�X޴�?�����$�V7�'>��I�?E*��M�k+�p���_"�x��dD	����ܤ\��'m�����Y��� �%�]�©n�wy[*�7��j���'���0?���r��K�>~����ަ��'��Ir���	� *R�L3@D�"H��bw�HX�6c�nՎ6M�O��D�O���Q�	�ܑ�D�^��x���]��@z��5�Mk��_������M/%L���%G�	Rv8R$/e���n�����	�4���%���?i��~��C�0��BΌ�v� �i#�����'��@��y��'���'lz,$@�[P��G)�8h�8(��Lu� �$E�!�ب'��	ҟ���xyZc��8��L��2g`Ȏb�a��O^A����Of���Ot�M�� �����3�uR��SK��Ys`�� ω'���'QbV������U��$}ꡚG��"_�t�p�CҴ�b��������Ijy�g\6N;���7Z������TP��j΋S����?����?�-O���O�H�[?݋`B˸MÀ�4�H� a�	9�G�>��?������R#�%>�Тa�+�j��Q�F
 �@	s�%�7�M{��?A)O����OZ����?�9�z��#h˧̔�x��L�W�oZş8��ry��F�U<�Odb�O-�X��枱	�f��t�u�ḻTa!�ľ<��-����)�C��UжO�Tu ZSaí�?1,O
�g��Ŧ��O���O-*��R�E�Øh�����Dp��njyRʕ�O�>A� �H�oo�T:FCJ ��q�	s�B	�٦�����\�I�?A)K<��jDl�CW�b!Zu��$W�����iO�i[����!́nGn�c���!�t��!̓�M����?)������E�xr�'Zr�O�U�1f��-/�� �옹6H����'<�ÌyB�'\��'<Ƥp����"�lXR��_N�a{�z���{E�t&���I۟�%��؇$��@���w�ڹ���T<��7��On�r��d�O8���Ovʓ1r����[��58V��$�\d�ѮJ� �'K��'�'J��'W�A�1J� ڒ`u�øu�n�R�$��]�����x��wy�-�*)]��S"��a f��)~i،8u��@����?A�����?I��o���C���"��=�ve1�+̅B��V���	��l�I\yr/�+.x����b[8>0�iw.�.C�� ��W֦���D�������`��W�Ā�C�H%��+��F���s�!�fS���'~�X�Rٛ�ħ�?Y��K��\����M2�z�j�9>�K��x��'��U.Y�O��e"`с��6Al|j6U"|7m�<Yv��0e���~Z������H���W�*X"���낇��	�Ӏh���$�O̍K%��O�O��x��!�V�4� �d��$%�̉!�i�&y`jzӪ�d�O��$ꟼ@'��	A�~=P����[e��4L	�QbE�4m|j�#����S�O2C	�D7T�)Ef��G|��hM�!ז7��O�iR	ŀ&/�O����O~�	�M�QЂɉM�(�Y�H+ö6�)��Bm�m%>��	П�	z�l�"�폨�x�x���5G�`m�ٴ�?����,m��'�r�'�ɧ5Ve/b�Zi�rչB�&��4%�����+���d�<���?�����!/Jf����i8��ytF �;�AEd��I�����v�	�����m��V��B�r�9�
L3,H����yb[���I՟P��my�'�J���S�b�]���U�h�06eֻO�O��d�O���?���(��	�O�Dh�0nQ:r�_�I�F�Ov��O����<a�V�6D�O2Ђ5�H<g0�aA5ŧ?gи�7Ls�d��O���?���c�������c�-�Cg�/J��H���[g����'[RY�d����ħ�?i��k�I��U
$�B�[&i�SH�\�U�i����I�(�g~��MSE�T\\�2B+,GV���EaȦ��'�����+e�f��O*"�ODT�K%8���/�ҴJI*�\�oZǟ����i�V-�?�g�I3)u>9��k��S=���� ̵+b7�ŗp:, m�ş,�Iʟ`������?��V�P��p�qn�?s���A e8�&l×�O>E�I8C��� �rό	R-1s�Z�4�?a��?�DE� ��?���~�A�G���4k��R�X�"u��"e1O��R`T]��͟��Ix?���z](�`�@%+�8XR���c\���'F���dV�0㪟���?�	56���)Q�͍/����8��(ӪO�� �8���̟$�	qy��'�.A8�U�R"�_�d�2��� �ҥ�*Oh�$�O@��?�	Pyb�W�j#�=�B(B�'�Y1󉑚bj�)�� ���ĝ���4a �T������� J��|ʴ�	%1gL����~�R*���B�<!�R�F�z<1���l�D��a�g�~����JӠ ��#H�U�\)ktK�/�}���J?<�����@P"�a��[�-#PEcS�L�a��D��p!f�zq�[)�6�����|(�]�W�T�K��"�쁋+�ވ��Oǚ)��#ʇ���!���5/��EӾ}��'� !��Ĺ��A�l�Ʊ��*�;S|過ߟX��N�uw�(bV�У�Jt`Q��Ɵ����O����%UB����E��%ܟ8�'Xj���PlX!)��L��j+}��%w܀PE#�bs���c�@����F��X3���'(��h��bJ�#�q�#X�4�Tx�O�Z�M�&�i�T#}2�'y�0�0��Ƹ'E<%a
оUOBi��'8 �z��	�1�3�"��s>���	Ó2����c��X�!IV��C�#5�
����@��M���?i��01��2�?���?Q�qC�.�9�xwk7&��l�f瀬|E��@�BG��6؄���v�Ņ%��v^��q�R`�<��IS�Ck����I+)�up�4ux�����~|XJ?=���\�N�8U�Y!���4{~��j�"Sm��D9?��Iß��'@d��)/=�,Y�3e
�EΨ���'��0h���s�a�/9���r�O �Ez�O�X� ԍכ,����k	�4Ƃa`�
:r�âK�����	ϟ����u��'��5�N��F��/��*�!�S��Ӂ3XF ���W�"K��V�'pV�� \�����?�ny�뛣&Bb� WN�8Zb�h�N��8�|�C�B�D��(�6 ğ	�qOMoڮa}�,R׃U�h*F��aɕe�����A	O<���?a�r-V�s�t��4F�8���9P�X4�yb��|T�c/-��y� �Ƴ��'$���R�54JLl�؟���Z�S��va��3�4g9&��I��P��AI��|��ß��`$�^; ����WP�<�S'�4J.�`�}8>�X&I��pb���7�ɸ;��Q��ɨ{"`�%��8�cI��"��XY3eEN�� /��r�i1H�2��$��a1�O��������;ovfMk�*Z�? |��&�2q��'����OV���O���w��A��d�>v�Zč�>_�!�DʦM�2�_�Y����AċOSh�y�%��M#+O\<�'H��m��ӟĕO������'��rg&[�P�����*Yj4Ei �'2��Eǂ�D�_�"�v�;���O��Z��όI�.�3p��qG�u��
���Ƀ	�\@�W͘R�0��\�O����ɬPp�yEAX �>��S�\9����XF�t�'�4\����.|�u���Ts���y�'D�t��o؎p�TMcQnʾ ���
Ó <��8�(Ƥ*;΅肊�6]�A���M����?A��DFpx�6�?����?��Ӽ���"�fY
�% =д4j�a��8���s�^�H��/S�<��b>�O�����&�^}1A@��V���
GK�'���'�y�tl^E�g�@&�p���O�a��`n��:4(h�4Z��v�'�(�[w�����$�O�Lbť�2O ���a�3vq1��-4�)ѧ�4�����E���u�"?yb�`��W���F/ -N͢�aڭ-�)�"!�:>-&p�bG�p�	����	��uG�'��9�Z`�3���]蘱�쓦
nX	���!(Or������<�����[�x��,��#����Ę����Z��3� �lt Ӌ�W�'����B��rU��D�W8^ �r1D���?i�����?)����'l�4 T�"{e��@Ѧ�:#���!	㓵�(ܔL������@�ىR�<�<��i:�V��K�"�?�M����?�B
܋F���Tb¤y�`7*B%�?���Q�x���?a�O�"�h� �lWR�i�\�x�S�Qn��"be��Ъ3O�0�J�rp2YZ�A�>�c�64b�*�cۚ4�\<�Q�]8�̨�*�O�'����C5)D�S l�B�,�b�,D�H�U RV��H_3�6l`bK*�hO�Ӧ�{�%�!u/��IC)�e�.|zǄ~�I*q��r�4�?�����i��+����I5JX��+��\��%�"@*!r���O0��)Q�>Ut��3��e}�Y>m�OY�����;*�ƽJmI"g�O���)�;d.L�	�?!w�<�d� c�p��K?����;'���qEc\��1( ,>}ª�8�?��i�J7M�O��?�(!��5 �%��$V���S�<�Iٟp��I���$̪	��|`�	�4w�i�Aܷ�0<!�i۬6.��4
Ht�G��&��(���L|ܤD��$�O��OP1��J]-En���O"��O�@��N>�d�Z�>�Bt���
� ]�d��׎v����CH�YC�$�!���O-p�'ajl��遀�����ƴ=��JP�>}����)Q�8H� �ݭA���掯|�ûi����;J���A�L��@��Gpb�`V�ig,7��O.X��`�Oq����(�����x���jL1D'�E[q��Yh<)S-�| 0T�p搯!/F�Qh]�<��p���8�ʗП�'���*͙%���& T�(�p"�D3B�t0B�'?�']�$mݡ��̟��'5��ɇϙ�6��e���:#�=�&G�N���j�k�[�P�w�Ü3��f͍�2S&X��C���X���D�J�2���e��m�a�E�^���k�	߱�a$�'�\6֦q�I@yR�'��O,4� �u$4�g�N�'j��t"OY R#��6����s��#	�b`� ����~RP� pa�α�u��'��	ćH���Ҥ T#ľ�P�G�d�B�'��Y��'�R:�\�'���5�Nh��	�S¨܉���W0R�iCQ�	R�@��,-��qF��(O�yѾn�@i��Ƥg`=pV'	�������%D:T�D,�S)��W�mT] 1��W�mr�#�DP4R�h�T�ɚ;tN���� �!����l�ۇ�ƒ il�X!���~!��ۦ!j�h��Qgp��h�/��� �Ab�I:ՠ�ش�?I����]���
X�h-h���7DB��2BK�����O�`:7����q�E�WD�������i�|*���z����U�ϦH\"��F)�y�D\�{���q�K^ Ud*�ⵉ;�',S�	h��y�(�V�ԴL"ɧO�A0s�'O��O��8VG�\��i�B�&��8؁"O����@/Gl�6�t��Mz��'��"=q��$]�e�4- ��4���'	����'���'%�m��/�O��'JR�yg(�*���1"گoN�4Í�d|��ۇ!hy�u�Dq] �t�I�D�$��IJ�!���0uv�Q)u�	x�T[����u"ң���*�D�=i��$�|ʠ�iN<��{�? �Z�h
:	�b�)mI;c���(���I�4�?	����?�}�'�RE�xݐpzG&ѧu�2���B&�����?���sR�
�"8�aԥNb���O��Gz"�OrR��R���O��
�`�J�T�5@˻[��9��������ɟ���<�u��'fr4��k�kPH.���N�55o~l��LE��ԝ��&ޒ{�ԍz��ʫ�p<y�$[N��'�d���P �_^f��c��s_�T�%���>q2��DN�C?>��0j΂�Gg�/~^!R��'�6M�T�'F�Oz0�6$}&�
#��OL��s"OT� '��l�"1"e@���`P(b�\Ŧ���_y�N�(6��O���^N�z�س��?r��[�"\���O��(���O���y>�q ��0o(��ׁ�k}bh\�<������R���2�ǉ�p<�uhYς��$���dɸG<��a֩R�u�4W�S��x�����?	������;|���́��J�'IR�'Q�O>9[�.P�J��(��J\���+�Ġ۴Q>�"�һ j�͒��	9��̓���c��UlZğ��I^���J!�OՉZC�`8��$W����&���2�',6�o*}L��i�nM"`����~)�f�R엜N��ay�)ڐQ��%�p�>ɀ�(ΰ�Sd�4o�RE�ЩZ)��O(` ǧ��&�T1�FG,]�*�O��"b��O���G�[�S���0�?<1�K�d����?I���䓡�'?��ǥ�%H���I�y�P#�-:�6�z�&�O��#�@E�*����
���vj���5�	ٟt�����@�����џ(�i��2D`0B>(�R�[?8���rN��whF2SB��fQ�)�Ǟ��|�a�>���Ȧq-�`[�7;��q��<;�Vl*���*/b�� �[�
7�h��m��H^�S;�M��w��I��ݵ49޼���7Wa�d�h ��M��V��C��Oq�b�'j��K'��eÓ�@�a: �A��#���d%P�&|����6��b\+�d�O��Fz2�O�]�
�H�T����@eV�Vw��uɓes)ʰ._�\������i�_w���'b�)чx�p���g��9��`k��)�`��O�q��I�/r��`DD�/R��T��(�=<�!��	�/N�|���xx�:U	6|������'���'tX�\�Ϙ'��m� *6V�@uh���v���	�'�<@@S�U�#A�(�Z	n�y�Ǯ>I+O`�;�c�ݦ=�I���,�3H�]	3��;=���ڶ��۟x��(萈���<̧`jL=�҈Ű�,1K�O����Ţ�Z��DA<vPv�sE�'���
2)�<��FX�T�EJv�a(Gj_�=ڜ��'& OV�i��'��V������;T�Q�D_�vb��a*j������,�?E�TNƣb��ّM�
E�5(���?�x��y���K�#YD�\-*�.�}�H)�2O����2�ix�'���97�J��	�A6>�0Po�)A��qz��_�\��I՟�r֎�>�~�s�a���T>1�O�r�2�l�(p�,�V`�9@OL�iL��PgJ�-c�n��\U�O��4P �72�8�r�ɈC"H��L��yV%�O��n��M#���O�:��B'�3}�b{��)Yt�j�y��'q�y"�S�V�l�jR�ڻ`$8�Gl��iў���HO 4�EY.�]	��������Læ��������Hޔ��5���X����l�������=u�x	�M��dt�:cM�'�< ��֗����q��I��'�&�������e�pM2�E+r렔���L>T,D��X�)��ƹ@��:m��mǛ��z�@��A�h����Y���I��ֵ��ŕo@�m!d��	���)��O�6�Jv���u��F
b~b#ғ��<yX-�`�$Z�
,� Hť-��c��D%�?A���?	��SٟL�'?�:)� ��:H��H���&l��n5*��Ҡ���2f�M�u���&�����@��x��'d�-_��)��[�c}�%�%^�}UV5�6�R�Y���� +
�Hd�d���BAQ�Y�d0��R�k��2c�'hr�'+�]����_�=���j%���P'rXa���8͘H�ȓA�VR����U3O5���ėP̓9ʛ�'���,�8�Y�������C0"�8�:��T*�oK����OJL�׊�O���a>�"����F��a���U.�l�s�(k�:�;�AG,_�L4y2�M1*]`4�����::B�1Ӕdś	z��!�T1@�`�3b�54<�4;��J�d����Q0Xۀ��/ڸ'�m`��iE���>�R,\�xU�ɚ����iv �A�[̓��=���F�Bd�bN��hH��E�Z<0�iHB���#?���O�U6x���'�O?�I;*�\�!7
\����)��2k��B�I��X��ç�M���p%��1��B䉪`2
H;��ݥ9d�p����3x~B�)� ��`��%z7��ֈ_� �b��"O���G	](I���� ��p�v"O>�"�Eyr��c�مq��0�"OȤ�E�(���F�^@�a��"O�����:|s�Ͱ&�\�L6��4"O��R�a�:i�d��DU�
c3"Oh����H�9�Ai'Ú7M�ƠYr"O�{PԜG�&���"1E�ɠ"OZ��ٰTZN�k�A��""OD1�����B#T�k�A� øe�$"OH��/�H0r� @B"U0�Y@�<�5IN�cZE�w�W>6�z�Bq�f�<��F�p) s�%����B�b�<�1�ˮ,����G��~�j@��d�a�<�X��e��� :\������I�<J&q6��&�FƁ ��C�<��b�:ZB��vLY9[�����g�<�an׮}�p�*�gԶ-��ɚ�jPZ�<����!(��STN�8�^e�_�<I�	��C����K�C���IA�W�<�� A�E���g(�(Z�UqGPk�<)�gM�=�lAF��'?s6Q���d�<��$�u����C�0��xMB]�<��֥���;w@��h�ش�cd�Z�<qg#O��^�2�XGwX����Y�<a��G1v���5&A.:�[&i]W�<a�N�+_��	MW�Y���C+�j�<��艎:�He�""�#i,��Q�g@}�<�R��dH� Z"@��Q�GB>�,H"Q[�$��D#�9%�$�O�h��Y����9������	Z�J	����$�34ޔ�gU�[� ��1��31V��c��&yj@�$g��I����ָ'm�rB�����$Kx�O�����"�=
�qB�=,�>�$.���TxQ��	ld>�w1&	�%��*}�.��!�e<��|�x����
+ [ӧH�&±��	��dx0B�Yk��q� ���'-n]:�f��`����H)f�#L<Y6��3��!B�t�nEAI}�$)P��Jw/��(��I�gy�I�-E�;QDESAjɈ^�6����0 ��q�W%��;\ŃhC��	F=���(��E\�'����/ؖ0r��T	ω5�,pI�A�PD���.m��I�O:��&b�'U�vh����:
���
�*O��4�cA�+"�!  ����'D��.]�
`֍h�Ê@�'v�dJ�Ӻ�X� �']��`3�Y�t�0�)ă+�HO�_�B�pp+�wg<��q�,Br�M��,���й�s�:GH�c�Ѧ]�2��������yPS+��J�\m!��Qil����ұO�`C�#��T�*�p�m��^�D����x�F��S<m���P����"��J,2��-���J�,��H0�O�l� ��4O"�����.�YIU��gn�8��� ��d3D�Oj���xr��c�؉�@_���=�ՇS;Tj��F.?!��en��i%�r� (K����f�9�RJ	'�����"]���?Q�\x�)�,� ��D*��nQ�xR�U\�(hB(������u��W��AQ7�=t�h�ԇ���Mr�$4�(O�4�4��i�;>Y0|]���0UH��s����1 @�h�w��8�O�>e��!FR��]����0��� �-�8ޱO�aI-��X�H4PriʚV����x⮃�`a���#-W��}��O��$�D�̹zuMG-)L���?>��%�c�ŋ+�jHc�M'!A�5?FeR�pp���	�PM���0�aP.�+G��Q�E!�@�'�2��I��<�|q��.OxaL��eCT�(��q��^���W["�q�C��#v��8�/�p��O�eA�%_!_yza:�B5M��L�'H6�O� ��B�f�bԃ�*1��4���D�;k@��b�y�``I� �?�0��D~����j�9`���ƴ����0>�����Z�`Px�d\+^�.-�n�/+��S�O��D��N����g�<SJ�y��p�2������G9c���OL('��A7KēWބ���CD�2���g$?Q�펚�Usk/<+��ן�S׽jn���o�=43D� kO"q)Z�,]�T.tP��D�I0��#���eL��I'e*H4ڄc^:f��I�W���L�ip��1b�ՙM�",�����S>$�B-.?Y�a�H؁J<~ƌ�8�!Ld�'���ba��F�D�R#�^�py�}����
a��H($HU,12���g?��T>�Ӽk`�+^���:��*?�d�Ѧ�`�cN�x-���5�ɻZ!j0�tl���(d�ʡ=�����O4���!�\X�	�G�iZ-O�1��w~��梆�PĜٗ�W�zxh�A��$:P`q-O��Q�x�� �>:�37��/v2̑Ʀ��v��I���e�/O����ǈYy"�]m�p��x&�ԫ@�j��1:��^3{S�7͔�:�)�,O�ؙF�W���J$��^���'���=� ���ԩ�D�
��w�֪� ��OX%S�_yN[�_:�D{B�ԒlAr�J3��"��`�f��z�L,˒,֫0�΁jR��,v�p��`��<�;O�+��=�p�@9z���~��V�k"�<�㉡������'�T���D{����>��fZu?��]�؈�O���`�َ!!��G<��.��>LFD	K�>廠�E�F푞4h��H�A&�ɇ<�4�jW�L'��C*�#d���]�H`��S���'�h)R�h�r��`�H�{��<���)Rۀ�Ă�JY^,J�"_u��Cb�O�B���Ղd��ɿ`�XrP�O��R���C4�`��hU�T4i�!V�(�j]��N
YVd�DM#?��K�4�O���P�?���@, �]�3�:Lu�p�w�+$@�������ޛ{�� 	�P��G�	 �&dwN!���"8����Ć''����At}���f���j�aYe(\����dV	��h��O�y�������a�RL=\	7NL?(�pEx�	.a�����ȅvz)�f����$K7{�����c�P�׉�Ȣ����$_%V� �ӾA�(�x�H�8m��T`A��l���1��7'̙���H�`��s���Y���{wʌ9,���n�W��l�?��O���$�F�+��=2��ZB
e��
�Kx$���C<\�!�@j/���W�o<��<фKV�\X�k�LN#�F�IdV?8dT�?�O�+dLO!��O�:Ї+ ���5ʃ�q�����C!=8a�ԡ�z�'#<����?�yL�>ChzՋ¬��OE��ǌ8�?1��ᓢ J�X'B�8��cL4���@'�^�'hD���F�v��pxgָN��e~2��-&h�����iW���!�	�V�5҆ƛ��L���M�y��A�s��*�r�Ul&h\:6J�3s�1AW�@�!9�L� �[����,�ID~�̓�!�,����<}�N�F�����d &{s�`9%�1.��-� iX�Q���F(V����i0N �{P��;F�	)b�O��9B�i��i��[�f�11'�!����:�H��a=S�Q�|C*�o@���U�uq�f���Ir�a�_�p�R��I7��Op睴1b"p���.��P���@�"<�
X0)��E8�j��P��%?�UϚ_�Y��k��y��x��,�Q~��<��>���9:�y��$��u���oE,q6Q��*Q�,���6��@~V�cK �K,��0n@�'	�e;�/�Uy��4��(���Ȥ!��<�2��;��D�4W��I�7Xz|b���s�'_�C�>'\�h!Iٗ+�:e��y"AɷkB:d����qT��E��^}-^����!y�4�Rn�5�p>���Z�V$D��4�8X3�_���Er3�5G�� Յ���(O�4�O���I=�yw��:L爕���$z2 ��J�O@\�e�ƃ5�)�'� ��OV=Z����i�l��%!P�	ی@Y�>��C2���S�$@�I[�A[dŃU�����!,��,2�X!pN�!�C���j��F���~RI<��l@
��O�
V�ڄF�"|�g�'J`�k�[� ��E���(� �A�]���I?t.b��Y2$��ʝ�}���Zc�W��'Y��X��4�|�ir� ALUA�]� 0{��W�fqP�D5��O���1�G�.�#D)��^Hz�I�%�Y�Z�`��N[.}dH�)§l� H�mK�/�,(Λ�"_�MT�ӆ�O�|�4�˶`�(X0T�}ž����D�1.Y�eK����EӍi��B&�~Rf���!pJ�J�d����MíF��Ђ	SXc��'�Uz�z�� <o�0��O�;�B�Y!�W�w������!c�����'�R�r��߮"	L���Ѷ!����Y/��j���� l�CX?��05�Όf�Q�
�T�nO�;�K)hN�A�ƀ@L⟠�'G�8{UK+�ħJ�ꍂ �[ q��E��/@+JG�H���H��C�,�:x��p�Լ۵���*�D(ީW�x`0���'�^�
E��~��	Ǝ%0l�Z1*K�pY�̏�]�U�D#j}�i��jD�n�����?k; �'yhEO 2�D��'N8>�	�����'�H�P��@@���h������-%J�eDg��T���!~�yr!��Uq�#]���P�/�'0p�v!Ou����F8k��Q�ͩ a^�;�A)#Z��&��axޝ�E�P�0��1/�����Hݚ�j�"�� uH�&>l��ХI� -�(�4�[*�lc�[��X#@Ҧk�P�Ӽ�OW�#��pa���6"t���Rx������<��&��X3p+�gFL�"� ^,8�B˓pЎ9qq��A}j� �n��'b����;(�e�s)�ED��b`^fd��Dz��(TQ2�'��)Ą�>��fތBv��u�K�	7�iD�&[d�I���M�5�N!t �b7gV{��ɀzу��'�D�Aɫ#w����;o��
ش�h {q�<y�nF��剒2�~�bK���"f�6�X��D!��G���`�e��������ۆw���"��d��YzY�6ʖ��	a��N5`m�����Ey"�I{U��>ͻ=�4r�.l:�!��Z7R� umZ�Nޤc��'U������$���(~�z�C�mY~���C�"X"L��	�i�R�'��������y'a��}E�<�(��0�&T��EΝ�HO�E؞���Τ
y����J�Ԧ}3�͵A5d�xg%X�jC�4Ѐf??Y��Z�U剁]��-O�ik�	ݞ�?�`H̀#��a���N2Tr��g�����t���;�Tr�n�3�?QA/	�L9����Ã��)�$y ��3<0���ǫ�Q?� ��  ��Ic�p��5�)� �� CEJ�|����ϴ%����
/rԤe�@��L�U��)��$�|��y-S����:��GX���a��M�4H���#?�u�E;~�I�%c�� ��[7�r�)Qg�6���k��](B/�I�>æY$��s��4��4���Z�+��5QČ8 ����R��&�����D��*����sb�'.���⣜:_��I�@Ş d����O4��?)��'�$Q�#9����ƛb��@�d�� �P���H�"2A��ɔ	@(��Ọ�.?A��
��-8��Z ��Y��@Y�D��@��ӷN�rh��F�I�E�O4 ��g��O�ڴ8�o�) >B�'FB�'�ў�[M8��J�~�
�/سr�ꀲ�L��a��고Pq���'ȓ2t���,Vx����N��93��9W��D1�S�O٬)ġ@8+L ��@~�E �ƎL����' �Ba�U2LV�C���%���#� 9��p�Sڢe�JUD`�<���D�;\�U��`ɌU&g\�`�x�Bu� �O��\��Sƞ�p$�	'Q��c�5P@!9a�)ʓ������C��	"*djV�ժ\s�z��U�Ф^�9�A���:��=�?q�f��I��ԡ�&I�t��8`�I>w�Q��E{�O�������:cAԜV:$����:�.�2��P�s�Q��Iļ�$��w*�C̈0�����O��N���'Q���B/��K}�����3\�tg�	S�kĘbƌ�LZ.�+&S/GLp�%��r��[�qM^�+ �ƪl�v=���6O�4{����Z+�����"*�%��"N�L�K,��Vz��.��#�����ΛTA"Hha��:*a⨅�NT,��U+	������i�i���(�8����0tS0�Ł�%>?j$Gx2E�F�� �"C?r6�4*Q�X��B�	.l��}Z��y44A�/*����2ėeh�O3��?5C�'
S�ݚ2"(K�/E�U�Rt�eB N١�d]9QO�["��&/����O�U�di0�}rO��=�f��Ԛ�"���ēR)l݈��Z���sfل]q����:+�b`gĉ9$�v��D*��e�O�?G��(���	|�@�9�CL�p�qPB��L���~X����N����ʠɞ�V%�@+� $}�I�-J��R����k�J����'�5���� <@�4�Z0���Xǆ(�	��R���&P?�aG5E�U� ʚ(S.�Lc��=6�<YQ�FKN"��DzZw&\ٛ�������ԀV��]�uɟ2<Б;&�*Lj�Bͥ��I��ugb@K���䲩�S�V�@P���ɩZ��C�	7s�&�0��N
q��r�Ȫ?P��D._��k&NN3��(G���!�D]�@f���6j�.K� `f���!��:/�
��U���2��*e�!�C�'��P�7g��e��FU�!��"�2$�0�L,����Q��K!�$�2&�F�`/��fF@��Y!�d	2�	�ê�);1:aA�TW!�E"@*
� �c�7W%�1�@�!�!��--Hޝu�U0xl@�D�s�!�$M�A8N �bƝ	\�>as#���!��i32�����:E,@�E@ �!�D�/nX��C���>�����R�K�!���%L���p���O�����c�4)�!��6W^��#�L@e��CF%�!���g�Y��We�H�!\=1�!��� ��aP�m՜cM�1�ď�!����$��E(d�O�l1:��1��q|!�$KnK| �gO�/��у�>l!�$�*1�a�&��3,�٪4�>�!�䏠f�F]�FC��C4M�;;�!�ē� ��焜�L�$=�v�q�!��,d����� 0ЈB�)U;P/!�$��Z��1�F�ޝ�h�جg!�$��l���F
  ���Nߛ�!��ߺf7��2!I����I�rK�3h�!�ėah�iQb�
o�ZEii�>�!�H�"V 	��["�t���G\)n�!򤔶O�P�H�;,�fef��<�!�D@�iߔqؒ��/�V��SFe�!�d�X�51�2t���J�䔼q�!�$��D�n-���P�&�YOŢ9(�B�)� �Q��P�.P��ܸ}n�k�"O �Q�a�3ll�M0T�\�F�h"Oz�J��i�j(sp	K�z�UA�"O�x���6l��!'7p�|�3"O�a�0a��Ls�B�GU�eQ���"O����AE�Qq4�!��@8 �1"O��;�K\?�yaw�
;#����6"OsӥU�u4�= cNG�J���u"O(�J����ۆN��H���"O�����$�c(ۍy�P�!p"Ol"��%cxi�@��[�]�"OD��ǪH"���ˇ)Ƽ�jt"O�̈���0W�¹
Rk��Z
j0+�"O���3��6��a3D��l��,{5"O^���
UYtF<O��s"O�<��#�(P��ṡ�B3���9#"O@��f �'mr�ڵ�R8l��e�d"O6������7X }�%�՘wϮ��"O�m��k�\`�!0�U:#��2�*O�Y�a������gC�
 ���'mN�ʐh+'��$0�����
� �'L�pYh�;Ѐ�s��K��3�y"Ǒ�l���Bd\�q���/F��yr)U()�<1�bnP	X� 1�L��yB�I�F����'NV�HP�4�a�ց�y2#��^�"u�X�=L�Z����y"��Ql�E��@��J`b`�F7�y�n�px���O�z4�h²�N�y��Z������C9k���p��T��y��R�]�l�҃�V�ZEh�Jr����yn �fΠk ��K���d����yR@�? ,1K�@��&��yRĂ-L}d��A蕋��1s�M��y+����u��-y��[%k��yLݥ&3z���O'A�4A�T���y�I�	�,�	j��8��\u���yb��J�4)��e];nQ�S(�;�yL.+�Pl`��ޓ,a�X#�ğ��y��E=M����dbC>+����a���?9�i6�S�OԱQ�"����`�]�2���'�rp�cL���/1�Ke Qd�<i�Ŝ�Z�0�١4j�0I��a�<IF�ϐS`FAu�]Rq���b�<ٕ'S���pE�b,	��n�^�<a@�ƾG\�� g���?ar0�R]�<���$7L�P�-?7�\bddDS�<I�D%L�"��w�|���T�<�Cm�=7Pj�Ȅoυ��I+�WY�<9��X�U���8���n&~5c��W�<�CP��h�)W@� �i���EM�<�t�V�����@��\qgMPb�<a`f�5*��q���d�}!�]�<@&�qXN�qxs��5O�O���dM�(���� aZa8��IA"'%M!�$ү
�p�:3L�@,�]��A��>l!�Ť�r�0,~8\��bO)0h!�]�`�� ��ۚ4si���U	,!��%P�I��@]�q��	�:<!�[�ge��RP�Z�/J�����,-!�$S	-��v�N<��ۆ�$)!�$�����ǈӜ���Q�Á�D!��K@�2�82�D��Zr��H�!���/?���1@ d�Lݳ��[�z�!�ć&�tU*���'c�\��$�ݺIe!�� V#�I<@eP���P3D�D�ۅ"O�I;�&�z�Rx�����j^�py�"O�9#�BѤ
s��IG�Ğ|_Vds�"O��� '�=��( %+�-OB��2"O�<����85�܅Ћߎ'K���"O����-p�5�3�� �&��V"O�U�
�E-`� �OTM/P��"O�M� ���l��h�U�I>\*���0"O�%ɗAH�&)B	�L�u7��ː"O��$��:q�:I�1F�G'IrU"O�-��R�3�ʜz�U~8���"Oh4`҄�Bp��{u&�N�`Pt"O��ȖO�^�\%���a.P�"O&a���ӁMd@tR�iD{&H�p�"O��Q3�C�W8LHCҨ��'Y�7"Op����0f�xH��̨QrJ�:�"O��V��t:(��Tf��
ml��"O,�A�,N�R���ʔeǀ|�m�p"O ����3)�X�ّd�dH�k�"Op�jU��U:*ݰңG3F@i+e"O<���Y(eC�l�ҡ�"O�}C�B[3@�ƕ��'D�"���"O���Qmײn���a�K�ڡx��'��D#�dő$��b���/@-�YSC�J2^,!�D[,q�,8vf��H�a(�"m-!� "V�]�K�6�l�񂧓�3$!򤈧jh�(�ޞl(�(�ƼX!�d��\hpa�c圜r�`�3�\=@�!�� 
m�0k���,�A&&_&P!����&XE�;�Г(��!�dF-_��"�'�t�6�J�G	�N�!��T)�x��$�øz݀��e��$V�!�$M�?�f�	�#%y�|(�L��]�!���:�$(��S�ch�%��b�!�ܙ;�� �sÃ?5O^����"�!�Q,_�z�u��0;����LW"F��IW�����Ձ�6]=xY��HT׸���"O4@���עڔ�3�E���50�K�HH<YEeV��Щկ��=��_j��XC�}�C3Q eЂO(��pٕ��M;�O,b��E}��E���ƧϚ#.���ǅ�y� �Kи���+�@�)�.ñ�y��*^���3fS�[ � ߯�yb�����4�JG@`Yّ/!�yR9��/�/|���1$�y2+�9���D�(HD�P��N	�ybfK�66���V&�t����Q3�y��Q8H�h�p ZT��������yB�?��c3&�AX�Pd��y���<z�2�I��j&Ba:���p=��}r$^�h $�Ed#g5�t��'���O#���9�X�lR�0ltXw�TL�<1P�V ����Ub�:)�愂nUJ�<i o��p�p��ȹkq��cd�G�<!5��W���D9Z���3f��O�<qE�9'Lc�jX�z�|uۃ�I�<���(�\DI�eKGf�L��#@�<��S�eF�dɕ	L�p̀Yp"��}�<�W��u$��*���!~�p�_�< ��  `���g�-c�K��T[�<I���|�UطkԚ8��b�Ҧ�G{���i�x�b��sZYS��?*�
�'[�%�vŇ�=�Z4�SaD<8�p�'� 5���F��������>.j�!���� L= f�A��9�sGH�-f
xѷ"OXX���! �ٚ��̡wj� �"O^�(&ˈ�;�+�Oz�8W�K�<I�lE�=�θ���Ñ�e��"Z�<��Dq���Nb�H��΁<�L���e}��Д|��D���K�Db\����y��]���J��)2R�j�F���y��W	id�h�,���F���y2L�76XM�%��v!�o�hO���$��8@�}K��T0P��M9�ɇ(r�!���Z�̓��>��u���8I�!�\0j����ME4U���B��-�!���)���xW�+2h� ��(b�!��i�ȑ��E���D�u艗!u�|��x��֏=&��i�E�]EF���6�y�� ��a�gV�\^��avHݧ�HO�=�O��J��hy����B�4#6���'��@0&BB�LZ�t	.�����'l�(�t+Ds�>q
����+Y�AAV�)��<y�	��aP -¶Y�"���s�<�T/�<q�u��ˮ.�J���!h�<�`���~��H��(F���f�`�<Y lC^�f��E��-��|8��_�<�T�� �����.<�XlPQ��U�'�ў�',&�	T��B���gH� ����=�Q">8(�j&&�Ħ�p	�'_�{�	�_������>�8���'���rĕ-J.vYY �Ff� �-Oȣ=E��V��,��#�w���$�O��Od"R�K�$=#���4�F8[ ��W�X�<�%�ܠ\=�1�Z3?^���#�V����>b��!�:�!s��.E`��H�I^{�<�!B\3���"J̏Sb�A�}�<�V�R�U�$A�%�ē�I2���d�<��F70Ĩaq��З"*����5T���F�T��4��b�Ȁ��X��n7D��4
� 0�L���5I�P6D���G:Q�b��G%
�>5P9��4D�TAW(��� ;/�J��1D�H���ߗ`�,�"v��;] �ത/D��Sa`Ș�t�!Ы�0C���i¦'D��z���<����$�n}H�&D��R�;/VA��9m�4�A�'D�i mU�u�L���L�6س�*D���K�	��0�ɢ}E�BG�3D��`��ϙ����F�_���?D�,""�=L�:5�Ă�A00�a�)D�tJڤ&�ț�lB>�����R�<�1B
� �C�,>�^����Kx�<�(�W�P��K�}�x�f�H�<�r��f�~���Ѧ3�v��f�A�<��o��7��՛5��d����C��}�<a-�7#�*��2DQ�5
�Dr֪^{�<I ��4y���A*E:.<�tE@�<�`��	L�5 E�I!4��%;a}�<QpM�;(T���T6z�wE�M�<���3Z��uω v"�d �F�<&��(�x��%C�Db�B�<Q��*�:m�7Š'*��w�FU�<���48$�I�/��]#�5�P�<��� `���%�́'�,ǢUd�<�g�Ȳ@���&�U��`�
���g�<�Q	�H����	-`H���n�<i�!�%f��P��\.�e��d�m�<�  � �E��"�ٺ�OGC�t�"O� ˄�ó@�Xk�/F�K�6h� "OP� ��ci��8���|e��J�"O %�Ta�P����7�ӯ^؄i "Oh�*$�BCF����D����pu"O"����2owX�їH��N؎!2"O�(�;p8`�&�Ќ�$��%"Oȱ��*�j��Y!��N��8I@"O��j!l�
d��	D���W�	�
!�Tq1Nh��
y���Qv��!���H#� ���U+^�Ơ�6j��"I!��W'}*��0�����`L�,�!���1j�a���>~R��Ԭ��E�!���4I���)t-]-s���(����}t!��٥r���g�˨C��̐���*q\!��Ŭt'�� T�zou��՗kY!�dN�{���	탚i��z���_�!�	0� ���4q뺠��"��L�!�$�;0�R�0F'�+Q��e��"gx!�D�?���а/��'���v�ըA�!�ď�6! |	�*[�� �zrnL)@\!�$H(L��ԡ�|�nx�E�W!�ޟ�<�7��_��i�K��(�!��:|��H��@�K� �@U
Z��!���4������ k�a�b�Ǽ�!�B�����Ĕ�@�ԫק�+Q*!�d��{����"\�~/`؂'��;!��;�,x �%k)>���JF.�!�]�E6ZU��,��@P�
j�3l!��~�8Q4���O��!RB�_!�d�,^k8H��ͣj������٦oM!�D�1�*щ\3B� ����#J!���2�(��&^�Le���)t*!��%C���Gd=
������7e#!��ٲbv�Cdd��v��#�A�7"!�d��Ґ��a��<!�m�W��=?!��dQXEi�)�<���ǈZ�V�!���!��\��G�
F4��!JV�v|!�DY�,V2�I1-�� =���,Wf!��]����C��1���h!�Q6x�a�Z8 ��U�0$�5W!򤖨y.E2A�ڕMj���E�H!���P�
�B��߈d�HyA剎F�!���n8�y3Qo��M�Z���Ò�s&!�x��u��Q+4L�(a"O���"jP���������"OЍ��d�i��gJ
g���"O�� V%�+a�!	�6`~��"OT�b 4[R)�&9Z�ԕ��"O���)hD����*Z&f�808�"O ���)����	RJ�]��"O]y�*_r6��VF˄M,|x "O|1�h
 �Mj����A"O �y����r>�$�	�N�A0"Odx��拋	L ���B��bd"O�h0�,q�Nh@w'Tr��i�"O����."�fY��%�p	n�p�"O��+�FW2k�
�B���-��"O����CL�P��u� t0%��"OrtQ�g��!��r!I�lY �!"O4Y�2C�6�����!�<+��3�"Or�zfl ��mh� �5{hl�"Oqh�C����hb��!Q�j=��"O������VY�([):�v�""O� ^r��͈J��(Z��͍��$1�"Or<[��I*m��	E�С�&D��"OD�0��W;]6*��҅20��[�"OQ����l-N���r��8�"OZ݂��]�>�� c�m���J�"OTy�wL�e�vI)�̳*�r!0�"O�YR1��N��� c��URXi�"OE�%U�`W�Y�7n�:C��5C�"O�!����=~��[d�Yfmj�#�"O������pz��T��ne�쉄"O�E+� ���5�
,O&"O�@�����.�T��W��w#�U�r"O�0�5Iײsp� Z%h��o>�q"O6 #�g��L�ڤ`��P9Z�+�"O�m�Df�j,��*.e�\HT"OX�Hc��F�̬Q�1Hd��@"O�%+W��B8�+1EB�P� ��e"O��{Fؔ	�"i㵣"�X�3�"O�!�'&�:堳#��:� p�"O���V�%>j�����.���S�"O�y{sO�.>��jF"��N�"	��"O>�K���8!�l�Q��w�H@`"O��I!���3a��
qD]r�"O�����c*씢��ӭ\���#"O�y��mT>e�P� ċ�X�v�#&"O:�"��I�,�Pc��^C�P�f"OdD	ٸ=�]#B�6)4Ht�C"Odd;�Z /� ��ǆ!�DH"O���@�/� �s@��۾�J�"O��Q#��!oZ<�f��)8�fLx�"O�����2~��h3��7����"Od��A�n�Y�c҂!�z���"O�=��;\���Y!b�� k��S�"OhQ��E <J����4w[�,2u"O���� Q>��ap�ED/�d�<A�H�??��H�ۃr���MT^�<��(
�L;�M@���
� 1�KZ�<ْ&
. �b���	�_���ƆR�<� .�= Tm*���e�!�FQ�<�c�A<iW4s�\XB.x:$Jg�<)��+'���3G���"�t��H�<1ah�}켴�	^�_qb����@�<��jݮ����@P	h� � �@�<����7m�4�P�O�r�� ���}�<��: wfi��.�j��@���v�<ѢIa��a�%��lO.����q�<	����z��mk���f�&P��(�q�<х�L}=�bMM����m�i�<�ƃUjx1���<5Ŋ�86c�M�<�aB�	���K�탶cB&�pF�G�<�D�E��Z=Re�� wHC�<i��&?��d��	S:d��ɀ�Ā{�<�gS2c����kܡ6�60��<D�$`0�Hs~|xsK���p9��>D��Ӷ��2�����	p.@�J<D��z7(�6/�$X�l��(�C�>D�ూN�%������ly��(D�0
"�^z���C��2�:�m;D�d[ 	�#q�5JT��UE@Y��.D��f(r� @xq

�2~l�BC+D�ĩ�/"T/��`��;fvpY�'D�̲5,�a�9�G�Y����$�y�S���w$LdeP��Q�
�y�j�t����%�O�%��- !��y
� �� �M\��,lÐ��g�% �"O����(ڈ,ô���S�T��"O.�6�w��,3a̐�$)�A"O�	�B��k{x�b��.�f�"O~\�5HF; Ef�C�	ێ'�.p��"OA��`ǇPi0��V�,n�L=�"Oh} �ʋ�a���ao�<o�̱sg"O�8�&�N= � nh��T�"O:��G�Ǧp ء3��@8]��"O��C�@�J�LDL�I}��"�"O�a�� ��:Ւ�����%N`TQ*�"OBeAg�W%c�r�[�/H�>�,Є"O��P�ښ �Ft��96��Dh�"Ox��w�A�fv���$�E�!�r"OȽ�gj��c�� 륡�;C0Ĭ{"O�Z�g�~$�(�!�Y	h� 1"OH�P��E�+FY#��A��.�y�A�<p�� GG�!f&�Q����yB�˽r��`r��Ɖ[(�`�E���y� �X.��$�ݶO;⨛��1�yr��!���KK�]��i�SOX+�yr
��-�,MKS��P t)Q�eʗ�y���b]�bV�4\tL[$W�y�eƇZ��a�VI/ ;>�RW�P�yBֽvA�������L�6h��y�!�%;f�Fꔅv� PsE��y�o\26ٜ���B�=ZBǛ��y�i�(ܠ���g	����qj���yⶰg'�ez�uR��X�j���'����+S4q������? �@��'/��xr��h6]JQ���5&,�R�'�V�� �6�t땄�72P\c�'�h���*��B�]�$��U�b�
�'�,w�@6h��D¡iW�Ib��'#�]8vHϕid���eK�:!����'BxQ3�!�>5"!��;'����'VF�b�K�V��(y���)4F�8�'��� 'P~zY���s��\�	�'e�e*�d��w2�M�&�H�4��<x�'"}���M���sc�3}ɚ�c�'}xUH�H�V�x��� HWؐ�'Ī�������)���'�IJw�D-lR����Tф�a�'EN ��a�0u��ѸUI@0v�V���'��PI#兓/����D�ͯ]��8�'j��b� R2fŎ8{��XYݬ��'�Du� 䍠{��r��]�6 3
�'���s�f�
(�B1��"3NA�'Q����� �yh�T�'_�̈́�3�'�T1z����p�4��N��e� @R
�'j�h��!)?Z��A��ƻ]X(�1�'�ȭpi�4J�݉$`V�m̈��'Y8(I��P�y���įM�Ps>��	�'�F��(Ew��pv�>z�@�
	�'���Y�	�y.}�`�w�x*�'m�SFE��ObKo�D\����'�ʝ�# ؂s�ొdi�;f�|�
�'�big-�el����Y�d^�	�'�H�臂;�d�ƋB�T9�tA	�'���a���"��s(LSpU��'j�y�a2�T��C��Q��D��'\�
ϹV?��#ӭ�]�
�'n�ūa�����h�d\�&?�(�	�':����#z@HI �"U%��:��� � NG"w�"���n�%v�h��u"O	06`ͨPe���p�DI���E"O`Y7�I7�Jh���=�>5�"OLR� r���a��Q�wN@�"O�X�%�)"�,QF��Ud�*"O����iI,|#0'��EJPe��"OX��]%zb�p��"k��!X�"O^T���<w����h*~�"O
i8c@T�;�]�Dפ"��t"O�e���#r���ą��)����"O�����ъ���!�d�xq�Ja�<ё�;��p���/|<(*�@
D�<��)U������676b��B�A�<ف��k��q��ͱn^���$D}�<Y@倅7E,�Y�� ��49F�]y�<�C�X�+��!p��Չ^,��8U�Hr�<q%bH�j���
D�j�aq�<��՟L�
� b� q=,�:��n�<!�N�4Μ�0iA4<�2�걋�B�<�c ��N$U{` ��!�-���e�<���\���[��@�y�Nr!˙]�<�v#�0'��a 4dY�Ա�4��Y�<�bDbqPI�fo���l)'��m�<�$d��/��A�W՜�����d�<q��LGvM3#\�x\L�I�b]�<�B�9f�`��@�>��j�r�<I��,M� rJ��X�AoOl�<ه�G�%i Q��͜~<ȸ�m�<�'�Q/9-\Yj��G􄰐/W]�<"�	]��$K���R��EV��W�<� ��3\D1��`��L.�H��^W�<�� Ű*wT�N �gr��T��P�<��Oa����+NmJDq��H�M�<i�dX%5 d!(1vH����a�<�"O L ��� ֘L�9q���\�<�&��9Bm�lh�J��m�#�\�<тi�%h�Z��� �80I��QX�<���T4��SK]�G���Ԋ�o�<�ׄW�HKP9�'!ƻnM�$`�Pg�<�#B�p:�� e�#r�j@3���j�<6�&0W$� �N�;H�p�"�ψg�<q�Bرv�
�:��I�&ihF�TZ�<a&lT�n�0��+Hi!�d����W�<A3��9~`r5'Q�3`� $�K�<���s�t���@���qh�H�<��O�O7��r��~��#��E�<�FϽA�"����<(�M��j�<y���yhBy���X@�#b��]�<�7NýJ48e�Eւl�L!�ĈZR�<aC�,n#�8q� 3Nk�� �P�<R)�<}O�IڤK�2��P��ʚI�<A���Gh�%��)#���R6�C�<�T��Z��$a��M$Ʋ�)�)��<�aY�d�R�IH� |׶Q���<U��̮�#��@�΀��(W�<y'`۲免0dMDl�t�G�S��t�ȓ��Y%��U��p!�F�f�U�ȓ`��L�FX�;��Hc�D|�J�ȓ%������ǀ%�����8?RP�ȓ\S,}*� ��~�޵���6�Ё�ȓ"S��RiP�Ƣ�Y�e�=^�(�ȓ'~�)��@�)	ХA0.��}�؇ȓW=��
�הa���*��gm0u��c5p-�/̕!)�i���Ad��S�? >��Ղ�5	�UR!H1l���[�"O$m#�ޜT���䍘�$[u�0"Or5�6$�l�Q���*5Or̡`"O,���M�V��"�a"E��"O���OZ.���А�<a 8SD"O�p$��B�J\�� ǁ)LH���"O��P�ᄫqJuRV��&:&�x�"O�ţā�#���e��bL��x"O&�p�o�|�~��b�+(CdH�"O �hC-�7t�셻�,֍|> �)�"O8�i���`P���$ePW�`,x�"O�)[`���
�.a���,E�`� "O2��e�M}�����##w�|��"OTUR#l��$��C#E�][�L@�"O�py�����)�b�HM�aa"OV��)�*]���)t�9p2:yʅ"O6���-Z%Y~�m�Έ�ٔ"O���dQ�4�R-^( ��,�"Ol�P��K�9R*��q�?p��Y�"OňU�D�K�%q�	A�J!<��"Ot�4ƚ%*�����BQ�"O�I1'D6ب�U&<Q��Q�"Od��Q�#���`H�hD�d�"O��2��,_��飓̺/��"Otp�^bN�]�F î�,Y�"O@}�S�m*DO�a���'"O�@����5	����=)~��˱"Ot�FnZ�C_@�q%��?E@�q"O�8 q�&0��$H��Ϫ/.p�"OB	�S̘ZnЬ�f瓾Ar� �"OX�#�^ ^�@Zf�[l��)�%"O��:��^P ���%�:Һ`S�"On�R��]�i����T'ʡ,���Xw"Oj�!g�ǶFy��6�L{�jd�2"O�E�iS�T�+MW�LzBQ;1"O��	�"@JTl�r�ʑ�k�-�F"O��Տ3�N�����2���ad"O"\�Ъ&,�.����Y�d<��"O��#gT1[A�ts�-C(ر�G"O���i�.g�Q ���
�8D�$"O$���YV�t�`�O_:���"O�ш��_�f��S%��Q��!�7"O�8�Uo@�'1"������	�"O�фd=5:.� �)zR�m�"ONU�2�[���/GQRw"O��c�傚!�V$�n�,k�*t�"O$$���!󍛼7�T�a@"Oh�����E_��s,ڈl��݀'"O�hL{��e��*�<.��I�"O�����sX��j�L-],ѫ�"O�,
@��v�+��Dd%ܹ� "O��z�C�2/�xa���,>��d"O�`C���?���4nQ�n) t#�"O6t�UHӡB��\[�-�TC�mh"O�I�a(��z��V6���J1"Opy!��չ}&@�Q��џp� � "OPY���CL��b7�?!�J��"O�5��Bh�(t3��_�9����"O��c�Y� >~x{�C7pP=!"O� !�o?^���,ޭ[Ţ�Q�<)��*=N�5��`1(@��a�D�<Y�(6=�1`ըڰ6.9[��Bk�<��]9����)B,@Č�R�bOg�<�K��8�����j1�h�e�<� ��zf	�,���1Aʅ{��<�'"O@p��M���*�U@
���u"O���/��0�I�u�TJ�Љ"Of�z�	�j KQ�h��z�����yrC���	�b�Tx��
���yRJ��)�`�C�Ð�Ϥa&���y�Lёye<ٷ$؀4���D���y��,)e$���K.n��xt��"�y�c�7wF9��BM#/� �%��y���*q
��7-���L�I��Pyr��
U�Ϙ�&���%l�<��F</�H�r�C�mN���sC]�<���<_>ݛ#hZ���"��@�<Y�N'�~�PE��g�Ƚ���L}�<a���J�]a�9>Q&����G{�<��b�1O~̱��Y�v.��tʛP�<I $/T��c���k�"�JG �e�<i��8��Y�D�ƞ+�nI
D�Vd�<Q�aT
Q�d��&
ě*ޞ�A�Z\�<Y5�@���H����r�TY"%�c�<ab�3;|Ma��hT�񸣬a�<1��<� U��d|E�K@ ߍa�!�d�%8-61Y�#�,P��/Ӄ*�!�$sH݀��s��S�"C�!�$�*:`�Fm�'SzD��ʠ�!��d�*1�we=�h�9,[�C�!�D��hzR�P�B�d�4�c��+a�!�Ĕ�s︘�U	M�vd�a֪�+�!�d����@#@@����5J�#�!�dUGF�����k���#BY��!��=tl��Ѕ�����B�@s!���zD����\K��|XAH}m!�$(��!�� H����B&M=m\!�_- ݹ'��4*x<����M&MU!�2����(UgX�@�!e�!�$֮hmt�Ղ?Br�@�"�.f!�_�*NT�#&%�F�aD��!��l@r�2N9L�B�	�"J�V�!�D3?J���=
HԵ�@�Ԫ8!��
m��
%��!!����Ⱥ!�D�'��coׅ?t���l!�D�0?�U�`*M{�{qⅱ!�D@�$LEbqL�C�[���5!��:mQ�`���4N>���ہ!�dԖ+褡���0,�(X��..!��aZ)��gQ
8_a�V�
-!��C�<�U�R�^^��y�� �!�Z�s\|�����
�0�l�
4�!򤘶0iB�
���4�6�0�JC�!�&$zv9��!]�8: �Ĺ&a!�Dƌ!��!��RDG1�W�H(h�!�J�Mzu[�*ށ�:y��D�!�Āp�D��6JɫS�p�9B���!��؜d�$r-�18F`�Q+��Z�!��49�# .ȳ]B�}
#ʔ, %!�ĝ�$rd�ÄT9T`C��H!�D�	�su�ݢ.��@��d#!�D�:������c��m#�[#�!��ct�B$� .�e���ɬO�!��`LI�$A�u�9���&�!�� e���K�J,Ɍ�񐭁!Y�!�d�"pS�hQ2�P*`��@�%G?u;!���!���-�j 5�X]!�D�XЎ�1��K�.����E�
!�� �U�G��.`�yBO�Ux�ٴ"Ov����h/>� �,J�28�d��"O����l�\6
�o,�J"OF�{�^<H���{���{q8��"O���5��.���p&�������"O�-ZB�����(��!���b�"Ot�Ѳ]1}��V�:g��d֕�yB'�-D=��~���ۓ(��y�+�:V����ƒE)r�2�,
9�y��)VF.TZw!�<� J˘<�y�i��2}��FH-@0�i��%�yr��f���v�B�m�d*��E�y��̙�,q�'�h
��;�gݏ�yB��1�H�6�_$
%9u�)�y"��5=���(�6[ՆM�!�=�y���#L����Y�R:`m�d䕧�y���-�����P��m�`K�y�녣Ki���F�!A�6�1R��,�y��!]�$r���$��@�1lW��y��:i��	�/[�H�0
1�D��y�Eu:	�GQ+3T���l��y�j��h�������S�Rx�P�̌�y�M)����A�DDx�G*B�yr�ԲWV��W�P�%���Ӧ���yӗ[ �x���	B���٤�y�N�9=O�$�օK��	�!����y�`85.h�;�㜩Lr;��� �y�`^�O��u�7�G�D�ҍ�F���yRȇ9"k���ɣ7$ԙE��y��mDAr��ω)	:Aڲ�M��y"�T:xU�pM�,Y�qC듬�y"�şZ�����+0`���y2I�׊Ɋ��ωO< 	2���yR&E$;��vA9b�680
	��y��Y���!+�jܴ	��p9����y䗍i=�|�Ak��ގB�ƀ#�y�d�6v*% Po_�u�<H	�A��y�T)E9TI!���o\�U�K ��yj;^M�ak�V�w^vݨV����y�h@4������,�|�ӀdV��y���4I>��+R��(��0�y�h=p���5O����]x��]��y��(p}B��$�r0Xm�4'���y�dG��(���+y����T:�y�$�	J��3�]�i�<*.��y+�5o�9�G�>���k���y�b�,���I�7�ACh��y@R*�#� C4��kuE���y�d�R�o
�t��m��%�l��ȓ	M^U�W�΢SB�:�A��8��t�ȓy"�%�v�1�Xy��F|)���/X� ��D3����Ֆ#��x�ȓ7���4g�,}�LY��P'j���l"҅H�@Ħk�6pBf��6<��:��xp��u�0�!�D�g�R�ȓVS2M�ѧ�i�@(èL�쐅ȓ`V8ѵ���©���lt�ȓ.r��
CK�D��G��YZ����<������5���t�UO%
��1��xs6�M5$�|��I3n�&��ȓQf��Z�^�t�\�h�VE��"�\5��!¨8�������be8�8��]�WZ�8.V.����Q>hd"ńN�'%ԨP���T��5��S�? Fie[;.�2mذ�Ǡ\D���"Oj���@X&H"�(��P0v��u��"O ��R�&Z�p8�楈�c��@"Opz�⎩Z�����@1)��ĳ�"O�l���N�:��D���6t�!�"O���s���B9�J��n�`D�"OHf�֝e���蚺0#,:�"Oj��1m΋^�.P#b��6́�W"O9Sn7~��!�#L�T�nȺ�"O8LЧk2J|��6{�Ȉ��"O�2}׈�X��"�(!��"OZ`�V)FZ��$�	�C���Bd"O����o��2Y�)��I��}�F��B"O~}�[�d���_�m�Mb�"O�}�"�8� �vύ �0���"O*%q㥟�( �d`���89\!�"Oh|hFJܨE�"�y��\?$���"OH�v�<k�A��ҳ6�ۧ"O�Bš�r��y#�&O�U�'"O�u�T�ڶV4h$� ��)ֱ�a"O��q�Ɂ0�r�`��L�y���"O����;-�u8��7�7"O�U �p��e����;"O�b����ʌ���ʃd��|��"O꨸@i�
i;|8$*�8B��c�"Oĭ)��}�څ(T �&�K�"Opi��G�h�#.�;H�E�u"O=se�ʨ`�x)Q�U0>�%�r"O�b�T,:�s��� ��p"O�H  `͢�ٓ�!��N����"O�y�!K�#8��J�MBE\��"O��K�� �g �2+�[-
��""O|�y1�ɮlH�����T)z��"O詓M�PgT����e	DK"O����9Fa����?!1�"O��bm����� &�`(�"O�ŀ�HͳU%���	�=��U�"Oй��[(,�4�iQ�_'c�����"O�Q�ܪv5�\� N��"����2"OL��P�H�OW\40׌���"O��еG\�m�ne1��83��"O���/�c�\a;`�ߞn(J��"O�M�edý[(��>.lĐ
�"O� ������H�C��Z
BK�eAC"OxK��%Ml��(�N�=ۂ sc"O�9�mU��0��$G2c�����"O�tp6"�mz�����(A�΍!$"Oذ�f�4]~
��!��.l�� ��"Of�˥�� Na�`Z��	�W"Or�Î ��8@!�̖Hp)��"Oܸq!D���VP�Ui�<e���w"O����"��
�6��a�F;O�By�P"OH���ש_�����oN���Xkd"O��3O�o��|�s�ެu��$�0"O&eA��@U|��^2V�P���"O�	7EH�,������tt�8�"O$3$��.�d�a $��x����"O�,�c�ޡ��,�RcJ�z�\ �"O(�BI3r����A�Bb���"Oظ�E�����b@�w@�+�"O:�(4π�(�f��b�=09ڐ�"Ob,�c��=�T�E��LÌ��"O�i���̒�v��I�Z�p{Q"OH��#>&�ƄYt��+���"O� v��ԏǭ	�^�BE��s�^��"O�-�J�v�~���d��<��"OZ�ǌN,���c�.9��H "O�A�d��{�|��g��;��]X�"OԘׇ��	�U�P�[2;�ڼ�"O��H�GV�i�t��1!T�{�@x�W"O^��+��.�B��`*b^����"Oڰ	�E�k�"�zrA�`�>�p�"Op�
�(w,���G@		@B���"O��� n��69
���j>��"�"OJ�����[�4uY��� s+��P"O~�G���$�����b�aѱ"O���m�4I�);%�+#�L�"O�l���`��y���.)���2�"OY"D�,i�(=�׀��2���"OX��4.YC)���f ߁_�����"O�xJ��8�D�Ѳ�Y� ��"O�q�p���";�Y۵iɴ5��)U"O�u����E_L���f�rI��"O޸�рD�� p��<?�Z\+p*O���� ƀ%����0&�MД��	�'���ʶŗM ���f�Eƙr�'�D1��J�P�ܐ��Kr�^�c�'����q��7�-R�i_�d�* )�'��Q�!^ܭ�wFE�d���h�'��IXj_��1{ �7_
P1��';j�(�a�@�z\A`EC2Sz�UH
�'����R�J�x���i�I�^��'���Z#K�~��I����'Iz�"�R8,*@C�%Ѭ:���+�'z�Qp�~z|:�i�-�Ṇ�'���� Qd  �pa�)�&�H�'h�ab���r<1��$�Zy��'�lqH��8T����D	x���'��yQ���0�z�0���!
Z��h	�'�b���aA�G�@u�h�I�U{	�'p�&A�*����!�c��{
�'VZ�;�ሽI�fh���F\V^��	�'��ȇ�F)0�v���b�!J��d�
�'s<r�Q�I?zy��ǒ@��
�'����.@�X����j1b�Љ2�'1���DV�%��*�圽j�4�z�'�EXeG��j����Фޞ��'Oxd8�χ�L��hwo�:r!���'>`�3d
�\��H�Ke5v��'�H=i��&����LD
u,���'�.B�mF�^x4�#�gS�x�h���'�,H{�i��ga��ӕ&�!�;�'GN�3Q	�ZR��Ԍ�,m����'FX�c���.P��m3|m�Ej
�'QZ��1�K�(c� �Bݚ)E�8�	�'jd@����p5n9���5���'D����1�|�p6cW ZHH��'�bm�1ω>ej-�ŉй~xx���'��aMM�z��#�k�\=�'��u�P�T�� #3g��j��a��'��U�R0�=sj��g�����'{�T*�HݗXv�Ae$�0fn�9�'Wp)���G�L<��B�=�2	x�'Ty1�(O�n��P��$tZ|��'z��BC��378u8�)�)tQ̙��'�dA�T��P�T��wL��j�r��'n�!����m��Y�&�e�����'��3��.�@|�VoO�]���� �����\����'�q���)3"Ox���,P�z��S>�\Y��"O�ՠ "h��*�CcF�ҳ"Oh�5�ِv�J�����/Fk"�)�"O��a�v�"�p�J��p�=(p"O�	�3�i" �ȲKS�`�d���"Oē��$��Y�	�,뼘�@"O�M�Ѓ!���"�Բ1$� "OHݻ��4PE:1�k]'��;3"O"H���G���5�@��(��ȳ�"O���bk�$egh��bH�3�J�b�"O�P�����+�-�0AI��>Ta"O�];W��&W�8�#� �+
��D�U"O�=Rrh�+d� �C�a٩ZԬ�6"O΄�e%>FB�-��ډU� P�"Od8X!e�.���	�J�4p0"O�آ�]&B����p��Z�z��"O^=��*_�?e,�p��Ӈy�p�"O�qf].a�N���ҵ�t��"Ofx��d�2mVRQ�6BU�8�U"O��K&	�BP�җ++5�:�Ap"O&´ˆ	�HȘ���)9���)"O�iS�Q�3�\%c���W��U(C"OXh&+�V�C�_� 2`�A"OdؓDB��/���r��:;X�+6"OquC�9�θä�H;_�Rœ""O(L�4gWD�� ,g��d�""Od��$�N�.���"�*�#��@�!"O��P,3w�2Q����B�� h�"O�A�L[�@�4p)�ǎ-�tBC"O�UB��'�(�"ɛ�Ya�8��"O�R2�0a�&�c'�i�vy�"Oj�(��,,���T��!
�@�4"Oޝ	¯�<��0R�>��A"O� �u�]����A�6�V��"O�0h��P8=%0e���.%*֝�%"O���dփ`�hUIaA��."jr"OJѠF�wV��������E"O���D�P|I��\v��"O�%I���N��dK.M08Sp"O���Tf�0S�`��{<�L�"O2�B+L�b�[5��`3"OD�qM���ȸ�T�!B��Z"Ot %� H���D@�p�u�"O|�<g' �0.�';MHq"O���n�^���FȦB�>4��"O~��`�������I6�@��"O4�p7#�)hNY�����<��%"O��3Ō8������c��hC�"O�H�v�B�RD�q$U��$�"O�����>+r��2&�\,C��Lb�"O\��.�+�a�ԂU�K�� "O���V&v(�JT�٧?q�T��"O:�0��P�'�֩pb<g�T�"OT9��/��#�f "W�rIxyJ�"O��0RN� �����)�1%"O-�V�t|ޠs��P�xe @A�"O��÷���[x�qaoK�1}�[@"O�]�WK͓�xE�D�r����"ORa;�@P� W��q�.ʴPc
���"O�R ��*�lM @���D]����"O¸��H�6w�8I@UK�&!U��`"O��e���	k�%Zs�vR�5:�"O�iP�G;�D�3�׸{�DI�"O� ��Y��&> q��e�	��q�"O.����Y�8�@U��
F�^� "Oޜ��ƚy����)��bg��"Oܥ�Ɵ ���2e�þ]�h�"O��F�E
D��M��a̓C��Iq"O$4�Q��x��YQ��Y���I�"O�tJ���B�y�N�# #�U�C"O�	[V�(p�P� �t$��"O���v�A�+�PQ��H�;���"O$:r���7s�\B�%�F�Xi�1"O8PUȊ;s��]�r��}�n��a"Oh��c�9@8��5#�+.r��4"O�X����BUv-	��O;0�b)�V"Oz<;�)\��p�$�ѭV��l�v"OF̺6!��} JP�*�44���"Oz��2/F��i9VR+�0zW"O����Ke�R��0�ξQ�h��"O��ȅ��lh�Ŋ1x�5xP"O��qB��	!d)�Pő�j��lb"Or,��XjpQKpc�_r�dr`"O~$`���0qΘ�9�E_�L1�"On���0���a˜�$g��Ф"O�t�w��,(b1ڑ�
�X�t"Oz9�U�#y�h1�4���Z���e"O(Y��L�Π�����Y���	R"O��ei[�]��9��H�
jf8�"O�� �O
e>8�CŲQ�L��"O�����d�^�zƄ�F�v�J�"O�yآmP&b��)�!Uef��0"O�M���1Z!A�RV8�2"OF];u����m�&���8R>�c�"O���7Ov��2gC�B�$1�%"O��G��/<�h1�*a!�0�!�P5 ܨ$Y��"��,)���G}!��< ϖa�6B �*���wL�E�!�D�T��#���B,:��G�B>L!�d�$`4��@�B�$�`k_�A�!�d�y��Y#��M/Hd-��)ݦP!��/�	������V݁T�!�d�)!�r�cU`؟y��z�&�j�!�E�K�5��m?��z�!�$���dy���@�n�l�r�!ݕ;�!򤁞&��,*�� Af��!�/�*�!�dǰu��������V���B�2^!�b@��HP)�,N�tUz�ۆEB!����M��L�=���'̘!򄄤S7��8uF&d�6�Q3YZ!�۱��l����w.0�T�ߛ(!�D�,&�#���<�X�@��0 !��.;��*��{PK���G!�Dgtn$��BL�� :&��OU!�$X&�@-'�Ւ��=8�HL�'$!�D�0�R,kF�rQ�"R	�G!򄆠�@�R�:ޱZ6˟�	*!�_4*f
m"��Py��'�!��ɤ��{b��2,�x��1����!���\�t�X�B��~�`���gѼ
�!��3�LAZP�Џ��h1���!�,w��]Yf���o ����H�!��ۚ@�����Q�Q�L��q�I� �!�I�@O~P��̊�H�y1�0|�!�!'~��0�:T�����m{!��� �%ʅ/�Np����0w�!�@p+X��a����u 	qQ!�� @��ᖘf���q`U�G��u:S"O9e�ςv
*a���.-,��"O� �CꝸGM�a"���g�l�ZC"OV)��.�=��8�ծ�&J�I�"O��� �.x���*��ҙBɸ�Q"O��XqAP+j����� rc��1"O�|q¥W�W:f��F���|f��S�"Ot����V/ F�	�bd�Z||��"O���F(���\5rFD\9qLZ"OZ ��ϴH�83���ZuN!R&"Oƽ���-LąI�R�����^�<�� 2O����Vu���]�<��-M�5$�����ۃY�\#g���<	�*e���s�V�ni��:��{�<�5�
�$�*Tc�E%} UB�<�sE�9,Ι+��:n�6����A�<��g�"lJnYybDW�t ꓡ�{�<1��K����YQ��N�t�&*S�<aS��oID��b��`K�4S&�u�<�!OGX3��U.�~5JLV��X�<�'�Z�.[U�$HӈQ���!�@Q�<��Bφ~��!te ��-I�	�C�<a6㌊�,k�� ⌵8p�
A�<A *��onx*GN E|hUc�|�<�����p����;%��98��Gc�<�U�7���f��^3p�F��]�<)#��0,��܀�Ě�\mrE�vIV�<�S�&�B��pJٞ��+��*D�$�T��C�N,뗠�	��0�c+D��pQ�$��SI�qb�K�6D�,{����xBp@��C�	*D���Gi ,��{C'	*�p��g4D��s��	�nؐpYE��#,���f�<D�XF/M��r�,1=\�` �E:D��C��R�R|���&�;sl�"5�6D����$j�pU��e�`ي�)6I3D��:v�]M��@��h��vG��Xpi/D���5j� 4 ��1]<y0Q�,D��{�	� O�$���[�^1�ѡ5�+D��J�o֚Ch)���'7=�u�5�*D����ڻs1�蟇HcNaF=D�L��c�!���rE!msZ��p&<D�L�k�vn`����W3-��8�f8D� Z�쐄E���+�%V�W���p�4D�L�q�N6�D����S*{�\�Ro6D�x�fg.q@`�1�	v�< cFK/D������Б����]J�(��yr��=f8�#q"Q#2��$�4�y2���(�D1�EOP��H��v�Y�yҍ�FT��+G�Y�t���ɥ͎�yr�E�2(Lk5��5��Buǎ��y�o D�: ��a�1^ԡq���y��m��!I�D��.�Ll兪�y��Ŕ=�P����XB�%�た4�y��<gJ �A���XFk�$�yrɇQp@�z4,÷n �����2�yBhD+6E����&m/FI�c�W�yBL�F�ȶ��)b0r	�b�,�y�ʀ{^��T�²XyKBCZ.�y��M5[�:1(\rx��%�6����ȓm�x��D�H�-4��"��Ӌ��D��/��,�aH��
L���[h��ȓ�v��ՍA�tq�c���9�ȓ]:mK j?+��IC9�)��S�? �A#�)tp�< S�!�yQ"O��r�ЫE�����\�\���)&"ON���Ǆ��Q���ʹBdM١"Oxe�V��&`�D`A����T��"O�1Y5)���`�1�Q�r�<��"OB�e��' =�v�ԕ	B��p"O,�a�iĶ#%0L�T�@.��<��"O�|�!,�*t� 1��̴]�fP�"O�Y8�Mb��l�D�$;�$e#F"O��:�kSB���I��sS��h�"O�d�D�ۙJ �e�
���P!��"O.�u$U+l<��jM����W"Oz���9܌أGR�$m�hC�"O�Q�7,��]Q�Ϸ2N�I��"OL(�&,��Dxؓ�!	3��Ȱ"ONT�%���H2���c@�x0�"O.�$	�~�LQ�EM%k ��q�"OX	B��o�h}X�ߓ>H]+�"Of�1�%�
E>��v��8e�d*�"Ol��T�Tޥe㈶PO�0p"O�5����<
8� �g[�8�"Od�F$�n��KY{(�#2"O��0$��-�m�J��x^̜J�"O��`GK�*?9�-;�铪f��؂"O:t���� ix���(�4w8�{�"O"-pBc�
S�cn	�}�j#7"O:E!B��@����1M�sw>c�"O0�hE��;k����"R,v>Q��"O� ���HBf�顮���8��"O���efD0:s�A�ԉc�pv"O��caK��W�9Q)�7)���3�"Ol$a��G�)/����jMt��"O"�� c���$y ��PR�"O�E�QeݥC5��c�+><�� D"O�L��Ǿ��a���26x�Q"O<��#��_��${D�Rw|�H"O�E@�a�2:�6 �E�уxŎQY�"O�����6մ�d�]�%��Y�T"O�q02"]�(��%᥹��!��y�)!0i�Ј��\>DQ:��$�4�y�"�}����Ldp	X�ǿ�y����Iv@���[�V��� �y�B5�]���D�w��zV��y���0��a@�sPB9�^��y�(ӌ]5��*۞n�,��"��yrm��^0dP�ү^�t���j��R�yRG7B��1��)C�աf��4�yҥY�vr��W���K`��DC�>�y��ķaҊyrք��*m)͜��yR�
#��؛,L'l��t��'�yrlRw�"T�a+S��P��m>�y«=��HpE�:|�`y ��y�/˨K���	��op=�q���*��~�O$���k�4\�� �Al����4�PxRk�)�
�p'dN&0��ā�̢�y���V"��[n9:˦Q��ΒȰ?i�'U@��f�� �y�Ü�/,�W,�/�S�'�8��?3_2I�`��.&��݅��F�IYy���Xټ��G k�4��c��yB�ԖLl%IH͈d�r�ը��?A�40�@E`��(N���a�ǊG
�z���'������ׄG
5'�,{gɋ6e�.}��L8��{���Ob�d3�����9 2!�6ZM  ��'�~D��	�O�m������29�C�O�O�(�d<lO�ӧ� �]�F�!y���Z�_�\�C�"O��	U� !����g]N�L����Q>9�G����Jw'N�s��X��>�y"��Q%�Of���x��V�e����<D���R��(����J�*}�IJf$8D�"fd�r՘��ĝ���14��<�R���w�҆s�<\ �H��g�*e��'#�OH�?9f�T��2�����T����x�'����ŦU0P�Ӓ9���eD(Q��y�n�O��=E���E�;�Ą@뛜 �`�DMا˱Od�=%>M�1��27�^�@4��	}P�	 �':D�Tz �͈\�5Y���^���9D�D���;�����Z:<�X�jw#1D��ڡ�Ì9��}hT�U^T��e1D�DQB��vR����Ps<��/=D���En��Q��G��+,t����jy���I�Qp�%s$�؏y��Lp����.B�	cv�YC����T-��1�	�>�B��EX����
O��m��<W��C�ɻQ��ݢ�HлT�t�襥�*,�C��!Vyҹ82�MNՆ��gZ+ΓO��
ۓ��HfK��#��Q��3l��I�� <��[Un��'��D��*X0w!y�ȓ"݉$���/�h���Բ��E~��	�?%rg�!(AV��P��tA�š"D�<JD	�W��Z���~�(�!"D����$��1�t�c�R�J,�����!�O
�"���B�I� c�v�a#����R�'��E{��D�t��R$B�Z��Is�u�!�i��p�+�8u�0C�!�����0�E��X��9 Fƀm�!�đ�I��xe�˱�p�샚�!���t��Zb�H}���f�W>h/�{���ۈ�Q�b� i�l�G�3�a}B�>�n�8�e�E��y�-8�nK|��&��P�J�K4��!Ȏ�����:D��@�D2 rĵ3R�Y1��i+��8D��v�¦i��I����8�]*��*D�|"7,A]��]�f��(t�j	c�)D� CfC+3#����E�/�@a�c'�ɢm"Q���	�A�91>���;����"O�EI�A�\�x���(�r�@��fX��⧁
�|TC o�(J�dȲc�(D�$���]�-��ۑiY�x=�VeK�{��@��f-!�^l�8�١��vW�z����� �Lسi�1\H���	�,:!�$��]�<1�L�	7��2EV*h�OD�x�y��)*���$�&wXI����6l!�d��>6�Xt�E6Q�n����γt[��/�S�O�
���I�CA��z#K²S�L�r�'tq��+���8+b�Nb�T���'��:�� 5���@4D�'�Щ�'������:)����æ� �\+�'�t�rҰHJ�����M��i�
�'��0R!��j�\4h3$W�}/�9
�'�z�3r��%)L��2��
u����N<���p=1%J���y�#ؙ &��j��p�<)GeZ+L�h�I�c��BR��P̓��=Q�!���e�c��8m���z6JA�'?�J�M\O��$�"��Xx�ϸ�<��	6jJ.dy�+Ͽ<�v���`,v�O2��dҝ��!���r�����+��'�}��+�,�?��)B*��Q�>���#D�t;��Qi��"�Q>F�FpB��5D�� F����ۓZ� ������[V"O���� t(��;�ȃ,@`�Е�'~��T�3�߲^�r����λ/�jТ�p�v�=E��4]Jrɐ���T��QᏱZ�%��F{�����8ht�z��?h�f�ص��y2�L�F�dY˲"­N�xՇ���'k�!��ɘ7`܍���2QX7�U6�bC䉛7�*�P�DR�~��tk���N�$#<�ϓv���l�P�H��i�>o
-��I�B��d�i;��b*�,�
��A���{��O���E,��qv~)ȅ�_�(=HQ�'u���
�����@��b@W��A��1�Ob��z�h=ڇGL�f @�&�V!���Ily��O��x'�P�3 �6xOV@chRzw�J�M6D�p@1ͧ&�p]ҕk�+T��]h�i���'�ɧ���
,V6Э�s��<���d.��-!�Ě#�$�&�����H���;�p�=E��'ϰ�ا�I]�ݸ3�;d��'6r y���-���3B� X����'�V}��R9�����B9��"	�'��(�f�6=�<�����D�@��'�j:�ʇtD� �D�g��j	�'ʬ��+��D?N���m�0s�[
�'���`H�.6V��Y���`.�'��pIg��5�`s��WJ���'$P���-Ŋ&;D�y�����s��?A,O����K�W	4�Y�iB�9o��c�)LO��aƼ}��V�	MQ&I��"O>h ��~�IV�/`OH�G"O�E/����$�RU���
-#�I���'���58c�� )�'�LФ���2-!�D�-A��A�B$E f�f��Q�*(���u����?Y�J-{���S�R�Նw�T�'��	1+�^�ɔcN�^Q�CAǆm$Fc�"BN�<AO<��O^�Pw
C� V����N�<y,dc�1�p)t��Y����J
�Zh�ㆂƙj��B�/�Z]�E�+N�*x�qd��gC�C�I��
�*� Rw"؁��j�vC�	�cA|��DV��,H�����A�Z��3����`��4R�l�U@͘Jp�U���N�	�b���e����E�@*��<.���#}W���!�3J|d[��[��T�� �O��`n$�@B�7����5�L���'��ubώ��I	3n�����'��lФ��(P��̚W*��H�'C��!��(5�)G�}\^�
ד��'��5�"b��~��8F
H}�v�9�'���3�V�eJ�`���C�LĈ�"OF��p��)n��p�U%F�e��"O�c�o�xYF�`.����"OtYpq%
!@1
��K�����'v���R"_"$��a���JEO"D��JVkŚ:d����U�Lj�}�����Dp���S7�V�p!�A�N�xaP�\�Q�C䉦>�2�G,p�u\vϰC�ɗ{Wt���%Ҳ^�X1�W";�C�IP�PE2 �ϠW|��v*���C䉓b�\5:3�$J�*� ���Hg�C䉤O��WL ����*9i�C��R�h�>u��}��NBq�()Q"O�X�TE�E�ҵh�-� h0�!"OV�y
�J��8+W�DXJ�hB$"O��F���M�k�M㲭��"Olx�tV-k��0���2L���"O� >�dI�h:U�#Ä?T����R"O<���64��b4~�4F"O�04T�)ht�ǁy�~u�D"Od�C&O�jU����
*r��ys"O�Y�nTkpe�T�eǨ}�q"O,lk��^!f�b�ss��~m27"O���W���Xm���#y61b�"O4DR�>G�#F��j�LA�"On���L��PWN�cH�-:�|�3b"O:�a�#V4��h��G&��"3"O2�˲/��q{�=ۑ��C��b "O
�32f݊ S�&B,��"O��J'�_<� ��T�O��C#"O���犫&Y����o�(R18���"O~Q�!��-)8�*4@R�D��(��"ON�yQ��F
AR6O� �^��B"O��gmK�!�<y����Os8��2"O�<��d�	J<��"r��:Gs��*�"O�iz4��E[��ɤ�70ZY"3"O�Lڳ���Y��@eN�S�L�$"O mR@Q~��j�L��S���!�"OF2���#}V��X�I�CR��q"O�@��Q�-�l�xcܳq��qW"O`��&�
�@Q�h���e�aŞw�<a��*ۢ�v��<!�j"��l̓.�1��DE�B͋�g�P��<)���/wEy��J�P�`E�d�<��D��L�bB�$����g�<Iǈ�x��lI����s���^w�<��1w;�%�d�,w	�Qc�%d�<1���hma�b�*R�ԥ�uC�h�<���>/�`QgG� En��J`�<!�m
�_M�!8�j�<\�M�l=D��;CN %\h��X���yn.D���":\-2B��J{�mp�+.D�4�2 ������'FҌ�s!.D�H�2��d�
�r�o	�<��<9%�2D���Ģ� �v1ZէM�-"�@`*D��C�x�@,�ưl�[&%D���aN%�e�!�+κ�c�@ D���c���c�Y@�ý�p� ��=D�HiP�\�;������Nv�Kg;D�����.c��b�ꙇ3x0�ڤ�%D� �ߔY yjR�I�<
`2�I/D�4h"�<?�&��\�u�W�*D�h�v ��Q�
����	_��!�%�=D�*`�J&��i����gb&D�AQg6$�|�3hN�rC���0%s��HȦ�[�n}�!GN�<E��4� ��q#R pl0��#BOOG����z�.�1�P{rŉ�+@�bG�ت����7A�	�8VD�-��O�1�ta@?.����b�<3�*aAE�'w��#��V��!�4��z.HI�e̤y��T���A��,[���T؟,�rh
���U��*�,/����R�<�	�6������ +(��-+m�� ��ڜp��K.Y1�xe_%B%��(�"O$��5��u��mI&�B0��0+RZ�ZiG�Y�g��5 DC+�Q>��;O��h� �gv�� �67%�<�'"O�2[E�vA@Ҭ�0)$��J�/r�Ex��'ʔC�R=���;ړ;RVi���:<݆�HZ�g0
=��I:=߀�:D��d7!�S�U�>+���n@�^2�a��	w��ӂ"� �5�'�zp���m�^���g�2�F58J>���3�J- ��5�L�&}y�<�0I�~�t
�Y
�p�t�Bgzy�g��I�<�]�U4�k�!��N3�xkM.c��%`�=r���É�T�4�&�=�)	�W�<�λ~Ǧ�ـJ�N1ХU8&��)j���ЁƓ���ub���d���B��b(��NϏT-�q�0n+N,����A��(O��6�ؒ-���zAG<K��[��'ZԵ���B{���kl�8g�r� h��  �@�4���'��ޭ��ć=LT)-�(�p>�P�Q#	��B�&�<UtT����T~��ͺx���31-�
$� �_"ʀ��JΫ<0�=�'
�|`�Wk�4�>���nU�l���]����+5b�Uk��C�9��p�P�M�_�*�8�^�u*��J�^��O�p0s��y7���3��iq�+C+s1�����3�x"�<2�.�y�&
�9v���L|X<�a��6���*�"��d0M�tǄ�$�A���o�'�,	�Ԧ�,@�L�
��{uʵ�Ó7b6�ЩVP����/o�`Rs��F�F�{`�ϼ?���#@��0M��X4���U�����hwJ�kwO?nT4�r��.B��	>~ޮx��j�Y�4���-ϊ|��ųW�K_��q�e؟P$Ƀ�]�u�ڄ�d�4�%0"OJ����g�����#K b\P�BD�;;���N�X1�,(��� ,B��K?m	�"��(R�/7ofA��$F�#�~��B��/7m`�RE� ��P���i�7��h��J.Tt
�� M�[��LӀ�����r'���Q�`e��<^@��D>%�tdPbF<O���b�M"�5�4c�6馡j���+$F�;�ĪB+`�hSc��*��0�F�"�U����&�-;�L����*�|��'t4,�p×!R��(3�W�&��l�]�	� 㗈!W����P��cӕt��`Pw��>(H��;��X5.��C7
��guy����Q�5�2H>q��X6�:��O�Fh��Π�y��Z�Qx��ʁ˃:@�J,R�����x��i�<ƌZ������?B]��"��A"`˦i�aX�}y��cT����0"�,�V�'����F1[�6�B��" �\��	��b�	� )�9��3 ���3�+�<y�P=�u����H0��ׄ �����hU3Xa}"��D��pXT#�,\@0�R����O �8���$���h��f��pEC� 
d�'���bÂ�J�8Dg���x��u���YQ���&�
�|eJ��ȬŖ}�p��
k&\� �f�O�xm�,ԍӓGGp�Z]���ݫ4a"��:�乀��Wo>�z䣉�V-����.�
�Y�F�(E;��K��
ۺ���$ɡi�Ndb��|�F��Uj��A��{2.]���:D�ɠk�>(yVL�|鲳͘{���J��Cf�&Y��	cpv���=Px�����ϊd�j"<Q�,�'���8��z��PcO~A��3l�ZR��3ĦP�eoZJ�<Q�L��
-�d���ӯn �%A5�ܦ-0E�Ř-S:u��-@wy���iٴA@�gC9fDq�� ��U��A
�'R`���Y���?8V���E�Ph�����9j�S�㕭?\��`ÓU�� yPM�<P�L؅HtD���		��	�q�N�s�^��/U���Ճ�͏~ 8A*t�S��Pq��{�I8�+&^��&Z�� Dx��,�4�PlF�WM�2,�2"�k&e��O^>�C"O�10⣟�[L�8�
!��d��C��Mj�|�'�%p7m�/
p�Q��O#�Nd��'�<q�bLH�sI�RÎC�?)*��`�S�-��`)��Hر�2/B�}cfE�(y��ɤ<��]�f�z��� \�=P��ʒf��m���J��!�݈���aMl������4!Ӊ�ƚ_ˬ\�f�|��tᝌK&�T&WV6�r�X,�y�%�/�R]�v��!K-�x��M�Q��$�h�Df����ēt	�s��/2�f��a���ēC��0zS�Z�L4m�u��<lw2,aw ͡2�A���HБmӡsۆ�B P�T?Q���'@�!�%��`���*�P��B��=�I�w$΃d�!��S�FjB���M�'����cEV4��'Lq�w'K.3lɧ�O'��a2��5_	v ���;v�1#�'p���E���t����
�3��p��XN�)1��(��L<ɐ���%Z'��_y���TeSYh<a��$�X��4
��t�>��Q�G��y�,UI��H�W����5�%��?2�1\Ox�5�&�D%l�ޔJ�P?XE�2�ȊGq!򄜻�`�3E�]:,��L#�o�`k!��&��
��t\HY��1T!�Ė"Ge�dI�n��W�z��r�<3�!�$ݾ=b�"$��~�`�3&�k�!���� 8� �H��L�k�C�o�!���&���z$�K&�ĬBǩ�71�!��	%L�&���c�
��G�E!�� ��Q �K�{'��#��!!�"O����%F�tP A!ǐ�L=H%�"O@!��H�>�Xm�Qhϣt �}�r�>���P�F�B��?����΂�yBfL�
R�E� $D�<Q��ß(Μ�K`��"m�y+�X$��E,Ҵ�F�q�g̓ v� �!��"Y��s��0G��4��	�s�<���,	J|e�e�T�P�L��ɑ�9Ybݺ��v���3��ކa�Sc��/��k�O#�z�Q8d�����^>	�5-֡ �w���"���` D�@Q��F5Y�X{���<`��@@%à<)0�����R�?�����bPY� B� h��+�.?D��J6�J�+袠�c݋c�lUL��a�L�'�T K�r]�'?� r%�ή�,��ƕ1Ӿ�Ic�<�O�J�FO�2Ք�!�Ϲ�^�P��K1�H��W����.>�8A��H?e�"�AK><�?�D��'�d����/[��$Ȝt��ÞG����V�ŇF�C�I�1_Nxr �]b�,�Q��/��ʓ�|��r�F>��#���9��E��@�� 򢌡�nJ+�B��? uD)�̑ {wv�"`Ȍv�L�3�By2lK�$?�Yb���y�ɯ'�&�RFG��E��`
�x�I�#�:�7�Hg̀lࢆķn4B�Q���}��y���\�Ƌ��j$-!�H�&`G����4_I�!hS�I�G��5cD(�fg�^Ԃ�x$��wB�Y�ȓ-����H�!K���h� �k�էOHi9��1X�`�O��M	���2�����"M<B��&"O��	�dU2��'���+�J���8K�����L<������(�U�_�[���g��N�<Q4���=b��L�u0�4Z`SH�<ѓĚ�&���BA:s��$�v�p�<y��ܮH�� ��ލF����1�s�<)E�Z�Z<��ϗ�$7��Z+�j�<��au��S��J  ���+͐�y�dO��RuY�AV:yox<I�)U�y�ˑ>|R�����+|u�3 D?�y	�u}j���'	?$D�[0	��ybn	�,y�T�!A�.N����ѥ�y��*�JZ2��D��5A�#_8�y臋r�����O:�"I������yR��,���#̝9;�l͂գ�+�y"��	��I��OۤC�4$Z%�V�yrA�պ���
��v�t�I��4�y2�M$,���&(�,` ��!�yR�[�|�橠�Cu*�R�[��y��:M(ʔ;��D�u]�!:  ���y @�ns�蘒�_�-�aG��yR���I<�bK?C�� �B�y�	���Ʈ?�������y����4�A�5)�6�L�0W�,�yR	��\4I``�F�)]��W�@��y��0����2�Q(����s!�E�Tu�ɵ��Ze�s�O�(y�!�$�6e�(!�`a΁K�n|��!�/�B��a�"5�$��6���[!�d���v�k5��ܡ`�P��!��ܩO�uҷ��,vw����hN	q�!�A9����̡j���pAgJ��!�H�%"��+���1�>�zv�U�!򄅮<2�=`֣S�/r����р:!�K8O���ꀯv�� Rk�P
!�DD�:������6Ha�-��䞻G+!�Y�n����]�ot�[�{/!�B�.*
�&nt���	�� !��4c�LM(���&@nH�xGč!�D({L9�T`�	�&H����O�!�� ��2V�b��)t���i��䁖"ODj��Z�;^�B	��Tp�"O��0�e�!u�6�
\�$�h�R"O@h��C��a,ŪU�/L�b�"O������$ ��QQ����YhR�jF"O�D�@��t��%+ac��hi�k�"O0इ�?!,q�B�K�L!$�h�"O�!�䞈L�(ie�܈v&d���"O�1�����w�:�(M�XF$�"O�� b��p��R@��k��Jb"Ot㦆��`Y� �׎ֈm.t�B"O� 8u�U�dV<��ը�G_b ;V"O����i։s�$XXQ��2A���g"O���T�ŜR���[k:*��4"O��z�#ki�5��,���d )�"O����쏃X��dȋ�N�,S"OXM�0䛌���q筕�Ib�e"OШ�lU&L[4բSK�	7���"O���nY�4�:X�s���6���!d"O���4`�q"��E��	#1s%"Oz��W��0fr�(�0��42dx�"O�ʦ��,�N�����y�p-�d"O$�#�ʤmjJ��ʖHtbj%"O�- `��3k �J�/١Tu����"O�����V�
4�g�E�z|z82�"O!1��J�TT1��M�0��2�"ODY���Ȇ$\I����>n�N䃲"O��R�Y�t�|�x /`:aR�"O~��X�F��3�
o<��V�#D�@#B��ĸ*�@C�] �� ,-D�0Z��J�0�'/�/ȞU#�+D�@��3]܅R@/A.!�$LH�&D� �1i�lyl��lp�|2��!D�����P��c�C�*�X�$c<D����ԙ��Ä+Ė{l��R�>D����#�.���3+''�jA�<D�� %�</��sE��2F��B׉?D���� ؠG�a3��!j�q�3D�d�*X�jYL�Z[�W5j	(d5D��ɓ.�;^���d<{�P�Cd+/D��*c���A܌I�虚��p
w�)D�4������}!����=������(D������l��(=�0��'D���v�9\�~��;�D��i"D�L��DX�u�~;��$w	��Ї�6D����S��*G^�h�{�`8D�<�d�+T��e���ՠ_'2��0�8D�����:*���Ŭ�_�T ���6D����a߶��1�CC�h,���B>T�l)�E�v�nx��J�m��"O*��g�й)��m�7��_F0�K�"O���o�d���CLA�@U i��"O�-����I+�t�P tV �;�"OvM������,@d$�eTQz"O�bqGB�T�D��	ِV�a'"O.�R���т�Bҧ��3��q"On|��Ά��DC�'�+38z�aR"Oz�ۀśW�X�C�߷L�ȓ�"OX�򓮐�O|��V΄�b
�t*�"O���XFj�AǮǱ��<Cc"O�1P�^��F����$o�+�"OJ��(C�H\[D�=x!��k"O�(s)�6�V$��(�wp`�"O. ��*��x#��=��y�'"O� �t���U�M�~�9��V��J�"OZ���2N+�`Ђ`�f� 4��"O8,i�!(wR��@�-#��$�a"O�!��. 'qn�"kO�5|���b"O��y��'mxy�0*�/eV��	�"O�@����6�!�'�>X��@�"O.��'H�1�Nɠ�-J+$� "O~Г����cw@�s@nU;}����"O���d���t12�a��],Y�R	�T"OAYB+Y/x�� ���5y��9�"O����@^�/B>PI���?��Xi�"O&�a�ƌhˤ��e �	\��0`"O(q�bꏣ4	��ZR#�"8�4�9�"OV�󆧛5F��qR�L�a�.h��"O�yG���1pPo�o�0"O�I��ʑ��hUj��I��4I��"O�RR�U���<0��"�8�i�"O����e�,q�4�A�u0��"Of��TKY�
<�
*!:����"O�;4G�1<h@���P�g����"O�1�MгJs:���
3I7���U"O\�����!g��?�<\�"O�ph�A�G.��f����"O����ŋ+_ԅ���_n��Z!"O�)���uP��"�m6n���"O0���׫!��@��L��I�"O��	3M�/VJ�� �E9)��m��"O����yV~��M:S�|��"Oʐ[�&-DD��đ-\H�9D"O4-q����F&��8��()8��{�"O��2T D�
��!ؠ�2]����"O���6�!+	���,��Eӓ"O��Μ��0�3PL
m�"a0B"O�S,�*�����.����"O�H�B���݂'Q,M�>m�"O�����V6i���7�*�� 0"O:yQDJ�w\@���_T�4Js"O��#f��U2�q&�D9����"O��������,3��4;��؊�"O$�a5c�>A^@D�ӋC�^|�"O�P�(��P�XdeI3 �2ĠC"O͐%b�36L@,�r�W(q+<��G"O,<��הVbk1Oȩ\KG�BS��j�`�|�'bt����S�I��7$ٖp4h�'V�]C��+��U�FW�/������wwpu�
��j9`��'�F�^���J$�*@Šm���.�4m�5��N���w�n�;���;BJM��F�x�!򄕎H����vH6�!�{�'�DH���4$&ɧ�O�RiS� �(K<8��K�<j9��!�'^�Q�-�zD��fʪh�\��E��u��+k�B����L<��Ϯ��=�`��	IU����	�AH<���Fs	�A�e�[-yԝZ��@/Emx�a�`^�p?��%�IBϒ�>VH䣢��RX�\��d_�Hw���O�����#<<�x�OI��\��"O<�J�_yH.aZ�O�
�"8��x���C�iH"�|��aڬO|�!���?s�fՓv�y����½��㉚yp~��!��s�.t%���Q�����2e�a�KU(T��
�o�^ن���T�s#ܵ`�@����$a�P�(��>0�U��I�3,�U��Hчu�Q���Y`R����fW�O	�P��fII3
�L�Uۄ"OZ�Վ�_� ��i&6HQg"O̭`�*� Ѷ���4{*�� �"O���-�2r��3��I5��"O� ��E�N�?�D���͍8"��]G"O�ݺ��>\�h�۲�H%[�,Tk�"OxqAd��)'m |��e�O"b�03"O�(A:n'� ��	��r��"O�	B�����l{rB�<v�� "O�D�РӌK_�3 �,��eh�"O"� @]��rɛ��$d��٘��>�O'I�.��?�0n�3�x;� ٦8��aJ6D����"S.-˪5���v  �Sȯ
*�y�H*���P�g̓8u��z��1m٨T�aBĘnɎȄ�Ɍ9p���r���ep�`��&�#Gx8�硊)��LrF�LF���Fk�>ZX^����k:��F3��p�dA)Q/�)H|���_>���9@"�8��M� �Qҵ�3D����W�>�HiV`(!|P�f.�<1��؃s������v��?���K�+(��f9��h�M.D� �`cڊ1@ҹZ�L��kTځ���
1���'P�A���.x�ϸ'Uڈ�cC_;^r��CrNd�(��3PԠ�&ی�p�����g	�sZ��Rd��x�d���'�J����<"�M�eN��'����D�f���M�: є��O�P`�b��Tjj��n�Dtj�'s,���(/V
="�(��e��)O�P���!w�R�a G\�O3N|p��'B��cb#��A6.9�ʓ{T���3�ņ@�l����nW�ȃ'����_�ou�mI�������e�2)ǥ&F���L�f4!�����Hs��ԐWI½Ȗ	�,V�tthT�6"�Bi��'����Z�0O�
�/сP7vd#
�հ�A�h�!}��'�ޙ�À�Q�P%�c��T�X�	�' I�a��t"�K��\4��H�p!ֈҦ*�:l$��?=#��ʙ�0|z��{�&!��e=D��"0'ެ�PEmȗa+�,*p٣۸'u(��1�3���d�$Ӂ���成���)y�!��ߙ[̠��i\*���6�K0�!�ę�F���9��eT� ��DF�!��B�tC> �5�S�i;bA���b�!�V#A�����?R��Po��T�!��(.�"���#(,1�.S�w�!��#�(�� �M{�d"�R�_S!��ޫ2JJ�jGn?>mJ�PtX<�!�D#Q��t;!�P8��A,J��!��[�j Z�9��˂$�^ts$�ݝsg!�$R���EH�y`T��Vc
�f
!��#� ��6yS.��iV��!�$	'�I� ˈ;0D�!���7T���
|�'�M���`�;�yB/_i����1j[�N�ءi�D� �y�ʑ�`W�����8Xb��C2�y��V^��#�Ȑ81�(i����y��(<��L��-�L�;ĥ(�yON Axv��h�?&���Y��/�y(ĝ��L��W��Z��c����ybnL>t�48%���M� B��y����h�-�C=n��/���yr�T�)��燾<�1G���y�aӴ�|a�R�_�X��=b�K� �y"%��k���p�^5(J���yB"�.�V�*�隆W��m�D��y�*"�R�t���@p�\$�@=�yBO�\?�uP ��< =R�BΗ�y� ��=�h��F�+k��@r�^3�y�/�~5�C����V��y��T�{X�]+�@ �ظ+qOZ�yB�[
{9J�⢂
9x0q��@��y�]�[K�:���< \Y��'F!�y"Z	D'�Pzեԍ�R�0�($�y
� �4s.^h��X��C��2�"O��Z�%�T,�`��k[��@"O4���WEB"�R�$]�M��EH�"ON ��흱%N��P��1`FaZ"Ol����/t�UJݴș�!"OjQ�a�,ⴑ���ՖY� qQ2"OЭJHZ�e�.��(Մc��y �"O� "��V�.&��S�⟧}���"Ob�� �J*�i��I�o�>�j"OB�BA�t�Ha�0��}���[4"O�e�����K=�a�`	J�0���g"O�X4K\�n���a�K�3I�Y��"O�C�G �ӗK��:A@�"O�R�*�/ ��s	@.ز"O�U�¦_ۦa��	��c"Ov���:+���r�b�p�@���"O�<8d��� �
����ɝ�pȠ"O� C3(�7gΠ�q���
Ū�2�"Od�Av��)]P��.�N����"O$𱐭�� q<ICc���"���0�"O q�mI.2��2��z!Fİ"O~��.�3o�!Pc��"%.:��"O�1aď���
=ȃ͏�=�1�$"O����F�zB)pb��m�"5ڡ"Om	���/��\�@(�x����"Ohuӆ��<)5��î��Arl� �"O�eq�,�H:��+O��{���b�"O\Xih��9��8d���h���C"O�ř����x�|Sf�]
Z �5r�"Oj�P.E�
-�%��4"�0�"O<ܠ����Ho�oNL1pF"O�U�T�['*D	���0,R"O~��p(љ5�(�;D�):����d�.4� �s"�
��)CJC=DK��OBቅ�K�Lh�	�����A���I�P�`J���S�gv�l�$A��)?Z􉓣�@��D-�S�O#,���M��Z���ċ+P0��ӏ�d?���AT�(N�����w1��.�S��[*" Љ�*���5� �N*�'�ў�>-jW�L�Ls���cJַ~���a��<i��>9�O���+�8A a���jS%0!)�	o���2%�S�\���I�N|c�����0�0yr��J�ǚ�J�>3�%\o?��:�~r���)�n��	�rn�4l1�pjr���ME8�0��n5�S�s��5�!>�`����d3ՖxR�Mb���OрYs�ā�V�q2�/YC�-��OV0����$T����kV5d����&�C�d9�Un�zɢ.O��,O�?�CB"�[dzEk.R��h���H|y�Qxy��(���4"�`_��s$�Y8WD�q�����'~^�DyJ|�d����yqE	ln [׆N�I
�Q�b?5(�F�{YFA1g�I�0Mァ�>�"�HJ���S&���E'
� ��p�H&K�@Y�E(�`^p��-�i?��J��~��鎀)��jc,�U�n�mV� d���c����'Ԁ���v�Q�K�cA�u�׍Ӷof��!��[����+9b��ru�V�`p� MʖN�ΓOb�=�}r�
3�:2�M�Qp�w�uyR�)�'��(�%J��{��u"�A��k�X��B����^4���%~Ț�Jf�%��"t�u>�z`GW�Te@��V���b�-�I�Ex��!�ܔrpg�5d�&�3� G�w  � �	�4  B��|M굆��{�<��ve�V��C�ɝrO&Ȉ�/N ?aZ�����Gs~B�	��mp��ʋ}�ڸ�"��cRBB�	&��*��]�MԴy���i�C��#���΅}�l��4Mލa��C�I:}ξ�V/�xDb�kRaNi��C�)� �p� �'3R��'!�����U"O�	���@eF)r��������"O4-��Aսyh�$:�o����a��"O�Ib%)߯,Z0�3NE!g�����"O����$���mZ��#s��L1"O�Y�6�3�0�ʗ�O}�h��"O �Bfď�a|����hK3q��+�"O� �߃2px9���֎aDQc "OV�#ҏL~���ǖ^d��C�"O�a�cg�0�XM�)<�J�3�"ObI2� �-g<!AƔ(@�ܻP"O�S���l6����__�蝃�"O��WO�k�qCu�ض*���`E"O�d����A�y��nW
V^�ё"O��H�;M��e�'���q-�D�b"Oሷ��&ϰ`(EH�5�"��E"O��bgi�#`��)��dJ�i��"O�A!��AV�v��"�:uE����"O�}�v�v�XJ��G�B2���"O����Φ'�
QPw�!Qr@��"O,E�Co�RL�XF��(�tX)�"O�:gfS(U�y��[[�>�yt"OpC�kQ�,�=YvG�d�(�Є"O��a��D��x7���G��1�E"O�H�� �6����Yc����"O\�B1g�,W�򵈂�>-�t��"O�1B�� �܌�t芹/���q�"O���!�VH�M� �+N�L�<��՚B�$�S�Q�pFZ�;��^S�<!�ɳc��I*�V.]w2�H��S�<��fl㐮�"@�bL'D�pq�eՇR��9��ИM�tu���(D�ģR#ފP�Υ�I�(Fi{��:D���T�2|vL��M-?A\����8D�X����6�)�Wc��B�P!�\C�I|a�C͈�M ��[��~�>C��D�� #�B#e��\PY�!�6C�-m,HE�%����(��C䉯� pp���nĔ������ ��C�	�[	Ε���)��Y�ɚ`�B�Iğ��L�melP B�m^�X��'5D�<*���7]HD� A�?/z|
7?D���eg�- 5ތ��Oߪ7v
�2��>D�H+"���*���E^�F�b�=D��*��%
0|�U#�/\ȱ"<D�(�t�664�X�c G�V��b<D�� $��0~��O�J�
a��9D�xAC�[�K��$�F'�+�`��$D���w���by�1)W�c����#D�D�Q��)~�U��I���sS
 D��Qd�Nq�8xs5�&)_��Ҍ8D�D����.m��I��J	Tp�-��k6D�<�$��L�CX~?h�V�3D����Cی=�|��T�í>���B��1D����ǋ�#���k��>����&n.D�8�6i�7�);E���kFPj�+D�$h��
$L�ְ�s
Y�`R@��c$>D��`�0Aj�c�Q"�:@kw�;D���h��(�X,цJкt��r�G8D��[��t��`i�f�$^Ƭ��6D������R������	�h���y��)D��Öj�@����EF=�nYI4!'D��p��RR�H��ӆ3w*�b%9D��P�'L0u��堡 ¤mr&�rf�7D�� ���g͐!*�p#!�n���u"OhDx�B�m�pA��%��Ѻ�"O~�qFG՘c��1�6f�$�&�)"O����
4��<�`eՋu�:87"O�8�7̏c���D
&����*O���nֵ�P1�a��_Od$�'ܖy��L�Y%e���%x6eX�'}����V�tz$�@�B%I�:�i
�'oVI��̜X}�lk3B 2(���
�'�q %CB�9��E��$�\]�
�'n��	Z5�Zq�T��M�f�!�'�,y#�uQN�ЦF��H����'�&�i�,��D����J\@�x��'s�0R�&�mm@8�K��5��(��'��5�0�^8�6-2����cAx�
�'�� ��|

`�K_G��	�'�� �T�R�l�y����XU��k
�'�rMxԄ�2(��AkEg~R����'}.xr�#cW�lځ$Я�H��'�^��娍0p`}Q�LW#4б��'��51̖/^��%��^75�@�'����=g�}��!�"D<��'��-�p�%' ����h*�h�'�����w�b� }T�P�'�6)ɅL�<�( ��'#G�}��'�0`q���~$��CB��$��'I����e*n(PS!\����+�'�����cB1V*�x1$�:�jt��'fb\;4�΂7μi�隑B���
�'x��-4T#���K��s�4�	�'BR����6/_�x��,�/]	@��	�'��ysU�Y�D�0ʡ���Z$�l��'�`���T�}C�����$�6d�	�'MZ	w �5*@�2���I<��'�axt��dO������0�E�
�'F�LzBI_K���2�T�r�l�	�'`N�p�*T�]s�P�aH&.�5 �'|��pR�C����`�(X�7o\������f�EKV�DyO��ª���y��W�l>��)�M5~���	�y�i"SP�q�'��x�8U��C���yRB۱ "dUq��h���%$]�y��3G�Q0b'C�n9��It���y�fRq���h����A��@�yrDi��D�<ip���ۙ�y�ʸ`N���M�eq���4���y��T5Z��ph�L�a�����ȿ�y��U5_rPT��/ǄJ6��0���y"��%��G�^�D6� p+��y���9,VҠ5Bv�d�B V%�y��Y�O�Z�T�;�X�ZB+��y���?�np�� �<[�P��ӹ�y2��_Q�E�OH3PŐ�bHS��y2�Z�{`X V!�7Bq�b���y��I=�f��:�E�V��8�yR��`�x؋��-늸�5���y%�@m��KeS��T�b���y��PB����GǠ>j(Q��.�yr,U�F��-{��mI��H���yҫ	�nB( �'eJ�7ۢ�j�I2�y�${�0�� �B"$�z��ʶ�y2"9L�A��
Bz��a� �y��X�nIkR��B��I��*ڷ�y���/!�����o��=�r5�� ��y
� �0S�I��;�Ĩ1tF,Br}(�"O�)Z���1O��$�4���Yw"O�Hx4Ѣ e�=���׶1�$���"OHD��K�2_�JM҄؞p���1�"O��lIؗ=7^���T��A�T"O(�3`#G��m�V��i��S�"O�ف�� �`�8��*�>�y��"O:��Ǝ�||�iu)F�r:R�Ae"OF�0�蛴Xn�YD�2RQy�"O��-�CY�E���&@>=�"OX`ap�	,V���T1^��u"O�2 .F�� $Z� �TP�"O���Eo��JF�&nH13"OС�P �v��V��m�`�y�"OR�z`Q�HA��@d��/�
��!"O��1�FM�{�Z0��o�:���S"O�h��J�k�N�*B� �����"OB��d&��Vl\8R.�0Z]�e�#"O"@:BFW�J�hMCƇ�i\����"O|����"�+�#�� �3"OBX#��?r����L�m���+p"O�]�g�8��[I�A�aڇ"O��SwᐚE;@-1)��O�tt"O"��C$�.G�����]�R��u� "OP���Y=&ܨ���	_�:�>} �"O�UCt��%�j�fH�\���
�"O`����C-F�p���P=���2�"O\�kb��7rV�1B�L-U�z��"O�0`CB�1��H!���="O��%(3�J(�� Fm�.d@u"O2-c�B@(R:�h1�-G�}� }X4"O  ӵm�s��%ا�G4)�U�"O(�j#��/�8p���$L�왴"O�<#�͜w��%�t�׫�5H2"OR� ��'����6���f�8�"OvH�-
��I�T�V�d�!p"O�)y���/������Q Ȇ�Ѕ"O*`S�C-{����qêr��5�"O�$K�H@�D����t[�)��e��"O���B�*3�")�3lZ�n&�)3"OA��#!���bȓ�o�pr�"O��A�&�G�Yv)C2iග��'������b�LM����'�t�jF
�a�li�%���Y���	�'#�( ���hXL�Ī=ͨ�#
�'� �"A�)��A�IE) )�	�'��M9��[��I�E.�%k�'oRL��⓳+X���$Z;n�1R�'!���/�0
�&$���f�~p��'6��-�7rd(�AɇYM��1�''�]�hy�t���|�p`K�'�� (WD �U;
��e��{l���'|2�K �G�X�L�@�S]�L�[	�'��A��A�S�Y[�#[��ة�'\b�!nX�d
�#��`���'1��+�JM���'S	x����'�*Sd3ּ�{#�޶g��ջ�'�.ٰ3nV,��Y6�V%+lfp
�'lp��U!��n��1�]$��� 
�'����J�e�I�����(�h�'Ȯ���A(��d�!�,>M�k�'Z��F�-8hR�;D �WJM��'
|i�  ���       �  %  �(  �1  }9  �?  F  ^L  �R  �X  $_  de  �k  �q  -x  p~  ��  ��  :�  }�  ��  �  x�  ��  ɸ  ��  3�  v�  ��  ��  p�  ��  ��  ��   Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�� |d��"O
`�(�;���8���-0��1%"Oj4��ND^[��"3/9�0|H�"OB���H��*�ʞRy=a"O�味V�!X��!&F�:J�$���"O,��a
���C�Ą�M�"O,$3%o�-���p���+Ն�:1"O��ݢ1����`���y14]2��i�<�6��{_���c�H�`�fX�$Kn�<��A̼VI�xR[�)�Ć�pඤ�ȓA5��('nߡ4�� �)˩%� ���,��r�؊b#`T�eT09���ȓ!�b��g��}�8�F��-? �ȓ
K|m�ș�VṔ���2�%�ȓ"R�X�j�4JN�1�˘X�i����̹	_�jZ��1!g��zܶ��ȓgil,*�J�
j�Ne��i�J%b���f	�(U��:���G��$Y^م�~r�� S�%T"���k\�jx�ȓ|4�1�îJb��@ӵ�ݩn�V��/[`�"�v4�R�!ʎ<��M�ȓ`:��z�ؚh�J�Z��$HY:	��H��p�m�C1��!��B:��0��EnjZA V;9����J[
2���	��4'J�EA�IVW&��~�(aZ��ӹ�>� o�Y�|�ȓ�f�A�
Ο7�H��M�$�����mޠP����/���ANXo*�ȓTv�����{ ��-7�*h��I��sB�8�8���3����ȓNe*M�悡;������X�o��!�ȓ'lj�#F�m�+R&;�|��2)n�C��0S4���T:
b���:�0!��e֊��)��ͷV��,�ȓ0�&�8#���� ع�L�����;�P�AFd���,w�6d��r�EQ�( �gVlɦ�M,H��,DP�	��|�I	$G#\�������?!��K�;�L	��<5n�qV��Y�<I4(R�)��D�⢔� ��ņA^�<�ukλ.&`�e�"y�r�,M]�<A�H  �0;r�W�[3�W�O�<�eW�Y>̹��;9j$����P}���$�=���DKFj�@{a&T�Y��Ĕ&~����3@9q0#��"^���$����'�a{҄�L�<�ۗAx�T�a���yBf\<�YWcK�rt�0����(�y�d�Ko���1�f�䈋��p=��}r�WZ+�Tfd7F]�I*�yB�
����eS�<\HْLV���$|�l#<E��0lA�է	]��� S�ب�y�"\�<d��(aD�@�b�x2i�y���;rDT���o?,�2�0�x��'���礑(1��P��.	�#F�݋	�'�2�� S�ܬ"�#Z (��Q;
�'V�P &��jw=�(�	�b-�	�'��@�.ۆ<��Y[2��Q���'�b�'��'ّ�t96��.}��{�&GI�<�X�+D���W�� e9Xĩ剘9!u)A�7�d2�Oļ*��F>|��j��o��y�w�	91L��|��O,��� C1�9�ehH6B^�����ˑM{
C�	
Z�t����o�D%��N��C�)� &U� ���6�` ʔ$R|��"Orݪ��GC*��\WM�\�d"O�٧�ۖg�"���jN 7�=�2"Od|(a���x�O��@@��ix��5G�F�d+&"�N�z����2D��
"��_�m��d�<V��Ko�L��IT�*9��Ns���9}����$=��͒x@��S�\/���fR�8�!��������ZA�Ӳ��.`�!�$1.�d!e1D(�������|B�xb@*;�����A(j�y�`dӋ�y���N�Z���#�@z �W;�y�b�&.��=��@ Tݩ�eמ�M��%�\؟��#�L,z��m$Yphhp1D��pFu�����KD�[]P(�si<D��;�+\0#�$��1o��W�0�E�ODʓ�0>	�h+70`q�g«7�>��C�Qo�<!r��-0;X		4+S�ht}(���R�<��χ O�rJ�o��@&�K�<�ET�P,Ѓ��'n�� ��O?�	��,b*\�8��T��?*G{r��6�D��Z�
���"|`\t�G2R!�D��X��0ӫW0^��y@��^�L1!򄌙(˪�+S圾.��hA���!�/� H��"��'ְ�C�����>QW�Z�m�j��`܆#�(8Em�'rўʧo��A��n�$L�1x ��
D'�y��F�q��%��
�X�+Ʀ�C�Py�ȓJ����,$²��=p�&���lǤ�����X�pqȴMK9�N\��N<��˕*8��a�QD��+�މ��v}H�!3���*l�rf�4Hc a��H�c��^�~�pɇ
�O�f8��	Y�(�x��	I-@XN��G��@�y��Pٲ��@O'Jtr���_o3�a��l>v���dN��RTH�)[0�Ȅȓ��,�@�R(1�>�����4RF����?��&�]�V4`�T9H~Mx�m�<�F�QZY�� �\�q[P���k�<�a��v�\J�O�x���3�g�~����>����f��tnҨ/4�KR�Os�<��f�,
A�B%@]�i�"��7�e�<��D(u�  $O�!��Q)��c�<q���EO���'T�1�<�V�<ya��$M����C�b��!�O�<y ���`H�`�u����s�TH�<�ƈ�/%� �bi������%��~�<q��?3�I�G�#Q�x2fA�x�<qŌ�\���� Iљ{,��"4*�p�<	��V/T	�L����7��àJA�<	pK�'}��I��@�A�ᶂ}�<���=t���RC.� M�9+�+^w�<@"�I	:�9�K��u�:�r�H�k�<9GdNahm�dnR:O��TB���j�<��F�h0�4~h�kQ��P�<�J���� ���/��d���L�<�dE��~1α#􍅮_���a�@�<9R��y(������2
��my��~�<���@��]y0�O�c��MiSHZ~�<q�MJ!��G�� Pi��;T����J\�4p2�x�H���Y2S� D�<�/̔i2�[%�@	t܈� �)*D�c�׿�qXF�1 �V� �(D��@3�U�\����Όb�b��$D�� �������<���6`���"O�e�QoT[xZe���C�r��c"OT��kLԊ�	c��#r����"O��ա����A"������-D���vʝ�!���L_�Onh��F!D����j_�}��k�͂4'�ٖ� D���S�� ��p�ƌ�1V�Xs��;D�<��
�jS���dB^3���6�8D�D gM� �\Q�猜4x��e��/#D������*Y�mx��C��Q*�I!D�\p��O�E�����瞤Ce�aX�`#D�<A��05|�(�C��T������6D��K�!Ϯ9���'�4	����f�6D�ԩa[`ؤ�a���5���2D���Ǐ/v<,�1睼2��V-<D�<0*CP��!��2�m���%D�\�#��r8��JE�ܞ�0� C#'D�8��	 @�$�zv�\�8�)?D� ����7q��8C"E�`��c�d"D�tX��,����GB~m�@@�5D�p0�k<?����V�͜x��-�7�'D��9�jٲ+��� 3d �P�B��&D�h 2��,�:��	��P�B�;��)D�PRE�J2	�%�V�#H�|�sR�4D��P��G7����1I��!f�5D���#P���#�	�c�Aqd&D�H��h��J�B���T�8L�h%D�<Z����<V�L���:��T�!D����dWK�J���r�]Pg?D��j�ރB�������>B20��/D�HIM�AL��"b�> ��bAc,D��2-�Ls^��f`F	!+r20D��jV�_+�*��@jE�qH�$�R//D�eC$.i�	��-؛@4=���8D��#7��NtH�I�~P�@�"D�t!��B��� �@�,|���2,D�p���" |���)_}��U���+D��k4M�����1BH��^�+��>D������(���' ��3WN�`�"D�$J��F�@�~�a�BXc�:b��>D��ґ�.,,�� �դ,A�pa>D��0�M:*�m����hb&�(aI9D��17�^v&��*��+4�y[rm1D�0��N��n`���c�N�X q�uG"D��� �<9��h &K��`He�>D�h8�o��ƖLh�j��N�� g!D��y�K�2�KT Tr�0�@�?D�$x�&Y+�xj��TbT` #D��p5�Q*=��)�	�BM��i!D�`�Dd�7 W�a!��~zPU���?D�ts2�U#<��lH@���0��9D����g�
� Zc��<�ZY�`�"D��{D��J0h]R0)RX�2�C��!D�x؇d�VYi&h�
��ae�"D�(�6b�+D���b��vM>PBb& D���%D�<�(�èS"~R<x��?D��/�#7� ��Q4���E�<D�\mZ�7�� C�xr��p��%D�H@aa\%:7|E��F�, p:|�D"D��J�`LLUD��ś*(D[A�?D��f#o�pB�:�Xm���W��y��Y�S4M�W(��8_�x�Ğ3�y��[��MI��	�`�uiG(���y2��*^h�#j[\7�u��$Y��y
� �L�aV�|�\Sd����4"O8"4B��<�X���7J�B}��"O���$� �2db�41���"OʭZק��+drK����Q�"O୨�'G�~�P��k�)����D�'}��'�r�'�b�'��'��']�5c��$�t�IVj��<�uc��'2�'�r�'���'���'$��'����N/6q�������3FL�T�'�R��Ml�͟��������ڟ@�	ԟ,�惈�<�E��� �cq^�@�ן4�	ßl�	ϟl�	ҟ��՟���՟��i^./��1ض.u�$���Nܟ�Iܟ�	�������	���ޟ #�N�O��=CTBO����@����h�������ϟ���ǟd��ϟ��I��Px%A�.������ԄI�V����O���	��	���iYm������,���U$X�E�QH.�}�`�Tv���I��	џd�	��0��ȟ$��ş���1g�a3�e�/k�e�b\0g�"X��ɟ����I䟈�	ҟ����p�I
.�"��ۛ ��E��F^*m=�i�	����⟰�I�d�Iޟ���@���H��t�@.nM�C��$u��4���D�	�\��ҟ���Ɵ��	��	�^S�S���p7��p��^R�x��	��T�I˟ ����������������="��T�u�ŒV8zP��e]�����������������I����ݴ�?	�4Ɔ�(ː��6�sC��Z-�m3p\�l�Iuy���OʍmZ�rU���HX2E�v9�u�,X�1*�"=?��i6Ҙ|��y҄|���yP�]p�nT��ːX�8P�kܦ}�I�Th85"�}���	�@�=��  ���cV��s�A��е"��ѬJx�<)���D.�'Z�&6'[�F�\R&���d���(u�z�ze{��6��	�Mϻ�)��L ��F�L�@ڀj��iӒ7�c��է�OȪ|9�0�y���D���aV�\���з�y�ϱa����ϭZ�ў��ǟܪB�/u�����NEP���f���'�'��7��91O>����L��T G	_lw@�#�I���֦�ش�y�P� �&�J����R�g�v��u`)?��,��l�@#ˊR�',�xIqC뀒�?��	��r���He.Q i���b����<��S��y��ؗV���$��: �,y���	�y�e��܊$���Aߴ����d	��
�����'rb�M�R���y�k��Xn�ݟ0�G�&��.��t��O�H<- %J=j�ZP�W�O9�|#�E�k�N:�y?9b`�/xQZ�>�Oi�4�ҖaY��h�k�#Z��HhB"O ��&�Ζ &\�2i�0a�7&�jN�TqP@@"�8�06�1ww:�
&�J1lĀC}�`�Ӷ%�vvF���ًa��!���%�̀�዁B�pm�� R+(�¨��M��H���ҝ<9He"����1� K⌏^�t�[�I��JMv�ao��fh� �2�	�N�!p�HNv�1�iG��'���O���wI �#5�P$8l�h�IB˶da�'��F�`�On��xR��e��e+ƃ��Y��(Z���!�M#�D�:ƛv�'�r�' �$�8�4��,���>*bu����@~n��QB������l���<9�~�j��@H�2f8��w��)o��Xr�i?��'�r](�O���OF��!:��I�.ƋtNVai�ƃ5tO|`o�֟��I�� 4.N��I�Od�d�O(��zbx��}X�id��U�Jb�M�V2%� �I$&���9��5+�e\�f�d�Q5��"-��7m�O^��p��O��d�O����O��'�?i�DR0;ovP����,�p����7��<sĖx�'��'�'�Q5z;."�2���ķ1��20И'b2�'�^���������oO/S���"DHG�ﮤ������?IN>����?��j}b@A�j�d���dU�nUZ�YBGͱ��D�Ot���O��AT����D��r���QB�!b"L�K$*�jlr6�Oj�d$�$�O �B4�i)����IƃvX��(T�EI��8��4�?	���d�5fZ��'>����?���LC�&%b��B�ձA*�dn����?��JD6ȑ��?�����6�4�!�+�#�� PCK	1f�v7��Or���5sd�$mڥ��I�O��)�R~��S�?���9TLE����������Ov|HT@=�	�?O8�a�Q�Iqdd�W♬+�����i�ޭY�En�����Ox����`�%��ӻ ��$J�H+�v���*��0�T}��4������?���?Y�'���|���
�/:eAVɓ2^�
P�����7d�v�'���'τ֝[yʟ�'9�(� N�X�Dl��`9�M<Q�(�z�B�'��ĕ����E)�&{����Ɉ�����'(�Q"�T����������oN0��U;Z�� ѮȈ�M���RX��J>���?����U�2���ړ�--U��K�}F4�ϑl�ߟl�	㟤�'��'m*A�I�ld 30����щ��=��T�,�	�x��SyR�L�oYX�S&�\�e�`�謩g��0듪?q��?9(O����Ov����OF��c`�o��T�.Vp�1ɂ��Y}��'n��'�I�Az���M|��P-r�^��5F
�	}�ia���N��V�'�"Q�p�	��Z�dIϟ��<xbE�>*��Pf�}��\,�M���?,O�i9�TU��֟��s��d	�+w�lQ��_'t^�%�֏{�.˓�?��gM�Q�������q�? a��n�?�4�ڳF�9U�pD�ёx��M�n�H'�'���ro�4�E�O�R��u��'��ظrBW�J�Ic7��T
ͻT+͎,(TAy�E�1|����$ҹA��\�C��ml�#���|z-{�(ʀ0iJiau)��u���.L/a�<��T!�l�X���3����&N�@�	��,�� -���R,I%u�Laj�"�vW��p�ї��T R�-��Y�1��|�}r�L8
��]�"�'"��'g�'r����˟t��H�,� ��c��MS�x���?�p�M�D����C�i���3ړT���Vo�-1�\�A�i��*iu8f�'�`������$��]F{o�/e��!����K�+��/]�_�a��am�?��?a.O���-C8��aTl�R��x�Q"O@�F�	p��b�Z* ���B�'������$��Nxկ;>���Slݗ �V-�$J<j�L�����?���?A\N���	ߟ�̧	2�sC�s�d٫����dFq�6���HkfX���)غ� �G�<��O�!��T�jࣀ��7����A�JI�c���I6��S�ƽy�R�ɚ���@�{-ڃ�?q��ih��7Ȱcb�%�vk-h�iVbjӔ�����9O��ScC+K�<��㌂��0��"O~�������l9깪�Ŗ�ynӢ�Ĭ<��	R�6f�V�'�[>�r�H4.�<8�`��>n����b@�'�t��Пl�ɭk&P�b��䜘p�^��?�O�ly;��T�|i�a�:Xֱ��WPϴ��T��b�|�h'�3񩄍A%ru2FaB$!���W�7�Q�k��O��<�I�O(�Q�b^xR`4(�D�B0�1�Ek�O��"~Γ/��$�{ZF��rD� .F���I)���L궫ܺR��i�C�v��͓k�J�%^�T��F�憉=���'J��:i�h�qF��-=H�Y�K��<-����W�������q�vD(�,�~����;u���u��&&[Vi�!썝M5<hQWOBonT���X=-��|�'Ń�E��>�.܂�⌣e� k�;�M�`/�)��(�O����O���<���Y�/ͺ1��l(Š�5MI�t��p����Ax����#	4!FJf�ϰ*\�a� 2�@s���a�!Rܟ̈�i��?�Μ���<� t�F�ݟ��ɬh�8�y��Aӟ\��ߟ��ɻ�u��'G�K'[�4]�����2�jw��:�原6T��I:��LT�"�� H�_���I,y�J\$�f|H *Ԃ;e�>Ě��Ľ[j0������֨�*��D�C>:�x7�Aj~�ٶb�z�&�� 2èH
�����~�K�7�?Yr�i�."=.Ol	�i�[����\��I"O�3Q������T��%�b�E���d�'-�I!@p@�	�l=�`��˘68��x-t����џ��I�8�Ɏy�
 �I۟����|A�4�Nҟ��'�3 Hz�Dj�:v�)[�k?�O~���H�m&IBc�^)<ӲJ�B&�lK���u"b!�*�p<ɒ-Y�@�ɓ|�z�D�.��*j֓{���N<	���?��ʟ(@C��f4���2lS�=����E>O�AEz�����M,���LĮC��afl��0C�̦y��4��D[q-@���O����|�p�I<I:}1C��X�BJ2h����?���3H��B�¤9i��P�n>C�.�)�j��u@��nv<��R헤��L��I�6��曧~%�$�1�S�&��sʔwfV����F8e��c���70�p����[U��~������M��iq"[>1Ҳ���<�Υ�U�.H�	j������ɟ�����Sf�'A��;%DըS*��6映2�OX�=ͧכ��hӄ����������@?_���`7�G.m
��M�����<Q��^�(�T�f"D=l7�aᰪ{�<1Q�.Z��e���ݼf;�Eq��t�<植�"���s�˻GH���Go�<I�!N�hM���A��0~�pOUj�<���_�)��JB��v22D�g�<���?eQ�+�B�T������Ub�<arȏ��Y`���Z��h�wÑ_�<��IDkH�R��A�D��y���C@�<���?c�T1�C,��h��PCz�<q2A�cԜrOI?"th�w�<)��Dzö�`�Q�L�0����z�<94��*�ޘbb ��w��'�\�<)��#a���b\7�,�`dƂV�<�!��^�dճ��P��|D`�.U�<ɠ�}a|,��S2h|̍�6.�R�<��	��Xr=��I%Y�nhh�C�s�<I��	A�c�釞 �Xh � �l�<���|�%p�Z	묵���f�<qd��0�3 C�`����'��_�<� �Bé�XɲaY��
H}�"O��F�eu:Ļ�ʛ:Ҩ�b"OR����Vb��"׎U���L��"O�<������Cc�r�`��4"O�س�o�7!���ed}��Sj�D�<��9��qd�h'���U�<)DG�'x���g/׿yL�<#���U�<1��FGl$�`%k޺�f�!c!�e�<a�%��B������gp�[Ջ�V�<��o�C�F�+�aܳT���sɔ\�<�$��%xp2���O|�y�k�Z�<�H��Lʌ]��燩c^���E&�Z�<ID�e�HD2W���~<�{4�m�<cK��ZI2԰��ߞ~
���u�L_�<A6�H'���hdiX�I"V�؃+�u�<�Q*۬=i�F�s�����!x��h� �Wզ̓����(�6��e�G.2���B:D�Py1$�HÈ%�2-X�� p�@*9�j���a(ʧ>�����LS���Bf��8��)�ȓ#y���HB�1��I�.~�"��]$�gi:�)�-�\�b�Nicڜ�3[)F]8�ȓ��K� �9
��RZ�T��'���.
T��4�A�P����s��%n�$�b!OB�Gީ얹k�DܻeM8�C�O��3׆`;�b�<fθd��XG{t�:we�S���$��ox,ѻ�kU-.��xa���e��Ɋ�bP��`A-,K�$P��:�p�O�	{2��q�K(�=��%Z	N�!�d�&Mx����-^����,N��vi���׉o�>���|J?U��I�
���]���}B�,��u�>� ���P�B�I�V0��X��Ј<R�x҇�-���3��8?�����d�cNKY�\�o1�X�5(`����PȰdM2����I!cƸ5�@�R�e�9�al;L4�2�7
H�@tB�>7�R�IP�s��q��, ��|RHE�!�`#a"� e���HT�<���T�AJXX��-9����0������t#�� �P�~��EQ�6���X�'�1(1��!60v@[e I�a��ۆh�ZaoD�S�dY�!s�ٚw�zXi�2��i���G�
��
�'uzYkv�B=&\k��р�|Ej`'����dۓaۖ����^]U��Ȕ��(O�,���i����$��(G��1��'��M1�YF8`�Ĕ�F�x�<�L��#*Z�e;�t���U4a��W�{"���79+z`3�hЦ>�u�-B��Z��|)�NK��δ� k]?&���S���}�&��l�$�����]L~C�	�r��-!H!_3��0U�MS��)#��"2A��3��?�2Q�]/���2e��0c��}��C��ݍe�HB�	%� N 5�&ez2=y���e3?��h2����ۆ"�����&ʓu �LڴO�9[�D@d�\4*}"��Ɇ=�����-�M��+
��pM*FC3;�B!��탿8rr K��b�41�W#^>��dN�E͢�+��`�V�2%�^�X��I�@��'��-i�EQ�dBН1�)P&��I�gT=[:pK}!�&X�֥լ�B���+g���<(p���b��l&^A:W3J,��<�O5HK�d��+��8a�M�c��@
��\�j��lN���2�.��o��%�JR�R;��U3j���J>E�ܴB���M&٦$c�!�&A��D~�.�1��b�Z.uaG�*�B���b�L}r�:�<Q[�'kz)&�9w������=Y���y�Oȸ��D������N�Z�X�mt�i�6.�#-�P�!%��&����ȓx�ܒ7��l>��S��G�r9��9�0H��;Ozu����鞧r6F��<��[���SD��,�4б��	B��)�w�8	����_�,���.��"�Mx'OΤ*�J�����I?��`�9�&T�i>}rKJqܓ`R�� .z��[�0[��EG~�OX@)(q���l�� ���N� қ6}]YS%B�o��X�u
U�#ϰLBC�i*�A
�Ŏ1+0N���N�!�.P�d�B�V��� '�N�E���괐�!��<*f��0*�(��l?��'�XU�'h�0(��a uD����I��"OV��pG@�	:p�jvKS|*��k�n�H����N?Q�'h��OMnhȆG79��杷���2!��D�z� A��>���DS3/���p�C�N�)B���1m��T��g�j?q�'G� �W�ο=�"]┮�3
а��{
� &l�&�OC<�5���&#j ���	)���5�	0N`T4U���7��;l���J�:�^��σ%'s:��� �N*�q���p=���%8Z�����2N1��o�A}�*�%6���u�Q�|C�����~"�O���%%��E��XR)ν�F�ص@����g�$�S�9��У"M�fV��m��0��U0��F�<y��'N|�?ѡ&EcӬes�w�Y���7G�� �sk�(,DD83�'DX��Jο)�`�Sˏx����U�B/�����O�I���ͭ�.����?a�W�R0]F͸@�gi�(�a�� ax2b�%J�9I'LI�H��!�O��@��|w�dr(��1�(u�d�@d���sO\�a�{���+]�2�*W��,iȼJ������R �{�쉥E��x�KeqO�dCC�X�l�0��\e>P���Y�<�s�׻5^� j���9�����	7~�Y�-�fO|q�=�O��P�aዳ�y��H�^֌*����x�ܥ��� ��x��X��6U!�L�$l������C��\�I�+��ۋG�ܻ6kʆj������=���k0V����&	�&Q�AF�;u�����ĭ7x4HJ0�
,r�ި!QL�X���� �V�4�*ʷDE�����y� �kABC�|!�����1C�u@C	�#y�FL�Ԭ��j)�	�rz��"�O�X7I'��IB�f������ERye��E� Ly3�J�^xL,��^ (���ԂO��M���յ$ ~��yqH,�`�nӺ���ԯ9<@Q�O?�S26I�-	����ǈ�n.�u"�'�u�<р#ͳW�԰��жg���蠄�[~bk��-O~ԇ�ɍ>Y@,���C8f���G�6�����ݔr��7M�@�e�5j�
aq�╆^S!��"xO�` SmG�=ؔ���W1 !�d� ��X7�WU�@$ޥT�!�DA/�~͙PCW29�����%A�!���m4� ���6=�EpGć !�d��5!Ճ9���� 鞷'�!�۫5�Xe�FǊ��p���M�!��݉g\�0gN^7}�" 
�i�l�!�@6�`�C�bED�L�ӥ��)r�!��.Q#�� &���c�����H��~e!��T-�P<�s�G6K�|���,�2m�!�$�?��k�喹0� ���2�!�Hj�( ����ju����	:�!�[KX	��"�F�^��@�P1.~!��Q�;1�< ��1
�]q#�z!�X/q<����ͬI0~�s"��ks!�Þ*pN`:V��7)+:p9kK�\b!�	Z+L�HB(�f 1��A_%!�䍃1��m��я0�,3a�x!�Y�����L7��j����)
!�dD48u ���$k�pB.�!�$4ֺH)��#v0Tr2����!��APU�t)Ȃ.��(�;r!�Kq�� rM�'vĐe{�Z6K�!�d�35?������X��]aU�٬->!��_=&~�PESfE�)G@܄(#!�Ā�Ua��i�݄<! � !�$�7x.5��G��2	��蚇4�!�dە�z�
����*Ĳ�	��Mg�!�JR��Qu!\�	tY�EMӍ5�!�$\�K��h!�"ٷҐ-Ʌ�U�U�!򄔄ϸ�)��\?!���o�v�!��4 R���Q�p�~qQ�ʚ\�!�dR�[,ԕ�gj�~�4�いB!�$�(P��LrA� �pz`�׾"!�d�-\w�L�cE�4����	d!�D%O"LK�K�0�ƭ�� K>h�!�D��� ��ˤ)lr AD�m�!�G�AT�d�6��A���H�$��j�!�$"q�=��d\-�%����!�d"u ���F#P*Y�Q�_>K !��I��13���	4E I�W'� C�!�� ��r�ƚ}X��(�c��;\N��"O4�p��(-���w�O�ID��u"O8iQ!-�+F#@�㶁=2��J�"O`0@JP)D�}S��V�9��h�3"O𹊒�4^ �;��*#�f4�q"O<P�͍�K�,A��P�;d�qW"O���&��('�\W-��Smrj�"OTA1� ?M��aW͊�:��\`w"O��@B�=�
�yg R��aK�"OFP�M\�+�<�f��3L��!�T"O����%U!u��j���Ce*�@�"O�����9`w�C���U���"O\e���*�d�pt,K7�p2�"O���8@q����j�9�z�Ip"OVY8W�M�mJ
qb&�k�Vx�'"O���dϐy�!
� ��0��p�"O�ȃ��F�+�z@����u*�I��"O�A���(�9B�	B�^��|!�"ORU�vA����p �'H�,P3"O��P�F��!pF�o$r<3�"O�@i�(I�-n��A�d/G	��Q"O�,ʑ'*
�:�y�#L�X�tٸ�"OH����Ju��l8s��9��pP�"O�u�J܇`����*Ko�R�"OʽR��& G&���C���Ȩ�"O���A�Ų0�b�b�	�%�3�"O�<s� �8u���E̔;q���V"Op��5&�:��u�����V[X!�"O�����B�'	>�[dA��TYB�(�"O�A�j�+b\��z��4?n�!"O�,ѣ.L�>#t}I%L�_"��"O<=�7 Z,Z-d���J56`u�e"O���i ?2x�Rw�#z�E"O4�4
H0N`�Q�_�4�DD��"O) �
��J-�:"�.YC�"O�H9���� �4,L+!@J���"O��S����p�1���
?�a"O��N� ^2���Q��0;>d*"OL퓖�3K��W'	L8 H*S"O�u�.|��BȚ4G|r�P6"O�PTeϦcb��W&ܳ_Ϛ�!"O4��-��y{��L�����"O�W�ôtRP���-b���1�"O �Z�`��U��$#��_p�Dɠ"OH{��ły�L a!׎/T��3�"O���r@��Y���6o�MpJ�Q"ODcS�U����Pb�Vq||�{"O�����u��E�7jP<Yp���@"Oz� BX�f� ��@'�UWB��'"O���Q �IGԕ��gEcTp=��"Ov�I���?}2�t�цŭK�1�"O�c�A =V�𘻣��;9Ęg"Oj�qĄ�|��ag�#{�~�H!"O�	�U��^��"�/�%x6"O�z�gۍI���s��W3$�@��@"O����Y�[T�[e��
o�̵�"O֕����LW���[,j�"Op�6ؙ�I�[n��  X�;�!�$�"w$�(#1N�80��b�B<�!��46�-���έU�D)V�ǵP�!��؍vn�1�HBU"ES��H�U�!��9_6�lz���xH:�2'I~�!�˿P��J�眏W5�%R�
��PyB/ݘg�.aq��ʬd����'D��y
� �	`���7_�	�A+��G�h�!"OD|�
��F�6�G#U��,Q�"O*�20�({�t�ddC�]@t"O�T�.�> <���Xj��C"O~�KA"
 �r6���2�M`D"O�ͨ��^
G� ԓ�B� _��`�"OY�6k�$�uk�@Hp{8�ˡ"O��P�٫i��+���]����"O2aH�H��!n|�����=
�$I$"O�|9����촳� �, �)2�"O�}	�\�6���e ]�D��PT"O�Ъ��]��]�w�W�� 7"O^ѧeߞ��+"cL�bH��!"O�� �Ȅve(��'�°/���(�"O�5"�E��j�2��ց��W[���"O�)�g�J��ݰ憁�TSJ��W"O�Pf�2�P8�L�rJ&�"O�0�a!j ��#C�)Ռ�i"O�Y���<RƨJk�-vʌ@�E"OD!��!؁�,@d�U�޽H�"O����d[%k@ay��F&��a�"O̤��BN&ǂ#��x�D=H4"O�����0��i2� ��NЛ�"O��.!���6��W�����"OPe�ШӼD�țsD�?X�H�1�"O�Ӥ,�>�h�@B�܇�~�E"O� �����V�Bv�R�p:�(R"O�t S�Q�uGIKqnU�4/���"O0�A�+�|�XU�Ά/pZ"O ��Fi�3�̳ �	$n�$y4"O����G�"'18�V+�[t�k""O���K��m�v�-�܈�"Ox� ͉!K�:�J��-2�|=��"OZ�ř;�"�c	@�$%�"O�s��Z uE���3Ȑ6[�š"O]ZFF_�x�2��S`�F��l��"O�ѐ�+[�D�)�17�إa3"Oұ�%"Ѝ �6�cd�f�ԕ�r�	z�OBѫ1+coT(BF^�8)B���'�lE	
ij�Y1O̯]�6���'��1ҨFTʖ����[���+�'��U�F�V�D�9	�U����'���:�[�6Ɠ/�Pq��'���B�a���9n_�)��'�Z��ǂ7�D�B ͈�G"�h�)��<��C4R�ʔ�M��$����I�g�<�,B%M� `�#�-��yE��c�<�t!�� �\��a�ؑ ,����z�<)'+�@���Ve�0%�l�3*�}�<9Ҫ1w䆤cd.��*�����Is�<�4�O&oTI�q�T��Ļ��o�<v�B�E���!S�\�jpF�ӑ�l�<q
����.B�$9v�
f�<���"lMҹcD��>o�Z$Y�i�e?�����h�d�$�[�
����5���8�"O
l� b�AY�U�����J�<Uz#"O�@at(�g ���݇X�8ѣ"O,t���80�,z2�'5�H��"Ov��c1ix�[���f�ظ�R"O�E Ԍ�%�BL���_�Z� �
�"O�-X��`��U�wᅠw�0�"Oԑ�ՆV p}8z�o�0�ʬ��"Oz��ַ:̝ZS�(��[t"O��s4Ǐe<-��F1���pG"O� \٫��� 1_(�����*լ Zv"O^q�4!�(�����ϩ�X�(E"Oz��+�(��!��hL����0"O��(#�\� Q�D�nԄ"�TC�"O:�h�U-c�t�s���g���D"O�݋�.�<p�� ��!|=9�V�t�`�'[fU�����r����d��&w�l��
�'|�Lj�	�XRP��t�C�g$�5x�'�(QR�U=#Ffձ�.Y2dZD�`�'_ti8B�M�OZ<�1�$K)(V���'%��#��I��i:�kA��VA�']@�	�F_�xp��xA�W� �!
��(Ot�E��-!���S���a>J$"O��@���5#���R���I��"v"O�%�фT4L^�͊���*R���"O0	aA����4b��%�q"O&��BCȈLϮ��eW�&�Z��"O���W���M�Y�3�R��2A��"O�:U�E�e�D㠢�4]1����"O�h��5q��0y�����8'"OE0�,�_�x]A�ˊ�(~����"O	���$O]�3������""O2I`�%�*FΌ1�C�(,��X �"O>���Fܫt>D��I8/D�]a�"O����,T��`��ٌR<�	zT"O��g�Y�@Yqu�	/���P"O4t����=sN�:���(f��"O���v�	�x�Fh���ΰ���"O����� "^���9P�V�=T��ɴ"OZقC�A.�80�甀qe�p@�"OVu�DD�TT,ӠfHU�g"O�����%F�Vгg�~��l�%"O�x��oS�4����悺{`��h"O�X!$&��UW�D��F�0!�0�b"O,HUH�K8��p�+P��\���"O�A�P�N;���)���>S�}�"O ͙fψ
P+�{�O1�R�Q�"O� ��a�1������R�\����%"OZt�"��T�X�J�<�:@k�"O�H#MY�#�lQ�N�,^��"OP� ���&�v�X���*d�۰"OrI�ŋ(�� �-8�~���"OF�YQǚ;*>]!`'Qe����"O�5s�aO���H# ��=hbv���"O�qAw/B��}ū�3V̰��"O���6,��"vҍJ+�zdTa��"O��HU�([�lc0�Ĵ[[P�U"O���B+Ɗi#X���8V��e)@"OTY�䩇�&I��Q�]�B6e@"O@L �莩J�
hX�2]v���"Oti��bB.ĢP�Q�M����"O8���);�x�Ck�#|��);�"OtȠt�jh|e��d�`6�c"O �h1�D)����ļRM*D�0��%� w#|y[���V2�Y��%.D�x��!
�ׄ(I���q��)2,?D����ޓl��1��
X]ܪ!@e/>D�л�J\�Oe<��r ل=�z�	C�0D�xb�I�*-$�"��ة6b�q6�+D�d+w�V�e��cuBѵJ���5�-D�`0s�g4�HA���~�a �,D����� E����`H4\f��� �+D�p��g_4E���y��E1*.�K�$D����ɗ�SN0��C,A0�@�,D�� �l���B�Z�¤Hr�ҁzH�0�"O�i�1�$n�pX�H[�+�\%��"O|���Ē7r)>h�C�ɏ&�5�@"OJ8x���T���˗�v��q�"O�����
�8|bA���T4"O�Ԛ%ץ~kT�3�$R��Ũf"O�A�bǔ�@��qjZ[�T�:"O��Ð&I7)b����4'����y���h���5j�M�@��J�	�y]��q��[8�T�
 AN��y���)x�v杗 m��g-�y�D̶v���rՌ9�yСE���y2�E�~`�U��<~:2$;�nJ�yr��5.������J�}x�I頊�$�y�
�g�p,+�b@u�2�
S�B1�yb�)S�~P頇��nZ������y�J��]��0��P�O����F��y���R�tI벼dy����3��ȓz��h(��/<y0@b1-��l��,� ���0��4J��8�VQ��TruX�1ttD���BB�	�X��	+��E�ސB���M!�)-���qi�s��zt�¸N_!��l	4��c��;*O|�ɰ��(�!�
!f!�����T&bh�W�H-i�!�DO)4�p42�fR!d98��ԎǗa!�$K�'��:�+ �0=�h��]��!���*-^�h��~��8p��8�!��<3�R�r4&   bF�¯�!��Y�L�aU�q�u�W�U�!�dHiE;�[�h��1�kӿ/�!��xn|�#���g�Lr��W�e�!��N�P�͐*���$т7fµ%!�$�^p�e�]�3m*�&�I�b!���d�ra��E�,m�8VٰVb!�� ��Ä@_�Hd2� ��Z�wX!�D %D/�� 蝬&Z|eۅ变1�!�јQ�=`sL�
��@��mE-1�!�D
�u��r�O>DbN��PG�<�!��;����	�Mu�D:4'��y�!�ćnҨ0	�-B�6�h�@fI�H�!�$�>��uY�KV�~%��[�NW�!�䎳)�8�AI��x�,0�C�1�!��?LV�q�R��D��O���!�$%h�~|��
@�.�lJS��'�!�Q��mI�P m�`�R9�!���j�����g�,q� 	�\�Pw!��z��9�'#�|Z��:�^h!��m3��:�\f�\�*�& �!�d��,ݦY���բN�H�GH˸V�!�T�<����Ǎ�"�!	pGµU�!�D�'K�@� � �����!؁2�!�$������U�H���F9,�!�D�4>U��8Ed��� ) E���!�a�t�wO��)㑀a�!�ޭ�tuj�-қL��[�bFV�!� c�����J�C˨UhV��0C�!�DY�s�f�3SFT�B�bX����a}!��K1��KmË@G�%� ��o�!�C�d+��y���& �X̒��I�!�D� aݞ�k���6�,E�t!�D,�t���EA3���e�ן.N!��	&WwzL����Y�`5I� mM!�9�B���VacP�+p��_�!�� ��b)��;�>�C�%wu�:Q"O.�Y#�C��8�!�*tNX*�"OF䢀m�':i���n�<jB�șq"O:IC��� ��]�a�D�})vR"OV![#ٺ�t��i�`��"Ot�i����*P�d���,^�Ģ�"O 8�Ċ�'J�z��*½Q#��+�"O@�Z3�
3�"	HUl�# �F)*�"O`�)�V&H�X9J�m�$�BP2%"OԻ2	�*�6���ҎG�~�cR"OHp�DM�p�F;d�R�7����"O$}��B3�u*}��d�1"O������A��q��枷 ��sq"Opx0��� ����Ae�3aNR���"O�d��d\Bg��Æ�X�"I2�r!"O65�p��zy���#�!H4��%"O����χQP<���#43\���"Ora�oD*{���*1�� hI�"O�@�c\`���j����AZ"OjԲӯ�n�$��"�B��	Z�"Om�#�H�ީӱ'�-J��"O:���e�=-�$���B<�&�k�"O2ȋ�/ʇ{G�H�7�ޭ
�d�9"O���E@י�X��GI�1M�L��"O`t��g�;$��w�"{�B�a`"O���n�� �,���E��=b�"O8d�W��Y���A�N0d����"O�-3�E�u\N����B�$;`!�$P�=J$�g.1%z��`��Z!!�t�&�` �s�^�0�(�5f�!��I�=������m������h�!��@{D��6�U4��2�="�!�$��1����b�@��;�fÏ2�!�$��FYvt�����A��0�!�d�:�@ͱ�g͓{����D�/y�!�$��Dúy&�=L�|�WL�v�!�EG~D�����7T�	f����!�$�m.�P����"6��M=!�D��0R
 i���3�����,$(!���f�F܋w��Oxv�J���#!�D@3^��u��ʖX󮙷D!�׾x�&%�Q�<t*��Q!��
�|��u)UFB�(5@c2BՖ`G!�/xxPMkbNM�$~�����xL!�Y4')�+4��l�B4I��O<{H!�ĝ�Uي S3�$�̘y�#R@!��3�����IP�E(!���/�!�$�)*�����Z�-vB<�ЏF4�!�dJ�=W$�Ԫ['xz�Sr��`!�M�0�b� ��S8t_ȹ;CN9I�!��l�(,1թ5^(T`B0�TX�!�D�O�\��g]�D
����B���}��ܦ(����
^$l�C�I�N��<f���;��ΘT�B�I�D0X�W,�m�fJ��=kV�B�	�5����Շ}�`Y�T�[�jB�I�n2�A��%
�y�� �1?Q,B�	�8_�Xhe�\ 3uRM��ۡ?��C�I�iȎ�y�I�
1�|y7eN�8N�C�	(/�P�¬��Q0eR�)�lB�Id=�e�ީ"Ĩ�"�ک)�B�I�8��+���o��1c�$X�W�B�ɸ-)t�s�6bx��� LYB䉪I9<Lk��L}l�aIn{�C�)� D��̞�7^��6#J,�ɋ5"O���N2����,0�"O�e�7i�Z[,��e'Z�t�8l� "Or$q�Bzr$2��G�_� �c"O<}���*6��]��Ï/����"O4��B��yK�U�&@�,I�lX"O*��Q�=@\a���>�|� "Oh8K!)���nyq��΋kO�!+�"O��0�hߞW�fp+�$WO;�-�F"Ol]���/.E���C�e#�%H"O|�U"
8ab����lK$���yB��c} �Zg�D�aU�ũ`���yr�ʦr;��YĈ	w"5S0�_��y԰NG�l�W�E ��X�bP��yrc7(��L�֭��s'��CFm�y�̓6`�-�ˆ�a���+6-��y"�ԗN��kB�q�4���_�y�f�Jh[u`Q�T�b=�d�K�y�	�W8�0��ޠQ��KD �'�y��D�A�x�2���7��ykCl-�y���r����E82O�E8�oP�yr.��B�Q!~<��y���~y8�'�<P�����`�x!�/�tg�E3�'Հ�j����oAb)K�͛�6�<a��'�D���Ų;V�)؀HH�(���'����;h(��!Cj��JR�U��'*�X�r\h�� ��ҚEi�8��'� |� h�	���;'�Б6v����'����#��]H��hQh�4zx�C�'brDs���9Q��+qo��A�1��U�L,k��ͫp�
> �G�=D�*����r��1�
w��)3�!)D����!_���X=-#��6�&D���Ĭ@��]��LUײ�*3D D�D�[+;�P{4�M�N�ɣ�<D���C�7~%�=��f�)n|I�p�>D��+a�G��=ۂK�{ҦȨǆ'D��0Q
XZ��&���?Q|�a&:D�l@��
ze"�A��v�l��4D��c��A'F=0c͘+ђ��FM(D�H0�L�,�Iړ
؄#�`U� 1D��a0��0�Acs��p$�H�0D�����EN��f��t��ͱU/-D����Cɇj�����C���	I��,D�(
�Ey�^c3�����LIg�(D���d�~"L��Uk���||pO+D��e��a#p0�׊?�J��W�5D�X�	��׏�wNa�3.D�).M6�,���摬!ƊP	f�+D��ۣ�c��蛠
%7]��'�6D���с�1X�H�ȓ�D��5��9D�2R�'����D��=O^`�CJ"D� r��Ɔ8\��L]joV���  D���$C�L1P���[J��q�3D�4�Q�C�g ���� �$�J�1D���� �K�$��mͰ�T�s�.D��!��$_*�Q&�L�8�R��6D�`�o�&73�+�zȆ	2��5D���5�	4^�m��"Ť[�@,�@.D�`����<,�6�2�'վ�8�#/8D� 9v�V%V��a��k�Z6��B�5D��X!@Y�a�0�a�D�2̵�F!D�<���Ա� i
w-3G.�f�
B�I;8 �q�F�S�5��,ΫY��C�)� ��;!G<o� ����U"�J�"O�A����}�ŏ�8o=����"OXf���Z�6i`�mWZ�`"O�X17c�3�����5Y����"OpP���WXn�x�&D�����"O	�	�
�ƭ�1Oț���"O~0�	X4cM0��ë!}T0�6"O�9��+�fV�E����]����'"O֩��[d��\Y�I���V"O�5�R,�� _������b|3R"O��Q�b_%���"��|�d0y "O�� �I.9���RUG)pT1�'N�ٓ-�l2��RS( �д��'� ����6�0qK#(�~<Y�	�'켭Q +��YtF��B�@<r�`���'�lu"rc��{��a2.́U�X(�'w�pqu��&>̺-[��/
�ԅ��'<��1��'�&����ϻb��'
�ݐ�GL|���h#��%H\�x�'$��3w�ւ\�R�Q��B�S����'�X�b��4����X�w�<��ʓ��HP@�A&l4�h3���n�����@���!ez$-[��V�2.��ȓK�z<�0+�8Yq�X2�5M���1�(jv��e���իF(!�&4��RI,|�el!I:�i����Hk�G?D����#V�B3~x��.E+s�� <D�H#AY:[���� ��%S�0D��o,c�(����*�ޔ�0.D����P; :�g/�5;�e�E+D��84�S�=xu��.PM�Pa(D��	�"�<<���р� s�&D�����̳I���Y��T�\���4h"D�@�,��j�L���Ԭ`؎���+D�@�&S�
l"�� �S$F���,D�|@5�-0��C�������+D��I��E�#ቜ�hM�+D���g�?
���k��[�"E�+3�5D�T`�ʛ�nfti���(9:4(D�t�`���u�\�����5�`�!&0D�<��cUL̽��Y1�~( i,D�4�M�i?.@��N��s@�P��)D�艶f&Ye�q)Sp�6d��D'D�t�p�'"^���@����T�#D�$h'��7�(�
 T���ka�.D��J�/}yr�`� Ϗ~�Rt�Ѥ,D����,I�^)੡Ql-<�R��N*D���]�	K�|b��!x��L�F*O����"F19� ֢PF���""O���QkW�wwl���d�9+|1�"O�ɺ���pNzM� .\�s8}h�"O\�2@�A@z`���@8 �4 2"O"�X���J왓pn;���W"O�ط���:�����W&���"O�0����0r� +'�F�00��P"O*�)��D�c�>����	8X�T�a"OʔI��Q7�v�X2ˉ? ��"OZDr�ay�I���,<đ"O�\bf��nH��H،TF�4�%"O�H����)SKD�(
P�#6�P[�"O��R���+�\��5
� ,� 3"O~�cF�W�c x�y@)M#S `�q�"OfdHw��!;�5����P����p"OΈ �NޫN���+�@�;�h���"O� ��
�F�-Z����<�:{w"OD�d�5�����7!��Xj�"Ozx��Q�{�-i��ݛ�h�"OBT���m-�舶��q~�;�"Ob��됧k�^ի������$"O�q��'�=��i���r�l1�"OB�1�S�R� ��/b`��"O����N_�9'�xyt��eP�*�"OLu#M��&H:�`��T�Z�HD"O�M��hզ@���7.F�a"O�!H����B��Aqç�8�Z���"O�kP Z
+#������%�>���"Oh���
i,� ��k[�x�
�d"Ox��Po�=p&�P蔦n��u�"O"�)CO.F�1 ΃:?`�4"O��B#=G����I.
�p"O����ʝ�E�dДs�1Q�"Obڱ	�.d����ܼ;
�}��"O��z��Ҥ6�z]���6u�
E��"Ot1@��˕*�ؠpS'�&'���٧"O�l��C�#������!C""OJ�[s;�� ���P�b9�R"OH�b/��E�8|���4"O�M��Kd�^�vkX�{`xi �"O`�(����I]`��g�x�
A"O���!b� 3"�bF��)N{���u"O�|˖&�2 =����`P����"OPd�!X�{L,h��oD���-��"O��� G�d�w�Y�m�b�С"O^��QgH1���ǚբ2s"O԰x��A/��@�F%X�`F"O�9��>;��)��^E΍#�"Ođ�!oN3�(1ge�"f:<8�"O�@��ۚG��H��݀J%�l0#"O! �霏ؚEȂ��
�� �u"O���q/��'*؈�� "�>X1R"O�E�T)� l��Y�i�7"nI
A"O��r�Q�vyI�G\	"��a��"O>���$��1%O�G����"OVd�"pE�$y�$�0��*�"On:���}��� ��p�"O��#� 1S/B��M����"O���L�>R��Cp+_/El];�"OE� -��/ʰIY1��j>�D��"ON���D�"X�gF# |S�"Oh!	�.�+g���Տ�"?�d�"OtIrB%��T�	�P�]����"O� ��?l���M�:�4�1"O��IC÷&�6L1&P7*�"�x#"O\J�M8#d���n��)H�"OС� �W(;I�q"��m^��2"O(L����N���A�,<��`�"O��
D �5�`�
ƻx�|��"O�U��C$1ƴȐ��ԉL����"O�d8^ɶXceǅv!F�1�"O@MA�N���E�%-�*q�:���"OzEr1�B�����k�6�J@t"O\�a�oN2M�p�I�(�*-V�s`"OLATh��9� �p手USq��"O��r&$Q�Z^���O�*����"OXH�B�G.H8"t�U��	J�"O�e�`��'p�Ҍ^�]�d�:�y���
�^�i��Ό��&�Z0�y���]�` k�-3|L�!Eጰ�y
� ���*T_�. �%ڐ'����"O�$���x)p�&d!$� z�"O���+�w�����Z3C�:'"O�T�f���}�8P��X�F|�"O�)	�4t���$�14m��*�"O��J׀O.�m3�m ZVLiy�"O��dA�2��(`p.ٌLGL��#"O�kg��^܍�0(�7H�J�س"OU�&�=2�f��?(c�R"O�=Z��N7Eq� [��Pc�@Ș�"O��r�*֑REכ��@�"OnY����v���R�Ƀ-%Tx���"O��x��܋ U|:5���`;v���"OZ�#�P���C�B,`��W"O�Ip��зnl�1��8v�Bt"Oq���� @k�c��O-m��� w"O��Ab-=&r�D��dI�E�e �"Oae��T��r��S� ��5"OHláBT:T
4���A�])�d"OL�0��ٜ�1Q�H<P�>�"O~&ɎS���PD�0H��p"O���t�[�$�C�!7qh,h�"O�8 !�ȿd�<,ҡ���/va�"O̔�1���Ԑ�G�'*_ ��5"OHuC��U�xFL=a��(Hp �"O.�	�.�������% .9؊�"O\�2��ۿ\4[ʏ�a��dA"Ox��L|)�	��g�|qz@��"O��2��2:��gQpx�'"O���0
��1��զB��Ur�"OVL��K��5Dڸ�b<#����0"O��!@72�W!_�x��e��"O�[��µ/46ÅT,xC!�<t!D�
��\�;���R�R!�d�?&=�xg�
�j��j��Q�F:!�D3J@�Z`���HC�����(!�ǟbW�E:���:8=�E��3|�!��o��c��]<.5D1��m�Z��$���ѣ���ZFI���y2ݵ7�&�J���A�%hC8�y�#ţ1�P�p�ɗ:���4D[��yM�����5��!/M��$FO�yrF�X� �R$��4��6�yr��x��!bS`��E�pA�#���y�]�YY���Ӎ�)=�:�3���yN�<n<.!&�+�Vm�3���yAч� ,a�*�8��y�b�Y=�y�-d/4c3H]�^�tXYB��
�y���z�������>]�8("Y��y�d@5l��2�6&9#B ȳ�y��̲:�L��ʊLi��C�:�yriʵQ��GNBlƨ�@�H��y��S"Z���ԃ;	J���@Z��yb�_�]1|P"��	�����	 �y�A�:\��_4�J��mT�yҏ�:nJ��b��e���J���y����X�z	94��%l��{e���y���L���X&�(Oda�'f�y�@U-�eɑh��E $��9�y2
�Z���0�-X�E����y2JM�D�9����u�@=ҥMҩ�y���m��X�S��j訽r����y­U�f�� N�f��X�T%��yR��KƐ��=)Ťɲ�W��y
� \2��ջ@��Y�ā�iF�*�"O���eԯSA��r��܅F`�̓"O�|
���;DO�1"����$OF|;�"O4<�eE[�e^���>4n�	3"On��t���j%>�2�	V��%�"O�)�sa�xX�����\���kv"O�dpBG�n���#�!sa�"O8�'��%}V��!���2`��Ѡ�"OpY�$���tM�Q&���B}13"O6(��T�y�l�[wn��zAư��"Oz�bЂ k���`��Z5rA�P�"O��k��׊lpZe懼lY��i�"O��1Ҏ�(C�yQ���'?�[g"O.%�wD�a�p��S�.:.z@�"ON|Ȥkb��{т�#B�a"O�ό
k�J�r���j��U"O�5��t����Ã^8q�"O(�"���)M�,��W?A���"O���wB��?�l�ˑ�:A�%{0"OP|『�oW�@_�R��"O����NS�K �I�C�Hlj��"OڤyR!O�6��'�, k�%�"O���H��j*��U��"O(���"O8�,mr�(.�8T�����%�y��7)�XJ�����Ba�F	G��y�J&(_,A��ŋZ����%����yB��Z�4���N�K�1 �6�y�nӗ!J8��m�3DQL-�W��y�*R�I����$�'�iÛ��y"����Z�(W:�%�1�I��yʡ`�����r�;a��y"�ۉzT����@�C�*�']��yB҆e8 ��旳$�!5�y��2|�(QcM�1�Lq��0�y2�)Sp�kR�</X\Q�'X�y���l�"D	q�7'Ί�:�"���y��Q�5$_�rg�xr��܇�y���nH�FF\(o���C����y��A 򢜚�Od��P�3��y2*ܧ
]��D�W�Z?�5�����yb@�������X�VB5�Y5�yr�<�q���g�p�cM���y��IU~��;`gY�a=t)�c���yrO�,m��ɓrg�"y�1'L���y@��h�_�1� A��N4�y2� �2��x��JI%)�̠u.�7�y�T��)���A�3{�}�$���yB%�z6��K��5���9�J��y�G�$��
_�`u���sNR
�yB�^+;�-Rt�0/�\�Ӓ�k��'Y���T,�_�T4�b�W:+ ��{	�'8��c�R���Q��(�����''�`���-c�j���C> G���'a�jp���f�x�<B6��1�'3H�8 Kƫp�|�G,�9�<S�'��MI�E����\k�H*�J$��'Hj���L��q	0�Q��)��y)�'�YB$قZ�pi'��D��'��I�E-߶?�-;&�& vT#�'Af���$�
{'�]╠Q	 �� �'z~}�6̛�&+Ϗs��	��Έ^�<�F�U�V��-�DG��jj �z�*	s�<�7�'Z�HqpI�"r���C�A�U�<Y�N�U"L�"A�	*��01�EH�<� "-#jKT("��o1
�av"OΝ�=7F~p2�T#��K�"O�����܁d��|��ƈU(C"O�lɱE�/6�.�#ԇ3e"%�"O����,,�*�����;���8�"O^�C��8 A��� �*t"O�8�q�Y�I!���!	Y�p� �r�"O�tȁ*S�q~���h��\.J�F"O$ �  ��`6vY���*�DIP"O����M�L%�J�=X<��"OԐ���J-W/h`q�"ȝ����"O� �ƀ��N�X��� M6'��� �"O>���� ��E�`��	(Rf"O4@�����Zt�
�Zը�Z "O ���D1��j7gCE,45�0"Ovݑ�C�]0��ehԙH�9��"OdtcՄ��J�±1pF;P-$E�"O�Lڠ��0����$l��"O�0�R,D�U`|��7��g��=�"O�E �O�*!����G_;y�9�"O8<x��ޤpaU`̉U�I�V"O��T-� X�ɋp!��n��"O��S4��Tr�ţE�n=�|�"O0�k��6�`��0̾mܞ\R�"O�t�4o]6�\qfŷNش��"O�D�oJ��8�B�Τ��"O��mcѸu���I��~���,_c�<��A�?G�j	��)WWh�:5�Xg�<!�˳B���i@ҕ2 ��c�<!�I�;Tz`���O u{��y3�G_�<��iC�Ͼ=�&E��!YG�^�<!b	27o�U�@������s�@^�<��+�v����`��v�HNe�<���]��\h��L�x�[W��G�<qVj��B���˒*�!b>L�Ŋ�\�<1�
]��,��S�4@6���,�m�<i��I1N�D�"���n\h��S�<	&��Lޞ�c�xx���z�<�h̵'[Q���I��F���Lb�<�	�J���\�BU(�
A�V�<��%OC�����U2��7d�F�<A�+k�H9T�m�UP��D�<qª�;k�8�����Ft6X��D�<i���F��6`�$
`��_A�<�S��_-�=*�o�'�\yp��t�<1f���A�{� �/?�0H�� Kq�<A"�YwL�I��̮g,�P��fIV�<�UB�?q��yɰ��2	��&�Zi�<�#Iw
X��W�=�:��r��f�<.��z�H�[0֦El��vL�a�<Q��ڤ.��P����7&J��W��Y�<!TJL�e� ��c�X�9�L�G�W�<�g��TÄ�
���D�K�<!G��aY<�)�,рeS�Ͱ��M�<Q���<k�L�k�H��l�
��AL�<1�V:�.O�:WT͓3�J�<Q�&�*� "�L��>�d�Q��E�<I�Yuv��k�&<�&S��EG�<���������ƺE�(��"��M�<9 G%~���aƐnΪ��d��M�<q��ɍ=���knAnݰ�H�<R���={|ppń�rZ��x,�B�<1��I�L<p4|
ؕ@��A�<�d�$f��c��_�<)p�f�<� 2�RD �I���C�^�Ԅ��"O�y1%����E юԋa�n��"O��`Q��4�!���	/�	9F"OV��f�� ��i���:Q H�e"O�)!���+|VɛRg
�=	���"OP!3BF�&B�@1f�;���Bb"O (�Ʉx	ö���n�J�x"O�(p�A�H��q�N�ry�q"O\���%��#`)�!�ؐ�"O2���+ �uY�ؘ�0���"OR�UG&w�$��$?�8d��"O�D����q=
�N��pSP�"O�0���~4��Ƀ��6x9�=��"O���%E6R��`����@!����"Ol�sq�]�Q�*��M�*P�""O|%1����<��1���^���rs"O:Xk�d]3`�
���¨%����"Oz�cᓹƅ�.�[FI���!�ڮ�������S<Bp@��0!��"Q2E�AT�u/ne�B�9t!�'/.�p��ںj��Ч焾Br!��Ԁ|Hm��
6:��U����/hH!��@�U듪��}k��3��	�W!��^��m��l^]Ă$:b�1>;!�d��|Q��X�A���@*�6.!�/ ���U�w�u����~!�B�9W��at��4os@��ȇ$�!�$��f a��5qr|!F���(�!��P����u$�Z����W�s�!�0��!�">@M�I�8��� "OP	K�N�Cm�l� �.�("O ����3vf���s��~���cw"O�T�E!:�}0vƀzn��b�"O֬˴`:(�Ƞ��?A<Hء"O��S�Ew$|�x��ǉ�J��"OҬK0	̞i�|E!���Rа ��"O8|�b��<0����ʹim��k�"O�}����r���e��	 �×"O�Y�����mSJ֗KK�|1p"O�)*�h�'��(1
E�rANթ�"Oh��r�>�r-0g�!a�0m"O,��CN�Kk�	�D/�<G{����"O������2�$4 H�N}xp�"O�Yu�C�~F�C�Q�Cfr	��"O\�q�G�!\��g��)`
�Ѡ"Oȱ���؇c��	'��r}j��""O&��lA�^�� 1� 	�w�Jt"O��I��E  �n����6F�
s"OBD�!]tXhѫqOֈO�@�(!"O��r�!��@��#���@�"O��A�o�I<�1�t��l����"O���Ǥ��P�\i0��s��ixc"O��R��eH����AZ�@H�"O֕�P	��V��Cp���=ӂ�I�"O֥��<O�T	�'C�omP�!�"O��vʙ�Vo��zw���kb�#�"O��#��0c�6qH'�̢u]��$"O�q��@�-Z��T(�[�Qj�5"O��Aw�E�s�􄉈
G�(��"O�Y�f��NZ���E^�b���"O� �;!�h��pD�62`�W"O�҄��TIF1�5�ɯ/��Л�"OZ��F�x %��B�;'�00��"O�0�����6n��27_��up "O� .�ʅk��\�.�Rg�G��z�s�"O�`҃�&]#q�{���R"O�	#��C,��j#M�[g|��U"O�=��8�jp�G�)�2|�q"O��cbk�'C�N���\�4�`(qs"OLu	��تe�v,S��H��d��"O� 3���?~B�Z!�#Jx�u�%"O,���h.,��d�ͯ`¬��"O���V��>�	�Nи9F��@"O�X����)�涬Bq"O|pK��Q� &��6� ͜�b`"O5+�ިNsl��gV��<�v"Onȉ�BZ2��d#��J��ԋ�"O��c��&V���J�+s� t[�"O>���+� /�
i`G.gF�e�t"OJQ�$/M7\��Ź�M)��a�"O�|�uNN������@�Z����"O����y�d��.P{Y�t@�"O�Q(�c�R�p����(^���"O�4Ύ�kK�} �lߡD;��{"O�<P���\�M��,��G6*D�B"Oz10/W�s��M��jZ�{�hbu"O(p�t�I�Pِlx���D�b0�c"O�ha��9h,��PW%Ei��aqR"O�� �� E�V�i�Dه�=�"O�A@k�jG��{ 
X1����s"O�L�B�l���PD�*x
�"O<��đ+9?z�k�f�3/#���"O|(I���R�L���J�)>1�b"O���҉�2A��IK��q4"O�	��N��k(�7f3h�p"O$c!j�$t���J	 ���r�"O�����ސ1��A[2"޾<z����"OM�1�;�m�疇UM>�ٖ"O�\8 �ۏ;����S�Ӳ\F�j�"OJC#�%&�>���& y!��b"OP���_2.I �[%A2]��"Op�Y��8�����պ10�(�2"O��z�e��/@b��5$ׁ-�-��"OJ%��bO	{�D�Ʉ�!��"O�YXtl�:Usz��Bh��* V�x�"O��0M�1�^�`E04-�p2�"O��
��@hjd%	E���ap"O�i7��(�d��ǣ�7��;"O����E �I��L��嘽Q��W"O��zBe�������MP�ARLc�"O�4�$�P�V:�T�W��?^+r���"O.yM���BW,�Z
D#"O0`1��G-��(cJ��G �ٓ"Oq"��؄����)Ӷ"Opq�b�%Y�*�ԁ��D�y�"O~0��8 ��D`M\���y"O�T�bS5s8�[�,�z�x3"O�Ay4��7f�����hR�+�"O&�3�W	Z�8=Зe�'^@.D��"O�ٺ�!��*@���	L1^7��Y�"O"\I��&Q��!��b��|�"O�Q(��͕c¸I#�bMSlLl��"OBX��j�?^�D��A�L^R��"O��:���R`*��Á%C�D!	"O:4�lΚD�5p�G
$� c"ODa��S48��X�J���"O�D�!���F�P;�fǈ|TL<��"Of��q�K�%l&��&��-?\ �"O� ��¢M'����'v-��*"O>��f/P\z,�!�F�<VM;�"Op�c�Vs��'(���"Ot���:.DAР��<[&�D�6"O��Jo��f;n	ƀ�!ԣt"O``����&d�n�FM�2Y�-	�"O�&�Zp�:��Yڐ�""OH@cb(C�x���{�T*a�4c�"OVD ��4�&|b�g����*�"O* �Q"A�����DF�����"O0 ڠ�S����Ӆ K�����"O�a��%&GNd(��A��8�#�"OZ��K3B�N�u�M�F�"T1s"O�e)mA���0A��O5=��(q"O����#5-��HP�]ʼ��"O�5"!�3<���PcȾ*dT�"�"OBq2����#!"rŤ��gO:L��"O �;�&*�͕ۗ7HPX�"O�qcT���L�w�-�|�	�"O6����.��qw�ũ+2N`��"O&��&O��Wg��z4�e��L;1"O�3&�K�< rl� [��q�"O<����=F5��Y&j���)('"O\H����16��,��I���b�i�"OL�RE<�Es"Ո�q�"O8�0�̒	�:���fJ�g$���"OD�D�� ���`7�O�贄��"O`���7U޾�q�a��R��"O�P���l]*������"Oڵ����<�\�&kK%Y��,y"OR\��lR-lZ>Q����{�ni�3"O~�ňG�T��<qR	M S�4�r"O�< �	�3a#"����:x� �u"O��gEG�l1$]�qGX�g�D�"OnS�ꊌ�.D�R�G�SN��[Q"O������NE��E�<s5D�`�"O�H�f��O�,�dR>�,�@"O�őЄ�[ohT�f$��u�i�"O%B�'D�T�xU%i*�!�"OXX8�#N�TO��Pg�&/zP�"OB��	�m���c��ޯJ#�yP�"O0D�J��4�ލ�'C�2���"O�Գ�Ù�[�,Pb��4��tB$"O�qRk�-���(��f�6���"O���E�ӷ+�����D8�2"O^q�Uǐ?(��Y��  3��ۓ"O! �e�
P�t�pq˕<�Y�"OHy��W�X�L�"T	U-G�b��"O$�ꕩϧ(�F���=�4<i"O���C���aE����'�'( (aT"ONx�E��k}~� �h\�(�l�"O��%�}�u�2hT�u>��d"OZ)��\�F	T�K�E�.$ˇ"O.�BР�6*�Ό�G�h`�q"O�l)%�K8T����qB ]�E"O�"�Ɯ.)E>� A���̩�"O2��M�<6q��Ž%b(���"O���t�g��8@�m�u{,\��"O@���
ٯ1��X�,��%n|,�"O��g��8��C�;oW]�C"O&�3f��*Vm�У�1DZ�w"O)���2-�֩�T�¬@��%�d"OJ�Jc��"W� �ʖ�j,�u�w"O�]���ĺ]��=�@�BGу"O� $u��B<O��x��V0").��c"O�E[�J9P���N�<"� �"OV�1ӆ��a��JW@��YPm�3"O�ՙg�Mg�@1��#+� �"O`X1��<Tu$�:f!��'�Ly��"O��8V�M2Y��y�T��G�p�z"O.L�v�ԏװИp�
4�p��"O��$ Hɢp��^�*��iyc"O"�8i��B�� �/�=Vk��Q�'��%��#�1ŖZvb��-�q��'|J����zΨ�@���)޾���'���2 �ܬp��9�E�Ͱ)s��J�'�4���׈t�ɉE�ߺ 3D���'/dq25D��^�$G�AWB@��'b���SCY�X��px���/)����',��#���^�R��#!9*T�'��}Z��P�/��� *�67�̨��'������u�Q�c��29�����'���B���<,ƌ���g�2=(�{�'�쐸� E$R�x�kcb�#lĳ	�'��d9���=&��<)�.ػ"�d	�'F4tƧ�iM����"�,���'��9�G�
�"�����ڜ��Ɂ	�'=����*�$T$^�����|`���'>BI�V٭]8T��%��z����'l=0�mۛu]
��a�HkH�K�'+�MA0�8e�0��Ti����'�^:L:�,�H��)`H蔨	�'�T᠍�o�Aa&�]��r	�':�i��!�,n.�D�PG�]�����'-�I2S��5�~���&M�2A�
�'��ifeY�Q�$�qGF1O-�IB
�'r��f��t,ڜ��_*^�4
�'����Ʋ$V�����
Vd��	�'ǲ����/ZJ��SP>(ك	�' �D0�Έ~�TXOS?��!�'Э+U���1RF	emf�P�'I�"m�=1��5�@C�S��@��'�lCƃYX�� ��������'F���W)�-e-���d(�BB�"�'ݪܡw�1������^�E �4��'IR�bph�G� i�/·iZZ<��'3
�1Ɔ8R��2��0L\X�'��i���@N���rP��8'�v��
�'�>��
P�g@�����<,c ���'+�}�w��Y�4pSnY� Sr�
�'"��d��!�y����C��j	�'��[F�K0.�z`9�i��=	���'b���
��L�Z�pF��3g �	�'H��� g�[��9C&@B�7i��'�v�q��Z�a�8�eH��`����'/BQÖ�P ���eF:)� k�'����䃇��1��M:OT,k�'~f0�L�iXz���kL�L����'X�	��^9j"�`��l�w� ��'�d& 
O���i!�+n��<y�'pb�Y��ϱ.@�Y� 
5P�~4��'펀��&<�:�;�LŘG���'�a��kܺ��C�C��1[�H�'yV4�򨌄7<����=F)��'�d1��H�u�lmsd� Bw���',<�Y�甩{$�"�JR,3O�Ez�'*yz�M8s*��z�)\�#QhK�'��T)-�<7XEрE� |��
��� �U�K�k����D+Ա=5��D"O� ��2�<l�p��-(i��"O�0b�F�-r`IR�j \�BA"O����e�H��h��Ȟ�^��� "OՈW�2O�����V�"�!�"O �j$%	!qȜjU���r
e�"O��C���P ��ǉ�@dʝ#U"O�3��ȓ�F���Qb�3�"O��*��?jĵKa�lB���q"Oz��H�f8R��cA]7��Q"O��xB��qB>�:���$'�(P��"OBĂv�+	�ԭs��O6c�t+�"O 5,L�(D��b�m[�]w���"O��!g�^�i�X��4lcZ@��Q"O��2�΀D�Mb+ݱ`+��`"O]p�IY&!�u�T�S�U(T�v"O\�� � O.`���,,���E"O|qرg����	((�@"O��"�aA�e7����W�
�*Ҥ�y�n�I�����C"���%�y��ެr�L��`H�5񄔻W����y"F�wt4q���<'h�uK����y�+��"
d�r3�:b�)"#��y��=o6��g.�Te
rh'�yB�R�V��A�||�Ôm7�y����̴`���L��ah4���y�$��I�d�0��4&�D�s���yr�!=��:@o�Z�b��	�yr�ѝ<�u��� 8���/�y�e�_oa����Z��3$� �y�'E@���T%�	��p3��
�yBlY�	�D)����y�����ǲ�y�ǜ`�(�$��wo��ӑh�9�yrꋖI%&!j��3AN���!Z�yR&�;-p,X�N�=����ۊ�Py�0vmK�LRF��L� ��f�<��	�w$8�z�m��Bxa�Ad�<�6�W��H�ir ��(��p�b�F�<!��E ��i!�ˑ�NL9����L�<� UO��I9��ӂvd��a�[m�<�S��)G�԰ٕ��;�B�3rB@k�<Ip]�
Β4�cKA3+�V�� �m�<�g����0��.yvz�)Q�^N�<3�\���0��VKN�9"�M�<!F��P����Ε4�Z�)SA�G�<Iu��",��K��l�j��cE��<�׀D���91�^�4�s`�C�<�dmĶ!H<��M� wф22|�<Y�BȅE����&'Ð_�M�W�B{�<�GfүȊL�Bӊ#��`0a�z�<����"~�d`{DK�DȄ�e�y�<�g'6��X�B�3J4Ա��w�<��ҭ@g0��T��Y��	�5��j�<�S,Գ,��-H�E��ݩ`�Wb�<�U��*@=G�	B�e�<IeF7�ͩŌ���i�I[^�<q�I:S�,��� �4���`�*K[�<�N�=f�5�5�[�f�48uj�B�<q����`SLi��Z�W��ː��~�<�d+��j)�"�b�ީ[�H�y�<�S��_vrd���g`Y��
\w�<��� ;��1R�bܛ]�ybV�Ks�<�� �[H���C������F�<�KV>MY`���Ɩ|:���Ō��<� l-#6&��6t�EV�P�<�1"O�m�d_�\X�2d	0s��)�"OЌ���ɔ����ǩhA�"O���Vꅇ}I$�Gc ?B��e�"O&���/�,j�B49V�  C���"O���f+x\i��V�G���"O�Ez��G'n�t��@�W�@�A"O���UJ�R�C�N�eW���F"O�Ȋ5
�8Z����V:E�pJ�"O��K�'U�yX���������e"O�I��6V>|�b�oA� ����"OD��̀����g�#&��E�6"Odl��M�.iHLh�&�	>�h�"On�s"-�#��m�$���1�v$;c"OH��wI�-ֲ�X��ڵ�*l�"OD!`s�W�Y��ٗOˍ�e�"O0���NF6Q����%6�	�"OB�[�����r P��9�М�R"O>d�S*_	z�xH���&5��9"O�����`ʂ�SgdN�>(��"O��&%�e�P���"K+9�X�"O�$�Ž_eܽ�r�ć���:�"O|8��l8 ��Z��Xy�"Ozݑ��@^��o)nkB���"O���n	+w���ƳP���Q"Otb��O�-��C�1}:�)P"O|y�E
]1e�䱑�㗠V��	@�"O��1��J8���b�9cq6��"O40QQ#X�88���N��8z��['"O�DKD	 �C2��)�j<w��`Y0"O���"h�^
��
��FZ��`�"Ot)��N:���J�UR�9(t"O�0�F�Ïm#��s^�*0��"O�{p��p�FD�fA,`t�'"O��#խ�i�H(��.χ֖�J"O&��ck��c���ڗ,uh�"O`�҂� -˚��'\�Z[�a��"O(p�#n]7��2�ZP��E"OĐIUMCS�� �w��
L����"OԹr!��9(&�`��NBL �p��"OJ�G��K��a��5P�EX "O8쁖�ϊ1�L�"ϿHPE�3"O�"�E�%d��Za�̅n��Hc0"Oy�1���t�pȂ%��	1�pŬh�<y��L�a ��R ,,g/���$IE�<iՂ��?c�|J�#)F��Z$�@�<9�)ҽ]��`�Ћ�;Ą�����x�<I�F�77L��F�=-Hθ���M^�<	�ψ;������5^� @��/�Z�<t�Z&>��Ԩ�#�1{p�!QŎk�<��A]�\Ř�M0#�n,�Uhmy�)ʧi�$Q�@5���*t� NL�ȓ.8PсqKO=h�`��@	�*��!��m���A�2��VAFgAvȅ�JB���R�]�_��}�(B<�<(�ȓ����c#��v��H7%r���?���)�C�X���M I)A��9�!��(܊(�%�',�!�&e�6�!��O�z�� �W�\.�٩ e�4-�!�͝y��QRĄ>p��<�Wn_,�!���/�
p�֩ڠ)Z���.��f�!�$ܘ����� o�U�b��H�!�$J6J��Ԑ�O�L��);QΈ�>!�$����a�Uђ5{�/F��!�� L��R	B��%�Z*&�>U��"OLx2E��|���1Ê�gd��T"O�@��\"ڢtA�	�M� �"O�Z��ɀ7�r9��JƬ��	�&�'���8wbu��E\+h���(/��!�$�F����GN�U�j8�N�>(�!�$�o���C,#y�yrw��	�!��ͿSp|�rn�8F�,J�F��v!��ћz�0+6h	?�$�'FT�bg!��+Y@��g W)}+���Q劔$e!�$�*
/x8�3�ߘcBl�3b���UUax�퉇7�DD���J�F\@)B�B޽�<c����I4Y)��sC���>~����ދn�C��($�| �Ԥ��6���8f[%X��B�	?	��%�A�o�
�R�&��B�	1H�L}���4c�H�4��"S��B�ɮS��)9�Dֺ(����#O��vB�I�{�X��
��>���3R��R�H�?��**�'��{�H!0O4��1)Ӓj t$�t�!�'�
Ԫ��J#T�qA���L�\Yr�}r�)��P�~�B�,1Yv�z�Ĉ+8�$Q�
�'>ȩk��	R� 8��`�56 ��:�'LHx�OR;��Y�� �@��1h�%� ��(�6D�8Jf���1T.�H!�
�3�� {����hO?�ă<V���q�*�����ш#�!�DG�.����K	�Y:xTML!�$! ��Ż�N_�k������*F!�Ě�j�RI����G��j���G@!��2�HE�GLS�fQgBw�BB�I	*���)İxY<�X"� *1�C�Iͺ��ĥ:�Dq
f��I��C�Q|����L�q����*��C䉏+p�1X��	�v}c�	P^B�ɕ'&���3��=#\�i����bCZB�	�8 `�xV�PI� ��B��C�0b�������p�J]�TDԚ��C�	�t0b�RVN3'�"���FP��C��!l:�	���Ҍe�E�(��G�C�I?*<�Y5,#Sd1��R̦B�	&(KFmK�޾j���֍�K�NB䉯\JN5¶�B���Y%��
:рC�e 0h��QC����VM�0>�HC�ɤ3�|P�Wi�/�X�B方?����5 ��@#���҉�JѸ`�!�D�w[Z�Y���w��<�@$��!���GJ��umOp���&�Z!�!��2��E��*ն]^Z��qOڲw�!��%	� �BڰQ<�W�L5I�!�D�8*�$�`\por�O�H!���r�,����R=m��83�3�!�d
�nAX��@B޼RqM�!��E�'��,"�����:��;~w!�$�Q+\�aE��j��p�Jk!�$V
@��I*p���X�dtӠ���f�!��5"2\��&#�����+� �!�䃹#8,���'�`���Y��D�=�!�Xc�HYC�#G%|�dCto��V�!��+@X�9�-`p �p��}v!�č�+�P܈�K��xq�h�5�Ӱ0\!�� ��e�ՅJ-{����p(!���o�@�ۣ�No��au��!�d�(��⏋scJȨA�E�dW!�2ZN�*�l�0+�;�(�.r!򤛬h�tQrt����H�`�F�j!�� ,R��m[v�eG�rw�1��"O�e ���8Y�<�v���x7N�2"O���$0��#䉩x��hi#"O���fŔ�#�$� ��)�ƀ��"O\�j0�H�vnX�P�A	:n�ژ+�"O`H��D�f6��灈�PS��j�"O"�G�d����R!���Yk"O$�Q��A�#v�X� ]	M5*���"O�����@v��W���-�4y��"Ot�QfdV9~�2�g�R8o�bE� *O�H8@� �R�lU(��J�=��D�	�'��	aIH�D�S $�3�8uS
�'P�`y�i �)x��p�4�f��	�'ŔEk��_:` ^���%�,汢�'��=+l�>44ȝ���K�up�r
�'�h,2�X;G���Q5�D�m�&p*�'��� ���1;��#���u�̌H�'�bu+�g^�P�n�K#�&[���+�'<�U�w�O4m�",W�<M��'��IuH���h8H5�"0��!��'~�@J���,M 1Q�!��x���'.PEj!+K�ra:У#�M���'�����B5`�z}0�$\)q��X�'���"-X�fqz��%Ex�����'�5:a,�h�	���yI΅�'�\���G��B����`�!f��@�
�'Z�h5i�v
�H��+X��Q�'
r��b�P���]�0�"J���	�'��ݢ�A.;��8+`N�;�&i��'Ѱ���Z<��ՌY$]����'ѨȱAдUi��ߑb:��
�'���s���8��.iԑ�	�'z�rG�T,]ҨC��d�c�' ���«ٷ7Mh�""Z�X��'���[%YF|� CL�Qn�8�'Y��N��Eqa(�2+Rqh�'����n -��q�����`q
�'5z1��.��� � &��|�	�'>i�uf ��M٠�
0ā��'�����$)�p��n��1�'��HW*	�O� ��(�Yp�'�`�a���g�,� �-u��\*�'�%���"{���
*t0L��':.�����O���8��2|�V\��'������I�d��C��@lթ�'a��׏I� �����n�U��'�FjU-C-P��;!�V_G�p!�'� ���H2 BJ�
�DY+�'L�퓦�e���1r=��'^:@�ŋ�k�	�U�[�b�H[�'$�4	B Z�|� ��yO�H�	�'��Y`��+g�������X�'���R�+��Q.6,٠K��RlIJ�';& �ϖ*
�`80�H,�	z�'�H #������WF��{Z���'��ٲc�P13��As�Ꜵ|!��S�'�`foĎ���`�iz��i�'p�#'
�{�P��߸^=���'�8��@*U���,d��T�T��J5"�&� �\��!d\#]�`Y�ȓ%N �����` �@̾U-}*��-D�T(fAĦX7�mb���G>8J$.-D�(�p�ܿW[�i�AU#-U�����.D�IC�T,N��-{���99� -)0a,D�� &e�ehT�N�\���m�y{����"O�q�-��8"�5h��[�"O`1j#���6�T$x���@Q�	�"O�����ڼ��A�d8�H�P"O4�9fM�
`x�0��	^�ca"O*����(N����f�T�>�2�[u"O~�8�FN�I=2���Ƀ�B�A��"O���&�!�
�SFi��#�8�)�"O�����E�����D5s��c�:OF��ꜮXVVhK�H\�Q���U�	�8�di�,jq�@eML	�VC�	�^�Y�=oT�F*��;w(C��fI y��
�#6�
W�ܠY��B䉮Vc4]�`^�b�8\�� Z�(=B��(�4�@�T6�^���_�t��C�ɡXK��т(M����eݺeO�C�I&=���z��ݭ9!(��a�T�"��C�I _Oؑ��G��h{�~�BB��Vp
��I Ø\q�/�3~^B�&`�,���S��!IA��m?B�	�R�D�Hbe[�$�vEp��X��C�	<�iqb��2���&D���fB�	�|6� �B�4�%�?O�NDJ�"O�!˵	C�/,aT�7�Ɲ��"Oht����"��M����n���� "O&�8dү)�L�QG*�� �R"On0�p�L��h�M��'��@J�"O���-��z� �`�?��Ѩ�"O�� U'j�@B+�?zq6p�f"O�����HM'p��R�2D�YUeDz�<ɵ"�'g����,s����^�<A�A�WLd1s�,R'\�(š�@�`�<Ye��ʽJt��Y�&���\�<���P��SU�>:��h��NIT�<���%j���5= 6Q�q��P�<)C�
~@��5�:�IS�<y��J�z�h�a!�7�����V�<�p*Qj�8� ���-2��a�0ɘQ�<ї���R$�&d�-U9�0��V�<	�͌�K��EEƅ�F`(���h�<1j@f-�D�nֆm�ʅ�Vk�h�<����|4� �,�8K�Ɛ��N\H�iЗ C
�ֈ�d]�"~�	�=H���e��`:�}��	ցu B�	*�yqdg�.�S�����FtB}h��Ѱ�V� �>O���!�K:��D&ֶm���1�'���ʆ�#U1���uC/Px�̣@���� �CF�_����'�|���HB\&Ri,�0RCԢ&���t"�	C�x�C�#�8�j#iD�1%>���޻Lb}�g �V!JL���"D� ���I�@���yf�S�N�N J�d�\9��8,�d�4��t�ĢN�#|J�੟S	 ^��g͉m(�Ah64�ж)�9u i�U�HMu�ń�m��h���_M���XI� ��I�V�'C���Q"��k�-͝W�A�˓:�@8!�fۛ8��R�H<g`0�%��i35��,��j����Z
e���1�O�į�5\�Z$�3%��Q�h�J7�x"'�4%�r���%����K��u�TSʗ-S��)-x����26��ˋ�$�!�䄥}�V����^�u����0�WaBD��H�?Z����/ɾ�v�!� �~�T�'~���s�a�)ńͺ��k񈁄A��![�@?��r�� 	H |
1ᝇ&���0���1�� ���C'�Q82�A	�(8!shK�N.\J��<�I�.����իɹQk�m!��W<e��D�/'�L��ǅ]�Z��Ih��
?c���$ˊ���ܻ��Â |�|є���J��� -?x��{����-�T�ê�&x��I��ǵ���L�6��r��n}dD3qBouL�t/�?+�����<�"r�ϫ���0���"�&��F"O�H`TJ�+��]C֪G=}f�5�¤�C��������b�l��W�\3,M�FhW=�����{�Ā[�ei���P��`��3 OQ�y�˦m'�O�ۖG�	��8v��+|���@�I���T��%ޏc�>��W�
s�a�*�V��héx���(��&��S�? �=�#�J�pp����g��s�]8r�#Ռ1�cCJ�rt��Бg˝v�iH�m��99F��D�!$��[�LV>��S,�|N
j� ʻ7�l�Ї�C=�ax�Ji U[c��]F͒(i-T��Ԧ47C"��5��*�pI���Mg:eä^AٲR�V�k)Z���K  B`}��k�!Pe�|�"FK�`��2�'�0Y�g��yan�Yr��zP���!�@rlЗ��#j��Y�I�(a�� �xaj�yJ\���w�Ԁ��ĀV/���R��2�MYߓ.�lM�@�ܖq�Ġ)�jU;h޼��o$Pu��'� �M{'pW䝡�� >�t�B�蕫u׬]A�E�N���sWi}2�>h��ɀ�� �K���H�n�5��'K���F��y��Iہ�A �py1��nI𭃧-C�GHdf��1kL �`�֕~&�A�@�c�D�P���NbE��BY�'�F��\I�N�:"����Ұ˔/?ҭȴ�/G)A�Q�̢�Rɚ�A݊M�^�
D���$�0�,81�y84�&����$H���͠��A����	�d���/��ś�A�zɌ�i�!%i�"�"�^=�-ȗY�D�vN��.����@�~π�؅$sqÕk��G
٫e��Q��Zۓ{���C`b�;\��$�6+�"x 0墎8%��T
`�V>|�N��`A�V$�s2jN%n���id��A�}�	A��S�������x�[�홌i��1��ݚ^ 8��>a�&W�M�F<���a9*��#fзult�ؤ�Ű�����Ώg�aYD��#B!4�s��+	���@�/ДCjB�R��������ϓ7L�E�$L-�:$���ϛ-c�(AC��]Mޠ���B0��bO4K�]�e�/�20��+m�sD�!%���
����@V�ɑ]0�"�٠�p?	ծ�	AÐ0P3LG�3�<4֮��R�2���2�h�r�.�fઍCu�B
Eʊ8P��7�(KVn���P�I�(���*W$ϱ~~��ir@��a{07K �Y���e[�9���E� ��]�&��e���#åI1O�X8[���iM�TK�i\�2^�۔n�1!��M�vN7g���;��O�MJ��>��d/�b��T�"�"�O�u1𬋵M@��f�&x��3�ĚξT���5I��l���<��l��kX�f1�6���2�� 8��D�Rk��e4�P�����0��5��	�T�b���*5*� C-�(� -�7�Z!T�D�b��1��9آIS�U�B�!.<>�@c�/u��sU�	(0l
 _�1��r�)�p؟�X�M���R�O>?ʵHe�ݦɠ�,7����Sa\
Wf��h����B�Ϗ��MC�J����&ϭ~�;��G�s��5�P�]X���T�h��{�GV�r�&�c/�X� ���HM8��� �M 9������Ѐ�Is�"��>���£�W�,��ܛ]���EyrhH�?�����mڔV�(�|R�Й�V��㉓A9R�$NV?��*�K��тH&ps���d�Z$6j�g _0�I����;hR"C!7y ��%#�t����/v#��:b˄�C�H�s5w>>���%[7} b 2�'��pr��R�@����n���kJ��rC'%;���K�' LY(�{�':�p�Z�@�P���I��J�*N���b��TH�	E���Ԧ΅mcȓ\h��;��Q��!�K.D�p����hAe�DS��yV��(M8n��ȓ[^P��VjP�}�x�������ȓ���z#��F8s5e߯)�D��a��T��NO���|�(��S����XM����(EA"�!�8ɇ�Uz�H���Ηh|2Z�n�!0ڊ��)�B�wō��,�a"���,
���I-�͓u����6+�� ���X�܄ȓ��������
��Y1
� ��pFz�'QMp�G�4��]AL�J!�|z��h��ҏ�y���G�(D�n�/kX}�$�<�M��чm6��"~n�P�� ���6�@1��O�u�~C��	#6P�;�\�bJ9��L:Y��j�D�H#J9|O$,+`-%P�\+��S�$�M�P�'J���AXğآ"F3s\���g+Q�U����¬3D���0'L7ek���
*��9y֌0ғg�Nl�C�;�'���1�͢HT�z���&S�,�ȓ`jdIF	A�H�V�6��oV���e���?E��_�Bm�<cU�ފAԘB�F�'�!�䔢3����N�lڠ�e$��R�!�Č�@�F���J۸9�����!���R�� �0m�(.������!�%T\f}�$ʀ�A��ZG�ܵY�!򄛾H�xՊ�e8؜��.�%]�!�$Ȳ(�&d��	6jŔ4�M4�!�1"p���m��x$񐍎�p�~r�DBǊ��� 5�*Q0Q��I���2w��[�<9���x�� �!�6�YpU�]R؟�Cb�ɟ�� |��g�65ԑ�1*���� ��74���e��(ꊅ��+W�C�.|z$B"D�����)�&���T�sF(����"D���#�52�h3ϐ�3�ƨ3��>D����C��]��R�N�xB,ڷ�=D����e@X�lk�J��k�x��g7D�8�É�)��)����$XĲD��E2D�|�u��"1D(�'�*o��@S6�1D�Tأ��&H�U�e��$:d<��.T���4@����y���63���"O��{2`@	����՝6?��y�"O><�A��tǰ�@�ՙShU��"O~H!v�<h�F-!�E[ 2�PB7"O�h؅�%7<t}�t!Љ"~Ը�"O*y[g�?�ت���x� �0"OZ�eK��/0xA6�N*@�ً�"O^�4FGtYt�� �R�B�ʰ"O֬���Q"���y!�E
&�v�S"O�`{�F�QH%�h�1т���"O�Ѡ����8G��!�ϸwǀY�"O��&Ā� |��K�G��>)�jr"OH�G���L+�\Y2̗'����"O�M�b��t\�f���!;P�
t"O���UB2~*���p�1%Q�"O��@�ʇ�t e�s� <?��Z�"O.���8Ė�� ��E)ҡ;�"O�U�'oÖ*4�M����5R��|5"O ���CO9\��1��'0��q��"OH̪)�F�ʭJ�9��K"O��R���P�(Hh�,@-D�P��!"O����D�E���#�����r "O$l��ʼ4��B`�$pi˵"O��� E�t��zF�
��1&"Oڥs�gX
S��r�!ڴ��"O�โ���EZ"�ݾd��9��"Op ���M��PD�C��m�l�i�"O*h{����T&
<[s��Y7B��"O�`��&G=O�a�l�1DɃg"O.��OS,c��i��\�!�Ry��"O���Sa�����&������`"O<͛%�̆"U�u�6l���ɳR"O��8��4w���ŉU�U ||S""O���OU��=�4�|܃#"O�K��Ĳ,��1Qg�M�p��"O��c��,nCE��70n�s�"O�pyÛ�F�[2�!O���d"O��*2��8�L驐�����!e"O�t"a�2;���:��̙B�~��"O�i�`A*JX6\AA�-A� �;"OlT���U\}���ǒ���"OL= V�N�)�n 2��3���z6"OX�*s �0>,� ,:@(�}�6"O�I��N�1h (5ѳk�y��pW"O�h�a
 b4�q�SJ=+@]c�"O M��$���CF�Ҝ�!��"OD�h�GW�6��[���{�,8�"Ot��D��v������<�����"O�љa��a�0Xq�����#�<I�o$x�I��j��7w蕉w�l�<y4���ML�H��$��t/�Pɰ��f�<A�j�Rv� V��W�,D��U�<�C&^����(��F�y��j�O�<�@�׊q(���c��{< ��5�@�<�p'��yO����L�d��%P5&C�<� ):��P�omR a���0�2"O>DqGf�+	/T�h��f�ИY�"O�����	��|
�OBK�})"O�8�I�'@V0S�E�' ����"O��A�J"��Q��o�hw"Ov�+��K+�X�T�BjĚ H�"O𴣄+��K���C�?\��A"O���P�F1Ct��dWz��"O��0��ny���E�T9ȡSD"O��ҕ%�"!��x����!'���"Or)뒍�8(�&H��Z a���"O.9Ib�E�W6�Ԡ'挭�鑧"O�� ���`��R���"O���W��F���Sҋ3 ,��P"Ov�4�ɵ"�@�!6�+aӦ"O��b ���83t������s"OVp���ۧ`\Ԁiģ�\��"Of���b��-1�UJԂH6z�`��"O�!crJF�v��Ӵ�ZoL,�&"O�(�Ίp��(�Ѧ��u\"\a�"O�Ac�%T�M�7��[B��b6"ONz�޲�l��֢W2c��1p"Orq	��ͅ!#� %���]�`�"On�����Q�h����B�=!�"Or�*�$C�`Ѻ�_�E���"OX���bF��9R�� V>�!3�"O��D��!w^�����ltV<A2"O�T0��H�U�Dy�A�Zc<��#"O01�R�Bq��	J��S53d%��"OV����G�it1����r<���"OM��k�{R���.^4WGb%{�"O�-��� z��@��1O�<�S�"O�	� @Z �y ��+ִ�KQ"O�H(�!�:� 1�RS���A%"OtsMU�B*ތ8��,��ċ�"Op![Tm�0X;����� -��q�W"O\AI�9���C�)�<�B"O��P�����������>U��"O�ic@ [� ��I=���D"O����*��
�h��aG:Cޥ9S"O�9�g�\(�������Y��"O��R�U:��i{%���/���"O��ˑ/��	6J�s���r��i�f"O�8��d޹e�&��V�|��Љ�"O|�q�f���m�!x��P�*O�y�U�V,��1W�Hs>\ �'y"��Z�*MD�w�#ua��R�'oT(���M�4G�Q�H��)�'Ll��G�Z�y�Fa�}Y����'�Z	X0���+�S(��Z��?D��J��Vg �a���=L���+wA=D�|����=t[�A��+�5B`�r�=D����06D��`,V�K�@�s�>D�Ĉ�C�I5h��IN�s�>D��*�F΂Ri�u��a��#
X��c?D���D�����<C�8 !A�:D��iaG.�j�ri��XFB�C �;D�@B�*�3=ځ;Q.�B���)5D�tA�ڵEk�}qG��.K��5D�X�#j�-dD��c�	�94�Y��7D����aJ,,���$a!�-Y� 3D�X@��I�e��i`��̇	���uL1D�D@��
z |!��� �@e���;D��ba߸ ��p�`M��A�����K%D�� v `�H����'�*u1"0"Od��v��'V��I�L�)-w�Ⱥ�"O@Y�fլG*Ш�lĬvE$�(C"O&I8TBD��,%aj�/��X�"O�ѫ4ǘep�+Ťɶf`L"&"OģuF��%H:�� �@�]N!�䃄L-~�V���i�r����A�x4!�dȳ$ �u+#�|� ����:!�� &>�"eA���4`TB�> �!��wI$�+��H��SǢ]�t�!�D9]hCI@�P%1H��U� m!�B�T��F I�&aԫCMC�1>!��	�()#��7B\v8%�
�x�!�$�6wE�Zb@	�Zdr��*N�h !��R�l(,ҕ$�|f�(P�^o!��%i�DrJBW���f�*F!���mP���;!�*�!�D�F8!�$ڈ�:�ࡧ^�?�t��ƍʫS=!��6���0%�H�<�����!�d�	|�|p9W��w���I�(#!�dƴX,~�W�x'�ΰBw!��2�<)Ѷ�^�|�`�;ׅ[2n!�d�h�n !Ei�T�&�r�D� �!�D�[j�s�Ǘ,;=��C�d���!�$�v�
R$ Ё`n���=t�!򤏨&Q���0K�>a��<(�!�䕃f��K�a�7CQ:�ް`��B�ɼP�0h��I?l�� �%P�Ed�B�I�@�\u�6��6#�\!#�01�B䉹#X�y�ܥ���:�%�i�B�,`ު}� ��|�<=k�b�J�VB�ɔl�L@ї�ͫ	�A�"��?(��B�	$d/4}�����2��Z�ʂG��C䉎A^�Ը��1<�l	�Î�<��B�	�/�p�[�Li �YVn��/{�B�	�k�1�eYV)���?A�B�	��\�Ц��/-@	Q�k��C�	 v=�8����_�U��B���C��"jY\���K2oq���%��qe�C�	'�YE�"s̐(pf�^�B��	Z�bE��i��6l��"ɉ�|�B�|2����v$2u�'}�@C�	8?ip3�9V2̘6(T<�C䉁
�<ey�h�,T���� -�&B�"D
Y)vMG�,+�	x`�ˊ��C�8L���B6�
m�|���F"��C�?F���T�A#21\ /C��C�IC�$l��ؿFj� �M�:�vB䉊y��shܐEyz�A��bFB�	�"k^���%� ;e\}X
O"V%B�I��z�{@�O�&#~�كo[�Z�FC�I�KY�1[�C1PZ,�����8�^C�	s���"���5�k�\>C�	�-b��
�*Su����
�C�I�luJ��eCU!� ��K$r]�B�I�/�$ء!��>n��ũԝW�B䉰b���!�D�I�RT���^�B�	/n"N�9AC<:�*��f� �JB�I���(R��B�(�fE\�E�dB䉕������T3P��BC�6xfdB��9)�� �AJ���	�cĜB䉟Q����>:��q�2XB�ɶ���z�L�rG�ijB�	�ȡk��${�)+�cF	G�C�)� �ѱnI#���#@H]c$X�R"OJ�CD��pR�D[	�E)P"O�9	֏@��F4�'O��V��u�$"O@���. (0���\>s��X�W"O���h�
^h`M�'3@���"OP!#BN�9�@��@�YKvQ�t"OV}3P��1-�T��r艍�|��4"O8�(b&V H�^��S)ֆW��!2""OD�(%W-0�`5�敯����"Odl6oBf���>w��h�"O�Yx���,%�2�����m����4"O�@�RK��>�^Eqg���E��`p"OѪU���<�R�� d��q;�"ODMs'K8Y<1�a+܅ڥ"O$Ey���:���AdŗZw2}�"O�-�۽k��Y���$2*��e"O̰Jbb��3�ᓣ�9'2A�"O,����V�Rh���-~�("O& �v+�$_��e3��5�IPD"O��0��D�Z��d��z�A2�'���bY�t��O�+v(j��'��1x��K��YI��Û�����'����h�EW���%�#<R���'5J��1$�*-K�F� ���@�'��m�����g�P�yyV����yrA�=�}�� ?�B@z��y"(Z�%�4^*�P���T��y�-	X�:eI�эT�HК��yB$XynDk��A,p��Yv,*�y�D9%V�p��ₖv�f]"�O��y�I�ju��#��6~m������yb	Yfha�)Z�y���Q����y���
JҸ�'�{Ȳ� #��y�a��QcC��{���kqd	��y���up�� ��E��!m(�y�'W{`�3��U\����yb��"6s�́�)M.I���[qN�y�" (j�y�NX<3�4�����y�O£Q �$�`ID!� h�W����yrE��0�n�r$�&l������yr�W�U�d��Q�ӻ	䞵6�A,�y��WމIP!|@�����y�-��4PS���Ɯ�X(V��y��͂��ի�P:2�M!E���yB��	BE���P�@��0�e��yB���9g�,�媑-)ࠢU'��y�d�>"s*�
!��?,2�je�H��yb.7n�>�)R�W-��P��D���y�P�,��u�p@��-O|���y�iӡ;y�x��l�P��@�� �9�y��/:�z�JȡKr��׮J�y�F86@�9��4C�b- G�D��y2+
8 4ze�V� ��%ֳ�y�	]<5��xD�!>4|��L�<�yBA_�>�d�:V!υ(�=q�jA�y�aT̅�w�G�T~�����y���ؑ�c�@�@M�YY@���yRe����b���/<k�e��/ٕ�yR�_�q�Du���ѫ7��Ɋ$�y"/3���s�AMVX�@�4fC�yb��3vۂ�Q���H(�]�@��y�Ĉ�&v��
@!��V�!�b���yB��Z���!5��Au�R��y���t,���!��r�xe:bŀ5�y
� z�ѓF�Ŗ%���/O8H{�"O,���"2������JGT��"O���IZ�*I�:�jګ&^���"Ol�X�I��p2�h�I��Y]8
�"OHh�eh $'+ũ��Z#@��"O�ݲ'��k�)3���^$)i""O!&aÅt�~e�P'B�l�E[`"O!$G/o�Xy�bH���� "O̀��%V��H(�4�Ys"OXBT�M����2(�&��g"O�Jr���:������ �&"O.ȸ�ͅ�$�:<R�j45���p�"O��ra.ګ|"�8����9J(dͱ�"O��0fN�r1��zBA@`��9"O���vD�*V��x� ��&by��2"Ox��3�R�.���+��˒~���1"O�X��b��I�J����b78O���K��9� uX@ ڪq��d��M��M�t��\FZ�ʳ��	in ʓ;Qpa����]+t�<S�!��g(.��0OD�ܱJ�)��%��q��B���!0�O?hݺf`�&L��:r�
<�+壖-k�i��I�O�T�C�0�0|��	��2�:��4ď�a,MY�HU�/�� 3�'B����E�Va��jX���_03n�S���x��������	#Æ�(\Ł�..��`� �2n�r�=+}D���K�
�:$�f�ު)6�ܻ�g ĦyE���k>�ZO@9tBP,SfE�2x��i�I� �nHʦ]��,^)p�Eb��)ހTa`���o���Bc�Z�A&F���1�n>*5d堅��P>-��Z*9�̪4�Qs�|�Fτˮ��s��,Jb�8����k�N��	J
B�"y����@O��!��(��'Ўe��������@ �O�5A�ᆁ�ё����^��s0I�l0� [�9�(���]�B%��>���2T̀�QpL���D�T�l��3�Z�C�|q %gӶ� �'z���p�Aed���ֽ=�����ڹ��Xvaf� Բ�����t�O��0��HQ%2;tL �A�A��ъ2���5[ax2��m�f�6Ǎ4�x���y�k��3"p�$'��.�z]ڂ�Y��y� �0�x��a�t.Ѣ$���y2L�=��P&�:<�]9k�6�y�郦YR$���Ҕ��18��F�y���zKеcg�ϴ�06�¿�y��̓R�Z��� �b�{�@�y�-��0p�G.�.�5N��y���,(�Q C�Y�b\i�	��y2�ȸ�n�����%|����!� �y"Eϭ*:����n�f�����y�E�)wC"��aܐaR�P�>�y� �UO$��O��1�24(��B�yB+
�Y;x�B�*$���i6@Ʈ�y2%Єn-�5���Y�k����D��!�y� M�j��q@E��z�Rœ%l��y�f�-?�[��؁wόl�����y��Ǳ%�!�&kA��B�y���< ܎`��@�>��8{t�W:�y�B0�R���V���uQA���y��S�,�a�G�=D�nH	1ȼ�yr��U��iH��@�@�����ǒ��y���mrP�i�BY�3�$16�\ �yb+�*O����,��2� �"*��yR���F>V�a@ǋ�0.�8�"�y��F%X��9[0k'$�%��e@4�yb�Ȑv"������4L���H��yr�Y"I|���EH�j�p�I3�y�n�<�Ȝ�@ Gn�"C���yrVK�d���4v.HX#R�"�y�&0���9�h^��z��\4�y��y���B�+6���:����Y��,��-��Q*�6���G�Ъx����S�? �}k��ƨoa�܊eHE/b��@��"O.�d���[�^{���04�l�K"O�U�ҢK�M��8 M��r��y�"O�0�(R�u�Df��1_���5"Ov"�ʛ�=0�EH��ņ2U|�KC"OF���,_
#�P���lI*@^�9)�"O�hz�� ��0��<E���"O�͸3	�="�-�#F	Un�A�"O�� ��4U	�1��TL� n"O�)�m��K�RE� ̓sL����"Op}�3�$��kF���0�"O���ÚS��l��GT %�C"OX|hԡxs����U<=w���""O�ԃc�ʩ
B�A��r���"OJ�-ެk��z���-A��ZE"O�]��MӉ)�L��1���P�lp� "Ot����^%u��);��Bm��"O�d"򤁻O��	u&�.BQ~$��"O ]�CV7)NN�1[727�e�u"O�]c���l�hwd>:h��q"O�#r�AjB�(�A��e/�X�3"O�ͱg�0z�␕?.P��u"O�ȳ�@H�&����,0~3A"OL��׹!=T���8K�P�"OԽ[d!��P�T�s���f\��@U"ON�1*�C���J��5 �p�Q"O�ȁ��Ƃq���Jf�\��}�""O�m����RO4pR�$�':��t��"OZi��5j����c	(j�2�"O}��,�4]�zQ��E0-b���"O�t)��;!�p�w�HIGY8"O2"�f��@p!HB̨|F�țb"O<�ԍ�9�d���\-)z!��"O.1�&
}�Y(��C�e:����'r��"/�pyvb�:s�Ru�ψ�s!��_�)�V!I`��!y�m�.�s!�$��E{b����� 
J�Y�&-z!�ċkL1`a"
�4�RY�t���2_!��ʓB�$�b���$��4+�/��w[!���_5�	{6�I ��I2$R��!�9]�z�����%r�� `�ҫ8!�G�hb 4�����r*��Rd#ãK3!�D�v\~U�t�50���Θ!�Ւ�����gy��4kT0(H!�䘎Ƙ��A�\�b ��[�YQ!�dH��-#��J�${�׿[M!�U�,s� ��P|#H�WLb-!�$������Т v`[���8~8!�dA$�Y����@/����cC�SG!�d�]@*�BYa�Q`���4:
�''^H��D2M@��Ԫݎ'T�*�'i����FS��Π�iG�v���I�'er٠�HBV�8b@A�2[gni�
�'�h���,�#qΤ��6��a
�'���k��K� M�*V����+�'iZ1���ÁB,�I�I� X����'c��2!���Ql��K\{BF��	�'���SGMM�T:���sA��	�'�4m`5@� /H��؅�^q�њ�'�\���E8]��b�E�$��'�F�,T��ضⓘ�������yrʞ=,A�m��"$�$1:���y�ɛ�v���	���+0����:�y'�`J\1n�|�Ӂ<�y
� �p�kC/^ƈ��A
n�y�f"O�)+�L�NIz!Cm��.� �:�"OP- �&
�L(@����~r�
F"O�T�e�	�A ���bQ"Op4)��2M%L�s�M*�5"O�U��C�F�n]��!��bE#"O��t�)��8��:]��a¤"O���D�C��4�m@="���u"O\�w Z/C�XHq��,Q��X*�"O����㈊
E� k��±[�"O�T�NL"HP��DG4��ؙP"O(�B�Ƣ'o�<�$Άq�>��w"Ox|ې�-.�U�WP�P�"a� "OpQ1ee�(V�z�X'��14o�iK�"Ovy�p&�\����[-8Xz�a&"OX�zw�G�}�H���ѸM� �Qt"OV�{S�8,�X�����k�"Op��+Gu�	���\�6�H�"O��R�K�=-[c �C�T�kc"OTG��z)���@�TM����"Ohq�6��:�>��T�^.>|��"O��X���	d�Iq�Z�KtP�"OL�X4��>��� �������"O�MR7L�q���I�%��"�8c�"OjE���S���4A��K��`�;�"OΨA�M�++c��s����r<["O�-�.� �<�"��61M�a�"O4�I��ū��~����gBU�!���
��4��W4d��e2�A1 �!�l=�hK���4ݸ�s"��\!�D_�X�@݃�\��4� ��}S!�Ɠ_��1B'N�cѨiVEa:!�d%'���@�$E�n�7!�� �125E�8O�03Aбq"!�DJ�T�`�£�58��}b��T!�� f� ���Aо��a�L�U�!�]1:w�Y�ʝ'���Z<#@!������#p�hsīМ~�B%�ȓh#RY����E�@�A)��M���ȓz�|
�B��u���b�ǔ5j4؇ȓ!H&��raL�)��īoT+����ȓv�ԣ����x@�Ed�X���ȓ,�V5§i�*�(�N*|¼��"l|�1�����b%��N����B��4�J�b$CCiE�B*��ʓP� Ca�uX��	[7��B�	�u�Ƹ t�C�C�
�0ͅ�<��B�ɭke&���	!P��2�)z�B�ɟ2���BIa��(&�@�\��B�I�<e��3AK��	�p|�&7�B��9P��5*��V���)��٦{;
C�	2ZVt���/��f�%S#��/E4C�Ɇ��,k�j\�X�A�pXȇ�Eb�@#-M%���Rw&�_^��PB�{F�������
�^=�ȓa����U�*^O�X���8l��؅ȓn�hA��BИ}����G��Q��C��}bӍ'��ː�ό#*F��^lX�Q���7h:�1�d�%�01�ȓt���w�E�ZY��XHF&l��9M����Ԛ.�Bx��  N�j���:o�ݒ �*Cʺ���MR�Z̅ȓcv�3� �V�EZ�dM*�X�ȓ7�,X w��CT�̙e�]�'�q��S�? ~9��#͡K��w	:'I�]�v"O>�bp"͠Ud�b7�^$C	Bذ"O�!�f�גCc��R"��ʝ`�"O�i�K^ 4�M��B�UZ�	ؤ"O6��BDN���'�Xg�T��"Om�ցX9�<��a=,���y"O��@���py��rV0��"O�Q�n�%ig��a��Z�"�I�"O�XҴ�>�p����.�4��7"O�[e�T�u��RL ��w�{�!�D�����Ew VPҁfP�Hq!�D�(u��i�#��@.��C�猟l!�2�,͙�S25Re���w!�$W/800�U��00an�1#��"MK!��E'\1�B��ˍYN�'{^B�	y����fCL@�0��	VE�C�I�l����qˉ�^jy��ŚCڶC�ɼ1��`8!�Aϒ���k��;�VB�I�2B�b��1���E�Q6 �B�	=1X;d�ÄWyȠ�3��B�I 
�p0Ů<4��R�J6b�C�	 K���r�_�er]��oM`c�C�Ɍz���3�oЊ��Z0�]-��C�i��?΀���	�?+�y�q
.D�x҂�K���٣�Ľ&BL1#l(D��.K$_�ra�c�`�9�%D�LqUG�,f�REO�*cX��Pa9D�$K5��:sy�ȱ���8A�H�+6D������CP��y�AU�b��Ѹ$�5D��F� ~��5�rō9^l���U�6D�zcĂ�0�&T� ˄_D����"D��xc���8�ȫ��C�s�ơʆ !D��2�d������l�jhp`�>D�X��K^�y�ݣS�Ƒ;�hh��`0D���CjG�O���a���ۜ��2D�0��� �`b��Ǿ9���s֎1D�x�p��/LKbJ[�`�l9�P�/D���Uq�ѣ���EvrlRE�#D���EBϑ1M"�§�W�tؚ3e�?D�����ܭo��@�SM�4�j�*D�X�6�!n����
�T��a�*D��s���.���Ԉ�m���r�(D��KH�G����&�7d����k'D�l�u
r<�A(�
�rBC%D�g`X7%�@��c�G?tK��
d1D�8¤�@� 6)��K2t���) �/D����   ��   T  >  �  �   w,  7  tB  =M  oW  ea  [m  �u  7|  ��  �  G�  ��  ϛ  �  U�  ��  ڴ  �  _�  ��  ��  (�  ��  W�  !�  ��  ��  ��  $ � � # i! �' �-  Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�� |d��"O
`�(�;���8���-0��1%"Oj4��ND^[��"3/9�0|H�"OB���H��*�ʞRy=a"O�味V�!X��!&F�:J�$���"O,��a
���C�Ą�M�"O,$3%o�-���p���+Ն�:1"O��ݢ1����`���y14]2��i�<�6��{_���c�H�`�fX�$Kn�<��A̼VI�xR[�)�Ć�pඤ�ȓA5��('nߡ4�� �)˩%� ���,��r�؊b#`T�eT09���ȓ!�b��g��}�8�F��-? �ȓ
K|m�ș�VṔ���2�%�ȓ"R�X�j�4JN�1�˘X�i����̹	_�jZ��1!g��zܶ��ȓgil,*�J�
j�Ne��i�J%b���f	�(U��:���G��$Y^م�~r�� S�%T"���k\�jx�ȓ|4�1�îJb��@ӵ�ݩn�V��/[`�"�v4�R�!ʎ<��M�ȓ`:��z�ؚh�J�Z��$HY:	��H��p�m�C1��!��B:��0��EnjZA V;9����J[
2���	��4'J�EA�IVW&��~�(aZ��ӹ�>� o�Y�|�ȓ�f�A�
Ο7�H��M�$�����mޠP����/���ANXo*�ȓTv�����{ ��-7�*h��I��sB�8�8���3����ȓNe*M�悡;������X�o��!�ȓ'lj�#F�m�+R&;�|��2)n�C��0S4���T:
b��|�O���;�'t�4,`v�K)�����Nk� ��+:�Zwd�gIv�:�OD��|\�ȓm�@ � Z�n��=�䢜5P^ȕ�>9������C�z!�1��ϫ>��!ҙ�y���pE����J;@<b�Q�A;�y,֕~�詑s�d�� ��'��y�i�6���.�	�I&�A.�Ң=�;�hO��T�W�{�h��/W\}z�6���'�q�"Y�3G-LJ��1��W�|�6()�"O�)23��5�ڄ�p.�3{��[��'����\���0�E�
���V?f%��}< ɓ�d:�r�$�)�8�r&b�'y*"��R�D/v���@^?z
	#� [XC�2m�D��#ޅLؐ��p鎹kR<$ϓ�~��퓟(�	�S�٧qFRC�� �V�IH������W�qJ���h\$]�p4L��'�a}�,�*�a���V��<�tM�<�p?��Osd ��9Dp4�5.�.{�zB��|�'�~�86l(1�,8��Ύk�(���'81O�u�|rL~Za�%�lm�_���/U?p��C�I�Cw�xY"*�GN�qJ�'���˓�hOQ>A�%'%�x�P�K$!{<�9B;D�Dz0l�^�j�4�ڵV^��DW$���"��?�HI�jݍY�����(%���f�<���L_��:p욫,�$�⋈6~�R��0?y��!`p�TZ�g�B"�h��{�<y ��,E�`b�㉙-}F512��k����'�:�Ѡ�6%j`�i��9U^hS�'OqOX��d��_9Xd"Q)��FǖiEL�;&�!�� \��q�W.fk��Z;2��(w"O�Y�t�X��"�!� ^�����'��V�!IG(��I?!�T���j)D��A�H�X���'fG&�.]�
"D���kI
T�v̒ab�K�6�#�O>扔	Z�L��LG-k��a���1X� ��V��h��`�ɡy�!2�N��pxXD0��'J�O t��AG*d}��9���<?�ɻ�"O$�4.Ư�^��^�,*@���'�qO�!sk�:J��qx�O Ud!��V�܇�	YRXjWA�*�\�m1g>`�<a˓�Bx��nH?ŀ�f�5WX�5���F?��	�<!:�Sbb�)y�� �o�[��B≊+�FQ2�R5h��b���4C�	�6�̡:��C/:n�����,cVC䉂iX ��@&U���v��;,(�0>��4%s�`�rB��� � �@!Q���ȓH�hp�A��uL`ȐFY���4��C�4a�"c�V��ٻDN:/�,�ȓ?|�i�E���д� �A�~;\8�<�����01��� N��u�
�
��˳O�qO�����L�O�ԭ@�{������rD���Ѵi�8��	#��lQ3�>o��A��(=XJ�<���;�$�.kpC�`#Y��H�yb�ʿ.���H�b�Hb���oA���+���>}�V̉�>NlJ�	æ����<D�Lr�H�=(��sI^JOHi�CF:��<y.�y*z9Hv������e�<qn��q��T��\)9<��F�L�b��"~�s��YS�C�� G����\	�2��)�����[6`�!@��,�X隷�.D��S��J4ν��`қT���`@���hO?���=3�`�����d��ȃE'�;�!�$U%!0в$��*� ��"$Cd�!�D�Yڮ$ȷNA��X���E�'9�zb�V=���{-�>W��i�6��zL!��],���3� 8��y�&o-�	�<YW��O4�S�4����S�N���&��@��CQ�<!�F�' fU�ll�(#�+*�@X[t��	t������G}� ��h k`��o�~��� �yR��2���`��C(`H��,���y��&	LY�B>�Y��k[��y��\Ψ��੄�{B��������ybJ�2B�p��I$xJE��O� �y����T����̡"��eK��/�y�!9�~�17 ��iv�A�M3Ǔ��'I�R�(M06�1c����%�y��Y6{C8��1-�0"I� 閧��'�ў����j!f�q��O[-	�c&"O Hj��۳Zdz�YQ�Wj� 9Q�O��:�oL��ˆ�&l�D� ��Mnp�Ey��Dܖ��)�]x���S�TS_��c$�ҋ%H�5�O��Q�&� i��1���9���4�IQ���PCΉ�C��Le:%��+a�!�$F�R�~��(~��5ԉ��#�fp�ɖdQ�"~�d@��0�9k���#
�		��4�y
çu�.���+� 3eJ�RE`��y�A��Du�92x`���͈��=1�y�`���a��Zy�b+��y�	�&z\l�r"_vT`8"b�B��hO,`D�4��:��=:��%�����y2!���sHM�t��D�PA2�M���)�禝I��8
v��	�4g��]F*(D�����M�:D}���/8Д���>��S�? �4p�H�We��ys/_�'S��Q�'�1O@���GE= `�:��'1JȕQU"O�	c�����@P�+E��|�>	��I�7o[�\�/ξ\�\5Ȳ��|'!�Ă�e�} M�8xje��d�7U<!�A5ʞp�R��i��t�3$
�9%!�d��s1�4�*nڎ�q��"��;'OxH1�U�蜸E��7)�qҰ�'���:	�!z��P7'�]�h�r(C��RJzУ6���E��2.� *C�ɢ5P��`E��*�9���&��"?���	�!�ѱ�eI|4@ic��Rl!�d��m�d��D��Fŉ����8Q�Ix���佸�T�!|<X���b���v&"���"|�'w���D@�c��};��� .|J>!�^s��aG�'��MQ׉�L��I�բ��Ď#��Jѩ�G0�{�f��!��\�We<��d菞5Q�lЀ��E�|��x�`۪`r��S�xT�qB�ڥ�yB�0��P"0�׹���g��y�D)*�t1S0�.y����#��1�S�O("x�E�1*�|�aQiַQ��01�'��u"��*�� �P��{�"ݡ�'��y�ꘓa�Hi�G yN����'ab!ıY�n�X�jN�j���W*_�p<��O<�'������-q���t�`Êy�����
���@��h9uBރV�E"��O��=E�"�I�h�'�Ȑ|���5hE�^V&l	J�8���]�˦j�uu�����p���OD%�=I��d����샵���"=���@@�	1!��I,DXG݂~!D�2N�Q�F�To��m�ܩS%�\���&O����x���7�X��uK��6vy��L	�K����>��'�2��i�'*Q.e˃=�P))d���!��*=I�cΒ���ȋ�!��Z*A\�@��Y�d���b�U�)�!�"8�Z���fK�N��|��&Ia�!��G$�|��O3�a�0慐\_!���#�؜	��g|@ydG��!�2$�x��a��K�]`g,�t !�
�)i&�Y�� �lB��".�3)�!�Dd$�����ζb@ܥWo�!a�!�$ɀl����-JR���5��r�!�,zԈ
Gܽ�*0퉏n�!����
�t���E�r���-�&�!�D:�l�f?P�HD��,2�!�$�	c~ ���I/
�D5hb	�n�!�Y��`L��o�9v4��D�D�h�!��@�XTR4KKd<�C�Ou!�dΚ��ġ�S#�ɨ�uu!�D�6,���0�[qCN97n!�ǝOR����Gä+�	���z����i�t�c�.���<1�P�ȓ��S��=_fq{4m;R2�i�����cD�_������.Za��]\p���l��3���s$�,:�V��A��h���[��[��߂0�j���Y��06dG�++��%�X�@ *���.�!f-�q��@�%:ir �ȓ=[�0��M�?_�p!Ʈ�2Fô�ȓ�<�Iw�A�d04��Y,/�X�ȓህ�Z�!�<C���%,걄�K�����K�$�ؑ�$T��l�ȓ��8���m��a	!B�8���S�? \E;Ǆ���k'��Ci�	W"O|e`�FJ�b�s�D��Sx2j�"O�lq��U��Y�c�b9fY��"O�(0r	66�����<&��5"O�(@� GN�� EI�4Z<|��'��'��'#b�'�b�'��'P6���Z�*Af�*��E�!�,��'�b�'���'J��'���'*B�'������G9��ؖ�����Q��'��'��'N�'�'���'JB��"�Y0T=�	��h�&Ղ����'$��'y�'?��'J�'���'8N`��C���)�$���dB��'"�'��'e��')r�'���'"Q�@f�9l�P!�� I�.1�U���'v��'��'�"�'�B�'��';�4��ͳ0�@$�3":P�A�'t"�'s��'���'�B�'���'�� ��O�Z�l3��:�5i"�',B�'wR�'[2�'���'A2�'o�`��dH(��p�"H�2ٴ��E�'�B�'��'"�'���'���'� �2�-�H&�I0@�
�]�2���'�"�'���'�2�'�R�'U��'( �
bv֨XJ�JK�Mb@���'��'�r�'���'���'h2�'|�z$��9���Hր TD�b�'��'�R�'���'�r�'
��'����±Z%�� $	T?f�	W�'_��'�2�'���'��"t�L���O:����D���$��D��9�<	��]zy��'��)�3?���iw u#T�2J�z��'�s�qag�)��������Q�i>�ɡ�Me8t
�y���G�J� ����'���'�^\`BH])�y�'�|cr#����#�O������+MP�i��$�%y��2��O�˓�h�Lmit&�k�4�&V��2�b!,�Ѧ��Ҫ0��i��:��w�
-�Gen����(T�P�x�P��p�(�m��<�O1��1�g���b�$���,?f�� I�OJ�!�18�3�
�\���=�'�?�!��,K�(�(�9 �틀N��<�*O�O�XmZ�FKLc���g�S1&���bA�Y������]�j��I��M�Ӻiv�d�>1KCU��b�i͗	�ͣ
�]~b��2(�Za��T��O�NI˗a��@U�� c%ʊ�+��;���hy�����dU�rd
}�Ơ�o>Ԙ�%��o��d�঵ s�-?96�i��O�i�3v*���!E
#hhp"�d��Ev�
٦�Cٴ�?�1���~�ؽ�'8��^ ���:���Nj�HF��[+ƩI�@�L��H��Ȕ�L�䞟^���_�~P����Ιw|�		DB�t���Ğ7���⁁��ze���7l\5�� ,5$t�X�'�9t������#���VM�l��. x]1!�*s��4�7oS*\�I(�$�M6�R�j� q��R�䞁\Q� x��Q-c����f��#t��hT&
�Q Fe�v��		��q0�#h� 穀	�а:ӧ�1�#fA�|�2x1���%Q����	5|*��`f��ӠP�r#�.�H�$�w�xA�@xB�Y(��ۧ~���B���M����?�����>�b(̤G�$�� <>\� z�˓�qDx�O9�-�.�C�����I�#a��>In)oZ�''����4�?���?I�'{t�'��`]��4��b%�(v�&�aG֎9R7�U���3�I����d�جi��!3B��8]t��L��M���$'d��O���
�4�~R��(ĉ�!�@(1�����ǌO�b�H�#�3��'�?1���?�嚋VM�]��F�U�s����"|���'��5��*��OZ�$:����iZ����%���I�2U�-z�U���`2�����	ǟ��'<�H�(��`��H�E�;2���̳CEDc��IY�	Dy����b}��,7ΌCRi�:�B�y"�'	r�'���'�`���'b��Ѫ�>��A��NFz����&o�R���O�=���O�DW�uz$
¼i��ˑD����1��Wfs}��'D��'�I36+�`�I|"�#-.�N�D�B�'<��W�v0���'��'���  �hb�`%��IpR�����lU63u�y�&��O����O���'
�|B.O��I�Q�p����I�&C=�@�&���	Ɵ�Q�M�1(Jc��fyۀ�ÀWV�K'F��}��n�`y��6��7�h���'��4F;?	E
�DsP�}�~i��nZ|y" ��O��~��c-W/@�e�eB�sNF�#ǹiX�(�5�')"^��S蟠��yyRy�4��B�R m^��*�>/��7�8c֨�W�������+5F��/W�������M���?I�:��BG�i���'�R�'�Zw� 5�87T�A�ə�K�@ѳ޴���ѽ01l�Zc9O�S�?����$��|e�Q#����1r�^��M��d�*	�V�i�2�'3��'�J�'�~R øbY*��O?�4�Y.ڔ���MC1��ԟh��Ο���\���/\�T`"�i��m����Њ&�>E��'e�8�d�O����Oڤ�Od�I�8r��֏�p�� x�ذ�@��H=������՟���۟�O�N�Er�|�C���b��jڞ,���$�ɦe��۟���䟔��yy2�'zAY�O��,�g��<g*��G����09� c�����O����O���O6<�b'S¦U�������蝗kd��#ƾ	��cS�Ԝ�M���?������O�Urr7��D��l��ۻd���A퀨��'���'>��'%р&�{�,���O��$�T}#���P �C>�QY�D
(�xo�ڟX�'&2�ɖ���|��M� �<�6���'<�|�PÍFp�5��i���'S�5J�dn���D�O����f���OH̀��0)��0B�G$b��!�
j}r�'�\IT�'U�\��Sq�	 
i~���*����CI4V��v��wr6��Ot���O����
���OZ�D݁'��i����r�z�1�U���0n�\&��I���D����'�!���n`d���׼q��i0�Gt����O���z�nZޟx�	ڟd���֝0`�ĴP�_����3��Z6��O�˓+s�%�S�T�'{��'��|�X�c���p7*�V�8&$hӂ��`�Hl�՟��	ҟ8����i��L���Ue<m�u�CX�����>��CF�<!���?��?������Џ#H�9��
D�YKE�\�&Z�Y,1\�6��O<���O:��I]�^�p�I7y�������<X& ���	ʂ���a~�,�����cW�Gן���ҟ��)[�``�ش8�93�Ȣr��u"���_�P��i���'���'��V���ɦz����Q��LY��[��b����݋`�9ش�?����?y��?���^]@��ֻi.��'X�ػh�,D�\MHǣ�35���/`���d�Oz�D�<���QΧ��:u�,�`o��-���4 �/(��6M�Ob���O�D߀��Tl�������!Ȟ,�Sk�-G��3,]�%b\[�4�?I*O������O���|n�4����'O$n� �I�F��9$�7�O�����N�ZmZٟ��	ޟD�S�?����g 8 ġR�ay�D��nP���OH�DL"W����O�dC��I!�4�8Ġ�+׊�$?J4�(���M�Td�����'��'<�4�O�2�'��N�q�����:����$Z�V�6��f��$�O���|bO~b�.���%$��̑��Z���dJt�i��'�j۠KqH6�O��d�O��$�O�

w����2�,X�X$?Û��'���=z�x������럸���O*�93�Ľ.������<j�X�ڇ
Z妑�I3Pn����O���?�+O������s�:�����hV6B�H��i��m:����yBZ�d�S����Iiy¡˚H��Eh��K�4c��(>��D��>�(O��<���?a�����pwF��7P�����|���3G���<�(O~��u��OB���O��D(	\nڻ3}���HR(0�V���!$�(�۴�?A���?���?!+O��D�F��7qwZ���+��#�0�v IaMBY}��'��'��'ݐ\��b�t�d�OH�H�$ �r%\`�$䌀�@X��\�����ϟ���wy�'��%`�O��O�Us��լy-���f��H4�2ҽiT2�'��'Q�fjm���d�O0��㟼�Y��7�jd�&m��*W��������ry��'zeɞO�ɧ��4r.L	r'
d����A���]�xYm��@���\�Tѣݴ�?y��?1�'����,��������.ia�F*7�P�Y�S�@�ɕoM���	j�i>����C�DP L9*��+"p�t��f�i�$�y�Dg�8��O��$��j���O<��O !AůJ)yv��BN�,M�����SԦ�b/�Ο�%��N�� (u��:4���{��QT�@!4�6�M���?��6��1�i�r�'��'2Zw�*�!��0���ha�����O�ʓ��Q��D�'pb�'mHT�!���A@Q��!Z'�a��$Q�&:�l��P������I#��i��$���*���C�P]��2��>��)��<�*O��D�O��$�O0���?Fb�@�A��iE�f��P	���$˦��ݟ���ȟdc��˓�?���9-�Q���8S��:�F�89:������ON���O���O��l&�}sZp�/?�,�A��F*x���@�e��d�O2���O��$�<���:��|����E$^�I#�F�w�D$+h�����OJ���O��O"X�:��f�|��Oҹ�猠+�qƚq\$D(2�֦�	�\�I{yr�'D�]r�O���Op4���7E��(���æXHˤ�i���'��&XˆpHL|������Y##g���4^�˅�T�8|�'h��
I��#<�O	�e��6\��L5GÃx�	��4��$B>@�)l4��i�Oj��@B~"��O��84a25v���N��MK*O<�s�)�S�z�XL	 ��J�Z�{�#d��6͐P}n�ퟀ�I������?��؊}Pc���&X����=W��Ȏ��O>q�	l��ݱ`��n��0���_�����ٴ�?q��?�qf͝==�'�'[�*t3Pl:]D�)�/(hM��}��@�ߘ'���'��nƖQ;�I��) iǼA�W�]�)��6-�Oxl���Aw�Ο���K�i��Y�.�,(���02ҙ��e�>a���R��?I��?��O���EY�+$)H�F��;�QjZ�v��c����m��Ey�O����Yr'�">Q�k�LZ�FzP�)�y"�'m�'v�;DIZ�O9��@72��قC��1dP2hɬO����O̓O�˓e��m�'7ą�n�� �T$+N$�O4��Or�Ġ<��D\�5�O��8��=G��P̴��e#�J���'g�'��I7dG�c���#É�B���Y�LK'28{��t�H���O�˓t����֔���'M�$���\�2�O	+ۖ�aS��( O��'� =Fx���3E�8'a�1PR�;b-�D�i��I�l��q�4���ҟ�����D��l;L`�fO�G���d�s��]�$	R!#�S�'5����@�&��)��ʄ+�,0l�<3�1��4�?���?��'B|�'r�G�tҶ�:F.�5
���� {R�7��r��"|��|[� ��`��l�x`G�ڐL��8:��i&��'���$@��O����O��
р�㗣ǅv���8Rń�f�,c���G�0��$����@���xOp���`^m! 0w��#�M���*e��땝xR�'�ҙ|ZcL�����0#lahFӟl\88٨Otq�����O�D�O��AHb�䦁�>�����E�R�CB�#(m�'�B�'p�'��0�p�cR@:i�abC'P���>���?�����Ǳl^h�ΧF�<�kri؃<3M*`c�b\�'���'C�'�Q�P���N��tY�S�P7��U�E��>���?�������s�&>!��K�-d��Ӳ�8� �G]�MC����p<�eT)�$���A$^W2Y�̈ݦ���ş8�'EX����4��O��iP)&$��s�	Y�%6�p�A�I�T��%����"|�0l�dȂ��%V0�6M3?A�J��M�T?��I�?��O��,�&�2�VoK*-�M:�i�ɜ<�*#<�~j�I�t�8�"�J 8��0�	ٟH���W���ٟ4���?�1�}�w��d+U� �P��c���w�6�T&-��"|"�{`�9���N���vE�.Sy��x��i�'�"�[g�b�H��Q?a3j�H~X�)��V�̨��Gv�E�F$�<����?Y�1w Mʄo�0]7�L���Ζc��J±i��h�n�c�8��M�i�����π%� a�`��/L���:���>Yt��Z��?Y��?�,Oi�P'-?��4چ�G=L��c{{���>��������ߎYB��Zbi��d&�D��F"��A�$�O����OD��ư�e0�H��ő*:u��
���#��x��'4�'T���x�5��e9��{|��ti�'�Q�'���'��X��1�A΀�ħiY(��v&�z0���F�m��	ᦸiV��'�Iwy�"P���Y��S�����e�J�ki0pc�-nӮ�$�OR˓;�(�������'C����Tޔ�I�S�̓&�A�(p6�<�*Or0{S�?��|nZ�T?��S(WU>���e	�'V7ͧ<����/k�&��~
������P�Ư�/ ��t*\�n��-�p'p���'>m�����Lk���$��r�KZ�m6��oZ�s8��ٴ�?���?i�� �'\�lH5�fiH'�ĐQ�p=J��6+j�7M���"|��k��#�ܒ�޽� ��8].)���i�"�'R$B��O$���O<�	$�L+�$��^�4yX`MO0)�c�H96M-�I�(�Iٟ���E�HBu��͙�BV��`��ʻ�MS��T�` 3c�x��')b�|Zc���VE[&P������İE�d���O��g���O*��O��bxds1���$J�"�v`�bb`�5s0�'��'��'�	�f�*l�0�L ���	�*�����/�ԟd�I� �'�����b>�(2c�`j3NC[���Č�>1���?�K>9/OB!��]�8��>[4(��̆t�t���>����?����,K;.�%>=8���(W�@7%�Vx�dC��M�����$]�Mo�O���ᖸ5�j!��͋�� Qиi\��'[剧j!�H|������/�R����άyR���ɒ�+|�'��Ɂ?�\#<�O�x2�)��m��k��Dv�f|0۴���L�P(2�o� ����O��)
{~��U�t�dX%n�B��3����Mc)O�d�C�)��R���Q5ί|��  5E�?4J�6��E�<�m���H��ҟ���5��'��Rv��	,�Z�z��r��Z�j�D�Y��)�'�?A`(�,�x��a��ӅImN���'���'��e�#�)��ß��]���!"�')D��R��$t��d�>	�KXz̓�?����?ab������w�*F'DxQ��#+֛&�'�F0#E�$�Iҟ�%�֘
p*��ф��(g�4D� o��`���U���<A���?������%QD���N�@��m��v�6u��A]P�	�l��r�Ily�&�	���`��@�v3&��c�Ƈ8{���yB�'a��'��49��LZ�OU�Y��b�W(� �S]�i^�Q�O���O��O�����''��*3@��yZ���R/K�@�F<H�O����O�ġ<Qs+U:W�O��� ��Z�AB���7��#����	v�:�D,�D�<�U��S}��H��	��阆�S�E���m������py��9d�8�ퟒ�&��=.��D�A�yp�<�qPt�CyR��O���#8��6�dF(@B�FU�P6-�<�e�	Z����~����⣚�@{򌘓�>h�q-�^r4�� ~Ӝ�ަ�Fx��Tl��^�ȴZ�IG�?�������M���?蛶�'�r�'��dk=��O����/B9���',Z�L<|(b&������%(�S�OWB�W�T��Ջ&,3wQ�0P�v\7m�O��D�Oڑ�%�Xk�	ԟ��Iy?9��G�0���x�j�Ao`Tjs�[g�S����<���?I��	�x�Q�ڝE�	j1��N��Y$�i3�BF�@O`���O����<��1Z��q�E�'*���&�;��'�Lx�y�'���'��	�� D�!i�"f�&��3�tac�bɳa��'3��'��\���	럨@W.ֈ=��1� i߬~��i	@̌��c�d�����ICy�Q+7�@�.-d<�`�c{�T��%#l:&��?����?�)O�d�O@!��\?�lO
������0�E`��[	�I�@���ؖ'�x�v`*�IٞD�
��`��ɷ��l��X��Qy��'�RAZ���Y����Ƣ&I�Z�M�.�@�y!�|� ���O��_M�I�M~���B� �$<��Q;Kt��Ϗ�r�'?�I.;�� �?�O��C!Kцj�P`+B%۸{� �4���^׺�o� ��I�O����}~�g��:Д�W0�����&�Mk,Oz08��]ܧi�����l]�p�v���]e�`l�5dي��ݴ�?y��?��'j��'w��DE:!aӦ�kAB-�r�G�T
6-�
�"|"��/�.PIa�Ð�I3��2!.��u�i=b�'e¦��5A�O����O��I�}�=3槃�a����/ɻ<&�b�l���.����0�Iϟ0p6�^3t'9 ��'|ytl���*�M[��Ri3��x��'ob�|Zc�V�c��-Y�}��ɩ4{�-x�4�? �n��?A���?1-O8b�f�w\��Z�eޮ��@1�(��"d�1$���	П'���IП��ǋ�*р5�6�M/`�6���c5DL�Iby"�'e��'���6GR�h*�O�"���KB&9�0`���(���O���O��O���O���;O�p��h٠qC�a�l��*'L`�n}��'���'��I����H|z6H�s� �rc�L9�dz6�J9��v�'�'5b�'�.��'��b��w��h�:�g`�zμm��	Gy���s����$���E��8D�b��nЄ�xU�KO����;%�>�?�O#b�8P&P�T@TJ����(���4���#~ Nl7��I�O���A�D�mbm�n�z}��{'nܳ�M{��?�@��?qN>�~�Ć́:Ȋ�qB	18�\�0��ܦ� dȘ��Mk���?Q����x��'k���ٳw��1�w�S�aQ��ȑ`Ӗ蛅��O�O>���(fTrͩr�	�]B���_�%vl��4�?���?�u�_�q�'�B�'���1��truD4R,\	A/��(��|"	(4P��F���O,�d�>izvH�g�E)vp8�LZ�x-*�nZϟ�J�����?�����۴��:K��8"'�7��)��/�O}b�!4��_������t�	~y�Ą<.B��"J�A���Ub�8N� 0aM4�D�O���8�d�O��Ĉ�Z�@ۡLK�V<����2w�l��8O�ʓ�?���?�*OH9���|b�H�(���V��LŮ}MHh%�(��Ο��'e��'(4�#��B鐱,SsfP	"� ��.ap�S���I��4��{y"A]F,�`,{��O�xd�@� R��p`�ɦ}�	˟�'���'�X-y̟�ɳb\�pY�?� x��̡`k6��Op���<���2Z[�O���OL�t�!I HR�͖�hIT��z� ��?A�������4��6�4h�c&�ѼH^�Ъ�C�0�M[(O�t����#��������'T2�0�#��3E�H c9*�ΐJܴ�?��16��*���� ��aST
y�uQ�'@t\o�Pc��;۴�?���?���d�';"M�I�'�ۻE�<�P�g�sV6�E�t��"|����&J�i�05��P��?6a��i��'�b/�K��)��S��Dѝjp�1���C�"lF��L�)��b��!#Z���'�?����~�I��	d$ �&���pUͶ�M�]�f= (O�-�Oʟ�$��%��˦�Z�<T� ��M��\�'z��NU�����Ov���<i���(@@2G��mt�I��V�|��!�����OH�d�O�s���' Δ�0�].��d��d�x��&�/#�"	�O�	�!B4b1���Qˏ|����2��C<ϧq��C�.�	*��$�*0���ȓ5��y�c��3���T��'"�8��=�Ԫӑd���V�
���h�O�p�M�V �`��A�Q�G�J����O�*�~EҀ(J��0���P
�bM���sïD�-��e;G���FF�ÿc���Q�	:xv� �CFP�"I����$�`tÁȵ4~>ʲ ��T�C苫%)h��p��A�혲.�:�@T3B�'�T�ƈԩ:��yS�i�W�d����'�"(W/��p䊚�:�~��U�X�:������2�]��l�X�h�#/���Ox=�"6)�pIcB��Y{�xく%��!É���TEu|�iI��� }/�ؒ�M��@�\��ۦ�Y��i��2E����m�])��S�I���24��"Kɐ4@ �$�WM�ļj�!OxYFzB ˉ6�����>PP��g�S�A�7-�O�$�O`�+���T2���O`��Oܭ;Eef�*��ܹ6��ʑgP$�Hx"7`�<2"�شvP�,*$�_�1�R��O�%�"��:kr �6!�?,�����+=��%�o����6D�;n�d�B�"0����8N��ͻu�D!ݶ6Wބr,U;lR*�(����䘪v��O�ў��6�P�[�8��bH�g�!s�b%D�Ls8ƣ�Y�\�C�����]l�����'��X�p������Y��C�*A+�y0�% [r����ٟ\��ß �]wu��'��0}��yb��F�1����SN�!V���j�az"��X�? PZ�"P1oeйj'>V�V (F�H&G,%�f����9J��VQ��['+YeqO�i�wsh�! cZ�	�x��w��$�������?���q2�����qӑLLO�<�aFX'e��|����6�� �gMH�i9��^y2��Z�p6��O<��6%�bI`#K�Ȑ��@Dۃ4���$�O� S��O����O`	0M�!�z8�@F� ��Z�O��`�f��'�H2y�P���Y�{q0��䄣dLQR�%	�0X��NN�E�J,3�E�F鮸1diS�=n�l�+/4�A���ΑCO>�T]����M�.��(�M�27���Ck�4:<��(O��$/��؟�����\��6F"ҕA�
�exXX�'N4KB�	��M��p��R&b�+<R�Pi�;U��6V���O��M[��?a,�B=R6n�O�iC�	N��<�[�n`:$�6(�O��ɗj�b)�d�;~�(�p�"�П�'���C"2.��ؓ��!>��ų���6��kvA��0QM0�A�����H�4���U���󆂧����>��͟��	N�O	r���hdҐc�)93�\h��I_��yb�\�BMz��1ψz��E��0<���	��L �UH��"�A�b�<��Bش�?���?�sE3>ݐ�(���?����?�;l&pR`��l�� �ѮU	L�T�z���<<���+fV�qÂ�%�3�D�� �|Exq'�4�z��a�H!)�$���Y]y�J��@�}&�VäB=X�b�.2�$aI��ӌ.tb7��˦����IYRL�)�<��
�$yxf��L0\Y#�Ղ*�.�@	�'��̩- &&��p�,��T��z�O��Fz�[>��'�Լ�5��%�$�3�f.t�t��-Q+�8B�'C�'���s�!��ӟ ͧNÖ%s�L	iDJ$9�́�*�X�5kL)}��d����=Y��M�0���e�
�}���R�O��n���X�ܣ��M"n������O,@rGc,�4@�)M�N��Vf�, ���'T�'�b�'J�OҲg F=@��$��E��5�g�'y�'l�̺rg��BZ�Bҧ��ZFh
�y"Hs�
�Ī<I�$_O����']����`=*�^�_^��v�od��'�2A�'�B0��KD�; u�a��i�>D��;zb���S<S��q8�����+u ���MM}�/��x2�M�v�ʽ7�F9��+�+�p<v��ԟ@
M<�A�ƚEeR���)t��I���e�<qb��0g!\0����/�l�
0�E�'ў�S��?��e@#6ݺ�ۑ��(T�c��s�<k�$�۴�?�����)�F��$C,�&�b�+ԻL��9A0B\(�d�O`�O��>�(�a�^}[>��O,�����UUOtݚ�h��b���KO���FnV��Ȭfs���ME6o��Q!M?I $��_�d�y�?�ti���'}�&���?1�iTf7��O��?��&\��u1UMͨ]}#K$�Iퟠ�	j���D��%X�KY�[-B��ejѣT�zt��	��M�7�i��'�=I� _�XM�xk�jO/l�*�"&CZ�D��'�b�N3[�l�!T�'���'v�bz݉s H�[�9���];��p�b ǥU �Fᐓ:; q���u���|���>����/�
�[5/=��1D�ۗG
��� "g�0J�N�{?�M�Ɓш��S!�M[��f����jW?	RZx�$
�U��9��lĸ�M+�i��$U�{���,OH�D�(t������̺o@�أ�Lͬ	6B��!Hx��o�*�(�a�K���՟|��$�7h�X�İ<y�)� ���zʓ;\���s
�+4t����N��?)��?��.���O�Di>��!� ����J
�@ �@j�@�k�+ @���Nkb^�;C&��8��c�=z���cgAY!@�pl!�'����Q���i�-I�x��]�/E��?鷿i�7m�O���?ى���B�\Q
$�SuQr�3��/�yB�"ξ�a/D(f�^�dj[��'U������D<κD���?)�J�"ͳ$ �XN�k$� 9��ap��?�Ģ;�?����T�{,p03�! �6�I�+߼*��:ƊV�!=Z���O��<r���G�YŶ}Ey"�֌=�	�p	Ԇ<�@c��6@�Z���#LD�@�1���QW��hȂvVLq������'QLQ��#щ'��P�Ӧ�Z��q$ㆷ+�F���'�t����2
̠�s��A�[I�u�
�'g�6-�'%���I�/cM�4iV��|Jp�O�!�TԦ��I�O H:2�'�"����!f.�(B��QoR�b �'_bZ�0���٣ ��uC�O�[�Ċ�'q���R��.��Q.��&jF�q��	L[�����J�O��L�Ò�^yHܒ5�T<�ЃI���%��ON$��?�xU���nX<��B��s��8�!$D�<���J"EϞɦ�(I֤<�E�5O��Ez"	'C�j!J`
E	\�9���*��7��O~���OV=y��s�N�d�O��d�O�n�(NF��#FJ�[�P�H��ٯL$��CwBU�Q��Ų�.��p?@Y�7D.�����M�ԎY�J\��0ǂ�!,f�L�c�T�J�~58���g1�+˄�?1/�VmZ=�� !!��P�s��]:D	�M�J�"E�UҦ���4�?��H9�?�}�'�bF �#R^9��ΜF ��I&֭N��	4i�J1Θ�M'���Db�80�D�Or�Dz��OL�[��Rs,Щs$&A*>-�(#���ri����t�������.�u�'�8��ă��ü"3�Y���U w�%�%;U�*�e�-nz��[t�]��p<�юA�hZ�mcs!�����-��EG���-7=���%�P����
t<h�g�P-'�>d�#FȉB$j(@��'�*7� C�'	�Ov)����b�����O�)i�Qzt"O�psc�[�U\J����6IgDQ�c�d\ɦ���FyR�J1@�H6��O2�$ˆ=R`jW�u�Ir旁2��$�O�9�g�Od�dl>%��䑞T�ء�]}�n'q�`�c	[��3�#�p<I�.�>V`��0�����'/*��D���"�B5v�L�Ǔt�u�	��@�'߈�X5F4>~��
�	L�i?`%�'�r�'��O>mC�A)��jDm_*i
�Q`"�&����4#E�=S���'4��F�K4f�Y���k�|�mПX�	T�D�D�K�U�L�Z8�RDμt�D|�U߬	���'Tb|2�,ɷH�<M�r�Yx��8{Aã~".�LjR�'>��\@t�D��N�"��>��OD5z0�&�|MXY�����O	���ɰ8�N`y����u��EKJ������O@�D�\��k�S���eJ�?J��R!ɐ[U*��?������'o��"8@������)j5h�Ó'��x��OR�a%�X/x�|$�%�P%$�RIZA�ݦ1��ӟ��	�H��c���$����p�i�	)��ŕMN��R	d��"şfXH�7G�1+��Q��&*rf�|�>�'"��#�Νe6�e�����y�#�B� R8�i�jQ2i�?1Q�S�M�-v��z��=$L�mسC�1�EZ�+k�f�<ٰ ���>�$�OB�D�I�~eif*� ���	��A�r��C�Ʌi����#j��^DA TA�f�2�	��D���"���<ɲ�^>">� �"�X�İ��+�9]��B6����?9��?Q�#�.�O��y>M��ת"��҂N� b�pH�ű־C�	�v��q�&��R��Q���L�B�z����3��y�F�d�(�RK�N\���D�S(XW����O����O0˓��󄙾`�2�m�/B�PRg!�>H!��Ē@�ڙ��I�������V]1O�8�'��I�6HV�y޴�?)�A�x�c�,
<XSt,��.�s�,�{��?!"!�1�?Q������D&fH���j]�B��		K>ذ�AJ�5s*=9�lҩU���䐛�>X��ƌ/Ȫ�(�-G
ݫB� �3�c� =;�u���)u����Od˓K"����yx�-c6.@2a�|-��?������&�0�̬�~����0k��{�O�%o�r;"ͳ�i�Q�DP`������Iry�
x<6�Ot�$�|B6�S��?�Ul�!�2k!��U�X��?��.]�����D�a��Z�ʧ���&�t4چ�؉D!�ՠ��e�5d�k��I���l�����-xs(Lk�lؐ}��1`���-c�� ��a���M�U�i2�i C��;'�̮c�B�Y����d�O��D�5�4���͜ Ѷ)��E��d7آ=ͧN2���2��	S �����5ю �|�F���O��X0�X!"L�O����O������I���#Ą��E�4Y 0(�MU���!V� B��q�g�	"N"��BW���	iǅπf����x����S��}&��iB��/1���XǢ��6#����T��M;�i12��C��,O����23�rESf��?4�v����a��C�I-hS��r�A��3���HJR��z�����O��I3,��M�&�Mvl�as�	jN|L*p�Ԕ�T��Ο�����<ڮ�n��h>Yy�l�#��*� ^!U#��T�Ӳ<��1��Kh�36 X�~������o.�X5啊J)��y�©t�J��ЂEPB��bP�u��K�ɚ�\�-�G���'���� =5� a�w��8�%J���?����?�����D�O"��j&��"�2=�UP���` D�hb��Gg�bkG]�2:�t{�o<�	'�M�����@� m�O�B�[�(̮Q���9>3��Ts$��'�����':B4�$�����/t���[�A6h�CN���7I�,:_`����M� �F~b�Ȧu�Q�a큟}ꑐT枘$�t	�t��c���`��ua�H�Oרtd<,�E*QQܓ1�]�	��M#W�<zU�!-��qM�1&�X��&�"��r���s�@�2���F@ԜhfDPXd� �8�ݴ h�i
�"	6��L�$�Q�<�?����9O��k�h�#T	A
��+&\`)�"O��`��+�4��X
?X$1��"OT\3ƯIZ��* $)�� "O� t��3)_�9Vm��l�)>���@"O�l�hDV�5�2�;X*xER�"O�}���t�څB���.O�����"O�$�ÍN�;�*���
�|u��v"O�}X!G�!6�8��;PBt���"O��he%��p:vt����#Q�ѳ"O����ϥ^��M �YWf�"O��ы�{��T�$�[�%F��"O��ɀ�=x\�	b"U���� "O�Ժ�KO-������L0!"OT�6�E<ie��c��V�pې`�"O|�*�Ǩ\���I��R?%����"O��X��ߦ$V � �>I��|�"Ot�+ BH�oZ�{�g�wæ	��"O`�P�"I~p�hb�$$�21��"O��T�Q�\�����!����"Op�E�Ϫ�2I��Y�3A�A#�"OT4YÄ��a��%4A���"O�ܸP��-�ȑZ�OV,-����"O`)�/�.C��=P$���_�Z�h�"O� +4�7I��HIïW�֝A�"O����ϊ�V�`��c�,u����"Oά2a!����X��Үi�	� "O5��і/���Zbc�G>���2"O6P�-ڶq� ��Ed/r)ӕ"OR�Q�H�a�n����ˍ9�E��"O��#�J[��b��Eƕ53���B"O�0�
�y9���� a�P+$"O0�j��@��`s%��Z��s�S��* �7�b��1G���S��	Ɵ�aq�޹|��m�3�� ~�A�׫5?�Boq���p�Gv���9��V�'f��JBmZ0
}�	Z碑-MS��(e�;i�p����?	Ӧ)
E��Pr�
ؿ���`-�-��R�'(��Ey��_T��d%s��q�L�1q�5&�����ʶ�2�8I"k3 �^DX#��1#4qG	P*e��O�P �BI�ML�Qyi��:Fp��d�x�[MXxbPf�6J�N"!��6��'玑�GS������-��9BN�-��!8g�G#M�  ���Y�̅k��W�~5�0i�`!�Q�L�fq*�F~򯉖9_�H�r�Y�m	s(/9������T}�`[�Yx�3�oE�O��u�Ĥ�,��'Q�m�&Ժ��$)2h��E�ر��-�mCV�[ud�����H�@�E�@a��2�&�Bs���.d
P�
� m��#=�;F��� ��cޕ�a!LƂ�Z�i�2ʜk�Ǿ�`s�(ݠh����TCy��Tn�����T�_3��e
 S�g>X�i�}��/�ڹ`�B�?M`���!H ��B=� �DD�+:$�Y{��"�W��$:B9|e1 ޟ���fM߰`	���#�!0z��k���#eMT�Z�ҝ��W�c8vP�'PVD��! ͹�z"=�ק�#8s8� 7`��>��&K�Cn��$�.VKVlS�{�d�cp���ـE��b٪m�*|���dM#z��TŁO#4e��(�/ ���Gy"bU-L�����kk�e��?��-��K���\+6��!�/��z-�D	!�7�2�e����#�'���y�����RC��<�iC�ë�?��놻}��0��Z�d��{����"\��5,�&�eɗp�:��AB���`R�芘F���4�O�e��L%�pQ`��+xj�B�+AI�b��uAf���+t��P 8Re��5|�\�����@@��(����@�ܡ���WQ 1k��ӎZ"pѹ���-�z�!
�6�:�!
}�'"���@��	��1�FJ��"�"f$ک3�6��G%$�x�/�	"Ƣ�8�aS�Hap9rPJR�w|"⟘�E%-l|�ɱfc�!dI0�r�˙	��81��S<~�hh����c�`�O����3��E"��36Q��� )O��m2�K`�Q����:s�6P��wL�xb�B�	��YQǇ7o�=��l�t���75=�X�dգ����y`A	�y��ej1�A9��������'st�A"d	��@���ܟ�N<p܀�.1���	m�@�5��  7��� Hʒ��-������?1HB�T��l���=0�D�H
�P��P���i��"2JQ~��
�Y-5�Db�e�7@������M�Ch����x�\#LJ����Ň}��PQu.�P�H5��4b��1j*΄��&X�MEx��ԲP{ļ3��@�R�p�Xe��>*H,	1O�9'�4ku	G����ɂ0�D�2��H�r��iޙ�-���z-V��:�"!ƉmӠ�qp+@��p<��L�DX��v�AN�5��3�E�ӄth�'� ��C���dǑ_dd|У�>�MC�hj�q�C@%e�r�!І?e��=rA 3�B��#��<�����E������c% F+;�ʠ���ԛ�6��'���CՉŹ[��$<,Ŗ'g^m��!O�@����V���)n�
(���k��q�����D�5D�0�GN	LW�e����~If��  �P���O^dyau��:e6�"�O4|�&�Ky"L����G{��ƙ"gz��)`<d5�2�B
�n�+�.ТuιB�CF�lS*���s��<ͻ�¨�D���@�f���iR�\�IlZ8uht��'r�x$E��X� �ǂo�Ճх�p�pQ3GÕ�O���N}�ͽ>Y��R�>���␎,jfh�̻#]tH�saχ�L��L��`b�Dzkֱn����'A�hT]�]Ϫ�Ҧk�����S4�������v�M������s\�H�5�� �z�[��p{&I�O�)h�ٴy���#D�f�X���'��LY����8B�E-�䈘x�D�c*OJ$��D�8p��)��z�pqq��F��C#D�Oذ�2��IS���E�6/�5��&��֤��^5j���ai��Y!-�*Q�,OP,0�� b��i�i+pa��H5�����8���#��&�O�@V���[Z
]Z�bJ�)�x:��F������鈄�?٬Oe�Te�JO��IRW�닏�<���QR.Z$��UXu"ϸB���S@?Y����L�^�����4?��+ai>h�6k�8�6�����8;'�D�>�/�	/���BH�OZ��X3�׏	q"���߫&.�*qe�^�H��9g�����P�R� ��D�A�Z�1tnX+��O��V�`��W�N�7k�u��e�K�hPp��ym�z��H7������%GXp����_��(O聡`�Q�^tK�ņ8o�N=�V�p�L�t�'�NTDŇ:�ħH�A�	�"pV(��$,����
4!�+o5���@�6�����%h"ZD���-p6nБ� ��PD{����/G(����T�X���*�ƅ���iz�J&�P���!ω61z�CQn�+�X�'��X �S����-��-�Ҩ(OL�,��b�)7zzM����65�� �T��"F}�E�C�k�J��C�d��Ib�M�z�X����!8�d�C���D�����y�hl"c-��ol��1 �<�剕־�+bcԠlrHi��M�Zȣ<i��VS�E�4�U�BV����e�Ojt'����m6�Ӽ�DH�$V�M*@�����U�lȑ�CfMɄB$�>Y�%O5pL���;L2���õu��Hȵ�� �h��,#�~0]%�h�;8P�PC(F0X�3�,�0<HEx"��'i�<����n?1�$�P~e�PV�x)s	W�R�X=� j�����%�' ����'?X<�b�!��(1�K:*��%bD�U<D��S�c��!ĩ���F�o���O��%�ם��Dԛs��"�i?L���E�;��	�d00˓7� �xw��HO괊�?2��m��$ġSr3$�$ԁ\�r1 �^�X��!���ګ)|}�r,�XN1�s�($��|�`�)@"����i�V!!���f�z0��V#F����a2"HQ����&d�zC�n�Aے����R4|I �{�*,7��@��֠o�$#��O �y���lه(ԄDu{tJ�@��s��4}���J�I�I	���#?���q��Ķ=B�B�j��
}�(jf�� Ѽ�q�D-i�ԯ��&���׬s��'���J��A0��
�t��f�HGv�↰<ѱC�{?)��s�FԁV	%�G�B���Ȏ_"dR��ک~�|�s@%DI�ɉ>|�>ͻr�����̗<�4�ĩ�,9S�+#�n@�}��F3�j̐7�ؼ���|�sW͇�]N���џ�'64�2��G�~���ط��M��. �
Fl�D��2<����6��bԘ��M \���(�
v�x9�'�T=�1�IZ��i'�L�N��H��'�0�su
�b8Ź���aLn\��FœX��*���z�.�NJz�d�Q�J`�)t	ف'j 렬�>��'��I�J:uI@�O7kI��˲iW	f�C �R� ,�t����lv��dn�D�*T��^W�'8��Pi`�4�����,(��π��'��	d��2��ޱ4P�t�a�,����Ȉ:N��I�_'.�6Aˎ�D������1︡��F�'�dt�C)I�C�(ae�'��	NA
=��@��"|���-v�8����53ذp�G�
@-*���U�PpR#L_+�`�4H�U �	�.����� �pG?^5��'���y�h�H��G48)@!/ПD���C�F�4�5x���;���
�!D?�� ʒ-լ*����"�� �Be�w"�lYR̨��$�>a�ӚoGJ5�A&�3�V�*s-A�9� ����UY�=�aՈrW��¸+�ZGzBꅮ1�N5��E���IB�ڻ$^�W�D�Y���c复�a䮼�'vU�#�����4�0��G��򔄒���F^.,s&�'�.-q":Oz�wďO��sV��8���F�����X?�[0V�����"0N�i�:+��n-Y�,��JP#E���S/�6�������4�剣6����O�(P��ghĉI���G��8�+�@}"F\�v&R���\i)K�	�Syb@2#Tr��ɬ+x�s���$����&>^<6m<.2�/O6���i�uy���"c7��')n�[&ND�D�B�ȴ��q��'��$J�<�p+խ1KĢ=����%���j��N�jpP­K�K�h�YR����I��O�./����B�'4�V�CР8l���2�R)��	�F���b�'�d@�"c��v���X5F�E��ET}2Fȉ'����`�<i�o�Q��ݠ>�V��w���Ix�)��(�B�f�<A�CI'p㰺inj�а��@bƙ ̎��^h��Oč1�}yR뗦E�x�/�м�6��Oz
�KG�a�V`�f��jy�&�iap�6��JyRÃY���!+�O1K���a}"��8l��%W�0��2�A7/�Z��4�O�;�@�iy�a�-��D{
� ���%)0V\��U+@5�D`�/�!!��Tٟ$R��X$���|��y�j�2R�P�д.T<�$�YA�E�M[B�
�]�"?Q�A�UX�bn��h��G��=��
�j,-��D��ɾR���$�$��4����b߸(!,RD�ܴdpX��$$Y��qX���=c�����2S�'G��&��;�ܤ���ՑE�t�a�Oи�?)4�'��)jql���b芐W��!r���J�7Ȑ�i¼C"�>\��°�`@Z�t�Q�4�'Z2�������5���C9O7�zH�\i��ϧ2n�Q�H[�2p P��%�I�d���4�|���X��=Π�K��*�Sz�*O*)�)�f/T�;�L �P�'-�v�2+vB亏��O[L�@ټ�׉U:@H�u.��G�f|۶џ�F{��)��S�8i�F.�!!z.U�E�Þ)�K�}�o��:D���
�l��Pi����:uC�@�2>:���#��N�
�'KQ�$���ߧ�0�
�×9T��Ѕ��d��ԉT득7��|�Um����H��]�5>�{W��'U6�DyR�����!Yj�|F+ÿS����p5}�F�?'d8����_���# Cݲ��' ��ڰ�
UX���&&"��b
<��hO�靹VVtXz�`0���2H�}|ޘiaM��'�Ʊ��0��?��6X�=��nP4G�ְ�qF�@d�t�%�X���$�& ұ���ױ@<��V&�Tx0��}��5^��J�7Gz� .K��ē���h��>�}K��'D9�Ї�	�I"����%�;8�ZFg�-` [?�8���ڞc�n�9��F���Ϡp4|��[䎬s�S��LR���,h��`�@����'��9�CɈ�x��(Pg�	���!��$�jeI0�HJ�BH�$e�1 ����T�"��]�Pؤ�	:7��c$�OZ"��YL(mP��{���!d1���#f�Hx$�O�2FX��Ɗѷ�
B�	� �� E�T�^�s���8	���S�$^"r��US 1t�PpyE�վcX�'��Y���Cz�څbgG�j��d��O��@i��=UǨ��AJ!�����2�$����U�)��XS��[�~�,!q4DRl�\d�6 ��<�W]&XF�q�%#ʒKZ��Q�^v�DV�e�)!���,t��� �.:�OB�	V��'?ڙ��垞_��)�,�|ܓoo�iZwA�#~��h�C�8H��B�c�� �8�@�4���.5;�����E��y7�[�:�<9��##6VE+��#�t�w�޳c��V��C�ø�M�'RK<�K�O�q�~�"�Ԅa��q�,�q$&�w ��:�^QppE�ȓ+�R
q�A�y��x�����E~�����7o0.�ՠ4�ܕo�h�'W��P �	{v� TG�-e�ΙP�'�V��G�$�"h�  Ć���*�'Ò	��8S*�����!j�'��&���UVj�r`�����lr���6�	*�XZ��7�����AQ i�'*�]�����F2��ȓ���cvf*�0�	DoW$���(	�(�-��J�P����B��ȓ8��Qe���g��A$G/ �ȓjG���QG�����捗!���3�="A�ͫS�:I�򌝷D�T��B�IƠ
�q���G� �Y4r��ȓ6�)D���	��+d ��	6���ȓ@t���Ŏ<d	���Z
�U��;�faK��9`�0�Q`��7U� ��g����s��$��1�� �$}�ȓ�40����˼�se�'I�B��ȓ��E���˜rA\9J��;~�D��D� �!�ڈ�:R���!8�h�ȓ$�pi�OG�+er�Y�K��G%�T�ȓL~�"�퟈
�4����_�,i���I��}�0�_o��y��˼\����4M�5��9��@����+�bM��h'8���$��`5�R'< ����8�c�LH�GM<���j��o��Ȇȓ�d��ƕ30$̀u�$O_�ȓ#�Ф@f��u���@�ͼJ(�ȅȓ ���I�G�B����i�;Z<\t��Q;�M�3�S�w��ӯ� "Wn ��S�? :� W� (���/�	���Y�"O�2�׾g�|�p��L㬕�"O@б+�!��d`V/��U�D(�1"O\P 3
��7S�[�j�YY "O=�G��D��u��Bo꙱�"O�*�G׳E�p�F�6���1"O�#��T5D������Od�ti�"O:,*v�Zc�x�Z�#W�-�V�{U"O�Lzb�6c	ly��AK���H�2"Oj���CJ�JzrB�'�`�"v �G�<dV�2>��FOT#��`R�A@�<��*�!�ڄ�Q�fxJ�*a�U~�<�����3 (EB KN�T�p�<I�hܶ\<0����j洡��R�<�*Ch�L����r��%
E�b�<I�N��4���Z�`�A�`�<����&�T�sqeщw�����B�<�@����iЗ!��`�ʱp3e�~�<�QBq3j���!�B�L\ �(�P�<Y�a�;N#�s+	���q��u�<����6�x�C P�+pio�<�A"�f���R6�N5&�-ʄ�n�<)���^��!�fN5֖A����k�<!��O/<Ѻ��S�z�څ�Cc�^�<q��?eN�r�Ꝼ�a�g�W�<皃[x`śD$��juR8Ч�U�<1� �$:�caޓ)oB���o�l�<�Ѫ�5z�����g,��ps��O�<9�⛛GV�遥@PVk�mWa�<��d�M/J
f�ݺ):d���ȗx�<��O3(�Hj���}�J��f�	t�<�7�ȭE�
���憍dN����$�q�<i���:�6E�W�C�wt����'B�<a��X�rv��P�Iݚ@aVL#`��~�<���'^�8)'�W,W�H��c�I{�<���R�E^(��e��!�����m�<��j�e�Tp��CK���e�c�<�ߢT�8����ۓvl�0��_�<�j���u�f�x�XD�0Jݟ�1�)ڧ.���z���!�0��TM��9E,��oo�I��W�4>(]`(�$�=��V�`R���JԪ�90D^"�|��ȓL����L�a5D+c�[�^�B��ȓAu
%ё���+�(ɚ���3]i��p� ,���AX�A�qv 	��$2��w�H^9D}���BAUͅ�T/VA��<j�~@���lr̩��*� �-�$|P�t�%�f�d1��&T�� ͼoF�ȗ՜B��A�ȓ1f1`�׍E����/�k���0u�=B� 4�t�k�B�^��P��`�Ƙ	Ԫ��G,4,*ƢO�v@�ȓ(/�!�0��Db>�1@�

nH��?�
�	QP�� (�(4ɮ5r+�f��ȓu�(1bw� CM�}��I�Fb:���S����
�*�x-:5���
M��	�������,�8с�U3�ąȓb�L��ë�,��ȶ�җ_rI�ȓ3�,�%N��Cu�}PR�V	Jjm��m�*���$��zY�5�UT����ȓ
~ �Q��>ew����A�$��@�ȓu^�]�ض��E�&��({�<�񠌅Kv�;F�?�����^�<������̅0�kɹ* i�a[�<�  Q�#�Da�F�#D�<cG\Y`"OV�s��-:���KL;.g��"O8����߁Vw�M8Š�l��y`E"O� ȤNޮ�q஍�%��I�7"OL����X	�Ջd<S��x@4"OBAkbEI�s`�QYR�A�Zy��"O8D���)e��6c�v�p"O�����p�
���S�X���t"Ob�`�dE.1^���g]M��R�"O� ��/T�~~>����<E��"OYt���:P��Xg^'5� ��s"OV�{�j=<�� �E�cqȰ��"Oz@���N�ʁZde�Lo�]yc"O|0�+�-��@�dS0�x��B"O�@Ō�2I(|D[5
��0�hh�7"O��hӧ�j��J�\�����"O^2������S��?�^��"O����G�>,���ˈ�T���"O���@�Ӗ#���3țf�fCP"O��� w�Ή�!B�+)���!"O�`��H�t_���	�Z���F"O�a�Ŋ�l5�Nǡu�fa��"O�U��F�GjX`]0��e�2�'G�(�d�����W�\�{�|(H H��^!���$tl`��L>�� �%V�k!��C�M��P0�� �T�e/��+!�D�6��y#����u(�L����Q�!�D�fm�Q�ޝM���q�/�2x�!��ҰS��=�0C��X������-!����i��1�>��W�ø4!�[�.�4ڒܹ�H����a�!��	'6�f�Q��z���fU�!��	}���nX�"�h�PƘ�]!�dڠnXp)���G�l����+2G!�$�/n�6�R�b�|���C��A@!� `h<�0�m�#V��<�"�@[��L����X�M޾q�T|9[�>%!�����y"���Fr��h΋O�N��#�D�NB��3=�d
�̆�*�3e�?%���$	H�2+�Y� ��Tْ�AB�ۂ?�F�m�c}r�$<�I�8��ّ\�%�� �� �������ox�q*�KX���d��y��r�� 9Zp
���,��Y�ȓ!�.��OR�D��#��Ѭ|&�̇ȓ4��Qs��&T�6y��%�)`�,�ȓm�R$���&|���Fj�(H�Ā�ȓ_��+6!����V w䤆ȓ��Ԃ&b�(Aƀ�t�Çv"r���z�n��1o�����J�C(l�ȓ�h���0R�b U>����	K�6W��B, ��>���]�d�.|E}���/��بT��2i�~th@.�19�B�3	+�ش\�<%:�`�A��m�
�'|B���F�-���*��� ;�!
�'! �#�Nؽ��љc�4';��A	�'�n�1��K>N���k�(n���	�'X¡1f�P�M�b���x�����'�&�u�LrI,�p/ys4eX�'�Ԑ������b�qM����':p�Re��k�j$�O�bt:$��'ْu���qئ`A%�9ll�D�޴�hO?7�^1. �RV�Og�f����(O�!��W�f�5+ÁZ�#��h-
�[�!��V+D�e�@�9Y��tAu�M�i!!�� r��*�5ra��MC6R�T��@"O���+Z��V�r��ߡ�� u"O�z�H��Ij(���aX�ݰ8sW"O�23�;3�ޜ+��J��6Y23Oj����6zbܐ����=��(�r+Q1�~�U�L��ޅNDܼ�TIʹ&E@�ۆ�&D�@
��O�S�0��D�A\.�zV"&D����_��=�Pȇ9^q���?D�������İ�#����F(2ړ�0<�P���6�x�Q�&*��-k��Ax�<��a�,0ïM�Bd(�(P�<�*C�5.IXc�T�'kژ��mWM�<��\9����2.E;0���&�<	Q�يt4�P���٬ҀL�ѣ�a8��&���@�W8��z�V��DQS�;D����E/Vm���b`��_k�p�%(8ғ�hO�{
�e�c+h�l��c
)�pC�	:j�|eh􈝋-��c'II�`�B�I�}xrXr��\t�p�!c�y�aE{��9O��+ �	cJ<ɠ�<�@�ː"O��T����!���N	k���"O�)�HJd�|͸1*6!����"Oh=SŃ��T�´kqb�0�\�""O�qH��4�8PB�9\)> ���n����W\C��Q�*���0EAE!���|��pQI�IRq��)v!�ĕ"r]+Oخ=���t���!�$<��M��D�4?�.#��K2H���O��(��9dE 3�҅wHV�ZJʵ�t�	}�O�u�d����%X9F�,`�'-l�ن
��鬥�C��3.9:�����'���i5�Ɔ*p��:`�J)r7���'��Xy�cقxZ@����z����'���H��j�K)B6B5��A�'���� bTz#�i��"K7+&L1	�'l��S�`�� � �.�dj�'YrԈ�--}��c����4�8�'�r-�J�u�� 3b�,$+�'�j���h\�/4L�"2,��T��
�'��	��Fѻ趌��L��L,�
�'R}b�]�6w�p��r�ܭ
�'�2����ab�hG���mNd��
�'��p0g�ߠ.����a�g̜p
�'LT�#h6kw$I�m�2H�2Y��'r����N�)��0��-[�wr�0�'?�h!��%v!xd q�}HL��'v��R��f-R�P��\�k�.��'{b�&kߓW�51E�f&<j�'�Tɻ���#��H�D�Ө)��D	�';�����ª�@<�H� Y�	�'G�	����.i��ЬH�<��0��'þ�2����6;�0Q`�ĕ,2�k��U�K�w�H�j����E�?D�Y5�
&X�i���K��)0D�`36=�Z�af�4>!��3�/D����A
.��6ˁ��v ��L+D���5�6�ҵ�+ob���)D�䪥b�$��h��i4ȸ7M3D�`�Q�'b<�q���"����t"7D� +2`��C�<]"��8M�ĝs7�/D��2� ��1 �v�ȝ|�!)2f;D���SJ(��Ĳ�`m�F!(�7D�,�Eǒ��`8���E;
�9C�5D����BY�7�t�j�)�R@��b	2D�� �t�Q-,7"eq���/���$"O� scT�Y���4$�X��z"O��+q�(.�E٥��(Jl��"O��IB�@�j4��K��V�4�z�"O��{�a3�.�rsDؽXH��"O�qJR��$
2�9 ��#����F"O2����<Q���3B��	rn�Sq"O�qg�^��4+��7a�uV"O>��Հ�3�A��	y�B"O굢v�Q.~�f�C'$��H9�"Ol�9��Q��Y���JE��х"O$ԙ@��$��=�N��y5ZԚ"Or� É�|�~0�W�O0 L��"O�lj�Д'�2��E���?q��8 "OY�ħ��6H}�Q�B!/o���"O�B��[�\�6����fTE�#"OP�)Pl�^Ў�hΒUI�,�"O���va�R�n\��"��	<��c"O�jr�J*J��bF�1���"O�ӧa��.�b��\#�}�D"O�IA���t�V�/N��a"O�(���Op!:�:�ȫ4�=�"O ��Rh>"��0��8�cU"O�XVX�^��A.^�v����"Oj�@ܕ��pzQ&�]� A�"O���1�?m�$��
�#^M{�"OX9�������H�3Xj�"O^���¢��P��DE��YA'"Oҽ���?U̬�e�TLʱ�"O�0��G�T*	@c�)S��u��"O��[�,�,��r�ƦR�h���"O2���!B�� �"e�J���y�n �K)�I	pf�����*�y2-*
���ԊJ��Ty��D��y2��0x���)��d%��EӺ�yR�ۓBf|pZЎ������d����y�b��\n�V�@A�����OR��y"�ԭ
Y�|�u�V�=�V��o�y2$�%��`	��ý0@�=�2�)�y���l� �rI�<�J� W��yb��>���o�>D�d�*����y��
�*���Y4��9�����y,�۲�S��(e��V΂��yB��3,�I�$J�P�QEe��yB�M�g7X��#�/bp��T㟮�y�O�o�ܽ9b�H�lu^8�+���y�ߖ+1�r���]��[��y�"˧#�<q+c�\ |�����yHӑ�Tk���?ɸ�����y��R#x����ƍ�b�n���y"k߱f|��" {>�-�%a-�y�kW�Z�0�,�{�����['�y��Wln�2��>x��<ps	��yBG�)s+��>`��)���όu�$B��!BV M�0��@����[��C�.h:4q���E��[!�H�|v�C䉿A;x�)4mսqbj�kR�?��B�	�l/&)3&�_#�\1���Ƶ<��B��!>����&`Ak�:�(w!�#R��B�iE��(O�R�*���aȌ#|���'��d�o,C���p�!N�&b\��'E��I�J��ZF,����(ҚiS�'-���E_"�̈���3,x�'^a�O� �*�;ъX�>������� �-{v)��~�h�#���$zw>|��"Op��t�U�U�.<A�a��Dh����"Of@i�M�*1�n��ҩ��p���Qd"OZlٖÜ�Ht�](g��r45x6"O`h(�I��:���
p뚉!�<��`"O^�ѡ�Y#��f��.�XrT"Of�0h�=�
]C��ɠ~�DPr"OZ�(�(_�_k�@CA&�R��9�y"阿��L���$s�qi$��8�y���3V��c`�%�"����
�yBFS�{��{�Ԓ}IXQáP��yB�ڀq2�l��$^4w3��!�S��yrĞ�L��!$#PdL����e�$�y�	�:X��y4`Q�̐�y�U�&s���wN�0��[a�;�y�.47P1�žt�4�hU���y¬�4`�bA��#��@c����y��Sx��a��G2Έh����y"0I�Z��C,��`'̘*�y�`ݵq7d8S�k�
:&�qd�V�y2�E��E�
��1���fI��y�(R
O��@���wJ �7���y"�5� =1�P��玽�y�9\Ǻ�f�
�]�����Ȕ�y�/�$s,Z%�0��Kc��"�ybǞ�sbDc�DT2	���i���&�y"�V-V�{���Tl�(�V���y���(��c.4E��bB��y��F2%���kd��∩#1�ל�yr �=�E��E�^"�@0�&�y�l�29��A0@ʜ)@ͳ7�]��y)�5w�~�g�S�Th�tA�n���y��׈��q 
u���S`L��y�e�O�]xw��m�Z��#J��yR�ם;��+BA�k�;G"�'�yb��Ca�p�'��)v���ԁ�y��U�hd���f�P��󇊪�y���"z3�PC� K�LD=9$�͢�y��U�oѠTj"��vTm�F%ǟ�y��$��� �-~u
,	���y2�M
�q���<q�a"1hA��yRƞ1�0l;c��ph���[��yR��	z訠KA,Z���;d���y��_�V ��"�Jh��z� ȥ�y�O
��`P{4FK'<�W�	��y��W=�|��AфvNŹ�D*�y��E(d��̅�t�@e*�fU��yM˽X'V3��کe������޸�y��L�qY�X��^gPx���y�5t�$ @�\�J(�w�۸�y��7wma��c3Sk�0�g��yr������$��N�xP�����y�*K�K���cwl>��KJ��yBG�T;���D�""��1���yR���KEF��u�丗�@�yBlǄN�V�T����ث�$V�ybc�#���f���w`*��'�)�y�E� ^�֭�7��1nq�Z�B@�y�ER<= ���@�g��@œ�y��U�A���t�-t��\�$���y��8 c��Ҩۼ{˞��4'C�y��|¢�q����%2=��¼�yR+��#ZhY5��+-ཻ�)W1�yB*Z�k@�c�M�O���D*�y
� �aأ�7 <]!t�0L���J!"O�� 0o���������x�<hY�"OH�ە�
O��LO�2�q�d"O
��CA��<��e��*Ǘ2H>���"Oh{cn�kO�,(p�֑TA�l��"O��`��F&mZ�K@m�"%.л&"O�а�i� '��)I��U�A���U"O�8!$I)ϔ�Q��ǽ���"O~d	w�'�T����#��x��"Or��Ö́,���3o��g�4M�3"O lr,Q�-�Lz�O²q�^y¤"O$��直0T��9@���2"O���a<?�6�{$�>&��p�"O�F C=k&�;�C�-�r��D"O^�W-��J��=Q�ǐ4�L� �"O��B`�M�
�X䓐�_<j��[�"OB�pc	�_���Z¡R*q~���"O��I[Y�(<���խ��\�Ru�<�A� ���C�&E�,l�ٵ�Ok�<�dl�3��cF�*�|�� J\�<���@�Sz���I)N9H&G�T�<Y f� �V��1��*�mu�<q� ��LZgA�%
� �t�<��M\Z�=٧fݏ��j�J�r�<Q6!G#kr����2ܤ��jEr�<�&IT
u+l�T��/ʺ��t�I�<1c��1?d���k��MP��W{�<��e\�Q�.丠C\9��J��t�<a�A�p�H	��F�Y|� ����u�<�2ʎ�G�t��Fӕn�`�S�]p�<�Hк
>��J4m�b��3���s�<�#U�_`�a��P;g�8I;�A�o�<���@�R�x�P#�ԝ0k�l ��b�<̚�Wt�@bd-{N�8�`_v�<�$Et2����xJ`蘢hZp�<�a406<ܨ��ڗ.��Qk�a�o�<����h°�C3g��6<�tE�m�<�$O��m�����!E�;˴�2��Rk�<�a-��,b���s��O���!�g�<%&Y�w����ǰ_��P��Io�<كE�R�|�Qn]5Y�D�᳋�j�<�4�|�d�+c#�.���J�l�e�<�4��=O(�5�2��-$5:E����V�<�Dg�+E{\P�$%'*���xn�P�<��/S�K���Z#M
:�V}x��S�<��H/��:⍆!���uL�T�<)2b?)*�,�$`���� 1v��R�<Aub��o�E)��H<g��Ѓ��z�<�ӉҪ������5'��(U��{�<q�GB4K}H��gP]d�9�!Go�<�q�*-v37c��b�ĽS@bd�<�M�24��ĉ�i�!Z*����b�<�b��&D�����G�m��9�iF�<!%%3\�w�a#��Z�`�B�<��$�6l��&9�eZ���A�<9˔6p�h�bF��W�Ĉ"��z�<y�G�>a4`�[� �!|M܍�d�E^�<)sZ�`�i��W!S�N��Sf�C�<��(�K�65ٱ�Z3�I)�L	v�<I�
_�(:@Kҗ�����Po�<Q�hT�u,�8#B��d�wHF�<��-�6x͒-�!��6fP��%(H�<��j��vP�ȁ
���P��FG�<Qro�$㚠�jגS<2����@�<� �{��R�x��9 "�ي{s��"O.�P�ަ��qgL�Fsn\@"O�0��r�<<����,&j�0rC"O����Z�SxP���mR�s���"OVC�*�),'d�� LP>��*"OИ
WKj���+" C�o���"OT$;���;F`:�.
�E^��s�"O���#��{h�I`�-A(j�;S"O��0V�R�:��mP	s %��"Ofq���U*.�fM�P,�ff�D)�"O���g(<x��1�E�_Wh��"O^��p���|��j���9��p��"O�D
0�Eb�x|2F!H��,ɒ�"O��(ˏ)�@� ���N���"O����`�
F`��OY:�� ��"O�i���;$>��o���(�t"ON����)S����CUɊݘ�"O��j����a.$E�a�C!5�"O��)�B��%��b��2!��(0"O<���*ɘ� �YVo��Xq�0"O�,i��޵w,���ؓ�عp"O�}xv��5*X���Ί� �>��6"OL3��[�A$fE�"G����AF"O�I�#���*��Ap&lz��Q�"O@���c֐����*K/��ܲe"O�K%(���r�Ęji �s�"Oj03@&[9/��X(��zE�"O��3��88���sĊ�	���"O&���P.Y��)�0JT�q�v�T"Or��T)V�Y�Pl�a�X�[���#�'P���!8����F�75����'p��$n���(�aĢ*��Mr�'=Ha+R� �����]�1��'0>�Zs��yL(��@��a�ΕC�'~0-b4c�
 f�����6H��r�'v�)��P@�����<<_��;�'���:'��N��p��C0:b�r�'�bUA�P����O�-�LP�
�'���M��a��%�P��3� �Q
�'�� ʦ%�0%$Z�Ϟ7A�M8	�'�4]���@d���e�1LƁb�'0m�Hw����R�:Ι�
�'{Fh k	H�	��k���
�'���Dj�4b��(�wǋ�܄)	�'p�٨� �+�v ��*ϔmZ>���'\�x��N�5��d��a��x�'>P�	G�K!0�$ȹ�ȱR%,I3�'�>@at�y�B큠�H�M�2�',�tF�TN���+�	B2|� ��'��Y�r兑�0�-��6���'U�1�&jX�.80��v�Q�
����'��E#n�G؀�E�L�9͢�Y�'�ty����vH����&��0��q	�'p�4�uJ�%E��+�����a��'���@�ʗ�A�X�zT��?dh��'��(�G#L��R�Ha��!]��բ�'��S6�Φ.d� ���,����	�'bnDX	��٨'��&4*�x	�'�J�)�M�2	���\�պ�-S��yb�X+?�����˝�7��µ�$�yrF�K/Љ�`�ԙU����yBG�/i<�i�G��u�������yji�Ō���M�$���y���*+�rx��d��pag�y
� �x���0 H���w��k�"O�MIp�Fj�P���@hh䱩!"OT�k�vWh����0a��V"O48����8G�����'5E��ʱ"O<Yg�^�V�T����Q��l	@"O�Q����i�x���ف8�R� "OlQy�	�� ] �'���R|rD"O���#� �|ꣃ�&҈�v"OdLYS�=?���`aE �Ԙ�"OZ,x!�U��eoE�l f9�"O$��E
�1:��:3�X*p�#�"O�9�C22\�M�2�+(ʹ9!"O��g�M<x�k3kE�A>օɱ"O��)���:[2a��*E.4�8�"O܄��T�I�2�/�,�8p(�m�!�dٺ&_���H �|��y��)H�!��J�T��D�F�	v�H�fV!���g�1öJYl��8Xņ�E!��D�T�,5��"K��i�&�e�!�,u�e�PC��w�@�3G��X�!�$�LӮ��C�� ��)b�O�!��יR�bD����$P��C[v%!�d��� ��Rv6�T���ƺ
�!��_�0�`lC$d�6{�ZRb�>i���0.��+O��1a]��y�E��<�����h�|����y��d!�<�f�G?XO|�k�$Q��y�鍿rʸ�� �:L�Z40C�D�yb�'l���#��x��!�qj���y�fK�5Ƚ裃M�p��X�M��y�.�c�Y0���V�0܁��!�y"�8��p��ǒ#cZf����Ż�y�U/j(���[Q���I�3�y"�Y�j]����Y>��P�*��yR��R؀��B��R;��p��yB×3zR� ��>4�A0 ���y�gԥa+ t��K�:�f�0�e@�yRo2?c�z��У"�|�Gf4�y��� A�p���o�4k�_��y.�JiZU	�@эgb	k�a��y��]>����'[�uv��Q��8�y���M:�����i��y�BE%�yr� G� �f�$����yr�Ѳr�X�xvK\�_(�er�cO	�y2F�wq��S�
�]��JAf���yB/U����kR	F=�I��y���~p��TGZd�)��	���y������kJ7<jQ#vF��y���S����͖(-,%�U�H��y��z���
�EF?�n)SF�֛�y�k����d@��sf Y�� �y�D�8/�(#��-s=L rVEE�y�Δ�gD�#��^�98�����yB���R)H��E݌!�<��0�]��y⬗�>�
\t�U�=�5�g(ą�ybD	X��ą�r��u���y2l��~�4�`��1?�x�N@��y�A�" �d�I����k�R(��y @���XAc.a9X�*�E��yLܦzr�7$ʢ0�^������y�����"����ӱ-n��a�c��y�+�h;b� _N���A%�5�y��8?dְ"�N6M3�E[1���y��\�Xu��GƋD4���@ N�y
� �qR�R�I^3RI[�$!�"On٫��� ����GMl"̃�"OBi��l�)x7z�"@��DnrLr�"O��V�B�`���	7J8I��"O�	�Rc2<��N"x>Rl�e"O�:1!`|+A&��,��`"Or���f}>,�z'%�O����"OH��c������y� �Y�2�!�"O�q�BNS"E�z�s'�5��"O�m{#΍c�hM�F��ͪ�"Oظ!�GI+����acrڤ��"O��h�$V�3p�A)'(�a��\Ȃ"O���$E'Nt��	Rg�}Vp��Q"O��g"%r�V}KU��fO$��"O�Ųrl(l�x�X�'9�a��"O�QaCQ4y��&BɄn���G"Ot���O_�(��!�M�K\�� �"O�Ʌ�!T*.��D�Z4��R3"O��qB��S� Cx���T"O(��,���:�Q�B�6NT�Rr"O��t����b@ ���l����"OV����
-��=atj�m�@�A"Oj<����x���'�yb9�"Ox�2�n�9�|���h:�K@!�y"�*��a���'(�@ȅK��yr�T�0 *��=  |D�dI�
�yR"��
�y�oƘ�1C�F���yB'�6s3�}�3�S�vކ���BǍ�y"�&T��@�B�j�~���Ï�yRGA�z/<� UA�$hB�+Q+P�yBgD�d�p8*��9\���+�G��y�.) ��SBdS!(�J� �e��y�'V�b�)+\y���С�zjC��2oBnq@�E]�W[��xEd�%�tB�.�����|���N )�:B�	�b9H��'��E��	!�o��qP�C�	�u���BL�E���ҩ�xz�C�I1"_F1!s���,ٻu��8v"O�$���%(��}����5so���"OL���BߊF��@͙�^<��"O�3��F���mR��I_�h\�@"O��7)!q|�������guv!�E"OH��'�2\na�d��sp�}`�"O��#5�*f�Z%�6"j�X��"OL�w���A�f��b�*OZ	B"O����#m"�}qd'G�A�"O~hYD@ۃ*2hp�H#*4hh�D"O�\2&�B~�ሆ��	Z�
"O����C�[9����ۙI��0p�"O훐��]�P�*q#L���q�"O�逖B��S�4��B�%�v��"O�[E��O��BG��,�6=�Q"O�<`WA�!�Pg�f��C�)D�� d�?xܜ�"��&u��:�%)D��Pf��M���3s0��!��4D��y#�׋n�j��a��<5^�!(D��ՀB<W0�`�
IL����+D����+*vm����!f��58��$D�L�oJ>2m.��b<Wν�d�$D�PZ��F-s,�4H�H�J�Θ0r #D�p����h��ї�ۜq\z|�5d D�P�1aȠz�� �7CZ)�:���L?D�4@�gУ94����T:Y�PcW�;D�|8���0$ ���t�Q2@�����8D�� ��&�z�v݁4�2C�F,KE"O^��W�W�G��paH�1RDLK�"OH�;6m߲2�8@U���Pn��"O�ɈejX*41�w�Q�k=�h�"O�0�@�J��bWN=-�;c"O =:L��S%��y�n�2RAb`"O.��3��}���3eB#��q!"O��rQސk�|�v��8�L\�"Od]sbE)BY@�KC��t��"O<�	ƍ������
���8+�"O��2a�%|�y����@pr"O"�a�n�	�d�a%V8L��x�"O��%Z�|I��	�p���7"O��KG�Z�"�X�+5�D�@u�U"O���?$9��vM_� �j<�"OXxQ��\������-�ĵYS"O�8AC(ӆ4�(������E{T�"O�(���<Ffȑ1�˟Jp>�*"O�jRA��t(�!�Z�{k8Y�5"O�$�����!�*�;��rJ�a��"O�u
)J(ie"�w��!e�\��"O�@[�矋H�b���ϛ�<��H��"O��P����.À�Ά���U"OX���#�,T2�"��tʁ��"O����(\�ڜ�R���S<$53"O6�V��*`(��%K2���"O>�'��2�6Lapd�9.pYj�"O�I���#9Et��I�J��"O���ט	��y�b��2%�^�c"O�����γ$q������x�>�:p"O���L�>lQ0͒��J0PB"O���'��4�`�2�� ���"O��;s��2$���"�"'� ��"O���#%[jHs�"E�VuV�{5"O��WdP+@�� 9�B��ym�$"O<��`�؞Cި(��
�>Rd$ucg"O��K���57�5cA��LP����"O�M���',���$��>6ȑ�"O,��� ����	A��1Q"OPl�p鄺d_�9뒍�=\�>s�"Ox��C�$A��;I�!"��"O����G4|䍫q�U�W���!�D	j�\�K�87\	pA���!��U.1�(�U�X�9	�ArS��}�!�* \L!��D.��Q[;�!�$��r��s�J�褻�o��b�!�\80�d!�0�ă@�(��!ʔ@�!�J&_��p hY�@����Vm8!�d��r��d��
6��H��P2!�d�&(Z�������b�%E=!��P�nYb��c��ŧ�f1��'Y���&"1F�ѡ �M����'t�%��HL;ڐL(�@��d��'&�-*���|�u�&њ
�x���'��Y��o/15.�Q⛹xy�!��'���Cf � @�x�O��`���C�'Q��3fɚ�?s
dk�l��V��L�	�'�R���	'�B,j��8Y�(p��'�Hp��e_VT��F	JT�Ƀ	�'��0$jŒO�iZu,X*0�lI	�'�<�Tz������� ���	�'@���Q!�!d��PB$�0��'�rE�q�7�B�ӐKS����
�'Z(�3��C/X��9�n�Oh��	��� ����H:c'd�+��ۢ����e"O��*Q��r%F��$GEF?F��1"O�[��m>���GZ!�3�"O@�5C�<3X幠`@�X�A�@"O�Q-�4V�f�"0OG�j��u"O��AD%�0E�$���<`_�,(�"O�0�efU	]鲕S���zUd�3r"O:ݣ$��uC�i���A8W`�i5"OVm�A��y��]�SC�5E:B�x3"OĈq"��43�(��(6R�""O���|6��J��L0t|K�"O����x��YAʊ�rH�A�"O�$ P����IAR'�� H ��q"O�l����7��T�F%m!�B�2R�!�ݾU�݁@��.5�D���S�w!�D�4�P"$���h���_� =!��+h����S,Mg�z��!�Y�&���)��M�.: �q" g�!�ą�%�,��'��J���q��!�	GJ�C��۬qE�,s2`�E�!�$L�
�� ��*G���d���X�!���=b;�0LO)ܹ;!Nɒe!�ę�a��u�b��MZ��*��4<|!���y�ش��\�fE@���@]�d!�ǮjژѲ���&�J�X���!U<!��8�����؅E61(v�R�	'!�$�7ΉhG��Nj0���d�5x&!�L�C]>tQ` Lj��酤��P�!�?Q��=���Jl�p3dD%z!���$�(R�+��%{nS�C��9k!�0 /d�)��פ4���h��ۏ\�!�G&+���'ș�j�q�ē�~�!�ړ*�L� c�c֥8���5�!��U�Q��'4�|��	�I�!��>농�DoȩI�fY��ň��!򤖕nNzu��$��d�.�!�D��U����G�*�ni�FA���!�X�["�	C0+e���Hrͽ�!�d\�F�}qm�TyF<���Y�e�!��*Q�LIyd�%m��a�6	λG�!�3��1�-E�6q������|�!�-Ez�z����	4�d� n�h�!���+|�9è�L�ք��
^�,�!��"��PS_���y'�L	�!�$��mm��3���!
���hߧ#!�$����Y�HBs�H�h�[�!�d�`�$��E��2:ܐ�!��L@!��u�n)�uOB34�ɉ�
6!��,A���/VO�E�e�:4!�d��6$��Arm��F,�\82��!���2i����3%\���G(V�!��3 ���t��X�䨔��!��l�l�q���v�
A�0�T�Q�!��);�d���m <F�ډ٧��2�!�䛥�R�`/(a &�Z�!򤑭x�p|y�L��L��a �E�^�!�d�:n�Hh�G�-��ztDT�L�!�œ^����X#e�*8��R4)|!�䃯R|8T����(�$���H9!�dP'2����#�Tj-dкaH�0�!�dB�&1����O%�9z��Uw�!��3Uv�z � �(	v)Y��S3�!�dQ
&M�$���;3�L�P%D���!�Ν":�A�mةN���[Gcŷs�!�� t����3u�i�'H��j���"O���W)��I��p*wkJ��� e"O�XrU&��xqz�qp!����� "O@ �2��*t	�h��0K��qh�"O6���AԸp�B�@�o�,��xj�"O�x�(\�Hj"F$]��L���"OJD"��A"j���[���&"W�x��"OP�RiS�*��b�N9�d1�"Oε�E��dt6}1�F��81q"OZY�T�A��^Ia��/>����"O��'&�80�X���ň	���+�"O�䩐��S�8Ȧ�U�Z�"�1c"O��k��D�� ����2�>�KE"O���7I�/B��q	W"%FY"O�dK��!,��!m�;���%"O�X��N�E �B����P���H"O��{�Nw������KR	�L��ȓ8n���w�%1l� ���� ��ȓ^|�f�1o��0�E�*2S����`D���E�x�L0���|D���ȓ�ɳ�gC�l���;Q$��{eB��:�����M�{��%�b��3�B�	�%s$���kͦ���w�GR��C�I�n�~݃�#\�Q�rY��k�ylC�I-2��z3��b���%�?r<C䉮c�(EBt�A
uZJ���iC䉄M4��#�X�q%(��&��FC䉨im`c��L�>��ؚ��;&B�ɕjF�ͨs��2ǲ��ML3a�B�IR�b9j�NѲS'���+���B�I�1q�0�v(Ɲs��Ӊ^��nC�I����!u)�_�dx��h
��XC�I�n����Q략gj>ԲT��r
C�	�V��aåß#��9�Ը7UC䉬g�EKp�Y"͎U	�����ȓ{��I���*Vp@�ݧ�
ćȓho }q�R�ܥ�N^%��P�ȓI��A�)�N���zb��$j
���z��5Y	�Bgʧ�H�2�T�<1�����	@P0JՍX�<qщ��z�� �!�0k�^5��
�Y�<y�N�r�^�#�F�3�Z͉dY�<q��f�~����[)u�xhင�@�<�a�h�-���!+�%�	R}�<��g�V���Ƙ�;b6��y�<9e�-c�r�ځ�U� �BI�7��r�<�C0�4IWH��	v�hGn]x�<9�^�H�X�JE�9!�\�"FO�<������P��5~���%@N�<� �[�,�k ����E�p��c�<i���n*f�bu�g&�-��Fb�<Y�
�B����x z��Ex�<����/�a ��	U�T��p�<�'�[�s��(�I�P]���eRo�<aՏ�7*�`�CR9���J�g�<���M!T%+T��4Q'vm���a�<�?sf�蘷-�����	6��a�<	�N�Q�h�RG#�'@n:x�f�
`�<!�
٨/�!:B�cN�"l�\�<i���1`�A T-!&+<@�D��t�<��#ڿ9�t;�2n�A��Fq�<q��P*&�����ݻ�C�l�<���B�Ӓ4ZwJ�t >�[f	Rh�<qfٝd�29��n؛&m��QVK�i�<� �-��/,�*"偮SO ��"O�Ize��W�\0��
Q�3 ��"O���EHЫCY ��ki�D�K2"OXu���D��.���Y�_���``"O�0F�1U �q%)_(Q�¡Z�"OԬ0 MP�P����4<��ɘr"Ol9x��ݣc��XhsGP�����C"O�\��h�Y�l�WF�W�Z8�3"O�!��l�o$��$̩er�ɕ"O����"�\E��+z�ѣ�"OFذn]rzQ��dB��"O<�C���Jib�M���^9��"OEIVH�$f �5�6@�<B0"O���ĢD�]Rxx']�9�6u{4"O.���k��]�~,���W�ls�"O������Wϐt+`dJ�o� ��"O1*�m|��[�b�t��*�"O@�:����8pX�! F�5��"O���R$ .5j!/�1�#f"O�I!m��ʔCB�������"O�\˲�ݞ0�8��ǂ�\���rc"Oț���������w�n) "OD�*񬅘��p�dLV�2"O$����Ww� ��CO%m	��"OԜ��"�fMSVg��q��`��"O���DߍoF^]1��Q7;Ra0�"O2d��呧xk&8�Aȹk<��q"OPܡ��#�PH�T**����"O��d�>�6� '�Z	;�X�T"O���&ā��P� �N�����"O����N_�����×�:�>��t"O���Տ�r���'�q�p�;g"OT�+�ₚU�N��Ñ�d�2�"O��Bw�W�(ɨ{�d_	;(��ӧ"O��%�1m�)���
M	�"O���fK��6	z=jS@�
9J^T��"O��j��=c��<
��	}p��""O֕;��R��m����9Y��Jq"OB�[Gk1,Fp1t놌a����t"O<�WFA�^n��bkB���\�e"Of �H�p���q���)�J��"O@%�U�O.?=��hN'TΘ��"O1�ԡN�2�N<���?�l��"Ol�B�fװlL�����5cp�d"O )�e�Ԟ K�P1�L��\"OXX���ԣ�xis"��>���k�"O�%����4��٨��^�$�e(�"O���� �nJ� �����w���@�"O���7"�oS
Gi�4"O]IG"OzmR'	l��LZ�%��$<:��U"O��!�Z&t��*�f��1�(I""O�0@��89l�B��$xR����"Op�0�H�G,�zE�Ce�p"O��Q�BR�>���1C�v��EX�"O8��D")Y�,��"��Q~�qPp"Ov�z&C>h�̓%+JCl�ae"O����A�% ��qB l��	T@�"O��1T�c��%a�\�p��P�"O�jc���a%��Eǆ��` �"O6����i��� �|lR("Of�ȁ�%z�*|C�ɰ��9D"Oh�0��[��򷡏�;M��1U"OXe0�,�7���Z0��'�=��"O��A�
��N��1,�(Z�TaI�"O� �����'�H�ZS�EH�l2�"O6	 7'�	�`i���X7rs��0"O��8�`��
���"�IR}W�m8S"O^��'	*+�6m�6
Y�S��z�'�v��˻\z���4*�|q�'�Z}��j�1O/��#�&k��I�'�0�؆/�F��pC%C)��xX�'�d����:+�-�hϴ�2��'��E+S*L�j�|��^�)f�j	�':���&D��)f���3��ȓi�qi��Н9���IsN�$�f$�ȓ4d8Q��/K��y��'ҀR"��ȓmnp���z3��RG�_�b��7z�p�.�4d�Xڴ(=���ȓ[j���E4�����!� �^`�ȓ3���u�̚Tx�T��,;m]���ȓ{l��X7�_�|�ĢaA��v$��ȓc�r�:Wa��^�<C!i��JkX�����]2U��'��p��(�=U����/j��8�c��q��S&�q܅ȓH��@qON�� i��B�L'�مȓq�uH��L c�8��H.l���ȓQ\�(aAΎ�T�����_Ӣm��;*\ @'�1>ȵp@�#�6���)�J���ᫀ��63fL��&|E�C�Y �>��-߂2�d��f����@9fG�mC�҂}�RD�ȓ>w
�iҮN�K
n��c��V�Ju��;��\���з~{vyb���e��B�ɷn����6T�t� �� RdB�	=i�z��!�0c06�  �Wnd,B�	�3�h�Ҵ�[&l�<��� T�?��B�I-vj���΀XQZ-��,W�C��49Ղ��wO (8Dq���m�*C�	��ꀃW��"r6e�P�Æe�@C�ɺ>q	P0/�3���$��b� C�>\q��1@�L_��Cc�?�$B�ɯH��AP/dD�剎�E��C�I�9��-+P��9% �'d��C�	Gv��gȒ��� btd�2~D�C��6|�(����%	��D�P-� Y�C䉊
X��@��~>�\���,[">B�I�1�6D���.���kS��Y8B�	"sXZՊP&�9eP|`"�@LD�C�I>��a`�ùc��ѲaW��B�	�BU���DT !�`i�HƂ(7�B�	�\�����^68�r3n�!,-�B�	�tB�D�1��8~azR�ަ�~B�F��(@�`Ml
�كL$?~�C䉕R6���)Ԃy�Ԑ �.g#�C�	�A���H� �t )S%��[�C�ɺ%����K�q=���O��.C�ɤZ�<�ؐ6J��9 ��� [C�	/jjĒ4��@v�6(�5mC�ɮN �`X�㘪M���	s��u}�C�ɤH�HY�i�7m?�T(a�)H(�C��i��H��� d��d�mלkֆC�Ɇ)p�����ǜ6���a��	?a[B�		^��M(S+Đ'����s+�	��C�ɲl9���N�Hm~�+�`ƜE�C�ɺ]BΥJ舏?� Xd�% ��C�ɜy��,�!
��a����e؍M}�C��([M �h�Ą�i��%�Ճ��B�:�e9FG��E��P�A&m�nB�)� ��g ^3���POH��"O��A/�P�h4���qv�1�"O"L�.�)s[>�H���=BV��B"O&q���	'֞��N�����"O�0�Â�F}��r�mȗ)�,��"O���a�?xH���I�}��@��"O�+QKP=&�:�)2�ҩP���D"O�8 a��
\kr�
�v ��Җ"O��� �X�"�
� �v-�"O�m�f&��#<si<S܂\J�"OA�S��4zk(�����(��`#�"O���E�
~ތ%#���#�:�`"O�(��0��C����1�b"O�Tr�X1R��pI��\괌�Q"O8Hҗ��D��ixA�$s�p}B"O�x�K��2"��r��D*)ԮM�4"OX��C+��NlLj��Y4Y�� �"O�!#s��g݀|�у�+A��! "O@T�C�H wi�-�$t@�"O({���&9���3�')`\d�A"Ov�s��]03������ŝV����"OJq"A$ '*��]�'Ȏ�9@t�'"O ��k@'�fh�P�Q�@��Is"O`=�p$�u���yG+I�1:���"O�q+��%�5`H8c�L#�"O(�1�3-G�݊���$����f"O\A�0ƒ�-�D!Pfn٦"���R�"O��S�@�Z� �9o۟Ji<�"O��z���1eb!�M��Xz��@�"O$���#U�k��$�c*K�/\dy�""O�%0$6Q�)�uHG�D�0A�"O^���) �\�q酀l�}ҥ"O�,���>+��y�����d���)D"O� KӦ���!fD��"O]!�d�D���q�K�f�V���"ON�A�c�<l0�jԌ���z@ʶ"ONة���u�`�4�ӑf��ɣ"ON�
� Ԯ����Fߎ^n�X�"O��3Հ�p���uٸat�A"O�Y���u2��"G�\�,r�"O��A6�M"w��̣�G�	Or$�F"Ox<��i�N�~u�3M��d#�"O޵����UF̈a�Ř�hz�՘�"O$�:�QI���
W�Kvd��2�"O,eGDّ'䈑{ n�oʽS�"Oh�u	ɞ('�5�A�i&တ"Ox�dM�=~�i� �v�)A�"O�9z��ڬ<$��i�%�2i���b"O��hs�СL$|(i���`�֤�S"O����)?N���"��A�D��"O ���ګ5�q􂃁�\�q"O
�1f�$s@�$�R>1E��"O����-W���w)/J� �:A"O�����	$�Y+T�ˇt.�:�"O ]hC�����GH"!jp�`t"O�y�U*@�AԠ�!��ڨzKPD�s"O:@b��
6L:�h��O}Dx���"OTUI��P&#�P�t�P�eGz�ɰ"O�����k����A��5x�!"O �{�d"U�ed �>4$<�"O<,+c_v�pH2��j��L�d"O�X���9��
�Dڊ!h�TXr"O$	�s*���n���(]$��К7"O��bP*F1B-
����þm��`"O� ���H�y�Uɧh�>��h�"O��"�l�Xsd��Ǉ�k��Y�c"OX����	�
�����{����t"O���(��L!��'%5:��u�3"O���o��Q�8 � �BX�(<A"O�h������&��ec��ve���"O:`�2��<?���2eD=d���u"Of��v�OA���'䎺n\>���"O��q�	U�|���4�nͺ�"O̤K�3���@���n�b䫡"O.Y�!KҭjT"%�"A�'t�Da{�"O�l�B\&^�^��ro�C�$���"Op��R b�����O(}Xڍ��"O�-*E��xQ�*N>�R"Od��$(Ӎ$S<����U�'>�r2"O����rY`����t#�Ё"O&]��Z�o�\��@�P2s�`r"OtL�u@�A��@�)�'�J�b�"O2)��/�,`����v�>�b�"O�(�㘋�����<H@�1i�"O��CЌ�oz�-�k,����"O���3�s��9�O�Y����7"O�񨆋
$Xq�:4KHD�^EJ�"OT�y��>Sd)�5���L�"O(�h�N��{���CĽy�.��c"O��b�˛ �<��Pf��P�>��B"O �����K����a� r �`"OZ����"-��8Kw��#�V�� "O���]k@�RV!�\T���"O,tc&g�2G����F�O�O?�}ȶ"O2��@��B�NI��8�T���"OL}�"�غ�a �E��2�"O 	��,z\��@�D�*���"Of3Q	U��� �ћV"u@�"OX<9�!Twp!ڣ�Z%n�ڜ"""O�X;'�S�j�y��H#9����"O�r�f� H|#%`:J��r�"Ohm�g �<\C�	sD�-?ބ�F"O.L"���<��)���ގ��*�"O�PY��K��|�+�a�\Ě|��"Ob�EzҠ�����V����"O��*g�o0,�'ꜻ=g*	�$"O�y��e�=#��٫Ĩ�5Ie�(�"O��橝�9&r-x gߐv+�4;�"Ol�9���4E�Z\A�/ޜI�Δن"O^)�����*�����A3c�Lɻ�"O`P���;4P@*��ACyL���"O��L
�L��H�
Dc�Y7"OЄ��U�x(.�x�W)]H�1��"O��r��߬*0����[�$��8�"OTQQ����?�H�ҖM��'��L��"O*�������5+1�
�E�f�c"O,��+Y!9DhܸPD�*��PU����=a���ϫ��Y�� �'aNd���
!bS��
O���N<����S><�U"O�1
��8B7<9 �.V�XG�'��d�;uQ
�������ϊ=k��&�8D{���V:_e��y�i�9���$����0<�J>�*O,�ǧ�C4�)G�-t~��B"O1*P��g����F�+l����'t���}��	k5��D?p���a�2%t�00u��z��?�2����f��-��="��Yd|��<����ïT}
I��C2m�f�KFƟ� ���A�0?	�n΂*�` 9B
A-Ok���`��ݟЄ�Ic�� ��9���;#N,��W�S/�l���"Oz�P"@0���P"y�,A��I|>ȡKgQ����E+NH��m�>�yb��#��Ǯi�tmH�" �>�Zq�/D����ӌ�P1�����K�0اN.D��rH�#�����/x����6�<��.�ڔ�TaډJ@�:VS�a^uI�'A�O��?A%L���D�{��T���i�K�'�����}�FBWT��#%��^�x��m�O�=E��˘*.���k�
�l�:@�?o�OJ�=%>�
��A�%k��yQ�(4,[��&D�@H�䘬A@]'ؒ;%�a{� 1D������~z���B�s������$D�@����,˂��2�B4)�\�!#0D��� �Z.yg�4�2�@S��0�-D��A�5%̈��`~�|L�kk�����%Hzh�h�OD fm����ΘB�ɒnNy#�֤*�<�3��M5OnB�	%yfv0�dLծa�E�w�Y�C�	����X����UA�Ɲ�,p�B���@��KJ22�ڐ��NݖER��O�1ۓB?��[E���6��qs�A�T�$�ȓ8�d�p���� g�B���ȓy��ݪd�5vHXR@ӻRӚ�E~���?���K�_oҥ���j�آ�o$D�ta�ȏMP֝cjn���Ф-D����[:-����K�CH�IIl+�O~�(J��$��-ؒHk�5QT�%�(E{��D�"f�>}�c��G;0=kѫZ!�dS�&��
F�O����i�'{�!�d��N˨�V'�J��RJ��!�d�-%@U���δ
�z �ɜ!�D�<��Y�2�_� ����׍7��{"�J�9�|���"��uW�a���	�a}ҕ>�ĥ��38aӢb���b�W��%���ݓ�%�P�Ɗ?Tt��)D����G�<,򏄟�N��� $D���'�ȸW"��{R��Cb!�ǩ.D�(J���7�]��߄{	%��J)D��pr�ܯ���a A�� )�4�I>:Q���mr㖆r��x!�B�.Y�p��"O~�*��L�>�<�PU/��fT�d�1ʓ��<y�߯=���A��:K��D(�]�<I�@��D!��z�Ց@q���w�W�s�C�	�_ 4�B��6]��%�<�*��D#�IZ��@��[g.��c��,+�C䉸E f��A��z'Rы��H
rc���:��v\�@�($!K�&���,B�	(ST��)�dG2��`�#<���j��h����wjM����t�w�@�"O����cʬ,bSN�q͸�:�"O���(T,~Eh� 6NW	 ਁ� "O�-
�ꞦW=���  �t1��"Oz�T(��aZZ�16nږ�T�Ke"O����Y6Z�����C�f��!"O��;$T"jt��d�X91��`��xR�'/�z�#A�Qn��WA�1~�"E/܌�y"�]4j�q��h����*������'��{��"B����E,t$kv����O�"~Zsȋ��=�e�[�hJ=�C"�M?��Zf���R�(D,q�æh�@�$�D��	7IL���X�GDUQ�̱z�>���(?Y�iҬa ���kĹ!M��(�+O�<����`�
�	4H5_�H���˅c�<� $$���	-���p�� ])BH��"Odk����������� @�!�'T��0��N�b��9�%���V�@Si�$�=E�ܴ��Z'�ԽA��=r�ȥL-nP'�F{��D�=�t9�D˪;�Ha�T�I+�y2�M#@��g�ߴ.춙��Յ��'�����Ʉ5S�ȫ����	_��;B�P#a��B�IE�TM1+ �7��k�>P"<�	ϓ7��m�eg�gA]�v�94b���	���C�\�Â�L�ZtH|��! ���O�%�
[(e����9p��a �'w���1o��D!��	G*����%�O��I]���堄!V�P��E���	|yr�O���$��;E��-�!݀HA���t�&D�0�6�/˔�jl��m�Z�h�Hd�ܔ'!ɧ��Ĥ2O�}���0�@�g�A�~�!��#Df:�+3�M��ؙ v�T�d�d�=E��'e�
B9m�@�Z�M��h��	�'�и C��t1��-�n\b	�';dぃ��~��@�q��)��`*	�'��,A'ӎRm�`�����¼�'5\��l�:E`<[ᇞ�����'�l��CU�7�2@��97V@���'�m� ��^	�)5��|@�R
�'䖼�t�&s ��JcD@�wkTH�
�'�zEk#�R,|Pp���'l��}I��?Q.O꼑�fO�7x��҆ܥW����.LO�Uo*l>���Ń|O��"O�J��,�Z��&�
|j�$i�"O��zr��l��Y`.		���%P��F{J~b�O�(9���0�Ρ�G×r�Ȑ"OX��X*U�z����Ğ���( ��x9p�)��?�\�B�`���P�H#+����扲~~a{����؄�ן\�4�k�$z�bm2�0�?L�������䗦K�- Dl�0a9D��j��*<�B��=|�������=W��@&�l�u$,D�x�������%�G�A��p ��+D�l��&Q�=x��ԅG�>d� �f�*D��3�V3xj��l���S�'<OB"<�C�[�|tUڕ��R.J�`uJ�K8�@$���"@�(&-	���Q!v��q"$,O��'���O���b��R�*�iGfw�,��� ?��ٌwͼ����ҼS�Th�S���x���P��}a�jMGܬ���P.�yb�_+�X��L�BYH�pf]7�y���X�z����F8@(� �P��p=)�}b��r**�|��48	Ӵ��xF�2|�#wȓ|�Α�3��(J!�$�6Jg~��/V;&s�Y�C &5!�P�[��q`����4oz�?y!�d�{`d�F��^�@ �FJ%��y"�	">���Y#�Kb��diP�	.\�C��4
l��a���#Z�Hʄ�ɚV��	�HO�>�i�&���@��gI�|Q��:D�XGj
vTx� ��(2Lx`5�3D��(��`��Ȧ
M�;�
I g6D��p� N�I�RFI6��t�5D���cu��x#�j�aT�����2D������"����������=D���E�ʐ�k��B�$�r@&;D��`�ɮ\ǲ�I,���89��8D�� S�6�A2��	�'�(�G%9D�D���(x�!S$FҜI�h#�L5D�DddF�6ܙ0S@M�c�,I0�=D�� ƕ"�%ޫ^c4ĒA��3s��� "OR���l��M�<j�mҲFtJe��"O:��W�ҩxa)aF��9en��"O�4��H��<�nI�dQ� �"O]:����o^RV�LO�f��"O�m��μ<�U7I�7D��z"O0`K��Q)O���r��[���"Oy��n�h�p驱Aߴy��I��"O"��sF�/Qox��j�ښ\ڢ"O���BJ1���wi>[�A{�"O�37+N<(��i�aF��r�T�2"O��Ã��A������F�FYc�"OT��U�H�N@ZIJ��BT�<��"Ovl�0���;e���#�Jk���"OV��.ȏ ڎ��\l�"O�(�,�$q8u����w? U��"O��ڐeQ�i�4�;ao�~Z���"O��×��8Ax�P�ㆁ\#@��R"O�ԓ�O�?a������
��aw"O��2T�)Z6�`����c���@�"O�<�`i��<o�)
2`°X�|Yb"OҤz�
l�DP��E�U��T��"O�i(�+��D(��ՀI�@�"O��塝%R���f`��C����p"O@|ۢ O/xؽ����&�H�����"!�V���4*���ga�Y�1OX�ДAͣBw@r4�Ž?��z%"O��+�P�_�Y�(ܦmr���"O����.ĭy��<��
�8q"��"O��i� �?F��K7;u(u�"O��a�Iͩ:�e3$�\�M~l�Ѱ"O��r��`r�J6���v"O2����.Z&P!���"r����"O�{�Fǚb�p}X�Ǉ�7ÀP3W"O�m�17C��"���o�:u��"O�;�:{"�,J�k��	[@"O�	0�@�(}L��J2XZ��C"O��� &<�09�ݖQ2�I�"OB�����;�L��ͬ1"��j"O�5��/W�Diu��N��[�"OTlH(1�F=9��u���"O�<���D����1�b�'2D@�"O�h��=Y�e
Sj�X�4|�'"O��Y�J�E�`iA�a���s�"O(L���}�!0u)	0(��}�1*Oh��`������P�J12�',j��D�ýO^��YQO��Ntt�'���01O��zERq6F�Ɛ��4'���t�Ȋ#���(O?7��{xY�GC����(1��N�!�$���`���O-�&���ܦ'��DK]���:���_>�ea"(��l�A���z��QڱC�4���I�9��� ���n�Qs�Ȝ	gLv(Q�iL""�*��k��f�ȑ`��'N��J��4B_��� 3?���}Ҍ��bE�)�ǋїz�:r��9М~ZEi�I�H�����Wi��E+Gl�<�F�� dBf����2�rd�\<R}�P�#��|���فe=�hJ�I5ʧ�V�ɞm�n��5VL�0uf���*C�I# J,��1�8��G-a�!
�����!oS�Ҏ�9Vh#!L<F{��(B�1�DG�p��L���<9��E�h����&PG4�ҡ/D',�C'L`C��!���@��j4B�;v���d��9���'�L!0t�1@�Aa�' 4x�q���Bfh��Ë=~r|M�t�C @D�OT�*��N8����L����K�'`�P�)D\G:���II./ �г�a�PЈ儂�:�����>d�$?���b���y�)S��|P���:�}�h/��x�.�'���A� J��	�
���z(xr���,�d��e�4|�aN%��9�	22�i6O�=<��{��A�5�2��D>z|�Mه�܁'a�I8��D�? ���'��>h��eE@�9�� �/v\��Æ��p>��X�8�(R���&7| �wE�y~B���If�p���v���Cë�Ot��$���`��'���;���L}�]ŋ�np�ȓ�\���7N��4OO�'�x�C0�O'I�E�����J��ha҉����O��ᑲd���y'X�x��x�^iҕL���x2؇��A�u��f8�r7b]�F���Zd��16C#p-
��+U��Y�ƛZ�'�Z��E$�CZH�����
%(lXb	�#)"��Դ\�D �c�^�J�z��UD��ă�c�2{2L�pGAr�Nex��=?r���	�&HcD�$����ւ����I�0KF��uM�y2��Q�['Dz�XU�\�P ɗӟF����(9,�)ɱ���k�7#!�4;|�	���%I-N��S�сm��a�c石)�Rh��*9��֏�4��S)PxL-���)?C֢�B�� �H:��!��#IG�L�Ӷ��'Ȯ�@5�(3>�yQ��D�hP��#BlKR�D�RC�_�@��&�I !�6��2*�	�j�yWI�*���D�Q�\x6��fA�1NQg����t� :����̋
O�5#a曜J���jQ��p>�aꅙ7,Mˤ��6��l�D$�m~�IS�l���piH_0X�`SFB�o� �� Z������D���!�$�Ⱥ J�V���� L:$K�b[�T�q���U.K3p�3�DC� "��E���=�L�T�=!N8�Oq��E	��y���t�(�aA�2]��5E�5�x��i���a��gC4�9v�u��� �
���DuAF�Ӟg��y���a���!W�'iv���@8oW��0I8Ws�9��M�V%��w��CEGQ@nx���JZG3��GH� �쭃T��=1��}(��\z�����љA(dԡT�D� ���$H�@���ɟ1$)��)
S�E9������A� �OId)�[�4u��� c����y���J\@ PO�#�T��U\n�H��������Ų)��(�^�ѝ'�:��d��>C�n� ����n�a�'�f�P`S��(�g�)�46��U `�"�'��[b���.5�%�M+��		�Q���~"(��I�,�|\2����!�]�Sf8g,��F��v�$�׈;fАk��'��!
���/�DA9�aY$��Dx�����5[$*W�I]Ɓ�b���.C	J�����#<�R�Q����y�?SQr�H�/M�+@�Z��M�w
ʮ��Y�@E����s�$MB𢂳bà<A��!Us���"O���"ȋ.J��,[��Z�pj��{Ĥ�/��亄m̳7ޠ��F�FMaxR*�z�Xт�b z��V?��=	Q��A����0M��^D�0�$!EEJAZ�O��Pxb�
,U���J��N�v�dQ��7�O@p�f�^Y�,�Y�&5�S��m�`�������%FE�C�	 .��r�G.�E�]A�)rj�W�AF�|�'
dب�
O.D,��%ʏ�$�� �'���2'��3{�*����T��H����pu�-���R��R�霏)iXQ�Dʠ��U��I�Tܘ`IT�Ćc��8�D�&H*x[��όWc!�Ė�]��aR�蓢
S:h��a@�5P�'�\���ooɧ�O���"c�)CtĉQ���S��}�
�'a(Y�`Ԙ>�Ĺ1fM�%d@�5��O�h��Q�g�I���	9$�ɷ�@`��ǆ�zB�=u4���w��[�i��"J�
�b��X�z Y��I~f|��� �1���uk�3u����f��Ë6}����� *��{�:"$���yR��"t�(�Zr灂�.5{��͟�ē��q2Hؚ��S��H�p�I�X�j���k����pE���VdJx��bˇ�Ь�S'�1���׸��~&���킗gwR ��ɔGg:��?4�T�w�O%i�U�G*U+�&Xч�S��HZ�F:�O<ኧ!D~qk1DГI�<��'�\-�ēeӄ�A/��j�LhE+�`�p������,�)+�p��,ج�e��R�4�SN�!o[�)�C�
(TL���g���Ի�LҶ�Ȥ����ȓ���B�'ڐAh1*�.�!j�
h��LȜҦ�Y�B�`�qji�����R���Q�A�0m4T{d�_���ȓo�|a �J,>��ZU)�<H��S�? �(k��
�NK�qi��_0cp�W"O����D#NM+`��_}� �"O���úL@���3gs4mx��>�!G;g����?����6�AZg>Z,�$�`9D�H��@�2���{�GȒ����5" ]�% u���@�g̓c���9��]�"���a/0ͬه�ɽb���yb-/]v����R�3I콁��=$���ْ%y��𑒬В����n�zj!H��<��COV��F/9R�%��P>���Y�	H��Pc�6- ���)D��s0�Ǜ#Q(Y��.9h6��g�<�4�N�@�����.͟��?���Ʉ�@R��n>&B�h[�B.D�x�#a�8i��ݳt@�����$쎔;\��'86����%g{�ϸ'�^,�e��?B��u� fТ+���	��a�P�U�ôZ����S��0Z������6i"|��**:w�}�HH�K�ޥ��"X!����Q�U���O*�J�^�f� pr�#�y�t�	O�ܱ���(ؐO��yr�F�As����(m�Uh�X��S#
4�9���\d`�G��NB�Q�X�sP�V4^h���E���y�M�#Fߜ	2 H��U+�@�&'ܻݨ(r�]��s��v�jb>c��� �L�l�8���+ѽ`ƈ��n%���@�M>�Ƞ"������1D'��//l\�Q��'�yq`T�2�@��o11f.̸��؍�w�W�}Ɋ�'�UI��b���Z�%G*��J�'�Jɚ��C7\��T��\� �v̓J�0�P�O8pE^�$��?��ǊF{b@��.�4�ԩ �)D��٠�ı-Ԕ����$7�V)�-�]ܓI��6��x�ĉ��8Bb�-U�jd��EԎ�yߺZ�0�f�@����C�R4�yR��=~� �S�32��T )�8�yۚ0������/�6��'�8�y2O�r�h+0 ��T�X	�'$�9�y"b��\�P��T��A; ���3�y���)~\��P!Hӿ=�	��"���yR��
]:�@��|�iC��7�y��O�&$.���&�p��"��@�y���,i�xi4�YE�PR o��yB�M�YZ�բ�Ą/%az�Dʁ��yLkL`x��T0Q��D莮�y��f��1�`��: H˳Ğ��y�ӯ�&K��7#�%���y�n��x���y6�2�CZ�y�	υA\~%��arC��J(���y2#9[Ĝ�S���Q5~��u�U%�y�!?�$��diȮK,0��)˂�y�1$<�����$ ��?�y�`�������΋\C�5����y��<�ɡfY��|ܳ�i���y��ڇ-�B��eŁg}~=��դ�y���`�5�ɔ_�0�[��ʬ�y�]�5\��p�ӏHR� ����y��
��%Ag�U�_�99���yB�O�}��X@�~TL5�y�COWN�	�ׇxk�@�m�y2��(Ⱦx�BˈG�}�"�%�y�j�<�$EC��?��� ]��y�_�f~1��ϸ7LrQ"�yrH��'�T�Q�.�,<��@�.�yreϋK�@�Qk
"p�d!㬀��y�G�X��� ��Jjdyf����y�oŬ{�͡�n��Yp�*%��$�y�A�dAq(X$d�8XT��$�y�o�	n�T�䈜8�0d�S/�=�ybdͼ> ��Xva5{tlH�'��y��D�^"x��셛j��p��A��y
� R���-a�ݫ�L�  <9�"O>e)��}%h�J]�
��k�"O�����.pT�
�*�;�z쪵"O��꒳�ŗ+	�Y����7h���ȓ%��zLs�R*ɖ2�Jd�ȓJ]0Mӡ��w�p��d^�d,F�ȓVILԒ�Ν?%���w�%^P=��;Bj�@�f6BŃ%)��r�|4��N��M���,�X9��!��/���ȓ#q�8a�OG9?�ְ��⍹C \h��i2�)��]���X'�Sw�0x�ȓ����'��}�&a�&�]�Q� y��$�}:�)J5vg��9Fd�/�����5�E1$j�Ly8��LA>$����ȓ8�9��@��FP�(�-�O�F1�ȓ
�� ��^�>��l͜��؆ȓ#"ܣr
A�m�x�	��M`�A��v�����F^�E@�xi(�DJ!�� ��$���F������ǌM�*��lb��!�$�3$��(Hۈ3w<�ȓI�����H�\*ȫF���xY�4��^m�ecM���e�e����G�� C���8~N���6�a�����sJXq�Bv��a"N��W��q�ȓW(, ��I�51Vi����4/��,��=K�
� ���J�
e�c`Yh�<��eҁgr,��	yV\E�Ī�a�<I��#��q!.��p����c��^�<���t�(��G���v����i�Z�<at��L�	��l�g���kb��P�<��5
�up��K�n�,Xc�`�<)E�_�h��T:��B9U��
vK�G�<Y�) �>]��b�/K����e�<Q7L��]+n%5�*�Thr�So�<��X� �H�Z��h�yu��Q�<�Uʘ�u0���ܡ,w�X!dW�<I�'�=Y������{��̘4
L�<�d�8C �!�d�`�m]H�<�uꟈO|� ����4��e�D�<���ěE��ă�D�P�$H��#�D�<1�	�=�,p�BL9>O,�A� n�<�����xLt��r퐾6�0����Bn�<9�g߅!����Oâ0x�����j�<9�ūEf��sfے66�yxU�Cn�<1D�Žg%1�2.�o
 ��ˉV�<Q��C�y1��N�3�بwGCL�<I4��D��}�B�P�2�&I�<�W�T?c�lE�@�7F��x���K�<�3�̃et��kpk_�
;Щ�P�R]�<�hh�9���f���Ӡa<�!�ؽwh����#J�)�  `��N�_!���((��[��o��Hq�V�6[!�D�/D���'�,�\P���[�A!���VfM
U�	cc���� G\!���L�ڌ���{@Xä�ʺG_!��[-([�)Y�>�AR-�(i!��3��!^�,�eH��\�!��T�/��]2%�ΑVT���I�r-!��-)Y��P�-�o���e�7)�!򤈸9\�l�7/��L��D�5��- �!򤔡Y$�7�ѕ
��<�����DM!��P�{�̣��O��){��L)/#!�q�(I���2L��ѐ�+C��!�	�W=RH��N���U��уo�!�� D�Q6�'glrȠ�nA
``2��"O�Q��x�r<�!�	�K�Y�G"O��+҈ڷ'~��1T��:ms��
�"O^|���?#K������o�}��"O|��Q,"����"��(�a�0"Of�a1�I,"���PgS�x;"O�ŉ�a�7u}��S��׻]�T,�6"O�m"`̆nVbXbpM�:�6`��"Or]�&L�5��l�BF�F��CW"O�Y�H� Z���f�F49���c�"Ou�n7}n�уގ9����1"OX��O��_�L�"3b�=q�(���"O^��dQ+.PB��2$K��P�"Ol�͇�_$��d����4	�"O�afJ��<��J�-�Z�k�"O6I��_3OJ��ХK �p����"O��OF�L��a!�����a"O(5���]X����?N�,�+�"O�]�7�Ȇ8.�B�/�;]��I�V"OJ(��oX�Ti@5���K
	�Q�"O���Q�J�n���[9 ��)��"Oj�)Qh7e���[0��\�\I{�"O0D�#o�9>*�:�K]�9z2��"O��3D��Edp��7jA2t�,;D"Om�&�[��PrD#ɫrQ�y�A"Ov�����0C��
N�H3"O:�:�.[��H��=]%�YY�"O�i�	O�4��YƩL0Lܣ�"O`��(ʈ u��zՉ�:`H�g"OЌQ��.b�|��,0x,j�"O~I�Cᇽͨ��莕(8�i�"O���V�H<��bQ��,O��Xz�"O��y�.�����=f��P�"O�`F�Ա���U���U�B"O���iل]G\m��&�uK `cq"O��C��0(���dC�F2*���"O�� �.GG#viQc��kޖi�f"O��u��7)J$�V��K�|�P "O�q;����/Տ7�©B�"OhU��҈ l�1��Y@�^���"O���ل�q���9�L�	w"O����	+K&�}X��Ж�@9�"O$= �
,C#�ɪ�P���	��!RC�`w0�|�'0���×�{�ԑ�f�I�9�Le �'U�e���
=H�PU.�yٴa4�7+��T���!<.-PaM�26LB�˶�˷ :���	4gk���7��W��
�Ƞ�z�ڡHD����LF�i!�䄺Kt2�-W�8lC0�E,0W�' ~�6�	[dɧ�Or��{-U��^��p��"+�dA�	�'i��N�9<|�G&@��bJ1�P�I�|5��L<)"E�$@:�w�Ό\< �rLIH<����v�ܹa�$_-m#��{3�=G���8�+��p?i&HԿ��u��HR�0�s�J\X���d��>m�O\�Ys���}�"�ej��)Bd�W"O�{���~h^����f Z���x㑤
�^��g�|�����WV�]BfI��	��[c�6�y��$3�,��4�T=?�<|Y1�
���L&�tqA	�����K.�E�4斑t�|��QZ��Ɠ)���w�P� �2�qC�"0!ڍ�gL�x0��	0��Ec �6@���`	�e����͐rs8OV�£���Xl��5�˒|E򨰀"O�h� W1zmJ�:8�E	�"Oʜ(��BCK��p.�aw"O�r��ʪ]D0K�jB/$08�w"O� �����D�LqP��i��amd�"O������B؂<iW�Cu@�8�1"O����P΄xb�I�5�qɔ"O �q1b�~��B�&y+���!"O��8�.��q�3*��"O���Sǝ&�N�����%��mh�"O& {��ٮ4��#b?�ja�'�>Ag���:}.��?���%���"��$�K�\a:�9PK2D����n�-;?\\�S������G�RM��'���e�g�:7�IPa�����X�lM,����I;2�U�PMPb۞xҌڳG4�܈������@��x���R)b������C��q7�*�J��u��bW�WQ 5�VT>My�ǏYN:�ZU@gV(�R)D���4��%xm��8�T�Ӫ�<�孀 Ht�0�oͪhw�?mCqJ`��(���&,��Ѵ;D�ԉ�!I�?�xy"Fίf����5dZ�-���'pt)�EmD�'��ϸ'I�(@�O�6��4�X�|�4X��oL�  �,��W��Ҧ�N��%[�f��-ú�%a�)o�}2�T\dd��P	^8#,�1�Ɉ���Ot��U#B&~Q���Tg�f����h|ш� �3�~�����y�,3-��	�C(N	�3C������, d��u`%G����$5�� 4��0%i��y���҂��C
�(��2j�\�҄�1]��RGɫ{Pfc>c��&D��)�\)H+i�t`�5��FDP�%wJ��R(^��x�zuaET�6�
ҧ��/����D[�y<Xdz��@+�D9wcMt�ax�b�^T݀�d�y��ch*�pˍ ,���d� 4�!�J^�������d�n,*Q�M��1���p"����S�'7+�]��)�5Ly 	���>�L��GQ�e��dֆR��u�釜u*z�{�N�
�c?O����)�.}W����A/k�,h!"OnayD���:aaД��+����"O��@�͞<���⍒�<�p�"O$�2�)o*��1�FE�X��"OR��.�<��,�r@�Q����"OHc�� 'A$�	�*�pؼ ��"On�)5�Z_����7N�.%��"OZ �0*äDⓦK�ZJTU"O`5�p^�yƢ�H&&��i
���V"O�mP���,q��S��{��HR�"O�8��.��*��x��M�U�Ա�"O@0� '�d�j���6F�NX�w"OD����_����e]�XԈ"*OP0ʖ-S�l8,�p�׵k�=��'e���D*��[EpE�ѥ�:P�d���'���J1��Xz5c��:���'�T��DP/W���@��~ ���'���ɥ@�6[X ���S�q��:�'�(	�F��9$ �b�A7`��x�'[$�H��_����׮βb"��
�'Q�m�e���|b�&@ٙ+4TT�
�'� �j"��
0`:�ʖ�X-3$Qs�'�V�c��6F�z0�˄)��r�'@f�V��YC�]��&=&�K
�'�=�')XD�fQ���[:�֥		�'�J�Ǡ�5'���de� S>�؉�'�f����wՐ-�%�Ķ�F��'��� �g�9�x��#O
y����''*��&��_�hY�� q�d���'\�9���5Dpy�Gx-�
�'c^�5��X���	�F�<8��'ܴY�F�P4��r��+<�$D��'n�8Á��Ca��`Q�%�⑲
�' RLB��V+<�����L�	�lB
��� �1*�� S�h��%`Q�YX�1��"O&����`c�����m�m��?D�`ZfDO�#�L�f���UL/D��k�@�O��:��o���W�)D��Z6��>�H�	TB]* �`��bH!D����֟m���4W�$���8D� �V�ڭtY^u�Wb�3_,P@*D���-̊�̰�Î�xz�5(b�<D�t[N�:Ү@)q��7����i9D��2EE��/����C��3V~TH��6D��*�i�%f�� �V'��K�<<j��1D�D�}x��qmZ�n���xV�5D�\���D�,�T��WĎ��ԫP"3D��dƏ*-�����,sf��GK0D�쓱"�4Sب���\T����2D��¦_*G��D�Ɲ�3��\o?D�(���ք`�.�[@��-i�6(���<D��) dQ*�~!s�K�{�u�#J=D�� ���cs^�;��D�t����Gk?D��`+�An�����b�t��%9D���VEך?=� 
`���8�p�0%�4D��H�)6a��m�E�Ћ`
��8C�)D�X(�F�3+	 ���b�rS�$D��zdcگ"�ʁ�,�AF�Z��%D��zjW�i��7#�:@������!D���,Z��� �`/�5 ��I!N>D�L2���.�L�У���}�����E!D�T��D݉ͦ�aMM�(Atɂ�d<D� c���ED4b@��? �1�*O��
�k^�R/$���X<u(�+�"O�D�@�"9e̸���5�Q��yR �84��Tb�h»v,
���)ҝ�yҩe؜3�o�n�D�j&C���'�X�ƃ��=�fY!�@L:d�(Q�ƙ|BN"A(d�i&�Zg����V���s��(�^=�PlT5|��P��1��s��'�ў�~ڐ�@�rUi��+WT��D�\�'ra����'����!_�2F�Yc�K���'�ў�O��0���R�sg��U-�8�V��O>����)�e�2IJġ��n�+��3��I��Y~Zw!��Eb��,ۈ-I@u#K�G�b����֏ʰ�Ђd��8R+�o?E��&�Ӳ���?�9R�*ۿFo`�ɬH���l���O�����e��fu�ĹrȂz�4�p��=D�Q���d��!Ȓ~6��r k��V|nؔ�x� �H���O
6(���̔lxxE�J�9�^�8�O��h����^�����`�n��ՆSeZ�ܨ&!lӠ5�*O8(�*O�?M��D�ڨ�� S���(i��Dy�&By�+Z���'2��I�nQzv�8�G�5��''��EyJ|�R�$�������{H2Ī k�J�I�N�Q�b?�3p�9�J=���&
�2�Jc��>QF��M������F*)�V!���A5�)P�N�H9`��rIUR?��O���~������c)ܺo̬H[��6{�<,��K��yk�'�����L"#�ϕ.UF���*��h�^0����p���S�l��aі��$ypׄP�i�O&�=�}��- [`t�A`$v
���	Zy��)ʧ�@�P�	Z�ȑ)�dMU��p��L������F�ۥ8�^y`a�փc2�-��	Z>��v���� �G�%���J'�&�	㦡Gx�'t�j��f��d��H�ߑ��@����!j��C䉐�<��늼9��ę� ��MB�C�I�n���׫�X;~<��יO�C�1�Բ��cX��Q�S�\�dC�	�8U��0P!ōu����͘w,�B�I�6�Nq���P.k��b��FB�I#Z���7i[�v����g�-64B�)� L�,�w��{&	O���"OB�y6#	�Љk��4]�����"O��4��
d"x�I�EX��p�"ON ��@Ҥ�T4i��J`����"O.�� -�$)\�6 ­Kz�A"O*�i��S�B��d��+ɸ�ɒ"O���3*�&��H#�-G	��Zt"O��+j@+J��P7� �!"O�hAS�W޳B��	�{�<����}}<�����8�F�"Q��t�<�%���/GV�C��R3",�$3�KE�<)c��
OL�:�Ɉ�,�:8ɑ.LA�<iA�������vI(�B��q�<�E͈<DN��G�K���xv�f�<�U`�>X�.a���M�H�H�Ma�<I��K�/�`�X�+<>����D�\�<y$� raQ5\#`�u�U&@�<��O�\�6ia��J�d�n�;7��g�<1�0R�~��s�o�$�����`�<)�ȗ��M�cJ�?DiK��R�<Ap��ebt)`@mL�Eմ0s2-�O�<SdG�l�H@�8.ꡉ��F�<I` 5�.�Y҃V�>vb�4�[L�<q��˰�����`��n<�U���C�<IujK��ȴ�Fč�~�,��H�<I�-X/;�40�Ā�1"���FD�<I�^�i�
y�w&��aT��
�$E}�<�u�QS.l�0*˧5@�*��s�<��_�<����&B�|�a�jI[�<1��2f��Y9�H��U�ȉ	�f�K�<q��[�/| �3�� CJ��r�H�<Y��%H������"t� Mʇ��G�<��`��k<�I�6�a���2��Z�<I�7E�Q;��wf(ç�q�<)2�_<k�2%�F�
k<lô*Dl�<1T��65���IE)Q�)���g�<��IIW����(��� Tf�<1��'#���2�惇Q%���h�<)�ÔHG|ܳt��j��$*�f�<���MS!͛�<VQd]'��W<���!+���TCΗu��S҃ޅ�L��=�<]��cň	�^��&@�0ưE��mb(�r��kyVq��F�M��P��+`0K�)F�?j����!��iȢ��ȓW���YQ�Ӣ:��<k�Lt����lN|}Q���=kj�"�'�'Sf͇��`�3�a�/%�d�:@��#�܅�g��s-���¥��/Ey5�0�ȓ(3���@�uL"D�f�>;U���y/P��ukW�h�n��4c�uH�݄ȓW���w�]��:��r�͛�VX��f!�P���V�%�P��� 0���ȓyoP9�Q��\nn܉BF�0)�5��9�iꁫ��^ܤ�4/�2[Τ��ȓH�1��BJ�aY�@[�☇�H�Ԭ�v��!s����F�E�|͇ȓQ"ȓ�K�p.���B��-x�\�ȓ�6n�&��K�U^���Vk�<)�g���t����k���"���l�<!��](>/xT��HP >��dL�j�<i�Ɏ~����;@} ��3�i�<Y) �D��y`��9H��E
�y�<ak��]6�@��V�l�Z�I�D�w�<ٶM�.*~X�8�,ώ8ʲ�Q�Lq�<� ���B�&~z4p�G�
�dUv"OJ�2q�W�!�B���\D�x@"O&�zrM�&�.R��Y�r+h�Q"OR�AP��\�8Qʠl-T��"O�9�6�
`�ْܑ� :8sF��"O�ī�B]�/�<(�8\Z���&"O��BW��l���`�5#@�i��"O��&%M>~��(a�Ê4008I"O� y!��D�b���N�J��pp"O��@��<���s�G���43�"Ol�䎁j�.勅C�v�z���"O&��lE7-��@�L�E�T8!�"O�Xb�mW!^�y����]��(�"Op�BaL��Ia�@�lU#-D�S�"O yQ�FG�j{��ҥaC�2��"O�y: �B�6�ThQ�o-#"�:""OX]'&�t�b-�7nI�1�"$"O�-��zBT�����"��x#�"O�a���)v���%�̿'�h���"O��G9l�CS����@���"O�q�E	-��P9���720 "O ��X�Za@ "B�$&XБf"O*��F���-������'P���"O���X�6�"���0����"OZm�������a/�!Ƃĳ0"O��0��<GwT܂�n��^��0�"O�Q)�"߄�V:޶�;!D	�!�s�\�2��R�����(�14u!���%Q���Zp���vKJ0y���0�Py��W�&^fM��h7O/�i9���y鞓T�"�0a�S�ޅ�7LW.�y2��Ӕ�I@�0;d�:�i��y�&E"nY|	����0ϰ�Y5/�)�yR�A�Aq�P{��]�V䲝�`�yȄ�x ��20,�� ��ht�y�O�7'�Đ02���с�@���y���X�$Sd*�w�D�(�o�y�JP��$��El����-�1�yҪH��Hjfk�U��O�y�DK*# 0㒍X�9��"�;�y�Ċ�}ܰ�8�͓�"aؑ�y��#.����� �t�Y��C�*�yҩ_�s��t���	q�z�{�(��y#�<u]6i�� ��U��L��yb��!�X��v�~��s�4�yB�ʅ `9���|R��Z ��yRC��tVD*�$�)L�p���LŽ�y����%�ǸB4�t��$6�yr'X�Zl��w/r�R-=�HB�'x��S�;z�<��ڛ0DHl��'$M�5�̅Oz��JA�לtP��	�'x)��ǅc�� ���L"��pX	�'
d!��T�,��aE7^(�'�T�7Ś�	�Ij��7M��b�'TjU�1�^?U�Lܙ#�X�Kr"q��'��P��nU� ��̱���?�4��'@,�
��P�i�Pɐ�4@��X��'4v�j�/� h��U���8��X��'c<��׌�0�D$脀�2-l��	�'v(��$lϊD~V�q��R�$� 	�'.�p��V�Z;t R`��2���'%�m�`�ќG�&Qrd�\��u{�'�^�jp%O�H��`Ď�bĸ�	�'GV��`gO�n��q�x�4ͩ��� .�!��=X���I�g�E�B�%"O����N-~��1��ڪ Lv��"O2�wi��D���f�@0��#"O�Y�� 5����w��!$��8a"O��p��� �A�ɓfg���A"O�8D�u�9�J=_�8�"Ozh r&2>X�IF��z��8"O��B��g��'�_��@��"O�q���l��@I�Y��u�A"O�9KqŐ_V��B�¾	��ԩ!"Or�v�C�iC�QU%[�JŴ4P�"O&��0đ�x�F���D_�&�h�B"O���#M�"$���*��1"Oz�*ҩ���8(��`ݢ��Q"O����	H�-�~_�-�"O~�c�IpVZe@��OY8Q�"O�U��1cpY���H44>���s"O��c�R=r�:��׮RA�\� "O���0�T"0�Z"����Jrl�"O���&�r�����M�C�0`K�"OL���mbP���/	��@�A"O6�떷<95:���*�2�*b"OI��/ƾ�"=���P�'�*�`"ON�8r��4U���*�mK�v۪�!"Of���%Up L����d���"O,�8t���>�v��ΘC�BŰ�"O�=YF)���tuHT�]�F����"O���fB�%��p!���	A�����"O��*�M��-~���ߑ���Jg"OP��6kͣo<�����Gs�hXU"O�x���c��틠�Ȗq�P�b"OrM��Ӵ���Fћh,m�d"O�9Q�Ο�t �! f�<6wVhQ1"O��1U�IY����!��E���iw�(D�l���ˉWt�X�F�q	XP��%D�l�f"��O�����"� l5b�.D�ܢ���<.p��1�E�QNT", B�	�r�R	`�L��3��Go���C�I�^v��XOX��j�QqT,C��(3�p`R��p�hQ�Ͽ�C�I�KC2����͛1C�@k�i&X
C�Ʉu�$I+KM�.��;pʂ'��C䉘8��=���ϗ~�Պ!.��i��B�	�}�){�c�ZP�P�#ˏyZ�B�	jA�ԛ�Dܗf���D≿.^�B���Z�@��̄v���0�/�Z]�B�	��B-c���1�	�c��,�DB�I�M���ڈU@p�xTk�"|C�	PEN1sK�-w%��z���?m"C�o�L�M��BV���D��c�C��#d��@oT�dhP�g�'V�C�:Je�0�w�'#fH�I$� PA�C�#%txytj\������?6!�䜒 �˅�E�OP��F��;C!�DY47����� uԉ�ūÔ=3!�Ą R�= p�F2B&>��a��E !�D^"/lɃ��(C�T8�&(+!�Y�b��t��&(Ĉr󄉞|!��ZXv|�Q� �5&ځ�#B��!���,��<q�H�$"$�"7LI�P�!��K$L`��:�(�7�J'
!��^�8L�t tl[�tݢv`�B"O	a�   �\   �  -  t#  �.  �9  �D  �N  �Y  �c  /j  sp  �v    -�  ��  �  ,�  m�  ��  #�  y�  ,�   `� u�	����Zv)C�'ll\�0�Kz+�D������b�vgى�y���yfY$E+�D@�,L�]��
�I[2kƠʤl�%�걂��<�,8@�e��"��n�5v$�I5a^��i�6s�ƥ�����$n�`a��))x� ��m	��招�f|@��ǁ�$��]�ޝ��'�?�a�_? Ôr��$Z����6m� =8X�(BR�2��Vl\�9"7�W*6K����O��D�O���bt��`텒xU0e@A�
3a����O�m��L�'���,�r�'��I|��a��Z p�N���A\�52�'�7��O���O*��
?���䚁��B?H~x�15ɓL���YC�@��G���yr��,�d��.9��O��% <=�V �5��B�d H��Ԃ�>��'r�O,`�)D6�ƅ(j�蛡�Q�v���PaP 4L(� ��O~aoZǟ|��ɟL�	�?���y�9��<�tÁ'È1�UmSOn�f�'�\�5sӪ�oڃ�M����ɓ)�~��ߴb�� 3��X7���R�ڢ<�����L�u�.���H�v-�SM~���Y�d�:^�D����lͬ%�´�&�t��1���^�LY�M��x�C���M�i+�6-�
��'�0��df�8{�l��(��3Jh]��:A>��o�� � �z#��+��<Ić�q5�@O�@nH)�f�i��7�T��9���+q� �0��
�Gx`� {K2]�A�C�@s�4k����~�>��Ҡ�!4Y�=:��U#��܃��X-U:���$L֙�X�A���^�j�Õ:J�t��э�ۦ]�ݴ+��&hݜgJ�D�&�ͳ9�x�2����*�z�.��$]ʠg�&q��0�r��ě2���uT�3$�#�`U�&B�O�⟸��
�S�b h���9p���u�G�X�q8���������?�h�NC�q,��5F埔��'�?+hH�w���@aA������0>��Iӟd�	? g�h ŗ�:��� �4�y��H`W�=�"E�3d�|}��ع�0<	�T9EP�äL����$�0�( ��:V>��F��-:�axB����wy��xWx���CN2����?���?	M>���?�,O��$Z-}�*��g�%2��W�B����O>��,��&�O��9O�I�ҟ�".Q�Q���"�B�ʝPVh�O�MU���g�i��������M�-0(���}D����l�O���Hx/����b��\m��Kϴ DZt������$��i+�^�Y�x�(�ޅR���-�:qz��դ���㘩Y6`}�XwȪ 	wh1N+���F<;���YT�%|ɤMr��I���޴K�bNi��5F��5�
Q1����d{���)�H��E�'��O���bL�_�|k� Xe�����L�hOd�	Ҧ�ش�?�3�i5��'zz��sw��2F�xt����v�r�'��Ʌ��	��ݟ��I��'{E�W������ɐ2 �����}�& �p�� �4Y�@?/���?�Ѡ�x�/-�4��N�"�0��@2n*�d�3���]�,�*��М��pC���s�)W<	S�y�?���p�Aͤw��8,7#,���ϻ{��.�<1Qɞşl�@�L>� �X$�2����"�@�e��?�����D�O��?�'<��YR��-_���b��89��Z-OJmڶ�M{K>�'�2/O� �᎑(� ���/	��c�WP��'R�'��IG�D5�P\)�ɗP��U�
 ^|�RgL�x�R�8P�C�Q0tca[4S8D~�ƈ�,p�{u$[���z@i�1H��hf�A%Z@�m�橙45�Z��7�ړ_�"Zܓ	̵�dh^	*
��s�R�J4sA��ßT��4Pґ���?ٴc	m�H%�&�PD��
%��?���?1���K�	�k�ח�K���W�|��w�`$o�vyB�Ԁb|��?!���;h�޸�wa4/�"t��D�?��t����?���h�  2.�*��tb�?YlʅCP�|kR)�bnS�i��!��FV�#?1�,O�A�4 I�7m>��q)O>|b(�EM�4A�*	�剆�l�X
.a���<�ɰj�4���צ�۴�?���&����.�:��������$�O�D�OL����H�̓�H�9p� ��di� n1O"�=�O�6�Q ��iy0��9"��W�X��.�lZky"N=r��uP4�'��Q>��u��;w� )M���]_i��V����0�0q`�DP�_ �;'�($ժ`�Q�k~��O�|����E�f``!�G܋W�Z� ����q	�!#κ5��'ö'��W@��4�lV�X{8`�S�0i��Ӄ�#Т���
�@���G�U����M����$��߿(T1��7j!�Tc4���Y��'�|��'6BY�H�Q%lD}���A�`r��sʖ���OjQ��즥�Ɏ�M��A�^X��ҿ)*����E'2D��i�R�'��j��f�Pٲ�'��'��2���y8�Q�Ř�|�+��7o$�E��S�,I ��r�S�T{�S�?�pc�xr�ĭ.��ŀŠ��Y��l@j���\��	_li
;�H��=���)CH����:9�Zu�h��Kき�S�>(����B�.=�P����QSZ�p1D��O�b>��O�Ćdk�%C��4�¤�ۡi6��D�O����O��d:�3}�狘$WRH�B�F�z�	&A��D�̦��4�?Ad�iF��O��tX>�8�
O5����_���
��6�*�z�/~������ɲ�uw�'l��'Z�s*ܤGE$�BGC]�����[-�{��N�11<m�eL��D~���:,tf��qD͉#w@���&r�4�@B-7X�Ȩ�P,��T	mӨȉ�dŃ)G�O�ĉ6���6q�qc�,PT6�����@�L{�\DzB�I�`��Q�t�OCOl��/E���d8���O�4b� b!�'<eR��!%�%��\�UI)�D�Ȧ	�ٴ����j~��l�ß$͓%�P�"��k�2�pJܓ8��UD{B�'�,����8,�,/>-��"�� �����k�v��`�C)�.-�"AT<Lʍ򄉾k�6�c.������%=*e)�������v% 9C�T90dOߍ�
�����ڸ'�j�!��_��'�<i�#�1g��d¤�݉J�,�q��{�O��O�H��C[8J,�	�"#� p4�p �'�6M]�7}�)@�#��OQT��OQ�ބoYy�'׍a�6M�O�˓��i�O�)��-f(	���1E%ք`�F�O����8���W�@ g	h���oW'䝰�oL�rK�S:C;h�B�-]�N���d�ʪ�Nh�'��:�+Q�ES�U�1�c�h�����#:��X%���t��8���w�e[
p��I���D;7��sӾ�G�d8�d�s� )I2X
g�Ն1t�M{�z>���fڕJ�EZ���z(�<�S�:ړ�?a�idb7� �dZ�D���B?���{Aj�!٘o��$�'[(���O��'�T�  ���^� 	�E���,�4O�5Z@��#c�3�]`!�{���OA�&	��<u��'�\�
�nߎw4J�!a�� r��)�Ɖ߱'��m��Y)`I �i��Xϴ=��Y>h7��<^�b�]�Eyl��ƙZ����&�n����d��t���O��3��V"���C��c�4(84��3��,G{J?y�Y �cĕe�,t(�@�>!в�d�ONUn���M�M>ͧ�*)O���E�-���S���,a��R��D�����)�OB���Ol�ퟺ���O:�S>4�$�s`��9�.��P'�4U�.x�vϟ
'x��M =U��Z�����Ol�R�"!���Q��R���q���B F����0��?,�5A�T�A��c�91�h9a�{r�rZ|P����[��;6Fp�C��O��=��OyʢN%v�hTHE�Υwo����"O�Cb -T6����81�A9!�|Jh�`��<!�bN�\C���'�2#��C��8+�@�U�F��f" ���'h��:E�'+��'�`�Z��;h��,��;�HmXW(*?�.�S�nI��y1u��-]�<G~RD�Fk0Q��7#v�!q��N;�i�6(G�-��Ǉ��h1����P�r(y!&�wܓz:���	��M[%\�d�0���w
����ՠ�D��<��6�S�'���A���~�ԑ���X�jbŇ����M[��4n�Ph��L�ʩ	�ǬE���T�`�����M3��?�,��|���O������
�����Q�=k���O����/z���d�<����>!2g��W�œ�φ�f}
]�`J�T~���$��&�!hG��&�0J��H#��7(_a�`�r)�'��}���y%�V(�'���-G�$��� �)V�TWz3�F����'2ў�O��P�Q�R�ZM;tg@� s����d�����4��O_���@H"BT�l���ˈfPC�i���')�n�[n�����'��'�"6�X���B��$ɶޗq�&�K#"I��y��'jD�h�m« K�3�|�B%
ԯ> 7�v��0�A��.��s� E:��ތA��(��TN�g�A�h��K-\�p�S�i��4"���G�����g�#
�U���4�1����0���?���9?y�'�*��a�j�bS/ԖLyd�}*�6�d�F�DҦM�O��S>y�4���g�xU�� �g�H
�$V=U��@w%՟<�	����	�u��'R�'���h1���p98����b�� p��3�>ѣ�:�O�u�h�n� X)5V�����h�j	�w�˚z ^SCE)ML&��	�`��M`K0F���a	7l�p�#�.�O`�mZ��HO���$�?�Vݸe��F<�gFٞ"�(C�	7O� ���J�pA@����*yi�D
ڦI͓�M�ƺi�S�d���ݴ�?	�'?d��%kF�⤡Y/Z<�B\������OV��z>��2G��[	E��ȹwi�VLY�Z���k�+��J��0d���#�3|�Q�,�����UT�nӈT*���3GHEq�c�G������'M�||��X�#R�����ճ��!Q����	�M�r\�0⇄�ln�`G�'h���Zū6��9�O�esp+@�r(YQ�͐�%�.�)�T�D�'�ў��M�΅<8;�AG�]vrY(�H�#��f[���I��M[����D�|R�����1�08�fܓU"�n[�e����?��ˡeWH�����z��er`�_-��X2��UY�ąQ$,���]+%5@��%��6��I+`:�H˒�̡���ϮGt�4�"H�)�d��@��?�����S�(�d��%l+?1ԧ��ȡٴ->E�4��邳�H?r*��	0m�{�4#�|�'y�'?��	�X��QУ��*v�����%'���<���sc�	wy�3�=����O�p�'L������'��'��$��Բ�'�"�'��2�ʐ@ЮX�zmCP��y4d '�Q�4
��-�A��k,Q,1�p�%���P?��]R$F�/�����Ӗ�:A��ɖ�u��an�}�q9c�~r7�\�w����;#x-�sfS{D�1�逅aH��IW~����m��$G{�l;h�FG�E��� �0m!�U.~lhh���;$�4�KBE	剈�HO�I�O�ʓ/��U�g�\"$a���&��S��c�5����?I��?qw[?Y�	ҟ,B�#��]�r��2-�:�pGZ4Tač1��ҭ�f��	ߓ6��A� 
@��.ʔL�D)S�+<����	�� p��+e�8�{ kf�'lJ� լM�l&�@ʃ ^�F  e��'�%�?�Q�i�7m�Oh˓�?���?�̟j��6K(X5Lc�&A�iC�I{!�'�O�=`�D@�f���݂X��
G�|�bӰdoYy�`�PB"6��O<�I�M y#�mȅ���ǎ�Er��$�<����?��O��z!珥MG�yȠm��"L��8��נ�`�	$恐|Z��r@זZ���[2��G�'�d�iw`�K<R��g[�h�R��AC��u+@CfJ��L�>	y���"Q��l%�/d�,�YG�|BD���?��i\˓}|��&҈"(���1g�b$'�@G{���!#�Aè�+�������Q��O\�=�'&͛6i��I��[�Ɉ�Z�*ɍ!?�66ͱ<�7��5Fo���'R�Z>�C�o�`�C��1z�r���i�Bn�T�LꟘ��6���+ Ȟ"�^0���O��M�+�(ʧS���b%��,G�v�s��R> �Od%C��$	���-�^q�&�&ڧq ؙ֡��=��m�0� ]f�8�'~����t���>ҧ�����k��q4�GU9z�����<1��$;r)N��!�J��;r*�%�џ��޴\���针V�5��b؟<����拮.l�7��OZ���O�!��,���D�O����O���"d���V��Ih�\O�-B�C�B:^�(�ׁ��0d�L�b�)�ӡ"訁�O�(1G)_;� e�1���+5��@�P�*����ތ&�}�B3@�L?��5�˪+��8�"f�E�L�8��0�L���m���L�)D�O�3�D 
P���B�O�X;�  \�C�	6d�}C��7p�Y��^ @��I鑞�ܟ��'������#*�8�3WH۹F��qV�'���˒�'�B�'���~����?����
F��i�L�WO\�x"�@h2L�#W��r�Y�"��'�"@Ag�/�;���1�CD�:�cpB��w����6 �2;�f���@�lP�˗6]q6��0��W�z�BK>� �\x_0��&A�`�u�38	����n�(�4�?.O Ь���D�<��B:�F�ʦgP�{��u�C����O�9؊{��i����'�� o/|��6����W�	�8��4�?	˟���c�~"�W�d Uf��h�Y�S+L�t����?���I��?�����T���|`@Ie��:pݬd�&cA�d��#��͟P���#�e؊G��=�sh<�<  /̆��1��>y���'R6�A	D�}JN���
��_S����A�)��҄�:�	�KSD���O�&6rD��UQp��h� b��'����ɞ;�:q���;S"��4��/8��d��
ǁ@����F��u���O2�#
�Tr��?�����IJ�\B�$�=?$���#��B!��A!#�&}�H�D�Or�RW�U#���&*�&7tU�w$����?Yۡ �%u>�i�Q�V-��c��!?Qp%Z7m~b�1Ą�]WTD��H
 _J3A�@R�ӝfy�H)բ26l:�.Y�c��3glT��ןhF��0O<���k�#fv���@*rX��S"O�1H�)
�~p�I�+_�� ��	�h�m;�	A�Y��H�=>���f�'�"�'�bd�Mz��Rv�'��'Vb=��t�jF3��t`2�Z�!Z�$��A?zԾ���,
�u�1���|�1�
�&�h!�n�z>h��H�ސ�	s���i��_�]0R��j������~jaEU� ��λb3X�y����?�&%���{PP��z~r�	��?���hO���V��5���ӵ'�5&��� /D������v-�T�Uݕ��Lv(�<i��i>��	Yy���7`��dME�MJv����3A����B��7J��'9��'b������	֟�����!��JU'X�̱��bG�!C1H:!ڞ�
ߓ3�jS�Z�y ���Qi�'o����63"h�&eG�/����w,A�f�J��	�'�n<��k<������^�;�h�0WC�OV�mZ��HO�#<���B�p2v���"fu;�/EڟX��Ey��'N�s�4�<��K<qb8+B�����&M�ӟ�1ٴ�?)d�i��6m�|z��K�N7�f�'r��-p��z"�H�S�\Ѥ�� U�'�th���'�R3��]�ˊ=1h�q�_0e.��ޙ|ߦ�k��:2{����g_U"0�?��F��P��FɹW���	��=h6�
�A\R�����s�h����T_N��B;�I. 'J���OP�.P�ٲgO�ᮔ�#��$gj(%���IU����ujͅ��2ꌆYlH
 �*��F���	���d+ԋ�.g2�M�!]�x�&��G�ORʓk�Pk�iH��'���+%�$���*sD�*�(ʐ	t洙&*ޕ$���'�2�ʆ	�5�dGC-{Tr�S�d�?5�E�À-��D�L�\Z�T�Ь'?)�M�l�v�����V������0�u��$Ƌ	���c��.Y��J ����%3[k6����*�-�7n���C� 4K�BB�	
a��؆CU��萍U�Bx�43���O��Gzb�����ǌ)cc����W/#7m�O����O!cDeu"B�$�O�d�O~�+-�����.+�4��F�LB�X��bI�<��qd	 ��˥��|��'1JNOjȇ�^�gXL�!��V<A�Lt����J��J�G��pn,�S4/D����QL?���.��F��=� DHx0C\%TZ�3pB�,���'gd���'�`AX���?)��?y@L�B�����7�fJ�F��?q��?���?qN~�=a�ݼ+�
�uB�M&4i��_���������4�?I0�i���O��W>i��ЩMΤ��֩Z!Ա����3E��m�B��۟(��ԟ|���?�������'m�y��١$�ZT!���PҢ=�G��sС{Qkd5:H)6���M㑟,��)��W���E��<�9�O�jvH&��:w� �ق��S�&pȢ&I�`!@,�$�Ĕ�������,Y��SeK�q�r�J��'���s�'ȨT�7K��>�]{�cJ�Aq���'K@����D�>ӌ��)�@���M>a�i�BZ���Ŭ���d�O"�����%�T���ɂH��L;���Oh��=r�4���O����.@"f�Mq�ܐJ��S�-�����YT%fڠ�*B�,3���s�'�M�Ώ��t��.�#N��Se�ֿ]r1q!AL!W��U��#T`�j="���O�'+���� ��6mnӈ�	���S��]�z��G�EB��?���䓴�*��#F���,�ƭ���#�&�S��p�.��i�-I��D�F�?G��m�KD����>�M���"�?��?!����I�-�?I��7�L�b�b>=�Y��+�?y�^|�1�"%�\�X�CD��#��@�&��?]�O�>�T ��t��i]�K#F�3�OkGC�z���+2��j�@pJ�w��8H���8!� �s5IБo�~���zSA��Fc���Odq���'��S�<���i32�RH
�R��A�<	k��t���ۑs��
&K��'�R�}j$j�:b9i�`J�
/� �c�	����O��d[�:U2e����O�d�O���hޭj�[�$�h��@o��`?�
pD>-\�oZ͟�a �ɈqsF(��(O�s)�qҼQfC
����1��
��g�߁[Y��(��F5�1�b%��ÆoD1����TK:
��G-�����4�?�����?	��,O:��+~�f)0�4��K�36�����O���$ �P\-ɗ�Ei�֍`�+��j �Ӧ��Z�4�䓕��'��˞b*�9�HT�W��hC��FH��B�i1z���?���?qS��P���O��S�n+��"��%1Ԯ� TB˒�2���#G-\F�bH��zS~���?��!��-^����d����
'x|>�x5�&Qd)Tʀ�+�`ȋ����`��k� �t��b��K��P�J68\�aK�#
^�"C��0L��GD�� `��$$m��&!�" L�+&?D�$�+�8�`��c	0V*����=���Ϧ=%��R����D�O��A��Q�V����,l(;UJ�O\���sQv�$�Ov��Gh�,9&��7Uu2�ZVHN ��キʚcE��q��5I�}��o���Op�R�)�,1��K�n�IJ�a�U%�|O��b�%��Bg�dRǦ�*A������ԯ/*�q��{b�ח�?IԷit�7��O@|c�M�3��9:�רS����+�<��������۟h�P���,PԀ�R혱�1O֢=�O9�7��s�lU�M�&!Q��r��\'dbm�ry��'���?A)� d����O~�����).�Yg�[$*�!���O��� �L^�ۡ�+D�����̰3p�4`�O�哙Z�sAa�#%�IS���)М��' �D
�CatF�I7E�{Kh a��"i>*�0��oD��,ٓ1N�tC҄��3d��X����IOZRFl�@�m�ٟ�O�Аq�:�qؕ ӻG�X���Y`��jA�'�؟����>	��o��A��CEQCpAi��Q%@��T#�A����'����'/D맨��O�!st����t�+֊U�#Լ��EGZ�E��䟐��(xS�rWO����	���	��ԑQ�Z���9c��㧯�8 ���x�O*�Ppb�J;���qO�IG�9cgH�����E�HL�W��@zfK�P<@�`�m�*�Vc>M������ѥi���]�v~
C�)Id7-�Ey�#P�?a�'���|��0>Y��tᓛf�����ߒZj�T��Iߟ4E��59���"�)OD���Y(+W��'%�6�����5�M�)���)�|��oD��,�)��U"(�lP R��(�yX�M�?9���?���"��?ٚO[p�q��NsF$Hv��}�]�a��D0dRa@V�I ���bџP����ZT�cc	~���p���9�� �\t��7�N��GIQ�:z�] ��D�=��!�-��m��@��\%�T���'���H�'����D���a�B�"��TH��'~AjƊC���P�(R�x��e�M>��i�2Z����D���)�O�	�f��l%�t#�e�lR�����OP�$_SN�d�Oz�'[Q ف3'I|lm�foZ)h!p��%�k��ȹ�ͅ/:_�Ͳ�H�`�'Vrq[�!�� ب\@%MC9j����� q֭+�aH�a��-9#A�S��#`�x}b8�=)�S����IU~�!VcZ��3& ^{n(d
*���0>�%c�E��TC��եD���p���p��B�PRKƼ.���eL>�����Kyb�C/�b�'-�^>U������P��l����s�8C8erA&Qş<�	?��-z҂�=$D��Y��[�_�T�㨟0�'�.�`R�ސ13�ʡ%� �`4�'3��f�F�gB�A�Ƒ�-+jIr`;dJ�� f�PrcH��0�	�eWC*a�!�|~bLˮ�?Q��h���)� �q36j��K]tZA
=D!�s"Or��2	�rIS�0�*s��3�h�� A���ei^�v�Cb2 r��'���'h�Hǜ?!�(�'|r�'��8�X�"kײ
1����hu�T�WOɆ״���:�2� �aƎm�1���On��s퍔!��]h��Z�#`�8��%��P��%Ʃ��'�sA�ixH?R5#�
p�j�]� G:�뒮��BCƀ��N: Xf��%?9#�՟��G�'V�bdON�	-���Շ�7]h��"O��4A�}���=-Y�y*�R��;��4���$�<��
��!��Y��KL-�B}!"��\8T��aӦ�?i���?�������?ٚO���̺G�\�iQ�X<4�1�s!�:{�,�$dVa22�:;sџ
�+�-~t��n�J�R�@�?*������d֬��gS85j�h���\/���U�DÍp�L��!ڐ)��)�f��t0��'*B��e�'\�iĮI?θPC�`�Mt���'��`"�D�;�x0�$L�y��*N>Aӳi/�]�dˇ�����O6�jCdU�Z4�9f		R��!����Ov�dũ^ۈ�$�OX�Sm@� ��O�B�H��dM�6#Vr�nH,wcz])5��,�AO�N�џ�t��e�4�2(�|�r�hHr&��-lX�f"��[�8�(FrG��˖SUqO�y��'�ғ�8�a��LC���Qj�qm�	�&� �O\xq6�B	���<_�Jl���'Ң����G�X��/��8�̃$�u�^�H�P$���0�I����OND8�'�F���i�>}⒍���4g�1���'�"/#w����l�9�U���N�Z�'��	�:N&X�A�# �B5C&
&��	�pt@9���\F8�:TO\(�sf��f�*�P�ן`�ʷ���`�a`EI9NZ��Ԑ�����O���'�'�y�ȿtD����n�+�h �����y�Z}���se�7s,��q�I���O
�E�*�� �2p��c�o�bc��?��?��	Gl�:Sf˗�?I���?���y�@��a�
��b�27k���ň��gn�1�.�!VMֱr�EEo�T�����|���W�.��5%R$4�2QA�$v�*iXVh��h4"�C��^�iS>����XH�)�=�@|�08塚��Y�dk��3�D�
F��P�'��I�����Od�=�EN��	�"I20	
�gǌ)�u�B��y2�P<'�r  �O�f��L���G���_C�����'��I�S��Ā/<pZȵZe$	+n,�0�(J3g  g\�W�XE��nЎR��p�,º[��(]Y��D�w�
�:�`�J&Y� �'T:��AS�'�^����'��'�)����\p�����<D6m �g��'�քS6��,�s��胲@�'��Ӄ�JP�]�(�Y5�H��0�f��<2v����t��t�vf���s0�	 ��D�O�b>aa�l'u���7��f������<���\4���&Y�"� �eM7gGjP������dÚ^�
�S�<|pDc�L*RH��(n���I�<�	d��ߪ ���'�2C��QNx�4&ğ0� g�'#de��	Z�|9qb~j(á�QD��
�$5��� ���02zI�5%���y�hÑ)q@�e?��8C,���&̐�]�
S����\��k�ǅ�)K��s�ʈ�I�ՋG(��'9�)��5?9m��Z�^�����5#*-�(�|�<��\ s"�ի�]����B�`�'|\#�'ңu�^�cC��f�tY�Gg�
�?a���?A���"��H���?a��?I���?���$  �z%%�X�(�	% �>4��BR�7cl�!�VI�gd��ʟ�>D��p�2��O��]3ȵ
D�Hw8��(D��� ��:��-C�� �Oo>8F�1a�h���Z�C�ߓBF9��ԤG����' �� ���?����f�qW��jظ�saI(<h���A'D�Й6ۮ�hC�o�f��I閮�ONEz�OB�U��z�#
2\��ڐ)^�!R�`�nZ/Oz��C
�Iӟ��I�?�������'g���6Fe"!��BJB�Icf�k�ySW�Z��LQ	��ɇ���!��V���<��k�����xр!� �2p�lx��j�'aj�)1I^�.������D�L�
�&�����0r�R6����b�'�j���
�R%D�U�L5�$�r�<�s�z�FAQ$�	*5:pa� py��z�N�$�<����!W���џ|ϧio��A��M����`(�%���I5v�D��͟H���A ��gȯ,�J�.���0�腰��AKw��)]��8@�RE6-2$�_���K�ISWF�$@��?u�0����3��3���*$�D�K���q�<8���#Z�qO����'B�H�.J�b��bv�K&#�����n���	a�X'2��*�`.'��Y��7�Ob�'��3�T��:���!!K��(O�L����O����O�ʧ,-r��?`�	�40�62MKT��-O
�?9@枃\����B���*$ 4�7Z���f�'u��d��" e��P�k����ΓGʨ#��NV�*uI�nJ�G�>���$B<\�JY�4�t(\t�H�I��(��&�y�)�B�'*�)��7?� �s a��R��!�T�:[p���"O��yC$�D�`P�0�R�Uي��I��ȟ���/ �sv�q��� Mt��A��O��Ol�%���'�0�$�O����O����O8���ݨ!������_5/���3��#m0H�T2i,邡\�/�P�S��O��)Q�ޭF&���D��
`�׏���"Y���!jt��RJ��e��ӦiC0$Y�"�\����&��K���}-��W�Č7G�ɮ(��d�O��=��'%^�[� I#Bɖ��Bk�\��� �'��"eB��J�~UY"�U�V >1z��-ّ���X�'0~QADk��d��JP�J Y1uI�
؟f��p#�'R��'���O���'.�	�\R�!K7��9Q}@�X��D!d��x3�	%V#��	�������@T�'F��C�3��-	I$b��i��EN�=�Vl�
LH�b�-��UF�4q'�/W��5�=��W�*Ј��e��5CQ�/��9s�(���G{�	 ��c⊝;�*%���J6:�B�	 B�yuA����)��{$�ʓ>����'L�I�G���4�?a�����o�5�:�p⢊�,�,Y������?���܌�?����?iҋ�Y�MX��)�Ɓ�Q���:��`��k�\�� ́"�44�p�nc��EyBb �Y~ܸ�&I����*��Z�� қkJ|z`�Q���2�ďff��W�I<���@ �?Q��ԃ��UB��Ŵ@zt	�Ȋp�!�$y��􄛴B��hq�G�e��h9�	�I���B�] {Pl�W�W�]K���?��?a���?!/�x�'��f�,(�X��0�@�M:HD�&:ڧh):����M+T!�.��^�Ɲ�?yЫG�	TJ�P?���������1U��#��(�M{��ЂQ8�'�����?����?��'����b�^)0��do��qS�E�Cn	\8��'��3��'~��B���u��?��;>
*���ɛ�y�,�j���75�@����O��$��Ty2�ǺC��?�'�?Q�'}P؃Pϑr=�U��M�2X���?��E�u��rQ���������g��;�ꆜz�$�#w&TQ���2��ԟؑw�O"�D>.�L��ܺ{��?Y����!�T37�XI6b���`��P�T#K�?a��Ma��0bB=���4T\���޾�tըv���Jl�2$�\S��1O��V�'Crk����I�O����� ,;b������̠wTh��&��	Z�0�$�Or\�;�?Y�'��]���O ��ĉ;~��R��,a��d��H��b)�1�j�hU�	*�b��O�H�Ve�$�'R�J Wb�c"�Df�����x=�6ˌ~���	�z^Vel��M���?��'���1�O+��	�=G�$�1&E��1��i��W�h�z����������MS`�Of���?����Ma���p�u�܀��L� �yb�X\�&Ȫ%JL7A).5+�K9�M����?y��?�g[?Y�	���M����5t;�q���Cu���զ���ϟH��ٟt�	���	џ��ItB�/Z�6����JH���u���y��wy��'�R�'�"�'7哱:�����O:I��z�*[�7ꁻٴ�?��?����?���?Y���ɇ2��T��Z�4(��B����<�N�XU��n�eA����x|���i�����O>˓��D(�$��h�@+��Ex��ń7J����"z����<�/O�OT�d�?u�bϚ6,ĸ��c�6��<D�踵I���|< �ό�_%��@�9D����"��(�	�͋a�E�-D�ārƂ�r�%��M�v��eA��-D�Xт�@0���G�� F�rqL!D�pQ����ow�K�	 l`�1�?�
�$821+��~�,@)�ޝ .t�Pꃥ �>d�RC@)j#ީ(�Z-��KV6S�<��d��>A����bI�%���r���ah�u�L�hz1��ZS�	!F�9J���7D����u�Pp ��S#O���i"����(�E��.4)�d�k��B=�"�d���%B�(�~�ѡ��"�.x����Y������(z`9�L�^�(�Y��=Y	a�Ƙ
�h�`��̀o�b�c��.K�̀���\��l�9^^)�"�'�Xゝ3ͦ����?i &�>�?1�y*��	\��\��J_7r���ag���!�4O��:��)�S$T'�(���֜-ɬ�K��
�{j�O�I���'�O���k���2߂D�ì_�l���"O轲�.�?��RF�ʱEL����'���<� �<{�� �S�G�q����$�	�6-�O����O(�c�D�P���OP���OGH�#vƨZ�ΕBZ.�RE�&��c��ڑ�",O St�,2���צ�5T�u[P�d�V�ay���&(�Sr��Dq�Ѣ�ϒ�]�%�̂��Oq��'+@�k �&D�-S+È?��S�'�0��t�^����B�ȯ;�ѩJ�l��4��O�0��w�̩�%��
Ka���e��o�XҴi���`����l��
�u�'r;�� ���J� ��*�4'b���B"P�L�!��D�? D2��2K��{ӁR<AW�q� ��x<	��X�9�vē1@9lvI`dپ;���I��p?9�Ê52Ȅ���̄,�E�iI~�<	�bӏ�JՃ���q�rzv�IUܓƛf�|bAF�^=�7��O.6m,R%
e���9jb ��V�jRY�Iҟ(2 ��ҟl���|��(���(%�\RvAG��j]#���i}�pw�&,O�i���I��H���������B� N1ay���?���>�%R��b��h] !6�8���b�<!4 ղl�d��2*�"6��x8g&	H(<�weY�	;X�@�œTC��ӱA6KS"4�H>0/DR���'$�^>�8�HƦၖMW�
7������ۅ�
�?���	�����(Ǹj�������PY+�[�6�t�ҭ��I�a�[�lP<����<v�T�$�xr��K�)r�O�{Z�����F���0THq����%Q�����M)f�x��EB�2��Q�������S�O�4�(��`pb��1+�,_f�<�ȓ;�H�d₰P��Ū��=$����I6�(O4�`�͂Rjy�CG2QU~�a2�X��M���?i����i�e��?����?Y�����Ʌ1i֜���p�r�s!�1Θ'جUR
�J�x}�$�H����b]��.��>a�JeX���&LϢxP�ӏ�^j0tXA+��'m8th�S�g�I�Wf��rG�\�z@��$^�(�C�	�m��I���ܠh�b��cݟs �'.X"=�'�ēK��y�@[+�H!����$o��� M�!�\����'y��'r�O�2�'+�酩N+��F$V�}��������L��Of�sk�
>��axtꐍc�еc��NQ�!����hqQ�A�5�C���%&�?���'+���F�6r�R����N$1��Q�'Y`(�C�MV�~�[�mػ:DĠ��{�b�ƒO|���m�Ħ���æe[��m���r%�W�~i����F��?Y������?q��l�Z<��\D@��"
�42�R�,����xq����U�]Cdȟ�a��"?�ƠE�?ς!�3�;y�j�����8;�,	�h���a�Љ�8	�ҿi�B�� JU&�'�@���f�vkz�6���V���E�Ke7v���hѺ
�4�'b�'#�'H��'���i$ � ���;�F0�bԂ;6�ٳ�#��*E�HH��@�៼+fJ�:��#�FJ1n}��E�xx����xy�Á:v�7M�O����O<��!^�6�X�����E�(���3%�l�q��՟�j�'0;<�Y��U��T>}�O���P�8�L�!�q�d�1L<�T�O!��Ix!�Z娟ʸ�!�&wI&�cd���A��d�7�x�H�?�Ğ|�����F�"q#S�s�H ����y�-I��De@7Y�D{�Źyڞ�=ͧ�Q��	R�R�l����/h���" ʘ��?y���?������SN�?���?q����3"�^��pK�h��6�&��iھ��'����
˓X���<ƀ|��ʜ ���>	Յ�|X�`9��M?�j0-U;RԀШ��7��'ӈИ�S�g�	�e[�rd+�T�2��f�|C�I#/H���ǆq-4pPq�΋Ea��'�#=ͧ�ē�EH��R�VU&ы�L��O��n.JF]���O����O���꟤�d�O��d��LQ�5$A�����P���wLh1�%��C,5����3��O��"�e�2G�0���Ƅ<<���$E�-N���t,+g�\RP�ɍJ2� Jq�i�f����DH: g:i�c��JQ(��ed���\ ��'7�@�	��|�	A�Q�� ub�(8d�D��SR�����?q�.��|�����Z�GH����%,��'��7����I�'x��k��{�(�dz��HHR�]�R,(��pjN [ӂ�����̟���"7��(�	̟L�'qC�s3�9h�U�q�A��#bl\`�$��5-_�[�\D[r�'�<���ץ�%	��%�(Ia,�f3L	��*Y� ->�ayR���?���>1R�m]��E
�$bɲD��\�<�2�Y�c�L��1��4��Q�
V(<�#�_�蔠ҥ�f�C�.%�J!�#fH��c�v�s3�i"�'��29�l��K͌Գ!���p9ҡƍ -�jH���?����Sܜ б�<h�^d�r��LW��V�4��9� �1��,V	�HA�C����z��ؐ�%C96=�5�ҡ�R����M�@��ʓF��"r\�RQ8��tJU1!	LTБx"i���?��|���G�F����DX�M<x�%N(�y�eփ(�i��lβA�92bF��p<Q�wf�H��Q�F��`��gԉH�H�w�i��'�"�BDujP�'�r�'��;ak�!QTE\���I�JG?"�ސ�$�Ps1ĕ���r� ԛa�aj�S�?�r#������ t�2�$�
/*(�"o�@��!ԇ�:Pi803 �#�P(�Ƌ��Cw�=hfx:��� �i+7l״v-zP*0�Տ;wLB�"�M�[�ةs��Oq�r�'�&�%��;�*K$"i��X�>���G{�C���?)g��{ ��[�_�mf6<��WZ��������4�?yöi*�Og�Z?�ъMdn0H��̀�nY�4������P��Ȧ�?��?y��do��O���b>�ka�̶8�|sG)҅o�0��HJ(D�l��BB.g���yb �*(�v83����/��U�� ��	��x�!H;5��u�A�T.����(SqL��������c�I�^,T�@3�=�6 #Cͥ{$�h����O@ ����S�`#@j� �HQ���^�9ZHB�ɳm�ʱaS���#!L# �+b,B�p�ߴ����_?�oZbI��O�c���W-]�'F�����?��O���?�����*�z����4+Y�1UI� �D�f�h��øJ,�HS��\�>�d9I'oV�T�4Fyr@�?}@.�+��X"	۸���)�RpM2�hɽ4&0Ac�$kNQ@��<I�HdFyB�D&�?�����G��u�c%F�Oj^�#' ?|�qO��d?,O��[4���x��ѐ�-s�rMڳ
OЙB�B)=��̪���/��iȕ�K*QD*��<9A$�.����'U�]>��-�Ǧ0��ǖ��(8�cM�� ��� �?9��;z�[������Y�c"��zk���fힷt1�Y�Ѝ-�$&Y��b?��vbڃ(ň�ue\�l����k,�ʹ��)5��I��-zTI[��=�
U�S���#Q!��6��Ez�nɧk��4r��7=�x�*ʓt@��ضO[5v�ZQS�$V9$��h���j�����O�D�����b�O<��O���w����6G�NUД.܌`�T�Y��'o����,�M�.E 6N� 4Ďb>�q%�ٚ��H3>Pt��C%KK��)5Ií4�*���'=nH�4��R�xS�ɇ�~n�;|ҬjT.��"4��/ֱ$�L���I/��ְ$���L<��/�z�!`�.J�p��
�L�|�<�� -J��wFS_c�E��n�SY���$�xRFC�ts�� C��+;fY:qA�<NeblR�d]=?��D�O�$�O���;�?A����ĭL��ܠ:��]<T16o�3`\�"	 "T�np��ňT��yR��+"��ȱf�j#:���ÚP�#X)� �qXҘ���gM�qz�G}r��&2h�&A]�\�� �-���[��/�~Z��ȶ�E�q�� ���R�J�41��d<ص17)�C���ӥ��Qj��=��ik�'�����.�>ش3��1��,'�!E �p:$\8c�'�r��7\r�'��l��1��H衢��B7��9S+P�Q�r��e�
	]8�!1E㔛Nؖ06�+�L�q���Yh�Vʌ1`5�x�dW4yxr���I��4�F�^�q.v�� ��V����=Q��䟨�ܴ7�v�ix�pY��
�C̴ ⷧ>�!3���<A��ߞ��d(���)���,=���?Ɔ�i�f�I��|��ҟ���g��$�D$?�!��ain@�r��<��[��N�-����	Zy��Uߴ6-�OT���O���ϋm�p6m͍F��')߄H��I8��W�\)���	����O�ݦ��o	F`a�Ǆ�I��鯟��X1"��	��M��Ԉ+ĩ6@`9$���ңZe�����!|�=1�NVDܧ:׀yD�N��� �cF  �&$�T	��O\ $�b?q���A����s��N�j�O D��c�Q9�=`vA�%5!t8��<O�Gy� �X�a@�A	s���y�ǿ?C��n����埨�
A�%�:��	�����Ο��+��u3�ӠhV��p�P�@�y��]*�K`%�U@7�S@̧(�҅	��O�P�E,��f|�YR 1B�J��Fʌm��9Z�#��`��2%U�Zb8P���\z�4�U�F���,=F��c�'�%溁�GΙ5��͒W�|2�Ι�?�}&�d
1��2\ �㭆w#�@b<D�񧪙	
а')�(LT��:}��-��|�L<	�决,�ěL���f���
Е ]�8 ��"?���'���'#����D���|z&�+5����'^:3�q Dߙ#/(��N���1`��)�E��25�H�<i���k%�9��
�2�Rihp��$A4����V�?��d�Y�?B�hc�b�kC���ୂO�hGlM3�ϒX�}PQ��7n���p�V��C	�
H��c�	�Qp�{n�t��^:�-"h�iz0��'�n`�BE'�I��M�J>�bγc�V�'i�6��fi��"<de�x�䏽��d�OZ����O���l>u�$	!oH&���AC�.�n|�rh1��\A��Xb�� . ��D��!��	%$-S��L���ȲH��4��2 P�R����a�˦��O^��4�'Ml�'��]�̈́�v-�B�3p.��'>ƽ8������S�b��5!	�'��cΔcp2� � ��&`X�HC9P0�'����ic�t��O��'n>��ٴR�\rSO6��� ��8# l+�'�R�Wd�@���̾vd�;���O�H�4�G#U�����E�%Ȁ�����qp�  �� ;�6aag���(��A�@�ew�%�!K� "D�(17�x�Ö8�?V�|��� l����%��	�.�P�A4"OnD�߿+��L��g[�wt})��' P�<�Ç-nZH����fR)W��-k�7�OP��O�y�T"gѢ�d�O����O#K�X4��i"�лd�&�Z앣x2��N<	G��2G�``�|&�(
g�P� �~Mi5E�H!fa@���*P~��s�^���F�A�����o�h��%��11����#�S5)�����4�DS4)���L<17��8w~ȱz� ���ᲒE@�<�/�|y;�����X(�g|��Rn���D�x��GRX��gL�(���0)ս��[��[
Gr����O��d�O]�;�?������E�RL�q C&>�z��HP�b&�R����1�0i�%%��� ��ɜT�ِ�Gg�E3�JLS>``b�_ڠ�{5��)T��mPw�M�']z�`�	�)�#�@�f�������?���?���������E����LU0 F��o!��&'�4��rˀ�t�� ��	1�qO��o�ɟ�'�i�D�~ݴ<J@�1��#`��q��(X�y���'��mՎ���',��];Y��]� ruT���G��R��)�$]���#E�>{P��F�2�]6�lZt�J.PP�f(�|&I�$�ǲuD4X�E� k͜�q��<�M�U(D��O�HC�'J�\�,BW-�@��`� j����A�4�I��剃i.�H��È=��P�H��r�"C�	�hqp�J1T��q"�i�)�3���|�'*qk� �`������|�6�L�����.�=��8�l��������N�5*��c�&D��l�1��!��)�~b��@¨��HȰGxp!��MB�IP�.P#��ۂ�AJ�K�ֹ�}��8uJf�ش�[�lx��-�~�I6)���D�O�}�޴���с������� ��6���O:�A I��XwJ�1�aP'��4���'y��<0�R9>D޽�2e\���
�@ה(7��Od���OR��0�U�Oq����O��$�OW��~B(K��5?:	IP(�t�b�0��,,O��i1΅�W�ȡb5�թB=��`D�D�Jay��§��j�H�V*e�Ӫĩ`>1&�x��j�Oq��'��R���3;R4`�LU!+��Q��'��}�/ �!rĴRG�D� zM�t���4��O�=h��Q�DxB��S��dI��&#d��' P����̟ ��5�u��'8"5�r1�������'g��O�����&�"k������͖Y�l���E�T8������(O��*�.A'����R�J��ф�t��x�n���)bIؙ";�I�(A�(O�ر��:8Enq ���� �X�5,��MҌ4�O��	��A�*��$�p�:�D�"O����Ӑ1E����EϜ[��R$��Ҧ�&�l2�h���M3��M��!I�O�{��αP�z�S�	Y=��'��be�'��5�2�1l@4F�� W/�m3\�A����	�������4�+"&��s�R+�(O�	����� �f��L��a����R0�y4˟(YƦ[��\y�#c"��(O� W�'N��'_b�x���i|���.ӰW��#	�'��[���j�M{7/D�U1y��'������, �PP k�5>�,
��W:��'��5Ia�g�"�$�O�˧"�&���4[�▮z\ �y��L��$!��'I���an����z�*�b��z:�p��'���@s��R� \$X
��a�k���O����nW�'o��(�B<n%��d�͏���	���
W�뎐	[��T�BYb5΅R!j̉'�b�;�d�ɧ�OY�e�@
� �.�ۀiI�y�>�	�'�*0;E �BT�;SjŲr���k�Q�T
�տA���:A"����=ٱ��V���Ɵp�Irj*�I M�㟨��ߟ����]:6�L=h���RƬTT��e��&S8T���U���W��U!�k.L�Y�O���C�w~��R/3&��ƭL��,
�Hր2��u" F_�n��d�GL�[�F	(�M7
c�'l��;S4����'���S!/�5q���A�ț�M���i��m\�aW��,O7��x9�TP��&C ����V~xD{"�	]��#d��@�Ľ*�</��'~v7�Xʦ�%����?�'k(I+$�[��\( �c�"��&� i-�h���O"�D�O��[ݺ����?��O�zݻb+@Tȁ�c1`�������#�@��cB�:P<�*�lk�l�a�R�'�@}�W�ա]��cу�G���kr��<s|Z%��A�4WhR׈�$��̓TA�)jv��J�y"�*Zr,IԹ=K��0�Ą����!��~BIݸ[���ECr3���%S��y�*��`q�T���G�`��h����4Ҹ'�J7�9��`��T>��%H�=k�@"s.�3L�����l7�If؞�I��S<��8�凍O߾�p�$1D��"��!���"�»]�ēT�2D�����&^YD�� S/��-#h2D�� >ȓI��Y�!�(�r�ЕJ�"Ov� ��٨5�=��G��	��ib�"Ot��DS&Z�x<vL�3o$0���"O2}!s��-g�f%!E���W��1C�"OD{r��V�&$�6K�S�x��"O ×i�6?X��ڀ��Hlfl�"O�p���&'�"����:�, �"Od�"���&y6c˟�b�Ę�"O�)(!O���p�p��5��H�v"O�]�g�Ũ1;zIr�*Ǚw�
�iS"O�P��bc=�]�ֈ�
Vk*�is"O��j�{Y�|b� �f��,X$"O� PP*H�Al$mIC(� �L5�"O�e�Ő<\� �*6I&u��+Q"Od��̂�Ѓ�h�)J[ |Av"OB����v�\��`��_>H-BW"O�8p�dۅ10� !K7:3��`"O�Yp@�<)����aɸI*I�%"O��I�$�OF-�Ug��F�{R"O��Z��Ao��X��`�E�2ERs"O����̝�<:��/Y2
��q2f"OHbu�D#o5�h��M�ry(��0"O�M	�FB��6��p�]�Z�9��"O���$AC���(ӐND]P8�a@"O1`�Jb�@!��N�D� y��"O�rQHĞ	β j1�,~�ȫ "O�@��ID($T��B�@pkL@h�"Od�be��h'�h[��:ha�YbU"O���C#ƢPz�`�q�љxYV$i�"Ox��e�ܐ/�,�0k!,R�@+�"OQ�&׎s�����ȦyRዀ"O�b�M;L%��H#�,AcD"O�Yj�F!V��8��b��["O>�hB�&p���J3�"T"OZ`�iՊML��kA�ۺ �T�4"O�"��I<�^h�!ѐY��8�A"O�� e��^9���`��8�%"OB��R�&�<�Z��-��W"OX�C�.�/��i0��O&w�x�"O�帶 ��K��kG�D&m�u�7"Ot��7g��ca�l!�7!$8Lk�"O4Y����f���W����"O�K�)��4T\�0c�8>8��#"O��N��`�Ny��^�2�aV"Ot|B�K�E ���l�=(�ک�q"O�I��Y�qq$1���?�h4aR"O@cu��92(��jE._�G"O��!
{ ��K'�xE��"O����Ykkv1����A��x�"O*��W���tC�Y���(bp�"O�=���Q=�R��⦀6%��q�"O.��fdM�<�XZ��Z�}��2�"O~�`���CA����aM��,���"O6��E�lD�+ Yv�L$B"O���PA]�4#���D���ҍ��"O�ɉ�!��4�^�we��[ l)�"O���#뇜<n����eD�$#HŪ�"O�P��_�?,L��% ���9#�"O�=bW,ȁ̃��D,W�H}�"O"�aW6m͆��!|���B�"O���J
W�=����5��M��"O���O_>Q��p(�تMI�"O�eX����퍟o��a"OtY��!5DF�HY���J�q"O� �C7��-}4YW	5v��X0�"O�Qr!�� |-��G�R~�� "O0T�qM�f�x�0���k!�ՙ�"OF�+`'*ސ�jF"�
<���R"Ov�z' 	�BK�e���%B����&"O�#"����B0B�7a��xX2"O������T(�
܇$��ȨP"O�,H��ҼbU�
9O��$��"O%�W�Ýj �@i�=K�)�u"Ol�ل.�@[���Q��Sy��R"OxpB��!�*���G \Z|�"O�A�e
�r#��yp��bE<�K�"O�x��lJ|�|�0�J&d;R"O�l�P��<G�،����
��h"O����K?M =�.+�� T"O�U�v��3.����J�<N���zw"O00�Fňt�}& �.0 �"O��p!C��q3�	e�`XD"OJ���k��e������[����'"O����ƛ_z}x�
E<A�G"O,Uɲ��%A���a2ŏ1��1�"O�m���Y2of�p� �ڔ��"O(�ږQ*/P)�t�޲2�"t�"On8U�Խ�R5��D�?��lp"O �
E�S�>Av�[�3�2��"Op��7`�
h�̰����*�� "O)��)v��е�?]�,Eys"O� �!�/ ��05-@�?�`ر�"O|k�  yJ�˱M˂����"OHtҰO֥����&��%�x�"O�����8lv�1�b��~Er���"OR�)��������V��x�"O �a�-�%p�i���C"qɆĀ"O`�a��!����#��K�����"Or��%ԔY�$an��R~r�!�"O�D���0�RY*Ҋ�*L�)T"O��u'��_���@x�	"O��&��9HEv�q�������5"O|b�!�S�>	�Aa�A�v�"O��yԜ#��Xu�Jb�Q`�"O|lbg�80@�r��!Wvd3f"O��� �-7���h��S7)��t"Or)��iO�bjѸS%�.��"�"Ov�c�K�9$���2#˃>lFA��"O�,:�ѱz�|�K��/B�iГ"O>�3�Ǎ#�n��Cd,>	�B"O�q��]�Cr�`�,P�!n���"OLi��\�[��qb�ߛlbЭ��"O�I4I�y3�2�Ꮋ\�i�E"ODE`ץؒKu�MYc 
�^�h�`�"O`%g�R�V<�!SAJʠ{WX0�"OIۣ��"f�숇�Q�&���"O0PQc�p�4�I.�,�"O,�Fޑoa R,C�qvF�y"O���!ZآIs�
�~80��"O~��N�+?+pYq��t,�ZA"Ox̛7 ȓN>�����%�"�P�"O^�Ӄ�[	G7J=�BF��<�R�"Oj�����q��y�Gb_- (�#T"OZ��d��#:�(6aV(M���A�"O�Eh��S�]/>j��R�KO�
a"O:1Pb$V����;CV�=ۤ"OtEx3����Z� �k�'>��q�"O`�k�k�d�������$>�\��"O� �����[iU��8`) �5�"O�j�-�h��U[�ə��6iz"O�u�'̩xk��"r(HE�
��"O��K�L�:;K|��@��6��A�"O�8D�ק)5:�F�� 7���"O2�h�n��_l��t�'�jE+p"O*hZ�b'o��Z�.M�z��a�"OH�	Ѥ�E���;���\���"ON"�.�\>&}�7��0���"O�t�7DJ&?b.�X&�p��z�"O.�ThV;HZ�+%�ӹq��2�"O4�ht��m�HY{3l�+	"F���"O��q�5��x��-�\�@"OҀ(�Da�l�p���+Qz�z"O�H��Ԭ�4�Ń �?پ��"O�l��reX���L�>)`�c"OP����4��Ej��2R��� U"Of�BĈD2aP�,�Ԡ�,"�Tp�e"O�U+D��FW��Q�EU��ܐ�"O����7BK���R�˴^� 
2"O�I6��RxP�`@�en��0�"O,�ju�ٜox�I���X/6У�"OH� gܻ�>�� ��:0��"O�B��\��ܠ烏�NR���"O�$���Ư+�:�`3�
B(I�3"OD�0��̜6�d5�#��#��Y�"O��b�V����k�"D�j 9�"OZ,���ӗ�)+j�I`���"O@���E#fĝC�&D'�h�"OH��@G�:|0Z��j���"O2�� �2$�6��QD)uj�\�f"O�Ţ�FW�r$�(�ŋ;L�`�4"Ol���%�S�F|B��x���C�"OV�X�%�
Zh����]�`���"O���0�9I��1�@�R���d"O�cŉ�5mc�M����4aZ��W"Or`�pD�3��R�.�����""OP�bል���E�ޡe�0��"O�dJƌ�&\�d��TJJ�"O�qq�M%eq]I�֫;�ʅ�"O¸a���7/�@�0�<���1�"O��)D���/�ci�
Ҩвp"O��!¡I��T�(Q�T��yzr"O,�kIx�\��f�.м��"O>a�v)��_-4���f�j�,ܢ�"O��ct%с Dإ2Vɴ4Q����"O�ii��Z�Rʈ�S���*B�dxA"O��#V��h2�<"���,�
5ҵ"O�!���J�%BD(A�4®�g"O޸p*�P�ލB���+/���"O�y�
�^���+��u����"O�ő  [2-u�d��b Wc2��e"O��r��/#%�$�d`R'3`0h��"OBݻ`��<��dRr��0[DZ"OR�C��P7I�pT�d@O;@yZa0V"O���┉j,�A�ȍ7Ŭ�S�"O~��`�:4��H�2h�(t��"OHK�C |��}��6R��"O�<�h�20�a�^�G�f�P�"O��X`��<\ !�B��,��Y!"O&,AwNϥⲅ8�h�-b���0"O(5���}ؾi�dE�_��Qu"OJɓ�b+?�T@�C)�*s�@ے"O(`�⃍k�d�R')�OTPm�S"O� ���Bb�n����H�)-.pY�"O�%��E�hB\���ɑ�J'�Xa�'�`s��e~��ЕD����q�A�=�&��86D�ȓ��!�G��If�W*�<��a��X	
�:�GB/),���a��+6H�(�ȓJ4�@J�c�� �bĬ59xلȓc��5��H �&Fܑ��	tĄȓd��C"6
�@�b˝({�I��8<h�f�q�d���"����A� �5O��Qq.@90�J��ȓ��!� -��ʗ@MBF���ȓg��9�g^�{1�t���T�"�h�ȓs��C�d�"W���j�LQ>^Vh���w�d�Y'�ι6�����!��2쀅��p����ߜN���H��k붤��W�@����!L3�-#�Mڸ=,�%��nĔ�����K����{�	�ȓ`R�����$ڣc�0p޶E��D^�i�J�L%��ӲB�0W� x�ȓq�Hȩ����p���C�$֔;�f<���P[�I'�R�{� �,�^��ȓސ]��H�L��@��fф ��F~��-"Q>a��%K tb��q�6_���yp�1D��j��MPʩ�RjX/�^�Z6Dp�\� ���l%�t'�"~����%���� ؉��"�LP{�<��N��v�>�X���^��k���u}���
6�0�xt�O�=t�x"m�Q��[��
B����$�>y�eUJ�,�2"_2lM� h���8e @U�� /Y�$�
�':X0{���wH��R�Y!b�@!b���t�b�Jo��s�>��C/`5ԩzCc<�T���R�!�$Q	ch�y��U�9/"��VB�s��2�.�w;\���*R�(�t��s��L�n�Hp▁�4p�8[ �3D�,)���^���!��R����]�&�ѫ}���&�C
�\Z��d��G�1�W�8y���B�FܠJ�{B�Lt����i��`@���
�R�$� ���_B��!��>�!��6 <��T���f��=�$�B��O&�r��l[ �@�C�fʚ�>��҈�%H8�u��D�cDH�"�@>D�t�%"J�U�h�r�i5RU��K����[!�	g�h���'�#}�'���e��9���3�DV�S����' �E8$萄6����O�zR05XݴH���#�^��QG:<O1"&��6�ިВ(Hֵa�'�$�Кv�b`@D��3;j�3�*ã(1q��ύ(�d�8���S(�~��Աo�`�c�@
'� h�wNº��'�������'G�lR�!��B��� ��~₰� S�܊Yw¼�q�B���Ls����_M�@� 冺�H�#�����K�n����$�g?!����[pP��f��7d��puf�n�<1��] @M���$)�llz��B�3� Ь[�2��®��+����3�6�DP����xW��J�#G�2�vM��I\�ʕ˰cJ;�(䁓�U%h��q�t��Ek�h�3G>x�\T��	�4�0<;��]�%`$�a#���("<��%��`zr(�<�J�JH~�We��t;���.T^|2U�q�D�<qpjI9x�Y����	3 !�P�Kݦ-+g	��b�x��4i@y���iyt%��	�>,��iA.T�
�'�(�B$#��P��xɉ{���.OAK&�$d��Sv�'�~hyG�VM�����2`Q���)q�KۛC$L9c#6 ��ID*?s犜�7Dʄv�a"�Ïd�2�2u���[��0� Y�8��'�|i��*�EIz|����tM4�9S�C/��X��Uu�4=Y1Th
*c׋W0._��Q�J�C؟`R�ѩs�<l��KN�d�.�8��f�6e{��;5��&/�n6��Ā�QN�q1gW������̚7�y��ڑx��Yb�	U��(a�ǜ��.��K	�uaV�Q7	��M������Y��(q��ߍ?�p� �:!�D6M񳥆�����bUJ^;n�ƢA0^�T��Zu���JbÅ*��O:}�i5~B��'�+��aj3�'�^�A��|�����˅� �t�b)��.�hȪ��˃\�Jx�C'ւL��I'C����N�T���J��1r,b��K��!RE�t36�G)^��AHGkfӉO�f���C?�@�A�[�4N��
�'I��w∕D]$�(0���-���R [gXH�A
�"��Pjڴ%�>y	�O��{�G�2z�]��#~��q"ODY�ϓ9^���NL6 ]BV�i�|�xP$ϛ?a�؈���k��������0����A�S�ze[q�Nbdaz�ѹy�2��c#!���������*�A���0B�1z���.�O���j� WB��V�W$r�I����_4R� I��;~��q'@M�N|�"�e��O
C`Eȳ�5�C��!j�T�)��:� �rP��ss6��L��R������>'�H7m�v�OPN�s���A�lכ'JJQ&��y�zȅȓ�g�ۂ'NTы�nG�1R�5o�?��pZ���:Z�V�5B�FM�"?Q�)PJ$��r.0g@�R �c��h8
�`�)��m�x�Rǆ\3 �4]�L��*^8qK�D_;U,H5��\yR骗&W�6(Qr/�1��x�<Qp+��zxʗ#��Z)�E�d�¦�������n�찰Ԋ�p꘱"�"O�\@a��~wf	#�H�4{� 4)E�4vL��uc� r�$H�u�i� "|�P�����B�"�`����Qt�Y��4D���^zsd̚0-�0`�&ܡ��yӾ٪Ak��yS&�HՔR5"�	!.�Xxb�L-+j�Ij����k���������@Nĥtǈq8�Ā,l^!#�Yw̦��gn��=���Ô�b؟x '���%�x0@".">>��S�M?�	2~�R�I�R��[@��7��t�a� ���%��c�A
�y*cep,�d�������d��E�2�1T�2oF�HA"@,�MӰ����DW�ߌ�r�пw�qda�aK!�M9.d��6���"���t� �&Í���U3�E�/Sخ��q���O���5�Q���8S�_�ѻW�'
)���Y�h�*��y��pg.8�����3y\���bʉW�����G�@����3M8nk�\�����Z�!�d� o�h�5/B!M�CR�N)jm!�E$_/�����V�R�[��B��!�dĄkNZ$��@�F8�E��GB�9!�Ĝ0	�h����9%������:{�qOX��Ra-,OX��a	ޖrm ��:�x�R�'�X��e->�|P�Ħ[/�݊��S;����'8�P@D���.�PD�U�߼��L#���%Xx�UDܧ\��a�)ז')��`3�޽S����^;x�s$ �9W����n��22t��AP̸�!��'4K��h��q� �� *Yy`퀙#��|"�"O|���W�EmR8@#� �-2��^��K���CTJ����'�r�	 �UC�(5B7
��VC����a��Eْ�^ ro.i��!�6>J���+<���!�O���Ē9Z2��RD�9~�*�h��	�!;�Y0cK[�?1�gWE�4��P�(]ز+�	W���dN��y��?"��3�� $cd
��$�M��Gԕ8��`�\�!K�OS��M�����|�b���3ֲ���Ǝl�<�Eƚ:3�5*���� эG�d��7kH�b���x���.P]x���HO<�#��G'*<ĩ���O���i��'2>���3b(R�J�8|��f̶k@ݛ��K5!����O@�`�a}��_	z-�5@I۬S���@@7ʓL�t��~J�iť�Zf��D�]f���	iQX�k G�. ҩfO\��ybCF� (���,Ppt�=��Y6d5	�
�/oH�C��3M  �aK6���y��ρ3����VFX�W�L-��2D��(T�ќMsf�p�	�Et(Rié��4oF-g��U�P�b6��F�'�]��	ϧ���{qƆBz"Y��M�E��R�+|"� ��+\�4�kX;Y8�Q�Q ����m8�O�<ش��2�# �;�4��	�>�m����B��������,5�|� �Q�Cz�`t,��C�	�M(܄�AþI�	yp%�[L��](!�4�@Ɓ�G����l0�'7^�+��"%q��!� �n`�)�'�=�*�f�)�b�3(#>��&��?a"�@�r�v9�6�S����.�-�1B�&澕XteD�������'�|���!�}+�t�W��Q�����V�Ґ۳�8�O� �t��[-v�����)�!��IX��`c(��k@�'>{p�H)N�B�p�4C*@�Y�5D�c�-7c� ��'2x3�c�<ن(�Op���M>E��  _:� ��A�	�j���]&�yBCI�`T�,��D��x��D+��'Bd�Xf�'��ti�����DM�U��8q�'�f�SF���S$�]�4�AK�'��ԓ���8��Ԣ�CM�j�'b�)�&Y�!���y�G	�K�����'���/Ź-� ē
E�@y��'�T� s��@x����@��Y��'5�-˧M�
�D��� ¡{���	�'��Â��a�PQ���y\�	�'��e(�n׽U���h:u��i���$=pQā�s|ze�or�<)��Q+$��k�+�}�xq��PV�<Ic
�B�&KE��i�V�8��
N�<y0��pp9⁂�*lӈ�XUB	f�<�A��.���QCF$3L��nIe�<a&�$�M	1��r���q3.�z�<�� ��@B&ɇBvA��t�<w� ��8d�a��cQ�p�D�Ce�<���@���veVd���id�<���z|��E�X.�%�SO��<)��ǟP�JaK����[+�����{�<��ٵ"_���`B�p�,�d�Fb�<�戇�<�"%
 	�;v��!8��a�<3K�>xv]�@�?7&�a1 z�<i��5?u4hGMſI|����A�<���e�J���ݽV����e�[�<���=6)"8[PF^�'�2xc3ā\�<y��\<��:�퐤F013p��Z�<�b/9*���G!BXl��TQ�<��� �+Iz�ҳM�7V������Fg�<)��X�$�(�h�0Lu~�0��m�<a�c���QV�ƍ�Nh��#^�<��$%�nH�GS�]ZQpqfV]�<��&GV��3@�ٍj�t���id�<1�nإH���{3b�Q���H�<I塙�,�V4�p�R�b�
��ʔb�<i�'U�Rq��������UOv�<iV��pX�íK�#���	��t�<	��|�H���!(���u�<�0���b�!1(�3|u��Y�/�e�<�!@ś W.}�Q���2���jCK�<��v�F���oOF��	"�]C�<�4��4:�I����\�rY�w�y�<q!��)a�̡��ާ�t�w)x�<A7��T�E��v�H٨f�1}�B�I>��%[bK�"1�@��|]�a"OlUx�B����@�R�B�.��"O.��� �faD�Tj��X:ځ�"O���7/[�m�@��cP#x�� &"O=����<Zv@��,���`��"O�l꒧G�$�����ɏM� �(F"Or@�A#�z¬�AID�)��9��"O^��w�4 Ѯ)3�eO�T�1�"O�<����*����"O�XR���:w�bL�&*�63L"O$ �u�6)Ěy�8J>p(�"OH���д��$��ϋil��B"O4]r��w�J��/ޣ�.�R"O�!����'R�z�k��V�h����"O��z�%F.�:!	"�C�I��$��"O� �h)ևϱf�V����0Z���"O�m�BG�$�HGZ% �H�"O����"\rH@���a%�kt"O�����)K�^�pG�Q�8�Z�ڑ"O<���F�%�x��T)�/X�y��*-�4dLW�>���bVÒ�p=�W��_�ձ�@P�o�4,7jNq�*A�SiG
>�[c;D���E;Paޝ�F�N���Jץ%D�ĳ$L@��� �H��%D�p8���P� i��cR�\X�.#D�(C
ڸ�h�e*K#c��4�!D��*'��9Il���<mQ�����>D�h��"�,��q�$MB�j���/:D�!�C�c�*���
#=yx)�-D��z`�d�²d��2�`ES�")D�<kWʎ
[�\3�B��\Taq`�&D����*Q �d�C�"�J�*D�D��L:f��1��МR<�P�)D�`k�"�g
��"��p��I�6��B�	; �(��]�+�h	W@�Vy�B�I<o����W�@�����o�E�$C�I�vi4�yE&N<C����0��%��B��^T�C�T,4� ���l�;�VB��t�^	+�J��x��̀&BB�	������ ���d��u,B�"D\�<:E�8��1c�ܫSZB�$�0a0үA�E�f��B�;P?B��3w�D! A(��h�.\�E�hFB�Ɉe���p��D�E�Ԙ��
S:B䉙I�D�`��4"
%�5N�;U5 B�I�9�i�K
E�2iJd�̟h��C�	�4���Ѱ�K��}��`K�3�C��[>�b�b[:.���5�W�C�	6I��� �GY!T��t�����5��B䉿d��y�Oӥt�� X�"�LK�B�I<7��BF@�H�0���-/,�B�I'h��#"��=�dmqGM����B��F6usԉߐx+��'E'\xpB�	�K�N	�ԮJ�]�h���^�HaTB�;Jv��Y�B��	���؁=	>B�I�k�� bb)��c05��c֦I}B�IiX�)u�՚s�h�ǆ����C�	Z���G�2ĚT-L�,��C�	S�8���>Off�hFH��Z��C�I#2<E���D&1��*�B�]�~C��	�=�P`WX��� �˻�zC�I3�j���풵׮味JKAB�7aڞ��V'��.Vp5I$�? B��;{|�����	;p9;�h[q1�C�	'KO���#���q�Jt�w�מd\�C�I�;I�@�`��-
�Z��V��YapC�I�
y&�Svk�G�r��J�R�B�	D0����#�Z�BY�7-�K,B�T�F���3bJ��!�@B �C�	 f��,����1@]�L��B�	/b���&�f� ���"k�B�ɨ]��V�)Y���B��Ok���
�'x�3iޕr_FHr`7l�j�'7��c�g�1���BB��,j>���'����/���h���x�����'��q��(��*�(��i��'��8E,Z*��R2EY����ȓR��	�V!V(��Pj7cC�I<p@��_��ى��λ(ڊ�2��C%ֈ���S�? ��I���B6YA�HZk[� �e"O���^:R>���U��P"O ukRO\0v���4�ΜWZ�\��"Op�K�GZ~0[猕�+T<E"Or5�d/C5&*�("��I�G�s�"OfJ��_~9�':8���c"OpE`f��rUʑ���@[*�)��"O���f���P�"���u����"O�0Xs�`� ���'�}���%"O���B�6�����,���A�"O*8�v�F�O�A`K��!v8T�S"O^���K��/���*N<Y̡�"O֡����9B�@�jS4"n���"O4�	�a�QlňE�Θ~�8�Jt"O�-�Ө���6��8\M�MR��%D�d Cl�vU�)E�J�1,\����?D�(9�/P�H{�TV�6r��YSc;D���#G*;ڦ���c�2��k�d,D��j�z��vfíWk*�	��)D���Q̎%)`0 #���!ob�� K3D����"�3u" �	e�2��M���/D�X�u���BP��a��Z&N���@/D����١{g��P �1K��9& -D�D
�J�"</z�	"��3)a L�c�0D�ha�oK9
*�!F[pC�06,,D���,�?G�0̃U�����a�+D���禟����;�*�� A�-C!�>D�P���V� ,ʒ	��RT�91'�"D�0����,����6/J-1��?D�xz��R���ԃ� �F��`1D�� �@�7LR�Y����o�	2�$D��a׀N Ne$H��m;a@��+#D��� �[)F+h�&��%�>Xo"D�`��Y|���`p"<; �!D��`q��=ɪ
�BU&��T��
!D��	���Q5:i�E��_h��U�>D�D�M$_r��2%����i%�=D��y!�� H�5;��(v�G�03vB�I*J�6�Q�����sP�D�SrLB䉕j�H�2V��\@�� ��G�4(B�	*�#��@�Z*�PP�d$��C䉸-�HrE�pnTP'F%K��C�ɤm��y�c�G�B�l�8Mq�C䉀jl4P�� |BE�Ɲ�!�C�	�h��`�R�_��,����@8C��9Q`�(��[���T��G��]�C��~�Da�-՚,��ȻaE߸�B�	�r�9ȑ�0D��!$k�B�	�S�D�JP�4ЪT91�ڟ! C�I�hD�I�#jW�,���Ӥ?}��B�I�VŨ� ��N�@I�sI���B��%@nP��3�rM�wL�k�`B�	�;�p�P�� �H� q�<��C�I�2
<���J��5;N}:�M8��C�	�{H�@2�H�!-_>-�#�S'~Zv��d5a��À�s��Ej �$+G��ȓT'l<�5Eʑ�b�)K�q�ܜ��M���W���5r|hJ���`b5�ȓ?���,�p�� #>p�d)�ȓ��虶&β1��)3/9[��1��'�d�rH�]3NXЃE�'r���ȓ!m�°�_,<�s���33`����Yg�p��J�5�d0�S��	-���ȓz�4�r���<�vٳ���s��Q��S�? d�`k��u���KU.Y#�@�"O��P�g�?cV�=S�'j���"O\�#�F�o$��*ą>%�*yr�"O$A����c��g�K58�ڤ"O0e#�ƞ"b�&8A�ʕGv �"O�� WKL �)�G��v8< "O�Mb�� ��aYb��Wh���"OVa�CM/;�[@NP0h��"O�� ���>^h��"#���"O.�#�"#�����	^zzy�"O�e��,�<V�6e�d��yeD��"O�t�mьh]堅/U?7b��
�"O��B$'V'ʨ��`N^i�s"O�! t-G�udRUzE�@f�S3"O ���fEb^:(B���%V��V"O�ء��W8>�"e"�}�L���"O,t���L";�h�BZA��"Olcg���ܘC@AZ�K��y�ğa�>]��d�8I�ǆ���y"�pyt#50Z����`���y��^	|��-�%����a�͗��yr���S�B��"�w?ؔ���2�y�E�0C�x�b�kdF��TJ�y��]��M��ȡq�Q��yB)��o�PEfoQ� A"|+�B���y��A��`�@�kE�-n�uvϒ�y���n����%�P�&���ĩ�/�yBK�6Z*5 > �p��HT��yB��{�p�Jf�D?Xn\(���y�`�B��H���M���)B� ���y��B H]FQ�4I�~��Y���)�y"
�1j����oI/א�v���y� �%��{��ɧq%ZT9v'��y�c*<�|sa�Q�R �B�6�y�<�`�v�_�EG��B�y"�Cڐ��s�9���r���y"˅#�JU!Ң@2}v�ic���Py�*�l�>���O
�G9���ԨL]�<��ՕcX��'HG�% a��m�<��DŇp�,���H>s֎��Q�j�<�E�ݛP��@ �'�^��р���{�<�Ĩ�wZf�f"�>(x� �1��t�<�$��.�ノ�#	��h�m�<��E�VM,b���bL��MQ~�<y�煲��0!���
��M(~B�Ɍ��*So�Fe>Y�a	�2o�C�	�Lz��RN�H��R卒$C�	�W���0�E1y<hഭ�LC䉡xz�Yei�,s�*l�v,C)Am�B�ɥh�l��/�05�f��$6�hB�I�9N�	��ck�(�tf�+�0B�I�l���@��"	� �'%�5��C�I"������M)ي<�`@�ƖC�	�3��p��߽R� |���E4<lC�� �
`nC�p6,m�Oq PC�I<F���%����q!�D	k_C�	1+�8�Bc'X�`�q��B�zRC䉏h+��r���R���ZR]��"O,�5o!u7Fyz#��8�sf"O���%�Ήf�j�r#H�"�=�#"O��{��6wN%[c�_�R��$"Oܬ3�$W\z-(�>�ޜ�B"On�1Mu������2<�,��"OĠ+���3(�<g职�<}��"O� ��i��r}��g24@�"OTuYCꚾX�:,��g�0���'�2��g�L�4g&����M�Ql��	�'��]�7!
��s��_:}��1 �'}xa��oSL�p"� n�x��'$��{cg!4΁���*mzL��'1ʹ�r�S"5�����+�kDX���'��5BJ\�� �����)j�P-A�'�ļ�g�Y�H,T��f�k��Q
�'�J�@0�	>��L�$��g�Z�	�'OFy���@8O��4sDeإd*�Pb�'#*Y� Œ�� `��Ɔ[�vD��'ݔ�C�D�=;pS�L�`h��'PN�s��|��0�!�<��8�'٢Q0EHЇ
���"Yy����y"d��u4�:��Ѱ~���!.��y"�� ��4�ۻ_�49��yboO;8��*0-�Sg���� V�y� ˍeV`�e��R�H�a�ե�y��va6bÇ`h�ՙ�W�]L�8��'x�a��_#�*9Ie+��m��}
�'H�ӷ��?8D�P�F?^~r(
�'�n��!�kѶ!x��J9����'w8ؓ�!Q�X��a�L]�y6�D��'DD�bf![2�TH��m{b���'O(@�smJ"�&�H�L_�c��0�'sꥨ��%Iu~(s��9(�'W4�A�T�_�~�92G�yfX��'�b��W�N9~�UZ!����,��'�h`!�U�W
mzc��#NP��'<�8QKC74��(NԐz�@�'���R�a�F@��$.��
�'51����=���聯R=$����
�'i,QA����ru��։H�M�䀉	�'Z�lR%ɭ�@�[FǼ=*>Ÿ�'I�-i��4Z���˂!{�5��'��A�·C�IJ�-���1�'u@%���M>�T���?
�
8��'�$�	U�5ҵ (�0p���'��l��<�@�*W�.%�ƨ��'�B`;0�BI�j(�b��K��ps�']4H FIi�x��7�պ�%)p�<�J��6���9)la�bIm�<�ĢC�t�f�ؕB�|�� q�i�<i	��!3�P�F���"��"bJ�<uFY�#� "i�����W��C�<��� Ic��3�LQ�- QЂ3D��ԡZ�r���O.>��)0�2D��)t�τ1 ��,���1�1D���w�F(@I��c'$D�l��%�.D� 3FoNNz�X���.�|%bti,D���#��F�Dh�U�̯q:r���'D��b�� �X
6p��LW6DF�:q*%D�8��j��[��M�Q��NqS�l6D�PX�B���ۇ�S�6�a�`(5D��:2��['�Y�b��ƕ
��3D�����*���G�EU^xY�c%D�H2��uo��*�,ȖY�:��$D��za���V\.'jE�F��-D����h��Z�N��M��ʙ�2�>D������%g�azq��X�N��g�/D���VgD�c��ݻv꜇s]���-D�,	���=w��MS�	[�(����F*D�ăv����l���۹b�@K��4D�� �y1Ê�GJ��Br-K�onB,�t"Od ���B�ܙP��'Qg���f"OP0+���>�a����<�!"O��Y�ަm�F  ��N�x���"O
Ah�߇8��-3��)R�U�"O�%s���M���`T*14NY�F"O(����S6=��Y�@�	�@��`"O�s���5%���fN�D3�"O��`4���b���,�z��`C�"OR}��D�)���W����"O���Ѭ��i���᧑�fw���"O�-o�0��E3p.�bE"O$eA�Q��S�<AL+"O�I�7�� �)�6�Z�'���5"O�i����VLAZ�ꖱf��Y�"O�����j��q�j˘	�����"O�ȑE��c��̸��?jl����"On5��0>G��j�!�hX���3"Ol��#	�!Z@D�A~G͈�R� E{��Ʉ�>5qH#����gc�8.!�dڠW�t����H3s�x�P�5*�'�a|rF�Vj�*UG� ��A`�����?	�' L�=lMW� ������'��e���hмTk����dȈ��4�'t"�|��(��Ҫ�����3]N��[ Y�F�'aT
iP*D$7���~���Ţ,dO�i9���#f�H��ȓW�`�D��5��1��T��Le�ȓyH�q�ƕ+����N�b�P��t͢,�	�|i��ppN�;C��h�ȓ��hH�l�"W�p�U/7.���ȓ�z�ߢ��d�^�;��م� �"!rq�ӓ�[���Y�fA�ȓ 7���$���<�a�H�@���ȓ,�� ��>#40 ˁ�A�PEvm�ȓeB�:�m^�Dg<,ʀ����ȓ\P,4)G�<^ZQ�Љg�J�ȓ`Xf�1&ѧQ��!�����̈́�"S8t�U��9*�����	@�X,��q7
����c5E!�	x�ȓz l���D�#�y���`*�%��b�$�盌?��	���]�g����[���� �/Q��C_
ߔ-��y��c���	!�6a�E��!^ll��w����Eɳ27x(@��Ǜ |���^�te��mU�E�<Yc�+�2⥅ȓ���.�PR�����DS����"O����&�F�C���]R*��3"O�`�W���<�U�Y�WAf�Z"Of=rw-A'
�pq����/���"Ouh�&^4r��� ��K�;�y�"O$as��Z�cŀ�+��*x��"O��#���pQ��d��.\�	�7"O�@�$�56,yf͐q�(�"O8�	�2j���"#�&���kG"O~ࠑ"D?h�,h�T4�,e��"O���ǈ<PbT��@J==q��+t�'��
��(��.I/!r:���kޞW�!���;�R��]P����j]';8Q�`��H�w�O�@�J�*ݭ|i`Q��)R����'<�4p�Iҏ*}�L�3.ѶX����'ͨ�0�D@�S�O����@L
:�l��n�
Ŵ �
�'�j���
��Y��X$3��(k�O�9B�'az� �:b��0��EA�E��C���0?i�g� H�� �iT�1)h-����Ÿ&"Ox��d�D��85����>������!��4��O��T���}���s�L@	l�A	�'+6 Y#P�n��S�#_Q�|ќ'|��Gy���ѷX��Y�	��P"I��D�C|!���3̮U�3ɇ;rxԋFD��ɰ>��FK���2�'f��0thZ@�<`BH=Z>�Uy&��W�nlx�EAa�<a�ͅ�T�z��m�3GѪ�a$��q�<���"~h�j7��9+|�1I��j�<)�g��e*h�¶�C X�^MX��<T���c�[5&o��3@Kf�<�qL3b���E���z�R��KM�<��BK.hdi�v���4�a�<�4S(!�-� <͊2��W�<�6��Q֐�R�j�P�	�[�<�ׄB�X ��L��Y��W�<ٕ�;CVv1[��E\B9¬GG�<�k��kla�%�^�*b�UaX�<q���ua0����l܆���W�<�%�	@@����ߩy����'LIL�<�Q�^�I�A�E,�?b���0�_�<���̜P~$K! <e:81��Y�<�W�Ya�*���AF�#�؜P�R�<��Ȁ^,L8J7e�[�\0b��M�<�eʝ:�\Y)���7cr����I�<)�n�����1W�������G�<)'�'��$p����Y�aa�n�<aV�ٌX8I�Vl��)�R�b�4D���B.Ѽx߾�#��I�h�Bp3Q�&D�|���<D0�%�dɆ�;�b1kP�#D�<H%��TL�'D,N"�:�?D�(�O>@�Txk� ���Tq�<D�H���9Ke�%:�G��)u�T��e9D�$9��[D�
��tf�J�bU�!T�CO42Z�l`��=
e@"O�TBs�
dt�nL|m.t�P"Od�c@�Ͻs�6��#>H<^��"O(�j��^!^m!&���F�x��"OZ4�d�o�6iz�a̻w6��+w"O���a�JM`P�Ӈ Ǽ,����"O�Q;�gO�.8	+��/y2X�"O��h�iģ��˖j\�͚@"Op(;�)��]7~	@�@��#�|B�"O�!�%��dţ�oI�2ِ�"O�,�`G�M�F�ɓ�@a��)�"O�h��A�7 �[�n��
���"V"OvD�7���Pp>̢�̗�9�|Ũ"O�prC``�����K��V�Z��0"O
q���]���Ұ�[�*�H��"O(�;3�A"v�ٙ�K@ n� `�C"O0�� V������E(G�u�C"O�"�A·����p*��1�Rp"O\�Cc��
z�9�I�	֚mx�"O�!; ��:��@��J4�� �"O�L�%�_��Z�D�o:a��"OЙ%��M�0��2��S{j`{"O"}�bP�93����&^yR�zT"O
����A:E&�	C�Ą,a���#"OHȑ3���\�!D����Pp"Oj��R�-_�����T��2I�w"O�0E��r�y��5��CV"O�i��
7�nY1�6����"O�h���I�0��z���|h�)E"O� ��І�Q��"K�qB"O�t��H��𜃂� 
���!�"O�`��	��4�7
�o����d"O��;�X�~�N��C �>�A"O�qnH&|{6��W��|K�"O�1��"��f�`�S�@�ox>�X�"O���ae8�*�E�=p����"Od!�`I�2�����,@l!��"Oz\㒄�dN��)h��Z�"Oޜ3�W1 ��ѱ�[|O�e�"Ohs�.�
J��jF�ODcȉ0�"O�eC���`��,�u �38]H%B�"OD��Q�_w,"���̻A�H� "O@a2w!H1>cv̓�w��,z��'�4)������u��SQ�H�.`|���+{�����O��$�O i����O��D�O L���>�1K��42|�v�N=Ujphe�I"��䈰��гq.� V*�hEj?P^�YZe�3�����e�jU:�5��L�>�I*	L�(Q�A5m�*�kۼE褕2A��M�����$�O ��'Q)��ڋc����al8*|���?a�KV4t=� �L�|��D[��T|?1U�[�+u��U�l��J��uW�'��Y?U�tD��K�\�E�5%.�ˠ�]=&,@��?Y�I7�ό$H~xؕ���\](�1�� :��	��!x��B""�:X�����(O:�§�12 [qd�Mm��Ů~Y�X�F�3�%z �V+Ѫ��A0�(O ���'��7ML�I�	G�� ߗ[F�i!� O��X�%�۠V���!�i>�Dz��D]�h`��H�2`Ea��p>1װiCx7mz�Ƽ@�#�=x�%ұ&R�7�Jx��O�4�,��,�8��<ͧK:�F�x�!�L��y�Ƹ�(����:4�E���7��(
ڴU�@c�&�^��� "2���߭6.L/NX�p����|�ꑘBDk�`�&�ň��YPɛ&!sd�`�*r)����Af���k,�r���Tʖ$���YR�D#4]�� Η�?!ĴiNp��?�D�ܴ$��o��s.\�7�s�t I��'EBR���	G����DSl������$K��p�K�8�Q��B�4ۛ6�'�6��Ot��i݅�B��
%�8��iߪU�v2 �]��?���v���"*��?����?���Z���O�6-D&2z��/ӱ&<�0mҢM���� !���.S2��&�K�.�?��3��<��OF< %�Λ�
պ�TT�v�@�FQ쀺u'C{V�S#�Ɇc�"B�����PfL�BdW���G�Y)e�֖�S �I��A�k�ɻ4!��Dc��$���̟T�'��}��-Dt�x��u1lC�{��'j��r�ڨva4�3� 6r�T�C#AIئu�ݴ���|��'����(V��
̌WL|�
�?b��}��$��'�����O|��O��2�j�O���O�uJ%�A6s�4Xypˋxjx��j�7ku�U�H�V����*��eF=l;Q�V��c=�EK2�]�X�z-*I��44�H��fK�2H�@|x�;z�T,Dy�jł�?�QK[?.^��a��B8h�Ձåew����i��Q����{�S�����9�xL���L�)YY��C��yb��&X�x���עd��3AdM=F2�$NŦe ܴ��$�(��tlş���K�D�V�QSl1qS�D"\ :'�E�$���O^���OL����Ox��?9���K��߀ ��}��G^�{�"u�t�I�z��9iĄm��c?-�T������G*=򐑪W�3�X��Q����M���)U�S����Dh�R��!�s�8T��d7|O��wr�Y�2�T4\�q��,s6����MCA�ip�V�T����t���bw
E��#9��	��	@�g�ubf�� @�?;I�$����yrG,C����#ږx/�d���L5�yR� �2ڐ�k���%
.�֍��'�^}�� �)���:`�I�^�t���'\�!�P^�2W/R�P���	�'mtPD��[y���p!P�b�'.�x�//]b� aÃ �l�h�q�'	��i0�S�'�)C"�p���j	�'�X�v�r��}+2!M�b����'�
�x4ꒂ2���#�C�.m��b�'1�����:y��I1�(^����'���ć�:Y�$K�dL�RvZ�'
Bm��׈C2�1�W+�w5���'�L����ƲL��,!��P�k�V��
�'�3s���=׶�1w�
!`�i�	�'�m�D���|� �*�JA�T�Z���'W�ݒ���#\e#�i	�R%�Q�'�\�p�M�d@`��	W�,�b�'��a�,R�M 0�DaL���	�'��iRL�$-Ԏ��,���*�{	�'H&�8v*��5=nŊu�L �2U��'�(�C�^�|=H��tj���m
�'!ttW�^���M���Q�|׈Lz	�'@X�p� ����D�m�~U�'�>l�&h��L� ���
�.���J
�'^�P�9�x1!�h�.2J4���'�3�C�8F)�d�t'�,m ��'�TyudU�x�T� �u����'!�DB��ҠsPΜ�ob���'oB�+�K!
ۂ�!���9E�<D���	B�R)��$$D4C9�K�d:D��KQ#�w|��C%Ȇ>J_�ab8D�4R��E+�~(kC�ثF�}�V�+D���_'c�48� �S���`G�+D��5�"W�BapQ.U5[l܉�Fa+D��bM�6���f��xh�e,D���e-���M��d�-u�J�*D��ho'$��ө
�@�(A�G3D��k1ߏ<S��sG�V�a�`L2D�� ��ۀ�>5�Ft�w��';����7"Oj���.MZX�Q���r��U"O�`Cpn��3�V9K�F��?}�EH�"O�����x���K�ef4a�"O����AY�Fَ@`a�϶pG� b�"OE����D�,����'�"O�����T��U���j,c"O~ 
q���hD� �#휌��"OZЃ��9��l#g��)��=��"O�����Yh�= ��:��@��"O�EqB��Tֶ�y��0w�4�v"O��j��@�,5�fh�*H�4��"O<4��@�1xC�q�U.�7(��|��"O���H �@_�4;s�R f�`+�"O�4Ѭ���E�L֫a��ٚR"O���b��^���T� �u���"Op4�%�=V!B%a_�)��Xr�"Od��	��0Q���(��A��"O`{'�C5%�Yza39��9q�"O���x�9�o�o��*�"O0,��-I*:�&���94A���"OZ��#C=�Zh���#"\�@�"Om���'>Y��)���#%�IB�"O�����5l�Y,�2���0"OdTȀO�������M "O�9 �@޽U�h1��m�$T�p6"O2"���g�d����
�\��āD�'j�d�l���2��m�z؊�j�<N�Ix�����曏l���@��n�&E�q�&D�x��FE�#�2c��W<�	�h%D�l�����5Ę}�0g/]>�щE*O�m�do�0X��˱	�1Ԗ�Ӗ"O��r��r�*iY��A5`^ )��"O� �cYNՃ&G�7F�9�WO�$�Ҫ�-
BP!��f�b��ǣ<
�V��c��F>j�T��Jԥ#���6��=R�q5��$�*m~%��c� 0b����p��5��[Id���D����6�Ab�H��c�u���ȓ=���v̚%V�.�ci).�m��	�V���mC"z����p�X&�4l�������Ȕ�F��%he�E�!ni�	q<��m��C��O����3O�̰ل�v�v��2h��s{�LB�O�{u�ȓ>ް�/Ϧ=@�"wB�wp�A��W�|��ANȆ�%xP� 5/�j��ȓS�h��L�'�(e�2OW�|��u'�|R��:tx.��c	+7�4Շ�*���h'��[���×)%�꽇ȓuN�`&B^#��)�$Q��	�2ms4��`x���j\�~��E�ȓJ��!�H���P�7K��9����n������r{ru���9Y ���U��2� f����5�ҲZ�Z}��W�=��L�-@�C���.!�����a���� Q ��`�'���ȓUձ�_0x�Z��Z 3��1�ȓR��h���׏�.��B%��=���ȓvgY3T�(rz������kuր��"��rc����$CJ�Ң�ȓ8����BES�����	k����ȓ(�
ɳ��ݎQ�l�Є�:;�L��]m,�V�@�W�E:2�ۚZꀁ��Lq�+v)ӉZ�$5ja=K\8h��S�? ��AS O%�Ιh�N��-���RE"O�� "ڝs�>i2�@�.0|:"O�@�U�v�TD�A��y-�R�"O �[��Eʠ*��%F�2��0"O�U2%�� \��g�P�jh4"O.%��<x,�P	��|�T��"O��H�N���|-�<��oȒ�y���Z[~���*]67�2�����y������҄��@��t:3/A��y2�A  P�D�=�~4�#R��yB@ʢV0�l9#)�+7�	��Ô��y�d��0�a)I�!�Э2alӭ�y27's�0�2ܪ!n�������y�ϭ*ib�9���j�ц"�䓡0>	#!Yb��:qP�`8,s��Yy�<)�c��4Ɯ���7���2���u�<�4e�)�)C�L�;~���V�Ii�<��C���isR��?Z�!�ç�e�<q��ڄ/VHE�U�T��i�<A%�*G��5��;3���g�b�<i)a�`�D��}9���ZI�<dfOF|-�6^�'*Hh��^�<��J�("x�B�x���Z�<��C:|GXj�	H�=6P��F)D��H���>ES԰	R��#�:���*:D��hQ��= B�y#D�-̑:�(:D����B�8D�� ��#?Fk�,��6D������<(pZQ�f�66}��RuM�OZ�=E�Ԋ� Hh��K�I�e�4@��!�$�
A�F,�5��eO�Q�nN<�!�]�b(vH�4��ᤧXC!�$^7ynIrdCJ��H3ں�!�یz~�=�g��=�ܴSV���}��H ���?�%�G��e"6�Rd�*D�x���+0s��c�
�[������(D�tJ�n٪Ur^-+f	��0�Ry��1D�|;AXV��L�L�oQ2���o.D�t�!̝�l&J�Au(��ڠaT�6D�X��lW�Y�M��'O��D���4D����Ј2ۆ�9�o��M�~|�T�3D��:�����\d�V�B&7�� �f��OΣ=E���!Z8k����i�j�� |!�ӪxBܨ�3!�!Nl2Z�*&^!��?{�8A#V��Hw�m�!�-~e!����V�@A!]�`{�U7"AI!���n�|�"c�_�mwp�V!WA�!�N2s�v�) (]�?w��kGO��!���J��gH�s�Ա8�M��g !�J?�F��`��'j�p#�V�!�$N$x5�d��=jn��+RdD�!�D��O������D:�<R����q.!�D�g�� X3B�-~t�&⇆0}!�D� ��JfaD�5"R�����!�$Խ6�ĝ;��B�Gp�ïϦ^!�dְe;@y��m�=:���`�܋V�!��P%B��x!�ǺzR�����S�Ku!�d2_s� ����w�H�V��hW!�Z/�� w�ӽ�z-ʤ��!�����a�Ü0�Jz䎏Y�!�d�/_�"��+V�z��yą׆`�!��8 �Lx�Ћ�:m��He��!���A���`Ϲu�(���d
�lX��)�'p�.=�TˋH�� #7�^��\|!��d'�&�	%f7Xܐ�T;] ���"O� 5)�M,0tIҁ��N�%*`"O��C��"@2l����\XP��"O��ؗL�Ak԰bÆ,��&"O�(`1ʃ[�� �`ȗ"��Z4"O�(Xsa
 w��"���l���AV�H�'J�OZb>��B A�W�����_ #@�a�C8�	b��4!è�yR�P��C�'M4�Es$�!D�x�q�Ɏ쌱��`�%�l��Am!D��"-	�0�
2��oL��b!D�<h�ܜIX8�%��9A94�<D�\J�F�䎡�s�<0����"n;D�,"�ͱ/���1�nU�.��P�k?D����ʃN=��r��P�'��C�*�I]���q@KN��A�!1L(����:����'��	9`�����h�K̈́�K��;��\�̇�	 >�3b�]�h�n�����`C�	�$.d�K�Y����� B�	�-�b]*ӥԇ͖�� (��;I�C�	5"S��W��?A��0W�<>;N�ONʓ��O����|3X����W�)6PzQ�Ed(���3�$�<�|�O�e��o� 1���U �<�� �"OP��v�ݐ?J�@`�$@<�� "O�1��ͤ:;*��G-o$8M�E"O�a��K.(��,Wy|��)�"OD�@cO�W�P�� .A%yp�0��"O.�"$��l����c�2e������'Yў"~�b%��B2}r.�:�8�	�f@$��&�S�O��Ā��
Aq �����U�Zȹ���<�+O��S�:,9���9 1j�:W�%j��:�rD�+tNHI�� �����4D���隩a!>YR��.C���dM&D����hK�41���)x�|@��$D�X�jׁz_������l�>��)�O$�=E����9Qh��m��p�J�GS�X1�	W��(�4�2bcX�v�� �'�8J�:,�"OBm�FJ�h�ք�5�@�-sb���"OF�ҡfƫ吤���2i�]��"O|�I�-5�m�r��yI���"O�;�m�>t�b��1)P�W�<���"O���1�a��$)�/q��u�r"OP�Z6� �4��2HH��(�"OF��΂G�.��� ��b�����	jy�T���'M/�aReaT#�r�w�OE�=��wy�'ɰTڑ�׶DTaBP#�.���'i(��Ћ��b��Jd�AF|I��'_�1(u�ǔr�(8{P��,k�C�'��X�V�х/{X0�dn�#0i��'������i(9�Q���KF����?������y?�!:�b[���L�:��B�	5!���� O���1I�[I�B�I ��%q��׊B��X6�#lR:B�	�F��yH�$�1y�pm�����4B�I�~򶤻�-�#LG��ϐV��B�I=I��QE%0�}��B'7f�d�O���+��(�܅��쌉J��5-�>k�(�IY�����B��.��X��l��kV��3b'|O���y�V�5F�C��A�rfL)R�͓�?	)O\��dVG�U���\�\/�=�&�ݝF!��f�0��v�I>	�����F߸<�!�$�/ |
�lT�}�c�$/�!�)�N��h������'���4��)vy�Qm�?;��y�B�w������fk�=J��d����D0yEB��\��BG�x�z�9WL��B�)�  )2�c�"��C�"��>ւ�"O�T�Ї�8��ҡ����$	"O"�I���@��`⠇="�p�P�"O�A Ԡ�2-�xX7`�-l���D1�S�)߱��}���6���Î2!򄞳/S�7��(���l�>jџ|�����'$�Ʋp�8d�c�L��bx�!����'�a|�n���Z����bj��'"��y��^0"� �Y�'�i
�XG���yR�ض#c��1V��o�b��cŇ�y�fӦ���Q'F�tp�W���d�<)���[�>`�m�EAK�F�D��OT
E��O���d��N)򠅵�>�^r������O��.§u�6��T�\�]T��k�1yL����u_
m20�ٲ1ҺD�l�CmNx�ȓ�^��EY��Yq6�,-\���Uq��i��4�����Ս ��؇�b	��(�<�b��0bR'����+PbQ�(��9�����?w'�l��1	@5Z����*�g�S��P�ȓ�f�`#	3a���g�N.}�9��J�L@�"]�Af����q	
|�ȓT���a 7@@��j]�id`��ȓmX6�ٲE��e��=x��t{���S�l�J�E�6��QB/\q�<p��y]T�"'E�bd^�Z3�[�"p���Q�0��O�Y{v�����$E�ȓN��R�U>E�49��	� .L�ȓ@J��3v��A���]����`�n9,~��%kQ9(d�CF0D�P�āŊw�Q�q�j��q	�.D��rLP�����N�� ::�H&e7D��h!,[�u���dC:\82�2`	�<	�\��T �p���6$���y"O��B�D5(	�tb�C P�lӇ"O�Y���R S}��Z��;s�ՠ�"O�m�UB���jC�ժ� ��"O�@�i�9 c���0]+s���"OҠCC�9����T8��8v�'ў"~��֪B5V�هÕ�O�q9a�V�yH�,��F�6(Ɯf�K��'lў�O�B��I3}6u:���8B2��'ŒaJ��L�h��r�Ávu6`Z�'��zw�L�hV� �ҫ[o�j�p�'��h�j�{5�P��ϯ_���
�'hzE��"E�I1|Q�q�&P��ɢ�'P�,c$M�'�n�r!�J"Pu���'b�%�7^��5�� >���#�'}�g�Wu\�)	�-�x֌�'�J��H�|_ּ�a�BI	� �'%�,+��%8Z(#�cN,@�(�'*4]��/Y@��`O�>}��K
�'<6�x���x�C��6L]b	�'J922���H�K�=f&5ZʞD�<�ȋI����Wc��r�zm���Y�<Yg�Ҵ#{�9�聀+L�aZ��U�<q�����P!�'G�n ��H�S�<��$	'����A�ه/�l�Y&G�K�<�VJ9�(��k�|	�X�CRI�<Q%��F�"���g��L�| GK�F�<!�ʢ�e��#̑vz��:�d�A�<iE�!1B,��ӥ���2�{�<�6I� |H�����K�Nie� n�<!���n�|�)[ x�)��t�<� f�r�h��0s�y@�>�EJ�"O�`��l���y�NO�_%j�X'"O`-"
ݨ�-�G�@H�D"Ov �!A	AI�\�U�RҀ���"O8$�V�T5f��Q肏��5�8��D�OH��$�2����A�H?�^���J�0�!�D�-��m�A.ߏ��	W`\R-!��8�l��e4���Io5`!�ː�:w�<L��8!�-�!��ɥzg$]�5C�z:���3-	!�d�!}�*���#��^w\�3ka���9O�<���_()PzQx�-e�L�R�'s�Iڟ�����$ҿB��y(��K9.h�tAիň�Pyb/�=2�A�k��2\��I[�y��ȼeBbo�-IB�̛F��%�yB�IeNu���P:4� 	� N��y�(A�s���Zr�.A��8�0�۬�y2��
�� s��I�b1��r!��O��Ŀ<����t��:X@�tӃ \�^����Ҡ����<	/O@�--����� ?�i)H�k"O� y�B՜CG�Ae
�1�Ԡ�t"O�����j�����HC�1���ѷ"O�!��BG�;��b3'�q�
�(�"O��1�ƒ��E��1D�>�c�"Op��c�T�G�$��u,�'�m��"O�L�oC�3���R��:�4Q��"OZ�i���T[�Q���ް��q��"Oz���*�;'2|"�&�S��r"O�0���YE��y G�Z��"O�RuF�5Yv$K��ޤ�x]�"Oh1Ɂ˟6�Z����ń�6�St��ޟ�D�t�@3�n_�4����?�I>i�cB&�!��t�����C2Eʑ�ȓ�(C%�
ua8Ńu��*Vt�1�ȓvgB��bf�J]ˢ��%~?`$�ȓW��IGb�$ºq���$HƔ��d)6�Xaf�+.�`	����F)��0�l<�e�Duq4`�1E�q�`���p�'Lth��h/TT��ڙQ��L>y*O�����#lz��m�@�!Av	,��O�D*��9[r*V>c �)�B���XXke"O2��Bg�	i�ɹ���}��[�"OJ�T"��2��ű�L�=̼��5"O���t��&���(�j�F�ڝ"O:� fմ,��z��өF��H�G"O�D�a��EL��֋�"�֑�T�d�'�az�#��
&�Ʉe����́>���?q��0|2��&���aԅc���RD�o�<�Í�~��B��I)��AĢ�B�<)C��Z`\��aLE
-.@q�"NB�<�׀��s�TѺq��0���d/�s�<��Hn�jAؑ�+&��Y!�m�<�Ɔ�.pմ�3���wB	�ā�C�<Q��>y1��X���X��`І�Z�<1��ΦYj|iP�Ju� ���O`�<I�b����8p��ƒ`���x�<�wH�|�<�����!;��$[F�N�<I@f̸;��e+ ̎�J��R�(�M�<aP��6K\q8S�Ж �hP�PP�<yT�e�-�LLn$��nP�<y�.�$m��d�c���*F�A�b]K�<�[ `@(��	d��8s�˛E�<��,��s@��4��V� C(BG�<����n��%�bE\�j��A�*E�<� ^T�R� !a?n="D�B�ʴ"O� �&ʌ�v���L�L�-p�"Or����g(�0m�`����"OXz�ǎ2:D9��,��q��<Hg"O�i��Oފ>��s�I�M���hc"O:�J��E�
��!���.p�J1�"OܱyV�U�	�n4��I��1�:��R"OB��Ëъ�L���}�^ �q"O�L�eG�1 JUqf�1�ļ�"O�Lp6�>���Ř�cKl���"OzY�b�݌k��{A�KBE!�B"O�s�iI*T�ԠksI�I��I��"O"u@����?�eI���0#��`�D"OX�u�J>5ɬ��ƌ�n�2,i�"O�(0eʆ-��af��<n����`"O���g ��Y��^�@A�"O�����S���Ve�c`4���"O�y��!����pz�cߣ�$=w"O��i��Ǉ:�d�;f,M*u�)s"O�D�3L�P���8�$f�q�"O`(؅c��X]��)�K[�J�w"O汣���'&��R�*��i�B\�R"O�鑕M^0Vg(�qb	��+�dU��"O�1�0 I9;Cn-�1	�}��"O��᥅L�2���U�֬,Ԗ5�f"O�$���Ed! ��0s��	u"O��a`��Q}��g�ѺM_�<��"O���S�4��LӀ@S�,Ml��#"OB�����. �N���o^@j�$�"O
غ6�N�54D�x�̈́�Gf:��"Of���%A�pv�`�.~M��;�"O�l���\tqA��A�	�"O�i� ʇ?�\RG��$�\§"O�EꢌB	��$ Gc'^�#�"Od	y��BL;T(�!
�+l��W"Oz�w���M}X���oG
Yf���S"O�<��I�?B0v��=yԉ{�"O�hSs&BR�\����,o;��j�"O��BbNoDȰ�b�I�s��	�"OJ ��A{����b��0�6ͪ�"O�d��&�&����%gؠhGh�
�"O�,S���9�A`3��(r��$�"Olx�� R�8�t�B;t���g"Oܠ:�M�OvB�e��"88�b3"O�=�,E�;6X��ʇ9<p��"O8Yt�O�(��l!e�3c �$�"O�$ʇ��� ��j����jʱ�"O��i�hۭ&�8A����.b �P�"On�"��V )���:�Rl��"O���4��h���88�'H�-�I�y@\�J��E�R���',
QЖ�\�f�{B*�;kV�:�'�@��˷sk^U�ƌ�=_<�Pq�'��p!S看R<�xa$I"nR���'(���A�
7�d��!( a����'V�X�wL���nd�&A�2�J`��'4��b�وk��S��4�h�'N���+I/��Y	)ɿ�b5H�'߸���Ţ\QjA�5�I�oHA �'�L5��x����uJN�QJ�l��'�H� �74��]�s�NxV���'HHBc���a�bL6B����'El�p�ÊDSpy���F6�Z@0�'��-rTd<����-�2������� ����Z�582�(F΍�uZ*���"O
ź�B�	�d
eG"S�-"�"O8 A�B�9$=��¦��4d9	�"O����%i<.�����NVe��"O�iRc��3�X�h�i�;EK�(;""OJx4m�PT)�1sA`<�R"O hZ��γ4n��!�H�;6>f��D"O�u���ܰJHf�Hd�\J#*!��"O$�� d�$x*�ٰ$�A}�<A`"O$���暯
��� �%^�9+Q"O
(�fl��;I�yY�J��
Q�(��"O���O�Jn��ђ�gJ��"a"Of�*W"Ʌtm�h���)A�|��"Oh��A��	��5���V"��B"O�ub���"3u�$���#O����"O,q��Q#Fس�F�2PjM "O�p g��\.)�Dl͞B4��j�"OP̛���ݺc�94-�]k�"O@�B�۪)WpT��iY�g�hÕ"O (��e�$e�N�0�{Ji��"O^�Ca��-�xl��H;t���"O�ic���B�K��7h]0d�#"O$��¹�D����s0~���"O�t��P��*�e�?�ޥ:W"ON���	F��h��$�� m��"O���STC� ��
��H|bQ��"O�Xf���X�a�T�a~�"Or`�� @L��k�0TBA*�"O(k3#X�?�T�g��$O��W"O��Jψ��`��A�	0a]P�"Of}b���n�R��F�Z_$��"O���p�O��U�0,˨=x�lu"OF����]:!����ɜ-r���f"O�mJ�s�4�r`)YB��b5"O�ɩ���f#$�Q��d��5"O�HB!��j�!��!>SNm�s"O�5�� U:B�<��M�YQ��Af"ONX2Y�80�,��G�F�(�"Ox5ۇ���;yƁ)e��\��x:'"OR�"��٤�%/�*+�|es���y� .pa@�+�޿�J5��@6�y�O�
H�+�S0Bj����y".>3nf#�(���EX��y���! �'� )�y����y2l2���b��v|qi�[��yr�͓3�������0�y�gȿ�y.�J�A��Ȍ1
f`��
��yBM�RB�ձ��W�0�����yR�D7B2�K�#o/1��gš�yg_�8��h�!(_�FY2���yR�ڰR��d�2f�P��A L��y�C-w��1@
οv�><
aȇ��y���71}�uh��Q�i��uH���>�y�MԒ)�l	#�,�"e'���K��y��ֳ\S�a��
)s�R&��8�yB�K 8�����y*l�Tϔ��y�JK4I�,���f��J�;!���y�	Nq(� !(])����u���y�e���e�-���i:(<
P"O�Q��٦b�TỡF�`:�9��"O�����a�hq��Ե08fL�"O*�jQ�/5�|'B��%8@�v"O�t���C��L{p@�+*(Ry�"Ojz%�F���"�^�K!�U"O� nuCS�R_w&�p�� 0�84"Oz80#L�I�d�l�v DXU"O�D���Bvo���':lU��"OD�J(Vl	bc��RV��d"O��:�y�:�	T�T� 
V"OL�bt-���D�'គLr�X�"O�-ې��}��8@t@����9 �"O-h���As8l�6���2"O�e����0A���3 Бs�}��"O�qU�טq5j�e�n��D+3"O�t�F�$̨X)�H<u��i�"O"��'B�T&M�@�
�L��AT"O�����r/Je��ǉ�s�`��"O`�WB+H.�l��h�>�&��"O�ȡ��Q7Z�H���h�h�]Ѡ"OLi�"cBt� ����!S�hm��"O��p��:}x0Yb(�� �*2"O��S�B�?_8hx1�΍:Y^8 �"O"0��i�~�`��#�֚PM\0��"O\�3蔊Pe�d!O.���f"O��qcW8Z�<�qdS<��Ъ6"O
i ��G��8��G!�2ۂ��Q"On�����9l*t)�1&��}.f-��"O���+��d�N�J2�ϑ`��h�7"O�T���"unԁ��Q�U��I�"O�m�`�&EV�A1��C#O�l�"ODH��dUca*0��F�.�6��P"ONڑ��!��Z�EE(:�԰�"O�A �]/N�s��L��\��"O��B��:D�6���I�+u���"O�	W)\�	|��"�Kp��"O@�� �X�>̻$�ɝ=T�h�"O�]�&��G-J��,�V�zE"O��\	Q�	�K���rI"Oj1�ۖ&��,1#� (�"OTD�b�G��)���.0��@��"O�ݢ�#��`��Ԃ˺M�6�Z�"O"�"��Y�P̼	�s�0q��AC�"Oڜ��጑k�4��鉁;�(��"Oz��`─�!�n��L4}�a"O�<J#��#+����L,)��C�"O\�aԄ�N����B��?��`�"Opl�"U�:�V� B�'zȭ��"O�h@�I�90xU���M��uS�"O�+���@
�Pu��v�J��f"O&5"k�ԬK�EC;�Ёړ"O��QHݕ#�(=�ccR�삑8f"O~�p��ڀ.�P�
��ω �ˇ"O����E�I�F8�&�G���"O.�3&P�,�h�(4�RO����"O�[&���<f9��#�*��C"O�x�0e��V0r����F\���"O�- �RdG�C.1P�mz�"O�̂�N �<Sfm��B�@����"OP��"�V���qi��A�ϴ�CF"O�a�fĪByJ}:V��+� �"O #$$��6R����M
�`�|��!"O��w.�#"��BW��:`�B�z�"O�y�-	�"�\�0ɂ��	� *OR���"T�vy7�\:H�vLc�'rx
gO��n�!;�HA�z�ݠ�')΍�e����HZ�O ��@��'=p��c'�"8�ܬi�H�v����'�"��̖D&eb���#i� �a��� ������
ʎL!�ۨ�┈�"O�}��F�C��DRR+]�?4��c1"O�L)�.�]��Q�W���s�"OxYq�IQ8(`(�HvO4aZu�W"Ob8�'-�0'��Q@�	�4��<��"OL�/M12}�7e?U��q��"O�;'�ݣkodX���>�e�w"O���P.Y�R�J!��LC ;�*P��"Od0���F�ec�h��5.�~8��"O�`�5�B�	������6{J��"OݩA)O�$�xer"�s�N�8�"O��ʖ�$YE�K����nhp"O�� 7g�0W�`D9��`�<9DF{k�iU�Zھ��h�]�<a����� ��љ��
�[~�<����9��u��ǭ
I�p�AY�܆�e�4uʧ`F�MZd�"tڗq����=�
ۓ���q ���}��L�XF�ȓE�2M��c��:PR$��)���(
�!�_/]��<Bc�R�L�"I�ȓ2���@���?��t�T��T|���/P����ˬ&�Z��
��T4��V�p-xa�D]�Ac�g
@��ȓUZ�g�C�:�pR��Ҵ��H�ȓhjE�D[�3�5�q�0a����a�<壴��
�P��h��+��W3�`�l���Y"��C�@�j��ȓ���ኡZ��r���&LsZ%��**��gd�s憬a7��"4��1�� ����U�� #R�e���kHu�ȓ+��8х���ԡS�^e�y�ȓYz|(D˟��d=@6���b�ȓ������'=��h��ʓ+��M�ȓu`@�Y��Ikτ9���n}��������73����v�֘(cl��ȓdȜS�/�3}�,�x��V�,aP�ȓA�U��i.o��pB�F	]���ȓ!;l�D��WF\噐��D�H�ȓRj0Lz��X��M8�jI�+wJA�ȓ��ـ�
5X�P�m�59����ȓ�ʹ"g_����mJ�(V�u�ȓ(*�U��
6�r	�
E�6�����	� �Bb�(y',�,&sP��������N�FS�je��+���ȓ$%q���
i,�ց�1=��ȓL�n���ϰ9R�LYíҜ&�z���k����c�*  4�*5�ٛP�}���f�{W�I7rU�-��狚@��D�ȓ��`���FN�uR�I�.��y��&���֪��T�"	rn�=�6���VTZ\� �v"��A�iH~��P�ȓL0<m3e���p3L� Pe�r��؆�\��)ӀI 5��(5��-(4���7��q�e�2��� 1��؇ȓ�ݢf�M���9�H�Fc̇�~LT��mɎL_��P�%�&
.�ȓ ����`"�DUށR�Է!J���'_ў"}RBc�u�$0i���b�C_�<��V<�)r ��
}W6�j���s�<�$���(�����㇈P�pªn�<��h�\O����-F�8�~�[�N�U�<� � +U���e�N���%�DW�<��OF� �ڄv+Ԏ&Nڼ��M�i�<1� X��9"����+���	�G�~�<� l�Q�ND-cH��&��3=�>�I�"O��k�׻F < �����"w"OP��eK*qڈYi��#���g"O"5iFf��nm��ң��9[�	��"Ozqӷ��Y��l��K
g���"Ol�),G;$r��ň߈ N�i�"O��#r
FSL��9r�Y��K�"O�p���W�h`�g�)�V�� "Oh�)�6w��,�$��.!k,H�p"O��)_�tD�������F��	�G"O
�
VG_F	�0E�D��p�"O�X���ɍ,r�=1 �6�8�y�"O�T�pC��Uؕ�^�e��ͩ�"O"����?`(EhM�1:ꕡ]�D{��)� &�(�3�����t�k��ϓ&�!�ę�M"�sq�Y��"��4�Z��!�$� 'a���P-|����ƭ�	!�DCdVF�@DՋ8��R�� �!�FU�t��A�+'�,A;g�݄J�!��
� 4 퀠蒲1'���6��4�!�DH�5[D}���X���|+f���E�!��G��5�d��3m|6�{ .L!���e����A���N!c��Q�g!�DًwhR�bQ�a�j��!�d�<WSHa�1��/H�J�M�&�!�d��$P�u�w#��:d���M�U!�� RgV��R��0 Í�bmP�!�d�l�$9�!"2.�3f�?m�!�$��4� �3�n٧i����HΡg�!��5J����6V�L��� 
�!��Q(��e� ��jRsČk�!�dM�k�>Ƀ3���c��e8�AGm�!�]e�;f�,�X8��X>v�!�$�	L�5i�|�T5�#̐"�!���azFYs
-o��hu̓�1!�d�9e{T0���*@��� N��f!�Dіu$�h���<	�ڱ���X�1�!�D�;D�oD�������!�dY�&ZmzF��sr0�
�� !�D�54	*|+�̃Ph0pٷI_	!��5�����ʛ^����cI;&�!�d�'�N}�ƪ0�J�A�)]�!��/;_����Be_t�{�˳9�!��>�^�(�
�[��K=7�!�"J�*D�0F�{����1f�,�!�Ă�MaQFF���V��6Z�!�Px818�CL@���ڄ؀H����ܮ7��,��A66�I��(�y҄�|��D���@�,D��́8�y��Z��D�it�@6=!�����G��y��[4D(�&�B�-x�aA�f���y��+,޽��.ٔ�������y"� ,�lHwnX�U��"T�:�yrL^>'����hR�Q*.�p�敲�y2l�h©ȬQ�ܩr�K��yMڶPӖE{�Ǖ�:.r}�D%E��y� �\�a+ى4H���@��yb�5��\�@�K�0IԜö����yRg�("�Nh��)W�Ĺ�4�س�yb��#��0����S�X1P��A�yRD�5
r�+4�N�G��`�����y�j� �pX�v��v���2AI�yBNR4�D8j�\��"�ח�y!\2d�5��T�ŚV%���y
� p�2�һ,:��{�g�"¾$#�"O��)ўI��෨�W�	r"O�	E��6�|�
�Ʌ1T�"O8�����FdtMВN�oE��1S"O u�Ca�7م�6	 ��Yp"O���Og�:!�L&O tp�4"O���L�K���׋ǥi�RuZV"OF�S4�� G�x��F,)�$�x2"Oz!z��%m��L<Jf���"Ot�
6gE�HA�ʞH8��C�"O(���bΪī�k�#���"O������& �����F�¬c�"O2�p�� æ9�eI��Z���"O��#��M��uI�g�{�z�y�"O0��2�{�h9+Ë� K��	�"O�	��P�P��ʭZ����]��DP ~	C�I)rF���Q�D|¦ۃ6|���S���&��*'�y�H�(./��ѵ��l�u��.M��y"�%"|) �t����*dz	�'�H("-1��h)�b�3�`Ճ�'����Q%Z��1���=glQ��'fh�8Э���dikI�<k��9�'�謐2^�X��)r�A�1��I�'f�I��AK�Gh�$��)��`�'SD%!����<ÃF�*-��(
�'e��z&/C#6̸�%R�R��ic�'��H"�B�/cj!�A��>��[�'4��r��/l�����"�,m�4�
�'
�ٚ�m*Mu>�`#�%����'Fr`I0@�#ɤ�j3-ϼ����'�@d:e���b z��2�4�-�'X!��O�:H���2#��~h��
�'�Z|�Ńˌ.q,!�*%v��L�
�'A�))����S��M�u$���'��A��\���q#㘎p���;�'0���b&Z	>���AhD�8�' �a{+Q�HzH��U�8����'Q��2�#��.V�0�N�&���')t�Y@���!ڄU�mإh��(�O���[�J�j�3@ %�'i����K��}$��Y	G>F��ȓz�ISU�%���s�_�pԱ��4T��d�=e���l�]�3�	�$l��ӦLq��t��KH<jH�����B����7�ҽs���,�:���	a��0�&�[p��(�������{S�ٰ#o�1_mH"6#B-��tCP�3r���-擁iN��$�3VYrL"A�D�*~C�I�MC��CĂ˔]�+�W����<E/�\������)�*��i#�ȝ ��ac�*U�T���'9��C3�M;+���,�9K���O�QI�ʈ	CS�N9I��tK���5f���sԞ�N�测�j��Uך�"�E�2f���� ����A�A�)y���d��DyRF�	��л�g�b.�hք�7�I0�"O���'a�2Uc`�9B�@]��Q��X+z.�"~�3�<Q	�� X��0�4 ����5�l��@Ü�/A2���3/��ϓ6���
�'�.�� $LF���!�Ȣ�E��IF��'&�Be��T�zƏ�0��X��'�����3�@XC�$ߖ(=в���GX���ZE	�r`� q�R+|w:�u��k�<�$Iŵ&Ԙhw�G�o�VP�'��'L�\H����9O�����
7f�XՇ�)
�<b&"O�)�)�̵XT�&'�pE:�5O��a<�O<y`5��)����!i�N���'�Y�Z�Щ����oD`i��gi�����)D�� �I� �hw��)eaU:n��P���	�k�6�G�#�5O�R0у���t�Ĉ�y���OkB�W�ـ��I��ȉ�q}������s���W��F�	IE
;R*�w�<D���P+G"5��,a���U�5S�@}�,J��Sx�L��cѯf�ȑ�(B����Fx��F{ʟFj�g�<Q�N�Y^.�BwȌ�Ƒ1�En�<ae��&�쑗���`eܱI"h~2_� ��Tj�S���O�h_���ӻf�|QU���0?�+O�1���O��v\��]Q검�cΜ3JX��"~Γp��Srl�/�pY����r��1G|��u�-���>+��) ���*E���	����'�5�b"p�j�h��)�,*�N$K�Ϝn����$��g���$�S�I��$j�	�?��U�6)���R�c�f���/��o�ԔH�o��?iV�,�gy�e�Q$9�"]�NH0͒�-���HOΔ��S�<��e����[D��&"_��+���hK���bv�0��'�Ro�!]!	��L/�E(��u�Fx�O�F$
p�R�"[�1� ��5B�6Hg�Ӎh��z�.E6�pA�q�!��(=T)��+׼t�(!���T�c$�	�x�UzF��(P�DXRweǫ'rp��%��'G�6$ˆn��i���!	�7-������aH�)#Z�hP��Ju$����.(���I&�D��o�J�!���`�d���$�\��򃌇x�<�'
�}s�D~b/e>
�'��UoT6s4�j��2v����W�jr
|�p��.U�0[w�;z|��f�@7s6�j�!�;��pJ�G
�P.2��� ,G�����`Rũ��ē)�D���jS��@<���
>:���)��ה3��a�`��
�Y�c�˄?v]!C�	�F`�=9�哖<�,��*ƌD-ZY҇c@"�1�H5���0@0�A�+�j��Q��T���ȟ��EE\�__���ƈ�c�Hl{S�>��иY����^�R��1q��sk���-�S���y����p'�ʌ/Ѐ�5���fJ-Ո�8���Q�
�P0K���00ǃ�[�]�3�'���[�<��ӃH:~�)�O�U�0mpEM�94���SgZ�`��S�U�6��3#����'�̉��Y���A`O��T�H�Q�d�'!b!��A<ukF{ծE�<���0�B�<;B�%�"gN�1��l4Ճ��T�Ps8�0�2
.�' �.A����7�x��
A�m�dP�'x���D* ,��󁥁&M�jl22�L?@�Zp�?5*A��*b��|���]U\ ���*D���Ȃ>G�DT����/����:i�6�T�E�}����B ���~�����2����z�I"$I��(�74q)tm�{>����"&5���N�z=ĕ��D�gU���iģ:��\���
X&Zd!�%�:L�J(�C�/�����*E��S�LVn-��96�N�'�y���Y3]t�� �'Y5�u�&j�|nRlb���2Ub�u�F% �g������ŧ7La~�@q�la[�F, &&� ��,��$Uw����P�I�k��uJ���^�D�ig�Ȉ>��'_ŀP�w���t��	�O��k�х�y���$&xk0��cH\��	�'��N�Q�F?�D�ui[B�S8�P�5	��<��P�x�c��S�4�&���Uq����o�;B$&�{��^,�6�8���(rpdl3=s����҉&aj�w��7A#(�G|r�i'�dZ��z�`��a�;��O�����I��)�Ŋ�� �d���D[.����@�k��B�%,��%GK*'��
�~��a��O%B}h�y��\� �b�'����Gٟp֒l�լ^�ie���#IОXy��)�?����3X����,�9+'�}0@�+D�d��B=g��ѫ6j5_O����a��ji>�3�?i��M˅غ~jb>U�ń��$�	{��1Yt�)l�F��,حM!�_	z���3@(��L�8@֋C`�H��2D9�NU�dn��g�6�1+��/@����$
<Y@�I��20����T��x"(��@����#^q�b�V�8<"yY%�F�U�X�^Y|9�I\R��	�S�Z��B�8p;��r ��zlOt,�������
٪1V�a"7.ǲ��'P5� ��<#>de{�Iv��1������U�ݿ}Si+�
� ^ӊ�2Al��X����w�P6C����Hh����Ė�	��x��ѷMgوf��<4�!�D P�>��t��9.X��$Ȑ>��Ŏ�)I�����%�1I��[�g7f� a��q]����S�8&e��	�e�r�����HښՈ�O�6-5p��0�x�TU�D�a��l�ē�F�aQJ���1��mMxBq�?�2#�(O7X� ��0��jP�� �cV" `��J�5Y"O��� Ŋ�G�QO�=	�4Sr"O
�;�dʁ=�j�m�Q=O�=ʖ"O� 28�� ��k�L���Eٵ:S�!�b"OTxJ�Ğ.^ZA��	�DI"O�q��ɔ B����=-��i��"O&�t��Xl�pHpO��,c��3"O��F��e�jm�R�.?�<�ۆ"Ott`Bȝ@{�YR��@�8j�"O.h�g/��G���cP�_+R�{"O���1�K.>������$�^�"O��
��N�%(����A�2�J`C�"O(-��Eɇ]��K�e7��͑s"ON1��i���h�C�!]�D�c�"O1�!�4�8�#�H���0%"OD�R���/��3��d���`"O轘F���a�Q��KʬSy����������	Ũ��f)Y4]�J�$�Ȫ$wB��D�<�q�ܟg�~$�@��'s��p ED�<9�$1 I�|#G��4q��(ġE�'�?a���I#m�4���)�Ƽx�#?D��c�@�'~m��AÆ�?[=�r�h�xF{�����Z<�}�b��x�|X�8!!���Xǎ�`�+4H���3�F�75�	tx��ˡ����^0{���v�Դ�A�%�O��VN�����~,b)br��D�DL�����N0����iY�_Z��G|���%Q����'�OU���D�է-�C�	�R��W�j JbDŮ_m
-��"Oj���Ē!v��#�\-=���j�"O��Gd����၊�swΑذ"O�!��LHX���I�H�n�s�"O�	��")�(Q6�U�;�V�1�"O�d�ʧo�q�5�ҜN�*���"O�VӷN�-z�H'��+��[W�<T�<"u9�o�]���ca��d�<٣,X,�� �/G;���À�I�<��Ǒ�9`�@+��̈Up��7��D�<��D�L�ت������4��9��xbƆ\ⴠ��Ǳ/n�ZǬ���<���ػ8!�!��AzX8G"f!�$�[i X�EН?��xgf]2�'�#=�}:���f�D����i!�\�Ԩ�A�<�f'Z���%j��M�4�^l���p��/�y��� KZ�(����=F6�K�����xRID�Q�`9�b	�`�ʌ;4�JB�I)#�*���l��	ڕ$�(C3V��D�C�$L��s֪�8Eܵ�����( ��ȓj�2�
�$�3[3�1�흳�@�<	����F�fQ��IǠ�>�P��`j��!�D�h��<@� 2+�l����!򤂅$ �I��#M�qbyRv���d�!��[F2"�!��]2F\:|�2!Mz�!�IѾa��lJ�$]DT���E�!��T.$s��H��LL����ճP�!�Ć�^=�7/�/gJ���Ȟ�3BC�ɻn�T	�H�^$x�_:%ȚC䉑s|�+��&{֝	��6��C�ɃV�AZB�á(��sf�֤FdC�	�Sq��� f H�iT �C�	&�X��'۪m�8@#��'j��B�	;[��AuLM�2F�
��[�3��C�I% ���x��Ȏ��;���-B�	�k
���G#ll$�P��.k�C�	�'���a�腑&z�,�q�>R�B�	�jt���3-s��7���C�I�$6�m����$p�y&HКD��B�)� ��!��]:*��$jM/o�!��"O��Q�I�nm><��hY~����"O�t�w�O�h"��P���1�R���*O2�q�)��4���S"/��O4ܕ�
�'�9pb�?��L2b��2m��
�'_h��`�""ą"�Y7��d
�'{�6�-|�z�9��y�8��	�'�lMr��S�$!�"hH�ra�<��'�PC�� 6ji��&�oV}��'xt���0U-��{��E�aڑ��'��]$��(�Juzw�.e0&(
	�'��|�l��y�% %�ԙ^�Y	�'�䍈r�n|,1�&\���	�'l� [�L  ��:W���s	�'>��H���,N��M�S�H�M �	�'ilX�C5qエ� +�E��M�'[ ��C�֞|��i�G��r��'�t�P��5u9����Cաz2)�'ִ1B��B�bqC
-rt~E;�'����@(k�B-����j��!�'������,i�v����;t���s�'�ʵ��B̄k:~aZ�D-1h�
�'h�i�ga�6��L�Uh�C2�[�' �}����;��%Ʉ�kVHً�'p��+Pn�Z�'�}6�4A�'
<m�d*h�|�����8�I�'�����/uW�}��T�GLY`�'DE(BǏ}���!c���}��'�F��dc�^}F�c"�\?J�<��'���D�l�F8�Q��<V�ܐ9�'̘((ӢB�,-����s���'��V+P�f���޻o�DS�'�x����Q��5����cT�p��'I�]2��F�A�p�`f�*P;T�Q�'B*�y@�
;cB� as�ʧS��@��'Z��#+m�US��Y�;a6�a�'��q�si�F�� �Ǖ7�p�;�'�f��3X��	��j�-J�)	�'/�-�2i_�&6��qF86(d��'HԈ�ث;f�:A톨x�ڵk�'R$�b��_�v���Փy� 8	�';h� Fj��ʼs N�g]��a	�'w,�����:~��r�e 7<ҹA�'� I��U�wo�(�'
�(z֑��'T��PZ�4���GS��2r��y���#b�xBR�4`��I�C�<�yb��z�
\�c`�}���L��y�D݀c %��ƃt�ZE"u)���y��+�b��&���;4 ��O�"�y�����X��T�?�D(�����y�W�J��k"��)5���QiL-�yថ_�d����${�2�2���/�y�3Hif&���B����W��y�Bט~���wI�� ��Q� ��yBI�@Q��Q�B?4�Y`�&���y�N��BÊhX�O�z{P��Ն�yR��L�J9�T�a8DbTJN#�y�&@V��b���� ��ĉ��W"�y"AG�?����A͌)Uk>1�O@��yR��M��Yf���y��r!̣�yB�Ǐ<��L��le�5��j
�y�KؤAx�Xل��+���M	��y��J�J�fl��/ߙq��t+4B��y2�#^��Dhw��'p��b�[��y
� ��ygn���@�kw�(� p"O�ؑ�ULJ�Pj���5#e��"O^�Ip(Q'T�)�(�1//��3F"OFI���<,��R���U2�"O�d0©�n�\���π�\lM�"O�@���֗c�@ͻV��іp��"O������/�������77�]�W"OtҀ��֊H��lZ�;-
a0"OH�E��)	PpW�	(9�h� �"O��u��([��%�!*
hx��"O����͑[ɜ\�d)�(���!"O�� �5��3��A�_ON��B"O��+�*�w��a1�55�4 "O�i��jP�d'ZqZHU&�t08f"O�QLٜcl� sg�ǬE\.���"O藆o���A�1���$��y"��*r{��pCc�5-ͶxZ�m��y��˝X�XK�h�e���܆�y�"��$!c`�fz&����y�� U�ZgF�[C~���%R��y2M?mhu��lF:Q@�\!�lA�yb�>5긨���&BN5�c/���y�%}��kV�;��$hj�yZ�t��� :{�Y��i�:"���	�',��tME-ˠ����@��'���t�O�]�ؘ*���.2���'�4x���0MJ��s!D='Њ���'�Լj%�ͧ%N�H����njl���'��ma�Α�5�6���G��!c�'V��跡�//2����m�	���I
�'X����ҳme8�*��R��@
�'��1l�<⾝C��^�|�|HA�'LT8��)�/���A5�G�}8P���' ]�T�J����ib.�1lK��Z�'�t�aE�?�
�BQON�kα��'1"Qy��(v8��P�C$f*���'���F�E-%�u�^�g�D �
�'��p�v [&5}���Ƅ;Ya�%#
�'u��s�h1qr�r����Ri�H)
�'	���J-5@�H��ϙ��Ջ�'g����@O��PQ5�?'�}@�'W^�Y��']f ɀ��&
�� �'�EDd�Pd
�P���'e0��F=$X�Q�0̶S�>�s�'��9��ڽJ��� @ةU�}�	�')΀�Ti�5v���`ʵMY`U	�'�	Eb[%J��)ǥZ�9��@��'�����ǚ�R14,[�f���2���'厭����3v��T�UI���B�'ަ@��W�n�����nRJvP��'�8@�a����"�?S�X��'7J� %��<^� �V ��B���'�v��',9�� u�C�H���'��a��?'��Z�?_�p�'���W�+X�Cd_+0g`�
�'Vr�J3΂�,,m��
�,lDHP�'?.z��  ,��CmT7%���)�'�d����P�6��2�ցJ�2���'�l#&�
W8m��EW�]XT���'��MR���`Ԧ����a�h�	�'�X��Cb��8 h��\#��`	�'ϸz㈔%�P�p :@@�l��'nT�-��e�A�ǊZs�#�'E�a��4UeP�pB��s�40��� �`��攽V��	!�X�Wp0|ʗ"OX�a���oNxh����έe"Oܤ�Wiҡ6�I����H��5"O��e��Y� )��K��"(fRp"O��X� m:��H3j�:/&��"OZ���b�M�Zm����A��A4"O�-��+�2�k�d��B�
X!P"Ohp��ǉ[j�`e#(�έ�"O�-P5꟬%cĝx��.w|}Y"O�\JѩX�� �� �9E&1��"O��yP�ފR<i�֦	%�8�'"Oy��X�
b�)u�ҟ)P�:G"O��(��lz�����C��"O���p�̺I�2u8��ī18��	"O��{���~Yv���	D2�h�"O*��c�~vl�P�K:��QU"Oj�I׮�2]��%�G�R�/����"OX���F�`��BF��`,6�c"O4�0%g̏Ǫ�𦌗�w.�e�"O�{U��
gl��H�ם����"O��臃s�ָ0
��B"H�C"O��3�I�y��I�U/��u2d"Od훶�
X�J�'a�+iK8�Z�"O�m�s�i�옹$/Km,�"O"հVN�~��2ɝ�|�dEʓ"O�ps��H5<�ڹ3��$ �b�$"O��r��L�Y��<��:W���"O
i2qM� Z����%�� ��u�"O�a��+LN��y�o_�<rڄ��"O<%���>2�
p4�T-t�ȸ{�"O��j��GE����� o����"O�鸆n~L�!8T�;|]` P�"O�=)^�Wi� ��ܕQ���A�"O�H���5�i�ǩTa����B"O��i�� (oh�#G(�\��%��"O��j���;+j�s&f�� �� Ce"Oh�R��T
�i⅌
̄��"O>���$�n����4��a�����"Ox�srȝ�f�m�GB�̼�"OBQ@�A�4"�0��N�
,��"OF��h��Δ��;���"O�8��ٍ��ث�$W�G05��"O�nAW���?'Y�Q�"O|�f50�47E"���3�=D�d)s�ČVf�YX���a^��P39D�����+Xh��)f��$*�!���7D�؛Ge�3��|{B%�h���&k2D�dEDݖ=~l�3&�! h�*�,3D���B��Ln��X�S�=�R<��3D��:�H��J� N�RM��q�/0D��ɶB['q�~=G/��7TdbQ.4D�T{h�h�\��Ɖ�`0(�#p*3D�`� ��f���&I(�2l���3D��覅΋q�+��'"�T	J���$�y�o��L+<�����JX�ǡ���y�JP�@<]{���!6Tx�@�y��Ը�Y��p�A��y�r[���_�,Yv�U�:C䉑Q_<0x�H�#�����DR�B䉜
�ʘ���ВA��0�'�*�B�� px���\�z�㤫���B��F��Y�G]rR�r����6l�B䉬{Rdx�gd�Y�&pJT)Z���B�	6cJe���7
�Ԋ"V�W8�B�)� ���K�D0������ ʐ�Y�"O2I�/�d_.��$Y�u�J��"O� ���W)T{GE��Ē�[E"Ox�EMقi���u+�_�lQ��"O��S�B��N}Ť�XN,�"O LE����X�K �L�_|x�i"O�S��N.Ph���@�g9��h"On���c����S�@/ ��$"O�L� ��Y�= �.�G2���"O��sD��KW*�FMX8g5jM�"O
���k�6�&��WB2F�p�%"Oxa'BB�
�[��G/&v�T��"O4��4��"`�q�MQ�is4���"O���mߕi�MA��:�Y��"O8�"��QJ,<Zv�	 ?qp�I�"O0�������7mª�z�Q�"ON8���+E#�`ڷ
:HWf	�t"O����A�[�y�Q��[�]ʱ"Otܛ�� %�py�j�G��At"Oİ��O��^�+A*��-��qBS"O� �u�.>���*��3X�@`�S"O���PU�E��L�E����Na��"O��1ǅM�Mx��ف���.�0D�"O�q���?;����+C! ��1Ot��S
Z�n�,�ir��9j�M���:o�ҵP1@E-�@f%�;�����
�V6M��� �cG�_>U�d�� \N$����Aj���*�f�>y2)�XTÅQ�Şv���)��D�	�i&2դOr98�)�S10�t�����rĆ�'�R�	$����?E��l�3��Y��&�i�@�'#!��9K0m?�)��R t0f�Ĺ`	��"���r� ���0|:�ܫ;�)��nJ+v��0 `ܓ]o��J~�W�_�]�=����$Wby8�nHS���+I����?q�t��Sܬ�AD�X}��p+����vE�p�S�O}�H��aQ����Lĭi����㟢� Zò��W�H8�]HW�Q���'D��	#c����~*���v%(x�t�A+3s2L���b�\yiG��g?��AB�|ɖ���P/3�mIT��'e�FP�P)ڐ~<
��'�O<-{%��JЄ��	�'4����ц]�lw W����4 �RE�8!�*5�0⧴?�%Q6>��
f(�&d�lu5�Q�ZSa�� �-`��hJ���yʟ�)�kF�<�#��0>������i���i�]��w�l���çoUF���
:�@I�C(�J��ORԑj
8hDqE�6�R����)VTV��� ����'jڴ�re��a4�}�-�>E��e��"�� y�@չ%�J�1�FV5[��!�OG
V�S­�chfQ�	�'9E�<2D�O "�x��*�4��SD��!Bv��R7����Qj˺���	X�k�R�gE-~�
!jC����JxT ���*����s��s��bVZeiU�C� q�1A}�"UQP�
+,�Hp�O�"��+ ��p�?F ���q�<I�Lן^�8,�f�;4�z\2��l�<�!6Y�<Y�#��"C��#�i�<��+E?m��7䌌�D�)4CQf�<q6��Т8XD(��Y�,q�JM�<		 x �9c/�6�H�M�F�<Y"�V([L���`	��zX��H�<��D�p�l9��@�@k�A`A�<�ƍ>K)� �0�(I[&,�@�<A���U->���gZ�B��A��|�<93E)Y�Ƒ!��A*e���Ip�<9�f�7��s��_m�}�%IFW�<Q`Ĕ�./,����ͬT߆̓�#�T�<��C?%D�gL'�:�#��T�<�d��"�H ��EU+r������W�<Q��T>plD�bhͩ!,�1[�j�L�<9�ǉ(m~�)��(O�Z�+@�s�<�Ǜ�cRdt�&X���
Uf�<� �-� � ~�.ك�M�8mO�8�f"Ox�2'Y�e���&gZ�RRD�  "O��W�κ$@�ld�NYe��2"O.��#J7j�$��Ӫ�)~Q@`G"O,��#�Sc*���ț�c��5Rd"ObI&I�ƨ�r�̇f㔡��"OH�Jů֯
a��i͂j��A�e"OI3v?�6����,n���"O��p�@�.V�@�@��#�rmIt"O�(I���]W�����[Eĩh�"O�����s� @
��/A�Di�"Od��dLN&0��<Aq��89�`
3"O"�Y&�-��q�mթ)���E"OX�*��t?��z]J�%X���y��L�{�aJgF�(��;�	��y2�_7TL���Zi$lK�+�)�yL �rPc�I 9����W��y���FVܥ��/J'7ehh��� �yrʒ�.~����H��,ޮ�Z�	P��y��.�Lis�l������UKN��y�B��L9���J�.zD��,��yb�*}�F�A�㍠O����$B�y���wzV��UeM�K�`��L�yrgT���hÑ��;w\j�I�'Y#�y�l���x�D�8`
�PcG��0�y�$�2)ߌ�&���AI\���.�ybk0<�"�֣A�Kڐ
�)�yb# $���/ /?��*�&�,�yr/�y��ń��I�2|P���y""�~6��:F�R�;xX`XѮǟ�y�
J�&����J��Fa�� ����y�ȁ5�����ʕ-7`�͐�y�

S��R�(��������y�Bu@��ꄫ\������� �y�x��<_�#�l�X�MI,�y�gS�B�Ny��R��<d�A��/�y�aM6}|�A�Q�%
D����J��y�$N1oz
�{��	�������4�y"/�%U*��+&�]�]Q�
9�y����6xh���
�T���T��y�!ӸN.!1�a�¢}2�G ��yB`A�/Et��%/�VXɧ�V��ybdϹCB!�5A�39ި�iB/�4�yb�ri��A�$ϾE��X!ro��yB�F r�t�a���G���rQ
���y��V��	s��U�Ր�+N��y�Ǘ:(�)@�(S���0��ybbG�]�	�'j�,^S�} !e[;�y�G�%um��c�W����y�Â00ZT�1k P�����
�y��$no�m�C�٫�zl�7lM��y�"=����P�_�LY�*M �y��\�v���dL�-��⠊���yR��?'��@ �@
������yr��|��`C�Oδ3�Je��nǚ�y�I�hx�I���	���+P�y�	E�.E��+�P��~!�qI��y�ID�@6Ĺ��/��~�H�����;�yr��	t���V��|"�ࢊڅ�yR%�=]2��˥O%b�xU�[��y2�Ĩ0����(Q
}o�tR��٢�y����|}��FPvڄ��@8�y�Ή�\V��g��08"��s�ѩ�y"�^�1��Pe�I�ȹC���y
� ��ڑ�L��x��A���Jij�� "O �"tb���pF�]�%P��"O@<�7�<�\�aY9,�d��"O� +Ӡ�[�hZ��εg09�"O�4��hK�(�le��ʖ:&]9T"O�%�1�ѹ5l^%
G�2+C.�%�>�� ������5X�b�܀���\���G��$J�1pJ5����KO�u��_�&0Z�s����<��ȓn$��qf�e��F�W^|Ąȓ��H���J��|#�cÖ>�x�ȓB&������5b��ܸ ���V��YB�UH�-22,�d�F�3��͆�I4U��`O�e+�i����aQ��T ��g���v!�q�?�ȅ�we:����!yjPQㄫ_b0��Kh�B'H�3��L�����\1��Ge���V�EI�$u�� �%y����x�H�p�@�3�|�2�	I�l��ЄȓEe�A��ۜqA2�Q��0a�l��>��Ţ�%K$ �8ջ�+DG#(Q��Sn�|3Tc�Vɀ��jB:4b@H�ȓg�	3B�E&.��r	,.P�ȓLk�ܘ�E��1Z��C��Ɂ[B�ȓ���qQ�z�)��<>+>��ȓ�0�R�L\ &��]@􂂼&���64:���;)WX� +2-l��ȓXR���۫�aP#F�^*C�V��E��d�2Z������@�4C��D��ub%��	�Ɔ�
'�C�i�W��Q��)pbaζqBRI�e�7D��!�jQ'��
�I�af��j2B2D��q��A ��;�oJ�Z���P 6D�((c�(a����ۤA�b�P��1D�<�q�Z��`��Z�<j
h�'1D�,qt+��w�T�ӑ	)M��}��+D�lҀi�9���Q�W(XNz���)D��2��9i�I(d�զga"��s�,D��Z�g�*l�%�!@H���`S�/D������|%��:��ʫ(W��y��2D����4 �\M�a.	�[L�Ai�o1D���E.C�J�Z|�q�E� �v}���3D��iv�U0�+�0~�B��2D�\�D/��:�@!2s���S�w!U"O�A��\���`eS�=�,% A"OTP��"���bDA )����"O�}{V�۵%ِ�h��]�d�>i@A"O"4C3CP�/�T���@�k�T�Ȥ"O�Jb�� @�d��E]��H�"OLU*��`z 1⤎���L1�"O�E3�Q�THbP����r}��ۃ"O�=Jr�=%x�-�>}n��:4"O����o��Pm������50l��є"O��a�lѽ�Z���d�-r|���"OX2	ũv�V�
� �e^�)�"OrD�rjл; � @��VM��k�"O`��b��52m�aD�-A�8B�"O���C�L�KP�aa	B$���"O�P	��0#c��2��"O���F�S�8рC�[�Gz�%�"O"�1G�:2����!5^z��c"O-0���$
����0F��%"O E�H5/��m���M�x�"O��ìT�\_�}c� ެ=haI"O� ���B�W�t���-=X!�l8""Oxei��	��L8+��_W-b�2"OfUaѮ�v����3nی6�<��"O�<h��"Y��\[�j��g�dT��"O�AC�+;�M:CkM��(�y "O^�K�E�5[ŸxC�
%S�Yy5"O�<��}RY��oʫd2���"O������~�,$�r$	#$�R�:w"O�Q�KL�g�p3��Y��Dh��"O(t�U�
K�D��`Ԛ)��k�"O�t�g��l��I 5"B�8b""OJL	"�E?�8�Z=1:����"O,܋v	�oʺ}��N�\8�u��"O��+��>wJ�&Κ"_2m��"O�dQ0�J$��,��m�'�Ѝq "O�l��lőO8�C�.T�=t���'"Oe�� �+��(vC�aʵi"O&-��%�L�h� �M�^bD P"OP���e�  r��KR�K��H�G"O� 6�L�95 ��$*��v�� �"O*���.��쐹�5mW8հ�"O4�)2Ǖ�L>�sd��gS���"O ��7͊1��� #k3v�s0"O0�bfj^?4�896�ÿFҰ�U"O�HQD��N5~h�@␩,�f���"Ov��*E�Q~^a�����2R"O����,R���e�Av��8�"O��p�m��Du�`��&=N�jG"O4]�n�
8M�'$� [A��� "O&�!�Huiq%�7~* ��@"O�s�ŗ�]�^�j� �*����"Ob�����8P4Y�uȚq�@�n"O�p���p쵩�';�P#�"OVDcr�͏X��Y2��/^�NaR�"O�a3�n^�F��� $7���"O��s5\C����dC�<C*� "O.`ADGڐZ�,Ÿ��Q!n����"O�˵�˕��Q�L ����"O���S$�t�D��V�
�{^
Yɱ"O������JѰ�G�=3�P}��"O<��`�U���m��:��6"O�8�B��Ln�u����B�����"O8i���D>_��=�2'W�K�p���"Ol�-6n���P��މZ�"O ����̬"�`!��M�[�j](C"Ot����i8acU�����4"O�鲗�
'5Ь}CR�F-pޡ��"O>��E��v�H/юQ4ER�"O*y���[ݎ\kT$P{N�`h�"O�(��ևxwX;��I_Π�"O��vH��+������  G�d��"O�����ʽH�h��E'�6E��!�#"Oҵ�θ=�X��E��*�K5"O��	   ��%*�$XP���ɳ:t�S�=�?"$j�.C�����L��)�#��<A��{�����?��?�����dU`�|<z6D]�dL��i�e��˓���lI��O���3G��R���ץ��4�8���}�������?��?��'��4����1/�0oX;����d�'LΠ��!Dx����'(�8k�#:Y��!���\�if�0g�'2�'���I*w��i>����v� IAe��l6��E�]?d`A���/��'�?	���yr.
�F̾�s�N4~��e8�[�?Q���&xk/O����O���?�I-�
� ���ax���dE�4ʓT�`�8$�Lj~��'�[�l�I26y��l_�.Y��NT�xjőp��sy��'(�'��O"�$��&jބk�˄VhXe�᫄���U*S�9@����	ky��'I�1��?�����G�J�1�c�ITA���'5"�'�����O��˖c��lLj�I&��"A�5x�/�6��E�G��<����?�.O��$VE�˧�?Y�%7���f�P$E�h�j��O�?y���'抂Fu2,J��aP+P0+$��)H��������O���<��"}��,����O��)�B���ǂ�<=  �r5ș�fP�<�	�B�:��`:�?u�0':}ux�;'�X��:1��<��F�����?����?�����$W�0z��Ӑ��6��j�������?qF��5@w�1�<�}��	���")��s`@���ϟ� h��c����-O���O,�假F+��s��~ф��p��O��ȓe��O81O>�����z�KP+B#>�@XE��9pQ���	��Iş��F�[Jy�O"�'9�DZ�?��X�a�V�C���Z8�y����O>2�'_�DZ�.~�� D�6!�k�e�^p��'�F�jRP����ߟ��IE�AG���#a�>Da4t����	v8��'����!" �����Op���<y�#l�Q�e�!d�Z� ��
�"P�aN�����OF���OV�T�I*}%�aʐ�%Wa��3�x"��� ,�s�>��?Q����d�Ox;�of>���eF�KHd���DS�|�u��Ot���O��d"��џ���Q� �@�0��Ze�L�i��7u9���Hy��'�2T�P����4u�O)�e@�B�Lq��O.ΐ�`r�6n��'^�O��D�.a8b��6�>�7h�*@D�H�'Y3j���s���ݟ���Qy��'4Й#�Z>�������.#�D��LL�5L�˓�T:>M2%�?A��Y��(�#Fg�S�DoE16���I�n HNb��c�\y��'���'>��'j��Oh�I1#�"�3 `B�2�jg�D�hz��'D�E�~\��y��,X�"�ƈN�&L�` ���?y��@;�?��?����Z.O��O�|A�8�Z���dޣI������O�l��MJ"Q�1O>a�I$ov�C,O#2H"��-NfT����	��a��Ay�O�"�'�[<�a�ݲ%����qHR��$,ڎy�OYV�O���'��;'^q6��9�v���LكaM�'�ZY���ɟ��I`�|��	�扭
<(m�򈛈O�䡔'���3D&���d�O^�Ħ<I��i��9�F����P��%N�Um�9�FAW����OV�d�O����I�BMb��s߫%x\z�(޿F]d�ԕD���?������O&U��h>�k�%�YDkB��t gȒ��?����?����'}���(H2�!ע)��l�f�8;|
h[��ù4�	柨�	jy��'�p��W>��	#L�5 �D���\\x��9@�6��	۟�?i��J���@��N��]�,j��"�,A�	���D���?)/Ot�$ۅvV��'�?�����c�0}
����~N�ӵCJ-m��L�IY���g�2�?� vT�1H��e���X�$��8�vqz"�'��ɲ�����4����O����ny�(�)�d" GOws�u8���?����?�'�͍�?i���?����*��y��~C�h[c��b7�h�s*��?!A�]���'}r�'��4�O���'.R��j��]�@�8K1���ӥY�C�n#�2�|�O��O���
mffٸ����Y��"g��1 Nf7m�O����O$4��������Oj�d�OL�dϗ%�t��1D��
�K1�V%j@F�D�OD�D_k�%��b4���|��Ov�
g$?T�T!3����)yY�a��O���զQ��Al����	ڟ<��;���p�`q���1,i�ɜ.x��H s"�<��$��<���?����?�O~Z�L	<��rJ�=b;�ls@�Α�έ T�iS"�'��'�����d�O��C1�ϗ.<"���p�A"��+���O|�d�OL���O�'3Ϯ�W�i}��;֌�C��ƭ�~����';��'���'�B\����?DR(�S�@  XQCaV)v��a�7i�#����՟p������^��רrp�7��O���K�,<�A�`0"q3�B q���O���O�˓�?����|B�O��2'I%�F!�'P4�(�R��'B��'R�'`N��Ii�8���O�����LJc��V�A���
ư)R��O�Į<�;��Tϧ���|B�ε�B�*��ʩR���H_��?Q��?! �S��V�'"��'`���ODBm�0O�tx�� ]��c�"7���ˡ-Lʟ��'P"�+�O)��;q|�2Dƪ���Rw��E����q;�nZ�T�I֟���?��	��L�I�oA�!��.%6�΍z���\O ����JNT�'�i>��|r��1z|���EF���x8��8J��j��i��'�	Z5���'�b�'�R�'��S��/N�L
�'�5tn8R�0�'���O��O����O���[�S�E���,F���r#��O������n�������I����c��2�֖T�4��Q�ЫQOF=����<���<9��?y��?I���IZg�iA?>�B@��)Z��ل�Ц%���P�I�� �����?��i�L�P������`
$h��*�L���?)���?����?9��?i7�D�^ۛ�	7�RPAC�K�n�i�G�:��'���'h��'��ßBFo>��EkF->�����F?b��[C�^My��'�"�'4B�'�F(�Q�x�����OxŨ�H�1�S�⅙�l�ON�$�O��ġ<1�tb؝�'���-\�PkV`O�h�-��@U;���'H��'
���R׶iB�'��Opma�2K�N��C'�3�,��'��P�L��!��Sؕ��nݫ�,3�I�5��2�Ȉ$9���'��D�tH�6-�O$�$�O��	�����
Ӗ���H�>ap��G1*���?9�nɆ�?���4�z�0�42�G�b�͒m�h��L�		�b2�4�?��?��'>��	Ry҃	���5��Id�p��l� t�R��#�y"�'��	b�'�?�mB�af���F��2�!����8ݛ�'���'�b��O�R�'d"�'��U"kU��p���JF��*�a�;���'���M�+"����O?�'T�] t�S�R�2���Y�.���'�bӶt"�6��O����ON�DF[�$:On�9��GK�X�@#��{���&�'�IJ�����y��'�2�O�2�'��#HLr�Z�֑ ��ǦY������M3���?A��?9�V?��'�ҋٖ��@hK&���mv��ј'���'�2�'�"[>�Ra���M��6gA��ℨ0)�U�'�;�?���?��?����$�O��w?��Q�ऀ��Uh���*�5`���O��O ��O^˓LPR�C��4`ކk��'�Ѐ�@@E�K�>���'#�'���'Z�����'��	�P�&�Q����_^,�p�V4El���O`�ĥ<9��}}�O�2�O�X`Q��=s��qB�[%��}�g�|R�'�R��"�|r8�����H)He~`ʗ�ϓ �,���'��	�+�ةش��i�O��ɑEyBb�� �P0�	��=U�_1�?���?aE��,����Oh|UK=lR�d�±Kn8��l����c�i&b�']��O�*O�����m�d8�qbܒm�<��5s,n�Ě�vb��#��̟P�rBW� �Nqx�#Y�
�4�SCG��M����?Y��Y>��H`�x��'��1O�y�á��kWM�%2K^a��'�'�m!Ş��'���'b��Ҕ	���;��&���Ӆ�'6�-"�>Ob���O�Oǩ�7tH���͞% Ш� .����D��C��<Q���?����dOܪ)RG�4*�*��
|s� �4�P�ȟ�Io��ȟ�I�G$�}�2�_.M�M��k�.��}�C`�g�����	���'XHwk���@)^%U�d��[�4E8fU������8&���������z��9�'N�s���'C��( �څ#Cxy��'4�'��	TV���J|�HX�A�����.�7�l�$���?����?��Ê��=��@ۓ�pїOGp�%*��̟���ڟ��'�D��v�"�I�O,��Zzn��0E�'Z�d�h���a���Of���Oh=ڲ��O�O�I��(]yaΗ�O�ZA䛃[�\����D-�M�.���|�'�Bh�A�������?)�v� ��?��6'����Sܧ~��d��m�ԀAcؒi?��	&V%����4�?Q���?���lۉ'��#OH�n��!(O%H���Q�)�����T��G���'�� ���b�>�Y���+00}R�al�&���O�����}ʁ%�<�I����j�f�rmšbpd����38����m�:]WH�'?����x�'^F�[�ˌ,A#���&� )<`��	��x�d�����|���i��	�wR���mny���?i�-���?��?����?i����dP�=h2�2L�9������*T�m�p&^_��ٟ�F{��'���6).b�@�[����#K��O�O�R_�l�I� �	�����7$�	���e���p�,7�����o0�����˟���ٟ�'����ٟ���/��d�m�m���h
�.~��<��?���?���ex�=�*���D��1��(�470jI���+�����Or�O����O�ݳ�'��!2��8�EG�� �#��8�T�D�Or��O<�$ ��ʧ�?����b㊚�s3<m3���A��)���L����?��YJ0�Gx�3����_m���+�ϫ("pa��'��I)X�T �ش��	�O��	LDy2�өz�2�RU�;=� x9Sb��?-�M[�T��E0+O�)�O���>�5�!f�H`�`>f?��A���h"po��M���?���� �x�O���XcѮ���$��p\�8��'�(�r_������3����&KSp`�*�c�@���K�i��qU�E3$����i�8�<�V�	�\j\���ꟴ�	��C��z����V V�EQ�����I��rnc�\��˟��IΟH�'�-;���!_�>�C���=�2i;���?�ݴ�?�"�'h��'�"�|b��I�#l�K&��#6��eM
Lc5��Q$��9h]�T�wFŉ/�v鸂*�wQ<�5��R<�.+!���/�WG> �.o	!��9v	�7v�����\��+���5G� �'���8�k��<0&�Ӆ=j�1�q�H<�pkC�I�]C�*�.��M��)?[�@�zueݥ�
�{���4I�JA�A�Ik��jL2^���3�*1O�:���2����th& ���pU�H�p��Oʽn�!�Iǟ|�I���Xw���'?�)��Im�,��
�<~<�+�M(�;G D9}��H�U�a؞�Q�dӌ��x�
���!��&.\�q)�
��W�j(�۴v<�c�b'�-F6���]�k�H�Y� K̽(bbSǟ��IP�'G�O4�Rg#
z(���p�D�C�%"OT��ܮ<�&�����$O�vTPT��MئQ�	Ly"!b�6��O.6��X�t��a�&E�h��
�d�`��I�z�.G�����|�r�Ȱ'��t��ʌR� hp�#��B�<1�2��9
���"��(ZB��X'��f0QdiQ�y9g-BYQ�>�����P� ��CS�=`[b�@���f�/
n��D�|�ĎT0�2�P�cs8r%�l!�ě�%A4� ����Zdt�Wդm���$� L�P#�"��<�5�H�*�
A���4����P�A��O�"T>������5楔8L�	�%��`��-A��?��Q����~�R��#�?+*�$�8ȸ�sb�h�4Y����$�`��¸�YH��Ka�pD�T�G$5�ڱb�D?V��l�b���ē}�t�Iş0D�Գi��(�|x�䕝��q%�w�<���>k�$,�D��1��P{SNt8��h��d��{�xUy�-Ѧ3N�8s`k]V�B��4�?	��?���!6��"���?q��?�]�7Ҫ��O<�0\2�g�9D	@�ޚ,�2ĳr�'*Hʳ�L���ē%�
�b_h�ԋ�CI�C��A[�h�(vO*1�&f�O4h�O�o�g�	z"���R��!p��Q-V!lQ0����D��e�O]��zԥAZf�bcN-t^}�Q 6D��å��n6"I�g�ixT����?}� '��|�������ac��B�<k����a��6<jȸ�^'v|D��	�X��ȟ�JYw�b�'��	�?���P��B	e�Su��9
���S/��L8�\q��%UDz<�bF3�Ge����"Z/�H��E,�d�:��A^�%eÁ�;�^H�Q�Z�a�z0��%S�aD����¥ơj2�1�JиK�2�q��O\b�d�[��@��[�<��uf���8�I0�OXO\a	�ių�����/q���v�$H���&�@�����Mc��M�/�qLf�b����ѫ�.��<���'pP�`�'�B>��B�im��i67;5����Y����kX	�P�V�H���<)%�۩�5��ڊqMv����Ilt��ʃ�"G�\ʲ%הA�\����	?U|��V��s1�����OVb��Bc�,��a�'^���,mW�@3B�R+)�Ƀ�'��m���
��(;"R��1Y�iϢ?;�'^9jIo�x���O�ʧ��ɹٴN��]�"J><ဥ�t�R��$���'/�x���i��>x�]�1�G��'���Y����c�$�D{jp��Iڴ$��'�p��$��y��qe߯@�H"|��J)G�a�"g|P�WlY�;�:���O쓟*��ZP �%<��SAOre�� ����Op��D\20�� �8"�@E@���9��x��?ʓM8��2��H���O�P}h��p�s�����O��D٘)�d!s�O����O���w|�uK��'�!�#��Z�1��%ծTr� �f����j|�c>}�O� *�����9
^�A��T%F�&	��6l�"���@0��{��X/����5���?�^�l�r� ��3?ۄ�ᐃ��,���c�|����?�}&�p�s�̉ZLY��It�ʼJ�*D���*�1�=�!L=��8YU�(}r�'��|*H<��GQ�g}n��D��mJ�r�kHHJ��Цd^�@��'���'vl��ҟ��	�|�E�*��'��TEwV܈�A$#�x1��sP.@Q����
P�6\�č�}� Q��ZG.�`�iC.Z���i��ـ�b>�����"��Hb���0��Qx"$��Aʟ�����Az�F*��4�� "5��+]�1�_y<��(!�B80���=逾i��'����a!�>�۴< ��1w�ю*�B5i���4W.xȓ�'�R�Re��'	�X�U	b�(����F1��LSW��8lj�Y�c�05�̕ppMm�'�6a�倚$[b)%HȚko(�c�!��6{�y�LX�?�pِ2��!\{f4j�ўP�l�i��|�ў�?)��?�ݴqjU`B��W0%9�@�(=*2�GP�d��E�S��],�yGiH�;��`� �,jѨ�Gy��i>M��-�(5{|�	%��{�0��h�Fb��I@y��^=�|D���'_�X>M�׀�e��&����s^�)Q�EH��?y�!�.���
l��"P�ʧ��	Yl�q(#��ID���ҋڮ
-�'�VT�E��MF���B���8R�3$�P�2񅘆8���đx�`1�?I7�|��D͜4Q�>Ń���|���+����y¢E�*�ā'�&$މ�2j]��9��|���)V����ԈP��`�C�"/J%�r�i���'0"�)?n�z���'x"����FN�qA*3�`��)�P0	1X���;L������K��c>O�0 r�ՠr���
�@����u ��C����4cd�)C�Pb����'��R�f�8{d�'�[
Z�,i���n�X����xC�ER��%a��mI&`Z��Y��y��L�Y�Pر􇑦c��U(B'��ɜ�HO�I0�ʧ�
1Ɂ*S�=�*�=1�Ȱ�뗞~�(���埬��ȟ�Yw{��'K�)ڵmd�hW AN$ Y�F���<Z��F�R`�������¨�0�@I�'u椡�F�.�,�f
P:���Q����H��[��=� ��6���>Z(��=I��\9��5#C.Z2;��b��qȅ��"�p?�`��(pN5�����WЍ�&!P�<�!#�9U܄�H@9o*p	�!vܓj����|rLU��7m�O06mX/KDv�C���q��D2㝌hr�m�����1�������|z4A  �J�sI�܋�jЎy��ٳD��s��e�7,O�Q�$��5�^=�LڵL������z��@� MJ�R^��j�ą�>y1��*��DW����@��A�B*��.��HF�4{�!�	4����%b�3�Fd��(�ȡ�d�%[���Q�LS�%B��2��/@[�p��9���8B�tnZ�L��]�t%'zě�	��9���� ��&t���C(\�b�T��O�!�a�O�c��gy�b�l09�2
��!K��"��U,�ēl,NFx��T��Iy��PϦ�0���D�+��Nzq�	i�S�'r�\{���	`Wv�#�꟢'@pU��Ȁ�I���! ���EF��Y��	��(O�i*�MG-S:�X�N��d��%�M���?a��5�r�3�Ѝ�?���?����e!B�n���aF�W���n_RU.܈IVg?I�i?t���|&����}s�P�I��A2��;�����pd�͞���:�!\>p�2-0K^�M^���:�.�9��j�#�h&i� �z�0 �H���y�00�)�3�D��n�t#$�Z���m� ���(�!򤅟<�����
Z��=�D]��jK���S�	�Y=Ɓë��T�A�)K�^�X!L�*x�LC���?����?Iӻ�F�$�O��S�ZU��kĆC�؝2s� ;�U �Ä�V;�LQq�N�{RJاQP���h�;L�y:ċ���hJ����|qڧU�C�l�4�Ƽcў`PFf̎��C�C��� �m����D�m��d{��ס��E�(	�=(ֱ3�A%D������B@�A����!���
�b$�I��ML>y'	Δ[l���'�����**�l 7�f�Q'DM�U�p��O~����O��k>ScjK?/�Pf၍b�4ے�:Bd�a����
w�xq/Z�}]�F�	�+�\���(_�*�	��%ycB��g�1d#rl�@� �M7�!��X�1�����/	������$@���ڳ�� �C䉞v��q;ߡ;f>q�qb�3��C�0�>`y��^}���A��i�xm��CV�ɎDp�Eݴ�?������p�6���`��M%eܟ7n<�
\GZ���쟼A@^�N�����P��2�S�DU?���>�Z���ꌥZ��܋��<�}��e�t#V q�d��2f4��L1�� �H�g<6�$���%N�KS �	��xbIK��?��y��d�C�3��+���tEL*"���y��T$E
�A�ac�p+TE�D�	kX�x��$�A��IcfJй)�NŨ�d���a�	�����=e�!1�\����Iԟh���qɤAӵ,=n��tk*�t�g���:��r1�B�zŞt�CHIH�Vu�|�@hE�|���$��}��6a�0�b��I�P�R��㗶Z}�s�]�St�4BV�,��2: �Ҟw���Q����g�l������AȒO��������Ne��h� ����"q#F�hi�ȓ4b8db�_Xg�k� �̉�O0YFz�O�':9H�J�PLN�a��� �U�Y�vQ���Oh���O���P�k��?��O��i��)�X�Ⱥ� �gp�e"���,�������?[e� u�'�@q�b��.��($l̔s�� t`&l(�!�r�LI��'!dXd�Eo ��8&���^b�	0D���?i'�'ɚy[MZ,�SgG�"t����'�x�	�{zɫ�eL��Y�{�Ic� �O*53B%�Ʀ)����:���KMpp�Va��hр�P�e,�?1��p�n����?љO
��(풞Q��(��O5iJ�f%^��u��e
<[x@����$8"?�+ެ/!U��$�)_����'��M��\36�@g�%�� �'i@1�w�i�̂0o�]��'�̢����p��,غ7� 4DջM��d��=w.��H��!�)���=Ey"�i>!B7�tnia1i]_2��,�l6\U$�l�mD��M���?1*��tP3�c����&��4o���:QO�16�p��嬟����	(0�\�b�	ބk��=��Ͼ]�x$K"ٟ��'/D&��^**�Pi#�+�,g�D�'�����[8o�©q$#� �R
�6W�I�ի֐L-��K��O�Ԁ�!eKܱ�J�2��@Ζ��		��S�'Bf�$��i�2�j����2,�0��^c)�[k��a{��N�6�h��ɴ�(OVzơ2vA���p햱f�|q��"�#�Mc���?���o�f�"� :�?���?y��ߥ�F�6^���".�@W�91 #��h���V�F �P�A�f�5\�ʍ�D�2?!���;^M��igb�*W�p�s� Q�[!l)���_�OCp�F�л'f"���զn?˧u��V�k�)�!�>|o��BB�8WM�������?�O�<�����?A��MӁ$�6M�5�RCš�
�����P!��57�\����D�{4�փ����$�OD�GzB�O2[��Gk�n����a��)f�1��08�(ES'�Ԃ�?Q��?�k��N�O���~>1��+�*Bjd�!Va�
r�K5G�Z�Bb��:p�:��T8{n�J���݉^�H��eD$3��z`�4+Π�����cBH#��3c�9hP��h���e�H,��' DeۀmXr���d��ej��#g\��?1�'9��"�N ?�\j��2bUP�'��M�У���X���pl��{lz���O� �`F�������x��݀4Tr�)����n��'���?���L�2����?ٚO�����\`�8����~ܙASm]A��v�oK�cn4,O� Z��Z��1 �03d�S�&�]7*X��-U�>�" �.�jX�H�p�O�@�OĘa *������%**�f�:�"O��C�Z��PTH-k�X��
O���qŝ>)��q�拱:j��r��TWޓO��Yʦ��I˟ؕO����B�if���C�y�pAB"Ѫ%��m�gf�O��յsM���=�|�'5rP���O3)L�M������q�O<�F�n���O��J#+�Y�^y�����xO<����L>�~���;S���hU�v�t�w�<�"`�0y���O�8�M�$�Uj8�����O�*8r�&UM�!b���2<@\X�4�?q���?��Ɵ�ah��?A��?�];wt���"��[�(���d�4����GJ	�g�ޕ5�J `�D���O���eL ���I�v-��g��jƞ4���<��XZ���\n���G�\8��1K?��Kԓ�y�C��l�ɀdK�7��Id�O/X=8�&��idi�Oq��'7���rɍ0��1j1l�>1HpM��'䖡�n@�y���EB�0 ��xO��S��4�&O^���<.$��a��QH����60�%D�������	��u7�'6�>���9&m�d]�t$��\�BT�p�U�6� �#�Q�rM�6��?>,�D~�ň3�3ӀަK��X��d�ڙ1r��=@U���<�np�f|��@5z�Z�OhlY�$z먈��ʑ 2J��F�
�5I��*�O��ڥ/�D���k�-1R��-���'̉'��Se�,�td3�HG��
u	�{RLa��Oha3�¦�	�}¥�5f�2�S���{BF<�T�ۧ�?��G�E����?9�O��A�ݤM6���W�<�M%�L�k���+�XZҐaW�xX� ��Y%9�vt�  �Pϊ7MA�� `W.��?�\@]�ay�\��?ɧ�i�p7�h�� .��G,J5!t$={ѪIU�l! ��Yy��'(�O���5f@�P�x�J��G�؅�
O&(c��E��uEF�@� �2���~�W�Z���,��I퟼�Ob�y�p�i=�9!�B	d����h�U�#ԣ�OD��N�X�>�D1�|�'O�4���WX��*v�Ӭ9n��pJ<!�jY~���O�	u�C�c���1u����(�N<�#�^̟@YH>�~zdfR�I�*Py3�9Or`�pXo�<Y���C,�e�S��1X^K��"68��dZD�'��ӡ� �wx�C�
W0����=��ߟ��2F����a�ß�����h������AW,v� At��TNv� 4HV,�p�����v��	d�@����|z���)(�|��D�A� &���#݀b��x�TH���e�A�sH
%�nMP����v�;���5]52�Z�'�4��@M0�Ę ��L<!���KK0����V%\���KM��<a�C����8�L,{Uܑ���a�ēf���D�x���7RB����ʨ�A��H4	=�X���R+4A����O<�D�OV����?����)C+��U(��>Y� �$��Ǭ�]P�;��8$p���*&�e��k1/��;��	����*�3���8/�f���l߫
3YP�
^�,�Ej�	���㞨ؔg��*�Q�����#O�77y���PE��0ഢn�D���ѰH i0��*D�ȫ��<%�8����7Ry�\ȕ�'���M�M>�5�V�(��&�'Y��$��	�Z�����b���a��U'iHL���O \ɤ��OL��x>%Fd��ڷ@ ���� '  ��/���`x�'@"(p��$�%1aA���v~PP� �I�,��v���R~Ƀ�cĻ;�`]+��'C�D���ēp�^ѹƂм4�����'�7�@�ȓ.R*�QꙌu�X����L0k%�UFyb�i>�R"��g�p�ȉ�?Exmbe�oxB�&���Я���M���?Y-��q���vӮ�00˛2�d0#͊3x�	����ʟ��I��n��%Ѫ>kv=��i�~��F9\��A�,V��1g��A�	�o�"�qR�I31�"��@N")7t�X=N��ǯ�z�I�����O���r�b)�ag*:��J�L��,�v��O��򄃚��`��)�0���*'��S��xr�$�
S��(�`ܒ�ݩV��_�]�y���O��_e�,`���O����O��Di�1� �T	0=���� `Ņ18.��x���+8}�1���
d\h1���4.&?)�	 =�zHJ�
6+�a��B�Д� �C�g��I���p�����.������Q�w |K��5fJ�O��:u<��?�I�8u���x�,Ƶ~ֆ�1G� m~$!��$Ӽ�y�hڒ}G��`lӘk�����0��	�HO�>��_�����o�U��A�H	�Q7�9��0n���������Iԟ��Xwb��'��	D�P�.���EE�0Y+�� QD0iv�,<�=Q��_,pn��qֆ�J�'P�D1�M��Ē�ʧn�!'��fR�������v�&�[1��L�7��wF�y�I9�_
�@��V����,�S�dh��'�����-?�L��k��	?�r҅��e��|��x2N�b-~	�o�L8�xS��S�׸'�B6�3���#_b�l�埄���D !�%@�4-��}��_,|�Zt�	Ɵ��4Iş��I�|���֢O����&�6K�Z�a7j_�~�rY���g"�%9���5~Q.1���ɦ:�T<c�D�InI�q���e��DJ�cR7Bh���W]���rH��.X"!E�ʮxHqO��"�'�'�
�*g�Wg� ����U0�b�'6�	��@���G�T��:�'z��bK&p�
Qs��f�0	�a��*��'�Vو�Aj�z���O$�'��a�ݴm�>�č��Y�Ԑ��<���'.� R��@�j��[��`���2p��������(]�}�S�ҟNwB����K��'�04y�+\��E���+]������L��1sϜ�?�*�J�/�^![�̛f��B�"��V�7���*���K�y>.]����L����'� A!�$�M��� ��%.DDͰ��.�x�/<�`�� ��C?=�T��BO�L͢��o��$�O����q�X�.�r�'J����CEۦ9�P�8�A��#��p��-�6p hٛӎ��cV��Y��j���CU���|~©_!7�de�$��q	���r�D$)�5[��[y��X�Ƌ�!Z`���.9��67v��3�Õ)�I��ʎk��zdlX���h���)�3�dY'T~�Is�j�
 �mj���!�W,r`�`�2`��}P� ƺH��?���G�	�S[�ʆ��!V���$�`q���!�uLVU��?��?������O �{�������2pD���k�0E>��;��Ov�Ų �3L�&�Z'ń&��OJ�;��J	�<50���93�p�pY�#��eA���%
b�����˦U�3EZ�i�4'�H���C� �	��ض �v�( ���_��� "��K���l�#��4ڂ�[��'+�'�z@Kcf��A54��#�i��{bpӺ�O��q�Q�e�����2�-�J�'N�	~TL@����?1��>\:�����?ٝOT�1���	�;�ܕ'������Fp��5K��k �i
�]dtY�nۢ#q �"�A05����0<���2�,۪>%����_z��qw�Ov�m�*�~�Ի7L�)s��Y)1�<�rED���~"�'�b��	�<y��uҗ�@%UC����
5���AY����&7ұ�a�5%���I�'J�I1cwV�)۴�?9���)J�J�7mB-P�QA^ t*��;��<���ӟ��I�WE|i:��%�6�@��)t<�3�ԟ��'\�H��'�
9��鐡��y��A'���������ՍU�>(�A"�y�LA� O�D-��K�8j��V����ԍX�5�xO	Q��'�<�O��Z(�����h"uc	�O~�bR"OJ�i�,�-,����O�S1����'HN�<I��؋ms�Ԙ0\8(P���E�7�y"�|�e�w���dK�,U��H�	۔w�D�Тԏt�!�l��e`@/]�>��� VD�#��=��˙���9��+ʊgJ���DH�(�.�q��0z��U �"J
>�!򤋆  ���F�&q�G�,�!�ć�-��0���9P��!`Q]#�!��Y�HT�01�����Z�!�dJ�c��%�UM6F�uB�O��8�!�D��G���C�38��K��
�Py"��Ld	Q�@��j�Rw)��yB���t�h%�3�D�sC�ɸ����y�
�E��Tǉ�`��QW)@�y�'�guR��C�_2����ѽ�yr� -��ɓ ��M�!��$V��y"*�!T�Zd���
�<S��Ԣ�y�i]#Xq�樕�,t<Ht���y�! �ڄ\���Q$�\詓��y2b�r�2�@d��J�X}R (O �yb�3a`R�k���,�q�jY�ym��8�� ��L�}4ۓe���yR�:w��[�G�RSB} �
��yB΅)ds�q��C1O!a$���y�K4u�2Hҫ�(G�N�1���y���>�� �w�Y�4u�����y"o�G��@���,w8D鑀ٳ�y��WJh⼀�<Ű����
�y�N�jQ�T����n�H!���U��yO���,Q���^5l�P]�&���~r��L��e�=E��(�"b@�ó`8vu�Ea+(�yR���wnP��IJ$]��Us��ū���'(�r�g����<���Q&a�TcT� �c�$�9pj jX�L�C`��V8%�c�� 9�t#���Lؔ��Aĺ@;0�c̷B�"�͙:D��#�c�'#��	�[���x��U�
\�)ÁQ��<�� Y���@�IU^
�>5�0n��!Zj�2"��%�pyHc�C�
�$|���"q�q@".�5e>ر B��O&��1'���K�kW�ys�<K$B��03�Ϟ8W�~ɋ�4gh�D�(cM��{Ǫ�/z��QƆ�8�.JnϢ`4�ʷ釋n���pUd!&��8*F�iX�<�!R
l|�H���ϵU��*�h��/$�ȶ�̕zA�`;�ߪ#�!�b�Ro{�@�WD��S����(p��@��S��:#D\���2)1�O-ʲdŕL�z�QS�Ǝy�M�Q�G�FU���sj���a&x~�� 	��=?6�8�'�z�A��	�NY�sc�{z��WaL5%����ŭ٭V5ظv'R����ʚoAޅ�5�Z1X�l(�!-ΩI������;�d�5&�8z�~��M*3�ᑃ��\k���W�F�"����#ɒ1�L�f8+r��KP.X6aB��^*<DԨ"��!=�Q�R�$`9�����/b!���P�*R Q&�_�/0R����y5��X�	�Q�}R7M�Uհu����
0���+5�Z�u�a{2F��QZ���9A6�Y�si�d
��e�o�2�;#4:�R�r��XB��&����w-�P�@��DC�"`x0h@��4��T�g,�w�����ўh���!e�X�&N�Ԉ�%�+x�|�k��|Xȉ1$A:PV���J�!�.����]�0@�eԨ~�h5IxPƩaÄ��<_L�2��a*�{�L�)��Y�K���8��3R� ��f��D퍁uN0���L����I���% �\�V��!Z8b�k���Q��$� �7nr�4�U��8���!U��#�t�N<i��F�jdᰢ��D� ��݋e���9d�ǔ
#�
���'�Ι fC�dD�+A��	b���)���}�쐧�+Y��Y�,�2V�����`�}����.XT�ay�&��/4���$XR3�͘tPc
_��U{��&4B؀�I�2��] Q�Y�&ٴ]R#č�?13J�F�? {��/	~�,LlFT�N�1��Oz���'�1��ƅ�i�8;1�WI��C��؈�&�9�z���� s<�p� Ȁ�/c7��/5�$�`N��qe��w��
�)ë4�4��ܜ 9ˍ�T*�� ���!Ƅ�Yk҄AO�rO�X��jP0�U��(�N�i�X4&j�$A�m@�/J��iժ�0DތAr���`��dYV��{�-ص%m�8y���4,L��qM�܂�_�A3T�)dN�l�*�*q�[,lX��y��F�jT�&��-������B7R�	�Gg2�mִ)�l@����u����E#�N�\�!�JF5)2M�H
Y9��tn��(OT�)��ƴ.�a@�J�45f�Jr�Q�dր��w"�3�nH+���/ ,) �͉�}/�upӪǵ1v����e׌�]dʤ:֦L#�4ʒ*C�o,,�5��an΢<�f̒ ���Çm"ӵ���bf�9��=5BI���g���R
]g�
��$�B��Pޖ.W��0fi��4Cq�\�e���ZJ�f���SA؁<t��A��EX�,�z�����'
p�N���+$���#�X ?|��)g�]�"�R��N�>�`c�N2��8�B��h��"46j�Z
G!�����O"Hs0C6��>95	�bT����H��T���v�V�>uX��Yk�Ȟ�l4����tP�n(C�LLk��g�q2��]�Z�Q�?*��T	d	�O���Iչ=�ћBH���(O�T1	��6����eҝO�`d�aLB�	v��##@S:��NF�"���A�:?��AJ�hh�Q�/j����A�P6��čY�Cpi��@�p/Z X�D��(O�����أNn8	r���u(\H��	MՌ1ŗC��8�6��=!�Qrd�IUZhmpo�2m�l����$E�(y�%�E�(�'�Ix��Oo�C���*%��[��i���
�5����2cF�؆���!o�c�hɨ!��<���M���faUB�+֤~�JxKb��>&Ԫ8%Ф�`E���%��I-z͒����6���d��;�:@Ӧ��H��Y3O^0K������m����NΑ2��)��^9�:t�k�2M��<�;@�XQ6�M�@J�ES�F�<�'m6�3"	W�'�b� �)\�	9�G��p�v ��W7]�h0��srj @7��1!lEå@ ��-y�� q�r,롂W�_��'QT��N�;�@8PE�.@�S��dJ*@�)��G�ʉbE�"ʊ=��
�q�@���I�r��2�S�	�ag�����$h�=)��б�1t���ʀ�ýZ'(BFğ1oy@���Ny�ػE��#gC��Ƈ�=蜭��i�Y"$Z$�3jrZ��.�(
�.P[3�:�ns@�_/ �RL�����1��Ͱ� aXa�N�@�,��@�Z�m�`�"�E��KDn�;��v	מ'l p9t.�?D�$�� !o�h��;G��y�'T��i�I���P��I+0�d�3�J0LꐅI+�// �k���88� �T.�"����"�Q<LB���0M蘑q�-**��
' �ɨM]fz�%��qܒ�(v�S������3,Ch���(=��zUU$*;�"����@�t0��(OQ��D���0�Ȍ[�Ʊ?��dPŌεm��?�ck�$c�T��	R�^��:�Ûi��Q�xds姗-O����U$%l�x�[�j�5Wsb����IJziD�^�r6��S�$���'6��A��9%q|�5	�E��a]`��m��"|
P�E�@�G��1�J3�D�{RG7�u�aQ�({\�"��qb��n�V��K��c� ��$�F(�ei� ]����1W�{T��$C_%S���h��dy�gaTJ7�YU	
�\������&}@��,O$P�Bg���ԨЏ�hV�Z����:�%���|@.X��H�p�Y�S�_���`"#Ǘ,?n\�P�hW���
L�0wpղc��!�z�H1�Ix�.p�d��b����"B`���
�.+�&��&I>F,P�+B0QpuBQ�̱ga��c��*'Q���v*>CV�`��)��ZRe\~؟�0�h����!��5R=�D ��Q �6�z@q�!�T@^�p"(���a���6��j��Vd9z咨�aJI�\!��lOd��0�S���]��	���f�"RjN+q�Xh�@�����)lG)'���7�i�Vf��2{^(��j�(:��Y{�]��Kb�˨s�r��\�£DV(��O�T�R���(#����>Nn�����4/^�Ȋ7bG>!�V�s<�f�@��	,x"r�;i�91}.��h�6\���I*�lJ��ʩy�1hJE��ɺGR@�3( �>[.� ��0�sT�t>=�SE� n`d1pǕ"1ol�Q�@�1q�s�� �EH	*���4`��_�H�aD	s�0�!VE6r��n�DD� WNC�a]DT/%ud�
��G
%+^�c��1,'�=�C�f�1��&��Y����A���hfRA�Q3_l����'!�-Rf��M��P��G0t����7C�_3�E�t�ʖ�b4��M4*�EصI��tY	��t��̨�!��d�ʗ[[`l ��N�s�Ȥߜ���E}�e���a7@�	H���!X?����	p����%=�h���K�l�:��`��-M+:`�#�
&)R���֫��	r�ڔ�'9�t�b�J��M;w���N��u'��R�q�#�P?�@ȝ-8a���5ʎ�\����O��Ţ�f��Z��4���8H �Ɇ�F }���r��Gd�� ��Fk7p �g���tlY��L#8�f(�&��"x�Q�<ɖ
�qB�Û�aǸ@j%�o����`�>�?V�؁r����V�K�*^�2$[�%R+f=�pc�ؠ�l���AB�-�6��ED:�-J��G
+,��
ϓ8�=b����o��tK���-�,����`������6	\I�r��	G�qQ\�o��|kѠ�)�>8���]�b�����._0=��-����2�lP�▊
�џ�j��RMB�L(�ՊY/ l�G�Ϭu��DR���6����Uz��
�/J��?)+R^O��SŇ�/u�`[�k�2��U�Pv��bG�K6e�4{AL'[ܠ��3C��G���'��I��F�F�B�	�, e(���䫚6vtI�����)VL����I��^�&��3��la�(KPb�y�MS;IV�S�,I�����D(u?R1.�2+ �S���5K�p�r���"�2�0"�:E�y��G�t>b��
'�1�7I�f�
7�^3и1���Q�x!�0����%Y�-�y���7�'l�2�'D���3!��Ed���N=��#@K�� �dʄ@��p�K�3:��zD]�"K�D`�(��� A�K�F0B����o��]���I����&�ۗL�x�@�a�[�? ��c$��s��X� A@(;
��F��tGl+'�̧x�#�n$�����v��L�p��*=����pOZ,�k�".t���R�.?�K���an � @���@V�{�ʜ&Wn����:jUۓ�\!��xh�x�0 !@�6:&��Qh�T��7�B3�A������"<�,�ح�j(|�H�a�puB��*7�RA�Ҡ�	1+M<��B��L*S�<�%� ���i�C��F�*�6L��H�@���B�# �(awd��dWT�;P�s���[� [�Qݚ��e�;z�U*W�?�Y�.��%����9L��90p�*kFr�ΜL�T8f/�8B�΁zQ��.�L����(sɲIU
E�X�AK�����	gK�%8Q��x%����C@鋜p��U��%�Q"Vu��+�2���i��'<W��PE�M�B�=f�CՀD�`��!��L�{��dޔ�I�+�~��u1��j̼�mؙr�Pt���X�`��p 0C�J����Ŕ�2���t{"4��M�S	Bl��ꈿe�$$S��I�%9��3B�<w�h�%II�Y���@���:'\n�'��\����U"4��s2EG�}p�@����_���2�	�'W����Sn�����1$���eJ�=�F}+��'�D�CR�*�r�K��/���+��տ!y�ʱ솻%�\������'�O�P9�� W��(c]\Q;�8�.�J!a�a�H���bFX���'$+�b�Ub�����.CY�!���+K29��A Di�
��-�ല��0M^98dF��GU�	��)N
"!���@`�j$dY�B"I9�l�=geጏ��'F0��PdF8�dE���8�A1;)ad��h���&I�KXţ��]�樺Aƚ2fkK�R���)�V�<�z��֬��!��OLMBVKCZ.2;rÅ�"�0@��f�>��bS1"3PT*�!6\m֫�Ѧi&$F
�M�\c
^mz��0U�} NՇ#Rr�
�C��%� e�De0%|OV�:�ȖP������7M���W�)&�rih�����)R�r��H��P���AS�MBh�&�Q�/�QD���*ƒU�diB�B�PڮM�w.LO0&�D*i߶�cG�V3����h��mK�` -g�E��F�=x��]8q�P�eT��&�/o�����ކ�]V@.b�Y�R?}�����WٲY�Á^�0J:��xrǃ�d�P�n���T�J�6Ju2��f 
G�xAQ
4 ˈ-)C�،�DayC���*�l+��7z���A�2��*"�5$I���O��?����CS8Rpbpb�1�f}���@�X72	`���$�����9� ��U�҃Q1D\
���3�te���@�y.X\%�.}�BI�D�	���w��W��ɒǈT�(OJM�$����W��^�������k���
�*�_<84��^��*1��k߯W��h�CZ����Jғn����ꊇ^;6(Ʌ��(��Q��L�??(��J2n�":}�=��@���T���,g���QGՐw� q��G�$����rJ�Œ�,� +�8=Z3��W�@� �d^,z�0Ȃ)�5Av�3�-EvC���Gl�/�2!��G:Q�VqD��-�̓��5L���A��D���<+
�q��^�0,�/ڛ(�؋�@\�O��3���D�}�'b-B@VLr`��F�f{�'z-X�Z�D���8d�F1ew�e��"�/DKB"<٤��m����Ӿ��A߅JрH��+K4SHy�I��OC�nD"E��E[+�.}�Do8U���HvM�ÁF����a�e.<TI�@:b�AN�'[�#<���˷_p68�2
q:� C��$o��Pȱ�N�'$��Ḅ-Mfh�voI�������#��bć%m��ɋMx� �(����e�c O#�X)�".~O����+�ͮ|I��5N�$9�,P�w&�ԂW��^�L����yY$x@��,F���
�%3.Dj8����Fb��z�O�i"#<,8,*��V"~Jj��2�� 3�ܣm���������>]���ўF(��v�Z
p�qa��+q �	�"]�h�����`�<U���Q�D#�5Ҷ��=,�:�R �L��p��$���BS����(J�KtE�	�s1T�Qe�Pk:ظ �r�J�0�CUN�8�Ƃ�Dޥ`��Ō50Z�@�兌Wg&��@ĝ
t�V�pcc��u��2�%�������H��f��x�W�y+`\ꃆ! Z��� z���J��cPq�A=O� ���-sU(�@�Őu�봡�"���"w�R@?!���g���X�K�*�w���̱w�@ ������瀁7����r`���-��~8�o��J�ڬ���о/�&M��,a��e*���
	���2J�t�)�����o�$j'���� 7f�`a�e�,
��a��B�:_�h#�o2RȪ��]$k%�˧XC�da�w�$�p���8�rS3��!Jl��';��+c �0��wAњM�j=�0#]95	i�N^�s���Kֱ9ƽ  �4��c�T�2��/~����+'\��dI�j?LOF	��.�/{d��k���8Wܥx�/��:��qI&VL4B�M�t�rX�c/������G$D~�Bc$T�a��y��c�4�qO>��q!�m=(�8��W"����.������O�t���		�SQ�mZ��G3	K&4a�'<�T+Po�3\@u�� ��BQ�Ë5��5�ѵi�����#�px�F�I�[��Yf���v	��gp����hZc�<Y2ώ�E����fE��`Հ��LP$��$A�*jW����a���"WxQ��I���,��8��F}�=��$1D���Tc��wz��+�h�3�daT�o�h��O���>���߶��A[7bK.�BH
QmV�<�%Nu�,;#��*CR�r��Ux�<����?�U�Rc�lZL�
b!n�<ɗ�ʿv]Fq3���<l(Y���v�<Y�'��*(
8�c�ڄy4RD/�w�<�e��0H�A�g%� ��j&EKp�<��oJ;Znx PQ��0t�Ćȓm�>D Ҏ]�%���FfJ$`l��ȓ*�R�b�S�VI�ʁ�G����S�? ��� ,?hD�&��
JZf���"OLU�dH�"u�t�ԊO�(^�x˲"O���dfX&F*2a����;s1JyA�"O&�H�EL�B�	B�'�:3��y�"OJ�K!��Aĭ� ��0+���С"O���w`��r^"��d �?dU� s�"O!��3���p�Dn��Q"O4< �`�1Fz�#�&L��{"O����t����*@�1!"O���LȌP�xU�t�K>T��'"O�@c���Z�����U�Q�+�"O�L�u�� m���+S�Tce̱�"O6XЇ��@ִLB2gЖjg��r"O$����{�j��f�Ő(@`}�t"O��`d�=7��$	i���y�$ɜVl"��C�]�2��9���y��I�z�����]�6A؝Q�	�y�8N+� Y�E6+Zd@�&E��yrN�I��ppj�*&+d���Ǎ�yR�G���yj���o
���$
zf�Q1JX$1E�<qFѮw4�y�Gʘ"q���3ͻ�=�f%��y�g	��@`tn؀0\����BO �y�⊶|���!�Y.$�d�ڤ���y"��	 ��p��N���𓄠H�y�%l���+�	���ܘ��A��yB�B9p5l��-� ]�B-�S�ς�y�C���4�1���T'�Lb��L��yҁP,Nꔰ��`N�L����(D<�y���)�00��=W��i��
��ye��
@�� �� �R̮P^2��ȓ+kH@�Q�]�7�ܤ��) ,����%�r7@��n@���@�1��ͅȓn�ѐ��F�vU�I�5wO�ȓu�F�Êp\1)g�Z�~����ȓJ�|H��Ŏ��"U�T�K(���ȓj���s��D�<a`�S"�\��Pei:�	�s��|� DF�Rd��7��DnZ�[A��H�	��7���U���h�6/~ !���!l\��ȓABF`�5�V��%� �7h�0��	�:�����u�̤ qBT5)@ޥ���0,ӵ	�5�(} %M23����ȓQQ��ȷCRS��c�'M� �tt��5�d��E¾4��6LK)?R`ه�4$�q��(�1L?��{�#�`:P��4�2�w�
���"��4F��ȓ6�6��eJ e�ᡔ�P�؁�ȓ2�$4��G�\�l�!�؎�M���0p��1���qf
�|�.чȓY���zT��9���� �]����ȓJ��P��@����%��P �ȓn0���_�,#��Z!��	4.���R��qI��^*O�<aHOE�e��q��dS��ST�T����V>R���\� �	�  >`:�
B5s�^�?q�����Y���D
HU�y�	�|x�"o�=v�ơЅ�P=G X�3�"Ov�̰['���p��~�,87�O��8�d��k�|��mљA��HcCn(ҧ$3|� p !^�fiC&ʚ��ȓ}Ĩ�q�X�.!�)a�̝$��H�SI�Z�����2���K���T�)4���z,b��咆D�УS� g�(���
J���Q#Z���3��\�ij��EFI��4;���3��Ԙ��0lO�8zV+�L�-��s��:����'5`hEΠ ��x�!��C��9��K��,Y@)��x���O��~���ܲEM��� �S�S�B���P�w��-�S*��$`d9p���
$٩�'L$�Ð�Q�>q��O7VM�+���� NWΑ/>�z�R)H6d���D���� B�,Hܛ�ةcb�8��� >�B�
�NqY�$*�eA���c*�tk��e_�B�VqR�芪~.B��������T�I6Z��VSe�(`�%��rL�b'��<-�0tR��2O�42���R��x�g �2b�P��٨;a�ˤ���ai��OF���HMd<�<���a/�1�n:Z�CP�YK�uF}��0sPh�⢫E ���d(H�!��X�$=l��E��M���ס�H��
R�ײ>T�H�D� 9~Z7� ��ugcH=n�4l`��N%d \c�z�#��B�'�t(�)Ƈ/����r���<���S)�>}���F��ȐAt���?�;���h��',�Q���+���Yriܓ�(e�Ʊi�p0��e��}�>�96��S(y�' y���7��	"�(�s��^θ��(ك=KX0�$ʜ�=�l�'��B�h��y��A-cT�!�O&��pT%�7x���M+}���.ݢ\��G��p<�fH��{:���(E�h��І���� ���OB4��L^�<���[+3ء�1X?!(��nӪ���ZB1`4�P�j1D�%��r�Ȼ��4�c��K��
�X����N0bXw0AKg�W�u���c���@l��
	�ph��O	?�(1ID�i)0���Rk���b�=ۑ
(i L1��[��J�c'�>�Z=!�O*��S"�8{A,�#S�*%��A���	��D	���z��8�B$1�N��4-D\���4�uȤNȫ��
$��Tu�8��K��O���0�H�xu��JX0$�8�J�Ǐ<H�@ш�G.��;v�a�:O��0�,�fb����8���%rLq�1�͋��ċ�R<���X&�G��4�Uh�a�}��N@,p�	�U@��<���ʕ�y�����1��h�~
��
Ԧ	����=K� ��o~�P\1x�h!{`�[x�V�R`����!3��%I��U5i�a"��.|wb�;-�!.W�uѦ`�"*�͂�/�G�r<n�����Lԗx�t J�Ծy�&EЂ)���f�9F㠴�6%L0��$���2-\TN�����Z?-&h�a4z�e��?��a�p��I-N�s.�G��M��.� 7��Qi߇Y��)�'�Ҍ_h"r����=D���2�8R� �A��0_�qD욜o#�!1@�����y���A�vq�L�C1��K�3��XC��*������4T�s�#��L�
�d���ޕJ?N��g"C8���'w�U���#��L�^:n����K�/��oZ��TC�/6�]��ԁD��	�cX.d����ɡ#��kH$x�`�ȕJ��o��4�Tt)e��	dL���U�ծ)�f�	�KT�>X� ޴]����.�n���SH����S�Jh�e���vF2�e댈B@�*N>a㜨��(¨�����kc$�~y��8:7�.�̣�$@�b�!�[Pn�X�A�ËX� M�T࿠p�f�-��@Gx"+�<{�ikGI��2�&��B���2Rɱ󉌖6�i)�m�|y��<�&���M��0�#䞎Pz�X� ���,�ї$�	_��JdȘ�~�r��5��?=�r��$�>.` u��,8�`�%J��05H�'f�,U:,���� ���j�P�7M��?]�'�R�brʵ�p��6�"V�pw��C�� ZЅ�G�Iye<yt$�C�d��%/�-�܀��ɒ�CO��q�HW�zr�R��l�$y�S2y�������C�I�a��06Ȼ *�9ˡ ]������a>�M�L=����iN)#S��	�ʍ�\���b@�(0$�jL߀.;�Y�v'B�&���PKڢj��x��/S�b�T�P�K��OxQSWU�H�����#IQ mxg�5EP��� 
�,L@<�]��9O�D!� l�&��B���&qp�+�#ܡ2��tRҪ�%�� ٕ��f��<(��_�0>���`��‏-��Q.�k 8�䞠�y�@��������h�(�⁍�M���+��O�VL�ғ�Z1:����i�s�����*l�9)��_��R$�'+��P��C�'&XBQ;�+D �" �At5TY"�4��dGF& �x���̠����F�D�
���@�SBN@����/�R�ա�� �녡0'�������?��O�H@�)���3m�5�rY�f�o�2����<0�L��KCOU���&�^�|"<I�炓n��X�f'�(|Jy����4�.9�!�-�r��Ư�o���O�)L� yH��}v�`�N���u	��D1 ia��0����k=(Bf�3c�±;&����l1�Ё���t�l���`c�Z�cEbyE��nJxՒ��7}�z"��25�Es�EϤ+َ�A♨�Xls'!�4`GV��$
�F~�FR�)@�	�M;���V:� 6�"�D�1I����T`�>�V�9�@�)V�㞜I$��<�HX1m�B�,���J�O��'?@� JH
'Һ�&�V�x�ౚ'�6MJ�3@�Ԉ��;|�~�2��T��Ⱥ��G�C<d�yf���0���gH��iz�;�KƸ'vX�	���џ�g��|Z��E�M�:�����A	h��EŬ5J^5ڀ�C;�X��ĕ�H_ �"�������eJ�z\��
a�J���♜ߦ��Cɕ�����mM7+Ϡ|�F�
�p��!@E�[�1��z(L�$�PP�Rn\�u]�=��e�X���[0&�+n�2��t�2H��p��	�E���>A��)�b%�K�-��m���<�qO6�x�E��,�� �n�
���D""  a�|��"E#���y)+6�'bT� �ѨOB*�򷢛�d�fd�$N�@ �� �
?���JboV�p|��Ɔ�V��U�$��l]?D��҆ɋ$���B�\7R0zL�+-�I�5(]!j���q+�WA��g��?�:r��@eT�� �:P8��'� �a�Ëq`��8v�4�����o�����I60�R�`��'.z	����=��O�Y��A�e[>Ur�yҮF�1��#'�;>��`�bC
ܨOj���K8��4l8���W�J:�'W8R����K�j���Q�L��#�!\)����3LO� ��#V�F�Y���ȗ�|[a�O�̨��H���	"�n��Y �e��?A��ߒ7�������
r�4���X#X�,{��<�O�����M q�&)��`�WļJ�O�1Q��{�Uڽ'��h�Qq�Û
���)W(�?1h��	`��u�ƈ�'$�lT��)�p�~ �s�_7`��\2�W�i�'����lo>�F�/`�n��4O�PB���:��恕'��������*jL�K�G���/f@��ZI�$<�����[�(:�eɧ%����Fӑ]B
x�����ޖ}XU
Jz�'?��a�B�X�@	�"e	F�ڡK(Ob$ !l��e�<h��$�X��/G ¶i����2`����~4���"GX���4 䎕D�(�C�Νn����۽E��v�M5C���6�	/K,���ɐ.��uq`J�
l���D�ʟ]Œ�I��䌇�y��(U����"��V(-�C��<��Oq��uԄ]a��%��8��;O�$`7D�$Rnz("e�T	6�z,��O rK�mb�w�� íƠk��%b3L��?) a�D+r\j��2OTH�F�M���hY#
�U�� �?!®Ѿ$Ö��4�P�'��*I_ɧ�MW�L�IT�C�pU+��R 2HB��
�T�{ F�3(��*�d<l�A%�CN��eJ��C�&�ݿ*�$2 ��.&D�O�%0�{��7�ѧą$��-�>V��aӲ"�_�J]�E�0LO�h[�cs�)#�Δ�.I|4��3n��x15�r�Ԙ�L>�`n�u����>i�Λ�!��;JR\Ǉ^Yp��כLR|�G{�¤T���#��F�AT����.�4�yr�уP��-�Ǉ�51G�ͫԃ�[��=	g�iq���&R�����Qj�銸cP�T�EE�>��  q E����P�z]�4	ڟ B=�\�H�Ƈ@��|�D�����4�� �"��4%����iù�Ji�t�eӄ}㔪�P�>l:�#E	-���	9�(�D�
�1��JJJ����
$��A�T�ᔨ9M8��'!�S�[�6$�ᡲ垳N������3L����IV/w��8���'t4��af�?C���`cbI�6�L:gk�51
k�fr��U+�O.�pR�P3ؐp3�R�!���_w�2�H�<�u��������?��&$�"�hO�(�d͔�G���`#͞x�K�0O\�X�A�*L�T�q�['%Ϟt��5^t\���U�:�>uS��A�<@��Z�I�5��u�KeO�uȯOt�����e^8���N����'��Sbm�{������+>nt���'�9��?���'��D�ߧX��0ⶃ�'��<{QEQ�~|�c���Q{d%ԃwP#?٠GR����J��#^~���R��I�4d�E|��eg_>)8�۠O�����=�rIh�6]R��FA�>^��0�6��C��<�3�ѱ
����	�t��M#�yǦ}��C	���-���oӶA��l�%��0��/~P|��	��G��X�#�Aa�����ݗ)[ �y�����d��q���Ò�P
WRl ��	�"�"�1�bM�!q��b
ֵT��E�lM���x[ ��k��K~� m��I �A����o��k~LS�������$�D]�O�Y��H&$^&iӁ%Ŗ�>1���'
�`@fm�Y�BM����IM�X���"Z��M��H�#s|�P"�� D��W��E�D ;��ɀ�~�?���??�4y�Fm�d�tH��JV���C�7*T&YBA�&~��q�O^�0�p� �5u>qFi]����.��x�K�
gߎ9��Iq���$��:aS���;��ic�h r@T��n����W`�V�$�2D����w��.M������C(���!��_� 䪑`���
,q�0���5����� �*����'c1.lp�ؤU�](]�N/���[����� )Rtx-O�>ȶ�%�����i� ~�T�y0��O��R����8v	��A��G�ʲ>�'8�8�B]2I�����@�}L� r��<�s&�3�vL3#8�����,<���݈K��8aUQ)I��Pŋ�Q^ތ���3��P-�F�'�ʩI�h��Ǡ�r���]FX�aH�vcv�
w
��z��͸'�����"ȐYd%B�*<��f�l���*�ɰ�"e�ƛ>�S ��,D����'c�Y�U��!�AI��X}X��G|b$�+3�@q4lOh	VI��pR�I� L`����6B���ADKp}��-(�����Lo���?B[NL#D79�5{��&9}xC�I �H���˭8�����H�0�xC䉃p���Y'N;k�P�q�F2jRC�(2LC�a�=x�z8���jC�	)k�]i��
9�T(�MH���B�I�,Ե����}�8�j�m�D�B�4H���J�͎"A��s���3{bB�IK���)Ԫ��#����>֘B䉲mF����T��1
R��B�Iv�����ߕ/�`�fNM	*��B��?n���ϛ��.�tAA���B�I�M�L����Y���`����@=�C�ɄCL��^4���T�ޛT�RC�	!t�A�@�@?~�G�[d_8C�ɺN�%;&�4s�(�*����j%C���51���
> �HEӇtf�B�6g�Lh�ϟ��"�Q4��B�)� έI�Iý��`v�JFf�QP&"O���,NGHH���	7W�!&"O�����Az�0A��x@5"O����K��F�s��̇MD��s"O�{5f�$�P8����T*}C�"O �`�B� ^/��b�-�$)��&"O`��6J��J�z5��ꎿa��,��"O�p �A!<��l#�f� %��Q"OA����i�ڜ���Q�sՎ���"O���wo
�O'J|�!*�'�t�y�"O��Q j���ɚ7�H�x�p�A�*O�T�P+�f���	�g�]8 (�'��
0J�Pr��U� P�L��'	�p��C>L��j��ݨWA<�r�'�z�JvhǏs0�+c�O�:��]*�'��iV\;�y8ъ��B�m��'�B�3�܎*:0�`�A�n�
�'�2  ��^&2��gO V�Aq
�'�~��AȈ-��$K&bյ`�L���'Ҵa�9J��D5d̚0�Ds�'��0�VG�1Rz��X�G����'Y.���@�����VjIw|���'<8�Aƴ>Rz�Yv�!�p��'�,�2���"�<A���(����'��,�c�:v?0��Ql 4	XȌq�'.-:�H�7��P!��$lZ�P�'h���e@#;(��ذ�H
R�V��'�֍��ϔ�,��a m1{�L���'����k÷O�$D���߃hKt�j�'v���pI�� �ڝJ��|РK�'�4�Ǥ0E4��&F�8ǚ��'@Y��E�@�8e6��`�v��'���#�)P��f��f�@�1�'#�!�	�	f9h�#��Y��A��'}*i�&���C����Ox6�8�'�HQ2��_+�@�Y3>�vMa�'g�	�C�trf��T�	J����'z��)Ǎ-|��9�Θ����+�'\:��Io����ɉ4<0���'
�U�S3�ܠҺ������z�<���7�p=�_�"�i"Ս�\�<	�h�)�P�*�%�;.C ���'O[�<�Q%�ȭ0Q���ce��У'T�<	��(?�*p��
�H�&i0'O�P�<��
�=5����M����ۄOg�<���T�`E�]Q���6|Ʈ)�/�h�<�Q�+*��D���NA���J�<yf���R@R��C3͎��u��<Isƨ\��)�ĈVBR�;���P�<�5I�� ���^�;4h��'O�<Y"a������AR
iy]�&���yb*�3��]�u�9^~$vk��y�‷W���N�)O1�܂t���y�Ռ ˒�eo��LxXE(W��ybퟱw $݋UF@��
+���<�y!BR�¤�����{�O�*�y��##V44
3#���kD㞺�y�͚
=�y�Ήq*x@���<�yB��o~����ŭu�<�����yb��76e��J�	 ZZP�au��,�y�%\����E��U�`9[�BZ~�<qB�~T�ErPf�%]��X�Z�<�D　kT>��� "u���dNRZ�<iB�7��a#��I���R��}�<� x�(��L�K����� v�)�"O�h���_W6�(�%L,z29*"OT�"��� &È�9!��u�B�x�"O������W:&��r#�r��a"O��H/^4Є����äL&"O�({"P�R��Y�5��2�B���"O΍�&Ɨ�/�r�)�bG�p���""O��`Þh��ye�O'g�M��"O�"�k!Z�E���&8�	"OTUkS+� 8cl[�g���Z@��"Oj3���4�d��>���2"O4���̂L���rk' h�Ha�"O�u0&��Wl̑�vi��W`�q"O�xq���=%ʠ���%�H���"O�d���4;`�ѥ䔵{F��k�"O�a��ǂ,����V���f"O�0�G��93Hq�e�V�IS���&"O��!LP?  ,��g��1UV��"O�hBq�\%^��ˣ)+Dz���"Or8	��8d��(�,$-@a*O8{3�Q�,�̀qT�C�$��'��]�)HrL���-�:WM���	�'V��'h�7Y���E��]xZ��	�'���I�Oőy�֜��lI4V�d��'8��+d�S
Et&���߼d58�{�'PdI댭|Cd�*�&W5����'�b(3.N d�<���_J��'��l1Q�-H�����N����'K��Iʦ9��	�j��D�ڨ��'H���5KO� 6���ጂ=�E�'�T8���_6g�x�Yf�<��Y�'�����>>G�h�d#J�D8��j
�'���R�	ĸ&����V�<�XII�'��qsc"	��*���l���@�'V�-�р
:y�VM1�Mڬx=T��'�Z�b@�/���2�H4B~t$��'ܤ�R� LzI��9~� #�'��H3iƐ[l��Brڵ�.=�'���qᕭi6ܩf�ڵF	���'n` �-�ŌQ)�lH�)K�')��X���#���h$T�J�<lX
�'�
��R�-E@�ɶ��Q"~�K�'$��A�ͪ@��8�pbI��=�
�'�t��
2�ѓ1��l��'��`�'Lg��, �KC׆�Z�'��z0��0��"� ��Q�'�����@�D���R�C�k*�i�'�P�������{�
:m9z)��'�2�{�:� �L�xz��9�'V�* M��7�n����/rL��'#���[�r���K�m�	��'���6HZ�"�ڭ�T�E�赊�'F�A镌W�p�V ��B6� ���'PR�j�
�{����Gj��2m�}��'`�|)QC�#5��a��
-����'3pk҅�3�0I`'iˇ%���!�'}ڰr���`�4l�E1&��1�'ŮX0 L/k;�(x��@ (cD4Y�'�Ĵ�PM�!�8��0&���v�;�'�H� �]�f/q��M�&r9q�'�ʜ�c�ƈ9)�}�2�[J ��'fL�P�)ەjwt)���^�5A
�'��<CGb��\���[2�^=|˖�a�',�G��.`�13KVB���
��� �8၏R	���1cZ�$n ���"O���V�c��P��؃8�>��f"O��9�jC�+=Ba�T
CG����d"OD���$N�E�xY�I�n��"O�1p�#�6�n!pg�	�@�B"O��mO�FǦpJ!�K�u`@	�"Op�NS(:&�L�F�Vn���R"O^�I���:/$q�o�.MV�x'"O�[��K�2�,P��11.��t"O򄻡jT�8��f�I;|�EX�"O`Dx���3i.��DP7w0��v"O�eXg�#o��Q(� +�IyE"O��1��p�E���F:���
�"Ov�@��6Z6��hAz��qK�"O������3�����'�
mx3"O��!�ʇ�q�$��$K��H1*@"O� "�)' ��q��J�b��e"O\!�5�VC��]���301Й2b"O.]���6FB�rF�!f��-7"O�h��X�U���tg�]����"O����zr{C%L�C��i�%"O^�{��S o���"�B�8=P�"O&�R!�&H��Pjs �1s��M)"O����ţ���*3�Y�q��pӰ"O����!%���#��*��1Q�!򄙗3l(�bS���48��,�!���c���Y�ؒZ��cS�шd5!��	�K�� .rk��\T!�D^}�БbS�
��a���GqA!�&�Lh-թI�ؑh��Q�V#!�Du��#����[| e��E� G�!��*܊�/з�ҩ����\!�DM�j��Qq��N9R��X��$��TaB�O��a��>bθ0�h�+iČ��"O��(���jB��@�:�=���	a�O)�L�U���TAa�.��:��
�'�ָ��Ǎ�Jb�-H�	��$�
�'��P�A�Y�_��Q��-0*Z��
�'V����G�#z�DU��U<}S��H�'1�$"�C����R�\��<�
�'���b�d����A��M+���'���!�*��<��(R\*z&�@�'��@�ᚽ�H�;���A�8��'yj�#���9�B�h�	,e�'�����ĽM���8@���J6(	�'��໧�zʔz0C�*���	�'��sE:V�Ȉ�A�9�'�nd�
G8][	��
�:@��q��'z�=1�^���u��h��H\8 ��'��P�GEʙ����v�0�k�'��5��
��\G��Xd�>"M&���'v츃OW3܍CF V�L)�yh�"OT�S���5�X� ɣK�ZMӴ"O"!k���=�,����ߢ�'"O܍�5̐�صJ5��&q݌��"O�P��@2��Y�K��c��8�G"O���ק�;8�V��TK�y*�\�%"OP������L���(C�L$�X*"O*��s��#�I�1��_�9	G"Oh��Bm�2�L�X���t��� �"OP���e?dA�Gʔ�D����"O�I9�B�HQȽ:�Έ�x�0��"O�Q�
?�$��!�Ѻ{��=C�"OZ�p�L\�(��m�|�Z�0"O� �
4d܀[P0�:��M12�Ƚy�"OJ`ha��w��!RJ���NT��"O(�{�մ%$��2`2�8pR"O�Ѡ� � ��PX�n̶&��!��"OT��@C�|Д���JI1"����"O�����Ҽw�<٣BlR1b�n)�"O*j��_�|��M��m�/B�⁒�"O�H�Eb[#���I��8j�ȁc"Op�C���u��
�8=�"O`�;�E#	4,s��L�A��"O����
����x�&]�a����"O�s��j^yᴥУi�d�dk�<IN���z�A��;l��� �P�<�0�E.:Ѱ��"f	�#� ��VlI�<Q��߮5I�0�)E�p���P��H�<�Q
1��%��1[e�-�A�#D����H$y�6I�&�h�KCb-D�|S��ʖ쨙9��ןbl섡��(D�с�:.��uh�	P�a� <;��&D���R�ǭsgX�Dl#R���
��%D���B�;t!XD��j㘍��%D�8(��߿;X0����~�:W 7D�\�'XXr��al�i�6�p�,?D����/�0L��(A7@*�P�k)D��x�GY'-�.��2ˬ.���CI+D�4��(�MNT�c^��z� �'D���W��3,��M�!�A23���k!�$D�����W^�cċJ� JT�9��!D�h�a�8<� (+�Ȏ?��a- D��s���-��)��:}P��V�?D����N�l*�hs!X�@� #�>D�()#D�,>O ����?���q�)D�h��Ox���o��C&D��h��"��Ȧ,L�>�X	10�)D��di�0�Lj�+)f����b&D�����
��!{P�Ib���&$D�h:���]�09��Ɔ�>���c�
!D������-���q�c��4�D@��+?D��XwɃ�i�@Y
#`زJ�Z`�C<D��p�d�������fV�?X�2Dm;D�8���<XMHt��
��-�!*9D��	�	��s�h�2BN�QJ����m)D��F��4�PBgŌ�N=�a2�")D����猾&k� ��t�jՐN'D�@8B�j�h5�T�ƪ.7(|��$D���¯]r�Le�탡$�0��i#D�DÔ/^�68Z�Z����m�f���-6D�L���J�o��Q�2+��	L4D������n�h�F��Y��x��-3D�h����w�N�9'a�'W��pQ#=D�L+�)�����B�!
/.��i��/D�`�g�	8
+T������p��K;D�<*��X�{_�Y�'Ƿ{�f���#D�ܐ��k�ʸ���E&%��E��A"D�\�c��y"���B@�$
A,>D���$e^�)��	�_9a����u�=D�d31��03bn���,�)h��xG;D�4��(�?2p��+e.�����3D����f��HaO��&jb�RF�6D�0��ţ:��$Q1)�$�XX��3D�$��IH�(ԢѡfVd��)5D� 
Cl�"xx2Q)t�'��R�n2D��1��ts���#�ˢE���J ,D�,�Ы1�l��0X�1B�i%D�� N�D1� s�䐷;Bi[#�IV>��)]N{����$^4AP��4D��홒d:���*['؀2�=D�D�E�C�4g�mIeJ�/
����:D��S��� F�[��p��)���4D�tie�S-a�DB�؆=�ց! �(D���Q�%o,y��U����Y�!D�x�@��\��,
�����	p�"D�0E�;*-�S�D�5��X""D�����M �*�s�ơ/L�L�J%D�ت�.�
2�5DD�`��aۢo"D�(�#K�:�d(��,i�u;��+�.�S�TQ���ߪ)�(p��V���W�UbtC�h�L�R�06u��M<P����S�@�$��l�$�ēb��-A���a���+��F%!r�i�B��8A��:"r���`�]� u>C�ɧ����$���=!5��E�C䉤�B�kv�^$�f1!tH�?0�ԒO�7�<�S�'\�VU��A�@�tbA��#�����%&�e-�j��A2���+�@�?�
ӓI٢	���:6L���'��7��\�ȓ!^���'i�V-;�GK�}�����'$�B�����r7�7}�l��0cl��7σB�8�bG��I�n��p�UyB�]�pm�(��|F~��� Z�����U�C�)��Or�:C��#z^$�sF��O����#�486C�	8���&�f8�ħҎ�ܢ?ٍ���	;�$��2���t$�-�%)�2
!�X� !xuwᅷr����
��!�$�6K��
F<TI$�7\u!��L8�MC���	��!d�ѝ3l�ISx���'%\@�a�I: ���K�GO�H|mh	��y�%A�c� l	G�D��-�N��y/?��]8(Q}I������O�E��o#�Ly�Gl�=zW\�	��7�yb�)�\�|�C�ю\����b�{�$���hO�>0UmM�%d�
}b����0D�` #	^-h%��x3�T���*��;D�<9ejϮ&�z]fq3w�K�gVC�I�g��Ն�[�d9P��H�3�8˓���@����O�^��;�"V�jPz�J���Z�!�$���H� U��x؀|��9"�!�$^:�"5b��:3��0#C�'C�!�����%��4?����S�U��!��,X�$P�%,}� 1I6�M)~/!�đ�pR��K!-E9Hfb�I���T;!��O/~=(�bS�N\����:Y�!��Q�f��%[E���z�;࣓�)�!�d��v�����0�h�*�ͅ�({!�ĊArUqpg��f�8�
�Y5[a|��|��
TH-���O<����w���y�덮><f��4��"C8� � �y2�!'�1�Q Lg��h�(]7�y"�X�TȪU��R�h�����~R�)�'j���{gAH�=�$��'b .Z��y��g�	�&<H�Ҕ�'C�fUR�@�=��C�I51�l�g�5n�TI7���M�#<���?��l�+@���cRkâ,���)6D�4"�6b���	#d�%}�0��6D�x8&�O1�@��g�C��8�W7�O�'���炏� 2&H�+&\�A��'Ln1��E�o���Ŗ� ����� |L���I,~�n12D�	!"0l�"O���W�^��x�viN�z<t���T�(�p�J8݃!K�Q�R-2')D����ǔ���49Č)��pB!�D$˞�Rf*�"V�H䇛�;!�D�����; ,Q�k��� %҈�!�$ƋGt!C�[-C�Ȁ�wI�W]���CH��i�)4��p��o��sM@B�I3l�U@faG.|�<z�m�$FOȢ=%>I�I��<a��`ŷcy�|r�.�'`�C��b\���
.,��9�A$4s)���=ғ7�x
"J�S'vQ� ��T����ȓn(���#ۃf�s�g�|,9�ȓIr��jשZS�z�3��)O��X��q�b���r���	6���'����<��'s��3aG��e,L0�l�<	DfϘO6V�*E;�	HClR�<!d�>R `���cr'K��Ê�D!Q-����lK�0��u��(P!�$�#ux2m*����@1�M�E��8�S�Ov�J��-I�`����@;�ݸ�'����A�!E�������噍y�'�(x�dĒ�05h:F�G��]�.O$�=E�tC\>#'.�R�/�'��lR�*��yr���"�q�(V+��p�U��y���;EX~��%�)Fh����y�#�bt�<��U��	����yRD�� �TϤj��J���*�y2E¬l~�A�
�a���R��yr��K`tٳ%)�[�]��%�6��IJ���O�9�����U��y���H�0K���~B�	���� r�|	��H�y��G�TD�� 1 ��m�q�㟵�p=1�}B���el���B�r��Q�3l�'�yg�=N��!]/w�<���KҾ�ē�hO����#��_4F �&�Ej^|C�"O���a_9f���X�/
"|���"O�a�2�J�zL�
�l��/ �9"O`���je|
u��3^`��k�'f�?�ЇF˩g��l��-=,���4D�l��(Z�*�d4�3��7*ظk(3D���e�Z�Wߠ8���+e"�x�K/D�X�����pi���z�)a2�8D�<�`%@ �$E �+����4D��ӵ�Q�@�jP�@�D}��ăTj2D��"4�E*\�ԵS�%3u�,:��5D��P$(�>;r�k��� tj֔uI2D���U�ʃYZ��S�J�Hb�y1*.D��x ǜh�E9G��|g���7i+D��gKԔ:ݠ��HFb��e<D��(��z�$����ړA�Z�u+:D��3�$�|@p����8j��`Վ6D�t�TMϊ:���C�W�V�,�gA3D���4-�^���i�1����C�2D�,+�g٢JXa�P� | �!$D���%cގ��pЄ��'!��ܫ#�-D�����	�&��'&):Ȑ�@�,D�h��J�/�"�[G�ϑ>gX�� =D��y�Ŋ.zJ<��Gh�)�ȴ�/D�Ȃ�EG���\�q��j}$��CK3D����#@:~y<�E�\�`�0��/D��{1*.&���X���	۶�y"�õw 8��e?9]���v'��y�I�3$�`8���*Ұ#�@��y
� �!bĀ_'?�V��w�G��: {"O�ջ���5g��] ֌�)p�hi�p"O.�Ц� j_�ۀʹv�vyb�"O�S��.$�}d*�H��i@"O�pʥi�?M-
���)ݲ=�
1*O HC%GI�ol(bс�7�"���'��i���Ls`k�*\�-��'\|����'��b��
�,`<L�'񜐘v�d¹:Y�hi2��s�<� �
*	o����,�9|�L�;�s�<A"��H�v������s��}{���n�<Q@&�h�څ��eX����u-�U�<I#��4����!�i��]K�/�S�<���TX�M�r� /I������W�<��W�;`<���E�>�8x��)O�<����+#%����)1`��P�r�<��1^���SF�/T���(�q�<�'�S	!�0*I*X���:whq�<�`,�
ƺ��%��"c� 5ѓ��s�<�G�*[{t�
o�'�0Ad��e�<��ғ
��2r��'Ͼ!��d�<i��:܈I`�
�3�f�Hg�v�<Y��Ɲ��ڔ�,Ƽ|p'�x�<���&*��Aq��-1����kLr�<9�)��E�
t�G��I~#�jIq�<Y`"	bJf�� ���p?�
��i�<Ab��U������ѓ-����C�d�<ᕉI��������a�h1f�_�<�b �`$��фP��|(��Nf�<I`@�QVx�"נ݃/��͠��_e�<�VjQ�T��h�5���v`�U�w�<I��j�1�2TT�6�k�+�t�<A -B`����2��c�j�s�F�<1�R�~Z���L��.M �����I�<��dE�"����$K��4Ԁd��C�<�G�^�>�+!L%hU�4�5	�[�<1��'`g� iأ2� ���NA}�<Ic�8ŖU�� x��b�_�<�n�b��c)�fy�4�2N�_�<�n�/2��dKSv�4��(�F�<Ie.<��T@�Ȝ�&�pY[fCW�<���W�-����2��k�v��&)�a�<�!��@�A����PO�@��VF�<Q��J.]�t��m߃JR�"p��D�<�E��;K:B	@wf��tԼ�0NU@�<��c6w4~5���Tq���~�<���4nЉ��ڃ`�N���|�<I���$YE9���r�w�<��I�
!��K� H�~�*����q�<�v䄪$>~h��%��-/�cv�p�<�5JҜ"�F19��@�	��\k�$�t�<�UlR8E�p��g�΢2�nD��!n�<��c̜4eR6iԛ7Pe�S�
j�<q�Iާt��(�q	��n	��I�D�g�<����H0���N�d:40GL�<��=M}|�"G�ʳ�f���b�M�<i��<(�Tܯ�=����&�[�4!��\C�胃%��S���	&!��X+�`�w�,�@����v
!��	�T�fȡ�FJ��cw�M,!��W�D�����c�+�,�fHX�U�!��&� !���V�RXBc���A�!�Ӂv�$����1�T�(�fI,�!���<�@�9�F�,@�>����ݼqC!�� ������6Sv"1x��4����"O��5.�h
, w%Ц �*�jb"O<�ƨߏ1��CDT�{�<љ�"O�E���$=3.U�e�'S}`�9�"O\�Ӣ�t�M�����k���"Ob�q�e\�RT`�a/��Z˾8��"OvMB��F��^L��.�簴+"Oz��b��sV�p�T��n�l4a�"O�	񒇈aTm�ce�`NL��"O: ��z(��3��-��͡�"O��
��C�B �՛&��W�0�Sc"O~%`a�2<�f�i�j�:�R0P�"O�P�c!�
�(��5�Ҭp�2PA"O���g'7}�T�u�A%S��{�"OQ�f���"@µ��)u��@��"Ovm���H�8����ۊk��5�g"O�Ȼa�ȍX�^� d�3����#"O�pR�ݐhA2�f�C�����5"O�գ7I.��s�e�o��C"O~�����C3&��46te~ ��"O�xSf�V�&��I:�iG@��T"O4@�&Ԧ1JDt*�h�@��It"Oj�0�	��E�!���TIvF(p"O�\K���5L�T�_�m`�Y"OZhӅ��+_�t�A:1,b��"Ozٸg	K�H�,���ͳA�<)��"OVD�AI�/��A�D�I-_���"O���eI�.�y���Q�`��(X�"O�({G�ʱsv�0vj�)'W&d)Q"O���7�ؒ����"���F"O�!6B�]bۧe�+:!d48�"O ��)M
A�`3���4
� "O|�Ar�R�AL$ FE��L�V"OpARw�+~� q�q�<��	�U"OX+ �:]<v}�#���Q��I�"Om�Q�M��i��@A� �.�Hu"Op-���=��Q�&`("_>�a"O~Z�l��n/j�@�)A	Q�����"O)е+Lw�H@	Ժh����"O���ZGR;Wg�{��D��"O�M�u�H+
�|$�B�]�"T-��"O��*�_U ,;!��,}P`�"O��)$�� �d�	@&WwLH���"ODQ��"&� �G�h6XtA`"O�D�"m�� �)�c '� �"Oĸ��i�
G��%��O��8)�"O`��'�S� �>�{.��ڽ�"O,$�`E�&��8v��[���s�"O܍j���^�h�KrȌ@����1"O����ߤ��F�=�NH("OL �!$�"A��+`���Ҍq"O�|:s�6r�0ՙ��Z|H%#"Oؽ��aU�c�0�df]�p�đ+�"O�4Xd-S;6ʅ �gβP�����"O�L�`�W�Q����ݍ6۰9�A"O��� d����L�0>�8'"OP�x䎑7eA�)s&�T�)�,�3"Ota���2)*�"�/�3-�\�"O��P���9R�Բ䨄��01{�"Ov��QN�"������Y4!�R"O�!��R�)w�� ���+h��9G"O�5���W~�Ч�1|_t�0 "O&�c���Z���o�e�����"O�"t�Y�L���E�$Z��p�6"O� \��활s��]@Ac�=��1:"O佁�'�'���̲,P���"O܁�� ����T`]�_e|�:""O�y�%GO����@�6_X�a�"O�M���-z��
+O�a("Of��M(6M�D"�� �
�8�"OBD��Q06���R��O��E�p"O�8�a��K�>,khɬ1��-ص"OPIq��H���
D��p��K'"OLe�1�_�HN�hÆ�' ��q�s"O@��c��K6�l3!	?����"O�XP�Y��M�!�v{(�Q'"O�����Q�HAd�[�D�%ae"OԳV��>`�`PZ�*]�iG<	Q&"Oz}!��U�n��
𯉇Jnآ"Oq"f��{t�'H�=p9 qw"O���R�f��
{�`�r�ެ�!�DO�C,X�5]yv�	�RC�!�S2huxD�5u�1p@!��R�!�d��3<�y0O	3=L���"�`b!��JpH�v�Y+yk
�q��Q9'e!��	�4�)�/�@���`�O�`M!�$Ǧz����ڎj���#��[%!�U!�(�q���e�Ji�#86$!�Z��haؠ. �
��X� �X�??!�dWX�9���X?5� bcZ3+8!��G�dqt!r��U���x���K�&!�1䬰��G�Y���6��d!�d	a]�M���E�桱v߹#�!�Dʫ�%�@K�����D�>	�!�d�Q�zICfױe�^��B��x�!�d� O}�,�2���a�p}��D�2�!�DJ:G^��(Ԃ�`���@s����!�DH�3�\��\-j�|H�7�%F!�$Q]�^!@���A��C��S!�$�0���PqH�(Lq U�י_�!��݊<[�]�g�������bO�C!�dB3��h����A�hI����<�!�$Q�A\<`C�Pf¹B����!�dE4�Ҭ)b[6 dJ�h�fF�'y!�D�9�p�ihIph��+ׯ|�!�O9x>�Q#�۽<� 0ҳ*��!��k��h&�]�~�j�,O&]�!�D([��I� b�i���U�!�D�m�$��+���A;1��=k�!��Y��ȰD�T�q�ڵp���;�!�]Y<́!�mM�|��ٚ��Ο6!���:]��������N�[)!��9�"`1�ɛ4	�e�A��oE!�$Zr�<�3�������σuW!��T�t�v��ˆ	^��U��:%!�=��4��.|��T�d��3�!�$^7sm�����~�@y[f�؛d�!�6��1���D������ ��!��"V���8�h��}��O�t!�$!<�ȼ:sC�(�<!i@A�"�!�dX�q`|����x����� *�!�7Dl��v��2G�~�P'��z!�$�l@�X &Z�$�H���7>h!�BF�pJ'�ɥ	bDX���)8/!���#� ��ݽH��P"�Iƣ)!�D��B��Đ&U�[6��k��ȶ�!�*������c�2�9@�N�!�DV��F���C�"U��aF�ƕY�!�� &9���T�E/,uxP��E� -��"On�еhA� jְ	��1m�|!��"O�|�!�7���8&@�`��D"O:�G��>zO�̡1�{��P;�"O� ��]<7�:}B�@)|����"O0����L�(��Ȗ��i�~I�"O�y7��pDȬ��,������R"O^�"�U�}I���EL�>Z��Dx�"O0lB
u���L$u� ظ"O�({r���&��	s�� k���3�"O8��EN���)s�-3�H�E"O���2懠�f��蒢��I�W"O)���n91�G��,�0�G"O��"b �K>\���F��#��"O��q��
��Ի��Dc��%�G"O�Xpr�Ó��� "��q����"O�8b��$]�,�YZ�6H[Ċ�J�<1Ďܶ����䖡&(ЩC�f�M�<�s\�|8�#PH���T{B��H�<9����2����*�}�zQ�,�~�<ɔ�	
fr��)��DM:�R��}�<��/˷Xe�PG���pM����m�<A�G��ig�
N\2̀���f�<Y�C���Ɍ�j(h�뎆$�8����y�'	j��EF�|���K �Ti(]��'���{$�6�YGȇ(�����'��l���X�&~nH@r��-S� �	�'�A�dK8+2�!i�<�PA��'�̵!�b��1E�pa莮`����'H&-��bP�X�(�#J<�V�:�'*łB��_׆A��A v�$(�']�ᠠ��8J��B�V�����'��ܰG�+����dˋ9���k�'v!bKG
8�V�����8��E��'��Q�
�q!�<1@aب?�:���'� �FM�F��)�$Vh�0���9D��z�
�as�*��6X�蹂�8D�H���6]4���U>7�,:v�5LO��<�+D�Jxl�G@�e{p|��3D�����Ƞc��d+�AK4D�m1D�P8���4�B��eþ>".4�).D�0W��"K��/B�u�8�w&*D�XxFZ�b��q,^�:����­#D��¶��Z��4��%'�vdZ�$#D��#�U*Rm��1GY�,HP�3,<�hO��$'�� �D�aHq5�ό,\�C�I�#"^ ���A34��{Ck ��B䉣R��ҢM~��ʴm5��C��A\ ��U�=����_�}plB�a�:�k�#ݨ�\�K6��WC��Rk�i����I:�a��)P�C��$t5Bx*@iN�^��@C�J!#Q�C䉱[�T,���!^u(Г�`͒�rC�1U�D���Iڗ�$L�C��k0�B䉧~$��e��<��x�JՔo��B�	�n�����j�
d� ��nL�B�		�µ8��+s�e
6e�TB�5�L���#'�v��a��?pdB�I�B 4ŋ3��S����T��fL�C�ɺ[�����W�W)��րD'|�C�I�qB,y1@�ڴ	C���F��C��;X����fǟuP�� �_ `��C�	�UId�iRi��s������(8C�9z��{���L���5Ξ6yDC�)� T��Ƥ�#�ƙX��Oo�p�R�"O4�q���5� �--f�Q��"O���(�2ظUBB���dn")�"O~H�1�ϴl��h�0F^"k�\X4"O����$�+G�P�HE�݃-��|"�"Oe�ҏR�^�� �PCQ|� ��"O�s�a.�,��"�$�N9�u"O�컷#�S�~��èY�� "O�8���0ST���$Œ
���1"O���S�)	��8�#B�C�,�c1"Oj���LA&��[bȝ�bJ�y0"O���QeJ81L$BGG���%�u"O���W$��A*r/�)��h�"OZ9��"Ƃpz�	aaO	�}xF-Y�"Ox�q�(��XK'n3x(�Y�"O�4���U��u�@" 8���0"O�ah5��%}�u��1$|"O���B�A�L&�	$�H���XA�"O�	�W� 4bHt!�6�U:�Ą�U"O|â۳�.�a���){z&xh�"O�ibK�n�b�+q
Z�	r:ٲ�"ON�CT�s��(�r&ĸnU X�"O�1��̉pê�S�#�P���`�"Ov�sʓ�9"P�!�ȁ��P2"O����M%,J,��Ƈ�k:��"O�8!��HB8z4�ߤW.d-�y�ِC���p�	&�Lre��ybe��D#f!��CC�N�PEÁ�F�y�R)���r�qEt�!P�y�*կ��Q�aV6Q��i g���y� 	,����M�4�YUiՋ�y�B�	T7�5" k$E̖�H�d�=�y��73,<��-�Bи��V�_�y�Lҕ\�J�D(�	�,̸�$��yE��
�ra�u��K��)�T���y���Ztxw�D��I��ֹ�yb��^�lZJ�4�61"Ǌ� �y2��!�`QA\�}s���C�ޠ�y�'Z�7V*��c�L��q�d-�y�-�P��q���ǡ;���"g˵�y�ꎲ,�e
倗7O0��"����yR
�2=��ܫK�+f�[�@���y�̣
9,ؚtF��-kJ��f���y⦎�wg�Lз�	8(6`u����Py���/^h�$��F�vW6��W�<�D�*e�5*�#�.<�����Ê�<yw���%"Ü�nPX�� �
y�<9�� 'VP��CAۑ2�:���ll�<A�d��	�a3�eVBL'�n�<)b�_,}
-@�$�D��HdB�<i��F�G"ӣ�+/�y���z�<��LՋ-5*A��Z)a��`��N�<9�IB*.��m�RF�a.:�``�J�<a@n0�Ast��pk
����]n�<�T S⎀0@o�Z���hR�<yV� v��� �C<<Y��Q�<9��BK��EU#��v/ҵ��i�S�<���
_'p�1Z���!G��O�<I/M�d��c%���	���WH�<����4ze�	�1	X#�d�)"�F�<�@���4;H�g@E�Wl� �vh�@�<� �-T捠Q�U�eM��	"N��<��g�(o�*��dmY;�$ə ���<)J��X�ږm�(�(��'�<� �ij�G�7S�r���Oz�1E"O̽�A�W"W�.M��͔���"O��Å��~c>dK`F�k�n|�C"O�it���_�z4��S�t��uC�"O���G �2P��A%�f�Թ�"Oz ���&U��+2��3b��d%"O���%��SC\]2�WJ�T@�"Oi�G�:�\��+R�\ �"O�p�d�)E":<�a�ۄ|��U1"Oн��S�@�D���h��q��"O�P��Lm�R���3A4Mo"O��y0AT�D�Ъ�d�v1rAҲ"Ovɕk�5��4�c� T �]��"O�5�Q��.�B��ǉ�9fܑ�"O�a�c� V��ᆟ4p��0�"Oڈ0)R�F��$K��R)Or�y�"O��s�g��@�x�#:�¼
!"OHh��Y9S q;U��|���Q�"O\�F�,I��Pp�4*��U��"O�]��M_0���¶�Y'?�^@:�"O�4�bMN? ���uH�}�D�q7"Ozx�E���Rh�"'�������"O�a�'��
I�PR(
 p��i��"O�`2�0_1>��fF]#[&��ZV"O8�*�$�J�t"e�P��פ!!��d�Ɂ5l($��[*;C���"O�� ")աt�����/������"O�`aF����#g$U�g�B���"O��d�0(ʀ��q�� "w"O�а���.�zYc�M=+�҈҅"O�$Xge@��$ɑ��ֳ9�8E	�"OZI�OM+�!8���`o�9P"O詹u��=�4虐�O�,�p�9D"O�B��	�Ht��C6Ҫހ��"Oj<"R��*�l�b��K2�hr�"Oإ`�"H�4U�}�Q��11 ���c"OT��gŃ�y�2^�x��@S"OL��0��8$��B��Ӏ���z�"O���$�!��ʠ��]�ݣ�"O���P7Or4u�&�NJ ��"O�pS���=��ȣe�	\�Hhw"O������Kv6��#�K'!V� �"O\n.&���A�lr�N@@"O���5�ҘK��\�R��`�vAY�"O�C�L��j���:b"ON��h� Z�|��D�����"O�����
 ��L/:���G"Oz� �$X( �Ƞ{C)%`�X���"OX�A���<F���$��9!z�홳"Ovl� j�xΔ�@{T��H�"Oι*�k�O��c�[9/�� ��"OF��a"?GH<���Ä�8��"O0���\{�<�2ޱ6w��c�"OQ9�	K/��1�$��Hd��"O`��@���>��4�d��Ym
��"O>Q�R" �N���B���Gm ,��"Oza� M��;�RC	R3m�|��5"O�� �g�`�*�"LҊ��V"O"� w��7Z���J(�����aB"O�pTX!_S�DFޓF$Se"ON-�U � ���Q�d�7O���a�"O���v����D�CB�C �"OP ��J5}?���N�,!�X|��"O�9a�e�:  �a�K'?瞬9G"O�  ��U���5iO�v�.H��"O<�D	z�����ԹE�.0+�"O��h7B�#P���q&�::�P�"Od\j�*�5>̘�c(�1�I9�"O<[�\�}G(Q*"����R�[�"O.�)�xg�};��
3���h�"O8x!��Xj҅����?Y}��# "OHp��I	E`��KRd](r�tx&"O���Ν�c��C�P�y"O| 2$F�8�"�*6�R�!�B�x"O��"D�I�pJ2(@D㑄�XH`"OZ�ۑ��G���)�AW�B ��"O����'��~up����a�j��a"O�D�F��)�X�ǧt�ba�V"O@!Q#C].I$R���nEE�
��"O�I���!���4�p��"OZ�TE���j� v\h�xU�R"Ozzf��|\k5��w��*�"OQ�"��(��@-P��`A�"O@4�SnD���!33��(�Z�jE"OPTQe$�WdP��K���rhQ`"O�xP��
�+���d���d0�l�7"OB����<:X<��M>c�"O�Ya�k��� �-�+�L��"O�3��̢Z� ��/��8�"OF ��I3b���)g��k�4K�"Ox9��(��}J����MH����"O��7�̠$ӒYB0�,TM�4xS"O$�A ��(c_�5(呿
�t�[�"O�D8"�O�tc�xR���s���3"O�RAN10�q��ɞSzz�h�"O���+#��\���X&s�Lr4"O�������S$]CLٟ7�@!q�"O��2�(T�	 27��:@�Rđ�"OX��ta�e�$�4aP U���5"O�XA�BΑ:^��R�3��7�'D�`�O�N2�+�i�Z�\�2gE$D�� UTQ*�a�+��e�)��� D�i��ݹ!�!q���R�>D�pv�:#HR	�7H�E�q#$>D� �C�üZ��r@E̥a�f ���<D����8V/"A�� o�:8��/D�\A�@_9VXQ��Ʊ&	(<B�f,D�������b��U& h�Ĵ���6D�pBGF�)*~�<S��*ʞ`p-"D��"h�k�Iƌ��'7J��,>D�X����[��9� Ԧ�*�Cqe(D�ܒу�X��'J�.`�L����$D��C!�:�<DCn��[R��a#D�,����"��]�'��/ �>1CE$D��0 M�
̩ҥG�M����2�"D�tۂ(\�.y�x��	���# D�t �lLXm��6Á�Z~�Ca3D���r(�+�P���Ӯ`T%p��/D�`�A�H�}�:�2��T�
�jT�+D�H�Ӈ�4jS��R���7$
E�cF)D�(&K�K{�`�q�!"�u��9D�t�a̟�%�l�)Ţ۸S)x�ѷ�2D�p"��A�\Jݲr	w���iġ&D�t9R�<C�
5�4h��d=�͈��"D�X��f],DXV0���G��|}C�f D��R��B�&q�� ��P!��h�S�=D�@��JӾI�JDP�A�-���b;D���͌�1�U:�L�?�Es�>D�� �TJ��>="���aJ�{Q"O�hc���'��IÜ�d�(A"O �sk�f�0�!Q�L�Lhs"O^�X�B�	��������*}�<�F"O��(&j̉9� ����7���c"O�K���=�>���Ο!F�,�S�"O�X�e-2��H[ƱCl��"O�Pg-ߞ��n�(c��K�"O8=�&Nн���X��-J��h�"Ol\���
�����m�2I*����"O&�9Ck�?g�%KWF�-�<B�"O4dx1��<cHεJ����I'ޘ;"O,x�6cdq����,Z9̈Hu"O�uY�KQ ����eE=U*�K�"O�$�"��J�j�2�,oqX\I�"O,�H���8��ci�T�V�j�<9�.��D|��	q�@��Dr�<9�o�6C���(��, Ժ���O�F�<a�`� ~��B(Yۂ1�Rl�<�Ņ� ]@̡Q�Q�\$�����]�<!�a
t����h�Fu����J'D�h����4W���Yv �2,=���&&D�,@tcP�#��<��J҃+����$D��s�̍�q�4��m�~�Yr�<D��S�eT']�ش��ڭ4^E���.D�pI��J	w��iVl�Z2���-D�T��K�p�l�s!Y�w& 1s��+D�pSe,�u`t��N��yp�(D� z E�����
�v�椪G@4D��i��a��-IM	8J%x���0D��`����uڀ�����!�x��"D�Dʀl� f12m��K	�9�n"D�P��G]�
԰e��
I�wT�U �."D�� E�Jr)�u��O��(�d>D�
u��;_X�!"��v��$�d ;D�ԢTj�k@ �X���O
��&!7D�p��)��k�Vt���i���W�4D���WLP	@��RdȢY4.��N8D�rE#O1	��Уm�J��W
5D�� L�6��b`���$�B|��3D�8y��F"M�\P�ț!WH"�ʳ-D�Ls�#[34�(!��D�$&� pM D��X���
/dp�25�A8ܪ$; �>D� �&��;:BM�Q�_T^�ZSd"D��"��L��!�e݃N
�h���!D�,��@�)��$Q��=tZja�%D����JMx�
��A?9e�yjp�.D�T�"-O��Y��<��1Q�>D��	� ��&y� F^	(H��0D�0�ċ߂J�x��FLֱoD���)-D������VZ�Ih�f�2}�*@�gH7D�x��fH�_�a#ǣq���c�*D��r�EۄF�<33�E�/s��*$K%D�x���(�r�S�.C;c��cè"D�{��=|�Y%��>p�( D��!�Lq�(qCfά@ 4�c =D��#�f�B��}��� 	8 ��%D��J6�Ԇ�(D�di��-��=��O"D�`��g��[m�	��ߣ[%ɠ?D������9cn�[1�]�c�&�[��<D�l0�� �,Y�ܘS-�U"1�9D��PFi^qda+ɖ%0���hP6D�DB�'��K5R�2 A�NO��*��9D��z�E��'~*I%�K~Vl]�t7D�� ���$�ԛe��ab�DU%"���p "OƝQ�%�2_���"c'~x�"OX4J0�_,k�h����?psژ��"O�$��*[|��S���.i�`��"O����B�(&! q�'Cg>��"O�x�EEm:1�2o�
Z?��9"O�����o�P1��M2���"O�Y��I��w� �`1��&�,��"O�;���.~�Z��!D�5V�Z�"O4�a��Ҭ<p��BʊF��1 3"O접���{���!̓�b�T�:5"Oxm��m��<�gM*�x��"OVm�����"2���uL�R-�9+t"O�Aҁȑ|�l�+O�I"r%�t"O��@��f�>���J��${��ص"O��q��F"��ǉ��v��1"Od�"�*L3;�j�[�,3f.�S�"O�dR�� H�>$��%�*a�,P5"O`}�D��o��ԡr�X'���&"O��6BM�djǆ�>��*S"OXYط��&)�9F��]��"O�gC��N`�ZEoč{�,��"O>x���U�9������ ���2"O�$�EgI�[�L۱�\�C���`�"Ot�PB�?������IC�C�"O��H+3\�p3� .6��J�"O e[R螯K�pyb�Ł1b�T"O���l\�"+b�fE�P��e"O���D��6�1w�P4f�T|(�"O"Xrv�˂Xs���)0D눼H"O�,*��-	�z�"�3��́�"O����I]b��2�NM{&���"O��@JCvOx���'>^�j�"O�tQR�Ť}-��˖�R^�X%L`�<A�c� _"�E�`H	\?�SC�E�<!$��!c*���ViM�@���3B�ND�<�AT
=��˥, [Ӡ؀f#�B�<A �2D�����D�9s���1��~�<9��ƅ���2�MN2t�Z����a�<9�-�l��i�#���Q���Z�<�ã͍6|�  WB�i�m��/ET�<�$�R|�`�	�A����E�AQ�<��i^�����RY֨9R'�f�<��K
� a���G	V� TM|�<�C�H!����"�\��!p�Ot�<��C]{]1#�(R:6��-{u��m�<���Px��
@�;fɂ�_�<	�f��\Z��q��+�j����Y�<�R:7�d�xhʍ[\(��aKIR�<�DdD+���	%�Y�v_:YS�K�<� �%~e�}�HM�h-{D�D�<9gܢ8�6Q��F
�'��	cf��}�<�Dbԏ)�i�i^3�LpG�x�<)��M�h�t���%挑`��J�<a!�N;=����]�$8p��J�<a�野:X8up�/�\*����"�]�<��(7)j"\"C�,>Tz���\�<9q�C�?�����\"��) �O�<i!�Z�;��� _�����
C�<�w�t�z\PA��VC^Ua��j�<y�aD�{&l��*�C�X���q�<ٳ��#r�U��f܎F����d�<�Ef�	7�${�l��=��,ǩd�<�W�K$[=ޘ����o�����KQZ�<� 8	2� �D�8��O�T/���B"O���*ѩJ�.ds`އo8F9��"O<| GBܖ�݉b��E; ��#"O|�ؕ����P�!OG��Zq��"O�%3�*-~;:�+&-ǘ=��`��"O��I��S���c�L᲌�q�B�<�H�:~�1��H��%C�~�<��m�K.��"�
A'<�()@c�O�<��O�0kd�`�^$s��gH�<9����7CFx#o�&n�8p'�k�<y��AT:9�������XTČe�<����ms��BW��_.�p��c�<�a�C�9K�/ѕ?X,����+T����O-H����S����*(D�l{�c�^z0I��L�h���P5�3D���gU�w?��A6�3
��y���.D�0З�ӷ4"�;�h�(N�r)T:D����*��_\��ajڡ|]��f�:D����N�g��d�f��1�Ԭ���8D�|
Bo��N
��h���U;��9D#D��3D�+�V��PKX	3����w%#D�8	�M�	>�^�9�h��f�y'!D���d\�<=��)�"�)7}�?D�0� �F��81d
9G��h��<D�`��a��pd��3D��~�Ԙ:��4D��)��ۋc���c���dq�0)��.D��Ȥ$�0R�B�B��']��P�&�*D�Hi��Ȃ}0v=�B*��A���e'D��t%1�	y�B\:x����@%D�Ȁ�Q?������ى@z���##D�$	�.�rO�C�,s^�9�F!D�`!� �A�A����^�d�N D�La���/+h9����ND�5�=D�<Ip(0 �^؂`c�D��T�5g)D�PhVfl�ɂ��R�*���K��'D��*�"ƓjN�\�%��[��ԋ��&D���%�.*�8|a�m���2ӏ#D���ƭ��=`���,:�p(Bk�@�<�#锱k�Z`��%YZ)��i�w�<1�*פ�c��P.�@�;��@u�<����p|��ë)�#E��t�<1�F�]P@9��;}�͢vn�I�<i� A�^`�1�Ԝ|��ґ`F�<i�f�+g��.:���SiW�<��������N% $mB��R�<1�+	�>@���Ҥ8�쒅-�O�<�R��(%� �`�$3b��rD�SL�<��΍�&�`�Ҟ$0�\��^I�<1Ӭ��,"���A�$�|c�E�<����"�}C�K��
z\���MB�<Q�̽�����	�-J��<���IA�<Av��\�4%s��T�4&`���!�|�<���~�D�;�CW�[.��آ��d�<)Bɂ�R�\�!��(5!���E��^�<YI9]�p�[gG�/X�JjA�]�<)匂~�4=3�i��;w�<�3�Z�<���ў@��q��-��/$��{@F�S�<	���8f| G�U9uΆ�A� P�<9��K<�\Yx"�Y�}�čS�MPJ�<!�C� ��0�fa���>�d%�G�<�F�2X9��@�oضW�D�I��D�<a$'�*���ᑁ�.�p�7�H@�<q�O �8����퐭8�� Y'O~�<1�hS=j]j�:�ի˸-+0A�e�<� �Pᬇ�hB�!��9��s"O��(�<]漛��^2a��)��"OLR��?��1g�WL�~�j�"OR%��C���xam%S��81"O������+@����ިC.NEz�"O�@�G>��Lӕj�o�<s�"O�x���;7�f��l�"x�"O2����B7h[V 
l�9��Ĉ�"OZdSs�!�f-0��۷)�a:�"O�9�4�R�<��iDD��!� �"Od���eH�RP��z�C��P�0�"O�uA�)
�2�X
��  ��Yj�"Oz�#!-&ܰ:�Q� ���"O��R�U|����&¶#��2"O��C$e��.�����Z��yu"Od���Ċ�,�j  �ՍW���7"O�����i��[ �~�8%�"O����)D4KE~P��F�3��""OpQ�e�B�dBY{�E�R�:�)�"Ohaـ�S0l��a���r�@l�q"O2l�S��;.�&�(5j/"w&]j�"Od��� E�.���ҋm�0(C"O.�'���*񧄃�f�hb"O8mر�M!��X�'H����"O p�#�[;��T��֕�&�x�"Ox5 2K&Q���P������"O��a���37�=�I�}Cn,��"O�p%��$YJqJ���P'��j�"OP�"e��0Tl���B* 20�"Ot�re�50[ޡ���J���"OD�jFl,Q�H@b��׷=۰D��"O������,�H�bD^)a�����"OpѠQn��sApP9��g�$A�"O��g�+`��W㈈b�̭�&"O��C �H )>��ꆣ�Q3b\��"Ot|�g	�c�Ma劀!���"O���t�
)��*���~]95"O�������qa��"RA�ƾ�"O���'-��0x���6��p%"Od��v�ى����&���ڕ"O.(���P�&:&�`7m_�l���`"O��I�P��8�+(pW�q"O~ ��&��hj�K�&=W����"O� yV�V�	��tJd� H�D��"OXP1�<�����Q>L� x)�"O�d�4G�W?�)a��V�I���ju"O,����8�!�c�ٛI���[$"O��(B��6%F�$S�GF�1�՘�"O�D; ��!@��0F�a<Y!7"O(��Ï�O �u@ ��a�%��"O�4��dݰ�h��C��J!@@�"O�ەK�;~���TcY�j~�1!"O�9�d�ly �{s�H+j��C"O�T���BU��в��QȅJ"O�-aT'F85p�Њ�H��T0�X�"Ot�T�H�B(�u��"+QF��"O~�c�"�N���D*P�L�w"Oe@��ټVG��xV�MO9�,�"O��9F윉��р�F��C�
 �"OQ��CbUr(IYi����M�R�<�'�ъ'3�aP#�1u=��	���H�<IV��*/u�륉L�j��+�C�E�<I�,L�'
b��0?�ѫT�~�<	%a�<0Q��BF�!�����*�z�<� �5
IN(��\:��[�9|lИ�"O�XƯ�fd���a	t�xf"O�d0�MV�>���w�@�?yB��b"OH0	`�(�d|�p��h�d�"O��&+Ǔ7�UKEEB= ��L�"O�a��M�sji�F��P8�@"Ox`���<<PBâZ+V+�D�B"O�Ë�8P�;���e^�q"OZ���Mçi/LI��.Nr��"Ot�8���6B����D7!^<�5"O����*M�f"�mq�CVZUz��"O���cG@}'p��B�aQz(�"O �	��0�FII���׾I�"Oz��Ɔ�`�d٨�"�'#�]�`"O*1ȅL?t
]2�"YH5"O�����:4���nK>
�R"O���$��p�%k�p��Yw"O�dJ6Ά�	Ĕ\��D�e�0�"O, �壑�SK�(�R����!(�"O�@٤�.o��
a�N�6��퉶"O�hhF$	�l�R�c3j�4�Ԝ��"OV!(�A��w�ԋ��G����P�"O����ߙX����kNL��P E"O�t�GG5'?u@`(W1q�^��"OLը҄V�,z��տ9����"O$����"0e�7K�Z�.$!�D�4����]�e�te{��cQ!�$�d�8)��O��������� �� $� �G��{�g�6f��=�ȓs�2H�5OOe[�8���J2K��ȓE^��s�b�!�&"�e]<�ȓIajpH�b@0k

Q��.Y�'�$݅�h��l�c`ʇ`a��k�3�Z<�ȓ-����	�DN�5`w�� �P��ȓ
2Iy��P\�D��B�JΤ\�ȓI��A�,' U�a���FV�цȓt�HeZ4Il�d���nKG+�8�ȓ W���"�5$R������ ���,[�	g��.�J1��N����#l����B!G�x�GC
lԅ�$M<A�E���z����M�^ڐD��&,�B"f��	&�QX1�C0u�8�ȓA���!%��'K��1❒5�y��u�|�I��+|1S�'�$4.,���X��Z֊�/g���J��"	�ą�]��%�0.�-R%�|}4��ȓ�������	.$������ȓu$l�$�;=���1c�53����z�'�F
]��ِ%�5Y�0u�ȓ��[OVb��t�u@�2E�����*�5�Y�qeV� ���#��ȇ�_gl�EÊ/�n�Cpc��f쾱��-us��S��"�8���R�8��ȓ��J��-+)1���T���ȓJ�|Mh$,�_�RlH��T_4u�ȓf|�ܑQ��,�l�yS	B0T l�ȓi��0���dV��&���l��̈́ȓj3���!b��$~ɠrc�
!�����a�֡p��Z� � JN+O�I��!��QB���)����CH#~K ��17�-x1.��hwb��\Nt-�ȓ4�
�R ��Nk��;�Z�JX,�ȓntX	���'����Ac�,Y�A�ȓx�����<!��:��ۦ;�bu��S�? p���L��]9r����M��0�"O~�q��ЖP��=0�A���ԑ�*O��at�9���ĞCYP��
�'>�GDE	(ܚݻ��þ6t}(�'�\1:��єw��P���'�Y;
�'�vQs��un���Tx�4<�����a˿6��R��͂j�H܄ȓhC0̋Q�W�2& �#�
{�<��ȓ42.���`��u(҈��o�:
>N���*� B���?�EKG��I~X�ȓt�C6��6r´�c�˪�0��sJ���7�D�[� u�E�%5�T�ȓ�R�R.q���E�B�W#��ȓA���1qh�2.ت��%	�qZ$�ȓN�	�(U�O���Gٞo�X�ȓ,��a0���iPB��
�H{�ȓi2�@���ɬ=K�D8g���X �(��4q�A��匁Cb�Q�m��[�̄ȓ=��pi!)��R@(����+��%�����a�ě=}4�Qf`[ ����m�����#W�Pg��`a�,"���v5�paN]�^f�\j'�X�(�y�ȓ�֬��m�=/�����9�V��ȓy�����LsƎH3'�х�.�̴��.2x�b(�\Ņ�D�0]��eN���bg�5�책�'��A�6N�,>�}�7n��5JE�ȓe?�� a)��w`�D�wJ�~aB)��We\���i�SL8��ċ)dv���E�lJăO�\SH8b�C�n���ȓ7�6�
�CȘP�R��C�\�!��l�ȓD�@�V)X�7(���3ɢ��ȓX1X5 �L�:��%�� G�:D��ȓ���cgNޕA�
�Qp������9��QgY��fy�åd�"��ȓ1ᔌ�G
�`�4)�*d��ц�X�h�C�:1'J���ўHY���T������%A��!�3�W�{/|��ȓ,�x,�e�3v�h�`��=�l���yt��z�A�G�]�tń�E�<ЙU1嬬r�J�� Z�q�ȓ���%l��l���,k=�4��%�x7��V���K�@SN��ȓ	a�ɕ�a_։أ!��?gl��G�`騁V;x�FpбO&X����ȓ`�@�z�È�kd�`�&U(r��Ʌ�T�Bl!&�pv�X�PG�;O]�)�ȓ?d]���)|�a�Fg���N�ȓ<¤(@+�"p)9��/�ȓ<Dv��&������@�G���ȓ
0ĉ���:yjl� %��	e^���u���S C2l$����5��݆ȓ ��{�M4fT �{���	$�:�����݁$焳k��X�cG�5�̇�]���o�nA�����Y��8���hK^��A�҆zjnYiu��l0A��]
b���+A����P'+RR$��Ldb���:5��2 ��<���ȓ;NF0)�B�zQ*�5g�Vl�ȓ/�2���`�z����/��X�ȓ?���2��:�t�CZY��0��,Ј�Cr�B�l� p��*�A�4�ȓ�xH�C��i�Ab�O:t��ȓ*P�
W�e#�(�I�7v*,��S�? ��KbV�uj���"QVOj��"Oڡ�&Е�h؅�^!9Ox4f"O} ��I�V�XA��2�:ّ*OR%�Ӣ�'�ʀ����=o���'bd=F�ɤ!�dp
�3����'���(���u���"R�
b� ��'3 ��G �@�¨1ũ�Y@��'d���	,�l�W���}C�J�'�t�ċU厨@�@��rmrQ��'3�9c�#Õ|5���D���h��'�F$��k��X?r�+��	�1�'-�)R�疶o�9�Ʉ�h�x���'�X4�Ʌ �Q(q!�0\����'��q���W�I�S�^�W�
���'\a b�)���bI5���'�$C%S:ZT �x%��yZ�'��)�SN��g���E�?rh8�	
�'L8��V�K �ొ�k_�\�	�'�y���_.6�R�C���mǄ���'n�t{DiV�Og�m�0G:_���	�'>���.��h��P!��~X��'���HC�4�J4`�ދQ�:t��'��b��Z��}��̀!B����'Ҩ��S�]:I�`���5��	
�'��xGJ2=�l�*�y���	�'���c�j/8S4�"��8�2�	�'kaB�b��2��a�@�����'g����g���Td&^<�X!x�'��q��B�X_8 ��S�|d�s�'��)�cU�BYR@j��^�n��'*���"�`�~U�#��V��8��';$0�����4��@��7���'�0���3p��@�U12'� 
�'�8 �Ɛy;9˲�' �8(9�{�F?\OX�QjȒaB�D�G�Z!t��t"O.QB��S�G#� �w���~�Dز"O����Q�r��u2r��'G��"s�'8:��=�e�R=W;����߻ ���c@K�d�<���I Π42��A�g��U��Lj̓�hO1��5A�(��u{�Ѣ�l�9V��t"O]���-]�6a�U��54�Y:A"O =ٶ�]|Zp�Ca�o� Xc%"OxxS0&['~]2\IW
.8E�=ѳX���	7W�&��V+T2�6�Ѧ��:ekJ���K}B�ԍH�F��!�N.�<�����y�'�a�L�ɴ��2L� ��2(���y�Y!}�
L���8y�hI�B<˰?�R��OFI�q䕣k_2��V�%9P�m��IO>YXǮ��[����1�X=�; �,򓧨� ��QEV�m6Y2�3����"O�0���-+"� ��4]�ܣ'\�PE{��I��X���SO�$ی�P��W�n�!�d��l�^5H�A�^Ͷ��t�܀}M����
Ǔ��V�v!F@�b��>����a-��a�w� hA�9<��#%Y7"����$D���shL�V�8�ōۺ	����� �!�?�!JO/S`���FN�KX��Am>D��Pm\�9�|�X@+0�B�4i;�Hb�4�l1k�L3r���0�A�f��$�O,��$@J���C����&x
���8D�!��U�~������S]
��� h�!�$��m@td�B��-FZıAP)�*v��Iu�s���I�3>@���.RKyZ�yt(���!�dh�@y���+onm*Rf�1VL�����s�� r=:�$��g�N��U��%HM�@��'��O�49�nW TyJt��H�A�0P�0��ɁX���ˣ�ɍN6nT��ᆗk�@B�I�u�nU ���<,e	��)�B�	�c����J �z�ګA@���*��ФC��vn\��F�:i���B!/O#=��W�-�����i5CZʕZ� �W�<A��G" �0T*w��$_�-���Xl�	W�'���<a��Θ~�Rd�,}ؼ���L@�<���4 �5�ք����5;��'��s��S��[N�q锡��7Q��87�94�h3���;�� V�J�LM�d9M�/�?��J&�S�O/�T��쁢~Uѩ�ˇ*L�M�ϓ��O�r�䗹8t�Q���C��XH�x��'���p_���Q�2�W�qY�q�'���x��0r
"0�Fh�p��	�'����A@)!��R`h��b����'/D�˓�P�9�L$hB��`Ȋ���'\�1o���x%(ӆ]w<QC�'�TrG���NB�tB%�[�(QX���*�S�tBEB��1>X��aj��y��Z!b)xX����<x�!ّ@�ў"~ΓHJ:�h���2+����6�0l�@�ȓ6���wKC2E��a��3zL̓ta"�ڨ_������#j��82#���y�F�H6j$;7��=b�x!Cg�����[���Oy�`i�E#id��
#���*nV�ˌ��9�w��DӶl
�o��E�L7QkN��=yۓ?2j�;��(-�M�A3u4��' x#=����^�tw@��c��^I(u�rG�R�!�U�| ��J
XZP@���-|!�	����#,�֤ST��
!�dY�J}8�F�?K�6��$#N�u!�$֐WL,9�2�H�,)L R�z�x��'e�O��+5�z��JaX�J�]�C"O���!C8�F�y����mH��c�>��;��|ʅc	Ϧ	��ӌA�w"Tb���%O��|�h��qO 9 b��8��p���\�X�H����O�������z@�!��l��`z�M���ݥ/I!򄅭a�����J�0qt4�qʟUDXT�'�ҒO?��%m��3�a�?��-Kw�[12 �ɞ��'��>����0U����f��;���UI�<a� ,z�u�#�뗩S�V����'�ў"|��V� �H��8WT�0� �.!�d�O4@�$l�rb���W�ِyQ�"O*TS��\�!�<%j�b�'l��Z�
O.6��n�9q�&?��2�n,�!��.q�`�AlC�,(�ˈ�e�!�GkL�	�&R�X���E��:���Nx�� ���n�#�����K��3D�(���	h�*)9��'wX�A!�-�O��d�yQl P�@h
e�	������K'��s�޺/��Q�r`�c�NF~��'Ԑ����U�8y0�Ц��P���OY�	@���O����C K=�F�� ��T��'Y�9
�-n�jm�������i�'�H�YclZ�T��ʀ-[��ܠ��'A����U�o���SgV e�`0��`_h����'�z
mB�kD���BO4P��Ó�hOJh�䈬e�L-��Ăk[|�"O�(�n�n ՓF� hK\��!"O��y!l��qw-;�B��_C�4�|�"8�Sܧ�6�0o�?

���0!��)�R��ȓ����P��e;&+�4�,��>Q�S�? �E��N��6 ��5n��_-�t�W"O\-�``��2�R�+��R�q���"O�����J�%���Z�\�m��F"Oֽ[��\wZm�#�=~��T"OjL��F��	�Ь�RH8ۅZ�3g!�N���t���͹G��iQw�][!�)d�ta�nY1|6^Y�1@Re!��%3j�}C��7@�82���
L+!�D����@3����XT�  �n�!��;)�4��iR1K��!ΨZ�!�d^���І�Z+���C���!����-�L�$I�#��`��C�	9Q�Hx��wu	6�\�6MvC��-�6�z"�6]��T��`܇D��C�ɝk�K�fH%La�����Q�����ZO2��Sŝ7J�yP���q�!�$�t����e���>ՙ!l%�!�ִ%@F����g�0,�e+�V�!��"9�q��N�>e�RЈ��FE!�R[R�S��ь"���㦏�%-�!���(A&ș��X�Rʒ�eqI�'p� �λb�be��d\�:�t�h�'�|���j�%���p�)�.Cl��'�jQ��F˙h�d�Ȋ+p��h��'q�8�w�M�E�T	HTO�e��Xc�'�j���,�p���_�\��H��'���$�@"(f�H!`��V;� �'�Ȅ�Fc�r2��A�Vs����'����uǃ)<���B7AC W�l���'�\��ԣ�5�@�o�\~���'u��8GjÖkH	:��AZ���P�'x
�D�?H~�{V*VNX�
�'[J4��E3X�MqEG��G�b	�'<��"��tu������O����'�|��G��`��[э�=H!XX��'���{6���`hP��A�a��	�' ���E��8�T�X0�0Zz���'㲐ЩL5h�qbF�SJ s�'Y��0��0���QnϠEۀ-��'��ܨ�%�b�n�9�,����8�'y�1���ȓ?�pd�R ܸ ͸=0�'E�qـa��_p��dΒ&&A��'"����1FP<j���~*6)��'tX��=4�f1��u}�E��'�}r�H��38N�s
������'�`B��'���UF7OҲ}��'�h��J߀�H<QUG x�[�'��=���ǎ<�0�q��_�o�v�1�'
L�xvCQ6�rQ@d�D�nB �)�'�ⱳ�E�n�~1k^�`y����y�<��#�����G-^�x[��1��\�<	�`��>\1IV�_�>�v��PQ�<)�̀2���� )S��ț�M�P�<�Skџ���䆘��Q;# �v�<)�Q��z��I�5ju<���\�<a�E	0�z�7b�.bL9Ig�]�<Aw��#}ز�Pl�b��8I��U�<�%��XV&m��Έ�"���8��|�<��/?9����#�`8�)�|�<����\F�����{U���OMy�<YSE	)|ED����CgV<+�(p�<y��ޣ{k� �3t�ˤ��k�<ɀ�>`��XPQ��0u�Q�	A�<�u�A�;x�����\�|�1+�%Nz�<� j�@�K�(�j���,����Z�"O&<��J�br�!c��/H�����"O.�x磇�Y
��H���%O���7"O�Z��Y�9#��I�*Ih���S�"OT$�L )���L��w&r Z�"O�(��X	���i#��N& (w"O"д��,w�����+"�}  "O&���̲>�b�A���r�*�:�"O2��*ϡ*TtKC@C�d�Q`"On\0�G]M����#��a�|z�"O��B�`Lt�i��+�&m��"OZ,x�&�7k���y�
ʻĬ�KC"O����Q0rze���Sl��JG"O�a���1A2��c4�� ���;P"Od� e��<~XՋd�R1Q�����"O1%�-%��8��Xx�P0"O`�3�ܵb�@��KT�|j����"OL�U$	Z}�'$�0h��S"O��%k�#;��bw�� �:��"O�䪣�\�y��	���vpt�V"O.����ot�$�w�β$1���"O��)��aĦ=#���*PQ�g"Of!��˸X�h-����6��3�"Op���dOr:������a�f�Y�"O��D��	l���:�C�ݴ�ad"O�y�*�	$�x���q0�"O�13��=r2:�5
� ,.���'�d=�)�2Fu�2	�f�ء�TA�5".�"�'ZD���_μ0���
%�����'�Դ�Ư
&rp�LǮ0��	�'(aC��M>Z$�$;��ϱA��a��-{>�'��� �� �2����!l��*,*���(/D��`# K�3>��e�
(o ͡��7D��b0�W8r�=R�$Z�fE���,l����E��;Zq�Q�S'r�����U��2�ȓJ^��%�6c�6��P�I>Bw�p�zvd�<�e�		6����MO�6�c�@Q�{z����>Y�k�jظD{#���~:i`R+�Q?��4���'��a�gP802�A���Z�4�	�')(�!	;Vٻ�ǎ�?Z��'�,ucG�S�v���ʁCЂd�Y�{��)��B���	X5_~H`��6M�'��|R���q]�l�4W58��=�`�Ţ�y�B^�JȚ,�Ǡ�.�����K���y�Ι�h3����#]7 ������[��yR�]0\��,Ih�9�ن��Ok�ӝ%��ũ�*%}	H��D���C�	;�|�r#+P�Fv�[fL,~����y�'�ӧ��{�$�U�N>QC�,��B��!Q���y���R�����i�p$�b���ē�a|�Z�VC*�zt�7qЅhVM����<)����� /ā�d��"Z��E�H8t!�dK�C�Bh��M���z=z��=d!�wk���W�W�\U���	PV!��Л~�a��Wsi2\��ې@K!�D�8<~]�(]�'�t����;<!���N��'��s��7�|1!�d	:#����eƇ�8Ơ��$0!�G:�.���7�8bgU�hqO����ԃ� ��C�/ �����5n�!�dA���A23��3�9�gdۮ�!� ���MT%h�4�@0#�n�4D�ıi�~0���?|q8嘷���c�N��
�'C��1�ȜC`�Y��/ξ�9��� ^����_�0�Y ��W** �"O*�ɒ��4=�`���:>�1�"On�����(���p ��6�2�"O��ңQ/i�jݑ��9oD��"O�R��M����P�L'-
e�':���S�I����J3%�$qwGA�	�,���L ��G�<L���
Y	
�pԇ�2��� ��[����̔BT�p�ȓ+�	�)ĞP�P�S�S>th�bL(��x���K�T���X�صigB$LO6�4���B�ه�ޙ W�.e�B�I�mE�|K�!7U�}��MO	#��b�PD{��d@��,�4 ڿfS������(�y�jV�� ��צm3X��%\��=a�y�پW$.	�bٍ^5���J�y�n^�<�X8�'ȩ~��1A%��?!H��n~x��PD�	��������1��Y��%$��hO�E�8� �CH*Zk M���<Y�bC�	 `�.С��=D���G`ѓ&� O����'D�'���M��x��-}ZA8�É��yr�ɑ}n�	��e�u#^� ��y��<:��:qJ<m�ܡӲ���y�$�&(�ܩÀ� g�<�Yr�V$�y��W�T�Yk2��!$޽A�HX���'���`�O�����*R��E�Ƽ(9�'VI��dL�F�0Y�U/ 4i
�'Z�����@����'	�w��`��'=�S�"J"@���{���1h
��	�'��� (�&<N�ʤ�D�_*��	��yR#�(S�} ��I�J\\!�&Q�U5t�<y���O����BİJ��C`�Қ"�r%B�"O����"Z"����$�d�R!�"O|pҵ�TPMa�o 14�T���'��O�'�%bq�� 0N�4�rV�'�!�$�!p&:� ʊ4�80�%��L!�ʥ*�*٪��M����3�A�]�!�ůE~��rE�  ���e��DDBR��G{��ԍ�}�B+0BX4@�
1�G��y��tC�� ��X�$M5��B�y�+V,�m�A@;(��A��ϧ���,�Ş�yrM[�����������vͨ�yҢվr~�����ɪIJ��&�$�HOv�=�O��7bȵUb䫐	Зh���b�'�@=�s	�q��]�!�!O�V2,Oz�=E�$%�� ���A��G�R�zS��O�y�-�x/��)ǆ]`��І��y�Ȓ ��р��')&���3�ē�~�7O��4�O�<dI3c�/Ҍ��@�E{Qf�A�H�x��_^��3gO�P�l�h��yB��p� ��ꆠC�d��
�y�+L�E��%�b"�@�ȱ�Љe�`G{���i��\A��K~� �CLȖ4^B�:�'����5H~���,ƿ|�J���'�4؁4f�-������&&�P��Oz�=�}۴N��wj�b�p��0�����i��w�9��ؽZ�H�U�P��ޱH�y"�8lO֌@����M:���z����(�O�X�47'�����X�h@�!xP״2~T!Dx��)���ʳtɬ� �a��.݈�Z@�uX�PFy�2�Q!'-w�f�Z�:�y�ȍ�	��mc��J:rº	��nٗ���ē!�@�>��ODځ1���s܀i��JSH+B���'G"L�7/�>[���t�S���y��d5�S���5*� -h���bL�Q���3��>��O� 0�Z��&�у�H��Z$ޤs�"O�<�6�P�.�r�n3���"O�͊���'���S�͗�hl`�6"O�1�&�V�0DrF�تH[�p�R��E{���B>n�ʑ򒂅/#5 �-_ �Q�	�'��b�]Ί�1Al�6%G,M�	�'��yk�lĞr�RY毘�!�4�[	�o�(c��Z§H.�
��Ė�O5yf�!D�`sዒ�%�L��Ӌ>�"�`�i,D��;D�5`�hB%�(w�i1�+D�0�d*,Ez@�u ��yh
m�<������߉;. ́0B�
�"Ԅ�H�ܸ�,'4�`����K�t�ΰ?��A ۂ�1�I>v�0%�F�<��eĂ"�N-�3族ed�$��ːn�<�R�N�L6�T��&l��0y�BJt�<W Z����aU���lb�Zr�<��?d]�����T�B��D��b�<a�K�4䬐�D@E���b�<ipݎT>�y�s��M�\��u!�F�<9t��W�:��珃}v�9��
|�<I�� _<�lj��?UJ��x�<�T�݇4tv���c]�.�H�r��s�<�UtL��t`ڼG/2�3bm�<��Ԁ`�8Z��FL�>d�c��h�<�����
X�e���|y�A�@"
\�<
ֿzXH����P&>�nq#%�V�<�1n�0mȰHyS�!����g,�w�<�uᑬ*w>mz� �~�����t�<	�H"�T�Sdh�Ui|�z���u�<��Ɓ*%��ۡ��o��!��K�<�UlL6>Ȧ�b�A��9q��c�N�<B׈4��H�"Jl�IP�ʏM�<yB��@'��7-D�:�����n�E�<y!�)B�>�Ɯ�N͌��P͊�<��!�ho�S�����)��s�<�a��h����NȪ?f�'�Y�<ٶ(ʠKC,����'5
�\p\�<a�fи7]�LK��_�w���+7ƃX�<)v�ٓ}N�٩C��K����B�V�<�R.I��O�d$�0Z��J�<� C�H?5
WiG�~eQ�`�<�e,L����� �hp �	Dv�<�t�>'��2PG��F/���U`r�<9�͖�)�<�Xp��U�H��u�\n�<i���0=`���65$�|ӓ�l�<!�k4D��Y�6MO�-�PkTn�j�<���,k(�3�*đzg�`RB��d�<)�HV<����dу/������Y�<���_�0���[�G�=Yh��F��\�<IU+H�J@
����G::EU���s�<qs��)t߬�A"!E�&�4OF�<��dC�@��0���U�P�Q�"w�<9��*@X��a�n]�%��d�g��s�<!��a\0H�]�-�~�{�%6D���2kL�k�`�0a��yE2���T+����ͅ
h���mx�T��$��7b�		�mE5@�4���3D�t��ę
�2�C�arD�+t�.D� �`M�'FPa!�@C\�1,D�A���']�`H�w`�2	���hc-D�|Yj'9�2�)CFԸR���Q�&D��*֡&2��U�p�H�Q΢�(�M(D��0��($ʨ���`
�B5^Mڠ�&D�p{�G�C�H�e�ɞK�H�!�%%D�� di#FEJJ�+C��y&�a��"O���!��4X��=Q��C2..,���"O��$FC.Ei�e��k@�	��J�"O��p%Jx2��k@�#�\q!"O�I2�$�+Y����v�3h�|m�"O�!�ةIB�0#��N|����S"O6�0�H3Vc��d��.'Nd�"O�U��~�S�A	k^��6i;D�����^�$�]S'��_E���;D��؆ Ed��P�S�=Z�K��7D�Ē�ߒO�z����0 �>D���� �!I�´QR�
�I$����+D�T9�A�#Aή��C�I$z^�R��:D��6e�-���p�E/�$!�W�<D�<���y
�*�	8�REx��=D��
���g�Lp""�.Sx�*WM6D�d�vkF?�
-��]� t�wo���t(Q� �qO�>����O(���V�Y���6D�4�P���12Z1�V�ѥe>�j�(�<a�용F�d��Ԋ-,O��ȴ�6���s�H	
�H�J��'>����5�~ػ�S6�$X��#M���L��
ɽk�>m�pi�ş"p�L��ԫ�IJ��~"őh����4M*s�Y��(O�]�ae�k��:G��'�ħ1�b����3`��(� >><���a�1��M c�D	�Ã� z�f�	��1ړL��9�reQ�r�W�z�}�T�[&P�i�2�W;4��7,qӈp��ܳ.V�
� �@��9Ҧ	�N��5���������o�<������ؿ	Y��xq
[��a}"���6h����kN,~F��w�
F���r��I�����}g�\HTLM�5l���os�H�o���.�Q`����O�BN-��a|�QGغ��TcA�4[dL�\��=Ս�1�t��UB�-<<D�ꝠPފ���_%I�r�B&��)2�-�0�|���B�)4,d�J�4AҠQ��c�1�c +�`�'f�+DOU8o��m����b�.�3���;B�H����ekNe+��\$&�X�ˆ��7� x1F&U4Ws�m*Bi;o :	+c(��`aZM{��D��O0"�	�A�"8
x��hd�U�t#�F:@"�A6�ԑ��F��K8,�9daC�'4H�@���mo�y˄�_�l36��K��� '�?Z�D{�Ä�T'q��	�}�&��oҦh�V�YB��{����	CF�:m���kb�קs����ICG�8e����UiBj#�]�0������yF`a�LZk~9�-��q��k�-"����HW+D���@�%�ɘS��+b�~q���T��
8"/��<���6��&^)�A�A �����˨d�dM�1�20�؁�E���Lܨ	�iX�k�qOt�d��7az���fN,.��D��A5M��i�G�l�x��U�qm�GL$,�eH@r����Es٤�0d$�]�L`�-��X�)�m:�d�q�Ⱥ��85ި��EiŹ*�:aS�/nG­c���\�@����7w��V$\�0Ҿ�ۅ�'�$a+7��q�Iy�r�D�m͋U/|4H�H#�`=a�K�r�д��I
Z�bxbe+E; 0���.a�P��e��T�R�ۧ��(��$�^�zD��:}'2���՟�,~1�ȋ4ɘ�A�@ F���l0A�	<ȨO�M�1䌄c�2|a�hǐ"���˔Iɭ$>�SRk5x}�Pт ���� Bӿ'�.y�G�
#v6M�XF`���W�m����b�.�%�h�x �U��/D)����6��Rox-RA�/␹�H�w7�zefV!l`��2���[��\;�W7`o���i̤qZ������)u�tq{&�	���xb�E�*B�jg�׶ch��3��%r\���H��1���!+� �`tE�S��*Q�w�^5�2K��BN0k���)��q�U (��@�q��(M9M�l���_�H���j�8�j�3#A֩��)  �\��%�s�?�(Ob�;c�V(�R$�
=�
�@�!3=�,��D�	5j��NA� ��4zS�J1Z0���G�9��P
L"2<��݅�"�� *�5j���tM��x��A��Ϻ�F�<� �D�i������z��a�4�8�Tt��g�0\\ة�eќnf�	�b���mr$Pc�ğ[��F��(|���S1]\แ呝le��r��lp x�.�pZq����W5,��FN^Ο�@�|� (�Ó>o���@�΄!xN]��aL�R="��.�V�DrB��*�H<�2e�<:�B=��HJ$C�Y��E1/[�؃�
�O�|ab�?��>)��(t:��F�;Ѹ�*�8W���jG C:h)��S@Mˠ/���h��L��܁mWUQ}�`O-Dl`��BZ�;�2`��k�O��b� 4z%����æ�(O>`��kܢ��.5��Y	�o�.'Ǣ�Xp ì�b1�t�\�!���RBl�*�r k�L��u1�K�&è�(�@B��z�oE�\�2�f�F,Z�+o44�R�Gy2KE<T��Z2��C&L�"/��5�^��aG,D���AU��[}��e��R�b�t��W`&؀U�UX*���.C���i%F�<��&������j!�hp}�/[��i���O�	BĂ�:;_��jbK^'Y�d�P�!E#꨻�٪ ��7݃)��; �Tm*x�¤�O�F�I�g���F�؆⇯Mx�ЦON�ʁm%��O�!ز��Pd�2�
_�a��[oZ,Z�: �ƪC��F���� )Q�8r�G��M�:d���?�(Y
c��)L8�#��}I���_�4��РgQ� �bn�?N���Ko�<aNX�����+�����r��k���4��Ra`a�-L�q���;���:�.ܡҁ��^���_W~I����"l��ƄG�#g
">��kJ�j8����ߐ��#D�/���nH�[ƅ���a�4��#C�vaI1E݊V�Tq&���88�C_��O p�A'L�����LPNMC�=O�xڤ/�����D�T�%�*h�e���N���a�H�I]Tyb�CY� lɑQ�W���bd�H3{��4�����|}��	#	W��+Q�̭V&!wlY�X��9�0%��=��"5"@qǒ��e�ڠ[��Kᣍ/R"'�=Z��睢�v<"�B�}��9�@�fD*����%D&ᘄ�0c���ȑ���yr��L��<K�N�@���p�Y#R�A��ˈ0b��Z4����e 2U��#FN�0�2�s��q�M��0<!&�b�x�r.>M�<X@g���u�|�24���:v��D��І���gh1/yj�[�����0<ad�	$������D)7����#��?�.Pph�Cx5I%��Q|�q-��,�����HעY
DT�p�j?(�i	�m�P���hH0���3p���f��=R�M����:?�,�P��i�@����[jN4��(�8�ib7�`B�W?��k�����p��S�'qj�
6�
�w~��-��Bl&	�a�P��!g��:yt(���d�$�ؤ�t��AǵD����L�&Lc�I;Q��(C���l�����9T0�"?�5�Gy�qk@��܉�Q�*XJ2xy�n�]P�Ux͆�t�l�B7���pM�Ue�d�|	,F+v�>�?���2��)�!ˎ��d��b�\}2�!\z��U������Px�� �E�]q:�S�K��ņ���OJ�v+`����[I����6M9���`��j���rB"Мz��r�/ٜOह�&���$,��砘,���.ۨi���*�BQ~��J��y��i3�wh\y�dX�*Ђ��,.���	�c�p�I���9 �����[��} ��$E�n�C��3_îl�ʘ%�7�{�HJ��V2.V`�j�Aȃt��L�$M`@L�vʴɅ���C�XF}�(�|��3g,JX�]k`DͤN�,Ap]���9�#�3iv6`h�/��f��:�`
�r;h ���BQ�za+����F{B�M`���ek���a�D�<�~R�ŮX�D��e�1#R�:�FΰWX�OR�$["_�ta�,�1 �7��]%j�\t�E/��\�h��5P���$�$)6��5���/��,I K��&L8��0���Ӆ�!x��"ȇAF@z�+:Z�1b � ��];UB��8ũ�VݬUz$�i岱[�HS�a{��u��4��"�B	\����+U �Y�I�Z$PYd �
����!��:�⁔GP��ыJ�V�Q�O%@1b���(f-�"˾cH��Yh�'�� BW�E"��s�L1�S�|&��!�v�
�!��͕4"D�Ba'C��Z�Y���t��T!�"��~"���u��aw��0*T�ٴq**�GݰJ( 0� Eo����B�Az��B��G����.إ�`�L�5Iz�k!!��F�y�����?(�#�D�t���ӑ$܅}`����B �cNey+�?L�Q�剫/��La�6�*�j�6$����L�t��C��X+�`+.��X �(�z$*�6$���hL�h���!!�qPdsǌ�3�,�˦+�Ŕ�	'�'�(���덣v1l-��]�L�U�4�*D9b7�V��Q�t�L���a� q1j-�A	ݗI�qЄ�*E%Rg֡�:�SV��.�f�k%�O�!�Т?� .Y %�����?��j#���������`N��fޗC��X��ڟ�XF�	l�y	��L'5����W�aL��qf_�E��lzc�K�}��ڥiܥd���r�[�Z�K�p�3���5�������Q�>����Q�L K�+��-ʄ
ߠtV��`N�HJ���.O������=d�h�Dᕎj��՚4��#yL�Gxb��=f��J��\\��aG^�����I�@C`��P�D����i�e��
$DV
WD����Z�����Z�$U[�t��PN}�����ӷV*�P�d����q�������؁#n�=��0I`A�
�TPXaa�`���끉�܃�M�Ľ���+���C��LnaC�D> �>\��I61�@�K���6.��%��P�U�pT�	�``f`�6ŋ?��eɁA܈C����hQ�؁#
�Y�<H-I�bcnxӶŊ;�93d�x�+Ưp�h�J��
W�V��L����kļ�P�,Y���0��-d�1�vlM�(�^���&h��7�P"�Ȩ���w��82��y^�q"��+�P���$W�&����'�� 30f���)�'�t�P��߬~�@=b�C��}�P�q-V�"���,��16h��	 ��l�0�K o����1! &�e�D�Jt��(��O��2	�0:��C+4?s,���ąaJ�R�L38�8D���C�?�^`��c����A�9P�!�b2�~��X�%��܃�(�G�D(���+GP��dD�
d��� ���pU"0ʑ�U��m�"@�L�V$���q�YD� �˃�9���0�B�:޽���� i�(L�c��M����fmR\����/@X}��FW��������Ȅ�R�ʫ1S���PiX+2NS��ݱ�
H)&M�!�q�b�8������d�B�s�葕)[�����	�"=���Slh ���k�K�6�"��ŉI/6m��o����t%D��4BRi`.�����N�,�JB��
M&*E1gʌA�FL���
o��5�\�uI��HČ�% ,����Țe��A!!�Ƞ`�̃���o��v���4
��<y��8��40�,!�ҢCD���'���\��$�$D6 �ZB$��q�2���#��3šN�wf���πV��DE�oiA��>� x3�G�+@f��"���sJb�+�ρ5s�B��*7w4i7$?�TS�ň[��`14�X�X~�Mpg���'ؑa�'ȗ"j�#�e�g`v�i���Rp�P	�A�Sgz�:b'�0�h]3�ᜓ5-�8@�FV�%x� �1�� �	s"Qbt�r�gHr��|��0��.تk�X�"�~��w�L"	z�FP�F)bQ�gǁ�x�����i.����d���y0�63��X�@E��D7�3b�S��ة� �˧_|%�C@�!E>��D˚P�p�e�=L6D
� #R��Q%���qQ��oZ	ADn�{��K�1��4@��}�~�H��>@E�dI#j� �����Ԫu�Y�A�bz*��$��DPr�@�f}&< bX�˞�J��)#�I�m�?��A��vJ ���ٴQ�T�SJ�˒�
g��/(�mK�̀�<�Ш��.��z�k:L�������q���M<Y�%�S�:�K��[~yb�	ܞtZ�A��!��å@_������dÌD�:�{-��~��Ak�I�>@*� 4.B=�B!��_7����3�"�)� P�xQ#V�2Bh=�N"J#�ѹE*�9v�p��WC�,�T�^�]�J��C0EbPd�
�M+���%���=�tB��G�`��(q=xhYJ%p�� 4K�Ts�<A� �p>~dI&j��t��ZD�� j-`�k����f��t��j�(C����> iF��� ؠi(t�s���a��h�Ѫ�*Fe15��� v� ��%5"ܨ���d���(Wr�k��0���aGI����0o���ɻ��3��x��Y�0�jQ�����x�`9�  �	A��i�� ���WL�1�P���5�pe����'���'�_�C�xF( C�(�z����Dϋb� ��qaC3!���w�߮ F�0�(R�"SM�[��5���O�`��悔�J�åi�]g�|��H�9h$P�p�|��̘n�'�f\[5�D��a��a��+�J  M�P��th��ߵ:��,U�pl+5ˍB��]�s���u� ��V��)�z���*�L�1gz�{�&�3��僗-\�#����5$Y#@j��g*��b>+�-Nʼ��r�����׌�6���al9+���� �yƌ�9ӭN����3��=sB�5> &�b�/��\P&�ȗ+����p�|�KR����(�C����%z�8a��Ο!Z2�"��\`�b�b6�pHC��7Pd0��֩/Rl�'ᰁ�Rc�.�@!@��
I<�)K7N[�yb��d��<A4�ק����́��~E#��H@�taZ��@-j�X��ȗ�a�� it���������luC�N� <�>�8���(��&��s��SI��)Y!.��m�΄���Y�0$j�O�hs�Q����B=V<�J��V��X��G�)���at#��Y�: 2�l��n}�}��MD3H�����P�pD�r��l2��c��ESTp��'���`RM7maA������9C��(B"<���Tb�C����6���J�`�!	tu`]}��!7��Z�@���
�ȼ~2��֚z�<EP�>s�T���A�I�r�X��G�͂F"~��7KӅf�>�[7���ĢV�l��$���`K�� )Ate�Qö��YL�(��s�Ԡ�gB�7gz4� �\;P%$,�LL8,�\3��È4��K�b�i�ƀ�7"7f{�	O�ϻ,�:į� ��P��Fu��ȓ4��� �T3]�lfX8`�]	��N��R�@�N�Cc��;q���5���a�U1U�O�mZ�k͹S<xѲ��٦c�P�0��'�l�㱬0n�R{b/S"_f@�0��.>Ვ����.g0X�&�Dl̢c�[��{*���J̬q*�����'����`O6j% ,0@aEWfl�km^�<�x��'OGx!p���X8�b��-��*�hBa�ܪj�@p�D�
lE�L�B�H��̥�޴N�n�x�jPٌ�&z��e��A��.v�dy���50�!�T���,M�`JIX#��1�N�@�Q���p#�'�ɝO�΀Dy���mG���1�
0d�q�i��y��D����k��f�j	�􀊶�MˀH�<_v���J�Q`��tG�-	����\�t�!�D]4g��L��%�.p����1
�!�B_�Lk���E�x�S4"��!�K��b&k�Rg�0ʴ�Z��!�d� (�@�P0ڵX~�(7���s1!�ւh{�MĀ$Zʤ+$��1:!��+$�����3F
�U��9-!��R�<�C�C	N7�[�,��<d!�����H�*�1kۜ�K�ȑ-{!�dW+O�$H��ڇ�V�B�hϕe!�$��{� ��P䍬�l�Y�(�QN!�9�V1q�Yw�j�BG^`7!�D�4��	,@�R�wj�x�"O��i�O<���J�lB���'"O �`�Kd���9B�^I�T"On�9��ŭz2I�g�N�rq"O� 3���=!@&|���H̸���"O��+�c-��ܹ�)R�,�Z�"O8����?'��A�C���X��0p6"O��Q�׀\��)y$�;0l24��"O���s%&^�6��%�iT����"O� ��ق&2�Qkq�\J�p�Q"O�����`�\�.��_�!!�"O��c�B1�
�֫�)_\ݪ "OTp���H�9ɀ�*�L�AZr�K�"O
�R��<r�ѳ�	�v�f��"On�s�!u*8�0���w��eA"Ox:�c�� @8ĭ�"[A��Qt"O�1�S���6,z',�4�~ �"O@�3&�Ɂ;z��$��
����"O��r�#}6�]BT��'��bB"O����T�T�2z��ܕn�PPQ�"O�8e㚋}9������5j�2)�%"O� 6����@���2f@4��Yf"Ol<���8 �&�$�Ӛx"9�U"O�l`􂃖��XaK�*'aꥡc"O��C`��)Ak&�T���}��"O�u��!,�tݡ�`ە�pD�R"O�S!H<!�� ���2����b"O8�S�l�������H�LESW"OPQ����-� Uū�V��Z@"OP�@C�;hn`�BQ��(�����"On��&Q��<|
������Cf"O� � G��vͪ3�T�8 p"Ot��a�@�(<k����jU1�"OF�IB'^#�tM�Ҁӣ9tD�:7"OfYQ��t-�yKc���W]V�R"O4��W˘ Ni� ��R�'���"O�����ݙ��I�o�=v�6P9a"On=���X�"��	p�Ȝ�f��ͻ�"O�aK�`W!V 8�f�y��e�e"O±���ґp����$��Zz�M�"O�\I"*��ሊ�I�$�����y��!����w�	8y�G&�~��̼�Jl�=E��㟃�S1&�mN�B�H��y"�]8�Сk��I�v5T��T���'"�� `-�Ұ<�ũ3n�t���-ֽE8v)��@yX��0b� p�2Av��R���� �!�2=ju�\�v�Jua�
�qO2S�W��	yG��W�'K��I2$�����U�^Q���,���<�A�_�&���ЮT�\�P!ZĬ��/���B1F�!E�pi�E�ȝ��ب`�Bd��+�pI��\	�hO�̣!Ԇ4hD�;�g�Y��<#�AJ�{NqF�W{��5�i�6@�g(k֘�'*�3�ȹQ�x�$Dh�+I	{\��JI��1ѩGt������A���>�GM;H����m��ճ� D~�p\�Ca	�Q��k�>+F0�7��9F�� .مk���Ҡ�Ҽ+2@�)Ox`M1�`?&�v�CEn�L�4��K�v1r$A��U�
�PJRC�<-�IU�Q�I_�8q �'!9����BZ�UiI�Z�XR�ν(�Y&��MW�%x� u��єG�P����%�o]*"<�� ��)�sI�%�u+��˫ٴLh��$�N�F��C��8�ub_+:Vb�YB��l��`dhͱ^ ����e�� �Z%���N�'�f�p#�]�dG�< ���z(B<�R��4�ʵ!�� eԲՂ��(�v�0S.ݙ`N�`vMڮ|#Z��lW3��b� Jz�;� P�X�T$ӷ`�(L�@�W�r ��D�B��(1�Ωd��0ʓ�&N|b4n!��*�����6!)R�@�D��
�뎩�uw�C�H@�,I���:�(\�1�L����m���n9��ɶB���Pt�Z�" y��[�uu���>��S�-��m`�C�� �S ȣ=B�zk�sx%A4Iʱ;���P���Y�Ȑ2����G�(<C�L���E��'M��`�"ƈA�8�T�U;�T�Ib$[2 h��(��vL�tNM�VP�Y�F��� ���I��lr�%ԛ9dq��ߎ�lx���'[J�	��x�+-ט���$]K�hzgj�48�"U��XZd�`�5DϤr��h�s�R+݈�EF�&[@�D��?�"i��,�f��.0���5�ˏ�PT�sl߃`���@n�Z���N%,OJ]2GA	���0B�A�/��Y&t�$" IN"� ��'P^}z��� �� z��/���U'qBW��xuh�u�­>���R����R	��>�G �Y*���i˯�R�y`
#���D�˒!�>3W��(Zg��(�
C�<y�3t�Ա�ݴGX�;CHB� M�UR���8R�����<6�5�e���j+`�PFн �O.\K1�G�;����@A� ��ӆ�7�b��H���XX���nY�k�`Q��/ �Z�H���� �����c�����
F�Ɣ0���/h�|i�h���\�'�:��m�_��#R��D�<*êҎ[ӎ}�u(�%\\�"5�*���4^��B՟�q�	��z��AC�G��(�����0=���Wi��6�h��o�K�����/�?����7�N�=��Á�H"Y�q��Ș�"kb�#���(�8Yreۅy���YR��?���Ѣ�&P�Y��ؙ�u�玀;�pa����"<��D�Df�6�a���6�(O~a��� 8�<�$ Če�&�!%G״N0�!�);u:|��Í�%R����u'��$�7�,?ْP"E���]|��IS;u4x���I%S����Ug�������K�b�4HsR�22�HD`�'����O�6"�JcC.D�TW��)�+K�g�.|⫄�1��Jʱ2�z�{���!aa"�;���,�`��"��;:\9B�fùwv�b�'�|�k��Y�|@9�$�k%%G�}Lai��U� JŹ3�B9P^z��T�g`Fm�O̭���;��;�w�v����خ+o�ujQ�J����
����rFY�����(:ʓI��	��>h� +��C�+�$�E�җ]��Qf1r�6Ԛ2/!^�8M�M�b����,*�,ڥh�W��ca��n"�x3�]�$����`���q������i2���"���P��p��̹pf��t�HxFk8mpȍaSj��x�})�m��c�l��v��2�6!���p�x�yy�$�i]��k (tr�H��t2�Hq��?�q���0&T"wA������K�(q|� cB�$p<�pJ�B,��vQ�b��=�8$ B�pR\ �Р�)7n��S�Â��	�(Ph����)#�JS5��|���Q���a+�b��U�nP�w�Y6��r���+'�^(3��G�z���H�]�d"�]�e$�ASኬ"���D�,6���+���R0���PRE��� �j�+S�{Cl�P낀x<�8 ��)&�,���$��<8���ɂ;��*��S�zAh�`��z:�$�'�X��W�ǡ���e0Z��]��DЫ\���x�#T�!�čv�6I�
���/
�|]BEp�㖿K�Pՠ�dC4w���%6v��D���<A"d�!�Jx�'�R��_�����4�ֈ$@�؛'���9Q,��N�f�h2�X�?� j��ø���
"M�5�jQ�p�P���C�50�C���� 3���#�'�r�:���q*���3*B~��+#LW� ;z!['�H>�.��w�P�5�h�jp#ײt#���C��|��3�wD9qg�I�]�R돾x_z�0���$j&"��4���ڶ)|HRUo�5p4�8A���?�aK���S�h�ysG�0��s���#hl%��Y}�N jZLhEۅ9~�s�� �0<Y�"»)�,ȱ��9Xo�9��
�#Q�`�V� *���ɰˁ�.�j�B%��k�$�b�ٚ�HӒ*V���O�y���B�P-���J�\+D���$E�8�fp���L����r�K��6�B��jF�l�ؘ�`���h,[�,\26J*�Zg��83<��	�"�|T�6m �m���C9v)�� ��Ƨo����@щ(_:�K7�&�rL�f� 9l���ܭ��w�xu�P�[2b�P��5)�H��'�|}� +�	C�L��A�8j��`A1(�r�^�T�T�Yl��v�K���87KE�B�F��!��l��HAX��)Tʐ�	>>IJd�
Uj@ai�K;��CT ��t��0t,^�A�,kw�r��	�l��24l��f(�:�䖅49�L�֋�A�
�*V�Ӯ'ObIP��I�@�,0
u��(N���qg��;�T�*U"��$"[���+A	�Xq�" �7@F-���I�O���IuM5������A<�Ѥn__؟蠇�] S�bD0D١ 1��`��Ay�p,G6F�"B��2W����U�v`Sp� #6�F�����VKKC�nMQ��X�cΰ3��J��$��,)|��1B)��F	�F�:S2pX�w�'�� Y�iU�kX�#5�i����I� @T2E@۔�F��AY�aŀ<%	��
��ߏ_����!�V���K�V��ٸ�
H�8�I��Κw� �z�H��x���%ŏJШ-!�D5kt N9��D�R�F�mҸ�3�|6�� ��O��݁���������Na�ĎO�b 2����ŋ?��Xz�	��|R���Y�@��cI	5�t�v͛�u�@y0��	;^a��mԺ!IW�'[.9ʖNɞ%���5B.8�S"n��IRO��*��qC4�]>�&�� �楃�
^�F'4P�w���@�ӑcPE���J� O����� �:��I ^�9Q�@]�>���j�A�H��"#�6p��呃o�.A\�T+Ϩ1��u;gL�9���Z�a��I��2�|>��OS�-=�AA4�Z�����cҒbTQ� ����@ɾ����?8 )�Oo*�b��3 І�Ps�on��b�C(Cj~ b�X�0{:D��FG,/l*�r�&�!Ԋ���	h~���b����#G�J���T{�R��O��H "Э*��{ h�+lF��'
��BJ=�`��^�rxq�,��*��]"��E�!a�5V[� ��\�lܧ�VL"�c2�Y9Rl	�/�Q��' &XJ� �	�;_x =r�ȅ1czhj�唊�?饧��A�J��@�^Z�p�C8Zt9rhD�b{�a�"4$�$m�eFB�.���b�M@!�`��Yd�y��$�x�$��MW%R���%EP8���� KF��d"�xD!�IWF9 �D��LS@�'@V8ل%��9�/�sX�|�V��{|lL�`�!��O�iɲ� H7��̓�B���#-\�PN���ìu�q�a���+��3������2�'�5�2,�".3VE�%����-w�}���-��)KezC�X�A�ŕN��I������'�B9�6�W�=4�iw�ޝH6Ĭ�RI�1l�nW�G�';-�۵��`2�(P�͝8n�I�Ӣ�X�dEZv�S�����S��7>&�!�e.�d�'~b�#������� �X$(E��G�?(��1/?��m�"�&
xh�+�BA����X$6�1��;;⡘Q��p���Ag��7�pQHЋ�ydMa�J�wc�Ʉ�I3�!�(��m��	$�B�!�@���Y�O�
���X�@p.���D�4��4h��l����&�^�?�RT����K����E�:7����[�����=�B�Jj>�5�xޠr���j�
Ɂ��S�Y�N��M�"vN����Ql.�e�yڬ2w��n�Eʗ��l��+�g�7~���c��;�ɳx�~T�$�@.�6���Ȏ�i������6J�����8R5���Df="�2��A�{�N�3ec��-^�1f���5cL���Q2��Gx"�̝y�J�𤁊3<��B����6a���G+E�H����-B�|�:��͟}�F���!�2?��4�W�1i���gE�A�x�i@#�$?�R)�jф ]��X4�V�0�@��I'C13]9��|9�*�aH�� �$��4�ҝ��N�,�I'���q���qo�, Ui�!I�%y�H��qj��`0:"�{��Y	{����␉!q�yE&��Je����B�e���P��Wc�4�f�]$4q�N	x
�)��M�Oo��q%C�`���@ܦ@4Fީ_�, ��H%�ti7�*��"�La(�V��E@4�P,G��X����ܓ�ċ�O<�B�m0� M��D؎]E�̳Tc���L�h�H~A����$��J7����C�����`*ŋsQv9�Gˈ�<8��!	�=�\�h��V ��$�QÒ����*D�u\h��K�32,�����N���$	��^��d�taRֲP�ĉ�H��|�Onᇯ�(g�����d�<e�4��~�Դ
V�ȎlI�i`�����q�o�U���qH7!`�T9���Vd_�Z@�&F�=a������'S���Mο<�DY"�=�X�����44�2	�A�)��Ջ�E���DC���M�
���l\��N��q+61�"�$���-����0�Z��Ԅ���I=F\���,�!��'@&5Q(8j�t�KSj�7#�YI�S��F��F�ǣ)�
�I�n�$����^� �N��r�e
��и#Cѱ�IQ�+��G.f�[6��"X	KG �����"f�N��5#�8b)���Td�X/�"f��_>��3��i��T2d���3Ɯw��Dj3�!Jl(-�g%͙����<��|���I��|��I�'�Փ%N��J�D�:�lSΐ>o]�X �4^�Q�'��mK�-�MJ	:�e.�v`���c�? u`�߫'>��ݰ<J��u�'�n�8�nY!J銑(�q����I�B���i�iȈ	�,IV��=���P�
� ���ؐ�e�����I�G��9`iI	�
��O�����$W�"Qh���w�"�M<�� �.?�aZ�S�x{����JҤz݊Sn'&�<1��Tȸ���%����:��Y��L�>��qi��ݼ�0����Pވ�#(;��;}�1��aR%��27 �y��� �2�`ª��rl񷡀�z�����!��R����7@[+o�]1�>b�ܨQD'��<Hʕ�Qfܖvڢ���Z�'�ޤItGA<=JΑ�a�\"f ����M�3F�XP劳��,��<\�xm����X�C@��!a ��EM�0F�H�EK3��4Rvb9�D���M"dt�١ȟ�t����@�O;tdR�GeB4?k� c̍C�����vQ���E�{��'
'jx�tHp�
�	TL��'MA�{,�L�V�I�k���Ѕ���<��"%i}�T�&K/_2��	҇,��h��"\9
�i� �C�8�.e�̏'y(ҡ�`�Y((�SiS�(��d����=�I��%�9�di�Č�tTn-�w���q���9��QC�T���{H�oܞ`M D!e��5q^�P�E�_�iլ��GHM�H��wNG7[K�9�&m�~����da�|x��^�nٴ�����?O���N�^A�=;����f���Kq*�D�9zF��a���AVH����l��b�+$� #d���d���{a�+k��F�R#T��%��cC3&�⦩KgM2:�,�15"�AB�l��8I��i���c�G�%e4Xo�!}�X�dK��<����K���<�ٛEìF��Z��H4M�̍�n�>Y�2�R�O �"���h��-Y�n�kp$�epA1�
e�pͪuM?C�mZ��@���`֌�[��D��dsU�''0t3�n�<��}H��X�Q=x���b�e�`���� ���c5�F9.$\c6nF���yH��@�CG�=%4p;�D�w��13�@@;U�� ã�H�=�NDRwM\�q�[�tF��"`�Q�w�0�!f�~a Y��X�F�Cwnfx���F6G��j�$=p�,,�a�G{j0qhS$*�V՛E��7���	q&Û&��"
�6���I�F� ��-bR�<Z�̋�c.D>���0i�&MI��qI�n5��"Dۭ��yD		vqO>eZ�T?����S�	WJ����ݩ/LR�f�Oޑ��a�~����SF��q��*"Z�Ζ�{
:0afq��e,��0!�97
B㉍+Z�kP)��*�x� ��[���% >�,�1`R��M��H��/\�{p	�|a �y�FӋJ)
�z7f)J��F@���yR��}U.�X��:Z&���$�hA��ËC�޼��R�*��q rȗ~R>�D�-�	���q��ՒKX}�W��g�^��DI%��ԓ��T+^x��LyCR��7�B�A72٢��^�}�8K�"9y[8�(4Cm��l��,k����-� Y�����>�ɬM�Yc�˙=�b]['F�,m
��t��55���)E{��@�EO�=z@��Ҍ�!��8`�nl�$��D���*K�e�����J .7��<~�JqA��Ȅ��I���K����8V"t�a+H�$S�:��Gw�<��+0 �>�s(���~,�Df�����C9���I%3A��S LQ�j5R0$�P���#Ƭ6.��3�"D�(i�E�z/�����D `����M�2����������`��j��֏;��Q)Í��!�H�v�Z�Ą
mIrd��D��!���% ��dn�xY���l���!��� Xba��8+��K� <!��Ă|m"�����47Z	��-_!�D�v8��S��a.X�bf٣)!�D�%vNP[�D�(WV�8eʻ"�!�� 	�vٻ����`PJ�(D�!�ќdc�y��4J��b�A;<�!������4�S�t��q�GFC?!�d��UNP%�A�L�0zL��҆� !�Z����Aخ���i�EL?;!��R�������59Þ���C�r�!�D�JqJ�z���L���Y���vY!�$"S�F���皿k�PͲe� 2~J!�dD2A�����E�Ȗӕ�, (!�Ťn�\���Κ��
��G8	!�	re����C9[UT@�e��=�!��r�$�QdߋdF��;7��W�!�$�5f,�@�`@�,�6��s R�6�!�$�����蔮�8Ɛ�C��];o�!��	�*���G�-�8��b �ea!�d�!@!�̰���4[p�CVA��!�d��fp���](C����"3R�!�D�pLڬ��̺/2���c&�d�!�d�,n�=Y��['C��*�&�Qd!�$�86<���ăZ���VE�9C�!��L�hC�	�Ej�"g�Vq��cVD!���7	�lȵk����,kgO�7>7}c@[���)1q�:�?A�%�A�? [Pn{���d��7�L�"�1�4Y���� U�7�Rt�)�::�(j0&-�0[A
�A��	��'���E��-4O^��Ȋ)Z?�M3wo�M� D�t�Š���}}����Q��╦�3�L܊!. �9�|u��0��}����'(	h�	�o��ʜ���Dsu���)ȗ\[�QC�ݠQ �%��)ֲY��'�!�	�2٘��O�����N 4��Jj7D�K cy�&��B�@	�y��i-w:���`��&5�U�'�F�I�b��8jM`�y��)۬+ߪ���J M43ĢMEҰɲ����'�a��� Xq��Y�H�δ��S�*l$�M>�� �0|Jgb�=pҪ��'�ш
`��CQ�b����Qܧ�ħl���E�!n�5 DŖ6�:��'1���� H�Zɧ(�z�x�'J�L1H��?.��A��G`:b�D���O`8t�4�T4�1��Q�G�E9K L �/��=�`iV�Z�x�Z���>�¬4:�O|�D:�л#��$V�@��t��=�,A���@=;S�IjU�O,�yt)���h��D��Ge2�SF�>��� GM�m~�T|���5��)V'*�q��'[�lD��D�ߢ�'�B�K��6�)�'VN�`8�H'����7%�4��i��K#�����O+
wB�b"m��)�D���L�@K����{2� �0|�u(Q��*�k� -9]�OOP̓-8Y�o/�)�(_����d۶Pw�A mٚ�����D������8^k���&�-L�x�"�j�V� s��Jy��)R�e� �ܐR��ҳ��)Q�1O��ڣ�ϩQ�ax��ӛ'a@�`oJ95
%K��-�y�`�90QZ5�E:D(�<Q�<�yҋM�R*��ᶩ�CJP9j!㌂�y�7zk�@��^ +lQ���y��ݯ92�T#�fY���D�*��y�"�'&�N}q�㝰�⌑���y� R�"�<x��Ś�e�؍!҉��y�d��F?l룍�'XNԸ	�!�yBmA |��N�Z���[2��6�ybD4B�0+�)�,b�T���<�yR��`U�y{�ŗ�0$8QQI4�y���^B�Ȇ�N�U�(�a*J4�y�mLȶ%M�\�ՀR�y�A�!�8��flH�Jx�U�����y�K���J�Ɂ<+�Z�I�	�yR�3t�X�)�d�9Z�����ð�yb,�Q"r��'��?G�� �!ƍ��yB%�"X�,5���AAT�!R�hܿ�y��ަv2��"j�!>�hav�(�y�&�$��1����	��`Zv�G5�y���e1t��֎or`e��kJ
�y�I-����+n���Y�쐚�y"%�V��'ٕ[���Ɗ_��y"�Z+Q��B����	���Qc^�y7H��t�$f ��8&%��yB��n����@�6xq�����y2�� hB�q� ,>�W�1�yr!�ܕ:a �����C��]�y��p�h����\ C$�(v�G�y��G�&���Y@��V�P+ L[��y�&���P�u�_!%씵�0#Ǵ�y���,	�qb��%�(�E����yM�{%�� W�� �[%'��y".\"H��q c��*5�$C
��yB���C�84�C�7Xfh ��'���yb��4a��}�s�FI<jD`�3�y�l�P�����?�L`sE���y2�w��!����!>�M����y�$0^�x$�eș�Z��H� K�;�y2"�3B+������'[*�����0�y�i��9��T���Td��vg;�y
�  e��nY*+_:<�p�C���8�"O��v ߜ@dl ��,n��}��"O \��U�\
`i���	_Ƭi��"O����흃��욑I��!�a"O^�a҃�4vb�p���O�8��J$"Onep��0����f@ӯ4����"O,�����F}��A�\�j�"Oh=�G��)k|�t��i4x"�a��"O|�9!� x��Ӂ��2T�a �"OR�8`�J�����(͍J�ahE"O�yӷ	G,f��1{@��%|uDE
w"O(]ȕh�@�P-	���0n�5��"O�EM�,:�``�S�[���<�"O���E�>de�pe̅��5x�"OԴ�b�D:#޶$�Ф�'e:��)�"O�����&Yt|�����$)T �"OZ�Ѫ��3�eY@[�셐t"O�X��c+S������6:-�@1�"OL �F��;�`���Y3'|i""O���ul_�tV؃�ɀmJ�v"O:����[o�J�	�kn�+�"O� $ʙG&f��AJM��J�S"O�t���@u�	4
C�`���Q"O��"��
 ;r& �2����I("O�e`�d�bF^p!���Ds�D�p"O�|�c�/Cd���i
7lfTA��"O����hP���|�
�"Oz ��蜵&3����q��LXR"O���ƆF.A	�-8u��=F�¤�R"O0�s��#X�(	3�/�W܌B"O�5����='H���W�6:,�Q�"O��bd@J�H$:���K
�$�%y�"Ot	������P5\���"O�u�(��EFR1YpFڪj�Uۧ"O��2 |$~8
Tć�;[f(�"O�M�G�1d��r�I�� S�`�"Od��#UIxlr6�*_��<�"OD��Pm�sĤk��Y<y�4�zT"ODP��_a��ț*n��܂C"O��%j�<�0�Y扎�j��Tq"O�,��ą�=0ƁC�O�/{0H"O��Sr61X����nI���"OB�����'\0����["��!W"O�Ԁ��w��P�͇LP��"O�5�Q����is�1.�r�"O���A���T9�E�z~�zc"O^���cv~`$R��O�JY���H�<90�K2H��@���G:4��H�D�QE�<��-^	lNhI)GH�>r��(�v�<Q��K"��H��N�,�h�uLBv�<�c��!
9c,>�b�y�Lq�<��ͬ+�X�KDkJ�mDea��r�<AsI �J]�rE>��9��dBV�<!0
E�j9��A2�ųeV�@s��O�<q0R*$�
���+���eoM�<�M������}�X�zU�	F�<�Ќ� �z�'U�x�"��V'�C�<a�lJ�?� ��W��
q0dcCw�<��KٌS�h��j�/&������p�<!�����̨���+`�YE��h�<	d@C���Q�%%��|�ŏ6T�xSԭ��̴��U5���*0D�����Q� ��&��e��i��,D��I�*J�1������NdҗS�!�� ,y!�fF�&* � ��~��Qr"O��2�d��7n�x���]�ԨU"O|EرGJ>Mn��rIN��@��"O(	�NȳJ~��C��=S�*,A�"O��"q*�L����G�u�,D�v"O����	\P4Q7'��xvnys"O��d���T~��2d��3~��k�"O���)�BT�{�.Q�<��d"OJrtoD��]ᣍ�-	� �S'"O~pyeJQ�<�z�@'ЖP4"OB�9ъ���)A�ŋ�*��Ɇ"Ohi�'F5[�"Q+�<Q��9�"O>i��cF#Ċ�K��]�@��`�"O,��ʃ��)Cje�\�k "O���j	������*��~��6"O,�Bvh�S������U���"O���EJ�B;�d�扚�,�6Ԙ�"O� gnįLx�X�P�50�T)��"O�	b�M� lv�Ҏ�'V�n\��"O�H��J.^�4*��̩r�u�"O�1
㕝lQ4UJ��\	���V"O���5���A������9!2x��"O �P�fWgӪ���A��Fy6Ŋa"ONX�'�Z��!a�/�?n�1�A"O8LP`է5��J�.Nze�AQF"Ojy��
V{�L�4h� �G�g�<Y��տr}D(�,K1]�0� �QH�<Iv�E�P�Ꝺ�I�,f|E���E�<�eJA�$Ƅ�!�{��гC�U�<���y lH�t��5kL!���Q�<A4G8GRN��,ʴU�v�0��u�<1��-H�oEP3q$�A �[�<�QZ�(7��J�d�	o���҈�S�<��k���`З��vj�ك�U�<!����g�m�S�пf1�KF��Q�<�.�W;\|Ss�X�r\�! ��x�<���+u��T�wo��\��yP	M}�<i� �[��:�혯5��U�Hx�<�T�����Jɨb��L�aiYp�<�A�Q�%� b%NId9b���"m�<�p��W,֑���ej��x6��C�<A� ܈2���/|� �(oY}�<i��:Y�E�#d��TF���/w�<��%$Cb�h���&^����� s�<aWBP�!�0�)��ܞI}�J�DD�<�-Xb���ԯC�q8�!�f�G�<���W-��dA�u�lIA�FB@�<ѥǖ�:,p<��-Q"Q�=!1� |�<q�(Xe*�:��)�q� Gv�<9e�t�fS"&_�"9��{�-�r�<���;�����+�.�&�@`�p�<a�!�:Ep4;P��zhzeL�j�<�2b11$�H:�2�E���h�<��?1���ꑁT7
�Tqr��p�<ѷO�5Q��ՃC�N}V����c�<ׄұ�ҹ�����)���p��\�<	`!H3Q�, D/��d�d P�iC[�<3���m��Z�i��
�~�iC$@U�<Q�&;� ����!B�x����GU�<�G�[6��"rnN�x���`WT�<ѰlT�[�8�)ҌB>杁S"�R�<�J�)��P� �	%��)�O�<�oס7kz��pDX}����ѬTK�<y���!g>�R��X=D�m3e�q�<� Da����z8��@�E��0j�"OV�i7�[7d��o	�Gζ͢�"OB,��iԝH�<A��	7F�fœ�"O$��fL۠d�b��!l̈9�ȩy�"O"T�B� &z ��6K�+C �"s"O�<�&�ed�Q��g�_(�"Oճ!ʙ0Ү�efTvMZ��s"O��x`G[i�(�wN�j�>���"O"�C�/,�|��튊����"O��[��h�Ȃu�U�Q5�@`"O���, 4g�(� �n����"Ol�@]3
^�룍�l.0�"O�e��]95�dbЉ�-�J%��"O
D���X�;�R���!=�p˅"O����ޱ}wt ǦQ�v�<�5"O\�3�����FF��i���H"O"�P�W�AR���'�d�����"O��K@f����`  #�� �"OL�:����:���N�0B*�cv"O> B����A��]KvQ�~3��1�"O$�tH?<�jd�&��]%z�AB"O4-�@����(����iԨ)$"O L#�&:�Q���Gz�Ŋ""O�0��C�# 9R��7`N�woT�r"O��Ƞ�O�k�Pzd�چ*=:كD"O0|r�ٴ(�T���7!���"O��Dn�v�!5ɓ�J;Ȉ+�"O��1��
0� :�	]��p"OX��0�	�/P�}rUh���`�+�F�O���g�S �M;�O?�I�m�(�R���!+�[�:B^%ӆ�_1S
�aYcO_�bobA�P�U/Y���u`�Y�D�Ͽ�BlD4= ��r�9
wN�cC%���!��(16LhDC0kz ����\�����Cq����"�C�4t��D����L�7��Ϧi�`��O�QoZ����#|n��h��}sq��x�h�����2�N��۟�&����_��?�z�)9e��0g�'s&<�!K0ʓ��6�{���Hߦ��	�?9��y��Y�G�M���������X����C%�M[˓y0�Ig�h�T��R�	�c��N.*��um�3Ry�5��aͫx�tD�_�T�RN>a�g�v��[�Eͳb��hʙ��\!d�h�/_�cr!��T���(Y�~%Δ:��I�l�v�j2iU�1��� � A� ��K�j��	��M����y}R)؄/7Txp�g��yiX=��)E��(O��oZ ���8�	�l��>X��H���4�l��ՏC�M�W�i=�Gh���4�n��|*���5I����$9���{��߉.�*Æ���<q�.H�LK��X5��K%M4I�.��t G`��\*��f�`��Oԅ��\�@���(O��dg�B	��9��R6u*���t��2A��,�q W�uW*�;��еMp�DmĂ-f��p�{"��?Y�)�<��yp��P;h�"A��sVJ���x"�'���T>�E��~6���ť�<
�]YЪ#ʓ��<1�#��"���g#s������Y?�i`6�<�ԂŜ^f��'��OS�S��I�֩�X���9�{R�'�(0a�']i~��n��:��<��E�)~����6ڮmq�s8ܤp�#��(O�N��ah�I�&��H��I�SL��`�A��!����MA�h 2ǎ�<'|\[���:��'8��3��o��v�:��]ZKa��L���Өr��0�渟��?	��Dq�ƹqa�?t���h�h@\�C��'N�7M����m�(p�~��&-X.�D8�G������i�ĸh"�c���d�<�.��OP9����2
���j�!��1��30FA ��A&c�α ӤՅ ����b�ـe��]�-̞���C�c�"rG"V�;��7͓)	8T�s��z��˳aU�&2F��'��8�^�#O?��� ���7��0pa�qa�7���lr�u��q���'���iܢ�3C>[v��D�.b4X�'ў�}�⧀B��]%c�R����aR�'� 6�UȦ9��[w'�DqB��$���b2̛�Oo��r�<��EJ4`�&�'��h�d���҆�#
q´��,A�H���Z1�[��B�pܴYH���jEf�D�=�D�M���1��ȋ}1��R`.��8*hAhW	W�cK��@'���RT?�Z�"ȣ.�09Z�``�I�#�]�r�2g�֬�6b�>���Rʟ�`�4pP�'=��'��	�$Y��٦(��Tժ��3)�4�q�����'I����u#Ӷ=�昸���*!�n@s!�D_.��~��� 覥���?��R���R$�   ��   	  
  r     b+  m7  �B  �L  ZW  �a  $j  �v  C�  ��  �  ��  ʛ  �  O�  ��  �  '�  k�  ��  ��  1�  u�  ��  ��  ��  j�  ��  � � � ~* J8 �B 'J kP �V �Y  Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�� |d��"O
`�(�;���8���-0��1%"Oj4��ND^[��"3/9�0|H�"OB���H��*�ʞRy=a"O�味V�!X��!&F�:J�$���"O,��a
���C�Ą�M�"O,$3%o�-���p���+Ն�:1"O��ݢ1����`���y14]2��i�<�6��{_���c�H�`�fX�$Kn�<��A̼VI�xR[�)�Ć�pඤ�ȓA5��('nߡ4�� �)˩%� ���,��r�؊b#`T�eT09���ȓ!�b��g��}�8�F��-? �ȓ
K|m�ș�VṔ���2�%�ȓ"R�X�j�4JN�1�˘X�i����̹	_�jZ��1!g��zܶ��ȓgil,*�J�
j�Ne��i�J%b���f	�(U��:���G��$Y^م�~r�� S�%T"���k\�jx�ȓ|4�1�îJb��@ӵ�ݩn�V��/[`�"�v4�R�!ʎ<��M�ȓ`:��z�ؚh�J�Z��$HY:	��H��p�m�C1��!��B:��0��EnjZA V;9����J[
2���	��4'J�EA�IVW&��~�(aZ��ӹ�>� o�Y�|�ȓ�f�A�
Ο7�H��M�$�����mޠP����/���ANXo*�ȓTv�����{ ��-7�*h��I��sB�8�8���3����ȓNe*M�悡;������X�o��!�ȓ'lj�#F�m�+R&;�|��2)n�C��0S4���T:
b���:�0!��e֊��)��ͷV��,�ȓ0�&�8#���� ع�L�����;�P�AFd���,w�6d��r�EQ�( �gVlɦ�M,H��,DP���|�I	$G#\���ȓ"�)���E�B	yt&B�^�LɅ�4�� ��eëF�ڙ��n��R�p�ȓp`@}bŇ�=�$�AUN��P����L��p���_�a�)�Y�!��-��u�5���o}�`iF�@A�p ��F�\�0��[���IF/5���k>bTؖ�;K'DT`�^��@��fnV���Y�b�lI��	����ȓ,nٛ��Ć3���kC��8�m�ȓ'� I ���x<=���޳{��	���Λ�9L/��
�� V�]��f�4�yr�γ MR]�v��,,�|�u՗�y����|'D��"�8sf�:�!��y�̄�V�@��Hsg�������g�<�}���0^��0�2IX��a�e�^�<9���0W:@GD.�Ԫ��_���0=�Dg�FL���J�E$9�&JY�<���D�(�RÁ?g�v��PC�l�<��-K�H�����26��*�MLSX���O��	� : �`h���k8r��"O�����XhCH-�pȏ�6BQ���I���|Q:�M�<n*d@b�L!<@ �"O��t��;GM���3�T'Z��`9�"Oh�p��-G �j0CÒ�,ĉ��	�V�?� j�{C�R=1:�X�d�Wod�'�i+ў"~n��&v c�EX	Zߨ��k����{��h�<���B�1�L�9n�G %3�"O�
��^4e�ʔ;���2T�����>9�&�d��4m��fepL8�銎 ޭ��ߦ���OҐS��K?UX����\+&^�5��I>)a�I��(T*]����5��AV8�d:Q?����K�,���6�W V�"�,3D�H83�L�E�~�q!C��F��m����8����6a�Gf �>�`%!V*�;r
C�	1wb����(�4T]�v 4�ܢ?���|BV>��*�z�����T l�����(D� ��E�#J�t��*R�R��
��"D�0����y}�`@�O!~\��a �O�O�,ys�>U��6�6-[D9���LZ����Be�c;2�#��	E�������<	��D�?./�0�d矤#�]�1��'Z�5�OF�J3"�/g��:����`4�|��iݩ$� H
��Z�.�H�ȕ�H�f��!�:D�|qp	��ݠ�s0��'V�H	���=D���7M�1AU�C�ߤ���$�7lO➠k��7T��x��^�~�`��n5D�H�E�C�X���+�ȝU�(�3� ?�����.W�P���0�J�LO��C�	�V��X7��.��,y�m_L��c��h��ɒ��' �]Kc�ܸ��8ʁF�"_{�\�ȓ"g����E��;7g�zf�Il��p<��!M�6�* ����k�� Wd�nX��R��ט'�~�(��fe@���:=؄	��O����ɛ\g�8ɷEP؀�ж�W4+.JO4�Gz*�f�H��Q�b��MX*��B��` مȓL|>@`�	}ɖ�	�G�H�R0��b��""+K�W�\5�u�̚b�`�ȓv�}K�	���"8�f��7�4��ȓm�VaR2@��F���ҶIq6��-��H�"J�{;����I��
��ȓ{��4��l���HQ����)h��U����s���UꉳI���-�V�6�`��1D�|y�l�&
+0�L�M2���O0C�I�=�*)�b��u�4�#�͇����đc�ɹp��-�M^0��2G�7@hC�I��D�S�Z��v���m�a#�B��A,�jfh	q^8t�qM�(mQ�b����ɽk���VnH�,�	9g�lꓣhO�����?rQ��
�3a�	)%�9\2!򤆇7T�2	�(�
ɭ"��'��➘Gz�%G;|>�y �H(@.�c�Đ�y�=���J�������ɍ�yb��.L��i"EU���L�����yb.у>H�P�֡�{�8U�̿�yr�,r�s���G�,0e����O�"|���=�� ���"Yr���E�l�<fbV(Q�d
��Ph_D��2ǐN�:_L���P����'e�)2%X���Q��	�dgzm)w�^p<�W�̻�m��à�!�\
9.����O�b�"~��^0�E��t0#&m
0b؇�Z�8Ɇ�
�8�,��b��!|�����Uw���{VꎼA�P`��Z��XQT�<Yٴ3�O듴�I�o��	[ь�� ��=��@X�T�rB䉱�Zb��q�u�-V8<�O����K�$ ଓQ2��Dǘ8P	џ�E�ԭ�9@o��Qt��� �L�d��y"$Y��=���$۰�Arb��0<��$@0lʈ�&[ݴ�Q� !�!�� ܅�%�$=�΍1v�G�i�-
�'��I�>oU���H(��{�C��B�ɒZ3FtH��f����_�5%�B䉥��a�,F1O�Hm�F�*:��=�çW3�܃$���fU�QC��1��Y�ȓg���U'�5�H��CO��\6�%��?Yvh:�)ڧ=�2DBK�5y����ԍL4�=��/���(�(�%n�)���,����K!�l�C�]�J�hBJ��Ur`��ȓ����A��L�ɟ�H�����ɵ�HOr5��U�'t����e��(�Є�J>��n�/z�dqH�j|Щ�"E�<����ӭj���D�=c��� ��٤''�C�	)^2� 0'k�O�Vm��l
�n��B�I7�\@��V#F���"��M��b��i
ӓI ���֬%� �G�/��Ѕ��M�A�
��0��K�/v:���)d�<qt�@�O�Nd鷩��[���v�c�<iv��Xp��ŰK�������_�<�t腐w~�u{�,[L����F�\�<�W�&=�*���)(�Z�@�Q@�<�E$�=+_H�r&ԣZC��:���F�<�T�
:�y�O��.	�Hh�g�\�<�uB�Lخ8a�-�/s�h�C��Y�<!E��s�P�Q����A8)�H�U�<�d].]�����	������Y�<Y2Ņ�VƔ��T�||M�5O�X�<	�iT]����FZ1Xa��e�{�<iB�.Y'���FZ�����3�!�ۙYN�d;#�7���kL!�!��:���Fc+ԥP�+C�!���:��H��-y���c�	 �!��r�j��0��
��\3�Æ�>�!�	��:��3%Tw�I)�ͫ_�!�K�TZ�!֯�4@Y�3g�48�!�� �A��5]P���d*�J�!��"H�Aj���>ش)c	�^!�ʹ$]XD���CR(�|�g��-B!���-P�jU���̀T�\YV&�e�!���~�53eC�>uN���6%%Z�!���D,+6J��b�P�!�d���bU��x���z$�2~�!���68�&�kDK�f�F�SǯM�-_!�$1&!�d腇?7�fUK�-�-TL!�D4wKV���,I�N@�1{��\�,9!��6�1��]0C5��Zə�/�!��
b~�����4/�(F %�!��Y�v��-ڑ�V"�A7ʞ4Y�!�D��3G������5��i�	h!�D� e|dA+M�0aN��#(@7#Q!�K,"7�A��gF/FH�x��-5!��Uq�0uJ��e�d@��Â�f !�dA�/����d�[�m+�Hz!�d/zh�������zp�U�8�!���-���a�BՁy<����!�!�$T�&�j��5сg�2y��T�3�!���V���z�%�:P�i���>e!��V� `�0Um<Y �ӭi!�āSW!�g�ŋrWDQ3a
w!�ć@j0}x3ğ�$V`��A�X!��-=*l�`Aop��q@�.v!�dA�gu�I�3�G %v8��哑C:!�	X���p�Bh\�b�ν3!�ހHA� ��E	M�{�㉍1!�� �\��LV��y�
�B"XĪ�"O =��ƒ(ۖ�K�B=-"D�b�"O�ქ�\�ud$  3I2m+D2B"O�=:lF6>X(W&���i�r"O@��0�K	ն8�a�f#d��'���'Lb�'���'��'[��'�V�&e�>�0]�T�ٺR�6����'B�'���'�B�'��'7"�'�:�Í��c�	�!F=7����'{��'���'b�'�R�'���'I��4�X.�j�xL�t�"4���'��'���'4��'�B�'�"�'�1�WkWK�6\r�(@;z�B�{��'�2�'�r�'R�'�2�'��'�5:�E���`��PX�
��'4��'��'��'/B�'��'̣� N�E���:�̌�5�4�0�'��'�b�'���'�B�'�b�'b�M�s2"~\��S���%���'a"�'&��'6B�'3�'�B�'Ef����6x�P�#D�L"�"�'s��'���'O��'���'$��':x�������4���dۖ&��0��'���'V2�'���'���'�"�'����>v�P�#ׅ}��C��'��'��'�"�'@��'�B�'8��ß+0��`4�j���pQ�'"��'���'�r�'&R�'���',�I����*]�Hr�����@Y���'�'���'�'�B�r���D�O�Q���ĄT�h�-͛voܐhF$YUy��'n�)�3?Q�isDrmS9h�=`�-w���5D�:��$���?��<4�i�^I�݃\�U��[�Pm���e�u���Ĝ�w�b}kv:O����W�����6N���Q���@k��"1n��P�S�k�Dc���	RyB�k�R�X#iT(MI���Gҽ3@f��ܴk���<����e��nEt�8��@Y�Ӫ�K�e
(yցm�M�'��)��/VL%�b�����	���eh�����H���y  _�3"���a�D���t�'P���c�"]��0@���$�R=�'<�V� �M�&�r̓k̠q�q�ŪLc<HH�N^��������>�g�iY�6�w�4�'�ƽ��¬7�a�dA.>��D	�O:��� �<eX�p�)Q>T��r��O T�TM�m�T��/�b| 8v!�<Y)O��s��s� Z �&�j�H�[��XP�`��j�4Emf�'_
7�7�i>Q�B��,�jQ2�S�O滛��Db���4JB��'���2a-���Dϧ'Z<@;�FB�
]���d+K���0G��)����=��|�*Oʓ�Ȕ �U	
�t��Z�i9WM%��	��M��E�u̓��OI.�{"`�{*�(�6gj �䏫>Q7�iaJ6�o�x%>-��ȟ�2@���j٠�T-�	ƋW��bQm�>��Ű��p �
B�n�'f�c�zI"���#��H( �'��$0�����<9N>�!�i�}X�'��	3��H�EJqkXzNXxI�'Tz7-�Ol�O�9O�o���M#��"i����:|�=�"Éw�����*�x��33�(�pg�a�`�d��?���ͺ�Wdm�I;p��&HB`C��4i<-x�%y��IFy�P�"~Br�ߐP�0M#�eJ��z�k�@q�ƛ�P���d�Ħ�$�t2��(�Y#�	�7��$R`�<q�OH�mښ�M��6��1�`���<I���[f��Pg�_(1 �(� [C;�����I|�e#c�"����4�˓�?q��
g�#��$�n�P����<yN>���i�4�Q�y��O���M��s���~���7 <	������$N���I�4�y����O��x��N�'-�Xp�%(�^�j]h��s����9�',T�Z$�R�%�dYG����i�"W�B#Fgp	pR�k9��ђ˒�\�	ɟ(��ڟb>]�'�N7�W���A�X���	�d��`*7���z�4��'��U���GQY�I�g�#Z�͋�LR�:��7��O�J$�^�y��d�OƄS�(Z\%�!�	�<��ՃEC ��CI��A{h��`d��<y,O��O��d�O����OʧY�bȠ�֪t���RDI�Ait�iX�`1�'+��'���yRBk��.�/%�E��:u�ҵx��&DBn�3�M{J>ͧ���5,�+�	��<!Bk
79�� ��[+#�h+U�<��w)z���	��$��'-2�'�����m�O�L�p�[Ԥ�8��'���'@�\���4tv]��?	��)a���S+��$aR���B�2eӊ"�>ɵ�i��7*�dɉ@�(�06>[���4�8_����O�s#!W�u�ꕃ&l�<��)@�A��.Q�3���F��P�#BҦ�Rd�e���@������e�"sl,�&��8���)n��/-{~�r�
�[��4��F�Zº%�1��8�5 �l��(A�񴮞K�'�^� &'֝�8
v�ωe�T	94f� ���1��'��,8ɓ�Y_>�򱊚YF����ȇy��y�d�*�p��&��p�y�o�"-dx�!LU�?��Q�g#�"&܎��c��,u�n(g���l�,1:4�ȠNP"�L9뤆G��L� D�.a��Z�hM�th��Ϥz����'���#�0�4�|��O�˓a|dY��S]d���9BZx! �i��/�'���'/�R������

 �6�W�3�r�Ap�~0}�O<A���?�����$�O ���LH�C���5�f<Qs���h������Ob���Ob˓$"��I�>���[�"P�	F���f@�|*�e:T]�@��ݟ���ay�'w�=���ĚV��:��C�~��a�g�ȅa��	˟<�i��&\����J��'W�� ���B�
L�C7��z!�� C�i�r�'��I؟��I�2��c?A+t��>]y����c��;��\�v�v���O|�Sxh)������'��\c�N�1��ɟ#��ĳ$��L��4��D�O���M�7W>E�s�6t�Q�N�EY��+��ѧ b���V�i3剞P� ۴t����8��
��])�Tp�t���	@���+>i�6�'��A��>��)��g≝\іQ��$�?#�f,�f� ��6�� X3�	m��������������|ҷL�;x�	S'e̊81�{���OC�6SY��ӟt�I�?c����	<�%��)�-s����Phێ�M{��?���%+�Q��x�O
�'N ���d�<����AC�	a���>����?ّ�@o̓�?����?i��L:�M��E�06 @Ejĸ-����'i,ِ("�4�P�d�OR˓�B�h�x�0��f�@�c������iI�k�;�'c��'�b\��	�k@��pX2�	)���!��Z�m�4cI<a��?y�����O���� "rF�h�� �m��`;�d�q&��j����O����<��c����O!��N�_�ʙX3'�.7��!Kݴ�?����?Y�b�'�|I�vÊ7�M�Sהl���p��nޡ�ah}��'�r_����9~0}�O��k�9��p���*i� ��dՂ{07M�O��,���)�e���)���-)d B�#��U�� �S�!����'���ߟ��4�V�$�'{R�OKR�[e���d�s�9�|��S�!��	�,Sx lb��M}(�
�u �-��5j ^��'k�/?9r�'��'���R�֝�� 4Ң�.Mn�m�e\"^�\��?ѱ���W��<�~�3k^�~G&���$D-O2�za#�Ħ��	�֟��	� �	�?-����'�
x��/ҭM�i�5ē�D��7|�8���D��rE1O>1���H��a�Q��d4-�+K{�X���4�?����?�����4����O��	?6�|Dsn�" 8��7j̺:`2��y�����.���O
�Iw!�X��[���!�&2V�r�'g�a"�\��	ȟ��vܓya�x� 3�@����&m5T5A���>���3`�Ȕ�'G��'��ǟ4A-�m�LȀE�nƞ�xĚ7]�|��'O��'�"���O��1�`N���1��o�/}@U�E��vk�Q���<���@�'
¬*��邟5�����H^� A�L�4s�&�'���'��O��� ��24@�i� ��_�t&
1�
Z=&�0�s�O����O�˓�?	�m������Ot���e�8t���T�L�^�� �e�	C��?�u�W�-n�`%�\�@�V����ֈ'3��q��n����<���`��q�.���O��حKI�t���0���T�],H"���>q�qW@p�$n�C�S�TIr����q�ɰ0\I+�/C�����O�]�j�O��$�<i�'���岶�']|Pp�U"�5�hz�R���I�"�(S��,�)��Y���+��
oH�8��M�4^.6m^�B�����O���On�)�<ͧ�?�v$	�A�68{�_<w61H���~��F���R�	0�y��I�O~e���٨]�M9��T;����dE�����㟸��K�蔧�t�'r��Oec����"o����7f^"Ti��I�'r����d�O��ɱ_�pQ�fE�u;�$�J�G�$6�O4�XSN�<y���?����'by[����.~x�۷�%�	�H<�@��y~�'�2S����yI�Ac��:e�АqА)@V�������O��$�O�㟠��)�rɒb�V2� �RK��k���o��&����?i�����O���%�?�0�̙� ��DAE(FQPa뱪{Ӏ�$�O��$(�	ݟ�����6���J�rwg�h��8�(�\0�	���I|y��'ʂ�9]>��IZ�AP���B,��
p��9�b�ٴ�?9��'1^����ēl�� ��"�<nR��p��T��<lϟT�'����c����L�I�?�A� 9 FJ=���<b���x���'"�e2~�Ҋy�����TT0e������f8����R�,���(��!�	�d�	���SfyZw�x�*��W"]V��1B��*9�9íO��9m�3���)5F`�`�&��&��܃-ڵ2؛���k�"�'����?]���D�'���c ��V���Lp��`Y��&�͚'�,#�y��i�OhĠ3!�Z�������"� B����Iٟ��I H-�����'`R�O)�R#�b#L�*qU;$pX#�$O}�xf��C����'���O�Z�D	��/�k<	���iob%I�D������͟P�=�ge�&|�-s�یI,���	^}���.i ����O*��O���?�`��m�2�c����l�F5�5 Y.O��$�O��d;�	֟بԥ��HR�I*ڈB��Э1��ts�*/?Y���?�,O��$��<�l��9/���`b�h�0qģR.*��6��O\�$�OX� �	�)7� م!t�bp`$݄0�:��1%R�C\Pr�R�4�I�'��,C�T;��៬�C"`?���	<RU�gJ%�MK���'�"o�Xي�J<YA� 5=��a�vH��S�8lk�E�����iy��'"�9YgP>m�IƟ���j�:�kSꗁD���0�[�j6�x)�}�'�DE��A�����	�h�����M�#ph�Ц��f�����LA�D�(�I������?1��u� t{Ў��b[���S�L7N"`�_��	��D���4�)��6!���V&��0e�(B)�
J
6M�N�h�d�O:��O����<ͧ�?y�$C�VyS �T:��l�o�0���-�?k�:l��y���O�< @�j��� F�D�m)J$m��������I�r�锧�D�'��O@Q'O`@$p��{����[n�zDP�'���'���O�Ó�J L�c���� Q(��ij�q��	۟��	쟴�=���[d�t�y���BQ����.�z}r�Ɂy��q�O��$�O6��?�7F����ÖH�a����F���(O���O��d!�	ߟ���V, ���1�ؕp
:}Pf�FC��;��%?����?i-O��dNa;x����(����� L� �l#�6M�O~�d�O �h�	�q��qkt�x��A�@>�Ĩh&�N�/.�Tk2X�(�	��4�'�h����џH���6�HTx��T�Y[�P�%��M�����'��!U�Y����M<��jZ�MuH0H�J�Z�Ԉu�Ŧ��	\y��'O�%]>m��ԟ�Ӱ2+�5�B���h��g�}���}��' ��'�Ԟ�����ќt��D%��Wؖexq@´+���埔r��Ο�	ΟD�I�?���u�E'n����I
b`��;������Ot8�� �Yo1O��l4�B"�S�||!k݃i�l%���i�5&�'3��']��O��i>U��T�Թ���)-��\"�:d��u��4OS��Rj�i�S�OR�F�"��z��Ƅ}pceغ"*6��O����O��zd@�E���L�Ir?Y'	�M{x+��į]�������9�I˟���Y�.��Iɟ �Iǟ,�	��$��hɫaX�X�$��.X�6������M;�)�,2�i���'�2�'Rf맙~�`��eY������X�6�)ˉ��KR��$�<Y��?���?Y��������&�>`���B�8�`ňS���'6��'�r��~J.O��DQ�(�~Ir�
)
%4I��-6�"1��:O���O�,����OH�$�O2��{R�<o�/I�L�`DFX�q�ˣGa�I)޴�?���?����?�+O��$B�R��鎀YSD4�!��Z,Z�I�	_�T\�n�ȟ8��某��+��i�h#��mZ������F�)���DU�(R�]/ ��Zݴ�?y���?*O��D8g���OP�I�~��\9@ ՘�6����Bo�7m�Oj�$�O>�DF+L�(�mZ��d��ş���7q@�$DG�-�xP �CM0;h���4�?Q(O���O��i�O*��|n��{�q1e�17�sQc�@��6��O��D͖L!�m��\��֟����?m�I8Fn`%/*�Z�B"�܀\Cv��d�c}��' ��'Rɧ���~*��Fh;�Y;� Ƀ���ئa:�.C��M���?�����'�?����?�G���, �C���|�f�:փJbG�ƫԄup�|�Op�O���R�&0C���N��T�@�L�D7m�O��D�O`� 2�N覩����Iԟ��i��{�N7��iXGf�7�q���GuNm�o��<�OK���'��Nz���A%4]�k��/\/�)5�z���$JB"�n�˟�Iޟ��	9��)������,4���ЛU��i���>��Q~��'y��'�b�'iB��/<?���$�5\0��y����2h�s������O����O���O9��` �����B(� ��]���Ѳ|X��?q���?Y���?	���5'h����!ҧ4ւ�(�k�,Y)
��w&
��MK��?����?����D�O<��p0�$��Ԣ�
K��`��
��Y�遀�bӂ�O��d�O���BC�4c�,P�6��O>��Ί7.�B�&��x�tx��l�Xl������ΟD�'�B� '��D�'.��F#x���I���^=�a��C�?����'#��'<��MA�7�On���OH�	\6o��9��R�<�T��)T�!�nZџ��'�2�D�O�i�\\�7�ٍD����#Ӭ�Hi�4�?��T+�X��i��'>��O����'h�՘@�(�n�+�πv?�+�ͫ>���@�(������|�I?*vnU�5� @H� �)#J�bVed�t�#E�Ħ��ʟt���?�Пt�	՟|[uɕ��l�9կ;q����C��M�����?y����4�������\s��d������Yk�)D�+�$mZϟ�������$�(�M���?���?��Ӻ3�O͚L�G�C.z�"�Q�����	Sy�ѻ�yʟH��ON��O�"oP-��hޚc�����V6j�<oZ���!j����$�<������Ok$�>!��F]Z9XC:
T�ɉg��I۟X�Iܟ4��런��ş���-��`�#A*=bq��+G,t���ڴ�?q���?��PX�SLy��'�~�)�F��$
�������y��'��$^���'�imf���47&�����2��|��B��^j���G�i���'���'��U���I�U��擔Upb��5[�NH�����6,զ`H�4�?�/֖�?�������QԨ|��4�?���3��XW,@4R��r@PR�b�i���'S�U�,�� u�B�Sן��v�,�S!�ȍg�4� '��l�0�n����p��3���ߴ�?����?�'C�h��(F�J"2��2�9a��i�V����53?�P�'S�i>7?F}]������E�]��	ٴ��u!R�nZ���I�O@�)�n~��;@�J8��Z)V�U��Մ�Ms���?�=�?�H>!���0(�.uR�� �[m�<	�8�M�V�&%��'N�'��$K=��1(	��ƇZ�%d�Y���ߴbo*@C��䓃�Of"d�/^\ h���6�}RM�u�6��O4��OJ�"D�Q�����e?� (�T�4_"Es$�Ή%J�9���d�(d���O�d�O`��ǾGf*PR��-�D���V�9e�n�ş�����6���?i������jƘ`�x�B���u�R�Zg}"��2kB]���	���Iuyr�D�I�X���C��86h9�4�Um%���5��O���+���O��$�"5�Vt�F�Q�,`���^�z�5��M�OX��?����?i-Oġ�ċ��|2C*O�X��j����G6V1k& �k}��'t��|��'uRb/�y�R�@�|Y�K���Qc�i�bw���?����?�+OT� �b�p�Ӑ13��a2EG�`�Ũ��k�4�Zٴ�?�L>y��?�b�� ��'��<�v*�#)��ŀ�˒e�s�4�?i���D�-c~�]'>5���?}�-��/���i'�D�'� Ds�#����?��l�|y͓��S�T��>e�ȫ�L�����4�Q6�M�/Ot�Y�,��]�������u�'�~�+7�\-H"��iR!ðLV@Xٴ�?��Ic��Dx��T�ʌ7�Zq��(*�( DI��M�f��(Bm�f�'2�'���-�$�O����X����T�CI��u ����2$�P��t$�"|�ol)�UGQ�`<�!��8�����i��'3R��>�Ob���O,��A.	{���ui�d�戎8**�6�(�$\:/�?�����P�	�K킵q�G�3FN����nb��ڴ�?��C�f��'l��'�ɧ5��[�gk����{��%�ъ���MC�V[n=�������O
��Oʓ~]�t��=���R�M�h/B�'D��f��'��'��'��'��s��V�݆1�A�O�8c�9��%�y�]�X�	���'?=���TJ��=�NpHG"Z�7
����׻����O��=����'E2�?y�G[� ]Zy�D�ȶh\I�� \�yc��'�2�'"_�� �ڸ���#�"�-N���ٲ��;�Zu37˃ɦ�E{��'f�)��'��':�F�	�-\ a�0��ǏG1p���n�����IƟ���	v&��O��'3�4`�
KX\�RAP&{ԍCA��6@(O����O2�P���Fģ]�BkR�3�Բ|}���p�Sᦱ�	ʟ�`�I���p��������?E�I��֘/Np�mJ�9dt���%�H6-�O�DR�Y޶�b?��rR�˂�)RK�=q��Ni*�.Mp�'�B�'k��O���'��S
H�i(U�^���\т˃/u�\T)ߴKA��Gx����O����! W��h���T]A�P$N˦��I��8��=ls�drI<ͧ�?��= ��"�Z":)��@ěiئ�HWR�������	,���8��🔀L�bh����ؔ�j�����MC��-Xt$��x�O��'��bNތ�!�Q4�*P+�I[�u���kڴ�?a���_̓P>�3�΁QsعJ��G8F��E˭;�hhrBݚ!�޸�t��Pc�,�`�E-��I��b��U��c�w�'`���G' B�D	�T����I����8}wDNբLN�m��ݐs��s�G�C`���?b��dI A���q�S�lL�P[c��6/R�TQE �*�ej�� �
�RabF>&>,y� G���PC�bE�zqq���L0���� �O�B2�/��E5����NV"3q��i��q�U�X�-a���^0�
�q�$�X> �/W=x41��?���y��zr��7�J��$�>�O����΃�L�yk'ƙH���dK
@�P���6��nZ�#���129�V1�%�ԙ�2��*.��5#�割��d�O��?р�i��+�Δ�-ͣZ��páj{����	=��p�X YQ�CZL����D	g��4lҺu�3�ӂ�B�-���x�I:J��p�4�?)����醺/��$�Of��A�o*�`�2LO�"�h��s�8��ed�?�<�㏌�P X1���"�����w�$��4��%E���	�䍮�0U�e��W��cgKri*T{�(��Y��t��֥|�^)�O?�N�./��(�A	tc^pB�&i�$��b��O@E%�"~�ɍR����Ī^>�� ��0�"C䉂_�|hC�!�:����� ��"<�3�i>-�I(�Єۧ��� ��|��o�b�������pSS�o��X�IП�	�`�[w�w�n,�`ʇ�2�E�*'_r	`��O�t��ǎ41>X-2��������ў�(�d�	(���E�j���DD�k%�!��I��u�R����hO ;Ԅ
�_{�X�l��1�@L9��Ov��S�'��Dy�F�,do.�C㗄3�|��=�y��9�+� �8c�N^#fд#=�'�?!-OJ�cE馱�#�6z8�G(�!U���5��P�	�\��89����	џ��'}bN)� .ܰb�ݫ���x*��#�+|�l�8�i��]����TɄ5AVoO�n�*�{6nD�aT�L�,]&u�c�P�F�"ϓ%����t�1홊6:��S��p�����Bz�'�џ� t
��-x����B��9���5D��{���K �`�+��0�q&r��޴�?I+OJl��H����џ��O�uHf��)|l�T��'�-n��XW*Ib�b�'�'@�C�����l\5Nf.Ы�$��D�l�\p����NX�Ƈ���|Gy2lǬ^��Л��rӄ�6(��Ks�Q�
��w��[�1X`긊7��9j�"/-��'2P���a)�>�ɧ⏧6���rE�Z�-��!+ë5D�� v��ď�O��Q)��̌'�Z��d���G{�O��O���@B�;�l��r(�.@`���9OȺ�Gܦ���埸�O
j%P��'���'ʆ��EK>�HV艡y,�9��@�f=�v��/6���0Uǂ�M�OJ1��J��,��K���]���Q�,K�ZT���ضP��Фn��'d�d�g,�G�Ͽ{v.J�U|i��d�� �V���g��z��%Oɧ��B� +q�0UZ��^5x��@��nͬ�ybJ\�%��8�δZtĕ�uK��O�Gz�O�"i�?��E����Kp�Y�\���'�P��e�US���'���'z֝�杮]�%Acϕ�h9J)�����(��m��i9�P�K05V@
4TmF{Bn��y(��Нc9HM{��/k���m�5�ɓ0*C�P����E۟ўC@jJ>��SwLȅ7,QbuA��Ĩwo�O���+�D�O��D�<�F�W޸�YG)^s2��B�Xg�<	��.�f��f�(]��]���
O����Sן��'B8xٰ�k�n!b��<U�.`���Zv2�q���O ��Oh��T/)�z�D�O`�Ӆm���!j�	2[<��ʂ	(U����Bd
к�珺����_\�'��!C+S�6t���Ǝ|�˥�?m�0��ÂKǪ���Z�jNXt"��y����=�0�����0޴S~���g�4g��|���ثi����}�����"JR¥Q�jR�:�ńȓop��E�:�L�R�Xb^����V�|A�F7��O��d�|�V&�0P�W"X�@X�� D]�v���Y���?	�
�IjЗ��p�D��G?�m�CR?EK�	D�4>��C7�7����"ʓID��J��*lJ���z9����`�XF=���ӯe�.��	����	H�O�V41�eY�M��y�&��b��h
�'��<� �I%p+0��r��R�II
�\ډ'����)T�F9Sr��a;�'®��EI�>����iC%QG����Oh�TR���`,cd�B��FzB`Y8��77w��j4䎳Gln�����ؘϿ{��jt���p�ύp`IT�'Y<���A�'7�\ ����ڱ��j i�Ao��+i���Z�j�e��qfD`�Q�=�|����/^��d�O����OT"~�	p�F�瓀r�6ԳUO׽I>��I۟x���;�V�������qMՅm��b���	:�HO l���O�`�vfA<fH�򩅋P�0� 'e�OD�DZ��4��W(�Of�d�O����˺����?���>~?��3�*x"�4�'�^Q?�#F��9��A�s�'��<y���+��u��W=K�Ȩ4oVg?�*�&�ᑹϰ<Y�4�<�H����F0�4ʧ/Gg?�	Fß(�	�T3h��PݾF��tÖ�؄��?9��\���9���J�n���������Sn�	;\Ũ��4p(�3��E�x��Ɋg�_����?����?�A��?a����gs��DèQuv��&�C�(��MrFR�v�2��ɉ~e��QE�nLh��A��	����2V)l�<qH�&��p<�F#�ٟ��ܴ	�͡5��%zx0�Fƕ,:�(�ȓn��A���y�(�bfJ_�����ȓ�Te��kV
Q�\!"�
	\��,�1@�6�|K��Qh�6-�O���|� �Z�sȼXz�=�!s��+'�b���?��:�	SrB<D�fX��G)�ܽ�c�?�!��H�aq���+�%<)�&�3ʓI]�i �G�EB����"M��;e��+<n@6��?+���V��,�t��w�P���ܛ�
�OrQE���¼6�(�wGQ�s���тD�yb��63��](���*hj�ݘB!��0>�t�x��U�}��ĨmJ�*�J�[�*
��y$A� ޤ6��O ���|bg���?���?�v]"e���#Laj昂�O	f �s���Uɧ�I(��O:!��g�*�8��T�ˈeB<h���/���@^ OpZ�b�o虡� ;���U�f%%.�HQ0ǂҩr�;ƃ]�lR�@�	��S��?� h�
qh�T����ӖL�{�<!J	f�< �>@@ Y!�#<�v�i>��I@ۦ�z�]<h<xrm 0!~����H� �E�,��ߟd����0pZw
�w%2�`7~�c׮T��\5��'WfA
� �"	�慇�+����׊.�����S�̈́��0{څ�p�)I�.r�"��B�	�y�F�d+|O�{s�؋��ل�F�{4�ã"O�!��g�	f60D��F��244A2��}���P0[w�\¦Q�IG$=�]�f�ʇ[CV�� bKş��I��<�	"m~�x�Iɟt�'x,����B��f�4����9P��1�@�,1|Td���G9ay2����#���QRLR|8�Rf�B&p�4��H1<�K�B@=`l�Dl6~��3Q�&L�X*M��f"�OH�m�+v0�ZG�E,!��@�ǭT)B�	:"��9�+��NԘ���ǋ
J8C�)�  ���`Ӟ&�\�����Y2x�q8O�n�K�	�jO`�)ܴ�?	����)^+*�`	���;gC�1��I4F���Al�O��$�O�X�.����,fy*�HQ0t.��2��X��bNap��	��		7�Q w,�: �T���dNY@EA�ܺ��͐�_1��P��w������[�'ָ��]0�>-I� S	~9�<H��	i}�xi��(D��"��H&��ckZ�[���S�'.�OQ�p�:MD��#���v�^��69O��z E��]��̟�OB��a�'%��'sP�p���u�~��N�7x����3�Ȟ?SJYXF.��
ĂvL  ��ŘϿ���=����n̛fS�������K�Π��)F�n���E�G22b�(�7��﮵Y�oW����d�� ���暚W�~�D�a�)�矜r+�/�A��3���DO1D����_<LqT)��
L\�6o"�#���S�����ʼ:Z�����&N>�Fb�����I�2d:�R'A���$���T�	��u���y��փZP0��ʄ�{��uqwy���͈/�L��4�.��$��hO�"�̀��9{�'#���^0q�ܐ*����7���r1��%kr�)9��c����i�/6Zp��C�=�������O���䟎U}.�G�D�e�j|�C�<!�d��#�,�'jŜz�
�pb�p���Gz�O[�'���bӈ5���'R��S,���0����O����OR���!�����O8�S	3���{1
Ԛ��=y���1'�R�6�L�B'h�0�0=p��
s��a0�ɷ6���"$��� �l�*��/�B9���R�!���A�'��U>�M���H��b1��!Î����#�Ċ�"����nV�=�Z%��G-D���B��$��Y��Tlq����!-D�P
R A0"���K[�h�bBi�|K޴��<�>����i�r�'��S�el �+f��!�*%8��Ɓ>O��q ������Iڟ\��V^z eՄ�* �S�� �%0F9*0<����(���(O�i���5_��B"(ٸ<�|�qʇ��=�n(z�k@�B��H-�(O�8��'��#}zP �����*̒=
�(��y�<)��^	��[��	=�^PycnIw�zH<�WC\�l)�@�/�:�2"D�<9���H�&�'{b^>�b�C�̟0��柈�RgL_z��W�*�,�ZQ��,T���� O%hx��k/'�pm�!џ�b>��Ɓ4"zq�Rd�)�ty�йS�j 1�$6P8�ɛ*=@��m���u�B�5՜dB�Z>��#aR~��A�'t��A�B"u��$2&e�O�b�"~��$�dR�NǼ(��(J2b�>E�6C�I�H�p�cq"�=gv܌�S�l;@b�<��;�HO�	�O�:�o�!?��"� �+}��ȉ�!�O8���jQƬ1���O��d�O������Ӽ�A�{�l��Bm� 9d]c��=1���$˗�v,����5
z��'n�Q�̲�cA�' �ĸ�+	/?� ��j�$1Q�dڳ�	҆��"@M��:��7)�\���8�Iт���E��|^���v��M&X��.-�$�D�w؞lۑ��=gxX�qc�ja�y�!D�؂j��P���шU�l0���f@��HO��0���>YpEl�3i�@���
�c���$K�o�(�I�T�	����,��0�I�|j�m�8ꔌڥ��
y<xSe�V>z
EXE�S1*b��a��g��A��	�L�RqQ ��=T(���<Q��!MC�.xP�@�GP��@�"b��M�WC�sjj8QJ>�wCNݟP��;!�B�ȱ.��y�����☁<�0�&����ş��?�O�x#��V,'8����
@\�ހY��hOL��@iD'�A� U���|�8O��o󟄗'�"�t�`;a�'��T>qi@J�>M��,�c��9gx�TS�d�N��IП�I�6�&@��D%{��и��ٳU3"���pY��1�˓ݖD�F ]?�Q��
2nΕJy�!�pȆ��\�b�#�ʐ�bӪ-��@�!O�J�"jp��4&T�)KA��*�R�$ҧp�H�I�tz�S�'��h���ȓm��%��M�[�"����g����	?�ē#4�8�"��|�Vq‘�k�,=�T'���W�iD��'s�S�(���I����I�:� Ȱ㦉�i�\�q�-}��Q��; �Шn� �hi+�S����'���;@�Љ�l0�pӞvdy�	�5�
%��
�*6�iȁ��O?���6uk�N5��(E�ϕT���#M��?-�ɧ����W0��`1e��1�&��F�6�y�AЅo�v�Uj��|��� D!�O�}Gz�OBhO�ɘ� CC2[6p����3��'��XG� o���'���'4����������X�=*EF�1=p�I)�^����2u��Ȩ�n��=2���.����B��}r
��C�JP U$3 ���PH��~"��?���'i�p��2�R�H7��P����ʓY^�)�Eg��a?8��b&?ָa�)§$$������ � C)D+���1��!�P��"
�O����O����������O��S"���+q�ґ���
�*�%O<vIe ��q����D���V����EZ
��O�0�)Լv�<!+w+��b��!o�5�ZHjT�.������-��R�ɋ$�$�{�Œ��?!��ivj��/�\� m
3��<|�V)B�'B����9CP= �ŅG@�]�'��Y@�n&Y�(Y
ׄ�(1�Y��'�6�5�dA7*�0�m��d�	w�ć#Y�I���A�i"D�"G��h@bA�!�'"�'T4��E"֯-7���e�[B�HC�c�Krv!�
&���K�S'���"ф@r�'
֔Ruaj�
��M8v�μ�@���u7&��l4�+	)U�i��$h�h9���]�Kb�'�`9���Cc�>sw�[�X0g'V�D�@t��� D����Mٞc*�Cb��;���T�>?���4�%&��Rs��82��P�Y�V��ŀ��}��)�$Q=�M���?i-������Ox�D�O���b�<"�M� �Е?�䣗͓�OC�!��ө5���I�a�ʧ���?e�Jq��sᘪZÎai$��Q5�u0W�O�cf�6���y���'�b�qr,�,[��D�ަ8�3ao�'`RKh�T�o���G��d���󆞆2<4z'�3�\�̓�?A
�@|�a��J��nE��C�R0F]Dx��9ғ]0"��:�<85C!^���&-��f�ܑ��ğ��
��h���۟���ş��^w$R�'�`1S�N/:M�|z�C��]B�'��aH	�$���*Ǉ�<[�&��T�� K�Y���>I��ɿ]'<�1.�(l%�TI^"C���ɏs@��d؞`�V$��uB�h;Bn�(y����e=D����"��nI��# *�k �M��Z��HO>ᙆ�ת�M��D�9�@��(�*���г�?����?q�FŶ	����?�O��MCWl�"��ׇ֫ն�L�L*�A�C�o���RoR�Q���Ey��2n��L�J��珊A"	{A��'����N�@��F�-'&\<��/M��')���A���H���N0����,#F%ȹ�y�O\�/�9���1�eb���>�y���2��� ��S��������y��e��O��+���˦��I����Os�H��l{���q&{\V���䑳?���'� j+��q�@{�:���H>M%�!�'q$�Q.�7����G֎�ȡFy�o1C�,P����4�< �@��� %��FB�Tᮘ)K��l32��	T��(��DE�NPe����H�B�ȴ��e��Y��X�?f��&"O��""A�_��8���=q�N�j��'�OZ�V�\�&vZQ���"�X��:O�<��T��I�	��H�O�"�	3�'���'�r1��|�ޕz�B�3�^q �߈}>����MS2Z��|�����=}t��B�8�����1#��pأ�����5�PU��0�2"�������"�^-���Ⴄ��19v� �'>1O?���
Uڭ���?���{�!
|!�d�=�qgRe�<�����pp1O�Q�����'n�s��8�j%	���:٢m���'����]!����'c��'�R.v�u�iޱ�7/�0`T�����@u�tC���h�J�VӤx� ��yH��~I�xc��Y�[ĮD���-�~rbV;;�R�c�/��<-5�� �hޱdx�,�ǃ�6?�I�E�T�$�O�O\�$�O$�x��@�CM��b�pB�/ U� ̇�$�$ģ��]�5�<��m^�E���IT�4R������M;��_�Ieqa(�p�"\� F
�?����?���ؐh��?y�O��� 	�d6"���/M,�Y�4'1_����̈́�$�
�����x=N"?� @J,nJ���H��n�IѦ֊Xe>�I��O$J�q�!)ڐ.�-,s~h��\�qO:�q�'�R)L�i����Ρ$d ٰS��yRl�?`t5+���K�������y"���E�U�O�c@P;׾A��æ�'�xC歘9�M����?I-��5��P	\n(Q�$!2EI� �4|���Ob�D�ce8!1 ��eN���D"V�7^��p�O�����h�f��|�Ь�&>Z�(��DM����� �ىQ�ȼy�ʃ�W�@��T�8���#�7��x��yPģR(��eH0��H>�(�՟��)�U��]�c��:�Ÿ�J՝q�!�$�(S3�p6啀7��p�ש^&���i���h<񄏄��Gk�.Z�@�	�9M����n�
4n���l��O�t#I�+���'r�Ú%��es�G0)���a68ײ8���= ����Џ�F9����C2����g��13�E�z�l��l%G�=yf�(Z���$G��k��Q:�ғw�n���BԻ@uP���g ��/���`�	@~����="\��'���O?�$�~ELG+�V�)�$Y�m?!򤇪j�R���IY6}��ePf)�&^8��+��4�x��,���W�_�@�.�{��U\)L���O6)�����Z���O�d�O2į;�?�{�? R䢀���#������m�x�v���>[��z�o�j{�����M-X	�)J�'��(�EW�b�<�i0$"a�]���¨8YYA��]�|�vƗ?����J�U��S��k~�.<����plֳ.#l�`%�Z$�~RDǇ�?�s�'��M�E��3��"d�$;�e��"O���oьCa�ѳPI��s䤨��O�����|���Qք7-���v��+ײ)��HK�1Pw����O4�D�O��g�O��D>U2D	F n2n�2S�V���-�#P#�� �8H̆��*��k\��Ȍ�$�F���5�`_��s'H�>��\�Pj�\���&#�'D�M�c��8:�P�PfH�#ٸ'�H(���Fh,R�T2¨�9|�~���&��y�.�z)D��O�:	����P���yb'�>,��-z���}N�فh��yrb�P�O�Xߨ�M��?I.��H�懈�vuZHP������%As����O���	I�\j�AE-OU��1�O�/pR8��O�<�0-� I'2'���;�� ��$�V�t��ˇ�~AV��t��(�"��;>��A�	]Ke���0->8���+֓-�-(O>W�ҟ8"��	�Sᢵ��	��! �Jr�V�!�ԵW��2�^��\j�b������/�]2<�jP9t�ם|����b0MJ�],�b�m�ڟ��Iu��.J�cb�'���W���I���:{r�a6��N8��fN�p�B�L��'՘�?q�L�f��h�M^�Y����aL"�61�c�UB�<%���D�Wg�S���'�L(�(��]�����쑨D�`��D딁��&~Ӷ8�����'�(�@��B5x�D��0-":�d���'Lb�'�$03*P�O6��3�䟥5#��Q���[O�'�)c6��&[�5M���f��k[������@�gڼ]0��	��P�	П<�[w=��'1�8����N!s���:rܜ�b���:#RL��:s��"�J�1��t�.� �DX�1E]�&��rW��6P@K�*��	g�XPe�/]��Az��m�P(H#�9�k<?Q�R�&p�#E��0�$M�j�s?	��� *ۓO��%�H_��jǡ/BhY��6y�T��P�
����+A�b�8�d�i>�E{��	%�*������Q>�Q1��ʳ�yj7� �iw�	%E���a���y�@��~/6y�LP?E\��U�'�yb)��r��vHJ�Lk0�A��C	�ybl]�:�l�k�6?:$ Ƞ�X!�yM�8?�T!e�ȿB�����y��-<3�1�L��q�ֵ`�G���yB�Kp��J�'X�t$I'ڹ�yb������
�<nf�Za � �y2@W�k��y1��t�xP&���yr���.��{e M�p�M�D\�y"*��@L*�`�M�8]P�(XԢZ��y����t���QE\=&]�4�.�y��#
�D�r��i p`SF��y¢��K�li4nT�t�l��b�R��yrA	�B���@EmR`};�kK0�y�aB�T�t����v�Ɛ�A	�y�mY{��1 �I:�L�r�@�6�y���`����w�U1�|��W��y��N�r����n�
-�����aı�yR�@�4���� �ܵ(�Nqj�kJ��y�!�Ab4���Ǚ8S��yF�C'�yRBđD�~����X��O��yB@���r/�io��I煓-�y�jK&u>��8�U�N=�Qjq�Z��y2�FĬ����NQ��k X�yB.6_��	�	ܓv���0��.�y��J<�vM��^4R��K��y"�O�3$���*qf�z�D��y2/�;�BH	!	�������yB*оs.PpQ�M����hq�ݲ�yQ�u{����'1�0Y�ЌX�y��]����J{�@"��κ�y�N� I���"�)t �[Ϙ��y"��"ʥ���"tT���T6�y2��^�,��pΊ~�hq`�R�����Kg����'&� �#��Y�� �q�B�(K�Fe��k��M��"O�u�C�H-2�ډI���%�Ā��\�xT�� g���$�,@ZFA�)�Ȣ?	���Ky�ИR�#t��H��z��L�� �$�rJM�^���4�Ó.��x�������4�Z��:=��ɺC	�!sa E
zK�D[�)Z�C�@c�DY�!J�JP�9��W�P����]T���JE��7F��à�<K6C䉳|?�q ��/��1��'M��s�%b�\HjtJ� _��y�Ԭ,�s���I�_~v���J��1r���C���c9=~P�pW=� 8p$�MX��,Y����'���Y[�����W�I�X�a�Ø�=�ڹ�1e�*���OF��S��ݮiST���O����	�#%F���������$�p<I�C3B�pi�' ��pxtE�	�d��(�7�D*;Y����D?�pM��)�R�˦�i>���$^��4 ��8���C�J 9������h�y����
�"��S*<d��O?e��$�*���Lw���큟��'}�<�wH#(�TT:s+�Bn�N����ф'�,��狊N~PjbY�Lz6�hy�����f����-��a��=O8q��X�!)��	�x������H�tY������Qȳ�N�oa�e"EA�5�p<A��Aް����b���$*$�8 �'�5�@t���B	�"kP�!��OX�?ARs�k���+�Z��Cf4{]Ĉq� ܰM����Ǔ1P�t'�"0C&�!��c�ܓ1�|�09��	�D�����Q����h���	Ԁ�k��o:�r��2p	
�s�i�;�h�"K�	n�8{1�N8d1�`��y2�^$��a�U��
v9$���B��W���OF�{�M�n~.l`�l�-ak�=Y������f��Ħ-�l�cC�!`���r]�]�D
�2J���OP�q�,�K. M��S�(���8IB��`
�6{���2ᄂ�*���W���'�u�J�� ��@ ���.�T��#���5&f��:d�X':��)3FB�_8�D��O:9��g(:l�`�+�D�\���G��A3�3O2İB'�q���O��XA��#-Г>�Ru1q�n>�:���!bQ���'x\}�q�ŵL�%:�BI&t��
��m[D��fc���y�lߋt�
a^_���c��r%�Dߴ���vR1��qmZ)ˀ��Qߨ���#X<�QѤ�NC��t�
Պ+�P��1l��jRa����NG�7�^Ȱ��1eMVdX��_;S�d�87��Mc&�ȈCL�)��ּ�eN&B���L��:'��%󜴳�B�7if�s'�d����l��2^@	�"��,;nĜ�q4O�8k��<�cFͫO�%�$P�0 H�/�0!��p�D*LɢABa� u�-Q��$���DS��9R�����}yi�'�Q2Q���<��ڵ�D'=�#��_����M3Q�Դ��U�elM�BD���a��C�JL��,�X;��w}⥩F��3nX�P����`�00;OL���
!��9�0W,G;��Ʊi��	F#����S�tU(	���=)G�Ii�*_6�V�2v�0ғK��ir玴cc�5y�'-/+t�'����C߾0�B���(�%�6�hujѸX5��K۴tx%�ī�$_%^����=ᰤJ��@���?@��%��Q�*����� �6�(^>D�3�L�>��dk�����D���lܣ��4.�:��JE�i��R!	)�xa��R�(DU�")@�o���p�
|9���X��,PU �F����ɇ���I����$F*��7 8D5����o*��É�+�$��O�;B����� #�쩸����D��v'�_�p �eO�;�F�Ce�/��e���#nŽ5\�����^�t�6��Ԍ�3���?���%�]B���$�+-���@vX5�HO�X��
ÅF!^dr�6$mp!�T�l��ǍY���,V�F��4�Äx�n���mӒ�jS(U�"��A���[3��,I�vR�'"���EJ	�5�� ��X�o��0�޴p=H(��2 ��I�%B6&�Di��Γш|Q%%]�]�t��U�!X���4O�T����G�M�1�房
{�=C�� O�1Sm�+HR���A�Y�𼺵_1s�f��'�dl�x��u�u��.PPcC�48�~�m��*5X�)4FA;��C=&z���V��q�0ӧ���	���W�� �O;����P��<9��ATP�T�C�ˋ-��@����S'{����'09.�����
s�Z����<+����o�g�'�V���j ,���Z�ϗ=[>�S޴���SDZ���A�jYM��8�!HTplښ8�J'A�>S����(J<����P��)zR�iX��3(�h��َ��ɂp��@�CÈ6@Nv�2��ix4���ybdV+P\��F��W��jfE��+�@yXs���3\8�3!�_�"����V��u7*i��7=�k��2���"�@J k�y�����6Jp�"�"���yF<)#�)v���b@Ko�7��&�IB��=M6Pd+l	��4:�dB��>ip���Ȑ��Ľu���3JD� Ѩ�*�&�E��&��J,
�|"'$��&qIB�/yL1J��X�$�lD|�(�n)�A��-�	���섍�?�r���V�P\�r�Qک0P����h)O�Dl��J��mΧ��u;uN��hmT�'�`c�ZYzDURcƋ�K�@�'���ODu��p�Z`a�S�<�dG4V��\�bh��oNI�C�N���Aa��l�Y��鄤]�����3th֔���'�(""��g�0A�n]����Rb��O1�Pm�c���W�<��f��."���e�6~f�|2�߷e[k��$g?象,�W�L��wDΥ#L|L�>�w�3��'&`�9����24n����kC���
\���O�l�� �xlJthE#�x����'����J�K��ݳpHV_-�=9"�ج��'�$"}�'j���n�@����p��2�'z����h��PsoLC�j��t�O�f�Kɇ=��2"!]�����Wj��+1�}��)� �m0T�K������M�0�ʰx�e�&��ES�+\>ܥ
������"eBȘ�!RAG��FĔ~ʰ���I%��+J�(-�L4����gd��q!������F�T�oO�0{Bn�]�b�{����ڒ�JٹA](��MxFkY�"/�\Y��B	{W �	!ʁ�IOh,	Wܟܼ�nL6�~9�$�@�@��q�w����'r�么��i��I�K`Hȱ��*W@1�.��\�KR�e}�Q��4y���O��9v�x������-�	[�ĄӁɨ_切�E�ˏ�p?1ЉǠ<�d��a	�=��]9`�0Cx�'�vh��']�ɥ@�
Z��ٷG˕C� �;<6��H�Se\icT�
P� �ȓ"����b	�b��)���M�lS��k�<��GIn�e�p��~�J?e�t�\1U`�9 �)+(륚=`��`bWcä�0=�Q��0�'�2��RObe��%ئ0����jB���nڃxrq�!\�|4��T"Ӵ2�J<���DO�|ձre	���ȑb�ķgqO�I3S�˦s����'����'�>L{'��*z�ܐ�<hΡ0���gŒb"��-9a>��B�*Cz���:Ehp�a�{.�����݁^�.�T�� W�&��ɚ�\<�s�a�x)2ui�?������͡��D�ܬJ�bUC� `p���5[!�d�	k��!ygj��Nz�(5N�V��)�S�F!�!�ł'�Q�Fi�i2��.-����5f%��C��S�Ϙ�52Z�x�(n��DV+Z����"�?Y֫�&x�� �U�L`~�A[֯�6\�$8�"�T�����ch
�%}�m��B�n�H���cпs@>�1�L�#Ae�L)5��N��9�;#H�9P�x�'W2�����vTRB��(ں!H�0F@���Ňӓr�x1�MJDi+��?lv�����56,�>b���ѷa�VJv`�-�2���(-�� R�AB���L�24�&��}"r� �-@���;� \V ���<	�,կ7��@� ��i�B�-ɋJ��HgGC*���(VAY�5��y������W�J���@����Ӕ� �R�d�d�^)�b�J�X��=�sk�G���Zգ	Z��d��i��W3t�,T��
�'�n�O����%"l���'���O)�y A�R�}{�X#��W�Z"h���'P�,�۳��B�~��!�D��BP�� ��	
kX��k� 7���Hzh����E�<1�O��T�P���9j����o��4�D�y�u��m�7N�i�Tň�P}��3��H�)Zx� C \Ok��5�*�-C�Y�*\�u
��2�6�^�J�E�CI�/�΁QU"�#jui����u�(�������"X9�6�:#T�Ч˳��<q�e�0�41�"�^�#��� R�r�)���VU���B�=a���!����?��ɏj4 ��=��(���F7f�	�\8�"�)ـ?t�-�덁?Hּ��
[:~>�'���{���0tlYt���!v�3�'X`I��W�?�� �X�+���%��w"�+��V�) �0��h�Rz�)ҚB�j���@�K3J��?����a��ʃ�K+D��sP��$:G(aX�g^�x0��@@9O(l����ʇ�S$�l�rR����Q��A��˶����гP͝1Z%:H���,;*��i��bGS2�6p�V����1R�o��H
&`�JVz�9³i>T���X�u?O��E>	��YtG�Fe�e+�!Y�-�(��
� �ى��R�FӀp��Mu� ��oAJ^��s��aY��;d�ߐ��I8
ތ�w�����9`��Ox<�:F��p��Y�B���|�Üx�!��S���``��%O O�y�����x��=$��J�GEU{�R��f�'�-��N�L���zF���{�Ak���ډM�	�s���2ʤذ�'����P��z�m*�Dz�PR��ʩ��D����:2��`�˺ S�$�g��,ymz E#Ԓ�p=��HF�M��: �)+0��Cv@�`�&;C� �J��F+x�8�i7}��2aV���?�f�|��8V	O!J>�S��JX��1t��l�{"�=PjR�
d�V<�	�23ȵi�k�)V5�q�Of�i�d�&,��D"�'!
H��\1 Mڬ�3�*T�'��[�oD �@�lP#m�b�)�Y{ܧb ����^F���B��A1���(hًql�$c(O�}	g�3?��N� -/�yȅ���[�6�
�lԉ~m�	��J���*)�Af�@MF��~�L� �4&H�L��H*���?<yr`� cゥ�P���rz����i��9��L =��=��	��pyJ3�ѹc��w�ΣX��
����S򓃳?����kd� ����Yt����D֨@�*��u#ѹ���񫂢V� ���/���el	}T�h5}��2tz�
�'XD�>��̩���2Y�d��8���$��}iY�,^�!�ʉX�Ĩ$`D�Z��4`d��{�K�9ς�$�ΊX��`C�Ɋ��剀{�b"|�']"̋w�J>Y&J� � �?sZm��-Ҝ8w��a�- ��3��������	?80\�;7���9 B$jN)�$���3H(�*,�O�1�5K�;
�uP�'�/'O�;F"O^�ek{ �Ȫvl�$J8x��"Ol03�BO�.Z
�C�	�~v(Y "O΀�Ak�"� ����ȶ ��]��"Ol��mڏp�Hӧ�m����"O�¶�n���j�d[�I�愋�"O��-F��5�^�;o���"O��W�ѡ$5��Þ���y�"O� �b�7���{�7}d}�g"O`mJ�;-�z8b��٨Y��� 4"O����o�E����8�v��"O���g.Z�	�����o����pHG"O��j�jC��pZ��ë:\|y�c"O���w����M���-8[� �"O�2��-�%��A1&L��y� �@�gĀ��tZpg �y� CCԐ��nR~��3�3�y���'�BQSa˟�{��Q�N��y�.��<(��95��}-�mk�MK�y��4�$Q�"M5`BV��G���y�oבe 
�;"h�Y���붠E��y��ZS%��h��ZIo��7���y�L�%3;�T�ē�
���X�I��y��0	��U�V�7Oݒ�X�b1�y�	Z�`�sVi�<���%B��y�� #݊ԫg���{8i���	�y���;f��G����DG"���yB�M�5%� ���	�L�j���y��)h EIY�򝒰�1�y����ڡ �lQ�iy�@Y�϶�yB�8"ԌAA�H�7�$,� .���y��T(=�  ���H�)����Þ�y2�[��,�zQ�N=JlX#�f�*�y� =s�i:�Z>>Ȣ7KP!�8D2�B#〥X|P�3u �l!�ā[ҩI��I�H�ҨpP`6~!�d^�G,zp13�h��L�DW�)�!��\�fz6}Q����"�HIqf/�*X�!�$��ldq��$w3.�S���&g!��	�
M�@!�4P9�(v��e�!��66D ��o�:�	��!�D�2���V�-�����N{!�Č.&��CWmĐc�b���48�!�K�L���4�� ����I˅Q�!�d_���Dz�(�0hB��q�,:!�D<v�V��0[C2~�3�H�L8!�$\l�!�E��f.j��dEV;6!�D�(Y��]�1i^�9>�E�dW)5!��&����IH�h�&�͆4!�DD$�v�ZC��]^H�C�i�	�!�B�	�c[�@I =ۧ�|q!��"r�MQѡ��$(���!�-5s!��H	������?A�b<����/P!�D�;eBJ�aa��%n���D)i�!�D.�����E�cY���bHT�?!��<����e�s����F,g�!�$C2QR�Ab��X�6mXRDɰf�!�DP�H�@�!R�X�^�	%Q�!�DPPr��7F	�U2�!`�Z�n�!�$_�	�b���8BD��9W�!�L�G6q�BM�;LT<�p +t!���F�hI���̷0C�%hŎ�#2L!���;?�b�⚻AzR�BӀ7.!���Tش��b�9V@Pp�c!���!�h󎖺'�
� ��P!��)D��-�&
�敹�nV�M5!�D�s?2P�s�D2�TX���ʉ~)!��ǜ�4g�I�z�J��50!�dܙa�b�qw�
�Һ=۲$ˠ@!�$\�tT�p:�� 1�z����ѱO�!��F�dH��U��$��Q	�!�$�RD�]�F-:Lm�i��Ӝm�!�� �DС$R�8mz���F�t�L
�"O&I��b�* ��@
DV<�8�r�"O �y��Jd��MϹ���f"O���%^���c�Gh�����"O�P��d���+&��~�\�"O��CN�	��܃Ѥ�
w�����2\O����A+M�:!÷�(^� ]�p"O�A�D:Vq��hC#/3Ԍ\{R"O^�h$��X>��' ��J�uc�"O|�IiЀb%^�g�C`�� � "On��$�,M�bc��H�*W"O|�	E Y,(�pi�o��%��"O�T����Iv���$YS����"O���H�|��q)֮��NG@8�"O� �Jk4�x`Ѵ34\y�"O����.`���$
�E�$��"O�	HD��)P�<�	P�V!s��ON���؀2;�tƟ�Ct\�8`��d�!������0۠��o�%� g+u�!��L�T>����P;Zh���&��m�Q���ݴ�Q?�pA&;k��p��t���*.D��#"�J�P��a��(�' dt��a>D��ee';X�L�#�4�XQ$�'D����&S2~��@���ɱLє�AѤ�>ߴ��>!T+J�0+���ݏw�fAce��QX�l�O��HתF�D�7��/S�	[�"Oڕ�d�I,@�D�H�A_�i���+�"O>�]�*�nm aY�
���0�"O���O�,E���Pܸ@i�"O�B�D_"v��QI��L_�V�j"O&����[jܢ����\�R���(��IQX�T"���0؂�Aҧs܁3�;D���q�_�?�~�rg��R���AC�:D�T��[�RB�#��2����#ғ�p<SA�uN���(�:j̭�A�D�<�M��^�T�����7N��X�N�z�<q%�ERЃḟ���#l�LX�@GyB�B�a�5��B�)]Q�A!�>�ē�hO��Ƽ�7���j_�8b4 ޗ`#e�D+�S�Ӥ=���e��?�ԽXՍۓ0pC�ɼ���Uj���� ��M�e�ʢ<���'v��! $O��<����P��S�"OL��K�6t(���ߟ}G��rW�+4�H ōD�ָ��.�.���	�	7D�H�Wk�`��\h��+��QYӨ2D��c��	�x�&eG%����!�2,O��<I�Ҳ~��ѐ-��I������H̓��=�6-�>e�=r�i��j�����l�B�<��S5)��x���n��E��Qd�<��;Z�}`���#۬@ҕ�L^�<�T�O�`����-ʔ��c�<Qq&G)E���:V(N��a5 u�<��&J�e<�irQ��YA�aiҬ]G�<A�):7��Q!H+kt�LA�H�<AV�3h̰(�vNViT��A��A�<��iQ!���p&����z�"NI�<���YG���mR�q���ǒHyR�)ʧIeX�Ĭ��_3T�jtZe�q�ȓGH���JP�> D�J��Q�J��<�ȓ8ސ�ȗ*�rar�E�;Z�p!�ȓ5��0�:R-�4\�n��L��'}b��.�Z�R����>\�t )O��=E�t��*:j����VJAHL%���y��ΙO���&+�As(�����0>� �kraȂ`�\��発;5�xsG"O6ɊEb�3;�ě֏0<����*Oꀓr�"0���ptJ�4N��zN�F{��4I�.@=� �9p=!�$���y���3v\d��/�p��Rf���y*�s\��uh��yd�l�F���?��'��)jef��� HNT4]��MC
�'(�ˤG�I�����(B�+��U��'�2�J٫+����t��k.*���'�h�`XX1��
�uI^y�'Ƒ:wʱ1�<C���m��!�']r=GǕ?R���.sXv\����!�S��˛H&�!,X��!!���yrg¦iI
4B�"9z#an�3�~��>����~b�K n]�'@I.D�d��ӆKW�<�fD�|��@�"/��C�`�l��hO?�I�6d�C�
67FI0B�T�"O�1#Í�*:&\+%l��g���z�"O:(��̊�u��8�j��d@n8,Oj9�'��Ɋ?�H��� B挩�Hr�C�	W:j�@��P6��!�D�әaB�I��HQ���l��@��V2F�C�	�K� �Å�	XD��h�T,�|!DzR��{g	�4)u�:���Jms��'D��@%�ۃ	%̐ТbI,6z~��/�Xh<ieO�X7t�X����.���roH����<1Ĥ�r!|�Z@*  ��D{#�y�<qĦ�<��mH�G��?d6d�V
�����)������A ���Pa�!�� *����?t�p�A	�1jv1��|10��BۊY�.�kW�ĢQ|����;"@$�D��d�U9�oڒ�����=N@Is �M��1��G�%��}��iھ=h ��ts@ܸ��!N>�ȓ�� �u�
Rڈ����ܚ��Q���?�3
�(�����_:$�q���k��hO�O���*P�P{�X��-^�5k�'�p��k�h
�'�*��l9�'�ў"~:�A����Z��o1�a(�Ch�<vƐ�UP"�A� �_�$�dF�z?1	���}�g*� n���	>*���(
�R��*`s�e��
�Ș�ȓ��p �g��&�P�b[!j~���S�Իe
�6���T�Ms<���?Yד.9b����/��\ª΅u�C䉊2���rN�c� i�(��C�  ���)R�݂Q�`�ׅ�dp�C�IL :��`�V���അڟzC�I-)����`��Э�@
cC@C䉥K��	1�cSʭ����C�I�t\ɲ��$��y�E�^#3�B�I:�n��+��>��1��^38B�D̈c���T,�����NjTB�� g�H,JaB��8�Ұ�D��^C䉴{�jAy��U�J�n�r6D@�RV~C�	Cz8JA��"?*��(�h߻|̡�$�5Oܬ	t@�=5^hźTL�&�!�d#3��u��A�Rf8i!�KȄN6!��W*�kE�u�ɋ�U�!!�D_	`��s�Q[>\b��J	$&!�D��G�`��˞Y�1���!��;B`�`��?%�j3喏,�!��Z�9�=/HF<R�bJ�g�!���+~B��`,Y�%or�Za�Y�!�� �j�#�7��,��E�2,g�@�S"Or�J���3(�����fG��ѳ"O��H���c�����MI����"Oz�i�0	�)A�ۗX�"O$(���
5�P��q�M�j!�,[�"O*!����yv���,���R�"O|!S@�/2I����dK�{QB�[�"OH
�oֶ;G�ٕlƗCD��e"O>�t�"V�$Aa��Cv�10"O�E�G�[Z�	�۫"-B�"O�0��l�
=٘4�F�pz�(J&"O��0D�if�0��Đ
���D"O�D2��5 ��Ec`�2[Wꙣ4"O�d�U.�8�	�K�dV��"O���͗ O\�9;v�7�H�-�y⮌�S��Yc�IP�@-6A����yM�}���O:��=#��ȸ�y�&l�ܼ��+��3�a6A
�yRX�H��m �;-֞�:��>�y� �;�F$�&I''��36%�yN�"���!%#�fԛ%�N��yB	�=n,��m
��9��[��y���26[̨��a ���dy4Ə��y¯��U�@+� A� +���l��y��!3]��Z�o��dy��Ή�y2Đ5]� 	���F#z�T���@*�y��](@[�Q��&W�EJ ���y�!.4�X�����(�z��r��y�ׯ_̢����xz�Ɋc B��yr�,up؊��׊mJ`�Gl�yB$ÖE}|}�a��r��]'���y2 �=�AR�+@� dƀP��y�FVF����\�6D+E��y"�/�RI� �Q^6D�P�NH��y�(�| 0�b�~]��+�)��yReݧ`
X𧆈�K�� 끋��y��L�@�T�x@��d���Ɔ�yr-N�� ���5Y��r����yb�2X?$��uL�#= �m���y�������97V$��'�	6�y��QP��E�`�F�&�,5�S��5�y��(N�@{rGǼ%x4���e��y�Ɖ��^����"׆ݘ�߸�y2��#p򰸪�����0[ď���y�7z�Xx�BB$�Lc CK4�y�NK�̈́z7jN f��*w@X#�y"n�p��V��mx��Ӷ���yR퉫|�ֹ��Ąl�j�Q�
�y�.��A@�b�gs>̳!�O��y"��(,Ő90�)��vk^͈"�� �yB�0)�TI�pD��g*q�oI(�y��У_�L��Hg���"o��yB*�9
̊d���m�o�2�yb�J RR|��&'�	�����/�y�D��Ko��RR�;2�ej �R�y���[i��q5fJLr`9�	 �y�B̖*V� �/_��R�鄦���yR�/-��J�D1R^� ÔH۪�yrg	0U�<HCh�HSb��#&���y��ѿk9ty��]�C}&�P� >�y򏂈ld�����-�Q#�y҇�<�H$񧉎�!���z��yr"/4hx�toY0P������>�y�)Y2R��-U;E�� ږF&�y
� �)P�.T�\����?�4ٚB"O^P���X�Z�$(*3K��(�Y�"O9R!�M�i�5�-�@ʼ܀t"O8�*Ո(�Jt���t�80�"O���Q�6"|�b��<]j(�"O�]��]���a�/��*Z��W"O�A�a�ϲ6��)B��)b\�"O02W�)?>�f�U&�Zd�!�dŸ`����
R.^uʼb�鞙j�!�d�D��6���H�p�6L &N!���F`�a'eϋJ��e@faɎZ!���%LA��F�Et����� �!�E�:1���>v��:"�@�xw!��n�#S,�5:�MiR!�č�(?}�'�#D��UmS>}K!�$?�	@ńX��`z�l�&C!�Ď�V�\͓�lE��z���TA!��V;�������|�qI�(�7k9!�
[:*e�UΈ,S�&�
���5>&!�$փH:F�h
��]�
p�3��%!�D=h�@a`��r��M�7k!��W� �Ѱgm6�1�ƍ�!�W�2jHcU�4(�zq�PkQ�(�!�䘭9S���&�K��uajղ6!򄌽��	�S�=#��0�Ǒca!�$D:e��`g$E�X5�p���ךR!�dZ.��ABL�4���b#d�!�ك[��i
5掛�RA��"��T�!��1�������9M�X� Q�b�!򄛗pI�� ���)˦$��!D�]l!�DՖv�e1`���=�� �0�#P!�E]zH #�NI�ҵr�/��C!�d�;�0Y�eՓn�P�!�	�{�!�$�64� �*s�H�5)�EpVJ�k"!��ףM�Й��#ҳ	�"��u!��4d��%Rt�\���mk!�$M�\Dl����Jw��a�a#��6�!�$0aO$��IX�L�	5AZ+�!�>VI>qa'NR!g��2NH�!�$*B�h$��ȴ�:��F��^�ȓ *� ��N2�H��ɯ_]V}��
bB�bA�|UD��c�X*0����v����̏a�����MTpɆȓ����ǯvtqa��V�X�ȓ"c@��.E��b��� �=��?��u��K )b�ɒW�}��1H�(Ke�IA�v�1�� t��ȓO� �φ�V:̹7Ȗ�Kպ���#+����EX`9%G:���ȓ d�,� NӾzH����x�h�ȓvv�+p�� &���ǩ��^c�9��e�d��T�[�䒐�M�K��I��$��z�N�?KC��j4�YE�J���@Ѻ��?��m��ނJe�d�ȓaq�볯�!��� ϳPUX)�� U��x��"/���� �3A�B1�ȓ7B����B�97�p4SeŲ6����4�"��b���ؼ*C)Ϭ���ȓQ�n�5�Xwטe���2/gLu�ȓ2�C�-T�%c��X��w*͆�t�֌1ŧD~�!�W
Y�&��ȓWB��vJT$Q��$ٗ��	f^�t��s�:��S@_�x
��p .e�ȓ �����\�Q6��'��rY��S�? �ЋPNZ�.:�g&�(Lb�-x�"O�*�E:I�����P���0Q"OE�G�գ���O��}j�"O�ɓf��}G�Y꧊�Lƈ���"Oz98s��9�B!��(W�J�x��"O|b�lF�nҩz��q�P���"O�`�p��]R����%�*�"O����ԙ.T��kA��;�����"O*Y���C	Y� $���a�zLj"O�y�"m��n��p�=U��0�"O��B�1~xaF�]*���pp"O(��ql��~$���l ,`�Es4"O��� �}���a��_�Yr�4zc"O��s&Y�]H���ݎ>b�$ �"O���D�ɣ8
�3�T�MBZ��"O$��T.J6v�t�j�聀B��ۣ"O�%��eI$���v]�a�"ON�R��Z���/D1wA�i�"Oh�P&ܽ'����̒�0>�!"O6��w+Q/p,*�0�_�*����"O����"�\�0�L��{,�`"O�X�v
�%=8x��*�n^<���"O�%��!� QfL���T4-H�5�"O>`:�ܚ���W�ڡ:�r0Zq"O>,�m�
D�(�vFC���*s"O.L��D�<MURCE�C>��s"O��G
�u>��[eN	�2)Fb�"O:�v*F�mE�b�764m"O�]��"��P���L0w��D"O�`�#S5_u�xc
��J�pC"O�eHS���/���Y���` 0�rw"O�����0��� �ǟ+�z�Kf"OBPr��Rt��׫Τ+�p�( "Oฺ ��"kF���R�6WPEc"O<,���X)8)c�
ڳa��"O܌0tj¥} �0�
�5zm�"G"O�����C��l9�(�	%|dT@�"Ob�/��(-L�T	��lD"O��W?fyH�[���__"�+�"O�"t���w��K5CZ�[��B"O򝘠�J ��:��H$I��"OP5��E��o~�M��!Z�`=��"O� �0*β,XּT��-��4
F"O�jQ蟚~�bIh�ώ
Y�n��"O����)17�����Ǯ$���3"O4l�0�4N�$�dW;rϬ �'"O����~���oa�gy�B�I�Fc`uh�?9(���qD�"EdB�ITZ�u� �H�r��E8��B#?j(B�Iq��@YPi)i���r �G� B�I�/�����X%����# ��3�(C䉗=�>`&HZ�T�)�����+w�B�I'i��,y�_yQ�Ybv�_S?B䉎<��s���2jhŋ3�ޒh��C�I).j���oȕ9	 њ�I�$KR�C�I�f�	���A=^ʄ@lV?z�B�30{�U�6l]����Y �B�	�a�$!���]��	 �ۦ�0C�	5?D�[��aV�u���D�c��B䉒>A���Wq�y*f���uX�B�	-T�6��K�<���ĺO��C��%� ��MU5��qA5�N�ǼC�	="��G�U�@Ƣ]:��ϼ��C�I�� �C�?���1�Ҳ'�tC�)� �Ds�.N�~��Tӡ#x�}h�"O��ZdF��t�)�B�1�"�"O�y8t�N�Nn�	�*̣=�`�b"O�ɳ�K��4 @iT��j��"O��ɖ
���b�ۦ�O9Du�ea�"O^���s$�BaQ�]j|9A"O`��b_^�ݪWϟ�vX���Q"O����IO�b^T0L�I���u"O�m��D���9�F�3�Ĺ�4"O�l���ɓA���ВO�3W4�"O���U�U0Iʼ��D�L�G`� #"Oʁ��.����@E+����"O�ш'Ck�ꭘŁ�`&����"O����+��\��ڡ#Yj4~PɆ"O>P%חK�Ĳ��A�0$.�H3"ON��Ui���+V��'����"O$�I���D`�����Ō.J��22"O��W�^��<@M�{;����"O< ���.&
J9��E�O7T� �"O��e��0�D+&N J!�"O�1�3�]�I�k�m|��e"O��i IHf��*h�X�y�r"O��P��'��=i  �4.�D�{�"OD�Q�Ɗ'.l�	�h��/�J9C�"OP���F n�ՑP�G7u�6=�v"O�pS�3yq����?��@#"O چ���<A��{�È	�N��"O&h���cs*Dhڗd��"Ov�p�/C�d����aGs�(��I@�<�b�Z��rg�Z�/ɰR�#D�@Y�:M�t�@C֊-���D%,D�ؓa�X��L��L5jZ�z�-*D�,� .�:<"*8�+͚B��@��=D���U��hB$�Hע^�df���g7D���SoZ-Mj�b�`^�B��|���3D��1���dj\�A�@)`�TC3D�T�ㅗ�E�r��P���P�e/D�`s�iR�$��]!C%<4F�$*1$"D�����;4�h���%?u�ҭ D���/�{غ�PAa[�As֨�ï=D�����L�;�N7xC䬳T�'D�P�ҩ��:�|��UH�&(Y��$D�l���H��`FIK�&�}�sf�O|�=E�t�U�w!&�{��+IG" ��'��2!�DZ#l��ys��.o8�$�q&�1�!�ձXS�� G�,W"��#�Zk�!��u��ǅ18�-8��4t�!��V�������h'V�&�A��!���� 	�Ԯ:=r9��)�	�!�N�0�HH�T��!&IR��	��Y[�'3a|ro�F_��Q��A�L�و��3�yA��9>	���b�~HPԡĳ�yR�
*J�ʥo��iީ������y�(Z,�Fc��ۏ\N^|�ө��y��\$�5HV�Y�!�.H�r�N��y�F�BF�ط�ϿK0x�#䁛�y��A�1,佣7i�	6թ�R��y�O,8�� �&k�p��/�/�y�f<��(�r�Of�y2m�9�yr��˔#���\�Z�sb���y2&�j�
hH�΃Z�����֗�y�O�,߼��tn�O��i�GD�9�y�cPc���i#dB0 ��9��Z��yr��9w�#�㛅%P 1�0�y
� ��`J�H�:�2 E�g�c�"O*�:ש@��,�cv
��q���`�"OB��c�C}�Ԁ�Y�s``yT"O(���)[�w�а+���\���"O�9Ra�ϓx�(!�r�	n>�q"OJ
���yA@T���/&N���"O�T{��\�Y���K��C�>i`2"O\$;��/>}h �0�ң]��Ց�"O:������(8��̗V� �QW"O�Dq�.Y� R�W�L�D��0�y"�S���Ĥ��:c@\�y"'I{�����!3���в��<�yb�����z���7�8Q�
4�yb�؂rK��k�NZ*��4�5n2�y"�\< ��E����q�i��ȼ�y�'I]@�h�T�αu1Tx �#Z��y��j�0%��Ts��)��dӳ�y�$�Q�FJ!Ɠf?�` �EP��y�f*A^���*БXGb�y@CI/�y�KT�~��A���ѡ�۔�y£׹0O^�;d� Ԅ�C�ꆓ�yr*X65� R*X�[���I�N2�y���~88ᣢ���iBH��y�a)�ִ�l��c��l��$���y2cS�RH�e���]|b`����y��߾8�
h���Z�Y��Lj����ykaX�ڔj̹S�����	C�y2�;',�pY��͘�8��#���y2(�g��X�8di��	�y"���P2�t���Ϲ��L�a��y�l�7��ڱ�]�o��8�.R��y"��C�
t��e/,��XJ$��y2D�3ؤ!��M�l��A4�F��yr"Ɨx��I3�E.4@� 4�<�yreK�i%�A�"e/A�0�"+�y�	��f����+B)4��D1��Ɓ�y���<�t��B^��
Y<�yr��0h����A[���2*ǂ�y�N�@]�9s��S�8ubU�EU7�yR�ԖG�\y��!�"� U�Fƞ��y"mѦu` \xW�X�2����yBX}dt=�ֈ�O����C5�y��ۄ`c��[(qX �àǾ�y����*��q�D�j��{�ᄏ�yҋ�%��|�a��!eЂ�B�C�y�	��3QTM#��i���0�G[��y�〖!�D0��
et�z��yd�$F\	cf& :d-��:ՊZ��y��Q�̵j��9*�ʕI$#���y�*D%x���9�@�2�JE�� ��y�I#�Y��1B�5���X+�y�ء>�
�&��3f�@u�֭K�y��O�_s@��DΘ�Fm��P��yRM�6)�8���gǉF��H	���y���(�����_�B
P=C���y����i�6dyDBף5	��₩�'�ye�>�Hrf��!:�Z����y(\  �L�L�35V�!�V�ϱ�yb��3]��e��, ��Z��ƙ�yB@ Լ���`d�S��&�y,���t*&䕋�X��TǛ��y�����0�)Ќ"D��Tc�#D��y�' �6@ Yp�S%?�H�R���y�H
qD.�����
J�u���4�y
� �$�JI�n�@��玁,ce�pq�"OBY�j�0���6n�'C��� @"O>���Q?3�<1a/[�,�|���"O�E�4M� r��b�OX>��-��"O6Y�d��Z��S��^�c����"O�4YqG�|8�!'�1s؅��"O$#�E)l�-@a�բ���a"O(\��$R�d��N(Y��$��"O�@�a#�?��p�I's2 j"O���_8&M�*�M��w���X�"O<���Y�N}��6*�t����"OF��D�I~V!��d�]��"Op�����P��B��<9PF�c�"O�Xa`%H� ��� (|���R"O��4�ǮBA�Q�
$R�"O��'C-�8���	�_rZ=#�"OHȪ�ߟ��(Gi��L�~�b�"OZ�y$ְu���D��b�Vm�#"O�=���0_���F�
&}�^��Q"Or`�婂&ʹ{� �'2LP��"O���!�ǃiҨ%h���w���"Oy��=Ne2"֫]�h�Ț�"O�ٓ	�	h��#�
A)}�<��'"OHiR��QR�pCd��H�t��B"O)�vc
�KyHHa�,�΁�"O�PAUe�,Z���B�O��a@"Of�!m�M����֘$"M#�"O�,ز�T8t��Ui��:S���#"Od]�V� -���3C��l��"O\�)��1�(�����[m�e:�"OPt;�j	(/������([&�8�"O��	G�	=D �+�GML��"OfI��#dx��*Y7>�B�X�"O���02��A�B�8��yٓ"O��YW�PQ���')��:��$QV"O�y�/�]���'Ǻdm2�;"O��{dU��j��c�VZS$}��"O�1�l�[��$F�[K���u"O���U�TY� ��eH��b�"O����
�{�ۡl�5A,MK�"O���)�$C����̽=+B�P�"O�x1�#�)6��!�0 � ��"OrT���h�t��@_k�~U�"Oh�[$�
6N����pA]�^�
�4"O���v�N?��(���;°�K�"O��S�LJ%v�L��{B�c "O�L 7�3�� [�ϊX'��(4"O ѓ�F)s*X�֯��'�bts�"On���T`��)��kF����"O���e݂,��"& �XH�"O8�+'�Ɯj�B	�,�sjA�G"OJ�C�ͮ^�z�"��U���W"OD`If��n�b:T��+Ӕ�JD"O]�@�L)Y�Q�D��0�Z�"O��CA���\uT)So���J�X�"OT��Z�2/M� oö7��Y7"O`���]�uP Tʆ�P�!�:��3"O�����c��d�s͋7$���"O��9`KMV6JX��	�AA 5�"O�aKѣ�#�X<jw�ʌA�l���"O*`�Ä��e��o�s� �@'"O���bS-1�����HD�rU !"O4����%as�9z%�_�)��"O� 1��4U�^4����z�"�q'"O� �1�Cѻ�R��%�C��:�Q"O��
��G�+� �cǧ҉8E��+�"OƱ F�ڡ3�Rp��A#/��Iya"O��hC��.�R�2�%)�ҥA�"O��S�[$-{�m���j�&���"O�D�7�N�K;juVĐ���"Op1�D؅��M�H�8��"O�@�u%N��G�:oCֱB�"O^ii�EH�-�AP0GC4 cN�BU"O�5�"K�9"���Cݛ4S\�$"O���҆3���j1�C�#Y�R"O���� I�Q8��@Q���j"�6"OJ�['�E�P�6dHf��K�.{�"Or��;>:Q�c��k���Z6"O�R+N�W������˗:�>��p"O<1��j��Fhx'I��ܙ��"O����Φq~�Z����a�"O^��ŧ� z�腩Po�*xrrT��"O@$�+�T��$<:�У�"O�B�dS�~��d�#�*)�Q Q"Ox��*^�:ǎ�_<(2�x�v"O쬻e �)y3HQ�Q �4`(�3�"O��XC���_�x���ȗ��}�"O,]	�����}�R��7�*�"O�T���Гq�(嬎
069��"O�� ��C!N���Åلx@��C"Op�#Q���ft�!�18'�x��"OX�el��G����ˌ	�> J�"Orњ1�E�YZ$ոg����<x"OT�ьۛl�,��"Y�N��4Z2"O�ݫ3��}����[`ިa"O�l0�jV�L��02���!ZX8@"O�}@L.F��D�N0h���"OjT[sIP
lL��a*V.O���J�"O�А�0cD�]p�J�4p���"O0I@�\�8���:̡H�tUh�"O:�L��(uc5Q��R�"Op҇�B� Hx�B�C�F�V-�"O0���Z�$��`�>��4�q"O�%�#� $qk𯎽|��:b"O<�U��3 DU.�Ԁ%�"O����4v��GQ�g��(�"O�Ģ�j=8�D��"$�@"O��h�-ՏZ��Ik��K�B�sr"O�``Cե+�lP{4BQ' �B(��"O*=yV������P�J�R�dQ:�"OR��# Ĉ2�V��䖐K�vpRr"O|i�-^c��t�PD�o����"O.T�Tg���%�ӃW#�N�#0"O����Lx�Xb�#��h�"O����E�a�D�'�jԾ԰"O�i�װ9���hb��W"O�0G��`�2@�2f`�<s%"O$̛��ϱg�,Pp��.JQ����"O>��$�H
b	H$�fIT�pBU��"O��'�%g7��7H�P����"O��j�l����M�	���f"Or�������'a����`�"O�M��V�Lx(p��F5�6Ai�"O��qbf��gYT���S�^'"OZ�E��H� �͍��NM�p"O��+�N� ��]r�V�9R"O��:r�89�ź�kܑ�p<�e"O�!�Q*�������O �1ϸ5��"O� ���`F�z�^4�u��ּ`!"Ob��5�hդ�Ȥ+	�B!tY
 "O^U*#��9D:M�mY-�u��"O�!P��XBZ���ҫ��C_�� &"O������j�H]�&�J4A�,1�Q"O�����x���A�?<U}�E"OF\#�&D�dy��n0I���S"ODu��ŕ�9�r$0(1���b"O����a� T�Xu ��M�4	�r"Of�wj��V x��d,C`�|eX�"O\@���˲uc�B��F
>��}�f"O��:2�ز:��&��/\} ��"O\D�IS�~�n�Kb u=���"O�����' -~�Z�C�g &��"O�=˂���n����тJ��!�"O0���̀�����p�3F�>��"OB@83���eM��:���,j����"O���7E%,�Ƥ���U�z��h҂"O>��v�֌�RP"թ�.� ��"O&E��DW�GO�xG(
�v�"O&9;T��<7�p����.4�re�"OVɢAȅ�2J���%?�qg"Ot���-G�#A4��F�I�\p���"Ol)����Aօ���ʓ_B|�1"O4�R�j¶4"�@�UHڵN�4��"Or����H#V*�q&'Q�)�0�"O��H�␽4� fE� -��Ty"Or0ۆ	�t�)���.��p3 "Od-��*b6�$�B%�u��<9f"O�][s �?M]���YO�-Rv"O�)�����L�� 0�$ưJ��$�r"O�M�#c�TEJ�#���L*�"O�	q��~ ^ �3cP0N�RTb"O8� �g�`��x �g�mx��6"O81���Q�_�<�kfݮour"O������Nޔ��H�5l�xB�"O�% "�Vd�~e��č�\A��y"O����O�c����7��Y"Oܝ�M]�ozb,#7)3B�V���"O`�X�,37����M(bk��I`"OL� �ŬՄ {2��T���V"OƝ9c�E"��E�E�o>dM�"O��S	�4�`���:2-���"OH!Z�X�j�R��"���1��p�"O��Zc`L�AH�-�Q�א�!G"O �h�N
L��D�r����(;"OD��Q`����"��/\��,�"O�\;em��KX�ASa�
5U��""O|���f�F6�X�D��1%�"L1�"O@��en�[ӖL� /ʔx
H�Cv"O��"�aU��ESd�Z�O��iV"Oh��?W�d��j��C۞-oB�	�{J�m`���%%�t��'[�W�,B�	�t
(�`Pe�G�jPrq�5:�B�	81�����h?����׼b)�C�ɢ6�5� mA�EEԅ�դU3��C�ɼg��i��Z���u ҋpJ�C�I+�~蓣˜�`�Hط���P�C��2.����b��u>�p�5M��jeBC�I8t�M���-t!d��b�+�~B�ɘH��Ud�W�6T
6-N�*d�B�� �x���Q�StpM)tE;�B�	L��qf�F�l�PI��'V�$��B�<�[6Na/��A��#/��B�)� ̀S�e�^�\$ �33V���"Oz=�Rm�}��$�2BZx�I!"O.T�W�0�ӵJ�%Q�v)�b"O� ���Qd�ƅ��.Ӕ|�̹�U"O*�P ���Yc ��"
�AQU"O0X`��D�<�Pi�͘�<[zu�g"O���OH)D��-�1��)9=���"O����o��@�t��~(��w"O,�`dM�)�n�ic��~���B"OH�뇛Z�d`�1�̶����"Oԕ񨜧O߆���!
{}PTcW"O�9��S�k��c$c�=|�y�"O�ek�GE/`4�M�焄 ����Z�<	�_>va�	 ��k�>0ٓ��M�<I�eG�<Aio���FmL�<�C-�"Z�Lr�!�;J�<�Afj�F�<�c��
�tI�W�	���0mRK�<Y�Tl�ph]�r�$�҉O|�<�f+o�hK��	2��4��F�y�<I�
�k#��;�c�E����*u�<1V�9J5�F6k�]��J�s�<aE��u�V��V�2[e�E�M�l�<���:\�؃���0��*�i�h�<9�sL�("5n��B\H��Ka�<1`�m��l��+kF� ��ZZ�<���^�J��e4=o�a�VO�<�c��>4�I��^7\� q�Ï�M�<1q Ћ\좸�a,ƶ?��Yzc�u�<��%�9̌� ����yД��h�n�<1���g9��,���G��^tLC��$p4��a�#��PO�i����"Oh��e�	q�� L0V?¹��"Oz����D�{J�-{�&ڤc��y�"O���L6�0����8,����"O�iJ���`��dY𤀄��:c"O�\���Ii,���D�;3x<��"O��`��K"ɔdX�S�W_��ɓ"O�D���@�����g0~��"O2�K��4r�0���5~	��X�"OH��#k��H��ߺ�.���"O����E�T��M�)�����"O|���'�KRJTI���)��E
f"ObP���X'D��D"�z-	�"O�9��Dxh8��	�5
S"Oz��K�asfә6n��@�D�z�<a7�Z-w���K�B�w�����k�<��&EArތx3�H��%��@k�<���3F�5���<ZaKA"�a�<)TL��_��Bq��/#�@��dv�<�����F1�oԠ\���D(�W�<9d,�X� '���@���	Y�<9�D҅"�P=Ic�!W����`�<ɲȃ�i-���F��]r�ƚP�<A �Տd�����b	��
���I�<� �14����B�	N��=��i�_�<'g�87ct	��O��`|Pიp�<��.D)7��)W�5Ж�Ym�<�e �=���G�?��;���a�<�@�S�ح��٤<n���Yw�<�3iU�6LX 8U$�!Ԋ,9���r�<ac��E�����L
�OU�Ő'��p�<�smǖ)�j��RCY�}i A���_s�<Y�Cn�$ݠ���9v�bJK�<)D��>ۤdZ���#�HD����Q�<� ���%������'��Kh�Q�1"O^x�B��9
�&!B'�XI Ȅy�"O�4A���&?.X�����Ni�"O�P���D(n��T��e��Y�J|��"O�,��,Hr�2]�C$ ih��d"O8C�O�w��`�P g4V�3p"O�b��'ex8co�X���"O��$,�7o�Ic��1V�$)�U"Oʼ��l��e�(�,��*��"O��)8ph"^�A�f��"O��3/�p��$5�@Qɶ"O %�r��*)p<#5����A"O�y񉇂.�� q�X�7"Od0�P��:Lmey0/�-�r��"O�x '��)�4��ټp�0�0A"O�Т"��)bQR��# "w̚�a"O�i�t�Id9���</��ِ�"O҄yB��_R��̝v3�ݓp"O�T�;�U �2 ���w"O���P�^tf�i�q���K,R0Z3"O�Q�G�jɂ�z�g�	��T�"OP�QaO@ð���G�#{�1�%"O�F��c���c%�Ec~T|0a"O�-�PФWlf�2��ο8�Jp�q"Ot����[���_�4�<�C*O8�ccF�f�b4�T�ݙ?�� X�'TX���m��h�n}rds
�͇ȓo��A�A �L2U9CBڒT����);�Pb��/���s�n4��!����Ps6H��4�����.�%Eˈ̄ȓ;��ꂏ��*Xts*�"p���ȓbQĔB�h�?_��� �N!}ؖa�ȓL8��c�E[-P��{�Ȇ$��ͅ�h��	E��_RԫæR�v�(���]�j��t#�"%\t��uNB�� ��w܀(SI��Pr�s���>8��h�ڭ���59ܕۀJ�`Ɛ��ȓb�.hᔍ�3 �D%+3n�,l����ȓf��H��$ؓX�F��D�'QX����
��-�e�R,EP��S�6���Ep�S���� h����C�L�ȓRq�q���J�d�{�F��\|�Y��$��\!dL�}�ȑc��#Xq}�ȓy2��˕I]�jגe�� @+��ȓV~��k��$J}`A�Ĩz�t�ȓh��5`�⒋dd�;7��'E�m��d��5˰�'����,� +,��Y��� "�Ȫvn�}�4b�'�^T��=ۢ-�F�� Tƌy�'�|①Z<Wm4 ��3e�P9�'h@�P�`ώ��D!��V�b�'���3���1?O3�
�2 �H8[�'&h5�v�J�jX}������
�'�Ȑb��4�d@�W
�����'����'�J?�)�l�9|����'��L+���Z�z�ȵ�:?1��;�'�2]8�lت:�-�1��K�f�R�'�쉂A���L�r�E�-& �	�'�X��P��o��(1B�X�`�{	�'mRQf��z�+Ј��F�n���'��#%!Oe������T+��)+�'�).�<�H9�6��:Z��R�'la
fNL3c`�4�v �?}�%J�'>�Y�Q�]�2��M��m�/�9�
��� �R�Y�;� !�1�FPhZ��"O��b��6@�8�Qgw$�[�"O"�C�R%w��гB#8p����"O�XY�ΐ0��i�GI+`�e�"O4���
�Rb��:�A�&�$�� "O�達CBe�,A�K���T��7"OD�q�
@%7T���4�F0cY�` d"OZ�._~P��t�Υ)L.�`r"O.=������X�@.%Cġ f"O|%��&����)����
�R\0"O0�0�J� qp�̟]ĤJ�"O�b�]�6��E5XDJc7"On=�EY�[(U{�M$�n���"O,��C �a�Dq�C/r=��"OHm���ߌI��TáO[�t2p"O�Y��k�jž���M�yM��h0"O�õ�-j՚a�N��&�"O֌2'�ӖU�ܛ���<`6��G"Oh6KC{��Zp'�a��+�"O�"�@�;	�8���D���:�"O.)q�IJ���#��&Q*Д��"Oܵ���BzY�'�R�5��pч"O�-�!Z0-8���G�Hl��"O���׏X�A��ղ�Û:&�E��"O�p�Zn��m!���AĢ�pa"Op�{S$��XH۶�=�@ܙ7"O��C1�ɓ"�eb D%"}�1��"Ox	�&�}ň1B��yd��iG"O�)�׼tt�2F�1lFn`s�"O�i����J�l�)S�@�^f)b�"O�0+ $ET M(g�O���"O0����Q���wˇ�$�t!��"OR�hf� y��ܨ�ʎ�9)�1�"O�! �Я+��b�zy�"O� ����r���0@��x��%"OT�z��Q�Ӟ�jaܮ0N����"O��`���=8Q����`F7 ��R"O��hc��U��-ذ���Z�R��"O�qр�|.����"��i�X��"O*�2�H�5�Ҝ�!�.�|�4"OD�2�c*���3�A8��ڧ"O�}�rg�9q���U��2�V堧"Od��Q�4��m�O�P�fJQ"ON�x��$=��ѩƤ`�\R�"OZa�F��3��53@N�0Y<�Գ�"Of���`�f@�Xn7Qj�P"O�� ����CM�h�G��ULx�10"OF9ãV�H����D�L%:d�#�"O]�F����hr2�X�Jφ��"O�UkF$D"
���&ˬ9���a�"O�����A�l`򢃱^����a"O�8�T��f��5;�BH-!�����"O�-3qa��6����ug� 9���3V"O���$�D�;w�+��$"O�MZ��ǻ���eR�㖅E��y�O��`� ���4dՐ�d���y�k�*�b}��l�����$�ߗ�y@^�8��%��!��]/ M�C���y""�YUv�ISEVMR�q	�G��yΝ����5L��7i>�*�/��y`�����JI)b6M��FG��y��ӋC�Щ�b�9TfL���7�yB�~�� `�T��8�� �y"�6\��8����]��Ӣ"��y
� ��
tH�~ND͐"
�K<�t�"O�q�o�0L��F��/4�b�"O�k��GogfزP�^=�,i "O�M@a��!�����?e���"O�}��Ϧ V>��C��*h2ys�"O�X�'cM's��q�G3 隑"O���C]?<�䅓H�$#�"O*4je�;Ev�:gW�g%�D��"O0<�E�E��V ��D��l ~� �"OLͱ�.�H��#�aK09أ"Oju�U�Z�_�
�G� l��IY�"O��KvF�@��� �n���Ӡ"O6d`5��n��j���/%��iW"O��v�.b��[�Z�l܂5�U"O�p�"^�.֨��§�mƂ� �"O�<;�'�C̀M�W�Tj�f�2�"Op�'G2�,�5 ]���)u"O�)1&)ה4aX1�%E?��$�S"O�Y`��4�Șք���T1�"O��0�?]ڲa��-�l5У"O�M�g(�=g�,!���y&h�r"O�8���V���1#�Ǆ0"���D"O��	�NFvt$���W���`"OT��iQ
W �r�� �x�n��"O�\Pco� ,�����"�0��"O���s���DM4H2ǚ~�!s�"O��ڗ���)�f���K�3&�%A0"O>��1-�w�bY
��8��E�"O�d:�� ��ݒ�o�!9�(QK"OZ����85�`��F&_|��	"OJl!f��32lF���Nih�+F"O�� �ǿM��7!f��	#"O0@XV��?LTm{A�W`��@1"O���p�[3(dl�'O�,	U4�D"Or �ğ$#NqW@UC�]��"O����!GH�<��2d'|��"O�1h�-Y-	����>Pp1�"O�PR+^�i$�9�ӭ��DkP"O���Z<��3k�\x��#"OD��Ƈ�T��D𦏋�m�   "Od
ǹK�,��ѬJ��T��"O̠��&ƌ@�8�yq*Á7Ĩ��"O����N�G���sI=yѺ<Z�"OX��î��D����-ݥH[�c�"O Ԓ����{��r��)&Fl��!"O��j�@@k�p�V��X&|	p�"O�!0�+�~��H G�$K^�	�"OJ� �]���d@�@�[���%"O`��&�.xO  ��!I���y�"O��
��T�Բ�n�'� �1"O@��'h��#��a�"팂wS��i�"O8�(��Y9A <:�!��?�(;�"O�5Aga�F�u	r �3n��Dk�"O^�dCR*ya�����N����E"O�Vk>e
\����8���H&"O�!���W�n�8 �qPx)��"O����n� ?���`E�m����"O�񡢫R��,P�ȸc�~<I�"O�4���RF� YdOZ�@,V"O�T`0��'��X('-O�J�H�&"O*��ʍ4�~�i�;Tpj���"Ol`A�U$�P��c^}�""O*�r��-��b�		�F�L�"O�0��-у&�P��(�16"O� ���Pgݺ{���#�� X"Of��� L �4�'�=:���T"OLaA��}ȰɩfM�;)jA�"O�)з��5,Hf�" ��3;�=R"O��e�qm��
sE��Y��! '"Op�gmܤm��PP7���r���"O�i���$;���3$<&�D�Y�"O�� �߭4BIcw�ٹ'n�1b "Ov��g��2 P�ԿlY"�(&"O���K�ke<d��7�\"O����˨� E�� \�NJ "O8`2�oĕb�f��d������"O��FOP�%�B=��/�.~��XC�"O6u�	��,��.$#�.�q�"O8��ǝ�	��mb Z�p��ĺw"O$yԃ�<rZ�Ʌ��"��� �"O2��g�޿Sv<� &�ԡV� �V"O*�s���Cyt8w ·��c�"O�A  .�T@�dt"Չ���A"O�xR�nT01��uO[��A��"O����J��WB�����"C�j�[�"O���R�H�r��lIvQ�2�0�X�"O`�آ�
�$-3G�5+�B�"OJ䙷��c������q��\[�"OJ1 �c�PY�%%������"O:�ȗC�Tb�Jgv���"O>��Sm W�8�c�Ӑv��|��"O:)�j؏�t�Y��``t"Or�ꥧW�%��9�ꑪI��8�p"O�E��L@?	U��b�H@�0�\�@0"O�8�O�^�)�SI�q�mW"O����̣G�V���ƅ#vi���"O���z8��;��7@�`5��"OX�KS��9�D(��,���0�d"Otf�,g�, �C5
NbAI"O0\��k�)����E�'>��"O�qR���9���!F�NS�)"O�5)bÊ/�Ԩ��d���T$��"O��q6�Ȉ-t��Pd��3�<-�"O����oU�j7�h�V	E��܀K�"O�9�S
O�kڜ�j
�J�4��"Oʄ��/R�5-Je��ajR�{�"O�9a��Gkb�i0MR6s�z�"O��p���{��Y��% {��D"OZq�AD� `0�j�E�8I����"O�M��aT;�������>}Py�r"Oj�#aJ�!Q���I �~鉓"O�hb�f�D�PEQ�$�z���"O��:S�ޜJ�� ��π4��u@W"OP��g�P!$�@�'F+k0���"Ox���"�h_�{�dOnQ��"O��@��ء$��:�b��2l�U�"OfcV��|��xQ�� �]h��;�"O�IɁAZ�~@\I��@Q� ��`�"Ob���/Yaq��7�:er"Ov�p��"X]� �	 N����"O�����0��@�%eٝ%8��a�"O���Sf�aɾ�����;/!����"O�$pw�t�|	"bcɀ:����"O<�:Gm\4�!xs!PC�M�T"O�8Ӣ�>V�XjqN��k�L�I�"Ox�2W�֜l� �P0� �B��HA"O<�JR����x3��#��`�5"OTH�����*n�-�G��q��X��"O� (HgA�([�X����0����"Oh���"�*Y����P�v"O�㗭bS��9W�ߣ�0���"O�;qkѐ>8� 4-ݳi��C&"O��SC�.!,�!�&.��p	0"O��q��2Q�cCٸR�`�X�"O�D��i½.��=�;|¬���"Ob��@dƎ7g��×���x��"O���W�̮`d`!�1�B$�ƬP�"O�@(��6� =��!��alvi�"Od���M��1�̉����8`��kV"O.Q�i^T��1�L=6�=�t"Op1�t�
)V*�"A��@Y���"O|=�7a���A�&Q�/@t�y�"O�Zqfπ\s�\���#�X�E"O`��w�!�l�!#�"O� Zt���F"R���U�q��"O�j���#0�(y�ԇC�& Daɶ"O �p Y�i1��" �
�>���"O�P����!qT���K�:�MF"O�+���Q�.���M��R��-��"O�x)e���0�x��S��f`+"O8����A3v(�U�� �*�"Ox��ɃD@ ���ƤM	�$
"O�}j��01qH]���R�i��yB�L> P��m]>�s�/
��y����(��T�Q�JE�W��͐x�FF<��y7&�u�x�HY�>O��� �+��V>*��S��'Uz�Yf�:D����`��NH"�Z4e�^�YѬ6D����+\ G����VJE
�+6�O��R�cY8���i�{tK��ڣK*��J�܅�	/TBbn���%�ݒCZp�G"OJR%��(�!�"_8��O�Pl��Tp<���� 	�2��3OH�5�:#<��!�̤�����u;8ѐro��V$���	
�(OΘ�p&��Pu�;�*�gZ:@At�]h<�`�I?P׬�hE��^ fVX̓���M+#�'�'ʭ��g{=~<`��(��
�'b]��X��*d�����{���	�'���H��3��PqM�e�4\@�'��PFČ�IK" sP�V.Y�q�OL">�}�ۙ}���u��6U�.1�uhE�y�S��A��?m�}�$�V0�y�Cɤ92d�L	�m�tF�y�iGg�ĒR�G����N��y�ƐA��(��ƒ����:�(O�U��	+H��K���s2X9���D�<�W��>v��t,�5
�����b��0��?��	E�ɢKɀ�1��?�%�'�4�����@�n�0�a���� ,���
 ��L��LZ5s���>:�mӔo�q������#��e��5i��B`�
����y"k��uNԌ Ɣ�P���ph��yR�-9m�P�2KZ=u"�sJ��yb� -s�XiF��mM���tg�y2�яc�։�HW90�4�0$�
�y�gO1w���t�]�&�p��DL���y2"�KWP���	OҬY���0>�K>9��Sy��	�V��-?R�[�T|�<�ƈ�d�y�&���zZ��u�<��@p�-�ׯ� R�"���D�p�<���� &�}��+��8�P|+��
e��[-ў�i�uO@�iuB�0��F!op��S�? 8�!Å�}��䚕bʕ}p"O
�����_O�YH`���U�� "OHqHB/��|~�A��V�n{�,[4"O©P.��l�����@MZ����"O\Ih �ՙP���Y5/�2�&��@O��&�8,K�j���6	�pSΏצل�{^Q��CY"
�b��5�/�,�ȓD�b�̄irr�Qq�4F@�)��K�,C`�F/.�;�䅘"�ҰG|��)�'=3⬒b�M���T������HH��J����,�lح����Gx��I��i�FM��;~|�q�dœ=�C�ɣX��j#`�|�iXF�U����0?�w�ԦRd����;]���%��w�<ir��@ ܔ���42j���)�q}��)�'�H�a@�;�jL
d�I��F~�>9�4���ŇgWfa��� m�BlKKY��!�D��4O����Ƃ�F�R�aՀ���qO����fS
��ƚ~0(B�e,a~bW�� !A@�RlL!14��^M8炻�\&��E{ʟ.d�$؋}<��$K�@� ���"O\e'� a�,J��ϐ�ɤ"OLI�`$�&���EC0Qi�uI�"O"QjԊ��v=L��iIt�t"On1X��A�yc�(��bU4=��؆����'ay�&^���r@�B�D�Z�8Ћ��yb��.�x��_�8%�0i���yҍ��[�6Ĩ��T !�4�y�	Xi���(TЄs���yB��/���1X� q�����'�ў�ӆ8���?~�(�͍��"�ޚ�yҦ�E���`�A��= �4��dG6�y2�^%�B�`S�	# ��"$["�y�Eۀ;�,Xe��'"TB@j����?y��$,��F�R��\I�`��a��>�<���'"�&!(:��}�RI�>�����'��S��Ɓ���sU��'Jx$���D1�^μ5i!��1.:��������'��~b�ْqmx,Y��g�*Yi�����y�-̘4m�Ժh�)=����JX>�yR��"c�051q
�(S���&���M�N>������c�e�Q����6�z ��y�΋�V���g�[��������'�a{��Y1�$@(1�Z4��C�(Z��y�C�.b�DT�Ɏ����중K�4�Px���'M0�t[�N�Xʚ��#Ɏ�yR�A�en��$a6_�jL�P���p=��}�f&w-����ŕ}�@1D�7������Oj�	ϟ��|��C�vt�����i��OPM�<)&��48I�d8�H�p�΄�C��J�<Y&98� MZ�&���|�b�^E�'z?em��+��*]� p�FgӤH8bB�I�7��<r�!H�I��M ץ���B�9<A�EW�4��}k�D� �B�I�8Ҝ��k�<t
��2��N;a���D!�Ie����B t%�	��o�/`�Th���'�����<������ .L��فE�f'B���E��y2���SSr)˦d>JmV��b�K��'�<�DyJ|��	���o��1[�c�}]�]&�T��Ck>��1�?	^e�����?�X(����O`4H�
$݈	3RH]�)L�Iq"O��H��F9�L�f��Ȳ��O�ꓲ?�wf2�IW��8]�d�qRP�u3��[��4C�	p�҅	��2JS�a���Q�c�P��)� ,�[�K�B>biPe%�8b^�QȄ�x��)�S*���hDh��c^�r���6�TB�ɆP�l�ࠈ��g~�����Dpx��]f����
Y
K �ȓO,4�ۅf��:V�@`aU'p���O`��1e	���p��O�J���"O�u�+�����(��ܷ{���"O9K`�_��PQ�_pu�'0O��P���SĘa�3�D��8�կ�(&�C�	5R�a�oр?�z���,@�C�I.0��@Я,'�p�ю1aC���+ʓ`����F]�		��أ $����^�Lr��ܰTo�<JC�"W(=��	w�'R��!�$ބF�^�R�⁨f�Vp��';�Lː�ȹ0�\��cӔ1z�!Z	�'����ݥ!����()0�'��qWI_�\�X�xT&Q�AP�'LȔy�Ń'AJ(�+ի
O�m��'i^-X�*A?NR��%IQ	��u�'�jh"u�N!���Q���K:Q��'�-��eP�,�*���4y�d�S�'��E�%�!	J�@gΎ�E����
�'��q� �	�f�)&0}�
�';�8$��:ีC��΁�h�k	�'llHh��ǐKBz�hS }(�T��'-qt�������.�)�����'��{pl\-+Y&႑fR��|�B�'� ѵE<a�qCdE������'Ah����֦B���j.�*�"8
�'	�3E�A�GA���*}*��a�'���F"��wz<�bIFf�1y�'�-�
�b������6��$k�'�Z�����}r����.3��u�'?.��gm�Ic��:R��(?b0(��'�~�I�� '	�&�a���7�N���'�TyÄ��d���@��+1^�x�'\D�(eCؑ]�� �g[�$b��'�`��	� �T癤y�$
�'3
E����"�N���ϭ��!�
�'%̝z��6-z��@F��6�(�'
��K��Bea<@�6B:��'^t���l���e�(+"D@�'g&�z�)G�D�&@9��Z##O*Q��'r���	�9��j�ā#���
�'�px�= ��/W�%Ȭp���I��M�%�x��Q&(�<�"O`	`�.$��� �69�2"O,�5��Vَ�6@�?R�|@�"O��IՈC��dPR��#K�4��"OT�"��	%<�-��m�v;�:!"O�}���N��N���"O�ɖ�+/��A�)�8�"O
�(�!T+�e"���"&�%��"Od� %�G��ԩ� 	�
$�g"O� K&�B�%���2X�4�ȡ��"O*|��8AfZ]��.T�y�7�7�O���%K`��1�%]@���͓�9x�*�"O0A���>t��@�sK�"�px"Oi�f�Q�1K���`�י�a�5"O��#��&} �}:������1"O@��A�N�U&z��Yd��- �"O�x�Sׯ|� C�AɑZQ$�5"O0����2I�L|�EE�8u��"O��B
;Q�0`�R��HH(�R"O� 5��Ҫ	?4���킰[/��B"O��g��X~p W� r�!D"O���j`��tJ��ՊE"O|��@��Ikđr0�E�,��\��"O��g�C��(c��H�E����R"OhE�QI�A�x��d�"?L��"�"O���3�tmC�#y����"O,U���\(`��}㤡 �nƊ�H"OT
�ӔU;����O�}̠��"O�Ձfk 'qj�%��E'iT�ɒ�"O&Hڅ�:�U��g�EX&x�"O�TSQc�)0�N���]O}�=Ӳ"O�	@��]|�p[JP3cC>�y�=;�nU�a ��D;�͎"�y�j[�q��t1vֶ�|Ѐ"ǭ�y�G�Wn`��Q��qv�P$ߜ�y�$�CK(4���ơxFF�; K¤�yb��Q�J��I"`�$�xW�wWY+0�l��$��P��������w������.,Olm��!Ǻ����/O>Y!A�� E�&B�M�9�d<�V"O�͚Q �=PN��L�/���Ӗ>�c�7]BM�Cƍ=ٸO�����~�x��ҸP�HC�c�&�PR�b��(��ɴ48�d*!�'BX}�&%��t@>,D�X�9[��PD�kQ���rĴ���MX� �8D�"���!	:WK�.܆q�ôh�H��ڔrNZpk��.-ha���
k��F�Ԙ6���0f�Q�4-	DAB�h�Z�s/��cP��� � U�\�܀���İ*��F�$�,L`���5'��y�h���R�YC�Q�{�X����͢+���'��BL�B�F	?c�Lb��		8֬Q�*F 9���si%v?�� �#�D�j����/:��Az����<ܴi�ʆ��ē\������7��THvK��?��'	�\��X�DJ� ��W.r;v���`�%,��"��`�b�z#%Ny0�IK(U��JP�6b�q����7֠��@_]�݄創މ:�ݵ��D؍Ǿ8�c�J��n�5��Հ�,
�n5�5 PU+z⺍"�����<�v�ۃ� �ej\��,�����J�@�K����>I�+�1Z����`�� Kp4�2&]�v5��ZQ�٫���d�/m��xG������ n�Et,�rƝ�r=��!*Y��n䪦ᒾzk�}���� �[�	�k&��7�5{a���� ��`��!��OH��!_;mIj�P�Y�m�� ��=��6�
b���h7KF��A�kDp�8���~2��}�N�Q����`�l����~Rb�#'�$��yR�*$ͼ@.�"b2|&h�W� F(���%�A�-`H����Q�=aBe�aː[\X�r��A1��&�S���e�e�'�.��"��U[��̽*z����̓)�Z�1�됶a�ԫ��ύ�4���
U� � i#`��*{�����s�ex0��2w���D۵~pvL����<S�^Zx�H�(�� �HsG��:.�%q`c۳u0tг��5qF�ٱ��]0b�Ǽ�xQs'Ę�z@1s8h��@���rN��Z��/��I��̠0�*DX�/;�U(jL���ٺo3µY��ه��Q#ebG&@C�� ��O)l@A��X>I�	S��ˋ Gp���ԟ��@���GO��@�D�K#xh��<	C�)k�i����F��t��Ȓ�}�f�����9o��p7��;&�6��I�[�����(q���C�:~�v��E�X;j� �:5�X�@pX e��0u��4
�R�]3t �V^z)�l�J�0�U 8�^z�%{A��"k��P��B��h�r�'�������M�J,�����]|�1[h�#i��X�T��8m�j��5�N�P|��l�J��8bwn�<8��D��z��d���ɥ^p��!C�`j��K��h�$��5|�]�]Ҽ Z���M9P0��IĘ:�<�*֮�" H��CE *�T��,�c�6�I�z$@��F�U�j�D�]�
Cڵ�6'#���GЭ�F�ÃF�`H�M-ε��8ix&$��"liެ��l��~f��P"�F�9���N�hx����
"��9�ڣnoԼ��,Fe��H�ۓG�1�޴854��g��!�h�ӄ�ak���CR:j�ia���;Ex�Hf��>> !�gG�$�x��`m��s� &l|�	�wld��`%����:b&�A`��x�&�^p��ό,'n~��3��2�|���(�>>!� `h�#`� Ar�)ֺ����"H '�j-"f�P�E�t��1hJ<;(�Xb��c�Qjd���yDM$}��!��M�\�8(�siE�*U�G� �J�"��"̙X��U ����
�:!�$�t�������	���'$�!����\��<R��!~K �P�!�z���,O"���� �ʼ��2C����!E��	�H<9f��F���{v��2�=zV�@`���xt�d��Q��ɾT��*"!�sdT���$m���0Ř+!�L�@��Z�\X�f�����J��O:6������d}��j�.5o�]b��=�� Q��n�P�z#F^5!6 ��#h�yj]�&jD,7l�q[�w�@��#�NL����$��`�!j���?V
�T���'��|�Cʃd�����O(�*=��c90v40FkH�+���A�i8hd౧���r-q҅�U>�IB��qh�X��3T^���LB୚qM�%5�)s��? L΢=1#�|�rps�+�;@�Pi�/�������"�I/9�ؠV↥h�ͨ���"���ҳ�Kl.z|�& [;�|5!J>�w)A3o�I��U
<O �5#�N≫|���+��>9@�@;hW�R�4�b�xѣ��������|��L:"�VV�,���D?#"	��j	%!h��������D��
���ej
�i�p+�h^O�Y�`A��X�����@O���љ�k�����
�h
�����@�ҥ��X�Mc���
��d:� I �K�,4����B�'iJ���@`���B3��-�`X���ZY��[�7���r�G'lF����Pb�qp�W3ZX�C�bV � 0�'-|����A�)T'� �� ˔T�M<�@
Ơ�o�����/�2L)B���ΥdrD�V�Hn�� ��ԮO?�O�"�̤�Fj�m�(!��$D�l��͑U�H��� ���7W"Pp��ٝ\��xb�̍�Z��aF��9$�F�\�a�����b&m���'A�)X���*�@S�Q�XK��;$�z�5�B�5�
���=`D�1!�ݡ,�T5X��P[M��#�w}D�s, pP�������Bz=��'�~PAF���dZ���G@�>$њ��gA�lpv��(q� ӯ=�xXI��Lm�S���r��;H��i�'H
)����K��6��@������,+S*9$(o�LX���Ty\�3��(t7"���/��j.@� �8g	ިz�B�h�Tp���$ҡ������,!
X��`.Ρ"7qOjh87����@,�0W~=9pʇ�pt�A)�M��aD�wj9��.P�P<���ۚ%FZYS7���0>�e��h)�`Y6�7ldh�!�?U���g�U(s�G$*2�#%��M�Ҍ4
g���D��yGg�3W,��[1M�)o� �7- ��y���1���[�kOi� C�m�dT�,(�=����VA�1u�fAQ��
1���c��ϛk�<G-Wa]�0 #F�<:�΍p�� Uf<��˕�p=�4�UG��2edO�树���~N%���R.Oܤ���2X�7��M�Չ�
�y��O�,�R��A�r���37�4�\�⢊�(��'�X��Ҋ�* `�lμq�@�V����d�yȰ`�,a��Mp��=�LL[�f�'%�J�B�ꛇA��(��Zt��p���?s�X�)�G��ĭ	`�%?0��kw���A~L���0u��r�V�yt�E#Љ)`C��:;�R g�t�N�MI�lz	���(D�0��[�D���A	�2�Z�@�OB�!]�%��+�J,; lT	S�62��@����Iİ�\�X�/�� _�)����%5�ӗ�6�l���o#LO���ua�^��ȈA�^���fG�l6j�Y��	?b��(6om}&��6w���KI�g�������'����F�K}=3b%ܰ^��� ��1G1O��p�N�4J��t��!UƓ�����ɹ*�����[?AَY�Ă8l���2���l#��;���6N$d��F�;.�����B�1O��q6GĖᨀQ�FQ�4n@Rf�bx\@Ɂ���Wj���&b��agD夜FP�3|1,�����Y�~U�T�Vk)
���L~���G�A��ɕ�����y��w+�6�e�0G˿=��䘇�۱r��I+1�s���s�L}��=cW+^��M�PG>�M�Q�6c��P+7�? ��#Ο"�l�)CAVx���c_&�|�i3��k�ZlZ�m� C!��j����,���!ŧӐ)H�b+13�A��=HD
!M��A!��B�c�*�ꃁE��42�IX,�� ��)N���s�Ĕ�UKp��@�N�&��RAĆ@fHaj�D0��DN@
Lh�@���H��,����EV`�3���=����Q-R>-��m� �$?�@�Ï�h�d	�|�A�t@Y�*A��)��Wm��R��\J�}�R$��$\@�f�t�]��4oQ�d������)5��5&	��ʇ#K�U�`Й���?��|[򠘯x0���n�-E��3�'� 屳%I�v���'�	�P������?P��!��Лcx섀�45Znu�����0�!z���x�喦8p�U�Cf��X��)ՄXj�$�5��=�s�J���g�(n�\�ʀύ�K�ΕA���V1,�䅮
�� ��ܙcL�}�Cөl�V�L�O�ؽ	F$YT7"��v�D��4}�vDv%���r/V#�6#?I�i�6 �{�,M���,�dI\@�V�F��`����B��:�9HC��nA^�8V)��L Jl���X�0�\�ƄDe���t���	^�P�G��!v<k����W��2�*=H!���b�`���eˇ(K0�c�͒�<�'Z�h�D\�EHp�N��t7�&-Z#u��tE��,*ǣ�9dԨ�9
�{�.Q�E�Ke��q��gD�����^������uD6��M��֠,9��Gaf\X����#HQ���e�o~r�	E-�)T4lc��� ��>q�'!U6KQ*R�t9�E��W�dP�	#�i(��k�t������ٕFoΈ���J����M,YD�a1DfM�K�L��K�Z�S��tԄ%�gf�Q�'Z�4V"D^��,�>6!�LCe�9G�� �T���Nm�� D&1��oZG�&�8��+hZ���G�v�!�I@�����xb�&B>���M
�C�գǌԻ��D\�oT09��(�?c��My�j �$�u��E�I������&�)�	D"�-�gkX�:�����͙t�^R��{����sk\��<�w�	%B<�b[$����I�.}��pb�dR"(*�y���[9i�H��׈��O�f��5O8tG��(]� !�djR�%¶�@�CEGO�A��̏R�ar�ԥkL�d�� ������o�@��	�+�8���*+i�M���a��p�2��t �r*�nئ�z���$=Q�$�g�D�z�ƑPB.���#ϖ�'X�;�ɰ{��S��O�]��iAe�1�H�0�@{l�����%: s�OAC����G�jr>�Á��`��Az,�N�h�������I�X)#a�<q�#�$Jj�,�K�z����7r0�lZqWF�F���G�n����4��B�����B�?֊��(Z�K{��x� ��%>��#�X`8����&"9��%Ѽf�n�#�$	�<5nHj"�oW�#���>PL���s�$�M;�-�{����*�tp����ܦ]�(�cfJ�o��Ez�A=��i��+w��y�S-!~X���-�	#��:h����g�^ܽ�7\���v�H.&vD8�% \�+�,I���8l���2��E
b�ö�9=2xhB����=q����1S ����� F.*8�I`�Y�0�#�� fpyǯ\�AȀ�!�N�E6�@����u���Ĭ� 1�Ê�vPA�O��2�!�;n�P���T��� �'T�s��Gq'h`q]7)0̑�kP��Tء�	YZ�#b�~�M�!,Z}����֘mEtL#��ÙǪ����
y�v���ƶQ:8���ɹ���A,h������Kl;���0�@ j���ViI9:-������;�<���@�i�������m1��Ӡ�!� !S׉��[R:�����	w7"m�ŦP�t�ўx�����v�D����*��X9J�=iq��waj���d����ʅ��B�
�f�LN���l��]�1I�(D*ref��d$/����p��D��
U�9����R���S� ��l����4�j�/_����v"�,�
H����(u������D�@�㊷yZ�]����1A��a�qj^
5>�x�W%Y�;mN4[�h���,]���2웟2 �=B�������-1F���4eؓg�!��ؘ-:�R��ؾH_�1��nK������5L��řf��f�Y)7(@�C�n�T��$U�Vf��%���W8��.,��3*G��������Z�@�ÈVT�e U��@�2AH�"�#PVT�uE��Q�V()S-8B��PZ�EP��D�F� i0qҡU\L�xUe�܄y`���+N�X�Uk���"����ɤ5��@HP�ؙ2�� P4is!�3C{`U��(,@T��&�t&:�j'*���J��̝`0�U���Gqpq�"H��@W��1V�p.*�ZD�WLS�AjcB�U���%{�m�4Ii�](#J�2�ԡ���8��|�d��3�� ��'� ���
�Kg��pME&;�A���$s�O9ћ��0-^�!�� Bel�F�ô����Kz�KtިS�
�v��m�A��mX�l�ħ�9�-4GK��
��f�N�Kuڤ+
w��I��A�kV�d�$G�&�v����i~��� C��|ʡMw�����G0�ў`�R(P�;�h\���_�*��%�Փ�l]�D���$�
]��mR�Y�D9̗�Jl�U2��^�.�M��z�7��$HB�jTȨc���2i��T�#DEd|Gz��)p��4�D�1�lE�� '>�a�� ��6��S4���z�(��Lϐ,!�+�+	0G4:,��ϒ�{�����O�ct��|�O<���5hyz g 3$ā�D�Ц]�V�"J��i�ƅ�3�bCrcGm�<�t�Cc@�CٟkI&f"L����O�X`�c�ǂP�B����"?LOr=y(ɷKE��I�6���x��גt��T�đ	z��8)��_�2O��%#�V��&	m�|�q�'�6ݳ�K�%E�pB珚/c��Y	�_��#2V�~<�a(��L
r|8�50���у���!���� ��fר}S��
�?+�A���ŲJT��#G��:�� �,ў�h�l��H�Q�=�9 ʅ	�8�t΋�z���k �U�S	����)��Kⴀ��Ƹ� J�(nȸ ��)dp�	�ɫ
��\��fL
CH��R&G�֘��JN+jΰ$?�zգ�fD�#��-f�>�Z��\u�<Qt❦�
QaG���1#x�I�E&�e�7j�u�B,Sb��;���O팝pf�D���H�yqfm��L6�9��^]��~B�!�������`S�y��7��ɐ!��2M-�$n�:.��I��<1 ���}<�ۆ)I�KD���.�7@�?�r,��%�,�	�$l�*�'�(I���BNH�y҈Yk겠j�O�(����o�x�!%�G��0q��m���&ᓬ"cU1A�kp�A�@�@�)��C�I*6i�tx���v�����4��C�I�;q�([s��bt��p��_*%�C�	�-L\��J��`9���UFיF�C�< ���{d�ԽP�h�c"�W7sxC�I/0�h�GF̵�z���F�myB�ɴ)I�S���.G8D��Ջ��q`�C�I�}_h��1*���j��$�ͬl_jC�I1 G�T�d�_�C%��p1�K/���'R�K`��4a���R�����'��-Q�cX�FQ�}c�l
����
�'U��u΁Q<J�qQmȜ��m��'NmڒgHU�%�p#"O��u��'R�ނ�0���/G�E)�'%Z��p͇<.1���`�10��'z�$���$z2�L�M������'�t����MM�8�cԋ�r� ���'6Z�QU�� �ʑa��U�]j~H��'�
8��Rp* KK�U��H�''6� 	B9a�v���gɀ�l��ӆ�,�+��	b�����P��&�xØ�-h&lB��"��m�ȓĬ��1�=T�Y��I�{!�U�ȓF�J�d��0���b��J�.�H���]�&4�I�C�аRD�3'��ȓI�Z�j�LT�<�4�:�假s0��ȓk�zӣO�;�mB�=h ���U�d�+�o¾*�r�I�i�~&ą�g��D��� D�ؕ�r���/�Ta�ȓ	R�*��77�΄�'HJ�>���ȓ[�Z�X'/F�j  i��ȩ�~8��u�vP�0�ԏ]��U"���{�ā�ȓ+���1���1��J�� ����S�? �Q%�.
�æJ�-4�~5Y�"O�)�.�9	h(�+�
��5��أR"Onx�W�P-'��-R�i�����"O�d��JJ�� �8X�<��"O���F?t��h��MjAJTk�"O���ņ�S
����V��Y��"O�� G��y�<��1�VE�b�؅"O*�0��T���9%h
,�tܻ�"O���� �&���z�r�ن"O�\8@#�&X�vPcS��K����"O^qC��϶i3&"1�]�6mP�"Oĭ�B�u�����<%X��h"O�����T�^�y6��W0�3�"OX�[Ղ�g�,��ع0���.x!�� d=,��� j�b����şU�!�D5}< �G �����x��K_�!�X,z04��f	�j��fX�n�!�D4�|h󴍍#`��]� ��E�!�䚷0˚8`Ǧ��K������5�!�dCy@ִ�C�*H�-���_d!�$J %������'l؂�h�-BA!�dة<J]���ݹ\������U�/A��ڃ���p?���;�0���(�8<��:��OX�d�����Er~�eP��[u����}贌��PA�@"D�s�&�v->���ć�(
RQ�@�"}R�I3T��0��b�q�PU�`�B1vk6̑�)�,4>��0�)LՐE���8�8a����Y���'�X ���C�~-�tD� �;GHE�S؞�#��Xe�8@/����H�L��Y"�i tS���B��`����W?M �{eB	�1��Ѕ��a����۹R� �"�H_� dȒ���{���CEN�R��� P��y�t��7i�:T�(�
�����k�Y��B|	�+����@�m�.Fjџ�e��� Fd���6g����IF�V�uy��
Z���B���83hIQ%ɑ�Uz6�������#A�W�}iՇ�Y���z��xR*��` �<Q@�,��HG���D��������?Eg|���e�%
L�(@/��h6��Cd�G�V�պ`��%��Lb�'@�S�[�MS�~�z"�&BpVA>�����<l�2q"�V-��1�%І/6��f���Ђ#R;'��8�Pe�|�(M��莮_?<��� Xbp��m�N���jS*�*mq)��m)�F����'�B���,�Ovέ"&���X���!f둷�X�4'�a�΅�eMd�y��L=LwƱ
L�[���됵{�V����,�\$��@� ����N�/Z�>��E�/D�Ђڜ*��:pAų(�H���˙!<z�@hY�3�"dyDC�/��)��@W1���H��@> ��"�X�? n9Ӑ�	5�8P��O��d�5>7v=1��ۈ����O����ɊE1p���䎍ڈ|rժ����P�ƌhH��00�	�U�<�E��=���s�gڥXqN7�]lx����1r�}�EGs�&�ҍ�$E�w�n �bb�6dZd
�i
�_�FP;�,,����A����EN4q�t4���1kDX�I�-\�D\�;OY<<h�KƷ)�lh��舚&�ԭ��%C4�bt�
�&�޵�te��u 	J��R<38��6x{�A��59$�s��O���C�v��"0�I%2��L8u��tд��y�^9,���B�#��HR�<���G���"PfNUcj���	˝b_��	��<�P0��Jo�J�N��&�)��KE#;m��І�O�@��:�D�s�	e�<A	�#�5��4Hx���&�#s�lIq��U��ً�G	:b$rIח wxT�?Ns�����A!u�xm1��Q������N�6�yw�N��I��NA�GSB���Ru��H��鐖[�,!�E��J�&�I7鉽J����.��k`k�C�^����d�O�l�qjQ��F<~���I�I��������hd(#Cƙ[����tIO�O9���tI�7�Z�P`	� k С�D��,H�Nk���؛)J<�T�����m��X�*0HT��m��ׁ�,&���ɥ� @-^ �a{N�:R,��_�48xD� mġ�iD���ћj��4Pd�?�<��.�	(�|�O>����+�r���N�qHB�aʂ�H��b�V�o���fj��|�d�b��#yj��S-�k�8��ǩ��3�����:��ʓ}�`�z���x|l��cm@��M�É,.���˪k=��p�p�Pℋ
��p�2�[y�2hC��%O���[���,����'B4@��x�$�ɉ`~}@���vK��R�n߈�0�G�� %�a)��2 �>�V�I	`�����@���"�
5��d��V�9����!��.:*r�(C�i�8�
r'P38ҡ��'�b���6��-!u -��#\(B�	�R$mM:y	T�3_��9R�`Ŝ4� U���I$KݔT����b�z�C�;d�૒#\�=D����Ѣl0�u�+2��Xa���Q��0	��_��\1�q�4�y��'���!�h�n%�0!(U;%�|�y3�'��*tM�Ѩ#�6�1����'!�*�݌9b�x3�
5�Ak����mi~�Z�@�^8� ��5uF5���,FZi�Ǎ��~"��75�hc>yD⇶N:P�B�v��!��gA+dX�aDC�!-y�K^�|41!��K0H9rB�r��-�Qgr��!	� �0!���^ū��� ��.�|MpD����g�	%� z3!̑x��	�)B2?�8�p��Q�7��'N�� �4����A�!:���~���1�I�2?�<�X䮐#3�!"�N�^��ًa�ߊ*����䡏�#p�G{��׸}�p�w%~|8m�3��b���,1p�Bb�O6h����%�O�J 	� . 1�D�6��T��D���
d�c/�� �%���:d֢`y���Q�(���x�$G�@��ub�J� 'R�J����-Lp6���I�nt�D��C�\�c&��;d��0��6z��kD���`�̘����"|Ob��I��y�#
tSh��*�<<Y��a� �9��hGEV�*�h����Ȟ ���Kr[~��Rj���	(ՎG�1pB��I�}��XY1O؝ ���1k�$p����	I�x(��.�
�	�V�\t��t�F�i�H� �`ڰh�*h���^�H�r0��U���C�G��J����vLp͢#�4LOFa�6(�$�l)S�X��g�V��`c�A2sT�@%[�Vx��cաJ�5��a��ԈS\��0Eg
�R��@S�$]�8�#� ��fK\sq� �qO��(�l�M�n��� �Pr�Y
Q�
]�4���U�s���E�Ј���L�ƌдh޷8���d�����{�cΓ*�PU1��O0��y��8�4��-���$��JLBKLP���N�.�DyQQ�2��$Atd��yW�$u����!䴰c��yR-=�t������zm�m�'��*�6`�#�.xЈ��'fؖx��=-s$��O0�Q6�^"hI��]2kRM�%͔�0�p�+Y: (���կe���,ƘQ��		� 2#�Ak@B��F��ѱǎ ��ab�#�h*ԏ�x��5a0`p�':$���:/�]�`�ʎvV��"�N�#�rD��
qH ����:2��s�R�Kg��LG�)�����-@�"4�ռw���$�Y�+�a|2شh�,�۠f�� ʴ� jV�1ЈY�Vo��o��A��M��tQ8cmX4i���3I�)Ձԭc� CH���ʪ5>���Z}F�ȓo	c�ʄPd�9���^�0���11!�X F�b�P��o!l ;3"
Sc��,Z�$1��`�0u ��^Cg��G��0l'��y�'��ARWڋhu��a��B�sD�l �G��j *��w�>�w��p�x�Z0�i$بQ`.S�2�x���T�T
�O��c��76xՊ��ʃO�H=����J�M�F�`�N9��[3C�,��(�d͔��C�O0j\8����?P�!�3c����f�� .�6�c ����=Id�׾�*�Z��wR���/|
zU�kp�c�K��W�����' �?����80�� 8e��-| ,"�K��r���'�^�f�z�� :[J�C�4G���F�"4Bpع MΓ.2M{$.�9kN2ä����R6E�����D!2Id��p-/4AkY.J^�l��댂�v��pC I���d<Vx�W��'~�bM�"��9��li�>;�� �6ʖ�;�<��*��#�M�k�|���n"��� �y�N�8�������i�~��CM�;��		���9��!QoNJ�pԱ&�'�鏚M� x�L/eߞ� �ur�1��b���FmY�b���aw�أ�%0��ͭaא�8���5-Y�l�e���z�Zv @$ۮt�"�>Y��!��O �i�͋5,[�d�C�P��j� ��"ծp��E�#��Y	'L��b� 	=��-J���0�*d�$n�7���$�Ú[��]���=K�mYa@bI����>����$�4`$ؒu�h�C-н|L���Ő̸s�̀�S	0�ز�A�Lx�ĘG,�8��򥁉Z#�XP
_/�<�*�K��?=�I�NP� ����A�.E�qȳ� 5���*��0���>?�a��Ѝ�z����N)%?PÄ��AB�q�3�$@� �2͡��O?rL!�Jئ%�:�n���l���ژ!�(5b�`�%�u����3O���A�-�#f̑�.�t)ۄ� �&2F�݈#�Y�O��W�C#
���W�H |����	}p�t��)-Jz��Ф�Y������?�Ҥ��B8H�]s/��!�J�>P��q�X'�ơ��C&[�ةb���eU8��-]8{:Nm���^�CH�hVܲ��І.�L]�!U�QX����E,hu�.���D�;�	:mR��v!(�Xu���8!�&5�_��X�#D	 i �����V�a{�Av�8 �ꒂC,l܁N�-2���Ù���E"lؑ��- 2���Y�d=�"����J�cZ�U6�q����G$|���,Z�Bx9���Y}*D#��H�'�`�fa���a�ByZ�����f��(�2oM�g�����N�h&/L*��Lx&�JE����T��g��8�Bo�b���H4�>1H� bY���u!�.�^H�2��f}�,Ưy�\96"K5="�`���)�j��@��d)�\Y�c��D�yT���;���e��dU��a���E͌��#���Y
8��%˜G)�x�'��@R�!�*(�T�VjL�4w6YH���?'������j��p
��RG\�[�a
.&�@�V��$7u2e0�kW�V8�G$߲� ��H>�ra��ɾ�|A9�eY�"���s��ƖP��%dP��aB�\> ^n|iŁ�X@���� ���P��Z
�Хd�V��AB�U�&f���@��uH�ǃ��O^pAk�-�j��T�B�90��r�D�9�N�k^Vx�H�
	� �s�F�}$���Ć�$�&�� H���w/<��2�#�TZp$���E�C���*Qbž�@�ӤH�>	�Ј"�qض��$A�R��A�u��x!b^i��q4N�.,*����.O��Zր͒>z�̋Ň�#U�0��BdO�`�4��'-<O����莬-U��3�b�!b�BƅϬ^��䲂%<6't<��[�cU��E���}���D0�l��K^�J���f��b��M�:�h�a؟�(Ԧ��8=����jW 6,�8 �.>�>h�#�
m�hPӂ����ʃ�C;8����\
Ȅ� �$,��� !O�"($��I�A�l��w ܋����7�	'���q s*t�Z⮞�"pqd��(�Hb���/(�LQ E�����@"V0��#Y� -��
,�`�*2�'�z�H�oA�SR"���@�><a�/OLM��ރg�(��_�[#J����g�	`6�L���EBD*��� -!N�r�	�lK H��l�n�	ڤ ��
�tɺ��'"y#p�]�jw@�5&Y�$�4x�ӡҶ�ν���Yj�m2�C6?(ec��|���0�댰M@�M�f�&k����!]�k�k�Y���8�-Q��a|B/1m���g"Зk.p��l�8U\|�����e%�fmA0��I�R�B��@Lţ+�x��c�7t����T	�F�R-Q8_~0��ҍA|�^1��k +v�ў�Z$N�O.�hS��ߤVN&�2�j�)G�n�� "�8�M٨�АɌ�But����$p�l� ��	�Ҭp�W��6�p�gݤ��ɍ�Fr�I�q9�AK��$M �#����TPX��ݴfy~0
R�A�R%�Us<�aVg"!G2��aM�PYL�H�
���p�I�K�� &ֽ?켨!�A?��<�g���hr���.Od��Űq�X�i�����[�熼0M\#�T� �`���jK�yt�CCD�u�@�y��G=��!�G?4G�d���&�}jc*Y6�Y���?-ў��T�ɷC��&CU,挸E��v��#&�E��k"!�(U�CgJ<m:=9���=`!5�q�ӧ9u����SA��[�b��2e�Ç
�?f���֥m�9I�B?{w����'�*e������ݫ�E0�����K�5n����,�������{��;� �:Y��4�$F�*?rR�X�!�>UΑ���H�Nh�����U	$��kU���Z�����)������`&E5���B�GM�h�kP�bXJ�0	/s�T�f�J1�u��X�4�6�?g.es�e d,4�'��S�p��#z��A#�&�}P eF99�����t�'�&�@��'�L����"N3�P���"��q��O�?H�5��C��+Z�4�!���Pؘc�H2�`�2EJ!��]��D>I�8)�"PR�D��DW2f2Т�!�O8�A"jE �����ɯg�v���#�@$ri�4GJ���X8���(���2��|sT@՜w�q�c��&�8 "�IO�AF��Gؖ;���h��0��2wo�J-�����j���7�k��eYI���(�Ҡ�0U��Qy�N�"�NT���2�?a�/\@��q�'!�;+ �qS�˛=�����z\��ڴ;k])c��`�h۴W�x�D��*g.�Of�tL�^�i2�G+H$ZE��VEm� I��&�~��T�4IC`�TfL�^���)O,Fu��VBbT�§�H�6�
��G
ɴ64����-}���)z��HC��DE�υ�R���FAS�4�<P���[���S"��m.�rS�·=Ӡ-���<!9^̀��ҫ4�&h�3M�����U�i$��P,R%
4�B��ؑ���K�WB�'�t������弆2�K7J�,�i�h�;9�<a�΄�*���X����f��cI�0�J���i�d�jdb�=�0q�>��O`qj!k�QcV��'�ؗS���@��i/b��*(��4��JU5o�������(���B�Ut�1�X"�·������"ll�O*���G5�0=��kG D�3�G#)ؖ,�Ѓ�+�z�P��:Wq�<�BMH1
7��O#΍⣤�iG�A�A'm��9�΍�|�� S-��P�f9��,)�O��R�CY�2-Ƒ	$���.���e�?#t<��_Ex�\�B��^���S�R({�y@�g+�H��36#��h�\!q ���sM*�G{N��0����)�2TLȃ�	\N�6psOE
D�P�)�!bٞ��Mԭ:Ɗ�q�`4�O(�Ӥ� W�!���9U߮�y��'L^d! eܳB�&�sŭ�Vn$�XS��P�1�����T�Vj<4	Qe� 9�l �Ѝ�,0!�֕GWl�����X
�x҇l��=bYiDEV�=�������~�L�s�?k3�A�M���Wmd
�d�I�8 w�:>a���EZ�q��K�8v��j���|�9��.� ~���s�iL�"��^�eW�i� �'���@��?<F��:�eըm"��$UE��Q�'��!quD0�ư*0 �,R��:�HD�e}�hI�$LkH<���G�q�6Ɔqr�A�lLk�'�z��Y�O��m�q.�5�5�16�����'P���ė4f����fYְb�';rw$U�D����0샠e��x�'r����&]�O�\A��)Z��h�'��hJ���,���ST!B���
�'�P�giȁ--�|`���6��`��'��K¡Y��T$�f�//+F���'��H���2.�^�	Ɂ���'���P�J�&��)C��+
�̄��'*���B�5" >�a��H*<�̤�
�'��ǃ=^�4���i��A���1�'gL�XÎA�3ExM�gn������'��4�����L�ւ{^�a��'�HnZ�,c0� q�4@��G�5�yr
K�a��HK ��C�U9v�\��y�ˎJq$`��Y:�*h�5(:�y"L� �42�B
�*��LX�A=�y«�&_p8W�ά ��Pq�a��yn *m�r��	/|�����5�yb�L�d~RP�!��g5Q�m�$�y ɣ-U�w�W��N�mV-�yb�#�`$s�A��LN�Bq
�"�y�E/[&2q�m� y%���.�.�y�F��#M*5"r��&{�h�l��y��p�3��X5,g������yR��f�����}��i���@��ybO��2��y5�ItH>TK�E��y�'�N%*�ɒ�3T�h0��#�y���%ľ�B!�ԇ@qRDѦ	)�0?��aU�R�0� \ds`ΐ�h,�y���ԶvҼ���d�7AQ����ܡ�Q>�c �>Fl	��K�x<r�C�^�P0�I
�z�2d��}>�:���$CDz���Ň>/��E ��\+�?9T�|��` �S9a�HH4g�v�4PH����'gT�X�ۨO̬$>�S�4��W=�4�A����T�NY���'���[����d�\�F�̱�1*ޑP���!Ƈ���#�xቋ���M���A���AK�Z8l����$BO\����.��� `��'62)��L]:�\7�]a(�����.ZwPh�#^9TG$E�P�v��e'�6��'w����w�H�R����������$4I�<���L$5�?�Kf��+ ���':�B�[f%�ēOu�������S�'��=yd�֬"�T-�C�P��u�'�d��JѯSɧH�r���P{�r��̀R�%���i@�po.`ɧ&�(C���u� VT,@��"Հix�8��މdbaIՂAD?�C䑏@�N ���{���5�@�q<hA�T�>]�����^�$�'*�����OY(���K�&z6������4�u����N?�AͧvG�O>�� !����B�L�AZȹ�p��y���/�ا���,��HTb�҄�7�ǲ\B,���	�F�>E�6�,�����-�jt�̄\� ���oܓypD�
�'3�,��C	%�TZ��?�9%�PR�#˿
qOq�$��A�����X�n���I��S���gCE:M"1O8ʓ��M��'L���sN��U�`%�%h �W����ٴ��ɭAb�S�O�0<dI�,�"��@{����Oz`��<��O|(�����o
�T��@�^��`�'G�(AW�Ւ4Ş��6�$�
4��'8"u��b �,��@���t����'*����E�-�Db� \5eHu�'�`R���N}�����Jl5���
�'�lmɑ(����`�ǃ;�8�
�'�����gK!d���#
���A�	�'n����C� ����
�q�	�'7�ȷǂj�����>���	�'���ԡM�����E�D*��p	�'ob5It.�_�bx����$mĘ�'�-bS�^���`Sw�X��q�'
�9��l��O7$���;	2
���'(��0I>�j�%��"~Z�ܢ�'`EYg̖+,b�;��u���'�6M��mҥ2,EI&m[�g��8P�'��WlL��~�U�_�����'J� ���	
��8 �;�p��'�L�+�'#�8��"M�a���':0��0|2��Vbޤ.��q;�'mFqǏ�+t�~�cW"%�H"
�'k6�AB"2Pل0�@�J/��'�ly륯Z) (D0
�ǆ���"O�X��
�J�tВ'�o9��h�"OЍa�*^�>-:��.*�5�"OW�ͦQ� �"�Vs*y
�"O�$S����@|�Q�*N$� ȳ"OX��h�1�JU`��Tu��4"Ov�ɒ+�w��eSv@�1Bs����"O�(y%��='@��J�/� �@�"Ov�c�h�*b�T���e]2�"O��TX�;��q��Ȭ{V�|�"O��2��t u���U�Q*O��#��M�}/�R6C�-t�d
�'RF���  vzeb��gpƠ��'�.�p-
�^ϴ`[�#�'Y�F8��'��e���Z)���CT$ǦM��m�
�'��9�d"�Xg,�q�-I�M�P(��'N�m��-R?~� Py�۱C���"
�'��ty�D�EЂ��T�G:�X�	�'{����A�~_����\�;'* �	��� 2�
�Y'6Z��eX�Zl���"O #v`�<"�@��ǯ�=Hj(�Iq"O&�Xg�Ks\�x�D�\P
�t"O�A�����8 i��	�`L�"O��7(ܬkжs��и&4�s�"O�������>Yp�Ai�	���K�"O��+�R�+��i�M�%T��j�"O<��$�M9���x�,� 9�"O^�yƦ���|`�+�;J��cb"O�U`GMY�F,�b
:��`"OX����ʡ[~��i�Q�n9A "O�U`先
=��E�0N���e"Opux��2VV�وqL��8��8�"O�M��DL[�h;���4
�!b"O����kD1�^E�G��C�d�3"Ol(�W�Աa�����$V�5�r8��"O�a(w�G?S����Ēr�,�Xc"Of�􀝬z�Ӕ� ��邐"O� ��/V���Cq矇�-R�"O���\�T;h"cl��U���AU"O�����_4
��Iċ������"O&!������A�"�� �"O��4+ %^0�qϚ�Z"!�"O�����:���MD'eg�q��"O�!��ӟ�t�E�M���"OԹa�
�:St�kwꙐ^;0���"O���+�4ec��G��;~���"O���テ3��lQ'C�o�6e�Q"O��"0C�%:�r����^{���!"Ox�@�,� ��h��5�̐�"OJm`p�ܲtL�s0�Ņ,�����"O��h����L\٫0��)/��AYv"OlX��+��#p����L�6�H3"O���ee��\��b	�j�ءzg"OtՐ�nޠb�$�5˞c����!"O�Q{WD��$0E�I��̠Yp"O��`��"(��PČ�<B��軡"OZ�g)�)}���2�K�*+ٴ��"Op�`7!��5�@�O��6!!�"O^�[��͑wŤ$���{�"O��r�H"6�QY��;�LH�"O�\�2A�7R^�RơX�T����G"OAr��؀f�N���M�ms4��"O��J��nz���E��"|g�pR7"O2̱@��q\(��񏕁1~��)"O�9�����GD^����B�n}��2�"O*����[�],�I�E �~Ll�S"O�����OOϲ��&�X6l��Q��"O��BA��#5[�-�%���X!"O��A� BZ�ԬȒ�� ��A3"OD01b<ٱQ��/�&���"O�M���**����)5q�0�D"O���D)��q�<�:'K\<���jp"O��j��U�?���!!�A(a��4"O��ң��U4��r���xl�y�"O�YS�I�}	f�;��_�`\��1�"O`E��UGZ�x���-r�+�"O����V�" ��l��8�遀"O�a@�ߌo�V�"4��P�Wo�!�F�-!�$B3R���Q �^�!�$�n���7��(��4U΂�A�!�M e� 3�
�%3����쎻_�!�Y	�m��Kم�������.	!��_�"\4Nܩd<y�!�� f%���]!�|ԙ�唹hC�i�"O���7���^Jl�Yă̇['8��C"O(MP�J9@t��qc����43�"OBL	gčO��#Cp�qZ�"O�!hGY쒕PDGʄ8:2"O�006+�;H(EݒE�u��"OJ�3�GV+!��$��Ӳ��8@�"O�|(v�Ղ	�X\��%�q�Z�W"Oh���MK��%Y@dF����
B"OP�3��Ϋ?{���%�* "O
a��m�
A�.hт�c�\�D"O�`5�V��"�N�c���J�"O�Ap��J�'<� J��Hc	�YyE"OV� 7l�����hAOД87"O��)��	j,  ���,P���"O�-q��X"u��X��ݢ#3N�S�"O@ˤ��~#�ݢl���p�a"O$�`C�����c+\}�"OȰ1�ձD�J؛�J@�~,!`"OXTɳ�L�Pb1+Մ?����"OJ!�P��dl�����{
Y��"O�J���k(�{1�_��p�a�"O���4��EA�Yf�~��"Of���D��Z�j��E,�p���"O�P�����~T0�GP�z��pX�"O��H�-g��(���=F�6p�"O`,��K�K0ဧ�T��T� �"O�x��IU�Qj�U
�W��Q!W"O,@ȃNΡf���JB�ۙ��|�"OF��G�T76��̕Z���I�"O��pFHwO�^�D��������IǬ	�!�6FR^0S��+Y<مȓ�ri�1�5����o��2���+�y�E-x�ĺ�ŵ@R
܅ȓj>u��'o�I�040�̅ȓl��4��ZE2i�l��Iü���\�z,���U4��zt��*9�ȓZ ƭ��R� n����ťu�i����pQ���)w�@it'�"Ei����`��t؁d��!�\� %\m�!�ȓI�* �3��\2~�p�_.�ՆȓC���k��i��a��j9)]�5�ȓq��=�'ǖ�S��}�ui?*_�Ąȓ,9�� ��.܌u a��&��!��+��pZ��_;�R�xbJ�>y��ؐ�pA�}�)�M�&w9B]�ȓ�~�)�i�5��IK;X�0�ȓj��Ć�+��'��
J��ȓEt�`h��Ŀ|��#�� ��D��TXLP#���3T(�JV%2ì��ȓj7���%��1(`���j�Մ��(�k���.�#wW����$�Jm��D>���,��PX�ȓeN\c��
,RD!0A�?8�ȓ
���ʂEI#��h�h�$R��ȓ�~��c�L�X�h���ɠ
op���\ �� W�S-~��F+�_����ȓQ��`�MM%���PD���ȓg��ф
5D�RU��N�b0��,�ȑ��$VK�5[�,� m�H<�ȓQS����WL�p�RR��C�Y�� 4	p+�^�LJb"#��u�ȓ,��aB�
 9G"��Cz��0�ȓq�lZ��(�������,5q�	��S�? X8��>W���2c#��qL���"O�����#�!2�hǶu,�DB�"Orp���ܬrtE�6���/`��"O"D�1.^a�|p�g���%�q"O� �t�J0 ��I:I�z(�"Oޙ`��ɋ.��u��HS��@��"Ot�0g+Q*��A��%�'�*	A"O
��!�	��I�D�;}͚��"O��W��Y���"D
��M��y�"O��7����Iܢ���C�"O� +D��"��耂ވ9�H1�"O�$�7�Ĳ
��P���7(GH$"O��Ao� �`����GZyE"O�ة��Y0�dx�ȇV�$8ɇ"O��y@���47�AYF��yrd4p�"O����&m`��	�!b
��"O�U!4�O54����C*DUMx��"O������L*���iľ|�z���"O�%)!��@*�q筙�t�z���"O�@�-U�2P)U�� MZ����"O��hXuul�rՇ@�K2���"O��3��b#pq�,٣$���'"O�eH$�ŏ���a��>����"Ot�9��R51�R�����7���;B"Op%���#5��,''�*Sx�9*�"OPQy񉑍Ȣp�х�1�ȴ 7"O
��J�#!�*	��IW-q�V�@b"O��G��z �i�8�v��"OL4� �[���
׭#{^�P�"Oz�   �\   �  I  ?#  �-  �6  XA  �K  zV  �^  �d  
k  �q  >{  �  E�  ��  ѕ  �  \�  Ψ  ߰  {�   `� u�	����Zv)C�'ll\�0bKz+��D��H���b�fB���y���yfY$E+䈳k˹X��5�u@E�"lHn����r�V�<��l��"B���*h0�)ԪR�B�I�4czP�q��0�@ۤő4y�� R���1i�,��U��,=�F�����>d��)XB|$�)���%	�̟�J�P谆�MD�"��rB�>�TdXn=�?�3��y�*���9?����$oN��'���'�"D��ZI5��n�	Q�n)	S��a�bH���n6-Z�Z���$�O���ŌT�����O"��΢'�N	$(2?�8<���V�;n��O�D�Ob�D�O���ލ@:<��א1d%z"lX�g-����^'}k
pCpiS6�~i
�bz�\�'o��҄�	r��H���V��0�5�4��Ѣ1�Ud}R4O$�4��B� �lI3�@Y�<qt�|LZ��A�8`~ز����l��4�?I��?�������x�3tL�T����q�W�N%�qA�r��m�8�M�ûi��6m�O��m�5��`0ݴH*��:,���8����9V���p���@g[�m�9��$ܭN�� +w`Ε`v�e3�0Q�)�|N���Ю��D��k��P�S'��j�'ո#�P�7��ަY�ڴ�z�5�����[=g����Q�O4t�	aU�_�$)�6�i������'d� +`��]dIۃ�=ih�=j��nZ-�M�i�&':�Uh���,�J�ɑIأ3��Q����
���$�i�67�C��Ӂm]�� �cL"L�]Ф��	;�����G�@��9��0'-�9s�Ǽb}�ɱ3(O<K�f�e�0�mZ:>m�4�F��k��;R�5Ga�!/�TI:f��! �VQש3�M��E�)!�������Y��@�6.��?�" ճ>@YąՁlN츳���Y�R];P��B��'��O��4`��V]^��Ê��^�Rhr�XD�8h�x�ʖ�S�2V�p�����'%Jܕb$SGn^h�f�>e�hH�㔭c�&ab��	=�$hrL��cY��P*��{���瞃W�͊!̒�d!>ȃdK��dx��&�>F�R4��M H�\\ڵ����bL��t�p��'e�<j�!V��f]�_�őpMܟ����'�X�	����ޟ��'+�RL ��!f��e��
� isht��ɖ�M��Kk�"��5n3�hY��E� ����'�\6�˟u�0lӟl�'����OM��Ѹl���hWoWł�����C���'�� &*�_k�<8e,!^�P	Ĩ�Bܧf�d٨!�%M�=Ձ��}�BA��O�e���m���5k�0"PB}:7����K���6v�b��'+)��1g��:��*��Տtt���'��c��k��l �'���J'K�͠�36�`a���?	�����8;(L�&\r�\@E�
1H \F{�9O�6m��y�I�MÜ'_Fh�	V��IY�mф��4�ŵi�Z�P�	�?e�	�,�IAyBͅ+wj&��G���8M�'BG:}+�/.�\E�&� �{b\����t,��hF��DY8�lQ#�%FP����hUԍ�M�ڴ�2e�5'T� ��#W�;͊�'3�^���"�μ�GI��E�1q-N�X[֘�rR�M�CY��²��O��%�%�O�H�F�)
�!�?jx#��?q������O�?�O�� 4�Z�Yc�t/\*~ve:��'��I�>�+O �'�?�+Ob�vI/*n8��ȣu�( ��ě�H�R��'FB�'��N�T1�^�U���� �E�^��N	p��$%hС���DXq0H`N��G~���"x��ѻ �Z�l�R��L�J�JA��)
Iɓ��g�+��ʶ�E�{!qO�բV%ΰ$��pȆ���T�h���	�\[ n�$yEz���A�_7��B�:qB��#�a,7��d�O��d<�O4�v.ԭjh�-H�L%k&�!���|b#k�nnZhy�8/���?���OY<	c㫟��� ��?q�t�"Mi���?���O���n�N�Q[T�i�.�1�J�2�"0p��Mt�ax�.���P�べY@ ���kQ,c��Ǟ P&�'���l��}A�-�n?���I��M{0�i�2B�0f�ˣ��04@� f�(4j������ ��S2-~r��UL	s�ƌ�L1	$�����ͦ�i`
@��բb%[k����u����MC*O�H�I�	��O<�J��'?`�����g�� ��I>f����'��HÛt�|d�Dg�7N���6ǩQ�@��'��i� T�9X *3L�J=X��I�H�G�,���
j��!;��/j�)��P43d��av޲�����(#�N���N&[�n��c�c~2�0�?�1�i���c>i{ֻpk'�	�W��}��)-KړO��d*�	p̓ �8	"��\ ~�<12a�5e���'|�	�'���"�M#[��y��țv�'�^��'&^U��h1g�-Z$��e�����O����x��2���O��d�O��$j���48�<��w�	�2S�qPb ��@�ʀ�öJ{H���}M���?5Q �xDK���Ո����$�����g�)5~4R�L\�,,*t���[�Q*F�J#��;��+VJFyY�,i�)��A�:l`h����?
0!��IpuW� ᣀ�Ozb>�$�O��Φ"�۳�	��Zp�R��%<�:��O��D�O���"�3}rJR�hB�A�ȭ�va���|��Ɋ�M[�ip��qӼ�$�D�i�|�ꁡ����b� �:&��g�^�,x#5lX	�?A���?i�����?��O�������{��s3��*�$�sb�,ltz@Y�AM�bL�N�%CDEc�A�O�'ZzHy�#�n�9���"Rz�j�g��hW���ʝ�'�r�QQ���*�*�Pv�'9 e����DY���l�1D�Vй�'���?!�'�l�C�RD�$��h��dҨ��'A�HH+3�� ŇڃU�V�@O>�2�i��'��cE�~�/?�š�*��>���ӂ���P����?I�#���?�����ϔ@R�+ᆛ="��	"�Eр @EQ�')9�ūa�<L9z�Z��؏
P=���$P}��'�4oL�@[�	T?|$U�6���W��Y�` �m����._7ZT	��D��`��%kӄt�'rH���͉WF����ھ�dI>��?L���,9�B�I���Z������?iT��>` ���q�J��Ȃ��I�';\���*b�`���ʧ�?��(��.c�r�+5�:��	
�?���"	�R�F�d$Q�.��7P�CRAQ3"\^��O=(�k�MЩ?3���_��h�Z����b��7	Y!��O�G�f�K��H�e��T��ԑj�Ҝ�St�^p��E
 z���z�͝0l��B������M#��S�|�T�͂D>��Q�_�v*�H���~�'�a��@4{�=1%�T��@���T��hO��$AæY�ݴ��{�vIarȅ�Kt����-^��D(��iA�P����G�?��ßl�IEy�$\.p2< j��ٚ �^�R��te2uD�F�V��,V��;5V>��S�>*r���)���c�un��V��'|�l��@wP��Q礅�^�ԡ��ƍB���@�%MX���s�)�w�@Q�
Ռ4TS�+D�K��%�i���^"�l���?����{0d-Y�	�G����L,�&����)��NǞK�ZlP��O�/ت���?���!���rӈ�O��러ʓ�d�+��J��4�BB&p'��ӱI�=�?���?����$�|
�O�Vdʳ���]�̝�������E'h[�8�lѩq��qs��lz>#?I�D�f�|���[�	�0�P�i�z���U!<�h��ך?pU����v�v�X6�-�	:E;fH���bfe�#�a���˖��O^@l��HO������Ē\ۖ��L,.4(�넂�ҟVv���D4�Oxarg�I;%�и���Xy���|r�bӬ�o�@y�d@)~(6M�O*�ɨiڤ�` (!e��H�CcX.{�d�<!��?�O~�ԫ�.�pTaՀ˖�r�*u�?&��!楋�|������-u��@�'/��A�#�%K�Vt�V���p�ur�g�*^�j����DV�ػ�e߭n(CFO� ;���W�|"/ˠ�?Q�i(�mZ��Q2�I3kH{�[�!���%�tG{b��݀'�}��t<쩨�A�sA�O6�=�'_��vI��ZbR��e����8+�L81D6m�<��a�-&��'A�P>�K�& ȟ�Q�!^����RV�\�,��b�Nʟ�I/M
���֤6fp1T'�$(�`-{���h����O��-�լ�F�� �B$�uB�H��OJ��cœ;�H�� ��u�P�J���p!Z8�I?Iw��mPXh"���+����� ??�th�ǟ��ݴPP�>�ϧ^z\����D�!(�@��˛(`xч�Zxش6Iǘ6H�h��R�&���G"�'ڧr`�
�@
9<.�3�h�0��� �4�?	��?��Àm��x���?Y��?ٙw(~�X�k�z��Q�F��4-��y�dJ�<���:F�r�����ICV��cY?��R& ru��	g瑈.�Rж�=Xw4T v5�3��MEb-�",F&��8�'�{�4�m���1?�"�O��3�$47EyfcK��Ё&�).�|�`G{2��4'aLCi�p��f��v.N%@D�<�i� 7��O�)mX���O?�Sc�M8w��1p��"�B�T�d #T�Q`M��	ӟ��	��0_wJ�'���qf� ��G*Ŭ�����I���q�SV���dDe �8x3�]�Xӥ͉�Yh�C ��'�I��,M�N,��ߺ=�����+5�:�J#}�H�pWNNnZ���e���<q/O蹒0w�\`FƐ�k`��i2D�,[Q���T��$��i�2I�p����O\m��<�޴4e��[>�i�Ե�M#���y2kP��*���f�ҥ�c�L��?�)O����OP�S)�A#�UH4H9�b��t(���ԯ�p�X&n��ql�ycl��z��M����R�hehDE,6�\�s�ҝ�OÊf 1��B4QR��"��*��|!��0쌊N>	%�П,��4W�I�vD�1`o����B��ɺZ�J�O&��D�'X�^92��^�ђCԏ ��Ny��i>u�ٴ{�0訦�W0'Y\L��l?�n����iG�	�!�\�޴�?����	X3_l��X(E:��B���qv���n�i`��$�OlQa$`G�L���g�P3s�,�X�FL��H"��#<z�L�W �	E�(=`A�{~�JM�'����ؘL9�D��B�����2��~����WtnU í�(!>��ce�"���PBl��A���3���t>� % Ԩ~��I�+��0���ȇ6D�4�w`U�'�d� �Hvh�b2�*��>��&��1O|�pς�,�>p�PD�覥�IFy����6����'b�'*�I�bj�3�DF=Kź4$��C������*a.�����]�UM�09��At���O���$��@��]�.�jF �8ef����7�:5HV肴vw�A�&���
қF����)֨T���u>�
�#�֦}I��)�1If�p��`�X`�'<��(��Zɟ�'2��]�E{L�U��+M�����Ir�l+����	���C��%<�(�a�G�OZ����Y9ܴ���|��'��d�.#L�c`F�iݚU��u���HC�$EX0�'�r�'���`���	�\�'%*Ȕy�Iρk�!���N0 �;ن4�h����PgRPt§�\#q�R� O+�(�\� 6�a5�1@��Xy!-C%/��}�"��qL��3����[!W�f� `��d� Fm��z����,a�ԇ��Xq��Q��'��6-e�'������Y8]��*�4"����b�6D��(�.<�����#%�h���'�� ܦ���[y"�!`��0%`�/�) !�������'��	��p�Iӟ����?*�l���M�I��}�7&��2��1��MB���!K�/f�� �'Ł���<�΅�z,�P���
��)S�K	�}� o�4&-�0��i�6!�8���֪:��H������9�������MT�q�A!D����Ւ��>��;�On�	��Y0_<����	Q%���$!��|���'�(��Ѧ�,�$y�CÛw��(����d	�IB�Unџ��IP���B9T�b�&��]�vi�,h�!�'M�U,r�'��p#���h�8<a���6� �y�H�X�L��4�?}{�.�R��	�#A�Z��'?Y�O]�p�L��BђY#@��F��/���:�-�t뇬��t�����QD�q��*�$����)u���u���F�43�P�����+P��j�iƆ$�a��"OP�#��(���iOL�~�ɦ�I��h�VLH0L�x���g3Lo$�(#Jeӄ�$�O���Ԛ!�T�D��O<���On�deމ��*c-��Zbʈ�dy���Ō1\�tC����NTR����m�fb>�'�\yU��+�~d4��;pF  �,O�G!����=x��@D�)H�,b>�&���k݃[4�,��G�i��h�E��OF�q�&��I�����P��u���$ߵJ-r�C ���&O����'�J��c�Ҡ,y蝡�la�/O��Dz�ONbP�๷lħ1h`<��9&��%�uf׽#$Z۴��<A�{��1����Y�h��E�UnJ�4"�B⢰҆Ɔ/(���*��ԓ}L>@��ȇp�'ٮ��EJ���j���͉�j!̉��M�2F�ڤ���h�z��UĜ�h�(({G��
��u�=	�@�xg�s�J�.'x�(�D���R���I��MR��V�f$a{Q̌�`���a�%Ed��	�'.��k��<�;�ę�~�<�I>�ĵi�6��<YW,=K�v�'�'��+���dz:��K;+��'���#��'��4�.D(D	'r���AkF 0�&�.H1�c
U��i	HxQ��C�(Ot���:Jm�P���R��[�|�"�� V6j����n2t��$�:�(O.�S��'nn7�ay"K�Oĸ�P�Ǖ +���8%���� m����+�;mZ�[��2����Eߟ���Ǣ8�c �5$�t� U��OT˓��9S%�i��O������7�
�<<�0�D�=~�p��c����Ij'�D��N4(T֔���nQ��&	���Oh|��4*�D^ִb4E!>��!2����V��u`<�����/�� ���l�bm)�GI7�iϋz�i��\�@S�Ɉu�3E��I8����W���J��|>�8u(>4^�����6������;<O�#<i�a#&/������h���FRq�'�f7��̦��|רƫ{)�}k#	�gf��5��M���?��_
��G� ��?Y���?q��y7,ש ��u��Ѩ���2v�¢t��	��8p%�Z�c^����mdh�eܾ�6`=��]���"��(�V��f��o1���yU��h�,�t����WB�\	�`	Q���Z(Oj�J �'`��?�OҨR  A!I��D�]�9%�}9H�<9/O���]�wf��(νpuB�S��&U;��ئ�2ݴ�?�#�i	��?m�O�x��G��~Z ��D�lBi �:F	���'`�'!҆u���I۟@�	�~��)��[)=��00,L��ڬX�%Hb<qEΖ0Y���֨Y�f�p1�ӈ�*0�Dl%U�T� ߓK��`z��5I��5s�HƋ*�h�Yun������4i��TDxRF	�J�� Т/͸��X��lJ.�䓔0>Q�
�.��$��ϔ�{�8}xU��R�I�M�4�i��	lUJ5x�O�d#'+T	�ψ%;�4�R��,=z��D�O4	����O����OVE�	�ɦ�	'�D�o��I���0;����f׃F�6�
/jNH)�P�	������.̸9$��:qm̝]��d����c����IQ�w<6���Ȟ�o�X�0f����qOJ3��' 2�o�������h[p��	�6����ԁsq���?��ʟj�wNN�RQ�G�ro8I �ݨ�����.�Mk�C*tdp���B�6�Ek�ki	��4��*f�j���O��d�|�L���?)W��>Y��(��	`���I���?��ݎ� ͂�
��CAc�$^�����XZ�* @ʟ8|�,W��\9�P��������u'΍_]0V��9�Ny����2Pz�x�@�~�“	`�
����><�<\���JH~�a���?�`�|��)�<3�Zp#�V�q�O�!�;
̘)�2���Y��1�џ�ˌ��ۀgm�%�6O�T���

�m�6��O����O��1�\$E���d�O���O�]T�ܕ맢Ϙ�R�fɂa�`�@nS�H
^��Ө5f��F�+擱^,h��OE�c%Q�
"�hd���{w �u\,#�U�Q��|�\��w&�vX1��p�4Д�~
� �MY�>An�l�/^���R��/Z�'4��H����>wZ��d��u2�*
�'�Ji'A�
�(�B��\�n��p*O��Ez�O��'�j�A��>���E��6�� B�m���꥙P�'g��'�B��u޴�?I�O�b����*yr��V�Ti���Q!��h �-�D���r��:�Y�c�	F���S�j't�D�[#�d�0(�`��'"���C��ڥ��tB�.���O0it�Kj���{�Da�LJ��ń5���'�ўhGx2N[�xX�6��$V��y�.��0=�b*Pr�K�����)�J:<�%�R۴�?�+Ot��b��Z��'���� &9n��$�	 0�҉�D�'��ޢHC��'��)�=a2������'���Z�Ԯ
L���a [f���pȞ����0�(|Z#�f&��+�ȟ�{��PXB�z����.t�"q�'�Ş��'������?�O�!��kC7j�zi�U�����C��|2�'��r��1C�\��)�,�H���y��|:�'d���q�	M3���Wn��=�������$�A*��n��p�	h�t'��yB���7�l�RK�?(�:�P��&�R�'�fL*!_e�� ��&�6��|j+�a�E݄���H�=Ū�'I2?!����0̜�>x,�Sd�E�p��| !�bp����0bM\%��L�g~�+��?�'�i'F"}"�O�: "�'�0l�
��ϵ����'$b[�(޺=���ଟ�^^�*��&�8�6+oӖc>q0B�x�(�U�Z�d�B��W��O����O��D��Go|u[�,�O<���O��Dw�A9b�~ДJs�Y�rv��	FŘ�3k�Y�ǀ�P$���WtRc>c��HV.O�5Դ0�a�[���S��t�0�Q@������G��c>c���G@�@����:tX�L�O`�&���	؟D{"`ɔtuB�YeOSd�8����M!�1	�(b�͟��� �X?/�ɉ�HO�	�OJʓf�|��E� 'j )7/�� ���Ɋ[��D����?9��?�E��D�d�O���G����Q�YO��ń��=����@�W����t �7h%��ڳ����O� �D��� ���am�B `���D���#E%8�2���� ;���*P���O�,єb�73dXA��K�i�@9��cM��ZT��8PW�ԅ!@v��#��a��y�db1D��C5�[ 
����⦓�^�R1""�-�DLߦ�&���A���)�O� ��{�D��*�ؤy�M"9��'�I�r�'}b6�������<�$9��A����ņ�0�nT\��D4m�);ax2╣Bς`z5!�2[�&쨒�'8� �c��s�t��.^�Z�0R
Óx���I���'J"JD�Ì)hLH*[4[W�(�L>���0=���߬+4�X��?G�*�jd��T���:�
��X`; /��Ӯ��|��IXyb�ε]�x6�O���|��	=�?1�=�P�PV�M�he�x�4,��?��m���`�/{�b����S'x�*�2�'��$�(<8�H��Ŕ�KT���'(���am��F���2Z�3�>qJ��U�qX��G��-5v5�m7?��ş$�Ib�O����VX��.\+34+��ˣJ�!�䑖,�ą��;1XP*��Q�X�џ���)^:�"���O�IfKI#*p�7��OD������?���?�)Oݺ�߷oC�H�C&$%���X�%K�k>��5$C� +�H×R}lb>c�HRc�̻&����q��Ѕ�=%�
b"]՟�hTF�jhc>c���$�K�+$1��K�h%q�o�O��E���Iڟ`E{����f!�$�/���!I�Zd!��3s����PK���ĺ�瘪OW剒�HO�Yy����a��T{��|Ad	�d�i ��h����O@�d�<�|��)�"�(����\�5������=Z�@ !0-�#�m�4e�b�I�M��Xr�K�>�d��!�;�
��a �>Ad|YX.��Hv�@#rџ��`�Y���R�ݡD��RV���%�J�d�O`�8�II�O&x��1'�9D2œ��_��x��'(xu+b"�
q�����\{Rh�L>�c_� �'!��9��>��Vzx�$��6M�4UBa�фT��V�T���4�I���� BK�.~��s�ظi a��F��P�Ӊ׮h��$$��O�$J�+�<NԂ� ��	H���1W
�Q?ض����a�vԣ��{h�?YS��֟��	J~2�X�k��N�#x��	4/��	���O���D��&5��;�	5,�Ȭb0f3W����OR��㜢od L�p�WR鰽�Q�')�5lk�嗧�ɸ|��N
]�V%��m�0�ȶ��:n������?Y�Xd-�%��/���&#�.U��Jm�6_38"��*�̖��"P����H�ET6L1hݡ���[�z}jF`�k��%Hv��$���DZ@���'4NTS���?����d�� .h�#�L�6e<�p�H�Pn,��"Oڀ��E���A5�!_^�X����h����ƫ
����Ĥ_��u�'C�\K��4�Q����X�3>q)do��c����h/D� �&�U�YE�h���;��=�D"D�����M&�2��;7j�`��>D�@��S@DD�3���0-�ҸX�;D���Xtu��W�P�Hb����9D���3�N�0�$m�ĭB0Xgd�����<iC&�H8� �U��"/�\y��J�*d:�X�5D����E; 9^Б6	�{�����3D��0��$���zw�B�Ew&�A�$1D�؂�jRl�0i�e�B,S���s"K.D�\��ő�>��|��-r��3E,�OnP��O�u$���e�� \� :�Ҥ"O =��.]�Pnݰ�*ǜ*���g"O�����)��l��ٞw�0p"ON=C�I��#��Dx�hug�iR"O``"	G0D"V�1�L6`B"O��Z"̎=
o�ɰ�L?�PZ�퉔FLh�~�̜�P�&�T�C 5�`bT�g�<���44�\h�˂:5	�u('
d�<�D�N	_d��ɡJ[6[� $x@F�u�<V��es�d���3+�Y�`�{�<)���;S�M��(�0uތ�#��t�<�e�
, ��A�#CL�U2����T۟<�`#�S�O�f�c�ځ>�h��(؆+ص��"ORW)U����٧$̲`"O���-u�~L)��ޮ	|��"O,ţD��N����0�<� ̩a"O�S��٠U0�3CH:%�JY��OT��#jL�����F�U�^�c"9�>ʓ]p�kN�~1�
�d�?�q%���"�;b��`ƴ�����3dϓOty���?A�2�t���?8����F])c��1"c�� ��z��#�^$c���%IC��WJ�q�'��23�<�J�f�?~$ޕ�L��=��Y��mb�b,3�fOGL��y��^�'�X����?���T��a�|��u�)��1�C%���D6�OP)�5�!L�<sR���G��@��';
�\�P��âm�����!��}�'��P���'�R�'���M�4]��ş�ڀB\�+d��肕|2ԑ��B�8 ƈ��n���%
�9�����P��<��.�U̧"W$�a0%E-{X���H��}�.<��Q�� X�dDX�P,W�0@3I���>�k����T8	p�W�����w���PI�O���-?%?}�' ���Fo�L�"��@�O"�p[�'M��P��� �d!��J$0:p��d�l�O+�T��	�D�h�8���	,T�c��'���'�:�;q�\� �r�'���'���'����i֏#~����-�}.M�S
�'e��!�߳2��̐"!ޜ���gby�>ق�$L�Ƥ9J�>J������5�|����@��N��T�V?��OW���O�v���/{���Qg��R�T3ՎT��	�\����O@�=�'�D�iAj���pЋoJ����'y�q:EI�7E�L�?s&��r�,k�������'d���ʓ8^�*\R���{b���w��1���5�'��'���O���'_�ش#��1��-Y�!z�X�$�-�� t ��^5[�/�	���rs\���$����Z'�#i-�pSc)&dsR��F��.��҄����`j����]`,]���$�������+��O)q4`�EGć5��t�'��c��YIm �`(�@:f�A�'E�}�qG� T���ꍧ2x�b,O��n�����'L�So�~:������G!/_x���#}�l9��%�?����?Q���?!�iJ�m��;���G����� M<t�x�3����$��J-9Z�P���	�<�TEy"��"����`�N�;���I�
�T����¦e�L!K.�)���Bׂ\=a��GybfO��?�����O��Y��L:%Hx��L�;l�P�/O����ʁ a��eeY�0G��1�̚	��}b#�<�! �#_�:Q�2�SCM�u���iy�F��N�7��O��D�|
r�;�?y�wvq����%'�<�"�2%�~��|V0���~iz�H��^֡y3D�NB����t P�7�pu����"��aQ��y��Z
^���S񬙄$�fH8�&\&��u	5�oܧDo�1!�-8p�آӇ,���ΓQ����П��䧆�� �Y���V�z�KUĖ=
h��"Ov���(N<@��˃G�. �p�	"�ȟ�BP�әG;*�pNK";a����O
�$�O�3�>}����O����O�嬻�?qV�^k}Dȓʝ: ْC���k��5a����y����cـP�͟����)��	�j���ˢ:g�B��:�����ᑴ{�bТ3��t0�U��n3ڦaB�t���'���C���v�l��
�j(�O&`��'r��I�<Y��_I�L�q뗕I����ab�O�<�K�	0����BҐ]�5�����q��4�J���<a�!��K��d1�&·x��1ۓ��a�
=�3 �?Q���?��9����Ot��g>�R�oC+y�%�q��:;�͑@ȇ�~��	��ʋ��iФQ�9�Ԛ���Q�h	��;��saśO�D��@	2R2�!""��+E�PwK̿xF�P �݇LQ�`@���Ol(�E��.\��KH#8�����g�O�=���d��N��Tv�J(I��8�r��,o�!�䈴;y&��O��?���c��;x剁�M����DYA>0n���	�|ҧa?fg����G]�G<1YcLʟ�R����0�I˟�pU�O3L+.8����Gc|�q�J}���\�ź�лq�Fś�����j��ڹb׆�3d�ڱh|����E�%Xɀ���u���ʇd�>�y��͠.�jp�.�w�/�b�]���{J|*�
�ZeE�Ԩ֌$�`�і���?��������ɂ׆�SXT�XW!
�I�CDEY����%��&����M{�i׺� ���]�� ��r�(��'�f7M�O|�d�O��$�Ox�$�O���d>��f��:7�X��nF�Gr�Yq`���8�/ݱ��'&�#=)�DӞ+1хfH�&I�������'�P8�J<�q��Od�'&'� �N��y� �����pD�����i�R�Q�~��I��"�'��4�'��[
�UBԄ�/\ Ā��$;��f���D
���$b�ఴH�?7�� ����y�(�>�%�N�u�D���#b��1�	ןXWh^�<Q^w���'V���'��D9F����G����e�m(���k��'I��W�R;O��؟�^w6���d�P��f�$ex��Y��*2�����rk�h��ɟ�"�k��?	_w��'��T�O����V`X�s� �`�ɻB8�("���O��#��'҆��D{r��O�$ڐݟ���?��kwefO�-���Ə2M���ҬzӪ�I�@���O�U�W�?���˟x�S�EWNtʳ��>��y!�Wt���%��<y��_���u��'��^P�ih�>���˕"8A�s+Ő`�y(��K�7��Tm���?	� �	�(H`p���f���OT��9$����^�XL��؁JǦ���Y�<1��3�Mk��i��4�'��d�T{
�[^�t��iH$��huĂ�):7mAi�<�{�\l���:�4LN�$_?y���:-���d�E�=@t�+�i��x11�'��m��B���`��ܿ�l`ܴ�?����?�����ٟ���|��4Nzf��'FG�U�vDҴF�Zw�8n�ǟ�IΟ ��ן��	ß���ğH��Sp6� �.��]H�$G�inşl�'F��'/B�'��W>1ri������D䙩T � �ʘ�MS��?A���?���?!���?!H��Z�E��\B4�sP�Q�nY0U�8��Ie�������dD�d�d�&��3T(���'��]�Ė'��'���ԤD�ؐh��O����*V�|�� �?��OS����S���儦tΨ �'�$ #�U�uk��t�A�-��'�� �@D�I&RlZ���&(Ӕ��	�'��y��Kb�"a!����L 
�'6�̨g�
��1P����J	�'.���@4�������AK���F
u�Y�Ǐ=Ry�]V)��v�B�aF�w�Q�ɼA?��[4,�wL�b�W\H<� � �.z4Q у�"E_�ı#N�C�p��`���ı���~�01�BL=l�P(ȍF!�uH��YlW�8��䅵��l�T�Z�
�%a6$��n&���C+ÛrIV�	s�TP/:�J&㊫2�
̉���0R�h��\.PD9��훹#�����R����V �2-��-��beNK�!c��D�W�j�B�rӰ�`���<\�~�*!�C�|�(���ɟL��-1=��	Y�S�,O<2�h�LNN�K����4�xBȑ�O���Q(�$ޚ1<�r��T�d��x�"�?!#�|��TK7�<�*"��;W�Xe�H �yI�"����eE���}��"T��p<��I:Up�m��a��b.�}#CWT��<�i�"�'��!�tX���'�B�'��`���X�ϟYd-��\R�,�	��d�d�ayB�#G��*�JT��X����'H�X˓HG�D���U�OHz��نd�RԈ��,�dهd���L<�MU�s�z�@$U8@����H�<	�,�M[h�0d煈S���A�FB�$t���D�x2.���Q��@;�����ȑ ���q�LI$��O��$�O�U�;�?�����#6J\���7z�p�O�$�6P@�'�� <``@�,|<�e��ꅳr��q��@_<Y ��E��Z�"6��Lrą������p?q�(L@N����U/,ȍ S-�x�<1� ��{Gt�rA]��p���x�9����|�ӑ,l7m�Of6��Qa4��T�D����/O�S,���I������Ο��I�|��hYӟ�$��bg�zRD1E�- N�EA��",Oz�S��L��1I�K �<�ub��9I�ay�� �?��>��&�?)v<k�W�0�a;��M�<�3�J�oz��`�Μ'%́ɰ�_(<a�*�ʈq�u�C�T���l�W�θ8H>!&_Q��I����Or޸��i��Q#�Ej� $�@�	��lB	�O��Č{m�ԘJ=���B� �?�Oe�]\hJF���x�񍀡:N
O}��d�tܜs$F?�E�@V8Xt��Ž�"�Q� g$5�D��aȥK��U�I�+������ܴ�?A���M63N:�xO˰I,-�D�,��'�B�	B}�d�;e�IҢC��-М`jaB��p<�p�i�6M)��� <�҈T ��e	r������4�?���?�W�ƁK��I���?����?YYc�,�xa��v�Bla"R�><����"�	i���$��A�A�CJ�#����遗45�O����'��I�D�d6�)C�F��xg���iI@�I�zg����xB   @"�8HV�C�iF�=�f���y� �+0hm��,�$t�d���P���!�HO�)/��4l(���_�}�(eB� øQ�@Dȅ
S2������I��$������|�w�X""�H�(c�W�{�bH3-���R������P�d�7�����H&f̴PJ�NL<�$e�"x�D�p�Gt1�9�3ևp�1�I��p?g��'O8Q�T3��0r�g[b�<Ɇ �"���WjO+`�h�13��Wܓ ˛&�|b�K�P�7�Ob6m�4I(�X���\*|i"��[6&�I˟b6jV��I�|ba�9f��B&�<W��h��R$Q w?6�c�)�oX��k #D"4���"E��i��DA%۔�L�P.I������8(8z����rO"�?}"/E�n��Zħ�D=��P�m�(�y��0T����*�0?ײ�`V҂�Px��/8�m:��J��ThD-ȵpՔ��|R*Svז6m�O����|J���M��
�4�vh���U����A�����'i�9ˢ�_b�����.�.&���T>��Oڮ��c]�[��D��K�"�6!J<��O�Ne�;�◭#���Qz�d��O?���V2#U�h@fQ\܌ib�'�ḍ*�R�.��	�q�N�fHDk
�J'쏿6!���4���B�c[6k� ` �/C'�x��:ʓ ��䐳t7��Y�U�[�Ќh���>i���?��i�]	��?����?�]�Eo6d�F��&Š�rM����dp�M�z�`*���n|#�(C��韀@��Ob�b/,8;����KJI�m��[�>��գ�eM�\D��*k���J!����iڎI�D�ϻYfQ�C$_
O���`6&PU[lЛ�/vӨtm����B�ٟ�	�W�,O@��4 �+�K�J��Ѷ-ȂX-���*O#<���/ �OX5bt�U�-�B�#r���$�$�u�O���!�	by��'����'��	�lw
@	2vs�%����� b�-+:�䈅�'2�'�b)h���	���6;F8��$��.I��K����:�Xa �%ur��ȑ䍬��1�/Α"a����� �,R��q ā�.H�L���,x���%�ׁLD�U� �n�΄�۴k�.y�Ӯ���j�L�"��:a�D�����X%��ǟ�X�4)��F�'7�Iٟd�	c�I�z�f�3C�ر҆���2%����?���/۾@�2�O%¿i�EJ�	%}�H$ۑG�
>.�uP�n�<)��rԛ��'@�ɗ���޴�?��4_��=�E�+u��h�"�;��4��'��A�4+��'�Rk�1O4�aj�y�����tN�b��*U��P+R+,O�iV��+e����O���)VE�vjɠŉ*���vo��T1axr��?Ƀ�i�L�	7�9ق�P9q4��v�K�����՟(��|�S���P����X�Ob�A�	Nf��pH`�'�r�'��Ͳ�(U,B�&1
�Ǜ�S�>����;�\6��<���I����'�bS>��!h��!x *�?i��(C�.�+q!V�O�?��M�(s��p�<�9�i��Y>�O�a��L�3?��<Q#G�?���(O<��`�VR;I�+����q�%��f�����e��,��mqםxR�˄��Q�Qyr��^H+�l@

0B�nL�z����;}��'��Q���	���I˟H��R�<<�
E䇷�`H.B<�ּ&�����}������<A�4k� �R�O�~���dM�;�I�fnӈ��O���en0P�%�O���O���w��٩l��j.��3��L�H�ָ�.�z�ȕ�� �%J����� H��c>��O��`$���w� �'�����]G��u�r�!�I�2b ��Gx���ҧ� P�t/O:
.��K@�ԙS�$��"	Eϟ��'�I���|�����'��x;�g�7�E��� �2�J�'&H��GDC�m��Y��U.`Up�K��Ɍ�4�\���>9A�H�KkĄ2uJ��Z$\�������l�g��U���'J��'j��]�L���|2@kݧ
 4u#$����xAW��kw��F�,q2�\���G�d�ɕ�����-*Te�,y��8�� l��8��/��t�P���ë6�����@�<�t-JW�"�F�T�r4#Oi\@��@��Ҋ�KvF����G�4�R&��=؀��w�ӛrü���<X�X�G��!����_>���=y%�i�'h�@Z�j`�2�l��P���A�.�LٴRq�i�׏���I�ZE�a�	ğ��'b��t�U�kQ
�i�'T�i���=:*T��1�� 3��}
˓Y�8��e#5���b�;=�|	V�R+�HabIP�<i��PѠ��Y�����؋*TR@-}BbY J�<`0�F�C)`*s���y"�Z�2��3H�?�:��5
I�Px�B��#l��b�q=T�NZ/I���;�|"�Q�[��6��O2�$�|�`!��M�`���7��h�@�JǏ��	��'�^̰C�'�1O�<��܍o�l���nZ�5��9R(�T�	%�#<�~����� Ù08"�"A�� slO~TX%�'���O��X�z�N��5�z�#�@�7T0P�"O:4@L�+3"�p���ϊ9	.���'Q2�<���7�1Ӭ�,9(@=��J�md>��?y�s;��3���<�?��?������"�!P��P�ʉ�t5i@��YR��vg�a�^�M�5����.���߯����9v�*@:�ʉ�C�h�!JZ�c�fQb�L̿ZʜTA�	M�����ܤF���O逅�$*x�A[%JS>(�גP�X)����z�/a�x�dU�VJ��Y�nڀWtzT``߯�D5��ⓍD�8���?��j�x����>X��D"�(�?{��ݧO�QnZ9�MM>Q���:�ODɺ����^7`����V�枠��NT�9@m@�G��p��D��)�u��'��6�h�P�ғBd���cG�Av2��"#ߊ61* ��'�O��I������A��
_-MB��J�/�K���2	�b�8q�w�׳D�>�(��ɀU\X�8�%+�٠6`,\P����E�O��	&w�MѢj8l����� I#J�<B��6uu��`��2ü1saA�?���dB�4���Āٔ�it2�iI���6�-��Mb��+}GޑQ�d�O^��ɹl����O�ӂ�R��)�$��G��S#�ܐj�<���V�L�ayҢ����'{D�AU�@Ҧ�� �ց�U���U����j5*��W��92 ����'�JC��\^U� �f�ˍ;0�B���
O��{��K�'d:l�s�ʼ^8�Y���
�By��O~Փ��Z���D�'�SY�DmڱW��$�񢙐fl��F'8=���?��Z'W,��ݤf�N�3 �^al9�E�����)+d)H��B򠑆�M"ik�'�,8���s��4��N*-����d��O�Ԑ�b��AV6�XS�7d���J<a��X��8��h�O��������!'N�,�vP���@9I�C��������2# �YI��)r����e�'�pi#V� ?#���F�"��^v}"�'%� 8xd4A��'U��'�;'N���u�(s@,�*�*��d�Ñ m��E��(|�Nq�(@'O��?�N�$�"�uՊ�����9��b�A�(W�6m��j�P��A�Mt��C$Ȗ����
d~$��w��ɛR`�!ezBm"'G��d �S)���ݴ�?�����?�;��gyҿ��0�P�=?~53�����k�Ly"�'�'6ɧ��Y6�6}J��C(z�,����},\9&7O �$�a}rQ����?���[}��v��{�E�w�kNѬ\ B����1J�D�OF�$�O����?�����$'�^��X;�ܴBn�Pg��Zּ�����CF��$�C:n`�+'�OX�)�o�(]�� �'G{�胠T�`�z�ɉI.�T��G�:(�&�RA����|R�*%p�;7J� �<4����֨���K���fz�t�ę���+��&w�|A��ܛ	Œ� 2a�p>)K<	E�$(�x ��E�ZИgPܓN��Ny���k9�7��O�6�� ��d����4��܀�c]3�%�Iҟ(� Aϟ��I�|�����$�����O�n6H�z�#��Q�0�92!#,O�,��d^�w�.��A�T���c0�Gay�9�?��>�'5��q�g�89	����s�<�׉��I6Th��U�(�d��[D(<3�Gns�вb��zC.ł]�fp�/Bw�	�`pڴ�?a���)��8�7���J����"
��Qr�1 ����ԟ�3N�!���2#�@7z�d��!�B�(����~�1�J�"���@�4�\��Q^�ּ�!�]�,sLՙ����vB����fO a��'W�X1�,1xf�)�(#�J$��IS�O��&�b?� l��c�V�a�9�ף <��]C�"O�QRWG9�@��D�@�5���y��'��<�2�����C�W�rM�����"�'B8OL�r����'���C�H�QS�e�5,i|9�cD��:R����y���Q�;9'��q�$�|��_�*�k\�j�b����� Q��`!A��Q4qZ�� ���T� @K*�A�O?%�"�y�������;.�!W�֧b<�x�4XT剸3�(���'r�i��]ڢ�C&s� �;�*� '�\
��?ړ��O�S�0��Y����\25�%�>��i�n7M1�4���ɶ>��o�N�J|�V�A�P�h)��5	q�`z�&�jDr�'3�'�J��ӟt���|Zp�|�p���be��3�2\�4�C4�JE��r
�bx��c副qgyyb�DKFX ɕ@������'x��H��Z�3�4�XmӅX�y	a�I���@��$Wv(X��X�c��"uK�Ob���	S���p��6�ZT+DG�3C�Ʌpf<��a�̧^o4��G�GR���ߴ��#<�Z��i�r�i�
�`�.�2���QQ�G�l��P��O���]h���O���,�&����݀W��%��O_�I� �ر	�`"���C�F��"�;d�rr�I�J`J����qĜɓ3�;�Lس��]�5�>K��N:�T�IP
�$,�2�#@��8 �2�ğ~�R�C,�`�P��;θ���ANg�!�a_�I��$j�f	J ȸ q��dV�/+���`ա+5�����N�is�"��9��43 �"�O�]>i����y0��d�*a�ꋗ[�4(4����?A��6�x���ʎ�vE�(!e'� |�αc�\?	�O�<B�e�t��Ъ��߰#��J<9gC�W_����_<x��L;����O͸� q�ZA$-��e���2i�M<aD���D�	e�OI��D��>G���J�5gؘ��ݱKL
C��8VR� �
ղ������d����'n�uS*�9k������b����6O����<ɇ#��B�H#������7��F����y��M��B�-/}��	&n��yB�
�D*LAW�N���q�h��yb䘆�2ɠ@Ϳ�Ƹ�q��1�yR ߵ)�
`�Ջ�&=��!���y�蚋0!£ˀ`�<)�K���yB�\�q��q�uaS%��:���y�;~�R,*�G\/|l���E���y��S���m"�
�)�ը���y�h	�
�z��E]�[�� �m��yb�B+V���)§qv���Խ�y�i�Q.��&DʜmL,�)ˌ)�yBI���$��M.������y�ȩ�\��� ,���{4H0�y��ļi��+Pc��o,���#$V��y����l,s��C�7]�����I�yr�ˈ�DA#*��*���CG��y ʎ>vEj6�<:\ˡƞ��yR�TT�*�kg�3(۪�H����yr��N�.�ѤܱV�c ���y��G/\��'������W���y��g�HI�0��8z�Ȅ�yRkU2<�B�a��6<���R��y��V$V!���ch�,V���qa��yb
X�T"�@I ��xw�ͨ�yRɂ�~�l�"��o�LI��D �y��U��A���&Zu��p����y2�"f����K�:����yZ) Z䘐 
�K���!%�&:+C�ɰs��3�X. X�"F�0#C�	/���@U X�Z���C'�DU�B�,Iz�D��/��T}�sdK�-޺B�I[V�[��@�8������a
�'NnD�\� �&j� !�ѳ	�'� �,޴.��iǢ ��fj
�'�b�(TI!@��ɹaN=��{	�'��AX���Hn�M��c�媴j	�'_H��5��H���жg�'S����	��� ��ڱ�צ0����b1	��`�"OpH*4�ݤG�� �%����Jk�"O@��A�LCm�YQ�[�u���8�"O��ѥ�mZ�|��@Y<�e9�"O�$8�j?���ǯ��W��-b""O�h�B�՜b���3윓D���"O@�j�a� =P�J�j)�*O\���$A�x�Ha����w����',�<b��,����tjRy����'�e��ԥt)x�ӆf֒Y�veq
�'D�0yVm@*h?��{����9�`#
�'wD ���K8��5�.ĩ�	�'9^�����*:���(
�G �%Z�'cn%QVgʦX ��	P�	��q��'	`]��ʅB#>㤇�}k�=��':Dk��c� �t��sR.e{�'��� ��R9I�~���[�[on��'cHܳš��^d&qs7��j6��
�'�44���	r��N[�y��'y������l2j�ĿUB^AS�'���Z��Cw�6��Ć��GP����'e��S�(ȈAx�S쓡����'Z0`�v둿hwd`��� 6�9
�'UX���'�m�E���?i]X���'�p���ŷ+�!�ǎ7iu*���'P<��S��*?aH%�F�o �I��'D%�C�H�T}����/X�/�\���'J����!HL	��@�E�~���(�'��`3t�]����pOF9ôe��'�pU $�(]ڨ1��-f�j��	�'��J�N>HZ¼ 5�p.yA	�'ì�������=jG��fbh�S�'Μ]b"�.k�q�D�ZL%{	�'�*س��}d��dA´�,��'~����=	Æ�83k���� �'�x��oE����a� �?Gc�02�'��#�%�
-F�s�曱>\*��'gi��C25�T��b^	�[��'�\��h�1�ƍh���� ��c�'�-�F�L�O�$��'�W�y�6,[�'qޥ��$��rόX;�ɒlM�Ś�'�
a@3��!cb��Q�F�j�N@2
�'��l��k��fJ�qb�9c�lM��'�D�dӔ^4B��FjL/����'��(����5J�V	�D4�踛�'��кӀE,���ԅû0s$���'{>P)���3@�$QI��̇%�`U �'ݣE��%P�(Dg[1?�tZ�'��	r�(< ׏Z�$ݲq��'z^x�f�o �5GP"�,%��' �����8;`��v��x��'���r������c"ē�]3�'��Mq3�T�
&�q$���<��'z��E�Zh�2TaER��As	�'������)��z1o��YFn�b	�'����hQ6�QQ�6P׈�+�'U<q;��R$K�4�����O^�9Q�'�~��5`���xr�e�zG���'����o�4AH�懎� `��
�'^��3�c҆Rʺ)��!��K�`�K�'���s���9���!A�,�PZ
�'PV,�ӄ=��)�*ΔN���'���!�]���9Q��)CÐ�B�'�r�#F]�R�a��V�@�:a���� :�r'�*T�J]2�E�Ef(UjB"O��c5Ά>,g�\d�p�ZU�%"O��/]�lH x�οl(��*OJl!�� i���q��(`P�'�vi٧�ʙ0:u�,��dSn)��'����u�R�$�E��<$4��'?
qj����P�sP��>I�
�'�R�G�í;�1P��B�~*8��'����fN߷(��z�N�6%딍�'Xt�1�eˬZ%��ɳ�Q�y9�'x0%E�MM���φA�y�'�h�F�$�T|��� �R�+�'G�9��3}d@�Q����M��'�>hHv��L
9J��T.`�'t5���-.����~����'d�8�7蜦��!+F�Ќ��pI�'yr%
�C�n���B֑8��'8D�
��;������{�*8��'�d���\�/����R�!�����'X�(���b� ��7��O���B�'� 4�R�P�|��}����
7�:���'�p٠"������:-yz���'u\A�4C@$����ɜ#M�]�	�'�* ��hϼ"mXRQ+,��)	�'�t5�qHW,M���@�;t~Np��'�rF��,r�lTj 
Úr%��'`H��!��2�L��0���[yr]��'5N���BR�uu�ĄA)X�t��'����ȸ
Ve��Ӵ��d��'��$�Ƅ���&���˘�&�Z]��'\4ฐ(0 8:���L��s�y�'<���oH�L��d(FGߍĪ]��'��$�E� </���@�7�(Y�'ͨ�c`�Q�N�p��'�֌
�F 
�'�h����{Ա0��S��dt��'(���&�ƮO�@�6)��=����'��u�w3Fֺ%�@�(�����'��<�a�N,]Eީq��$��U��'��(�����dR��·�X���'�.��E�;� i�#|y����'�2�Y�m�PA�a�̄�`�r�Q�'��i���)b�B81&�UB�U�
�'����>S��E�ǂFL�
�'����
��>�B@�7s䀠�'6��E��m�҄��%��T�m��'	RL��ǲC/0��A������'o\i�AC�M���0�"����ě	�'�X��c ק1��m��%�66�Ԋ	�'�8�"@N�F�d�J�Z&e]��'Ǆ��5�	�D���Z����T�D$��'l�X��.�v̥�BML* ��[�'V���s@��x���q�}���*�'��H���	�8�D�s/d]��'2�Z��M�YKN�J�M�x��ɚ�'h&I�c�N0k:$B�ıuq���'��lۅ���'̊tR��mֺ�#�'`쵒6蟸SL9��"�f����'�5���P�c||�P�g�]bt=	�'���c8]&���կN��-2�'g�"�/�HE�2�\1��+�'�¤��ʐ��s���-i�y�'������.k6d���'<���'����g��m�R�[�lE���\k
�'&��1�F�L��)3����{�Z����� ��Zf%WKVY:t�-�Ix�"O����l_�j>��*�!�D�2�"O�%�E ^Q�@11�?l��X�"O��oϏQ"�`�AH�S`J�"O8�+D�%vR3qBI`&�P$"O^l��n�8\(����f� w^��1!"OD,(L�W�:�z��#-�,�a"O�]��"v~P#0�-$Ґ�r�"O̱0�.�9o�X��!N�k�r-p"OR�BB��0}�y� �L�5�p��"O^m���H�X���դ�[�jEb4"O��i�])A��='�2T��I��"O:�Ҁ�R_J`��#"��CR�mj"O����GقĕA�A4&��"O|�C�L�S-��!p�_,/��J0"O��jT�RX>Rx%��%|�Z	�"O>�RC-=�y��ܼi��"O�ؓ%b
v���%���8F��"O����I�*�D,H�P�Bк�"O����˔=��D�7�ɧI��r�"OP�[b+��,}#��?���"O�-�eA�,a���ښg�:��B"O�,�`'^P����孍�Z�Lm0e"O\ͱ5%�>5��-��,�d��%"O������z��a���6{},��"O��"���>\����㊹f:Y��"O|���F:�c\4SK���"O,`5#92�"�`�O]2���"O�\J��;��|��Q2�*9Z�"O�]2��V�
>�11�.��6u�"Ohe�C-:7N��T��N��#r"O>�:�b	�>�����&��Zp��si �-I_���`@,(<Ob\���Y$��HC/��/�9X�"OZX"�Br�@�4��s��X�"O�H���2,�mJ�Í!g�H3�"O��ëD�Y��0b���Jo�y "O�`7 \�Y��M!�J�S�P͘V"O�qVB��(h�^�t@2"O�Y#FĹ	68�y&-V-{ӈ�)�"O�5���=e�@���˔r)�Y�a"O��� ]��
C�[��^�I"O���aӟ[�l���ҍc�:�[5"O�١j�<r�h��R+ІQ��"O�-c���1Z�N�3�t�a"O ����
�e(��d�M�82vh�"O~���.��C�<M�`�&t}Nd�#"On�:c.�� 6A�x��h�"O�y�-��h|�Fݺ^��;�"OD��t	F:?�����KNS�t9q"Ob�Z�]�w޲�)��ݳV�BY%"O�:FL[8h!�,���ߙ;��	��"O4@��B=Kp:�*�@��]>^�)�xR,�;�z2�U�Vhc�jŘC6@<�JT�0?	!"��Q<�0N����b���#���bK>��x�0�tӆ��#֙����HO�1����L�:�k��4�zGt�X��A�6�Č� X�S�|B�+�����(A��Y��hY+)07m� �v�!�K�S��McI�<���"w,��@D�$Hy�<q\,L�*{-BN��A��?�P�ҐWP"u��LI�Xd��s����GeBy�q���LHAC?U7a|rhR*Zb����蜃rk���E�[�9�7g��zQ�����B��&Wnő�d�� :�G���'�򩁒)� 1݈ͮ'�ٔM���F��3L�H�v��	H*x"�"O����&B�f�`� (6 8%L��[p i �f�Hn ���'B�>�)� �X`U& �(��[B	F��K�"O��e��?�f0PfhO�h�`|���iܰ��O�,FJ��%��x�R?x�``�C�(?RJ#*����=)�W
 �D$���Z�pT���7)-�hF�H;y-n�+�WEH<�e�c�� �!���*v��C��U^�gn�s�/������7���@�����hB�P���?="B�Ii��)�B���P��W��浒"���hڹ�MY!:����5i.ҧ�~��W, #���N< ��f���yre[s�����/�5��Г�
u׶0#㟸x�]�U����R[w�Q� S"(��( �UJ�X�@d�/|OD܂�T��!Q& S�[���W�!}�4͢wHƸM��D*��۾��?��BU�P��]�c��!��$S��I^��$��8�7e��!nĹDϒ�����=��^�7o��p�.ǚ&d�Q�D"Ö��
D=?М��S�l[,���Ĝ�j,@U���)j�8�ʲ��O?�I	2:j$C�%F�����&JJ�ZC�I�[i]��'Y!u�l Q��+ek:D��58��P��25L~�P��SD�'���vn�{)�,q�:[�\\�	�5������CY���!�<u�6�q���8	�ң	:�Px��!�Y�6��_�Dр�(Q=�hO8���i�V��c��)F7+�bAA⣄6v���´��8/�!���J*���ئ�kek�$}��\!-��lh#��v�6Hӵ��jjH��ж&�B�&>!�C[�[Ind�#�� B�H�J�3D�� E�@��������IgB1ꀋ�p$�D�3�9�.)�r*|���&>)��L¹P̺�k����M�IC�A`�ӦrT\\���������d���y ���E[�o��Y[�x,^��x���e��b�����da�+��c$f�F�*����5�n1���LU��q�Cӆ`c�Y�6�K�9��Q��.�m	4B�U؟�h��	�+�v���K�=]��ۤb<�h�ڦfԟ6���Pl�Z�6���K^E�|i�`��K���Bٲ�y� 
 ��r'Ɲ��b	�'f^�rQ�����8W"\y�,� �M�Sᓈ�����%���S��T��M�T�!�$�"g#���@PHA���+�2z��h�=��+ -��a��Q�GG���OrD{e(�6>�J�g݁G�n|jU�'����ȳCw��+�'�;c�8]�V���x$lHSIK�M�Ȍ����5O���dG�1��Mkģ��J(�8��ಏyB�O5���=%F�4��ޢ(l:񉂯$B�	�� 	4C��p�)�9}!�$�s���;�b�VM8����b5�;u/��CjV	`׀��(͛F�.§K�I�r��X���I�bmK�D�bnpC�@��ѲN̶;Z�ب7I�,6MV��tC;����f�����K�ܠFt��cBA==�tJ��7LO��0���qF��P�OW�f�� ��֙a���2eRp�|PG��h����I�p�tĒ�n��[ׂ�b��?��b��	`���L�	�IO<y����w)`ӉO�����_�4��0���&G���
�'.�h�c���A�p%צ-��h����pv�+�/�-�m��46M>I"�O�1�5F0P����!TD:�y1"Oj4��`
�f�.m��^� ��}��i�L��Hѵ��
 ��O7��i��D��?����5�\=ΥPj�':az	�>��(��=JL�@�F�
�dIȃ�1�dA��6f*D����"�O�T��i� ��p1,�2���$�L���EDj��A��7��N|a
�}�jL�VNڌ(<�$�L�<���U�
���P�ϡdh����L����TU |K���ɦɰ���c}��h:i:5n��R(܄ؕE�yr(_��a %�k�Q���9�M��O�#L$d�p��1*��9!�Xx�'�h�r�T�O�\p�瓸 �Ȁӓ�8��M�/ �@BF����&��*�a�$�S���.81��kڻa�a��"�LY4agx���D��'8����@�CH�!C�E��eS��x�t�S �����(9p�b����NB�Ip��4#�B)
�:|���H�'�� ���~�J9*Һ|���`Ӓ%D��>٠D�?,lX%�8�.5⒉�F�<aA�2P�x�i��1Qp�<����Z�<Q�h�5#H�a��h	V�`0r��T�<���@1˶��n� E�T���OQ�<��i��8a�%iT#	�-��e��cl8����Am�4=�d����;
��ĮF�$t	��S�? ��D0E>�rĨͺ$�H! �P�D�$��vk�c��|�N�xN& Y!��'>]�L��C�<!� �fLp��ʂk�FlI2Ǌ_�F�EWȌږl�u8��{��L�yQ��i�h�6~Hвl,�O�-7��r߰԰ OS�.KN(��B�X��Q�[m(<	�Xc����A5Xe�w��P�'�B*���'"��0�~ʀ��p��Jq'QB�"@��o�k�<���,>�3J�w�&��d��<1�� #��s#�x��	L(|�-�
��=^yq��=B1!���,b�p;���>D�(�cg_�m���&��O��A@g��{�����|Fx�)�kLIzq�N��"�ƻ��>�An�7�8d�e%Gm���1�Gȁ
-�9�Vl2"r�n�p��	���:������V �r�A5f�#=Q�@.Sx|�p#��N�M;Ш
S���1����I`#�p#E��L!�D�6�v��D�9�����ܵy�\c�aǿ
�ђw�����\�I�u�Ͽ�d��"Vu��!Y
7�~PIU�h�<�Ǧr,4�s1�Z,�<cǋ��xm(�BCW3��0E��6<�'�HOA����Yx5,ɒ�(���'�j9j�����=���E(��F��W�0vmI"Z^^�ĄP�/a}""�
��(PcN��#��@��J9�(Ođ�&*�(J�)RgF��cb�A��B�~:���7h@:3i�7�l4��cX�<��H��y�(`YP�yt�bR�����2�	%l�"hS(��
QC�s�&��I����4&/m(0.���yҨL�)K��#S!V�bY��ʷ�W7`�U��l�r�b�*�횈<�zt�����p�얕r'�IC���9O�(� 0�O�)� -wJn����:1s4��E �Y���{�]:NH�7O3�O���E��U�"�s��ƚRFq� 퉀(�r�lE�H}�5���t� * �mRc,T�N�t��Ӛ�yb��6����C[�FԪ�����~���^ZR4�RmL�t��)ڧM�J�	GbMWjx����"cv�ȓl7��+f�l*�j�m�)�xX�r[�0�@�������e�~�?�����L��.\�#Hdx�K]n�������,��%��<f*=��
���ʖ��{<S H&2���Fة~"�( mBi8����Nx��^���-��i��"�l�D%�ȓ[;�M2��.��*SF�`�~ �ȓ�2��槛�.�nXgOڻ7]^͇�B�T�R4�9,�:��1���cs���ȓo�nmFMB�1� ��V�34�%��J-n�AsoȮ��@x2c�p~x��|ڴu(`�ГJsĴB�G��B|��\(إ���&���Rf��G���M*�5ࠦ%f,ԧ�tXq��d��]:t���p�	��Y��Z�.��"-ViL�����!~A�}��6� �zХ���V�AЄ��~��ȓ�Ȩ���
��iQb�1!n���ȓ=� ���8gvY��Pj[�H�ȓ0�����ͅU,"=��;cNfD�ȓ���bb�>ɐ=	�Ί>x,���8d��{�eH�$N��T̘�uk���ȓt�ZH�>
l<���:	l��ȓ]i� �g�
 [��{��B]�x�ȓl�RɁ`B�(/Ľ+á�1 �L�ȓ~��8Jr��J�"���݆/vx\�ȓ9���s��񪌫 �c�����!���Ua�0\�s�"R��D������$���M���J���ȓ7{>���A��EGj�ʱnX
F~p9����,8��5zw�-�`�8٤9�ʓX�@u�ɀl��둊��BB��(p�$B�4��0c 'l�B䉞ar�����2�� -I4i�B�*,�ǆ����B��5C�>C�)� &�k��$�j�ɗdU��:�3&"O\$!@�Yw���J@:��G"Od"�HC������B�9:\z�"O|	��$E�*06H��.	5$�X؃"OLE�6J�ѐ���	�s�"O��p�N�k^�d)��@j�61��"O�Hq���g����X'�֬�e"OVT�c.�/~I�d  F|l1�"Oʵ�!B�d�B�"5�O=%jzt�P"OT�B�\*	B@	c�#۫O�ؘ%"O���բ
2+4��0 L��)7"O�M��nǻ<�J���#��t���;"OVq�^/f��+�F(|�8u�R"O�hԎ��m�%��ǚ�]�
|�"O�I�GT�'��d1s& �a$���"On=h�J�R (B$L�}EB�S�"O�	�2�1Cb!x��A�[��ت�"O�pQ�D�w������ۿ^cr���"O�8�a�#e<V@�ƈ�N�����"O��Q���O(�M;`�0m���"OX�Y'��"�d ���;g�t��"OV0K�,�#bt�"�l��"O թr̂
:��g�B<V�!�"O|�I�c
'9_Bh���ٕf<&$�"O:1�SI,�2@Sȗ�%;08�"O"�W"� :�; �iTp)�c"O(��b�:�i��ZbH�{�"O��M�6z���n�V4x�"O�(�a�s�P��&t�R���"O�1�`��5" (u�e&��}޺��"O��Ac��6z&*v�D�_� d8�"O@mj�Yg�|��oԅb�<�"OR`���� �f%�uAQ�Y)�i*g"O���U�[/����@P,3�A�!"Oqz� �+F��HP��$Gl���"O4-a�葇<���	���;&  ��N�FɞyɁ-�H��b(<Oй� ��/BR�ɲ�cO�J��3"O Mi�Lܵ:��`�hD�.�.��F"O���(�!&)2�FƏ!�1�"O�T���A�WFp��&�$$, X�"O�@��K��u�B���䓭7�Hy�"O�|�R_����xピ�1x�pb�"Ot���H>���e��"��d�!"O��@D �!=�̩2��oA�qY�"O@����+z0�� ��3?ذ$�"OJ���C�5�6�'	��\�& ��"Of�uΚ�0���Z$��2��"O�!���P�a3p�s��$�r8��"O�4x�`]�3�bP �dh��e��*�Py򦔿@$�͚w��~&< ����Q�<A�	ˌW�9�ŸF�؃�@Q�<�`��S�:����,*�BdKS�<!�G�:r�!�4�� ���K�<�E�ڽ;M�T*T`�u�:����H]�<��#400�GL�w��2��]�<��R+k����BՅ ��%@W�<�a��=���⇏�j+�I��U�<�D�U����5�� ��×`�Q�<�7�43Bd�1}D)�'�Sd�<��@�:K�"h�#����A�A�L�<�B�۲,�nM;�A�V���wE]�<!qĕ�q��Gl����ҠGY�<�PlX���ۣn��	�a dl�<y�K�%�ʭ��J&Z� ��F��j�<� ����o�R��ܭD��	3"O��#�c�8Ӱ\9�g� �>���"O�M%*�80̚3'�����2�"O�@�IC1]�R�3�e	 `Sn�"O�� X2�N56�~8`�p"O��a)R
���1Z�"ONU9$M�5��pyA!�.0z4��p"O�,�3#�8<f�H��]$zg, �"Or�`��*E;��"W�!Ih��"Od��7�0"g��g��>� ��S"O���G�X�mj��իN�}�Jq	�"O0-j@�Ǩ�"P�J�$T�L)$"O�P2FᕅD��e/�U
��"O����ELP%qt��5�8
�"OK߱:j��ʤ�A;gd�k����y҉�=L��ThPb`|� 2nO*�yb�x��� b�V}���K�y�k�
L�� ����.F�ȰJ`/��y�C�)E���3`"��?�V�B ɓ��y�*]�&<�"��_�:����6$�,�y�oݙ.���KIE��bű��ٜ�yB�.=�2�R�Ǖ׌��^�y��� [\܍C�T{��D���̜�y���Gގ��Cc
2pk�xCՌ�y���H�p���5�8����W,�yț��< ���&VH,1'�I��y�k;8Ү�� �9
�tx��V/�yr�����1�G+������N���y+G�j�@(�A�DЕ�0�y���(8�V�@�d&v"<cM���yrc]"pU�=sT�%�6.=�y��Y����$q�	CѠ3�yR�T(Os<1�����1�ĸ�S&L��y����~!�]2cΙ$���#��y��D'CEh�c$	��tp�.�y"���vh~�I�'��t����jܹ�y�ɨk�~`S��H nG�A���T�y"aQ#6µ���==e.~�X��ȓFl`�Q��\�@a��M��蚀�ȓHbJ�1lTt�<�K�������&��WUƬsn���0��6����$q��|�C%�3 R�X�� �Ȱq��0�d���E/&�(���yt!
�+��X�Ƽ�(�?7L܄ȓXr��)C$�=(� *�E�>B-@}�ȓ5�Ec��բ��WN�F�"���S��8E��V� A�`O�CQ�Ćȓ��M�W��z���ӊ(-��}�ȓQ�*�ʤlM &3�IJ�)�${��Y��V���pw��/L�s�� ����ȓU��ۓN1a��Tp+ˈQ-�B�	�eԂ|Y�ƄtO<5��O�/&�XB�I�/�53���EV�Ѧ,��m'0B�	�}���#�	�����`U_�$B��9R3H���;}4Ҍ�OӍX��B�	�| ����f_&H������2z�B�	�Oon7m�u&�����M8_��f�$�Q$(�<&�B�z-ղ��'1D����Qz&|uHb�X�w�����.D���w�����������P�L?D�0%脬k� Y���1�(�bԠ0D�H�##Xj�J��h�"A2�0D����!�g�2p
FH����!o.D�� NZ�2��!��v
�Y��'(D�� p���O�p�,:'�M1�r��p"OnLb�&�Y�.5��'�)v��L:�"O�Ȋ2mN��y #��&�(i�&"O�T�t�%���đ�y�BE "Olmb��b�����٧@����"O��ƨ��0�̑�փGihV��"O���$�K^�8 �%�"-T\@3T"O���C(#�F�@�OG8E;ĉ�D"O��7��-h��b���<q�V���"Ol��q��kZ�` -/|���T�	p�O����l �	ƌ]*3��1�'����0a�}I�fM��bx��O��=E�$ �FԨHS��Ѽd�`���y�g3s~Xh�p-�*U�|�Y��T��ym[=�1k�A��T����@��yb�n�4�'OP��P[��*�yҧۍK��hq�B�K�ԴC�It!�d�2'�v�1D�a���@֨��5i!��\�1��0	����:��$i�2A�!��:\�Y���b�� �q�!��'ox����/1��K'���Gt!��^.a�\c�ǋ�c7�E�P_|!���0��@�,j0e�E)@�od!���7��p�-rd �ERq�!��O�X9��Kb�E�G��˶F�7�!���.�ޘ�Q/�]pЉ%��3�!���/�(��d��->�`�J�6m!�d��V������6�:�x�$R�zH!���(Aa��S)h����)5!�]�=y°�J_$^�2YX�M�"~!�ڥ
ܨ@X�a/@z����mʟ+l!�D��Me2��76loNȑ�LJ�!�dC�D�TQ�� {���ꆬ?�!��V�	�1 wM�?b�^���iI��!򤀔�����A9>��<i�K/we!�B���H�a(�L�<�R�ˈ76U!��O��17��-��@4���!�$�9h��AV"� )�a�E��Fn!��ȼZ�K!b�;��I��$U!��O
$�S�B�$^	pW捪a7!���o�����G�4�<�цk>l!��6`VfY�c	ܶD�0L�t�ҹs�!�$�w�4���.ÔZ�X!�`�Iq�!���3ɞ��6D]�)���;�
΅J�!�5q�RP�4�Ĉ$����&kL5{!���7;o$i:�Ҋz�x��iM#i!�ĉ�y��Pv��F�l3��M!���X|*)�Pa��ՈIkU.�!��<|�5� #�s����'N0<!�߾P������*bV��[�P!�D�(�¼�WF��]J�I�Ǖ�!��"�J�*�A4 @�u���I�r"!��X�
݂���>����Ċ�|!�$��6TT��_0g������!�[�s8x����{$2�&�G�[!�˼�2X[' ƖAgb4
4˅C�!�dʲ`��MK���9Q���j/�!�D�-�N�c ͚�K5�i��G1�!�ه��=���H�xpm@H��g�!�s�����*mH��7'�"B�!�d�5hp�!f��*/C �ۣH�u�!��k�F�J���_��6gH�lu!�DU�8���aK�{�h��GFN�N�!�T0u��hU���R��m�GǢD�!�� �tb#
�*&�� �J�+{��#�"O��'$��`"���?�Ƭ��"Oɠ+�=uz<��a�3M�� ��"O�<�&8L�8D3e���r��ɛ�"O��tMn�A�х�ky��!"OhI�D� ʆD	��ؚ�F
A"O�d�t�إ
��H��搉��"O��n���o?|l(��Q��^��A"OZ��6�L�\��D��DS%�M"O�p�lC,}�t,��X4y��qA�"OK�9m� �!CEH�-����A-�yr*RFִ��CO
%�&�����y�C�.�%�F����[U�D9�yR%�Q�v�ycd�~�q�eԉ�y�II�xޡ��*�P��sG�ݡ�y2$�YԌ�s��AAv�9$��%�y�@�`,=�� ��7&�Ie��y�iK)a��p�Eΐ[ USKZ�yr�͊"�����,·�PiID�	!�yb뀥s5�`�`��I�>�R��J��y�lŦ'��x#@�.]������yb�$�d��RC�,t$Q���y��?�hX�O�m�&t�+�&�y@"A�5��Tfbd1�&�y)�L^�F�SE��%c��yrL��()����b,r~y����7�y¢�f+t��&��0u�p��$��yB�r�f��Gb�}5b`����y�n�;(���;hH��`�α�y�p�&�
�" Q�Cӧ5s&M��'[���cH(����p�
b�*���'���b6�%e0���R�Z�I�'nT��E��Z��:��Y�L���x�'{P,[w��D�^1z�OP>B����'�Ѡv�O�5;�a��B_1��x�'��h���y���e���'�}���ʯyb��P�+҅� �'	�y���\9�������5SƐ8�'L:@:�١v�I[D�Q3i���'7(9������BV�'`��	�';�qSu�-�n�7a�����'<�n�	 ��0)�V�$�v��'�����Φ��C�ۊC�8��'�Z ZD�ߖp$eyS��A#���'&���L˓#�z�BP&�6"�R٨�'��+���]̊x���ĴP �'<�M��NǮIZ<�Hr/S�!|���'�x8 �68�.�B���!B���'E�a�K��mv��"%͈PlI��'c	:��A�C�I��~�@��'����P5�e������	�'!��K #ӌfDҽ��K�8$�@���'��5K���$>�t��A��Q��'�N�Pbɋ<�ܭ��cG��8�j�'
�B�+�Rힸ+�>�� �'��q�F�ũ\�>��@���
^.�i�'� %��Δ��x4k ���9t�"�'�(�,��j�!ӧ��z�aj�'aXY���G3P���l��y�6�"�'��Xb�c	00��j�ճt|Z���'g�R�!�+1\\��"Ӊh�ʡb�'�H�v�Ǣm�2�����d~��'�A�
�	t0���V�ԛ�'=��B�E�:@`�o��AC�Z	��� ���U���Xޖ����C#�b�Jq"O
�1��:$��v�U)d�����"Ob��ѭ¦1�FUG��m��c�"O�����\1
9�I�+������&"Ot�s!в��m��KK3�����"O`B,T01y �)5�V��|L��"O*�8R.N�0��=hER��4�A"O�1��ب*�	@'������"O�!`��0�A�O�(|���D"O���w�ӆS���H�1�|tzA"O�i2�G�.��A)��O(�����"O��@)D)nxnI�(�1��mIG"O�؆c)B�<�y�<��%�"O�� �٢u�h aS��I�� ��"Ol1�1�V��^�s���$7�<D�<�`LQ�B�*����(]�H��G�9D��XD)�4E[0��5�|f0}��:D��HҏUt�f���iM�=aJ�9D�H�r+P1<��h���	�U��"1�8D����������"3�ڵ���7D� *���1�t��"`�h��Hbu�5D�Ra��+!�T �T!)� ���3D�0�M�NwbE�+X�1�F�Y�=D�����H�D����Tn���i�Fo;D�,(4n��A.`!6�4�=��4D�h�5kY�ٜ=p���~�R}�U�5D�P�WOՕW=���J�(�l��S)D�`���A�p02���(j%0mPe�)D�\��'�0���aխs8���3D�(t,XWL&H����Yp.x1c`0D�$�[N5I4䊏�R�0SM$D��F���D�"���+��o�:aX"N6D�L[5�	�<��J��#T��&�3D��e��=��\v�-=SR=0cA/D����K�y��D��Y��*�X' .D��s�#ߗ�<� �F��N 2�-D�8�DK>8��@P(1f�@��.D���h�)��	����mh`�!D�HP�I/_��Q��� �9�.�*U:D�pyQ"�&��*��
�@��I�,D���D	R�J��� �ITe ����*D��`��M¤<xH�Ѣ��%D�|����,=����%Z0xt�#D����.�.~[6�8`��w#t�Z�<D���*^t����d��Q�d	��k:D���F��+��ar�
H�F��`A7D����B�>J4���J8Z�,�Q��9D�h0t��S���kq��6Y�׈5�O�i�P�hL	W��& (��LA�&U��2|�eS'��d���
��	��D~r�S�>�܁{�m΁dxj	3B�o�B��sj�5XQ�ʕB�P�Y��Że��B�ɱ��W��6�B�io��_T�B�ɍ9��� ߿`:���A }$B䉦_�@��MK�d�e(�cAf�B�	2(��������Lm���e`�-��C�INx{�&�j��[��]?O��C�h��t8'��~��6�O�A���ȓ}���� ��P("��
T`���9��y���P?]��H{2�/+W��ȓ!�H`��;Z���4�\�%���ȓg��iI�LϻDђ�d��sV��� (�����Y�H����W�2S����?���
�$R��MҠN�d@��S�? ��%ˌ�G5H �7�5��"O0h �āpm6HA�L�{�p�3�"O-�%�T���jr�(,�09C�"Or����6:�y8��0�n�"O���Ǒb.(1�U�S���t"O�r6ŀ�d���`��F�y��"O���F��J�m����.v ��H�"O`��qLD/j�,Y+��&P�<-�S"O�Բ�(aL�*��ȩ.ɂ$��"O�EʇE\�i?�` �
�v5��"O�|0�M]�N��ekъ�3*�,pq"O�c�[[,Ircʒ�'�fYb�"O ���E�+cB�Չ1J�;�8	�"OL!�n��b*ђ�  򨙷"O(|�sIř=�@1Q3͜<�$�{0"O�x@�ȞbT���T�kU#�"O��v��xF�0�	�|bɰ�"OPA+��K�� �ŎE37��r"O�a%$��^ή��$n[Y�̨e"O�L+!I�Qe\9�`	5�R"O
��S�P�� Ԯ̓=�QB�"O,�&�66�z��W�YD�=a�"O�X� /D�
�4�35��(���"O���J\�#�D��������"O��Bqo��t��=yы0sε��"O��r$�H&-x4-��ŉ4�0t�U�'���7b�aP�\�x�PB �DB�I�2��D�BY�R�Tt��b�&�&�=�#fAt�O����Ek4�T�@�A7����'��ᓢ�D`hEkqgÅ4��Z�'X>�Ey���C_5hܑ�)S,N�� !�K�F�!�DB���A���P��(�����O���y�(+!#T�(��B�G�&$�d��ɍo�v�*C0)�q��"אDYd�+'�fC�IF]V���r�n�)��K1e,T�>�W�ӍY���
T�=B��@4f��5��C䉕4B1�Ī����+�N8��I�!Q�#<E��@�cS�LM-�����y�bW�ðhQw����4���ɶ6Na|B��=/��@�݄p�.�#��p?�"`�x�����YyR�8���C��PP+-D� `�#��Ȩp� ��y��f�)D�w���w����B�W��r�)(D�ڥb��<Z�H���V)h��D,D�X��њS���KՎW�J��\��(D�[��@1E��XG��ü�p��$D��iH�kY�(P�/�3ע��An$D���VaVYD|��C����*'D��f�Wx�l	�	4a/�Q���?D�Q1��A6�G�:(p�!�`�=D�h�"l�J�H)��R�M��M�wK/D��Q�@�-�ftB�,�_R|��r[!�d�z��80��&
��˞�e�!�d�	#��ecɶS���I��!�Ĝ�#*aK�N��/�6(En\�$�!��Q-��R�JI�@G��LI,�!��^�a`�8z����BrU��jLG�!�D�2`�����7`��U�G�!�FTؒ6 ލ ���錄M:C�?~^�x�!X���h�lȽY�pB�	\�f�z0�ۼkϜ�a�a�9/xB�Ɉ �x�A����Dihh�N}�dB�	�:p�hA&l�'7<zp�@�j�@B�1���x��I�>D�p/@�9��C�)� ���+�/�0�	�n��p�p|�"OH`�C��\\��1N��*�&��"O�2� ��2���rnM�d�Ɲ�"OR5��!H7[X�e�K�R�Q�B"O�hE�M�W�jl����C h�a"ON	���50�i���#���"O�ɩ�k�����H� k ��"O:eq�m^3@���q�	O�}�~��!"OpMi���?<��Iqu*_�wʐM�e"O�9�E�9ڬ�i��[&
(� �4"OX���/?`��!���~r��"O�kV�W}���C��2`Z�"O~,��1oR��Я	&Tш"O`QJ'�ľ`5������_���7"O����ߔ�Q��/��AӾ�S�"Oȥ�j�N��	3���\���"O8Qb.�&/���#OH7�8��"Oҵ�@�����*%Z�Hǆ�!��"�4���))>���7��!+�!�Ğ>|\�r��&�E�4�C�/x!�!��2w��h���Xօ�n!�DL+lj��H�,�T\i���A!�d��f���b��Of�(s�Д!�!�D[�e̴�[AO	0�Bc��$�!�����PQ��Y��ջ�BM�`�!�$�l� Hx�K�T`f�� ל3I!�S3���s��-'Fຐ@I6Td!�D�&o�y�*�}����P*v=!��-��T�rg�P&0��t��!��3�Ҩ9C2�ѣ��e!��6(�~Ĺ��ƒg�!Y�`�3}]!�S��S��0uXh�� (q!�$�+7Ĥ[qdW�{�(3# � 
!�]�ȴ�;��ۙ��8��ۥgF��D1xx��R��A
��A!E
�y2
x�X"����~p{�h@=�y�L�%���q�1�29p�@���yBF��[8(����Ւz�2`��	:�y��ɄY��j�\�xS���@���y��Q�1ômI`@j��1���yRL��u�(M
vh�1
+��q����y��Z g���R.�3W��c�)_��y���y��Q��οHC��C%(X��y�ȓ�o` �1ʃ>@�@�j�	OY���>n� �oj}��9O�E��!ʾ �@Ct�{f�%�{`\"�ͩp����v����N�Gh�9�O���;�N@'���e��i�gG��ұm9;��${rꑤ�4H�3�  8�!S�.6����1�~��1�� Rn�e+�-Q�#���nD.����i�+O�$�s���`׍�;�sãǉ#>~ث��O��8���'�l�dC� ���J(���	�������ٴ�䓣JZw��<*�N��,�v�봧¿)Z�\s�*�<���È����'��x���ĢV$@�Ґ��ZFν��l@�:요r� 7<��&✳
�����2`Q�ts��|�,0��a��抮X�`��e)�_��@��,�yl�*��T��A���6�Q`�Z�lq�(�/O�m��@��8���:G�,�Y�X �!�O�(n�HO��TiD���	֊`���ǁ�zj֍�O\�=�}��,a�� �AP�#vHG%oڨ�nڽ�Ms��[����O��S&.�%�1�&x�������J�0VW ��	�<��՟��歁۟���˟��|��t-�xl>0����Z��E9f��Yc$��I�t�p+`�O�J4���� Pb����n��P	S�8��HqÛr�'y�9���4 :d�3;y���nE\�|��� �xN�v�'����4�?�O�$��D������D�I���b�'kaR�W�U�D�B!�	�S"tA�T�P}GI��7��<��@�!��.�O(��~�ѯF�|���\� ��)z�J�$
�'���'.D�2�\�a`z�ے���ȁӐ��-e��SE��6�L��b(�2YkF�(SB��(O ՘E��&��9�1n�,Y<P T['�Q����:\p�a
�![�O,ڹaʐ�(O�Y��'��7������m�� J=ۦۨGx�L)@ ϰp]b=S����8�?ͧ�HO�, DbK����`n�N>����'_6��Ħ1l�*�B̓J�Axm�`��$���I�.\���k�������	oӼOƑy�\&~�>�4��	|X��%f\6
��M#t�����f��\j �v�<��O���;R����BE\Ji�c'j_�wZxmm�:tX��.I�D��m�H�2�2��S�G!+�ҨY��~��@kʐ{��C��h��C�ݸ�l�sO��$Ӧai+O�D�s�`s�C�4 ��E!�ᐂV)�%�Q� ꟔��Yy��'��O�Lv.${6�� h�e�F
E�Dy2�m�bPl�����ٴ�?����uG���1���:���Gnf9!�^�f$6���Ov(��&HU��D�O`�d�OZ�;�?�ݴ0|:T�ji�l#Q.Y�%TJ��O=y�Q�Ƨ��Xi@�X�~�Dɕ�](�+K>yV�F8R�fA��� ��ȥ�ۮgֺ R�I�Y�-"RƇ�h�bq�O��L{�J��6/Ѐ���P��ju!/5{�lS�`���󛦩[�,O<��>A����;B��n�IHe�"CZ�<q��\4V> �Ҩ<^h��y �+��7�S¦�'���O?���䉏  �����)9x����W�<���';�fF�1p�i��W�<Q�N]�S\����f�xej&�V�<A��L�.�<IȦ�P������g�<	І�A�erN���q���m�<�f^�֚tz�KZ�0er�T!i�<�f'Y�)�%sۭ:~AƯ�]�<y��2�J���旨q�t1�.Au�<��($��Kء,�������W�<�sG߈&`���	�uZ�;wd�P�<�FiF�HuB��]�$�w�`�<!�N��$kj�a���g�Y�ծYX�<1K�o��`	wׇ
*���P�<�q$	!���8�ˁ|T�e�RN�<yv�Ǧ	������2?���q�t�<�bX�=�0��@�-���`l�<�E�ϯO5P-�U�U�Q�H`Ӓc�g�<񦄗�Sw��Fa�%},ði�~�<	Sn��\/,%�W w�]�4�o�<a�"4'�"��C�2m�*yjc�No�<a�]�{��@�F��. $<
��Pg�<�w/�%�d�d�G�m����'�d�<�g�_�%b�8�"�>��4p�!Xe�<��"Ļ@��A��f��lӦ�H�<9D���e���3c;�:�C���X�<��@���x�V�_?����gM}�<���p�"� �<)��@����x�<�3�H#	g
s���tP �NO�<YF�߰ae>��U���g�C�ɢ�& �rk��m���5M¤^"�B�	�E�L���ƈ �`��ߨW	�B�	�8��b%`=����h�C�I��f9F����4���8�B�	'�D+'ڇC�����gN�:m�C�	�:�,���S#N�v��V�=7P�C�)�  �� �4 ^DV��:P1l�""O�\rՀ]�:�!�	�2.HH��"O�	�
�<%KB-eiP-&��	q"O�p�!�ݽv�L��L�V]�%�"Oz͘�,X�7���ـg�
hS�)��"O
(�vAW�h���&�)'��R"O��a�PƍZ��.C��*�"O��kY�K��hهJ\7X��y�"O^�:���&>�X��D�V��"O$}+s�R�i��Yc[�h�8v+���yˮ;��H٤oK�O�-�r���y2�)�p�$C��9��� 5�G.�y����f5�"F���d�j��y��?4��D������C���yrǎ��HR�g��
p�B�y���9Q��+*zX��tL��y2�	_��P"���(�4@d����y���=YFY�
�1$2j�c��V��y��<)�E�7�Q�!y"�K`%��y��3I5�����"x���y�i^�m_��!�AÝ]�bxõ����y"LϻH腀3��Ok�I����y��	@�,8�"�LgR����y�CU�J�dcIXSV�������yA��}�N�A`�J�;�ȥ-��y"���A\T�FP52*� )A�I=�yr�O$Z�c�-�����y'N>#2a��G�G�M�I�yR/f�R�zU�W�ɦl1pf���ybb�".�Z�I��Q6	}�@�F�P�y2'��`��DKԄʉ|���Ԭ��yb.��~�tZ�i��)��y���(�yR��/L�^Qz�ѝ��� ."�y�J�3G#�]*w#R�
&:d*�I�yb��)��t�cG�'
�x�ҊD&�yBm�a�q�4a��x�<��(�yҫ*��j*Ϣa�N�ᖬ��y���k��%p�LL	��C���y�OX}���#��Ͱ }�9�un���y�g_��0���/Q�yѷ+��yb%��5�]p�A�,E���f&	�y����C8��A*�?,s�y��B��y2��7%J�1��A�U���@�yR+��@*r�rAf��R�~X�5��yr����aˆ0I
RB���yB�I?1򌼻�M�#A��AZq`��y�"�&i ��D��(��x7$���y$t7̩'̅z�v5P����y"�[m�� *�%.v����T$A��y�o'��4XXʆI��iw�<��P���S��|D|��"Ź��y��Wr$Ę�T�+Z�LyN��B�ɿ�� .�=��p�3$�, }�B�ɖGe>h���ՠ^"N�!�+�wR�B�	 ض=0�W����"�W�x��C�� �؝���� ��M��jbC�*P���+�Kɻ��Y)S	��p��C�	)jY��`��f�ò��	|��ȓ4R|xH�T8d�@�� ��5��
����E�D{huɐ�>R�\l��hs�ū�h�	
�;FNR AY���ȓ5<=H��S, ��&Ç8��ф�9\��[��5x���U6,�v��ȓ|�L��lW�1bL����H��S�? ��6�ET ��F�Q��� �"O8ȑG�W<X{&`��k]zǔ1"OM�'�;bh�A��G���D"O@��'��N.tdjf(N�*�t�w"Ov`(�nN�P^j�Ѥ&<��t"O�*WW�Q� �����0"O�)�A�bb��z ��,`���"O��s�C��:&��J%�B%URr�S"O(h"�m� ���H!F܀|Iux�"Ox�H�hƛ^�����
�"0J�R3"O��0T
ї\p��jf<�2"OXT�2oP�[��a�V�Z �R"O�-���c��P�o�Y�m�"Od���
�I�X�hK�u��,�3"O�H�ĞB�i�0f��
=9�"O�i�c��w&r�х�H�]��`p"OnMB�!\4�<��SJ�,k���H�"O~�)�J܏4� �cp�����"Oj�4��"(2��1Tg�>6��+e"O���2:*갛�%ŷ1�* �"OP!!#�\�G,,��VCC?$���"O6�+)�̑�5�U�Vx�"T"O�\*P�҉yBPa����< ܸ`s"O ��5E@��T˂�����M@"O��)G���t�O�kg�Ö�y�(�Z�<� ��L�l$�a��M��y��ݞ4�REJ��.s�e��l�y��\��B�y��: a$�f��)�y��!z�0�������h��yBl�k���A`垄O�|<b�* �y��y%��K0NP�Go�6� 6�!��Z������K��o�<́�׹x�!��V�Kv��A�
�<K��� O6�!���x�s1K�1j��qO�M!��*wP*���V�aP���K<!�D�itڱ��W�L����\�8C!���r�r	�7�D�踙��E�!�$��t�T���J�a�t+��U�r*!�%��]�OI�)pX��
G+&!��5_���S(�9�j4�bϞ�"!�ְ<�HC�"T���AΘ!�!��܌0â�t���"r�15m�r !��ENS�Ԡ�b�.m����K�C�!�$��h ��N��%e�0�`����!��6J\aQh�`H��bw�_�e�!�D�1Jh�Q�H�_d�-��&��	�!���Qh�5%�Wp.���ȳz�!�d^&͒eSuLU�n�Lqj���$L�!�d Ff�X�&�5�xڗ�]�>�!�䜬]�p�V�	�T#�a��E�!�D&EnNuӄ%�@�zݰ��=k!����¹#����%b�l�E�#pT!�d��~.FU��ȑ<Q(P�@U�y!�d��¡��l��ZQ6�@	 T*!��6p\�@�n
�wM�����@~!�DHqe�y����;Q���Ѐ_`{!��E��x\�B�O��U!��94u!�$D Ģx�*��e�r �2Rp!��TD�!8��T�DGn�3 �($<!�R,uz� � 0J���,�t�!�_�雳e��/PdI#L�na!��MeFv���g�&���#�O3]V!�߯-�`��`F�,�]��Y�*G!��׶v���IF��)[�٢
�z1!�� @I(�`�HĜIA��>!pi2�"O
}j�̟�Ȉ�P�-A�N��m�f"OdYs��� ��(Y�
-�:�IT"O�M%C�%�R�gB19�V��"O�aYB��6u�ਢpEX��"O��R�=���O��mH"�"O�)� m���pAS8����"O"�� fѽ�� � ����Y3"O�����Y�L�h-��	C&a�.E�u"ONxѓ,ۣ0����ĉ��W�^ ��"O^<�W�ǢOD�˕(Z��p���"O�����&ad�!�1�̇M���w"O�"P-��`۪���D٦=�pqA�"O00����/k1z�:F憪��00�"O�����HՌm1Ǥ�S�3�"O ]���Fx�D5FÁ+BHA�"OƤ#6L߳xn�1�2䊴:�D�Q"O� �R�"���C�
L�(�H6"O��Z`	�}6.���D�X�~	��"O��Ӡ�!zv�K�%߫=s�J�"Ot���T�=�w�iZ�e��"O !a�l�;z=�H�W �QM ��"O�BU%ͨ��ӄ��Q;Ɂ�"OP��e:DY�Չs�S�g$.]p�"ON�2��"|���o�5��"O�!&�׷m� ���4���{d"O��4��ai����4CmTe��"Ot �%��7R�$$+eɆ�O`��"O�d�%.z�Q��hK7����S"O|�2��Z�;C|�+�"�.�����"O���aJ�Vfm����-X^|8۵"O�`Cf�
+KZ ��ܚZD<��"O�X�R \
�U��HNxi	�"L�<�1���n��e[��݆���LJ�<�̞�@/��Q�W�&� D��aBL�<�a��7t��85�H
I�yj�f��<A�鋅?�z9;u��&�^)��DR�<��G��g% �¦�]��S�L�<i %�	C�|�b�ϊ�38j�TC�<1g>QЕO�w��i��&�B�<��1z�P��6�^!bt5{D�~�<����'\்́�m��H�O|�<1�+	�If-��*W�V?��8,��<���[ʊ0Ca��[@A ���{�<��)�z���C@����!87k�P�<$ ��0��H�Hl���mBh�<� ^2KX�ܸ��ΐf< �zp�R|�<��ꎟp�Ԁ�*_"/�e��C�<Yg솑]Dɠ�Ɖ)�8�H�D�C�<�"&[1B��kDq���OA�<1�K�.��<@1J�}"�3Mb�<)�e�6�����$գȝ���G�<�C�))�N�*$�"!}d�Y�NB�-`Ƽ<Z��D�xҨ��sm�;}��C�I�J]z���H���}�T���C���*���!Ǐ�~u�b�L�!��B�I+��j��)��J	�s��C�	� y>�#��E).;�i�&h� R�C䉓6�R䉢ˈC"hDi1+�#R.vC䉇f֦qx����b�1d��<UhC䉹}���% A���H��&]P�B�	�/�z|���4D�|-IB� $7vB�;v�)ȃ�ƳK���⅁��VB�	T������^
ȼ����*B�)� \�[!#H0%�0�B %P
��HB�"OB��u�ίM�W* �➜�"OP��У����&'Ք|y��"O�:��˧4Uʉٵ$ƳB�� r"O����`2jE�����380���"O�!"$�ѤkY�� A���H�Qt"OV��$�8�����!�q�b���H��I9=�`�I��@8�Ө�g~�C�	�}��Ȧ��q�xڶ��7$�)�"O�Q"׈��v��K3Cٜ1I���s�'Q�,kc�E�8�:mbcF2p� S.*�O��G����N�1s��!ڱ̂�vÞ\'��D{��nφ$�<�'��+D���:w����Op�F��!�>,���K 7~�aG�$�yBJ��h�BI���
<~�чN��M���s�(�b$�M^8r,���(�I	�O���2HO'*SA�8|niXQO���x֑o��4q�K�f�*�1ЬY.�yr��<B��8�eU.]z&��w���y�IO.^-F����$��ӭ�N�R��H���U�D�|��]:c��;q$��ȓM�F�!DdڰQp��d�(&08�=i�NU�'~�_G�hc6�02�ʄ�u/�b�r��ēE�(����dDdt�C�����O|�'b0�)�3��!�2 �W0�ČZDO�H��y�7�ɡ-�y,�GG��� W�Q�6Xc�'�Rm�;D���p�6�QS$�%�M[�OR�J�����.b>7M�	]mfi	A
�>(W�M8�� , !�d��9^H�-^�M*��QA	.k�d̓}��c�hD~����Gdq�@)�)P����>�W ��*a�C$8�S�Ԗ�] �g���*�O��h��ڹe�d$z#���[P���	�}А=E�4�Ҋau��f�";�ųBj��y�P�p"�M0�J}��mӢR����:�D�Z>�*U�ݍ �����	$!�d�aḟ��I_�f�8�	�H���yֈ[O���k|}�C/}J?㞌�'�6=������&�ԡ��2,O��<yc ��z� h+r�L.>,��f�Jy��'.��8�KY�rxI��#C�>���I�b ߃��ᧂ$A�h���I��~R�)�'Tc(��i %C����� ʎGxR�i�Pn�D��
� ա1��`�C�H�f����d}2�Sx�H��$�y��U�D�I���U�Ad0?���T?m�Od0���O��dC3�U�)�p���'������W����K��	�MRp"/D��A񪘇�BH�eɨ��ya��+�d �S�R��XcT��l+�1��
g��D��)"�a"@ϑvSXp_<��(��R.D�Ytf�9��H�dK����ēC|`𷂖���-�G'��>ܸ�#œ>q�"�O��$�R�!H��G�#�r�)��Q��D�6Q���s���Yb^t��!��X�!�Č�V����͔L�l�Ї��+�Q�X����@���Ǘ=3r �vD�/q�PH�"OTH��m�=إ�BQ�j^�Պ�E�U����r"ћ1�L٩V(Ի]��2
���y ��`8	1���|2��9z��y�d,{K�L�#�W{2�sr#�(@��zk&��W\��I�)� �+�L�R#>Q���C1��	"E� ���+��F�2��O �=%>��JL�X��OH�9+<��wM%D�<	c(�4�@�Qp��+���$"#D�̸��Z����I���d3-HN"D�PhP��0:S����ְ#��H���>D�� ʥ�&Fz�
pjSKڥsʊ}:w"O��
�Z�d�y�)��w����V"O���%�Ho�,	��ݳB�����"O���ǔ;�~p�ǘ�'��MH�"O��BB�C�Hlvy)�e��o(� "O �+4a�	�����bO�",�� "O�ر�,G<A�d�' ��s���V�|f;�SܧE�v4�$l=�nQ�J��\���������k�Y�٠��j��>Y�ΟCX�85��b��+�*�2 ΅( #D��+���*7�r &��>:�LXa��HO?�	�{и�z�76h�S �N�`C��Tq6jT�� ��h�3�RC�	�4@x�@�>WЂ8)Pb�2P�����<找
�x|��#RIe�$���q��C�:ɾHᶏ�8��e,��Q��<1��T>	1�'�m|�u�dG�l}�F9D��
�ݕXT<񙀢�	�}��.�hO?�DE�p��ǫ�;F� ����A3*�!�d�RH�L�����Y�!�O,�+��(9�2��ElȜs����"O^��%���~��'Wo� �r"O�j� Sv~}��)=H��=!c"O dp�%֚3��T�uH�:1��\��"Of$�s��-�<��s*F5?���"O��"�oD:��	0��gLq��"O �����H��H�^#A��B&"OF�sG�-�ʰ�@WH��'_"�;�/�z�t8Cv��N�vP��'e�����H�,H���"�3JX����5�Z�(�R�	*����=�E��cV �0.[�|����������n���x@�.Mv��R�E7�Z݄ȓ�B���Ş->���D���	�j��5`A�0�y�6�҆$��G��9��	Y���%L��QnD0'��ex%̄"$�!�dR
�t�Pd���H��d��÷
���@F{��ܭ����jvn�*��ޓBM�� �"O�y���N�4��@z��K�R.���`�'�IC�͈Ol�8�H(%?Na�@��)|t��'\��I,9��١N(/���[&��b$���/�M�G-��[G<m
��3As�O��v����iZ�P��A!h�6�m��혶!��^����4'*-�QH%mʐk���*�8*�N�Lv
��#�<gf(5�t�;D��+����NE���b��8{*�@!Щ#D��p�j���*y�)�e�|Љ!D�X���*|�N�"ne ��C<D����j�?6��`��b�:�����8$�,����28���mn� [�Ƙ=�y!~�8�(�_�\.
�1%�÷�y�d��ލ���ͪLCx�dJ��y��ečᅣ����dsuF���y����&]����*E���d�!�y�Õ��BI��M-Y��Q"����yb���bj�CDЍ;��m`�ȩ�O����9%=1P�B4|�K�3.uF@K�'�0�����b��dI��$0&���'�H��Vkŀ[.�Lg��p�� ��'�45��Hڽe�X��5]�3� x�'p1�ޜw�z9�`�.�`�K�'�
�zo� ]�8����&��
�'Rr+CMQ�>��Z����[(����'����+��"8� ӊ�8Y�L�!��� *���Ƌ�9X��WDö}��U��"Oz�rq�Ȕi� �$戧`v�l��"O~a�D�8Y+.���%w
���"O�řŉ�	Tr��!7�M�IY��9"O����!M�Wl���l\�t^&�Q"O�i�d���g�H�A�3a�(�"O8A���W``�
�<Jtȹd"O:��
7Vh|��AG���t"O69�g��(�������ب�"O��Q�Z�1t��1Vo�1	�"O�e���1���P��BA"O���j�~�T5�T��?x�0�86"O�U 
�U�D� �/\!���3"O����
�o=�X���J��"OX�@O<
=�р���?�T@Q�"Ov� cM^�X�9��EZ-1"O���i��V�$\��)J/@�:%��"O�a�W ºF���BCK�D{"O�8����;����bG"��Щ�"O�D	�a�?L;	 �`\7!����"O��р�a�N��f��	Jv�"OF�el�
D����.8yS"O�SL� }�$� �"r1���E"O"TjvLR�B�L���@(td"OX�DL�
F5ps�Y
e����"O� ��'R
T�dڕ/A%rϺ5c�"O�4�����k�.�R6�Թ:��8��"O�l��� _� a3���~��!"O��3�ET+�T�t��lg�]c�"O~fD�1�V�(%��3��Z�U.!�D�wx�B���#����B��Y�!�S�y��(>��4�_sw!��R�~�~����U?V�
ˁd �?!�$S+w8���ؘ8���U�ӗW�!�O�a����K�4��� �aG;`�!�A5Vhm�q���~�D"Q�R?cc!���(�����RG�L\�%Ǚ	�!��.ľeC��o�����cy!򄉰j��@�b��o��P�Wd"`:!�d�Nv ��'J9�B��EdZ� -!�z5�$J�Y��Ag�%dI!��!|���k�#>2�H�F |�!�6Znd� L��!��) &��f�!�Bx �M�.3�*�2�Ok!�$Q�l�X0e��  ����Ư�YX!��)%�ءC����z����Ø�!�d�#x�ސ�t	� >PڥzsNP1[�!�I�^��裥�P�$?F��1�.�!�DZ :��.3X�!d!�!�D�n����Q�^�0�xG@�#,�!�Z�P�"�Hto��)�D��!�d��_�,�� �[�u��0B��P/m!�Ĕ���9�0AA�=�@��r�9u!�$ËptFX��+4g��#ì[�:!���h���h�J�:\�m�Ы
P !����̍z@�N'��Qb@ՠk	!��Ƿ��ԃ!�6fP
��w�!�$ݦPT�D�f)����X�����!�$��Yo�8၃�1�܁� _��!�D[^v�qV�� ��%C�w�!�$�,�ݙ��J�T"��2�LD�!��^-�5�F�͔b�N�0Ǯ�;wl!��l��E��F�3b�0`���M�$T!��(����VC��FE~����&w�!�� XiȢC߸k���r2�f�Nhp"O.R�*@�U0gB
P>�`�"O���W�D=Z�Cg�#;8FX��"OB��b��m@6DzEG[�T0t	k�"O4 C���eӴ��Q���P�"OPb eHn���
RM�;5'jp�$"OJH��,t�`t C,)��0"O�b�E[;]:�����_�U	�"O|IE
�`�zH�TJ��	���zp"O�t�+#��a��?ǰ03�"ODX��(ĵ@=bD�§\4��T�E�OL��D{�lq�D�f<y�G�D�!�n���ů@�(	&��e� �CO�藏�_����S�T4���,�d�O�ʓ
5�Bb[�C��]{�¨K(Hȣ�I�Mt!�D'����"1-2,10抎Ib��b���@a�f�!$��SAP�H���0��2LO�TZ������N�xh��D,LO*lxu�f�hm�� 82� {%Ov��Q�
���2�A",$��@Q�[]���C
\�)en
�tq@W���	~���O?T}Rs����q�L�}8��	�'�j����,^���Ƞ�ɥ
� Q�'f�!���t�d �)P�d��Q�')!@`gC�1)����(@�ON����&\6^�i'��1Ǧi���Z!\��m�ԡ }�O��h�O0P2�+\W�]@�L+|� �g"O��q)��Peq��M�\��z�]�hΓ�yR�>%>�"���&'εS�h��3�� [n�Gz��~'�ƸA��l��\Kt�P�"p�!�D��-<�Y#bo&i*������O�ў$��	C�����ӯxL@��Qb�WUC�I�1��	���-_�ph��(J����$0?��,
�d����ŋP�ґ��O�q��� *]`~���Y��a>7�DH�����O��~�wb� n|��mW�{&�4��Ro�<���"�ڼ�%�6����Qm�<!aM�
fr}2�J�aU�}q@�H)�?	���9O����&����u "��5"O\!Y�%_9EX����9X .=Ц"OԄ�C��_�-��"b�$i��'���8b�O�/�b��v��|5>��4�<a.Oƣ=��8�j�(ߊT@#-3C��14�'��䁊6J�VB6V1jh�t�G�>��|�ȓ@mv5P���Qd�l �n>\DR�d�4���lӉ\׮��7K.3�C�S�9�˙�@����
�r���$��"~:��H�q^ 0� F�F���G:�yb�J~d��W���Fh��M[��hO���I^M2Pq�&U=L:��^�B)!�ă
t������L*���/��@8!�$���}2#蛶e�0�2�M� 5qOB�����J'�)��a����׾
#!��<[�ᙴ�Ѯ2���$@Y N!�Č�m�0��b�Q� ���i� w�!�|�r�*�+�%o�LA���%��D�<�I�LF�/ӢB���˝�L�)w����y�#R�L1����mH�~V0�7� �yRK�'PĊ��@Ʌ=qⰹ@V�@��Px�듶z�h6�R��es *R�W\d�(!O�ЊǫG�_�N�@2�]�ZV�JG"OB A4�ǋ�$�ʱ�E�X��"Ob�hCLU?��z�˸��A��V���� �@ xp�*N�V���@I�6�!�� <M2!��Q0Bp�A��ZukS"O8!�%��Q�sc�~q�t��"O�i�� �P���zARuVi��"Obab�g��т�A�~��!���-\O�Ԉ���.�(���)\wА�1"O�]��݊i8A' ��Z
�[��|�O���C�A�(���� 9tځҵ[�g�!��Lo�(2��@�a;�������Z��B��(����Ų���)f�� >3X5K��'{�D�B��@�]$Yz�����	�'��!��Îf8
I�����21f���'���:N^�(A�)�%�?0�$4#
�'�P�S�NX�Fm����*i���#�	�����'p�s�����T��> t��'��,�R��|��@�$dB�hn	�
�'j������=6���a,N�8�2��H�ә{��ܱ� $Zv̳T��(^���I�'�x�ScK�/uF��q�Ās��\(�'gl�@6�Ծ!}�� ]#	j���'�dZ5�I{|�8%l���:|H)O�ʓ�0=��A ���](r>�-��C�H�<�Q��r��X�G(���"E�!�Č�=���A�L��.�2%��^�[!�ę+z���X�@T�%qrDx���o!�@�xߺq�a�,�����-
,8f!���R[nA�C�~��{g-҅z�!�DˀBn4���=(�>d;��FM�Q��	�����	�`}��d�؇ⰍP&�W�!�$��]j��AG�=�Ȅ3����=a!���q-b�G��OϚL���D[;a}�>��`ʠ.'JY2E�S�P����K�<A6�%k�-;��])!��M+�Ǎ_�<��S �3,I��E�5@JC�<qpցR�>%�墕�:�P�
���x���hO���A���W?�l��ͥE1� �ȓ |�ԣ�(ιgԘ��D�ĺg_�H�'��ч�I7L�~��«�VP�Qjc��T�Z���n����V� ;����*V&L�A����q�'�������p�Xŭۃ6�s���<�'~c|�KTBn��ɔ�=#o�4�ȓ��T""\�gm�%�S����'��F{��D�|s<I�d*Y8O�|=(�����y�(�4'�� \����V���򤅃��>�`	��n�~��jόW�@�C�ĆU����D�HŲ�>V�@T ��÷uJP��ȓ:�n�P�ǱK����Dԯ!���$���'i�?��Uk��$j�ܹI�;I�8�1�$D�ت��A{\b�u��0O?B"F)�O�B�IE��W-��D@2hT<(�*"?q����;g�pI��h�����"�Ǎ�d��81�$N�6&��#��}` 1K%LO~�����
�R5��B�i�
��פ�����'ha|2制eD���#��u`��&��x�ɑ����2z����^��X	�'�V�87��)X("� ��� Q���2�����'��'���	�a���c�I�9o������)D�8��Q�A�`Z�ŋ�_���Pg�2D���@�
%:Ԡ$�@��k�x���b-D�ظ�AV�ZP��Be�7JI�㇦(��p<Ia��%�� ���^kv��O?qL��G{♟d�!>����5�^�A�l����%D�T���g9�0$�Ɋ?�>u���#D�4���9*,T����?��Zj6D�l�kG�xY<��bÎ�g$1���O����S�O;�  Ԫr%� ��xH�k!)��Z$"OЈ��	�+� ��0a��0��v"O��r6��H�m�"A� h�M��"O�����3U&°h`�ÕxR��A#"O����4Fi3�N4l��ڇ"O�0���w6x�t��)0-��"O(`wE) MHq%�H�gv.���"O*=q3���H�Z�ˡ�[?P<0=h�"OB}�bN�Y�a���8&-�`k "O��@e*H�x���!�G�uN�q�"O Ao�5��1�p��0i��S"O����U>8�~\rB�U�z��T�"O���QeP"O�쁣/M�A���t"Oh4;"aD�U��uA��Y4^f(���"O��R
z4�8r�`�F6l�c�"OvL a��u�7�Y+/=&<!�"O�����85����jL*ލa%"O�p��R:W�d�s�K�|f�)a�"O]�b��܄86���D�j� w"OzPs�nH�]�怢!���_Y�Mb�"O|%�D�ܠ2��%01ˑ-uW:�[U"OZ$�W������쎂AI�y�4"O0��!m�r�:�"T��N0� ��"O&����U�ȅX��h+rq��"O�9�F�/|��3D��i*B��c"O�ei��κs���,�����C"O�, 2�I�_����`֑W(�9�"O�!�G�R�nԩ��)<H �P�"O�q���NZ��ݩ?����r"OHEZ���sZ��V�`��"OX�)Dnݍ <U@���8�L,��"O��Z���
[V����>A��|S�"Od���:2@h1�G��t:�"O��J�%B0O�E8 $[�`}*�T"OH���l׼ZRH��a_�%��&�''��XufO���� �hM�d���ʢ(��"���	C�"�Ta�r��/�ɇȓS��<z��[*h� h�"K<�ąȓ,P���@�fžՃcE������ȓx� ��#�gtP�Pg�?J�Ն�%�(a4D�3�l��宖:[}���ȓTw����,d"ܩb��#pQ̆ȓl����."&�� ���#ƴ��ȓI>���b]�8�L�h4f�oM�܄ȓ/_P�MM�h������+��)�ȓ*cV� ���/~9�a��X=���ȓn�l�8�F�Wm2��C(0���ȓq�����%�Y)�DF�D����w�p��M�Q/ܙ*�'ţuZ���ȓ*8\�qT���Q�f�X� Ҝ�ȓeZ"=��E�q�N�X�IO�{�Ąȓ�,�����DYvT��;O�¤���Y�nP1`8���J,?���ȓBpru�A�f<��9�S�I'�$�ȓĽ�ɀ �� -!�g��2\���6嶈����Nm(� �7Op*�ȓ7�`j�N
����ԡ��ds���ȓ.84�$ث8F��s�G("��0�ȓ'��jK>� �8cN�)�����(1� ��&���Ȕ$Y=u�ȓu�F�0���(B����Y>s�Z��uj��ޫ�����K��]5����{��=��_�5I:,��hؖy��,�ȓS`�u2v*��u*���C�H�N��S�? ��'ˈ�'����'ّj7p8���i�f��$Px�taaʕ�>/�e�7��n�R�s��:LO0��pg�7l*�1��'����"��g��X2�'R\L��'����(gX�p6+�&,x� ��d(��Yp0m��@ĠCy4{pa�sy�EO��9�O(�a��7�P��)�;1�.�ɍ�D��v�ִ���B�NIށ�G���ڀ<�cB!!�e��k�n�H'ĉ="N00Rܦ�~bk�:#K��)B�P��x���2g�H�q"�ȌI>�d�½�~RJLc@l h�	�����@��e�B�Yr�J>�	D���?%kf�U@.��bG�Lޒ�r� �ViAdb_�:,z�����.�F{"�<TY��$��!��|��(���hD	p�O
Msf8 R(O��!X��F�����Ƃ!��l�P�P��txXw(6͡���)��S�ow����(Ր�,����X�������o�#UG��@���8��%GO& z����E؋Q��PL�Yw�pR'�{]��8����>��5'Ϧ&v���GEىU�Ι�pL"@
l���	1$&���)��GY�牶}��4 3�B/�z�h���"BL�g���5,(��ɗCS�	J��!J���G��;���R�U�W0��a܍z��`��� �+�^%K�e��N���g�M�:���bo��]�d�f�T@qQʑ�q�8�
��`v>x6*E�
�c�`�S�<��G�c�Bh)���8w�`5JS.au<@v*E�;�̱)��]�$T1�G��:TX��h��.���BGq4����E���'p0����dQ T���o�vɲ0�J/8�N�Q�.��4(�d�6�V���ܪ�7�.-�"�&o�pݒpK�9�B�a�N�5%�P����e���)��6��t����.�X�h����.�R�(�MA�7���+CK�+ ���a������8E����&˫�̠J�@{݊6�H4vZ�tY�b��Tkn5���ړw�Lk���P#���W�$=r�AN�X���Ф�?H0vl2��'�@���
�	@��ӄ���RZ")JS�^��PDϾK8b@ZU��1�]Q��6 O����Κ?�)�ӊ���eKr�H9-��s�2:��q���!K���BO�:�5�C:Ot!�A�ј+�*�8�A6	X�*U�W3��rE%|��ĩT�f	���P.�:�Hb 4N�2u/1T,�	@�W�2Aq��m�Ft�$����d:��b�L��E$H�F"A�|2��K�R J�I	77l��G��8�EoG�d��l	�#/(S`�ñ��^�h@
�74x�"F�� �����d��PI#C]?($� �̈́<�f���k������a��'���め�d�Z�{p�Ƭ���	�?)��c�C�2��z���Ȉp&G��95>�ˁcK,��7-����cbGt8pt����I2~�Q����$p`���"Q�}�X�W(Ԯ7m�Hч��O�����|�V�*s&x $�����~�D���6n�\��b<n+�&�*��$��"�:��w�B�aa�q���1@~}R/ҩx8�2V�٧+��8KDgQ$�,���c�����,\r��:"�̃4��Q�*mCN��gY� 3�4 S͓#b���Ƥ��^w��
"#�0��,q���+mBV ��6j��YK�E���+���E�RH��mGE���)ȼ6/�1C�D�ǒ9��b��HM�$���5A���t�(���4d�JT6�5�<�� ��/bA,!�󄓖
�L$	�+S	�F�:$�f��y�#^��ب�� ;6�X��6;�b���MN�%�n�c�#K�Tl��a��\�C�֘vdNT[��pV��?/̩����dL��(ue�	b�P��s�]�G�ڌ!6�κ�҂1�"�*� !����M��k�MC� �5"�O��╚v![6�qc��`�O&Nd��hƦo������^�(���Q��7i�r@��Ͽz����"K���IS�su�������$,6ƌ|�@�ܐ&=���:���R3��7�I�@��m� ��!X>�R��� �'��f \�
�`D�����w�� j!(Ģ�(T J� ��͝x}Α90�VB��2 �b0h�R�P�x)�)�:��'�ܚ.Z����E�<����3��6��@ϒ:{�ı���
�L�0I 0R�05�U3��ä�Q}����ϲp�R�j�bT�9�i'�5fF5��{�e���J� �
��x�� �u�d�e�S�fZ�0��M1dC���hy$?%A#�B�I�0�Re`�}/Z���Y�4�"p��*B+P��"ž�?�O� �O
~E�4[��i�L����;v��-�G�C�~���-�=���g_ }�4�B�;����D��e�M��P#��S[ȵYPǀ����r�����?1�%ܚ|�hP	�)���`s�\RY�$�K�F�h�M��;���[������@LH��<���=G�0��j		� ��O���'6�+C�R�y�����
�<MA�X�p�`t�àǣk�ą�)SV���	�9AC�H����tl^9j7����A��k�mn����G1y��yAс��n����>1�[�d;��� ���O?i/Y�hF�ۂA�`¥�"�+�����`�f�pq'b8Z�#���ip ����8Ô�#��D�^�C��	8^�^x�,�q�X��.�2!����U���	��tJ��G�ݭf&��1��"m��U��)2��EP5����%���L�8�ӻi�[�E���|��)�Rgr����xe�e/,�g� �iv�xf�qS���>zPt��矂fu��P�Za($��l�% �G]qT�-x�@Q6���`��6!��#��nq����S
�y��ӂN<�xJ�)�99�����T�U���3A }���_�ZL��=�-;1�it���3V ��k�F���n��ZF��� '���b��/I�ԫ��;ǪL���
$m!����&Z-@�̃!�/��P�*P�����(E,�A�"�^�e�)n�*x���qu�E�[��[�lW GP
��wm�T�H$�0j�%�5���g�8���Q��P�	S,`�ԫt�M8|������ ٺ1f�O�S)Vf��$I��5S�u
��	*!4�[5�|&@�v�aOj��r��:V��\��Bj�X@V�?* 0�sE��?(\$̒P	�)Yܩ���5EӬ���,�J��2e\)L�P[�-[�,T*آ@��*-P΅�DM�5G߲��RC�n��4皦Rj�I �%��`$��F.��Eu�e"��Ĕzi��8v�[:��<'Ϸ>b�0��-c�%݁Yp�1�c�2` 64gI��S��N�G}�H���̓6�Qs��K� �� #�&�ovAi��֓�̨0iP��(O)s�&_�zdnm9P�W�ڀ Y>����Q�m���Q0'��M.����E�5,�=�Z�[=���)�V�q��i�0&총���� �Ms��X�&Ze�Pl[<wP���ǚj�@"��Ϣ��E+Ir��Pȟ�e��GN�W��H�� 1oY����18��@B���R����`&��ZJ5+P�ډ!�Qp��Y:lU���1ғ8��t�3�I�0�٧3`�؃�ѝ@��,:Q#���U��ƍ:��9$̌#0�}�0�Y�5~���ȑ%Tt<R�F	
&p��E�2��	�%F�Qfx����'S(�i5���/6� |��ȰJx�I��*P��;sL��L@�;�$�F+~�:�H�7�b�����0Fh�DF�R�쯻](4y`�72d�gF�>j����`h�'�Q�-��򕓱Ə6����*�� �H2��� #/��1��S�$�Q�'}��"�^�?��`N�3����P!+���]��\ɓ��c��a+�

��ɑ=�N�(朡��S�T�ЌY�@q �t'T�����L^Hdr�Ǎ�y��I�B���Xp|��e��Dz����Y.B@��%�7ړ^R�w/.p������-^�DA%����i�7Z���b��������P�8�h��K�)+(�����̥Az����]/5#ڄ����w�@*�Ϳ1����$O������m?���Ɍ
:��Ј���?�ĀF�	#<�܄�LO�	���S��i8�����
;��N�
Y+�J6�
T�8]� ��7Q���D,v�A� �-� q��Ap�]��4! ��"ɒ8g&�9TGZdv�];�� )�8E��&C�G}�ip&^�#N�oS�s�nar�턭i	�kÓx�����S�n!bm�0�d!��I���s�a��者�5��'i�~�I0*��V8�K1�Z:P�&�����Gx�Č6�B|�re� @`��1 ����
��>�R�c�<`�����
X��A�(.r1 ToZ5�ZX�!F��T���a�%$b��d�i�[�%��l���d�%a�ܱ�n�@[7�7 �xRV�\)N�
�`&�7r��I{��b�ȝ��OPb�|#�j�$��N�~��#ńWiD�����p���,H�}�2 ��j�,��B�Ʉ
�~�q����H��� 0�\�`N���M; �T H|����p��3Jy�P��=�TX¤L��x�!b1�'��-�'�Ӥc6郐�
��d��\!2�V9�D�M�b(d�̿��2۴&�H��b^�����'o�Fl�B��D�
#�c���c�T�dߦ���D�pG���rC�<��o�=~�)��4�����5m�(��ǜz�� ��U�]@T�+K��@g�t��q��B.ڝ�4l0qN�Yg�'A�S�䀆]`؊@�k��� �DY�PFt�ǯ|����B�	{��Xz���l���PqdX�T�{��+p�|!G$��b�ؐ0�9�OJ �Lة&_�Y��W7�kC�A*��<p҅@�bTb�pa�0@���� &]�q�V�<�S[4D%(�� �*Ȥხ^�j�`��֋QI2�3�`#�t��A@'��r�@�"RI߳ ����״i�I C�ޟ/��$��2Wpm˦��6�����3h�
 #� 7o�i8�^�.��8�N��icGՏ6m>�(�9S����儽>a�AP<C�ܱ$E�!�����
G�3�k$��+G[��b�.Κ8���3b�sq0Qwj�'1ڤ�X��[�9+؉{�G�s�"YR����p<�T�ʤ�Rb�j��t�\�N��Ͱ0���&�z�0&ޯ@v�q�d�؎ή6-�6
���h�8j�~9�����p"eF��7S�5J��TH��ȇ�I��:������V�	EÈML�q�I�h��X�W[(����i!f)�p	҃O�&8"*���I�b��
�4�t�C�R\rh�(-g�vl�V�>`P#>�q�.��e����xY�w�
#���2�ZP���Ol�2TA��p{�U�UEh��4�̃P�D�Y'��_X΅��k��o�8�'���㧨 IR��!��+�b8��~��7�3%�Mj�Z��v!��Q����I�b�&Q�7��%��m���I(g"����7J4���!��X���"��ۢe�nT���K�s�xRJ.	��!�jZ���	��@A���"�@�1��%�!�&tTy�
�,��q#j��yba�X��u"ډ1����p#�6��$Xs�ء	v���ih�`nŀ���!T���F�62ft�pΈ#j8
E���Lj�I:�����g"�"U��4&�55vT���Iz/rI�^a* ��X;)���!�`:98�4OVH@3�P�tV.�C�� M*���ƄMLL�!��\��`y���*fXd��T�W���u���2�z���&�NFT�A�X)Z։'���eW��Xŧ��:�:��ri�)~�����>����!�J`H��w�3)�|���OKV�\��&�<`�)I�LC�%,���QKꜤS�L�Q�.h22�C�l�͹ϓ8Ɣ�H]�)P$%��`љe[�sl!�ܑ�R��j�i&E��=͎!��h\
/]0�v��cQ!�3,�!	����MI9���ۓ3h����=/��)	��P��[t	D��|hZ����_�:�0��]!F�J���%%4�����-�i�~dR�2�8� �ݡD�D�y�AЛp�����7DX�,A`b\�%
J\�� ¢2�`d%Qn��\A��D�����3mfj�B���c<�:b͊F�2��*E��`v��#%=ČP��mdb�z ����'Z���
^�	_� �l,kʱY�EX�S��^T�4���Q�i��y�ػQ��0D��hGfe�TU���
X~rm@��'WR�Q���=&�p�e'��DijX=�D}ً�DܒQ�R9��"�*�P�"k�;��1)E�:-x�邩)�~E�c�\�R�D�C�֜*�\�Q�6<��=�>��@Kb0�(铥*ֲ��<��艴%w�ĳ ܥ|�X����p=����-T �l/�h�J$�(��(���*�@�&����6�0&��(����R�X
!k�J(�HL )�ȝ��
Y�6�(����8� ���*����
��UO
�����j�8�X�#!L>X�����j�@�\+����u32�{S��6U^��JDaʷEGHi�O�����V�^�jB�
��Ρ3��(*Hhn �� 2JU�	�@)zJ7*
萫Q	$�@������T�r ��	����
�N5JA�7)���ѧ-��(���?<��`eB�+?[H@��
�ym�ͣs��T ���3��)�����וU;Ф��A�V��A3�o�$^�!C+@(�y%��6���xB�T�U>ڌB� ܺ��>`"�\P���&&T G^��!a���*T��6��xC�j�!+Z�����
�y��7\���;@�֙jeL���λ� ���e����q怓+��ñ�	�<wPI։��b ��"κ���g��b����ц�"����Ϝ�5�����+����"i�S���"Q�����"佣�Rz�[�%�yQ0�BR�8k��ȉC`� ���qb�d����AKʜ; �y�Hڟ"��,	Vϝ.����� ����yb�f��Ɋ�K�>�n�����1�.�e,�)�N�"$�X@a��E��L!&��|<*�K��M+�(�*�>l ò�
�3`)0�����A#N����9��j#ꚫl�(�$�L2��D�S�+4��c�8�ʃ�l*aSN�3	<)�0�Q�_ �H�&�7p���������
 b0]3�n�0�C�G1xE�;l� ��񧜩 �����L�#��LCR��rܱJ�؀��'��
��ˁ5(�x
��I�+A|� �N<{UT�n�<X[Z5B�F��ˇ%T�n�:��<�g�h�"��uEԠ#c����O>�8`��/ZQ,uR�ʌ0$̎ȥO�T����dC�1���B� \q��+��M�P�)�$ِ8#6�Q l\'<j�z�+ՅL��p��'�2��mJ�c��7�@e�t	�w8,K�l�%7~�:Ë����3��Y2 $_D���۳h�:7>�j@�Q��dރ@����ӈ
�02�b@��oG�P��?>������*���;E)�`���,�`=jU-�D�DY)��٢�H̡�nW�Rߤ8)�,�v��5���$G�� ���zЍ�@KY�$g�<Ygn�	�������
��}:��Ku㸘(��~؁���X'"m�!�.��Z !%��	`�:'�߬Y��*�΄�Vz� VAl�'�.,�%��>Z.��eƝ#�����V�s(��e�|zDm"�,W�1�d�;��Ҝ`[D-�BYZr�>6�b�cW�SdSX��'!�|�+���Ř���E��A�Й?~H�O�I��$�={Bq�ɟn��I���i$ �QgDȧ]��8�Ō$D:�!w���sK�p�ˍwV�TrģQ�q 
�y7��&\��'�ƈ� �=�U`��{���*���3g\��v˘�:��C�[�n���2�D���:g��ঝ�'Q���@#?H�:�@����3��
1~�$lӹrLi�(	=P��F}r�P�
�|p��O�8�R�_�6
��0���)��U��M�X��χ
�0�r�(�3Պ��`w� (e@s,�wCP��Z�Vg-�O� @�j��]����� �6�%�T��yJ>�@M�,ap�s����T�n0�c��)B�}SV#L+lه�2���#iL` 䴱Q㞚Op��+�H!=����4��)��<���C)�l��+S�b8¼1���v�<97�6�ND�ɟ>9�&�2qgF�<��e�+BΉ�W�ٽjh$�h��[�<�C˩	���%$�Gcl!�'}�<)$M��v��Tٳ(^?a�Q�BR�<a�cW,ox9��%G�)Vn�:U��S�<醈N30v�kchN��J�J�<A�C]�uP�I�CE�I֊�k���G�<a���Z3`,��B�0Jb\��@@�<�bn�$�t)[��2���"�(�w�<yt��,���d�24L�2�g�q�<I�^(=s�{j�m,���ƀT�<ɀӹT:`v�ŉ	x��s'[Y�<y^�~d�c�I*G�pA�CU�]��B䉲|M�	�'^�Sh�+gm�3n�B�]�ލɗ��
����!ңKlB��%:w �`������dk���!rjC�I�o�]AeH�aWx��T�.�C�ɵ �T\a�I�J�d�k��C�I�Wtˤ�#7t0ɔo��W͸C�I�jdl�t�3���qAS�E�fC�ɻ��-��Œ/v��9��ՈdNC��,j�3���Z+� �&H�'��C�I�R!RuH,,�h`cel��%��B�	�_�������t;�L"�C�� ��4G��HJ �������B��:��� �A	�5<��B�&f�B�	/vT:M0Åڑ%��)p��	��B䉣H��C���L�L���j�C䉯=��؊↦e2�X�.�2{uB�I�;�"�KC�?@��j�CRF�C�	�MvNP���2$�`4���XhB�I9fN����L�5XDғ�]�B�ɾx?V�e�3���c��B��0H[���b�šf��e�6�,M�
B��64�Ip��ۡ(s����#�B�����z�(�[����ae[���C�I
$n�Q�S$&ܼ]S��8��C�	3��B�۟�n᫣	�0��C䉫"����=�J��2��/}��C�	.x��ɔeޡy��ҳ�qM�C�ɂ|�-P .�:� �;蒒_AHC�ɏU��,�6"��6%�%���{��B�	�TTl̂Z�H�ksg]�Pޮ��"OƩ٦��R�����&��"O��CE���f�t���t�>]"�"O� �YKÅ��L�` �$�[ f ��W"Od�:�i�xԩ�5�ކk7|H��"Ov���[ \��ٰ���*!��"O|�2�gO{�h��[<��u�!"O9���X�f"��폰s�f  �i4���dx���S9C�̣�J�a��Q@k8LO�YIl�p�� ��'���reU�)����6�ƌ�5��'���#Kc�
�p'��[*����[�a3����I�0�R$�.�2����qyB���|��O���ؒ�Y�82p�{B�P "�c���D�%̔ȉ��^�r� 9 a�+M]H`A�HO�2�A3BRu�d�;E#�,6��d8 @Ә�~2�)Lh�Y��@��x��H'd�R��b��{��M4�~2�U
e��#-���I�@�}n�z�L��c|��k���?}�7&G!M�!���g!���#I�Tg~�g�Ѷ%ib6�ʜ>���E{RgU�ꑲ� c��@���;��i1P��{	<p�aX
v/X���������@C�c��hBԌ=��U9Xw��%� �@86T�M�� W��%;�GH$q�sSቁpm�`�b���C���oڟ A��y�Ό .T.���)��*��tK���jd�9�%���,m�+̴dxld��F� .U(���I,��\��nc�)�2%B�V ��Z󡟀,�ֈY�숞:�&牨4���M�Ɇ�CIҡT%��S�(�؜y��>�2="�BJ9�p���K�ؑ��G�)+�9��cX�@��K=~��߀1��	��	�}[B�I��ͨ�!=M�~,W�����HX����Ɓq�x���N 
�����Q�I�b(`�V�������4p���ŀ�� �XF�ҢC�����	[���A��a�8z@�0z1O:Z$�4p��s`�LR�)�D�Bp�GV8���YU�!J^�]�!��Ppp���̜S�9����Nh���Д$bڶL"�1��k�'Xh���қD*�y��;��F,�]��B�1��Y�ņ�#�>�)tb�f�V�����:��-�R@��x u)T��M��Ӵ ]� �/��)�нj���8s8M e��� �L�(:騵�re�/>�I���D���ɫ(R8�Rڇ9���ۋ;즕���R)5�iȳ��O���#.�u��@ei�0Y�HP��
Ta�`G �S�$�P#%��F��85FQs��x5	Ӊ2^�l �IPf��v�
��+�
��$H2�ˁOºm��T��G��)D�E�d��;�$���HN�]r,@�b��L<���9i��:#�v��D"Z�Ha��Ge)5��� a`N.�5��F�{^�zS�<��yY�"�K��f�&9!#
2l����2M�Y^����X5Y�@��إ�8��}Y�Q�����9��U�@.K�s��9 ���,7'���l�?eĨX�Xe ��jS�|� f��2�BZ�~�8-�L�gƄ5����<Tl�eL��q������y�%:�#4\̀�2��{��$��ڠG"d�����R�2H;�d̃��RDB<D0�!�./�`ѵ#ƍ?�����Q,̺�K�X1v��[��1�AP,��B��\8j�ȣ��2|1��-w���`@�:�>� oڗ"���B�̀ ��i¼��a�*-v��HR #<�(�ːo{��j�W"n�R�+�H~�:�"Z�Pp1��O�qa(�Ԁ�,u%��BEA�l�X��A#L
d��⚯PhaJVb�3-�A���Le��@&�`-D�nQ���f�"	c�Q��D0�"CQB^a]��x�Ä+Ym(3�׵RM��`6S9@���2�xU+����bX��pu�E(Q}Sl�4PH��Pf�̥�$����DA֜y"���g�D2X����>�D Y%=��	�@�ə5E�A��4�MKF�<N>���,��ĉ�ϋ8.���Î�n�� ���\�����Q>J6������u7gV�/���9%X�Ă2���Q[6���#۱Y���	,)����>5�5�E�8�ȟ8k�ś`':�XF�̇^)��3��0u6J�Q��R�d��X�e��=����r8Ԧ�-���%�����ʖWM��bKC��VA���y��da�L��>l� ��|�'�d���S~��8��.�6{���$ޠ1���hJ1\�2�(#�ΞKY�)Z�I���'j4e#D�a���q��ʹD��A�3($����%��Pkt�NJ̓$��D#���d�p�Y�B�	Bȍd�di�E�o@2�@W�"6�t=Y`�d[�%���R��؈h��V@�t9*����FkV��.�M�E������èG�>���iE;-}H��q��Q�H~"�^�1P]Z��X�WD�[!	R��a��`1��) �ĺ�ʟt��@�	u..Q�c"~�dU��QG�E��0?��(��$D��5p�d�k���A�1L�'(<�D;��>�q�K��<@��nq�:�W�&�*�gة���Ѭ%�r�bK������>�n9����[`�8�m'5Z��¥,u�n �2`1��eb#�ȭY���/F�)�O��d0-��F������ȳdO�!Ba	��[V���+ʉNՄ$k���Ԫb�ޡYY�oF�)c�L�I������!�a�d	4R�υX~��S����O�ѷ�F�M9�@pHȾ=d�O��h���0s��By��k�/�'<T�A�Ǎ�:,:(�W�ޱu��X�P6}�4���x��Ӆ��(��Z,p$�z@!�9bI@ы6O|ڰ�Z�b	#2��D�O�S�C谁2!��e��'	?�%R\l�E۱*]��|��P �7�*�������B[/7�'�������a-�'���h�G=z1Ǆ8?���#V��OԌQ��Fgx^���?f��X���?i�'E�8���#&����!� bM+b�-x�"�2ڶ�+�^3&иqF�E,��9��	�8c�q�Ǧ��c��p�Z-gj��t��rV0�h�ϋl���F��M�F�i.�țR�Cip���A�S ��7-e!v@1�P	�5�� ԴaBi�/�%�򤞲M�@-�mǣݤy0rI7�D�ӿk��}C�o˶8� �1��3]�0�o�:n��E�F ��b>RlH�˒'|�r��Vl�h`�if#d���I�]ڪ��*�G�$��QC;[-h��튙O��� �ӌ?�����O����p����.�h���&[RVY�4�����	�ҫ�%�4�E��Hl=;@
�2,�*=��#[SRI�D��d-��0�̆I^�����Q���px1D�8f|�`��N�`% �� O@L)�fF���F���K2,����W8�t�q:/Q��ڔ��8t����$��l���� �2Lʱ(C���臯f|u�"��)Ȱ �r�Ѧ��,C�i^�QE�fZ��K�#Ѝ\�:��V��#Zd$ۇJ�� ��Z����y��I6�h�'*�
1��cC��u�jcH�;.�U���=7���� �#b;�0���&Yr�#�+��u�Zf���8+�Yꥠ�=6���H�t�? �4�D�7z�{!��	D�ԃ�3 J.93gп�*�X��?�O�Z�$bA�&�(4ژ&�29�Q"e��H��Ã �\�˅J��4
��ϧM6,�YBj;Y�45�!#ғ<"���!G�����U�ЙDe����';�@�����0îV=�T�����V����q�L�7�x�����+=��G62v����M+~�P�2a��M�rh+�Hl\�3�JT�恘�DH4+�y���W� p��V枉	M��y��|Ip	2b�Xhl��� d�0"�Q�g� "t��;{$ $Yҥ��j��)ߤ`)�+��˹OTўTI�%�Ndm�iJ�'(DZܣ���/�D0&H�C�0��"D�??s6(����OzpAԍ�+���g�,� dp���G� �λ<�j�@�FӖW�(�#��0�͓o0aa���<C�(ҧ�)��RR@ A�A�x� ��Zc�����ٺbD�h�/�
��qF�*8�����%���pa�[G�'M~
u+OS����e
�=#��	�I<9���{E)#ԃH�F�x�A�jV�Zɑ'$��C3��r��D�n�DЙ!ƕjK0�3`�E�>'^���D�aX���	"!�l9�^�Ī��� MJ�XBAܢ#�|��/?X<�t�� �-2�(��h�^��C D!NF1��(MX�d��1�`׽Nӡ�$�-��X�����z�:�K��V�<d��P�����v�"��B�T����MOm��!�*�+�< ��*b��LЖMK%�ЬbvAD�5A[���0<)�2	$�����ڨy#vD��Fb�����G�Tg����&V��
�yGvS%�J5�0X��%��d��ո7$p�'�2m"���=n+ ����Lɦ���ORL`a�(��m	�g�$H�HP�g�:,���I�զ��di�o2��Q!`XI
�ɰ�E��x��]������`8�O�D�ba�l�0�����]���[�i6-v��VNiĎ��e	�;2��P��!G�j�*���8Z���S9�ܽY!��~��������jq�'�کi�@I3!4\��a�c��|��Y��k��Xz J�~�&���4aJt�@`��ZE�/�'��9��v�๥M^�
z#� ��y�?��GV7}�<�	�� L����6d� /t�:�j�/ml�9��@x2g������?Af���HBD���	�U\�����Ӎ��Ē$��=�8�B���V��yVF$��,��L2�cK�c:z�P�( q�����=j	�%��M02��(���sfvM�f ^8� 3�k
�	0� ��q��ɘ?V�!�D�>A���j�.�(������J���)ɩ!��e��Y�9[���@�=G���2R��U<�HA��!�@y��I�
� 0/��~�l�0Z� i�g��`��W�T8?�6uڐk�� u�(x�F�3y*R��S����q��l��BT::�,A� +�pࡡ��<iR��[�D��'��-��I�2��UY�.LL/�����W�{`|A��J�V�`x5���kN�ܩ&@�z���q��G�R�r�����o����oK�S�n`ȗ
iI��' �$8�A�=F�4��)�͎y�O�PI�gS;0�=���":��g� r,����Y#�q��@%�.ԑ�	�7]BK�=�4��=7��ceUd�Ջ	Ǔ#�2��"CZ��ta�R)Y�B� ⏓�,0�q!�֔+���RTB"�4��b���z}�IثE�44a"/R.jȠDYQ��\�ʼ2�(Χx�ҥ��L*�O�A�"�Jv�&�1t�YM�l3�+�0��a�i@�k-sӌ	��Ά}_����!� `ͨ|��Ù"Z�|��'H�
d\U��=|hhTkӣ	O܅�Iy���4�V�F�0�#�	&]�PD�G<^:95D�?�M�A�E�t�E!R PAa�CX5P��醽\6%:E��V�D�eTf��$b��k�k��kW1O��{�+�4�M3�,J�6W�ȡQ�3q�~���틜7͸h�5�U�]�D@�B�̌$���jԤZ�By��i�&*h��`��*)��xb��
z2�E0Q�R�g�<@���$�~�m�(��S��@8a0��V"�?�2���	��vY
���i�N��G�R$K���Հãi�����K[>(A�e�E�c/		_�4Հ��b���c6�P'=����u+�oJ�} �ʈ9`�e��	�^�0٠f$�f����;�:H�d�^�u�� ��hV�r��	�<?ra�T�Q�p�N1�q/VdN�����a� mSWʔ2�va0čzTV	y&o��s�Z���bC�Od���Ķ>{r�A��(���?�G[?<�4�NE'Y�㜬y�,���$iVda�m+"�\r�@�:���1B��B��R7�'��0#��Ҹ i~,��-��w
�u��O��HbG���x���\�`�mr�DL� �)!�@�K���yf��7q!z\�7dJ�J�P[D�'�!�dZ&�"Ę����k��@���R=.J�!R �K��T4�Q���
R0՛R�X!��ID��H�%R�0�2�R�ʥY�b	�+�Q�t��ɂR(�2'+H/Y����F�s��H&�ڈa���ѓ�ƷM��5a�c�	`ؾ�p&Jݝ;QzP�4��C7���Z�c��ə3�'��h��c��j�V���K �$��{��rQk����X�F-%哬Z������~���-у.�JA��$����g�z��`���S6XzA� �or������XN�u��n�b�ЅC��O,o�r컅�z�$#�O�W����6I��[G�U�n	0f�½;Uoίh�t����ʵ��I�6�ڀI "��u5��A�&�	� ��=kq$	m)2A���W-V��:���1��h����,�¥,E��	`c�O����ɎR`��F�"U���&��q���pU!�/f����R�-����@f�l� ���|R&фn�*�:�'�,j;*i��J	�mi��*���M�E�G+��$��E�3y�9SF�pLΐ�rOP�(C�O���f�uu�\В�Y�>�5�uCH:#lRLmڼ/p��%,��m#��d�B9����r�IR�( ��BÂ����峂�i��UX֍�; ��M(�cR8{Z�81C�$�t��h��8��л�j�4��Y1��F�<�R9�S�ʼ?�6ë��"����Kr�8�ɓ-S`��E�ǋ��s��̃;�8�޴i�r��փ�]HC'ۥ�a�F����f%�1T�>� �y"�d��� �*�J-T�J3�A�w�̦��'��é�K�l`��5S�>� �]�O�.ț�,ӈܤ��ǹ!���4N�?�$��@	>}r��]�J� ث���
Ơ�#gF�$�����X��B��#�\���J���XA�e�ݮ~ȁ�s�!?M2(�ń߈Y��b!'(�� ��3
4Q�*=�]�B��`��!<=�RMU��0T���S�HN��j��U�&)��C��|�Da�>8����UIqX*#�?�v��#�Y�0 @G#6���c�͖�<2�ȸ5�B�yL=B󭍽�vѰ���zY��]�(8JPsU�0a�����)��	�"��7R�pSF��\����rO]�,1^b��K`AhӎlR��0U��Q�N� %
,�Vm'@�5S��ܷ2�	@b�lݔP2$�Z�U��e�n$�.ڴaV"=� �\�'�=*p#�.Q��@��� ��S�i1��w�P
D��PA#�Y�2!M҅Zt�I�ꑰ>�Խ��Ap�"U(Q冝Q�ۋy�%V�!��8IDi�MӇi@�����4 �RX��I�tj0�O���哄6�2�8�*V�Z̰f���R>u��ԔbEK�gVڅ���E�;WD�W��@�rHHVe�	):D0ȓ�E�x=|u���bZ̭�" :V�t�VC�fx ���5��+��܂%��6K���c�0�`�r)-Z��}�T(�P�2�H3��&)���҅��4N���3��w�R	ɖj�:E��ȃiɐ1kB� RNl�Č;�/O>}�� qc��'�T�*Lx�'�D-�`Y.j�8��̆}��\��(���v��I/�x�gk
�y��-�B`X,n�(����y��|��h�,�!�D��{d�8��,K҂�ր_H4ѓW!V
�O(�R!��[���eN�,��l�e��҈�8�L�W�|�-G�_�\�!��
S�yi%A��hТ %%٘�`%LU�d2�͇/Y�L�E��{v<�)gj�v�Pm� �i��w�Xy�F��(CYP�D��Urp�t��/Z��	y��A<�JA:���V����i��S���h�%pu�`+Ŏ/[���E�,��)�Ti��G��n�&��	{���/68~��8�O~ �����4��'�H��^�<���P�R |�Ҽ�*�j�	��Ȍ�P �7�
8�DE}�ņ$���6�V	�t��^�m�$���&�'�v����TB≭	��:Q(e����Ȫ1A��F�	b��_���:#�@N؟t��/��2%zԠV$��Pb)3�I?~�T��ξm` 8Ф�у[�O����u��*?����>n�$���'"B1にI�X`�@���Y$�x4�3��`�F� E��t�S��y�J-o7 �j�/L�)��8�d��+�y�a¦}t�@��I(u��ŕ�y¦M�"�h�(&�U���Á ���yB��?N�
���G؄Bi��sB��2�y"�F�q�P��c ڧ(�x��KE1�y"+G�F$��V&a���*'F!򤗄���Xi_�d����J��!�D�� �$�ʆ�ОS�n]h�C]�g�!�H/Ji2�Cæ�6��}���c�!��:*ܔۓ�Қ$*h����,V!�N�V�(�R�irA���_w!�DM�u�p�ۗ�R�Pؤh�fJ� !��R�ob�x)CG�����d�8�!�$�7x�%D��q��� 5T�!�dڤ 劬!S��,hXY�㋛u�!�d�\��e�dc�uU�$��#�"S!�ݯjz(�+��� V�9����w�!�$�g։�F��]���f�!!�D�;9e4���g��~"��y��_)!�d_-mg&j�("��� ,��M�!��R�.��A�47�%J�B�p��~�坩sT�bs	X&{���4�Զ�0�@��lH<	�iެ:`P8B�U�k�ؕ#7�X�}��ɢ&���}�a��ʚ�Hp�#Є�0TU�	:tD�.���E|�BN�O(��pai�.%�yW�ە�@�Ӑ�\����Z"1}��O�baɵK�'��bҨ���0K��d ��(O�'X`�Yz�D���	��Y� ��$����)��+���*�BF�\�S`�6F��˓�t�t�E%ʧR��{��Z7FS~��eױcUPD�0�Y9OqO����-kw����@C&<D2��C�&D��غf�9�V�M����i͋�QC��ɖiI �O<x��(8�q�o�a�O����« �����?X� �O\	��T?��H<i��Ȇ$�<��#����d�7��р�'xc�"w��Lj�dRE�\:w��h���"�?ɴ�"qֺ�D�d� �(8 !�,i$j�/?�J���Cy���"���]���'����k/0�㆕�%�byS��ۦrg�7ͅC~�mE�n�ș�ᓔfJ���g��#�:Y�Rƈ�?��M��S4���2G��Ok�drb�5A�҉����'�� S��W dY	ݸ|��}�[���'���D�����4�ЍA"�08�&��I��#��*�-��Dr��O�+��`�V,Q�#z��g��7��O��w�OO��weG�&�kʅ+����|K�+����'d<Y"Ȍ=/$�quC�6d
y�'z\L���Ơ%mɧ�� d-���,�8�ۦ�B���U�Y���DOۢ�ا(����T6�9��gE�V�J���'h�Cu<�)�'z�0�+��G�-J�*W�< b̩�)�?��'r���(Z� �E�ĵAxB��r>�dK�K�* ���c�_'D:R9��%�J f���ד?�f���
Y���y�)6�FՄ�N؆@I��X�i�N�8���,vLra��EV�:oҜ0�l|h�.�%x��	�����)B�ռ&g�#2�L�y�p	�ȓ|W\���f�&+�]C#l��h-����e���ӣ�^�Q�|0�A ��$}$T��)�����#ߒ�9 #c
�+�&��ȓ(ּ@�GF��+ȱcdNE&�:Ȇ�FC�푵�>A0�`g�# ʚ���E�j8�8,�����ȑ��
��ȓ>_Z�@G���y�h�rl�0\h@��ȓ@�4����P�W{l��1�+4���A�ٙG���[q�AJ�%Ŧc����q�j%�/[�h!�9�#
���ȓwV�(�ppى�5nZ��ȓk�x"�ۖT&�)����]�<�ȓyk�|(�.K�M�0�� �%�*�ȓI`����W+�,Q��\8���ȓf�D��* 0�=���5<��M��m��(	c��+.D|i���<cTdȅȓk3�0 K�A���S�Dsn��ȓY��I��O1����ݍ��%�ȓX��4Gi��b��-В�K�d��!4��0%��~�E���oc��ȓ	�B�:֬�$3��"��
�&ԅȓd!\����إD|�9D�Z	r�21��
��8wO1z"!0�ƛ0�nɇȓ|�Xc�@�;J5a�&��q~���(z$����$�� �(��$P���ȓ5N�@3��Y�|<��FR�P�V!�ȓN�� �1%~\�� 2MtJ �ȓDX\Ct�2 a
�����#|��ȓ~��@k�_;Z�Z�Ro=��@�ȓ�@���[�S�24k2�IAz�ȓN D�Rς���j�C��L98��g����
��GϰHfF�:-�ȓ��ɑ�q�p8�G�@6G/`�ȓ�Z0цN�9ڂ�#��1���ȓ+kJ�h�-P:���7Lv���"D�T(�E��O�#�|��2b(4D���2���>na�Ğ0!ۚ���!&D����P�t�L��!W�\7��sR%D�X��KT0�p�1��^�jQ�b!D�@ZV�\ .<@��c@P~�yTa>D�$�P��{��,��M1!�V�ba<D�`���?��Y�@���2b,&D�X�a�D�eCN��gE-O[��'`.D��Ʃ��1�Բc*q8��g"(D��yW��Qѐa�a٪�@��0D���ȕ�a`�p̕���U{��/D��c�P
g��-�����Y�tl)D��C"�4-����nRbF�Uj�!'D��)R	[21b��'�����oRK�<i6���jR�1�N�NF��RA�I�<�qǥY�F8�hӻQi��B�f�A�<�L_�+�Hm��Ԟ"uf����~�<��+� >	ٵdX�t�dBr��|�<��� �&tx�:��F�w��5
tl�w�<�Q��hg�`�1��gkr�v�<
Y R}Z�#!�J�]CD��4�Vu�<� �x�`@��$�r���_����"O���B�C��i�d��{b��a"Ov�"��1L;J�C��@`^��t"O� �p#�[9�8�Y�,Y0i��"O.lr뜀$�r� P����b@"ONQ�!`�/"0��5��7�=�b"O�qϔ� ��Lꢁ��1	d Ҵ"O�!�R�R#O�Y`"�޶9�r�e"O>� b@��Vt��iA�X�/�>ezs"O�m�o]1��`�.�7"u� �"O�	C ��,ZD��,M�qrኁ"O��0���A��E����+i ���"On��!��Ҙ`�*O2LcW"O����+V�ct�"
I�_��`�F"OƥY���������>xK,�8�"Omirn;w��1��� I��Eå"O��s�ʙ#��M�`���h0��"O�5"��H�@�d� ��O(
���c"OR��!
�=�	Z��FT��"O�ջ���
�t,�ƥ
]N��"OU��ED;CDd���OC��kB"O���j�`��z��44��S"O2y��M\�b��:��H�^�~�`q"O6�q%E�~� |� g��O�����"O����hI CbP�`���5�V��"O������0�����zh~���"O��S��@��xX�rD֦B���2"O8<#L=��ȹ���DД!
�"O&IB��Y���Ic7lU#�4e �"OJ #�*_!X�a��J-6B,�"O���P�-����(�
˄��"OZa�#!�%C><0sm�t���2�"O���W��.Z����9�ʑ��"Oj������P!!'yĨ��"O���H%�N�GO�Xi4b�"O^ؤČ
и� c�gD@�k"O�4��ꄮ�@붡O�XAn͙"O���f	�	�>�K�퐞I��,S6"O��R�	��&lӆ-��El�LJ"O��B�jX�����D��AB@p�"O����'U4��c�M,/.����"O���e� 0��X��\#H�  �"O���6�B�|"���D�;u횘a"OD� �݌#�reV�ȉ�ܳ�"OD���1!�Z��%��v��"O�� 1�0+?�x�sBC�v�� #"O�-�d�S�_��i��a��J5��u"O�m1q��]��c� 	8b,���"O̅ѐ*��?���H��܎G��%�G"O09��N-K'6�8o]�YW�U�"O$ :�^9���f�F)!I���"Oܝ��Z	�옐��<H�8|��"OBm��Y4p�щEl��8����"O<+�L�:n(�X6BV+g7ʠ�c"O��8��U����V4"̋�"O&t��aF�!�������i��"On��bbU�'�*H�O��
���"O��3�� 5q���5OJ�\��Yt"O�%A`����z�@	)R��u�1"O��aC�^�|X��J\*K}�x3A"O��Т���G��!'�ʘ|M�"O�q�#FΡwSR�pBJP4;o��&"OH�)�j�
���B�R�<n��C�"O`���@Ւ��̐ag��7X��"O� �`8�/^RX�h�@��{͎��U"O����ݔJ0��)�^�(c��"O�89�M�+�,YȔ�LK�屗"OZ|�A8b�e��R
2̈��"O4�J�L�B8A��eOpFD�3"O�q���?xp��禛3B��0ʄ"O�isR�V��Y�KŲn�h-{�"O�m	�b�;D�� �D�Z�&���"OHl1��J25�
 �����.y��KU"O�Ӂ�$<�A��̃CWDI��"O� �TC��01ȵ���-ye���6"O�(�e\�	����e�A#E[����"OjuڲA��f�@�&3Ba�'�/D��� ʖ�_����.��Q�ƽ#"H/D����@ʵ ��,�$&�..ƘY��g0D�̀MW)#n��;B�]��-*@�.D�(���[�Tߜ�j��C�HL�#��)D�(JFR�xȘE��	�<N<�Q�'D�� �Dŉ4���Hr�)�n�1�,GO�<iML�;�(3ֈ4��c
q�<ID�ܾy�<��f]0�U���Ks�<��Y"2�|����;�Ф��!m�<1���o�B5����<ɢ�x"	[a�<Q�	2^�$|	p��>o����c��R�<�1-\�t<l���˖�l�ɹQ��Q�<i�JΥC��Z�k
�
�|�Q���u�<��Dr]J��@O��Iu�Q�'�y�<��gԈ+�Z��e��L�V��kDP�<��M��s��K�	лe�:҂��I�<Y6BE�+.E���y��`��o�<a�Ǒ	��$j�'�-j�J}1�%�g�<a�3!<���P	٩\7��$�]�<W�B4T��L�9�F�3!*EV�<9�a�'��YC�՘R�D�q·O�<��Ϙ�*�|��C�w.� ��K N�<����d���
DmT50���R�<��B�n�� ��o�Hȫr�AM�<QH�.rF�yC�l�t��9�u�<��O:���t>犁	��i�<9��3M��E)�
ٗ%q���@��a�<�Gͬ]��c#��Z��Ȓ+R\�<)� E;x.$pA�E�5$,6��n�s�<�wN��s�z��ð3�2}���o�<ш_$- �� M���� Rb�<�d	�VRƬ`���Z�~�K��a�<YF�ȷq{�5��[.x�ՒV��\�<��B��re2�����V��6`U�<�Q�*�R�1��/��i�`�{�<ْO����VB٧8C����q�<a��	r�&(��-�"ms|�!�)k�<I��=B�bi��E%�(q�B��c�<�k�El���$�O�"$h��_�<��,UN�h"D�	p�C�'�Y�<�-�Y�j��!��jDx�+���X�<1�T�l��̙T���1��xK�gGK�<i�H&|W$`�*��Xt�����<��*�6@�h��1	�]b$�sMK�<����~xv�i��I�~ ��a�<�T���������9
��]�<���Y�GN4����c���1�DU�<!��.G��9����(�3kO�<�P�H.?��aIֆ\���	�@'N�<ad��� �&Шs��>�*�� o�<�c_QKD��W	9ib�	7ɟu�<�  ��P焱c�&͠�`u�=b"O�uDn��79P�{��%:H:�ڲ"O��X�O�%����a�TKP"O<�À�\�I�K���%9����y��Ee��i*CE�u�"�1Q�I�y��Q�|N���A9ry�a@���y�dʒ(��]�5�S�x4n���O��y"��R��h)ȇi'N]�L��xB�'���k@�D���Q�K����-ܕER�mZwx���	�������ͪ��s�k^+�Q���8��s2�V����ж"V�; A���'�%�|�h���~�*8��Q
-|�1y�W�L���9�J(x ��!�я'��]i*̈́D�j➸��X�zL<hqQ�E8� �1��ڭI���Ӧԑ>��?��}�@Fc���C�9�����
�5���?y�43����5)���Ɔ6?]n�Cc�'8\6��OL�l��M�+� ���"O˦u���̉)1��})�]�GIH�BpD! ��؟4I��{�T ����2�12�N�j:u��ȃ'y��B���|� ����S�M��<�f)B��)C���O��hӴ�K�rZ�kbn'T:.8�RF�� �n@)fC����3�E.r����צ���'�2	��F ^��`����3E���{��'��i�e**�:Q�U(XF�{��u�ƙF~Ү��pl�+R��d�&ȉ0+��@\�j�.��ΦAP-�4�MC����|�4{P̵C���X�L!��/g9:@���?� F	!�8�B�w�
@l�b�b� ���4��Y0j|n0��C�4[\���\5��'*R\�0��zI��jE���V�&`�c���2�$���[�?M����1m:I �J�6v�a"	!�dΕFKs��>�I/�Iҁ*m���ۣ�4�1B%�qO
��.ړ��d	s��Rf6߮��Z��x�hu�\Ul�A�I=��y���@�ɢ�'ULJ@9�i��U��p"C�?AGz��R�-B�y��˂.h��`dJ�	�q�a�د��t�Fm݅	3��@p�?]�� <}f�@r6��P#����[+����U9+��� �CI�T�����$\�E�n��tI�R�)?�T�#��杅@���a�E�x�>	�w��$qxY�Q�iz2˓0$=�i>���ē9.ƹk�Ô\�9��G�,JG@9Ey��	W}�h�6R<�c�R�<��@�@H��'�M���iA2�m�(ʧ�®��)�e�'$�N8:P��v�B(@G X�� �4��<Y�&Z�I�W�3�F�Ô�� �}H�B�(�r@�I'L��;r��PE��(�g]t�'+eAd��=u���J�@Ȳ�&��FӀ�{�k�2�a�*]��xgH$�\�=�5d��*����K�-���Yԉ�0[Vx���M��Ic��f���*ל+ˌ�R�G�Z�AO�,hv�M:I���2��Df���S�O@���M�E�i��	�_mZ5�ܴ�?�]�$ p,c�e�1� qh�gbʢ>A��&�z��L�W�n6m@L'�����.^���ыy���𐯎��X� ��(O*���@�E�zq�S�J&�L����&��Y����+t�΍�^�n"*a��/W�b
25k�{�k_��?�1�i��	�+ת��DcӖaRf�#Ө�y�N������T���'�M+%��m������+(���'g(<�@��Fl:(�u#��*��i��]�-dv9P��i�rA}Ӕ���O���7���>!i? &  ��   =    �  -   j+  �6  %B  �L  W  a  Qi  �t  `  ��  6�  ��  ݘ   �  a�  ��  �  )�  m�  ��  ��  3�  t�  ��  ��  ��  ��  ��  9 � ~ 1- C; �E L HR �X yY  Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�� |d��"O
`�(�;���8���-0��1%"Oj4��ND^[��"3/9�0|H�"OB���H��*�ʞRy=a"O�味V�!X��!&F�:J�$���"O,��a
���C�Ą�M�"O,$3%o�-���p���+Ն�:1"O��ݢ1����`���y14]2��i�<�6��{_���c�H�`�fX�$Kn�<��A̼VI�xR[�)�Ć�pඤ�ȓA5��('nߡ4�� �)˩%� ���,��r�؊b#`T�eT09���ȓ!�b��g��}�8�F��-? �ȓ
K|m�ș�VṔ���2�%�ȓ"R�X�j�4JN�1�˘X�i����̹	_�jZ��1!g��zܶ��ȓgil,*�J�
j�Ne��i�J%b���f	�(U��:���G��$Y^م�~r�� S�%T"���k\�jx�ȓ|4�1�îJb��@ӵ�ݩn�V��/[`�"�v4�R�!ʎ<��M�ȓ`:��z�ؚh�J�Z��$HY:	��H��p�m�C1��!��B:��0��EnjZA V;9����J[
2���	��4'J�EA�IVW&��~�(aZ��ӹ�>� o�Y�|�ȓ�f�A�
Ο7�H��M�$�����mޠP����/���ANXo*�ȓTv�����{ ��-7�*h��I��sB�8�8���3����ȓNe*M�悡;������X�o��!�ȓ'lj�#F�m�+R&;�|��2)n�C��0S4���T:
b���:�0!��e֊��)��ͷV��,�ȓ0�&�8#���� ع�L�����;�P�AFd���,w�6d��r�EQ�( �gVlɦ�M,H��,DP���|�I	$G#\���ȓ"�)���E�B	yt&B�^�LɅ�4�� ��eëF�ڙ��n��R�p�ȓp`@}bŇ�=�$�AUN��P����L��p���_�a�)�Y�!��-�?i	�H���iD!���QԨ܈?�L��sֵ ��GO��Y�
Q��-�1ar�N!�$�ӥ�X�.����Ɗ�p>�H<Q���8fr�s�� ����Fh�<1�Mn����M]�$��8J$���O@�=�O� �HVhբc���Pf�=������O����&H�Z\�Q0�ӧ"qFh�p"OR@r�Ε_���*���v4�#��>����)Ω8��c�D�,j�^�`��ڢ
�!���:�&/;Ӛe�c-�%s�D��0?i��ZM�D�ǯR�D����U�<y��0`ka�*���DA�X��ȓ�6��B@UGZI�]:�Խ�ȓ9)��F�s��I��+H�?*,��}��r����vR���� /���鉾s��<�ݬ���a�lM:�$k�
	�C�I.^�r���%T�h�+Lr����r��*[���:}��M�~��
^�^q
���!�`��妉 :���dQr~�(��y!|�J3�^�h�B����~��j�H��I���y��j_:BU:��-W:�,�'��	A}�_>���A�|� 2��4fl����GB�����"OXLq���(�@
�I#��B��8�t�c�4�?��*� )،+� ���V��^(<i��_������^-���`a��B���^y��'�����F)3k��)�ߋK@0��	� f��{"�\�D�J�(�M�@#rM�#�ٽ�yr�ٮA���X!��B+Y$AZA�{|B�Sz��Ac5D��@y�y�c �-8b�h��I�|�5��,I�Jr����2
�`�'���'y*"}�'�ƹ곡G� rTlS�e8�t��瓧ē }Lt��$�?{P��#�da��l�>�V�����hI0��q�H 8�4��ȓYnl���@E<R��Y�ӂ��0��0���Fq~b�)��.>�A�Þ r1Ll���Z���dtӲ"<���M+�y��L�x�F�Z���wjs�bՒ��'	±��I�GmV�IaK`YX��}���@F{���6M��"�Y�5c&X2@�ı
�a}2�>���M�M�ڍX��+�DE��Gx�<�dɮt���W1 �`�@�\�'-ўʧV?�Ż����Rf֙UAn}��Y�hl���4H8Nm s(��el��ȓng<����7=�n��w�أX�&��I
`��L+.��i� Ɵ%Э���W��S1�!�"�-d74��F�q!��?	�jU��#[/�k�OÅI��m�ē$>���@��E��d6|����<!�}�i�;���� �>}�,��
'�yBb�-�Z�q��6q:0��a�����)�S�O٢�C�Í����h�HU-��ؘ�'�@�[�M�i�	�^�Z}/O����#?Y��5��2H�N��׍�o�����On��L�fY1i� �$%�'^��"�Q+y�d���i���h���$��ȟ�8��Ն5(Թ��ʨ��{�"O<�{��ߖW2�qpU�ϭ^�.E�"O�,H��BJZ����ɡ~���S�"OPISb��9}��L)s�ٰ<��)af"O2p� C��)�N)�%@�7O�i�"O���րJ0M��aw`��0�~}�P"O05sU�'-ᾠQtO�2([\�d"O^\����;&B�� �ٯ2B��2�"O��XfF�&X���0�[HX�ɪ`"O�ܣeѬ���)b�H!]NB�3p"O�5{G#�;U��aC�N' Dڅ��� �0|����:_j�{�%�B��dJ��p�<!B@��2��t AZ'Z31�E��+"�������O:�Ij�*3��}�g��%h��Q"O,Dx
�t��!�I�a$	+�^�����������@Z���=��C�I�R����̻>�0b�!=i��C�	��(�`�#��AlpPp�¥C������xc�,$�flj䀈?\pW�'D���"
L�
� Ԧ\!��ġ%OB�=i�;:k3��v)�Ыgn��<��f���J=1w�׫F�
`3T�Or~2�)§p>�Ѱ��ja.�Zg�G:�d���#_�Ũ7�ƻ ܩ��O�
\�j�&�<��"3=��Z���^�X����x`�C䉴r�f�
f��Z�h,�� RtRC�Ɍ)��T����+��\�CJ_� tHC��+L"�H�RNݜ^�MQ3�_�� C�ɖdGD��eMC�8�xq��tI�C�I*~�V�R �"�����L�B�IK��v��/�Ze{���_�DB�)� f��PZ	ҰH�i�-�6k�"O��S�E]2&y��ݔn�ֱZ4"O���Dh�K��*b����mC�"O<��%�B2j�3��X
�F�Æ"O����@IY����'�*�Ba1w"O�y"Ʌ<
�ܹ1�{�lhf"O�qy��N�6���)�9z�<���"Oҹ�aG"7˴蚂�
,OXq:A
O�7M�e�.�� ���#c�'`���1���6k�0m@Aa�Ĉ#'X��M�'%��1S!�z�:�#�ˏtPU��'bz��nC�4k�D ҌQ�ļ�hO<��O�b�D�=�P)�'E+��rC D� �Hi��	q�<ɀ��>z���;g+�/)A���A����B�	-5`t�I�!�*&.��1 �82��J��T>���}�d�kn�}��D�@?J `S���y"h�-H����a��6�ب3�I��	��p>�W'�7EJ���F`�W/<�!V([L�<aa�+}�̩���Z%6�8Ia�LF�<�SG��TK&q[a��it"Y�$�@�<��J>kBr|+b'~���bk�y�<iqf�}���2��G�hEAJx�<Ac�D�r��	ZW(S�Z����!�t?���R�����&U�)���r��C�����U*�qԆP�����C a#&��ȓP����qQ�7��:�Ȉ h�H��s�X�붦�6^D�Gj	�QĄȓWXX��#�=0�BQ ���ȓb�Tq���,	j�<k���Ia�������8\�`�[;E�\U���3#7X=��l7D��ۗ��JbZـ�
�����/D� �3��G)���a���=ȑ�a�-D��pV��Ii�Ab��4RȥJ8D��	�O������N�1+���Э5D� �톢;���3q�,;��]�v�4D���ud:R-��PB�,촑J�4D�(bac��h�t�į`�V)�C�7D�seD��V��QIM"HP��!@8D��[7�W�9rԑ)�h��p{vE(D���jN���j4LNu�$@� (D��bs� �"*1R'
؛]�:�ф�*D��&E9un�3�[&Y��}��+D�XXC�»t�T�1�L�hZ���'�=D�� @�'i
�vIgE���n/D�x��9dTtQ��~u��ht'.D�4�Gm\�$2jr�.A)YK��X#(-D�D�GC�x� }coѢK\T�9D���W�N�U�1T#rɻ�5D��H���.�(�&��Gcji�4�4D�$���� !����f�PrOT�P��4D��`˖<>D���M�5�ӧ2D��9�I@/!���kB���N��p��'1D��I����Z���S�K�/�n��-D� ��K�'t���w�N��L��*0D��g�ІnC���Sb-7�v��g)D�X�r`D�(������ wN��G	'D�Ę��Ȳ1�<Q�tn�QU �aT�!D����,N�"��F�ȪI5ek�h4D���Rha)r��B�f^ݰB�?D�����${Z�H�� rG�hq�;D��! �/k� I4�
�4�$�7D��kׅÈk � P����4H���8D� [%�> ��Dx��|F`6D�8�F+T�|�z��D�\,[�\�W�3D�� �x��J*i Fhc�&�8!b�HB"O ��͘ x�:5R����A�r"O����Ő=
���#I�~��|"$"O�m�"i�'ߠE1�녛nu�p �"O���z�}�P�3rL�t�'���'���'y��'Z2�'��'�KU6"�2��C�L ��Q���?!��?���?����?y��?I��?)bbɨ^RP�;Wg� �Hcq���?���?���?9���?���?����?iE��FkD%�D�
�(8)�&��?)���?A��?����?!��?���?I'�59�Ԙ
VjCx�u�A����?q���?���?���?����?Q��?Y�N\Y�a߅%^����ɹ�?9���?����?y���?A��?���?q#��	b��:&�>�Lʄ�P;�?����?����?���?���?	��?yQ"ՊYxH���D"*�,����?���?����?A���?���?����?1S�܄t�R\ �,�^����P8�?y���?����?����?���?���?qb��vu�l�RT�&1Td��)�?���?I���?����?	��?Q��?Q��ÌN��� �ĚF��b̞�?���?���?Q���?���?����?a�K*^�> 3�գT�r��_1�?���?���?i��?����?I��?ie�thZܑg���,�q���?����?���?���?a�H��6�'�R�T�h �`J���.tf�۠��-�N˓�?�)O1���#�M�1��#}y�[�+�����[Bg;31�'H�7M)�i>�	1�M䪁��`�fЕu��b%-[9!����'��uIcDõ��$�3W"�I��]����بi È9�"�ŔZ�bb����Ny��4%���pC��
 �q�d��+r�V�۴N���<�����t��NLB=$�+0']u�J:a�:SDQl��M�'��)����Kg
{��RDB E-�,�� �6���~��R�h���AoSj�����'r���l[48��hKQ�� 8���1�'��	Q�I:�M���J̓+��a�X��2E���,b��@�>a�iϊ7Me���'�^Bc����ڐ�O�{"J0��O���@!�!���&�)Q#��`$D�O�Q#��߁*��PH�.B�9���V�<�*O���s����e�3c��xR�e
_�,�3�s���4W�n��'~�6�<�i>�0ī��Ti���c�qk4A!�r�XAݴRP���'�R�2��/��$��e�Щ�Ү�v��4��HR�u�v�P��<!�>����1��]�ĉJ�37���i�2����[����2@65�nQ�a��-�<+v�J)���6��6Vǔ1`�E�\�BTA�e#Xo�=�5�hD�j��A"q�"4_�H��٨��#F�mQ�(#���K&J	o��:`�P���	���;m>��P�N���"��
��	��ms' O{��hz�W������G'�� �:�V��3k! 
�!�QH�=F����V�7�nA�`B�py��0�U۲h/2f�K3�y��D*d�]4m�d=p����HT,�;�y+0�i���'�"�O�@�@d��xw�٩Rq�xK���Il��oZԟ8��2e
#<�~B���/.lDN^7A �̹�[����B*�MC��?����
��x�OV&d{���}�`u0�F窜�Op��ux�ϲ<1��?��g̓��d�Y�~-0ir�*IZ����Ee���'�r�'��=: �,�4����O���@�>Z�|��˩7��}Ae�Y}��'Y�'ۥ��'sB�'>�m�e���'(Z
F�T@j"$E�X��6m�O\�S2HAJ�i>��	�'�yZ4��qnt �B���tsa#gӂ���_�1O����O��Ĺ<y� �.9��A:+Q�5��52&�-@1���d�xR�'���'��	� �	9l�����/5v�e�C�8����f/�I��I���'
�QBhf>�*pC_'J1<�+���hO�)y��>���?i�����O��$ɪ���+DԠ#��Q
�a�%�B��?���?	,O��RrJc��5ɼ�C�T��v��R@�lS��k�4�?�����OZ��B?K��� � ��
k��@D�N�:y�õi!��'剬=��H|�������@�����$�����,h�|mZYy��'|��_�����i0^�S1,�&a�LD����)��h���+[�����i���'�?��']��	#Y�H4ĦF9Ge�����u�6��O��d�E��S�t��ē9����'$U�}o��� �7;;�lZg����ߴ�?���*lZ�?�O<�'|��@a'#�8���H!94��i�:���S����؟��3�Iҟ`��H�8�,%Q(�=@�(�/��m�� �I��(��j�����|Z��?�G���\�vf�o}�@їω�'j�	��x����Hb��������}>�}H�C^�> Taq�OͲV�,trߴ�?)�eH)Xm���D�'��\�xH#i�v����dA�(�<1��n&�Mk��1r�y�<1���?i�����2?Dƀ���,V:��f�g�4�d�H�	��I��'�b�'�Xa��B53��"�����(���j����'�b�'�"S�����ćB$jaH1�w��R'`К��ä����O^���O$��?q�p�Τ�O�ޱIw�0�FQq�ϷIXX]Q�O���O�Ī<QtU)�Oh��j��\���Ž<��萒�m� ���O���?���:X��~��kŲk�N�Ð���B���bR�����oy�'a�h��R>Q�I�t�ӎe�����!�Dot�Z��R�Hy���}�'�Ġd	9����� �P+�������Mˋ)�paB_���	�Q9@��I֟���ʟ@�SYyZw��� &Rtݔi�a�?I<ZȊ�Oh�D�2�&���F+��t��W2N������;O�օ�)b�'���'�$P�����a�I>XH�%�	D6��C�M#%
�n^��<E���'���I��^\�p9Q��+pC
9X�~����O&��@�6� ��|���?�'�^4ɰm���<Y�ڰ8�p�k�:��s��8�O|����?��'���"�/� .����ԝd�\(��4�?9BZ���d�O`���O����XT��Zf
�>�μ[��>17�ɥ,���'�'E���4*b�%t(�[�[�P���ce�g�T�'�"�'=R���O29c ��(��t�3�;/���AS-I�]�Du������Iß�'y�&�mH�)��B͘�J� ��Z�^Q�QK_3X����'�B�'(�O���Z5�� 1��i��9+aBL�D��W��W(D��Or�d�ODʓ�?���N����O��8 g	J$�9��T0'�֦!��7M�O㟬�I�l�$m�.#�$��x��Iy΀Hۚ�RcDI�2؛�'	��ڟ��$-|���'l��O�=�Պ�e���#�3JN�Cfc.��Ry"e��O�. ����T�K?������>z����`�1"]��x�I`�	�?Q��u��X�:_�Ty4i�1I��ѫ�������<Y���j��ħQHI�*�5aR ��G¤/m��o��JJ��	��l����8��Yy�O��Bʑ$�� �U�g��]�U@�/s��W��Dx����'�������6@�J8��FblOe����OF�D)\o���|���?��'޶����˦-�4\�� Fm���4�IK��0H|����?��'�\u��ׇn��(�Ė)M�9ߴ�?�R����$�O8�D�O�� @�%"�(d*S;N4A���>��j��,f$��'��'k�I�(03�"hF�
>7��k7�; 6��'���'�b���O�X�J�=t��x��m
����j�-Ī ����<�Iҟ��'RBd�8Qz�	R�5��(�f!G�$���7n?��&�'���'��OR�ĉ�Z��y��i�th"��D� �L:f�>�p�O\���O���?���D�����O>4��H�!V�2�9"�1!��ꦙ��N���?y��lva$�|C�*o���G�E\�(��.f����<	��x�*�����OD�	
���� �k�f0[f�� f��>1��Gt���gH|�S�dH@-@� �
n�b$z��vDѭ����O��:"+�O���Oj�d���Ӻ��I�>Jm ��.�($����H}B�'��ڶ�Ʃ����O� u� �Z�(�Ѡ!�%k�p��4+ja���?	���?�����4�:�d�j,�P5��e0� J�L�Y��lڞ1e�iZE�9�)§�?���8M�����L?���2����M����'?��'�x���X��Sl��f?�b�  4�zFB
�?����!�ĊR	1O��Uu��ߟ���f?���JT�2W)H22r$oԟ��VHTy��'W��'@qOn`臫O'4���j�&ȨT��H�`V��q�I����?������O��rh�G �,t~q2Vc�)���H�<���?���'b���:Wj�a6 ��t�&���E��h��Й�Jɦ��$�O��Ľ<�����y�O_�Yo�5eA�-��Y�n8�ش�?���?ً��'W꼘�(�M�a�*EP{3�WuȀ�C)�~}b�'��R���	�+���Oh�N����I���6QID��M�W�7m�O����<I�Tْ��$�Ė�.��� F͉\b�e���@>Z՛��'���ݟR�W��'��OM�a�r��M�^�k+�&�jX��.���dRb$�|��b��U9
�z��S�L($�ȇ>l���'�����Bq2�'��']�V���Iu�Ԛ�U�<&(�� cb�8eT���ɞ�4c_&1O��
��a��?A�
���Ӣ1�@;�i,U�g�'<��'"��O��i>���k��*�Ō�H�b�F.KXq��4f��])��s�S�O�¯X�y�6����5��l��#ݨ</�7��O2���O�Dfǧ<�'�?���~�-YWfYQ4G�
(��	J!lb��3$E���ħ�?���~�$ͧUH&����n �9+w/���M��S���/ON���O���=��94~��1�'j��Z�|s��'O�A��W~��'g�X���	�c֎s��U� �h��a�o�MV�ty"�'3"�'��Of�D`�0��,�b] �0��ت���|2����@��ty�'� ���ן�������h�� �����S���9'�i>b�'�r���O��C?]��.�+�9���_�P:I�% 	7��D�O��D�<Y�uߔ��,���ĉܰ�k˞`#�ů*PQ<�lZ�,�?���CM���#�@�I�kd2ts1�Q5���ab-�/�N6�O�˓�?������)�O������d� +�<S�0@q6t�X�$^a쓻?yB�Q87���<�O�$ᲂ�=R�4�v�̎9���O��D�&Zi �$�Ob��O��)�<��`�"`\�U%>�
�a��C^��'���?5�`�y����^�hs*�P��U����0�-�M���?����?���
+O��O�EcflB�{�q�L)	��<x�q2ǘ5Y��y�9�)�'�?)�� �A#�"i�l���[\����i��'e2�.1��i>���䟈�7����f(� E��mP���P�>v��$>��	���I�\y��!���F{d�a�y��ݫ�4�?Q�C�G����'R�'���~��'~J}�#!�w)z�����]g�tb�O�4IR3O����OJ���O2�'�?�Ƅȏ �=�'�J�`�GC6H< �#�������@�I��������?�2#<�"Q�Ơ%K��FՊvn4�ϓ�?Q���?����?!-�|pJF�@ۦH4kX�3�y�t���T��ܫa�܇�M����?q���?������O,\zU>�k��2:�0ad��o*H- bK����ߟ��I۟��	ٟ��΍�M��?a�aC�O
�C�+w�*��q��++���'���'�����(�o�{yr�O���3Δ 1����OO�ȄA�7�iE��'��'}h@��	|���D�O��$��Ȍ+�M\�hk�H]1�\1��妍��ly"�'�N�O�ɧ�ܴia[�j��Z��H�K	�m����	
f�kڴ�?���?��'�R�2�,���-$ݢi��L��8a�W�$�I�o�:�����h������t@�:�b+PF2E\u���ݦ]
u!��M����?y�������?���?QaōV<���J�w��X���0m����6S��'��i>M%?��I>_�Ehfi��!�tڡMaȽ�ݴ�?��?��F����F�'���':r�uw� rk���.M-�)	�I�3�M#L>�Q�]�<�O��'����t̰��$�d��ˌ@Y07-�O��xp�E���	�����������IF$�,���W�}��� G-l4
�&�� ��?����?����?i���?�dɀ�zd���G&J��iR�a
>Gj�T���i�"�'#��'�������Oް�n�v�؝3a嘢��dX�!ۖT��Ľ<����?1���?1��y�E���i2��9�eج]$��k0Û8��*F#d�R���O��d�Oj�Ī<���9Lx%�'*��ܻ �R�9� �*�Q]��\�лib�'�2�'��T�T5�H|�1�.x���B54����Ƀv~�Pn�ݟ$� ��ݟ����*�ɯ;�+"'6iH�`�JE6	�@6��OF��<�U��|��O���O�ų&"M�y�`�'f��Q"�{��"�d�O$��[-0�F��/�T?�+ƕJ	��(T�q��z��`���V���s�i��'�?�'K���6!إ!N �.,s��$nw�7��O6�$���$.��)�*�҄���[2~/�kt#ԗfכƧ�W~7��O�d�O`�Io�	�DAj���*(#d�a;�DH L]��M6������(��Ǐ8b�r�M�@.��B���Uo�韬�	�0��'U	���?i���~2'�,��B6B���"$ZCg؏�M�H>y�C�<�OO�'�K�^��k'm�.#s�5�I�r_@7��O<�ʖdQx�I����f�i�ř�L�<��ʂ�$i4�Sdj�>ѣN���?�)O��$�O����, �gM3^G��`q,
�2A�H�T�U.s&9'�h�	�&�l�I����R�Bi5�ӫ!Ô�P2�X ��IPy��'�"�'@�I�1�O�:`
�o�-{�B�@��@�H�'���'2�'���'�v�˙'�����R�HXaB�-r|�ҍ�>���?!���dHCH]$>�t!��
���Y4s�t�ʡ��4�Ms����?y��Ed�L���I67p�m���"��͠G@ҿ��6��OP���<��cWLډO�O`�]X��SG��+��Wt�� �5�'�D�O��Dצ8��1�T?��"�0x����r�Q�@Ҕ�`�F�6Q�ZE�i��'�?��)g�Ic��$�3q�1��L�C��7��O&�$�ϖ�D4����o�i�������3mW�~}�F��
"z7��O����Op�I�o�l��XA�F	�wM�aR��=��k3�i���*�'K�')�SSy��'��J���Q,�e���Y�12��Dmӌ���Ox��:!�`�%���	�����P%Dɪ"�Q=OG�]��l	%>�mZi�I�i��pK|����?��Q�LKE̋�tL�S ϒ��z��s�i�R�W�s��OP���OēOkLG�9~`p{��F�h��q"�bJ�I��LA�IRyR4�"�'H�ɥp��[2��a�����X,(�A�4��ē�?����O�8s���Jqaz�ē7~K ���Ӭt���$�<���?����",���ΧvЀB�"4a� ,#W���~���'��	ԟ쉆�Aş� u@�b��]��øV�Z\�#Ө����O`���<)�M��M/�P��I�M(�ȡ�e��=���1$al@n�ϟ &����ϟ�(�h�8H�O�� "n۳_L|�2(��M���T�iR�'Y�ɐf�
O|j����"�A>s���傫]N�C��"}u�'���'�*���T?}#�E�m�VT33L׳3�,@�1kӆ�	<Z��S�iɰ�'�?�ƺ+d����3��=���S�LQ+K�8ӗ�g����OH4w�)��7��ȵ�9L�܄���gv:6�*��Lm韴�	ܟ��&�ē�?Y����Fތ�sDOƲBt����Ac��a^;�O>���7o�6���Nϝ=��т�A��XY�ߴ�?���?	%M�(7��'y�'~���pNl���67EH��QkI�O�O�]�W�$�O����O����ɋ0]��x;S�ߌO0<�ҩ���U�	�14��IƟ\��:��?��0YL�检J�>� �ʘLM�%�'ֹҏy��'��'U�'=�� V9逩�I��U�b�XL�pzrY���$�<q�����?y�D�BT�cGK-�N)���35z�����E�J��'	"�'��U��0�m���dD�<|���2&��!/](������D�O����On㟨�~��..��e*'�͐����0��t}2�'t"�'���'����'�2�'|p�a�#S�4ѐ�hx�}rLk����8�$�O�����(~L���x�M��#Q ^m��(V�0�M����?)O�l�Վ�G�˟���A0�[�'D�;�T�a�Ʉ�HaȼbI<y���?Y!f�H���	K�^,��� �K�=��q�+a��[�|ka	��M37P?}���?���O� Yc��yP���De��@���F�ij"�'�����i�@��\�c\n@t��O_�VB ,�t6M�O����OB�IEN��� K�dmP�+&凃��A�F�S	�M+ǀ�W��������&t�b��oj8�5M��-�tlZ蟰��ǟ8�C�0�ē�?y��~��Il�i1��5@.u{!����'e�X:�yr�'{"�'&q�Ҡ�F��lG���F�|����*,f %�0�	ן�$�֘���!�#U*B�j���J���M
���<���?���DN�$�f0 �`�Ь�AT�_!9�ڈY�j�C�I��0��v�	��4��-5���i&N���lpY>�TQ��f/�I��,�	ן��'�N�+�ko>�q�`����iG�Zs�$Ұ��>a��?K>i���?y�W}RG��i���Q!�(�pbʝ0����Ov��O����OfZ�|2�'�YĬJa�"��oG�
���۴�?�J>q���$ɇ ĉ'j6�H�	�;t-`��m��T!�E��4�?)���DN��)&>����?�H� ܀L�.Q�jF�Z<!�����M�r挋∟���8�~XɱmU6yt�hT��M���?aCC��?9��?����+OkĊA�)W�N#-������Wț&�'����"*�*Ţ�y��4�_R�����U�5�ڄ���0�M��盞	ӛ��' 2�'=��:�$�O��B��&''T�Ѷ>v0�q���}��"#�S�O�I�$
��sE��ޞmw\nK�7��O����O��X0mw�������h?�����V��̣�(,i�T�7Mp�/���<	��?9��k
n�Y�ʟ�=��*��E0�Pif�ih��;Q��O����O�Ok̏#o>xEK��h����恂4i�I�]	�b���ß �	vy"�V/\  �wc�6�<=yũ̈h��}��m2���OD�9���OF�D�.��U읽5rFL�>>2�I˖���O��$�O�˓#<�=���'݇ �\�j���'�H���^��	ӟp$��Iӟ$z�.�>� ѥ"�����_{�(� 5^}��'�r�'a��'�e��_>����K�ҠQ��&��r��� ���Zڴ�?aI>���?)S�C�=��1�)-<v��d`��z<1@���?���#�Ѥyv\XrD	p`T�O��.F���(;�:�̻}�����^sVZ��kX�D4&؅ȓ>m��jig� S���3M�b��FO)U�ԙ�F��"��uK��5u���ȟ�G��K�mZ�^�2�DJ#Y����֚bF���Re�"$~�l�毄=s��]�%c�9�#�Fσ~�r�ӗɛ�V~��`�4V�̰g��� N���/
�J1޺ZQ�|@��&'$�,s��7�UZ��.�Xz��?����?��]@�˂�8��ĩL�4�M�3��=��(�@&�~��
�hԤ/�c>93H�T��U*Rɬar��.N�0�B��O<}���j�E,:1�E� 5���r��ٶ��i�1:Ԑԋ�w<B ��dݹ���Z�l��/���Sw
$����/���L>9q ��.���S��[ �J� K�<��n�-�t�E��&)D�]r�I�<!�!+����T�	�VW�ĂAA��m�� %�R��Q��N�!zH�L����`�	���Yw���'x��!7�P5���͖("�a#Ì�M�R�"�8)�����6\���#�ir��\�n�.Y8 �[M�Z�qH='� ł�)ߝ�t��<'�>�#��z��wG��ҕP+������I1}�6q�����"�
!�Q�(��B�&�L4�:l �qP��.Bތb�,��4�� �F�qW?�	&f���*R퐓-�쵱��eވ���韈��lߟ��	�|��k�J��I��M4U�Z�Z�4Y�P����[s���'EO�SU�8���}ļq�m-���pp�[�s�J����ۂx����&O.O��'9Q���0�}��e� &���A��W̓��=��*��{���bȂ�C4�,���O<A0�i�v<��E�b*N��d�U��<YK��'C�I�7a*��ܴ�?1���	�E$���h6���E\����w��mD���O�yÒo/LA8��،CW��� �=���S>�9恏�8r��0 ңZ�l]�և!}��u�vA�����t��A�+*���]0^��m2Ю;g�����#Z�:L�ʦ&#��O�e�P�'�1O�v$��A�2r��d�ǀU?z.��d"O�@�"I�H[l�cƈ�A^%q��(��|���	�%���;!�(3G�$��� &���[޴�?���?�(Z/N�:y���?I��?�;3:�ȅ������4N�H�B �Wn�"U���'j����IY�����S�? ��ٖi�=u�n
��1\A���pE��}�<\2t)���P�VC�#>wq��'L�� @�Y9T5 $�E.פ(� D1��'���/HQ��4��=	1�݆k=xd�Q-� ^�)��mp�<tO��X!�����RP4�� i~�(��|"����J��āHt�rX���EÕ���'��j*.�d�OR�D�Oԅ�;�?	�����'�
<�FD��dҌJ�1QJ4��n�;^"d]C5�(S¤qP��*����
�.�P�����5�m��Ȧw�F�q /� k�.88E�/*^n�{��Z>�qOޭ[�@�6[+he�&�G�Mg��	��*	�6�O�`Q��% %�x��큾0V�ip�"O`P���D�ȵP��]�-G��X��D���m'�� �����)�O�	`Aϴn@f��jK\=���BJ�O��䖳g�����OT� _2��5(�L{>�alI�6���BAL:�tPJU� C6�<��'Z.����X)xfL��У��Z�zPpd���hG�÷j�3or��5cO]8� !w,�O��m�$���T9r�%0����lɚ(�=	t1O@��2<O����يl�$@���X�r΢�cAO�l�n���$&�B��4���n,�	eyRlV�B�R6-�O����|��NF�?i�g¨;�60���"�`!J��ρ�?���I�2�ٴm`�iX3�ϟA_V���ZdB(����Q�!L�}qp�\�C' ݸ�#}�U��ME�ǹ>��yP�aTH,�Ԫ�w7N�Six�1�ċ�Ϻ�d�ڹ[�)���"}�I���?�E�|���m	�&��]c�˘�i�)3g���y�e�(��}����g��$*5@��0<1 �ɢcό��G�҈ Z����b����şp�	a8�0iY���������i�abc�cW�h����y&�����?&����u�@�.E�����M���|�M�!�fec��!�.	0D@�m�����Z>���j��6'䚌��%}ҦʶI}<с�_4 �rp3֬�Ki��O|`3������0%�c�5�.�`c㑱���kl�ᄤ��1�Y`%��a�m�'؜#=ͧ��L�g��)t�4x���vr��@����wW��*���?Q��?Yw������OT�����&$ǟb����iU�\q����M�Xb�d(��#h���F��V�'�AP�Ϛ!D�J��v��,f4x��í��"�t�:���^وH�ĥ�7�џL�e�8|Pb��
n���;�k�.tH���`ٴ��''Xb?qa�/@�]�$����++�y#�;D�T	�+�˾�0�ͺ@�L��;�	�M�����
:<�mZ쟤���̝Q��u�ԨB4�M��<����qA�L蟸���|"�,�j<[�ђt��I�'�!y"̆�RtXLP&U��A��Ǽ=rP����v�P�e��.$��W�D;��MҳbSo�zP{����qAB*?�$G�?�|�+s�Ώi����A� K�!�d�(u���� +�d9K����!���ڦ���� J��$yک�F��BX�=m\����4�?�����I�>o����&#�*a��.ʀ�b ��7^^���OP�c�T�/Z�"��>�Oe�:�Q������	Ri��T���'L^�2� V���%{!����J�E�$D�y{�m!W�ɨj$���$*���	�S�@��`�)�Se�Ӓ����E#7����C䉦Od:��k��?�p%�g̦Hv���Gc�'������MCtc�%Ȩ0�T�y�
y�J��O���yO*1覉�O����On�4�\�{����hȩ��j�F� �A�},��'Kv�:R��������b4k�^����*N�W㔽R𫎶t��:1��+���|b�l32h`bd*E ��aj�3P}��O��!������V�K�HX�t9L�R�Rx�J9�ȓ.ڼdx
4tptz #=P�$UΓ�?���i>9$��3�!����ϑ�N�Ձ�n�310��/�����	џ��	��u��'�B2�^I3BSB��eF��Q��(�s�.FW�8�E>ha|ra�;-R�i��з&�-�v�\<3|��rCT�	���bQ�]�*%��e�6��Oj��Q���Yݬ< ���4�=��$� QC2�j�Θm�4�'�����E��t۳L#-k�#E�J�o�!�Dĥad`�Ѝ��~d� ���Ǳ
�1O�����OR˓`�]���n�$�O��(͍]����L�3_�q����O��D�>��D�O�S�d��mI�˨op~�d>)`�Y�7�2ӆ5a;��㉴_��!�F��N�h%�}c��f�>=�P���4Ҫ�00��#k
uF{�	��?a%�i%d�^긨@CS)�p�F��	/B�y��?Q����������+X4ܑ��^3"N<SfO(�l6�FI�GA�k��+�n� ca�d��Dy��f��7m�</�,�F�O��RN�W�,��
�U���B%�O4��	.=f�8�/�=hEc��^W�N���O�S�Kh�k�/�7d� {""^l�'��� ��I�sF��a`���EJ��u*�Q�@@�/�� L��E�}.mg��5(��ß>�t�D���+H>�����X�F�zajԈ%��# �NS�<1D%|KM��FI.�˥�FH�����͙b�|<�g�0R����&Ҙm͟�����(B�G�Q�>��I�$����$f�� PEɽ^.���< �f�Å獙0<L����i?�]R�[d�g�!K��Ep	ǎ��a	D`�6�N��5�1�����Q
��* 	95/���'�ur��U5X�%#P�H1��Pf9�DH0���L>9 �=7b�U��̑D������C�<�i�#X&���E�]�r�B��X|~d-��|"O>	2�O�X�L�îVꎸ�F�$viP�������O����OZd�;�?1������Xi�L"ag�LDݐ@ �t�����Ǿ&�Ʌ�(��{���\��$G�2�A�E��?S��q3S�X�(r�@��2O������n�xA�L�Z�\�C�ƍ�R�'�*�;�1c�uX��Y!Eh�A��'�����Y�1��`��HG(f�$؎yR�x��O��H����I��d@)N9;I�T�תG�?<�Ia�ҟ��I�`(�	֟�̧&>4���ʪUJ�`v#�7�:܃��N�.�Ц/
~֖�Tc�'_v��h˵��J�����(1"�I�s*T�Tb�P�Q3'��c��59@�A��4pR�A�����sV�Q����ē|��-BG��e�L��eC�sCڠ��`u�P7,J_��(f��b��.�hO�����能*���@��VU��G��'�8dz3'g����O,�'WNbԘ����a9���)/P����˨;���`���?�]��0�@�Ǖ&�"� ���ɮ|�v��=�� �EG��&�`��b��� wͪ� S�v�ֵ"��1 �~�IR��T�H�:a�_����'��R���?9��?K~���`ȭ��-�Z‥�i?R���i��?��?��@|\ٓuLJhf�9�b� ����I�HO�y���f7��Z��E$0�@�	�QئI�	��I����*5������ӟ��"�u'C�&�`��6�A9&�Uy���`\��J���1m��\�!��1M�y4�)��9�H�'�s7��<�d����]$����̵Q�5(���%�}�5`O���O��\�#�[�<a%���Y���z �;��Qd�K�Y��'��Q+�S�g�	�fJ^D��C��hŠ2
Kh�BB�b:n�-��mF�X��#�<K��0$����E�ɗ� <G��Xx��޵���	G.X%��ԟD���_wB��'��	�<*¸ȥ�${@�j3�%�p}3f�	w+(����:|O6,c�����/�=
 ���m;�xX�f��f��4XӣԝՒUe%�,ʳ��k��!b���EZ&ȻR��㟤���22��yu����s��ޯ")dC䉃t�X�0k^�*�F��[1E]6c��I�}�'5\y�7��O��D�3�xK�i`y>�;�-̹ �����Od�D��O��Dd>e2BoL�y����k�!4�D�lګm!x�w&�3A�ތ�.�"3h���R�eP�!l�pp�UPQPF�<.�u����!�61Ⲧ�3�=it�����I<���M�>�S��Ë�0�H�S�<�&�&�@�F2v����RQ<r�i� �2����P%М�F��y�@�-�D��?	,�n��d�O�Y(�,V�C
l�c)�/��q7��O���"
�� �A-� g,ח�_�ܠs�ν>E`h�+��(itE^!�S�E7�P�pa�>�f��X`L���B��|p҃�:u�l�5=J���l��N2���	�x��M�"e��'!�>��I�/0(ۅ�� m'h,+ҩˉ(�d|�Ɠ�f�[r�4� ��Ҝ(��x��ɏ�HOv�Puf�łk˧5��t�XM7f�l���П�s�B��G����͟������YwvX��հf�L	���K6'��[�扎^ޱ��&�!�L/u1��'j��	GK�&�$�C�P�)�����FB����"MƧ0 PIK�Ʒ[TD$>1������.�3��1j�2���"TC�@�ul���M3��e�
�(�S�gy�'�@y�O�B���P(0>naH�O���"�үu�޴�q�Xl���Ô�@���$N;�~2T�8��Ȅ3�B�ڰiޡYřV�H����������̟��ɖ�u��'�25���1+�^�*��`�j 2Lp/X:�2���(�pdv��%����p<�����h�lݪ!Ɯh�	!���>�
���ڥ0"����(�ư�@ΞV�'֔A[���/	��,��(�#|��� T��?٥�'ov�J f��J�t�)Ƀ\�ȡ
�'L.v%��ƅiܚ�B#�D�b�$��}���;C,7��O����8���KL=JE�-d8����O��#��O\��w>��Ŋ ?U�� 癶T8�E�B���l!�u��Z�)ھD��x��D�� V7X��A[1�V��"�#����@:��}I�����"C
�d�|�)� ��Tl�7_�.�%h	bO^��"O��!խ@"=�$4!sGˌ\FF��OnZ�5V�%��a�4.�<�GgG�&1*c�R�M����?�/�Z j���Od@�;z��`���V�P��5e�O����7��Ej��:@r��ig�'�M�O��+A���g�-��e�7�+2y�'W�Q�!��`�LI�nQ/�|BRhYF���xt醢y�VM9�z��E��/(���̡V��<DțX~��r�$��F�!�$C�?AM0��*Z>��1��N!ax"�=�c�)����i��oW h�!�iRR�'�k��4L�:6�'	�'��wJNH�҂0kX��8��{ELEj���̓M!L��Ó�Ե����3wm ��&F�V��=A�%U2�6���E4ʉ��g�";TѠ�b��b�̀���Oq��'?F� �D����@+R�N�i�'�pԺ�CN�K�\hU)�/ n&���O�DEz��I]0J�ڠ�1�3q�$��sL�	���j�ַ/~.�$�O��$�OȤ���?!�����.����M�$�(А���0-J��	E#�t|)A���>����d2�,ؙ�e�y�`�1��!8=�0(�:�9�,Ybqx͇剜�M�D�'P}���q�T,F2�+�m�՟�3�4�?A��?����?����?Q.��t���Ͱd���0f):Zr�y�"O��ғ���:F�k��$8�v/l1O���'��I`��Is�4�?��7X�h��Dlj�b�ҭb���?����%�?q���d�*
$�Bt�SS� cCa�t6�8����qEE"���D{ў�H&hNs�A�W��r��0�p��f��0��͡B��Djb���.���z�'�N�[���ow@@�h7Oʒ��n�;�~,�ȓ
��-q�#�(�� Ɂ����`��ud�f`Կ-Δ�#Č	ʖ���ώ��'�De	��o���O�ʧn��@`��`\^\д�I�n���s�d�:w��hX��?iVn%%L�0z֪��\;��іbD����|r��RD;$�@0�7V�L�ô%JA��� X��%)�C2�X�˃*O�#|��l
�&ɅU������_{��YCS�>ɑ������N>��2(�R��X�VbLQ�0A���<�Q��u�� �ckN=���WE[U�TX���ɳ%^�Z���rp�L��G(f�8oZ�����ӟ���E� �Iß���ߟ��/H�A�$� -vx��@��q�`Cဒ�|�ą���i���p0��ߘ��M����s�B%L(�Э_9T��WmQ�n��}�|�۶-������rc��jB�3���[�β��,� �|β�?�}&�P�F�Ƽ\�.���H�>�D��j,D�Ȼ�#�&�lg�����{D�+?!��)§tL�m�vdO:a[�  �)��ٰ�I�w�N���?I��?�f���D�O���Zznm��㌎7x9�e�I�=n^�x�b�jpyR��nVD�y�.�������Y�"�s�����T{��M&kD����[&`���j��'р +�2Z�l��j�9I�&D��A���?i%�'�V�22
Z��y��\A#�l3�'�(ec2G��b � +��=�HaY�y2�6�I�.�<-�ݴ�?��U@\j �Z)0�HR��G�ٻ���?����7�?!����TgW2Ob�#1�ކr���	�%Ш����N �TA�iɼf���ϔ�,�R�g,���n�4H��8B���܋%z̈́�ə4n���-��]�C�	�m��S�#ǌ�-3v!�$ܧ~�^mR��57:ՠ"�ѓdt!��ئY���J�*�'��$�NQ)4�.�	�a��q!ܴ�?1���	�y��dG�:�AV��.=�LAx��5X2���O���pI� �
r�c=?�O%�$?���v ��O���KA`F���'�Vu�bM�$@ܽ��

b�ܔE�D!H- ��u�3�݁i
��(��ӭ�����g�)���Sj]�W!��D���P��Q�<C�I�O`�T(ƥ��t~�ӡ"R��2��D�N�'��ecsCąZ�� g3�&px�|�x��O��䉙���(��O���O��4�|$ȅM����'dS�H�`�ab	�o��	�fQ9��O�g�I�	�QrP�ҾG�0�ywY.w x����V<��i�G�f)�usb:�*$��	�Y
ʍ�)͸y���#�*>L��M>�c�џ�>�O�h�7K��Z���mW�D���"O��c�Q�+.Z��-�-j��Xb��H���ᓳc1
����5
f���* s�sSA49lbD������	����]w��'��)�yn���
�"�ťTa9����bZ�[����oN�b.�ل�	�]��J6��G�����@ rm�5j�<gp��B�*�$�3��yӊ�2d���t��<	$��tnp)an@���1��螸T�`�� ��?� ryJс�?��p�̊�$	���"O��wg��x~�sk�8u]���]G�Gʚ�"Ǳi�R�'��B�E��p�$ђD�P�r�����'Ib�
�O�"�'��^�F�p�ǏB�.,���H�Bq<X�D@�9jϾ+񬇟h��r�-��*�p���H�|�s&΍��ҭ2t�!"|���@�!l�t���eݰqE���$Jt�'7�D��ى'ؖ�qi�4��q�7��(E��c�'�lu0�$�eVf,���	�;�F���'c�6�ۣ���H��ȠLƺ���E�!�L3+���;w�/f`l0��|�!�D.�P<�M]3a?��b ��(�!�G?wv���+������L�!�$5%*��2㇜y.��۶nɛ~�!��^/Q\���7c"<��-��Ai!��&=(���k��v�x1;S�[f�!�dI#@��5z�O��	��I���|�!�d�1��t1"�Ĵ�Х"�^'Q�!�$W*!�L��lD�3�R-@ �ń?�!�d���躤`�~+�E{���4�!�$ܐ)pHu:�
�6O�ysGa)V�!��+n-n4��Ö!��� ���!���+{���:q#�M�Bu���_*�!�Dھ^�Ԍ1'�ۍ$~��h�O��C�!�D��$�6�B��W��I�B[*�!�dJ�$�L��ĥ$�4pҦ�ծ)�!�ϯN�h\�2��'�4��4@�:p�!��1�f�r�L�w�4l��i�4D7!�D׼5 �@���ǒ�<�0Hه�!�$��k�T-:��l��mP3��-:�!�ΝtTX�z2�0��]�ݧ�!�_�*u��)&� 8z(�W�)Q�!�d�<�3�(9z4(tR�#L<$!��4(�T����|����"�!��N6�� �ꀨ>�(̘� J��!�ݛR�\@ hS�]��x��N�"!��6�r�#��l���&$l!��>V��1�ϠdHS%�~e!�̩N�3ר�!h��4�WIV7c!�2bE����t����Ê��.=!��W�H�`��֮��@�~�`6J4V!�r����6��%����a	��!�d��lB��7��*�Bez���!=>!�F:!�tA�N �DU�Q��5*!�.N���+�Y��yjv␑8�!�d��Z�I�����@h���b��x"͇�g�����&��	`cu�!l�@�.-�D��,C�I�qFҙ�đ.] ��$\rt��:�Y�dd��2�8�'?ˀSf���qS,X�"4��ȓ��ز�M&1Q	�a�����Ø{Y���,k� ��4�4�3�I$�d��C�" =����L��?& C�I0d$da�d��e�.L�5'���i+��0&�f�Zr����|b���z���sfjƠ|�~��%��<�0<A����s�QN��	<�P��¯n��IPL:bB䉬We.LC  w���JÂB�$�F��]c֩��AH��<�:���������%�ԫ)H`aDy��z-�����AL��!��K�D��z�B�:��I�S6�I�0,@�C
���!�M?�G��%��<�|�<�� Bd�Dɥkأ	
v՚wX�L�"%BrY�:�<��hG�9�dȌ�i�L�f��j�3fnɱ�G�L��dǺ[ ��2��D���je03�@�``��J�߇}�I�ƀ@h�[�'x>=�EF�ZD+�
p�z$ͧ:�4@#�П���<c,��/��`5�4� H+G5�ha��9F5ZR�OgAj9kV	 ?y�f\�SX�����U
����.^�G��48����,~\���fP�-`�D���d���o�'����@��>
��#Q�Q�x� xv!��Ot�9���R��� g�c�ȹć�a?�s���'ۦ!�J��C  ���%(�.(��t� �$ ߪ�)ˆaQ�\� �Z�b����;E�*��W�ѕL��$i�`���������)X�CK|D�OvJ=̧z�Xq�j@�C�
�yFu����q)�/
�>���;Q�VT�'�E�? 0��%�)|P�.A)B5�*���,� N\�V�z<��>�����hL�\Y7lR)
���B�^��=Ex��@�gX��6fɆ��pE�ܝJ�T9�'��5�p�+t�I `խ3 L��]�G����r��O���&HЊ�fA�fD�"��=0��ۄ�r�R5� #�P�����#�l��'V�|0F��k��r`�i>E���;����[�@ �y�l�>��pӼ�
 ���^A�E���$�HO ���`��&��p�Q�7�8����X��I(��i>	P��סg\-p�Oe�E"�D̮�R��&ĝ���@�p=���Y'5onYy	�����4����C:�N��'a����[�p<��jW�'}��Jax�yѦ��0`ڄ���*���SO�d��g�I�cs�K��<�D��� �6kHV$x��q�x�'� Lb�4��A�_$NT��ɜ�ew��H����σKK����iP���g>H�'⤔Rr@V
`��U��,ǷE�V��'FZ	e�t�B2gLNr}YPc?j����4��(:7h��4���3瘿(V���G��3ƸH'�Q�y���f-�*�p<��h҉ �:�bNܚ9�t�ش�Ժ	&�J�k���D
��1{Nɀ�i�>���x�P��`��Me���ÉK�Y���dC9(-�Q�Vo�%3�f�3a	��t�٢F�� @�A`����ō�"��@B<��?E"��DJ̌3�,����|���:��S>X�3uN+� &�h;�/�yq$l�q"�<0� @���<Q��D r����$,x�@*G9qD\t��8$c��'�ʈ!� yt����	�m�u����g�-����P �ծIJ )z�`�2zM�Q�0��?�13|@�r碖�f;��g`J%'�7�(n\�P�d��@|M��4O�39
��hk LA�qB���Vf�S�Q��	ٲ�M+��HN�z��@Cߨ,�tL)nn��p�'�2�W�K���;��Y����"�(�q^��f'��~b�)�`��f�&�T?��{�I�äK,1�b��$��v�1�v$��:5Gxr�A�&��`WAI��aa��X����`�4uCǥH\㮘���T<G��!�ACן��1暉��4܊�?e���;�Bd����%=lF�@`K[(<�5"T6[<�\��nT*��#<��kPL�;]	4	� YQ�HE
wE�W�I0ZHDs�'�\���1����$m��ґI�'�~qT��R�h%&�t�Q���ՙ@��1r5��0($9G�Q�b,�Q&�'��*�J�9%��0p�A���V���NǊh<^���C�.(��YH�fŸ�ا��-�SPD�S���*5�8��Q�;^�#<�s��Z ��9�b����s"������8A$-;WIQ=qk�aY#���R��ə

�Y��ӯ��"sc&Q�\�Q�`]�(5$�r��pb-ܥYE�1�m�O�O���bÅ$�fu8�	i}V@�d)�M���ɌG@4'��*(8�-"A��f�'�����aO�<��珂SEb����>�U��S)��):Q,F,�0|:�
��2m�%BYH)X�H�s����e�>Od#�h�Y��L1q~,�w܄h}N�ht�ߜY����q�L������̛A�~֧���j�.lȓ	K�b� l���=ExR꒘gZ���)_l����R̕�O����@坼:b�ܠF��:���
;I��ȩO>�ɟ��E���te9�'6��˓(D+�d���B]�<�6%�`늛|	B���A�(l�ԄɇeC"O����O*n��Q�T�k�Ѱ�ݏf����^�N��2h-+0��jaO��n�D}��^.� q��b��e�.9jgk��a��䀥���X炃66�(�h�
���Z�sRL��%�M�dD��K2�)���9�v����'��ST �~��Y�ԇ 1|ʠ���R����~� ��W�m"����~���A�*�I�O�x1�@l�W�'����f+�;HHT*��F�`�Y>����հv�V��Wc-d��ǨvӼ���Jyb(�����>��@2V>7�!
�|����<`\�0����b�,��Ç�	���-39{��"��2�Ӻ�Ӻ��eŢ�T��S�טz���3%ĕ<�V-�ɚ~x���ǋ�p�B]˯����˅��ii6=�ġ[^F�䢗�,љ�nÓ��ʓ�~Z�~R5��I�t����N[75�������aZ�eJ##�=��<����1!��[�8��xf!�~�����.)l�I8���N̓>Z���i�T���̸v��������	I��:l�!�D�z�6��t�PcI|�ʊ%
�t��=	a��Љ��M�+I�+h��4!��hR�O/)�KL.2-��	?�(�C\r�,�b�u&�;�햽����T
�J0R��O쌊� R�
S��|Fy�h�6��$��C���̊���ē.����?r�������3?�G�%L����<c��@"�����xr�U(��D8娑@�fH�T�˹d7Z��0X� �0O҄z��$�O��O�	*j��X (R4W�$-
p���=a{⦋�%��T�7��#N�T�a�F�.� �1)�=8�M�E*6�d�'�p�'�� ��H��'�!�e���
` ���=Y��`��}rCN�P&Y҂��^۔�)��_wd��'��$���]�5i���	�f*�-�㖟�!0/(xMT��d���)rp�L�f��T1�)ߋd��=#6��g�N%h`G_5C�Jk�#�?qL?˓Aj�*L��P��Kv��J1�k
�'+0@ `'ϒ07�y3M�2{D�#�
 6r,�	�W)�C�N"+�`�� �bd����z _�]��t�'��r��!=V�3���Te*�;4�G��9�pl�(s��0JQ���~�4&�#MG�'�Q>���E�	b�8� ��'LF�RO,�	�1d��P���%Y�|�tH| �1ABq�(x���Ct�:���者tGV�W��"Y/:�CS�s�XJsl�8�8)��I<rR^��G��0@ܴ���A˒� �霹,\�	�'�-�,A2�^��C��p�ܵ�1��DΪD�(��`�+�"]��	�Pq�H����ˍ�i*n��uˍXy�D��κ�M6I��@�/��H8��[�{�$N.K���'B&(��{8�T;%h
�@�\��a6�8���5��!��	`�Q'ks�q��Bc��)�
!!�E@âR�n���Bs!�!�*%)�e �'�n�������DY�4����Pm3}��^�l��hi�?�v�3�=��dV������?�x؁�X����I�?��8�Q��8
E)u��"GR��aʠ9b�������,p (�O�x�+��k����Pp���TLuz �1[�'��B��܂/u@�S�B�0Y�A<44�-��]n��ؐ3 ��G$����d�+% ܺp���n�dA���������R��l���ɄD�ʸ �**�c�O��L	V���A@Zp���J�4��YP���d-J���<I�k.o��`B��Q�
�c'�H���Opxِ�`&���S�	%�R�ѳ��R|��x3�Vn����BD�I8��)��ۮwCz��6	�-4%T4���������L s])U�6��,s�lCie&4��fŗHpx�'�bI)7��w�>�C����
�I���y��[.d�� J㩉�	c
��a���5B��8@C�&c_���4��^F��Nؔ^�h��`�:��Oμ���N��i�R�t�eo�q.N���
�.jBh�P�D�<���]��� "�t��O>U���Z�&w�〉��%q�҂�C�m���D��U.�ץ�\�aRfP.��T��Έ�G�^5��4Z,j�-��J����n���O�1f�� l�;9�ia3�C<E�"?���H($����E����+�� I��{C�)w�)�F�.���n��7�	�U9�!�mݽ#@���5X�tЅ+V5��I�,.(,Z�`��z�
�2�D_ j�F�ԉ� �;br*!G�K4W�,c��,B�c�� u��f���L��)�燀�-;�����=�F� B��8���m�p�<9��H���O�!�mщ�ƌJ�nP�?\�t��)�YY�jTg܈l��C�N%O�� ��i���[�Ow�٫�!b��
���:~)���֬#E�QQ/C�0�ح��I��56���h��yP��2���mI+%��H�����6�Y:t��-k��Z?iY ������y�ό$�}Vf	
hB�Y�$ڥ��T��v�@aQ��dY>�zcN�,G�
 �&Nx<3��]�>�Bs,�@0��2o��w��h���S��	�!��5 P6T�j0��74�]ɧ��t �����Z5}H�� 
8����g�)I����ܰ�@Xт���J���xʚ6$��?k�%3b���(O�e��F5u�q�$	�	
1�-H�H�`UQC�	1wΒDy�O�
0�'i(�Kt�V>�%�R�\�R]y� ��t��$8A#�w4(����3a�^�W�<�2b&ԘI!pĎa�i���1`�$�;���cѵ"s��� ��Z/<�����_�� �E���x�=ky�q�VSdIp�&��hԸ	�D�O�GGZ�a1M&�I��e��
A(����ȱ�. �kЃ,�9)l5 �|yBJ�`�䥲�Txs��	���f�=����GhY:���*�(D �FE\}2�'_�TcA)�w����M�t�Q�����ʀ~ʐQ���ӌV_��3*!�OF$2wiɵ|���@P�Ԗ+�heJQ%��wt
�˃�Y,D�Nl��&�O�yU�֣A��_��P�^���O��x0 ��A,���JI��i.*�^��@�ڱ%�f:Ъ��!��q�����Z�n&Ě�	2sk!��.t��; X%l` Lg(�],!�ҥB�z%��-SlIrI��#$,!��~�e��j.`@�Г!���K�e�`�#A���p�S
�!���&X��P���ٗ�
ɚ3E3�!��Q8��(eO5P��AhR�&^!�R��� ϋtPD$3ՍU�=J!�$�=p:��R��n�+��`��
�'�\B�S�"f��!�`�	��h�'L���l�y*Z(�3�%�ԙ
�'.L�����FUqC�-7"1��'�n�q�)U�Qh>t�1�ь�hT[�'�lp+�
l<�u�!N�'}�X}X�'Ҽ�ŬGH��A�P�]����'ZuI`ߨT�6���/�^b�5C�'�h��Z�,�ddY��Y��Ȩ	�'F��%�D�6��a��T�{x�U��'8p�J�/�$6���5�D�cija��'h�"`_�=�$���W���
�'��D)Wȃ&T�~PƖ���	��� ��x�F�Wy*�y��	v�����"OZ|[1��6rtv����
O��9�S"O��h��ob�!;ՍO�|�4��"O4�gD�M�|ժ�>/a^�v"O�)�Q��D��q��ԅ-�L@#�"O�mh�B�8#>4+��?�����"O<0ko��=I���0��5z�
���"O��mє7��B�.��~�`�"O�H��4�d�#�-�`(��JE"O�%���B?�`�U12%Pp��"O�؀cOa�x�kTɁ]@�8�c"O���1��)C'���M	%�U+a"Oұ���6&� �H[,}V@�c"ODtkr�V:�p���Ƙ,pj�+�"O�GKB��F���D6�P�"O��{��!j^�`�fj��6�q`C"O��SV��?T����.�::�T0�"O�)�
��"�
$�عv
ƀ �"O��S�C�U�D2#B�0�����"OL%
SdJC��H�a�'ۺ��"O*0����|Ӡ%�@��(w�r�hf"O`���M�7Z4�`E$؊L���+7"O��H�YR=���Ӂv�V`Ӑ"O(�*r�^jiX`�E����`"O@H�T�h-���u8#�"O
�[�E��@�ɔ��yj����"OΘrgA^'�1k1���t@*X�"O��2G��*G���*�F�2P��"O �:�O͗.��8@-�����"O�����K�-薚)�e�e���y"�F�cB�����&��s�d�9�y"H�#�0\���	�2=a4�B�y�F�5���҅����@#'Ĕ�yR�'=Q�٣C�X��P;�C#�y�L.?��	��z�:�{6�0�y¨��Y&� s��iD��h�cM�yR�,a�^�:�	Q]�@�5G&�y�!K*_H�y�fC�N*�	9�����y��^/ I�h�
O+x�s�����y��F�Qd|�b�΀�\W^�;![�y��U�+gl�SƑ-D�
�s�n���yR��+X�b�\�feXQp�臜�yJ؟�|ʀ�Y�N	�Hס�y2��h�P 	���T����!��yB(^*R��(%c׌Ea��h��y�UYF���j%:�RI3R�D=�yr���CwƓ�2��D��@���y�Ϯ:��#�l*��l��)���y��� ��-�uj(���`��X��y���*3�2�`!N�5j��@	�yb�=J>�ŮĪ��t����y"a��'�h ����;�4�G
�y�G��07�� $�
��aׂT�<���� �\Mr��� ]� k��M�<��		 �*d��c��O�nMRU�JEx���'�6Œ�Fθ���	3G��\��'f,��f@�8P� q�D�8c�'�$2�bP�Y�1y���4jZ\a@�'�9enY"W)@�;�d�,H���'Ц �鍍i��,������&�Q�}b�)�G(KfHmC�-� r��D�o�k�!�$�c8���wK5u���PB�*D�Q���>L>�$fA�c��y`jG%o�^��7��fh<1�nio\�" -�%k���k�����y
� n`��OQ5C%h�;�����I
�"O2Iѳj��
Fz(�@+ѕp��$jA"O�P���H�J���)2pB䠶�i�ў"~nڡ"����@�I�	�^гg�̫:�C�	NM:���Ή]=%
�A�>�rC�	!j��İ��A(?���Z�'�o�NC�ɤ!��0��a��l��d1��>����	�b
H���E�z�v��$E�5R���u����B�=:����Ē?�|i
w�)D�qD�Gz?�4��$͔@�Vk&ʓ\֪�D���L-D�3�E$	�,��@��y�&A?����P�	��m���W��M����s� � 5Ν1o"���q�;k�ze�c"O6�A��ǭ|�ai�B0kٞ���"O8��p*�s�����R#g�2��b"O�M#@MiH�*�HF��%�#��<\OLeb���(�du�HU4���֛x""�n�'xqO�Y���Ƅ�3
�W:��4D�ԹR�A�0A8�*f�2�P�(��2�I~����(�g�R��@�*:W@K5$&D�8[�DMa��AʓN�4�� �&D�l�&�ڵaG��J� _9�v�K�F7��f��ħH3� �FM%z�J��ă%$�A��1���)�!�['����٪hϘ���XvF�g��KBh�r��
�vp�S"O~���+FY�<�ŧ��~�0�#��'�O$� l�8Y����Y,P���"O���(YUȑ�E��#��d��"O̰F�K�֌ �� ��rF"OV��J�-���7ӏ#���C"Oja&�E��"��[��:%"O���w/LE�*��E�g�`���"O^a���C�9���C��R?Bw��e"O6){�ɝ��P�z4EÒWcx�w"O�$(EBԶ1��� tdP�i��	��"O�����ӓ2R���C؅0����"Or����Q�cY��kS`D��Dȁ"O����@��%�mK�էG�����'/�I�G��p�oM�Y��B���ߚC�I�Mv�VF�?
��c6bC�IF�0��@ŵP�ެ�qʖ��V�>���	_"�$5 �GJ0GIX�ɖ>�.�S�O�>�8�m��3��M�AC�+�Ni��'��EAͯ#��0!2-�-z	�'l�t�N!A�*�pv,țt�����'�̓t��:A�i��㊁n��� 	�'%�P�f�ɣ�0��'_3tT�)�'# ��r}V����� i����'�v\��@&q���k��T;Z�MQ�'lҙ�0��3.�f��`��A8	�'KNEh��V2��Pc �M�f�u �'�0�����,�����B�G�hq����9�S��G�$X�8�5��(��R'�G��y�LJ�:�q�钎��H"��
��yrLHUi��8Cٌf�p2���yZ؈���1r+��3"a#ZPQ�Of���_�w,�����s-������Iӡ��e��B`܃V��i�e�+z�S"O<ay�i��#��ICoق9<�r"O���@�D?<{$�q���dTCf"O2�6"[X�I���0ט�چ"O�h��6#�ܴH�˕6O��-a�"O�ltJC4ؕ�\�j]��"O|l+aC�+�P�iT ����%"O� P	�u���l);ǈ��t�$Y��"O�[�U$T�2���eJ`�&0��j�D���g�=`��#�DQc�@]�ȓ2 ��.�\k���
�y�p0��'!�a	��D#
���dg�#it��'�H5p�$L#� J���)%"4@C�'2�s�l������įҫ��K�'�H�U�(��|3D"T��ٓ�'&� b��@3K�v۾�1��HO�!���S� ���B�ƗU���"O���SC�5	��9rfJ�� ��bQ������Ӥ3�F����V�{���AŤا�C�I0V@Y��>�(9��֗a%c���I*9�� ��ǋ^���H  ��B�	�P�2������TZG��/E�C�I�ܮtؤ	ک412 x�dܱU;(C�Ie�&�ʓ㞰_�VR2��.C�ɛ?{J�(�i�V�.�����fa�B�IM�d)r��Ķ?g�#V��
d�B�	��N JA#J�t_�msv"[7w��C�IH��Mɗ���U݂��\\�C�<����բ�}�����X�f��C䉼f�,AYd��<&�J'i�Dz���5扃'�N���6>��)	]?�2B�I� 脱`�]�St!��)հ��c������t���J�j'�+D��|�Ͻ�yrM1��ycӫE�1L���L���(O�P�Mu�3��w�Xq���L=��G}��ӖH	|�a艪W��@���+6Y�هȓg�.�3W"��-ც	k�2���hO�>U`��0,�֌��Y�a\�h�1D�H	Q�Z̑��NY,kh���(0D�,{u��y�H�aU5E��m��)D�DȦC�8�$U�d�΃}(�+��'D�`k���4ψ�`U-,ڴ�@�'D�$��@�1�T��B��<�����&D����G�@�r`OP	X\�(�
9D����-�E������6p�)8D��r��Y�jp���h@��/�>�����;#Ϝ%,�:Pس�i�P�j'D�����G�9G�x�
�*�1%6!��'���1$�5�T���f�,�&TC�'j���d��>��D��#�� �'� �b�R�J��g�,i$\Y�'Q*�c���9�(#��O���
�'SL�@b^�.�m*��PjeZ���'�x�$AQ�
d�G͍�)@l(	�'DH��1��!*A��L�Q	�'�<��T�fY��}48��'L	�A��9Eeb\���_��My�"O�Ba�=i���Ä�?a��"OR�p��]�x���eM�M�P�bw"O68[�C��(�l=h�%ުW���V"O�ͪbk�S���K�� e�!�$���Z����r����P��v�!���L�ɑP���;X�ß{p!�(�M 6��n꺁"0�K�P_!�DX&�6-�7�Q�n�P�I��O�yH!�N?y'�t�s��#;�DDQ���x9!��*m��@�?�����> �!��58R�
bn�	F@i{0�� �!�d��RBr!���Ѕ�h��	.g!���x���k��0VԳ��e!���pnr��D�EP��(`l�s{!�� �q�v!G� �xP4�J</��=Z%"O\�X#Mħ��ԀWE��oy��:7"O����6t̩��V�0b���"O���¡3D}��kS�*�P��"O���SG�/u�@�
�)���dTh2"O�mѕɖ�-�|�C	 ��F"O�XS�iA�n����4�E#��m��"OL]�AB��t��e�9#�8��"Or�Q�"h��T�6dpT�ӵ"Ot�'�:�6�A�I�Tk���"OU���-*��Вw�U=H� UC�"Ov��TI��L��p��F���A�3"O����7L-0P吙&�hYU"O.��R�M��ad_w B��"Oj�Y��Ԇ3*2}
�i�"����u"O���A�aDq;4�=}��A�"O��IA��f�[ Ʉ�g@qr�"O���C�Z҅Y��c�: �!�dX�d���C�>9�;�bZ;+!�N�N��Kr��u�=��!�F#!�L ��kSFŷLaI�o�t	!�D
�tI�v��B|�Yv�W�!���K~�@�z$�	B��!�D�`��"��+�d)���/n�!�$E�*"��p�䋐]J�P;Zi!���&*��S�#`�S�'	,|�!�dY"?@qpfċ��F�n�!�N.!ڤ�ҋ��&"�c�N�VF!���P���4 �5E��`��QO!򤏊rV�1H��2L�)0C��5k!�$K�g�,16�8(�1�C�ItN!��;�6x3���Z	�{C/�.4!�O�hY4�#��Z�K@�!�ϻ%��i�"T�]΄��	A� �!�VuӢph�ː5 ��AqP��!�$�#���*�
*�ڬ�&#ރ%�!�$�(����+�? ��l����!�B3O�|�WYюQ���O�d�!�$����;���%[n��C����`!�*� * +A��Cʋ�aw!�ĔF
�!�l�& ?`%��)ac!�$-0u�Ѓ��i#z��3eKrm!�$Ҫ��Di�+�H��2&Z��!� �,݋P�ەO��-q���N�!��D�f�ii"LB�\�j��i�\!�$C&0+<�$n�#��d��}<!�?z��<�-C[�Pݰ1� �-4!�$-Ȱ k�جH�BT�w��&S,!�Ć�U�$ S��ؔY�@XG/� W&!��ADC2�M�>�� ��-~!��
�v��A˚�6�H8A��T
!��ǋ t�s�Ŧs�֝��NU?�!�F(�� 1ã�c�VL:6��.I�!�dϵ(*8Z�'��"��4����
�!򤄋;�t�j P�LP��C+^�!��G�Nʆ����<oKl�OO�77!��<KL��t������.��
5!�G�h��#���_�8�	��H�,7!��N�?��T��NƴL��Re.8FN!��<;:Yi��W=g�R��`�V_!�dx�.��#�33���k�&!���"4j-�Gc�&M��t×�H�H�!�O"����Z6g�`�U.�!���q<쬢w��8[d��r7�H�/�!�� h�V쀁�R<q%H�-aZqJD"O<8;�+���ڝ�d�.aV�)"O�e�T(�$AXh���xKz�$"Or ";\s��JFCF(F`Fu�"O�8��%���	�R�Ȏj�Xq�6"O*i����h�x7��
H�h@K�"O��p2�)1A�����|=�G"O��PKؽ3�,�ڈF)�A�&D�LQw�Z15j)�S
KN���a�#D�س���>^A$�
���c+�H��A!D���'�
H��Y�f�W!xiH��i>D� ;5dH�#ٸ(�@��Y(�/D�����'fNz��fRl���:Pc?D���*�+��z%	Х3x��2-?D����LT�A�a:��BC򒙨F@2D��3E�8W�bh��H�IwX�q�`0D�,``=��#�+(��.D���̓)|���] �� �I'D�p�� 3n؀@�5��Xʰ *D�L8T�9����cD�'K�0�0J$D�t�*�A�r%���h�t��ab7D��S2�ϡaҙ�6(��DPb(A5�6D�T��ʒ�4%�1�K�p�<��'4D���R���kn����*��XAn1D��A�+М���i]5n)(��a�-D�X�PKQ"�ai!υ^i b�!D���S$~A&Q��͙h���'�>D�L��V ?zZ�ȕ���hȤ�`�N<D�<1�Mܹ3���Y4�Oؠ�Ӂ9D�(`�Đ�mSD��u�]�Lzd-��3D��!eO�zN��XEn	�6�ѹE1D���׫�(-��DJH�U_0�9֢/D��2e��&�%�� ܳF�YiU+D�0��)@7D:d���pt�-D�2����u����f��a4���o.D�D��`����E��·�>W����+D�XY��6N$)S��oh� i�*D��O3���c�Χvz� �'D��CѢ�z��bh�8X2����$D�<��+H�bH0� tM/T����3�=D���ï��=�f�r�M�8y��;f�;D��B�!���`A��7���;D�$����G�@a8���&*R���n8D�ôdN![o�XSW���q��l3�8D���K�{�ֵ�`���#LIZ��4D���4T�|$�1��g���R%�2D��@�-W�SGˈ̴��0D�P��մCrj%P� ۥ�q��.D��R'�+C�" �V��q3�	�'�+D�<��BڮU.��òl�T��u:��#D�81"A+I��cˉ��8��2�.D���D܋4��i�	�b~��-D��)4OI	��T�T�_s�s��+D�㓉�G�B���%��8�� ��%D��Id��#\��2#�q�n]0V�&D��ZR�΂d�\���	2ovF%��(D�`��B.K�*�"&.R3ft�d+��+D��
���4o<&ݢ��ZR1r@�%(D��Y�ԇwjպ��ٛX:Q��&D� yE枸>�4�#�
�!�(�&D�P	��Cd-vH�6(��n-�y9fK$D��bP+��6�k��O��$rd#D�X��V�c��ٰv���V�Ļ�"D��@M��N�:�A3�I�h�NC�)� (�S'�E�~���u�?v7��y�"OҬ:��̵f����*A#3l�ك"Od�Hb3�j�"��<B,>�p2"O�`ꂀ�?���ɰ��z(���"O����bW W8L�5.� Avhf"O���$4zn��c��q�ٓT"O��Ί~��k�ň	�x�0�"O�P	���#�`U�$�=H��|X#"O܄Qu/�L �11�ğ�X�B��"OP8X�� m�-��\X�J�K�"O`�#�K� y�'J2�J�	A"O"t� ث! ���c�����"O�D��� ��e��I($4�JT"O�%;REȹy�T�1�GP>4��C"Oġ`A �2l>F��W	�FM�IC�"O�%0��0n^����B2�ze�w"O �&�/��aR��df��a"O,�j#��0Y	p� �ɒ&�>�ؑ"O�,�r�?R.�������%�.pf"O�(�g"��?�ܜÂgܫ+ʉ "O�����pv��"f׫>R-�b"O�h
U��}��eO�7V��r"OQ;$�%��'��Dn�
'"O��1�MH�Ci��A��(��A�"OD) E��br������r��s"O��S�O��@���/)�ƭ��"O0�h��%@�<�-�%l�XxYC"O����+Z�yb ���[s�l"�"OpX�̈́�B�<�g�	.���`�"OFt��D�>u� Ĺ��[y�pM9 "O2���OO[�s�(UL���q�"O���&�j���q5���n����"OZ���2�Z��ۙ{�rTj��G�<Q#OV2z�|�@��豃I��|�2B�I�M�	��X����sO�'m6C�	��(p��V?v\�`��3uTB�ɪ>^���F�!O�*�C�_���C�	6���!�mG�=��c	�
��C�	�t�d3� ����S�,v�C䉏_���kU�P���:��G��\B�	�`������F��ԁ��=
C�I/E�����I����q�B�	�4��4AG�[�D|rA�L0ʡ�d�!��ᡦh��?"J,@'�r�!�D˟<��QqƝCb,� ���W�!�ė��\myr��H[^��Wl�!�
��Q�d��Of`Q�m!�K�z��!�I��o<���я_�!�D�.@��)�O�\4��;Vo��v�!�Dʒv꠸"�.C	"j�9���!��T�@��+dO�7>��ؤKh�!�d�h��5RT��	K!�QА��p!�D�+0{����J�t0�y�-�[!�d�Nh��IuD
2y$Q��G0�!�D�,R��gOˇu^�!&�'&�!�D��a2��zB�L�	j ����!�Ga���1QL"IМs�ϕ�!�D��bikScO?<��oS�!�d�)Le��j3�I�<�<��-��"�!�$��<�3�`X�4��D�D-��q!�����C$�̚E^L��&9p!��X ��i!.H 5f0Q�� :c!�� ��\
�k�y��@��	Y!��M�@��@�{��ؘ$���(�!�� ���VI����C
ȟW���"OC�dޥU�����"|����a"O�X��)۰D@B$.p4"uj"O��Y�*
��e"�%H� �)��"O�o�>�iX��'���X "O�۳ �����i� ��i7"Oȴb��K�S��t[G	B�l��aD"Ol����S
�,�#�i�,ў�cR"O�l[Sm�)Z��0�C�x���z�"O�H����	8^lA!���bR�	�"O����N�1o���AdX CL�B"OƁ�G��0�P�q���-*LlZ�"O,����P4�YꔮY�4��"O���E�Vz���t#U�{�� "O���.H�
���
jO��1�o�<�/_�>�����@ˌ�.9B�$�F�<I�E��2B&-���Tuιy�L�@�< �?88S鐟m�HX�1(Ve�<�ej�eH��xv� �M�H)	׫�G�<�ӊђ�r(�I_!Ob �eMD�<��[�|��!��W)Aa��(���[�<ٶ���!2�)��e��F���KV�<����ă�hf���w�<�7*ǝL���!n� /��% ��J�<�*E�&����Z�mN�Y�C�E�<GK[�]`�1��C��Z �D2fD|�<�SQ�;��t�\2���kz�<�F���&"����fF�g����e�x�<	��!i0i�K�#B\h]�s+v�<�g�$�<����};����]�<Q���
a%`�z�mV�RVtɥ*�C�<����$S(L� J�g�$�q��<�A�ƫO�6𢇌��~0<�h�s�<	3��jHE�����t/Qk�<p�B{`4)��A�%x�21�%K�c�<I�GV"f"�@s�<� ;���^�<AC��2樅k�Kܟ0��[�`"T�9���$Z=���9Uʈ�
1D�x�Iԩ\؅�E��-njM��H"D��Y�*�n�ܔr��� T�b�!�=D����oT7yn�iE��3^�ĉc�6D�L�֣R+y� ̡X�+���FM3D�D𥦕�$�5��c�r����*1D����gJ �&�7-E�PH�C1D�xidK+�(l�W��Ѐu{��!D�����K\nxz�K�� JT���o?D����"h0�łG( ,>)jW�;D���B
X�{Vi
'"�Q�d �7N/D����JK37���W�J�v(i5c,D�L�ݔdfXX{�.#� (4�4D��Ud�@�xBŋY�Hc�4D�0Za,�2a~�h�H�C�n0�h2D�L��hӿ[�p�Q��/.���t"%D�����[�$F9��HQ�I},���"D��H� B6��Gůzi1�"D�p��b�,!���PkB<\{�0x��-D����J�:x�a���R.&��㶋7D���6	�LZ����'V�Ѩ 3D����F�)8]r��`M�6I�~� ��2D��Â޶f��Z��C�4)��N&D�DK�S2'^�`�H_$?����� %D�,��"N\gf()�d�2�@�bA7D�`{�.΋s��%{�A[�O&�r�k(D��ceе5[�ӡ�, ��	�խ;D�� �,������	:�����@���"O�Z��r��l� �ƿ �
b2"O8`�jI��t���jr򸘒�"O���@)!H�"� pJ���b�"O����'.�<��IWZ�`B�"O���kǴw�rɐCoŁ2 ܝ��y��'C*�|BBh�=h��dZ��W�y�锥3.���m՟_��*`��;�y�I��_1�i��G��,d�0�
;�Py��L!�vɉ⎗~��A%,�|�<Y�O�4 �~�[�*(l�
t�)|�<��]
soJ5�A熦c�\Y-1��C�ɍ9�~���D�{Tf�JC�?4�XC�T� jŭX5k���K��!$C�	$p~͛gړj;��З �{�LB��4f5T���v�sr� ��C�I�5�^AEH��6ˬ���� ��C��~�2Q��sJ�Y1�-R�C�	� '��jq4#��B��?�b-�1BzU6��g���e�B�I� �����)_��Y-A03�B���}�r�ǟ<���������͆ȓ$�j��3�!��I��cI:Y+�U�ȓ>+^����3g�9�4��9,��(�ȓ}Ҟ|�p�F%���b'��$R�U��f*(�MK Y\����h|����]���bv%I�D� <����M�y�ȓI�j\�����}s��� �^��ȓyq��$؝!Xqi1B�����ȓ`�¥���
�D��`1e��9J�d�ȓ>�X��6�#9�.	i�)6&aF�ȓ7�جR�V?tt�q�s	̹���ȓ&�4�)2✈̌���}���ȓm�Rc��,���)�M&F,�̇ȓ!	�����Ac��V+U����ȓ~&X�Y�	�<��!��]�o>ͅȓ6D�˖e	&����ȉ/u�H���xĕ�D��oF�u�rJ�,f⥅�w�Α��DR($cTܫ.�"U�����o�<�Z�I�0@ ��F��/��P��0�p�x��0R<8Zq
��<�ćȓ
@��0 �B�$�K5y�������� 1P �t�P-wn&���7x�C�Η �pԂ��H� �ȓb�!��mۆ#�N�3WJ�'�5�ȓ;���5�	r ��%���/% ���PCb�#g;��p΁�r: ��ȓi�R9;s*Ƒ$����o�%f'.؅ȓ..$�Cs׏a��A�
8-��ȓI��ţSG·KBP:���#Ŵ�ȓ
�,e���ˈ,��@�ǥ�)c�0)��3���:p&H=h�|U�W��*�����!$���U���\��X�fԧ8(ͅ�)��X�E�nID�q�ݷ3赅ȓg�6}v��=HJ�Ҳ�ќWj�L��%� hk�&�03X���6�]�=�̈́ȓA�-��EWU~����B꽄�-�}4�Q�(l(m`�d��<�e��0jH���@�nl����S,X����7o~t +�64*��7M��DŇ�?�b)BqM)>!�HN-�h�ȓf/����`KwɎ8�dA�)wfj��n��b\l�0�1"�"L���ȓ}�H(�� L��\9���
�Z|��S�? �H�A�M ��e���� V,i�"O�1��a�v�x5���2n$dD:2"O0����HMc�!K��եV� �w"O�Py�e	��XE��F l��"O�Q*a��)ֆ�����o�����"O�}k0����U�a��Q��Q"O$a�r�.z8��#�o��|�̜
�"O��kW�X.B�P]J��媍��y� DM2x��&ݿK�t[��J��y���Ft
�q�M���B@���y�̊?��+��h\��C��y����T	+V�)���q.Z�y�MB$r���3��j&a���*�y��v��
C��9RjD���'��y"K�6���ao�9VڼX0��y"��	G`B ��c�<Hr�\yPN�y򮄦fG�y��S%jSB��
Ҏ�yb�\��z�P�kL jp楩�B���yr'�sG�E�i�=f���i�@؁�y�	=Vd5P�
d0���K9�y��M�3�n�b�M��s)�I��yN�4���߆f_�<��\	�y2���d\0�q�� ,Q�Wb���y�Ev`�U84!^�r��dP��y2��#6�n�#P��d�iRG��y2Ë�Y�*1kC���iF)��yr� 6W�q��D2{����ַ�y��Z'M��<����{�rE�Y)�yrN�)=X5ҖC'oR�]�w�7�y¥�Y	L�YC�c.�F�0�yB/�>zu�\*��7]��p�G9�y��	�
b��AiN�P�8���#ϓ�ybS�b�J��bt��+��y�KnÅ �&;m�%j�W��y���=(�F�L�0��91goL�yN�q��J�$ӇV�H1L�7�y҈�a��`����U">�sGk��yb(�.+����dfğ8b���ʞ�y�'U >l��	�m�:x�� xq���y2��{eV�)�CלuLBiy��G��y��
"�RRp�Ҟh|�0u�ƣ�y�bV�V����4
�M&��	�\��yBn$)��Y��"}�z�)�Ȇ��yb�=-���iѯ%b�E����/�y�Iǩ�P��䍒72�z �G�̕�yR���
QR`)Z�#f}�6��ybEO�t��\/#��Y�EL'�yÀ�^S�M���
��D�r�D��y2ʝ
,h8��N_h QR)�y�Ş�+ټY�6H�eh����	��yr�B7i�`t
��׊u�PE�Y(�yҎ��4��ũ?����y�@R>@H���0$�x��}�����ybgψF�\�r!kQ�w.`���&��yR�H�'A��Y�է;L� #��yB/J�Z��8i��S$
0r#k�yr��05s��g��D3F���y���'"DppB��;>p�$P�B9�y���t�d�A�*h�ʼk�c��yr�wU$8��c8f�,�J�Ȗ��y�i͂S��Zv#L�L�ffũ�y2!]�z�\$c��Esސ	����yF�t��@��P�9�d��ƚ�y2��>A�d��j�|��p�FM*�y
� ���k]4t��	�C�����4S"O� )b��-m飗.��P{��HQ"On�� �� Bm^5c�O�4Gy�%z%"O��Ѧ�6u�p���0R<��"O�uHڊ s�i!��	4�1g"O���Teܫ	�4�` ,��v -�D"O���Dj��%
��B� `�"O4�KA*�=|�yaP(�D�BA�"O�9sP�n�R��r�s�� `'"O: �P�É-m�xePZ{
%)�"O6}�Al
�P�N�K�iK�$�H�"OR��R�$#�j-���$w�N@�"O樳P�ڛ:a`���gP
~��i�@"O>I��iF4`� ��1�C	���"O(�#��3����PШ14���"O@�b"��8� ��"[FB|ۆ"O�$�"�R�z�D�� ��`"Of�q X�N��]aB@�R�(lxs"OL��T�J�-D�)�aK�4�fQ�"O2�C��\�%
���u$$ۀ"O8𑖣�g��XS��Z�a��1"OR��D�+2��񃲮T�Q9t�)�"O� Ĉ��~5Y�M�;���xS"O@l("�20�M��M��W��%1"ON`;�������,Y�f��*�"O�tY7�VV��0v+Q)�b+Q"O�3�\�E2^d�R��zjQ�$"O��vH�YRiӕ��6Ve�"Od$A�Gՙ\6��怩ctRB"OZ�1%���6���S���кM�w"O�l��K7�� jG/,�h<B"O��r�K�bL���U�h�����"O2�EA֜�^ě.+,�|k�"O���7�^�Ґ�UЌh$��i"Ot�(��
�k�>�ە䕁A�T��"O4\����28�-Q6�7<���"Ob�Ŋ�(mfvXّ#�$9h�5"OD�٠e&�(g�X�yAb"O��:@+�J`><"����N8tizd"O�Y:��R���|ѕ�l5��J�"O^I8�ON�z|��a�M:`!:�X�"O2=z��K�~��bgDN+y���"O���1��G`�b�a�2Wl�Ƀ"O|HtaE&V��4�.çgC���G"O����HKrX1m�uj�sp"Oͪ���0H��ǔB��{s"O8���#y�F�R��Ϩ�+�"O
�jv�ʅyǬuʅ#P0���h"O�R����E��CFC�Y��4s5"O�!��7_&R�AQ�-���{"O� i�̎�2!+!ѢC�$�#"O�����g�x��j�*9(��!"O�m9��f4�"���<q�,��"O(
 ð;"�I��m�9����"O��W�G{P�Y"b�O�-��!��"Ol��uCУ=�&�����,]�4�2R"O�@����O�Ơ�S���Aa"O�}!���<pɪ���2}���w"Ot]� ��?����6�1n����"O�`@�ÞV�{V��.�:Q�"OЄ���;3^��$�pՎ�k�"O����8rz)z�dQ&�a"�"O*����Z�S���[#	%P�h�;"O����+�F���hڦ�p��"O� r�٣�3�Nu�1�w�j"O�٣�NX'go�,�F�����Q"O�)v �r��A�l
(M�xA0�"O�s6�ȇ;9��9�t�T%��"OP�j��.`��}r&�2��"O�� ��Z���ܲ��HS�q�"O��Ao�D}ģ֫�8�8�	�"O�ٸ'ƦK0M��
�#t�Z]8b"O�mDaL-��yE�͑^��	"O����_�j��֭U�����Q"ONt�T�CW��G*?u~p���"O`Q�L�8�D�i7O?Q�Ek�"O~�`�G��W����OF�Z�v���"O�\ â�6�X��wNĜA�X �"O�4�ď�����ƭN��8rw"O&��b��
�r�1u�H�tD,�"OX� &ʧ�"%����Gd�ģ�"O�q����.w�8�ʤ(�TX�Pb�"O2��%�q�DЍ� \9�	��"O����B�Y��P#���9�]`"O�ŪV ;�5e߃F�=qb"O��f'�(��0�D%J�#��6�,D��0���@�Z���g�D>.M[�M)D� �E��e�2;�1R�*D���PꝣQ�K��#�4H���&D���䭏�Zo$@+0#�W�9���(D�8�ѯ�x�/΅��ӡ%D�D��ɝ�@xRujǚ|4��*�6D��r�Zw��0�Z�P���F��yb̍~�dp� �aS�A�#@�y"�ÁFrp0�t��	f�s���#�y(��6$��r�@�2޴���K�y���#P��BuOM��(E�5�<�yr%��ĀA��)N�|$�LXP��)�y"Q��e
 I�s���0���;�yҨ�UW����G�)f>B��ׄ[�y���6���Zi�,Z���^�yR�Z�H�q�F�TG�� ���V�y���U��5���"jd
��4Ꜷ�y���î��5�a�&M�d��yR,��N����1Ds�D�̙�y��K�p�VeHe��C޾���^#�y�'��0%ݘ,����y��1$�t�ȵ�
-zc�d�U,�/�yR��3�*��&�I>t$�\1B�G+�y����j���+x	0��#N_����ռ8�7)ԍF��5�E�)kU:!��$z��K�Ƽ_AZ�k��ئT��|��W�Y*�ȕ�m��0Г �!k���]9�@$H	�B�E�ٻ����̌A2k%�\�#q����@��2#����Xd3�À�;�$���ua�yY�ēcz�DQ�ǶqwD=��c,!�$�6��0���;>�
�ȓ9D!j3�[9&�A����7
����_Y��b`��'����攱lt��̊��s�[�+/Xe���W�U��@���4�y�oʯn�f9�3.�`B��I�U[�`J�z;@p�`��;	]���A�%�1��20QH��ܼH�0i���նjO�RqD�iԠG��� �"O�\�!o�W��!��
+_y�mKP"O��2k�oV.H!�S:z�k3"O��D�_�0k^p��^0
H�F"O� �(�0k=LJ�${��S� ��"O
Ez�i��B`���v-�6V��z�"O䈸��J�^��8���90tX�Ӣ"O�k��W'/�hT�5M�n�Rp��"O���8+df`��*�T�"}�q"Of��mJ�YX�
�J�7f���"O"ej�"_�m���j�jU]2� e"OX��$��7'h�AV�O�G����"O
���)2���=.n�XW"O6-��b����DX��#E"O��U��}N8�hw�)'�DR�"O�H	�@B�~�\�'�S�i��iV"O�Pȱ@SQ�\�#�5z-����"Oܹ�Ea��z��٤eN�#PY�"O�U���I�x�2�PTCX (/F�D"O8d�,���a���{#�ԢC"O$:#�B�
�t�s���;d8�!kT"O��I�Ć�T���rA�	 \"��qv"ON���
�� �)�i�v1l��"Oe:1��F����vゟ/&䠔"O�=#s��;cv0�b��x�`�"O\�yF��'�6�i�cߒo����"O2��iP=U�섰�Â�v,P��"OH�1t�Ip��{�⑐W�j�3�"O�HR��2��ٶ#<Y~(���"O���5�T0�,Loe�� �"O�40@m\�X���9��O�3dn�zv"O�a�u�.� ܫ��H$e�tht"O X���ʆmv�r�"��<�00	c"Ox��'���>��ω�8h�"O���O)[d��2�Ŀ`L���"Ojl3���Y+��ɣΔ�e^`={7"O�8)���B�;@'P~�
�"OL��U)�{l���ڕDV@b'"Oހ)�$�	U����$V�r6"O���"B��R�ȑ�]72��u"O�]��	�����@!�ф��p�1D�pAo)q,p1`�ӕNm ��A(0D�l��L�s[ܱ@�̛�#��M�r�/D������z����֣;},ԡP*O�Yz��Vf�$DzsK�;8X���*O��!G� ��5��/��p���
�'f���D�7H���f�%}��y�'�~���
�*�s�u��m�	�'� 4�Jq�6�	`iG�L4�	�'��E"�NP�SH����|b�
�'�2T�V�C� ���{`��x4<U�	�'R�� ��^�	H9���ő">Z��	�'�.��1�E�-(�ْ�&�l�	�'
i�, )��U�T�X7���s�'d���̷^��\�Wߝ{��c�'{6�ZN��X����!wg��(�'C`�Z�g^�QS�<Y�m�&>��z�'@$P)g��>g����,�h���'k����oԿ`E��
��Q�<�1�')̬*qB�	�4�H!�Y�~���j�'��c�P�z)���@�WfR\�
�'��4�ȶb[te�wD�7^*\���'�B��b�:?�PlAw��W�(H�'����Q�M\U�
�d $�i�'����Fd�6#��x�m�0څ�
�'u�tj@��F}�"��"o�h
�'i^�(�F�ܠ���u*
�'F<rb�4�ސ��׳ L��
��� (hap�8N��"j؀5����"O>�����{`f `�GY�����"O�(i��Ą(�d���D:"�D "Ob��rh�i�z�L�<D!qB"Oh �&��2$'r�W��p���"O��n�
p����}4���"O9sS�	���r�
��Xzr$��"OR�xe+�^���Ӈ
�ĸҁ"OF}����+2��m��{�iH�"OL�2�C�+lx�	��)n����"O҅aP�M�fպ��傭ld$��""O��T�[�Z��5�.^Ph�1"O�$�Ffݣ%j(C��D_F�H�"OЉ��R�a�\!2��k9� ӂ"O4Ժ�hM�G(�5�����-�!�D��|�������Yr*�����?,N!�ȌHG'�����I7 ��]!��4/Le	�h� (�
�I��[:nW!�DUr$.��5APH�*��>!�Y2Z��=P"a�i3�AJԈ52!��`(>Lr�'F(�
-�c#ބf�!��(]
(Q�QR�<P(��
�Tg!�D�8�*�%)(Z8�y"B9U!��ΗLafirUJ��|�&=ʑC��!��6��Fn��{f��D�%s!���*9J��%5-j�����u_!���m�\�S�HڑR�XǗN5!򤉮M��|���A�L2�Ba�	��!�䏵k>,�%+*�j��]L�!�D�uܸ��Č�����!�G�AC�<�tJV.ļPiW�6>!�$ǻ'�6����B�}�H�(��L2�!�� o#���wd�v�,��U�N��!�$_,#������&_�@��
L}!�D_�R�qg��?6<��i�,c!�d�:�ux�o�:��đƪ�T[!��4ez�٧l�jeCKv!�\�i�Ĵ��)�}V4�*��$�!��L�X��)J��11�0�!��ۡH����夝� f�]���	d!��T��Q����P\)�%V�<!�3�zy��bQ�m� ����ȳF�!�Ĉ�A�Zms�W4D��8Ԃ֊>�!�dʤuj0����r�Dq����`�!�d�=wpҀ�%�"O������El!�d��,��	Y�G�T�҄S�X�Tj!�$
GP��p��<�����N
-e!�֠�L���֥Il|��ݟ]!��U�m�p��E��U��T"����{!�V�1�J��(Jc~���P��2|!��\$��aų#c�=��,f�!�@�W�6|;���pY Ł�aI�JI!��o|��eH^�T�ı�/ �!�d	��P�ؐ'N?a�P���#C�}!�%F�Ф!�ł�H�~�����&,!��0�>���.=_w�a+��<�!�$�j$��e۪j0�����s�!�d\��4����[���ņ�7�!�,#���FO�)}�<x��D H�!�D�1KTf�A��?}��a$d�!f�!�dlS��4D�;u��A;�#?�!򤀍c�J���)v��(��B�!���,��U�$	��c�D@�a�v�!�Ę3q��8`��}� t"��O7�!�� �%��+[��8��b����̈0"O�Q邉+ ��P�r`y�"O�l��Fӌp�Ȕ��&# ��R"O 
�	
�����>X�"O�K�BS�'�C4 H .D��"O�k�Ȁ8$2Ei���97�Y"O|\u��2A:d�B��"7���E"O����X�@��	�&��l��)�"OD��Rnչ(��e��J��X����"OТ�k%>%h����H���[�l!��!  �А�0tИ{uL�:�!�$j��d�k2�cU��25]!��@d���#OL�P��Ɉ+P!�$��Yg �$͂ΜdÆk�?!�J'��I� �C�Z��h@�6I0!��Y~�C%dL�`�08+���5>�!���5���CX@p`&n�1I!�D�+���	�m�4k8��'n18.!��N�'�b#F% �^��A/Ea!��'������¨#������j�!�$�Q/��Y4NĹr��H*��M�P�!���<az��1�ϡ8n�h1N^$�Py"-l�`15ɑ%<Y����yb/�.���L��X#F5��9��B�.�� �MW�'N�R�D��܂B�45^��R0+ƪ|mJ��g��,C�	�'Z�٦'O�Q9Va�Q��.R�B�ɰ;2f��Մ��dQ���S�Z?s��B��8E&\�P�
�O��e��.X;\~B�ɗK3.`�F�q��d��,7AhB��"A�p����7 �z��r���"O��g�ї(R����S�Պ���"Od�HD�
#M�H1�@����3"OX5��̍�fD�!�Ċ$P��L�s"OR܂��0��0�⥎�A��ͩ�"O:��f�OY2��g�����"O��!��S�~���+�%�6(��I�"O��x�ӧXl�����ţa�y�"O~0�W�Ǒ-���k$�\+o��@q'"O`�r'��c\������3����"On�K#e\� L,�@3a��]�$!�"Oެ��C?uJ�%s'#�)F���"O��8�'"XB8��0 �(ؤ�J��y�ֿw��S'��	���dIM=�y2�7˶%�ҟ~����F���y�E�&~
`	�a��{��)xé\�y�%Z�O0�E�uI��K�3!T��y�^�*�"�)��	�I�TI�2(E��yr@ ��)�Rb�=�Hܡ��ã�y�e�r�K���`��Y;�m��y��W�(:�;����W4��WƓ��y����3-�S�`$��`��yr!/I�+4Nf�qQ�#O#�yB"��zml}1��ۉC�p��to��y�����Ma�G
/�p�)�)�y2�J	l�N�:�$��)�>��v�0�y��@�!.R�����5*x�A�*�yB		(Ƃu!��ȖYDt���ܴ�yg�MyR��W��HWH�iu��y�3��Q����>L$��7�ܓ�y�jë~d~��hM�:��Y��#�:�y���V�d�C�	�
V��HԺ�y�  0�섳��Ř��%W:�y�o�l1.])�i���*("q�"�y
� NQ���>G>J=Y��D9/�͸�"O��:�a^�.@�#r� F����"O�H�küQ �uE� �:�"O@@�U ^�j�12g*P�F֔�T"O\��J���*1��Nt�� ��"O������I `͓>��py�"O�d��엺.PXX	�� �6x��1"O�u���Ǭr��(�3��Q2A� "O��&�� ��r#\+a�R�"O"�R2�B,W��Iq��,:���R%"O��Á_:6�3�F<*頥�&"OJq���P���Ӂ��-�b��"O@e)��7=���4��#m��TQ�"Od��v�ί\�b9XFǚ	�<ź�"O��{PK�jc�`*�ܑ4t�RW"O6̈E�!A�
�8'$�6y�}0�"O�]�7j�3^�hH�dݒ c(�+"O��p�!]+H�d�ɥ��:q�L��"O(Ib�	�`����Aơi`%�"O�ݳ������@Ea���3"O���s�/�\z��O->v� �"O�%xFßN��8�n�$oa6A��"O:)ZwƝ�37pp24M�!/aB��r"O8�B3ρ-:ij�(�J�*=���u"Ox�fb_�g�ĒTE�%<׊��"O��#Dh�C��0I��L��5"Ox虢"�R߆dˑB2(�z9��"OFa)�X?K�Xy�y�G��SE!�䆌s�qۄN P�d����$0�!�$��r��Y3�W�}�z��Č ��!����O��AE+�K�|�q���>c�!�$�e���W�)N�2t����H�!򤕌-h��vC��kn�!�a�0�!��҂#�'umb�S���Z�!��uq(�x��_mb`�4��S�!�$ˣ��ye�dU�Z!B�!�8|Y�=�B�Ɓ	��ȁf�!�U�M�.����E�[uP�iZ:!��4�*R��x��%2��m@!��7搨�'*s ��#�%!��vEN� #�ԍ|]����6!�d�6Nlm��� �~�$�!�&1�!��U���F�&)6��fH7!��6\�N��u':t&M�'ܧz!�ӽ��Y���*w
�yQ�(!�7yo�أ��K �����ɺ%�!�$ȍy� �P�_�X�̥@!n�!��*t@����f�����D-N�!��_�D�Bp���݃ ��2� �!�!����"Q <}ѕB>;!�D��A���)�<%�X��N��d8!�$��v����
��?������߇J!���1>{�E�K�P���&�;�!�L ��yc�G�)CO�Zw(�Y�!�B��a��
Gi��1�V:4!�dT~��P�7��de�	��F­Pb!��K*�����Q��HV�\!򤔐�6��;�ݑ@��n�!�$K6B��1X�v��U�p!�dzt���_2��(�7�]L�!�D�k�PA�H�.AA�5
%#��lu!�˚G�.�H��S'(��U.V!��ԑt�� 8M��a�J�]C!��2��m{�(L�u�����r3!�� %	"�K�v�JAZCDO7��p"O$�a��O�����M8{|H��"O�C��#GRP�MnoV��"O$9`AE�	��M��
�QN�}��"O���@�Ns�Ё��C[^K��"O��	�%�(f�����/I|�ф"Oz��ȣV���{�ǳ&+���V"Ou �nȐ*���F�5޽HC"O���g���"X�i@Ŋ����x�"O�0�E:r[��rV�ރF�ļ�"O�ÌI��s���� ���"OTI� ��1m�fSe�0nƵz�"OD�{R��O�<�# �7*	�@A�"OF���26��hf�{�y�"O<i�v��0�4qY��C�
}
�"O������!rP%� 唟4aZT"O|)���'5�Q��&K8p)BG"OFXh��Y�XN����ަ{�Y[�"O�Ě���P��U�EEL��r X�"O�=ٳ_��� RE�)P*��"O���I��
���N�>�sW"O�ٹ�l��� 4�ǃ�����g"O� P�Fb�Wb5���"Ol�C�cf���sE"�8' �"O�����A��U�Ю �&\{"OR	+��30���#W�:�J�pq"Oh�;`#9쪸;5eԏQ��舥"O�2r`F�V�l��@cx
�"O<����)8 B6:\��"Oе�gҰ� ����Y(�a��"O<d���5�~�	TA��Dź	 6"Orѫ#�<tJ�x�S�D��`�"O�#.�#}	��[r,�V"O��ck���æD_�
`X�R2"O8��	H�r��"�S�I�&�f"O�d�K��v�r5�w��ޅ!"O0|����Q��z6!3Z�D�å"O@m��im�$�r�A5PꆘA"O-`#�O�X�P�@�	6+Hp��!"O<�R�/�$p<虪���1YV|�f"O�h�񤀅t���y�	3$��"O����1.�a0K�-'�$%"O`1Rt��!S|%��l�
UI�Y�"O�B�aF%k�P)�IQ>+d��&"O�0�"�St��Cg�7m��0"O���v�T������e��p��3"O�ؐg�ȩZ�������V뚡3�"O(I�Ǯ�vi�m�եH��iJ�"O����H�9��X��c� "O|�@��R9)Z���5�\�D�j���"O���
|ұ��M�"(�.9�D"O�<�!�QJ\@9歌�!�:���"O -�ĥ��N�����ݣ5�~��"Ob�r
W`�Ty��8���"O��@B��@"3��Z`���7"O�=�w#BB�>� FÔ5p��"O�,
�b-�H$P��Ǵ.�p�	g*O,�3֩�9C8��4�15�Mk�'������߁��z�>���J�'���J!��j�VT�c�1/�U1�'��yR.��$����E"%��H��'��Ċ3�;il����^&�a�'Ũ4���S�Dq�����.����'Yf��p�[&S��,[���f� ��� v`J�Mȏ~�B�B4b���s�"O����¹�콻��A����"O��PG��{t��t�I�A��J!"OTб��/v��c�KU��^bd"O�����܎"8>�*S�g{�"O<�)6�U�Z1f�j��ߟ'�Is�"OX<	� �.|�d4��bE6E؜z6"O� a҈�>��]#� �`���w"Oh���̅W���� ���c�<4	"O���j�/Xϸ]ص�.i�\(SW"O(PF��2v��	�.H'U�B8���'�ў`�2f�2L���a٢ee0D��5o^ w)��['͎�&0n%�uK:�	f���S�6[�0�B*Z�AS��W"�n#=�N>�����S#��I0K�o�VhSS�U��0��P��f����E_�rU��r~�� )2!�N�kp; ��{|�d��%D0Z���'r�qɄ\!gX�$\�#`�'��$���g�ęR�hMA ͞.vhq�<!�dn�(��>�ʈpmڏ��O��=��490�H�s	�as4iʿB�&�K"O�݃`Dֺ0��3�;%]��>O����l�6t��*�Tx�\	bDOj!�ĕ��q����[i#"DɔGK!�DL�=gt����ʰ3V�@R��.1.�y�(چ�)Sm�Lܼ���žJ�H�>/=�I�|B@LL^�Y�$e�+u� K�	B�$#�O$0��&B��|��d�r��U���'��	�h���f��d�l�ذj�"�z6m~����ɏL^��w��L�T����&|�0���'rў擪Xlĸ�K�xp� ��Q���d���i���nO�,Aւ�Bg8E���4D���,P&L�$���D�F��A��2D�� צ�=h�
%�΃pB��D
0��+�S�mnhh'L@34���� F@��`�'%�9����S>{���1"�`�����X�c�4�<q�N��tᇁց#���L�Ţ��ȓ<��͹��Q�:�M9�d�!4lm����@�gD)g�dP�D�6L�*}�'�a�<Iq���z[Nu�$O�v��{tf�\�<q���8<`�uK�:j}���	V�<)w"�6����W�4��ۺ�hO��`�'w($HAΘ�r�i��5�樣N<1�\���*9������'���>ً���$�T0w�@�ұެ>���wME��y�c+X��B%K�k����か�HO����$f�A�/ƾ����^�!�䅙#�Th���y�aЁ�G��Qk�O� S�W�,���Y2���(��yb ��g�Ac��V�ȇb���'F�z2f�'�*x���e��,Q�
��y���#W�9�l���.��g'�0>IM>)6%L�l�L����
X&�Qq�h�]�<Y�.Z8CG�q��i�*N�Ԁ')�Z�<	%/޽g�Bq{�D�2G"���A�<�1H��*�b��V�v9�}pw�	~�<�&U2'�젪 �&98�=��':��$.}R�'Ş� �M'%�8�*#��y"&���'�2-��Úe!j��2"��`q�)��'���Ǭ[%P�rݠ��V��
�*��Sh���Q�ڼ�*�!�8e�|�U�Yf�<AjV�4hĹ[ �G���<�W(�b�<	7�eyA��@"��@�R)�^�<I� N��q�D��qI8��0O�X̓��=� 4�3�	֡V����GQz�8�2�"O�Y�7���X�4�A�țq�$(@"O���� JbN)�F蕀�R�"O����HٮZ�������fH	��'�'����p�D�db���LX�̉��'Yb9���K',��rb�F��1 ۓ�~��lӶ�Óp�z���m�>
o�9�"Od�
%��h�� ��yUpL{q"O��Z5#��p�%��RFy���i����@E���Ch��5�3���x���^�$2}��iPK��xb�Q Y��$rp�?�!�$Z����Aa��v��푂쏣�!��NLR�[p锏Xf��U�"b!�$�O�@�B���l���KN"t߬=2��x��B����`E��L;�i`��/��Y��,D�tj1�� X�6`J/ŀZ��:R�6D�����}�FpS��i|����<�ش��Ih��x�O�,,���� �0���$!�bE��'!������ �H�2��!�Hq�'`� u��x��	ch�;��8˓��$/}R��u�.����	�,n��R��5�y��_0{/�d����
$5"��aM���O��:���yBl	1�u��0���~�<����$Z�T;f(Gܾp����}�<���v�&���EܭXfB�jx�<)QN��z7�d�GD�;�L j��w�<��@�ҶL�@R�I�=)�HS�o�x��ؖ'����#o+2��Yz rƸ�{2�'8ay���3��P I��q��`��y�f̵	����w'J66�Z<	POH��yBo�0T��[��ޟ4��p�P8��	p���OAla�Pi�E��	)�m�^A�${�'J-��#�F2&�{���V"PL��'>���i�0|����sk��P�����'���jvc�8i�j4@$i�(tcJ��J<�
�0g�@V-OQ�,8*BB�:w$�h���*��O�!�)Q6v��Q�NC߬L��"O�p����@�A� �'�����(}�Dv�O��0�/�Q,�@�b��
Xq��'.���qυ�J��5��-ȧz@H���'��� �H���tѰ��w[D�"�'�n�H���p�9`#D�V�s�'Oa§�#9�`�*q�-Q�i��F���<AUB7��	�F�R�B�1��eZ��̆�TB�I�*uhD�R���I���h@��yv@b� D{J|���
wW�j(ެ����DE�<G�ӟC*P�p���E^&�СJx}������ɼV��iq�$�
 0]9�ND��#?q��)ٕ3Jz}z�1h�Bh�Q�|�!��A-���*�F��0�4�q���J�Q� �'�Q�����T�axS���)��a�)D��q�(�.e7���σ4K����Ҍ�O��=	�N��,�=YB�����e�G�CB���.�}�<i1�u�J'	�{�>��\|�'J�s��)خ8�.��)ƿ��;FЌU��TΓ���0�4��H�:�a'	�wA^�3D��M����s��pU�[~u$���&>`�!�"O������1霤�� ά3g���"O"h�f�%:F혐ďV�����'u���4����iҊ�p�� ���`��-�FI�8��K�A�Aߊ��]$��G{���� �k � I��c#X�H0!�Dǿh�i�͍�j��s1`�7<!�$ڿF�v��@&��O�̻0�m�!�D�{�? ��rOW�C����9	 �	�Y�̅�I$;:�%B��xJ�	�s�B&)�C�I��G�s�(f$*͢C�I�3LKũ �$ [0+�Z�q"OD%@#H�,SI��/եw ���R"O��Sr���Z_� Q��ԇm��-J�"O^�YD���	�I[�̷C�X��r"O�k�BME���f�:cR��'"O� ��D���AD�	x�ݹ�"O�ekR��"Z&0B��-R�D	�4"O�u���'z-MJe	�#c��Z�"Ob$���\%�Ze�+M4�f"O~=�3�O���H�`�'Ts"O���R��l�E;�埑t���"O��� �rdᠤ�"rĭK�"O2	b��ϩ+��!�����<O!�K��|��L�6�1���x.!��  ,\�I6��U��F�#%�!�D�6'�R\	���ljTP� ��8�!�DP,r�fu�qR�o~*1{��[-w�!�"\�i����ш]eAA�!�d�+��Q�"աj��$��OC*!��؞{9dm��a�^8i�/���!��:*0�\�A�G�<+���V [?O�!��)	~�AE�
�}y �J��!�ć0�x�0� ܎_��i��Ѡa�!��L���go�)n��!�ElQ"x!�[�VG�U���;r	h��SlN��!�	���b�ٗ{���[6��{�!���" ����	�r��\�Jú<�!�$" �z@���ךFD.Y��,Ô	T!�$ّu�t�a���:���u�E	;!�DH&/sb8h2mה<�́y�jߗk1!��;
y^\C�Տ3��AҎ�)!�T�M0칂aFC	p��1�R���%	!�$��b���]�L$*	�	�� �1O49qR�@'���a�Ǫ)`�I���d	���H%�Bu-l�IB��"=�!��7�R��
A����ڲ*� !��^Qa*�����U�r�h�+��T!�D�%�D� MYc־�S�o9*!�䆸~��
���?j����U ��7 !�ڟ4HL�f�M8g�jd)�F�!���%�@�H���-{���`Hܠ2�!�d�[���#E�ȑ.Ү	���فm�!�{��S"��,�fls�]�-�!򄒉U-�ٹ1� �s�F(�ly!�$�

H�pˍT�4�P�׮:A!�$3}�����2Ja����X�L!��V�>]�i��̰b`)�A���X:!�P'd8̸T鍿_��2 {!�DR=s��ʶ�
KHE;!�Z.`!��	�(���PPk7!��xP�J-h!��,�Հ���/p�"��!�7P�!�DLG8�b ��f������ԭxi!����L�BK®ׄ,��_�F!��
pGj-��͎��(ӄ ݑG!�$[d�򐣀2X��03�A�-Y"!��&vvԩ��6t�`�w@X5b!��?n@�ѥ�Wob����	)!�$�/'��P #$E�\H���;X�!�Ҥi�N�f,w�T���"�!�D� �N�����H<� ��b!�de�TIK�)_Qh(��Ċ3�!�$��LI�@N��Y�a�'�n�!�� JD���D�ji�K���Xa�5���	4Z�J̠��ӁkVf����_{|����	�C䉍0+֨b���%nsJ<�s�H6G��D*w��P��D��)�5|F�x���-&-Ʃ�'$ש	���"!�c����&,¡�7dW�������
��y�~t£�G~w���'�����S�:�����'2X`@3J�,�:�%=����ņ5����d�R�2[4�; �K�/1\hHK?a�w� |[j��Ц/'ʾ�@+CD�$���8%��b��'E�,��&�x} �5(j2'���૒�ղ^THrQ�� %wZqʾ(\P5�u���82!zן�M���(.�H&�ȧ1td��놅d �)y��jܓݐ��d�2PF<�D�8]3&<;��I:JQP-DS�>(�鱫��2�&	���
�:�c���� �R#�1*$ ���<;$���K+0� ˨��9�1)X�i9��3�(ʨ����'����c�r��6��]%�%�T���֣8p�������ؒi�wJ���3�e�:	1�IO [
�ūw�D�:g�\i�h����(� �~!@ԁ#��d�0q�}2%�9lM�­nf�F�F`�t$�37)$���&��d�tHhFH�8lY�Ђ,mf�3n�f�|8�3��'��A�֜~#��x8�XbJ�W+l��a�`ܓ���P�U<����a��R
����$�,F��E P+��Q#�Y9S�.lN��
T��{�bݗ5���䙬F��y��3Q!�qA��	�i�z���I+Wg�Q��3O|}QM<����d��,��P-`\�0y�J<N�$I6�΢+��z6�A {-��BTꑗI�T��%��Ux,�wb(G�e���Ĝ���é:�+q�*�f���+�
��`�Ī#f,*1��	�(�!��r˄�b2 G [�|��나Qxhy��ȩ&h8�叅�2�I�G�t˘�"��!Vz�B�N� \��e�/9��8�g��y����ċ]^��#��Ur ��N= *�'p�+B�T>��L�B�W$�̼�e"�'qD�۱�M/t`}��M\#|�CB�=��|�R��
�ڴ�u"W<$uN�c��G=�h% e���W��D"ס�:3�b���-� U��`��|�MׁV� �UnL'w$�+#�%Cm�!���M"n���vƌ?G��Z���*�����^,ie��s�m�Cm�)��m�o�ղF�G�
�t���5�@$;m^�I#���W���uVOB(Ae�����JF�	fc��+a�DR��8Y1�+n� D�U'g��\_p�X#CˏJRn�4�U�g��hq�/	�49�ȰT%C�ZA֋J�t���x��NXx�i��%!$`��Se��<��|S�,	N��MC�G9\��s�J�d�|��Ī�4%#l���Q�8��\f֋H��yr�F�[�.8(b�@8y�8�B��9�p�� b ���K��f� A���@�_�6P��:}�6�O4��%ƼpdX�ÂD���I �&R�{Yb�s7��9%T���_Rl$m��E>uzl�â���q@%��zZj��%�j��#�JN
4�|x�Ǎ�L_�P����&��`(�2'�� �I�1u�H�T%Nu�De�����4� m�&y�i��K��]��N2�tU�g��q�PU��~�Y��L�6\��)+ d��P]�ѣvdʪ}�*�rQ�G�8{�i��|B���:~�u�R$�>lH���W�B,z;<ʰpqR���"���'*@I��8�_{+h�lĶ|��J�%�+I�M�����V�\\���ߨV"ݓ�DY/tSE,E4y���ɖON�� 1)�Kݎ��,r�p�L���<��.g�6�T>��)P�c��騡-Ay��٦�N�cI���ǥk+��I�3*^`�� 2FD�;zR��ӓHX%>��A���#`A���E�}�/H�0���;"�ֱSv�l��A�������c2(�9`]�����S���pȮl���4@�$��b�'��I�eQ%��<�qʊ<:��*�*Lf[�AB��Y�Ek�Ċ�F�(U�����*)��I��N)n�H<��H�O�P�J��h6�J� ���B��ء?�.�yu�݋b��a�	�~�P���|�����.x��dʧ��z��Ǘ]�lI�䯙�w���o�#��uΙ !�7A����\m���#�3K@TCdII�2�:����8:� d%��n���i�$��t�8yz!���5�дѢMS�M��味�W�:��ٛ2R�M��޸<s��R��>��[ �1@ģ�Gf��� 
:2��|�5�A4
�0����[�hJ�Z�- �}B��o�X��7���м��퉟�j�����x�h�Z!��\Ֆ��aY����ꅵl&pUK�G�Y�ט}��@�✽2(��T�O�h��&�J�a%���"�		v��d�P&R:oR�q��ğ@�1$� =��	┈D5* \����4�~2ЧF!�I)���n���8��^�M2�Bۖ ,�A�F<�\��E�p �g֤VfJ����� HϮL�֠���	s<��$>�1��H/�b$�'�29�x�3w�\�M�<���ID�}��<�C��q��1�$����L��G.�8�1�F��W�i�H=�	A	\	�"� u�-R�*�d����'�
t�G��B�B!Q���D L�B� ן:4��`�$�Ye��>U#<��a� ��I�f��TN�C�S:*�2�ʟh� �Qu�dڤ2�x��ᚍA�J�i=/�ࠍFz�� ���/���������?��[�E�\�i��,����Fx���%[ ;ȭ3'D$j��ɘ�%?y[��C�<�I7p$��jOM��ѣak؟��7oM�_+"��S�?��Ĉ��|��BR.=�s	P�F����g�^-.�	�4'q ����Ҽ�G��w#�	�p�4!��!�T*�Q~¡�kEY���'��� �~�H��xM�e�񢈐.:�ЧŪ[�j|A0�4�2�Ñ
xR�n��l&�ԈӠF$U` 2��T�jC[�17�0��3���R *]�- r�R�+߭-.�9Z�I)�؉���5��Śr!1���
Њ(*b�r���J��i��\����t�9`5D���Za`�g�;����RD�����'y��=�ám�����XMD�p2g�,�Őf���5�H`�dU#z���hM#� D]%����ƒ=���0Q,G�q	N\���$�h����Ē*`�&�e�'Z���n_0D���Km�|qc��
]͜�K��F�5d���垞I�*��Ŭٺ6Bv`A�a:{X������YŐ�C�D��1p���_�y7Lޡ	�3-�<,��I��Š��$��{_����D��Da�Rb��m+
�Y�����Ar5��X�-A� UথN\&P�X���1�N<8����Qj��Fl��,��ܠDm�j'�ӿ&&�+�M�:B]�!D&�+u.�SR�=@�ԉst��Fh�RW@��$%��]�EQ�%*�ǲib��j5�C3GB%���S0`��暯P�" �đy�:�?�Al[t�
��sD"-"=�Qg�*/���x����:O���bR zα�r�v���sH#%:9�A睨)���8�)Q�9n���#0!��-cd�"3ш�"�Y�m�'�����B����5���Bi���aʨW���s�jɱM8��FM����eIɼ0��۴�h�������)U��� *��o߱1&t$*��?Vд�%�>At��}��u��N U��f�$�i� T���A�,�����. ���၎:_���ٹZ�<YA��[=���u�K�.����Վ�U�o�b=Ҥ7X���83�֌	�|�v�� Ol`���'n��a�f18�D5\�� ����p��/��32Lw]HS�22�1�%e����Ƈ0�(íѣ��<U�I�� �Q��*=ʗ*EY|ȹ%.I$Og�������v��^�d�$� +Z�� ��F^pܙn	���Z�T6���Ԯ�84��i��ɍ(50��%���c�H��p����(EshĽ�ЪM�r��(QW���^�)g�]����[��̐r��ѱHp`֕��l�m�5�оU�`	��+-(�i,*�O��s��0)�j�`T��+q���@W(k�ة� �R�l����\�o6�9�2j
�)	��	�ʗ�=��ѻ�"*����J<�V5a�  !�iҐwwQ�%�d�'��(�DF�h��aP��''��<�&�J�L�d�$ٶ8T,��oȁ�^�r���GE�M�c!�1*��<�1	E)u����Ŋc`���ሜQH���mWTvT��a�/��Y���-�`���	ip���A(}"�O�:�ȳ�/Q=1O��{ୁZn�P��g�=z����=V`aR��A�\%��C������� �rTot�~0���>v��B"�Z@��r��<$��
�4+Z�0s�C�N�݃$	² ������y�*a��]�TaX�ȥ�ٸz0�	����P�A`��ː]����g�C@{
e���$zb%	,@���[΢8���Jg�>a@/
�Ti�d�B�*$�A���w�	d��xf���.KF��A
e����X�g���2�~�,e�p��>i*��gF�!�� �׏��b��v�/Ul�
rL,��}�^)0����H4�I.A�Ҭ�'���ظ!N��G���"ti�y�N5 ��A�
4 ���G�̔���i�Ɲ��k>�p���4V��y`�}�x��	�Q���&횦֡�FiS�P*�)K��oӪEJ��ܹi�6�q5�0V�� �&mۤƁ��R/�5e�
�s>�RD*A�CF����AL6}K���!!�VY��F�=#�~����/-\\�)!�@^���PS��+�Bܢre�8���^4���AE�/ZL�y�M�[���xc�Q��R�d�6EU���ߥD� ��3M>E+����5{�N'�8���.S��%���3V��1��&&+��Ʉ�^=V�5"�#F4zNdJ"�Id��+���"0rd��A'%#ўT�0�"E�hD�X��V� A��$$@N�B����`�"
�i��H��F�x���F(������"�養�.�0)@6�YMH� A��K�J��r���0>	u��6x�B��ݠ������
���[�^�{�g�Y��`	WL|��c@պ��06����@0EĆ�?J��DI�����D�f��˓ ��p��Po$�8�oH�u�8�yddʪ-C��QG�!)�V�葉�FF�����P	tn4��IĎ�6�QdK((N���G�+�P��	�ݦu[��ϳ9��7���J�P��"�D�$��
�R�i��)����l|�B*g*y�����O�R��kJ',�d���D�T���n���h���K4��q"�)M�X�)��	r�՚�+d� E��YZdh8�G��N���!1���Q����e�F�y���􋍝j�(%�ލ^W`d ��ۂ�m��Ԩ<�]['O�GD P�P4hB��	�r��ՠ��d�N5 �	:7���"[�\,�qv)ԁ'��3 A;=!������f�D1�i�7���"�Y'�<bHU�F�DzĮ�AY6��2�'2�����?��\0!%C�C*������d�pM�a�ιۆg �_Ĕ@�!IԀ�n9v��48c��-;>�"��2Zɲ�#MN�2�%��%�t�92"M�sx���Bj�	��6�"��QP��901DB�	.�5�tp�Kt\l �@U�2�F8%�Ո1�Mb��Fex���UNH�@C��&BxD\XA�x���"�E
5lA�˘)��!Ǚ�+JP� ���(����a@������9ziȒ��+	��Q� #�l�^F(L��N���R�\4&�< 0�E$lOH�djx>q�sC{�D��%A�9(�L����>:*萷-���.�\0�'�:0>�_wjxQ�E.�7����0D�r�)����"�p���џ��.����֮s�B$h��ѹM�����v�Y�ܱQ�8; DJ�>R��0��T��)k�m2�u���55ZԁWf��w�Py��'�8:t#��3�5ɇ,R�HA:]��O��̓d�I*�I��D	�!��
���Ѥ!���R����Vt=H2hK�����1������ "�L���y	�6-WZM�b���~@�r�N4ݜ�� ��
5hn%(�X��(N�F��+׃R}P��v�դ�8�� 	w5B�:�&�5U��Vǁi�a��@����iEm5|O��͓\ԕ���O������t��nںyh�ڗ}�Q�c�[��{���x"��W�=�<֝�?	r�#�4mp�L��S5q����4�'?6E�'̔~h8E;g����@J��Sck"��Ò80�Ψs��w_Z�A&F��5:�C��M�BB:YW�Ě`k ����81�ʠkT�tWH��fB_�.�!�����h���66Y*��ҡ�T���R2]ce�[�>5���M�|�`��r��bA	/c��jT�;^�}Rw�#�%g�� G�d����P%q���q�u �R��9Z� Y���"$/D�V�AP�r��P�?�:�թeN\x�F�f~|�c�ȣ&*N�
�O�v��XwW�|hr�����E�-�&ā@T��W��S�o��J��(`���F�������9;�,��B_�h2�����[�ZU� /!>N|)��k��A�e�Ԇ�<,�@�C2���6�6Z�P]��o"?NDAԣ�h��{��,I�r�3%2�a@5�ɵ�j)jwB]�8����ˡ=j,h�0� t$��5�D�&��jw	�MZ�Ѓ��س_Q\���"Z)tҖ䪔%H<����Ņ%��*�ȬN^�ؓ��3]Vv�:�&ʫA'���T�O�V.NA0�Hǭah��R��N�K-�@9UBU4�h�Z�(G+��"U&\i`SHF/`hra�$o�*m�"�h��	����d��O����V�.ִ����KJzi�4/�o�2�8�K�I���/ޝ	SD�8��@�r&$�P���/O/�l�S0���O�y�1��{��x��
� 8d
��7^��7j���0e��{�y�!n�%�F�#��ڍVk�%�\���c�LǉF�y��r�A�<�6��A�@��C�H�V��DɎ��2�_+w ��#�](>�.7-�R�{N#��"+9�6�)EAI�b�ԉ �0z���W����> &� ͒1#��������F�iJ8��r�? �L�d���(qx���N��oc���p�K�NaȈ"G�i����֦�
\�d��& /~f����kd���Xw>���&�*dX �%L7A�pavm�n����D1]/�\S4@	�b޴�A&�.lH �E����M�rL�#5�D@'͇�8Y5cq��Ñ�z�@p���Q?8�iG�и�x GM�?1Ae�t�
O�K �	�6�`���D1�ih���� J
�x1�Ҏ î@�#�q��+�䀋�,�8PL
�M� � }��@��L�8)�b˘*�qk���!#�ġ�!��,�������7��'k��C���<W)��(CL� �کRSEG)K	S��y@ܩ3[j� ����.=��8eM̒�΁���'<�b#�V��! �I�XF@X�r-��5f�P�@2��R�F������%Z�Ef���D��!�b4� �(��#N��Xޙ1�I8�D��rIY�6� ժU�$E����	,��0sn��\΅�d��|�B)�:V�9k9b��Aӷ"�8=:"�sܲU�.���4/���һV�1{,b�U��4w���q����`��D�!�kJw��%BA�@Tn8HA��F���!���#��S@�a�y2C
<98K�
>���ɗ'^�4lؕ�e^�̥���~|�[�46�Ի�CA�~�ɺ4j҅ء�W�0%@J8Ђ�P����` �˲e�qB�g��,j#>!v��pIjYYG��� �M!~���s�N���bdX;���_�` �lI�!��y��fоVk�%[wȄ�{=4jx����o4<�3a�=}Q��K��W(8IR�ÿ�"��G!�����WM�
P�E��ͻN]ر��>OF��M��/	Ҩ�%]*.똘�wmd�u{4E6�O�f�`�(,��Q�/{.���'�ZD� ۡ,1Vd[6�	�t�bY�˅4o
��CŶd�lQ�n���3��"a�Du��AU�.�J! �mD/���$�"`�@�!�9{�]��Ε�;��;A�"�HԀ�g����>�R�)Z�����ֈSDU[F��M�<9�앬U�R���ѣ,Xx��KLL�<��R	wm7�\�b�(#HPJ�<��]9{�rDIqH�p.:�҄*L�<�ˮ_ul8*�
�wd�9b�Eg�<��
�2��{�Ғ_S���^O�<�4oG4N��hg
�3l*0�E�F�<����x�4`J��ڏD�`X���}�<�Ү��8V��E��h����6�\@�<�i�`~)zN�?oiQӷ��D�<���K_��x�E�B�`�3Rə[�<�D� @��y*�F	+	������|�<9$�^0�� �,���Q�c/M�<��J 1yq0] �#�)L����b�<�X���('S�}��@O\�<Y���> OR�`�a�`|,�b`Mg�<I6��m�8H����r_�!�Sh�T�<Auh��#���
2戈y�HY�Νo�<�C刌��ȳFE.D�����6D�|��`V=.[܍3ܯy�9#�(D�d6�Z�R`�g㟂]�ډ��+D�H����+h�v �m�Y�hp�v�:D�(�)�)xs�;�L��6���b!!;D���N��~yM�RL��J�~���9D�p�����|�8��]9�"��rO9D�l)2�H.���4��1c5D��+!J�&7�,C-�#3Ѣ-q$J=D�����٭<C���g�:��y���8D��C7,x�A0��6�!�#�-D���'M)*Qa'gP_yV�G'D�dZ���<{��Q3��c�*�Cn#D���`U�Q�xyG�2Uݦ|c�o3D� Ӱ$��4��USu/����1Q�j3D�(0�M'q�D�r�JCP�ɨ�#D�Dۧ%.!�1 bZ>?��x�!#D�\s`���=W,�#�j�t-K�@!D�8��ÎH���
�nN0R�P��%D�HP �s�����9[-�ܒuL"D�����_=L�P�V��k��=�$m D�4�$�pU� `^"6.m�T*2D�d��P=&kl	�GD߆Z��(��@/D�d���'t��A�X3���)V}!���$>&�y(���h+L�b��<MP!��@�Q:R�	�-�< �Qs�٬U)!�D��G����&!Q�!*AG�<,!�� 0��S��D(��1(Z�M�!"O�d3�a�=r.�EHch��`�0"OB�a�"%����=��C�"O�5˷&AJ��\j���
$y�4D"O
<�IB:�$Ah�ƒ(:oVuj���.� ��@ᓥj9�}!���u�B5l����C�	&3����q�ԳZ���3#��q. ��ۨ�H1�5����)�'o�8�DƟ�401��H�YO@0�"�		��u�549��ȴXN�'J%����t�f
W�y�˓R20p�eۨ^��h�,�-a��؈b&̸z���	�,�"��'슉(v�+:�H���-�)��p4 �@�$@_�)s"��8����e�\Fq"@ra�˿G��y�ϓFp&Hbq��>���:/�>���D2���3�	f��.�	�H,�o؟;�4�����)�$���O��ع�)����s�����lR0W0�ч�Ǎb�qO���⃆1Q�j���e��q���O�/;du��8_����qi�rL���J��+f�=�!�����@7 <N�<��R�������q	F壴j�~��D8Y���������$h� M�Å�xZܴ�شw��K��-�������Acᙜr�D Ô�\�	s���n���g�
��zCA� 0�R�ѧ�/R^-i�Z/2&-2c�՟o��ŧ�R�vX*�Iq�G�ЬZ�Mǚh�P4���0i�*�b�9Q�DS<�IQ���D�ްZ��d�4xteC�t� T�2��8C���h�	��W�@s~4[�^2�z�$�o�_5d�h7�L!m�PRv��<D׸��R�ŖQ���@���b�@�CT[�-�L|)%�蜣v�̱M �5��-��} ��ru�:kd�0��b_�.���$�nVج
tF��P�O��yE��!��	�P"p����͋P�Լ	�
�*L,I�Q=<���ꇕK�ȱa ֠R�h	��xl�T�]?x9ZU���V2$��A�FI�̽AP�!Q�d�v�ŤW��C� ����t�U�N�jLB`��ιT4����Z�椙֤%}P�#a�Đ��L����mD\\�p.�K<੐���*<l@�㗕�:����C$�r#�P4fi� .�
O,�� � �d
b��a!#�O��=�t�V`�J�P��2��	��͝�K�rp6De��UQ��I��	�䬗a�H�X���zR�R���u;���ž/�L��T+S�jC�#T�On*gC%J؛r�sN��*� p� ��K�AG2 �4gW��
  7��&�� q�d��Nsz��*� q��p�ˍEL<0�$�W�,�FZ�Fu�ذ�$�d%j=�Rf�@�ɜo�D�*���ޜas�(N��ء�ů\ڰ:-ص2�9n��=������Ű(�k�C��<���hߏXJ0�ҭP�&2�Q�N��8���堅1+�!�a��0ms�<X�Q:U%K�IY���I׊�i6��f�JY�b��/��H��M�`}�@��U�(H0Q��H�Mޒ��M��T��8�
'%�!cVa	�ܘk�ȏ	�ez��Q3e��A �H2R���xњ|��c�h�2Ƈ1!�b��d��+�hG�)�r\P�'7�Piv���c�~4�¨G�1 k��(X��c��أlYR4i8IޠUɖ���3����aV$A����t�n<��<�D��m,�{�C��rY:���qb���ͯb�I�`��8	&���Vn;��
�ц	�ۀ��wb��7���b��&���F��K�ɉ0�D{�@�g���OLcD�9d�Ԩ�(��'�� 3��4F�k�(��F���"�����q��>B}���Q�I,F�|`i�o�$���.����ƕ��a��_>Cy�����ȮC�f��b��\l�b*\��ȑ��*J���$�Ƚmצ=���?p��86
N}����4S
����z�<��-Wk3�q�Îj�bu��	[�f�V�=��јv���&���}���"-�@�@��5�h*Q��T(�%��oD)��` c@��L�R>��p��L.8��#
D>GQ�i�%� 4J�q
�D�h�,�xcD�CP�)z�ڧAMb�8���e�킰M�gUQ6h�0[�]�D I�	� ��L���	P1R��"�R��"O� @#����O�9��ް/�\�r����=/��CH���ՀY$(|P+נ"2���� Ö!n]yw��19���dn[�S�Mzw�חr�:�[�L�1 �ݧv�jQ�}�"�:@��6�
�e�Z�j�K-&q���vDxq���nE.w��j�4Ն���/��X�й��N@�[N�ҧ�{�dG;����ֶE��t`�F��#Ep�����uduc�H�pe��i��Ǌ8��O�<���s�$M�o�|ݚ�W��>H�y�+Ӗd��yɧ-�?qj�LY�ի��߶d��I�!o%-)'�@� >��h��Z���a!G�M�'bP���-�>��En�jD�7�]?3t�@�"q�� �T�>�H���H�U۰�2�OH�	✜FGإږMT:�|�����f+��!4D��o�N�ݔJ	d8�˘ F�e��Ǐm���$����F���"����'<�=���S�n�m�Cl�~������M&l�QG��=Ĵi���ݞJ7�|(�!vd�u�s,;�Stf�7���v��1�6�U�w�fLpw��>y�	w��2m�\�$�u0����.�u�����T+t�jHP��-a�iL���)�be�b�hCM��q��"(T�i���8�!�.���㟌2bЫ|6���B�Kb�\�g�Dǈ�����+jY&�ٴ�ȷ}�D@�`�'.��&%��Id�\�WČ�����}6J�2W�>M�4!�k܄Hz�D�cT(�t�?�3�/dt�8	򨖺��`��r�씳3k��\�(���5A�	7��O`\P0lč�xS��͑p�愫��B�m)���w���7�D[���h�X�8�3�O4�ɳ���
YX��T�$�O-f)ڠ��/F��y�P���|��K�����+�%K8Hځl��M�	ձw�~���ɆJ<���D;tLZE��4�~��Ҳ)�Ѣ%!��,X�&��:BY�[bfe0@;�.Ұ"��ʕa���0l��h �7- �Mr��54=0�D[�:T��#�$}*q�@pI�]j�� �hO������"l>̹��Е�7��>s�!�j"����~���;鑠d*ة�[�ڵ��X�w�:1�D�r�8�34Rt����ʥ3�N�?��n9L7�1�׋ߒ.���*��1���/˕(�a��_Ox��1��;��L�� �6mиm��$F�:
�����*�A��͚�[Gv�λR;���s؄6����&,Z�x��]�'oyq��6���ԊG�z�O��K��4<x��1��W21��L�J���`�J4C�eRN�L�܄Y��ҳ���u��Ȉ&m�'�0-�����irc�3�b��%mR I�}  �'6�-��8\�6=�pD]��qB#�1�v��eM��� X���(W,��	Ǩ_�D��a���Y�%�X�`�r��-�4���LV7(T�l�Ǎ�_�Z�h�aA)o�v]��Eɥ@z���˅W��V�4)T�xJ$'�[�L� e�+k�|Q����K�Pm�
I�w���0<IBg��T�RH�ը�I'|扞J;�0x�M\��ᛑi�5S8���CLe��E!�ؽ�,l��E�O1�H�-���탡�ô}V2�]+.��� 
ր1���a���6�'bR!��BϧE.�yH��|�'����g�<n4���Ը���y�6�#��*vɚ� ���:{.��l?h>�"�����'؎���O���4)�"M,:��Y�MX�rL�P�'������1�3AE�4Eڔp@J�-i�y�#�u�3V��/(��,����WuPl�Ч޺`-����NN3O����ލP�(I�.Qz�80��5~\�e�J�̀g��6�u���ďT�8y��y� �Oڴ}V� E��[�HZP��vU
�ڟ#�����G�ų�O�q�ɪ h�Y�-�]�����Y%
���Z��fݲ�0����m��(�+h�I��[	T���a?�4 �/z�l��E�\ıg�' bx	�.\�O��-S:B�t�ÈC�-N�D�tBL��<ɱd�>�&0���4M"ʤ�w��?H�@��³)I�'�,��1凐k,���u��
Qɶ8���Y�f�zM���
%�@t�kݥ��Y�V\<��Y�ǳ+�e��/+6 �T�
�Awd�����l�� �pX�H���2ͪ����+Y���%�z����LJ
k�ޝzA��iWj}�GMߏ1Ȭ��O����[=~�h�BPK١C"�YKd�8W:��w�6�P�&�
p�ʐ�@�Z�<���Q���i���x�l����m7r9lh��W�픑I%�շ0~(XCG#���93Ac�����gKJ��]؞h� I\1f�H�fك �����B*���p-[M���HR��B�$4�bIվ}���ۋ!���C� /��1� �[W���5>\�U�l��X/fixcȃ�3O�O�� ���\��!�m�r����#N� !�ϗ6ja ��(��U8�J�6�8�H��W���L�,�%�daI����OT5�b��5g���JB
'8� ۗ앒$�<3��ى4�(�H�ȳx�DY���14e��0SjÈ"5��w,�Ѧ�AvFϦX��݉5�P5�v��6!��ed�d���'� �)��V��BA�P�;Z)Ա��S�v�y )Ֆ�|��E�\�|�:�i W� �Ri��(G9Y,ޥ�_cx�)��X$����F�I�r!�6�?lO��SIӬ!ݜ�/?p��(�*��X_�a#���&��I�6�t�����7��l��҉�>�0��,\U�9��
�� ��A��ϟ��P��!5�e�g�M�x�dIf�5��2\�y*&B�g��,�Ǎ�4u�QPC�X'Sb:@8��z����Ī֓*��RV�&d�G�I�I�|���*���(��By�ў�Ԅz�ȼ��2�zt���0KJ8E��ˍ��z<k�NG%HP�,���y�δ��3�n\�T��0JE:Y�!�V�/d|�"b�ɜP� �t&�(x��F����>9ħ� g�����Bt8Ҭ�Gv�0殘!���q�D!� �xD���e�������Bp8������M q�|���� �2�{��L��`�üd����G$��@ b�1SB_�v�����p]]:dBV�4(�:��>i6РCg�Q$@!h�q�"+p������8q^Q4�ip89��Ɏ2�j��1���������?��dZ ��d�4��ucC�94�SϦ�dRa㏨z���ڲ�%a܁
��	%6�_`�2�'dƽbp��3��FzB/!=#�٧AM�.7��/\�{����|Ќ�R� ~�ֹӗ��#8+��ǡ�	-1�	��oݻ~��8�n^n�!`S�6�ѢI^�~�,���/2���88�Eia� 34���^+ ���#1���$C��%���j��:3�a!�ρ�<�)��ޫ"���?V�JWc�f�:���!��M|2��Ԥ&E��gN.d{�ɱ4�B�KJx`J� mӪɡu��=��x����I�������Y����۴P���[�5s���FƷQu���Ik"���qmU�z�68 �@_�p�6U8j�R�޴��*��@��J�i��~-Y�l�	|��I��^�v�"�=QF�<�P��І9��� fUo�h�X](�JW�3|��Y�A(�,��&��6�`js'\GﾈÐ��D�pr@-? n�!t�9ZH���w�dQ;ӂR'S��82�ԑ�z Qg�V41(&]R��
%LV-)��F�r�raS#"S$V��� �t݁��w3��Z �Z�!`ď�d̚a��'X��U�L�!���1�X�p��Q��_mޠRB 
���a������u��( ��ȱ�ٜu�$�� ft�5M�O"���&4-FyrbS�dv�Q�y򯖓$09:F��-�h�aF g�*��d�Q�j�:�2 |4 Ƭ)I=	�f��(�>)p��
)��Ѓ�+Uܙ���5J��r�ʽYR<�Rq�`�\��)�Ě�/ז�J`Y�'��`�m�&I+�Ս~��A�C;1�2���4�p?90	V��"1�֏Ƀ
;�3���������E��=i��F?s)��b�`S�;�q
d��x�kBm���u&t �(�P��E+��8K���>Qwb�A� A 5i\5`������v! p��M�P�ic�� �4�� E�03�@I��[42W�ChN�BZ08H�Í�Q�msӥ�5��8�eC59ڨP�Ԣ5�$�J��N!}H��OH%Jc,�0 ����$�QgI
���ՠ1�4+�*N#qP&�A
DB���韴&����F�(��,�U�����}R�YZbx���M�XM���鞶"��%��'�R�X�" m8�cSH�E<`�ă/
V�p!�<�M+3Bȇ�x� `>}���P�7+�XX��V�.j��9u'�?K��b1�� &�ٳ�Qs��d��'�	���D�`DF��L�8D��6ac�l�d�R,^t�-qGA�<a�Us��L%L0���gvV=��_7bc�d℠S/_u����5�fg\�pS��U�y��y!�[[�'-"d[��̆Ǩ ���(=��#"�50��`h⣜�
t(f��9;���C�T"5΁ � �`���(��;�^�i��xx���;?��V��Sb��w��q���Ѕ�+8ʔ�!e$̼o|E1g��Yr���#���PA���w����E���;Ϝ��M�jvm)g)װN^΍0��	)��d��sWv%�T�d��9q`�8GR\{�W0N_ʁ��@� $�� $�1#_�S�^P1��'7S�D�>�MHK��Fu��۱7N0�x�C�U�DxZ��%0_�%s�Ï9�9�B�E1H�-a!	$2������*�JDA3䞑P&�xr�JI�H/�����V�u���̞�H��G��\:�0�`o�����D��r��u�U �'ܴ��4��u�\>	�x  !��2ў�k�mA3Y]8��Ǵs���'T�(�b���ʵ�~I���[��<����ΝU��TplW?sRЌPr�[�D��ɇO��C��W�͈%���x,�}�ؔ{4�>vZΰ(��C�����;B�.�6�����LD��u�G��qy����h�PH�pN�%tp��8�'(����&LE��e
ק��tr���2��hv0IC�A]�1�^�a2L_o����R�b�P��!�챘&O�/Is6A��0�P�1��>��[3v�|qH$�_0|��KԹ��!S�E������(J�^�CP��1p�jY $K�Z;d���4s,M6n�\*�[棋,[�$�3%�X�h<�%B�=c1���oC�P��-3�}BoԬb�\��$'�
�8�!�M�`�:U/Ҽ\��!�sH����A���S�,���H"8��ء�L�n�B�/ӾX��	�Co�38�&2}���bU@ʝ���	�ptn<0�bL&`�hݛ�� :��7GƂF!Y1'A"�`CW�%�~���dL�r�Q�K�1v�*`!�φ+FҰq�A� �r4��C&�x��'q�	�TLۓ	ک� �]�8�Fm���ڰNƼ)��@]�	%���o�+��D[���]�w���+��h�6SbcΉ+Lzy�&�?'n����� =��BdW&am8�;R�G��@�Ar3�xq2���}̓l������"�� T���(=�'64a7�Y!���gi�So��P�Q}b�D�IȢ�� �(�8d�W��F��Vg�Y���B�B�~M܁Q ��O�d�S+�-��ׅ.t�@!ӯq�4��D�(tQ�r!�`2˓�f��A˄;Z�锋8)K"9�wu����;P
����%Z����d >Q���ۈ�i�<�:mqW���Cd�(+�C82p�S�v B� 4��3<N�S�0=�8�R8
�����do��
�c�M(7� ��@A �y���G�H!���p����u���,Qh�̔"J���'+�;\T���O?㟬�B�X�>�TXx�Z>4�I� �:�O���b�X"�T٫g���|A��I��
oB!��lս{���	� P�i��!ܥ/7����OA�o�6���F����3ȕ�@�B�2�iܿ~Zzчȓ%����|E@�`4��ifT��odY¦C�tQ��!�R�[U(��ȓS��� ��	ZZ4٫"�ՠ�pH�ȓ5ʛ.0�
�1�qapl�ȓ"$�T��+\|̹ ţҥh�ʕ�ȓ%a��&Q�L��XV*��$w� �ȓM�V�As�ϲ�.$ �ꑷ ���@>�9#�E*a;��R^��E��/̌(�G�mɎ�ö�J�*����P�X>�TA[��	��ȓ=�,�3��ɔNʾ`KF��5��!�ȓn3hTq4�]#&� ��ÆH�0�:���4nDxS3NZ
))�ԀDf:Du�0��0�@�c�R�I�,J"�Ļ	x.)��k^ |1�B
 	�U؂���b�����,�(�:��8V�*$p�)�3.H|�ȓnX�(�rl�f\,���) �l%��;�T�j�X=z�(� 䓘�*��ȓn�(�  5eBgB�G�Jm�<9凃@�TQ��k�>�(��e�G��"!$ٶE�~dY��Ua	�Fy��ΫF��*1�d&$X����^�6Q�WO��3��IN>�Go�3�����3g\��֡��~�:�a(E7�<Yd�^#3f^��Ɓ2����XAh������>�B`AJA��}ā�>%>Y�Vi�8\mjt:��К�Ś7�$_!�(O��2iV)�eB �21#�m �Z�,��)ҧyAQ�D�J�VĢ�@^.W��Ҁ�Q���'�X�𩊑W1�鐵F��p��pP�×�W��➬��k�+ɨ�����O*A��Qv�5S�d���F���k�����+�fra��L:H��h c_1H���"�G����dC�+��E���W�?�� ���HO�q���ݏr1 �Rs'��UU�����Y'X	#0�)�'rdp%;6n�b�Cg��d�m�	2�'�i����[c��Y�(�@v-FCTpu�<If-�CUr��i�>B��j�mP5~{X��	�u��'ԛ��MIR���	`�
����N������M�$)��J~~"I_�6�MZشQ��>���\��W/�&	����6ˉ6F2�+хQ�y�m�0�	ڟlקȟDICt�xo��#�{�����;��%2e)G<��#wa�Tʦ.<�sE�^�n�����D�h�J<y'j	�1a��C�r�½s��v�VbY� $��C� 	�bX���S|g�� �C ��^�"�m��of�˓�r!�6��S�π  ���l/��P�ǀ�@�N���'�4�`iO�x�O�>A���zRt�R��&&	R�[�i���Eo�n�S�O����1�T�*�	(�jP�w���C�K���'�R��I�A�(ey� �<v8�F��5/f���W ��cA�c�)���� �`C1�v5�0�tP.L�ȓaR� I�)K�Ĭ��-���4��*+�K�E׈Zz���u!�akȇ�^�����1O�eb����{9�C剗+a�fN�,�(�{�@�
|hC䉃��Q�1l��m�\]�cc�g�B��=gP@��@6�9���J4'!B䉕,�h�G�D�'�	��B6f�C�.���y!�W�@����!�/Z��C�I	��8��/+����e/�#Tt�C�	�J�J���:
*R͛G\�j�8C�	����Ft��o�=b�EZ$+5D��j��֌�X����L�����-D�h�`�����X`���\Ȓ�re*D����1}������f| �6K*D�x��'�	{C��aB'ܝ^�ht��f"D��A��=6��i�G˘� O^�@�-!D���vf,uX�����e�t�3i=D�Xq�GYn�d�XgNmQq��C&D�ܙc�LT>زģ�4Au�`��$D�d�7j��J!Gd;&�d�@"D���@D#_x(�#M�;����ĩ2D���mF�/� ��7?��p�7�3D��A��V#RrMڰ�W�H�A!��1D�0aU��-y�V�Sdϔ�7����1D���'i�fE��eM%xL؉ef0D�Tˠ�/R��L�'X*�,-;D��x*��l��`,93�$bR�5D��`���hۜ�"���<<�B�:�H8D��A�|@YڵŽ.Y�a�2D�(�B�.�
�)�� i�,�`�0D��q���+����Ԍ����a�E.D�d��K� x��R$ę����d�,D�DIb���1+�g���Y��5D��K�.Z6� ��A���+�C8D��5B�!B�F��Q��9v~��s"9D��"��W3�Q�m�]r~�8�6D�<�0�ęCQ�P�&�L0b�ɳ�&D���%B�_����s�	q�I�f8D�X�3�Ig ��Y@�D�3�m��k+D��pGFGu	.��4�µ`/�]��J)D�d���E�Dh"�`� Z|u3ѥ(D���rJJ�P��xK����:�tI'D�\�0I/� �!Ă�����'D�X	��8�]	8%lJ�Rq�&D��@t�S6����5k7L\�E%D�X���U�!�R�)�Ω�tЉ'D��TDƾ�.t�����d�l�1e$D���H�2İ�T��i�D ���-D�x6#�j1�ɢ�Ǧ#]<�' +D�@zU%��hFg�/p>UR�%)D���E��Z��y�r�Ơ,[>���&D�؀���`'.]a��7r{,v�?D���V�V�%J�
�-�$�?D��ʔ��,p3��$*\*�鄠!D�HK�O�X̠ B$m\ͪ�e*D�4!'�J�*	pMy��^�1���N)D�����ô#��t�Sa�%��c3�<D���H�>�T)�R��*[��u�Ek;D��c�(Q :�"A([�����n>D�� ~��ֈ�,W�M�l�'�R\!�"O��۔��U���$�޻u���j"O�L�h�c�<�9ժҌ\��Q�"O
T{ã���]����8�̚u"Om CL@�j�8t�QhP%���Af"O�ɚ 
3e M�燔k�� ��"Om���Q#gn���,	�*$y!`"O����E�K�4��ǝA@���"O�Ċ�"G��4`��R��q"O`�HCN�OBHt���ƀ)v¼C0"O�L�I�p[܈:ah��vJ��{�"O*Z�[7��hZ���\����P"O8-3�	G�@��gaC�&�8�1"O�ı���:���yt�܄�ŉ"O��#����I��.rF�,rQ"O�9��M�I' TP2<�R""O�5C��4��I$J�,L���q�"O��zq��9�&EуI�\���"OXq2s�Ҋ��b�aR�hn K"O-�efC�l�����.B��)1�"O��H�B
Pcy����)]��g"O�P�c�:{�9��'D,��a9W"O��7��8��X0u�T�p��T1�'/rX
`F 9$�"N�A[؄�
�'����]8jǴ][�]'$|��@�'��B�4%ٱ@Ü�V^%�
�'٤��VEC�n�ԛ�'F��%�
�'z�U�`�)/����"	�4i����'��rL���hX�j�Bl1��'R`z�)Z�G�QX' M�=�f��'�l<g��,/��G�,3.�T
�')�Eq�	(٩�V�-�`e��'��i�KL9��i��̋R�h B
�'�Ɖ�*V�RwhH[ �߂Wz-@�'�2U���X� �(��з|` �ORL�<Ac�M:Ez�\�����{R��~�<��N�1���P�ꛅs� �k���w�<Fm<E�����B^���ᰑg[r�<9�A%U.�0ʂ�Y��á��o�<iVj��G�,5	�HƜXȰ���f�C�<�,΁V͐0H&"���M�E�{�<��֦&�t�##�KwL����B�<!"#��,�*,���%�<���Y{�<Q&.q3dhCB�G_�����\v�<ѡ �!uq��`O:�̑0��q�<�th�)M6�2�
7�V`2�AC�<���Y(�"���h�!d�hr�LT�<�C,��-�B5
�쎜JF�FCP�<�dO��Ix�	�xM�Uz�+�v�<����$��x��,��N�:��p�<�$������k�~l2��Qm�<Q�@�VuZ ��Q�Ұ����e�<q�M$@� s��L##H�!'��d�<a�ǥV�~��䂐�KVة���b�<Y��:&`��F_#�,�J�h@z�<��������U�F��j� �u�<I��5p��-ڬn��iz���w�<	��O�,��Ղ�+�88Q�^�<9P#�	�p8U�R�G��yZ��R�<!��	l�2|�$͕�Kx(RcJi�<�����6�vM�q�	��\QF�\�<.�6qqxȁ�m�9�)�E��_�<�V,�tP=�7
;}T�P� e�<I�'Z=׈@j;	vH�!��j�<� Bh���X ;��@�O�%<�Y�"O���i,b��u*r�:M���'"OqA�
Yi�$P��@ƃU
�0F"Ozeul�Jt�X0�D�ފIY$"O0+�A�k!��ʝ�t6~�A�"O^0���
i� �@	�x��-��"O�[qJ5O	���:0�f̚ "O��k%�@��XېA��>c����"O2\���N�A��4��U�xHH��w"OHrBX h٘��$J-N]P`"O�dq�"�<*^,�r��V����"O�\b���	V/�lK�h[�@�&��"OF|!Ƈ	%%�9S'���
�kb"O�<�&C�=<��)�'D[�0�K�y�#�4ń��e"@��n���y�W:4~��8#�����rĜ-�y*��[_H�;pA
�|h��÷�yrA��w��%q���*w�:���d ��y"
�=���b
�%=(�x�MJ��y2�T��pܛm+,�PS
�$�yr	Ĩ*=`)��e��V�P�b���yBOL/<l�������â����y�M�5��0��.���qҡΗ�yrmE���$q3�̯
�,� �i���y��4�l���DZ����!�1�yb3%m�xb�%(T�¹�wiH?�y��]h�e�`���p�����yƦ4���u"֬U��A�!���y�*L�|�X���K��A�5�J��y䖗k'�AR��!R�d%a��y↟�S��a��[,L%�� ����y�	G8g�D�K-�,A'�qAC����y�/�5����MB5��0C�\��yBa�1L�Ρ���6u���Ó�G��yª
�4F%����tŖ=�� �y��ΰc ���3kҫfQ�@��	� �y��J&t�bB��;_��h�h��yBN�x�lhC�&��ش�����y�F/k9��(�I��Uy�(�GI3�y��{�N�)@M�Q5~�y���8�y��_�[�T���*��) �'ߌ�y�cWU�!3���gl�����yb� 8	�&p�v&P�����
�y"��n"ѻ­� ������B�y�.Ye�T�����IR2J��y�!����ᐉ5�̲q�V?�y"h/Eh�L��!��,�xp6��?�yr,�4`�������)n0!�@%K��yA�m�|`͚��.��᪐��yb�ɰeL��L�8;����聁�y��P�c��8I��֟B��]�g�Ǐ�yr@T>ux���+�1Qw�=X�
ٽ�y"Q~�MJr
� �Dq�H��y"�n�k����#�F�R@/��y���@�0ҧ�c2�"�ϒ��y��]���d9gkZ
DĤ�F2�y�.�����5�'/n,�%���y�o['p��)*s��t����4�O)�ybA�	�Z��`�\li݅�y�@G�b�BxgGˏ)����ؠ�yJE--�D�`d�[~ɋ#��'�yʶ~����	�3�슳�¾�y�-�%EC�,YY��ДQ�����>^ɺ���/n̴�(P�L�	c�H��S�? ���"�M*�+��	$KҌ��q"Ot�w+�i��� ��'@-�L�7"OĴз�N(~/0"$ڎD��"Ol���8�*�h�!_VXt�3"O�LzA%ŏN��La���p+ 8�"Or�����X�a�224P)"OlI����K�M���"��i)�"OҜ[ 	�b
"슧�Io`��"O|�ѱ��X�����38���if"OP�g   �