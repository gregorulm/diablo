MPQ    ��2    h�  h                                                                                 ��Y=Ô�%%~�[&���S��%6��8q9"��ʜ�a�����9�{�n�݅ZRm�#7�Y�-��:Rq"?r��e/�g_A����p,5���Ôj�S�hY�2* ��]�!f� H��#ƚy+˝*��װ�v躹V�wt�C�N��gmK��o��j
��솙���;��:��Xc�󆇏�3�e0�l��En���.&o��3��ʈ���ߕ�y�4���C�h��X�o�]L�z1+?����M���"K]�Y	|��nd�����>�#��7	,��3I�i�Н_)�G�D fJ�2�����P�rjiS���7s"#: r��aĚҚB	��X'u���@��ڗ����ٗ�)�m|Q�3*�_�9��-ٹa���m�I
%D�t�R?�#AA��G��H+�O�ϕ�����[�O�V.?B��Wt~1��iFܐ��F'$���S��R�W�(@�&�Ԃr[DV��,����Ϫ̤��;�^Fv���"3*Z�X���u֛A��!|������k��N�N ��,�s~�X� Β���W_�N�%3�Do!��Lu���2���\��* ,��&�O�P91!��.�T@$��/s7rђiY'�C2�����6���	{���;��[��9Q��M����Q~l���q�~ji�擟��-�Ѩc[o\�Q'�i�	.GÜ�5�q��e+�B�<.��������!�V�	���2q���u�����vo��sU�����ʕ��ɨ��m�A.oz�L�,U�G[���h��B�t�u��qIB�v�p=�:
��W�������	m�D��q��8�M�`��\J��\�~���ߡ)=�����Y�R����E�b�I�J��_�TL>���$#𷄐��L���<y/H��5�@�Km!�����+Þ��%1�8=b)4�L��uˁ\��y�$z�zb8n��*�4HYL�3�p"7�4�U����$�Uu��8��]�텼�e�*�/�Zw.�� qE99zc�K����Y2=����y�{���Y1��Q��s�F{��y1胁χ�;�&��i�'���&�x�"�g���^"=��o�o�2�[n��Y��;��s���Պ�R����F:S* h1��)yL�KX��I{3ډ�	�����I_ �A�\;ԕ|Pmx�?ގG�?��7`����
��F� ���9�K 7����s� $��U��+�>[	��L��#������_�7�6�P�7"�`#��m�&(@��#�u(0��ێ[�G�l��&2�Ͱ��c!7#��U�D��|��,���K��*Kـ���U����/���Rƹ�uW���,T��g���M;M ���A�IM��d	g�����iz��ƾ��|ÖP���?]M�p�}�l]��??�Ԛ��O���z�⁫bT���T/3U`�=U�ɴ��\5�����C�:�%6��QY?)=��8�y�gu�}(+b��;1ө�5��nHL�D�J�႑Ѭh�����saF~И�:���ik��r��W_̡	��4%���生���R~u��\Zj��z���Up��s{��G7���y �S���Ӭi���aHm*���V�����A7�߸y��y
�yf����A�w�R��,M;��^�9B$9C~ɀ�-���K_������W���;������c�w�A�s9�L[���.�u��fQA�P��o��Q�n��Q�`֗Oi�[�,�X%g����U�5�V��Ǆ#�U�[�e̽���пe ��@;wdq��'��U3\w��k��'s����^~eGգO)8ʽ�$L8ف�'��{�E*~���}����/��.K��w�w�!�3Q���1��K!��m,Y2��)�W�.�|�׆�����+/g�P�¢��t�4�����,�D]f�a���wk[����6-�����o��m��@��s,|���By��9M��N�ɼY��^fr�_)��`:?$#�P�N�)��lL���qך��5���^O*3��[�s���ލO����kj��@�E+�X{�	T�?�4��f�a��iл�QW��J�0�y�L���}Ϛ�i��xDl������~��ޅf2�'�*�z�������eǖx�M�����^�0>�,"%ț.ұy��uq��h�WR�f1�S"{��Q����	(��P�;����4���!{���h]�7���ڣR�;��r=GR�[�F��xy��DT2��QIs0#Q�EI�Z2k*W�>_E��c�)��^ǈ��F5�aЉI���Op_�@_�6�9�5�Kז�:*Y6kf�$����3K��kV�����~���w7�K:/G)¶!g_�C�n�#�TWz�J��M}W�Ha9m	��?ZH�b�7������z'J�u��>���^z��q�C<�~yA�:�E���#L�;j�<�N7�̱��r��M����iw�/U���; ���8m�-���AƇ\*��~��|)��>�h��*(}'ٷ�����	��ePfپ��>z5��m^�1�Nw��i�O5R�����E|��������ME,���Y�_K�{����|��.�������U�6&h��d4��Ӈ�t���6����r[�fԞZW�p�	f'�Ĳ���E�s�vT��Z���{�R�H:�ճ�7B��p+~ƞ�:u>Yw��,���-�*�@���<�\���[��Wd�6�)��s�v���2h��a5���z��@c�0�D,+�����)�	����mY;�AR1bJ�0��/<M�.�kQ��#(RL�z�#���5Za�*Y>��{�IN*?
��9i�r�)�Q�	!�q����̀�Zo�Ӑ�f�4E���G�`:,�JvФ�%�G�C�{1B��4��]���8��[��9bn1N��S��n&�⡿���R���3g���I��%��2�Xk��G�J���Iey�H�Vz�΂N����e;/�S�SG%��y�I�Gğ�63_���`�	f�z+�NO��3������v+���#?5M�!��!�b�*0�*uc��}`{�,�mZU���&"���-���$+e]�ĵ��=wB�����}�c���/9�c84��g��4p�_f"��Ⱥ�s���چI���07U���͸?vo���=��V �����L?���e�x9}�t�G���@���Q����î��j4��@�75������XY�dZ����[���K-z)Q�d��G��@�
+֓m���(֣�$۸,�=�oP=jL�c�T~Ù�����ޕ�Ifˆg8Buh�q��(7�2�V�E��<�F��FF���v��}U�Jrr����ԝ]�x={�:v���w�(I��$��ړ�q"_�i���|�x^�ck��IHƔ��:����؁:�prKa��܁��ݳ$|U�;�[J�׆%��5���Sݺ�,p��w!� ]YV��k �I���AU��c�,:6��T���!��z���Yw���Y7��	3Qhd�nW��*�\�	-�4��WsB"9�e^z��)=+�lcr9'�x��x�_԰HC��0!t����;���)
S�gr��'����xaOx��1<�ĩ��@�m/�6���@d���+N�Z��6���儺t���;�熝��ݰ�d�O��.8�(����Y�EC�δ7��q%ѣ��o��X'J��	I�ۜQ,�����e�=�7I��҄�U<���۵b��u�!��\+����@6�����D��H~�|dz1��'�G�v�#���]7�t,��L�b߱��=��c�nWD�٪�m��G/��E����/�sS^M�m�`�+�\��a���������U��i��2�bR�����W�������z��L��U�������P�`���/�w��,��m�o������@�%�S88
�4\t�����w��yR�U?�n�2�*�1YG@M���~��痑��$yε���f���#� �)e��
-/Z2�閚�E��|c�>��Gs���0|���{C�YLb`Q|�s�`F����I1�Wj���>��UYi̽��@��x}��g�#���M�=�f~�x��2|�7nx#Ԅw;���s��e�%����SU����S���1)=�)�;K3f�5��$	e	�6���_�l�A���=�PH�?Tc�ڂW�7����B
ΤsF�a�����KNK;R�^���t���	+��-	�mt�f#���Y�ò��7�2t(��7�ľ>��(]�G	#u������n���'mCA5��+��>W�#����\��w�씇K�A��������Q�0}��7,��N־��~WWq�����^���7� �S}�|�M��1��&�g��������݊�c���q���N��]�d;p�
}lf�������I����ӻ�&���b�>��l�/���������B,\�����~�ǺbJ%�e ��tg?��ϒ�΂�*}�So��s���B�59K�HG�,DMG���9	����#8�ND�~�:��CifW��︿C�$Q�4�~��u9� 7M���}urp`�jel٦/�U몦s�������A ��K<����i�)a�����tVl�I�A2��ӳ�4�hy�!��ZM����wN��ն�6M6�E�(vB�H~�-;�K:�a�(A���Z�6Yq�2��cX�A�9k�t[�{~.��"��xy�b�"o^�Q�K���U`�'O�&ѭǦ%bٮ�`�a�NV��"��b#��>[��J�["$кv}�1q#;2�vR��37]0���)���H����G�jF)Sh���{8��'r���]���s��������.f�=��R���\*3�S���p4�F���8���/�U�ҜC��0�I"���b��h�g-P�)�������){�gj�]c����w�b��|ā3w��Zf��J��J�mE�g��F/|GE�����T���&�㤤n�(Br\�����?����e�Dלl������է"5*N�meO����5�����d۫����:AE�'�Xv)�T^{x���l�����Z#b�g: �F��J5��y�K"�k��UCݱ�Y�D盿��;��K��[�8�a��'L4Cz��~���NeB��(Z����O�0��,}Y���y�z�q*+��2<�fl� "\1Q��A�d����S�V.G�g9��QK�6?]�b`�e�Rb���`�=�[��l���7������{�w�s�t�Q�zI�kB!>����!�)�j���jG!oa����>�?p:)_O�1��c�58`����*��f�rJ��3&��k���xc��y���m�K�0�)8��!�4C��E�h��糧�l�j�LWc�9�-1�v�+Hm��7�/��דuI��N��1d>�����l����Cw����J�5js�	��#^���,��t ù���t���ą`w���/͂�-�\���� ��s��mn(����"��7�ڏ7��L��q��C�e�}�>'���HB_� �,���Hѹ���[��S�h��G{��M�O��|?�M�ٔ|�8G��{%��E�TB<_�8>�YV��D�㉻��O�Zf�Us�hŔ�d�P��Bk��6O���yˠa+���lZ���]�'/�D߸(���TNfE�5S鿶��(Ś���-7��_�+&2ƹnu����q<�X�-,@�`�<ޖX�l{P���遱�V��c�v�߁2�a0K:��\�:Q�K$�,��������d�Y��@mT����%b?���B�Mi�Ck,�A�^��t�u�5�W��\2a�Y�v5{��]NU6�
$09d�ׄhُ��@q���D��%�o�=���E��^碻�:�8�v�x�%!�IC�.{ld'ݵ���X]�+�[ئ�9}-�1�6bS��"&�9O�<�-�$ů;d�gVE�Iݛ\�m �XFQ`G؂O�z��t5��QѫGNI4��s���zS�h��$��D�H���W3�1���	�Yp+�A��(�r�e���?܇���?�@�!�
��i�0��a��}������m���/&=K�ը��\��+��h�_���8�#�i��d�2�~N� x;�#$֞�}���)�/�F_����]O�����U6!$$?�k�U���ͳ4�o�v�¼\X�q[�x��'����e@�Tx4=�t����C�K�()����E�B�jϨ���37��6�;3N�sF�d�,�����Axk-,d�_$G�����֮E<�P���9t���5=)�iP8�zL_û�
����X߳$\9���9BAnq�kg���Y��`C<]�a�!珧�q�6}�0=��r�6��m�]05�{Ն��)��N(DX�$惟�q	uq=�i��֋W�$^06�YTIC��E'韧iH�UJ�흍��~8]-�N�bU�,��sr�J�ɴ�@(E59�S�@�gX{�` X<7�t�k�A�I�(JAО�c�$w6ƿ0��?!�Y �,;�wi��YR���f�h?Z'W�����v-���ϲ�"�^�V��+�Tc�B��DB�s�_��PCMR!� ��;պ�d����"ה�g�O3� 1W֮�$�^@�+/�Ur���F_�X��D����6�����;����ᰗ���������Cb��g� =r�	ꎢcNcў#�oC�'��	d���� }=Z���ea^��2�H�?�?�W�s��&�ې�=Q^.u-�s��bÄQ�&�H��� �gɿ���rC`���=z�4�"�WGg��ޢ��x��t|��'u��"g=",յ
�W��Ϫq���å�g3���)뮿�MFat`���\ �ҽF��#������e?�m(R=Y����k���'0��ˮL4G]��P���t�뿤��w/��ӂ���8"�mr6��`��Δ%g<�83҄4�;�d��ӣy��X�0<�n+˂*�S�YB�"�&���%���\$�f �h����Re�B�eJ�Z�C����E/�kc��q��!����w�pv�~{�AAYg-�Q�3�s�^sF�:�7�21�Ko�=s⇜4ki�sK����xXTeg.��Ŕ�=�%��Ӌg27.n:�OI�;�"s�Q���<$��݀�<��S���1D�v)oK�KeM��ڿ*�	����\�m_��\A+tԋ��P#��?T9��u��W@�J��
��9F��f�vE$�6Kv�D���]���@w+JJD	)?W�}y#��"���T�P7��-*���7��YD�c��(�g�-u^�X��p���60��\X�ͦl6���#��}�:���rE�������'�vc��~��rH��y���W�g�����W��CT= �����MO����gP�C�D���n��V��L�M��D]��=pַ�l�՜۵��
9���Ӗ��X�b�����8/�#�������6\+��س+W���!%H����1?�a⒮�Ν�o}�H�������5��HB�D���w���󉞧��)G�~F5�:3�ia0S(�B��Fڡ?̜4]��#n�;��HS�uzv�6j �ۦJ�RUfԇs�����-�A �K�k��A�i{}a>6g�ĩ�V<��u�A-;z�nLK��3�y�]O��
w�z?�Qw�M1��ͲB�x�~��-���K:��c���Nu�1)��rpc�cAg9�ׄ[g��.:��꜀h�]���oZ2QI��r�`��ZO�њ�b�~%]?�ǻ��!V��O~,#h�E[�=���mе��̌��;���.%��$�3cf@��]������UGKQ�)n&����8���'=>s�{�d��:5�j8V�N�.�F3�m��¸.3�*@�g/��A%z����Y�J1�M������M+G�&�#���gs)����1�*S8��9��WZ]��.��DHw!���7��N���D�%:P�ؑm��F��9�|���블$�o�@����ӶcEr�ޡ���?�������_}lB�謷���)5�#��hO�c����"&W�E� ����JS$Eah(Xq}
T�NQê.`�������BC�����J�gdy�j�Ij-���Z0Db����������\�~'�]�zsV���e�U����31�A�0��,ح���qQy�Q	q��m�F�f�"�H;Q�g��@�b8{�q�[�������O�.��]����uiR`��X==�>[~梓�:�z�����L�s���QV�I}q�k�L�>�����O/)�K��>kQ�,�apX��y;pԡ_�_��o�v5��L'*�C�f����?3(�ḱ�g��tR��-�5K�R�)ST�!]8�C����_ҊU��ܟ�/�W��9�q���iHH��7�Q���p!į+���i�>ƽ��T��QC� �����0B=�d��#� W����Dқ�Ə�H�]��/	ٿ(wT�"/�кH���1?5 �H��aBm	C���Z�e4�J��<O����G!���}]Ď��X<�������v�����4��iBƎ�d��8��Q�O�8���1��Z�|y����4�K�EbKA�O�_���в������g��T��E-U�Oh�.d�)6��o�Qx�,ߵ�{p�܈.Z�������'����s����r7T����L���a����97���@
�ԀIu4�^�\ּ˓��-�K@�[�<9��'!����6�,�O�vs�v2�2�tQa+e�0␷���flQ,!T�ci˗���+[mO=����b�����u�M�;�kd���>����pwr����Y��a#�Y4X�{y
#N�bY
��|9_����n!���q+�7�����oU"�͜-Eۅ
����:��Gvm1%�DC��P{����P'��S&���[���9�21D��S���&����׈=��ӯ���g�jI�e;��-}X!G�@���oeݿ���PN+�\�[��u�S���!���?�%�U��3�z��'	\�Q+�T�c�J�  ���(��U�7?�Tp!͕��XX\0����`�}�'��
t)�#���}��&X�+�#���7E1+�E������3UA��c �陯��{���7���6��15��*�_+M���D��������K�Ul�ͮI�oB+1�w�+��N���(E��s�,e��;x/�t;��p���&0�������W��jj`�~vv7�������юSRdP�q�y���|3�-�NO�Z~sGi�\�y����=݅��i�դ3�.��=�j�P3�qL�u���5֙��&��K4��q7�ݺ�B�9Iq�wU��ǨP��{�<�Ig���G�Z�!Ig�}�H���r����'�]��{��~�d����(?��$AeD�,�qX�i̍�2��^k(��XQI>�a�3�b��pٵhF��@�@Z���M�U�dE�ΩkJ�쵆[�j5���S�t���`u� � S?���LSk��I��iAK��cm<6�`�DVr!�'����pw$3�YmC����!hPW.�8����-�F���+"�Ny^�G��F�+~�Zc�k�Ů��n3|�f��CZ!�F��uO;�ӷ�R�ʝ�h�g�vu�O�}:1r�ğ�U@��/$��C�Z�{�T~r��Q�6�x�z�sqtp;6\����^��n�d�����^I���Ά�V��D?���J9љ�Gom��'�y�	]�G�X@"V%e��Y�-���p����rp��z�a�k"���uȦ����7����B��./�:KO�M^���0�zgr0��#Glw&���/�=�t����;T�'��=��^�	�sW�2f�,���#,�����nd���K�M�t~`�"\[{\ˍ�Щ��x����è�Ζ��sR��⁩�"s��{�A���L��ȵ�5T��`��3�/Y]0�f�Sa*m��[�y�W�O{�%��8.�4#�����yJ�Ynf��*Q-Y=�����ίe��՛r$o��p0��KG��V�Se��	���Z�����)E��Fc������*��r��R�{��MY��Qr��sv|uF,�Ҽ31�_�Ϙ&�W3!iJ��6��x3�gi̱�/u=�P�.J�2��nU���-3;��"s3A��[轇䗢S[�	1_u�)�z|K郅�	�Zlc	} �����_Q�1A7���JP�u�?�>ם�Hɗ���<g
D�#F�E���
D�OK�l���f���f�$+ �	D�j�X#d����9��p�( mް�7S&�t���3�(��K�5�u�����I�$����Xw�l�!���"#7�o����m�W�=E�R��0U���T��枇έ�P��=X���DW~m]�W�pĄ��' ����IM�3���
g�޺�Ou�s�Y���'U���S�]x�pф�lB$�p���%M��f(�q⮦�9`b%�^��|/D�N�n}`���\���؎�(�0-%�$Y���?:$5�i��θd|}��bC8�Z	{5o�UH=��D��2KB�"]�[��j�~���:�Fi\)�� M��j'�Zg�4�[0�y�2�v)v���uڟ��j۩��e�U��s��«��MȾy �����Q�� ri'�?a��w����Vw��AA(�f�����Yy����>�lNw�$���h�M,�9�o��BUȶ~��-1�JK�,�����(�(�,��amcΧ�A4M]9aMA[B��.uVN�7H�W��SoԿ�Qf�2�`g��O�����U%X�M��קXV��d���#Cf�[L����=�а�k��1�;�wIF{C3�,{��������	��o��GX )�����8j�e'x*��%,��!�����`�.�q��x��43"����<׸�����(�e�����iވ-`��]ɻB�g�E�@Yw�,ܔ��6u���d]7���ǌiw|���	�ik��P�n� ����m{�݀�Li|�	��sR�ɊLD��7�ZԈ��hxr��|����?5�2��[��zwEl�o�臊��K�5`˭�hO;,������=q����r�k�Pㅌ�E�ȆXl�4TB��e�����r�P�	�l���Jk3{y�����%�����{�D�����e��@���W��'�Gz.���:e8�v��7ݻS����	0],3"~�_q'y�H�q ��o�f�u�"LU�Q�m�����Ɖ��-����?���]�����+R�|����=�C�[Yf)�)�����'dZB�sa��Q)
I�,�k�w�>xI�4�o)�LHǙ��wX�a!��4�Cp�_���
�5��ק\*���f�nD@U�3ܨ+k�ͮ���o�܈:sKk��)n�;!���C�dF���%�F� � ыW�N@9����l�H#�}7St�S�kN���ǞD�L>���ϱBg�"C�ݯ�OG%�+:����#}���O�y���kz���ٺ�w��/C>'c����t ^ ��4Um�}��֋o�m���	�L��g�l��ɔ�bh}�i�ﱐ�����{E��~ѯ5��c���Ɍ�I}��uOF�����Ak|�k������3E��6�J J_\���iO���3������P��D�U���h���dE#�Ӹ��l���^�V�����Z(n��F'��h�.h����TD[<��澿,̀^$��C�7Sh���{���u�yT�7[m��S-bA0@�v<�k������nL����Q�"vmL29�a&�k���t���?��Գ,�m�>Dh���U���mJ�Rc�b{�P��bM_�k��H���#&*k�C냹�
�a>�9Y�Y�{T;�Nˮt
R�9Z�:�)�:��qF	��:���7o�y�7W-E֗�X>�:]�v!�%��C��{���Ђ�N���I�[N��9�
1�ۅS_��&1���r���T~���g�J_IP��c[�X��GNSf��h�j�A�g��GǝNF�M��D�P�S�NK���.�:�İ��3�#�0A=	��+r����~���u~��12��?f�!�@��f0gd��<}1�e�H]�~��8�S&sW�՞N,��?+�s���j�.������I��0����\�kj�挒�� �%N_w���$��s;�K�~��T���U�m�ͩ~do��m�2����Y�ncs��|i<r�eve�x*�t���+�y�Ar7�`ۯCܮ��9j8i�yAu7F����ѩ��d˞��T��Ϸ�-K��U�G�J��4�9��Uf�F��/c�i=_�P.-eL����%�֝g�N���ڧņ�OBFR<qգ�ʩ�cg���C<S���׈��������}	���m�r>5ͮ) k]&�{�~;����P�(:�z$�fɓ�B�qsK�i���0M^�:����I9���_M��3���$㢊�b"�{w݄�Uż4�)FJP/ۆv<85�$SnI�݈��HP� Nb-�*��kQ��IQA�ϭcHt�6<����|!� ��u�wߋUY����z-lh���Wi�-�8-����h��"j2�^ˢ���+YP*c#���I��i�����BC�Ȁ!Ō#�;�9ڦ/�8��Uu�ѣ�O�w1���3�@���/_�r��+[U��������D6(����8�L�;q���R@S��S��`�=���yP��]��֐R��y��g�єcyoȁ/'{Z	�O��K�3�U]��e�M|�(Z@�J�ҵ�C�M�����F�J�T�uc����·��x��v�6��ɵ��(�t�-��z�l���Gǧ��T�?��tr��� %�bE�=X� ��NWU����a���f��	$�I�.�$�GM|��`���\���HA����/�Ã�-��v�Rsv ��M�έ�6�7�˓�L*�Ȑ�ʷp�!����pe/�9��!y	�n�/m��Td1ÊH�%�8)�P4m*`�ڀJ��G$y}���Tn�[�*��>Y8Y��+ׯ ����P$��?�K6��*���&-e�^�Zc�#����E%cg�X��ݥ��H�mj,�={tI�Y�#1Q���sQ�Fg�m�L1ԓ���	�R{i@_��Lx�g��"�ʐ=�߉(�2�Bgnp�FE2;�&�snP���	V�Q���mS31zA�)e��K�­5$;��͖	x�U��_L
ARy�ԁ�QP�_~?�c/�������� �)
�$2F��m�l����K�7ǭ/�'����4+��=	_9��#?G��
8s��\��#��9f�7�1�ܬY�3(����{�u���������X�)��Zٟ͜�ϸ$#r,��pf5�h=����r�<�K�_�lf��������E�!���MWh�����ө�9�] ���-�NM�����,�gsX���;�.���ԅf������]�1�p�q�lwΫ�+�
�@��XF�L$��ζ�b��R��4�/�r��) �� �D\!���i�*�k�l%~�����?�Ȓ$���IQ}�_�=��ӕ�p5
��H8E�D^N����=-��.?�߬�~�QI:i�jiWB��8׿C���u"�4za�T߇���h�~�u��,*�j�xͦ��sU\��s�)�3H�c�� �O�Mh���z�iB}Ja4ԃz�V�Iu�A#��$��eݨy�5>	�وG=w���Շz$M'%���u,B8�~5]�-�?K�M���`.��'t�')��Cq�c���AO��9��[�_.�62��/p�2[�s=Ko�E�Q7���`B��OU�*��>%Sk��q�N���V��a��#�[�~�,��Ыi��B;c�d+��3�΂�������E��ʫSG�~)��`b8E��'�6;���+��(ݟ ����M.����c��xЧ3=9ܕ�ݨ7�S�I�Ee�񀹙�CC{W���Om�\kɶ��g)�f� q�� x�P�����]Ҁ\���&w�8ʭ\;�����E��S��(�m�,���|X���.0�ɥ��pF�5��٫&r-J󡢘A?�X��<�ٕ��l8��b}�׆2�5�.��hdO�k�G���X��;pЫF#h���E�I�Xg�{ToU�� 3��;�� ������\�J�y�����φ ѱ�jDXi��}�{����,[W�R}']�z�$��5��e��N��֪��@ ��0R�,��e��y`�q����ù�f� "�Q����ue��m6���}�r��岇z���d�]����+�.R�R܎�]=3��[4 �d&;����}"�WisWyQD�-Is%k��?>K��
�)�m�����2��a<և���Wp˟C_ ������5�F�ȓ*E��f��[3�I^kB�a�I��j�����pK&�o)�f�!S�?Cqg��^���Q����{��W�;�9�Y)��)H�}T7�Fɕ��{f�.��{�8�>�{��J:B9C(�ť����&R���F#8�x��:��T@.�S˪��,ٵίw
Q3/���~�J�'�~ 9T$(�m?����9`�����!��|��$���lxa�}�/F��*�Y���Q��*�%�*��>�f����y"�ѹVO���p���*G|o5��{�����E�bd�E+_����#���������o|��d�UD��h���d�<��s�ܱ���"~r�1�;�R��ZÊ]����'@���7����T�
���A�gc��L���&7��v�\�&�
��u*o�� N�	\H-���@��S<�����Ɖ�*�"㥣,��v�a/2Թa!�N��L��kC���\�,���?u�+�a9�mE�2�Sb6�c�<�M��ak��$������f�1F�Z�ϐ�aYV�Y*{�{/��ND
ힾ9U�wו����gqaR�w�u�t�!o��=�ҵ�E��v糯�:��v<�a%�e}Cpó{�f݆���I��줠�[	��9�*j1:��S:Q�&l�^��%�ůLZ�g��wI.Z��ި�X��G�뿥KGekb�)/Na��Q��+3�S3�j�W�B�5xt���3K�3K!;	R��+Mڇ��,X�6�T��ZׇaL?!�!�N��0Bb�O�y}��9� <���g���kp&�u�����v�+Q��0$w�)�0�z;>��������qe_h���O�R�g��� ؕ_҇���e������������UU��ͤ�Vo����{������-˸&owW�e��x%=t����J�\�)����ۊ��Ͳ�j�/��t,07�f��l�����2dF�a�/����	�-��PʦG��������ׅ�V����ۤ��=��"P)�TLp��@m�������8����S�8B�Gq��x�e��R�� <������ǧ�ȝ��}�,Nd=r����D��]�*{f*ȳ���{(5��$��.����q�/ i{@���^�l�*,�I4��V��ؐ���W^U[�=$���F���U�4���x@J�$����5��QSI�����9 I�B��q�k�AI3� AARc#�6wY��z�_!�#:�=Cw�KY�C%����h��W�e��ō-�؀�Ô"%6�^�;y�+4��c^���d[	��+C~W�!�����{;fej��Ӡ�Ŀ�,�AOd��1�i�ĕ�(@k�4/�s��y�iP;֧
Q�F{�6C��p�"'�;�P������X����y�,���w���H����I�4��я3Go#Q�'6��	�aϜ=����v�e2�V�#�oYE��p���J|�p���!b� 0u�����4��b�1�y�T�Q�v�0�����h}Zz�M��
�G"�:�V�����t�E��&�ߝ0=󅺵��EW�	s��H���ɕx�޳$�9�_ĨM�:`�o\�W��1����c�^]�N�R5v���!)�����'�L�-��k�������@��͖/6�� ��?�m�9J�/��5�%8�88$� 4�Q5���ā��y�G1����n�S'*��Y3L�7~�۞I�&�$e�& Ə�-o팑�e��vb�Z���!�E�J�cBJt�3�7�`�h�g��]{/��Y�N�Qh�s,*F�&B~1��&�N���͐yi8V%�,&�x�Ag��G�e<�=�"��&�2h�n����V;]ړs�IՑ ��;,�MժSч�1�-�)�9�K�!�p^_ڐOB	sJq�mD$_�+�AmPF��f�P�i�?���Fu��w#�[
��dF�������^K'�V��8��[���?+{� 	z��`{#�V�E� �!
�3�;7� �����J�(��e3�u/�	�³~������~��Q��f�n�#������c�2��8�-`S�fI�痥��@��#]$ҹ���W�
�Ӽ������i� b���h8bM �2��n�ga���u���Iۮ�OMo�ݢ��:Xq]Tp�~�l�z3��݇�[F�wk��'�w�	T=b[�ޑ��/�I�����;�G\�[�D�\ǦC�%dr��@�?����/���N�}�5������O�5��}H3�D�<?����X�"o���~�D:2�iR{H9���N����4����/�l�����lu��?���jQg���t@U�4s[�?�nu�U� ����r�ti].�a�S}�Uu�V�(��iAA�S�xR� ��y�����"L�w:�I�"�M"��%ziB��m~P�-'w�K�8�Vs�^�W�"Y%����cD��AjB9W��[�N.�6J�m7��-t�Η�oJ�0QR ���`�6O���3��%N1]��}M��V6G #���[ν��Ц�J̝r�;ϴ^��3�4i��d�.3��͡��%�_G|Ŋ)� ]��A�8 ��'�b-�Llc��O�{����c�.����DJ�S�3xp�8+p�2�J��$� �񛭀龺�V�a���n���7ɱ�g���o4�ɔ�:�+���Sߑ]muWս|�w2�	�h����F��Ӷn6�jm�S4��ғ|�N��-������~�P���)r�B���i?�5*��L�ٰ��l��6�=� ����5�du�Q\O�`��8�sgH��^:�!���^FE2�Xb9�Tʈ��۪���FIb��%�2�J�*Qy��[Z%V�A*U�5tD����X�a�7?����Md�'���z��4�P1�e.d����h�ɡ����0g),�jM����y"�cq���#�fX�"���Q����D���8ʉ����׾�{����R���T�]�N.���qRN���5Ռ=��[�&���9�K�����Rs�7�Q_�9I��kq-*>��D�j��)����O,p��aW�+�*�wp��l_;s�@��5����]S�* ��f"�	6X,3�
Ak}����1��ew(�>�.K�w�)��!�m�CL���E��[ 2�4[��sKWOH�9����būHٔ7�8s���ca�<�X��E>���v���Cc�聾p`�!�C�u�#�(��}���v/����[P�T�Rٰїwe�/�y��\դ��U 0_;wm�R���-�#�G�{Z�T�]x��/�Q�}.����-��c���n�E��ѥR��S��?�ЂU�߱��O��+<��Em�|���V���~E3ʽ@>H_�ɲE����k���ɻJ@��F�U߷"h��Nd�u�.>����b�����]̞�-Z^ŉ�M'�z�ߤ'w����T:�cС�Կ�WY����C7	gi�Qk�%��u��D���^�D�q-��"@�V<J��X�ˉ�ρ�C�c�v��f2o�7a#�A2\�&���1,��&��Y�P�"��v m@�Id�b����:�OMU�.k�U��Jb�YW�aK;�ڛ��7�at�Y���{
��NA��
���9P��Az����q|��3�O��o�;�m46E�7�A�:�k�vW	%=�CK��{X-��!�X�D>��\�[��9�iR1� �SÓ&�.��&�����A2gBдII���Y�X�hGģM��ǋ`?����bN|݇�̕h�Sn�޵�/�0���fߛ3��f!!	ͧ+(M�����р#�ϣx�f�?�O*!����0����J}g�%��O�4���j1&��UՔa���?m+��O�ˏ��$����KP=���A��I�C3�֊��Yx��h_-q~�����b�A4���*�W�kU��p͟H�oS�¨��ݳx�d8t˓���\]e���x }�tLD��?�wVĹ��e3��ij;G��o7�7���'JL��:Od���
�v�-%3-�v!�K��GzUX��8��0�<�2�f��߫�=��PP$O@L�VA��8Q��D�|��s����B|�jq�[�Ӏ����+��;$<I�������jR4}����z�r��t�_]g�{A�$����:(0�h$R�s�]��q�3�i|<���5^����I/�7�����/��F��'��F��"ݺ��U�����[J������5�*S${�S9��~� D��3�kǸ�IN}xA���c�C�6�����!�QP��0�wU��Y���pt�h�%kW�㴵c�-�v���"�Y�^����s+�yc����F�_z�w.�C9@!�x��S;A�KP���n�)�SF��`�O� 1�ڳ�<@F�/�č�K��e�9�@L6^c�����A;��������}�Qa�|p���	�S�{�ds������ Lъ#�o~@_'�	Г0����69eͼ���[�_K�+_��g��h���1�=��u��k������3K�4���l��ɫ��nI��SLz8�ͩ[pG}h������ th���Lw���E=������XW��]O��/^T��,ų�v�뚰�M�o�`�np\lnu˾D�1����%�9�\�YE�R�D�����p�׬�Ϲ�DL e��F,Y��cW&e��JD/jRG�������m��
�� C�%�N�82�4#�*�P�b��;Eys'��o�nl�*"�Y._���𧯖\��&�e$��H���PT�'he������Z���!�E�`c �n>��{c���K�{�ЋYә�Q�-�s��F�_D�~�1�[�ϩ�����iS���Zx�7�g9!� �=�aM�?Es2#��n���;��;8�s����,W��E���S���1�9Z)[��Kz����w�+�e	n	�ȸ�_�+�A�GG�wAP���?@��'�R���
u�F3��b�[3�Kb��e������w��+6�G	�����#�&��Ⲽ�B`�0�7��r�dA�OC(b�nh�u�!5��5���X�$P͒�9�D�#�.�����^�ʔN��ၟZ�b���w��^�L�UH��[1W������	|��/� =���IM����9g���0Vu�d?��4�øy��u
�]��p«�l-G�ۡ5	�v����&�t�D�b�\��T/UA^��`�V%�\�,�����%�3���?K+����H�	tS}
����j�#X5@0�H.AqD���cՆ�s-뉊5����k~2�:��iM���	l���'����4�
�'�
����u���PpjvO��Z5UR��s6�����r ���ڋ-�ix�7a*Hr�0�4V((�PP�AcT��qj���y���WT��z�wu�ս�pM��B�wO~k�5-��K��ՃOk����������$c���A��09�m[���.&W��_X�HI�)�o��Qm}H��3-`���O˾
��C�%I��'�:VV(��k�#Ԗ�[�ʑ�b�DС����BA;٪N����>�3~��,��ɛ%������G7,�)�^��Cv8��5')�Ӆ�?��|�u����U�.�*��Y�%�.ha3��ȕ�i[�-����uJ�>~����9R1E��9�c����ɬy�g�Z�qqO��{����Lw]��ո$vw�g��#b��ٵ�	�ӑ�q�mL���EC|!��K���k���@'����O�rc�h���m?F3�������Wl.Z��ñ��.�51�>��YPOLEբ��Rގ��1m����G�6�yEͪ2X]]T%��Öi��H���л��^�m�J<Vy�& �����s��P��DN�N�3��r��bh$�H��'C�z_���k�)e�SB�ot�\V��0��,D?5��0�y=�q�
�y��f�eP";TQ����+D_�N#���8@v]�V/���"j�,8]�x����R	i�P�=)U�[꥝�ڼ������3k�s�8�Qz�-Ii'kL��>����F)�Ǫ�z��
ar����S�p��%_vdȽ۞^5��l׸��*��uf=�(�	)3m��k�����{�`n�ܙ]�K�)��I!Ij�C'_��L���,����1u{W
u$9�,���H���7K�$W�\�����5u��>2���@	����C��-� 5b��}��H1#�k?���0��
:��4�	��-1٫�;w�5D/tG��'�!� �g�n�mu�����Շ~Z�6��/=|���������}�ސ�|v�<=�����`K�� P�����z��:��ǡAOW���*�`��|e(�1X��7g�E��g�;��_m�L� ���3�s�xIػ%$k�
Uz��h��dV�*���i���+������L��q�Z�ͤ��#'���_7Z��T��I�|4x���c/g���7d|�����@�Hu �>�ȩ��<�-3x0@��<������"�=��,���>vX�2
4ai���7`�ᄡ���K,p��ϔߗ�7����'m;�\c�nb�)�U��M��ks;���N��\'a�5}�E�a�r�Y ;{�N|S�
#��9K���K�k+Vq�D�m��*foA?��>EǍS�i�>:�H�vr}2%�4gC&q�{���ݼ�w�?N>�Z9�[m�9��10CVS�T�&��w�C�n�'�I�g��Id�G�ԣX�A�G�{����[�׿x�Ox�N���Gn���oS�����Y��+�3��<�3��)�A�	H�+���O�5�l6�����Qa?���!9��DRQ0��rŅ�}�)�������K�i��&��^��(�+ǖK�f8���0��9�t �gNI���ųZ��O��L�_�z
9%��x�����k~���&U�2�͚ݯo�<%�cۡ��jԭ��F�nڪ�@eGk�x��t���\!Y�����d �@���C�Oj�~E�jb�7W[�������3d<Ё�����h`�-m�F�JG�
�en��5^r��-��A����=0�vP(L&7!��$-�'g[����k	ц�?�B\�q��V.��ǔk���P<��6�h��Fa��5�}�E��ro��zK�]���{�Q�P�!R(+�i$�*����q�W�i�������^W1�`�I*t����N����U�T���,��U �U����:ǕJ��#��ʑ5,�S�g?���f��� ?���;�k���Iib�A7	�c��Y6�_j򰀭!��B��= wVbY��&��G�h�hTW�Ƶ�p -z�h�y��"���^t�o p+��c�Pk�O�Z�ґ�C�ԕ!�[X;w��ca�	���		���O�$K1�k)ċ�+@!%�/Ҫ����F����<��$�6y�a�fׂ�og;"ŏ�#�~��q5In�T��%|��8;g��0�p�j}�х3�o�O''��K	��9�3�K�U��eh�4�������ޤj�fI���!�x��u41��`�������<ч_�&9{�	\��I�zӨ�	�,G��O��m����0t��n�����=)�v����Wf` �v��J\�n�׳�g_�ռ�MM�`�u�\�TS�y���Lq����3�1,��\�RDj��c�߁G�gr��.L����!s�!������m/Ŏ��Rp���pm~^i����;p4%n#<8��4~ @�%��Qy�ɛwcnR��*�Q�Y)�T��p�Q:��A0�$[A��܏֏7������e��<,�UZ�k�<'E�1�c����h���)?^e�=4{�ĨY�KQ^��s�3F��>�(1��-��u�Cnbin�)�"9;x���gU��ś�=���ߚ��2��{n����;;�Es>4�ǭ5�o����SG�[1�eW)�x~KU?��2��Ʋ	i�#MI_=K�A�^���;�Pj��?{���|�L���z1
0�5FN����`|6(�K��� H���P�ғ[+��	���V�#��	����W��iJF&7?i)�<Ь��(=>@�-ue�X�դ��8��S���V���`:�##��A���Y�~���I��l�M���ZX�Rb�Ι�^���,���Wy�I`��$����� ;��ަMV.D��RgW��B����E<�Óp�����]�Tp���l�3C�\�����m���ݩ���jb�ῑ��/�XN�Z�S�qF\�v���kQ��c%O#l���*?�m�U+�$��}��|��b��FJ5ۊH)�Do�A��e��]��i��p5z~m�::�JiHM��v�t9����4��=��h�b���Ouu�)P=�jǤ���`RU̓�s�}��$m4m� ��^ӈ��G�i��a�\����VcG��V�A=��5�b��K�y#j1z�3��ɡw���XoKM������BAG5~�R�-�dK\ۃ���9�]����T_�c�R�A�U�9Mc�[�x�.a�꣦��ڷ���o���Q���yt�`�&�O
y�i�#%D�ǂq�êVC&�u��#���[8!ɽ��fМ|�S3a;��l�$��*3Y`�gt��d$m�ù��۝WG�)�����dB8��'d.��3{�w��1X�Lg�.t9���L�	dv3�>}�nȞ�(�L�Z��v�������	���tvM�-h�ɧvEg:�},8wj�ה���4����p]��ճ�w�.��:��s�<W��l�����m�rk��خ|i��_����`#�t���Ƴ~��5*r�	h��RN?�P��m�&��7xl�=T����7�5�/ ���@O��ʢxK�ީ����2�׼�q�AEh��XX�T�O��QH��#��<k��OH��I'Jסy���B�Ϸݩ�k@_D�V�S����M���CX�'n�z�趆)�e$c^�Js��?6}�0��',�3�K��yXeHqj��TW�f�J�"��VQ���c7�	.^�����&�1�݇+s�5$_]�~�<C�Rĳ��kOC=�E�[ťd��3��f$�?��WEsMY�Q�.
I�Z�k'cO>����")��I�McG�a�ߋ� ��p\Ao_�u<�v�T5�*���*v�fX�o,�Q3H�k��.�Y��[����S�KW�)���!Ć�Cb2txґ~��&����W��89*���Xt�H�"z7?}���МWBq��80`O>M�2�h��	C������ZT�+��#iΓ'G��������o����}�٦7�wج//5�φB��ih ʿl���m����[��'5��+�J͋�S��e���}d@��U��j4��ʨ�{�Kћ���ώVƵq���ˢ��E�O����9C�{$|�Q|����rۘEi�=�6�6_�.���k�NKĝ�2� (��Ue�h�?d�HӤg��]��\8����EZ�����u'Q���gA�0��T0Ż�W�+�b��PX��Ü7�宊��`�[�lu�哣�˺�`-��@{"�< �j��=��=�s��d"����vY�2��	a� ��\ķ�U���N,�[����<����2RGm6�k��cbg���pU]MK�kNA���Z�-W#�W��� �a�0�Y���{�>NN��
�9F9Fz�צnˏ&�sq��`�S�m�o|�ͣ��E������:IE�v��%L~Cx�{��:�W��:���5[:��9H�1��^S��&�"��/w�4B�]pg�՚I8o�OQ+Xh��G:t��=V�,��C3~{N�g���f��*S�µ(ď�&R]���3|����	��+ޒ���R���ŕ���+?R��!T-���,0�� ��}�*F���E��z�$ȟ&��Պ�r�~1[+������Z��֧ư�� u��r0�z�� 㜒8f0�6"_���y��0d*�7�KF}���.�U&�%͕�o	�b����B��Z���I��(�7e�W�x]�t#�������
jc�WJ�~Cjjq֩�e��7�����u�d� ���Z?ϣ�-�ې�A��G0�5� ���P���2������UX=��P�L�7��q0��B꼑:���F����lB���q����Y�O˩��<?�CL0���P9�}��E_wr*�,����]@{��N��g���(&�$����5Yqߛ	irqw�yK�^�Ý�XMI%���gQ�	�;���0�,����g,��dDU�\����J<zن���5���S�t���ie�N� :.���Hk=40I�g�A��c��w6(?�K�!��Nk�w�.�Y����f;�ha˭WU@L���]-u#W��=�"V2^7Oi�>x+��	c}ŵ��U��-�C�Ï!1���;�/�7�ʤS���=��O��91���ş@���/K�e�J��A���}�w)�6�{`���T�~};]�g��Fװy'���91)|=��v�I��B���k�@�QрcYo4'g�9	X뜮a+���IKe�7��gj��ҡ������I3۲1&��&uϣx��&b�s���FѢV�ɡ����޾`�zn��]�G3��@)���ht^�]�I�	�N
.=��x��Q�W�;��Ӽs�ez�����xz��M��`ٜ&\"[��4��gzġ!����˖ϓR�0聐U�:���"t��7��L4j��٧�\"���Ԥ/ ��X��|�m� K���8�v��%	"8":4هu�Ƌ�4�yi�R�rn���*X��Y$��H5y�8ڑ\�$̠֙��V�r��]�e����,ZO���W�*E�cc�"h��֦�1_�YN<�<�{`�IY	�Q��s���FS2ٟ�1����_�ه�Mi�Xh��rHxz�Mg�!��6�}=�?x����2�)n�g1�<;�VsZ�g�b$�褹�^�SF�1汼)QH�K0��!̈́�a�	d)��~�_���A����mV�PEG?�8Y��	����lYt
��Fi�]�X��=�K�8=���]����-�I+�lb	˭9���#��[��d���&��O�{�7�ID�4G�E�(�U���u t�2����D����e͈3�;P#^�؅܈h�T�N�{^�o���X���-#��ԑ$��ﭹ��PW����+�?�!�%�0 �;���M���ſ�*gr8��O?��g ��c�n�����3]%X'p�e�l�?��E������b7Ӹk����b,��T�/�^��jɌ�A\4V����W�s%�2}���]?Д���?v} ���z�Ӂ)�5vH$��DʄS��&����W�����K��~�
�:Ղ�iC�JZ�/�f��N�4�3����|������Vu����j��a�솗UHmms����Yw�(� �K6�����!�i�Fa �@��`�V��-�}�A7jߐ�:�Q��y>f��6��8]w�W��� �My��6G!B�6~�9�-�v�K7�A�����/Z�������?cu�"A�'9�x[�=..����>!��'��f�o{��Q�ס��Ա`���OAu;��3%?C���VI~;IV^�g�F#���[s�t��1�Зm|̮C;O�зpx�34&}��������uK�6�CG�Y�);����:8���'��<�G[�r�����H��5.#���O����[3)��	G:�#1X��xU1����I��/��_ޯ+��Q�ɢ�g��0���(+�Be����~]>�ծ�5wCjʙ�������Z�G=�Im�2�����|�%���h�v��8�{Ķ��(r�4?���
?����(���8�l$A��Έd�r��5gŹ���,O�?�3���Ȃ�'�����g㬊�E��XS�T���G��>�\���1�d��-�Jr7y���k @�rgz��ADD;6������r��Q�>�'���zշ���&e���%�B�z0���.0�e�,�G�P�ys��q�䠓/!7f	P�"St�Q~��/��X^��l�ۘ�K�f#���;>]�@����Ri����=V[��{�P�.����!�Ns�Q���I_��k.�>7���;;)�1��`La�"H���!p7�H_�D�0c5��n��*1l�fs��̦3#
k.�͵��V���Oj�K��)�
�!?�wC���m���,L(�����{W�.19E������Hj�7z�)�Zj�RկM���W�>hx�6��� ,Cp�V.��ƴ�W�#$QB! �&�^����4�%�١��wv�U/�BC�K%�ң �75�m��Q�1��4�ڬ�e}���2��@8h��}��V��N���L}�=�ٖa���\q���q�&|���	�O��\��閟v|[���)
�o4EL�1�_#���vJ��i�\�nRٻ�K��� qU��h�j�d���_,���c��<�˝i�>��Z/�̉�C'�gE�ն,�K==T���2�S�e�ᕭ�Q7��H��v�8u�7�~ӱ���&-i�s@v��<[�x���s�X�q�%䣘r�v��2@ĶaUt�R���WFי�9,gF��j
��<���^m1CwU�b"ٞ�H�M�b�k)g4����*�R?�L ���a�vYAr{�4N��
Y��9Aa>�5���.UqͶtc������o�-�>pXE�Ѡ��4:b�v�ţ%~�Cܞ�{	�i�� �5(��R[���9:�;1&(�S���&X���y�}|�����gsDI��>���XCgGu�/��ƪQ�=�.�v�;N�ܻ�=�6S�2��N�!0c�wW�37O���C	>r�+�e���%亢`��>E�w�v?k�!ox0�:�0���;�5}8�z��K�EuI��&M&�%�����YZ�+=�_���٠����������;�V�]�c�NT�;2��Ӝ�@	_>���R�Kp*���M!����yU�U4͐g�od��ٺu�.9$��g��$'c,Ce}d"x�Ct]º����Ȝ����R��+����jNƙ`u7С�X+�0BUd2�������6|-R���<�^G�մ�ۏ$�k�����H����ې�u=f\�P��L�Wa�,\q�]�&���2�!���?B�BM�eq�_ ���
����!<�R'����y�\�}�S��}
r�=/��]�ܶ{��ƭ�W�(!f�$cM����q���i�X��T"^�uu�RI �j��J��/ȁ�GJ_��k���,݋�SU�T��kJ�\���5u�S��)�2��O 5����:k���I���A-z�c�k�6c�g���[!�������w�'
Y����N�h<NwW�F�4��-p|A�/��"�^RJ�e��+���cJ#�P��P+uԈ�Cj�-!L�qu��;�,�?�����B��k$OP8�1��ā�_@�N/����l<cܧvv��2N6�7��\6����;��3�Y�$�t���'^�+*� T���-^����$��ַ�{��o��'"�K	!�D�)7�z?��7"e�������n��\Pxy�\j�ۍa����uj6È�������eF�ѽ�����o�ѾT��z	�$���G�ye��O�5P�t�_��$~�߉K =_h����:W7��#�怸�dс���E�K55M��U`���\}�O��$���E�|m4���;�
�Rzo���gq�(���b�R�:L��f��`7���(â�ρ5/{g_��_!��{Dmt���cñ*%�,�8�z44/ˣ��O�cy�=�-��n�t�*�0bYX���¯�U=�w�a$Qn��'��z���{e�T��cZ
���raE���c�UD�e	�̴�TW{�d�{oY$;�QT�[s��TF���t`41�w�Ϻއ���i����́xUr�g�����*(=��g�P`�2Ts^n� $�(�;��7s�|o�����#�乺`S�]1�)�7K݈\�y����	_^����n_��A��z�萭P �V?����g_�����X�
�z�F��}��K!�q�K	��6׷��Ƈ���w+g�U	�ڛL�Q#�f��1@��i^�
� Ѯ7�J�M����D(�3��&u�ʇ�w��F���J��|������#��C�w�1�O�:�_&����	��ӝ�������&sg���:W/� ��o�Z�ل��� �2N�T��M��ź��g�9޺a|z��+��;���I���&�\]��rp��l>lS������B�c�ӓMʦ��b�J�z�/f���-�ɧ��\�mذeǒ$�%�bF��M?\Rh�˦G�Z�3}{�����Ӽ\*5��H��D%2ų�P����/h�&��~�H�:p��i>���2���̡���4x���d��� �����u����lj=b��U�v�s��{�Z�5je ���%�^�i�2�a����D�V��!�aA
Q���5�yY�1p�6���w&�Վ�hM^���^B�F~�@�-a:K/� kP��v��Y��
��c0h�A��9C��[d"�.�w��ٕ�Y1�:A�o6��Q��z�oU�`�&hO| R���%:���8\�9��Vy��kn�#e�[�-��3��В~��	t!;
�4�j^�!f3�ݖ��D�Q���4�Gh )+ٮ�w_8�7'�S���zs�m+��D<���.>f���6����3d�b���-����*��t���-��������c[�ɝ�_g������������84�?T�]ه4թ��w�u�T��H��2R��"D�""em���^�|X���d��,���jjs�|cZ� �{r4n�?W���2�Xl�d"�f׭�5{k��4O]~5��R�������X[��P�烍E���XNI�T6����e��Y�Й2o$�?,�2�J��y}�V�޸�-���jD�?���Z�#�k3�l�9�D'$�Wz��,����e�ڃ ����J'M80��,U|���y��Mq>�
�fDu^"�@$Qyg��<H����.�P�=��ꇡS!�ks�]�:���7�R:?���I=��H[{㓋~������|��s���Q��zI�1k�5>r=���L)}�ǻ���2aÅ�GrpM�_'�ཬ��5������*��"f�cv"�'3�M�kig��P 8�Qܪ��K;_)D�!�DC��A�"O�ǚ*��b�B9LW;�9`�>�N��HE0�7�A���#�M����1��oi>����D�B^CO�`��B���մ��#��]Q�������m��|ٜ�w�|>/�pH1Ф�Z� ��KȬmF}�����"��g}��Mc�I��{|=8F}�놐�g9� �]��1�ٱ�ё��J�+�z��LƱ��tOhP��`�E�|��������#�E�L��,:_~+W�1��M=��̻����2��UK��h��dg��������;.�xXo�yp/Zʢ���'L�ߐ&�f�T&:D��¿��� *��â7u�t�|�Ƒ�u�6�Y��0} -ϩ@q��<��ƫD)��s�7��r�sb,vϹ�2�<a������W��#�,~�~�`H�<�-�h�nm,�~t��bݜ���[�MA��k��6�0�9�M{{�va��Y�P{v �N-�
�@�9<h��\����q��ޥ�����o�${��niE����z�:��MvÙ�%���C��{D��ݍj��0�'�k�[�d�9U�D1��S��&�#���Px�L�sg.[I�l��EYX�qG�č�R�L*����N�q]����rZ�SZ��^�P�.E���3�	�a�	��P+�X�� t�=�ׇҪA?�^�!��V��]0�7v1W}�����◠��ꚥ�&|jՀ��4�	+xcx�7~��N��A3<�o�V������B��v���n�H�jL_�Vcj��f���-2����CU\�͋\Xo����e�IP�Pb��W}��be�2x�Yt�����}�㞿� ���� "��C;j�嚙[��7h���a��K/�d�!��vzH��<-��`�78�G�ꓚ�P�ֆ���(`}����˄O=ʹP�L7����ٙxP��0�ܳ���z�sB��q�K�?nr�ŏ��84�<5�a��m���5����}�
�^r����˶�]��{�e��u ���(�$�J�I�pq�ih`c�/I^HA1laI�s�
}��X�-C�ű���2��X�&N�U�l��K�J�_��y�5�HS���?���\ 0Բ�L}k�/yI��(A�b}cjc�6����0w!�IB�&wA@�Y*���\��h�W����a�-k�'ϊN�"�(^me[��+{C�c�]��Hx�KoV��{C%p!g���Wn;��<@���j���ι��Y}O�b1/�:���k@���/��W��s�7=��я���6���ו=n�y;����	�oQ �������?����v���;���v#ro�=@'�T�	<�F��,�U���w-e9f�
�c 	Y�6O/-�ת��h��)8�u�创x�)�q� ����Fɗ{K�J�4���z��1���JG�i0�� x�P��tT6���#��Ĭf=��ŵ�i�WwR�I�������k��놡M~�`�J�\��m˪�������&å�{�Eb�R�쁆�k�uhט���m�\L��Ȳ���}Ì���~�/�����2��zm���vo��췅%?a�8�W4��@�<�D�j�hy_����"nL*���Y�C���J���䑒��$̪۠m'H��2퓆�e��*=��Z�e&��A�E|c����Z��g*\O��N�}{�_Y?�Q�'�ss�GFɄA�1�k�����t�i��]��E�x0�g���lv
=���߫��2�un�('�!;�=�s�KK՘q.蚭����Sx�1��)GG�K��Q�abڗ��	Z�A�4�_njuA�c��c��P�z�?,��M�L��%�"xZ
a�~F�TF�N����=KN�0������ؼ��+"x�	(�ǁ�#af��l;��(���Z�[F7pk�1��;4s(���Z��u6����@�������4��~ ����l#ԳB���J%C����1b��2�No����J�̊�Y���`W��	zEw�u�ل�� ��01M'��ŵ��g([��ə��ʥ���$��az][+6p���l���ۍ�7����ާx�nO�0F�bb/��u$1/�^�狐��M1\0؋)��l0% �ǝ�O�?��{�����uH�}�_Ǜ_
=���5�Z�H��D����O�[�߭d�v�4��F~��:��i9x> +���䶡%4�І�vX�j?� X�u嵻N�j���"3�U>��s�S��!� & �	�o^�5di�taZ?��H�Ve�*FA���F�����8yt���Z�iv�waL�)��M	cV��o�Brv�~�g�-�kwK��; ��e���	)��em�c�".A�+|9�<[?'6.��t=������;_o��Qٱ���f`d�<O����:��%5�Ǔ����V�~[�Y�#@BE[��'���Ѝ�4�d��;�Y�>TnX3�[X��5~��MI���G#�)F���8gʗ' v�S���h�w�B���}\�.Y�E����3�d��?�y�5��k���q��"R�%�����%���ɘ-'gK��]o��j��r�s�zA�]t(դfw�D���}&�2���m����]�m�#��QZ|z�����G @��bz�Wk@�;�"r��u��,?�h�30�y(�2��so���N����@��c�{��~-��I�)��mQivސ�#�f=\�$G�Ѣ���Y���}atlf�&��;]���{��R��k�*G�<�g���@e�fp��K�ox允��(��a�
-���8"p,Ś����	���S4>��50��O/RZn߱
C��z��Z=NR�E_�!�^5�g.�s�����1�:�,� �Ĉt�lw�7ZmgCDl�}��|Zu�y~�A�s<_O�tX�hjZw	�(�c�����/��AC}�������f����Q�(W0F�S�7��Y&�B����$(�ݕ���Y�FĠ Em���,���Ķ�6F�)(&�M�������T�O�c"N��<��]��5H�����v0P��G�O�h�B�|����3ԣ�ܕD��34~��1p�i�n! �`jPC��j	_��O���N�"nz�HM.��63�D�|!�(ȼ�@*N{����o����8��ݪ�6�}��AH�9g~䐧tJ1|f������'�˅㔬�]z�➨�@��狵�?"=W�GP�r�(˲ME]%{"�<b/��o.���7��l��{�Zp�O��������DB�e���7ƌ�<������n��-�_ �#*D�Q����[���<���5����~� VC�8�	8b��s���t6�j�0���9�M�5�i�i�ހu���-�̤pm�%=w/�����şq/{&����DC���q��'RU�3�R��2 X���T�����g��b�� ���R֓��kdvG����)�|R�/ɽ�&Lo�V�0��sy<��:�߬�!�Qg��>���-�Z�g}�yC���_sK�|��X��S�[�T:.��lC�a]��/�7�w`��-5P�S��_ػ�Q��&UdM�o-5�?n��;`�/ۅ}9��E/QD֍�	��#��-��#�я�2/P����TO������o��d��?�k�d-\5�6�	�\-��Y*�d�ۊl�Ԣ��]��H���Y�n�_����nVFϥu�x�s&�-���2u���V/мw�nA��Sr5�
��!�ȝyIi9
����@z5,�EC#�:�a�ov�ȃ�^���.ZY�Ź��"}�}?8���kZS��g�ufͯ�o��R�E#�"����4�b��=��|3[F��oRf�t����mhF �J�IG
h�|��!@p6����G��@N�7>seIR?���!�v&�k#p�$W�M�TQ7����ɦ�0%�_ѭ�\#�4!��!@u}
4�������>�#C0��U\-�B:�!W��`]�kTf������]��q���Y�׆��XD/���n���8��;0�r.^�Y,��܉E<)!�h��d�tq�r����/�T�	vAvU�	>ܓ�Fl<�3l���O���k������z[�7�>؏e#��P�
�os3����9�(����GM�݄�����e��֦$H����.�(��*�&����S�ţ��$e�r�*�(R79j]6ƅ�?�dg��Z\�#(W��p��G��N�L"G�mN�+?5	�D����DO��<Y�P�7YpLL����=~�R����Ɨ� ����^��n�&�jj���2��3���+*�Ch�q.׍gr �����M���2xUX�E`�8ω����'�l "�(%e�0�e4�}��Zwk�;E7�������˟p�����y��(�EEZ�n���?lу�e���AE��ZJ��W��1�מ8=N��<�B���S2 Y���F�9�%�Hc��o��5��\ƁOSf/�F��[\̧\ʴ�/���| ���?��h[l�	�T�[%a.����cl��75��v�w|h��6�{��AY�K�ª� }5��L�����f�?�ߏj���'F���f��s���șs	R�KF�Ǌ�pxC?�ކ�m�$�������D�29쩑�G]��f����qm�O�2ڡ�?|�>jGG�ZB�x���;�_�K��@T�V(uz�;G�7�L.���S���,\b!��IeT�������懎'��3��~�K7$�!2"�fyŻ���r���������������C
�P߯&��"k��������;i�M�'Wl��s��(��-�XD�2�����b�3VCU%�'��f��k����D��z�0�1
b��{�Ug�tjx�Zg�<�(ݶ�I��6��$i���-z�w��'�?!~�0�%�+ΒQ�Y��*	Zc�;�ע��D)�.@J�\lX�V�ۧe}+(���Z��?�)�3l�]x����-J��쾧��Ǭ���9�8�F��B�B^���?c�Y9(�F�UH%/��ON�ou-������S��Ҳ�][H�\6�]�H�X �N!?���hG��	��[Ո�?ԛ����l��5�v?�h͖�}�v���YP�`9T�Q��5�j�����r�U��8Z8���-69dû%B�=���̹7�~��c�ĝ��~�?0"�p^>yn��V.�P3Vm�B�܂v�m��0m��f���D4�j@��ɳ92h<3Q&���g3j$��w�uv"����h 4�2/W�!o5D�y���N�6.���Q�Y9��.R�x&^�ɘYV/�w���ΐ1������ �b�[��G���Y=%��)�+��֪�3�p�J��q-(���?Q���R61X&u���{�g��ԓҼ�߲��t���KIh�,r�19��g�B��o`K�<����A%,���'�� �9z��x'���Qd�l=��b��G�&c�e]�NENٯ�s� e�<fJ�T]��}��C	��:NQj�3~�`�gw0ڨ�X�I5�ɛ�f. ���'.�1�hu��Z��:��c����D:�ש�>�ZM���v/u��I:�!{G�z�F���O�!��y����Egpy��͋�a]{\�/�}!�kOj�T�����IT�^S)OG���F\�C�&��$ ������1���)�Tn�N���N�z]�Ht�+Zd���>Hv�mv�*ePC�鹵9n��\��UI7�a��W�6�iM5x�����Ojp�K`��݂TV��A�q��r���8�K�j�9H���G|^5����R��卵+�c�ͼ��	�)�Hx<$���R1���t�i��Vy�5
[6����ܑ[&���N�cGO���kƞl!�h �oj�0��s�Hwܭ�w@���I�Fbr�Lq�ʳ:`S�J����r����g��� @B�V��4t�/���N� ��Ig��
3B|�װ!`*����'	y�`Tp7^=�I>`�
������!��#�"�$w�b�tw�����K���0E�v���Z#�rި�#�u9�4��}���>�5�0cNU|"�b�=!!yf���kt���J�}6�ϑ,��1��צ6Xdq�|�����;P	��ҳB�+��ܩ�Q)A�Lh��Z���ro���ǖ�thva42U���>�Y��f���S:��ᴃ�AOu�Y��-٨>�u�#��P��no��Ø<�9������g�ݤ"5��KOe���D���٢�Hu�*�D����i���u�4�;e��*��7Y�6�??���\��Cn9Wœ_�2��`�LB��mn��?UgRD ���d�S�\6@2(�W��LlmG��w-�r���4 l�M��J���^�5i�FVj�y���T�SP�����cl��0S׭�, �5��Gm��Axu�mE�O��O�
�G BV%�{�����7�Z�Qc;e���%����f�����
�$����(�,Z�tؿ�o�l���{�a[��z$���*
���G���
8]8ف?j�B��shYY��~F�w%�J����o��e�ΪLơa�S6���f�[|*\�րO+��3� _	?8�h{��	ˎh[Eߥ��$Z���dl��w5�Mv���hx�1գ����Y���ʔ����5�b��<8���cG��	��R�
ɿ'fG�ԆZ�s�!�'=��#�����a��x�ͥ 鼅�<�d�X#�Qӆ��c'���vn{��Fn�3�b.������:���UO��8v""e[t��[X �28���d~q�YS��H�$��|�ϖ����ޛԨ�0���M"�bh���ڳ*nU�`�����bu`oO<5n��RwL|��*�
�^��<�,��y�������b�wq62|�aq�n�c�QQ�K�̶��޻)&0G��������D?�,�Q	A��6�=#e̻�o-�+��,g���eV��$����f��8z\�٣HX+8Ԍ�@�}���<h����F�ּ8�+�]��ʁ��)!�-��3�s� �~��A7���E��հ�M��`��ݒ�����h���hC�|��_69@_h�Z����1R�Rp�B%�ɣz�F%�)���j<%~�]��fF��� /ڹN�K�(1���|!
��ƓX�y�M�Fh&+E��XF�*ww����i�A��a����A^�M��p��m��:��x�ש�-�|�13f-�g ��Ej��*
���G!�P`|?g�CU%j�Z��!%�`&�n�7M��6g��P�z�{�җ�{��f���������o��6y6��b�Hb�'g^��yF�1�r�m;�!�՝���� ]��:M]��k2��=x"�F���~�D�0��Q]w�"f 8/�3�.�x:73�_�|�^�,?aÓ����w5���|!��DH��@&�ZK"���1�{P�m+�#�{���
/]�am�2�?/�������foN��ZP]c!\�,"V����Z�
�Ѝ����j*ip��b�2��5����vҁ���[�母������dv�������(SG(G�p"�]SQ$c���蝩���t�N�=�S~'$Up0 %�A����a6 0�=M
��Q\=(3�J��m7�T�4��y��(�//�cd�{E�($0�Ewь?Qi~�Ϩ�c9�! <�Ba�$� |��s���I���~y?�ߋ��� tI6BUp��#AB�t�ˆ7 �B�/~��Kch����ˑ�HAؙ�:y��˿�BP������K����9P�؏ε���gj��-�<_^2m l�ufj-��w6�Lvk�b� ��2��z��m�D�Q��'Y&�_�ǭ3��ª��`��!�aY?��Eӌ�]g1�sK ���2����G�G�Y&�G���5+�5����v3 �%4���(���HZJ���[��J@��{�%�3!N��Jo��~aD3ػ�N��C@_��eJ+
��1��B�T�v{�qX3"�җ����m�Q��F�WhS��v����)�>&Kz�\�����6��ۅ]�[�95��xBk(����G���P1�rwK�!��e��N �گ�>7���Jd��S,���7G���6NI43�ǵ`�4��F���I���%� IA��Ȑ��L~�unK��������v��:�a��kP4���u`׈:r �GU�F$�&O�v��԰��B�g��oT(4�</\�}��Oe�T�ס�T��2�s)������\H�/W���V�`�k�Q��)�� n�N1�2J!z�d�C*����_7V�Y��豋�g�w�VF���4�u��2,U�x����Ik��Nz�5!,��iv�x�j+��K{����%���B߯���������%8B�j����˟|�Q_oa�č���(���^��8)�	�v H� ��7Y�R��į�yi��VtD���]�c?��C3;�_i��cU�J�tI�vN5)�Ɗ57ܢyo"3�jϻ�K���ݡ]`��nd�Pq���o<����87�j7^B�'��|}��q0�1��Lm�����\��	P=�H�����X�R0���Sn�iϕ�Vvx5����t1��z<���(�c&i��Xb�k��Ql�����T���0ʣ"Ov��x{Fa�r�k�C���So�|1.E����x��Cb�
��i����b�C��r�E�=#
�P�X�����Ơ�h�Ҳ��7��rd�5�\,!��M)�+l��$�]q��հ���6��j�,+9Dѓ�þiT����6���頊�?5
>B:I��6J���� ��{��R�kNQ�w9�����"c�a$�Ӫ'*Xzg%o���.�1���I����>r���,�:f�/�2�,��r�9mϘ�~%�����1E:���h9�L،��G�ܔ��R�ux��E���#Cن�m�Μa�"�뮔rٷ9�d�&+$��}��b�O�auWb�$��3. �!ś;���<��D�1�^ �4���EH:5��e9�;<ݰ���č�@'L�4�7�V�tHH���m�\�ڕ9��V�����*�_���<D���A�q�Lp����a�1�����S��O�K2����o�A�d�xi]�þ��� �)�J�l1��\��mT�V�
���m�CXwY���?�������#r{V�-;�@�h"��ջ���\UQ�Q	�=_(��7��-����}�
���.��1�7eB>ҡ��
�bb�@�}wv�Bj�lO�N>�WCZ�ؐ�^
�hjoiޯ��q���!d��4�^Q�WH�&\V���}K蘏�1���#ddQ	�����N�"솾��:�ʕ10�zv9��ĈK��u26QW��I�4篣�*������y��<���/]aH?�(��m9&�|o=�$Ԫ��	TuqrFvSeG�D|_��aG������3���؄@�E(r }\�z䄨�9#��>�C���¿q�IĬ<x��EP)�z��,�ZD[����q�!^|=a�c&�D��+:E����k*kC���;�s/��t �"&(��0 �8�L%W��D� ,�!�s�&���Ui�<0Z�;M繭��Sm�>AC�ƣ���qJW���fO�1�DM��Ϩw�2�'6藨�K�ګ>r?*q��ͼƋ�*4^�oU�m'pX,s�^y4���)�L�����y(4�0c����ƐQ��Xݎ?�^��6��>F1�2y�R�s�ۘ�ܖ�8��us ��jο$���t������a` �-��r��
9���0�%�J������z�8�ٰ(�Be�#�bI�/4�z)���"���M#�W)c,��B�M��cTTc ��3����-o��H]��1��/d�7K� ��/i��*)�Μg\�A^F�.�8�.F�*��Wlk�iP�� ��;��\�?�iCr�wD�~�^�l�@���{y'�P?���V�C�������C�nT����^��P-@ouڢO�$
A��Ī��+��R�M&���L��������;�x���RJc��ļhM)[����Ѹ%pl���qt�O �I�0!�z���6���OZ�2$���� u���^���4m���$�D��a�<"��R��倬��^���C�puIV��L���Y�߽��L�0mDG�n�����*��W\�Z�����fJ�����y��b���QAJ.�cWSV�V$�_��L��똶}44'��s��-�Q?�#�Qm~��8#��S�u+�
,K$p��$����|���P8޼?ه�?+��a�$�}�<L�� �F�^c84��]�I��1)�ݒ�Ilsz������%c��:�I����߱�`�B+�����e�C�L���U$��߾3���1�B�p�mĹkP(zź:썊��N9g~|�]r�F�ac��׹�5�Ib��q
����| �1q8F}r+);�X���w[p����A�?)�=�|�N
�S�T��m$���О�CZ�ź�'2o�'�h���j�1m�+�2�T?2Ś>�?iG#bg�n\�`�_�Q�K�m���T�nu�uGUL$�	�آ�J!9�w�?�qTU����R�Ap��M�40���\!h�fo�b�^�r
���s���M���u������G�	ߥ��<�� -��NHC�1��M�� ��թ'%�y��)M-'��h����b\�kC˶��LȚ�M���1��49M���0}�#b<����.-t�.��4��ߥ�,;j��ݴqxͺL@��Y�v)mJ*���ќa'`/No��-�͈�xwń������A��[�T�(!Lcl�dNY|4�2����(U{�G`��p�,��c�Wt�߮��8��t���=�ik~i��p��+���X�axGaʿ\`��Qt=*�)u�aq�c�TV�����Tʇ�/�'$�e>o{���$��>E�)&����i s�s���#������$4�ɻ�綐����~�t��Mq��"�6��4�fJ�B�k0ˈ̄4�~7<oc* O��K�������yy����x�P��U$���-�����{�l��6�O8j�h��~Rv2���7��w�*joVxw�JIv-v�b� ��2C�헬ۜD�w��i?C��R�����a�W�yѣ�r��=YA��OM��Kn 1��&"S��ˋ�+�GF��Y(���6�+f������3�4+k���
������%"?@���M�33#Kи�҅��D�(��icN��@�$e2���� 1�����q�{�	L5����U�o7����4�HZ�hH ��n���D��@zK��:�c�����(�읡9���xG���MF^%�dac�Vd��w��9�r>��5c�����ψ���U���C���j�� ��JO�j11#�p�ш�6yzV��z�ޑ�ۨ~�}�]?PFf'��_x��Yᨋ�2�
fg��M*��g|F��4+6�XWf�w�u����A)\p�jX���A��a9Gmы��b��06��GYU2��Ƒ������w[m���2�3?>l>m�iGP�z�;q����_�fP�^#�_T��}�ϣ���R���Ce|D��l���N�O\@P�e[A�#1+1*�Ő�{[�H��h�
��5)� ���w�ThW�]��G���OMKK"m����,��>S�\�9��x���}b��)�Aiv���;�R�e	d�Nq�}־�L��#a�D�K=�:�2a�PҏN}��3*```̋2�����7I�z�#�� �B��9����u�9]����W�͇�:ݝ���-y6�{� u�?:C�0G2F5G�OT��%4y�/�g�)6!�˽\�RM}� O��-Tc�ա)#Z��\){v���A\9W�h����.gͧ�¶�v�V��)2-nz���#J�z	c�t��ו���%���ș"��8J��Z���eP&���Uu!��$ ݃���>?<?5$!�l�A�lj��K`Eݮ���K������+�*�8dK�j/�ϔlb|�%v@���~9��9�+��м���	��H$�ԑ�MCR�g�Ġڍi��AV�)95�2���0�O���Z�|�csҚ�E�jk=ğlͨ��9�� 0��O#BXxȬ6��kq����Z� 4|���E�F#��x�x^O�0/(
�;�i���/+���E�&�
H[����Q��I�����7}�#��Z��b(,n�
M�o�i�$ �q��e��ԙ�ř��g/,x��р_��u��4	��V��Vs�LU�>�[@�2 J����v_��3�͆ǈ���Y��r�y�*���L*���[<�A�$+.v�U�h���kW�c�iW ���#;�M\���[CfO�D�>�R2=۴���6'��9P3L���C���ȂsÕ7
�T�%o��)^|rP!<�uN��x�A�p]����V� AIi�gΊ����#�x�ܸhx^1��FԹ��\$J[Z��5k%�N����O��O<I�n������i�7הC5[��:��׵�u0E4^z���������bn�U� "p
���~g���_^�Y�Ce�pi<������Y$^�ș?��5"��>�y4�bj�~��Ke�-=*�F�7G
6}��?_Ӿ�)���z� W���R��s!L�
&m��?�DWU���&a�s��)�K�.��L#���C������-��>q�	�п^�����j!������ć�"ѫ�zR�'Ȯׄ�� [����`��j�x̵|E���!��h��1 �ߕ%<J���W��y�Z���;|��<����G�랡�ܧR(��Z&I^���l�O�\!?�s��30�eb����.��8t�r�6/�B�r��*G�Y���Fk�%:�2�/aoރ���v��x�S�a.��sp[�U\A� ��B�J 2?Gh2O�	b��[�U?�Jj"��5l��f5��v��h��ȍ���5�lY[Zv����5�Cz����6��2��V%�AG@'}�A�}B9s�f��`�=���o��Tf�a2WS��4�t��h#����r0�\��X�v��"�6�{�*w".��i�Lg:J���w�GUcvYu�[�} �RU��	�6�y{�q�G��}��H9>b�+p��w���0�rWL����Rb߹o�1��*�6L-h۝��sb���o��n:֜w�����*�2͏u�k<�>��P���s�zEvw�kj|�E�ɥ+�t�Q�3���)����n��I�� �?���Q a���>#��^o+E1,�DbޜS��;$��҃t�s81��: �+��B��ю}�*/<\���F��68��:]q�����)xi𒸾�s��Su����׍�5֮�]��v�`C�j�ȫ��݁Y���OCs7��L��+���"�5^1���p�����z����vّ� ~���]�|�F�?s�7��Eԁ�����[ 
3 ̓�,"��#pFP�+\V�X=H�wN$��XԤAO�G�P�jfĺ�w٤�<~m����Ǣ��/'�m2��{�.�c�;�۝�]mrsF2�>?�={>��XG6;G���6�3RB_�������T���&$�@WQ&u��A��এn,�ZϜ+��O�&O=��R2�	��7�G�anXJ�Si���eD�E�F�4'�i�j���7�@��!5��<ŕ<�&����vpoZ��#�!0"�Z��	��t��Z
,;g��ffD�oq�|�"4�'���4�s����|��h���o�
�tڼ���~� �#�I�6
�Z|$+!������>��W�'75S!I�0w���U/gњx!t#�v�$����k����U�|���'�0�=a�$R�#���%�u0�4����]�>Ik�0�K�U�$zm!8���w�kK[g��;~�>���Έ���H�X{�u��gY���~�͉;�D�	��)ym�bH��C)8mh����K�/r��2�KE���K�v���U3�>��=vQ�
���c��>F7u╋PW(�D�;>���#��.Pz:�o*^ј�I�9	�D�I�~��ݛ���}�0el���9`�i쒽���*��ɉ��y��a����e�pg*��M7�9�6=HM?v���c�:�W��7���I��L��m��r?���D�[9��39��#�L�\�O�ީ�~�K�Ԧ��?�4C�B�^��u�J�j�v��Iy��j����c��:=���
4�D<+ �h�]���*��x��yEw�u�˨��j��� ���%�FH��H�4vZ��;<�y���Ԓy7m�Mڞa��4�(�+�Z�ȿ���l�����إ��ѽk�%���0���rQ84����q�B����9�YD�#F+�d�����"L�3���|���Cy��p�j����~�7Y8�4�\��0�����O�<������U�TsA��:hJ&�5�UxcF����.ƅb��J�L�W�	pV��_ru�ࠀ���w��,$f}�Ð��l��j�T0�_��Cd�N��S��R��9����U��l.�S���<�p�B\���
�'�¡9��~�)����O%�k��H[���龎(��*b���{ ���Lq��ۘî5e���$E4]�$��.�� d�E��}V�z�/�[ۅa�_���`!m��s׾��;��:�H?��zA�C�s���K��+#kK����� v�X�b�t�j�XE����b�!?���Ny��!f~�E���.찏��֡h����Js�m�Lƅ{&�|�׳.JZ*�@���_6 3�=Mm)�Q{5 ��͝(L��GU�N��׀��M�W���}�y2���;�U�f{��':sV&定/űưMG���yG����FN�%�<� ]]�(/"<g4kG�-���C�	�y�ʺ<-D>��&��/(���e��z���/S	���NR�p��\LZY�M��䞖�����㒇[5��H��(�Jp�Sm��>C~p�����SWNB�|?b������/�|?AwU���&ɰ؊�j��V7|�9��Ɍ1ma��V�lη�b��9\�ۛ�{N��DF�0$V^!';,�h?�b����^cQ��ף�E�(X���~h�g'�}�:���기<����0B���`
j8�zB}dC�B�^O;��N�W�թ؝��
rs�o�>\�;��I�gd�;/�+W��,\c���*�L���X1ޯL��d~�w	N�a�j�g�/O׾e[� %�1<v�{�ۤ�w.��#R�������������Bl�ʹ�C(,\���]��@}��~Kv&>H�v=��A�E�B	ar�!�SN���1�]�q:�����cN���@�r��x�^ȇ���F#�!��k}��Ǉο���ĹP"N�2Pv,��{�Z�m���Sq�޿^|߁=n�3&q7~�x�M��H)���Jkph����s�D�t5�&�MW}e98z;,W')�M�/!�0)s��z���������N7M�E��@]�k|��fi�qW_}ڀp��~��Mo�\�u:����'�����F�X�3?w��캂|�~��4���UԒ�'xd),�PNy�޸v7%�L�:�4������b>�����i�`����F�.-�_(�R�4�G�ܣ���8��sM� W�翱R�$�h����N�P`-�^-5`��@;ݵ��Z��Y��*s�I�zH�ٽ�B���#���)z��B��hb�xY%�Į�9�Bt�L����TPt����}�Q�P����r&�����<W 筴i� *�;��\�A+L�.��;���7 W��i��,���;��.�CwC��5D����pۍ�y��y'�o(Pl���U�C����%���Ti�<�v�^���PZקu����:�A�m�WF�/n�:���o������|Y�UoRx�������	E�Uo�[s.�#�%=����`�\^qIXPc��/C��N�P�q|KΩ���P>Y�t��a��i����b:|�`�����U�����o��G�8A�w^g�g�5&j�b�z���е�S_��˦������N� 7�nu��[�nx�B:E��HW6��r'��r! �?{%�ے����Z���;���͍�֒J˪��Zʞr�����(@LZW���Eb�lYѡ��Q��b��
��V�y�.��_�48�I���ABz#|��	,YU��F\ %KS���xo/���6�|�	^S�E^��͜[�\RǪ�(/� vVf?���h�S\	3-�[�J �[��3�l�w58�>v!�%hi���[v�&�Yln|�2b�m�5;*�������~��#9^�g�-�r~'Ω��	�s/�Y�$=_0�`��e|�ac/<�5�7�$���Sj�����Mo�i-9v� 5ׇx�� �.q�����:�ý���Xmmv��F[���ÿ򧚌��*F�qgh��n�HJ�G���7���m����И�����b�UN�B�*֒A~J|�X1bo�Ko��ny�w��}�%4>*�/0�ƌ.<�K����X���K)�w��<|b����`��Q"�?��:`�)����|t���y�1�?P�2Qq0�����#�5P����+e;,�b���3�Ì
�������8�?��=+�"��p^}��<���TFV��88eM]Bi���)��2���Ys�Z��1�ʩ�3�>gs�#Vߵ��`TM��nE�.��i7'C����?���	���g�!WX1�a)pfm˹o@zI��쑋 ��Z*~��;]�-F�D���A�������}A�V7
엓��k��G�F���+��)X�>(w�襠	+9A �f�A�owiX嵾+��im(�����G��3x��b�I�n�����v�Wd]Mhf5u��s��=H�'v��������?P���ͯ��X4đ�U-'�'�,_�y�hF�OP����¤��4V+����v� ��.���+�9��	F��$Әg�R/�~8G�<�6���6w/�T]�;��R�Z�2ݘ'��͑���(��_�@?+��b�zJ�BڼxNa��N[1�-+1��|�w1s��yPwέ�Y[�xWڔe�ck>d�h �'�%8(Ac�G̟�p��x��c�U��Kj��$ڜt!�=�}B~Ջ�p�}�o�����a�ʫ���D�=<��]��e^BQU�g��s./����Q��{��s$��EE-^��{�i�V����Td��2�$ 	�'i"�|�5�yb~�M{߹g����6��x�R�]B���t���K�~#Aqc���;�������y�2˭~�Pj�X�y{Υ�t���������cj�������2%}H2*�c�jۛw�=,v��)�8 VY2/?����D��~��0Ҍ�q�a������^�я]���Y-������7��1,=�	!�7���r�G��WYe���d�+Rz���33�Å4��F��E�vX����,�4@�/�Ṋ;3Yظ��ۅk�DB2ƍXNj�r@͇�ex�;���}1a$����H{�l!�E�1�[2,�=R(�4�h�#)�Zy�����,��K(���l���)�ɺ��	q59���xp�V��� ��	(���T����Mef�}NnX�×����ū'��J�Zw׈眭 �Nz�,3Ǚ�`	�O��ĨF�8I�M^���S �}��6c�z��u�>�\r�5sͤ3�:��ޙGv.ve��qHuN�: һG�<�FR��O��Ђ���0g���Bja��\|�k}�6�OS��T�R��&ё�`�A)�<Q�0�\�����":�K��ф�i')o@nWj<��ۏz&$1��4~���k��&���i��v.���"��eCPUr�#yo���4����'�5A|1��*'�W�j�q�K��뭅�j�3��r��SH���(8��Oj>y�1[�|���]��~��V�B�L�ż�q	GlH��j�%��R����Mi�M�Vb/&5�a�v;�A�Ċ��Y@hc�q6�b�zk�6�l*s��O
��L0��O ��xEy���[k�P�C����|;�}E�	���Ix���	��0-�]Է�8w;���j�V��4���8�!D���� ���mI�|�K,�b7y��d��7p����4Kʢٴp�ƫ�H��7ԎO1�N�cF� F	VӍ=�R��E۳_���h�f��s;v��dI����R9���a����`�p�-c���.˰�GW�� ���X�Ry �z�U��+�B�4 #./��f@z$�E�h��f>"�r1@��NB��Q��9�T����.2:�H�V�>�2�/ö�$���q> �g�i���*$�^���iAM�.����)��7W�W7i��M���;����Q�C��}D=�9@	�{�)SZ$'y%P�ª��rC�B�ȉ�E��TWǢ}��^EP�\�u�J��|A����`!��x��&Y��jR�Ʀxe㇪-ǯ�	��m�[��HD^%+*/���?��5I�X���=�ѡ����H�����l=��0�u7%M^a�ǿo��р����u����"�����0�����^}1�C,��p�|�����Q�UYk>���0�=��I!��A�"#;�U䧸'���!�J�2,�H^(�M
�]\�u�J)�|W���V�i�_������)S�wN$y�\�iol��2���_���d�r�i=���9�ś���l��2ps�Ϝ��5�,�'��#9���~�����e��(��k�u:c�0 ��Lc��=�@�^/� yAQ�́��昶�e�@$�q��7�j.� 7��E�S�BC��7z��[�ƺ�r?��Z���
��$��v�6H2�z���&�V�^��+�gԖ���S�"��q��g3��ZXƋ(��*bC��Ȁy���f�2E�.hK��P�{6`��b_s�����{�1|�[Z.TL��3�@��_�e��As)��{�7� ��f�����p`-U����J����)'���<�by%+�\c��:�U���h$'�w&#�/X��@���o�yGo^���R���}6<�V�]��o/��4^�(����C
	
�(�-gN< �F�
����ѭ�Մ����h��	�oPN��V����Z��
�R�:䑬��絸{��Ǩ���c���R�����#�h�ͅ5l��X�0�������#Eg�Ⴅ��ự5Js�+�Z��)Âx� �����K��Ɓ���J��M�'��\y���
K�����<������=��T(��Mq���2�q���I��6������.Z�_���q6.���CZ����K\�L�����ܲ�M�f�/��X��E�\O
K���Qn�W��\��J%�rf���X�}�@��~}DI�J�F``���t%�8�r�P�+�6�j~�j�!��|d�v�P	Į��c�o�Փ-Yk#��M��]>QW7А��L�����R��*E����u�}�f��3��	��;�G��7�Y`�*�?���d�n\of^a�K.�JxSVn�(���v�ca1,�v)�8P�2��O�y���EN΁`���6�o?R�SZ�8���D����)zRݿ�_��u^��g�o|���8��U,T��?�htt:P���_g��lᬃ�jo��'1#Ab|_�eWtF�o�Yw]V���εj/RR�A�����&��ɒQ�|�������A㹳~���މ�2�;(�Ղ�u��H�ΠN��m~�,��m�2i�6t�.(�7M��.����0�=Z6c��	��Ou����
I���>��=>�P�b��=5��9�i��3@�܃fl���:�_ԗ�H!�d(`ת�_��j7I`�=甁�+*n��5M\�e6!u��*v���)�nbX{��*�����A�J6��?�H~ ig����91*0z������YչS�Z,]赂�����AG�8�'"���uN{�`C��`,]��"_�/�e%.N�G7O����H�OieH��8�4+�D��eNS746�<�Y ����x�~ͽ%�Q��D����P�>����jŖ���E�r�:OVq�.����bZ������蒞X_�o����:ϗ�� ߙN���:�ip�\�=e��r�k�̸`Ѥ�	|ue�x�Lq)o�B��ü9��]�u�<*V���Aۜ)O�e�Z���
형ҹ�K��*�B�j
��}�ӷ��e�G�*;�F7���6��g?K:��ɂ�fsWH=��|��vsL�{�mqU�?�zD�.Α�-Z�߲5�ښ4�L?C��}���cٽ��{�*8�b���]�^Br�����j�� �uJ��B�0͋�k���O�*w��8X�)0���U�{�5��<�2��a��Ԥ6T�j�p�H���g砐��1I&��f�����xN����]gWܞ5�o�?��W|o"�-%�T�@��-��(�]��"a�/�1�.mBv7N���ܳ��ZO���m������DBSem�73��<��a���[�ML��Ұr=D�?�o�����I{D��
����k�VЂr�6�by>��3����� 9��U�:�������)]�m�
�9�pz��=$&I���Ō�1s�!Ndo#�C�W���R��G3 E��Ԏ��}/�a���! ���R�D��1�dc�	67��1D��I'�����3����0�y�y)��:;ߺ��=BQ4R�>���v`vEgʓ�y0���BgK�u6�%	{ST�TG4K4����?7QH�`�x��~S[��ȫ|�?K�d��W-"�nJ"�`�⊅����Lx�QQV��F��pzo-�?��E���_�����������r�n��I�	��}kH���^5�I:v�:��Y���(<��v�0�53VH�h�B�ہZ��� n����#/�e?&%��%.52B�P���?��Bn���S��<�������}�i�!��@�fi�]\̒�]�'����e*Ȱ���̏�ZƯ���|�"*B�Q����PZ��egG��f�3�o"���R��"�W�f14�N$���#|`�x�R�o���t�����| ��I4K 
�|�Y!�bֆ�l����7�Ix�w�Z��{��k#�X�$d�7�u]�?r��XV��0R��z?]#�0���=u���4������>��0 U)�Z¯Ȁ!��;�k��k�����Ϟ����G��LXQH	���]�IY���;��K���H<�x��ܖ)δ,h�"9�a�3rz�����!�v�[VU㥗>��b����� @f�9�&����˝T�f}����>��#0o�P�{�o �I(o9_�\�_�U���
�V[-�uM���X�eM�*�5T7��6+p:?͛^�Wr:�h4�W�31]���uL��m�H?:utD�y����0�!������\jL���=R��W�ҽ����,�����>+n^�+��pj�������؄��=�(�踕��ײ�w IG�K0���\x���E�i�r��o�L:? ��Q%ʴ��jt��"��Z���;*5|͊Q.����5ӞO>��~.�(6[�Z9l����lV�(�2���9տGw�Ӷ��K����8"vp��`UB�	��oY2lYF�M%hf�;�o���36zƦY�S۴�ҫ$w[a�1\oIvt�j��� s�?=Bph �N	-[*���xLH��ll�55�&v�+h�9�v�T����Y������ʜ*58���A������ω�򙐄���/� '+N*��9:s�K���=<��ݙ_�2Ka �w�����!��A���zs��)ۮʂ���Lv����6�阊�.�:ڻ:��:��T�:9��u�lvG�/[9�$����7���g0_qD�M��Y,Hg����tԔq�j�Cޠt������ׇbM�H�_��*��L�/�U��bJ�o���n�Ćw1�5�B��*����#�<���~�F��R�(wV��|(�^ɓ�sرQ��-�w��)k*2,�=�8g��`$?�۸Qn���;3�#
�ݢ��+��X,�wފ���#��}�x��8&���F�+�p��[|}���<-*�>F�8u�{]v��f`b)�A$����s[������FJN�{���\�
�2�8`q�R��������f�'C�č�����?�w�>�h1w�Cpú8�l9&z����ηّ�	~�
�]?�F�Gf��7���V�-� �Io
�,�=�3	F>%[+
*�X���w|�k�F1�A��c���"��r���5�Sm%˥���g�����H2�qߑ\�C�)6��KX�m��/2�Q#?s�S>AY@G��!��^�!�i_d3�L��3doT�2uQ�|G�K9L�[�ʺ�؃�!:��`cQT�F��cv��>i�ŁeB��;e�!i��f��K��b�r}���f���(vT�a���[��H�N��r���穁����Q���MM~)��-lժ	����0-��:���^��6�b-*C�-x�MZ��ͧ�H3��8��q/0�%b�YǬ�4t��6N�3��ݍ�b���������@���w^nJK�B��J�a��N�X�-`K����w��ˉ�:u�b�[<xډ��c +~d��K�\���Xx(V�IG���p��va�cQ��N���D�t��=��~��:p�J��dxS�>a��ʀ!�|�=+������SZ�*׌`���z�H��/e���f��{��L$��E:�8�^�"��i��ܨT���$�p��؋$ud2�Pw�z'����~����.���#^�6��ç�tB�}�	k�%)�~��c�c������X�\Ny���B�_P��Q�V����#8��D�Rk��2�j,���i�2T��z̥xI�j��hw��Iv�A���s �)�2����o�D���OM�"gͭV��E*���`�d�@ev�YBiZp�3�1!��l��l��G�G'/pY)���WM�+������3��C4����k�0��4:���FF�@D��ᮙ�3�F��-x-�@��D� m�=�NVS@"��em�u�\1�)c����{m2w6����:�߰�m�2����7�h�֚/���%eD�A0�K�����*���^�X�>@p9xn>x����t���k��XJ�������
e���NC�����a�z�hBO?�lO����NOM�3<TV`�P=����I�:��u� ,|�(����mu �����a\�Ije2�%�D>����̂�b�+�����n�J�qr���  C�Ky����2��?�`>�C�GD��ȯ����`_nx�TL���LT�ǻu�=G9*Le�h�j�H�#��!�M�� f7T6�O��;���u�!�����.�Z!	O�f0���Y�ra������h���K�:v���c��f�z~���!���o�r{EM�N��J��~����-(�}��#�"i�b��`CL��������z��5ㅯ%p0��.b��4�L�tAA!�=���}�-V)���[Pj.�z@T�@�M*J�L|�ma1a(�UN���- ^�AD�wF)5�.��L�[��f�)�c�	�d����c��:3B(��NG!��p�^	�=c�� �c���t63�=@��~*%�p�A~��>��a��7� h�ɀ=�c�6:jR�w�e�wK�<���u�/�l���{Hl�$��E��<�����ia ��� r��E��E[�$;�ɼ�ﶱx��Nc�~\���λ��ìF6E��GoB��˩	�śh~���c�[��s���K�W��)%yz����WP?1��܎Y������<C���!`�P�\j̍�ɿ�2���]U�x��CA��̻[��h�X.L 똍ER9���!3��z�![��I�&���L��Y�M��2��*��Hf~zH�l�Z���+�LT�J����=ǟ�'̛kq�X�������bw���|��y��fŶ�E�c".E���/-��&0s_[���{m8o|��^.z^&@�@�_�&��(�)8��{V�t )�ͤo猤8KUqs��~>��j�������3yY@��q��"�U�b@"E'�|�&L��/9�t���#�G���g���7<���]�J/i�4��܁4};�*� 	�#�a��<�{m�>O�v]���খ�Y��3�	UWN�E3�~+bZ�o����ūۖ��|{l���Ǘ|���5:�,L���H�h���5 ^���f��� <��Y7��:�Y�P���J'��+��F�q4N����;w��ԗ];�ӤJo�j�[T�\-�>�#�Y�m�p�/��;Z����gҡ(��Qqk�f2�]A�[��I�t�6�5����a_%]�q�x�;�8C��<wCK��L�����z��+��/�ٞXC8P���_K��~���O��\��C%���f3�<X�N�}���2�I�����w�3}%��H�Y���A�D�������~�*�k�E��b#c!}��Gb-����K�Q��Q�����و�H���dsR!���C�)߉}Ø;fnׄ�"(���W��K���*)R����´��"f��Kb��x�;�\�.�*��ae2�*��8�,gOuĭ���Lε=���k��9R|��l�>,����|�^R�+_��c^��TgP$��?�V�`�v,��sQdt(�ĕ�ageB�l솹�*�[�A�*��t�m�L�d+������i��/�"�Ae�8��N}<璅�Ds׮�"������l8�d)�f*(���ɩ��v���m2J�,�d���'�6��R(�-�M�C��5��S?���O+c�����~��4GǾ�����������ʭiw�j�d�+m��MӼ��_�bN~̾w@��X�(>��j�b ��y}G�f�]�E��.�h͏gق�r}	�Ɉ1sb�(���{0�|"��.��G�6@�#�_�r:���^)�^D{�� L)i�'yT��rYU��]�!}#�m���!����y|�FN��t#U�k��Cc'��&�D/�+���*�̕G��G����o?2<�SP]'$c/, �4��O�����;	S���<�����T�9v�����Js3�9�	��N�P�ہ��Z#�H�ɹ4��OԖĉ{�����i��:z����ݑ�>�㚇6h���5����o�V��z���,��\<��$F����#dJ���+�}����W�OF���̎s�ԗ pF�J�j�>&(\p���vˤ\y��(�e�S�}���F�(��Vq�42_'��^�+I63�6[�(���e�y_��q-�Y�ޯ�C�C�3K�"�L�s�!��d�e]��/e�%XFܬ���PK�w������Z\�u&%U�f�S>X�E4}JZ����&I�u�}���%���I������*���h�����igI�ĥ��c����3-�Ҹ�����Q���Q��˯
�)ivB��:�U����}�-�f��� ���2��F׫?�*��óL����:f���KE��xJ"ʗ�?��-f�aȈ7��T8����.�Đ���V�X�!��T�CbR?�p���������7��ER���_�_^L��gm��bl��o����,K�uJ,ź65����Kp%��|0S}nf<��gC�F**8�)�]�t�=��)]݃�=��s��:�=�}��ג?�ST�	��`(5�MQ�������Cت�,�|������^1X�p:.`��<z�����e~�@N]�/�FQO�\���
�x�dW��`j�
؊ �蔉��F��Z+���XB)w�VǠ]S�A����*K�d�	񾤬�m|�E��
�����|2�\ّ�z��2�����m7WA2(�d?�&�>8��G{y��� ��5,_�I���ګj��T��:uH�Gp�L|�<�a����7!�k��:�T���Z�_�	%�8 <��-�<�!�3f�r�Hyrt�=����<��J�e����������x��������MiD%`G��	HC��-�Ț���9&�b��C#�=դB&�B��񢋦��u�\�0յ�b���#7|t�A�mUg�J)(݄�5�9�r[�%�@+�����J�����a��N�bq-�8�[w=ۉ�WnΙ�1[/.ڀEec��d��o�ߙ�.�(�ZG��p��@mic(߷�7!���n�t:=��R~�ضp
h��[�b*��aБ.��֫�=�G�͔��TUQ�u�2�S���/�?tܽa�{�m�$
P�E1��s�{ٶ�iX��˗;�{����$$����%Ƕ��q�e%~S��ߥ9&�z�6��-þS�B��r��Ŝ���=~�1%c��Ð*��ⰶ�s�byѾ��-PVp�|�{�e�e�\x�����ir/��j؟�֬2�m�4����j��wܱv�2co�� B4�2�3o�ND�����ߌ9���M��!Q���m����ܑ]Y����ì���p1zJ%�#nD��X�G�ѻY�|a��i�+��|��͊3Z��4�9��k�b^��Q�}Hr@[~�ᥦ�3{�)��`�ס:D.�2�p���7#�(�!�V��Am��R`���@(TdZ�p�@�7l�������S�]Ч1���i�����8�g���B5�����	Y��1F7�7%�8��o"o*�x��ٻ��h/S����Is�[�2\��zR �󖇙 Ѡ�?[�h��B	��[�J����o��15l
@Q5�gOvܶDh�	������Y�tc��/��h��5�ʲ�_z��Y�X������h���'��\�I��s�Rrt֒=��;����a���0����_��nc��4.�(���T�vq.ׂZ���!/.׽��I<���v-�&۔�+�FZ��]����x�?�O&�M�3=�Ρ��͡	�RQr>�QS�U���J�RF��7��뿿2���g��������:�W���uR*����G�ym͋�:a0z��6�T��Q�u���:Gh�G��aF9]
O�*,�)۹}� g 0����TB\��b}���O�STg[����p�ǘ)��m��41\�D�l9��G�1ͫ
ٶ`��Z��)�Kn~����{ zť��4ۈζT˛��&�g��<l-Ʊ�,��6E�q�U��8����dQ�A���y5(�����E<!j �K��2�Ţ��r�!፮�ٿ��7�8h��j�N�Ϙ|�|6UD�q�{��=8������z	��H(��l�\R�L��$`Ni��V) 15���<W �����ր��c��:�I�k��Wl�3`%�%�0[�yO'�-xL���`�k��P��?g��c|��7E-g���xx�W��4��
$�8i��ҳ�w��sE@�
LPC)�s�YY0�Z�ٹ�s 7�0'�gӃ��,�OM�O}�z$$��q�ð�@��I�u�k�.,��/ф-�z��8h`���C�Z���Ѕ�>�˶aAJ�l���1'�7��K�k��T�q���f]��\��RX�ӻ٪X9n�%�[��*�S��Ӟ�����q?���"r-:�A��:���cɭ�J!rv�B�i~}�!F5g�:��0�ٿALi�?��ⱔQhĵf�Y�V3��*���׆#96
a�#'"f��C׽9�q&<�Z'�+�B�O�f�a�}���+3�lk��N;�� <�!��p���� &�6L�}H��V�/;M�Q���|�KA�L#?�IrV���HqLkm�7�ڦQ:9�Z��*��a �����V4�>�����p�Ԏ�J���)�>E)S{��� �#Xa�ӷ����A_ŀ���T�������rO�]/6�mA�m�C�Vn�^��Bɫ��(򊛅]�����\�TQwV�;P�#h��_���Ѱ�b�Q��N�(&it�F�Ǵ�4}=i����!�����W�B�}���
���HR}��B��Oߝ�N/.�WT����O
qso����2޻mWd`k;�O4�WY5\�=b��p�	��1�
�򪷸d"$�	rX���S�o�	!D$��1��v���Â��G�zȾ�2�@�aаd�0�[������ @��u8]�Td�-�"һ&bs>�V8=Ƌ;��*s	�\Nra�Sr����ၪ�y����K���;����@0��rQ�ׂ��9Im#�D�����T������e��G�P�i��bZ�t�̹��q�>�^ Do=���&UW��TJ�F_����ko�&�s@�t1�&yϵ�h8�1WKNހ�=~!YNs��D��a�ō����;Mx$��d|��)�sT���q{>�$�Ի�[tMG+����|���'G����[��R�?�=�^)���)�4/��U�f'��,��\y�����}�-W�¯��4�F���{ơr�@�+���Ej<m�F�q����R䤈۩gs�ǹ��i+sq���vw��*��ȫ7�ȁ5��1`Q�/-ٝ��d-Y�= U��d���v���|z����_BX>)#CfY����zںއ�<|���y�h��]�B诧#H�T�r������t�|�%#H���Dሦ� Li��1*��x�8��AO\T.��_s��{bW��i��8�ѵI;c�F�07�C�CLD������۱4�I�'��P�k��-�C�dc�?Xȕ���T�-@s^��P��ru�۾�{`A����?t�S�ޝ�⤶/�����x𰪣j�@���	[�Y����%ag������{"I�8��%�ї	��t�� ?��#����Iu���^��f��YG�v^T�2b�"�|!��@'�D�^�:CbRup��::�ǧqY�����(�0�������%�k�Բ�������W��J�n_���_��ӝ��k��J��W$|�Vհ_����I���z��㦍�/i���F��y�,bmѪ��`Wŝ���9��n���t>�����J����
B��Ë���/k����L·'���Yʏ�xr�ӡ8�XߩJ%&f�Pe���5 �G/�ײC�j�r����B�:�������2Ar�_�"~<#���.�:U�4���LOO$�$���{��;�<$T����=I�_E7a}�"d���\9�N=&"Q��I�LO�;�a�']�{��3L��8֥;��6<���T?5���� �L��SHqF��|qw;3���{���LI�����-O@�X�c94x��[X���p$G���
��tF�r��N�Hk����0�5\���"���YY��[��P��i7�{-	M��.K�a�J���nȽdϸ�����&k\�+M2�d�IQؼc��n�:qS������u�as����i�w�r-�@�8D�x��Xg6��x��B�ȶ�Y�~�ZLw��=5f"0�k� Z&_gMj�f`��o��$�l�"�v}�׭$4$���H|fp���oE��t�yO� � ��I���
�E�|�y�!����Zֹ����7Q#,I�܎��Tˑ����a#c�k$�!���z�����0�ʸ0XD��@,�#t+
���Gu��4�j"�"�E>ej0&.�U�O"�5t2!T����kg?��m��0n�ϤZΤ���ygX�JS�����i�	;O��U�Eg���Ƥ��6)ԥ�h�4Ǳ��r��
�绋���v4y4U)t9>�>�Yn
�����"�ژ��������`;->� #�L�PLoF)D�Ox�9%ߖ��:���]�7�✙I�e�M��`
�����4�*�����fZ��'ge; s*�d�7l �6Y8?�s�H��ֿ�W��5�e��LU��m��?([�D3@���	�O����2�
۔L�[�k���E��gm��d��T�,f^���YŌj�D���
���#�~�ǋV����
��`/ �A��y������x�јE-y��]F�np Uũ��"�1H��?�:�����	�)���l~w_@�)�ll0I�VF���< ]X��\�۬`��u�����2'͊�:@:Ι�V�RL���u���:�u>G�L�F8��O|����o��g��J�~i�P0\�`�}��?O��eT&?�LJ��Fh�)^����\�W!k�D�&��j=3��qٍ�)�8n�I��=3z��R �
��ԟ�mВ�|��{h�4�����(�kl��A�U�� 	���f�%Z|�35'/��i:\�j��K���ݑ $�Џ��@�x�����JlF�@vW���3Y�~ܭm8�=����Bz���TYUMF\C%K�뭊o/��6E-�	I�S��]��x�[�
\R2j�����R v�q?��#h�v	3�R[�U��[h��3�Ol��58}�v!�]hi9��U�& �Ylٱ�2-ãm015;��������}'#D�g%��rI�'��O��s/�Y�=_ۚ`�!e�Qac�T�5j�$����	S�M�����MzZ�i�v���ׇ�
雋�.\Ի�&:�\ý��X؎v�Z�[�9��J ��w��*�dqg��n�HJB����7ľ�mqm��#И����åb�`$�BO&*�]�~u��X�bo��o�8wn$�w��.�%�*��O�ƷG<�����X윥K�Bw���|���֔Q�Z?���:��)�o'�����Q��1��?P�AQq�����<#̀���ny+p},��3����Ì5�����8����re+�*?���}w~<�.�/�FVn�88��]B�����)��+�髀s���漚ʩ���>���sߵ��`T�D��9�.��iC���Ǌ��@�����!��1�,�pf���o��zI�,����>~���]���F����l���t���h)��
�&���ϔ���F��m+��X�əw��H�	v9A �p�A��w�x嵉Y�ؔ m(V�x�G���>��2s�&�?iu�l����m�C2T�?6!�>d1G'�*����d�Z_ЧO�g����T��Iut��GF'L�f�b��&x�!=�B��g�TY׷�����6��d��8v1��!lW:f�}��r��n��,�'���ٓ=��K�)ݻ������R�Y��̊M���Q�qխ�zK���Yv-��9�l>�eMub` �CO���P*��nѻ��%��������0I�b@��OE�t�4��,����ݰ�q���۴�ZP��!@WC҉z��J����M�a�\�Ns�-C�c䉹wI#������[�Qڬac��~d��^8�c�=��(Y��G�M�p�0����c�l��cd�<Xt9��=�`�~���p��ە��D�1�a�@^�Æ����=.�x���u_M}"oZ�)� eʋ�0/�9�i�:{?$�F��ʋwXw��C��r������a�����.�*		�̈PGk6�Qd5V$�6& �IY�����v��6z}��5�S�()���t2�v��n���ϲ��%lR&�M���0h2"仃�>���n�(BS���19��>�Ȋ@SiƮû��d@G1���i�Rf��V�ּ�%�p�j_Z�����"�$\�Jx8Z��?g�fZβo���C"��ч�` 4^��ӊ��| ��z�o3�tp ��4� ��
I�]5
`y�|zD!���H���6�֭7�7K��I�Jo�7Q�N7���#��K$$\���W�����Rs���0��:�#��>�u
u��4����\c>�+W0�hU�Wd�o{�!νڊ͝ka�$����ª	��^e=Ξ�_׳�2X��U� �	�6��{�;}�<�_z�?##�8��V�)��Fh�]��!;Qr:����ˉ�CvnNU���>I+��S� ���J��K�������&0�ڑ�>ED�#�)�PP�o�,N�	��9�/�DP%Q���;���/eB���q>�������X�*ɕ��T#K� ���!�Deu�*%Q7&�:6S�	?���,�3�W��Yd��>jLA�mۿ�?b2�D��Z��w|�IB���ڄF~L9�r�e���%�ᩳ�T����f�2^,·��Gj�д�%� 7Ц8��P�L��"���NC qP��s��� ��x"�E�O���͗�:th� �%�q���X�J��Z��;Ra#Ͳ����]�P�w>ڧ�3�(^Z<(�ʌpl~LH��Ǵ.������c��s@��Du�8J����a/B?�#�@w�YZ��Fn%���z�o�1e�[�6��'SH6��u[���\�����[� �� ��q?e�!hH�.	8�[RO�ࠖ���ql��5]� v�IAh�����N����Y�|&�9̣�[5`N��iw�������*��=��Wj�'S)��s�����=dS17��tfaH0�����I뎪i�t�U6��i����썮��v�E�K���#%.����b;�: |$�b&�ĝO�vo��[ae|��7ϧ_	,Џ[�ql*���H�.��&�Լ�D�����Ȃt��R0��3bu-[���6*���<H�}3{b4 �o-�n�[wYm��ju|*�6�K3<�ۦ�\��uҥP�)w~K�|PHɻH�4�Q7�3����)�Z�T���<���,?���Q�Q��c�#24��܎M+���,�޲ܻ��/�����d8GA����+E ��h}�i?<U~�8o�F��8���]G��ʎ�)��γds��R��n�ף$�ք�!�Zd)`�L^��VS�������NC���,���4�gA��f˿1�^p�Ṕ
�z����rD��.�~%0�];	SF�V���ݹ���U��q�j
	�:�e�o���oFf܏+2ƃXӲ�w�Ꭰn<AA%'q����<�����]"mmM���z⠬M]�C`�2����FY�Q=X�sDhmJ�2�?��>i9G�l2�7c��IA�_���tߟ�[�Tuy�G���L�-����ث$�!b���I�T��W���N�f~�ũ�;E���!��f�x�� �*r�N���I��Pب��Y�����p���,헩���������UM�x��a����az�,3-����� ���bE$�C�	�u�]�3������茯�& 0FYb%����z[t���^I&�[��ݵc���Qٴ����>@�-t���Js`ڼ��Qa��N^--��N��w����iΊg�[@�ڱ;Mc(��d:.� ���7(~��G�׀p�q���cy\��H>�!��t���=ȚE~�Pp�V���*{�PaA��ʨo��zX=SF��m��KH����1���ο�p�/�I�܎�p{Ч�$�%Eb(�ī�J��i��[�|�K�L8��͞�$��H�D@_�9o��*1~�,�V���K�F6�����Wn��FV&(�foߝ(����S^RҎr�[���\��w���[� 6�?`.=h� �	��[mG���$���|l�N�5�N�v�h)^��Y����[Y,�G��N�-��5�F%�d��`]Ƕu��'�a�2+�'��Ԯ�s��=�f �l%Qa#�3����乑�dS�7'�yv�l��)�~v�--�G=��[]n.�e2��GE:�d�}����[vJ|�[�b爃ܙ�ZAK�ꒉq'M��.iyH
���B���
�-�<�Å��X���u��b�����*���>OD���b/�'ow��n��Twt����Ȧ*�\���Q<���ۡ�*�.S�N�w��|˶�ɖ���]�Q�>��u����)N�co��������I?�Q1S�^�#�B��h3+ǡv,�7Sލ���L��@���S8�z���+]+`.�h�}���<�ȁ� �Fx�8��]��ʩt�)I�f���s��:�N��i����Z�?'�u6�`b������� �)C�m�L�h:�߂�e��+1zΩp&rY�/�]z	�!�QX�����~@�
]���F�q(�H?�vFK�Pr���� 
����O˔u�=FA�+mG�Xn[�w����w#A�͚� 7~�uk�1m�=���������U23�͑���,Y3ۮۦm�ȭ2:_?��>$�G���Ȳ:��$�_�iTɧ�V�Tg��u4:gG��yLhP��̓����G!�4�1'T�8�FYL恨��$�Ȯ�W���!,�ef�+�{�>r`����^�ːM�d!+�����1C��&a*کd�'��M�u��M��a0�mX������-ki��,���%7Ub B�C�"����.���]'�x�����0��	b �s�_�tdg6Y(y��Yt�p���1�^�K�v�@O�:�Jn
.�P�akmN3
�-%��w	���Q�p΅܃[����l��cCod��u��W���G(@	G��ph2`Y�nc��u�#*���1t���=c��~�[�pvHP�G�Q�cNH�#\fZ[�vc���F��@%�y)-x̰���>֚`����Z�乕��"��$oݾ�h�Z~�~g�bf���o )D���"(�1�/�e4|i��hmB|�@f�p�6o��8tN�L�x� �^�Id
>C|"�!+���-#���Kܬ7��PI鎔��#���*�#���$���_���]c��p���wN0���ј�o#����S�$u$�|4���z#�>���0~^�UG�Rj!�@#�k|ak�f��ŵ�� ��b �����ќ�X�'��E�g����;[����5��R�VN�4%
),�h)�?� r�?�?tb�?Y�v���U�me>�C韱��J�����2)��#��D���	>�V#N�Pn�o��ؘ���9}RP�=��Aݏ�;��!e`�,�O�Ҙ]7]���*�R�2����;�e�"�*�7�8�6�%]?ؐ   �  v  �  �  �%  �.  K5  �;  �A  H  aN  �T  �Z  *a  ng  �m  �s  2z  t�  ��  ��  >�  ��  ğ  �  ͭ  �  ��  h�  ��  &�  ��  ��  @�  H�   Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�� |d��"O
`�(�;���8���-0��1%"Oj4��ND^[��"3/9�0|H�"OB���H��*�ʞRy=a"O�味V�!X��!&F�:J�$���"O,��a
���C�Ą�M�"O,$3%o�-���p���+Ն�:1"O��ݢ1����`���y14]2��i�<�6��{_���c�H�`�fX�$Kn�<��A̼VI�xR[�)�Ć�pඤ�ȓA5��('nߡ4�� �)˩%� ���,��r�؊b#`T�eT09���ȓ!�b��g��}�8�F��-? �ȓ
K|m�ș�VṔ���2�%�ȓ"R�X�j�4JN�1�˘X�i����̹	_�jZ��1!g��zܶ��ȓgil,*�J�
j�Ne��i�J%b���f	�(U��:���G��$Y^م�~r�� S�%T"���k\�jx�ȓ|4�1�îJb��@ӵ�ݩn�V��/[`�"�v4�R�!ʎ<��M�ȓ`:��z�ؚh�J�Z��$HY:	��H��p�m�C1��!��B:��0��EnjZA V;9����J[
2���	��4'J�EA�IVW&��~�(aZ��ӹ�>� o�Y�|�ȓ�f�A�
Ο7�H��M�$�����mޠP����/���ANXo*�ȓTv�����{ ��-7�*h��I��sB�8�8���3����ȓNe*M�悡;������X�o��!�ȓ'lj�#F�m�+R&;�|��2)n�C��0S4���T:
b���:�0!��e֊��)��ͷV��,�ȓ0�&�8#���� ع�L�����;�P�AFd���,w�6d��r�EQ�( �gVlɦ�M,H��,DP���|�I	$G#\���ȓ"�)���E�B	yt&B�^�LɅ��|��B�,�r�Ռu3�h�C��'8!�D_��p-���K$��aU�/ �O@�	i�OOx�h��	:T�)�"��,n:�;�'�ś ֬y0<�Ɂ�މu\�	)�'C �8�:\[B��@�׵olV��
�'(��#t.\Q֕����c3��q�'�F|#�άt1�@+ 
�-W�Ɉ�'�|�Q��I�A��A�Q	5�d��'EXհ��IB�k�	K�PV�%I��hO�!�s+�'\�F���ز=����"O�Pr��� +�Q[2�[�_�� ��"Ov4�m�?Vd݆p:D�D"O�3��S�( ���1qZ��Q�>yG�'�j�AF�O��4���E�5�t��'Q��4hV�0i�tK��*��m:�'�K�N2��F!�9��hê�\����?�'%��)&Β�C´�;@�C%IK�a�ȓ`��s���8!m��Ks�%�t�Ў��s���Ū�1|_��z�%�"e:"���4D����Ƣ]!.�c׋X
[��Zu�����xbB�6����MT��
�� ؏�y2�*=2D�w���2��5�*��y�?@��2�r@@0�X6�y
� �E��U�x��\z��P+E<b�"O�0�䌆�n[�!�� �Tx��d&LO���h��Ԩx��E-�BG"O�D�������Mb��XL1�"O�	�F��;(�bhc�-��H \�"On%a��Y�l�{$���BS�"O�ఢ#̷F�0 �G+�VX�"O^���Æ�u�n���Ɉ: @�I�"Ot�!�'BR��F^�P:� ��"O�x�ь�(v(���{6���"OLH���Ti��a�dU*'�'�!���kP���^\��'� L�!��[5	�V����:GPƠ��e�Q�!��$
�
�"�Zi<`�G��.'�!�d)Bà4�cD����<!��� �!��1E)�)�ի�':昌�̘#o�!�dN�|4X�����W�M3��k�!�$��DX����-���VK��?�!���X���`# I���_#+�!�d�)%_�ʆ�f

*�P�2C!�$Yh�|\�`��� �Z����=!�ı�n�7F�0{�xu��M�<a:!��* �6Ҳ�]:�x4��!!k�!�DDL��y���Xl�Q��ͯYta}�>Q <hwR�X�%Ym|,[�NA�<��FT�(�� �J>v:Ț�LM~�<�"�N{\!J�#;5>&�$�Iw�<�GZ�F�Dzgჹ(�v!�t�p�<�Aj��e��,9��5}:�d��h�<y'l�]&
�1$�q�i9���c}
���hO��b��1^h@SV��>3��g�'�MP�0A2MB�Ni�����1KF���>��`���j���|6��s/�30�	��J�0H����+����glΕz�"̇ȓm�2\��L�x��\YwKő2OZ��<y���	 7��L���
u����a�k�!�$�g��e`	�9�i�� �n�➟����锅0�t�:c̊@����2���C3!�$�� �~��T+�6��uH7&��Q��/e���N��V�n5� ��)MZ�͇ȓ]�.��M�������@�IM�����z�E,f���9R��.9��s��)�}�Gԛ���$.3����C�y��	@lY��d%-V&Y����y"ݛVd&�������TPg���y���%mB�`��GS z%�uK@ȅ��y�葎�=��L��C#Ԣ�>�yB��l�|���i��?Ĺimޛ�ybo�o�d�Q���+:b|<�U���$�O��"}�E�VWB�ု�.��� ,@a�<�'jަF�7�ս}S֙j'.y���=��� d�ZP��n�9/�Vi*�SL�<1�鐡S�ʨ��E9��T2 ��|�<I�i^�%�>@ ��3o8��e(�w���?Y�W7U����)Ӳ!Z����z�<�G��U��j�L5NH��2T�,����N�����Z#�$[$�9D��s�ʑ8n�
-�Y-����/"�Iz���)�[x
@H���EA��d"D�x*螙HU���'^�Q�ƜR�o>D��[5H�q��iR��-��ibi/O"=Q6��\�y��bԺMw�հq�u�<		C\�z�WO�/��A�5��h��hO1�^0�"\>�T�'�
$��"O�  =�r��xN�1���>�1��IyX���q��<6�B}Cw�"tM��Q*:D�D"6�_m/t!�b�#��>D�����P
����uB7���O;\O<c��W�;t�ZMU���4��2�h9D��2��N*O��t��KԵhɶ	"��7�	]���'b�6y(6�mwJ����ߵ1�lX��*L=��ʂ�W�����k�1m ���6�\h�S���k�Q�%�)i�!�ȓ/����l�r����3��0cI���O',S����V/j���ɭ  �P�ȓG�H�FÙ�M�D�׀�2����>߰��,�TJ�I�w�[�v1D��<�����ӻ-����'�ۆ�>t��'Q�E�!���DfNd�W@�y��ђ�!�e_!�dR�^����;p� �@c�0P�!򄆗e(� 
Ãٱ>�TBGb�	]�!�;n� b.�6�I+u��G!�@<�Xce�1!�dU��	�R4!�DVD�R�#�B�E������~|!���9_�$}aFOڵL�pϋ�s\!��ܯRT4�&����$:���ML!��G�-,�e��j�і^=�t�s2!��$���Zv(M+6�*�l�Y�!�U�yF�X{�E�(:"��9Gl�|!��-r�<ate���(F�$�!�d�'J�L�W)J8l�*ؑ��I�!�d�G�X��M�L��I��)�8Bt!�	�z�;�^�
�� Wd�0s�'���%�=-+ΐ��-�w[���'�Nq�g��^|�EG�&q�"�
�'�����J(pUd��g؞d,���'4�ЃRD�#kĞ��t�U#V��<P�'�V�D�	<`����K��0��'WJ�`@LW��p ���s�;�G�<��+��@6ё�&�+�f����F�<ɰ�=N�"�B�	rH(E�UA�f�<!��6W\��f��6vz�Ѥcw�<Y)I/V�*�ȒH��^dPE��k�<����U��C1��ҤX��Ag�<A��?B�^�#�w���g�a�<q�Y�.�����1PO^(�R��[�<�Fd	xQR����O,�8%Hb
X�<�)G^��!�R�|�G`}�<)#�9�l�l��bi\H�v�^y�<q�K��s2$�0�j�5�@L�1�XQ�<Y]yG� '�ܶii��4h�j%!�D�
� ( ���6	�C�ªg�!�Ć#H�Y�2F�
�E0`�dJ!�DP�=���Z��8~���5P�!�D� �,��t�*�����m�!�+�|2��P��uصP��!�D�2��I�H<L�Z,pwL��p!�d�E|T��CL�J̓%�Ƣq1!�;4*�����[���`�G	�01!�d92�8��F�JH4�;��WW:!�3b���O_�73N�K�S�s�!�D̵i���ku�ǩS(n���8+!�d˽]Z�D[햻p��Q���T�!�$�i�<��mι �\a�-D�m�!򤆫	Ǆ�C�C�(��QE-�0Wi!�dªc�0�[�9�fh�t�=!�dK�]'�麀���}�J�*c��`X!�d�l�����b�⼻��@�2?!�� X,����� 	��+�h@��"O ���rZ`��G����	�"O�!��Nױ{��E+^9LC�0�"O�u%�SUE�{�ކ(/�� "O�4��j�WE�|3�ǅ�j<�]8��'�B�'l��'��'ZR�'�'�Zl��R'$�\P��'2U"h���'d��'pr�'B�'�B�'Cb�'u�d���ԾvR����E�tp4(#�'#��'-B�'���'j��'F��'/��2-��i�V�+���;[����'�R�'0��'���'���'Qb�'��LY���r��gW�"�ՐC�'��'���'��'t�'��'x!��JܒH�
�#���fl\ ��'���':2�'�'�r�'l2�'��u�W��>&adCϋ%D@=#��'�2�'�'~��'�'N2�'�ܰ��T� �x���6Qr�\���'���';r�'(b�'b�'xR�'��X�OɨZ��!��A8f��9�'�'�2�''B�'K��'l��'�dJq ` �9oQ/\��(��'��'���'��'vr�'VB�'u(�J�d�"�U�$����'���'���'(2�'Rb�'R�'�^H�F�#��sސ0�t�'B�'��'0��'��'��'q����,�ѲQ�T��7N1U�'���'�"�'Bb�'o��b�����O�hru�D�N2��R���!�� *�fy��'��)�3?!Կiڭ��M��FCp���`d�4�S��	��禹�	I�i>�	ٟ��)"H(,��E�N/kG2�J�ERџt�I0r��oZO~9�xU��Q�)ی\�~�S1+p�c Ù[}1Or��<��	�>0����U��-L,13f�=d|�n0Q��c����U��y��I I,DX��D�vp�$�[p,�?a���y2T�b>}�����͓^)
�iƢٻlR��U��"X�yϓ�y��O,���4�x�dT�� �#B�.�pA�d�[���$�<�M>y4�izv�яyB$u5n��W��!z��	���IE�O�@�'uR�'o�D�|�4!�?&w�Q�A�P�`�qW`/?���B������W̧B������?Q�b��-����� �DOv"�g�����<)�S��yb�^@�z�"�8N6�)�S 7�y"`~�<Dxe��l�ߴ�����j�?7��$)���@0MS�'�y��'o��'+ni��iJ�	�|���O��\��ׁ�hyZbY&~�Ԭ�aH/D�`�c���\�H s�l�t��);D���FnI�f�Xy��KAw�(sQd�o���&�<D�7��5Y��Y�o�w����IDc?ƈ3�f�s��d+��	ou6-��AH�`�R��@G_�\5�IQ�މnq�T�&��h��j�C-�MHWDM�t���EX�@�逤d�}�nX�!+еP��d�l�s=&�	Dlɪ �����	5x�iB� Vg��)ɞ"�C�I�:���� g�a�V���
�b�ɃK\-crePe��d풀� ���*��e�q�QK�`藭�X	H�*,�,)m+!d��Q�q�Z��ˉIx}f�H+�A *�,���*zj� i��yycT�
�`>����,3��%"�N�\�@�4&@US~�3�/Y�'K(� �/AןL���4�	4�u�'^2Ň"M~��30#��#u=S˞�C=�����O?:(��K���;C�"���O&�����Y̓�p�a1W$d���H���s�L'��BC�5��=���mB��֘~r`��>u��D�L�b���Gʮ'�� ��Uu����<SR�'(b�ħ|j��
�~b�� �,p��Yi��Vi�<!u�^,YX�:��'R�ʠ
�L�-����S֟|�'��t���l��``lD*�jɻg�0T�^����Or�d�Of�d�������O��e�h��C���<%�T���f�!�
C�dɢ�型|1]�"�'x�e��LH��	7��D>�mwĆy�2�0��D4�(0w�q(�8�t)��'�i�=��C�ӟx�	/�y[�Ƅ,d�T�cE�N�d1�Iw��h����(���X�+Y{n�EC��+V�!��#V���e'�j��x$"�a���W�����C�S�O2Xuz�\��ĀB��0j�p�'9&,��U��ճT�ø�JD��'/ 0��lW�#㐅�3��0pt��
�'�΄�T]!E�F�r[�S,�̃	�'_4��#Oǈ䶝��b��@X�	�'[�E���]=(�.�.ԄeQ#���y��ˎVA��aR#�=-�u���y�#F���c�M1#Դp#��;�yB)�Q�,��u���z�a�E�(�yb+V	��&�Ҝ^�t�Ō��y��@�ĥ���=P�\|���Τ�yb	_�ʥ���67Dh\B��.�y"g 7�� �ʞ+2}K����y���z�D&�83pڱa ���y
� 4�p)ߐ/��xR$��; rt(C"O`y��'7v����lɱB�j��2"O��A,O�x�K��7c�ذ�"O��F@@�X�a��$��ju�v"O�0�F4̞	��E�,��"O� b�/N�>�hbC�/,���f"Oh 9`�Ơ��ʒA�-,�j)ʓ"O�1RB,N?�h�2�!��%N\u�"O �I�'#�i����ي�"O>�i!F\�V@|�".�4P�"OV�F��8�l��/��G"O�tz�E�> �s�ēA%tDIV"O>!��HݹQ�����Ⱥ`ī�$"OHJRKRA�t`S&A�7u* <��"O�m�ċ�.�<�:�ʙ�t�%�"O�d�2h�+'����JN�0&�R�O��W�׋(��;6�V�V�
�K5�F�<�6��=%�1�E��4ӆ����NE�'���j�(�S-0��U�C��u����cX���B䉪C˞؈�۰+˜�������8\�\�>��<E�I޺Q����!\� ]�Ê�.�y�iT�H��h���َ���Fh��]F�p5O��j��^!-6��I?�4��)V�uۊ����˒=�`�Ӑ.!�O�hJ���1HP��# �tLX�p�#~/J)�`�%~��IÌ�jX��z�MV-2x32��!2@��`�(�o��H��U&/�F��5L(Y���
Z�"UA�a
Y��RB��"C\Lا�	`4�H3�F9�%1O&�QA�Z�a�����a��M�?qY�OQ4 'zyH�GK�P��0Sd3D��3jG�s��1���Y7��؇�s!v:3��J��t��=H8ʧ�OxD�"%�*���*Cc3w�c�'ni)��HҤh'oL(09.qQC*�e�@�� ��6rƅ ��7u$���d�2�A�Ƙ.	aКǩ� Cl��`�h9>�[gD��p�h��Pap���܃ _���bA@�LG�i@�a�iL!�$�s�� 	�G�A�B�9ǟ�`2"��p�DL &Խc���"+�1����)
���,���
�#X�S{� ��#D�09�M[�>h ȿ��%i�e�s��%��4m�����d�M��Or���gՠ<����_rb�LAd�'�!��kNl!2q�X���Tmޢ*��x"�Sǰ@�Q�.�O��(����nj<5B�ɒp8�U�A�	]E���E����![ט��	A���1�A@'��9�Q�H�!򄇚$FĠ�G����!	� %�dT,:>z�KaO�^�R&��z�O
,���u�-SȜ�5[0x�'��``S�V�n��(�D�@�̩�ƥ&vj6��S��i���US�3�8����L�S����/�����I�2�`t��\A��!�:f����1v:J����:�����I�s�$���jT��~�3�0XB�=	���	��&U���ORjiaaӞP.���E��	K��J�'#�����Աh���!���#q ޡ2޴{���8ň�y�4yy(O?7� �E��<�ڳd�h�3-ͺ-�!�E�2�8�۲��!>	�x�s� nA�ɶ5��K��#lO�B'��d.�U@զ��F	���'������<h���`9J�`���
P�`�'D�� N�wU
�1 %G1u0@�.3�7\���I��v2��0�ݤM7:u괏��	h!�$K�J$�H� �0)r%�;lb�V��<S�c�"~nZ�4V�B��7Lx�7eM�C�I��	ɂ�y����gްZ����8�A� 6|O����HZ>J^5Zb��,���;Q�'����s��M��l��2稉V�P6~�ҩ��VS�<�'!S���������l��Q�'Ȍ�!C)O�Q>�X fɒ:^��h���h���
*D��AH�tT8�zr/ϊkJ��Hq��Ot�IC�C�gw�O?�8ccN[_։ғH4W�l1�DZ(<�5/4W�d��I�?��0��ڮb��@�OX	d �U��� �@c��V8I�i��#W�JU�1���'7°J�F#?��,6����.�,p~�a�V>x�8��V"O�y�D��Df���!J�,7�)���CMS���$�s�0G�����Y�d��$��+>������yb�E�'���W��v�2�rg�����̟*U��i��k���~�<�r�rM ಶ��8Q|r��ōY<�v�<$`�u)�䈈P��	V`ĺAN
dA^�Lx .H�Qkaz�@!7vz���EI�j���bW`���0<�׫�=m����^�Tp�  0���	[1f�Y	W���y���
|%���qB8/���V�����(0���'��&��B�~ڕ�uU���Ɵ�(���6�H�<Y拖�*� ���ŋ�2����O}i�?�^}j�'n|c>7-)q��S(�"x��k�D�.40$g�;V7fB�IG`"�{��Rr����*HFu�V\�FH~Ӹ-�$吪A�R�Sa�|�?�A��2� q%�c0�!��EL�\�I����X�V�xс ��p,vd�'��Rx�$C�@�P	�jW�92|�#Q�'��t0�U�7�,ф��:;�H*(O�Yi�L��?�&�v��Eb[���g���d�I���3P�Jp@m8�	��yr�Ӫ`���9�ؖ&�F��<{W>�£��S_��9v�T?mkd�� ,��}޹���
�$i.T(�� ��w����dLW�US��� &S���Pc�}�P�J���Ц��'�jm��'
�)pt��{�1���-{JZ	3r�R��=����/��-E~�B��s����ɽ-�~p�bf��MAD�	^�{%�[?j�@C��P����(��r���)���r/B/��AJW�wNj�8�z��5Oz�qVK�4��	 \$t�i>鲑�Rsግ��m����Qk��$D�<9D�_������ѵJ�l0��oͳD���E�'o��q���~z��J��9��I��ɥg�*���� �x����'��Y���!�${�g7���:e�_�!���.��O�<�ቹ,ňA��V�xe���|�#?)BZ}��$S�NP���O��l*$��2���ȶFv���b�O�����'�y��ua���ӄn��|��OH�	'ȵo&u3��۵BC���4�`42d�ܲ";���g�X�v`�ia�"O��Ģ����>����ra����a�:��Ѥ�^�m��T?O�Β�O �ػЭ!��8(�MNu}a���=@�RӄYi��ڒ"�1ְ� Su͘扈��'��<���>��a��{1&���+�q����3dD�-;��݉5)�Y��1�X@�%f�	b�4уE+?���Oą��I�|�.�#3��_B:�8d�R8qM�ż����[i&(^^�O�����߶\�DP dfE����'�!`�H@�n�()%+Y��#"6
d�I1�MS�*����gܓ@Rܹe�%R��T+�	�ȓ2V�T2��;b}�=h+A�:�R�mڹ
�<�sC�P8��c�
%F\���@�_�4x�pb*(|O��J�G+g&�牆�
�B �����X%H��~B�	"�B�j���Xc@�}�l����'�-n�\�F�d�K��]��
�f���K�r3�'P��{a͙�k�5fN�[)���H�WV���J<!��>!pD@��||��X ��$h �OL�<�E ��ij,e��$��D8���KRȦa�7E��l��e	�J�Q�D^�"E�,�ĮW�a"`����"	lz�"
��<5�ːy�(�k ��<�0�,�O�<���k�Tu�#��Gs�ӑ�s�'p�H��d7���P��D2~4�⡯��j_,�ȓz!�0i�.�v����&��}�nZ5f�ބ2�}���i�v�ä��{��逽���3"O0-�I�.���tI��M"��I�]��r5���0>��ˁ�Pl�f�n]�ᯈ|X� ���G!�y��<z⼹��݁|����lY�yb��>*U2�K	n����!�HO���`>�h��RP�4�H��f�[P��$h�"O����da��V���=z �iþ�B����������O�e�څRF��.@����/��yc��r�t��/�Pв�X��Z���Ę�����'l�S�m�1�zaÁfWE���
�lJn|2���O� �x��aO\�<1�桒�+x� �B"O�e�1�[+x�ļp���Bo�2�鉁m	2���i�"m�\d��K�|��	�!K�N'!�S)�ƴSQA�	�����M��&	ͨ�*c�"~n�m�������=V����PHL�C䉉{�d�d�B�"�ġi��=���Sֺ���'��w�D����3!a@�@eU�� AJ5�7O�S$��-��PSĴk&eAS"O\9�G�"QP���&AT�Z��ɢnŠ���U�z��<���,b� ��U
(�!�d7PK$E6mD�Q3�\�_����O?HWIZ�^�x蓅�)ց�pR�<��G��8�ޠ���B�&��H�z�<	�!��8��I�̲li^��3J�a�<�4��1]&-À/�J��jK�_�<�ƠY�L��)���**��M��ÞY�<��b�2��!�M�|�Pi�-J�<��M�]�Ē�g�D�\���nB!��P�C"}ȀH�$	>�K�*��0!�d�I&x@��M���2!	I�!��Q�q��I�d�A�}�ܭBWH��]!���&=�W�]�� �h6�
��!���

A(@O	t�hu�R6!�!�ā�oa�~�PLӾ^K�9�"O`1�u�Y:^��4����|J��r4"O]K3-��RAL�Q4�2 ��(Ӥ"O>�9�펊_��l�F"\.8���J�"O"U ��]�	S�#v !K���K�"O<́�b�&D�`�"�ٽg� ��"O��Տ��z��h�BκR|N�#�"Ox,���D;(���с�� |��"O��0�X�S����� ¼f���q"OzH�����*G���oהR�:=�u"O�I�wCP�l�a�D�B�湑�"O�%����v)��;e�_�����R"O(��g$+u!|�֬ԔK^�;�"OD��ÃǿI,Th��쑳cYl��q"O �@"�d��t���Y�X"�"OHX�#dQ�E����3d��Q�,�$"O�i�W��K̔DbvB[���L��"O$�HǍ E^�{�!�P�����"O\����rg�B!J���-�t"O�ء2��01���o��[��p�"O$<2a�J�L�p0�o�2n��(�D"O8 s�LG������B�>�;C"O���V��G(ܙ;wK�H�T0�"O�(�0l�Z�Dк%c��n�xV"O\,�t��,$����b҄q�J�f"Oʈ�%�8:���c�����taxd"O���0�ǀ7��T��CҏQd�c"O ���9S'̹:a(�jl>���"O��ܬ]vd���=
,�`"O�����O.4}�ɱǅs�|��"O(,;1C���%pD�/gHqV"O��@w�Y�p���$6_��ra"O�����M(a��M�N0��q"O �0�Ôr�[X��,EN��"O8)���PY�)8D�U�P* � e"ON��� t��L����5�"O���ԋ�E���j�'�6,�`"O����R{X�0a�{g����"O04��e�::�� K�O��n_���"O�L�1C�f�a�&��;9m y1%"O�]F��\�X�а$<�Z"O� ��:tGј[c$lq���&c�� ��"O�c�/
�}�9��@�.V�0�"O�4��ݘ|:I�@�N�B1 "O
�p�G� DvU�0OPs�����"Oڍ�E��M���A̛Z'�P�"Oa{fE�*U��l�e��[�Xr�"O"2uc��4�K�.	A(�H�'"O�YK����:�3Ռ*472�A"O��j���!
�1j��c��Axp"O��ϗ�@�|}����_��ĳ�"O��aCV�P��PV�N�Jq���"O�Y�ϐ{��$YA���Rd�ʃ"O���W=0�ѺR��L� rG"O@�`'�Ɂ����bW�-����"O�dCD�7��m�7A��??ޤ�e"OTUSCL��'5�m� �K�lc�"O^����=F��F�-NB���E"O��� 3��t	�ڇL �`�"O�[��=�mr��ME����D"O�9
#���\�"�a���8��e�q"OP�[�L����G-�I�����"O�Wh��3:p@W��n{ yaB"O�ps'eы+	 ���/بK���	�"O.l�� �7|�jq/I8T��"OT��rM�h��1�M�_GT���"O�pHT��.
���Ro]�@G0�k"O�3��N(5Fp���^*/8�dB�"OxT��L&1�L��b/�AXi��"O2��"nY�s��"$@�*?��k"OĠcAB��b�
����:Z���
"O�{gG[���������hy2"O�� ��8%�,; 9��IX"O���엖+f�H�f��i]��"OH�[7��*E0���<%(J�+#"O��I�+�0f��=x�e�*\�0�"Ot���n�.I��١^��!� "Op�(��-:l�u	����Ѣ"O�5(���J$D��R�Y���qF"O��c�Nтr�ڲ`S��"h[F"O�8��(�|�2�U;(b^��"OEƩ.G��Q3.�t6EJ�"O<Q�I�=>/R`J���tZ���"O �ߎ��x|������!��R'~K�\a�R$B��t�LW�!�D�	]lp��_&���t(�!�,}��sF�LJ��Ti�([�!�DŬ8�l�]�&=0�yV臡Z�!�U)�\�R!bF4O����F�dD!��Ɵ~ˆ}H���j>ld됧J�r8!�
=;�~趡��Dݻ���;i8!�$D��m��%wP^�;eD94!�DU9m'��K3��;v9�����a2!�DJ�no�bUaD�t5���DmZ�,!򄊎&l���#ïv'��r�&"&!����bi"�.j����"IP�!�dP BM�%��ɫr��mY2X��!�D'g���p�����*f�D�Z�!�A;z�@U� �%'�e�4(Q�Q�!��,^Al@jʖ~re�A�_���)� ��9�&fjt=[c	��)��H�'$���A�<(h����@'�x��'kT�բP�6��AS�:;�8��'��|�g��m���rGMH�J�!�'�
�����]D�H
���/�2	K��� �4�eDYB�z�.uF�P�"O��`���.�t�6��Hf0�"O�@�3!N JE8����.(*`ta�"Of,�%��W$��!�n�bf��"OB���Y��qaA�*] � "O��H���>���3O"@�X��D"O؈�ك=q�HAc["Q�z=�"O��t��2Ŏ,���e��D�"O`	�%�1'��K�G=OY~��"O�i�d�ل=�4���KL�$�R"O�庲(B�����O�0d$X�"Oj�y5��z�3�G3'^h��"OfYI���z��1�/ÝÚ�"O���JD+v�R�#��P*�:,��"O�U���� �}��튏!�,T2�"O��toF�a�L�a&-ЉQ.ΥQ�"O ���ЇF�X����E$=u���W"O��d&��<�:"tW�`��"O��������U!���v��!J�"O�	���Y*�=Ib�<K5^�"O
�R��Pф����|��l(#�|r�)�Ә9pR ��:K��i�%؋^�B�ɥg�^(!�HZ?̚r���B�75BԬ��#\!��V�)�C�I!�p��u�"/�2��@�fB�I)"$�+`���}��٬xH0B�I
&U����.M�ča�܃{�C��[9R�T$ �'�!�a�tn�C�ɹu�F%y�(�?-Ƅ	�`�U;TB䉯��\j@!ֱ�B���6~ B��m�� ��Ö;s�a���MYB�I�u%�%��k#o��D��;N�PB��07�|�C��d�����X.b2B�ɴ�� Ba� Rit)����:)A2C�I���ภ�
}Î	�*�C)&C�I�{$Rd���J�b�!a��fC�Ɍq��!LM�p^�Y� R�öC�	/��YWě{ܺ��Z��C�ɽ+��Hb'�
�F� e)Y/*��C�I4u���-ѳ���HE-�C�C�	��4�!��ʼe$PYjC�N��*U#��nTrD�L�HC�	Aո�� ɕ.�`��	(��C䉘	�:��b��:_""tɁlݭl�rC��8r��ъ�6u{NLc !ܱX94C�	 l�y�5_3d ��iX�R��C䉆�b��g��T��Ÿs�ոQ��C䉢E�"�+f+Z�Gev�k���C�6B䉸?|.QI⯅�4Ɯ��6�@��C䉘7\�+2 �N��8�1*2��C�	�f8� Q�Q���*T<�(�5D�8#P`���l�����!k.D�|�������;�BJ�j� Q�-D�ă�l�?�`��v�U
��S��)D�����[;2r�r���Z��ljPH(D�,z�\�<�@��^�J����t,D��a��8a�!zB��(+x�)ʱ�+D��x����88dd#D`4�9�P�'D��C��)�=Q��;%'͌�z���'�
���lV+�����	
F ��'�*�*_�6N�
$��'R(�� �'�j��!��zTN�R�<8�$"�'�\�O7D� $��(3:2k�'~2�	�L�K0L����K'/������� �H2G;.Kf�����I��y2"O�yg�ƃ@!]*p��1RIj�"O���Ӣ�t��8�d]�RM�0��"O45	v�=J�i� �>B5d��"O0]��B�K���R@o֮;&�]�"O�x�Iۡ2���S-�A��]X"O�ܩD��s^��cËH8f�:(��"Or�h�U/FL��S�/T�"��Q"O`HQ����O#�M
��Ӵ!���j"O���)O�1��P�5���P��"O
����"����0��=!ָ���"O����	1�@�IF4�RM�"O��e�i��h{�G�4���Q"OD��f�L��9(@���a	b"O��J�-�/�T)�Q�W0\����7"OX�wB�=Th�HAW���;�L��"O$���_	oWZ�QB#��x���q"O`�3�̕�@���d�
j�Be�2"O����e�/p�18�l(xx��)4"O\p��:��H�E�� vY�"OL����2:�X�PܲA���"Oƈ�4��4[y	��
5�Ԭ	g"O6�@�ì2���֏x��� s"O	r�ꚴ<���f[(n�E�D"Op���䕘C9�����1���Rr"OV岳�W������)'����"O:Ј�BB/Bt���C�jp�1""O֭{D�i�>��7CW�O�l� "O��j���;a����]�?\!��"O��j�Jh�go�h�c"OJɛ��T��������273�m��"O���^f��q u�B�t.ZM�"O�shT2r0�f=(Υ��"O� ��V���[�Vv��0�"OzIC[4�i���2�����"OVEsKή!�$���Q�KG�(�"O���8u���Z��J�j�&�!q"O*iS�A3b�Y�'�W�x"""O�0;��WmÜm3e���5�ɑ"O�(Ѷ�.P�pX���E(r���"O4};u摪\���"D��ά�as"Od ��o_p�Ό�0o��k�ԍ
3"OF���eȎ v��;��I!x)hX�"O�����` ����]`d��"O�p��m�LE�A�҄Ўr��%ɷ"Or�A#ۉ�
2W�T	 �|1��"O�8�܎�G8�=�Ս�Q���J�"O�܂�C��i:���*���`"O>�2��v��|��ɘI��q��"O.5�Eϊ�h	v�i�J��D-x�"OB�Sq�z��J%ǵ��0��"O�1�% �=zbM�@�@4d�F��"O��B��Z�B���F� �Hh``"OT}���W��]�UI����5"O,�����K����EŘ�;�LY
7"O��±'^�<�!&Z�(bH�"O&xvLŇj���Cv�]U��X��"OƁ������H�ش���X8�p�"OH��L5�� �K��A$"OXHUgT�;MZ��A���q�(`:U"O�!����4��U��цQ��i2"O��z�Z:4���D
��%��hrT"O��*C�c�l�zsɔ�;�&eb�"O����%6d�$A16ꕨ/��ݒ"O� �	���F���1���A{B�)�"O`d�k�b�&P�b���Nc�ܢF"O.;1��!/谣���,D�8f"O6���)<Զ!����5"�:��v"O�IX���sJT����hpށ9�"O����ݸe��)AbW�Y���"O|���a@7"������*C(�H$"O"��D�	M�D�����L�a"O� p���_������ (8��c"O��S��ʇ^��0@2oǪJŤq�a"O��K�D����p�gP�e�@��4"ON�+�G��j@ ����W*�ZTY�"O�HZPA�/#��)��A�9�$	"O��#��$��P%T�l�R�B"O��qD�����I�d��X�3"O؅�$ ąUK��J�ͦC��Ř�"O(`:�[�!�A���`�)�0"O�d��
2iܠ����#^�=p�"O,��Bi4�l�n� AB�"OjX�dԤ|���x��%��\;�"O^�:�.,Tb�s�1_L��"O.e�d��-#h�ʡ���4Y�#"O��TlĭSJ�| �e�K��d�"O�+ǂ�740��C�r�\�S�"O<���y\aS���hX�"On1�QaɡY*��7��3ȅ�"OPL�$��)�)�|�Z{`"OԄk�m6b>~mk!��"����"OnQh�+�P��#`�7(iPLk�"O�u��(�-��=�R���K�j�7"O\q���'�y�%UDI,}�'"O�C"1�!aU���E��"OF��._8/�]��B�H�dXp�"O*D��,T	����P�n�6�� "O&��a�^)w�\��+���"O U`�
{Lq�*ByF�"O�%Se&�u�1ɂ�T�Dր�"O�=ã��:%׮O�	8�8�F"O6ٙ���"A��11W,3��{�"OT��k��@0�kLPt2�s"O��Ҫ
�_��]��d̕2���pp"O0�����B��=�@:��tZ�"O��!�մ/�AKE@��6� <��"O��p� -DZ�HJC�ӱ�ѹ"O"��(�5
���<�4�hq"O\4�f����QA��S�K�N���"O�p�0�E�<hh����/8���"O
0���W��'ԻK�QW"OB�{�b@�ZM�S�ӌ,�`�3"O��&�@�B��m
fW(P���:�"O�4Z��S�J�F���K��`�"O����>jm���_�i#Tm�&"OZ�'���	���DS��Y�"O�uZ�$��<>$p� ŕ ;�.��C"O����׾B����D��d�:�˵"Od��C
](�N���R��r�"O��"�	�@�ȧ�ƿ!���)c"O��p$�Ƥd{�܉4����:aJ�"O|c���nZ�)��-�2�I�"O,��B ˑ��QC���!N�J���"OP�Cg�o 	�O�7�C"OʱA'N��wmD�Q��\Y�xL�S"O! ����* x�ݠ]��ѐN9D��!,�H�m�Q;ܵ�6D�� ��b2��!XH%���_7�:eB!"O�s���I�*<j�)����P"OBE��I@�����"'��Р1"Ot"��9Q�$��m��v8d���"OF�s��P.�$����Ȏ (�p1"ONM�
-2��0���$a!���p"O��;���!�`�[3�N`���7"O�,
$�,/C��G��'�vE��"O����AF�/��E�,�T�XLQ"OVlX%�<l2\�B��/r��$"O�JՏ.�|�Aa�Շ��i*F"O:�(��H,h�I�V)�>"p�"O�� ��s�BdZ�H;���"ON���M��|��=<��M�#"O��y��1xP�9�6��Y�|�u"OH�5��W*�H�E�U�Y���"Ot��C�(�+��Of*Бa"O
I�D�)����%�2����"O�{ �Þ&���R��0RQ$�?Y�!�d�9:�q����f�aw�S(�!�˩ ���)ŠT1~�$����p!�D�;��eET���(U���Q!��<3��j�Y�z�2�����8l@!�d�Qv����m�V�q���61!�\�>-I2�ƖzR
��.
��!�$ÉK�l�b��FQ�y�`�ͺ�!���78���KZ6K��y�.Z R�!�d�10���9��ߚt0�P@.A�9�!�dەjg
 �tBǴId����N�!��$O� pa�	�<=��BŒ�'|�@(�7Gc�<8��"O�4i HU�i���R`�B�L�^�s�"Od ��,��#���J�&S��)"O�D�Z�9rHsu�{�J�2"O>���@� �8 D� Q���"Ol����A��L2,^V�Р�S"O|Y+�^�!lEzīB!�$��B"O��8�.(���B�K^,j�X��"OH�c�,Ӗ����E��p'I(5"O�0K�j��'��AB��č^� h;�"O�Lig��W���B��.~�J�"O.�bFCǬV̔��N�$J��"O^���"�&Y���O�9<hYd"Ofq!�ǅ=�X}��GT.���""O�TC�O�J�R��c��",~��"O��3 ��: �2���.C�uY"O���� ~%�${�E:z��A�"O�p��K�(s L4�#̳0��H�"O�d�@I�8���1�3U�"���"ON�� CB)!�������X�p�Q "ON��h� x���K6-]��"O4�YtB�27�y+Ń�� ��"Ob�1��J�R$|�#M<%��}�E"O��@oI>n�д���Ԫ¬}��"O�@�t$� H	����7!�@"OZ}8ЎO���@�5��q��"O�m����8�`
�C�`����"O��T�T�!g*@DV�LѠ��"O�lI�)B2;&�L�s���v-H��0"O��kS�&H��}��@�IZȢ"O��ZUFE8�h���M"<��G"O>�����259� ��$�z�x"O�j�C�5� �h�O�E�n̲ "OZXڎT���x��S���	2"O�  ay��ݧ���5�E�\�ZUp�"O<SW�ݸ
��#����@H9r"O�P����]Ք�1Ck�"3�t��"O~d�u�ٗsĮ=C�&`����"O�AkWdO�3-��i������"ON���G�*Q��ň�u��("�"O.�S���0pS� ��^�bt�l�d"O������U�L�b�̉0Q,�c�"O�IIV�M���5
_�_H�K�"O,%���S֌�P^aȰK$ܙ�y��Tu��� ��H�
�S�#�y� �=�@Us+S���\����y�J�-o���h�!�$8��T���yB��x=$z�+^t���)ٕ�y��d�(�Ł�5ePR9�)���y��[�)S(�4FIL�pAQ	���y�ú#y\[c�U�T� ��@M�?�y2oJ�z FmB�6�0%�����yRF�h�b�b���0���;��
�yb��3<�X���'\���a��yR��֞@U�M�%tؑ��y�>C�>�S�L�p&8��m6�y#ҥ} ����з;F�Hc�L#�y�GǌULP �(:נ[')���y� �)h�+#�N�Af��yVN��y�g�Q�V��G@�>�"�j����y�
��=�����͇:�N�D�9�y���>m����`�8�J�&�y�	D7n�|�s,PScT�ї��3�y�j(,� ����-txi8$��y���"zجKR,�l��Qs6I���ybA�?���%��kN���  ���y���KR�3Ңu5P��ɒ&�y�5!l�p�/�?��x�2G�+�y�G4(i�FkhP�b�K��y��؈UD�Rk^�+@�1R C+�y2��9�67fS=~	�(j�yң�v>)���`[�5[1��+�y�c�����^ۦ|�☌�y��@�G!�cO��V�"m�`BD��yBI�
 j��K���'G� P���ܟ�y�2�0��&� :*fݲgÄ&�yr�D(+xI��H"+���:��Ҟ�y��T�k:�3OH���lb����y���.0(PzPeS�b�F��q�8�y�!P"WW�az�	�6f�
D+���y�N�7a�����H�V]IT�Ͼ�yr����h!�:��:�!�>�yRF��,B�m�D��L�ai1���yb�͇r��AP�C�8H������y"D�
%�& �t�B"{�&��DB޳�y�]�(@��z���p%0����yBj�d{>̲�b�
g��-��_��yҫ��d��@�Y�r����A��yR��#=�2Be�ͪ=q���\��y�DF���¼a�,y�a
��yR��"��U;N�XY��b1��y�DS�{��U�g�ڲR�ܙ
v��D��L2X(KÌ5��a���L�8v�ȓo�*�IUdѕֈ4b"�� X3䔄�U�p-
�\�ׂI(7�Q�)��~�⤓'�P�Z�(�;�#� r0�X�ȓ'���g��e����v>�L��+@�A��%:k2�_��T@l�<� ���1�)ņH�j�p�5@"O��J�T�Q� ai%*E?W�A�"O��[W�� m��4٭2VN|�b"O�bc�-~/PH�ūCjتB"O@�jE�R�G+HPp(�9���f"O�)��!��&w�զ׺U+���W"OX�УG�H���C��(fN���"OHY������	�q.8v*<�5"O&��eS\J�y��A���S�"O����N<0&�ŉ�*y�v�"O|xRK2����K�0Q`�z"O�\�&��΁!�O]�R�|�!"O.d����"\s�}�w�@�CA����"O� 1�NMt���p�L�_��$��"O8)��ף/x��0*ٷR��hr"OViJ�J��`���:�I�/�Z���"Oⵁ�m�Iu|�FD/cШ�"Or�3uOQg/茑�e�L⼺@"Oz90v�X�T�ʄ)2�U���1��"O��C��\6I�X���e��L�U"OD]h�	@8+~=*�K�Pڜ��"O���%�֥?��)�`�/-`� "OL��s�ڟJ�Uʛ�|�� �"O. �g��$�H�FĊ�(�PhR3"OJ4�愍m�� �dE�<R��&"OD%z�E1+hδQpc�?rD�d�T"O�b�ѓ��ԀpK

��"O�ثMU-Ƽ��
[�A<�T�%"O^�/'{ ���k�<*:��)�"OX`1H���0A�b��A��H#"O�$�D�I�0��Ô�`]2�"O��A^�s؀��D52Q�X�&"O����G?8U0�(�lѫ=N*e�"O��+�Œ"��t�Q�T(F@�˗"OF�I��,1�8�a��N�gݪ�"O��;�K�O�D��U�� ! ����"O�1��A�2>,0��8I�@YA"OȕcR_G�Ω�ƙ3��u��"O��K�Q�Xn��ö̆�WDH��"O��j섰@ᆊ�@`
|c�"O2I���؏p���aV��5d(�	W"O�5"�X\�0xH�ؗg��:T"O!u98=��3�
@�t{���A"O���l_�),�Y���
VK�a�"OZm���A��A��x= H�"O��%n���)2��Z�0"DDQ�"OJ\����.��1�iF (���4"O`P��F(8���]�xa+&"O�A����10��`~͊\��"O��9�$,� ��F��2m�@��"O^�S��J��`�R���U�"O<I���*f��t� ��4�x�B"O����7=���Vc�a:b)y!"O�,��ɇ�i?��GA�2܉�B"O���!��h�ԁ&B��s4Q��"Or6y�B���F.^��NŪ-!�]��Z�QOP٫�&U�{ !�H/2ق�3��Y�a4��SGFG�!��F�(d��r� ��2Yd�%?�!�P���Fk�(�Q��!�$��@��Q��闄M�n�����9�!�DJ1[��1����7D�j���GF <�!�� !8�|��Fl�FF�&\�!��`��� �N���	�Mu�!��  ����]� x'��v=��H�"O�)��$��zd3v���r��%"O�����N�?b�x�.�>�xE��"O`阃�Մyy���r��1�.xR"O`��G3'5(��L�{����"O�u�Wꞹ?\�h"d*_�Qʆ �"O�xX�N��>V��IG��T�U�a"O~�kp+R��r�M[B>r�4"O*�È�j����e#��n8J	�B"O(�S�/�I�ʶ�##:8��"O�x���'�R��
P�4
f�""O$�ӒF�!X9�@1��L�^�<��"O4�I�+H���y�a����`�d"O��۔�1O � � �"��@�"Oxh�&��_r�SW/öp<�X�"O2� pj$�4<��M��al��"�"O|1Y� ֙x~�$[%�jW|�sG"O�Ps�V�g<�(�i�#aK�
V"O\
%��,_@H�D�W>g�`X �"O^}����=A��p�g+i�pbF"O�H(�/�5�@�2d8c����"O�M+�*�>��i��ͥ:�%H�"O���&�9hz�|bb�4b�&D�w"O���LLn�(�`��u�$�Q�"O�d˂��U¦ *"o�$<�~��"O$@;��f����������G"O\i{%A��5��0M_<WPza�"O���ҢY�p���cY����OL�<q"�6e�j8	7�"!F�P��J�<�OT%m�b7�@'U�l�0/L�<�e*n2.%�b��%����L�I�<1��*D" �q�D	`&�@S�i�J�<�2 ,�K��L�~�{�l^C�<�MUc8%a"hK��Ġ�GOX�<��"�a�So�p�={`�V�<ɂ�^6۲�FÝ�"��`1�Mv�<���23��8���O���EX�<�&��t 1����4�
#��Q�<q��m*�%�S!i��#�D�v�<��BN;n DQ�f�J4<:Ako�<�@"�;O5pY�ȃ�i��x@Q�<A�΄45<��@�.��s@�i��Jx�<��I�~��������	�}�<�3OC�k��}��-��Z"�K�nSs�<�������;7��i��кI�r�<�é�*�PԨu��H��$J�TU�<����*�YR.Ɣ8n�i �N�<i��0LX��S���h�0G!H�<1ǋ�?V՚q�/Ն  N���o�C�<1� �.qr�����?!Z҄Cg��B�<���K�Fu��S�7G��8$MZ�<iVH�<;3���r��5 P���JS�<�7.�%O��Aˑ�O�X}�f�	N�<��#.���S�)^<5g2=y�k�I�<y���� �8H˲f�0!�V	cA�<�E�N&�l��H�-?d.4I��@�<��	��"Ҭ96oΣ/��8'�~�<Yᤆ6.��ys�B�XfXhp&�S�<�6gS�Aº�h$�B�nի���N�<QE	C�?������	9�d�#cGV�<���6?�̨KCOQ�t�MFR�<�֫T�0��E#W�d�5�i�<�d�)ltAz���f��$���n�<�a��#F��R��&J��C�i�<� �ʂ��M �� ��c��E)v"O4akQ\�I�He�����w*O�d:R�� �x� �4u�L��'�`JG��]r��P��=�y!�'�Xݲ�˕M��@���F#~�v��'n$�+[�o����r'L�|䪭��'�y��Ɓ*A�"�̀n|u�
�'o���"=,��Y%����Ҵ��e��4(��^=!<�laD@��l��ȓ̼e����;v���	g�0�ȓv��sr�O5P�j8�6o	k P`��?��=��AT�Xp��A�w�@�ȓ<JpPs��� P*�@�����A<Ω�ȓd��s!�a�âCUڨ���Dמ�1��Dϔ,���D��P�ȓqW�P�?6���TH��.Q��n-�U��V�It�r`G�8]���j�����,�U�@� N!�s"O�H��[�1^��öeݵp�T-H�"O�4�l��&n8��e�,PҊ��"O��9���3'ر����,�'"OR偛a�إk�"W�qu2e`�"OJ�8e�T7�(��� N 	��+0"O
x1���3i��[�o�%2⮸ZR"Opx��/pv ���m�
@�Đ�"O��K�f�k�p{q�\�nL��"Ov��Z�J�K�+t�d]{"O��1�A�s��srk��F��A��"O���. ����:��	*!�Z�1`"O"�sq��!��¤
4Va(�"O��t��<3~F:���
{�jᚵ"Op`0�D0\�x0�Q�V5�m+1"O��� �N? dB��N�L&>�;�"O��o1T��sB7;x�M2"O�d�V��#�)Ò�5+ÎX"OD�"!�!�|��C����ٴ"O~Y S�_3F�ȑB^D��}y3"O�y��X�V���ۀ;�R���"O��H��C�9��R�Yw�P%1�"O"�{���+ ��Ѐ�U�/��"OZmC���!ف)O)�&}�"O�	Kt
E�$th��T�y�hL�4"O�\����G���PT�̱T�htS�"Olչ�;"�f໱C̎b�I�e"O���ʀ�N���C� S5[4B*�"O`-Q�f�\ؐ} %O[�2�"O�d��)CdQ8�*�c 5K�3�"O�u��]$#	z�����N�.8!"O�H�3n��9��ţflI6i ��3�"O�m���8C���B$k�\���"Odp�R�Ɯ*猑h��W%}�U��"O@�#s��/Q�ͱ�O `M��"O��f Pp��k̂-NA�9ca"O@��,�~V�زQ,�����"O6��s�I�,#��"f��Ȼ�"O�M�M�&z{������9T���P"O�D��o2(H9�ʟ�q�zG"O����*�D��O��QE"O"���㌄Tr�M���B�X׀6"O�`���2-�� ��j�&g�"}P1"O ��b�V=8x40� ��lr���%"O�<�P��f�*��O4<�2�C�"O����A�5Y���kU���=�*���"ORԪ��;����.i�*�"O�  ���Z�\y����jB�,���A�"O��J��.DL4:t#P"mvU; "O��� *ºM5رA���!"O�M�t��<���"�\�a"OB��gM�U9��I��{;�DA"c"O*��$	@4P�:sHJ& ��|��"Ol����N�`PH�XE�@N��I0"O�4��\�H5���=3���0"O���n�3'��yu(&�"O�t�I	�B�C�iT=��u"O(��#`�8~�I�w�[�hH` �u"OV���� s�$��p��H(`"O��x�Q���1R:���"O�$R��$]F9뇣��6x��"O�a�˃�
�Je����pE3F"Ob�qd��X�-�V�U���	#"O��k�(�#NV���A�*u�""OR��gW�O��9 *F�c�p[s"Oͺ��_�.H��J����`%��y*O�"%�N���JV�I��`�	�'�̴z�ږ
�v�+��]�w:�H��'�:Lx���+ �Н��b�0D�PK�'��!��:12�uQ1Č�9�h�Q�'��	�kq���p'��,�����'-�x��BN�z�.�[Sc#�\��'m@���H�[m��ɦ!gH`��'��N1
)��R�H/(!p�P	�'F�q84��s����!d7+^d��ȓ<���Bǉ)]��y�Ƿx�J��"D��x�ƅ
���!J�9���,D����&��q�Q�݊)TTr))D�`"v&�>q��ER�"@�,z��2��1D�p��/�M�xE�F�%ZT5�5E/D���"�~o�pc�{��M3�N/D�P�c�ߋ1��㇈�8n�ȡ[�!D�r� ��5�Eg2u�z�f$D�|Ȗ�[Pl��R`ғr���`B?D�t���&5�tUiu��D���'�=D���1�>�sv(�W���XE#;D�A�$&t���s ��8��c�4D���T!�0g�d� 2'ό�P\J�o-D�$��`��
��C�m�~W�3k6D�l�q�Y�2�"xkW�Ӡ+BbHf�4D����CW����\�4�J�ɲ�1D�d�Go@�p#8EY#�;Wj�j��1D�@��6Mr�(H4m	���y�P�"D�t��[�+��U��f+4]pa���<D���TCI�pc ҧ�B�!��<D�pQ�E\#`�;��ёl�؁0)=D�hP�OT�	����R�4��ѐ�D(D�p���O�@D �@i�3y�|�Y��*D�`��J*2����$���\�L���'D���P��(Htը O�.�2�H �1D����%7 Ac�� yYS�*D�d`�:-�c�e�z����`)D�T���ޮ/���[��Z�I��*��4D��SdJ�b Bl�b!רX�x͋�/D�t��"D�xKh=����C��u@8D���u�D"u0'L@�@�t`y'5D�D+��_c�c�AZ.'�@��Ǥ1T���!��4<L��R�I�eX�0"O\�K�
�6*��2�P�M�Xp�"O���۬sh�V�R2}���+D�L��uH��2�
a��QD�<D�� ,��L��[mx�,��:\6�x�"O��V�ׅ��0�ˏ?-9`@Q�"OR��P�M�6��(@�CRf�۴"O�	�%� i��3QOR� �[�"O ��qEĄN���@ծ�.���RV"O�u�
&�ܝ��-���AZV"O����
8J�PK��ߙp�,���"O���ӧ1#�``���Z�~����"OLUA��R��6p��P�g���5"O´�cD��}��<A�l�3Q�j�"O����J8c��pCta�&�Ԛ�"OҩGC>C�z`AYu8�B"O���+1W�Prq�F�c�"O��Ak�'�\�d�$TL�C�"ORB
����S�I_�;0 �V"O����'�o*d���T�B}@���"O&����J@��TÝs�j�i "OܤIg���yYxp��D�,�D��5"OΥ�d�υКd�wI�:�Ή˃"O\@���(tot�P`�?H��B"O�Q��@0Be��Yu��90�L+"O�l�"�øXv8iCG�r�z"OF��DD�^�b�Q�Ȯ#�a�q"OrU�B�4�@���o���� "Ot<�7+I���%��7u��h"O2��0㎙z�Z5AU&Z�v˺�h�"OԀ`u��_�Rg%2h��8��"O�(�d��#�2���T4zeZd"O6�k#�G�{݀Q���L� Lа"OXH�/�GIu"G�W#g,uK2"O���Q�;=H,S��IU)�l@�"O2��$YJ�Y�nĔd���"O`8s���9�a2gߜf_b9J�"O
�sF�^�?���;aE[��&	�"O ��E!u�-[�"T+e�\h�"O�y���1vB �G���t�j�{�"O��� L��a�J�İ?�FU""O.UB�P&|^*Q���%1����t"O�q��5L�UC�Z�gI6�2"OD�Q�D�!)��=ɥ�3w/�0�T"Oe7�QN�p;���?Zp�"Op(iL�6}K3�Ο� �"O0�q�G��\�t�+��E�f�Z1"O�����+fج2 �<�L���"O���2�ŽỲ�g�� n�`l��"OzĢ�n�y}:}挏|r^}P�"O&MC6dX)k���"�E�#D �(:�"O$e+Fl�7���&�n��W��yR��$����#�@�d��f�O�y��=5pxVK�L�6�)�����yBd����<U�ߓZ�b���]��yb տT.x�j���N���$(N��y�o���H�)�D�}�$���'E��y�i��=C�<F^f�E�����y2JŐ{\���B]: &J� �?�ym@�M�.I2EȚR���o�?�y�"�2*a)%�5�@��I���yB�"a����eʗ3�) 4'I��y2�]�x�H��2B��}�PG��y�h׿<�4���L�iQF4�7c߾�y�d�,esp1+�7Q�}[�o�6�y�5��Q`��7D��&���y� Y	b�T�٥��4�`́�+ ��y"C�jW x3ׄL�*�H��<�y
� v�#E`�/R�"�w���6�, D"O lp���e�1��L3� �)"O����
��a
#�`I�"OB!�7$χWJB�X1OHi���"O��`�$��v�<�j��X��P�"O(1�P���,;���`a���
�R�"O�`kG���f�H"�"h��ɩB"O��҄H�j�\���+ܣ�Xd�S"O�i2�.K^�� 	�*E�Tih���"O@U�U��R�����H�</U��"O�}
G���k�zaG�G�a�"O:u�EI�e��dߡ>��p"O�m���$9ݙ��Ř=�x��"O���e'9\���;�E@�b�����"O�5ړ��%,�HP�@�<����"O��4sHݩPƋ�4�1"O���@)L� �Eٲg� P�A�p"Od%�3A�55t	z�L��H�v�B�"O4�6�5��t�Ǎ1:8�)�"O�5�@-��4����FK�ZR(б"Of)�FHT7'�.Ezd��;4|�5"O��#�	)p$s3FR�Y�Z��"O����(Ӹ9��
��I�لb�!�L�>����m��JN���j@*�!��]�3��yS�f�44�H��
��-�!��ޒcg̥�U@�/3"���j5w�!��.h>��3�X�%�Läǁ;T�!�$�d!��`��9$>�P�Ʊj�!�$S��1A��W��L�q�ɢ%�!�dO�o�h��	Y�4ga�&܍B�!���w�,�"pL0��A��<8�!��Q�	:�����"|���s��!�ρL
�H)����F�DJ��[�!���"��3�$�>Xh���)�!��+�,ZQH
;N��VM��!�_�~$��C�-���'*�!�䛢F�x�)��!r���l��HB䉐��lp�ˁ`@18���8?:B�I-2�zUa�ȥHq=���
�zC��/i�`�儙8$m�1I	�9�BC�I-ޒJC(T�[�I+�ğr�B�	3 �8��r��=K��8 bgf�B�	$ZxB�����q�����l̸t C�ɭZ �%(�d�=/u412EE��!�JB�ɤ��1Jef�]�$��%z?LB�I4P��+EƉ�D�UY�_�E�BB䉚 H�S�'̘
�����N\;~�B�IM� �QW
ԉW�zɃ,>4B䉄):n-�f*�'�H�vI��v�RC�I#x�.�G)X�6��aEv3�B�I(1�jԃ���#�Ɯ�-ɩJHC䉣<�4�;䡄)qZtD�$�/?��B�	<7�@��T�ǿK=$�qa�fsJ���+�X� O��/��sW��S�A�ȓUf���G/s_G�	z����i��L:1��)[.�ă��Z+j����ȓg�d`Q �U�K�.ŐeP�=Ѐ�ȓm����T�b�,=)��$�F(�ȓ&���1�A=%n���s�A���*D�$�Ş�]Ϻ�1'D�!Z�+�g4D��%Z��zqY�I3(<0�N1D�Dkd&�6��;�(S�@�:��/D�X�w�R��Ɖ�2%�$b��+D��&KB�D��5�$����0���
=D�� p��ӭT4ra&4;�*\�A�N"O��
'� s�R`��#��u��"O�pZ�C����iW� s�J\Z�"O~����K4G��4J�b��
����"O��(@M݇1��$ca�Qo�mC�"O���B�'�艠�NӬP0�5�#"Or!X����&P�[w��"O^X�c�6+˴�Y��S^^Ih'"O����Λ�XBԁ�"Ϟ49Lp�R"O0��'��`u���$I�	:"O��{v��'j��P	࣍�L/M�s"O6���R�A��тޞF� x�"O
�'
^���Ѵ��՚�`"O��5*ߨT��4�rԓ5���q7"Ov,
���'ܘ�D��,�����"O�ҡEϙ)L8�K֚z�r�6"O`�!o(~���'&�|H3�"O�����B�AJl<Sc�/��q�"O��)q�ߕc���;�섅��pV"O��ApaIvwZ����Pe��,��"O�I6ϖK�2c�ԭj���`E"O\�1�<6�����
�����"OD���D- (�,�"�T�"O�i8�+�Y��u2�A�{����"O6����N8U�^�	E��^!U"O	s��)肴!�,��[�����"O��h�O��wh>Z�EQ*\�)t"O�,�`g$U��A��y��"OΡ9UZ�a�!"D��HLp(*�"OB��q�۬37�4Xd�Y�u�ӱ"O4�!��?N]Ѭ̤7�r���"O���B�6n��Y�,�%W�*�[�"O��6-á��y{gP�|�p:�"O�J�U�v�%���X
	o�Q"O��3�WX��h	��Z\�HQg"Oh5�R���q	 %�gS7o4@Ap"O���"E��@D�H�N�b	�x�"O�u��aB�EޚMӴdT�M
.8��"O����R������2x���T"Ot�cڄzT��GM�(�v�4"O$$�3h�\�&h#b����	�$"O��p&mE t'�D�di�^�Vq��"O�!r��j��4HY.M֜#�"Ov�����ER"Up!B+��3�"O��M�,t@ȱ����a�c?D�x��d�z��oB�a5X��>D�D�P�߆Ry�i��:u��`�<D�8�dA��"�c�3E��i$�:D�� $S�K�\�O� ���ᶥ2D��5�
67X�
&b��	C�*D�x�T�#R&�MRu��-Or�B��)D�@1 a��������Sm�`�$D��#h��T�4���D�1��˰�#D���B-42(@h�� %��@36�#D�L����+���@#�� -J�!4b5D�����V�L����$� bb��G2D�<�e���HTH�	W8Q�B0��3D����,S��T��F�� J�yP�6D�X �j�le�`c�L$�F�p#6D��p��$k6Z�;g/�'I�`��f3D���!�ID�U����t�W
0D�� �.M�qqv�As0�v:D�����N� К��cҕ5�*�
�/7D� �����Ar0ą*&L�(6D�� �i���Y�J�rU�ƍk@���"O�=u��>"e�O�
��`�"O�q��n�����O�Z�<��c"O�8�b��#,�p�+�M�?D�)��"O&X�#�%
nLP@Í��:��r�"O��d
#(�4}z�ʼP��}*�"Ol)�S	 ��[��OKŚC"OV�w������� a����@"OL�����O�d]ا�j��,�T"OBpPa͏�8���*�HvP��"O�* ���L�n �0郍]xIg"Oɢ@y��i  h�;#^a�1"O��c��A]ϖ�J��
	\�EY�"O.h��	h��	��4��<�s"O6�ag*ěuQ���	/2���5"O���6B�J�ˁ�O�h�Jp�W"OJj�F-Ҡ5��ú@0�0�"OD�[���vG�����=s�"O2$�ď7(�>1��c�:Q/��p"O�&�	��α@u�6TsV�x�"O ���@	�4���];4p"$��"O���C�/��\�6NM� QZ��""O�����һ{j4$X\ʨ�"Qn/�y��-��%s��B�^k�0q�� ��y��)I�����-T¸�@�Œ;�y�iO�1.�+'hL� �ڱ����yr鋥r@�٧�ń|!&��&�ˋ�y��Ջ|(T�b�	��D�0��m��yr��BZl-kS�
7��D	���y�M�#W6��Y��Z�8��ٔg�'�y2-W=l�xh2- >-240#	���y! �2�8��t.B�:R��`� <�yb��89�.���4g�dx�'���y���n4��Ѐ�ɹ+�ֈ���	�y�m�'1o�����*�=Qf�W�y��������AB���HƆ��yr`�T�TYh�MS�$�DM<�yRN��%�W�@�R� �5,P��y� @�jA�K6E1�����	��y�K�]�ᐡh]!@�4�	�e��y��B�a�F��a��6�z�3R��(�yBJ�a�.��4�Rk1f���yb�H��䰻U�S0^�Q�a»�y� \�{�����敢N3�f�ܵ��'�t�_q�Y��ҬR�\�k0�!D�`�鋮`Z�B��ԉ;�@#� !D�T��D�`F��+ ��/A��DZ4�1D��h�����nXbt��"�+a�$D���
A�(��ܳ�B����9s�#D��`���J]�)�$>��U9�A?D�xe(�TzθcAΤDh�9t*D��qQ+z1*�p�iW�sy�����$D�4 �
ߚH�TI��d�+�M#"%D���4�+o��jb%�,�f�iT�#D� �`�=`I����_�#0����.D��� D�j���hޠĬ���o-D�0�dU��<AW�F5ug�-�2k0D�����A`�ࡁ*�$\�B1��.D��q%l�k����"_ pD�kf+D�������$۰��W %Q���pb�;D���֧Ʊ*�J,���$6aP����7D�0+Ƥ%\W�)�H[�\�`a'�5D�b�I-8�d-�`!�*!~L9�5D����#(���Q
}x����3D�� L��L�s@Ȁ�!��B�\B4"O��#�I2���E�t	W"ON�0n�����d�&>P�P"O�q�S�^���ـ3��6 ܨb�"O�y��hA�P��	���M\`$��"O�q�2+D�.|���"O:Q�B�)��@��e�i�24��"O:�����P�V��&�%$��y�"O��1(M�rQ��t�#7&Q��"O\bg��f�����5�ذ�"O5���І-θ,��� �l�2�"OL�1�Ö�o�zi�7-����E҆"O:-˒��R�Di�bW�]]�|HE"O �ԁ@<b���;P+��tSpxS�"O�4%�S�V]Xث�)#"���CP"O$�2V��L��m %	�L��J�"O���ư%�]�2��5(�֨ �"OԵ��gl��"��B�|��M�!"O�}���6!n��[�e�3I0���s"OJ�h4�
�3|z	3��o.$h��"OrH��
B ��@�6 ����"O��8f�MxL sÀ�w|�6"O�� Į��
�`ďĳc��1F"O
�rd�G�S&`-ɤ�� J�Q"O���pe�TT,ԿnZ*5 �"O�TʗG�����Y]�4��b"O\Dj�ߣN���˞�z���x�"O���%-�9P#t`�dLb���&"O&q2����P�R��1%vL+�"O�1ʗM�<V,81Q����h��"OxD�B�� %��M�����"O 8#��-v9�2A�R"r�|�t"O�ja���,���ւUH��2"O�y{w�K���+��X��"O��kPJV�a�0Qƪ�	X�j97"O.h´f�!o�S`�ͼ!)�e"O�h�ݵ"�&p���Kn(S"OB@uE�� J��:3�¨r}��"O��+�=z��H� Y�ob�0�"O��I��K�v��A�!!�p��"O����
�@|v!h���d���k�"O��@�G�g�)k�;֖�	"O�����׀��p�4�_
Q��	��"O<���@sg��g#¡O��9F"O.�P�CA�#*^t
�!�g0�+1"Oeٓ7W �@��W����"Oyq&h��?��QP�� D���!w"O�H#� ϴ�(����|?�0��"O>��4���\�b�kS�0���r�"O��Ð�k֘��)o�H�m��y2,���B�0E��L��Ӡ߯�y��V:�P�%�@�}�"i �y"@ �Q�8�b �bo4H�5�@$�y2���z��)!d�
hd}�3�U��yr�?pz�^2,�rC���y�8A��HS��՘]a�\�#T��y�j�nЂha��ƥT�O�tWl�ȓ6|�`aG�I�����hܤ���c��RQ�׮.�9���F�2�t=�ȓ_T���S�$aC�Js�^a�ȓHb�f�
�vO:�P��ҍb�d݆ȓi��P�jj���J�4>h-�ȓUW4�s�#Ȋt�����M}7�8��6
#�ڶ	��t:!��@ ��S�? LQ8��H�#��A
2I!q\�c!"OBlct!�q�|a��.����%�"O��&J�7.X%
2�;>K0X0Q"Oz	Q�GU�p*l�1uf�7�v���"O���&$V�T�8U@P�J7bqP�"O�u��� QJ�Y�GͻjIzD:�"O��s���Nf^��F��t��%"O �FI�:�����ѳN����"O�$Y4HŦ;���ˣ��d��R&"O\K�O�89���耋A�j�LŹ�"O�-ش
\��	(��67L��"O�h��#ʜb����v�0TI�A�"On=Ia�))�|��A}=Z��"O$���I6�L @�q��@g"Oܤ�V�:@n�ԺGn��*����"O������D�CmلI��!g"OT���E�%-���[M� L�Ĵ(�"Ob��� �d��M�<�����"O&�#���4納a%��'R�`r"O�p��$+6Aps!Պv:]�Q"OZP����ܢ��v ����"O���DOQ�t�n;7 ��*��"O���"BLm(�$�2<�\q�"O��֐Q�N�aIڊO�H�"O��bvNE�R��E�ć��-�L���"Od�(��,i0f탂�U����R0"Opt󀭆�yZ��B'�����"O䜲���9)����P�D�b���"O��s.N�`U��ĉ�4yy+�"O��R��yf�L�GN	-<�8��"O[��!̅u�6�W�}�,�g"Ozl�A%y}64+@�S�L��D"O�ctf��}�%�VnI��<u��"O A2�L6=[��o��D߄��"O<d�%"5n
h�*ģ�72��E"O���� ��mر�_�`0^4� "O�h�"� Ah6��e'ӝ["��bc"O�	��k̸jJ(@��D�F0R"ON�x%*�0km,e2�T!E�&P+"O�˴��O�(��B?|�X�P�"O�X�-�!Q� ���<��r"O�<� HS=�t�@gEh/ج�"OP٫�G[U ��T��=��9�"O����N)
д\����7eG����"O���P-T�&��a�\?5b,�w"O>|�t�P�Gmf���GZ:G�3�"O� C�a��%ـ��Ȃ� ���7"O�	x$F�(</B�!��6?��})�"Oj$�£��B*�fpP�c�	5;�!�DS�z��M����ayRL �h�#[�!�'!B�B#.S9q��¡�E�&^!�d�(M��Ek�j-'͐�;�وQ�!�D��K=ĵ0����Xdo�>�!�dF1R̮heBV�a�Z% W�!}!�$ m2q�!��|H؍K�#T@r!�$P�,xT0��,��,LP��fCC�[�!�Y�D�P���&B5����0�!�D�	l��!��R�5��Ȱ�
$�!�D^�k�B�#Y�$R'j*H�!�dH\�ڼJ�	�D�=*	��"(!�N%z�L��"L7�|M˅(ҥ!�B�<{w�ԑK��)��a!�dšK}ZL�E���>��-÷�V�kf!���;]�\�f+U�?�|Z��qP!�� ��%WG��U�گk�&�i�"O2�B�G��i�lꒋ�<��P
�"O0�6jZ�3��仠OA<����"O�i�6ƊbP��ƭ��� Cv"ODm��˙�s:����,�+� �@�"O�@��Ff���s��.q����"O�
�����;T�#|�B�Ap�<A"*֜pb�pCW�H��`Q;0ɛi�<9��	/pP���@�X�u��y2�g�[�<ek�CT.��g_37��hQ�SV�<�U��2�Zp�UxT�QB�H�<1�d�7X�N\�C�(Dh�Hxa	�B�<�7��/Eb���O��
o"�� iI�<��Ɛn���y��\�U��e��#P�<�𠗳D�������jAb$��J�<��D�;8��
��եj]PG�q�<yP�@�,��pⱅ�r�z���END�<��Hؼ'y�`��+ѿ3~�(D��@�<���W�|q��ip���7T1�%{�<�$������I�P�X��t�<�aU�>@�5�Re̾"fV�H'��Z�<!f+	)p\hp��J^duh�S�<�t/6�P�T�YUmMht��e�<)7�K�o��B5f
S�Ԡp0�i�<�nH�(j~�����  �@PR��J�<���W,T��I<��ѓ���I�<9��Z&z �������|#�O�}�<YËI' 2���TN�[��۷��x�<� �ȧ)���")CJ��ѦMr�<v��k�$�Mrd	�$C�f�ȓ&к�X�*ǹnY�<���V$h
0��ȓ_&rmy�JO�~n��Z��TE�ȓX�6�сMF�f]�A*�@���V���YP`��?�`u��Ǘ��p��xM��l:$��U�%�@9��E�R�Z��v=�"��~�<��>,(�2'O**cy�T�f �ȓD��!�3~.P�v�F��dU�ȓlO�r3)G�q2ꡨ�-��z|���6�ۇ�؎mj���6iѝ:=���v�Q[�H�@�Xq� ˳7P5�ȓs$�P���@��dz'
*mh��ȓ/�2	[���#fu��l��<��ȓ}��d	[T(���͌b������Z�q�Z5� ��-�>�T�ȓnfj��b��Oٸ�[�������ȓ0\5)�
���� l�60V4�� h��A̚�@�<0�/A�D��؇�a�8���
}s
���W�%���ȓi�B����+V���m�!Y
���M�P�tE�+S��\B#�Ĳ
К���2l*�oN��RQ��,cZT�����<.To�pu��O�%G�����:����Co����P�U���#�PX��r��r�	�\�,�LX�v����ȓ\LX�i��ڢ\�.�z��
�hl�ȓ�:���q�Be���݅e����4/D���&�� �&o�>D��ȓV#�h�FLz�LU�n��yN蔇ȓA�����V�W�u$Ň�b|R�@�i�#k�b$C���	9�
��*�8����v�fA"#͊K��ȓ��Ȍ>N>��Si׿^����ȓXۨE�Q/'DnK^�&|:d�'D�� !�`�%X��0��s��Д"OJ=���ɖ|�����B���Mz`"O�| �%ͨ�NX[����pyX��3"O�˶	�����ɕ�G.$�B"O���#C�ӄX�U������ "O�MS�`�X%�Y��U�I���a"O���#B�t�h!����Qچ ��"O�XC�$W����Bg�	x�F���"O ҕ��,���6�W�T�����"O��C&�K��$��Q�-�(YJ�"O��x�o^��c�E(%`���"O$�(�S: 9jq��nQ�~W}�4"OB�w�N�SC�p1ůA;2P:� "O�`���k0h�vN�;n.`��"OddrebJ��(� KLR��p"OeX�$�9Ŷ�{d1@�1�"O��2����Nd6u��'̇ƺ�{�"OFDq!�:Rs"U��g��L����"O������"�䙭I��1�g"O
��j�orb�#�dO�K�tT��"OJD�6w*d	B�Ú4.�R%)�"O�7��72�̌�%⍕;x��0"O"��B�ՁzT����4Mc�zu"O�MA��_�T�C�Ըe�p�"O�y7NA�Lj�I�o� �YD"Oɳg���-���4�4��A�s"O��g�P�ol��3bZ�#��� "O�q�l	6l.A��X�es��0"OĘ���P	�ٱ�"��P�G"O8 �M��@ǺY:�I8y���)�"O�Ԡ��R62�A�`��|?,IѢ"O�	�Lݲ|�Jɑ ���]H5r�"O(E(Ƣʈ|�6�:2a�1nF��"O�H
aiү@�!�o0���!�"OdYYE�y	�= �űq��`"O\�3���d��Y�67�"O��)2⊍#�P��$�H1pހ��"Oz=I�(��k?��K"�O�R����"O��Ydo��L,�� ��%L��	:"O�����ĺ8��=)���I�T՚�"O�uj��2| (����!{uF�"O���Ḵ��"�͓1�hAP�"O��02)S
<�X�S��B���"O��aU���H	�P�P��(��(��"O�<Jt�Ji�t\�cBHcz����"O>9r���_"
����,��sd"OLaP�DJof\�z`a�RF�Ɂs"O (�S&ĭHJ�
��6W��J&"ObH0o�7fI2�P�NX=�"�9�"O�uB&�Z>TSx�)��e^���"OR�R`i&���$_D��xS�"OLMc��*kr�ģ�t���P�"O� 0��2S=��+ �I$.6�-q�"O����험XӞ���NB�65n�p�"O�£ W%"2�x!��?P��"O\̨�mC�@���XQ�F�W����"O(�˳$)�P٦�lu���"O�!����(Y�*�.mR@XBw"O%��/J��1�`̎�k3���e"Oa`�&��+P�U80��"O�9��M%!i����G�U)~�	F"O�d�V/,\��2���+��"O�TC�5�~a4 �+BB�`�"O�� b�bS|��D�_)k2��s"O� ���2K(. �5�i�(k(��4"O�)4�D1>Ƞ��ĜǸ��"OH�që܃���*��,I�>x�"OZ��ƥ�8�B����(:�t�+�"O^(J��F0k.�5Y�Mys���@*Onh�$.�@�!h��-0�\��'��p�	3P�l�E�W/S?��)�'1�|x#.;F�ݐ�i�%9����'T\�'�� rG�$�`J!I�l��
�'\���B���(�2�f��jRQa
�'�h�h�f�,�}6hF��:�a	�'�Du
QI����S5p��'}�<ɶe�#L0�IƉ�$5j�AB��u�<��K�X�9 "��������r�'R�M���J$Z�Ib�x��A9�'���q`�ǲ`����	>z�X$p�'"j���A�jEy�K?p?|�h�'��e�F��))�D8� �w�(5��'K@���e��J��0�GD�:�����'�LL�S#צ@
�$#A`�??�h��'0��B�7g|8kq�H�`N\�	�'��kUeϟo4�$� �E_$}��'cf�9�E_�h
�gτL��=��'R4���/=��墡�KT���',x�G�ݞ9�,�-�~b6���'r�Ԫ<0|�ͪ��W8��i��'�(�8�a	 &�zTÓ���>6�B�'�&�X�M�W����e������'����%_[��ٷ�ڋ�4�{�'W���TdR�ǦS���r
�'���Ä�4���_�bO��R	�'���Wr�5��d�8QK�'�4��w��.�]�D��R����'�$a	VA��L�!��8��,Q�'�ĨRc�*���#N�M��I�'��q2"���XR�;H^���'��0e���H�}A��w��t8�'�$pàBM�H�LA��� i�$K�'�(
�oP& �����/W�U�&(��K�a�a
�[�0���gK+K��방��O{┆�IW�>���-�����j)1-4�bՊq*\#�!��[!E�V٢%��p�t��	��B��,���se���uG���]j� �2��dߤɐ3���ykp%�C߳e� I9��*�5B4b���O�b�U d�1�1O�� ��׳�2HѠ�_6�4H�4�'2����۝2�,��5��6!HN���O�{>��aS�C[�`
�[�&��$�ρK��q�mV�Q�D"B�5<:�:w��]�tH��O��Sh��W����6X(X���'`�|���WT�h��=T3�����j.x=P���r��+��*lf�tF�D�F,t<��+�EK$��FK�!��΋��p�C�]�$����B�8������&;ܵjb�X�8"R��cX?�Ey�hF'x�' �*:�D `�ۉ�p>�#���m!�)�a�Qx�y �+�,h�� ��
.̂5yu�݄%�l���'�����͊#f�t��/]� ���K��d_~o.��G
IN�đ0e�8X�y��O�ۅ��� c��Z2B,��X(	�'��z�ј*��1��]���@*�*4h��1^�$��Uή��F�$0�� $ӽhn��h�"N�W�l�xS*Oи�DGV0)2���)P��@i̩Hqfӂ�ޮ{|�
�����t�q�'`P��f �I5�D�s`F�t�	�:j8xa��mJ��f��p1�5(�̧�(��� E��r|rǣQ��t��I��x�"P/K4�Ep�kU�F� b��B�hQ��|(�ej�>{o2�pǡ-V����6"\E1G�� "�|��pk�h-�ȓ�4� �6m:°Cs�XZr�|(�H��z�T�V�͸3h�9Ʌ��0c?�I�1�q�E˗�p�Ӓl�1"��F"OJ�@�ʆ{:�9��P�����&	U�F�\��di3�,[�k�J�ʄ�(O� L�Y��6!\YB�
 TL�R�'��`��(����(J�̰<<��An�9L�|��Θ��rѱc!�4���*�O�(bw��<vU�mC�0���w��W�{���ԥ�8l����ӓhl��7����-�&ѠdK����fL�9��Uo�<@'��~��LRT$ǯ���aP��}���)�CNd��p�	�]d9p ��B�Ƴ6m��.��qz�'�|!!�D���!t�I�儠S�,OX�ұJ�G��0����(5l��b�Į���y��d֑z�r��X�Aô1H�E�&8��z� ��nFIIiO3\M��S��J8Ǹ|�OԱnQ��q�����ȸL˶�a}2���z��mq�iC!e\��j�0Ӹ'C|3�h�+��K$�
L1�r$G0��ʲ'�5�fbY)A������
�!�$�'��	��Nj||�cA�N��`
K[{�͑�G9@��qP�S��y�o�)��  6�h)�f�A�_
|�ȓ}�: P���8cܚ���l
%D���爃�4�B��m��*��@b�
�?�>YС�,B�!�Ą7B>�q�fFAe��a�41"=��KP���Q��E;t�x��C�^B䉢ewd�rӉ@���(_=0��<	c. �du`�z��ө7�F`y"K��i���!_�o��C�ɷ]�ªmcX�Ct�C'b�t����<�f^���JL�IZt���.�s���`n��ϛMu���ȓ^��)Zf����0����)����ȓmQ�rȎ$I�x�N],p>���f�R܃Ņ�,%���M
�*s(��ȓJ�+1�<���t�#Ы'D�dj��L&֥�$(�,}bX�y5(7D�`s�D�A���db�����'7D���C�W<rJ
�a��$p2��V#2D�L��Ȃ[w[&��~
�țg�'D�$�`�Y�f�АT�~0"����#D���S.�"�x5��F�kM|Ib��2D��!��?L���a/�1ٌ�� @5D�P��ˆ#�Ht�t���3��#�B0D�L�����0Nl��ih�4�TO1D��j��C&�\����	�(��6�.D�
���%v �M�.����!D���G)M-��Qg�����c <D�H��k?��|A�G�V�Ľ�S!D�P���ԅt ��z��ďmL�y{@?D�di�Æ
#��e��A;�36s�̈́ȓR�bٱ�h���v�\RA<<��I��Y��kϣ_$
���%�s�Q�ȓ|��ZE-
1!>�K� 9Q�i��E�������&��Kц\�tҐ�ȓ	�p!���J+ve��S�ۏ%h@��q���H��Lh (�"*�!�`̇�a��i�c�Ψ4��!	Np�����:(�"��٤���gW��d�ȓ$� �;3��+Z��DHۍ8k����LC��gc߽&���f	��/�̄ȓQ���5M�������<KTe��@+�b�׹M�X����Bl��'��1��	X*4N$(tŞ�}H���LrJ�HC�p�HY�HK�%by�ȓ��3!��+?ӆ@��A��+>v=��h�Ą{2�C����e�M�:R��ȓm.�*��D��ȕ"��JX���S��e��J��
�z�C���!���������?h2His��%N����!02z��-_񎜩W%��4�ȓFWX|8�ͼC�yb ýpT��ȓt�x�p,C
|����ա��n@�؆ȓ�4az�΄�#�&x�f[�>e�u��hq�<H��!pՠ��Q�K]\���S�? >L��/���FA�$�P��"O��2.�\\\(r�@�76��咢"Of1��&��8p�/Ş>�(Q�r"O(-jc͔��D�����+5���Y�"O�@J2� 3 ��A�R9��9�1"O]c�H�/n֕���ɒ|�0ܰ�"O��
a송<���qTʒ=)�T�"O�iѩ�"1^ꑻ���.j�ٺG"O<��J��o�R+s���ZZ6�Г"O�����v�$%��b����2"O�=�c�rБ:U��<�$Q��[�<ɖ���H(���r����@N�<���R�j��(E� o��EH�I�<���O�f��Q� \.e!�/�@���5��"����#V��z#�'���#ǥ�R��C�	�g���kTi�?K��́��b/`�DB�1��4#�S���؈�@�	^�QPo�{�B䉡o�t��L�F�\�5!^%C�	�f�M�/��01�'�(:0��>YdG�'�4p��\�^��;qAzH<��cF�l?�%��O:��o�=?�`�����>���@�+�p=af��`��aMA�-* }b6�yX�Ġ�Cڃs]Z\¤�Zq�
�0c�Â�b&;#��Y��'��y���*g�\҇��=�1�$�ø��I,rS2I�u;�lPe��J�>=xV�ҍo�tI¦C2����"D�l����*���L�I��a�4O��Y�쭁�l�x,΄��*_�M�$�>�O�PF�ǰ_�",s��:X8>%)sO�HmG�c���Z���`��ٵ���rz8{6�-`*��zqX\	��d�@�2��R�Xp��7-ӱ.ax��  ��2c�o��QY�B!xT���`�%�Hm�)� )\��Ox��eIO	�<h;���GH@�ї��|�6��z���*C�,z�<��`!�G��Q5�LdoO����'��]����%��|�W 7zk����\$!��3�I|fP��_�^B�Q*"�r�'��WL����x�Ա�aX�d�X��TD�h��_�?��H�"�Q�F�T2ew��� ��"�� qb޵��<�FA����TS����D@Z2�i�@�D�j�*�x��TXA��J:q���eȎ`O��@�^�b: ���(��E�*R:���D`M�I���')$9��i�n����ŗ=kXIZ��i�"G6����t�~	[ĎJ�$x!�Dݵ+"����J�ABhH��_�5k�u�b�+(���4K<��`3��|r��>N��9C��<"���b� �PxR#ߧ<*؄`��U��٠���`�$��c`�I �9����h�鉶S#�A��J�QJsrψ}2���U�&�� �^$�t�FJ�8@x���cgZ�;������_��t��ȓx���N\,htp�DM�iN��&���0�#זp��#�3�ލG���E�D��Bj_�y�����I��yb��d����kP�~��Ŋ"E�D6=`�J^��	4+t)��O�7E�^L"�IG#J=�� a"O촛w(?�␊��,{nFU���x�V���K��y8a|"b��@���b��Z�[Re'��=y�<%T��F�
��0́0�X����u����ȓ+��@���?�Bq��E������ȓ'��(���!	cdD?!F.H����#H�`.�1�i�^x��ȓr�"q�G �@ u�n7���t���r���eCg�Q�`�ȓf��t3c#��W:��OH�FC�Ɇ"��@U-�A<�=�e@	G�C�	�o�"dw��}���*��]~s\C�ɴk!B�A2�]8���C�߾n)�B��+�Mb�/�`B�5_q�B�!o�	�KC��ZqB$W%�B�2c�X��CjK��T�X�C��XC�I#
[�06�yz4릧�9e�C��$� �B�V�(�Xa^~��B�)� f��Um�
�|��a�<\F� "O�I����Cf����
pTQ�U"O�ɒ�Մ4
 �6k	1/�1P"O�yxp�K:�\����T(@�"OL�R89̊@��*p��Dcu"Ozu ��P�ݺ��G&R����A"O��5A�l�����χ!�dS�"O�lpt�ȴR�8����<{�uAD"O����A�9����0�Oh���t"Oz�z��$�fE���${d�(�e"O�=�tbP�9D20�a�9Qrh�&"OJ�����_Z<T�kM�C\�1g"OV4�a��,x\NIӣ�YgL�\)"O��$H�,CE��P�j�v~�@�"O�i��1nl�(�éB�Yɂ�iT"O��j�� "Fȸ�*��&oH�!"O�P�CA�*��5q *ۻJ[�{�"O9	�`�S���0h�REI��"O�0�D*D�O��@')��Q���;U"O
{Qo��F��w�A06�hw"OH�nĿ6vL�`&�ad�:�)9D� ���кD��[Q�ɰx��0��6D�@�s�A���%�P-_��`��b#D�����)<˖�j� '�DSæ#D�8���P�]����UD��Ͷ0S��<D�Dx� Ŕ�9�1�L�'��,��C8D�̺�X�/0H�w
�'td�a9D��RS��ht=�w�ԟL�,T���4D�����Ք9�VX��:tTB�K'�3D����dƫ40\i�I�<�05�3D�0#��;ܸ=I��D�a���` .D�h��Y*����F�b.��2ea2D�$�D.T�f�dC���T���f.D���ceW�P�ve���0���q�!D����([�?�DɛCiǤbrA��C(D��'IL���)���Bz�03D���R���z
m�O�<|��Yr�1D�ā�N�'��p��̄b��!�u.*D�#��Tr̆�3�*C�PKԝQ�/D�Sq��7�V��n��	 ��y��(D�8y�)��L�NaJH�y�i�Ū*4�`�T�G�b��8��e˙R�PXˣb֌N�x|8V,/�O�s#:^"�(�U�@s�����'�B�qd+ 5��	��8ڕ�pd��r��&(���Kw�!:�G�?'TΩZ�F��!����O��s���xE��e�O� l6�W,`�$�e���
�C�'�
M8�ʋ����6��p~ 	pDHP�q���hܸ��s�@b�g̓P� u�T���]d�"��Q�����IQ�i�Q�H���� -V%�.$�TdǕ��b�+�`��d������5m[�0R<A���A�]-џ\�G'׶h�d��嚯�t���`	G���Q��`��S�B��<�}�Sc�O��Ð�~����<7�`j�Ċ3K<ɲ��\=	�?9S��ߚx�h\�N¸\!�9��y�<��h ��-ڮ��p-ݞL�4\�"H�)���m����ɑ��v��	�&&���n�4ڍ0f ��,�����X��`�gf�M7�#����s�M�'s��`�c
�u�Jh��~8��qT� #�8�r��:�Z��4�?U����H�-H�)��
s��#e�?9���@J5�&G>.y2 �)D��if� \i��d����+V�D�d��(�Ƌ~Hd�p��=g�B�IF�ɼ�b���F���z��K0i�R#ѥ�F�<	��@+Ij�v�Ûh�$u�M�&����mL*��f)�^����Ld�<��lܭp+P�T�ҚU����`YV���y1��}�Q�̝.'��i`�*��1U#��f�B�A ���M1�O��d�&6�tM	椝���5(��d�=n�@1��S���8���Yp�p���?� b�+�`�h�Bݸ���Wt<iل"O��rU��8j�.��aєW�nC��+S\̹�Vyq�OG2qk��b��$lۼ�5�O.`!b�R���+
^��s�g�C�<��KY�o������Q�>86�R`�^�:����<� �s�������+!l���<	���@���裂G��\ڇ�}�����"�,4���C�ϝ%I���F��_�0�pp@��v@�n�k� �����p>��@�y� �б��8/b
� ��C�0h���B��u��Ԡ�`�IIà�)l"�	�$z@�����B��m2eB�%�!��cԸ��@G���9A�L�U��h�mڣInx2��X�a��;�`،��O�^!�;4 �)��f@x�|Qy��T�5Z\��ȓ
Kpթ��=�~�S�#��0!F��dWk�: ��IV>c6�C�B��
Ix͑F�#�5�.���@]�+���X3��d�~؇�	0i5���I�:��t�E� ��LQ
\��j�)N�}it�[����I6�1Y���o�b�f�;9���4k�(]�K�(���� v�XH3�P25���G���!Gq����Ō&��C�	����(cl��5ڢ���HM wp��{
�1���bí��+��jg8�'9��Z�H�Y�m�<{X�,"�0}�!�U�U]B��p��F�ݳ����T�P�E�1�{d�<	�,E�`�ϨO�Ԉ6'���rJ�C޿lɰ�s�'��ik�E��iIlH�c�R>o�r�S�9��ɰ�y�a�S�lmqal�+e���"�@C��(O6Pk�!��R�niE��E�?l%��u%N�^-V�Xֈ��y��L�6�<$s�Ǫy���FF�yRm�d�~Y��ဟ,���ȁJX6�y�/�4h�6� 1# XKLP��y�g��l�.8�C�S�k
r�P�5�yB�K� 	YB��v�Fi���M�yr��O�hmi�%�k�v�W�<�y�.;�b�jt%��h�D$2'�\�y��D'�Q�#ʈo��4�ŉ	�y�+C(h-T�sB�)Z����5l�y2�0F
�Y'L�e��{U'�9�y��SN@��#T�T�)�N���yBOܸYպS�:Q���&ף�y­6��H:��<<*��;�[��y�h�=7���F�]�(pT(�`�A�yBY-��b��#���Z0b�(�y.�]�D�j���$�i���y��?)�F��`� 	�`l��+�y"�Ĉ�6����K�!�1.��y2�@�6��9��I�}��l�D���y�e4NR0��π?sB���/ώ�yR���@�ۢ⋕K�ʆ�^'�y���J����
��˕B�y��/���K7.�0�8��
_��yr�Ku�&�1E�ֶw�)�"��yB��-<���EIЎ@����U.�y�@	z�Ҝ˶EA7�$I�g��>�y⍎.5�a+t!$�y��\��y��śr�xK!l[��`�Y��y��׼;�f9U�7'Qz8�FA��y�C��[ L|!�$w@����V��y��T.i��qkD��
�e�H͝�yRDC9N�@ �l�xN���bܺ�y��^S�Ԃ�����|������y��E1�͙�l
5�J}��B��y��G	>���._�0�����݆�y�Z�F_�1���T.]�mqW�yB�ܞX*�$�`bJБV�ޣ�yR��m���4����i4�yBg
7)�MA�I	�6x�vU��y�܅rf �Ӳc���p�$���y��F�xBT�Á���j�xi�4a�3�yr�@�By"R�7uJ���,���y
� f�"�ĉ\��X���d��P"O`��׮P!)D2B�B����x�V"O )����g��ɒᄜTΆE @"O�JD-�3���GB�*+��$�"O���@�H,pҖ"֯�6��"O.�q�3C�b�2AaيZtr)��"O�T�rg��/r(=$FD:a}��Ɇ"O�H�1gF�V+:-S�&�`�j1�'"O��I6���;�0�6�Ͽ�t�zE"Oj��u�
2N������ʒD����yB�]3Q�J-�W�?��\�B��-�y��OtH�bZ4�J�e���y�0��4h�B<��ȳ͇��y��Y�s� ���!�|J�9Q��߉�y���o���q'OW�sw0��e�7�y�E�:+�jT���_�[��8�"�1�yIH#����bSx|��F՜�y�W� ���U4s��C��y�KX�KT�ö�"x������y"Cϔ>����5�ƀp�����Ո�y��ڷ1�h�s���!h��xc���y2��Rz^��4j�:�)
1N܋�y�/�f�2mZ����o����e��3�yR��3���#m<f�0B�폻�yr� �'պ-8�n��S	�)�P���yr�>�tek�ܖT|"�Y- �y��h�4�ycm�*�fԙ1���y���:��M��N��fZJ؎���S�t�B�ش@R�f�ˋ@:4��ȓsJ�����F�b��/��s�4 �ȓ&�=S�g�^Ѐ4�4L��ȓ	e@q���@�x0�0k�D��ȓ�l5S���2��Y�P�N�{����ȓ?�Z��4Ɖ ^*^=8g�/i}p���}p(r�C�9��`���Ϡ�"=�ȓPR���c�0da�X#��%6����^�P 
�M��r@f�:� �q2�y�ȓV��M��O����CG�N��`��դ	��hG
|B�LR%��T��z��#�G�,��@�ώ?~���#�z�ZD,@%��(���8'O�1��	�0�'cU	���!��1jP�ȓ0�ֽJ��W7��dY��\純�ȓH�l���}�8��U&P������`�Zv�X&��d��@P�rUD��ȓ0%�I؛�"T
��p��L�ȓUp��o�2e�n�)�)S��fهȓ�ɫ�B�b2]1�"��w����ȓk�}YWC,zD&�h�lԗ8���ȓ��ѥA����] ֮Fy��ȓ*� ��GI���,�c�F�q�*��ȓ�F��n�jO� Zg��,V��9��E��'F���n��NV�݅�5������¹XA��B
�a�ش��nb�y��Y�;	����A
{N���k���Q�Փ
s���O� I�ńȓ|�D�����K�f�;��a��I����-��]�B�˦ʔ@ L��ȓGff��ȍ#�����(k.$��_��(&�_{F�䇓+��P��}y2��D1?$ {��n.D�ȓ]C` �
�l%�a��+U+�M�ȓb�
�3%ʘ�)�I��X�4��n���CD5%X�Y0q��u�&h��S�? �-Bs�׭]�z�HdF�����Q"O(��#� y�Ɲ��îk��	��"O`�1#�5�|�*����i�:(�"O0M�3
�,51� e�%IH��b"ODR��א~�V鲒
�2�ܫd"O�|¥�E�)`xI
BOP��"O��x3Q�ͤ�ci��L'���"O~T�d�jQp�hJ��c"OL�B���c<��*q��!X�p �"O���@H�nLPB�Q�u6��"O�*�[ m�n�0��:#)���"ON �ȣ3������t����"O��BUjE�k㐔+������"O䁙�E�u��]PB�2>��m��"On@cto] ip�ѡ�M�7H�0-�f"O�ʠ�|<\k���-�����"O�P(��1~��O�i����"O^u�,��i;�Ͳ��[�W�� r"O&y���6{�,��8k�ļ��"O(��bE9�`9��'o8`�"O�YJ��W6�`2��ӡ|���V"O�e�D�ΨWN���!FZ�l��əs��7+��a*ȑW1�tsaMѳ>|0�ɰN�h�&o�:1��ę�n9T&�Dʆi��,���: ��H��
�<Ld@�V��?y.=���t��D�O^,���b?�+d�6M@�Xw�D>q�6A�$��9B�rih�O>i��i^s���S	����U4TX�P���^��q�H�����I�,�^�H<�}2QN2L��9JܔO[0�I$��ly�P�qR<iɀ1}r�!_�� �c]�b�\xR�
�7A�6M�:�x��D��S�0
� b�o3la!���;*����d�ںGx��ƱH6.H�b��1+vj�ozxT� ��۞�2O�3��|�'l�0��u��l٤�]61�@��'ݞ����}��O�>�@j�+
�h�c@�CR������ɸ�:ҧ�'8��O:8x�eʜ�4��)�VΛ'��H��i�N���ƕ�%���	;H>uϧ_x��aQ�_͎�Q�E<vԌ�q�E�.���̈��M�׮�\2���S aH�RザF4�B��=<�F F����M�ƨ��U������Ḩ��ߟ��ׂ\�N9�0�'�2�"�w@�কc�	Ǟ&Q� �'a��I[�TBb0�tc�8V�����LL���B5F#I6���g���d�?Q��C&�p�H2��&��z%�T��cHB�.$�|�i>�����Nx���Y��!���/`~��>���KX>5�v'P���Q�OM2g��M�@�6��3B�$`DxJ|��j��e;`�z��ٖ@�����g�	3-�"<�~�r��1\*�A,6GU�бz�	�:����<|W���Z2t��Ya��?�(6�ʴbu�"���i��a�b�GEx�`�猶:.Q�l�ᓸM��u�o�yV� �Ŭ��~C�I�X�"a���*�z�#G��HC�	9#.<XD�Y k2v��!��V�C�	G��@¬F�izF����A�g�C�	3�2��$��kfx}�b�+HB�ɠ`��	��׮�m'�	��hB�ɐ.1F�t*
�{)H0��G�u�XB�-Yfya�T,��u��!�d�;�>͉���q{2YA���WG!��W�b��<y�B	$Ӕe)ԯ�#0!�$G�M�ѳ��H�%��� ���4!�dT&I]:���P9�hI>Sq!����8�ṠӃp��]�(�/�Py"�O��&�sQ��3L�j�`����y m�p�"l�=qP��ҤE��y2���v۴�z���>�Ur��� �Py�J�+$Ɂ��O�cŦ��'J�M�<�g��[LV`x�"ْC)���J�`�<� �
�K�����J�O; �Ƞ@�Z�<�R��,
4�B��IZPr�UDV�<� U�v�.�r0[��_�D�)�%"O��Aƀ=s�m���ϒ3}�1��"O�t`��\:b�#�LZ+p��4"O�U��OX!4�z5@ኔ-L�)*E"O�,�u�5A��*�#�MI�"OB������A��i�>-��\
 "Od�ss,'!��h ��[�����"O�ta�ҙ��5�B)M�K��B"O�q	���/:'$�B�M"�pA�"Of�2pbS�4�6Sfm�/�t���"O:(�eO>u�����ڟoȴ� "O����@�*�0P�R�Z\�i�"O<��1�K;�N4y����HQ�LHb"O��Q�S+2��T�X'c�> 8�"Ohq�e��.\���+�s	:U�"O�p��L��R- �3t�A�<�4�K1"O�́�-�]n̸;���0Ǌ�H�"O��0Q�Wʶ|a�dW=c�v�9�"Oh����$!#�ʄ-n�z��q"Op�R�n�.
&��ɡW4:����`"O����btlظ���� ��	s�"O�� {t����ۛ2��i �"O�x��ҥ\
"�D�7<$	 "O2(W"V�,DQ���Kz��"O@�cvHM��	#��ħ\�N�Zf"O���t�;H�F��G�#j��$"O�U	L�z��@L���KP"Or�C�o	�*�`���6A�}hf"O|�{��:K9�t�G��*l!bPe"On�`�E�y$�|₌4[��Dڡ"OްB�.�L8��Al˪2R�U�"O�P�E��5��x�"VI����"Op�*$e�v�0��u�[�S=����"O���i��M�-���p,�q#�"O�A�&/]&J�p��3Hʕ|!y�"Ot؂ԂÅl���sA_��� r�"OHP��	�(Mh$AJ���P9p�I$"O,���'��T��҇J^3h8��;f"O�5�@�CV���;D*���"O�%�`b�67��@�bI��l�u�"O���V'�j"�x:���	�P��"Oh��F�#D?���f�-|@ɢ�"O4�bg�4DR��0�G
Q^���4"Od̑���v�)��ɘB�N��7"O)���`�0X�e䑤t���Xc"O�@	�艖LR453�(^�`��M#v"O�a���L]�j9"�,f��$k"O�X	!L̐Am]3r�U@�"OND뀥�j(�� +�9��z�"O@�ȓ�E@�(�s
N8nMD�0�"O��P��+J�,�/�;��؋"O�����/1^��`�L_����"O� �%���R��$����"O��3��\ ��,C�#�Z�:A"O�AS����{7�4������@&"O�l{T�3�`U�k� |`(���"O��4 I�w7���ˈb2�j""O�Hr����%pJ��q	�G�J1�P"O��k�$�vĘBh�Q7z��"O���VJ�8Ey�<
��F�*�\�"O��.��y����r�_�S�xJ�"OrHy"c��	x(dJ�����Е"OT0�tK� k�r &Y���[C"O �Z���rm��EK�|Y�"O� ��qr	̩��A�Ŭ�:d��q��"O Xq�f�t�YH�DC�fĠ@"O���#H�pG��v��7�:�Y�"O��X�c.�9��b��h�h�҂"O ,�Ҥ�+/̖-��]�S&L|{�"O�l �aЅt�D(f�a��3"OHY���E�LE<pA邪<���1"O���5b=&�nЁ%��^���G"O�!�7��/WoByA��	���"OR��"��}��i��J�+����`"O��x5��	I����#H�O�L��B"OX�;5�+'S@���dE�p�.���"O�u��Ńy5޼�!S03�d�"O`M �@G�=��qr�^�"O�A%���$q�O�{yʍ�s"O�5�!h8���҅�˩"�\���"O�@s��$�J��Ra�� �w"O@ف�fҝi��J����� q�"O��iքf����5�Ϸ.N�}��<D����� �P�q&Hѧ{�VI�Չ D�HaB��,\���"��]�1-#D���իJ5Ztb�8u�:��đD�"D�[��KF �g]6D���TL6D��{��U�_�@-�e�NUx)���!D�� �� $vI���Q�03~��A&!D��b����q,ˈd
0���3D�|���:�xE3Q�	���5�+D��KPN����� ���r��YX�)D�Ȣ�N�	�D@@fŌ>�d\�!�(D���a��|4��ђ�r͜���,D��;��V36l"�RvNJx�t����-D�+'a��lj��zc
J�Q�\8�ׄ)D��X�#]�_ANi�gƺ�H(2��(D��X�J�[�4XHႍO^�/X�C�I�f�!b�#�NٹQ@D;}gjC䉙e������9���c4)U�6DC�	�A.�$���(|����g�s(C�	G�"�@�] &F��2cݰZڶB䉟�x�2f�$ Xt�S��d��B�ɍ:��xFd��{�"l���b�xB�ɜa��qc ӣvT��`�J+4B�/[~�}� *V�q Rx�WL��l"B�	-K��2�&^�	Cl��W+�B�	OjL�3�	#��զ�F4�B�'xBE����,����6��;��B�I~F�1�B�J`&<���G�АB�0Z�)@%��,���C�F"D�VB�	�?�2��Âe~�EaE�?V2B�Ɂo�q2�N� ��C�KúgZPB�5J��ze.�������*A�dC��u-�͙�e�.OU��P��=ZC䉹okdh�ɬJ��dK�#	�p��B�)@L��G�S�V��: b�Y��B䉠[���� .���j@�~�JC��/����(�;`h�"�e
;!K�C��/`.{��:�8�g��E��C�	 w�T��ך^P줠�ƅ�>Q�B�	sڴ9gϙe��th���0I+NC�	�Nd�i�LǮl����W49LC�	�"V���nS�J�����9BDC䉾w����@)����y�DL�C�I�U!L�G��h�b]����l(�B��1u���X���69�"DfH�.3C�I�$�d����/O6���F�~H�C�)� 6`h��O!1��ňE=#"OI��o޾80h��T�϶I����"Ov�q�O��.� dA2̆ N�"O"��W!��#=����J^����"O)сȕl�H��
�,���"O�@����-��hعYvf)�q"O:y��(_�k��9yHėgBܢ5"O�]�� �,�XY �ُ-����"OڐC�@� Ek��a��<{U"O챉F_�-�����X�Z��"O0A&�W�Q�$4��Q�:�zj"O� Ζ-2�R��G�\���"OR���%��W��}I�-M�;ߘ�0t"O�S�A7��
w�^� ���'"O��Y�~2�t�O)��q"Oh�0ëO/�D�A���L�\h�"O ya(LV���)ܶ/�J�r�"O�E��oӜ�dܨ�-8�*�!"O�Ui�-��C*δ7R�a�D"O�����"��!��I�8G�ɱW"O �(�$�(Y-n�pT�P�
��e��"O\��u��!�2� �HO"C��=ؠ"O��)qf%^������](Yx�R"O�<���ÑM������gT��"Od�ٗlӂ(�R�QL��h=t|��"O�ܙ����@��d�I%'1��@"Oh���,�aӢ�>}��� "O�̓%�F�)ZD�c�M�D��0!�"O���R��"L�u��%қFY8"OD<��B��`�>�p�KK�=�"Ozl�Č�{8`���*6�� "O��pqꉮo�p3�kV�>��͊G"O~ 2i
� ��� %��,����'"O�M��5B|���3i��H���ȥ"O�9�L��Y��M��h.'��ڑ"O���ֹe�&u��AA9+7�a��"O��I��!R:�ȁIj�4��"O*1����]A�@��a�����"O�4�s��ku��B'U��\+p"OƁ��~f0M��H:B�ܰ�P"O�$9���lPL�c��ϓ+��A�"O�e{��?����#����"O�K�j���Ǧ�;���rf"OP0pt�j���4�҉L�8-A'"O&Hs�CO�O�|�	�h_x�p�@1"O䨢�.�P�X��pmM�a� p�"O�i:AoE�g��c�k۵Vt@@�"O�9B��҅� ��Dʄ ��"O��a��P0|�R�	 �?��Ƞ�"O��{�c^�PD�)"�IL�_�{�"O�q�T�Y`´�H��,Ԁ�"O�S  
  ��     �  y     a+  �6  B  �K  V  �`  �j  �r  �~  @�  ��  �  ��  �  (�  j�  ��  �  0�  r�  ��  ��  8�  {�  ��  �  ��  s�  � ] ] �( ]3 �B N 6U x[ �a d  Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�� |d��"O
`�(�;���8���-0��1%"Oj4��ND^[��"3/9�0|H�"OB���H��*�ʞRy=a"O�味V�!X��!&F�:J�$���"O,��a
���C�Ą�M�"O,$3%o�-���p���+Ն�:1"O��ݢ1����`���y14]2��i�<�6��{_���c�H�`�fX�$Kn�<��A̼VI�xR[�)�Ć�pඤ�ȓA5��('nߡ4�� �)˩%� ���,��r�؊b#`T�eT09���ȓ!�b��g��}�8�F��-? �ȓ
K|m�ș�VṔ���2�%�ȓ"R�X�j�4JN�1�˘X�i����̹	_�jZ��1!g��zܶ��ȓgil,*�J�
j�Ne��i�J%b���f	�(U��:���G��$Y^م�~r�� S�%T"���k\�jx�ȓ|4�1�îJb��@ӵ�ݩn�V��/[`�"�v4�R�!ʎ<��M�ȓ`:��z�ؚh�J�Z��$HY:	��H��p�m�C1��!��B:��0��EnjZA V;9����J[
2���	��4'J�EA�IVW&��~�(aZ��ӹ�>� o�Y�|�ȓ�f�A�
Ο7�H��M�$�����mޠP����/���ANXo*�ȓTv�����{ ��-7�*h��I��sB�8�8���3����ȓNe*M�悡;������X�o��!�ȓ'lj�#F�m�+R&;�|��2)n�C��0S4���T:
b���:�0!��e֊��)��ͷV��,�ȓ0�&�8#���� ع�L�����;�P�AFd���,w�6d��r�EQ�( �gVlɦ�M,H��,DP���|�I	$G#\���ȓ"�)���E�B	yt&B�^�LɅ�4�� ��eëF�ڙ��n��R�p�ȓp`@}bŇ�=�$�AUN��P����L��p���_�a�)�Y�!��-��u�5���o}�`iF�@A�p ��F�\�0��[���IF/5���k>bTؖ�;K'DT`�^��@��fnV���Y�b�lI��	����ȓ,nٛ��Ć3���kC��8�m�ȓ'� I ���x<=���޳{��	��6��(� N�����
�y2<��ȓx;6q��I�
=  yG�O�,�!�ȓW�>���.؜ɰB��;�����`9"�ˁl�$@��- G��D�ȓ���zF"� ~\�`%�[�ل�E�1�N�;f��PG�.
�T��=���!k�AμO�~m�ןOP��ȓ[Ȧ8vh�;Q��;�ȝd(���Y��������O\d
���v��Ɠvĸ{�`�?t[̥�2wp�yJ	�'�����K}�&�{ V ��{�yB��g�O��LyD�K�gj��B a�5�
}��'ЮH� ,��`��J��hE�I>����I_X�%��cH1d�\&�;�!�� p�Z��  h��ŏ��x���i��Ć��N<*5���,��|	��J=si!��' �n,��,�F�0%%Կ>S!���2W����mI��2�e�?M�/m�|�iW�l���vO� j�<����0>�M>�A�7p�-�$ؼ]�4u����K�'�ўʧ�*]�`�]3�ܤk&c�ypL��?�`�'�?]�V�I���F蟒 ��]@4��, ��"~�	3=L2p,]�MC�uAB���w(n�=�Ó#�
̱v��(I��G��' �M�!��~�R7e"T!ѷ�B6*����1�0>yJ>YbJ��]�*�iB#����iL�I�'�a����3�ʤע[(Jj�r�eN��yR�21(���0��1�	�-��?)%��a�Ob��jC�S�mD�%3�fE�"�`��"O�m��"�]�,B��Ko��c_��Y�P{�O(�^w3�O(�s�(�,������;r�&�&"O�ͰQ�N�}R(�qV:5T�IA�x2�<�S�y |�e��'yT��,�k��م�2VV]{َ-��9� 
ƕ3Z��ȓ ����A�-+�őסO*�@	��<A�d"Тd�La�EB%XUՇ�Z ����5!���R����ȇȓ2��JX$�����c^q�ȓ9�����g��hc.�P�T�:۔��=9�;;r���mԜX����F�E�%���	~�'8@��b)!Q���!�G<<�8s	�'�"aq�$ω�0��G�&�zH��B��4��O��ᯆ~�i�q��0Y�n,0�"Ol�	��˗'ۊ4:%G�~l�8���1lO���ܷ=ʈ���d~h��"O���A��`�^`h�BV����4%s��"~�	2�A�.�?eAB8�#Ь_|C䉡_�e�T&S�<p����)(gDC�.Sظ�Ci��4��)q�k�Eɂ��D{~2�C��N�r�	�sͦ���ɞ���uX��c�M[�@t8��1�F����RC%D��s'J��1f��nO�K��?D��� %��x�h�[4#�$>*�lP5J?�8�1Oz�'u���7�21C�51f���Z�F������w�ǽs?b���6&�(�'���>a�"0��,�	�^���K�N]�H6j���>?Ka|rU��+�i�ji1`��G�Ty���hs�eB�')�����#~Jȱ3B�_Q|��d ��4Hs�����t$����V�>�
�7q͢��F) ��@P�Cn�:��O0��p<YS8�xX�A�,j�0�BA��܀�'�z@� �%c��5B�ʗ�.l�u��'X�`�U�v3{�B�1.[�H��'����*)�b�ς'��y�'�Ty�m�9:��Шc�%Tr�!�'���
+��_5�x���Z�y�D�\r��r̋�,��`���/�ēu<��b?53��'�����b֜�%D��c� ��d�`R�zv�<{�,�>�/O�'��g≠e6�8�$�R�ԩ�êV�q�:C�ɪ�B�O��P� EbdO$���	 #p�H!�� 33|A�nt����d�>IS�	"y���H?�d)K��a�<1sO�#7 �K0�W�$�h�k��DG�<�$�/I;0��$�44�{��B�<��&U>-&Qф��H� +��i�<a�$�,v�Y�ק�h�2��ol�<I4#�8�0���GɚhA�`P���h�<� ��7+ՁF"�E����BQQu�'�$�%� ���K;�����"�!��|'b<�B���?'���"�\m!�1��3��T5|�]�0bڊOd!��݆ �y򧫄,��qWJYc!�dS�|"�u8 ��Hmv�R���s_!����y���Ti��%4H,&B�'R�'.����
/\`�w��C�pQ�	�'{�(��⏣CWm�� H�nm�	�'.�ɢAˀ/8�4X!DA4-�ȰK	ӓ��'��穂�B,������"�T���'��	�Ubڥ/k:(�G�K�Q�'Ƙ���Cߤ*ɠ��G�L�G�1q�'dr&�|�����zjX��s⌗�y���]��ff��F)"�1��$�y���pI�����D�9Ɇ͚�y�-�+X�!�W�P�ZdĻθ'��!���!���u�� ��IN�	�Y�!��*��1�$�2�̙����y��O�=�O��ԐJ^`�D�d��P2��'�'�v���/3O0���%:���_��%���O,��B�B%{S�v�*2�I=����H����G�N~���%D�'?��ϓ��?��M�>�!�dǘ�Q����N�y+qODm���'I���!!��@>&8����<yx�2�"O�T25ˎ/5^(Qڵl��{qV�a�A%�MËy��?�=�%�Յ��堓�I�E9���[G�<�� �~ш��bŒ5h�$bL[�<I�f �f�8��ኚ5t_t�z`oUM�<�R� �o�!�Q,��>q��$� H�<I�j�/a�H�rp뇥FmZ���A�<A��0j�4��;o�>Jc��E�<yRK�2gU��f �9Y����I
y�<i��_5,ɒ5r�X�f���)1�V`�<QB��87�d���� �n��`�<ѷ��I�<x G�\��X_�<��iR�t4d3b�:��Rb(w�<��m�;���(g����q�<!U���h2d9�FC��4:��s�<Q�h˯=*i�gǎl?\)����n�<1�IHZ��*R�
,)��l�m�<)w���v�8�3e�x;��	׭Um�<١�E�A������Z��haҮ�e�<�E�_'np`��MΝs��)Q�ke�<����8����7ڑ
}�1RS�d�<���]�Ĉ�咲''�Ʉ�XI�<��L��?=���e@���LԪp�H�<��L�5����e� ��%�yBN��0=b&m	�^%�<+Q���y�C�1���� "K��@���	6�y�ϔ�	j� �ňY�JLmzb�y�,ƒT~�q;'n�YZ�!��%N��y��Hg�,�ҵ͜�I��C�l�(�y�	�M�`}B�ݰV�Np[6C��y2l��y�M���Y�@��`���y��*q T�1�X/W�X��㟈�yR��(S��7M	"��j�c��y�e HT��˥@L�~��1���y�D	s��W�/]ʘ9�4�:u��B�ɏ )@M	5�O�HK��yA��<w�B�\j�U���C b�0�!ǣ,��B�I%��8�������$��ӦB䉴���S�IB&;��#'�W�<�B�I:E&�h�Åז�"�rTnA� *�C�)� �Q�gQ+�T��'J��mv�{"O���%��ۜh�#I`�4 pW"O�@�nߧ��0�ǖ{��M0�"O���w�HRG�וB��<(�BN��y���v��c4�,�J�D�?A���?y���?���?1���?I���?��B7"�v��"l�Go�̢#,��?���?���?���?��?9���?Q����4<s2n�$���F�'�?y���?i��?Q��oǟ���۟`�	Q�3��� (f�,.Ab� e��O����O���O��$�O2���O��D�O��ˠ(���QC�X5�=�0%�?���?����?���?Q���?����?�!)J>���S�-Nh#�X{Ђ��?���?����?��?A��?���?)��2$��C��h��e��[�?)���?Q���?��?9���?����?���0^J��4�ѠU����ug�.�?���?���?��?����?����?�,�6q���kL��d&�J$������	џL�IşX������Iݟ ��0��u�i�9_H���GQ�p���������	��	۟ �I����֟L�Ɍb����`Ys6��r�	9����ϟ������	����ӟx��ڟ��I�G�,�:v`B�p(\x�@�I���I�0�	ß��	П�������Ο4�ɨ&���
`�һs�h�iA�[�%,�)�	��H�	����I�D�Iԟ cٴ�?Y�	~xc�Ր�@ũ�*��,J,фP��Iky���O&�m�XT�Q!K�.^bА���I���>?���i6�O�9OD�n�)���G+?{�\�i����+�M�ڴ�?g���'��Q�Aȟ-+h�)���H���W�T H�D�!�v�d�O˓�h���f�;� ���RY�����b�'�u��6���w�<a � ]9���$$#��+c�sӞ�o�<٨O1��`Y'�qs��:�̉"�o�%L�S�O��6M�(r���
�Ժ}���=�'�?	'�O�l��@�`�ܒj� �k��<�.O��O��o�
sܞb� � H�UQd�F������oV@��a�I�M;'�i���>)r��gdh�ݫXd��Ქ�b~�DP馤����ΘO���xZx4�D�'��M��MT*
��gm����^���'��9Oްi�̼��A����(';O��nZ;h���E%���4��#dk��r| �$�VfưZ59O�]m���M#�V���b�h~�B�4H�Z��^5[�P�ɖF�[���`�$��&�u
��|�T�b>c��`t�G������*��[�@镇.?�3�i.nA*�'7��'i�4��@�JѾ�!"��$8n�!Dq}�o�*-nZ��?)N|r�'�R�A�zr��iDX���#�LI�h�ggG���DL3-HQS���*u��O�F�lxٲD�!�lQ#�9i�L����M�ߵ�?ɡfK�.�TH0��@5A� B����?�E�i��O�t�'B�7ɦ�H۴S�peY�
K�0�	+4��(4��T@��Γ�?1ڜ
<I
�BՁH-��?��]�J�y� Mu8*�a�.x�D�Y���p5��6W��%���{�fh�`H�ϟd�Iџ���45px�O�26�-�DŖ?�!I�h�]�ɧ�F�P`%��۴j%���O�戃wFͮ�y��'���PKG ��B޶w�4�RE��8.�8��e��&�ڴM2mK���PĈA���2 ��G爔��ǈy���� cQ�u��I~��c��W"@㨰SUbS
{��q���"L$��cw>_9�Pw��m9
�B��2`��D��(��rPB��2�K ;'�Q���K�v%W��+��(ңBަu0J���U�~Iv��
�'+���F �O�&�H�� 2 �H����'2�]�p��L���: L��@@�#��ت��1��0@�A�\\Pꉠ0��� ��:�� X��Ì(�� C�O,M]�X�pj -*�!q&���4;7��2u���m�۟��������<��@�I>S�I�o�TW�DHO<���?	�^���	�-o�)�T� 7?�rdLQ���VR����O��M�`X?]�	�?3�O^L2Q-��z�M�X��d@�i���'��� [��S֟��3�d[�<�||���E1w���*��WX�v☰(r87M�Ob���O&�I�g�i>Iyg�J��k�k�GW@�	��Դ�M�tO՘��D�O�����1O��W%)�|8��W 2[n��j��T��n�ϟ��	��RU�R���|����?��!�1o�v�!iW*Kz
��0�V'L�I�P�ɻ=�c�������7_����e�ߑ02Tb$%�'74����4�?����6����$�'o�Y���5�*r���˃�4j�8�H����MK��XT(�<���?1����+q�
�z@
�P���%��u�j��P�m��ڟ���{�ZyrAޓU��1U/®q��%���r��y0�yR�'���'��ɂ:`�љ�O�i��E+�	��Ì�J���[�O��d�O��Ľ<Q��?1���J��Z�nw2��3G�X5���N�����O\�D�O^ʓH2� ��ԥG��Pbg�ձa�5b�
̬a�P7m�O���<��?�`�R�rrJ�
�h���$7BH�Hf�nZş���[y�&]>�r���$�k��:-�h�C�?�q� $�-	��VW�|�	ǟ�xe"�ǟ@�s�B! �l]1y���h��t%Z��iA剗d�`�0�4bn�S����Ӵ��dP>��8i@�^�.P��ː�W�9a���'�d�)��g�I�,�8x���Q%�޼b�o�s�Z7-Q��1n�����	柴�����|b�� ����N1�hUZ��Ҹ|�Ҽ12�iL�%�S���	џ��3�Iڟ���K�Z�1�O�9s�4e��&E#�Mk��?��
� ��,O���O�����\�r�	=%ѰĠ�/׳Y�D2%�֘'���'��Oh�$��|z�Ñ�:8M� ��	��D�U�e�|��ָ�2��?����?I�{&�+BG\�dg[�K{α��5��d�	���!����I�X�'�"h�j��=�b�T8Z�!��c5dE�]��IΟP�	p���?�Vf�&M7�q�� 8^�	��". P+��Po~��'frT���	�/)u�'#��k�/\
��;��D�<.FUoZ��I˟��?a�6R�������!�Krh؈HPd�,'�Vt����>1���?1/Ob��[b�ʧ�?��e�{�NX���%#��{u���[��v�'��O,��%XRjqa�x2�ΕP+f�G�{��]X�`���Mk������O�*�Ǫ|"���?���#�유�ʆ�c�y���Hg�l�d���Oq�ee��dE1O�ӂ�N�A���t�F+�<�$��?١-�4�?9���?�����/O뮊91~:�o�3,��a
��'*���՟Рɕ`��b�b?�B2`��oF�H(��P@���B(tӴ�m�OH�d�O ������|*�����!%�lv��X��R�t�jXq�i��l�r"Q.꘧��d�<^�Tp*���H|FLN2x�nƟ��	ȟ�K��Zy�O%��'x��Pj=SL��ڀ��,K�(�<Y�˅-S��O���'��$�C�mKS�_�ngf�P5�*���'�hh8�\�t�I��p�	wܓ/6����&�=!��C,[�{g�,�'ꄱWGG�����O��<Y��g$F�	��z�l��3��1=r,$���H��D�O����O����	2��!R�'�W���p�A�x�W�ٝ���?����d�OnDA�?Y!�e�	1�9b5+,Q8VpSB�`Ө���O��%��ty�,_��M��� |.T
�i�'=z��P��z}��'vrX���ɾz�&�O�rT�",�L:ӮD��"�A�)Ϣ%��6��O��0�'F�,�I<Q �F��Q#&��&W�&d�Φ���py��'�V�svS>5�	������t�P�r��N�p(�$��73:=B�}�]��SD1�Ӻc��P�f�(a;�n�T�:��D}R�'!�<�D�'1�X���SqyZw�xp����b�Z�۷
�Q�Ot����ExJ|�W�Ɨ��p�k�T���b������q����	��4���?m�����'��{��K�F6t}�5�)i.�#ƾ>IV�S���ONr�K�]��(��C�mGH�fc��gw�7��Ob�D�O��!̬<�'�?��~.�*4�,�YCK
s�>���k�H�#<���d�')b�OT(�ނ�R��A-K�@
�Q��i��-�3!�I��|�����=� ӊKP���2(�#i��Ż��O≓8-���?�����Oh1���E�c�B�p �YZaӇ��	Fzʓ�?Q��?i�R�O� ��O�8������ԟ�&a��ict��O*���Ofʓ�?y�������N�r�9�S�M�,���� 0�M���?!����'��ɏh�7m�=%�8:�c�?EA@�r���_.�I����oy��'V�X>���xC��S�+&J���E�B���� �?���a����ƭTo�	 (~�p)!�/6�`��ûk��7�O˓�?�Q�����I�O^�$��܀�O��_�.�SFF�8� ��r�WP��?���Vy��<�O݊0�T�	]�E��7VH(e!�Op�d+|.�d�O�d�O��ɰ<��g���k�^�;��Ȣ@�S����'��蓭&E"e�y�����9�"�j��wN��B��M+6f�'�?���?1����,O�)�O�ȡ��^��� �CÜ,�TJ���M#�!̭E�:�<E�T�'���y��9]�t@j7��:��pu�|�����OL��H�`�l��|��?1�' *�H��(�.���&�t�)�O=扡t�,]�N|���?	�'��`'-�*�>Ma�N�rJ*�޴�?�ADA$����O���O���(��Y"}a� 
WK5e±B��>)���7%V��'���'�I������?J]�0O��}������/Ր$�'o�'N����Ohy���H`�tj��K]I���A_,lDs󙟰�	�`�']Rӏ��)�,@�0�$!_�+���Z����'�b�'��On�D@�M���´iБ���ҩ���W���B��@��D�O8�Ľ<)��)%ڼ[*�(���4�М�b �#-��J6L��lZ��?A�p�����w�	.�6��
��$��mܲT�6-�O��O��$�JRn`n� �I��4�ӳM�fD���=
0�4�ci��j����4�?A(Of���!��O���|n�:�0����0 ��|�ѭ��l6M�O��d�9;��n���	����?M�	=7�h��&�	:՛фՕN�^گO����,uŬ���Ot��|�J?�
��">z��Ά"}]LѠd,sӶ c# ��=�I՟8���?�����������68$W��=%h���"S��M#C���ĭ<�g~�O�r�<2$x�QF��9�8
C�},�7�O��$�Oؘ-ZԸ7-�O>��O���O�[#
8MC�mW<�s�j�),�IRy"a����4�x���O���� %�)�sH�C�(��?<O��m��8Pt�	��M��?���?A�T?��S�? ��@�oUq�4�pE!x��qBW�����7?y���?Y���?�/��ԮF7,����bּ\R��0Tm�9�yoZ����ӟ��I7��)�<Y��6َ�Q���|����-K&u,�P�%�<�/O����O��Ŀ<1�G�Z󉕈�r�%F�N�X�R&�+BO�vR���Ivyb�'���'s�1��'.��Z�/Vd<5w`B�k���Ajg�����O`�D�OJ˓P�ҵ{Q?��i���2���@��3� �i�� �sd���D�<i��?���<�����4/�D��7��d�TLi7�מW8&qlܟ���ʟ���1�")�ٴ�?��?Q�'?:u��; ��]"�")pnc��iT�[���I4{ <�n�i>7M�>�y�Fl�Vł�y�Ն	��&�'��
�(9��6-�Or�D�O����@����	��j��$&�ز�ʒ�[��@�'!�["P�B�'��i>]�����&�O�<>8}�so� &_�D�@�i��xzP�gӌ���O8���z���Od���Ỏc���
��� ����p`��9� ����'��u�S֟�@�
�8��-���*�ȼ��=�Mc��?��ƶEp�imR�'�"�'ZwD �p��ح�6���'��R �m��4��5K���S�$�'PR�'%�ͪ��A)��� �Դ�:P��im�����+a�nZ⟨�I���	������x��	"C=���� 9?�����>YNV�<a��?���?����s�TI�q�Bb4����B��`�IJ��Q�	��\�	ǟ���&ʓ�?�cm��T	I��ĨNj,���ʈv��͓�?���?���?a/�T}�բ���=ph�	A�Ucv@� Ӷ�Y M��M����?���?����d�Oj�#�1�V� "M�4R�tq�bw��	�Ģ
ݦ!�	��h���P�I�����Mk���?0MN�"e��U.�N5���G-|����'2R�'L�	��4� p>�'��鉔�ы?oz$�)]��&�fm����O"��Oθ��)V㦹��柌���?%q���Z�P�J@�Y@t˶
T��Ms�����Ox���0�D���v[>7M�|D��&l�� �����=U��_��3��M���?�����W�֝�Q@�a��6T���A���$67�O��$�*w��D$�d=�S�"��ѓF��4��u��+Ξe�(7M��At��m���I����S���?�����]�쐹1�Ҕ_l*��v1��,��yқ|��)�OXU#��_*c��|@�D�������(�����ڟl�	�%#�ُ}��'h�����I��l�<>+��sUf��h��|�BK��yʟ����O����@@�q�e� ,g0���"^8Po���|K�*���'��|Zcn��C�8Z���Q(U�@H8��O���1On˓�?����?�-O�m��EC�(_Be�6aK�;�<s�.-QPĩ�>���䓇?	�%M`���B��
���PMʸ�4򋅨���?a��?�(ON�@��|rt&��z̙��l�.fr�{���`}2�'���|"�'�NK�cl"NW�|��s�)A�Yϊ��Q'�R���?	���?a/OH���Q�S2&R(��&_
;�^|;b�KM��ٴ�?�I>���?����?�H���ab˗S�Q�� S<e~�x��c�z�D�O����p�����'z�dc�g�j�q�.۪6����aN�m�Or�D�OT�9OޓO�S�QZ� ��I�J��<QskJO�6m�<	���P�fΠ~�����7���Ck��5D>M(2��2T��x�ah�b���O6�z��O
�O���<�"�S�Zy��cۮ]��i�d�Q��y�j��O��D��1�>�"�?|�f4Ȗ���>2P�!�チZw���"�O��?��	4E��,��	�m��*q�_�4d�۴�?I��?���0p�'�2�'q����n�lR�
\�mXc`
b��|b)�2��|���O�����-cJEٳ�8n���01�`r�4�?MЇg!�O���;����\rp��1O�ܩSK�`R�� $��]�	H�	۟h�'�ey�/�82��!˵�<X�v�;�Mê`4O���O*�O���O<mѕ��/��I��6;��8�;�d�<y��?q���׿J>��ͧj
�yt��.mt�Q��4.}n��'���'��'���'1���b�'�<����+[eX ��@����dG�>���?1����$�(��%>�!�!�=G�j(U-"o:�CǏ��M����䓮?���h_���>1��
���fL�?} ��5ÚҦi��ڟ��'���Bk%�i�Ob��	��F(kUf�0a<!.M�$M��$�|�	ڟ候ȟ &��'!�����!�:��i��5��'�"��K8b�'q��'~���''���D�$ٳDa��wx�2�(�K!���'�b*V.g��X��y��4#�L?jHq�C�-Wҍ��ʒ�M�v��|���'���'
��=�D�O�`�EbJ&hȸ�����Z�I��}���-�S�O2�ɎKՌa9h;3�V����1k�:7��O ���O��{�͋g��?q�'���C�bS(.��h�O�=�V�b�}�̘���'.��'�՘�<����J�U
�"0 �)+�6m�O6��PJ�]��?O>��,cr����
L-{�	N?s�'9|�؋yB�'xr�'q�I#A0PeS�ֺQN�\��'��t� uPq�T��ē�?������?���U���R��0JE)Qф�� GB̓�?����?)-O,����_�|*��&��ɃR�\>uv2�B�.Ps}2�'���|"�'�RgL5��� ��B�A�6�f IP^�Nrq\����ʟl�'��7 �Sɟ��ਅ�E"D�3��@y�*t/�*�M������?��MN9��P~�	�~�	��m�� 	���C�9��6M�O��Ļ<��ܼqɉO\b�O�y�#CS�H�t����ÝQ�Z��6n'�D�O���I��''�½%CC 3��!�!A<\}lxy��!(7��G���'���0?�bi�}kH9��4L��9�b�¦)�I韔(�#+�S�'Uw�x�f�X�v��*v���4mZ;8:�p�	��,�'��\�<�'p<�C+���`�q�O�c;䔣��j� �B�E��3�1O>I���pt�PA.�$G4���ᕗC\aIڴ�?����?�1�(HJ��d���'��A��.����q��$J"�U$�Pgdb��qa*\��ʟ���ן����5۬�	��ak�nH!�M���|��!�*O��O�|oM�I��T�ߟO�ځ��͟�	�6�Jר��"�Q~R�'�BQ�T���a�j!�׉�&j����js� !0d�fy2�'br�'��'cb�'0�[e�+b��A��A	�qeG_�\�A��OL���O��Ĵ<y�iM+O��i��06T�d��4- �)��f�>���Ov�d-���Ot��^<:��I��LZ�o,r6a��-S��?���?�*O
U�S�Pe�'�6�1A��D��ϛ�8�F���4�?	O>	���?���Mf���(��F��8%���J�X�h l�ԟ,�I�\�I:7�����`�'��G�#r�� ��ɜ B��*�O0�$�Oܵ��/Ȣ�1O�S*y%R����+g��X ֣U^�7��<aդYT�����~�������! Ґ�豀��*5ATO9���A���3�$O �����]$/�f�p�A��6�	�]��'+���?1��ß��'�@ ��*��:)�t���
<�,���*k������Z(Q�1O>����l�P��Œ�f^�h#�ȍ>I.�aڴ�?����?�W�OO�'�"�'���Ǳ�h-�N�d�[�E�Ρ����A�zG1O����O����dNEj�.߂m	�,Kd��C���l韴����,���?a�������g�"d����>r�"�)Kw}����'K2�'�S����J��;�4�@�� T��"k[؉�K<����?�K>���?�`��<k�-X�5��UP��=nĢH�<��J�S�P�5�Ob��R��Rj:�|�%�ƽZ�����=k�l3#0wi�j�
ˤ�����Oʠg�Qꅣ:�*`s-���(O|���БG/P�G�0c������1\y�����[��
q
�<3��Mcզ�������\_nA�cF,�.-�5��#��h�d�*!N���hߩo��9����k7�� Q%�2-���Z���&Kdi)F�_���ˁE�=^��s�NK=.е� ,�D��ٳƥw���(���1���62 �JS�!\���#�&l����\b^��H{�|Y���?Ic[�nW�H�D#�f,�hP����|Ruƀ�q�pd('��(/��!���ZQ�$a8�	;��� ��P��<�񟚭P��8j��I�f�ߘ%�D��%�>���L֟X*�4�?)����'�?��ˌ'��� ��ֿH���tּ�?1��?����<�W�Ո+�Tĳg�&�hm�.�|������I�qZ:|R%/e��}#�D�4#���mƟ�����c���9��D�	���	ݟ8	[w�8Q�dW&�a�F�)�"��^(_K��2��O��ѱ�N3p�1��'��ڂj'K��䩤�8/�"�qf�����̓GExjܑ���ЂN��4CI?u�t����.�@R�С�H~yF� ����-���$�O���Ԏ@)6��Y�x�I;�.U���g<�@�ꀁd��Ɠb���kg��2����տt���'ς"=���?y+O�}��=чm[�
���B��ЭE(ubU�K�{���'KR�'���]��X��ʟ1FO��Xl���Qc L� �P�}:>����'���S�ʑ;�"�!�ӯ1Y�l���'E�й � ��Q��ɣb�B� �BB	N��KV(�AMj�(��O��l�x�'��O�'���$�k�fɝA^�Y�'�%3����*&V�$3�"E�m�� W/qE�Q������۴�?�,���ۅgFߦ��I̟���Mٛ�b��W�I�yW�݊�ݟ��	�.���I�X�'"�����H�Ɍ2J��ZwL�<o�x̉�a���&��*��O��W��V���1�S�@7�8B�'YR}*��p��'�V��6`�f��\���9��'� )(�(\yDq�O��O�Y�'�7m��`$��H��<5�C�ٙt��O`u�.����Sڟ��O��	�4�'U�T*6eʥ��䊑V-tp�jS�'3r���" �mC�A� �cՅ�O�S\�D*��as�p�G��4�w�Y���;Q��� ͪh�0���]�?��S���~A��ץ�e�q��)}B�K�?����h���D=;��I�D��h@�M�v�W<!/!�DO�1G��B�#v5bY:�&D�w�ax��+�y%*H�V��0a_
D��AΏ+�<��G�i�2�'�nZ�=������'�R�'��w+b]��	J��ҕc���0,+�Q#c�8���V4�0EF%�3�DUQ� �Y(�}':YrC�H?--�y6�_�/����6��B�hB�;�S� (D���5��  t�Kۀ3�VB�޹:&�]V�G�	�8&����|���H���
 ��.�d�9���y��ޟE (Q��7����R7��D�^���� )�M
������LŰ#�N�ȡ
A2�� ����O���O0�DKӺ#��?q�OV����7,�1��c��L��=2�ʅ&�x��,Ny�G�͐F{M�2CEe�x��'~��bD�v��aV$�-D'��h&T�?)��Y��a&����TC�FMc����Tx"� fH_�P��� -_��D�<���i�'�.�@�e�6���O�����P�4�h@V@Ȫ37j�Z�h�O,���Q����O��?���)�є�<M�m
�%$(�&���|z�xBmZ���'�(���_;&�`eQq����Ǔ�$�	��x:����J�OU��D�R"����.�I
�BG9A\�H��͊s(8���Q�6	o�u0���d����`Kű@��'
|�ke���d�O��'1\R1����Hx�X�c��� N�U+&�����?����8v��a���,�h�1�%t��j�t�ȃ7�r�a���K�	�o���9D�����ӈ1����ݵ��l�D�:�i۝0�P�s&aV=z"$��2,G�9=�{�D��ɽ�M���?�M~b�`E�|Š��2��9 gaٴw�����?i���?��?�n!��"�	q{� ��d.1 :���	�HO>ђe�Ǹ8*���v�L�w����R���Iޟ��ɱ�B�j�m̟p�	��\��'�ue�-�0�� �9Ө���ԑ^)\�O,|�l�~Q1��'�`��M�I���ђ��A�8X�U�*���%v������L>���`�r��ui�i!ĥ��M����z�z��؈q�t��Y���ɃQ4�-�恟|.X4b���6f����|ܡ�$��=p�!k���`�܀�'�#=!�'�?	*O�-s��� %:�U�P,AȖ�+f��_� q��O@�d�OV�����#��?ٛO����DZ("ќEi7aӟ{j�My��_�x�W3�f����ߪVl`8;�C<P��0�'�n��`H
��� k�.O�L{�(C#�?	��'*��T'�5X�X�I�_g�r]�'e��� �5$X �1G��Y�ͩ�y¨j�2�O"D�զM�	ҟ��Շ"kK�h�GBJ�Rvo۟`���O^|���0̧H$n��G�I�ohX `փ�*���p�/JJ���d�t��O�л�(5� R'߾;z���'��b��[��'�`�!䧝D�T�fjA*����'��*�'J�vB�-A�;�^i��'b�6���av^�I��ɽ}o����ΛgnʓO��8`��ۦ��	⟐�OHT���'7��@���Q��!$$��L�*��'��l�	w&"�T>�a��� =}�^E����do���O����6�8Р�*.�'W���[�v�H�pG�=jxi�OV����'\�O�az�#sn�X3��T6V5*�"O@d��lWS��́�	��������'D�#=9Q!��n >� 5b»H����4��'�v�'�b�'+�Q ��m���'���yg�@-���dc��sT(�r�m��~g1O�`��'2��婅9U�^�Y�C3h	
�:�{Ro���<�g�(*�	���4�%(�;����K>�#�ٟ�>�O��Q��C�ϰ�x m��a&"OJ$R%W�&��� �(
+���1��4���Oz�'/�*d�6!�aԣM&^p`3ah�N)1���O�D�O&�d������?Q�OGfu�6��	����_#{���	BN _�&�ყ޺}_:�*�)��VEџ��'@ےCv8{E� �$����(f�j�X2�
�G)R��+Ȳl�6G�9]Ba���A��)��$�1H��������tӸ��"��T )l`H�k�Ip��D��yr�M�5�ЧU;���C%�N6�'N66m�Ol��:@�Q�l�I�@ �Ѷ�R(^�����f8ڶ���ݟ�PDl�ܟt�I�|J4)��`���]��d�3�4�⡸ �Y�lEL���m� �:O┒�*��~�,u &"Ĵ\f�7�k���B�ΰ6�:�25�R�j��x�+E��?)���?��F�RD��G�3" �D�`n�{���R,O���!�)§R`N�A��r�J��b��z��h��-��FO�z|�aA�'ӓF;�U��P
�y�P�h`r�=�M����?�)��	���O~��b��Pq�t�i�l`�A��?�o�-A��1y�ģ�	؋Vm*�ʧH\�@p��ٺ�IXM����O���6����Q�O�#}Z�Ɇ\���؆�O�X;���'�E���T����� ,�τ/��i���:vZ8��"O�IRF�,/j 0�ǔAgP,�#�'�"=��'��% x@�+%9����w F$}��'���'A�f �_A��'��y'*�$k�R����>>��)��<v�^��T�KR0�C���) :�5�iW	)t�pb�'m�YJ���'Nk���#�V�D�$ �� ��ͫW �,SBT�"�i�q����I��yr`��%n
<�'�ݕv~�����C
;��O��Ɂ�����t�2\֡������@�{갆ȓ5?��أ
��7�ҝ"�oʤ ���'�H"=ͧ��O����d�(kA��.��r��:M��9D�ѫ�?I��?Q��)B��O����O0��Q#ΛK�|�C�G^������Bݻ9m���
�'7,ak�ȗ%��<��c���6���#��@�2KP����ǆĒG��4k4��A��	%����ΰ3��$K(��Kd;c!�Oo�#�M����$�O��X*�K�9$Q�4`B�W�Vѩ���@��
4�	g�IO�I#~<�Y�T�B�H0N�׈�'4t�9���������M������ �xv�0l�\�I�v*�5�UMR��6��Ԭҕ{�ڽ�IǟdC&�BΟt���|��_��$� )SN� -�05�"� 1�Iӓ;O:أ��$58R���Q�8�$p�M�7&��x��?iM>IÁX#G?�т�C9�����u�<�$� )1NַA3f��(Jo<	D�i,��!rEO�B�j��ׄ/f�h�y2m�g�6M�O"���|jԎ���?���
	.T��A'�"�ȰhV�D$�?���&l��M�Q�p�g�	�y*���':s�p�W�W@W@8+6p��O
<aj�(��qV��n��>u*r��/�Ԙ�'hf�����:}���?q�����'�P��F�}�����K�p�:��<����<!t�w���6��	P����M@�lC���
':���K�]=�X�ʁ�	��Tl�Ɵ4�������L��[xT@��џ��	��(�\�a��'gT���C�&j�� ��M�&��X�b��" :ꥣv��[�'7]�j�*�h�
ٛ<��I(*��z��1�E��L�H=�aO�&�N���\z��e��]>�R�гGl�nŬ��ТҢ�+_.��=Y\��-?�/����>���O^�D��c���єOI�X ��m��hC��"s�6��$!�.��!�4�B�"�Sڟ��' �x�m�9��H��l������A	��'ib�'.�Mg����؟Χo+����{�f\�.��}r�5��Ć�ni%��n��P�����M���qa�NN>$�un��0���8V�C:%E)��a��O��@�T+8l�QD�}n���"o_6W'�ɀvlۨx]�-"�
 Q��$�L؟�(�-�(0�hH*6(H�$r4a��>D�dp��?:���f�&�@���1�I��M�I>y �O�B����'\�a�F�� b2@�)c�L�r�%KCW��'?5[��'Tr3�l���Q�e��4sG�wYh��^'HզP� (>+�mBg���p<��O��4��Б����`w,�����@��IB��S��"'�(��Й�4	:H=�%�Nܓ����I���r�N(�T)֛7X!:�L."�P�ȓv+0-�� �/�� �U�'O����	ԛ���E�� �6j�$I>�dt"U��'�.8�u�&�$�O˧l,���<�N4��E�6��q�@�9z,���?���W
�)��"�4 �N�����i�|!`̌
r�x�iM�{��	* i���
�bu*e/ĦiO��ǅ�( �=�SHX�x��躞O�B��><��j ���&g֙�L�8����O�'��?����=4����^�5R:�#�2D�4��˦Vs���S��l����j0O�HEz�.�/n��:!G��Z��-�"D^�p6��Od���O�QR-]�h1����O��D�O��M~�́eZ�����C"�1\�`p�RQ1J�B,�V�����-�}�
m�<��k�8X{p���E�;'"���J}�Pʆ 
�X��B�D��]���OC��lÒ�y���N�4�H���d��uO΋Op*6�fyRO.�?�'�J�臧*�
��FH�� I�A>�y��Zn�������Y�U;R�@���$^t�'r6��O�˓u�$ݨwL��wj�p��E�,���[3��`��q���?����?�g����d�O���J8m�ת��@�H�	���j��ؑ�߆O�
ݙ'lYD��p�WJ�5y�luiri��J����w
ű��]�����8���	�I��@R�o�?1�^�a�Ȉ]�[�h�O����ɠ(F.�:f+pe�k�@� ,��C�	�t!\����_�!6� ��>� c����}�#[%6��7��O��D��aDZ�.�Șa����Y����Oz�˨CDN���O��ӻI�x�ZG&��o����1@F�� ��s6��Ӱ�	Z2��3��,O@e�HÍsI�IX���� ��ӥ4�Ls1&��h[$	��cÊ:^���>i����V���j���	���J�#�M�0�bh*tܭ"sJ���S�? f��
�=Z���FS��XA6O��l�G�l�E�*~�S.�$~�$�<*v�N��M����?y+���{"K�O
�P"Q0��쭨O��8��Ƃ��?I��$<�ۧ�L�/��[���CF*�nʧ3V}�2�+:c�`�%*i���OHؠg%J�}p �2�f�s}+���|\dC��h�t�E��d4TE�6D���EKB���I�o���$�D�)�C�\�'n�b���0�D�=�0C��84�JW�Ȋe������,q����E�'r&�rsl��L�4���$U~����Grӊ���O����#���06f�O����O��4�q�`�1P��}�ac�XP�{5,�n�z&n��(W�e���ٶv��c>��N���C�ta�!��N�^�� �\b\.���&-[���-�(�5Fd���)�`J| 9�wM��R�@�}�#T�$A���hRJx��l����`I���>˓�?y�c�!��+�ƅUƨ���ǒ��xr�Ҁh���3,�|x�B������[�'�"��w�'��;FF��I�䍄�a 0��!�+�7tv�4!f�OZ�D�O��Һ����?�O�i���9�t��!_�?�&� G�Y�8��;�OC�+�2Ų�K=,O��P��Y>7�M`B�Y�0�p�ǃ+V�z-�/[�4v�1�W� c���"'�p�Ј{�쑓`Ob\C �HA��Up���&e�d*�v!a�%�&:�8C�o��pS��y����y�D�T�:�3��h"l�D+O��'���Rm�ɓ]uhmCڴ�?q�`R�,B�-O��@�A� %q<�y��?	Q�M��?y�����(��)Q�|�>E�d��E����fĲ M�w�B�㉏EOԬY1�)������(�j��̠f!�`��3_����FO��]��L�>/^^��c^v�y�p�mZޟ|R��3K��0�7�@W�:%A�Jvy�' �O>��#FU�m� ��\ʌ�b�Ҋ9�!��]���W���ڲ�$8(؊���՟ԗ'��q��
VvQ��'��	�i��-�|�	vlO�O0��g���g�j���ǟcF$�N�bMԌ��� T˂���i�|2�,��VUj�����)�g�H�D�R�Y0PH�	!rB�#ш�1�U^wD�͉�C����))d�p
ՄZ&1��+�(6��ɵMb����ܦ�)H|�L~��B]���*�g�B�$3VGDA��2۴��<�j�27�xY��D{c~���a�w�D"���)H��x���UH�U�gܔoZ����	ܟ�0�8�P�	ܟ��ȟ������Z񏚋}8P)IE��(x$�[�EG5'�z�$Xw��3���f�g�ɲt���@��:ce�Gb�0;�J6��k�1� a�*[/Α����/D���O����f��;Ɨ>|����B��4�c���'��4��S�g���69���V� �¨"L���B�	�zA�%S�ڮ-���a��B���"̑���o�ɉzQ[1䉛��9��|n�9��)��w(����̟p����HSYwd��'|�Z�r�ҥ��,�X�P��dH�67X�!�/]�m��-��,��z����ĕ�[b���U'�)�W`���r5�ȕ B\��5'Z�wi�1@�LY.q����bɷf`��L>��b��"up�@$��0U�p+[|R��IŰ?�@KW�Y(H�d��b��ѳ�E�<A�C�e��D;]�Z�R�lEe̓"L���|b�
DM�6-�Ox�
:+7��h�m�M�� C&*�w����O����-�O��d`>�kùN�.�B'oŃ �<����@g�z�A�L̾`pF�	�{f��F o
豃��=�1,�b���B��H� T87���L��i�d�	*���x�I�^4�r��G�f~� 8 n͛W�B�4o��k$�V:���A1E���B�I��MceiTm�������d����L̓!����ѱi�R�'���l4~��I-`�Ȁ�oT�[���`2�״r�2���ԟ��V&���*6N�*|� �S�$]>	�C��/�<�3g*$W�R�8(#}*Y/z�r���4���ӂ\�F�Hg,��`�^uڦ.�� h�'Ʈ����\ɧ�O�*�kDȄJ�$���C!v���yr�;�>er#�؂S���Y�̛��0<��	 ��3�Z��!Q_�N���	�O��$�O�pc�(0���$�O���O�H�k����d��?g��
a�P��V��7��� `'!D�%Zs�(�~≚h�HUG5A��0a�oŵ%U����șc0R�m�M���:�<���� <t�!Y�$	?{Xl<��T�.0����4|��ɝq���4����>��-kp��B�O�4���7#w��B�	+l>���h�8}��	1��Ҋ~[�����'���Ɇ$�<RE�A� y�MW�M,���sK�=J��O"��O�8���?i�����C��n��!�-O��``"Iը0�h�)dZɻ�ˍ*g����I7\}�����//$PB�DF#V�P���]�����f��VmʀP��'�p)[�,�	2T�fį7�N{���,�?���iWn6--�I���O[(�X"J.g8I���U������� �h��f�A�F1�l�6_{�V�ZM}"Q��s�ȓ���d�O�h��/W-;�ZxjQm}W�����OR�$��!�n�d�O0擹
��Hx�/�mv  �N��u��鉴'H�	�b�RF�Њ�'O8ı���!=����J�(sh7m� 4���a (�~��&
�j��xb���?����$�q�(dk`cQ��i�U�@/Y�1O���!<OĘ��!䎙�N��*��3�O�9o�6��y�RnG�P�@Y�C���0�oyr.ߜ F6m�O*�ġ|�pnU�?1��Ŧ;L�4�B��
��ɂv��H`���?Y2IO�2�2��ND���T>��Oh%j@��&��c��#� sO� �@V�lc(�Ph/�����r��[�L��B&�=$�I�O�X���'�J�O� �Jq�12���@R�L�Դ�&"O9�Q�'�0أ����W��<���'P�"=A��m'��9��F��ੵ���	ӟ8���Y�� �����(��ޟ�i��3 I�(�>�!�R2Քѫw��$0���ѩ�&.�6��M�v���L>�f�G� ��y�b旹c�X������Y@8|BQ�/
�7��3*����L>���U�_D�,s��	3Z�H�#׫݉�6��<)vb^���S�?��?�uH[�@�m@�gW�nT���VJ�<����av��p���m1}ӥg�C~c2�gs�IvyR@��\A˓ �� �yL A��"�B!r�'5��'�֝ʟt�I�|��O�1n���P��o<�r���3y9܉���MwDI�#!��"����v#��Y����ơ�}<�c!���D��h
�vǠ��K�)`�I���?1 �.(`r��$�L3|=�b��^i�<a' �YW���g���B�D* ���<	��$ێ*?�n�ҟ��I;=�Xl(�GM;N(<%�شK�ri����U"�d���|1�@�YW2&����Hj���@��.E�Z�c��7O&}C$�bܓ�̱"��E�5�ħ�#y%B���	PdT�D@_�	�7�BȰ��6Hz�7���B䉇$����$ȃC��sp����B�I8�M���M�g��$Kf��a��r4MAU̓F��C$�i���'��,a����f��m�fꄳ_Q�%�Zh�$����xÇ&�]�%� W�=�S��R>W��	ld9QG,in:Z4f��I�o�tH�nH�>2���#�'xT��b��[���R7�(�O �E�'1O�^�C@��<��}J�Է[��A"OX�$e��N�<�6@gr9��'d#=!�AEx7x�#̓Z"҅��e�6�6�'���'8b���U4���'���y��R:YXp���>-��\�Q�Wn*��a��<���@�e�|&����O�-�0�S@_�%rM2�Mjܰ�`)Ot0G������9d���4�=�t�35_�)I���?��Pa����S�gy��'jH�i�a��)��!�ǐ+IδS�OF��,�?o2�����7�>Ѻ������d\��~2Q��y7��x�u��baB�G�^�G�F�[e��ǟ�	ן��	3�uG�'��3���{V�Z�17N�`� ��
l�)���l�!����x�;�P�]�@����=UP��Ov�;g�7/(��d��*	�Z]�aO��S�ҥ"�OZ��w� :{�vtj��h$�1ce"OL�keIV�e�����W	��"��d�L�D��	*!�iC"�'m\�����>g�v@;�̅�yJ����'����.u��':�i%Q��m�+�K@B�33���V.,7/La�t�ޣI�m��(+��0tK߽B���bB�S%45��@��?aƠ��Bc�� �._�1y~">ɳ'�ٟ��H<��o��g���zT��m����0e�`�<�aH��
u)$E�H�Eu�U<)��i��R�*�z��a���2��1�y����7��O��ı|��h��?�� &:<6$a�8�b���mG�?��nXUɐ/R�\��6�Ϗ~p8d1��~�.���q��B$b�0XA����,�H%�>� O���)RL �5��)���O�2E�6��
z2H �dؖ)����L�h�@ �O`�mڂ�ħ��YĚQ��`��+�
���%2�@�<�����<	Vŀ�mR��� �G�Qt��t��h���9vtB0��,��w��y��/>�L�o�ɟ��������r����Ο�������݁|?z`�ڣMC;qeR�L� ��$�i�h�;�O�W�����2��O`J�'�J�o��� ����B����w)Y�Q�z(�l�7��L�l��ظOl��-O<�脠�8XƙQVo"M6�r��ʦ��(Oa�A����?A���?��:EDX:��8Y�Q�S	��x���8qp#W9n�bi;��T���Q�'�Zy
� ���t.�7l���s��ސj	6�j0g���V���n�Op���O�����{���?q�O霸�CL�$m�f�@�K��r�0`b
Д��RdLJ�F��Qc�	%,Oԙ9V̓�q0ށ*�KJ� ���ѷ��75���fP�(ޤ�z1-�}2����	��� bBCJ5~��j��d��)�T��O$(o�ē�?y���'.n����$� m�cF�T*1��'��=� �?xla��,�P�����yBƽ>�.O����I���m�I��h��H�4,4,YC�l��B=<-ʆGʟ���V���I�� ͧ[�9j�#vX䕗'bv��H����g��7��m�ǓZSȜ�g���b����' ԁ����P}p��x�!�=B��Ij�ɀj,YX媇�~��@'A"�C�I=
� `�gG<*�Ay���&V<�B����M�!�
o���a��13��h�⡜d̓Va�8��i?��'y�Ӛm�>��I`�^��"B�T>a�5.�0J�����$P�c�_�Ұ�w��Y����a���i�|�Ph�����swL� sx,�'�r�P�w��8Y�C6La�Bec�O%�����Ҡ3������o r��J��SE)�O�c��?���'&��m�F���{�`��7�-D��Ð	�?�4P2��δQ��A�M/OdGz��V41�r�X�aݰ:5�UC�(P�j7��OR�D�O��2&�T]oh���O����O�.�U����U�'o|u0g�Ad�0��h� ��'ZiP��T7����=+�IPe��
�ԙBi$X<��r�Sa2��H
����c�%�uܧi��L�����=q>Dٴ�G9t��Q{є|�LG9�?�}&���O�	u~�m
�PD�8D��j@�F2J�ɛ�.�X��y�`;?i��)�'y��ܢ&K�VbZ���Ԋ+�p̄�g��؄�Ɏd�L�C��	���ȓi�4���P  ��lã
�']�
��ȓtj�; %X54!+T)X�.MT�ȓZ���T抩�hl�f�Y�"����ȓK����eE E*J�r��W�%����ȓ]�h�hL�?Kpa�@h. �4��ȓ[���+"k�p�A2���Znȇȓyz���U�ޞB���$AU(yμȆȓRyl����=6x���ۡac��ȓ5}���g#�;%�mb� j��D�ȓx���Q�mӂh�4!�J�g����-�fy�E�ʅK�m�TF�D�潄ȓDLH� QǑ�'iR�He(ȢlB"���x�9hĮ��y��[tǕ�_�ȓ4݂�p'���(4H�%�
Dd���-�.�q��ғA{nu��F��^9N���wö�r�*�>n�Υ�EoV�����sP�Yc��ͯ=�NL���H�3����ȓV�� �� �'�0����4K��ȓ1]`�q�2PH�c��Ħ�F܄ȓ2^�`Vf�ct�$�$��D�ȓ���7�\�d �	���cu*��^z��q��Y�0��Pk�f&⑄ȓb�!���&|K&$s&Q^ܜ�� M�D��	����L� ��?��S+d�Q�wo�  0氅�g& 8K*z��i$Ɓ��Ɇ�G-�P�gdQ�T��S��N/�@�ȓpBe�$M��C�rx{3K��V����g��d����.�6�Z���x*���}��ET�ϵ6}�4���[!�^��ȓ	}̑���O_��[C
Q'wԅȓ$�B�{aa�$6@��Y<L��ȓ?+"���\W�n���bq�͇�Q��
RH�L�P�K���#��Ox�� �j�F%R#B�
H��įWi�1&�Q=���ҮH�rW�C䉐hҼ�P��Q��� �-�ɔ�"�[He����`[�@��D9�n��R�̼�4�I�Q�pb"���E��C��8������2�SɀPվ��g�~0�y�"�%��
Q�yx���C�:l����smشJFu��*O�`1�/ξ+C�T�4���N��M��� p8a����K3��k·���u74�t�DΌ�`��@�e�Sh2���#2?���H�HPd9(�W�nȘsD�4��O�I��H�qL�L@�aU�?����'yt Eۥ0b�p�ȓ5(�ظ�O�4�\�)�/w�<X����9��O�'���P� I6y"�8ò)(]T�A
�'
��R�MH�a��03�!Q0[�E0f��9R��[R�S���fH$#��y����a�T]�G�m�
�0<����\��2�`�~��a����b�=�-�n���;oԶ�@m!
�'1f��I�1�ƽЗ�k���+�O^�y�'�a^���S,֌\�0;&�%��Of�
�q�t pG��.u�5��dF�0Kp���'m�(2�h��ǀ{�qV��f��9n<(��4��uǪ�p~���~Zc�6�c�@�,0�y:BߌH�r�s	�'6�aF@̛g0n��oKar�ek�-ҳ?�Ľ{��G3��I�'��IS��|��.Y�U1$I��
9���EcU���%A�085nq��WZ��a��T�@� <����]\6���S�'�:���c8�p�0�"%���T�w��(0������a�+�$	l�a+�O����*G	��m�ҠS���1�+���@��@uGX�L�L���QV^5�
P���XxS��G>�@�S/ã}��O�����6�|�@�!��f�{��Q�=�^�kg��/d��ڥ`�j�nN�S�ʹ�udb[w��7MH�V�:��W��-w�p�N�h��Uj���8%\�p��0<O�Ŭv{��q�NT�q��A�=h�X�h��I�<)��\ &,؁R�s��IH($v�Hz��Q?_�僄ޙi�ax�O«���� dp�M�",2{�I*4�P7�h�(3h��qCs������q�|�Æ(5�~�O��1F� T�]��N
P�E)X��HA�ȸ[���0⌓���17����X�@�~�*I?����p��91��AO���v[LA)EƟT�D<�8��fZ	r~�9��(�G�O�y�p�H4�������=��E�M�eQ��J����kN��N�cQ��M���禍��6���FH�`|0�abДkc�8���I�+�	������ʛz�r@i�L�H �R�@�a�����&�R��&�R* J���D�F��?�ȝ%G�Y3��єi�ޕ���!lOz<�6�Ǚ��"6�����	�.�kZ���IH:Zd����PhBX��=O���#E�c?��4��lP���4] ����̼��B��kvXa �K�~^�OA�֦��^�$2��
*��So5�6-NQe0�ItJ-���Qb��{��TQ�6Od�@`K>eVH��$_5�0�Kp�I���1�e�ݓ$=��+�cK�*e������<K�˙Y?�R���a�iǂ�2f�ԯ]�,�s
be��J�2\����@��l��(F/T(�q�'����lK̼S ����Q���D5;rhTʀ��(E�-�E�7���G�N�����qm���O轘�=?�v���L��XY��$�?k��y5�:�� ��չz�B��60O$	 nZ'q ��2-_�p�zxI��A�@b�t�Y!.S��\�E���mJ�Li� p��M���r��F�ʵ�˘(��JՌ]=l�}e�M�����v�P���~��8��h�hQ9C <�C'+�)A"��� �O� �	�L���$�4���,���w���}�J��e��5+P�¦ 	�yx�	C�t�[���E�$ �<��}x&M:X�P���T�R�2��4#ɧW�ҥE�ƾ1Z(��b��F���uz��G-A�5�$��LO� 4�xZ#��~����%�������|2OI+t���`Ƈ��%�C�r�'�r	[���`\��ɜ/#�h �,��!��(k�`ޑ7obY�1BXJ��)��<�{�.��Z��D�H��O�(,���N0bpX=�	�[�U@�i�|f��1�N�AR*��q�O'`��b�o֪_�������TB�a�-�y�O�QK�����ߜM����&��D�5�mXB'�7��:Ԡ���ў�B��@QtHc����˗	R:����DYTゕ��~�1����R8W,\T�\?���X�x20��,[�[�v�{UK0���s)XKџ����EH0Ur^c|A���Q�>��M hR	[�a�O"�d� JA�f�@�ԟ~�	?�*h�K�8�����E+�ޗ�L����a$Ւ!C>�zq���*o�DS/.<B!ڊl(�u:�N`q������T��	�B@���ѯ�ş@Y��gq���OܟRp^Q��Խ>�\��\ `��k��7=`H����	��D̿�^P�O>�g\�T��P�Y~��ቶt�@Qr�-[ş�X�헡H��hI3$Fx�n��+���{Q�3GJ�a���41o6���'��3$�=}rE��1���#b@�L4��$W&(����őF\�у$m�*�rHpa��H�^GB��a�����t�Q��oS�d�	ya.�vzl�p�J�<1#앙���1�
��)��4J��l�E��P���$������ቇ�^mɦN[
*i�i����M̓)��I	�m��hQȝ���L4��[ `�s�!p�$�A_�D#sF���O���ף�=P�飣�'!�D{�B� <�������z�Lql��(/�W=���a���:�X1˃E5?4���^}�l�	!��|�P�G��ϲg'�ޟ��̟�L���;#�:IʔX7O����˔m�@牦Hq�T�P��O���c|:h��$ߟe?�P��W��<|XEN�J���6j R�h����O+�h�IY��5v+�HX�qϜ1Wz}3׆A��?IM<�b��>��ɯ;f�o7"�J+_��,9�5E¿(�����a[�O:m�F�^�.Xpbc��?Q��)��Є"B>�y*��]$���тJ.�"˓6p���?E�#���4���{�P�3� y-�WT������V��!��QQ�qyA��y� 9;�4\8"�Xc*O�!��ئv#:@I�ˈN4���'��lh3��T?������#��Ol\*>2�@��C��X���օb�p�")O��"�4��'�(�2�3O�F��F�\i`S�ϝK,a��%V�#��ր�M����w����ňp�-��!;�K5U�xX�F�
id�����#��U%��	$���<��>O��;��X9g�@��g�	�0�ʗ�\|�"<Q����h��M�����?	d��9��ϓ �P\�LĄffv1{���>!R]	T��<i�4&�6���?]�DԤ�v���~�R�>v�4śU� I�N/W� $(�0Z��(@��/g�P�"����O$|81���'��Q�0��:�8���8p��j��J�J6M�6g����'-���O�`8��� ێY*&n�$�,�pC�S
�| �鐅"bmB���O�^�ֽ��X4���m�/H�e�(b�HJ/9����%�O�����/������+��t82��:l�MW�K�A��\�<�ܴi`���KW�4��e����� W�����)C�&;݂ͻg�I�7Th��ű?���I,h���s�H�?���k�>+/���B��$9�����v�����mDH��⌜]�`��㞤�T0qÄ8	w�@x�T����F�p��$P�D��ǎ�Γll�	�$���P��<y޶�j��@�r�j)@p��qnZ̑�e�F�%+��'ݠa3�#�(�%O�H�pdb�'����7��=:����R��ȃ�< ���*�*\t���D*Z�Q���m5��P��I]���~hH]%Ca�x�� �8"	����7�@�yaǀ�"����\�����+{��kF1A�O���Zw�1��T��x"��4 "<���4U}~-Qeȁ����%ۓnS�)�FN�
�8�
���nΰ<�2�2-4qO���FpX�(�y'�U�:�:���9kHY���+��d�u��	�Θ��Z�"}bdM�L�d��cT�_$5Br�ӛf�h�P�Z�|�� م�t��J�
���,5ʓr��Y� A�Dт�s �5h]T�ΓZ��eH!g2jP��'D���$S�Hh9�U��n*f���4=e )!�/>�|��b��(=�a�W�2Bz2!���7�I�0�ԏ%�)�1H�+0k�ܘ��kJu8f�R�����_T�]�T��c�� ��u�~m�Ņ��~�Oֲ))�%ővp�)�Ɯ=]gĄ��䔨P�,dPT�S�C-��?1�d�ωb-��I�k��w�\���	���*Ҫ�$0�h;��Ĉ%���s�I�C+ց��g��:� �$Zt�� �f^8��h� I�G#ƶ3~�%�*Ț� a�!��L{�'y>QC�l(/8�- o�9U����򄅅{y�Ґ������QoK5HH�$Vm��J��56�ɝ|1�i��@�o0�����
d�,����Q3+@R�i��ʪ~��;���Q��,D�F:��D}b&��s�:9#�X!/,�X:���1$�Ƒ��oN�sh;��O� �2�\�?�}�'H�)�,�`�	0)k�ո��O��PC��D���.:�������f�R�LF���&��q��B�>�)&D�2���v�
�T��* �S�b�B5+ǣ[3jO�P��O�S�"\�Q����y�"��̣�hˡ$��}U�ۑ'�|r��*�HvS���'��dɷ�M;���.�Z�� �[~��#w!M,U[n9���E�= ��N�<d.���b�C��1*�# ?�EyB
�u�s�F��`=�� �(O�BE'�M�R�U� R�'0(q2ef٤d��m�k�7G�������l�Ɇ9#?9���n6�r3l�	<��D�K���؈u)۟���G ^�+1�6���>E�R�\ˡK�<���yW�Я��Hb�#�z�5xF�9�0?	�͌�b~�Z��FZԒaI���2��A!q�ϕ���.X2��ϓ:_����$�����\7�X}��m�[�z�p�I�xP�W�C�(��I�W�.��4�!O���(u��!e@�6M�'K�#!k�|���HG��8$10D2��(�ͬ4�z���Q2C�� a�c:�:nlBv�7-�]O@�!n�}�$��}�����?�N�M�nml�+vJ�� /����>@p���ϱ�))h��
 �p���ߑ�p>quBٝ!�T��d��C�b�[0�I���;�]%��d�,f�ў��;5iԠ�ta��-�J��
���\B�d� D�!n����L�pl���!�YV�'�8r�˃�<$�);!s�Nܷg6>�R,�)�x�	C@X�|�e�L� `�剭y���cSd͛$���3u�Q��vx�'8��Ĺ�"���e�mo�[��N2#�T,i&��:�h�Jt�$2��ˠjYm�@�F�� $��XG4Dh$�
�:��-a�c$b:��qLS�r����d,�OB�P��Q&�y3�d�~�\�"wW��
�ŀ�)��pq�̽���S\b��oF�AE*!��"3dMr��ȓp�F��6lc�dk��N$;t�,�ȓ_�.]�A�_�yIb��Ve����e� �qch��5���Ơ�i����ȓhn$�0ܐ&xH1jV�ڗOa`І�V_�����T�$� JSD�ܸ�ȓ?���(p�H-i�X/�.b@��	Y���e��q�n�[�jމwB���ot"�1KΎ-���f���A���ȓd&������Wp>�ȖƐ� I��S�? *��1G��K���r�+<<�Ԁ�"O��bF,g�\�I �M$.Z8Q#"O��"gФ:����<!��CS"O �iW6T��@hA6B�"Oz�(�	>
.�Ѷ�Ԓ<p8�"O�4R�ƍ�w#a��
L P��Q��"O�����!EL��f�]��  g"Oj|��gHS���"pn4�v�0"OB
u�ǫW� )5��� �D[�"O�qQѩI�B�^�`B�� U7�-��"O�A{�a�)j-�m�D�Y�@"O�xvk�6p����_3Dn����"O��i�o̢_�,�A�J��G�(�$"O4Q�7f�8Aڀ�⌡I�<Ų""O�58��:�
H�b�0;�|D�v"O�$���K��b�Kb�>Q��$�6"O��b���$K��@��r� ���"OB���:7�� b� �a�|5ڶ"O|i��f��J��H��2#�I S"Ofl�"��
�5h)����e"O\	!�R�C��ċD�=��5XW"Oh�!�L�lA�eb�Q���}��"OP��'��{�������\�\u"O�峅b�|�N������ �ʽr�"O�D*N�Q�0�p�a�2ю9SQ"Op��J=p�4yAQ �7,~�@�"O"٫�F�Ys����`%}��4"O�����@<�H�@�.x|���@"O�m�ӣ�+F?V�����i�5�!"OD�A��ϻE��KĎ�6�"�"O��6��9Hp���EN�\oF���"O��ZB��5v{BJ�̓�Q��� "OrU�QHG�A
>�
���6՜!��"O����������űB��Ջ�"O���S��x���ԴqX`����.D�C�i��`�b��I$-Xu*)D�LS2�ý>����e��%8j�+a�%D��JU9��P�C=P��hzR*$D��K���sњ|H��K(��i@)$D� �b��s@��'b�y�x� %"D��2D�K�Yhp�f�H���� %D���Q.�%$��!�!�p�B�KӅ=D�X�N	:{������ͪ()���(D��K2,
�;�"c�^꽲��!D��q��Iu�uk�J�> ٴ9#P�5D�l��C�Z���a��aA��� D�8kSd(Z�����Gr��,Q��?D���w H�H7��A�(�-"=��!M>D�,S�D�) h��Ǆ�d�%�9D����9y��S%��$�	�	<D�@�����,��!2'� ��4��->D�iu@�0&�����!X���V�:D�,;���	/PI��.jDf�;D�Т"�G�)�8A-Y�OD�2�c;D���lA:l����$حmp.�
C�%D��Ӑ�ǘLBuK�
:����'#D���UN[�:\r`���3X��8H�H4D��Ke�U"���N+d:����<D�$h�ܞ7BIY�� '�b��u�;D�P��I��j��@C�H�2�J8D��0G�T�|d�b�[�I�u��2D�lBt�L;,ڤS��3¨�P�<D��2�m��uӤ��� ݎ¢T�i;D��S��b~��@�^tx|4 �h,D�� ���E(Ť}/��B�.��\5�9�A"Of �էC4�\�&��/+�Lu� "OrSv�@<wՔ�h��̳B��P
�����	�4����7�Ŧ7�}Pǧ+݌C�	�hTL[Ǩ��,���Q� �p��B�I�Ov��p��Nd�!ba��	qlB�	=k2ia�V�R�킄,R��VB�	!#Y���G	`
@�K�m��PB䉩09������|Y��S+Z�b��C�Ɋb�� pW�ǌYP�mU��
=��C䉢gV�:v ��yČ,k1&��tC�	iJ�Y� �X&>g\H��%�B�I.Xw|��ʄn�
8(C�V�PB�%!�2� T!O�F�zbLZ�Rr�B�	 hv�ĐB��>p�a�"�C�F��m�'(W8� ) �#s,B�I�^����G!��0���i���B�	�y���d��./����7(7H�C�	<�r�GÑ��(�;�Jî
��C�	��X)2�5n�\aE�R$�B�I	 �44褧�%c������:ʸB��l$VL1���"����/�<"����d<�I2{C��cs��2��<�d���h��C�I.��1�T�%���Nܝ#�<C��+B�(��i0;���񩟖A�4C�	�|Y�|&�6pa��h�h�&t�n�'�ў�?���!��2)�Y�cI�c��y[��1D��E�5A�`�`q��J�IRA<D�̛q�:Kb) ���*�g(�>��������Y��l*�9��h��W6�*�fK"b!�D[�	i*T�(��f4�8���h��-�OX|�!u��v��(n	.��'ڛV��C?�ŃL�@F��UФx�<P,�n\��1�������D@<�p�e�C�6U��I��!uDs*�A��g^����ȓ�����;"� ��`�Ȼ�H���4�O?�I&���,���A�K�~ʓ�0?5�^(.�Լ�I�;j�����N�<ir��>s�
�iJJ�G� ;%�GG(<۴om�m�)�LJ��᝵����ȓv��j��E7O�ޝJ�,զ'ޤU��n�� q�+�#A����У�.y�L��J(<)����
�t+��M�xS+4�O�OF�b�(�lu6��Bi��� Q3"Op�SEIHm���i�J3fk�d�g�x�y���O{�9٥H_7]�T�bB)ۡ'm�8H	�'�����(�%j;Ѐ���Ǔ&���!�4��-+���S�3�dӲV鈗�3�R����]���Y���O,�q�C��>�B���N�  ZKa"O­�t,O�9�
�zC��R841��"O�h�gC:��ț2�R�J#.�)'"O��`��F��qg,R9VH ��"OX�����N���!U&�=[��¶"O�I���خf/@ؑ�do�]ZB"O�,@�_<�A4*�$`-"On����
E&�3�/H,/�����"Oޜ8�!7m΍P%�Х3�Pl�e"OT��ra^)aβM��n�%�4��"OF��� #*4J��^�>�KQ"Oz�pF	�2	�.�Y�L����["OX��c��0��� F��N$@`"O��A���H�����M"�<с "O�Myf��=e�RTja��t=�%`$"O.����$.��H�&�2O�8�H`�'g�� x,���9r�N5a��9�2�rT"OJ�c&��$<��r�OC�<L"�"O2����ȵm	7%�Q����"O
�S�U�U[2� �1�VL����?lO���/�y��<�� ߀�Z8K"O�1*iX�/5~�8� �k�BP*t"O�x*�FY����A��&�"O���)A�n+ִ��O���x)3�"O�����75_R#un�Aa�m�E�O*�=%?M:�O`I�W�
>lg����"��� u"O��{�lؕ&Z�p�0N�1�����"OX��pJ �����U73����"O���-%���&��22��i�U��6lOV=iw��Ƽ��@�S�|䑶"O�)�.P%��R�' ��\��"O���%lT�,���˰w���Ad"O��3�/D�Lºы���>�V�i�"O`h�j{mvۣ.ڨg<�ْ"O��R'�KV]y�E�A�VY��"O�-IU
��^��(�H��V ��h"O�1*EfT>��ٳe�TL�Y��"O���K���p�
F��"Op�NN=j����
A��	�P"O����ʒ�)���riR'c�$P@w"O����� �^qP��05h$R`"O�x0�k�7y"�8xs�P?���#"O��� ���Z�i��'ю1�h��%"O8�� FT�Z�qf��%I���Xq"OZ�����|Ơ����,9���$"O�A�BJ�|�pز�C�,au(��"O����N�H䎵y󢊄Brz�k�"OZ���!
02�%�W1n�p§�|R�i;��>��PAT=\�r�鏯4�L�gN?D��Q*�&C�=9'DM&{�����>��y���c�iI0�b���n�`Ȃ0�?4�\�'Or�2aPKWiY�٪�y�<�u�G�tG�J�@�	��X�j�y��T�>�fE�.z���Ie�M��AT��v�<i�FWe J!�'j��Gbg�<�D+�;-�!ct""wE^�#�a�{�<A��	0@�L���Ý"s.�{1Ez�<�sI�̅�pʕxo�P3vA\z�<���&%�2�S��Z,�@@ÔD�~�<��C�7,w����J�Q�`��UNWc��hO�O3��U�B��0dL�H���2�'s,���ѩI ���ےC�,<�0�+�I�C�Q����;������z�vڮ�Ґ"O^&E
���*�,�=�@��c�'1��>}��'[\eA��'P�
�+]k��i��� �D�O��Dc�����%O�h�BM\��*�+D� ��+ y�
	+S���n�$����*���,��U��)��M������<qg"O`E�Cgי��P�ϕ�S�`�tb\��?�Ê+?��t�$�9O������J�	�Q��>�v�J�"Oޥ��˲-Af���DX�L��3��'�!���!r�FM#`Æ�U��A���
	!�D�V�������< ��ˍ�!�DV�@��e2G�δ<脬���[�!�$�+�����_�^�R��d���x�!�$�='h���sDD��I���B�#�!�dA6y�l�p'��Yy�X%W�a�!���Bq(���
u��[g홷�!�d�x� ����~o��C��{�!���o0ٓ`l��-��ų�v&!�� Pɡ1�*G|�d7���|�Ȃ"O�I��?P�*��P)�/(�~xh�"O��	��R*Ck~qC	V�ؚ4�"O�р l�>5����ځ
e��[�"O�i�t�F�ڱP��I��A`�"O,$�t��e�]�҂�������"OjU��f$�D�#�Ɠ
�ұ�"O�T 0A���� X�#C���"O��ZfA�L�Z	4��5&�(ň�"O�	�陭 ��a��	���Y��"O|[�1C���!�)w�PeK�"Ol�(D�cun�g�O�~����f"O��a�:;kv����A?@��@�@"O��Ӈʛ'�8����6LfM:�"O%P�� `����f�;h�qU"O�(�Fn�:2T%	�Ǥuy��"O�Icf@ʄBL�]ĉ� �U�t"O�HɅ�Z7`hx@x"b��w�6�f"O��f�ٍ�̄ʗ�ύ5�l�y�"OZ)� 8P2v�*�.W{ ���"O����LӽZ2�L;�٦T(��"O|m�t)U��,um�V
�q�7"O�Ha�F�?,B\*��?O	B̳u"O��+��J+azq�4�٤5��"O��`����ਤ�ݘB͞ �"O8TQb ہ9�0P��a��Dّ"O`�գ�""w~͹��	A��U��"O�=S� ��`	�����Qq�"O�лV)΋'k���B6-qA�"OV`��K�l���P�c�70RpD��"O��%�8})�1b�Q1,?B2"O$A	�:����a��};�4�"O!h��@298fb�-OS�L$"O0��+K1v<f�hׯ��gB�h�"O�*qG�4zfD�W-MĖt�P"O���mV�]��QbujS ��Y�"O^`��ݐ����FS�T�j	��"O��c�B���$�
�*Kn���"Oԑ���[�ɹ�lR���r�"O<��C���`��I
�KAQ^�@H�"O���H% tj�
�sT�T�'"O@�2�)L\d�$��k�'0�x��"O�Yr�D��.|B��ȏ.	.0i�"O�D����XE��hQ@�<��XG"O2�K���.@3`��,��ݛ"O4���L9]=j�DM
gx�h�"O�$Ӕ���eA$�Ӹ\VR�"O�z ǂ!A����h�%=,���"Of�B��b��4���3;3n�C�"O��r�GV�M��ՂG�&<��"O�$؂"�:�"-��L�(%t�a�"O�	�D	��=w��#ik��t"O�1:S�
Bjp,��X��d"O�H �Q�I�^Ep��πYW�tr"O�v�X���a���	M9s�"O�5�]'.Q�M�eLT-4]��"O`��T�m��lq�/r@��5"O��K���-Q(̈ ��	�"O���6�:Q20�U;A�x�`�"O���#��&.��+��L��|��"OP]IU���<���E+C��1x�"O�1+AoW�T�@���D#bX��"O����� ,�h�+ �4 �C"OHѻ�&fAPphP!D���cP"O� ����8<���򪊄 �|���"Oh�B��½��*�!zM.�0e"O40q��H���s)�?J�2�"O�-鵮�-;�d��r�S�p �MrB"O�!�⒝Q� !0g�F��M Wb,D�)�*�[����Ǫ�&�o$D�$�f$��i�p�ba*Q�e�@+� !D���A�(X �8)��\:w�E�qF=D��2E.���XE�׽z5���:D�8{�	gh�AT@لn:^43��7D�誶��	I�><Ө�f	�`� �*D�,�bT�y�*�:�LRb,�iq'.>D�t�GD;6=,%тN�Wԡ�d�>D�@�A�;�EX���&X&�K�O)D���3�F�E�TR3D��2��b��1D���Ǎ���|�!��/U�98�C0D�Tc/+6�1C���c60�/D�|8��\�
M
3��4�D�2�,T��6�r�C&"ώW_����"O~T��W�jff�0�&ݕT�xt�T"Op��&�Y9�v�Qq�U!^���
�"O=a�����e�B��5"O����-P�J��d�#p��"O�ȳ�U#O����oPx|ۓ"O$ݫ��/M�(p"��	;|2"O���ȕ�P+H�Ga�g$��S�"O�<���3@��֊L�C4�-�"O�$Z�A��tU��+ˇ�22Z�S"O1`���
+�IC����(�"OFm��K��>w�!����(q|,��"O��є�ę %x��0y�̝(�"O����!�\Aİ�C��+�|�в"O6��G�BV�mX��M��h"O0 �5D�B�(�Y"F�0B��["O�!7�����[Rd@.At �X�"O
0�CE<����C IǔT��"O�����-�Q�!,�]�"O"U�B��7x�֩Y��Q�O\H`"O�JԩϼYet���\rDl�`�"O�)���.e�z����}��9"O���C�K�DV
|��޻=
�$B�"O�I��Щ;Ӻ��̍�j(fu��"OzTb� N�L����L�!�d�r"O��&Āu�J�9A,!&��	X�"OP�B�U	j�-��{��"Ot�J"�"r� �WFJ?:��D"O�m�=Z�\+Ђ�'h�N���"O`4��Ƒ�k� a�J0f2�"Ot�񥊳^,���.Ot�"O�!����|qGM�(OL��ء"O�"�h�
N�L|�����P�T�"Oz�97��8>�<͚F*Ęa6��#"O<�5�� Q<�����o2���d"O>��F(̘T.����[�l)
��"O��� ��U��9btG��!4�A�"O����r��x�`K�,�c�"Op�y�ˈ�W���
�n�aHb"Ot��'��qs\�A�`�c1"O��8נHږ,��\��ҘZ�"O�#�`9�<�,Һ,�:��c"O���S�7-��z,!j��J"O��r��G#P��#扚*���"O�q��&,���b�R�*9��"O��q�C[�;z��b�N�31lMy"O� 84c*M5$���pF.@5n+v�a�"O0�2����I��n��+F��C"OL訦MJ.���q��ˇ҈�`"O~AH�KM��i��&,^#�p��"O�@��C1V��X�G��66���"Or=+����d�R'-��4�#s"O��Ku��QY��w�6�%HH,�y��5;F�"e��M�M�Fd��y�Jȱ6�b!i�DCOJLc�lQ�yRO��H1%	h���P!�yD\�W?���V�e���b�c�yR����D����c�Pɑk��Py�E-7#�XZw��S�����d�<A�+�"nj@u���c���`uLb�<��.
	�=i0�U�\�<�e�(\;
|dL�E� �XQ�W�<9'��-�T��U5R�P��O�<���8@4� !琐\�P��Uv�<�c��F� #�)�#^Wr9j�	�x�<ї� �x�"5��*Qb6�$�tf�p�<�2�<
�t��#�\�
q��!2�t�<��E�����'�M�X��đ��V�<	��:Y(��[W������[K�<لH̛X�F̠C�0�H��U�K�<�ׂ_�}z>�Y7��<a}8��Ĉ�J�<�b�-M]>�9�ߠZ@H��g�H�<q�)F>�`3��"���GI�F�<)r�C3�9�#�P�<��ö*_{�<f$!"��3�mRE�8�P�s�<�DL�=�� �@�ZX�	�0%$D�����Y4����4,���B"D����mȪv_J푠�'=v�M{�I2D�S� �S?��Z$�[�X�T��"�.D��g�Ԁ6w�(�ׇ��B�<���)D�P��銊V���!`�u��躡�5D�X�  �!F��˳͉�Àq��.D�D��2Z	��3*F@�r
�**D�8��l��<�X���=r�ɂ,D��SA�RY��I�$L×4��k(D�L��ڵ0�\�w���8����Gb9D�D���/�s7!_>yn����:D����eɈ8�N)�1/�+>����P&:D��p��M"$L.�*<&��*%*#D�#�Re�CW,$�v�Ҧ("D�$؀��;|��"��ӱ0q ��!D���3�ZL�d��*����5D�dk�Ì�Q�eB�J�v��Vk2D�L�RO�$ D��#�w�^D�B/<D�\@.܈%�\��զG���Ue/D��毙�Y=rE���k���ɐn,D��"`HG�:�����f�h|��+D�����K37s(\����5��G�*D��:�d̙2�X��`P|1�uq��&D���T=v��@;Aǁ��5s��1D����'S��(�o2o��Ļ�("D�$�2N�b_�L��k@�,s.���?D�i¡�2A`�H�*^�@ʁ���>D�h�b�B�.�#pa_<}Q���� ;D��P�n^g�ZX�׉�"W��Q�$D�P����<���z�޿Av��2�� D��c��
�W$�w�ѻb���p�. D�X�p�%D,pZ���)�H��3D�D�"���Xr&Κ}AB�8�).D��Q�ED %��O�� �q�0D�� x���o��fX���D�Ҩ�c""O�p1'̖&�Y�6Ę�=\H��"Op��c�V!`���P��%`�$j�"OY3��7B�fE�Ri���"Obty��Q�T��jD䑏{�ؐG"O4��cݡ*�j��C����T"O� Q�AYA|��3"/�h	p"O�y�̜�!l�� Xp��)��"O�iH7gYxVy�o� 3 ̨S"O,��a΋FKZ��3�X�lP�Y�"O������>Æ��,щ^�>�"O���O%��(��I׺n�0��"O����kP����w�Լ3Ǫe��"O�TH��
�6B���!L�j��i�"O���@b��1��"��D�����"O��A�|4d����B?quF"O�U3���W/>� ���IZ��*�"O"1b%j�8 �X�RIQ�U=8�t"O��:�h�,�Ĩ���+�����"O�T�R�Gf�Ș�v�[�w��"O�s�/�켨�$	C�|qJ�1'"OtD�@�
�C��	3�H� O2�9�"Oέ!@��c�z��@�Ծp4��Ӄ"O�U�a��73�]�����8�'��ԒA�˸\r��I�m��[�ظ�	�'��=��텾;:��Wm�R�X���':�T>W�^�$��< �����'�:��#���*-+c�K�B��x�'V ��A]6��%�gF�2jRB��'�����-xm l���Xg�y��'� �ҡ�d0iG��2�L���'\�y���K�=��$|��
�'i��#�<&'��c`	�r���	�'�����d�ѓ'�I�e�$���'1
E�S���24l��C �]��\��'����v�Hpa#�'}3X8��'ڔ�{vK@�n`H4��E	!|H��'Y�8��	�"M���<���y��\=��a{&mX�!���P�G6�y�l�K6���Dҟ���Ń �y�l�fj3�띰
� 4\��y�
J?�N%�$���ab���$�y��Ĥ�B�{2��
��՜�yr��1W�N�9*G2��r)��yr��W_z��l
�w��"�L#�y��M�pф���Y�o�*�I"�C?�y��ã
�(8p��)a��a�	��y�� 6M�UbP�N�l��9Q�X*�y®-;X8��>3�9q�O��yҊ��:�v����'s�[�$U��y�%�5�x<aQ��-sp0�B���0�y��1�D%A�WZ��`b��C�yB(ݐ<by�`(E�z8q"�j�<�y�j\�C��m�g$=��R��
�y�cJ�U���U��,l�����y�B� s�P��	Q.̀ʤ�O��yb�1��냤T�����4�y�ϦOL��bH"5ֈrD�E�y�Ł*..�����ݯ�V�b4Ƌ��y2� xZ����-	�.I�S���yRB
�5���!ag�k����I�4�y�H"�J�HQ;�hl����1�yr����y���,�����N��y�#M<\G�;�� (�"5���y
� �����,�L9�AÌ�Y�0uHA"O�a�c-�:߂�Ѧ��s��\�"O����Mz��ɆH�-@�S"O�����VȐUhI�]\؄�G"O>��2MؖM舕R#
�r��"ONA"��[h4;�+�ƞe�E"O��k�I0���&Ŝ[��Q�""O�,*���%\vl����5B�f���"Oz���bâg#\t;boQ�q���@�"O`��@ƽc��0��͘/$R�@"O�p ���~pr��ސ8��-"O\U��jӾ�����̛���Ѓs"O�9���H�J4��ć<"�� R"O�*��(P��i*V�zL��"OVQH�@�S���h3I�s�H�6"O�l���� ��ҀEǕR�:j�"O,�Y`lM':��C&��F�L�
R"O������0�*��@f�V�xT� "O����.��!6  ���%�bY�"OԄڷ��X0	UX<��ZB"O͈3�[�>����"r��ܻ%"O\{����_�D��AÏB���"O��8ǨD'-)0H���,$��Zv"OZ��Sd��8�3"k��9	d]��"OV|brԢ%/\�4�C;+RiP�"O�T�gfO+e���2��X,$���r�"OP�u�PMƴ����B�jȨ�r"O@�)''7F�����@9T"16"OZ��%�o�H�QUΓ6�<���"O�U�@�
�?����6;�>���"O�!���H�(dQc�C�b�J�&"O��qdѲPRFh�N¡���A0"O9��lO�<u��/����̣�"OvI��r:(�(.�8=b��v"Oh�R�OP�oR� CU�|:p$p"O��!�˓4>$=3AC�:9�!�"OBh��W��<W��,p4BT�3"O����"[҂q����#3EC"O�	�@m��W�]���\�Z���S�"OX4(�F�%Pzq 艄K̤ʠ"O2�C�FJb�fo��r�"O��`�_�tM�����[����j "OʝKBH�-_^��p6lP�E��y����A	 Q@D��)`� ��l�/�y�c�aP�P�N�V��ljË�yr�R�y�q���aa� �׋X��y"j��(�`���Sc^X'(յ�y"	ݭ��8!���MȦ��6���ybjߗ��!R0�&BI����yR/�j��P���)3_���.���y����|�i��`a���y��A��y���`��g���j�Ҿ�yBT��tr�L]*X�Z/k�B�	�f�,���`�)I�09 ꉘaH C�Ɋ�L��&�U���4��DǴf+�B�'5�e�6"�3H�D�3"$G2�`B�I9U� �chH.0fBY���ĚxnB��$C8�	5lA�b{wD����C�	�"Z�})��M�b�䡫P� -��C�	3|x� e�c}��%I� JvB�I.u0�,��U�Lxz�.E5�K�"O �7�מJ���i�����"OfY�d��=�T��	�<���"O>l "��
Q�*��������"O� �%31nM�Z�P%,z6]y�"O�lRC�X�z�}#Ēonĭ��"O�����P�0���$�|���"O����d@� �y#�؋�>���"O�*�k�Y�ERL?D�
1 "OX	8�@��ae����mX)r�:�)s"O�逗��1���V��V�XI�"O��K�J�8�n|�"$P�t�4�a�"O|\�#�' pq�!�G{��=C#"O`v�{eDE�A��"�a�*�W�<���N@$:1F�V�\A�!�]�<�ei	\�m���/>Y���X�<a�gT�h�� �w�ӣ�$a��N�<�En�hr��fѡk7�Pa��I�<9���dd���M�%[��Xt-n�<���XފiH��E�������k�<A��O�2gEA�zz�%����}�<	�A�r��,��y��uz��T�<�1n}�؅XDD�Q���22 �{�<�lB�CKd��C�330�%:t��[�<@�B	�~=!D�խ_|:�S"�CW�<���o�h0Fcπ:��wo[T�<�EGH�	�|��Oι^i��ʄjDR�<���Ԕ6�Mb���/(0.�j��K�<��X�1�b|3Vm�,*��Jp�`�<��%��!ה��Q�|]Jժf+�s�<�bNN����c�X`n8\�5��f�<qE��v~4��:9{�h�"QY�<��h�t�h�
4N����x�!�X�<�� $F@C�#�d��}�A&�M�<�l��,���B"P�x���M�<�T�R�Wʨ�j�#_=�*ᐖ*@�<�W�ւV��cnP�T`�#K�<�҄<�������>2}���D�<�!B»c3x� 4�E�3���5'�}�<EŞ8�	x�Nf�,�j��Ws�<Se�����	��]�K4�P��j�o�<!!~��8�T��Α#��Ke�<9cˊ/�<���Ɂ/�*x�6�d�<���F&!�
�	�,lc@�����]�<��0{�N��ui$)&-�N�V�<���"u�tݩ��g=ҝ4�T�<�UC�9T���;�ď�vI�/�N�<�dK�'t�)SCƽ��9�Jp�<�r��9��q���Լ����f�k�<i[R�ŘЬF"j6� ���@GzB�Ih�5��$F!�����T���D8'�`�'N��s0�H	��� x�!�X�7� \�R&9 �kQ�!�� �S�!`�'@�JsƑ:*�!�̾ye0��"j��'!�!�T1����3'4�s���(s!�d">D��"�-D�Xl�p�Z�i!��6:����"C�����ظ)?�B��+}dM��O3r3r���!O�C��S��u{��E8�2��D�[ND�C�c�RQc$(Ͽ0������C���Z �>sY�t��n�jd�C�	oz@��*N+)��v锒S��B�I�]�l��V�L+U�٥�Ў�C�	�;�`�[��&$���4bC�I�W���d
�7.��aʗ���vp�C�ɪZ�$<�E���~ǦI�� AdC�	%%WȀau���F�	+ǎ�es6C�)� (<��.�62n�;�Kś#��Q�"OB;���L^z�B���u��ys�"O��r"m
0�!s,�C{,@r"O:��\�a�n�1&	�lsD	Z�"OH9/���T�FF��k��ԗ�!�D�(:N��e �9��)����a�!��˫-�̕Z��UG¼���W�!�ď�f��iL�M&ά؅�R�,�!�Ě�.��H����4P���YI_!�DMV��)`7�Ѿn���ȧ,�!�D�!t� �A�ėJ�� �Q��!��l0�c [�AoRY�#CC��!�$K��n��[LH�04����!�$��2d���GO�=�F� ��3�!�^�Y�LhY�m� ������J�!���c��6�",{�Iـ5�!��-k[°"F�"c���:�bJ�
~!��Tk�-W�`�*���!�mx!�$�I`t�uI�q���AG`!�Ğ2`(�0�U��Hq&@�:P!�d�)�^�¤��7]̈́�@�`�v!�䈰M�p7LQ�.��d�����!�ą�t�����ݚe_�M�ç�*w�!�@'¤`�&� �/Pnx�ef̼�!�d �`��܁� Ց5=��}l!�$F!],�m�A!�]��g��^g!�dI$k�v@��`���+�!���7}Vޜb����(�옂�j5N}!�D\�tɾ�q��#�L��f)Gv�!�d�(^1�"3�
�sǾd*�ɉE�!��Ú((ʭ��
�84�D���)��m!�dDr�R6bܞ]Q���[�~!���Ci��[�L1{c%͖�Py�c{�L�Å�ٱUNd:Ɓ�<�y��10ypd�u S�d+�	g��y"�]��X��^)�a��l���y�?Af��;W�����@"�y���T%���e?U��c���yrcG�z��y6/A�7Q:��3��yr����A��� ����Fp��ȓ*5�a`�L�(q����G�@��ȓi�v$�&�8|4ҩY@F@</�̇�`@����*D$�lq�g�4b=��ȓDB�A�HB�?)R8Q��J�	�E�ȓ=�Xx3�X;4>�4��#�ن�)��0$dٿr(�9�$���i����c�¬P��R�v�`-X��(��ȓy(Jٱ�F������˟v0��ȓd���xCW�I¬�g��+�Ʌ�^����վ|���b��RG�V�ȓcJZ�곩��^}�ɊΘ�7<�x�ȓ_��5؃�1E$,���w�Մ�  6� $�*|<ҍS��0$T �ȓ���+ul���r)�5nK*@Q*�ȓE1��ƫޔFe��J����Za�ȓD$ژ�%�ҽ�*�ZÌ�!)�x5��y8����Sܨ����T�\Y���$Sƨ�b�܉I���d�CP�pm��0��uY�cGD��Dp�z6�ȓF���W���. �F�?9 ��B'�y�w��`��M2* �c!l��ȓO��|F�/�Bx5h����,��!������×?�مȓ<8,؆�H-i���oU#�M��S�? ��h"���C�<q���'��@�"O���5 ա$R�'�H4[>u�"OXɈQ*Yy��Br��^c�\2"O�� -b�C��3"�ĩˇ"O4����?bgN���N f��R�"O�((�U.����AL�	��T��"O�H��
��RD����2V,��"O���ǎ_(
n���v�f��U"O9��H�g���H�!M��
�'�
pQE����	���lt	�'1|@�0�<
����{(���'��q�aU�zF�Պ�	��}�:ȁ�'��40��<�$�G�ĝv�ι�'	8D0�lȓ9p�,����q����'���c�V]TI:a�J�m��)��'|.�ja�E$NPH��Ё�5c:��'2��z�a�y\"!ѕ����y"F�.�2(����֌���Ϳ�y��J&Ir�y�WJԛIo�B�ۅ�yrh��/�9�e��B�j*�bÇ�y�#jI�C
2(N,��$h_��y"Έ9i �%�*�9��QdN���yE�)=�V��VIٞ'�ը���y��ˁ42$!����Rkó�y�n�xf�+Q�*�Εj�B���y2,�����v�Q�m?\|�f���'�$�*1D�>D��x�dM�\�i
�'���r��'^��0b�]�B��	�'+,��PM�&Z֐�6	G��s	�'3̼���Ϻr� ��'��Hb(q�'��͙ue�>GB��G�i\��(	�' ʜ�W�N�S�Xs`'K�j_�=b�'ɖ��Uė	C�Tyv�mth��'��!:"%ec$	�5��+4��"�'X�FN�)p���K�$@�@�f4��'4�P���Uq }Z��99�`�'�@�GnM�l�`8`��j���`�E�<����=P�l%�@!!.��h�|�<��F0>k��)���V���l�{�<�!2[�hp���Tj��U}�<�WdM|1\A2b�ͯb%�%+�#q�<9���7bú���#I�@Lp�:��HH�<���r�Eqa���M	$�2 ��O�<�ҿ�7=�ux�aU���P�$"O�8"�&��"R��p� �a����'"O��X��
�tעT����JM��QW"OlzQ@����3�o2t��"O&ѹЉ�*Y��P:&�LQF"OH8#�gȪb���j`�$J����"O�����(,C0��C��pЗ"O��I7/�7��k���[yJ��S"O"9a�Ϥ9��u���m��j�"O標�Q$M0Ā�@[E�P�"O����%��
8X$��C�Q���g"O�A���!	��1j��* ����"OZA���
? =���m��=����f"O�q�!��F`��B��K� �T0R�"O�9@�(o�r �q���KG"O�-�%��J�	襌��}�*���"Ol��oE�|�8��L���R� �"O.��^�E��!���R��'sD�@G��t��ԡ��2Q��(��'�0��r�(#F�Q� ���G�H���'_ �p�썮|�����;������ nAz��ȑ"J�����7NM�h�"Of`��m�"v��u��?+\0�	v"OQx�����%�B��c&ؕR"O�웕��E-,xЇ�!* �a"Ot,A#�Щt��T1��d��"O���e����`6G�	R�U)"Op�z� Ѹ	���d�ۥX���p�"O��ۑ��a��X�0��,�����"O����ㄦ1�(svE�%@���C1"O��g�o�P-��^�]tF@�"O�+���o�t��T�MhFᨀ"O�B���i޼YB pfh<[�"O�x���#'4JQ�U�&Z���"O0��B�#�U�,�7LJ��R"OVU����&A�Љ;e�@H9�ؓc"O�ԂR�τuj�y$ ��5�q��"OL�11��82��%�N��z�ґ"O8l�V�s5��'+
4h\�Ճ�"O2���D�:��xx�
s�B��C"O.��.�;%������0���3b"O��v�?e"Np*�._ �`؁�"O���d�d�,f�
���9""O��S���c3����g�! �"Oy����>�&�(���g���S"OX�����g�0���S%$�)�"O2M�.��ԕ�F��K2���q"O�a��H�M��=+�K+��rv"O�؀7o
�t�zla�I�"'b�t"O��A �l���  *<s�Jx"w"Oj5	��A;m�0�h0��y|�x1"O,��gJ`��2Fߵ�P���"OD��o��WL ��qŏQ���"OL8�h��l�&�����o4I��"OD�!��.N���Ti\:Tw�,
3"O��$.��|(G���aFA �"ORh(2� j�|�ӈ�>M��i�"O�!��	ǜ��٩�%�4IIP���"O���v���HQDdS@AV�+�"Oތ��%I�z�#�Ë�6�Z�"Olt�T��1˚����C)u�.�A�"Or� 5 ���$0��(-�¸��"O
͋�ߡiP0ZraC�W�}z6"Opm�Q�57��W`� �0��T"O>9�l�-A��PAǠ�2`ȈQ�"O�X�6�H�DY��kT!W�u��#U"O�� �BM)2�y���,|����"O�"��8-��B�
ߒ-��m�'"O�b�kW=1�\[�/��u���2"O�32��
'�HH�����Lh��"O|�9��tZ�Y �Bǻ+��a�"OBP0�j�Kf���C��)�"O$dQi�R����D/�Y�̘g"Or�3cU<YST�Z�$�QD��B�"OF�r�3_f��hrE�((Z�j�"O�b�K߷_��eS6�Q1yz�c�"O:p��F��ܠ�)x�$�"O�؋�dK&HRQJ��W�`u�	�"OD��Ba��I��\CF/�
vK^)�t"O��H��!u|}��W:�!�s"OĴ�QR�tO��@p@�;�,qK�"O������s��=J�͘F�8��"Ot�v]�s��`��ۯ��\H`"OR���ϱ+�f K0L�Ds:��"Oz���d"����_�|�&�0V"O� �  �J3 %�,z@CHV�jt
�"O�11�FW�0 нb�We�ly)C"O00pFO�+QB�C@G�i#z(�"ONm��p���S�%wDAK4"O:��K�N�&a����:b`�"O�	`)� @c����ʞG��;�"Or�Y ܸ-���u_?i��YKE"O�\IE����*�H�(T��|#�"O�}ا��v*�<��˕k�̀�"O�EH#`ĥ'��0�UAGx�8P(#"O����$1B��/�N��!�"O<��B���A�|DR6�Fnl�A"O�
�	XH�:��NyMps"O���E��^���`�Ĉ|vЅX�"O�<�B��j��3C�Üx����"O���6GV�"o8�Zf�,s����"O �g ��l^�q�Ď�,��)P�"O�5HNL��tZ�ү
��Q"O�����'�DГ%�>��"Op�[cۂR���D�Z>��4H�"O�	�SH˥!���k$��ti#"O�d `
��>&�;�KW�?�py�"O��Q��3�XI !+U�ީ�#"O�D³��(2�$6Tm�xÅ"O��"BL�,K#Te�cC�(yQ�|��"O&5��MO�}�`��_�G3���"O�)P�F���Ff(jw��!���j�Ղ��
/�� �e���k�!��ا,�h� ����W�B�e�!򤖰g�渂��Y��$�"���su!�$�7$��T"�Cז�҄��'=t!��vJ����]X0,H�� !!��ܑW�����+Y��$C�vR!�D�J؞��3�U�4VN�"m�9Q!��49de��͋;��T��l��L!�dB�32�I��6(�pXX��ZB"OrP!Xp�F��4�Q�?�^�k�"O(�8�L�=v(�0é�?bD�
�"O@�kS�E a��@��	Y�d��"OH�s�A0��t3��&9��X�$"O�m "l��?�� R3��41� ��c"O�٪&l�$
�l��-�
|=jŚ"O���aI]�X#���C�,���@�"Ou�l�}��10�ݙ2Z�i�"O����邆~`��#��ux "O6���-�q�`�d�:#X���@"O0�H�~`�f��#*�����"O��� �BV�zc�S
P��dR�"OT�SĐ�O��aAN�e{�A��"OxpI��ARNHa#���@��"OTС�S#x[�]����R���R"O>8
!�ƃ`H�׊MXX��"O�́ ��9&H�ŪO;c��2 "Ox�6 D�Y �hE��{�(���"O*`��'�E����+�r�pa"O갢����G6�aPc��6<�A@S"O0��ס�0��)���Z+2����"O$$ qʛ�q�$8AQ���Y�հ�"O��gG�m~$�g��J��y u"O8�kP)��B�X�yP�� {��Lz2"O&=��%؆2&����	=���hw"O&*��֍(����W�Ҽp�4���"O�}2��n"Dj�� >٪�b�"O6%P���8�z��&�%M�@���"O� 4����u7L���e��,�8P"O���
��T���dR=f�p��V"O
���
�������'�0u F"OB�{��ٯ9\J1#��W7%b<�f"O���ĮkNX�%���*�}
"O�Qc���"T	��R��]���� "O�Z�@�[�9`�*���8t"O���&*��6r�u�Pd �O�؈��"O(��P��3�xׂ�>J��<�q"O���A��+J;z�K������z"Oj�t �$�bH"��p����"O����#!5����%�4I�"On43ѩ�3B$���T���`"O~��vȧH�8�eF�uc`T��"O4b����g�|E�fոY
�k�"OlQ�M�
!~x�hB$G�uBt(z�"O�8Å��P�Z���	 3-�Q"O�i��E+������);��b"O֩pp�N(t%���@���)y�"O��C��� Ya@NDU�R��"O(�mT oLa�1���`�.U��"Oҹ��8v00���? ����R"O�9`
)&R�Җ�96�h��D"O�,�&$��uq�#�h��^���"Od���D$FXp�m��?�����"O��N�}-���-�63�u��"Oh�)��'X����5�K�A\:ų"OF܁�Iتc����!�JN���"OX��c\�E�H e�.>@p�U"OFd��_�N+��їCλf�����"O*8�!�a()����'j�B�`6"O��g8*Y�8V���}��"O�E����� �8QTN�O����"O���V�Q�U����m�4�L$��"O��ȃKà \���BƀK5x�"OL��R�]�v�ä�O<U.Pͳ�"O0I���_�*Wd)ɳ�*l,L��"OZ��R@�7�v�t�� !#B�t"O�� 'ɖ�E��b��ԙVH�+R"O\�+'cݳH,�j2F��RjT���"O� 0C��^��� ��)UW�L�"O4Q����8k ��:�ɑ�Y�� �"O �Q"�;�樒Ү��e h(�"O���rτ8cg��i�mH)f��đ4"O�3AI�H�� aj=�r�"Ot�
tN�O�L�b$
ɣb���"Oj4��l��X��2���2<���*�*O�m;i�,^>�MJ�(0Pf�0��'�m".4m�а)�ۜ0�$T`�'���H��ЭB�8ȢfaZ�'��dK�'QTh�3�(�t����q�'0΅
�!Кt) �q"F4����'!�a�q���
�P�0%7%pM�	�'#�u2BfǦki���JԠA_�A�	�'�Vdi�T�3�F�Z3�ɝA�,y�'\ }�A�G�<�2ƪ��i1����'+VX���аy�J(CTihZ�'5��G��3j���c�,���'��\�!gK(z�rfϏ6;R�Q�'�HI��0)���+�e�5~�v$x
�'��:��Pg�,����)C�ax
�'(	+����u�@s�$q�hȘ�'��-�$�V�%e��a�Q%4w�5s	�'�Pu���"h�`���~��!���� ��1��@I�����落C�"O9KE$J�;T�q1jДjZi�G"OJ̀���.����G虩PPZT"OfD����Uqb��`MįGb( W"O$�3�ꅞþ�	�J��h�T0@%"O �z���1��!�ȟ]��ԣ"O����T�4|2�d[2�b��"O�H(t�� ˌ���A�W�4���"O�(AlH�y����� ݼ��p�"O����&�!m�ޤ+�*��UِU"O��I�ٳ)E��Rҧ�Q_�E�3"O��Cro�(!4����K,9�^iW"O�m@����f�1��T'�xX�"O��R���k��q�(
�j��U�B"O�qd ���$��F��K��]��"O欓A5�2d���\�4�t"O�5;e*�,>=�yX���ȭ��"Ol���>�q)f�!��KB"O�4���N��݈`{�l�"O�p"�(^1z�����%��W��2�"OX�uNY!S��d�4�O�WR��!"O"5j�MZ�-a�����0� l��"O(Q���8����½Ӡ��B"O��0'��<�<�2Do�q2�J@"O�ͪ�ǣZO������9x^}Ó"O��r�o�&3M0�B��J�cY̔�Q"O*2�,��_a�:q�r��T"OTh��/z�  ��L)m�^	(�"O`� � �G�H���%C�S��٥"O��@D�����q�$��9�D5x�"ONI��c�7��,@�>�>lѠ"O�=Y��	P�lH�! \��ȣ�"O��0�� =��42@S�TVj�В"O&p8UM��".�0����'Ql�`"O��y�L5$Nع
�dό2��"O�ܢc\0,_�
vD�9��$	�"Ox�9�!�#M�Ѝb"���s��ԃU"O6�Ф`��*9���Sz�h�d"O��Aq�O�v���wgE|_j�A�"O0`!��g���Y�ET?z�U"Ol;�ᙀX%���V1.d��y�"O����a�0�(ĂaK��FO в�"Oz�����
@�41�jY.@T��""OB(sW���A�cĆ�07S�t "O\��ȡ-��9+�d�Vh����"O�q�ꐃ�8�Q��M:h�,hr"O�Q�a'G�S��tW��43��"O���%�* ��!5R�`�z�"O���4��4;��H��76��"Ori@�!h,0E��/)�`��"O��Z������� Y�DY�1"O�@�ǌ9d������-/ܥ��"O�����ds����� v��M�v"Ol���d׍: ��B�Q3�^�f"O���7D�oJ��f�DrB�C�"O�P�G�F'ٸ��#��hh�9��"O
�� W�� 5�D�g�^e1"Odيc��2�LB�hI2|�� '"O�x��'; vt���Ĵ]�Jp��"O��0d+�lv�����۞���*�"O�]��i�-u`����_�B\�"O|a�Boϥ9@�	 *�4���H�"O�y������Q�C}F�uQ5"OZ4"�E+�t�ڐ�/@58�"O� ���L= z���N�=i-8Tk"O����A�,7xu���1}���U"O�A�@�*g��p4�(]�.���"O��{ ��?b9T}k"�,ڤ-�p"O� *�;*��M�P�>c.ʠ�"O�I�$h��\�.��
�!v���`"OfUx��̄<�n�H�R��"O����o�(� �q�&�'m�Z�##"OJLz� J;
��t�����˅"O(01F�(���%4@t�35"O��gE���� �!t,�H;�"Oj�h���tVi��͹	��� "O��+woI�W�a��#E� ��"O��a�:V
�v�٣hB� @"O�};"��8r<�r��;	S��+�"O��@�)Ez�h���I�E�j�"Of��ץ�!:@r�	�H�}��P�"O�݀�E�LZb!Z�F��F���RU"O��c� ��l�ZD�P�]����s"Oͳ�g� R����C�
`���E"O�U3�KǨ�)Xaa�#��Ƀ�"OL+�/�=��&f�q~L$�7"O�18QE&���@��Q#|j��"Od�9���v7��C �W�:�n��"O�,p��L�����,L+$��J�"OD=8���w{�X`�	JP|���"Ox쩵l1a�̪�	�C8:�;"O�h&CH1d���u͎4|QA�"O�����s	��℞�y0愁3"O�@��%�� ]AӁFi���"O���NO:!_hEI�@υqFy�"O�1��%��W@�0�^\��"O��Ks
F#�.]���9/�j�*�"O��a��]�8��0�-H<vx�"O�!�s���B(�)@��Rβ�@f"Op�j *ҤW\�E�gI�O��P�"OP��gQ.JBDKU��9贩�"O.Er(A<X�I"�&�q�H�S"O�H����>��M0�J���8�"OZ����M�$6�p d��zJ�"OH�&�Ň����"��m��q��"OR�jY()WH=��.�ʬ�V"Ol,E1B�R�:v�(s��J�"OD��!�B�[�t0�x�&a�<U� C�I%m�D�p��8rj�2�L9�:B��?T�$jD(D�Zq�11�e̠_�&B�7�~\�0�Q�vIu��lM�B�I����D
�S�8ՙ2�j�B�ɀd|x)��P'\'��Gn���B�I}�Hb�A�<���rEgZ1SrC�	Pj��Ƽt����P��B�I�Bs��`C!�n��<i��¼B�	�X�Ȝ3B�"yHtI���&��B䉎/��}E��'i@�#S�<��C�I=a1�MCV/� V	Z S�q^C�I�$[���T �==��H�F
�V�pC�I�"�"��S�E:��q!�N &C�I�;[~T�v�k��X�&��B�ɽ  ��"w��UȜx�`��#�B�VjǊ^�F�)�E�$;�B�=qs��xs R�P2+� ۷*�FC�I�"�8v�r�𦂘�O2tC�I�"m��:D��3U$���B�	7/Of�`�=*ΥZ%h
%((hB�)� �Ģp���w����ʪM�Μ	d"Ob�!���V��Z��V�?U��0�"O�q�d=����B�Q��Qa0"OȈ)�ߪ4��M���۪�"���"OH)�J[$G����e�i��X90"O��	�KOn�\�ʁ�I�T"O���C�\�/�����
����"O�����p&$�SD@0T���7"O�M����O�����R�����"O�kf ϗ!�x�B#��_���[v"O M�ㅨ. �Pr�+�(��AV"O�M�ָ�<U��jI)�@D�7"OrL�%F�0�ƍ�`k�\���#"O$Dp E֌oNZ!`5
��{�Ex�"Ox���Ȅ�NX���'�w#�rw"O*�
k�lL�����-C�Ej7"O�����3A�xL���E�����"O`�q#�n�(� �ϬC�b`�"Oq
ȓ��ȩ",�G\`x��x�)��gz���!�Ƨ~���Ȅ�'j�B�ID���rB-C.$oF�Q�"L��C�	4�����R;Ό��e�%zEBC�I1z�b�`b�I�l��A4M���'>a}�nȡ$o>hzu
$9�9;�O/�yb�u/�,�DG�iR����y�d�F��YB��	CB�rg�7�yR/�3Q�(�N�7j��f���yR�2 ǘ\���Mzv@̢���yBB�,ẃ�H"lJ|�u�Ф�y��Ӎ%'�ɡ�		d��y��ܨ�y�e�?j�.��
[N6d���T��0?1(Ox�6��=��� T)C_$L�#"O��2��7CIdY��V�U����'=��Ǌ�	;�d��קc����b�oӾC�I9��� ��-pt���cF&CeC䉼I2`�AC�SV����WӨB�I?b8�\�7ᔀ�RY�JA�B�	7nt@�G��U�<yZ�M��n��B�ɢz&�H2�F��aez��oB�R��C��$=�RXp"�&N2�q�����x�NC䉢㥮
9�.�#��S3�H���"O�x�Re��]@�4��6Ȓ�� �'��O������@�8Y5��N���"O�A��"�,O&��T��	q���T���'��''Q>�q���9��YJc�3Hm���2�*D�x�$9�Ll�,ٝO\���h4"�~��I��XM���"Y�
h(�CC�z6!�$�s���h�J��3��,a7�ąP��z ���\ä)���((v,k�h��$F{�O�R�%}��?-�R���9�IjD��yB��[�X����+s`�� פ�HO��O��>�D�&/~���H�&ux���3�O��j�qH1�E0Su(���[.bt�x��S����8�D/-�� �蓿Cl�s�1D���r�7t�8��"dm�/D��b���s�؀;Pj̧N >aP�L��$G{��	�.eF���)^�L��a�K,9�!�dQ�a��ᄍS,,d$Bh��}�!�4#BJ�j5�.[l,��R�f!�D�4C���[��VF	^��D !�Dس:��S (0���P��",Bf�=ͧ�hO2]�&�0Q����h�*��Bd�|��'3��G@�T�b�.Ů��x�'f��:A�S*ݑf"�	~�p���� *�G.��i�l�%O�+�P`@F�'����|_��O���S��l�68@Ԩ�Ё00x�>A4(�'̀�В��Y@���3$`��'�R�D6�ɾ�R=� 
 $���	����$<�\���'�ƖPWXzPK2a^&��1�*pGV/`©�C�1b�.�ȓfx��Qn��[@$|h�犵fi����@�HK�;�%<2�V���ɴ��֙�����x� ��]0A��az��8D�\ �#�=��I�WZ���D�7�IŦ]GxJ|rr
���X{W��/?bVY�ĭ�S��d���O��xp��;*��/5(�6"O��0�_0?�ȁ����c�i83"O�H�GJ�&fJ�mYQ��DP��9S"O:�h�B��m�|���7A�"}֘��	a��8��/�[�����e� ���`#D�l*��T�hMAB��j6N�Rg5D��8u`��gDL����[����=�O<�O΁���Ҝa�1��թ&�Lsc"O*���.�PR�X�B�@�z��z#"O�-��OQ�಑�d�Z�I�<Oj���<9�U�\$"�͝�Z>����".oj`��	�<��{�,�@.�Р���Q��� ���y����ZG��p�����㰋�y" ��Fd@@D�VEH�
�2��)�S�OL�mp"�L!�fى4 �+n�\��OP��$�&x�\X�.�6|��Q���%`���|��H� ]��N&@�f�R��3i�b�
O�6�D�<0�}Y��-��t"`ӠF�1O��'B1O�O�dɨ���][F�s��)P���'Nb�I#��
 ETj���蠉�'�@e�ƬD"\dp�������4�hO?7M��s�@�2	>z�� yu�~|!���?QD�ܹW*q]
HQD�]
\�'��|�G�~����%ǫ.�R�e�֢�y��Ɣt<�!kѣ����Z�.µ�yB@�)��$�sʌo�%�b�y�iŐ�T�
׈��8��"�y⇟�)Re�A�C�֡��\�y�K5W�|IWMil}�R��:�yBGU�*X�$[�
 e�K!�F��y�٘`Htv ��~�6ȰiX2�y�LO(E���*�BD�Ln�\�b�	���O\㟔�O
4	��ޅ���b�ٛ(S���'f��p��*Si��ĥ���4���'�|���d@�C���{��ʙ����'��S`�О{͘�8��j� Ĉ�'��<�� �/�}�de�uPa�
�'�|��&	�}JQ��i���c"OBX0*I�-�(s4��l�Z���"O��`ѭc��f����"O���`$��{!�(*r�+bP��!��0�S�ӣB�<ٷ�O�sꂹ�FI�c�B�I�/���&��*�qI �\�5�듅p?�&ȆENLl*6GXG)z�*��_|�<92j@�"Z��B�%4n��A�ֵ#�!����\a 6N	��Ҥ
�)���k����EyBF-)�h�R/Δ0j�p�%����O�~�3��IUa�2B�Q�M�g��Z�I�u��#=�M<qR�Vy� }1d���o��T1��P�hO�>�;�'S�HA�eG@*�-&J6�#
�'�:�P%�Ԣe$�ʥb���╚�O�c���'���~:5�� XfQ�A�/TV9P��r�<��͑�`E�D���.]RYZg���q�<�5�O��>��� �!DF?q)�X34f�=N����"Oʙ��iG�X��@K�*�?;����"O�M2��R*hq�����?e�ސ����m�Oh��怉;����(��4�d�8ŤX֟<����aO�8	?J���P���44jC䉒C͐���O�"�T�1+�s�ZC�I[z�}!M�p���j��ٶ 5��Ҹ�u��s�I��O�G��ٺ∄'y��8��0D�d)�o���J���	 ����J0D��*T ��)A����_.$�B�d-D������XV�T����\<;a�+D�d�f��_"LzS#�J���GJ)�O��O� �*K2&r���C�-�1�i���' �E�Q��2#����@L!H-d��	�'#�a���:J7����K�B�@-z	�'�"S�R�qV^ ��L��q�5��'�~I�WJI4��4���ns�8��'q�Yh�ɥ3��|�%�o� MC�	x���⇕������O��/0�B�II��� ��3��|A���:<^�C���>8BG҄��U���ĬI��C�I�ZD�1�'�͊YK�u8�/,Q��B�ɉ�t����
�#��*E�C�	�ԁ�5"�^��c��@�>!C䉡aI��i���%Z���9��B�68���(� �3i�}ɕ��ܴB�ɭT'<x�F���&AµZa�F&�HB䉗)��ᑦ%��)AzA�J	��B䉲,�TQЁ�غiy��yboԚN($C�I�r�]��/�'��i�%l�<C�ɾP���ɑ����S����B�	�h����A	���"I=ʬB䉻(�|U�3!Ĝo�@ 9%�,V�^B�I�S�X���d�-Wd<��oP:U�C�	�\���bs�^P5:p g���6�C�I8�ب2���=t���k�)BZL�C�I��d� ��&�@�m�?R:B�	')	�����!��s��%tR�C�I�qv�IÃ�~�%���8_�B�	��x���G<e��`�g섅e��C�IJQ�l22jX6�>�H2��:��C�ɊW����㉧E�|�i�"�`"�B�I�,��͚��f�{���`Y�C䉤Ww�`q`�c�6�&�T0dC�ɦ�B�j)Z�t� 	xQH�A�"C�	1=BP�r'�:-���ۯ%�C�I�aF�� R�m�����&D"6C䉢iP-�0*ǔ2
RՉ��ىP�B��8;�T�JF�L�����	%q+�B�ɃUW8 2K�1��!�uh
GŜB�I����%'� 9V�	���݁RabB�IZ��!�K��b)[#��,FB�I�`K�pҡ+_�9�R��E n6HB�	�OXd�a�H�<<�q�êjZB�ɓ9d�k�(�6j��p�KԚu�B�ɾ�Lp����@�y��0d<B�I�^:� C �9B�I��1�B�ɄJ����R"$6��%�Ci݄B�	y�`��u`V!jI�ȁ��.~��B�	%	�4�5Ⓓ>�p���7��B�I&�و�)Z�=������	_��B��<az�9s��2��8��9L�.B� @��	��B;)�N��)LC�~B��7m���NA:5'
hcU��9�C�)� j��UL�j���i�/�'�컧"O\lq��ßNr����I�P��"O0ܺ"	�D�*�Va�4����a"O�a���'��H��WJmt@"Oh�����h�<���ؕRd�"O����AL+Y��)�+Lm�TҔ"O6)ISn��M{$=�`��<J��t"O�q�&�·N^�a{��6O0�)&"O�@n Ā��A��Ġ�V��K���qOQ>a��b��b/��t/�-p� x��J*D�@�Um��M�m Vk,�h�k�-}�V�%[�:�d�[�Q`ݒjт8��犸BC��Sw*+�Oԡ#���3��E"  �"@��E2�d?ca����%]� ��$��/�mɠ���M��)���'-Aў YVf�e\<�Xp��~ˉOl�=Ð���~v���Ǌ kt$�'�b�	��BM��
�R �� ���Td�,Ld��
5���"~P�ӤP�ѡw8D�"e�d��y��5�����S��tQ�B=cj�E��E�D{�+�@$������|���N�*1"a�.�!�a`9�OF)jPÁ�J�"�ieM�
TĤ`�ֈܯ_��[b�@�S��hul*�O2�S4�^t���R�E�"����I.&��	J�C9E��K�^b��Ny@��)���z��)��9>!���G��A���^�"Et��Fn�*i%�ƈ�kq�ä��U��9@��u.ڞ�(%?9��L��s�0Q�Qb��Mp�O��π�(�/3�O�M�5IıU56��!ҍ�!iA�4�?AE�C�*2��������*�����I &-f0�V$�̼�a� b"����,�.`Zp$vИ�JRԝ	�ę=q6���q`�{o�)ea�yr����	)
��b�l޹�����
S���wǌ'��90�L+�"=����(s���k"C�o��j&�>i^�2׈��Y��qcfџ ҴY�G'�V�je��nN��y2[%~qN�X�o'[��Ez�OW��M� R���S�FF��?IQ�Q5*	0�yA��?7h`6�_�p-b	ڶ�i~B 
�?����5��T��c!�P�AN���� �~ 8������i��	��ꈂKH�A�GX�@��݈��0M��0�$��7p�E4�ZͺK�* 8mZ�8¦*T�f�ŊP�%T��O�
�3��7�0?q��7Z�I��
��\��MD�M[ Y�G�5��,*`�I�z�X�ä�%z&dK��"�ug�7�$E��Ȝߋ�E�z8x��-�l*�'�NI!����f.H��B�N&�?a�JT�lV����@�&a�9^v�A� ��ne��-Lj���Հ�x5���W��LDy"D>�z�a�
�IB�H��]��+Y=��~B/ȉ)t��"3J�����$a:��b��?%N��%G�=:P��P@P����+2D$Zx���bzp3U��!X�^� v�A$Ȑ���R�=�EI�d,d� L�axtl%�P�]�����K!��'n:H�1�Ա���`g�+A�<� �']T��G�J16���-=V,MʵE��zq���#�1
x��s���[XPͧJ2<�S��/;]8i��w�$�HR��s�6X���'5
�  �5�%mÏ!�~X�akŋo�F��BP :���"5�G��X���KU�-+�é�*W�lx�1��k�R����|�H=��	�!��:$x�-"��B!��O�c��0e0��c�O�A&}H�< }@��"�Ph-jiö��1L�3� �*�����6lY �4H�qX�,�¢	�gC���5�\d�@&-p�4k
]tV���O�b���0bK�̰����^`�H&M�+'�h0�l����̃ ��B�l�@��J���xҧXh�Ɓ0�
�(��!��}x�e��ȝ�ẙ���C����Ƿ�B�ⅺin. �oj���]�h[�(�P̾#�4�)7��9B� ���\���#�O�!3��:��!YӼ��ve�w�%8t�Ȫ��<��-�i[Th���]�F0��"�\ئ���%%�U�FXY��еٴ\���n\�cD���jV�S4!őd�Y��K�N�8�q��Bv�@���9bFT��+��K���
��b��遛'�8Ԃ�I�k8��u�í:�R���.ݶAc�gI�[A2��ST;�n�D�4d�������?�Z��P�,ٲ�'#n5��HX<Z�H	 �R����r��c8������I� ���}?�+Ύ���Q&�L�	!l e�P�����q��L�(m:�&��|ʁ�c��Y�t/�' m���[��sDG�4�P{uaQ6\sd�'h�-��*#o����EkYc�dM�@�n���K�2FB&�FM��?�&	��	 }��D�i��(��R����0�'CA �v�>�A���'��,V�2T E�P�~�d��Y����Cl)Y"���':z�h�eM`�@�� A�?���,i�$���)\c@땦��w@�Q�E�'���	�S�p�1PȽ��0�UR�:N|��R�ʜ2Fj�!�Y&G٨b2A aĆ�a�(%lZ#5��0E�iD�1�تJ(�d�Y��y�O�XA" nD� �YGU
K��9CΏ.w�HHp��vvX��d��]�$A�:���2�IQ�>n����	
y�v�G�lƨ��.o\L�X�̐�h0l|��l2�����'���ǅoǲ�q Þ�kT\�`�,P�j7p�QB��n�<35�S23������a6���o|8:a�֬2M"����?�0s��\�t���"�H}1��\�$(�tɀ�{���mZ�.��+���#� ���;O��r �8�MC ��/����؃��n�i���/t���`׎��a� n��,q���
oځ��o�i���*y���f҉��j���K�)�
�ZV���IO��e���C�,��ZU���CG��n���K�)�
�ZU���CG��k�]g0�����8hb��?f�Um;�����2bj��8a�^`6�����4gj��=f�Um9���`���ZZz������3�p��h���WWq����3�p��h���Q_x������?�|��mI����v����4պ,3�N����{���3й.3�K����u���8ص!?�L���Ny�,���{P� �D�I���Ny�,���{Q�$�L�C���Bv�#��~R� �D�I���Ny�,�s��p0g��`�xd/y��s}��w:l�
�l�s f#q��xw��r8l�
�o�tl(|��s}���ڸ���
R^'���|)c"��Ҳ��	� U[%���z.k*��ڸ���S]"���p%g'��Ѳ	^��e]
ŋ<&yhX��LwS��lW͍9'yhX��IqY��g]
ŋ<&yhX��IqX���08����		���sv�5>�������wp�?4���� ���rw�5>�m�
O�9������ܺ�/�)�n�G�2������ٹ�/�)�n�G�2������ܼ�(�.�i�D>ki#�FǷc�r��Nm�9oo*�Oͽj�u��Li�
<	hi �DĲd�x��@e�;jj���$��[�bӷ@~)	�����$��[�bҵB}*
��	��� ��Y�bӷ@~)	����x�o^M"J��W���H|7,��|�hXH&L��\���Gs;#��q�`^O'M��_���@{1(��|�h<)a2��&���PJ��s0�9,e1��#���TI��q5�<)a2��"���XB��v3�;/d�(N1�Y��1tyV�ݘ�ϫ�!E:�SŤ6p|S�؝�ɣ�*N0�[á5q|S�؝�ɣ�(J�,�����H�@���E�؄��N�*�����M�B���J�֍��I�/�����O�G���@�߃��I�-���mьg��;ꝉ�	���d@	��jքn��1㕎����d@	��jքl��7䝆����cH��b��U�tA?�Ag^�"m}���Z�r@=�Be_�&fp���W�|K6�IoU�,m|���R
��}�4�wJ��W�Y�)?�Y��}�4�wJ� �R�Q�#5�P��u�>�}C��U�Y�+=�Y��~�3Ҙ�]�*��`tQA��`*:�ޗ�W� ��by^K��i!>�ݔ�T�%��hsTB��c)9�ڒ�P���Ǖ5��Y��UP��e���͞9��P��UU��o���=��T��\\��j����G>�K������9����K3�H ������3����B;�M������3����A>����~��5�7���,�(�f����q��?�>���+�/�h����p��9�:���)�(�i��������̭#����zo>������Ī 	����zo>��������*����pg4�������"�з���}����kp��-�ڱ���y���t�ep��-�߸���r���v�jz�t�'�鰪3d���gl�� !��a鰪3d���bk��-,��kạ>i���bo��$"��a貮6k5���1#�²Vf�D��Y�d7���6!�ʻYl�@��[�i>���;*�ǶRa�M��S�l=���%����.����s�D��rrd�.����%����z�D��{xk�&����*����z�I��{j�-��J�(����s�P�[���K�+�����[�Q���A�#�����[�Q���@�'���3ÞeYcs�N�0�@L(���:̐lRkt�E�>�OC(���9̓gZ`y�J�0�BI"���0��:������g�dH�l)k�H�0������e�dH�l)k�H�0������ b�l@�k/l�@�8�����0BL�=�id
�m���K���3@O�6�ei�c���C���8JD�6�al�k���O���W�+T��,�1��H^/�X�KJ�W�+T��,�1��KZ*�_�LL�Q�,S��*�5��I^/�]�HH�W�+U�������S���9w�ױ�����Y���4{�߸�������Q���3|�ڼ�������,u26^�9�����c�����+ }:>V�?�����g�����,u26^�8�����f�����&R������ʡ�񇸠��N�\������Ũ�������K�Y������ƪ�������K�Y��� #=����N��`��k��"!<�
���D��i��m��" =����N��a��g��%$:��И����ЪЇ��_�����ӛ����׬Ճ��^�����ӛ����կЅ��W�����ۜ�-�lR1��F���wyc�9[��(�nS1��C���qk�>S�� �iU5��G���pqk�1S��,�lEN�tJ�!�E�H����$�EN�tJ�!�E�I��-�NB�xA�)�@�I��%�EN�t%�/�9�_'����MmT:<"�&�3�W"����Nm[40/�&�<�]'����KjS=:%�/�j}}��W���vypѨ�#��Wmuw��Z���}sx֭� ��Si|��W���vypѨ�#��Sh~y������H|��ko�;��B�����Jx��af�8��G�����Ap��bg�8��G����ux�=OF�B��&i��_xb�u{�;JL�I��)g��X}f�t{�8IL�J��,`��Upm�||�;�9�0>��-}O�)1"f��:�76�� pE�.4 f��:�76��!s@�&>,k��1�?�i��,)�Ʒ��\����l��-)�Ķ��_����a�%
,�Ƶ��V����k�����N�e���@���}�����N�e���@���x�����B�o��E��������N��S��}����P��T��ic��^��v����S��Q	��gi��Y��x����P��T��ld��S�y��K�'8���MK!��r�f`�~��A�,3���JM$��r�eg�y��K�'8���MK!��r�gg�x���r��gM��1;�]�EMY�x��gO��;2�X�G|H_�q��mF��83�X�G|H_�q����c���y�1�a��v��<�� �e���s�;�i��s��<���g���q�>�a��y��6����jE��j4�� (YHՁf<�^�o@��c>��	 ^Mуg<�^�o@��b<��%[Hׄo4�V�h E���H*A���f�z��B���zM/E���g�~��J���yN.E���`�r��E���|��>�W�x�#�߈�5�_�4��>�W�x�!�ۍ�2�X�2��9�Q�}� "�߈�5�_�4��>�{��K8汋�f��9�"���O:泈�i��		=�&|���K>ⷌ�a��8�!{����R�j��8�E���{m ��U�o
�
�;�E���}d*��S�j��:�C���tm ��V�G5���O��*h6!��t��@2��O��/m3&��x��E7��J��/m3&��x��G3�t�b��v�o�z��N"쇛u�~�k��|�e�|��M 삟r�v�b��x�b�y��N%뀝r�y�b�Xlh�R�qD��q~r��W`b�Q�rE��q~r��W`b�T �{
N��xvu��Ubcv�r�1.|-,��P�E��g]�s�{�8!u##��T�C��cZ�~�{�:-~"%��T�F��d]�v�s��:�z1�����K�D
���$��:�z1�����N�L ���(��3�|4�����I�@���"��9�{!�2~I��p��/~��̠%�6uE�}�u��.~��Ĩ#�1}L�w�}��$t��ƨ#�1}�ށ�@_�j���AV��@cu�ӌ�KU�m���@P��Mgp�։�F[�h����E[��G`u�Ս� zt��+� K85B��
�{�9�3��4?��)�!Ē!B�d���Q�:ebD���d�4=�1P4�B+-�,0b=�0��&�Dt 耂�%��I�Cȃ	f-`\w;����@�:r�$� �B�F�F  �I�D 2HТnLR�O��j
Ј��S��O �+��"D�~(��)�<Ee�	8@��%>@��!�ΆV� 	�)��L�8C���hX���4���`aOT 5H�����Ru�9����\�x�ܺ8t>l�HD�2f�Pg�;��Ɉea8�j�O�2z���G�L��P�î�8ӧ:vt�PP�Qu^��ᅣ'�,3��G��h����.DR)27�Y0$�	pW 0�b�ġ#�84[���A���ta�-��u�Uͅ�MP���/�Hb�b��XX�\ �d���i�H���!Ư��U����1IY��^w/:A�1���U	��T�U���02�0~�8m�����WPX�E�X �2�Gi��ia%�5�D��T%�B�#
c��3�,L'3��K���e*�0��4y�����柳e� B,�A�h��ʘHk�%SF ����0W�X0AE�ލR��i)�A�K��!3U��W2��8�yB�đU7�� UH�<��4���h��
?F��L�7�����ɋ���+� �2?��Mѯ����lږ��!�Y�i!�P�a֐;�#D,�zL�op6�!�H>	�/�r3�5���	0Cb�ǕR���P�c_�
<�)�A��@�2ZS"�=UU�6�Αf\1T�"3+`���%�i1�y�!FE�.9
��V*<VA���Opta�n��P��!3��K�.��l��gO�$UΜ��~���?}�X07E�)p��re�JP"��GOvX�����1�)��Zl9>u ��<i��.���) �H7�.<���2�Z��p��qOba�'�F"�$IFĈ�r	�	Z�V|4,�IT�ȒfA��a7�\" �lu�cBE'�)�$ɘt�b���{9����R2 �V�"G�E���鲱I^�m�0{��)v�Vh�x�9�a��x��q��F()�`'�"��Ѹ�N�L�z��7��&�=�Qn��U�o�y$�\j�g�o�(Q����(T.Hh���+'�\��Ʉ'��JABL�n�$���S]�Yh�Eͺ@�=�4�	�S$m�u`&]��S�j� I!���\�MH��:@�%¤�Ȋ	X0IIa�Bfn~hIa�;��ԑ��XZ�'*��YA�ަ���B��t7�u�-��4((M���JΤ�c���u��	��L�/>lm�����H/_� X�r�W�Oİ�#a@�N��ɣ��ǡ/&�}
�:�U&�x"j�;�]�1�'�|��۵%��-�ñi3l�7�\9fhT�Ap��^˴�@K�{޵#F� �����;lO@ɻs%�4 ��Z�8&@<;V�ĈQ�0��ٱ��ձ�� ����05MC�_� j����&hG6X�-�"�&c� `�'�÷��#`�� Y��K�x � �Ra�0~��<�*ϐg\���g��O�ӧ�~"7o �^�NG87�Z��'(Q�P�(Т��&L���D�x:�+�H\�U��Т�ЖDBE��"��mS��ZBaQ��y9 �3�<�X�P��Y�?�A��Y#Fd��$AR`�H�X��,L�nVLh�E�" ��ȗn��|�FeA&qa}"e[�R����L�'��U��e˧�y�Fo�BUi��M���]�y��*
θ�t#L��uRC��y�m?8|qtȇ�T^B��q�˦�yr�V>�lat��U�L%���P5�yb΅&^��#�n�>p0�s.��y���dk�s��O:x�bLP�ё�yҌ
m�J p��T,��)��y�0*w� �q	�.q���5��y�׶s�e��閟rZl,	U$V0�y"�B`�����׬ftp�J2�yē�m�~�A�-T�vD$"@��yr#�N��Xv��80��ԉ��:�y�Q�C�"1R4��*,�)������y�BO�\O�q��(�u�����+���y"i� |�	0��гa����!^�yb㏉]�N)yp#�c`x�����>�y�NL6!qN��#�9}�q' _-�y�@=4Ɇ��v	�<�`�1�����y����v�܌i��
�{)z�i�m��y¨���$��͞j;!G�ǧ�y2%64�L�X���o��Q� �,�yB�1
��d���5v�\Y{��R�y����G�a"m�)F��y3�iX��yrFN�!ǘ�b�V�E���H֠G��y�H�C@̩�E�L/*M�`�u%I�yB�W�3Вt��Z;S���� �'�Py����E���aY�=o�(b%�G�<ADjK�T���A�����Q��Nf�<�6��7WZV,�N	�A ��f�<i�߭y�u(1�>���:�A�c�<qҠ�-��� �	�n����Z�<"��^�N��Sϗ�^2dY
R �y�<� ,�R��ț`4���ū���q�"O������X�ؒ�K:>�mx"OL�y��
�|4��#��3)�)��"O�)0��Х'6����C?u�e�"O.��U'5:�4d�	B`�|L�0"O��,�9�Su"R�(�Z��"O��Y3�0݈ԡ6B
;#�X"O�Q(7��U�$��aA�1�>D�"Ol��k��NDY�F�Aײ�:�"O�wɌ%p5�hE&�Y���ї"O�����ğU4A���l���;�"O �RaJ�� $9�X*�1��"O0��%(Ŷ�VX;0X8qa�	�b]�`RA�@�`�qOQ>	�P!V'u�x�S��v�}��
8D��H�G�J޾x�ˍ�>(�����"}�k�~V�ie��E���Ç�!+e�@xv ��4���@'�OL}�c��<�r��!�@]�����z]vi�R��0�B��D�	Q`����*J��R�C�6xў| A�{���
��;��O���iP�H�b�	S=8�U!�'?0 �G]�6d�� ��z��1bv���nB$:~� �"~�Oɻ$�V����ŋ@�`{玄<�y��0�x|�ρ	kjjȖ�����7[���6�W�i��LȨ����;�I�Y���
����uaB�*�O	â��|lA��F'&�J�<*�m���qcz�YRb �O��	%m��A$<�"@��^WP	7��8@S��e��`1�%��o��H{3Hk��b�ԡ�'U{!�d� a�Ƽ���G��i	 ��$@Z���4����� �>(	�$��u'��<5<($?	;�m�R:h-Iҋ��k�t���ܰ6��0��6�O����G�L�\�s��?< �@j����?���<�J��� ��rH�)R&xG�$�X則e�,i�Ơ:���!@�#z��d@8E��(� LS'MhJI��Ec�h�*6��#?�(<��\\VP9v�-�yrh��Ha���z6`��HўA@�ɎXP�����W%!N:�n@X9�#=����+YHH0U���$�� 7 �,�|ܺb%-0?zy9�h�� �J�q�����
��W�y��e��5��ώ�2;|qEzҠ���A����,��-)�@��?�q���]��ȀO\��6�3)<���D�i=��3�4��9H��bX�Y� ̛|)P|ɥ�0.FLa��V	Ȱ��{D �U��-��i@��\��8��GD"]��R���Z��U�Ӻ�� �e�z�D<Eo�<>M�ŭW  ���BgYd���I�Z�a~2&�-i-d�*`�1N,d��KV�[���$�0gŪ�T��&�b�2�%��Mc�fl�1O�nǯ[�^HQ�R�"ˌ�v̓?1fl1��*�$L+�	]~&�>�0#�`�!m�O�)ɷ`�
<|��aMV�T�V�R��@��[mT�z�z�+ũT�.�9�!:#�\���M�-V�Q���ǟ�kQ�	��'�/
��`�<I6(��y�:�I�U���#��˱G��˕!��TeXj�	�\4�)!�ZP	�`�8A ��%�R�8 aٗE5�OXE��SM\X��E�38K��w�'�>�	P�D�oPn�3�� |TY�qL�GJlmZbx��+�?������9�<�H�`��5�TX;b(*D��H�kQ:�.��q�^�`��(�ff�	����S	Y����2mg��P�;�,����e����fi����:~��4�[2d4� �5�O<�P*�> ��(R�ܾ+(���DL�� {�ڲ@"*����J΀=J�gߨ(�`�b�?)/Q�,�B-R�$�>�C���pdʩ��`*�V�]R��y�Hyc�;0�`	����<��si�4I��t��II,c���A�Z)5�J]�d�'�M ����s����K�`��E��'��eG�0#��*�)X��yh˝�w��<K�NK-a���#; �jG��+@@6��f���x�|��%U��C�"V�B��i�+<(�x"�]?2l��j�n�D��3`B����F�+S#z@��bUv�ݐN��(�w�`���Y��;�O� ���lA4Iw�_$#�\qa��,�Ν��nc�E""*@Ũb��U`��F�ߤ��O���g�/����7A�v���A�M��1O��a��̮xl�r˜�}~�*׉�2����A�٫[&�̻%�
]2uX��j����Ţ���0?iѼI۶�X�(y.1;�1��S35ٲI�l�d����B~*#Sm[4`��0��ҍ(9�陛oц*]`-�B�s���Ąs�ay�KDV2�8��X�����w~�i*Q���T�� F陑E&�QI���%�2�U�ρ`��QD2��}�.��R�� f��Q}b*� �g�%z]�%�$g����J���{��;D�R��?}��r�6�)�JE95
 �მiZ!���Aw\��БG�.��ӖhG�8�lĹa` }�mQCrT���))��򢡆�L��h��i�7E"��B�/-n�	,N�!�0I���|m��O���N�4�x�C5� �;@c0�A��� G�>hhC�P:6dʓF����M`�矠ð�=��m9E+��+�|��gD�Ա��}�n�:c��Mb��?q�w�^b���S�#��y�? ]�B�΃v��0nܻnN$��iP%-�$PW@�����N��Q�n��ر3g�&t�<���'*�x��T@9r���K��K�[��u�rj��I8�#)�>$y���}>���B8p���2�J�_��i�2�8r`j���*K�c�LI��MӇo�T�_�l�����%	Ҿ�@7��w{Za��k�<i�ͅ��u�mHؘ!EG���2�O�M�C"A�0�� �҃�Vš�/�>#���'<,p���' G(��P/�?zͨ��ğ.�LbЄC,�\���욠;J�1��� 'E*�S=g���� x(%x�Rl�n� �8v|y�b��v�0	�V��Z�{�W)\ (wKRm���~R+�n#�*3Y��4}�p�C�|@\�ö�"4��Y�R5}.��w$�8i �*#�7�,A���~B���Ka>m�FF' ���k ��D��DӴio�Dj�H�<��(�'��ȹT��|�9� ��y��|�6�	$�Ru t�\�~:بkp��n�ıb���D���'c�;�X��Y?"&�F=`�	P��5K�N(���ę�ȀC��5	�43��Yg~"�F�iZMp�BʱK�L�@sbט2a�6PC�03Ÿ�·�*Zm��K�*5�s��
�zT���F^��,|����6�b�)\g���5^w�B�b�폢�<K5fD�"�ؼ9*�-c��z!��1VaB��o͙��ӧ`�̜0���5BJ��e,I<��E`r��]��|zE#Q>c ���؆"ob5�u�'5�� ������ɽ�F ��T�"��щ	$�m�F� ���x�m��8�80B�7l�\)@ѫ�R�&��A� ��'Z�dE���Λ: t�FO�8~ A�M!���� ֢i�n*I<��A-G���4��'��Ś��Ǯ��B�Q5φ�%A�)1�p�� �K�/}[p�غSp�:C��ƪ��b��ǒ�s��ƫ6�t��P�Ԓ�&!h��6��ɉ5�'(h�'�����֧)lD9a��w��i'?)Y�J^��v��AD����7�A�JG�����\^��iK
|\Xۄd߾�v��u��@����GA7KE��&_$��5!��j����.P�@�I�%�\�\�V�٩a^��*�ޟ����J��Z)�RFרt��(Ѳl��Us����7,0�J=r��]1��ʽe�la��`B�R��c�Us���mֶ��I</��H�I�J��!H��#���:w�Υx�u��ۃu�I�KJ.v.�H�'	�K��=pw@��!���"${��ŉG�R�4���P.��^�IBO�{>!����()�>QBCG�1��K�JK�	��B�Zx�#"Ƃy�qZ�ɊI`�ͣ0�F�8'd ��.�'5\����F��^l���"ǀ}�Uc��
Im�����K"L�$�S�L5����e���l�j�R����rU[����l��$�&�)���%��9uW68�( 0f��X��WG˺�Q�Cִ9�,4H�bE�Q1j�P���T>lYӃ�Áa%D�I����FȲ�a���NuNY1�ՙ'�|)����7IPd����6�@�)���3k+�Xä1�JUs�T�!�`�&�H�NLD��΍cd��*��6D� u!f ��+���3�j%��jZ�k��<c��͖pdV3j��O��8ffώTn)��k�3�R7�!L���,=�U��We,���7Ǒ%M{l�Вk�Xr�Y6�yt]��G	)�Z���L�3�t|�D�[>���J[�D �,G7PO�'Y�P,3���m/�q���' ���D�U�92���Y':��@" �X�KT)�C�ڝ4�M�'�$-U�Ϗor��+�))8�,rF�̽=�T�#�%-[$�s������8J_�h�W �/���٩r�֠��d�D��c�D�9An�9L��E�G��3i�.��3	������H6{Z,-�&��
?�R�i�.�;H��U�e��m�:�ȳI���#���O����)�8����@�6qș�$(�t��ܹҮ�-�����&D�X��DG�uh�U��0�aؓ���3��#U	�o˲����;�p���#X�W��ة�J�5�I�3-'�.\��j�Ю`��E
y��xQ7�A�m�����˗y�H��wK�taP���ӨH�W�e��CE����'\�6����Ꮑg�YYRO�) K�8Aً��>A�"�=�qz�ɼ2�� L�`��Q�-�;)�T��&F(��� fj�dܘ�Ӓ��jn(��d��0v-�9-�D��V�+���(6�$$��q���%�lA@U	��h��'=*բ�jҽ������6��I����m�Sh8Z-�q�@t��)Y�PS�NHl0J��V�D"����L�P�􉖣�25v�	T�ȨZ�|;5�i:\!˖�N�a.r$pb`��x����aO�?n��D���%<��gk

�駟hb5�i)t����[ >� �� nJ�zkT,�c�+�Q��$�G�� 86	�A@�0����N�`L ؈y�.@��` `䌌J*�dFI	�^9<�1(��D������`�����3�pX��N �HC�I�Z1(�h�b�0H��S�D�K�O�*U��3�aM�W����ļu�qO�zD"���[�ʓ�v�8P�G�0h��#�@�����ư>�pc՝bl ��]�2�8�c��6\�	F�ᦝ�U&�x���
���7��hύ����w�=D�`��T=	bi2ħ ��؁�,ܗJ�X�� W�Ay� @ˏ���I�$ȕ�?fm2��� ��Ĺ��|ޭ�0M_%�l�:�j!FFh5�=�Oҥ�pퟴ6#FX��H�#_VDm���W6\�|�$n�p-����/Kza�E��54&Jx�F(֠Z\VM%�􊀁�4e�ޭ*Sm�e|Y��3O�!K��h�� �X���u���X�ZD锗f�>��&��!�c�E(G�^Q1�N��U`B0��i1<OF�S@J��E� j5Łeb��!�x�J
�.���i��r\������E����7~�@��݃SԌ��)۵zd�qU��2�4��aOx`�ǡ�!dX0�i_��0hֈ��~��C↔�����q�A�a�bT�g��8#g\�'�)�;0���PŜ:3��)��
����tS�AOܓRY>�?-qjK�0��E�nL��鍢j�`�  U��f �48���&@͐!@2�%\�m
d�c� n�'�d�u͡n:��WAK�Y0�c	�Y��c@}yB ��d�[��A�C�q�x��.&b��qǇ"^����5�ԤzY�I�2�֨n �5��;X�@E�O��T�Ru�敪to���y�m�;7<8DX!��a8X�t�;��S�#DPf�C�MQ6 �Cm��4:0PhQ b6x���8��c��˪C�����'Vs��H�n����	 1��@�Hpz�mAU�5ڧAiڝr*R2��RG�G\q9�f]�"�&%�hA.s˜u�1DBn֍3r�R3��b�XFX}��9+Y�:�%��:ͺP�������@[j�a�'�~HP*�*[��O�(L�Q  �?yq���-`��-�Į�8�>t��L�5���:F���H�F��@L&\��9��-a��=�������[���e`Ё6�H���TM\���c\T9 ���
�DI�āՙ<8��U`�7�|����6eXUf�r}^!�#�2g���t�|"����Ó�i1L#&�H�L��m��(�d�݋��7�nX�b��c�� �Y�Ũ^R0�Jdm��nP�aL����/B�>�!H�[�
����_]"���C� �j\�5�ƔIؤ 3C4:=�Q�9V�&�hD$�J~��F�p�fa:(I�DR6�纣��*^�Z(��ŧ���BCM�=Rh�
g܉R� ����ê6��`��F+2{̙l� 6� Ph��Z�h|�� ņ�;�D)P�I��P��!(�2���lv�C�c�6Wg�4Ң�Ӯkʆ�i����2>lq[%�	 *�6�����t�{�c�Tf�4��*��Fs�L{�!W�)&�	� 1.��)��I6bdͱ�#�R�ɰ.��sBl�:9 ���'Ȇ5�$d�� 9&�x��c��>u�hh��;��K"l�:��Ӈ�1�0L郊:'�b5"�Áq� h&��^�(�ڀ� �8J���'đ�0!�`�ˠ*���p�� !|h�m��k|�,b�&�~��=jb��f�$!���� a��G��$ zmӱnw�4Z���2z��"m���i3j�����˦��e�晹��ΔK��ڃ�W�#MF4X6��Z��T�� /;���:W�.H�����\�N�R�Fψ�qb���D��?d����Do���j׆�L�쉻3�]�K�F ���.wo,�i��E�y�-ʒ�Ƅ#3�r��C�C�L��7�Q",	lH�^#2�	�{�	�" �'>�=�;tq�7FG1�L��l�j��y��$L�~cj #��I�]ž�&(�[K���GF�3�x�E�|R�c|�� v	�B���{!Ń:l��[6'�`�ƈlڿv$�T8wM�r��4��LS����w�˄s�J�+�,n�d��m�+Tl���.��lp�GO�/�VQ��Ň�=�da�<�⥇=?�h}�F&�p�nڣ<�V�I�Lگ?sִb�@�m0��s��3Ǹق��(��c
�9�J6�X4]~�a ��3�vtQ�GS��(���׽$eʠq��J^��$��a��J�\����K ��?Ar&L�tR�ܱu���4�F_���M�V"B-]v�x4C_[`�	� ���h$8��RE�F1�e�%&����e�&���,^|�8��]k�!qdk��HR��iՊH�*��a��F����
\?Ae�x�D�5%�%+W�"�Č�P�Ĉ7-�Z^rĐen��e�~��栏�C$���n��Z���c&LF�o
��Ģ��7�\�����?c�j��� (�d��	&M���pĭͰ �h��B'�h�$��C�� S��F}+�`*���$K���d�L1�j�7=(4�)�"��*kB���:D�H�����*/���T��p=A��]�
��7Kق�x&�V]�T��@ѿ_�a��M�c
~���(��CA�Z4Oѐ� ���[�J�����.ވiׁ��N%LE� [�7"���Ԅ���Ac�<.܎͠! Uh�2�Ѐ6}*�4��L��o��Q�!(CCOuH��� �j���*ū� 7x&<���Ս^���Ɏ9 l�0�$i�'L@�&ʓzd����n��(y�钥|J�0��A�=�2�i�cV)E/�窌�<R�kR�1<`�J���#p���Q�H���2�PcC�+@%�("�*,�I�X�@0K�#݉T�� 	�+hF�O��06i�	kB́��E8څpuf��49�p��p���v�����H�a~8�14/ǜ�H�)��Zi����'᪕�b�ƻC*�1p	R�.��m!3���~b�A�J��i	��˘r��\�sc� ���tɛPȼ�G�ƨ$�!4P�hW,@�0 ��Q"OV�c���^���8cK�*b�z���4�v�����2�^��b���{�.'�De��^����0~�&'�E�`���DwbC㉯"%�<��B2Жp�f)H5G��������dD�ɥ!�����	?�:ᩰ�s7R@�5����	Y
;�����!6�hJ.OP�� oD�F��@ФM�`8�d�-�B�{�kI�Ͱ>i7oW�\:~!�ԁ�3׶ ��gFz�<��kA�dj�	j1B���u���t�<q$�R�N�E+Ԏ�C�G�r�<�F�V/0(��A�مh�����f�<�;ka�>V���� ������'�8��3lS�Y��pI�q��Q��'(* ��'R;D�;�c�Pq8�8�'�$yB�O]�Rf���?}����'À9�#�=l��I��O��h<b�'6�1��P�~��ip�E߾1|x�
�'V������ Nn-��qR���
�'�ecA���`i9)�21�X]�'��4���ܟ#;|�	���,x�eX�'28�3cf)k�݋�e�3��Z
�'�rɻe�C8&29��n�/4R8:	�'�9�4��*���O�*��ȓ�'h*��f��L]B�A�;&�p�{�'�:u�"FՅb�����,H���b
�'zRe`��9cʌA�a&�&
�'�|�!�8ŢY���y���'Y�� M��!'�t�3��:�TU�	�'m���vJZ0 뒡
$IH��¼9
�'�&� ����%9Z	D�1P�ܢ�'�ny��f]y��8�( ?����'�-�cKL�?����p怑Ql�d�Ǔ1����GD��'A�Av
̫&� �uh��E=�䎙d�¸bb�I�X��)��U�f�X#mQ!e�Y�����R���QUH
5���OB���'��l8�-Ǝ^�,Ebf�)zQ:�����?�%���y��[>5�W��&!� Ie�Q(1X<����K#�xi�*��<+O1���� �!f"�0�����S�B��8��Θb'�c�<���O�������0`�Ɓ�L���d�R�L��İ�'<�@�C���E��|P�!ß?zͤO����)��%~�h��.��$ᣧ�'�,�	3��=E�4��#'�� �te΢0` |3��;�y��GO?���K.K/R�*� }l��� �Y�'�G��,�>T��@�c�%�j�ۧl����S�x�o�4;8��}�O|�cA�0�6���nF_( ���z��PvG[N�i>�~���E�N�H�Dn:��ckw}b�Z?�L>E���ֿe�R�ȥ/�5IV��aX��M�L��t'�"� D� /�F�[�S���Y���~"�|b�/�ٛ�O�����.����A�$0(l���O��Y�')�O|dM|
VD��%)���a$'\��Uo��`D&�P���!H������o	�S5�EꡨF�e$������=�41E�i<�ɦVoa���r���
���jlv:@�7m.?��Y�䉈��@/�ReP��
0?���*���a��`��0�0|��nG�fpf�3smF�t���A�)��,�t�cG�<�&�&4�a��mB�QxЋ"��,*vT|��.G�$�$0�'���Y�E�:Ȑ�IԄ��L���g�b���%��R�T��,�{4�"ֱi�&�B*�
sY�!q	�'51
�x�h-1A�� &M��wfPa��?���fI!|���$JZ�r��@'V�Z��Q�N�2�#��g�zD���2Lp�2Qv(�a�	s�*D�ȓG�� �����؜�bK\H���~�����F5IpX܉�mZS�B̆ȓ}��G�ɭ%��,R���7i�e��M,FDR"�ѡ����$�� P݇ȓZ��J􀎼_��XS,P�`'�(��ֶ`ku�X�{.~�:��M����ȓ0�"�8䩆�K=hгa��P��0�]��R,Sr�5����3Ǧ�������֫J�e.*�j�:a0���W�D�F٤?��D��B-�M�ȓQ��9"�ƙu,m+�ʐ \'*��ȓ|9�� g헮��Y#��ޕsڜ4�ȓu�<y2lL9H��eGM��(�ȓ���b�%n��@#��l�l�ȓysܳpDݮKC�D0�ȁ�~�����g N))��G2���ˤBn��-�ȓeiZAX�Ì�P(`�M�%���ȓa�BQ�"cO>@	�Lp�K�^vT������fI-8R0��&��Bx)�ȓ�z�d��K;�5;��]9�̄�.nv�UZ��d�q`�,!�����o?0 B�D�X�T��v�G.�����X����B#�?�,��ƀi`�]��Ŷ�8�^q�qkR� �w��Ňȓidx��J�`�ڝ�1��9:f]��(�z�У�ʢef��b
#f-�ȓM��
6cߌ*��*�h�8����K�$���_s7�A��O�M�h�ȓ<0�U��Ŕ2�����E���i��j�0l��=0 0��$qF^م�8�(���e�L����A��N6<Ņ�.�2xz�ȓ3*����O ]�Z��j\���@�D:1����T,��ȓA�tHS�^�.�2����Hqȇ�\D�i��K�d���-o{���ȓ9�X'���JקLH�(¦;D��1'O;sl� C�жgP<J�;D�()�	������C��w)���S:D�H�c��7�α�'�R�vUr7'8D���Gm_��@u��ŝ��l�A�7D�LQ���"B&�x��]1
q!��*D�� zxr#��\�����r2���"O �cbb��A~(�ˤ�NYZL��"O��ӓc��Zf5��e��8H�ܙ�"O�Eڇ�9���Iˣ'4b�	�"OX��p�+:���6NC�8JF"O�����2D��"d�>W��A0"O8d�R�[sXp�U�([Ҁ���"O���5�I�^]n����9�����"OP��C�؛i&p�T�ޗr[X삄"O"�z��{�ЩRA��_g�Z�"Ol��#�J�:>T9Ĉ	S`�L+�"O�x�,3?�Ȱ�&[	���R"O���ʉo�h��Y��(�"Oĵb�AG�7�X��G��X$����"OL�xt��/2��D�ڼJmvx��"O�CF��-J�Q��aP�LB���"O2�����c�|Yp�F�`""OX�c�c��4Ux;w��9y��"ORu�e)�zd���a	/r��b"O���D`C0}͂ҧH�C�"O�����jV6X��%��L(T�@�"OP$�e|(�Zg��y�x]R"O��a��
���d��L�|U�F"O����a�ĩ䁍<2�4� D"O9�a�:+XB�is �#��I�"O�Pze�͡&�R�+Ġ��7�RI�"Oz����3����{�QXP"OR5�g��mB"i�?���)�"O�%P���~�\�CǈNČ�9�"O�1ɗ��7��9Z�Q ��Җ"O�� ��O�褭s�F41��²"O��gGP+po$Z�F�e�C�"O�t(�b3b��J�:�y�"O��Q����\�fhDH�e"O0�4ةJda2P)ˇ��
�"O(�Ҡ�[°�S(1!{$źE"Od���c��|Đ '��5��ZU"O���PF�.���թ(�ڸ!"O��pg1��A�M~���"O�x�@e���G���pv�z5"Oj K���^W���5�=3fp��"OR�5��+E�x@ˊ�4I��p�"O�ljUz���S5IE="�RA"O,��PBQ�:�� �I�P��Q��"O��QӢҐ:]T�2���Y�"O��C!Fmc��Ծc�ډX�"O~c��	0���HR��+H���(�"Ot���
�.�����]�t2u"O���'�&C�⩘��D|�@�� "O�5�n	+F�8U�R��1J����Q"O�ѳֈ\�ae"t��ӸX�$���"OP�����}\zLi'�1�>Y�"O�d"�JЍm�(�����r��i��"O�-��H�2n����GkU#Y?Yr0"Ỏ��e��<�4�\P/潨$"O2�hd��Y|����F>a�(EJ�"O��#�Cv��]n%J�x�x�"O� �g��5�X���޶q�)S"O8P�O͗k��9�7k�:Kj�c�"O�=��%JQ�iY�)�86C.BU"O�$K�'��CV��r�a� T��K&"O�亅O�Z�,�+������ �"O�9 ��ӄ!����S9��"Oj)+r/�vt���V�o�z}�a"O� �T�u�U2A���a	�/C��DB�"O\��$@�6 ��
�g^�Ia�"Od�$	W�Ԁ@�R�q���+�"O|���舚�2�#��N�"�� ��"O(��#��%6vt�p'Tj���c�"O=a�aV-���8�����dBF"O~UI!�h��%�f(ܑ[r|�G"O��Dd ��a2E��2��"O�D�@�7>rJ�3��0Hՠ�"O>�;jD��ⱻ+�"�Rx��"OnP�2@�=x�f���I��u�8Pjp"O���R�̋�$��ϛ��i�E"O�\6�A�h�°)�Η�| �'"O�"�@��%����ț�~�X��"O�ѳ��P3W��p�fN`!Ç7*!�d`ajU:wAⰁ2�5n���"O�1������$�H�SS��B�'���Z,18��,#A��-�����'���G�³N�P�E�V�Y>^�3�'`�Q�3 Ɉ�`I��m֎S��'V.m�� }`v����ԬP�8��
�'�PT(�ʋwn��r�ڈ]�:��'w�9�b*�%P$lp
G&[�L @�'�VPP�>\�<� �I�R�8�;�'�p[�\6N�^=!�Ǻ嶭��'��Hk�FN2{�.䣵�Ŝ���'�I��z.���ćޖ��'�\9���ڂan�z��X+"O��ÓI�1;�tT�-IJ&�	1"O�ܲ�(Ș��qr�D3.FJQ("OL��H�7)Wj�xq�.Y20h�"O�T�B0KV�RN<7 �C�"O4I�7�Z�)�	Ak�/s`ma�"O�0H���%Z<�Ö�L%+U�YA7"OҘ��m c[X� ���726�e�e"O�e[0o��M���A,�>"9L �"O��!�b�_�ͩ��X3p8luA�"O�,�u��Mߒ��&�K�z��M2�"O|�����'�@����]�V�-�"O��ʅ�+Q�x�M��z�aD"O�tr3���$tT
��������"Op�1�E>v����g͖wq��K"O�\#E�Ӂs��]Xg��&��� U"O�m��Nݝ��|�⩃�d��1��"OH9k�ñ8D0��S�$8%"O�a�J�Q��u�3�T�S�~�h�"Oҁ��U�aZ`Q2Ӡ�"���q3"O8���ꉼ`MX���Z%=��bV"Oʅ��`�=���YP"?<P�`E"O.u� u������֕X!6:�"O�- ��K�m��y@�*b
	S�"OR0����-��!�q��1/���C"O
�b@ȩ[��K�/�9!Խj�"O�훱�������H�s2�)�"O����$DE4g��N؅�"Oʜ�vH�&fPh�&��M�ލ�5"O�XHe)���r`�w�T��"O��P$j׮{c�
b�O6}�T��"O����Œ.���#�LU�6�d�C"O(!��!%%|�P� �B�y�|QY�"O t�d��xmB1;�ׅ;�T���"O�`#�&]
c#��m~��s�"Ov�Wm��5ȸQ�c�5�L!A"O ���U"U��9��m
A%Z�{V"O� P�i'W�M9<��\�\�LF"O2 0Ɨ�r[�M�"ˏ18��"Ob���Mu����i֋C6�xzB"Ol�BS�����x$����"O*p��% ���F��UR���"O~9��
�k�cË��_�&���"O�]KĂO�m�R@�T�6j�@��"O��z3l�h���~�ؐYS"O��i ���KzQ��.*UǊ�٤"O���
nf��OL�zD�"OT�	֊�(s@]�҉ϋ{�>�"O\��6S����*�Xi�<��"O�u���%�A ��c�-
�"O�����������87:)+�"O� A�áT�	��
��"O9w�ܡ7�p�g�("O@�:`f��}�h�@ӥ�5 818�"O�,��m�6�@��
D�v�"�"O�|J�e��,�/ƺ5�p�"O����7Cs���Zˈ�	�"O���63J�I��\5r����"O�<J��Jڞ-��H�5�J�@�"O���Orp��"s�����"O�l	%莐��\��R�\�ܹ�"O��   ��     �  Z     ^+  V7  KB  �L  jW  �`  aj  Jr  "}  �  	�  x�  �  U�  ��  ܯ  �  a�  ��  ��  +�  o�  ��  ��  8�  |�  ��  �  � � � �' `0 X@ �L uT �Z �` !e  Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�� |d��"O
`�(�;���8���-0��1%"Oj4��ND^[��"3/9�0|H�"OB���H��*�ʞRy=a"O�味V�!X��!&F�:J�$���"O,��a
���C�Ą�M�"O,$3%o�-���p���+Ն�:1"O��ݢ1����`���y14]2��i�<�6��{_���c�H�`�fX�$Kn�<��A̼VI�xR[�)�Ć�pඤ�ȓA5��('nߡ4�� �)˩%� ���,��r�؊b#`T�eT09���ȓ!�b��g��}�8�F��-? �ȓ
K|m�ș�VṔ���2�%�ȓ"R�X�j�4JN�1�˘X�i����̹	_�jZ��1!g��zܶ��ȓgil,*�J�
j�Ne��i�J%b���f	�(U��:���G��$Y^م�~r�� S�%T"���k\�jx�ȓ|4�1�îJb��@ӵ�ݩn�V��/[`�"�v4�R�!ʎ<��M�ȓ`:��z�ؚh�J�Z��$HY:	��H��p�m�C1��!��B:��0��EnjZA V;9����J[
2���	��4'J�EA�IVW&��~�(aZ��ӹ�>� o�Y�|�ȓ�f�A�
Ο7�H��M�$�����mޠP����/���ANXo*�ȓTv�����{ ��-7�*h��I��sB�8�8���3����ȓNe*M�悡;������X�o��!�ȓ'lj�#F�m�+R&;�|��2)n�C��0S4���T:
b���:�0!��e֊��)��ͷV��,�ȓ0�&�8#���� ع�L�����;�P�AFd���,w�6d��r�EQ�( �gVlɦ�M,H��,DP���|�I	$G#\���ȓ"�)���E�B	yt&B�^�LɅ�4�� ��eëF�ڙ��n��R�p�ȓp`@}bŇ�=�$�AUN��P����L��p���_�a�)�Y�!��-��u�5���o}�`iF�@A�p ��F�\�0��[���IF/5���k>bTؖ�;K'DT`�^��@���)��x#!�|^lz���6T��jC�:D�$�"����!"�g��p�D!���;D�p���Iu�4Tѣʇ.E�(}�!�$D��!��pζ�`v�G�� 50�&&D� �dP]&�1� �� 5�Ɯ�f?D��0#ҶEbybÊ�
"ܮ\�@�)D��9g����^���H
'kF� 2�(D��2�OhL*uY��0!�/�&*C�	8�$jM����Ph�6�>˓�hOQ>=%�N�~ b���
9� M�r�3LO���i�b�f�qG	?V�ȱ!Я&D�0��A�0i�~����������$�d=�Sܧq��y!⯝0a5�8 ���9��X�'��~�[=\e����� �J�J2Ð�<�O<)�O�OaʓRVq��ɨ<!0��F�b�ȓo��!B*.�"ܡ� ? �	تOXqIM<���4�F ���T%y��y����?����'^�)� �= �O�bش�RaE[�%�A�"O�#aei����/��6���V��D{��i��s�Z}@r/��t���׹
!��r��u�|�,�n�4w������Dx��	�Rr��D��z-Bv`��زC�	���� .���(�EQ:���S4:������dהg�0�H�94�!�"O�ۄ`��6Gzl���^:]%T�9V�',��Fy��	��$���I��ޖ_~
qEᗽ��?y��	ߙh��<R'8~ 0r�jɹ9�	sx��H�*^��v���EQ>]�(U��xъ����"y�tE<��؂���h�C䉠S^���"&3ҀXE��k�'/a}��^�Jv�r�▦4b�q8��2�y�� N
�2�<]�<b��&�y�ּC4U��+J�pxC�߁�yR��O!��ʱ�B�udh���^M���Y�N��"�_�x�X�!��A��!�dSe�``1p���?��U����=%�!����`);Į��d�[�ARBe!�F^|���./N�4�ªE�!�D��b��=�@K='����D�8"�!�dC�D0 ��֗d�x�&�K+H�!�D+v�1FM�T��!�Hm�!��	Op,6�����#r�[�9�!�E+����� <kp� �
R�!�d=e��[�C��G��f	�Q!�䐴.�9����_+�Yx��X^�!��3��Cd'�v>�)�̒��!�$ή˂)�<U7�Q�A
�C�!�{�d��v,�<`��R(I'`s�O�m2ĦI9*. d��f��u �����s}����!�D�B�Y}T�چ��>�!�$P]"�,S�)�#Gd�;��J�2.�'B�Dn�j���O��V�\
pY̴jb���QD�	�'��i�M�����jA���H��Y��D}X���adϵ�����!*:b�i�!D��"���$2��`Kq�¡�V�s@>D��Yc÷&Ez��LXȂ�� '>D����6*Tx$��
��8U;D�(�C WP�� ��۶p4�h��8D���&ʇI��%Av�zH�+D���'�J�\8�u���:l�:�`&��O��T��@�,�
\уgȮ=H�����$D�L��\K��:�l�D���W$D�����&ci�)Js��7�b�a׉ ��ȟ���p�װg3&h��LܮJ@y��"O�$�s-�
���3K��n)�d�O��=E�D�Z;2�  ���|�2�U�B��p<���Ʉ{HH�-�	-��aY��B]e�B䉎>���Fi̘����BK���'��"=�O�
ʓn�h���ņ�	(K��  J'2=��� ����-d����e��E|�R��D�$C��햭���ëS�l�xA����xҢ�(eF������Tv^�22�D?�O*0Gz���ֿyVN�[�mSy�1�qƒ��<Q��3������Q(C��ab�(n+F�X*�+�fL��!�7X�F�z!\�0T� $��z��)�����ڽ� 	y���_W�C䉿M�=��Þe��MR��H�P�f㟘sϓ	S��ךm��U˳ جA(^��ȓnpx�����x�2��Kܑ/q�\�ȓ-���:��u{�&�#Fl@e����M�&�_}���[�~�PF
�y
� ��p�l�>*�"���*��y�6�a��'�O��C�j�~�:}��S(�j	"Od��$��X	�L��B���"a"OT�r�fˑp�����HF�'0�e3t"O��#�Ѹ0v�$��/z�T��"O��Q��]�=�P�����1;τT�5"OV��ѡz�H٢
���h��"O��@Dҏ��\�d�b�P{�"OF�+b�ǂn6y��DS�'v|j�"O�)���J$"��͌T�XhG��?�S����?sx���[5\^�)G`�eA!򄆟w��pP��V�2�rǍ��( �Gy���P���W�.Q����:�����8D� �f�f1���i�%�BJ,D��⡍ߍ0f��P�W�MK�=۷&+�O�˓F$��J�A>2���F�4	�*���N�L"��J5?��%�!��E��C��?�Dy�#�:>��p��B�gh�Q�M�y"�_?<F��@�$�HAi�o>�y2-]�|'�x1�E[�M(:Uω��O"
��R+$��	�f�A�a7�F�<iES����Ŏ�VOxP)���<�pC�|��\A%Ɉf��4�p��|�<Q��6	�`j�.F+l8��f�T�'�Q?���X�vv�#�*G�Z�[�D(D���CߗZ�
��0`�eq��6͂B?�L��1ON���Q�m� ���]Hx)uO0(h���#/�q��1JyrOTX�P���R,�*�
�B(d�4���'�O��{�'�D*����2$��gד(cPm��'��Kg�P�<��t(ޔsg��2����B�Ow� �u�8UMh��n<m�Y��'V��2(.�Ԭɤ�V<cʆH�'�p5+�I��x��ղn��1J�'c����**|m���ؿa?.,(�'-.� ��GἝy��JSÔ�J�'��a�ٻz�D���<V�~�s
�'�@��C6z<���!,֨U*LЫ	�'iBt�An�$1f��a
C��
�	�'�H蚔�Ą}
֙(1��#rP��'��}��$Ϝ q�x /Փ
3��`�'W��Ia!�3z8�+q)��|� ��
�'2P�� R	/��R0��E`R�9	�'���!5�х:@`jW�TS�"Ѐ�'D����C�Y�Li�$+ך���'�2xb�GS�Ur�9�Vɍ-~��'�� �e���6��c�yNl �	�'	 ��H���B��B�E8u��Hx�'��(��g�;5�
b':gb���'��*�'�Xl�}Qa*�X��q��'����rP8δ�B�˿�����'<d+GD�L�r\�&� �rl��'�<f��7<��A�C�'���'>�)� Ɛ^6H�� �:y��'��R'\%-�Js�	�-iHո�'�z�KW!
K������!�B�(�'P�@"#�,gY�H8D���>��'-(����M95K�Aɤ�^w��
�'���E�<"z��飏��,�I��'���3V���3�n%2�&� 22�I�'�����޸L\|Pϖ.r�6�{�'9fKP��^2���JO%���p�'���3ENK<[`�I@� 1
n^�S�'r��R�㝐=��ݩb�	~k��� f��'N���^10/:%��"O�,*��8|@��U�>P�T"O�q��H��Lܐ��B���p!�"O���� �J@ʸC��׹�f]B�<�'OL�$��iX2���R�rq�Ɵ��Iʟ �	����	ʟ��������ԟ	'H�"� �x%��':�T��fD�����I������`�I����(�I��@Rc($[$ Z5��P�P�J����I���Iҟ��	���	ğ��	ៜ�q94u�6/2D�ٷM���	����؟P��ޟX���p�����0Aڋb��#�H�:'�� CX�t������	͟���ʟ��	����	����,�::��c-޹I�ިP�ޟ��Iߟ���˟���������l��̟|*�#U2s��HSKݺN	�DҦ�T��̟�����(��֟�����H����x	v��bnr+~����F�j=�Iȟ���쟤��������IΟ���	�F�h�#Ƿ
N�B��Q����	������p�	��	런�	˟�I�|��x��9��x��n"6�"��Iǟ�Iџ4��ȟ`�	� ������ɄK�@�QaM�#;C��;���*d����ҟ��	��	ɟ8�I��	蟤�IWC.�!c���h+ƱhA��� ҪX�	ߟ���͟,�I����Iٟ��	џp���H�
��7��T40K'�{^����������I�l�	���A�4�?9��:��V�t?�Z�6N\����Q����Ky���R�8ݴ9�t�c���j|*�ږ��$N���҂#�g~R�a�&�d+�dYF}�)g�N`�Ǌ�D|\�gi��옗�\֦��IJ��%l�L~2O�%F��sW�MP�)(n�Ȕ7��i}&���F�e�1O$�d�<)�����6�8m�&�c�̍�����Lo���b����¶�y��L~��lBv����6TГ���T��6�٦�̓���)��qL�7�b��ڡ�#��A�R�O#�|��#t��"���(�,���WP���4�'�8BG�ŷd��Z�ŝ(��`ß'%�W���Ms�Ez�� �A�j
,_1����M�2��t���Ž>A��i~`6�m���',�p���_��'��+�O�ģ®^�bj"<���Ѽg.���?+T�4􁲄��}F�J�c׶��$�<A�S��y��޿z~�I�)˨:.�P@D �yRfy�Beq��� �4����T��7<`����[�8����KE&�y�/vӴpo����/�I�'��m��L�$h�"�{��[�V��I(�@�c����Vc�;sV���KҘ`X�Q%�I<c)�ӷ��f�|=�@�O��4��a�1g'&!G�� �t��؉k��]Pu�lx����&F�j�P-��k� _�Ƞ)�Ƙ"G:�w�ӟG����	
�x@�A�N)A�:@�tg2I��z�ƣe��2���&@e6h;$]�Y�VL��ϒ,U�rآ养]Ψ�:��éy�ty�%*W,>(H��iτ1͘0;�V4Iފ5C� ���.����m�R53�,Z6'�(ZplĒ%���{g�S>U��Ճq(�9뢐"ueˇA�t*�`��P i�7l*JT��I�Ms���?����jU���ۖ�_>���Ԭin��k��{Ӑ���O��d�m�po�����?�����rᜂC3��h0+Vp�N�Y"�i�r�(��'NR�'H��O��Ix���Bb)���1*�J�&=�d�بT��6��_���������R)r�|��q�J#�|i����M{��?���m#4����?q)�t����,"�ߝ?��$�45"���Y����'�
�P@$��O���O����%`����S**=�[�K�z}���.U��My��'��'-(��u	�*�X�i�>� �>AB�	�2��'���'$R�'�2�ڮ7x����̪Mf��:e�ZgA~���'�"V����^��ݟ����_b9ہ��˒�Y�Ο(M-���4�b;w����	ğ���֟���Z�b��	b�,�(�9�\)h�睶GH�i��4��d�O��O��D�O`$�Щ̑9���%�0�(\2 i0$�c������O��D�O��D�OF��n�|���,J�i� 	�5�hY2�I�k�� ÷i,��|R�'-r�+}���RN<df�?��i3U���\�ӖI���U���0�'��I��?��O����bty�eB4ڬ�s�G*���6�i��IޟT���.�<"|�����s�|I�v��SR�����I�ϛfR���r����M{�\?]�	�?	S�O��h��>N�8A���ΚA�Pذ��iL��'g�	�!X��&�Xe#�Q[$IQ�N��:��M���v�BY{�*S��I� �I�?őL<�'�t)h�$J�q��)SdM
��ba�i����!^�<�I˟��3����|`r�
,	)��xT�J'�]�Q�C9�M3��?���5<@h��x�O*��'�$j�i-8~�
W!�J���G(�>���?�6�s��?���?�4��X�T��*[�w�~�X��*=�F�'CHi�v 8�4����O�˓X�)A�)
2�)bK���a0նi�E.��'���'2P�d�@� K0MhMȅg�����!ډ\�ʨ�L<��?A���d�O���\���K�B<�4C��U��pR#���O��D�Ol˓��$��9�ʍ�cBY�T��0�H-}�	 1X�d��՟`�IHy��'VB$١���Q�>��8��ŵٔ��1���O�I��IIy��'"T��Q>9�I�B9�Y��F46_
=1F��n���ܴ�?	�b�'���Y+���\ȶ�� W1�b	�;;Y2�m�� �'��H��/��㟘���?� �j�)դr��
h���F#ر��'C�.��rCX�h�y��� ���M�k����Bb�j=@PT�����'цD��ş��I͟��`yZwȀ�Z�bN#b�̛0�_T*���O�d]&&�<]���)�?AaDl�6�D2w%Li�&��'`1��C8J���'�r�'���_��S�
�ARK��v��pFO�6��albO��!�)§�?1A�	�96<(�mA]stIr��.x����'L"�'�
��^����L�I|?�"��,�̨��/,�ʍ{2��R-1O��@j�����	e?��&н.F�{�I�,,>}�&��	�ɿE�"M�'��'�2�Va36 ��oaEH��Q+�9X��	�]]��е%0?a��?�(Ob�ď��a���_�kb0br��#K�b�A�i�<����?�����'�Ri��u���h�mҚc���Ʌ�%C��g �0����O*��<��S*�O �C�쒧e������\�f�,Yڴ�?���?)���'͢�㵋ַ�M�p+[ F�d����eR�BuG�N}��'�R�`���)�e�O#�-@�q۞���n��mR��D�V��*6M�O���'��h)K<i�B�M��d�EC(.���j���ʦM��Yy��'��8rCQ>M�'[�T���^�:`q"��8$n<9#&|^Hb���'&ĝ����5"pn�!6~��i�"��D���R����(�z��	��4��ڟ���kyZw��=z��44x��&:J$���O�ʓ2�j�ExJ|�t�2S2 Řq%Y$�KV47�P�2=����OZ���O��ɸ<ͧ�?ɁL�+S �,�����}ʆ��,�����^#<�|
�u �uqQG��M����?]�8꠼i �'^�ͬ@�i>q���p��,�j��`ƪ-��8�g�)t ,15��?�ħ�?	���~��]�,s����-)�|�1)�=�M+�0њ3-O���O��6�3/HZ`
J84D��)B!�.O��s���������'�2��,#PX����3��Iߕ%Y��IT� �I���IT���~�c��J����cʳT&���#�Mk欖a~��'��_�8�I�K��=�'s�~�qw���zO�T"����~tm�͟��	ɟ\�?))O����i�+@2;0��@��
@�|@h�
�O}��'BP����նq�Oi/��!	ࠪ�ᚽn�N$�D"՛��mڟ �?I+OX`��x�܈?��ã�,
��M�tJ��M����D�O����N�|����?I���*�-��`R���n�`�H5���O��4K�	1O�Ӡ\�Bl���E�[�Hz�%Q�-���?Y�'
8�?���?����*O��J�JD�����. �*P��fS�F�	���*�Þ+KdDb�b?�z�IG25��!�kݵI�~I�SJs�QP&�O�d�OB�$�����|"�X:N�9 �Į;�ބ���S�#� ��i~�!��$���d��b� J%,Z[�wK�>/�]mZџ��I�:�)�sy�O�r�'���55c�ٲ�]xB��D�Ө=R��<A�� B��O.��'����&)_Fl�u�k~�	U��H��V�'�x��S�`��ԟ��IH�v2PA4��6 u�0`�׬vD��'�X��jޜ����O��D�<��"���Ǝ�u�,�v-��m�@������O�$�O:���I;��`��
�-e�z�i��U�Cba��d�	gR���?����O"��+�?���� ��)k��Q
��q v�p���O�D#�I��Zb�'Q7-
�4�KV�^�Đ#`�ǔA��������Sy��'�*���[>)��S���×0f�T�pd��h�ߴ�?y���'����F��ēZl�C���7^nJ-w�F��Xl֟Е'6�Ŏ�1������?y����1()8�T �=Rvb ���'��@�!Y8�[�y����1aHZ+X"�{�P.	�"<r�T���I�vGl��ȟ���ퟄ�TyZw�bt�VLY�nhp�z4bňD���#�O@�dP�s9������id�ݳ�MT�c�l�B
-U؛6�� |yr�'U��'G��V���Ꟙ #���g
!k,�[��_�>m��۴դ�ٓbZ^�S�O���"$1ѳr�]*��V���4�?����?A¦)��4�,�$�O���"�ؑ�vH�vK�%��R�TIFڍy�,�6O������O���/M0d�vg�z�Hs�	��\6��O4Y���<���?Q���'�6Ej@��\���`�JHA���O��T�ڄB������	`y��'-�4@2͝�����Z�dcq�����#��I�����ǟH�?��>>�	2�F�4�t4A��\�Jw�#煇�\Δ��'��'��I��$
`�YyRí��'�Ig�R�:b��������IH��?!7ɽ_*�lZ����;2��h'e�	{L���?�������O�Xh0#�|*��F��1�H��Yg&���e���T�iG2���O� 3T�_�O?�'|ց 卄,���b'P6�`�ݴ�?����?���:Jd�C6�iS�'\�O0@�X���.j���J�j�q�챹1kr����<��P�Χ�?A��0	&!�禑K�.�9f������,G��%C�ap�����OB���@����I��|�I�?���ΟLH���8D�$�P���Б[q�ĳ����Otu�6��O���<ͧ��S)��eI񁛉I�$d���]�>4�6 0K&�}o���H��ϟ���?Y������I�{�dK�e��UZ����gF���ڴT������D�(��)�O����O���Xr�? }c@�(7+♺͕w]����iR�'�"E�$%��6m�O ���Of��O�N��x����&O�A��hQth�	d���'��F�R�x����)��(�d�O��ʖh�,�f(:%)��~,��hSk[Ѧ��ɣ^h:���4�?q��?q��t��St?�K
�Խ�a&�>�Y�d�OO}b���y�\����ڟ��O~b�`H��¥B�;��@��g̪({f�dӺ���OR���O̝�O2�	�0p�E�.�֤ٳ�߻p�>�(�FY�L��۟��	h������	����U�X?�M�EC~���:BĨm�V��$d����'N��'���'�����g�n>�37�̹9 0IܐV�D,��+�M+��?a��?y��?�ׯK�U����'��.B)5������?X0�`K�!��6��Oz�$�O���?�Ei���ķ����/÷i��}�7�R��l(7�i�V���O����O|�r�e�ƦE����x���?�� ��$A���H˱R<>��բ�M�����O�2�����<�禡��O�L�s!�G:v�H���FdӸ���O>;1��a�	՟T���?��S֟��C���)��i5��E܅1!@������O>���<y(O��]�B���I�%Q)f8�+�0I��6B�])n���I����?-��ӟ0�I14,@��$�۲lQ��J��Nȭ��4}��-S���?�*O�I9�I�O�A��h��j�
�p!��D(��C�`ئ�I�<�	=,�4�?���?����?��X�4�U.�:[&��ˠ �J&B)m�ԟ��'Ĩ�ᙧ���O��d�?i�ǌ+[c�T#�X5x�r�8"ݛV�'�hmX��x���D�O����O��OM�$�7}|Iq�'ٕ���x��d��I�P��	Jy�':B�')��'��0�㖗^��z4 ȦI�n(� ��4�h7��O����O��m��P��	�q�x�xad�45��P��N�)Q��7 a�P�I̟�����l�Iu��@�'o�7m��D���1� �YG��*T��o��p�I��p�	ԟ�'�b�&��T �[V`�����Qo��t��
�7��O��$�Ol�ăs���Y�V��6��O,��� 5d}i��ҍg���A��i�*�d�O���O���?�RHZ>��䢟�*�=pLz@�̑!a�xZ�q�z���O���O��B0�ʦ1��������?�JEN�-�YxphX�J!�b� ��M�����$�O�%"B2�����Ol�ʇ?��6ʏ;8dqr㞵��$a#N�(�M����?١튕^o�&�'6R�'��T�O��&\w��8��\�T�޸kb�lh꓄?�v�ieb�'�2ذ�O7�Rz,أ��ޕ���g�Ҍj˚�l�`;���4�?���?a�'�Z���?a��� X��G�M�б+� ��#�ѳ&�i |��'�S��f����t
��*v�`��U��E>��#eI�MS���?a�!>IT�i��'�2�'�Zwj8����f%�5�Ґb�@�Ц)$��0Ee��'�?���?y0�=>�iK�I��N�Yp�?"כ&�'�� �4���D�O����O���OM�DP!4�d0��a�6x蜱�e��*g�ɷB3���T�Iԟ���s��4dr���ݗ@A|��ԜqN����V��M����?���?)0W?Y�'����O�0t���о9��pi�B���O|�D�O��D�O���O�����R֦�����8���#ns�lB�!ɚ�M���?����?Q�����ON��@6���E�U�� q�b�Ʒc�0�J��Ԧ��I៤��ԟ8�'��YJ��;���y-4�Pf�X�X�>�w�FFߛ��'��'���'V�	+�'��'j��K5�D$X���@�X��qo���Iky�nN�2���d���Ӧ
/?���$J
VȜc��r�	ԟ���:;3����r�~��N_	BJ��g�	
�<�k��֦�'�]��|�a�O#2�O���Pz���G�h�Ç5"E �lޟ���VP��IA�)���yRG� s�D�Y���"�46m�6Z@�n�����������ē�?1PG�� �����%M����ƀ��
5\��|��	�Ob�6oљ?&�)�dƟ�A�ZAAî�æ�������I��ƕj�}��'���J�W�X-P��K�L�j��	)��֚|2C���yʟ>�$�O*��7r��`�6�K:CTNq��N�!��o�ӟ� d˗�ē�?�������C%Y�ɻ��/Y_`�����k}R��*?S�d�I��d$?m��#ŜcC��H��;S�ز�U�V�L,"N<���?�L>����?Av�@<��ۗ��Z�lc����2�tI�����D�O����O��� �jD:��-R7�DSp�}st#�	
H��"�Y������$��������U_ɟ���ůD:���k��|6p*�2���O��$�O��U;갰����+��#�iYE��1- �u���y�P6M�OH�O��d�O�Y�v��Of�'��x{�`�#�eA�DDZOZ���4�?����D;9pl�'>���?9{o���乺 �ſ2�P��d�^2���?���R�� ͓��S�c�}����g_6&��0$���M�*O�LI@�P�yQ���������'�yp�X�p��8�Q�]7+ ��4�?��e&�����S�'b��@rfd�4]Pҧn�Nf%oڱG�x��4�?����?��'s҉'�"R4^g�����Y�xOX��b���O7m�l���)��S�!�5>��9�K=R��X����Mc��?��yTԝ�xB�'���OTt�Ԁ�<������S�J��Q�i��'qv�
��>�	�O���O45���3ErЬ�� Ӗ<W(�p+���	�A� ��J<ͧ�(Oj8kaBH}R�m��d�^#�ȃ��i,r���U��Y�l���l��gy��!� 
����,{����N18 �H!�ˈ�d��'rR�	���hG�OJ��
c�O�*�(�Q�Z=̤�I�X��ݟ���ϟ@�'v"X;�v>1h��[�������Q�z(FM�>���hO��$,���d��b�����L�Z9��R( J&�' b�'�"�'�R�2���e?�p�$um���H�{t�{'�ۦ���Q�I柜�	3mĐ��`1�$ݖ#����f�4`�\�KM�}U���'��V� yւ�+��'�?!��+��`�¤�G�I�ڜG���؄�i]�O*Y��s�^-)�/ < 6�zSdZ��+1�i���'��@P��'\�8��֟�i��w�(���xtcK4��A��gӌ���O����i�B�1O���@� Ǐ�U�Q��Z
v~�KE�i;��*�`wӴ���OT�����&����9��hy��B�^�P,�hYs�ߦQy��)§�?A� ��q����	��Z�����R��V�'>��'t�9��0��O������2�[!PR8dbW�ֵd#$�)*�I-��b���I��P��/n,�"	&�8e���1��Zߴ�?0��c��'��'�ɧ5Ɔ%9d��˓�P-DB�X`	���$^��1O����O&��<�W��;t����'"(Wz$�Y���77����0�x��'�|��'"N��d�"4:�m ��Т�)�6�Q:�y��'d"�'��>]x[�O	r���TF��)�4� �ʭOv���O`�Ot���O�q+�\�@ ��|��Ѓ��̕q�����F�>!��?�����X���%>���J�h]��<A�
̣�/8�M#�����?)��Nn��>1�*T���$Mg�ȼQEiO��u�I����'_P*5���O����*j��Ĺaϧ���)@-J�� $���	��@x�/9�S�n��n��3`
r���ը��M�+O����_��������
��'������9)ą�3�ܭK��� �4�?����-Gx����Ȁ<A�\P',�8� !�&�7�M;��Y���'F��'#��D=���O��q`��X���[p�E�3�\�Qa��U�FM9�S�O+"j��/���׋�(�l����F�.7�Ox�d�O�,�6�e�I��0��C?�WA Crm��oߥM�H���`�n��<���?���0�����&�z�)�'d����i\��>7FO��$�O�Ok�1m��1 �Hvf���G� M�ər�b���I͟��xyb@��A�iܘuv��x���b&ص�`)��O��$#�$�O��d��/0����&ފ�p� � Q�J� hs%��O����O��v���C�=�`�:@�ƕ�nai� ʃnN�2PV���	۟t$���I۟��°>ICGH�&
�ڧ'��Z�≹#M�{}R�'���'��I8T>�D�O|
'� c�1jTc�@�jؙ6�� d��v�'��'�b�'�B�x�}��d���C�.nT�A�S��M����?�(O�)�a�r�ş$��dPA9$h�#�I�S�}-d"O<����?Ic��"<��O��X��Md(�bB�s�90޴�?���wv�u���?�.O��)�<�1څ2Ԃݟ	���#	8��n����'�&=ҏ��DJ�'����'�$#J*�  �\��MSTM�|���'/2�'f�t�/�4�<y���	g	��۶�.��d�������Y��|�<���C&�̊�Y@*@��ϔ+K�����i	r�'�"a�)?��'3��ܟt��h���lE$�N苰$�3u�pr��I��ħ�?9���?Y���pv��  ț�A�����A�k�6�' 
m(�M(�$�O��d9���,�B�̀.5��YiR\�,
��1�Iğ�I����'5��y���:H���hS��+5�&1��d+0��O��O*�O�$�Ot�XR�P7'b���F- H�]���BT/1Ot���Oz��<�E�0󉕚ey,�SA�%�Lh "��$Z��ݟ��	U�ݟ��I�(X��U���� �_ uT���s�i���'���'�rU�h2�bK)�ħ2��ڑ�N2��p��":.,zB�iZ��|��'["�D���'�8�����Y��AI��_��`�4�?�����W-�0t$>��	�?���
�<����& H���M�憹���?���uEx������c�<`O�k��)uy17�iV�I�Er�ȳ�4mS���4�����$���xz2�d�< �s<��'N2Ț	�O���6�G:�r��!#��T��i���A+g�����O��d����$�����1]yhS�H<-���P�_� Ĥ���4m�\pEx��I�O��qv��o�D��GC�Ae�Xd��즁��ȟD�	�N��M<����?��'�½pKŧ7��q3� F֝K�}����٘'���'����S�xi���ǻ���9&n�`d6�Ot�Pa��s��l�	E�i�I����<j\P�*�y
$9g�>��Zl̓�?����?Y(O�Ā�H�'V4�DhU�I+lTZ��p�քZ��t&�������%������L�`�G7��<1T��[B$f�#�$�O��D�O*ʓ^o( �>������
�VY����*YJ��`�W�������&������$i��>&�]+_ZU�� 5H�:ň�ǖ^}��'F��'��I2)����N|z�� 򰘓ҢX88����~�`pS�i�|��'��&��'��,w O��&�����4�?�����[�=Xƌ'>����?m�I���U�u��ZoR2������?1���$Fx�����c)*)�A ��%P�A��iw�	�S80-��4d��Ɵ�����DP]Ĩ�"�g��w�~d��LF���'eݗ�O���P��o�50�ܢ�.W�y`><`�i����v�'b_�X�S՟<��|yrG�;���u�<m�~�;�f�6���LS�Dx��d�'�����˟xa�&# }�	��eӀ��O��$M	����'�S����I.q�R�xJ�U"�$������2���O����O
)���Z��hW�CQ�zd�����	�.8�	ϟH�'�|R�J0@f�mcS�0d�@�d�Q(h-$����,?9���?����?��A�.��"���F�pt��4m�Ɂ�����Ĭ<������?��'�L(�rLP^����ґ:B��*ߴZ��|�'x��'�BP�,{gH���D��@�N�b%�2h�(��c������OV���O���9��~�ǃ
�d��y�G�ܫ�:X"�Av}"�'���'R�'7���s^>%��h���	�e�$Y���b���%;�^��4�?L>�����d�,#ɉ'FPq�Z�,d`Q�\�� �s�I�}��`p6(,��Z��A�	����VOh���a��^+p�th i�~��x8����(xAG"�8� +ېx2�נ,�V�[�ك�f`�1��{Pt��o�� ʀ	� kD�N�GĔ�!�nɫ⍝��.��@i�ox$���dð}&��N���\*A�W!��z$���1x����3��<�U��*II�QH�1�b<�#��C	�|:eK���ƳB��x�T��:�ĹȂ�%{�����h¸w� X0���*(r�'���'��֝2��)b.� |��p*ӷh��������?����b��Q�g�I�J6�Q�T�#`����R!Cީ�g�Q�~���[�U�(U�9�҂WzDd�O#b��Ӣ��[��=K�L���&��;��!�!�ŭ�?!�O8�C6��퉿 �ZUZG����p� xY�B�9-��e���K�dG��5�P.%���a6���S����'���"�2`�n<*w�@	QLLsWŚ�F:� ��'&��'EB+mݑ�	˟�ͧH���!ap���W���c����Pa<�aB�SO��P�	L/�����흀�&u��PK�\���9th�x!�
�T���+����<���t�M�Da��!�L5�d�J܄ȓ|�̓wB������wKG/e6R��<)����^$mZ���	�H�t��Nё ��Q @(�0��I䟌#3�ڟT��џ "U�\$S�)�#��������هH`@4p��Nu�A����� >G���ɓJy^L�񢊘����'��00*P�Ɖ���	g���Es��{D�B�[�8ua��]Jg��'�|i�J�O�o��M��lT�	e��Dmd�&�]܂E�.O2���Ot�O>QQ1*��-��i[6�̇�`�I��0�X��4j���j�HW*;e��T�z���I�iX�I�'�ۅ �ȟ��	[���:6"R�1�-Z�nQ�M;�-����dS��$�O69�w�O�b��g~2�$#��$���>7`� �I7��ɲx�"<����N�$ժV>؂H�Q*\i�D-6x��4��i�Xr���G��DiI��f�!�J�@`��a��Te0��&���F�ax�1ғ?=�P���ҡo��	���ǳ{=�U�óix�'�B���:ÒЂ��'�2�'T�w�.Y;2�ùa�,Z������P�I��3�,R�(�O��+s��1�1��'(���h�5M�����C`B �G(]�V���_�[�5�D��4[1��PG A��yΚ�a6�[1�O;�hP�#&ஓOf@�=O1��'W�-�1��! ��P�+�6�n��'�8|���G�Q����#־%|�M�O\�Fz��i5 r!�p�	.V�骂D�?8�B��7��}��D�O�$�Od%�;�?9����t�R� �$�@�E�.� W�׈Y�U0!

��0?q�C�X�hHR*��!�v�'���&�$��EE[��H��B�t,���ARO�� 5�ŀe(���O��D�OP��?���͙j�ٹ�FA�N]������y��R�3�$���\Pڤ���n�-՘'<Z币�'7�	8wD�`]w�B�'�,�:�!�yo<�s4����|2�'2M�E�r�'���]O���|�M�	F��jN()�B�K��T��p<!g��r�h��Řm
�
Ȩ�֩H5Đ��ɵ+D"�dg≺H,@Pi,e-�M��#��,%&C�	�L����C�+:ͪY�PH
a�C��:�M��ƀ=�aR��6Y��ˢ�_`̓~.<J��i~b�'u�S9
��I6m�h 怳�:E����as�L�	�xS�/^�Z�>9(5eƯ]���:�S�V>�۲�78�Њ_�Ourm�e�)}RD��2d����F:���V�K�@��[����7�H�̧2`��&#D�c�&��'�ހ�O$�Ї�')p�O�� ~���bC i:T	؃o�; �t|2q"O� �	�{�Y�"�߻j�,#0�'7x#=�2CܑA7�0fg�4�!c�̚�-2���'���'-ZA"�!���'L��y7nӛ!O>\�Z�9i0���n�>��=)�cξN�bݒ�&��n��T�!��KA��UT�JL�@ǡ^�dU�
��oqU֩@�7k����4^��E��M�#)�2]-���;FK��yH�B�(� �Y����"U�3��O
��U���P6��3N��1 �ا2��a��Cx��[w�Tp�L��Lv @=�'�"=�'��:|��Р_2�f�St�B ��X��猄z0q��?9���?��������O��b�1�
���\��IĔ#�x�Ӷi�j��`����1�	�犹@����a�#֦*9&) ���P��B��&S��
Ş�Y��������{�DJ	&���D$>cm���$9K�`���?IN>	����y"�_:J썋���1P�<B�k��y��Q�� �1K�<(�1�B�͘'��6-�O�˓l��᧶i#R�'�`� ���
6��x�c�ϙc��)T�'�R�/<�r�'��IH q`x��+��c�>�`��z��i�TF�8O�������z�0 `�'��!B ���x/�E����C��Y�3d@�@v��3�7Iu�l��	�,�ԘW@�#9����=`őݟ��K<	TO2K0~5"�揌^p|���ʖd�<1��ƺE	2h
7��SK"�ːd�^<�T�i{�"d�Iɣ����oP�\�|Rd�r[�6�O��D�|bWᆖ�?i��W�* �:�":I�l�W(\��?���j����&N�q��a�-g*��˧(T���,J�?nh�q��)e��q�ORl٠�s�*m�S����Z���c�q�w���@���6��a�@�^9���^��y���>12`K⟌�H>�"��R�W�d8k�����f��J�<��H��a�{�N<��	�2�hO�GO�'����%_�m�p�Aw��!�jphqkӪ���O���D�3!PQ�)�O����Oh�4�F��!��ġ�-=R_*�'DN�Kk�y��c��/�z����d�:}r�	�{Xd�R�?.Ȅ��gK�D'BDxぅ=|>}n�;z��h��z|�O�&a���H꼫�Q/M?�@Qa%ʾ8��\�"����<I������>�D�O>��	d�����
t1F�֥�6%��B�ɛ=Y�Q��!�M=�\�bꈦ���1d�����՟l�'�`A���êq�,���M���(�#��7��,9W�'�2�'R�c�y�I矌ΧA#��$K�70�D���5�&0Se�W�N��+�g�y��`�m�ĝ�s�!U�P��%ӉL�����@ #6Z�E�0?2��e����3M=E¾��9��<V=iF��R�	���<���$\S؟��B+�}�jE1��X�l*Đ:��+D���QjZ�#���#*��l���A�=�I�M;O>I�Ȅ;�����j��)ղ5��i������I�"�x���ҟ��' �V�H��� &1:�`"��8�MCSB@�t6�`��/�
����]s8��Q�BB�b��B��6N��Y��^�I��tg��,PL ;�)�:Y�GȅqE��X1�$E�"�"-x�h��'�fxq�F]�q}����N�'�+�y��'��yBgD�^���cxJX��A��x��e��1��͔'e��Ʌ�Jpj����O��/ �i���'��S�O����I"!�F��K��1�{���r�`�	ȟ�"am���<������ ��u�c�8�F�g��x��R��1��?s���E��� �,�A�(<�# ���T,��>�)���+���Д�'}��R�J*G��B�I��5�.�'Uw|���1Z/���DNa�'���AGEh�8�po�?l���S!�l�����OZ�$�]
`�t"�Ov���O��4��q���۱%��9�� �(�@T�2�Q��2uB���?Y���jG�|�oP�2����+J}��ؗ�_�O��E��Nװ�`���DM�h�H���SզU��{�1	�oԸT
��"�JH9��x�k�������H���ӟ�>˓�?9��*�ve�7셓e�|��
���x�؏n�!��H�KjP5��^3��ąn�����'��I�l��'�ӻz޺\�B&�H�l˰Jb0���������_w��'P��5B�Z}��44�N,�#N
-5�<�VO��c�K�:->;�̢4º�i���`�!�� :(�\��>�b���I9-�0���'����IJ8���r�L�4[`h�7NSm�!���"9� R�	[¬
3���c�1O<QmZI�GT�ڴ�?���I���Jӥ?���'Ikap<2��?���?������޾S{����!M�\ ��C�B�� ���6%B�_ӂ���iK�$
�A�	�.V:��Ey�'m�Z��oOp�]0��3V�� Pa��buT�2�؟i��Q)�,�O�yGyra���?q��x�
��xh�HǠ�:J/��0C��y
� ��Ц�Ճ;1�����*bT���O
eoZ�3�����`V��q�ޢ:SD %��e �M��?i(�n�eb�O���cv2,k�I_1$������O��$#A�<��/�|�'�z��t��4����K�F���!L� �;�S����tzk����Y%5@���O"��Q�'��O�T��B�jZ֠���B'uo�qh�"O������dz����aN����'�X#=Q'�ʠ)� �e�}���c��Q�p��&�'o��'����e��C_��'����y
�Fܽp���**�գ�#�(p�L|X��>�&���%#Rj8�|rAșO��1���H�y1�0�W�ʘOxH��W� �T��ċE�r<���L>�V�*AlY�c��<pى(-�?��Ov������'l�O��(��!18n��Ɉ�vt<�p"Oʄ�\� �QG��
�F�C�&O��I��HO�5�'��I�s����䊊�JQd����2|n-�s��uO�,�	��P������\w�'��	�ro&y1T�ׅ6"q����,k<0)1��S*�ݨ3�_�e���	�(�l,aEcH�N��Y�0��W܆�´)�	`X��-��;� ����(4IW���̡0�m���I[�	ӟ�شBM���RS�'3d�Ó���������3@����ȓ	w ��fg�$�ƌ��)FR�� �<q6S���'���Vll�^���OZC$%��� �#�OI'P=���&�Ob��W!2����O��S0��B���J��$G ��'嚙he��p3`�-I�F��v�-B_�x�'��K��Uc"��	�ԭ� U�p�r��g�	7F�5K��}���I�$��Dj�	���d��#���ug�o%4C�IJ����͟>cV]h�h��=�$C����M�D� T�h1ƦH�c ��#��d�� �3�i���'��!)L,u�ɂM��y��遢c��Y�wlͪb���h
яKǖE��~�!��L���I�|zSg�ilTJ���/�����X��K�os��a�藃&�i�@~F�b?�  �R�[��� B$�a@�)�L5}�H��?D�i�6m�OH�?�h��N9�~�����Z������3�I�P��	28��4�p銗-�H8�0�I;j��D�y�'$\��o��s?`��u@U4$Ou��`b����O��D�3Ipv����Oz���O����� p��$ڸ	
���ƒ%Tt�0�ʏ)~
�f�28��!���%�"b>1$��pK�6�|��애	�x� T�8��P@�=	���ӱ	�Hg�>Q%���"�8О$[e�uM�1��iL��vI�!�)�3��̄z��z�@*�M��$V�'Z!�$��k�D��U"۫[��Сʔ0���	�HO>��g� �,����"۠LN�H5�ǜ6���c���П�	ǟ����u��'��7�T`"q SN1�6@�����CC���(c�]�3'�\p$����jD��l�(U�rh���������y�8[&-*|Od�篐���a
�@��
���'��J��=�O��Ys�X�0�� ����"O��A'�	됔�fO��uR�g�A��x����i���'��rpʘ@���6�Ti�H�[��'�Ǟ�mr�'��)Pv��|⠋�O���8$� �"�`�n��p<�Qe�I�iO��e��w#�k��QuE6`��I(�����_�	i��H I� �F��_�7W�C�I-)�0�jUc׶[�4�;�b �*+�C����M0�U�y<zl�L��L��D
�e�i�+�rԊ�i�'%�S/�D)̓wT�9V@H� :U*УBG:��ITH����8�<������s�J1�EK6>��5b�F5<1�O2�Fx���-ՆV�Z��C�˻E�^�C����u�����Y�)�S�k7�h�`.�ɺ����*\�LC�ɧS�d���C@��!��� =�L��Ąs�'R�i#D�8mĂ��U�[�@$�M��~Ӕ�d�O\�$��{���f�O����Or�4����K�
3��	".`��m+�ɳX��Dײi�P���'C�`|x(�C�qO� c��'����������掸AB�%�$�<���AF��L>�c*�B�`���^��)R`�a�<A$�_y_��b���X��9Т��T~�+!�S�O�p���g�mx�`QL�}��M9`R˼����'�R�'rGe���I�T�'j�Hz�j�:���!��sf�}<A��a��(BI�x�ԉZAJ�������b��U`vo�zy�[9;\�T`Hğh�	��Y`x���,I?&�\�����B�Մ�S�? �9�ň�c���F�_�Y�ΡҲ��]�+mX��p�i�B�'�`H���&���#�	.m�h4���'z�@W13Y�'��iLh��|b��� �\��v�^�w��饤Z?�p<I���D�'�L����֓C.�aBΤb]L؇㉳YO�$[Y�ɚlv�����X�_Gd�� Ͱ6x�C�I C^L�1��\��D��^i��C����M3��X@'ɣhC��O�q�?�K�iG��'�哇��-���+�k�"��2�M���Q[���	蟨!�2�,�h��4}*���'e8�72����e��&�h�N��p���?G�m�`�O�,�2@N�}�L����3oKp�(M��j��O��l��MK���O��,�0��F�Q[v�(nT�p�y��'0�yR�ͰB��`K�R�h��f ��0<���ɇbϚ��R+Su�8�Q0�8D-�|!޴�?i���?'(t�^$a���?!���?��;>z�Ѣ%�
yR����5���h�y���.��<Qp%�#}^�� 7N v ��b2�oܓ#*�����xg�P��,*��SuH�+TG��O>i5H���>�O�	��<v����PmU��"Oֹ���ڙ78�"G�:u;&`H����Y���2�����E(t.�G�O< M�A�n�f�̅������	����]w�R�'��鐡?<
�HUK�{�(uJPk�9\��ЅO�T)�@9H��m0f��7b�2l!�8He<g��G���4E�q����']�����6{��(H�ǒ����a��Y�!�$�nI� +r��kD̪fG��zi1O�1�>IR��kM���'�bM* ��3�C`�=B�ĳ5��'�,A"f�'�2>�� Rr�'�'Z�8� G��Pq �[m�x�{ǓFL�T�?A��͡.Z���Q��l����KA8�t����O��'�0�v��Tܨ�խ��"�ƴ��l!D���˗�(ӂ��G�m����'4�$��4�8	@E�L7�� ����Sf |�<�Y Vg�v�'�2R>m� n�şHY�A��'�vDz�na��JA˖�@X��'��:��'�1O�3?�P���Pc!�;%e�Xx�v��£A.��?�@d�!k&�,z֤Zs�l[I:}�,I��?���|���M�*(��S�U4R��̋t�­�y2πy���68��<�#g���0<�3�	,��	��ҭ`u����z���ش�?y��?�t �zj��q���?����?ͻ{t���*� EV�Q�CvV�E0�ȘSe��:%��pc�����>[D�����2t�3d��%���A� Aނ�P��#y� �{! D�g�	)�2Q�`m��vZ��e�-F��URH>��e���>�O���
>}�Y�g�s�TbU"O`��w�]�����Sg�.?�F+����،��S4&Դ J#�3����� E��ࠥl̉V�J���˟T�	ʟB^w�2�'5�	_������N3I�da����2OR�@SG����7	�%�g�'���q��,i�X��:�F)j��4��E3h��%+v}R�j���0<Qe/<�
8YJ��*�G"C!x���)�M#`�i��Q����M�����"pR�O[	�Ji�ȓFfp�$�^�t^�h��<�"}�<av���'�$\���|���	ퟔs�l�(Sdl�r�D,��q# ���I�D��I��0�'u�� o�3�J�"��O)T�f��'���z�@�P��[c�>O�����Q�9��Ik���-A�TU:#g�q��ՓDȴs�$���	P(�D��ݘ�4�?1�p��,q���;�D��d�X8��d�O��"|*�`T	M��1H�&ǎu[��*���h<�a�i�2���<��aC��c�d�`�'��	9+�hI�������i�T�X$t��%�nY��W|��(f��!��'`������r���ڳ��=��T>ݗO���ca"ݿ-�|��dH�W7��H����Ő�����"N,��}�CN)�.��6l��'��4�``y���-kK2� ��I�+��+F�M�d�D�a�J�_m!��UY��dڇ��:b��phޭ/Oax��,ғ^����4L��<X�
A�T��kŹi���'��DűO����'*��'_�wvU��A2`���͍�&V܈��$E�)B�y���o���x�_`�$Avi�
Ǹ'L��ϓuJ�a;Q��'A( A�$9&�m��yb��$�?�}&���PBM(F�0<r�cړKjV�@�<T����&����1\��$�4��� ���3� "	rW� �v�f��wŏmtވڦ�LYAREkPI�O*�D�O���B�����?Q�Oz���q	L���Y b˒F�����ϖ�x�A�q�4Q��#95���3Yԅ;�'�<Q3�'W|~H(�(�����_��?a��'p�,V�P�zL�5���5}R �
�'\�L����(y�n��$	Zu憙Ȋy��%�ɺ��qٴ�?Y��o�t�J��HJ$��$�J`I���?AQ�%�?������?K>)���3T���EI;2�a�`�U8����(�I�?m����Πc�M���^Ҡ���C:���*���,A(�)��+\fm�a��LB!�����[�e./-��QN�u!��TĦI� @O! �Z���`W�/i�`1��
5��lZ����	N�D��0�b ��C�Hy�@N&W-���r�r�'j���'�1O�3?a��R��}���.R�X�0+A�D*j���?��M,_ ٪Ӭ�0�(XI��>}"'Y%�?���|���lU*Kڂ�ұ��>-H�jaK�y��܈Tt��b�gS�18�$C1/���0<Y��	�V� �@P,ϓ𢄙�D�/�vp`�4�?���?!��XٮPX���?	��?�;���҃*H�20�ph�n%*���y����<є�B���W	&W;�=�bB�v�>����	�D�v�{P�Q�8O A(pEN�Z��XL>0EN��>�O��;3��r�0�b�[T�AP"O&�p��@�e$De�!ξs�Ȥ����t1����.��9b�E��*	��(3�lZ듈\��D��ן����xj^wR�'��շy&9A��3�J(W�[�j9��9egt����k�:p�t���B+�D��i�
1�!�\� �i���/�Z�ybn]+j~����.����j)�!X6�ľRy��+��'5Z���>]N��J�z�j<��銣)j!�DނH���H�P+ZpԨ2�u1O�)�>΃�k˛f�'��nQ&x(�A�$.b��[�5��'�<����'f;���ID�'h�'W>�ŋ�$[|��a��vF,ya
Ǔ��a�?��B��"a�aZ�!
 ؆�a���P8��i���O4d'��q��\�QC���)3 ��{%`)D�ĠH�2;�|��͎�J� Bf�9�8[�4o��4��տ`|��/I�MJd��<�⮝�EK�V�'�rR>��!���(�	I�v�ܽRƯ?a��Bw�����ɯF�ra�	k�S��O
��b�3Ĉɢ�Kɪep���c�>��K�K���OY��2 I u���b�S�3��x1N��CUE�Op%��?�)��ɑsQl-���H(��<��6D�s���7�xs�.G#oA 8i� OAFz��۷�6���L�'��Z����y�H�!]'����+��	�2d��y2�C�&b80�T�	fQ+�E�:�y�K�!	X�Y�I-L,�	��y"fS�#bz-@����p��8����yLƕlkZd�D�2ml�+B�
�y#�O���a��]�n���]��y�'�k���G����(�yBL˪�u%�O��HS�](�y���K8p� �&x�Z�w�
��yBF�G�h����A����_��yb��6G�m�%�	&AuPx�A��4�yRIܠ����%l�@���[5�yb�� ɾ]�#`BT,� �`0�ybh�(|L�X�փ�h��A㑤�y"�z[���d��(f�����y�'�=2��Y1�� �MHf���yr�V5+tje�g�^<��n���yr#�/Wd`�Q>���ufp!�a!D�p��	�N��[%�� �zyPl D����Y5.>�ñG�)(R��""D���6MþD��I�6�$C#@�8Ƅ>D�`�BHZ�7~С*D�Y��$�O<D���r�%#���2*L ?��}p�o:D�� .��#(µ�.p:cE7s�D�jr"O,�B����+i�ѻ3Џs�����"O~�RUM�(P�I3N�+� ���"O�s툹l�A��q��"Ox�rM��&I>��%B7I����R"OYsf	�>/`x����9�h��e"Ohh&n� t���"�9|�f<�&"OR8��E8��ǀˎ���pA"OmH�M�y_�]���[l�$��6"O�}@�1An��T��d�&=�&"O�)j�k�!./R$���ӣ	��,�"O����UJ��)ZG<c.�#@"O�L� `����a	�F�>.�K6"O�{s`Ղ!�,D���)v�i�"O(�3BH/��e炏�;�"O(�k��ښ�z�&�Z D�4�a"Ovp�7-�4�T#�7T��"Ov��)�-Wk�&�V+CR�"Opl���]9�xY�
��Ƣ��fO��`G΋#��������\E�q�.6d�9PE�;<h(	Hۓ{XEQ��C2UP���.)t3�Ȇ�ɧ$*���7M:hf-�qۀ(���x�N2��91���4?���	�'�	�ŗ"��@KF�Jp��'��ҟ�pҥD��Q���'P��z����)ҜG%vAR	��0�쀛���:a|b̤��$�aރR 8���QDm� J,- J�[Z8��H���� �
@��9&?O��E��O�H��/w����I5"�~19҃w��%�$���45��T`��eY��)�[�o$)R�����&�Y�퍾"���ҊXN�d�#'��I��<%ǚ"$L ���LY�~�"��`�ܓ�~���yV c�''� ,��� �x�1��F�p��	�'�p�r�)� �h �b#V2	���x�'r,F�6}� .���@�l�HJ��k4��Pt�|)�F�^n.���-��C��A�۷��O��pwA-��F#�\a�'+Ӄ%���FU�:���6=22<Z��/�Td�=���?�����&0Rr#���	8��!��"��Π�Dx��	�Q��
BJS��%?7\�Z��`��=H����m�z�D�=���[����}��@(�G�E�TC·&�	]�|���@g��|�g����ɓc�=��T?�I�a����ҟ.�>�2� �Hʂ���G@
w��A"qKU�?\`አ$(.��rc@R7TT��]?qGyb)�%�
e9d�E/HH@������y"�H�����M;b!�U��el�����VO<$� *�>o}��6�,
>��1�M�:�ͱR���!3�̠���˻}#�U�)�,K5�5��
�C9��q#o �jK��[�@�{N��:�K�?w�!��,��5�g�����3�g@�t��Q_�@x�\$�� ,�$x�#<�b�~#����ډn���I	������T�E鐨Y>���\-"��a3T�M����B(y��`�	V�t@�L�za�gV>���Ɵ�r{&���Â$�����p�|�)�k
��-K�%I����Ώ�2����?�������4m�8;O����n	/\#R��c��[���
�|m�р�*D��m�O�Q��i7��3�p��hS�u|��U�|Ӧ]{DfT�?)�ʈ�j�)��O"q��`C�F�����M�2۾��tc�3,�湪���� ��1��=����g��*�Q�ȫN�3x�8���gW�#�*���l� =�����<a��u8����~�@ ��q��Ӂ`�u6B�w�T!�OI*�
Ǫ�$~s�:\5�g�ۙ�O�p8u�O
��H��y��s�n�a��̞cp���O�J�N��e-֨���;&׸���TZ^r�hDW?�
�/]�6����OG�GN�~<2�N��޹�4h[�$��i��ށASn���S��!#�G!J�����o\T��'"�9ӳ�ϝ<�zy{vNG�d���F��}�������#od�	ĮO-��S~�'( ��m�:��d�D����Y�
�����C�h�~Pȶ��E~B
�HQX���eW+@a`t� ]���M?�ȃ�%���IDi��O���ӈ��H��(*��$TH����t�x�I	�Pՠy��\�=^���x����/Gd�̱r�v����&��R,;u(�'"�R#ӭ�d����R��3p�HF����V��Q(ǉ� c^,��ꗍd��|�a	��L[H�6��8�n����5� و���~b��V3�в(�ƽ�婉�k>�ړ'κZ���{k8^iX��K�]��Q'Ǡ�b�B�C3-��}��/_�?�+O�y�'�;�����b����HM�S�r�1J��X�c�C�$�말(O�]#'�2N���j��� w �IE�̥p�(��·�,Jql����/3�X��
�*��ƼR 	**��E�d�b��\`E`�)ʀ�!��X�*q�L9Tg���j��'�~��<&���/�>M�<��i�lPJ�b��=uB�`I�Z8���T,"h��H2\�آ��8k܃��R�8$�����o^8Q����]�=S_��'xx*D��I¨��	ޚCjR�д"�8$/�r��>i�f��>i�GJ�Y~�KAJêHb���yB���n��4�A��9R&��C@���X9���_��h�a$m�*y��x�P?�Fy
� <��V�!.,��ͻ^n�;��<.e����Ђ~�н��FZ�T?7�~�E͏�	��ə�/�=X;�k�*��T�I�䃉�y{a|ZcQ�ģ�+��5�7�U4#��U`���2���1/��	s��'s��M�?š�X��,H;�Ő�D:���m� ��<�rΛ	t)�'�$�%��#NڈH�v�^�2V
\cwnP��?᠅8�	1��r�F�*����̀/$�ğAw�@j�l�=�
5*Ukݖ**�'��hP�ƚm���vI����g?Q�ǟ�{�&5�S�+o/p���`#]�>=q�'>Xxy�˗,D��ᙃ1�+��DN�K�M�a�~�l���		�ɵ���0�s��`)x��,Orٲ�'A�Ul$����\�;T���E��o��)Z�N�)(�ʴ��Gq*1#�-�	y�x3ҤPi��9p�S}�̋��~��,O0D���|Qۑ¨ai���X}����B�Tzc����y�ʂV�r�H�a��<���"۪r.(E.��p�V	i�OF�3hA�����i馉�2��� �R� ��h�([(�X�$бu?����y�,��5���P�p��*G��o�'�fq�u�Ըv>m�q�T�-�<  %X�\�+c��4Y�Zt�f��#@��P����Z�'��tkQ.v�t�t��6*� �)��Q"?5�⇬�P+A_��A���U���4.�0�i^�M�wQ�B��!��+� ]ߐ���Z�9W$+0"��Ot|A�C�"+����Hl��Й8��Đu��0�����$h����i�>Zf�8�ֽ>���OC���-_v�I� 5HL��v�P� ��#<�,�����.qIŢ��)X~<�,��¹i�t� �� ������{��!ZSN	4� `�>�Иv:X�'x.�����0 Ƶ����Xy*t��g��$�"Dȇlc���U����J�x��\n]��n��ZHXh觸O߸��@B��,���gN��m�,�Xw��
,T銦	�-?n�X٢��5W����퉇Kop$����%(���_����҇s��ݓB�R@?b'� ���i-���rk��4
��;\��E��L��Q^R�-���X�P�'L�mM����	�&z� �K��ߵȆkQ���T;��BL�z�(��[�,8���^�WD>6�R���U)��t7O
@�S������S�Ҹ �i0JqF!r���O�`RR�f������C�Pȷ��4��tm�E
u�"���x����D+�P E�ФQ%h�(��sB<�y�S�
E
t��h$��l���d\�ba ��'���@3�ۿ��4(���D
�|`5�-tC���u`M�&��H ٦�>����ܖ6��{�*U�tLۗE�>"�M)���C�ʁ�Aה=	P��'��t�'��� �/���`SD"Q/6!�X,�y��4A,�fʖD���<��0�K��N�6�=
�/ֺ4������tO�i׈/��kҍ����������k>xi�D%#��y ��4��r�w��T�O�����+(-*��A�1��F��.�~#<q���-�VQXPdߣR�b��-�\~B ���ub�
B�?��i�����O���ըK. ���D��f�]E�'���a�ŀG�:Xk��ؿM4�%a��>v.Zzp�������@kH2�0<�晥�$L�pbNE:����G�I?�#i��S�
)��Dŕ}�L� ���`�'A����B���A��F�J� �A����xOY6��"��5y��E�Ǎ2q�d���>�0<ɗ^
�n��;-���0�v9Qa�j��Ƹ	Ӳ	�-O3�pc�+ 5&.b���O��$�'���sDj���@�	�m¼#�pp��$O"NΚ�9��/�6�>7�_�R`M8FOI ��]q�+_'Eg�U*�Ƥ#t�����5w8�tPp�/�`8�HE��;:�U ��@�� ��������M%��T?�-�x�(u>-����Z9��AB�G�.(Ѓ%�2����	$_L4�ej�%[ M�$Ǆ�IO\�I&6X�X�Lx�
��o��O�L��O��5���Dǜ!q���%6�=96(H�	��Bp�	r�'�0�������@({��
�銲G���p�+~g�'*����|�I�הb��i`�L�����fS!Lp�Q�+ړn��"��1ҧ51>�SU%6����"� ֐Y[�<1�fk����@ !+H��]"_@���3��v�="��Ұb!BB�	�j&(��(�?��I�[�8�`t2�}R)^X��4*
� �Q���fb߻7ִ����7 ���3�+O�1Z�j�#_��1F�޼�M3�'h�n9��`M�X��0$b����#o�����
����0c��w�6Ii�� O���'opl�ֈ�A���IG)��7�fl�M>��O� �f,����,R�$˂d��I���!�WoY.`�pJ�״��0��C�m�'9���!MS
���F.!6��Y���\n���O�;`���P)����v�O�T�b]��H-�HE�`�쫔�Y�ꌋA+�}v�ӤW� �7&�d�����F��@{*dx��0ʓ�05p�(	�tbDL���Zm��iuC#G��J#N4ʓ0�Tm�V�[T~"�ϧ'��K:{i���Tn�}x&E@ !ܰ��$׼K'(�Cld�$��8�SB�G̓�(5��B�E�'2
�+%�S)f�b��587�!C���h/>	��/�|o���e	��Ey�A�m�H�oZ�U�䬹�E�u�� �ZY��p3g� ��'��Qq�o�y�nuS�O͓{Ȯ� 1S����삑K��q*pG�y�<���>A�C�{���1�I �NAIr��E�'�\$�AN�2��Āڽ:S��[T�T ]l�=bw����ܩ7��Uџ���)C3'L��r�Q�X���Þ~8dj�Y��P���vP��S�? �Ax�n�4j�����:Ñ%	�woa}�+{�}���1We����K��]�h.�	��}ARh���(���|�����I�잣=4�d����gZh���&]�2D���u/ۍu�9�F��tib�#v�a�6u�ǔ#5p��+��e�P� ��>ilG}K��E�ǆ.v��p�Nn��cu 8��#H����00̚ e�d	�'���:1���!V)Y#CБz�Q>��Q�):̵���	-LZ���"�5U�6����LI۞��`�y��d�C��>Fp�!�퓋��D��@�����'\m�s.�/g��i�p�#������j��J"%�
X���/Q����i_xX�J��lhF��-R�x��'�\�Ԅ�$H�
'��@��>"VeXC��2�ޜo�f�C�?D��#�
�:Z�l ��"Z��@��U�r(p��qŶ��� �܎�q��'��!��j%��1��=A����'ט�9b�M�U7�1�+��cl8��'Y�����5ZDд��.`!�\j
�'D��K�J�_K*����G'\�t�	�'/\��T�.,"T Q�R����'��ʧZ%PAl   C�8G�<��'� +uE�Z�u�TH�#0=�9�'3t�3m��D���8G�L6���	�'.$�Q��2Vs�b6��*dG�H	�'a�I�V��\�
�:V�b@��;	�'X0���Jݡl�\(�d�P�����'ؠBs�̨��Y�H�!���3�'A&�#cb:2�]���&�f,#�'AV����.l�┐���� �'��t���gx��24�N����h�'z����3J]F��I� e*D1�'B�t	��w=�h1����W'b<i�'��(��Ɇ,���j3���$�� ��'�BV�͞D��9�����u�
�'+t%槕�Xd�f�	M,�]c�',R�(ΰnHv�a���EHR��'��	(̤y��Z�e�N�R���'�B�G
I�~Α�)A�5�hD��'$P�v ܰm�0PRB��2I���
�'�~���@3.�`X���R�0R�!q�'| ��K�>1��YP#�#"����'��$�$��h�t�EE���
�'#��Ұ�U6VX�x�H���NI0
�']��Yd�/"�<�ĉ!\�ŀ�'�L�tk�i(�:`�ÿ	!���'�4U;��J�]��T�tΗ�yh�Z�'l�"��Q��B`�L;#{�U��'�:�rD$t~,�W��R�^U�
�'-R��5�\��@��CE�`�
�'��"�A:T�0iV#˲>�	�'�����	.��bcY&��b	�'=h�k��"-�I��\������'5ց�D�t<���c��ؚ��'H��ՇJK��+��H0/R	X
�'� )��=��	���+��ш	�'~R�`�I��+�Z�s nT�'�l���'% �S�ܩ8��)E��� 4C�'tM6ɐ8����5l�-Ƚr�'�Ԉ�MטN�B����x ��'�x���#9�4���D(r�R�'�R��S*� ~*���/�4��4A�'^�T�ÓR�|����.%��͂
�'��m���;r�rE )�ԩ)�'`V�}~Ќ�,	b<� K<D�$2&9jn	��'�(>N8�� (D�Ț��=��6L3���N&D���!Wc�2�k��V����?D��k@EMc>�}k�oM*K�jЙp�!D�� �YR����'p"�%��4,�P"O��	�.�(U�(	åM=���@"Ob�
� ��4�zX�S�U���qg"Ox0����'K�&��f�ΥS��̋�"O
}�%��-<����f/��x����"O����+Z�"��Ȃ���|=Ne��"O��VN�$0Ө!:��Y$O`���"O����[�;ЉB�&��I�<�b"O����+�HU#
:Bv�"O�@
h��Z�NQ9#�� ��	��"O�XiëT]©aF� 3c�a#"O$�K��TG����
�<Wa� Ц"O@�ҧ�\��9z�C b[(�"O�d��?M>8��g��2[N8�"O�� ǀ�^X��:�̒ ��|�t"Op�"H�4"T�2i^�G��г�'����
��P�ƣ�*D|���'�j���Ʈ|���E�^!�V4��'���JCR(y���5 ��x�TY�	�'P�(��Y.:+8 5J]��8���'I����Ă �0I�Tń
^�%!�'�[0�G?J�  ��s<���'��x�G#U���:Qeò]`NQ2�'���:@/_�K/� r���C�9H�'s�ݨF���y�̽ eF�?Lּ��'UBX"*��B�F����Y�zT�3�'`E�v�^�\"��F-{�����8�'�4Ĳq�@V�"Iy���,G�v��R������A�D1��Q�2®���hO?��j�Al�a�e�HxR��,D���&B�� Ȋ@��(r���K�,D��9V�*N�(Rĝk�ݘ��(D�̱F`T0����NgD��S�G(D���Ѱ|6�HF��\ʀȕ(+D�`�ӦM�%�TQ�`�d$ɖO<�O��'�"�)�酰���Fo���P���'qp�s�5P�d��H�>5M� ����<щ�����,4�*;�e����G�!�d
.B���%��"BHd��&�#���G{���'���wEY�xV!�bə�|=���'ў"~��N9G+���?߾�K��X�'6a�d����dbC�W&�j�dT;�yrgʌi6���FQ!�� 2ƠÎ�0?�*O2�DX�Z!F�k� A.=�`���"O��4����b��X�vr����L>]�ecČ<�<����+|�@��	,�O�u�윛�^���ئ�91dę��^�ѧ��=a�JH�$ض�Ҹ�ȓWݞl��j��Q<L�[�gаuod��23�)�7ֻat��ADT�|����hO�>�B���8��A���Y5:�"􊗉4D����"����SHY'?�c��%D�0�d�N!m ���AF�2�Ӕ`?�O�'}B��ظ�"�I_\����'?�,K���:X�M�5�߾	�(@�'�8<ST,ۖf�6���(S��%��'k �Š�87�⹩��	 t6�i�'�2yB�>#Xh袩��x��I��'���M
>.��@s�@�l�,<�'{�0��˝qa��A� ]��us	�'����O"Q`z�7Ǒ�X�t*	�'
�Ҵ��/DH
�I̦��	�'q��Q ��0L�[V�B�vIp�3	�' T�iC�{�0���}q����� ��+g�/#ۘ8q�.���H�"Oؑx2o�=4�d��mF=l�
0)#"O����c|��R��֎Q'�Y�"O$��@��e��hfb �>�9�"O~X�׻:�|y�$դs� �9�"O��AuJ?wV��E��2,���:b"O�a��J��Z�6��f�:�0��"Ox4���ڢE��k6h��z! UQ�"O6�вǛ#FF�CD�àV
��"O��F$�Eg�����z���"O(!�!>���X�䖾<)�4��$}���剸ZC8������R�aV�� GN��?)���@*V5�T��KJ(��ػ���d�!�dW�a��\���0��&%�;U\azңf�ΒO�t9�&�RD��3Ԥ�"Op�kƎVI�5hvČ�>2��w"O��UG_���рC�%�n�;�"O��h��U�u~n�Ђ��X�:��S"O���&I�9EtΩ�B�,	�U�#"O�<��@�q���h����P����I� FaV���5/� "a��B�#<Ob7M)�I8?�^�����Zg�(i6�U�b�.B�	)��j�e@��0�1�Ӡ2]
B�ɖ3ʝBE �	 �$
��h�C�I�In�{E./OX�a��Ŏn�@C��7aE��(�m�;��msq��p7@C�I��^����	�_2v����B�	�ROF��íQ�0:z��DƉ�Dl���̓�hO�i�*Ba���D�V�@� �P̞�-"!�D�!L͆���C�U�f�0�*�6b�!��
�A2>�i��y�b��R��K�!���3襉�R/� 8�R�
}�ў���I-:�dj��K.@nM1�+�0&�ZB�I<mx���c�[�5$�$CUR�ZFH�ƓQ�V᠅�F;[g-Q%B�!21(1DyB�'N�D���(���q�:p�6p�'$���F�&kljp��i�O���	��>�W�>�S��{L��P���(� t
AJN�ͅ�	#=���>!��6l9��� ��H��8�Ga���z���Q��2��/R��YG:�y��K�>����2$�b`A�kA0�y���P�0��a W�=N����';az�5'e�E����w���z�f�y2" I��"�햲X�^}XѴ�y��.�N��*�Jh0�Aѣұ�y�#�D����/@9?
�E�Ci
�y�'	�\VE[%�_�%�R�Cr#��yb�"<B�\��@�/$���Y�y�/>��A���2lSBв	���y2��e�i� �̳f�N�;��D��yH��;F��*�*��mVP9�S-�y2��=e��@��mH.Y/�U� �T9�yBE��W��E�'�>��x��(��y���v��cP������C
���=��a!��/1��+��<�N����Ƥ	l!�ٟ$���	�K��,���J3b!���n�Iw�A�<��=9r�ٝ x!�䔴Tw>]��h]�Q�Z��d�L�}m!�_�n�8PY�i[0�p��\�Dl!�)�,�Ń�)UN�� ��&&WqO����Q��E��5J�8�V����lE{���y1I^e� ͒��..T3T"O��1��ݚ��(��J�/(�xT"O�����M�#����L!]��Ġ�"O� BuP��M��DIC%�#4M)�"O��w*T��F ���4�ɳ�"O
��!��T�i#BH�%i��a�"O����� �-U����5��"O�t���P*h.f��G/�4F��p�"OP$q���(آ��PE���W��pF�T��0rqp���J��eC���y.��	��+��E�IrUM�~2'.�S�O����.3d�y�)�L�2��' �W��?3YzdL6B�XŚ�'60(�Am����Ųd����S�h�m��U����~�v(���Y���|i�M8�ŉ,&<�-�q�ă	���ȓ)V4%��I�T����u�A)n�ȓQ�l�a_�f4�����x��"O>DX%bC�I_z��6jX�}��G"O,�Ȧ)̫,1��1H;1 �*�"O����+<�����Ě2$9bA��"O��)�X?� Đ�DT�$F��P�"O�h�ֆ�7!_�`G��J�9�"O��� @���\�u��[�Fi�q"Ozԋ3cP�
�h�!֩z/pM�
�'��At)[%���Y��L:�F�I�'���{��A"^�b�s���Fh	9�'�0���W��1��
��
�'<\�*#�W�U��)�G�Q�0�
�'32��6�J (s6�Y��4�|h�') �4�	%B�u������(�
�'��бdV�C�8ؖ��P��(
�'=d �Gėb8Dh�ׅ�^�!�'��TZ�l�6r�Y���o����'vѣ'!bp���@�5�N���'��"�'��0AB��N������'!���� �M�W�ǌ��K�'��: G@�8F�sׂ@�
���
�'|�BҌ�UoR�`ԇ{��l�
�'n肖�6I>b$�@�ż�x$�
�'|�@�ϧG��H�"j|����'�l�82�	FkR\�B�_	��X�'��@���0 ���/�>)��'���ѥ�*{fxٴ-��U�P�)�'��6�ܮ�c&Q�U���B
�'��5y����"(�W
R;�΅��'D��3g�++�LC��Õdz,��'���0�j_�P��閅ՊY����'{.)㤄84>|��a���F���'�f�b$�	m����CW24���X�'� ��!!P0dRq�U�W� l�'�����B�d~ke�ԑ��H8	�'�D�ĮS���)��U2>a����'H�TF2^y4� b�<ڞp��'>Qj���@}��)\. [�0��'��X��gE�=+��C��(���'�Pm� �fyVa��,� �̜��'���e
Z��:�)N��dn�X@�'�A�Ճ�@WL���
�ND���'8���'�s��U�Q�x���s�',��z$�� Ԛe1�M۴Cֶh��'�[C�ҬnԖ�j3m�#>iD�k�'a�UP�'N�8Q�����	�p�*�'�dI�T��	�r�;S �R&���'�\8���Q4d�a�Q8�e3�'�H���*Q��� �D&~]��'C`�9�+�"i�Ec�I� n6d1��� �\��R3XF�"ӂ�N5X�"O�M�v����t	�^�I<(4"O�Ej�X{~DU��Ϥc���{P"OZ-����/F�aԗ9���4"O:�����Pj�*dOlw� "O�أ�[~�Őf��xo���q"OX�H�f�s�A�69�a(�"O����эN�`����R2|2�}0"O�������Y�\�Mȱ`�"O�б�I882M�'L�0B�\W"Ob	Å�$-�\9#�$�M=�ءD"O���`F�mNl�§�T�dP�'I*�X"�F�	qı�6EN�Wu�i�'�`(�烢_C<]Kfc�2)|��'o@��&�η?K����VC|E �'.��p�*�>;$��4��)�'l�p�Q�ԅl���[�(�)+�
	�'،�:�N��^I��#'r�]�
�'O2�X�ֶWC�c2&֋$n���	�'X(�r��7^�8I�C8'2N=��'�,��Oo�b�`FgEJ\.a��'��0C��}���CU�mJȼ�'$���I���8)�N[�i��3�'o�]�L�����7�SOR�\��' r�3�)�� �U҂X�s#�M�
�'����'F�P�d��+�0sv�̣�'�|��e�Z3U�d��f�;�]3�'b}��
�6f��9���N�}��ԉ�'� @J$��׺d�we�	h���
�'�z-���Z6p�PZ��e���'x��b��7fޑ*�N�[5R�'�h�{j��Q�L�!̯F,B$��'
:5	V�=h�a�CR�H��}�'�����$5�IH�Q�N}j4��'R�,K�JPH��(��K,N�N���'�\�� (W�P�(Q�SEF*�9�'j��SE�*7aTq��,ќ;�2)�
�'�!˷M�aC�Q�Gg	`��{
�'�j�!�м�D(��	�^!]�	�'����M��L�L�jT�Bm�-X	�'@����O�7�z�I�$W������'�x!g
�/ؘ�Ӯ"����'00��/ٲl�<ac%�<0y�A��'��M����a{p0���("Z���'e��� B�'~���럗��U��'.���未9��� � ��C�'�6xK������A՟ t���'�N"t�� ?rr-���?��a�'Wȭ��l^
b������8� ��'�2��� �&��8A�U\V���'nJ�2�^,\ZD�p�<��
�'�H�R�"�/{��(����{tН��'��Cp&��e����V^)s��O�<1�/�&��)Ri���w%�q�<a֏�^���� �h\�bIk�<A#��50<���DL�jQ�8��k�<�2��1��#�fY>q��x��@@d�<wȅ7FV�IvA��V�4�*G��H�<Ɂ3.BF��P�Q�\A8\�F�H�<�`�4\��q�2�St
6l�m�<Q�&�4Pe��/r1�$+ь�B�<�`!� g�F��C'+ ̪���h�<��kѽz�z�2S���b:���ǂ�N�<I�'�5C�O^�2a�Eq���`�<� 0Ջ��mF�0eE�=Ld��q"O�Y)1�v�&-��,(���K$"O�(wbޜ �ڔ8���v��Di�"OlXP��M����ˡ��-7��L@�"O:���F�T~t�e#I����R"OL�i��6va����	G)����"O���@/�2���Gj��6h�� P"O�d�`̀r�<)�D�N�7���A"OD$P��%`a��g���6�!�"O �@Үv��p�eA�g�$Q��"O���pL˩I],�q�%��rv\I�"O�mB�-1C�~��$��s rM1�"O�1q6���g�dQ�pd�A��IG"O@	KC����4		�M��.�i�"O�4�D"�.`-���D��&*i�0b�"O���DX�JV�-1���XJ4@9�"O���ذi �hcܛ!J
E+R"O�	CU.��k8�yp���-Jd<KQ"O�
�P�3��9���N�Uj)��"O�I�Tj��ҽ��+X22�Ese"O��9�G��8���9�(8K� �"O�@��"�!�0:4ԧc��a�"Op�2&뀣P�6t�dΛZ�� �e"O�-s�j7O��Ƀ���)�l p"O"��gE�;���蔈Z�B���0"O�Q2�BW4�v@9��_G�HJ�"O aH�g��9�h=JMfP'"OH�toױ\�����"2�4Cq"O.��E��$-�޹�$_�Z���"O�57jC8{�hQ3 Û1Y1�u�"O�tk�
�+�nt둧O�K����"O�!4'��!��p$\� !��ڦ"O���"&̯T�HeY��2��"O<�$!Pylr5��R�ih"O���&�
O�d;����;�x"OV���/mJE��N�0!<�H�"Op9#ш֝>.r׏]����S"O�����_�a�(�)��^�P�΍�#"O�5Z3iȃs�J�3�
��A� �(�"OX��o�%�<W�%^���"�ZT�<92�;A�1ȳN�<.M����L�<�w\5IaN�6��T��$-�m�<a�j �/T�d��%u�*$xU�Mp�<�`��n
= 2l�%6
�;&��b�<qpB9I0�HP#Л�N�t�<��D�����["nn@�i��Wu�<y����p\R�#"O�`%��t�<�'B$
���Ґ��Ve��ѥ"�s�<	��!�(���
Z�d!�$EV�<�#!S2!�yxtJ��$q�M�<� I�#�XѺ�@��S �%�&��n�<IS��4Zԛ�k?0��1P�ll�<��D԰f|�"Dj�< }�];t�i�<�S�0�X���9>|��)	^�<!���"Xʑ��lK3���\�<ٰ�δݨ�pbE2EP:Q� �FV�<�b��q��9��A2)�4d��IQ�<�P	�#C�|���hT+6�ڍp@�w�<	�Ƶf��:��[�خt�W�~�<����g6V���JX�z~�5�am�{�<y�-M��m(@�E�!�:�9q!�w�<����c������A�d�Sfz�<��K���K"͕� v���m\l�<)���X�xҐ�Z!G�T�f�	j�<� d[�	�:�إ�"��V"O6��U@I�#��P���;mP|`"O���)�V�qj��߮b��P�"On���J+��)!�D�xU��:1"O�-��Ϩ8<p,�'��87= �q�"O��9qA�bCF��e ��"O�%�%d�9h|�v� �l�n�1"O���s����V�S�BX����K�"O�m�2,�-2�|��b��n�� �"O���G<����*8d�ntP�"O�,�bϴ5�I�"/�`��%@""O�eY"���'
��ZrM;[�%k�"Oܭ���b[A�&"�v�,��"O��`A!�v��t�V��+lr�c�"O"�8GB�&PX�is`jQU�	"O���cZ<h����IN�98���"O�$�3A >���p(�T�����"O̛af��~�@3꒙`p! c"O����I�lr��q��^"`���*O�4��M�h�Y0��#�^�c	�'v���d�5|�4F�5i�ы�'N�9�E�K��t(C`��Ě�'y:-�IL0���c�L�B!��+�'Ң��#�������j�0K �+
�'��`رb�]��b�@�h$yX�'P�Y֤	�\�L�g&U�{N�B�'>B�8�7j���E	� O��I�'g�ݸ�o�G��l���)�ܨ��'��	��+
Tޖ`�-�$s�%��'���GCɕiX�!���oh�L	�'��͚��9T&,���c�p��'Øt+䉟�+��11��_��h
�'|�hڄ�M H�Ї/O�":|�X�'"�Q����z�z�b\(�2ͺ�'."��@DZ�j���Wn�S|*� �'���w��5F��Y6J?�@D��'c���g�Ж��XI`��Y�T��
�''��1�*��v�H4L`����'e�iT`�/:�yE��7Cv��'��LJ����4	�8c�K�'���GK � ��r�i��.���@
�'"�5�)�,l|�q�e��%��
�'�������=��@E]�-�X[�'�����V�C( �+p�71�����'�E�w���-�z�7(S�����'aؘ�g`Q�Z=0!�H�,�*A2�'�T�2�T�>ob|q'��!*)`�(�'�&�AÃ���>�	��ZZ��=��'j�9�`���F��@��U�FAk�'i\�:���"m�*�qd�����I�'2�Y9Ċ�2%�����X�d�6H��'-���&#	�?A̙;�&+%�Z��'9�6��,m�Xd��DK����(�'*n|�ɚ/.���cv �FeJ�'��-��ȬOu
��%N	8
�tB�'Up8b`�}�
�ⵢ�Q�dc�'��8�cK�>�]ٕŃ�P|l�:�'�� (�!\�X̎}هɞ�7@I��'��Q�$I)@)*�� *+��)�'�t��`�o=�T8aĝ3/�B`J�'l}c&���C;X�"���'z� à��Pr�xC�K?|�����'��c5�Y�Q^�|��dK���s
�'ݨr�_�_��#���1P$���� H�:c!�QpJ��ä��tE����"O�!Gj	WT��+��<̎rV"O܈8%���\j���aǽ^���"O���d���g�գ%�� ��Ȃ�"O�D2��Y�3�.���$�L�1�"O8�o�yqd ʓ��s�^ a�"Or��adE�3X6�S4�q�}	d"OP���'#�\��Շ�7g$]�"O��p�`E-P�z���5:�a�"OP3�@��pRA��+ ��7"O��ڂo͸F2�㖯P4��"O���DO[�Ĭ)0.)�p�k�"O6�t#E�6���D�7F��	�"O���W�B�V^�=qc?OI�(s"OМRt%�~���0���s	؁%"O��s�S�`ԩ��%X��U"O�Qc��mJ�x#��ګ렔��"O^��T �xn���#&^�Ψ�R�"O�\�0��
�*	rB�a����"O�ۥaK�*��k.~�Q��"O��r��l42 b�$\�ct��@w"O������*�.�ꤍ��$Y\[""OZœ��r���"R�-j�i��"OЄ����jH�!�Ų�v"OV9��g��Q|֤�	��D�
�"O���蚰/I&}�0�,5��u"O�H[ %� t�����GC8��q"OZI��.\F��wf��04��B'"OLi"�N�_�P�PC�-UB��r"OΕJ��-vv�!1i�7n5(a�"Ox0rBg�V��0���˶9 �,�"O��bh��iQ�\�eFPrH���"O��󵇅e����
�w���"O�4�����e3����k����e"O�s���%t� q��k%���;C"Oz��R�3�t�B��F�k�@y:�*O&ų���3Vg�}�G?H��@�'�t���C!_Q���F ������
�'=&�cu�_TAh�x��@�2
�'���S�(ޛx��)���_->4(D��'\��J�.��ؾ5I�Q)-�:���'?,����ҹdh$�O��<�!
�'�Bik�$ت>���L@�G����	�'�tȒ��:z�c�Տ9����	�'���92�^�TIB���2{
mz	�'r�0��H�1y3�5�����|��(�'s�죲�ɐQ;r� ��]�����']BL�u.��YyvL��S�ʴc�'�� �jT7$	�ևϾE�4$��'z�,x�V� �m85��$51��'ܢ�
��֋W"x5{4 �X�<��'��y�o�
Z���bD��/K���'�@E��� ,2`5P4�D;�.p��'�v��0=f��JG�3$�r�'czљ'��F�Eٷ�τ1@Hj�'H����N��5�6�C�)"8<*�'8�ex1b�P,θ��3U8X��'�JЁ�/�/��9A���0'6�
�'0�	Ţ��'$ x;��
�!���
�'�%4GC(ABȥI�O��R�U�	�'cz�Õһ,^��B Z(Ҹ��'���!$ö\��Y�I53��P�'�.�H��:5����ϓ>'����']�3eǱV�P1��	摒	��� p�*`eӚyd���$#į)��3"O"��K>a�l%�WL%b��H�"O�@��˓� gLij���"kɨ��G"O�cL�u@I�"�� �(=3$"O��� $!�J�7ɕ�4�V��'"Of�(�mͺ:Q:�;�H�<���26"O>�@G�lӎy�4���O�X��B&D��b0ƕZ�'��Q4/%D�p A�uTN �+�Y5�y�#D� b�J֊M��t*"> ALY"@?D��ɱ�!�0�ү�[��I�V�8D�|�D�P ��A�H�w��C2D� JR� s�*)�U
.��h�q�=D���"���0Y�ƞ�����'D��i�c�K48� *[�"�e�8D�H`��C�gQ����X6��!(7D�P:���D�d���� x��ᛤ(5D��˖�
�����r��*}u�ձ,(D�<A�ioPP�� ��'2|�;�L!D���"Â�&\2�8�=��f=D��Pī�(B�%��%#w�ج�0.;D���W�,֌�� ��?!���+:D��xR�B;���S hX��H8�`L4D�[���>W#��Sʖmn��"&D����FCf<f`S�ʓ��ܱ� �#D�8z�T�X>�T�$��x>�"fG$D�8�e'��w�˃k�6\3
���$D����
kS��q�,��wʭ�w�<D�@��%�:�ZY�BԁI�^yfh=D�l�Bв����Љ)%^ �Pl/D��kgk�tR�A��Έ���I��)D��vC�:��y�QCL�=��� �'D�L�eSj�f�R7KK0�Ɲ+� 2D�,��
@%�a�v��Y���yg�4D�$I#�O-O��ę@�=n�z���4D���∁�g�V��A�.p�z-	��3D�hSWk˰0g :`Ӵf�\�T�>D�����H�@�d�0FCPf]\ma�k0D���}4����"b@A	r�;D������]�� aM�3�&�zĭ5D�(�%�.؂��&o�@%�C�3D�$�R � t���E�K�H~��g�4D�(ö��N�����(� =X�`r"n1D����	yF�]���Be�HX�-0D���e�(c�	K�Ɂ�C�(ir��2D�$#�h^�MU��R���69��2R�/D�����Ξ;�9�T�ތ��$Ifh,D�0��A�ceJ��۽=g��B�-D���S �� mr���*���,D�D+����I+��ړZ���1I+D�l�%�^�V$��SIN�=2��B>D��V��4H�6W���o��k�&?D���b�]) �:� ga�v�p�@ 0D���F�,��E�W�ir�`#-D��S�Vxp�R��G]�\DZ /)D�����V�L��A��R>yuH��B'D�H*3e6�Zh[�F�����U�$D�l�sj�1�lH�M��Xܲy�'$D��0��C���钪J�]r�y�Va D�,�@�]9'az��-�����e?D����aN5`2���`Rn�)c�>D���P$͛ �4��@ܪ&�r��.D�d�S.Y8&`�ؒS��I�v�;��?D��a���3�\�a��m
l�ҫ?D�� @��&+B4z���/[#"��E"O���0e:̫b�Ӡ�`�"Oʄ�!�Zp�:��3NX�R�����"O��Irj��;� $1���@u�E"OXԱ�$_�'�X�$+V�>X�	"O�xi�I�w���{�g�kPL���"O����F��x�QT�H) V���W"O�K�l� :>:AQ��M>��PT"O�',¤���T�.^8�"O~�Q��$>�e �e\����"Ot@3 .�J���������L:�"O�(��$G� `*؊�.!?�� p"OJ���J�4�W�E�� �"O�iH#iHG6@�s�T-����"Of�����F��Y�B%�`xٶ"O>,�B���4����\�Μ��"O*2`D&�}��g����E��"OD�j���Ѣ�fZw�iҠ"O,p;ǂD�BU�aB��luB�sp"O��dЈV�줉R�@4^�tA�"O~�A  ͳ����LA�uD�|f"O�9 �G�sɬ��cq��kt�	��y��q�Vh0Tn��Q�A�c�;�y�kQ��r��1E��X�Xsl���y�k�#�&T�pD�;v��6�7=!��j�l�;�)A'j~���B��<)!��?mo�����Z>,KE���\�P%!�D�$Ⱦ�l��[������/!�N3fԘ��eh��*(]��"
�Y�!�D�2"��X�h���d!մ�!�d�%yeyi���4iJ�� S�ѫh!�d�-x�z��7%��s@v�3`��5A�!�/��(X� �Y:�)������!�dʋk� #!��q����L�H�!�$�$!��sGȒ��J�[�Δ�!�U&��0��ͤ��h �F�jg!���|��Y��٨��}�RǞ(8{!���8���L	W���pH��?q!�D؞-~��u!M)Y��|���4 !�ē4�jȓ�睬����$�ٛn�!�$ί�"�p�Y����Qe�%h�!�DD	�} T��4����-&�!��A�y�v� ���	���!�6X�!�!B���Sg�ii���\S!�N�g��i�`��nl��ZW.!��^.)�,�cJ^�/�ji�C�ɷ�!�1�Д� 膰_[HxKE�4q|!��"T�\A(jH8U�m2��Cc!������XMZ�z d�3s !�$��x���1C,�V4{A�ʦ6!��*\��8�$��(��UY�@�l!�$I�^>�U��!M4�"���e�!��V���Mu��(L��qcH�]!�û_36���CaWZq���+A!�d�?�:�c�X�.��$kA�ߜ?S!��
�h���b�'\��r�7
H!��W��L�P�f	�9@!ɡG�!�$�An}���Z}8��[��Y�A�!�\�=�Dʤa�x4h�jE��d�!�ξ�<E�
Z-S/��:䂟�x!�$�V'�:fb�>]T���>�!��_�sR� Xd̜~r���Z�F�!�$43%��0bD�38y�ي�/u(!�d���rUbիV�w��C�+�+8�!�� ��&߽^� $b�W�X���
1"O��p4IT>X�̙Ѐ�?��@�4"O��cE�J�#J�h���2�� *@"O�I����u|�� ���S�f��w"OaAb��,{b��l�� �>X�G"O�r�AZ�N��KU+����"O�Sa��\��V�.��3$"OrYb�甌����2K�0B��11!"O�A�J\�d�@%���6i6�!F"O�����<+�=z�c�?��8ѵ"O�Xt�7E;��sR�&`U�Y+q"O�I�c���J�x�
�U�u��"O���m�8o��0�1��w/���"Of�
D�@ ��Ys�'�1U q��"Oxa+�l7>>��� �O8I*"O�y9�j'Th�0�`�s�� �"O�A�R�B�D�L��ͤd�ʼv"O
X�Q��q��U�위6�B!rc"OL�ӡ�U;�F ���~��	��"O��Y4ㄧb0����h\
{Dp�"Od����ʢ'�f-R@�ܹi<\AF"O��1�%�C���/@0Hk'"O��H&.�E�gޥ;���"O�L��ާ��exP�3���"O�Q��.MTĩ#��
����"O��ˤ ^hH���T(�q>\�9�"O��pǬ
OZt*5�ܔ&�̼��"O��q��hU�$�&��.b��eJ�"O�,�#�cdk4&�7� ��c"O�(����Τ�w��%�I�"OL($���pƵi��;����"O�0f�Ѱ"�@̠�D�&k32�@"O�QI��I}��8��V.%"�i��"O���c��5�,Y $��"�Tbf"O�U�����M0�����M��D�"O漪��V$E>4��	�T�X�"O�<:�#ͥ'�
��(	�c��P�A"Olęb�ʳ}�i˃�����"O� (��ݹ����0Ŧ�Sq"O2	����0%9ǋK�j�|A�A"O�]{M.�u"��	��h�b�"Ov�8�m��=���� Î-'`���"O������gC�A��AYAjTE��"OywaIb'��iB�ݝ*\�Kp"OB0���0<5�Ģ�=A�y�"O��z禕��\(��s  ��f"O������z���C�׷6`:�"OtQ��˅fo>�Ђ�f� ��"O`h��푍R²��G# %AЮp"O¼�&�\�� z�I�^Մ1��"ODВ�:��Qe�wo�1��"OPx1���vްk b�<q��U"OH�!>D�ttS�@Ԡ?hrEB�"O(�X�C�aD ��N+a֙�6*Ope{0���7l�Æ��q�� @�'[���*գCd@y���@���
�'���'�߅Qw�����.���

�'��HPюL�g��z�a� �҄��'�TS&f(H�����N@&�(��'�:`C�O���c7�Դ&[�8b�'p�l�Ǚ5j�أ�"�@��'zΌ`�&K�W< !�������'pz	�'l��P����o#;����'�����% oʡ�BOLIUv@��� �]!c�Z @�:��Q�?e��(��"O�m��M��	��5�`X(��@"O��a�T���� jN�?h����"O�	��'زR��"GI �L8(�"Oʬ���!ȍ78��7"O
�;�aX�\�X�h��+Hd)��"O�5��E�A0"p1FռT�D� "Oѻ�+{t�hcO���>X�"OX<)PˑB�"H
��|��r�"Onݣ� C�E�Z�@!��?���s4"O �P 8V�q릇�&?�N���"O,ٺ�'x��ucLĭp��8��"OB�"P��bP���ƫ��m��zV"O�}��#�8P`��� ŌT�¥��"O*IR&�5[a��!ЏӨ���p"O��� %N[�f0��-��@���a"O�؃����# ���Ӎ���є"O��
�U�1����Q�Q*o�� �"ORܛ�DS�sS0)c�ς/M�q��"ON!���խ��Q��o�1�@9�"O�ICPe�/y�Ix䎖�r�U&"O��HGϏ�7@�u�r�͒R:�p�v"Ozq�w�>�"Y6�D�F'l��"O�eK���1e0q�G�lV`w"O������<<��=0`�J�tiHu"�"O�)+t/��fբ���
Sp��b"O̸3����I1E8��=�a"O@i2-�"$\S�KRmb�{&"O ��q$K;,��e�ƁWx�u��"OV%� ��z4���Aց
N�j�"O��#�\ ���#Q&p�b��"Ob�:g`�[]�(��� 2�ZP�"O����r$�
9o;ą �o�&!��F�<���OMƤ�����?	!�D��i�Q�ή<�~@%`G�!�DD�I��+q���j�@/ ��!�A m��a ���Q��։I�!��Q}���`c��?Y"HPh���=<"!�d��6�<Q�M�C�m���O3!�DL.o�P<	� I�Io
����Wb!�$�'jg9�@ȓdc���$�dC!�ͭ-��X��&;���`��]�!�?]b��1��M�}B2�Jfኝt!�ٸK�z��˴,�b{���2�!��G4���q���6;��(3���)#�!�D��/ �
��p� Y��!�$٘l���*e���[|v��'O�Y�!�d�C���k�+c�`z���!�N�d�����R`f�ȷ/R��!�D��y"x�c�ڀa�:9�g�]�8�!�$�42��L�R��6K�3��t�!�$A/5Pe���TVJ2tq���5%�!��@1Z���E��245��zqH\��!�� �L��@�>*=���V��l�!���a�<��'�:0��� %
K!�d�5�v�Iw�C���5�b!���x����wD]�v��X%�R!!��Ǎv`���2-]�D	�%��Eń
!�H6?`��9U��	3�n�
��V<!!��ݝ;�x���������b㝳�!�$�{\`���A�[Z�8Jp��5N�!�Ξk�6�R��ap������[�!��!!>xX�D�.t-�` L�J�!�d�@8L@�&��,_bz�*��U�k�!�� �}aG�D?4�`�d�@ {�<��"O�x�"J�U�"�����3z�VUK�"O�@2�m����Z�bT(>�VQ��"O܈+���(��3b�3��uG"O�aj�^&;L��o�h{f	HT"Or�
4���V�UಧB�'l���"Ovtї%ӑI�ལ�f�xA0� "O$��3/��1q QJ!�"O�58q�Z��,����"'��r"O����K�(�D�N43�))�"O
D��ט=��y��j��4�`�"O� p,���������^����P"O�)�a��6�rT`0��T�*p��"O���0�1I��-`𧈘}�^q�'"O�d)�ヸ3�XI����G��La"O��8����
���"tF�+����"OI��*[1
���Ǔ�21��n,D�x�u
E�=*R���hO�L�<�wO6D��BC�LE��s#�+{�YH6D�x�$�Г#b� ��7|\�ђ��4D�hC��J+�����&��g���c��(D�H�����w�̉*�Ȁ-w�h�1D�(�O�
�4�qa��(��c�0D��P�&�vD����"iV�E��,D��AB�E]���T�%�X�"�*+D��
W`� p���zgAވK��h	�i*D��3���n��!��DZ��t��&�(D��0���.`����)�	�M&D�$'F�w�@�+��8Y���[[�y��®ΜY��[<B��e��	�yb$T1����!F������Hݴ�y�lLt��q�i����y"e�c��)C�&��$~\+���y"�+3�r�BG .wnep�gK�y��/�X5���_�-�ƥ8�G�.�y�)U� i��Y������"�yR�0X��@	���O�F�zC�ٱ�y��`1 *�>?�rt	c�1�y�ˮ#b���F�=���8��D �yr��<"��䁕�Hβ�2��0�y�˻v�v��Y�1�`�R
��yb��"��Z�Ҵ'��0�HG�y��D;h2@��mڜ'��9�V.=�yr,R ?,4�סIcx��G_��y�o�*#R�LPŏE*!�ȸu���y���~x��2e�%E�2�H��y2��<[�h���*�V%�gl��y�F1k ���`J��q���zǦ��yҎ	f�NmY� �f=(�3cN�y"n�%i�Yӄc@0��c�)�yB�ڔB�PD��%݂Z�&�q�G	��y���v��$ۖ��N߶����X��yr!_��n!!D�E�=gH�R��yb��-ʶ���(��E���rb��y���	!����.Q"� �q��yr�,�p�v$C�|��Fn��y��+V��� �G�4Ϩ0����y�a�8 �6�R3z/�M�#O�ybk����X��O�[�<uRR�=�y�bJ�x��`R���X�A���T��y�%R�yr|� ��8O�1�����y�.�9c5B��˅xQP���
��yr"���JE�FE[�b�,�fhW��y� '�]P,��T��1�ʝ�y
� �Q�(��)��-���7X1���T"O�3��'�*��6)�H�� ��"O�t��
S7 �8���C�?�u�"O�X���B�����#�?��h2"O8x2�Wt����#��V��"O�-��?2��҃���L�"OV���n]�N.���mI�=ن
�"Of}J5e\w��]���I�/�&��A"O�G	Jo`�7I�'x8���')�,���U�����m��3���'_<䊰�@���%�#��4��)��'�$1�Cd	,wÂ@�bcտ~%v�r�'�����Mm�T���.pr���'�(�D\�-�f9��Ö7��a��'i e�Rh�Rj���W@	�1�L��
�'�|{���4�4Ђ�`��Vl	�	�'����	
�(y&�DiW�a2���	�'���$Ay���6e�Y�(�*	�'��,����]���@�6���j$D��u+)t���#nA�)7�PKG$D���$���M��h�,����"�!D���G@����2�.q�8�t�4D���W �4>�*p�ޜ*���Э/D�xSR�k�j4���[?k�ԡ�$�:D�x��*�)>4�2V��/<�`���%D�l�F!�?�&ع�mĄ4�����%D���$����iI��C�����k6D���1i���JiC#.T�(k��4� D�<rqC)k�6�"��R'�9Pw�8D�`iu��t>��TT!Nn��
� 8D������ΌPׂ��ٻ�'(D�c�'�6H,^�뢤�+D
���;D��)�	'�`m��
�}����f+5D���c`^)O����bK�v)̐J�5D�p��%��Xy2��J1�\Y0C4D���dOJ>�fi�3�9yC!1D�h%I��U��A�w��?Y�ń!D�l��H	<~e���or�۲�>D�,���R�#��#�Ћ,gډC&�<D�l�Q���	�6耒��N�- W�9D�pٵ�+6�� fg0jڬ�Ш8D�`[w�+������
V��A��5D�8��&|>A���.�p�3D���ф\�WeTX;2���t���1D�L��mC�Yi�h��C2B�h8IЁ5D�$jE���Y��\�&, �0�l!��h5D���	�W8��A���i۬��#�2D�P[��_�-Vy��勡hlnA�&.D�p��4n/���I�D`B��%�)D� ��*��X ~x*��
	IU�&D�t["�C<I�P�f��'�4i��6D�� ��Ϥ
["\�G�v����T5D�T�f��kB�#')Y���HӤ�8D��PaM�nʬ�)�bU�;Q)�!D�(xw�̍C��͋��
|R]���!D���ǎ�j�N�z֡И@�!�S�%D��г�Д$�9�	̢m���`�-D�T� ME)M-6��&�`3�9���+D��r�dE�UX�Dj�`&d}9w�,D��K�.Up`���f�E�F�� *D� r��� <�Z(��"ҍ?�*�4D�T��b��M#ljs �!u��a�('D��cg�T(4I*"�_$6��\8�7D�|`bOK�5V�p!�N� 
0 �(�`5D�� b���H<P���T�S�J�s"O����	be���lҾ'��E��"O�$�S+�"v$��[�j[�1��;B"O��;��I6ir� �	_�-L(2"O�E��j�J��[�bۋ��k�"O(�C֨<EX��/�g��e�"O�hf���� }�� ,˚���"OT|��N-ZZI�5�����u"O�@P�%�fI�aC������ٖ"O��
f��N��a�j '�DY"1"O�9��g׬2�4��I�v�<}R"OR� I#���0���#� �"O�TH o��Ku�d�5��+U�vܲ�"O@b��Q�*N�2�W��x�"O�bk��>�B�B�i�w*DMk�"O�$+�
"��ảC±%�5A�"O~�tLȌ0>����!e�����"O������!d��҄YE�8�`"O�ô��J}l���J_�x���B "O*�(#�{���!.�u���j�!��
&	��xᓅ��.$���J��!�DE2 q&9с���� �G�-�!�܅"蚈*s	���D����\�!��4,����Î˧2M8��&'I�n�!�dC>c��!�(�,rK
�94&̶�!�$G<oorԡ���7$��2�H�7�!�dI�/�X�������֛Yx!�Ą3G/r5�5� 5! 8�� r!�jlC�O�F�,=�c�Zj!�V�lN��n��,���%�E!�D��|�U��U�c���:�"H�!�d�*$�H{cc���e���A�k�!�d�0{���f�sFF�{c�A�E�!�D2+�P˗K�:0����}!��`;^���E���Ĉ5N
	e!���1�~�H'%��?�=���	L!�7a��u15 �>a�02�l�-#!�d�9:��.�'w'N]��HF!�d�S�p�pOM>"PQ���dX!�d"j"���6-�H��3 �"Q�!�p2�q�i�{
��׭���!�D��9S@+Շe���񅍡!���#$�$��@�3��L+%�Y,u!��XqM`�i\;d�1����`,!�	0[.�Q2�A�6>D}�Q��/!�Dֺ��|�rj�"�ZXR�i�T/!�$S)"m��)-��t��F-!�ׇ��9��cV�-�m3����>!�D�P\���A�8 p9�RD�6p5!��H�MS9�#�T>�X�PB��n!�ć�M��0;��R?uW���`ʃ*#!���F΢lK1��kS�1$!��Y0%U��j��1�v&F0!��I^~Q
 �rG
E���_,�!�5�����`X�1+����*�!�dNe����Iј}����"�)�!��L
Q�%W�Y s�z���bӊs�!�D�gh�+��J0 ��yP�!��!�Ȋl~l��R�jDa���L�!�䂵���',X����*K�4!�Ḓ�����*�� 1����!��0�t����!��I� i!��P���YpK�1$0�<���?h!�d�y��9[ U!7+6v!�� ���!�ϑs	�4�0�ܼd�P|e"O��*�]���U�ܪ���Z7"O�<��]�Cf�1�,�:.ٖY�'"O��k�7	��
s"-u�((��"O����)�SQ��2��b��pb""O�}�c��J��r��r܋�"OB�b������M�y���"O����\{�L���.�<`˄"Ot����%9�ry�QeKh2��"O��AE�O��8c��Ɋ9��Yڑ"OQ +\�S����-����"Oh���BX4����#��|���#�"O�y�Q2m< ,�ż+����"O����	:���n�0YJe��"O����_� xz�"�-I-i,��h�"OL`##ոMU�`"�>g���4"O����mT�'��9P�!��s
`�Y&"Ol�AT��t�(���a׷5���0�"OD}Y�L�8��4�ƀ��2kE"O�ʎ��2Y��J[��(�"O�)�ʂ0?���A $,P��Bv"O����%nh����,�n<p�"OؙS����$�t��^&U��US5"O8�����:�HhWO&j�����"O�˔xol�w�.^�jtZ�"O�����w�p�{&� C����"O�Y�񂎪)�D�`��c{�� "OT�C$�, .T�w,ʬj�=a�"O!u���@�z�±���"%`""O�hK�`U�)GT�"�G{ŪŪ�"Obm��#�$��Ԁҁ`Z(Â"O����H�-��]#� ШKE&M�g"Ol|S���a��($��� 2"O\�+�ܱ�ȠD�U�p�R"O��G�;>����^��Ͳ�"O̜��  �?J�er���~y
�"O0���	T� m� �$e�8�8�"O6�x׭�*4�Z��&Y�]kƔ��"O��1���w�����O�� �"OV,�UAԬO|�$(?/��2�"O����AM�9�Y#�F�8x�	��"O���V��W�&\���P�2�hf"O�lh�Nم=��-�B%��M8�"O��R(�1HJ	DG��W��l��"O�5� ��$U4dC'Gԭl��"O��c#E�]�)�e��0�C�"Ox��c����J^�7��� �"O�p�#�=��9:���&అ &"O��Q刉&�H�!A�̭�%���y�Ô�a9����e���Jώ�y"&N����C�ܚa|��bܔ�yrL��2����G��Wy�ū@�yRF�O��H􋞻Z����U�T��y�l�+{;�ђ`S�Y��!���*�yB!�%��1
���zFʈ��
Ȫ�y�!
# !i�`��e���R��/�yl3
���%,'�Hm�+�y�cʬ %�����s�bI�d��y�g 8�Լx� �7ehQ	�۔�y�>Y�0���3�� �@��yB擷�|�إn�S��p�M��yB"R%p�zp�wKb�A�BƁ��y�)��Z�T1�#��1�h�B��#�yb�Ǽ&BBU�� �' �������y
� ؅��h��SlA�ɟb��:�"O���ƆY.wg����F@��d�"O��B��N%���JdfO����9&"O�p����qĎ#�ը�h`�u"O(�rb�:x���CS<M-�]�E"O��E���f̐�c�0% Ͱ7"O��b�e����$��>L?���"O��"�1O�8���
A����"Op䢐aAgh,8§�1_��%"O�A��$�����%4o�
$s�"O\Y��@�st�B�0���"O��@�FB:#���fΐ�N�r�b�"O��2���1a� �9�TL��,��"O(ժUm�����`���{J�1��"O�(�&�����p{���Ͷ�2�"O�J�mx��!f� �|L��"O�(��}["}�ĝ�F�J�"O���RH�(h�5)�"��`����"Oc�g�?#�Jl׃ݨn���Q"O�hfH�*3�����	�Te�"OĀҐ�
$����D�c>��st"OT]�T	V,,č���X��"O�(d�$�a�
ٴ� "O*�Ƥ�}�dB�nNT"!"O49 ̄u�(��! �VTt��"O�XxBA�Y�(I�ː�5Tp�"Of���
�5P�u��ʏ�$H� "OD�Rw��,��T{j�j* �)e"O��2�+J#� P���U7"��:�"O�,�U FmJ=�n��r�("Ol�fN�/�~ �$�B�c,�Ȅ"O2�IJ;d��x#���l�i�"Ott�CO�V�Y��?y�m��"O� ;�K?4l�hh��+~¢���"O|\Ƀ)ΫDWB�{�W���Y�"O�ت���0K��,x��՟����p"O�����$Wѐ����@U"O��#1逤e�J$�̈M��hi@"O>x��:��pH�Z6
��5"O�UsO��E0u��n5%�Ykv"O��y��N�w����AG!+x�h{�"O.͈�&���	��ȝFK<8	�"O�U���ֱ�\�v�g9�P)v"O�	Q"JD�!�9�-��.�Ȩv�����I�i��JqN�0d>:�������C�ɺ;��t��dD:lc2�R G�:_sC�I�N���J�%Z	��&�"](F"=�2�$�'��i3��&#5�t���חq�����l*���fE6C3~}�Pѻb�Y�I.I-Q�"~��M>)�ݛ֭+wW4��I޷�x�H��_yr5"�DV��Yx��SA~C�I��$��bg�<(�pWB�L`A"O���1˖:/���;�2�hT"O�b�+H�w�p5) -B$a<��z�"O�i�e�ز�iA��Hs3X��S1On��DK(�M�g� {N�c�K�'萼�!��@�<Yф���Q�eGR7�@l0�G}�'<Bn]�Oٜ��`J�-��<Hi
~�v��O<��d�m]�ٛ!�s�р��%]�ɰS:Hq�?E�D�P^	d�شA5ʂ���Bç�y�G#<x0� ��U��1�CҸ'�a{aJ�n>V��-ČKuvY�JO&�y��I�5ɺe#V�P8�����ۣ�y�Ip��>M3�I|�j͢�l��	54D�� ؼZ@\�����#&��U�iE��Ҧ�������i^�d?D�eν)� L�"�U�y� �<*4T�T�l$ ��#�?��'�{"AI>�R]je�ڽ0�� �����HO�%0�{R�?q`vo#UL��p��i($P�S¦A�	m���ʡ��Yd1�uIM=��Mx��=O�=!�*ڿz�ȍ���&����CkPu�'ў�&�:L�A��%cW�=���=4�Do]�Ē�?��s���+�G�//b��PR䂯.��J�"O"��� U���EC��0Ff�y'�?|Oh0�$J+�ҭ����6y'Y�L������
�:��Ս^Ν)���nD�*��E��xb ǃqS���f�2�v|�4��=��{��
 ���Y-1:��h��S��y@J�Z7����%?�2��S�P��M���5��p�'��4���?7�D�ލ����Z�L11�H�P�!򄟎��u
�IP(
����,a�!�_��T����~���C���8!�Ds�`�o��u�X��W@4a�|I���if��PX�hI 	]��I�=[Zje8�:D�,�ԍ�.<����!"B:�^9��m4D��2�I>fĶ�A� �=(�Qp�&D��A���Hm��a �V�V(4C!���$O�ƑA7�чJ�ZIH�fȆZ�!�+/�99rC�~��LH�I�d!�Ʒ/��!y�JQ${v�P�D�PF!�$ö�,eQ����rL�wIW*R�!�$V�m�f��`�@-.�,0�(W�k�!�*d=�d�I��g���f��c�����	�=q\0D�L��	�f��<C�ɘ�h1�0NF�<8�A�c`<C�8*�zm��H(�ea�My�Xb��D{��Ԅ�H���rI̊{O�a��jY�B�	�� ���X�:�xLH&Nɧ �:���1�r�"V�Y9��%d�������I��Z	��������x'��E{���aƭk'tx�W��6��a�PAJ�yBD�B������4T���1KD���	�'�h��
�(@�32��>���O��x�=q'cx�"�;}���{�M�v$��6x6B�	�a$���ee� Xl8��iC���	-(n�Ic��ħu�xL�$T�#f�:�@TY6L�Dx"�)��ٹY+�|k$#@�A}���b!��?�"�O��I�<	��9O�L3�*��5��Y����kt] �"O����	�JBl+��F�b��"O�@��-!HΠ郅� ot���'V��i����-7"��d�.E�<�Bf�=G~!�yB�`Eb� .B�8S$@@�[�Ob���|B���"� s�k�w�)q�)LXH<ٱhN#Y�R��&'F��%I�iY�vd��'c�'n�>�I�\M�[�'�2h&HQ�E':"|�O���{r�ӷ�����j���H��:)p�G{��9O�iy$ҥ(l��oV�R:�:$3O��'�<p���Izy2�0G��2Q('����&���#�O~9:�ʌhAZ��ѫH�B�TA�0�Ŧ���`���@6-�'�m?j���_�b� �iV 2 ���_ce�M��|O��xB�F[���c��p��͇�k>U�sE�0�Z� ��.k#�L�'f�}�����@�g���`��X��yҮM�c�����E6yu�p�
Ŕ�yb��-Qtli�u#m� �3� ���5�S�O ��9��J0W�֡�^�\I�'U��1敲W�p�ӥ��\8����� �+��C3E���QJ�.ON] ��'���'A�D#t� -���I �̏�!�䑀		v��/�;.����V7~��ON��N�$2[��_[� ��M�{��d�0�p?� �)p��Eضk�DSEM�s�<q3F�p�.,�cc��s����MG�<)5m�W�r��M-N�0��h@��hO�O7�$�S�)?@��ćP�H΍��'D�l:4�,HT٠KѢT@�X2
�'t�9)O�
������C[D���'�$�#��N_�Y�"�P�@��'�ڕ�V��()���;��ĐH9���'�6b��ʬ|���1o�7@ƮaZ�'�X�B&��Vb ���`���RDOm����I�,m#l��.e~ ��ǔA$�B䉀q� �@D�:���K0�Q<B%�6m<�S��M�Q&�_���Ӣ�Չ%]k(L!���O� kr� 8��j���+I.ݫ "Or �d˶z�	0ԉ�*w���{��D��(O�O7 ��W�C
g�Pe���&x�Tr��~"��Bk�(3�hƬMr��A(����;�S�O�0���*�lh�2���-����}B�x2�S'#���f�]��[��F�lOB�	�`���cuAFJ�:�Nϻ:��O�"~�w��,m1���G�nRP�f�A(<��4qN�h��͑?���K�"{lE����s�J�k�3T�`��D]$��4; >D��s�A;~0��@̜�[��t#�L0D�<KCmѮ$'�̀C��9c	�k�'/��<�S�'[h��B���PEt�O�*���<Ls1FV�x�4��ˌ
y����ּ�B,�,u�Dk��@�E:��ȓz�[Uc]�q�BLv��2�ZD�ȓ(���Zb���}y�$��]f�@��(�"�sƛ�rF�#�k�:'�h��ȓ�ʡ��$H�u�@�u���ۆ�]:^�ӰӶ0N&в�G��-,��l(�!��ϗ��`��õ`9�\�ȓq�8i`�17��̰���5V�P���j��o�R�F!wǟ�DƆ\�ȓ�^�dJ�:�����<�D�ȓ	"ej���*iF(�+�^�Lc��ȓ>S�| b��l���O�K�Q�ȓ^zh4z��ĵkE��"ABC�*���ȓWm�����N�.5�qOڱS��%�ȓ|פ����:\N�uj�dիbv����kˬ��֮�l/�%�&���|0��X�
��Ө]i��Y:�����8G����
'AGn���BL�u����Fh@�V��qԈ��W��.��̆�gT&@"��~��4J�L��7��x������ɗ$�`�(�F��%���;��B�"}��h��$5J�مȓs��ɔ��
��� �"HE
���(Ȩl*Ӡ~�ȡ��ǎ).d<��
�'/Ұxd� l�����ǘ=1�Y
�'�x����90�$ܿh��t�	�'�^ �K3`�p ��YJP	�'#leB��� �ne{����M��
�'�J|�` �?�F�1Qa��V����	�'���Wj��*7R�0eV7G��a�	�'%6l�`���@i�7�GW���']�3v"E�0���Fc��?=� �'q�Ygh":�̕�u
�@m���� ��0k.��iPꕃw�a�R"OZ�pPm]�^��A���q/;D� �T�W��rjH�'�L�2�7D���V�)oZ���%��:��҄m#D�<*�Ɔ#\�1�"@�e�
`��  %ar���0/X!�H!LOMh MÍN��
V�����R�"O�mH���I��ZU��=O���"OThD/��e���2NBT�"O]jr��SNrY��֑A_<��f"Oz�%G����;NMbbS"O�y���ҲK<�h�?�,�X""Op�Bo�,E��Ve�	��,��"O�e�MV.iQ��@d�)!�	�"O:���� n6�<���B����B"O2�kƩÃ��c�� {l�*�"O �
u	l��AY��'B��M��"O`ɣG�_M]�8a_�ϢU��"O(��g��<�E@��(���"O���L�M��]�G�x���B"Oީ�ԇ�b�`A0�-E��q�"O�}�ňU�y">�j�ș4�P��"O��s�@�%��1�%B�)�b0"OFq�o�]��|���>E�,* "O�u9%a��*� [7D��JC"O`̩P%
+sb��(�� �Ci6��P"O	�o��ĜVM��i���'"Oh�5EN�x���G��'Md�!��"O��ABx�|�@�!n=vf"O�x�򍚧N���� ֊e7ډс"O����ݘ�"1!�e��@8Ё[0"O��wG����`��c@�SQ"O�����
3*��Xv�%3"O&}�Ξ/��P�EDV2�Rd�C"Of�aG:cK�, F�AA�v����O�K�%A��0>)�i�2 f���Ǫ�-&S�C�jP���r����	9ǹi��"#��i`��GMB=h'���
�'1�a!BcЍ=�`�鏋r��c�}�"G�k�R���ȍ@6Q>��a�LE2� ��Q�B�$h��	=D�`v�F�)�R��Bl�,\����baf�����,���	7NvQ>˓M�J�cq푉5jMq�e�������M�N�#⣐(C�B)J�ϊo=����"<��+��p���flXC���c-P�t�0!��ƀ�α!�:�0�iQ���C�b�����˸�+#m�d�6XX�E�2[ lhaF*��7A�D��-ְH �M\�7lv�@W�G���͓B�µS���vav\).�+ݤl`��:��O�a�$ٯI�p:��D&f�a�g`7J����^��!q3ʂ�ƞ�� ,Ŋ�$$�%hX�1�:��!���\�H`�c��2R��p��>1ৌ�hz^�-�1!c���ab�Yx���!�Pvژ���״���Vg �^�P䪤��.OpQk0*βkx`���/I�� ��$�<y��֢�.˧L��t2���2��)q�&Tk��DzOG�fd*= �� �ƴ�0�R)3�dDzfƓ�zhn�B�Gƣ0��p�S�RQ M��F��uyf�ɟ{����r�:�3�Č�?�^W��M����F�+�NQm��v�0y���R��hHŀV�/j��9w
Ӵz�1���Q�Á��t�B}����X�]�<�a�>C�H!0�~�vT�"I�s�D$i���o�HڧO�'/��,+��E��F��Q�O�|����r�F$a�K�`�\���F���Ӱ�J>S�Kwj�}8�h��I4�~l�HԶ�p	�I ,���x'� ��	�3��2����,Zw\�BRo2>
�D)IaӐIC��
�QC�TG@*f
#�#�,fE�E�]�l1$����I,d�����,�����banǴT�r�����+U���fip���|t���V�2�!P/6�XX0���f��;e�C���O"�SB���t�����	�A�F�c0�iK��aN�;*Ɋ��_*x pmh'D����3AS������ քsOƵ�a�^�${͛7$��� *R5�US3dԺqG~���P�ȬmZ�v�,@�ۈ/�`��S�-kHH�����r*��;+��
@&�7t�83 N�(�j��C�X� fZl������BٚF0+2��S 
��q�D)Z(��Ș���ө�0  #�pY��Ǜ�x}!�̛�I�~�3 ��h��i��TƬ��l?# �T1k���ha	��/H�r�sb��qآLZT%�<�.��)��t���M
�GQځ�S��9���YǏ�=p۪Xj$�݈?�>��щ�p��;�mJ$yBp�3Q�94�i�5O	������9
6���#�X��@���9{G~�{����=<1O|��>.L���Y���&�V��G=*I{���Y���%�\��L7#
O���Y���(�^��K1&C�R�_�Ix���d"�I5%���U�	W�Ap���g �I5%���U�	W�Bt���`'�O3"���S���ey���뵍�B#�EU-<��op���ﶍ�F(�J]'9��ju���챈�K*�HX-1��eƑ���g����XɠFrƑ���g����P��NzΙ���a����XɠFrǓ���u�jxgy�!�HIئ�*���~�n~g~�%�JLҬ�&���z�ewjr�)�MJڥ�-���s�co�:9�,�ئ�@3��qG�e�20�&�ߠ�F4��yN�o�:9�.�Ь�O:��sF�j�9���ҙ.�38��6��q�Θ����ՙ)�96��<��{	�ɐ����ؒ#�>3��<��{	�ɐ�����c9l`��t�r�-��`*�j0fl��~�}�-��h&�g:ni��{ �t�*��o!�l7a|���^���L�jjH�h��.ry���R���@�bmM�j��.ry���P�H�i`@�a��"~r�����$U���H��B�6��z+5g��*_���M��A�1��t!0`�� Q���M��H�;��t&5j��'���GfP����7z�;��YY���GfP����0r�7��TsR���Jj[����4{�;��YY���D�}�`�9�Ld4t99�:+RG�v�d�8�@k8y;<�0'VF�r�o�1�Fn=|?:�9,ZM�{�ir��|������)"c�3y��s�����-+i�>r��}������$#a�;p��M�mI��!.�]*�C~��M�hC�q�$(�[/�Dv��G�`D�t�&)�[/�Dv��AK���uΑȾ�?������B�	��ŝű�6������I���~Ƙø�9������K��T������|;�G���?n�\������t3�A���?n�\������|9�K���3b�V
������������K�6ж�}T����������H�1ٸ�xS�����������A�>ڹ�W�����R�e��G��)?N�Զ�2�S�e��G��-9I�ܾ�;�X�n��O��+>N�Զ�2�S�f�B&��$�\$&��uփ(�H!��!�\%(	��z؂(�I%��-�S/#��pы"�E.�d�3̞�@�E��@�p��*c�4ė�J�M��A�t��-d�3̞�	C�B��O���*a�0�q��Ԋ�&��A�]�NX�IT��Ռ�&��C��S�ES�DYt��ށ�+��K��P�ES�DYt���h�K�h�� �#�xS�� k�N�m��)�"�t]��
a�F�i�� �/�v]��d�B	�!4$-�?[4;���H"��,;)'�2T
>3���J"��,;)'�0V	:7���M%��*>-��>Ѱ<8��	�;B�ȍ����5۹4?��	�<D�ł����4ܽ13���1I�������8Ԏ�ub6�ڼ��;	����.���ub6�ڼ��;	����-���pg3�޿��:	����.���u`�f�A�� �6�`V�y ���j� A��$�:�lZ�z���n�@��+�0�fQ�q����b��+��~tw��Et�ȯz=X:��)��zps��Fv�ɯz=X:��+��~tw��Aq�Ϩ};]>��#�׭j�4g$���'�+�xc[�)x�h� 9j)���+�#�qkR�#r�`�	3`#���.�!�qkR�#r�`�	E�`7������]7tk8�E�a6������_7un=�zA�g>������V3so>�wM�f`�񑆬��1�"�%�D8��<h�������9�*�"�@;��<h�������9�(�!�C8��}=i����l#CLa�ډ�Ȁ�J�R��9�o @Ob�݁�Í�G�Z��8�i%DKf�ߏ�χ�O�U��=�h Au��pP�q��y �����<t��pP�q��y�����9q��qP�q��y �����<t���M(%~����h��5Շz6�I)%~����k��<ݍr9�I/"y����o��9؈v<�L*N�敛aM���I������$H�ᓞeN���I������!N�敛aM���J������&F��+j�����3�#��?$c�����0� ��|<&a�����0� ��|<&`�P�T\@g�Gl[
������'Q�QVJn�Ok]�����-[�T\Ae�C`W�����!V�Vu�[������i�Nߗ�p�X������i�Nߗ�p�X������烦c�Gא�t�Y��2��O�}A���(��`�T�;��@�M���"��k�U�0��M�~@���)��a�Q�3���\�D���9(-��=s*��W�\�D���9*.��:{#��\�T�A���8*(��:t-��U�\�����K��yZ�;�	T Z?���G��zX�;�[.V3 ���A��rP�3
�X,V3 ���u�9�Hy$֭PQ��c|~�r2�O|'ԭSW�a�y;�H{'ӪYY��f~}�x�錥=��4�uҞv�v���|�䁪1��1�pՖ�|���{�怪1��1�pՖ�|���{�公}x뷔�����,\����y ~췓 �����,[����z~곞 �����%Y����~�����ɷ�ƴp����/�n���˵�ǵp����/�n���β�;}����$�f���΢�W��@��XL����Aջ���P��M��PF����Bֶ̭�V��@��_O����Fв˥�����2)��^��gkΦ�F�����2)��]��oa«�K�����7*��[��kgª�L�����/��PW-f!�����l���)��]Y/g!�����a���+��Z_'m-����i���.�Տ;Lt�2l����Qs?➂6G~�:i����R|=㙅3Jp�2l����]~=���>Hp���A������!]�����F������,V��
���C������,V��	��At@n��n�.+��W� ��OyLe��e�)-��W�#��@vLd��e�+/��P�"��Cr@3 Y|�7k�-G�M�e�9	Qz�?c
�+D�M�e�9	Qz�;f�!N�E	�a�;V}��P�e���:	ٌD��5��Q�g���:	ٌF��2��P�i���?хN��?��U�dۖ�o�����Ztf!��z�dۖ�o�����R}l*��p�lݓ�j�����_vd#��{�dۖ�c;l���jC���Z*w�g�g<i�hN�r���]"~�n�h3f�nF�z���[*w�e�c:n5bߩ����h ��R����8iա���b+��^����5bߩ����h ��S���� 4b�|-J���j��l`��b��v$D���e��jg��g��|/I���b��jg��g��~,L��W�ߐ��0�k0bLZ�U��Y�Ҝ��5�l;mGP�X��^�О��1�k3dMZ�S��X䱟�8:L�?�6�����_/��?2F�2�<�����_/��?2D�:�7�����Z+��09Y���Sj`X�wż�c�u�d_���Qke]�tǽ�f�|�oR���\hc[�pͶ�n�~�lY����CӒ���%�D�'�ʯ�g,	�CӒ���%�G�!�å�k'�E֑���/�N�-�ɯ�g,	�CӒ���f;q���J�*��b�naC���j4���J�.��`�ehM���o?w���M�-��f�lbF���g�������c�<���������������a�;���������������c�<������������>{��`��h�����ER�5q��c��f�����@T�=x��j��d�����@T�=z�@��1�`��ĐZ퀰�J�D�9�h��ƒY聶�I�O��0�o����S⎿�E�N��  � O�C1^eyt�:q�D���D�xq��TD��H<��H�(*�,�{��)���ɲG�(�d��bLt� �� -��8Kt��Hj�`Fd��,�B��1B�:!�4&��fE\����")��<k䋒�=��:� /62>q�X/��K<��鋅�18r�L�����ʑ `���"�O�p������;jb�H�ț�@��8��L>�М��Ld�����
}��3h̺kf��Z�C�L�a�1�ޜ�c�$yw�(!��L���I��Ib(C(4�P� f1|���o�"�&������aR���Y>a��Q��A�o�s�E�+:��#&,���ƀ��bU����8�*�<����gZ4�('�:�`�*� >��C�B�H�Y"H�3�H8�cl�+�a�dњ$�4�H��ł:����9&���j  L�,���HN!v��	.�|��e�����#(E����ܢ4� diFo �j�LҒ�_]�9B�Og���f�!/L������!3� lI�OA"b_8�1��C��H3!�ܣe�����gy�bv�1�������:��������L��98�(ވ>Ѭ���*H8|G�i��-�6���3��8�������M��1(�H^q�P���8/R�c��S��"=��'�9w %e�#�;��իntz�{�:&H�E�Ű.J�0!���?{��a@�^T�B T8���c��?M�e�E0��'J�yb� � ߲�� a��^\;۴O/XPԣ��4h �nn�|˴�AC7�m�ABE	쭐&�7K%04jPE�Q.�8ەꑑ\�^m�D�� ^P�KE��1^��דwXJM�#�[��Hԭ�Om�AW�U�9e�Hz�ZC�
̀$F��u]FQ�S�˧V��@��A�On�mR���]���ؠ*�k*��X� �6t�ȅ��l�6p�c��<6Z2w	��l�>��*ʣQ�`���"w��Xؖ	,��b�N�41Zb���i�0��jJ#S�n�(��T�u+�}�E1���RA���L�4��/OL��
E��y����zrm���@&+�N$��f��N������*�A�����
�xIS�^���:A�զ�be �E2Ir�KT4P*>��R��T㞸[椈AXU��$5/���r&�zӞyBhC�o����F���]�tp3�l��%�,��F+ȹmQʩ�UL�7q��0!��v��읉�� ���.��@˖�Y�΅ Ь,��PI�OB=r�����$�̂�[�oD���JN�u�괱���|)���&DZ�Y��@I'�nC&��b
nE���jNr�����h��0IW�
	rx}Y2G�}�'�b%��&�E�A�r��^]��a o��Yf�@CMN�J�# E�L�}���1�qɔ�U;6	B`�0D[z�@s��J�D�3 �'	K�M��N
�4�ґ���D=k�%o
�l(`x6�'�Nt��F�X���j�悆g�֝��L���Ms"+ߗQ!�p�:sV�}x��#z�HJ� q��|�Uaׇ&B,RB�H�0�ux�͕[x](�ē�&r�h�}�!s"�� /	(u�x��耇IT�"g

�*�w!�H�NX�R�
�*�+�7�L��e�)%�]���R,n1�	����!6�v���$i�$��v#��i
�#>9��R��"���;��y��79y��!G��0�J�Kp���5�y��G�r&ҬI��;7��9S��6:��7�V�+�cQ�.��݀���`78%�L�Yw��Ģ�HG�w�t��B� 2���';�|`���pɐW/K�Lzs��ڨ q�JVx��@Aq�$6N�`��J��j�������M"`��D��xAP��㟓�hҦ�E FE�6mȪ~f���S�F�D� ���O�.���0���Q4$(���OL��Q���_�uң�یI;�ơ�������>�������t��!)>v �[�T���ء9�:��!�?�#���	�ӡ ,3����C�O�H�a虢?�R3�^�+:,��A��x�F�u&�$"��\#­9��=)R�M4&�>���h��md�d���7B���%����L�����H��O,k����5$�4�6��a�V�m�(s�E�2*n:M����#^��J��4ғu��-�"I�2�����EJ����A�L�6��b'H+t� �'���)\]��̓+q��z�+�O�#�����C<�0+�Ph�qAD��@������<�DE6JTha՛|D�a�� �C�m������~�]�5�B�HIS� Q�����y���[�:�{��Ûe�p��AG�S[<����<�փΌ8���&�8���9���λ3.�Р��P��|!$�Tx����I�Nv|x�!	H�V)��!r�]�*��H�%��f�ZhY��	Z̓f�^`I��)�;6���!o)��]���c�v�F}r���P-��əU�'}j�K%��M����5�(y+d��ȓ2F	���*L�n�V� &?8��'�2y�%@u�S�O�����#�*+�=��$�׸0�'�vHXC90 D�dC	�KTv�<�&Q�`�q��!�d�N�3�U~�<!��[7*�ȴ0�����3B�y�<�bK�W_Ƙ�Ul��=�A;w+�q�<ɤ�[���ec��b�����%�o�<��Ηk]:�*]	��s3�Zi�<10m��JtЂ@GY�v<��#�k�<����6���`���e��x*GTI�<ɗ.#�r�0�B�5*6P�%g�M�<�b�Υ`'4�l,@�i�eCv�<A�j�a��%S�F�,J��h�(p�<!Ơ�%����٫�T���ŋr�<駆�
��ɺ��W����RB�F�<I#C
-T��R�Ҟ
Ht��L�U�<��K� ���6�Bm��	�jP�<9î�l�
�`�&��v�4t�׉�x�<� �E��.F�^�eF؅IvP2"O>x��Թf%��+t�@�� EZ0"O�}[�*@�s�0(35�A,t�=� "O"Aw-(u�`�;O�+�~U��"O<q��ō|��kS��bq�1�a"O�xa�˹v�VP��M@,�pe��"OR��1]�wt�x��� �*!"OpA��H�LYhvѵ#bu;�*Ot�%F�9z�t�!".�y�r�
	�'�.P:u��(c>�Q� irpaS
�'�1�SI�@������0o��1	�'�x�����C�p��	6gw¹��'�����B8�ށ �L-Y)B��	�'~h��6��d�,�"��*R�ȍ+	�'����p�_�g�h:���A�v���':�e��B�*]4Q��;bj��	�'
����>?ޝ��(Q� �%"	�'�p�Pd��	T��[�MO�`@��'	vU{���zŮ�∐�
ple��'B<�RG���z��O��v��k�'��)۰嘻H7�c�Սmʨ�*�'��9�Q&s����G ]�j�B�'rH�Fd��-O��0Q2́Z�'B8N=`�����e��u����'�,�*�kضg!H��NX��$�'nZ=�!� �Cg��r�C.��
�'*� ˶(�\�����n��PX�	�'�y��f�*b)nX�7Bv%��'�>YP ⓪JWڄY�L |�~U�'���p��_8�]��(�%��e�
�'��(�uM)���'����
�'<�9�%K�g�������ƎA�	�'��b�#]�Cb,	��"#�����'�49�� \X��S��^�B��2�'a(�р� 	 ,�p���ٳ�c�'uh�y�ċ-�ЬhG��,^n����'���;sAPB�kAJYbZ���'A�����7R�X���,Xx�'<�����r�8Z�Γ�n�<h!�W0b�����;|O~3F�I�-2�1R�4�tp%#4��[r�G��|�ȓ�P��n߽1s�
4GײMӪ��>ٕ�5h�  j��:�(�|���-�ēv�Ԯ�^��R"OnaC�@Wxx�Z#'Y�[��k�lV7W	z��Ǭ4s�d�#�(�� 	���%&q�.��P@�`�~���� ���0/K�-G~�IW�ݘS�� ��.��,���֞p�ЕEJ/LO��ҥlC�
D�����jÄ�
D��+\�0�p�^-bd����)D���Li5��u�I1qT�q�W��,��([
�'��5A'K̰~�z��� M ]� ��'�� ˇ��k��`��.��	���1��^��&C�rv��	M�J��4*��n0�a)��'��9�d˶:
!��a_|������5A�@� #P~h�ɥ������2܂�Q}"���Hy������A�:9��OZ&��>���ڧ�
�ˤ�
)j��"pB��%���)q���"��"F��(�}�ٜ �	�i�Ky�%�<evL��O�⭯�Վ(G"ĳb�P�E8�(�|�c�GE�oM�a��3u%��ӂL�=wp\\���44<�#�L�nL����aB�ZS�O�|{�L�=,1��'�X�`��w�0PA���.+č3شx t�a��,C����cĺt��ҧ"A��c>��w�ӻ.A��;�.�=k+L�P-j,4�����W�>ͫ��'7�\�D�V�d�1A��fr�`;���H�xi�a!�#Q`y�@�O�h]x`@5�@�56��Ǔa�Mp%٨ ��W�O���>��0ON� "A�@��U,�:9 ��c�TDL�� Q��Z�Є��Y�<�PDğ�D�mZqzN�5������!�Ȫ��H�HT=cO|@��%�H��#=����qN|���#62Q��L�~�^�HWDF��k�7K�UPw��hoę�Q���M�q�Ԩt�bq�V&��
d���ѷ��'՞4�w�;[#�M��� ����4F���!�+�OSt�Հv�)O؛v�Dd�TQ�C@1��D�ق-ۮ8������Nb��;��[�+լ����N/,|d��Dӻi��y�t�Ɋ){��:�H�{�"���jOB���"�X�t�*}�w��:k��m�$d�/~��2�h�'}�0�� ��rWEQ�Vd	���/q~*� ����8>Bӎ����	aܘ�2�eD?_�iCd�)���`�c�F�3�5N��ڱ��oNdQ�k�V�]i��H+���@f�`�V�sP��y�tKԏ ��Bd�d�%��}0��w�H�>I`���m��	X�c�
J�������j�lA��v����V�.rHA��B)1���K�<
VxM9@"F@C8�B�l ��b���y�, ?���2,�L�&)2F�F0X���qI��)�������#`�~,ۥ`J����r̍�N�4j���2]
��ñ	L	NՎLD$�?  �u*��o�J����ɦEL��;p��
M>Q�D�<�0��+n�H扫|��A�6�۫H���x�2@��W�]�o$���IΏ��,Q��D�y��q����J���0-M�2Z����	:�.,K,��
�x��t8�� }B��K�x]��J pU�:P�N#
-F��w$S�b��a��^H$a@�)yA0F	�P��(�u��"X�ʇ$#g��Q�Ɉ�_M*A@��D��P����$�d�SEGH����4N9f�X��'u�0��
�:��Ɇ�D�ԁ��' �R��eb��݀��r��*JBbY�w�ʣ������/w�*�Ҵ$�}����j#��*G���OHv�';��˺h&5���׻5(.�S��O2ࢄӦ�ѱn�v�[�>C��H�nK�n/�F��81%4�;1�N�1笘�!^�pp�2�-Z )��`�!S�,앚��F�Ҷ%�2��f�ďP�E���H� x����O8,�򏊉2u�	�ė�y��	e�1.�h#Y0AKv�H ��RQ.˂/�0q�C$��	w�	�%�)�&�sř�|��cƆ-Z�X2���FAǎW����$�&f�D�$��r2���'�� s�(+��Ȕk7�TsW#	�xV0]k��2&�p�6�4u2����œ4${�<3�h?�d���2c�����"^��G*��Cnl�r,`m�<���'�(������iل���{ �!5�Aqf L2Ry((zU�������ڢh;��AEǂ�V\u�P�� H��9��C�P~8 "�!�6	��,O@��`�4)��y�U�7�H�kcG�hД#��`@�Z��2`|�1F�5$��!1�T/1�^��F�`��XS�?�d�Ԍ�s� ��ŸR"z1p�N4KŨa[�'� `iZ�:�$�MD�!	��Qa.�?i�-[�o��4��e<e`Ę��>3Ш�Fl��[�{v��N���3sڑj���!%��ah����M�2ڸ%�PO��Z^huR��C�^s.0��(�	��	�v��@Dơ �*����l*<�FCR�_f��2����"��U�"h4*A�ef�,t���ɰ��_b<0���[i��
������Zi$�VKמt��Udq.��x� J�z��w!��~���L�O r�]�b"��ǀ�\x�:6��IP�o�XH���K�"eA�mڣ	(���kH�Yoj]lI�1�� �9?����,��g�ۘD�ZݪƧ�r�����B�|ð�iD��-kyV am�=%��g��D�R�."&�����W���kB#�#.�R���T�!2,���C�� 9,��h�&�V�K�#Ҟy?�TO����$��<�|�\�� o
�/#����i��r=��o����$�bb
�,�
�顎VӦ)iҀcT\`�W�99��b2럑"���A��-=�l\�q#+~�ñ�?�$Q#*|�ˉ{J|�!R�l��!�������R��-8m�v���Y�P��aL��$}rų�j���M���8r>.(M�Lpt��IZ���)�)��<�5)Z�����r�ڨ ��P�$I<i@JuX�N��F!F�2�f�8I������
���('gb��d>mGDi`�N��C+RO�<�0���8�sG��#6�9k��'��љS!�i�A�eH<(Y��>y<�{F�ћDfLKVd#��b�B96=��[5 �-���IH����poԂD���cv�DT�E���{F��y����26����Ν8��1D
Z�J�n$2S��(���s��F��I��-#11�Ҡ;��4��H�`$:�m��t��`$��Kf5B�N�(M��'Jb9b��ݩO�n�X7�=��蒈��Y��(2�T�r���P���JT��V�ԅx9@�3���w�|)���*i�@I��R�Е�7�{�V�"@"�,��	q����x��w*o?i�-����/'�ܒ�J�f����l��6 P�ɐ�D�Y
6���H\#�`T��?�p�\%a����03
@�᠆����3R`4JW&d��ꂄ��(�t�	ED�`(�	�-L.���0;�D<\w��!�+J�¨t�U����fF'G�t����C�xl��4BI cd`|zDo��:���yR/׈�4�ȇ�׭M+�f&Ƨ�2��aM�q�����#@��["����	y��4�A�1=�}��C�+�&����n�y  �Oa�z�9�f5*�p�	�NU9��3}�H�� ���P�=��ԋ�fE>�8����")�q��')����/cx ]��ٴ~����0}g���!K�I֛&��<L}MI�O̲7j)��ɛ�[Ĳ�ӬO�t�U n�.a�1T� \03h
G�J-��J�@��	S��C�2��T)D���*m9�.�S�4H 3�B�Z ;0�R�G�-Rb��PC�0R��D1�6�@tN��&�^iY��
�&�B[��1�J���L՗v�dl"��Lh��'��
�Ta)��G$�0�	�ć�xD����U�r�dt �қIf���T�
�����@X[���!���}%P Q���\
���u�ʙ��'��Ăť�k���C1B�.���R��f�"�
Fۛ5[� ��/��u��Q�i/Re��13��	�@��Αf�&�eF�4\�ؠ/X	w��<9��3f��2עP�0%��F����!1�I*��=v栄0�,���M$�G3J����w�?�{E�+(��0@A��3�����Z;UT��	 L�[3�Ȯ?��KU�),��h�a��0��¡�:VQ�ѥ��t��Y �F aHfl���Vn�
�L��#�Vl	�,��k�cK����BɈ�l��b�bd�!G�<4N�X��c�= nhE	!AQrR�SäI�(9�SP&0�(u煽6K�P�������ykhtKW��W1�;��47�YX�i�4r�V,��Z�P���[#�hp[�ME2S:��!y�`t�`d��o�E��M!7r�÷聽|D0��cӖX)��Q�#V8x��Ӈ�>��d-s�
�/��e�p`�B˅�q��IYdF��Pp�hc�싇}/X%��Dd��u7O�p��bգp��}9��I�V|�p#u�
�x'L5
n�m�j�ʲ��=2�De3%`� "�,�'e����jA0H8$�U\�5���*o� $`d@Q�7��I��T��ԔN)Hd:�Č�}�E��k̥.�Z}��bD$7Gބ����'K��D�ү�O+J�]2�k���P�t!����JZ�		���5�b�+F�r��EXd��V��<&?	�h 0��4U�i��]a�*D!>z��dHOT�R��Y�2�ZbF�F�X����,1��QA��D#6j���Of��FS�i��p/�G/�	 �]�o*-��/�
q�2}R�����]�Y$�pӧ�}�:9r1�΁I�8�`SI�6~�E�dƌBf�H��;� �� �dB~�Pt�ǈ��ܪ�O�����C,�����^�](�2�.XbH`��o��"4����Q�d�����D�J���q b��!��f��Z`Vh���* ��0-���>��D��D«6���1�D��6�r�ť'?1S	3id�ʅ�
�,�D@u�V0̌ ���� �a���G?9�H]��$$B]��q �$,�b���O�	J�@2dś�I�HǾ:�DA���O%@^��9�w���S#��y���2��؛��a8�� .[�K֥8��?]*�ONک0�I�=Y"��cF���8�0%� �1<�-vf���!γS�ksC�b��=Zf� :�{�A�76�w>�6`�{�ޘ���f~��ӨU�m&��g({3D�p�GQ=�L9� S���@���0��)C� Rϸ9�d�D�wM�i���v� �Ӌ�3F�DD:W䛔{X�m G�B�7(��(�f�N~r}j�8OD�Z��ɈzR<��۔ǀ!��D�A���ȗ���}X�A!��ws\�
4�H	xW�GEZ�͒<��D/E�D|tL�T���F��zm����xR�H?�� ��M�.�>��P�w�~�۱f�$����Ι3��!IW�V>f4q!���`��q�h�r�j���F�!���H��1��5q׫׼P@����B�1i��	��v�5$�/k-�5,��*�_�^� 흹`ǬaBٍ��(�U	�)%�~�!�Y�\�bD��+�d���JF�=�E���(��<!iO)'�p�ɡ�XC�֥���ƅq}����&e�qAݪH/hH0��
�SI"�O�Ι�t�Gs~��3�A��%b�8A�� �$,5��*nHZ��'��<3
 ZXZyu
��R�����E5�r�A� yhz(iIĈEBv�i$#(r,$�'&F�H�p4�G0�Z�A�}fh1�	E
CMj�ydc@�����Y� 2��`�S�.U����1/Q �!�-z��#����L��@báH��4�7�X��L��T!&<�th�{��!K ��?H�������J��0�꘳����W�.. �x��DS4<LGz�!چm�% G�	x���"�+�]�&�%J(2�N]El�3�L�y��p�$bR#��-Q�&A�:�ڨ���%���DoqO���	�T���B�~Y�U���ed��@�b��{R�yJ Ȁ?��䱠,((\��Y$��/9����E��_L������>P�$��V���a�X�����I�>I\%+����L�\���cr�#�T0!��҄�	�|�z��@��<I�LH�"�(�#b�ޣ"��)��WC:�3b�B�/���_!`�z<�CÔ�8��	}K��c��0?;
`0�eF�J�"%�=��!ӓ���5[p,��)[��C��381|���F�`�<݈H����?�
���[p�LppS� #��O/n0�� �qsN1G1�Ȃ�c�*�02�џRJ@yGJ� ���P�tW��Pĕ�M�1`#Kh1J������RΕ4P9�=i���1T�}r���P����,Q�y"�@�9KDT�����zP�
V*�&b���D����)�GEX�a�hTr�ҲD��h5�
�&<0,q��&i5.���	Pؼ�R�cCR�'?�e�C�1C�����J�~)
r�`�� Q�/I
�>���B �z% �ːc����P꒙z%$z�@����1vHE@�ՅS'`��т؀
�� �	�#
��ڲIӱE�`Mh�¾`��j �.q	���3��I��ɫ� M-"k`0׀�+?S65ؤ��>n��:��V�q	����� J�������,'gx=P��XSlma�`�7$Z�p���]�O��Y�I�'�`"�	I(�e��hڵYPdyQ��hӦ4�b�D9
�Y�+jq��B�&�lid��A�3�
��j/�d��CN<Y�DN97�LD�vM$�p)���������A隄'��yЭD:3��� �ϝ��I���B�ÃI
	����1��(����<=��谌D����G#h^�Sr��'qX�pA�A8b�| .hZ�G|��D<L�<� !��!v9�&�(H�ڤQ�@η��	��֠i������
�HC�O��	nRQ&Z)J�ּ͓��1z�W<{HN��䞑��ڀ�<C�#=�P�^< ��8��I�RtaP�O���k
�6�P�I ,z���:QR^ٻuA�2�F�Q ,��$]����=[�a#㩄ʲ���h�MiE�Vl��|��L�e~1�c�Aki�M@���æA:��-s� �m�5
͖��i�)c�K��'�hSM0'���	Qʝ0���9D�>����u�eE��	#��k�
��]�P!@� �?Ez���E����ˁ�:�أ�DIg�Q�I+/�h���Ҥ�K��$�ߟ�J��Ϲ��!�نy�8�&�&EtT�q���m��IEc�Bm�{�W<d�pFE9`_
R��:$��l��O/[:�����fX���F|v��B��2* )o����I�wɮ����6א� � �CN���6��X�'��`���n��aP � &}�6n�`$Bp
ҘzVG$%gH�jB�#��)	���)��'K &����<q�h�k1�-����H�1�Ռ�ş��VC\@�}���]���O��b�NJ%���O�����X/b@*0�
�Nn����"O� �� [���`�7��]T���Jr?�&fӽ�.��R�G����*�b����y'�V��B�Ƃ����o�"�0?�"��:dڡ��R5F�5��&�7��T�ԅxW.Yk�yB�T�yU,]G|���7r�浠�L�C��M��cR���O�u3���l��0�����!5(y�5�Gq�9[v����y�엚�&����G�	�@��'��d�**]���{��ixΖ�����l{�p��j��M4!�P>f<[�f���4��Q�u9!��@��fmypM�)ze ���D!�d�.)��d��4iU����Y��!�䑏L��I�5c

C����kF�N2!���!F0���w�Y 1h��㪔R8!��j\3�dX�$�U�A��==�!�$�C������Bΐ��Dۓ.�!�dU#[p�{�LÇ0����"�W�!��Z�rEq��n=H�Ո�!�	;$>DJ7b�B����$�!��2x%D��"ǘ � �����=�!�U�z#�š�ξh�ʼcP����!�� 0p���1[�Aj�N	��ՠ�"O 41��j���K7�� �,��"O�u��@�%Ú�bS+�T�>I�a"Oz{D쏟1�Zt���H*t��b�"O^� $N�1D��y��8o
�S1"O�0�I��)I\8{�MuZ Y�b"OIk&��&���aCF�B����w"O���F��;��'���:�"O6d@�nϮ3.T���!��&p���"O@��Ӎ����b�Pq^T��"O2YP@�;��3��zhq�'"O���3eN2��d��h�5YR��"O�e��
:oz��g��[X,T�����S"��F#HuE�u�'1z9�pC�+N|6� l �fk�'y�� �gX5���H���01[޴����X������'�
i�+�~�b�] S�	�kB��A*A0(��:��l�D$)�>O �ᓥ��hF��B50X�Cg��K�\���yB#�5�y�d*�`���;�MB8\���#A�<�� ����P��0|z�oݲ;(΅�&ӛ�����1]&�'��h�I�㘧�OV�����#8��2Ď9dGVr�Oš�!w1O�>Պ��v�0��'��,V��A�t��8
��s�1O�?��3�8A	0H��3qza6������y"�$����W៖���@]�#z�=IB��ȞlN��r��ӭhCp��3Ɋi�<p�B��>}O�p�jŜ/|1O��(d ��ýP1$��V>d(Q �Ɵ�cB!<�N�����C_l�4�?N�p�������F@���Z�K�,@�rY�2�
��x��'V�O�����OP����!��8���%q1��h���2�S�[8�IJ�A<'���e.M�@�'Odᓋ���	�E���x��ZK~�������D��\��b>UR��Iզ=�ӭ��`��+�[<X8Mʅ�vӸQ�/O����I�<E�$MX�:~D0�g��U�<�$)�?҆�̓yg��Y��M��������ԟ�ɋ?�����\z �SCI�J�ꍺ�M���'�la�,�-��#]�a<�j�Ȃ.j�0M�ךx�х]�fc�b?eyT��QG,��#͐+߄����O��e��,/0ВOQ?�0�M�1'K�1�m��(�-���N��{��<A� �<E�Ν�;�]�rhۡ"�(�� �ލ����%*��&�"~��"
(��Xĭ��\d1QM��B�I.q�|����J�U�(�"�n��B�	.aЎ}���/	H�R4�T�~�<C�	=Y����C D*�s�jѺt2pB�5��ѧ��-�@k 	�<fPB�	��U�n�0Y�!����yIdɺ�'������L�}�0P$
�$�|u��'���Î�+d�~��#��<`�	�'�X-c�'�>,4=h�����A
	�' |�sF�^��.K�^?9�B!�ȓa��Y3�(a����`���͇�z����1��;HVd��N{:�-�ȓb��0
\/A3�t��i������^2���i�D�2�$nZҼt��d��U8��B0Ql�HEbS�)90��ȓ0�������m{����˺,t���C��9q%'�/_^R�)���X�ȓ*hH��Գ!"܅�3��L�Ĕ��K|�A��M����я�uAby��Z ;����/'Fa�#̀Vؤl�ȓ;��1G

>�����~}ʰ�ȓ;�إ#��pF����ݤ@f����8�i䖥d�@��C�	h���Ej�e�J�!f�%�vL�u��9��9_@Xr�m��,����#F�H�֑�ȓ*��$G�`��!�*/"�JE��it��q&� L�}c� ʧDi�P��S�? �ͱ6AJ���DY=/�T�ٶ"O$�2��*T2 ���!nIT9:V"O,�R�`�=z�b�� "@�l��q�"O��kֈ�A���C$��Q�"O��hC��ix>8�����ʲH��"Oȥh oߓ*v<=�� �2�{�"OL���j�>TC~�@�L�-�*LA"ON"� B,���prO��7�X"O��Ar���y���$��<'f�
�"Oܘ부�	�ă��U����'"Oq�Td�ls����A���@�ӥ"O6�H�-СHjJ�� ћL���C"O�t��W�H�9%FM�{y0�[F"O@8
��M��f��E��E�!"O�HY�˙A�9��,�_Z��1"O��ЅGI"=�����J��V�$��v"Op �!��E<�u�
�q�A�"OՊuIA<|�[pɎ�9�R�#"O��ۗ`H���!��*��u�Bx@R"Op�h��V�>X�8����O�`�1�"O�r�V�I��!�5\"t&AQ�"O�- �C֤e�����Mm.<�w"O!���=��R�M eB�\kf"O��a�AB��t�ʎm(���7"O�MSFi+Ę�2�͇^���"O>��C
[ ����Ι�y��)�"ONͩ5B��)�2�6��b�j���"Ot��L�M�rh!�̒?m���$"O4\���H�ZD�H����T��t�"O`%�ԒLEf�s �Ŭ��"OtYZ�^�
z&��G��$;㼜��"O��E�X�`��a�H$	Z�1�"OB�K7@�o�p�fdL�y@|z�"O�����)��E�B�W5�t2�"OL���,��V�p)��	54M+�"O��@mJ����8�j�:g>�R�"OM�=P��ت�	ȣ �h��5"O`��s��+��A����+�ʹ*F"Ohic��@>ʤ'��*y�1��"O0L�Gʐ<a�>4�bm�[T�0�R"O��ш��,Rl���'0���g"O(ih��rEppZ��		��	� "O�Q�^X��h�ueͻ���:W"O�š�=�hqI`O��J����"ON�J�OP01{���'��hO�$2"Ov�2d�m+�����0`����"OP��H���X�.�U��}�"Oz�21������5 � ����s"Ox��vIÑ+�C�Lߦ{���"O���ai�< T,�T+	�~O�"O(d TeR�F�v��`��)��4;�"O�� ��N�4�T	�B�����F"O�5�5�'2����a�"	o`���"O�`"��`�*X��լf��ջ!"Ol�L�eSֹ���-�.��C"Od0E�ߵi��+�RG��,+G"O��{��͏Z>R��2�R�X�<�3"Oly�!�_*L�Hq{v#�{J��KA"O�,�WlI?N����S��P�LЇ"O0��sK�*(D$��Z*���5"O�9Ӑ��18>��d���|��q�"OBA�c�S29L��� W�
|�"O�ʇ`5�$|��2��X��"O� HA�ؐ=Z�0FACi���@"O� *={��V	�����BT{d�p�#"O��Ң��6�+U��M�V�P�"O�����-Q�(=JF��{D$���"O.�r`ж�h�H��>0:�`"O�-����m�#H�$F#��{�"O\$p3�ّO��+A�P��p�u"O��k6�V�K̴�a�%H� _0�"O8�+�f�$~¡ɱ�ZL\"��U"O�QB�&ےe���qcY�c[�)q%"O�A���B!_T�|�� �11z	�R"O�m:w��S���k�R%m�渳5"O�����ӥF�2����2rvt4ba"OvЛ��.Z~����X�v�Z@"O�lp�گ7$Ȥ����(�tx2"OQq䇬k?�(�ȗ9P@�<��"OR�h@��/��+�@�&�IF"O�Q��g��5��eK g�.uhB'"O�c
G%h�����q`<���"O��" �=D8�5CSVƑz#"O��P�o�c�>M�'�!3#�l��"O�5�Ҫ�%!�"���'^) w"O�a��"V�q6��� ��a[��0r"OJiA2��
L�J!GK%n��a�2"O�Y�c�
�y���	d���>�:�&"O mQÉ#r�P��ge �u"�jP"O�=c�fFn���͂._]L�:�"O�8)��V�-��2UMM<	[H�1�"O��� �?o9x�vL�kL��z7"O���c`@@~��G��;+4,z�"O���4l�!�dij0�;!���"O�` �#OI&5h�B	�8�M�*O���$��$�Y �Tt��db�'�����+O�t��������[�'K���fN�����a�����'e�-�5�8x\��Ң
�5�x���'����	W`,���˨`4lh��'(�� ��-`���@[6�^��'��T�#��4Z`@�1|�V�'��)A�LqT7�����bS"O lhpʁ6z���͓�b�4L�2"O����(�q��ȑ�G��X0�"O���'�� �0��k��*@�X��"O0�CO�/�H�8S�A)~�q4"O&�:�c�NJ5���V���"O0�eN��\�uPV*�I �I�&"O�Y�k̀I��rH��$�,8��"O��R�J�>��d�q��ٓB"O*�a�D�I���R�б}b !�"O
]��-ňWÚlb!(t<)p4"O�Q(�f�R�Q��G�l]L�q�"O�l�D�Y'�Ґ*G�PWJN�RW"O�Y�ТU$HN��6N��3�DH�"O������LIz�[֍��r�� �S"O HKS��6RJHꦇ2r�&<х"O\� ��ۏ�.Ɋa��p���@s"Ob-�쑪>�ڹсő97EJP�3"O����/�A�e5;�Q��"Or}��^"/t�XŢM'44�r�"O��Y�R	_�^,y�N$ܡt"O��#�&�7e�*!�+҈J�下1"O�L�o^�_"[�I�b� �"O�(v�pa�H5.�� � "O��F�L�Sՠ��sF"t۪�h!"OP�
��R)9��3�H}��"O� �����<��;� �
��!�G"O��U��!-��
M���"%"O��V+�)({�� ���o���"O�@C��E�C��w���c""O��d�J��y�1	`Q4�bF"O栫E�O1ݤ�ӷ鉎s�L��@"O��F�O6&�|�Q�[����1�"O��bAhG�'r�HWjĝb�jix�"O�Q�6O��44�#�� �`@q"Oz���cͪ	�<��g�+:��$q�"O��d%�7x(B��W�F5(9z��2"Oڴ�Ŏ�+�a�2E�)I"t�"O Ǎ��!��k���-2�I�W"O��1G�Z�y� �V�K0h�,��"Ov����:2s��� F�P�t��"Oz���ŖSi2A�4�2���"O��r"�4*��m���'�N�� "O�x{�V�c�5·��B�6��"O��b�XTq$�[�D�(L����"O���ˋ�=��9`�K�c��r�"O��Q�ě9S�aH׏��n�m"5"O*�y�fVs� ��!��ca�@T"O^hzb��eɎ��\_�T"O�-��
F0N��d�%�T�!�y�r"OXа�Ț�`�!��(��f̀��"Op���aզ5)���GD�=��|��"O�P��$� ݈�$�8%����"O���#ɥ06�E؂�*�&�3u"OԴ����5R� �2a�Z>	���W"O.�8G�ɨ}H�������I� ��R"O�%�Tj�T���D A�u��p"O�e�2�
>����O
#`T��"O��S��G~�0�M��b3"O�y��ɇ:��A��쌘�*\k�"O
)C3J�� ��X�W4\�Հ�"O�D��NJ�+)L��R9_~Ѹ"OP�F�J�O�����_}�����"O(�BҀ|cr��AVKUz�s�"O�8P���nl���W�xᛐ"O������&m � b͌(��1�"OZg�ت.��1b`j�O�����"Od��r鎸U:h�0����#�"O����   ��   �  �  �#  ].  �7  �B  �N  �Z  �f  ?s  8}  ��  2�  ˜  �  X�  I�  ̻  ��  �  Y�  ��  ��  4�  ��  3�  v�  � � > | � " �( �. ?5 �; �A H �N �U \ Kb �h �n Su �~ S� �� Ց �� \� �� � 9�  `� u�	����Zv)A�'ld\�0BJz+ �D��E�2T��ƕ#Ĵ�GN9�?Y���?��FJ%L+��s�'Y<��i��V�8 !¢!�b\�Aʶ�֘=2�j��F9��P�
�)�b��IK�y�fpq�&K�l͂,�+[�X�RtX�˟/2����I�K���Źt��ƥ�y!�'�?y��$q��R)L�ƘQ!'�L��p��)x��S��C-��G#pH�`9P�i��p�T�'���'AR�'�d�B�
��}"J���䑙O
!���'�Zb���Ӹi ��((����?�	��|���^��,`����l��3��ߟ@��Ɵ��������䟐�rj�E�Aπ7}B�!	�>?G�E��:Θd:��0SZ���c4O �`�������{�����ŋF������n6�%�>��'��O����/	���v�r��ʷ� �$�����B�<�Z֏�OP�l����͟����?M��O��6�޹(`�Z	f,�UI�@�^� �ӵ�'�:7��mAڴ,ћ6�',7��%Mpymڕe�~yW�(Ѱ��f���w^r� A^�"� ����h�DT�E冻/�Re�0\�Y��z�]A��#rي��'���:��z��et92C��
<�����要��4L����O���	�Dۃ��;�\�1���!k�qQ�I��ؾ6톫s��5� bT�R��-���${n�:�#?, oZ�M�ŵi/�`��I�<@	�D�?6 �E* �I%F$8P*ԩ6��7��)bڴ"�
U�M�ు�SAOd��S~I�EK��.Q)���;'0`�e��Y��(�i��6��ĦщR��[�P���aI/=���
�_Y7	�44"bȅ�P�M.��b�i ����K�� i�,ڰ�E=\|~Y	d�'��Od��@Q$�@��AN�kr�Y�k������OD�D�O��I��`	��E�B���tk�Ox��j�S���h�3��\��
�Oʓ�?a��������^YB3�c��6r�i<Ш�SBh�H��.�]�]SR�'��3���(g�bM���
j�����_�
 CSNU�qG�4JR���Z�`֯�,��)�=�w`�ߟ�1�4 ��	<#e��P�Yd�E�D���(�h�d�O���:���O���OL��g>-�t��)����I/0܍�vm%�OZ@oZ*n�΍!�
*)��(vfϹ{.��޴�?A·i��QCS�~Ӓ�D�O>���bE���O�$s�U�t��=P@�м?��U���O���\�1z�͋���XR�$Ô�t��˧��	ٶ��Pe�I$�ȲՈV�A?Z�6��`�m�!�(��
-� �b�ȁ`�����?]7��8}y���Q�D�@�(.?��֟(�ٴ�>��'1H���c�l��$�әUev����F�'Ԍ8ZA�`%��� O�oR|H��d���y�4��O%��3S��3ߦ�7�V!��;���?�/OF ���O����O&�D�<9����1�Ā/Q,��*י"�p��+kmdu+�&A�	��Q)�6��� ��UR�(��kf��SD���=,4�𦃄*B4��U�i��)b�eE&�L���R>a�(��!� �ݒ_mn ���W�jl�ru]6r�!mڱ���W�3�b�O.�3��F7�X��c'�3SH4�&�ۥY�����Oʓ�?9��L�:V�V�>\��
Rp��W(�<Ǹi��6�4�4����<9ĥ8��x�K��(�Veʔǌ"g��X�W�@�I��|�'���|����K��ȃEN�-]����sFZ�I����%n��L�����<�%+��6,q���R�0��%*WKȍCK�uڳ�ؑO"%#0�;B�Nd�ߴw�ؚ!��x�xly��K��r�Y�HQ�Z�&��#I���4NC���?�' ڛ<�,X����LY�@�a� �?����?��>�X��Ug�=/9t��F���8�&�
޴pC��S�\K�d'����O�|���݉w5��je�9w@�1e��O���J�a{����OH��]GFD���!ˏ�0�o��m��v�v| NM�Tye�2ON2�垝cT�d��2{�v)˲�,1	b��cм�f��*el �ѧ�.���{B����?Y��i��7m�O�5Qf<�`Y���N7���ʫ<1���?���0|���ʐ!���aÓ
v�*!�sh�y���kٴ��x��c��< ��@/�M2Y��i�ɴ��Ģ�4�?i����L��2a��<�e�w%N͙Ы� F�����O��$EX��ȭKW��2W�֠��C����X>���ߤS L��5bZ�.�b��L�v~b�I,x1"E�ve�9[H�w(1ڢ�*GCї@O|����OzV���@_&[���b� 9�`l��O��+`�' 7�I�|̧Qgˋ�;��p�lCi���3@)9�$�O�� �<��ϒ0K���@
݅� ��'py��ݖ�~��i��q�Joş,��4�?�Ǯ��	pl싰�@9��� %�S2e훶�'Z�I�eA��ǟl��ڟ@�'��G�B�d���ŏ@y@�i���`��*��s��	�����˧|��OZ��Èy1P�,�49����,˨YP@�1$g�,��Q������Ȓפ�|�e�	`&���;>�(HK+ؚlf�Ź��V��}m^����:{>�d3��OD���O�,�t��g���j0b�S0$����Oz�d�OH�D�O��?�'64@���y�6�I$n�04(/O�1nZ��M3��"U�v�'����OE��+8�YA$=;���������	�0@����� ����Y��<�$�O�AP��8,�*��L+|�
��M0<�%� F�%;�B���ć7@������I���%��.
��!Щ��ৌ�,YF�|��cK�*B���	�~��l�ff��>OP�O�h���W�S�6��k�2F�X fN�L��%� 	�.6M�O��?���<+O��"S�P�\��P 2A&P*���f�,?���1_��Tl��?��	�<Y�bM�OS���K߷m�:�)���Vy�'H6��O��h�<�Q�iq�'��y�"	@1���B�@*
h�ѻ��'��&�+R���4I
+-)1��� �h�W����� VH����4�f�@<b:�at�H}�'����k)[w(i!�'>g*6}��,����qi�u�`�j���F�\qP�h���E�ĝ|����?��i���Ft$l��] @�Ĝ�c��
K�d'��EB���	�Z�cj�rF�r>�Cm8��~�����n��t�Ӽgd6d)�&+t�=�&XϦ=�'����%�iӘ�Ĳ<�)����R�O��q�'�Y�E*�P����W����O���B�E���+�y���lw�'O��9X�͞�"p�Q���n�k�On����0T6]`��S%>.z}���!
g~A��S��d��O*81#��ۇ|�z���)��[����sӸE��7��T{&`*m�2T�G��ȉR4�'�O����3X��}3BbU�}�=���ٵ�0<��4^,�&�'Q6�x��{�`ǖ �n�1���I֞L�V!�����I��P���>N�� � a���	���	�#��n�8��]�p�0�NV`y�'�@jǡTeX� xA-��tzp���	XU<�P'������B����M�q,��#���|�<A��&O�Z`��厧cxZ� 2��%�MC]���b�ON�I0&�`��J"��6T�)c��d��W�'Daxb��sf6�ja#��I���	�)����D�Ȧ�0ܴ���|��'��$6,�X�A�N�}ȰE��j	`8C��������O���O�\�;�?�����i	��t�"s)\(�8d㖲h�̜.?V.-��̏8d6\�R�,��O��(GƐl�Ӏ��.9P�[�N ������U8'g���昧/�6�?i�$��� �֗YK�bQB/~�����?���'�>���3O�f蹕�XiH�u�VH<D�\�gꇒk�zqSJʺ9�P��;��Ŧ��I`yB�	�F�*6�$���?ꤡQueѦFaz��🨕'�r�'��� ^T�X�o]�}�\�NX96z�����R���i9���]S<u�HW�'�Xՙ�hF���L둯��`�d�p��
 �1� ��nyk�Ŕ�5�b �2!S}�s�|bA�?YD�i~ʓR`hE{���9q{&ݻZ�*�%����='���Q�=t�h��G�j-���'�O��m���}Ȏ�-�h�p��g��I�۴��^���<ߜ���O��'�$���+݊)�P$��M^�=:#�:�8���?Q� T8p1���'+�`��q1L=���^����N %�J��e�� jC�XJD�((��b�^X�!Q��X��)�d�j�k�%��O�r�yv!�!]�Ȋ�J���a�O>ԑ��'�7m�p�O��)Ĩr\����n\Z8`p��&���)�'9M�1KV��	hF�i��)lD.���M���id1O����e
e� �J�c�-�
<� lyӠ���O��D�O�i�'�O��d�OT�Dy�q��FD� �v�YG�/ ��5����H
�DЎ�Ʀ���F�]Z�O:�⟨ӑ/Tv4T��)R�<*`�
�2<���a'E�0�b] ��@��D-B��~"CA��Yϻ��]Ǫ�&*E�1�5�L�
ͳش��I,(g��dV�w��g��w	D1�M�8t�ԅǢ�R���?�+Ov�D4��N��e 3�"-q���x���!e�b�'~����|�����D��S�cp!O0lul�SQ @<2�q�Q.@����O����O:	���?�������K�|��H��*M{���G�3	ܤ�lN˲���]$��s`@�B�8�Dy�n�| �l�#��Q8�5k��۩5$.�"��J+�5K�#�.zM�$�,( v�p�%)cR�''~�X0��m	n��%፜�Ƥ �D��?9��'w�!r�h�#DX
)1�I�<;��݁���'<Ny �Qfje
u��>qf�[K>�i�'ȮY%${��d��X��b�-[I|�,[lz4���ay"�'B4����V'7���'��9+\7�R�C���Q̑@��@Q�i��M�~��LR���&F��y�c�!Mi��H"���� �� �԰Iq�hw��p����(���'�jp�T����<�aQ�W�nI�*�ig��:P��K�C��sg�1JU�@�䀪P� �QC�<�
ߓ
���@oX]ց���Q#�> �6�<����N���'T"S>��� H�P	X�m+&A�c�)����F������ J=��4����>a�J��YBl0z�(L�'Xu �N[r~�-�|z��s)�,T e�#&�'{y2q`�߄s�r�r�ƨTY�@�'�2����+��&}�<��㟄Dr��~Bq�C$~��M��A-�.�",�W�	Ɵ@��ɧ�T�h���%� 0�菅 ����<a(Ok�iߔ듆�dk>9HƦC���CA��c;(��b&�æ���ҟ���7�fLsp�ϟ��I�<��׼��-v�N���"��_]�ƍ\i���AOl������g�,�b�h�f���
��IO^q��\�G�Ei�n�!�"���N�'̉'op8���P�4�Ѭ9�"�ke�T&Yy���<i5����h�|�����u���k�V<`���ʈ%�6�D{��'�Ȁ��� y���g�ۓ)�#,O�nڌ�McH>��'�z*O|����L�`�ʑˀJ �ʡ�M!6�8��!��O���O��������O���Ͱ����GKَ9�`u��E "r����ǳZ�LY���'����� ��4�X�?�y"BŻ7p�1�ġ�;s�E�3�ӛG�zSAPM�'�ڙ� ��>R�\B�b�8O\zp�Rhʐ�?9�P`�'��'��ON(K0J�j��Q%Пi�f�#ړ�0<�0aڸf����d$љy:0x�&TG�I�M[R�i+�+&Wx�y�4�?��f4��P��+��싑!��$HD1��?q��N��?!��?A��ǳ#қƓ|�dQ�;D��6L-pM�VH�=cfaxb�%H[z�C��L,rv�U���k�Pe*�@Y7&g���&+tT*D��'˸1!��L��fmaӾ�� 3�V�H&b��ޠ���ǂl��d0�^��.�)ʧ::�l�ԋ��>�1����(�,��'��	�D�TL�On10t=ɂ�����
#�DQv�'�	�"՚�P�4�?Y��?y��_��0[��En�S�b�7!��Y�n�1`b�`��?�BED q���a` ��4t�zbD˪kF��������b�JsGlY�~u�Q�Z�0��&k�8��Ě�v3�X�7�ؒQ�Z���/��r�ʅ`��?I��j]�H���+ˮI�j�=?Qoߟ4��e�O���ܿEҙ�WD�?$<��ɤ@B�x�!�7a�6�c��o2�y3Џ�7l�ў ���HO�9Q��ɭ6�Id2<��$�5m�ҟ8��͟�;`�($�x	�	�����X�;|9�|��&ÖK؀[�� CԀ'��kuɎ���<�����q��d벌?,�bxj�[�pO��z��E+��ƀ_n��B���yr��(35ȑ
w�^�H^p�il�7.f�Fne����ӗq��� 5��O���O��20�.z4�����mT�]B�4|O���y�-[���%IJj��(BD��?Q��$m�Izy�V>U�	Xy�İ����C��3��SOݟ0�δ�"%Ύ<��'���'�D�̟L�	�|�!d�)m��AwG� |�5��*^*M����F�GW���K�h�
�4�ٗ.��<i�ř+Tؼ�)ßXx�:�mY�-����RE0�DԩGI�D�~��l�:� �k����9���wgU~Z��0T�
m��#����Iz�'��H(�.��v�[�m�,l�%�b
3|OFc��#�,;���afL8�Nh�E�6���Ǧ���yy�h�6����?�R��(?���8u�,QFxE��l͂�?q��T��r���?Y�O�`��C�%` 8�T�C˼\� �H3$��!�DOU�Q�h�(7a�(�R4�!��y�'��I���X%f�(��ǖ:���"
�,��ٓ�OM.*��!Î#k�,ja��rǀL=��H�0��I��'t� Q�a�/������A�>���K>a�A"�,��lҶ���W p8�|�?I��4�@��	��&1���Ԫ��5�%F�<Z�@�D�<q��r�V�'��X>9�G+˟xJ��Au�ءr��=�n�cTD�şT�		;Zx�ش����>Q0��p�2YcG�E�@C�N�~�����x��iӢOf��;�0�'�rU�@�И�	M!/�� �T��}~"'�?�1�itL6��Oh��O(��6|��1d��W8|ї�٥8�l &����l��\��gT���R�
Zr��� B����D�<��+Z��ty�1�YS�H���i5�[�A���jEHq����O�ï�`�Ơ�O*�d�O�Ds��B���t�D�{c�B�l�~h�3�7D����d�$���V�Ŝ=>b>��Ul�
s�D�?`h��Pm��/�-@0bB`xLaQ�K�1�J�Yb��23�@qGŁ��'Id���\ܼ��ĕh�h|jrF�
N�9�P�Q
��M�-��`�g�"P��c$)N�s>�R���k(&Ņ�9���:�m�'�-���d��I����4��O"lk�n�1T� }P3b"^�1��, �f\����OT���O�������?���#���U�ʰXo�0Y`ιt���UC2��J��'��KG�XZ=��]#f%:(Q�)�{D�8&�N5S(5�e��0<�3*G�qT<�2���j�U!W'Y�ܐ�I8�MC��i��X���	H��pr�&lQ��Ԝ�t�=�
 ��x�Ñ��<h��µ=�p��D*���M��v�vӖ˓G��l[��i���'d,�� ��af�0i5��Q��'"*R?���'��)F�[��Mr���7�Z�V,�O�|��͒�)��(���ƇQ|r�z��'�"��G��'S~��p%ًDnp�6:���B��!�z���Px��2@�=%}�=�ֆ�ß���Z~rO��Q�0I�-�"�nE����䓡0>Q"�?_V��Iю/�Z��F�����b�����Z�l�ظ�Q�A�L���Jy�AH.~�"�'aY>�2�f�ȟ���D�.&��9�(� 8����n�ԟh�I��ڭ�P����ݨ&b��?�Ox�S�?��C`�0��0P��
0К��C�'@0�@T�
�Hh�XKQ���4\�P�OI����E�b��Ik�Ҥߖ���O&a���'r��<��@O�jM�]�m v��P5�u�<)��V5Z��H�"�B�x����%�x�'*��}և
�9C�M�È�>8�2�(��ȟd�����Ip���H�G
���柔��̼�T�	�\���&e�P���Fz�
T�����M�	�a��]Ј��y�H��3m���S�=Sܛ6�U�>�ti��W1Ǜ�@L�s�:�
���ʧc��,�ļ� ��{�`]���adƐ�q��Mj��'9�I�"�X���O�=Y@��؉�(�$]T�@�@��y�Y�'���O�����7�?9�����˟��'�K�2���jd�&�©����]��e����?���?Y�����O0��r>�UKK4o^d�Rl^�W(DڗˀSD�� ȏ>�$�0��G���i2�ZoQ�(�3��)kD�4z�&6D�E3��K�n9k��źqlM#�b,(/��lڰS��6�	�l��'�L�AA�K��11���k��i��ב�?q��'1tD�"������0IW�9+�9�ߓ��'\L�N�k/�u�&�U	fi�e�I>iѽi��'_6��գ�~j�� ��7%_�jJ�� F�,\�rTh���?I��=�?�����4�R PV]C@W8h˘�A�(LJ���$���p�����c�2�M[@�1r�`Ey��D�td��e�,d�r���F�蔯z
�"F�E�p0`G�3�ġ�B�i4��H>y��ȟT�	P~b�V:�<T��OU	�����+���0>!��(7N5����0a"�z��hO���,p�BK*~�-��* |*��@$�O�B�N�؂�i���'��S�v�t��9n�	�&��	
]�.�>[`�%��ȟ(��&�o�"Q��+Zy���(>o
�����~�4Uǲ)B�b'�i��C,��	�yX���T�4
@���Mԭu����G�& ��'* |�S�Γ� �2��D��6gB��'�e��/lɧ�j�F��&h������#�""O"�K��@�g��m0K��n8���ɍ�h���yUo��}h����P@L�9l~�����Or�DRplD�ش*�O��$�O��q��&0��YK��P�f��B�z3��z�).DN|�	�o�Q��'��t��+m���#����l�	x �E���D�[�M �E�4�Z	��x�$��_�';���u+��lQ�&�g��EX���b蠈c�-DV�I`��D9�3�		q' �P�A��s}`�B���q#ZC�I�3�r��L�PM2�B�GT; T˓O����f����k��J '���)J85b�%�D������8�I矬bZw��'��iU�V�Ft�R�%D'zX�A`��^���d�A����MȕJ�ؑ,�"�����	N\���jY`\K�=l#�x �-Tb��G�8,�re��
��} V��6�(ODys�(	T4�ۥeG/ ⽳Dj��_2�#�O��zo�%HE�@��[7A��"O��+a��
�.Ș���yy���� 󛆗|2aTU��'�?��	ӏi|�T��-���M�>�?��\ (���?ћOD� ���5K��B�ˆ$
��f�<Qf���'ب[�N�C���ak���F�'K�ѻ�٥I����`��C�qJs*�U��5`3eUV�9�^�<�*Q*&��OΈc��'�R���bc�k�J=���8��Q�.��5�O��&M���xHӱIp�h�!��'4�$�VϬlZ��dm�i��h�5,�r]���sC����	��<�Oc�0�r�'���2,�9!Ҷ�Iq���>�lXzW�'�"l��.>�0����S����̖��|@2�J�	���O��D2�F�e�̥R�#E.w�����=2F��o�-�7�{�(��Y!f
����	�?]� imJE��V��9�k=?����$�Iv�O���<B�=�N�*��qQ.ѩ'�!�$C�Ҋx���_0%���kT�2`�џ�Ѝ�i��>�P�Q��J0����V��|D6��O��$�O�!S�e��Hp��$�O���O��#L&x��R�TyT�)6�ÙH�õ��0����{w�As���U�wM�i�ԭ�1hA��#��uł�~}B��#�b�����y򈄫']�\i�JQ7Jtx� bԝ�?��O���u�'����}u�P�!{�-�F*�qO��ȓ�|"�����5��D�:�(@�O�xGz�O��P�D!��Ʃ68d��g�M���IP���`d�G蟰��؟��I	�u��'a20�����dĔPzb��G�G`x���j�<���T�
�kj�xcJ7S�ޢ?��e�}��ѐҨO�XB�5ёJ�+� 1��(��R�3�"X�*ۼiБo\Z�'�E��V�`8��\ݒG&��?��?�����e��m�SO��m���2�\�&tB�I�#��HzvES�o"V�����O��mZџ��'Y:�(�/���>���S�/�V�l=q'#یT��X����̟h�	�O��@�W�"hoLY����?1��&.��*�	o:�@Sl�e��i3&ʯg1�yR�J�T������F�DK��	�n��S���?��Ě*o2�'*�I���3W���#M���3�� \��O����M-t�<�'�"��!�O:4����Oف����M��L��n$C.Y�S�'��	?�M�����|*��trT%`��M�+�B0�f�
�w��u3��?9�	[9t� �.Z�q������xcT�߃H�(	��Vi�h�◟k! ɶ�
IaCY�iF��
&LoH$�s�I$�aV�^��
�H��'Z�>��S�? ,`J�� /�U��I�%~��� "Oҙ��$�?t'ȱ���[�2����-�h�t���!ٗ'��铋8�`Qu�'�l����4�Q���e-Hj���#�c��3�=D�TB%*�:Zr�$�.Q�a�^�i�E9D�K��R%_�楃#P�.�+cd3D��B5F��7Ř�
PA�?�v�!��1D�<h �F2:��җkK!P᠑�)D��Ӗ�V(,k ��	�"��󤩧<��KAY8�����Ä��_���e�R�8D�l)�nؚ~$x��.2k��#�7D��
!�4=z���w���/D��E �z�h&��H�TA/D�b���!$4��U9VPD��q.�O�X0��O y�˔�o�*X˦�_�Rx��"O��1�
�k���Ec�O�j-A�"O�1��O9�^���h�;;�B���"O�g�bjI����Q^-��"O.Yr�a�I�@�DD�GK�Бe"Ol� H�1	<��J�E^�W�6����I�|dȣ~��W�7�<+$� �n�I:�͌i�<�aì;8����a/x��/Ne�<ɢ���:!���ԯ�' {�p��^u�<夛� p�<1v�ʧ!\��o�Z�<q� E��� e� $����ec�U�<auI�OQd��`�i!�Xc�� �)�S�O?2D+�IJ8׾�"!xɑ�a���y2g@'x����݈61<�s����yRĔa>���k�zZ&ljrbŪ�yr�]�#�f�T�V=:'���1e��y¢D�T3(��!8)���ݱ��xB
J�Y��b���9W��X�
^�C�F��5��!�M���ֶ�p����l!d��O�8��b�O�N��*�B̒!m�< �8q�҉9>���Ծ���O�����=�B/%K �Y�/�9Lfݭ�d:`�ϪD�����:z�Hl�6�[K�'`eYj�"sg������ M�H�[e�� ���Ȯ=_��&g֜b!���#lY��M[���:��7�t��I���|Z`�ǈ/u�1�3%�-V#<���ky��'Nȹ��A�"�%�ҫT��R
A��i���d��<���/��
Vk�#�8pRW��G~R�Q�?SA�?�,�XP����[#\�|s�!��
T͚q'�o���Dͣ`j��[��X�	?�ِ�΄#.2讻r�Y��$)��O����OLFp�4o�y�t� T�,x��eQR/"vj�n�8�ug�I$}�品c�< ��,M  ��e��	�A�
���O��S�}~򂘱%�(�*S��Ewܨ�u��y򁊑9p;"Ē�j��l�4mZ��'��<��|�.�=��}�@B��Oq�@;4&�lp��?!C��R�!�'�?���?�4���d�0w�l���^3)p8qx�@V�J�ڤ�L,�>ɛB �'E���$-�ԃ@�9!V�'���Hu�d���t���\D,(�f9¸	c] @�A�&���哗B�aR�ϚY���JF�}����%��%�nCO?F�H�Q��؟$E{�5Opp32kQ-$HF5b@�A�=�Ovݡ�����1�rN�%&��sI�O�lDz�O�2^��r�/�($x�L��};1�7e&Q�Ě�N�>5�}�I� �I�uw�'��:���A�!�̍��i̼(���F⚢=� V_CU��ta�^$F��P�ɬ=V�kU���(Ђԁ���YrAY�16H�C��rk�A�rk\�|�c�e����x'��{���O ʗM'��*�[�!?>IVE�O�=���D�)$�4H�b��Y��]r�)J�~<�y��I,>��P�B�_�~�q�"��Zddʓ ��V�'��I�g�(E�ɞq�ڬ���|"p�ʀ	9֤�@�>I�u����|��Mɟ���ܟ\��%��WW�,�B�>��q�v���u�.O�q����WJ}�}j�%��<X k��H�|��A)[np�#eÌ�+��]���@� �n�jM�s��P�H�C�ii��; �|r��?����O� X��L�#f�!�p�{)O6��$�(P�h\2M�Pf�Š9I�'�ў�S��� z���'.N���x�!Z�(��	1-��y��9n\��Iv�$�D���'��DYB��j8���靎[։�C�'��PEf^��i��F�3	JbD�qoo���eg�'9��� �;G���"��/�6�ϓ)�
��ʢ�h���Iޤ
�M0[w�����*ā)�<$GA	������$bܲp1O��9P�'�2����$�S�? �	N+K�|��d�$ ʴ�"O�9"�G�0*�9��hL<n���3��D�O�IDz�O�����ӺL��c^�+t��C�fT�"�'�Rt[�oY:g����'��'d0�䟌���Ȗu4xۣ�H���A�mD�9G�$��*'{������
g����O+*̠���X��U,7y�����#\�j�(`�@[d�us����G��9j�j�%�&���g�|b��6mWJ$S^ļ;��+n]�S �=k1��p7����|���}��g�	�<)�ȟ=M[�i�'M��?a�C�_h<��KY� ��cwc�JV�YS���?���i>���qyr��7CJ��C!Z���%ջ#W�����F����%��'Gb�|�i����ͧ�|P���:*
�#`XuQ2���Cv�Z���`nƝx��su��)�o(ʓj�n �Cf܆3�Q�sg	�<.8�Ӂ	"lE�,����38�8�bE�sZ����Ò ����H>����ڟ�2}����+��!�2Q��H��M���X�')�)���(2��D��y��a
ϓ�O�acZ9G8T|�s�h��[bQ���4�?-OP��b.��!y�����D�'"�#�I�M��e�D�J.W����#O���	՟d���cФC󆄧]�.�pǴi�����O)*��1��12:�����h�F쒏��ƚ%�R��-�Q���ȥJB�i��e;�t�3fB�(�`C5+G?�PP��AC��I.���BIl�0MlZ��ϧn��p�1fC?���*��)f�b��I��I� ��C���Đ9jڔճ�J�N{�53��X�ce�������`�4de��ȴ�Χp{�$hE�å)V�	3+O���W��%�����I�|��ԟ��'+�,����A�t1� b����'���)�y�"ғ%� S���ndF�6  ;x�L��2��h����~b��_:)�,�p0o	"�.��&�4ћ��'�)A�2O��)s�'4��O!�=O��K�ܯA(�����+\n>����Ƕ_�R6m�O�b�"�O��I^���s��.CB�wզ-!��Ժg�A�IT��(Hp�矘�ɇ��Γ�u�'�"�O�b�OV0QG#0�y1&��I��̈�D����U�E�4��h�N<���]gH�d�		ΝPAcU&Sx��qȒ����d����'�,�8ь�O���ǟ��I�?���s�V�R�b�81b�E{��y	��"(&����@��ԟ�!�`�8���}	W�"Szhc^"*+.h�f�A���`�4�y�%��?I�̲��O�"�'u�T�����)Ҵ	ΎpО�"�N�z3R��0:O����'I�'eݱ���<a����شQ�TuI@gM�'�lSd��Ug�%�v����O�s2�'��@�	O�'�?9�#v`��uF�0W������`��)h7�i�ʐI�:O8�5pӌl�?��Ʌ�?y/;�JA�_y�N��ǎQ��`Pf�M�r��r�����>�p�Oě������?e�G� �P�Z���J��KԠ���G���y�`�#�fi�����2��,B��A�M������O���O����Or���O|ax �D�M-&�AE�FF�w�Ц��ޟ�'��Iȟ �I�@�ɉ&,q��B�&J�x+1�̢N�"�2�4�?���?	���?�)O�I�O:�d^B( acY�n�i`��]�}�dl����	՟8�Iߟ�	vy��'o�dVEФe���h�6�����jx�|�'3�l���ց_�+6��ez��r7)1��?i+Ovʓd�Rx�U��5�uc�ʜ
�V�ؗ'4�	ퟤ�'/�i��a"B��	��i����AV=�ȓ]���	D G�"Q#�F�+ѲY��D�ni˥�ܗ`���Z4�G.-h)�ȓaI�0�!�3�.��ь��ž��gC�Xr"X�m�8 Ea�',�-�ȓA���A�/V�Ka�$WE�8G~2�'���'���'t�	�F`�Z��
��-=$���MS��?���?���?���?	���?q��?�hI�j�\˪����R����'���'���'v�'4R�'��Z��M�a셮it�J͓Y�\7��OJ���OD���OJ�D�O��$�Ot��ڻ<�P�Ô��#c4L�h��"�n����I����������ȟ8�I͟�ɫr�L��R���b���Ai�Xݴ�?A���?���?���?���?��U��z��QJ�؊�nMRlq 0�i�"�'"�'�r�'1��'���'�b��䨎�;+�E�c ��lHP%�$r�R���O��$�O��d�O���OF�D�Ob�!*W��X,W1ʼxq'�'���'N2�'��'R"�'z��'e2�z�Fm���O���<�A��3�6m�O����Ol�D�O��$�Of�d�O6��٨84؅�S@ �f�\h�Fˎ$E��5mZşh�I͟T�	�����ܟ��������P�&ͪ�+ݾwt�(��ӓx���ڴ�?���?a���?Q���?����?��9�0�x`�X�*y2�Fπ+s6:�	��i�2�'�"�'�R�'�')��'R��1#aMI���!�i���H_�M��O���<Q��)��o	9{�d)���A������7-�#[+1OT�	!��F���λ�F=�։>t"�{�mT>�q���Mk�'M�)�)�/B��!�ON(�7ʃr�H��5`���`�'�<����^,����i>]�CӸL����8.�Ľ��KZ������Ty�|"�w�ۙf�d*� �Q��-ST怰 gM���=���Dfyr�'r�V6O4˓lF�ݘ�@���3�ϗc<�'d�3���.�����O󩍦>	�p�x�ĳs�M�&Fl �b��
o�P����<)O���:�g?�+@,;�H �(�nNHta�D� ��4$���'��6-0�i>�� ��L�E�)\&Ny�W��<)��M���u�$�C'PI~�
�=PK��*tj��[���H�h�r��Xb`�5� ��d�'�bU��|�¸����X�E-�)8�Udy"�oӪ-�b�d4�S�.]`%ɖjȄ-�0(#�%;Ne���)O���h���N�O�X�3d�;O�v1�䅅95������"m@}��Ov�aa�(FWҐbw�<ړs�	��Lׁu"�@y��H/������ĵ<K>�d�iL!r�'q��'�U�,9j�T��;I�X���H����'�ɧ��'t��iA�ό"��H@�5�x��q;�p�IҤ_�y2����胓&O������]�?����X.d�3É�i��d'F�':@�	��|�'X�)�'K��]:��B��5��i�C(A&���ش%v@�'�6��O�� �N"�Nנ;�Ț`��3b��$���Db��oZ�<i�	�:���iݡ[s( ���)W��E2D��#	��5�Z<�Q	�X��[4�xR����dyB9O>�����R�D����� ��pd�'	�'�,6��'^11O��':f.�ӂfG�&X��P�-˼Q�'���?�۴�y��T�O�|	 T%Λw8F8���Z�C�U�����C���P�D�~¨C��u'������p�'9��V��q��a�\.0|+�I5l��|�'5�]�x'?�w���]�bf�ȶ+ץx�ҔC���+���
�O"1ln��|��?)�G�Ip(��D{ ]��d�$�M+�2,�y97cO�<��$22��V�� 4� �'SL�����d�H/-��ʷ�'��I�����ퟸ�	��P�	ȟ(Χ ���CA	Y� YJ��J悕x�4D��-#ф̟�?q����i]�<��R��V1O��D-9X �"�!�A��)Ki���oZ��M�0^�D���?��S�k����G�u�P#�l�K���2�ռ)��Tğ��$��<����s�Iߟ��	���	�zNzr&D�3���%JG�~IZY���������M�-O<n�)2� �����y�XU�&Uԥ�-�*q�"<&��&�Ԡ�4T��֫�O�7mh>��l�6���A�� �D����OV���N��(�F��	a�������]4P"�!�''6��uƀ%u��{7G*<�	���?i���?����h���]�Ať�M��H��"7���d�ɦU�$	s�H�I؟ '���<��O�6<qXt��D�C"ӟ�q�4i囦�d���#`�X5|���O ��� �	d�TS�%�*s�tI�Y���
�M5�Z�+*O`��O��$�O$�$�O��d�O��D6ESf�8$MN��<�贎�+V}�!�fG�v�Ld�'���?��q>u��"*]r����&/\Ěү�<�0�i�\7��|oZh�d�Of�$�Ø��z���p�蕺�P&5z5+���'3��I�B9D���:E��d&���'�����a��̛��CI6����'3��'A�'��W�āڴ4�\�͓=?�ts��	1C��()b��r�
0i�t��DP^}Rnӈ�o=�?QՏI!oF�Hr������M[
���6@a�����~�P�,C m1F�'���������/7DH�ݗ`$��%�'���'9��'E"�'U>�B�kL�q�*��AmQ�ps$)�O��$�O(mZ
n�(�?]�6��5��t{���fX��&��������>���%�i��D*	�*�"�O8R�@�R�l)��� R�Ep��&�$혔N�#1�ؒO&˓�?y���?���z,4�C�"ƂO����O2��x���?�.Oh(nڧ��	��0��C�tg^�c��y�a�5�����AH����^}�/eӲm���?ɋ�dL�&��x���&8a0�`�+Ư'�$�bjC5[j��(O��	��d��1#.�	�iۓhԼ&�܊wk�&�r��?I+Op���	�M�5K��)AR�I�,׏,u�$��\��)�'3 6-�OZ�O��Od�$��}�� �F�$DdA�6Oҙ��6��O����U,�$�OLw���a��X���K�r�>��7ؔ95���e��k�ԟ��'L?q ś��x��r��s��i�slTæ���G:��?}'?)�ٴ�yG�[;*���t#�nn.c��Ǖ,���i��<���?���6N������P�O�% Pt�X�MJ1[<�.Mӟ4 ���Ӈ�Sj����4OB�9 �[y�h���K�/%�4M���'��Io�I��M3F�T�H��D	A��8$�ڀ�%��)#�i��� F�Iٟ�nZ�<!*O^=�t�lؠQ��$��3���A�'+1Y��!)Bcܓ��d���	s�9>��	$8�x!D�:L}.\5-xl�ʓ���O��}����&��<�^�5�C�Y���	#�Mۑ��J~�k��D'�4��: 
r��\1��\�\��r�x��l��M[�k]h�CQ�H�<��Ip����8a���ݦ�����]̾h)`�уg�b�O���?���?����?���!�-ܴ�[��A>.�nr�f���dKĦq;��p����џ�%?�Iu=���`)˪:٨݁æ �4{��x�Om�5�MK��'��>Mx�
�Zd@Cꎋt�%����cנQ�1��\yBf"M�ʅ+�G0B�'��I�Q�$���׽W4�Axu�ȂT����Iٟ(��͟���ß`�'�7�@�MA�� dDؐ���t��Ȅ!�--V�1��'JR�|"�'��	��MkԹi�b��I�r8L*�+Eq=�!x¦�BYP8�eK�!�y"�'��S���X<D�*A]���S�5�Q�e�H��	�r$x�Q�Bv�'���'G�'�B�'1��j�Ȅ������c�h��k �a��D�O�m�A��)jH>q$n�1-���
���<��5g-"ᛆ�~Ӽ�[Ϧ�(ڴ�"!kT�=L�|ϓ�M�Gܘt��hP�D		��P-��
���c�+!B\���|2S���I� ��ޟ��vk�?,nu�¤P<L��6�ǟ���Ty��qӘM�Ԡ�O��$�O��'h�|�#g���fcx�@W�9u��8�'�P�R���ds����Ij��?��S,�`��Kw�|<�:UI�=!D�R㙳t ,��'��D��M�����|b�)|����	P�@Zr��cgM�b�'�B�'<b���Q�ؚ�4�$�U�T"	@}��ʑ)��Y�(F��$L�m�?Y�\� 3�4q1мYWb�w�Ĭ�P�X=��}R��i�H6��W�j�#>O����KQr�C��B�!I ʓt]�0���G2�����a��I?��*�����Oh�D�O��$�On��5����6��5��LO�
�hJ	�M��� `~��'��V>I��ǟT̻y!b%T!6��mH�k�$��)�44w����OV��:�'��D�yL���dG����c��>�����RϺ���?���M��\%�QN>�-O��D�OJL)������!�f� 3���"�O���=Id�D�<Ƀ�i�@��O:�I���J��v�N�ku�\["ГO\�D�<���i]6�����*�.u���TXLh:3.�(�>$�1�'�2Ä�$ZF�1R��J���?U
@eB�	(Iϓ.�u"g`9C�\��ଊ�q�b9�������ɟ ��`�O��d�%'�t�ZU��%XW~�!��i�~�Z<�e��<�f�i��Or�	�.Gܶ��
}�� �o֌8�.�d¦-�4#���n�4K?|9��''Q�od�5�Wn�؍�$AU1:� ��uKC�,�`��u�|R[����ן�I�������h�6jV,3
�gc	4B&�rE�xykv�P�Qa�O��$�O���d�k��YA��+ �uʣ��n����'��7���Y
��ħ���'.e;v ��!] � B�M2i�")��h,lJ)Ol�(S��}���I(��<���$s�\@cw΁�v ���Df�?A���?1��?����Ēۦ�!#�d���b��-kG���� '��@�S���D�ݴ��'���,��i�$A�	)>B��U�-��I����(|A�Ԉ[��I$�~(!�cM���t$?2]c,�a���MY8�+.R�%�`\8��'Y�'�r�'��'�i��h��];u�������w��r�'k�+r�r���3O��d�Oz�O�UJ�ȕh�:ͪ@�N�{�^�M��TmZҟX�ڴ����Oܮ����V��y��'>*�!�-
�J�w�A?1�&�c �L��	
",�-|<ў���sy�=O�YHD��6�I�e2~�h!�'E�'�6M�67�1Of�il>=HT��1|}����
N����<��S����æ���ħ�JօV�|�gi^�!#N�eoRx]�hq�	A(����'����z*�!�$Ϛ0@p�h��L�+�@U�/B�	�'�����ͦ�� �"l��1x2嗈��1�n9� �$~��4����OR%�dU1�$����5>�-�0u����8D��=8#<O���� @�ȼy֮*k�	�wd2�����9�hzV�f��qG�|��'0�IL�O�X�3���j�T�0�|��'�i�r��y��O��OD�7Myމa�	�<0�� #�L|XU�蟔l��<(O���O&B���Y�8��'E�0j�/^�E����,��tx�˲�'��Ea������uJ��i>)�n袜��$ܫKH�e�t#�'���iy��|b�c�>]����<kԀ5�0�>��y�kIA*2⟄�*O��DlӸ�Uy���>tR�� w��d����?���Zw�5P�\��''��+�@�zue0O�|că�%�Xi8�+�+1jE�u�'�2�'���'e�>a��n,���� DJ�,��Md�x��,�M��c����Gߦ���\��?�*�@W�m.1
��#R�m"��	��T�ܴuʛ��a��	�B���2fL@5����,@��p��W
|Čܺ��ƹBi��7kS(_*�O���'g��'
�'���'{X�mI�2� Ҏ4%4D��'�)���Ц+��ZƟ��	��4�Z��'��Y�w�Ωko��AGǧ�$P���>y��i4�6-�ğ�&>m���?%9��:3���S1XV	��!��%	s��<SeU�Pl�ȩ�W�2���O�h�+O��������z� �4'R���
�<����?	��?Y(Orp��:����2�(l�kҋ]X�P��F{&��D��m�?��]���4Hs�fg�OJ�k��%BI�sf�4QX�A���C�@�a��'T��]�
�E)��O���?�9�;1��P�7��m9|���.�h����'���'q�'��'!1�8�U��7\ Z��� a$�-R�	4u-v�8��'u�arӲ1��>O*����Q$�th ���;�^9�_�ͱ�E��?��O�!o�<�M��'��z�A�<��`)�'Ȍ�Cp뛐v*H���S��!�1���?���?A��?Y�;@A���8���#M$^���K΋_/�FS��R۴EB"Y����?mp�2�I��~k��ۥ,���@m�.JA��a�O��O
�mږ�MsF�'�vX>-��'��\Zkɞl0 �pk�'%W����˙)
���& �WyB�O���H���T5�'��u�#m#G(t���Af��84�'�R�'Z�'��O�ɥ�M� �܂��f�.�Q`�cj�Y"i%K)���Ms��`�>��ii #�%�2#f@9��/��I�r���Ge��`o������Cg����l.�ĺD`��*�&]�'Z�H��h[�	����׌@M����'��	��	����� ��A��kˉ1����C��[���/�"�y:�'J��'(7g�X����	8� �R�V�s�L禝c�4`G�W�����?Q���(�1�m��
s�F��h� 	�&v�С6�L�0l�[�f�9{��yB'��G��yy��'E�`�Q�
m����fV*��'���'(�	�M�T.�<I��?	���)v��iw-Y�9=Ūs���'��&ƛ�$|����	X�t�#\G�-���i�Я�1�?�����L^C��w�{y��O�<��u _�7����l��dn�(�TO]�l+b�'�B�'���S�<�7�R�r��]F@
:�IS"^ԟ YݴW�0�'7<7-)�I�?%�wdٗjQ�EN|���џ��ߴq͛q�ȁ�D��k��ID�H��oz��S���u,z��a�I��]��1���|��'���'j�'���'��qq�ȺPgI��0�I�n�q�I��MBN�v���Oe�7��9��'�	Ipl�b�F�h��5���k��)�M� �i�8�Db�˧���'cD��p��2�J ��aP�{���cj$Xݤ��*O�5Ҷ��z�he#&&�$�<�!��^j��s��M�@kK<o�'���'��6�A�T�D˓F���i>l�4*�L��&�2���k�c� l�b�d�����<���@&�I��M�T�i�$�D؍Bm�"��{�j!J����X����Ѷ�y"ꖡt+��8�@\ h���6O�d�%ǀ�X�I�NHD�E�x��d�F��}���I����I��<�i�m�ȟd�|zsK \�I���CR�����_�*,��I՟4�ɽ�M�uE �<�*���$�<�b��jZ�!�X�0r��a%AW� ���i��h�x�lZ�?�lk!�:O���5CU2�15B�f��Y��N�K� ��ƀHv\a���4��<9��?1���?A'2dXqP ��a(`���׻�?A����DZɦ����y�0����O�d�R�D�"6,uXP�Z"=Q���,O\L�'��6-��M`���ħ���n��FQXb'凮İ(�ԋǹ�F���`��dRL+Ol�i�J׈Y�1�<��Y�v��*fX u�c�-����?	��?����IkӲ�pϛfO�#Wֵr��� .\<`r��/��IB�'}��'�'p�'I�7m�3W����b��U�ݱ�`�oZ�Mk�T�R�z���?�a#ܷ6��Q�Q��B6ywDp����+�(�EO�9Z]���<A��?���?Q��?!͟�� `M
"誑���X�K͈e�5-s�T�Q D�O<���Oē���T覍�5���o�(����B+�1W{�M:۴A�&�O���z�'�
A�.r���͓aq�4��;4��L�F+�,���g�x�Eh��Tb�
K>�-O����O]p cP��m�7hJ5LPxt��/�O��D�O*��<���i6�+�'tR�'�:-񢂌�u��ȋ3�N�p�����Mx}�Hj�6Lm���?/�T�#�蛳�&���sȥ��'�o�)z�n��C�ܦZ��I�?���p�j�ϓ
��u����/�h�`�c�ty��ş���ڟt�I]�O����'�x�`ȣ6z�%���I�J\���;G��EO��y��'�$6�/�4�t��O'&m8U�Ǎ:
��bC�!d7���D˦�
�4[��mƃ�8y�'���@?�L��, M���X�I5��G�V<.�#Ǜ|RP���	�����ӟ������3"�H.W ͸A �I���@��fy2 o�>L�G5O<���Od���d_�<�2A$'jD��/��+�Be�'�6��٦�����ħ�r��:�Z5T&��)����$��=	�ɩFٔCe&�)O^$��e�9�	qH*��<�&L�z�K �ފ-n|8CUǴ�?����?���?����dȦ����{�@e��&�x�U�"����k^�h@ٴ��'p�����@�<Q��/ݚK�(�#6`V�� AO
f�"�B��y��'��hvH�a� t"�T�@��-���p �PL��:T�χH���R��ៜ����d���� �IHy��,ݧI��Ga:H�^p�
��?���?E�i�Z�#�O<�mh�`}nm��*]l��p1����.���?��O��m�.�M��'H�s���<�;��e�t΅p
��Qu�U+o��p�0;�K9`�G{�'����<a��^�~s��ÈT�'
���3�Z� '�0�ٴF��<��'����\K���p��W��P0��8��$�ty"�'9��:O��0�I+^Iz�2"V<w���+�o@7h�b�DY�pUN��V����ӧ_� ���
~�&�4JC�X|���E#Y��	�'�r^�&?�Yh���E�t���C^H���Ru'Z��~)q�Oll�ݟ'�泟��IPH����@`ز����u<�0lZ���K�Y6@�ȟ�j�"C-��АU !?��*	0_��2��IQ�����?Y/O�"~��G��`a�i�p�a+�)�Ћ���M,�|̓��O��6�c�<����l����I��Eb��Xl��<�(O���O ��@�@�*���'��Gm=l�̨��mN�Tۮ����'�V��$��J��i>��o$.���@?<Æ���e�C���	Jy��|��gӘ��u�$E	6	 �E�	cp��X� s֦�D3�DMDy2�''�V>O&�MHd)5��<(�� gfV�m�:��ğ8ȃ��+h���&?���aQ6���m�y ����ѠN�^� ;�G�+�?����?����?q���u�� 4����P�>����>$�@ 0�'��7Mч�D˓xc���'��'��ī��*s�s'
Q��|���>_|2h��hlZ7�Mk��U?5��ϓ�?Y%d��4Xd�Ó,@�,h�t1��	�{Bb�Bc�$"B9qJ>Q+O����Oj�D�O���O��l5�Pa
��(p�J� �<	F�i��!��'G2�'���y�S�Z�V��+ߐO3ؕ �:[��|��6Gh����~��?q���, �QCu�%f0b ��+ʀ0�D���#�T�l��'.� h�O*_X]�U�|�_�Pz$��mB\h1��@2T�NK5�����	Ɵ����(��yy2�|�f��i�\��N�Bf���W�؂#|����O(l�s�?a��!�Mばi6,���<E��I�΃�l� �B���J@�:fȝ��y�''��хe�o��U�X�(�S�������B�DТC ^�(:J��7�ʟH�	�����쟨��ן�G��)*Z+�;'�8ݱ6'M�`�<���O ��UΦ�$�Gy"Gq�Xc�؉4��(��8�ى>��F��ݟD�'��6������Sl>Qp$a����0;uX�P˔c[E���V
�h�Q�	<��Y�-�^�	}y��'���'�"%�.J��]D�҃|�I��	�A���'T�I*�MC���&�?���?�̟���Ȏ�qjB��B��7Mq�8�F\�  �O��m�Ms�'ŉO�����x�t�S�b�t�m��ʦ8�hQ��ʂ?4dBS����?9'T�x@Q]�ɿ1��1E��&L��.U�/�p����@�Iğ��F�STy��eӦ�0p�-i���H��жY������	��M����'���+�M�3�˜b���W��#R����dU� l�:�ٰ�W!�D�O*�HG��@�CK�<��Ԓz���l�?w�R�����",��x�
)`�`�C��Y.{����'Hc\D��� D��'gB��a��g��Y�c�3ɺd��'{.a���7WР�re��20���`#7����3�/ {.xJB ]b0~�����#o�@b�f��.��Fb)#2�XIEnQ
���'N��$ d���.]hDV$��HC����ʅ�^���ǀ�qjVAk�<�nЊF�L��[��&]���Ň�),��8Z�D�O�����$����w�6�	ٟ���Yn��3�9�$��NS��J�BO��b� �ӟP�	ǟЕ����'6R�'��I4tvp_}&��blΡu�^!�'���'HbY������I�[��m��<Ǽ ��\��� �����L� D\�W����?9�ş$X� ӳA��<���?�4C������f��Y��I65@֐��?���?	���$�O8˧�M�ծ�&݂��ddX���J#$�6Z��ɛ^I���C��?�O�#�� �+�Q�dV�w��%b�"O$�˳�B�`��ËC  ��#��,S��BF.,��&�'}w���`)?lV��e�}�ɲ�	9�ڥy��ۢQ�y��%�
� ,^�M���{���]Jf�#S)#1�
E�g�Լmk�)8e�?8�ځr�)!Kq̥zE�ŕbz�mq��-C�aR�F_�]���@EA֊/-P�wG�y3��n��l�㟬�� ��85mC�~oH�1�!"����ԟ�%� ��ԟ4A`IE� ��؟��+1�`�&��\0�x��ʟ�����������A��M�.�:���x]��M"^T�K�$���h���&��Oj�dM6$�n���O0��"��)��^?�m��	3LQИw-럌�I֟p�F�?�M�,�����̗'��g�F�-	� ��a�:Z z��?���Y�x���?���?�M~���;9~��KC�I	.)>����[�?�#��Q'�f�'���'���$��|-B���圤)���!��(D}�	�h��)�	ܟ�����%?��O��dj�a��%����Ph.OA<�!�-�"n�JIM���DXy�da�!]�)���K���O��ON�
�(�!�� �3ô���n��?�����?Y��?����ښ0��̊`ǌ3i��(��
A�ҟ���ȟ���|�IƟ��	�Ex�P�"��n�2"���MY�<�Iğ��I꟠�	⟰�O��T��O��Ą�r��
'"�6h���0' �'Z.���Ov�O�I5N^��J����Iv�(�	.Dxl	��O\�m���!���4��YFA�/$Ƭ����31�"��ILz�� ��X�'-�I؀ʌ`�B��䯓�*�Is��d�Ue�3d�$z�,`�H؏�8���uF91pʍ+sb����4E]�y�&g����p�d2x���Y�Y��π16��e�*y%(���\���#s��MC�1A��ǈF稵zAO0${R�{t%JRT��tn<U�ҁ�ۡ|�p����s�p�Dv��X�w�˙f�3�"P��P7�'���'9dM��e�<�r�F/N�l����?1�ń�	1�D-����(+�z3�#ғ{|@��@U�0�0$옝sHj�ˁ�ǲ�,���.nG4a�3j��!�(k�c��0�M>Q#_韰��4<wq�څ 7D�vt`U�!9���z�O���"�OJ�XD�_4R���*��${�(��>���4��$�O���� +6�� ����,��!3��O(A���Jզ�����O�:�ۂ�'��i#zM�喠:Y��@�Y�f􂝫7��&5�	ڐ���|V�	���zO��+�O�1�kl	�I����$�.�<�  l�BכF-@Lģ��5&e\ɪ3�Z�]�����į]n��3�V>�.G�]�1mr(�geJ'}�7m��K3B��s�"lɢ ��HV�� 埧bE2�x�"O����텵}��t�ãضx5jE��d�O\-Fz����.�*�^z�jm���H�r�L���'�r���p���W�'	��'�Z�u������Q/<�9�5^C��  4�k}�LL79���r' D29c���ĄR�.�`��$��,����7���*OR�p��\%�~y�}|��b�7����%K'?R1�'������?�H>����?)�O� �$��PI�z�0��H#Q�Ѩd"O���s!MkV���@CY$	5$`SI�HO��O��+��a��B)����Фfb(��� Ϭ�J���?���?�g U)�?�����EM�2�ՑA�,0�s"ϸ<u*��0�]�l�Pg�B@�yB(oݰ}x��O��jA�CN˄N����q���`� �V����G,-�vl�bV;��'�~l���8�j �h�L���mǜ7@Z���8D�01��M �z �2b�/WN Ka�7D�h���Ѓs�J��H�-u�����`��}R!�2>6-�O��d�~�S�ӖB��*��
�(�VȲBB�9����'���';�����
�r�dU2�N����m�~·9ú1���g"T<�X\�'�<PzbK�Q��J� \�'Ez�b�Y+W� /��a�B�Ê5��Fz�D��?	��8�z ��*~��4����nU�B�I_H�*&��1w/�l� ���C������_�ē�(B�+��+F�LA�E��$z�8Ym֟���S���S�&Y��'��#�lI�t"m�!n�|Q�O4.<��U�ODb��g��?nԫ�c¹6�PQ�ĕ5��oM�"<E�ܴ=,t�#3!F�KZFu���5]�>aoZ�zd.�DHh�)��M�"�nL�A�B82}v*"-8D��Z�R�1�(P�UN߁A��%�pJ+�rX��ʧ5��@��F;$�5���Q��Y��'@��_=|rh�:e�'���'k�o����ﲠ�4��e�*������(nT`��-�h�Ig>�S?#=���c�R�(uKǀ?���oW3�`�E�T���1�F^_�v�On�$���M���4�'�u�@D�c��<��.$�
�K�O�c��'�a{�� J��Bэ�&Fϔ��E���y� Y6< Q�㓚>�������sl�Dz�O�'N�P�p$�`h�@�@?�LpW�J	<,�8h��'���'UP<$���'��	�
� }B�Ί�a���h�'\�hs`��vܜe+�m��1 ]�5��x�'� ����8}OT�hw+F�.��	�@��:�ր��%�_��t�Mp��� �Ҁb\+Ҭ9�ҁb󄙗2d�	�,Kz3~����6\_0Նȓ2��wo
}�LT8��̬2J��ȓ[. ��(��x��MP� ���:���|��Unj.6m�O����~:�!�57��Y��*�8����5	L�S���X3�'�r�'�NxYV\�5�.��$�T?�K���Y8�ș̟5�z�U�.�a5c�G7/Jl(��˃wK=/>��@�@18��	b�+ű����IB"4{,�P���=�S� O����R?�́�OV�	[�B�	�z��xU�9�Q⒄ �^q���d�m�їg��]���Xi�x���O�=>���~��Loݟ��I]��hÐu�'?�����<�	�A���z���%��J: ��h��*��b4�H>2ݰb�N8��t��ȍiV���8�jm[w �.(v�1�i����'V�_���Gc�76*>@2�LIqlAۇi*d#�s��`!.՚"��[GW�@3C%W��M+�jMП�K>E��4+����v�Z-�rmK?7*�U��S�*ĸP�ŠKw��b�eV��N��=���#ؑ���AZ�˚�Kq ��r�J�o��YVA��?��`��v�D�?	���?q��n�.�OD_0� 6��W8:M��T���ث�a}�ެ#��l*�O5y3�������:H�a}R�G�RdH��jڱ
w8�]�����O�Y��N��m�q�R����X�4IzC�	5qt]��H�a�������*om&Q��)�'2�=�W'P{8���f	�j����N�!!� ���?	��?��Q�?�������m�P�D�ƹIzl(�P^�����"S72��'��uw�y��9a7�x���ƠJ�FY�劏)<�X��!�B�7�q§�,H�(�"K�'1,��pM�{�L}�I�U���ٗ��_�Zs�Aӗ6vp"O:�(��~\�I�aϫ��xi"O�,�#��c�:���09���
Q�O��l�[��1_(2U�ٴ�?i���)X�y��`C�̸���-�==�����䟤�	័�!�UƟH�<�O0p�r��!�>��ުeW�i���S$.ܑ?1��Z�4���������Є>ғw���I��(�4����TxV�b`��)S�t��"O���0��= H�䁀Dq�+7�p>S�>��'<(@8�Xa�y�QF�&a��I�^LF y�4�?����I�1b��O:6��԰yD��P�a���G�*<`�� ��<���'_���fcU�A
��a��
����4��<Gx���i^X�N�;D��Z5oR�wy�\zٴh9ԙ��2��S��MkF֑(r;�$t���r�<� �AcQb�*B���%h��C�zВf�ɒ�HO�)z��hѓ���5q��k!�/l�9�Q�Mǟ8��)/g���4���@��ß����uG���{�М x�AIM*���EH�O}�$��>�e��7CL|�)V>c�pDӔ'KQ}����>	���f5zl8@jV���R�I�O}����?y6�'���Ŏ�N�<���T/\ \�	�'yE:5�ξGF,����f��{��[���d�|Rhɟ� �z��a�������9�p%���'�R�'���{�'�:�|��s�6��� Wc.%���Y�i٘N���v�cX�t��k�W��(� �#
���9fJ\�$���C�"��>��&�ޟ�8DA"��h�e���&��m��%�$q	�bJ<a��?��*�Ҡ�6	��m��}RcC¾,B��2"O�`����%M�I��b�.K�"U��O �n���'���תv�0���Op�LB���
9S��胩C��R���gY���'��H�|Ze�d	?��9O��PK��s��2@tI c;gcZ"=��ł�`,�҃�4If�%>���-G>N���G�rk���5ғF�n|����M��?���>TCD�L
w�Y:gB<]��U ��C��L�	���I֟�O�'뾩I��ǫ$���*�\|B)�	�)��L~�L"4b�V�>9�6��*G����Y\�:��i���'P�S�8�a�I��xl�)M�A����c��=;7N��	ު�� ?�?1�y*��OF���IT TM���^�h����it�9+���s�Mh"�-(Th�r- +�4녻iJL@��������� V1=���r�Ўa��Y�`&X��yr��t46X�F��^�������(O��Dz�Oe�ց8Y�xɨ'�N�&݂E#��V	G��D�O��i�jD�]oj���O����O�A�;�?�abAJ 叧x94 ���$5��ae'90z��%�!(�n�`AŴ~� A^�vГO�C-��Q� �"� ��G,�����%	Ԋ�ZD�����(��A� ��'r�"+�$�2zo�в5�X�	a~98��^�Db�I�kƲ�$�y��TK����p��(;���sd�(D���w�H�q,��SI-���3g9����x�}�ƕ3p�K�m�@|���ǝ>�P�)��!H���	㟌��؟hZt��Ο���|`��E��T�ʞ�=3��
�|7��.�`-XE��
�qy��۽D�Ԣ<q6̀7� �iGD..p-����=���A'�v�.0�AS�kSd)� 	��+��iT�,�	����DJ:*NQ��Õ	C`���P����3�'yn]��J�-ꊉ)3ÛA�@���'ј cj�5f���K�l�j�4��'�R6�(��;s딡l�ӟ\�IV�T�yy	�b��l��/ٔX�yz��Or���O�Q��Oc��'J�RY��j��]�$��Fs��Fz�	�u��AJ�Α�`~̉ؗN,҇�P1�TY�ꆑv����IUi�'�B��uHQ>�bp�W#ZJ�"��4{���X�I2D����"�*Rҕ�	�>�PIy�l.}R�i>	"H����>W
�H J�B���%��@� C�'�M����?�+�ʬ�E�O �ddӐ1&��bb4S��9G��m+��ax�Re�g`h!�ɚ%b�Rq����c>��d�,t2d��._�����;�7�]x������P�\nz�a�E�,ɾ��rM�)41�\cUf�	�lE4o�L�R��1E���kٴ7����	��M#P�i�R�s��<1� I)���RƊхp��ar�Ol�$3�OHM�0�W7^���ɖ�;j�D��2�HOZ�AJr�`���	���!�@�����|��2��hXTb@����џ���9�u��'Λ�&�2Έ �ƨW�@	�N�!��#��*l�ZQ	�)��`������������@��h�"�D��}��,�7��q�Gn�K0�̐����_J�F�\�b�	�V�y��� l���	�4_�x��h��,L����`����T<j�dٸ�
^<<<z-��-5�to�9>b��v�\�z�֝kC��>|���i>Y'����������tf�%,�D�ьŤo	�IUo]ϟx�Iӟ��'0
���	՟��'Lf��C�yG�E����Y��S��C^�QZ��.`:4�f�S;��O���oA�Fv �@�H�a�x�0Fq��:��WQP���ۻ9c`7�N�^��y����P.J�b"E��q�Ak׵�Q���\+
��ȓdT$m����;�Ty)�s �P�ȓ�H�2��{A�Y�IN�]D.)�nЛ�|��@(¢7M�O���~:�L[�yf��Sq쎓G�e t��c5&����'��'�DmZe�kFl�#
 �W�t��g.�?�idh;HN"D��`�&A�ȗ<���3t��?1
u�Sb�`�Xw��RD��ixX��è�c�U�GƋw4�I���+��Ɗw0��+ʧFpqE$N82fL�c7��+�ц�&��A[�m���f��#�ؾ4W~)��I��)� Dx�6$�H0�t�Ƚ`�hi�f�Ot��C���	柜�O� ��'��i�FٱEDB5}e�$��&�
.�&�Y�iV�l(�T�Td�;y+����K�R�f�OL1�k��)�h]C6)��z���b˯+T����Y��E�t'ܾb}��gCG�S~�ԮI� ���~�1%�H���'�#}Oj�b�C�	�6m�(����M�)�禍� �nM�]IU��'Q��f'D����a�	f���"�!�����y��%�(w���ܦ�Sb��q���]$��E:�G9�?��tL��Q�� %�?Y��?��+���OG%�:I�ĵ�v���X�b(����OT�Z��'�
)�KC� ;YAOU�0�P2�O�����'bl`�����/RU���Z��8�O2l���'la{�j�	6Qޝ7�B+�
แA�9�y"������"���T5yq��%{�TdGz�O�'�Ru2��� Yyp1�UgJ�]�f1�F��@!$���'.�'��m�YsB�'��	v��\���+	������M44𣲁�u��U3�KAH� ���F-��i���L46m�@*;�Ҩ��MּbC��L�?2HA���Ò��O�qD�'�f���[��-�@,
6,�J ��NI�<�¥�4QV>P� �<P�����YF�<�v��FrpY� HJ�@Z�h(UP@?it�i��'�Z!�4�h��$�O�'F�*(9��X'N� ��H^S*�c�[-a���' 2D
"pJ�m�T/m�°���ĘnC����tL��q���,2Z�F�(��#=�6�O#&���Ч^�8��1
@���u�釘~��`$�[z�+!��*m:HqNL���'�8"��u�Q>����M���Jdzl��&'D�u�D�F9a�w��)/ P�kA%�OB��O��d�	K� �Qg�ǵ17�����O$�A�j���u���T�O�F����'�b�i�����"�1��u*Y�?����`,\.}@��Y�!L�xu���Q�:��1�O�1�k�A�4��N� ������V�i@�a��J�@
�Ō30��،v1���~��E�X9�� �H#dU!&�  l�*e�4�W�)��1 �˩��1���Q�3- �ꅢ>D����� KIjĘF)
"J�d��$=�P����S���D�-B�p��ϱ;������?��q�^�dc���?���?���4���Oǀܝ~�
y�P��12�8�sa��#��$�L���XG����<)$!
2�j��Cb�6�ӵ��fwj!#�
�`u��k��o�P1�O�"< �p`��c"��.G�L��P},�?	�'LhSE%���|y���).̋	�'�hQ
f{���*�"�J�ai�Z����|��͖G�*�D�� *z��RG�1z������L%�'X��'�n����'K�3�(�c�V^@&��f�^aJ�U�I&��)�%U�	~�Ă%h�x�?9T��Tf��"����,�É��\��PK�5S���"��!���0�4flj�u�bܓ5�Ҙ�I",��]P/zUhBKV�(�n�#"Oءr5/�!�\}`t�T�����"O\�` �U���91!����C7�ONPmZ]�<w���ڴ�?a�����¿R5d|��&ē,a�@���ȫv�(`����	���R�	�6�.諶�����S�į���cR_|����Iâ#�Bpڲ�;�HOVU�r�4.'D���܊zl���`�s݅3��[�Z�R��2��+Z������X%�K+�ɏ}���W�O ��C�Z�h�����iE,
V���
�'�����T5��*�Zl�+���{��i1V����V�
,|;���\ƈ���i���'A�K������m�!h"\���l]��oU}� ����.2���#�;��u���E�)�v��s"�H ��3A��=r(��̦p�^>A��� >U ����Bͺ3��],���k�>2����N���� Rl^�"������?��|���i���wcB- �����;P�>�#�'?�*���d!`��p�)K��)��D�o���4�iZ,���N�79�Pڳ�ؓT��C���O�D�N�Bi�O8�D�O��d�ӺC����P !��q���_�@TD}��KX	.d̔c��i�$�p'CPU�\�'�(O:�@"ǌ���[ah��"SBt��םL��`���8,�p$��\��צEZ�nI�s��U���P��H�J���șj�*@�'c�DZ��oE�z���HJ2���e�����H���y"f\7��t���RV$��J҉�! b8�Dz�Oi�'a�Yҏ�?2�|Acm�(��<���&P�8��'��'0�V2���'��)=f�`}!�n)�U蜬a�	�2a�K��	���2A�qU`2�n��
�B׌<��&I�%��5h��L��t� s�-Y�T�X�nR��M[BQ� J�=��(Yџ���φ���[𧊇q���u�K"0w!�$O�(���#fJ*7�l��i�E�!�D۾2�r9f�=s� �c(�Ud�dΦ�$����DR��M����?1��� `���B�1K�T1�K�%q~��(0��,��4��ן��	!������(x:`�P M��AX���O4��^�v����,52�ŏ6ғ]��i��4]�d��1�*w��r\ws|��d��o�-1��Q�ƲP֍�,u2�b�{��:�?��S�Yj`AJ5��E��u�"h�6"m8C��<s����L�dQ��k��ɶ= ��DF\��7"�nA�DN	`�F�zp�ҚS��Ě2vo��(�	c��-���'����^6��9"�	VO��{�-N�:�����Ta�@�!�\����M�T���\رg_�2~a����'�%�i|(\J��˧fp)[fI*9�\����q���Eu����7ꋺ x����ڥ[����Nצaq$�O�Q'�"~n�7�!�����0K�@���	�' 쁳B��l�R/�6��4z��\���t�i�ɑ��\��d2��݉��	����Oz�R�!o� �O ���O �$�ɺ���n��O��0AdJ<��"DߙW��M�tKv�|d��E�.,��(O:�2�Cã+ƦF�1ͪ�*����cT�<��״	>�#�	��d��Ħ�����&�F���S�ʜY��3jQ�1����'Q�̂���z�늩<!*�1fC��&� ��y�-�P,�ad��	�*$��Oӭn�L�Fz�O��'�ޝxu�H�t����� �BK���3�O(`��(cW�'|r�'�ҧV�t�b�'w�I�3Vji)�lUn�������jK�uȅ
�1v���U&k}���%�^�''"8�@�$V�Խ���Х~��(9��3AUh
�������M�q��9;W�Ϳp<<�Ӛ|"EͿ�?��J�MbF�g��Q�P�s��K!
C䉜C���O���RI4��`����/�?|���Ir��U�VLF�Y@��� ��֜|b�D9d��?9����E�EY��!��ςLDZ���_M�V���ߟ��ɿ> ��g�	�p�h4 ���{%�Y���_�y�P�ыز\�b �S��9Th��$,ʓ
+$����:u���Pa�'X���A"�,�굣RޟF�����`-$Tc3�A16Q��%�M���i��Y?��D�%=5�q��I�6n�4����8�?1����'"���8EN�Z")؏6��(��� I��(�c�;�<5!2��SH���7�v����ii��'�S�+����	Ο�l*f�:}#���$�H�c5�
i�0��K�,0���1��Яdi�y��-�Z��}�nJ����5FD��.�8�/��;��j���5�M%�>`���s�;e�P��UƼD3�K��3�s��1㍛M
��q��R�X_mq��zӲa���'r��O?7�Sj�1R���H��	yV@�k&!���%�HaҔ�O�cr{vF�mQ��@��4��7M�1��Q��� ���s7��5^t��̟\*! ��\���|��៘{_w���d� ��Z�kS��V�@1���<x^�ѐ�@%Q��iɓ��(��ӟKf�-k��|B�6\r(8"�K[p�t ��&QX�b���bҐ`Y��>֠Pȩ�����#1��+4��f엡��u��K6|��'��@�dY�z2ES�1�P���4~�؜	@�@��Py�K�)c�>tJ��һ�%��Y;vEZ"=ͧ��]5��#5�T�x�<����Ĺ$��q��ȆTT� ���?)��?��IV��?����dŝ����d�W�_<��h̔o���ـ���L5�f�̫�"��E��7-���R���#xP��Ҭ7(U���,\��Qq��H��q�3�^^�'�x�[��KTX�(�������QBשr�|aU/=D�ԸC�͡|�h�����`dQ��/D���"W�+F:��hО Pd�P'����ݴ��)��𰅻iU��'��S�J��)rmS(6�"��!�?δ�7�S�?1��?!aA�N��uxC��3
�"���z��S�8�1�rƐ�I���S�%<̞"=Y"Q�?�F�8"ω=`.����Gv"y� ��Pۂ4;�זy�&)x��L�鑞�hGk�O6"}�T�۸XP:�:��E+8`��(@�My�<A@��3:���*��Ĩ�3֨@]8���K��q爓�r�c%H�4$ݬ���e����,���M���?I-����D��O���q��-�rOC�I\���H�~��p%�& ��\�7#X�8�<)x�ilJ��S?�'?m�1)<(@'gǐ�؁�׊E,8mZ�?� x�D_#C�ͱ�JM�!���&9OV�q��R�oo�sӠ���-��C��2�-׵<�́�i���A֛�oj���$'�	�����b�z�!cLV�P�D���4��𙳤֟p��P��HO���2��6~Xy���%�l�剤�M� �im1��7�f�!`��Yk�r�� zv��A6� ���U� ��ݩ���O��T	�5z�A�7��1%�|I�y2�)�隴K]��"@o�	��]�@U�
��u�$�J��h��$��}����a�@�@C/�!�d���m0' ��%��0GL���!�A���cÇ0|�L�c�b�	G�!�$�;����ԅ"�@Љ  S(n!�� z���[#��=��R�!��xZE"OR!�7�h��GC�M�Jy�S"O��)e�K�Pq��C�3-�x�!"O~��I�^����O��pq�"OQ[�P>T�z��5A�� ��R�"O2y��$ X�&�>1uZ\�1"O���g�͢�,�/]���S"O,Ȱ�� �f=���-9Ea��"O<,AU�C��K�ǎl���C�"O�(�
ފČ�b�Q'C/��"O���FlT�B���0��\���"Ot� �v־��D�tv=�0"O�ɑU��-M��HQ!Dղa(.�Yd"O*�y�Z�K���Qbe
�;�F�#�"Onhr�aA�>�T�C��+R��<i�"O|��C�'{��)&�A�s `�5"On ��˰<T>�0-Ɏ�ei"O�أbF�(r�Fy��,˨0�Р�"O�Y��޻|7�0�#
���w"OJ�1�ȞE3����*Պ���"Ob��)��6�T19��P�~�@�"O>XRQ�K7Ad�غ��(8�8)�"OH(i�� Fy�1BB���y��"O>�デ��
�:y�F�G Got颰"O=��i�^X݀PjU�[F���7"O^i�#֦ ��@+SI
����D"O�dy��[�b~�`�2gޤ5E�IJ�'|��	�nŔ!�rA��-m���'Eh�y���Uk��s��FN&��'N���G�J[�XtY2�-�0͂�'	5r��(un`� q���)�'$�懘�a�� �L�B��+�y���%*���~ҙ3��y2�O���{DoOl��Zĉ]��y���VU�����.`0��2^'�y��_ƪ���叫X�� Ye`�%�yBe�/L����A�F"��ˀ��y�E��^dƹS�o2Ij)y��*�yrE��$%Bc�`ƣ;��1��y��_:x�
t��4�Y�u	��y��ǡ�<Q�9S�Fm�t��y2��%�8�F��@���ZC$[4�y�GVs0��玘�B_PԹb��(���ԋG���+�g�� ��kR�P�J��f�z���sV�Mm�n�Vԟ;����ȓP<��7k܋!h�c�K�y��	�<����i�O��YE�M�3�bM��քR�!��M^�zt���X��`x`G� 6eI��牤]q���]>xY��E(��B�ɒ&}��ȍ,*�v5�A�	1(�B�+V�qa��$D^���Ɖ/(�C�I�@_R���❒e� ���;Z8�B�I0
�((4�ީ:P�0�퇑d5�B�	��J�3��3[p�۠��!�lB��4+�.	Dl��{0����@�7�PB�ɑiE^�b�G\�Y���
� ߞ�"B�d	d|�mD�E[`���>�,B䉥W�b(��#��P#h�3 ؚ	pB��9%@B0
@	&}&A�o I/"B�I7Fp�%"1�@'y�<���K�0".B�I�i�$`�[?$^��i�3z6B�I�L��dq��P����s��8�$C�1$�"��v��p�����A����=�I7(�*)�ĭU�}�~MR!@� �<B�)� �Qç�N����b)��UEx�0g"OJ�Ҥ�S�%�����fI�7<K"O��b�-�m1Eϋ�s$d��5"O��rwL�6h�$��ðezl	�"O��k�`�)&ж��4d4�AD"O�-hu��n�J5�U��U?��6"O )f.P�b����MÆ�"O��I�F�$إ�G='���F
��y�ʔ���QЧ
R�Z�*�'�y�P�6!��l�N��m�7��y�D�'K�z=���֍0���f��6�yR-�<=��IP�-1~_�ݳf� ��y��0a�\Bŉ�nՀ��f/�y� Y�u�@r!�Kb0���J���y�@ĺ~P|Xʉ�dFt4��o܎�y�̆�)Qe֬@_���ړMU��yr�ɤ(���2# ؒd�|iȗ�S?�yr	�(�(����	�N�j��'�y�)xe�I���C4<BR��O+�y2�Y7cͲ)�"�x�Hţ鈋��'�,I*��H�O.�`r�;2� {��D8O��%��'�&1���Y~n��O	�� �d��M>��O�,���Y��;�8gx�V	Y�g@lh*g�3D��YT&_�B`;�F �w,Xb���Da��P��7j�|����t���H�0�������<	�"�68���d��y���M@( �p��2vat�5��y��)XaF�eN�}9�a�����|:�}��ȝ?z\��F$�'k�P��b״/I�YӲ�_�G�����hʦ�'��Q\�L��A"T��\�v�˽tDPx��O�Be�;�3}�'��\Y��'Ƶ<�f��H+��?q�B�.e����|�de�u�X!�cҷ53���KI�NT&��퉅(t�{F��y�h��eK�h��>�g�;d��ݠW��Z���6���u����KCfx���ݲ��5�eF�5�y]3)�0\8%�ʐz���s�,$�~�B�T_�؃4�)`�4%Y���d�>�D�Є9��LD`K�N`)��'D�l�^H@�D�՘b�������M�ŎKwZ�1Q�ȫ>����0�t����~��]��/7I�8�Ո�nr�~2O�����Y{jc�Ҍ8�.P�D�� r葫�' �4U*��$�H�	@Jf��9�R�[�zqQ�p����DtxFm��)V�a�O�������-qT:��-!��Q�'0�<��-��.Iڦ)F�&r^t��O�i�@	�O�=���C��蟎$��T(UvQIl[8I0�<@�"O4��է�:R�@����4>�a"`"Op�``�Ym"��%��>���HQ"Oةa��>Z�&<+'��b�t�g"O�A�b6����<�xIp"OB���Pg�*�H��� zT�z�"O>D�q=*1��q�2hH�ʥ"O����C T�9�e�+�8E˱"OΨ��ǒ#�� ����u����U"O�%���M$QЭH��Fx�a'�'��(� n��� ���6*v�yˁ�{ֺ-h-�Ob\{�"W��	kX���6E9+J�(���%
"��C�-.qj�ɡ�J&sT���C�JL3�f�����ΧU��a�手03�´�0銱Jy!�?Ŕ�bD�)�,}���X�~����̉:"B��b꒷=ʄ��w([>Ɛ���i��Op�E��C>2�j��I���z�ɖ!5D�t�U%T$g]R؉����x^�b7�6_PJUb�+m�]��/w':u�uE�$eXX̡��F�I�8�A煛U����J:��z�"<�:��0aN"T.m҄���ep�P�F<C�4���ׅL�2 �&qb��c�+\Ox,ӄ-�x�� �Lȩ^ N���dH)_D�9"��0Iм4�ר	1#˖�����$lr<ÔM��CY�����0Ƀ�1}�s
�'�Nh�5��`�(M�?\���
��^I�A&lR5�@�O��ZL�U$���i_�5<��X��ȸ�� �8f^�A"g��I��D�;}pF1�c�Ɨm��`ړO=����gՁ=ujH��KM�9�P��I �|uJ-��h��b�� �1k�c�;1PZ�F��͈��c�'J��P �QU�C+N�i�J�Pm̓Y`*�`�S��R�
�7����f����UH�i��3K$0���6qN ��h2��4t@ �P�3T�ܭa�Ⓛ�>�G�6%k\3.%$�hҩZ&e:Vջ�цZդB�I(��,�p�ߑ}�&�-Q{��p!%�}v�l��I�j��܃#G�
^h�ק	��哞-!VT�;e��hUe�*�(@�#�%�X��Ɠ �� ک+���E!�� �Q`���­L#vV�Q)��1��F�-��<�=�4�N0H�
�K`c��7����'Jux��S ��3��=���7M*�{�)Z�\(�d��NޞC�z\��,��-��I�
���ď'\O�A2I��Nԁz筂������|��B���[D �!��C��ݨu� ����I�#N��;
�~�K�&�=JĞ�B`W9Fb$��ȓ���
6���>ٸ���H\�H��mȠj^�e9�L��M))����������N~��
�Ǽ�F��^����``,��ǒj�<�%΅v�z�3ABʁ
��̓�	�	^�\�Qw>,�<���̽8������t�t�o�Vܓd[ �CJ��)��	�Ƀ�B�j,��ɥz�m� N,��y!�C�EĞ�XA@� ����ϯA��n��*���'�ў��p�'~y� �X?.eЄ	�%��ɸ'iƈ��m��F+��w�ı�Ph�$"��pPyqq�gN�u���IF8��HP�K,2,�)�OdL\�*���
V���Z�@�&����>�	�/O�}�%� �k$a��N��v��{�4�Pxbmٜs0��Xv�F5'ר�x��^-�y#�d�lXkR�
M���'��KAA�����`AK�-i�
	j-R�L�Ō8å�'h���K��͔W��0s���5�S�ӛh�ER�" ���?N��B��3&���!$:aԀ��S�%��"=��$�8�0�kv��[q�סf�,��ȓ@1F�
��X_\��ף ��N����B�a���d����ʟ,s�e��o4�D���7(Z�
7 I�ȓ]�x@@���~�q���(Ui�Ԇ�:^��X���	*���k�������T�@.�I�r���ǖ<J��ɇ�J��)�äZ�r�^�`	qP\���mߒ:M�F{*�����2��i+���EY�s��(�� �gl@�c�'�������1�h��� T�@
�'�J�[#
�6<]k�KȰI��)�	�'IHr$��;4�|Ycda�!D�6�J	�'^���f��|N�����Q�F�<��'�.��g 3x `��N̽e/.Ł�'m6�Q��m�h���iB�R��j�'=lz���8C��f��W�h�'F}җ���
(��i��z�<9��P�0�+#5�IP��Nr�<�ƣA�`}A�*XC��m�<����:lRb�A+�ћ�iVa�<�̅�������S��3��c�<i6B�#T���E���`�
]�<q��P�:����K#���S��^�<yCK�:Z�@k�ND�xєYӔ%)D�����ʻb8"���L W�v����'D���F�e��HY'�4 E��Q�c"D�(+2�%nMJ	�.�)�|���%D���B M<-
�h�gIۃ[g4Cu+#D���b��~e����%ם#p��y�!D�P��S�h�"��0dA"V"2YBu� D��C2C=<��	��뛐a���O>D�$��,^�kp}�v��<��U���?D��37�+'��R�o^0�QHp�:D�`h�Hς.?�m �M�5~����;D�8#F�H{5h�CP�$�����*D��0�C���Do�hh-��&D�ؘ��M�p3�Fe�ޔ���F"D��C�"2���vZ�(�f#D�@�eԨ-j��#$�W�\�[� �7_�^��Rf^rx�� r��3h�=ob�
��6�����"OPzf$֌S����"J����""Ov���h���x�@@$��PCG"O�[5M˺ /���p���r��"Oxy���۠L�r�I ��.'�|�2�"O�=3���>Gp�X�2�t�(�"Of]W�(de��a��t٦y�t"O�����/-����IM�نl�"O��i ��<<��b��BJ���"Ỏk5�� >��+�i������"OT��!�		t�Iq��[��[1"O���2HՕ�Uk�f�\x���p"O����� Z��xW�
�d��"O�P�s@��\p�dk@E٧$�ʡ��"O<��Rk[�"<^-؅$@/Sب�`"O x�@�Xz8���;&���C"OF]�g⊄Jy�1���E�lwQ0"O��Th6$s$��I:��"O*XH�O�#]~,A�&�_�&�����"O��H��AVܵ�2Hw�lv"O�A�	+K�.��3Aѓ>�0 E"O��[��P8�n��@�%����"O�����:*1��E�K��k�"O�Ex�e��Yl\ ��.��d��;�"O�9Ҡ�1�4���wA��"G��B��n��!�E�{���ё�#�FB��7A�(t@�/���+
37�B䉠#�^)��Ȇ�R��=��-,\ B��=��T�~��0 ��66G�C䉮/�da8��В#P !Ja��	�(C�I�,~�X3��J)>�ecƌ��FC�I�[�|����������;J�B�I�u��I��,F?e�"4��dX�i�(C䉗��<	�ɛI�,P��#$C�	>lv@��e�6xIZ�Rч�5�X#>����^2���'Y���N�y� V!>�@dze��i� xe�Ĺ���)" �J���$+y,�5J�QtX�b!#ªN�D�liA��0�ƀ�S�O�ⱐ�J��qt� �M¹=|Vj�c$HCo.pZ$����8!!7嗯[n�c`�H����'?|�p7�#3��AH`�O���N~��F4��M� OO��:��!/<�q��o��p�B�0�� �B�����I�Qe��'?$����nz�xu��_Ֆ�{�KB1�u�(�����n��ٛ���K����󄝯Pˈ���,��]� �C��i�1O���#W�4�k��ǻZ���C��M�4d䁣�M�?��p�AN�U��'ڄ(3D�S�fűG�ƙW�� �E��:Tk�(@<;Tl���ɬ5��%Yub�!��
�	2y���X7�L���9v��0!��r��:��![�Lm���H�b�	�'} !�M�3�$m�E�ֿ2@d���/<O\1��%��"f��#%!Y9tl������<6 [�i����=��& k>ZJR�2h��4��,�r��B
�L6H�롘|B�/�H��@Q(	����F%G�'�N}� +H$��a	q�ԱTz�5r�}r$�>-ܬ8���`��Y!�-�9�ē'��� �+��Q��0��C!\��{ Y+B?���q,>�?v4�Tp��
:n���+�oד$Լ����|�gǳdT�ل�_$hm����e+eF�Y�aF~"I#�'�D*W(K
s�m�'U�X,����'��*����b�B���E rJ�1�xM�v�I!	gR��SŔ@}��i>9+ �\�P���
B6��0Ԉ��	N1���K>��^>qi���P $Sx8�K�hܓTk���CN��Ȣ�Q.u�"�'���I�jXD��b]�Y�~�c�AO>SٔO��S")^2]�	c3*�f��4����e�$1�-�v#j����<)P \.��Q�DCGWD �"ʒB���P���	���rpM�oB�x�K\	q�VYٳ�T�8YT@ǥ8�1O(yX�@���E��ح}� �I��A�WVŢ�!����$Y�F5^|Z�
�p�؍=��-�FL�b�q�q�
(,{u�Oz�ɁR��a4��;�����q~�32KH�Y�����_�_8��N>��O������c3�5��%mܓo4&��b۞:Yに�G>u��c�)ְ��O
moڇWxm3�i��Bd�N�)� ��v@[>u��h1�J��Upp���(���Q��6cЪ�C�{�O�3l��ı���s��!wG��r0ƨ.��9(�@^�^ps���M��G��x��@��$�Y�}��ᑎ��<1O̡���\����S~��LZ>��uc�+� v�"aI�[�J�x҅M�,��艀- .kLJ$wFr�bQD͸Xkh�Bi�����'���;}�[>�֍�:w�6-���X.1�,�p��b�ᙦ�5\�bN>���E��`kߒN�P	)��~�`�Hx�y6�	rE�L�>��'o��'Z�a��)>��̂���[���N<�M��-���@%�-;"�$H��Q�K�j_.NԢݰ'*=�����T�j�f�0��O�w�f�����X�N��d�,���y�d�J.��	�\� 0�"� �)�.3�e�H\��G~�O�=�'��)���Y���S1��1��Þ��I��ɗ��5!�ȪO��p��U�q+�ǊR�(}��c���Z�	�Q����>Z1h�'����~.��Q
_�{��(2�A�B�t��*�OB�p��^�*i����b������ ��Nɐ0kT�C¹X��O��$�O�q,���&j� \�(f�
��Ҧ��@�C�9�h����#��q$eJ�O�:u(�˟�>�?Y�'�5lY�%��
�FB���	�C�4X��ڪ`�j#0+O@�p%��'@�h������B�a��+���'L��ƣe��l��#>F���ݾD�h=��	n����G�.4{���%2
9�`�;��Z�I(��m3�\���?�d^?-�,�K��YR�a�4HA��f 
!��*. =k��|"��
F� <i��P�d�e(�`�и'^���&A+�\)贈�]r:}`�'�X�DQǦA�!��'fހ��"�i�&�����'}e�G��-g��xb��Y�P������@�<��p��vK��F�r��c��^1?��T�G]=qJ耱�B.�M1�聳Ǔ:����3	G�=�����肞 ;���'.!	��N�[Y�}�׌�
��)��"Ond��eO*�*u�C�x�!1KL���j'D�=��R�	L�Ұ=��ON 
>�KTb�Hh�Bo�U8��
��G��TЁ�|��W�AxU҅���`t�S�KK���'����N-{���B�'ӫ	7�}��}�bҭ?���t"�{5��8&������Ѩ��2/��B�*�X���Z�>!�&�����<+}&Jf�_�c�R�ğCuɱ�o��$���:'��j�����	&&1F��ĩH=;!t\�[+
lC䉄X��#I��16�@�� 5'LH�Ɠ����A�dȕQ�"�&
ht*4�>)��UN���H~�=1�S�(��ƐT�t@26�l̓tA02�`>��%�۫�j�<y)�=E�J�#��B*��|��dܓ������(�Rb]�RX&�<"QN�}��	+��C�:��ňg��R���g��R�>����'|.,20�Ɔd�:�:��W0X���*���C�jmJ�C��~�*O�j�B�?��y�C-�.7��p"3D���H\���'aɀC<]"ݤ0`ay�F��e�h�p���5�@��tb�y��	�E��% �����9 ��P�L5i�ɹ���7B��PZ!3�]u���D�|��E&����@�2_hGaU���'8�1��4�2Ṙl�D�Q�}b��T�"� X&�,m���X��[�l%�03�-�ᄄ3'	�����\ٲ1�	�2�����i�DM���V�Y��p�E�>r ��C�$(��Թ$�T��㉳r(�U"��Y׬13�f&UgD�ȓG���{��ԤB����J'� p{��'
"�K�����ĵ���1@"F�l�A
(s#l�I(Al}b�P.H@�e�\ �b���'�bu[�� ��А�#��xD�Ak�E]�8��@i�M�5lޡ�D-)��L��
�V��J�(�1���`p�m
C���P�C�<��������~�⌀�LRd�j��wbU59�X�S%�(XK$tCR�����O�Q�;�>�'�>�6��r&V	�OZl ��\:D,��Ԃ-�\l��K�Ī���]OI`#?Q�jӔ@�J�"R�ȼ|m�˧J�D2 ��EE����'�vGN٨��'$rn��x��;a�ƒEh���:o�]�ň�
%���f�j}����T)��.�CP4���'���y�MG��`I�̦6zu��Q�Ɇ?�	xq���WYt�e"����ɛ�牆t�$x{��".DT���S$��hJD�W?q%�}�ɫ4���~jeǃ�;;L1"@�WD PP摓�<9��k���pzA�������ѭ�M3&H�<y�<���Ӡ.����a�1�����"Ƒ>��kF)r��|)	�5�8q�1��h���A�sy"�3�'s^|���=�^��'�f�z�:l�t��L~�T�\ ;[f�P���d��Rb
	����D*�ۇB�	 �P���8�:���&W�l`:5��74��w9�ab˙a ��5�|ꃕ|/M��͚ů�\]���</��h1M>	���o�i3�k��|�X����X?a�I���ek;`����
!d��7�
9,�� ���P?	%�\]�	� ���~:�g��!��`�nԝ=�d5Kv�V�s��hv�[`F���G����5@Ӡ+����Oj�{�? �q�C�	?��h��`�����x�(�1.A�HǓ�����≅��������i+2��'nX�Bh�xܞ��'�p�zf��qpbpx�f�j�bV<:Y2[�,�5�jd*��R�f��d��XW|=�����H�Xz���A�
�>�6h�Ӫ�r�	�OX��ML]��˒�U ���ߨ��g�hk6�Z(����O�/#��
��.�D�cC����&s�4���Op��14@�0nh0�~��*DFA$��\���]�=׼ ��k�M?����N�Ir�*!�~�r���,�=i  Q�3Q�~"�dސqMr�ӗ0��1�1	f� ���� Ӽ�g�ܛ���%�ºB��|�pLFX�DX�5�����(O�Řu���.q�u�'|��[��N�y�P�+��'zW,q���s�"~� &���&���ĩ����

�HUd�'�Y��Z��(�!Q�Ʈ�a �֤B���y��Ղ�~j�"��L+v�G�w+�-I�_�&k9'��Y�,Ο"��p�H�)�hhP����{4�܊kx �N>y0�̪+���&�ș�C�
�'SJ���k�|�iS�ƉE:1C3%�xz0��U͞8+�J<�1��1�V92��X&�E�Gf�I��ji��J [�LYV)�
�@�����n+�дM۴U���L�{�h��Rm����"�����m�8�&MY n�4�DF�N����C�(R���G����d��''X�i���;g�T��C۲X`P�{p���F�޽rL�!)}�-�-�g~B��?v���01���X���q�J�t����Ԩ
b @f�יj9v��6ZTE�gnʃsg����0{�$E��E]�X�&<9u��/����L:�N:���DJ$��D��N��4&�a��ҷK((�)q�_����(�+u�O�ulT�Jg�]0v{�|����r|�X�B��T�9�k�:Y�<5-P�$�uF�b�� �:5Ɯ�;�c�.<4{t�0��?�`#H�#"q`�jև��q��� v$= ��&=�ё�g	�	c%T��O�̨3�f�6E��-YW��%0٠��RƜ#�lQ� ̲5�*] �*,OT�#���abHؕW@��B�+2�Z�$��}��[��~�%��I��uid�I�YXB�cCː=v�a}�;l��6��#�Req��:���{f�@�_�x ;�%�O���'Bʜ'
�����)�'=-�@Dj�\�����'�T�G{BG_�@�S�
W+�l&>Q�8p�P�D��Cʡr� I1e~���'�mV�+G��ϸ'ab!�S�0%���sE
���%���jQV �$�PK����"|�."S������'�<�u�F�B���2M=�<lr&1�O�s�JN�Qwvy�W"$X�f��l�<��N�D`����|�m�}�Y���L4� NQ�ҥ�J�!��G�U�0�y�
��2��#D��!�M��9Pe�5d�J�"��L�>�!�\/1�$��'��?3lr��	&d!����t���Z^H�x�Hݘ|�!�dػ)�*TJ�MN
QKHm#�"ÿ!�V>Ŷd3�앳S�b,�S���!���9�1�nͭtx�	�˙O�!�d �oؠ|���EF�6*7O�!�d?<K�9Q���T/���J�,�!�$��D�D`!2�D�P��<U�!�D�8+n�(cn#4��@�s��!��GdqȈk`�/��ɠ&�E@!򤆘&�K��:�m�嗓+ȴ|�	�'֊  C��/�j ��Z4J�[�'Q>�����GsHe�7�ӃV���H�'E� �����g^�,�gh��I��'Y�;SL��z�['�E�$TH�'�&p��EP02�+��]p� �*Op�U#M42�^���l��
8u�"O$J�.�rOf0;G�U�D V	�#"O�+&]+J�t�ݽa����"O �A`ȍ>8�$hlR9��""O����շ9��ys� �2�DY�"O2��r�
�$S�CUK�&$����!"O�Y�#�Fr�0@�TJ"X�"O����i�+ƺ0
Fk�!���"O�;!nK�v&�����
L�Ɯ��"OV�q��^�}� �k�g�h��"O�9{'�	�>bJ���܆6y�4#"O !�+�Z�pB �Q�>F ��"O���f��(¸�/�0z.���"O���FB*j��x�/ڕ����"O~�9��Eˈ�q�΍�q*ʝ&"O� ��Qm���	��ӳp��"O�1qDȞ�Ȁ�*��U���"O�M��
�2,�z��JY�"8��X&"O�|C�.�.�2-�'Ǘ��đ"OBy �N��dPW ��{��\��"O��X��[ŨE��a�<>�x�U"O>�1� �?L~Uh%`R�]�\�u"OPa0AJ	+n`,KtMӞL��4`b"O\)�c]��\k�,ћRkb�8�"Ov(�3�A�3yd@��qU����"O��"�!{�p22l�+e��(��"O�Ԣ�,^
�j�*a+]�t�py�"O�IQ�_�z�l��0!��'h>4Q�"O$��FP?U����fàFJ�T �"O�p��N
+h}S�c�'T>�"O����f��6����b�	b�\"OBM!&�W7"�A�gQtR�d�"O�� %a�T����CD��C^�D0�"O��s��`=�D�LP��"OH����5F��⩙�D��۳"O�A;����P��0��H��4.�d�D"O���!Jtr��v�1)Xm�"O2��ɛiIf����	(Ib5"OT���P L��k����G��{ "Or��4�]7$�zh���׫S�P��"O��k��ؚ%�����CK�K�P��1"O��	��k����9�P"On%QS�ي�49cL�t丝`1"O885+��Ν1��1���D"Od!�ƭ݂0�Uk��	�v���"Op�Qd�#C	���C&����<�"O$�b�L�&\��%@8W���3�"ON�&�O	rǀA d�M�y�"Oj���!^��lA #��W��(�E"O��j�+�r��	�`��B��H�"O�rc�*6�bə�� ?"2lP"OH�b�D�$,��gk�;2;�`��"O���i6[�Ni�����0uɳ"OB���"H���X2�-����U"ON%��G��1k&}ؒƑa����"O�	���\�1����Z�~�1�"O���3d��LMr���ґ�l�w"O~�v�ԒI�T���>bA˕"O(�رa�p:�9�#ISHU�h��"On�����r��M0rʑMN�!�@"O��+B@΋:K����(�NQ��y�"Oց��v�҅���N9I&8*�"Of��Bטd�R8��ֵ`��"O��r#�
�9ԫ͢
��%"OX�{q�O�	SPh�ǈ�r�|19%"O\$QU�X�]��P�1F�4M����"O*ABo�	̵�r'��R5�Y "O&A"�ǒ��	��5ց�d"O��
V�SO�0Za�D%(�T�U"O
��tL�(P,�� �A�Pd(�"Oj�j#��VB�U�� /��|��"OL��D�Bf� ��B�T���"O�%���~(�\���mQ.=h�"O���`ԩ9{�x#!K�/Q�ԣ "OH�ccPL�x�AJ$vW���#"Ov���7�tI��i0k��aW"O���U0��$h��xT��"O��` ���3f��դW�<TQ�%"O�]���S��ePS�2I2�f"O� ��+�
�?X��uX��L$)-@�;"O��I�&�E��h���\	�8�6"O���7Ǟ�4�	$B0?�ԍ��"OT�x�ÿ�	ʇa�sHR�XW"ONX�'X1ߥh� ��$qQ�8�y��)7Z�����LYA@��y®^�J���3.[,s�D��B��y�P�~I@3KV�uR	Hբ ��y�íI�����H�DsШ�I��y��L<�,�ŝD� ����.�ybg��Gut�b憖�d���Xf����yjJ+ d�D��	k�mb�%�"�yR�yR��E�c����!ޝ�yb��+�V#�!�(H�f�+�M	��y�HU�"�jeZ��,`F�ȗ����y�gD��r�Jdg�u��`	��ӏ�yrCΞ ��%M�p"	��X!�y�����*����>m6
�9�'��y��[�uB�%QS�۴-l*\gjܚ�y �gC��"�
���������y���>��(��\4�|�2� �yr��6#�	;@����DiZ�k���y2C�`:���q�p�2m��yR*A^��҆�=aȼ�X����yb�\�w�0��*��V�hh0��3�yR�׺~�"^�z�d�2�d@�y��5���b� �[�l�C����y����#�m`�g �YPL��CK
�y�eݖ;_x<�gܶg��B�yr�Q%n��I0$�/I��;�̃��ybO_3_2�I�Z�>��!qA�0�y�f_�<��7J��4��IǣK��y�L\����e�Uw�����y��gO �L�Uͼ���2�y�DC�Xo"@��M7��-qK��y�Y�3��A�'�������y*rU��p�5���Y��yB�ٍJX s�E�)mz������yrDF7���F�[2z�����M��y�R�a(R @uG�vx�b���;�y"��a��@X��Z�G���y�5)�AJ�G��~������	��y�c�!���Ձ�5B2QF�ù�y�bW�R��Q�BE�6x��j��y�憲St�x���C�h��M��y��4W���; �\�)ٌ��wI�5�y��A�q�H��,�� ���ЂC��y�B1rF@� C�j\��I>�y���b�J!PQ�̋e5@u`�����y��d�h�m"4��̱`P��y�J��bk����P&��x�"�Ժ�y��^�H7��ՠ�+��`��6�yBˢ*�~e��	�.�4�U7�y2mD�epJ�"t�%\P���yR(��E��$�0K��	PP�34�*�y2@LD�M����}T��@���yr�\*�vؘ��B�>T�XS�E�y�C�+/B]���>������yB��Wi4���=	,��Ɂ��y�ŷ0Y��W�ѫJ�$l �y���AȠU*u�A�x� q`
:�yRd�=X�f��R�:|���E�y�S�\^��b�0?����BC��y�b��pp����,`� k����y
� ��p�f�&1�(4Cs�16�6x�"O$���ڙ`��8�!��x���"O\�6�[
B�ڜ��
�:�P%B�"O��Ҷi��1p�P3O�$]����"O�X���R�rs�4�¬4,����"Oe��kE�3ƠU�w̃�l���E"O�ep͐�MX<)wbJ"a��j�"O� �ӭͪ
{�вᎶ^�T0��"O���&U�}���R3#�9�	E"O8$[ J2 ���&H/r�@�"O�����י�<���OK�	*�aأ"O^����Â]�yb��#"��"O��P���)�Xxa(�&R�s6�O��=E�������E
L
���_�ҙ��'���*�0�d��#��	Nw� 8�'`zq2D,�s:pu	��@�47�(	�'�T`C��pyq�`L9iJ�z	�'J^�GŌ��*�)�H)]u�Ј�'F&�� oD%R��;g�����'kb���\3 %�H�1OCW�ε3�'�zX 7K��
��U!��ՈO�R% �'�^`{Q��}���3l�p��'��ZUNB�CP�@#k�h�@�R�'��݈�B߸Q�����N��Y�'\�u�E�MU����v���c�'�%j֯����tȗ�_�q�'|<�(#o�3A�%T*J^��I(�'�\�q dW=I�li��Yk���'LN	wo��2
<���E!eoR�J�'��u�g�'3͔e(�h5U#~p+	�'!�h1�l��Q��mS��@D�X�'ܮ���A+
4��L=2Y�aK�'i�q�%$\<�0��,-�R�h
�'L��P!L�7P��c�GS�!]�!��'��k '7��ҥ���H�H���'r<�)c�,a�<����U4\��'�-�rE�+�dxRR�
�R�\h��'�2E
�E�<
.�AĽN�2�Y�'�T�6�\��ց0�n�[`���'�p�߈E�(� H�_��%�F"O��9�e���W�.Z�*Ȑ"O�I��΂u�92���0)�)��"O�*�햇��yb3�6���"OD`{��ǓQ�����ք`���
2"O��XQ��z��(0f ��̼J�"O|X�`L(���A�6��Id"Oi:�ںz��oՑY1r�(�"O:Y��Q',U�����f�v,�"O�EȒ��F)>]i��O�wyr��P"O�AxE�Dt4X��F&d��`"Ox�
r��/3��e�'�O[K:�I�"O2X�D�-�ȅ�226�1P"Ov8���,��A���#F����"O�Y%��� K2Q����>+��2"O�]C�g�m�@���	"`A �"O\�a ��]C����Âp�̸x�"OtE 2�3^H]㴏��վ)9�"O��Q.6h)�I:+ƺI��"O8���6J �)S�y�L�C"O�̘��)�9[�胏@���[�"O����E�p=�Q�'2�t@ "Or%#Ӄ��L@��a��2F�:u"OYY�W>�~@x]I���([�<�g#��X�;�l�,��QU�<� &\�`ဗB2&�r�aܚm�r)R"Op�a0!Q#{��=�����q�"O���#�ɹ8�*��$�Y�a}l��"OT��t�ˣHv �!e4bkVEn"ORp�򍟍~ڸQ�gתoSfP&"O���F�F�B�)�`�+q��8"O�u�
%@��]9s`� :���b"O�8�1�W	s���˷�ϳ��92"O�mK��Jk���K3��q�"O�	�0�+9�>�j����x5�)��"O��Y��!]2h4��oX��Y�"O-�T�����W�#+���"O�e ����I��H�R�^/~�ȁP@"Ob�"���&�JQ��[�j��"�"OX26�P�|bl����:["i%"OF����A �-L)]`t�c"Ot@s曵X�P�t�&j!� "O,�uBY��`;TbČ�P%"Ox�+wd�)Q�R��˞0t�c�"O���@��9F�xBL�u���3"Oԕ+m�)'b���ˋ�8ͣ�"O��
��V@l8�Y��I[�O�`�<I�c,"�"U���Rm>=S�J�b�<A���Q�`�xנ,�D����Wz�<I�+Q�B�|X��gJ$xۃ_r�<�s/��N x�9��#I�X c�FIJ�<�-D�W��¢g��@��:���G�<�CŅ[U�PJ��;!�4
ҹ$C�ɥVc��£Y�(�����$c�C�"3�t�z��NV&\=��2tF�B�ɮLj�`3hV�:^T�qЪ��XC�%z9����ܾ}��9��M&�>B�^����_?І�{��`�vB�ɧrhD\�š_0����H�Q����d9��B�\��<`�ŵc!���I�g�F;#�:���
ݍHS!򤗎�ȕSQ�-1匴�`�M<17!�.�|e���@�O�ƈ�G��)'!򄁸c����	�S'��v�� p!򤏍8���{C��_��\�!�$
�Td-9��S�wxX�c���cw!�D�z��b�aԍKa�Z��`!�Q,Pj�I��cW?_]f���	�2QX!�d��g7(`h��U';�x��'��/Q!��A�����J� )�hN!��+��h��K��a���a@��Xa!򤛺k[��9�f4�H�P��6B�����"y�E[���z<I�i���C�P��z!/�>Ev �G�"�C�I$vC:qK���d6i�EӓϮB�I�gy��8�Dϕ'o�h@�co+�B�ɨ|�xQ�d���/�p=3�雸#u�B�-������*8'�pB�G�
D��C�:t�䨡'[8A�r`��B�L�B�K�e�/�4�`F��j-4C��1nn���7�Bt�c$�=s��B�I=R����+D�"�0⥍��C�I+y�MR�AGV�P$�eH�0.�C��6?��#d��Ra���`�:CÄ�PD{J?-��I�D?̙�3F�!�0��7D�(Q�@X�킥��$EG�uj�4D�t{�O�q���rG� fX���C/D��(�<,������P�r5�-O�=��
B� �t ���;]s�1�gW��hO�π ��v�5�x�Pv���:�����O���D�'	"�Y��D�6�1����0���D{���,9֠@�8�V��%�I<4焄�"O���ч[�\D���]�|ٜ ��"OP]h���	 u��b�к5�H�%"O($8�ir>����-h�ܠ�"OJPc��l1pY�CG"���2G"O��{3�J�H�f	b�@ �J�U"O�LSp�V'���;Zw��"O�):�-��f����dT�z�h�9D"O�i��C���PmH��`~��"O^騵A�$j=z�����*�Mb�"O���� ��C�~\jĄ�H���"O�0��?���{���5u�(p���IJܓ��'yZ	{�n٫%l,+%��r5ڌ�ȓR��2K6�l�DC!s�V1�ȓ>�
.�9%���RgkZ@V����K�P�ׁ6](�ˢ��o?��$���IH��(�e*�<Z�� H�Xl]�P@k$D�Tx���IiDQ�# ?HU
��>D���5"	��su��?'�2yॄ<D��b�(��/)��Z�nӖT���l9D�@��V�Bz3�)`X�ܻ׬2D���->BFf�6.����aԨ�<
�^j�3�� >|#��#.C� �$=�%�'���.}"=N�(l;��5���wcF6�y�j���d�ڛ>V�A�a�%�y�L�,%Ǭ� f!C�?ў�9r���y�\\�-@R�7��Ô�]��y"�pE�FE{�戲1 Ѷ�y�@�;S1�4����(��:q����ybF[5!	vTq��	N�vd� ���y��O�g�z�Ȇ���L�R9��Z��y�*��'�(��� �1úS�����'�a{r����J��ڟvy�H�e�A���'�ў��e#"��Y�6��7������v���Ob��D�	\{F��s�R+ ���$0��Ā5~��pa&֕'�F �a�7����>�C�
���Ƀ"��ݣW��^�<id��?�u[���>>8]*���V�<a�kB�q��y��+� ��QbS�<A�́��ha!רp�RLP�+Fh<��JY�!�dȦ��>%Kh�7�S��M{�'�Υ2����-N����5]�);��y�$�9|{>����1i䔚"΂6�yR@��4Ys&>	���
�;�y�h��r���',^�J�l�6�yBj؂�jh��Ÿ&�f�y�
���D>�S�OvF �"-C�Z;���ʆ5�lҏ��-�S�tDϚ#0�����ȿ.^-������KX�\�r�-~t԰:Ǡ
�{����1e%D�|�X�u<����m̼E��b����	�	=$"�T=��9�g��J�Z
�'/tD����1i�	&dH$q�'�Z\cf��L���b�(�/.�����'g|���Ɗ� 0�AoC�n��A�' Z=��^�+z���_�r�:��'��B�^g�µ��aP!?��M3
�'��L�-,&���:�㟞1ƀp�
�'���¡�L3s�pHJ&��ĩ	�'���e۸c5�@�@
�"��x�'��,iVJ�6��A�q�M4#��)(�'����&dуr�����ѷ&���'� �ɃJZ)t��`�0����#"_�<� �1����50:\�(��A�N���"O1��-��/J�WL	�?�.�Ab"O���Ë�k�\���K�Nж)h׺i)��Tq��W� g�d�����!��6-Y�`0˃�d������\_�8��>٢NѰZ)���!G ?�L�z0��U�<!b�R�qE#]C(|z�b�P}��)ҧ<fX��"���7g[�~-~Ȅȓ;�8beO
n���𸜄ȓcW�i��$Kf���NF�OD$�ȓE+K㍃&�"Y�xa��ȓC��i�5⓹+�llKc��\J|��+�R<IbK�/eF<sV�I�dd(��I�~�ō.�(4���1����a%
�y2�߂R(rE^)���o���OԢ~�C-�
3�4��l�E�F��A�<��#M�bN���ж),���Z�/^j�(�D�O>���I&L��s�*�[5�^)N�{b�d@!*H��,Ab�����1O~��d֠N&�P[D-�!NH{b2sQ�HF{*��5A`k�dM8U���W
Fͱ4"O��BHG;���J���2���"O���ضIԔ���# ��k"O��AT���kj�,�5aR�5��)Ęx��'L��y�91�2�+��)i=�3��?Y�4����T��A�(�TQ̕��Pp^�r4o�1@�؅��Bu�1��g�ڜ���Λ1,�����E�w�䅆�u����f�?;z8Й��J�W����ȓX���BD� Pp�0!��	�i��e��2Q!�x�����(�v��)<b�1��X<?\�p��6�����o������xKJ���Ƌ*ü݆� ��a�T�E |����%.'�ȓ4��e3��&z������L�`���v݈E!���%���h0B�D�����BKRD����蒤��QEM*4�ȓl�BL�� `��v܈LB4��a����e���s L�4.: �2�(D�T�g�� L��h�)̨�@a�d,D��gH��XP��������y���*D�`��91.h����? �h@�e�&D� �"�]��i[׌��IL2�N&D���SÇ�@�� �!��
�n�S�K$D��"�˝�iHp�� ^L��Ю#D�$�(P�7�8�����9K����F%6D�d3��
)��B��
����5D��+7nS+5���k�.S�Nl{`�8D����數8e�}���,�ИbV 5D����!O?az�Pb��F>#μ�`�1D���eS�vN9��#Еb�|ʀ�#D�̂t틝a��XIA��fD���"D�BgcA�XdL�bCT$�V�j��+D� ��F��]�d5{G#
�04���*D�0ٱ�D/ޚeJ���w�L�2�'D���4iעX�%�![�Vkр&D�D�P�GF��"T�����y�L$D�tz�J�L ����I]�HEI� D�ؠ 8Q����C�3y*)Pr�<D�xc��ޙ"���;����[�35�9D�T1EHB5N������d�.#D�\�@��2dRbt�E*o����.D�(��J@�4a@�JW{��x��a.D�,�Qg9`h�A�N�~Ѣ�*D�� ĩ���M�,P�f&!�85i&"Or� /ٓ	�<T�AEZx��|"�"Ol`0��I��z�0%T�<�~��"OB�yg��/[0��B�ǾV���"OY )>4�t�c��\(s���q"O�h%�M5�D��X}�U"O>P(&�͝�,}��!�uK����"O�����T���2V@KJH�!Xd"O��������4���@+Z�C"OQG˟��������" ف�"OН��*�^p��#֠�1k��"O⼃ad��v�h�`�	�O8���"O��Ca�K1k���o[�K?R�SW"O� Y5X�;�p����C?�p��"O�X��#
�G��h�!��v��(�"O�У1KL��r�, ��&\Ye"O�9�%�݂u�<�@F��c�\���"O�-1�i��hR��^>D����"O���a��@�e�NA 2E,���"O�����	CJ�B�d�%Ӻ��"O�)ѩ���Y�1�ݖ�p=�"O��	,Ļ2���D�<�H��"O�I�C��5	t1t!�6�6��"O&�����+,:(:��� Xfvl��"O��I kħ-���� �\�ax�"Ot�+ց���Д��(L4e�T"O,��0��Ny����k�YY1IDf�<iĊ�*7[0X��U��BY�RX�<9e��� H�3ؽ �ZZ�<�����D,X���_Q�N�ad��V�<a�GV�6�xa�L
b����Bn{�<�G���~ ���_�?f�v��B�<��� ]h����V�6���S�ms�<1E�C�D�6$���D�8o6�;1�p�<Ѣ���n`F�>`ܑsr̕a�<I�݁ �\���±�R͘�"�u�<	b�W-4���i|X0�.�p�<IWARxb�P0�Kξr���0��A�<�b!
��x�롤�5S��yxV��~�<	�K�a�Rp��(�+�>���cV{�<I�#ˤE*��`aH�-D �{�k
Q�<1��2ZyrF*�%.�Y�d�Me�<!�23\��'��.�08�0bBz�<�2(:(pU+�B�'w�����j�<�B�7q����!a� l��E��G�~�<�	ٷta ������,���B�|�<���]6(��M�~ȌS���|�<�f�
�)R���@}�Mc�DHP�<�.�&V���9��^T8�J��Fb�<1��ՀnC�� ���,uLxM1mOd�<�U��"{�]B7�0ɪ��7@�f�<1 
�&)�����|*8��va�_�<aPKV�CB Ͽ=�t��g�[�<a� =�Z��DE�eE�Q#g�Z�<	V
^2IR�\�C"4a^aS�@�_�<1S�P9z��$0�� TtQ&��A�<���J� ���R"���s���e�|�<d��D���䎴qb2�b �_u�<Y"D��iu���eʸ9�����A�i�<QVO?Y�3�g�;*�s��Mi�<�s垽K�R��'��l	@l�d�h�<�D�;�2���5eռd+BcSe�<�'D�n�� ��D�RK&��o�g�<�f�E�L�@cұUZHo �y
� �#@J��5N^UaL:,�bm `"O*����[�{�����2Q�p�BW"OnQ�n�f�V��듗5�M�d"O�U�� ^T$r!�c���:ti[�"Onͪ�JK;g�9�х�9 h�"O�%D	�b�n1��d=~���3"OF�d�� F�9�AΚ��4u��"O|)Â�
�0M�E�B���"OF�t��H��@!�+�L�$4�1"O����˟�ez���$�6QO� �"OP�h�݇qΚ����Z9�tx"O����v�z$��C5k�f��"O���I�m�PAPX��X"O�\�ʑ-i�a�"/�+�*�0P"O���"܄dRU��[s츻�"O�q��jjD������^�҉S�"O��7��z��`��!�'{J:�S�"O�YQ&���ؙ��i�t�`�"O �Z�*�s�����.�fc4��"O�-J����t���0'��r���"O�l8����3��` �Y�	c��	�"OB�(D���8��OE3_��1"O�-��Ӵ��ѓJ*X��"OܳP��,��j��:h�X�p"O�h��/$Bq�*��	�
���"O�HA��(N�1�~�rU{U"ObX��W�h}P�S���<C���r"O\�0bR"Z��9Jæ�=>��'"O�x��Ń�Mn:<���x�E�&"OjM)��<HOδ����&t�u"O��Ff��Hp�� !�6�|Т@"O�����2���4`�bՔt@5"OT���J�>q'�iIs/��0�%�"OJ��v��S�ґ�/lޕ��"O�1'�Дxe�%[U��a~�Bb"O�q��oH�G�Fd�ebJ6P���x@"O4�;�υ=��l�r!�'i��2"O:,��I�3�� S&J�2a�����"OLqp���j��a���W�z���"O���w��et��`4�د�.As�"OV��.�>6H~��"n�.B���i�"Ob�����%$s����K� �J`*�z�<�l@Q[�,H���B|��7��x�<��C�^� 0�A��5,���H�p�<�#�	îh�	�h
n���%�A�<ɒ
_3
���Z&�ΉGgڨ��QE�<�(�VXV�h�#E���vH�@�<)��Ҳq�f,0�$��.,�݃�MT�<�������X�6�A�Ut����V�<��h��Xur��w�W~�����Q�<�A���̨JF ��,�B�K�<q� �1�$!� �ۇh1�K�I�<�@M�М��l��Xz�كH�[�<A�G��S�F�ۤ�ѳDz�x�í�^�<�CJ�^A�@�9vJj�Qc�Z�<y�	¤?:['�ڸ������X�<�ǢZ�#
D��S
N: �p�T�PV�<)��ͅ|yJ�3���8C�H��`@T�<�m����l��B�(�Fg�<Qu �P��@�b���la�<�� \ �%2ҐY|X9p�"`�<�U���2� t�&�1�����k^�<��aG�zɒa ־(�f�U��d�<	�wy�A��1[� X`��_�<� :�'�:�8r�44��4�"On���I��3ϊ�p�~�A�"O$�KR%@�#�U��^9M�^�y�"Od-��A��U��(8�f"O���M��<,��W�G�^��(�$"O:��C�3����to� Ԗ��"O��H�FS4y(�X��C�tВ �"O.�xǅ�N��X�2�H]�D��"OZTh�*oaF�y�.�	Z��T(�"Oƍ뱫#E�
��9�n�i�"OL�����4���W?�Jic�"O�5[2GS�(�0�Ȇ3֖Y� "OH�0t�٩߾b$��=��lr�"O��@�J�4�b�AB�H�� B"OVE9��j��}�d��)��M�"O�p�t��3
f,hpt�9[)�)�U"O�%��`X�9؀�8���4��\�V"OD��t �4GPFP[�D� .�~}�g"O"�3D̘0΂�2��� e�ذf"O����A�h�8�J)ؿ�z�(A"O��CǇ��$�p�Bc��L�q�"O�%��%4�$Y��G�!�tۥ"O�܃3�[�`0��Fȳ{�t§"O�I�Ɇ7ת)f��oz2Y"OV�4�Y?�M0`Ɨ9��)R'"O�L�'EVk&8h�`����"O�s!n�]�Fẳ�N�x����"O�4k KU'�LpC��C�'�\I+#"O��� � z�#`�X"#�Zxإ"O"�ai�n!�-�s���$��q8"On�.�>�3@6)ք��"OR��b[�pD�����	SQVa�R"O�pp�D/ 2V�
���6<Q!��џ^$��0��r�`���<�!�$�45���@��QUyr���*�!�%>I(�+B�5���is�ζu�!�š̍"t��^�ޤ���֭a�`C�#����,��@IV �<L8&C�I&�fj�Q��1PԢ��R�<C�5�\ ��E�"�ԁb���:"�B�I!��K��`Ů��!)�tզB�	�>�,0lȮ"��� 2O�=�ȓ��P�)�9G�r�+FIQ�ȓmytPɧ��I�L��"bP0�R��ȓ!{@T��)�Fh��j0�c"䠇�0*����cO�~p�fX�D����Rf0���C��S�Z-FO�+o�t��sOr9��M�Y�"�r��́*�$܇ȓ!��5�v%
�鐶��el>�ȓ4̆,��ī\ed]�T�ǂ��ȓ���#L"e�x�)�Å�?�xT��-��@  �5M:�8�� ���ȓS����J��o�t@��B��A��`���C !~��DZ�lمȓNU�QPsE�YA�xU��59U&,�ȓ0=��Q�+;���P$c�1'��Ȅ�.�n�р	��6��t�7M�)մ�ȓAq���R�7o�* �ǎ5y'��ȓ	ʎL�q�c �=qf�.0�z$��!z)X�"lŘ�Q�'�V��xN6����&4lP�@F	\��ȓ&�"[ס!'������~0�`���B��n��Ի�)���%:D�Л'e�<OXV�y�aʛ~�tɡ��4D�� �@��,�9-�0a���J{�4ɓ"O����.Vc�+Qc�c@�i5"Ot! A�O�k`X���ձMD0�v"O��ag��+ �0��ұ;�b�(�"O���$o�7*�t�� �����"�"OB�PuE�vp��A���L��1ys"Oʵy`��#��u�%枍w��D�""O�xXV9�JaȻN��Ty�"O*(��#ʑ����GK�<\��"Ot�(� f�QJ毖(5�>�)�"O���E@¦G�>ՂWU3.-��"O L�6 �?6[a`A�,�h��q"OzYX1$��`Q�<�T/C4}�:�"O��yD���
�x��wN�#o��Hw"O:���3(�����*6>,�Pv"O��ْ��M�0��($J;�J�"O48H0�P
XN(�c�Q�qH�B "O�0Je�Z�_(�ɘ���1�l! `"O&��e�I%A���8�����}"�"O�d��JѭQ��j0&U"��"O(x�/[�Mf\��w��J�R��'`���3�X"Z�"ӡ�ѻh�J�@�'}�eC�����ؚ �4
����'��IQ`�`��J�DU0Z�&�R�'�L�RV�<)Ԅ�+��OXh�@�'�h�)�b��f�@�����OP���'l֐�2�I<;`Z5�Qj_
G�V�X�'?��І��7xĭ�q��',��z
�'\���o�>,%>����Y�$�~4(�'~>����YvH~@���	�?\0��'_��#���H=�|Z��ئ�=�y§ޅr6��@�7֞1��	3�y�FБ|
l4�A��4+RHbRe�y҆_� ���t��<d����c��yrf7QMT�VaJi��L�A@�3�ybBՍ��ك�]fQ�1����yҁΣ�L١E,$VK�����O�yb	�+T���cg`��^���[g�P��y��=:l�V�?+؀-f�8�y���<%:�3�-�*\����`��y2b� 5�$I W=D����y��50��(��K%zǈ�p2��y�N��h���Z6#��qq@t�����y"� |qj�:��R;J�cыX��yR�� p�R�`���F��,f�̝�y�jR�nKZA�vL�(����JM	�yR�!��%J�/�M\~Ջ��S�y���m��L3��AK���1cH!�y�jYya��"G˄�G⚸�޵�yrOϟ|���1�ǅM\���j���y���*t������S�AC�K�y�fߔw����	@S�q��U��yD��j����+E�탲�ص�y�IΡ��J�!NR+���־�yb�X�cODuҥ�x��O�|��L�ȓ}�=�Q������
Q�S$��i��U�:��O�5W �i4Dԅȓ`�)!�\/6��C&@>^`�ȓ|�����02�Th�O�	H�p��S"xsg�(;��u!�BN�Ą�<9x9���T"n�&�16e
�5��ȓ%��m����;$UFt9q	W�V�X��,��A�SgX021� B�1'|���v<&�Qpșcؚ m�2�Lɇ�S�? �� q��S7T1tQ�ބ�`"O@�P��يZ>�Hcdl�
��#"O�U����j���˚�?�����"O~���a޵n@�xئ�>b�� E"O>U#�Z%�
9���$�\���"Ox���iV92����ڪ�~�d"OrqƮ"6�D	)ł5��,��"O�Q`b��!�������r"O�{��־Xh�6k�-Zr$��$"O��ۂ6(ɪ�B��Δ5mPA"Ov!���
u<PBT�ۙQJ zf"O�5�)�~�+�@�k���R"O�x��K-��1�CtZ�Z�"O�e���G�cd X9U@��k^�D@"Oz%���7Ԅ�Q��xQ��;"OV""i�3 �dÕh��:�`�k�*O$|(H��9K��X�Ϩz���!
�'�<�3�@��`J:��GA[~x��'��q�e�(��:�Y�?4��#�'�:ij�L�)l����f2>>\���'�P���d�C�n0�`�+�D�'��0�%OA"l�(k3&\�+�J�`�'���IF��[�ձC����b�'�1�N� z�a�@ �/HI�'��S���;]����E�/6IJ��	�'��Q:�F�a	�vN�%F�Y�	�' 60�B�R�R(:a�B@�0,���'^*�)��A�0���Ga�!*�=�	�'��I6��D�yh"�%# J�'o�@bI8�����/	�f�*�'I�A� �Q�k��ZfD�}�y��٧q��+3�W$5�@��BgՖ�y�
�8 VIs��T�4/�uAgl�yB�K���&��lʝyEǇ��yb	ݷ :B� 2��.j-`%�t)G��y"�D7����L��rƢ�JqN���y�I����Ej[,fR����;�ybg�q���{R��mŦU� f��yr�\�k����jBV��ha 	
��y"F\���L�\)�tR� �45#jC�W�0�͇H`��,�2Q6�B�I��2�����$eP�Ɋ�\	=&B�	)� y�@�R�(A�}�f�Y@�B�	%F hȰ�9k�j}���l�B�<]��d�
�}��,��Bq�"O�h�g ���2��T�`K%"O�D�AΔ�i�d="��Ș�`�5"OnIB�@�Y���򂃋�;��� �y��ӡ}��C�/g�>T�ceѴ�y�� �݉"dT��H��c&H��y�Ē�d�Y1��#(ܡC�$Q�yB�ʹN3�=}d�<�Z1��B�	�H*�Q�#I ���U�ՐS��B�I9~�i:��ː�����jMHC䉎Y���B�ؠC#B����G�g>C�I�g���ҁ�H�q�P7JB䉕nLR�����4��j[2k`0B䉺u�����͎�f��mX�eōm�B�3ˬY��P�&Qcn�teB�"��Ɇ/R)t��8Mߝ>�!�$\�l�q�ߤ9s0��j��!��ЃB.\�5MA�o]�e ��+�!��B$\\ %�M`�X�&�G�!�ʈ��=r.@�4� ���h!�� &�2׌�	yƩhb��1V1T���"O�B-��ZLj���O� I"�"O��BBlK4|�xb����U��X�"Od� ��>$�0�1y�8�6"O~\�J�	$��Q��ۮ"�����"O�)�`Β�3E4ŋpF*$����0"O ���hLc,���1WL��7"O��oM�0�v�?{@�ѥ"O&��$��/\��	��ۍ[���[�"O��qEo 1���V�1hb	��"O@���D&�����-h?HEX@"Ol��*O	p���bAↀ`;dT�"Oz��g�F�! ��Z��U��"O��Q�͛�Y����"e[
Uv�}R�"O��!��� 1i���P��e��"ON�!� �Pa�!C��	�4���"O�̈�A��v�*���5Ԑ�t"O�5H�O�%#��u#(�F�n�C"O�}Q�陣��H�� I��9w"O����dcf���2��,:"O(�zB�����`q'�+}�ru�f"Ol!��G:Ͷ�R$%u~� 
a"OT]���ޮ�F	䄽-d� 3"O��#��PH��`'bʪ�L�b"O<�bA�	N��1!���BZU"O�!ĊկW��=�E���_��c"OV(�1��3�H{uK�Bh��(f"Oބ��g�i�ԘP�	V8jX�1�"O+�%����'��?~Z�P�V"O��9#@ 32d9�J��N��q�"Oظ��؝	t�i���5WD��E"O��[�&����b�ّEZ��
"O��#��,BQ"�eĕr��ի�"O�X����F zuh�b��&죗"O�`���*;	m[��Щi����"O��C`�	j�p�3��%l�~)p�"O�0(�I	�P � �������  "O�@�ƹ�By�4���P���"O"8����\J��Ԭ �x�V["Or�P�e��:���J\�
�t���"O�!"�H�l���*w�$5�܈�"O�y5f؃m��9�+N�urn-�"OHp�wbAf@��Bg�d*"Oҥ`Ҫ˶ʸl��'B	db9��"O�%�#��$�McV��� �Ј�"O�{���	'@9�g�Z��0���"OT��We k��t���T��;�"O<��B���>2B�k�����,
"O��3�A�t$ъ�O�Z�d���"ON]����42���
p�>Ғ��P"O�X��.Ή�x�:1�@t5��"O�ȪpA�i}�}��� �r�*T"OLi���G7
�����$���I��"OP�a�\�.�T�z4�_;FQJ"O��Y��P�JZ������U�޴9r"O:yY�T=S�)b�LE���Q�W"O��;�EO& �8�4ˏ�5��I�"O���EΈ7�M`0�]	d����U"O���$X�Tv4�Wϝ�IlŢ�'Y��2�b�pAP'�V�S�
I��'���(�
�y�=27��twf,1�'` ���a���~ ��`ɨq�
u��'�0�r$!D�-W��������+�'쾼�&�F�3�ܑs%Z�}"dK��� �t�3�������@5���Q"O���gް*"����1�e
U"OH�����O��QR�d�8�B���"OJ\���5h�T�#FG!���6"O�rצ��i�V5ze$ÒxS�h�R"O��C$��5�Q��G;O"�C"O�t"�ސ4��)�,UD�Ȩ�"O�X`�#4�Q��F<@�J�"O������	x�� C�w���;t"O�� p�h��)��h0P�"O
X�o�
v��@��Ơ+f����"O�|��V�L̰��M6dWx`i"O0�ȣ��/pX����U%Eؤe"ON���/�'x��y� ��v/�}@�"O-��B�"X��@�f-��iic"O���/�J�1��돭v�ЀҒ"O:� 6-M�x\��+F�dM��H�"O$�oO��*`�w
�}��0Hu"OLA{#�� �
����n�\Y;"O��y��ֆJS��l*4����1D� �oӌ#������	��p�n,D��b���k	�ըu'.=�pUP�'D����#Y�;���'CCg�JUcu�'D�lTl�{	�Q��䟚'��)〮7D����%;NH�h�%`�"@��x��/D�P�!EW}��jµ1Ѿ� �,:D���WMP>Ya�@(1X@�j�j;D�����S���pr�ܸ*�
t��9D���J �I�i�d��	&��A�6D�0Yd�%f�$|1��0o����O3D���#NQ�,2-�� ��G�޽[�D&D�(KӇH2%�00�!/èI�&D� &mȇO�}�߀��ı��7D��"���4����2/[K��XPG4D�Ѓ֠��~+���� N��`0�$D����I�8��Jf�W�|�\�b�.D�h���ӯ6Z��g� ����E*D��Xe`��S$�)�P�Q�x|(�S�'D�)`劗��U�ѮL��w(D�h���
3%�Yr� $zmP��`G'D��H�m�P �1� �)��$D���7�\k$-rV�O	s��슐#D�tY#��_|ԁ#N�K��HT-D����L�/0����:������,D���SnV>x�hd	��T1LI��+D��"ʎ0t:><���I".�B�A�M?D��re����"��qvPL;4"=D�,�� Y�fy��3�Ƃ{g&XJTE8D�`Z'G���Pe�J� �NpkÌ#D��C��U��pib	�78<BQ�$D��@h'a�e3W�/2����$D����w�	�D�<'���@�7D��I��[)uj6D��τ6��0◢ D�l��g
3?�e�b��\̘H�I D��zS
˨"7<�{I��r|�DA?D�8�`�^,JBz�ۖM�C,��tk=D��y#�6,�� Dk�<���(?q(O��$�<QI>�'z���7�����E�����AS����}/�K�TH"��ZXfɋ��MT#��J-����fx �0Sa(C��hZa"F�5��ȓA+5�/��9�<���C֣%ּ�ȓ;��\1�C�!(a�u)��1�ȭ�ȓP�� C �9���+4�Y���YD|��3� �� ʳ�<������xU��"OJ���܅!�Y3�05�"@7"O$�PeIS�o�8��u�ȿ-�4��"O�ݚ���"�l�.�<a�ʨ9�"O��@H'�rqm��R���0"O�,P��I6S7H��#g֚!����"O�����6^�b��a�4�4�+���<��ɕ n��5@��ǌf]�ĸ0�Ǟye!�$و �X�r7���r=q�9v!�C��ʦC�=�
��$H�7�!��Qj�(<
'&Oo�K��@�2�!�D�[ׂ�a'� &���q���p�!��J<\�`��<<VNy;œ�!�d�9�@]RqgS�zQLT��M@5>!��S����H�$���Ԗ!�^�
�~��;S2z4�#iG�\/!�$@�8m���A�r!>�`6�4Z	!�ĕZ���x��]�*�B��>!�D��.�%	�ڡЫ�7c�!�䈷�2Ds���;�TY��i�!�Dϻ0�"ܱ���� 2���`
L�F���Bx�\`���#;����J��x�4]锦'D��Ӈ.
hNL�S&�ߩ^�PI���&D����a/Rľ����;�.I;�%D�T����B����a�Ӱ��-��,8D��!(E� Y,1ƭ��p����E�8D�p�ĎƮ.I�8Ҡ�D�;rE
�6D�葶�����10��,o| 5���3D�@��A%mY<U���<^$� �f�nh<�05w�j�R�ݝ.+F=!7,Sc~�D�|+O^��]�p�DI��^4XT1Q��J=V)!��^%,=�
��,�x{�nݺ�!�M5{�zM(�Π*b��H�*P/K�!�.C�B��7 ut(!�i)G�!�$6s�B=��6�2فs�Q<U��	ԟ�F{��D��x��A��Lح@� I��N&�yR�]jM�#@�-@������&�y���=Ҡ9sp/�9/�5Z���y��Z/v�A3��,1�KR�nڊ�ȓc�f����5O	�q����;V���ȓ:�h_y�4��E�/�����4R��@2��1���TA�Nu~��ȓ9�f���5?O���LX�*��ȓL	��Z��+6�0Pť�[���'h�}y�P>�'?a˒g��T[܍"�jIP2$�,D���F����t�6#\?��}	��)D�H���@^|�qa͆���E{�(D�l"rgC*h���ʰ	Þ9D99��&D������-y�Qq������$9LO�����$^��tYT�^�]"�y�';D� �mּt�Qh�)�}ʥ�8�O����<	UG��R,ѐ6`@2vdʩQ&�n�<�gО8�H,(���9�l��Î�a�<a��	�29� åĬ5ltȚs�]y�<a�g�^�$%�FhƦi0���n�<�P?����b�6+��={4 �5�!�D�0�+�ժhN@���흼h���ȓ}��r�R�RӺ����C�w��5�'���jy�Q>A�O�"�+��1e�ϔ
$H��J���y�G�<�)j"LD�EԁA1b��y�)��EV�ɂ��޷G��P�B��y��L�)�*�{��}��z�����y"�˘(��3M�
�p�Q�&��y2�O�d���Yo�b�p7(X��O��=�π z���H��MI�.ֆZ�O ���N/�4��4Z��i����,jB�	*fi&���?J�`��*U/^��B�I�@�!�#��:%����ծ%�PC䉒`��s��Q������q�C䉳�(�A�'�2(��LB�">���h��[��*G"`�	3����|�k�"O(y��-���r��R���R�pp�	\y�[�ЖO�RK@��y�� ����Bi�.,�񄇵?D�)��Iْn�=�"$�<uR!�$��0������*8ۆ��A�S�"!�$-�HF�5fqFE8�iA�D!���7[���p��eQ.t��)�.
az���a+|M�ѽ�3d����_!�d��C�V(�ՙ,-B��0��&+E!�dZ &HLH`O݋(	�\��,f>!�d�w�i�,͚O����ͯA9!��Z�f3n#E��f��mC��(!�d�r��D fL���4h0Bڇ!�D��Ou��'DS�1rv����7������%SCL<�mǫrҪ`���?S�B�ɳfu蠉B�y��-qeJ�`�����d�<����'ˬ���\=o���I�J���\� �'Æ��B�+t�}��˙��lE	�'�TL
󎅏'Ύ�
���'�	�'�L@	�f� �ڐ�D�*�֩��'{n���r���b�� f�����'�y���nr��+F"AR�Z�'f-J`�>4��hV�2/��)x�'�jM�F�;��yb���1!���!�'�D�s�j�X�r�q�l7��Is�'�6�t%C�q(qX�D��al��'��:���g��݂q�h���
�'{��A�X�KR�H�
C�N=��
�'��:��:�	���D�~.�	�'o��Sn���~������C���k	�'�i;��� gsnua�儫3Bx4��'��}�"��)��𻥬�!-��p��'�,�*�ٷJ�����XJL���'�B�Sv��zK8A;!EZc�R���'Nl`*���%8k���-�(g0����'%�gcǚ�vx���F��a�
�'�JXC� ug~� 6�JhƴR
�'Z����ݡlTH��՞|�ZD
�'��tBUMG�E2-��-��uG�z�'���С˾m8�	�@�g�h}j�'b�Sf�m_���L9[��X��'`X��Q��'4l0j%dL��\H �'A.�	��	�K���6jθ��u��'p��af�U6:{ء�5� �x�:�'�i�A�Ź1g\�b����ؙ��'^lͪ0�ϵS��-���)E^�q�'��d[&k �8��*!Y�����',�2��F�B�`�A�$w�%a
�'��|�雠qb|!�P�KϚ�C�'f�����#	0�p�%K;,�N�y	�'�t1�c	΃;� �& `�ɻ	�'�ne����ԝ�W��"�
ܚ	�'����f]��էC�����
�'��x��V��%k�~��	�	�'��Y�o�P��dr��	"c���	�'�@��g¸T>ԛ�-�/�H4Q�'#�P@�4̠-p� �~�
���'�1)�A�\�.p12�֑.������� �D�d�,�JP���<g�"��P"O�d�e���xjzuȵA
'T�Th�"O��k䭄8Kr��)dA��mm���"O����"C(����b�5
�!j""O$1�%��!��@��X�{�b�h�"O���S���Cd��c�Z���"O>U��.D#��Ӷ�ܜx�l�XV"O҅���Y=nj���r��>�
l �"OѳG�>�@����6ds�"O�!%��~ER"�h�����"OZ���Bء-��S���w���jB"O.}��`[U��y��ZӦ�z`"O�,�t�ɺ�>���O�8*�
��"Ot�s�ٺdϖ��Σ��0��"O������?=�a�T�R�Tj���"O$Q�%[�D��a��\�Aw"O�,�cN�� 9{���N��)z�"O�H����u\�L�����y�u��"O,�TdS�4���V��(K���y"�{1N�"`Q�B^�"�]�y2 ��Q젤���u�pA� �y�f�+R���� @;c�$@&�P��yZyi�D:��K�$��`��LCdB�I&RK$� �-"f��E[����ZB�	��
�x�`������/\�fB䉢*�NHbF�5�$���-i+,B��/y�Y��&�L�Q�vG��qK�C�	+O�"�*P{�0�F_-%��B��^���-��3� �z�B�	2P�hhp� �-0�
��Z�t�B�	<p�:��l�0C.��Ӥ�� ԘB�R3���n�a0�H���E&<�(B�:$AB�#H6<Ӫ4�ä�E�>C�-^i�uX3�^��lP�UdM�B�	����'
�I�,�'A��xC�ɪ t�=`��·g�RЀ�L�~5>C�Il�lQ"��,}P��5�J�-KC�	�I_l�@7��3-�D�zk�� $�B�ɥ6����X�$�kw$�c�"B�I�#h@0!weکd�ZZ���UHB�ɦ8�d��n�)V� l*T���C�I�tQ���cM�w���Ö���N��C�I<u@fcBF庴�T �e�B�ɳ:R*u2���6ì����-�"C�	9�L�I�g ���#@ E;(C�O lh��/I�x"n@�� _C�I5��2B�(s�F\i�k�>Z�C�I=B�4YT�,8	h	%.R ��C�>0��,�t"�0=�!e	U�4�fB�
.ݳ����}*~��E�,apC�>;Pvx1%��/MY|�@�،f B�ɡM�\�Ḋ�Q�r�13A�&�B�ɧ8�	�V"U3H�T�`�BI-�B�	U:���A�:=��m��ÆDo�C�	���}r��0��i���Zf�C�	9RXD��5�4D��i�gT>3��C��/w|��0v(�nٵB��C�I�^Q�T�����MF�yf��1 �B�%S�@�W�,����uH��EIxC�I�Q��l9�ʝ��\��d��?�XC�	�d���DP'a*�����:')|C䉚O$P��G��zn�r0 <�PC�6j l��㍝�wJ�#3
-�:C�ɟX9J�H]�\��pue��8�VB�)� JU�6I�%��e����<w��,@�"O5r�<=ٺ�;�KM?�(�A�"OJق�e\��4Q�6T��9e"ON�KQ뇑`���Ø�#p��"O����Fɲ7p t���=g�	��"OpM	m�<\�d"!,�@a�`�g"Of�Qpd� (�9��u\b%	"O0�3�dڂ�|��IS�����"O`S'jR�0E���	>P9HB"Oj$4iNf�69j�U77�V(��"O��낃�S�J����݆`�Ġ�1"O��Q�d�0R�M)�d�7�4`;�"OJ�be^�B΢��D#�e`6�4"O��2��>[��0�h�~^LH�p"Ohq���ٙ=m@<A��ÈnjDL8"O����	; ��E1 lO1��ɫ�"O��eF�2C��jV�����s"O�q#��"�BL:!�X<~ A"OTQ�t	I�]�9��F]�D����"OL�&MX�(e�L`�,�0k��LJ�"OTtȕ� -�j���\;"O��ps�]�@��c��jN;�"O��g��D�0��ŕ��ce"O� �%�D�}��!�9zPP""Ot�G��6\�ڰP�G��&*�M��"Od�J�D�/�܄�R&�47 ��a"O�5��㞩����N�� �"O� 31�ސ!2�ItHK3_���2"O@eKP�M�S~�*���r���b�"Oi�QJ#���D\4i�FhS"O��8��W0H���IFF\��;�"O0e�Q-F3wr�ғ��M�A��"O���KT�$TT�0���-Q����"O╛�
� q�H��Ä7F�9Yf"OX�E-�P�������"O� �CH�	������eQQ"O�|+�ϗ�a�R����#x�h X%"OL���Ř*]�pt"Z
;�ܝ+�"O� �d�*~���R�@�J�̰��"Onto�E�
-C�i��"f\T"O�Mh��M�{�:��꟢f�tPZ�"O��+1F[���D���v�C�"O@ya�?:eX$3f�\�
�I!"OZ��3c�*h %;�K�#[���A"Oz�K�n��IH�|��d�&TR���"O><(�*�6lH���L0:��E��"O^��Ą��<)��S�A�<w@�� "O:���{�T)�c��& ��b"O�$;D�x�R�@3`�'K� �7"OZ��Ö�19��B���=WM��"O���JNp��Bb���ⴉ�"ODsЅT7N��A��
�)��Q��"O���E�
�*)��+¶F��$K�"O"���Ċ	��T+O�,��ܒ�"O�ڧ�5"�&i	A��6|��T�V"OR�*�
�"$���пJ����S"O��㔌��[V�S��Ûk{�i�a"OPq����l�L�bs�D�G�Ɓ8R"OB�	d?=�@HqBK� y""O^��aE�n�PK��\�T:%"O�����S,&S�"�'�T�ب��"O<XRU	��o�\����b���[r"OB͐#HD�	��JVd�5� ���"Ol5{'e�T�+�-A��RU�c"O� `�16��%f���F&�%�<\�v"O��s��SP����X<�4"O��[�D�m��h����N@�"O��i�)����	d�y�"Oh�PQC�5C����G�CN�4�`"O�`�ˇ-���S��:��"�"O�բ���)�D��E�Yɶ(��"O"9Dk��d��)@
"U���"O��{։Й���z􌌚_���k�"O4�[1a�:�,��W��c5\��"O�x�B-'�Qс�J�@2NX3 "O2H!�֢$]~�R��^TJ�"O,�3H9$AUТn
�sP���"O�Q��aT"]zgoZ#����"O�L���D�sv�슢mo� �"O`a�����v|��e���j�hw"O� J�j������� �"���"OP��BG>��� ��084��%"OB�� �JrR�C����z�pt�A"Of��5�^�F7��K�AN�͢�"O�)f�U�d��Q�R���̲x��"OڐA���YA�0�/̜Z�d�*�"On=x��[�6��;(�=���"O���E�!3�  ��H���"O��*!���RTС�[5m�,l��"O�	�"aϻ�L�T%]��0)��"OX�{WH�7d��3KT�s}���"O�q�ą�_ ���/K0k09p�"O<�I%�
B8 �����
k�9��"O��.C�=?hI��NS�~�!�"O�,A�g� (�<�ږ��3<u��B"O��#� V�BRգ�	_Y�q�R"O��xp�@�H\y�ӟ�h��"Ox(K׷�.���'܈w��X�"O|�C��c>Ȫ�C�m�E"On��M
 �$4{�'�)��8�"O��� ��.m���(�,v����$"O�i�u*��"�z�L�"OȨCq*T8���[ M��#�~5��"O�8��B�`��[n�z��� "OHT�e�H_�ȜA��17����p"O6���J#Y �g�(w�Г"O\��T�=��uƘ7��+�"O�}sF
5l��!��V	 y@�4"Od0`��ՠ*[j��#C7_x�9k1"O�T !mD�<�V��sH&O^��A"O<�!!)N4����3c�D�˃"OE���:�%0�`F�{:4�"O�%��oa< �eO5od�Y�"O�dqba�'L���T��j�,��"O�(��ܬ*�(B$�;I����"O�=[E%B,`���ŀ'D5����"ODDhuM֯I���9�d٨V�Xq��"OTE���ڤs!��R��3p�荩4"O��"��
"Z} �X��ΒW�*8�q"O8u�DN�:-�* �1c�)B�f�T"O�[�`Ϋ!0J����G�� �"O�0�Ij���	�Ҝ��1�"O�PhS�g��x�v���
���V"ODe�� ~�J�cB-F�O}�D�"OTA��$��(���A�]U`��5"O$�d��?;�hI-�D�/!"s!�$�2Zг���&v�u�5�]�hi!򤖁gY��#/σ�!���h�!�� DTc����q~��҃	P�?�&���"O�	��bD/�X�k��ӃtКDK"O�*`�=0F�n�Jۀ!Qv"OX=x�L�0�z��܍<_� �e"O���cI�V{��,�0_�t�A"OZLxs,؍���"G+�|t�Q��"O��!'�եg�������%n���"O��$A��@�����8k�Y��"OfPA�͎*e� 
�E�^����S"O�p�&̗W�)��Nߊ���Ѱ"O�%;&���i{U�Rmvz�RA"Of���	ZU�>�s�e��~y��"O�A��
?[��ݙ"�9H�l�U"O HS�h�77{*e�0����r�"O��h�.K�Pc�����^�zvHZ�"Ol�Є�="VL�F��8��+D"O�-�©-=�h� g�ˡN��� "O���P��uOd �!�x�1�"O$�0t��-d�J(s��e��H�"O�x5%�zBnI��d�#~�e��"O"��v�'@� 1�#�4m0���"O�qKD?4x7�C�<��t��a/D�̩�C�2a䨼�!@XZ��Y-D��1��Uc|��å��5����*D�HPW�Mk�u�v*�'���K�f'D�Gd�6:l �E�>fL���%D�H�'KD 5�QQ��%U�H����9D���#T9k�4H�)��f*F��7D�� ��Ȑ.�X��SET�6� T�4D���Î'�Z`��/�>�*Ԃc�1D��(�m�B-�uQ⑅
��=� *O��S$F3\������Z�e��"O������T��y�f3�D�P"Ovx�p-{�x9��c�b<�X�8D�����RWv����!4IYB�5D���"#:P%�J�--pbt
g�1D��sG���ü�cW8K�J<2�$D����`aL�R� x����C$D�4sU�փ$��8�'ў[�+E@!D� � J��e \���)5�(�á�*D����*ˢK0X�Z���h��u;�I)D�T�EN�D�dp%�ˆ~�bD�q+)D��ɡ;C����
������$D���h�&|�lR��zZ��0(D��Z��8tC����,��I�DH�v�&D����t����(�+�py����<�W �+L�^KҌͫU��d �f@B�<)&��)F���1
�"a�� �aP~�<ѕJ�/shi���)�~��� V�<ٗ��u�y��ϕ��.}��%P�<���Ά�fM
p�L.�pmä��w�<�M��]�{�@}ۤ�2��q�<�b�����L1E��  ��[�LAG�<aҭM�a���RF��8S!�A�<���*~M����os����F�s�<)�hC*EvH�sņ�0@p��	h�<��d���	�KS�VəR��[�<Ʉo�#��j�8F&5��V�<�ɐ�\��e�J�:J�l��!�Q�<�� GB`���Ϝ9H�NQ:�Ct�<q�k�'٨��d�\�*��TVͅo�<�v�J�x���:u�U���n�<as�ds��
@G�{�����/�g�<V�(:��P�kM�A�0��0�Cb�<� ��(��t_�+q�]�/��:�"Ol�c2I�%�,�&AK8 ���F"Oj��c � +��<���'�~M0"Oؕ���3'�d��Iz����g"O����(ʘ)��]F��e/_d��9�S�'+�X�x׊P��DX�� Po<�ȓl��!R���l^H �؅)d(��ȓ'CN����htl�7.ҹBT�ȓX��ك@�Ըu�Dሓc�aA45�ȓDΨ�"�91��d01	Q9F����ȓH�j��f��'�jɪ� Ծ0m�������,/���@�V�X�D��';��6lO
`:��K�]&	�9n�5S��'*�D9��[�X��8�+[*a�z��"OT�,B!�6`=�S��b�Ш����c�!򤑭-��S�'�*�x��u�ϲ�!�$K7����@P�r�E��֟�!�D�O����ɡ2� �k�	˄'��DI�"O���'욿|Y�I�5i�?��� g�>��.�S���~y�햜x4z�����4N_l �ȓ��ȡ���'P�	dcU4$�dx��j�2�R�͉# �=�b%�39�=��4c��O��ɸ|j���Ri�t%���8вc��e�<��M �1`����O_N�fE��Tߟx�<�6�)2�e���l��/� ����p!�Z�<a��'$=0R�։^��kwcJ��hO?�"(�Ɓ[� �a�ؘtHC䉺=|ʰ���̒2J
��@�R�2�m؞ 됭!<Z�x�kX����X��1��p<�S�=t���OMhe�g�ôK!��+P�:�@!�W�%:�+-N�p @��>�������EH'hRT�c@�(��U� a}�>�k�#u��[b',��4C㠘q@�F}b�	8{�
�Jr��h����֞{�B��0@7^͋��׊r��Q��y�fB�I�������
 ��=�$+L>-�#<ъ��?�$셄R�"a�G��/t��:."�Ig��|���Er�]�')H�/�2���'%}��Ov���|�RU*�c4)l��'�V!���<��$G�w$
A�סX&0a!�ԮR����r-�y�̂���4{!��N�n��Tc7�ɻD��/�|���)�����O����tA�[΀Ѩ�O1D�����c� "v��{a�5�&�ώ�M�E �O$`�#�w���
t���]�pN���d&��6@�TӶM�1F�4����,m���Ɠ_��H�G�S�M���HBc��A���Dx,�S�T�e�L����v��yY�Ƒ4��O �~�G�h�ʴ�п@֨R�%BU�<)7%�Lddڅ��=WߊL�ƆZ�<C�<h&�3�h�� l8����j�<���V��@A�6h���!�d�[�<1dbL���u��)w��	�	�B�<Q CF�5��/� �|̓+��7m�xi�"��q�չ����z�v�y��{ܓ�hO�y`����R�`� �ރdp��p��L�l�p}�
��?�}&��������s(���'3ʓ{y���(O�R�T�>M�T!�(ļM*��>��m�I��Ԉ6Ȑ:��jL`��z��+ 
zP�	����Yt��������G6�������~��X�?���'	F���iW')C.���S+c��`�'�j�ؖ�M�PH�AiB�����4�Pxe�"�D��%�1���'F��p=Y�O2�D�O� �i�4�*y>���R==4x�0v"O")K��ơa?b�	+�3/ ��r���F{���F� ��e�4�]@`�H�N0E�zb�'��'06X��%��d�;F�E�e����'�	G̓�HO()Â@K S�2��+�,'�րHB��2�S�	�=R�J���$v�,�3fN%G��'��S�3��$*���6a��7�mx�.��c+�AG{����<���߿2Bb,!�'�Ezh�_�<�k�XR*��am�R��mQ���U�<�$S�iވ����,�n`i[Q.a{��$�7g��M�	~ߎ<�ЃU�!���9e3�pY��BXҊ1�v�v!���b���(N�R��i��蔧mb!��D��L)F Q*v�.�Z��J�+vaz�����l��7�8���S1u�!�.;ϚI��n�Ƅ���0��	c�����ajם=_&�H$�?<D1�"O:�*�͘n<���0��3/7nQ��"O2WY&s��e�ՠ��%Jq�p��M���:`�O* ����[��!���*.��(C�"O�\�E�)3�(�@�L ;<�th��"O>�!��U�?檵@���npؕ
�"O����(eB�!��	�i2xE"��'�!��ߪ3������6T
 ƈa{azb�D��^����Bl8e��yJ�N�)^�!�d.t\ȅIK�h�*���o	�b�1On�=�'4{�	%MF��2��L&�q��^�`�
ʓ�hOQ>Zw*Q�ub(%�bf�������8D�c�ў`��U��6��a�$n<D����
�(M @�p�?f��v�8D�@���;�Pyw�AD��@M7D�D�3�E�Y��c'̒�L`��e4D�l	��Bp�>�#5oί0j���D/�O���'�Jj��Z���ÇV�E�jԹ�'�	�(O�nQl]�!��0<'0Y9��p�H��$��Zep�e�4Md������!�d�$L��㧍�C�ހ���A�t�i�:�D/�)ҧN�.B�A/OB���'Y>_Y����j�-IXx�t ޡI��<s�-��7P�䱟���I��p�X�\�RY舳a��("gN#=!����?!�̚4�>�`�Xv�H˃I�i�<��m�#��I��H]�
eL��⦁�<!���ȟ�V�ѓlw�����ϨZ,�ʄ����y�ć'Wۢ,A%AVu��{�h �M��D��7-!���	�H1�� 0	�J�DipG��.2J���k�0�I�4��Y�����b��[	P%�B�0;>��{��ء�b���/2k2��!ғM͚%h76oO������.� 	��=���%�@\du���r���������q��84|��@U���ȓzv��;��5$�X�%A)e�X�ȓBdؕ��E�a��	k�ǟ$l������a�B�zH����ߺ#�����w���baN/����@�Z�@0���y�0��� �R[�,�@hٞ �ȓIʨ�C�H�pg���p��}	8(�ȓ-�jq��o_="E)g(�(-v��~�b�3ALͫJ�m�3�T�ꍆȓ_�>H�r�}�0�I��� q1 �ȓA��`B�`�#\�yyf��;���ȓR�D�Z�H$immd �5�h��|�^ـ�R29T�-9s$O/B`2��1�̽"�}��=�łǩ"^|�ȓ5�9�dNٔZ	Lmy��ΉE�Ն�S�? �$y'M�\,�ԛBgܚp2��3�"O,;t#����Ϡ8���Q"OXm��H0c�Z"��+l8HyQb"O��*���8BLM��![�K�)��"Ode1�����[�#�  6�e"O,(�j?Wܙ2G�G%���'"Or�2�e��>!��pB�4\�j�"O>��g�G+&�.H�Pa�!-����b"O�`.mr��J���,~=��Z0�y2�\7it1���z����C�?�y�c��TzZ0zC�ɻB�����y�a�h@�d'L6q�0�:�)��y�ǁC�d������`�^�y�Og5��5j%-�J���(["�yBe��bz��Jc�!,32���Py�	P�N�HTjVm�t��"co�c�<FFI�#��@FC;�h��`,�c�<� �$����A�ޔ�qjJ�<I"d^.>=(�
�
	��.�2��B�<Ч�8��U٣�Ͱ13F�K�H�<�(
�,X��J�j06H�MZ'�n�<q�Ȕ��Q��P(�F,b&�r�<�O	����T��V�^�A%��p�<��B���G,Ĺ7v�E1�Q�<�V(� f�����e��<|)Q���B�<A��R�04a���5VfHK��E�<!�i�+)��q(�Ř3�~�A�j�G�<R�+d�y�a��q�$!Y��GC�<� "�!@����N9�~Yx���B�<�B�M�^�92�1?���-]~�<��@6A��UZ6��+o��Q�c��}�<��-o|�zD�v>���}�<�����scB����	cH���Kw�<�eg�=$��E��EBv�I��L�s�<��D�,ysF����G�cN�Y��p�<a���Jg�� !
F�P�
u�<cL�$���[�Y2M����/PF�<	�͓"s�J�$_/��-�@��h�<C&���`�1�)%<4@����^�<��L��\��E�Zh0��]�<q�S(/.hL�#-]�fv�i��S\�<�#��N� ��+^.-̚r`Ft�<q��8:c��"�)a�L� CϞm�<�dj��P�4�����>�\}h��Ik�<I!�G3_�"�0@�w�X؃.�j�<i��F6q�D��%ÇA1����Üc�<���Y~4ܛa�0j�2�i�N�e�<���Ou ���B^�Bψ��H��z!R�X��=3n��`�)�&߶0�ȓ)Z1�pe�|h�U1���?Jd�=�ȓe���郯7�ʠ0J�"e�:e�ȓ���z�牋`�Ha���ED����l��0�V��U��& W=�VX��55l��R1n��٨�F�X1����l�`@�B�$r|8c5��5���ȓ{G�#/�*5F���*3�0d��1���ѪZ�z�Fi
��X%B_2���S��r.�8��	@�)>vȅȓ/�n��t�O�D�����_�P�،�ȓs\t0�6*�~ۨ�C� ^
R�X�ȓXNظ�f�°1��U;�C�i�x�ȓ0Y�r� ލ(�8��s��
y2���8�VM�'�
�y���ʑ��
x����ie&�ˁ�ϐ`�R�C�'�\݅�S�? �%�g�&��)(5n�?"D5Y0"OZLr�LK
�f1ٖo9k��Z�"OL� ��	," �(U%�7d���=D�t���?m���Ǡ`e�ਐK;D��9�$���}�Sd�-���R*$D��jR*�w+F(�Ų(�8l"��-D���V�ŊĐ�T��6D�����¯u|���ިn�8��1�(D��83� j�eƘ�v�e5*D�(s&>vL�2h֩p�ΠT�5D�hcSM��&W�u#$�;/ vlI��3D�h͔j��S���W��K��3D�Ⱥ��ˢ��93�*�.=��M�f 2D�Lbr%� B��B���5���s�.,D����Ņ9�\T��)TU�����/D���p�.�B�B�o�6�Sr@/D�b��ϠY���r4�2W�)g/ D�,���W�_ƶ #�)]� M�G� D��y�dܻ���:`�آ|v�$��m9D�غ�ױ?rt$�L�2z�d��2D���$�3c ��ϖg��!bM$D�3E�^�T� NGi_ԝ��#D�|i#D
>&�P̲c�)_�I�F�5D��8�8y|�cfoǃVmJ"�6D���%d� @2Pi�e��rs:�@�k1D���'�G@��f4 M	P	+D���BhC�r\���B%q$�P�ԯ,D�P���'!�������y3 � D�1O߁Z��I����0iCXuv�:D�$.Y��|�g;pK������x�!򤖸jsV��'�ّ�U�*G2E�!�Ē�B�Z�Rg�.u��=(���m�!�dVI3d�գ(�&��`UE!��BΦ]�s��%%薸�D� �B9!�$�U	
�u$٨ݫE�E�99a|��|� �)[� Ё��^���qi�9��xr�V9O�Y�@`�89���(ʨC䉷|����G�2�jd�7�C�ɱ�v�&EÞ^^� ���p�@B�An}��e��Hppr@��WA�B�	;0T�ɱ�"�a#h�{���B�Ih���@�
C�%���8}���䑘(�(a("%�U���s@K��!���z� ���T�[sP(�$I�s !�$E�dz���JϹɈ@�&�!�dX�7��T��i��'�Ũ�fD>!�$�S#��QB��vH)#��݃_�!�D�e�IvI��*����Ť%!��Q "�D�;խZ�J0X[�O+,�!��ټp��x!���nT[��ҝ�!�� Դ���%
���Tɕ8?�!�$S;aܢq�p��6�
�@�܉i�!��`*~�(�@l����H͟w�!�D@	0��x*,�(��Ѩ�U�X�!��ЪLc����S#�|5��'^� �!��C�/�f	Q�_.X�*ۆI�"�!�D��{EB��ueӗ��,k0葐k|!��X�h4�T�VQ�T��I��5?!�]���R$Wp�,E+T(B�"!���O&�c#�B�Z_&��G�L!���������E"KJU�B�B*!�$K=j�]��F�t�0�Z�商i�!�Sx�uk&�*q�,��t�ϘI#!��N<l|V@2f�Bb��u���@�!�� =��$®x�����Đ.�$���"Od�� �#vu*�S�ڌ<@	G"O�8��]�z�Hq6�G�����"O:p$��D�s��q��`��"OH�;���6��`z"+��"�t�J�"O��Q� 3g�^��1�u���P"OZ�5%H�K��0ju�ȪL�6�"O`�ق.�9�x9ZQ�/L� �"ObZf��7t��A�51JL��"O��z,�:r�)�P�P)^+,���"O��8��	6�n�(�iZ+����"O�<���H�d����+�<w�X�"O����4ظH(�V1=�P +4�|��'�q[3��#K�z$�H3:���'�F$	�A o�0�y� U?B�2�'R��k�a8�h��`m��5S�X#	�'\e"t/A$?>I(ЋW�4�t\a�'d ��VG�D٘0@�A:/��%��'�RAB���o��ih�A�)~����' �!QB܉J�D��&��vt<�H
�'��b����]c�c�w�.�C�'�ҸA3,X�B�8�`�mA^٨�'�|XR딺B��Ф+��6FDy��'��x3���s$��b�J�D�RL��'�
Ual�>@��PpS�A�<���J�'p�fT��y#ӡ%Ȫ�Z�'��TB�B��Au(ܮ!&���'��׍˻< �Pݖp���'C�Aǚ++c�Y�Ē�nl �';�� ���r�`Ћ�͟!e�V,��'� }tgZ�w�*T
W�4���'�Xe�� T���D��@�Q�^x��'!v��H��/޵�@�|���	�'��X�J�D��ɑH�"N@�M>!
�2����A�w8c&f��665�ȓQ��9��1!q~l�®�&c�*Յ�u��cʎ	�l�A��� �b�ȓ{��R ��N
()D�ܜ� ��cb���G�4xՖ)R���)��,�ȓ
�Y��B��{�N!���H�N-��	7���g�ߏv�0B�FE	-`(u����Τz�)����$�n�����n�<92�T5�R��7�L�6.��a�dYi�<��(�H��	���߉ �����l�<97�0h,�k�Nď?t�sWf j�<�v�ɐ\��{&�/sXA�'j�O�<�7mQ�j�v��P�]�8 80sRN�R�<��Lیi�F0�vA?�,	�F�/T�����D�B�Fp��"Ҫ�N�!��0D����� ��H{�k� �I�"0D�$*VI�L���Wc
?��=X�/-D���܀ge��j"��>CQƱc�G D�t�RG��K�� w�	*u�ĝ�+D��9�`��~F�BAL8`��!�+(D�8���!	�%+��B
HQJd�$D�|r��W�;�
�'�~y2�!P�$D�0��M��]���rhH�NP�CW�=D�P	�'�$~�p�Ħ	��[rk!D��{/�+[�ʔr�fB7"4d�C�>D��a��0����g8[��Y��)D�00���q����@_>Y�	�&D�ɑ	[%� ��
�.V��I�$D���W��R���X���p�L�un!D�,�@������ɷ>�`d1�K>D�� dU����b[�)zCB�Bj�F"O�,H�/�u�P$X��\0	OhuQ�"OX�F.p��܋�!�#K]���"O�����i~<�2�2~>��3u"ODeC��ŷX�A"��]�K.丒"OVx�$Ő2(4f�2�K?>��8��"O"�{��
�C��B���>��U��"OF]��T�eFT!H�������X�"O.�	�`�	.uī���8��"OT��b��f���H
sl���D"O���dT'���c��1#u��"O��	`��&b���@lݥ�x�"O0���W�^�yF��5E�8�#"O,����p� �����l(a"Ob��TbH c�X;S��p+�Q�d"OxD�E�)s��A	ȟ+X�"O��8�7\�bp� �A�:��.�yZh ��tq��Rs�I�:�H�'Pޤx�,փC�	2�d��gpx�X	�'��&�0z�� ��g��sl�|��'et�z�N�톽�w�/g429��'�J Eǆr@���̝hH����'�!�!G��A�n�WX7|-y�'e�����E(:���fMa�0P�'8D�3n�r�qF$PSF�(�'b�X�l�����L��Q:�'��X8�N�%gH��ӎ��C�Z��'c���fO�-��()���-�Ph
�'�D�bhB'���b�.(f>!�	�'U�m�v�ݟ.Х;�\*#Vx��	�'<:���W�H4����	�j��b	�'Y�����Z�\I"2.V���	�'��X�R��?*�JJ`��U�pp�
�'� ��e��7ݙG司S��0
�'�e�0n�����L»?%0A2	�'D���@�����&�ĊT���Ċ�YTS��'z��k�H����@1F��\|�':f�(����Cd�ՃG�,kƴ��'�n� AѠgj9Fq+̙��'C��J�JM"}�i��
�s%�lX�'l¤�@��+:��P۷Nʜxf]��'>��Xg Ov�l9ReͰv\��
�'�(�sGL�v9fi��^�d� ��
�'�bM����Qo����[0���
�'7�4�4��2"��b�JDH*d��'��A&ǹk`��C�-N�� X�'���gJ	]XpU3�M�N܊T��'�A�P#�.,��ٷk��?�����'�$eI�d��w�E��,��'��
��*�|P��g�9LJ A�'c��j-�c��M�7�O�{Ř�p�'y��q2��P� ��7'.d���'g�])�/ē0�@�*@�)���	�'Ēi�eCmS�4Z%(Z#I4+	�'���`!g� [��$/��p��#�'?��H�*��>��� ��I�̫�'l��Jk��<�u�K�V�����'n%Sb�'1?T��N����'���s,�<TT��#JΌR��C��5)F8Hj�#�A�%��?�C�	?��-h��6t���
q��3qL�C�+ �=`ăP�r���Ɵ\�pC�ɻ3���Yt*�z�x�S��٣LC�&*38�n�6$���p��;M	^C�)� �]륤�1Nh��ĩ5nlY�"Ox����rs���Ń�=�<E �"O���1�	6露��Bڢvt�p)�"O��(`�}i0�B9{�]I�"O^-�PK	��j��� V7l�-�"O��h�s�$�xॗ�u�0�y�"O�}����r�2U#��rU��"OШbc��4P<�u��Ǆa1J��W"Onh��EλK��y#���.P��9#�"O���?>���Os����� $D��k�Z�rmcQ��-Y�|�s�#D�Q2e���#FXQ�8�xW�$D��c��ڱ[�4�e��xhƬ$�"D��)smݣs�&���׹]Ό�q��!D�t7õX��m w`2��=�U�=D��bc�Gv�&�(T�/~�x]��%D�䫧iL�K<�lJ�'΁*�fŠ H"D�,�p�75"�ag�n�
LH� D������ DB�K�^�u����0Fzh<yѦ̙�@�tO��Wmnx�Pm��D�?!�n=Kl�a@��B�ؓ'k
l�<���s{����Po,9���l̓�hO1�JEԥ�*-���'�j�<��"O��e���0�R熈B֒ ��	Rx��(b�",b�J$O�J�����M7D��!���R7�%�K��$m����5D��;��Ѽs�\a+!`��||�c��,D���vH�d@�jW̱#$�Q�'D��xסU}D���JD�����"D�k��8s:TɄI)���3�?D�\0�W����!��Y�L2*��?D��Pf	5	�ܜ�c��8J��{T%<D��h&	�rT�r��`z�.D��/��@Ǻ�"jדQ�I�7�2D����_͊��B5JF��!l�FC�Ib8�Kb��#P�򘒀'X'T�C�	�9v���3�^�w��@#�B/L,$C�I1U���h��()�H���? /C�	&aJ��@ckL�S�~qQ����M�$���4��b�Μ`��j�np�Q��^rC�ɋI�N�+qɒ�7�~��#�V�o�B��M%`(�3�'waR<C��U~��C��5H}����FմFsV���S�`�C�Ƀ[�����/qjR�"�P��B�	�3�0������¬�V'�C�*B�	ߊu�.,0��̰$�J0�B��?+n��C�	�f$�Z�b_,V|�C����ʃ��0g�f�#d�]- q�C�ɹ��٢�',s$�T��on�C�I6|� :�CQ�X�x�g��n��C�I�� YO�s���Ju���O�C��>g�l���=
Ar�fS�xŔC��
>A� �畫����l�j�<C�I�:u�Ժ�"[:x�(P���(B�I�kj��W��*������D�B�I�Ux�fUg��p���,&�B�0M�J@��DPqolh�EA�B䉵/�2�2��WN|�t�$��<^��C�ɹ1����JN�O(4XP�҉V6�B�2zְA1B�0`���ů�6?��b��;��O!,��?��M˒N����� �$m�}��2D���3�@�;\�1���O* ��j`T::���K>aPa4�gy��'�4ۇg��7��Qa���y�A�5�PX�W��+[N4�9c�
Z�hC��}Z���)�  �9eO�16� d��ꋱK�)��'�tô�ʳO�9�:O�FE�Li�8��R�Y�X��G"O��E��=PPA��(*�٪��|�H��)���0��]��D�T"͇Oj֩3� J�V.��y�-S�
t�1���9��Y�G��V�(E� ���I�=L���O�H� �b�,a�N�(���'�d��E"Q����Z��ex ہ}����E@`�e*؇��퉝H�HMؑ�}�Xpr��c�֣>��h��1�뀆!��p	�,��uWBgJRA��Ҕrr�}@ī��y�,R�:�$��eGаj����3m^5�~a�>��Y����l���[vIƝq�>mX���T��E�Sؖ	��=s�D%D�X�w�Z6��a#�&z��j�~Ϧ}3�
�0�v]��h@��X�O`�O�h���7|&�l��H֜R��M{T�'��!TB�6>��Yt̟�Q"�E`Ma�#Y�F����A�1�O��肣?~�ȝ?��Yp���,?����� :�ԩ�#,�E�t� U%��rf��:1Z��*Р�y�ǂ$ zSCi��Dv i#f$ı���XH���d�1"#�����Ƌ%T��C ��F�����9Q�!�d�Z�U!�-�9��ͅzc!򄆟Q�!5G??ђMH��N�1i!��<ȱH�+J0�؀��6Ti!�$Zs�<\��%�[�bT�C P�O!�H5mt,,�5`�?�R�K�FM=U?!��գ.��:Q��7�ܕ����)c�!�䍟\�.a0�+�3"�U��?$�!��+0����><�,;R�9 �!�D9ˈ :�K�5{)��iԂ]�uva}E;��,�	��L�x�a��,���f$z����&�$��^�ԇ�3�Jy����q�<�`JC�
�*#<p���f)���r!�O�`�A���]z��M��9!����õU>a�����O^�� �ʣ���B��35Z���2��
��,*!/��*�=C�e	�,T��0���?�O\�]�K(���ïS8�±@�,'�C�*P�X����'n�ȤaWHBo�:�	��q>`��+t�r(1���P�^�(�`æl�qO�*�E���d`�0xJF�I�'�HQ�q�G(Ly�Y:��M�>�b8��ְ���g�$0F� �#�ƒ(;b��䃕a+���iѯ%��at�N�
�1O��y4
�/	�.xY6"��>��
 C�����L��`*%�0!w�tP��"�C�4 "OT����ԬR�\��D`�-�H��2��X&Z�z�9N��(�B䀅"�-S����=\L�ݣt@Pl�.	�DL�I2��TC�I�Ept�c��6c`���,L����J`[��N/Z�l�I��\�Ds~�[$ �fk���<I��̽R_|�����9#��YFm8�x�U'��J��p��T+��Is��B��q�!�c�2�{5��;�TXD0��a��>V�az�&ߐ<_��Ŏ> �q��J���>#�eӁꋫ�e�I*��i!ׂآ�`�U�6����6�9D�����U�ND���Cc�<1�\�x ZQ��`�X4:����Vkڥ��`�~v�c�Vth�杈{^U�O~"p��0�&kA��(X֤���QX��cO����|W�)��-ǋ6 �u�w�DI�J�ӷ� -�j�8���}B��T��y\��b��ь��Đ`�
 .ұ��ɟ!,�y ۋ(�nȜ''�(@τ�m[��񒊙1��Z��X�(Fx��eJ+��E s@�)�p=ɵ5{��i t� �6\#��C�I!�<DĐY�6x�gI�@�&u(��C4qO!Е��rt;`��=Fl�l{U���!��D!�"O���WhЕ�oL�҅�V���KrH�a���FS$ h
ɽ"�t��@U:��0Q �!?���JcO�4v踚q"O�8�P���Z(��.ɤQj� �����0�T�T2�F�2s�0�aAR����C_@�(
�_�<��ć�/u�zR�1�&��%˜P]m!v�B�U�DM1� �j��|p�/Ɣcƛ���()'��IX��ħl7�=B4���[y�ꑥ�G�~��=�r�#X:�p�1OQ�K�
�����V4���?Ġ\�G��HOd�������+	(YTr��&�
������^����U��� ��9OB���C���Q�sd��EY�h#���e���b\@�O+*���� @�F���Γ�����.�>� �=1�B�'��YQ�fT�8����@\iX����8Rg�哙X�h���AN)a�`!*��^���'�ў�t 2��.W %��*�
n�9�e"O� �L��(�`H)N3MT���U8�tHq$�EzQ��W/.�<Q�a<D���S��O�Ь0K�ʘ`0i)D��p�#��pn>�:���D�d�G D�@�1����e ��7h��2�.>D�@8w嚟:b<z7�B� �%Q�#D�NW�f4Ip�� �
S��b	#D�HQ��������g��5	�m>4�������b)Q�J�4*N=1u푾.ȳ6�S�����S���!��\)j'Zh`MR?�
�h�;D���Ư4-��h��� ����-D����D�&��M܂o���QuA=D��ZE耖�b�;"�ڕw��)'O9D�P"���B(�!i	Y�Ql��)D�Y"f�1mZ4�÷o�H��A�g�0D��aɊ ����C9
(hᣲ"D�8�b�ʴfI���Cj��]rm�v�=D�p�$v0&<�2�Z�P56�3s�9D�H�2�;$�-XC�2��ʣf;D�T�n[T(<m2�f�2)�,i�9D��c�e�)���z��v�Xac%9D� ����
G�\i���ir 1��7D����E�<+I Qb���]h򔚵,8D�8����CB<u`CBI�Ь �8D��0W20^6X�p�D?}O�AP�8D��a�%"Bl�u��4k8VԸ`�7D� ��D1;8��٧l֟4�̱x�-4D��R�C<n��8�1bU�^� �qE4D�d�r�c44����W.�����&D�`� �Y,J����_����E�3�y�hՈce����T�k ~��dB��yBa�j���V!�#i�xM!Ɓ��y�M#��8P�^�+���y⃙�?�y��Q)\�P 'W��y��~b�B7��Eߖ��tn-�y��H�o�=�&��4�۔A��y��<���fY>|x\J4��
�y�m�/z��e4��}��,�0I2�yr	u���Q�F��8 &�ـ&^��y�%Y�$�A�D�5�FCB��y��sg�K���!>7Ь �� �y��מɜŉ�bj�����W�y���X�P��غA=�EX�����y��Ȋ0)�$�d�Ć`��ɑ a��yr�;��Ɇ@B�e��@�Ϭ�y�@�4rJ��g��+Jˤ��WCѕ�yh��L{�e0U�-N�bE���y"˟+4���x ٳ0E\@��  �yR�A�K b��J21<���yC1� ��T�
=xT��x�N9�y�L�5=���>{c�{��	#�y�G�"��׋�!RVPaRn�y<d�&A� �\>�����y�h@�~@*d!L���0I�CQ;�y`� >L�8TE�{�P4�͏��yRo6O+T�8gd�*:�rD1WȊ�y"��7,�^���R�D��� a��Py��؞i��1`m�?��*Pew�<9P揟lS�Hإ�I� .���Dm�<� �� Md����.afd��Tg�<���O[��A��B:lƼ�`���c�<i��΢U�ġ��c_�r�l8ᥖP�<�b�J�y��YS��[&
Jl:���O�<�FN�71b9 ��ϧ^I�Qa�!WF�<� �!��! ��)�N�m��C�"O>�zф���iSp���m�Nd�E"O�p��NS�uئ�Q��؜r�M��"OI@կ�gB�d�CF>�̘�"O���t�["�}���݉]� 1A�"O,�hU����!nO� p���i D�0��I�TȠ��VN��x�Ь#D����-H-֚厎�����y��e�*� �K�m]b�`�%�y"�A�u+B�I!��~< ��f�ʫ�y�L؉F$phf*S%r�îA�y�i
y���;�(��j�& cpH���ybJ�)�����Q"d[&����y2m�6yTD	F$I�MŎ�fgB��ybI3U��r +IE����D_�yb���V��5��L"A�fx�1K_��y2@R�=d=��E��IA���y���<.��I��G7b�)hq�(�y�J�S�0U�d 4�li°���y�ɚ�$�� �#)|[�D�.�y"��_���A$@�/��l2g���yÇO�%P��.�U���'�yr��f�u������\�e�5�y҉�(��Y������`K��5�y��}��i6��-*�(���J��y��/mo��@B�. 9�����y�� �q�0qkwa�'R,���'�yX�(�$���\�% ��y�O�(a�3u��
��qEA��y�H~���k��+�B �'��2�yB*�E���Zf��V��hӶIݩ�yBbB(3�r5HK�I�6��f�S�yB�=�I�˝1���qw�^��y�f���Lp�ܿX����Q+��y�
Єu�LY)���ָ b$�4�y�H�kLx��˅;|j�qy�!�yg�M� UI�Gԏq"2�P��y��R�|q�$*?r�V1�ЌF��y2m�8��-�����g<��(�y�aE8g��ѡ�NJ[�'�'�y�B�B����c�����-;~�@
�'/��	^&JYX�rv'��(w�i�	�'H��HGG^85��A�b	t}�`+	�'�����/�1ld�a��C�� <��@P\�0���%z�) $�����ȓ2e�Ib�I a�|u�"�G�yH�̇ȓ_����f��m�J
ыri�H�ȓ3|���aI�N�n�9PA��ܩ��:���jC�۶D��KTvi~��ȓH�����L�P��8*B&�?R]��t,��⇆�~��)O8rp��ڙ�cJ�7���s��5 ��q��CF�]����$HN��`.ͷ���ȓs����$�.7�h�p7��*
債�ȓV��`�(	�ఈA��E����ȓVĆ�H��I(o�X�a���,���i5�@�b!�	CR����{�����V�*�"a�K	Q\���#�.=��ȓIN|���*n��$�c���r��ȓ*�����F�9�f��a

P9*��ȓi���w̛/&�5�`���t:u�ȓiE���'�0(`�P�4͉7$2��ȓ+�4�R�/�z�ʠ�B�4���GgL�b��=Mc�cg��-3*�	��S�? q*AC��[T$P[3�O?s��48@"Oؙ�B�խjS���tLͽ���y�"O�kwLǑ%�R����@!t�m��"O��R"��++#|�@uK�#��P�"O�a3�9i�d�r͜$)�!F"O�-:B�@��i�1kU�e-��y "OT�R N	5�ZU��+Z�C�zhz"O�}�7/U�e�L�q���K�,�"O��!5�ލn��( �Jݨ�#�"Oa���v�r ��� =r�Qf"Oh՘aOBl��9yu/ڿfJ����"O��(�BQ�Z%|`�O�'"�	�3"O��r��	��r� sL�<�6�y"Ob$�pn֥�`�+)h�l�6"O���"$V�n
�Ĭ��g��d"O�Y�b�Q]i����*ϼ՛"O���m� ;=6��&K&F��`"O­(�o_�I�P9�A܇@���#�"OzB���)mr�uR��F�?FxH�"O�ͳ�L�;-"���'F�
)�]�"O�#�H�c].�;�P�t��"O�$�G�BL��АEJ�L� �c "O~�WK�5x6���܇8�V�I"O��
S�s�����*76/Rl��"O�d�"Q��,a��ƃ9M�9��"O)��0d Cc�V�Z�I��"Ox,�1#V[e麃)�y��Ѷ"O<Q{��D�bה1�a�O�Z�r��s"O��c�G�S������ņem�Q�"O T-E�89(��D�P�B����y2���mIcf��B��v�1�'��<!��B#m����fƒ��'a��A� ��|z�Cׯ�>��'��%p���%S���J�߂|�6ݸ�'~��1-Ñ� ��&��7֢���'<J��$��PD��e܈#s��;�'��XT UwSd���i�!4��E��' i���(�*��+#W<\��'��* Q�Q��I�B�K���B�'`��)��&\3zl��C�����j
�'f.��#Ǜ�}�`\J�P���eQ�'jdd��Y�(�$=3Di�|؉�'Ҏ���'�+}��9���F\���'^P�*��S�@"�4����6�49��'��y��ǔ<�1�*#x�FP!�'tȚ�	�c`0�#�� B*X��'C��a@٘!�5ARL]?K�(���'�ڝ�'��@昵 B�%F�̐#�'���pV�M�j�ɸ�ES�)�����'@��@$�D֐yhe)9���s�'��	���;�\��� ��0q�	�'�X�w�4f��8�GX� �FX�
�'�3��g��z�`M�?"�=BD"O��#w��.>��dj��K2Fx�+G"O��\~i�r�M9\$�H`�ZA�<a��eU�e3��)J.`�~�<�7�ߋ���Ǜq;Ls�'�s�<q�A]�.u�v��g��4�aXi�<)��ҐS�Z�hP���0�����n�<	��
k�<��,	h�0q�@c�v�<9�'װ*`:�A�
ɋ%ժ�I$�Y�<��k�:*æ�l��B��Q�Eh�<Y��=s0���GŅ]�l�(�is�<qw� zHD��b��M���8c�m�<� ~0�W�8��a:`-O�i04�"O�}0.>B�.1�T��m)f|Yp"O육u���0�
4��[�@"OH�ӳaJ2N���q�C*��4"OHl3$ͯtL��CP v�b�)�"O�tЖ�9y�����B��R��A"O�� �}0�pR�X�}�d��s"Ol<`֥D]b)�`��5.�@x�2"ONYuL$d���b�\_���"O���w�.YQ��aM�~'���#"O�3��(�d���#5/�T�s"O�p 0�9�"U5$�#Iz ��"Oȹ
1#ކiR P#S�����"O<0"�镍/�\�"U4Jx�5�#"O"!1J�7Q�Ԛ�$�d�-I�"O�����4D���̓a��z�"O4����'=n�){�#ȭU���"O~L�e)3��H���� bP��P"O�0�e�D�-^�ۥ�NuV�U�p"O�Y�1KU
	P�@��C�H�	jS"O�Lb��F�)=>�S@&[�bo�	�!"O$�;�k�9��h����,zD%1�"O��IaS"1*�e�e)��ҡ"O�Dy��
l�
�D�%B+�b"O��"e;H�����aD A�>���"O)��D3�VлՠԤh#(8"O\8���;�B�*3�"�	ض"O����	P�>�z#O��+�9�"O�H�H�)>���`�π�sB|"p"O�Y����B�:M�D���R�8�'qXPJ㊜�F/Pey7[��x�'g�92�J��7x`$��$�^6�@	�'�l���W�JU{M�$!FD�')�Xq��[�5�A� /ԋ&�$X��'ׂ�`�.i�`2ЮP�5�m
�'c��z�M2J]���b��, Jx�	�'o�P`S.T�c������^��'6L��J]_���ĥFAA�'.�,QG��:к���N<*��
�'���  D�UBL!�2O�����	�'����4�������&D�e歐�'~�(�G�R'}FL�f጖[��P
�'ˆ��+��`��+e҉_A��
�'䠪Fi�$y���U��P��Ir��)m��q��'���� S�4$���	f�ʝ���K("r
p�%�>15]�t�5�Sw�ĄK	wٹG��G*�R�eߊM���>ѧ"��i�B�^%2�:4h��@�8�2��d�3$&������P3b0t8u(]&k���J2�xb�:L��O����Ҵ�x��1�G�d��l2�T��S���I�S�O��1#�O��R�ZD!
�$2���5+�X�S�O�@�Y-עWb��=!�".�[��"Ca�Ԣ����qѰ�	+�.q1�O6��']NdɃ����8ld2��QhW��B�3��.��84"�z���d�G,�:��t�G%�I0�B����'<(�"}rsb[g�r�����-j:*�#͊ŦiC�Ln�S�OR��M�#:���$L�"h-��{0%�x��za��.V3�d��G��"@�,��f��?��'a�]������K'NUP�{��@�pа�e,S3��
�e3�����K*^Tq�?f<&uYD�P4���ʋ������r��-��2{�ŀ���]l��gę�h7�� 1���˭Xb��ԧȟ����a�:�j��*T�qP������?�@����I��0|:�l͢���C�v>ͱP/ 㦩Q�CR2��ē�� 0���.��p�cR�M�D\�p��(Or��6�0�)��Q6&lZ�*F2H�	�cO�,j� �V0�E���� l�y����=�Ĺ2��ͮ`,�ӗ�i��љ�����H?>MQ���	��D9!RW�]���3����$e�v��Ki}��F2,ꈬ��m)ksx�`'a��`l ˪OJ]'�"��^��8ЁFǕc/�P�׆[k�<ѣdh�c �S�%���E+�"OFm����?
N���댅-�jEi0"OR���ۃFM��pc��*z���"O�i�!���-�pY����Nz��"O���OPxr����H�[���r"OpL�#�NN�T�Awg
6Bϴ�a""O0�QBO�A���e�k��8w"O���ښd2<�6��&����%"O���f/܇ֺ-(6dL��~|!"O~-X��Gsa�"N���A"Ot���)O���b�K�&�"ON8y&���!���i����jA"OƄ����uf���! W��)Q"OԩZ���Q7�� .���"O��HSf��c�(�!O%�xM�q"O@�!F�Ǡb���pg��[D`z""Ox�{�fU�Y��Ae�G)Z\��"O�́N��4��3 8D�"O"�6eh�]�`k�!
\��F"O�u[�j�W�l�+#��/.N�"O��� ܡ/M���j��6�"�s"O�8��(~��Q�P��4|Z���"O(}�fAG���x�f�9v:�B"O��z�f&(2ih憚%h��A"O����ϵC��9��ъ5���ha"O��*"���^�zX�6D�6g�b5��"O`��6)S�@�⡍D!k#����"OЩɗ+�^�&Eb��n|���Y�<0m6O�q`�ԇ6w��d/|�<�T� 0R�u�0a=lqʜs�Mu�<�լ�2DdTb�C<�V�1P��n�<��[=DJ���1L٭<Y���'O�a&G�B�LxڥB�c���	�'?x�2��F�?V�Ѹ��X�p���0�'P�5iS�lY~�4"	#`��� �'��Q��[�r�,%�lC)RP�Y��'p�A�0�Y4f��46`�!\
�Dz�'�����k���
���ȖR�n$�	�'֦��!0T&(
D댿{\��j�'W��1`f@"VQ�`!���oC�']��蓇�-� i�<&�l 	�'!��'a�*��I´g�1rL�'.��%�EHh�Q��#�`]R�'�X�[�f��L|h*��K�1� 	�'K�U8�K�?>{R��OP��4:�'p0���N�	�~�
WKϦ����'/"E�Ջ�8�h����2/	�G�<�d㐮�6ȃ����D���R�<!�@�eE��(0���.��7&�T�<	G��H6`ac�05N	�C�k�<��M�Q���@a�M��M�ňc�<1��RRJX��F޶i���2�o�\�<�䥞�M��سböZs��٦#NV�<yt�2a(�+a@�.����)�S�<	�C�$�y�(/Ɖ��Pd�<yBh"T�A�kG�vTؙ2a$�b�<Q��
?�k��I�y� ��Z�<yT�D6�j�p2n��^���v�V�<qg��$K���ja�('�K"\�B��u1��Y0�4ڕ�	%aۂB�)� J9鐀��2' ��r)C61���"OX��O�?���{c��h�x��u"OZ�:4���"H�`s�C� ��xP "O^8�bKH�.u{�C[H�m3V"Oޜ"���8����&c�
r�H�w"OƉ��Ӎ%�.��!�k\���`"O��G�p��	�ņ�,NG����"O~D!g���]�Z9u�Y��TBF"OB��P'ϯVM�a��6���y�"ON��P�;5h�Z'�<-zH@�B"OJiS�#b  ���ɶ9�R��0"O�Ez�V7�*�H�#��4٤��E"Ox�y���3X���P�I�4N� �%"O�T�eЉ/!�A�A��:��y#�"O�@�奟�<=J�A��1F��8X"O���UJ�a���)�lۦ�{�"O����H6&�*c� ��±�c"O�j��,L[dq�)R���Z�"O����K�v1\�3ցY�-�"Q�"O>`�v��6v�J��B��;A�&,*`"O��I�ݪ$�"d���8J��}��"O ����H�qGF�g ��0"O֭t���K�d�%"���Ӕ"O~�C��ӻ�����YR̄U��"O*�xs�C5s���k�b�: ���"O��BU����C��;b�rU�G"O���b(ٻT�8���\:��H�"O��j%,�186B4��Q�nXi{"Oj!�T#H�Z���AE�ɕr���"O��r�D.��$��F:m�Ƀ�"O������ j�I�NS�pҍ�Q"O�mXP�Y�vVQi�,��AC��yB	_�km����o�1\��q(�ק�y��6�"�ՊQ�E{*bE���y���
���O	K�IJ%����y���bm�h�Q��x��1�)�3�y�g�%q�d[���@��	��lǜ�y2�*iZ����&;��K�ݛ�y�&�+af����(.`b���A��yR�N�o�����~ J���^�~��'�`${�%I������D�)�*}�	�'�&�yBG�&����mͨ9X	�'a��԰r�yZūíp�f���'vjtZ煟1h���*��T^0��+�'����"�/���r#.��Z:5��'^|00oF4���Z�[*U�j���'f�HfO?�8���xC�Հ�'P\TC��ǈlꔃ1�YZ�<9�'[���퀓pip��W�JN"��'���g�W9gt-R�A��q�h�
�'�y�)M�v��@��i+��
�'.����ȃ4��i,��uĽ��'�&y���{m(�����sv�Ո	�'��Y��ۇT�L���!�ƭ{	�';a���C<$���$F
&G�Y�	�'^�������%�hܱL&�"	�'(Hi���+?7PA:����7g��+�'��i�!�\�-��*Ф�=-��C�'FNT�A�U�n݂v섻nJ��'𚑺��,��;S X�Pv���'����*��5�Ϙ~7�H;�'��y񪑙D.4����c/�!���?�,(2�Ǩ'����m�S�!��U��|K�b?̀)��
X>@e!�� �yZF�N�3{���eK3|�2��"O[�%�5G���� �R���1b"O��z��V�y��X�zt[�"O�����;@�1��đ,
���"Ob5ud�>u�(��
Ê��B�"O���ĭњYUd4
�F�C�e�"O�0�&]�8sB@�ˆ5"�����"O�p�$ T�<��1V�Z���C�"O�Jt%_�_�X�u AI�]���i�ў"~n�=w�����
W6��}8�M�!��B��<yɮ�ׯE�>�z���ř�jB�	'l�t(�'��)��j Y�E>B��/=hR�hga݅g�Na��M�*B�	0f����u��*�X��d���"bB��UR.(��b؝%�&<�C*�FB��tz��ʇmL_����G�gL�C�ɾDo�aªS�
��;'���J��C�I"qn��	#a J��H`v W�(��C�	>�ƥ��D�D��� �Ɉ�fC��6ߤ�2�c�!v����e�1d�B䉸���!��O3!��p�"-5��B�I�Yk�1�,�z���q�m�"O�X�<�{�%�6if��v"O���M�>rs~��CD�/9��Y�"OT���5�f4j�!�MH@�ѕ"O�X�cB?�*8+�@P=a���"O��CE�O�GR6�i�.�Z$^UY�"O�e:���}��ۤ��4
(��"ON!���F>|ڸ]9c(I��H�"O��xg��0-oR�Âs��YV"Of푱�K-&�yhC�R4B�FL�'"O�ۗ�A"I��h���z����"O,4;g�E�6��s#�!|�"���"O �P2�+3M����ߺ ��1�R"O
�Qf͗t�TkЦ�uFM)�"O��j$��7� ��T�l2X<�v"O��VE�U��<H׮T�: �!�R"O��#��S?��Zwn֗@��Z�"O�����^+Z\ɴ,��c�X�R"O��[VAR�@e��r��ıI.�
�'���Ё�0N0�����@ 6"O.�1�W�T��$�wҰS�"O��3�J�
�ı!�`�0�R���"Oh�{�
�,p����a㰄�"OԼ�֦�
|�l�z�\�_ؾ�Q"OL�q�bY�+ڮ��A�[�hB�"OZ��c�,����'(����7"OPك�kD|�<-s�d� 
"O�� H"���6�c� ��"O�]ⵥL�q��-z�
]���U"O`(�'-ͫf,�	{'��V܄�#$"O�H"�R63bDSp�΍A֎�p"O ͩf"T�O�T"R'7I��q�"O2����/ZU"�s�L�;r�r�"O<�)&�"}"1[FF�,j��b"O,�1�ͺK+H����� aX,qW"Oޡ��	_/�T�e�!fE`�h�"O��Q���?&��!H�h����"O�H�Q��fo�e!ҦI�@�f�q�"O`l���T�8(����N�$ْD9$"O���g>rx�!
eNKD��:�"O88s�
p�N`G��+֩��"O�-���9.�8ql� �(��q"O>�#hЙ[���6�� K��:`"O� ���"!ZmTR��.�Hy�!"O0ۧM�b֌�3DF�
ڔ�b"O�8�6o�5s��R�E�b��[�"O>T����"�X�v%��$en�g*ON���O�"c�<4�ǚ1.BY������`�dЯ�%�P��y��9-��)����{N�,�cf%�ybɅ@Ő�9�f.ne��+6Ζ��y2炳]P����P3r(�^to�c}2�'�̝Y���yb�
�&��Ί/;k�DARLX�쐢r@�R���#` ���i��?]���M3�Al�i��ï'6h���K��ʠ�b�J=A�Xs���yyT 2�ꆺ,�$̫� s�	ۅB?��ͻc� ��˨o��qI XYfY9f�l�D�'����S�����ͦEх��; Px� 	�E3��Y��G���'xayB�.GFȨ'��Za�V��􉽘M�A�i7�'���O��41�L�	�L�6)6!���D2��G�Nj&�&�O����O���_º���?!�r��%{f�>0�*]Pw�)z�68�o�1nO���뜞BU9�dj�T���Be�b�'t�L�4oH�b�Lx#SD�?@*�ݠA �M�� ��jH�1M8����.a���7�ŹrƆ� "΢tE創�����#MD8`��LX�?p4�
�H�OymZ��HO�c�t���;M�(d 2�GIs��spK }��'��Ł��$�DIh!eCfA�m<���ߦ	�ٴ��D�-!�m���A����{Nݯ6&z�Ғ�õ"�Q���ɼT�MK`�ͷ��\{�J�(�p�%H$�t@��ד+St��ƌG�l섐k�*ʓ�j���LZ�;'�����[��\Cׇ�SF�%�bN�SGiҦkʮ@�6M�b�'�P(r��l�����<q`̈�r��i�l�!��83�n�l?A��?A���d�� X�BI��'�xꕩF>x����G~��ںq���9�"�/,���SE�P",���׀m���B $�g�iR�'���?"��l��d��4j�拌Z����rƊ?e��#��?!uL����r%M��R��k@`ŒR�<�� ����YX�8�[<H��h�#%Qe�':H�x�%K3Z� �z k/+�y[����r��"�j�m�A��(l!%p���z��&E�O %3��'��6M�`�q��oHƜ95��Yn�-�ҧ�#ʐ�'���'{�'��OlEғ��	5����En�2�р�Vf����rӂ�n�y≔<�����R�O����!�9��iv�'��)�)��AS5�'��'���Ƭ����o��pC�ۚO��5�#|��kE!��Pq����H%p��O2���Z%R��)��������~�>�t+��42�UIahĈt9B�H�
��q��+S�3�Z�#�I���I�! W,�̻<�܌�@�;#�:$��ݘzX�S�m�ޑ�'���H�S�矘�I��2QFԌf��`Ug��x�d�{��/�0=�{��Fc�,��74� �3�LQ���ɳ�M��i��'��O��I.7 Z���/����L�H��:�/
�D��1���?����?������O��� +!n4�юǘ+z�,(�oA�L���	���s�&�&D��� �jO�4i���Z�8�!N�y;A�5K�a�E��Q�!� Q�h����ڦ�p�,oӠ�9��|��0���/l�R<�Z�nmh�a�;���3���'�4�!z���jSa�$���'��y2�x�FD8[��jlD�m�|����]oJ�O��m��M�M>���?�]/�� �  ��       �     �+  (8  D  �M  lX  �b  `m  ;v  z�  \�  ��  I�  ��  �  /�  r�  ��  �  6�  ��  
�  h�  ��  ��  .�  p�  ��   �  R � � � # g% �, �2 29 P?  Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�� |d��"O
`�(�;���8���-0��1%"Oj4��ND^[��"3/9�0|H�"OB���H��*�ʞRy=a"O�味V�!X��!&F�:J�$���"O,��a
���C�Ą�M�"O,$3%o�-���p���+Ն�:1"O��ݢ1����`���y14]2��i�<�6��{_���c�H�`�fX�$Kn�<��A̼VI�xR[�)�Ć�pඤ�ȓA5��('nߡ4�� �)˩%� ���,��r�؊b#`T�eT09���ȓ!�b��g��}�8�F��-? �ȓ
K|m�ș�VṔ���2�%�ȓ"R�X�j�4JN�1�˘X�i����̹	_�jZ��1!g��zܶ��ȓgil,*�J�
j�Ne��i�J%b���f	�(U��:���G��$Y^م�~r�� S�%T"���k\�jx�ȓ|4�1�îJb��@ӵ�ݩn�V��/[`�"�v4�R�!ʎ<��M�ȓ`:��z�ؚh�J�Z��$HY:	��H��p�m�C1��!��B:��0��EnjZA V;9����J[
2���	��4'J�EA�IVW&��~�(aZ��ӹ�>� o�Y�|�ȓ�f�A�
Ο7�H��M�$�����mޠP����/���ANXo*�ȓTv�����{ ��-7�*h��I��sB�8�8���3����ȓNe*M�悡;������X�o��!�ȓ'lj�#F�m�+R&;�|��2)n�C��0S4���T:
b���:�0!��e֊��)��ͷV��,�ȓ0�&�8#���� ع�L�����;�P�AFd���,w�6d��r�EQ�( �gVlɦ�M,H��,DP���|�I	$G#\���ȓ"�)���E�B	yt&B�^�LɅ��wyr*\(u�@ UV$ED02�-Ə�M���sӀŃ��L%'�r|�f��52���5"O���BO�876A�%x�`J&"O��@��~�nW�8\0H�teE�<A/�6r^�=��OA1 D�k#AX�<�A6I�P�j��B�0�SJ]�<�t"�>{D$1�dȫK���b���bh<����d�n4�s�C6P�NT�T�E��y"�')��m�):T$X��䔗:,.mi��${��E��$�@�Xe��_�F�:#�_�yB"�	s�9�1䗿E����A���y�	Ǌ"�
!�حNn:tbqa��yr��ZCpܪ��Csld���W���=!�yb%�.��m����=1���*��yb�խD?fd	$HZ���h�E�a�\QEy��9O6y�D� CqX8!��A=	z�!#"O4l���	�/��]����n��DI�"O@��B^XX��V�m(=h��$�yҹi)�c���SJ�ODIi���.h�xsQ��E��B��~B�@���!���D4a��������(�xźgȒ�i�2I��cD,cĸiQ"Oиc`�A�*HV!���A7VԌ	��|��'K��*ͦ���"����� �m��	�վ��1EʓH�̒Q:O���d�w��� �D��(4z1ڴM��IZ8��$��Q&�,��P�$F-@�h(��j,D��Q�nE 7���F!Q�	�Z<���<�'/�{r� "�li4��*:��$�����p<aM<灵��Y2��
�d ըP[KF� �hO�S4U���a���?��;���P�C�;��$�RI�&"i�<�g��E��C�I!f���"��5I�d�ɋ `���hOQ>��I�}L�� Q���ը�O�B�I�E��+��I3|�b�nJ�1�P����p?����<8j�y�Hύp���Ɏg�<Q��KX�� 4/�$H��-�4.�a�<9��\�\�� S	�
t���`�Z�<qg��Z�����-<�@��Sܓ��=��$�FHUPơ�'Fa4-r��N��4oZ~)�f�΀.ל�rመ�wt��Ө����>��OH��<��L��Z<Pv�@���i���	
�a�m ���0	�xⶃaA!�dV=�=zv�ܼ(\a`�ۄ
,�	��HOQ>�PQ@Ъ��83Ff���*��$�IQ���'DŚagjP�a��:5���e��-�ȓC9�=a��ˈ.~��j�/��l�& ��Q9�-���
���Ĕ�T�l�ȓb�zT U�R�h�>X��O!\P��@���@����t��l`)ϨV߼����6�H�'t�i�#L�(���I�4C�^��.��S�O6�=a���6�`������?O��=���OyBK
/���@��$��t���O�x�3�'��v�i��x���<&æ�B�O'<����en�����؟��.�S��mܲ1�Y��悽9&�H#@��,+���Л#Ы�,֛F��"7�J;�!�آ@Ӕa�q��@L�K��P�!�d�Ȁ�[p�[�X�4����B��I��0?Q���rA�u�u`K�L��ܣ�m�h����'
j �S��}
 ���ć<sʞQH�'{�m��ꁨ%�v@i�m�Z,b��$�>I����O��y���%:d e�+^�Л�'�x���j���I��ᖒQ�؉�'Ol��T��+{.�q��ӊb���`�	ş�F�4TJ� s)�+Ԟh�P��?�y2�'��#�@?X����G�n�x�O��=E�'̯/r�}I@�Y�I��jց�9tq�'Aa|�%M#]��R��+>��#a*N����'6�xQ ��H��I1�#ʟ�t(� D�����Q,pv
����cW(D� (V�Z0���ʖ�EK�(%��ȟ��	��1���dlz-p�"O�)��N!A��ѫGI^�L��"O��g
�2P���	"b΁j=��"OF܀����/o�	Fgl���w�IU>�Ƌϩd�B�ҕe�.[܍h&�.D����A �lX�h�,u��ժ%K6��0<�Ō��~��j�Z49[r�^Y�'ga��.�"dh5�޶@:�o;�y2dD#2'X�p�`�����Y$*N=��<i� 3�	
V	4h��Ǝ�Afp� c�h5(C�I \/��q�l�FV�(ʣ*K�MC��6�m 0BֳM]�ר�R������IgM���x]p��ϖm�U�/D��D/U��t�g��9�� �d-ړ�0|�W��._�������<UZ�3dl^�<ٲ��8�1�s��3
�z� �&�؟hE{�O�f�ȨTF��h!�J�j�t!��+��p<� ,��@[�t*̕J���-$����5"O@��*�^f�2vB¨;70x�3"ON�X cZ��11�@$*����CH<1$U�xc"�b�c�n���Wb�<5�KP�L|ab����4}�!Q^�<1�f׀�>��'��y����7�Yx����R�֕	����U�j���ε�y���cmrl��Ε^:"Y�J����j�h��$�m�dǂ�?�9�u�X)d�a��O��H-�� G��V��c�`�;4�i�O,����Y��	"�3tR�`��z]�t�4O�̓"z��eꝆ0鑓d�<*�O����D��),m;g,5O>p���>������'��RK�-��Z!;�-i�'}΁�dF3s�-��� 4���O^�q��c��g�I'�|͘�@�&lD5ۀ�H������O��b�]8��dr�oՈWk`��1��2�MS��;�e�̬`�nBZ�"jS���������=���L|��!��C�
Kā��k�<� ��E��;�m���<cA)�~�'Nў�WYpL(���vI]����t�Ș��ybZ`�� Y�hQx��%CB��p�Of�=���N�����s�H�2lt��B s�<�uսmE{��H)5�U83F�k�<�w&M���I	p%h �c�<�#K_;T���Pf�ӳY�2(�q+�a�<qq��z| tY��A�����Cv�<I�+B	T����
B!<��Ѓӈw�<� 	+]�ԍ!Ӥ͝&�3eJ�t�<�BKU�o��� �n�gxU!�u�<��Ph	,��5͔�&��#�NW�<� �(��}����
<�L0�� �T�<ie�Z �<���*׾�0��\F�<ip�Y�t���HDm�iW.�DH�A�<)k��dR��
rΠ��E�z�<	r�X���U�B�p�@pC�x�<aw!�-��V> R���e�^�<����6sh�G��T�Â^�<eaM&l���@0!ڂp%T�3rn^\�<��芟_���pl�}�0;�l�Z�<�Ǩ.�(��`������wBN�<!�ə�lVU� jݺR�j�bRF�t�<���ʔq��Z��5o�Ȥ�קp�<	���x��E���F��HF�<��i�ny���Ei#�z��H�y�e�/LB���8/�$�S��yB#�>@��`c0�[XR���:�ybU87���@5i   ��Ӿ�y���'`�mn|fy1��%�yB U���`��L��S!�C��PyB�+I�F��a�W�\�XXu��U�<�d��E�I�H�%� ��nCF�<�����_����E<Z�.�R��G�<)CJU.F?b����:i�TT���@�<��B�1�4̹%ڷ5�<Ѹ�WV�<уB� cG�X�	G��C#Z[�<�#'��E�
L��[�ab|��C�[A�<	�Q�YN��QA�OA֬�!զ
{�<�GǍ�U�2PK?e*A�#��x�<�A"ޅi6�ύ�h",(��I�<��^�cl�b �Z(O��C1��`�<97b�)p%�aA%��QM�\��]�<-����tC��@�x�VER�A����ȓ4{��hؒ=9���拺|2|��S�? �	W,��|�u�fBu�h��"O �Їd�K�8�),;Y����"O�d�B`��
��-�q���T���R@"Oi)a�E�F�FM�k��h}ҹx"O`貦�҄Z����Ԫ��MuBLRA�'5�_��������	ҟ<�������6�YS�C�xu�QZF���s6��	ڟ$�Iʟ��	��������ß���4nv��X%IU#s�@���
~���I�������I�d�I��<��� �ɭ]u�)Q5)ї���Źc�j���ҟl�	ٟ���֟��ȟd���X�	��L@4��2=#�DRǫ��f����IğL���d�	؟���L��某�I�~��@܅+ߪ��4b�.,gx��I�L�I����I�����ԟ���ן`��-KC2���\<Y�b�&L�2��Iɟ����8�I���I런�Iҟx���J�����t����FH�6.��l���'���'���'���'��'���'�8�Z8D�W��9�D8�Ǎ�+bkb�',�'���'j��'�2�'`�ǐ.^��99������dʓ!xr�'(��'G��'$R�'���'��m&H��T�F^�!Pb *J;R�'��'�R�'�R�'P��'U��k�T��Um0���Sw�����'���'���'*��'B�'9�+��n�`��C��z�4T�!cߔn���'Fr�'7��'9R�'66M�O>��ߣ6�b=�1D�$:�.}2&^,%�88�'��Q�b>�S?�&�?x�>!�%��<�ҙ
���.
#��O�nΟ�$�泟8l��;�6颲������q$E�+�n�^����e���8��Т�V��4��A�~R���)~ADY+gg�C�M��NT��?�.O��}j���a��	H���4�R)�6����'�񟒬nz�M�����䨈��� 3� EC����?�ش�yBV����	2Bƒ?��d�E���0D�Ѥ{�N��S�:��+c�U�7k)2�=�'�?��@�GM�%X��N�f��Aʇ�<q,O8�ON}lږ�pb�d�AD_(��"CG�n `�S�v�i�Iȟ�mZ�<��O�-¢�>�n;�X�]�ֹ3w���2v��
~5HW�)�S��%hg�	���pȆ"+��5G%X��Ӳ��IyBP���)��<ٔg[�G���Ya1�@pR���<9�i����O�Dl�i��|� �(�>K�Oҗ<GT��m�Z?a��Mc��^G�t�7�G_~r爞R*�󡁐:��-ˑ[�FF��$Fw��i>�'H�OaL���N�T���%ްF'�r�OJ�l�x�c�4�SV���Xh$d֐��.L�Ղ4�*O4�Dd� �W���?����Y�`�`ᚌa<��ڄ鑒E�����B.%��O��,R�ƍ??xi��m&ړJi|%K�@��,��FC]�>��l����d�<�L>�g�iM~���'Pp P��G�@�*��úZ)|�'O�6��O��O��O>�D`���L$1��U�BF��}b,��k�+A��h��̀,m󄃲����.F%2��EX�O���̑�\c�d�@0Ӻ#E���i��R�����'�BT�\�����]Y���$VQ@x��̙t�H�{ ��IͦQZw�:?1��iN�'��ۄ�+&�v$�u��MJ�|;�=O���M��i���=Bp$��'J�\;F�MN.�<�ԥCoF��T��*C�,Y�GH�;]H�:�x��uy��'~ʝBb.�C� 0z�E�'CO�(��'��'f 6�I�oL1O�ʧOR�%!D)I	Z�t�+�l�E�N��'~˓�?�ڴ�y�����OQ��j�J��3�xy�e����3ƅI��q0aW+���蟈Ta���/O����?i�Ĺڢ哄A\(Bk,�cc�1�?����?����?�'.H:���hyB�c��	��ųR�1��	ư�
���Ƞ[��D�O�yo�C�i>��O��nZ"����@2��r�+�2	�۴S�F�w���'�2K�#l�@�`F�J=l剗Y촵 ���vH���/�6*�	Ky��'���'��'��Y>y�AЂs5��Q��P?~�ܘ:�ԍ�Ms�?�����?�ȟB�'��w�D�!�I1�µ�C⑋2��Շr���m�'�?i�O�쟮�	�A;65�%;O�Y�jJ�_�䕳"�E�g��c 4O������10wP�p�5��<q���?�v�3����IϤ:����NA �?����?��������4�2?��	�.Ã�y��`�L3b
���H>	��b�	6�M���i8:���>饤��/]�����������f��<��=��@�� 
�^n"�.O��i�
3�`�!,�O��EF5"B섐a��	���)5��O����O"��O<�d$���H�M���wl�XQS�V>$N���EّwT�����'w��I��y"���4�|�^� :�*M<Us��sf��9F�P㟈�4)x���|� �������Oh�3���9a���J�08���
� Э
�~s�O��?���?q���?���K*�Ipס/�R�2AcY:@t��.O�0o���������IV�s�D{�I�n�a�bJ1*�Xh$"Ɇ���٦�۴A�R��t�O���-��F+11G놌+c�<ڳ�8n�L0�c���w��94B�� ����EL��&��'ئ��DGlؐ1�bd
cOFu�@�'B��'
���DP���40�(P�	��Ht+��fm��/N4;	1̓'ߛF���m}��yӬ�lڂ�M[Taݙi�x�s�BX��53�-�r!t���N~��[,mFjt�qM���O�.�8� �t��ͣ<X؂��=��A�=O����O"���O~���O��?�Mʨ{��]{�F
0dah2�z������,��4Lt@�'�7 �$/r�aã�@D4ࡀU(�� U@���v}�c��poz>eԳt�Aԓ�P�E$W�av�ba��e{d�z���:'�.P	Ý�#$f�G{��'��I՟��3�߭0�����Ѽgm��T*u��&���4 z���<9���zCEX?So
J�E�+�*���"d~2��<I���M��'��Os��n΁���6� `���e�S�:��\�0�űz��I�O��ɒ�`�X-ؒ ,�D�b\r��%
�>"\�ł�\����?(O1���4�MBa�&w����CÔ%�N)遈M09Fx�'�,7��O�O��O*6̀�?h�="D��ީa0F/D�X�mZ��� �hއ4�����{D��+b�s�c(?ɦD�#<_��R��6�ʡQ�Kc̓�?)O�}z��PR0�Qpi�8�x@�"��F	�$��'.�T��$�z����P�	���Z.����@��;r ,�������O��T�'�zЙ�lǝ�y�hʬB��W	��a6l('�C)�y���s���4��rCў���|  $	]QA��+�!ы�fk�t�'��'4�7b1O(����ل\�	@J|l
t���O��O�Օ'�iG��>�K����M=f2���Z�<�#>|��NN�Q���']�T�x��]"�'ʨaH��-�2�G�a1�!��'���'4��'A�>	�I�\"(��"V2�k7�i�!`T���S޴$����dG����?�;=�D,� �8�luy��7[0Tl�Z$��|Ӭ�o#y����3�������g~rAXb�H�H�:Yr��+�@q '-D��'��	���֟�����l��4:A`�ȳkЅOWB8A�N�W�޼�'>�7�
|q�	ɟX$?����F�n�0���RX�J�`���Ts�O�InZ��M;�'��O����O�ԅ1�$_[���q���6v䐠aY�=���e_�lؑ���t'\p�W�fy��'��I�r�*�`�oǾZY���F�6�^}��ԟ��	՟�I��M�(O�Do��6�R睒&��eI��̑@ͦ��7��n=�����MJ>ͧ*	�	��M���iS�6��
so�E��W�/��b� [?<�t�Q4�SH��h�k�6v	@�q��� ��	�2���(���E�)��f�W�l ���:O��$�O����O��d�Of�?�̔�WC��� �}]�ӧ�����	H�4Kq�,
(O�pnZK�I4�K��Z�4���U�]�ST�l���d����`�4���P#mD̓�?�!@_�b;z�k NT&O�HLL� E�0����N��Jd�O>�(O����O����O\�����~Kp�2�[_y`ȑ��O4���<� �i��Tk��'�r�'8�Ӱ ��m�d�Ғ(��X�'"�@� �@9����M��i�6�'�	���Q�	G&=��J$П	�j����^��%�W˄,��˓����8��
L>��*W%yX�R�ݦUP���H3�?����?���?�|b,O��o.Y: �8�.��>]������n������O��lʟ ����
�>AA�i��Px1��Y��i�,����!�i�z}lZ=`�̬�'j�4�ɵ�:�zc�?J��'C~5�7`D1, �DH-6��'�	��L�	ߟ��	ʟ��IB���G�bi��J7�$��  W�t6�^��I��0Χ&%��ş������m^r>|�h�$T�nڠ<��暧~�FaӨ-m7��4���i�R)x�d��k��d�/d1�tڶ!�i��]�b����I�=5\� 7k�$1��OX��?i�~K���T�B��-Y&`�4,�������?y���?�(O�=m�qך<��ğ��I4N�V4�4d�*L���Q��E/b0�U�?��Z�4��4uӛ&g�OZ�[�:� H3sL��@�ȩ��?���w0�EHn�8���t@E�U9r�n�$D;l�MrM+ ��hW��&���d�OH���O��$-�'�?�d"s�dώ\�f���dE�B�49���3��$Q�i�M#��w8�D����c7��
�2Y�dK�'N�7�HƦ1JڴT-��$��<��GI\t�R�'J�]�6�l|�Y2�L��J��"���䓆���O&�d�O����O���XM�����>u.�x�@�1����F��y�'����'��T�E��#=5L��EHE�e�`����>��i$86��ߟxD�dBݧLZiɰG#k`M��	�#	�D����	�'��r@�TZ ��'!B\�4�&� [�D"�9y� A2` ��h�	��4�I��4r��WyBt���b0�p���O�@x�� �H|z@kBA�OplI�i>��OblZ'�M�&�i��4��; Y�@�GGU9#{h�)� _�}�&�K�'DƲX�ɣveB7 3�I�?U�_c֒��p/P��Ej7��*�,@��'&�[�`����ҕ�s��+$@�c#P�@h�ڥ�$���5�)?���i�BP����]����ƶv�P��$��<�-O�7��Ȧ����8�
��g���	*} F��n��t?�X�l��{m|�yt��;�Lj�@�u����W�L�I�y֑�х+>cJ����An�IY�ɷ�M/�ּ�<�/��dK"i� {��H�c��Kn�� B���+O|�{�,�	^�S�?!�!��f��%"fb��fqxe2��)�뛜ad���CĖ";�L��K>QW"S/��u��\�*��m�����Op�S�g~2�n�d\+q �8�� a�2��ܡBm��.�I�Mc����|��M3hqݲ���·�c��ԉ������'�(�s��yb�'�%��D�/��5��O� � yBbZ�iw�X�I��ua�T���d�O���h�8�jA(� @��}���O	V�$�R������3�IG��H���w9�0Q%h@�3�<6���<Ap���O6�a�(��j�'�?��I�u� �͓-�(�J��ȳL�h܃C�ԊX�|�	�*!s�J�(:,��M>a.O��O�h�.�shmjc+�=��$e�O��$�O<�D�<��i�69��Q�l�	�e�F��7/ڵR���ƠZ��f�	x�Ʌ���]�۴[��T�ࡰm�)x*��
��9�1�Hv� �g�Ϫ`�����vI�Ӻ3\w�� 3�Ή�@���d�5EbF���D<�^��@@�)I�����O�D�O6��-�'�?yǌ�9��@;�G(|`ȻË@��?�"�i���2�Q�� ݴ�?yL>ͻ%<��b��|E�ԁ�;�N�̓\k�Ex�FqlZ�:��ǂ�y�gجH�8�V�[;9Op0�w ğ?q��!��D6d�q�Ϭl�j�nʓ�?����?����?)�K�8l C����J-n�R��.O(m=uYf�����IM�s�������Upa��
S�Jia��	������ܴ!O���t�Ou��@�p�M�1	ԆOR�)�Ć�_��HDBY(��IR�"�Q�g�`H&���'�^\���M
^��sCDGb�E�'`��'{R��R�HݴB��R�=�N%�7��o���a � �R�ϓۛ��$�l}R-jӂ�n��M;!cZ�8��!i�0���
��Y�2y����<A��OL�u� �<��*Od����;�L8m@08w�< A��BeF�<���?���?!��?!��t��!7g��`F�y4�[W�T���]rc�i���'�n6��v��d�O� l���'�ȑRg��/%n~e��:I�f0����O
�pV�Ơ`�\�iQ����?Ox�d9�v�1�,S2�Z��@(�������H�:����8�ľ<9���?q��?	��&�ҥ� ��1
J��E���?�����$æ�Q��ny��'��e��Q��tAli�I�'sl�c��I9�M��iD��0�I�`�SD[>ղ�����OFJ��ᡇ97;����ꏈ���q��=&|�#O>!��T�jeA8A,��/1,MIT*9�?����?����?�|�(OZ�l%CX���ŷي�#� �9v�q{ FEzy�y��㟔#�O8m }�R��	
b	J0�Ò%؊u�ݴ^뛶@IJ����'�b�kbh]��J !g��!���Z�S����yҶ1۰H��Wj��a8Oʓ�?	���?!���?Y������
X0'�#r�p5'�$h�nZ+
��I؟��Iq�s������;#C	�D��=+�_?7���Hw��c��"sӸ9�	n}�O��d�O���P�l��y2,+S6��+����H��0$�'�5Y��ԃ{���Kq�|�S�����h���Q�y���D�@ب��$���@��ßT�IYy�/t�nE�=O����O��X��]�4�F��l> Q2��+�ɴ��������4=�RY���Y(�A��!�����X��5B�$y&ʌ���]�N~ ʓ ��]���fT*�TD�F� ���K�eѲ�S��?Q���?a���^����'�����ȋO)�-�L,��M�F�'�*6-0![��O4�d:�4����$7��A*�����1���L��馅��4H�f��}.��'���A�l$�z"��[mH���C�@͞�Ʌ	�*X�`�|�S��	��0�	ɟ���Ɵ�C�&D;'��'I՘%\,#���hy��u�$��ضqD�$�O��S�?���O~${�eϱHN��(�~8B� �<9��i)(6C�,'>Y���?%(e%�U�m�q��"2����)W�yQ�M[�<1#/К+���F�W�i�O`AS+O��B�Kçk�	���J
y�Bi��Ġ<���?)��|�*Ov�mZ-�� ��"]�Z����N#�B�E ���,�M����>y�i�p6-�OD�d@�l�kԆ����86`�8�$HT��D�O���#�XRY�t��̴<��Kk��7)�z����ȃj4��S%ǛqQ��O���O(��O��D �S�a5jЉp
J@*��K�`��ܟP��;�MsuɛM~"��ܓO �����*y��=dꊙ��$럨�'l�7�Ħ=���(�n��ƥr���I�W1\�Q���">X�����q�����g-�b�UCy��'��I���ϟ`��95{���Eؑ2d��S�͝�W/��I��M#(O��o35r�$�S�����[��C�n��)�\<h���"R��y"�'��F��։dӖ�o��ħ���$�+@�E��C��h��t��xL� ���U
<P�q+O��)W"M ��4� ���.�,Q�chT�M�^��v��Z�t��O����O���	�<���i	5�#e@�G�IBw��&TT��j�;?P�I��M����>	��i	 ��� �N� �eJ�	`:��Uf{ӈ�ndT��RLc�$�I�S�^�p�V�+B&(�'�@�����X�V(:EM�|ʲ���'��	ԟ0��埸�	�X��`��@S�Kw��2��=%���-e%�7��Z����Od� �9O��oz�A�E�I&jR�쓵��1C�HM���M�!�i�b���>ͧ���'E��D���I�<!�+�j�� �%�&��Lұ�<��ɘ�;��40�Τ�����O��D�4r����B&M�`�FrU*\�P\�d�OZ���OB����2�yR�'"b�.$A�X÷FK7rAB�N�p��|b�>Ƕi+6ͅ�h�'�J,;�,Q�x�m��E~Xة�'�r��+�at����?-+1$� vx��� Qt�a��q��(�!� �I����Iٟ���Q�O����t��h)�b�I��T�e)�/��g��h�@��� ڴ���yWD@�r�V�Y�S7h��dJ)�yR�a�^�oZ��M���:2*�̓�?pC̮@w&�b��O�? ��؅J8@�\؃�
���:��%�d�<i��?A���?���?��F�F #Ӣ��Rf"��R��f�	��M�aZ�<)���?QI~Γ,|r�N�'y<����.G_섚DQ� �ش'NvU�ڴ	�O����O/���a�!�X��ȒVh�4j2�%`���XbZ���K֔G�*	JdIz�Ty§�3�&p�R)�F紝
�oF-v:����������fy�q����>Ol����^?dL���gH>?���6?OdTn�C�|��ɸ�M�G�i�Z6M%Z��Ip��vJ��/A79Lr��$͚7X���Ot�&�-A��Y���<I�'y�kLą),�M�S���fHh�=f=���O�����i?���A�'8�9�&�5�*c����4sLE�'U�6��O�˓@�Vq�X��S�W!/��g�</O�6�i�@!�'L��kO��yr�'�2�`��(�>��I�Gx	�Gث7�"� �h��ў�Qy"�'��	�jN�L�I�q�����'��'�6mӠ%1O:�I��B�{t�
�x`�u/�.��񣅓�8�/O���|Ӏ�|�S�?Y;��M/}�6eI���V��E���E�c��  j�������b��)'B�[L>Q�ݾs��I�܌I���1u�߾���O$�S�g~2Jr�D�e�]
a�H@hC���||X�nF�a���	�M����~�i�V%0!��KH� a�/�8��Hu�Z�̄,&<#f5O����u���F�³{_�	�y���C�_,��dIʼYjc����|y��S�1޲h��%A�<�#��FDa��45���<�����'q回w��`��Z�B�3�C�t�d@T��O�7�j�h��R���?���®C��s��<�� D�Ä����8Ee,ΓR��S�X<�[L>+O�I�O��6iC�k��У���/r�"4���O��$�O��D�<��iI�]���'S��'��`�w%5n��`�bM�0�e�'V�'�@�R��"pӈ��IH}�U%U��p`��[�����y��'g�A��uҀ���\�(��9*~Y#��
�\p�X8i��̓G��/l1L�
�ן������	�TE��'���S�B��')�Z!lV3Kr�i��'�6-L�R-��6��V�4��z��H�]Q����6�)*&4O
HmZ5�M�u�i�Pp���Ճ�y��'�n$�7�ףuX!��(ZK&�����L~���a3��'|���������Iן��	? �����Ǚ��9����oζ�'N�6��%��˓�?1���M5���@#K��X3���}$�yٛ��l�R���E���?���6����M��W�h��@�<8Y�Ĉ��W';[��'���b.*J��p[ϟ��T5�y�&ް)M.���߶c*Xs%��y�Cνf������U���A�Ü��'Mj|���x�D��#��VMK!"�2F�a7 7R�4�Pwn�m���9%��w5��6G=��{��� pfyY�CP ����DУ},fk�ᛒ?/,u�	�,!X�% H��z5� ���q���qC�]�
ƨ$kq*T&ƦHpt���t�KD,*ݴ�ۃkX�}ِlZ�41L	�@�9gdXX'@�m��t��O���O\�O���O<���G�O��2�T��1��J
��a�vmMզM�I|�	�����ԟdB1�
/�M3.��̡g,�!A��9�o�L�x��o�Ǧ��	u�䟄�I�x�v��	Ɵ�	�C�|�zҏV�A�4�B�f`"�ߴ�?���?��8���X���'��4�I�f]L|����w��q��[���O��D�O.����O����O��d�?)2��=wj`��B�p���}Ӡ���Or�Y�٦�q�����Ꟛ��';
tHG-��]�����W\cR5y�4�?���C8��j��?����?�M~����'Jp\���,L�,u(��c4\��07@X�r�	P�dQ�L@q�	b ��BӲw�ƥ�� ē9G��-pX��s�/ B|�4 ��T�!�J�;��tA��;��	B��d	��	O�|11�E�rA���N��HP�C������V���Ip�?A
y����){��(��Y;I�CQ%��$!�ǋ�U!�e���5
iT��S��'g����U�^1aF �G��Lg)*�b)ܶy16�&&%�E�R(��d�O*���O,-�;�?������E���[Q�-t����C��Hb���S��5"#���\�J}0w���"�@��.R-W�]�t-N�DW�;&`�}���bӆ��}����W�S�cr������4�&����l��<JX�I�'ڭĨ-�� ]4���ަ���4��'�hc?�j��/��t��0 �ֽ3�%�O��OL�"�;R�$}�Q���2�9��dަ)��Py�j�
8E�6�O�� ��H-�o4np�C$�Y����O�
��Ov�$q>Ur�+��'�����onΝ�/^	+,�"U�ԫ% �*�	>/�0-����ݲ\�^�)�OY	i2�8d�E'Ej\At� aFE��dʦy���cCK	|ӎ�c�aZ�&z�O��c��'��'x�d���M��u�=?���
�'�`�����#R�hQ@I�7Ă䰊��9��|�i\	�`�1B_�|��.*�!��|R�V��7-�OL�$�|���=�?9vd˴n{�@��nϖG��ja͙�?���q�.�pw���!��-X�B�>�O,�
#r�������!2� ��
��	���' �p��4u(IZ�b"�D��t�DiS"of���E䂀H#j�O�L�U�'���d���H�)H� URdGZδ)a����'�2�',�M���H�uX�ų��͉a{���1���c�J�9�����8~J1HA��6�M����?���)UR�¡*�?���?�Ӽ� ��K�@�&9����&�o�@�%h�'pw&�# �B���u��(g��c>�O|}g�������6�
�j��<�AjߌD�(qk�hU�mxXДȎᠱ ��1��+܄Z�]�fd@�+H9+q�G�*�@I>1�ٟ�>�Oڄ�rO��I��Mi���xt=a"O��r.T�Jx��c��q��h��ᓜ{��h��ܴDn�ٰ�m[s|Hq��U�I�IƟ��ß�`^w�2�''��" ��)����`�����f��u	�h�̚^�H ���f�!��I�4�N��m�1s;RHБK�|ϔ�S�o�
7���r�e��=ˮ�P˓j|��6@Y��.-���3	j!��N��d�	��?�0��#��+�p"g@''��D�ȓE��(�E��B_�1Ð	�"Y<LY�<9g�D�2��mZ�ɘ[�lቀ�Ch녭� 3���	ڟ0r�.�� ���|�r���<'� ð錏c�q"7#V$:�y��;O�0؅���9I�:��ף_��y��D+)�xB/�.�?�G�x���h/%�$mW�aCZ��@ F��yBoW�`Дq�\(V�r87a�%�x��h�H��f��\� 6�O��r��D�s�&�n�˟���a�GM$_.��ʟE�84���
'C<Z�2�'����O�T&�p����
����i�|�"C�(��ؘgk!"�p+G��@�$t >��U��64����ц)ӊ�(g���W�J���O�����["�M��#�p�2 �H���$��O�b��?��" W5a�,��bgF1c�H�Ѥ#D����E�:���i$��!D��l��  O�(Fz2�B���xzS��Eq�|A�懵w�(6��O��$�O�!a�7o0����O"���O���I1THyN��E���y2i�� �2��u狏a���+�_�#���{��>����ɢw�$���	)0�=��F߶�V���!F5�V4��i��X���UV��1V>M;`��?l��<��0G
ʦgx�$b�ʎ�I���%�8B�Jn�b>�O��W̄��XyA"��4#�r9��"Oָ�
¾t�E�EQ�W�V ����p��4��O��	�*GQ&"�X��(��H�M0z����2�O��$�O���Ϻ���?I�O�6��1ə^��aGE7h\Z0�/sx��F'���R�'4�,�#J�
�n���ᏼp|�󦠏�4��ax���|�h��#Xy��A��5{�]��{RJ�go0�	+R�B䈥1CB��OѮ�S���?��@AM�MB���4W�����K�<e�ܳ;pf�U LP2z�J��J̓/͛��|�C�*A�7M�O�d�/��Q![2� �� �^����O*TJr#�O�$`>�(�'N%[H�X��	m|��2d_2I�cf��<�t\� &Ϋ?�$������(ɬ\ �^!4�a�'i�59�m9c�CGZ�0��T�(}4X��E�33>$Y��>)��O04Y��'��O0hp�ς�LN���;+��Y"O�Yx�  "O��O�A\2F�IA����"}�ԘYa-\qO�q臉��A:zjBo-�d>2FnZ؟��Ip�$��x`"�g�`�뗤�r:J�*A'Ćx(R�'Y�J��'u1O�3?�7�Hi�8Ayw�6s ~�IE	x��8Z���?��dN�m� �,ԥoa�(���>}2NY��?�p�|���2H�d�a���G��!󑯝2�y�I�
�u)4��.B$�!��#�0<���	$
���X�KC&U��03ԧ�+�B8��4�?���?�p-�6�������?a���?ͻ��A�W��-���Fn����	��4O���A�'�@S������(:z�!E:P��
��A�Ȭ�#K�dЎ��B�P�����A[�x����"`N�yg��%�f��GSv�`6N��O�`v�����D"X@� kưמ����MY�a�ȓU˴��Ţ
b�9gCn�"��'��#=�'��*}�B�d*��(�� B��ˀ��/P�@�I��?����?�R���D�Ob�ӿa�X ���.:�&�p�G��R���j@)�<�qG&u���@�x"y�B�J�j<B��'w�f�Ǣ��&U)��Z����A���OҌ��I�p����u9;����1h�,��'a�؈�"ۃ$���0�Jܸ?��T �y2�c���O�i�կ	Ǧ���̟�맅�􈄸"��3�������I7O-���ϧ8�P��	q�//�Ґ:���<J�n�:2D�@�����58��O��Х�� us�gG
ZVP���'~d���+�'���j�I(w{.��3 !�Z<��'9,�X 爗����ň��
�'��7�Z<p:z�j��5ɀ��-��>��O
|HD����}�����O�^(���'��	�[�@2��O�^p�J��'M"b�0i���T>�S�? 4�+N�K�����FmH��>����t���O�����;b�����%��i��{H��a�Ol<'��?��/�|�S5!R5Y�B���4D�0Ѥ`�}L��s��?NHL��.>O~Dz�O?/�����`�(/���рǉM�F6M�O����O�\���Ɲ[���O~�D�O�N�pi����L��RZ�`$g�"	��kL<Ynµw2���|&�0��a���5E�� �����EͫH-4�%����mƃG�q��'�j2VAߞ?�@sq���m/V(qV�g��ɗ'_�mS�S��t���傐6hT6ex�əC��xd��~h<�d��e.�i&,�*�l���B�l~"�'�������d��t~��󤀄�[�z���+#?H���$OF���O����O�读�?�����Da�@�8�2�
O>yujj��աC���8g�0 �PD�d�[;�0=)�,�S�nE�s�P�<�-�E�S�G2�! ��-(G��Q �[��ۆ͔Zr��ǮF5��!���Įy� �$Gݦ��	����	ӟ��IƟ��IK��^�r�|�'�ܸJԾuZ��W��y�k��8�虠��5�@�H���:Ԙ'7�6m�ORʓXC� I�i��'��U�9)��R�҄8e�Ubt�'R�P�+~��'7�	Y��|��F�f�^l�@*״"6��0Dá�p<AC�p�WD��p���ؑ�FɚD��p��	,0P�.�DEy?&�3��E�]d�hQ1�`-!�d���Ds�Eׇ7H�x`2���+�!��Y�����O%�.�����67P�v�{�	�z����4�?����� D����|x<\����w�fJ�ɚ>�(���OX���ʡ"�pq��)^	J �ǩX�@���3"�|��5>ϸ�b�"<�w/�\ �O�}#�A]�WB:9@t�Q�^Pq)V���?U�ϟfa	�i��V��q��
�Ni �>iE�P��H>��d۟:y��k�;��y�FK� �y��@8*#�m�Ď��+��,�3���0<���(;�x,B�N�=�$�a��%I��۴�?���?q7l�;/�>� ���?I��?ͻ9����c�1��(�ar&�Pʙ]��aNǏE{T��A�"��O��1%�O�<��(�2b���2�\&"IԨ �Z"9��4��D!F�����{���nn����,q$�J�w�J�wj� i+8X叁$�h��Ԃ$�d�%���L>1��<]P�Jbm^�p���G�Se�<AK^�)���ɝ�>��݀f�Fy~�),��|�K>i���<u 8-� k�&�`L*б,Ql�B�n��?��?I�z!��OP��j>Y�Bm�+NTlNض-qr��Q�nC�	�y8F����"/oX�w!QE*�a0��S5 �Sa���oD�1�
��jT�t@Η'ђ4����G�uJV V��r
��`����*91�|2��	�Y|`���E�H��AN��~�p��S��6g�vc�(3�4��*����v�i���'l�|� k�/u���  3���E�'�) ���'T�	A��,̩�� (����C?chȁ痟�K`�ג'ߦ�R0�(�~���a��mk�"%J��h��F�&$��|��'W� ��h�!�MC�cR�u����=�!)�۟��4hЛV�'�uFGW)�j|�Eĝ�3�0���^�T�IZ�S�O�$��APV(���ؗ$Z����'��6휉��8��OсT�p�h�D������<��g[�n1N<b���?�-�~�æ��Ot1aCܸ�������w]�M��O��	 (����gP�qت���\#(�H���l�@3�˧m:P�W���t3k���O�US%$V7YD�r�
��Dф�5cR��a�V�
�����x!��=h#*�8�E�97k��'�NT���
oɧ�O�2x��0n�]�cA@[�(��'^�3 @�|��mq��� ���9��i>���$�O���pmL>[<�IF΁�e~�l�������Lc�H�uaV}�Iڟ������3iJ!�a�k��as%%��7�X	�d\// ��i�M=�)xFHŅ��J���=PL�y;g�4�Kb����Pk�bӯD8�b0��.)q�X��l6����������ZX�t�&���p$��&	�Oq��'�`5�mGW08d���Q�H}�$�'�ڈ��ǘÂ�1"󀩣3� ����X���$�|蚌sLl�&�-,���"��Y4��m[��n#��'R�'mN�ʟ�I�|�E���:���s���	wI%^5 ��qF��@ p���
	G�xЃ��d_����FZ�_��	��� P>�"
r'�uQD��)��(�cn�N�� ��L}&��!(�'{�F��3Z�);�԰P��uAJ��I؟�K��ΈmO�)f��#QdB�[�A'D��c@�EuN�Q�" )*!�I<�MKJ>q�O��w��6�'�B"�J�t���m�9ct�m��R}R�'&�`��'�1��|�"D��q*��_P ���#xc������'��Ҕ�*j8�?��lO�'�@�Q��L���Q�&2� P,!��
t�jAP.En��r�EΦ��.Q�8�&㞐a���O�@%����y즬�3mܛ!3h�ic�*D�Hp�L�$BX8�@����4�+���ݴ*E)ÎI!7PpL4Εe�j�I>�f�Pj����'.2U>و��Hϟ�s&��3�fxa"
�]֒��BGX������2Iz���l�S��O��2�m��
  R����R̡E�>y�"YX���O�R�@�#O1R1��S�T�N�+O�4B"��O�b��?-D�Z[����Fa�690�!��<D���$I�L�H��e�ZO6!�7b:O:�Ez�Y�tᚱIy��mPИ7��O4�d�O���E[0��$�O��d�O��Tx��pE�D��ƽZ&&[5{F�YJĂ�`��8�cJ!RzU�d�2�z≔!��u�������e�ӛ$��(��0��<i��W�K	�-H�',��~�I @xj""�v�Vmk&��;)h�E�I>Qf�����>�O
ɪ��F������@9t��q"O�����1��a2��V����Ě��ˌ�4�ޓO�=a��6��u3Q�+<��H�a��	 W,Hh�(�O��$�Oz�D�����?	�Oa��00�S��EF��$�h�a'H@	1���Hk�j��#�O� v�џ�3��[�l
f����4�������5B�y��U�D���+�-{�n�mڮ6�Tp#��>Y*�[s!�}�@��BB�f��D�$��O@م��Ge��a��_���D�2B�.e�v1S�h��;Q&�yUa���'��6�.�D�"=;,Emߟh��-p`@qo��s.H����m.�$�	Пxq-���P�I�|J�����*H[BԐ��!J�/Rx�R�bP�:�y�'	�@~F�j����w���s��,gI�I�	�n�FQA�L��s$�!� n �7=P�!D(z�p��C	j�K�{�G%�?�'�x�	#6�U�u�@�4�\�H���y2H��0gB<�D�
�1}2�a����x§zӮ�"Ѕ�s��I���|q���:�d�+�@u����O4�'!U����[�p��壞�:z����ӭ{�������?)�ÇC.�IӔI[f�T>ٗO��:3J!�r���$@ƶ �K����D��|�F�A���/_/�
 ղ��O�`SbȬub�5�P�φ<�N��K��K&!�OҘ&��?���`7_Zʌ��BT*o ��K,D�� '�ْE�N�a"ԩ���Ȕ�%Oh�Ez��ѐƮ�Z32]ӂ�Z��*7��O����O(���AF�G?(���O����O���ў�Kv�
3dF(HB#�T
"��pI��R�6�2u"�X*�8��/�SS�	��rM8��ˁo{�����
�r�\�쟙E�(�U!Vt����
#���OޛF��"�y��O�Am~H�S�L!^2!4�_o��O<!t�����,�X��Z
j��A��ٓ�=�ȓP����.�x����a�`1�'p"=�'��:�^��v	ٖg���d�]h!`�bwB"_nxq���?���?1f�����O<��*�x}�����V�v��"Z� b��� �o{�Di���*l	8�&�d�'b]&J�H����P�lO̤��E�j�(�X!Scmе��)Y�vJ-��3�{R
��_4���A̻wĎȈ���d�D��la�Ή�W���C��6��X1�W��y����`�N�����)k����Ș'Wt6?��K*��l�����	�@��%���yv��E =J$�I��*fȗӟ(���|��k��b�<��ч�&d� G�T6
h���ʫ"4d-۠( ;��d3��8ˊh�D���#14��B�@�jP|b��	�u��hC�t>���Ak����)��[qOt����'H4OƄ����27�x�q��g���2"O⩹���&Nj��R�.�x�!�EOTn	IY����`��Z����C� =��$��B����M{��?a)�T%6��O&H���S�D���y��9��s�*�O���M
 C����!W�����J�s��p�O���1X�1��V�Q(�bp�I�\�'���9� ��=�������` T�����W
�<V��)�W���� 6!Pi{6�B��oF���,��S��ަ�Ӓ���Q��Ӡ�w4r���,��6H���ƴ���v*���	�HO|Y�^#E:�5��SJ�\���צ����d��<`���D���\��͟��i�	r��.�t�{f� X��hXDE;:�T��L�-g4(酟E:��|�O<�G�� O�4���h��M_�$�r��LBh[��N�8�]ڤ&E�%TdT�L|�	c�r�0�2ﾜ��P4J�R�k�gԑe �d���Y�	�g ����|��R� �x�P7K��1`(��ybc�!K���Hq���L-2�y2���E~���Ē|2.1?��vKǍs�N�PeM�Ms��J��%l���'2�'!��]�����|�`�ĵMnV�"���F���y��;i���`3a<����G@,����ۛ3�<`�ף�g��.���1&�F
Em�2!I�>s�Ѫ4�cp��σ�kR�!H�{�A�u�? ",J�
��R�����m	BԳw��O����I�K�Z`!� U�B�
�{U���S\8B�I�u&��Q�,�O9��k�oK�b�8�ٴ��U�"�0�iW�'��q���)&���ipfN�?��|���'�g�'lB�'��	2�C!�B��R��1R�~�YY�
�>2�����F5= f {�g2����2G��9(�x�����y8T� ֌J9>p<5BL��.@U!��M�� N�\"l%�=A@�]�|1I<gk�}�8Z�OT�v�����g�<!`�@piJ��R�Z�C��;%�]<ٗ�i���kZ�<��`��j�R���|�e\-J�P7��OH�Ŀ|:&�/�?A��A4^�>l`��H�6w��T(�?��MV�Jp�À7
 ��W-L�H����W?�O��-[��%�0{.Bh��@\���'W�\<ё]�kR�ڵO�+1=R��.!҈zwG`>�w��x΄81䴨�x"��1E�@Jt-�i�N>��f)\,�x��)\��iLM�<1�$ҕ-��9�M�)E� Ia�K�����$߰p!��ǚ)9h���ł~a�	o����	⟠�r BH��̟P�	ޟ�ݡ	8&�A� $|���e+^W>���d�)�j�A�K�:�qUg�a̧|��!���k�B��(!T)����8�Z�1K5dN�-��d�/*+ʑ��M1�T��U>�D��6!�N��;A����3���0T�>�n�&��T�Oq��'m�i��ߌw:��Z�
ѓ%�j�@�'ΐ-8� ��k�n��5�[2 >XD��' 9��|M>q��=H��$�ʫ%�M��Jȃ;5D�3���?a���?9��2I�S��ϧ;�����i�\�R��!�:}��i�:��x $,�2U"	`/�-O��Q���#�/��X�/�<2�]��n�7&�Y���Y�q�APQ�Q	��Bs�ֿld��QԨ4ʓE�JQ;� "R$�,��[2_�R9�֤Y���9ݴ1����'���П|�?��AZ���!�(��Y� ��Kr�<aUO5l�Ơ����Q�H녭F�}����'�剑D^�X{�4�?���b]��e�M���@s�K4F�����?1SB��?����ԁ�U�dh�Ϡ#,Nh�1ڸS�8 ��5]��@x�S�zyq�H��;I�Fy�M5o�<� t�ב7���Xn��2�tMD��X	�`��	w�	a��ڤ{�B9Dy����?s�x"FJ%n� ��c�$�4� ���y�L,Qx��@�	5,�X("��� �xb�i��qd�t��Y�VC�|v�)�0c>���>B�-nZ���	o��`9��E�4kA��1�+��i�&�)Cd݀eP�'�l�k��"*�xTC��YS~E��Y��|XPT>E��@ _,����&n�@i�M8}��K�������!{����dśv���pW�L�d�ݖyk`ЕM��x�a2��I:��$L~�)���=���Q��^���(�T�fC��	k��AQ��Ԛ"�(,9�L��*���UE�'����wCB��~����v��k��j�z���O���F�2�x����O^�D�OJ�4�±�E�4��k��Z�0�x��呒%�h9@�ʢ/�ns���7?x�c>�&��`4H-db��b�o]	I���u��l�����Q�>��N� @F�>U'���b9k鉨��B�XO�$}$��;B(�Oq��'s~��h�������=>�V\�'Y�	5i���0�'���3�bL��O��Ez�O��'7"����̿L� �����?�@{�IY�X��'���'�B�l��	ퟰΧ:�!`SHGo�H�T�7��$B1L6���iT�G�����'+��m�|�1�#J�Lن�Hq�Le�L�5,�LrP�E�Փ#�n\�� ��hO����~�:�>�2]q�Hɞw{B�'h�m���\O�]�C,�3j�t�'~L�h�+�0uɖ��抰W���yb	u��O��qd	Q�%�	ԟ�0�W5��19����nw^a)B	ğ�	�F���I՟��	�.�Y��S�~1�Ѱ��i)�1��aկF:x�U
�0c�5� HT�kuџ�1�i0,����G;bu"ePƬ��N���v���l��L�`C�7A� h�fW��@���I�M�i���ONE<�QG��Z�jA��f��'a��'(��d�|2��z6�-Z �Q!v����
�y��'j�6�E7�J�*"��9(@�y*Ƌg��m�Ly� 8p/6��O�$�|jv�(�?Y#�@o�9s��	��D�?�Om� A��y��	#��G��B�DJ,y.�,�r���HS%^��|���u���U�>��gN<L�칙��7f��ѓ�K}x���GW ��ɜ]�<i��J̒8-�y0�Lm�&uZ���{�S�'6�l���e�~ĺ�;#@�6N@��ȓ(<��A>Fm�L�pdZ�q�!��	8�HO*��%_F���i۲B��5�u;O���dޓ)��x��;a3��e*�f�!�D�oE�¡�6)06%��(58�!�$��H�ZE�q�I1&Ł��V�!�� ^��-S�г�ՠ^�l�PW"Oƈ(�
�@`a�^;_z��
�"O�Đ�j��,�H����ߔ}���(d"O�`���h��= ����R��q "O��p&���1;���hY9~X�]�r"OڅrB.�39��XCb�ۇY-�Y��"O��	#�R�~��2� 7��X��"O�Mi$�6�d �ʖ8n4�g"O0 RA#�#q�S�("UPE��"O�h���y���2!�B�Q :�v"O�Q5�W���B��L�2�"OZL" p�j�A"��h��	"ObQQ�N�'�Ta����1�n���"O�hB�̺%|�J��ť����e"O�{F��7b���S�ؿepY��"O���'�ٜ7Ȗ�pf���R�Z�"O9h��ǅ!��Q���@�~�%"O�hK�Mܰ9(8c�&�!�}�"O�$�%Р2��
�F�<"�*�""OBP�a�O�!�L�E*4� �
�"O"� � ,��eJ�y�jE
�"OlL"2�&������yE�-X�"Ox��w]�c� �c��#4���v"O�(����Y���z2-�@"O.�����!8���#��C�r[v+�"O\ԪC,�"&b��e�!�Ɓ�t"O�����;Inɣ�/Aj�,mct"O�ܺplw���Z��N($��ّ"O���qn�b�����&����0&"O�{�hѻZ4 UY���*l�"O.ళI�E=�H��)��u�p��T"O���#�	+�^��ǞI݈Tf�'{^��ώ-	]�Ub7O�]0@ZS��jq'M�|�ި����%��tR4�V��z��~hӲ5	��V�O�|��-��B��ēy��Yc��sv lX�.1ڧ, uj���w�H[��-l�%$!NL{��{`N�e�'>�[�jm�MC����(s��Q�e*&�Ң�O���4O�s��;�(���/=cp���GP"����2���&���\(����2xin�AsdZ0W�(8"tX�)���>tǦqI?�)��Źz�ɸ"���J,�$�ܨўru��?'��	���T�R0�*3"����7�Wt���4�E�iX9��&9�^sF�傞�UF��4e'�%�$,�1p�ˎ+
�B�b+�p mZF�xس�hU�^�d-	.d�X#?��e�iS�5+��M<$�Zt:��Y?���I)E�� kѪ�pT�I�6D�T�'2�����
Q� "W;O�e�"�O�:��Dá0^���'H:����C�4g�iK��񄇮O��̻|g�I��5�Tt��T'�����7��C.X�YL�Y���#(��sd�V��hOr�	�m39�d*� Z� q��Y�؛ghN+JH�b��!� �2�.�9�u�����0��!n����ɴ	Z��C�B
Z�H��O�4�&7M:�\I�EI[?I���ۄ�Ƅ)��� ���3~Z�[e�ٓr��Z6�-].0�=��9�g}�L/{���kՙmb؋�C��v\�����)���qOV٢G�՜!�aӉ�+]��)��b�:�\�v�>Ot4�h��۔$R�N�fmC���p�A@��fܓ�hO�i�%�Eh�C8R%l���-�m�-�� �0�HO� �)�R�T��Ė<��c[��W��7*܋��ҽ�bl4��?�S��j�݉��"U�Ҽ�bdD�gX"$��A�mW���� c��I��(Т�h�K8"� `*�	�H{B ���iB��&9}���� ����YY4 �s��~���c\w��=q\h�Z1�G+]��hF�EKz,pX@�X5�d�Q�B�I^�)C�H��ߏ�n�B �D4ֶ��6,��< ���ǓSQlY�v:���}7<�
0c�␨�Q���?-9�F%��~�!~��s�Ê@��ʧ/����;���p�&S=n��I������2ĎϽ<�d�I���b�ZQ�>I�퀲���3J��V�� ��I�(��4y|V�r���O�d�� '��
N��:���+<n�	`n�<g�l��ƒ�I�,6�Ӎ��L�㤎�2��Y�0��%�qO<h�P�s�(X��PE��2�O�*%lP�摂�?	QL�CztA�V*��=P�(
�hO�U�.D>��uM-S$X��u�N%!lB�=yħ��~b�OH�g�? f��$��1�!�hO -vF� �m��h��# O�����Y�kL"��hW͐�s��1T.� !,qO��	k�ĳ| �� ^�D��SE���a��OqS�(q��p�'���WM�1[�`��Ga��̉^}b&q<��	�.�� a�6�,�?K�����'��{!�$Q���2��b�"�u�S%�%��!YF�,�M�eI�N��%q�, dK�݃a�d�'�\�!��ġ��I0ٻ;�0�����:pb�IF� y�j��U�|���hOD���f�^�j	1���K��pF@�j��G"�O&��'� i+�O��2�D��%�H�h�چ��x�*��'� `��b&�5��~�P]h3O��!�n4��B�8��'��D<����D�$j����3�U�=5
���mA�Gp�#�/�a�ZݛբƾZ��겨ЃM8^��'�`Y��㏅t|��+sIŝdmP�A�{��'��B5_�,���N���%i�b�?���E��q���8�0��զ�x���b�� ��'I>G�FU�)�D�Lsq�B�N]bS�N�	�PC��'g,M+���v��E�4�Lq����V��8�N1	�l���
��⯅ A�џ�>QM(m0�����9 �n�
\Q5Ѕ�+��p<��#80�DԮ18������4�"��n�О��=a��'�~��l<&y�͚��FHt�Q���I�>i&��t�=ғnf�x`�zA�A�ìV�t~A�'uJ�ѷ�K*ޔS�nс�j���y�f�Oj�nZ)yz�xKAʋ�!��v�OӺ�V�'�����}T�5I6[=Z����4P�b�Q���fI`��O6QV@G~2-�(`�x�b����U����HC(3Ӓ� 2�$���(��I�gl$U�c*���vۯ1���y�NB���?!�L�{޴1��
�����8O�-�#�];�p<S+ܚ+b��Wf\а J,n��}�V���~2����{c����i�nߙOH��B�JK�'�Z�3IN!?g4p���d�L p�O����/G865���H�?vH�s�I�Mr�aWK��Z����g��pw��$VnB�!� O�C^��+���Tn�ƥP�sd�+v�[3�vt��]���Ortj�Q�$5H��g�
zK�c��O�$�EbΘ|kV�Y&MD�:4��	2l�|�q�ޟ,�<S&��
[M!���W�Q��~�oщ*����Ë�l�yƍ�'y���A��0?1rHM�R;���Q톮�^`PS�V+c�(�k���I��H��I�r0x ��*
�����d��=i�l�<L0)�G���:���#�B?�'��3"ֈ)�,�;�J��� a�'}��sN�:qe��zC�B�w�"�'�h�z����^jt�����zv��4�4��C�6�bq�V�5���D~2�M;�y0�g�V8YR�؛�~b�ޣ� 9���ٲ
F�]Ӯ��hO��p��FVpL�+4�J�CUV�pc�(')h�����s�i��훬 ��I3�+�Q��:�ǀ/]�Ȅ�I@#(�;&����"�:J����� dg�0���9n���٦K��>�<��g �
�>8A��G���88�AF"_Ԟ|�7F� ����>ɢ I=N����l�H �]�d�
}�'���� aٟNK�A� �Ε	V�����UslQs��]�D7�)[��)P:�o�*������eK��1Bט����d����I׈�y�@���-f�"p����̙*�@�h0a�K�X�ԥi��"�Py��DǢ9�(�X�CG�A~ �[	�a���,lٚ]Iu�ΥT*8��P.�`������ɵ��xr�S�x�杫l�.�*�(�c��C�^�z��#B'��0�\dys�G���gyr�ئ%ޒ�P�䜖5��]b��А�HO�%�Bd�2/I~�CvF�:m.0�QP��"aԠE-�e�2��nH )�0I�
B�FXЊK�mc����	2T�O�tAA�|"�G�v��keB�z�2�;Q�Lꦩ#��!-LisGK�:�
�KA?�y�8��Pl_$:���Q���6h������v�h	����O�KqҪQ�n�bT?<�h��T� �DR�A<��E��뼣@����,0AkN�K��9��E>J� ���"�p<1�D�Wy�.�I����R��F�B�.A� kqOd�K��Y�u!�I�3Ե���<	'�
�f� )cWO�#q0��Tkn�'�p�eP����/��x��d��OXؘ�)�G�p�	D��SaX��t���Y�x@׸ ��̆K,�'���R>�@D�A�����?���9F�l���4��X�����O�OH�3���K���܋o

�!%� �$="�b<ev�����0�d%���?�Mx�i(Hi��� �#]}��o�`��р_���拀Pt����r���6�Q���X�����I�aW� h�g�=�p<���Wda�N���D�"���- �X	W䂱MBBGJyb-L�KF6�f��H����	'��0��~"q�Uk+m�"=�d��3O �r^/�ͨ1��V}�gK4 ��,`B�~�r�f�Q�*��E���"f���'T�K>�����<Z-�ic��3v�qX���QI�F�Փc��e�Nk���1"Y?��OFa�m]6������	�wˈ)��h_P�b�(��`$�gyB��2Sà@s!k�/ �Y�NҼ@)11:��->L�oU	s�<�6��e���&]��H�I/�!�GdC�n�����$����� �����^�^l��@�1V������+>��Sf�\�H%x����Xֽ<1��U�Z�s.��2T�JB��r�'Ք��pɝ�-�8�K*Y*z$#�'�\A H�,	n�TB�Ԏy!l̩�c4 ɐ�N_$�@�I]��Ov�	ek�|����
�\�a�.�*��ҡτ��S	�+r,֤�T�����Rp��O �#�f%��4v<�$1Ո�'�&�9���
�PIc�+\r�JiPH��'v�,��%3$E:�	䇕�x:��9e��|�B6�@7�|��O/��?��0�8��ϐI<��#��Íi��HeC�c+���O���H�:�ʘ#LM a��}˱��
Q�٢��)r���"z�Da`#�C�ԕ2A� u�*�8�{��j�n���"=ISo��3X�����O��H1D�����8QE�%v�6�X@ ��@j�a�b�M�'��2Tb��`	:|��C�E�O`�:	�%]g�9���9�\2`�iG ����\'u�\r'뚥+���s 
�+zN�pP��5W�.Y�`���uG�N7r�͓ �BX%r4-ո�~g�$9��,�"��))ƌ"U��&�hOQ*&J��Z� �sG�1�c^��#lD�c�J��� �JV1.K��4�~��O�x�OݢPߨx�'��L>�	 ����^x�,�:O2��"�����:�h]"ibp�2�ɋ�3��c�FJ�C�V%�$_;�<H8�e�+v.$�Ey�JR�IV$y'��ĉ�B��T�x5��.�{�')޼��目,bDL��H5|�Er��ŋX9>�A���@���#���J���b�	
`���s�@�\�D���@��Oxt��G-Oe�	�扙-�z	)$�i��ᡜ!\�=2�	EAE�����:^J9�!�3s���V@ ��uW�ޜ5��8�ӣ���b<��J��~��Ѽ^|$Z�Y4z�)ag޺�hO���N̼b�"=B�ՄH��r�'W+D�) /�3T��M��C<G:���Fܜ��3?�0��?&tm��F.�4 aBũKS@��gJ�fX��+xY�u�J�:��@C��%e걀�M���E����O>�RV�+��Y��O-tݨ�Eқ�*E��K�@	V�i˓w�T�4��z�צ�O�����2!��!����ht aE�!n�*(V �9�~�	(�H��ɑ��tP��
 ��4f�rOB<�1`�|���8�(ƹ�h� =�p��� zXy���H%V ��w�i��Lo����ux��A!ẼX+�e�*k1�@�g�8T��=��*�<�a����A+�Ħ�*e���5�^�Qu�,�U��"O�HqJN� T�˗�� �Ȱ#�"OЅ
��J2*�8s>%����"O�x��eՀR˄ I %�Uެui""O�mɗN��	�v�3D
� h�AB�"O�K�@�!D�p����T�B"O� 10��\��W@A�\4R	��"Ol���j�*/�y��Ă�o+��8�"O40+!$�]'��J��W*4���"OH%S���U
�-�(r��"O�m)Q���rM��"M�D�|jg"OZy($��(Hz�ɵ���$I�"O�� Ɓ�6�60�@��*�u١"O���mi�,H���V��5a�"O
�j&T�?�"�8�L�d�l+�"O�H�Q�>k�L��1O^�f��3�"O8(�C�^�E'�-��n��Ok�}T"O�����J:��r�	3�b�Ad"Ob('+M�x��BMٮS|a1�"O�,��d*
a��Y��2����"O��3Q���`�&�22i��xs��r"O��a3�6 f����C	k����"OF��`D\��8c�ȎVfΐ³"O6���dǷMa��8�G��vW��g"O6 �e�S<M�p��E$U�� pr"OF�)q
��̠�������B)D�|��#K�I��st�(�w'=D���ĦC� j1����1!~ڕ!1D�X�e��%������Q|��Yw�*D��6�9q�<<���,0�vIR�e*D��ѵb�,3��Ra�ѝ[�TU�6�2D�@��$NQN,��c�W�a�R�0D����=����eJ$dݮ����'
���ik=t��gC����d��'�=���H�5$t�ڗ�Z��8��'+���r���)܊��M
#M�(��'>4�1�'GB�)�ӯ� !��� xܘ��Ұ$,�2\
>�� "O�x�fM�H2fD�')��ބ�S"O(�J7Cή+�Q�pH�� T��"O�1p�·)$�$*&��>���XV"O�1��� .��p-�-88F59"OZ���,I�����m
a3ț`"O���w Cd�p�Yfo��T-�%r"O2�3��GaR��Cǎ�8��("Oh�b�&�{��| �nϸx�\���"Oʰ.Yn�QwLC� �V���y��� 2D��b@Hf� y6�$�y2LM�Xm���rj҅Y)�@l���y�	45P� �-���ʙ��)��yb��(��Q�(��;��3�&��yR��1C6�y!�0�P�!oF��y�oT�X7�Hɑ�½�ݚ��C��y�+N�c V`���ާWx(%'f�-�yB!M���PgØ\�`�S���y���&����D���֭�UB���y�-��fF�ѱOE&P��:6�^��y��·H)^�����n��!���ڷ�y��̜3�t�-[%Xb�5��-��y�N��3�:�)�%·V�x�QJ�7�y�� 5wu��k���E��S�g�)�y�K��7���0��D�T��fQ�y�]�ӄT�bGO"��cP���yr�	�hp�10`O�;,`I��y�9i��l[5;���׏���!�Ж	���JI <�`2F%�6
�!�d��h!3����&��T�!�$�w"B@��%|�p1�?l�!��4����pj��c@hb�\�!��|v]Rʞ�Pi}�G�mũ��7n��ɟD1�I��G�D�����.����W�z��� gR�Y�$T�ȓ9�vz$B�d�� J߄}�pՆȓN� �Ҧ@.'k�� �G\�BPXԆ�DG��+�Յ	�����Ծ6I���ȓq��#	ӕ`2��!�E)�
ņ�sR�)���M�<q��'M�m���hO�>II��p�<��l͘r;t��Ŋ0D�h��e��W;��BB
*^����k:D����"�;F\�6�XxE�C�*D���ł��	SD x��	.�BჀ6D�x҅�Ѭj�l�����8Nf�JA�)D�p�H�G�m�!�A�,
�4D�<�,X�Z�4`�*��L�6Q�D�2D����͏s�q�$�8Xb]+H<D��� ��/i��ر!�Y�{�r!Ѵ -D��W�f�xI{�&qep�iuD/D��Cr�ľg���@�`�n���-D�@� `�xS�zw.Q0~�,���C+򓿨��P��I1Pn� G���d�"O��#�M� ������0�QS1"O����	��С%�	d�\�"O��97l�&<�4=�aJȯ48�J��'�1O6Ā�DB /�i爛l�2����X�O����o�\;�K��Af�a����'��>�	�2�:z��ŝ`�@�;V�ώc�
���1ғ1�p����\Y�^�P���c��ȓ?����!m�G!@�p���d\�ȓ,�)��F��8R`��	� ઼�ȓQ_ l@d��nI�Ě�@H G�H-�ȓX`��j�s��)Jt�f�2Ɇ�S�? ��8�FG�':*�C�����ò"ObYbea�=H��qTg�'L�8���"O^��1ƣ6��	� ����P"O�|�׋X�divd����@��"O�e�ā'X���<d�"l"""O�I���)h�H�"�[�4�@�`"O���#&�b(���jB�=)��'YqO��	�{L����L�:	ĶE��ǄZBB��+R"՘�r"x�֡9vB�ɒ*G����)͓�h!����d��C�	�7ߠ�;����-rBq3
�pz�Q��b����I+|���
�a� !h�K'�FH��C�/KK��Ɋ-A6*�ȶ��N�C�	2%�X՛bj��,���0hC��C䉲[�@���K�D��RS��c�2B�I�<w� (cE����4���	g�bC�ɿ2T^�3�2+r*�jL�m��b�h��	y��,j%��4�D���I�_f����<1�'��V�Z�z���!Z�W�F���bR��yBl
6��z5�3|��آ�y�Ǒ�-�p"A*�M�|X�QL
"�y���~�h-C�!K��ٔ.=�yB*��^Lb�3W�r0hc
O
�y� U�4��r�l��R?������y��D�`)t��@gD�!���	�GF��y� ��>T �A����������y�ͅ� �X'����0�Bd��*M�ў"~Γ,h��g.Y�B���x8bф�i�'@�?�+7$DG
��`��! �ԥzGHsӌ�$&�)��qy5��Jz���Y=[��2D�L�[�y�1�|��p8j�\f�	R~R�'-�p� ��5�:��&N��0�
�'���a��n�\K���*M�$	�' �Ȁ��'.:H�� ^�9�L�)�'�$�yc�2�p<X���$M�%��'w�<��WW�Ը�!)	r����O6 �OX�"rG�EP*A��	�H�nEX�"Op$����/OpJS��Z���`V�i��$�]
d�r+��R�O9"Q!�$DdM�w�Q�@��Yk"�SC!��h�Q�L�3�,p�K�:qOҢ=%?�
Wop�T�Q�_� �#�����,�u�(��&��s9�����ICx�,DEZ'&�\d��
��$[@��!>D��1��8G1,̛�넭$���c�;�$(�O�����lY�!1����!�(�ᖛ����I5J�VJ�b݄k�}k��_!u�B� l=$1����/��ÁJ�+'�B�3m����Ϣ5$���a��]eTB�I�0�҅ �Á3l�e n��B䉧� �@wǘ!̨Y�a*�5�C�1Lo�yr��٧+�AZ��Am��C�	$C�j�)�"�be.,���S�t��B䉳f�<��Y���3N�_v>C�?zB�4p�	�$����:�
C�ɞ	�<��p^05��2��ڦ��B�I�3��S#�];5�� �G٪.i�B�	2���C!��A�Vܳ�H�>��B�	�~���C_
=��S�Ή}9dB�	�ww򅮊~Z��ZFnK�S�*�'�a}�n�G������^ri�$ּ�y҇�bp��A���dhP��s�ś��'.N��$KN�,�t���N>�BDH��!�G5h�����k�r�:���8Q�qO��=%?� |��U#�eI�8���Y$V0"O��amưyD��C�D�h����`"O<ݐ�!�4�hy����MK�0"O*��5��'pa����ő H'��"OP8B��dy(!hRP(4�ʁjW"Od�c E�2��Z��9ӀbѦ�yr�L�!P��D�O8���N�,y"fB��j?�ɸt�R �E���n:����+����Y�U"�	'Jh:FC�)��B�I%��yr&_�C~��t�N�o]L�C:� ����O��r����!gǈdҜ����~�D���Y���p5�#�hO��𤙋F�N|:�b; �,�pI� &3ax��I�Mv\�)q�PE���TM�=�TB�ɴRs Y�iOlT0c �i�.B�:XB����`�hi<tφ��B�3�Ub���H�	0�T�aQ��剖�hB�M�"12 �r*V�F�B�	-L�fXPTF�:i*�+n[�]�IR��P`�d��`3�n:�~�'D�H3d���t{$�E?R��$D��[0L(a�F	��!��B$���"",O4�<!��113�@���Ȋ �Ri�~�<�I��:�����͇/N�A���HQ�<��bb�#�ۿyF�ٹ�XM�<3KJ�-È��f��=TIc��G�<a�ӽyF$h@ٷ$4��:7G
D�<�@T}s���ЁC3 �Yh�u�<$IU5o����-�=U�tz�C@s�<9F�-P48X`I�g!&���b\r�<٣�@ r�,)VK����a���F�<Ae-�:05����'L�S=��"ɖ|�<I��4G����Z�S�a�Qcr�<)�����[q�S�R�˶
�X�<)���0Y)�!#�K>��Zp�Q�<��a�/-D��q����M4 ZS�GP�<)!G�	 @�t�qJ�3�\Ա�O�I�<Yr��F���぀�8Ch��eE�<� W��Ӵ��>.B���<��`D�2�� ��⏇,ll(�Bʘx�<����%	 ��8�A���3�q�<)e.�+l����A�.�`�7�Ci�<�Ѯ����K�[�x�6
`�<	���Iv:�h���!so)���]�<�Q�ߵ9��C��5M*�����Y�<�U�;k.��"�M1� 㖣�@�<qT��H/d� e��+p06�b5C�f�<�'�^��aiH�P)��j��]�<ٓ�ŘN"I@A�	i�Ztb�e�<��	�	4jĀš>��	7&a�<�f�Y|x�2'F�Z�F��n�\�<�q/�	 X��K�lD�D���N�<����8����u���F��3�LE�<�"��;͖e�C�]-Yݚt��`{�<���=
��أ�J�=lP�QV]�<I���=􅒥L'0dY�o�S�<�r�N;/�2�x�E	��(1ʌh�<���TIH�� ��#�vm��`�<9g���j�D��d�3tЊ�xV��g�<Qe��z�:Mt�29�t�h���`�<�ǨU�<��	[�AF-\K��uf�B�<��l�;P.fq`��ѯ=&�3w�@�<�L@��nu�vnٵ2A�a��͑y�<A��.g���W�p�1�C�@�<� ��S��Pm|�,�ӌO,.����"Oz1�B�F�:\��sL�%�]��"O�#"��*0�@�l'�VA�&"O�@��G�T�����8���ʶ"O���OE�6���*�D+�"OΝ��$�,hm+�/ؑa7\DK�"OUɡ�Y�\n�TZR�	Kru١"O@�8e�Xt�R4�q�*:�l+�"O��r�D�<T�q��� 1I�"O�a$��e!vԀ�hB�K��a�e"O�D�R+8��dk��?2���1#*O�H
�dݸ0�a`gM.�p�'<n�A�LݴglD!�e̅D�2 �'��88"���_�� b�J[5��$Q�'X���%�L�0��Ҹ}El�	�'�Z�K����@����o|�q	�'$H�4d��/�0�Ae�V�g�"u��'{����HӠM�v�CɌs
VZ�'��1���@�P��&-Ǵ2��'�0�
&��"7Q{�A�	Uv�!�'�R@�����h�X��.3�T�2�'��(F&@g��DK��`Ep+�4D��Q�/ȝp�E�*s@I�7?!��>f�-�͖)5�J���Θ�.!�dM�Ez�x�����ec����!��J�n
I�̆#:>�E���ф;!�j�(qc��GI����#_��!��)5O�$p0l�-��(�#� �!��;����3jO3���T,�J�!�D��	�X��$ͦz�T9�l� !��Y� ey��0����ä-�!�d�	X��s� >ڮik%J�iP!�$�> ��Eb��"1�1��+rV!��"��-@[�,��@�_�"���'�� ;"���y�pX�+�PS���'t&9���'4, H1O����ʓmr�at	��F��A�q��B䉿~v�شKE�!�^� ���T�C�I�&���H�6=0�;��\/�B�I-YS�<�T%	� �9� b�)+��B�22�,0*B�C/m�܍E!Y"T��B�Ik��4ђ�	/�ڡ�ꓶxӈB�d�:.�~�=HB�Ӥ<2B�I(n�2�"��ǩ y�t#@�Й!��B�	\J�$��k#��Ph�
� Q�bB䉗J 	 �IV�W	�S1&]V�VB�� ��)�f܆^�����]��.B�	�	�EL7Vռ�jp�2��B�Iz���`��2ص�R�Zs2�B��4n1p��T"�-���+�E*R��B�ɛZ���iq%m`p����p\C��up��H#@�"2Gxd��߬2C�	�E����E�0^9Drt���7�<B����u�`\%!C��6�ٳsI�B䉧r��ƄG�c���1AA�=�%"O<��Lz�:f̻8фR�"O�4ȴ��5|D��:J�e�$�� "O",c�\�JF���2��>Ɋ�(�"Oj��s˘��(��&قK�^�5"OΈ�1�
1b@*�%J%R�X��"ON�s���FuJD�A��h�`"O�`Ԩ��P��X���/�XB�"O$� �@`[��2ăL�6V ڦ"O�D�C�݌&�4 �chO�D���s�"O� ���gg�K5=��,"C�j�*�"OT|��DE.W`�!���=H���"O��ؑ	G����نn�T�H��"O��#��G*iN�9˕�H�_|ڨR$"OP�ٗ,��>��<�ł�cz��8u"Ol���96�� =gϞ�a�"O�13����ص�'`ҭM�F��"O�+6	�-�  ��Λ����"O��@��]�!Z!"&̂juJuB�"O�Cф�}�����aT]9e"O�)�	���00s��W EBG"O�E��NQ3lB�S�ć�+�er�"Oh�Q� �G�L��`<~�J@)""O<R�H5�Z���H�=�z�.�yR��!�D�����Eq M�vaĹ�yBJ��<?��8�$��s��M�.���yR+�y:����;r��\Ӵ ��y"@�%>= uۆ"Ͻ�R@��/��y�f_�Y0��E�X؅�GT|��'�F�
�����C'[?�� j
�'�j���"ˢT�Thbn�>��	�'<�ҧي8sp�9rd;8��%�':��kǍA�-�0���5�z{�'�ѐN�`^�bB��+��ً�'�T���Nzfb1x�M/'�`0�'��Yꙿ}��d�q��! ���'�(��@^�;(E���{v~�;�'(	��
�� �I�ʝ�!��a��'K���I�.'�(@��ȡ.\v�;�'��s��&[�����V��'�����/�)�� h���h
�'�|ESY�P��,#�eÑS�#
�'%���dC�6զ5�R'�(I	�p��'¼h��$ʞ~�Z=qRf�0L��q�'�Ԉ@��gp�hA@<��\�
�'�E�bG��0��y91�$��e�	�'^�r�!�+h:�ܣ�nB��(9b�'6��V'��P����1��'�&�I@B��I��=R���'|�P "����|�ޑ
�'҅E�&9G�eyfj uǼ1	�'ڦD��R2�jT1G(X�i��TY�'��|Ҋc.LT�e��\`l���'vXx%@�=�$8�v��6c�R�'C���k��<R��&��3�u��'�]a#+������ć�".j�<h�'��RKڌŪ@���%t��'}jaq0J[�q��)st��Sdlj
�'g�B&Q�k|��D�غ�
�'�ܑ���xXԫ�	_o�[	�'��� ̂R-8�IѯA�θ�	�'�4�:Ƌ�$ax�q�R�<���'����JU	�n���H�-4"M3�'�����M�4!�~u$Aɘ!ɤ�q
�'��(�ƃ&W:d9SN�+��	�'�T��פ\�Җ A2E 
69����'�^��r��:1���k�D�,- ���
�'`<��`��Y�84$��� �܂
�'��M���	�l��ň��*R\�;
�'�\ɋ֣�8p@H0�XKo�ъ�'ƀ��\A0���O%�xS�'�8M�W�D"j���h��˚3r���'��h���������,XT��
�'��  �@�v�hi��]�N� ����� P�����J����
� 6���"Ob�2��=_bN�(6>���b�"O���>9:�%݂d�*��"O�};���I�H$�b����Q@�"O||9�ˤ%�5%�\�7�p�#"O�]P$ä;k$���^B=p��F"Ou��*)3������	kAzm+r"O*`z�c��[<|*�i_�l
c"ObĨ�睢k�z	����"�F ��"OBLq�	��0�2�+ㅗ�`���t"O<�dF=I��L1�N߄Nq� Be"O�D�aʎRa�qʄY�v_�X�#"O`tҲު+���"cH9UN-#�"O�7�D�ܱ���KSP�G"O8�pO�!�����G�TC�`��"O��A�IO5Z�LXC��5���IP"O�����6��v�wgHѪ%"O�t���U�!�@��͑�8afyд"O�L:q s$\4�Rm�mH0i
c"O�� ��F�`زS�P��R�"OĴ!���*G�\���E+���g�<I'�u�,��d��m  �R��Ҿ�!��)��wDIH�d 5�QG�!�� �2>�ŋ]&'��=��G�Vi!��G�J��J�I�*6��U2�JPxu!򤀞hȀPZ�@�rjda��IG�Xa!�a��1u���|�uH�OV�pR!�ǋ$d���4�߽Bf�,&h\� �!�D��y����5a|x�U�5�!򄘗=��8[��X�V<�yr��!��:}pX;V��Z,�x�D܀�!�D�@�j#�ϸI�իW�̾e�!�dK�#�P`���
s_ �6�ȑ0�!�DP>{̼�b� ݩ`Az<2T�G5g^!�d�S�
�KdOAz:$=(���fG!�ǧz~�Yk!Ȍ5ؼ [hC'S!��C�%&�tx�(a͒I��G'W�!򤉙e,r��Ն@�1#�t���a�!�$>�\��g%ۺ	d��BD���!�dP�J�x���@'~��A���:�!��R�+9*���A�Z��ݐ���M�!���s��9��Y4x�V8��
!���*�r����K���P2슛K!��"C�` w�ʯ7{�|ZW
�*~�!��Cb)�����"bl�Q��S�-}!���4>C��:�F�T%v�(�n`!�D�4P�X�я%�89�v�JB!�d��{�2�:�����}
��F�2!����v��χ� v�����9}!�_  0 H��Y�ael�)1�]�]!�\U\J��2�?r��Y
�H^�|!�9��3�/A>�\��Ǚ�S�!���#�b1�V�A#k4���R'+!�$TC�)�e�14��r��4j!�d�&<0�y�t`H����9�E���!��4?�إ�pB��-fX�3pe�T�!��1H� ���L�4`�2=HP�G32!��X344$L`��A(�Fi����!�ҥ6P�����<���9S�Ut!�č}���@ʟ�:����S/;e!򄆕01�ɩ�e:~�x���,�eF!�$J��h���,y�����:_!�@�p�<ك�gC|��P%�hJ!���--��,�:O
�Pj�;E!�� �0���n�$�00M�h�bxk"Ol��A�J`��`A#>t�"O��6k�5r�x45�X�&B�d+G"O:P9@e�>`��`5	�9-+� �"O4T-�kmf���FJ	bE"OB��S�ޣ,>��h'��(�l��"O@��JV8`�����*�(�Rt"O��A�I�
$�PՠJذ
���w"O>I��c��?k�����MOS�C�"OP�K�.H�7yNA#�AN���S"O��K�(��S[���U��,��L�r"O����ü0�Pz�e�L��M�c"O6`覯�2�yy�	��L�jd!"O���M�W�$�r�)͒T��\0�"OZ����e��	/�W��!hr"O�:>�4
���r��4�q��	�!�$�;RW�dH�j���9q��==�!�d��䣕-� ,�<�C�P�r!�ĂD2���@�8CT��vO�g!��ɘC<��Z���&F�"�+��Pc!�;:��"��8æ��w���W!�=��]2Q�ڐ��\�qʍ^S!�$Z�p�����ɺ`�L�ʴi�5	E!�$[� _�}Xp��y�x��V�5T!��<w]�d�����fpq�K��8@!�D��|k�,gğRxl�3���4!򄜰(r�� ��'2n��jI:<!���{��C�E�9>��iG��@�!���8 l�%n�I/��2�X�!��J�X)�Y7!V�S���P�_���DF0I!pe�BҲ4R���ӧ�yr��/m��U�ޫ,���+fM�%�y�	-�Y��G7ٚM��υ�yB�H�'Čr���|�۴O��y""I\�2�^�!��8�a�-�y�� ��y�A[��Hp��$D�yBj��� !3��U��1��oט�y�n�:�;��	�>��e�Լ�Py�eV'�ܕ��έ�����Ut�<aF,���6��d��<a�9��I�d�<�r憰K�6���X�>k�bS��V�<����%���h��J�,��4acF	T�<is�K�����5��݁�d���y�f^����#"UQJz�<I��%�x`�O��3���BS��l�<I���*-L��!�}�B�8���o�<��a���C�L
h����b�NF�<�gӺ5-ع4�ܞa���MWi�<�"(��t���EP����
h�<��E�l���Θ�M�^y��Jg�<A�D-]Zh#! > \V�x'�k�<�g韜$�������!G���@��o�<�d�	�c�f���WiZ�	��IG�<�1!j�٧E��B<6���C�<�̗�{�J�c���?\���%�F�<�VK�j%>��4�����[��AN�<�0�]Fw���3c�H�����^�<��Q3DH>� �lԊ8 c�\]�<	Q�θK�JQaP�߅#�f�6��V�<!0/��dCV(��j\%��T��F�R�<��#2�q;��,yr'�M�< �� NY��]��`�X���I�<qD�\�z�ى�hV-����|�<�F"�: }2�P�2�2A(@ �y�<� �bN�S�FI�"�Џ'�8r�"O�Mp�aۿ[ԱBi��6 7"O������]2��5IOx�VTP�"O�H�5��gp��q�����"O]��B�S�`Lj /�d��-�"O�@pqCF�/+�i���4xنh�"O�����͂:������,6�4}.�!�F�Q���C���0�h��"HS&�!�d 2jՌ����)c��9�HXY�!��V�N��,�5�+tH�{��X5(�!�Ă3�
�pv�UVaP�;$	�|�!�DE�<�@�����i^���fR+w�!��zb:��>bP\�G�3XM!�܆��M����QC�y(P%��X3!�d8$�e�P a�ɨ�֧t�!�Ca�B@2���"��N�}!�d��C��Q�U�=���;e���e!�d�Q6ٺЀQ?=�.:b�E�}!���c$E�@��.!�F[&��$�!�$Fie�m��V��}�T�!�ē/�Vt���e�L(2�f�$R�!�����3�OP��ݪF؊_�!�dԉS�T���b}bZ�1r�"O��B��k�02��'�f�""O t�3J�9M]�Qacnٱ(��!�w"O&�����o����0��Q��*�*O�hPw�z�ސ�4g��}����'kP�G`�o�Z�Rs�q^����'{"�ժ�=Q��.i�j���'ކY�f�͢L�1ĀI�H Y"�'����M6w�i�rJz�8��'�R��jL�j��1j�.V�hr1��'t@�CѦO/B��̸f���$���'XX�eh����(C�D��F���'�i�U3 �L��~` \��'��Y�G�7va2��
tRH��'L��K� ��:�	��l	4�{
�'f8�r�O(H'��X��'��c
�'>�4���>u|�!b� 3�Qq�'����	�-+r�x�O�8�mh�'
�hZ`������ߟ,�J���'������%��:�	X-\\
1x�'	z R-�[�c�+��X^��X�'�f���F0a>��׏T0LG��x	�'�E��̝&BCA�B(:6���'�` Rσ*Z�dI9���:��\!�'�B1SB��/?�eQ�P�DM�لȓ�LX��ʥv�*\���
�/Z$�ȓi�2XQ��M�]]`�9��P�#����bhz=��hA�-D2Qv&��No>�����tA��׃2�Z�!��X醐��v�Zu4M؋IB�Y�ˑ��ȓ5�
��l� w��Qq�HY�v؆�gBP��C;&�.)E
�Xp�M�ȓ	�"�#
�0& 0ځ�ώO6
Ć�}Q>�զ��n�4�ȍ
Qb���G�\es�(	$F[� Á��
˂���b�XK"� �}LL��p��0d5|���?>LA�w�eG�Q�����=�ȓmM�Zdk�+o�СS��%�\�ȓuT�8�7�y)����
H��d��u@��@!-�tx�r$gR�I!x����m ����֨ڰ������$��aN���R ;nx���S�? @� � [�7v�Բd+K�y�F��F"O"�3�H]�'"�)��K#]�5k�"OfHr�狑��l��J���U�"O|�CˀAҵFI��&�ĘY�"OpY�g/c�t��qI��(�T8�"O�ыÈR�Q�L�p�֞b�� 4"Oƥ�en����(�e��G�J1�1"OH����_�R���*˼]3��"O�h6��gI�8*∉� j 83"O�i(��+��袁�I�z���"OJ�K�@�;o����4⚻��퐱"O>��f���)�#�Q'alU�b"O,��ѥ�T�A���ʠ��H�"O,��W"hhq��(��P��"O����_?!��I��d�8ئ"O(\Y��Χb����r�_�$f�Y""O��PS�gi��7d�u����"O�چ�}5�Pr�Z:4Y�r"Ol��&�		����6�*-���"O@Ia�
�m4��I�܊i�N��"O
݁��8�$PP��]�W����"O���U(Q�>/��4��O�F�{�"O�܉�˅�}t�'� @�BH��"O�)��ˍ9I� �edF'_Y��"OB�c��gJ6�	Q��C�tT�r"O��Y$��U�Z:��	�@"O�- & �8�D$�a:��x�r"O�����6H얥:�k�(+��i��"O���$Țg*���ԩ�D�5��"O�0b�ɦW�0x@)��i�(��&"O,��u��<\R���4H�=YpTp�"OL��G,\�ޭ�ǑlLѦ"O�I`ŋ�K���Z�&`9lp�6"O����r�f����4	"$B "Ot���șE���F����@���"OPt��B4hקO�t�:�P�"O�R�,W�3�S�X69�ܴ��"O"���D�v x�g&�f��X��"O�����?gȥ0��@�xuH��"O�y�)�!�ִ�c��6eXAa"O:����_�~A<1�����thN�S�"O܁Y�Vi�1�̷;K���"O�Y��*�=�y��	�.JiC2"Ob� D�U�H�P&�Z�%�|]qw"O}���ad<y��$r��a��"Ob��AW-i�(r�d,5�Z8)�"O�L9�-����a�P�.�x]��"O.�[��� 1�̡�A�"����"O�Uö�υ/�� ³�˛V�|9��"OH�i
I�E(S��:�vl
F"Oİ`�"͜]{�1C���/[���"O HjAB���~�`�f�LK|\��"O\�sU/ɱB6�!2Do�d��g"O (q1�qY8,��-�d�pa��"O�,��F�>��@��Թa/�!j�"O^U�T	�~>L2⡛�" �"O�=���F j*H���[�u�ƴ�g"OF�@��	."~�a6/L�e�,K�"O2�0�O�4'�jΝx0p��"OZ��A��6tsBd��K^�h�"OP�34&S��@31�/�np��"O��9�hG�u 	b����~߮��$"OB�"j �:7�����]*���"Or�Y2k�/s�� nкvxڄҲ"O� �1G�ԦS(��95;!t��W"O��A�J.r�kVkL�Ru�� �"O,,�� �6h&����˼ ]>���"O�E��3&NLӇ��AvT��"O�\����:�%[�*�i6�A�"O�K0�]/uV@�*O�	
�"O�{��vq�O�C�:�+"O`����է-��	� I� ���"OD�y�J�kՐ8R���T�Dd`C"On82�+K�H9潹��	��B��b"O�!�R�$Q��EǺx�h�"OH�#���97̈�f@�'�̐ �"O�I��Ҫe��i	�؜I�n�w"O��sC0,���Wߓb�� #e"O6�1ѡ*a��0Y �ɬ�\��$"O,)��iO���<� ��'���"Oh����Q2(yt<x�	��t�&TqU"O�U'e��(�FTYѧR��P��"O� ���ϓ*M�ī���|�F�ʥ"OD�T��9g��%V�%�B���"O�A'�0L��Y��dD�&sN�a"OH��ƪ�50r��c�\�vb`�"O�!���R�rԸt'uk6�s7"O���!| ��`K:?_��"OFu�C�A��Ђ
E UI�k�"Ot���<T�`[b��=AP�K"O�qs�H��.��Z��*8J8�a"O��Q�䁀?�(���"#�6�
�"O��C!�B�v��P��Z0��'�H�P�K<�n�H�R�S�H��	�'�UzVbXx5�=�ՎN"�ȍ��'� i�r�W\� uip��%C���'Ɛ�y�Ǎ*+aH%�T��92U��']��
1nEf��P9���Gv���'�	dׂ�L�ᩙ`ŀ�J�'�����̮Q��� &��[L����'�h1�e�6�8�j7/[J-����'�ʸ���<]*C��SO�n�{�'�}8PB	�X�P���D�$]q�' �BtAɢ1�*��u��sE�=c�'7�t��C�6a<<�#��s����'�Q0�:$���rȎ�bmS�'t@*&i���q��"����'D� Y��_�I(vx���&{S.�
�'u�P$�ޏH��h@�cO��y
�'	�`V�Y�i���'��1*׼ő�'6U+t&ϹB�@�ag@# 7:���'4�Z�*L#-��8�AB8��9��'�d���Bܤz/,�f�@��D��'ߚ�A�TT�����8�V�����䓓�4��ʓ��D.ʤ	b��
���E�s�!�Dͩk-LI�����9Gm���!�$Z;z�ȇ8v
��w��d"!��&"D�hʓ�O�کI1�N9I�!���B�8!��ֿPub�h�@VBA!��!��ңb�>�rP�Q>'6!�d a�q2G,��Q�Z��7n�Q��y���4MYK4����(�/^��C�I�_fv8Q�'V�+�ЀQ�ܻsbnC䉂(}FT��
�j>���oZ�&f�B�ɏS��a&LvW|��D��xB�	�__��B�T�Xl�QE��CDB�	7O�J�$ǭ?�0p�����J�B�I7l�D���VU.�� gǾE��=a+O"|� :8�o�(?.p1Q*��m&�<�d"OzxKU��9tI��Uh�Y��2"O��Q�7)����A��^�h5"O�Yq��15���T#݀fȶ�W"O:  6�O9x�1�2�� =��9X"O�u��
(�|�RF���k��q1�"O�dH�OF�;�"Y�b��Q"O00±)<&�j�����+5؎��t"Ol�牀.���O?v���Qc"O�4�P��*�g���'����"O"ea6A�U�B�Pr�C�*b-��"O��C\�1V���h�;e�D�W"OB4S�J�"ײ�[��iΐ
5"O�qsP4]!0��%�̕:f�mA�W�0��I��rT��[�x���f��#�B�%X ��Em�Y4���%�i��C�	'@���hpJ0�����]7$ �B�	W��	w �)m���W��-!�B�	�.EB0r�J m��	Ტ��B�0b@Q/Px���P/r|B�I�!B��@C��3y��	��HoٖC䉑_<d� �)��^�)�C��9n˓�0?iU-�> �ȱ�f�a=(p�f���'p�S�<!�A�%d� 1f��]$L��3�ޟ�����.(±)�G�0�[E�<j?"���Y��Rb�D:i���:�*P 6�d|��Ѯ�A�	���L��#Jg��Q��0��tqO��#��m"`
�/OH�E{2�OF�±�8a�>-+�B�"ˤȩ
�'Ȥ�E�?Ԝ!�$�%"Q�9�'�^�8��%&<չ��@�N���'�P��1C�Ola0Ԅ'4xTI�'|�%/�]�~u�,F�>�8[�'����Fi�ft؛k����'!x,C)�*�]�G �:3��T�
�'�� ��\!L�~�"lN83P`�3�'W��4�S(^���E!�1����U�l�'��S�|���M U(5���J�o�0��'l�_�<��m�-09R4T�=�>���AT�<����_v� U�O�Z����.�Z�<) ��l1�us�P�?:�*��@�<��U���PY��$O�2F�Btx��'d BL�*A�HR� �
LC��'��i'Ѐf⽊��Bu�P���?9рRѲv� �c��p3�%�y�!>+N2T8�/�Y���1�抱�yb#[W�r���ąU3��	��y�Ķ	�Y2鞣=电���P2�y�'��X�d��	��I��rM��=��y��9%V�#��Ӳtb�����y�C��V��0�Ñr� ���� ���'}�IzyZ>�ͧ��@��φ�4�Z���N@�f�p���e<I�'�yB,mar�̘���r��Z�<iS�N$W����!N�H��L�&��P�<�7�T��bpɡ�U�yd���$L�<�у7;�
P媖
�ʙ a��I�<Q�	�8�H"���U��{���I�<�T��;:�Y�&GBZЋg%|�<Q1�V��H�`��	_��Pۣ,B̟P��c����b�٥jyP�!'���'�%D��p��_6t�vy(��@�W��Z�'D�Pkg+ڊslμ�� 
V����-$D�Xh��&���Ō���)�Ì%D��aT
sJ�����#�p���>D�� ja��KV�C�8�"��(*�Z�1u�	}y�Z��Χ/ö:e��=-!� &��	�r����d��ɖ�ؼ���D�G�n	{@K��EW�C䉏7:��P�^�xtz���C�iaEc	4�ؤ[�C�/O�����"O��1嚤w��I�L�?n9ط�'��	r~�L�!^���@�ӡZb���I"�C�	8q�H��ALG�&'Py"�aY�c��C�?>�} �$�9a�$!�։k�`C�	$1|ղW���S�3��ҭ@8C�	$k�(U�QƗ�{���hP�&C�I�k�����L�P��)%�C�ɬbH@0�4)ݔT��� ��K�)�2B�I$fpH� �C��y#���K�*B�I�&b:%AqO�(�I)�n-�L�ܕ'��`�'c�hx�!ɗ/0~~�'㝂[L��IT<9�9q��
+ğK�<�A��i�<�Ùy�f�kq Z	:^1��i�^�<�5*�,�Fm�w�ڜ^��y+�FKX�<�+ղ!��ag��O$��:��Q�<q!� �B�ƥ��.Z�z*�U�0'�B���͓H���pe�?{�
����B�B��ȓ��+rC�%\��O�N�.��ȓ�9Y�Ƶj�u�螁�����	L\�L��HD.@{��˱����,��P��6H�Њ�HO5Vϊ��ȓ�R}Q��T�\�'�*q�����r. �����x�"W$�-O��]�ȓvB^�s@�SD6�h*�`Q�E҉�ȓ|�p�`%FB�:�����P+!Hu��{��4�Ƞ�$u��$TY�|��I�N��7��W�<q�dL �L��+E��2��*�ǙZY����T[XC�E��V�1�S�&,�ȓdL�rb�� q��[e��/K�5��n@����nۓI��
^�b�؜��X�8qkL4b@�	��?\	V͇ȓ2~D�2)�)LfX�s�Sj|�ȓ��I����d=�(cc@�8��e��qĈ�FZ3%�� B��J��"O��j�C��2�`xP�L�1���Hs"O�iE b��#$�䡙ӬH>7!�DS 0dt�2�*r��1si^*�!��H���0�˜$J=��;�%\�XY!�ӑo0΍��/ȧ��}��gJ�>!����%ZL��T[6E���T$!�䊰(b0Xf!�+k>�x�T��A!�$�,MAH%���K91%��ω�P!��ѲSt�9�$\ ,"��N�S"!�Y�ü�c�I�Q $��G�1!��]�Ê 	&�Ā{� e)�`�
6�!�$�:����듁g�`x)5��
8�!���i��ITM��	��ʎ_�!�dܭK&��gܒY@�m�M�&w���
���훑�,c�9�y�A�o/�()"��a����yB��x��53��E*
�@\ ���y��^;lz��F#�Q�ZT"�,��y" \''"�����1�h	����8�y���,	4�*V�^�/���I�Mޮ�ybgӞ7�>�9@�^..�F�P!݈�y2B�E8�чOYH���O��ybm��IlƩp�JSE��} ��@/�y2!_:P����d����x�����y
� $R6Hͳs��<Kd! g�!�0"O����cD��,����U�L�@�"O$�a�L��!|�E��o��\��[�"O�M���S����ӖhСnL)�&"O�u2�B�Wz@U�4��%>w	+3"O��1�F[�9j���4ɓ�0 � 0"O��*�h� �H�i�%Q?%�D�@"O�h��J׉��8:&ʔ'�h��"OL�r�$fF�t���}��	�"O-3���at홓0Ƥ��"O^�k�	�'%��+_;��;'"O@8qs��/|��(C�)��q"O����ľ2K����c�:��"O�\)w�Ҡo\��J�m[��!�D�5o "���q�<İ��� {!�d��q�Z���$���v�ͭ4R!�Ԫ[yV��`	2�Fp���\�JD!��J30$��XƉS�H�lk⏖�.�!�D�R��q�ς�`� ���/ڦw^!��^& �ځ+P܆�����!��D�hq!@%�b%�nԋ3�!�D�S�rA�s�(p�X���@'Z�!�$S��Ԉ��ƆR�ƅ*�N�-H!�DɅ�}�q�W7@��1��G�'G!�$%Gp8�@��Q�����A!�ܗY�����O�;PdF����=KM!��B�7��[kQ�j,���d�r#!��F���@V��D�mp�G�.�!򄔉���:ԁ0Y�X�}0!�P�K�v�pe�.8�t�'�A(A!���`X��ұ�Q���Z���
0m!�d�rm�\3@N�����P�+�Py�I� >�05m�6=!���!Y��y�#H$T�9K�,O61��2cV��y�ŋ�;=t��ЄÒ*��rbOI<�y�e� u�z1*��-�QX"L��yRM�yT�ٸ�a�i�5��yr$_u
|�B���u���u��(�y�*�o0LE`t�'�PP��(�6�yB"T)�d���=3�ɰD��y"�ÕW���ZS�
3��q��L��y��H7H�$�7�;1(:�ӡ�ڛ�y�"��UN��CA�֗+�ҙ��j���y�0xp�܋UO@25��ȫ�J��y��	��Y�V��&�NX��lZ��y� ��M���/I�ބA3��(RW���ȓ`�`�0i��l�n|����2
�̆ȓ�>�#AH�N/n���f�~��}��f�` 霊S�~d�7*�7�rńȓ6��!W"�B���[�C��"��ȓ;P�FMƑCU���4@/�y�ȓ�:��
�"Hi�a�W$�����R� 9sb F�\��%��N�T��W�ңM�����E�z�����B(��2.@��J���G�9kgXC��3w�ּ�@�ƹ 2<��1@Y.C�I�=��m+����&�4)�1���~��B��#���nځ5���k�B��bz!��|��4��`��vة�Cǎ�!�d�)�)��Ĥ��ȥ� -�!�D�X�.(F��'�v�)�#��,V!�$L�T��3�Bٕ3N
]8�9B!�$LB��8v(?[�B�j�m�+0Y!�dޣ!w*2���w��]�Ď:z>!�� ��x�	ư%x�-� �4<2�"O�chZKM.e�,ߊ(}h���"O�A���Z�l���%f��"O�1ICM���p��*	<VLb�c"O-	!dʲ�^��f�Ȥw�2��"O(��c쀥h_M�t�� '���"O�z���C'�8���)-,Hg"O�� �%�Ft�{��m	x��"O@	+�(�&�d٥�U-L_V �"OhL�⣀j��J���l��Yk"O �c$�ˏ>�y	��S~}�M q"O���G���P���Q�p 8�"O�A� �;U������K�:��k@"O�``��J�<��R��2}}إ��"O��2'�M$�Pppϋ�p��9�"Ox1�e��0��%q�S"/h�p��"O�4����Q���
"PL�0!"O����/8�*!;�HQ-@0�a"Oȳs/���m��´��"O,MI�M
FV�����"�0�1"OV��RI-y��̨ o٦S
���W"OD	Q�-֦T����N�^b�Ç"O�e��F-/V@iB�Y�Bp1�S"OK�.��jd|D�ŅN*&�}kA"O|����#I��:���Xĝ��"O�Y
4
B%a� '"է4�����"O�YAR�֑Q��� �����۶"O8Y,5�*�U��4w�D��ְ�y��`�f0�%��k_�a�`�ӧ�y�@��#.�(��Ba%��M��y�l1$/L� O�]T�}D�[�y�h_�$LٸDgȶSv��j�O�y2��
J�P��F��_0<�h$�yR�� ��PC0oV (��|{Vm���y�LCu*��g�)%���`o���y���'bJ}��p�h�@ţ��y"���CsΙaDпl8�4A�H��y����\�y�����4���yr%+/��:�!G 6���T/]&�y����i۲pf�B��B���yr&-�������7/HJ�4�]��y��УZ�B�CU�T�����ϓ'�y�ھN$$����Q��p�ī�y�aVct� 4D��=!��B�:�yb!S/t1s��?c�����!�y�$ӜcFF��P�G�F;D=� d�y2���>!��Òrj�1c�X��y�a�!��<H��E3n6�US��� �y""N$�6X�dkf���c����yb鉊Kڠy�@F'&�}�êӏ�yBi�&&�����$GZ}�SK���yRBC*w{Z�9�S!4z��i�,�<�y"4AZu�!K��.�Dbcaآ�y��ԛ>�nD�"0^�
@/˴�yR�ܗ9������^�%�(ѣ�����yB��9��zBlC.V�H����y�1*������Qp�#��y��FRvN��΃�h݁��ߘ�y��m���1th�}|1�fc��y�D�	r��P�zO��Cf��y� ��}Vt�4σ�tfڌ+7&�:�y���
?ڲt��Lr�R�R�'�y"��@0:5�X�[3�Y�Ȭ�y��FƎ�P��P���Ir�[?�y
� aʴ���w�vA����A��Aa"OڽfK:��TB�G3
�MC�"O���f�2=,M�MK�i�4���"O@��A9Z�u  �� t7����"OVp�``��`�p�*��H"��u"O��j�!��K�:uk@h�>y2t�0"O���� vƒi����[O��"O��s�ܗgT�t�T�Fn��j�"O�(�NJ�5�	�eҩ[kfy�T"Ot���P��DP�G�/J�X�ڂ"O�4;�_����c G1EYP�"O��@%�,Ð����f]��T"O`�+DI�T'��Ha̤'�<��"OXI����:;�4���<�8�( "O�p{"f��Lb��Q���i1�"OF���fF�:mB 벬V/(&<9!"O:��Ƥ	&u�M��K "��"O�B��H�,���ϥ�0`�0D�2� D"c�L�7�O&y�&�� �"D� ����V�,��g����)4D�|ӀUTp�9!��|.���0D��4�	��J�" 	�$
�)F�-D�آ�N�X�"�;1�M
4��$�+D�,����;CD��G�M�^��e���(D��ss�H�@�z5��K`�Y+�1D��+��Q
H�q�H��L��V,:D��)���5{*��U��w�:`D8D���@E�u������N@2ȸ�+*D��HI��h�1 kH,G} ��$D�������1��pSd�Q�{�d!R�"D��c��		P\��Εh�P<�U�!D��x�׊:��E���P�F�(@�?D�tqܼ!M % 1)�~��j�b=D�, CK!���FJ��=]��⣊<D��
2��r6P��������L�r�8D���,PA��S5a�o��܂7�7D�l����_�t�0�� * l�x4�4D��5���Fu�U�E�i�EE4D��x��t���IxS:]H��g�<�Ge@-BPvq���+Mm���RC`�<QR��h�ƩA1�ی.b�E#Z�<��g+
܊�Y��]�MDn8���U�<9�+;O:Ըr��:e"��1�S�<1'�XƆ���]�`;j��1�X�<�Vf�I���K�E�O�Q�<�$A2}�đ� ��N^�h�c�<�U�n�r9P��( ��h��z�<-5*�yB	��!��:	�lB�I#Cj2d'[��������{�JB�ɛt�X�����P~ԍ��D[�1l�C�`/�ͱ@�M"E��BAGU�|C�I�>,�4�C�N���0���u�B�I !���·7q��Zo��-Y�B�I$KmzM��B�	���G�j�&C�8Q�x�A���˘5q1�q�C䉯2x�!�ԊN�?\vыg �j�B�I%E�j�̔)DnE ���VC䉉]�lL�dI&g�(ʷ�V aVVC䉜K�,����� ݠ%Rr���lVC�ɓb:�;f�S#�Ms�m�}�@C��"�����)��Iғ��C+�B�I$j���"��U��9!���i�B䉮��1	3NA=(���9���d|vB�1h�Jp���GR��%⛝-�FB�)� l��	�8�( ���,��e"Ory��c�m�����N�h�.x��"OЕj���:Y��L
&BV�U�$9�3"Ot��N�]���1G�I�2��3�"O�5!�`Md�8sG#�) �4M3�"O�-���h�`]z�5��uKR"O�H{��O�S����֢�4>d͘$"O�q�I�C�h�:��	907���w"O���wm�f��db7�B�y2��V"O
�+A'Ă��E�7ʗ�?s��!�"O����ĉ���!��̨@[6B"O��+ #0�h5�q��qL����"O>��t��y(dp1a&{�2H˱"OfJ� ��D����T�1��ٕ"O�9�b���fR
���%3H����"OD�(p�M&	�|�ِ��,>:V�0�"OHi��P@��2f�E�&�1�"O4��v ��5X֠
%c	��e��"O΄8�LޕA��!"T�C�M0"O �+rH�Di���`�<\�9�U"O�YP0��"5R� b�Aύ*{�}xf"O��JK�;ƙ��-b��@�"OV�#D`ܑ\��uX�-83U�;�"O�� 0YZB�{�mZ�D�-�7"OY�G�@�+��1
`��F�ၓ"OJ���)[�?\rٳ��Y�sa"O���-ŁŨl��[�u�(]��"O��(UK�b��Sף^�m��@0�"O�����(z��qu��	KG�I��"O�����ZU"$L�7�W-����"O���d c�]K���
�~�ځ"O�y�$��4���;��3���� "OD�:��_C*�Hyth�����:�"O��c��:�*h��GB2c���Q"O��*�;h��1Ħ�2E�zAq$"OL1��P6k�l5 ���]�:��w"OV���&ǔ&�XKva]�>��"O�1��E'�R@��oL-� "OА���ȼad�t����>YB���"On�4��h�4ty�U=D��Eq4"O ���(M��E���	
l�~i��"O��ң��<�w�L1����"O����4�L5 B$hx�c�"O����-ºU"�P(�C��fp���"O��b%�=o���'h)�d(D���a�4fH��c��ę����d%D�|˰�ț%!�:�J�E�� ��$D��k¤�})Pš� �����v�=D��q�i�7p
̱��[4l���V�8D� 3BjA�`��`��#X�c|�8K27D���5�F���iq��V>@yh��4-5D���%�P�)i��U� �@�bAC7D�����Z���B�@X'F&=밭4D�� ��(vX��$��l�=	V >D�"U �1>�<��!,Ǫ2�挀��<D�8�Vk�/n�p����e`���'�=D�죅kU�o�B�p���v�Z���-D��Yq��3fQ� �h��@���+D�lz��\5x,d�I���mpp�q��)D��k��\��؍���3"�
�.2D��0S�c�����W�}_ޭz�*O@ѱPl�(ZzL	�v�E�@6��"O\��t/�1�j��t��=F^pA�"O�}u
�$O��a�5�:�ؘ۷"O� �\���a.p0�	oК���"O&���aA�P��{�"��I�"O�d	BdÑ=�\$p�L��\��"O�A�
�B�0��B7+�����"O�P�HF�9�}���9R�z�HQ"O��#֏�+[L��kS䚀x_B�f"O�[2k =�Z���I2P�t$��"OHP̉0hy{���Ѩ�:�"OF2.��,���"D�q)�(1"OL��]�n�B���B2uFXYv"Oj�z�'JyD�0�@�S���:�"O���6�,tѢ�*Sΐ
9��1(�"O�t��
/������=,ʾ}K�"OB�a��n0���肔5��Ii�"O���d�U�+Ȇ!Yv���$ؖ�G"O �3�<~��y���,-�\)�w"O:T7�߭yS�1yTe�/��}bD"Or���OK
+��t�@J��A��Y��"O�vg�+2�,��$�ж"O��p�Q�_� ���
�B����"Oމ�����'aTȘ�=7�$�"O*9���b�(���5����5"O:%3�Kߥ\�\P���:;���"OB�Z���RS��a�DI<WoD��'��?�fHS�ʝ�p@3��(g�!��X�pP��K'J�~���
�_���2�O���w�n���!$M]���p��"O����	Z%��rk�k���(�"O�Z��ӾC�X��a�FE��%��"OD��f ̀%Ġ���j 0"O�|t�\
nD@�Z�_ ��"O��t� $CF$K�Q�fِ�"O��S/� x��M����4� "O��ũ����4� )�_���Y�"O���*S�28�𧒼M�Dh�"O�4�T�SY��ąR5j)�!��"O�eł��	�m�E (޵R "O���+C'�,cq��^��!"OBLKǉ�>+��p��,ܬ.�:�R�"O0��OKg��p��ʑ=K�R��"O�U�7�OfJ\��*�1�|��r"O���JH8�\���q���3V"OX|�w"����ԇJi�t��"Opl���g� ��v�K���)f"O������+nY��u&W06��Y�v"O@�2�B��K�xx���a�t�jP"O"��d��!JVY��R�]�r���"O�L��AN-<2 �dC�2u2��t"O8X30�=��d�D `B�I��"O�Lz`��=��5���ܞ;�k*O�p�mA�S���4/��v���'SX�(�d*e(�t�۲��!��'���Z�d]�]��M�s������'��I��!/���R�pJF�y�'������ք��'~;���'���% �<�q���#oR y�'|B=;��AX�y��G(`��'�;T��,#PYq���X`��'�"ỳ!�]Ԓ鰓(���c�'��8	V#��i�0HS�/
�v�i��'�aJ%�¬j^�X#o�:#�Er�'��=�%�B�jLu�l��{����'�8UJJ(�j�S��rƜx�'�N퓃�۲sAK��*iH������ ޴���*Q�`sFB�%ז�ң"O4�ӱJ/q������Z9b��"��N8�QWE��|�2a�#=�
pBJ?D��IӦI1����2
�"D��k��:>�I�gL�4�P=1�5D�@��%��thP�Y�V�h����e5D� E�3��,��`��e4��&9D�,��΄�<A�e* 2?J�hi6H8D�d�f� �BF_�0�0��^
^bLC�6,`0PS)\ h�J�"� �<��ȓ9\Ղ5
C3$�2��n��
m��7G��)S�'(��Y11	�?Z���2�.	�A���%b��4 :
�e�ȓT�V�t�W(>BRD3���d@��U� rDN�<%��EGO�:M�ȓ����r�M&O�� ��Y�L��!�u�p��l��%���A� ����ȓ"Î�Aaӑ��لHFi���� ������K0ٚɈ5���ȓƖ��󎆊r����Hҝ����� &L��%�U|h1Ţ��L�ȓ���q��BR"(���ДD�& ��n�F�yA� �4�0 E҈:�>UEz"�'�ܼ��b�;>a��ƪ�	�'_�p�g!�0tjf�MOV�8��'&(�rlɆ{�&\w)ٳx�!�	�'��5��Fk�A���C�H��'^v��C�&j`� ��(:�$�k�'^u��l@AN��I���5D�=��'�
��̔?`��#��'�fL��'�����~-�Q�sC��a�'�vIɰF��.[h �cN�/$����'*ȵ��J���f$��)n���'�4ڶ�^�pZPl�%FI�/����|H�C�A�2�P��ń{�цȓ�(`9���@}�x�Sc�[���ȓ\ު�x�� U>�u�7+Q�&����|�a����DH�# �]�f�`<�ȓ7'�5�e�87�� *�E=��x�ȓ^k��wD
�&[vTsbH7�	��`\�p ���4rv�c��W"��s�6���#=2���@�Ru)�ȓs���3� f[ ,��ޖT����ȓyF���÷?�|A�B"�)X�h�� l�����\����iL\<��w�$�&oZ��Z�ؑ}�!�ȓg|���Ț,�<���=�<�ȓ1\��0�Dc� i;g���u�ȓ8����3��3O���_�]�N���QBͫB�L@TH�e�p����&P&!��N�%l����a��? �=�ȓx��Ȫ��O�?�,�U!)C� ��|JV��D�U�����>B0Ї�#nT�%��A�����S;A|f����d�SII3)𝱕C�3�|��HHT0zp�W$2Zx�hq@@�I>��ȓQ��}�L�h*.��.B�U����'<���aN	�@ln1k�LÏt| L�ȓ~t>�B�K�{��+��N�5~L��ȓP�B����<�L���!�����Q��X7&�^�t5���G0�����^�T��B�j��.�Q:4�� On����ӥyn�Hx�F�4졅��@�Y��͛�&@c ˤ>;|���S�? 8�S�g�&���APX�yӀ"O�� %A{�F8X2Qx*O��n��4���f�#.=Z�';
pZe�9U,�#���/n*��'4&�z�,��b�B���Ɨ&N]B�'p�e�$��;-�Q{$�/!4�[�'�4���
�WF��w䅧��}*�'��04��	�����q�\8�ȓ=���N��A���c$�Z������#��C&��O�l4�TFЁH���ȓ>���p��Ň�zy#����>������z%�"�J��D��;w�H�ȓX��h��V�Q����!һx�T�ȓP�B�����bw	���L�H���-6
�+��|����I����ȓT�	q�E�)�\��eM�f=�ȓ�L��/?Z�	L�d���,Thhĩ��6Ȗ,!R��V�����B\q����N��ǹP��H�ȓ(��)�ơ*鬁�BEP�$�$t�ȓ/B�L7��1N.���dV�d�v̅�
%ؑ��nG
NјYSŭ�y�}�ȓӼ]�!��K����P�Z=g���F��sT#F5G@E�lS}���ȓbD�Ib��\�*T(�h�N$�Ѧ#����.�"E�|��I�d�t]�u��������q�B�ɷ ۘ���'"��� �K�S�ZB�ɂbDȢ���|D�R��=InB�I-�P�I���v�Z�hf��C�	H9������Tx�8B���nV�C�IoY��R��(	)<$Z�E@�[$C�I�?��yYcCH<=�<�Y!k�qC�	�?�բ�͐�0�A�"Ü7�B�I�GA��rq�[�;8�Ѱ��91��B�	�;�(	`��Rn��;�lC��l �����L��T���0c
VC�	�e�%�C펪fhJ��V��%:�TB䉑��JAF{l0U!�'�tC�*T �����k�&$� k��i�B�	�G��C�.�|��"�$C0pB�ɏ
)��vQ���գ֨%grB�	")��a͝.��� ͛cf�C�	�gNd��bM�@� ���o&C�ɻ��u��ҭ�>�'�����C�	�Kz��G�	$i�u	"���=��C�	&K���T�B��;RFL�Lb�C�	�v3�40w�ŘA���]uQ�8D��RGa8V�љV�̭E���8D�6�ܻ�J
f��>]�u��`�m�<��#�m�,9�6-�9N�z���k�<A�I�=�����4&�Jq��g�<��"\/x�tQs�.W?Yz�Ѥ�LV�<�(�5F�8Qɣ��8R4��G�W�<�F	�;o��%e�3~��}1B��S�<�#d�B��)
.X�o\|�#˗K�<��eـ3d^5@Ԯ�"�z�Xw�_~�<�fK�9%����儡S�&���B}�<�B�!"�$�g�""2%�5̎S�<�nC�T�	�N"��k�H�<��Ox�����Fk!�%<(5:1�ȓk���S�%�'U�������ā��W�Ld��"�&f�����J9!��f\X��!�2y��=���3)V��ȓ~^LQ E^��Ӂ��e�}��S�? �� ���?Y�
�僠�	��"O�}iE���S���̣\�9�"O��CۘS�4��%"N�L+j-�R"O<�	u�	\�r�Br��4aB���"O8w�	�L�����O���x%"O�I G'_nZ��mħ<يiy�"O��#�#�Uk.�`g��^|���S"Ob��"aԖ�q��:c�$a�P�T��ɗm�4+����S���7�O�����8?A�'��[�r���AR�u�dbKV�<9!�\�'�8�Za̭ ��2ÂQ�'Ga���Z����1�ȭ"�}b�J͸�yr��L�⥲!�&G���Ģ̓�?����S&6�n��KH���:�r`�ȓ7�%��i׶KB�k��Q�إ�ȓ&��z�㈥d��@o��
�h�ȓc���f�F2!��X2�d���͇�&��-� �$7ʌj����Vهȓc�\��D��y���c,߃|̴�ȓ;|�񐦯�Jt0��!��s�Շ�o��<�Ӆ�Io���l�1b�$��$�X9�ᒞGb>�Ơ�
&���C˞�ٔ ��ZC���F��r �ȓux��z����Xi��.;y�,�� ��@*�q�\�(a`��E:`]�ȓw1���FP��,���#Y�";dL��,�؈�ƟD{�!p�'Hd����ȓ<3a��E�	jQy���q�P����xyB��a89�bl�.ҥ�b@<�yB(��
�xk�e��Z3�^��y�CQ�p�<��&蓴&b��A
ԣ�y� I:Z�D��qN�?��ʆ��y�B[,4V��ʋ�q(���Ɖ�y2j��?�x��`�		�|\�E��9�y�	Af�܁&C��y־=�ӫ;�yB-ȿp�P�]��8U��Β.�yB�-��AGQ<nh��1̗��y�׫@��ݭ$5�h �##0�C�ɴ+<�x�#����qc7�E�R�C�	mbD�P�IJ�|�ր���@!QդC�e����7�� th�I4D�;,˂C䉡~֦]���HL�.W��C�I�d*�hp��rPL�w��C䉻(�虊������*GJ�(e�C�IZ��U@�"׎.��y� L5m�JC�	$J6����@ C��sF�2@f4C�� �&�T
�1ӄl���'��B�	8V����v:z�g�T%C䉒��\���B�r ���7(i�B�	�+%"D�c������c(P�G�C�I�v�	��DY>B 1O1�B�	�t��@�����B�N&%�ts�l!D���d��,Q��3�D$ِ?D�X���A߮TXR患g\�r�.+D�<Buc��/��3e
�$H=p�%�)D�@K���vEy�I�j���EE$�O��OK���Ov���f��,�Qw"O�s� �5��$h�ER y�����\���)�1e1J]�w���#�X�yP돵9!�d�2DN��#K
5#rHLv�L��D8��_쓭�O|�Y�`X�2� ��E:�²�'�v�R��F�d�4g � >_���i��~��!�O�d��'ү�&8�@��������M������{Җ��B�77��4+̉HH�6����y
� �EK�
<g�|H3'Ȋ2P�� 1r���'t�4���<��ռ"�����KۋM��}W@ z�<!dg�'Ua:#��#�2��D���Cq� "E0�O:ё4n�3�!J����'b����"�e�� �i
�N�:,4�y��
@ !�D>du�E�'�ɱS�]*$ː;qO*�U�"�)�I��^+�aK�P�Nq#���!�D��`Z�@�Cܬq=��x���E�!���}��@	R��b�6i"��(�!��u��9(w�â,�����T�1�!�D�/�Z}�A@eP�Ӂf͖�!��_	rF�^�f`��_#H�!��2�VXaG6墀�.�"[���*�S�O��E)P(Z_kH��T!o$�{�'�Y%K�0� ����h�f	
�'��P�o�!i[�(;t L)d4T�	�C��Rf����XvƏ�h��D'ҶFb ���\��yrK��$,p�q�NL86�0��C�ø'RM� J!Z!")y��+tc���ȡ��:VXd���"0����&"O�88 ��#+�\��/N5Lr�p���J��2(���5x��\�$'�7M�>�:�:uB5���LVa�d�&��l��N�,�ip�1Z3�4�Î<��e�g��è�e��E8���m��0<	5���Rj��-�W�QX��)�j�-=jmk�oB!��5��Ɏh��Q��A
zx��3%�#y�䘶�'P�$9�ܞ�� �w�M+��h�N�t䏎�Sni�v�J'�N��a�A��%>�0�C`�1�"b�KJ9D�|�	*JT����^;�ltp��[�m����ġ��8<�E����j�c>Q���Fk���Y��p���,>��Q��EQ�4�!���X�p�V��5�0P` ��q<�9��뗰iCAS�(�)�C�2x�x�����%#��/@�evІ�}�џ�h��=c�e��`Z��bgE	 IĽBQ(N=Z�X��	�k(<E2��ܪ��Ї�ɂ�`��ꌕrL��R�GD�I�@�3T�!�B��4QS`G6ch�ze\�.���ɟ�LZ�/V�hz���0��O��0`"O(�Kr��������)8�p��ÿ!\�- pʉ���1��C�e��O��-���щd��6u!"�YsBV��XQ�V&[����7w$���U�ӕ �����O#k+�^���rC����U�1^t�E-,��O���
��x�a�}�Mr���)/:<z���/k_��s�i?)�V�x'�*t5�@ϒU�l�CA��w��j��I���C�a@M�,����H�$���ɦ��<���^/ 6�T[�G� �IpP!R�O ��B��7��	�,<dã���6%�y S����!��ţ���`k�� L���q�}�Jjq��	�n�[r���,����ܞ��<��?O�=��.-,�A�Ã0+�h�{��'H�-��N�9I��p `
~��&���%�@!^^xP��9��}[gn��� ��{�Z��i�y8��(�
-�B��%�%�}���C@�,�.�jN�?bL(	�K�{�d�	ނ$�zyJ1�ϙ �L��Ǐ�'Zў��D�'��(�O�;1%L�瞚[��ɼ�̀@i��~`x�Jb�- xᓀ������O2� 䁰z�T��׫X�=˼�R�'ў�}��Ϙ(���a ���w
�o����,ɖz��@�#ۇu��ڦ�!�)v���a�Q�	����%cڢG��x��ȼ����n���+��S�8��Z@�D�;\ Ȃ�d�yI�p3��]�-Z��cE.mE6٨�DJ6>���=q�O&q#�Ď,f]@�Y%G5(>�D@��	:��e)��u���F��h����/1n�d��g\�oj|`u�B�w���"�f�6�㞔E{��O�#�$I� ����/V?F��'�r���\�p��qI u����D)!{�����SAɢ:�t�Z&�@J���Å�O�=E�TH�v� ԣ ��f��h��-��qX�퀼	w�h� &��v�"�B���U��Ӈ3ed��4A���� *Z���o��Qn��V� �hr���4*Ǯ��v�R䣣���A�l1��C�q��tRg�ſ8�LԀ�V�'{�	��/[�[&�J�FJ��˓_��+��H$��*ɏ9%|�̓��ha��*\�Q�5G�N�����@$P��Sd�<A1�Ūn)�K>9"�*j9��R){�9*w剔��OV
�Z�)�`���Tʊ0�����'�j�rGf��+����� �
���Ɇ(u`�h��-Ms����������S�T��Qc0��*�oM7( ��a�aU�^����!F��s��`��i���j�nj�H߱&Tf��-����)� $��=�fR�ʴf%��'i�H��!�"A� �
�&F�i�@�Ӥ-Ƌ]��5��ؾ:R!��1p�Ԡr���T�i���!\!�$т!]|H1p�ʦx�
A�Ed��	G!�D�;>�
�R����po�� `L[!�d
�@SaN�J<��s*X�[!��#iPܔp��� ���!N N.!�$	34��T�����6kь�2<0!��F�h#AX$rɌ4p7�~�!�Vk���f�&�@�����i�!� �F4$�bʆ=:�԰I�f
��!�Ğ�tI�%��@�tH�$eP�q�!�D��p&`I��� )�$ ���C�!򤗐	D�p cI��5wd����'�!��\�M�T3"@�7}��i�H��!�d�%l��m��U#c$%��->1�!��ݝ=0�t����� �@A+4"��5�!�d�9�TY���;k�8��@�v�!�W�-�ԪF�D���u{�L(�!��+L�8��J>�­i@�Z�f�!�ċ����z���"�D���띒_�!�˻\��k�<j�T��I�P%!�զ�DX'����|8҈ �M!��ƺ^h�hp�DZ�A�&��Ç+l>!�Ե6}�lYЈA�3�����I�<M!�D�3�L}�%ḠR��t�V�m�!�d�L�fȑ+��J��}˃+(�!�ݔM�f���ɿo��T�P ��
!��.i֜�+˗kڶ�`M��
�!�D��l��\i�]>*(��[rc��!�ěf6�����-��PB�&D�!�D<.�Y��A��н���;�!�$	`��GIK�x>>]aPfʧv!�ޫH�&)���/+�����I�!� $���b�ϓ2
j~8�!-�7<�!�D��<�,�"Ƃ�i����U�#�!��X4`!�)�3 V4]Vҭ�t���N!�D\@$��� 
��>�)�B�&?�!��'Rd�l 6�ɂ� �]:�!�^(y�Q�L�W՞b��E�	�!�\+/Ɋ�"sa�(�
����4M�!�䖑QY��iE<J�^�h�L��K!�d����i���D��q����!�4o�eb'��SՂ������>�!��i�H�@{.p�aGC�!�d�� cL� R��٧�ʎ�!�۟f�Y[s�S"%;h��'1!�D�2r��x��C�[��d`1�+h�!��&.� ����HH8�e�ţ*�!��� ��@:e,^���s$QT�!�D�?1A�(	��5�������9]!��C�?

YҡA��=~T�@"��!�r�ȡB5�3}m�U��Z��!��(3�>];B�.B�R\��Κ�xs!�(|#��@#�+j�l|�E
�''O!����@,bs%��T�IBۨ-5!���U
ȉ �/8s�S�F6z�!�DI�*��q�7�$~\��A, \�!�=H��� ���"07fX��G6V�!�D�+�-���S+bͪ2n`h!��D�8Pi�N� ��i(�m�pB!�B2sEi�7�0h̬
�Ąn0!��!d����DaF�f��KF�YW!������ᖜv��� `)�]�!�� }�Ǫf�����	B�A���!�"Op�XƩг;�j�!Q"��c�+�"O��ceo�5Q�b)���%�x�U"O�@�ܼ�^����-B��Is�"OPzV�B�?���1��͙N4d�%"O^�aqPg�n���/�~6j�as"O�h�͉�tc�e���";�t�D"O����Xt���)X�1��M��"Or��%�L@��B�C:9|H�"O �9��DVl8s�	*Uuԍ�"O���&��2�^4[D�jԱ[�"O�� ��Z�f��)�AG�@Ft,i�"OJ,���ԖY80�sw돈=P�h�S"O��tg��E�^�x1��+}�"O�}�V�W3Dti�Ł2x�`�"O�`������#�%M�$벝*�"O:�j��7o�D�X�E�0�����"O�p�.@*�,����F�'�(<xA"OZ��V�Һc�p`�Qb�=H�lU�"O�p�_,b��#�R% ��(! "O�Z��$$*�������Q+�y��۬Z�z�6ET�H���)qG���yB�$L ��i�F����`&Ͱ�y�=-A�MYԈ�/�`��O���y�mv����y�(#@��y2υ�D��1���B=u"��zpA	&�y�m��#�le�m��<`dJY��y�֝T획j�;e����S ���yr�[�,�b���K��imDQ�JY��y���[\��K�1r��q�Ŕ3�y�i��\R���q TyK��G��yrNף%�j-Riأ�^��5G1(B�I�
�<5�ԤK"P��8�'>UlB�s(��a�R�t��9� #[,�B䉝L�n��1�*׶�Fo�E�RC�	�ct���A�74~e��/A�'�*C�	�O�ձ�eZ9�4�F�J��C䉣���2�A^�$��j0�_%]�B�	*��▫$�0�)�I�a5D��PT,y��)h�"��V�Fq�1a0D�@�����y�M*���oF����1D�ԁ��t�Z-�6�B� �NM�@#D��/�.��NP�!������!g�!�E�^����	"E�1`o
�<�!��&_dhQөZ��ce�P�:�!�%�&��Ԁ;_`}�w�K�!������_�-�`�۠OC-\�!�$�	,��s6�	3�8���#O�!�_kd5��è&�p9�2��)�!���$!XRQ�� �+^� #`�ʁ�!�M�3;�l�L�d�xXh�iE�g�!�ʔ$��L��~��\
6-��!�d�B��k2m�x	�"��Rw!���.�3�K=F��`�N=+�!���3}�|���T]vt�Sҁ�&+c!�䖬E�d��
<�܄��O�0	
!��6\�Ej�N �8��w���8�!��L�F�SW��'}���F)T�~y!�D�TE6Q���XbA��i��4F!��� �P����W9?U:�	�\!��I�!�͊,՝-Crt���M5�!���P�&GJUM����#
!��oa�oʼI���e�0
��&"OT��H��5�T��q�>���B"O� �ЛDeԠ3�hŀ�F�
	�"O$̑d��[�v�jT�Ӟm����"O¼�s�ݭbp�
�a�{��=S"O<��BDϸx��G K�B� ��7"Ol<R��;Z6��@Jm�rI�"O�W�"cp���սpQ���Q
Hr�<��3r��+�,E0UZ�J��o�<Y�$�P���GA1*A��J��e�<9,#>f��K�ʒ��N�<!q%
P�0(5MA+%�� ��~�<1BgҩO<~��-[;�I#s�Qz�<'. �E��$�ǥ�6`>��M�<ID�S�p@ڽ�`�8�h� ��P�<�f��?@42p��� TR�J���R�<�/�)]�6�X��8j��
0ǒe�<���οI8��+�;	n���e#�b�<w,L?TD�AF>C�x����K�<9C�]%w��|y1��>8�F����C�<���?h�t"�+��^s�9�#�{�<1�[=lh����հ��Zƍt�<�#�&3b�ɦf����H"p�St�<���v��q����|Ir4�+s�<�0S�
+ȅq�(
�i�N��0�V�<QR!4l���#�EX�W$�̑D��e�<����:kf���`C�S{vĀ��J�<ᰊ��Qz A{,�Ц�S�<Y� H6�ތiU"cu$�xB��M�<!&�F5S�.1S�Z)�ҦXO�<s�\�=0!K�ޙ*�T̻�d`�<QT�CS���gj2d�ˆ�Bw�<��BX�u���3�t� �� I�q�<)2�Y�itX�R3}��亓L i�<a�揣N(��A�+k��é�H�<��F	�l��D[���t���[��G�<'�S��P��W�Ϟ$����M[�<A�K�@7��Eh��SQ���!�RL�<Q�kM�)��m����<��@3+c�<�#c��eh@�P���/j��Z�<i���p��!�S����u�U�<I���jb6�81+r��A�%JT�<���~�(�h	�"����#�Lm�<b\�e���4想e׈�'%�g�<1�D�"w�!!��-\`�b�H�<As�S�A�Z�@e��B����&��F�<iT��j��-"�ڦw�4�S���I�<��i��g�F@Æ�&�l��k�~�<!�P�l�1�n�\#la�7�u�<���RF:�Y��à~2l���%�n�<�q�#{&��C!ܪr���`��H]�<����Z��)X@�E); ,<�uJ�B�<1g%��+�@��e@�G���!"*�j�<���/j�q �U�OhQ���d�<!��h��`��-X�V��8�`T�<	d��
I3�̑��[:I��L�WM�Q�<�3�D�7֔U�0�T5U�ZXcä�O�<7�?E�@C
�$�p�+WlD�<!`�4�.-�`-�	Pf�3)Qk�<�֦Or$ 9��^�Ǹ1�%De�<Ag']'S��J�Z�,@$���Y�<	Tf�I�����K� G�*a����L�<��K͡"�t�h�غZ���4BJ@�<	��'D�P�FQ4d_�d�mT�<�8X�r��hT2	��t�t�<��B�r�����J��L)l+���M�<� nI�q��.6�vDZ��E�0���s"O�q�����yAPp蓘cK\E��"O�T�#�R�J�0xY�m�_$����"O�9���6K.��{�*4z�xH�"O6X�"Q�U��|��+C�\�����"O�% b��E��1��@�B�n��"O �R��Wa½�$o:\���"O� ����5�z0�O"`�"O�u�� C��bv��y$ E+b"O4<y���rpہ@�6.VXI�"O�ũb�+i�&XBA�P#.�� ��"O�-���O�~t�EN��,5����"O�}���ׅ8����®DC�"OH��W�]�f8�`�& ���%��"O�ȨE@Q��<�w�ؖ��"O���6+Ӝm�A���O�.Ya"Or�8æ�"w�"e�sMɃD�60j"Ob)[���&�Ȕ2�jܮy"���"Oإ��l��:�M�P�!z8��e"OĠq�G:p�0���X���"OL$3��m �c��OF>�R�"O�u��(�:N��,Ө^"r@i�"O0�*u�O6P����J�[ �Mav"O�{�-[${At9J�G���Qc"O��)ɰQ;��8��T�w�ڄ�"OjE;�(ݧ���C�H�(�@Zb"OTlQ'G[t-'`,�`�Y!�W�?�2D��W/�� 

/j!�N���yd�O�:��<K%�8%G!��	��!(S�C�)=%Q���{h!�$S<Y���'��	 ��PgK�+Y!�ɝ� l�E���+&�R�'�!�UR�,X*�Z2PU"��#��c�F)Yu)C&er�{��S�8ay�������5C[KH�H���`才�ē�i��D�d���u�VݱƮ�T%�#�O���Q�K��k�8b�"~�R���S\J����|�NM�F��+��2����<��dc��ݻi6,���Z�ɋR�C>�el�$o����g.is�!q�>��49��<�?%?�S�Ù
]�Y�p�2r��B:}R�Z�d��O���i��X;$)�33�=�<�Y��O�%AE8�)ڧT=���y���KH"q�\qKų�������1��`W!YCň�!2��#?�Mщr�Gv>%��(�L��Bŏ�v`���Q#=�I�0Xn��?%?m١�
�+�o4K��$I!�9}Bd��h��O�D��˜"C�&Y�R�v3��H뼟,:�O�U�S�O�p�6 N�I��Jr$P����p�!Hk�⟢򖏐�i��X� �K��,��+�o��Or��ǧI�2	V�Z4�F��2��sL�|����H"�i�0�(�$5�7. =<rZ����ʥ��d���D��\�V��0|���[��rW��-j�(��XR?7(�;�?q�d����𩁖5�֐[�/w{D��4O!lQcNM��x�g����$[�f(�pA�'9m1R�ݪe�D���,\>] F�G�hX!���ؤ[���'�,Z�
��?%?Yi*�?m�ղ�F׃|��=Q��'}r!�.��O�}��Ѥq�A�6LV�r|Y7�O$���(v�S�$+V�D� ���P*:�&U	��bsj�Tu��br���OOa9�f :N�0A�6SpMy�'�F�'�9b���3�Ǘ~'�`H
�'ܜL���:"�*H�Ǉ�"��
�'O8ia�I�	,Ķ�At��L�Z��	�'�"�Ё�&#9b�[V�T�5T��0
�'[5�J#�,���,%�I�	�'� ˅�'���d��!`0
�'��T�g� d*�����4n��=`	��� &�
�㛡��m� �_2Uۆ��g"OA+-�*d0��L P,D[R"O�M��t�1�A'
C��Ea "O�ȃ��:'�lL8#aM��I+�"O��E�9	̥�3�/ d>���"OVa񵩃&
6�8*���E+�hS�"O 1�D\�cԚC�P�1'=�&"Of|b��C�8�'"� 3�"O�ȕ��:�Z��DG�z�iAs"O�C�_�D��lԦw�Js"O��rd�8~*���ۂ%����"O��J*���B!k�*3Δ�p"OP�Á�
efv���fʕ7��=��"O���d�8E�L����)Zv谧"O8�+�D��6Ϣ���M	3���J�"O �hgE�2cp��l�>�2L��"O��Ssl������z`��"O�g!]n2�c��ë=yh���"Odi�a�	�2�����,\��r"O�˲ ��^����4U����"O>��ҪR�/���$��EQ��b�"O��s�J�'؜�F�3�}��"O C��@����A�U�����"OH%+��N/"`B���G)���c�"O6t��.5��4�$�_�p�R�"O���]4���;��а(t���@"O4|�o�!�A�D�&h���"OP(p����+N@ia��_x�aX�"O^�R$�B"X�>}�&����:b!��Z
0�R�S� � w9t��S��`O!�D�b�<��ƅ-Y ļ�M�7M!�� &2��SIN��M�R�M!�[�uQ1�N�:�J�Zb)S=e!��`�$��q�@�B�P"Έ;E!�$�o
��Mۥ+"D �ԥu�!���)���V%�75%3rMA��!�$Z� ;b�Q4ŗ�p��8�˝:-�!�$�j���YVʍ�s�@IG*��!�dɳ;�����5���"�06�!�ݐm�0�V�6x�R!l�8h�!�D^�C�e�Dn���� �+�/Gw!�DƼyU�\����K� �V�_�!�d}K�-��ݎa��5��1,�!��W�cc�����xU�TO�A}!�$�~\De��6(��c���&�!�7A��*���7]:�"#���!�H�uN�H4o�W�\h�K˄�!��;p�r���cL�U
ep�a	.=�!��V=b��)ɒ"�?NA}ȓ�<!��[�+��1nR�=��!��b.!�C�J�2M@o�{6��qNY!�d�<:>f)I�B։c$NA"L�N!�d�;r�d]e��&@g	��C�!��
���!ugڳ ���R	��__!��1�x"�в?WlT�c.A2!��(o�du�󩑜KT� #���9/!�γGL�x��л7��F  &!�/�uA�"(�p��Lm!�$�����:mZ'�S4`�!�d�`˼�Q@?��9��B�!�K5O�
p�O�z�N�8CO�#o!򄜣fҸ��$��:�&u" a`T!�įj%B�JH�P��(� WkO!��vH3d�C9M�:XkQiL�?�!�� �m�e�׻O�֌�c��)J���"OL�X���OM�X��/-�X8�"Op���Y{��0�M(X��"O�J���V"�`s`�^!Θa�"OZ9z�Aٙt�$\r��Ķ8P��v"O�����N.f6�hr�s( ��B"OX	�N�0-�����D�%{^4"OX�KfdI�?.�ir%�\�Z�h�"O"�!��=�~�;�*�I2�U)�"O�����Ǆ%n8����D!l�C"O�s��،j�2�6�G�c'�P��"O��ZQ鑡�]�Ҟ? ��H�"O��J��]�t�)6�G5�@F"Ot͢� �j���@�f�ڔ�d"O��+�%>h�6q�ӎ�{��!��"O�D;!E�8Mͦ4r��0���E"O�p��!Т8��M�Ǭ�<3�)V"O�U�@�Ϫg�4�C�JA�Q�H��"OZt����|����T�K�y�"���"O���/��^)k񩐎;y��"O�}�X�b��܈���	n��$0""O|4�1hM&�l�P��"�d�"O�E30/غz�H�5�Bl�>�;�"OJ@8T�S����g��[�����"O�UXpHAx�F�"�͖!\���V"O��c���
;��B #����"O�9s����@��W�m�����"O"�J�Z i}����C�:����"O�ht��>6N����U5xmB�"O���S��J��L�����!�"O�`���(wA"R�ӖIh`�"O%�fW�>�9BJ�sQܙt"O�|{�b��p����Â14�\J�"O�<#`N����X�.�<�$��"OV	��'1��H[�mH�sw�<�r"Ox��Jߴx��C!g=Tl�h�"O�\S��E�
�&��~�R��"O�%-�#����&G�'��Ub�"OĀ��(�+K�<X��.1z֠��"OHQZ�
ނ | �Q��b��x�*Ojq���LD`C`FϽS�D��
�'v �U�ݐ3�K���Ԥ��T�<!��z,��"�]�@�����v�<1�&@�g�d�d����	U�r�<q����j�`�#6.V6M=��`0c�r�<A&/�3zIR��I_ޙ(�r�<�J	(]>���do��82�ZGd]V�<��5m��d�)��T%�j�F�R�<�# �T�Ն�fWnA���N�<Qǂ)F�h���
 2����_�<� T�6�d<B3`�Nn~���"�X�<i�T4p��y� �ZѸ$k�<I�A��xX�`{�Ȕc�<��mR�Q�$	�V!�| p`0�(�[�<���ލ,M�;A�0`s���6��S�<QłW5���E�)�v���-�Q�<��Lנ5B��w�K#G������L�<�`@�:?҈�E �"?����`W]�<c#��ML�|�d��m�"�խ�[�<A��Zaw�ARv�ϒu��$kEZ�<y% �YZ$����	x� 0�QR�<u�L��9�.,cVf�K�<��a��D�IX�oV~~�ApUF�<yw�C;���pi�:}�[ğA�<� R��-	�v����.�*؈3"O��@�kľI׶Lz��5�q9�"O,9��]�%j������b$a�"O:=	�m��XhBeJ�+��QS"O@T{�F8x7`$`��_6cǶ@h"O��'JP�]�7���1���8�"Ob�҈RmĶ��Y��u�"O��"!$
](CՆx��y�"O��A�Ez�|%ӇC
	y��p"Ol�KdN�2sPȓ¼H���k$�O,�=E��ek���Q��4z@6\�#�H$�y2�;	�|L���m|���#J��y��Ǣ&�l���P��: ����y4:.]�֣>������y��EL(xcF�[9�<y!���y�f�%g�ta���ؠ7��z$�ظ�y���2\�V�@��\�3�Hx�H�y��J	��	��!L�1����3*���y���J�pF���xA�s��yB�9�0L跋��\:f�{����y��14�#qW���##��y��E�P[�4)g�>'��-���y�8lZ�h�(MQ��@0�O�(�y�j����S�
E�h��d�yҋ�<��D �M�	f�ѠU����yJ�Rm�L(']4�.M�u���y2�Kk�����L�c5���yRMHG�`� ��^��-�o���y��V rśf+�
ҸSFȈ�y�	z�X�HBI�~�z�3�	ӽ�y�mJ�m�$�x/�&�v��7h��y"g��C�n�K #D�o���wIG��y�M̴$�kv�o�;�hV�s�����(��۵h�Y��}������؅ȓS����Q(ڱ$�|iCS��EuT �ȓa�BXb�R�H���Q�)�tX��"/TE���8?�p�cP D݊܄�G�:L���?�j��Ŋ��.L��4
�p� c��(�3+�\a��ȓ ׊@�s@��suLdC�N�Q�^���q�:�t�4O�P�R�M�[���������ݚ6�t��4j׼ �lt�ȓ�$���Ҫ5j9�K�0���� �b�G	�B�:��V+���6��f�Fh&��քɁ<H�4�ȓwTv�+"T�%�<�Ѥ��j����s�*�^��h��Ȅ�G��ĳq"OB�JQ���UA������"O,�rP���.3�ћ�[5q�r�(�"Oxq*D�^�|	�a��&��6���"Ob����,A�H�prˆ&I�
f"O��7̊�iᚥa�)��	P���"O~�ӳ�F.N:��iT<J��2D"O$\�&��@�dn�;12�}�D"O�<���~���a�M&+�Ē�"O�+b��%6�8��քr�j�J`"Oj5�����uf��Wj��0\ �"Otx�#�
#���ױI�D4b""OB��彰�n��sIz{��!!�GM3�z"/�f\2Л��3�!�䄻"JЉʰ쇫-��1կ<3�!�DNN�Q�p#܉b'.+1�!�dLxR @  �զɣU��A2$�1ĠJ+}33͚�[���<�U)��B:6�ad�M���'��b�R����=i!���p)}�($;&�ďr����B�
����N��f�Z��g�<k'�V˧:�`�2*]6�IQg�Ğro��Fz�dY"yAUN������"λ2Ep�q@�S����� 
�M������P�'��E�P�Y��t��D�I�k4MP2)Y����@
��H�����$��i��+X�eD��d�5P�xŇLvj7�L2�|��RG��茉R��/ެH�	��)h���j��*�6�.omJ��ʙ�Xk��2��0h�W}����5fA�,Y�(��NYZ?U��0
x���p���,:�Q��gF�a�\٩'�	�pi�2��Osx4j�J}],帰n��)?�U�$Ǉ#c�R��7����l]A��NL��@�/l�NQ�Ub�U8��#%W�]�1I��n�h�q�jZ$\x���+��P�0��mF�7��i�e'\�H�6�P���n�r�S�[�Yr���KP�:ɠ��
�Ob��`)]�V\�*aY��HOH`���%4xFU��_)+	b��g,�^Fh���ޣ ��c�$��9(���K��	r���<'C��� ��Q���ޣ!��3Bd��r ]:&�<�����#�A^�dlZ�J�n��wCѰ3�h�󀨊
9�p��L��z:!k3�9���� �N�H$ �J1�|��|��\5Nj3��:਷��[T�A���'e2���oԙ� 1�%�W�x�
�fR=l�^�)`�[~j���@ѩ6`8틆�����-z���Ӿk�\ɑS�OJ���ٖF�THC�'�>��F\�:u�d����
L�)���`d���e�oZ~���`I�$e�F�W�\��V�K� y�дeb���'oX�QTn�d@��oގ@τ��`��5k��Y*ĬB�q��ћ��25|D�F(�����Z���	[��]ҳ�yK~�q���@Qe,_�?<�I�gDF���閰}��'���!��\?�GD"�����'��a @���#U EQFތ�4._� ��)� +&�Z�U#1���tNO#x�E�6� $m
r��ޢK���7�i���d�gC�<)�oɲ˒`���'���0�$IF�8K�L��=���X�eF�(4/0 ǌD��/�&���h&���g���];lP^�sD�A�h�a�3�.��b�+M� g�K8#�6����Y�l,����	t꺀Sb��c�ɭ�h�.����UI�&62�8���E5`���@�a��kk���B�_�,�F}���a��^)hl��C"ZY�:�B��ڈ.�U(�H	�|�Eu��_���@"]�@���ۇ.&U�\P��H�>-�Y0�(	��e�<��B��=��I�5��7W�����a?	E͒-:~��� �aby"�ĜU�(ղ3'�)��v�Ѧ�LС��S�f��D�L�5
,k+�N,u+�kHn����`� LO��8�/�<ߪ�Q��(��5{�yA�P;9ռ-�q�B����ى�
��c�G���#���%���pY�kF:Q�Ѡ�}x�Tˁ`�?Zh����H�=4����ʄN\����I�-��K��@*=O�@��\,��S�2���C�KU�0�e�H�)��b�)'Z+0II%-��@�B�)�VC�b�(g0�tES�-Y��#f�hc�)6�����k��E�<q�	A74�P�ic-���ni dc�@+Ci��2��Ԙ1�x2̔�Hja��38C��U�y�%�~Ix�#�0�F)h�LՀx��`2�ʗ�9a���F�V���\]/�e�&���&� D��5��!�uY%k��!iᏒ	A�\Q�p֠��GG����S�.�)�R�X��[�ksn s�)�G�Ιra�U�uܴ��6����O�]+MM2OQ�9a�&w�dy�K���(�4e<lOx�У`�� �A���mb̢��4Z���pÙ%l%���6�i����P�3n4��m[��ॉ�+m�%j�A��M�P����-RlH�%b
�E$ � ?�3\�d�!eL�VdQ7�	&�cC�L�R��a�B"Q�$)������+A��Ĉ:16�}���YМq�P*T��+��Y|��!�jyr3�D�<�@�04�_�!���	`#�Y��ģd�r!Y�Α�i�,�I�"��g+H4zFT�9���#��T�& L�cu�H��NűM�4@�k	�B��N�D<�D�������j+`�6U���9@"4g�~-�3*�c�8I�S�L�G.��p�?�<�B��?a�6�5��j�'Ta��:��M�b������.ci�y#��(pMԌ#דy���vj�5RB=�#/K�C�9����w��PE�T?�����1C�	����h�.�Z"g^_	�{4�^/�`Mᆊ�91vո�(V?Ej��$��
Y�L�?�u��#[�8���Rs!p�b��^����ԉF�H�x���
C�B�����H�|��th��> "t N>I����i�>K�r��J� G���D�'��<��#�WX���0E?/j�4��O����aI�{U��9���a�j ��˸^����卜By�����oiD���I�
D�-��#ƫ2^�Պ&���L��\�*0|�JC�,jcV�Dz��D_��c�ȈI�"@CT�ũ*�Zx����7ݞ���	�5G�N��DZ�$�&I�B������L��D?$ ���8�H�y�H,�rA
���h�����1]�01+7O��1���V,�th�1��S�w�:S��>9c6e����'(QZTH�gD95�L��e����.љ�~pq�k�5[v��ؒ�,O�e.Z�x�ђ�
�5H8�sdfТo\��ˏ�&���.S2zf
=¶�]�]��
�� �Ў�1ze
5��Eݠ^��:NM
�&�7P�o�L!�Dڔ6������!Hx$(�O<��I�A��l �S+$�l۲F��:4�!�4�d	�	�0���	0�z�*!((z��t����z��L(��Ƭ�����/H��:����KD�i�@�������v�͞����6.E*Z,H��X�m��Y��I�k�P�ZY�D�S�G7y J�۹�R�n��&IT��bLX���(��T��T@;2d��.Ì�דdB8��*Ϋ"j�r���h��m�aD2�Mk��,^
�ɻs-\�L9Ȝh��T�UL������=��-���ek��"%G	,it��F\$+�&)�דqF�9w)�+J�4�w��&clH�Pb�ƌ7"B�0�S
O�q"�iH���!D(c�dJA�<I�Ȍ���JhT�bF��$���t���(V c�p��+\VI���>��+_^]�^}�H �/Fu���ގ��"��+"�=� )��La�}�W"��3�2l�b"���d�4&�{",��,B�.+�%�0	n݁�{�`M!�"���*.�`=�CjP@�L�Y ��%Uן�13��0��HBaő(UXe�&˹<)�I7f���klP��U�m�AW�G�.X��a�0=m4%i�4��䕷f;EӲd�QcM0hB^Ev5.�P��7m�Q3"��0��Y��S�خ5q�LP�M�P�fJ�	��5{����<�tMԥ:�;V�J���4�� m�0�����5~�����h!��@p��(��ɻ�N�@�	s��ˢI��y��BhQ4)���sЬ�C��ēN�*��BF؎}�a�J���d.�� r�yq��<�TfXUpb��B|�km�Eo�i`e���pЇ���U�6�tF8&��ɦ��8cH��o�6V(��B�j��,ڳf�0X����
f�Blӳ��Ar�� k_"m�(xVI�<ے�Qf�]ny��5!
�(��	g�1f��u���R�����'�`c�Ɉ�|�݊�D��~8��;��6��|��N�?E����عc�tu[q��&{���^;z3�����tZ�.4=��1�֋7+̤@��7,O]K����k[�}�D!V.L��!#��ˮ@Z<��A7��kq��)A;��:� �
e�Ё?4�r�K/�?����7
��S �(C8��Ą,I� �I���Ѭ�K �Ji�I�:�y�7`_W����u)Y�<Jq#��|�M	UȈ]Y��Ba���	*%���1g�J`�ԥ�1F��H�s��*FH*Ev�$IX�?q�K=� ������֟C�@��0��""�H@o3{Np�9T�U�����
��w$�F�^�9����qW�M�g��ql�z���w��a�eY�x�"5�	�Z��6L}3�,��cAIJ -�@Pi���7#�"81(�D�! ��P{>�,�C��N@2
2 Q�l�
��̃�z΅����2D !��b3O�Yh��C�`�m8��
L�f0�0�� >�01��߃/���h�-I(K��9�a� /���X��	�J�*9���K�U���r�`Ԉ��dj�;�Za�G�'<�}+2GR�[�v�9L����O&A��R#�@P)��8�$��kO�|R��Q�3�,xe"��?a��k�#�1+�@|���T4i�8�3��7:0=��8�Be�V�҃9k��[�#3�	"1�8�Ag�V=�UڐU�d8B-
�蓠wp%x���v��LƫAhmJ�㏭�l<��!��c�j�
��Q�{r�jfd&}]~} "�%|���W瀨bNv|◅WG���P
E4M��lc�a�)?�D��2%H�Jt�D�43Ь��iś-^ؓOʜ�	Ę+R�EфꅵO�z�o��"]~m�����,#є��ą���6��&��\k�C��\t���D�	�d�FA��'R����JOj� F�o�����[z��D�t�6AΟ-F����
O�X��n,c�8hG�ǐ܄�J���&�x�2n�e� ���֖�z�'�ɩ�-ڡ�u&�F8̚�	�`]8߮=�����f�x���	�����:�{�t��i��Wc���*���6w���oO)r2��aÞq�h3�g�j��"�C }b��E��L��
Z�L�@U�\cQ��x��L��0?!`�?�.1ˀ`�kJ��P�����Ő�LS3
���F�UĎ�z���:�4	ː �nE��լ�C�!��x���QCY P4(v%�S�h�BA�.R��� �%��Qa��#_��[0c\�AT�2�/�v�8�
	39�%+��E-&�}	GN�!Z��C �3@Z��I;~F`�vG�_�����;fX�"<q��K�r��(�m�1�<�A7sŠ�A��H�
2������I>���..a�p�)�f��`BE�����S�1�����䅈E�h�A7/+n�ӷE[� oZ�p��X#>D�⇺~S�MZRƄ
F�`�·-,~��g�%%eN� t�׿��d�r�X/ yXCF[#ut`��)��-:��$0K��O�~n��ҋ^0i]2 �@_�bU�w&	�-��5�v�C3M�!б��}o� �r��1jZ�� ̉�"ΣvE 	c��^y�u;��'��ؓ��#z�PuQ�c|�x�٨,�lT�d��6o���:��FQτ��2/G�O�i�V�)er�@u�)-�hX�4ٷl�B
U�J��� ��7'w�,����(O���%�U�N���;@
@7%r�8�S)[]�Vu�4��;9�A �a�
ԩ�,�+i=*��c��U0��! �?Ǵ��Vc�81ўt��#ؒT�]�����A��ك��V'?9�= e�`h �/Y�ijjy�c��M��#@����/Mwd,ۅ�X�� ��A��"��y��˘�X2��ь����>��f	6Mq�R���`����yIt�i��i��X"ra71�o�?�H�R�K�%����c�~g�--�N+kC�J��c *ix��s J٩g��j�O�+]:]yE��[��l��b�������C��U!]���ɵ�c��?"a�+$�b�8�:O�"�)�^�ށ���j��I��I�����e�x�W,,�����xuyz 	C�X �$�`
�og���'�&�8ȪU�
3R�,�f��,f[�ش)B?n¡hU��mR�#?ɢ`�I��Îĩ6ӌd��.�3,
x9Y4c����P�(��\�Ӵ�WD1B����p�0��1,��=�V@��Y<���`b���b�F������8{���6�^�Z*1�>����?t?�a��"E
����2"O��o
�|� 3��W'֨BJ6w�<4!��'�.�H�B�q����O䩛�K�_�Jl;u���X� Z"�'J��{G#V�
�(x�1.�tMTä�I�W-������%�x�Y��'�ea�-�r��	 ��̕�p�Ӊ��ŶR.ġʦ�ݡ0Q&4ҩ�@`1H�$:�EJelč.鈘�"OL��#$��5]�i;d��%O�2�
�V�pїmаY�2e���R8�?�y�LN+` {q�̮Y�zM��+D���ӄݥ��9�q�^�g|8�Rr�G>N�Y�'\�����<��Ϙ'�ԁ���H�"�Ό��H���
�'���qC�P8(��k�c��2������X�6�����|��|2�_�v����o�/f��d�'<O�� �/ݯ�ēN�QPÆ�/�*��#Z�(�\��G�:�a�aA�*���bIL�\�8�ȓX�Ne�����.0���p��4Y���ȓ~昅���]�|���kѬ�h8�<�ȓXj��V���+�b,a�b5a���ȓ9�a�aϛ�v� 9�BĒ)U�6�ȓAZ��U-�!lH���k��X����ȓ	;jp8��l�n\����
��I�ȓ^uґs�䂌V�L��$� b�̆�|:�CQ/6���q��=\Ȅȓ8:V�ق�\B�)s����v����Eƨ������ {��:�"Oa�lԎir�c4&��6�@�"Oj��`�Q(&�I'"X(�J�h�"O�@�V++C�L��4d�8|6苡"O�l���By*y�VE
P7�,r"OX�`��,��yQ'F6a{"O��R��k�XuQD�D&Q>9�"O�����?~&��%�
]��q��"O���s���.PҨ��Øo
�"7"O ������iA�ο:ۈ�a�"O��3�mY�P� ��i� ��ebd"O�����Fy�(� �X��99�"OR�+$R����A��%J���V"OÑiL������C#���B�"O����G�O�xy��C��
1�� �yҁ� ~7�E9u�ˢO�-y����y�b�5hR���k߶Q��t"l,�y���e�@�H@��U����ejVA�<qӠ
9 ������=	�XZ�ĐI�<٢ R+��0�n�81��+t��J�<��m�; ����sM�q��-]j�<� 園>X�%�G��"-;�%;��j�<�B�'Th�c� E'�U�E�`�<ї/䩑&��>Q&�s�N�a�<9צ��V��H���V�I{%B[�<���[(y�n��Jс~���c��Y�<A#�P��h8"J��T���F�[�<� H-1���B�C$+$F���R�"Ozt �L����ܡ㪌aq��Q�"O�-)��˼G׀Y��fE����{"O:=��KN��8��t�9zB"OȰ��ϊ%x�҄hsǄ�cnpLk�"O��A�	����s�W�2W�i�G�	�T��)�ᓚ0���3)��=����BB�I�!�D�{��N8 �x�PTCʮL��dT�6�������)�'Q=RA`��ǳ��=Q�)C)4+"
�'Gv-��t�Z��&�'/f�ժ�4%�v	;�^
Sܮdʤ��=Z��Su��O.ai҅�<n]
DxƉ�:�j��4�'q5�%H_�`����,A�����]!W%�õ���h�|�4�ߜ;h�bu0\O�h��Q�8_��a�g����,9��I"�tZ"�P�<X��y�']���8��I� [�D8CGK
�.��B%I�M�D�"O���EO� _f���&F��$Kq��H\��BR%�kdl0� .B0����O/!]d����3�j���ׄ���c��}⎗b�T9c#F�j�g҈Y֬MPA���(Z��"0v8���ݞŹA<��B�g��\ݴ�O�"���t�¥Qc�Ȥq��hB���/x�YO<٤h#_'8�ʣ��8�M;��.3�Q�E�{5��S&a_f(��������'���g�A1����U�v`��'|4�B�AR�N��Yg͊_��5k��+G ]�� \�vը�E�2t �:4�'H�4/OhuCg�@I����wWj�k�L���:�J�'��0=av�@�D�C��Oҡ���|��u��fY����dݺi^i��ߥ8b����_3DAȕ�Q��}��a҃�������wnԙ��~CX-U�� �t���$�#XH��(�b����-C$�Z-�8	�b���$X�(m�PFXi����C) ��t��S���*���=%2�B��$Z�$M��&Y��ē|(t,��Z�Em�ܪ���"dЄ�w"F�|&��y�4[PZԌZ0�D��oD�2��,�!�$Gβ=c0OČ!��`��C$�츶$)C妘yC�	�4M,�¡�nA��d.*�(d�xrC" M�\X��V�9�ji1�,���8"Č�w�r��co�`͊U�1
� %A�P`��<�naql��R�D)o�PQ2$�%Jxp��1HKV�`�����T7z�"��)�=���H�e̩I7H�ɀ�b8| �Bܰ$�:�Q�e]*74�q#F��]2!�(��\�18�i&c z/�=#���PTƹZ�Ǝ�p 刢U���-���	�K�˟,J�G��l�,����ۑ/���Hpȣ��4OGҐP�UgD�.K � 'T�%�Z� �̸&&J"d�E�p^5Prɕ�?ؤ[2"�!CT^ĉp�T!�L�X���z��]���̂$*�N�� ]3�x��%M��}�,D�r��
 �c�O�[�ꀓ��C�+���C�v������=��52ҤȪ v�b�
)�n��H#"N���q�(t�����)�d�BF�!'$zU�Ql��"N����h�b���,pr�E/k���@ȅ6"pyÑ́ #	���j6h�L
[�fPH��3tAf�ė�g���6� �"�R�ظ&8���k���S�D�Ҭj����� ��va�&S�fE�Ɍ�j��!,�i�t
%�6E�дR����4��	�Q�h��5Zb�`�C5,tp�+�)F�w�pS޴�x}�&�O-y� �H�n�o��O�0�0TNChƬ�ʱȕ]ը�pVL��$Q2�#���P��%͛c���%����ɯi�`sf�O0�ء7���鱅I	�}{����p�����E��zv�8��8s���Q n�X��p�G�1
�`�)��H�&84���	9aq���'6�O���'#�]}�@p�ܚR��C��ݤ>���ej�� �֙a�N 9"�Y�s�L�\�R�z`�\T��KJ~Ќg�n�`��2�2U2*�
�B8Gz�ٲp��Th��n�&��~�5@!!�h��v�@�QQN����С[	2%j�,�j: Z�%T� �' �d��������h�J�P�ՄN�"��j�?`�Ftm)�Լ�@�ۆF�J��G���/Ң��ɟ8�2��4Z�U�c�bB�`i������v���h�h�䊔 ����\�n����d)e)$� ���t���6�Hy �J�"��QN�${��Q,i����B�g,.�(��J�r���f��Nw6�z�B�b�|̛$��愑��L�ʰ��D��yC1��,`-�VZuGze��,� )�R�2h���PG$�T%v�2j��+n�V�Z�wBri�R>�i�K��Lq���A,_�tE�5�Ñ��Oz��Չγq%>ؙ�+گK��h�W
Z�&yf$^5'F����ցq�(]���ӓbL��D+_�h	 ��~��'T�x�&�L��(�&���c��B�i��l ��U�� h\�L36}1䤃�	�ӡs�$�$%Q�M,BQ�f�\9�"����fb���նm��5Г*�H�����I�?�I)�F�d�q(��H�j����wv�0 �؇#XE�dH��=�]���i�M`R��J�j��S��7�м`т�����A�c$ �����n&���V7�Q��٥ER��Hvˈ�ib%N7�YR�%X`���^wN�X��ea�QQbY-"0��i��^�*��0��L-q�dU�( �Q�P��@���"'M�'X
�Z@͟.j� "�@%H:8yLY2]� G���%fD����rɄ��@I�t�l����I>�s�1Oމ6+P6%�H�ä+�1\�@�#��O�%Y&$Yq���j�*�^1˕(Z�d!�u��GX/p��5�RU�]�*7B�,b�$�#6 �t<l4��� �v+$�b�Nýa�\Zӓ2�n�K�A؍dl�E��nO�=��c3�G8r��vfؔ(��`���6�z�+W�`h�M�ObX�p�kM4A�̋�$�_�8r�e�)b��}��(a��l+p�)fIp�-HYG6$���4`Ì�j�d�&#ߎd�E�B_|I�OKTB2M�_L" �u�6d˜�*�W B|���Zޖ����ʍ؈O�"�C	�3/"�᫚R� p���ѭ4HH1��ߴW�άl�������s��Q�q�PE������?		\`a'�^�])x�j�o�)� :�yf��zT�ɀ�J�
�5B$>O�q�7�n�zԫ��C�"��B�_���6
Ǽ��Rb,�Lq��F��thIH��M��,� p�+��E	K�����Z��ax�F�.�\��	� Xz爅Yf�X��i�w�H� ��w�X@�eN�+�tPGn�w���Y�ܙ"� t)�i�E�C!K;����(`���^�LU�eMr)t99��_;�<���+m�R��s��7���A��C�-]*�^�rR�<y�YBD�>P�ʑJ�n�,8��-[7��0^�Z�FE5J(�F|��9g�V�HfK�"G�ʀ�֩��Rzȡ3�ô�*��S��
	��q"��
�I;4T��Z�tPUL2c_�l��RF���C��V�(5�ō�<�OF1y��"�ë<��
3$�f?�SE�N�Q'�U$�$����8\Z�Q0��tZ�Q��S9x;�5�S n�R�P� f� !��<���6J��c�
92vSV0>��@*�eH8|�4����\�~TJq�!cE.T�DF����'j&g�d��Kk�|Q��Xަ����C��T�@�!Zr�d��;�~��1H.*4ⅇ�.A��zRDB��v�!�
�  ���81&L6s�2\�#'�s��P��}���NW�jw�p 3���D�A"�l�dI��GO�7�B5�`Jךf��u�����[F�F�'j����a�kU
�:/��7"��Ŧ�-%$�i{!F0jH�sn�!0� �2�b�A|8�ք!>�L5B��&#�uCd��i@%��Ε�6�4��G��4��G�3q��,"&R����8f納�,'d�0C�b���Sv.�G��U�Q ͟䪇$�)vF6=I2��.-�cÑ.F�"��!)|-���7:��7dѫ�HOtЉ��ɝ"7�;��b�0uU�-���A�C��8�����U�~��B������2A���:'�OQ�pE��v&�o�lht��ş_*sw :�p=�Ɓ-2sL��g�["oSn�갊Oh���
��E:z�)�'s�PӔך9)���M6+�pE0�'ȵ�u7f�9��<ۥd¯f��5��_����ɒ��#� ˂Waf��C'��9ȰzB�*d'pܛ�/�`x�b$K�%Ӱ�b&���X� kP�A2�Jr��*e$z��EOS2mn�"T��&�:LX7P�	���i$��R�L��x�\/|��j�dC��("���0��DJ�(1K2\�	�Q�`�+ąL%�dY��H�s�6(�ϗ9C_�LJ�ΔS�TY珃 U�l��%���'��<{6B��D�A!�*�������b)�PďЕ 4t�
q)���+���B�aRc*����`��a���&oѳ7��pR��"���#�Ћh�+�Hʦw�(���X*�1��a�1Kw�-0�ǂ�Z&l����æ%6	N���T @KA�,�XD oãa��dK�
N�� T��5n#���r��T0f�2/V�q��	��I���Ի��\�m��6b���-T�=i������7g��YXشD�@���Ե�n�ȶL��hC�Dx�Xu�q��j�N�XcB(D��π�O�"E��-Y��`�yR�J-[���Hu$5:�T��џn�*�E)$��yRퟹ|_���dަW�Bap�nU�$��ge�?BH�yJu�ԇt�F�*��8~\��ݒ��';�t�a*��==�2��-=�h��$�������e����x:���?9��'rh� &L0`�.���̍!J�:���ǧj�(k�I��8�����'iF��D�F6h�(u�2OV�Z�|ЗD�N�xT󦎒�.�r��5�@G?��c�6w�8u�L.~,��S��Y�z����u4�"��ןp�B��
��|���:��
�<��8�y����b��M��)Ҷ�L?A6��0J8mz&�5YTr �F���T�4[���D�Al���37�W�d�tQQ�d�/5�k��%d2%jU�A7K��	2h����ƒ�PT�Ԍ�2I��ON�)0�M*b��H�L�$��?�"c�% �TA����F�L>9�L[OQ��&���Y���� )Ʈ��](c��7�B�Z��5hE"�%���+,�52�(�����W'�ekꊴޖ�R�˜P�|@E��P��h`mدv�ƩN)LO�	 G�_ }�<�yFOQ���!�;���3 ���n� �whU�����Y����Va1{�H�h!,]�8����	.>W�%�� Cx<:QG]�"�r��ô�&� ��9#OP�����?<�	�'ƫP�f	�� �<T�x5�H��:vl�2�Kց~ 8��V09�
���S�n���R�W�t!�#�gpM��#
%yb-8�M�Z�,l%�B ��$'��i���j�|@�� ϤIz��/,��ڶ
�;7�r�B�`
E�2�1����J��L��DR�@�KÚ@3�0�1
չ4�z�R��dZ���8҇b�!��x�3 Xo$��:!I��~-����&=	��fB[(���'"�%��l�3��m/��B�	H:Z��јUɄ�fږe���$"���eh]�_�\�B�-9lO��i��EV:�[R�(z��X� ̓��Pde��"Y���G� �E� ��)��C[$�3����}��P@���U	����G�^���0�N4<O頴��.]����.ԑ[�J�#/8�Y"D+ b���H�#\�z�aR2,@���/�=�Ej�%""�	��D)%x��gС_�p|@�KJ�XV0!C�0c@ ��"�"�0bC��rM�&��l�5E�:P=[��A>(� \r�
0"� ������+�j�s�HPc�1�P��1��=A�<Ap�G��<6�8�N�}��I�vy0��#b��`��(�~舃dW�"��4:/Ά��q�!gO;L�fepB�Ϡd��H��ȝ�u���Ԍ�&�F���(�\x4T���S��Qbj�9�҅��'�U��J����T'Щ`� �i+����#,�EՂ]�0N��F�k�	�6	V���B	�h72���1�R�Ӧ3h i�O��9p���տ���Yĥ̽f�v}�D���>��鶧�6��B+J�$���(��oy��kA/B�xe����;���Ƨ�3��d�O����&
��F��KM 6p<s��0E���[&&5�J�XU+L�3z.$C�'\�Y�u�ƹa�M��)��Q"s�\�[�f����t���_$0T�y�I&ғ)uP� Δ�+h��H�O� X�͓r��!�^��"f�W�d�RP��?,@�pT(o��peo6}Bf�8��&�]��B��h�*|c(���	�0?��bQa��������!��,M:\!�y�a^�xq�R�jٱo�֠�u␟d���ׇ�����,�����æ7���/G�h;ge }�02�;.�ŨD!�KR!i7�'g��b�WVޞ�@�ĕ�v��xb�,��RJl�Q�MICF�.�%b��z5ė�Wې��I:G�U���3����"��H�#<�'��p���Ԁ�5a��̄$z�6c�Hb�? �-�&�ݒmvT�J4���Y�P�TA��i�����B�5�ԝN�!�V�<�3
�d��Ӌo���R�n��/r�+��O��"���M߬6��̨���;7�t��Sn���#��)y�c�N7\t�� ���!��iC�M�F|A����S<H(��I:\f�{�lȗg�<������t�CeG�E΂P!�ahuv�P�i��<Pr�3D	�e�,�V� ���ݍL$��^��|����T,,�n�����lA�ףǤ�Ƽ�Ì[��*�� �ʀ>���JT��?Į�{�iÉ�0�Sl��D̨��L�?�&��0�J ?���b$��O*����B6[g��vJ��:�{�	9�&���C4_`��6�ϟ �0�c1킫j첀�$�1��5x2*ē}A� �JH��=c�J��"�R����۾��T�;ړ�ʠ-,l!H$%��ѳ��ڏUg�3�"�G�*A�7�޽*Ȯ�@uF���MH&N�P���E7�؈���),���&�!G$f�3���(�����b�1��>1ڈLW��B�
�<��R�$�'$G���dem�PeQ�C;\D�,��	�����%��z$���ɐOI�	(Q��ZV�]>kh���!�ܢ?(�}2�\">+��
�셧.X�J�+�p%�8�'��/lNX��bE�G��t2��|nbP�b��g��$��Ը2�l��y%��7(떬@O�<J��xۇE!�Wc,t��N)�DK�<��x@w��2%��H!��%�X\
�C��ۤu
���D�A0:_x��%��E}��N�Q.2�
E-]�J?贒 ȁ���O^�Z�	�*l�a��T�C�|hV��z�&x��#�3�azgBJ�('b���'=ab��4�.8%H���q�$� ����C��h�,B��%EG�@��iK�'W>�� ϩ�����LE#$�\��/]��h�FD�'W�Q��
S����Be
iF�$ۅμ�a��	J�3�Ɂ7��eؖMR+7�D�Wa�:\�����ܝj�Cr T:?|����|�z�	4��� V��Cgk����Z�F�B�,_�L�ny�H�!(;џ���x�"���e^�0���E�t���N;�@�I'�Q*�fB�3O�hu����?d2���U���V6���d B&E^e���3�7ʄ�Ǐ[\Pܑ9�N�vJԅȓ.�]�����\��HQ���1�l1��lQ5��dU�~�̈����dÆx����HǤ�tZӮ*C,��D�<Xb�x@8;�YA����w/�8�	F Y��� �8�N�f<X��(G=[��Є�Id8P���xR���PE2I)r'5~`�cb%���y2iU��t�I���%N&�ʆ�޺�yr�M (��e��)h��a�`䀉�yb��Q1�cC܋�x�ӐV��y�,�/�} ���5r���	��yb�ƸSK�|
���$��li�'�7�y�ۓ+���d���	#��y2����2'��� �S!I�yr�4Q	�`q��{��k�F��y��Ĥ���3!j%�}� �d "D�4�Վ�16�p+s!W4bġ�1+4D�|�q	G>��ؘ��b���0�)D���	T�2]�\X�J��AK�(D���2�J"ϰ�h������+&)D��S���]ô�y��}Kf��a�*D��@ȝ4`n9���٤S�|	���+D�Dqvl�?�2�Xbj�O�~}��#2D�x�Rޡ!�BYȒ��"5`�j5�-D�8x'F��7d�*�hȨu�*]@Չ/D�C*E�����	�7:mF�ʃ`/D��I�҅�� ; #��:�2d�&D��#Q� �7S�y�Q ΐx0��2��.�	?��Jd/��|�%Y�
�b��AS��OJ�q�.K��0珞4D�$�X�OD"}�Di�^'<ȣ���`iHI�ri�H�ў�:�'��m͸���X��5��+�m�'�ўʧ>�ΐZ$ͮK��`A�:< ��,��<E����&N���+0@�|��A��E�=���h�e�V��= Dl9�
����6���>)��f�O�B�g�85�ARAo H ��}~�R���'&w>)B��XVth8��
y�t�'��I��'�`]ٙ��	(&ع���S"D��FFA;}[J6�<�H>E�ԠS�v�x
��[�vr��P�lS���$7Z���C��&��)§=��aXhT%��I��K+@����@�8,�o��<_���OzH7M�*~p��0�n ÌZeL����/��؉Ԓ|��� �%货��u�`�'�O�n��Ā��Nz�yRO>���OXBC�hѸ+�ހ�2���D��I�%p��D��AçsuL���K��_@�q���mn
$������7��&�b?Q#A�>^U8���B�M�� ��>��)�4}��`J>E���H ��(S�#{�pT�BS �M�)�3dH��<�(��Ux'�H�NC��']LZ��P��wS� �$�[a~8�'wSܑh�M։[��b��ɽa��� �]	6�f�l>Tm09�'l�>����R�8J� rlN8b���VaD$h�,��I� ��+�h��`D@�����,9��IG�A�f��zy�H#ƀ���v�ɷ;�,��SgZ����(�'_]�<�Γ/}��)Tn��s�z�l�G��}��Oգ1��	�b.��������Ge[
r㾸bS+��T�`�p�A�~U��('�˫6���C�S�O�L,i`fI�q-�X�Qh�
�ޅS7�g� ǂΕ�D������y*�2e�Ոm�!����=KD*�F"OL���ɛi)���k�8n 2p��"O",�S���A�Ցj��H��"O��C3�ϽE�&�Um]�2�.��"O����6��S�
W�LI:�)�"O�}	��K��nT�≛�TB�@��"OVlH�X*���T�(D��"O�9�FւX����(p.�y����nް����Q*X�@��Ы�y�	�Ch��(eL@�OqJX;Ba��y"(xs���I��R?��c�.L��y�)Ƭ6a8p�#��Bj��P��;�y¬�]�>����K5��0�@�9�y�#O�c,��R��I	�ț��	/�y"*E:! �y"�*��zH�Aʀ#�y"��)[�e���L)VR��H@?�ybm�v\�
%����ո��c#!�Ď�%�]��Ã�z& kPc@�!򤄓�2yc��;����Eh�!򄆖:v�Xcs	�.���a�`�<>!�d
]
z� d��/���V1!�$Y�G.ȍـN�".������~5!��H�8Ū�s��e�(Iy@�֥D'!�I2G	D��7H�f),��O�!�d[�a�;r��,��A��
}f!�$ė��L*�A�,]�Ѕ�)^�!��!T�@���.���! 埐 �!�d�	6��鉧C�:A�J��񦆺!�!�E3@�$�� O�CQ�l����&�!�U� ���*�n"2ꂁ���Y�R�!�$��_�|Ӡl��.�F,z7�.�!򤃲RN��Rf���!w�Z�6~!�$��34|	kV�Z�l��ѠbËK�!�I28Sd���N�u����Ů�?�!�$�:�jc�
�"���'kU�!��7w$(��%�4-�F�Ae�!�$�4E|�+�#�@��z�▪N�!�&9�PP��ke+�����ַMi!�D��O�i��N/:��83�>F_!�dی%)����*.�B��i?!�$��Q�,�a�ɊJ���C��&�!�N"jԖ��c/�qﺵ*DIG
�!�ڡjG�(cg*�4ؤ%K�(�!f�!�$F8S���p`�*`�dPJ��X ~�!��0��a��ȑI���	5��#n�!�$�5l��0$�
*�kG���vh!�ګ8t��h���0;��ےZ)3!�$�z���k	�zc����CI!�@�t�X�U�$N��S᠓8@�!�ăM-Č2�C#?H�+�J1L9!�K�.d�d�2�
�2PRq��I!�D�}������#V��Ru!�� ��K0�ǟ}?�{2f�lN��"O�)�W����-sR��"O��P�̐u�����-Z�H���"v"OD��תT
x� ��;�n}��"O\h�Qff��ԉ���<ۆ��3"O��Kcܑ5"(��E��ld�	3�"O�4��i�77L$@�ָqev��w"O^t�A�(L��P�L3]��� "OF��Ə?b�T�6hܳ�~q��"O��k��ٵkc��z���^�h���"O� 1�@E�<O���p̉q�q�"ON� �NϮw+J���I��1mY�E"O ����o�,�p���W�-g"O�ea��
� 	�=Sa� 5�RbE"O�	�K�w&�!#m� 6� D"O��@ �8�H���EٔY�JAb�"O�P�p��7|���n�� (�A"O�T`q��0,�Al��~س�"O�}�4�J�W�P��5�=��%A'"O���k:h��#�I���zp"O�����t幡�>[���b"O�pf�W��D=��A1_����C"OB�@�s&�3cǇe��d�d"O�P���V���C1��T!��"O`UF"W$_$�h�φ5�1z0"ORp�Eǵ#�ly&kP>|lbA"O:|`�e��
Ci��1�lXkC"O�D�/
�BtУ�'�8k����"O�q���0r�M��蕂GU��d"O ��g �Mz堷�UO���"O"�F�!7p�i���@p��"O2��PF��N�����z8�1��"Oہ&�[������	�[��v"O�9���f��I9�`�Δ��"O�q������`�2��$k ����"O`���F78Ŵ�3aE-;�b�"O�C*ǓO3 ���ɇ6�E��"O�%�U�Ӎ!D8E�U횿6Ș�0"O��4@�a�n����DךD��"O�Y���R�>��l N��q�a"O2�!5n��0 �m��R?�yB�؋jhzA��R5`�����Oé�yR�K�T�,���	�Jacb%���y�f�;g�H���K���y��*��yҊ�OM�w�Jr��|��O^	�yU/{���cH�A��4c�䀱�y���o�:S�ǈ)A���&e���ybG�k*h�UPL�f0SF�W��y����`1"�A�25��/���y�BF-U���2䎓1H~��e��y�b��������-��a@0�]��y�
E�v����%M�/y�A����y"K�1	Zd�c��Ղ �@��?�yB�݆4>� �Ōҏwd\Q���y�m�١Ћ�0||��s���ybo�[��2*κd������*�y�(� �۶�U�V���q&���y�� `{����E�F+��hAJ0�y� 2O^H�1"�F�NP�$ӗ�y��%�A�sl��B�rm�E�Ɩ�y�F�1�8�k�Ď�h�Z���y�ρZI���
ء/g���S���y�Њe����ԫH2)M���b���y��P�=��z�Kʑ'�2d�tj ��y
� ��(��#B`���q�����r�"O�I3#�=dSxIz�,��"����U"Od���X9.�&M
#��AK"Oʴi�@8z�4Z��}�j��"O��Q��,j�%CcO�2=�:�4"O`01����Qw���X�4�(G"OV���U�GQ(�H1�2nZ���#"O(�p�+�f�};%�������"OL�Q�a�	n �]�*�%=�&���"O0���FS6u�s�<'�8�"O�0���9^@��KV�K��"O]�D��SϤu27�Bl	T"O�3a���{�riJ�ct�"O�A@��õ<5��2O %�d"OD���m�v,x�TLM&8q�"O�H1�(Պ Z� (Jr��"Op�K�I��$��+���$D�3B"O*�`!F����U;b >/̐ "OTX8��uf����K�uB	Za"O��K�C�[A*�##�2|Δ��"O��ꃪ7�>�jp�O����"O�};�E�1 2�11�^�&�jղ�"O��J��U�*sd�I�g\�v�}a�"O�t���K����"$	j��u"O������%4��٤�Ϳ~�굙B"O���C�C =g"qt��/8�D)�S"O��S�hйH9�@:�f��i�l��S"O~���C�3(����D.n6z�"O"�b0��Q��pq���	�2"Oց@�L��B�A�Bߔ3���&"O|��]&w�[ck�DȚ���"O�#1iH�P��ZC�Q
�H�Y�"O\��ӤW�K��`+ǢW�y�̩�%"O��˥L�	oT�a�B>	�J���"O�5�` �2(U*.V2�
"O�5A"�A�vF�N>v8�"O��B�#O`��]ҁ$� 7Ba3u"O.mA��ߊu���+�JGh1��"Oܜ�3���rO�7bF>}μ��"OV�*c�T#7�hK�۸#��y��"O��R������-¥ve��A�"OlZum�:˂ݙ��4$ņ�;�"O>10B����ћD��9G���i�"O�m�P�W\�h�L3���S"OJ�µh��QidC^#9�.�x"O�ܚ0��q��i�S���s�"O�,#��M�V�HP�A�GI.�v"O���AY���P��
"��	�"O��S�OS�S��(����LҀ�e"O��+f�ԣ�>� �J�H^�ɠ�"O�`V�6���+qZn�#"O�!H����Ny�M��Z�Gw�<�'"O�����x!�T{T�ޗ@~޸j�"O$@�-�!-l�`	�Xltڂ"O@�`��@�]�A���\%FKdL�t"O�x�OKA��%B����B|��"O��Q��$R�z��̷YؐL��"O����ʏ/9%&���M%�P@�"O�D)�b�-+"�J�m]�����"O�i�uk;@�C2�K�Y!t<R$"OD|!��H�F�� p�[h�0I"O���S�R�!��D���EN~b��1"O ��1A��/���5��&@cS�"O�P����5��@g坌U��ڕ"O� �i�h�o��0�
K�-x�'"O(�X$�T�X1�ら�{݆ *�"O��xu)X;1HhT�,|�b=2�"O�m�"��Y	�O�<<���F"O>h�T+өbP��(!˓'�*[6"O!��,�U*Ì�@��Xh�"O�8�A�(���+�+&րi"O,U�aF��qҸ��cbtd�%"OX��DExV0���(*�y�"On������~��a�H�1�nhR�"O8QY��P�b��
L��8G"O:���ՙ1�&��VnĹjܐ�Iu"O`E�a���S�B�"F�װq܂q�b"O����F�7`� 18 ,�-�"O�����5��3R�C�A�N�8�"O6����<y�T�1g��,]�,��"O�9p�Iq�:�i�8M��
2"O��   ��   B     �  �  �+  �6  �@  �J  PU  `  �g  s  K~  ��  #�  ��  �  E�  ��  ʪ  �  O�  ��  ��  @�  ��  ��  
�  M�  ��  ��  5�  ��  G { �  v `& �, �2 �5  Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�� |d��"O
`�(�;���8���-0��1%"Oj4��ND^[��"3/9�0|H�"OB���H��*�ʞRy=a"O�味V�!X��!&F�:J�$���"O,��a
���C�Ą�M�"O,$3%o�-���p���+Ն�:1"O��ݢ1����`���y14]2��i�<�6��{_���c�H�`�fX�$Kn�<��A̼VI�xR[�)�Ć�pඤ�ȓA5��('nߡ4�� �)˩%� ���,��r�؊b#`T�eT09���ȓ!�b��g��}�8�F��-? �ȓ
K|m�ș�VṔ���2�%�ȓ"R�X�j�4JN�1�˘X�i����̹	_�jZ��1!g��zܶ��ȓgil,*�J�
j�Ne��i�J%b���f	�(U��:���G��$Y^م�~r�� S�%T"���k\�jx�ȓ|4�1�îJb��@ӵ�ݩn�V��/[`�"�v4�R�!ʎ<��M�ȓ`:��z�ؚh�J�Z��$HY:	��H��p�m�C1��!��B:��0��EnjZA V;9����J[
2���	��4'J�EA�IVW&��~�(aZ��ӹ�>� o�Y�|�ȓ�f�A�
Ο7�H��M�$�����mޠP����/���ANXo*�ȓTv�����{ ��-7�*h��I��sB�8�8���3����ȓNe*M�悡;������X�o��!�ȓ'lj�#F�m�+R&;�|��2)n�C��0S4���T:
b���:�0!��e֊��)��ͷV��,�ȓ0�&�8#���� ع�L�����;�P�AFd���,w�6d��r�EQ�( �gVlɦ�M,H��,DP���|�I	$G#\���ȓ"�)���E�B	yt&B�^�LɅ�4�� ��eëF�ڙ��n��R�p�ȓp`@}bŇ�=�$�AUN��P���Gx"���z��:DJ����,?
K�`�P.B�	�#����E�/�6\�&�S$|�8�	؟8q�� 01xk� 3O�:}�C�2D���F���rN��� �M
Љ�s�4�d��?�w�0�3�D-��\����;ZUؕ#�LXvIax��>9O���2��Vh.4 �AQ�*G�$#V�e�4�'����'�e���������S<^��%�	�'�ʼC���IP��I�M
[@��B	�'z�"6�R&#V<UI�a�4W���ʈy��)�����E@���#qaԻ�,B��B��E�-(r�@� �<�.%��'���y2�V}ҩ��D8b�H�4�Ԥ��y"Ƹv�>�c4�O�Z���S�7Wr$C�	�zz�� �cĘ%lRݫ�C�0r��D:�S��4O@�'�8R�� /�F�rB�a����A0Onb��D~����K�Bar2Ƙ ��ٗ����y�n�#��!2�"~d���&����~m9,OTO���D�jfԂQ�ٿI��,Z "O �Pd� �e&��G܍���%"O �J&�D�fMe�R�c�B��"Op�+h�,/�*���-��	�����q}��� b�9�@�>����숷q�Q[��Oz�	�.Z�؆/�/*O��q���/����+�����6<Ύ���P�|U�'~2���R�B\� �[<+�8+q�Z�	u!�$���.I��ȝ�m7�Z�A!�$�~�|�HD$ ._���ܹu(��)�'uC*q�4�Ԋ8�#��<'�i�'��H�꒡F���LR
1�b̂�'̎U��fS�`�D�B�DXW�A!��Ĩ>�yB:OLq�6cɒB���ȑ��T�0�a�'N�˓N^TX3�Np1�U��°<d�1���S�'�y�3a�O��p�4��Q�u�'�ּI&a���8�4OZ-x�f����x�
6P�5ȇ�M_<bF䇉��d5�S�OV�-�����hov�3���-^����'좀��l�3K�!�Ѝ�V��$h�y��OV"<y�'���%�;7"q� �V#n�!ՇV��y�i�6H	G�U��=�BT��0<���P�d��q�O��f}�e(� (�!�d�"9�*��'���&�8y'�N�Fy���K�!e[x�����2t�� �(Z#�y�$D.[�T�[EOL�|��!%ĥ�y��&
4���)J��p�Q���y"��M�H���Du�,����p>�I<�ԇ��Pn�����_4h�$�ic�G�<�gGRF.H���$ڰlcB}�vOCB�'�?�&�?��u�V&V�)h��#�R0�x�$��[6��Ф�aLD#U����y҅Q�0���H�B�S=t��C�^��y"��)z�\��+�u`������y/�Y�X���bϿr�Vt�E��y��8�$!�*�,a����V��y�&�<"���D�-`�t(�4aW��yr���^p������[UH�����/�y2�i5a~B�W'~��듆�"Y�l4B˔���=��y2�K�}8޹h��8#l|s�f��y"�+~�Li��lnM�4�p��.��'�
�$���'�6�O�N}�����2$y&��7�2x�
�'�i�P#ј�*3�,-}���d�>1���i��Kʙ�U�d�f���,1[a{��$��$9��@e�ą�|����䓹p>1�m�1g���HCZ��Ԙ���|�'�p�~z.�/gY~�z��SF ���B�y�<aE��)��ik�A
8f��H�wEt?!d:O��`��ϸ'����᫖��h���&+��!�
�'O\�C�	 2��i�b��l|�'zBm"1��6���p�D�(����'���4<J�T ��?�p���3$��c��66�бFS�M��X��`,D��
#��eCz���� r��E�B )D�����ĸ��I���&Hʌ)��+}r�|��Z�*m�ai�3r*�T�̋���B�IL0|`F�
�l\E(�A��a@����S3��A`'�
x"(�³�Z�X�rB�:�V��)�����ԢS��B�	1F���-��͈��?H8���d8?IO�$c���O�V`�C�*��`�+D���qK�,G"D4W� H�S�-}"�)�S�w"�"gͼ9$�8R��
hRB�%�"�qLN �BŅ�%�$B�ɱ@pN��,V8zd�ě`�:��<���T>�3� 4 0a2��0�\9�D�*D��`[!sÌ݉�/�rA�j��>���?	�' �f�� ����/��W�i�@�V��y
� �t� �ݱ�����&� j�8k�>�e�D��H�ʬ�$A	0�ܕ
��oP�ɵ"O�M0�l�'
"��B$�Si���j��iDP�	k���O�¤��ڼ@�,�pby�T(�ۓ�������M�R�F��+V��P��/�S؞D��h�8�@��G�)��d3�Ho�"r�0�G/_�9���'!��>Y2C�	/)�<����pR��B���m�(C��?��D���*G���r�%�HC䉁C�H�@�����1K𥞋�
�'ў�?2��#J`���va�a$�-,O��	E}�OD�1+ݝtd[��J�AЌ2s�'���v�'�v �u�5�#`Ѣ���'�~l�����A��<�l[®;�'�������2\q��Q�\���Co0�	�<ͧ�����\J���b���J�x�$���xrcJ�n	>\�BjY�Jh��Y�#X�C��?�� g���iY�](�H�(D�B�	�U0IY��.�Ua�I�mCt�Iڦ�װ=a� ��N���a��#,M.�X�T��L�&�EҦ	��ۄ'��@��� pږ��>q
�T<9Z���Y��AJ�#&�>�q�>و�	?��``p/΀�
�(ġG�0!��_h,@"Z&��d���X��hO�̉�c#�W�bU�'C�(�8T"O�� �i/K	\�s�(�6J�J���"O���䎁�=ZN{�_�F�Y�'�剢Z�`Y�d�M�tB��4O�C�C����P79(�m��'Y/�����N�����O`T ���>rxR6�\g�0��'bh�aC���	�`p�ŨD�e���'��Y�!���\ (�FĐˆ��'����nL	Dd±0R	$Q�>�s�'̰p�%[�/��9A�H`؎�@�'ҚABq���F.�U`gI_�*��T��'�0��CI�% ��<k�*e���'�v�p��	U�`�3`�� e8���'f��2a1*�r)9�J�8צ���'+D�ԅ�.F
��$�ho(�B�'o�h�VT����M!h�
�:	�' t���H��4}�]�e��2J�>���'�f� ��$[qذ�t`Z�:�^ě�'���e�ΝV��@4B�1h�
�'�~�s鞡��4*V��J�Y�'�4а�b&�ړkѹW�M�'�r	�`��e��A�v��VOj���'�8�iR!�O�l�Jvg�xf�0��'^P|K��� �<y�cE�vd�
�'bd��w��3|�]����n"x���'�< �$�7�Y���12�|I1�'{�a��C�~K��cp�Ҩ)&x�'��)SEN�^h�����tL{�'J��aX�v\���*/D_ 5��'=�����)f����➹h�ya�'����6�ZD��-f�(�'x��f'ۖrژ�$��x�u�'��Ɋd%��6:�,qɒC	�(S�'�$\�������q��eB�H�	�'�Dm9�E��=���6�Y%uH�'�|� #ͻ�>X�5�K�~u��'e�	�7B�8�^1��nR�J�x��'���/�]�&pjE�F�@�ҽY�'������08H���#�L	�'�|(�bl҇:Ɣ3V��MI�`�
��� �ՀE�*��i{c�z�T;�"O�0�F�b�ٔH1zul͚2"OnU�'�0�j��e��!k���"O�9�W��"^�8�F�]��"O|��J;g�
ȑՅ�L>b�00�'�]���	ɟ��柄�I����I.��ZW�e;�IJGj֌:���������I��x�����֟x��۟��	�e��K ύ/z�}R��	9I�T�	�x�I��	���ğ��ӟ��I&zԮ!���<���cc�1;����ӟt����h����x��՟��	����Ic�ApW�R������B�R��Iӟl�	����	̟l�Iӟ��I�|�ɓ_�����HH�)Ad
a��x�I�T�	ڟ�	���	ޟp����x��Y>�����)#m]���5��m�I������L�����Iҟ���֟X�	�z���G#��E�0ٻ$�H5_�J�I@���<��џ��ӟD�I��|�I C��mᣦ�![)�u�'����ԕ��՟������I�����ꟴ����|�	�\� 5���&�P�&-��P�� �IП������I���I����Iٟ`�ɍM���uj����-QҀ�-��q������	ڟ\�I��������؟���Bs������b�,�:�暧Sh�e�I��L�	ҟ����$�	��I蟸�	�jtTM2��4'tP)4��
^��`�I���˟���ǟ0��۟�#ܴ�?���e1̴�deG�%y���h�ZКS���IBy���O�lZ� 9���D��s�j�*42�� �,?Yu�i��O��O 6��D<�UA��9(�D1���pTo���DYg��¦�'���z$�]���`Y���D�����4{ԭRW���O�˓�h�
�)�`P��d�2�-u�q�˦�
 g?�	a��r���wK<Pز)!����C�J�� Y���O06q�\���-Ā�۴�y�d��)ظK@
p0t��i���y��̸XC���{�ў��ҟ�S$ ��=HE��(W�^�1��s��'��'��6-�j�1O�v�.S4�����۔�^w�9�2h�<���MK�'I�I�4X��͋�*E�"�,m��NH�M82���|j�"-�uw��O@$�aފ*�IiANT�'��t�%'�<	/O���s��Q�d�LV|�C�Lt k�<H޴W���'J�7�!�i>uh��0.� �򠖶}���:�㶟t��֦=��3N��n�V~Bm�v���!I?hs�paub7�l1�WAf%�� �i>��'�Ok<:����Oo��X'Ykd��O�n�8Glc����X�M��9K�E	�X`�a�!ղv�&9/O`��qӼ��x�S�?��	�]ލ0GJ��%�p`'�Q kL��a�"q���J�4Y�j6f���ē����wO�-*�ÇvN�ʣ�c8��<1-O:�O6�o�'>]��	��J!�(�9C��8�'�g�`�	��M3����|��?y޴�?��i�Y�l˓���hmꁋ�h��A�&e�ش�yr��<pR��,S�f�.����JZw0}�1? P"� v��3	���T̓�?	(Od�S�O*
|�M�Rt�3�BK�z����y2aa�J-������4�?!-Od���B&Zޤ�%��$L�d��Cc�l�'Q��{�D��ԭR �7u���֥�,�ة����/x2}�d*)r��Ô�ïhiV��"�g�IG~�O��LJ�咸;|0�v�Q��l��,b��'��hٴQ�L�<(�D`�k^�{~����E�Ijqњ���,O��${���Ig��?��'䖠]{ة���Ctl1���
~�`��b^0�����Ub���u�&#��ҌQ��!�"�:_ �c��հ�d�O���O*��)�<I%�ij�J��#YUF�J� ��0���� ����d�����?9�X���ٴbe��E%�=F��y�ug�)&(l(3�i��6�ۍh�6M??1t%� ��-�5'���Ě�b���z%��F�H2k�(W1OD�D�<q��i��M��9���;�i�ҧ�]�<|l�?pc����Գ�yW�,�J�� ��+��"�.t�^��tӎ��@yJ~ZpG[��M�'<b�b�%0~V(�,E�V�2���'��9����Z�k��|�R��ݟ��(�6+�� ����W 8��ޟH�	����Py��`��đ65O����O�x����p�z�(���� ��膍,���O�˓R(��a����I}BGܹ55�Mz�,���j�n�y��'���ҐaϰS>�@�Q� ���,��1�;4u�i�yp4�rd��B�ߎk��}�r�'6��'J��'��>a�Ɍ3�V�����HDNR�5���I��M������CǦY�?ͻ
?����y��p��LI�%I��̓*�6|Ӵ=o�+m4�oz~r�+G��a�?1�l�ፙ<2Y�e��@Ż7�|ɨ��|�P�����l�IП0����G%1�P�9W`�(� %B�*_y��v��(�h�O����OΒ��Ė���@v O�U�,D��;M�4!�'87�J㦑p���H�xX�F�#� Qa玈� ����qN��S�� ��G�<I�264��Z[wz"�O��o��0J �e�v�pv�,s�|���?a��?	��|:/OzlZ�e2�I4Ǵq�����`c��HC4�	�M���Ľ>���i(N7YΦ��VnJ33�������"s����0;L,?QE�H<V�H&f:��'0�k� �1{S̄�y��1�1��	gR���;ON��O����OX�d�Od�?!i��L"Q�2U &��8N,f)���`� �IƟ|k�4>j�'9t7�;�������S��)H�ܑ�Iô�ʔ��x}b.h�t�oz>	(��Cæ	�'Q�e�"*󠱫�G���(Ui���
p���*�ўl��Cyr�'s�<�F@�c�|���G���'�'��6mJ�1O�I�t��b]�1�t%��
�=��u��X�/O8�����I|��?�æ��&VaD��u�L*�:��Ԡ�4l�"�[�2]������_�u�$�d	�l]�(�'��I�g	����?(O1�����MK$�[J��N�a���i�\RΑ�'�47��Or�O��O�6�78�:5jƫT�*d:��\5X
uo��8� �V�MΓ�?Qt�)3�^�ЉNF~R���Z�c�(h�� � �Ø�'�2V�0D�/�!ؠ���"+\�`��HKM� 74z1O��);�)Ȧ�8F n�(�֨ᄈa��ϥ3:k��M��'n��"�)�O�8 ��e���	 ��jqϒ�8%�j$C��oL��ɯ'"D#J@�b����'z��腌u
$���E�~6�
�'��V�	,�M�!��]̓J٤��ES{nHie�0	9�9����C�	ן�m�<	�O�,�P�#$l�bĘ�/��<O��d�6@A�4S I�	A�	�?�XƬJӺ"�'[�1�C��,�6���+�"��� �'��'���'�>a�I�=� "Vh�?K���$��x���I��M�bɑ���$P����?ͻ\z|�G&�pa�:k^y�~z�ƀhӜ@m�
	|�|��c!?E˱ 6�-��'W���!Ł��iK�M9���J�TaJ>1.O����O.���O����O�Q��-n� �2��!��s"�<i!�iXЄ8�O��#��'�Tq$�AV[���N��"��ؠ�O�inZ4�Ma�'6�>�(���
e]�-�G�D�Tz�)��)���`��<!��9?�a3  ��ã�|�]��� �� }��d�����x�
�*��̟8���� �����RyRt�d�S��O�m��R ��<�k=��m�";Of=mZ^��O5�ɔ�M��iƴ7M�>(�9�g��i������!X�����f���}�����LO�h
2�H~��Ɯ�qP��h&�ipÂ�%*�࠻�6O
���<�+O?U� 'N���Yf��|�V#0�3�MK$�Ma~�%bӞ�O]Rf���(6D:�'�5���Sfr�D�'B���� W(ě��t��!N�z�:c�,��F��, ׏\%�8�w�04���&�0���T�'w"�'Ϯ����UC��ٱ��A�P�Jr�' �Y���ߴo��Y��?!������i�~9����<
�2 )��P�#�I�����Ȧ�ڴ^�����P�.��C�EY�Єk��A�+@�+��T�'/�ũ1B�<�'9S
��^w#ҒO��c�K�%�M�����,B��O ���O����O1�X�w���Y� v�rq���zR��s�)(�Ua�W���4��'R�4����ʿ+/���F�ς(�:y�m��c�Z�o�yA:�m�~`�3	��СШ-:�ɃV�<���R�`LR�2�M�
~���	{y��'c��'���'��V>���Y�t(�֊Ē:��I�s�ρ�M�3��<A��?�I~���?�;U�zĀ�(Yh�N| Fc+BS��i�z7-�ៈէ���O����E�8-��4O�a0�D�2����<�F:O>< �#t��Y���-�d�<q���?�#^�1	>K��L�u[@5�eH�%�?!��?aB�<��$֦qY䃐�?��	��ץf%�}xU%�NL��
���X�'�2m�>�f�i_�7���'a�ar� Ҿ�ǯ��M�"�	�'H����gbTչ��¸5��?���C�ֺ[�'/�n��k�(x�V��&�Ǐ.H��'��'��sޭ¤��;J�פ�0����ď��P{�4f�,�'��7M:�i����k���&����h%�z���4f�f��p�P�rӚ�5�\KֈԠ<S��|q��#��t�U���������Of�D�OB�D�O��DAs 13%N�!:��{3��J�ʓsכ�3���O��?Mˇʔ5>�Y���_�8�؂�Bɿ��������ܦ���	�� as
W�p�f�	Q�L7W�:-�p 7K+�˓$�4}h���u�"7���<s.�'�@�eĽI�D<�@��7�?a���?���?ͧ��\���.{��r�(ɨ&���:�n
X��9�o��|{ڴ���|z�T�`2�4��}�,�Cg�7U��s�#.㞌�u �!e�7�{���I�qRl��m�\���'�dI~�1��@;�<��ơhݾ]�D�i�p��Myb]�"~�A�� Hf8cbƇ�;����AMJ̓%՛ƀZ.��Ǧ)%����Ÿ=$�dC,c^�ӷE��<�)O�7m���y���:�<nZ�<���z\�0@A\�B�5�G��Z�;�#��)��9a�^��hO��<���x�\i�k�N�كa�@�fИM���x�����'���O�޴���i�t�M�y<1�Oz��'��i��%�I����JS㟧�r|�5��q�:��ج\2�m�K�D	�I�?5�P����K�|"�&ƈzF�P7-�@�%k^�s��I�8������QŦa�'J20ŻÝ6,�L��N����{"�V�'�ɧ��'���)�X�P��]�qE�	�THF#��7M�Oΐ�7�q�$�	��iC�^*v�l�3?� �(w�?r�놮!w���I7��O�ʓ�h���φ3=�V��`��? Uʘk!�I��p�7��\��$���w�I[�Օ �Z�G&�&�Q�M�OR7-u����r���?�����M�'i �"�m�9�ڨ�1#_ R�����'¦���j�27�� u�|�Z���ȟ�ą��^�yV��~V邓���� �Iϟ(�IyRhӊ=k�O����O�������ș:V�&-��1�)�	6���Ӧ�j�4w�r_�\��Or*����8ٶ��e�??&ff�� Q�+D��䧍E��㺫c�'���"Զ4�b�X#�0��=
sY���'���9O�V��FE*�Pť�X�xk 5O��lZ���y=�V�4��L�*��6��ƃ�0����E�O
�$t���*W2d7m$?Q3�]'M�hE@s�Q*ah)[A�0� ��� �z���4����������udBr$H�{؎�'H6��1Or�?�����+&qf��Q,�9f�pb��[�����O�7Mr��G��o�.Q��b��Ev�EKEj� 䭓c %����4_G�(��Ef�c��kw2O�s�FǁWfuR	�\U\��@"O.���kC:1�� #�[	�&@�����i]HP�疄qi��1�A�3�0���[gF����]���v�E�"�\��W�L�x�q���gt�"K�H�"�Q2�i�d����J�ެX!ԮA+���kq�A�5n�i��5!V 9JMD� 4��'��E���߸C������"��w�^/	���d%j�и�B��lp�8��:�ٻE�l}2�'\�|"�']"&D|�ɛI�Hq��iU�-�|5Qbe�g�B7�O,�d�O����OB���XH��n�ԟ���(R��iz���798��Mխ����ܴ�?yN>��?�ׄ��?	��?���@J�9d�G$N�B����.n���'���'
RG^��b?���; ���M//�:Y����w�bH<����?�Pm��?Q���?L?�r7`Ʀ21�aiaD�8`�*̩�@s��D�O�x7��ŦѬ�`�D�jU�'d�����ד]��p���Ƽ~%�Aߴ�?q����P���?)���O�f��(Y�QQ.���$�*%#�H@�W�}�٫��@?G_��
#�2��{vM\1Dy~p�5'�$9���!���h�1�aB�P��DD�(�MqҪ9D�`�r": [f�F#���F�23��@� �o�@�Q#cN1T���� .;H���A?&�t��D�8�-���R��,C��Y�&��@�)jnb\����5.1�����S5�MJ'��F������E�V��uBڣE2İw�\Ѭ�X�Ƌ�>�S�fR<I��@j�E�ʟp��⟄�	��u�'��>���Qɍ�N9V� ��Xea3��$x��p�e�F�,H�f9<OR̉�,�Y��:�
��<'DI4H�
m���aC�W��L���(<O��Agęl�$���iK�].31Bժlp�h"�O�a��� 6O �q�r?���"Ov��,�$�Y��!��y� ��v��M̦&��ǉ�����`�4�ō	�@��-�>>9��3�n�蟜��'1S:��	����� ���ӣG&Xu:HA��MK@ \�
Vxp��gP.5~����ǎN8���vߔX���C�m�8��(�É�2x/F�+��غ mP��D�'FK��'�<�Bs��0
�O��)dI����-��?�O�"���u'���</%��f1�E��'�!�D ��r��:_^U��Zw㢜���M�.O���&������8�O��m���'sP�P@�И�R%-9�>�v���?���e�L���+�\,P␤�=��,QU\?]�O��&��b�A�!�L���N��@O{��"��҉DJ 8�2�UW�'Q���&��p�mR�U�M�����OL%��?��� #]�"-��hfa�2�3D���D� ���5G�z)B����.O�Gzrl-D��S�'��2 .\��7��6�O��d�O����f��b�D�O����O�F%{�4���B�3`�d�2�P��̳�ߢx�����'����*&�3�D\qq������'8F��uoI*X�u4@G�	����ɋl�^$����|���Ӱ54"	 ��=�Ah��!�>�O�-������Y7!1bx�ɑn~��FWn%1�@�s5ơ��-�1�@��'�#=ͧ��S��� �H;Dcs�W�'Xj=pA	Y��q���?���?q0��4���O��Ӝ f)P�aα)���MZ8|1p|q)WC?8�����e�䵊d�
P��)D{�$�z#��2�ȕ�1��kƫM�p�d��Gć�t�5X0�v�hI� H#ў��aȪ>�6�"T�Txr��T�����m؟H��W�P
�+Ǩ	6w0�j��>D���נ��O��E�4&FI���֮?扭�M�M>��h�Tl���'��F��yaL��'X���`�&s��'$hq[B�'"6�����4~	h���K̤l�*���6���� �O�|`�x�kư��x""��e�M�kV�U���'T<m�FԚr֖(��۹Z�l��Ri�5��ݟ�'3��e`RvA;�HܤOΔK�'�'��O>��o�5 �ek�/$�z��0�8�i޴ ;���P�:��)wdD�!")����4g�Z�lz>���U���'L
� b����;gA~ł��،`�hЃ���O��䕸y�T}iUL�$h��a�Qd�!P&^˧����%na�a2B��?��� @M�]��2��xD��"Y�G��"�"|�uA�!�0���@O�+O:X�᫙}�dA�VV��'!�>��	�}٠t��Y;�^u���=m& =��Ehn�煃b�k @
\n$��	��HO4���@O�����bjЉaRLzӅ�Ȧ��	Ɵ����X����GAܟ8������i޵�#k�J]�A���36@qt�m�$�N�|1�	�Uh�., 9geķ+h��p��i��(EԴn,������ʥzT�ؑqș�D����0].s��>�٣M��L�K�][uΖ�0�P<u��q�Q%� ;uH�Oq��'n~��DC&��lB�j�3l���'d$p� ��R�𠄉L#i���!�O*�Fz�O��'��$��7p5��hA�2eG�Y ��SC�'���'f��c�}���ͧ6����q[�c���Rs%�V���e�a<���ֶ��I	��]�Q�
�k���O�X�J���PO
�k�.\O\<��	ˤ\�Z�[��L11�� ��ҫ
��%�O�+�'�= ���3E�T >�{V"Ol�3`<eq$��E�PPdÍ��1O.�m�[�ɗDt~%�۴�?i��J��
wlF7�@��ą}*|�����?dKū�?�����K,s��<*�	 �BX�Y���T�H_��&M��\T�&��� �a8�#�S��!Gy�O�,�ԪE�^�����$��8Xa�2)ճi(�$A�:7����EX����Fy�OX��?5�x
Z��� J?�691�ƾ�y"R(Fw��R`��0݆E	��x��m��p�*�$!��J�.��`C�>�D�dm����	h�$�E:0��RE�!�"`5E�lLX�#͍<�R�'h�2���r�`KG�T>�OmhXq���+����$��R�dh�J� X��E,g��Q�ע J���t��`�1��!ɖ��U|6��5MY��z�0��>Ek�󟔣I>�jWf��c�h30@G-+*��6$PK�<w�60����+�&C�fu��oXk�|J��G�F�~�crbP�>�^�������DplZ͟���៰P!�4���I�<�	ϟ来J����[b\�{���32d���
��fI�M�Dvv�"� �e�g�	0 �nm�tF
��A����2CN��}����L8:{��!�<�3�$��I(xұ�̅I��IF-�E���%��iF��Oq��'L��!�
1�����X6�v=(�'�8�"���<	q+Q�[d2)p�OFz�O��'�zy�aۻZ�P��}�3ч�\����'���'�@{�A����̧gp����dߝgЄ�� ��0e>�!�Ê�>mP %ʄ6�M*�`]��Ot fa��z�猄� i;T*��'r6�Ӏ�2KΦ�	0��y���?�$��3m�	����:��b�ܬL$!����?	g$�;sE����eأS�*�3 �`�<Q� �� 7��0�I�4���CD�BH�Kk���|b*L�v��6m�O>�D Bj-qB��*7�9�pt	&���O2��6��O��d~>1���O�O� #��لDL��5<�vQ���'T��P�8\���H Q#	��H"�挎�p<�2"����YK<�鉥t��T�B	ЕQ�	r�)�V�<!T��zY�����#V8����f�!�d�ʦ�@�f����H��^z��D(IH�I0�y���|R���H�MZ����Ø�jq�Kd�f9����z�`���O�<8�
[4�X��ԫ�%-��P#2̩|b(�V))�@�-4Ȟ� ��|�tq�>��W1>��i:�$�35��l)�7�'0�v�맥[_��JF��z�O�ț��'ǔ7�Qh�Ox�D�ɍJ4u�u��O�J�	��\k���$ޤ4J��B��W`P���B��'Z#=��֖h ��`�O˼yD����̶Q����'��'��\+�_�/���'�"�'��]�y��q��,:%6
��H�AוJ�l��`S�
K�6�+)�h�L>1��6$p��Ԏ�U��	YA惨4��t�PD	{��7�(O����L>�!hK����7���*�(���@F3��'� �Ȟ�����<5���B�#�1y��Ht�ȓD"��ȅGK�)�����&�F4�'��"=�'��	�N�����;.ְ)�n�[����h�h����?!���?iý���O�ӢrDx"c��x����R,Z#�=3��M���?�"�Kj��hB�O�
=�8K�ȗ�1^~���'Ӹ9��P�DNH��a�Q����̣֯�?���'��xS�m�,J�f�N�ZA��'�VTZ� -wH��b@,��<�,䲎y��d��O��S���ɦ��I�D&�
C�hiÄoۮi��7&M�����vr������Χ`��	`�W�%�=�P�� >�Q�f��;���r�Ś`}�@�v�'�0;�ƹ/fm�1/�8�1���-:M�U�C�V�S���)�����D��B�j�ORX�W�'�8O�%(���^��1�u  9grġ�"O��qA�",6L�tJοGKj���ON�m�
Z�,(�F��6Y Y0��G[�(�$��z�IΝ�Mϧ�?!.�j ���O E˖E�B&��F�7Bk�۟�?����t(6�2���w
�>�O��pj��T�Ʀ)��5Z�G^3���' �=��	�Da��ʥ���J10�b���d����NѪV�>���̊ݴX	�>��Ӳ��O ��4!��;$;4�@����`��|1��E�`�xH�P,8On�Dzb��Tu��6D�N��QMӿ�86��O���OP�X�AOA~�d�Oh��O�u��)OLA@�� �p��.
�ؑ�y����<�w��G_BЗƗ�8퀼�~�U/��I�JD����)QQX�!R"�1ت��L>"��>�O�Q�tEA0$P�+�'{� ""OpŅ�m�\��B�4tlܼ����Dӈ�4���O:A�e��t%�p��\�Ȁ5�5���O�d�O��d�ͺ���?��O
�����(���¸P<��$�W�C�D?s��42��^/v'��!��f�'���֎_�e+��`���OX����n��d��- Մ�:԰ ���G+�����QY�'��a�NF^�`�H� 2�d:u�Z/�?a��'u�n��Qݘ��c�O�H9��'yxT�ÏH=1e~�e)A{�b9��y��~�̓Of�b��������П���P�/����f��V�"=0�o�ßT�I�T\H��I����'�6��	M��I���Q�PF�v<�@��h����
t}�OP��`�H
뢸��Ŕ)�x����' ����tK�'� Ӆ�B�$g�)I3+]*oڴ<��'�л��ٜhD�#��fT �'$�7-+	j謙w�ML+�A[V���_k��O��+"g�����ӟ��Ot�x��'�BQ�B��:J�H �sJ� *S��J��'D�m̹�"�T>�8�@b�L�0�	� �?-FͧO8ݡP�)�T���4�^$J�up�J�%R���'�6<��=�ɧ�O�Эsv�؈�.�iD�|�a�'H ��WAD�LZHK�	D�b�2
�uݑ��� ɑ�u���
$8y p�Ћ�Mk���?��}3�<k�LQ�?���?Q�ӼS�	�)^B��V�ێ]����Vj�1B���Cf�XX�h�h�m܏e̬%Z��䫑�_�r��	���3�ϖ!l��Ƞ5o �'�h���[/	����E͇a���r(�m�'Zl��pg${���&g?I�v\qg��'F��{Tn���E�� �)�3�d��H��\C�MF#rƛ�=�!�䁄9F�Axwm�&�1�m��	��HO�;�DB*MM���b��;RЕB� ����'N�i�x���O�d�O�����?�����d�c�2�X�N�SB ��
�$��)�'��\1��G�lG��zO<A��;����x�kG�m�F}�.B�C�֨H@�B�����k�ar��{��i��iِ-У�-�y���'�.�H4D�����c�mM4��'6�;�؁j_<l���0�I�Z�z��6��X"�p�U/_��(��(���ҟ����|��D
�b�j��s��0f�46�G�b�b��栏�e�H��*J�� eZ�Xa&�<�����e����S02-�q��	�pQԲ�D���A$�ݙ
�̨#��M���<�p�I�@&���SDY2Be��bh�8�n��7`!�dQ-���mۈgH�Y0#��F>!����SQ(�0��h���O|=T��q�ɒ{rHE
�4�?�����i�_!��$ە�b��$�}�	����2
��$�O��g�O:c��g~��S6 �����|!��I������R��0Y ]��RH8��Z�85�e��JⓄHm� ��K�����ׁǋ!N�'2%��IBɧ�O�f �: ���E��?�N��'�j�je��TЃE�35�j]ÓD����pPm*A���@p��	[)��@���MS��?��_>\�0���9�?���?q�Ӽ���7˂�[��
D~��a�i�#j)��Y�n�$HqIĄ�5���Ԓx��A0'ˊ�	���..�{��̚C�����$����&Z ,)��L>A""�G��0	��Bi�(x���2�ia47��O~1S2��Oq��Iڟ�2�MX�#x[!& �
�����fh<�b�MyEE`���'=�����ao~2m:�,}����DƱd�$��ˊ�]�VW
�-i� d������?���?��2���O0�Dl>Q���?�ju%΍��Ԡ���̧O��l�PM۞A�6���h@��<��'7� �l�sE͉Qy6@`��Q�N��˓mǆw
��M�������"���,J�S-�IE,�ȟP�	�,�Lb�aL�3�р"*	R̆�B	��d/�M���8�i�,�I�<�e�iX�'��0c�lӤ�$�OR]�F�$y �b��.hM1���O���5?����O>���PC�A7x�c娙,^!��Ѷ�͢k\�b��)[7�0��	�Z6��%�I�k^��� �0Kq|�ӇK�oo�T�%��e+���J>#, dȴ�l��L)U�	�PE���~�ɗL�����ɀYW�)"Ɗݘ��B�I�5Ms3̀0k�z����$)�B��8�M�SdA�s��l��.S̵y���F6􈀾it��'��ӬN2���I�8�5�fM�,��l�f�W�)t�l�I럌z��/l�8ͨA�b� %�_-^W�5���U�lҸʧ���*T�&F��衉I v���O���E�����C��ӅMנXj��_�&I�x˟|�R ?��I�bY�VuH��>��n���H>�J3���"�qh���;��Uq�G�Y�<��h��1�Й���U�m�������}�pڈ�ĝ�A����/j�N0��7&���mZҟ��Iݟ��@"�	!�����̟�݉9�0<��dA5=����k�vmL%�0��^#����O�> i7��I�g�	hR�C�`�h�BL7v3 0�`K26_������b�E,�3��A/-P�5�4��3X�P�v*�"c�&�L�v��Oq��'�tm�cD�\Q��Y� �H�@�����٫� R�bMs����4G� �'[V"=ͧ��uȌ�r��={�`�z��A�s�6|밥Q)z�����?����?�����$�Ol���$����29ۆy����HRz ����]w�����ƊA�.��wbI<��%���#S|�9pGKO?��Pd 3L	�JۄP�>DJ��B6e�����߉i�\�q��f�<�3r�:���dD�'lXȱJ�Ol�oZ����?9����'�D���c���Dţ�*�٫�'�, �S�V)1��Ș��5Rc$8�yBb����<i�bWl���'����s^�}r�![:!���@Ӧ��e���'�Z�1��'g;�8�2��>ap&tӾ�l�(���8s�W� c�����L�u�.���i�(H�������R �x!L
>w�$��QAKW#zi2E��B��4l��'&�u:����;�h�)��B�(�` q�j%�V�<�0咛
�2&�Y#L�3fɃ^<QǺi�
�3'��
�!�SM߷fH�e s�|rĝ=nV�7��O����|��j�?!�� e~.��bB���G-_�?Q��Fm�d�҈��A�8���;U*���'& �� Í�k�^�ID��I�L��O��ЎԵ��;0��8u�8�4�] ���S!�4#>��ݍ@N�,��l�)_ڨ<���ņ/��'��QY�c^ɧ�O�"4;U�O���(�c^,%)��"�'�I��(F�4��+"̈́�� �
Ó9Α��p6��,A8�-�R�Ńt ��2AB��M����?���F����+�?	���?��Ӽ�R�X%V	z�bc��x��i�	�.Uѳ�扴�yE�4� Q���L>����;j�i���<q��qP ���i���+^"ij��\v���MU���9 j
`�w�����%��1q���`hP!�'�9�D�`l��L>!�eI�O��5)�� .i�>���$��<����*6��-: OS'(0d�z'k�B~��!��|�J>�C�0i�p�2'��$R*�)*S ӿpp�Tɠ�'%�'�|�,�O^�l>}��蜎;������գ^�Q�h�-_^鸒� ����6`�lx���QI��(�A��Y� p����@��[A�Q`#�A]QPu�!�Q�Z~Fu���6��@&��`�e0eʕ,0���@�(=�R�b��'�X��I�HjA��ၢJ��A��{�!���i���Ӧ�ZIS@1�M�5BU1O�n�H�	�0�sݴ�?a�2H�
��!m����3.zF�����?1Sι�?������:�8�����X�B1Cm��C�۱�v�8��[.C@v����X����F����-�[̬�R�N�C+�P�gf�,a��if��v��Z�*����O��&���l�u� yR @G�,� �'D��Uo)�6�Kb�]�G,9`�H0�h�ڴ<ʈ	dg�+[�m�e `��K>�4��o�&�'��X>��G�ܟ0q�@�mhZ�	�D�v6:h�E�џ���C!��mZ=Wr�X�&���*�6�'F�`T���LQ*Y"`��i���O,���iS@��F�3H��3���}���ha�:c�m�;��l���+?�XAr4#C�`s~t�O&����'1O�0�T�R �9�ԇF\xQr�"Oʵ�U���#�t�Q'��
vaD��7�' �#=q����:���*�	9-����dH[�&�':�'��,`�g�uy��':���y�c����kHB�[{��ka6n$PpB�a�+d��� D�ϕ^�r��1O�5�c�H�}�z ��zd 0ђ�T+/H<yTIX(4;:����M=�h�+P�~�p(�zl�=� ��C@(:C�F(F�Рl�6�� �O�'��Y��S��h�	���30�� �$��-�*d�2�g_���<�p��C����#���X,���a~R(t��<n�L�i>���CyB#�	)�,�h$h[�(-�$u��E�X���aL�D���'���'�.��L�I�|Z�K�z���c�+W1,�0 ���еQ�k�^�
��L�V�g��؅�,my�}���4�K���C�lP�o�)��iΣR�>��'�b}���!(�qO��В��2D����0R'tȨ��Rd�C-r.-�O��7(Z<O�l)n��f�{S"O��1T�؉J�����f̰~�j���Ϧ�$��H&˃��M����?i� �O�b�sR��~i���U��?y�y1,I���?�O��-�Ø�1
�钂�X�>i�� �
�<)�&F[�3&�����p<�Vb��=��3J��J�C��>
ژP�D�i�� �L<�]p�E��%=��0e�(��YO>	%�ٟQO<!rP�=�T(ʰK�=$��MS,�<�&"| ��PD
�)�Hu�r�E}<ѽi\�1�恬j���)3CǦ}"H�Օ|�-c 6=����|
�&ۯ�?�f�<;8@�P�[v�Թp�.]��?����z��ɐ��=�E�F�W�6-�~z*�4��d���F��AjѶ9+�a�d�k�n}���a��pz��Tئ�~�����g�� �&�K'S��4��Q^��ؗN���{�j1D���OQN��#Y�T�#� ƦItx���O�p�n��7$,YӐ�т t�$*d�'$�"=�4��i��D��Y1z��B�ʄ@훖�'�R�'� #2�'���'���'��ם*=����@?L<���M��k@-R�l�Tf���ߴg]����՘O8f�9tM��<�^�]%�`�"kR�^�"����U��0�C���,����4�iP����e�Nɬ�'z����lv�E�	�(�lЦ�D�S��
��S���P���)�3�d�l�܊�e�M$j �䋅)J�!�^#�X��N֝j�Aq�6f�I�HO��1�d	�-� D e,��T<���տXP�j2I�p�D�O��$�O@���?���LĿ$�(��fFk㒠���\��h!-�:	&����E�Z�(��CF�\�B�Fi-�,aP�kٳ"�캳)��7)��pqK\XX���u:(� ����0�Q��[�CJ���]p؟��CMO�:W
aq��Ԇ<M��(��%D�p[F"�:�����Л��+V�8�	$��'�&�)�hx�����O|Yx	��pz>����y��rL�O`�d�ju|�$�O�S.G�Q��!��Z��S�jަy��v��e��H��y�:OT1��'�:���/®^�-i��*�6�	��xI�d�Ɓ`A�-�q�y��0��{�N���?�қx�� �H�jF������Mǣ�yJ<q����	c�9ˡ���x�b�8a�C��Z]���0�h�Ʀ3��4J5�lo����M�T�4��U�+���Ί�������"D��'�
�B̔7Y4�O�˧�򉒢U,A@��`$�\�^+l�����q'�b�֝�'�D9�R�0��Y> l���!Y�	o� ��1��I��	��D�޴�?i��t�	�<��89$��#D�`����
Θ'���'>�_�|��I����R�"Ɯ;S�
*�m���0<W�i�7m1�D�>�u��\�EʽcSDH,X�حm���h�I�pS�a��t��	ٟ�	���Z���i%���R�x��/<1��5���f^�����ZP�Ḩ��Q�Py�c��h�'i�D�Z�j�	��	$$�2�'�B��u�}ܧjĘ��6Ls��!��^.|T�*Ǐ��u�\�(f�K���v�\��)�3��;U}��o˖X4�-�D��6c,!��T�4t��@ H�:%�pq��A�d�I��HO�)7���\?�`{Q'�M�	��|T�D[ă�Rq>��O����O�d���?���?��ɟ�i�.,h�eL6\> ��.��T��:E�?zB�z�#�f��ybO�:^H8;C"̌�>�`Ʈ1j�E�aEH�?,�XC�ޗU숍���*1��[���VܓC܅�G+қ F,�I"P��{�����@ "�<�M[�����e�Fl�?i��ܷ<pL9�[���ȅ�w+!��	���[1!@� ��d�U� �$�<y���1P��Q����A9�u��'��D����S��k Oݎ � $���'�Ҥ�����':�	�e)
�bi��������3��ybA��@�#�okxEƈ
b�%���bM8�%�:X�љU���&��P��8 x������kr����-C;�rm����׷$��1�$3Q�)�`l�>��q�Z�}y!���g_��bF��l��eJ6��)m!��̦%��ƈ�0k(��g%âN!���b�r��6[����4�?�����
>8����X�$e:�� �K0>p��/� ;(�D�O,���e'X�6ѡ����q��S��]>�R�t��� Lؤ힙�rl1}R���{+�2�9c�$�h�Ξ�u`NŚ��/I9j��'`?P0A,=���!ׯs��Ot\Y��'B�O�� I��#�v[8X�ӷS\����"Op(VăBO̔ ����j^(e��'�#=��!|�-*�b� ��4�wnP�fz���'|��'��=��恦	H��'`��y�a���Ȱ* ��Cjt�b�A�-}�<k�@�4� �D�,Թ��|�m[�;Z6�t.�kш,ɓ���^��R��1z�(�#UJ�3�BA#�U(�˧$*���+h�m���i$�Y�sN�	[�,B�$�9��X�<�)�3��Sa�$]�����'M1�!�$�39[��X���E�:��g5��I
�HO�3�dؘ9�܌��K5d�v]�3�ˡl��]劙�>U��D�O����O�����?�����ᙰ͢�#�F�R9p��g!�k�J���'�|��oJ5��\�#��3&�����˄,�xZ�� !fT�,��T@0C��<��B���͟�
���|1��b��E��K�&����D��֩� Z���%�;T����<�B��ۈ�n��d�I�af����I0W� �˗�Y;�����˟��փP����	�|��DƟ�'�D�%#Y0Q�xp����"�v:�B&O�I�����r�K��Cx، �(�"/C�x"�	��?�#�xb��8��sC�@�9�\T$`�/�y����^�<\X7k[(B����aӣ�xbDc���Vi_�%!�$��h�%�X�G���dmZ؟��B�	`	\�Z�u�E�/e[�A�����'�~� L�uw��y�J��!��|�(��y@mö\�P7�ŧ[� �q�>���ŒO�Ƒ1!�!yn�Y�u͗�]��taw֟PB��ӥ+U��#��ďd��-���� ���'�fY{��xɧ�O�-�R#	'>J 0q��6Ye@l��'��l��Ɩ�=�q���2%�V���II���)w�Ǳ)T,pz�!ޔn������j���IzT�pU�U�u1p)DǒGאB�I�_�(�N�,!;PT�R�!��C�	�)�x{g	��U�&d���æG�.B䉵6"�QÅo�
�Z�Ґ�]�7��C�IUQ�T#5A�RyK� =otB�	=
����E�c(�%XP*֨a�JB�0e{��+�� Ip�h(�'��q��B�+�����k
,?�2s/��d�B�B��p ��$�D�'�חg�B�/�T�q��}x���l�$�C�əi��X3��
@�a�3��)qXB�IE tp�ʙ�^�xeKV
LHB�I6Vz�4�U�Y
ܘ�Y�X�Pp�C�ɴ=輢T�=� �s��P�-Y�B�I:M�.�@��<@ �ʕ(O0zF�B�I�U媄@ѠPP��%M,5�|B�I��r�c��P)18��M�P\tB�ɶ&�q����j�l��;�>B�	01����Qy0 �����#�B�	*�L�ʠH¾Fm��ӠD�P]�B�I�k��ŠQ��14��1yc��?��B�9Ɓ�w��6,N8y� 	�%7 �B�-]�a`G�k���[�I��:�B�	�_� �0a�	�$��۠+� E2�B��.4�v�@+5R�����
5��B�I�+�n���O6b$��`G2>��C�I�#~���`F71�A��m�v=�C䉬�ҳ����-�,� �ć�d<lq�-�����	�mD�(�ȓ>^(��.$�t9���? n8��Jb������R���Ww��F�9D����bQ����@A]����8D���O2t�b�̑��t��I"D���R�Tx��ѐP r6�A��,D��.�.o^0�+tj�W5S�>O�x����}�
]�D	 ;sĄI�dH�N��ɋ��4 ��dP!Ψ��'YU�7�@�ae:�i#'/P�A�O<�C�4`U�����(5���١�~rG����K�?�����Z��O(M B��3��T��Y�s��1���$���8'�\�o��9���9�p<� ��:rF_�z[j-!�+ӧ\����DfN�c��d����2R?a|Ro�<T]�5�GB�3
���jdKˤbuȅ���PX��%��0�:��o�x@�u�6�&|O&Њ�N�(�jY��-��Hj q��۽Y5�iA��(>d4�<�GN��� p� �˝��hC��HyҠ�_F>���īd�-�����O,�0���^d"gdA��jT�i�� �3��d��4�uN5q�  3
 �IV�S�@[��D3�0<1�M��"b�%H�"s��YGD@_yB�ɶ`U����n1A��iQ!����(O��{HE+͒ɚ�Y6
V\����OР�s !� i�Th� Θ VҴ���k����N^�v��d-=�9^��r��;���X"~|n�]������V�����E�S�O%Π����4L�4�s���	Bn�X׭�#~���{���)\h��BQ?Sܩ��+?i��eN�T۷c�9[],}Ⲣfy�mތ��'��8�eάAnlt���۪Z��A�:T�Hs���_��#��Z ��AQ�WI�Q�ac"�Lq���+*=P牡)ba�B-�5�F��qA\�N?�$&lTqOLӌ�9O��e�ބ���$��&KZ�T���Q��O�J1á<����h��B�=i�L}���D� !Xɟ����E}��'ZL�C�w)�<��Cۂ?l�G/Hv�i��i>5J���B�:y�c�RZ�4I�o]�F�Ex��ψz�t��φ�l4�k�Ϛ��$�h����i�4q���pw	iў����cdpD�4E��s�ܜ��eR�(P��P	aވBi
�H)u�1eX���d��zՈ����ቡ}Uk��#Z.5#$(E)�����Ӻn'm����� FBi0��z��r���-d��AfLD
�$Q�'���@R�'�1O��J1�ҹ?Yn�CfkB��X�RoJ�T�,�������O&��I��hu�n��l���a����\1�� 5�;=D�O���,f��c��������?if�)`���#�)r<ejFBp�'M�I
�
ܦ��)&�Wd,y��O��Z��DY������b5�`�O�ɔ'E:���OT�nZ�-�(�²iq2�$��&T�c��:��-����Z3����dR�)�f���ɢ^�<ȩ1+Z��0<Yօ��L^IH���Fc�аc�B��M[�Iit��`\6Z�lPnZ7B�N1{��DB&}�XP"�-Z�N�buY���7R$e�S�'T��>��"&X���c�U� P�,"#J�}�B`��&ˏz�Z�>	��r���v�������������>1K�?��'C���@�!|\ĉ��B T�
�1I1^�l An#M��l��ǥ (��gk�,v�9�'�������Fw��K���VW@���'�铖?��њ�jp����`	iq�~*���1��^�`�Xr���䄬qp�,�H���eg
��DF�:G�*�@��)��
X)���A+F������MC#�"P��<j� F�v��խ;?Q�$��D�Z"��[�d�!_
���O�`oL��d�����'���ɗn\>>j���� �0��-De��|i���N�N�'��`ɢ���3��,1ЙiS�̝�8��[��'}���q����n��f�Oh�p`��[D<8�h�	]o���6�I�5Q�`���H7�!zt��6S:��Z��I`./o:M{AH��n�8��?Q���?�$�L,^t-��:e]2pzS��I�,� �-^I�F�ڰ���`�L�0#�R,Y�$��eT�M�Xr�D(�0<��%�>Ic͑�cD-��H�d�ԟ���<9�Fu�v��$�fI��-�>	��<����-=!2a 6 ��gMn��g�I-9��݄�_�/Z�j�C(�����D�:�a����f�8��� 9�\�$Щ�	������� n��r�mл�	�C
�a���'o>�uޕ���*�p���l����X�&�O�� '�+hՒ�XC�ɚ��5������=9�x�Kσ�@��ya�k�)��O��ȋ�#O
8�LlZ�W��N_�{�fI��y
hX���D+�5	c��q�0@��H��5]�}C��J��0<��-�(9@h ���-���QF*�៌��6�I�/�Q>��¥ٷj&D�s���"/�.Ġ ̀#y�B�	E�6��ǡI�7���"�F�0��pR g�->���yW�Ɉn�l��"z�Qӆg�c��<�"��9}��!��;�O�Pтo��D�*%�1��A��d����	Ĩ"<9�5	�TH�kڝK�t�D��{~2�]����A��Ú/���'���O^u�w�&O�Ѹ6J�(���b�蕌d�h���(��]��<��d�$k���J��X��q��3�FM���;O$�h�@p�=��E��Q㤀).O`�+��J7F����I��E)�I�Us�1�����!)��[1�S�$/}���R���E
�HҠA��1I�G�D(��L�p$��I/�>q�1��˰jaG��P��'YS��O�<F��O�a�]����7�8��I�剽tX�c�M&VV���3�>x��ʓ9<�mK%��${���&%՘Q�B=E~�gK
)0T$��_i)ƍ���<�M[#A�;�@�X���,,��q��u�d�� �U	.-���A�[�豆�I	|�@��N�e�8y۲Dʞ]&��z�����e�2i�v��SH?�lGy"m�y����ë�,�8]�G�&lRɒ��� 4��q�A�xa���gK%�r�P@E��[7U��_���O��R#�(E���6!��0b� C���פ�)����7v������D�T�jP�F�߸ �8�Y��	'u�V�CSM�D)�Ԣ����1���	r�t�E��,%�L���gׇO% Dҭ�O3�A1qΆ��>��0h��b�8�ⶪ͊Yk&4�k`��2 ��.+ڭ��nR#!a�Ѻ�C�ax�5`�*�xa�U�3��b���:���-����c��&+j��AH�
�Q���РX�2�@)��):�~��C?N��B����NE8E��6% ��qaFP�[��K��D�hlQ�	<W����o޽�sJT?%s�t�F�J�z3��	�/��vA��{E>��a뒕~��/0�}���:G� 5�Q�O�96�Gx2O҆<�`}�F�5X@h�� ����
-9�J�P�Lыd0r�b�LZE�ѐG�,5K�J+�M?Q�g�	�&R�)��3�Xq�'��vx��FNފK�Z9G�57��k��-d䬺Ч�p���f�lj���Q�&4!:�S�a�O^�Êy�i�++���I-+�tB��ܢ���1eU�NEҶJ<�OD]9�wL T1�����C��>9��شj� ��ē��O`��/�#����C��	˅-�2u�(��*F>{��F}�猐X�(aT�>!p�'�Ӊ@�䕻�˖%7I�x���$�2/r.�!��S^�)s+���I6p͎|Ӥ�z���g��qD y�OT]-m�(��N�����HC��Y�49� �┻��L5,����A�6���&^���U���'��la�{���t~RЄq��]�2�J9���S����3���T� &���H(ʓZ ��K_�u$�c'-��h;
T���\ܓ]��"=�����C r������C����Q�	D�S�r0�E}r �Y�1�a-w�	� 4y�
Y�c�45c8���H��K@ �	�<��'��aQ�
w�I��߅��O�x)�!y���3/(�P�n0S
��+ǿhqRA��Q�^Q�'�a���H�"�q��\�f ��k,O�����I�'��k(O�4 �(O�0a�`�)^�<����Ү������I�L��AÃ-M].�x��9��F|2͜92'$ �T	o��hB��{��}sF
�<�ڎF~��z��4�W���(�� j%\���NW�6"Hq$�m�'^�T�>��w�X�@@Q�l�zq�η"\�޴C�	
&�-��ON���JԡKQ䰬�5�|�ؕkV��FH��9�|�OV����!�,q����U;��!�i=��e�OPx`v��$$�I���XL`�&�)\�����	����� O����4��&�Yxat��!b�:8�EDC1� ��M�7W�#����?�O�!���?�@���+j*H�0(��yM�$Y���)$x꽠���K�(��,Y�E{�#>9� G-	�h  �$Nj�9�tgA]�������A�P�D�<�G\����������kb=���,� )T�	�ð@��dE��;����\!SNt5����"C��wDO8.0�0�L'�o:I"6�@�C����z����c�S_���Q`�b~2��>�>x ��Ȩ�h��RdA�*q�ux�%]�K"�H��C0��#<	�ꁕb<��F[���E��,	g~���!Q'0���I-}b�խɉ?��OD +��S�3?�$��{;>(��G�b{:4:����"&�)N����%�_n�bjR���ei�M��`���Fv!Q��%�7���7n|:��w-�<�yR#�F�^#f�ө�*:W"�A�)�ubj��䚌8 � B��
I�q�r�D�u�Ȋ�I(# TS#K.N��I<�T�C�ј�ɰ7lǄn�����X�y$�K�).�;CvM���߼���/0c����D*1��!�+�V~(�t"���An_2�h��}Rr� >�l�r�D��f=��g��ux#<�r�@���H��K�H� �x2c�\~�OF�` B���I#,`{��'N�䔥O�X����o��T�"_��y&a�5� ���RA����B�P�>�Iw�� Ơ����n� �1�Ӹ4�hYf�+�������P�Q�����#��x���1�����KL89֣��W*X'!��P��剚|on�h'�;>����3��0�����o�'�Z�iƊ/G3tO� b`fZ�Aj���A�P������F�$���q؞��Y��eClR�%��.��t �*�DJ��U�O��������@_Ҁb�MF0}H��s�����f�;�z�KÓ+�xb0L�v�����M�~���K"�PK��,�q]�h8�i��M̓Hx$i���d���`�ؒ\��t��O"}�.UA"��˝�s�*򤉞�����)g�T2�AC;��¡"X_1O�ã�G����ddU&#���ҡ[!s���x7N� �Vd0f��a��0��pmДÄ��L�P�/i�fQ�� �&�L	�%��+��-��	�'�DZ P��!�s��5I
���E�<���ē+U�ų0o�(�V�@U�O�����j��p�#jC�?�x0KW��$�"|���N��MQ�k��	�+�,W�,a�ȓ B�Kf��t*#&gj���ȓ5OH�W�{��R��}�U��k��8��J%�iAfŠh�:���.	a��Ѣ1^ja�ɖU�ru��S�? x���ҽc7���→W�ܥ��"O:D33�&Z$<m���H	f"O>�s�O��+���(J�K���(�"O��h���iN�9W��� ��t��"O$�٢�?HA'F��Г�"OP��$�:%�zԧ�nQ��kw"O�(yW\�Rs���c��!5�h�c"O�e�C�u ~	KԥB.(ʁ��"Ox0��A5z�ip�F��L n]�'"O��(G���y�"��$e[�E���y�"O�(bfٙ@���eIF"O�NHXT"O�� W�̅|u"�Gޞ3�Pa�"O�iE�;I֝k� U6?�|��"O�h����;�
��D�r�~�U"O�Y�ѩQ)vp{�H�lL-a�"O^ ��h;dxԪ��H�XW�h#'"OJ`��E��ZYR(��H,���"O�-�J�'G�A�'-L�U��"O:��
�&��j�CZ�'>f��V"O�!�w�GgTd!��<#�=Z�"O���2 �:��p�W
�k��R�"O�a#��׍b�<1�� ���""OxE0�&CTij c'm�/jaH���"Or8��KE�"Z�s$m�;���hd"O�y���1n|t��Y2vw,Q�3"O�=�#�6.,�1gG�lb(i�"O8��$�Y�e���1H�A�I�A"O$\[�NȎ2�$���;2��a�"O&�2P�9����)���"OfeH�(+e0Ȅ��y���%"O��pTFu%�y���_�4qʱ"O�)�6g]NpY(�I($?fPc"O.���Zh �Z�+Z'4�a�"O�8��/�t�P�2[:Poe��"O��@�'�X�"M8 ���bm�"O���0%�.6��9M��`��"OrE�MI
E��a@�"<���v"OF-� ��}���ycK[��J\�e"O��S&ř�#���H ��N��D�A"O�xb��;1�H�2�߮�Z<KG"O�p逭J�L͸rÁ�M.ȵ��"O.E�w&�2@���(�F�7���"O�I#Wl
�3�ha�ʝVf��
�"O6�F�@�_Lj@�&Y���"OpА����Q�$a�s��:L �v"OB��s+Ƹ@���A�p���"O�i��ۼ
wd䫷.
X��r"Otr�IG�2{HM��_�(�w"O|9��1���@i@�)x�$"O��smNf(��ς�sr�� "Of���%O�!V�x#�]>Lm�F"O�*FP�G�����n<&;�Hpc"O��P �B7?)xi���(=�r�8�"Oz4��잾A�ѦI�}����"O��I�O�
 �@���:j6<U��"O�01vhȦB1���G$��0��"O�DHRg��.uvа$��cul�f"O <�4=,ԆY+F�ޤv^�-�"O8�#�8]\�P��R[>��z�"O|�+�;8is/�,0�e�q"Oά�/���i���3.z���"O��ۆĔ�5���f�
& B�i"O��4�� )H6@�ԝM�^(*"O�и��@̚XsN�kf�zE"O� ��Jb� �.����fS9mA^4؅"O��Q�ڎngz��T%�+G=�ĺ�"O�YږjQ+6R�-Э� Z6���R"O��b��'`�pJ����qbc"O��Y֮ǣO\lq����$O�̂�"O2��h#��Ї�_r�� "O��"�-�&]�d�3'� W�JQ�"O�Q(ՂC�s. �a��z�8�R"O���)�<�\2D_	J��*"O�'OL�x�.Œ2)��
�\�x%"O�����D�'P�(
��&�z��W"ObU�N��1��P����;W�0m�@��b�O��<ɠ�<
�y�ri�e�a�'x��S���&~P٠�
Yh��L�m՟T�<�SU�?�b<�G�݀DF465�RB�ɨ@2��B`߸)=B�p���D�NB�ɵ:)XII�+C̍��G������3��3#+:�Ã�P,��az�BdB�I��؉���H?㐍3����_��F{��iW,�]@`��{\L�U�4�!��-�L���IQ_RhA����;��!�S�O�NP�q��	LaA�т���'&���c@�Sn�!h&��.C��MQ��d0�S�T��
}���R�R�^����I���=%>A�<��fGL�X ���F+l��-1"��K�<�Ef�<�n� ���?�F��I�<Av�G����� �ŝ+��0+F_D�<�q�_������ (`��B�C8�p˕�y�Bh
6͉�L�	�@/>�O
�	�A5�T����r�drL�;.��C�I�J3�H��ĳ\\���B��	N�C�	%>vhأ��8:
9���b�C�I�F��]�Q��%o�(�%ˋ?5��C�	�>�z����4���"M	�ki|C�Ɋ1��d�4��*(�0z2H G$B�I	�8`G*֛=���f�6<.B䉽K׼�e�Ԭ*{�a9�ᛝ0(B�I� ������a(�Q��B�J���4��+?E�䍄X�̍ʂ*@�x�"�;��'�!��U�tt�+��b��!(@�O5�!�9N��	�����r�8`���~�!�$���� v�ҬXW�|P� Z�3�!�D �g\�F�ˌ Q.��aǊu�!�$Ba{���MM]P
	���	�D��'?ў�>-8���]�\��k$c��I��B�<Ɏ���tZ0U��=F�d�dZ��C�ɲ[h�jAA�h`j�-\$�c����I�-s�f��*L�����B �J�H�'"O��D�T
/� 6B�F�ڽ@�"OQ�4Hljp13"S'���0w"OĕZ1I�.O~ڈR��A �	�"O�%Mp��@N���!`"O� �V%^1�be�mܳ&��Y�F"O,�S�D�um�j��Q�T�6�d/�ŞC��M�Β�m6����ә!v���ȓ�������%L�6X3#FK\4���]�Ԥ�0`����N6+�E�ȓO��t���F�n�������{�Hц�=�X�鵫�N6�Ӈ�K9 d���L��{񃄮o��i3P��=sV	�ȓz� �#t�\�o�L���Vq+ �Fy��|B���>VjJ�R�\�v
��y�
Nm�<�u U�`e��oǤ82��C����hO?��F�liPsn��`�����С,R�C�)� D�;�� �g	��{�f��^��9%�'j!𤛀I>V����`&)8GG�7Z�{B�?�dSy�
$0a��;P頡A�TR��*�O��2q/��[�~�*U�&��щ�5?�ቚC���sE	_�~�X�Á�[�JGC�I�\�����[Cf��!F�:N�B�	�
�d�Q��D$ODH����V!bz��d��<�b�Z)��!��?�V��O�s�<ل�Ѕs��+V�T��qrU��o�<qҩ�%��̑�I��?���+l�<"Q*j��𘡆�^���ƨ�k�<������%�
	��G��P�<)s� yz��Hs��8�����Mf�<���'�.M��놖h-H�Î_�<yF�[�4N @�¥F9� fA�<I@��LB�j�΍1[���� ��h���$00� �l�E�$�JP�Ʌȓ:�XX�FܶT�\j��H'D`5F~R�.,^ �@�� ��t�lQ>`�HB�	8Q�Q�ֱ03�N�K���h�<a�����`��F(���kk�(��B�I��z竞�-)�LP�Ϟ
��B䉡_7>-j�� sQ���a��*�pB�I7qWJ%�fjH���%�FiJ�L��C�I�o�}R��wa�������4�*O^�=�~j�(Вy�B�V`�*~�p-�CKQb�<Q����>$.98�N�/�T!�j�v�<��"W?��
��c���o�'e�?�B��&��lx�G��]�y���9D�lrP��8��DC�GTm~q+vG2�O�'�6ZG�D�YR6ϑ�XQ0x��'r �� ���%y�A8����Rѱ/O䉍��K����d`X��v�R&g� 6uxC�I^���2���PrRMR��ODs�B䉵:B^HWIĨ v�cS͐6B��`�DQ���o�NV ER���"O�X�p�43����Z`��th�"O�D:�I�$I|,�a��/U��X�g"O. *�gm��X�A�	*3U\0K5"O��A�>�rк�*��$lv�#s"O��1�G�?i�l��7�)M����xRjRj���O����� �7�0�C��(NgHD���y�d38�Rgŕ�Hג���mW/�y�똞E��à.�
 iO�kr�4�<ɉ����aƾ.I&��"R&9%Jτ�&B�I�z ����+_Ԝ�7ďoV��D)��\��\�B�.��E�+rR.M��x���[��� ���#�	�ٕ':ў�|jt��^�����10@��(�Z�<Y��K�_��"���x���(��<i��NqHD� Κt����pb��1�����@��ΦU:�/�N'����)E(� y�,D�@1B-�,3Nz�1 mߨd��)a��)�I}��G�O�nX���Ȣ��9@���z�����'!"�ǈE�T�w��rCnQ�
�'��s�b4J���R4F$<�l0
�'��aB�SR�����D<��4C���2O���ɃI����$	�){ͮA���'��O29!f���K�H�6�f�2�"O`��u�N?	7�8r��O5C�H���"OH3����"ߌ�xA+[ "}"� �"O�Y��\>U:�YQ��l���"O��X��K�b���9f߽]���g"O���C�@�ay��C�?D�H�"O� ��H�F�Y`u�'h�8jC.!��"OLu�L�?Ǌ����eC��C�"OZ�A&i�$v��%�PF�R?��[�"O�<�eN�����6断U"�E�"O�`�e	)?Z���ۈRi�"O�	�+�da$��ǥI�O� ;�"O\A��$=�T8���Z-D|k�"O������䒶/��`��m�T"O�����T�$tYo�*/��=@�"O�� �J2\�[�-�P�t�3s"O~I�Q�d��5t�F�M�hP�ȓ=�hv!(�����M,G�fĆȓ5���*�$	)�d4�w��(tjh�ȓ
�Nq�"�h�XQ�%��<:��|��7�@�MV���i�D!_�G��-��rӤ��*��X��ӫT[�L�ȓ;����4�Kb��cl��ȓ&TI�Gg�"u	*�(F&{����T�
�$ӏu���d�%R^ ؅��t]p���x],��&�C���ȓi�2y��,a�0yHr�B�/蝇ȓ4�����Η1JB����6.���b_P	[��Z1@�VŊ�nߪ<�=��W6(���Q.̓���P�V��ȓXv�M���ۇ~���rgB���ȓ84xQF�Q.d��/�l	PІ�<�T)��;M<1��,�tVf$��akz衄h͞5�u�+
�dW�1�ȓ�f�!�o�$n�n��l�o@fه�58��S��2������a[ꠇȓW#����EJ�K��y���`Vpq��q�L���]:3�R�)%!������|,��C�/u0�(�)�Z���cǒ-���-;�ε`�/H.�����%�M�dF�5[�!���A/}�1�ȓu�@���W�j��DS�^�<K�-��"t�U+bN[�F��S`&��C��هȓ��+Sl�7��p��lԺQ �`�ȓ<�h\�C�D�A���Oصr]�1�ȓ ;����ǧ;@��Tӯ|����h �R$d�r��%�B_ t��ȓt��J��B]xH� ��͇�@�*�����4��\8��"���ȓ �3A�U [�D1��kd!�Pu�<�k[�7OH��#�ʹR�0���Lv�<�bփO��(jp�T�a�P�㥡Kp�<I%�p�T]�pJ;J4�9�B�<i� ����z�" w��Qy�JR�<��F��L�A�94j��׭�O�<A�lһY�B��G
�6D�f(Y5e K�<��(N�u�F�3�V�B�HH�O�|�<�G�� -<؊�A�8V"��CXz�<�kH{���sF�3
����͈q�<qe&93��E�� G� 1t}0���B�<Y�À�[���p����T &C䉺e�60��U�m�t�:����>D�x�6)���lpB"Z�y�~l)��8D�X9��ߪ`j��1#�:\���
0�4D�����Z�bJF�R5ʳj0N��?D�� �A��1����=�:)��k:D�$y��RjM�!��x��:D�@z���]�Ll�C�?K%ܬ��,4D�,bi�~�D�Cq�X��@��3D�sE�}z�I�w.ն%r�:O1D�� $՚/�?q��H2$B��th��"O�p&@�(���F1U�\h	�"O�]:f��(Zψ�B�� u6\��S"O̸��Ӻ��p�h�_��`jE"O�%�G���G憳S�2$�D"ONAˣe!8��Y�G�'#M��i"Od�;��5Cbi2���+p@���"OV�X��Q.WX܈cE��0bMXs"O��MXp�'�]����"O��mR�&W�P���[��Ջq"O:ICC+��_�A1�JG�y�^���"O@����!ru�L�D�=�"O���qe�{�x��Q�#6�a�"O�0�3N5DIbd��g;|���"Ol�1�$�bz�d)A��$���ZV"OҕQ!m"��sfm��B�"O�i8� ��1���i�߳vq�U0�"O(�y��o}`�;��v�~L�"O0�S��1&p�������-�T"O�����L4s���*P�
�s�d-Ab"Ob�hW?O���nʑt� (�"O����L8;%������dVZ�"O���]T�)8 ���"��"O��9Q!N�L`��ۓ!��h���Xb"O��*�3�B�ڦ�̢�qD"O�Ar 6ZA `�	�0�TEHb"O<M�@Α2-0TQ�P��m\��"O���4��0k�����*�~^��X�"O��cՀe/�,"�(B�UW���"O 4GJ�[Z\[j�V$���c"O�i)G�~ز܈G�ݗL+��"O~��a阜hD�t��)|�Xq�"O܉7H��\'�����J�dz��:5"O�	���48�E�/nX���"O�<I���
��P{C�٠s.�h�"O&L�UƝIb����I+zY��"Oܸ�CL%"ʺ!J4�v�x�3�"O��
#)Gm��	��*��"OV̲�%��D�D4��LV�>�(�"OL��O��T��@�m�g�*q��"O�UIY��~��g̀~vYE"O�a���(ў8 ��MWNI""O�9��hT/D�~�r�LÊ5Jq��"O*�"����ժųoShTː"O֥wJǢ/�0����S<6�����"Oj�U��Z�T�סM\�� �"OB�bSA3��IE�ơ3LJ�q"O��%	E�k��Q�F*�%+�n�2�"OV�`��+r�r�A��p�����"O�Y���S�U��!�X��s"OZ|��( /��S�NR=��"O�y��ǉ�n]���N$a��U"O$8�_#Uh�M
�mJ�k�1q�"Or��ïi��T�Ҭ�7 �x<j�"O�5�F�,-�.��¢��Fy�"OJ�$�5�@I�#�,yސ�+�"O.頡��5\���P��p�uR�"ORD�edJ�~S(���&vԶY�"O���O��ص�,�/�R�Hq"Oȱ`_53\�-{��V!Y�VHK�"O�y��E
d6aɗ,��"px�"O��@@��cn�y��kܩ���;D���po�/S ��X˘&��%�b�-D�
�BO����閌�ȡ�@�*D�� Q2���)x,K��K &(`K�"O~`���1���{ti�'% `�y�"O,V�Փa��=�4+� )����"O̹��'\0p&�Մ��$��ʖ"O��2A90� y�8�ϒ|�!�$.,w����(�X���U_�!�$�d����d�"#W�E�!���'���P`��{��-)�Q�!�d��(UrX��F�P2$E�4W�!���uz�1�5�QZ���`$ȑP�!�$4H�`@rO̙@	.�*�b�3�!��3@	hS�R$9�:ёSoJ&G�!�D�-J�f��난eΐp�ׇQ:t�!�dJ_��E��r����g׮!��ײ=hyK�	�.�rъ0$�+!��[1�\�i0�6:&�aٱ�	�9�!�D��Z���G@�	;�$;@���a!�N0W�N�S��K:c��u�֪Ġ	.!���q��01J�8F�\�Pugǐ,�!�Du�^հ5aW�-��H�E���x�!��7���P�r��]��_�M�!�d��u����BϬ!2` ��N��j�!�D�3x2��%�|��M6+z!��4+�̱���5��Tl�:�!�ʯq�H`�3\��q`@�U�[�!�DJv�
���#5B�i�����B�!�d4d1l<�s�ҕC=�"JD�{�!�$�r2 ��$&S!D@�e�1}�!�D�k�H�@�f0��K���Z�!�D�&�TI�C�L�'O��J�!�*J�����p"��/'�!�d�7,�E��TV�1+�k�*o�!��H�cj�A�@�1u�e*j�.4z!��<��W�a�8l�{�.���'���:U�E;!�g��#����'老�%�5(�)ď��m���j�'�*-���Wb�A׬�=;\i�'~J�a�k���b�"2�i�'�4x��� ~\��CH��
�'�Z�S0-�j�HI�gW�:"O4Xr�Ȑ+I�Y1c�7�@�"OŃ��2^�RP"���$"^�:�"O(�0G!�
D.xRr J�d'(��"OBD1�H���0��L=9& ` �"Ók��߹[Ad����űw��q"O}��$WC�HE�m&���"O��q���v^�*���?�M�"Oj5A�ߡ}Hh�qA)� 2Z�s"OH�+�1�\S��t���"Oą�����7C$�2�k����+�"Ox� ���=!�a�(60����R"O�`���t��E\/�ZqKr"OJtz#L_ ��,�f'v�Z��"O���ac��2&A��"qv8� 1"Oą�DhV+Y�h�����<jDk�"Of�Tl̀{��bAJ88V=3�"O��4.�"=9a�H���r"OV�W.�^��:�H
�:����u"O�@ِ�.~  ��4_��D#S"Oɲ��F�u�`2C'�*7��#�"Ozpc3���l`�XR�G�:s�|��"O,��%�25��R��:^��x�A"O�A)�'�	S^QbE!;f��%"Oœ��iC�t��
WR]��*�"O� 2��e�&P�� �JjSt��"O ��f��zNn�K!�M�I(4c"Orx��"�_"� +�k�;f>,ʂ"O,�R��Qn
R�rb	Z _"쬱B"O<��׳'k��	ª�>�� �"O��Qa�˽+��L�� ��
��p��"O��q+�&AЀ�1/�`�aÄ"O\�:�̈́�K���S��,r����`"O�1�$"�y54���
lm&3�"OXZ7�T�4�! ��f2�"O=q��D��$�u��(p^Fi��"O�Qg
ь_�����9H~\��"O��R$��	'��YA/�ƅ�"<�!�dD�|b�qrP�l���ҲE^?~�!� 5����Ŕ��OL�!��Mo��eh�?K����@��!��]�)��o]4�^]�Q�2|�!��J�����!E�k�.9& ���!�G�0�3΄����qd]6ix!�";@���3m��Wʕ;T�ƿ0z!�$� U_�p�U`
Ն���Ŭ8x!�ηe B�H�.
�x��Kҡچfn!����wMR�A��T�"tK�<bZ!�ґ
��83 N��E��8	��ѵ,O!��9$� 8���/lyb!�dDK/tW!���5d����C��Uk����ˡ-o!�3r���/R�DMTP"�,j5!��L/&	(�#B`�&B�y��X��!�I
M�1;�
Yd$X���ĽZ�!�&+����A叁� S�e�p!���3'P�+�������t�B�Ah!򤝑H��JSZ��-��W/r]!���ghp;����>/�Qr ��X@!�d��U.�	 �#m��2�OJ�`�!�dG�\�d'�NT6\j��0y!��+5��	�4@H>
S���D�9cT!�DR6�ؙ�"�ߡ&B��yU��,!���a�(��?)�<;��_mw!���0�I� ��'���BZ!����j�K��(If�PHE��|D!�d��rax�c�N�&��u�0툞O!�$<$ux���,f�T%�$,��a�!���WDpYQ�`��0��hJ�Kެ�!��EQ HCm@8��Ѣf�5�!��&6'�0b����SlhY�^%�!�d�;�4��� �.$��4{ï;!򤘅nlX	&"����y��/�Si!�dF��"q��1Fʒ<��L�5'�!�dր7���+�I�_ph��@̾n�!��H�'GT=���H6Tx�a���y�!��`4�� �gY�k>5T@2(�!��+M�!�V�l�~��rn��t!�L���Rs$]��:t:3@"A!��)K���3F0�49� ��t�!�DX�s���m����&v!�S=�l��&g&�i�e�BJ!�˘Ŏ`�F��$GT�h��<z�!�$N��� �#�@�e���8�!�$_�������� ���33���'��	',�=TzhȰEI1����'KfYHď�D�*I0$Ӱ/�d�x��%�0l�`�`� ;)\!��]U�<�7&X#\�|�7ꞧxtJ%���J�<��h\�0;F��)�#u�|ru,H�<� ����M�~PY
��� d^��q"Oy� ��"��фK4����T"Ot%��cA'��8
�m�%Iuʡ!�"O؜�!�B��U�aB�>q�c"Ob%y#�R�X 6��GG�tn� ��"Ot(R��5l�H`�u&�}���2�"O��a��A$�Hѕ��x"�a�w"O����#S9���f#Z�W �t�R"OAQ5�ٟE��ܛm��Gv�s�"O�( �ϳ9}��Zd%�3]�r�"O��I�FH �͹ Eƹ7g.Ҵ"O6`�EZ)�n�X���Xc��	�"OTLb���d	����&q��e��"Ob��iӜ;e����g��8� �j�"O�e���_]�¡!L�*�("O�5��]6#z�+f��*��P"O��2���,<�R&ڸ]�Pj�"OJ�	�Q�lֺlP+G��3�"Ol��_D��Ě�ӆ���"O�u����@�0�$Α�-�d��5"O<<� T#���am9="D��"O�@bX�"d�JCF��)r\� �"O�A�GhӽhF�Ƙ"^���"O4P�ˋ+m\��qe�8�䓇"O0q�*�$$ԖhT�M:���Hr"Od1q�V-!�������?�<}3�"O&x�`O�p�nI��IG�| �"OL�#���!G��(�B�M���s"O���ϋ^S����8;�,��"O֙2�n#\\��*��:� ��"OY��IJ�ŲQS2���_��Kc"O~�S��B����P��('��e#�"O8�cb��^x2C��~�]*6"O((� 5"��)��oB9�V�Ȑ"O���0	�V=D��4�z�H��2"O�Q��K��Ad �I�/��W�p�9f"O�UB0�5��iB��T�����"OX����"Lo�-HĀ�' ���v"O @�F7|m���8��Py�"O"��E��XJ�"QH��K�"OV݉`�߅b���;�ȏ<�JT��"O�X�QB�	/(��d�Yd���"O�}���>f�Dy�PS�Y�,��a"O!@�/~�����\4y�,��'"OȑQ�TC.ya�G�[�x��"Oj��Q�+�J�j���&n�q"O�fU�}�1�I
� ���&3c�!�$�A��Y᠋�0bVX���/{w!�V&A;C³BJ1���Q!��5
�� �b �+`rܱ��:!�Z�Du�Ċ��5C:i�gA�!�D
6&M��gE`,ȖET!�D
R�zW�ܐ6�t�!����!��׶Z�PuR�eM� /�]�4�͍z!�N'R��J��<��"gA�x�!�Dε|���Z(&�jd�&cN�n�!���I�6��%� 4�-"0CS�!���@�SL�;
�=����:+�!�Ğ�<3��Z!�s���0n�T�`"O��P �I�~�h�4.�]*(��"Ob�PV�I2EN�dJ7F�FH)P"OT]��!�&NpZ�Y?S���f"Op���d�pM(�Ǐ[{�9""O@��7^}�)��D�6s\��"O� ���jǄx�!�u.�=	���`"O�s�(?����ucI/N;(�;v"ONX��c�;�b���'�wL�"OP�ZwK��o�p�����A�L�T"OF5i%�(/��%�����"O����b;ܭ�!Ł�a&XĚ"Oh�y��=���fM6!��1"O�|9� >��1#$��\/��""O|����8�N���P1r�CV"O��#�;:I�4��.�=i���"O���'
�?<, ۃ�\|q,�"�"O&����۬3��Itf�	h�t�"Oȹ`*�V<�C�߳U$��"O�H�g[�]j��%�3H���"Od�J��-2��2%��*@T�'"O�8��zEP���=z4���"O���3d�����n�!jm�w"O��X�@BעMSwmW�)a�� �"O|5�^�8G��0O2cz���"O�P���J1;`"�:ԫ~54�Q"O��˳fL�i0��k�)���� t"O���Q�r�I(U���b�)�"O�9I��>+��b���/|����"O 	�ʕ�* j<j���*���"Ov�����<-�h�BЋ8P89c3"OV�C�@�I`5�W��3COh��"O0����N����B��J����yR�\�ld� ��FZ�u�TI�D�R�y ́S�J̠��u5�4 3%���y2O�i���+��� kdP����H �y��.m/�4����k����ǒ2�y��O~��8���4��y�cF��yr� ��x��ϋ "�2 �g<�yR�[=m&В�/��me���G�ǳ�y�l�/@�n��F�k�:�w��yb"����� ٢jl�q��:�y�lӂ$ƺ���O_�f�H���Σ�yb��ZT��#���6����,�y�U�UҐ{��ZWg��P�.�?�y��h�'��TA�䒂���y�&_�5��|��� F�*�PH���yB��<r<�I1raϵA���CE��yBF�c�D)�q�-�fҁ�W9�y���#H�0@�.�4bҤ�B�N��yR�ǩ2�P�dB0 $d����y�=��x��2頑8�G��y� �.i1x�eB��(p�h���y��Ә��!KĘo��ph�h95�B䉂$ ���ۺ$S�H �\��B� ���R`aC�#\�0"�,�OB�IM���&�եv�a�)��gLB�	,���cиu;(�f� �e�B�ɣ����Q�Kf���^�;��B�$O�0���,]�Dp��Z9�tC��I�T1�-�+ ܱ��icf<C�ɐ<���ҷ�V�\���	��Q�>C�	�)T�X�Tv��
%ny��B�I�0���{��FJ��¤�}�rC�ɩ E�!G��m�]$M���C��,v����eP�(-��w
T~C�	�A����jJ��A��"(rC�I��u��*��Hl�C�`P�TC� 4��|��a�Z��w+P�B1�B�	�+��xyLY)1����.�}��B�)� �d���TK��1o�=��"O���K����L��l��/�0ɘ`"O5��/޸�R�k�O�(�F!�"O�8�$�[�\��q�Z�t�<�u"O��a󀆂|
�˃��|�*u0 "OĔ�pkW�x*�`z"�¯Q�����"O600�H�ܬ�L�y���0"O����M�w��|��P|cRj�"O��BRh�,Z�O�LV�$�"OҔ���\�b0T{b��� 8t�p5"O�[�����(Cq�(�=h�"O�H C��Y��K��,&,�`F"Ol��E�H�r�J;�ʅ�E�w"O<�b��"5��"+��V�l�5"O�= P���zk2�!ȍ/4$V\)%"O^�k��l�J��@&R�8�.�c4"O����E�
����`*@�9�,=�!"O��+v�5���;@�@�q���"Oި`�OK78��,��i�����"O�10R��&p�d��+�0�2��"O�ik1K	F:��1j:טq"O�@A�V#� u���	$O�:�"O ����,	Ҽ
�G�i��L �"Od�EE^�N�p�)�&�a���@"O��ˠ���u�$��/:���)7"O8�
���qcN�`K�,5���j�"O��B���x>�xrb(�4�\,� "Op��Po�J~@�[���I�H�{B"O}�`b �+�,5;F�,1�6��"O��	�!j��9�N��W�����"O�E(�B_"6Z��bv��a��0"Oz�*2h͈HI�4���ߙ=�\\�"O�2���8y�]���
�H���ô"Ỏ�bfR�i��/����b"O A� DO��f����<D��Y�"O�MAU`�=�*=��z@v���"OJ遣��k��%��Kձc5f��"O�lА/E;o�@\
)���ev"O���rl�=R��
	���"O��R���&��gفQ��|a�"O�Ea#&��ha&��z�΅�"O�3�߇?X(�h��	1{���z�"O�m�r��3!v`�z'��p�tI��"O��b��
q��=���'@�2���"O�|�T��19�����Lˆ,��	bt"O�qx�B��d�v�Yu�٢d�0|�"O��xc�ƚ�Ҥ��ɗ 8��$��"O*��p	�	*�![s��@Na��"OJ�J�d
�
,��#G��"b"Z��!"O��X%��O�hᣲ�¿x
�M�"O$ �se�W�$���D¼�`�u"O�J%4>���!�R�|���1�"O�X���4d�ě��վ8�ڑ�'"O�ɘ���#t1��0fĀf��,p"O�E!�B�$L%FJ �3O����`"O�|{d#C%$K�	���<=��%��"Of!��&�)C>�8���O�K��P"O���h��	�x�V����q�6"O�+���2����F�Yg��`"Or��鎋5���xgS�|� `�"O��3��I;��S�"�!9$"O��єaQ�+W��;s�*�37"O����7hV�9;��,;}x��"O21)�k�k	fU����Sa`�K�"O� 6(�̟|(�,QA�u] R�"O�X�ބK]:����53]��!�"O�m��.i��f`����)�"O����& �v%�/..ڼ�k�"Oj@�����tT6��QԜ|֎|+D"O����%�1ln|+�/Y�@��L�"O��i��MA��qʢ��@�´�"O���ƅGGY�y��Ӫ\7>��"O���04��Kgg�$�ʩ�"O�8jF��F״ݐ�(�A�Z�у"O��i`��9$'��I�G�j�F��U"O���F��LH�)��[4h��e�G"OdL0��� &d���
?�U"O��Z�HL�άZP�DD��҂"O �X�l)RB�a�5oś)-����"O�Q�I�eRX�b��Ԅa����"O�P14)N�<I�V@�~P!!"O�Պ�LY(�TZ&���nsP��c"OL���T.nv�Ȧ�Ҫf{`1�"O(�ҍ[�*��A�S�*�����"O�("�P���A���ڂ���`q"O��#����Z���TG��q�JUXc"O �!S�_�4>���#9榵��"O*	X�G�-�<���F+02R��"O<P��A&A<D�Q&�O%n�Z""O��`b�N�_Z�aJ���T���q�"Or����G�QQ�!�����"O.@ł[�t�
�����l)�"O�A#h��� ��FM4w�jC�"O&Z7��m�4�wO+/غ��R"O�z�@�d2�,K��ɚB����1"O����	
:�૵��� a��"O0}����gnΘK��ԬF� �D"On�iU��f�*��[.���	A"OV�"VO<������z�D�p�"OތGH��Y5�8[�%���JD0"O�,�4CC�P4��&CN�[�8l�'"O�Pئ�� ��јW�<|")I�"OP�HQŇ#x��j`�
<n����P"O�AJ��Ÿc�":�֓L���(�"Ot!��H7#oPI  �X0m�T+�"OЃW��pv���Fx�$�(�"O:����#FtʜibÌ�}�
��P"O���S��C�t�Q���
���*O��`
�\QDي�Ha+�9�'�d��C�b:�]��J�/�:Ua�'�D���/I4V��d�#$Ӫw쒤b�'�FRN9P��{�X���I�'x���& �\����f��Yv~�S�'���Kp��2��;q�F�LR�'�4� �ׄe���
�7�Ɓ��'��[���,�͙0�ޕ��$�
���y�k�B>���e��i���̼�?�-O��Ğ/0^�ha�HâI������N!�S�J^��6��I�P�1
�!�ĕ"i�-��i���#�(�=�!�
}�ukWd��%��q�4�AR�!�ˤq��ȖB��n��L��>�!򤑓�U��,+{��A����=Zn,��_�>����׸T�TDC�9|H�ȓgԅ��h�^j��DK+�}��qQ��2F?�>��͍�\�tT��>��u@�œ��i���р^2��ȓ
��0��,ȌEƬ-��e�?�u��S�? ��D]�f��d���7r!�"Ov�5�N�J���y�Z�[�81aE�'��Iş�)��!@4~EW�X�4��0D�G���=-nW�1u�* RUlT"���6"O(���F�pj��ۙD�����"Os�|n�ЂI�5����V"O�� m-F:@-F�OF��!"OT�ō�}w�	ZF��+!"O��0��g�HU�@B�?Ք��S"O�H��]w"�#�`�.7+��C�"OR�gԤPc��bv�\�=%@�"O$����8X����Ûz��8I"O��D�ȧ\)�a��^�.�i5"O�e
�7��t(���0�B�"O�D˷A3WB6����
[���U"O �b��[2H�B���N	Y!�'n���<�!M
�z� ���CI�l�K ��x�'6a|�jТj��CD�L����"2aʱ�y��h�ĴJp�N-V4Q�F�y
ؑJ<��D�������ybO���:���gT���+�y�jS|s2Y�ч��.�|�2�`L��y2,	�]����L"�����ګ�y�E�Uq)A�%ߦ>�|CT���䓱0>��(ӈ]z�3f�\[
$lń�h�<������)x�M�<�2a��N�c�<1�O��s��[("�<̙�j�]�<)����,�҂l%∍��,�y�� PB����٠?�ЙC����y���bWР�B�F����zi���?��'��1�C3]f��ٶ�� 8��e����2�O��S��H!�|Y��A6S_h17"ORU�U�X�^���ˤc%q�"O2�BC�1O�Lu�B�F�s�"O�8��dߥ��8 �A-D/�\��"O&(��2]K�=�U�-#@�'"OԽ"��W<�<�QddÂ*Έ�c"O��j��Q�2E^|kT#��>�ԍ�"O
q)'gݞpʰ��<mv\b�"O��ja��r�i���!G`> �#"O�� +3n�uK/�E��q�"OT��#	5�Lu�#��=�R"OX�HUEA(5�v���ǝ�L�e:%"O]����7jq�qy�T����(0"O:��r����ї�E8( e�|b�'̪�B�_wr�P�K�"'�����'va��a2*��́W2D��'X���'I�@��̀Wd-(���'�X���]�|*D�Jw��b��*�'}�9��\3U~x9 ��V�|K`$:�'��)Q��
mWX��v�G�c�N��'Khl��c�B���T�[#/� �0�'m^ʄǄ<T;�T�1y�88��'PF}zfO1k=�a#_3Y/H�"	�'�*I�3�	�&�HQːUf��j�'W�A2 ��/�8]qU�֕H��,��'^ʨx��"?0X���Z�LI$8s�'y9�P(J�_bN���

L�ҍ�'�� @O�"�����Ę�H��Y	�'	��8��,�^a�U�߁X�����'`\�ĕ<G�����JX��t��'	�c`���rt��6U ���'V�D#�KO9rX�ơ�"_T<}y�'5^]J�!�\Vv��6ɋ�^���
��� 8���KT!h�5��-�p�� ��'&�,���$���&�.U��3�+D��8"�ˠOt����W��\��T'D�9�A��M�pr�? �X᪣*D�����l�>�3��!i-���d�#D��å�C�(Ȧyy��S�q�]�T�&D�P#6i�Ez���v�У���;%�%D��1�_$aQ�@a��n�To"D���ƨK,�h@��
�(�N��Q�:D�`�e�9P�eeȷ4��(!�;D�|S�d�W@h[b/��^p��H��;D��A�IÒ%=  "�X�5Q�;D����j��HI� �4�[�Ei�!H�,D��#���y`�Ы��%N�uqd�)D�\��A�)7tXS�E�%�J�%D���綴����߱���uß�s�!�=* ����!����l�&f�!�D��Ke1�##��d����)s�!�O"�8�q�ܫO��k���+)$!�$��p��4⥣��=�� �HY�!�((�"�S+
>|�d��H�X!���$r���ig��ke���p)ەnN!�$[!�ucᢚ9}k���a�¾ 0!�Ā *���R�����r���\!�O'U�}�U�J�q����! !�d��C��k5'�8ּH��А�Py��!1,d�7��OvPj�eW��y"�C9��EB�O�u	����Py���x��|ZT�� 
��D	��h�<`�H>n�����+.XȈf-�}�<�E�R�`{Xp�|d&A�S�J{�<	Q%��1O %r$�T�b`����u�<	�k� ����Dd -9S� )g�n�<Q��6��Mۥ���(�S��s�<�Ě�.ݪ	zv�ɳ�U�D�X�<ɲ�%d�ص���2:���&B�_�<�b�R�	�)`�I1N�)��/�]�<A���&	2x�"dʘ_�P�aETZ�<�	R�n��7��.�p�w�A�<)$�W�@��,K�#͛{�
�k"�y�<�T/���9v�H��XU��*o�<�+�-��a��w���ঘd�<i`d�#��D�'�n�V�p��g�<����+�t@�E�&UHC'ʜe�<�r-� Ɏ|�c눨$���BG[�<!�.;>� �� �/'xf�z��U�<�aEK���D��k
�y������Z�<I��x-��dC�,rzP����X�<q�ɚS�&�Y D*8��Ap^T�<�v
ӗu�<$A$�Oea~�#���S�<�"摾Sԅ�!�A�E�� ���P�<�á�|ِ���[	R���w�<��`�,��H�r��C� s�<�!��6=�1Є�X/e*yႡ]l�<Y��Z���p[��?�ly��o�<��پ*)2�룧VIAb�Q�h�<�W���a�.T#6�Ȁ !�e�<�d\Rm�X�Ă�\`x�@��i�<aq��13�T�ӭǫN���k扞e�<5mM�xYr��}m��!�`�`�<�#�� ="	S��*2U0I���[�<QA�ߩI��F*Trb)��ΎW�<)3'��`l&�h�M����V'@T�<)qំ���Kচ� ����J[�<� @��F P��n\2�/]p0m�v"O l���TS��6 2�XC"O���ىjz���&a�P�s�"O��e���n�t��a-���8��"O& b�҉!*|����J��ɪ$"O��IF$�1�a2� ����F"O����=�@�@����pU0q"O~����űk�L��咓���"O�M�����V5�%�<,�jQ��"OhU��4mK�nχP��	�d����yR��`ﴅ;`�W�E���"�GK�y�Ļ$��Xa�[�<M�h��o�<�yb�&�-܀��eo
���!�'��䢃�^�;x��j���]1�'��(��@�b�z�SB�J�FM��'�`t�ެ'웑a@L���	�'?���w��3V�Nq��.C�8ܩ)	�'���y6�>TJ}��!**����'�DY��I���$)!%*(�4	
�'Rn\�ơ�>&��#�A�8x��	�'��I8�iP�,!�-��휱[��]c	�'נ�z0���m�+0&�
JV0��'�X�E�����y:&`K?�90�'�Rlb#��_���i�m�)HB�*�'E��3B<�,IL��x�Z�9
�'��%zViZ���a�o�q�l�
�'rT`kQ��`��8=\)c	�'��e��gM�b��u�`�$:���'�n�dE*r_ �h �ѻ#�Y)�'�(�e&�p��p����s��}K�'4�ʓ/R)7��u�A͌< �ܭ��'L�@A!@�-��Wa�4��'�(�P��Er��g�)u:
�*�'1���I��Ι8 �tJ^���'ɖ��c�:	d`,+
7qz��'�n�`�!� $���1򂄾x2}��'06����'f���Xa�(�$Ĉ�'7��l��BЀ��EeU�~x�E �'2x���ot` �1��2p�(�'"y������DU p�Z�)
�'�T��
~������)���K�<ٕ���F�N-+��#!0p,�ħG�<qQ�{F�XP�M�Bo*��!��B�<�@�Y�W��PD�D�mv�Q��x�<�S.�,?�̋�� K�|�
���|�<Y#��5xA�3�&�h\�
A��t�<��$��8��ԇ64�F$j�O^r�<�z������
�8�t��m�<��V1!�l��6$_*$>t4�G�~�<y�n�T�Nl{ń"s��i�\6B䉼t��`�D%C�l���S�$��+"B䉽&�x�ˇdK"Y�f�������(C䉺����@�~@QiW
X�B�I�4nr�p�aT�J���@�_L�B���=�1dP����:�X�4��B�ɕ@��Y@��4��|PB�5:��C�I� �eE�Y���re۝M)�C�Ɏ0� �s��#))4�Zac�~��C�7*�()1!�aq�4h��<KpB�ɂ4~�0� |YBj���dB�ɫU��G�Y�#��d���BB�	�G���fi�Yz$ӣ	�o�:B�IOA�a`��L�%x���nüB�I�i���v�I�"����OO�B�)� �jp��l��D��m�0�^ J�"O|���}+���S�p�6�;0"OPl����,�m��nݞm��L�f"Oj�Z'��<C���MN?�J�"O,�p��]#*�����,��X�r�IS"O|� ��5�.���X��"O�q�MWK���E,�"А�"O�,��&��5&�3W�-u��H""Oڱ��'K� ��<��Q2"OP��W�e$ ��ޚ^�ތ�6"O�D���ܒ���oz��"O�p��C*J�,#�jH�B�0Xca"O�лa�Ǹv$@C&i�X��E�"Ob%�Ջ��'CZ!H�!Ա�"O����H�F]��EO�8�ȅ	w"O$�@���-r���CB�>
i�"Ot�t���E�9��>$J�K�"O�q����.�J��� �A[�"OZl�O�R���;	��)ѧ���y�JT�h��<0%�
�n�p�f)��y�F܍I�΁�� ��nO,�ũ'�y�&Sqz���/S�b������µ�yRb�=5PlscÕ�j�|2�$��yR�Y�7y�D�S�E�_��]b�c���y2
��_��%3E�	�F��b��^,�y¥7l�F��5mW��h���2�y2�/=��s�-�<r?����4�y�UpoL4"��Ըn����"@Ƃ�y�4<g�0`�@I'�,�z��0�y�hYA;l��ő}��e����2�y�A��D���d@��w�"=��a��yR��$-�Iw��xY�t��e��yRk�+ �^Pp@]�X���,��yrb�1��'d�.y����y2�
�=�	�B�V��UY�[2�y���꼹���Gl�lIp�L�yR���p�<��F>wg� (��y��>!,�G3B�l ��
E��y�ֵW�<+�i�6�$ ��#[ �yb V]�Z��ԭև+n��0kQ��yR#]�-��̲e���t��T��y"��&�ш�/®������y���R���k���(M���*v&�)�y҇|) Y���|#�qnף�y�L�5c
��`h ?�t@�ʝ��yb�����p��	�:4����T���y�某'����%A������J���y�fJ�~B�s�)FzM` A��y��U9J�@y�Cg�f��N��y2I߆<��#!��qOȡ�5�[,�yB#Ɛ�0����x	j\�$g�=�y�!+Ha���wE�q�@� �y�n�S�J�Kd�H$B�D��S�H)�yR�J��v�G�#=��Ը�׷�y2m�U�bH��>?t��dK�>�yb���4���d��H�h(�c���yҭ��#'�I�ф��~�A����y"�=Q0�����z��Q��	I��y��75t��i@��y>h��b#��yri��P�*��.��Y�N���.�y�!�>��E�7N�W�T,�Qj���y��n�����_�K�����#�yr镪nH�Y�`֪Jt��E���yb�Dc�=��,��<S�q�E��y
� �D򁯙�lN�0(�&��>�@���"O��(��'@���P�H�2�6� `"O�X# �QP/�T�SGJ���|�u"Ov�x5��:��q��8�Aˤ"OPbR���`��C�T�:�0�˕"OVL��q�d�U��7dq�Y�&"OE��*�+��R�C uYX��"O
l��c��-xi�t�����I�"Ol�Y�&ϋ�X���.N<���b"O.H��͙6	����完��P�""O� �aI@�lP.8��*ZlF�#V"O��a�*�c��ɑ�a��L�t�f"O*]jc*�[,���d�=pkz�B�'ܤi���%��c0b#/@6Ik�'L�aB���/(���g��"I̩��' ��� ��b��h
����%d�\�<9�%�&_��VɆk?0��2��T�<IĈT�F���@�m�)�6t0�+�y�<��ȈI#��0���<+�2���(y�<1�a�C��A�I\?��DY��Wn�<�g��W�0�0�P�U�)���u�<��\7%@H�y7��E�N�8��M{�<IO�wȢ����v�yX�Ns�<a�m��LX �O�4V00�`�Rm�<0�#W"DdA�@��{����@�f�<��^�}��$q�nܝ�&��.�W�<A	@3<#0���Tz� k��CT�<YGa'K&*��Bę�?8VH��QN�<I�n�*S�]��
�	44H*�!CI�<Ar��?��-c��V���%*�`�z�<�v�*�V���ү �����Q�<)s��`w��q���}��Qi��u�<YA�B�;�Ȁ���]_n��tf�V�<i�F g� #LW/p���WjZX�<�ȇ/\mP�;���+)��p� 
�W�<Q
�'j
^-����_�	�1BBP�<��GO`Ű�i޲��%ˑ�P�<Y���(����C��0���F�p�<Q�f	�
���$��&2!ؼ�ℊp�<�V�@#A0�3�f��t�0Pb�j�i�<!�kS���^83�{�J�d�<y��I�*��p ��V�Z��]b�<i�ā��JU�qQ�B�����`�<!�Թ$ ��Iu�܅S\���5��\�<����`7<�R5Lӄ[]�M�P�@�<�'ქ���"e��I�|SF�v�<yGj!tCe�҅w�6��sf�u�<Iī�M2�C��y�[C�G�<A�Q�@`e��
^f�3��R�<9�0�`e���h���B,_|�<1&�QF���c�����<$��Zy�<��lD�:K�h�@U9z>0��A�v�<)$ϓ�;$]�1c��U6d`�r`�I�<�jO�K���� wKZM0�i]�<Q�a��*�*H)�ͺ:�hV�W�<y҂�'2s��1Ue_�`�UZL�P�<T�K�C��i�gJ//�ez�s�<��K���V�[*,$t8� �H�<au�Z?w���Ztj�"Ê����D�<����YwhA������ئ��|�<�AI-yު�j��	�ZB%Awc�<a�mɳGX�tBa�-\���Hvj�\�<��g�3�vP���+�ę�7�M[�<Q��6\�AY�a�{s`���ǜW�<� �S�H5.���u`��A��)j0"O@9��+կRN:��/'	�X̋�"O6��D��_\|���G8w�,�%"Ohl24�]�bWn�BS��>L9
x�"O>	��.ѰqC��a�W�Z���!"O����B% z@@��ϟ~L,ɘ�"O�)J�C�=��!fj�2\G�P�!"O24 �7/� =���&Bj��"O��R5�w��U��

m=@1�"O� �˖	H%��H2#.lų�"O@��%.oӪ�٦��d���"OHIҦ�1{> �2���>g�0a�s"O��9��Rxt�,1��5-4�[�"O���b1�T�f%�"y�.p{�"O"��a(Κx�@����K���p�"O����T6B�Y�G J�<��"O02��Q�\�89b@�:QR����"OF�X����22�£	N��T"O"��$ �<����: U�@�"O�1zdȁH4�Aˡ��49�X4� "O�Q��/ȖT��@C� �8�|<P�"O�i�4�)W�>����Ϝ%�м@2"OP����]RvY�_z���B�"O~�#%e����0�^�^�0��D"O:�yql�
MRSD�.��
�"O�|�Ɔx��ta�!5|�:"O\��4�Gd��r���e8�#�"O�8C*������:m��2"OH�J&j�5	|&��oV=NvM��"O������R	,q�r/�'Ct�"Oh}j�����h
pIZ#z9xr"O�0HUJ��r��`�2f�~7�zW"O�uJ��PH^Y{�&LN+.䒵"O (�ReFeq�I���	:$���"O�E�����@�teHL*�"OE�T	�9)�R�!A��0i�,�`D"OV��c�G9_��0�`"Х[VBK�"O邂˝�Wo6E�B��|b$�*a"O@0�vC��. ݢ�[�xY��"O`0�eɄ�;�d!�5mE�{=��"O̤)t��h��HH3���i��1["O���7��12`x�FkY�^�4��""O��i_��U N�Yv��%e(�y�	��W�ْ�,W�<�e�̬�y��Ӟ<e�v��T�D��G��y"�!)O�=����Q)L�4��$�y�e�:*Z�$�5�֡̮YXg� ��yb(ܬD��!e�Z�"�(հ�-N��y"i�*Z���ˆ��	��K0ƞ��y��]{��Q���-�<<p�I��yr�ܷAL8��Q���x���+�̘�y�@�-��q�@�^�t�F4�����y�[f�v��!,lxVx��"�/�Px�i��z��L�w2��@Ό-Q�8���'{n�8�CޜAa$ۥ���B	�|0��x�ؖW��"�M̷_r�Ⓢ[�y�)g���b��P�ShZA����y򇗹 ::�a^O&�e*����y��<rQ��Y���N>8D�'H�y"�1t*R�$#ʒ5�M{���y����S��\����]$�F,Ҩ�ybbG�ll��S�~``\��H>�y�:/BI�G,�:	�)���yB�ѥQ�n��"�(}�x���5�y
� �����Cq��C�J�_F� ��"O��C���-+��{�E�=BLPA"Oĵ�Њ�
dx�aB��$� {D"O�i�d(�9a(Thf�0.|U��"O�bECۯ7J�̒wɜj�Ȗ"Oh����6lM�m�&��3O,M@�"O��H�+R)g�)$��=7?��"O�`4DKxB��)�	�,���t"O�X��Β�fI�ɀ{	,�s�"Oh�PaN�?��Pw뜦D��A�7"O�=j��R�S��t�/Żn�j�"O�u�2B66�"�c�&P���B�"Oe�ӝol���"Y�B�l�"O 4c��ދJS𬁢`$(��8U"O�6O^,���Z�ŀ�U���#"O6��qԆ����'ĉ�(��}��"O��@�ŎSO* �#IŐ-��"O1�b���0�t�rc/�=����"O�4cDڕ*��P9WW�(���"O���c��.(a`�/��j����!"O�e� �N|l@��]�u��Hz�"O
���
�Z��%IϮu��ACv"O��a�O�0�a��6K0v��yR���5P�
�Mܽ2���/N�y�T;HԸ)��b�tq���	1�y��5�Bmap��b�fy�(Q�y"+C!8�\�e"
�#����G��y��/]r�I�	m��p�����y���y�ꉙ��/y[�,ce�ļ�yrh�(0~�%!Vh�s� ᛧ�T��y�n&�P�-�'`s�aɧ���O���P�-i����h�(����ϐ"�!�$R+S^�*����r��âe�!���i�&ȹ6D�X@��K��� !���
[�4��u���`��(���@
!�<5;$�R�v�*�hV�d!�$�W��ٰ��Ҹ,ؠ�ՐLM!��B��3������m�fC@c!��	���=s���\F$�hbK0 !�DQ_��Ee	='��S2ȅ(e�!�D�Z�i��K�n��X7M�;5!�$�X�@�-a�Yɶ���'.!�D]S���h��F�jM�Y��Z� !򤛍VٲG�MiAl �!�	e!�Dʃ<��h��@SN5�AD&�5�!�D�7gr4����nx��VGJ�HX!��hz
�#�*�4F�@�!�R!�dڦww�T�b�0�(4��!�$�/T�}[E�T�}E�5�fm��!�$�[I,�H �p6�y@K��!��s�I��M�s;���`�N=�!�Dʷ�tcB/G�cPX�Pa�ˍNj����	�P��pš��T�p��Y��B�	2�1��>C�캱����B�I�k;��*$-ßd��<�"CR�M��C�I�<�`R��
���/ܟ,��C�ɪL�
#���''�X��۫A�C�Ɉu#ƴJ�$C3C�=�G]��C�	�SQ\ЉwI¨z���`�F�$��B�	�!��U�Cǲ�N�IS���sϤB�I�4��aR��ܫ�*��G֔c�xB�	�9u�|i�1au���EC�I.�����!�W��(
S�;@��B�	�4�YP`eػAΎ9T�A��C�)� @�h��;Τ��Y1GhT4��"O��ρ4�E�ԂÔ^xҔ��"O�e+�I�0a����Cbח^u�%S"O���)�pv�iS���sP����"O�E���_eX`�����8KӜ-�a"O�$�U��$7��+��ە�V��6"O̙c�)i��y���+�d%�"O&����ǡeN@�膎A�O���"�"O�H{��0-*&�G�<�,ܩw"O��##�)d��ᔀG�#|(z�"O�	xׇ��`�
@�B/�,e�x�$"O\b`-��T�H �~I�)s'"O!ڂ<"�p$ 
�;��Xw"O��w�؇
��QK�.S�&�z�&"O(iB��]�\�|u:dG�:x�p�"O��: �԰o��T"C@$[*H��"O�t�Ҭ�������$��6"Ol`p���nKTx�.H�0�""OzP�O �0��[�O:1�iz�"O&!�!�R�x#$l{$M�;��9�"O١AbR,#�\��#f$!"OP���&�K �ݡ�k�fTT(�"OLԹF �R���s	��E�Q��"Ov-��(�Yax�.�<�@��"O`]��>n@ȁ0�B�$��@Q""O���"f]�c&YA&,���bу�*O��`�Q�f���Se��5k_����'�f��ˍ�T��[U�]=g�hѺ�'""�����	�K��	��(�'�6�s���q*�瀗V��*�'>���	ܰ N e�F��~��'�nA�#��T��9�C�%�y��'��MHE�i���Pa�q.�u*�'��"�l+hX�6�[]'���	�'�Ƞ�!!G�v\|1���!S�|�
�'x�ٛ!��9
��źD�D/�(y�' �a)Wl��|�X��t	�D��0�'��4!1L�Mo�<��d��?8�
�'���ɣ�#pv�!3�B8P�({
�'��7#ɑ`�dt�5��2Ϊt�
�'ؠ���^��N�+��\#e�mr
�'EV�a$���Z#"W� �	�'"�m:@oȘd�j�F� 2�F��'	)9���hz�g�&W��<C�'<���3-2��B�W�LGL�(�'�X�чQj����`�tƊ��	�'��E��h�g?XU2C� �nڦ��'�M�ؤ����ʒ�b�<�1�'��}��"ec���Rk��~	 �'�t�Q�f]�T��tr��3{�	��'��s��=1���kw��#�\��'��qi����9�t�g�*M����'f��B&�s�`xC�M�D�$���'�6Lj!��3,���B� 6v�`D�'�� �r���+��4ӓ#��v�N�;LSp�@m� |�ȓHW2iQ ��_BH�&��
.�\M�ȓg����3G��>\��q����HL�5�ȓH��y{#��A���I��$4I
|�ȓ����.\:@�d�ω-��Ɇ�=b�p`�J}`�a�����H��ȓ,��H�n�<��IU4�֬�ȓ'<$\$eŲqh������Jo�a��6��M��"�Iw^D���F �؅�Y�x`�+ʬ	�,a�5盼4:h9��S�? �ĺԭ��Ԅ�G�?1�z���"OI`��
ҴQo��X�D<ۆ"O��i�  �*�� ��e"O�R�o�P���BA��IWp1�"O��I�$�;o"y��\���ܣw"O�  $��q�FXB���2E�*�"O� B�'3�����'g?ܢ�"O>� �l;"��c�Λ3{N,��"O0�Ga��$,��u�T�%��"O��T��\(f���3Y��"O�@�F̈,@(�)�MX�aH�Xʅ"O �f	O�"�6	���Tn��G"OtIEJ�s�F�1h[�[<�g"O���Wc�, ������6J���t"OAk��d����s��~k���"O�}YT���$z���U�U"O�����A%
G-n\l�چ"O���ƪ�����/$6�'"O��@��;�R�q �>�
�;�"O,����*pi��'�p��c�"O�-i��BO��Bu��"���b�"Ov��#�.�K�(�.`��8!�"O� 9�(M�C�$��Q��0u��ɂ�"O(�["��b:nE���6��w"O�ʰHߧarب+DF� ���c"O�=!��[�i7�U ��+@X��"O��s�S:+D�����Y�]@4}ؠ"O� ��펮?�$x�6G�|T�a"O&����	Q-�)c��vb$�	�"Oe����~���Ȣ�K@WFey�"O�L�R�@~��!߸ ^�q"O,�%O���M+�fںl�ȸ�"Or�:���ҽ��F��m�М#��[�o������6My�A�S�ZFbA���U�a���h�N~��o۠{_ف�����!HQH<��ą�i�:��`mD�a]p�!���d�'�Q��&Bu�'E��q�C�ۮ./B��ƞS��ц�t]L���D�:�8P&�W  PX�'�|[P��U�S�Oa��`t!	�\r����Aـx�	��'�TA��+��D��S!-/D��݈K>IQm�-A����C	��y��
�T@��ƞ�P��r��
�X�yŮ�հ�`��/��0'$�YH<���-R�ZiP�ҿD�A҆��E��:�*@��VX�qr0`�8t�I��+Rc����U�@�k�~!Yc��8��	�"O�JW�ݰ6����*U?5����A"ON�ô��<d	�҉��}g���"O���Ύ�I�Npꀈʁ`<Ct"O���E�7��ɠP&=\�%�E"Oz�c�F��]*�:��C�h�����"O� +�U�jG���Q�1�R�6"O�a�A�Ő��<��%�:]b>�(0"O���R�k{���v��{cj�0f"O�\�$�J #�]X2�ʖghف�"O5�'����R����=zܰK$"Ob��\"��;����Pl��B"O�|��
F���"�"Znr��"ON}�`m�<�(��
�Y�0�g"O"4qq+M�A��"SF_.s2Ta�"O��2�&��^)y%�Ńy�@�"OB]�3$߰)�&�3 �Ÿ
)�@��"O4�7�����d	g�)䳶"O�p���4{@pъS��#�����"O���G!�\J�|���G�Vϸ�8w"O� `	�ǆ>P\Cᡂ:(S�0G"O��;v�@�:V�yCt
�hK�M �'���jTn΀9��Y��,LB�
9H
�'�X�cD�0��Ęui	�2+�1�'ϖф��iP��S��,S�X�'(9A��Y
Ҙ��Sd	7�"d;
�'t��`˞5p4r�� �>�K	�'��}�FS4�h�!����#'���'U���g�7Y�B)�l?:���'-v�9�ˌ.<�M��%�v��Xq�'�5R�fY]P���
Q�.��H�'��+�G��Y�X��Ub��J��'�$�[DML<>n����5Lޱ
�'z�EZ�%�<]�e�����%lGQ�<)���U�
i gB�,k2����R�<�$��/*ꖩ�/RsH�'�M�<q !��9�p��7퉯7�(�j���O�<� -X2+P�P �iW��zYJ��E�<��C�_X��� ��8 ���d��I�<�����<��H�IL1�C��<��K�`SH)�b�~7`�
F��<!���  ��T� �ed<��o�<y���?D"��c �t ���R�<��%xVB(d��?U�vX�� OW�<Y��"��}���7T``�Y7��N�<���x�
ು
�1?{�@�$B�<16�V7�"x7fI)b�.Q�W�<i��޵?�H�ˍ-Yz��@��YU�<��P�J��&_|�]h�DCU�<q�k@#D�Fp���m��5EUW�<��ˌ9.e��D�0Ex�ԳW�\k�<�勆����C@͙�~��S�b�<��`۝l�^����^)-{f�����g�<ъ��Ŋ �C+_�L���	\�<�w`��-�Ź��,y}t8�3MMc�<��,�(�"5V��F�f$�#o�q�<�SE�\�6���%	�> ��n�s�<�0+�.�8�4���J�o�n�<�4-A1eޕ/W
 �t���[s�<��ǈO�FL�B�d��1��c�o�<��Iُ-n$X��'��<6�8(�\h�<�b�Ѳm�0�SdF�\��ucD�NO�<i
�?ް	8�&_����!c�J�<1�	Z.~2�C�H�)P����ğ��7�1U���Eoy��)��)�����+#��:�T-%b�C�7����HV=M��2`��|��m���<�`���(��<��w�?�=�����vq��b��&$�]�B�B�01a�B�#[�Λ�Ixڽa� ��s���C#�;��)���]w�~"��9���AUkT
--\p�G!���'�,����0q1Ly3�
֩Y\��ҟ?�;�O�MYt`���U+q��ek��.D���G�۲->,R��S��ܙ�Q�y@�9�"C#v�6}��J���D�DAo�)�B"T��05�P /����#D�l�ď8n���v��rE�՛F��=A���F, �ka��hפ[?jr�m�#�O8�HOF� !d��zMf��G�H&%�:�3�'���;�ӓX���Y�j�$��8����-y��,k�f)_>N�H��J�;
�̊�r8�,á$̡_g ���S�@C(JĈ2�	�A@8b�H�B�4���
G2M"tDA�E��I��E�����y|rY0#��v|!��ϛ��zc�ºs2Y�̎NU��ɀ�P)3�>�S�#��a���T�O���O���5�@-��e�=Q,D��#��[����O�� �a��M�aZ�A�=q�T�ɆFZ���s��$1P�{'�ԛia����ݽJ�#<��!�Tz�d����E�sx�j��Γ��-R��ǱM--�ǧ �H��)��W?�feWfE*xv0�T�ݣ�tф�iP���'� ^H+��Hp(�OD�Ȑs:ɶeH�yކ%�U��6!��!��r>�uI�!�FH
"��<�*8���%D�� �a���&*�<h�I��a�(y��ط�:E��l�5G��H��S�Yp�q㡝�DZv�N�IM������Y��l� �а2a��䉌"ܨE��,)f�c1�6N� �!B[�L�ʢfQ8�vP���Q�.��ŋ$�A��xQ���n&�9�F�m��I�j,��^C	�Yc�	Δ*Z�$�1���#�L�6-���E0$�AA��x�T����XB�*���j�~��)��]h�#	�|�q&_L�r'���i�r�!�i>�G"�l����w �9y;"�9Da'D�l��Ҋb��S�!A8g'ji�B@G�rt<�p�a�S
�+��W�/tx2��2��V&,x�݉y���B�	\�gH Ѻ4D�)�C�I�]���b+�#d�J%��� �e�Z�,�t�aR ׬B\�M@"\���+�Z�'��9jf�>)�D���c�5M餬�ϓ)�B����4Iఄ�L]!c����Q&�\Đ���S�9�h�B�Zb���l+�0>�56 �XP�hқr��Y`d`|�s��MH�>NXTx3�`�6��I�D��ϧW�F��Aˆ]��`qT�O�>�ȓg>I�3b�TИ�83LN�p�`&S�?+�����7��l�$�e:M'?q�DiɼC�,�)�'ɇ~0(h(E,�I�<y��� lB�`P�b�.����K�V	����eiF��˲,q��iN�<�Tc�{�~U����)�Q� �N����˕\���{��'�~�����Q݈�t*z-�ALL�y��! �T�#�(���Ɋ~Ȫ�+���4��a!� ;bH�㞴 C�0&�\�s6͞�G�a pf�0��Of��2 +������ܿ*��\9�'N���n.T4X���	�Ip��D�-�|�ru��)�d��d1]OQ>Ýw
�K��_�|��倗.��؈I��'�p�:�LR�0X�ec�Oߑ^���{FK�3� ��%[���	��h�=�2��$��bH,Q��
s�.K���5�a|b��"T������T0&��bΝ�&x(��-;P4�R@+7��M��	=��Ã2%t��I��bM`�<!�D�=�����2'p�	K|*��f�@�*�ȫ ���ԩ�a�<��/+�Z1���!t���������Ҹ�,:VH�,��)�_$��i� &&�uH$ꔜ|����'�d#3�ڃL9��r�=k2R���'������k���g�ߛZN�A��'2E@�ıL�����e� ��'�����Fւ4-����W�0�k�'1�WV -ܞ����- �Y���=D�0y��.ۤ�U �(l�����=D��!5A�_�1J� ��0-'D�| R�`�h��3kн'|.�`�*!D�`�M;wt�J�Ña���!�(D�h�R��rX\y٢,��l�T"6�'D��d�О�d[��X�>M0�H%D�Li��D�{P��x� ��^��u�6�"D����EۅI|�(0�ktM����"D���$��k���AlS�}+�5s@�%D��!a�V�T�$r�Ӹ\"p@�k!D�d��O�nd����Eu.���=D�t��_�Rd#\.�d1q�8D�xi2���(�mK��R�t���l9D��j ��Yv"В���<�*X�S�6D�$AEӽ}�H7/Ǌ<T�S�4D��b(�i��pK#�ūC2����5D��0T%�IY"�x�k��@otċG2D���j		gtd1��f
0R8p���0D�H{"�Ma@��a@�m~N��d�/D���K�#V��9�U��~_r�)��-D�����Lh�䍍��\T�*D��b4/� w��t%���a�)D�xӃ�E/Z�p��֌[�r�x�B� D��h��]�5�cjWRE�M�a+D��X'F~V4����+3��P�I%D�l1DY7/�j�+�G����z��"D���b�Z/E��¨mg��z"� D��;�Fڱ�����c �=��q�b(D��!G�P3��`��IL�4�)D�� �IF-��
�>��@��o�H�c�"O�pc`K>V���ʱ�F�<Ղua"O�$j'�[�
*"�KC�
xТ�E"O^i0�a_n��$a��0�"OӃK@!�f�`� �8=QP"O� �K��7~x�0R 2=��|��"O���B�͎K�ܼ3�@�;0��U�U"O�����@<2n�
c�4weʙ��"Ove��H�{~ʬ���tS��2c"O�lKF��}�u F���Q��s�"O(�S�jG�\ |"dK?�f�*�"OZ�r��]����D$)4i��"O���"5&�Ja�.فX���p"Ob�� �6v����m@�.k���"O|H#0��\��lp�\�YC*�x�"OB|�2e��^�Ȑ�e*@ ��H�"O��J�9Z�Y�@�@�T�M�p"O�����(W����H1�qH�"O�)��ʍ�"D$]I��N'jY\��"O\鋇�GK?fXJ�⟐5���'"O���D��1|��7&�c:���D"O�(�%-� T�~T	椋G��J�"OT�cS,��@q���bc�{�<eb"O4�i���MB 0Su�ܻA�D�"O�]�c*�=wU�
P$��t�TS�"O�ss��@�AK$D�9�
�B�"O���f�]�v	`�:{��q"O*��s��i^�� R�#�\��"O���q+�Ƣ�3Q�ؤ3�dEʖ"O��Z�!�+�̨���!%|�=��"O)�6�]&_'���P����"O"HъH�\�J�ȁkL/	�JzF"O��;��*C� ��k�4<�
,"O:I�,��`�Zի�߲��u"O�y	��P�p�H娤�ɟ/]�3�"O�M��/J2x�>���-Q�SN�Q"O�D�E�C�2L���-�3 �����"OPtSSÅ�s��Q;4�1Rd��"Oz �dB2w��K��4N��*V"O�qCQ�U2`�)�k�*'����"O.��ׯO�X���2g2/��-r�"O�xsOܛs���"Q匧D�;�"OJ��Q�7C�xA��ӆ����r"Op#"���L�t�"�Ӄ3k|};�"Ol]�"�Ҭx-v��)ޒ5q�*"O��(��N/x��R�K�`��i�"O��S���:4�Y����"5�"؉�"O�aŇ�.2�����dCI7��rc"OD� É�=-\�H�L!T�Xs"O��.�(�Ɔ0O"mZ`ƀ�Tg!�de��	�!n�3��9�E�'�!�˅ -�-ٰ#ն	5��zGF	1h�!�DҹZ}�e��O"rdx�숋4�!�$(k�ZQ�IX����$�(�!���#���ȱ����AS�+�<�!�!}D�̸�lM�1=��z��L�p(!�B�D��b��ǦH>:=�FI͢A!򄋳+8�}x��=M�J	s���2x�!�D�%4vޕ�q/� ��`3'ۥ&�!�D�3Ū����ׂ?��p�_�!�$�(.�0���ߑh�(y�H	�<P!򤛌A���%�̰5�*92�,$!!�T&����fƇ�k�.p��dU;c�!���k���R����p��X����=�!�� ��+EjK�m�p̑5E5*�z��!"O�����5d�ĝ��BK��p9�"O�-��I!��3�/J�E�^�p�"OVh���7>�X���Ԭj�J��V"Ox��/Y�\��h0E�3a�X�d"OJA��ס�zH V$C�x!(�b"Ol%�w�
A�����+Z�V�*"O��A�$B4F�B�HRc�(=o*��"O��R��TO0mS��HO��"Oč �F�'0P�`F-� ["O��ڳ��=�|,)����Xr"O<��u���g����D���g���r�"O�u�B�3Ra��%ͼV��F"O�0�I�!�pԚ�!Y�`�z"O�̨���BV�x;��W�~��"Oұhd#��13�@Tr�d�Ӄ"O�<Ȱ���:�h���+[ئhP�"O�Y�3Xg�"mƵ�b���"O�ApOÖ4��$�����,��"O��
�KUXV4���MK�)Y�ĺ�"Ozً���Z�V���eW:q��ZA"O�$��iT�#/�x�-�Z��Y��"O����G�	`N顇���o��h�2"O��( L� �\��K����W"O���D�+64d����58��"O�<��<����6�>I��@�"O�9��"������A�z�pL�p"O@pr2*jW�h9���u�>ų�"O��3á�--�.��V�1h�.�3R"O@�$�X(����� �N����""O��K�!Rx� f�h����"O$���"�N]��AɈ����"O��Qq�O�^\q�g!�E��\q�"O��R�MS���z���U�4�J"Ol�X��P�;hR��JH�6�h�"O���Z^�24��J@�M�
H�"Op�D�$vJ(�����8B(��E"O`<Gg3;���Pt�^�o=R��$"O�,��*A�.zNp2��̀oA��@"O~���h�(]��`� �9'7bq�B"OZ�0P
5f��yғ���~H�ip"OZ�p
J�(�n����c�T�`T"O�d���J4m�,�	6�;Vʘm�"O�hJՌE�A��]QF`�T�4��3"O`@��,�'4q��#ui�W��"O�l:Є�8��	ɗJh r"O(�@�0G�~	�J�5t#`�@R"O`�!�c�t���j�,��ct"OX\3�bB�?�&���$�#�T�E"OH����b����iE%U�� �w"O��qHRq�v,���h�`�"O�A�G��-�H|jƖ�W� �X"O�yɣ�T�9�)��ݬ�~� �"Oq9s),����u��2��%�F"O^��Q#Oud�:���+|6p�"O�<���/�j���A�iU�D�0"O� Xv�D�yy�=��K*�����"O�y{�b�<t��E��O��#f"O6UKD�<g�lhp%&HSVM2�"O��C�	��X�)TSw]v��"O�U��8���b����3+���e"O�\�Ȃ$��L*6�џgj����"ObSER3 �,X��O�C�<�R"O��1&�(q�H�pb(">xI�"O� ��W)J;|}����A�(�"OP�[�hڗ.�j�0�O ��1d"Ozx�B��1g�KQg��}��q(�"O<`��L�HC���C��iv�dh�"O��J��CFh�d��0�ȘK�"O\�t�Pk�ѲMʆX`n)�V"O؝���ҹ>��h�1��$d&8Qe"OxY8G�S�jHF�"4�$kA�d� "ON�i��h�q��̪D�8X'"OZ,�7�%K��$Z�"ZԨ"O�IQf��2xڀ��&ȬNq�,z�"O�1��ߢ�)Ҧ	�6@��"OJ��K	b�*J�[��"O(��ի28H�� ��y�r��V"O���"�XG�x�*�����r�i�"O�P���K�,�� ��`v|E"�"Ol�W��5���+6��PL���"OM��[�
�lc��I 7Y�a""O����(@�lO��2C�I�,��"O@8�$!m��8�uc\' �8U"O�,r�@��p�D!��n �"O<�p6�:�E�� �*&I����"O���� k���@ͺ,nX\ʣ"OF�q�-��'�t�B��J�6�Ē�"O��賧�';���4y+�"O�ea�[���P@�LԂ<La"O"$��i�>砭e![[�"O���oƈv(��C �4)�vt��"Oz��e�H�]yd �@�T���f"O�0!F�����5���JҞ���"Oji�6�ɭg+\$sckb3��86"Oh iÉӖ7��=�'Ʉ2��)"O
�����Ô8R(N8�Y
�"O챂���� �b�)�`6�4D�X��'ݵv��yt�8��s�,D���N�8 �u۳l�M+(�X�c-D�|���8>��BԀ�~E�q
��(D���� i�
X�b� 03��`�j)D��8��քB�
%�1��C�M��a:D�ȊE(�>3�N�#TF� ���G�-D�Њ�E�jczt�(��L$`+D�8�tG�Ɉ8STY���De�+D��ٱ���k�N8�V"S�|�2D��ɶ��!"�c�-֬1!:cu/'D��閨��1��hŇ�!g��ӡ$D����h�����sKI�RH��k��7D�dSRA
(`\V�*7���G���s0&5D�3���y��\{@W�Ҹ�1D��HteU�"�Pu��)]T�q�C+9D��!)M�p[�aCJ�=��eZ�+D�Pr��x��5@&��2dZ����*D�4����8-�j��+�R�)D��+���x�	¯	+����%D��ipl̴#lN�U��i"D�c�#D��AҊ�&7���X��f$ȹ/5D�@�� ��<����e��qѥ.D��'FQ'0ĀˠHӄ{5� Qf&D��[��Y�(�\AB�J�-
� $D�(���؀~�zg��79M9x�a&D���M��eL$2Ы��D�*�{5%D�L��ˎ���@d�ن��8��!D��R�GA��L-��NV�J��h�iݮp
� `(�;�z���	!OH�!��_�`cr�2f�2`Tx�	0��!�~��ա0����� ���)I|K�.�8�a���!gE<7ɏch�����3� V�r��ѫM�"S��ԼG~"	�2�i�<Fy����~K���5K -��`A�,�v��<a��O.R�÷!ĒW ~H�ibc���}��X��ħu���2.(mr���b��t���$����)��f�0�RQ��:\D�9�cџ=7f�r$ԣ<E��gL+]CP���=L���{CA���Mc�K(�S�OVpY:�������pŚ�4A�X�w���0|�5/�G���vs��)�	@�5}��<%>}�t��*U��@�+?�$�b`=����(O��J�W�5�8���@�BE����_��0��)�' �01A���b���� ��rLnZ�&�Q�"��i��s��8�%n�8K��L�!��:�(OH���ST��(�� �.b϶	��E\��bb�xG�Oz�Y��AZ�O�N���	Ubj58C�@�1UΥ�3�Ի��������ӵ>����ω)<�����FH�r��ON�'�������P���5�"�3p�'a���A��E}���@�C�Z��'�j�b] �
�<y@�O�Ā ��P�a�"�|�B�}�(e���'h(�sD�)q��� `V*v��$�,��)��;-|>�Uмg(f���i�d�^�:��9Gx�O)d�&��dG��d�2a�/3��5o�<AwƽBv� ���D�F>	�U��ZWj����!�*�@t"D�|�g*O�v�\�3��-��b�&-D�D���Ԟh6�%��2o�8 b�� D���"E��l��s�-��d�Wd2D��1��L84_�`)�?
=y��0D�\#��(��K!�I(�Mp�+/D�L��Vx�d�@�F)Q�!��0D��"�>'�@��O��D��@0D�p�P$�f������ ��	*/D�XtdD|8��@�%A�5Kv2D�T���Yhm�P擏N������3D�����Ւ7�� [J�4������/D�@8F�!:��|�a`C�H���+s�(D��A`�w69qJ�)8��3D�x�B�M*X��&�U�hN�8��O6D�XI��3f�� 2�Ӝ����I5D�xrr��-&�
�)bI4\�nћH5D�H��ꏝY����%#1R�$	��%D�PXƋL~&6�Z�!/�ld��#D�����o�8����1A�JL�#M7D��{5�]��!�F]�-�EkE(6D���[+?��Z���{��)*��3D�p@7J�jQ�� 0�ٕFB��(��3D��jS��fG�q��%�]6Ƶsg�;D�(e�
��!��jR��Ě�7D��z4�7L�i���bb��G�8D��uՓ5<���͍�OQ�<��)D�XY5�T�� ���$CM:��2D�\)2��0`�	�ڣk��8�R�<D���Qd��:�A�g�V �!�9D�h1�2 -Q��ʭb�p�ӧ�9D�`�'�6q�P�#"�9CL�v7D�Т�� 0 IY�Q"d \C)D�t[�
�i�vX8���??�SF2D�)@mO�*;d�{2P�n��,��%$D��`��C�'<T�0�O?��E(�?D���7����93q�ΝA�ru"d�>D�p9R	�V��AcR���hu��i=D��ۀj��
����>	^�1<D��z!.�Q��b�q�\���M&D�`KAF&��z�	1�)��Z!��\ﶀ��,��Ԓܲv�ٖ!�U�2�=;4��j�9+t�^9!�� ���44JhxᦍI�>j��C�"OL��2脅��H��M$WT"-��"O��Z��УQM
� ���KQvD��"Oh��
A�{"P�G�.$6�	�"O��pc�d a��7\�"O�A�,9���{�D�)@��y�"O�0&��.-�H0zu��Y� �X�"O�j�yi�EK����R��y�T"O��B�&8� �jbD��Qo����"OZ�k�L�6uM�U���S�Mp�"O�"1Ȓ�z\@�#\>���"O`(b���'i�"��R�	�L;V"O�x���ٛC��|a��|�~���"O�p�K(�,P�4�k�&Ȩ"OBtC�Ά�aV�Ѐ�K!�N� �"OLUV�Z�&�!@�?q��%"O�t(0�A qZp
b��9�VQp"O�h��ғ)H| �Ĩlʘl"O$%��ߊ$U�腮� W�JT�"O��ShC�JE�8�P�T��"OnI��N���y�ƌ�'+hb�B�"O|d��K�P��E��Z�"b"O­z���v��5`�kcH�Y�@"ONmx���:W����נ$Fe�q"O�P3����6��0rqf�-k�� �"Od�a#�ʱ>$�Ca�r�0f�BT�<��@ٍ1x$pⶦ�aC�܋���F�<	�O/����fO�)�x�sr�G�<1""�1F><�r͉*�̠�h�<I3�סU&�Y�&L�K"�d�<����:S����Q$��#
�݀�f�a�<�d��3sA�@�PEM�:�����g�<	�79���Am%T�Pt q)�}�<a��.��ٳ�Ȩ4���1e�M�<�b*Z�	��+!XT�U�f+�J�<Y!  .$���CNךJ���Ed�_�<!���19�@�`�Я8�@!r�͖Z�<)�m��	#�.f�t{dXl�<�i�w"�@���0��`�<�#�v0���q���k���^�<�di@�K�h׊	U����P^�<A���?��m�a/ψr�|�s��^�<�0I��P�\|���Ǉ_SN�x5�HY�<�Ƭї^@�hu���jH8� �)z�<��e\p�!�� :n!`�g�k�<�j�M$R�I��	5d�ض̝h�<�����%~X��B�3tݲ(��c�<qt��,���EBY�e6 �sɘi�<�`aH����r�՟��ᡶ��f�<�_"��P�c��$2ӂ1�Ec�<q�i
+tq�
2��!�Y!d��s�<A%�N�>�������(�^i�Ue�n�<qRH�39 I��V������j�t�<i�G@�D������Mڀ�`rr�<Q��ψ9�n$��ޖw�y0���p�<�D�T);3,\QP���<���{��VT�<W��HI�`����M��ɪ��ZK�<!g�8W�~��3L�H'�	&χP�<��k�9J��P&W�_fB�h1`�L�<٦읙r	l���<TR�ЁN�N�<a�cͺ޲��sg��}+��h���M�<��EE��s`fB�١�L�G�<���ɳz����'J���*�F�<�&:�^52!��D�	��Lz�<� �ɢu�S,gC��[��U�S90"O<���!7l[|;�Q�k5d��"O��l��丠�̽E�!Z"O��8r���^->�����+ZY�P"O��;�k$zH�T��#��rS"O�1�3�������ޱ\��eC�"OV9�A^�^["��E��%��ɣ�"Od�
��<]��	ŃY�X%+R"O"��EU�"q�e׈#����"O 1ѷ�Z�Xs�q!qe�`�PP
�"O���jM��X��d�,B��9�F"O|x3"�z�@E1$�T?�&|�@"O��� j%K@���-�@�1A"O\��B!�+v7�R�Tt�Xz�i%D�P�eO��c�8��7N�3ۘ���6D�$�4 ǌM���Xǃ�"!��ـ�8D�Ha��.�����U8g��ʱM6D��l焱#��x*�bi��;�2D��;��A<~����>kbr�'�=D��%$S��KB���,�V!	&&D�� �MED	�.)C&��N"D��r��	��Q ���ü0���+D��8�i�Qv*a� ��hE�.D�P��F�!�0�a�@3Zq(TH�b1D��Ȗc?	ٲ�oL���S#+D�ҧ [.S�>���aW.fU|���O4D�4x">R`�AI�d�n�����-D���Ɉ1^�`�O�}l��3�?D��1S�ÇI�h�g	��;����?��V��8 �W��@���\
�����0D�x��@C#.�22j�q~��*p�/D�p�.O2^d����-E�X�����M8D���$Ɠ3{b�s��.sT誖 )D��@�\X�y���E�HxE+'D����A^�:���i�1N�3�1D�D1�goΒ0��F�Q������+D�H�T� � �@u���{D�@s�e7��oZ�n:�wJ�W�v8 �E�& �B�I�H�V��ώ�A����b�O�8C�Iy�����$Ęuj򐂒��#3v�C�I4�� ȿ��"��.��C䉻n�и�c���v���5� $>}�C�I7�R9R��Qe|�{��_6+4jC��,���4Ȟ+>cNdy#)�(�~C䉈}ʄ!�ݿ+�z(@������B��r�+��F?MJ,H!�R���B�I�Ox.x���A�@MBTz�hM�VB䉂E����CB3�h��BJ,P��C�	�I(q�g	ӊ^�$銃H��rɺC��
Zm����d�7��d�fF�&��C�IIξh��-�.F���R��`�!�Ti��0�7���%2H��+d!�$�4#�����U
,
����o\�!�Q��Lrȝ���4�t��/�!�$�6#b�9�GQo����6��G!�U��
�R��R��L� ��o3!�ڼ`�F\�"ˮH�ĕ��!�ǩ1"��Tdӑ�<����A(1�!�$�0C�޴ʦ��v?P����N�!�d��x�~EP��Ǧm$�q�$ٶ)�!�ć'�,�[��a�AA�9�F�	"O�x�q�+l�HxQj������"O�h�`OJ1�d��.\��"O|(��o��V��i��ʿd���J3"O� 4 �bכH( aS��ܭ��"Ohy���G�)ƾ����۔8�"OֵP��
}��t���s��Uz""O-��Z�bB��@�(I�8�"Om��K\�G�j1�s�#��A�U"OV8��DCT����),��Q�"O���g�$*�-[�ĉ�&�B��"ON!ʐ���y�n��̈́9x�<X�"O�E�+l<�D g�y`
�A�"Obj�� �#�Xa���<;V`]�p"O����*F�iFR@Y���%=<8�f"O��6��>#6ܳ���&>��Q"O8� A�R�8!�`�f����H"O\��͏,i2���(Q�(غ�"O����Y#��x!��Uh���"O]�Q0���1�_�9�D]��"O>AiS�8�REiC�Ēj��(��"O��
w��
m������(�֠P�"O����.y�iP��ι� ԳC"O�Lk�(3_�ٰf\no����"O�t���ԆU|%�ц[�h����"Oa�0��A+0���\.�P�*�"O&=�t`B:Tp����U����"O�q�\j���`C�hx��R�"O��3Th� ,��$@��B��"O%2(��<�� G[��`�D"O,D��$F^��&�#^(��"�"O�i1   ��      D  �  1   �,  �7  0D  O  �X  eb  �l  cv  �~  ͊  W�  ��  N�  ��  ��  =�  ��  ��  H�  ��  ��  �  S�  ��  ��  �  _�   � G � :! �' �/ k8 �? aF �L �R �T  Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�� |d��"O
`�(�;���8���-0��1%"Oj4��ND^[��"3/9�0|H�"OB���H��*�ʞRy=a"O�味V�!X��!&F�:J�$���"O,��a
���C�Ą�M�"O,$3%o�-���p���+Ն�:1"O��ݢ1����`���y14]2��i�<�6��{_���c�H�`�fX�$Kn�<��A̼VI�xR[�)�Ć�pඤ�ȓA5��('nߡ4�� �)˩%� ���,��r�؊b#`T�eT09���ȓ!�b��g��}�8�F��-? �ȓ
K|m�ș�VṔ���2�%�ȓ"R�X�j�4JN�1�˘X�i����̹	_�jZ��1!g��zܶ��ȓgil,*�J�
j�Ne��i�J%b���f	�(U��:���G��$Y^م�~r�� S�%T"���k\�jx�ȓ|4�1�îJb��@ӵ�ݩn�V��/[`�"�v4�R�!ʎ<��M�ȓ`:��z�ؚh�J�Z��$HY:	��H��p�m�C1��!��B:��0��EnjZA V;9����J[
2���	��4'J�EA�IVW&��~�(aZ��ӹ�>� o�Y�|�ȓ�f�A�
Ο7�H��M�$�����mޠP����/���ANXo*�ȓTv�����{ ��-7�*h��I��sB�8�8���3����ȓNe*M�悡;������X�o��!�ȓ'lj�#F�m�+R&;�|��2)n�C��0S4���T:
b���:�0!��e֊��)��ͷV��,�ȓ0�&�8#���� ع�L�����hO�>���DR�r�*u�c��;ֆ]h�)D�4`��o�z�@$%*]!v�#}��'v�8�⬖�D��U�dG�3a�$�Ey��|� �0"Q��EC@-^⒍Rfh�[�<aG&^�5c�@z%��'C�(����GQ�@F��'�t9[�.�����Cdh�*5�LM
�'Y�rŎ��+"ZḖb^F��
�'ga"�H(8�����3d�dI׭�y�.H�o)H(xt�rG���.B��y�₸1
���.�^��錶��'ў�����85j�h� J%Y���v"O�Is��2�Q��/ڮ%~8�"O�@B�	�6b��6o�/t5�}��"O���h:^WHIz ��-'@=SҒ>��2������)���y7G\�v��ą�I��lZ��~����2�؝�փ��9�~�oU8�y�aP[kj�P'�$�8�Y�f���y�iVR&��â��(�8$)�F��yR*��z�&�&W.��ץ��y�B�E4)�cL���7���y�ϴ:��Pq��	B�b���AG�y��˱c�~l	�P�I7��P6J���y"iM�~9����;� XȖ*��y�� ��	1`��9�l�1#�ޕ�yR�V��~�ٕ��6�Y�B�ӭ�yҍ�,�`��� ��5HR��2�y�\	}*��0�
DCXx擖�0=	*O�S�? ޴9�F\&M˾�넭V����"O��s�B�,R��FOL�Z��)���X��?��{����M=}N�I��ۊv���К�y���L{�� �k�� �.��d��'�yB)�A��R2{��t��dܰ�y�	��Srd��6eޅl^��:�N�y2e��f^=1��e����cj��y���c��3ǩZ=X>��JF��|�Ԣ=E��)R�ᑈ�/$p�� �J�Z�|xG|B�S�>bL,r���-9�>}��CW�w}��$$�|C�f��Ŕ I�-҉M\��bJ8ʓ��'܉' �ժ&�]:d���T���NBf8��'��\1'g�!	��#�g��e�^P�-&?1 P�\G{*��������v��C;BP�B"O�!��=1�z����3$��1E�ieў"~nZ4t4�ջg�	9?�� ��-G�>�d#<����?Q �*��"R-�Ӊt����v��>)��f��w�R��PQcFX� �v��	�6��1�O�Br2�Ѕ��*r�NF{�i�Q?�!�Gf�ɒ�э 1b�Y��-D��� !?�:�)�@�23�����-�O����S�O	�9�#˘Z��apE��!"O�a�A��L:�3p�8TQ{�V����O���اu��	A�F����`Q6 ���P�>�����	���R�&�\�
6A�C����	7O2�M!G�>vK�>i
Ó:�f(��Nm�j���OZ�7���.ʓ�(�	W��X�M�� �0A�~�,������lP�������Ay�0}��ɔ8hA�T�3�7���S�=K!��:�)qT- �}2D��!c�0���=?)�Oq��'W�P�#�&�j���C��0	�'K�x���M�B�����=^���+�O �m�g�'H�OB��)��"L����Ь���'W	�'fvTx�f�9����F��U�!�{��)�i�jђ���oz0���P�)�ў�@�R�O*�-��ő�����qdW����~��'z��e��+����&�=J��98��hO?���=���c��vR�1�h�z�<y� ��CJ1�WIN�oT"�`�Q?q��d�P�'�(Y��`L*����/�Ht���d9�S���$S��qgޱe���HE	������<q�yr��O�r��A��e��,8�ߍ8�ў"|Z�4J2v7�!-J�Ȫ�WM�bM1*ЧC�!�D�y����#�8#�n����ʬF�$(�	�<�A��!��P|X%+%	Az<a&���5�^Ѕ"Oԝ��Q�W%���ȁ-�\!U"O�!0'`�h��e� Ü��b���"O��A剚ri��d�J?�����D#\O�m��c�9�ƀŢw/@���'���'6X����E�T�DLh�C@[\���
�'T��e�6���!!IVR�j����D�	�0|��&�N�S���L�n$��� T��HЎ_r�ܠ6
�53d���b�1D�4��%�d����(�$_�fᄂ0D��DlΙF~��У��p�Cᣬ<�� B�jW,Y]�(0���[h�F��w�h�
�Z}
5Ƞ�c(��ȓs�p�ѣ�YcF��C�#�	��[E�u1q�]8U� �ViS�6��ȓzȨ�HT�@�GMZ	s��u��+��9�OЮp�L(��IET����8؛�p�E�eP" ҷ�ǳu����7O�\��i�j+&u�q	\�#��|!�_�<�?ɋ�)ϔs(��ɓ�$�ᩡ��_�!�� ���I)Y����53~({�^��E{���D�	�D�JD��>#�I"���C�!���Oh�T&@�@��@ڡ����"O����5*U�!!/�>T�u�6�Iԟ0G����NZ, �N5m�L�hvl��yr��:{#��t,
-l����f�I��y�.�	��A�u�^�p��C�?�M#���s�@�8��B>��̲�*��F���'��N�O����d�X T��p@��'���@a
4.���s��*k�\�`�'�X��"+ƈl�q�#��.�k�'"T���)�q�LP��c��X�"�'	�	}���ʢc��f �x��%-�d���g0��hO�өn
������= 	bф��=̪C�I6V<� �E�\��lI��;c��$?�S�O*��wF�9uE�D��n�6�@�j�"O��Vn�����B�]�Lf����g�x��?�O��s�=W498���
,�:�y��K�$:L�'%E�-�ژR"����'a{�߉q��ň%+:"����y`�	P*�t�E	�7���!Ac�h�<�G��?��[3�M=[D�iT#�l}"3�S�OWvh���ǣ(�|<�F�U�T�'ot��%
�7h���G,�8`�!�{28ғ��'m���KSj)YJXx�B��<l�ȇ��?�Dc�/u�1� �9!@lr��O�'�ayrO݁nf�5d��(g���V�y��Ӓ/�$!cɃ������K��y���Ox0u�eяH�Vi��y2���HF�PD��|�������yb�	-M�t��a��Lȡ#��y"ǐ�^��ԇ�#J�����y�h�z�&�x���nL�sG �yb�<�Vqb���0���� �yB&]�v�Z��'C�	4��:qjO2�y�쑣\��qUBz��9ҁ!�2�y�jX�'� D���H=q� �!&���yn7y���C�@@�^���"���y�
�^�����T�Zu�`I���y�lډ�ER�k��[J�5x �Ό�y� ���u�>+�P�gnͪ�yR��6ߔ`��<��jW%��y2c��;��m@��� �z���\�yr��A�fhK��U'1�iA��y�+ȯ�Q��.�c�tC �l�<q%��B����w�� �z����\�<B�'��i��Ϻ2���`��X�<7�R�-D�4cwM[�x���D��X�<i �5T��u!a�Z�[q��붧JT�<�5k!fq��(�#��8� )&�Q�<A�K&	o�0 ���E�`a��&J�<qu�&9�����D��~]�H��o�<	��>@���K�LȨ:�8� �!V�<!1��g5v�	�O�!�6XXb�Q�<�f�/j�t�d�kK�)�4+�M�<Y����l���D�A.u��Əq�<� �97���J''�9k+�|��E�f�<ٴǟ0?jl��1�5i�*5�I}�<	�"��lC�"�0N���i�g�{�<ie.�=\�P�ğ�&�f��G�t�<1�&݅Jr����N�g���{DBU[�<y�e�z^���A�(b���C���Y�<��&̠d�FU��l�
z<�q�sɅ_�<���L�B2�@&��N��e;֡�\�<� ��r��W*j���@	"6���w"OL(��㖜`��-� ��4Ҙ)C�"O� �� SC���Ҏ�h���3g"O�dZ��^�
e�\#$f�90$���y����-"�2� Z�8i�c�� �?����?)��?���?����?����?	��� ?�rS�іn✙��Ѱ�?����?����?�'�?���?1��?#Zǎxf��[�����?����?)���?�'�?���?q���?���B3*�H���CF\�	��#�?���?���?)��?���?!��?ف���E�FH҄�E&|4�4��f�?����?Y��?���?1���?y���?��!bJ(!�/�2q~���ᢁ��?���?Y��?���?���?����?�7�X!z�&���B�7}�4�k�▸�?���?����?����?����?���?�$�(��ؒ�g�//�&�@m���?���?����?!��?���?���?�u�H�g��\���H��x��ο�?����?y��?1���?)���?���?)&F�w���i�1u�z��2`E=�?y��
�4�?A��?����?���?��Y�9�A'��չ�Ɵ�& �����?����?���?A���?A��?i���@%a������G�%	�����?A���?i���?����?���?y��K�\���AG������ ��D����?���?����?9���?᧻iAb�'  �+�Đ�8>J\Zq.��3t9�0"�<!�������4F�:�ːF.z��U� 
T?�M�թ�x~�is�Z��s����4.�ʘ{�fg�x1�Eр=}�����iz��1,X�(
�O�����V�3&�`�N?��a��9NvܛG�
�_I޽Xs�<�I����'W�>�S`�ItH�p�J�1S���Qa#��M5�	h̓��O�&6=��m�Ɔ�"Y���xAB�mRZA�Å֦QXܴ�y�_�b>I��ˌ�hB��*&$v)[��5*�F`�Al�

��	����bm��f�D{�O�򡅁<�8�T�&΀W�H�v��Ay�|BckӢ�
��ƸK�@����b7�[�Λ�l�b�l��O`El���Mc�'U�I��HJR��;)D��C�=zE4�v���eƮX�(��|R5%ǰ[�����*[~�*�kv|�YU]�k�RD�*O���?E��'�|Qq'�� q� ��b��cb�x�'pn6M mX�Ɂ�M���Oi&�1��8+l@Zr�_�*	؈�'N7m�ͦI��b�h����*?�ѯ��8d�izS��\]4�HT%�?@b��Fe�5$L,5ˍ�4����'M���&R�6X��)�5͘T�'�:7���1OJ�)3���~��(rp�X�"������Ȃ��'x7���̓��'���S�.�
�JF�i�4�x֎ӽHk��0��އB��L�'���ZS�h��z%c�t���K~r��1Ͱ�D�ɲb��k���:&�\���''�'P�6M_�=p�X�,��I�3BK�m먊�B�f��?����'Cɧ��'��7���E��3m�Lu[��DA(���U�¦��3��'���I�X�!��-iϼmk؟2�ij�Eq���TA#d	0#.�q�	�����3O��Ĳ<	.O?�YC��'d���6�,G��t	� 3� �Mc.Fg~b�|����<Yu� ?�X��r��=aRi8 ��#�y�Z��۴p��f�'m��Q��D�yr�'��Tz��٭O�S�!�.mTrͫ���-8���:�aH%ў�SUy2�'D� e�ԮF��ە�H�u桋�'��'F�7��(�1O����ؠY�T�`�H+��%l�R���,Z�O��n��M��'�OG�������X�m̒dy<���%�X-<��m��[��hX�O�)Tr�6�Y�
/�$��[I��zP$�g~4��@�6��d�OH���O���)�<����&�m�� ��dU�V�2�KF)M����'!�7M9�	)��D���7�E�7uP#�<R��U�⑑�M�ѱi�u��.�yb�'Y:��4�!C�D-�G]�3"ٯG��0��_�Ee����t��'���'���'(Z���c�:Y��#��3��} ✑�d���4#ob���?y���.��d�Ȧ��4�֍y�P;(�%P�-��XLش��f.*�4������&���� �GN�H��X#I�;1X���2X(�䄁%����DU�R�^�O���|�d�V�Ӵ��&y.�`S O$�~5����?����?�)O�o�P�@�̟l�	�r�Ƶ�U័�̯h�2`��	�]��N
�I��Mt�i���d�>��H�Ð��7��ͱ����<a�<�U C*8H��*O��i��O �$����O�SF��gY�CO�+S�P=�3n�O���ON���OT�}λ~�`��
�L"\����0	!���7f�FA
'���঵�IE�i�E�����t���,��D� �uOz��4rɛFq�����$4/��O� �@���h��P��d��ϰI���M�б�(ʄ>��O ��|*��?���?���..>�BfP"�����D���x3*O&al��T��П��	i�Пp�c��xq� ��7S!| [4KY�������}��4b�����O���	U+�pSՇE�6� �g��*\&a�R��,d9�ɗE��K�)ļ=ܐ�%��'d9���	k��w怖K'���'�R�'s���\� �ٴzGb�3��h����A�q/`����	]����L'�����G}&oӦ4m5�M+,ȹFz Y"�_3	5���=X��<˰���<I��p��m��E|� y(O����� R]ʅ�,y�bI�5I��j���=OB�$�O����O`�$�OP�?iH����<�a���d�ܡ��Ɵ4�	ߟ��4R.|E�'�?�W�i�'8(u{B��_:�1��n�)8���X��|�p��m�ş�r@U�a�h��ʟp�J$B�����_dB~a���K)1%�D��!j��i�'�.6m�<����?���?�1�	O���UiϢ`�8�tA_�?	���$T˦:�o������`�O�2�PdT:�MZ��&jr�O��>Q'�iT7-(�4����:a�`N@�LN���2}�ġ�T�7��x��"�<)���z��2��L,���{"��3 wzy���
�A.�,*�Þ
�?���?1���?�|�,O� l�%.U���O��}�����eЧj�z�*�m-?��i��Oz��'r(7T�[)�M4#��q�JՀ��ˊtb�oZ��M㑌�84 u��?��=��5c���9P��A�`��w�� �=B��d�<���?����?	��?�,�bȁTje%:�3� �D�D��G Ҧ�A)���	؟�$?	�I:�Mϻ�ҵ��&̘������Ô�N�%����oӞ�&�b>���bQv�	�%�ၐ�H9���S �ߘ��IצE�D���3I>�,ON�d�O�i�Ĉ��VjH��A�0Ŕ=����Ov���O$�D�<A��i$]� �'���'�V�8U��?�b=��M�O$Ĉ���J}R�i�(�n�v�Ɇ{z8r�E�?a�A��ϔu���I쟄���\�%o�`G)AVyb�o�Qɒ��u�h�	qj��j�3{�����N p���	�@�Iݟ|��^�Ocb�js�LR:�1�BK[�eT�,��'5�6�MYZl���OF�mM�Ӽ[�GN�%��q�$g	$��)	>�ɲ�M�2�ib��	�^��ȹ�'�f��h�8�(φjM��ST#��6����$�'H8D��P��X�4����O.���O���OZ�Ȕ�F��1�ʓy#D,��.	�	9��3u�f�˛pK��'�����'�~���2p̱)C`M�o%�m�� >�պi�@6-$�4�����O�8��HS�2����VJ�>c$lq�(Qz9@R��O��3��c���b�2���'�Vї'S䌸�F�<+�ll�ǆL~B����'n"�'r"��$W���4k4�A���d\���B-�5(4D��b^����t����J}R kӊmZΟˢ�6qM�A�D�gv`��$�;~_����p�P���L�*|Y�ˉ7r$�I�'�0ם�߹�UG�By��rT.4uz<)[@'q�8�I� �������۟����c��ӌ0�I�E��pd�:�?����?9�i&�;�O9�%u��O,�ؖ-��l����!�z�`�L2�$Ц	`ش�?��˗5V�j�͓�?�u�3,$>�"р#G����V���}f#�1�1j.O@�o�py��'���'��c�)(W����DG�Ŗ�Pb 0	%b�'P剄�Mg-��?����?1)���k�:�𑮑h�`�a�&�u~ҧ�>a7�i��76�4�z��(_6p�S�3w2�Ǆ��N�6�ҟ4%�%;�<����ҥ�3wP�ʓ���G�@�<g� �3��\��/�3�?���?���?�|r)O��o��?Ҿ��w�ѩ_|`{q�^H�dP�
�ɟ��I�MC�B�>1d�iMV�і��.,���1�'v�$��f�D���6'A����8O��$U5cMZTX4���{�˓=L%˵�ӓBH�Q�Ё�,yod����i��	şd����L�����Iz�D����sq&L�;�x �FY� �7-��G!����O���:���O[nz�P�z@�����>.� ا��M���i)�O���(���	��'?O�=�G˳/�iSee�O���u1O�<��C3F.��� �Ĭ<	��?1�C˼ F���(B�}��������?��?a����d�Ʀ!Z�$������ڟ88ь�¬s�g^�r�b���  B��v��	?�M34�iI�O��[�)0_�0K7�.w���s7On�$bӎ�)2Ǒ#}G&�'4�tnJ{������'���"��V���{Ӎ��?B���'4��'�b�'��>]�I)�T���3��a��%�2��Ɍ�Mv�Wr~Bnm�l��]:EB� EGH5xP�U�6�P�6��	�M��iز7F <o�,�:O*�$W���� 0�������Ⱦ>�J%�֪�+n\��2�7��<����?	���?Q���?ᖁ����	�*N&
z�����DJ�� �??���jJ~��0a-���󫋳���%A�c��	��M;��i�&O���$�iE���0��@+ބ]Q�
l��H�*P�|��I(�u�4ۡ�^$�l�'/��5���|!��F6I$����'`��'2��$W��`شe���la��*�߲JO��W�9s���̓t�f�'��'l��g�f"}Ӧ�m/[����Nҝ*������M>� �F�ކ-��������`傀P�t��2I�My��O�n�2s��l�s�R{�Ѐq�N$")���`��ݟ����<��V��3�tx��L�.ؽHS`M�4�f�͓�?��)?��G����ɦi%����@�D���%�D�U�ʄh��ߪ�?�OR�n��M�'c���a�K��<	��C��A�����ibv�Yՠ�>/b�� �?A2y�F������D�O��d�O<���	;��J���e�|[2F��>���OD˓0�v̈́�Lb�'�U>��u��![��yC�[���`�u�7?�W�`(ݴ{����6�?�j�GhPJ �ч[�qs�젰��妥hU��21(�j.O�iG�%04!`�_%8޺E�>Ӳt
�+	�����Z�S�M�z(��!d0A�N�4�˄�=%����n�|��r�^(0F�RAĕ����25*֯w��#?� BW
 ��hƯV�W�b�3�l�Z�܈u&�:d�U���TI8�Ad�΂BS�x#��U.B<З�* �p��C�dAr��> �X A�<��� ��T���o~�f.Y�'��=��B��^�h�1d�w��ҏ�<�Y Ԩ-3��:dզ���d9�H9c��Y�:;Jp�	�2Yv\䘳�D0
��O$�� �d�O&��F3E�
���	U��z�C��۰��95��O��d�O��O6���Ot�DB"W� �Ā���b��R�~��![�C�xmZCy��'��'���'��ZF+<�Mcp��>p���"�ǘI�D(���m}r�'|��'LB�'��ek�S>%�I�}08]���W	4�< ��={�,A��4�?�J>����?9'x?�e'����&�1E�r逡e��tХ)�Ga�Z���O����O����O����O��d����ĉ�������{� kQ)G@�	ϟD�I���+c� �~�2-IN��лW钐Eh�PZ�c
��!��۟0@ ��ȟ$�ISy�O1�i��R�O��H�فH�hP �gӨ��O�ո��]�r�1O���,!��B�%�؅A%hT�eӄ�V�i�5��'��\�L�SGy�\���$�@FO�hK�h�02d�(���M��̃�����<E���'k�z�D�J��L�=N��� &jxӨ��<A�+�3�?�����$�O@���4�L��L��T����\���$��yRʓ�2�����On��	sC|U�e �	"�ċA�N E�hPmZ���!�ē�?a���� ��!2���΋_�����QQ}�'�ט'��'"T�&�G���7E�����A@R�Nq`x�'��'l�|�'m�@�oZ�Q�C�+�8YFn�SvH%q�|B�'L��';�	��R���L� c(S���<bU&֚q$Yn�՟t�I��D&�p�	������>�t��'3��$!P��i��cw}R�'5��'��I*|�(�O����Z}�\����'��h9/J���7��O�ON���O���O�2_���I�/��ap�Ì�x��Aw�.�D�Or�(��D�)�z���OX�)�26���-[�����5n�> $���Iߟt�WlJF�S��b�H:4��k��'� ⅆ��M�(OT-@���O����O���|��C�'��`1���H(K��b�����I� i%�S�QD���ČY��{��Ϋ~�l��?�I����ΟH�Hyb�'>2��#Lf���b�,��9�M�6L|6MʡqR�"|���=3���G	�>� 9:��u�w�i���'���[):����$�O2���GV@2V�ٯV��ȱb��{.b�ġ!WD�ٟ��	ϟ\y���ް���ϑRJ8*X��M��H��!+Op�$�O"��(���,�ِ/D@�܂	H=r�d�dQ��B!/�d���|�I�'gڸ���ͪ\ь	�P����t�2�B��]�������	W�����	�rJ�Z��P0Z 8�kKN�1@:�@�Jj�Iȟ���� �'mN�۟2�Q���X*eCP�)k�)��i���'$2�|��'%�a�:�Ą�G��h�Q�[{�웻I=�	����	ҟH�'HBpqQ_>Y���F/��;�ɋ�
���.ĜW���ٴ�?�I>���?A�����'�:�(#L�0%B�'[L:rL3�4�?Q���䓠 J�'�?����2P�Q.+� d�g*�\
�!�3CQ�g��'���'?��I6�T?}+������Y�1Hچ�eouӐ˓ND�|����?a���?	����Ɛ8be)ɺ&�ʍ��_�0��2�i���'��lf���_�LZ���s�˓>��*�!�r#�V��X�(6��O����OR�)�E}BT����	�#\���͛�p�.����%�M+ I��?��Z~����O�1H� ;A}��rĀ�3B�C�����U�I���I�{���O<�'�?)�
젭Xc]�<o8IPQ��-QU�0�i`��'+�I���9OP���OJ�DI�2�"�%�sɣ&��<1����Ìs�*���]۴Q%��S�`�IbyaG� ����ANU� �~` �M�o�7-�<�����D�O����Ox˓_��h���*
�@�5#��j-�[��C5?�'���';�'��i�A+���J�t�ԀC::B0*�Aj�8�$�<����?���Ć	xj�E�'E*��� �Q'bE�p��j�hh�'�'w�'�i>i�	���������X����&
�LZ�O����O
�D�<A"@R_�O�@]�a�<��Xǈ��4���l�n���O˓�?�)�D��1��C�=�8��@��T%X!(#����M����?9)O�91�^���s�=ӅΉ�����@ǹH��ˁ�'��<���?�L~�Ӻ�E>i�r��u�SE�6]9�M
���'�$��j��p�O8��O���J�"�1t���+�- �W �L�ldyr�'�Ҁ'��>��i`�X�OъX�:�bv�F�2j�L��4,d b'�i�B�'WB�ObO�ʘ)�J}�r�haDH�D�!+ƅl��,��ß���xyRZ>��O��������h���SS۲�x��Pbb����O���̀H�S�Ԓ>Ql��UplM�/�*<�xAǆ�n:�$��4�'��DB&uR����ȳ_�څXp��X��6�'��H�[��r���㟬�b�V�)%$<aq	���-�gO)��� :궡CS��O���?I��� �9��.g��I�pl/%�4m`)O����O���s��OS����V�T�q��#�B�KV���2&&�	ٟ(�' bb�F)�)E%Y�`���P�r��z�EP�����'CB�D�OJ��α6Ҩ����� ��а�ɞw��� �&B�apP�x��'���Ɵ��1L�}�D�'��"�ɹ�(��C���M����v�P㟠�I���WI�5��O
�� T�}�x<��(K7 ^�+�i�R[���I x��Ob��'�\c_�HٕLŊl���ڣlK�>n5;M<���?��'I�VDlT�<�O�ĩ��À�%^Fi���Ұ�ʀZ۴��䚔{��Plڻ����O6���E~�mԖ>�\�jD
���\1�����M����?R���?���D�O��sӾh���ڣ]A�0c�b*�����i6Ш4�kӂ���O>�D�6t%��s�����g�P��0l�Z&FP��dӤ��0�O����OV������g~�
Q:b��7�Y�0L"��÷]�>6�O����O,dE�
G�i>]�	՟dS4hU�K�E�3B�� n�Eσ�M��?9�K��qQ?A�O�r�O�l	��:"[�zD/��1h�[�iQ�0G��I���)0�	�>��<:C(@Q���.]�n�H\��O�u9T�;���8�Iʟ��'���d�;((p����#�~=Ij���0O��$�OV�$�<I��?uBSy(TRb旙<���Żb��x$B�O���?I���?+Oz�Z���|�Ҧ��ww�$�w	�-H*�j�&�P}"�'�r�'���П �	!����O������6$Q��UI�J#�O��D�Op�d�O����!B�nݟ,�i���!���~	��hV��r���¦�������LyZ�M�4�ϧ�򤰟\+�I��V�1`�E�S�5@��`�N���O��D�O,��FN���I՟h���?)��iX�6N���
b V`!�*��M����$�O���!:���D�<���A&��K<TA���VoL�!��|���D�O*��&jW��I۟�I�?��lJ2��A����
|�`��( ���OBA#4"�<�(O��]�+��D;$*ʵC9 Pį�(^�6�Z>!��HmZܟ��I՟��S�?�����|�I�#�4�@m�r���ٗ��:K`�\�ڴH������?I/O��#���O�\�NZrB}!��R7o���pӡ�ݦ���|��3G�$ԡ۴�?����?y���?��P�ڠ3�lї@D�Po�Fk���'��I4�v��|���?��6�(�ZV�Qw������M 90F�Ї�i��&֒; 7m�O�D�O�c�4�O��y�%�
�V�h��R�¡X��0s1O��$�O����Or�døh�Tt{sA�4A�.����0]��2I�����4�?q���?�]?u�'8�������GS�o��� �_Ҍ��'m��'�~m'�'���'l"A�w��6�T�o�����ӌ5��H�C�V��]m��\���<�I����'��E^6���Ǘj���īI%p�|\1�ϏS����?Q���?Y���?��D»=���'�2ȋ�⥘φ x�^p��9M�t6��O���O~��?��&��|����~"���m��Dh%HА K�-˂�M���?��?i֠� e؛�'J"�'I�$c[�f���s! �L��@Po?t �6��O���?A��G�|�/Op1��&�E<i�2��lL�5eR�`���M���?YQ͞�o/�V�'�R�'�t�Od�@ڕc�������p���;����?q�S��?.O~![�=���O�|�`�f��@�2���Y����4,2�Q뗲iER�'���O�D�'0b�'q�����z�,����)L��@�'l�� ���O.���Oy�0�������΃R�b���dX5K��$����{�9mZٟ �	۟��WF@��M#���?1��?��Ӻ{Q�<To��HC�_A�f�����٦�%����Jv���?����� $N��0!���7p�iI���M���_#J�QǶi[��'���'����~�̅1|�fpsN˄4G��[1"�����ݙx��O����O@�d�O��$�OD�K�'��Q���AU�]�(1� ���4s�$oZ՟l��ן��I�����<��ct"��m+"�K�pp��
����uLD�џ(�I���I����!�e��M㷍ٵi�Ԃ3�O�f�Q�,L;P�V�'y��'��'�������~>a��*��m�*�j�<o�¬ˆ˖�M����?����?ђ^?������MS��?��!��df AF��������Tԛ��'��'���ҟP+�j>��'�6u �@3vp��!��]>���2�`��m�r�'�"�'�|����`���d�Ot�D�BPD�bP ��q�F�~<,ld`����{yr�'A���O�bS��s�N�B�	|P	��.7ɢ̘`�i��ɓu~�DS�4�?	��2۴�J�\��݂&�v��ԥ� �9%V�p�7��O��$Fp���O.���O����V�0�@! �BϚL���4rg\�2"�i%2�'��O��D�'��'�#�k��K����PҎ'* ���v�(��W��Oh��<ͧ��'�?�c�F�H��,<�RmR�ǖ�#���'�'�����t�@���O����O^���6P�1�U�­�i
��aT�i7�'�x�⟧���O����?�h��P#s�(Ua��!)�B%Ilt����K$i�Йl��������	>��)����$1�,�Ju"�B�4	���>I���<)/O���O��'�?)E�]1>��B�]�<�"��%�18�(#ֳiC��'�2�'�z�'��D�O��Q3%DL�(���W?�lٙ@�ƌ/V���O|���O���O,�')s(-��i 2@J�aV=sQ*d�E�ݎU���D�d����O����O*���<!��F����'����%�6�X�e�Uw�[$�iAB�'���'�D�D�V�XR�i?"�'H�\*�(L	z�ʩ��D���RR�c�����O>���<I�~$�	ͧ�?9�'p�`i3�E�bH|�P�Ùr�a�4�?y���?1��b$�%��i��'n�OH�\
�̙�qpR={a�� ����'`Ӓ��<��>���'�?���%2���� ���J�*JXQ������b,��i�B�'�\L0�p��d�O����V���O��Z�ϒ8Yx�a��p�ء��t}��'�\QZ@�'���'�B K�OT�'F�H[GG�z�t�P"�MG�ƈlZg��`Y�4�?y���?)�'Pȉ'bBD�|t���'��?b}��g�<� 6͋�l�f�/��.�S���HGfF/.	��`��\7��u4���M���?���@��(���x��'���O"X���X�t�����@;�,��i5�'��l����	�OJ�d�Ob`xF�"]OfT�j��dq���ϦU�ɋs@���}��'�ɧ5�@C��^��A��_��#����L�sRD�į<����?aK~
� I*HU��r�aP s�����愵[�t�Bc�x�'���|�'��dڔ2�d�.�'v��u��&���@�c�'��	ڟ��I埰�'ʹB�Fo>I���J:䡱��`w�Iapb�>i��?9K>a���?�'�Z�<y� Տָq)㎛�>�~D!�T���؟���ß��'��JU�<�5Z����fĄ�5�d+�g>�"8n����$�@�����1"f�\�O�0���y�( '���5��i��'�I�r1�]XJ|����z��^RX��E	$^�,��@r��';��'>�d�'�ɧ��A�l{.i�ਂ�C�1o����]�42OM��M3BZ?q�I�?U��OI�͏���a�B�~��X[��i���'f,5 ��'Oɧ�O5z���
��JqK�=P��۴�@�t�i�r�'���Om(b������*d)�b2���E탻�M����<yN>1����'V���g�<��#��S�
ò��F�fӨ���OX��S�$Ҹ�$������0��z�t��g��YEz�+q�^:f��(m�C�	�=�t�)����?����Ƽ:TD��*�,��ɔ<�r�.�M{���Z:-O�A�OxB�|b�H�v{�sG�� B�hy��i���?%,��<����?����?���[ZzH���ia�q!r�.��YB"�T'���Oj�$�O�Oh��O��{D���Z|p@�*_��P�1��� EƅR����	�����Oy�.)Mb擯%����ug��n�y�
T	 �j6�O��$�O�d;�	% <�*fx�@��R
wZ������'a����'�r�'�r�'=�e̝*����葯��VnvXX@h�?h�8�H��(�M;����?1�QL\(���X�*�b� ��P$E�p#�a�	1o46��O4���<�@[$2�O�O�b`�&�U�Dl�QSs'f�0`���aӦ���DW��3?��]�Fc�`%p�nL�|��ݓE�j���O��*a��O`���O<�D�N�$�OkL4� ��%�ݸ"D�ps��-Eᛖ�'�r�͐�O��>B$�&�H��/ȭ@�L�S&$�;,LlʲWa묄R�J�1svJt��Gé2���w�#_Ϩi���o��`�,͠|ڬ���O�XV�a�[-�y⍏�� d��"	F�26��5�JX�a`�N
�|2 EK!u�b��/��:��H��,~�D��!���p��y���;`
[XǞ$��Ƙ"K�RA9g����� �N�9XA�����m�<{�\D���#U�](_��yv	P���\*��F�-���8`�Lp�H?t+r�'j��'���ȟ4���|
�F�d���y��<t��[��Q�/����G�P����>A�����O��z��`���Q<�A���y�t�ѴF�-��9G�J�����ɷͰ?�!�!� X��.�,D.�uB���q�<)t��6R�� �N�B��i0$i�=��O~���O_}2�'ƒ�q���F��ܓ��Q4r��'}�l�O���'��	L�|����eJ]��^)sT�uӦ�$�0Rb��V
Q�r\B,a`�'{���W�sӊE R���^��6��Lm�H�l�0v"�a��'��p<�-���@��Ry΋/L��ن}%RY�7�͡��'#�{�能W���V�zx�K����x|�����A6�>qh��p��T3O.��x9$�i�"�'��ӅX�p����}��=P��ѲG�]��럎m�$|��۟l�F'֝}�$Y�O��J��m�S��S>�:6�M�u��t�2䕀"��Y#�?}B@D7�9��	�l�ĵ��)6���b!A��)̲�_ ��R���	��M��i����ƚ@
�����ˌ�o��X#��O���$	S������
:��Ĳ�J	@�axBi!ғH�
m2a��$j���q��)]�f`�5�i-��'s����D�.����'[��'���w�"�����)"5&�[�K�3y�n	�b��=i�#���O�����;8�1��'��側ȁV[Ű����kƀ�PR�R�n���`U�O`��%
�����r���T�Q��i��A(l�&8ae�|�gA(�?�}&�ܻ���lBf8�i�Yn�R��(D�(sw��1o�:�q��:J8mȷ�3?��)§Rۺd�Ɛ�,\ �C#P�,�g�9U��}���?���?�������O��S%�ĹQc��E�ȭx�ƓN!����Ɛ̰?Iq�K7���2�K��23TP�"̪B���_1@�B؁�I?�&`��I�G�n\�&��8F��"P�X
m�n�O
����"!��1�� �d@� )>D6�C�)� ��p��=lB��!.I*�
 ���j�-:����i��'*"|��A���x�jՈ��ZE�'
҉V-�"�'d�)�1�U�b�ە(g��#6�'C,P����/>��E)�_�O��Ǔ"�&02�ģD�樐VN͟ ����-qz���b	�8}8��1OT��A�'�6���-�ɓC������+hd�Hۗ��.x� �'����
��[�D�b:8y��KL�B�ɵ�M6ꏈ|���%j@ iنHɰ��<�+O@p�偎z"����O�˧�<�H��H���S2I�A�T�ےE͊Q������?�D�ȠY,h��Ȉw�]R ��;p���h�d,D:йQ@EI5r��Y���߳��I]�@���c��w�d99�eŪxN��~J�E<:g��z�n�F�
���o���-d��-���Y")���jd��G�̥Q�AL�e�!��^9��f'(w�@x(���{�ax��7�[)��!�Ǧ��xb�A��
����i���'��	�-��m���'7�';�w �h���Q��*�:�A���>JU��D	M�q�DBo?]1��OX�"�LYa݊%�VK\)u9X��h�2b�J�`կ�)W�9*T��7�q��O@���7k=8��
L��Ĩ3��N����|2B�.[��hk&n�&.,��9G�0�y�	Z�H��$hY=�=c��V9���M���bq���`�C?*mP�)׃1�A
�@�O��D�OR��ZպK���?Q�OH�t &��A�)k�G�B�HL���G�xrj�Pc��,~�����^
z�`���'��P�I��VL 9��B]�x�F�Ɖ �?	��'D����Խ>b\��6��'����'��p��p<�I&����y��>�I�:�U���������h���v����D�Æ7�"u����0���X��X�I���ܺ_���'�`w�G�8ܙ����-
���O5O����&F�z� �%"lb���_�S:����_�B�p`��p<9bN�؟�����M���_�	���(�d�U�W<:b��(O���4�)")O��BM�<ZY�ɂ�j�~�4��uO��nږ�4Y�S�>bXQ�`�	�,��ٴ���"}^Dl����m���Z��� T��p��D�|���S���'�����-�0=�1O�3?�6�\?H��suc� '�>����{�w*(�s"C=G��Mz��~�O��uh �؜w�(0����$8k:��I�L@$��ORp&��?M)%���1�0x�@�)"������:D�h#�CG�Pz0q�����1`e�8O�xEz��T�a&�Õ�X;6�"hQF!I{�N7M�O��D�OT%0���	2��d�O��D�O�P"+<���tl��)f�ԍw�%��P�A؍6c>�O�Eya  ���Y�o7${�q�чM�ɦBq����|��\(l"D��憱uO�$��n�'F�ʓO�4�������k*=(�	�x���[�XMu��QX�Y�a©/� JwM,,px��'��#=E���W9P��Q�	^�:<,ܸ��-�P�ID�H�C�2�'��'��]�d�	�|z��.����e��T]�����h����F�+G�P�x���V �'~c�hb$F�`<��E(��w�;w?T`����)��	���?!A�Vx�$@"�Y�X �4(�	�S�<�d�V)_},��$Z+�t9q�/{̓r2�Oص�`	�L}��'/���#O�ZI���D��*m�5@��'�ҤXE�'y�)Gc"�������t�	taE�_pٱe� >2訛��$�B�Q��-�,`t�`h	c0$V`�\������8
� q!�ЮT�T��A�knF|2a��?�����dM!o����r�F%�N�{a�߻r�1Od��><O2ա#�:3��84HB�ybO�(nZ�Q��h���.T����f��# 9��nyB쉛��6��O��ľ|����6�?�Cr>�(+D�"����n���?!��Zv�������d�� ju�[G���hP�H�<��ɏh\�#<���J�)`L yd�O4?�ƅ���P|��ʟh��'p�O}�O�8��
�`�Zu�ˣ�JhP�yB�'��y2녊P@�u��N����eE�0<Yw�ɡY���Y1��1PfX遑ؼw��<�ݴ�?����?����]v�ys���?���?ͻVV�B���P~��M���<y��94��mT�'T� ��7�1�0O~��ʘ�~�P�B��&|8�|:7���5Ɍ����7-^�ͺD�ŧASq��O���f~�މ�4��DT R�Ş|�	FT(���|�ˠ\�J�{��̄m�BTRU���yb��2��-ʤbu^�1d/ɠ��ąk���� �	�DjS�&�İ����9`~*l���%e�@e3�i�O����O���ǺC���?�O�J�
^�~ӆ����`IUq��ӄ�x��S4���r�K�b���闒w)�t�
�'��尦K	xDN�j�!Z<x���U)E/�?�V�'����p�M�e|���F	((����'������g#V�1vK�s,����y��3���_�=�ܴ�?���-â� R��H�ڥl�6�D=b��?	���+�?9���d�_�2|9+��C�#���c#�X��d�U�TBs�P�隫��0�'�u7gC��v-k��X��#� � ���o��}�v�\8�L0g �O̼&����녆5��,�ƕ�/{j<Z��?D�X8p�EKR-Z��@+ON����=���ߴ)��d��N�L��D�ʄ3�� �<����7��&�'�B[>��E��ן�j�دV�Բ��W��$�Kv�Q�|�I)Ң�H񨌥]����)�|
��S�b��`c3@L�<�0ţgn^\��I��-3���e�)�S�Hk6��"̵ ����ڱe�h�'@ja���Lʛ�r����;�Ӹn�=s��^sD��6I�,bddc����fx���T�'1y�8��� �*m�b�3O�tFz���� Y��3w��9D��Y�l�aQ�'d��'�����KN����'f"�'�nם-��R�-�IΖ���� 9���0���3B�B���� ����R�g�ɸE^�!'Þl4��5aĞ1��1�RF\�'2\���{|�|�;�3�$S�!մ�����1�.�q0��*e�$��Q0d�Oq��'<�E�	׮����d�&q_��{�'��tY'�F�j�G�4�~��O�)Gz���۰~	p;Ĥ�
:s&O���vAx���O���Ot���?������g[�xX���؄4-*�"6�P��,	�޺Y(�yA0��.U�5��GǒJX4Fy�^�~j�YRX�{�,�z ��+^�Qy��F	s�Ѳ��ު0wh���M~�DEy��K6]l�e-yY2vB��X,�@���a�%6h�V�ƅ��I:ت�aݎ�y�� 7�B��e��$r�,V�)��q�<�����\��o֟��I�
�|���g�*z|�9B��P˖�I�X�q![��	�|�f���&���t'�`�"����
�5Ce�8O]�3�$��]0�
��К2��2/�*��x�� ��?�w�x��F�r��e�55 Igo���y�Ƭn�$��R�W;��*wbL��x2�y����ƪחv�l1�3,L�v��Q���$�w��UlZݟ���k��.t� Ps�y�D���ƹ
��Z2�'Q���sh\0s��3⚰gB�T>��O�� ��%�`��G�2Pą�N�L�#;�r�2��G�D� ;�D���'�Ms"#����N>��F�)���R��)�!�M"�������GZ�B�	�J��)!���/��_����~�'��HzR��n�L��⡋�y�,Iөh�<���O��PN�'��O&���OL�4���gU89Pډ���-3�X�Ԋ.�I�ݐ���S:��v%��}5F�٠LD�6?qOh�1e�'6~<`��G�6�*d�_�d�8 �_���L>���%Oh�׉� 2V\��HS�<a�� BftA��s����L~r4�S�O���Qb���:��q��EG�8��������pd�3�'��'��ݡ�Iǟ,�'T��hB"Ô1�Y{��[(�]4:N�����PX�(P�A�7<��)�`��N�,84���o|y�`���>���P!���0GU=��A+1M�m���Ʌ��?Ƀj]#I��pKD�26K�L�ǘK�<��,9o4X����B�m �Z^̓=�Od(�6�OŦ=���PP&��_�� ���3n��c�h����t��ퟐ�'|�<y�	w�I�v�4���@�c?��{@R�L����D�85A�O@|'F͚>�d��T��3zЩ�W�'l�l��ZΉ'!�ᩇJ�?���c�+�>� )�'0�����F9����snG!�h�	�'�p7�5 "Ԁj�$ْY�\ѫ �'$1O��9�FAӦ���ן��O1�H��'9Lh��el��sW�_�	3|�A0�'8�&Aq�ŀ2�9�T>ɔO��y�H��� D�[����0O�\���c+(��b,�)D�z�]�%:��5�9G�&��`M��f���O�]"a1O��O�X�(Ɉi�<MQ��U�r����P"O*a���.����P��M&H r�'�"=9倾x^ �Ȇ.#&��S�<PQ���'N��'���s���{,b�'&R��y� X�S�Ȁ;x4ZE *ٽjY�M� ��.\��p�'�t�P4�������L@|C� �J}J$�[� Di����#3�I�X��8���|b͝;�x�W/[>P�����%�6[ޓO��ڠ�����1@N�d[W�8��-A !��D��t8Æe2й�� O���'��#=E��N
+I�rP��+9�B���2��}��oO����'8��'8��'���'�r���@�);
��ϟ*h$�r�mK�{g\*!�T���c�.<O��#�` 9�����6b����U--�)���\+�݂#�T�5Ԁq�Q��2Qh���ė�23�)Uꋀp�V����[��\��'��$�D�O���0���O*Q �O
$X��dH @�脪w1O���D��x��AX�Gʠz&X��7iȈQ(~���ƦY�ɬ�M�"�i���W�z���4�?����.h�tʝ�\����$�TQ���?)d����?����.��pf�'N�8AT�ј�)ϮT0�%��������}p�KU�/�J*H��σ�\?0�D�ً�fW r=r�j�C	?zx��0Poͣx	v�#W�'_JV8:L>��0L<	�@�&M:�ZE��py�4���^L�<�B>2���ʑL�z�|y�YG<��i1���r/�'^�`C�?|�<�(�|�m��~�>6M�O���|J��	��?��@6�2aKp���6�C ���?a��B<�C��<6|��i�M1�*��' E$@z��I�X��1M�M�&�O>�r �7z�͢��|����3ge�Q���;a���өsh�|kQ�M�Iq��`��V�I��'��TQ��'�ɧ�O�l�K��&�Z��Q�^�S����'��(��GB)1k��QJ���Ó@푞�$'�m����#L�"A�����=�M���?��.p
F%��?����?i�Ӽ�r��2 >��6L�-I�D����9:�B���E^5\����7^_$	���L>gŕ�w�B�F���$���H�Iv�ed��0\�PR*ñ*�d��t�[w��Z�c'6ɰ�w�Qi�#Z��8a��T&r[e(�䘳T"��L>R� 1=K�0qs���iO(|�aM�g�<�%���t̸�{"ŀ;X�Q��SO~�;��|�K>���-&��)����Y�<Bą��X$LȺ��Ա�?����?	��%��N�O0��w>�I�-�'��t� k��/�]������y22JǞ�T	�3��8�<ɖ�Y��`�Z�䁵$��s�dRͤ�R�n�-T��Q�#]36tY6JZ�� k�&+�v��1eף}���$"�@�I�`K�O���D�&N��A OL5p���h�o !��]�P𧌾Z��yq��#2^1O1n�c�8�jܴ�?���?t( x�"2���,�Dv�I���?���-�?!�����$�:k�a���F>t>8�L��$|��%�8�Iv��(!r��s���\HD�ū����@h Oal�pmS�s�t� ���2����7�6��-Y�"�J�X��l�OVdl�ٟl��z�RA���$q N� ��Щca�Y���|�	ğ�I]�SO�	�VA�9�5BelZRSC�ɫ�Mk�H�!,1�}�'`�4o���p�N �?a.O%8�D�զ�Iܟ �O)&u`t�'���򈐲�*��E�Y[�E��'��J��)PT�T�S,���h�O�V��5^�>��#J[~QtѠ$ƀ���I'�j��B�G(��U��;	���(�3.�Ա�f�޺�C�7~_�)��NUdԱ� �~�$W������b,�q��D��Cp�p��m!�dK3o�hzU�@jΙr�I$�ax�,�$�j`h�$�4Ɔ@���%jߒ¼i���'*r�Z7htx�`�'b��'��we���9Kۚ�9ӌ���������w��]�WKU�ne�c�*d1��O��#��X�+�xĐ��`�h���8E"R��	_R��9�Fɘ0<R���xB4i�R���H%u�0P��eO��O>@�������1|���lR�6�HK׭t],�ȓ$n�p��׿jb�\Jqo��n�l��'*:#=E���]�{�.ˤ�Q4��͠U
ém��qTn�+J���'���'�,����I�|��Bܦ]���4`H*S�*���	WH�~��u�ЈXETl�N"��<�m��^����C]*j�)�W'��9��m�F����<񡇂�#,v9*��7����U�u��Y�	R��� Ղ7;$D�i6d��*@"��� D�t��h�.c{��!�Ɣ;g���j1h=�I���'W�P�df�x��OX�ʓ�ԇ����@�	!ό1���Ol��^�99����O:�H�"�����7�@��p8O���ĢP�z��Pp#�vn0U�'
4�L�h�ٲ��<��͏�0+Ԡ"+��88�4Dq8��p�
�Op&�[���2w-��x�o��_},|���(D��!*��չ��G��$�J��$��j�4F���q����>2&Q�J� ����<�K����v�'q�T>Q�sB��B�ؚJ���ɖ=x��T��,�I4<��I�pa�H�S�tT�� ���c芄$.��jF��ٳ�>�q�ٕU ��<��1�H�Ha*U��H';:�B��u���Nr��+��	V�U�ȉS�� �Z����W�+�!��6}�E G����|�����&2ax�=ғX@F�#��Ѡ_���R��(�b���i��'h�BP��
!���'���'9�w�,I��C�<�0)���](?1�A�D�3	U�y2�
Gjƹ�f��
`�t�P��'Bn���A����/.}j�i���7:l���|�o��?�}&�+�ɀ�)uNd���[��a"N<D� Q�!�8$
V�bɥ/����T�>?��)§m#B-�s�
�x(�8����mfv�о sz����?����?�c��n��Oj�$t�V�� V:	h8i��Փ>q����ٻui�%�r`-�OP*`䍎N��EPDG�J��Ssg�'"޴���ڔra|�&?2�\�V�n���I�]�.���`�aR�-BL�Y��3U0`ٷA��y���7�H	��i �1k��ȝ��'�Rb�<l�=�M��?!�IB����Qm�5�u��'�?A��`���?��O�Z,[���cLU�q'ʜME�!K�Pk&��X8�����?��*1B.)�i�BZV�[7�
2^�x���̦Q�B@=��#JS���@�6o�|Ts�eC�+S!򄀌	�j%�WJ�)���A�o�!�d_�cS�W�ǲ��A�8�1��1�I�~.09�4�?����	�b�������|��4f�Ig���%.͈b�����Of�� �O�b��g~,�o�H0�0�B�������#��I{K�#<�*���)I��y��D�@["S�-�l����;����':�V��'���D�J�+��l�!�7
�2���)Vp�J�k�9aaxb� ғ9�!:��E���8#�+M&�1���il�'TX�,O��*��'�r�'L�w��@�ѳ}Պ��B䖱x;�A@b�^�N_����I%%.�0#@g�(|�e�gA	d�.���p&��p<9T 6[
��s�U�KvHp�ψ�P��'q@p1�S�g���<b�],t�1�և��'�C�I6"���O/?p�����-(��O���"|B� ҃.��b,-.m�@� ș�B�(_���'?�'X������|�*D�v��;'K�G}��;@�'҄6͐�ia2���NB��0=a��ڗ({Μ�"O�&c����B�7\p6�B�c_�, ����0=�R!��bT��F�%��T��$O=�l�I��M3��iQ�Q����I��},��D��'O	+�D��&.D�|Q6����,�)�5$߰(�)'扏��$�<�`����'B����w�^��1L�=��Y��a�C�'�����B�'�	]+�n�"��=Z���N9���
<L,�/�<B|���I�KD8H0��Ҡ����'
��j�!�j�ȸ�'�D�
���sت1�ɐ�ē�"�j����1��%w�~��ȓ r�ݡ���9|W�1��ɥ9-vh����V��>k�v�)�l�4$��b����'��9X,q��d�O��'!�Ph@�P$p�T���t&��J9]�(�i��?�GF�!� �k܆of�|�-�������Y���l��-��>�6
�z��U�Dᆩj�������(D��]���� 
(▁U�T�~�'A<���<���dqӢ�"�S�&�1��hО,������!��b�,��_x�\�3gQ&)d�d!ު	n�	��)O�FzR�� h��w��m�Z�r�-T�3z7��O����O�ђEfE4�x���O,�D�O.��Z�|p�t�D��+k��X�	f;�c��!�-8<O�0)ų_��[3k�-t�eb��$ޡU��y�h�{��E֭M��m lK2��O�} V����� ��a`ԭC�l�(�)uN�_tP�ȓ6/���;�=�Oڥ(]�]�'�N"=E�D�
Tf)�W�$D6�1W A��| �N8x���'Vb�'^d������|2�=�М��º�4��G��1��p�ǂ/|�˳fB
/>�������7*�3@���n���͜�(�I���N"t�]J�-�$m�Bg3�8�LXB�hå�|��.�X��eO���	��i�&R�r80q�W�j����̎w�<���"'8@5�3+��
ƢKq̓LԱO2\X��S��)����c�:a�v0�FC�i�|�YA�����	�_���ߟ�ϧB��P�� Z��mP��W��M���6��p֨�PX0�&WZ8�d��DU�i���`@,�j ����� � ���b���7�P~b0��fú��Of���'�O�A���T�h�(
t��'K݈�B0"O,��c@[�J����(;j���O�m�s��I�Қs�&���h�,U|�c�t2����M���?�*�^��p-�O���׃ =z`AW��� န�'-�OH��E�D "y
#ˆ�G���ԁ]�k��x�OA�>ոa��JD��dܬ^,��'V��2�Σj��P��!��>e�����U���'q�fd�2�מ:8$�J3��>}����OtLR5�'~
7͌�A�IX��a��H�@�Lܶ�J�Kݶ#���<Y����<qRd��\/ P�(ʫur��+F%\[����$�q���qS.�'t���j5�K9!"�l��������Ad�4v�b�I�����X��?k8���pm�k8��f`Kf��\��%p~"h��,������L>a��y�:�D��>(�0��h�:��O��hO�����-�H�gB�tdMX�B�`���P������d�����?�����-ȃ�O��Qg�&"��x�'<2��Eݿ!��M�X,A��]A�O�8Dz�Z>�'�J`�`S*h�(�*��U�;㾡��'��=�bj��8��z4�P�'�4��m�2)fG ����'�:�[�OSr�:��,�,�!�'t����BEd��7(ϡY{��	�'�����2zP+$��Ml���	�'�< ���Hk��=S��	�'K��)a�(r��� ��]�'O ���'��FKVd���aA��!����'���k�^�9x�
1��	�n4a�'UR9Ӂ� 	*�ʩȱM��61�x�'�8]�˓,����g�(�"��'�]YB�qV�6 �.Oߞ�
�'I8�2�A�e�|�v����Y��'<,U�s�$�B�BrH�W��̈́�i"͢�,A�w�`�
$_�F����V�{�*��oE��#o��5�|I�ȓM�.�Ht����H��	�Pb̈�ȓM�da�E�
2jJ0�Ǜ{ �� �Z�2��F=ܐQ�c�[��,�ȓM��m�K�n�0�xL̈́�c����W�P#a������#n��E��z�����fQ$K�T��☟{��,�ȓr/pi8��X/6�M;6oR5
"^Ԇ�aG"uB6�?q��:�L� ��(�ȓSl>�Zp͍v����(�
��Dlq�H�!+���$+(&`f]�ȓ_7"P[��W�p�h�A�N�N�:��z������o��.;�%8���](<�O�H~`��! �,7dJy���\d���<A�����O�ջ�GJ�=@w�G�) ���'��q�@�X�*w:d:čK�*���уg}�u�v�S�s�����O�d�.	����Rp����C�4w�I9I,�m��L:�&�� ��S�t���oZ�L��]J����ul��s� �$'�nB�I�G:$ͱU�T)�N�
4.V?g��$Z����P���a���~�#��u���O'z���L�Pc��H%b�j5��'�j�ZFc�7FLܠ���=Xra�����.<�i1���/^�����-�_�Y��k�6w�Lݠ�����':��q��KR�( �J�Ko p�Ó0(�}ІOQ�:]x��]A�9��@, ?�[�ω5 qj�*��,��� �+J�Qq��e��HQ%��g��H"���:-���0c6?ILAe�JUK�i�i*$������T��V�u���&B�+��i�%5���s�9TbԔ�ȓ�D�'@�_.`�s���)��F�N���
FgU�����p�<�4/Q�|rR�8Oλ?ih�7@�5D`���eݳZ	�p��HT/<�BP����)Un<�����E��$�lDn�P����0h[�'	_ BQ���7�	0)��j���(�Zy��D5i�*���G6�F�J�d�HYP	�T��Bck$|�m�ŉ	p�`ȐA�t6�@�ďȆ[��0A��'Ҕ�ROՃ�XA@Q��J�^-��O�����Z�]@�X�E��4��x��>�O���s�iԣ`��c�ϥo�t��'
,5:'�ؿyX�0 �AL���:��B�3b�����U.��)�I��fh�	q:�� ���4,�y���v�:> ��O���0�Ņ.�����Zq�i	���%D���T�0V�Ɋ�E[ N$, ���R7�ў���>\�B��@�ܙ3��a�$O����&
eΝ�t�+@��ъ�
�PZ%�BAȒ�L��5�.L`P
�E�k����?.�!3��9:�^,c&���3�J�Z�DF>�:�����$F����M�S��%�bMHl��T�'��P�!򄙍f��T��(j @T�W'R�5��j�G^*RУ
�O"�Y��3?a�ɛ8��|�'�ȏ���8APa8�H�i��b�R ��$�p���U��H(u�C�(D3 kʙ1������3��RC0����E�Vq���/)
�C� �$|�,�W.?)��F���[D�<���!M�^�'����v�����I���GC"-�"
*G8y�#�'F�� �?TR��T��-�p{fl^�HR^�A!폨���+�\��ݙ^74q��/(>v��C���0C�C�ɹ�4|@�AA G���pf� ��p�#��'4��̓A��O8�����s;H�q��|"��X	�HA4&�	7�*t`�%�}��HN�q�N�+S��o)����an�X0�%xB;��Ϙ��h�. �]� gP� V�7(�8���	���`�E�U)��6L�}ۢ�R+R�3�e��qz�D!G�Κ�̼*��ē����G��!e�ծk��(���N�d�b�u����`�;{���1�dܦc.P�Z�'�!�f���A�;S��l8���d>�B2�\�p�$�=~Ȁp��#��@�O+�	2�,QY�(ɲ&����"ߧM�D�Cd���-iƤ�`��|��B6,�}n�B�}R
ۀT�҉S�ޯlT��䃂X�ȒFT�"w~�b�J�%���_u$Ks�̝=u�\ɆjSiZ.H�U/Q�t����Wo޵,(6�g�'���d���q0�$�h1ŝ�H�Ɍ�x$+G�	.��`
�z�L<�'+�#F���L��o04�@r��0:28pd����>9��k��⇴}d�`lL�s��b��Q�~I;�OƌAF�c�H�禵λe�69�U P/�> ��	jd*M���%'68"f��&q��=�A�^�b�����$"jl�σY$�� G�&�O��*B#8��mQ)M(���tϜ!�XMpˑ� X�ЀJ

ẅ���$w1�	��ا�I��Q+B@P��Gr��M��c-�6bU(HJ���@f�I�rm���$��2�ɽI�&�q�Fѵ(�.M�Ȑ2`���dB<7���S50�O�=f��_رs��(?��1�c�ɓ!�J���gX���{*�@�a�v�U0�k�9_.v��_67c2(�6C�<��CH��?ɤ��,����i�@t���I;D�(*�g�+��c�(�o�kL��@o@�,��IP��O�9O���VE��� �fI(l ĉ�h.��Oʧ�M�� �#v����'l�,	���S��Q��H�_֮e��(ڲ`�Zl�4�M<.���<���L>&����[(����GH����Cl�#{d`Zʉv�;�daX�K��E;%�@��r�U2������o���*8��k�5�Q*��%�HeaSL1�'}���]0��l"csr�c��=v��Y0��d#�r�ʧ>��q�w��Z�� 7A�&Pxe�68����!ePSDh��yrkA2���ɲDclވ?	�p�΍_�=�<q�ޭ><JЉ�&@����J`̓@LN�z6�зMf wc\���HD��c[]��fPv?��$�\��n@#6����5A���^��Cŉ nS�*rB�:7�՚���zԜ	�2�Q�b��ͣw�NM̓f������O�My����͘�&|���(L�^����Ś�0'���͊,H31i�/>l ¥ꁄ-�I,�`�y�������hΌ_Ĕc���shώ[̄�b	ǟCa
"|겦PR(J�Rb�_�N�T#Ӧەn�
T#���eF��I��:�|�B�]��ywϞ�Kq���#�Z2j��|����oj�z�'������Y��js�J��P��W�P�Kt���d̓�t���
�vG����՛<���<Y��؅ xb �1'\�	tر3����!}I#�<;R��y�	�|�R��ƏC+�6���7@Dᢱ�՘'������.4I�xyLZZ�{�A�L����<94E�h�\����S�T��Q@�1a@n��& �O��[S�8#�K�[���(���`��K��e� ��\ ;h`TH'c)�I2 �t	�g �+�)8��:�'2>}����,�l���hG��IR%��'.18��v�F�_v�ʧ�.��w�( ���A	9z&�A���5���Ŋ?Ԉ��!cK�yң����剭l7DɊ��'L���B�D�D>���<�F�T�����rK��(� |� !@_�c~ڸV�7H͒�Ȳ!Wk�
)r\��!jQ�rK��D�+/����E�#��8,�̰�0�L!4SD0q�G/�&|�%��N��@7M�Q~���d2�	�uOD`ە~:l����݅��%���_�j�^�ȷ�I���%��`�g�*"�ջ���z��IT�$��D��$�Sb�I�&�A��b�hꤦe�Px��+D�E�#|:R+F�����:���U�\9e�ՈUnP�hE�B���=�OE��W>�p@�&Ƅ:r�1 �F�!/^9���p%�l�'HZ�䔱+0>˓v��HB�A28�P\��CG�Lp�1 �y�KW��0&��dd%���%�?��<�`�
&1�e�`ڈy���
��O.�A`�c^�����M��X����D��	˪=_����?ը�g5%�T=p&#��H�&i��B�Z��PQ�@�#'�2���e�O.�3��?� �ɂ�m��7oδ�1@����i�,�t��OɃ�Hң|t>��ٟε��{���4P@�7/,I�\��P�;�?I�	4����I�W'"�,�"�aQ�$|R<!�Z�d|����!�<V�i�D/�Q2�b��	�O	��s2?�r@�c �L%m`�&��
�>I��D2�?q0)�pr�ڐ���?�3'��<涉��(R^��!D��)�HON(��G>�hO�!t��
g��%�GhG#?�< +�� w^�r2�N�9v5�w��6��H���)r�;>�x��G��&(�'�æ1bC˗>/���2vɔ#%p$�q�$6�_������20���7-�+y��Pm��T> XNb��!!>�IV���ɧ �7#*y�0B�89Q��b�A���<�4J�y���yj(Rr%���K��iĶ�e����sd��ᑞ�iS�l%Gݠ	4��s�56v��VA���GyD�I���	�N;ʓ� ��6����ts�B(�6��d&2��E��e�1J�ND����Dl�'��\���$45v�fg͜3�jEA ��9Ξ�I{k��Ӻ��'t�v��s�$Ԉ���	gKۍ��t�#��5qȺ͚GhL�06�ܪ�_7y]��ˌ9�'��	�o�rW��!7ZV��7N�֢��2c~I�ai�	>c$Yϓ2����g�t���E��MB̻chY�4�B�I#b�h�IVy2tyb`I�tM�*������1`h:!�J�7�\@�O�&�G� ړC��X��.�+�.�ۆnF=7n��&
H�6���gFFy$�zy�oV�-hQ>eچfVHH��sF�����F@'6�Dx�̖�A
�b�I~ZP��������-q��Iԥ��B�ө):.��͎y?9J�<��.��%�V@��?��Ѐ�L���Y8:�ː�,.79
����Q��ᛁ�C�Ly,��v끃��8��	Ur\��U$(pN��Z㤎dG\���1��Y=eH���B�+8�e�҇˥29�PpB�e�hS�	��](��<<O
�(Ө�>�[�q�x�ksc�y������!0�T3���v��p����M>|�
�;L����Ff'?2��ь�7*�n�Gy��?Ȉ�pȳՠ/4���%�͇>ߐ�ۢǞ�HO,�kԎ�hf���S�/H�l�gW��3��ch���l	3���v4K��Fx�O����Q��2l�f����?QᆁCW�]�>j(�S'�Ӣ5��t��N��꧎Ru:,Xw�_78��eAS�����?��JX�(�.���+M&�Pw%�z?y���*1!�
�k��Pr!�L�n`�?(�vmVK%bL+���*2��5q" j�n��ƵD}�	Z������8ɸ��ۧp-�4�D��%	wn��Ԇ��[�|ӊ:�&(ظ �~��R��^m6�;פ���B��<�p��F�T�M�O��zC��* )�c��1^#�"<9�c���p��Z�~:APf�PٟXkq�{-���� q���M�>֖��Wb�<|��<$F�#;#�({��ʲS~J��h��-�X��C��=i�j�A���8�ւՊ�ܑ���9T]�A���i%H������uO�ls�Ě$}�� �W����}�AJh�	�G|�|�EZgͬHг��8eh���#�	h0�!�(Պ|�h�s�ŏy���R6�B�������)�'c����m�7H*��@����p���\���U�h"v���Xt��%܁�G�3)�IFZ"6!��" ��@dR��DD��"8��Q>bhء�Z;W��+��:��p�$�3�|�ҴK�6.�:S��a��V.I��@��_6�`�O�H��� pA�t�'?���|b��9A6�ň���8H� ��(`1�)I4Iy��4��{JP��&h6C�E���\ � ���u�-��B�,�������D�;��lz৖#A:��r�Ȑ��It��!�J�!�F�|��>�HQ�=J'S�U*�e��)U�Q ���ͣx"5!�N�?RD�Ol�����*U2��π�I#ҝHa�,��IY��Y)�aZc�*��&�.9J�e��Q���F����萧�H�]>t�8O�O;q���1'��eݞ���R�.�^���"O�h[%&��y���A�O�=?���6O��"9x$��O�"~
����р[U �C��G�N��̇ȓi�4��2�VG5l(�tB��$:a�Oj�R@� s�H���.q�z$a��d��l�����!��]}Ԍ��;ւ�µ��G�!���	!D�ȃ���Y#p̻�*}E!�DOK v}��FڥS�R*w#I�P!�d�b��E� AV�����@;+!�Dփ'�$Zv�%��Z�(S6 !�dP�>"�|�%��c��񀩟9G!��\�^��5*U��'��D���*e�!��L�t��p��Sb�LX�b,є&�!�Dƹ�|Mk��I�JBQ^0Vy�)�ȓ`Uz�10�A�`1�,z5j,�bх�[b(���N�F&xɂ���J.jŅȓ_!ܤ�@j�R��q�E�Bx�H��c�h-�Vo��XT0v3d6���S�? l�Y"w��ѣ�Z08|��"OhA#s��|�>iBe��Y��@:�"OB�#(�'R�:|�C$��1��4�T"OMV��-j}����ژ{T"O"�cË4'����!c��yՒT��"O\Mɖ��'[,0��,AY���!"O�Y�d��-4��䱳,�>7~|��"Op��GɟP�px��9a:La5"O0H�tʇ}�Q�g�?6�EA"OZHZ��(h�@�J@.v�)2"O�}q�ȕ�pֶ3��"8*j�"O8-�W-�@Wl�14P#o6�K3"OV� ��:`&�izt�ۘk�4z�"Od9"B//Z�!�W�O���"O�L��l!欹R�D�"��"OX̊����p��
Nk`���"OJ�9O^	��x�n��6rX�&"O�`��(3WH���ͅ?X�t;"O�CQ�E�F�"A���@�oR�H2"OFm醯���i�"˓�虋�"O�Ub�Ŕa��X�K�u�m8%"O0��];��f�4F,��iF"O�x���)�r)1A��esp�7"O4U��>x3������h��+�"O�����>�Ѓe�YRpeY�"O���2�K1$F.�8*��Ը�"O�}����/42���O6����"O��)�EX�	o*�p�&I�v)�"O�-�㯁B�~��Z.!��1"O�XP��D���Y�A҆z����"O�`���y��8�4'L:��Q�7"O��x�JL��8WG�5nLm��yrDQ`9��ֿ>� {d_:�yREX~,��ca��)ֲТ�c܂�y��$���b#癨ln�e�䉹�y"M�Z��q��˞^$uy��K��y��b��1�tWFt=s�/_�y�E��Jc�.L%��mu�Э/��B��<4p5´-��
�j51Wț�$��C��-L��zvK�.�4��,Ykf�C�I5t��уE�҉�$��C$#9	�C�I�J��15��/u8u����A��B�I<�z�kPd�|�N�s��GN�C�	"N�V�Af��=-<�:� ʙ9��B�ɂ�p9hu�� ?�\Q���Ɂ}m�B�I�t�(	r0�V�kW��w�H�}NtB�ɪ_�-��%��L�)VXB�~�Vh@����`�9Q�LB��\��0�$�4�"��� ݼ"tDB��3�TH�s�"B����!��\E|B�	�u�����������;v�
B�	�S�������䬻�"P"SB�	�q�1��Í^cx��,�+��C�	���MZD �Bf��"'�u�B�I,c�!�D��
�1k���p�PB�	*�0��Cdݮp"$��p��w��IJ����H��jƖ�P����=��]x%"O8�Q���$6u�\z�mF�(�2L0�"On$K��n˔��LY�)U��"�S�I��RB:� s��7�je���C�!�	HAp����	�t�� a�-�1-ɚE{���'��!#Ոkf4�;R݀�P
�'z��
VH�^1�XSC"#j�`
�'и�q1�Q�{������P�	ۓvt�0AJ�� �Aw�B8~@��df��4�	�"O�)H�舗x��|sw��T��D�0"O�H�g�X� ��H0��t
�Ӣ"O�\�������JJpS�s5"O~5R�虠. Ѐ��@"9=r<��"O��p�Y$
o��vcc��d�G"OP�7�*Ru�Dx5a��w�P���"O��R)	�}�F�aℤjH\t��"OZ����7�*�Jcg�B�tP#"O��Aa�)Os،�Ѧ�Lh4I$"Oԩ(TH�$��y���)P
�z2"O��ˇ��6ʹ��L� 
"Ot����9*�5��iJ g`���"O
43���3�b�X������p�"O8���+i�p(� �R����"Oh�rV��$�Ѣ�����$��"O���w��1>>D�R��HzQ�*�"O�ʐJ�n�`	bu�6eI�,:�U�h��ɔ>��dk�C _�F4QFJ�>@W�B�"*8���
R��:���� _�B䉓,�
Y�o�+\�H�%h�b+L㞘G{J~b���"D<YsA݈g7T�2#g�<a�&8㞅	!�V�HJx42"�Vb�<�� ^�����8P� VDb�<���Z|@��ˋ%����WE�<qAB ��zu"�d�	;����֎�D�<�R�/�����S�"|v0H�M^J�<	E {�|Hcd�P��iJ��[��hO�ON��˗��9T�T��JN��-p	�'}����kY6(A90uE���:���'"�pC�T��iӴ�>T�@l+	�'�1�4	[�,��4���߫;�) 	�'w��B��D�T���7J�ҭ	���\ (A��TT�hx��C��a�ȓZDu��I�/D)��C���p5���ȓq�K}���G�O�`��'fazr��DH�ɔG�`�#vAۧL5��p�9D��f&ŷja�����'8͖Mjs�1D�\K�
ǎ'��N�0s-���'f.D�h�QL,Z�>u���M�I\p�jT-?Q��:�'(f�%I��TZ��Fƕ�,����O<�o�s��`��a������ON���' �'đ�[G�K#���a�D8=�C�*.4���,@�d�bi��|���ˁa�<�'C�.�*A��H�k��:� �^�'L��'U�O}�J��ˉ\�����*h��'a��]�Э �J(
��`��!��O�#�u� %Quq3�Ë�X?�U���N@�<��
��~��ު^��"NVyr�)�'q=$�1�MH�ynh�R� %d�V5�ȓ\Sp�F�٢'��T�r=$���Ɂ'��D2V�-�L)�HRK�R���$��l?����x�u��OD!Xe0M�Gd�~y"S���<E�$�>wm�qD�5J��!L��y"J��-�L�Pvh��~Q���7C��y2)��p��U��Эgi��Mˎ��sӜ���ȳz`�k�0@?D�A�"O.I@�Z/%&����j��l.�˧"Ol�s��	My M�U(^ q�^��#"O�/$���@Ɗ]�l�w�P����'���'���gh_!!��@�bǞ�@tX\��'I��#+.�a�a�S
�\�����y�/�#i��Qy�D	n��Y��Z��>AK�,`��ד
��=IqΚ�b�nQ3��o:� V�����-�F���L��O��0�3"O�=�6*�
j�ag�����!6"O��;�lH������ ;p�<4Z��!�}�����Γ�b��A�릸��	g~R�tL�r�*<!Ǥ���,�+�y��$T�jD��B����w�ϣ�hO����փA�� Z�'�!����G=�!���~Z�+ԇ��:̘}�"$�@�!��i���)u
�R[�X�a��P�!��ڇJW���B	�P/@%����Z�!�T�h�Eb�">)D��V�ˑ!���%�N��J�:,�u &� +}!��[�4��A�B t�0�k�eA!��	}8jq��9t��,�' �4�!�d�(�>a�5�z �/��j�!�;8�D��va�
R8�qsn+|}!��6O�
E����4�j��]�e�!�!:�|5x�F�1v�,�5O�`�!�$ށ_
�*�)�"М��g	�!�D=v��
w&�����Q��]�!���/-'0�s ��G`���$1 �!�]�,�n0{�a�vl�TۇaD�!�!��ɓX��)�7�η/�
J&�)ϑ�G�do�8�����h�Z�xi�2k���yB��?;�0����J�S�AB���y��!������Lp6 rD^��yB �&,��(��E?���$͂��HON��T�'xf��LZF�Ny���)E��]x�'<ܕ��+N X��9C��>�*Db۴�MS��)ڧ(�&�(��DL��1f� ��M{�f	������<0��FH�<��&���^��Ȉ�%��e���C����V��Uz��x����" �7|���{"��� QMB��t`A�Sc ��ȓ*�P���ͳ0k��r���'hZ�ȓ90 �Ȑ�� 8^9��X4j������?ѧ�V 3na!{�2i��
����'�΍�ʂ7�<՘��=��p�
�'�vT��
@�'�0��3�ǀ,*h���'a�E�u�3V�p�k�4T	i�'�,���!��q+f���$��'!N�@�'�Ȱ��&e����O��m���'z�R���8r�[��M6e�FH�}��'}���+AN�2m�P�O_׌���'�������"iw�U���/T�Ԇʓ%��X���U�zA��@��(�ȓ-l���M�z������E�ȓ+�8�B����|��f�0[��L�ȓ-,v�#ˉ�7FL�;��	�hs �ȓj�*j	0����!	�!� �ȓ)+~|����a�ر�Q�N�T|����vP����3� �
�N�8��ȓ6�<j��ŠN|(
@IR&� ��璉�K"�����؅ee�ȓi�y� T�6,h�y�G�e�`d��2'~�2�,ްF����i�#��^[�<�.��h@e-�"/��ez��N�<��J�s�"�p[�oN�	��I�<�"��>m=�L�,��1xF�F�<nT�%�F8�ɮ����4���<��D4r��ɀBIH��-(u��v�<aaKΕ"�Ɛ�3�fIErc�|�<!ѩ�RK��8�-��p��\!W/|�<i��$P�(�Y�+��H�
�;� �c�<� N��C�H
���e D�5�J@�r"O���T�G�8�����Oűl�>D 0"O�T��O;m���*���$W,�pP�"O�t!@�d��S�hO�J���"O ��I��I�01d*�p����"Oi'EY�`�T� �(�O��z"O���0��(a�lӧ5�$��"O�`��8?�FxQA)L?'�
a7"O*�;����JD� �����"O���V�8*줘��ą�Sd=��"O�̫�球h�FD
Ra��X陷"O��h�l�B�l����X3h$�y�"O��rc�:H��oѴ>�`}��"OpD@��1�<�î_�Q�8��"O�eI��a��Ųo�^h�IK�"O�(+�aJ-C� ��ډUH��z"Ob�zWGW�2�4	�.C�,��1��"O��:��CRT�¥�R���jb"O�� 7OZ{6n���jաR}���"OfX�iQ��Q#
TmC�d�D"O"x�1�N�0�H��p-2��A"OH���N͟$��%*7��,o-`��"O�|4N�� ��)�/!"�×"O�(�Ř$mp�Ua�e�]3"O*�j��^�Ng"(9��.\��	��"O�����/�bdÆ5}UH�iq"O�Y؃�P�sJ�;3C�;X�@�"O�H�&�L�:�H�Bi6����"O�=����D)�� #k/��	1"OF}pd/�i��8+��:xzd��"O����>�đZ���&o��H"O���9JUY3扡nh��X�"O����
^%�<y�䆱g��
�"O�8[���(��#\$If<x5"OL�)��T7"dhT�2k�FZ���"O�}8�.(nI���SL�
dB�L""O��3 �V�t,I^r.y�am߄�y�/G�j�i��7*��l(эR�y�f#kBtp�C�L�� I���yb�C*&!���әO`Hcw����y"��7����k�I���X����yb���c;�q�@��T�x䠃�D�y"!:}~�ث�FY�L�dh���@�y�%K.F�ȘۂD�H�VZ�b��yBn��4:d��<�,T�����y��C/�����6���땥ך�y�䁫 '���U#�;6a A���C��y���8/<8�9��R 1�&%3�Ւ�y�gE�Ț��#̗:  ��𤒬�y"��b8��y�g�"5G"�h� ��y��G0cV�J�ƜC�nɈ0A�yr�	��I�J+S����N�y��>1rP+&�үta�%ʗĘ�yr��dQ|�⫘%Z�VYʆ��yB�'Q3t���z] (JE��y2��=j��#�Z�Fc>��$@�!�yRHe;'"P錜?{J��AN8�y�L�D�Y�F@�9;��`D���y�� �%{h�����;B�|)DC��y2�T5+pٓ%%�2b����ˬ�yr	���-
B��4*���#I�#�yb�c�r�y��M��<�����y�O��v�2a�䠁����#��ճ�y��U%Z�Z�Ó
}j���+9�y
� �@����x$��\<6��\#u"Ob�J�� ��y��Ӳr[估v"O~@��ϩ'X�]ᣮ�</HZM��"O�8��m�|t���eWl��"O:A�C]	S��]�U���ڪ��"O��U��?M(H�r�v|�B"OjY�kP�@��f��^���3�"O��C�1<.����o�.7�x0Ƀ"O���a�#0�D���""t�*�"O6us ��U���гM҉��"O6��F���e�PP��:bʔ;"O`ZP%+dfȡ�7
�>s� ��g"O@irFJ�,\ڨ��h�=��,;�"Oʙ�ⅰeP�gA�x���2"Oy
���L�9Q(�@�B���"OR��b��T~�@Ȁ �Wy�y�"O<Q�!�ɓ ̤� ����t�]Y�"O�@�2G�P����GlD�07"O�]�e�	Q5��@�/�!]e&�˂"OԩEk��m�P���㝌W��zR"O��aE��8<l ��`ϚT5"���"O~X��+Z�F���P�%��d4�"O�q�
שXSf�bE��r!��6"O�Ek�����3c_�C��%(C"O�T�B+���x0��<+6e{�"O��ch^����.چ &�0��"O��s�]�e�Th���<@�"O��qR,����qH�n��`*�"O&,2�+ʾ=�Z��tN�'�0�Y"Ob���.Nc��DAE@�"��x�"O�1XpÂ� ~M2�Ԩ��""O�ԙUk�C�ǯ�D�\e p"O�����y����.\�{�X� q"O -ag���Q� F��O����"O��K �T�Qr��`�K�U⤐I@"O�ɱRT x �0�d��<�L�K�"OV,�F�U�Q�Z�3�,_.���s"O�+)N�#c�-A�,��H�1�"O��bU�:��U�0y�Xa�"O8���Ow0)s�d�v��r�"O�A��&
e������1�N\�c"O:�x�/)�FoN>��c*Ob� 	�qZ�XP��7����'쒗�Hm;�8ibb͹R"Oj)sb�B&`��h@e�"U���kq"O @��,�"��S���x���S"O�� ҃�6I!�X�"DQ�ymT�R�"O��dL�v�d`�� PT��"O0SEjѧV�fd0���O� ��"O8��mS�R߸* ] W�>��"Oz<b���1o�bPC�	�O�V"v"Or,�B��v~v0���J$r|H��"O\�1 Z�"�.MU��CzZU+�"O��R'�.%�y��K�^^x��"O<y�3oJ\����"AvP�"O��0�cl\!�%�C*q��c"Ol�Q�cڹ}X]R��S�elfL�"O\�Zr/UUD�ȱ�!S/i`�QJ"O����+k�le��ʔ�A참�"O��*��r�T|��Ɛ.Κu��"O�q�ίdp�2�w�f���"O����S5lj��9Q ��Gf����"O
�9u
*|�0h�$�~r�c"O� Tn�=c_��T
A�+>ȹj�"O� �,��Oф{\�| c�\C0�qZ�"O�
P�җY���p�Ì�;)B̈�"O�䩖
 �<�y��#y��"O�%����K��3cC�X(�:�"O����aζE�X�p����9+ "O�1�L6�t��1A�;wZx��`"O0q�RJ� ��	0sO�uDd�kP"Oh�if��,Uib�2�?�mP�"O���HG	A�ȡ[��W�Xx؊"O&$��7m��#F�,g�vAY"O��8h Sl�xk�BA$6Įc"O��ѠI.�bԚ%!��
��e{�"OR-��֛ B:Ȑd�M�,P۱"O�LYJ�3$z�rG�ުB�
$�a"O�H���HOvN�8��
9H��÷"Ol��M9k4^-�n�Ԝ��f"OHQ�A�ʼf�"���Y�"��"ODd'�O0/���$�|�M�E"O����A�9p��S/_�_��K�"Ot�����o�d�Ӂ��/~8tA0"O
����qPTE�0��(`��4"O`Kcd !�*I�@nS"R���"O�PAkЩuVlH��]�_�v�H�"Oh@��K@��1��,@�a�B)��"OʐB]S����j�% ���`"O�9�m@a �)
4�	�MǎA`6"O.գP^� j�����f"OV%H'�@�E�0�C��ΦT�&�1"OU�s��JЉB��\/�f���"O��22�6A�:��T�bk�	B�"O����˟"�F�Yd�Z��l0k�"OX��B��+qֹ�T��� z�1�"Oz��pė%1��1�V��B�"O�y�C)�'Qƙ��LZ:C��a�e"O\�n�-}22�0F��n�;�"O�i�&�k[0q�KG�4$�'�d�e�
i���B%Jۨ]����'jNI�cW�(�0ŊCU�UN���'@�� �S���2U�Klh��'��S4�ոR��@#o�=0�Ls
�'
l�A���/��kGm[!6�q��'�x2�e��%���E�P��a��'/`#2�D�+�d<Ѕ���Z�I �'!�A�AR ���o����I�'��K�<q�e� ��*�'��Qpq�P�v�,a��P�l����')>�Hģ�J
���Y�fT�h�'�P�j�
^��p|��I^�W0�r�'������pĄ���UԐ�i�'�"U����\c���.��ct,���'��ڀ�	�h���/�����䓫?i��L�� &�ڏ~��1�h�IT�m��7D��B2�X*A�1��� (B|:5l(D����aJ�v/\�<�d���UM�<1�	U�����(26�(���NK�<i�q�NIQ��9*���oO�<	Q��,�� ��8G�2�"ON�<�Q���U��{E!�.d!�%��\�'axr�C,�Ja��/�|Ћ(���y'�n��A!�"��=��%��yjˬ=��x�%N-�(�����y�C�O��s&��xP���8�y��-�8�{ �ܺ�J��E'�y�Ȱ'J`2����=ɐ�K��y
� �a�s K��F	0�؋6	,�O@`�t�,���X���;Ҳ`��l�Oj���O�����$G@�i!�AF^�9�b�ڡ|j!���;��yr6��g[��2wf�$}f!�źC�RDR�,��WL\,�����;�!�[E�T]��Kצl��qG�]��!�d�<	��I�A>-��!3W�A<�!�d58Т��G(b{��ᆇ_�
+��'.�[P�2� ����b�+��'�!�d�%^1ҘA�a/oH�v%�l9!�D^!qɎ�C�#zK�-���E�;2!򄝝����G%K�wF��{�n�8!��	7&P�B�܅T2ZV ގL�!���;
��
S%¿4&p�D�O�!��z�d�Z��J�)�V�2#EÔ��B�'�F�􈀟1��pT����L
g�'�O.�}��2k���N�}]�ykFm_=zxȓ�D��9f���zƃж>��-��8���2g-
 N�N�rdӳe�5�ȓm� 1 F�(����a
�cc�5��g�-�7��Z���SEJ�L��ȓK�P�{�iI�M�����!p}��lV�ࢅ)�VEkr"C&~%�h�I`�����?W`��y�d=]bE�o��V�B�	�v��Y�ƫ8�6�J�E�4zR�B�	�r	�4(dB>d\*''�  �B�I�;��$�pC�'�̡�	�T�B��	4�bAUhR\�yag	H�Z�B�	a$\t�A�	�U��Qq��V�B�I}t����'w<��q �>Wu�B�I&k��a���.m�h���B��B����ʯ7"2�Q�L�1VHC�)pn��
֋A!���0�F�"C�	7�u�'%��"�H��t�P��.C�Ʉ�xݨ�@ i>A�SGC���-Yज�}}�fХ)�BC�I'˦�?X��
uED�	~�L1q"O8]XA��h�LD;ƃ��qkTE�U"OT5�goSF$�$EW��i�s"O*u��|�L����;}�����"Oz툵(��"q�)'	M����"O�F�p��IJ!n��t�ƨ�a"O�(p��9u�h@��5�F��"O*�R%�б5ȠP��d@"*���q�"O^����ʰ��f��U���"OZ��!��/���!�u����"O"	�QG֜%�n5�V���KoR$��"O�p3"!��t��0�  8����"O���b�Z�4�Va!�*,,:���"O������1��ѡ�	��@��d���D"ړ��$R�j�P�����+y�UQө��0u!�$6(��L���3��+��/�!����{fKN?�^`���P��!�[;Cz��8��K�v��%c�*!�ĝ42�����@ �~�ʖI�!�d\)C/B��V
�:z>�RAJ�8�!��W��ˆaڌF����1��`��'/ў�>ըT�3v��D��o̱���N1�y�$��
�����)�3#�ڍ�1N��yD�-^���+�/��!��H�[�y���J�(r����f��@Ɋ��y2#�"sZt� D�Jr�`aS��y�m̷M
`s�/M�I���PC��"�y�B��g<(�k�'�M�H�Z1
K?��'�ў�π ������;���1��1}�6"O�YScΔU�^��C
�'����"O��� �D�e��qP�B�4�hi
"O�Dhr �R&G��dzS햝�yB��!#$��^3�\8l�T�y2i^!|3�]��h\;����4��*�y��!+���A��Ic�9"D���y2�լF$�v��n�p�[bG��y���%e~�f̎yd��!���y27��x�`�y��cċ7�y��{:T����u7)S����y�+�@F�x��УrH�*�+���y�L	<
 ����S|B�{��;�y�	����z�KA(rf\XQ���<�y�g��^kzb�O��[N�r��](�y�g%F�x�B���K�|� ��ȶ�yҩE��D�ȱ%4���BK��y��M�s� �+q�*o��)��P�yr���To��3����s��jM�y"�'p�2x��Xės�J���|��Q�%��>��R���zΊ��ȓa'z�h����qh�
�A�^�l��Io��h��$��4��-����7*mXB ��LE!�D@�
�pQP�ȌL����[!�1q2�E��mO��a�tK:<I!��Z�Z 
 �E�]TJD��H�9�!���>�u�v#�,>�SfI0\n!�@�E���b�M܊�ô΁�vZ!��Ű$Tbm��K[����@�O�j�ўp�ቋCy�w�ҤF>1P��O�&B�Ɋr�ڸk3�����3�aK��C�	2`"DE��뗾xf�U�1�Y�e�B�ɬ���CEU�zx��E��8�C�I���lɂ�I�|	a����cHB� ����	�(|�μ�"��<��C�I|+�)H 蜋J����
�C�	�7��:g�U=Hip�zQ�Ne �B�I���xH��E��K�c��B�	� ���BE�s�����H�l̀B��r�zAZTmȴe�p$��!T(o�C䉉U�� �(H�e�Zx(�����B�I����s��\+>�2A)p �C��/@��򥋱d
$�bO��jQ�B䉋v-�ܛ�/L�T^��+2eضn<~B�	/��1l-b�S�	�0\B�I�g
He�Wd�����s
�*��C�ɾ|���[q��>�|����JJfB��+����-�1nbf�*���U``B�ɚc�"�krc�[xNL@g/W��4B䉈�:�� �8��D+�\�C�ɀSA�a+a��^�\����Ng��B�����eRC�d�z���5��B��6\�b��&�Q�J$���׭P�|B�>x�Mi��W�֑#4�һ=fB�I)q�а���]�Q���*�V��LB�I�?0$MS  C(��U��n	�2\B䉃}5��[��JV4��	��LLC�	(j��b�^�f����b�5�C�I8X��\�Y&�-��ߴ@�B�	�~ܖ���gЩ$2P(��I�D�fB�ɳE���
0,	���z�ϒ,� C䉐'��E*WjIh����#�8$`�B�ɖx�b�i���hR!i�&*�C�ɲt��kΊ&3\��8�AˎG�HB�)� �UڇÈ:y�LD�ѫ�$C�x%"O�f"51�`�ߖc)�ɹ"Obd;d1 􈁏�-3
pA��"OLM+pޘb��
�Ā�a� <�g"O��E��s9�i��⑵���b"O`m�e�E]p��t��e��A5"Oda��T�nV�����#-< {�"O�DPSD�.ԼQ��c$0R�"Of$hH��m P�óg@.�$Y�"OPd9ƇX�^�*m��˅	���p"Ob� ԥ�+3�>}�e�4H��"O��eCBarl����[�U�.$A"O��ã��D�)
F�l���"On��B�C�p�ʗ*F+T���y�"O�U���1D����=KǨ}��"O&4���ӪS
�	��]����"O��ZĊ*{8Ĕ����5]���t"O��yu�-]�hH�5B%tJ&�!"Oh�i�r���X��\�E82,� "O`"Cn
�tˠD��et$��c"Oj5h˹KTh���	Ցr�0���"O`t*�`�<���N���	�"O^�i��S�o��Ӎӎ\�6� "O�KU�5|}Ԕ�u�H6Gd�E�A"OB<k��*�M3��_1,��v"OR�E�T��,@3 �i��i�"O6�jw����"��2(�ޜ��W"O��B���e*����m�$a!�"On4)e�*m�tAԭޘ[Ī|��"Ob�┬2)�$���1\�i�"O�Y!
�9��E]�:�H�"O^�@rㄞZnf!��&�7���"O2�j���9C��ZXHu�Ư�p�!�_e����CG#eh�0(��hA!�>���Ն�G�u#�'Џ>�� (IlX9r��	hgR�г�7�y��D2�d��e��1gH�C	�yl�7 �d�	h>�Jp�$���yrϫe�`X1�ېc��L"�cS��yr/��5���+,%��`7I��y��=.��s��lp-��雾�yr�Qj\�QJS�Ӑ��;�k���y����p=B Ct!�	z�#�j��y��L���	k"Dݮnb�Y9dJ?�yb�W�+.� 	�Ju� �s��y��S3+g�y
�� np %{Rlޢ�y�F��-��hüC��pq�۠�y���lJi�1銨G�P���y┶B�	q�ł��H[!#Y,�y�i^g��q�	҂Y|Z�� ���y"j�$��<�`��A�q٠� *�ybƁ+5T��+D�;�D�뇆��yr ͝c6x}��.L�I�Ă��y".��<��MQS�4
Ea2�H�y
W.{��҂�y�6��T�D0�y�MV��Ҹ�0)�uKv���Ȭ�y"��H>�� �8p .���V/�yR��:��I� �ڡU���:��F��yR��>N$lɲF�/!_����-؏�yr��3]� ��v.�>�b�kuH��yң\0��d�0��r�K5�U�<�G���ܕb� �x������Ec�<�#�4)�V�Q�ϳWd�(f]�<��h�@(�� ӭL4�ɀ�mYm�<� �)��ꏧ���B&A�-e$��H�"Od�+��*�����3s:����"O&����\�}�Z�Jr�'j��)r"OP�i��3t4̑à�>ؖ�A�"O���mE9_�ٺ@� �j�u"O�*�"Q;}=��PփH($���e"O@�a�i�� #��`bǷ{z(+"O�@�!W�t�P�[Ţܨd���P"O4�7�[<@��$��L�o�T���"O�� ��F�*��	&�ͩse��˂"O�d�/���r�P�%l|!�"O���2�:*��J]����"O$͋��H�q�N�`Th��"O�d���#D� cfH CSN`! "O�C��<|����j�[_ ���"O�K'6‡�Ϗ�ٙ�"O��c�䁉[@y�,pG$�1�"O�1��F�m���9f�/Ҙق�"O��`�C�0�"�˖�:�B�0�"O �����iܢ� J��Bİ4��"O��/N'dTP%A�)ĭ/�T=�"O�QRW��L@\T��M�Zx�1@�"ON�q����Ss�D&�x�hlK�"O�!@g�M�i�nyȆe��N�f�k"O����K�@���ɅD�:�؁�e"O|���l�&V$ݱe��@m��"O�-ykD��02��4#�ɑ"O����	�6m~R:`�T�r}0�2"OL!��������EA�����"Op8���_1�d�X$މi9��C�"O��&ˉX����t%�7|p�+v"Onq�5.X46jЃ#ȧ-�VA�"O�I`+�AUL9�F)�6m�\ ��"O�yh$`�Uh�g��&j|be2"Ot��}8= �ړJ��bS"O�DIUI���0�����
� ""O���3���#0�5� ��?5���"O�M�e��5���f�E���U"O�ڇ�4a��؀5�RB<�S�"O�� �U8H��m�$���y$�i`"Ot�B�4H%�A*��R4@�8Ez�"O��A�T2L0���T"O:e���F�J{䔉`$�I�"�"O��S4�-
��8[R#S��V��a"O��*��M��|z��V# ,�`(�"O���G�M7bg�ȑ$ �r2r,�e"O��ӧƓ��8#��Ѿ0��"O`Kad��<�|�i��!`J�i�)&D�SB����Y �G�Ըɤ�6D�HhW���q2Ř��� -E�<XS�1D��q��<ن`�0D "U@\`;�"D�<[E�n�VUH�+��,|�c$!D�|)Vk�B;z�#��ϖ0�j��K?D� +�k�������F�6����;D��s*V�&Y(����Q��4(;�-D�|�,P#F	���e�O�"f\�rt�6D��(1G�1g��y�*O	(.5¦$'D�dÀ U�5X������hP�a$D��҇$H�q�ؐ�V'�2�0�B�(=D�����4A����nP ��u8T� D�H��"M>F���ҐiɴL���ⶩ0D��0�E�;�1�iF=U1�T e,D�0 �	8판� `qq�l��! D�PKCL,R|Zx򰇟?��d�s&2D�� �Tȴ.
2��UŎ�;sO���"O\����1u��f-ɸ~E��9�"O �a�����Sw,8A�0K�"O�th%SS\�*��S^�P�"O���K�!���2��,p���"O
{���2Jj�:C�׿V�F��q"O��1��C|xQ��$Q8��"O<9���ǭW���P7h	 Pr�"O�SԣL�G0m7�39�h���"O~�f�	a���&@�ܓ�"Oz��WR�`X��
��C�6X8
%"O���/L�,�h�!�c��@h�"O"��V:R*.=��V�*ꊤ�e"O̸��F�*����cA��4��"O<x�Ůs��ȥM��7@�ɰW"O�p�_p����A�2&Ƙ��"O2�su��@�)��֫>��1Q"O�Q Cꔷ/�\�ۋ1��$`�"O:���ɖ a �)C��1l��@"O�S�jӧfN��Wd�#N,��""O�ಠ��m���rÈ� sΐCt"OX<h�dV4{>p7��_� �Yf�"D�aF נO�~��KE��u8��!D�4)p��i��]���K��i��?D����G�{#�}c*�%cJvM��?D���Ri'~�±I�9W�Ȱ�=D�tx����[�F����=:78؈'�:D��h�#0NՖ�FZ*���ul7D�\r�#H%�D�q�̮+�ȁC�4D���ㆾIv����L�)#F�2D����JF�^$Đ�7�.P��]!D
5D�p���I	T�<��/�B��!�0D�<���!~@�3�^�4�Hł2D�l2�� @Z�����h�0�/D�XQrl��؀@F*֚�vh*D���D&��u@��%��'�)D�А�����	�K�~d�XBSO&D�t၅�&D�jQhG�ݎ f"D��I(��+[�U`b/F�Fv�h�'�=D�$��f��F�0]u䃼#���Ig<D�a�OG���0���P��|!�M8D�0��� �I��	�c��y�L���7D�\a�Ƚ=����l�;
=+0E D�L)v�āM��A���\�"D�$��bW�8�Q�ժɂO��u��H D�|�W�7V���D�0
��I��!1D��x�̄+"�4����>���N"D�<�ϔ�'P��̍1_��h��>D���dލd&��t��X����,<D������6&+�t���E(|�l���L7D�d+d�3+����4��͈B"0D�0��
I���Ł޺^��2�,D����	Ko�PT�>ts�Hkp�?D���UNۄ-���,(C�<Y��;D���tc��0>���7�ƈ��9�.D�L�T��w�L��i�`Gx�9�-D�0�֤�f����cB�� �!f*D�|�mB�*
�ˁd=E�u���%D�̙��*NϜD#G��%,12�(�#D�� �-K�"ly�M\.l7&T�%-,D�l�1!��Z������Z%7��m�i-D���WJ������Bڂu@b�z�� D��� �]�̶UrE)�g/4�A�:D����B. -R��E���b$�PYb`8D�� ��A%L�.YU�E9�π2�d�q"O���%7:��h���ʸL[a"O�0�$?&��{f<Q���Z�"O�!�n�+�`QW�Y�u�����"O� ʤIW6L���𰃗�<�(���"O�qQc�l�d:���4WJHC�"O�`���Z+kp
�ۧa5N�T3�"O���G��goґ��@O"i�葐�"O
��0c�Z��� W
&`ȡ҇"O�|H��SxԄY$�6
�t3�"O �ѢE�|��m��t<j i�"O�-�Ā�"!@u���H	$JEr6"O�h��g�/IR��(wE�97�� "O��y�)^����D��@�(hU"Ob�{!kܜ�.�J�h�2Wu�m��"O�bROD2̈́ w%"6Z
M�"OzdP�P?��X��&�uT�a�"O<�q��t�Q1Ѕ�VQ���"O�����"�@K��X
O��J�"O� 7�C3Q{�b�PB�kw"O$`3Dȧs�ٺ �O�>H,@0"O�!�Ħ���>��p��Q3N ��"O���d��"o$Zp���ћK�x5"ON�q ��	���K���\ ���"O�A�DoP;shl�A����bF"O����V�g�p͙#��'7ܖ��"O�9���(=2�5`w �̎� "Oh@A�ȁ8|%��r���F�i��"O8�K�"��JA�0�f.2��d�#"O\2�,)�eQD�ۭ0^�,@7D�X97��p� ��C9���w(4D�X���Tm�L�U��#��<)��3D���L�?nTm��$�谧�0D� h�`G2-�(�� �'Ǧp��+D���O&��)�g�4B������*D��S�Imk �wg�8�����f6D�̊/��I�����S�r��`�75D���5�ńN��A�J��1i�e q�3D�T:�Û8�\� ��?�	ˆD3D� �3�Ӭ����l[�oֵ��b0D���I�x���� 
�Y&�5ؓ%/D��q�E�>�ڵ#+�w#�U�	/D�4j���!n�K�#��&�΅��?D��X��U��+�� .�0��n!D� �O�`{�D��ީl���b�a?D�,0&A��s2 m��.�7w�qjf�*D�`s�g\�g�`�Z���8h�e��#&D����U'.hQ�L�x�@��!D�P*R��1���X��Ё{3� �A*D�434��}�H�3�ۢ!�
5hS�+D���7���,|�tAeiZ;<J%���(D�T�4�J=Q �q�WK4` �`�&D�X��r�j�s�χ�Lծ7�ZM�<����l��@�ӌ�1��Y���^�<���]M(�8��JRѬ�꣦W�<�$#�.�Q��a�.l����XV�<���� =�|���p��婇�g�<���C;?~Hzd�� X�혶/D�T`�jԩ^��9Qȇ�y��!�:D�pi��@�9)� �� D�X��m
�8D���c��L_�8�A�­WZ�5��!D�(3��Q&ǧ@�ql<h�a� D��0��X�ec�T���3f�>D�d�Ʃ̢
����� �gq�YC�6D�� j�Hg��`�����sA�};B"OD��%"B���q˰���1)0�!�"O؜�ƋUC�|ݢ�c�s~并"O��P�A�;���v�?o[A�"O}Y��	!�:PgBR3.P0�b"O�`j'�])>�c�@�	Q9~�""O�Ձ�Έ�n>Vа7�Q�5+4̰"O��W��rv@�-{y�b4"O�R,�&`����h� ^Ty�r"O��
�~�"r�M`����"OTA0C#�s��)�ET�v�p�"OV� ˜)A�$�҃R;�@=��"OV��ŭ�V�zAX�̞�2���0�"O��f�;Y�^���DD�����"O4-a§MfA4��&�R~��
�'�f�K��¶s�I���*����	�'��hS�d�V�{��p�'��9��Өsiz0c�<Dv~!�'�8� �ܽ^�h⇅0?���'$�\x�o[#4��+����; j%�
�'��[T���k�D��`
ͩ*�`���'�0`���"qrp�2�*	�X�!�
�'q��t��3w�Q�w_���'[���_�=�J�	�V2i��$X�'��q�f�PH ,A� 
`�VU��'[���Q�%-�r�t�ԃg���)�'�]l��I�����+[��X�'�E��o݉Ql��i$Ï"*-�y��'$8y��l��y�,z#K���H�:	�'����ĭ	�5}��Ys!�7|%��C�'��9aШ�*;L�Q�m�t�
qs
�']�4�G�^�lX�LrS ��:=��'����L�=I�X�q�֮]|Ԝ8	�'�0�E����s�bFQ��m�':8
Dj��[$�%Z�-T�S��Y��'�Na���� �J��B�MpЁ��'��� �'��`�d��A̋;��(�'"0);���"O%�}Y��Q�D۠,"�'Q*+�S![
���;,����'Vl�V��D|��$ݸjV~h1�'����G�L�" �N,,�I�'�TPBt�!u2�y��Z�]��'Gv��Ui�<��2��
:G����'�h-��M�4�ҹK �;^�P�'~L9 ea��L����+l�e�'���C�4LL��X�F%1���'��19f��tw�	jAh��"N�d��'~Π:�C�7׾q��&�j����
�'�$`�v4Ъ�fyЅ�
�'\�8��+��u�`��`D�\�>�0
�'We�G/D�B��wLx�	�'Y�����ĉj<`�p
�yG^T#	�'F�����RL����`聰i(�'��}�&�(h����zlz�'xʁQ$��S%�q�g�V�'�lH��'�j��!�N`���(�E�22F���'R�N�>	�0#�J�v����'(��@Bͷ7��PI�q�ll;�'�T�z�,^:N����0\}l���'��P#q ��F	�չT$ؐO�����'���I�'��H��Y`��9�%A�'���4�I�Q�4�f+O2H��	�'��4��,B�HƩ�Ģ��*O>�@�'1�xs3�Ba��!��-�v����� ���E�3�����@H�B�#�"O��Qi��^M��pB��"���"Of�����b�P�2��Hl�I�"O�(
4�D�J��WF��rx���c"O��B�,M8Snj��$���rlq1"O@x�%�=5��"�b*��%��"O�QD�1Z�\l�֠�j��"O�Yt뙠=���KGe�7.c�8��"O��#d�A�c>��CMiM��j "Ol�h��
x����oL$DV�c�"O���1��4��u�� N*�S@"OQ��n.]��H�.�/.U��"O�=@��3L�t��P���&p�f"O�, ��؇J4$0%�6F�ƈB�"O����`Ї|�Qsc��N�b�:�"Ò�d�V�!@(�HB	�0LoB�2u"OAc��1���2�R=_�i�Q"O���'��%|̤�w�.Xܠ�f"Or)�nȴd�`�%̍O�C'"O�8!�G�
���N�z9P���"OX|&� ?�4�Rっs�z`"O֔�D���\�H��� F�L���"O���ۅtt.�	�����q"O�я�Oqh8�qAޞ ��bS"O
��P� �5�r�7*́l٦d�"Or�����G�FD��)ͧ}����T"O8"�C���⤉��C��4�P"OR9h��#2o��
���H��Qh�"OF�P���_��r�Gާ;�n�b�"OXUJG�3=@��I�Ӂ(��1"O���rB���
C@�'ג (S"OF S㗒O���["�YϾ�#�"O�Y���P;��	]����+ZU!�d�\& 8��̸�R�z����eI!�B4B�^cҐ8l 1{��6v�!��Z.Z?*���<6Rf]�֍��!��M�ܥ�ԋR�:��A�`����'� 9�@�5&@�0S'��:�V�c�'��IX�����Jtk��u��]�
�'a��-7'Q��
��t��j�'$�m�L��
r�j�GK�W{��"�'`�j�	08D�c����T�	�'�Ԁ*�4-�@��̒ r����'�z{��ܥG�1ա�U6:���'�Va���O"*xPa�w'VI"�b�'��æ�=u�P�6)��8?`t��'��A��.w�z&� *g�@��'���1L��[蘸��ѻ)��LR�' z���IG�gʖ|(E��UTXh�'ݪ�!`�ӛ_̀��4H���X�
�'@Pv�� �lل��7}�m��'����1��N8��E
�a=,E��'0��o�*^����a�����'��ɩg��Ѣ���[��i�'���"!��+Vt������1�V��	�'�-`�ʋ� �	��A�L�8�'X�
v�T�U[��#R� ��2�'�VL���(���".Fv.R(��'32�+�dG�&*�a��<?ʬ�'U����aC
���_�4 �m1
�'֖-��f��L���&�˟c��	�'	�� PK߇l����)s �11�'�ؐ��aˀh+��N�m���0�'M<D�ԣ�d��cl^�ze\�H��� ��mN�m�c�f�7d�x1"O.�c� g�b�'��2�"O��10���p�	0Տo��$� "O���!� $散d��bS�P�S"O&d� oV�K�:)�Q�4`5��"OD��OtF�5!���:}��"`"O�mhvLߜv �G���8(U"ODDcn�;���(t��1C�N �U"O2�kJ���a��)�ѸDV"O��C�ґ%��)�D/ܖ.��Y��"O���dN�T��A#W��
BZ�QE"O�9Yc�ߝ��#���&K��i�"O6�J�M�*w��%˓ǚ�f�c"O`Y��ȸ5ENTk��M�E�X�0`"OZ�Y(�y9J�1�]3���"O\� @�^�a��4��dOK�����"O\�B1�V�ud�	l@#Xܝ3��2D�����2w�F�qq���QߦmR�E2D���$�;R3BD��$F"=F��3�5D�4���!gj��&��FC:X�#5D��ǔ�7V|��m��'�(��'D���*�	�|����H�k�X�e1D���j�d�G�ˈIp��q,D���$K�v�� �EE�(\�Q��7D�,����6U�s"a�/P�6|�sB7D�0���/5+0���+�" ��+D�Ȫ�n��h9���i>^@��'D���V����`�ڳ�A�c%'D�0�G�A4Q ��z��ֱ*�P�x��%D��@Cm�>Smx5��G��6J�Q�?D��`�0Z���O�4h�=���;D�`���k��J���2kR���V�'D�`�T�T+dv>|X��N5F���%D���S��R��������|���.D�(0@n�HB�� ����uL+D�����٭;"��:��F���4*)D�,	0"��t��TK��d9V��c�'D�(s1T ʴ��Vj_�#��0r�#D��S�
X�	���{���([9�����?D��Sa-H��pɖo]�~����7D��F�A�w��	���2Y�-	C9D����$�(������2b�3��,D��@�,]=��E�b�$��C,D�$�5�N!-/���ڦY^�����$D� �ʔ.s�D�q���	�����B&D�����`Ҵ(�T(D� 1��E>D�h�3�ܖ8�68r%>w��"�B/D�$��x�&x`��A4,�����%(D�Ģu��Q�آp"�dB ���$D�����t+���t�<����'D��
C鋟NX1+�"�`���eC$D�$@�T*I4�s�Ղq�iC�"D�H	r���w3`��@�E8���*i-D�l�b*��K1`��2������W(D�<B� /e�e����[ۆ�C�1D���lRl��9��&`��0D�$�HV��Ma�j�=hG1D�|�5C�4��� �ĘQrVD"W�,D����U�}�rP�� <�H�)�` D�i&M��~��QaH�0B`��f#D��W�B1Z`p�%a�=@qZ��$<D�tjF䆖#z�%�DI��#�b�*Gc9D�4�Fܔl^쐁tD7pBL��"D���G"ĹeR��X@�ցb��!�?D�� Dh����beJ�� a�9w�x9�"O�,��֙	�2�� �@ڒ��2"O�Jv�͡J9�8�!r��"Ofc�mӾ*Q
�¬�>B�	:v"Or83��-��Xy��V����q"O��pDI�,�^հ�C�\�0<Ҵ"O� z���t��w�/	x8�Z�"O���Ia�<�֎Χ1ohZ "O��9 ��

e�+��8��I��"OJM�2B�w�HudŜU�\Y�"O�X�+X�(�"]jX�r"O�aV�)x��2��\@v8�5"O �B�(]�q���a�]�=|��"O�Xb��(�C ��k,�y�"O���͔��� �Q$���3"OX��p��i�n�$���_Dhd"OlX�DʛD�K^�vBN��2gπ�yb�!]�V�jѪ֊i�`]����y�N�r�De�2Ce�1c����yB�X0��0��oX$n_� �D���yr��2�12�1^B<����G��y�N��T��%��j�xb 
º�y��?l�6y��gF�u+�i�I���y��n&XR�\#j�F�ɇFO2�y�DB6S�0�`���;\�R�
i���y�@O�;Ll}���K�S��{0G0�y�j/x;�̛���a T�4�]�y�
��p���y�e[��X�Ӆ��y���>Z�( ��W�΍��h�yR��W�\qRfɎO�@qB"��0�y"�ޣ3��K�I&Y,�2bė��yRm�Hݫ��ΗC%T��A&Q��y©L�6��	A��>Jrara���yE�(���E��<_�������y�	��,�x͘� 3@��S�Ă)�yr�7ؤ<N��#s��w���y��J�k���b!�"H�����yC\��H����R�H �+J��yBe\2B������O�<�ح)�;�y�Aիj�|�;�)�"b6�Q����yᗶ��%X0���j@�3AO��y������N\��D��&~!��m���+��̓'�@pC��!��,b�*�r�Z�0ߔ�PM��$!��[�R�����+E{��k�K��M�!�J�aQ�k�_b1�#kJq�!�dݏ=�pX����ZO�� d��!�䉌Ah�5�%F�+o?��6��2t�!��'5�2M�҇Ѣ�Ժ�!ɖ�!�D��R�(�f
�|�4 24C�(�!�$lϞ,� �@8u �/ز�!��/qʙp�c�#O,X#�D��@�!���	)�iӄ��^^����Ƹq�!�W�`%�1�Tcνc����cM�Th!�	l�����Jٵ�ұ6m
`Q!��>J�q�d�uj����,�	�!��3c\�Q���#�:���KC�!�/zǼ����fUF���	t!�D,r�j�!�3lŹ޶Oc!��D�9�P�°NV0� :fO��.Q!��i�����X��0b�I�=8!�Dڜw�8I�E�#x.uDb�#q�!��ޥmGD�1�NQQ X���R�!���{�, �6N��3d)cġ�>f�!�� ح��.� >F�a4�
�h�$"OL��GH�v���0wM]
O��e�5"Oʵ���ʫ8�4��v,P�u��}�2"O�Y�a���Ɇ�@�y��0��"Ohmq�� (�x�b�U	%���6"OYc'#ɛ[�|qr�%��q��"O�, RC�:0[�	��/p*q�"Oyp�Ã9]`��hY�G�Mk�"O���c
oV����i�CZhW"OTkb_U��1K��	ޘ�0��}���7�i>9p����X`�u�S�;5��
3�O �/�¨B�L�6�uJ��ɡJ5�H��#�����V�)�6�v�E�MC�F{b�O���ɖ ^��Č��H	(T��O���F#b����^;q
��h@�Twh!�ɩ���KT�5)T�Ys�P�V!��^1c�)1�Gڜ���� �Q!�D�(CV���[�]��qb�F��?_Q�@F��[	<=P����pEv�j����~�'LVl��JɲxvT��'Q4F��9�M<�	�	 e+�Jy�i2�fF/l���nwTLHkԵg^��l�
��'6��v�)ҧ1�Jl�GkJ�]	r�R�P��xT��W@�Ӂ��Abq���\ ^�ipe�<�.O��%>c���R'�,6Z�5 K9��zA7D�H��EבR����3l�qZN���s�D��=�O:��V/ܻ7�$<`�m��(��a �"O
�1�u%� �$���`��G�'�qOa#Ud�?s7��:s���u�����o�'ّ?Y"H�mN���	�H6T��
5D��j1`S�
��{!EX����1o-D��ʰ���,�` ���R�m)�.?D����c8���$fU�wBZ�y��:D�P�'{��T�В-��9D�xʠ�R�N��Y�C̳\O� ;e�%D�\Ya��p]z��3��:%���.�Mx����G���9�E�+ =PA�ȓG�NE��Q���F.E2[}�axdY�̄���wh���MR��)0��٦h�B�	0'��0ᶠB��a"�*�6��C�I�m���E.����#T��hO>���
�7^��!�	�o�Z�J�f9D�<P7�O�+�j��8Q� ݘ �5��|���IrǑgf�uA!��&/�awm'D�胴i�=:�TIЧM����;$�&D��Ӣ�V���qHs'�<K��B��(D�,���5p��QF�U9i�̻t�1D��Ӄ��FB���E��n*��S�e1�"�(O����s��M,f���8fB�2WC��a"O\�wꃔCˢ��Fጴp��8��$2\O4|�T�U�U�x��O4R���:�"O�y�B	P�@H�!$Z<S_>�u��L>Y�s���&����4����2�*�O�'�2�A����+P��`m�,o� ������'�8#}�'Q6�р)@�,�2���e��<��'�<�0A,ǎ)F-Х�_d`Psڴ�~�$<�O��
��͞[�S�$�?`'��#��`x����H!c�2ဓ���:3����%D���nƭ:�6D
#b	]�,D#D���siO�^��U��䆥��â�-D��T�ГQ�|UX-� ��d*�I�� XD �(v��ٲQa�����h(D�8X�f���0���;,�9��n%D��cA/@�03�.�f8j	�@�%D�� �t V&�-MrN�R�K� �ޝ�@"On��ə�w�Z�z��,E��š�xb�'T�5���#��"�A�D�.���'8&<J���PV�7#�
:�#�'����w�Ӿj<0r�тD���2J<��e(����	���L�7{�Ԅ��K?���IԬ0�����m<�"5`e�<���-[���Z�g-V"A2s��`�<ij��[`dhk���9�4�4��\~��)�':z�xs�L�@@���$�A!{�J\�ȓ�b��DnJ8@Նu��D�]��h[�y����<�}&�l#�$X�L�t�hVGڠ_����g;D�haW�\��tRv$'j} �S`I|����IvNd���>
���d�Zv�C�ɴr9�dx���.e��L�dl�2�C�I�*�0��L�<B��1d+	2	��B��vYQ��e�&F���F�>:jnO��=�~zש��N�	q#ϺelD�R��s���=ys��2N@J	�3`S���D�q쓞p=�!Gī
���Z�	Z�+2�|���E�<��@2Yo¤8�)޲�p���,�u�<�p�@��� ��'c���I$��o�<�@G�{���G& w��q��P�<1$Y�>O29Sn��T�XI�%	P�<�e��S�V��e� ;-�\C&��L�<�g�V�@ ��ڐh'ɡ$,R_�<!� �4]BU�C��"Z��MR�@�<�돣+�|�dU�b�H9Q!Kw�<ه�\�l���{�-�>����*Yt�<Y�l[g4���qJ14�t�V��o�<�d�H�J��:��Q6ۦ��E�h�<)$e[,I]:���nɭ`� ��+HN�<����,Eִ��͓�x�N8���t�<Ӯ^*"�`�.�;JI��� �w�<Q�ck��� *K�=3�hRV#�k�<�q(đ\T�l����@L�p� �Si�<	*I�+��C�J%wz\��h�'��x2j�����m�)oF}�b�,�y��].U�8԰p�ߤi,��I��?�M��'��1bEB"����EN��� iY��7�f1Y3��+GJ��0d)�6��O��Q�*B!6����e��Y�8vpX�HFy�ʞ�`f��O3
v0����y�!;#��8#K+$Ԓ�;QR��~��'/�d �:�Xr�)s���瓞ē.�H �Ӫ�y4��x���6r�mZG(<���P�aC����Q��[d\�'��ɿK�>�e瘸z��H�G� S�|c��(?A�+�����K�-Ǽ�e5.�<d�Ʌ���r���L<�C�^f����ǁ?)]�d٢�PT�<9�g�s������;A�@)�휌��	W����}�o;#�؀�Aɀ&Rj	��ș�HOأ=��'3���
+j����V+f��EI�O���D�in�(��K�n|���U�"-�f�'�O?7m�)[��/m�Ⱥ"�ƍF��u3�OV̐`/A)E~0�J��QTuְ� ��?��|"�O0�#����;��C�Kսh̺M�a"O"M:Ec:*P@C�L��du��러G{�'p�FBG���g���A�L���O�	@�y�>���O����*���*���8S��ae �Kg1O ��$�=}fx��A9#ABaa�.�`,�v�'�4�B�4vX��u'W>ӧ�#wc��)(�"�f>�JqCR�](<��4��A��K�S]�T����1C1"�͓Z�X�<�{�'g��(�o�lZ�x1�[�`�.����HO� :M����7�0�X�ρ�~��@IDN�<!M>��O��R��$ݲ��3O��*�\��"O2D�6�9|:n�A��"x��Uf"O�PY�Z�I�!�%&u ���"O�X!�Y!&8*i;�K@�r�+e"O�B���3b�\s֪�."8�H4"O�]���F����-g	��I�"ObI����$�$���_��Yð"O�I+��ʐD��-A(�k�^���"O�,�+��s���F��*[�Y�&"OJX�gj˨w�8��� TH�r"O�����N�ax6���@!��`p"O�MÐ�V$b$P30h�/gz��7"Od����̇Ja�ݱ�&K�ƨq�"O�0�B����ÒE�9?��9yg"O:�s�ň#�] ��Bj��a�"O�q�V��	G;�����j�0��"O����⟗a�Tu�A��C8���"O6��'K�i�56Ǆ�J���"O5*��[7o��9�'օ]$��""O��ۢ%�Uɾ�J�K/>�z`"O��[�R�\Y�\�t�	1'��"O���'A14�@��ߡL `y�"O�ě� ��1���:��"O�����\��
�u;�"O�4QP <��\�q��;��2"O �jp�h.�t�����L|�Ჱ"O`�ः^#H�@�0��9g_�p��"O:�B6��=�}��DT he� [�"Of	�7%�@�@U����e]��"Od8�3g�E�,8p�"��4a����"O~HywHR$$��} u"1@���۲"O�d/*��Q����s����b"O %���ѝC̔a��8�|�30"O�c��2*qz\hêO;S����"O��aWy�0Ab��Gl��aa�"O6e��]�_�DP2CU�[����"O����1#��� ̀�WY�zq"O$��]Q�<�5@��w4&k"OL�ᱠ_�pa�))GNM].N�jt"Oщ@@>�ص����� "O��G��?7_l4`�l�9ftU�"Oʬْ�0h�<��B��zk�=��"O陵����e���;g���"O�e���L�D���/Eb^����"O>D @�&L	 O2W�P"O�L0�MT�%d9+uG%E�l�'"O����:�d���vb\�b"Ot���(&K~z�*@�\�5~�w"O�X�W  {+f�p���^����"O�����D�d��f�Fu����"O؁�W	�;�z�s��~܌]h"O�('%+?G,��Ga��2-ن"O�Ч$Ӳ�4��u�|ʎ1�4"O6��Fĕ�_� ����.��C�"OX�J.�M�8!�vF�;��y�"O�xH����"e�� �N�#6"Od�bWI�&�>���'ަb��@�"O�L5��4{8Mi�'�/r�°��"O&M��gM�"6&-���
�`���cp"OH��p��׎��m�;��p��"O*�P��W�w;�8b�O�8d$ u�"O���g�6b���F���c�� �"Oʱ!�O�e�9�7n�6R����"O� �Q@v�A�4fT!+S��1vA�X[�"O�Pi��ҺҘ���E~����"O�����8�$�I�P�
܁"O杣�(^�Yڅ5o�� d�S*O�}��.��2Rf-�7-���9	�ܰ�����<�Ms�*�=#/����(�rHS�l�G�<I�Ň,�,�7���SVD`���W�'��-��hˎ\�]F���ʦ}���b���)g���%��yb	t� �R�C�/��(8���x��R�Vh2��*O�}� ��zS��c)	Q���!�`�� ���Eb�K�*�DC�-/R8�I�X"&y�$�CO2\ц�9`Sp�(C�Oώ��VHX&P�����H�m��UbuL�cVte�$ѯPV�Y!i@9�t���$<D�q�JԴ!ʎ�w.Ȁ%H<�,4��O8u�'�\q�\e#Z�>	9mM6[����SH�!B�&��Fg/D���Ro�5T��x��Ş9<s�^)�^m#��X�T��h���ī$4�b� d�J})�A8X�H⟀G�?�g~��ߢA���"��U}�Qs�?	�+�.G�ܩ U���<D�_e<� ��ߺIV��y�O� Q��h�#/O$Qa���R�.\�ǃ�*8Zֹ�d'�?Ekޘ�#�$/�d��DX>@`ʄ�K<9�R�<T�	s���)4|ۥ�Jb&��<ѥ.
a*�
�c%�	]��y�(��}��[�mߟ|%�Y3_���~"�ekq�?�)�)z3$ ���̈́~�!�R)��!���g�B�+��L�O>�G�±*��D�|��~4ll�ǀ�W`I`g ���Wp� �Z�2.�\d��e�#z�{�O>�ScLF���ԛg*U�"J�O�y�K�-&��I&A�,����3�*%��'M<!2� � �8��Oq�6!
�'�Jֺ���d�a $�Q"�'��Ec��|��7|N�(�g%���I��@�'bHE���/}"��kD��o&���HW�u��8���78�:���]et#��ʍ��xp�I��*Г#&�;�����.�O�<rwNR����f��3ry��'Q�ѸF�6|u�'F��ZT�\R&�hR��L��u	
�'*�S��M+Z1T�;D���q�^{I>)@F%r�PC�/�':T�P�"�7X���ya@��8ǘ8�ȓΖ��uEf"@i󥅂1Q5���8��P 9G��O��3���k"�A#�C�$Eh�"Otr&F�P���+=�"�V"OV���\Uk�G��W�˗��y2�R�p��Y�&:�ҵ�d��y��M��A ��Ӏ���I��yB<y`�+G@Ѳ8��� a��y¨ D�T8�4M�`�3����y�� �RX��BQ�t,��  �y�f�y��t��&J�t uʛ<�y"e�0C͠���%ئq.��T(�;�y�eH�3�",�TLK.Q\z�1�-��y"�w,��T�@'e�f5�B��y��D�T4��䈍v_�!��Ǐ$�y�f#l� 8Z��o����-*�?ɖL ����DJ �4+�����2����a{��UC�H.�~�J�0��񫥧 > (A��.��y�f�
/�������" �d�e�O(q3� ��6��������t�j��w hC`L@63mv��"O6t�ՈIJ�����0O��%d�5]��|�>O� �DQ�^D1�1O��21�@L��ӕ*�KL�@��'���Ah�lpLݒ3� <���@��S����v��.>�����d��GV��yB"��(��1�L U��1iQ����O��
��I7�Z��6$�/H%��U�f���J�/D*I�`�*Z���b]�@�fA\���<���{�n ����%!�\��/KYy�,V��P�@�K�*i8},��O���"&�@�sᮏ^�"TJ��یSXA��xH<�
�.9��[SM}�8��$A�U��Š����8�G�B:N�$9�
X+3��{s�>Y�wΨ��u�էP�D�a�	�wˎ�y
��5J�M������a`:pO8%q�I�mL�P���@
�C�$�R�đ�?��i'�)���W�d*�,N��z��X��|"?��f���pY����f�bU`�π `q�.ջ	\�`m�<di�T�xQ$��62l`�ڰ�'m��S�ހ�Ρk�d]}�H�[�O8p�n�*&�~�#v�]�7cq��	e�D7��4!j 8o���D�
xS�I��D�x�� �V����� בC��}rGl�z �s�ڟTOZ�t��h��A �S���ɂ`7}?�`-Ӏ�B�`�b�R��!dÔ�{��'M��b֡�&
�hsB��3&��HQC͂K��y��@J7'�(C�(
���ɔoKB%h�������d���i�L�s����� ��?��/���իt;JL�C,���d�mC�9R�
�`�^`*�����ĕ6@Ć��t&#<Odi8��N&Y�a��+�1:��0�Q��
��[&\樑�eD(�<�d�I)�0�d���Ԅ1�kԪa���ʅ(]0�yb�[Qv�Zg
6_�H�A��I9.�5)�/t� i�(�WR���J|�>yW�T5=dE�B�b]���n��@�K�(PYF�����#2~�p'B�2eZ�I@�z�CG�u&�&�j�ǟt1O��{!f@�`�"h�blP�x��I?f��@�OG�'��LyV
U����:�����@<kj4�v��$Yhk���h��"MDԤ1@��'�jr���b"F���ѡR�%s�'��;A���`���@L1V2)����@�X3�Y�B�84{�l�A�&-J�6��!�I�w�& �u˟aH<Q��ܠVb����� �R5z!N\2�%*U�X
,��9�j#���q�]�Sh���Т��B"᎝ݼ���4�"���)W(��R��X����w� �<�`J����E�+*V(X�g��8B�h�#L\0��BB4x�*�q��K"�	���j��$vL�r�%Z�#�X(� ��0P!\�>i�AT)tR��`��(�,3e�&sJ�H�
<A2��Q�HD7W� Yq�Sw���+��v�\HS�K���<a#%�-�yu��w����^`?Q��ө^�K6����b��p�4��q :c�R�PЯ/�`�@s�K�L�2p[�H
Rn�{�G���x"�	�<x9)T��l��y��D�f��@ѡ#W�G�D=ʖ�MKZ|*fI	�6lM"m��a���ŧ�y���P��XBⓀm��5��l͹հ?1�
Y��,��$�'/ <򄬋������(JGv�s�B �Nʰ�ra]�ɁI��6=�қx�������Q-N*Q�8����;��O pbp�Ǵ;�J�� �ا�
�;�%���~䂴AA�{�LPQ	V�<H��J���"�,��<1�K��5?ޅb�&�q��]�E"sy��Eα2e�
�D������g$x7�ǝ'/%�����ľv#�l��'6�Y�G��/Ef�ܠ�I�j�.�;Ń�~�^���O�Z\�4i�?����}i
iXv�H�xQ���Qǈ�l��b�'��G�$27n�(�A�C�|с�O]�p�dUc�O�'���Q�E�Q�~D�C�ǕN~�Z��>LO �)ԃJ�>A�	(}����ǉV�N� P�$2ޓO��d���� U�!�>�)"�@ U��������л4�\?Ϣ`r�A� E&\y�.�JR!��A<+�0�P&�J�̓�m�Ma��\I�ɏ0�"T�}2v���]�Խ���E�(K�\�<I�Ӕ1Kb0����nE{c"�f?Q2#�l�Ұ�W:}��� }b��ytɌ�d@l���3Q�!���f��2	J�@ԁ����y{ ���𤟻lQ��tmL6�<q��@>m�Q���6��mPqO�}�uO\�.����,��m��d�2 �;�\8�t*�xb��:I�L�g�B�<_�%"6aǭi'���l�;pS �೅\�crԚf�ٻJ�T�s�E���Iz�i�2��P&�)�%�@+�8S�	9D��ЊęF��@vI
 #��$s���J�Q�M�d��8(�-L�Vd��i�H��R,�B���'����W=l�p��B-5E�X�ߓ-о  ���^���ue�F 8�ڤb׆.��r��cTR�x��Or}��K.oa)Ó��8F/��PrN��̍�/� ��?a�E�31:L+!��8V��x�O�$��a�[	Z@��bp�ȫ_�65��0{aX��U��n<1'`�:��1�����Dq��"%�qrp�S(޲k��u'CZF��Y�Л|Zc���ǁ+"hZ���Fc��'<��r1��uJ�L�G�O6c%B0Q��v� G��3��Ot�0g�H~1�O���W���X`$V��PT�'����^	AS��n�}q���{�]��+��cS��+�&`�ג��<a���,'����|��4�'d�&~�<��W8ZL"=!�d	��)ag�mY�� ��A$N!��T0C������Bq�1��9 �L��cl2OX�:��Ӓ��p�H|�;B��|y�fǮadȴ9�HϜ,�
=����=ᡧ�
��L��#��l,�U�I�|:pЀ�M�+9�Ӻ�s�Rf������&Ǘv@��:D�>��8FI-D�l�!��U�=���I�*��=KC�<�����!���k�l-,O� <5��,Z:���J �	�e�}3��'�acNR/�\JA��#NobpU�Ǝ�`B#AeH<A4͈5�	v��j�Tc�s�'�Us�GÏaD���~��K[��&�0�Z*�s�<!TI��`$hYZ�F�1]B�����\BV$h��5�>E�dAG�G=�]�1��*R����:q�!�$�6V�Ld�$/\�.""YBჭs�	�AYNP�`ĂGx���GU�k(�q�'�E5�\�5�?�Oh�7b��U��l02%��Qh�
Ga
7Q��h��'��)iq�*LRRPYP+E���*�'C*,;�ϒ9Khc��J)?�pli�'0jeۡ��]�������*5�ij�'�x))�[�A����"1��S�'L�5�b�_�v��FǏ2$�Tu9�'���9��Ә��� ��Cz��P�',(������y���6D&�"�'ṮFO�*F�X���$����	�'\�8��D�`'ɂ7DO�):2���'�t��s(C�͌�D�2u6�h:�'���ц;�,�F�����'~Xa�e+��c*��:QOJ�	jt���'B�EdI0Nz4����9u�����'�����jː2����g�43&�`�'�"���)NZvf���cҝ*j���'v�0�sJ7V��-[��5	t�5��'��2T�
2�%�%��+ǖ)R�'� 刦�ԡ,A��	��	I�TE��'�p�g�ǠUA��J�Nܲ8k����'��̩�k�?�ph�5'��=L@ �'�p�ZgoG�v(i
 BF4BX�
�'����l�7��z`��'%��`�	�'������Y��X��ˆ1L\h��'"2�Q'��\��b��.��9�'�T�1P/ۂE:RL��	Z֩�	�'d`���eke�KS��R��}P�N"D����/@?��#�O�?|d�U�<D�HЂ�F�N+����
Q�l;�/=D��d� 0J\�5����%,D��
��сR�,�!$��N��ٻ'�*D���4a�\ɮ�����8k�b�t�&D�أ�l�-�tC�]���P�$D�����a8��Z5���O"D�,�D��7�x�
�N>�5D��!��q�z����L*E|F���b>T��xA.Y�z����&����"O���0.Ƅh���)B�c|Ds�"O��s��0x<<�v��w����"O���d�ʌlג�(@��7{���aB"Of��2b�c�@e��L��p3�=h"O�M�!�/l&`��5	�#^Cr�1"O�L0V���k/���j��R)K�"OцT�+W��C��E�9��a"O�$W��-j�ͯz{T��!G�Z�<!����J��U�AfI�gg4���[�<!�'[�Z���6I� ��aB�V�<A���?r���B
�z�4AI�H\S�<�&�1H��:��I��8�r�C�<���ځCq�}��"�� 0����_B�<Y��L�>�G�Y(b�� n�|�<�pE�!\=�k5'��(����C�<q�B��:����&M��**�OJG�<`��CU@K��{nhHy�K�<񁣗�zH&H�2�L�d�u�t�	F�<q����(��$"	��<Lq'}�<� ~0S��T�C'�%���T.0hʥ�"Oz��֬t�|�&bK�7Gh���"O
	SA� t�!3�N�6LZ [s"O�Ly@��#6��ƯF�WLA�"O��JA��+�萐�Y��<y�"O��r�IH�DD�C���p����"O�d�����/e��r�G��Rv"O�� k�2}$���Ӟ�xR"O
Z�U�p��5��3�^���'�hk�D����i"y�Pǧ�2��ӥ�yBl�Q.*4qQ�����Zk�0�Ob%:V"�'�T\`��i	�@<�@
E�݋{ *���"m!�d�>Q�ya!� 
���Q#w���#�nX�E���P��G��'Ե�U훜,r
���*e� E�'�����|�8�X�̜nE�(���q.F�7�ҏP�������b���9&��,��5]}�̄�I2R�H`������C�L)E�N-�E	A�
�&�I��C�<y�HSZ�.J�-�&bl嫃CC��}p~�  P�<��I ��i!<�8�@�M�}�@�HL@�o�!��;M�|���X���d�E�4,:���4IƊS��rAX��D��'Ңt��f����3�h�]��0��'8�X���`�J����E���h��d�Y��5F@Hӓ�}
Q%S L-p�5kF�B��I�[�jX�`ʄ��y����/d�������
,�%��K�<1��5I�t%�
�3L���B�B�jT�<���R�A�fH��h7�)E$�yw�WԄ�"�G";0���X��yRMbb���Ā�li�%PT��`׌�	��F�lO�O����ƯmM1�¤�>^��%�F5���;c����<uNƏ0���3�>��=E�vP@�(��ڂ�n�<���ۿ����U�-�:x���|�.�,D��Z�y�?
`h�f`pz����zל̊��=D�l��.ȣFx�-Ң��1�F�R�W4l� JL�� E�m�g�$��@8
�pFS�U׈ A�A]Y����gK������sJt9h��1e��`(F��8�8]�P]��9)!U���2�Æ�G^6D��ɡV���
W�$D]�I�Y<I�Y�g1��0W��	��B�Ʌz�H(�ϕ�g���� �;{L�O�������|BH���I�'>2� P��U��N�	Vś�-�!�$��5�J���M3J������t�vdx3�4��Cv�>�F�Q3���L�<���# ���u� Ԓ�W�?s��$�[9yP(�ȓ$���CIWC���s�ɳ����6`�P���^�]C�\Yc�.5{VD��@�@�Z'G5d����5�ǰUƬ�ȓJ$(��G�E�pn�3�ЭKY ��O��%ٰ�!I�xLa1C̩G�,��ȓ[�L<Q���Nsh�x0̏"/�$��j�ƈ��A4��1DkH� ��U�ȓn�bg,ej���B�TB�$4��sб�JS��%�SA!�2�������C�d��T`�����ȓv\TIZ''S�rܐ��<?k���*a~��GE��<�H"�N �T����xV� z��'P@})���3J�I����6�2ѓۓi5z((�Fئ�~Rס1�l�`$ Z�����	�y�)�wh�0���Rʮ�9��ϝ���#��U9#�8j>����q̡�s��!"��t��a��C䉌^�B,S�6����k	�-����k�0f�:�8����R�?�3�`)��jq��]��������d�b/������
LC�`0�ǩ�*q�k^�y����
�!Vx�PzBEB*=1Ob�����5`H�V/ܿ|����iѐ	io��u� �	7�P�|����{0HH� LL�l(:��Z~"A��,�t�@d�'���ì~�J� �	�G5���)O�1���3 ��h��m�꒟� V�Gm��L���Dcj��GMA�H��hG�B�x
� ��0$�_�=���*��ӤHT�iTe�F��]���'6Qj@�ԘCP��p��ކ9����O���ʌ�'h�����F����$ɒ�Ҹ����"�^���,��a���26䝸�M(�����N� � d
<�a'?*�o��H�* �W*J�XxѢ��y�'�*�꠨ޫ,;j]��3�����(|r<H�/�
����_
��dU>0�� W��<���*H�x%`eD��4x(\��My���"���� ��:E5z �}�����3�8iEDO�`���K�S�M�@x�E�^6A�B≻∵P��A耉D!�.K��'����T
,O�����ٹmґ�I���;5Ҍ�))\�t(�5mˤ4���iDШ`��A����'�V
>o0����
g��*�.x4f��K�8D���^�Pf�AB�ģ���p!Q�4O!�Z$���RgB����3�-�"��,l1�%�',Hx��iqER9��,�Fn�:N�h�C��$�Ol8!�E�I��A;:)@�Ů��H�2��'�x��D▕@���E�k�'�eH��#^�F����ɛ+���8
�'��h�"��tQ>�R��
�a�Qk�'D|�����b�S�O-�z2p\�5e�9��	�B���y�䜥>�Z)B���27m2uJ���_�gk�p�4<O��o�.`���F�
� ��S�'��#n@J�f�02�6B�p�k�U$^�� *�HH<�W��mo�����u� ��� �]�'t��)Z�h�b�~b��X=	��!�*k/ڄq0 Ul�<!`D���@w�� ���3ܟ�c� �r;��P�>E��/�4 �4�)EG]�(���x�eM�B!�ƹ%,���Η�)3��ՍQ]G�ɻ]���+��Dway��3xv�9ǖz�A�դ��>��D�Q��뙑�؇�A>O���r�IQ�D��C�ɫ/:�!�`b�'���C"�R6Y��=a�*�dB$�(�I$��(n��uq�&v�l�����9x�B�@�(�5�E$Ez,0�)b�$�^%R�y2G���)�'< �8k2@іGr�T��h�0p|���
�'����WE_��d��L,$[�O2p�F)�4 .��D�*h���AT+��Rb�	�����Ca��@%�S�4̆�cQ�ߌX� �b @�'�vC�I�@���T�G�
��C� �O�zC��;sD.Yi)!*������FC�ɞ@t�r�J6XAXq&P�K�PC��.0��ڃ��=�"�AH�$9�2C��1p��A�S�)	��;��L�%�C�	�4׌��5�e��ze�����$��5Ո@�dML�Q����K�j�:�$ϐx� �:?�h#�5.����������O���q�[C���>��vi�Q�ЊpG�(+k�\�1�1D�t����*6T�w�B�TT��'��Pa�a�>X氲2�>E��HN�?�����V4y&`��ׂъ�y"�1Ґ�c�A�~�P��'��;��	���"wO�u�ax�#XI��Zp�"z�ZX:G���(O*��cؘɸ'��L�Ѭ�'�t	��i�4�I���u*8����@<Q�e
>y�ɺ��)<)�����Z����,��Z���QǙ�nF���O�R�	�T�6O�W�����ػ�y��.����ߜ8��X�q�	�?��b�*�����4��I�BR��Cg�_��rB�"ņ�tL�4y�ᅅt����DH�tJp�(� �M�Ս �-}n� �
�Q�(XI�L��#�FyJ0�?�0<��%ϥ`Ƽ@�!LZsI�!SE�� L0L�@/�HĈ��<l��O�Hr�z���t����Y��p�Ѐ�W/�x�_�(6��q� �eܸ-��,T�}*p��"
�'�����Q &���X�"!t� �7���D0�.���y��:�t�rF�(�詡-��?�s��/`���ڷ
 ��/a���ʗ* �$�0�(r�	Ǭ:TU��H���{b��4�0yp�Q˦q�Q'��/9}��"��K��2?�N�&@�E�ϓ1&%�a��~�
��Q�c=���?)WG;"lTb+"ғ�����Ϛ�Nݒ&�L�J|؈AO�agP�n�� � y�*�� M���c�)R��'"�K�'�T�f�'>�=� �y��H�4�� pf��A�r��G"O�0� ��[�p�Z
���$��'p���u�F�a�J��O�.E�M:j%M~�3�s�0��6H�TnN�x���4�ybMѿ�B�X�h�0I���h��[���$�"j�<�s�BE��<ibg�(n��ӥ��VCyh�d�px�p@�$׳ zB�ZIհX�8�i"�K�m���#��1�!�3N�(�P
ӘF�B���*�ў�§��%@:���i�/S���A�R�<��hw�!�dX�8��U*��	oln��S���}���q�������|��S�S���H=e��U���?��!��1�n9 �`G.E�.�ca��Ms���'��M����?F��y�J��K�#�nRh ���c��p?C+PP,�QAh�4])���R��T8��?D�tx��ă �wŅ:z�i�&b.D�|�pH�o7�,�����g��9a�/D�|�7�\�D���M�I���H*D��藯�~	����Z�Tri�r+D�<Y�̺KX�*Ao�Y��
��"D��jU�~�+ǏX&s�!���; !�߾4(=�$nI2�����I2w�!�$>k[�u�'	!b�b��r�EW�!�D�k��A�QH�3@Œ��!���� L0��;�
������!���P\$���Cݹ�R`�%b�39c!���9�6�s�־Rn��9r�ߦZ!�3r$�9��0Fy�I �㇒En!��C��I땊ܹp���b�.1�!��[4#ڍ85�A	% ~���	�<!�d;7nⱈ��P�w,tIz��޻R�!�Č3��P���J����E�sP!�D��a���rrhK�L`w���W!򄗈Nf��֧�
�$􃔮�}B!��T
�A�AH�Q�+�?Bj���aG��� 	�z���"�E	g�ȓ@mr SRG�8#������w�m�ȓ.6xz��ՅC��)р	�f}�������΁8��=+S�j<��ȓt�̄z��
W��5�;񪥆ȓ��9�i��|�T̈4BX;v`}�ȓZ
�񠐈��u�D�pBJ��+^�ԅ�6e��h%ǔ�%h�A(�	���ȓ�\$�BhŤ+6A��L[�9�D��ȓBb�]�@)�����K��0Y�N��ȓ>A�T�6!ӱ!4e)��ٲ$״X�ȓ$U���d,h��ȔJ� 1@ ȆȓW7�\ȶ�B�NLp 1��81�����V�Ȉ���4	��e��3V�d�ȓoY�ɒ��7v���6��-W�Hy��B�q˶�߷�c�I9�Ѕȓf��,2b�� vf�Z�O�N�,�ȓI�P�@�O,"�q����'1B���!+��SP�7muXDaq���8�x��N��J���$�3�䤒p����j��W�	M��T�2i�	v�׈xD����%-�a�,��t� HzC�T!g��X2�J0w��A�/�$75HzV�ͥ � {�����-Id��C䞰_�����+�CߐPH�ǎ�M�߱v�~�Kd؟��i�7�6�*
|����Є�	5U�R��@�U�8�~�$�[z#}p�T�~��H��8L�ԡiуH*�J1�/�\Aj���'<����S�Q�`���;��ܛ���G��5*�:k�5��)iʄp�!_>�ȟ������+�q�k^�R�����A�Hh��I(��A�7�ۘ
�>y�O��:0�Po]DU�G!�4y�Aj#;O
��y2�i>E�/8xhb}QE/B�O��ˀ�*�>�O���e�~����/�?�6��"O����C8l=��b�G++�� Z�"O^`�bB���<S��7?�%2v"O� t��k��W���UŽ36��h"O�y:���h�,=2�9r�"ON4�"�\�%�ґ+��1&�j�X�(E{�􉑏�hDz �;����B�,M���'�?���-R�i�e�fR��>��� �	D}r�O��T�
�0�;��M��OF#=���	ւP�<A��)`/�d��OT2;���Sd����D�PR �)9��Q�b��F�z��Dh4ғ�0|ʕ��]Ȇ�3�AE,E�a"-�_�7Mў�'?������4]�$ݭ{m���<�����^�W�p�5�4��\�W(�>z��J��n��6���(O�d�!d���i�6`(� &��x�oB�8�l��K>	�O8�n���1.��<;�鐝Sh��6+R{!�R KH~�#t*ڗ#NV�R��ԫ�!��R�*t�Z�L�� �.Ł��E<n!���$�R`���߫N����c�	.Q!򤎗/�\�F�W4x8�p��I�3�!��G%e�,���Ȩ+!z���1 �!��/���y�灓:�IEGV�r�!�Ҵ/�:�ئk��~��BH�T�!�/I�!x� /!�&5�g��//�!��Z�	;��%o�� �R��DL?g!�d�i!n};e�N�1�N�{���Ws!�D��TW�a�� B8A���9TBBn!��]$>����%c�R�R���^U?!��=pA�YPF� ��LW0f&B�	+�\����#��@)��H�ƞC�	%z�݃��
�6\9"�z}�B�ɯ*tDՋ�G̪k�R1
��|B�	;R� \KF�֐(��YHS�#);*B�	����� +h �)���.B��!Z�� ��H�����i��B�	'����ha�-E�\7xB�"c=`I��ߐ��� �	�!xB䉍c��ܳ��˲IO���pď�	`B��D�F(ae�<G��9Ѩ��c[�C��>p6�KTn�Z����Ϝ
p�C�ɺk��YJ���&]�°ȣ�-=D�C��df�E!�M�4�R���a��DrC�I6QZ���GM D)"����ZC�	�|���c�/Z%
a�p��g�]�$C�I/�X03`��>:�x�F3[`B䉕�8Hإ��-G.������MFB䉅PP��oO�.(�I4i�@(B�	�z��8g�M$=$Ȭ�m�r�C�	#F?8��F���ytA o�B��2PT��K�5��(��M�;#�B�ɤr��x��	͢��P��J�t��B�ɒ/]ܜ`�)�*u�A�'�U,fB䉃;�~���F����DsB��X�C�ɏSČ�Isa�o]�����R�C�I�l2HBpL�X�D%94��B��J��`⪗1f�m�������D@�,}�#)T�mr�h�f͒!�� +x� �Ņ�XP<e��lڿ
!�Қn�*$ �K�R� D�sҜ�!��� H�IK�j�+��xplªP�!���%�r��Ƭи+�ڴ��8�!�ʽ6�rx��� w����Ŵ:�!�	(y}�J��Δ3L�1
6�ՙ+"!�D� ���,�.K6rM�F�T>\ !�"[KXt�BC��fPxu� �`!�$B3 �ޙ����5?4��0̟�r!�Yr*X9��J�?3��xCjC�K�!�� F�
 ���������S���A�"OL ���Á��K����0��2�"O4#�NR�,�di� �ݷUs +�"O")#`g0f��]`�%�6r�~(P"O����.Z���Q"�}�J$Z�"O�p�8zQ�@Z���-/���"O �
������[�/� �Z %"O"E�b ��g�����g ���"OxQز��+=��u�4Ý��I�"O@}ڀk<((�i�� u�@��S"OZ(�`D�wz�� +�+'q��"O.q�R��
��YF�8m;$���"O�Y�#E� �IK�jN���ã"O�ak����	)�Ȣ��O�4��r`"O8���%�S9FeKw��nh�*'"O��Y�^4b��X����:T�=�A"Oޠk��άe���A���	'"O�q$�1p��P�Oԭ}�0��"O>-k���)Bz}!V%T�q襈�"O(E��#C!1��Y��EI�cF%C"O ���:RRI�e�C_�x�"O>�Kר��!�� 0$Ke�(!��"Oʹ�+�'�Ы��hȸ��"ODa����"�$V����"O���<%]�Q"K�H���#"Ox�����QH(�`2�����V"O"5�u��xP��1,^�eh0��"O�8�i\6�:D� K\|�hC"Oԩ)3�K�;޹p�X�zh�@�"O��q��4����+c�\r�"O|�k�»p�ᗈF�G��AЁ"O����6ܐ����N<��
p"O9#m@�>�Z�S@k߻o����U"O�AQ�C
	Z�~$��i���n�cF"O�M#���vC�u�Q��50�Jv"O�! W�<k�]Q�蘮o5�X�"O̍"���'e�t!��Y'd*�rW"O��B !�n����&才=`,�p"O�,0�h�#3sfP궄�����"OV�zaD��M�ʉ#@�2K�ڀ�f"O.�[uH.��$���{� hȳ"OZ�[�H��%H�ƍG�&�б"O,Xď�!>�#�X����k&D����gL�)������]'j�H�j!D��b�J�Xy���R�R��d� D�����:��%��N��b�*p�"�=D����FӇA��@���Rah�}�g@'D��� ��[y��(�E�l��v�'D�X3�[0SyhP�!�����;D�`�w��h��uK��܁E�^��ȓr2t-項�(M�a���71�I��/'*t�w8��4�ڊ-����>�R�!p%�%�`8�I̓]}�ȓ<�ʱ�"҄Ij��!м9� ���X���OiAn΀n��I�ȓ�$m�#N�A �,�ǖ=�(��FR�1��e�8i�4u(��=w>d�ȓRZ|��g�Z�p�����y�l��t*�� �ԠX�D��Ƙp(^������6��G6�+5h,��ȓB=�'jS�b�H��U�\��^Ԫ�37�q���0eP��͆�{$<�4E��|�ԘВ�N�\����)Vr�@��/M�Z(b�B%|���S�? h�x�m�.-����6�p��"OZ}[��N0�)�u���@�"O��ړ�єN�֡��S�E��p@"O��s�_�G�Vp����2�Va
v"O��ARDQ�l�d�c�OR�|P+�"O,YZw��!UJ*�qb��j����"Oy�Q��t^��aR�,E �(�5"O*PZ�(�h�Lـ�<BA�P�"Of�b� +Ί�(g�c2����"O�i��ґtLPM�&*Sl q"O��P��60u���9V�4�g"O��8kE�X�803)Z�+�(���"O��A8���C�4��{"O4�H��ˡn�ق`Ō=&��Xے"O�w�d�T���W�X�Za��"O�UXǈ�����P�ju�q2"O.t�X�`���ѰXSb��J�<���I�y� "%/#�p�^�2B�)0�p 4꓋^��9��%̉4z"B�I4#��FkJ�@B<1��V�@C�I�nt|��7egz�:@g�� �4C��h�m���Wo�
�z��@�Vl,C䉓�i�T ^�vsި�n�+m
C�	򬱲ԮS��P��͞�$��B䉎��Y2�?��Q�͜�a{xC�5O�(���٨ ��S@猧;�XC䉦u�6D��V�k�-!ȫ_C�� 2���3��T@�'�ӗC�C�ɚ�T�6�����Ti�E^�C�� 	�'��%4�{D��-
h�C�I S,�a��
7�E�4�O=�C�	�6\�C��R�H����K�NجB�I���)L�K�2�(���

�B�	�V�Р��ˀ1+��0�O
�f�B�ɲw2X!��Ŕ)7�Fl3f�F7X�4C�	����0�H1f�L���8bC��@��9�'o�.
��)����,C�I7�ұSU�V7i��XR)�L�B��$Ra�4h$�E5=3�h ej\�e��C�5*g�P9�&I�|�td���W2��C�I6�0<�L@��&�c���$�6C�8�^@�v&͑t�V�ff^�2f�B�Ɇwt*��
�wS8��'�צ�|B�I�j��1BݾZhS�┰H�B�&o70�:��VA�h�D��TzB䉪5R�3@��|�0H)7�=6�C�	��\}b',�$��u���RIjC�I1>}X�ز�\�En�1H�F�9~B�	�Lr C��6G�H� ��2�C�	�)� ���]�P�̲�P0*�B�>��H�a�ƩX�H(�+ܖR�C�2!������N�x;$��>�C䉂&( 	ٓϋ�7b(�2"��~��B�67�lhX�)l��8�BӁkĄB䉉R/���'O�<W�)"K�2e�B�	�y����#$L�d��Ah�&,�B�ɒ#�d,��M��|�� 7a��nX&B䉰:A�5)�P'U`)0� 4#B�I�=���3H�,e\6�Ҁƃ{�C�I�B4�Y�1Α2a�\�s/�O��C䉶a�΍B�s��|12�A=@��B�I�/V�|������S�k_h�xC�ɘy�ptc�)�%4%D�×�?hbC�	�f�V�2��h�T�P�(C�)� ���Bi�._�SuEˮ=�z	KP"O6i)Ţ�j���z2�Z�{���"O�`��T�#���C��c�fE)"O��	.�x��y�&"M�4�����"OQ���+q�*�`1K��x	�"O䙩FJT�H8$!��'`Dp0�"O� Y�B�	�x��Ơ��9%�2"O��gT<�����(�J!�7"O�E��HW�xt�3E�$=,�A�"O>mҷ@|8+�l}:�yU��k�<���G�p�KB˂�4lA�nm�<A!�=��0�g��$3���;օBg�<i���:��[�aR%	}$<+R��b�<�S��7�
	A#�{la��N�j�<��
�8*��s�,W~�4��6��~�<R�8��E�(_�0!�P13 Eb�<��A @  �d   
  ]  |#  ).  G7  �B  sK  PU  *`  k  �u  �|  ��  C�  ��  ە  �  s�  ��  ��  <�  ��  '�  �   `� u�	����Zv)C�'ll\�0bKz+��D������b�FN9�y���y�FJ%L+pL���ҳB����5�� KrDE�Ƨ�7}�H�!A�i�d-Qq� �T�nʭr��	W�T����ۃ_l
e�N�E�YB
�"sIAyaa��C^꽂�%O�^���Rw��zqB��;9�V�����?��
Z�?���Ke	z�-KDL�[E��z�k'>�Rk�:�@���xOT7��m�x�$�O�$�O��d� Y�浣�e�-'"�	�:B]��D�O<�l�N�nM�'�b�6��t�'L2�����' P `-�YD��%�R�'7M�O�ʓ�?i���Ϻ[�̧K"P��
%mj�3P�N�-�$؊���
8(�@�v���'rtR��*G>���ɮJY���N�o��H fg}r<O�⟐��N�[�б���<E(Κ,�d��G�|�T< 3���ڴ�?����?��������|ލ��K8A U�@�'��:�F�O<P���	�0nZ��M��l��.��>�nڝ��h���@2�!�%�(�"�ָ�����dFs�L�r���rK\�F ��|��p�M5j����8 P�m!�JT@:K��\<Lt���.6�6M�ަݻ�4��>�~���gS�w�:P�쑭l�|�B�� }m訚�i�Y����H? ��42�����ѕ�ԱW(�7MGۦM��4y�Z��7���`��Z>|�N�I�Y�'br�CT��=m�Cr�b nڑ1��A"��6��!���N�E�J}R��]�'nv���د��xFʐ�53�eb"iGZ���q�4���#m�j5!P�S���x�ǌ���Qu.�] =[ @v�h{Dgy��p4�i� ��8����c����* �'��O(��)�=}�|��CY�1�����Q�7���CŮ�O4��O��)�������R�.<~�x&��OB1+�R+u���� i/;��`�O˓�?A�����S�_�l`3�̎G  0��i��8g �vesǉ�58l��'P�ف��%^Td1���p3܈�"�̞G��iť�LYt9��G��� h��܌l=>}�=aUn��$��4n$剷WbZ4@s-��K���B� -��d�O��d(���O����O��n>�օ�fgd��"�O.���'�2�O&�oZ-&��d����3P��5�����zڴ�?y�i<����c���O��D������,�O2� 'k�1wK �0sfF����A�Od�$P�	�׭QV�HA��K(w, �'��i;�*]�B�c��;��W�����U���֧+m�uB�a�>x9��Y1K�"Z'R-#c��?ձ�i�.6�������S���P�7?�q������4ug�>��',���9�� m��9�,K�)�B����F�'�t���]L�àʿw���@��d����ش��O�	��� T���D�M�,������?�)O��2��O���O���<��ALbQN���o��4�е��l��?z�,��c	>�ʽBs�ܠ[ʺ)�(�b�	M��ēcsN�3'�H/=��z���D��A�6N�BPۀ�is�ccИh�ATY>u@`���u��])/n��x�C�1�Z�I��_����n����d��e���O{�3�D�q�fH[�(Ƴ(��%Ra>���$�OFʓ�?i��L���t��J[\�0o���%�"��<�&�i�7�<�4���ɭ<���˳��0S5C�a8�Ю hl�r���D�O��<9-���S =��,{4�WU�Z2��C�h�I��}s�qV�V������;KJ�Bs(͛:h�s�.��o|@d��	)��	Ӄ�&7�(]J�������ᔁ��D�pjE�C$>@Ñ.�)PI>�[���!�����-+��$:�I��l�R
G��N8�ƊO C�j\�I����	@�¤B
�:�P�	f�C�0 ��h��3�d�����4��$�?Y?��'��FJ��A3r�.E&���Z(;���'ӂY;��'s��'�jŪY0��@�2nh�� ����p�R�28���ˢj��:��'30CGO�D~�	)�`ٹw���A�ƒ�,���Qdʾp�"���O�B�Z�ȉ�D �=Y����$�ܴ
�6�';D(H�! �r+2�[!+M������W�\�����W>�xW��K�ʔ�a#U�T}\��U",�O�ou�<��h�S"���t�*VX�R޴���aa�n����	]�d�����&�f@�$�o$dX`�\-0���'�d�H5L,Ac�ϖ�¨@��M:+�X9yRoݭ1O��х����P��D;?aS�Gc]��o�-o45�$����aF��!u�D-��R�[�tjp�����X�n ���D��*o�n|��$>��|��m*oFy9�� Jl��Bj�w�I��(�?��y�C��_@�yp�(�^�G�����d��3���|ӂ�Ėצ-�ߴ�?Q`�i�2(�O���[F��'L?�< �e]�0��6��M{(Ot)���������O��d�<����&V��sǝ;&=@��gŜ8xN��
���1��dO�E���rY>���r��+q/��Ԍ<&\�ɦm��vC0<j�dZx����$P��bE$�3H\�S�-@��`�q�1���\( ̨���6\�<�IÊCզy{&Q�`ӵ��O�b>�$�OD��׷J ���"�_�nPq Uώ�Rhf�$�O����O��$7�3}�K̕X��}(�J�D��vK
(����ݴ�?��i���O��dY>�ڷ%��\<L a��=�ZE�%��ڟP�t��l�I����	����O(�$�X��X�*ׯ �X��ɦL����IBǺa�ab��ch���wG����O�s���-�V�>y������<W��pIK2�}�TJ��r��U" cͪ:�R�D2�D��:�X���KwJ��ۆ�*��P��'�l��'`�$��<a��ʓ��ğ�E��A����:O�4p���;S�J�Ӳ�4{��➼n�?����<��._����l=��C�hy"�'ML6��O|�C|n���i�R�'�0�p�'�?%Hxyp�ˀuP�P�'l����[��'4�g�%l�HP�1���S#��k|� �=����mͲ�(Z�5_���U�ZM�`���Gm��U�ᔟ<l�؆��5h#�XeI�'aRx�t���vG�q�"�t���Ǻi���N>10��ǟ@�޴,��ɹ*�8���B:_r�H23�Y8��O��=Y�y�虜+8����O(Z�8��O>��'�ў�S>�M{�h��+�2�rX3��V �4%���\���7�4�M;���$�|2��(O�1y�`���P��Q��Z��?��oͧ<��q3&(L,g.l�öi0���b��?v�BQJދu�m�w�-?w$���X��S�	.��T���eFJ�Ζ=��+_M�@sE!U>G���i�� )Ҡ�~�i����Mc��S�|��icl)�#[2��۷`Iџ�?����ʟq��`�]�P����9M�j���|Ӳ`mZ蟘B�4�y�˄��r�G"����:1��v�'���'�&D߄���'���'��7�b���/ �jl��*��8*���'m򇔄 @*x����������#�P��/	���D!��Fj�Xp�۴j�(Re�J�g̓0������ l��p�X�;�|)۴_���R�X����j�g�ɋY���Zʏ	<8�{BJPkQ�!G{2�'q�ё �.7q�Y��\'x��a�-O"�m��M�O>ͧ�Z+OV�c� 2����2��<��k��>*�D S��O����O~�d������?q�O��xQ��G�)U�x:Ä�L��W�/Dn���q��;�duQ"i�!G�lh3��S�(9Q��Ѥʾ#Ϯ�c��Pbj���e�+���3W9\:-A�dD,
T�L��pUb�F^I��$�2IK���
-��9c��,4 �Y;֬�O��l�!�HO*#<9a,��'j��W+��"��檑y��x�<��2,����v��-R����d�N�I��M����$��HЪhm�|��ʙ�t1��9#��!%vy#Ą�?�/O^���O��ӘS � p
ȐM���@A"P3P?����P 5�P�mN(W;"q����*��O�-`��ˀV��o���Iw�Ƶ !��@F��0~�=���.j��
@���Vt~��D�0�$M�Vx��p�nP�'�`E �3d����	�(�x�K>y
�, ��(�b�y�U!�܋���IBx��9ݴf���uҲ�1��: �ӵi��	�5����ٴ�?�����i	�x�����\�t[2 �J^t$�׆צ4�\�D�O���K"OM��K�ni�Bcf��;�����ܧ��Ӏa�9)gG�rL6��Ƀ�a���'�Fܑ�A�b�&�p�J��.1��H�!T����t9�`��!Ƥ���ܩCo`�����\y#��O�n�H�`�'|>��y#��)pz,�g���54��+�S�OA�I��}� |�C]+v館:��'C��Cc�`b����	Dr�!��h��]٠@̦���ܟ$�����զΟ�Iʟ��	¼{RB��t��zP+ʉE�X����Ѽ7g�0htm�5�M+��I���,�p=�?	dBBy��k�hTU��Y�Pd���t��,�E�DA�%��G%,���A�J�z�wD��3d;�p!#p��d��K��i?��y��h�I���������BU�v�ܭ8`��n�2�j!"�'��S� �	H�'���=g��y@��J�����J�~6�D�O���'V��t��'_��>��1��M�����)�,<��=h�gՆu,f�����@��ǟ�Yw���'��I��c�� qu�%nQb�*�#�����@p� ��[8m�N����:X�ܘp��$Eql��2�+�-D�\l�m�U��#��(D�>��eM�[�
��f�S*o�43'��%m���O�$3GMQ=@���Z0bͩz��!ue��a��&-�O��J�GD>m~�+�I<F(p��'�1O�tC��E�ny�'ֻn@�E[��|��iӂ�O���f�Ӧ1�'�� �RHؖ.c�aR�a�@D��#�����O��d>][UC�w�ɱ��\	���n��fR��[4J�D���S�\�%�V����3e�♻VB���,	��H.������K�^��� G�< ��ӎ��c�Z�� i��B}qO�|�t�'��6�[iy���p�Ό9vm���L1��,�9���0>QG,�%[k�LSQ�@"XQ�5��Ly��'9*6-�8�(����@M�d���#M+:S��n�ay���6y�7��Ox�Ĥ|��N�?��sD0@t��U�Dc�ӓ�?1��H׶�F�Y8A�zu`��q*�N�?��O�F!jp,ۻm�8Y��'�:h��A�O����e��5�Ъ�5hR��$�<+F&�)-Y����iŏ~,�<�u��0x�Ў@|"�	�Ka~���O��}��'��[�:Ui���o�X�'������̺(<A�f��1����O��Gz��V+n���*���}� *CXqh7M�Ot���O����!��V�f���O��$�O���	2`V}��'C�m�LHÁD(:� � �ݎ:0 ��ɉ;&j��ce�|�����Oh����2�J:�8� ϯ8z�r:S��А���8 ���`�|BE/^�(�̻\�0!b�ҔW��)q���na��Mc4P�,��?a�����|�ĝ�mZpX�+ !I��lsƨN����)������m���"���/�x2����0�	��M��i�ɧ�d�O�	�P#����\
��1P�2�� g���ԟP�I�x�XwK��'t�f�� RE�A{�^ػ!��'
8PIeK9EK֔e�B2�c�.��,��� .E�d�ϟ"���b�� '.(a2Q�a����J0N���Ӣ��+��/qO�����M3d �'	L=Q����i5��'Ob�D+�'|N�!��C���y�WF�_5�Ȅ�	O�Ƃ����y(��6fq�$��ٴ�?�*O����X���'�Ĉ7��M� �PG��u\T��'s2d�vx�'��	]�w*X@afA �V$���� �J�y�7@^!G�İ!�.N\�yb�Kw6���dY!J|N|����;�xC��6qx	ATc̫vhN��0�@hP�h�6,�tA ��J;�ҒO��'��6AVy��=��(�n��-5���9���0>�'J���b�3�8�oJh��hO�ɋʟ�#5�WbD�F�ҝ�SC�OZ�(l�����?������;3L�D�:^��Ts��X��b��i����O�A��L5�<����"h����	K��?]�-�c>d��S��k� x��'#?iS!L�8�4��׃;�b�;��(z����� wi*���':~j��BlJ�3@����UD���'`����?E��:OTԳ$@͡8Z\d�cΓ^�<`�"O��T���y��U;FW+$e���	��h����)�V}��K�����L��r���D�O���O5q����N�D�OB�D�O��ݓQ�~�Qe]�
P�!$��|�V��O�/<
��	�,6�����8�Q�/0}@@���A�hT�����v`R�H�y��8�I<�J����3
���Oq�4�2)�;�y׏�7�*d����2A�<���B��?��O�x2�'?��ɛ+�R]QT�X��8�b�G=J�H�ȓ,����.`�P��'�7��e�Iß���4���ĸ<�`�!lS��O=�@뗭��r��A��?���?I��Z���?�O�����-*��Ar�E�;�|=����>�$Y�1�u<��Ƞ�'џ��'N
�/���U�N�}X��������L�5rd�Ȼ��՟���������� g�	"�TZ�ζ|���fF� )-���O���-��O8 �V
_)b�y�G�_����'t1O�m�f�"gV��[`iR�4�N$�|��m��D�<E��<,��ן )d˔�P-K��֔q]�䩖e�؟H��-�d}�	ݟ̧9~���QJR�B}h�Ucpܦ�	U�N�L��<ɕL�j�q��&b{*���%�Ӣ�ń�S�b�R$,���� �K?����K	�|:�	:�f�&qpA��עZӔj4{�	#[�������+O���vw�Z��՛F��t�|��'U�!��(ob l:c�<L���C��i>]x��2".%sg�NK��BU#���l ��fy���46M�O����|Ҁ��?!fMK7}�B�	���2N����3��<���H� ��G��
%n����F?d��U8�+�*t��˟�i�RS�	��`ؑiʿjx\*���l�s�ߔH�. 5�Y/{vn��e&P;Z�逴�7z̬���]� �x�˘	a<��5�L�>�d��`��;��S�O1�\��cɦyN؁��C�BE���'u�� e ��!�f,�$��8.�P:����O��Gzj�<�<�W���:��-���,����?��7
|�V�?A���?����y�	���@9����{��!qnB�#ώe�2Ɂ�wtR	���(�¤:+����ގ)<���G��'q�L�*"��	d�=ّ�M�4yR��
�"?l��#�N7P�˓0��̐�/�*.�6���J˺T��A۴q���'�p��"�'�1�����<(�l�L�:$��Ȟ7+:Xu�	ǟؔ'����>�R8t���KA��R�Մsy�ce�Z-lZr��?��Sny� B�P�6,j5��h������m�a���âU*��'���'�4֝ɟD�	���'�:Q[&J�9[��}�%�N�d볥\.W�a}�w�>��D�D�$ �0��/"#�	����zB�0qE��<��8���26����ˀ( VMb�&ڣyy#Ј�O l��M�����d�O��,���a��5�5��eZ�T�C䉢-���ȡA�5m<Jh0Ԥ�0$˰�O�%l��M�.OP�c�
¦U��џ ��G�:���xCl�#�і������^�i�I՟�ϧ�pm�F���Р�Ğ&�?���X.ZϼmRW �!٬�����q���J^�5�r�ȷa6t���1*�#j/X��g�#�xS�dрF�l���ˣLν�������'��I�I�,s�0
�@|j�	D,"(�OL��d�PӄL��Ķ �YCC����O(���#� �� AX�kx �5�'$�I��H���䟼�	Y�D�ԡX��:�
�!祃8&g���� -1l��'N�4����{�PR� ����T>��O�ʈ)�O��Ԉ�r�5F���O���Q%@paFeU�K6��ރ(V�x��?����ś� ��MĿ$��c��9?0�����	�O��ס<��\��䐚��0EF		�!�$�%x$>XZ�aTe�f#cC�c�џl������)[����NژT�PI��M��'G��'��bv�����'�r�'���:5r�,����E�
�#�/d��(qA�:�6�Z�,V���6�3�	s��Zt�śT�.�0e�K�ZX0��ֹs�� l�8m�l�pI8���B/�v�9!cO>]B�� h�WꖙRyΘQ�h3����'��	�/f����OL�=)%iy�̓%��s}"�����	�y�J�Hdl)�@��/kD^��	�?���u���������'��ǌ�"/P4h�≄��!��W%x��,�b�'�B�'�b�h�i���PΧ|�8ɺ�L�XjnP`�a��Vm�$e[[غ�DO�w �N�6<���B�,�[H۰, r��xY���B�J�rVn�9�ν��Hph��"7���M۲�W⦱za�1��îDkT���c@�:����0"�̙���' ����A8w"p�!�,�B �Qd3[��{��O�D`��a�'M�F�!�1��'~�6�'���3B��p�O�2b��O]� ��#\o�'��7{���'b$=�5�'?r9�@����_8O�e8���*@�z�[G#w����P�67�E���R��`1`W�(O���` ݁&Xd�!A�K�i}l��F��wcb@�F�'?I����h�B ʡxw˟�M[w�e��>�B���O��;w��C��J0in�6�Z`t
!�|R�'��<��I��F>�!��,�.Щ��i>���d-�QӂF>I��\q���Iqyr���Q�7M�OJ���|
g"I"�?Ʉ�UMCLM>w+��j�HӲ�?Y�|�
TR���a�te @��W#�̊�@>MBR0c-������
�vS�[�g�d�r�{��.?iE�¡?�<Y�����H���p���BE�\�p
:��^�+�\��A���Q��1���=
�r�:���:�ƽS�N	#$����L<�C�141��2ֈ�(����H�$���?A��� E�MЇ�Q�>�i!iϵ�	lZ����䟤�th@�cj*�	����I�4�;�JY"�1�����EAH( �B��T,``o_[�	�D�[��6���0�	�~R�Ɛ0P�YҶ�O��y���,D ��_�<�rFI�/��i)����D��B���{@v���d^8o�����هs4���O>����Ɵ,�|�<��dH2>�ά(m�V7���ȋu�<�1� �W��4�jE�-y��"��Jy"k ��|"M>�Ģ�K`��E���]�y��%���Sj���?9��?��la�n�O�$f>Y�D�׏>��d��#M>�0�#���hX�#��,lL�3L�����@ȏ	�Q���NL . �J%���z��̈m���rFA 0��%�%Κ�\�yN�6g@¸q��Č����f&��D�\AW���g�NI���'�\���ҍ�ʩX��LP�{�k��E!�D� �����m\
7�<� �_�0��'�
7m4�$�+7��O�BM�8C����1E
8Lpu�gҗ"��'��%��'p�7�niabo�)*.��KRA�Z6�Y�1䑡�N�#&(�c� �(��6��hO�l�4�
{:1R`y;4�x�oڠv�JmR��� $	f$A��U&/N~�kGM�&3T��d��Ov�d/?tJ=2�xuh�J�$O��h6��L�	H��pA	�B�bonL��%X����ԟ���fͦ9)�<����i ��2��O�ʓ��H���?�����.��dϗg4��AT�g�B�FĜ*`^��D�Od� �Wd1g���((h�G��Pժ@x��<BS��o�F-�B
58�i���B]~�`�:�p�5i�	R]ȓ+��%3���� �$m�2��'�<%��(,�.H�I2����|Yt��O��D(ڧ�y�*T7X��)��)��M�uA�<�IB-n|� "�h^*�*s�y�'JF�}����2�B���!�k��X�
��M���?��RFB���#Р�?y��?����y���k
)ڱ����Q����V|�|�S��>iunXiv�|�<�G�ݦ0�ƭ;Gf��~|
��T�KB�{ ]�\��Ğ;��c>c��{��?:�*�rs���U32�q4��O��N�f��Iӟ�E{��,k�i�0�L��pcG/k.!�D]8V�&m�fG�*`��a�獧x��D푞�񟀕'x%JT#U?!�����-U���F�ֶ^��ܙ��'Yr�'ru݁�	՟��'s��a[�1]m�TC$�M���b/G�X��ք�
*R��7oё��O���F,V�Z�� ���#kxx(rUQ�������h$��8�c
�6��	�6s�����'�S��,�6��eRL�Z�n�O2���O~��F��O�� s������Ό�bl6D��"¢ȼa���)R(HN$t��k6�$DצM�	jy��ę71���4y3��@G�p7�ȯ�	s��'����������"���Fh��	�)H�V�N���VT�`�� ơk��U�8y�d�ቐQ�I3��
w�pA����֟���燃=��dbg��^����2O��G�'�ҙ����o��v#��c�Նw�p`�o;��5�Oh��S�YH) 3��]�V�'J�����(�fn�,PN�)�r�ۘbX�|�E�Eyʟ�ʧ�?��N� JALXA��l�4�p6�G=�?�����p�����P�8�j���:M&��	�7<�Fq`��;����]�,��	�@@|e ���6�e�Q�O�l,��F�-M�x�L�Y"B���O��3��'�2��<� "�P����a�����P@��"O��O%�T�9a#W"0�$�ɟ�h����h�qp4}�!������ԡ3�Z��|Fy��9�$�Ȗ��l���J1�yB-M�?5����X-�t�Z$J��y���,���`�'z���jF�U��y"뜘^\.9PtF rytѱEoK?�y2���ؤ��Ƙ��1�n�>C��,:��3��22z�E؇�O|&˓P56��ɑ+ǈ)`�K#>h���?S�B�ɶ/2�Y�_?lTĀ�!'��B�ɺZ�~%Z "�+rl���5�@B��.&L�2��	 5�6J��TXB��4����l�r��P@�J��J�����V(5!���|�8�ɦ.�b_���J�I�!�$TKW��� ��3V���ӫ�+Fu!򤌼z�l���ƌQ��� 
V/�!�D�� ��Pq!�\=J�-�C(��x�!���lM�4l{:�a�̑d�!�D�2=H�@�I1��q��A+ў���h3�F8�zu�]�5��2	��Ǩ�u�<��h�������̓B,�Xƥt�<� e�9�H=C�!��K���xԁ\h�<!$aY: *�k�F�^��݇�m��iq��$#rD!�s�U�7
�ȓ]�\�h���PK�����M6C����6)��"<E�D��c��W�;Ŭp'oE"{"!��^B@�5�t5k�.�W<!�$�`����b�x��������!�D&��HI�nA)y��5%;!��;�(ɘ���E�X�V�M	i��Đ0#ڌ-�skA T&Rq��0��S�g�<h�b4i�"A��1#�D���nc>i�)����.��l�9�NJHAp�b���~g��Dթ����O���ʇ0��!K��X���F!N|�H[w�@M����4Y�-�$������Dܳs�(e����`�a@�b\���� x |(7�R	�.��@m �,p��F��O� p��'zR�	��< �U"��)�Hx5,O:z���I���q6Lݩ+?:i&J(tkl1`��:�$+��|J2_���f��".����gŃp�8�P �<I�x��I����S�t�[�`��'��X����d���� a��t�%�'8��FÝ)v�� $.@�N�U9%GNʈ�T�]�mٲ�+�(�	T=V��#&��y��V%F�N8�e�-��p�Q3Y�|��t�DTM�`��P>1X�
�4�����bH��<��f�T����O��$??%?��' �l�t�� O�j��`O�2���	�'��`�)�*SS�o(��qꝄ��'6�!��|��ί8�i��~?�1�)۵�?	��?)�g�J�Es���?����?��'�?a�Ƞm�6�D�p��j4OE=i�8�5ɕ�E�9��V��T�d�?�J�}rY�	�<=��K�XfIA�-�K+H�b��8���h%A�s���i�R>�kd#۞nr���$A|����R�Us:,xT����Z'�(?a�����\�It�'��$_�Oʔ�S�A��'_*�����m���Dؔvm�����4y��YR�� P(^��DP���D�'Y�It�${����*DB�IE��O�RQ��>ߤ��Iҟ�	�0��̟�I�|
�A9`��u�� ̹?˶EW`E1f�~	�w��!-LH�pj_6Cd����I(p�ub�ߣa��l��S��U���|6�d���.v�M1���>:��T��%N�' Q'�H��E�O,�!����m|X
��Q�Fj�0{G��Ob�=���@�FkNR�DF��x �l���yR�#5hpzB̈W�����Ǆ˓\����'��I�=�Z�ʬ���d|>UX�h o�����o^�j4
�ONM�V!�OV���O`!��X5N`��3OPc�,��u�Ät���j$�^�c�LAS��>ňO��9)D�hT�'�2x6��4Nڟ	�>�K5!E
W.X��J�v4�mH�ǎ�c���#/�$N�c0��'=1�Aq�/��G)�|��h�4j4��R]����I���dX�JQ!;�Tݘ!��l�OD�=�'9��=i~��k�m>M:xDE�?�Z˓{���h���?����) �GR����OVMC�1ܝ	tP�p!� �OP�h ��wGܭ@���>���J�"����)�>|8J=pfcjAT��7��&��]_8ء�I�]���C���&JQ��q&D�]A�$��M�|�uML�Jdy�3f
MzԠ"0���<!�DVϟ���O~J~R�O� \uzP�͂����&����6"O�lc%JR)~r�����(fܕzd���O�Fz�O�ڜ���Q>(�6�s�O�4Ot�y��'��'����1,��dP��'���'_���'�"�!�&�^"���Į��}�����2&H����t���ضg�3�����'zꡈ�M�z�AW��]�̨ a!���@��#��N���OF�SK�)CF�Z"#l��#$�mPu!��+Zz 2��	�@�T�x�����D{b3O\���yj��1�M�@,0���Ö2�XA �DX���g��	�c/�Ov(Fz�OKR_�,c��5��L�祏�S��B܁H�H��*�ǟx�	�\���?I��ԟ0ϧ`���yR�
�T���M�V��PC��ہ6����MOѐdC�,E/L���h6�͏hLT�rdN�M""��&T"h�Ԝ��#�*m��̻' ����ʃ#S�is�@g�I�
S��d�u�T�#F^�iK���G�G7A�r��'���O2%�1�OJ8 ���".����'0�d���
oƀ�r��?j�:�y��<���ilP�x�R(�M3���?��O�^�x5h�>g�F��"o 	�.)���)J��+��?���$�]��D��U����ɓ���� �-؎�b�� ��b�zs��	�3��M���v�'�b��bU�:PZQa�/�j��"
65�<<#R�ӛ��Hya�֔*�n�/N("��`��|�N(�?!��)�;h2@��+��{�ы�̀�r/!�$�B����O6~Vڥ��늷7��'^ў���Ĉ,X�p@���P/oMf��kԿSD�֟t��������0�O��Ӎ@��葰�Ǩ!hv|�&�4*˓a\x]�<YS�	��,�C$���)��bY� ox�?���p�	!y��W?�X����N�:��$i  [%�M���P��C�'`S��?a�'�?i�'l���`Y:�Pa�D��3A`�[_1nZʟq�Mڟ��Dȴ�������8�L���kߥa��e[c�A&���#GT��?q�26 �'}��OJ�$�&�Dߟ�ZA�0 ɠd��'���
�����"�d�O�p�J�O`u��0#�^�s��nƐ�y�T�	&)�s��l�p�eaV2�R�?���IPp)v�'�n�O~��������e���%(\�/�RH�E�K岽�I[�<�D�O^�����O���	+���sӰ����3N	Y���I����0mZ=I��m��<ဉ�Ɵx�	�1'���?����B%��d�1	p�EZߠ0
uU	~U��x�'�NtX��?�U��@��`�p����?�mڋ2;��	�| e���\�Ft�t���M��' :S��?s����Sڟ����!�r��RHN*Y�5��-A /_.���4[ej�'�)��i� 7m�D�$���B��?�N45�6D��C�=]�����	��T�v�Cx6͗��pn����4,��^?a��B*P�� !a ~��b�@���	�'/p��dB�����鎖<pf	��4�?�+O����O��d�O���O<�$Y�&
:ds����c��Y�"s�`�nϟ4�Isy�X�\���l�I�x�f��9&����V�-�'�^
�M���?����?�����4����O�͡P��r/N0◫�&�@��Hݦ���ş��I˟��	��Д'��O���kN6u�\8Ӷ"g�ȓ�S�����py�!V`7��3R�)p�N���ӯT�"?�����$�<�.�f�͘���9H�8�����*g��cybQ�x�Idy��~"s�N@�TH򅑕B�%�$��a�<��,#fh���*W4
�B H�<i��K�hZe���$y�\�i@-�x�<���O�"T���e��&h|���k�<3��.���c��I��qqWM�j�<鑍���nQX��סv�J�XT(Ph�'����v�Tm;�	I3t��!y�N�rVv1�Ղ�2�e�Y7��Ţr
X�d,�� ۳x�shR9�!t�	"F"
���-扎b� �"5��6b�H�ʃ<k��b��� � +<�1ˤ�՛Ԗ��$
��qR��F�K�O��=Y���N`���(S�Xd��PD�ؔ[��aꠅ��� ס�{�`����8�!/^�lbM���B6Dr�L�'�S>Sj�12%�
/� 4�4�t����c�f laю.q- Ԙ��$fi�@+@�雦.X$*=d�����/D�&	(Μ�P��d�Oj��b�M���Y?4�B�K���t^?�Y�d���@Z`J&G�����-�$�u�%�M�jp�Qs%	rn��ȴ}������<?�H?pTP;%CrH1��*8�D�<J��-w�2�%>�&>��0�%�
ix��\?x#V%Q��;�	�h$�������''t�LD,u0��3�ςO���ǓN�"r��O>L�Tl�q N,5f�p��Qk��
��M���?I�uu8}p1E���?)��?���5c��/fl=v�;$��fE��D
!�CcZ�[A�	J�&Q*o:��B�E=�1X:,Y;�'�=A�?�`x��͡d�4躅�V�*1X@��7
�BL�4[f�����B��0?��睳	(����H �d������9�j8۴�|�
��?�}&��0-�'� ��⪞#�$���"D��ʁjڅr�L�aI���)�+����	�HO��'��W�:�|ceQ4h����1�)H<|y���H�2A�I���ӟD����l���|�B�ɘ HBm++СJ��[tb�I"B��'� &�`/� `ײ�{���jv��_Y<� ��;ND�ɉ�#( sM�e�U�Qњ���>�p?�!��g �y�M�	�X	qτs�<1S$�=E2���-�(�8��FIG�>�Ɩ|rb�rb�'}��١��T1 HE�� Y��fH���D�O��&l�O���q>IH�N�O4Oʌq���.d�@�#�\7�(r��'젍}�hٳ#�.�� ,ޟ����O�&�<1%���pI�����I�V\u��C�a�vۢ�,D�(�v#� w�� &�%d>���I%��@�[/1�H�@cwZ)Į�)��&��vF���M���?�)��mB��vӀ�-�QɞQ�$@�D�4|X ͟��	�$ڄ��G�S�,O���	��<��Zb�2a �I��x� &�O���TcG��/XNBpsWᙏL$Pj�x�.�3�?���|��ģ�;mK�]��M��i�(I��yҩ�H�����/��]@�� �p<ia�	< ഈ�nƍ{7�Ƞsc�?i�as��?i���?97�<^)J�����?����?�8F$$ 
"B���ŁS J8ʺ�k�y"�G��<���^=9L\L �2I,1���y�(*Tp��I�ME�d��
%�hh�@�[�E�`�|����?�}&�4��� I�����1M�BIr$*#D���1N�N�p���u�V�sAN6}�� ��|RO<�' 
��Hͣ�ӚA��X6���}���æ�H���' ��'��D�'�4��uڑ�_�Fl�P��U���z1�ϋ+�!�$�6|ᔱ���ӡ}p9�+Q�Nֺ�TO���t%X؎P{v��r��yQ�킽IQ�*�O�p��ħkT��9vOьG�M�r"OVUs�¾Tf�)��!t3‚a�d�Ŧ�&�Pkd�Cݟ�������FϓV�409�˃	�<Q6)]��?���}v�}���?��O����`$�(G���3p��%��ki�4�g� ,O�\�f��ܵ1��Iz����)0�L�g�I�g!ay��M1�?���>��g���~ ��B�]4�-�1M�<�!�)�%C��	�~`B�	9$�t�Aj��'R`����3!{�M ���;rI6�'�c3l��������<�OZ��i�\p;〓s�����N�r�(	���O���ɿ5"��(�|�'�>��#�z'x�A*h5t� J<� Y]���OZ���(RU2F�V�L�H<�`d�@H>�~�֠Zȁ�T�l�|(v�MB�<Q�IԔfN6@ك�c8������<}�^��34��M��\�`I����4�?���?qS��3:�j��?���?��'=�a e�X�k�DDr@DՖv�&|ڋy2�؍İ<��$�4R�͓�AǙ�\�A��}�4�@�剤���y�&�. ��̓'Oߢ[��I�%�|R�ߢ�?�}&�,*�Zw�6WI� �zزvC��y��J6�� ��2eC �x1�	����HO�) ��Gw�b�m��Y��X��/��F���#�!L2$���I� �����j]w���'��iP�$�0��!&�"uu��̔4)�+O�tx cX18@�@*�Z��pRt��1V!��X0�8���S�V6z1 ��\�ȣ��'��D�8� �X�m�?�@����ʨf�!�X� X��(�KZ;:Q,����u�qO|�o�M�I�M���	ϟ�n�2'���!�[Ur��S��G׌,{���?Y��H��?)������
��?�K<a�b[�FZM����g�^ H�HOX����-��}�X'jܷ7X^����ݼ�V��Թoi2�%}�b�$�>h ;=�8�坨�yb�S�<H<B</�� F�B�Px2F[N�,�'Aġ��.-�F�ട|2��,�D6-�O$�D�|*��X&�Mk�Ia�5�g��koN�*We�V�"�'��е�'T1O�3?��K9�9��*Ɉ��(�+񤝉's�b?��f�N9IE��{�� �#�dV�!���'��	9L��p��d��"����g&�01	�'����I�<p�A�d:�9*	Ǔ*�Q�H�ĜM"r�@N�+�u0�!� S��'�R�'����%[6;�B�'7����D�Ö �,u a��`���B�U���<)��|X���ËO?}B�  C��!=��Ea?�I�uK���� �|�e��@B�
���40�QS�Ʌ��74�I�)�3��(W�4Ag���*聡�ӵW!�P�p0Вh��䙒�\'7B�v��i�ɩrn�U�-�&,e
���aB"d߬��s��5_�x����?I��?���d�O��,@K�Oh���̺7-v%�(&�0kB/ԽI�M���G*Y"-��C�	�K�����F �zULĻ#,�)<B��ш�O-��ɏ��t�㏓�Rzr� w+��5�B�ɕ5�,) ���m>@@�&�SC��\��4��%�d�Y�i�r�ik����`�?w��[��=iGj� ���O����
�(���O�����2�d�z��ԛ$咶k�Õa	U�ayB��>��'��%����;Ī9�M��u��LC�t�M�����6h������:�!�/@�fU�B�
I�����B=f�.Xň"6�B�I� 0@��d��A���/B��q0�AB���,Hyش�?�����	�1n	6��=6���D+�>l������Z
 H���������Ɵ��<����O'
F�����e�t<"�D�.�'��YY�����U7�Щ7��/��(B�ػ}�'%n�a��3ɧ�ODP�3q��>��i�U�d&���'0���F��-.*�d�ƚp��B�5IQ���c��%j�X�"�*=i���o�:���'�"�'�Ҭ��E>I���'�����{sGPQ� L�q�F�j���T�Ӟ7v1O��'���F/�_&ȡ;E�{��e��} S�ٰ<i3��5n��%8�ID(EA�@��6kړO�P�����ēg
�t���Z��i:vgS@H�p��f��	��Y%:�!�_pD�O��Dz�O��'c�e�W��&I�H!4��9��a4���'9MiC��Ox���OZ����+��?)�O�@\�7@/a���a�-N�¼ۃ)Ϟ�xB��Of����)Z|�1��ʲV���'	nEQ��)�h��!!V�7/<�w�@�?ٶ�'�~�GU�70VV�;T��r�]@�<��&�#1O����Ɂ&Pj��wIzܓJ��f�|��ؖg�(7��O�6��<A$[Ӭ�Mzr��we
1\M�I����R��ꟈ���|b!*ײ)�8�tgБ>]�u��Y5=��#b$a֨��N�~.t�LM��<i""=a�謸�LBNB�I��,;v���m����H�a���h�
$�'�΢<1s��h!I��+�m��lx� ��@8`|:�B4D�ؙ�lЅf���N��I��qI-�0�1��Y�D��ч��)�V��@�nH�%�i1aB&n���O�'�܈P�4rH��Q��`��Mc�	ܪ˺�!W�'��),?��Pj�X*ZdPJZ��'����S�l���e�4\$̹R��E($]���`fJ1p�ϲs��Y����Y�HTr�'T�@;R��G�P�-V&�uf��a�b]�� �<��O�ɺ2�'62�Ӧ���*KJ!�ڗ���8}�4�	;��x�a�<<�w̚���y�CH�p<	��I�Dg1sG��)y����4�|Jq�l�����O��D��C1*�b�L�OD��O���w�<��w�>0P�v�z����^�i��<r�����%JR�y��i<}RBӥlV�D;ǧ�j[�j��i�(P/^>*L%�R���:t9�U� �ȵ�qC�|��4���ݯu��q`@�R����M�b����D[( %�O�D�e��!��'Bd���*�)�s!���p�wFI�Z��fBx�am���SݟH�'��%R�状E���0� ��$��q�b�W.;� X$�OJ���O^����#��?�On~<�!�ظ7ބKE&�-�R}�5�H�+�R�K$c�iPpk�
j�џ�R����Jr2|��^0(Y�h���B &�V��I�l��HP�&��|R����$�>V�A��b��?ä�Yu�{r%���?)��?����I\�&i���P�wF�����m�!��4>�@��; q�$	E�N�qOF�m���'8��@�m�4�cӂ�`�H٤	`v�+v�ȿU�� "W-Xß�I���������'*���I}�#^HP�*0�C�*|�i�*۷g�l��
�*1�O"���m��-�	���b���sR�'\�	�D���2-8�e�U���#/Z㦨��je��ct�)���#]�X�i��M�ʉ�V�����"��[�O�-�������:��)[�i�B�'��S;K�io�DR������Ia�YZC�Y"�x���?d����r%P!���q5*�*A�AzY��Oԙ��IȾ(�RY��̊]L�k��D>�'��(+s�ؚ0�<ؘD�U�YV(����x�V�����<a�p�g`�!ƾP�4���vO�m�F�'�L�O��� �0p�ŦGp��`�eK1K^�"O�����B41���԰lT�A�"-R���4G/ʓԱ��ѣt�x(Ճ�%]��Apa}�J��O���U8L䍘D��O����O|��w&ԱE]�/;2P
�A�%�l����{>囱AI�5�|Pb���Kv$�'�������a�Iy���/�@�����L�1�&餧��`�*�F�#W�Π��H�y}><���%Ht�\߼��ť�: �6L2
�lݛ#�ϝ.�v�Ob͛C����ē/ �a``�b�z�L�k��܈B�8D��b0��`���T�H!�X�!��5}�F+��|J<!�	@@;|� ���m��8��d�%b�X8�PR"�'b2�'2�4�'�"0�����ɍM.Z,��&"#Z �aEV�b���d�
"�f�#ㆉ.V��?�r@2�	BT��%2+�M���O=[\M�a�[�G�`�Cpd�'d<�#޴PIL�j��P�'�
��/*^!��؅
c⡳%�O4�$;���'.dIg�4����5n�=a�J{�<�ШU9�|0s�U�V|H515g�`ܓA[�&�'��65��)ڪ�h7MH)V��u�A�ĆX&��/Wф0�Iß�Z��Q՟��	�|R� �3r6X��`V6a�ĄjvI��/+��Z4�����u��m��h��d]�8{���g?nE[1�IfIr�`	�\b�s$�nBl�j�di�h쀢��B�qOxL��?��O�M*Uĕ�d}���t�(ab�v��/lOC�M@�n$b���gȰmS�A8u
Op��V���v���zT,�:��kR"H�A�����<!"�	�?ͧ�?�*��뇊z���1��?L4r E��"%\�{�m�؟p�IX?�-P��Q��z]P�Y�|Z�E�����'���r���L�V9RK��*�6'��a1�[!Lu0�)���i�|���_ֺ;�ɞ�Azn��7'�4@0`DY�����$
�bO ���?э�ie�v� �bc���1��(�,�cd"O\$��B��9�U��%�*�4�؁�'=�<���a�脛�HW�daJQ� ��Z6��'���'<�Ԋ5HF�g�b�'��sQJ�_�^Q9��F8�v8�%L0˘}�n�#w�<*2.Cf�rA�i-}�_�8`����&��`�d9��]�d?$��b�J�={�I�<�;�&��'�M;$�t޽"�+�/�D]�ԌQ��V0���+�?A�O����|ʊ���y��c�-g�!�K!�ː8����ȟ�,D�ʐ� 8 �������t�'�����/M�MRU���
'Mz�2k݊B���)G!�O��D�O���P���O���u���r��+YFd1�G�'h"]�������JE;��� Ry�'�����D��DE�u�C"5<��gf �S��	fK�I@���V-֒lB 	��{b	�~C��y�P�������=,���I��`F{��$Z��("��9K�l�a��$K!�䂠\V�e!aɀa�`�Q��TXXqO�lܟp�'�t�u��~��4j�\db��Y�YG�"��V�*!y��'��/�T��'��ɓ�c���JDNZ�	D�ɡ��ɽ's�h;rJ�ZO°*u'	e`\�q1''� ���p ��OU���,�|ȧ�c¼@Q1�� ���ˀ�M�SKXK"�=��O|�ķ>���R&�tT�`O"5��݃�A��=	G-Yp��ų2��/��5h���b(<Ya#��tBT�U(��(X��1�@&X�ֈB�����&s�r�4�6�$�|bP�«�M���_��ʔ��I���]�ƍ����'�TСW�Aؙ�HR��,���~R��z雒%�=wr��@�f#�����x�����`�t+þG?jȧ!�cB�Ư�Z��O�8����  �
t�R�R���ibN<�0�O���2�'�Mc�O�,�|0��ж]�<(x��MW�<Ys�*�܀�dG�^t�B��V8�@�����(r;�q�t�Y�]=���$J������Iן4�I�b��oE�5��ٟX�Iğ�N�$i�&x9��U�$1u�h��T񣵭ʊ57�C��\�K﮼�BL�ḑ��v�⁠�ǌ/L��Ш�*b�)�/��0��L��BÐ��y��V�L�M���7�M��y��m����eH�C|�{���P��D#?���O�i1ғ pz`I�.+�5�5�	R栆�#�&�ˆ���#�i���{P���O�}Dz�O��T��SB����* ��tVqH1㑼n�|Q����?���?i��"���?�O�B�b���J@��SjS�M.��e/��Re��g��_��E�v'OZ�џ� CL_?>�r��E�N�I��+`JJ��@Mu�d��f��5Ǥ�m�$INY)�I6�I����y��>q|�$ �,�f�#�'v��	J�C�ԑ"���J��A���%HU�ȓ&�ʅ"(_�!5fLc�')w`�8�=	�ia�]�đ�$"�����X�UiБ]�Q���>Q���y�ʍ�\�I5ǂ��	۟xϧu~����*!b�Hd ��$m�<}K��I:�f�#��5L�����߷��O�;�J���eJ���o�t�Q�EK9$��!��]28�Q�^�\P6��� 4Zp�$�P?q�����E�Jj�m�k�����!I�M�qO���� �Ap��I�A:Y�G���1�
O�E��솀mڥɤ�ζ
ۊ�" )�0�l�d�<��fZ'�?�'�?�)�A�0�dӆ��F�G��z`f�މc��t9�d�ڟ$�	�I� 9AE/ˌ0o
|���.�� �����'�Vt��Q�t�sdW�!�`&�����ǵGcF���ԑ8]���b��#�,\`�u��"X�~��j�1:������Oz\��?1���vӪxY�l�% TD���N�,Mص��"O�u�%*�'j1FP@R @3M���G�'aV�<	#L�d�专BT�>�x���� �B�'2�'k��	��b�r�'�������a����܀FA���Ix!�֝v���%��xYv��.T�-��e���i:}R�PW	��G�6Zr��j0�Q�?��}p�A*M����6�#1�(�`nz�'�M3g'b�Iؒ��.`v�,k3��>9À��G���?��O���|:��� ����E����Ƶ(0�@"O��*ߥ~��a	¦V�xz2݋��>9��i>��Iz}r��'*:���m@ ay*����y'隖Ŗ7�&���O����O(�I�O\��w>���Q?Q����y�ꩋf�U0m��`"�y��)�t
ע_wX�F���.��]c��'�qȵj��R z=�A)�<�J���z�m)%�iM��� �5��'��9Bh�=����F �^H�j�Ǳ����R�'M�OPx�KA�u�K��̻Iڔ9�"O�q9�̒��&0�@�[Ҭ�C��d
Ҧ���Py�'�A�6��O�6�Ѫ/F\�E�E�Ym�P�����ȟ�#���	�|"�"H(=��i���5��Q�qb����{Å�^}�p��;?�DX��	����� �J"&�Ti��"�	g=�@�ऑ4^`R�Rq��iP@U;���>N�I�V Q6/vؕ$�T�V��O�ؤOl�J�ES���="񄑵=o^�� "O �d�A��<;�#�9���@Q�IO�����DoBԩ�H� tp1 G��z�,�J�|"*�.6��Ol��|�����Mc�C��'n0!j2��ypd��T64��'����$ǽQ�u�؛k�ˡ,��yb�ػ�S?٘�cӶQ���b���6�!��-�$2uv��2���kelX�G92%cRF��)�1a�e+U�^�~����Hk�'���H��ɧ�OҰb���tP�:�Y�0w�=��'K:�C�I�W��d��-A#���3Ǔb�Q�$s���~r5A�Ɣ-1v�"&�= ̛v�'0��'>�J&� ��"�'�v�ٖ6�P5��'@Z@��Pe�qT���nL8j���7�99E�keW>�ͧ3��Ę�h�O0l��N��9�` �'^�+����_� �� �H�6
!�n�4.���>Ap��T�y���
�(@p�aI(5�D�2���3dhL�$���o�Oq��'�,�`�e���(Y@S�ek6��'	��bDO� �`�P�±Ŷt�M�<���4�.O�A˶�ـ]|�<Y�@�	f��bWZ�?tUHÇ�ПH����t�I"�u��'"8�X왆����E���� y(I��ӱPw&1���S,G`����dB��?��Ǚ �� ( �r�d���E�E�� h�˛1rXј�MR-�0��D�(Y7��F�;a9��
�n�C䩓,�?a��?����ۣ.z8y,B�M�NX ��s$!�pҨ�%#�&�������LqOv�o��'����~ٴV�H��S)M��QF��j궩h5�'0��fHr�'3���}`g"�@�Xi4� ��ĄP5�Ή;ܶ{��TR��!�D
̺��L�����N�0S^���U!�x�mR�{�"��l��OX��S�'u�S��Zh��PQ\��d�@]HI)��8�	���k:���	�<�бv!�$�`�3u�Ϛ5I�R�
��9�H�f�O��oB��7�?��_�d.�=3�����(W��`� Y 0��˹=zp���O��"��V�d���کw�T��WN��U?�qOZ0xˆ-�&ľ�~ᣲ�.�$ҐDv
Mö�A�+_ �
�T��\��ė�$GC�dy�\�EOR�NU��j)��7����ҟHG���i�dIE+�����$h��~��4�e )$�B�M߅PFj�kb�Ҿc�D��)O��Fy���+z��T[#�T>LRxXJԯ��n��l�џ����D�2c�32���p�I���.\"�p�!�eC9^��]�tA�aׂ�a
΁R0�,�vIP�\��XE�U�'nx<�+�O����cd� 5֐�IԎ��P��aۗ��n�P�f �Wz�m����<G�j7e<�iB�f���λm� �6�6.�$-YŤ���<��H/�D�����L<�C�U�4�E��*ܐd0α�X�<Y#�M-o�d��b��V��i�E�V�$o���d�x���Yv�<*SKS�ef���`�@(,J& ��1M�6���O��d�O�<�;�?y����dd	�s��Z�#�/'�y���@
t�!�'G�=bY��W�I\ؤDh�AZeFy�E�)k� 2��X�0�BX�FU^�-S  ��k�a 0I���Ʃ�2?k�Fy�f�mh2� �[rtL���ٮVrz�8��O����&A��l#O�Y�B�k#J%1iC�)� |hC��Q�:2R���;mp���� ɦ�%����b�4�M[��MR��.��$cOM<A#�iY��� �b�'�98��'u�'� �1��cV7B(\��,юBY�4�ӧ��>����Q8��<b��� S��S�!غJif�J�Q�Y@�$��eь;rh�X�=��m�&��>1Z���@)�	�-�����զE�ܴ�Mf��0�$�A�>-�ƹ�ӂ�a��Iџ��Iy����	ʟtnZ5ܥ�ެ+�0Aqf@��s�TݹSO�m��m�T������?9�j_'x��J��U\��;g�ܸ���y��򤓘$��Dn�ҟH�	�����%@��mڗ=[�X	���� ��a�Ǽ3�}���?���m��lz�L�;?��x�i�Y�����+^���f1\�� Te��ēEڶ�8ӎF2����ɫ`U\#��
8�L\(qM��hAPl�U�h�j����sQ�(j`�x�$I��?���i����<�ɴ��k.2�a�"����9&��O��O����O��v�]Z%@�wDؘP�ա�t��I��?Y�4��XY|�����w�!0�OT x�02T�gӔ���O����,4�.�3�o�On���O��dm���dƂ �H	��"�1bIb<:˞�x l�(�
�)PC��"���+�������˸���I18�Z�iF)È?� ��	pv:����AT��i���_J(����jܧz���6���S�T�:�*Y��P�z�c�&����~��)�3�ğ�Pϼ�31h_"q�>���D!��2c�l�6旫�F$	�U��(ґ��R�IlI�mk�iF�h�<�v�G1���X�GݢW����?Y���?����O��B0�,��̭wJ~��A@�0��&�0� �,^�h(C!�Cm� ��É�|�C�I-\�fY�Tf���t��	0;f���Of��ɨ+H~���_�sz=pp�@/�B�	<Y��4���I�vP�H�Ē AR�X�ݴ���F�h\&���㦕���(r"�šb�θ5^T��BfM�?��T���?��Oe(u`���ē�hD�ec҆�.u``^�>݄�	5:G�c�t��NJ��@����0yM^�Q�#,O�����'z��'0�(�6���F<��kO5XF؅i�'�������Zez��E�<�j���'�|�fȅ!Q�]��\��<�ɖ�Z�jw�'zܘ�6�z���D�O ʧ:<@��4n��I�L���7��t�!c�ٟ$��^<����)u����R"x�����*&%�O��r�HW�t`��Oۅ8�VXI<��㒯�;��Sjβ������u�ʏ�u�%��o�����Z^�5�1�WgPl���x��,�?��|��D�M�1L,�H$G�#)\ �/��|��'�����!�/n����'L:&:dZ�(��|r�If�t�0�[�yyX�GI�d�,�p�i��'�2!j�6�'���'��;����T"W�SbFd�f�-l�`@mT1gJ��8$�ɊW�n�"D�1���'�ƠKqAH�4Ҝ��V�Z �vQ	t���CZ�: �S�Wj�QNחv���b�i�$d#j8���%ŉ\,1���F�lY�4͇柼�'(غ��|�����'�,��aD֨�}���B'"̌�'�~�r���Z��=f�W�����'R>��|����͉u'���A��<T(��l���Є�	5�q��� �I̟��^w�2�'!2�����$`��* ��\�Ƌ\%t�I�"I�936||+�j"|Oh̀JΈ���gI��y"	�%�L���!j���D�^�Լ �G7:^�{3F���TA�%\���J<����?9H>a�4<��Xd��:�.�Sd�_���'s�㝄:9��'3�R?����x"� ">��s�@r���P82ʓ�?餻i��P�6K�A��q���M�EE 
*~�����i���� �^v��'4x�f�'�b1��%�_T*�ö���F��(�C,�Bc��e���Gd��!!J��
�`�@ݞe��Ey���udl��B'�/"��I$fQJ���
��?7f�ZGn�A�4��7��:>E�s�2B��'6E����b�8pᦍ�	?��4�	�u`��ȓ\�@�h�,XR�F�ba�f�Fyr�i>a���N)��!��u1f�2�TA�0�%����V��M���?�+�Zj��n��i!�8$T"�'G�+w�x���ҟ�	�9���`���Ry�D�O
˧���Ǿm�z튇%�PvQ:��,ى'�.��'D�q'&�X1z��P���O�R�"+�VG��Ip��>��I<Q��N�8ܴ(U���'ޱ�l](sfU;h5r��w�X�x�aR��$�OT�($�,A�ᗝ����"�1Z�����/O�	o��M�M<itF��ܥqp���Qƍ�M
�aQv6��OX�D�O��hּ*��O����O�֘7T�j���7a���E�@?���#�A�=ltҜ�A@��gV`q�N���O3��� �����#抃<�  deE6oCj���$1� a��8h3��B��4%0)
#a���-80��w�\��D*o�*	�5�ԓ��A�˔K�	�����xҤ� �J�:V�"�E��4�y2�T���.nr<�f�ő0RM��?�g�i>�$�� ��Ś=~Ε�d�q-�c�D�d1�Hɟ�����<�	��u��''b8����X�'��h3A��5%h6�`k\�m`\�
��>:���Ѡ^�5���F�ص�(O �
�Ɨ�p_P]EĜ�j�2�Y���F{��{��0LN�7��=�&܃��/D�`8�/c�I.F"�Xx1.��F�ԪN�)�Xer ��O�e��Ia�.A��ˇ���0J ��#L�H��$ �DΔQK @��kA0 E*4i�'Z#NqOdIlc�	� D(Ț��?mcO�M�TȀ��H���!,}�'=�Ik�OI��(�����6"�-Aє�K<��`��e��>��*f�ƚ;p���6���� /J�r��O�~$ԥ�ȓ b^���͹&fX�W@[�?�`�ȓg����rjH�=T<z��� _CL�����qs��(�n�QL��9�Bi�ȓ=����L�T ��q�O�Ѐ�ȓK6��q���xͨ��d���8�ȓ~��=�dF�����R��]lЇ�O�(ݨ���Pp�(��Z�c��ȓ�P�!K��*H�����ݛ�Fe�ȓ'�l��IB�;�h�(�>V���ȓ]���j�a�"���ǖ5+�t���{b���C�.@5@7�'h��%��wRH{���z���+�I\�G����A��ar�˪bd|e��"[&r�:��ȓ!A4�b���7+޸�bL�>�Ҭ��,�4�
���'?�f�`SIx�@�ȓu�,L�"/_�l� MaQfס#&Ї�Oy�|R�P�Ott��HG�}��d=�(�B�	)*545���LSX���P��]��)��l͈U6��Πu-\�I�7�(�X�8�E�f�<1��ϴK|�x�B٘#��0�׬�b�<��J��n����͓_��l���M_�<�s�0Z&yk�A_�����(�Y�<w\;�$�#!�)Y�ni��n�L�<@�߿��$(��>'�h��bI�<�t慠b�Rqz&I�� eV����OF�<�e��*CJฐˆ0E����!�B�<	� �4{�@�����+M�RĈ&�A�<���zy����dQ���%z��z�<�o'������.TϪ�����r�<��.I�~r��ql�)vQ "D o�<��\&w�iKq�Ռv2܁:�_l�<IA�^�rƪ��PFP�m_2؈��@�<9��%?W��p+�\�����p�<Q�ޗl�.,f�hRIFo�<�V�B������� ����a�<�L�>K �jWeˤ'�`a���[�<A��='�8���$mn୫�K�r�<y$�Z(�X��W�KaH:��gB�n�<�"n�W����o@�q�(�0�Hq�<F�6|���a"�;31���x�<�@�&Wo�}�!U�+C��ʗ.Bq�<!�cW�h�r�-�-�l!JPih�<9G�:26��sIC�u����d�<��f�:ک�W�%LT �9�.�K�<���[�:����R�НI���i���p�<Q��J;R/|�PL�H)J1�ao�<�j\#(���kS��� q��c�<��. ��^D E��_���(Ё�_�<�Fo${K�ŀ6"S� �{'_]�<I�ԍB,�T���n����CX�<I�Ǜ�q�1�Q�Nf�X��w�Q�<"�&��Q��$Ű���yR@�1I����
֛l��������y
� h�i�*ԡM6��ږA@���"Oz�)@D�(�*����l81g"O��T/>w�	����bI��S�"Ou�@h͊�ܑ���*1R- e"OHe�`��AH�{��>����"O1DJ��(Ze0"]?��xa"Ox����ڔc�h�B$��wrұ�"O�����*��c$J�/�R�;�"O��ӵ���z�J��X�k�Z ɥ"Od�����+��Ӏ�T�2}`5"O�A2�%��Eɶ8�1���x�Py0�"O����aɮ(�
 C�A�����"O�� ����h#��'�⡑�"O ���B�/B����
�8u"O$�EGU;@q�MC���s��st"O|�����ȹ�E�9rڬ��"O�)�L[#L�K��D�=\��`�"O.���Z%Q�ҝ�A��U����"O4�3��I��&���Eÿ192�KV"O�iÃA�?R� �ŮDz<.��&"O]���B��a[����R"F���"On�s2��$�j� %�Ťo\X"Oҭ���N�Z�R0Pk�E��r�"O�|�F�'v�p!0jP9|O��Q�"O��ᢢ4${~��r�	L����"O"�yVb��fӆ�vD��\#pa("O����W�X�#D�,�=�@"O�8�#�/M��PB���'\��=��"Op����6)?��p"ٻ���P0"OR�1��/e�Qk�f[2[��� G"O�����+��XB�ғ<�N<��"O��[q�U�m������8�Dq�!"O��3bQ�
�1�5�]1@� \��"O��Q,ǹX3zA2�T�E�g"O�MJ�n�Y���Y�C� բ8�"O@�0ˌD�.��[�ڸ+�"OTL3fJ�(� � &J�|�Т"O���`#�U�RlY#΁�w�PK�"O��S��2V��� ��MTN�S"O����+Y$Q
�;`�4��у"O@ܒ$�#w,>36��Z��
�"OАⱤßx� �jd����"Oʱ"T@�Q�� j��Ȯ�<��Q"O�H�%{딹�a��!R���"Ol�Y�+эw� ʶ�>4�"%b�"O�I�b�5�B8�E)D�6U�26"O*��S��Cx��r��9"앓�"Ob��a�B8����T�09�����"O���f�o]h�	�M�7� #"O(zvwMN B�+2״m0"O�|+�K#�ʉQW�	z���"O���Q�X�G��1DK*�����"O��Ć-;����0N�LW�#"OH)��(O�ư�7�Җ/K�� 3"O��Z�n]��V����e�eɓ"O>x��
6a243*E9yS 9��"OV�z3nL�i. ��
��5�H�а"O��[3��m�40�����dP�"O`�`�ӧh�1��.#����"O���,�=UXy����Y��9�"O8U����:g�5I3C��*�𠢴"O�DCŌ̶c�ĸʦB	N��C�"O�9p���.єx; Aÿe��"OL<;H^�K(��/9a��2��y
� &}c+�:)6���x5 ��U"O �s�ߟ@���Ȏ6�5*2"O�b�o�~�> a	�=(~�D"O�Ⱥ��@	�Pq
��ys��x"O8}���B���M�S�[=-d.�"O�������x��E�;=�"��"On|��ӱ�D%�$�X�W�-q�"Oj�;�W�}�b�1�������7"O���g?�1³�77��d�"Oč����;_��5�ӥ �d ��"OrA!kQ.����3�U��i�U"OT�p���1zBl�F�U�r��\��"O�����R�1��:Ul�
f
fU#6"O�, ��b��%R���%��B�"Ot,�,�T�H������5X�"O�T!��� \�����j��q�"O�|y�hΦkbU��*Hg"���"O� �v놓��<���&�Z)x`"O��;.�#h�y��Д*��- �"O�59f�U30�rWF�^�p$"O��qJ@(����D�%��"On({���,;��	�#� �I#�"O�9c���VztPB�����A"Oiv�h�P	��ͲB�I��"ON4Qs�A3i�|l܃=I����4D�,H���qh�p�D�(%���1fM(D�����ԏf��h�5��;*ct�8��!D��@�MZ(f�8��� \6#�<+DN-D���6�]�Sve*!!�]�h<Q�>D����K�,3` ��b(ѩ1K�xv,=D�Hh��Dtex\;bdN�S^H���;D� k� 4�x {u��<�� @6D���2F! Q�d��i���,Yd8D�<�!4
�r�C���)��C5D�|p�$�;6~& �2�
da�$`(D���.@@-�c٫"B����'D�����\�kE��Q����0D�*�@�=C?� ��X(cV���)D��� �[���Չa��F�� ��<D�4"�nݹYnʵ�rh��A��hH��:D�h�%����FNµN����pO=D� :�#�1X��%S����5��C9D�8Е��<V�F��G�V, ��A�,3D� �d �o�|��D��F�e�'d/D��
d�Q<�"Lk�.Ѧ^L\�3 �.D�8�C<�@RS�N�>�<�j�I)D��Bw�R69��caJ+	�Uya&D����)\�%�}���I[��X�eH#D���֌�&h8"iL&�@Z�4D��᱇�� �g)��a0+2D�`j���)\�!@��C��HY�`/D���g���eЮ6F�]�gC/D��H��L2dn�ђ�A�Y˖K-D����N�!'���a,V��5�f7D�\*u�B�|{6=����-���3��?D��{0�U�QL�8���v�D�6
0D�Af�R�%�0<�.
)a�$�:D�̘�.����i�K��q?�ġRa<D��i�#h��`Ó��+v�J�S�E&D�@��� -a���'㐹/Ak��!D��BdGL�dy)PGB�:���FM%D�<��G׸�ny8�	�;E�8�h��7D��:'`��"7HuA�ޫjB&5D�xH��JqtX�@G<���7D�� "�ӈ].�ֱ��띥J	*dт"O
���	�x/����;�8��"OD̻�F��L��y`��1��5�"O6�!�B[+)n@	3�l0w"O戚щ��v\��;��׮zj<rs"OZIV�K7NX@=�ģ�Jw�l��"ObȲS�U�	����;jO~�k�"O�D��H��s�>�8g*�9:2yb"O����^�%�)�^Uɬ���"O܁���P]@��� ����D"Oಖ`�der&��� �.eK�"O��qUB�|4´��͛]�>���'�8�q�b�o��q;t�]@LD��G�L@8¨�ãM#n�>��ȓgXYx��"Na4��%�\�(���	��ɺV��.v�ɳ�Ɏ{H\�ȓ(-H	��dN@:���	���x���t�a�(�tG�qIq ӑV����H��ӧ��?��MA (X�hbp�ȓK.�G	Z�/m���o-?Jq�ȓ=��	�4(�.�,���׳:�8	�ȓ3�����Z�j˲P�V��B�S�<c���g4�<2�&P�l�����R�<�2�[���
��\��Ƞ��Q�<a�+O�"�0����Q��B#�Y�<i��J ?o��	੝�'w�:�$�T�<�BO�~􀝀l"|�Q�kT�<Q�?_R� ���&Ui��i�<aä�1)n��p��y;n���D_P�<�Sg��1t�4R G�;�LAdǞu�<1�	� �$�;#-�Y;�Z�#�M�<��ś4@ ���$�!C�2����o�<��N@p�F(؈S���bm�<����7Z/z B'���4�h�!'d�q�<��¾y���FU�'�GN�<1�.	��8�g���@m!��G�<Y�@�Fzx�a�S�L������F�<�CW4xxC��H-u[ �z5*�[�<�	O�w����[�
��4�c�<�q�u��IQƘ��X�4o|�<��NV���� ���0$4"3J�l�<��AP*n�<��
�>=	r���@�<IM�.M�|ē�
�:���ól�^�<�r` 4d�)���[
 ��Rp�<��ʈ�2����0�zAZ"��N�<)W
<D���e按)��A
a`�M�<	'l
8��1�Ō	F6���dTr�<�#��6G8]�w��9��EZ�B�p�<�Ӧp��) ��s�~��SgD�<���΅��[2iS�9��ٱ�I�k�<�,ur���֚>2��`g[g�<� �;apu{ǁ�x�D]��w�<�f��_�pm9qC^�/��!Q#Kz�<��ۻt�QB��%Y�]91�r�<��ʹ���b`�ƒ**�%����i�<�We]�<iFx ꃑV�x���d�<�t��lg(����*m=n�b@JU�<	gaD�'y����%�=�8�B1�F[�<A�(�qfb���j��B�/^K�<��bK$
�����)}	��q�D�<�o�>h;�AXǩ�HV*)����h�<���i@��Ҁ�7.�J�� a�<�d�Џ~���%�W��*凗z�<��j�y͒�!���G�n�g`�m�<1�KK�qcl���[ b��tk�@S�<� x-�8H6Îc��0z2"O4(:׬Բ�F� ���`���V"O�}+P�J]'����£;ޚQQ"O�E�b����PSY�:��`B`"O�5�i�Wbn���
Q&1��|�"O��@���b}�b��C�`�W"O �d"�&V�� �W7V@��#"ODC$�Ӝ2.�l��W)=Ox ��"O�Q2�#�E24#��(��]X�"O<��#�$����BݼD�� q�"O��1�G=z�)��1U�QK"On�Т�� KK�����\.9���"O^t�$ ���T��h��D�ib6"O2A1�jȦe]��倪f~���"O
���EY7S(DQ�je^��r"O��H��-u����#7R.K"O ��(��}�Ib��N�H�b"O �&�+2Jm�e��)"hU��"O�X@���H���JR�5R�6S�"O�pD [�*))T��?Ȭ<&"O�|>.�\x5/�&Lmc�'ͼ肧e_�KwH�h�q�Ҡr�'��L %Hַ&i԰��	i2�!�'�.�9�-��3c(��U�Ԫ�&���'��4�r���@�t	E�Y�c����'�@$�CaN�.6-�d���D��	�'�,��q)�v[rQ#ՠ�4���'uܜ��J�!�� !"L֛�rDz�'���S&n��5���(< �' ��8#*�I�D؄.�� >j<J�'j�����Ĵ
�p�%�إcoT��	�')��Ĩ�H��%pA^�qq4	�'�jD	����h��h
�Md�ꘚ
�':n��U+.0�V(E^�`�'���k�Y�3��D���*2<�U�	�'O�u�'�Z� ���2a���k�'mF��G��Ef����:`+��1�'�Ԕ��EÎu\n���$� B�e��'fJ���� �N����c��:�3�'8F=@@C�s�@���#A�>f6���'ڪ���hF"�d�@`� �=!.tC�'�F9���ǒv��Ѓ�z�
�'܀�	þ2�`$QB��R̺� �'c�"rȿej��e��r�(@�
�'θ�0�UOW��[E�[�p��AK
�'�Yk��B�F�"�amT\4P�'�20Ӂ,�iq0�6����0�'ዲ�8!�(h���ƍ�F�p�'��	�3/B�-���`�Ÿ�V�	�'�8��RH\�]��s ��31gd%�	�'��P"�	�0�i0�ͷRI�<��'R�	H�ܙ��ó.ãs)Vx��'r���**��i�ʎ4d��@��'����CR�yp������F��B�' 5���E�o3�}*�@�J+X���'q��Y�d�0'$�d�)�X6��Y�'����G�={�2�N������'y(��lª#�"�i�س9J��8�'d��Ŧ%��HbT�ߒbg�%�'���(��ǝ��-Cԡb~䑑�'*��������yː�^2(���'+>e�r��(C
��.B�z��<��'� ,��v�����3u�ܜ1�'j��s )��.�f�9r/%��X	��� \�`�������$L�h����"O:a��� ,���DY�H�l�E"O襨�J��<TYR� ��\ؔ"O !�,�0�"p��+k/6�#"O�J�4f�q�s�f�RQ�"OlԠe�ܻc��h��� �+3��'"O.<�cM4��m�&�(��"OB��dL&6xU�C�<0crA3"O@�j��E!e��M��߃~P���P"O�(B�ɝv��8[�
�I��鉱"OXXQ���&����%jA������"O ���_��
���n��E����"OL$F��P-���ǫ |�=��"O���-�o��ba��7x����"OBIh+�x(d}��՜w|,��"O$ӃIU�0��졧DN$MT4�R"O���7�A#�@��K�K�10"O�m@.I�]6� .` ��8T"Ol 9VG_=�E	O�mZt�p"Ox�:f�;J�x�2(I?N���"O��a�&De�P�UG�"����"O&��D* *�� ��+��e�7"O����ǚsz~���쀦8�T�"On�IӺB��!�������
�y�.�6�l,�����hc&�)�y2I��7�" a��
x�Pvb�4�yD����,��&�(	p �s��«�y��
g���D=�(I���O��yr^5Uj!A0 ܼ7�X԰#N��y/D��\(Q���h����^��yrF>}�|����m�z%J-T��y��è�|-B�΃�:�~��UfH��y��g5�M+�Ǚ�?�����.�y2��w�N�x5&N
ω
�yb�L�1�|� �H��`ˀ��=�y���"B2����B���<A�l��yB&�;l����ף��-����&��ybbC;�"`vEA�MU�pY�F��y�&�(F����C���I}�]T��y��Oj�Ȧ.Q�B����`̡�y�	�	y�4����
���k�F��y�J6�2�������!&�
��y��7$(��j��A2L��ߗ�y�N����"h!���`ȕ�yBG��^}�V[�1���Hei��y�ā�JݚlZ���`�(\���7�yBO�_��蒒�V�j̀���y��1����!ۘT4jֆ�y�S�c>5��JW�;(���V#�y�!C1	�"Iω<�.t����y��"pUfH�V��69�F,�� ��y`8HFD�5�P�1WZT����yŃT�"ESv�Y�ԀJè 3�yB�����\>%o��0MF��y�BC�N"=�V�պ2w�Y�*��yba��_�4���� �2�`v(I��y��M@��Q�F��6	�Qj�����y��[�%*�1�qg.�|H�5+��y���iH"�(�D�$�������y�kڇlMn0�P "�IA���y�L�h������ѯU$��@l��y���&%��q�Ҿl� ��?�yrI=M�����Y6�	cd��y�a�7&[�1����,~?���4��y
� Ɖ��d���4�J��;a��,��"O\L�^*�8�
��� G ���"O"5�R�.Xa�48 -�-=�F��3"O�h8���^|<0�"�'��e"OBa9�C�>L�@Y���>f��2�"O��@���Y�,r��L<>_�e�q"O�u	%�>�*���ƥ~�pԠ%"O -�tJJ�-�ru�A���D�h��c"O��b,ƃG����!o�j5J�7"Oj��Ň �3��B��@�	&j�{"O���3�*]�W)Ҁ%	�d�f̚G�<��)�,����Vi[�c?�d�C�<�P.Y*d|�� `���h�$�]�<�dk���6>�V�0��=`�&�����x��扅A���"�.S������셠�@W�&.فI��[�	��ɗk�`�g��d��ز� �h�h�D^�K�N��ƥ�##t!���g0y��`��R��z���c!�$#<�r��NJ�G�8�Jg��!�dMY6,�f�M�R���W�V�!��5w��Q�*V��6�5Uz!�D	�?ԅ�g%ײLX�U�%^!򤐌	SH�q��w�\��r�T�N!�'bu����Q��p����x.!�M�P��Bu����7���9!�d��q�~䲱�֟3��̰���X�!��Ut�C�ˬw��ȰQO<!�!�$��L������P�qFv��!�ߓvd!�D�e��R��V�?����^��!���%����g�G�i[dT��쇻Y�!��C�]��Hc���"$����IW��!�D��e��M�Bb�'֔x�ϴ}!���~4,�A�D�R�(�*q�ʾNp!���:�����퇕b��0@Tg�$]�!��/�Ɯ*M	�C�`��&��N!���kl����7?:�����rR!�䙾v� q4S�@�0{%f��!�$[�k�R�8���1^oHٗn�{�!�d��j�{S�ںIF���@��~!�\�������-{0���Ί�`!�D �I(K1cNRZ�8`��PW!�d'̘��D�͵s/��(���R9!�DF�T��`�|�؅����@-!�d�[E�`r�M�5R���b���wv!�[�@`RGD�t[�.�|�!�ܡG�:�����Qy2$c7�=V�!�D.8�
)s6fўGdB�uJ�?�!��N6OD��If(@(SL�嫗��+�!��S��m�S�V,$D�������!�����=���M'	h��	�;S!�D�i���k�jX�z!Z�)�W�!�D��zLh�IU�
sjH�'hԛz�!���Y)JR�+�-u�Bd��!�H�1�&�S�JKh���K�0!�6��%�1�"vꁨDAT�G!�$,�
aȃ$��`c���/Gl!�!	BV�j�ˑ?ZJlP*�NB�!�$%�T�8��-��[$mɦpi!�Kz^�����3��U�V,5!�$�xH����׍�走�&89!��Ц`&6@���ր ڴ�I#g8!�dN�|�,\b�&#M)�	A�)�!�D�6+��GG^`#j)q@�[�I�!�$0zƌ�H��թ}��sc@6K�!�� V�J,�5����f�/E�;�"O4u�t?���(u�
-j��J�"O]G�Y"ywPMCW'�mۆ�ó"O�t�5Җ1���C��*+��A"O���U��=
@�<��f,h�T���"O��V�[�sLX���H�H�ڴ"O �ԠK$.T �-�x	nY"O���En����3N�:��D�S"O���T1*D����"����"O��Jtm<$��{ehD�k0�!�'�6�a���Kb p�p�Ю-�TX�'C`�#��)H`�Ç?& J%�
�':��CeO�XH��!��U	�'E�)�mQr�8�� �+lK�=��'UV��!�7$�Z` �ҷs 8`x�'��̃3n[��f�IaA�%X#L�8
�'I��a��{�Le`�M�8L�	�'_L9:����%��qW�-K_�1��'���Tիt��6�)L���' �|##��%f��PabD�G���*�'b�їᇜ�E�1g�%=���'6� 	�E��Y}� -"	j@��'�4����5Ad��qÃ7�p��'��uB�c�Z�.h��I��a�(D���h�"�6���i�&ۢ^ &X��{��x��Ře>`م%��-�,���JB�����
u°Đp�C�e�*��ȓL�6M"����h�ژ�\��5�zq���6����w)\=��	��4wԈ�g�Gk�X�3�::d��F���weJ�*�D�D��iQ8$�ȓc�T���  L<S���,!�x��5N�Ep�\ �(��4	62���,�ĝ1��'=�� $
�z���$����I�+e��wl]if����=9�FB�I���e�;�l؉b�A�&�tB�I�����a�[�<�h$����u�B�ɿ^4�JG�J�g��T#�=��C�	�~w�Q���y� ت2��&MD�C�ɀhm^�P���8�K@�!�xC�1&C���C��w}F%�tF��BC�p�R��q$�^xh�
��yJC�Ʉ/�=p�'l�4T B.�ZrB�.~�6�1.��i��0H�abB�I��sfF���@z�Q�`�fC��fQD���ءZEd� SN��NC�IK)���0�R�M=��'.Q��&C�j����e��Xm���`�HI�C��"E6B�r�e�sl8@I�j
%t��$H��`A��!���:(F��!�D�iQ�`��e�$`��
��!��Kzॉ����6�a��E�q"!��9h8��� CO�<�u}!�$z�����R�~M"nW�!��;,�`89�ǈQ��m� .2!�䎲r(q���-n�4�!���3*!�D�v���aV2b�v�����z!�$�t`|-h�W��x���Άjs!�D^>Z��Ƀ�KJHg�ѱvb�Ll!���fM~�7�\6=b2�8�`ͨ0{!��Y�i� P�bm��$������U/e�!��W U�5�(��}����g&�!���u�(dX��(
�n�i�%	2�!��<<*�:���l�lrӄϳ�!�� $`���Z�	u��z�gUr�,�R7"O`|{��R� ���[�E�>�	�"OX�X�A��H ���n��0Yv"O����J&Q�`���:Q� `y1"O��!'U:3 ) B�rX�T"Oޭ��FG3۔��"� �{s
���"O�	3#�� � r���OU���"O|��D�7U�$ �gfB3O�&"O�h�ǌ�!����Ɣ�VЪ00"O�]bT˓.y���
�E����2"Ot��G�2At�A*Y�^����"O����;�v%i�Y��!�g"O�d�UnS�3�����A�##d��"O���M+l��-[6׍iA!"O\�`#�H�c��ZB��)'	�+""O��IR��7X�PX��G=`����"O\���BM�Q��X���#9�v�f"Ox}S��L"yL`��c��V�"@��"O"�#�lÐ}�d�P!¯0�@� u"Op�A��+R���:*u�6"O���-X1w��Ƥ^B����"OnL��Ə�8�V�R��'1�Z4�p"O�(��A�"6��s	��<\��z�"O�dsb �}~��S�Vt0P�"�"O������j�^�Jc��>&Y!�"O�ܠ@(ˤ8+^��5g[�4��'��"Ba����`÷>j@��'k�	�e�+U�f!(ҋ��!~~8��'b:��S-��"���B�@�	�����'vܪ!��/$SNX��Q/����'l,p��ߴt<z�0�[�Ψ���'�*�ҧ8���{��̑���
�'܈�aΊ�)��H�Sx
�
�'�H+Ɗ	6j,���T��c�����'Rr ���kXUB��.��(��'���2�/&h|���]175��B�'~:t(7�i ���b�<Y:���
�'~(�� ׊B�挢���U����
�'�>��&�آL ��Д �6q�ȡ�'?�ȗ� �h��S� �!��!��'=������ڈ��e�@x1��'6�]�IB�*Ŧ�;�!G�u����'˼���k�=W_"	y5�Œ]��]�
�'yڠ3���?�Pj�Z�%��@��'�P��c��4a�bP�EA8����'�4���Q��Pe���` �8��'���1�o��U�T)���?SV�!��'�T�sƈ�7a(L�3d� �h �'4@�@�&	NHx��k̮j���'{����?i^�$ԏ�f�N���'���q�H�R�$�N8^�����'�6�*��V�搜�4���h���'K.��w
Ӥ�:dd�O��|k�'|Z�������ų����P5�M
�'B���47�P`��,�<D���'�ȥ��U����(?�P�'�.�(!��4����ȶgb�H�'8ni�A�N�茸��U6b	���'�|���
�Jh�#'�1Vx�99�'dh�tf{��hƣM�<�P�A�'�Fe�k:0�ܹk� \�3�2q��'��e E��6i:H���G7,�$L�
�'_x�)���k��`�@�sO�q�	�'PMyv��-�r�2GK�6������ �(�7	��9౥�HRk�1�"O�<h�e�$C
ĵj�,�"O���Ù�^��H`�H�
'"O��dʁ~��p(6��c�0��"O ĲĀ�d_2��5f�5�|���"O�d
AL������ET�H	��"O��t��1T! A�a�ڐ)2�2�"O�(:� ��2���	�* "|b�"O��QO�X��]VKh����"O|�s�c���b�KƦW87"O�}Gz�@�����a�"O,��w%�{��̗I�a6"OV�E�W/g0�ų+�/�]bp"O���7%�>.�8]S��k XUP"O��;�Ǚ;r�v5� ��e�V5��"O�9�͙:KH��s�A��!w��X"O�z&��Aa4�"ƀ�JY��"O�"х���2�[D�D>u�\��"O�ׁ��	���%Ŋ}��ѡ�"O�
g�]�G��9kʊb��$s�"O�� E䘘l���	>&�u�"O�M2Ae|�ru��"�����'�PI�2���J2D<�gúB�X�	�'qD(�E�]��T*0,R/5G��;	�'��\P��������G΋&����'?���K|x' $n�J�'��q�
\�sv����CG�u�`��'`h-j$E����e④��l��|��'3��o��y���!@Ae�piq�'�t��%��lXP��������'�� �i {�($����q����ʓ*lօq���a{t��C-�~�tp��A����JB�1�A��ğd4b�ȓX�+�e��Y!��$?��E��,8  {t�Q�*}�Y§���@�ȓn�F1@����  `'��3��ІȓP�J 	�;&��f��O���ȓL�����cC�&�0�ٳEN&j�L���I0��d&M�ze:\óA����ȓX�,���#��-�|��-�!s0̆�Zz��"���fL�v�7k��,��M|�P�����n��Rc�a�@p�ȓ�����7��aF^7g!�y���j@�M�c�U�E��:�, �ȓ.�N��,T9 X�Ǣ%N���ȓh ����&��_�ܑ閫C
��ņ�%2�Hk��O�1�hP��f�A؂t��B���$-��p��$�W�C41�@�ȓΪ]ʆ)F��"9�g��E?NمȓCĵ�
	~ۄI�b�]�݅ȓH���2�l��4�%䇙]�8T����I��O�>: �k#f��Dμ�����5�=R( �4�A�i�<��4)��q�n�}��y� 7V�T��1M(��Q`�Y��9I��-A��%�ȓTɪ$��@;C��� /�<����Y��)��
�t�q��(����M������T�?��	��a�$mΚ��ȓw�D��gAA�Lz�ي���&�9��U^�mʒ�I{�]�e��+rnH�ȓv�0����K0)qP�8Q�'u�TQ����a3�g_���8�Шq"��ȓR`D���؎���Pή"κ���*(nd�����wg�����Vgpx��S�? R��@�Ԇ9^,0���#+��峑"O�A�%KN5c�*x@�KG��,��"ON�8��-Ph0j �N.�ك"O(���]3�d�k�i�E��J�"O@�@���9������4��&"Obe���y4f��s�ǂtc����"OF�e'Iy�`�����!� "OR��$��6G�N��C�ЕV�ԀЗ"O���S��j�͛�U��h�y�"O��SFd��@��b�O+��e�"Od���!Ȍ	��<�ƃY7yg��
2"O�yaDQ,1A����Z�Db�u	�"O�l���֝<mX�O�W�갰�"O���dFRu�4-�dnË(�jPPb"O^��q�H�"��K��d�!�"O�|�"CDL�b�⁫P4!��k��,s� ٜ)�	iFꃪG&!�D��XT��h�@�H��)�2�!�dPi��UB�C�2���ې�ͮE!��y��\3���.��p�E�68!�\�C�\e�'�.C���1*�/Y$!��P,D 8�ˏ?�� ��A!��/T����9�����BH)m�!��S(<����,�|�3ᣕ52D!���ks��С�u�V�{ÌOw!�d-C�)e,̚�,��q� �R�!��Ўq��M`QjN�D�ܹ@Ѡ�8t�!�D�" �\s���v���07���!��Bvze�Vh[#q)6l�C�B+h`!�D
�J�d ���"75±��_�]\!��ܳ"�8�hr��r*�� acұg-!�"�`+�W=T$P��h��)��~�KC�<Q�猫^���*�O�Z���	�j�<��Î7�6U��=F�ΰ����i�'{�E�T$��G��};��Z&z$����ʨ�y�L4�-UH���Z6YA¤��~�)ڧM��q���&~̲s���L���� AF�(yK8��lҿy���}�Nd���l�"�������H�|���#LJ6%�E�Blnц�N���P�F����j�b�Ȇ�]���+���}u(�R��U1����~p��D��9D|����6q��ȓ;8N]�� E�"�`���C0�\�ȓu�օ�H�?�z�2��\VH��ȓ0SV���E	�0'OCkbi��F�<����G�H����"�0,�ȓwH��D��Ҵ}hg �u�vm��[��PK1˙oAt�Æ�y�(<�ȓ!�|e��ܻb�
���ޒ'� ��ȓ�|8�5o�4�F��crs�фȓc��Ա�i�2?$�y�C�6t:݆�K��WDv�J���ժ'7�JC"O�eж��<�\�8��8E�T�Aq"O���'�-Hب1�F���3�"O�eys�����6���\܋�"O,`�5��(H(�"�BM"Fv���"O�m�� HD�kR�v���B�"O�H�7�K�7�8��?]M�E�C"O�E&���J^p��� �8,9P�Y6"O0T�����,f��:�gC�iP"Oؙ�����8�
`@Ӿ5t̛�"O���E��Z"��L�x��u �"O8i����e��Ah�CJ�`�L�R"O� Z�U���LZZ�'�
��`)c"Oh�:�!ͪb�@8���Z72�~!�>��(Ef��4���Ж3Y�u�p��c���#�O�P���'^�SAM�<?~ �)�D�`�x���'��s#dnhT��ƙ�P`���W& $�#}*���!t���J�j�9�u,Ps�<	4�W�q�=y�Dٽ?.BU�i�o?�3�����h�h�#FJ��1n 3`�����"O�d8�h�q��9K��C1��� ��>���)J���)�t�h"���j1����=*-����V�+�܈���XeJ��@)]2'a�I�.��!�<!l�f,�	� 2�͊�Y����a��d�OX���'��T�
i�&���b}�d�'Q�Xc�$Ų�:V�LL����'|ў�}���A%2[5���^1��ڕ�A{�<QSZ=��ZE�ׄgu�$:��z�I}8�q�̔�^��d!��[5	�Hh��'�O^��'�:9��ل6���sc��' *� a
�'�r��S�I�G($Uk��C6BD���$[#���E�ď�1����S~�p���9�y�aƤe�,d 1	�O��i w�F��~R�Ѧy�>E��	f���j�`�q��=��hQ��yb�ހn�"EHV_o4;�B٪��'X"��dR1L.��`ޡ�l��
��!�D�"&���`	���*d�C4�!�ϓN%h��i0B�U�H� i�!�DH4潱Ј�7�D�`eG�&�!��M�
��%��+��kD[FۻS�!�=V�l�q���E�Fy$!�ֻM�jŚ3�(l���Xq�(O=!�D�����[l�\���P72(!�D��o�:��f��]��I�u��'�!�D�xdm���ބ{�|�&��5�!�$�����v���&$�'�6�!��A�a��pQbl��K���	����!�$� [F�hU�4x�'���!��ʽ�h�\\j!���M�!��m9���"Z�b�<*��ڮ/~!�d��P�����߰���2$�=?b!�D�:
^�IU'�7���7�գg\!�$��*||��FF�Fq�!�L�^?!��E��� �@�r�
H�����O]!��[�i�.�G�&chp�Iw���M��ęX�Р1�喕y[f���y��D	�E��H&�����	Ǎ�y��źRi�=�'��8�񻴈���y�d��o찤Y�&�;2"���p�H��y��;�a��jE,x6��Q�fS/�y�dT
x��
�%��jD�\��y�(N9q"���c�&,6������y�(�$&����@����
P%J�y"�#����^
��%��h��yo=X��y0BL�6�u���˫�yZ�С`C��WO،��K�>8�܇ȓ!�n�K�mW�Gil�{��<6�����6��u�B?���r%B0bm @�ȓ>*��۱�	%�Xm1��!
tv%��s����k�Z�f�8f/�,�*5��%�dx��`��5&���g�:�Tp��z���1#��8I�.9����
�Y�ȓ��s��ݬ�\(�+UA��=�ȓ-b���Q�Δ5b�a��Ju��@�f���ş$8F\�1�ݫjK����c����E�Iڜ��s(I�9	����S�? zik�S�TGđWc��N�(��"Oڍ����5:hq��Lm�r�IP"OR�1�c���P͓B�A�5�h�jS"O�q���.Yj��8QBC+<�td��"OR�hBGД�bM�րMn-��i"O�	 �lB
ux���� ���"�"O��{5#��'��M�� �9"~�8�"O�qIPȎP&XzҌT'+#r��"O�x����@t��%xj��Ѱ"O�]�҇��HjTsPb��tj"O^a1D�-���D�_�	�|؀"O�Ĩ�'I@���@T��8�"Ol�U��~�0�q��M�`���"Ox ��&�"�n�p�l�_�5��"OHdS�W+~:m� k�{�n�� "O�m)S�ޥ<����Ȑ�j�n��U"Oftcj�,������QcY�ݙ�"OaQ"�|_|����2(�N�(�"O��[����\��m�l��Q��"Of@c0��
hr���+F;<�ʹ#"O0�å�	-2��y���ȟJn$ȳ�"O,dh��D�yⶽPd��
	dtaG"O���̈́��d�y�L����1�"OT�lD:R�r��Ơt��}Keo3�O
�d��@-Z�Ps/c�h��7K�n��8�C�p�����֟<U�
�B�(iR�*&�L��#��$pH�Чo|p`!A�Ƭ>M�$�ٴBi$Fy���;��\�A`�,����$
F,31$5�F��J@6H�ѩ N�pK0D�(^Ħ$���MxܓcQ}�	�O"8�����jT㇄lE���7&)�ē�?�����'��S�Ti8�(�e��Q��Ԋ��ٿ-�B�IG�&,S ��x��:���]��I��M�Ѹi]�Iy(���ش�?������̳(�6x��ߒ\�*��ef�ʌ�`��ӟl�	����to�ȸ���e���:�ř�T�\���д.`&���ˍ�nlF�ڕX9�ң<���>�z��\�q�vxi�EH�� �ph�}���P[��׏�*���#�NQy�*\?�?Q�i��>�!đ�C� $�6A�Z�]��G��xFR���`��C�+T!-y�����I��|2�dӶ�n�����5[`.�`<~��<ȁ ��@نOч�M�����?�'�03�Ʒ.����L'n1�ܒ�!05�芑��4(�&�㶥E0kq0�A�a˷dp��O����2:Ł�J��f~�Ƀ5Ú�z�R�oZ�Ѳ�'
C:Cج�3�	�1z�����\��}��hΰE�'�a$��`A �Ruoڶi�
�$�-KAP��	9��)0uOV;,'�)��h�g��)�@�� ��S���A5�A�`� S�h�R�\,o!�yDy�m~�t!o�B�	�?Ѭ;:<�p�g凚0(J���MTr����'�(��y̘1��'ub�'��l�I�	ަe`�l�&�{�#ʚJ���+B����~�A�Q&#<4��mD<c<eh�'_�er�$�H�U�����<a:�	���=�$hpf�B�6k�����0��(�3I�~��4�lچ1��ɔ}��
�bԋl��Ǣ��%���^��I��M� �x2�'UrR�d+��]73ߒ���B�B[�j7Ϋ� ��I����$T#T��JA�KU �����/O���d��OT�)��jʓb�2���P]��"��_�m�H��_�'�$�����?����?e/���?����?AG�R!c�4hk��Պ�L1��-@��;f��'^ =	��T9/������Y/�EEy�g�2�q���b.�C�ZQ�d tl�
k�X��F��2d��I{�,7�baܪa�<1F�����3p��(��YFn;Y����'��%�H<)��?	�*��� �K�^颔b�N��<��#^��F{��I׾m<�1o��-���+s�~���ʦ8�4����pF��'�T?i��)��/"�٢��YQ/���2��/��|����?��%A��P��>9q@e[סY EJR|�fi>a��V�
���Ձ/�H�@�%ғ_n�wIלe Ju,�zF�l��H��� 
M��Cv�:bI{�ፘ��hIO>q���֟�R�43����'��\���a�.�
AEHi�삋Bz�!��������!�8��C�ȞX�ژ�W�ɺ�p=q�I����|�$7m��H,h�$���!Ő�s	ۚ�qO��$"��$��8an��   �4   
  �  I  )  4  ,<  mB  �H  	O  YU  �[   _   Ĵ���	����Zv)���P��@_zX�B��S���A�@�8K��$�.?�����ɐ8��2��]hֱ�'*�01�fՓTE�<6D�'�_�V���
>�O��7��&��8Z�"�e=<�S' ��|_�Uz�
'<~�I�B@;{ʈi7�_���b"$�qld�#��`g�Hs�����rA@<NI�� �Ɇ+y���PS(�$,�EEK�h�D�27!���J�C�5Oa��('ʁ%e����D[�/����(q0M"�"��i�B� 0e>����A��'�?9��?��\��O�qڰ��/X�ΐ��!<ǪᲵ�P�;�*m����}x�Q�v)w�qW�c�u��Q��O�94"��/Dz�����$ u	DG]�kO��ұ �'}�j�:��Is�ӂo�>U���`1��l�6Yqt͈[謻`(^P�漗'mh-���,G�6 �d�O�d��$����+��ɮ�m�0	������O��d-���� �F�D*cŊ�@�FR��7��Q�ݴ��������P�]A4��#�yV�٢e+I^y8��	 "5����O����Od%���?!�����IkɪA�D`��d'B�U�����u#ҭS�V�aՄ�c���f^�eGy�!R�a�� �b�/2~z�svG�tԠц�?ˮr�	�U��˗WaI�k� �'fI���D��S�Ψl~���ā*&�q !"O@�Q��.<�"D�)ܔ�5�'UQ��y4o�� �RI�h�b$�@#�>)c�i �'0�)j��'*��'v���z��ҁ�ή�Q���{�����=W1�'�r.V6lm�ԟX�W�;4�n�xa��-��y�ɭ!��~��hֱs�����	ՂR�r����Bt�'��5��44>���O�aR=�K͕_j��v�:D� ;��+j�R��w��v�@D�WH9�O�|�'�u����sk
a`��ҽ�x9i�O�u{���O����O<�'re�@���?�%�G&�$��`�٫I>Y`�n��)����T�%wb�T>c�T��g�67�����&
��Qj�O����)�M,�RG�԰Xo�0��A-�����vPN�	1��S�O��ܨ�/ϣl�@ ӑ&J-1����"OT%���ʏS�=S7%���!0��>�ȟ��wd[�_a�06���-��h ������ʟ��Wg���I�� �	ڟt;Xw
Zc(֤#�$�.7�ԥ`f)x��h.OR�2��';�Q�#뀂?-�e
�F%C.<��-Op���'j585k�>��`��/#?a��-O�J��'���D��lj���BּyR�	��f��!�D9i<�<@����[P�	�w&�\���b8��|JM>id+3n<X��!�vC@�
�#�@�rAI��ބ�?���?������O��x>���#�Oj`��˲Q?�|�G��S��Zx��*�&���X��'���)�3Ңe	�
*�O�u	��'QL��
;(�(�� 5	�h�da;D��F�(�!���È�@Ia9D�4r�X>o��`�g�( �4��b�>�ӹiG�'<2<je�'M��'h���K#D!��@�4E����"��+~��F]�f��'>�V��ԟ*�sG�L&����)�^�R1�		=���~�ť�E��Ő2/n M{6ƐW�'YpqY�b�>%)Ƨ�e<�	���˕{I��sb�&D�D %(Tuit���Nɑ9P��i1�O�]�'��=x�fu<t�1�ȽQH䬡�O	(`�O��$�O�ʧ0�� ����?y�H��3�TC�"Q�b�Q�
/T��V��\B�T>c��+G���bu�a�kS�P���O*��r�)�')�u�DZ�vR<��Y�C�t���bI�-��1��S�OäqR�-:!��1�!�8jdL��"OD8s�cK
���t��m98AC���%�ȟ�������b1����)OF��4 E��5�	��� �f�5f���ϟD��ɟ���ȟ��Q�f���!хFaKB�x ���vX�8�� �O��I��.���%�4]L 36U���E�:�O�K�G@(��X��o�����U�p�cE�OvA��� *&V�3 dE�
$ʑ�1�ۿk?�B�	�sWbmyl�
@�=q���d|�6�S����|r�P�\U`jF��D�2�I ��-j��q�K`��'1B�'(��ڟ��I�|
�BDڟ��ÃH�,���-Qƨ���^���>��#Sn?� ���=e١N/��!pJgx��p��OJ|�.W�N_,캓g��TPa�.d�<Ѱ���V�J�7<*��Q��^�!�$ǜk�E�6B�!¾pX5B7Rg�I�MJ>�"dR�ݛ��'�bޟv�aኾ��dC�q!x�)r�iǾ��'�'h"�'U P[3�'1O��T�F�D�q	N0L��w�ȀCўPV-=�g�? ��A�ıF� H���_-�qx��I�%!N�� C�O�Ie��Sװ�R�T����b	�'ܼ�X@Můi\Ra	U���0cH�	����3Pd��b!��:B�d��t��>n2�+`)����?�����	�>�����O�^a��y�gMR?tȲ�c���3Ѫ�؟��<���'��1�� .ʐ��&�Mʌ��� �đGx�����dD����9[~`��P�ֆ��FJ�2�%���A[æ�'4 p2J[�AۈІ�z%(�25�@2��� �^&0Gz�n&�
�tPho�*m?VSbh�6}^�v�i��'�
�`���"�r�'��'s����֘�}�t�ٵ��BU�q��BL;kq˓A�ń�	�;w�y(vgU�i�V�9'�}��vn~���x�&�#���t����;תʓU���I�0=ٵ�-R��ѸGШ^���RTa�U�<��=W�Աq҇�'�j� 3F�Ӧ}H��4�֓O�i)��ܽO�����V>]m~��@�GAb� C��O���O\��Y�����?�OB�MH����)���J��Y	���}� ���'�X���']�( ;]0ؔ�%d�1j�q�i�����#R<�AaF��Njy����j�X0�'�J����H�&����H�5hfn= �'4,�R���YÞ�BċRb6A��O�1m�k�I�1�n�k�4�?I������
�7�Y�b��:��âR�M�e��"�?A���?�r#��?I�y�O	��SP#2=��f�4 �|2��$���Q?���OQ
�
ᨖ�Z�b�[�M?ړ~*(��I6��de�@&�_���`�_3x�4MQ"Op=b�$>\,�t��)Ɏ�уf�'��� 4Á듞%+�ղqb��E�.��'����vӒ�d�O�˧|��@���?�7L���]aT��1�Ԝ��&�9\��fc��"�T>c�ԁ�`֌�x(��#��>s�\�%��O�qɂ�)�Y� !)׬=�ɹQ�T�Y�fa��q�:���>��S�O�QD��?�L����� )s"O����"h/v�{s`�%��� ����ȟ~��v)�|N��(��J�n�T��Ц��	���[b������������"^wLZc�t�����8��%_0^�<A)O�|���'2X�@f�L�?)2�Q�?3���(Op��'��-a��Ӹ0m�0eԖ!\P)O\@���'����DV�0���1�ʅ2 ���Υ<�!��15�����:�P��ћVN9��|
H>aĀ(	4F�r$CS�U��݊��'&���K��?����?!�N���O&�$f>��7	�O
���L��q��41͏� i*�JP��sx��3�H���r���O��eU��R`+��+�On+��'����l��l@4h��@�)D�~���=D�\�T�S�}^zY�-��vZ*��)(D��@�I�Pl�)� aq���d�>��i�'�~i	`�2�$�O�0I���f+O&cT*1n@�~�6힁
�z�$�O�ѐW�&��7�?��G�S�2`3�+ߗh �)�tN>ړZ�&AF�$hS���q��J�d�`��g�hO����'��"|�%Cq{��cN��M��0�!��t�<�U�*bn9�S�	�]��)��!�FX�L��O|� �LC����@�R��n��VQ���� *ߴ�?I���)\4\�$�O@)K3�ޜ��7\&���LJݦ�i�G��5��Y�ɍ�HnB��@�2~��n^���O
�z�8|L.\
1�#A�� �S�'��8��d�-'5;WHC�R�x3I����}���޸����'zr@���8	d�D�
\k"O%��S� n�Վ��"6���@� �xP�ȓ)9�����*����M�r���GzBH!�'g�����kA�T*ҋk�� w�i���'� �R�*׿�B�'���'4��]���X�+�v�A����>�b���?����C���%�T�{rj4Vg�|�O�|2��$$2K;�aνf��8P2#ʧi�>��A��,s% �e͒&
�r�X>%�PH�$ .JT�����<�c�A�`����,��_�����~y��2�?����?I�bӟ��3�M,}�@� @�'^i�G"Oq��@���aE%�"q��i�D#=�'�?�/O.��D�M�F���ɞ��0D��m�*����O��$�O��$�Ⱥ��?ɞO�p�3�Ğ-f�M(�M�.Xjxx����R�!��5��qhp�-!џ4RB`YBg
4�DC@7n�,)��΍�p(�$K�d>d���X�a��oځd��i9�L��g��m�I)Հ ���U�K/ 7D���00����imr�/��u[��N Z�FڸUo&�Q��,D�L��b_3 ��B�d�b�\;#��>���iI�W��y�����I�Or���JC������$��W��>I��6����$�O��$�2�`�k"-�-y��P���D��'8R����!,��B�J�l�5G{�ivd��'ϣ5Z�1`i
�N��̈��@�&��(�a�?l5���v�[�Q�
(�Q�W�D���Iӟ@�}"�.١uq�9GL��Cr�Cv�H`}b�'}�|"�_U2�Uw��@0���>�&���H��<��I��/}� K�>a7�~�v�'��_> 1i�ݟ��ɶwj��У������[v$F�)K�� �4=J���������$�3�(�H�Ɵ`ƎpJ���HH�m���O?a�	#�A7%��-�$lx'�OП�"*�O"�&�"~"���3�M���= kҠKpF��y���_�J�;`�A'x��Ì�HO�)E��W��m�T�l�>�p��\$m��6�O��$֚O<�p��ON���OB�D���{����[�>�밎�L��2��Q�uޞ�6��6��m�-8c��y�O��$��m�ɺ98i��ңt䙓䀢`��-�@�;*�F�{ba��&�x��|��41:Lm��Z�L�ɍ�񲁈Z�(7HX���
W.�˓i���I�0=A��W�c�l���.-T{d�sH<�UeO�`�	@��|�p�\ěV?��|J>��"���}k"	H�D�^$ه���N��ĺ� �6�?����?i��%����Oj�Dw>a���ŰT�RУ�ᑈ:�bq��ǚ�H+R��^4Y�9ɠi\>l@=�����NQ�#bR4-y*�X ��J�^T�b H4�Ѐgڀ��a��Z8�ԩ⯊+7u,L��,�I�8��$���@H[cʅ�y'�����V�ȓ_��qi�뀮1��р���J��]��^�Ik�D�t�V�0s)X ��'��7M%���?WI���O��ԟX$���N#�d�A@'["�Q{��i��, t�'0b�'����APY$IBW�=^����G}>��Dh�H�M��_�� %�<Kʵ��	[3�l��B'H��Zw� �Hs&ĭm�&�B�Ę+V$t���A�C�{�@����wܧ5dؘ�geM4}�Jy�!cL?lx�P�'l�~b�Ӷy���D�C5�)٢a
���>�E���;�!�0FR�Aa�2;b����>��N��?��?�*�����g�O��$O<q�4��`��1���%գlWJ\n�?�hK׀W�Q�htW�{�.)ટ�c>�xQ����1���4L?:""��ɟ��(<��M:2�	B��ɺ����*N��1���T�H�"q�"XyT�9� �v �O�%���?��O�O��j��3`��#'�RWGB�ȓN�h ;���7p��cGG�><�,LGz��%���1օDev�A�3e��@v�i�2�'v�y*�'X����'�b�'����'غ0P$�9)Kx0��!a@:A+qHu@!��dD	����b�1�ʧ�O�+"`��cC��`�@�Ĥ�9� ��\�;x����H�{ �S�X��ȫv���Bv*Y�ƃA���L�5a�
T�' �	��PF{2�O���Q��d9�<��
�y�8	"OBZ��"\u@�k��ܶ)�����i�H"=ͧ�?�/OPm�#H̶k��9A6�̍Y{*��'��J��O����O��D��c���?�O B�P/7A(.� �d =.���Be�� �F�x'^���%4o_џ�P+M�,Y<ٲ!�B��2Vj�l1��j�J��.�m@'m9T�Ftm�	a-�9�[�qO���1�]
1��O2�����i�ўPF}¬����֌��D� T�K�ybh�v܎���QǶ(�E I5����঵�	ey�� =T�'�?��O�h��A��*��p��+Q,v�ڴ/4����?q��i l��^�8245�f��AÄh�&2����� O�_��@�O�<[�fY+S�I�_�:����5DzH2%m_�n�ʜ�;CxBX�Q�S�H5���@��o�,� D�#��y�=1 �O��4�t�,y�Ҫ�<���f�pw���p?Qd��]�Xu���չL�`d{�AP~X�<3�Ox��u�J�y.�p��l����]�h�&�Ɵ`�	ܟ��O��X��'Y��,'��+ν]eV�фC�"03�6�F�	�yȴiA)ܚ�8�O8n��Od1��8��C8&H����f�*p����O�<� O�AX�-�Zպ���i���Y?FB|�O:v��ĥ,�U�ÎW4%v���'�F�I��p�䧦�	%��p0&MP�s
���ߕC�hB�	08$�4� ��<�@�Z�T�`"=i��S�;�x4����&,�{���M3f�kٴ�?���f�$;����?���?����B��IxR�P���!fFl���ݪ"�ޑU���C���c���]G-R!�k��R�'�썠�+����(r���E�n���͚�
�0�P/D�,�N�bJ����lӖ��D-Y�iq�	��BRn�cx&pQ)Xf���j9�d�O��=�꧀ �H��\0~LH��D��t��"OV`rd'!e4�� /�4}�j-zb�i�p#=ͧ�?(Or�yA��S�~�����p7 �B�C�.�Nh���OH���O��dȺ���?9�O�P��Y?(�5�bJ�@���Õ���9��� a�"M~�a�M�'\�џ�QcN�Z���h�K�i_B���@��q7b���$��TTt����zoTPnڐO;~t���$�	&�~«[�o@�p!�Ie�V$�B*W5C�7-:��Ot����ڑ�tb�9��83�"O0ȩ���(�Q1���G�:��!]���޴�?�,O�e����u�$�'s�)�1S@�EA"��FLs�HK���A�..Y��'nb(��Ys*P�s��h�@�+7B��f�*s;
t�"&S�A���p��;'`�=WL�5��4�ש�@p�h�	�u���?~XbG�	�5�tL��@2Xf�뢠	�ϸ'��������}j��͂g�> �ΒNb\�jgP}��'Y�����!������]	)�	�cD��-�h�1$ю�8�y$`��1q���F9Q���?������	�&���O�D S���9*e��X�ʉ��a]��%�$F[�p����i$g�v�ⅯL����+�S�A�IJ�ƹ�05`�k��7~X��0S� Z���&���rAέv����;!�J�c���r�IR�6L�S�Œ�2HȤ�FJϩe8�$�y?������4�>!Ƭ�<q&�Q4C�����a�oU}�<�ޜ]nY�wHM4,�pd�F��5�HOP�F�dbR,��ɖ�Onip� ���1bJ6��O��9z���ɕ��OD�$�O��$�(�D�\~�@��G�)�0��a���..|���B�_��A,^�+V��ꃆ�L�D�	>s>�r���E�\���1j�`���_�J��7!L�`"�T
��|�ڴ0�ɲ���d}�%U!V!��v;̹pW҃��d�x?���hO2���ʅ����O=��PuIo$B�ɕlH�ً3��,N��`��:�P7��N���$�'P�Iz��!�bE� J���(��I���b ��|PL4��������H^w\r�'T�)A�f;XY �L~@6Ŋwa�D�,3B	�}����U�^�hZT�qBD!�#�k5@��Hv,�x�D?���)�噿r���QFbԑAW `�`�P��Mcd�X���@�=�D�O�"5CQ�ve�1G��D��.	��mD{��ɨs.<�5C�+����A��3>$C�ɲu< �ʴ@O+p�,�aLR@��z��f�'���5H�+����$�?E�nF�[X�#'^$d�"�ɂFqӪ$8�A�O����O�h󧈇�t<H(�r�B�~���s��|�u0��5JW�E�%��rR^�')��H�Ł-]�M�R��Z����d�&��ZQаF�G|�(�tˌ�iaԴ8&�$t?����O������fpE
T�4ņ��O�����=GV�Q�F�L�(q�D�,ma}�6?I��O�xv@�R� �_b���B}B䉋c�6m�O��$�|��
��?!�A���BOV*����N
LyE�iNf��L�nU�����M���X�pBSS���Do�:N3���F��oA�}�0�E�B�C*kZY�ef�-�D�PDH��|3(��Fէ2(�iX>�H3I>V\�F�P��	MΟ��c�OpY$�"~�s��Ĕzv/��~���'���y�[>�8�"���L ��� T���'6"�?��|§AO'�ș���0f�-ɡ�� �v�'K2�D ��Dˆ�'DB�'�rgs���i�Ÿ�肬k9a�-C�R������ ��L{"��`���XgJS�8o�ם�|
�W
O8�����i�D;�`2oF��Bu*� 2T��$L�`����f�哋��$h��x�õ\Ol5��A+nLn�5%����K�2.6LO��R�T/d��PҠ������"O0t����p��FD���S��iAB"=ͧ��|uH���m MNha+�O߱X�(h�,"�����?y��?���� ���O��1޸i��� n �-�>gd�A��efq	aD��ء�0a��(�x�!��	�e�qyb���m�UA3�ꇣ ��
-Q��W�cc��Xs��I8�C��;6��ĆT��e�c�Ë���O׶,��݄ȓ:�P� dd ž�Qd�'jń��)�3O�c͐�(���=����']n6-)�$k����O�R֟r��OR<|,�l;�����i,\(���'b�'	iC6D�)9ƴx�FW"F*����w>�uO��5��9#��X��ź��3ړf��a�em	2T�`Ă�ƀ�CÆ���O�8A�+j�8CEkɶz��pa��d�'��'q�:ma��
X�nxRT�T�%�%iS���Ic8�ت$Ȕ7^K��b)یY�b C%�O�8�'�&���A
$!\P�1g'܁����d�{/�o���,��p�t���s��'��|�A�Рi'���+1'l$��gb�X
�-�ܠbdI�S�\�i��Lz��P�	��]�4,W�"�l�$�,?D��$�v��u(#
�`�nt�Baǵ3��}��O.U��zPJP����[��?)`�����c~J~���~Ba.2�ʌ��Ο�I�"LБ��y
� L�Ӥ���lS�݊���:.&y{u�	�ȟ6�T�>C4rEZ@��#,E��P�ꦅ�I�2� αz�������d���l1Yw>�M�{eȸss$˵.8(���L'e��e�Vc'&��zqO�?����-�|R��_�;��0�o�)~�I���+BU&�9g��C���pg�C�^�['R>�BD�/�	�.OZ�Jr+�=?��#�FD�Cn�7��������	R�������[�x{�_���@/K��y��$
ԉ44�q��ی�M���i>!��@y�`ƀZ�F�q��']��Kڴ���K_��m7M�O�̬��?Q����ԩ��3Tx�/Lnx�p�fF�4��M��KB2>�2A�� �p
f�Љ�<"���FybI�2������P=c��1��L
�i�C�Ǡ|����W)��d(���)ɠ�˗�4��3*���d�,R���Z�(ť&\E��cH�7�T���,�Bq�3��&8�Tp����]�ȓP���r�ԵOI��&Ɔ�N}���'ZP6-1��_�f���n���0�	{r��� �I�M� 7"��I�J�Ȧ)i�� �����˟�!Ȉ��J���(R02�����&�T� B�
5B�J�Dv=���� ��\�<1CG�
Gu{��N�ET�J`�-'u\��cg�D4�e��c�4h:6�c�.����<�С�ٟDC���V�O<	`�0"i��
4c�X�!�D��{��@�g��:1���&ǵR�a}¢;?�T�F�#3�x$%��Ga^��Pv}��,*�(6��Op�d�|�v��?i�+]�i[,��-�Kf��� W�i�.���C<e�87-�L\�n�t��Y>��s�VC�L��(�;T�ѕ=�Bhإ�'���)3�\&r���� �@�M���
�2�(e�G�I��Y8�D ʡo\/32�]�G"V�@OV�D�Yb�}�hMm�П<�O"1�D0�j�$�B`c3��x@���g��>����?i����D�O���O,ܙ���.D�:�X��8A����ֺ
��5mZd��䐭�2ʓ�?��'N*nl�@�Lv�rQcW�G���B�i���'U�]���Y�?J��'�R�'��םџP���B�V言�B�G����g� ?���S޴�[�*n8\��� �F|r��Oz��+��ʂ����B�n��}���D'u�N@p@����U�-��i;!��N��B�O�kE��\��j�g�(��i�%_��j6(�On����?1��~�k֔Ch�
�jƃE��=i#�R�����OT�D-��S����hE�I����e��#��7M�⟰nZa���?!��ry�&@?��s�h,�Ő�hL�H��%�@C�3F��'�B�'ȶ�]ӟX�I�|Bd.�m�0!� �oo�IP��Օr����6+C�7"�;���1/�]�-@�[��<�7kC�7P¸
ơ�
���G������À,<b<qҋLK0.�-z(!b�i)�S�'Ǻ�OB/�H  EIϗjm���O*D�`j�g�<H���Ge�f�Rv�"D�,*`Ã9PƝ؁G��TLk�`�>yűi��'�T��c�f���Ob��.�z1�2hL4$~�4j�BF�d7�9W���Ob��^�#1�$1�?-�E���3��.M:��Q5�<�hO�� C����A�g�B���$6�@�=9�Hџ��I�?�8��t��L��R��
�!�䗿Q*����fH�X�	����S;a}�N0?���hg��c(��f*�\��AJ}�̙�MBN6m�Od���|*�N��?!�\paz�LN.FL2T��[��)���i_u���'�1O�3�I4 ����S�@�yY�V�^�8�D3[��"~�i�Y�H1`���:�c���?�����x�I>E�4K
0qg����,U���B�iC�S!�$0/4E� ��q��p׮�,38��d:��鋃@���e憴|P�5�p�_7J�>�l���$�I�>�Bl����ǟ���՟���9�uW�5FF�g@���SP 	5���!1E���*T�E�S�ݪc�Ƹ*�t�`WF����/	6"�� \��k�2���Ɵ8)�� �r��$s��9�a��J���i��%�ܴ"�6͓"7�L�W�F��F��6�֨8w�p�'�V�+��azBD6r�,l��Jrp���Őx��"N�j�(���30�H��OoBG)��|�L>�bER%�
mz�c
(����]�P^\¤�P'�?!���?������O��$i>YaRnM�t��`���͉=����۸@L�/1\}@���6Yr=F�� ?��uqc�+-�� �S�T��!�
�?��e:�o(��U�'�uɠ������'Φ���~���BH�LT�;��ܞ 'XU	2�i���D1��]��i�G^~�����י����&�z�� #����h����Yl���'�7��O���?�G�i���';�	#K��@H�jS'��r���&+��
E2�'�b�W�r����C��; &7��O(���!^�t�׊R�ҕ��Ā��=9uE�2rJ��`�
c>=2��Vt�� X��w/� 4�&ړ�̡�'�2�^ܪ���zV��ܪT(wD�Ŧ���h�ß(��gyR�' r+-@n�Svŝ��~|�q	!L�"6�25�Y�`7�D��4����'sn� �p ވq�Dٵ�@+U)L�¤P�Ի�D)�M���?��:"i��?��!ʭ1��ff�����W�g\9)P�i�Pa���!l�<yz���6`6��P0�����ݎO{�Ġ�kG���"D ,x�����v�0FC'�3�k��u|��L�,�т�|b�=��a�	4:�BH ׆���?�P��۟`9K>E���pyq*�L�3u�lQ�);^!��XO��$aWeǠiI�ӄ�<��O��ĐB����i����+��E�I+�	J%KS���7��O���ؔG��u�s��O���O�����K����*�f�� �"��`@�[�����<�$�@�R�>p�yB�%3*��3�Z�U� �A�F!�1�a�
�v�Qs��9����/�Q�0��N� �&�����2�ЦkӪ����5���Hܦ	Q/��Iן��I�Ҽ�Ѯ˿n���Ę�+�hq'���	-4��*F�F�=&�A�ER4b.`6-_Ԧ���4���*�����H&0�AN%Z4,hE��"N(�$�!`���D�O����O�4�;�?A�������M�� �ړ[���$�6kx�yS�A% .�%�띴f���a֟
���Gy���%2.0�h�-(���'-FbZ�K���^�*=2`@��Q7��w`Ȣ^t����+��4h�'s�����p{ ���
85�F�Z�)P�JI"�"O`�@�cB*2��0���)e�e�'lQ�S��LRE�Kf�m�F13gó>�e�i��'�}�G�vӺ�d�O��;�h�: ���]�`�r�a�;�B6�F�!2��O��$��?��k!��"�iᆯC��9�cg�*xl�#f�9�&���z(�a�I�*z�l� �K)��pxsH&(﨔�bᏬ=v��e-�/g��ɑL�7/`�H�3e�6a�@'�T�3��OG���ѫc��8[�e�(0(����0�y�&�[B�pI��$�6�b�EA����hO��|~B��4k�V�CCL���������d:"ڭ�B�Ɔ&���b`�%~둞8ss	�Q#|�s����2D����d�.=o����@!u���	�;D�d�R�	fR��`'�&g[�,���$D�X�
�#�L	����mPH�W�8D�)C�C.E�:����rQ��%D���ȂgD�)5(/q箴��`$D�H�f�K
����?t��;�!D� h&��t,�dG=P�h-�*O�i!���O`�B�#ʌ!���d"O���+ٱPi�I�EM�ZS��"O�P�dX�Xd�a�t��/l��3�"O ]�b靕w����0�A�JS��"O�I�䋑�n�N�J&HM�NL&�V"O����#�W4:4�Nĳ i��"O4-���;k��	v+��m���҄"Od)�d�.g�b�@��L�Br|�"O��#���4���� �:�l8�V"O�JV6))���/>�tp�"O�噢iX+gH� %E�> >����"OƑ �]����V�5o[�2E"ORa�Ge�!?��` ��)0I` "OV����Q�+��0�r��%�@Q�"Op ��&�:q����J�A��]�"Oj��D[%k�}��G�]ߨ��`"O�bB
�a��Ag�.7����"O^Pi4A�#Y�<ti��#�´�p"O&h��'a�f`��O@@D=��"O���5�A�D�mp����h�"O�(��L\`!@�LnBn�"OU�
R	&M!ӫM
rN�5��"O:���$�<��dLfUR�"Oph1�I9y������O�F�X�7"O���R�	'�,QZЄԶ�d�h""OA�Q�L�T�0*�s&X�1"O의0��4��)A�թ�Q��"OZ)�ש!{�t=�m5��;f"O���쒁�Y���5l��j�"ORP�#��7x��v`ĞPB|���"O^�(3�Z�8k
R��"�`w"O��
��Q7d�2�b����݉�"O� `X
�dW'O�9I&�t:�(3"Of�@�E�]�H��1��A|pD�&"O�����
z\��/a��"Ox��nЗ/���;�d6d�4�b"O�����.�x��w�  h|�<�"O\�2��d��S�)��Xd���T"ObA����#�< (��X~�h"ON�I�����⩞$��e�1"O�q���X�CI6���Ȅ"Oh��6a*`�����A��"O�X�]����p�aOC��ae"O��s"�Pa6v�4�A�7�"�	 "Ov�iu��j,j�!H�,�-�g"O����g�'p�Z���^�� "O�q��ǅ �$K��&��%�"ORtcŁ��ZJ �%F�+��y��"O�}#�b�=����Jm���� "O��p#9�t�"���W�nE�f"O�}�u�֥c��y{Ca�e�l� #"OR0�B�I�Ul�b �"�"O&�8�B��L�Ǜ$�����*OF�W���5�t�ёeÖD\�)	�'VL�k�Ƈ�;��` T��"f>�;�'~,
Gk���ν�G�f@ �'��H#�(K)[r��ؗ�̈́==0i	�'f��D�M1'���g�/oL]��'/b��OC8p�)� *n�P�'��R�P��A{�K���i��'4���P�$>L�E)��|�#�'�8ً�<c�z��o��I�',��H4�ѲL�pB�܈W�Ƥ{�'ЈI��^0�� ���~��ف
�'�����^�hN(������sk�\��')N��!gI6cf��A�3p���'��a%g�;F�4H!F(��	Z�'���:��<R�D��EL�	��'�
$�["u������<S�lY�'jbP��N�s4{D��ĕ$��C��3h4.�A�#�p�K�K��%��C�		�*�P�J�q'�B��T�zB�	. �X{�L�T���&�Q�O��B�	�:��p"w�_�_�fjb�Sh8B�IQ�X��#�	�0�XѠ�j���RB�	�yw(-Y�`�
�4�sO�p��B���Ɯ;�[()U$р��@�Q&�B�I�l�)��Ό�$�ꆉΩb�C䉵l��Q�� j^ x9��P�8j�C�k)vQ�+ϰ(�����B�I;v'x���*��2�����<�B�I'�H�т8������)
�C䉾0}囇jB�4LH񀶩��Y	hB䉲-�����>�j�sS�΄u�BB�Iv��t���������./(HB䉢1�F �Wk 1����� #�B�	@e���#�	�h��y��IC�B䉷F���Rq��~s\����G�1��B�I8~�ɓq�@*���u�B�I�N�n�I7l[������Ϸ��C䉬R�� ��r�P������C��(yp�� r����p���J�Y�ZB�ɂ^�����)j�R����M�B�XB�ɚt��+�-Ӧ$�6����# FB�		��}9��# �P���ÒDh�C�5"s��Q�h�0`�r!ĝ �!�� �}"��['*Y�3C耜Ty2��c"O�]��]�cq�x�6΄5Rs���"O�: ���G��m�q�="f�D�a"ORX�g'֑vN���� \�D3�"Oz�6�VkjT�@"�%d�j	 p"O�����B1��c���6~�~tt"O���``��C��ʄS�$Q�F"O,�7��)d|�l�bC�<����"O�YK�E�F�ik�� 1U�X�2"O�)��GV�}�C��s��`{"O@���>pax�)*�|""O��yU�׏k���'�Ê>4�}��'m� �ڗGA�4C�h��~L0\�'_D�%�Fcr����0#�t�
�'$&�q	��::=R!��X<
�'@D/���懖��yv��<�yR��,6�4I�F�ؑJ���BȤ�y�.�1T:@�J��<�6��!��8�y��$V6l��b��3�:,��!���y" E/EZt����&y;��20N�!�y�пZ��s&,[6j��)(o�[�<a�mT>d$8*��{�!q2fXk�<��KҜ5F�cle�����h�<��M�/6�	�Å(u���@c�<a�#S��RgL�g��aR��Fb�<�s(�2UQ�J@�V:{��z �C�<��":8|��v�ڵNt�S4jy�<�4��Q��-q�̚�OLݘ�*�x�<�С�.6�l��g�ؼnY~zRgMn�<I��&M�\�G�[�q2r��i�<��F��ԹB¯4~��*���d�<9t���;�$��f�қ7�v����Y�<i6F�8f�lpf�'o��e��T�<q6'��Y���@�@�Ht8�D@R�<i�@Ё-���2EɆ*�:�{�al�<�p�ȳ{ȄXj��5(�1�6��e�<�S�3ݨ@ �� }�d-ӕ �l�<	f�U�kmT�;�&k^�Ę^_�<yW&���Ѝ��hp�l���X�<��A�7P*e��	L<Vb]�g�P�<-�xx����l��GeYt��H�ȓY�(��`сx_^L��nƗv��1�ȓgW�2�DRwȸ	%�
�_����ȓn,�R���y�Р� )�/o��Іȓ��03u)�4n��BP8����<�:7gb�Q�'�p�Ω��Z��@�����k�8�BP*�-8P"	�ȓZ��%�B�[!b@j�C�&8��-��S�9iCʎ� �|�V*$M�4��݁��B��"5#\K���6��:ꔧc�ȣ@K<<��ȓl�#��G�NxM[���s@I��;2���E۫0�|����^[O�y�ȓ;n(�� �q��m&�{����x&6jQL�3����bx��ȓaIl�A!'ʱb���ȧ�ʉwv���0�t�k�_A-B�X���>Մȓn?���G��A����B�(Z9�`�ȓm%Τ�+	|5:2f�W#=����X��`�'�V4����8�쁇�-��9�*�&�����Ͼ������m����]��`�	&x򖨄�e�CR���&�9V�>9��hd�GM �+T�Ls�˻s�0-��S�? ���0ΊI�PdF�<����"O�-� l�P�(��BE�)Ǆ�p"O@D��f$qT6��&���F*.S�"Oz�� ��+q&�0a!�U#B( ��v"O�X�)GC��*�A��5+�/�y⨝�1�"�4��?�f��p��/�y�"$L�Kɣ
�������y�D�1�F]r��#8y���c�F!�y§Z�J�tPtI�04@� k �H2�y҆�?b\Ih��'���aPi���y"��b-���b�U�#3��ss��yBE�2ƶ�;"�W�\8�@�r	Ӣ�y�%60�×��4��t(�=�y�'���ăS�f�x�E1�y�� )<AeO�G��p�tJ�3�yr,ݓd禜S�@;|�X�r�đ��y��ۼ[��trN��q쨃WI�*�y��ǩs�l��4'��rƞ���ɡ�y��Z8�1� ��dk��I�Ý?�y�%(�عP2���|P����yR�:$�b�P�F�9]RL�Q�O�y��"0�nUB7�L�8s�+�͚3�y2��8�j����X(�`�x!I��y��ؑ#�����U��\�$H<�yҧӐ;e6���V��z�{@Ø�y�i�B�2�2Q��h�݋0+�'�yR�o$"����[8ފ �C!�yrȘ.<t%���� މa BV���$ٌ(�J0�8fHϑ���`��C�����	zivhD�<D���� ��	<]R0�M�i��r2-<D��C�4Z�$���gK�`�BH���:D�0KbmK�5�h� #����Sl,D��Jd ��y�t�G�Vj k��?D� ˰�P�1t+�)H$E,�)��0D����H:p��U��C40:�xA�#D�Ĭ�
(2\��E�s������yR-'<��P@���.`��b��y�dΥ
�P�B�-]�*����	+�y��u��){��L����RV �6�y�� f����e��}f�Wϝ��y�EFl��FnZ5V�
��V���yb�Ű	l����b�Pr���6mQ��y�G� *D0�W�.>�bF#��y"E�z��Xp̃�/�h�����9�y�	�{.�AY <��Q�����yB؁7d$+��Y1"X���ֻ�yҩ�*�|�����(v�(A��yb
�'q#�,���'o�H��ž�y�G���kDo$>j�{�8�y"�@�i���bI*N$ @���y獐&��4�5�=lY��֯���y��'eb�aQ�іg�a#/�y�Ƙ,#B�`��+��y���y��0C�8�d�˹ ̪G�[��y��,'-V�aW��.|�f+���7�y�oB\u)s��t*�!�!��yҧ�1#lN�`l�p蘐�C���y���U�(��T$B�b���c���y�B1���(�5W2]1�	��y�h۫-�&Ă�Q1S�f� ���y�hu�vh������5�q���yR��;�0��E�{M���@�S�yr�T����� ��u<:�z��y�@�	�5��-��>t���ɟ�y
�  yi�2p͸�̄]�*!�w"O������7@��� X�@�6��6"O\�䍘>yl�����Ԉϖ��D"O��b�cG�s;�}aDK��af��"O$d�Հ�)���Q#JI[��:�"O�h�Sƛ5h�Lx�MeXTQ�"O����邡?9ZB�Ϝt���"O��!�.�bQa�a��:U��2p"O�}�e�q�ؘrp�Ϧhd����"O���J3yᆤ3QN�	7Lr�"O|l��*��	|� &�:<ڽS6"O<m�b(��$�V�P#�5(Xe"O下ա_�E������'-rA��"Oz�[��h�b� `��{,s"O��c�KX���*!/��_�!3"O�5�A�!�<�ԃH�	�2L�p"OƭU����@rP��>�J��r"O����J�2,%zոE�-I�"�"O��$��\Ȍ5�u�U�CJ��"O����	#w|����?h#B�s"OT�#q��d$Y�6&1{2y�A"O
�9'L�ml�,�u��^�P��"Ot�a�ȫE}>�P�FH7`���"O:]�����INdӅR�,,2!"O2��k�x���T(�fM2�"O���#�ύ3��4��)+Q�B�R"O��J���8�h�Wo��Gz8�"O3��ˀ`V���C�T����"O��!k�l[�0�,�'D�<��'"O� �!�8_��yJ�/(�jm��"Ox����n��I�)÷M ���"O�,�����q����U�t"O:��Rg%��9A 'u3�Qď/D�p�c
O49�����' �"�Ľ�`-D��"6ʅ��dI�C�ߺy��m�b�+D�`*$ʡC^��ccO��7d���E5D�P�PM4DaZ�㧠w�>�#�h2D�H��/��,�n�I1Ǟ�wH��0D����X�vr��&J�7H�a4&.D�$�7BZE4�,�#��Se��HfG6�I�\MQ����#��/z�Hk�n͵*�n�X�"O\\hv+],&'*Ma�d�4(6� qw,*ʓ]��>�x���"m�;5�0t"Y�8�@؆ȓ�8A/M!��r�iA3�phFIzӞC�iiI�&�y�~hʃ�ʪ�P���"O�����ÿR����%ōz�h��"O�+��ǒ3
�X'�^�d���"O�X�d�&y�@�ZB�Ʃ(�l4P�"O��ѱ#1Z�J�z0a%��t1S"Or���
\o���i7��(�  @"O�!��G�_�,���!����p"O�u���=��Ms��ͯ7��M��"O�����-Lc|��QbE7 �<�a�"OJ���@,
�R6�V.a��7D��V��j,Љz�.ǹ~��c�g4D�|;�ɵC�5�C*������0D�0��fH�
AK��%x�1g V0Xo!��B���1�E� 1]xx��@�4g!���[�D��@OՊK�D�!�V9G`!�dM�|w<%�p��05f�x����I!�D]#i�f0z��
U������r!��T���u�\���PS�`��[�!�H�wy�({�aȝe �<c5%��!�`.1�Ȍ�D�$(z�4"x!�� p��������{�&��`��}C�"OL��b�.H� As�S�s}^�� "O��4H�/u�z%hgA���z� �"O��zT-FAƌ��\ºlbU�.�yB�ǔsT�s`kXMze�����y"��=NX���ʍ�g� J �҄�y�'a�,�
S�J�Zj�P@L*�yBWGUH�ZS.E�$��H��_��yb�ȩ&�`�)�.D�"͖���=�A�V�I5zv|ȸP��|��J��B�	�5N�:GA�< za
6@T�[O�c�h���<�S�ӻe�ă�+;���S�#�lC�	���!ba@N�ZD&RѧљR^���$�k���Di	h�
ȉ8L�!tAuNC�	T�Ar@K�*�.�C ��R@7�=������y���°`�31`��#%Si�a{��B�a2�˩O@�3��9e�(��d�@G\��f"O�0�q��.8�dzĄ�)�t�Zv���Zö�
çw�`-��,�2�$pcD\�K��t�ȓFV�Ht�
*B��['© ��zc��^���h��D�=X���є��F�by�u(V�:N!��@�+	h�a`(˗�TC�W�R��f
O�љ�Kӈ 'd �af��Kc����',1O�અ�S�\��׻�:��'"O.S��(����sɉ1�`�������(O�O���bde+�.,�,�0c�"h!�'�	���.y&� �HW�U��`HVǐ���'xP#}�'��sC�N�p�(���'O�B���'g.e Wh�X��ՠ�(B)I\���4=��7�=�On�1�C�0/ޱ*��<o�6�
C�'���F0�e�A+�&e`�%X"ܸU��X(hh�ꎛH�P𻦇��P�NA��[���$�'�A�A"�v�Ą�ȓd�"`��j�IZv�-YCf��� "D���gd��>��}	0�7.��d!D�H�O�����s�`�-��Ds#a3D�D��ǒ�];n�4�M���$qХ,D�DhWM�A��H�EΘ�k���)D�L8wj͒>�����T�=��q£�"D��s�� }�TX��>��!�@�"D���
��*L@��t"���p#d�;D���!�J8�U#����7��pSҭ8D�8��20H�a�E��| w�4D�hzpN��I�p���$ǡ# �d�V�4D�����%\��`������6D��!�D�?]�,�8u��aJ��f4D���v�Gtި�%H�%"F���7D����̓�M3�)ˆ��u&�%�(D��K`hS9,e88��M�+jD��J#D�|�R.��`�"	����YJm��-D��S�B2"0�c�D�G�D-���'D� Q�,��ZZ44�Ջ� u�ИvC%D�t��jW
s�U����-k!�ؑ�� D� ���84
d,Q�(��O�����( D�,f�ȼk8{Љ���/+�B�	�j_z��!�1��e�e���C�I GK �r�G�=l�����'�TC�	%r���DB���A���/bs2C�4$&�I��I����1ReԎ}�C�I�Zn@��I snt�r3��/B�*C�(���W�ͯ|�F��wj/Nb�B�I+E ������<݃tf�v~!��/��0)F�C%Y����+t!��ؾJ���s�T.��5jgW�yb!�� �Iڕ��*��1'퀒kņ��"OF���;��X��K� a�"�v"Ot\�w�Δ�Nu�BJZ#7�2�5"O漊�f�/35�R��I@�hM��"Or�{waJ�V�2:�a�<��T٦"O|�xk
�����cKћ&�b��"O�=��+@�R�DS�N�L��&�/D��b���
e�YU���~i�d�8D�����K	�����vl�-ö
6D� Z$A�,&1���en��(�i ��.D�dsw�؂=����q��
p�z�)��-D�@�GF$Z�lᶯ3@�	��*D��[CL
�5j؞9p����)D�,�!��
6�YS�4w\U�)D��Zc��^��D�3:� �gk(D�����4	�r��t���(�����/(D���V����!L]=�pLcu�'D�̋ �R4.Yp�� B??��!D����`ʲ�Z�Z��/Z��]0P!D��q�N�11�t�v'�����e2D�@Ho�)��:���X���9��B�I*h�܈�&�J��l��AH�R:�C�I�GVdp��Kk8E0bD!��C�I�p��(�AY�{20���,4C�ɡ^<����ʌ�,��u
Q"[�Z�@B�ɷ(�P9����5���P�A�H(&B��~��XO��<���s�{��C䉽L1>yj�.B�c�b�S��RC��C�	�NZN��f�I�A��V)j*�C�I�L(����Z�0X�@)�����B�	�^�̹�D�*�x���$g~�B�ɀ3�����CR<�b$��!\�B�I.S��   �O�_�h�W��G��Ĉv�m�<��ͽ�P���ELv��3$"�N�<9��
��(A�u����G#�v�<�w��3ªMyu�K�ۢ��)s�<q�a�2v��o_k@=�GHg�<�DeW�0:!�4�B��[ePh�<���	1|��k��J
a��H���b�<��@Üz����,ʜI)o�y�<�vO�-C�p�Xe��|b�����k�<�Η.lr�p�G�t�Y�bb�B�<a��@���1�O���%S� s�<)�(��#mҲ2����ȅr�<�Տew*�IBC�M�#Z$ȓg�����ib��Tl��4$����:�,y��A��\�wIG�f4-�ȓk?X�����XNƽ�sDM�&��̅ȓW����&7|@�( /�?���ȓR�f�4�L.D[��𔬃�C6�,��ҨH9�e�����3��#?��e��ؕD��+k�� bM )[u^�a"O� F73h�����2or8I"3"O`��Ԭ�&tIpL�ǈ�B$��-�!򤍓[��a�ɖ�k{���dE!�1z���B��
�<Rr�ZM�!�Қ9��0��!�7Yk��â%�!�$���� R�̜�Đ`7��((@!� ����f�N7 ٘ax#�ENX!���$?�l�Z@�׾C�T�a��9G!�$$@��K�=��={�I^�@�!�D�K�,�@�����vX"#8�!�� :�ǅ�tD�(P���!4�R�"O��#v�0>��钣�K�T�*�"O�����K���YH`bQ8q���a5"O���Q�u	��5Jz��!"OP(d��RF@���?Ey����"ODx��`��q�� @Fm\-WrԨC�"O�U(4��	xYL�烕bo���3"O@5H1F;s�>�[!��g�8��"Oڙ�#ŝ� (H���SO�ɓC"O�t��^%K�]��]�b�M��"O^�*bOD
�\�r��.\���s"OF�C��Cxap2 ڃ4Zp��"O�<H1G��GA(U����⦐B�"O��	6��|�y��-ϢX���ӄ"O����eɣs�nP��+1����3"O.5���p�$��bCE~m,D��"Od<+Tn�q_t��@ٯSQ�e"Oҹ�v*ݵ�T0r �U3�d��"O�M�2GL����i���%���"O�pǥɷ91���� ١�N�С"On��u`�&[���0��J�`Ӛ��"O\�4CF�@$I�9�a�"O�	�plV^&`����$�R��3"O��3'�>p��,�db��S�^��"Oj��4�H�8$,�Bb�X�,��"O�u0#��!�H�d��m�Q�"O֤a_��� ܪ4�R�e���y2:�HsDޒ&vd�z� 
�y�lR�v7�|�J\�"
�r��>�y2�]�X�.�����g�N)����yr�=��g٧[�P����&�y�GM�{�d�$���>�f�3 (�;�yY<��T��%�61&xx�T��&�y�fC�d	�a��9%$KS��-�y�ɰv��(��� ������y�!E;X���*�.sj]����yROȊx� C�$Śs����J5�yr�O�X�f�I0LLi�F� ����y�I��\\p��a�L隇��3�y��R@��P/���qoQ��yr&N�*$�J"�^�{������D��yoZ��b�!�Ül}� ؑ�P��yr_�I�|[��P6,$u3"/�yF΁t���b��*(�v�bQ��y���	��\[���,�j,�q���y��D0CVmZ#�"B�B�B0�yBm�.8�-#!���r��P��	�y��ԋ"�|5�h�0pL� �ð�yB��,-$ �`�\Dd!`����y�	Y����.�3@���y��B))R��⏍ 2�)��-��y�!L�m]���+��-a�߿�y���� u��T�?$�(��Bҍ�yBG�B�P�y��F�g�NY0r'���y2"F+�ș� m5�Q`1.�y2ņ�d��8s�L�<a�|4kU�Q��ybF@�i��y���	-l�>xhR,��y���z�\�Jb�RcA��SG�_��y�(GP�,'��m|躶�B��y2��SK� c�B�3�Rx*���7�yBġ>�<h(���#*|���
��yhV�O
�Ф�܀�p�`V�M��y��{X�B� P���(���y"�[+�b��&���
�*ե���y
� ��E*#�t��N��*�h"O:�����&R *��(G�:|Qg"Ov����9�\A#n�)A[�i[�"O�L��f�=6��r���1x<�"O��8�ͅ�%�f�RS�F�G�� ��'<l9G�D.6`� �WD�c�0�`�'���5k۴N�\ڇ��?M�&8�'�R��b`ؾ�A�DLC�v	��'����pz*%��c��?����'  l��e��X�,se�������'�Ꜹ�=!5�t9��>�0ĳ�'�긺1���9D�1��=z:���'�A��">t�M�%��t��'r>�iE��	�:t��f��gH�c�'8`y�W%�D���:�!9L ��'[L�u�G�Q�l�:���[���Z�'�~$��C�<""��p�
iOxa	�'9�)C �ZAd� �@/9a�2� 
�'Ȩt��"':e���fx`4�
�'��%��O�$+�
� ��7e
���'y�����h����עH
jc�	i�'��0aǭF��.L��ٖi�|�
�'W� ��'&b�e[�ٖ{zy
�'n�y��[E�T�ALH�vJ�dc	�'A��huh��Gy�L�Ь(s���S�'���1.���!R�dܚ4ḠR�'���C���E������W+ў��'��@�AOgy��+�n�� !�'�T��be
7G��1�
I?[1<�p�<�b枼	��) ��KG�����a�<�f��Cc��Kd
,q���I�IRU�<��D�.��[����^02��R�<��Ǻ	*@��b�HF�+�eK�<!a��t�J���J;���h��LH�<)���yWV-2va�=p�� `d�L�<���&^�.X�Roi���hvf�H�<�W-�&{/���ҏV5:���Im�<�O� @@p:�+C�n���P
_�<	u�,N��d�3HW�Z��d�<��
��1�u� ��18p 0 U�<iG!2��5ķCLy��.�N�<	2��RZ½���s.�\�Vc�N�<)��#و	"�Y�)&u��	�r�<A�jS	�l`���1 �B��"OIp�< ٮ&�mB�*W�0G$H�vo�<�"�ޗ�hٶ'ףH�p��#�A�<A����WRV9;��ya�,QV��t�<9�D�2��(�Ac��@A�o�<��!@�;��|��HG�,��F�d�<c��J�L` A�t�lqS��Yk�<q�@�*1:z�!�c��)���d��A�<)T�B�H�di����,1��I�T�L}�<IGœZ��5����tM��΋v�<q3��wN�C�F�� 4�����p�<��٪s��M��E^+Zň�!C� H�<!c�\g��)1�^#@��,	G�<��A��|�T<Xd&��S{P��dnWj�<�bk˘��@�ʗNga���f�<i�e÷J�h��K>�ttAn�n�<!��'/��AGN�h��x�Cf�<�YRV-���T���8�DG1��B�	=Pք�0N�x����iĵ]e�C�	,����:̘���vC�	 J�0(��Z1{��|����1l=C�)� ms��½70�,ar-��Y3�x�0�i�ў"~nZ�E+
X����6��� ��I�.��D!�I6<����L;Ѭ]Z �u��B䉗[���Z� 2Xr�A��e�ڢ?ٍ���oτ�g)�b��X�Y6n!�W�K4>� a'�E��`Be�ob!���)voD0� � X}��E#��DEa��O�d0�*�>vD�`i�g�g/��H�"O"lʰ!�,5􌡓h\�^�"�h�"O�0� ,_�-��(!��.\�t�+�"O�8��,� ]hY�
�"Д����p�O�n��֠���t�0Ѓ	g�b��N>�	�ca��È��H(Y hD�I�|���u�b�2��#0��RҤ��BJ�0��6�`���͎9괵��X)7z�O���D5">�p�͎+Sp:q��Xt�	N���R}"$[�6�.�Hw*R�'��O���yr��2
��5"V����jF��'a{�Ği�!1�矛*݀=��C���=��4=��\�f��1y��!8��<�L�$�?��O��餉�5h�@p�Q��='Z���	�'n��9(	�Fh:��`�I=�4��4�hO?7mH:�P�,В&�!�!S�J
!�O�Q�2q�C�V����y����!�d�&y&2�-��G�P48��@ N�O��=%>�PH�%��s��X�F�5�0H)D�����ǻm����e�W#Q��� �&}?Ot��.�D7�I%Ж}���G�D]p�(��G�g3!��s۴)��@l>lT�����-1O��	R8�x��� f�:uz��G<=�|	��5�H��D-���&K%���x��@�U��6mi<�����Ɣ��"�\��R�D8�,�X���O0�ʖ�[���A&	�.d�b���"O ���n�={��{�bN�%�������h���	��+x��Z6}Z��s�&=��~RZ�8�I�F�,�P�!~���(�%���'u�i�]E{�CM��V	q��:k��q4&�0$!�
�M�`�I+� u�~]Q�b^�)�X�	
��?��j�H{v�8Q`�(s�za�2��v�<�v�O�5��D��ʕ"5��|�Qe�G�<A�!ӗBn� �!��I�Z���@En~b�[8�((�ذlmTe� O�i��� �5D�pK��^1�蔃���Z&�1�$!3D���Ě1�"�����{ V�fβ<��y�H�G�O8P��@n�z#�e�%��M��my�'��T@�Ǫ7C�[wI_�Gt����'{<�I@eՙ�&]Q��
�v�J)�H<�	�K���ba�BJ��1F�[9U��'���ڃ�I~�'n�`A-�䠡���<�^(��y7�s�S��@D���d��<��OB,��	���<���6]nP񕌉�?�4#>Wc?�( �\ba�Blhܬ�weӵ`���ȓ�B5�Vg�$���&Lb�Gz�'��`jDT�B���$8B�R`RJ<Q�D�9�KF�����!���)�nz?I1K\+��=�
����&(�T�(]iiBP�<Ar�����X��V��)�5�J�<�Â�
�xp��=�1V+G�'YX4D�4lɨr�f=��.�^}p����
�M��'�*!CdF�Wv�5L������hO�py�)�{R�2�*��g�. P"O.Pa#��:'���P)ƿT�.0��i�ў"~n��;�Y�N��)�,�G� F��B䉷^�`H�윤Wg�=�!� ���p?� `=�5KN�y֮��7M�r�5�D"O�a�N� %�x�P��>}IJ�y�"O��ٖ�Mi�2H�9�yJ�"Oܝ�E�mS8���k���Y��"O��ȧ������@��T�*a�8f"OX����9%�<B ,��>V��Y�"O�uK��L<p���G+�1L,l؆�D�O��$��aj��0����V;""�|�ӓ��']�tځ��T�N�k'KC2(����'�ll�s�:!�J���⍨ ��l�H)��h���§j?��P@�81Ҵ��5
�t9!�䈾t{켛�ቫ?q*����K6�viϝwh�~�����R5j��%��Х���=�����ɩ|��,�P�#����t	>�*"?i��I�:i4���m�l�RȐ0��!�6Z�8���f�Y�b���!��]��T���Т'S�@H��nўą�ɛ.�(��(	x�!C��*7I�B�I���1��2zx��pfƶ>��@�C�'$�'Z�dF
�`|�`U�ȆJn 7��~��2hld@�V	̘@+t��!��=�S�O�����S��PX�
;Ŵ�j��d)�'|?&E�C��@�j�"u慗1��1�<�ߓx�4y����CZ�+A��Xل�In�����R+|1�������e��pl�{(<� ��e]�k���2ȵ�`ΖA�<�������Ć|J����!�t�<��(�v3�H1�mʯ&��fiV�<5��/�t�z�N-4��)��
~�<ٕ�TU����g��h`�)��Ma�<if.ĵYAl��۰G"�%P��y��kl����A6��Q@I&�?9�'���SGg��Rq���N'���'C�V�� 0}"���K�������~��6s
,�� I�R��S`��y�$��&*�8[q"Br�0�����O��~��,=l���ݟ:�9�f(�|�<�P�
0*��HZ%f�PF$Z6bC`�'}�?A���p�0��D�W�L���"O.D�8� �u�
���� a���`�-D�P�sBÞ|�0"'%��� ���*D�t���z�r�P��R�}�Dʁ!gӀC������ګ}&6���@F0:�J�)	�'`��4Pڹ:���7I�
�'�@���0Y��Z�!+qVPb	�'�
d6g�1����	�3+&�s/O��dқ���bO 'BJ7�E�0K!�܂� ��q	5j�� F�+#(!�$C(fP6�E�a���vÉ*Z2!�ğ5Z���A��R�P�t� ��7!�$�O�e
�F(x���K�nT�G����3"O2i0¥��X�v��"��%��]8�"O��1�ɱN�ҹZS@C0z��h@"O<�i�/?5��q�������6"O��DA�y�xbc�C> ��0��"O�%1��L�c�)�g�B�|�m�"�'	��:�S�'��9�s@�V�Jm�'��'��=��	h}�G�HYnY�%�
Cl0pT��t�<�3��i�8|��B-ZÚ8���Uo�<fO�r����k+�����[F�<�$%�f�Lu��a�c��hر��F8��Fz¨H/[�p+3∜����p�^��y�D�$��`�'@]<:r,��	����1�O��pv+V�H�SǮ3+�`ѳD�'��)� �u�bl�?d�����/����ݢ���$lO4�r� N�g�`������*C8X�"O�)z�C!+@���@Ζ'1��)3"O�E�5���0
��k(Fq	@"O6�iah�?f�:P�ԡ�6xd�S�"O�E ��H��	*��*ff2#"O�����.94�[�ᕣk+�5"OZ-�2��1W��XF���"O�Щ����4A�r/�j� ��"O��xuJ��V�$蛵�ڷ]�2��q"O�uvEm�H�9Ei��H�e�`A:D�� ��"�Le2�@G�C2����6D�0AqiG�(�>m`≟�it�}j"�9D�L�g��Q��\-*�:U�6D�@��,m����ř?N�,���1D�ؑweɔoɾ�o&4��Z��.D��"��ϊY{�@kP�S9�|�q� D�X�2��/i��M�����*�>ш��<D�T�0'�<`_6ȑ�ž]2�*�:D���!�3c	��� k��RN��5
7D�h��L���C%���썈�0D�,�F���rHŲ-n�уt�\^�<��FS�hR��5i��$z �KO�<Q@%
�T�)7L� iHt���A�<��?"e�0�,@�$I@���{�<I�"U���%3H�P[��[`�<a��\6 �����꟨8J�ty�L�@�<�W�	�Ya/A����s��~�<-Ґ�3�	a��uA��C�Y�J5�ȓh� "s��zv��E��
hV��ȓ*��A�e([3z8�Xqt�	3�T���.!~�k��۳E!��AF��]��& DX�F�Ѩ����3F&�@�ȓD�q2�H����0�L*<hD��hRn)ZQbȒ+�ix�`;�^���"np[G��/ �Hy�2ɓ�\�������,�cZ-��Г�C>+���S�*�<��B�� >��*a�ų&�(53'�o��C䉩)Sa�ԩ[�,A�!i�v��B��0�[�H��|Ԑ��?��B�	�p~>����=?$�Cl�sӒB�	  V`����ڤoTH
v!	+JxB�	�e�b��0mB�$t��ϒS(B�I�^`2���.I�{�*���C�356B�I�*0%�;\�P��obJ$�� ~�И fH3��yСM�#�L���H�n�
�&T�p h�n��(�ȓ]��ѣp(Y�
6�%8DH
�E�ȓL�����Ցڪػ��˫!��ȓttD�%K<,S� 9���33	��ReX��$��1.�"���O�x�ȓ^LL�BH�[O� �4ٖ��ȓ�t�Jh��t����T����X��!�^�1�*��@<�I��p�U�ȓZQ*t���)4 483�k�$��Ev�X���ޥXB��Õ.��fхȓG<�����Sd�y�Wb>�Ȅȓ{0�K���#t]@�c�`�$JƂ��ȓ3�����x.��g ։%[P(��9il�Pa��Bh��
I�!��|�����1�\9s�^8�s��F�HL�ȓ}�B�В�N�jf��G�\?c���ȓ�x�i��Ԫ0��q���7P��x�ȓ����F��~B�|{G��j��P��S�? �h$��>��2���E^�0�"O�4`��^�}.��鷤ԗX�l��"O�Q�@��h�����œ[�H��"O��Rg ���4Pe�U�-��ʴ"O��s�-Y	,���f�fa�١�"O�M�q�K�C%�����zR�"O@б3A��"�&��.�eb���"OT� ��d�@���J�_�8�Rd"O$ r��U�/Y}���J��"M0�"O�)��ޒjd�9���.4�.�s�"O��rd,K3Yz0}�6�=>�j1�"O��a���<�IQ0B�\�µ��"O$<�r�,~�r�����e7��RQ"O��5k?drР�P�"�xj@*O2tX���rP��l"�ib�'��5[�?;���&B�$1���'�\0�HĒ�l�&��9x��'<�;3*Y�R;�QV��9?�A�'��1 B �vbPGز	�>���'(�-!�h� 5�5ї�ֆ	X��@�'��Ż�A\Y���'�3xP��'�D � ��*$9�q*���M"�'*�}(	f¦e�ф�/�&Y�'�P��e(`RLdу��R�'��$3�ڶf���	Q��vb��Q
�'"8���a^�{S`��N�e�=��'ۀP#Bhs��d8�j�Y�ĝ�'
���p�:*ǀp���c��2	�'�s�&���@*Ha�PkX��y���(q�L��jO�5��<J��� �y��Plh�Τф���\/�y�&�Dn:�3�,�)d]{r@���y�
d�L=��ʃ+O�iz�'��y��+I��[�͚D���ȑ��
�yB�W/J�x���9i�Y�iB�yr��9_\\��UŃ�3����aÙ������:YW>�O?�$Y;*d�٤!�\��]I�dK#1~!��H'dQ��j���dq��	��ވXm���bF'�p=٣��-0і]���L��y m�l����D�\�֨���ҭ^|�k3�7nd `����_�vU��Wl���͘�79t�C�C�7~s$$�?醯���� xA�0��>u!r��4�Sb�/<��,���'��x���{�S�O��{�x�P`p��ǈ;��0'��X��OćJ�I\��~�N�	dpI]���GJ�H��ȮO��B�#�:P�����2.I&oP% ��3�k�N�C��a��9�� �qO�a�f\ _��h���le�X���+�5�m�n�A����ę�,�^	pt��v4�S��P�+���ʔ'��7��6aO|�ɱ6��;6�>Ps%���)}R�B޼�DC@PO>U�Q�\�1�Q���l�K~��u��1��l�L~��)7�j�@�(?�^�����	>l�`Hd
F%�x��a(��M���I�Zx�+�`]�45날��%��m��e�?�=bs��<��'_�7hL����'�����:Mw�<� ��W̨]���O�}�g����rӓj#�!��I�RP�c�-M�2,�x���Ѱ�140����>���A�X�HU8��5eȐ�"�jP�$Y���S��Й�P^J��b'���M��_"n(!�5���)u�0��ځ��lV�Da�7(�D�E#��Im 󎝞%|m��LK�\��%��%3�~r��t}�\�튈	^��K� ��]*$��.Ѱ���aD��|�O�u)a�"��O�  K��0�Bհd���	�c
����X�.R�
N|2��@'FE�RDY������/U?�`�$�����$LOЄ8� M�/�2��O6.�ၲi��!���r���B�yJ~ڐ�B�=0H�1!*�-0'ș�B[�x@��Wȁ�g�*B�	 ~.�qQ.C}T�	�(^	LH��ɜ�4���2�����"{�V�q�NL�� �<�K�Mݑ�fA���Z�c����D�4ʤa�h�&�2��l*����DW%V/�ar���+�N�
Z,=Bv�'=��D���?�Ґ�A����АT#�1U����?9���[y��AW�Yn1���� ��'�6F0ȳca��
�p��FQ�� ��ޜ	�PP��	�V,j�K��<���!R#D�MI�b��0%�0�3���=&1bQ$?��G.��ºiHXd����,���0��NW��(�'l�����	�^��jA�I�2���fY�4q���z���D�S+nlџ�{�!�>t�.��f��+���t�<\O��s7 
�D�.1p��\�8�h�����;J{P��X�=��C�H�|���D=TjM�Cą>zdȰ�#&��!�qOZ�1C�ߒj���2�K�&&��s��0���O��i�ȟhF��9���C`|I�'_���U�׹B2�xgI1;���e[[�l���Ҋr�:�1�cJ�OX���EI���iL(=0u�ֆW')b=��&h0���5��'B���DS���Ţ ��<�ֱ �2��,D0�D�$�M#�B�E��x�u%B
#˖�t��,c@2xcԚ>9ri�[�<�i 2o�i�"g��)�NXj4�|�S�,�Zt:DjS^y��ݦm��B�V��X��H0M�9V��;12�ҕoÈKǞ�`Z�ah�#c��81�� 5��,"W���1Q�:�ᄁ�[�8�%*M*Bj K�LC]?��ٮRkJbӀ��e�X�0�/R�f��Bb���*a� `��Y)XK�P��I$}o�D�>G�^�
2G����O�����<��H_%9�հ���ϰ�ۣ��E��U�S!ۏ^��شqy��Sh�=Ou>��]�B�YQGg�&e!5N��U|�� 1 f䍺��DҖP�
t`��ѭ&,[ƾ~�Po@�R2��@��z��S�a���:�Z�10I�V���ρ�U4O:��[c�I�S������J�*�v���҆x��$�_�}��	?z�"�TA/���y�"M�'HCaST�@�з
N�@�&
9�H���qM� �؀&k��F��L��ѵ��3̆�2Q!�5\5^��T/۞_i���,i��#+O��֫��;c����m�r�H�wT�m%�A����2��b�#�'��b�oΔ�G}���/�(��A�^�z9��x�FOQ��9�b��k�����dn�4	U������x:��h�O��-���m��聧�m�|>Դ�؀�ӰG��G}�h�d����	Z�O1X�a/I��1@�Y:-	�''���d.�����Ӓa5R�:1b�o�R҇d�];�8�D�2�R����Es?ɱ�5!�����֖��~B�����-�f���"��G��g����$���7M�s��X�{��iR�$f����Μ�ڥl�mA*O��L�i���;�ə2�| �=�;l;̠P0E�g���4--?z܆���Z�|�i�· �:Up�����8���Q�v���'�LI"�*�*E�k2�RT4f�����ܫu����)�0 K���H���M�aE�a޾B�I�F�-�f�G-"�� ;�i�;O����Ц@�41�'A�:� '�0��#�=B�ʡ�	�'��`+�ˬ#����������$�����v�?�'	��R�	� 2�d�Ԥ.y|e��M~
�I9 �P��FL�#�dP��g�l���>����OPx��#��R�2��CB.Z�t�"OP1{r��8�  #b��2��y��'e� K!C�4$ް��I56���r.�V�"���:+�(��dB(b���ӂh�MS��	g�Y���n�
�Rq��a�<i2`�/[~  �'C=h�H����J�Tq,�0!�A�\��"}��&�Z��`9׌��*� 
Fo�|�<1a��J���Y3D��ة�L�������7A��h���	d(@�[VA�-R� $��7	!��{׼朢`=P��"O4e�RM�Ek�J���O؞�R��ӤW��M ¦�}�088��:|OH����C`��Zڴ0l�����Qr5#S�F=;�b��}�S�������8pd�Fx���Z�8p��#ʍ�t�/r� C�+�;.C�ɽ$�� ���f[a��h@�}���CH�#y��"~�ɍ�8��2,

5�X�!Aۡ:Q�C�ɝxr(󗳤i����n�w"O��3q���c�L1��m�D�0Y�"O~���GX>�����2)�䜻3"O��2)C#_�����^q����'�T#4%R�A��;'	�3yrpAy�hɬQr@�Ɠd�\lP�#ϙ�l�Zd/ӎY�"�F}�Ň'=��y���*!SƑ�'����d���Ѵ[!�d�O鬡R@��8:Ac!GM�*��䚚"���㐴��)�'B��D@��a6���.��/�r`��Z��X� �
o�F�1!�2}H<<�'�� ��`��p��ɯ���9�O��?z="��֙#�Z����i�f�h�����\8������Łu`�m�	��� �\��`���d��͟E�����	�h��Q-�q�>M"b�;$�BD�m�_�̱��"O@��J�;��0%,�1�x�j<O��Kq�U�- K�"~�RB?	"4\���35�jk�̋m�<	��ʼzO:4A奆�C��A�v�Fl~�J�'�L)� m^M8�<
��t�
���n��%n|Eqo4�O���W
�1<8��H�=&$8T���Y��Mp�j��Px�=?����WZ�S/�:���˨Ox�ӳL�>~7�c?�;d'1eP�@��B�V|�$@3D�|�T�Y6/�V�j1�_�o+���ƪ>���֋H�@�"}zr��[��� ��ûj�����I�L�<��X�jp�bcD� ��Tk�s�<)�B˙h�2�k!	��'�p�!Ro�<���G+mJ�p��,c�Q'&�A�<9Q̬,P�3�)��

4T��f�A�< ��Aq�I釥�9e�@<��f
|�<�0��cڪ��a�Զ[�`̈�}�<�ѡ6M��CK�e�F���mu�<9u����]�w$�/G� g�k�<I��_���0�]-$�DhxB#�k�<qc�
���jjA.e�n�XDnX`�<���ۻH����u
�n,�p�o�c�<A%P�tp�m�/D�����Tq�<IP�� D��C�,�"o�)����m�<	��7�8��ܠT�Zi)��Yj�<� 'e����+�H-�-a�G�x�<��N�(B⹹�&�8b��@�FQ�<��E:��p
0�ȯl����Nu�<�wI�y���D$Ez$�@��r�<��J�:,�6y`�,� ��Ey��ZA�<A�I�I�x� �G��@m,�h��g�<�+�;
�L��%��=A�� s�b�<����B��`A��[������X�<���@�j�@-���Х)q�<9�KA8	�HԂpcZ<̰��%�n�<���Lsq�e�UiM�>�	��Ck�<w _$�=냀ϵ��9�.�g�<��$�7�Xe��D�
7:M�b��_�<���4�(��$�l��P��Y�<�K>zr�@`M��7D��zT��U�<qA�Y��t�r��ڝ�ph��,�V�<��	8;H�C����v��B�Ic�j �DO�E���)����P}�C�	XWH8�&�W�g��C�G�>gVC��/~p�8�d5LpRa���ߜM��B�	zl>A��.E7�X	ˤOP�C��>!�,0��[�*U�7'�<*��B�	�Uf��ㅢ!+:	��&��/�HB�t�t��
��mR)���
C䉋8Fv\26#NVriې�W�B��"ₐ�cg�{@Ѹ��̱kt@C�	�n�`��Ƀo��\Q��/?|B�I�?o��#��Up~,iDiJ1I��B� 	��i��M�z�&�i ���B�	=�p�d+-6�n���C�T3B�I<B�j��Մ*F%��N&>P$C��;0k�KF�ųN n��D�ɭB"<C�ɋw�@��[80��$+ڭn�C�I�C!"�c"]�D����D�tl�B�Ia><�+Z&c�Hd����I�jC�	�n����BD��~�|q� 퐰d�vC�I>QB��Y�HZI2HY �j6^�@C䉸(N�S�Dm:q�Sd��!�TC䉈@�*=H+�]��sK�m0�C�)� ��@�F
��q+y-`��f"O֡ �*�$U�xu��+>��"O��@� ?SѴ�Qg�P�6xʕ�%"O ��oE3t@EJv�ݹKP���""O�$�G>z�`f�B#Y��A!"OF�VgF/<�C6��[9�`"O���$ȟV�,�i&��0e�:U�r"OV�b�!�ePȐ�#���ʶ"OR8A�ʕ*{��<p�Z;[^8��"O,5����A)~8�eH�&[[�I1�"O40C!�t��E�G��S[B�"O~��� ���(��>]����"O�i�̟U��0a��Hn=jp"O��!�)���a��%X�|8�"O qA�0�`�tD�D:L��s"O���)�9�TT;&��u,�0i�"O���$T�WXh	��L�5&����0"O�iԃX;'#dЧcv�"Oh�yr��'��X)�&"J� ��"O:�sb��c>J�"�jׅ"Kr�"O(PZ όr8}ȁhO�?<Xp�"O��Z"$	�9\x�v�٧-8l0�4"O��a璄9�veQA݈`>"�;�"O��q�cƑ �6M A!'$���"O2 ���N%E1� ��F�=��"O�j���8m갻����Qsu"O�����E���a��K��� �"ObxI1�B
�u+sϛ�S��u&"O�A��>!$����.Q�lf�$��"O�D��/X�un�\H1/��(X�a3�"Ob�"�|����/��,J��U"Ot�`�dƄ"UR\b�@N$<!�"O���"L�,Wt$"���
��*$"O0�c�)I��Q��nY��"Ojtbr�X�4��%����2*���"O ���
��n�=��&�_�\)�s"ONp�ER�@��F�E��ɋ�"O.Q��V;p��`��KM�r����"O*��.��g��Q:gA#em��r"O����ƌ�a�v0�$׸l&.��g�;~m�`�,�A�)��`�N��*!�����ōa^H���9D��*0�E�=Y<�rkżz;&L�Np�P�Ӆ�2)�\ܻ��'��D[1EZ/.@��	�}�����z��Y�7l*��LS�a"]c�Y����f���yB�����٪�	�+h>$qe�ʤ��'�M�Tω-.&u�u�ӑ`K��R���}�()C�̸Wz��$-d�T�ҏ{��	�.#��,��Έ��~��&*���
"O̱=�P�Q��<a���O:<��ޛMꈄ`��׊i�|�&T�hB�D�d�RH��əY��l"�$U�)�^�Ũ�.P��䏧!CJ��*��S���|Q5��Eb�h��&�-u~<1�,�&�`D�S�^?>�b�q��'��鳓��Q�(-)��(#��䚡�J�X����'߫j�H�O���w��j�Z�b2�ȯ��UѴ��=��ɕoD7A��}���	�^�<�� Y�~.(h�_H�z!0!8� X�3�r�H�}��P:�)P�})�O�%��L�O��B&��O���O	%8Y����Z����Q�J��� B�����?��&��Kl����>�w�	�d����B��V��)ؓ���~r��w���
��A^��$ ᅉ��%��i��r����~��ᑫZ��4YZ�
 ���5f���(4���7��'�`����J$�1��(�(�F�I�,��@�f��M���
G�X�b���" q��MX�MB�4AN,�%3t���aH����4d��.�m~���9U�<@�2�&1��~�	�2��Q�l��7H�#���@�hQ�E5S�H� � ��>ŀ�O����& ��O�xt�M�T�jL��jĶ�r���2�D��jҏLRP��N|�� Y��h)��	U!,0hX���q?!��H�I�� LO�X�W��,E���8���jg�'D��r� �%*�����o?%>����ڬp��D�wd��?3*\!ciҵdw��bG-O!�� 6�с+P0�lP���%(�К�B�>�Ԡ� -��qaeּ�������I�{-�n�/��M��e��E%�,���m�}�` h.��R�$ISf�+Ƥ�U�깻���#x�JE�t�V<aK�%K��>�I*���2b#�r�B�J�%L;���/�=����kI!_��b?���*��t�p���.]�7~�]s$F�>	���t�B��ד|ʺ���`��C � �L�d���	,r����3��S�'
����oyӨ=Ya�%_PT���X�6?t�R�"O@8��a3Դ�����1���X�X�Gނr��p�'���Q��#*���Z���FJ��*�FH���!�f:Yy�"�L+t��W�K�;n���G�3$�XҶ&�*Gr�U��0��k0�>�K�ސ�eȮ��O������f��5�5�ŗd>r���'4�ѓ3)U�H�0Ő��S�P�E��=;�Xq��Mӌ��'�<M�O��*$�F��]q�8T��K��$�:�@6�*LO�1;"�R�U�T�i�[�)"rԜĹ�H���Ez2�� 6؀���	g?���cM�� B��b(��Z|�O��Z�H=_r�`��	X=���iD�A25e�V�v��1�3.LE��0C�>E���C,�P�ǖ1��Xր�	v�Pa��òF�dD�6H�[Gd+��S�U��AؒkL�-  �
g��l��D_k&DQ��W9��O�]��Õ,	�&82vK�>�H� �<٫��C!f�
�K��ɇF (���ï��U����"j��J� B�"�����	L��҆�(c,hS���L�t�C�[�Z	c��N�}� H����(O^����]�Ts���ң]	&MrB�¡q��4Z��LP:�$�!��� i`���1�'��n�"Pr���R�`K0�x��1d��RUG�k���O��!C��Fe����u\�V ��1C�4�I.�Z1; �h�g��8�M{e�Y�H���s�&Y�h�"��T�$��P�0�>q��S	ؾ��%�8R)�e�p���$@����JV̘;��F�$0v���%��D�r��%qٴE���T�"!�Ӝl!3����9o�:���Y�n>���0��{ ���K�/:0��	�,�Ba����}�O(�)��
[$K1+"��rH��ਟh�)G�J0�#��Uy��iHR��D�D
�z��� ��c��͔I�4��=E��؊'��0�,�	V��cNC@����'�z0h�O�ju���O�aV�@�/~�H*i�1��K��'���֟-z�\�`.�
m��"�4x"�����U����V�J�����l$�jb1�7�+�6l���3��O�=�$)1,V*<{"���S0b���'�`��a�kb(4��%ğ8<��#�}��pƯ|�0�#�YU?F�qD��Mבּ/>�!�d�ys�, �T�/8p�T�r��P��+���E�4��'��lz���h��	1쒹�y ÕP��f��	U��a�RV:D1U-�;bT:�'��>�	�t�X��_�s.y!�ЈC�I��x��\�+L�pj�5"����W�<Hԭ)1B�5��=Y���?"��d�sF�EzZp"�GNY���s��$Ds��q��ir��{T�(�=�g.SDub�{
�'��D���6XY�L�vB13�� �B��L�نe�l�O����lw-�	v������!�'���1�O@�5��ܹ6�7[� ���o��c
*}��P����_���E
�WJ���h2T�	��� b�d5�4�|�#�߶��M@!f�p�T,�V؞�:�_�i��׆�$ �̘�c<|OzA*2�Z8̕2ڴ$�����L� /������OJ^��ȓST��b%]��2��Q�
e\ Gx2���b��P�a퓃H��Yင��N9]��&��|��C�	}������>g�8)��a	0 ϾLFz������OБ�d��6SZ}�@�L�in��"OV�GoT#S����c�;���B"O�!����\-�}�����x��"O���#��,�>9k��%%� ��"O� ���<,es!��='�P�$�'��\QM�8��c6�X�b]0d�ȅ5��U�Ɠ	A����Q+n�RE�i0�G}�?=;���O|\Q5�ѵr�<̹A����l��'a����I�T���kV����x� �'���xըZ�e̜�O?� �XDi�d���)*ի�z��"Ojd¦j�8mњe@2�TK��b��<��dU��D1�'��i�e�-z� ��ʀ�wn�1�2���̹eؠ��ҏ5�9�2�
^�m��-�<��B�0:]��I���(hy �e/�&vP z�'
�;��>%а�%<�L��#�bx�$��(D��,/���i�!��s���y2���Sd�A�`z��y#V�@�C�tb4)�E!Q�B�+j��a��UV(+��.���� �$�#_*.����)#�Z��a(J�%������a~R���j�@)7�	y��dp�nāxn^�{�!E�4��4 N	���ӥ$��Sh��wޚAE}���m:4M.��O���c��x��e(0�ɃS����'	�Dҕ�<S��k�W�H�t��Oz���߃���H�L��&9 ��ׯ�5��ٔ"Of@�3��T���rΘl�~L�d"O�1�FO�4aI0/�&�8�R�"O����	p?�9�`�V�%B8��c"O��;��۔H"��#��ؾo�LqU"O�UX7�,c�LC��U[�	AP"O�صb����{�N��M�@�"O�̸��е�6�E��w��6"O�A��jL�~���]�5�@U�`"O�8��A��� ���Z;���G"O�cd��&T���jSB�(�,a��"O�\1f��>*B�#��GV���$"O�@��I�W#<����Z~�4ٺ%"O�ؐ�R5�U $@C4G���� "O�Ё����&�Z�0**��"O��aj�&	B i:�i�T��e"OV���"�� �L��`���"O�x������ ��dd��+0"O*��cӧ5n���K�%d樈�"OPp�P �@|*ٔ�*A[V��u"O���BA�Vg���I�$CL=��"O��@BL×S�$�	��I�v2ŋ�"O�Q��P�0Nuya�\M�d��"O,�*�AX8ux�y1��Hp����"O�ʌ�@dd�2�21|9�"O������$��`.K1�� �"O����=���g���Q1�"O��{�
��o��H�`��!^FfQ�7"O�)*���R��"d��OA
T��"O�ep�E6z����$����'Ll�#�B�A��D37�b\�����A=M�*���'tJi@U�κQ�R����YL�b��'�X�;�)��z>R�A���l16Q��' Db!��6�H�j�I*UI�ex�'�*t�b��D. j��CV�@� �'^�	�σQI}Ɂ�ЖHV8|I�'�8�"%��V=�� �@�*+�DR�'��sǤ�'u���Y���#���
�'��P��&�l�¥̯拉i�{��O�O�de��l>Q�@��Y�܈�O� 0� }��S.'= }�ƉX%c�ڵ�d����F�'o��Q:Ɗ;K�;�o4�'�D�I=!������@�	���iW"�$ �B��똮oo`�@.]v$�I`4���A(Z�1����dN``�I���������Y;M�7-̸ ���~b`�><�k�ς�C�T�qwL�'r4㣰i��]��'f�@��~���ᲄ
ʘ�S�$Q}�Z�ߴ0]����ELٷ�u��C��)GC����_�.3�ĹQ��)�p�9lz���"#	~E�B�O�du��LJ�@�Iٗv�`�l��%{���):-�����L�Q?��53uzk��Ȩz1�f�J1�U;C�W06M����Wi�,���?�"���>h�.�3ӧr��ťC�r�8싶�ґ;��I�.�O�q�ŐE���7�N3M���H��_#����'�4Y��L�>� �aFi�[���
�M֨��A�??(J�x��Uӣ ����uB�^�$��X�{Ⱥl�v�O.��7a�(P���Kƕ��}�u�N�x�:c
K!s�r��q��^f����/3��:g�'���'��JP�у`�Z�)D#J�ek@/�+�9 �'Af5ڱ�v>��Qa�vbl�S�ml���D�����1d��֦]�HL����QV�
5� ��?onYQp�6�!�$ܓ�V�Q�@	I	��k���{!�dG���{�c��Q�-���K !�Ԟh|y���]�	�`Tڡ�T!��.(q��P�>ނ�`����8M!���j~x��nްM�&Ի�oOm&!�$)M>��6���_�N�x�ˋ�E�!�đ�i@. ��X���T섁�!�d��"Z����[F�y��lZ!�ڧ/M���l(�]��0Z�!�dE�Y�Lu����r ��0�lC7U�!򤇌
���:ȘUಔS�,�%(p!���ƾ*���.;�`�`!u"Ozk`�C�S��0I�ڶQ5�!4"O½�%͟*��Q:7cG����yB"O�t�G.ҞAQ�X���5C�|���"O�3&�
7�\S���%=H���T"O��/��"dK����V���"O�$ J�h��Sg$��N1��"O��p�f�Ǯ��U�B>D��1��"O^D�$�5�@�'"�5"�� "O���
�"(��`TʊtH"Od����Dg$m�ʘ(G�xzd"OZx����?�Ry붮X�)O���"O$ಲ�ɘ_��I���4H>�6"O�xX��\/>�0���\0�x��"O��@2a�R��HtbE(f��9�"O�,
~��R�A[�Y���"On�JT-8a�J�j�3R~Ń�"O@�r�/��80�\����"O��k�e^�1B4̕�H<�qQ�"Oj91��6�Ժ�K8���b"O�\F#T�V9j���ןC�"O�zB�0I�9�(Ж~�D��"OXD;�'�9������T��K�"OPh N��>w�8�&��8/M
��"O��c�I�S*a�L�9"����"O�y��G���L4�u �.P���"O>�0�C�B�DH)v�����"O�I6�I�E���x��M�d��Y�"O�袮�T�̝ O�DBh�C"Of���㒸q�d�d@ǔ"��XI�"Ob�Kp�J�NH�� g`	Y��p�"O��CW��N�V�9�X!��(QS"O�`�	�1 ������LP^y��"O���󃊡AJ�Hj%f06�+�"O��2C(áB�<1i��(5z�<�"O��#�I��M�f����E@ ��y"���A]���Aϵr��p��ġ�y2�H�	����Ԋ��#��`�y2�]X���@,�����(�y����y����1L>����<�y�� �H�����G%"⨝
�/�y�m�:/#l��5��1�n�k�T!�yBϓ9���Un�.�r�8P.R=�ybŘ!U���J�>�i�v"_#�ybƟ6+X�ّ����d��l;�y������X�D�0^�H6���yB@�3<��9V��ƈ� ����y
� 0�r�ǜ�B��E)r)Dzo��c"O��I5b�4|�E���_�f`=�"O���)�L>9�K�y���u"O�i3��dzX�c��v���`"O��+A�CQ���`2H9O��|�"On,{➑- ���)EB�x�"O��1,ʳtl.�HǏ�6ؼlhP"OV�����8@���C��Q���!"�"O|ar�)N�g��y{%(ˤ.��M�"O\�q&�@�&(�G�V)vf(�"Oh�IE���`px"%�s�7"O��" #׹a������V�b-P�"O\q���ϵs��<a��	w��(8�"O�0��J�T����U
�2���r"O>+0�����U,K�P��ջ�"O�i(��<O_
�K�`*"����7"Op�C@��r��8BUB!E|D��"OBy�b�@�X��V��b<�x0a"O�<r��f�4y�&KA�ڴSQ"O�� -���Zp[�CƻK�4t��"Or0Cj�i����+^.~��"O����C
$�@-C���I��;!"O̍�C����$ ʒec�Rp"On�HB�'b���3�!Q9 ���"OD�	W�ɳLN�+.V�E2"��*O��1��^�`i,jơ�P�'Lva�U4w�ݸEӤGn���'�(\�t@���`��B�{y�p��'��x3�G�[��4���v��Ѳ�'�6 A$(&�4�`"B�f��
�'�J����Z��U�"GX!DN��	�'� �҇�x氵xl��?�ج	�'_�b�'�r�ԅ��@"G�5!�'��@�uÇ�<T��(5����K�'4FXgh^3 E�AԈQ�C��E�
�'�|�R` �B���j�.=�P��'p�� G�N�t%챛0�Ԉ/�xH�'��8��J���> ���qd��R�<�A��q�n���J4V��q'�TM�<�Sc6(�@�3�%N#,�ؐ	C�<Q��B<=,�R
X.H�XC��z�<1t�@�y��P�E��ٰ��Ӄ	s�<I�Ǐj����2e�&e�&|Hb
�p�<�THӹ<��(��&MB�4,x.P��x<j��"l��T~��fGU�w�|�ȓy�F����<.]D̩$�����ȓ�v�UB &M� ԓ�_�����ȓW���T!��03�^�f�ŇȓbY�$5���}'J�q���k��̇�.����@�m3j��3��9ԕ��(z���HWT �3(��0e �ȓB��r�"������`���>���v҅2pm0 ��e�DǒL����_Y��qG� 1Z<�qd�0�^M��c�Fe�t*C��;7���A�hD��� @��%%�t���%S�-w������HTO��|�z!��&@4I�V����4�:`i�@(�lj��D;-����u�$Y*�(�
�(���(7��ȓ�"�0���w�Fi)��4�q��cx)3V��txİن�ݞn}�(��>����	���cSq�Vh��1���H D]���`9��Q&Q�"��ȓl��$
 �ͩI�x�R-�%��M��S�? �!k`f�I���tA��^;p�(v"O���c���F�P @S:� ��%"OiZc%�5[��;�.Z�2�R�Z"O����>��c���)d���9�"O(��Gc�����K0�ט%��њ"OLaeC>��@��] SE6��G"OΉ�&	Y#��9 #�7&Ԭ�Ȕ"O6�aSC؞E��<h�dB�e�h�@T"O������7���q���u�0X"#"OD�"�h�6QdQJ-��(��y�-�569(FhD-N�^� b(�y�-D@�)�e\tF�A;!����y���]�"u�T-6�x���܎�y�C3"и� �-6�T�A��G��y��џ���9-�
̡�	L��y¢�6Ȇ����)SpQ�pG���y�� ;~�8���"'G��q���.�y�i4a��%�g�E�#�����F��y����?��]�������nǵ�y��ޙYl,�g�G�~}���DN[�y�"C�J�� ���s?�E dhK��y�	$w�`d褁 �$�&N
�y"��!zk�U+ƀޗ�bX�j��y�C�]v�h(�NR�\!�Mq��O��y�>p(����Sj���hȆ�y¥�&1�x'B�sR�)��oܗ�y��؆mS���ЀI!z�Z�C��ɵ�y��_Ҕ3%�ǃ�"=I"M�yD׎
7����l�zI rjY�y���!���e� /�4���\��y�̓p�I�D�O��H@tQ�y(:�i�BJ��5�P:T�A)�yb,��WhX׌�<_�.0�6I��y¢�7[cz	�@�^��0�p�.�y2K�%	�-A�KR�T�T���y@]�`I��[ϋ[��a�"�y��Ι`!6���N� ����H��yB�L�UOf���� �T��g�yb�ǌ]9����#P��A���y�O��@�h��`
7��A���C��y"�Ղ	�I �5G�|9�����ybe֟/��u��ۧ7!2I���y��>A��|;�`�;���j��E��yRc�|��Q@'�I�'P��̊��y�Ä(*�h7�R )�y��l�4�yr#T}�H�y΅��V�gA �yB�^�u���)��I�Tp�뒁�&�y"�Ӓvl�ڐ(�TL����N��y�#Z_ 2M�R��3_���+�yB(^�}�t�C���SڔрelC;�y�#�P�%���V�9�����lG��y���vO��j�+�4�F�:���y�"��FYA�cU�C�njЊ��y�a["'g�D�旴R��K#!�*�yR� b���*QǎG��BF��yR�Ö5��Ó��kU��{E�߃�y����?b`�D��ڭB@	�#6�!���'tZ��@�Xb��i��ʾw�!�Y] �i�ŵS�, ��怗r�!�ď�1����3�\-��+��E�!�Ւv���`�ܧA��̣�I�[s!�$�zTlqzC/U���Ͳ󌏯i!�� $2����\(Sz:�p��?r!�$źC�HS��$���{�  �?�!�� ��۵��"2"���
۹+v���"Ob&���g6��H� <+��{ "O ��&��$�<(�'@3 �x��"O�� ��r�H�ɦ�@O��`�"O�-9���y�8�J�i��T96�j�"Of`��	�
 ���ɇ�0А� "Oi�qG������T����"O�myʒ�h*8a�b
�7����"O:E���(�ؼ�"�e�`T�"O�ճ�   ��   6  n  �  
   �+  7  �B  �K  �T  �]  �f  �p  �y  ۂ  ڋ  ��  �  ��  ��  ��  �  ��  �  R�  ��  ��  '�  h�  ��  ��  .�  o � � � � # �* ^5 S< �C %N U L\ �b �h k  Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�� |d��"O
`�(�;���8���-0��1%"Oj4��ND^[��"3/9�0|H�"OB���H��*�ʞRy=a"O�味V�!X��!&F�:J�$���"O,��a
���C�Ą�M�"O,$3%o�-���p���+Ն�:1"O��ݢ1����`���y14]2��i�<�6��{_���c�H�`�fX�$Kn�<��A̼VI�xR[�)�Ć�pඤ�ȓA5��('nߡ4�� �)˩%� ���,��r�؊b#`T�eT09���ȓ!�b��g��}�8�F��-? �ȓ
K|m�ș�VṔ���2�%�ȓ"R�X�j�4JN�1�˘X�i����̹	_�jZ��1!g��zܶ��ȓgil,*�J�
j�Ne��i�J%b���f	�(U��:���G��$Y^م�~r�� S�%T"���k\�jx�ȓ|4�1�îJb��@ӵ�ݩn�V��/[`�"�v4�R�!ʎ<��M�ȓ`:��z�ؚh�J�Z��$HY:	��H��p�m�C1��!��B:��0��EnjZA V;9����J[
2���	��4'J�EA�IVW&��~�(aZ��ӹ�>� o�Y�|�ȓ�f�A�
Ο7�H��M�$�����mޠP����/���ANXo*�ȓTv�����{ ��-7�*h��I��sB�8�8���3����ȓNe*M�悡;������X�o��!�ȓ'lj�#F�m�+R&;�|��2)n�C��0S4���T:
b���:�0!��e֊��)��ͷV��,�ȓ0�&�8#���� ع�L�����;�P�AFd���,w�6d��r�EQ�( �gVlɦ�M,H��,DP���|�I	$G#\���O>�=�JTf*����)GѸ)27n�\x�lExZ Ɍ) ���P
�ԠmT��y�Gq��Qi� 6�LYq\���'�ў�O{�Q9��R�[�d��a^h{���PD,D��:�aO�$���^!
ӞT�t�4|O�c���p̝��� ��_ƁáG4D�<�f��zb�Y�g%�Iy3D�@�Ăj��p�ф�.L|ZH1D��I���Q|���"�;Y6H*��\Jh<@W39Z��bȂ\��5x#/r�<�$D�;]1X�
�_�HjHtKC�\��?�	��|����D痡C8��d�-l1t��O:�)�Q�$Q&�E0Uu�i�0o��1 ��y��[�'ɕo���! ��Y݊0%��E{��d/��
�*�x3\�1`���y�F p���
�G�.U���y"׊ ��P� �S8Cg���m��HO�O�Ly'����zI�-D$Ɣ�"�2D�� t�b�k��,��x�0G/��Q��ħ%�M�i�I����ܘ;�ȓm�i��EͰB� �@C'X,C��مȓ/Ǒ���a�^UA����e�`��� �2%s!��&j���F�$=�����B<Yu-��,1�d�b�ԐE� ��*X��`�'�>� �ia%C� }��\qtL3s �+"O��#����z��q��,���q�O���>1iQ�b?��B�*qz`�#6kK"����B 9D�$ٴ'Y(l��{��#9PH��%V��x�`@Q�~��4e��N�`���yₙ$
�>�V�N���=�y��]�(��=���V&8�Za��yb	A�Q�.��޽(y�]hf
H��y"�P�!��,bF��&_���E;�yb�!R���KP-.�48��Q��y"�k�[E��]��f`	�hO6����T�8,�բ���!�qLڅl~���G��j�U � �2^�@8a�I�y��D/[����֔I���؀cW�y�ȅ8j>��E�0G�ڨ{��Cn�<12�H�V���J!Gf)���)#Q�	u���?1�>��欄2ԍ�X"ك�&пt�lQR�'�24�
7�R����tY�}Rd�8���'Ќl)�d��}Ȍ䀄�z�rX�b�)���΋|4y�R�R5*S\�␠
#��'��"=M��a4�'��P����9g
$���,�$�P���O�H�d�1s��`�1!3}��k�7D�0joR�U.0к��B�M��!�7}G����=���8�R�'/C�)�V�W�]�B�I ��9�Pl��Th��qV�$w� B�ɵ%d��H��RB^� ����4�B�)d%��
�+�"..>�z�@
�h)�B�	��b��cj?%^2�s�[,dn�㞠	��)��ً�|iA"ǫ�F����푞0��I)C��(���%`��P�F��&�Σ<I$ 8OpaZp��2kF1Zb�^#�����'���(y�B�v�U=g�2P�b�^R������Gy��䇫@�L��#��7�d�c��Ә_�!�M_L����L��T�嬖+^�!��k1荘��OjD��5j��t+��0p���O�!�*��s�\Q�G�m����"Ozq�D�&O��u�a�],s�l�T�'����)��w���/��S"CK7=P�9���<+��날� ��=��'�I�Y����D+V�j4�����$EN�'�ў�?I����0_ބ���`;EJn �G�!��hO�S&P��I�B�CX��qѨG�4���I��~2�i���>m�1�T�

�W ��`��"�I)�O��s>l���#�`���e��ZƤGx2�i�ax�bC��e b�E�~�p�qEʏ�(O`pD{�O�j��FG��hpW�a�`���4D�Dh��+T� ���4e��D!1-4�	�<��}�x�@>q��e��k������
��y���j,  ���,	� `&1Zz6�ɜ�a~2Oʪ��Sj��$��y�L���<1��?.
zx��F�+���4g,�ZmE{���'��T($�H���d��,˵0��[�{��ZA������hZ�tcB��agT�K��5o�������'Z�ɳ�@�J���;��-l�D��$����HN�8T'U����
�:�00���$:���AQ�	�� ��&�(,@$���i��4D{�OF����a�}<�BC�>ن�*�'��|�����X��Q��g��Ġ}@d�"C�2i��?ьB�	�E)�01(�N�.���m:�O&\"��d.��1�D��G59��hB�ф?��	T����V �ip��c���,@\y�ď D�@҂C�^�Za��Y"%�*�b��)D�|Zp��4��9b��#p@�����%�IZ��|`��f�j�kf���>�T(� /D�� P��?vRN�E���D`�1c+D�� �b�%^;v��+Q"�%�@"O���E	�F/���Q���]��9�`"O��	�H��w_� �΢v���T"O�X���m�,�'+�&+���"O԰��ޒp)�e�qIP�B����"O���t*��RP�c�f$� "O�ɫ���$(��v��T]�"O�$�/��Q����oV\�Jy"O�|���:�̅�m �m0@���"Oʕ�v̌!5�����2h0�"�>!���	 a��xb�瞕g����o��lE!�$��6vdA�U,�����F����Ġ>�DA�Od ��eW�3 HP��Lh<YVE�1w^v����J82�=����3�y�	�8���{��;��exp����<��d�4S�B<�AF�m[�TC1�޳3&.6�5����
]��l��2���iO�Ic")(�	{��
 �>�A�L��`AC:����W�<a�A'}
s���7r �u��{�<�fW8.L�e-�����C�x�<#kNM*)���q���l�/�yҥC(^``A*L'3�ر����-�y�!(���V@?Xsgc@��y"���L
����T0׆8�6$ȋư=Q�{�+�.)���'��:���#j��y��6F�~U)� �13r�a��y"�RK��Xc7��Y8B��v%2�ybm̅Tj���FfI�Q��E�'�+�y򍐪}lh�b��C׮�I*�yBo��e�R�򌑴mt|��'�0�yȐ/c�VTi�O��
_ʨ2V@��yBL��_� aJtc�z�R4Q��ybg2��1��2kzr��PF��yB��Z�Nz���8c�$;P �y�n�8i\倀�G=�ة����?�y M?�CA���\k����y�ʗ�a~�$� �4-�(���J��y2����J7�R�2�n�9k�3�yR�Ϲ,� $�6��6<�c��:�y򏚹2�(҆�(3���,�1�y�͜�]�m+�ު l)�Q��y��H�$(��q��^)
ĽA�c[��y�Ϯ>� ��4/�zr�g�+�y�#ʊD08�Ɋ!,%���aH?�yR#��Z �"�R�;��ޘ�y"@.Lk�0���J
8�D��KR��yRe߻(��E�NQp�M��yR�ռ3�j�8woA���Y�&&�yl�4o'4�+��K:���k�oP!�ybGS<�Dۧ�̻	���C��� �Py���T�0���+�u���@I�<q����Q��[�E c���QWk�M�<Q�����f�B�NM8o�8䒖�L�<��Ě%�΄�!�=L�2��J�<�,��FO�s#�<yr�M�<��J-O���bƺ6��5Y1B�B�<A$a$> �/�>&=� �_}�<���S��Qp�nN�y��0PF�B}�<���:��Y��>J�� ���A�<��ON�z�yA�Fļz'�8�ʎg�<�@�<�b� fJ� ���3rh�a�<I�f�&y��5��K�6®]�E�E�<�C�;�Љ��ҋZ�6��s��H�<�C��"1�ʤ��Dw��UY���F�<� j!�!�ڧDײ-4!.R��"O��A�F4Mw!I#���B���Q"O2�r�'_�f���T�u	���w"O.*!-E�]���z�N� F"�I�"O��c�Qr=IC���τl"��'z�'�R�'���'��'���'*(|`��C%g?p�B 	����p�'�'�2�'��'��'�2�'{P���(1Rr�x�KX.'�m��'�"�'���'��'N��'/B�'�SQ
�>`�h��F�D�N����'�'�R�'�r�'2��'��'9��K��Y&J; Mç(M��'�"�'��'iR�'=��'m"�'���9��R��z��^���W�'e�',�'T�'��'���'z��ȶaͪO��5`\�P/�Fv�'���'���'2�'��'�2ԎB|p��Y)  Xibg�I!��'���'y��'���'��'i�k�/"�t��ܤE�Ĭ�d+P�5tr�'�B�'���'���'���'� ^>8��m�Ӣ /�̕b4��%m��'0��'V��'���'���'gb/��<�p ��%@�f���hK["�'d"�'��'���'���'u�χ/��נC!G�����)>v��'��'��'���'�B�'|Bk�=u�z�yH� ���G%��w��'�R�'Q�'���'��7��Ol�DlV���ϚU�6��H\�q�J��'?BP�b>���ve	,^�i���]�������Og���Omz��|ΓS��B�*�{P��(������~��Mm����{�-��q�'����Z�N�����.�A�P�ǉ>��8����O���h��%	�@ʄk{ȓ����a�lPƦ����/�Iq�����w�:]��p��u"���(o(���0�s�\UlZ�<��O1�bi��m��I8����5K�8d?�<#�C�q� 扆ZJmV�G�3�> D{�O�Z� Z'��Kx��㉟V86����D,���ঙ£�'�I�"Ǫ�6j�ntRdІM_�]�?Q@Y���4cݛ�0O,�6���2��oRR��eA�2�2��'��$�$�P"�!��cLl$��۟�����o��'�W�%A4mWxy^� �)��<�F�49�����M�_�Vк`�<���i�A��On�mZM��|�V,š�6@[�.J#�A+��D�<Yƿi�b7-�O�أ�Es�$�U#KM�A,Jx���',p����]7�:a	�d� ~szx&�l���$�'C��' ��'��U�$dK�+K2m�k��Pf>Șd[�0H�4x�ҽ*��?I����?ᕇB_��P�"T#-X���A�/V����M�ǲi�ɧ�OI�Ɔ=<��x8�7	i�H�F.�Q�`�j�O�xQp,�.cۖ�];�䓱�$ĔSt��b�G��i� )�ff�d�O��d�O��4� �^ʛVƂ$1"��R &�٨h�!R���z���?���t� ��[�O�DmZ��M��0Gp�f�� :�x�B$@x�b�����M��O�
��\A����d�w=��AP���b�T���`W*ArH�'2�'r�''�'������p/����S�\jr��A��O��O�nZ�Ur�Sß�xݴ��p<1�[L�H���ٕ9j�k��x��%�M+�����A+���������i�l����*)���13LD�֠D�:��'�P�'��O4��E���0O>�K���^��<xu�ɏ�MS�U��?���?�+��CЂ�zJ��է��1�ԟ�xc�O0=o�&�MsN>�Od� aBW85m�ts�c�;n��i�BF�&��J�̡Mr�i>�*�)��۴�|R�\�Z��" � �E���PS�HB��'���'����Y���ݴF(p4JB����Xزc[n��=�L� �?I��Y����N}�#xӦ
�"P��6a�!��^��c��%��-MN�n�r~b��p��P��V��K:ZKz�����1/g\E���ֈWR�ħ<a���?����?����?�,�l�b@_�%ʀ��ͷEZ�ɷ&^ڦ)j��pyb�'��Om��h��n�9��
���#&�� BNZvum��M�L>�|BT��&�M{�'�мx�f�8lJs���a�"�'t�p	���5�B���|�^��S�����V0r�.����A[�(���ޟ������	TyҊv��١�@�O����O*�2�Ft��Ӫ�,Bjp�	2�����D�ئ%hݴ��Iq�)���W+�X�Iܭ �J��'�V�9�W�Mx��;���DJ֨q~������w�w$de3ЀK����v�6D�H��HΊ}��2@��k����G$�ǟ�Yݴi\�\����?�g�il�O�.��y�ڤ� �\Z������̒s���ʦ�8�4�?	C(^1�M;�O����o]�x�΁%- �:��}0p�!��l�3M�*���O�ʓ�?)���?A��?�BJ�����5C�4	�A��D�0��,O�LlZ��T)�I�P�	D�� ��K_5N*M������a O֘��d����4��Şp�� ���ߌ�´E��	�,c� �@�L��'"��t��"��ΔC�	yy��I�>��P��⋁"䊄�\���'r�'��O��	��M;����?��v��e�g��>i֭[��I��?!мi5�OΉ�'=�6i֦%�I��0!�ў+��)¡��
�B�
���i�'�*���%N@�}�V�Mf�? ͫ����%A��,��+ׯһD툘X !G>	h3Iؾl�Bm���>�ФB��8���kV�٭h��� ��/ST.��Q/:`YBŭ�>�R���Dq@��ca�@��2O�bܓj�h��~�
�)�29�rm�C��Oxa@7+ҟ$��3�ћ!(��[b�zM邏<-�"͹���c\���35��a�Qj�,� ���6>@A��N�	�.1��	=cAV�CB9)���;�i����V�W/���K�̽�&B�^F��K�&�M����?� ��u�-O����O�����c���,$�%NO 5�@�S�J7�	�"�5�D�OB���O�зOr�x��"�@�Xt$�2�"���	���',2�'R�|Zc�6���\=e|!*�'_�ZĴ���O ypi1�$�O4���O˓l1`F�۵\��Uy!��T��-���܀��D�OX��O��OZ�$�O�|@�B֑;�:�ss	ܿr�ީ� .�sl�O��$�O����<��I;������@��)0 @[:��e.��M���?A���䓇?I�^.!K�'R���O��A1G��(1T= �O��O6�ġ<qD�0\������o� _>y���Đh[P�`����M�����?���P� �{��N��(4Y5�ْ���2�l�,�Mc��?Q*O~���G�|r���?��81l5A� O-T�P�ҥ�
	c�X1@�x��'���@��|��ZlÂ��6l�#e
�Pqr�ib�	:H�N(��ş���̟P�SJyZc����Nݰ}�4,8���o�
��ܴ�?�$������S�''�©"���3�̤�S�C�@N8nZ5U��Iޟh��ȟD�Sqy��'&Mՠ@��5� FǭbdJQ�&�ҕ:I�6m�+j�"|���S�z��K �ApiM�8�W�ig��'�Q�@=�꓅���O<�I����$"��CC�(�Ɗ���b��	G��A��ܟ��IƟ|�W�Y�0}�KѮIyh�hvDH��Mc��q���,O���O��7���F����<7�||	��<�Ή2�R�|��*'���h�Iɟ��''�3��-��XPC�s8z2)B�D��	�����ğ'����ğd;��ě-W�ـJ@2#]���sy�%����џ��Yy��R�\���:��BƔ�INj�[$��KC�V�'E"�'��'D2�'�*�b��'G�M
� T�l��h�e��?�1!q��>���?9���đ�+Bj!%>%u,ò�u�T��u�Ũ�M[����OD��|2����	)4k�I��(u)W�'�7��OB��<�2�H�`��O�R��5�T7��@��6򎬈H������O��0�9O�N�,E\��b"WAQy�UF¯Л�X��˥-�M�]?!�	�?A*�OLQ��,ʤ!-2X����R�E�6�i�"�'S"�'���'��|n�?_踚�oҙVf� ��H�r��6-'B@n�П��	��t�S����|�B��/� �ae+�b�\� ���1����'���'e�R����y��'H 94Kچ�����'�9^bA��q�*���O���ʙ��=&���ş�	%i��]@��$"�@�Ք&|@���4�?)����@_�TV>���M�wl��ir��R�E8����Dܦ����$\�'h�꧹�'��$Д�2mv	2)�L����6.��<����D�O:mb!��L�0����*,(�H5�S>�lʓ�?����'���O$X�t�(X� rI\#p�8�i`���y��'R��۟0��ar����X����8&��������u�	П��?	���^�՛��G@���R朅j�����NU)���?�,Ox�����.ʧ�?�!�FX����Q���d��Aƙbܛ����O|�bgX�'�!�̈́F^��f�P/q�TzU�{Ӓ��<���|.��/�����OJ���5Vk]�i�ذ���0D��f�xr�'��I%�"<��"�*bÅ�Wn1��!U�^����'/��M1�r�'b�'���Y���v.%{�MڡRPҘ�s����7��O���PGxJ|Ҁo[��Hh��&�V���u`O���p�D^ǟN�a���?��'��?ik�����x���(!��
�"���$��r��b>��Ɋ��	G��"fP=(��9W��9��4�?����?�f��=SӉ��4�'��"��Ҽ��4Lf��x���.,P6��O\���<�R?��?��XiL��fX3P(R�B��	��h���i�B	X�FO��O:�D�<��f�>k�r�k
�o
8�94BҲ%��F]����jyr�'�B�'��('VDȱ��;6f�C	8S)썺d����ē�?��?y/O��d�?qY!�U��0�1O��a_Dmh�f~���ĳ<����?�����$��%�
�ϧ�$��#��l���N�v4�Mu]�d��矸�Ihy��'�����e���ˊ�󺅓*U����'TR�'���͟���w���'8(pydß2k��+�*ٕW��\ӎt��⟰��]y"�*�ēw���sF�I�f�RiG�5zƵn̟���lyb��/�f�p�D��kl��6)Ӡ� �P|�R-D��6R��	ԟ,��ß�$?�i���q@�>/��P�ܝ0���z��HN��6�iz�맅?!�'���3W�Y�EQ6kY���4 ܄'*47��O��d�O\�$�f�s���M�K�2t�+� T_�rݳ�f�}�ec��M����?����b�^��'~�*������c�X�Q�D�n�0y�P1O��O��?u�I�� 9�4aϔ
���@�B������i���'�ώ�>X�꓊�D�O��ɣ\� *C#
"��P�Re�Q��6��Ol���)�S�$�')rݟ6(����p��%��?$:`�%�i�b��)������O�˓�?�1��i g)�rpВr�\�f� �4�?a7O��<q���?A��?9���򤍦 �v�3��NHz|j�G^�y/�Л`n�]}RS���	tyB�'�R�'bzX�#/E;L��sEL$O����S�_��y��'R�'�"�'�k��t�O*�РI#ay΄�"oԬ:+ܜqܴ���O@��?a���?A�/��<!&A��N�:�B9�J�CG�?1����'"�'�2V���DD����i�Op#0��o����"�#*�U��M���U��Yy��'cB�'kT�S�'��Ovܩ�%N ?�1��N�Z�.�� �i@�''�I,xi��Ҫ�^���O���H�X*�D �`��"�A��Y�b��'��'���y��|"۟�xy4�\ X{�D{��ҁu&���i��'J�CP�dӪ���Or��������O�̀F�E8�242�n��G��I8"OHp}��'`(x3��'Eɧ���~R�M[��8u��З�ց^���nڟ~�t=�4�?����?������?��q}0�G�9��83�T�ERjy�źi�R�9&�'e�X��\�㟜�P�A%~ܩ7,��w�T"�����M[���?���4dR)��i���'���'RZw���Ȓ��\d�!��v�����4�?�(O���#<O��l����U&��3� �#�۹?f��t�Ɉ�M��
$�\��Q���'u�P���i���wlĮ>\�*u�@�hv�UB2�>�Q"��<���?����?�����i˨aczQa���;��3��]�^��Ħ�Ѧ�Iȟ����T9���˓�?yV�23�D�P�cܑx���4.��+B 9�����O4�d�O���O���WЦ��BW�2Z�A� "9c�X��'�
�k�O2�d�O���Oh��?�r _�|�U���Eì�� ɮWR�AeA�j
���'��'�B]��Z��V2����O�b��k�L�7N�D�p��������Sy��'n��'
��k�'l��Ol�Ʀ�q��w�ټ'w��kF�i���'���'h�i���m�����O���򟌱q�D6t=��U'�@��Ea���㦭��\y��'��x�O{��f�ܴ9�����.Ģ^LX��\�8Ǵho�uyR�ǁw<�6�v�$�'��D�(?� B��2���J]k���
�M�	�l�1BD��D%�b?-z�ބi�����ްQTT��$�qӬ����=�I՟D���?q�O<���5��H��=nΠ�R�N
�B%��j��i��p��'Lɧ���d;�&	a�g�I0!ہN)�hn�쟈��柘C���ē�?9��~����f�9�Ń�]�ճ��]��M�J>ـl!߉OO�'Z��J�0��ǄG;XUp���J�ʛ6�'&����*��O��+�����A�8I�F�薊_���Y�P FA��Ĕ'8B�'��O�0 �����>��
�d��l2��`Q�j��Oj�$�O�Oh��OB�:��	_�eJ�b�	}��QQ���$�<1��?�����ǤH�̨ͧ�� ��0(����¤�W���'���'��'���'��-+��'Y 89�㈑t�>(6JL0�4{"e�>����?�����̈́M͖D&>�8��N�iuDT)��
7vZ�YP�Λ�Mc�����?i��Z��h�����	�dd���,��=ʹ%���X _�6��O���<��%��y��OZ��Od�x�@Û2T�ӷm�h��IU.�D�O���� =C��>e�|����9��hxR�A�c@r�m�Uy�̂-��7�\�4�'� <?yq!�~�i�L�+�ґ8`��ܦA�	������u��&�b?!�a��X�����̛�t�B�Q��l�8�/��o���T�I���ӣ�ē�?�vM����=q�(n����!�d���a�.���|���y>A2�yq�����^�`3
��C����Y�����I
n-���N<��Ӫl�[?�T�h���2��*]�@q��צ�'��J��l��'�?a���?q�'>B��Ar�J�q�v��� KO�&�'dl�4��O
�d!��ƈ8)�+�`�(����P�j\+7V���&�ԟ��'b��'KRZ�d�Q�0j?����Ă9a����A���ฎ}r�')�'6b�'j>��/��cY�lJw7�`�4��'P��Q�����L��Gy��X2J{���IxP���(H\XE���-�듖?�����?��4��Xϓ<��{�@�(`K���$�^�5L�v^��I�$�Ivy�'X�_v��0X1��5T ����OCN�	���u�	v�I��p�I�C�����h�dQ%syh�÷��[DؠI3'��-��F�'�b[����M���'�?��'{y�\��%�M]�a�bX�=Wv=�חx��'z�a҅s8��|����ذ������ϐfA����i剶!-�P�42P��������Dޠ7�8	["�Z������Í�<*��Ry��'a�O�O=����0V؂�C�v���4�2D@$�i���'r"�O`�O�i�-UX\�3��I�lh�s��Ν0X���'W2X�軋�I�O��f	ٽ
Z����B��9P!�DҦY�	��I�\{:Ԕ'�������@����:��%0-�)n[,���I���'�?���?@B�~�������'Tp�p
��x:���'	&Y
R�$�4�����O$�'Y�h�� 
Fc:آ`�B�J�6�a�O���d�O����O����O�,� �8��+F��(�Ǫ�>Hh�q��D���D�O*�$�O�O(���p9�b��u񆨉`"���Z�bӦ1hC��P���4�	|y�B8bY.��+�޵�#&N��.����� ��?���䓰?���f����'U�'�X%&�]
��,0bЍ�O���O&�D�<��N�?"�O!�9�R�Ă���.C(k��h8��}�H��:���OJ��H�O\ #6#[mǎ�EOD�7M�{��i���'��ɒQ���I|b����6C�-%�l�s�o#6;�1 �։'mr�'2~ 1��T?��(-:�i���
{�l�z5�s��
]��S�i�<��?���F6�	Q�\D���.:���07��O��� (�b?)!G�A�I�.�� Fl�|��vӠс�IŦ��� �	�?)��}R�AMp�Y( �y<���ޟRt�6�ǎ�������-Ϛ��C�'P�"	;W� iF�l�W�iY�'�b�GJ	�O����O2�I3D��0���?s�y����v�*b�$j��=�՟������j3�č4��큦d-_SPp��9�M����6pcқxb�'~|Zc
@��^- @�� ��]+P���O�9a��O����Of�"�XjTP:I& awi�
|t�JB�F�:6�'���'e�'���'�8չZ�h%��m]&\�HX�$��͘'���'G�'�roҡM� e��0�$�4N����&���7��O���O�O��$�<�Q�_ͦ�W���2��]x$MW=�p����>����?�����κ"�t�&>�B W9����*%C�D�ᢉ�
�M+��?�����>��Oɀ�$���B|⹱@I�9�n��4�?����?���!i0=;(���$�ON��B�!( hjĈğ0C�@su$�&�`�Iby򯌜�O�g-�4IvL`��D�v�I� ���\�b��M;�Z?)�	�?���OF%2wiѤ��|6�F�yP���1�i���'fV�����	�1w�Hx��"����3��:Q���JQ��\6��O��$�O��	IK��蟼���X�"��#�Dƿc���zw�$�M��
JI������M@���I�\
�
b*$p��o�ٟ$�����C�����?����~�m��a�GD�>N�V5�GH>��'h\�
�y��'X2�'E�q�u���	(����$b�<�CW$ӈ���==��%�����%���C� ����<Ť��@�M�bJ��/���<���?1,O���U���|w���Z�:p��q���"co�O����O����O��O������Y�B�_?ĥ��I�2�����zӀ����D�I����Oy�a��+7~8�"��A.1v��bU1r���?������?��{�F6Z\h\J�莤j!*u�kғ��D�O����O�ʓIQ���c���֍P��{��R:����ơ+�\7-�O�O���O�	v��K��V杴g�DԪ'�AF��V�'��\��J�/��ħ�?��'CK�6 ��qۂ:5�`@Ӡ#�:�ē�?���>��Ex���uG�0=��k�.+a��؆�i��'(� e�'��'b��O����5&�ë��h�Eʐm�m�N�$�Ms����"���*I�d�/6����˕H�LEH�iu���)}�*��OV�$��Ψ'��S" �({��74-�`�%$�t�޴f��,��Ϙ'�b�]�!q~�ʶ�f�^�j��P 2Fx7m�O���O�����Od�D�|j��~��Q�bȻШ߲%s@m�A���,A6#<ac����'���'rDE e@�F�$���'�<�t�[ܴ�?���A<�'��'�ɧ5�ߴB�e�dGrq��,�;���=X1O&�D�O:���<��OQ2:�e�͒6��,
��`ǶY���x2�'�|"�'��W5��U�
�-��1� L(~��y��'��'�B�'��ҟ�u��f�_j�����3�PZ��i���'Rr�|��'S�	%+�6P/|�����؎�4EQ��<)p������I��L�'�&I�q.�~"�z�X�m ��x�w�M!vж�A�i^��'��O2�d>��:KT�rE @���0(ŚGy"�oş<���	�(�2Y�I�����ʟ��C8�9�5
jȣ�#�%�l��K<�����$��g����iT�ա���_���&"D�F�\E8u�3�L����/@>zD�LW�Yv�@q@̙s@�� A�R�,����<M*le�Q/e�(�QLҰ��	P#̫d��ŐG�'�y� ���x2W�Z��B��>Ѩ�	74z�Q���C�x���nѶw�]C�c���ŝ"�.+0��0>qq�MOF�(,�cl�O桃`��Q�"�{5���W��h+�(\*�֡���̦a��X؅h��<�����?_��ܺ����C���k"*�6��AS�K~�L����T/0� S���<GV�H!�[���^J���C�O��d�O��$����?��M�4vz��bIC7;*n\�b���ԝ*TZ,&�6L����נ��'�b��G�?�2\��]�� +e����`M
_��������*���9�4$��'�?��X�`�1O�3BU��bP��oآF�>�R�O���'���IKyr�XO.�5�¬#J�ȳ1jM?�y"��]Z��� 0z�Q���['^"=�O�	fﲌ�ڴb���b%�ĕj�4ڕ�B	L��T���?����?�'�?�����cO�z��QUN�<Y���b�=d}$����բi�sc"lO��a`F�/��@� ��q�&�6�nu��C��/mD����=�ťM�����pp���m��kX샥��:Y2F{�I�K��A���D�$8�!�^��C�I�f�:1�V�ӻH�*4�q �)���ɼ����<�H�x,�F^�t�O���[ 
�4�t]S�L��.4S�F&�"�'"
�����T>���C�Hd�!�Q��;w��Myqg+�4n<E�$&�OѨ@�͔t��e���ś�(OP��b�'Ȫ"}*�eƟ�V�R��ͷb�E��T�<�p�;*� ��i�?�P�X@mi�TJ<y�.�6m�H1��`�!.���e���<�R�_8Y���'�2T>q�fQԟ���ßT�Q�B
o����ņ�$G��0�4�N�>�8�5K�4��S����'g�ɚ�J�X� }p.�(R\D�t�մp�<��<���O*�ʑ`7��Е.Տ.�B����(	j������ٴ�?)���'�������3�������%G��h�'��'UH0�H�U�|���-��8��d����Kk�'�哾%�l�y҉44>Y���.��u�I͟|���4#��	�\��ӟP���
�$ˈ3����62��;r�3���f����cz!�%��Hr|��&^�M̾�sE�ݮ �w�ٕh��x���~F{�M����A`-h`�q7
�=�2�X7B�'���d�O�ʓd�d`G'	s�lj�/S> ��?��f�U<��򥃪!�
��i���|ʟ���2���M�����H�����1��T�?q��?��}ڞ���?��O�Bh���?�d������ɾq\��P8����<��ͬ�����C�69�0� F8���(�O�yn�Z�t:Q�̻I�~�S7j��t��B䉿����_.:	$���M	Z4B�?Q���0�P�<��10�"�y@<�I�Bǲ	�O&��|z���m�4�!S���6[@�d�ǻ%9������?i�Hżt"QE֐\�t�`@Ʌ1<*�(`H�l̳I�J�[��L:[�:��T�ɾz��)��A�Y؀h:sA�c�5i>��:Bd� QiԲ�WN$�<�4A����IL����e҇F�\P�B(Y���ϓ�?y�xi�JT�͍wjY���{%�i��ɂ��#���#��#=L�`���}l@ϓx㰥�Ӽi�b�'
哑D4����韘�I6�*�c��WE��x�q+[*5�"UXA/����<��O��9�Q�)ٴ4��K+�@�K`��	d��#<E���>���S㬟�av�8`P�D�qe"��-�<�?1u�|���'l&��HY%G���g�^�xp�e��'뒹P���0M=4}���ܑ�v!��$Q���I��F�Pp�o� ����t����O����Gu���O����O��;�?�;"���K@�|ۈ�� s��m�u���A�n��$�Tb>R��eX7i���	�n�Z��d�.3�1P�cI(�� ����d��O�/ lO<bw*�'x��y*t�241(T�"O��X���$<��v���2�`����s���((Y�i_�9A�U�X �,Θ+h\�RA�ӟD������ɚN~~��֟�'�<�Iџ��`ߢ=��8��j�@�Yk��;�O�2'[���	�$��ᤤ��S�=S�%=�O@%h��'0�6�ooB�:�(�F��)��D4�!�$�y�D(ԋ�35?`8�6��r!�dR*Hlc��Ԃ<R��*���dI�b<Z��V�i�2�'��S2]5Fm��'E>H�H�ѧ��4������ԟ������y��R�D�<�O5"t������E�Ԉ�8��d �5Q�?�X�8!����P�au�\�3�=0��	��H�����	N�A�� C5l���*"OF����F�9h��	~������'��O�1��L�7D���pF�J�4$�`4O���#��ަ��Iȟ�OI~�Ѣ�'B�'�
Ј�B�4$)��(��g�ӡNȖ�b�T>#<y��A��ABezY���݊7�$`:����OF�05��#x�@)A`e�8C~�!`lQ�6���R�)�矰�r\3h�q��N�+l,�3�5D����Dx�;p�N��Q�5Ñ��'iP��j.O�T�Pq�3
À`�f�J��?!�&��8 ��?i��?�#���4�N����o�~ �`M�s��lk��O>�J��'�b� a�Ą?�W�c ��p�'`�L��S�? a�R�O�`��-�.N�D	0p�OlE�'yv��� 2㜭9�n�-���S"+V�w~!�dضѰq�PǸu�� ��*�Yix�Dz��i	IH�im'&ˈ�)q��@t��8BH�9�t�IП��I˟���-��,�I�|��E�\��a���x�c̼z�9ّ���9����)���Uh��D�yHJ�pF!I������r�'�&��� E�L# $�va9�'��@xC��JF� @��Ů%����'��+V�����C' �k@����'�b�� �&�M����?�(��0�h��9�����)�f`c���f�0���O*�dħA�x�$#�|:��)u"��"G�=D��XZ��~�'�fQ��iU�H���ט0^�e�1]�Q� ����ON�}�)I�,/�\2��F:<W�9CTv�<q��##2�%�6D�����n��1O<��`˳$�(Ei'�\�f����5���<!B�Y�wS�f�'�rV>E��������՟x�h\#���j[:C���jw �#r����I�S���D�$�&m
��E�U"���kC�P���>�S��?ɔ�D�|薕"�Ƌ�q��QQ�ʎL�@���0lɧ����@��lz� 0$"c�
��y�n+��M!�O�)��ȳ���O\�Gzʟ^�"ǉ� ;� ���{#��O��Dد~D����OJ���O��������ӼS'�?,h4Y���7(�b�-�O?��%�{x�d�#�K�x$�QKX�|�6�/��@s�5�Ol����	.	e��U$P�:� �C�O~Y(C�'%P���w!��Ņ4;�����!v�!�D"zr� J�+�;��+6a���j�Ez���@�!��%l��6;*}[�M��dx��2#�Ċ7����������\;���՟����|��g�/���X�aڛA��5[��� $Z�D�rφiz�ixW� Ub���$ &!zQ@V'Q5M��� �Q6ubd��R៛&Ǝ�9"E 3��Z�|m���Oh���#Z�����ɕ!g6�"ѣ4���O�x�G/0$��]�&/�7$���"O��Iw�f5�p`V��w�	a`2Od��'x�	�����4�?����F�`�P0�D��V���/Ne
�P5��O��d�O��)e��O�b�ʧwt:�	�"�(,(�k�fI7.��pEyR����ljvL�c��xY��*v�@����5M��0ڧ@�H��a)Ѥr'H+D �M�(��]V`�bmɈF����(�fń񉑁ē9� x��Z7,�J�ʆL��B��j�ƹ�"�i�r�'"�NTM��͟L���gb�ȳ1N��r�2�� `�6��BԠ��l�<��O�蔍G�l����f�:JR�"��y��"<E��� R,2�O�
%���a��m%��
PER!�?ɍy���'�9je  	+ԍ��`�!dV��'䔰�& �32��H�� 6�hd
����r����ׇ3z������(��sR �S�
��O  C�	�r���Of��O愭;�?�;H�����I�? i�r*�;y�Q�#�m��I�0����a��AC)���-��ɞ9/l��d3}t���ע$-q<����6`u��߾���'�ޠsQ	� &�4A�"�X.���	�'�HX��/۵aXxxsb��V6LAIbg;�S�O�ٱ�tӼ��`D�vΖ����������O ��O�D�.,,��D�O0��/$�\���OJ�,��#�p!�N������'V�l3+O6@B��91���a��5���p�'#�����?��B�g���#�ޥW�H�s�<A�ƥGViy$�ɟt`��
Ty�<��F��M��U�������i`W�<!s��<��n�䟐��W�D��9�&Ac`I=%�<�G�%醟�?Y��?�ǉ2�?�y*�|i�ᜮ"8�X��V�EO^�k��.���J&�<z6��^6�h�HE��(OZ����'72"}�g�BF���,�t��K�{�<3Ě�EI2љ��aO��:�c�t���M<�At��#�8�` +ŌY�<�t�0���'��Y>���ޟ�����MC�}E�PD&5�RM��Q��t�	I�S���$�)�tr�$ûv���GiJ�tsb�{��+�S��?QqD�]���Y����7I�@2B�G@�<��B[ɧ��
� �$� l�wg��{����}�$"OB���gآ�BfU/I�X�I��ɴ�HO�/���I�`.g�,0��e͋W��I֟PX�"E�3̸����	��4�^w%�wW>��V�R�t1u�`-�3��y��'��
�tV����oI">���.pt1��^$�a����+14���*L���Ӽɂ�	\pX��@w؞�Ƞm��n�A�Ԋ�$j#����%D�l�v�U���0Y��J'sZ���)9�HO>��w(G�M���=P���.)^>*A)WL��?)��?a��l R�����?�Oy�����?A$C�7X�9!�9PT�[�GY8�\(b�<�D�*B����V��<W��s���W8�L3SL�O��$Չ;81��i�!�`|���k!��D�*�`(�΂�4�X$s�)T��!򤓃��(�g��e۠i�c��U ��Q}�l�4�jD�i�2�'/�S7s8m�	bF�)7�Æ�4�a'䟰��Ɵ,`��N�D�<�O��i`$W	6"�L:}��P���c��?�!@�.^f��YG��,,l��1
&��`��I��H��h�D�T?J�d{r��.t�,�3�"O��#�G
G���9�eg�+���0>!&�x�o1(�*4+ ��8+|�����<�yR,C�6��O����|�
��?���?#n��L�$����]z������T!8���������ቂJ#�)ٵ�
��Ș�ʐ�\((��d�K�����B�J����S� '��%��ȍ=-:Q�T�'�ҒO?�$ԧ-�y"`��{�<�{�Dӹ}�!�ӂ_j !�~� ����n��@���?����ѷ$�b���B��*����@ܟ���U�u��������,�	;�uw��y�m��d�@ݢ5
Z�X��ԙd��4|���d5c�xՋnG�m�x����hOP��B�'o�
�`c/ě���s���ɟ0�%I� ֜$�@�'$�퉝X��I�C�ۋ L��k �qP�	��\�d�O&��.��A����x���blK��¹[��F�y���y��e��J)RU*�����"=�Oa�	�M����4u����-ϡF�����E_�!0p�(���?q��?y�kJ��?a���Da�������i��pf4�Ƭ���ݡ+��X	�Q�Js�A��Mk��C����Jp�-�N8��,�H8� 3��O�0o~�
}��h��H��2�M�B�2x�ߴ�?)O���>�)�Ǭ�T�&�P�A҆W*̉�E�@�<�������aEDV�u �q1C��<qvU�P�'� ��$�j�N���OJ�'p+��	��`��y��X'RP8��NT�?Y���?���8�?Y�y*�&qc�_,,mܼ۲��5z��i��I�W����B1x�(Y��f�LŶH�@a�'�2�֑>�H�Y�� ð/�l�4k�.D� z�I��>d̰$bǺs�p��b"�O(`$���w��B�С� ɵhBX2���r�C������Ot�'8t�����?���f�Jsw$W���wU�g7�&Θ�@+�U�(�M���
���)&��O,�`�F+mh�)���&%��E��wj���;<���3������'<�՚'�=$
)sȴ8�b��>H<�ٚ7�'8���������<A��Ҿ;�2T��OH5:T�1��^�<���ݷH�I��E߮4�ظ�^u�'|�"=�O���;�!�$t041vjC4J�
�'X��2j��� �'���'bJc�-�I�R���naN���,���(P�fᡟhr�D0�Oz�Z�j�f�)��U�o�,|���O6�Q`�'n:Ȧ�A��l��HS�a���	�'9����2�a{�㓖SrLi���/��P1孙�yg8��u���� *N�)ڄ��X�X"=E�d�ip�7�KX�l�P�΋F<�q�iߜ'�����O����O��"���O���f>�`o�O��Č�J��	�!�	 �[U�o�r�'����(O��Uo�:�D$�3]a�P	K�'b�Qc��,)���a���"�m����u"��y�S�h��ЪT��;0I��`����y��5�B�����,���y��;�	�����޴�?)���� K�q ǲ[;����oP�j%p5[ad�Of���O&yӕ��O�c��'Ar�u�Lы6x@T�##�3�
Ey�O]��n�
�.��M���sf/���x+D�I�@Df���Z�O(
����Z�\�´q�Qb�e�
��� @W�5o@��ҍ@8g�D&�'�<O�:�Q�x��K"=H��g?O���'͗��m��۟ �O�j�V�')r�'��y�MϼR�,!�cK
-�����
�L;�,<�T>��|�	�JP`�N�rn"�M�?'�n�`%��h@J>E���*�2E��bV-HN�*��G��]��S��?����?I����������� �,
3t0<���'���y��'��}�� G�b͟!l��ˡ9�OjFzʟ�{S�V�8��DP�v��q�d�O��$H?b^~U3���O����O��dĺ����?I��R�s0\E�C�n��'iSN?���Fx�̒�(|~i
cN�7Nb�SrO��\�0�?�O��*3	Z't����%�5l��Y�O4�+��'���$�Hd�pz&S��=[��
T!��>x�D!�TĹkg�}�`�Y�<Dz����*q��oZ$-�^ՋvIǯs��薅��d���4�	ϟ0�D�䟌�I�|jd^�z�>���2.i�)S;V�h�҈��Ff����^�q��Ȁ��q���3I��=�pY�C*J�!�H����*im	��� �h<�Ɋ��OpXI��'��̓�\�L��n½B�^%1���C�ў�F�D[;w��(�1�`h�Qڧ�yRF)(^���,R0����ȑ�yr�>�.O^H0�Z���I����O�ZM����
��)+r@�8^�4�6��b�'gr`��]��T>����g���"mC:A��MQd�9ʓf�B�E�t�!����7BV 6E�`�c�0�(O�3�'p�"}J"hN9t�"����'
T��f�k�<I��S�#�r8��N�/1�d�寝d��rN<�6�XVFб��
V)�|�û>��6&Hn%l�韘�	b�������'��Cņ��9���Ix�,5�v�/�Щ��'(1O�3�i�\MR�.P7��9s���m��@��-�?�O?�Őg3�Y9��S�)8BPY6c�O�A%�"~�	4ptʔ�Ƿe�9iU���1��C�	�6��u��jJ���p:A@N�i��#<��)��"
C�L�٣���)x�!Pr ۈ�?��T�@���W�?���?��)y��O�n�F��i��Ξ1�Ry� �ۡ^.��BW�И�����yR��3��b"�ز7i�M��T��~"̚�*�89��/B5��<af�J<.)irC�I��Tу����?������?Aƺi�6ݟ���X�'5�5�H]5��H�J�%�.9��'8�lc�1��}�7'ٸ0	wL1ғ
u�I^y�H!j9�֝b=�����;2{�́FC�z����	џt��؟��+ޟ8�I�|���Nß����D�TaIs�V�Z���Dݱ8:�����C��I�}�F%0�F-�\W��sH����\ gG�@�� acg�2-�6@p�
`N��G"O���P�zThx��E���3"O�"�����`��eM�m[L��:O���>���\,-��f�'+RW>�J�D�e���1��b+:�7� "�����l�	�XL���	Y�S��.H�K���,,
�C�mF�p�.a��

 ��?�Ks)GE�h\h��5&�B�PQn%ʓ�V��I��H��|�j��NμQ�C��z���"Of�q�"C*H8�B͠<� �yR�'��O����fz�\�w�X,��3�5Od0ٖ�զ=��џ�OA$Y���'r�'E��i5Â=L��SF�TҎ�R�ǆ`Wr�T>#<����n<��p�_&�dIR3f[�Y�6Pۊ���O����%|̋&�š#n̸uBٰ/��|�)��h�D�8���Sb\!<�P��!D�8)CCB�R���� Ed:����?`����O�!҆i0;�t�H4�}L��R��?i6(Ξ[�&D����?����?Y$����4�T���h����P"�3�l���O>A�w�'d�`���j���V�L&)��'�FŹ�)"Hy��&^;'ќ$⒤7z���4��)�	O���P��_�V�V�	wM	�>����#)D���f�D�;�
qcB뚭�jq+ F���HO>�+q��M[��Z���a���:
h�����?a���?!��N�Ll���?��OY�(����wѢI��蒖P�:�z�	1;��D҆ �T8���A�h��#өsP\V�@>a�`��gQw��|�㞝�?��ixa/���ل��:2.:6�#�$�O�d>�)�%�	,���1U��V��Xo�<� �xc��?+͒U�`�K�N����;Od�'�b���4�?Y����� /$$ �ǘb��9��I�'�d��"��Of��O��:���<u���Ey*�(��P�$a�����C�]M�l���	2N��l�!��8#�~��L�;����/@��52��@c�'Y4��}���g��ĵ|�ŠD�p(v%"3T&a�a0��B��?����9O\��R��$a��:��S�i�'�O�@� KY�U�֡��
U
�`�:O`K�.Ym}��D�O��'z�b����?i�����;"�-;�L�BN;���p����?��y*������/���yG�Q,�\A�TB9s�iGx���'Ǹ�s2/��#r"0����T��1!ul?'��"���O��P���B�����A�\��iJ"O��A��@:*�ިS�垆(Bx������HO��$d�����D��p #.�#/2��I֟��ƫG�	�h������۟$+[w?�w,zU���Ne��a�K�ks��k���yQ��Yȝ����%! ��T�	�!�`�ۦ���|sŎ��=��AS� ~�RP볂B.G�xmJ��?!Fz��W&�ZHR���=~At�A6�,O����$u��hg�J���O(���O�d�O���2'C�R�
A���D�+`x!���M�6��3�$�в�R!d}�MEzr��>�)O|����D�E���άe}( ��\(`��C��ǟ(��ʟP�	�e��L���,�I�zG��Y�-��q�$�s�]1�`���X(<$�P$�L26�>��D�v^�];�h@�O\L�(%�P2읇�p1�\�0�zuP��T�'�> �J�F �s�<�����2eB!�D�,d@6��O*ʓ�?�*O"�?ikG΀�.y�P��z"hV2($!�dQ?V��q:!"�����W'w���ܘ""TnZry2C�4c����Ɵ���\����)�PQ�D��\F���h�8R�$���'I2�'��)Z֦F:!�����O6˧5�
�bfpz�2�L�WT4Fyr ���<;� L�V�y'�Bc:����'F)�d��#Ƌ@n6�*M҆Fc�Ey����?)��Ff�v�'���7B���B�K�W�v-������I#4`�_�Ӻo�Y�'���(�%p�+բ,bԋ�i���m`�$��Zζ�d����S��C`��L)q��ElZП8��[���AE2�'0��B�P\p��E&9�t�(�"�
e�|�ǉ�_皴�H�ʧŘ�?cӬ�aYR�Tߌ��i +aw�Y[�l�t�ŤO?���4�vcҁϢH�8Y��,¶L�^1P#��O�un���O>���%�&���8\��d�w).��O����V	AF�P8DB��0��Iksi�C��pa��D�|�'�޲HgL��@�ظ=&�TR`hļ�?i��D�,�*"N��?����?���<'��Oj�B#�H˒�F����d�<H�D��2P�}a�#"Lz�i@B�
s����~b��(��>����*nOp�o�h��;���~���;�?���'���Rg �"D��ȲK_+-"��	�'����t�tuM�`R #��y�#3�S�O\�(c�l�.��C��={����	R�I���b���O �$�O ����^ǟ(�I�|����p��8@�Y����	"м8�L"8$����)W���N���!!@��]��)Q�S	cU���DD,N!��s�q�F�*��ur�'�m���V"Or�)�boĀYd�� !k��"OL�0���!u��x�6aN.}KZȂ�8OR��>�P�A!y��'L2P>ex��ß^� ��H�89^ ��h\	E�&��	���	I��I]�S���T7n������J�Nɪ�#!�(O�����O�l�%�F�d��"%	�,��Fy��.�?��j�1��-W�4�U���;�,C�	$+z`L�4Y��Ȼ�˜'1q����z�&.�Z�yRÙ->���׮���'$���۴�?���IQ.=l��$�O����R$�e�(JP�� �B#QU����O�c��g�'<�;S�]]��A�&�C�P�
�Ã	���"~�	�XR0��Fk�0@`)��mR6M֔0�e�� K>E���¬m��J�;��pԣ�-�0���8lD�0��̟LV�O
 w#��Gx�;��|��[�8��F�G!V������8"<�����?IWEF)%�+��?����?�����4�,�sB��r���#��� s�Ox,J��'W�!sK�M���H�k�C<	�RC����.��D��3&9��T,���:�F®%�	�h�[����6v=��i�� #�NC���ȋ�ًS�H�i��>D�| �Fɪ�j��֭�`�Ʉa��HO>m��.R��M� 2��D
 <�e�3}�@8d�O����O<��L5vk&�D�O��ӢJt�D�Od5���מ6�*���/%	�< ��'�J��)OJ�X� ӧj�2�pu)�0eb0R�'Ŝy���q,�V�K=%Wl�)�"Ev�m�@/��yR�H�!���ԫV	g���5�،�yb$�-!1���a��^t�f�_��y�%��[B�0Kٴ�?����ɖ���7��y@A;$���W@�5%����O���]	Hi���+�|b$`÷j��h2�W�Tp�y� f�'ǎ�C��	��,�A�K$P�Ⅹ7��Q���A��OT(G��5�Vq�a+͒@����M��y��Q�8����'ɰAp��@�Ă��0>y��x��ֺSn@,	%�=%h��cԉM�y¾)��m�؟���n��'Ч#br�'�B��PH]1`��i�B���C�*�v��C�'71O�3��x`�P�<�m�w�Ֆ5rz��'i
��O?��O���Q@��)��d�
G���o�O<c�"~�	�ls�l��ʁ�k}��J��� ��5D�,Ce�����]�>Cbɀ�1fϑ��'z�X��.͋D��B�똧q�����?IAJ6;~XM��?����?Q�����4�^�J􁙮�H�:��	��x1g�O�!��'�=����0��`�*N�L� ���'H`4��t�zi��D��c�V�`�j�#�tX�$��IH�����$*d�d�{ �J�࠻�3D���UM\2��P3�ݓ2��p�".�HO>���V.�MsQ�Ƭ\�x �U�+>J]���?����?9���jE"��?��Oy������?IVk��3:�x;I60$�`�e�@g8��I@ú<���q����(ըu>M��F�f8���4��O�4nZ
���x7-� *Fx��!��B�3��Y���̈́#��Y�*ܜf��B�{r��+��ߺ,�LsG@+T��	��'C��`�`{����O�ʧ��pn[�rޜ��ʉ$T4���q��=�?y��?�5���?I�y*�
����ш5�T�[�D�|�1�w�ɲN{¢�B^�i��)rCD��B`��!HR~�'�,����h�^�S�'/]���EA�Xr�H*c"O��j4��4 ��x�풪n����'h�O��+�P��Fa �G��1o:d��6OTdQ*TƦ�	ϟܕO��=��'�'ep���$�$�J��w��.D:���W珳)b�T>#<��䏢+n��dh��cbd��G�W�^	 ������O��g�Vv�(��R$T(��n�x�`��+�)��DB1Gڙn��=�H�$��8KT�&D�@�VC�u��ؚg#ͮq&�H3f)|����'x��ʂBV8`��Ȑa4P�v-y���?9�����u��?����?����T�4�ֱp��8���'(^�@����O�|�7�'��e:P�A�8H���Z�,
���'I�u`	�P��Y���2�,<9�$_�%#����_騅�I+��=�`�9��tkP�0:$1�N�d�<QUg�&����	</��h奍�*���"|"�ձUt��M��DCp����^�63�xc����1���'�2�'���q#�'Q2<��j��� ���`���i�"T��D��^f:�PA�Fhv���'Nb�����8Td�w�΂�pQyw�˨f@��j��O�8�!
�!�D��I �M���-Sr]��FȄ��I��?���?���?y��?�I~��S���J�*׮u/� P�
�ZY�ȓnnѻ��؎zؘ�d� 8t���^��	@yb�A>X��7��O��|BF�O�mx�B�C�� ��Fz�(p���?���	-��O=8�;F��*����C�3
i<eJ�5{v�I�W�>Ѐ@*!��+��Fl�Ӟ[�B�fӅM���_$ei��<i֦�ߟ4K��i�3K<\�L\g�dl����R�!���ruP�,��Aq|�H�͝A�a|d8�Dȡ2�
)��T39b$\�
L5Y󄅕9GH1oZƟ��I]��	A�7��'"��E?�0�Z���'�|q5�([И�0�'}1O�3�v�xIz�(́6�(��ͤM^(a�h���O?�$�*���V(�$Q*~PXQɍ�
1"�b��O�H&�"~����)���5!,2-�"�RB�*bE�4ϝ:ma�YqCS�n<:"<Q"�)�eN�-D�|�
R��"u��n��?��)�FQ8�C4�?����?�����O�� Ԍ�g�֠�>�h���*C�Z����O�)Q��'m"�"�!8s��2#�J�VIX�y�'��q��n���F�T0/$��j�?B�ʤ��1��i�I*а=QѢic458�@�!b`�u����yb��!2ip(�gQ�X@V�xlG�$#=E�� D�6��6hH"B��O�Z���@
�+����O����O�4 cB�O�p>��F�O��dx|�Qȗ���
��aꇑc�|B&���򄋣p8�yVh�,l��l�rg��w�|�%ʝ�?I�i(2�����PQH��4yT��'[���C���ݸ Ě+
�t��'?J`�c�1d��:0왜?���'Ϙc�h 锳�M{���?�+�>��eW-VJ8%�S�^v&�a�lT`���O,���1���$6�|b��}��`�LB�,�^�9�)�p�'��B��)ЭlQ��G�
�a
���FIQ�Ȱ$��Op�}���*�4���
��)3 �)��]@�<ơĨ;e��۴mN,.��S$��R���J<A�܇V��!g�L*��P�P�X�<��ꍏrg�6�'�X>a倔ȟx�	�9��޿^�M VH[�<�7	��2m��D�S���DL1M���pDጕ(R�ԃ4AӢb�J����)����E��7$��o2gb܅Z��J!JXt��ɂ��S��?10���.+��߱(�z0!@��g�<� ΁GT�6��3p]ιxa�'�<#=�O+����J����24"F�Ip�'���+bζ4�0�'!��'�"�sݡ�i�uȧ��y-�ɔ)Z[����!�N��?�%��L�nu�g)�	0�3�hg�(i1Hƥ1��`�A�Sb���5�'ĺ�; �vS�1�&ĂCF{��G���aA��4!r
�V!��~"���?AߓR�A���%`����F��m�ȓ�ĕ��"��(��H FU�7���g�)�'6,rt��i���ڕIġW����s��9�}k6�'�B�'W��	-`�r�'��iL"-���'�J��pd�q�B5��%6�2�-����'���7�DP$���C��^w�I ��z�����M���t�\!;$E�-/�t���c�<I�3�8����L�*h�$B�`�<�e�
.6lKcd��E���<Y���^�Ao�,�I}��OP�+Z�M�҉ �A��ܚ�\-Ŏ���'���'hNi#�'P1O�1i�L�����u �k���:2�&�<a�h�O��9(��H�e$9��F��B�q������(�'y)�4J��Q-n<��YĤ�E]2ćȓY�-��8�~Y�-W�/�ި��ɋ�ē(�p����@'$�� �؇%���&dR��IE�ԊF?�'1�I�7�J�ԇX���L1@��@����{\���JA��~*��b>�d�T$��a�Ȝ�o5��tAװE�6$8���!�i�E%Q�}p���O��`5aߋlU��`�{��؋�LK�WZ�ċզ��(O�O[�$W��,�8!?<䙀�n�� (7D��ⳋ��L�I���c4D �!�w��D��OZ�-EX���`�,eI�8bu�¹���'ךL�E�S�P��'8r�'H��]ß ��'Z��$W���
8����IU���	)ejvU�bK�|�Y'�'@P�"��@?�T`,�%�dɰ�'��۲F��pAҩ෍K|�ܹ��H;}�Ł��¨I�|Q�%���c'��O�I��\�R|�&j$W��5/g�B䉃<�D9iV/�i�M��I�$��3���	P��1��4[��=���߰*�ɊS�،9Ա����?����?9�/P8�?����$՗�?��h�QPv�ċO^,�À�?236x��ɒ5� �*�P�"��-��%���X�.���	�a��d�禡X�"Ͽ`�2�1#c�6�R�r� +D�غ℅�l~� �)G��>$I��(D���G%��JѨ4H� CȨ#,b���}b*b��7��O����|�VŎ/9~��6D`�M��w�:����?��x��IZ������l x�@4�Ƌ?P���0 3pQ�,z4!0��̲}�@��_���ik[7G@UDy�T��?�W�S� :pM��H�%T���v�7	�B�#b������G�z��F�9Y[����O��5H��]S.�&A�P��F�W�7�"�	(B$�lܴ�?y������o�����On���D¨�0$��j��U�3A���,�9�
�O�c��g��� t=Z�� �̊��_?�xrD2b��"<E����F5��F��Lm�t�>�nˑ�T�?!�y���'v��q�I�Qք�
7C�t�jD�
�'�6p� � �͈e�A=DEX�Y��D�t���)�+Nh�P�ȋV����e��+�����O�q:7�lk^�d�O����O���;�?�;CFf���ρZt\�PW�F5Yv��l&����ʝ=@-�f�Y[F{�%��D�0��ϋ�-y��`��%k��C�J��0�c�	.Ô���hO�� �٭N�֌{�hQ��K��O`e���'�j���8q
����ϻy�ipA��_�!���0	Q��� $��� �(���Fz��IN'h�UmZP&�� hZ�D"|͝�e�j��I�������sp�ߟ,���|"�K����I��ur��ڱkf�5�p��92���]��	�A,b�JG�a�����Z0w4�����j��Jp����'�4��CGْǸir�"O\�rd�OI�@��U�{�^}{T"O��!���j�vIp�_��X��<Ov4�>��	��̛�'�"S>=�bC�p��)A�C��>q4�vd�sF,H�	П��	�B(�]��d�S��ˠF��0�* 1D�RU#�/���(O�ՋW�8{'�L�0��rh05ST胡h�L�<������G�d�ŴA}���Ó����c�"E��y��"�p����I�D?R��Tϋ��0>f�x��:N��p3č;P}��H�C��yҦ��vB�6��O��|⳪P��?���?�i�+/���B�U�^V��B��Bט���Ԙ���� ���p��T��m"�%��}�0�8PN�S����"�)ـG�W0RF8i��߶AR1���'ux�O?�d��_���Pd��s}��h4l�!!��ʄ-#�pC�]�w׾��6+��g��xh���?yq�� T2�E��_?J�S $�ǟ|�	��4P@���L��؟P�	$��9��l��%������ʆ�^D�r�O����Ŕ:�{�
��/B�2�.Z6���B�d�-�~r���G� ��	vEh���]��S!m�b#@A���rЊ�+��?��S�'��R�Р�#ƍ7j	���ğhU�`�'�jeP���Cf��1��L�	��mK B)ғ��<�3Dn����3�<�&�F*��c��w�����?����?�FG��?���������?��� H�e�D��7�uFI>|@H���ɴ:�8�mr��1�ƭsʀI�W�C�t��I�\����O���NP��a�Tz�`�sb"O��A�(
?-c"L{ �T<D�y"O�ո�'P:I�c���aq=OtL�>��`Ě��f�',"_>幓dZ�O�f8v�%o�=E~��%�������hAUȟ��<�O����fo��Tvx���H��	u|i0��$_%��?�b�
�.������nڼP��"ʓv�,���H��<��V�U������B�c`��a�"O X���O*9`"���B�j]Q���'�O��9������"'�(kG�`�1O��)�l�����ܟt�OF�<z��'Vb�']ֽ"�׆iؤa�%�-�l(`ф ���T>#<IF�I����E���P�Աp�E�d�Dɋ���O��Ŗ�����"ٞ��HGK�c[d��o�)���p���+�� ',��[ x��f6D�$륎��j��D.��W�� G3f���oY���ҫ�5���S6��7=f������?���$z�I����?���?A&����4�eI��?}VQ�6�6?h�Q9��OrU���'��`����xBC�$����'@�h���N��&횗V�"���X��i��jӼ|����=	1�@�.�e)E�ڀYD#&c�K�<)%��m� ��ȼDN�x̞-]��"|�f�ѕS���beN��ȑiN5� ����*/��'��'T���B�'a�;��<`�'%�b�?��}��P5���F]�p>)� OAy��M�b�P�2kT�nJ���Y��p>������	�Lըx�R/��^�M�sO���C䉀a�
}Z�ңe��		����C䉲EWJ�Qu�^�`���C�
���ɢ��'�`\��j�����O�'ye&;��׭}Ӗ���k�D�(�S�_��?���?�T��)	Ej�2�|*�hD
�+�H�A�3��;|DQIv�^K��J���A�π h(��H�1Uf} �щ)	h�r���-����Oғ�f����8�@b^3/��If��-�p��7�)��<��NS?1 �S�0#�ʨc�Cv��2I<�я�)��]��a	�>�ʥf@�<�E*�[��'��Q>%��W̟ �Iן����+]f�pz���g�x`��J[�P�,�Ig�S��������� �嘅���s��}���7�S��?p���w���:���5 �`To����iZ��ʘ�����G�  ~���j�*�&�A��y�*^��\�*����[�,�����O�IGzʟ\��"ͽ� ��h@�N��8��O��d��z��w��OH�$�O��$ ɺ��Ӽ���C���P�H �v�!*k?�eɊ{x�<tU/��A��<B����.��\2K"�O��w�G#���8�e��6n 0���O	�%�'o&��d�q���˂�	�>4����>mg!�TybCF`�'x�A�2� JZ�<Fz��	��Dd�m,5ѦT��ѿs�Z`(�6zђ����������;�H�����|J��H�c�D@b�+Dmq�9�	&1�xu�6E�`@�塓~��P��)�>V`���Ж'EF�˱�K�H���Dʷ;�� ��*LO`m"t�'t6�	9V�l,��Oތ,P���NV|�o�M�S�>物
d�:���a9&yz�"O"txb�6b�I;��՝&� Ѵ2O�a�'�1OH"}r�%�f�*�#C�(n������_�<�c��n��lہ�K�i/��s��Y�<i��+,�v]��=}IT��b��S�<A\xRDz�`Ʉ�����N�<9c���pO�]І�R�|[�(Ce�PK�<��@ $�y��cߡ)&ʡ�a�C�<�C��:�9
d#f�� ˕Hy�<��{w�@3�X1f�䪃f_�<92/ËPE�x�"��5��:f��_�<��oڴ~���u���U�*���]�<9�`@�z4���4ᛧ.�Ƀ��m�<Y3	
�r�>��@�D��9��j�<�w#�0d�a���i���IDD@�<a�٠I�,L:RcZ�k��Y��s�<�GN[�h���+;^ư����k�<��W=K�`�f� )uj�Z�nVa�<9�I�~
~%b��D�Q����b�<1������4(�<���َ.g���ȓG
�qP7��*�8��Ț�A���$(v��ktF�x�\)$(��.�B ���A�>�[%�փA&ܔ��N}�i��/C�!��%���r���TC|l����>K���+GO 2ü�ȓew0U���ݙV�T��A(	�-��a�ȓ�q�r��11�|�LS�[>��ȓn���2PJ��(�����Ǐ�lxl�ȓX�¼��ݽu��u�R������A��)�%܅�2I�1���<�H̄ȓc�@h
��HUfؼ���������@���X�'K|�=9��٢{����	�V����ØGO"�3u'�F�B�ɭP�X5�'�[�v��[�$�0O�2➬Z�N�<�n�D�d�M��ā�m�2��2�ǚ�~�.<a}�����P�e!��b��$�,�l\l@�C�u�IXY1�
�K��~B���mix�Q���]�I���X��yr��,.�*�k�Ê�M��(�D��.������ҟf���buv���S�āֻ=Zv406dְ4�FوT�V��0=6cH:#lE(a��������ݰ��F�/Z��k �/�B��^�nY�E+�w��s���E�8j;΀�p�I�g��C+>�I�'�
G#λ�Q?�(��ɵ=H� ���!��!1��}�\ه,;�@�V�'�ڕ3�� W��3�G%C'L�*åMS |�ON�Q���
�	k-����,A&p�Ç˜-�L���p���;���CK��L��0�'Eި�Q�O2��Z>ӧ���a�? �yr4�˽8�H�� ��k���!��'$�{�M�^��)�V܀�¤f�֭����#s*��Ff�m�����	M���=�@��.$� , !��07r���@I�w��
��P�LdJ"<��Tǚ���=KډX-\;	C���~n0�ӷ���UQ�����;��*V-R�7���yHG�p(�!U�ڀ�O�'0�� �'
&�P��߲h���!���NlE:�N(��K��l�8뗥� `2ژ�%���n�Oڙ�!��F@n˓.��Ȧ�6dA䏖��J�;%F߇!]��:CSs&��p��N�5'���4�[���`Hf���L��/�޽�ëQ�R��rl�Q���0-OL�I��ۑ=LF`�g�ę7o��h�D�8 ��1��U4h�a�FG��znZ�B�N?fQh%r�H��uG���R1�b�0�ы��]���(S�ϰ -�Tbf�;\=��QG[�re�	��'V����Ÿ&P	楈 sZtQ�h��}\\�im �$֚I�<i���;#&�a�w�ӛ-����y>����_�3ۦo��8����6tJ�*���O6uV"�/^��	�m�XwAJ��C��_2����N\p��!�2�H�#�d�'��ā�?� Eq�K�>i�b���j/.P��FV/X7� F��7b��ad(d�	B�����`�8A#'��[���	�/�eVTE���,��D��Gg��Yb�QD-Ɇ�\4:�t����y)�S̓8�<��f�<?���ӇB�(n*����L�6���c�*��{r��/@|��)2�\��&�M'�y��ѷn.�`���j̓��Ͽ�P��m��IG'̝4�*���a~Z�b9�T�
�|Fd�(�P-?�j�  �2B|�y&��"�	����I�^ j��R��4�ƈ�8y��:Eǐ(r����'j6����.��O�A�;zD���5Z>�d�]w�T�KQ�֔:
4��F�D#���Wj�P�zM�$�Q��C0
ب=%6�����M�]c�mU�w�p`Z@�H�(���
�/+B����":�rE����Ʀ}#vmT�s�pA��Y��y�_n	�G�N@�R󑈅�q��T�H9�Op��v��%�܁�%m�+5��8��.���Y�4T1��2!�#@��C5O��'�0Hs	u����X6���OF-0� ��O/�O����K�d�nM�F��&=�R��dC�^�xK���o|��$�P�&e��I��$tnL�B��}�ddB���$��L��,� �}�Ğ�����z�h�'�\�狨dv�d�^�����W�lc��	p�[��R5���Z�O3n������@G����"E��Ot�;#�;L���o��j;�T�'R�`��8k�T٥��Q:�Ok�t�%��ܦ�9''A�+JЊ�aK��R��$��te���4�O�\�3�]�@�r��W뛎s��ҧ��{�����_t��!H�<9���oZ� _r���O�У?� [vN�u��9 �!4�xC�'^Ƒ	�d�i8�i�G��pUT���eӌ ňE�#�4}yd˓��!��h�O��0�T���]>�n�1IE�x"bQ�"���_Hr#>1"�X2dB��%BL�q�����
YΟ$i`m~�x�ɑ	.�Y�M��FV�P�ɭ'�t�B�u_T��'>��<I�K�32��A�C ._��!B�<!g��14� ��
1Y� �H�C�ӟ�3�ɸX�h�����l��yX� �)-����!�H?�}2%��kX�O����̍&\D�ź\P�;�?L�����ĝ�ZP�9���?��;���$mю}��醣
�~g��'��I��Wu�'}��+F��#p J��C�� n<5p��ÓO���Z��$)JԂ����;O�>�"�NQ�u%��TL�R���aJ�F|B��	j3�%�Gk��)�ꑰ�*\	�y�kɗ/��Wh�$N��钴��8��DL�M8\��C�:.c�#>���۷8nj���M%&tYC��_}���m\4Q�EiR�u��I��Oߍx�j�F|�牖.���S��#�0�څ,� J��i�N<15X��~r�;z��=	 ���g\ ��_7\j����@bh	{��b���1Jй"��>AQ��F��w���0�	�~B���t�L�E}2l��)�L����/�=[T�+��t���P���O���vlP�JX�a??if)\�+�J}yc��70B<`�uh
E�'M,��v�E�o�,��N�',2L��'�<����<{�����q8]#+O7���	y~�O:>� �s��rz<����bit� �b�m6�Q���y�N�/`����bk5pL������O8��נ�~6���,�7f��,�')����W�o��iT�K[����=���[�]�d1zW�d�Y���\��d�aGC��ϓr�40d
<;t�$)�H�i��x*#�[#���G�Y�"
ģ>��A�ǼK2��*�zAdL@:�*mz����'x�����E�T�$���ō�N�xD �wS��
�"��$�Ը���ȉZo�	Γ}�
���I�&C݄�!�@O�i��'��"�)E��J� �:���Ph�&?��(Qg�f�����Hg�l�'�O�R�v(b"���}t��T`%�Q�q&��%5��,�AnP3]���<�Ef@H�����0'2�YP��?�+JԼ��S��9�������1n�`��@�ˬ~���f�:��˚}���@`�rI|��b��Sܸ�ۣ��.D���#��Ɂ+�F��2��-CaٳYд+%)�}� �?���!2�0b�Vur!�_;[� 2�KּT���Ƣ^"�$�i�i{�� �i��/���[�lB�Y���$[�dD|�HȪ'��͈1l� Y4H�3��B��H�C�� ��x��m��y"���x�>��ZV��4��(��O2�3S�������L_	@���C�DO"I����G*Cs�>Q9t�ʸ',�A���T�����������	0d\1J��N�J�	�ʟ,�I K�Q�*	�d�t������"�L0)��H��Q�L�Q�P�e��ո���-h$�x��#~�!��9��B4��	MԔZ���!v�����͏8:V�B���+���l8��7ǋ?q�t���&�Bl9Da��'6�$B7�ѱT&F�cv&�v�'oRM{�a��#>�$@3����F�ͻ{Y�$K'�P�4�dYVU�H�"]��/ے2(j���Hڝl�����ϸ'n�I3�/�����+�N�!Q����'�l�tg^;p�� �lww�ѓ�W����A#ŀH~�g;<D�H�8�QۄOF??���G�x2	��zv�-�g���[�B� #H�C�I�G^.�K�i�	Ⱦ�RCΜ ��y��Ҙ4f���J
e���Kƀ1�/�x��ܫg�`IK7B �/�� \��ܝ:�
��4�����@A�'�!̻JϬ���j�P	���Բj	���p�Z�'�>��B�h.�t	�O��_y1�͂�k�5.���X�'h��WG_u���XuO��y�~@��10j���G/[=q���$a�TЙ�yRɂ%(D�ۅ��M~⪓	B@��7V�_#��_�HL��(�n�<y��p�d"�oF�s3���%h��+L��'Wftv{�K�\��	�[���1�×@{pa���3_�d��5�߬��ė"6d�@qc��fp�^���`W�����F�_h����:k��a�Z)lB�����^ax���Y32������9O�,Y�eB:>�\�1��+��æܲu�&���+ڵ[C,�������~2->�.�`��O�#�n�)u")�o����X"�����
�'��\p���)l숁�šOa��O0�JgoOTn�}{�8O>��sR̺���� y�8�v\`c�+������T�s{��K��',v]b�F*�q#���8@Z�����U���U���&�/l���d+5OB����S@�O�PQ%�N;y �0*W�J�MWx�RU�'���ǭՄo4V����J2��	:��jJ��i�(��	@`p�)��3 ���,�}8�p�E啺�p06�L�O�h���/�I�x�@4�%�ި���7�N�^@+�q�A��*���¢\D�D!w�F�Z���V
O�h�H�l_�U���V9W!��Z흤D�����@%H��p.���Ni
�@�(,ߎT��OI|˚wr�$�U/Z5t���q�Q�z8�
�'��� ���1�R�@R���.��H��̐D��1Y�+u�ت�F�;��Br��U?��CT��M�$ƨg��d��D[�dy�� _az� �i�"�	gHM�O��A쌨?I��Z�%�a�8m��#Ԡ:^���H�u�2�r�Æ?�B��	�b����@�S�b�h��w�b�� `��_���kR��i��y�"�FIfi�w�"}��P� o��Q�r��0YxC
>Ke!�d%C���)V�5p�Tp4��8e��ppf[�\Q�$�KP5'S~�l i���!Fp��o�мC��,e<�@��\�{Vt��aGf�<i޾���ye	f{q/��6�p�:ҫM�#Y��a4Ct82�j� ϜC}��;�m9���'�i Aʖ)�Jd�vDS��� ӓ%�"py&!����y@�P3ip*��q茹
n�����)P��� �
�}GN���.�1iY�� ��8O��sD�<OH8[�ᄻW��,�U��̉9��h%�!
�`�{D��"n�\��#jɏY�8��k��o=t�r���iN�w��
<6B�	�lh@Sc��0������)0䑋V�61�ʀ	EÈ9l)>���O�,�hAQg�H�	����&�зS�,hg�T�#BoJw�<��XC�$G��2�@��ƞM�42 �Q2 �$�C5',4����}&���E�^
j�:U ��N9CD�3D��UA�l7:eA#�۩
. <�˲>��!:1]NTr�!<O�%�d΃�Ԛ�����gjlTk �'O�٪����Xȳ� >C�L項I�T��Qbl�eh<���H^הb���h岬� ��X�'T�AIs��+�0�Z�fֳ>�*e�&
R�W/d�	R�W�<�sт�.�B�-Ɓ}VR<�6I̦!X���%��:��>E�ܴc+pP[�(�F,���#�'Y:�)��7p���R��7�����C�?uOh��'��;��G�^�����ɼ@*R��FM&JaB�!�n��&����d��f+��	�*U�5R\��C�8C8x��dL�s��B�4}�|�x!��- M�=3E�4%n�C�	<'*@��#_*a��)A��.��C�I)��	j�G�?F�����F�;r@C�I�A�VEK2%A ]�>Mx�á 
C�I'�
���/ǇJ�P����S��C�	�bz�F�>E"ś��K�;	�C�k��q���/��,	�	7"aRC�	�"�����W�w���07���j1NC�)� ��
Bb�}��:tG��hSB���"O�`ґ"8�2�O/�F�"O~�S'܎ZhP��%�&"�"OZ!D��(j�uK�.�5;\4z�"O^���Cء@����� h�|��"O����&	o�*LZ��R�t����"OZ��4	�8��f�-A���[V"O`]C��F)9nZ58�#Ք�����"OҬ�%�V�:��$��v@ڵ"O�9��F�h ��">z����D"O��0%Ǎo�#�g�� ���"O��@vN��(U�������	��:v"O���cÅA	,�WC�
�b�"Or S�G��K"~@AG��3I�d݃V"O�@y�T�[�Q�t$�)1�:)8"ODɗ$SԠ���>��<�%"O8UkF��%xDn�k���p��T"O�$���
�"�9Q�Z1��"O�xP�a�p�(s/�D���b�"OL�Q�
�Vg2��#�3U���V"O���nM>�V�SU-��o�&]"O�I�S��	O|Pg�2��,�Q"Oz�`'K�o�EB��X�W�b���"O���BL�	N8�g#�\�K���yJ�#f�`!��,CD�:�5�y�L�_hL�i��H�V�����	<�yR�=\W�� u�@�Xb�Ј�g��yR�ѝo(��b���Qъ��7�̗�y�4?dܠ 4�_�F,9GA˛�yB��� �	�hT�+����?�yr�V�$��5@�o���A�6G�yR(��:8�â�� ��h&_��yB	Fp�� ��vߚ�Ye����y�F�E{N����^$>����֭�y�MSTq�Q�/A-E?�!�p%B��y��B�$̍{ 	ζ>�x���&׳�y��7X�t�T�W�a���b���y��+�ȵ�q�V3'@���` ټ�yr�'>U�u��F�:.@�1"��!�y"Ř�S���3C�-�,p���-�y��6Ǻ9x��҉O�4 Yw��y��+st��'�MLHɈ���y��ѫ�l
3)��E�lS�Dѣ�y��J%Q{��/ټTP\U���y���#���B�G[�U�X�2$Q��yb�R�A{P\�v(�N���B�hJ&�yr�X 0j���$nC�V�*)@����y�X�\J�u�u�Z�7`��j%�y�6'؀#�W���r�F]�y��R�|r�$�t��u1a�B��yRF�<A�:�"'�a� p8PlE�y��Ɠ��a"�=Z�`RV���yb��/F��vdHF��ڦE@��y�*<K2�x�@�?pt����֋�y�-S�\�{�@G�dDX�2�铑�y�FS#�.���!��lG0�)�n��y�ow<�Ue$w�{a�G=�yR�޸{�d�S��$Y2�2�����y2��k�~����A9|]f4ɤ �5��OZ�~�E	�7�����(7��TeLV�<!6 �	�I�"_Z �a�ŵcG��zP�a ���vB�!:4P'�y�k�3)<�ǡl�.4	4ђ�y�HE�"v�Ͱ�+�j�!Ѷ����y
� �E��UU��1�QM��]e&��P"O�xY�c���Y{0B׺FV���0O��=E�􆃑a�&���cG��aB���yBJ�3L[�Sv�\6}m�]�@f�y�J��Ĭ���	��=��"\��y�.��S���r11pX��	��y�E�wU����,��W�T������yR)F�r��ukS�WZt��c���'|�{�E�.^�ʰ3׍K8QEs�
�!�hOr⟐�O��H���<y��
!e8]���Z�'�5��	א�)3 �)Zʾxش�Px�ȴUɾ=���Z�>�ԛT�Y��y��$e@��%�;j� )+D�Q��?9�)�'e��""S@�� �0��9|���'�|��6CϘ
ꠕ� ��2�3OU�"�33�.�8���>_]`a�Wj6ғƈ��*$���ZU.	/���$��s8��0O^!�q�Ǎ=t�p�D�<O�l�$"O.�@��	W��$�wDД����"O0�k%(�.V;�HA��-���"O���vk�kv����1c*ʐ��P�E{��	�BP����)JьTc�L��4�!�$�+.0�y��fP� V�4�*1R����'��>���|�lh9�ɓ,YZw�7D�4CC	�f���bţ��2D�	%A��`�,��bC(��HS��0D�t�$	�8|pqiV����s�O�<��'�h`�c!PF�8�'��',-�����d�
��FI^�8�����9Y�C�>YV����R��4��%��#/�C�Ip`�}E� v�nؒ��5[��C�I'�0m�嗓 ��ià���:�7m;�S��MC�̋�iOpu��T� 9�=sChVw�<qDHP.d���8q��0Jm�<��˝�Uftt c�02x�+�j�<�%Hܺ�� ֆ<r�4x��_�<1�%�&��a��݃i\	.D���$�@�r`K2M��1�Zâ?D��ٿ-_rL��k��j���IW���~��>�~�1N�
I���PH�1qha��MK�<qW�ץs���Cl�.O�� �E@|~2�'��
�>��z�L�d�0I�O�c����Ӳ~����W�O�*�(2n��Ff���0?�aC�3L��U���B�%��Bj�<�c H3dP�Kܫ]���aGFa�D;�O
���l�$9P`�j�����"OP�@��޹g�|��s�O:O�h�"O(Ԑ�&/�Q�h"=	&� �"O4h�� 	�2j�,e�U�?�BPpC"Oڕ��hӭG�
�Xr��R���""On8rE�ߞ`��"a�G-�`2D"ODЁW���1��Gj�6���H5"O����.Ü�[e*���0�|B�<|O��zGOу<�� P�*�9%wl��V�'�V�"	>pqN��O΢P��������ȓd�`1f��h�xce&��_+��G}R�ӡM�L���7��9��#��B�%�*�!�FK:��-{���h7��'I�f�'#�����$q�R���� �a4��	�'%�����[�P}�4Ȃ�b�8,;�}��'�r<�3/��w4Ju��턇J��-*Ó�hO>ɉ�o@��؀�`ŝ�&`N��"O�J�$E�B��oP�=X��7�|��)hn,i���Ͼ�s�cʛa�8B�)� R��d��AB�-��M�0���ۄ�Iq}"�I5�>���o��z@v3��4F�����>��DC	|��q�fΛ�N�&�X���U�'��"=���y"t���Bb��9���@�M�8B�	=� A���l�0a0�
 ����<Y��ԟH��GlH�c4�ĩ�D:[�
`�⚟�E{��S�"P2���(s.Y:�H�-8���m}R�'�v�FƄ�_ ��跈�40����9�S���v*f��l�r�^ѹQ�����IX��ɀ��#jᆰt��2�(����"}R�)�����I�:`��R�ǔ9}B�I�'�\�r�#�(^R:�飦�c�qO@���?I�,�/߾x��L�+l�q�#�x���ΓmTQk!@	�@�AK���Q�h�<����I�vH0\�~��,Q ȴ5���mt�x!g�]�D�T�Ԕw����2��|���$j�;�%F77�vyS�GH^B�'��O���]V1(��'T�i��e���'���O� ��J%OH��F�M*����C�W~��xb� ��ߩ�pG��lXS�K�bS}��� D�HjXqF�Y���<pF�K& }��)��n�2�(���q��U@����B�I-9Ν�$�-9~�]Cb��QtZ�D7��qS��!<|�.T_�(��-%D���ǆ@ ��E�6��)!����g D�� � �$\����C�R�½	T)?D���g�"�XPӪ�+Zg��k4�8D��a!��"N�����%d��rd�6D�t����a�X�" ��kΨ�r�(lO���yčA�-��"Rˢ.��堂n%D� 1�ٕs�l]�3��^~��h"##���HO�OR�Z�N�9qg�<�����t�	�'J���h���9w/;#`�a���ј�0<����z�lE[	���U�fB^�<�ǭ%?���R&��n��P���ݦ-�'����Pm/5`ŉЈx�0�8�1O:��kI�v,:�+M���*f"O�T�Ў]nT�:��F�K�����9�(O�O�|\kq���~��"���T~�Q+
�'�+f�Ť��	�kh]A�H>ʓ#�>�'�O�ic.���\˳m <%�� �"O��z���<����,�g�}Y� ni���O`%��d́����"&�"I]x��דK�f��By�J!s��� ��p�1�c�ސ�OT���d��F잨1Ȳ�ۃ���~c!�$R�j��ٰ�ۧxX�	q/K�!�K��Ց��J
z���Se�ݫ.@Q�PE�d� �Ȝ�Ac�8zB2tb!�˂�y2&˗D����L��u�b�"��֣�y�"T>N�]�$�
�o�|!Y����yr�B&�GKA�[ي�R0͘��y�g�=S^�Wn҂U���ѤE��y¨�~A��S	��M{T9*D����y�ۼ��uz��(؄�8�(�'�y�
�"R�����N�F�Hj�� �y򠇪r#,d�A�8�8�`����y��H
T*!���L�f�,D��-��y����#䠬�,ƨ��ݒ�c��yҌ�2�X% ��u�9�!HE�y"F������jϞ�:�L�y2ᆣR� �h�Q'Fx�P�M���y�&�cln�K�H�y~V4 (	'�y2����t��b(G�"����nG�y�I:Y6ƩgK'ͪl�c�y
� �m��j�!{Nd���;y�̰�"O�p���"cN��n��j-�"O
��Sk�]r�� ��p��@"O�8�a��-n�.��D��0R3"a3�"O��sn�;�dz'�����i��"O���dN��2� �CDk�0U�g"O��aJ�B�JX{� +"o���"ON(��t� x%Λ�Zs��U"O2���˗�mx��Å�c�qT"O� 5	?6H0��,�g5�u��"O�8� �6sxB���2o�T�A"Ov-0��?I�2����A�D�4�"O@��0��M(��3���&���"O�����\3|ؘ��	�ȑ"O|� �E4.�^-�B%��U#d"O �cQ��ԄY�ҩ �t(R"O��f�ƞHY��0�D�t�rQ��"Ob���$5����K6v"�"�"OȔV+�%[ ��ڔ��%8i�t"O��x�c��-D,�
���DL��R"O�	۱a��H*�iש��	#,D�$"O�m3��ݦ8�r�I��w"%��"O���a/�.V�H��hےB�t�Z�"O=X�e�)L��� ���O�\r1"O����i�c
IZ��2!����"O(e�IY�`��Q8�
ˇ!Z�E��"O���@Z�[*
��g@
 ;¤��"O��9Agۣ>����,V�
�ȬR�"O�x΀>�Rl` #w���s"O*�;��/f�B0�J�'q��xv"O�HJ��
�q�����S�~T.�p�"O�Qځ#^�0و�(GE90�m�"O.xᕄ]�BK��- ��"u"O����F�_�́�o��tI(�"O
<�劌�^��@�!X�����"O@u�#�#%Bic��S�i���8�"O��{D�O�D��i��li�$�"OH����W�.2�Q0�l@�L���"Ox�[t#/���0�K��Ԩ䰐"O6A�	�H+~=����$�!"Oބp�X���cl0:�0mh�"O0��ܰ|_�5jT� �*�8	@"O �a"�a�=����G(�n(D�ܪ%��a��YƝ�>����"D�(!Gf���� �G�!8�pLK��>D���ٕ*�����W$(��L��'D�L�f��,$�H`E�C����('D��`
Z�Jn��W!�.z{J��f2D��˅J��}�8�c��
B,�X3�.D�<��{�ʬ�Ah��3�@MХ�*D�@��)/N�AvgK�R��1uF!�Y����1HZ++h�y�	L!$\!�$�n|rY2e�r�J�x�
-rK!�4v�įQ8e�-�b�@F�!�^3l���-�1*k����,��EW!�$E
C��3�d,`=d���lB;!��ܻZ~�M�q��R⬚V��b�!򄙑j"��)����mh$h\[�!�DY�.�HSNְ,��+�ՔzB!�$�MzxY�fӉ��0�6-35!��ٗ$��1e�B�X��Ha%:�!�DŘ"6*���ξu�xmk&��5�!򤁠>;�p����3i��9����B�I6:�P�j �9M(���ƌ��B�)� ����J=>�)i&�� l�ٕ"OZ `Wc�+�L���Fћ4��su"OT��d���d��eW�	*Rt"O84BÌ��GxZ��JL�b��LA4"O�YX��ڦ^(��C�~�2�+q"O pˆj��p�3n8P���p"O�݃ѠB߲=��Ǵ�t	k�"O{�F��P��P�zD"OHᒧ�ݫ ��:�h���|��"O�!0���^�@d��l�+��,X�"O�XB�@��`�ƜC��X���"O����J��7���s�BA��
x�"O�@�kҦC�`)��3x���"O֩r��2��;��6DY]�0"Oh��	'R��Y!S��7$O��:�"O��Bp���"���zv��.;
T{�"O$��c� P��[�ְ(*�R#"O���q��eC��c�g�  �Q��"O���&E����H�G���P"O�\��D>Rn��GV�/|x�J'"O�M#� 
4�9B�ϓV��(�c"OP�B�o��HZ�3P�@Rݺ5��"OX���%�>[�I���O��, �"O���*^2�����- �K��\	"OD���d_���9�B��
�D-��"O�A�֍LMfa7Ƃ���z"Ot	S�hU,@���S����X���d"O�i�/By����KM&�]�!"O���G^�<R�"�56@,Pg"O�p`��K��H��@�!2��m D��P�׺}�@�RFް�`hy�)=D�����W5bڝ��υH��- q?D���!o������-�����4�;D�̈'	�J�d!۳���st!��;D���t����%��^<r[-=D�+d�U9V����cGÈsǂ���?D�xR�&PqP�Se�?r��3%8D�d�
Z	�B	��?�.��r�7D�@�(D2%���gF�Ȱ���5D�\
�o��m9�)�3EJ
B��dӱ 2D����ï	7�\
�(��bʮ\��5D�8��El�
��WhI|Dx�`7D�`�w+X�Ȓ���ߥz_F(3��4D��	�&Y�NB��cuA�8 �Fl��3D���`+�)u���ר�<�\u˒�,D�(�s'�"5"z9�%��YG@ղ��,D��uDI�5�\|�b�%v�F�`�>D��:t�G��Y����� �+Di<D�ر��;V�0�2&�Ǿu����E	%D�ha޸.�z��C_��1pf�#D��i���#Oll�#s���:*r�Q�� D�,��/E��*�I��3�!�J:D�ThQ��L������D�2�P�8D�,�7��2^�H��,yH���G'5D���
�X�.ȑ��T��8)U(1D���b�ؾ �0���Z|�J.D��"Y�=�He�l9� :�i-D�p�Wb�;8|<e�<���!6D����_��8����J|���F D��R"H�u��)rAҁ]�����)2D�t���6A�<D�ɐ6V��3V'5D�|��]"�@=/��E*jL�C�I.�0��IO�XYu����C�?uQ�$ ��_�b�s0m�t�^B�)� L�kbh�4�d	db��L�����"O�m�JW6�ToU�V��(��"OH<����,`|@��B$�<0I�"O��Ն�"0G��$L��mr�ё"O�DȒ �B�	W�^<eP��"O��з�G4 �-�g �g
D!c"OR���[�=�H`sG�.U�)h�"O��C�R)2�>�{��Y��͓"O"��K��|�t�e$��J�����"O*��SOB&H�qQ�\�����"Oh�k��#r��
��	�x�'"O�����K�^9���E�r�� ��"O:�׈�1:j
��$��x��M{�"O ��0���0y�9�ċ
.}��%Q�"O� U䚮 � �Ar!��)�<*�"O�]��	6��Us�� A1b�"Od�)�hü%�z� ���y��	å"O:�#�.'���9` c�� T"O����ҭ1�0 �'��"Or�ҏ� 6?h�r�o��\ b�@�"O:ܠ�%�JV���?
�6]z�"O�U ��Q�5������I�G�Dy"�"O�Y�0��HN�*vE�3F��Ē"Oeã�ƑS=R�p e�[�֨K"O>Ek(ھ*��kS�I8B���"O���a�=�*E�C�a|�ѹ�"O�� bΑ�y�P$4�mC>Ĉ�"O�k��ǰ�"�Z����2��tz�"O6H3���w����I�#*��P��"O�xqF�[�~����ʛ*�]��"O���"�j�`(1�)�?]�<�y"O~��ԃ�����DƉ�j���a�"Oj�x2�h��hk�j�y�d�&"O�S��]$s�>e0���2���"O ��)0��r@���z[�Db#"O&��� ^�X����C��KJ��"O���g�6\(5��@x*p�h&"O�P� �F�8J�x@מ{6��#"O�8WN��Ck���Bi�;��@�"O��[@�;���&�Gi.@z�"O�Yz�ː}n�E�v�ϻ2V4(`�"O�9�e�M/hT�d��mN��`A"OƑbn�1��(�ʉ"[K|]��"Oh�;�mHY9���i��H�3t�|b�)�ӆoGL"��L���"��8,��C�I13&�<��\�J�Jr♄c��C�I��f	i���^�|�B&Vw��C�	�z{.��`]I6������C䉝t5�%���y����� ( f�C�� ��u+&�~Xx��>-�fB䉭v���Ǥ��M����'@�SI\B�ɢ1���@��S0Wԁ�wjߤ^�"B�I�n�02D�;uurȣ��B�I�T2�"�c�'��cRʕ�V�2B�I�Y氬�G�V*p�:$`b@�M�$B�	3Z��LcED��ʈؕ�/^$B�	=|�0�õ�T>� �Q �dC䉾Ll�`C�i�����Lu�D�d5�S�O��yp�dL�4����b��\�h0�"Oĭ���/�T��F�`q���"O�2p-Y?I%J�s��`b�u�s"O�u���&9�DJvŝ�{�t��"O�Т��B^��"���S�l�S�"O�($�IE���s�Y�5/�S�"O� ,�"M��/�P�ՍJXur 6"O��f@��<�x���Zf c�"O$�����h�"�*�kڲ#�N�
�"O�|��h�$e���#�i��8ǚ �#"OfÆ
� ���@�Ӌ6����"O~�J�ʁ�t�=�a�  �XH�"O�p(���rG��X���:��\�"O��:��^�P�z@��X r���2�	t�\[�FH�g�<SQ!�?Z��K`)9D���0)������e�ǣ,yzqZbk5D���BԵ_1Z؀V��+c���A�2D�����eMVzG � �Vx��F0D�̋�̗\���5��:��4�Ѫ,D�$��݁TN�p�J��wn/D�Ԙ �}`mɀ&U���<Y%C.D���GM�!j�Bè�U�Jpq B9D��
s�� ������> 6����8D�T�4��9Hu��k��L�.LsE%<D��aġ�\ @Q3�Yt�	�'�7D�x��Bّ@Ǭ����O��|��3�7D�HZDO�/��Ԁd␎<�T�j6D�|�Sf�ty��gC������bo.4�0�Ϟ
yg�@���Y�f��r&�U�<qc�߾?|�p[3/* 쬠U��E�<M�}�� �ŀ^����F@�<�%���P�ie%G9.W`�%�}�<S��r����V��CE�c�j_d�<�Q΋4gk�Y���ˑa�l���.�b�<!���5)8�	CuEz,���6�Z�<�����p�i���
]p �r�B�l�<Q��T� b]�V�	?KnEHC�k�<i֌�=x� `w&��|�hJQ��h�<!#�JD�z��dϸ2�^����N�<ၮ��'�N��ھK���AM�N�<4���9��HD��W��_�<i�&C�{x�X��`Y�~�ճ�[�<!�C�6�^|Kg�M�0Ǯ�6G�K�<A.�(`
����R�AY�,r`��D�<�ER��8�����	���XY�<�'�O�+̂���\�R� �PS�<��e�,���h�9V�����O�<1�l�x�P�@�4O" �d�I�<�E�%��\�/�-lb<KETz�<�4GZ7+�j�Y�i�&rܒ���Z�<���Ҟ9�H����d�r}J��k�<YR�`�� P3(�E[�xzj�a�<��	жZ�8����̟�4����D�<�w�!?[�U*g��pv��) �~�<�b��6��`��_�U�>i����v�<Q��='B��aԫe.4�Xs��p�<Iր	��ȨbT
�y&X!@�ITm�<I��X ��׊�� >�x@ހ�y�	9�(I���O�wb�uk���yR$@7"������Z�~\�8�M��y".B/�bPb�$ğf��	(�y�ꍓX�̱)c	�[���T*�y2�kr�����X�j�c&��yb  �F0F���mM�IA� p��Ha�<�b��V	ˢd� {�T��%$Gt�<��*t��i�� P�M!S��m�<�!ոg�YYq�A+R`x�HC�<I��"Y-vax�T�w�����v�<y2��q�,B�B6[�����+t�<I'�E�x����h��=-�`+6D�� ��k�g,n���v�R�(`"O�Q�e��?$ʼ9Q#ҞTzn52%"O}k��|�>��LI)a^�`@"OtA��ӡx���
3u�J;�O#D�|`5��x}aW��Mw�d�F D�0����"3�69�Aa�4}ȸ9�,"D�4c�I�%��� FU����c?D�<�b��Y1~�v�4P:��b�@?D�D:�M�6-��qmM�u^��7N:D�t�,ʑQ����v(˾VR�/�y�"vɪ�S ��#�a
 ����yҦ�������/ń�X��B�yr�Q�׾�����)���&Č�y����Mh!#!��q������4��d(�O2����>6��}#��9�pa"O��yD� 7y&&���B�p���"Oư����|p�{6������"O%91�_;�x�'��=#f���"O"�r᫓z�މxs&�|�ȕ"O��aw��dD�R@�@�x�ʧ"O��#��[�ht��S%���[D�|�'�QA���:9/@@B��%Y�!	�'��I0���J�ܵ�ѬX�PU޴�'(��7��0-���MZ�r-h�9�'�i"c%�~� �AՋշ�=��'z0�V��E1�Bt���BH���y���.�viJt���}"�`� �yRE�b�zAk0m٘�,��JD*�y2��2� uӁ �\#@�b��W�y2��O#��A���&H��I�&S��yb�ѝbj��� �ȵ|ډ#�S��y[&_z<#�+\1д�`&"��ybO� |�$ Iqi��ٲ� �9�y�u;�R���1~l�Y�u���yb�!ʠp�r�n�`q ��M���$&�O�^	JVY�r,�!y���'@�{�<�4��ZlY`l��30��r�g@u�<1�C m`\��E���Ȋ��y�<�R�L�}ͤ�r	](p��qJ��
`�<�3��=:�Y�b��&yh.ĢB_\�<Yc���Y0�ؗݛb0HR�`JB�<) ��T�PK�	ѓy��,��E�<!��H�O�4Y�F�y�X��@d�x�<��k4�Y���χD�����|�<�5a�8�R���yd�-�獜B�<y���5H�]SwEޕ6?B��.A�<i �U}�����N%-,a ˙f�<�p��I��@t ��A��Jh<�2L_8�� �і�
�����y�薌"f���1n���V���ˇ��yц$�b$!���{m�0�倆�y��E"U�b��R�	�d��|�a�(�yBG��9���t�Ʊ0��)ժ��y�ȣ1�4H:W%�^R�aYA���yREӦR�j!SC([l����L��y��j� ���h&P�^!��@��y��@�<Q��*]3F����"ǚ��y�,[�+�V�X�]7�R�#�Eۛ�yB'&����@i�+P�10�V��y�َ���Z��W6�!�W0�yR☢-)��
$b�/>���/��y��xn�s�/�:!�,��FS#�y�	bD�c@ɹ	�npa
0�y��o�lh!�u9�IB M[�y
� �P�4Cp�ɉ���2R�qZU"O� ���	�2lbn��Q) -x�"O�`	�O�L�8��GU�%"O�Q��/հ%��čH"A��y�"O�1�w
�B)n%Is�C2q�8Љ4"OQ�p�$a���c�]0�&hIp"O�h�c@ْnJ2�a�^�D�Re"OT���ҁ.�R�[��*{�t"O@�JBʀ".����OD�[��a1!"ONEƏ,br]y��\G�\��e"O ���+q�a�o�F�ʓ;D�� ��
I�t��P/ݍB����A
9D�,�C��@%P�Z�۸ax��p�:D��!+RU� �����
��H9D�����|�� ���*�* +�f8D��Q�F%`b@Q��H�PiHL��'$D�8� ��+}�1P��E�|����� D�| sV*J� 4�R��y�PR��*D�t�r(�){d@��8O9l�B�=D� � J�
�:X�� �))�X0jQ�=D��	�E�q��(��i:;*�FH7D�$�B�ʵ;����D�����7D��Q�l �T�ŐY4��a3D��x`�́6�:���� �c�X�!�O>D��@C�Śk=(=[gM˶P,�S�?D���d��9i�N�j0lH��l�3D����(�A%�DxTlD+AQ�|�C�1D������<���A(`�l��� /D����hJVl��柖]ܚ4�+D����o�0O���	r�]%@@�<�e�)D�h�B��VdV���	�mxؠQ�:D���ˎ�X�tt2��5F�H��#D�!�OP�f���Dr�,8�&>D�h/�+|�2�0f�A)���p�"<D��cH>Y��)X1J��as�8D��r!+�\h����>���i;D��Z�-0g$��*�$I|��A�9D�� ��H5����*�� pfe,D�l���Ɓ'�R�eZ$$�|��"�4D��h
��������?_d쐆�3D�T�-מC�v]�GT��L �=D���3cT,Ok��p���k}T,"��-D�(
�h��H�V����P�jqT����,D��
��^�u�xc'� Y�,P�V-D��{b�B�;?���#/pް	 ��6D�, ��I��)���"D���3D��h1�\�.�*�[V늣2�d�`0D�h�Wdƞe�h�2�bjt(�/D�ȑVe	c�r�l�*����-D��'�$�����"I�s�}� G-D���o��H�����
C -D����H\�l�P��#l�!N��09�@+D�,����U"�� �#{��j��(D�0�`�=����$%Q�\���&D���w#�5l�����N0l���q�i"D��(A/��yP	��@:n��JW�:D�����Ra��}ɶ�@�^���F9D���a,Ӑ*]�p�[�gtj�;`�9D�|���,J��T��(j%��8D�@�� 0A\x��L�)�YQL9D����X&{_��	W��e�8U
PI9D��3L>O?@أ@V>
"X��a7D����)��3� �G��2��<:��)D����iB�F]h��@���J��vC)D��  I�qNG�S�#�� 0+��"O9�F.�,�aAU��Y�"O8�{��YY�ބ�ǭ��u��"O8!��f��#Yb��s놐c���[e"O���I&)�
��ԩ��5Ѯd:q"O<���EƇ�Q�Ti��5�R���"Of�Jum	�*�|S	��@Ÿ���"O���f/�$\��@昀?҄`�"OR�� \٘�:�$��64!�"O�!!���6�=��ЃQ���ۥ"O��wgƠ? 
���Hӫ=�<u	 "Ox����WP
���sܴP"O�<CG��X�w�ŸSl�R%"O�8���шZ���s5$ON����"O���VJ٨k���/��xѼ���"O*��J)b}��bRo��U��x��"O��C�+����q쑆Y;l�%"O%�L�1p30Q�d�]�;(��a"O��ڠ�
U� �8�ʃ�q�&)�Q"O�G��.�x�q��>4�ye"O.x�b�}����H��yR���"O��J@�&2�NT�F�G�<{�"O�}Iq��,���c�:V>Z�"O��!��0��`K�A��SW�U"O@�[�`ƨf�L�����YNt耇"O�`r Ń7�\��+݁YK8){2"O,��V�ߑ;�Ĳd̒�I��1��"O��Y���.ɞt�vj�1#���*"O�Q�Gf�v���O��c���"O� *a�3m������(_V �"Ol\X�g��a&"��G��Q�����"O0��`�8CwDp`����T�NX�<�3o��)C��z���#d���aA�O�<!D�(R�B!�g��dP���J�<	����j�������/���j F�<QAMQ�<�kf9V����!�f�<�5FU	MӐ���		Vձ1Md�<AUń�t]~$1%i�T*$���Wf�<a1�(��H�̑b��XC�_F�<9��W
&��Qᴭ�\�>����CH�<a�gʕ��!��%�8�8�D�o�<�����H�E I�>�a��Xo�<чA�i�ƔYƭU�v���_�<!׏��\sb P�MK�:�3#[Y�<!gcܩ�N5I�呲�ś"-W�<���Z�"2��H�T��c�/P]�<y� �k&�̓!��q���Ba�S�<Ap�����{E����
���M�<iE��g�H9c�`B�+!��t�T�<�3G�LWF�����V����UP�<q�
H�F ��#���h�@8�4�VQ�<i@��d�hE��=+�j��i%D���&Μ1Ԑ�� �>]���q�?D�H`�K/z㾹��!^G�r��?D�$3&��(s����B7j?b���=D���'���"�V%
�l_�Q���)��9D�Tؤ���B��Qr���&C�����5D�0*0�� 3֪E���Z��H�D�3D� �1�܀rɦ����_�b7���&�=D�&��

� !�I%h�����/D��a�,Cآ%���
�N��q!D�<��޴:TFd��Q.6}n��ł4D�p:F�-1��Y��dΔ\< �6T���6
�(U�(5*�]�GL�1"O� ��;��B�:AS���2�±"O<���7�z�R�N�0ȼ�:�"Oh�Hf�ƑQ��Y�c5��"O��`ؖ_BPc6m��E.�,��"O� :���
3AY�Lˎa�p�"O�=
4�!m�H)��77Ｔ($"OJp�dK�*j���x�g+*��	J�"O��IV!A�Ήb��ML�m��"OR����W�h-���X S-<�Q�"O��d�Ռa�hܲ�a�'G�A�Q"OV�0��U�0P�f@O�4 ��"Oj}�P��jB��ۥ� x\� C"O����4�vѳ�oR��5��"Olu@����r��h�	 ����"OVa�_j`ppQmT�~��c"O��&a���er��; ����`"O��Qa)��!f�I(׭�AД��"O^�zҌ�*�ީH��5�z`�"O��ʐ�}6�#�@�p�^��f"O�`��W�j��5����溁˂"O�lA+}�b%ɵΏUCVYAF"O�Uw�R��	�E�K�S��� 1"Ol�hD(��6}
-���r��C"O�h3�c��.�,{�K�`�	�"O$d�!�1.n�i�0�N��Ĉt"O��c����-blW�<��Ƞ�"Oc���',�Y��W
nL��
7"O@9���#��{��A a/0�
�"Ofy������j�NH�f�`��"O��ꇄȮMu��+�CM�#��ye"Oȱ@�aÚ��h�-��Q�B="O���k��f��{�A�L�½cG"Of�┣\�1K���pa+ pAX�"O�A-�ARl4�A�	t��%"OJ��r&�2l�$�#���j��"O���M��R`@�D��u<�L��"O��1t���>��(��)�d�:�e"OZyi�ϋ�����a�"�zd"O� �[T�D�r������P"OZ�:�����U��(Ixñ�"O�L`��:x.y���ƴ'uB�r"O���.+d�8؈����@@d�4"O�����
D�ȳiԎ.@��"OL��aNϹ�����-�6i7����"O��ϔ){)��SDlD�ZJ  �C"O���E�a� XT���V���[�"O�h��N@�`𜓐J��9��H"OD[���0A\�+R �2��hp�"OXt��KK�\"��RnҏgY���"OE9�#S���y�bl�^C�ī�"O����J�k>x"�
D�R~��""O֝sL��^ؤ�a�fE2d	�V"O��,\���ec.~Q�Q�K
�T�!�ݑ2C�0K�!�a�ƜR戆.[�!�$?$/\�J�׷�n�T����!�D�he�ܳ�˄)>�P�TfI�,!�䞄S��H���Q?*i�l2EoI>�!�8T'����"�R��i�v.�K!�W(<�Ph�@�Xy�l)b�E�!򄇖v#(���iȀY�R����M�!�עoXάBs*5F��E���է9i!򄔭rKp̲G�Fq�.�  XnJ!�1`b���cˍ't�]c����N4!�d��V)���T� ҂�HV�j/!�� ��������'m	>���"Oܡ´&��K��8$�02P�4"OƐ@��7Gw��)ʂ��fm�"O�f@@�]6.���ލ3��"O@�:�A��V,���!H�ܺ���"Ob�+ֈ��8!܁���5>�0 yf"O�+m��W�$���(ɒ`w��A�"O�L� ��"�v��@�Я7��1�F"OJ@���Tg��c 0gM"Ojë�� c`(��
[�L�*u��"O���E���D��!+��V��[�"O2�Xg#!��l2�"�5>_V�"O��FK� �i:c�N�`Y�}��"Oj�E�:!�DX'���W����"O����eҦW��{��5?���"OP�#��L�m�I����Y$���1"O��z �לGIBM�uo�B!�`x`"Ol���"Z}��`�nI~��A�C"O�Y8�=d�~S�CO?k���s"O�$��M�Zṟ��"�~טp(�"O�p)W�сnW8P���Cdn�Ö"OX@��԰ײXX��X����"O^@G�H>���ږ��G�2A�"O�q�jZ�`��-�P+�6rDM�Q"O��A�/��/s ���T�SQ99T"O�0����+x�c���K��B�"O���)�g�1+`�|z�"O��@_*<U���)K��+��$D��;��S�R�И
2�+d�@��M/D��`C�N����u�(_��)1�h,D�����]%^?�bG
�Y�$�2�/D�ı$P�L;pH#n��\�^`Y�+D�$yU�)o�4�"n��D�G/D�@zvh�`� �`V&�)A(���/D�p�F�<*��b����O"�%�G�8D��˅�$��95K�3!*�a�u/6D�������s�j)B�h��(��3D����Kךja���4�C�<P��"1D���qƟ��,�a_���t�0D�Јsd��
����ߐ$���7�+D���׫ʷ@��#Ԟ��'&D��ɐi]\$��ԡ,�~����0D�(Ё���<�����R�f`�b�.D�\@��J�<�h�[c�"y8t:��,D���`E�;7e�����;c�l�n*D�hB�eq�(�ɑv������&D���¢�H�$���-W��$���$D���� [�Ƞ[��O R����'#D�`C�:clh�R��s���e6D�ġ��2�>(�`L2��c�l5D���b�0T�)���*Ѕ��'D���So^����r`OƗj� 	A#�#D�0!��	6��Ȳ���, �c%�>D��jR��3(V ���bYN��PPr`*D��rweJ	z�B� �ɉh�����*D�����^�r$�1��6��pI7*OF\)�oԀBz�'�بW��"O<0	 !U���*���uv~}�G"O�$�'G(%G~�a��X�|a҄�"O���G�x ��pgP~��$"O<�򵌜�]-j�À#��@��Q�"OZ��ag���8���rP�:�"O�3g�;R<�"sЙ8���""O�	��FN������\5����"O� ��
�'��8�*�i��+"On�h#(#h���b�į\�b�A"O@<86.� �����C�Y�q��"O��K�I	�^��(�VE�G,N��"O��T畽I���C��:̝�"O���4�I�u���@����ޥ��"Oة�5�\�z�������[� !��"O�Tg_��h��1�`�Pz5"O�,���Ǽ�%h˿K�	3"OQZs�5~�4PP�ϲ�8Đ%"O���M�68�R
��Kj�(s"ORD��BξdjH�*W�Z
uM���"Od���MP�y�'QI�l̡�"Of��4�����('���l8"Oh ���>c:!+C� ���'HDI2�dʿKv��#����<���' ��I3'K�@$�� �_��
�'2� ;��3MU��ceC�^�h
�'x�x�5 Y����ԃ|�p�	�'��aģ� q�3���a��*	�'��<�`�K�9ހ�Cd̠]�q	�'�J=�ҫ (�U�#�ʯ 7�e�'It����o��U�硃�f<��'Ď��AF/��HwO�)_��ܠ�';hP#c�<:a��)7��?R]���
�'�xm�&�/7�0��C�4���	�'lc���o*5k�j�2-�`QS�' �`��,��ٹb��'���'դ͈t
��XZUp�X8i�n��'�̬�t��.g�ʩ�QoG&^�б)�'�B� :7��qa�ͨ\v��'T�bm̑iAJ�Ȁ�PB���'W*c���'D���I,� ��'-����M/ljp�I?	�:$i	�'�.0�S�S<r�̙�kt+b�`	�'�N�3`�ؤA���D#��4�*h��'�T�ZQ�Eu�<%��iR�,.�A��'!@e��֋X/
�)��H[�h��'���æG�8�-�R	�N[�\@
�'٦ؓ�Ɂ�$���r-��VτE�	�'V��(3�ٯ{�J�%�аTF��'��-��=>�Pc#F&7�j��'B,�6'�.pxi��(p�'�L$��
h���㌋'�p k�'�p��:0��`�@_�!�Z�[�'�hr��I���b�.~���'�4����٪&�8��\�x�]A	�'_P�-U��V�O4�Y Ek�(B�ɞ4dp\y�
A�<��Q+p*V�t��C䉖%p� ����*�H�-P��C�Iu�uK�GŅg�(Y��	�5?NB�	- @Wĝ�XdQq
<�,�	�'٬��e��1��}2��:u縅	�'������RxL��w�ܭh`BQP�'�^	sDk� $��͛+g���a�'�p���\�4Z�З�o��ٰ�'��qB�
�+��% g��n.�I)�'��YA��
?�����(0�"@�
�'мi`b��{>���c���!�v�;
�'���щ�8��HKд�/;x���'ˮp���F/���7�	2+�$5[�'�v�t�C#�fQB'��9nY,��'9��m�d
f� G�9i{ƁK�'$�����,kvt�Cq�Ϯ`�hI
��� �!���E>���c��*�� p"O���P��xa�7�j��"O�zgAArr}�u Գsc����"Ou� ��^u���)D�$h#"O.����ǫ��:⍒#;���"O��䋕�8���+�f�m�L\A�"O|�`��]���eRW����p��"O�Հ	YB�&iK�h�4A���0"O���`#�&H�9c&ӺG�@�"O�l;��^|#t�A����\���
f"O���#�'ONlu")�N��6e/D���GïZ9��ؠ�?d��C�e.D�°��*	����Q�A�-Q>�!�`8D���C��$;$�`P�I-'��y�G;D�p��Y�>8�4�@����)sC8D� ��
�m������4ԝa�8D���*�%-��#����g�Ν��6D�X�C�B�{E.J@�V/M��cC�6D��/
�U���A��5`�*i	��*D�h(2�Sq>l��̋�Cb��9'�&D�@��oK��x��F� U���a��#D��ӡ	J)��<[e���q���3%�#D����֮\Y�T(݈_��A'� D�{\I�2(4M�;�ĠS0�?D��9¬>�0˗(S���;D���m�$'��eѳ��$�ؼie�7D� �d)��$�P�R&�.'���@�4D�\Bs��p -��Kz ��6�?D��:�ˍ\p+��QM֍���!D��rf���
r�-0Ä�>��QC.$D�4pA�C��MXpa+q7޹J@	.D�T9�['ڬY� %�:u�e;gH&D�$R'A�F���XQ-s ��K1D���O�;�$H��j	�bO�-�3�*D��z6�A$.bHK��u���&D�0��OیF�l�q& ,b*�[��7D�P�J�`�ej�F*lJ�E;��5D��p��٣t�z@� l��d����6�0D����$�D����`�9#���I�o,D�|`����qn$���'j� A�<D�,���H�T��-�&Ɋ���-9D��b%�	1�h���Y�
 ��+7D�X �,���X�5�Y(i0�{0�'D�L8��D�����^���R�(D�L�Ǆ���X���=2� �2u&(D�DZ�!B�n�r ����D��2��3D������?ZB�u��H���f��46D� �@(��X�8Ir!�g�3D� �$�	g�J �X{�
jsA7D��j��@K���P�C=X5��05�*D��b�ҧ#cީ�P'��	��Jr**D�в
M��z H��V�,`��d'D�xy�HɻZJ|0h2�N��X�*!D��	t�Ȍd��(VI] ���t:D�8Ȥ@ D:y����?8��-@�3D��i�%X�X-  2��.�&�Rs�.D���V����L�y�ަa��@��� D���E�ސW������|J��"�?D�\�4�]//϶�����7\��V*O:=R =��K$0y�qw"O��-\N��1B֑Q2R���"O��q�H����xE��Å"O���!��m����6�֖Q�N�[ "O$aRE�� #wu��I�@�4�(�"O� lD���˷�M2l
�[�v��@"O�<+t� )[f:�8�G�3��@�"OH�)%̋-Y�YʷfB<���SA"Ob�J�O]�T#�03��[{�~)�v"O�����ͧ`��1�)Pu�����"O�y1A�@I�򰲧���F�z�"Oz(����P� Z*K�p�q�"OdA�g�6ya�@�����0Ģb"O!�7	�;:/ր�5�O���g"O��v��E�"�*�LħkE8pd"O���E�J�fy�()���#y9�"�"O|�B %�Iw�eLD�z��"Oژxb�:p�L:�j��+\��"O��Ye΁)gخxzv��;3�t�"O�t1�mU�#\�9%�c!����"O*���A"x����u!��̩�"OL�{�膟+ ���O�(M�恫�"OĈJ ���-(`̛�F���"Oj�U�U�S�p��A�8$���"O�	��ME�
Dd)s�b؁3��"O����C�B��Y0�B@�գ�"O��El�i�z��Q朎F�n4��"O���Z�(]Z)�4E�)����"O���J�2^��!�IӘ7��)�"OH�ᑁFH��2E�D����G"Od�B�j�!mXi��k��:b�!��"O�T�0�ʁ_�<�i�*�RI�\�U"O&q	RkTC��@���/%��"O�Ay'(8,���_n\��"O|�ďK�(��g �q����"Ol	8 �P3P���I��i�� B"O��I��/a��IR�I],D����"Oq;G�1:e�����> �t"O�"�	O��D����Z떙�E"O2��_̒�)gw�y۶�U>�y�� /P��2MB*X�d�PQMў�y���3b�%s��]'[�d{��y2�L�D|���!��I*v�む)�y�e��PP%�%m���s�4�y⩂;��M#A��2(Xf����y�̐�/ΰ�"�+�Xc�!����y��	Q�ݡd�̏K�֡"���y�E��S1���G*:��q����y�ς
���㍍.M:U1�L(�yB�O�� 4P�G�Ux�Pp�����y�JA�Z:ݱ�"ԗJo>�*F��y��Q>g8mp��I@�)�E��ym<��1��O�,`��Ĉ��y�Y�,L#G!m��x�F���y��H6r!������D��@'� �yRJZ$~��9˕���6�����	�y2D��+Ѽ�A�Ƒ�{��u�b���y2�ה�1r�Fix<�����y��ޛC���V� \�|iqvFK��y�ݥ�X8�&'!:i�y2d@��f�[�n�91֬��	��y瀗�  �P�HZ"h��Rl���yrڍ`��}���Y�(#�B#_�y2/�5~Jq�C�RX�ܐ��լ�y��HR�|�S� <Y>|\��(���y"#�+HLE�j�=|<����V2�yڵw�Y�oCw������σ�y�	0T�����m���CE�Ω�Py��^�4Y�'-��[���s��Q�<� $-�eƔ9a�9S�φE����"O0��ìի �x{�d�22y��"O��� ڝc������T����P"O8�`�>#A� �� s�4��"Op|afo
�*0N��k�8,�`��"O���ʙ��Z�4|ym��"Oz��E����>	�V.N�,�qs"ON;'	Т�A�E��l�J]80"OLXѡ ,|/�%fX ۄ��"OJ��v�Z#k���BE[+c�D1"Oa�eV�vDA����.idk�"O�\���	�<�f�P*� m@M �"Ox)����K�f|a��������"O���&�*�ک:�nҪ;R�U�e"O�@A��ˌ7iBT8 ��@+P���"O�LB��D̉V�F(Jn	�"OX`��ӕM�
L��\��"O�5��@ӰZҊ�â�>3E����"O�yDV�YԮ%X�#�\D��k�"Oh�`�J9D�[�BAR�yp"OQ���	13T��a�OE���"OP�yՇ�x���D�Ni7����"Orц�P�\| B�ݩgӢ��"O��NN�`�x0�1��r���1�"O�@d���DJ&)�q��D����"O���S���ɂ����(���"OM��A�I� �S�<��m	P"O� Ƞa�:,�9��[�=g�}C�"O�a��Ί5*nAA��ΑG��P�"Ot�Ja��7�j��B��!s"O���r�H�N�΍;� @:���q"Oz��1�HL�+�`��k�@��"Of0p1�5-�^Hӕ�R�8�*��e"O����m�^N���3�\�8�B�{�"O��h��9��8XR��-�~��"O��C�k��~pRqnK�L�P9��"O2��g;t�9�kK�v�I�v"O�4���%XNh0�EL�$cN��"O�`W3��Q2^���yy!�dA��nY��bܩQiʭpWiM�xo!���7̀)XB�QBh޼�g'N"e!�$S�w�9��h� UU6X �&�v�!��#GGXy�@�0�x�	�ڀ3�!�dI7Z�QA�nC�_2�CFd]��!�հ=*�Scd�2#�䋐(Y�!�#3+d��@���z!�LIŇ�3tx!��̈́&d9���G"U�b)˵D��6Y!�G!j)V�B�@�Z����l�06X!�@�}��MX0Eٛl�$2���R!�$�1M���!�� e�� a��z�!�$�K�R=�%�4?��"�/Q�^�!��8Z���q$ś]m��S�NM�!�er�Sb��mM<�8գJ<�!�D�\j�}J� �,W�)���R	!�dC7#<d� iT;��I�ɞ�[!�$ی]O������$=��iԈV�4�!�d�(��b�.O\�y�F�_�!�!��-(ň��F�TV��a#IX:�!��P�]
�J���r��!��^D!��,e�X��l�ܱ����f�!����8�Qҁ��D�٤�#�!�G�[.2̐p�۳�:<*a#Z!��7*�\C��M:7L�G�!�Ã/��eWj��j�<e��d��8�!�� ��AcJ ;v�[a�� BJ@\# "O��Y ���I�����善%<�)1"O.V�)L��bTmP�]��lScmV\�<�"�P,b����h�H����Qf�A�<i6k1LD4�pNH
�JPP��H�<����*FP8F�j2����JL�<A�4�����¾S-b�S��E�<���>'��ۆF�%S��#��@�<aW��A-@|`���,����}�<�G�߷M�<��l��o��20�|�<�G��g<t��a\�1�x(�COw�<I��e|�r�֡�΄[�@u�<��Y,3(�7�NE9�-�2f�g����'vֽ�d���f�.�Bt�u���'^�	�׍�Yz�`tM��r�¥c�'���ƏY�A���i�$v�$8{�'��8��\M(S⒅C�D1�O��=E�dm¼0צ��5Gj�	���1�y��@<T�4���.�E��l8dGA�y��Y�V� I�h���ps����yr��J-0g/�o+0U�U���y�GZBHH��c���$�M��y�B���x֣�,S��QNՊ�y�3E���ԝ%x��򰉚0�~R�)�'⺭���RT~�xT�ǷFU�5�ēM��6�+]�x�*�K�!VW�(�M0D��j��pQ⥱�A�	���`g1D��VM��:*�YL�{�z���m+D�h���,p�z&���_��#*D��A�e��k�j5��E�H_ �Ia�;D����e�F0�5'A:>��	��b��(�O��DâT�R����N�أ'%U�3�|��x�e�2͚u����"���0.X��ybf�$�Sc���h�B5E
��'!�'þ"|%	V���LJ�r;�`G��a��&�O� �m
�z"�h ��3WP���>)ٴ[��d/}2��Ƙx@$�`O]%cB�\��d��m��D�* N�!�ĉ��!@�����ً�'��	�,�)�L>ysb&C.�0��O=W�"��j�e�'{����; ����� Q�J��ҁC.Xu�B��!+Zy� +μ	_V�+@�-Ӿ��dQ����(?1s�T;U\Q��ݰ|m�0V�	W�<1uA~�VDs"M'[�|uIT�D{�<���O�.l08�-Gw'P�#U�y�<9Q$T��F���P� c��˱J̟�'��V�^@}J~&���A]����EN���xs�'$|O�c�p:f�ϰ�C5��G�\L��j#D���槞�Y%n��5��1[ T��"}��O�6-�<�p�r>��?	�ՀQ, �]!S	�	 bN��o D�HZ�i�L�%�%`��-�d�<��hO哦<���C@�έ=J
�"�X��C�I�K`:s���\y��ɇ���bX�"�%�S��?VᚌA>�uKsA�v5l�3�D�<Y6d�%d&��=&���ůQt�<��m�Hw�T��Ô�F�3��s��hOd�T���T	D�~�±�+h�8p�G"D��H��p���7%��+q�?���<���8k�����+"p�h���}�<����>P��q@
c�o^y�<�AC!4d��b		�V�sL�v8��EzRHBA��xyF[4 aRT���y�,� ]�I�e�"|�A�\��y��É<"V�(��C&�I+V	��E��5�O��H10�
t�b%P7�as2�'���� (�� �Oo��q���%x��XE"O`L�r��4?w6`�
退BQ�@D{��iF/�����_�J��MH#%�!�Ĝ�t���#&e13=Ƽ�eN��J2!򤙗s���!�C~/�����4:!�}nz��t��)!����l_�0'�*�O�(ؓ�U(�x��T�=a��"O�<�0�˫B����a�`f�"Op���`����x�P$��3O�=E����!1��X"hF%3�4��+��y��	j"�t���'z����Q�C,�y��)Q	��(N>u��ŲmhK����ا�O1z�ѕ�C9���37!-	���
�O����@��ځ���!t����%�����y���0��D�yI!,N���$*nC��a��O����[�%��d��
�o�N�
b;O�b�,ק����/hJ,}#Q��N�J,�lùu�!�DŶp���A�-1!��Pe
���	Ix����,��uX`I��F�>]�aH�O8D�xr�Ҫ�H��뛏vR��A�#D��0��[;}~��f�u���k�!�OXO~����>er���?W�]��"Oz�#c�����Xr�T�Da��<O�ʓ��S�$�|�$^��zd���ŘO�Y8�G�(�yR�� ?�*���aį{Tꐱ� \���'��Z�S�'OuBU	PN� q��o�
 ��yGz��7��;��
��6�*P�d)�����d쓬y���O��k�"l֬�4K8A&0�h��'��#=E��U|h�K2��+$�D�8e�� �!�׵2f=�dƙMv��Q��(�铅�=�ݴM΁�Q�V�Z�;�*!fX(���	dy�Ϛ :��af�E�Bga!�@���O"~j�iDB��b� '��,x��Uܓ�hO��ǟA�ā�rO�� Y ^��S�>?Y���&�"�Ŋ��]�2���U�	���Fy�)�g}RƊ$v��h:M	6i� �je�F+l)�'�a|�M�+�nm�!�<"4쐸%HQ%b����ԣ=��BH��<�p��V}��§�k�<IV(�}��W��U�j�2p�<u��'e��4qWj��G��_,���#i����h�|�� �r�XZ��L5�� �I�<y	�F�.#�\�q���ɃnT�\� Y��	G�\��˄(��i�&ӱ^� C��86���W�`R�"�+`#�C䉘[x&d�u�S/d��#���ǺC�	P  ��#薞.�)�P"�"�C��n��d:4,��J�)9i�%)�C�t�
�ۓ6ǼA��C�/E���N�Mݤ`�i]�rFl����3����c'��F�#p��熉${2!���TU�����_咹jE�� W�az2���j���!�/W��1���58�!�d�7��!)��K���ʱm�>~�!��0b��D��I���x���B�J�!�$� �%G��w�YP��+w+$]��'_D8����C:B���>qQ���
��~LO�!L,��E�:���O��yr�Ų���[�g��{�X�b�oS*�y��X����Vz�R��V��4@�')�T!%*"a[��z@�P5r�1���' �9㫚�r;�0��,��Vdr�'�j�@ΘcLd-!��D*4Hqh�'ipD2���u�D�R(��8�Uk���huR@�6��g��x8�&�}��S�? �) �m72��i�BT�wX4�"O�ڥb�'	��F"�R�];�"O�u�R�v�z]� �<�$�� "O�D�f��r>dB���h�����"O��6��n�hz��1b@dr�"O��儇1$�&�I /S[��8$"O���#�F�P#�QkWT�HP�K�"Oz؂E��SD���4�	��U(�"O��;@�l�@慖�x��"O�����-1ҍK#�V��q�3"O�m�4-��\�
#��
,riu"O�E���0�2��2��%H�}"O�K �Шql�+�(�;XV^(P"O�-�#�ju<�'��&�p|��"O�X�D���L��d�Z�r�n�!q"O�
R��/{�f��e�YEp"O~d)�H�3���XdJրj?`��"Oj�Z��K_\}��)ۣQ:�C "O��Q����cA$��c��a�"O���
Pv���b����(�ą"�"O���P�\Y3�[x����"O�	�"��}�G�M#i�!8r"O��r�E�&�d:&��Eص`t"O\���J�s{��r͜q���J�"O���̖&|^�q!&��E\� p�"OL�ð-4gXh����2oѢ�"OnH#�E��F�ऑ��)"i�\��"O$�ң��$2�1��A�:>���"O���ǂ֔P��Do������"O�mJ��84Q^�t��o�u�g"O�0�DJ�5.�	�6OY��"OZ�(f@.L�J2A͔{:���!"O^���ȇ3{+��b`ϼ�dJ�"O��j�I����i�L�m}��B"O*�0.Q�|���#a��D,�y	�0{j��I���+6����X��y�W/��}`��6���;�k[��y��%M!:��O� {�D�$Jٗ�y� ���Ы� �oWXl��HC��yR柽gq�$k���z��tJ�L�3�yr͒#ШAW(ϒyh��Ro��y��e�L��r�I�
X�R�O��yrd_C�쬘T�ͣ@�z��c�
�y�a��~T�J�CAL-Ҩ�ǉ#�y"�4_瞸�V��40���H���yR�Տz�p��qtl]8�C��y�蛜@���5,ϼe*9�'C!�ybK�@@���#�[/]���&�]��yB$L+:�~���ߗY�J�#@�����O�����sQ���k�*V�2OB�	F��&f���O(W���t"O݂��@	9
"x��im���"Om���(K�:|�ℽ�P"O�|Z�/�)c�F�1� �N�0��"O8���̕�b�K i=:P��"O��Г!�B�\���LW􄓐"O6xQE���9�g�On>�g"O�j��F�Ju|<�&Y�qoD�V"O.�I��	s����b%X�y[���4"O0tX�iV���WEPr��"Oҽ[g�ϓ{��Q1�`Z��@�"O\@��H N�=Ä,L�VY$�u"O.TBϱ�$��������""Oޘ�e-8/-@�I�e�	{�.=�v"OR�(B��j��	&BP�"O� N�2�ȸ3R�@`�2f��PC"O�+�Ơ
)�0K�F�;}��堶"Oꩣ�H9�B<@"eͷz.�(�"OJ�P𡇂n͸��2�+2�� �g"O�8�C��A�޸�1���"�fyʇ"O�$1���.f�Q㏺C���z7"OR��F씤�核�E\>%�Q��"O�ڐHY2�� �cߋ�����"O��z��z���`� U�l�R"O�Ѡ�m�U���Oq�}��"O��`�I>Lpcr�Rgn��`f"O6畷2,�hC&�f�H�cL$D�L+ë�i.�49�꒵A�N�Xs�/D�d�"�I6�!&��\B�E*D�d��J3e�\���?���ÒK(D�hQb*��Tͨ�	�
ߴII|��&D�����%WB����z���'D��@�ϑ�Y&t�F	�=\�!"�8D������{�X`Ei�^����r�4D���*I�v��5`��Q1h^��Is<D�̻�K�96�*X(P$��8��Ѕ�'D�4('��fu�l���'�u*�J.D�x��E�,���R�E�Y*h�X�B3D��+cb�,*Ĵ���6 <{c-0D���BOc�a�r(��q]���4(/D���q��lɸ�{F�?�pq�A�#D�<�Fc��+�R���V��6tB��<D�L3^�ڭˁϞ��HrEo�^�!�����;+X)g͌� �/k�ar͞)x����^(Z�^����
=p��|��[^h<�eȏ�>`H8I�DU�2�$����o�'����S&��eI���Ճ�V(�L"G�T$j [�"Od��hA0��$�E��p�'�l�1��%:��,�O?�
f�2	�:X:�m�* Z�ݩ�/2D�(����L;�sK�!��񺰋6?����I4�5!7O.�b���@
��5dX%@�X��'&�X�)01$�<  ���pZ�15+D>N�i�3�NC(<ɀN^1Gnt<Q�l(�!�A$X�'��{&(��B'���}�&�ca����ɨ:�l�kD�Mc�<!���Sʖ=�&
)};��[���<!��Y!n�H���C;}��Ʉ��)�D��@��(�@-�`�!�dš�bAȦ��/�tM�gͮI��ɩ1Y���g_��x���dSp!��O��4H�a�<�0?�`��{x<�&(C�Up~�)�Z>$�V���vhæTrz�!�>���4lM�\:��1��4��F|�S���)ˇq6�ɹ�F�~b�d��p�:=1r.��nla`�R�<��EO��(�EO�_%`=(b��<Q�d�
[���u�V!��ۖ�+�'c������78�����P�T���^��c0@Ԍw'�drh� y�%@>@7̈́�N�
9:�����3�	�YZh�9%n�$�.LA�
��V
���d�+��؊CmW*l�]c�c��3ԹsP�ˍ9�x� _�>B����w��}0�aA�;91�͇�az��dɂ(��cJ?��ɛw-�݀f�ߤ%�Z�¤��j�<�t˘ Q�U�Q"��t�C0@O̓u�0#���M���~��⇻%�1�cLT'TNK��E�<!5`�$8��#wkL��^x�d�?T~�xң/}�-���I�A!�X[T�S� ���Ҥ��C�Ʌ�&��r.�V3~l�eJ�; 0�UP,)놀I�i�H�c'@�q����ƺ{�T��lB6}�ĵ`(=LO��A�a<o�� �.]�0�M�0�@�o��a �"�p��(�c������d�^�����l��`Q��)h�1O��H1�k��I��h)R�� �a�M�ӠR ��&G�,�$�(��
��C�I�H��J3M�E���j�@��'�R �T�� 6��Th��s�c�%�'��ݢMs 8CD�@�S_4(� !�� �=󥅲spJ��E�.�zb�Y#0\^ +Wg���T�Pm��"��NLW�'�|�c��	%�b�ڦ�?wI*��W����"��\�t!a��8�R���#%?юu��.���#i�Nx�Q���Q���XsK/�)CӤ8�5H�!1%h�7R���8ӫٮ�!K���!!�r�%I��ɮrO�P�s�H�Dn!�䋅.�k���+@��-��C[��P���2�\�B�iY��
|��BQ>�&>�ݩD��й�m�+X4�z!��IeC�ɼt2h�A4.ܙZ��xq��Q���+�C֛G�̵Ʌ��uM�<(�I�j�i,O�1�O,����}��&�j�7�'i*	��ɉtY<�Q���*iv��Q��'x�cV���]���R��:R�i�' t���V6!9v��f
���.��x��O�Q�\�&�tjJ�I1�$(Ń���:yƬ�KS�- ��(S��M
>ܨ��'��T��EA$|2��%�_��ɹ'��
Tl�7���[(q�����y���'8�S���U�m��	�d��=aKGB�<!�[�>A�Zӏ��$�32�����s�O�3�,}��NS?%τ-��:<F��;���Z�Ь�EIh�p���.���dQt1�X�`���Y���9�ɂ�P��,@פ�)A�f8s#��E�"!�/�B~B�&OB�t+$v4�%�P
@�x"t��t�d.[����EH�K�p+�AT�m�F�'1:y�R��t�f�:�[�!�m��3����7}�pI�i�"���k�&֝0\�e��IǑ7�b�z�J���M���t���L�s���"�#]w�H�c �o�!�7D�|!�M(c�� rG��l|C�axޘ�g& p��1��ēB�Ոd	�ɟ5b�X(� �#x4U��	��A�ӘL�̝(4�EI�*͹�|�Q�G�J�̑b#�|�9O���G���bQ@U�_�m^B!���� ��xK1o�y�� J���'#9l��LH-tH
��Ȑ
x	��0��6�hAV�3N���Z�P!��ŗgOH}Y� Ę�X\��h@�X�}�P�����Ünܖ�x���5`��e��BǄe�(R�Z�����[�4�
TLؖ�V AU�T�^ID(����?�>���U��<��ƈw!�̲g�Ng�v#�ĢG�g�I�u'������&x�>h��	s3�٣`�D
E��0i��P�S�x�7�=dJ➈����@@�)x�*�.� z�#Y�\]��!$�=}�lǳ:��`[c���	�^,	"�LG38���]�I�xM��#<R���!aj�+��0�@�)�p<�T)�&3$�1q�iY���%-�F8�r�S��! �P�G�0M�rN�O:}�Qi]r�mͧ-�L �BS��b#P�V�N`�K�)lHh�@�&O�d��+܈5�\As��>�@i�7Q�2Bߙ~Zy{.N?�p�#���k��[�q!z`�����F�OF�̧#h.xz�M1����*V�u!|��O�ɳ�U�*�Z�P!D-�'c&�U5���h�`ID��j�m�6�2 �-�.��S��M�U�A�t��a`kQ�Uv�z��_�hbW^��it�мs
q��'�X����\'ha&Fo(i�O��Z378lS�W!l}�g�̖U)��j�gUpX�+\�|��\95��0<��*�^��k��]�3���52u�Y�I�����$Pk~���S��Nv8���[��R�aD�	&�?c�2�Gz�韆p�#)�N�'}<(KU�Ј{��h�Ɲ:T����Ox����L�v���C��"�'_��d�SP'}��V�0\+��nZMtb#����K���@�熠O>�(�|2*�PƁ�w�7C�J�HXY���@�>���1��O�@	r�"aj�҇#��"n ���'ԭo/>��R�ұ
2vQ3�FP̦���M�?X�Y��ɠO�4D��8J�,����#H�pD��
�4`�$���muY"�Ò&T��g�N�'X��f�Q�@:&�X�i �PҡG8��i��&�<(��'v\5Z�"Q�"mԈ������ԡ U�fA�C��@I��	/�(���ʝ'�4Mx��%�\a�$�fH �'Ҙ[ ��>���ȃ�D�	���£��hBܣ��?.@���-?֌c���2��$2��4l���J���z"�B6�gı_H�$R������fEru����;c����Ϋ��>!F�P)`�)��%D�/ڲ�B�~�l� \A��2,�D!��Θ)+�d�֍�W�$E���u;���) 8��#�-�y"ă�dS.���[�\p	���_J( ��C+^����.H�i��#�ӳ/��Ε�X*�ዴ�!�r1�U�N!�!��
,��a�h�4(���q�C�*�h����7X�HU��
�A6|��ҋ�
-��}Gz"n}X�5_5{G�P����Ұ=�Fo�(E����*� ��M����;Ƙ���9d����r'߇:$��� �IX��J��e���	a���D� 5
3�,�I�Gc��Q�搢�tݱӢ�71��QrV?�Yӱy�0��%h��"�	�1S�<᰿d���n����ԒT��pp�G����K��+2�<9Q���/��}�=� �h�r���?�$���d�(`�H�� "O�|�*μX��i�� j�(=�E`M�\��̓ej�L"h$���[�I>ғ\�J(R�
0#��<ZF`��I��eȭx�йP�FO�U���D[��h9W��' d�PU!�	 H��d��d\���͂4��<������������3&�y�GF@VW]�c_>-�����D0ӷ�ڄ�(?D�����=C
��Ύ,aB�,pF�qӀP���Ȁ}H��ѥ���N0j���i��-��!�,t�����*.0 (�'�N|b&b@�'����3 M/c���rm��?q�(?�X�Bf����I�r���k�OH�N?�KcI�N����d�O���׫�Eb�)�BH�y����n�e�Z4pt&X":#���$�$�I���p���bC���a~���D�3�D "�ԖYm� ��+��L���j_�g2��ȓ8o��K���S�t��FP�8�� �'�������5�v��O�>)���I%f���ʰq�z�)J D���Ee˾y
08BT �%>��5 5扥>��%�'C| �b� vO:$�1(��>��%��'��uq3A)^P��F��0�<�
�'�rP˧d��ZB�S�P+G�N�	�'��I��'�c-z��ڰ9Ud�
�'����&�&&��\�1NƏ4�X�	�'�����1A
����(�[�F̀�'��S5hI
}{,_^��s�'w����ЗE��ŁQ?�К�'l�����	4٨�"V��M۞�j�'K>�h��M�f	>�p�Q�G�A��'�j,��$F�*S�-� � H8���'���B�П6�X���A;2LN| �'66X0%��Lt�+�%�^g�<�A`�]ӌ��R�f��#�k�<��"z[>�:��D�,5��{F"[�<Q��02�Y��L�ҽ��͏x�<��i�	_֌�#!�]oިy���{�<�aN�A�ЋUnk�u�r`t�<��HꌙH1�C	0�leP4�k�<�"���8Y$��Nȇ@��*��a�<�Q���☬J�@7qO\�G^A�<��n1t�)���%%F�Xb��^P�<�7�O6�	
q��"gx�U���L�<��g�<�MI�'�[`�%��
a�<i��,Lk���䧛^����Ј�i�<���1uX1���:Ι�dkk�<Q�@/����R�=oX����TY�<�� r�:�qT'���#dTV�<��E�h�-���'�@xP�M[�<iҠF
��� ZY}��TJ�<a�!H�S�r]�g���9?�8Wb�~�<a�ɂg�J�F�i�i{f%Uc�<�M�
��h����I� 	��I^�<�E��Cj$Xq�@� �>��E�1D�{�%��7��3��.� �ġ.D��ӵ�ģB}"�9�@�:�pԊ/D�4��bק]|"�i%+E�vƴQP(!D�8*r��U�젋���3*t�Z��!D�X8v/G2$ HT�H<iX��3�<D�,� �(`��D�K&r�|}� 7D�D
���I�vU�&fgN�p��i0D��{��͝L�$�(dIK=�ư3��;D���T�N�"�uo��r���u�8D��u��#,�z�0h�4Q1z}jv�:D�`�1?A��r��ͼiမ�' ?D�db��1�^D:�$��E�peSv�<D�
ѯ�,�P��H	�\��a�'D���Tʕ� �^)!��ƿX�<i[�I0D�� �8�� S�I�؝ �m�U|��"O����&�%B����I�r;�a1�"O4�#o��#��ɁS+B�z?��[�"O�D�dϓ�nt���U 4,J5��"O8I�pi	uG���τ(-�(u2�"O��FM��4��%Z��Ĥp�"O��wA�sz�As��S�]����"O�ԩp@ͥ(����ڨV`҈҅"Ou%���C��)aU�Q[�ɋ`"O �*��tnDM��[�5��DCc"OΜ�v� %c�����K�9�$1�"Oƈ{ �ꨬ�	��K���"O�4;��Q�h�����7�|-�u"O�A:����H�p,�wHpI4"On}�X�S��x:d� epѹ�"OhH�4&�$��h�%ꛀc��5�"O�U��c���ƉBi�hd1W"O�@S����G���)4@.L)�"OF�Z�,Z	�ā�ۡ6V��"O2p�@̗�}�,���b�<X�ڠ"Ox��D��)�@��`�T(l�T"O�`pv��.�`��&� z�"OV��"�]{b.�H���"��AQ6"ON��U��.au6M��+�8l�2�C"Ot�p�2�����@�8~	H5Z�"O"!p��$~"ʔ;E�צ&��3�"O�5ȑ�F�Y�$5�U�M��haa�"O\�R�f��4Hq�pCZ�u�*	R�"O Ló,��K�u��=)���"Ol����!8L��3a�� �����"O�m�&h�H�8Z��ۖ��@"O����D	(
�@��.^r`�P�"O��� �I/��<b�-�^`\ �w�'��ċ���B�(�DI[��]��ؓ*`L̇ƓQZ���ԩ�1Uں5Sr��Z7��E}��M��C���@q�6�Ѷ܆y����0/N�!�DٸF����8�p���>
��D.IP,�s��/��)�'96�J��Σmrpx���S��ȓ aL+;6��=�D*[� ��'n�];��մ4)Ht��;���Ǐ_'��a1&
 Z���F�'�I �o�D�Va��AtL	ЕCح9x�X�'ۆ���#tY�4Έ�F0����$��!���$����O
u��Q�fQ��p�Ğ�`>Pb�'d��s��sL�%�Y(��'��`�_�/��P�O?u�ሐ �l�`�>[/b�*Rb*D�@{�N�/֝�aF�9�j���=?)��B�|
�#k>O ,J�� ^ܒ-i�-��8���'p̹��P�mW��3!�w5d\��������E�!:V0aG�'��i���)�B�k��۰���q����:!�N5iE�_	~�te3V�P�T��@F:���}���y��`y��P���u�-�\�Sq@�<B� ��^5*���.U�����R蘢~b�ꃣ,b0Jef\>sB�9�@iKD�<i6�
VJn��� Vx��ڗ#��cY��Q�fӢ| ��Ͻ\�z�H?㟸��`�!S�0��J�7��R��2�O�QbQKA�hNh����3n�6�J�I'"r�\�6  ����6i�|��C�ռlj� �%���1c*���0=�Q�N�K���	E����b+֞P_��GIq+�T�i&D�<;�J=w��M��F�@(t�Qdf+�7B/`�1�&
2!�Q?��MJ�3
\ʣ�G�Y���"D���q�ØJ�؍RC���}��Q!*�[*���>���z����Z 5bi)��
,=s88�ڗ5!�$�m�f	!�i�Qpa8��Z,6%�F�4���
ݴń��p�%O�C+G8O��� D�� Y3�X	��'^Zbt�F�`�lZ�}*T�ˡ�VZՋ�5M�z�2� ݦC��
� *Mk'H��T�1ҪD�&w�)����$q�5��R�w����a�� �N$>I�c��D|U�!aUM��@y��?D� �D	2B��gjT$ �8hq�FN��1�/P�}�R�� �5b�|b�O��q效~�K�)�6<�ʢ"O�"�u�E��	�>aG$T��,Ϡs�4Ia ǘ5y�|�C��C6?�뮜r�';2U��'�-��c�P��)�CIdd���O�p��� �v�P�vl̈́>N�`����[L�H��@Ux�Pa"i����8��2#�/�2��,a�ᗠj��8�Bf̓>��:��Є#td[�HY.1���J���"O�Y�vD�*����OW*^�f� V�n@PP�`��+�`���*fc�QE��w$tQ{��<��yS�o�W>����'Ӑ1�@��ג���C2J@1X��������ѭ�Ȗ><�Dᔁ��`	,ғ&y�[�+I(~6�#�BG��}��1p)d�{`P�"���B�?l���_,u/�u����k4��F�[�a}�chVq�0��W��pJ��C��'kzl��"�~�ܸҒ��)J�b}�䦇G���
�:а�%Y�S��D�5�ǎ�y���9Hj�OW��IR���:�@��D �;��@ �J�&@�3��4�'�y��[�|�'�D�@X�Y%'Η�y���B�����+��=���U�b��(
�d�S�;�Fi�'C��#=��X�H��53B�V�t���#v��r���iWH�;g�H1�r�Y�d�ҹs͋dx��G�0s���2�m\�22ش�	�l�6�HW�+af���Z.?��L�?�ŧ�Jߐu��N�+P�8��?�p�'��`c�ޛ��[0Ŏ�m#�)��=�(l2㊐�r�x!3a�Q�<���C��1� a��0L��#�鈟�䈂~Lb��Wm��o�x�x@�_CJ!�d���1cP�A����d��.>�A_2r�� �/O��ٲ�ϨOZ���iZ,e?�����iT��q�'o6A�v ��R��u��qU�SGF����i�(w��xi᪀�)Ċ�����	�٫���)	���A���,�O���BCY����.UbQ�K|*��*��j`�B�"D4�h�WF�<A�`,*����e�IQ�@ k�VB��b(L�\�	��e���8D��'�Ȍ#`�92j�ua1fR�C
ظ�'\R�z�j_�]]�����
b�eE�&��=�Q7{2٫�*A��F}B��"\j}�bBV�nD������V�jL�׉E���W�bd�W��AҜp��5\rpď��,�iGMT��y@�� E���=���)v'��# ��oV,  ��57\�J7��{��=hn���.�v(����� ؓ�&�ܼk6 �58�lP��R�O� �A[y�7H�4�C�'�Ȱ �H�1�Dģ1j�蒄C��A�U�<
3�����YѮɸ�?�p�"2�Hг!:���k�
��Q� 2�iQ�l�`����K ��q��"���0<AD+G4jU&(��N[-����#�Y�⃃�|����ģ�(T�����7�&B����\��>q���>QE;�&� �KԽ@���X�ˬX/�]�>���P�_�FےȒ��ȟ⩛'���\�K�G�#'XyC7�i�έ���d��O?7�H�E�x�Y���(}�0牜#V�4
T)�]yb� �"~�h�}&�	�
�~p�����e�
����>�����v �� O�z�e�%��E�&	�8Ѽ�#��=R~�1R�ئh���^�����R+̐l=|�9�R�
)R5���bD���Ó]�N8���`3�O:q!�Έ#�|-"`'X)r!�2C�	���1�gE�P��2�@T��!��y��� �q(l�ؐ�>��π'�^ĨсϦ�ȟfӅ�ՙA���0��  ��v�i��c��x��Ot%zU&Я�8H%>7-��q��d����^:�Cd�Y�Fo�9n/}��J2Z���p��Qf����&\8Q���WLr9��*��o������0`'ђZ��݅�ɡ4��`p+�LZ9���� ��pQ@!��$0��@�W���� ��"4��Á���@�	TO1s���s��Df���!�P7B����@��[�lТC�QA��!����rblU,Z1f�	�Ȉ��(���"�Xʅ8oaV=�&G	�i|��i��ĪB��,�QhAƏ����ͮL,��B�Q�ltԘ ��*��O %�sï�n����N䈰�:\Odm�`���6:��VɁ�fԋ�Kգx\��0�o5D� 3
���z��'�Hx
pM:|�4�Vj�0���z�{Z/f2aq5�
J��G�P�C�@�&>E���!{����/پ��$�'L D�h�mW�}���4g��bR���i�b����A�^EXy*�-&��|r�O��g��
��$-��#"O�X�si�2~����9ag���N�=��0ۧ�Ўr���S�&J<{��\D~rʆ��J�B4��
\�y�#n�4۰=Q�K�Mz�y�F��L*� ұ����o�t�c�K�3d[�p�T�ݚ[�����)�l�:��K�DH�B��]�d�㟰[���8P0��UH�x�:�RM~
e쎈7��4w�XЮ$4�@���B5k�#�)�0Y�6Έ�X-h��O�i�-�︧�O��T��P�j��|�pm�`$�}��'����Т5B�����'d�(�k�'̤!UXP0����RG:�I�'d��uL#`7l4ѣ�؞SC�l��'��+�΀�K�)��	H���'�"x����;L\>l���;\\<���'^��R�U�$�RI_5/���#�'��ǆ�U�DHR��Q:2����
�'Q����fA�}˾��C�, q�	�'&�d�ĥ�%�:H��e�<!�����'+p	�����~M�A-M�$A����'C
�k4ö>�V���L��0���'! L�2F��R��W,�{�ys�'S�y"N"TX0H7��e�l�!�'�&�ʱF] Xe*��Q�O�[�v�p�'���ϐ7V Xآ��FR" �2�'Ԍ�����bQ�����	�'`�0P�K@]<��ZQ��:?�����'�ݐ�*S�*iJ�����z��Pj�'K�yJ�/J�D���Q'��?u[��b�'Ҡ0!D���H�ڹ���LbY�c�'�L�"ԤJ18��z�W#ݱ�'�T�L�.9����C͒L+,��'%�ieI�.#�2�X�'�9 ��	�'�T��S�娓][g�$��'=�R'�ؒS�^�;��J&]��'�F�g�""@���Y&Ca���'�Jd9�'^*"����
�8�����'��qD,Ќ_��E��
�*gڑ��'���ۤG�����U r���*�'�֤r��ڷt�Fȸc���P3���'�8����4WΜ\���EC����'� D��	�-m�I"�W�m���S�'���8��K�VZF��"�[�ZX�;�'��Qx�h�j��䘕0�p�
�'F��)�S1P᫰�M8%N�9
�'�, �ЏX+RQ��g߰B��P�''�̹c��	f��I��$ɻC�`@�'|���BZ�]V
19�l�?6H�x�'���3��v�b��[�9���r�'�R�r�i:PX�={����=lP��'�fтt��v���J�"}H
���'�69b`H��͘���zKx}Y�'I]c "dOt�HQ*�~Z=�
�'0�����9*���`&�ijp
�'B�$��Ax2�M� �
�|.�L�	�'�>�@���H��"�O�6` 
�'M��;p��G� 	J���
h�%�	�'�z�q�fH?0)��;0�Z7E����'=��%!K-4��MӧaH� �@ ��'=����o�R'�D���@�
$ S�'���c��\;�(�À��
��'϶<Z�eH�^�ܠ�So^/z�J���@��491�su��ϓ�;o�U	T�P:s�U@����s`-A]�S�v@�6��'"��ӈA耠��=<4����� mw����y��Oa����3`ٰ�nB2цЫ5BQ�M�OF�H��'"�~j/O�S��4I��ғx㘸�P*T,�t`qٴ���şd�����m様O�2�SAI]2"[2�K�D�JLF���O�`��	 ���JA�O��L��EX2U�PB�������^��$��%n�y)OQ?u�"��r�=R�"R�HH�E%7�?0g��u)����O%�̪�π fi�D�-�0��bʂ 0@sVjֶN5�� �')�(0"C���|zF:��	��Zo*!br��s�L�A��*�I#ޜpG�M�O ��4�L�	���,�)�f%��x�ر�S�`��h�w?i��ZL>��3�7~3�ɡ��s��IP�Lpӄ7��L?�r�x���O���0�/
�q-�8�ЈY�W��#�OXxy��)�'a�"J�!ѶI�\��ӥClZ$�iGx���B�E��Y��ɟC@\p)��l, Q��)�2�;6�O~�4��(Za�n�A��I��0|j�$�p���
�C�u#��t*�p�2���֝'��"��A��Əb���i�<�0�(�Z�S4��<E��kZ�4N>�[��C����.9v!�Op�-��%��b��D��K)4��9����ŋ �,Pܲ	k�4;��\��b�8xf9���ax���IУc��Tǚ*%�:��F���Y926
<At��Z���h���e�Ǫ����W���04�E6T4�#Ь��^	��s�*��C"\d�Pe��0|1 � P�z�yc
Ca��.Kԉ�b@�{�и�1��!0mv�%����T>AI���!��U�Cj?>Q�,]�n��=Y��O��DB�B;#��X1��H�JLX���%$(�ᓢAZ���R�ْr������FB��4x�D
~Φ����Íp4�C��"MIĠdN�N�p9���%DC䉩��1��1w��u�� 0u\C��;��|�Qf��&�MI0P%FZC�ɗD�<y���3i��IP��όJ:C��=e��<�wH��~���	��M�{��B�ɛt��L*��\�7&dE�6c˗$
�B�	4(4x��P�$=6��I<{bB�I�Rդ��7$ѻ.�(�	�C�B�I=����
M�/��̸����ij�B䉚$�"a*�j�'�(� ��[�"�bB�I�D�F@Z���{e�����1�C��>���n��F0�b�T
"��C䉃Sю���cH��1a��S�P�~C�j��a��H��1���P�NbzC�ɳ,��!T+M>{	�R��V�C�I�Zp�M;v�N~�ޥ2�Q�<�:B�ɹ*�B�_�oc܅Q��͉F�dB�I6;h,h�dƯ����P�4�C�	41��I�����\�v��C��C�>=���$�8*�{e�L�F9�C�"��3!�Q�$��M
�#SbB䉽G�^�;��T�Z��J`���L��C�I�Zf&�0&�l�ɱ�  7��C�D�YSą�;G�N�C=D�<�!
�'}Xԉ��gw�xkT�T�:�P�[�'�<�9q	�:L8 ��1�T���'z�KBkF�"FYp�	U0��a�'8N����_MU.���$rE�\�'N~�I�*��.�Ęb�ˡl>���'�r�d�-7�002A��g�`	��'�J=9&�����	��Js(b�8�'���iW�^����B�P�},�c�'�4����[�N�tMq�h��z���'E�l(v(�Q^�@{�)� Il�ea�'Q|%p���$S28�KȽD.�@��'��=��,c� ���.={�%J�'�|Z�B�pۦ-;e�.x��C�ɼQ\n8�S�]��B�9�C䉧P��M�2+�R ��r���2F�NC䉭B�\Ej�ό��ٰ�E��yC�	>��� �E6�D3c�͝R�C�ɼ;��y
4%�Fs�)���A�Hh�B�It�4*�OË���c�>s��B�Ɏ=�M{�BÇU�@q�'�q�B�I�i��9�@�R��ŉ'��ޡ�� ����,� +RE�j�c"Ox�l�2B�hz�*�@v8��"O��p�ЮLM�)jՏ��� ���"O����n	l"�r�T#|
���"O
,�(�����R��]	�"O��4�X�s�f4�"�J����"O�9+��ɑW-(��*�Q"ODlض�ғD6$U��ΩY��a�"Ol�`F	�7���1i��.W�P�"Op�b���gXТ`�$)L<d�"OV�@F���7s�t��a��j�Dm�$"O�h�s�F�^Q�b�>�hs"O����Q<����o��G�^���"O�6✃($� )���Bf��"O���j�g��Ps�+к&n��[r"OLT��*M�UB�1rʘ	�Ƅ�#"O�m&m�2��0µc@�\�5��"O�t��)F��<����r*�I�"O��Sa�Ŀo��0bܭ96|劣"OR()g�(ux���rb�(�*���"Ovݣ֯�3;��Ca�8l�\�"Ob�{�M��W�lM���Hc��M p"O����lW$�Mބ$��5�3D�L:��	��}c���u~E�.D�D3�G�J��I��ǉ�S�PQڤD D�xQtC� /H�h�S�҈'jTjC?D�x�I��,ˤ��UR�+��1ɷ-8D�l@Dk.<�J�$	QP�h1%�+D�d�Т��t4�fM�gW!č*D�d3�m�(`l<��F"��]s�)D��I f��IQx݈5I�#-l-��l%D�EA�
,v�z4'C�F:5W�5D�lq�Cզ7��pR�@
v8�IS!�4D�<�M�Z�^(j���5�����b2D���-C��:,��]�~8n+D����,X�r�T�C� ��z`�w�(D��k!FMs�flQ��#���%D��8!��,*FE#��+X�!	�=D��k lG�u|v-Y�D0 ��D1��&D���lJL��Fb. ���P�&D��ѩ��?t����݀ ���)��$D�\��!�(y�)���T�!D�C�'�POB ;6&�0 � �f%!D��Q�*K�|�`��lܳg徔Is�1D��+���=M���)��`�L�R�.D����%���`�Kb�t	 �k1D��A�O(D�a�c��g�Pq2�1D��Ô��9I����EǺ	��y"$*D�����8c��(ȗ�&Y�!��.<D�`3A��2ت`�FJ� �� QA�5D�|���Ͱ_��á26#�1D��9a"C�T�kP�S=@u�a�V(*D�\y����X\�Wģ[l>-�s����y�� �N�P4���DbЩ��_�yb��?_���*F&r1<آc�V��y���6?8��FH,X� �j"!U7�y�I
4�h�Z3�-H���a¡���y�⃡:P��qmCC�@)5���y�
�?';���nپ6���AW,�9�yR���+j�	�c��E�M��i +�yR��Aκ�JG�8A0������y2�W�'�<8C�b�&~u������yb!�Ԍ�PW��%8�t '��yҩW8�$%�r�J?�X(��@�y
� ��W˄:���V�Q|��`H5"O�T���G�6fE�5#O�sx�ey%"O��ۄ%�%c���p���\lD"O]��K?5QP�Q Z17R�@"Ovl��mα(��l ��>_50���"O����ɽ[�F��B�G6 �J"O�)�$��'uipA2T��9bX�b"O<|���F���1ˉ
g8�r�"O� �Qo��$ �]z��qY �p"O���c��iS���􂞑q��8"OTP!� �"W��ʅ�MuҲqq�"O6� ��A	=�j�� 7�X��"O����@�t��9��^)m&hAP"O&�I�SY�$���2��h��"Ou�
-��ܚ��p�l�"OD��3��+��@h��nR�"O\ i3��Q��mb��#8VDk�"Oإ�׃t��г@�d+�XT"OԌjB�@U`P�Y��GE��"O�13�ь}����A����7"O�l�u�Y��K�T,D��TD#D�`�e\36\�$���KQ�Eac "D�$��dƠ�ҐK'��au��b<D�8��$\5��%ptn�<�Ҍ��6D��C�H!5�NP��Ʈ[���q�4D���J;>�Z�p��I9s7D�1��1D�<�3�L�u�x,��"�:Q�\��!D�(s�N�x[���B9�D�u�?D�X�7eÖ@���4IA�p7�Qà�<D�Hr�D�1hd�Y!�B�k*Q�ӈ:D�`���%�
9����8خ��Sd:D�(�v�S�<?�hf��"<|A���9D��QdЎ=����m�9nj.��E�!�\�L�Y�4C6`��ۦ"��8�!�DN&^\(��&�[>
w���6��1H�!�$ĕo�@ �ٳv�x�(�D��Wp!��?-� ��4�ҩs�2�`WI�+7[!�DȬ�����%R�-͆E�"��/e!�9S����AOQ*?��ŋC�Pg!��͊ج���*�V���Ia�!�nF�%��'0����'M�̬��k� �ёsdh�9�+.z��ȓS_�\�d"U"����C���ȓ+�*yb����e� 5bj����{��z0�F
�j�6��n���ȓ
��2%`*��B��'�(��ȓ7��0��`��i�	���m,R���E��	�oE���x�Fv�蜅ȓ&uB�nШT���7/�s���F�\:��H�K�1���~~n���BgN�V�������&JdT��V@�S�<�t��K��t��!L K�L�;ĉ�P�<i)
�Y�%�����x�V�<yU��	+�z�J
 ;(��;f�N�<I�f��{B� �ɤ;� �� ��F�<YР?[dUA�Idr�ɲ�w�<���Q�Jl�CCb��չ@��s�<!��W�sD����N>H�JD��k�<��@�=�DHAFE&J	
��d�<�pM���~}p�(F �Y�@V_�<Q"_>mJ��Рe��u4>��Đ`�<Y�,��M���"u�A>�>drw��g�<�b�):h��펍�R�ɌY�<1'kZ�'CR�@�dQ�1�V�ė`�<� QRW*ѧ"W�T��C?z�R"OT�� �HR���憓���r�"O�)��/v`(��U.p��(��"O�ueg��;�ȡ�'�28ꝑw"OJ�[�o�>�18R���<��"O)�ak^"�2DYt/Ŵ_�����"Ot8��iQ�WM`s�MB+4ٔ|�p"OH�ð
͓S�^$hg� Ҁq��"Or�b��5;W�ݛԣ@-A^��ʔ"O���ƢBlG@%#&�ԀnD���"O��t#_�PH�����Q5�x�T"O�!ڧ,I�z~x��a+ңZ�z8`�"O�(���ST��!�lÆy}$]��"O�Ѩ bפ=Ԗ��l�4RWX��6"O�$�#	�r���U��-����e"On�R�� N�IZ�,��/7ָ�"Oz���٥/�� �+�]f0��"O@I����<}۱I�e( 0�"O�4+r�]�-��8� �ñ�Y7"O��P��R�=���z�~�d���"O�T�q*�a�&pS�A;͢\,�!���94isV��4C8�!��/! �  ���1 0A
hp�Z�j�)�!��� �6��/@�fƞ����39�!���F��[�AW�4��ޖr�!�@�%��q��;�T�� ۱>�!�D-�8�jeII11�h�� Η&�!�B/۞Ƞw_$�E��!�!�$�	\"��S�/a�<�1���1�!�Dբ�RM��O�7X(��o�%)�!�_��¡�!A�vH���A�T<_�!��P���XU�΅:�$�W,F�+!�� � ��~�@q�]g��s`"OЍ�!�����8g$f|���V"O�<K�ώ�(�����T�oa61Xf"O����H4,�.�3A	�m�z0"OR�b�E���9��=��Q"O�}h�,��LA��ئ.��>$Ш1c"O��x%f�~bЛ�)B/h��"O A�d`?r��Z���8��<��"O���f�8)���cW�A �|x"O敢m](.�0��2/�o��	�'���kJ�4�B���ù�>�S�'>J��A¹q�� fϢ���'�n`�f�[Y���գ�Xܬs�'Ұ��.L��"l�uO7\,���'��E�\��m��(�J"����j��(O?�$B�J���@ӥ�&Vn���iR�(�!��K�+�"�$��W#��r홵_��D�Bg���$�s�L!`��m1���&@�{��ڴ�D�'\d�j�j����񆧊�A&�%b
�'F���̠Q|(�M3E� B���ՁG��\G�d*	��l� TO	C6m�P	M�y�"J*{����Ĝ?Gk����i]$,�����,�B��~��ӓB��@P� J�6'\����/�y 1F�LhR��3T�J�sP���?yD��"�h���ɀO-h��$�:u��ᖥ�$o�{�˟m_rM�'���2�]hE�)r��W�Ro�d#
�'��L1�mִR�VĪ�l��Ug�l��I��0|ҧ	�a�F�XTҲ}����w�o�<A/��t8���V)Q���k�e�<�Ҥ��t��d1�D�g��!Ӳ]�<�����r�l�;��'y;�5S��]T�<����l�|�@b�*[��Ђ��T�<����,>`�Y��K�+N{�q�G"�Z�<	��O*I�Đ��?!��+т_Z�<�����x�Q;Ĭ,�@��V��h�<��Q��4�F�қ�)x���k�<!�MH.^X=��'��"Z�ycJ�_�<�$�" �6q�"�/g�!y��XV�<iq`܄x�6q)en�H⸐���o�<�`�a�����D	#@�`�{o�<I�߅.Έ�� D�+ތ;3gMN�<��\T���/�^�u��A�|�<)f݄\bZ re���PE���5�^w�<����~��p�GV�mo�I9u'h�����Ǚ	&yf�'U�>��(��MXG�4[�.hs��?5�B�ɿQ*2��&n�H@(<�GoF�!�p��b�n�Pm�4��}�b0
˓_�,	YԮ��NE�0� - �����	�#El�V��Bt�W	H;B����e����|{ �x�*�3�
Oh%���[����"C)?�g�|2��>�7!�)�E
���?.31���S��ư9S�t)u"��>�(h��"Oʙ�1�U(}"xT�D�d�D�B ܘuR��G"�CD8R�/��( ����-O�)�%�
M��+3ϙ#�\E�a
O��˂�\q���J�\�rW ��6����58�jɯ{���R:h'�*�N<�C�xf R,�f���&�1/i�ą�3�d	�e�ݞ5��eqS�N�N�Ȑ,)�B��v�_�t�!��͋-� 
e��4�p�|�x�yq�H��TɃ0kG�	�4d�heiR�bޞ�����t�Q1C	U��J�Eإ�A
v���f ��& Մ�d����@�g�!������1l���S-c��9��&�\ô '?%���']���Q�>�p� ҎQj���҄$�>e��	6P�6�Pv�!`L�q�A'�%Ww$�##ʹeb:<BVd�6q"�g@ ;4�X{�c�'.(���'��~`\���K8peV�����I���C+�إ9b	O�h�@��o2p)C'��%N�,3R%[�	R��#7�OԅIf��(
���V��Uv��V��J���+F���rl�)k�ʃ+A)�A��]����2��[s ��d�DQ�)ݡ�y
� R��֬Ǫ8��`.ֺTZܡ�ak�9n�d�R@#�)�t�S���*��O�d�c�ݫ��Ļ	����<HݼT���-I:��c�:�Q����8\�̥���X_��tȤdەx���ݹl'�9�E̎OL�M�p�/p���.�&rH�hh�/�.(b��?�����y��=b���	"��|�L�a�R;nX�2)f�hp+T?"���m.ĨOš#ʺ���� wݦM�'��8�fD�j��Y�歚�<r���I3mF����?�ېD�7>���Y���9w�)Ԧ<D�ȱ�l��`1$�U�U������>�x��F�JC5��0���X9{Ul�3��	�z����Oɐ]V�mz�CL�Pd���۝x������)k����fB!ی�P�ʏ>tF��6�K?k*�=��Y�F����s'$�:h������7FYF�j�F])R�p�F"�
(�y!勐p�^ٚ�돘,+�l�t���I���%�Q�T�BD�<aǎ�]���Ӂ#��`��iB*0�RY��d�<Q4h�'�̨卒��`�XB��A�|��j�;��)�
R]I���fvhhv��R(!�d����$)�,"�bH#Ή�7u&�Cq��,M�@�b��7�x[3��do�5�pK#7O��$N���`X�A7
R�a�O�.�@�pQaK�D;u �� 󼌢u��]��I�W�1P�)XCH�@��D��lxX�Qy�>�z�΂uaxr�C�_��ܻ���u�3�`I>n�.B`Y*���AG�k	�=P�hR ������"��oA�	�ap��O���'�P`�T�D�+$�;a��9(rA1 �O�0��w�Lqڬy��ü	�' �%��nO����� T	)Pb�|�*��D
��x{�LP ����O�'u�Uj^��U�d�P(,L���?4�0{dV<'���b�s^�0�R+��`�S0b�s(�|�eɃ-�v<��	#/����!��VeJ`��\�"�����3'6r .W�u��P�~��)����pcm-���'��!"T�T6�6�z7N��msx�Y�{2�G�8� C6n�!K�v���I��5��|�Q�F��	�:�!�E-bp��H�	b�f�@�,J�Q�Z�2�A� m��(�[��F��'F�I0�S�X��ғ�#l��Qc�'e����¿�� �f��Y�'x��A�`����X�K�4QC0�A�'��dW(`+�1�Y�x�v\S�'��`����4pk��ٕd*d�0
�'��p���H|�v�Id-�m6���'���s��/����[�bp����'�,���@n$����*b��'	$�#��C vg1��=2D��'t䡚c�ޚ^0Xj+9<��'�]�)4?��b�$�	cdEP�'���F�"~��0i�!!8�@K�'Ō�C��)Bg$�Dܯ;}�$b�'�4�x��N,<2����[�`'n���'(�\�d;6�"�AN`W�a[�'Yȁ��#�Ơ��L`�����'�����Oąl�f��%a�]�,t#�'�Tٕ%�1~Z袔�[�6���'	0h�+� 3vq���X�L�)�'��|���a�j���]�:$��Ӌ}2��z��xR厂V(�\{7�Иi�8�#�Ŧ�xr��Ubi!mR"+~���,A�7�l��C���x�]������u��P��Aܑ��Opy���F�w�c> �o��i�6K�A4xU�%	.D�X��)^�Y�J ���5/-�2�L�<1qdS�n۪�@H>E��F�9����Sm�쉤���yb�2`�f졅��@��ly��D���B��P!#��0<�I̓@g���k�Y����{�����)MS$2�*s/׹dڈ�9��	��^M5�l<��oS�IN2pY��C�R|���~�'(�p��N1� T:�J��d�zH"![	� ء"O�0A�SN�P�p�X�HR��P�4��d�,	$��|Z$��_Z�b�8V��C�*�A�<0�M��@4��4��|�R-�F�	56��T���_F���4�ވ����D��X#��#���d	>� ���թ��_�j�;�A�,}����C*��]�!����^�yڦFZ=;TD���#�ay�-�5{qO>��oF�I;�)���}��A"OJ�YS���l
��ʡ�оY���"O<-	G�@�T�,�q���z���"p"O���)X,�fQ6�((��a�"Of̢����'-��RB� l���B"O��fI	�O��� �3~�A�F"O�)�DV2mfl�F�U��&�14"O(������t�af�(*�X4�3"O�!"2�ú
z t�u%ƻe��8A�"O���H$��h ȸm��y�"O�Uì�66�$u�AՈzv�H�#"O
Zb̚�Z���	8d>mC�"O��c���wJ���ł7.w�k�"O��c7d�*=�h����]����;�"O��x�IQ�w�.�q$gRJ�>d��"O("��Ųa�@Fεi�4�kU"Oz�t�?���LҴ`��xR"O*�z�QhBP��k[6g�f5D�h�ըLL�yg�n�|Y���$D�LpW@��D�����P�"(��� "D�4:��>i<@=��,ѲJs6���-D� �cFڻF�p�P �'lp}x��(D��{#,
+=�`2F��"r�\�r�4D��R���Mje���6���ٔ�'D�8��@8��db�E�b�ƭKd�"D��@�@~��8h�ʃ;qFt����<D�\��AG�@�CA]/*1X�CT�;D�,R!*F�^�x}��ݥtll���-D�	�40wb��V�D�l �����-D�4yÉ��_l�ɷ&��h`P�4D���G%�V��s偸<�NHhv�2D�<0��8%�90D#�b?�qd1D����T7q�$���$�y���/D�ĨTbUl�<do6W��1Q�K(D�Ċ��a���p#Y�Hu�4��%D��p�(���R����GA -D� #��O��b�4EԾ!K���gL(D�|���*e����0"3��H $D����%>A&��pK�5���pa
 D�X1 ��`8y�Ѕ�6w�p-�!��0G����[&.
ڨ��Ǌ|�!�d��bEPmJ�&<��˂��?
!��O���1����`|(���<k�!��I>]���ʰK�X4�G��6�!�$֨2�lstk�+?��87��)�!�d�Y�8i�闫KKx�JǠY.!�$Cz�P���7�r2 �U!�Dzĺ��V"�*�:u�Ѓ3!�$� $�4m��=K���PE�ԐP�!�R;�$�[���+qH��v�3�!�dذcije1ч
�M�6���J��Lg!��%a�h��!���,(��7g!�d�aL��ԍ��o�ԁ�3�Ļ)]!�d�v���&�Ԁp�b���-��Pyr�H4W�@@#�Ĥ@PƘ�R��y"�k'����/7F*�� 
�yr��x�.pC���%���l�'�yBH�dFz��u�X���(�яQ�y�D[p��};F��t�` ���y"_�0Y�}�"6�N�(��)�y�g��I�4��1�-�f��yRP���� TlX*c�\�rU�y
� �\(�
��x=�Q�K�<f��CC"O����L�-q�$:�V�>��Ct"O�A(�GM�I8P��k���g"Or��λ/.dY��&��D�*O�-"1��<L>|�rQ�>D����7D��c&��j��T��J��	9"4D��"�W�Da&�I@fT4s��px�` D�0х ��h��@D�.Ҧ��e
%D�@�c·<-\����+y�VMk��6D����'L��Za6fX���0P�j>D��i�ɒ�&R�U8#L��z�x8�3� D�T�
G�-��!РR?:�|��g-D��Y��3x�����̟�]�(S!�+D���e/ݏS`����F@�'�j<*C�&D� � ԧD	����j[[�|4�`+D�p�3��(j^<��\p�D�+��&D�0��Dڋo��P�H$nT �d�%D�0�5��A����R��2B���"D�)�@�62�	��=R�^*u�"D��27`��i#�ٓQ*	�z��7D�B�V1zq��g��(�@]��5D�|��Y�� �Pz���*O��(���-2���qAŖ'tڬ8'"O>�0'���O:���f�A�D��5��"OޕÑ舝e�����ǟ><]�a�t"O�$�0�_�8����<�l�@P"O��a(�}|�!���ʉV'*��"Op��À�
r��!BFN+q6�k�"O
����%��c"ě�%�*��R"O����l؀Z^�Q��=N� ���"Ol(�C�ڮd��5�%&��"O��e�0-V�3 �:r���T"Ov�xU�2Uq��JWNٽJa႕*Or���dƈ8'�d��aG�1o��3�'���0�ŁhGƩpU��!5����
�'�$S%%��'�x`�6��8��'��P3��H"9�b��!�p�X�']|B�iʋo	��2�Q6t�Vy�'����	)%`%�Wo��H��'ߠ<�rX-�s��K�Y���	�'��D�$��rvZ���)Vg�x��	�'+N�b!D2��PQ��R�@ub���'�P�	��T �5�Wi֩C��2�'�P�gJ�T�\�B �G_�<��'����+���C�'�,.�t;�'�jh���×L3(P��
Pٻ�'q|����Km0~�`��ݗsX���'kP|СF_z�p4'�Av!j�'u8d �S� �s��<rr}��'T�(�g�;�ܰ ��Ӽ<�b�{
�'��H#H�QZ�J��όocR	�'3�'�҉D�!lٴ`��'�8�S0%L&g���r��8S���'�:���-�7�Z(����%&�u��'�� R�9�p@k����(��'j��b��@f���h�+f���'�(k���G˞���*\K3

�'���ҙ!eh�-~�;�'x.����>c��h�N v�N@�
�'�4`���Lϔ�:Ԫ�e�@�0�'ݒ����:l2(0����,|2
�'���p��p��!b"X��~-�	�'�|�Ч��pJ���1��2t��h
�'�*%�r�̱��m t�԰a�6����� X����	�L7�ДMͦ��&"O>��I�y�D�&�sS浸�"Ov�(e X/Z��� �� {t���"OƐ��MD�bx~���Þ9Rg�T"OR��N� ��<آ�ΐ/^H0#E"O��+���5KX}:��J�M��]��"Ob5�0摺.�P����מi�J�"OT�`�@V�,g~�����9bֲ�@W"O.m �E
�_݄�у%D<����"O�@�5��:56ҥ`s�<G��l!�"O��)�]ݬX�υ�m��送"OR�6	P� V~�/�-~Z��6"O�-������o��#�US�!��!=�T�c̑�*�h*��ҏ d!�d��9��|�� �(i�%@6
E S!�DVJU�� C"H�qV�l�`
�9~K!��D�7}xݸ���[G>�z�ڍG>!�I
PO8Lp�,55J�m�eț�+�!�ϰ�����.�>/N٣gڧ&~!�D�Q J!�ՀZ� @ �D
g�!���i�v����N)��#c�\�<Y!�K7]��'lѠ4��`�$�<4!��-���#&I7�� d��f5!򄐅?�Jl�R��-dDu���2&!�DʭG�.A�ԀS!A(4-��	 /!�/N�5)��G}epiQ�ظ?ܡ���!:�����b� ���y�bG��<:cm�y��*����y�e(X��"��z��qc���y���W�Na�1A�s� �`@�,�yrh�H\����[�s UÖ퍧�y�`�G�D�W�v�|	�E�8�y�d�#
|*�w*J�R�V��u�W�y�W���k��PK@�EI��T��yb1�"��C�%L�>l#��^3�y�țh?��8W�
G=�ݠ3N���y�f&oF|i�F��9@qKCaߒ�yFG�,C�9�s�=:����HC��y2HǲQ�Uv�� )ڎt�1��
�y�)/5�n샓��t<�SP�S��y��I7J(43��4W�2Z���ȓU�.�ဋ�(�D��Y�H�ȓN�H�ĥ�3�)�q���a���BI���H�,Ҽi��@�\�ȓ-�(��Wa֚.H����e��l(��|�ĵ�6AF�%���A씿b((��HU��'gҊb)(F�; ^Ԅȓe�����̓/Uly�D�4��u�����ې:������$"���4TR��&X����'�[(<���ȓB�l��%
�)Zm����j%�P���:�2Ǡ	ۨ�C�J42k���ȓn�vĪ���3��4�J�dUZ8�>6����p<�0Ȏ�4��M �LS y�����\<� hN�9����,��yA%�q�Ŷ���s�\k<)3�_8̸$%I�p�� o�A�'�S��'�1��	q�,7X<H�a�wŌ"�"O�(d��N?�uYwo�,p��٥Q��xw?.���&��|�Z�XlS��� ̴ �fnV�<��G	)~Gᳰ	�;`��]�fg�R�c��q�ƇR�<[T�T8<�,`Q�ֻj��չ�k$�O@ ���3H���G�8��m`�m�0�d<��hW.mADmB.��d�M15��6_�9IM�8٘Oc�-+���(v�\ �(�1!�l(C��� e�� �K*N1���� C2�;�Y�� e(R1x�$��|�DL6�������`�m�`�<�Qo�&�b���Da�1$TV�I��JI��ĔV�Xi��:`��5�6�C�mnx��:�PqRL��utL\c1a֬9���v��!V��D`�$�4���ǉI�p!R �¦Ew�zd'*,O�b� :�ɔF$i�'�,8ɒ�/�bB��]B�A�b�(=�6�H��r?lB�ɽ5���̗l���N��:B��'���%B 3<4���'OB�C�8vA��o#�~0��d�6�6B�	�A���ŮU�I�ZD��ԊfI�C�ɶ+IP���1A�<�S�S�1|�C�	�[mn�s�/ղ+��;��P�VB��+u���hT�D �*@�Q�nJC��5W����+T s*.Y�"C䉨m2�x��7.��J7�Μ_a�C�	1?�`$���T���	�O�8B��C�I�!l�����V�	��U� %�x}�C�0F.u*�!�;�: )Ԃ�=b^hC�1^�����M1E�����ߖP�C䉞d��q�6��z�=Xè��G�B�;X�:,9�d�7C�eJ�$�=W\B�ɳ_Ѱ��5�S+5>U�G���F_,B䉧~Y��qa�$�(Ԑ4I���B�I��.�[�@G/{�8��D4Z�B�I<,=i������U���B-24�B�ɇy.ʩ[����<��=b��?S�B�I�Plr�_�L���IiTB��-D0�!����*��PӃ��)6B�ɑ2�$�V��}�bp(#/ķp�VC䉵_�6S0hM�~�\��S2bJB�	�r�>�#�[)F����٥k�.B�ɰM�8^�s��=J���`(�C�I4S�^D1��E�u�je�vI'v1C䉺Xg}���U�d�RaT�F�pw&B��&�=�Q掕I��)�է�X
�B�ə�>��lVVd�"��1ǂB�	n���[�D�)1w�=��?+�B�	�w/1h�ʌ�U��yB� �<�xB�ɫR��`��,�Xp�_�%�C�+��x����\�#]8�0C��%�:|2���g��H� ��fC�	�l�����&i�ސ�AC�8U�B�ɇ	*7EI�uL��O�2}��B�I�h]B�3g��`H��)É����C�I�.��<�lծr�*-�1ϛ��C��|���@�H�V��I�`�@�VB�	%L4���'�/$��2@��%MB䉶	��h����zn!2�j��nC䉰ϼ���5)u Q�jP�B�I/oj�Z�ؙ~��, �S�'�C�	��T�`�9C�@�4
1B�6;v}��n��Fcn� �)yZB��;P�h��e��E�	��珒k��C�əM S���X����*Cv���$��3q�P�a%�ܘB��_�J�O����O�t�Ѧ�_�
Xs5�ƺvR���}����O�O�04p��߸]��4@�+����M�K<a�hT���O�(�!�LԯslV|Rf�V�u0E�*O̵Q	�k���Bs��S�����9l*���I{�y�ڡ�P�),e�}ZWT(�d�iў"|��O[^���"f#μ(���<^��}��' �O�O����W��Kc��v
�/���qH<a�����O4�EJa�8||��!6z�н��O��+��A��� �� i
 +�-��c�?��$�"O6m��$͏8�v�Z�U�w����O$4� mL� s@��%�i5z抎~�����aq��0�iF�P@��B�X�0v�� E%�#/O`q@�'�H �OQ>�Y�.?� @x���+��|Rb@�O@e��'�jM�������X�[6)ԟia��2)Ӓ �&��'��H�=i��I˗f�Vi;�
�B�h@EDY�6f���j�6f�i;ҧ{��u��Tg@|5A�
�l�0�g/�D�̟�`I~�0���8)FĴ��b�y�.�p��J!��DB
!EB�3*��)ʧ�KQ�L�y�ㆩd84ac�O�����'9l�B����~�3��b�� dʔk^N �a�Q8�*��/	A����	&�'/
�@�@ ���p����	P<�nڠz
�'$@������ʅUƼ|qS�D�T��M*���:��}�/�N}��Ǜ]:RP�Fk�C�,!q��ߧ��C�.�<�SR��'-�J`�C�ɅQ%�4�����>9�I�&D#<E�T��$hӎ��60�hUA:�M�M��#>�O����<�d��5�"���4���aF@\^�����?��ȅȓ2ɚ��������
լنȓOJ-a"�ǈt��|�4 ^A4�ȓ1�Y�d�R�>k4#������`�)A҈ȹI	2�:�̜y4z��ȓ >���/Y�re�`Qi�7~���ȓi�*�JEnR4O�*(�7Y'rd�ȓk�@4�]aN���_4+���0D��)m�2���L�Cm̠۶h2D��K�B�W��MP�\9 E�����1D��X��:�{��$z�<D��	��΁2�"Did��[^X�w�;D�t�e�'�]xE� Vt���7D�x ӧ�,E�-#4i�S�. iV�4D��F�O=/�J��'&05���2D�����Y�r	���O�[:�{ �1D�0�L�N4���I\�SQ�����-D�Pu�՘?��YR��V,��q�n-D�кS�Ej��	�D��6XxF�B�L>D�� ��ǻ`����C�@��@/=D������eJ&�٦��6KѠ�u�;D�����Ƌ��ԩ��ފ�����-D�TсcI�i�����Z�a,DJv/!D���6�A�8ruQaL��a^
,P`b D�*u��X�|q`�Y3e��݊S�"D�\�`-�I?f��嗇���$D���D����v�I%��R�,D����Þ'�tQ7���)� ���=D��Ӷ��9�X�Kt��0� ��� D��"��"=�N�B�BÛy��!Y��+D�c�͍x��\pqϸ3+�	#!l,D��7��s��(���ђ��B��<D������=O.�x��ӱl1b([-?D�d9��C*�-�s�݂ѐy��i2D���K�s?*xx�M1D��(��2D��Ǭ��c]�� 6A�!d,2�A]�y"�
e�$�˧EN;�@� GW��yBl"Zay-�3��ɱŖ�yB`��1쌰��'@d�]�yb��3�d�P��?���/�y�C��<�$�.sm~|X�g��y���qf|���5t0<�d��y���z�����U�9 �}���ڄ�y�D�)%�@�{���+�X�)�٭�y2�M� g^�r�o�'��R� �y� ֋d�ɥk�����Z�c��y�`+"�z��c`K o�Sc�H%�yR	KV#2�&�֗u `X�5�y
�  E�@���.�¹�qҳ?T��ӱ"O*��`X#ž��V���>m҄ 	�'^��j0���n�;�c�*K��		�'���1K�g
"�8EI	t�HmB	�'x�E���Uд���ȵpm�QS	�'���B��KUc�����ܻS�6��'K����O�1<�x��F��7]���'����\�<�{&� .�� �'��8�a�3u���§*[Ǧ�j	�'E�a�5��%.��ja��
K�R ��'60XB-�!W{��*R��9FF� c�'��iz���%?0�(תN�uo�(��'p��A@쎇+�Y���Q�gu����'�V�p�T�dJrY@FɈ3It��'S��RR@�z�nT�ulXE@�Y�'x޽
5MV�g�FY#U�H8�*� �'X��ZU�Q"���KA�0��
�'�9"7N�"9eA��2=*nA�
�'�ڱ�!�ɋ&������ύ91\�

�'���$ͮYS\4s4�0�XA	�'s��A�=P�J��Sb%S��9	�'�CS��P�ր cϝ� � ���'�� &IQ�n$�:��'����'aDd�g&
�q�-��!��LN�y�'Ҭ���N 5�a
tA͔ZZ#�'x��T�;1�B"Qo0���'�h�9�A'M���Q�iV�OY�,
�'Ƥ5�e���״H��	H�b�'i�P�#ž9D�(+���sF }��'�����ہ*�����.lq|��'w:����1�:ɰFI�1czـ�'D���oc��ȡ��M&W��@�'ڀUd��]��r�U�ZPH�'\D;��K�\���"_�MG�-�
�'�H�4�DD��Q$%oj���'�r�{G�=��{f��b���''�LQh<HX%Q��ݏ���
�����>d�I�Ҭ��/Ҁ}����S/!�d�z����ǗD��URQfZ9a!��""����@��/��QR���1Y�!��4�~� ���Z��G�VX�!�ē�c�X�spE�b[�pP��SCx!�d�bZ�؃�˥vLKXR�!���6sP�PGgٔ4�����њ(�!�d_6_L�(�gW,H�̀�&�!�d�m�(��-��+-F(��Ŕ�n�!�D�7Q� ���
S��:��R�!��؁_�0��g�aݪ�G��c�!�F�A���#P@* ���BJ�!�D\?���j��X-��q���ׄJ\!��Y"dOP`q��&| ��+�02�!���,q��.2�
�@SNu�!���8
�Q2��4�M@�o��S��C��%��+�[#W�f1(�	�j��C�A�x�Pæ�.LJ�:�c�5X6�C�	x�d���o���$9P�/AxC�;#B,�� �K�q/Ĵ�C�C�	$!�.PN G�ȵz&�S
V�4B�I�)��[���I���S�H��,B�3h�,X�#E�U�rA) �H�@C�	�`�J=qQ-�1WZ����	�,�.C䉽t����ᎅz�|,���P�
C�	
v_���U��'I�F(J"�J02��C�	�L�0y�4Ly���U��C�)� �	����L�$���ʑL9
� "O�(�\}��}Y�ӿQ��T�`"O2`�0�M[�v�a ��-xx>�S"OX�٥�GɈi�i�	iid"OJUd�N�$L��bJ�*S����"O��b�k�J)b��΋�L5l��"O�8i�'
i���F�$-z���"O�3�)T=��A�KQ�����y�b�;U��[R&'c��Œt�!�y���!K��$��\�WЩ�6f���y�Ry$��JJ�ps�?�yRH�d0���$�Y�?}N8�щB<�y�ڸ0|����7�
���J:�yB/�Pc����.�+���G'�.�y�n���X���&��� ���y`��2�i��k[W�8
�����yN��Jꤺ6J̡z�X����y�J�?~�:�೧�8[^�k����yB��6_�r�ᅯ�7M��8�D3�y�b�=Xy<
A�@,ta�!q���ybE�:
+�tj6S�d���2�)��y�X�T0|1٢�P�2V���0�Z��y�e����A���,W�x�L���y�"F ��ж!� �N������y�+�k����M�"!� ���^�y���s��I ��&�\�ç�T�y���^����tls��B�y�f
X�HXQ��f��ɳ����yB��,%��j'�̬j���3S͇��y�M�&k��\�@\�R/nmx�	Κ�y풀`���5�W+0�ˀ��y�(��":t��u�_)P�N��D
�yb�Y�+4ܻ������D�չ�yR���(�j�P�
P�`�S����y�}D�1�	 f��Aiш�yҭ��{���I���F��&C2�y2��3Y��)#Fk��?�@{�ѧ�y�n�& �%s"���h$��G���y�i��Y�X$C1ń�cĸ��EL�)�yR�r�x�
'I$FE���k��y�+V��{��t6�e��ߝ�yR�͞Skl!2�ꇣ�,M�fME5�y�S(�hTGG!B��m�u(���y�A�-Jqő�D�bUj��y"��,j����):�Ȣ�!���y`F���1-j&܊�#���y�(�Rp��u-/��pU%Ö�y�H��D6�Ȓ�͕Vz=�4h��y��Y������;^�����4�y�=]��P�� �NNё4��5�y����<�(�R��%J�P!�P��y���8�LC�'��;��PC�O��yL]�T�p�k�N�C/����[�yR�\6p��PBk��3�v`S�V��y�/�'�}���(����y2FD���ѪG�V���\q����y�@�T��%J��
1LJ�e
ͱ�y���
1u���'�H�'��}�.^��y2O��e�z}���O�k.|��v L��yR��:�A��Ɋ���Í��y�!
����ˑ�V��z����y�e�j�B�"�b>�!홆�y�ꔑ:!h����ݷF�H���m� �yHE�\n���;`k�P��y
� N��č��r݌切F) ~��b�"O����������Eν&p�8��"O
i�G���	,$�1�Ιp��S�"O�y{0�ߥ� ���H��R�i "O�V�M8\�l]0�k�hG�I�V"O�a���!I�XD�%K�5�X�"O$ [孙sm�` U��H���"O6H�s�22�rT���/'��)"O���v��`�ʌqǮJ7w���4"O�P�QĞ�	��Ea.C���9�"O���ʒ�O���YtJ$[�N�*e"O�X���z��Q�S�{|���!"O�I� �M�d-~٣��1|.���"O �2�&��r#��s3���\"�"O�@�G��@�yRh�?e��6�4D�p�&��&*�����'��p��ڗ) D�D�� �j�J��&m����;D��[��ƽ#F�Q���q�̤a7(6D���ħ��7{r��A��#9f�XZe+5D� ��V�w���j��S.l8j�f3D�4i%���J�x�S ��X���o�`�I�_��-ǻi2�)��#�-9�iJ���s^:":(Q��2!����$�O���&��Ux:/Ƴ8p�Z����K3��W���sÈ8Xx�DhL�3,d]I�P��PQD��rʙ��Ǧ?���N0	��@U�b$��S;*""!)�(Wmf�UqF�����J }��f��OAm�7���Oı��Yh׆J��"���"X���>	��hO(OJ,�#��H��:���6i�X�I��MS��i��Mx� ��{�5��N�#o,R��M�bۼXJ��D��?�+O��A�iU�����O����O.�;�M[��Ѿz9��n����GT�7m�]��̑	�U@�U!:�����r�n�r��i�'4���-v��xAO�[� �� �{7�mS���>p�eʇ�-G�7g�|�5�O�3B��D*��ґG�U_v0���<Y�N�̟<������?9��M���.R&\�gG�2p���g�t8��:�򄂖˪�P3��U�[���#��[ݦ1�ݴ�䓊��'��]>
�x� �;��Z���,!�u�ǡ�:O�.���O��O�X�;��)�O�U���5?\^���L�1[h�d�2i� ~8+$���N�����,�4�z�`�)u|Q��{��-/��0�3�W�&�*��'�7��	y�������jn�M�����
p�B�䅸S/���&����%���B|���dA�-l�@�$J������s��?I�C��T��I	�ϊ�2�r�%}�'��D��)��fl��V'Q-�m!I�Tش��]�d�3D�4�M�����D� 0u�
.ҨA|�H86�H
|$H��m8���ǟ �ɀ�1@�dٳx\|��5�ŉO̬y���jy`ISE����4�J*F�h�e�;�xsT�*f�N��tva�`�fN�ǥAL�Pv42���8�p�7'�9?�R��ܟ]�rq���mן��	� M(`g�!&t��&��k����?*O��S�Ovt�k΀�rs��W��;'�4 ����M���Y(��<SЏ�qj��җ��	�t�Z-O&�"`�X�x>�d'���Ru��fӒ4k�e�2�FT"�� ��)	�L)��J� ��8�j�@S��Ҏ�F�kp�<j]w�r�R��^<n`�Wi��Ɉ�O^D�"�.|l��E�L,ZW�)��I�C�T��'��)G�تE ��:�&���$V��������������b��柚Y������(e�$h�f#Y4�p<����?)H<�"m�mW t%Q��\X�DQ�'��7�˦��~:�
�7F{�-*�,&U ��r�b̊�^�@[��<+�T��	����	��X[w����0K�HѠ�ںB/� dP9FÒ#�@~#$�!NF�b�Oi�d�:!��C)O\M�r��2�$A�W�����X5����h+���(k����è�b���O����g����/��<�q�[�"er��rA  f���U�i62�.�B	[_�<����M��	�.��AV�8�h�#BR\�'$ay"�Zs�`<�w��|��n�~�Ls���nZn�I�G߮���L�I�6#����7Q^x�`��̴�
�'G�I�@  ���   E  �  �  ;   ',  �6  YB  2L  &V  �`  �k  qt  ��  ۊ  O�  ۗ  B�  ��  ɪ  �  P�  ��  ��  �  X�  ��  ��  +�  n�  ��  X�  .�  � � � � ! �' �. E5 �; �A C  Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�� |d��"O
`�(�;���8���-0��1%"Oj4��ND^[��"3/9�0|H�"OB���H��*�ʞRy=a"O�味V�!X��!&F�:J�$���"O,��a
���C�Ą�M�"O,$3%o�-���p���+Ն�:1"O��ݢ1����`���y14]2��i�<�6��{_���c�H�`�fX�$Kn�<��A̼VI�xR[�)�Ć�pඤ�ȓA5��('nߡ4�� �)˩%� ���,��r�؊b#`T�eT09���ȓ!�b��g��}�8�F��-? �ȓ
K|m�ș�VṔ���2�%�ȓ"R�X�j�4JN�1�˘X�i����̹	_�jZ��1!g��zܶ��ȓgil,*�J�
j�Ne��i�J%b���f	�(U��:���G��$Y^م�~r�� S�%T"���k\�jx�ȓ|4�1�îJb��@ӵ�ݩn�V��/[`�"�v4�R�!ʎ<��M�ȓ`:��z�ؚh�J�Z��$HY:	��H��p�m�C1��!��B:��0��EnjZA V;9����J[
2���	��4'J�EA�IVW&��~�(aZ��ӹ�>� o�Y�|�ȓ�f�A�
Ο7�H��M�$�����mޠP����/���ANXo*�ȓTv�����{ ��-7�*h��I��sB�8�8���3����ȓNe*M�悡;������X�o��!�ȓ'lj�#F�m�+R&;�|��It�'m"ui��G:�X�yc�\aR:�HJ>a�����(O�dD�'�H��kO�j�8�p�'���_������ؘJ&"�1�d��w��C�	4'��b�b�K�,��+H�"^
b�hDxR��N�/a�!��c@�.(��������L�ē9t�]�CњP�~�"a�ǆ8de��[l�A��ˏ�e�T@B�k�-����y:8ta�BI'4(��#�K*����	�'!J�ss�V�3��(
�������'���ق��v|L!���b���'�XA �~� g�Z&x0�!��o\Q�:0l�%�8�X�	�9~�E��?D�|��ɟ2��}��B�z7���F=}��O�7M6��?��H:�yQw��5�,�ǀ_�"n���d�<٣N_&0�>=QeD52h��;���,i�'���S�g��f� q��π(G�F) Qj�����|���"�>>��%%S.��0?�דT��IC�� 7���b�7v�άZԖ>��O?�$V6l'�c�+GZ �Ϛ%CnNC�I?�*4�J��|A\٨DcZ<<�F�O���$��B�>xb�ԃX�{���o0!���{��I��I�P�)Pv1!�DT/#T��R�/�q��!�e�y��ɟO��@��	�/�	��B#sS�B�	�3�Lj�03��-�gOEdʓ�hOQ>{��O�0�(!(��8c�#D��ҀN8^�>U�6�L1U���%!D��)r�C������y춐i @?D�`���ïU���	��؊�?�;�S�aW���D���(�f�^�D
���S�? �4P�Hn͚��h��{|P�&"Oh�� �J�)��L��m�@>�홵�'��0��IӶeL�װ��'�ˌ",H��)K��s�ܖ ��\�&�*Tj��?Yٴ�hO�,�����K�p��B���U�B�I>m���*bΛ	y��<�ť��E�PB�I��vH���U�dSU��3{{�K��)�矀�"�:` ;��D8$�=HEB*�Ű<ѳ��=y0Pu1��� n�:���S}��'���"��|���H(�V�{�<��K��={��B�ƺV����ܓ��'����v�8<\���,͈Oi4�1�O(�����MZԐ#�X�c#�P����>���M#�y��� ���q���:!%6�!��[�{Q~P"Ԉ�$	�
�r��B�D���_x��F��I�μc��إ�$�3�.�>Y�O�b�"}�͍^���hD�F��*�dr�<��Z�A=N|x�-�$5Q +o�I�<��	��^FL��	'�����Hx�(�'j�Y�v؜Ds��Z�㎞J� �������4n�rY!��N?�\q�aE%�Ɖ�ȓq�@D���̇[N��KC�ޡX|�'����I3����xOd���(�*��C�I�l��uc��.<�8#Ѐ=��B�DN�!/֤%�|x�C�P�.��B�	�5ݤ�z�`�&3<���O~��$?���)�b�#�#N����Hf^B�	'&:E��o�0}������U	2��G{J~:%��^�=��F�*/Ո��H�'�ayB��O4P��GL�������
��'}azBm�l�^�(P%��p��yJ���$�y⥗�p��kS��9a<�܁BF���O># fH�V^9����F�� �/�zx�@�'c�A��O�E%.��q �������'��𯌿L&�#���]r�J�'H�8:g���쮱��Ŕ�?�uH�'�heQ6�X�ނ�Z7��;�"�K��wӔ���P�Y�����t���q�T#v�!����P
���"�(a�w��/��N����g	K��TAʷ��I�x|"a`6|O�b�Ȋ3�ڏv��͠�Z�U�B�Y��4D��CǍ�,G�U��Yz|>��@.��蟶̂!H]<n�V5�����a)x2�I\�$�B�@h���(ݽG�<B4#1D�􊒂_�q�T��@+�Ƹ���!D��p�'�sFHq�I��� /#D�ĢR ?��̫T�)\٦�ZE�%D��5��?���p�[1g���A&�?D� ���«�8!��$z�9�u�?D�z�B�RȠ�:�"� J���A7. D�"v�'J.�(�!�18}(���j=D�X5bP�dҀ3TG�P@��f<D��1s���ܐ���ů>����b�:ғ�hO�+N�(Y�J=��!�#�ـ�vC�	4G�4A�G�I��A��#�f̎#<����?m�T�kg�u{�_! �H�"�g+D���Y蜩@G�9j�r�
V-�=�,���dn��%��*kJ�����?�QL��?�Jq��ض&@�T����w8�&�t� JH�G�`�P��0@�ȥ��&%D�<hSD�'�v,`Q��4L����(D���%�Ҷ/Ѽ�����1璕�s�&D�ԛ�,�S�Q���,�>��#M"D���&��T�pL� C-s���!�Io��� �)*`,�;L�m���5tU6lY�
OP(��K�xq�8��{�$�+���&�y���)w�%(��ʐAټd`�����<9��D]�q���p`��&+KưX�!��44���#8Ƃ 3���9��d�p��������߇]M�H��+`�ʦ"O�b ��l�q�ھW]�L e"O�h�u���'��j���Y^rpAG��>⓸�I/��3W�دC�`��f
�y&B䉈l�,��,A�4@��D&'7�C�	2Bp��(�iޥ����+M�y�C���4�s!)H�T��hBU��n;��=Y�'����m�7d�a� K�`�ȓDr�#���I�BX"��ŠCT�Q�'�a~��lH�vEƙ=݈dچ�V=�p>1�)+?	ŋ��
%4|��OӯM��U��CH�<��(�j|�@�@������MLA�<���
<al�B̝�s���#�u�<���_�h�I��&#^������H�m�������̔;`�2�_�5Dl�9�'���y� Ńo��Q�/�db���N	��d/�O�q�	���ߠ�HY��Z��P��_�O�Y��"m�(�������'��TCSc��!�P���t��I�����'ڱO0� 4�?��\�"��-�L�O�('��D�a����ژKB�]�d�O���I����E�(p�`���	���3ʓ@K� 2��S8<���)g+�,��>X��&�3�J�`砚�lytl��.HbDӴ��=U��={�G�g�-�ȓ�dh!�*��7��	+��R�|����q��U��MF�t���ˀ#�:���H��2$�1x�H\;C.Z!@�(9Dy2�'4���F�-t��mf�	9�jԙ�'�81P��.cr���.Q�.$���'2��2���v��X���XvD��naxacn��-�tl�r��B���ȓo˪�X��f�$P@GP�-p�-��E[ԐʠlE6
vأ�@��'Nb����p��$�P��~��K�~��h�ȓ�N��6lN5T�ɒv�ʷ'�ȓ RFY��n��U�p���@�+]S6��ȓ2���훸I:���LԪL���ȓt��!��1h,.*��'* �ȓb��"��'=|<�eEP�u�^�ȓ3�(����~6���0�ȓJ�D�! ��x<2���;>ȓ-�D�yҡ^-}�r B��C읇�h�S�
;t ���c�L�7i���?<� �l�oB y)E�+Ch��ȓr;�<��G�c��D)%� q��=�ȓ"�r@	�H�F���-_=|�
��'+P���g�(D��"�u9Z���'��U�ߑSo��O�rRʵ��'5��TjQ�Q���Ȣ�}��1��'�p�yR)M�;2 +S+׺|�i�'&
�K�-"(ՉC�RB��L��'�p�ٲ�T,P>�I�2��@ЦA��'k�%�������ȴ>����'�$��g���Mz�kݮH�^$"�'���0G	!tV��<1��@��'�2��c@�g�DE��52/2!�'r�mhcRk$�R�4|��S
�'�`���C��{�P�*��u.]	��� VE���	0S����$�=@���"O�HZ2N��#d�+C��r:J���"O��Ӡ�(1�QZ�kޱ>7:�s"O:Ya��G�"���k�!N���"Oڱ�7��
�Д����Q
X����'X��'���'�B�'���'r�'C�Ը��խ^<�b�Ӹ��,���'���'���'���'��'��'�,�e�úB�g����Pi��'r�'���'���'���'���'N\@0&��x���Wd��!�'S��'��'��'�B�'<��'tѦ�M����W��Vq���'�R�'���'�B�'���'U��'�T0�Ν�'O����)�s&f@��'���'���'���'0��'h��'�,�C%%��Z*�@�&��>����e�'\r�'�R�'���'xR�'���'V\�Z���Mu����+ɽ?����'P��'���'	2�':��'ZR�'2	P�I +ྤ�P�j7Hhg�'g��'�"�'�"�'2�'=��'ip\���dz����\�I�N���'�r�'�r�'���'lr�'�r�'�ڵ	7�]/C���3�	��'��@Ȁ�'��'���'���'���'�"�'� �	"��YC�j�˴0��LY��'���'B��'^��'U��'�2�'�ҝ�D�Ūt暑����T��AX��'���'���'���'X�bӒ���OR�	�nJ�?��!%EE�s�������]y��'�)�3?���io\��/�y�XTq�ƹ,GnQ��ŕ����ئ�?�g?y�4o��d�K݄@) t8���n��idB��a����������!��~r�L�C���{n��fH�h��P��?a,O�}�+	9mΙy!S�
ō�-����B'��'x��lz�a�EG�8w~9����<�-��&�?�۴�y�R��� ����i�
�I1:�����چ��Ø��	�y9�x@�͂X�-E{�O��čt=�L�%/��9��̲�y�S�d&�x��4	��)�<y��Ap�B�/<s��)��Mn�O`1�'@ҿi��ġ>)�ʛ#PB����4[�2I�G�e~b�jlt�bƏ��O9l ����ɡek^<� ��!fʢ9 ����*�'��I�"~Γm�2}x�.$d�a���J4;6f��&Û��B!��D���5�?�'f-Z� 7X?�l�:�b�6'� ���?y�4�?���D��Mk�O���m#Kg������0Ҧ��sŅ/z�r���.��X0R�Op��|b���?9��?��L/��Bd �:xj.�!�#ںqà�.O�m��ޅ�'�b��4�'�Phqa@�K�VM��L�r���a��>���i0H6�Y�%>����?{Q���}<�;���!�~�8�JY�:P�X��ny��بqE�@� ��ذ'��'����$���u#Q@ńR/a�`�']R�'G�����P���4/��t��S�"��B
��)���� TT 8��>���
i}Fw��,mZ��M[�&�)�|�S,�����m&�q!�4�yR�'�:@+g�HV���R�����5f�\[��t+i��ͩ��Q��y��'��'Y��'��IR< 8�!y���x�m��FߢJ �d�ON��_̦�Y��i>�����M�O>������{O�6,P6��)W�;�^�`��4ݛ��O��up��i���O��k0ƜA�`	��L)��A�CޢcBT8F	�Yf�OV��?q��?��[p$Z&,W�C�]� � �
�Z�0��?�+OnXn�8�
��	ܟx��E�$!�0Oe�t��AI�Q�V� �ϰ����G}"�gӤ)mڙ�?�H|��'q�x1pG�Zh7|L�'� !jT����V�l�*�5����d��*d�"�t��H>a���C�\5�pJW�$�z�Tʋ�?����?����?�|R(OL�S{���S%	æ`�8�xF�7 �t%��O2���ߦ=�?��R�X��4fu��K�?h�ѣD_dU&lKb�ib7M]��7Mg�0�	�X��=+�*$z�t�'JTyP	O�Hq��kfNJ�B�ԕcg	�1���*�ڿh�4�D�X2 E�0�"J�\Y�-+�MM�^Фu��e�%yiP�ϞW1��dˑ y-�qP��#tּ��"J�F�p�0�aM:�mQ�%��I
�H�|R���!��="���)>[�L�L���ū3
�&\���B���19�]q N[�$���b4��#"c�3�O�	��e���tfK�L��y�pA/�"�@��g��Ѭ�:W��bݪ`�C���`:6�PN��e� ���,�6�X��54 �m�AmJ�S#Ќ2�K����<kUh[>�M;��?������x2�'���$jϗB~���-]}�@�!�~�<��t�i>���ϟ@�	����Cg�]�t�4
izTYW����M���?���XA�-� �x�'1��'�v�K§�8�����ٟi�"���:��1��b���	�x�I���[��΂a��xBF��|99�O^)Q��O�D�<q���w+&<k‍�~T�!�D�×wf��HU�$i���]�@��?)��?q/OR�JV��M�T��BG�7.�ui'Ð�'��$������'���'4(ꃋ��ⵈ��V���VSmܓ�?���?�(O�
7���|
W�ݗE-L��5��<z�d��͉M�I�$���' j�x�O�It�ςR%ʕ�`�I�UZ�pR����՟���ӟ �IVc�x���(�ɢs���ϓl�h	R��۲yf��M[�����?Q�S>�SKH��	fd"&���t^��+��ϔe��7M�O\��<��B�G�OJr�OFXar�E���@�
\� �x(�R�"�$�<iEG�_���� �Y*5���[� L�V;x顢�i�b�'w�p`q�'�'�2�O���5����}޼t�@l�Y�dh�`h1�M���?������<�~�+�>}���jF�v�̀S&���1��5�M����?���0�x�'R�sv`CG椓��/E��%�Ddh�J}��)§�?q��B�T���ξgu�4z�އR7�6�'{��'��ىp[���O�r�O�3���0!&�u��f!	�z<���F�Ѽ]Z6����'^b�'�>��dl�K�И���|��0�cdyӚ��(�p�f�j�d�O����O ��OL�$�8`� ���Q�>F���O���ɟ#���Ο8�I����I̟�O��s�߸v�q��'�u�N����S6�7��O���O����tW�x��9�"�+X��V�P��I�#-J9!,�ȗ'\��'�2�'=!Q�U�7M] Y$2�J��ɑ>� ��ى<	�m�۟�I��p��ß@�'�2�2��t�V�j�fLj�A{���F��W�7-�O����O����O@��ư*8&	mZ��<�	��֘����:�����^X�t\�޴�?����?1.O��@7T���O*�	,<5�B�W9I���a��7-�O����O��DU�z�unZɟt����O�@�aF �|��Q��&�T�v}޴�?�*O��D���I�O���|n<�T�+��d(�cS�Q�q�L7��O����1Ob�4nZ��	ݟ����?��	XZՒ���<+V�!WD�
죯O���@[����Oh��|"H?��A�}?�hb̞�(E�iҒ�|Ӏ�G���I��ӟH�	�?1������	���P�؇q�� �.�s�x�s�O��M3�"�
�?���?Q����|�I~b��� I`��Womԡ���
�8�HŰib�' 9Q6-�O@���O��$�O�.ս+��`-�.d��[��J>���U�ܬ ;�Q�4O�S�?���ڟX�]�� �(΀qw�X3��ȓK��n���i�)O��M3��?I��?�T]?���2m�2N�2((&I;��I�Vr n�R�8��o��'��4�'�B�'Ү�-p�z�8���99�(EU�(�<s��g�����O����O���O0�	񟄮�
��05��(>`�KԈ	��ez�'p��'�R�'��'=�͖C�7�P��򇌌}r|�F��!��o�	֟��	��'YbiZ��4�}�P�*A.(F��B�s��7��OP�$�O��$�O���`^\=lȟD��9ۺ���o=���S�kn�E�4�?A��?1(O���X81��I }��S3v;���6*.!�V�+��:�M���?���?)�L��v�'���'��ԍݖk���e��*ZH1g�	Ol27M�O^˓�?Q e�|JM>��EӱK�/m�|���n����c�t���OJ��%-�զ)�I��I�?����QgKK�Y��`pW��Kn�K�(���$�O���A�O���<�'��'����k�R>��S��27J��� n�������P�S�?����d�I�h,$�9D�T�V� ����C�L����ش�@�c���Q�i��-�I���T��,� D�6
�3�^�*7���!�	���.=���(ش�?����?���?��V�&U$�Е-�xx!����k�i�bX���c�r���?�����m��aY��a��+rڡ:��G��M{�H�|�@�i�r�'��'��'�~b�O�U�x��͝NԘ 3�%��M3FE+E�hUΓ�?Q������?���?iRF�v�ja\���Rl��1M�)���i-R�'I"�'��'��d�O��eٰ�H����Σ6cPÃ�C�&b��O��D�O�Ľ|��&�򙣧�iʆ�pT�B|���!�O�t`aٴq�$���O&���O����<���L&*�Χu�����4z�LX�u獑9;z�röi���'�R�'o��'�x�&�n�����O*E3`��h�đc& C�oP{ �J�I����`��uy2�'ļ�9�O�B�'�!�E W��}�2��:>��mː��-'b�'�b�'��� �Nr���$�OZ�d��(Db��� �1z$f�K�:qK�
�̦}��]y��'銄ИOrɧ�ܴ:lD�C�@uC��	c�j�l�Ay"�A�J6�H���'���$?Q�lMkI�liD�	�8Y�XP�G�ꦩ�'b�Q����i�M���p�Kd6�!qO��8s���Sz7M�OJ�d�O|�i�o�	ܟ�*5�L>�\0�(_� 8��h�C��M[��T���:�Ęhp��FZ��B�c���S��nşL��ȟd�����?	��~�*�}a���G��;h�ęa�ˆ��'=:{�y��'xR�'�M�#�#��I��"W(�M���k���dĀ+���&����� '��X�I���P�B�2>�r�!`�Q����S�l�<���?1�����\�6Hhp��"N}�R�s�H%�oZD�Iퟐ��|�	my�����C4�H�( 8���A*n#V���yb�'6��'��6o,�-C�O�| #1�#�`)qU@�=z�\|ӫO��D�O��O�ʓ��U�' h����D�BEĤ�5`�p�O���O��ħ<A�%ǫ\��O:6�XvmYQ_�� Pk�(W>L�$iyӮ��/�d�<��$�L�5��[7n�/k���最7�x�n���\�ICy≏�+����D���[�T�P=���)��:�`�#h�	lyn�)�O�S$e��٧	Q-�x�e�LR�7-�<	 h[�Ad��~z���Zr����WH��K�NUQÏ���; al��u��EDx��d�:�5��\:_�!�NR�M[�N�<0z���'@��'O��*/��O��`7�1fG\(�7��r"/�@Sd6�K�T6�"|���<�� :T���&�Q��K���L�f�i5��'��	�nJb�t��N}�@��9r�L˪L�sqN�\���<����?Q��}c�H
�ARD=��
e�SN(ta�i$���PiJO@���O��Ok��7�����V�[�2Y��b޼v���3z��b�$������	\y��\͙���c �/��8��
΂�-�d�O:�d'�D�<�"��R���g��ĸb��99.�0�y��'|��'��	�\ E��O�Z��e]�g���H�	([jJ��L<������d�+g���	Ђ�zW%[84�&P-�4�Bǯ>A��?�����$Ɯ3f�@$>E��Z�Qt�\s�Lߕ��| ����M������DҌ ��O��* 7_�V�5�� ?J@U�iI��'��I�7�d�L|
���*!h��|"l�&͢��ʣ=��')�I-�#<�O�����Z�a�8���[�F�F��4��䖅$��8nڱ����O���Wc~�LAL/�,Nl�2��8�M�*OH��)��0.�������x0{(݅D��6ٙ���mZ���ퟰ����'���`��Ci$^��eB�>4~�i`Ӵ\З�i>���������|���Ơ�u��D��427͗��M���?���4L��RC�xB�'���'�2,�S"�\�b����1T����+�ɕ%H�e$�L�	ş �	�l�&p���[�]�Щ�*#4��Kڴ�?aԨ۰o�']��'��Z���s���*H,(H����H���Ѫai��?���?1��?Y-��y��ߵ&DRM9![�[f��(�o �*�`P'������@�	jy�W�dz�B))_0�Z��lf���ц}k0�&�|�	ϟ��	kyR�W;C��7��T���'�0���LL� �J,4�x2�'!"X�|�'ff<���xX�匱[�2��`���=p��r[���IԟH�IWy2M�4�j�P}�&�ĕi�ʨb��K�QV�i11�YϦ��IQ�	syr�Z ��'�
�� �1��s"AH�2��i0�4�?�����$+GS�%>��I�?�
Ү�ׄ\&��Pf������ē��K"���'soօ��-��\����&'N(hn�zy� �;D67M�f���'���3?�`�Z1���rdJ�����e���U�'��`���Ɋ'e8�l[���s�.8�d� ^{��Hҽj{�6��OL��O��i�Z�I�aAG�n��H��J��HUH�9�M{��d�����$I�Dc�		6D�s\M��mʶf�(lꟌ���܊s	M��ē�?����~��԰&e�*�L4B0�4�ϐ��'<���y�'jb�'8�$�S2����Sr���@k~�,���L�%�L��՟H'�֘�Jd╺3����P�M�z�M{�m�<!��?�����t�� bEŅ{�M��&Yl��'�K�	��Ij�IsybLܲ'.V\æ	�	n|�`:���t'<�"�y�'j��'��I�}f�=�O�8�W��H��u���Ê\4P�H<�������3y~�I��\�ʡ�
�p��<�G&�j��듥?	���?�/O����.Z��!Wt������h�<�C"Z�s�>�4�?AI>),Oz�c�$�-"�fA���A�&�6�>�!�iZ��'��	�r��L|b��"S)I�X�*�z�V%�Ё���V��'+�	
m��#<�O�����\?rmZ�Ɗ+!�ʐP۴����uXmZ����Ot�ɘP~��=Mh�z2���yA-���M�/O���3�)���M�.�B, �4@ 7��)6-ֺ�`�l������T����'�.Lyը�"{|�ɧ;u�P���~�P�@�)�'�?	�(Ռm ؠժJ�`x$Χ+��'���'&<Ջ��=�D�OL�䷟[ �'� �y��&Yɴ�)�D7�ɝM�<c�(�	ڟl�ɤ6������L7��L[�@��2�4�?I�MֲD�'���'�ɧ5&-Z2�$�Ӗ�6\�6����0����,:;1Of�D�O���<��i0V�̖�3��er���L�A�x��'���|�V�P�r�M�_��@�أmFbX�3�����b������4�ITy"ː�&x��3!Ĵ��&��f��Y�	�=�vꓶ?i������X)5�I!`�V�9���,n�*�+�dj��?���?)+O��xrem⓭U
��j���x5]�ÅQ��M���������OI��'ؓ)���8f��"Nu�I�iP��'��q8y�K|�����Ǟ]��98R/
x&Ե� �A��'��ɢk�V"<�O�N�A�9��M�`A�w�ظRߴ���1�o� ����O`�)�{~����>��<�3oűV���6Ñ��M{-O.-�v�)�����9��Cw*���n3��7��tI�xlZ֟��	㟀�Ӭ���?�[�\��lP"a������l [k���N;�O>��I)F[��1'�`�l|����b)J��ݴ�?)��?��*h��'���'���_��t�L.���{u�Z�:c�x0#2�������X��֤)�p�
�/؊P=.�����M��, =�&�x"�'Q"�'��i�US�@]�s%�`�ԃ,�	x�����<����?y�����Z�? ���e%7A�Z��䉁�H�Х1v�F#U�OL��*��<���9\����C�ڬ���3�~�<����?)����
z���'H�seاz��e�6π7�^M&�x�IE�py�$���XJݰ��I�-Q&:�#����������ܟȔ'n���$�IR7I�(�:�(��o���X����pnZ���'���	���ak�ܟ�O�ٵI4*�,0 m������i���'�剼.k�L�L|
��Z�)�):�9��e��O�����C�{Ɖ'�b�'M`��W�|B�~"$D#'W�I��I�[�$p�VC�򦁔'���w�{Ӝ(�O���O/���d��WN��)C0�#�3=�R]n��L��!D`���j�)��I��IP-/X���PU	 Kr
7�IJ$8�m��P��ܟd����'�����C��zpKѮ�C�@Q�jl�ީ8w��OؓOz�?���]�Z,r�ޔp�Yڷ�ַPp�x(ڴ�?���?YP��sF�'���'���b���Ȕ�Ǒh��DZ�"U�$K�֔|���yʟ����O�Di�^�H��'W78��N�<6���4�?Y�#��`��OT�:���TLbd3(Ե	�)�T����V����🸖'���'��Z���c����*����,m@���!����I<���?9M>����?i�!O�K�8�b�\B{dh���4JdΓ���O���O�ʓ\]���4�*i��"�3YJ�#�G�$O��]$U�8�I��8&�<�	��x�s@���b�BC�e}r����T�l%���*�>����O.���O��/Aޡ
����i�o���p%�~��d��_�J6M�O��O �d�O-J>O~�'�l%��J͉_) �(ӂ��v.��ش�?������S� �B|&>����?e�LС,��9 e��[	�aM��ē�?��~(3���S��.I-:Dfq�aON\���7l��M�-O�U(������ʯ���d쟬��'�����
�h���g�ܒ�Z�4�?����I����䓲�O8�4��iW�Nͼ š�3~���۴ss>���i���'.��Oc:c�(�[$5�Tp�̯M�D��W�3�M�����?�M>�����'�� B��L�#6�[C��h�t¨n��D�O���;N��%��I័� ����Zg�����Q�F�mZU��}���)���?Y��+�`�1�����I�J&mbr�i��
�F0O���O�OklVe�������|�n�q� �4P�	0o"���	sy��'���'��1q��,Sw���zT!S�W� �<mc��Ȍ���?������?���*J.`(E`D�t:�訥��#]D쪄-�����?���?A/OlM!U���|����t��[ǮE:�Qg�W�	ɟ0$���Iɟd*����XS#�ن#�t=���FeL .l��)��3R����� �H�/�P����
�*��� �,�(3cM4:��P�BJ6Z�:Q��b���\{TA!s؞ y"�3���S
#"��'����ܙE�\8Y�lN?>��|�1�����DH����D�2h�*G�5��ݾn}9h�KԘ#���u�\�WI�]�᜞\ά}ؑX2c�$�r�ҠR�)%�ق�ԕS��W�{��	�H�>+�2��$O�$?��N�Y��@K�JM#u�|�[0Ɗ6a�NxF/ͥ��	Ԉ�O�$�O�4c�'\�,D�;�燔+2��r��#?,��B�Ǩ.����D�{�d���8*�����n֭ZT�8���\0���OXxif���ㄾ7��Q��L�H� ��%a;J�0��w�|m��G�a9���MT(y��IW6*%�'���?�E�� ��ԆQ�&ˀ&Ώyªب��?QL>!��D�>I�䙙t3v��!�v8	a'��L�'�6mNӦ��I��M�(�P�IY�;z<*4�P�p5V�X����) ��D�O(%�]. ���O����OH����?��'���"�I�"��JF�.�F���'`Bb1I\"#d@��	AF{2��q��w�z� چ$͗G-N�d��C~��F� �I-�0��hO�$c�&W<s7�]X
[�1g:�3r�O앻��'����kyr(� jz�4h�+7Z���q�#�y"iթ/{"5�v��>KEHU���Lm�"=�'�?y.O�x����ap�.֓]@�K�dM�I4=@R�\Ɵl���D��$8N�I�Iԟl�'%&�݃4��a3��0?�
T��$ʳ|�ɛ��E�s����*���O|-giZ��� �b:�B �o�U�c�
N$�B%�[Aܢ?Ai�̟\�شw^�9!�
x�|�k7�_�<ѐ���p��7_�,�. 2���>;`M�ȓcz��#�,˛Ptd��_gz�Γ}3��|�'�-P�d6M�OV�D�|RR-KX�6�Z�B
7d�Y�(k�dP����?A�Y�0�Վ�j�v�#��G-cz*�����	S���"��͞Znm��	�l����C�.ECv G�S�bqL�X�M�/~F)��V�<YAaU���S��)/%�2h�q�Y�=�h�*u�@�!��,jΗ�\d�S�_�'-~��M �'8H0ĕ"]a����ҏr���c�'�����m���D�Oʧ.+�D����?��y��#�Ð1?�lEa��\]��y��РuUԙ� ˒Rxm�tiS>4aR���b>���FpX�FSE;��.Mpvm���b��zTቐm�(�da@��K�&{����0cLv肪�#H#n�"D��3��'Fn6�YmyJ~��'��� �u�6E>|�b�cQ�]�mW�` "O��#�/�@�����7S�,��!�HO�n��S`-�=Rx��ID��'hHB��0�IZK4|��&G��d���T�ɠ�u��'�rG�1eX�l�#��i�R��&5 �X�3�6� `l��a+p�	��\��Iʄ"��X�+�o�b�̓3�|�)��	�/�����U�'`t���ͱog�R����6���'j�}�z�a{�a �Ph�|�S��J��P*ࠑ��y�f��͡��I�.���*��-�H#=ͧ��XRQ���iƊQ�VkE�h�t��EC"Pn� r�'�r�'H���$��'�����'BR�Ф@)2�L-�bU�I�5�	�v����'�p��P�j*�ɇ��G�.�����	<�M�a�]�R�Q�_`� E�s�<i�+��iي�0�ȅ8t���o�<Ie!T;8�)7⊊G�.���V�<Yv�i��'k��t�x���$�O8�'H:�k�u�~	�3(Z%��b��n!��?�ߦ�3��V�Q6��#��T>��I3'5�0�Ǻ@H��"�6ʓ]�i�rM.P�����	�@<r\$؇b�<�b��������섾Q�1��!!ʓ<,��'�H�:l��쎈]��B�5�*�� "OB��#^���pQ�����'ߎO>���&�@& NK�A�
պ�<OTx��A�A�	��O�p�`�'���'d�`����^Z�tЧ&�u��:F���(x��T>#<�f�%J�vX��I�(��<vO
�la��'jC")R����o?E��e6�q� �-|�~-��de1�q����ɧ��R*»Uk�c �B��Q���6�y2-�;1���g"���xti�&K��O*�Fz�O�2�	��ة�Q�f��Aϓm���'� i�'GQ����'�2�'�dם���)i�K����tI�O�rh���a��X6��1h��1 X�r��q7�l��yR��Bg���V�fQ���@	�tBR�!��8�Q�P}p�8�O�\9ark_{̓A��H�6JL5v6�� U�H���Rf���ɀ��=9�d[��J�D���z#�_}�<��'�2LE�����K�T��YE�u����Sf��x�!��4#f�k�ʀ�=��h�� &n��:���?����?�fB/�?�����fZV�Dc!�W97#Ԁ��n�(�DU�1�>��8!d �,��yB%-��b��l,��p+X�A��	�F�Xz ��ư8���BԆ`ںP��&Y)
�'ݲP���?����]6��`"ٷE} 9P�f�J�<1����y��0��6y�`dXB�<���� ǀ��BI>B��L�O�<�i��'t�'.gӖ���O�ʧZ�t�ۄc\�@Q��#m�2YI�,J=�?���?QvϞ�&�~T��e_�i��`!���i(&z�aE���	�
M�@�
�]TQ�<����T`��9����Ћ�|26��!|G<�*ӎ 8<���	�KW�'�lq��7F�>�����+��d�ۢ*�F4D�$�`��k�P�Z��9/�=!!�'�OZ5&�����j���Ǐ�+�-Q��e�8I0����D�O��'l,����?����~%`�^X�Ё��2Gݤ�A�Ū)1�
(����&�,.��Sl����J���9ޔ�@t�ʤQ[p��r�C,=cvPR�/C�s�fL�V��@+���w �H�"Hq�M ��	�0! `O�h�'���'?�D�r�� :#c��]�1j&M���O���䜃l�3��8W�h��	�RG��Z��D����9O��-;��#�I��(]��N�D�O�͐J��(����O�d�O,M���?���pώ(���.$9�5ʥ$�!+�\�o�����	�Fi���?�A*G�N<���b�`��ğ%N�%��a�>(�Ȉ���?���,�2d&lO�K��Me[�F�
#.hmk�"O~%;��ܘ��|ڠ�33��lY� �M���d�|&��7-Yi�m�F��5*��R�+$b@�D�O��d�O��z%`�O���b>�+2-�OT�$ڀD+�P{@�]	n {����|��5��d�k�0�#��5G$�pʜ��|��)�?ɣ�i��i[��V�[�~��t�HI�0�'�h�9aGX�^B6SU�ڨ4M��8�'Y�iP�㏅dR5A�Z6*�N��'� 7�,��߁[�n�۟,�	l�DĂ�^+��`dɓ���9�#�=.�\���'J��'.d���EHN6HX�CE�%�xl�|�	A����Ɉ'��p�B��W�'c6����v��Z����8�O\��k�fU�8�)0�~x����!XR�#�'6��D飌Ũ_�T�"IǸI�x���S�? �b�뇣I:�銧��!6��9y&�'R�O�BF�S��4I��Ǭj���ɱ:O\��������Iҟ`�O���p�'|2�'H�(��/V��z��ڔ[�l 
��G�t�04c��T>#<1ed��>:�35�@r�B����
�F��O?�D�X'�Ԛ�g�$�Ӕ���.gt��u"�Oެ%�"~��5.�ђ.H�1��	X3%�3�B�	+<]��� i��\C���"�#<)��i>�I�Y�3J S�2�� D�8����I��� D�I�)>H���d��ΟĪXw�w�ɸ!ܸ#l��u��zi��Ú_Zn�&NČo���p ϝ;xO���)FC�غF��Ȼ/���c6M�c��Ѩ��V�)�Bl�aO�fޔ��֌��:��Ͱa۟b���X�ј'���sd�,?���9�U�*���'�l�i��g�a{®[�2����됌+BM �H1�y�f�\:@�K�F�"^=`H��BT�c�8#=ͧ��l�0Q�#�i+��iB%�w�
��P�R�8����'cr�'�����i!��'��i���'�Z ����&(�0��O��l���0�'Dz�@�.��A��A�(W$ǖ]��_E��I/�MkB�D-IpB���H³~�����~�<�Ԅ��6I�4*�/n����lw�<1u���4��t�����<�JD����<�Ĵi�'t$1��i�,���O\˧_͂��ֲ{��pQ'��3 ���AN���?���?���$.�н���+m�z�Γ��镥R�H`�U�O6Ƞb��.g�Q��e�Q�a�������9X�R���T���c��[�Ҍՙ�I�� ����Y6�r#<���󟸰۴WG��'��S ":$ ���5oR��ϟ7I-�1mڇ������9Oz+W)@�th�M�к�	ϟ(�'L�6-����	�u���B;���
��;�D�I�m���;0�N�IF���><���'\I�ksN�vM�'H�t�*�(�S���u�'�1O�3r���p�#�^��,j$d��O��)o��O?�� �j4��-v{�`aS��� m�q��Oxc�"~�ɦ1#���+Y+WR�d���>��B�I�/Ј12�)K
v��A��0;�"<���i>q�	�\��$����,8�(��
O1x!h���ǟ�J���4�-�I����	�X�����cN���	�XT��Ax�ɮWB��I���f9O0�Ⱥ�tБfڲ"8��rRf��Pj0� �� ����U2�)b�pI2�5�$R!h��Ф�4 86��r%��n� ��W+MT�dN����t�'o�P�$�#���rģGD�-����s�9���<���$]�2���T��p��GX/dΛ�a|Ӧ�ORdi����s��0Z���MQSn_-X&�bw�O!X�4p�Qj�O@���O���9)���D�Oh擰o�đ��U%��iJ��L6,��Iᴄ��Ԑ���=t� �Za�O�'I��bagR�c���s6l�O)�����W�C3P(k"k�W��8Ad�5n6џ�`�,�O�n�+Cv Y� xS�ܐ��T�V:�B�	�u��D	 O�/޼�����;�C�I�/3��JD�t�R%�g*��dW��	��McH>����9l<�f�'Z�_>-:����T0r����H��0aKׅo$��I۟t�	�0٬���$Ŗg�0���Ȝ�?�O�$��5��]F�rc�������D��y�$y��i��{'ʉ蒅!'�哋5�Bب'N�R��X�&dL0�<y��ʟ�G��~�X����������ѿ�y2DI0&��iJ� �?�r����0>�c�x���<���f@�(���CH���y���6B&6M�O��$�|Ҥ��?q���?�L*(X҆�wجQ��G���"��8S�K�
r	����L��!���w�&ݫ�(�V̖a0,˞n�����la4�g�p\p"z�x��D�*4�q�wU/P��`Gɓ>�0\ Q�
w�^�RA�'�1O?�D@�I���9f�G?EthA: B��	�!�$Jw�^q�1B�):c��P�@������4����(UZ�k�@1>��2u㚪f�^�$�O��)��]�f:����O(���O�Ԯ��?�;L�̈�V�9IbҬhWk��'��@�Gه���v�|0��AF8k (:@�.U���I%;^
��B�^ɸ���
�(.�bC�@�l��D��V4��8lO(��"�_�Z>$�(��1`^*$"O�E�qN�.	�|h(��S�n�ĉ�3G�[���4�|R	�.� 7�CX�H�"��|b�uKC.ˢF�z���O��d�O��27��Ox��s>i2�(�On��;+X ��7��d_����.�),�|��Π���>��Ձ��|W�|#�G3T��|�L4�?�iKt�C�	�(+]��o
�fY�mj�'&8d�w%A74 ��O(唨*��� Ω@�@�%Ix� S��6qbؤ�E7O
��>ap��h���'<bW>� WA�%f��ꢎE�!��@��/n�
��I蟄�	0Zvh`��l�S�D*�)�BJ�c_�%�*9p��Ϯ�(OrP��2j�,`��H�,2�v����p探<9'��D�D�� )�[1��HjQ	�e���y� � i3ɱ�͂�A��������I	��9(��WjU#fWBɉ�ʄ�&�|�D�t �fU�L��H��B�?���'X�/.�h�3��+�Tq��^���}s�� S&<����X�-Q&�T>%�|���0@�-�El�-){����͂b��ɐ1�9o�va����/��؁U̒	4>�Fݰ	r�Ͽ��G�s�(�PFKȑ�^�C1�N�@n|�2�C��V��<%?}�SOy"���b����"� ����&��yˤK0�C�Oݫ��֡��OĉDz��}�����i4
5��L�-b\ЋdR�vN���O��c�W}�0���O��$�Odԯ;�?��iuNl��b�6^�TL��K@"�ϓzdT��f,Ͼz����	�p�HӐˌ>jhzG`�>XƄ9䎏.���k0�Ǩj��&J�?%����MF�b#ɳ<y��A�9:F�{��Փ(d(�%k?�埄J�4K�'���'��	)��Ɉ�l�?0������yI��	R������UB#d;<���V�� �HCٴLl��'V�7��O����L˧CڔAf�i3,9(%!��MY�l͚'���:"�'#��'�RF�4%9��'�����EߘR�|��P���,*�i��c��|x�a
�+���M!�|0���	;rpqP�F���[,��<�BA>��X�7�ݚP�Z%X�hE���'��p��?y��M�>�ەս:e���G�<�J܏b�2�b�GH��\�©�F�<�$bV���ms@Ͻ+;�Q�Ц]�<�f�i��'~jlQ��f�R���O�'%7��2��ݻk�vx�a-� 3:�UpTE.�?���?���RG0��rs	л]��x����I�	K�Tb`��B�B���AJ}
Q�HؤG[�3k�c!��R��ea���ȺCuj�r�<pj�+�,s�i�ƘH�<u����{�w��)�����'?M�	�d�n�3A� f�4UыI�|������S��y�#��\jTe�'CT�IU��9Rˈ��0>Q�x�LL��d���g��6�<h$��*�y�
ý)`�6��OT�Ŀ|7'��?A���?��bS�R�`��C�k�x!��FF�k�e�NH#8c
� �i��T>A�|�	�Xbz��҂N&;�d v�j�ѱ� �!(Y�8a��[S��gՆazA��@�I&�Ͽcs��u����R�M�>�� O^-6��q�-4ɧ��$_�7���a��-�>yI�M��yR�Zh�<����G�#;H�YWn��O4PGz�OdbM-��3�`�'��e�ׂY�"�'��,�R!�~,��'���'����ɟ�]�L4�+��Π{L$cV��35 2��q�6��w�	�Ty�9s�tF{R&Ϗ@�|1BG��b�0!��< e hi�,�!Br���&)[PIty"�O����)s�6L�'8����+�-U�z��H�S� y��'6f���:Fa{��^���0���+>8��ᄭպ�y	��@[r�Gj���b��"=�'��=�ѿi��p��$�� Q��7�jѨ��'bb�'�����'��IOZ=�#�C�Q��xw	���	�J nb�����A�n���;+
bؚ�HS�Q�:��w�D�-BX5sR��;L4V�� �#Cπ�Ca�ٯ��G�=���O��'��7��.ExMI�k�C�>%��MΧ1v!�d�^������[	 B����ʙ�\~!�t�T�A&�ߚN���0�)��d���'�쫔�\��M����?�/�.i`&Ό#ւ�8��4P9֕�n��#m��d�OH�d�f��6-��#"�@�	�?�Oa��XՇP:mZ����0	��P��Ds����]�hH-$Ps�p꒎�/�Q+D�ףK���G-�O�jX�7jթx��'�D�7��O�G��b�iq<�;u+��Z�>�#'�ڵ�y�h�!;+Z�9�Z����"�� �0>ɢ�x�E@i���ٳ!D�
��,G���y�18 �i�"�'�ӡ"0���ϟ��	HN���+K�����iǞ�����݉?F9w��9����S����'�R��A���I��E9�oEM~X���M�+8h�w��c��ĀSB�`�PCB�{�r�0��|�:fg�0y�"&z��0�ݱ:tH�[6�ҟhJ>E���8myAV$8*)U�4l��E��AX�`���z\�Pᯝ;$�<XFxr�,��|�3BD:Eh��+/_����/�!�?�`�
��f�ո�?a���?��!^��O�N�+�eR�sf0��ϖ�^
�������`:梏�8����Пў|H�Z䍢AjT�c��]@��E��D�S�#�r��_$���<=��Ѱ��(Y��ɣ������wО���+����'ި�dm؞$��Cލk?��FD�1�$)�Fh:D�l�bM��wa��e���HO�/�D�8"�]m:� F�is�Q/�&�� ��)�.�s��O��d�O��dU�jD���O���������I�&q�	�P�N�
��<�r�L��$��F�?F��C�'�m�P↓r��L	�&��qg*Yrp)W]BAK@D��e �>D���E�Q]� �{�B�(�?���i��K�䈑C����O�E3
L�� xӚ�| ��9O�9p%�&z$A��i�rj>(H"O,0
C���yڦ���'A%2V.iz@<O�qn���H�'SD��t�qӰ�d�O��'~�\|�s�[���E1�e�;�6	3���?���?1��+�nبB-��%�����O哈Y:��!��Y�u|��ÌFc/��<	��YN�= �e��La|$��i�ZK�A�C�/jQ���cgس$�H��#nE��-�5�'�IRƞ��0�'#��#"�Q�		2�r�D�@]�̆�(Rl��#Уw � S�!�;o��؆�I%�ē8j5u�P$8��Œ��7*�2�I9d$����4�?�����#D�2���O"�ē�%����A=��dS�L����!A��`0�@smH���S����'P���0`|�V��ÑZ�d�3eP3<g�d�oA%/x��lK#u4���E��*J?���*����O��L)vՃ�IF�|v�,Ƞ"�O��'�"~�	�/6(��oԠoD$� ��)SK"C�ɌOǒ �g��?y�*��K�"k��#<���i>��Iyg�И��͈��qjCh4!�^h��۟Ȉqh/�Lt�	şP��ȟ b[w��w~�)�Ǘq��� �\T�
��̦��)N�e��xy�o�:`,��I
"L�B3��(2�Nu1a�"�X���i; ]k�@�! `�[�bWPF{���#=��j�+#"<�b�(� �~�DT3�?q��i��7�5�	�����f�Ҥ���!{�4��*y�!���m0��BCY�^��%Lި#BlFz��>-O���FX٦��eY�s䪕"d�d�r�XT���	ԟx���E�R�����ɓD���:',��||%�0�F3$��PeH-nV��6i</��z�4q��mV+�f�'��;'��,���ʘ���Pbkf��;2�G	}�N�����5�qPU�(`��@��|r�(�?Q�iy����_zL���-Gg�Y�� e���Į<A����'jB�'��}�v�� ���g�R�3�B�(T�':��H�d�:���!`
�H��Z5�y� eӬXnXy��B�P6��O@�d�|�SI��4�h졦�ߪ,a�y�Wn�v�2��?���t�ȜA�
��(���N�"7 F�K�X?���މs�>�c�͟�N>��>�
�2a�c$S�s����[4~~�������肱=��eAF)ר�X)B��I#f
��d�q�OK�}��TN
�I��i)8��)��'T]0�b�!;~����͘�ZD��9�'aT8�#Y�9h���)��W.��i�'g�-�@Gh�,���Oh�'2�4����?	�/!"�Z3M�9K���C��ҩX�as"����%�g�ףd��9�V����2��OH�s"�D� ��&��2]>dXe�T.�����FM�J������ϝU�en�]��*2���k*B��4i���:��%F:幆���?)G�if"�'��Opr�'�B�ұp�^ai����}����>s��'��}�D	D `W`<d)X�b��X%�O��DzJӚ�DR�/�P����B�c��� +!%$���OҀ���{��$�O��$�O����?!��6]x,�3�X�Bj�u2a�3-��5)@#ˉb1� �< �P���)�GF{�Cܹ/.l���M�VK�A;fC�"YR	�����	����Z'SX��
��hO܀y��L�,���Jѳu�J�"!�O X�tk�OD o�쟔�	��IΟL�i�m�u���(�Z��`ɇF��,��7D������"�:M�������*e'
��HOƌn�̟�'��1h������V_�)�B�Y�rjR��u�ޕ�?	���?����8i����?��O-�D�W�(I�Q@U�}��a��Mh|)�K�8I���@ӓ)[f�ҥ�=P���(hU!x��AƮS<o6 c�T�ك@AGS��J�/ ���8Y��O�lڛ(+�	�fC1wᢰ���χ+�C䉂h㚡#D"J"n PA��Q�"9�C�I�>ߚ�[�/),+ Q�u �9Hv��M+M>q����v�'�rS>5���дc��0�� ������AD}�I͟���sA��!CٯY��A16BQ�<�O�����)
x�A �6(�򤃱Y����+4:o8�8`Ϭ�B �ƪP Q�����W+X�n�� �& �)�IL6��'햁��h��Ƣf���|
&g�6��@c���3\� ����N��?���9O�tC�GX�k��h!�Q[IH칆�'r<Ol�A%Α�+��P!��B�w0�@Qq;Oܱ �O�>���O<�'~l�T���?��"��+�b"�<�P%�9E ����L�p+n!b�ţ;;��� ��)%��O���  �
p;�8��چl9��Y`��.8n����aS�#�|��喅>� <��eY�!d��g��w�D�a A;q�uyVI�j�������B�0���O�A&?��A@1-E�5��%�#"OP�J�"^�	��x�k0.���u�I/�HO�)�O���֍L�2��5hD��@���O:�d!i�F�S,�O���O6����S�Ӽ� ��f�Y�T�9�-Ni��Mb"b�([�t�r�� T�:p15��?���c�y��V�p%��,�_g(y��N = l=$�9V�`��V;\��TA�OC<�r�eMt�R���с�;"lᢢb��'ɞ��0P������=���H�n��2�J�%�
uʁ&�v�<�6e�E@F)�@ �<�:`�Wi	������b�~�9��4d)�����U�1$6*g��%��!H���?Y���?��Q�?)����k�>}�֕ T��$U9��!�D��4ـ�i�j��D���QX��C9
J2ͱ��G /��7�%*�l��^�I�|�bD_FêP��eE��'R �����?�7�	#�>y�.�ED��I3�I�<I����x@�͒���x���B�<Ae�M�]r,��%R3�=I���<!Ҹi�ў"|�2��-U��h0����Š���m�<��o�l�D���� Py�l`f.�s�<�@�,� �a�惛�` �eJq�<y�J���A��6#
x�HEv�<�0�P�B���4I�-6�<�Rdn�<	��X13�tE�&���G�z��Ղ�o�<q�9:�£�PU*Dp�+�i�<Q��W�k�$0RN�JVlAC��e�<y�EP?Q
��n�E9�y)`��h�<���RR�ؘ�f��x	�)�c�<���((�~|`�Lܚ-���G�Wa�<Ip�N'+��5��#�)r4�	Wna�<ѱ�P�qt�qkĻz�pi��aw�<yՃ�.!���P�V?E��K�y�<! HP�@J��wA��!N�����`�<���Q������M4+��a2��\�<�G�S�-K����ǭd>A! ��^�<�w�:������'���藭�Y�<���N�C	Z�Sq �=8��0��^R�<��� �Ly/\�2[(�����Q�<�b��$!ҁ���2�L�<	%JV�f����������2fF�<A5�>I[��)�N�1J�t���#�Y�<$
W�y)�	��ΑL	w-@�<q��H�	�@���[�BU����Q�<�@T��p�`�1<<����S�<	��ŭcX`�v�$zih XƂQS�<�V*�nKh��%^o_`��u��N�<Q��:Ju.�ViDz6�	�Q�<au�R#PCcO�� `3�CN�<�k�6Y�^�h�$� \���5�C�<��o¡_�UU�`��U�I7g�b��5J&�q�ܐ�P�	Ky�'Rjct����g�NT�@�M������9U�w�n�P��8�8hx��)�ɖ_���[F�x���;hm�a吰ٰ�c�����=`�[��b�p�a�'$�|���`� AƼ��� �,�V}@���?�p<��*[���"Wf��I�]�u��+J<��S�������r.����h�`VF��\����ʦROjVS<�@�B����1�'�f������(�L�ˤ��#vq|MYT-��轸����xx���>yuII;~����b%��i��"�*]��M��@��9^�R	��KCM���>��@�$�6|'C)3gxpH!FX�I2<��u���-5�U��S$ea�%���J�8�PW&(�O�6	,4H��,�P:����fP�*���C�1|K�H��]��O�Ι�.|�BU�H�''(YC���=�!�$Ձm�`��7���.��AU9Rڊ���?㰸U��/1P�S��w+��A�
�b� +ɇs���{Ò|#٧3C��y��>~h"�2��j�H	���f5~�r�H#?�hAfMj��ᆁ&�|�YG� b�?Q���'*5������ �P�I�+ ��OP�K�#a>y�V��;P��Y	Ƒ>����(2�`I��S�n�(Y�A�!-�� ���0t%��~b��ٶ5�p(�MA�"D%���#I�lY�"�BY��$JD"?J"?�ݍ9�����'VKڀ��d]����}1�Y��`kZӧH�U2���o���!�+�1k&��@E�x�����X94a��5fjɁ0g����ڵ)xj1�	�!�
/O����4I���")yD�S��yr�`��{�2D'��c �8ywfd�"-�(<�V�"&G�<�π dq!CԞzPS$+X/J݆��A7rD@�'=(tf*�f��HR/*
d%�,�D@�9
R�-����8����@���Ԝ�$�ȒyQH��/O�?��J�"5w��:�I�(*��tMK-/4,Pw�Y�S����JN��S�����H����ċ^e���Ќl��A�#	�t���?!�m�D���8�B�׀'�lP�2��j��$�7r?=s�h��h��N���c4��e�P�`0�ש��A� I[y�4'>EJv�b����'�;�.U$ I`p�CD��,�������↏� =��ģ�-"'V��,|~*�>�լ m�~ I��;AX��s�M
A�O�@��~����4@Z�H��*���a��;|+^l3sE�(fTK%4p�����uo�)���V�D��U����ʖ24B�K��M(�L�XA��X(l(A�(��t�؅�e�i�=�Wϟ� ��ȳ����4�N����[cH��M�ĤRqNЧ��$�:�ll`!.��3>�H���CF-�n)f�Ǵ5��1��>�`�d� 5�!v�MX� �h�j�G\�$I�Y0`�� �����P�D�A���H�e�܄�I���D�X "0};���Qjؑe'�jg#�p~r�ĐcKNJ��V�� �cߡs��ԧ�)!:!� �$��r��THU�%���*�`����N��'2�B	(�%���ɖ|�6�����N:PY��O�sg�lˣb�o��,�b��UO�)���Z��f�V�tͳ��5�± kNGz��c�D�K�^)RG$+"0�us��i޹Y�핒 ��8V��8 8d�p�h�(�F���J�˅�Z�o��I�tB�<jPO$T�}�'��F�P8*!Z�P��Ӛk. 1��b�a�'t����-ݼ��`O�9�
_�5"L�IGǙ>�xՂ�E� T``d�'������o� �>%?eZ��ށ4;���헫F:L5�&�HD�O~�h��D�,��ǳP�z��0�<�Oh�JƬP�X�9�WCR�(����g��$L
��Τ��W?eʅm�#9�$O�B��S*��ѻD+��k?��������4#�/|�X��'o�>��䙴!�4�1"%D
0iJ|�)˼��I�AC=c�B���ԗ@�ͅ��ﮄ��Ә�z���H�
JH��7O��Ǣ�E5�f����$�:�rЬ����O�0@���'�ԯ�V�c��;b��D~�M$~����-3�L0��Y*D��1�1�;4�@�V
S� k��i����$J	��s2�)��~r��H. �)��=�l�R7oC�\�i�'� ��fƶ�8	Д�2X� x�!�?j�lj�P(�72�PyK����UY�m���Q �x%�l���|"���
YZ�m,}2OI%>N����=o�@k��ϡG3U�eHÍ�l��u��{6GYE�g?�Jy��yH�m����ㅍ!$횳�7P T���Y�y�^�F}�w�lA�hZ3g�\ҁ�������4Hb�Mj䀙�/� T0���$����� �d$/?)�-,����;-��!�W�E�2p�>�ƉOH��d��}�eh�ȟZ�$3�°>����q�V1<j���>�֍^�x�zO>���xX�^K�|djG\�M����"+s��pP8�#�U,6&���e���,�b��'�X�'Qy:-b
�X�X8�nF\[���ò��ɬF8�=8�O���ᦙ�3l�'�z5�p�E�Q���G�d�+��G#h'��HiH�~�]p�C����O����A�ڗE&5��˻���r�k���|�TlB�L���a
�p<��V�TU���9)�1��)?�Mi�DE�I�ސ������k���,��Y�O���	=�D����PJڬk�*D�5���d�/T�@(k��E�PuV�z�O_�al�ɑ "�!�9�y���N��#�$ةh]��������I���p�'|��r�AK�QG��Q�Y�K�8	$��U�I�KJ8C�W���q�IS_��4JX�N��W_��4��q�Q>J#�t���� :��4h���|$U�c�.�I�N�u�b���܃��]�5b�ы{��)�5���`'ʽ���K�A�{�>@P����?�'J�(,9�@�a�� 
�"T���A�3��Y�N�+A"��S�'�y���dUL}j�@�L��ʠ̇���<����*��I�/!�P53�ևY;0�*sAQ2/�� R��`|��'
ґ{e%P@����]j������&8�-
d&V�=����0/��'�z00��!�������H����o�8�v/!
j�BD�Ӳk�Z��B��� w�`���T:,�R�6�dH-A��y�d�,	P�
�� B?��P���g�&� =\ "��)������d��m�=C���A�bI}@\��^�_��1��K=T�������L]�%��4W`*m����9-�Xi��O�� Wa�--��j��Z�V&�?5Ad
G/�܈�w!��D8&�9�,V3��OzJ�N��KI�%�5�݁$1k��|��͸4(t4N��a�G`����$�l?�u/#��rh.��tܧ.�J}���
�e�����d�Ny�'���B)		OI����-J�+	` qM<�O�.���L� 5���b¯�1O4�!a�R.OHt	R/O<�ʂ�5b§3>e��'e�t8��=V���"F�R��E�P�X�3�z�!A`K��)��ҥU%��'nU
9hAĂ9<pҖM��f��R���V�@-���-Y�5XEe6�Ӽ�u�T5�p�_�J��#�IX?��쐫Pp�uP�-���8-�B���I!�I��gtD�%e�"�Y�`��<km�8��DW���C���>��K9m����߶:��u�1h=#�6؀5bA�(@�l���H���1`�-�������� ��^�t�wF��rsj`����7��<[e���2	_�/E3V��au��S��ONW<Q!B%�&{�6ܺ����ӣ
�k��k�ݦݸ�������c3�� $�JPd�@��8�cdѤ,��1�fKB�D�6�Pĝx�L��'6���E��d��|�d�!%T0СPeS,�LU��j���^PF=J�6����D��0<���j��G� �>xR��v�U�̸#է�:d!�/ō-g^8S��O���]�I�
�b�^#`�2p����0!p������v ���۬>����ȷ&��kH�(����jWF�z��ٰ<��	%��Q�6*�,M��I�d���ɒ�'t��9B��05a��[2���I�!��q)�l�y��X���^r�h���\)��@�i�<7T���-�6"Pʤ���� 6�qG�'^Bi!�	H���Ɂ*��d���ʄxvN�s�jT��f_�=�M�c��Olq�B�8�qG�4�$pDg�&'й�с<}�V(�u�Q"���jv
��Z�8���d����O�nO#j4��G��/~::�2P+�)��5��H�?d��࣫SC5☀��Oy��x#␓� �p�(���
ʰ����$� D׮J:袤�w��zѢ�J/�}����t��x�'c�y����#'�����V��Qx�S�'x��(@�@�4>��B�
dg�l�'�h}����5DH�E� ��<Eɑ�Sܧ.M����L�2�p6v�����l /!�!Ȑ%�͟`aC�L�'Ap�'��b���
d���4�F�e�Ȕk�%�&�ެB�c���?Y��\���O�h%��|2�j pe��"n
�.�q�T�U3*�S��;ab���&���\�>�;`QgU$Y�~���K>]�L� �( �1�PD�!���9��сĴ��?�λ|h��� P<?��m1�Ҏ�xňď6�����E�6�.��d�G�ߑ�����`@Ia��,�@��P4~I��	#���b��G��I[�C ����O$kՔ�S��79="Q����"��/�zE�歇�kĬ��`��2���o:�*Fd�����r�R0ġ
��`@I�y��y+S'u�8u��H�r�' �'s�D��1u�~����T�:#�;�B$��Q����*Ѧި{D�c?���|R�Ĕn�Fxp��ѓ~���ҹ�L�c�'w�<��H=�p<�1\crhʂg��2��P� ��K����1.��l�&(B�N:л�����?�̻Y&>u,Jc���¥T7E���qU��L8���ǣ�]�I��E�j�L}��M�O�� �4E� D U	�٫_�a��i*!(�Z�,H^���� |����&�,_�q
©�%�!"ֆ��Ib��l1FL�M��eP��[�8ҧ��I�N���y �A�������+�����":}2'[.�2��G@�@|�I�'�~�2�fEe������
FN�y��W���SP�9���)�����f�r��l��ؕj�Z˸�j"'G a��pÒ�i��ǊN�C�XQq-��PlheǦ�<QfMՕ "B��I>E�TG)�����wNm� ��x�$G}��	l�r�,�&O ~���;i�h��Y6[�q�v����r �O>�r�ѦTVr���i�6M��X���֝BȺD�.6B-���t12��!Y�l�X4�;��ԸW )�?�j8rvgS}J�Is�k�r���?yF���4�r��ކjz�͑��x��N�"^`b�ς�VL��BC� ��*��f},�i��'Tju�)bQQ�Ս�A���IU���� - %]����I䧿����� �(�ja��)[~�1�FJA�<�����A�=s��gD�*5��8iax"���C��9�$�E�A���3w�Θ�4�Ή-��f�P#��z
�9�X �O�(!'��8g�+r�t���:�H���W#Nr�O��� ��5qgM^�N¾X�U�$��u䦆��Ѐ�E`G>�l�� �+��:D�D����Җ�:��Rvt�*�&[�{�QC�I�% T�!aO׉2���S	$a{­'y�`� Տ�xv�	T
=?\�q��+}���o׽ %ay"� 3w�`���M �&�c�f��Q�d=�O2�ɹ���I�
h�pg� a8LC�M����{QS
H�l�-�"Ot�زKQ7Ֆ��&Zx�I�"O�Q�'���b*��"e�GU���"Oh1H �ËQ���	w�@�L%�"Oа������ �0=ܬ�g"O���G�(�N��R��fv��"O���� %���H­ȡ�"O9��qa�$9���6~�(��"O�%a�94�����.�����"O�ե�4B��PE�Ԓ�����"O�����
��@rB� �&4ѐ"O�y�2�	0���Վ̃N��Qa"O<���h
@���R�L.+
 @c"O���a*ʊ"ޖ{��Nb�lU`�"Ov�DIS�H����S �	�Y#"O�P9T����5b� !��Ȉ�"O��(F��2�9���JL��"Oސ;�D�F`� sw������"O� ��� &�$XƼ*��ڶ>�B@��"O�S	̩-�� �V�$x93"O���@�ޚ*(���� �%s��uj�"O:���I�{%؄i���=*Q�1�'"O\x4 @?#9�-�%^@�Q�"O|����l�ډ�G�ҟ+F yc"O��֋��$���ª8��T:"O����ߴW{5�Pb�)|urT"O�y�cH�9C`|	QaJ�F��$2q"O"�Sf	��?KxD%+C��-`$"O`���kƛU�B�Y'��u�R�&"O�I��R;>�E�d��<�� ��"O��A�x���"$�?ޒxP"Olh��`�;Kʑbc#N��""Ot!q�&R�_P���oR�"�`a�"O����ƐcH�ɓ�hº+�H�Ҡ"O� �%4T������&��L�"OAQ��X�jPΨJ6��g�P�p"O�U�&�Wk8m�q�[#r�"OV{���+/��a勝X_���g"O`�b�@6VĤ ����h���"O�(СDR� !�,5pU.��S"ONؔ��,4�0�!KմN*�"Oby@��ގI�R\Iu���P��Ð"O�쫃�q4-���I¸�D"O�����l�:e�Gh�c`,3"OԄx��i� ��$ۢDT*E��"O�IK�@E�1��*]1�@ذ"OND�ө�)z�t��&�Y"��8u"O�X�/0�D� �;0���"O�1
�Jbl���b�ą��d)�"Oh��Ef�j�(�ՂS�`T���"O�$§oص&r��a�E�l�<ع�"O� �0b2N����ׁ��ڦ�Q�"OX�
s��.�t)� [�t�)*w"OژJc��8��/|4q�'"O\����7X�Bp/nl��"Ox��4�۠@�ܥ eo4f��9�"O�h�GD�`PzeP�#Y-CF���"O��a#��0	�y!���0d��"O��� KpXx���r��cq"O��;�*��AF ��ұ�2��e"O��gk�1^����A�]�\�R�"OdP3%74�A��"��'~l�c�"O� +C�YIh�ĠʘUl���"O��	�"ĹX'vpv�GeN�K"O@�2ׇN:k��vl����� q"O���!�&l��#�K�d�xi�F"Od��wԸ'�"��qi�\5�E�&"O� [���'!teB��' �  �"O"=��ΙE�A2F�G\@q�O��'q�c�)���Sx�hZ��D0C-`�e��y2K\� F�����V#D����H�&�y"�E�8��p�U$ϼ)�VM���ǁ�hO��)�z�p�c�o�rN Q�r���w��:�S�O��e��Iû,�4��dG�x�HQi���+O�k2L@d�	�n_��l
s"Or���>bR�h��	�>�Vu���	L���)<"�vȒ�ʵ~l�Q�%jǠyW!���]��U/�Z�VF��r� �D{���'����$���:�@1��.�>8�tA�'82XI�Ƀ�4��{��!i�4̉�y��'�>�CE�? Y ��I&fᖁS�{��'��O���]w����i���T-_�R����ǜn�� ��� *t0��[�FfZ��6��+��UA��|b�O~��$�,#���(A�5��-k�,��?>!�䁫юuIo���>�����b!��7�:9���Q!�zi2��%_�!�,E�T����W#��� W��$(�S�O����V�5^�c�ːF=��!�'Ո���B
S�<�7�
?q@@9Z�'kX���O�F����V�[�b��l)�'np��������}�eMR]1����'���m�	L�����D%a��eA�'H��� ���tbu/�-i�dB�'�h��c��wh��H�i��+��qx�'�I�@��F�ݐ/-(��(i�'�>�(LI���UjH�rf�i�'�hi��.N�^M��@�>m�����'��]�!íy$<��m��@P�'��3TDű�* ��H�`�P8�O>����I��2�1��G�;����z�a}��>YVAͤZN��T�U�\��T��E�<A(ע<x����\�qr�34"H��?1��T?�GajIz\y��	��E(v#}2�'�(��'F�lR�.M4��}U��k�<ɦ��sf>=�1��v���j��BNX�@Gy���6��5p�`F�-���ʅ3�yr�H1l�<�d�	�ma�)�yr�[:&%*q�4U�'���h�=E����T� UD��,�l���OD2$�ԅȓw������9F���ۤ~� �ȓ^���إ(�?Jz����I�a ��'I�U����V�P��"k] j�N �ȓ,6��b�+
�$:��څ.�b��'!�}b�[�=��MzD�)6�]qpϋ.�y�l]��F��G��5�u2����-�S�O|ny(e(e�.��	zw�}�'�0��`E��rp��bD��n��'d�M���??�`�+n�IS�B�'I���e �%xUj ҷMÖ8)P�s�'x.5K�#0h���M�6#<��'�c�AT�Up�Q��G�6�^���'$z�S���,^��Q�m�2RҀR�'�� Q�U^�6 
�`ژ&�`���'J��h���qjF	���v}�
�'LM!���Mo����D�}�@�
�'�Jl�C�k����@�ʋ��$D��*���5kbT%�X�ߊy��� �IMy�S��ʱ�G�(pyP%��(����5ʓ0�Č{�Ԃ(�^)�[JJ��W.ړ�0<�D��$�֬�V��7%R�M"��E�<�&�Z?`ՠPIi];]d6��v�V�<�S$��\@ViI@J�:m�|Ը��UM�<�cf̃mti#���G���8�K�<9v*��\R�(���V�fqt�
R�<"CB�<>����"_�v��P�'c�d ڧqFQ� YZ�r8�A�KK�@�ȓ9���s�J�.�L�Q/�D� ��=q�������+ܐ�#�C�w6H�ks�P��y��J�IÂ��eAV�tT��K��~�'�"�4	�	#�-��V����/�y"�%Ml��T���)F5�yr� ��1 l�N��	�LL*�y¢	'y<����G�t�pR@��y']����bΌ+��2eݍ�y�lFh�(R�4$z�q�C9�y�(��y�`�z��F�R�p9��f�y
� ���� *��`2	��Qz�"O�LB��V$t�A�$��y��3"O�<`U��*L
T��C䙨CjȩCp"O���2�'��9��Hi.����"O�X��@�L���H�a׌�*�"Ox�j���gR�Q��Y�E���I�"O�)�d�Jgs�}$�0{�,���"OAƢݘc�^��A^�R�
1�"O�,�G��"0�V(�8�����yB�-8����	�?f�PA�M#��I]���Op$��/X-Kͮ:�Ș�'Sޤ�I\`x��s*��3�^�!�}B�'��+W4��b��,#��s�O���\�^��ߕfKT�I�"Ź�!����cbzI�
R	Q/��c�ñ:�!򄀱!S�IQ27ĄXX�������E{��F�
�jX-f�o�P��U�$(?D�p ���0�bH� �S
�����=D���$�.dh��sO����B:D�B�ܲ^�T��a�ۆb��i���-D��ca�I�7��Xc\	Sv6|� �-D�41a �Sr,�ʑF+E$�сS�'��'��D���l뀠a��{�P`8	�'~
�"�*�bB�A�C�~y��'iT�s�%̗>]ΐ��!M�Pb�!`�'�xբMIY(�l�"M9^��'K�L��
K$3�m�P욃Jr=)�'�0H�s�M�y@��.;K�a�
���'E��B�(�1�J�2�^b$��S'D���J�f~���	�8kjU��&D�<��Cn����ԍ��[3ƅ*� %D��B#����Cƻ'� &�/�	r����s�E�;�LA$,ãv��!1�.D�|��E�=0È`��n�1�����0D��Y�-�/��u���Β/<%0�.D��;�@��
�0�"EW�K�(�)D��9�ne�yJ�
J�/�+%cfӒM'��'��>7-H'lg�`���7hoX=�jTz!�Q4G���Ơ�*:o��p��zU!�B8/Аh-Z^Tu8P�M�m�!�ݵd���+�C@T�Al�4j�!�$T%n,���OU G� 1!�Z�[!�-_^ƙ�,�>f�Q��
�,6h!���?x0���!�m��&G��q!�Y��� �Q�Ur�)&�Im!��W{�0��'gJ� �)i�!�DЍT��ٷ����e9�Oӽ��R>O�xĦO-�!H5'T�'�~ٛR"Od�SԨ�u�nP��`I�(�Pp�7*O^�#l�z[�Q��6Gk�8�'�
x3,����h0�Hux ���'�t���͙a��͑�E��rI���'���� �_|�얓eD��C�'����6g���p��G8`ǰ�*�'Q���V(S?Z������Y�0z0�'��8*�K�s1�P7��+ ���j�'� �J��j�#ͩ�(Q!�'�B��ǉۊ2���s$��~��<��'�������1�ca��w3zP�'Z2\�@Ö�c��U�7ߴ7���
�'�����K��d�s��6}�⥠
�'�:�90�������eF+	-&z
�'�0��e�31j�\�����Vt�	�'��ջ�¬R:�t,	8e�Y9��� ƜIR)N*L����֎?n�ܪ�"O�d+��|XF�b��kn�5��"O썘`�	����U}M��
""O0�k!�;8����藃aG.�j�"O����2Xn�A���51T�
�"Op�g̉�4c�UB �S.���"O��K�ʈ�ec��(L�~�Z�"Oz�	%�՛+���P�a���A�"O�@��BQ�#(�!��w��D�"O� ��ӎ6w>�҅
�1/�h�t"OZP�dk�
��tz��J�]�"O�K���3!=�}@�Ĉ�.<Y��"O�@%êe���,��Qp�"O��` �I��(�O�t�r"O���կɔ/F��֍H23�r�!�"O��Kǯ�l�aF���3�V�S�"O�A�S�@f�ڱ��w��7�-D�tx塕�PD� 	=����'D�Du`�!�$�dȢx�@���'D�4�7CY2/�ޭsVbK�A�t��?D���7k'�RhAoD�?���Q�#D����@�	�2=��IO ^�tr�	 D�D�1�R�(�A��쓷�:D�(�͇/:'�u8')�T`6��.D�����B*�ࢫL�ow��%.D�؀f�K)����<2:6��P�/D����!��vo�Y�2�
�b��'!D��;ce�9T�D}�a�i��SVa:D�xI��|��C�p�P��7D��b�4@�6Q����8I�zM�P"5D��H�h�% e�@r-�5	�
t�$3D�@���?=�Td: ͬH�8<�$0D�@��[L^��Њ "0�	F` D��S��}������?ѕ�?D��jc!&?����b�7��׃0D���Ak[48��[:F��q:�K<D���w�1ҤA���%Cx�H�+'D���d�	9U���@RCT�J?�U���(D�$P�i�:!{訚3R�Q!��PF%D�4��Π���k�M L��Z�e$D�<)��܍g���Q��	(5L�[��#D�0{�+ʁRbL�ꃇ7+��,<D����\�PY�����f�N����9D��H%��(3&F=�(ҿ|�L��$7D��A͊ �~�@@8�~Y˷�4D��j�E�wD�mXE��V�$u��. D�8�/G�q���h[����M=D�p�oT.,��ؤ�&�|i;fD.D��uk�Sxa���"�>Q[&:D����	�0x�� ��+)�,Y�a�;D�@���AsJ��G��T�A"֭7D��a�e�sh(8�$%J�D��5D��J# �Qy�D2;��\��,0D�T�!�ܴH��`ae���xUi�J-D��j#� ��@�YbI6�@S�+D���go'\�}8��Y:PZ"h�.)D����JN�&]��BTE`5���"D��a���H%2r��0c�����,D�t�
�M���3GP"G��݈��+D���e��o�$�2�I�
�r�{'�$D�Ģ�B��:?V�R�%��iH!D�h[��T����|�b);�<D�@�$%Ɲwx��$g��� ����0D���$o�&���a�H�����'1D�� x��L���9�KK��J hv"O(4�"m�8n����Z=v�2��u"O��e�� o�&L�D"O���9JE9q�׺S$n��5"O�0Aa�D\ Ԑf��c�5�%"Oܠ�1L�7�8���VЃ&"O�QKg���lޝp.o���RB"O�`Bf,)w��k7ʄf�(0��"O@�
C(\�_�x�
al5Js֕��"O0*����D�8�?M�H�jQ"O��*��$ �(�n�`~F��""O���dV�+-Ѕ�dN�d����"O��2n�S��1�AN��I��"O���C���i��%��KF� @P�rB"O��0�# ����خI�j�2"OB����xd���.Ͷs�AC0"O�Ah�YʶHsED� $�=(�"O(�
����F�2s�L6RPQ�P"O�iB�,�3�N���aD=2�B�w"OR5;R��|�ᲡR")�A!�"OBqh�JƗ�t�pܷ!�D�ڴ"Op��T$�����P"�*t�NH��"O@h��J��@(�����f�P$"O��1P$Z�@��t��`� L�(0e"O����W,W���ȇ!�ANis�"O��9��U� ��r�@N/N>� ��"O0�����X	�M�BO�!�x�"O"�s�J�KLz8��-�&h�(z�"O�]Gb��>:D͇7!,�p "O|������i�qǉ�*�h��"Or�#��6�%jU3C1���AfQ*�y���-7��*�?��`�m��y2��.�,��ҮÇw�&�9��y�J
�$��J�	$���
#�O��y"�ӈ"�ֈx�j82��H��y���¡��A�yH�ؐ"W*�yb�1k�ɋ�D ��wE�yҩZ1q��u᠁�L�y�R��y2��Oxݛ��5u���N��y�gL�b�>`r.�"4�9����y�ꗡn�"�X�-&���4d�"�y���?��Q"[�;�0�d�@t�<y��Y@��(��lVn�°i�|�<9�n��n�AE	أA�
l�u��m�<!��
��:�f�
S�z2"��s�<�����.h���Bc�d���
g�<��$�r��������pрNd�<�b��\Rޱ��]_ΜɅ�F�<a!��|�+�/�p�eT��}�<��Z�O�`�@�Rpu�@��'J^�<q��#uN�������BD�ai��Zc�<1�����bNY! q#�i�c�<�cl�9�jԡ�aP��ΡceK�C�<4	>.��YUa g���1!��|�<I2�r#����ȋ�:T��y�<A$`�4X�e����UVxd�qer�<�&��� �ʼ��ޕ��]ف��d�<!���'��Y���pLҔ�Ҍ�c�<I�AQY^�
%(��{��i��^�<��	G=A�p�G
@�Zh�b���C�<ɱ*Il@:l㥌�t<DВ%��A�<�&�C�\W�|�ǩ�<o��-0b��@�<�Fk!tL0�Y�;��AYP�z�<�С��6%D����(�^� �H[�<� >)pC�ɩ-J���)�k|4�"O� ��H��S ��1�۟H|����"O�=ha��&T��l�Q���8$�K�"O��cp��KvvJ`�	��6ݺ"Ov	i�����ϞK:ҹP�"O,�S3G�iAv� Bd (>��"OP�K�ܧ�0�Cq��"G�r�!�dYu^�$���Cl��a�#�J�c�!��SM���dL[�z��!����S�!���8>��n�-a��\��)�!��*��Z� �w�(��
̚~�!�DJ�I\�e�7a�Ԑ H��L�!򤚣X�ىª�7E)2�	�L�#�!�$�&�X(�	�'8,�b�	�D�!���FS��QG(t��!G�P$<�!�G��0;%��`(��s���5#�!�C6g��`[B斦?��SC�œ_�!�$�&���\��3I��W!��̨OyB�eԉ)��uz���!���!Q9����D�k������1-�!��Μqv` aab�MX1�!�!�S�_�x�aD���5� �1�!�䊺vC�u���3�������"!�$��W�Ȩ#� a^" ����"O$�)�o�� )9�%0��a(�"Oj�Θ�8�ॱ��ׯu���0t"O��I��^.f����J�k�e�"On���Mi�<�
!�_3� �!�"O�Iڤ Fo�8�#ë\��h��"O(�3�oV�?�lp��'ϋ ��*�"OT�P�@�9(���4��$8�<�W"O����A�! 3���&&�b�ni�F"Oh)86d�'h��y�D
ò|""O,<�G�Z��E9�C
�QT�-Hr"O"�����o��T"c�q�����"O��#ڬa7^AI�L���p��5"O� E�)~��Rk�����"O�A�1IP����j2Ҏ�S4"O���pL�FN��ֆ%,� t!"Ox���!��)P�EY�;�
P"O(MDL�&���#$��t� eS"O�=j#-�-8���C �8����"O�pH!�R�(�zX��H�q�4�s�"O^ S�
@8 �:ЀS�E�XW"O�M�욑��E��	N�ȕ��"O.�j o�#rCn!(���3�ڽ �"O<���a� T0+�W�G����4"O�=��<�q4�=�M¦"O���@��(J9¢
��
Ԋu��"OFy���ؑ1UHMIw
��W�ԝ��"OZ�(�
O�F���U�qC�-P�"O��"��џ|ܤqQ%��c�"O�����ջ���Z���?>�Z��"Ol���)�2�($֏�j<��"O,P��������[�:��a"O��B��JRR�j��Q	1v���"Ob��o�7s�iÁ�O�/� �:"O�x�An�/�=Bǭ� rBV`G"O@i��'WI"4MC:{9���"O��$'��5Q�p�$m��0��5ѧ"OVxc��3l�Ti`�k&Xd9Q�"O@X�s��0!Np�C�)�nՉc"O��po˅E�� ����\�  "O�=: �t8���lM�D"O� �Y8���8CѠX�F)�i�b�j"O\ xa�*?�t��\)=o��H�"O���Jޢ`-��qV�W7*g�� �"O0h�v�=����Bg��Aa�lHT"O,�� ��ẁ�p�����E1C"O�a`�G,�:Dp�f�"9����`"O�-��k��1L"�%�d�|���"OZ-ze��(�d��CΖ/�h%��"O�pJ�!N�j*8�HuDB�9چ"O^��R��z'�y!�k����b"On��6��'m]��rC���=�6���"O0Xá7/��1���Z�8Y�'"Oܡ�W�^vi²�ߩB��@�"Ob� A*\�REq�0Qp�
�"O
��C�˹u�<Mz��=p\�p"O��ѧ���H��ч�2QuQf"O�LV�,�����R9L:v�A�"O@	�(�;<>l�X����|D�!��"O(I����ޠ��A��YO"�"Oh����n)��%Tzk~Y�"Oƅ���#���B��]�8aZx��"OV|ϙ�J!ř��ı)]��2�"O��x�[�qe�\G���p|	�"O���K����fDI#Iך��7"O�=��iB+SN�`�tL�-��!�f"O@�Z����qE�+�$ڊ2&��"O�)��ފͤx6i0T��"O�0����w�ܤy�ƌfp�0"O�U��@�/wU:W�ݷ���;t"O��t᜽9- ���z6H=˓"OI��>i�x
��-+/|�"O�tB�OZR���s�@��!N�c1"O�����LPܹ���	*K���"O���5���"_��R�W3L ��
 "O���� ��{E�)��>)x�"O�L�$��N�:�hR�T:*^��`"OuzҢ�!�m�Q'�"^��id"O`����W=QC~�X gӛX.@J"O����FF	L	D`�"��5J�{A"O,��$P��Y3!ֈN\��t"O.I�F�nt\)3��C+F��"O�D��¯9�\$�%Ɩ Vru #"O��an�}/HA���VC�"O�L� J�4�X�CT $ȴR�"O0u����.P�~Ai�� �'��x�"O��[G���~��aE����}"�"O6�@gҥL8�u� j�!&"�K�"O|4`�N�O�JȢ�jX�q�nx9"O�t����rr��1ț�t̔Eq�"Op8	���0u��QG^	9����"O� �e���'_~��eF�#�9�b"O*4�.�%%>\��R;si���"O�-�7m5�X�)Ԁ\~�Xr�"O���ǋ���X�[ "����"O��H� �'\ش�釨t�еX�"O���3*�\�fPY	՞b�U��"OIicC�7�<="��ߋaș5"Ot C��v���Y��4S`"OD5i�Y�����=G
܀�"O�Z���u��tc&"FB��t"OZ��T�ص �Ɣ�� N 8���{�"O䙫�!��{U� �b@ɗWg �hP"O�T����"2�4tX�N E]��q"O�ApW�ӯ�j�:g��"o�l�C�"O� �,G�ęH�@IR�Mg�rhk"O&�c"IņB�@h�2�ň8��	3�"O(2kȘ=�<���.>L+�"O"8cA�SEE2@S*�)-$*�j�"O�b��K6k+0Q��HX�q��m*�"OX�� "��}8FL8�f߳*�L��"O~Ep��8n�&L�t냫-�.	3"Oub�$�#v:R1��)�-����"O*�"� �%ne��ǨI��b��"O\���O�(Gv��'Ze���"O�h�dM�7*	qG�� �
�"Oڤb'�,bE��c�WU(3�"OR�H����0F�%fF4��"O��Y!��L�z	hEP=���"O��J��!Q�Y���8P���ۗ"O6��e�V���ˆC�9�.E�ȓ+h��jTOH(e!�C��
"2���BΌm1�
�1#=�\��k'����*08�1�(7T����
Af��-�X$X����>`��GB	
���� �H 5��(uB^���+[�S�	��p�q��׿}1�(c��E�>��up��p�Y`ڜ�L۠ �y��e�49(��#��8t��{�����M��l�4�F4\��L9WbՅ9*���%�r}۞�&p �Ҕ&�;
�1�ȓ$����v��3Ns��� �4|���ȓF������n�ޅArA��L����ȓy����GJ Q[be�B��p���ft�[  
�u< I��	_����y�A��aѩ9�%23�	�P�|��ȓf`PY4!�8H�5���[���ȓ+`NH�r��V�a3-�ht���<�8�4#��*�K��VEXՄȓ:y��+��M�N�Vm+���3��Y�ȓh����99�yIq	P�m�Q�ȓG)�@�A�J@	�����J�n!��pY�AZ�jT�Ym`$kr�M5�� ��y�8��kL8@F���Q:u$��ȓ0j�t�(���VQ� ��w�!�ȓM���
UN�e��]��ۯh��m�ȓ�ԩ���+0>�Z#����ȓ8�*�p�E l�V���R pT,�ȓDո�A3�н`�	!�*��L��ȓ.�d�a7 � F�Z��'��AeVi�ȓj�8�Q�%9��X1Jۘ|����ȓm@Pm+��Šg�|}�U�t��X����� ��7�r��
�K�P�ȓ�\�CՂ"�H��F�;%y(�ȓ,�.h�����+��o�67����'�t�Â�O�p�*%hU(ي �H�P�'s��ڤ��/h��Q�nƾ`�
T�
�'��M�F�/�yٲfR�a���	�'�B��'��>�r���*ݦQɎq	�'�٣Ane$֥�����BnE	�'J��Y��"Lԙ�%:p4���'R&H@t��06����#��8�؝�
�'�敘b&���2���<0~I*
�'�E*����a[�kg�K�s��5P	�'���J3fԎ���*@�n8��z�'�NX������t��,�"b֠��'� ��ӯ<�����h�i�'z�H`⒞	ze�u&�~�4i�'L�1:�ƆD��e��ڧq+�\��� 4%� c�\�$9��Y�n���"Ob5��2V��ш��;�&���"Ode:%	5,�l�D�U�CS��"OLJF�S>��� EH-%\tX�"OrdX�K�O>F�����~�!�d�8D��A�T�)^�r��$� �!�$��#�H��Aj��${���!�$��x��Be��R��%	��C0v�!��َH&(��(	3`�� 0�ö�!�PJ���I׍N�Ϭ�S�#��]z!��Oـ����.����q$ 7z!�D�M��8�Gf	
�|�*�CR�[�!�Ĕ��d�(  I�������&
!��ƽ:F�XBB�]'f�& �� �8"!�ď8O<���&��P�� ��.0�!���+ �\�)��P�^��)��Kإ1�!��G������5p@��j�5y�!��Sen�,g+�V�H�;ϑ?2�!�D�R;�]3W�S�E�4���-D��!�Ĕ5X��U��o ]f��U͂�!�䙪%_rq��fs��2���/c!�d���EY�K/5�X5�3.RK!�D�:6>lj�kJ�P�OQ�N"!��EΨ�Gh@x�Ը��U!��]�s��U��L!���跫K�!��6yh�R�'��1:X�W�C�:�!�[�*Aȕ+���
\r!�@�"�!���1�eA��]�ht���!�Dx�5 C���L��B�q�!��H��: Sd�[�Dܨ��)4�!��L��,��m���%R���l�!�dӜD�⡐&�
`{@�
�Ý4�!�d���{7m��J ��IUs��ȓQ̨R�$
xuI�������O�<)��9Ȁ��g��Ora�We c�<�DD��4�L�j@��YV��Fu�<YSd�tj��#��[v0ZH�Q��j�<Y74fp0�bb��(Kd�#U��q�<�b'�~�8�q�?�p4�� Po�<)aˊ�7
��*�!M5fn0l�(^h�<Q0&^&Wb su�H.Y�����	�`�<q�K��2�pI�.B4_l<#U�_�<Yq�)?v�A!��JEw*��P^�<���܂;͸m�*D�U]�5s��\�<�Gg$9�RW Y	
�^��e��s�<�W�N
q}rɨ��
j��b��e�<1��:q?�L�����j�����Kd�<!s�]�G+��q3�F�m����`�<Q5#�>���b�\�m�n�����_�<	ae�.������+pzPpG	w�<iB$@�$�Y��U�~Ћ�#Bo�<���u^h��䗸>��p�Q�i�<3*/&lY�1j�c2h�	%�^�<A#�[� ����Vc]�h���¡�V]�<! *�� |I��@��4`��\p�<9�㊲[�d�"����g�TC�h2�< ��X�~1�\p��0��B�ɐ�D�*b$(2�����-d6�B�ɽ7��a"Z.{-ީ2���2o�B�	Edp�ġؽ@�┢�"T>�xB�y�8�����8��I�l�^e&B�ɨz�p嘱��&�,�〉In�0C�	"E,�ذ֊Ͻ��	:פ�/?�C�I�|�ũ�BH�9��%�0m�y<C�)� $��lȂ>�4���W�<:�(9�"O�AZME0^w�U8V摨Q(�1"O@�c�����e�q�48�c�"Od%�B/<�k��E�"!���"O��K/�V�&U��)8Lhh�@"O��&"N�u�T��DAN���"O���fn�r���A�
�6׮�a�"On��w��C��|pC޹P�,8��"O��s���	Z��M���
�l�n�`"O^m;�84Cj}BB�Z,1����"O(}��,��́�`�$���<�y��ڏ�M:iT�"�v`��@�<Y�!򤐤�:]8SEɪ5��%�4�Q��!��-eCV���"РI�LP����!�d�O�����|�p�r����
�'F�a2e\�5�&���@P�]g����'<�u��/M�&mL���*�L�1�'����t�U�w�R�7gړ 8z�'t�6�"M]����A�)	P�Q��'���C�J_r�\a�,�S�� ��'��t�����i/R�ɐ
�<�H���'E2�3�AF�z�PY3��mu��(�'�Hi�M��u�H��Kєd�DD[
�']N��OZ���x�#H�F30B
�'n� ASk �ek�/t����'��(@�ںMq�"MJ"a��z	�'���2�	7IX�9�'����-�	�'¼��P�D>6����w�
	��0#�'lQtF�&z�i�0
�'�ּ�w�L�)
dI0���	�(ѩ
�'q�U ���	yC������=4r�����8A�g�iFfX��[�X��I��$�(�!l&JZ��hV`��q-��q@zsdִx7�0!�5F?H�ȓk|���.�8G�	0�D�5�<�ȓZ�ި����bro�H�20��*�:���=�y&OQ|k6L�ȓP�̫	�lRD�wF�VÚ܅ȓ7C���C!����Ζ("d�ȓC[�����gaV(��a��z�ȓI��I���H�+�|hRʞ� }"фȓުX�eN��S�b��bn���e�����a���H+Zl`�"O��ՇȓrP�0'(�%
r��H��v���4j9���>W�lӁMEZxP��lF�9@�یW<��4Άe�e��6C8-�0�D���3GU�&�����
KV� c�X U@�sn�*H���B(�b�J�^�x�	��Z�΁��i3��zrƓe�*9[d�܊@#�d�ȓV�@y�C�(A������?7��ȓ4���/6�ЅZ�%��gLp�ȓg�(�T���U�ʜ8�g���&���/���aRJo��1��^����ȓ>vx�T,�Iz�i�g�Ya ��l0�裳*ѳ	l8����̝*���QL�I��$O�+�� ��W�ъ���=�fTS%d)/�]�p�HYaf��ȓ=_����	,,B���AU	 ^��ȓ&`��Z��?b+���A�y�v��ȓ8\���*�9{ ̰xDOC!_*����S��8�R#�^
��4É7$	=��C��Hxs��&O%ȵ��6o��ȓqs�	j@+h`����_1utP���S�? �9i�Ϟc=���u�ܒP�l�P�"O@8��/E�!n�����VN�
<�"O ��jH�خ��C�F�$�'"O���D�>7A�Q���B�{K���"O<�z橊��������g_@m["O���@�F���[b
�J$��1�"O�Xa����@(K��G��j�)���y�I�Us�m�Ō���0S���yR�H�JT� ��d�ЂB��y��?1���0f��/����!��y�
�n��H@`Ȕv~���Ћ��y�ǘBR6��A��_LVi����y���iS��P�'�>+`�r�	���y�M��di#���.<c�
(�yB�ͧ��"`��5V�Q���y�/�Ą0sb����5`��Y��y�A7�B%�q�щV��	���9�y���9���Q�k f�$��ybA]$7��ich^�V0{�V��y�V1~������ �5o,�y�KQ�m/lY�o�	u���eB!�yN
�j���/Da���H�!�y��c��̑��F�Q�|ؒ�
��y�H;:���u�*N:���Ɂ�yr�?e�� ���r��(%E��y2�Zr��w�f��2EaL��y��^��d�k��e�z��!�%�yr���L�~��$Y�(6�Y�eC=�y��Y��zEj'ǾL�l�0�\0�yB�p�8� G��UѲ�UJ��yr��-
q�!#� QP<��doҶ�y��ڎJ{ !�����< \(�E��
�y"��Q����4B���K*�yңͯ{<݈D��%��xpJ��yr�g&yrE&*\@�r�eԴ�y2a�1:�z�j�'�3�ʁ?�y�L�ы�+�x|#1���y�L�z]��C�l�X���՜�y�
��l�QA��Y����d�y2b��H��e�G��Vyl�P%/D�y�N��Md9eȒJ�\���.V�y�D'`Q��p'f��:�(�:D���y�I Qq��1�*Q�%ۓ���y�n$����KҜ{�X0��K 2�y"�]�b�T��¨J0jŲ��V�y���'��x��h�~0:�;�y"�ڝ��-r��:Z@����0�y��*�r=���	�Q�.��p���yr.��|�1W� +����!C��yb��B����S	R*�����9�y����0��H����WJ4�&���y� Cn5�&%V�~U�(+�\�yBC�2�ౚb`�y����%���y­D,5<�y��Z����@��y���R��I��)DF	�r���y�c0V�Dyd)�+�pd H$�yR�B�<��%"���"T<��$���y���vT��/nf8J�����yReČ-¼ 	O^�d�f�z����yR +#E��/U`����;�y��ˍl��jq��0>s�\c�nD/�yBb�M���Sŉ �4���V\��y&ӓ@Z�2Q,�r&H�y�\�3qta�΋�)f�ؖ�ڍ�y
� ���*��+*�� ��f�$�1w"O��S�iL�L�C�G������"O��w� e����Є�����u"O����L*�R����0�
��"O���E�j�܈�b	�w���u"Op����"���6陃=^��2�"O�	t@G�o����%��w�Q�0"ON�냍�r�˴��t
I�v"O�<$�# �W��;{�jH�q"O>��քA<:T�]�ƌ�r�@a�"O�8y�J'���9�jI�]#J�!�"O��h��80x��b	F$H����"OB��l��I0�<{!	<7�Dj""O�p��ŗ+b� �8�A�N����"O��C�䉪�lm�D��<(�dq��"O���vG
*
(�D�ɪ5�,MyQ"O�}���ɘ���H�HId|�"O �Y��%~ ]C�Ȑ�u��q� "O8mЀ��:܀�fm�<s�0�p"O���v�ٕ�m2�L6]Ȏ|C�"O���fLy��[Ebڿg���:&"Ot��7f��ICQ���]8�,l�"OVM!੐�jq^)I
D"_��"Otd�ef2P�@ظ%�-(j�"O��鄸9�t�"��M�(V�i"OPA��I�L"�A�0��3:�<��"Ol̊�&��VA�g�Rz�Q�"O$� ((Ę�'�jd�"O�1���[G�Dz��ω\��(0"ON1�0�"]�p�*��E-{�"$�!"OV|��掩cH�,[�g�5I����f"O��� E��9�`�eF�<X�A[�"O���
9U\| k6�$4ȷ"O��'�A�Bi����ƐT;�ȂF"O�q��P�K,��0l��[#~��a"O����V�@�IC�K�ef��@��	L>H��ս5�\s�T5qi�Sk6D�|�Њ:��H��cR�S=�����.D�YBGE�+Z�sϑ_w�9�v� D���%�i=�)�a�P�)��:��$D�#ģ�6�bl�B�O"�t��I!D��(��O�AWnH�ׇM'v��)D����
%�L8���?��j��'D��c��@�.�z8{@aʐ�"1��8D����kk���抂�p�o6D� ��ɚL[<�����=RJN���!D����e�\�`��\#\r��"?D�d�'GI{>�d�dU�Fc>��R�?D�|�P$\gh��ä�ӓ3Pp��*D���$/	X'
,�Vp� �1W+=����,��'��7����L�Z���1�"O����P�F�v����d�r"O�E��ɖ6�h8��I[�<�Z��@"O���a����.Z�p�B��"O�19a�33;J�;u͏<ME�P��"O��!%H׵	l��s,��{?�A�"O�@�1lJ�� �3�XF�N�c#"O��b�l���^�b��ݽTv�y`�"OnH��B�(��PC���RgL%"�"O����Aߤ�sE�eH�)(�"O~L���4Vv^� D��:h/\�X&"OL��nO�<���C�@&'@J�"O�8��Gu�`��%cw�P�"O��g��.P�I����Fl���"O� B,J��ِ�^���@�9w���S"O���P S�n�$l�,�63�f���"O�Xr��7�4��N�"��EA7"O�(�d, ��Fn�>�D�B�"O�z)�� �w̗	~J@8�"O�U�Q-ZG��t�g)�_:�;d"O��Ԁ�5V�-x6oL�FK
��`�IN>�PK:p�R�#���L�(�YWB'D�����\�"-zW��hd��&D���!�	J�,ajƨWax���6D�t��W�=j�R/��<��5D��qp���E�ԯ�UZ�a�l0D�\A��̈́���a�H��,D�PPf��dD=�� ��px~ܚ�,)<O��$>批]�܊�D�(�0��@Ʉl�B�I'��9�-\�g|�q3U��36�B䉷;u�����[�"�( R�H�9�����&��R$f	xIed��k�!�� ��r<�C�6�ykP�ۖ�!��T�A�����I��~�J�e:_x!�d
쐹c&H�t�N��f/�Hv!򤘂N(�$K��P`�*c���v!�D<l��{� �cu(-:#(��~�!�D�"� A�1E����F@%`!򄁋_����Q!<'½H��D&!�D��iQK�5T�Q���!�R r@	�q���G.�<.�!�D�z�����'���fyW��
D!�d��M.`��똗QaPU��L�,U.!�ǂ{[4�5 �%1�"1ڳ*� )!�D?RX��A*׺�<`�u��
Ci!�x}�HZ Ak�:�
�G-z_!�³}�|݈�J;L���鴇�2@!�ޗl����Pi�S�F��"��*=!��U:v�A�)ǲR�в�\�w#!�d�V`@�gn�'��$ʊ�!�+�z�	�,�L���Ȕ	P�!�$R�7.��� AN�PRAʅ�/�!�� CƦ�@`�/-�&����h�!򄐧}�|a���ʹ<��6#�Z��C䉷H�l�d��5��򮂉@x�C�8{�^hCF�S�3��b�<o�C�ɹ<8��#�B]cvF�ӑ����B�IE8p����y��bO�C�	t�{����G���J �B�h�C�I�F58r�ô~������C�7!���3��:*cj4Q��A-n�C�ɨS�p�bR�Ӏ [L��\�C�ɬȞ�;��6y7�1+���G�B�Ƀs�,�h,��BL�Y#�9|C��"9��7䊝��13R[2t��B�	�d�8K0#�+x_�`����'�ҥ�եV�.�b�F��^�	��'�`��o�	v:�l�V��_����'�@�#��V�|ڈU�SoD�J:�'M�-"#���s�
I�u6�[
�'@�� ,�e�<��O�qv�A
�'�.\�Ԣ���=2��D�T�n(k�'���B�D���j�NE@�P�''x� 'թ:Rφ�@�H#�'�dj�^ƹ)��$�V�`�'JH�p쁾'�U����!�ZM�'���W G 8N�b�CD1����'�ҡء�V�j��m)�J�5��B��� ��X���S	�+�L��"O�P[�-��H�h��5�H�)�<
�"O>x���W�L���M�v���r"O�q��~-���S�
�6�"O$V��2�z1�R�v�@-+5g\J�<9$�ѹOv�����G�<�ŔH�<�$&;=�%*���4YZ���!A�<�%%ܦ`gbY��(�<hbD&	R�<!�g�G���c�ɒ0=r��(V��D�<��q@y5�G�L�~	1���00�!�d\8o�"�95k����4�!�)$!���d����5�rmqT�I�6!�d	 V�Z�@��("D�eR!���b�
u!A,��:ˆh��ʼ4b!�d��y�yC��5�T�`���23Y!���)u)��r�g�C�VM�t��%V!��ݷ"+�z��F*42��J�)x:!�DNf�X�+�J���'�`
!�$�+�ԋ��U�,X0@��3�!�G7;��␠�.l��91�l��i�!��N2`7F��bhМ)��aD�+�!��N G��`�P6I���.�h�!�d1��$ B2�`k�c_�!��$upa�n��b�!aG��2W�!���2Yd���D�*�T爜	!�dǏ<r�l�����Zq�����r!�P�Ryڠ���G6,�90g	)J�!�O;F�8u F2ߜ�1@�Y C�!���0�;�;V�l,s��Rs!�ĝ�(�����$��� �'W�E_!�$��C�,Q��		�L�J�'�!84!��-��8�f��m�8�0e["S!�D�* d�&Y�M(�h�:X܊�

�'j0�Ss�Ưr�A��(��z
�'D��97ɉ�%�����V&zL>�c�'l8��%�"
�!+%%Ƭxq��8
�'��p�F-��p�
!sc��v����'utm�Nׇj��0�c�p�V`��'b���� *OA���T"X_��Mj�'�m�7;6h8{�E�dw��Y�'wpu��'V��$�G%![x!���<D�� �^�?Ȳ�Ѓ��LlP��'*O�̱�!Q�O���`�M=q(��Y�"O�Y ����$�F�Gcl�Ղ!"O@���Ν[W��x�ݞ�&��"O�a"�h׸q�ڼ[�;*":�H"O��sv�Ϡ~P�5����M	tt� "O�&8O����� m�6�d"OV�0�]1p�T�Ȱk@7�2x��"OD\�"�оp+�ɰ��s� �	�"O�����j���1f�l�tThB"O�4��#�Wu���hλ#�FQx�"Opш�b(]����A� y�x��0"O��9�*b� -"PDĩMQlh[�"OʹS�P�X4jp2MP�(3ڍ�B"O��"w�۲x�X���<�ΉZw"O��k<dZ�=����=j�Δ!f"O┓6+ y�~����E�N��3"OL��:cbĒ�R�ČC'"O`����ۚd*�lC�E�-"n40��"OP4.��s��V�D?SiȱV"O\X�"'�0E�d]��$S�+Pb�S�"O���Ѓ�>X0(BCVLv�f"O";`�=g ��2���zkv��"O� @�W	B�:v~I;�dMjgv��"O�|�L>=�`�թ�cC��"O�q��=�d,�p陯{H��� "O�h�Ԧ�%dΕ1D��2I��� �"OL,��@�I8t��td�#!����"O��`DmV�A�� �cI���u
Q"O,ٹ���%LH,���w�d�"O2[�GӀ~^z�j�l�%)¤�;�"O
<�&�û
Ӥ(���=u0@Sf"O��a�
)��M��F�<=�6�B�"O���\'_I�qse�V�� $"O� ���X�!;pd��-�6��w���5�֑c������3�^�W���ȓU�R]�3N��n�5ʧEM�O8�ȓj&��r됳1}� �e� n�%�ȓ{. H�F­ El�y�k�BF��ȓ_�ꈘ��F�����]x�\e�ȓ�Ԩ�M�'�T�'��mta��D���B��3*���� X�����~�0��G��e��(���j��0u�,R�DfhX8R	�8TXVE�ȓ�)�7��K����A̿�(�ȓ[YP��k��?��|�f�Q�*�VD�ȓH#nŐsɌ1"��8むܵ�d1�ȓr/8��%ŗ2@�R�d: �ؘ��@u�Y��J������۶#F��q��!�$<�V�ڂ�Z=~���v���peċ��6AA�!u�A�ȓ@\ѡ���#Z�\�:�k�9T���ȓҖD�F��%��:/�h!$��/��Ԏ���Y�`�AP�*D�pC�`ʉ54)��U�F�Jpl)D�tI@E3�x�(%4l�8q �:D��b�W�It�ګ#!�(�
8D�@xC�Z/g� ��'[�\@���0D��9����v����V���:D�|c0��*�b�O�>� �ho9D�X��	!殰�UC����/8D�H)2/?X��@�$N���ތ9��1D��Cèm�<hh�����$4D���f��J:԰iq�R�]�t	0�$D��s�4�0��A��bئ���%D��!���2l�RL�a�lQ�g 'D��13��3�ؙ��)ϚV����R�$D���n\$6
PD��A22�­�g�!D��x��·a,�Lx��^V�9���>D���F��+* ��bp��;{��Ex�g'D����ϗ?"8�pI�>L-[3m$D����B�-F�=�&�90�(��f�"D����G�zA ��kE0 �|[�!D���$H�
`T��fC�%�����=D���աZm��(*��@�����O:D��9��M�2U�m��F��*�Q��9D�����ݡD�$
��p�؁�e;D�8K��X�v�D�u�� +.�) �
8D����ݿ!=L�;���G���z�`;D�|0��
�[b�c��3����:D��p�5-��!$�8!K�lQ�h9D����N�(�����NZ@�8�C8D��je@D�)��� @��r��m1D�F���0�&�F>0r��.D�0C5�J��0h��q�����)D���bc�?9ބ|��	݋��i�d�'D��Y�K(K4��"I,ġ�S!D�� ��qP����QW.�n��v"O��*⅋1o�v����r`�<��"O������B�"\��NN�t��=��"OP �F��?~�aRЭH�Z.l�"O�m��U<�B�IЭ �@L�iW"O�9��!�~�Y�d&��`Ag"O�Y��;�D�XkE�4��7"O
9�7���{ �9&BE�6aP"O.D�`J��2`hk`#�e�<	E"O0�a��w_ޥ1�'S�l�fH6"O� �@�&�.���d�4�^�y"O8m�P��TĮ��QD��ϰ-{"O��b�i\*=�92��t3�"O�����\X�l�C�E�zz��[�"O�I��ʟ-QPִs�M�:�b���"O }b�D�3��p%�	-5�f��"O���g�F,�,�pA@���~���"O^��Gn62��#O�p�>L�A"O�5(��$�I(�� U{�=�"O&�&� Ԉp�VZ;���"O&�{2��&�dD�ѣ�=_�Zūs"O�%��u$^YQP�I�����"O������k�f�0a�4��`b"O �N�����W`��@��%0�"O�Q���ĴC!|u;�/&dj �"O�53��� f��k��,�,�)G"O~{h]�+J�(�q�ܻh���R"OR\`�E3�֌˄�ͤ�f�Q�"Oĉ� �;T�|Z��+�y�"OR�/P]0d]��K1q�Q"O䬲`�����z�u�`T��"O�ta��Cڦ��W/ȍP����R"O��������i5N=���h�"O*�@%�R�?S��an܀'���C�"O�E'@���`�0�	� "O>�ȕ��UY5���~�$��"O0�"�E�7`sqHI�D��	�4"O�!�g�	z��ыb�s�t`�2"O�(G�͊k��pҰ�]�`��lh�"O���L�0>t��!E x�pc�"O|��K-/q�g-mTM!�"O0ț¡�'	��Q�G�Q$p�� �q"O,-9�ʋ e(�;�����8$"O�c��&>,��RK%D�`� �"O�,�m[H+`�4J� )�"O6��͕R�xg6�T��"O���m��B��|qb�8<�T�"O��#�C�R��ey�斲g�q�t"O�ɲR��.����%]$]O��A"O�)d��>r>D�@G�H<8 e"O(�!Q>���Δ:Wt$�"O�Y�P  �;P�hsuK�)c��h�"O����+$L�J9���;�F)ش"O�hCc]�p��PE��R�4��c"O���!�m�Zy���  �"O@pI�*\=�������<?"pL�"O��
��P}zV	��]��"O��q���*z�.�8��4w��y�"O�Zc,X8_%�x� A*\:բ�"ODU�ӫ��?�d�A�m�xnu!A"Oq'�&oZH�M�h9��"OV䪑D�H�HmA�
�8H�psb"O���2��8B�THԯH�T�aR"O|@�����UGh�:�A���{�"O� ��閂�y (	�%��W��ͳ"O���doÓn�
A��o�=P/25hB"OJPRR�&��`�E�}T`���'K�'����
�><��ʲBΙ�H��'�R@��HO�������� 1C	�'���[��G]Zr��E�3~�^���'�B�P1$�yf��L8e�M<y�C��L!4��9}�Vx���#
� e��n��]�<񕢁��j�[D�Oxc�5��e�c�<A�a��z�t=�LUk&V���AG_�'�Q?��J���S0�J5mѲ-�IB��8Y�JO	E�ֈ�sG_�� k���G{��IŜW\,$8��	rbtTR�EW.M`!���
<���d‛fV���F��,���,?�	ӓ)<f�u�D<H&�%���6��y#2h/4�L�򦗍.�$d#�NX#=`1�`b4D�Ċs���P�����B"��P��2}��)��+Z��놌�"a2 ��@�(1C䉰`�Ь��c֓W��U2�(�Y$C�ɸ6\���O�O�����֚Lf4B�	?�JIP���"@|)G.Ʉ^�B�ɼp٤]c��ǵ|�N�kc`��=��C��8i���cQ���Z4L��y`��'�T4:k�!	�B��Bl�ê���'�!��JA�) $�"�J�i�Ly(O6rӈ���[��kt`��B�^���ˋr*!�C>;����%�"Hٌ�a1J�+!!��Y8\L�f@έq� �]4,�|x�으��Z6�.~݈��ַ�y��AC%�� �ƚ*�����؛�y��̖G~�	6hѐz������D��y��ʓc3fՊ&D�o�4��eNλ�~��)�':~���T�$ąQoH�_�h���][H�S%��d����̺(��ͅȓ.@Ђa��QV�̰�)���~1�ڨOv"<ith�6��$`�
C����	���Z8��&�l���"o6��#DW��KqJ)<O�#<����QFp�(�]�(��йQ	�B���<�O>����XȚI�&� 0U�.��v,B�˰=!�׷.D�D�oD!wϾ �w�WB�<� ��*�@L3�I��8
xY`s$~��p=�W�Z�9�|�¤ٕE,d��{�<)�(1CN@	���K�"��Iy����?��۹Q��\�M\�Y;��l��<A/O�O�n,�')�\hH䦓Jb�t�Vp�R��ȓc�b��2��%e���+�Ⱥ*TB�I�n�8s𬗷������ّu[�C��$�`� ��3',�����*|��C��q�,����4a��lc��	�>��홎��)�<�5`�,�  ��nB.7�b�h3cO@�<��-M��1A���0pp*����
}�<�FH��>r��y�GT0]Du�5+ t�<�t搀M�$ݙ�!
���dɄ�_o�'��x�OZ,�tt�[+����,�y�%5�@ ��� �@88r���yb�:�0�%!'��q���y��ޕFx��N/;���s�,���y��F�!�%x`Ɩ�d�8�-T��Z�'�D�0�S>��� �ҢCE���'|�sB�o��l�S��06���3�':6|�C�ۃ9���3&�<0��5�
�'�v����>�ъD��&�ZA+�'w$�u�D����T����a�	�'��yg��#��mS%�R��$T���� zQ��l�Q!l���*� ���W"OT�x�+�bd���*�0٤��"O�m*EIG�5? *� �}ɘ��6"O�\*1��tJH���� �_�tE	T�xR�)���w��yw%M?-��0�v	N�!��7�<�DVi��;��J��ǘw����<D�\x���5TdySl�:Ӱ��v";�O O��q�iT�G��pv%��*n�M��"O�ՋU����0L?�i6���y�.� G�B�#��̖��c���'}�ў"~�m��h�Oۄ+�V��A�/��v�>�H�"~�	 Fπ�@�+�&E
>��1��Y}dC䉭z�8m��4[���c��.�B����'�џH��mQV�����`�9�@�0�3�O�O�Ex�j�M/�9�4�9,s���R"O �z#���*����:mJ���D1ʓ��w�, H�-��)�$�O������D5|Oֵ�©E;G��F��B��paO�p:DH�6�M)����8�KR��`�<Aԅ�I�p��.F��PS�bG��~��|R�~"�ʆ\��E��۹m"5�b�Ua�<a���ZN��[����,mLlȶn�E�<�� )pP�²��.�xW	V��>�J�L���x{Zh{3J�80��m:�O>�	N؞H�O�$VB�p�@M��r���:��hO�����$�DTm��fł���ȓ}5���v��%$�V)C�}�@���Dx=80�V5^�(�5���0��//��͊N�Q��Ǵz�����ē���ӡAR��pTc�Bu.�9��W�a��C�I���R���Chm%��9dTJ�O2�=�}"¹r��������8��Ín�!�ܞB�"��b�*W\� �Q6O��!�O�JǢ�Qd���k����i��'��)�3񤈼7%������'	��e��)&�!�D�b�D�cs��O�A�����B��>yL�𤎄^�j�
'Q��C�ɷ]t�mbf�;Mހ�4� Y�v��f��h�x�@�E�>�b\9eiB$%�
��t"O^���Z�#M�Y!�F�h���ё"O��`�^�'���a��H%�~l���d>}2�G�q ��I>q�)�=Y��9��ɋW�|�!�D�O�ys�܃x���&B 7��S��>�B�����O0�K�#��	PnhI�^-zD��y��)�v�$�A(��Nw���ǁ9�����p<q��W�D0��6�қ|�}����V�<�VnE�G�m�"�A '����l�!�č,VO$%�7AX�)b؛ i�>E�a{C]�I�]�|(b�)��G� �2� WN"C䉀u�J͹2�$A/Бq�A:g��B�I7ƾ�f�H 1\С�Y�d��B��G���cf� ��]s�N�m�B�I�R9�Q�Jӂ=j�F�mv�B�I�4��&W�ҘѷI�;���	�'¶]�6�D>{�m�t�Adj�`��'t�d8�Oء�[}~�@�!��I[�,�dx���'tI1`�� 2��,�8.���'����'d�8#T��T�M*��`	듎�	k��B�n@1L�ʴjF솣9iB�3��0��_S�� Ï��<BJ,��Z������<��	�䥜�(�!�]>5`���ǖb�`�Q$=�!�$_	U� �V�B�!%��Q�C�o�<!�(ͷo���*G�4n&��B ��n�<� ��'Ϗ� �z�b�&�"��'Hў�:�=+����Wȍ��|���H�>�' a|�a����Ӆ� ���e��;�y��,X��Q� �F��Y`e2�yR@� �0�SRÒ��na*�%Y��yB��;j��4�+�;<V���4]�y�%��{/&i���&
�� d��y�j�u��ݺ���$p��g��y���%:4��K���@0TBÇ�yҩ�%e��h����-}��A�B����y���O^"4�0)�5tк!�b�	��y�"��!4�ӥ�6���1e-��y2ą70LUشL�6|8�8dnF��y��̩S�
 �U��'J�e�f�ט�y"d6
�֙�' � �$��D�ۑ�yb��hӢ�`���2�qd��yr��5>Tu������X����yr�{]ӵ��%�Ό��G��y��`���	@���iԮ�y�1a���Q�)ŷ~r��S�
��y�J�0�̵���'� ��a��yB�Ë9N�drAU4O\�S1��$�y2!O�wo"�rɅ;i��I⌥�yF͐#7 �S�Gկ6f&Q��.˪�y���>$�0�rbK�.�8�ԇF3�y"ek�ر���2*{j��$O��yrʟ4_�2H��Ě5)tҍ::�y�O2O�
A�q(͟(�`������yR�H8o%��^( z$�bH\�y��������a�gl��q�ߘ�y�#�uDĕ�ӈ�x���j��>�yr�3T��f�^' � *���y���P.�c%�D4/)¹�B�K��yҍ ;=`tE:��}��ݡ�f��y���	��K�DҔ��`Wo �yB�ǢXO�H �y@����/��y�=3T-H�j��s���E��y�k�?:�(Pr��G�l�V)�0)Q��y�jRC!$i`�kL3_��e0�m�3��ONqr��E�
cf���?i���0Ol�k7��!�f��R�TMn&�z�"OȬ�I�Lр]�1�@� Z����"O*u+ dO�E�6���S$=�P��T"Od8C1�ɭn��ڴA�� �z�:a"O�ٻ%K�=ks�D��Q�e˘���"O���ղ3=�BB��%8R�j�"OP�4R�]���� ��5}����5"O��Z��NG����z��)R"O]�r/ pc�m
u��X�=��"O�dX`�6zBL;�`�8�q3�"O`�;G�N�*��	�e�[�$�:c"O�T)�ǖ-1A�*׈^�=-`�"�"O�Sa�J� Q-��~
4+"O(�����z�T�j�H�&.ic�"O���p�&h�Х�_�4�e"O���(\��)��55�~4��"O��ꢧ� .�,�h��- �f�x�"OX����~��m{DG�w��-��"O&(S�(�=h�HK�	��	��"OXs������X�(�&#6���""OB����̒ErT:'�=*v^�!�"O8�KW��0\[RR�'͐3BM"O�h�Rf�,s����D�W�.��S"O��4`�68=��,�5�&�p�"OȘ���(N|�9���ťYu2K�"O� �3*b��է�:
M%��"O��6�ڥ
t(]�dE�$}Y�}[E"OR����6/w���㫕#<A�PSA"O|�S � �U ��ze�`�"O,l[#��7X\�H#P�ѓ"Ozh��$R�S�͑�����q!�	��Q?��,�]���KDI���i@�m8D��hp��$9ꈄ���- .��P�	�O~\���(�)�'b\\�Չսi�΅*���>k�>���'EB�`e��~F�zC"B�W�m��O��S��V��=�I[�/�D[��9�:��[rX��Š
5g��ς,qk��`��S�B`��a��y��&'�Y�Q!�����`í��HOh�#R��h��PcEb9Y�Υyq�T�^o<
�"OJ�i/	��Y����!slx��iNN��!�t�S��M{��CC��h$�>��1��^o�<��J��TyS�F���1ĊGp}�jq0h ���^�x(���X?�l�4�P�:(��Đ� 9,�I�*��әP�t�$�T8k�vB�	�E�naQ�mZ�p�"l��U�2VB�I�_�|�Y��fLIa�(P YhB�I<I�1"������t`K�N�B�I�G{(�i%Ɓ/WG�9�"I�=MJ�C䉝�]��h^��ps�D���C��	H�6���[�t��ҍ*P�I 1�(��@ɗ}�*ل��(L����f�� �5iS�^��$�e�"a�s�+P�40	���`�K �o���YSNߡ1{Cቢ�ȅS��y�
��%�����d��Y�����)� �KF�i�1����H38&&y��Ā�
!�d�M�z�ZVό7���a"M�-�@��D+g��hS��_$�\˲�Zy"@U� ��UHFA�)v��
���x�a�X4�"DB�;ȌAuoA!cƌ}	��,G(\9�C��V�*F��W�'����A��"WU$��p�8��9˓E��D8AA�:&v�A���60�|�B	U�q]6U����&�&����&/�T�Y3���gӓ@��)��'ҹj���O*eC��O%q�x%�S��?��}Jr(�7\�L2ϟ>�Ӳ��>q��K��ȕ���!�"OƘ�����<��#�H��&�(�pЦL\�(X�C菳a�(tPB��jq�6<��Ă�y�������0K�;���x���2�x��	��dqA��zAH1I�&�3��Vr�|	��V�08�4��»a�nA1퉀44ڥ5�:Q��pթ��o���E(X�ޝz5�
*J��U�`�����Go ��c4W){�,�i�m��`��>�O9�G'i�L����t8��B���"��)8�P,��*@�,;��
V��(<�t�O"�]�AeO4-���OP1Yb@��'rm�"S6T�>� ,O_?��.}�"T1Q�)Q�`I&��NF��H~B�'�.JN�ͻ���b�T5�x�e\(N���������K#�� {_¥ѵ��_A�!1s���4Q�%�GE][�bU��D��7b�yCe��U���*ҁ��Q�ZIH�d��h�d떁-O�ꄊ��$Öm���ٴbL%�`$_$4�ԭ�Q�A�7�*`:�eX�ez㌝�f`��	�M�v�	�b	9S�P ������)q���p�U�07DYiP�[5mBɢ��	^?P� j��9��{��ϘI��B��V�5��Lp�fĠҌ�$�%H��|� 4���p9t|q�I��A"��O?͸�,�k�:��BɌ�
����}YG�U��8B�I�C͆�S���?^��GL�;"�c	R�LѳG�)x����Ca�>�,�c���=zUQ��	7P<TĈ�u��_&��a�1O歂`��.x�,�J�)�u��K���=<P��Q���n��Gi�01ʊ��c%Z7�d$��a�l\bA�0�l��qd�!~���'`��p�#@��!0��TN�t	@�[v8��)��@�r��r#��Z�հMM������T�<	�n���"�*�`��z'Hu�p䃿t���H@j�ti�'"F4��.>�D�ĩ,�dȟw���0D';X�%a��;VX0��'���o�V~t�S�Òa���E��	�Z�I�'F�1�"��fI�X�p�Pϕ�Uyd�Gy�cN� ���h;q�*`Z���p<	�fǢ����iT>o�*�X�c+��	��D�\�e�-��)���"���!LIإ�'|>ġQD��tg�QB����̆H�D�%,��Q�(_�{0ؙ!�M�wa�Ab�B'����'3�ظ���"ə�a����S�? H����rp9#����\�}����5I9m�W�2qJ���A��Y_D�L~��'Y_�n��s/�����Ӎ
2�	p�FkC����=e�X�ɤ�Q�]�P�B���O�Z�Kv	�O�m��E�f�� �D�E=�?��剎E�x�V.@�6grx�ǉ�m��̛2::`��d�4�{��z1��$��p�T)|$����M��X版�p>��k��	�\���eT��Pb�|ܓ*z�0�\��\��7"��	��$�!3�����U�mfe�� ��yB�W�P������D��N7h�z��HP�I��Ka$Пp�F�7���NV:~�n�H�stީ���%`�!�$1��щ$)bY�*�,���<H��@���HO�0�E)u�z�w��!�ū�3�y"A��<r%j�31�ҭ򃈑 ���|x���R.��$�Z@�j�B?Ā���1�O��pW�U`�#�$IpH�B�3\1���<{�+� iNq�v�^�;�ڀ2A��U��=(�F�n��9-�ڈF���Or+�c�5*, �d�74�"Ox [��L4jܲ�i��k-��s��G�ON��t��,	�����?v����$�"xa�M�ƥ�y���F�ۤ4�a|��O6;� ��&�<1K�P��� �uh:�0� 	"0f���$�%HK��Ikl�<1tO�1�kӯƙ�HO̸¦d	57Y��7K+�S�&o�!%��:^>6M�fI�,$�`C��'>��c��` J@ ��
�B�IK�Z�At��F�*�GcM�n�!��^9FR�R�_����å�#$!�䛞E�,�v!�ev���.W� !�ɉ�bd�e�I�B���S׭��-�!��ݤ�01��
Hn�E�wk�-�!�d!:���	�
;�4�pH�|�!�$@6~�\M`�MI�O5�h�2z�!�\4Q�ve˲)�+C#lQ;FH^2x�!��	o�5��D9.�2<2#g��3!򤚭�DI%넨��H����`#!�d�N�Z�{��ĤZL��X���I�!�^<ql�p�G�ҷ5`�P�Ȏ5;�!�ӛ;> u��GC�aFD`���&�!�d�L4
T]o��5)�=1����"O��J��\�B۞"n6͢�"Oj��FB�,M�m�pb�7Z�Ը�"O�E�"ꉰLJ�Ha��.Ԕ�%"Oh;"��6�������08+��S�㟒��� c���
�ꤋ�Y���e"O(�pg�-0�m�V ��Jc��IaeR��'a��q��>1�ΐ uZa�Q��0�T=���]yH<!t��.,HAS����`/��^�F����յ�p?i��[�t���*��T��؋�kX��)�Ȕ��f��OvH�BI���sA`��,�Pj�"O*��f�/~���bvn� x������x����%+5�|���L��'ZR��c�.u����jU9�y�_#�T)��w*��� ��"O�-%��À�%����2�:��%�X�h.ҝ)`D�Q�r�ēL���ҋ$Z�8u�P���h�p� ��/�,]���k+X`i#O]*Cۈ��g��&����I:W��=c%/T|�d� Xx(���]�U�J-r�K�� "!����rES�mG�=�J0@V�Ɔ4�'yl�X ��jɧ�Os�1 �"vWN�r��O�FG �(	�'�(h`��C�rM#(��>&�	ڇ*F̓?%���L�`C'��-�PM�5{�~0ca�=D�p��
 c���zG�٢%-����d�� �t�@�VX�-
HX�(�vI&ɇ�>S�zD�ޫ\������3v��{��:�힥 ҄���ąO����ȓO��sAÃJ�.T��*�]eR��ȓl<D\��'ķV��ҕ��8�( �ȓ{�$]��L�P�<���bW;y�Ѕ��S�? �A��LШv�8��H�Mj����"Ol�*e��/^j����,Sp�ӄ"OJ�ѱ)[8��	[Ola�"OX �bް#����e`��p<8��Q"OJ)��3fJ���+6�h%"OZ�;C��I�H��.�D��#"O��(pL�:nu(�;w!&����b"OP`�ӍU�o@ġ"T!�4r��Q�"Oru�� ��p� ,��Y�"O����U�h,|��_�6���"Ov���@����Z��ہv�`p�"OHLʥ.ƻV`z��E�
O�����"O�蹇�	�p�
�$�"�����"O�ek���Q;��x6�K�a�`��"O`T�ץ��Mu���π9�aC�"O�m�!̛)z�y���¬{���:U"O��Q��*p�lP�hOJ\ Q"O���:n�<1��P�Z�a�"O�*p�90��ӡ��$r� ��F"OĠ�G$�]l����,F�Ś�"O��*g�u�$�l� ���"Of���d�g^����6jc"OJBo^7�2�IҊ��j��Գ"OV��G��r�̡"�&[�`����"OX��FF1�䤀��)C�^�"O.�rͶC�1�t�
>~>xD"O��Ɇ#�+Gq����)K�>V�T��"O ys7+P�Al(�)��[w1��"O���0d,7�piK�#>h4��ˢ"O�x��� 0jXآ"�0u��̸Q"O,��c\1<2\�B�Pr�ZU�"Oj!�b
S�,����ڐ`��a�a"O��H��)�h �)¡T��P:"O1Pc��l�(q��8b ����"O��y�m3M_d�C�`0=��5"O� �`gѤS�n!iF/��.K\��y���_`DIp�Ϯw~��`���y�YK6y�R؎q867G��y�l�Qa�x��ϐ9Y;��:��Е�yr�C���I&
Y�t�R�&���ybʖ�� �q�K��T?��S�9�yb��tQ�:��ץV^�Aɖ/�y"d�"�(�hp��J�܅��y���7g�E�c��+jF(��%"���y�4(":8"��n���5h���y2�ߵM�tH�����x��E&���y�E[�D��1��-0aP�ҔO	<�y��\R��2r��$ tZݱ���"�y����j%Z�K#J�T��w���yr�7}�l;�
�>%� ����y"�1>�&�Jᨐ�0[D,�H	�yɐn��Vß�F�ΰY�-�yr��(���"��&:�������yR*�44h�sE�ޅ>��U��&�yR-I8G����(\̍�5o��y��\,R,&����/Fpj�+�y. 5l-6M 1׎4�p�Q��E2�y�������%b�6��:���yB�_�s�x4{A��
X5��XT����y2NJ�.v���Չ[V�$�#'H��y��u��4G�20J�ZSn��yR���炰n���h�Ž�yق�y�Ѕ pv�$�r�]�y�#�8N��(��9�&%cǤօ�y
� �#�	ʵ
�
�{pfY��`�(�"O�1�O��P3)cq��֜��d"O` ��̟?0&�z�W��ո�"OޑE��>Y�H��f��'3���"ON�@�NJ�wv�8ce��,V�Vy�"O�A�LR'!h�����a"OB$�E���C�P���@�D91�"O��*M�;~�j0B�4�LP��"O��J��Lu`BY���R�:�"OԐ�ɛ ��t�� /��K�"OB�rK��.܄<83쟪q�*�h%"O����n\�a͎,��)O�.I*��"Of���h
=N1�4
)�|M�""O��&�`�2�u�C�r�DT)�"Oxb��'��		bi�>:Q,�AD"O�u:7�fp���7&J
w
<�"O��25Kr)�b3x� �h_��Py��L�)f�q�!ȁ�5���M�<فM��<Z4�f�i��#�o�N�<�E^�5�8�&�B�$��d�I�<ѣ��_�^�qM �:�%��΂D�<!���k�B� 	��Y���Jq�D�<ɵ��8dp��sK];?��j!��E�<qǧC������2�U���x�<ɇÎ'!@b4����y��*E�r�<	g#�,/m�	#р�v�Y�+�@�<�ӥנu���k���?�����.}�<�1 F��!	�܁n�re�%�x�<9E���&�i��\ @��u�MJm�<qS�F�u,Q	�$�	�,����^e�<Y��ӣ� 1&셑I�۳lc�<��
�-���2n�z�	�ŮWw�<I���z���s2��wK���2D�D�<$��5[M�t��OQ�O����
D�<��70o4��FրFt�b3�n�<YeiגLe�l��O�T?�=�3"C�<9S�"RV�� �\�I´�B{�<�A):�����G���6�q�<�IS�e�N8��¾&� C⧛{�<��,��}�Q�&���o�)�GI�<��#&M�ܫ�LZ���*! Yl�<�!�._����/�1D�|!���YU�<)f�Ua�)E��r)��jW�<Q#�V�r���8��A�_L��I�#�J�<9����j�I0���07���gPZ�<�C��./��xi%�.=�T��n�<qw�Q(���iKf�����\\�<�`ѩeen]рH 30���w�<��(��V��aA��}���S�#�v�<�m*'���kA������k'�Vn�<��
�t���3&�;�VU��
\�<��I�U�	���Y�gi�_�<1�
 g�\�s��&��ey�UV�<	Ec��G2�-�J��EF���O�M�<��ۏ$[,*'D!u2��D�O�<�6�J�w=\5Z��P�Dd����V`�<���.LI����CŨ�^�<��ŏh�;A ��$D���X�<�U���T��q�]�{�9�2*CV�<�B힨�l岢�ȩyN(���nT�<�w�T4k\EHuS+.+���B�P�<�m�m��Ԙ$�O�H��]R�<�ӧ�/n�`C�&]2w�0K�	�e�<�� P�f�my�h��~��F��g�<� <D�3':^��tk3�2�x�"O���"˖5h�4[rKG�DaA"O�ɋ�Q�N��ebfO�vuj`"O���%��;qj�j���h[�"O��Z���O�:���ˉ�=�4�"O.��'B&8�DM���R����""O���ЏX�N:R���,W�����"O����ˎ���P�&n܎t��0�5"O��᱈L4g���)t��I� `"O�Aa�V�6�Åȥb�kp"OT�q1n�/<�s�ЧH���"OԭKW��X^X��B�(?��A�"O�(���̧c]��P�#��$f"O�E�#F]���ytڃv����"O yq��]���ڑ%��d`�'�4٫�O)y�|K1AC'��!�'@��;���,�20( ��:���Y�'c�z�[�Y���L�� '��
�'���O�TQ`$���1#
�'�&ThTB��K�H(�(õlQ�	�'ub}�'��7FP��g^J�xp	�'Lb)��R
rf��QB��3+"-8�'j�Y�5,�� ��X�.��q"�'#��XD��}�A� �0l�'��͊Fڎd�^�p�266u��'�2@ra�~	��Z�>m��'�X�F�"�$�ɔ��=k�:�*�'�I�+��B��z���m\�%j�'��PU�=AJ�c!a]����'�9I�f�̡�IC��N�p
�':�t�f$�SxF��BaUx<�̈
�'}����Q�3
�i����y�]�	�'�%C��Փ&��ٲ.O��@�'f�Ke���%� x��@ ����'dva��O�Y#l�`抚-�h��'V�I"�)ٯ3EP�{׌͇Wڴ��'��D"C��A�9��#W`���	�'���p4oK�: �������6�����'%b5�AO,����(0�|�s�'��A���y�F����&��K�'�L<1e�Ь<����B� GR5��'ڮ�� " V���� �^5��'d� F��)r�R4e�H��4p�'��A%jB9S9�����3n$"�{Rfǘ5�O�OU�\�&�S�z@� �W�U,̺��
�'�����` -am���C�ڍ"��� +�J̓#�����L��$��0>�|�(�茀z;@�(�d7$�@�$-�xc��@�*�[��`����ї��L���c6&V�G�(���ۗ{�@(f� ,O�MPGK4*�>�'~� �N��|�49��׈
$�P��'x\uC�Cbv�Hw`WT"`�H<���?��X�L>�~Z"���� 1%�G �����X�<�ӧK�k���BÉ�1F50�-Y9x��O@)`vm�C�g�I�[ޭ�7����a�T�V,B��t(�����Q�,1+�.x�(]3�O"<eՆ��tN��犂�c��:!	A����>�0 +�2}l������0O�Ƽa˛��y��?|UF��'�O=�h$��b�)�ē%Z��#��S�1�85��'�% �0PFhؕK��9��"4�� �K�sPВ��� �����y���#���7��!��>b�LP������ȓn�10e��5����_�|q��9���Rta��]6q�����O6�ȑS���y�'O)9�`�8Q��*TCФ�1�y
� �e�s�C�݌H0p�]��:�"O���q�!8f��(�g�&S�骃"O�1�U۽Ac��R�`���zL�"OQ�&bS{D����Ď'Â@!U"O��i2�W&$diڡ�A�>Պ�J"O��b�@@�J�U���$5����2"O�ay�L�Y�����i"O�ɳD��7���1��3F�DHɷ"On�j��Ӌk���$��.Mp"O0���OH7X!�hD+t �xC�"O�|{J	���$AG�Q:.
\��"O��y��g�jX�dޭm�\PC"O}3�"��(�]�g��H�"O���U�ߤr��{AL��Q�PH8Q"Od(ѤǻOX�%�0�L�a�a"O�m��{��jv��/ (��"O��3��6�(����)��`"O`�b�@�V$�rDd�`���rU"O��A�
�|$z��C�?��d"O�Z�KW�skuH��S�T����b"O��r$�IF|��\K�8y"O��S�/@���I�@!I W��u�"O��1�ϠzL<����G3!��H3"OڼI��>0�~Tau���d�'"O�� �L��l�4�sĮ+�j���"O�3ы�q�����mA�Y���"O�p �#��u�6����	�F2T	[�"O�5kW���2��PƦ�,ߐ`�r"Om���=D����3�:"kN"p"O����"	 �p�rq��&"]��(""O�	�DزJ+h�y�� �|:�ػ"O���Q�E+X<�4��nu��lh6"O��*wK��`1lp�mĊ\�&�Xg"O�1A�aG7jذ�I��^�)x֠1"Op�0�����`��WEJzL0�"O�Q�E.�+B,�ɡDZ�='���"O� C˳et~%���!��s$"O��R�@��^:>izL]�����"O���t��s'��ñS��@
D^!��#%�x��,���)�p��/$Q!����(PIܽ������ r=!���`��Y	M�;�|��E
٣aC!�dʤ0*P�S����ȑ�w�H;8!�O,jN�Y2���+������*!��X�#6��#	!�0;!,W�N�!���<�;��C�4
!ꁶj!����yy�e�&S����	�W���"`3(a��2�>&24"
�M`"�T���H��_E��p��LF̓E��t���4��I$l��ьV�F-n��t 
��
�'�X�X���	ǹs�d������0�C�����Q�"}�#"N�@�D��ŁЫg�
W��B?I��;�͙�O��P�hN�^��P���)��Ӝ}���G�n�,�##�V"r����=�����'#���bA�L@>�S3�ğ>w��O��D0�)�S�^��C�,�l�`y��R�V�*�Iʟd�?E�4�h��k�c��=8j��3���B�	��Izb�W�`1�p����>W�HB�
��px��U�9�:�� -��C�	�+����%�nt	�`�4!��,h���!��S�O�ʖ�B�(��a�) �P� �4Rذ���F��S���i�T���甇d���ʈ;3>H���'�>�Dy��iu��yis㊠j���7��$t_��7��66qOL���2d��H�'7�p��
�>�%��x���<����I���M���>q��i�'eQ�7�	�9��d˼)�@�S�π ��a*Tq�JZ�(մZ�YР�i1N����C*���O�?�x�� �G�ݪ'�J}[����?q�!�-��Gs>1)�(�)[�t���E��H۶Q�m|�;u��h�V�O�c?U�����h�8i�f�w�P���K¹!x�'�a{r
[�L����F+)�!��F@��VP�<�~�������RA��-!�@�d�Kr}ҦЊ�O�>����C4-\�t���ՏX8}����k>@����!K�\�(�� 7@���Ѓu%�C�I]
��7��XB��"%�v�C䉂���%�>TH�݈@�οSPRC��!΂�����MB�a[ƢE�$C�I�|�ԡ�"�_�s�%I��ɥJ�C�	u%�E���ԆB�l	�T�ܕ8E�B�o��	!�k�����J�-͒�!g"O� q�ˀ8d�2�W�'��[r"O
��b/ڬU������r���yC"OdQ��l-ǎ�;Vm�b��"O������Q��x����.��`� "OR!�e�@�k4V@ ��s���"O�<[vb�������'�3X�6�õ"O��I]b��$�Q�F�#��- c"O,��W� �R;��[���,9��}��"O�����u��a{��˔$����"O�l�B�[wʠ9q�'�6L�U{ "O��t�'g�m�`��/�2��g"Ol��5gR+D� �����|��"O8	��Y@֚s�}�l���"O��� iK�}��#T!Q,�T�"OV1��K���Q�c�?qyY5"O�q���K��F�ѕ+�rPl�"O���e�Č���r�
���"O<�	�
��
�`��(5�a��"O ɫ���A&P���WlF���"O9�`k�<e<�e��64�9�"O�I�!k1406�J0��n{�"OM�fˑ����q�/NYxL`k"O<�3T"���Z�m	T��X"Of�rw蓡y���m�2�� �"Ov����+N��L��,��+�^XA�"O�`���ӏf>�jC�E Ke"�b"O<A���,T�*5q��C��4$��"OĬA!��$2��d�[���Ӥ"OJ�We�o~m� MU��q&"O0��'��4`���	B�p"O8��FN�m�r����"��q"O�H'I�LǎΟ���`7"O�q6/�"~��#�l�*A|��6"O>4`�g�2Jɒ����
\aP���"O��)p��#NF�͠���eP<�ʦ"O� �#7u<�z3i[�Nih�"OإyrO�!>\F̓0�/6�`�"O���D#��rb$J�n��e ��"O���).6�3m���ف"O(��4�� �@��!P��Ek�"O����np$�dcJ�;���"O�ɠ/Iq���paZ0��@��"O���ɘ&����ETZ�Z��U"Ot�����&M��� ��%��U�`"O
Y;G�ɖx�L�2N�|�*�"O
a+��	(rz � I�Z�@"O 3��^�R��q�䡙:Z��4PV"Op�؄�Y"`�xmH ��>����T"Of�eC%P8��xaǕ�H�<%A"O�ђj��0��!�$M�J�6Uل"O� lQ�ńoh�rUn�5{�[�"O��pw̍",/Z�Ru*K�0���"O�ܻ�&	��)��K��iz��U"O}��Ė�2����1K[*J��x��"O�1����x?�y`��\�1�M�0"OlA�jɅM���ׇݺr"�K"O4�����,ZP���eȾa��mpW"O�����bsV�(uI�5���"O�z���	?��l a+��;��:�"OdH���{3``P�+�8N׆��"O>|x�J[�`����VC��j �+D��PDE<Q$��.�3qq���C+D�,hA��?h����Pd�0*��p��@'D�$�ԦU6H�Ai�嚊'�D��B&D�4���2i>�-����h��b�.D�h�TM�%L�����-��pߘ����+D��2%�·"{�; 揤d��ERa�.D�!&ő9Y�b��UG8���#�,򓩨� �⃣]'&�]X�E+MͰ�(�"O��ꁫ�7�� ��䔴��
q"Ov������i��d{��πT�(ۅ"O� H0�B6��u�b�:r�a	"O퐡N���t#\�pkrձ�"O��3F����	��/Z�HN&iC�"O��AQ
2>c��`�n؛zKv��"O���N^Hn�U�*q˖"O6�rA(N�G�h�AÌ��"�<,a�"O s� �
 s����8"�"O�=S���eǢ9�$�4gq��B�"O��Ѡ��i,�3Q+�	;>"�s"OH�
զڭp].`d��"z,�"O��h�HÏ6$8����N��"O���ׁC ThE<0=�&"O�I뵎G?{j��4�13��(��"O��QI�ꌻ�	��q���#"O����1DݪU�aI�7��Mc"O��#�I0a��E:�'0��59�"O�(�B�5u���4�G�ΠS�"O�9t��/�LL���K�h�"O����m܀�`��o�&�&L�"O������9H`����iRD1:"O�-��k٥|�HY�T,ΧZi���"Ob*�j�3���cHW�RZV���"O��a5��,f�����3Q����"Oҁ"f��q`�`'HP|�"O
���K�B�nh)�&J�($s0"Oj=�t�\:��J1� ����"O��$iþ8״Tf#�O�T9�"Od8G��D$6�2�'چ��	��"OΌ`�@Ѧ\Z���B�o���2"O�L����*2���咆8 |�$"O�\�0���31��
F��6���"O,�ySL��@�����fA�|2	
�"Obȋ&l��:\�����6(pM�'"O���s�$jDB��ׂ	3~L.�yB��R��h� �1x@��EF��y2)#Oq���a������N;�yR%YpЉ�Rb�q^��*�1�y�KCC^�a�3k�QҜ��WI!�y�(���� d�96�Z�zw�C�y2�|�����N @��hH���yR��N�L�y�B��.��y9��%�yR��4��L�ĨʸQ���S�	��y�cO�Ll�+pW��d �H���y
� �	�u!�8N*��ӑ�î^��1�"O�����:���"23�VAA�"O�A�����gp�YJ��׭�v�҅"O>�a��E�|�Pp�jΓi�(J�"O��Rv�/P"j�(7
�4�X�V"O̝y2K�S�$���è$lH�1"O���CJ_�#0Z�t�I�n�dT2A"O���j%yKP��I���+"O�A�3�K �)UJ�(�3"O( ���5A�2i"RkRR�Z�"O:\�F�Ȣ;����u�L#�"O�*�)�4���q-A=�LA"OR�K�I9z��AÔ
O'@XU"O*�c�*B�~��y��L!Ў1��"O*@1U�\�?f�	`c��Ƽ ��"O���I��S�PU���*�fɺ3"O����O0�%�;�LY%D��y��֭>bh�[A�ށ%�>達���y�'ܛ*؞�T�h��@��\7�yҧ�3��#Ѯ�:Li��QcBR��y� ��kC~ �JW�>lflX�iG�y"�՛W�\�F�[0��<)Ɩ�y�͉�D��v̚�6?�8fE�y�E�f�&|z��U�+�8\Kƭ�yꜻ4̌!��P:�X�Yd���yr��	|>>�z�N0)Ҷ�����y�VW�0=��)�&R(��GM�yra�&3��p�ӑ�hY��D7�yb��0 %. :���%4��u@2�S&�y��թ�~� �@L�)��Ik!矼�y�D('�dQ���	S�V;F`���y��QK��E�k�NhbݲUDC��y�K�|����.�?��I(f�]��y"@�>����Ӣ��4S����;�y�m�8�U`�N�	4%�yB	�i98��c""l8x�3bR"�y�	�s�0���1T�&�s�2�y�Ȟ�$`�t˒��c+0y/�2�y�k̾w�u���Ǉ*��ظ���yR� (X��#���IH���6�y2��'Of*���"(��񻥊��y�뚿1C�
�*��p�Λ��y" P\a9c���ş*t��y�ȓMB��UM:2�r���Q)Gr̄��}rˑ�5��r˖�o��I�ȓJh%`���g�D���B��jVfm�ȓL���UG�M�����b��D	ʥ�ȓ!xHXB��6A�"l`D�%j?���ȓ3�^��&�̊��lB!�]�>*p��!P�&Y6l�r��AF#Pz���\����"�4F �A�g�%sj��� 6�B��˻ �.�!�k$��ȓ�4��vC��n�۠�ӏ/�.��A�ᐳo3Yu����T�\�ȓ]8� �:0L����\:cF�ȓQ��iV�ָ��R��� `T��Q]�{3+�.M�(��*��Q�ȓ � -3�l�4p�,�iP*�T0��k�L���Y�Dl��!�*�9	�';�X	4�O{�|�YBb+	�Pm3�' �y��YN��i`Q`H�z��=�
�'+�%�B���/83"��mo�=�	�'SX�3g-�� ����cC,1R�s�'8lTq��۩t��mц̅�H58��� b5��H?B��9�@�A#	>
�A"O@�(���%KS�]��lV�=�btPq"OV��(R�5��h�I��Vt���`"O�y"��R�c�(03�[�^g�噣"O�% �$�,4fꝰ�cˌ�>0�7"O6Q��U&�������q�\I��"O���/2�	�C��.^�F��U"O�(�L�26ez����I��b��f"O��bGA�9b� `��v�Ԣ�"Ox��f/�>V��T�U�q���"O����<El	�T/�3)�l�!�"O���f%����v��e�@M�"OR��U 
  �   /   Ĵ���	��Z,ۇ� 6v���C���NNT�D��e�2Tx��ƕ	#��4"�V���D�az�m��@b(�BGƛ�O�}�'Kf{�<0F撃Wf���T���M[�ڦ��Wl���\w~���%�ORU(U��R�H��$�|`��t�о\��,����2��$ã�&�S�i�s��A�E��3�$g�옃3	Sb�#fL�`�RI�-O�XR���G�Q��R�k�(�<=��d��>���'
��a�QUDx��R�w<�Q� A��ēH]��K!�ħ!̢9
��A?�9�qU*iH�pR��B�z�O���D�M��'Aй��ꅰB��|�4@���M^�,X��^����c��TJ�!���F�*��)�I��I��ʙ����{!Ä�o���I�+A��堈1���D�IKVd9@��[���� A*�l���;�V�(�2�\�%>j�;ε?�?���p��<���o��tR���6V��1`F��Ȓ��$�aC��x��a��[4'>M2P���
���ӡM��O�6B!��0q됈��$}�4�������	@����C( )|\���U�X�u9sǁ7>�I����<����9:u.�SB5��<bd�<�]:��϶KV�x�i�=_L�/�R��@ˌG��dS�<�a�Xd�G �)�p�r��(X&��1V�'$cцZw}��]�<�D�2��	4@�aA�(����K�F0�V��/��b��,Y8Q�` f�{��#i��ɥ��	iJ�'��P ����H�VmQ�+ӗQwɃ�'�޸ExB#d�ɜ����d��VP��A+�H��4f�mB�ٻF��!�q��:BT{�H��댥��Z��$���?���D;X"и���:a������	o�9�R�0��!z��ycҒx2J�&5��5F����U�s�@-�TRb%���,K9�c$I�����s�@�t���R6�G7�`��D��y�&ϡs d  ��&�2�
�Z�\�J\kEF/D�X�1I؏+��(aVe�b �k�n-D�����67�|�B�������� ,D�� �)�����F$�u��AZ�"O���0Zu���2E�[�k�"O`Q��\�pJ�����2�'"Oj=SDja2<��i�Yۀ�A"O�i���#G:��sOG� /!"O�M�RJ��ebV� �E@3��� �     �  �    @)  "1  �9  @  pF  �L  S  GY  �_  �e  l  Qr  �x  �~  �  ]�  ��  �  $�  h�  ת  �  ķ  N�  ��  ��  )�  k�  ��  3�  w�  ��   Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�� |d��"O
`�(�;���8���-0��1%"Oj4��ND^[��"3/9�0|H�"OB���H��*�ʞRy=a"O�味V�!X��!&F�:J�$���"O,��a
���C�Ą�M�"O,$3%o�-���p���+Ն�:1"O��ݢ1����`���y14]2��i�<�6��{_���c�H�`�fX�$Kn�<��A̼VI�xR[�)�Ć�pඤ�ȓA5��('nߡ4�� �)˩%� ���,��r�؊b#`T�eT09���ȓ!�b��g��}�8�F��-? �ȓ
K|m�ș�VṔ���2�%�ȓ"R�X�j�4JN�1�˘X�i����̹	_�jZ��1!g��zܶ��ȓgil,*�J�
j�Ne��i�J%b���f	�(U��:���G��$Y^م�~r�� S�%T"���k\�jx�ȓ|4�1�îJb��@ӵ�ݩn�V��/[`�"�v4�R�!ʎ<��M�ȓ`:��z�ؚh�J�Z��$HY:	��H��p�m�C1��!��B:��0��EnjZA V;9����J[
2���	��4'J�EA�IVW&��~�(aZ��ӹ�>� o�Y�|�ȓ�f�A�
Ο7�H��M�$�����mޠP����/���ANXo*�ȓTv�����{ ��-7�*h��I��sB�8�8���3����ȓNe*M�悡;������X�o��!�ȓ'lj�#F�m�+R&;�|��2)n�C��0S4���T:
b���:�0!��e֊��)��ͷV��,�ȓ0�&�8#���� ع�L�����;�P�AFd���,w�0dFz��'��܈���h��;�3W�����'���tą'i�\�	DkI�.0��'�1CeKY�R�	T��L���'7I36(�z�R�`r�;X�xt�
�'U�9�.ӽR�p�Ph�Oh	#
�'� ��nS�8�H8���ƗNG�q��'�n]1f��+w��A1�F�)E�pa�{��)�)Ƀa:Ԩ@E�'a��Y�1�!�ę�'פ���Q�֩
e 8�!�$��S��
ce�p�-��bT�k�!��j�x��4����sB���!��(3��pv��/ %2�ږ �5�!��D�Fv|�)v����t��@�'�!�ݮ*H����H�[8��Aw����!��Q�Zt�	�"Z	���\�b�ab�O� ƭW����G���1"Oؕ��DْvO��l�ץ˴�hO�#=��O �b�Y&|Шe�1(^0o|@��'@HqGR`�90 MH%hdh��)O�=E�īơ;�@e�u�E�	�-A����yrߝ|N���W�7� KU��m�j�D"�|&��A3%�G���Y�"R6Dp���#�Oj�i2����'L�40�	���<�r��Of��9lO¼;b��&��9Z��E�NvyI��	ӟ`�=A�O�H@��h�.`(r7m
��Q	�'�R�؅͚#-�pr��ܾԝ���� <1�q�G?$L�m�S&�v�&�Q�"ON�0�FȢu��󣚢>�j��֒|��)�S(iѼ��#�Zz��;5�C�I�3�M���� �H�c�!�|�TB�I�	֜���d�Є���]?tZzB䉚��
�
&a/�8±�]�2�LB䉧r��t�u�T����J�ȫ<Lf�=�ÓN�n�뀃ݶL8� :p-��F�Z��ȓxN-���t��5�E�_XzB創)=Iq�����NGfh�ȓC(�� ���	Nَ9�'և*��9��)��X�.k5@MS�CF+t�x�ۢ�+D��!�.1
�NP(G�7���פ)D�\y���w�
�:��@)>j�s�@'D�X�ꉂ���2"�_x�ա�)&D�s��ޕc8L�G���t3�̛�f�OzC�	�M���7$��K]�v$I������<�@�.V�-9q���pqlO}�<i$�@�V��TgF=INܛc*ph<�C¶y���G��%TY��x�d��yRgA	��iIr/�^��HS�B8uP�=%?I$��Y��	�bV����S/a=�!�`"D�X2�Î�oT&UJtL�(]Q�	{�M����	�_<�2�A]�\�����h+��C�ɅX��ec!_�1M�'$X���C�	7 \��#��2�����Z�
SN���<2.ނG�=*����:�|�!�[{�<���խ_>Q@wb��tY*ѫ$��@�<�2fF�\`� SII&qz�%	d/�t�<�"�D�A>e���H �����d�IA}���(�	�g��UcM�(DҔ*OD�>E�B�ɠk<����9.�,�����D�.B䉃�2X�!�I�DϺ��`�+N�4��$*ʓ"u�a���|A8�coʽj?�P��F<	5DXSV��"��<V� U�7�RB����<�©�3S�x�Kڷ2�H����y�<��g0B��1bpU?`P�5��)Y��$����'��SL�g?YsA,Lϒp �� �EL�0#Zi�<��c�y"��bfDx�&򱊝h?�	�f��+�1dr�(v�Ǟqs�	���)�'4#�#Ho�����#,����'�N0�DO�3�����"��Z$
�'(����Y̔3��>%��"	�'���(�ٗ~x�;"��5q$-
�'X>��Q(�6|i�9��E(p�\ �	�'�ih�FG�+�[��̧`Z��'�>	����2���!AfM�Vn�z�'��pq@)�,�J$[��-&��S�'��	�&�^���Pr׍�=kֺ���'-Ё�)�p��q蒫8�ؘ1�'��A���U%�f����������'���9�B�,P=l�O�$��R�'���b��t��� �jZK�t��'p5a&MM&7���{�hYJ�*��'W^�pSlEr������ؠw�X�'������:H��|�f�n�
�'8���	D	' D����P�FL�	�'@L�AR�n}(r��ގ5�8��'=��uD\�P0�	��EB�7�(i �'O&������m⬱��6�
1�'�f|�E��b�L�ȴ앇]+Fp��'���*��s�2�	�o.|��'�֜8#Ι-�\�xf-��~̀-�'_��$/Nn�(y�5�^���+��� 4�F�n��귩N/IF�"Oh��$&փ{,��Q��0h�� %"O��
�D�?J	�#_�:���g"Ol�� �%8{๺ ""���{U"O
X@�M!ib�;`��'�� �"O�Xz3G�$t��DQpʟ/ݤ1�"O8��  G;r�I�[�*��TbC"O�4�≁��T���OE��"w"O���	+f�2Fb��.��R"O8T��_�W��z���YA$��"O�Y{���R�s!�E�)�\x�"Ot/O?,J�m�r�|�$"O�0d��f��$kǫ��p��`�"Oh���h��Ju��8H�"O��
����V�DP� '
)��,�"O:x��+Z)J�q��L�@� "O*��$�G#BD��Qf��&�����"O>0������ ���e��@�$"On�)@�A;~;@������B���"O
)����+F�|`{"�(
��af"Ot�Kf+ �~hPG˭O6|)�"O����"�d���G)v&�)��"OԁQ7/�2#f֍б�˩D�	S"OT�i�ˣP�*��$eW�"Q�5��"OȌ�����8�P�	�c�?�]�����y�B�K@��7*�2��3�ȕ`'����G�Z!H�kC"h�L0��V�j��!��Xj��G���dm
��%�-$��ȓ!;vؒ��X�O�d\#�(�4s!���ȓo�-�W ��& [�+�n'��ȓp��5`�E�,ut<I����/]�ȓi�����X�@5!�B(�.%�����Yb
�m�|M��mY'f�7D�TBA�Ĕ%$����X\���uC<D�Pۆ �0��i0��ק2�����6T�PxF� Q"�Cg��09�P	�"O~<`�L�5�ꐣ���$�N�{�"O�ѲI���j�i��Cr�tQ4"O��@�Oվ@��d�B� �g�Ĉ""O0�Ґ�-A_�%9W[S=4U9�"Ov���'�Yuj�B�%�e*4xh�"O���a]�C����N�i\a��"O�`z���ì��n(T	L1�"OZ�S�[�'��la˜nI	��"Ofܑ4�B�xS@,	�jY	��p;1"O�-���� 4;�GU�q�.H��"OL)��M`���C*� "O�t!���~��Bg�%'t�Xi1"On�J�L�9^WV�E��
]��"O�X�c"@:T�
�K���l��y��"O�4���Z�&�L#�C�rz�`p"O�d8���l�h��R��煐��!��զ(n�iҲ�� �|�0�,(r!�d�m��c��L��,� e@KT!��8[�i��L!N���3%���]#!�D�]'�d�ì�:%FQ�� ��X�!�dH�XA��V�(R#��)�!�M��X�;e��@��"c��i!�Ď�=P� (�FZ�
��pCBL�@�!�D�#_�L�B��/E��I��Kт�!��C4DDޔ��/� \�:�iWǗ<�!��C }�9G�9�����є%�!�ăx$Y�������Å�p�<��Zzn�� �`/�; &Xm�<� Pс1�L8Lq�a�&+[�f	���"O�$ s�/@$�1E�Y�V�,ũP"Oȁ!7,��c��8���]a�D�"O�+�(U<hBJ���y: �p"O�	��W'��sGFP>1�'�R�'c��'v��'5��'��'老1E��T�� �m�{;T@���'B�'��'ZR�'���'?"�'Z�J3��B���h�Am�dq:��'%��'-��'Yb�'�R�'���'� ���j5(��3�����i,k	B�'�"�'���'�R�'�r�'�KԺn�V�6g��P�4�O=>m��'��'���'�R�'���'gr
G?  t�!8��E�QB� <�'��' ��'%�'���'6�ݗ~<Z����?�d���&,2�'��'>��'��'��'&Ҡ�&�	�BlՖs���9��ϚH���'�2�'�2�'<"�'�b�'�r�Zv:z�0t�ʂc�D��s���R�'jb�'�R�'��'K��'��L�[�Zk3��%w9dlq�L����'�"�'���'�R�'/R�'�2o

0�á�2A4z���
��@�R�'w��'���'0��'b�'��CYi��U���XX��DE_o�'���'Q��'���'��'e�jZ2>���ۓ+Q� u��a@$ b�'���'��'�r�'�6��O�����t\Ɋ��ѣ
Ԕ�`��יd��-�'�rR�b>�49���� Is�a�[b�R�/���>���M�g~� |���s���I8f�9�&ZQ��()7��#۲���՟�Ӧ#�ԦY�'Z�)��?ɤ���ZiϮk��������0����O��h���׫ƊFw�ڂ�Q���I`A�֦X�N/�Ia��!��w�V��+eh��A��8�ƈ���'��7OL�S�')��޴�yr��0.N�a�@@0b��T��0�y"4O �	].ў�͟H��
Ypΰ�DB�2T~T���~��'��'f$7�$"�1O��ʇ��hX��Ε�K�<u��.�	����O��dw��'���J� HA��I��(c�*�b�O���11�\U%�]��?%h�OzY�2o;;�\�q��T� ~l ��<y-On��s��Q��CB�p$����!��(cHa�L ݴ<6�`�'��7M"�i>:`�aHʌ�A��& ��IRz����ȟ8�IC�,}n�T~"8������B ;##K�^hP���� ������J�	AV ��'���AV�[y�g�I�Hk�!�O�gM��hE`̵βC�	#���.�uz Q����j-�b��-�be�a�_��K�M$��i���P�R�♵~���P��v�����]�o��0C0GQ=QT��7s���5�6g,��5��B�"�SV�Cǰ��ET7E7$�Ke��79�`��%)ɶX�4��6L]�6��"�Y `�j�z����k0�7M�Ot��O��	�z~R�h@���`f(��b�=cE�D�'�rO�� ��Od�9O*�$
�u%� ��!F�z�4L�i�:u��m�C:*�s޴�?��?1�'͉��t ��|���Z�G�2(�`t��Yk�6-�7c����3�ϟdҖO�c��`=�p��� �M���?Y�ՠ���x�Oy��'�>i��i�>Ĵ�1��>_�P�;`ag�.�$�O���P?"��O��'��'�,K#��`�XZ���'��p3Vd`����ƀdfb1&���I՟�&�֘&�����[-R�N�{Bdے/'�7��O�<#D��O����O2���O��'�?Af�>a�n��o��.���k��Q� �~���x��' ��'�'!�n��G50dk\�7�r���/�1y��p�y��'���'��ɝ\K�AH�Oe�pqDkŒJ��f���(�~ŁO<a����?i��eۺ!�'
��c!*��2�{CdݝX�tm��O����O��D�<�&̃l�O�X0	E�,c5��yCo�)]�|<�a}Ӫ���O�O���9V1���^8}�  �Z�z�X&A���Mk��?	-O�Ȋ��\�ȟ�8�q��# ��FM��O�F�N<����?��N��?����?)L?AS$
K4J��)B/��i�at�F���O
=s3cY����\�$��f8�'�1�0�o1X<��B�	i�^tѯO2��J�bL�8�3��A40#�C��RC�lG0F����dyz��i#��'��Og�O�	P��|�q���S�����gZ؁o"�n �Iʟ��I�����k�t[>�C��(|�`'!Ƨ5�VE�f�P��M[��?A��V:�)"+O�{����2��/'�*E���M�b�H48O<���7lLa���'$��Ĵ�rAC�^�^�� �g�(O����'�L�B�[���<���'H��0��rՏD�}�F�e��M��>d1AM>����?!����e��H��$��#�}c^q�lP��#R��'���'��'��ɺ,� i��T'S�)AW���[�
�0c͟T�'���'B]���$ѱ��ć�Cfl!0�� @�)������d�O���Od��?��/0�����Ժ�͉/�F ��FUd���R�P�p�����by"��&���)K���, ���i"�[xt�q�����}�Iٟp�'>��'R��6�'��'~ƪ��f��E�4`��%n��$o��L��Fy��ݨe=��6���k�51�J���_�8�\YS�&��6V��������!cӟ�$?=�s�� ܵd�R�x{��M++�dd��oSV~g�V-�-	��1���	$Tj�x�7E�d�]�ŧŞq�!�O�\�p ���?xlP�'ˣ#��d���5l�a"7Am�l���L-L�6���e)l/<�%έ?���b��6z���C�̘�b��0b�7r��4N�%R��9��?^)��� V�,����ǒ�2�`�9n�|Uµ���J�%��#G+.1���G@v�aGo�O(���'\!8P"�$�O4���O�į;�?��L�L�[���gLM1��c���G�'h$@[ńܜt���)LpF{r◯V���C������m��_I��D��@��JpID1E�T����hOԼa�� ��58# I�"U�h�&�O0��'��{�'��v���&��vҰ�R*�%�ybU�KĸB�%U�:̀�P��R�U	�"=ͧ��M�PS��iAx8!1�K'F���b*׈"! ���')�'�ү���D�'��I��B�9sc
 ����[FE���r% �4��A큰9$p��d���h3
���P��C;B��0� � %.���.B�n��;�'�(��?�T̃�A���T2&2��;���?	�����O���'�2h��N Iڄ����ȓ7	8,å�/N��RI�$)f��Γ*%���'0剌2��m!ٴ�?����XB*Nu�S)6S����֧;7��q���O��OJ�
0�C0����L.e��)㖀`���Ƃ�v�i5�2o��d�N]�(OZ����F�º})g*��[�d��Ȱ~�R/�i Ɓ����(e�$����_�'����b�>�z�Ő5}:&8qs���i�5u�3D���� �5\��];V����� ���;�O: '�عeeE�(�PYC��`�*݉��y�l2���M#���?�*��}�e��O����ON�h&�h�P�ӕ]�L}����Q��q��	&]:ū�%�7;�5K^�_�Rb>��ȪU�y���K�>��@������#�+��(�T�1�Aԑc���#'E�U����b��wD��"��AM�	�Nʂ)w&�9A�K)b~�,���O�I�f�U��\+���M!0|�b"Onh ������@���w<��q�I��HO���OP��%j�@a�+�3T7��  +�O���5���1C�O ���O0�����Ӽ+��9SJ�y���(S(X9%��t.M� �D��"��Q�F�g�hi�'
J ,я}2`�:@>�����MRjPi"���
#>:g�ߩ�&���c
��H��O���QF��K�*�96�

f��Ro��A��DϰaR��'�V� !<P�*�*�NZ�l��M/D� S���m� U��aA�6����%ۍ�HO�)+�$V�w�-n�URJ!�a%�x��2%� �R��Iʟ@��ڟآ��͟��	�|����4h�P�f"�<�X� 6J/=[�,Kd���A�,�d�鉳TB\qK�TH/��@���/��miJ�16y\9E�� ur����<��'A��2�X0���%$р"�L�Z�'�htBClW�`)	�O:N���
�'�r��ĂJ�Y�mPb�"K>eZ�'�V7 �$�-䞩n����D��̡*a�9+�N�")^5��bW�� 4���'Z��'<����'k1O���h�!G� 6���Ss�o��<ɔ�d�O�� ���y��{g�]�6��y���\�w�"�,�'<Z� ����W�M󅌉8=6��ȓ|t��1F�?NF�j�
=����񉬪ēM��@s@G,v��k�e�4."x�$9�ɂg�i���'���y�����՟��I7�d�� B̕H�����3|k�5{S��jܸ����T>Y�|���X�p-�4����ꁁ��<�Fy����N���4M�$y��ˣhپH���p��w�JlKvAM��xᰒ&#s� �A�Nķdb���O�}H��� [bL���^'��,H�"O|y����	� P�%�+��A���	��HO���O:��P��5J;n����̜�&=���O���J*gH�x4I�O.���O���ܺ��Ӽ�"��)��2_s�򂪜T?q�+�Ix�(yQD�{�fZ1�ǧK�8������
�%܊IS���W'I�5�ax�'7�{k�0��y���_��~�l��?�'�'DP% �͐�C�-���d��i��'T�-SC�X�v%��P��A>Z\l�(��&��|*K>��$]:$ʛ��ؑC��U�@��mP���U`Լ:��'��'���s�'�"=� ���ڂ(�@��f��TVH�/Ռ>"Z���k+j1�a��u�`�Ƞ�(O�ۂm�7o}����@��~
,��W '0�l��2y|P-(�!Θ^��yA ��(O�h��'�R7_5F����>(�� ~ !��DzW�=���{��8Q�
�U�!��DM���Gp��`�&��!g���Ϧ�D{��)�m�t$���I�8���A]/)�!�M
�dH�&��:���1�!�� ��`�L�n6���2�z�=��"O�I�jſ�x��ѻ<����"O��@@�e��rS��I@�5)W"O}-+?�ȜY$��Q6H� �"O �NP�/��p�J%z%P�C�"Oƀy��ե8��(�ƌǿMZ��
�'I��''�Q�����V+�&���'�L3���A)R���A]*h1�'ݤ��ѣB'6�8�M� 	,Z�	�'U�{0�R�F���G�^��P	�'�T�`"_023��J׃
�9nY��'	���L�5Z]�4��Ő'`��r�'
�$#��%�l\���>R�̘��'JX3ĭ�_��"wȫO?��'�hi�Q=u��Ma�曕I�&��'����-ں+���xڀ�
�'@N��-�I��aeɁo�V�
�'��Aj���!V_!��E�����"OjMbf���P���e�>�"O�r���	*�����J����"O"��	x#P���ސ�2��!"O�#7�I(U���TEF�����"O���O���u�3^sf�qW"Ox�7�ۗ8�|i#��DȈdX"OV!��%�B(��`� Q0�R�sd"OhEPQ��	oΑh��˄I�0M��"O�)هH�,7�#d^�QĀ�3e"OfT��H�����-������"O�xP!b��1SLu�eN m��W"OԜR��@�h9y �	���!�"O�9���,X�<�t��y6�a"ObP냎X�m�����$X�,�2r"O�4��b5>�nPؤK�P��Y�"ON	�qN,P <Y0�����>!�H8��=y�AW>12���թ ����F�N��xq'I�O:����� ��1����ot�a�9D��#qb#K���{$T&8�<M���:�=��-abA$�'t	��Z0�B�;4�#O�&�X	��~�
@9�]�G�	ɦ1��ΓC]P�y�&+�)�'%�8���D~�
p�dm�O:v ��A;��8�cCG�mJrًP̴>i�a;Z.iQ��N�"&���o�'���f�܂/��U2@�;pa�	�se}�A��!r��څӽ��9� W��HA`���&�2×�s�p����@�J��䘯�h��toT�+譢c��'#�\��HM����?�<�{��.�ԟ�b��J�G��ȣ���kc�)�*O�ZtŕS���RDD[�hig-ьE7�]:C��N�S�TLT7W��ik�w[����1d `a���G�RwZ]�
�'���b�͹U	���"H�_�z�����5���]�2�9QkW3+DL�;�"���(O�Q���
�x(�y�ffԠ{�0���'ְ�A�ǃs#�q�M��q��¸.�2�"N(5K�=z���W� ��!S.ar����I��u���
���H�Z�0�E���X�5"`J�ϋNq��擤'-\ub��֏D'���F�v�B䉭5
��0)KJ}���5㎌8R�XǨ�lS2�����?��1랬x�R睑vb�HH��E�;�[�n�>}/RC���6�YԮߺ7��zeʜ8#.Y	�'/?A�
ҤY�F]��_�b��Y��'�Ls��i�L]�m�Hi�����g�����I+'j�l�BB�U|=�ң�Y���h�%,e5�ѩ��¥)�� ��fȭF�2�PR�	�J��|b���~�����,\�V�ѐ�n.��$I�h����%��,>Lp�֣J������NS�t��$�@Dӑ�(�Y����y�C�
TO�]�%���	���S%��Q�4�B���<����=�O ��Q!���yϔ9�*E��Ť��G�
�xǄ<y�n��ggA�]� 0kF�!`��#�O��� �A�Pj�6MQ3n��coQX�'�`	�Ɉ�"�l�zU��'���(
��[(O�� Wh3La����DF��.(Ru \56E��iFT�$�qI�J8�� mK��%	�p�+g,S�k�\���a�����dCUn��l��i�D�ֺ� '��}�#[7qf�4ie�q�<Y񤚢����m̒h�DӒE�o�ɸeQ8��-����UQ��Q�~b ��oa�Hw�D (H���^l؟Љ��1*S���!E	%�Ly`c�D�~ޤS5��{�R�R�Ǆg�)���@���,1[�͘�(̬��� @�2��d��ve6�Ӗs���.��8E�)�� �>[���49�+�D	�p=�2��8�X��'퇎T*(!��Z}��)�t��'�͢1	��<�'F��9�'�p�3	��'�uiWBH 8��H�"OvUa1ֈJ���S�&@8��i���`��
��~"a��vT��?�q���ɟ�s���'n)n��G�!�ਘ �-�Oؽ�#f��*:����Ǘc8�H
uJ�
ըx�	,�~�NB�bT�ڴj����_ߎ��=!d'�$
����r���
Q�'�$TǸ0���2����8Ԉ��4a�2����w&�U �G�E�b�� ӹ�j zc�M%"a|����'0f��e-/C����ƀ��	+ax���v�d�ZP��K�N�	e?��'ؽ[�%�������A�ei\;�"O�i�6��$��BL�]�HTB!O�.��=CF�Q?Y�'���O܈���c	�
���]}ϞU��BB�)R�i�C�.�����A�dz�<	���:P[��
+z����JX?��'���3w��>ja� ��(V�NT(9�{�G�Z�����V�E�C�Ѳ��O�𐄍�h6,�q��P�lӧ�i�6�2u�]u�4���r�wgCS7�$Sc�_�+�� ��Ij���{�j��+5��1TN���˓E[��C�@�M+0&���<b��u�B���0�&�Gl�H�M_�P=���p"O��pa�>u|���l������i�.�ӣ�����ś`8� 2�S�������s�-� 	��tЈ!�m��.�Z�	�6�,�$2G���W&��*�y�G�?[up�'�*T0�D��?6��BF�}~�e@�B���<�5#��3�� �C�η�0<Y�!O�YA\�� �>2���"Q�έ���á&[6i�4��WH�i�]���_\�d��FC*��=�e%h�"���I�B��DT~���L0
7 ��ٰ����N4`���5m��(�+�4�x�A�	�.!�Ė� �4�J�,��h:"Ȁvrl8�E�!!$��V�T>��pL�Am��]�{Zޑ��C����ɰ�F2�C�I�;��8Z�dE�؜�7,ei�	2�#,}"gHNJ�i`hW8˞�"� ���'��Ĩ�/ wD@2����]YÓ=q �q$Ⱏ �rm		w�*�[���Ɣ��� �drf�>94�\�?(���dӢx@��4�	A��;�H�h��O���5%�'��)�Y�v�	l:������md ̨a%H�ynB��6��5`5� �P� ��(��*�I#��	���S1e�6�P0�
�
�4�bB�68�B��:7L�����3 ����@�?UX�'�"���'���IE^9�2�6a�3a����'��� p��I2\*�Bʜ\9�-(�' j]�t���Wj�xB@F7����'kD� �KHfj��آn�i�b�Z�'�P���� &~�4���.�]^����'��c$Y��|�{Q\�H���i�'w
}��+^�n� L(B�T
Li����'�P`S�J/'XS�P���'7�Т�S�0t���sH�EB����'$r�Y��Kr��̂Ȇ�:y����'3��+B�B%Y����C�'ׂ ;�'V�]��GE�$�R9O��h��'Z����
�I��TGR��9	�'� 8�&�]J������@
`q��'�$t����908,��5NX$�l4��'!�5�'��6U���4oϦ�xٲ
�'���!^'��#f��
�u�
�'��E9@�:\֤I��T�q��Q)�'݌yJ��ɽ�8<PG'n�$�!
�'�,�R�B��� a���RP�<	(ۈ=V�B��\�!�.��.At�<�-�2>�^(���Ň����u�<Iv_�xD�hR�c��D�0p:���s�<��I��^�\qk�'Ҷ$��9��/o�<� jZv)F�@x�P��1O� ��p"Oq���=�PE�ը�'.tƥ�"O���h �"@�P��:
]v	�&"O����#�~��5b��c�R��"Or��K�2S������Z�E��,�"O��{V�?kz���o��l��""O!��ʢFQ�U����B��B"O�%+��L�X���v�V���"O� ����D"HX5fE:9)�G"O�P��iP�HD��e׮c rܙ"O&d�P�ɧ	f�+/��h��"O�t
Z<A�mJ��G�Ye�z5"O����hӏUe��)�L�>@X�+"O4Z@�)^�6��V�M�#��Dq�"O���"+P�j��=��݇f��} �"O~Xq��_f] ��g�������"O�e��	�tU����,�n��c"O@�I @F�B�5m��mK7l �?D!�$�Y�ީڂ^�{t�Q�	7!�$��n���C��׀RV�
JއQ!�D���~8RAg	��T���Y#!��9��"4��c�vmbW"ߪL�!򄎬4�|D�$�e��=�!٦!�䙟4��Mj��D���B�8qb!��Հ�z0�����tĚ`,�6ok!�����8����N��0swK�L}!�dR��F����GŤh��	.f!�G�dy��J��YC��MR�!�ۤr������L␱&e���!򤑞Z���h�=%���ېdO�U�!�$��Y�n\s"d�"e��Q��Тz�!�$�0��lѵC��	�H���/��ms!�d�h{���+_�tɆ�`GJ�wV!��T����v�<���hI!�$�>*-�,�!D��!Y�	O�S�!�$�����bO <P�� ��t!�䎚>Y XJ��s�X�%'0'p!�D�:/��5�,٤Q�F��q���dk!����n���/F�3t�!ӆ\�~!�Nd���R��{g��?p!��E��D�(�gWX�n��D�Nn!�@�;Ȏ� d�B7e�����I�Q!�J	
�0I��٬s�d��ɗ�R!�ę�	��mp@kC�o��-*�E &!򄜲[��d���0����a
)!���"o�ЫҋZl�!g��_�!��f՜Uk0�Q?m�@�3��1Q�!��x9���pC��V��+�P*^�!���9(<���eI"O�4=�u�	�G�!�d�&%����,ԗv�nx�&���v�!���9^������P6z�m�t@I�Y�!��J�e�1�##4\�>РBB[7�!�E�V8.���K%<��B�M:F!�dY�XB�H����4�'Z3o�!��P�>��s�Ľx�v�7@ІS�!��V{Zh�в�(2犘k7�A�!��+H���{�o!zDb�
���q�!��ֆ��9;p	��^Y� ��I�!�D�-`(���%�Q�5?^��Ǯj�!�T�p $��DT-&��I�-�=D�!��͇�X,sE #vqTy�mÎ	�!��
�}���3qa9aDyx�'�M�!�D] n*������#�n)*�#41�!��(oʹ)� 
R*�F�`&��Ux!�� ���m�4 �J��D�W(i����"Oՙ��T�~�X�ئn�&��"O���*�V�����l䶸��"Od#��po�%��ǀ2�j-*0"Oh�A�CE/>;�D��ݑD��i�"O��3��*q�Z�
�̅3{U�lQ�"OX���b����T��ƲBR�ىs"O�!r�M\�S�����C�Y�-��"Oj�S��S�����Z��Q� "OX��� /�~}�1ܮZ�6���"O�s��V�$�tiH����2`x�"Or��1���\Z(@�L:.�jP"O��� ,��Io�P�.�!ƊD��"O��AP�(���U�D��1� "O�e@�,X�wI�%��	:
�젩�"O�XyedG
��Tb�Id��R'"O��	��ݍ2.�)��`A>(k�1�5"O��Y&��6@�T�v�QL$�X�"O�U��n�!xI�@b0l�)hI��!�"O���W*�}@�M��@�)8� �"O��)�hк- d�ұ�:a3,Ġ�"O�-
���#��}���8
+ȝK�"O��%�ܭ$O�\;D�I6� C"O@Ԉ�#�:�@�p�a�-H�"O�)��	(Td�-3paޢ<ƌɓ�"O��L;>��(b�NN�.���Yu"OV5a�"H�dt�&�������"O9���S�Q�̩ a�C�(�"O"�)��^;:�����	(%��d"O�D��*@,((��Y�0�5x�"O�\Q�*�1��H�0���gڄ�r�"Ov�9��X�#�2eb�g;U��9J�"O���7C�5~vl�rfހ��u�3"O�e	&��w���E��w�^<S�"O��S��'c�0���/	���D;�"O�qp�+D�z46��UoH&9��ͳ�"O��Td@�8L�:ϙ�%���+�"OD���F����VKU#(B ��"O���e/T	{�F�x	�)z�&Հ"O���A�1�r)��g͒��|��"O�p�տm�@e��K)����"Oƈ𰀁�BO����E �xlKB"O>`	�-;!�TY�7kڵU�X�y�"O�Ux�d�o7��qd����L	""Oµ�!m	@wP�jF�ͩx�퓁"O��
U'����)�0&p��7"O�@K�(��5f�v?uP��А�(���3Q2��9 ��'���'��TC�	^��}àC��N&lX���fnC�ɸ>Μ��,H41Cа��i��c|2C䉼w��-��Ag�Z���JG5`C�I�EH���!�4}Nm@rh��;$ B�IwsH1�9e��@"�/%�PC�IA*�-�2�۳m�4D�§�C䉈cT���lJ�$x�c������F{J?�8��ӹHh@T;���nY@�S�h+D��05�D9ZHl�l�*7�j�i��(�hO��3c��*�1�t5x�ヿU�C�	7i1���]�~�j�R�/B (7FC�	�ⴁi�g�YB�Rf����TB��$D�wӓ�k�]1kVnC�ɜTô�	@%*�����I��H�v��D%�7���S�F2�����Y
��C��hܚؠ���E�M�`�A��#=��S�? f9��1.���se\��I��"O���U�K!DC��GÚW�z(�f"O��p��I S���v�J��(� "O��"��t14p.Ihl��F��1�yr�]�J�Ua��ΩK��K�`Y+�y"΅?e���K]��%B%���y��Ku��A��Oٚ~kf��(�*�yÅ0d���� �-�����A;�y���P洬��,ˆ"����`h�y2��S�|�y�E�o�p"@̄�yB�20�����>ce y�p
��y���<Lbڕ�� Z���[!�Ӿ��0�S�O�H��-�mS"�aBJ�Y3L��'���{��<MM�	g�i\@#�'Cv�k4j�	1����+D�s��x��'aƠ�D_!Ex��C�u����'����kQ=�l�b�K�JY��'����L��"pb� c�a+�')����+�.B/�Y��˨�~	X�'��))d&��r�b	�a��k٢�
�'�(��w��@�:�bښh�"U�
�'h�-�u/w8!��c�Z�"	�'�X4赩��Z�)�C%M���	�'>B8��	8��u Ĕ5p��	�'��Ԏء�ar���pz�r�{2�'*v��TP�4��<a����Pc�0��'�R@��K��3t� *��ȁKw��1
�'���w�iL|�qB\���� �'�L!��R�]����q��Di���
�'�q �#��x��t��&��Hڔ��'xP�&Hǳ~���;�J�%X`b0@�'���B��N
�i�JgX��'I��b�k2����֤ш?e䝋��2�S�TI7x�V #ŉE!vS��Z��	��y:Zt��d�S+j��补I��y"M�m>̨kF�d���ŋ���xR�
[�IÓFB-� ��&��?Wj!򄇐/X��kCM�y~�'�~ֵ���d?iłǠ8�(�`m�5��I�&�
}�<��ĕ�Ȅ+T��3M+�
��d�<�2��,K\t5T-\޴����d�<)�M��6��"3).RR�`�<p��0T &���E)1��
�HMZ�<GNI+,��]��(�^�* ���T[�<aT�q�e����Ԭ��l�<�1ɂW��x�d	V�Wx�����~�<��I\�Y�Ɣ�5��,	��+���{�<)�	
R��EY$%Kf-tm�ċ�u�<9�O�v�� G�'2Ĵc�Vu�<���ηYA�H�$�
 Iw��p�<�2���4��!�CP�6mȲ��i�<ADc�`�>L�&,U=�L`�P\�<��e��Q�
X��c�M�Nݳ��L�<��)D�1.ƵQ�a��q?�]�HJ�<)�AȇeD�L*����
��l��!I�<т�,O}h��@!�|4�1#I�<��H\#�Q�bN�ɼ�&��F�<�-���%���Q��Aa
[E�<��ٵ�2`)2ីO��pt{�<�Ȟ?z8��b�2=ylؑ��^�<�0L(>��,���Qf��\�<)4 of\����,��KT�<�q��/3T���R1K-8�Y���Q�<��E�!m�>���-��]�<(�b�i�<� ��zQ�H"}�K@�	6 K�"O�[%�0p��j%�ك3,YH�"OP8H�kK�t2�A�2�Y�B+��"Or�f〛ep��f�L��S�"O�=�@N�-��Y[�Ê�uK:�*�"O��>���AR%��q9�Q#"O��9�\�/&�RŅ!rhx��"O(���J�ZVt�E\�e�"-
U"O��be޵/��x��Y�\]�"O��
�+c�1�B;�`�{U"O���Ǌ��@�f�	G��� �l��f"O�1Ƞ� �K��`M����"O& ���������.I��"O�h(V��(�gP�b5���"O����	>�����=<Иu��"O6�Q1���3�����LU��$�1 "O��pgaS�
��3aR�v��0�"O��P�D��\X \@boV���k�"OX���G�Uw ��C�E ��8C"O~���.��x<h8@@K�m�n��$"OV���X�$+�8V�y9��d��'�0T1�!]N�Y��☇`��k�'�V-A#��"
}^<
��I1C���'�r�1��ɀtHޕ�1m�,uĘ�
�'�X�h8	����a�A�&�x���'��|�gⓌp<(�Aö%lč��' ���Ǣe�h�)���'q���5��4b��I`˘)B�@:
�'�(���!�>4�a�H�����'?FU��i�/�����d�`	�'S^��
�.�l�[S-����'��93�hZ�vڐ@p.��|���z�'8�pzw�N'<m��8�oTsqJDA�'��8 9*�4�(�\pvy��'7�ݘ�EA�a�0�I����	T�i�'�PC#��8f���30�
2	X U��'�|@C�gE�A���W�	�
���'^>A��(ѪI(�Y��E�UY �Y�'��D�E�F�l��B�J�^��'���t��h�۰�R gΨm�ȓTE�)
�\*W��x��b�$xrv �ȓT��݉�JϲP2��p	G!A�"��ȓ<�Zip@g_ R���0���JFt8�ȓ(�Ʃ����8v��� ���ȓY&�U  �bn p�D���$5D�$��;8��y��ꈚ=���2��?D���%	Ѓ}$��@ Z�u;�l��D*D���Cm��A� ����54̕���4D�\�0N
* ��x0aפ9�I9P0D��A�`Z����e��b����/D���3�ߞH)�R�4�hi���8D�L��f�
KXث"���`�X1��#D��*a�B 0I
���$&Pu���;D�8(a!��)��9����"1�E��f8D�$r�V^F�xQ�菒#~�U�6D�d�2왦)X	z��*Ҭ�Æ�?D������ak�-
BJ7\�|[�f>D�Hу�;8^�yR*G[B1�t'D��˒��}o��Ф�:lM��%D������g�diړ�ڹc�����D)D�XHb �
J8Q��.���V�4D��Z� Ő<�B�
d5'4��"@1D�D��T�-vD�:�f�E�@=���0D�|*�-0tR�� �	uI��e-D�� H����1�)�1�[�l��6"Ovqb�¿H��������Qf��se"O��B�+e�^<�b�߭$_ j2"O6�8�a_�#M��S�Ką Z\���"Op/M!�*MU�R�Y��Q��y_5X�
���B(H�:*b���y ֔Qr0Mk��U9P�b���y�-T�.^05.Z7WX����,�/�y�)[�'� =Yd�V>���#U=�yr�K�Y�jw���9n��+���y�dB.*�	�KW�&"C#Ű�y��[l4����Aަ$4a�J��y�m�h|�8�R얳vl�SD9�y�"U&:�t#�T4f��L��eL��yR�ǩ]`�P�,Q�`���L��y�s�V ��b�>.G�mxs�̄�yr�a�:J�P��8��OA�y2��x��ѳ�%�J����"���y��P�L�s��37=��{B�%�yr�)yLl���ڴ$5�X��^�y2�˖3"��z����D�I2��=�y��)~�Ƥjv��U�%h�۠�y��&�l����#~�Z��7	�6�y"iB�/�Duɳ#�sζ�1���6�y�����*�z�
��*�yBOH|Ģ�ˇ���c��W��SPC�	�S�~�c�"ƟP��Xx��]+E&C�3vw���oB(d�|��
`��B䉩[�%�&ݥA�(�����B䉔@q�y�4��Gs�U��V�o��B�.�!��%�6��eJ"C�%L��E�ԁ��(�IG~�CBů()!�DEBې��I�.9-2��!C�<:!�$�o`&��f�[�ABxI�B� J�!�$�����$H�O�[���A�!�$��N�F,ydH6`"������o�!��l��ѣbyN��X��	�A�!�+x�>�
֪�	|�z�ٔ�:�!�D����d�ٖ �ā�S��Ci!�D!┕����*%�"U��̕�?T!����8��䑞��zQ�U�p�!�$�.2�5���+K$>8��iǑ�!�$�$(�4�H".����@j_!O�!��5T���T��l� ��IT�-�!�I���	`w�6��ر&ĔE�!�d�m��a`��zT�)���o!�dڇG׊)`uB��TZu��*`�!��*F��L��Ė&5d�h��0;�!�)7��h��A H�@���l�!�$�A� -��|��D#L1!�N.X(�ʖ{ ��
0!�d�$3s�y�gJ�l���0��	5%!���p�P�;f. �<fp8k �B7�!�E�[yt�.G~�PQJv���!��:0L�wś?�t{��9E�!�M� �`�R�$�&8�M@W�f�!�D�?}�u��#M3�8ӥ@��C�!�u@<�T!H�K�zH�H�%s!�K5�`�!Cl��w%��ʖႛ8!�NG�4���N(K
ʜafB�%!�M�O��%�/p�p�A��N!�d���PU��{�q��`J�O�!�d�y�� �F��3��Q/N�M�!�ć�9x�`�a� TD�Y���!�� vX�@P��,q�DZ�z���U"O�e
,ܠ3�<�j��R�k�.��q"O���b��=��Ȣ���0|�UB�"O���Y~a9'�G?l���ô"Of�����Cf �eUh���"O��)@b��%�n��gI� K�\!�"O��I�KFT�=³@>��4��"O\�GI	 䰹.Lp��(��!�!�D�.i�8L�R����c��d�!�$�8YLԙ!��-* NV�3?��}��7aBwa�d��ܻE�n��(��!'�dx`���jq�CK�=,l�ȓG��"�CE�gn|sq�7n�D!��#�Qzm�!]�b�Iq�J�q�����q��\H2%���mY�cةY������lk�*дe���)m�H��ȓ'w�,ڒ#�'�� Ѣ�\?��?��b$��	W�Q��KY[m&1�ȓkVv15HO�N��R�-F�9C�1�����1bN�_�̩��� ��Y��j�HB���T~�0�S�7?�-��%
���@L�h����U�CD�ȓY���d �7j�YSg��d�z��1�n�	�jS���/4�]ؑH�H�<)��e�&��3@ �C��|�<y��O�&p�.\�(<Y�F�{�<�&D)��c .E�-Ɉ��$��t�<��a*}��X�	2����G�<�� E>��i�Q��0�� 3�XC�<�@!�0"r�d�gjӄG�8P���G�<9�����6H�AI�00H�V�Z�<��f�P8d�پG�yT��k�<�eE�q��y�Ԉ=/��Yy@�k�<a�c���kQƊ�S��DQgk�]�<2DZ={��0���1J6Ή�t�Q�<-=�(�dm��R�8�C�$I�hB�� G�$���CϭΠ�@EE�Q�C�I�3X�l���;�Bh� ��?e�
B�	�S�V�X�
��!��K�!��I��C�ɶN��2 "4T�m2J=y�C�	.(n�3d�=>��<ڐ��W6�C�	�]�hH��*N�V �=a��a�vC�	�Z���M�A��LP��R�6�C䉇79c��C�����,�2,�C�#	��`�c �;4F}b4nH��B�	�4�(IB���kX,}������B�2E�;�.ґo�>������B�Ik�!y�g\=�d�y� .��C�ɪ@�n��Ћ�Fd� ��'\ڎB�I����5��
z��@���F�8eZB�I� �|!�ϒJ@�e�F$�:m{�B�I�kP��"��]\����dg 0OV�C�I�F	�u��[3]t�ݳc�B�eC"C�IB���ф ?f�dP�B}��C�Ig��]r ˯2��R4d�/0C�C��	2L8PE.G7j��찢"�0?�^C�I�f�(0@#��\4`1aA�,7hC��	��I���*+HT|�!��%[!C�I�A���1�(�BЛ�G� 5�8B�	# �sGY�I�4P��_.DZC�(��0��Ն�.���ؔ3hB�ɇ+�MZA�N?���a�֕x��B�	�bP���#�%~�{ѡ�;y��B�/F�� �tc\#wQ$m��f�#@2�C�)� F|��᝜X�x���'�LyDT��"O�%�	?�bӅ��8?T�D"O6�!���LQ��EFN$&,����"O���e]�"���f��#88�` "Op�H�:j��*rf\�&�=�"O� z�l�
�X�4�@�p6ȹ�1"O�����ގv$&ш�Ie�K�"O�����\�20�5r�_y���R�"O�%�#+ |ˠF]h�4"O�bf�T	~	��b�BwB��"O
�� �5�HݙE�n���[�"O6$� ���}�(� ��r�P�"O:cO���)�Z��,xe"O�pQ�HF��L"aȓ?ϖ<�r"O����'qP<��l��[$�p�b"OZ�yS�$��apH�[!¨�t"O����JC s,T���h��)B"OR\��@܋FN�b(�����"O�E�pkļbBh��>͠Q"O�H���cƀ\aBg��O|���!"Ob��3�P���rЭm<A��"On%��ɡf�-�AÉIk�UBV"O8��2�F�8�K���p��A-D��J�嚒O
�J%�B!n�h�	-D��PA����ұ"��<�d�,D��(1�E���<K@�PVpԃ�f5D� �1#�_��<b�L|m���4D�d���ٖYH	p����tpZ �/D�Pk��ņk�L{始�9�PR��*D�8�4L�=݌�〣��=n{�('D�p�GAM(u��A2dF�T�P���%D� #��)|�xHeC&��tp��$D���G5Xs��c�T�	��Ƞ%A-D�hء�Ny8P)�f�"��:�*,D���(U�L�mP�Ǚ0�t��*D���q�A���9�,��8��J"(D���Ս^�F��u�W�Q�´ �+D�$3UG� ��A��,/ن���(D�d��'` �	�eҜhĜb�%1D�@B�?����Q#H��"�*D�õ����9ℐX0�E�#J3D�pF���W9̀���~]L9W�2D��p�Ɛ� \Z\�P�ȮJM�u�6D���$�>8R�&��N�^��'�(D��Ҷ�?-� ����:�i�,9D�p��Z�/D��d�W<s�,Jo9D�<�E�4r֒�����3��D6�2D�܋Q�@�m��e��4Y�1D���ǌ48�� ��0uG~0��4D�\xWn���`�*Ƃ�jؘ0/2D������)AY��h��P�r$R��b�.D�܊�V1N��L �I� 	7Tu�r�'D�4�'�˯+��0�	�	���('D�,�A95���Q$J Z	2�+&D���P& �d`,<�Co�=��tB7�%D���g$B�ky.��$��9n����."D��KƮ�s�4�D\(>b�]���5D�`3��O#%�lq�4�s{Lhz&i2D��Z��ż$,a��˔�CT�У��=D�HB�/��Y/0@� 
=��T+4I:D� Xb-�N�pE2�iS���I�C&D�����۝UR(WD��(z\L��%D���&ht��wN�g84���l0D�T����t\�m`�Ӂc����/D�� ͋�'\�9R�����<:V"O|M���$^� ��3lrc�	0J2D��[QlǮ=�����d�:zȰr�-$D��pA�����2*��Z^�Ը!j"D�\`Ǭ/69��!5�]�0]@�c 3D�@#B���b%��mۃ�.𺰉2D����+ؿ[�<���aV�	.�={D�=D���'�Kyа�����CW�i�a;D�T)$�@�@"%H8%�9��;D��`@�6@c�ѡ�AO����32�4T�Ps�EQ9i�4��3( Z�"O!���	v�||�u�Q�cͬd؁"O� i��1f��K��v�0!r�"O��;�K�H�|P�$Q�v���*�"O�m����$kf�&,x��`��"O =�ƥ�?��8�̅�s����s"Oh=K ���bg%��\Ѱ�"O0��F��
�%3��U��9a"O����-逍!4$�"|0D"OP)#�"�/��`ӂB�f��+2D�Hk�>;3��am�h$K
 d)!򄝑����@�ΌN{�Q� �u!�$I��;wh�&dE*@��fZ2x�!�d���HaF,�W,$�ʰe�2v�!�$��V�@����ݬa��1A4ɎB�!�dHj'�+E��0�B���d� 4]!�^�:%T�p�W�5o��!�M�/C!�D�Jt( a1'�\m� (�/O6!�=!�����w�pu�F�'L!��:>g�m8+�/9��Qk�ٰR�!�$ǉ!H\�h�l%:Hв%�>7R!�ھy�T�+�oP�^�H�5�D5#W!���i];��@$e��u�P�T�.I!���"a8$��s�?��](E�ԥP�!�D�IpX$�a��m��H�!�.l&����IȻq�LB҇E�!�d��S�Lic1i�8j�T��'�&�!�d� �N��C|��9�b _��PyH)2����Cnӱ��ԡb�[�y�eK�*�v����J)h�e��+�y��M�G�ll	o�+u����6�yr,JvP�LQ'T��\ ���yR�1c�$�`���\y������yrCG3S�lԚe(�(9d����Z"�y��PB���/��A" ��yR�/�$��tg)���Q��N>�y��?�(�3!W�	����@�J;�yr.�q+j4�&��Qʴ�f. �ybIS� f�B�M �A�(�9�y�S�4��0B���[<,���3�y�
΄C|����ҘK�F݈�o�$�y�Gߝ=�Љ�Y�D�� �Ə��y���S#�y�L�CmT8b�E��yR��s�Ɣh�r�������y��R�	��my��Z,{nZ�F�y"D +@�.�����w����K �y�̋�AYЉ@jLDE��y�-Ήq9��嘘�$�t�I��y�AӏUҶϐ�`��s�K��y�L,-�Ѕ��K݅]�b;����yҫ��>m��#��MAnx��S2�yBNMt"���b��x�,�H�D�yr� 1��bC.q���"M�<�y�D�</�11�O74�,�Bm�=�y
� �P��*H?�e#�㗓s��E2�"O���u�>)��M�)�6��H�"O)%���$�V����		du���U"O�Y@c�<t��T8��OOx�1"O�e�f�^�Um�0�cA:'�k "O5����]��W�&5�D
"O<=��!!Ϡ��"�2*2,�r"O���IO�2 Ƒ���Ͳn�й�"O��R���7�Qhp�V-S�<���"O��)�ņ�E}Bq��>X#��;t"O.Ma���u�X�m�?�D�Rr"Ox�J\���%a�E6���a"O���&�[w	^T���\x���"Oz�&I.TQ�h��x��p"Ox���I�[_ZQ3 n�}��S�"O�3�ܹ?�L��#�)Z�ܱ��"O�!��\4F8R�V�ڇ/�-�D"O���R�8O�N�̄���5+�"O��RL��3Ҁ��섚�"O�-��F"4yZ}�-J�!|��"O� .�0�9P�Ǚt�3G$�0�!��Q�8�{��5���&"&qk!��8H��Mw��E,�}C7n
3q!�dS j\� �T�¬;~h�-A�!�T��mZ�c����2��%US!�j�!R�C��7�T���M%!�$ԃOO�� B��I�న�H��=�!�H�a��%���T��݈�&[!`�!�d�^��Dn�<РY�e�Q �!����0h��p��1����儜�!��G?@�A瀉�ja�A�ѷ�!�L�Fk��ha� =��|��	�:�!򤃐#��Ӑ�R='GB��G r�!�"`�V�Y!�V7C��) ��ӾW8!�d��H?4�@7�\�i�. VH!�dGY���k��5��LIzD!�H3*9"�!�,�+�LZ�GJ!�D�.~%� ��M���N`��ˑ"	+!��ЀY*b�)5��<Oa�	+�H\�/ !�$���L�R�+Y(�uxw�܂�!���'���Iņ�J�5q aЩ�!�dY*\�dp�s'�(rx��ꑆ��q!�$�*,?phsp�
 #f���Ce��mi!�$P�Y3�A%2K(h�BF�`W!�D�(�J��%�:6,��!ŤJj!�DYV���cS�߮}nU�bo�?�!�DZ=(J����'kڑ��nC�^�!򤕚@
�đ��"��ա�M�b�!�D]�	��P�G�ߪ���] �!��'*M����R�k�p:�,��71!�d�K*҅�U�S�疭���MB!��2��d8P��*�Y��S� !��UÜ��&�V�d���rJ��z�!�d�!������{��=�V��!��v�^�#P�H99�GʖX�!���rX�@��?0�A��^�g�!�������ВPN� U�5�!�d�<	�mB�AU5�1��!���w@�ĳ6(RK�A#�B�.8�!򤌩kw�h:E��-�&XYs#W�:!�ޛg��" ���薽r7!�d�����qϓSڀ��5���2.!�DO)e��� �^l��l�,�#j&!��S*]� � �A�>O�L�Q.��h!�� qѵ��1�d`�kW���"OB��	�72�� P��1M2tX"O��A����2� ��9Y܁�"O���E�S��\��L��9�4��"O���`^-sz%���&+q����"Oh��`��-bx}I���tt�'"O��ɶ�̩#�t�j6MD7��Q	"OX���$ �f)�Y>s����"O���<t�0̊�� ]�rua�"O�-BS@Z�%:|`��'|��B"O�`3*�!��i�RI�b� �"OPL13��#�Hq{h�4FQ ��&"OD�!�.�{r\ s�g_1��D�c"O� �J�+��n��?ɜMz�"O��(w�_ca�D͋*�� y'"O��a��ǭ^���Gc�#G�!����:ɠ$X#
�r @��ʥ|�!�*
M:g�͙<�����̣b�!�$�)5] hrt��<O
8���7�!�ˈh���A�ܕ<P��a0�H�!��xf��j�6G* �f+@�%N!�Dx��p���;<�=�p�-?k!���p�peP�%~�i���3�!�$�H!���ANR$r�"S��\�!�dUQ �l%dǉ1v0��3O�l�!���M��	�n�>T(P���|�!�$E�FLղрY�87�L��bٰ0�!�O�$ܰS�1/�@�A�q�!��W�N͸EӳaL+�2�j�Aێ'�!�َ�d)Y"�ܡ'�d�#W�P�]�!�ǬF�l9�)r�"���!�d�7H�@i�#�[�r��)g�!�d3M��Y ,W+�����Y0@�!�$
�ȭ	wi	[�0�zQ�^�Q!�Y�0�25�#		�0uZ�:GK!�بX���[p��`i�L��,�K�!�DV2%��۠ƚ�DB�����ʪ-�!򤆀x�.M�ŌI����hwkL�s�!��×&��}A4���W���0��1�!���be^%�% LByTX��IL)!��K,l�H�A��|l؂�iB.!�$��Y��X��.Q�"y�T�FV�R�!��ED]�i!���~V|t�昒K�!��
��pӡ�j#THc���q�!�䚺w�p��1�;'#��i��No!����EZ�o���]�e -�!�$3!��2�#OHz�C�0,�!�d �lPR� MP�r�&�����!��هv����7u��1(��K0lw!��H�h� Ie	��E�~)Z�A.K�!�ȓC.�@в�ĒU�N��V�Bvs!���'W������1k��� �6q`!�M�L�w�\�n̎P��,R!���^�(  ������,)AŇȓ��y+«�#T:l�r��*
D��DW�ݨu ]GFD��L\�?0������{6(ȫ\�$)k4��7��}�ȓ�!K�!� ,<�"$m̘h?�y�ȓQT����L#�e� ��T��ȓ~��a��S?p&��R�@4�t���9UTUfZ5M �1R�C.T ̈́�#�t��C���ij����]�Ԁu��:H	������Y�@��t� H�ȓ/Q�!C�D�~ ���M�7"��(��S�? N<�$��mU�Y�"�ɠ���"Ov=�DKH���Bs�ƍ����"O>�q-\�:��yrc)H�d �"O��[n7+����%Ȩ1�&9�0"OT�!f���8�*�;��ӓ"O@�����v��u�ѰKb,�B�"O�U���ͱ>3�XP釕3_�2e"O��!�Nl�~ #�gkBh��"O�A�7	C���̨1�N&��"Oy3"EI@�1�O��� !�"O��cNNg�����N]�p����"O�#��鸀
�N3f�S"O6���"Qt�k� �5�t���"OL!u�ܲ4T�\�c�<���� "O�����U�D��cB�L���"O���b��/� �?=^ �"OV=QC"�rkm�C	'=j$	�"O�Q���Ld�@���S�+I��"Od��A�ap9s1l��z���pG"O����"ŪD��	`��ؔP�jI��"O�`9�#N;Qzd8�0最s��՘�"O�@*䌛^ `ٲ��I=>U�c%"O�@�O%d��	J|R�|X�"O�U�ѩɁb�n-Z��'dg�92Q"O�Pĉ�8^,���0"Yx�F"O�� �=}.��$ؿ]��"O��k2 ��,���3]�U�a"O�)�B��/ʌ{��i�q"O@9 6��#ɂ<�d�"q(��"O�t`��K(!�H=s��/D\a"OF�UƟ�1�@I������"OZ	��:�>�2�3Y��h"O�m% la�ٰ�/B}t��v"O�܊���D�`�!�%Z�-y�"O$�S��5�V!	��� 8�H�"O,TbA�%G�4ȁb�$�r���"O�( �̣9ҊT�p���Q��(��"O�1�Y�V�PA�ɍ�@?�"Oh�ӂ%�x����'Η�+�ђ"O�a���A,��A
N�.2n�H"O�0J��OuHQ���ɭ;6j�""O���a�],=J�1ԋL"~�Qɤ"O��D.M�}^�e8��/Rq"O�XA׈Viʴ2dH&)��`t"O��v	�*���)@A��]\А�D"O��bf�<�Hj@"�,P
�q�"O:�[�H�$�����)���t"O� �#K?nQ ���Q<s29%"O�h 4$��jt�Uj��p9����"O��@�ÓCPR�Rs���,% m"OnA�BO� 8�|b$�����6"O�y�2��1D�ȸ 0�.z��b"O\�'�M
����.%f��d��"O�xyq��4���\�x���A�"O.I�LHr�8"a-�}Ҭ��G"OP%�%S�P>d,��ō9N�j<��"O�Q�f��H|�����O3��"O^} 3�ƕܘ�j���d.� �A"O��CP���G��=�!*�,o d !7"O�|�Վ��$Fz��(ĳu�&��d"O���W�b� ����'s��v"O��M��[�<ؘ��ްc�\�"OD��#J�R���3E+��0W��Zu"O!�$ִF���P�S�.8d��&"O� h  B�ѭel���\"T}��"O�åY%|��3\�ԸP�"O-qv��_4N���ȱ_���0C"O(\*F'ѥS	�X���ۧO	z���"O��z�ŕ���1��E�v�p"O ��K��C_� �́1��Q*F"O&�����#p.�\����.���"ON��3�]�D͚��@�f�4Xs"O�8�&j�%|��ѦA-CMf�� "Oj�5ȶ�RIK�͒s/���"O�4(���
x:~�*ê�H>��"O���ӥQ�\f���ގ!�D1[�'�:i��E�}|yۣπ�F%@<{�'����)J�	�R�0���>y�=��'dA�e��L�����40�I��'U�3�kL�K�z,�s�P�/�x�
�'&}��F [ՎHZSi�&�f�`
�'�j�Z������"dQ��*a
�':D�I�^K� "�l�2��-�	�'�\*�e�	��q�5g�)Z��S	�'ڐh��!�{H 5��$w'C"O�q鰦ٍr�����<]�D���"O|�˖.�V�5����Vr([F"O4�wG�v�2s/�	Bi�d "O�=1��я�0 ���@7Q��r"O�(��0&���3�O'i9�tCd"Oh���E��������,J�d"O�
��M6L���)����"O0 ��E�B=2艃-��~T`-�"Oڬ�@C�
~q�P���.8C,\ç"Ox���F�/!�$�$ն���F"O���S��p9�J
7���"O�d����e��"�_�it,}	r"O�q8cmG?is 5��@�\��Ғ"On=��Ê�v	���X�8Q�W"O���F���B@l�SԂ��j����"O��X�B�=r����kDЁ�A"O�q���_��M�\-;�-�"OB�gD֜)�2�͐�|��+5"O���p/�<0ä���5C(d��"O�}����?5X`�&�Y��DD
�"Oΰ+2e�V^��#m[ =�N	��"O�,�@��H�r��V�%�Zĉw"O2ܲ� �*q��k�a9}9Q�"OL�
CC�q �� !�=rh\��c"O��r��
L�g ٕ'a��`"O�d0#��7�Bh�@SX�M�"O����;0p�C�U*�4�U"O�u�.�2cq�(���-E�"O2d�Շ2, ���*�~=x�1"O̠�$�Q�m�(Ci�"y:P�5"O�8�&;2���.�\����"Ox(�
C Tۄ�۶͍L�DT�1"ON4����>
��S��M��:�"OX�����8J�W�+<(��"O���a�]����*�>}8r�""O��q�Ͳ1�0��ꂛj.Y� "O4<��)V�s`\Еi�;M��{&"O@���	V�8�r���J3PRmi�"O ]A&L����1�Ȕ�?,�I�"O��B�1<(�0U�Bg>q�"O�4�#�7�f)Jda�*ΜB"O�����
~%Ơ�$��W9~�T"O����u$T!R)Ko/�(�"O� �Ӑ��,�R@���B*:���"O�<�6�=��xZlMh>�	C"O�2�l� Q30+ �P0V���"OF��P�a��@% �!�pyPF"O��8���|�8V��'�210�"OZ���Єb�
��P'� w��5��"O8#q��1�����
}O:
T"O��"�!�I+ �V�C9
�"�"O�]@/�&x�Z���	;"�ly%"OV��@`҂�֬��+�l}A�"O��*!㎴N,��c%A����+#"O�Y��5_��P*�����"OI��ɞ�s �  ��yfA��"O�<(��Uaڨpt��9 ����"O��v$�
I|�0��e��I\z��"O�BO L4�1��Q�$&$
t"O�qF%F;^XL��C�&�@�c"O�m*�F��U�()��V=:��ԺD"O��$�#�E�w�
�A���B"O ��H�\@���ˌj�F��"Oi��C�����oBV{䰀�"O�uR�U,cZL��&��_k��b"O:�����fsH�*b�P?D��a�1"OL;&ж>�>a�G��3U��"O��R�)  }ba�gjV*pAR�p"O��r�*�G�d�{5�P�>�:U�"O�:#��g9<��E��3�� JF"O.ݣ��Bň<#NT��l�(E"Ob�
rĔ�R��U�+��2����f"O0��0��$��2�X�8�k"O:I� EːSs�%�Gފ|56���"ON���E	Y������2|���Zc"OĨ �H��Ee��iSg�c��x�t"O)P�\�#@ ����8)��uk2"O�hǭJ�&�
4�"��	���@�"O��� kγh�-�KG9)fN���"O�l�T`�ΰ��4IE)��x
"Ol<��mB
I���z�	�2�����"O\�Y0nQ2V�Qa�B�w�� "O�a�UI�2s�:�#U)֑mn�Y)�"O�ر�k�Z�"���		Q��X��"O,y�̟��D�
�A��|�Д@4"O6 
�����Э^)`��Z�"O,�1�	��f�l�XaM��Q,��÷"O4���	ӭ _��W��/2/.��"O$ �"OH�Q�q:��=�>�A"O�d�6�F,�p`�BIڗe$�l �"O޼˷*�c��iR�ʆdk;�"O6U;V���:%k0n^�IP�{Q"O�t1q%?1�
0�� R2�Y�"O�̢�J{�X5%E�P'�Q�q"O��G�06��#&�`�1 �"O,�Ƀh@�
�;2k�k�fI�4"O�)�w�ۺN%���i����H�`�!�ηHm�]����,��B!�13v!��ƣh�F=AMV.T�h����&d!�Ą*���0 �Τvʬ�¯V��!���<딴Y�O���ٓ2��/Z�!��� Z8�U"�
%e�h�-�B�!��ԘA5f$bp�^[a��x�Q�-{!�D[S�����׷n[L}�AYj|!�Re�j�jqHI*P�r�ן!��K��	�QB՛T�\H它�+�!���=q�@�0��p�.�sT(A�~!�� ��Ɠc�@�+��[?`(�i7"OX@��	;2C@�a�-Q�n�� �"O��&Ɠ�-�����쇃G���k�"O�\؂�+^��c0̞� �A0P"OF��rfK	W��Xp
!�$Dz�"O���d��l����^��n8h�"OP�ц�B� �l0�$�Pr�lYS"OV02˟=u��PP�ɑ�"O�,�#�q�����G�p��"O���4�^-+$D��@/0�ˇ"O:0�eg� I��ܪ7	��e>� "Ob���$�2Q��ԑ�g����W"O�M#TO��py"-�օ�� �s"O������đA� �FD�4"O<q�!��H�����]��U�"O��kC�^4$4h�!B���
�y�"OV��v-¶0e(��P����a2"O��� �CͨY��)^�>�x��p"Od��Ӣ���B ��1,��y�F"Od|�G�ɓ4pHS&�\4{��S�"O�p�r��V�`D�O��ț3"O"@3U`��
	Aam��{^h�"O�pbA�ɝ|���Sı3nHʤ"OV����l�:%�BA9]5���"OT��N�>�z�)�
��p9��SS"O�t�f�m�����T�^9�"OF}92R�IՊ�bgI�;�����'�|�b�ņr��� ��T�@��}+�'��(���Z�z����/��>� x�
�'��{0Ň�q��4��,ض2,Л�'�݃U��*eU~iH"�ć�^X�
�'}DZ%�� [j|�����
0�	�'��(ׅE�'�.ݳT@^�6��<��'��$��� h�]�c�\�Y���'�&mP䆒WC|�B�C�y�

�'��d�	F��-�0<(��a�'�Pu����{�`�[A���7<R�
�'�4xu���,�@Ca�D�.��i�'���[���o0h�s�� f���'.��f�!�0K� �:g�Љ��'��I�Aڥ}Z�Y7�8Qc�AA�'�*�`�/�!�~U���ϢO�<��'ʢ��M��[a�Dp�Z ��p�'{ؔ��0j9����� gj���'a�2�[^��cQ�~��j�'۠=k�.�����X�"n�`H��'�̉�S��;e+
|���x� ���'A ��ul�=�,\���ӡtf0�i�'��I���2t{f��E፞x��)�'?֩c�ѰO�a
�8bL��'(���o	v�4�%����u��'L��'�׏-�LMB�3-߃cO�C��9: �X��S�T3:����\A�$C�	�AHճ��:�(=I4�D�W�JC�	/0���'/�.B�He���:Y�`B�	��
)b���+12	c�M�!7�~C�	+�<m���ޔp,��&�V�LZC�I#^�e�c�W�.	� ��n� C��?#g�0�v,�6ˆ]�'b�a��B�I�{u���W� �^��� BD\B��;*�n�x���e{|�;7�[�y�Y0@��)���`
r`���y�N�>
vQp�	1 
i@���<�yB!+��	C�	z�XY!�\��y
� 4X�`m�*76(y�6N�&8����"O�ɪ-j�� �1�%��Y�"O^�ia �!ri-C9O	`"�"O�,���g.{Pʏ�M�n��E"O�YC��΁fnE���9�Ȃ�"O��{ǂ.z�p�!�\%:�.�
"O!�C��<_�{���y����!"O.��	�+x��!�jؙ9&H�g"O�����D�H�h'�����H�"O�q+���J��q�G�	�z�:�"ORM�������A�e��ͼ#"OVuk��H�~$�	3��.���k$"O@a�D�3&�f�e�	 �
�Z "O������M�$�+&,ٲ���q"OQu�$n��I;g�� %F�-��"O�d��G�栵�
��,��;e"O��[�g�Ir]r2i�0m�jQQ"O����:�rL�5g�;dgf3�"O���
H5S�X�B�oÎr��Y�"O��K���qaIKo
H���K�"O*8�B-84Z<�F�	��x2"O ��b�3i�LuX�	?���2W"O�HQ2o޿L� �s&R��ɐ"O�u�d�P,[ZRh�G�׃%A���"O�͡q�R�"za�b�7�+�"Oh���)<bdl�P�lM'Ȱ��"OR�k��NY�����[B"O�0Xf���?R|x����`p�uP"O
EhW�1>��3�ϿnuL*�"O�,���T7 �iڇoԻ�,��"OZ	ia.�%d��X���M�
�3�"O�<�T��e!���D�ܳw=�݈V"O�������C�h�U/nPs"O�d��cD/l�EbPȔ�I/x���"OIj�$H�+S�A��g�	;Z}"q"O���.@0s���%6�D��"O�( �� ���K�sJn��@"O��8B�,`�8P��ϳ.?�q�D"O��Q��#z=ڂ�ϸl]$(Y"O2�bu�
��|E����TCD5W"O��>=����b�6?<k�"O4\��!]Ă9���?#6�`�#"O��j�%*�����U�+��i�"Oԡ@ǯR�P���À���w@�0P"OJ��֤�7 � �e�\�)��l��"O��3%�� А��#���:f"OZ��损uTL��V�\CV$�q�"O��0���8����N>i@tt�"OF��N��z^���N�0;hġ�"Op�:"ML k�@��&_s3��H�"O�x��#P:)���#���1�8�r"OȰH@Gd��3u�D�Lvr*�"O�
J��T8�	9��h"s�ʂ�yg�1�!��F�b9~�SlP7�y���)e��@d�Y�ر�E��y2O�D>$`#Ve]R�4���B]�y�SA���[3v��,�fѯ�y2
2 |��r��k5�E�͚�y���:�RԚ���]�N�!C�yB��1�yX&� BW2�#�U�yH�
Th	R�H� dQ"�+p����yf20:��W#��j�R��G-^$�y
ޟ$����%�G-h⒰��T��y��B�N��뱨3WS&@@�e� �y
� �l*AiɈD!�9�F�T�Ya�� �"OF c�Cʛ6e�Y���R�2:��Pe"OL1��[eʽ���+kώ #"O0Di�(�g�$�WIm�P:�"O����ޅV4���$�2vi���v"Ol	�#wR���(A�Q^lcr"Oм8�J��[#�:b�هbF��@�"O `:��U\c�����$����"O(���2z��)K��K���|q�"O҈ѷCȦ.Ҁ5�EN�l�`Q"Od-�d�� H�T`3��ܑqx����"O��P��>/���J ��c���#"O��3�ܰt��d�'��s�.T�`"O���C�\9v�������yZ��	e"OTj�
Q�4 ����In�B�"O0@���]�}�y�t��8M��3q"O�Ԙ�����d�@OK�i%<1��"OHa�!�V�D�\`�ۧli�j�"O*���@ !H����T"u�h��"O�+5a��_ڨ�roS��QxD"O(hp���D�z[�(]��N�9D"O�\9p�W<2����6HY�^uR�"O�́tɚ�Xغ��HK\mK�"O�(:f��L�u��C�>WJ2�R�"O܈�T��0���@%P�S:\���"ON���C:���w-�3�z4��"O��X�H\+9��Ŏ�
���"O.�P��2����7M�$d�2�cR"O��Q���z  ��d��d�*�c"Of����T��D��l˧U�}�$"O��3!��4�"�ӳ�A7k�1��"O\0�Ó,��p" �ȸQ]���B"Ox�c�
G!���sď�eT�E
�"O����6~Z&�&v*���"O���BB�k��t
�B&)�e{�"Ov1I�
�2�v5��::|��"O�y���� H�t�R�ƓWFH��"OP-ct�)_] �;�@D�1&h�"ODM� -�kS����ό>O	��ӂ"OZ�b���=��`��B	x�S"O$�h5�^GW�`��ժN��z�'���ß&#�칑���o���
�'�Tl��,��9���t&�b�,��
�'>����g[�"lH��U�W�^�-x
�'c�%i��M	N2Z��q���_О]"
�'�$��*��G���hk�#U�ȴ�
�'��\��`Ҩq��i!�o��Sf 1`
�'wF���Q�!fU��%ƚD���	�'+
��!I��nm��jD�R��u��'qĵ��n*�B0��N�Z�8�
�'���+B�[�T(�X���T���
�'�p�`4�v����P8D��U��{�n �7�A&x=���dȄ1g�:u�ȓ�D��iͧ!Cxt��HL.k���ȓt$8x�R�������	�C��ȓr��0�3>I����Ŕ'\�*@��:Z%R��H+p�cťO"qa� ��eVM���Q��L8H4*[���ȓN��4ق�;,Xm���Cy\Ņ�-�@ �&�ܓB������crl��Wt\}8t���ab�h@�^�jR���ȓ[��)	@�E4b&,�6�h,�ȓ-���Xr�H��d�س&�V"L��ȓB�2}���,@�L�b0�G"^i��S�? ���j�c��{3jO(gv΁ia"O8h����HwD��T(D>S�8!�"O.ȨV��H��U�B�ǒyxZ	�"O<Y�mJ!,&�
Fr��kB"O�M�7ЙI�5{r/ϧ|F(ȱ"O��pN[� 1���Ύ�Lh戡�"O�i )�:�̹:sD־Te2���"OlT�C��%C ��ׂ�H��@h�"O��EA�T�XRaGB�	h�S�"OE�؜ʮ�񦝷<��"O�*&7-4-룥cH2$"OT	9�E�+nFdЁ�{x�� �"O��#�30j����I�0��c"On� �e��*8<}���L�Ք��"O����瑦3 �$��,|���)�"O����Ce:�S3�8)�"P!�"O�i�f��4u�t#����W"Ov(�t ��s����k�y�Z 26"On�fm�"B�,3%H���Є�s"Ox)��^�"�]s�ǲK��	�"Op�Z��T�݀%z���+� �� "O"�3Rj ����XiU��Hẗr�<��G'��I�fE��.>q� ��G�<�UƇ�o����u)B+p �\����l�<aC�B�G���$�����f�<ѡ���H�{���m/tqra�{�<apNIZ���8�i�
qVLR$��M�<�7��Y����d,+�z��s�L�<i0h�}���Ӿ�L,�nYM�<�b��/��`���W����^�<��KW�Bn��.�K��Pc���<����pH���^���RJ�`�<9)	p��ȠV����I�3"_�<&.� F�bd O�=������@�<YP�J+/M����Y�	baI�y�<���Ƥ�����0G�ř$�u�<ч�@/��)�P��4�	��n�<���N&�xbP�̀ozM�ī�g�<�S"����h���IA)n��g�<q���	|����ȋ"��@po�c�<1�kc:La���O�:h@�M�z�<iWfH'j���*�&� 	��ɱ�s�<1��.M�e) ��;8�$���T�<9 V0`mR���^�G:�i3 BOF�<�$`D���!4|<��S��V�<i� 4��W,�,V��Uãi�<a�ٝRs5�6nL(H8>m
���j�<�CC��09!鑦+;����+n�<y��W�a�u�Q#Z	���s�^o�<���C���+N��Ai$�i�<�uh�,x�l[�K�Dj�LɁA�Y�<Y��:`�D���b�t�J�YsBS�<aw��=ZVJ�����L�s���T�<��8⁈p'̳^x��#'�_Y�<IW�ߖk��m��AO�q� ��JM�<	B�=>%��31E(/�8<�ny�<� �W$S�f�Gc֎UХI��Vr�<�1��6��CNҿ6F�P�Ѣh�<��ES�,x����ּ�ht��DK�<���v<�IKչX.t�`� J�<�am�Q��Ib3�(؄q�+\B�<y1�V�D	*s(և��!Ș~�<�`KQ&g�,H�fM�3�HF��B�<�R蛍^�H%�E�7��q�j@�<� ���T��(�XQ��H�t�b4"O�eyV*�=Y8dkgn�s|����"OH顡�'�!dn�tPظ7"O�aQ)\�6�i��._7.�L���x�O��4�ʺ6xɋc�B�H��'�`�cf�p4������k��R�'sF�S �E�T[���L˪5�b��ʓa�b��׮C!L~�EX�����ȓC��V�2�*�+����){�Ԇ�I}̓^���!,��<�׳�!	���O(B�I	s�@h ��9ox�sVMM7�`B䉘م� LYjIZd�@E	�:҅7D�B򩅂X�&!ۢbZin�Ѫ',)D�����U'Z�g�%7"D��7%D��'�� >�*�-^�i~��' D�ر��I�wq�g'^�/��$�ŭ=D�"�%(#��|�%
9� 2e D�T���	\�m��g�)�&�+$*O�\��øC��A����`����"O�x;W��
A��6����s"Oh8B��9��H���Gxܥ��"OlA��Ɋ |+� ��m� �њ|��'��p
�V߲\�S�
`�Zt��'aR��C	��P��x�K�P��(J
�'AZ��Q�LI��X�b��Fu�!k	�'�<�C�S!!0��UoB6-����'Of�dG�KN$1��
!��@��'�6���ݞv�~�U[	�����'��GG�Bt ���Ѥ9��Eaď����#�S�OE��K��
�@�A��֟ 2 ��'�0-`�o]���Y �7P`|�
�'ۢ � e�MY�-�&Q�)+���'���! N:4��$q�LxB\��'��Hq�غx~p�Aa&O7���
�'�`iS�8��������r��U:��I`6�֚5c>�{�$_���E��N5�剎|�Q��|:R��5R,���&�qaܡ�`a�a؞�=�n�#Ye�� ��Xii0���L�R�<��N�S�˷��[88<Q��LM�������IP�?`i�hc�K���ؘ��cBdB�	�-�a�+R�بA�φ?9�$�<Q��T>}�׎ N��$��4]j`��%?D���^�{��]X��˵;EV��Cl'D���Q���Z�b�ؑ$��4Bb��e#'D��D��01�'
�Q49@�'D�����8�RdЧV�,�2Yc0K*D�p�vy����X��e"D�,�@�2���eJ Y��lh��?D����Zh�f��D�H�[B���'E<D�� Ư΅Qk��bD�.bD 7�4D�X�VF�8s��L��:aǀ�� 1D�tp0̆#:f�]@�*����/D�����	��0�X��X��2ɰ�l"D����]�9Zl̻�Ń�f�,q[��4D�b b�7H&lP��&>Ma�����=D�t�q�A� ��pRf���}gѫ�j8D�ts�[W-L�Z6I�>���4D����bQr(�Ť���᱈1D����Z6C-�}kpB^�a�ʬ�*O� �I�+R'��1R:�g"O�PB7�ߏ5.��-��>:NmRu"O���
T+.��`f���jp���"O��p�<-�j!B�IW�Xp�q"O�BS���$:bIX�(\{ "O� nPBN =u�$@��A�Y�# "O�C��wY�e�@M߮��"O���HȢ���¥L��Ii�lئ"O��2m�"��|`�n;+SX�"O\lIի�2(�x�˂6`�V ��"O���9w�Nܫ+X�JOܱj�"OZh뒦���D`Z&@J�M9�X�"O>�`��>� ��Q�-i(�,{"O��8R�I5�"8� ӥH�)�"O����jÛ��s)�	kZt{e"OVpz�ݝlk&� Q)�v�J�K�"O����+��
���S��3;֝�3"O�P�2�ִ)S�Ԃ0a-.3����"Odu���<[�ԥ)�Ƈ�2)�4�v"O��)����"o�<#�ƕ !:I�"O���� 	@� ���`����"OQX�lL�E��󅟓K�2�j�"O�d�5�<�9�. �����"O��An�_�d��G�T�#����"O<D�L�W(��D� ��S�"O<��ήv䙳��ɑ!"�s"O����
�R5T�y�ԪA�L�"O��[�&-`ph���J�7V��#"OhxR�!�s.2�ړ���^�H"�"O$�82+�V��|�&�8{m[�"O�x�KL	i%TJ�#�@��"O�U���	-V��z��,~�ʐ�f"Op�:D��0�z5S�c�b�
�*7"O�����Z��d�A�;�����"O��B0Ɖ7{��8E�q�
}�!"O
̙��0 �ԸӮƙ���X�"O�L+@C�,Άܻ�l�>�t�"O��qB�<+�"yʄ��b���"O��Nĳg־e��!��� "O�e2�J�Dӈ�зJ,6�J×"O~��d�6k����Ò�8�r�Y�"OtMؕFl�V�V#�+�*E��"O~E� 
�'E\��	B����9�"OT�q�x_��xE��؁ҥ"O(���(�?2�2u�7��.�.r�"O�Cw�T�5kXZ���'�n�[�"O�q���"{��qW�2�"<ѡ"O$����=-���!�ļ�4��#"O����ט� ��I��Q��"O̩�T�OјU�"ID4/��X#"O����[\Z��7a	�Z�!$"O��H�"[ sZ�A���x�3sBć�V���৯�eDh�*�A�(X@�ȓ*>��0� ̉u��\
#Zr�؇ȓw����ћ@�h���`�*X^bP�ȓi��t`�*���� �q͚K~$�� ������+B	�EKbAT �y�ȓA�f�����  �p��&��ńȓ��)SЧ�7�����%\��f�����/�\��9!R�W�\��8����#D[C� Txcl��UI�ȓ$4�,�Vo�.D���d�=X��ȓ(�@K�ƕEs��c�J]<23�t�ʓ5Q05�%n�:�|�"�\�pB�	)P6aHu圮z�bu�tL�2�xB�ɕ}��t�aJD�?�<	UڋS�C�ɏu�P+��.��R��g8DC䉵^]"�Z� �	hV��ҖoכE�C�I���)HQ�
>6��	�A�O,�C�)� :i��kL8)d-�./z��u"OB(�ŇAd�,�u�^�9��q�"O���#	h�u�q���p�ֽ�"O���*
�Ly!�^ y�A�b"O��[�)D�{z� H�ǚL����#"O2ȰJǽ�a�g��9c�01Sf"O`�r5��/)��Q�"�JhI""OR���)Lo��Б.f�"�W"Oh�X�o��$���(o�_�L��"O�D���	G�dX�VoK�O��l��"O�tI�r��0e��[Ӡ}�%"O:�
�n�3;���6m��v+ �0"Om��-ܘ�d�ڄk�!&;���q"O0]9�D��$P����t*@�q"O>�R��_-]����t�e�^�1Q"OT`B �ƛS�Љ�i��^ḕ"O��խ��!����� _�`Ȫ�"OBu'�	o�n�j4�)�\aA!"O �'b�~�80�f�'zn�r#"OjQ�Rѐ�J�B Ȕ m�!7"O�Y��d+s���� �BT��#"O�&�Rr�$ԋ��F9"K(�S�"O"TQ#  R��}QVN܀G���"Od��v�ۇu�|�
�b/.~��A"OT8�`C�\N��!�_BQ� "O�H�	9�i�V���o��Z�	���iZ�ƺ*�`���UD|�ɢmw89�F�Ex��!��Xff�C�<p���Ӑ#'�Eb�+"3 �C�IHR�<2�>v�	���BڠC�IPD<���ą�oy(����γB
�C�	/5�4��K�w�L4(3k�zX�'K� �ӡ�()�@f _>�5��'p��H�*^���%A��]��'�@�7-\� <fHC�l=���
�'�40V+�;>�.p�KL)5F����'��A`W�&>4�0I�S�����'���'�;���*2�X�@���'��T�!enU^\(��O�����'aP��4ծ^�.h*u���9h
�'�l�a�@�G%���d�c*9��'���Q [(������'���'����p&0X�Z�w��(~�x�'�P���e�]�b��M(#�0�!�'/B�����#1�㉒4'��
�'v�	�b2BL%^��K ���y,h�2="�&M�)7*���"ɧ�y�E�0otJ)�@&�jѸ �y�b��?��]	�H�@C�� ��C�I7"����RK~���-xC�ɚs��x0�J��/U���-0�rC�I�]�8�03	��g���IJ�]$�B�?�z��77M��Y�I\��C�� R;XQ��)�*�)g�8B(.D��['��3��a -`عt`;D�d���K(L>�Չ����W�F@�m8D��ï��_.��ے�5 ���`�9D��V��@�ҁ��+�0(��!��)D��-��R�ْ����1�px	�%&� [`�m�P�ݚ���S%��	k���(l@h��y��v6Fa���qf_	t�d����w5��%f�	e�H��h��D �%��9�d5?�+0L�0�!����eb�]3L�HYz'�C);'m� ܦW~�%���u8���g�'Y��e"�&��<�aN� Ͳu�ד'�@u��@2n�(p9��:L4�r�i��4�,-��T".�����ǰ?� ����B
�)�'jC�2����DÀ3��+���b� ��  ��x�2 K?�Q�)�l��<�S��+ah�)c�-D�`���	L� `��&H�����7"ڐ髰d�u��H,q�d�?����<A`��b�	��[�4@�M�7�\CH<	GDi�$��剴R���a���)W]L��h�y^�T�O۞EրZ�E�k��=��
([My2&����T�"+�oX� ���L�a��EW[��`ys&�#8����G�^&@H�D��C8`�$�SKX9{U�}�-�=W�(	æ/߼�L���ܙ��	�x,��c`W�7s�A�w�W�e������(;~��O�hƠʜ_^=���P�9I�'ר�m��仔��p͘�0�۲�q ���<OQJm(ǌI�ժ��Zq�,I�y*�.[=T&]�@(�$i��[�PxW�]w�`�������wF��n���u�'XE�蹑
@+}l���-A&g�'YD��4�0��)"��� ��53�Ĥ�u<O��P�@�޴B#��6v�"�&��/�xm#� ȼE_�}�"�r�H��b(�7`���θW��`��*w�r�$C�d��$˟DP�[ċ������(Ol���a�9D�H��I2mqĹ��f ccV�Z��ͪ5��{r�ø�yR'��Y7Œq��Y�deӠb}�����v�NY�h]MT62fg^=U7np��U�4�!�y���\x��g��hNУ�%�p>)Pώ�-��u؁E�e~�)`�l!l�8Ӕ�#x,LQ��[ sǈ1�aFϰJ48�G"�fy�	(7�b� �T�3}".TJ<�rǀӘMY ph���g�'L|4�d��&��lp�N�&2��h�$�H޵"N���B�V�/.��A�kf�m�"��)q�Uٕ�V�
<P�F=�%�H��r�H/�la�i�C4j�YB�
*1�h�"I�D�j{���#�R���*�pQ��1A2f�iNT
���KT�2=t��RfB�o���zaK�?��?��3l��.�k����E���v��=e[ƥ��2O*���1i�&�'�[�o ��9s�B�-1l�k�	�n��ڑ'�b����,A/q0"gbƯ o�9�`�N�tFx���¦P�:��F�C?9�놓H*�J�ɏ�4�xp��ʸ&�~$��!���dɄ|�����	�����Q�O���ׇ��!�9:ӄV1 XD�"JۈzrPl	�a�{�����FS1h��,XV�v���w�ߨ{o8	�V� `�HT0�X����>i���$ƒa�6IE\RP8X��٭Ty�a�L�k�B\����6��"U�[ πA�F�ņ^W\3��Pp�i��
_��
�+&��/Q32�KG_)+��A�@�0�Ot	i�Ӝ#[6��c� L0y���E�"�A�%Þ?�lP"��$�`%��&X6���&G$Y�A��ub��s���`1�Wlr�h�,�f؞�2�"�/ǂ��4�Y�(#@��BQ#�� ��ҳAF`��ѢU/,[
x2�$'4=D��?)P��у ���B2B@l���B�̼�� ��Q�Bhb���8��>!u���"�R#�ˀ6�R�2�	/P��4(�BP)0��L0��G�d�^�#'F
ʬ	�@M�ahv�p��>to|�P��*�X��$�5ALry3��_� Dv�pP�aBH#D�V��S�D����9F�A4BJ~a�	_�G~�@�+��dM
lK\Q�W�
���냄�\���H$!xЦ����8L5���܈kt�X����S���`Ԓʅ@q�
rqڵ`�܁<Z�aA]�el��݋T���SO�}�䏒h�����/X�`�i���'��%"@��
��U���E�$�1Њ]>��1��$��QT�R�ĭ�3/�曦$"<��EJS��0x��C�C����O�i96��r���V�͓kH�I	�bM�8+���f��R�.a1V�̛&Ֆ��"��h;�A�焪�P��vU�<�G��4xJ��a��1  'e�~��E~��	FV���י )D����V��@4E�:ph�9��D�}n���	GT�����wݡтGX7N�AB��Lߌ�ɇm^��Q�V�پu���购�[��h�V�շH�I�F&� �SC����x���kb�m����5��x�@�6K�I���Ɵ�Ks�o�����D��� ̔�=���ң�,�O�|�c+�0�~�7�ٹ <@��@(�3:8��q��<p���cD�	�:,��C͡��m�3s �O�h�B�a�-R�h�6�Q���G
`E{�Ő/F�|�4n�p�,B�a�V��5?&�)�L0Wm�P��ܧirB�-j�k��MEX��A�/G��9�T�.1�^Tz3K��<���	$�qO��Vd���~�F�2���Qe�0|�9�PMƂ,�\�T��Y�<�3N��_����6N �E���V��\�w� �)�{��4��h�e�B mǐ�����y�횧wZ*0؁��U�88�G�B+��'�{�AU\���amɾt���fH�*P`����-��Ƅ��2B�d�B��$h����@2,S� O�ਢ�;j�q8�o�(	<��g���0�?��5�>��}�'Q�6_dؓ�0	Z8&��<�ظo3���� �,<�lIwn|�	,?�tQ��� �R5A|�uB��4�>���|,ޙqpiP'1EC!O;(i����¤s�C�	�B�DAz�扡Ln���2,�2=c�#?�F*�3F m�~�t�T�a���A�N�K�/M/'�!�d�:������%K`�;�IM�N���n�>uB�d8�)�g�? r�шˏ�Bd�4��v� "O �걍�;�ęc����  �`�G�|�dX<����ټ'&8��D�9@�8���e�=!�ٽ%%,�TB�<$�с��>zF���E"O�T1'u�B�K�k�?$b:�"OQz7�B�r[�Ģ���jLl��"OJar�CN�[x�ӷ��:�L�1"ON�r�cیM3b`t�P�藆/!�#X�� �6i�n�d�Q66!��ʦT��p�D�4"q*��؂k�!�d�;�f���
� �Y@T�?u�!�$@�*�4���&C(ΪtsQDV�rN!�$�VX`�C,S>,؆9�ä@�2*!�$�g�p��4�I��4� �$
?��D�3ZTf����0'x!��Oj�%h�'?����#w�,�)�jΥB,\ ��'g�!�"��_��ܻ)/^y�'OR���Gz@���7*$�	�'R`���ڄ=��e2���;D��'иi�p��7���u
L�;c Ԡ�' W�T![4T�b�SX��'�XU���XdЎt�&�-x
J-��'fu��P�Μi��ھy��d��'�����)\|ԱF�A�q���'�h`c�M=|ǄP ѩI�;j��	�'�9�3c��K�"` �ƉF���1
�'��hk&�*g�%��W=��	�'φDQS�C�M�h	�4a�=|.2�a�'<d Qs�_�D��ĉ��e.�U��'z���u@Ѣb0�U����^ 6X��'t�Z��WE�X�¤�DX�'b�-�%�M�)"��C���<rl�U�
�'i*5��!zV��,S���	�'�.�#�!Z(\�Id�]R�;	�'��x)f��[Q(y�#��ӎQ@	�'��}�n�,Y�ƈ��`S�rʌ��'l��hU��|S$�j��1n=��'�l��(�v�Bu;��
�ea�Hb�'F *ĤܠUf$tK��Zhw����'gh2�Pph.I0��0cd�]2�'����֯�.]���!׀	,[N�;�'�����4Q�45QWL�+V�@���'�0�5�To�]�ƧO���]o�<YQ�U$��,J�0g�n�	֮Ni�<9��ߺG	�Bb!W����a3�_�<i�-O��Y���'<��U�SV�<AG��<��yV'�!�Ꜣ�_x�<)7�	1QB��F�3zxp���v�<�U�ݸJ��aÄ�لq�0��b��j�<!��̽M+^#`�(�����HY�<E��,AB"P�%��o��e
���Z�<!��Dje�cX1:�Z�Y�M�S�<�	�2y�2�+�eI-�p�4�R�<��Kڴ��HJB#�(`�E�<�uO��F�#�H v�j5	�n�z�<���S�<����G��b����4�v�<��cQg8]�g��a� �G��s�<�����D�s����m��K��^k�<�F��?3�PHF(և:%�X�A�J�<!$� vݸ�3a)��hMj�.�J�<Q�#b�
@�"^:(9� 
)SA�<����1"���4GP�({hyrP	��<�ЦѶhΎ�0T�D4Or���\b�<���	-�h�ꓬȷ@����.	f�<� p�G �50�\U�K���"OvY����s�f`�� �/��c�"OFDs�-թ�%�R���=3d<X�"O \�d�2�����b��õ"O��s��	O:�$��a^?
N��"O4��G&�i�T�;�`�"v���qC"Ohl g��Q��u����a��d��"Ox1sr�֘?�|!��֓B��0�"O����䅌q)��Y�.A�?L�p"O~9�e��-#c"HC�o�1}��X6"O@�)7"�Ѭ]�Ԯ�1
�(Rb"O��Sd 7`��@�G)Z�HQ3�"O^��� ]1
P衹���(ߠ�#C"O�T�(#&��I�t햖nd�(�"O�ͺ�a�N �Hp����HS""O,�˥��0&v�q�M��Y�QqR"Or����T�g�x�f&tPX t"O�� h� 5�"� @��R��8�"O,q�3-�6I�xa�Ҭ>�����"O��	6�N��d�x��<��"O�ś�H�N�q7�ۣ\�3r"Oz�)Sf*~4&l �I�-b8�5 �"Oİ T�H�|Ў�A�h�1 :��r�"O|-Q��M
p�\j�aR<s+I��"O<�1S���p����V��L��"O���E��"2L����~�AX�"O�8kq��,,*��`E_�
f�R�"O���u)��A�8��DI �����"O���B I.|$�4�׃�
S8`��"OV�p����-�p�P�F;1�E��"OV�9��Ӷ@|�l�F�iH�S�"Oժ�EO	�.UI�P��.�C�"O4X
`D��[-�����Ơ,��Ic�"Ol��D�]���f�ڭ	Ă3�"O⠋���~E���[�1�zlA"O�٫���:U�n4�C�
.A��"Ou:Fο#�M��G\ -��1�A"O���`D�Z���C��P�n��4"O����γ2���%��E�$�z6"O�MHt��Rl�Q�
Y�s#Du�"O�p�B�xZ���*h��D��"O0Ir� v�* �6�:ٰ�"OP���-�SK���6���&u�"O�A�4n���2����S)�R�@q"Oz��A�D$}��� _tð"O4|�wa�m5ҁ����+
D��"O������1a��N�H(Hٗ"O���`/|� 	9��-�P"O"|���M?Q4	� ��}�����"O��r�,�4@�L��5\� �{"OFDäʙ=6�tɀ�l��8���"Or�Gm[vub����DI0!"O08 �E&Wߪ%j��S;Bw\`A�"ON�S�Λ�%�>�K G��h� �"O��B�$�>$P�L	�=��\��"O0	㤂�V$�qj鄁|Ȕ��W"O��
և��S>�=	s�Ҟ_�8%�!"O>5K`�M&i� �6i�����"O��1��	�%ʞ�ӆ�#:$A��"OR��*��h���J0�V�u�Ȓ"O|�1��'=ĩ��ӣp&@K�"Od� 梌!/��Y!�̐�r��*�"O"�X��*���EZ *�fhB�"Oލѡ��-,��XB��H�vt�9��"O� �@�Ʊ�.�V�L,{L��"O���D�}��I1 �=�ڄ��"OXB���=}��ks�W.2vVHku"OL)��m�8@�p��H�wT��"O��#��):����5HעZ�ve��"O X#)R�93��T�ح�W"O��rD�Eo��pň�h$QP"O !*�Ǟ�C�̋bDV2Rx�ذ'"O�}���er���ߌif�*5"O� X�Z`N�Y��%�	t_���"Oj�x��L=`��p�v�S�T^,���"O�!�+��<Z�:C�׍Fa��C`"O 	���ѬF��<Q��9/RL��w"O�m+0��S���OBjCV`zp"O,��@�B�-�|؅�٠d:\e�"O1�҃ɾA�4-����
H$舋"O�
�/������
˽���"OQ���l��	t�`��"O�%��,�K�9��Xp�P��p"O>-4jM9S��}+ >����R"O
!���		=���%�K�<E�0��"OZ	(�*��l#b�ʑg��"O�
����jaZu0J0��p"O�m8�`,E?0�ʥ�R�90Z�K"O&�H�MN�.P�Hy4�T=q4�}I"OΌ#E+A�[�F��׃W��n9ڀ"On�ɴG��(��`"�� s�d��"O��z�莫UID��d�|�@P�"O$��pK��R��,�i�`�&"OdM�� ƹ�%�L"l$�H�B"O:��e�K;u���狉3x4��"O��{��[�'��,W*׺s,2�c"OΕ0�ׯv(K�j��:�#�"O��+�Bʍ�	Αz`X�"O�dXtjI�~ʨ2&�JZ��]ӷ"OT�y�M]�Z9�ā��N5&��"Oj|�!*�+2���S�-,���"O���dy )_
��k�BX�y�M<�8�n��S�V�p�߹�yh8\,����r�JЃ��Q��y2��i8���ȵ$�N�d��y���Xqz4)��ǦJ���be�"�y���&<��/ǖKwP���yR�߰f��=�뒮C�<���bJ��y2K�@�TBQ�:�Vi����7�y"���]��=Z�o	)c�����y�+�B͒0��&�z��p�c��y�-��)�cюJ1"�L�cE��y�īX�2��¸aP,�f��yҫ�Vv�X�Ǘ�X	G�@�yR�6�XM�
N�A�X!���%�yB�ưf�JE��E�#D�F�ЁJO=�y3TB�Ej�?`v#q���y2��+���6`��sqI��yҀ��.W����&^�:I�P��,�y��Դlٞ]�B�5N��m��ϕ�yRė�{��-""��s	r`�n�.�yR&��_�$5:��X2D��y��cO?�yR$L$y�`A�J��D�~�p����y���15d�0�*��=�"!�P/P�y"N۲+�@�	��șd=��[E&��yb�b5"�9V@��^.!+1�y�G�J��+�/\|y"�iECY�C�	� ��!1��5ךԐ��A:�BC�)� t���,�|j����?����"O��%�>=ؤ��V$\,�2�a"Orl�n�$5�t�J��N:JZ�"O��"���p�Rv%AH�	��"Ov�����`ڒ`�N(&Yɧ"O����gXH�҄�؄|�.D��"Or��EE��d��)��١X�txC"O8I�����x	���v�L��^Ȼ&"O2	��S�O�$- ��A#� l�p*OhL����o���r����BϞ���'G�H!bCפv���#(��;��-{�'I��I�LH�2pԑKd��=9�
�':x1�m��<ElE+S�9�V<��'+�����­s��\9ff�����'��S%č&3�]	0萼p{$���'�J���EX�>Ƅh��e��q��� �'�ZCɛ7pT�"��˄��Y��'*V�I��^&�Y��g�0��t��'����%�̂\iB\�6+�	3�@X �'�@���׋O��lʶ���9�����'�|��w�G��)8f�ھ"� c�'h��ɕ�
�]z0U#ħǭyW$���'��UHp��/`��x��G������'E����� ?s&�R�Կ�^u��'n��2ER�n\"��E7
0���
�'j�${3N�ʔcc�
�J� �'�,p�S�M�.���E�;rf���'Pp�P&�ٮ.��C�/�3K�X��'jr]i6ȏ Z1X�I�Nt��' ��q6��7��)J��ɘM|p���'��!�%Y���"�o�-<�4���'!���LN�&��Q�'�P0�'����5'R���Ğ��|8�'�H��M0^��7���$X�'�*�A�9'�
���ߛ?���
�'��&厒"��Pꡨ�,x&�	�'SV�Jr'�$6���V�Z� 	�'lH�q'3\E����B�#W@Ry��'=B�2$N��9���0��p�TI��'�Z1�B9�\���B��}6z��� ~$!PM� �Xl�����}�����V#\��A#M�(t���E߻Qs�ȓ^'0M�@��	V �I����-a�	��<�
	{��Wc|�Q���".G�Ԅ�{�T�Y�d'/��]�tj��eqꩄȓ-�����,�/U\���B0 ,��ȓ2�t��Ӯrp�#�	)P�u��M�^��Ѭ�=
�,���ɯ\Z���ȓO�F����*_�ppV�C%�D�ȓo[(��'b��5Ӓ�y�CG!U�5�ȓc�`��!�+3��+��`$j��*����$���,��Ӏ�v���4��(���'d7��c'�Ư!�hd�ȓU����� +�@c��2z݆ȓu��(*�+�{F��&BzŇȓ6l����XZ�s�W�r����-I$|�D̓�LM p�gm ;����KŢ�ڴN�^ؼ��wĎ�<����"툍spD��	���@�HO-譆� ��L�3  Y��P�)�8�6��_
�M����MZ%�T@T�ȓ%�@L8�+Y��b�Qь��[����ȓm^�I �I��|?С�#)^�Z۲����Al�PpE��1 �4�en1D�� 1j0n��ydP�2�G�0��Y	�"ONYP�n_�R��+�+\֒��"O@"�& �)�
��ve�����3"O %;dUF0�F>����"O�T�T
k�)�D�ZsX�r�"O0h����A>�`�-s���"Oܼc'�O��f��9g���"O���bE׭SR>���▂ZI.�u"O�L!fa��b���Ѣ�B��&"Oƍ�t`��m=�ಠᔬ]�����"O���m	=q�jT���ֶ�}�"O��Xѫދ׾�k��
4�(��g"O�%R!P>���CR�� Q�Јc"O��C(ÆL��Qң,��_x|	"O���#ŌY 0q0���'e ̢R"O��iyu��:�C��.PZ �"O�|Q��48�������oA ��"OT5c��G�ju���!�DO��ce"Ob[�%!��)8�Ь>0��� "O ��d�8����A�'Jn$+�"OJuJH?FWz['N��2L�u��"O�-��T3X=�dU!"�"O2����0(��5H <0��"O����-�Jt�4���S�z�$�"Ovmɂ��	/"M�է���V��5"O��CB��?-��k��8��Y��"O����LF�Y��I@��F::�D!��"O�����@�
[����V�
Ɏbf"O�XI�#1/�03K���أ�"O�8Q��[��*QeA�rXi�"O"���E��W�D�ʳ�ڈcg�塠"OU{�c��0$ku�G0Y��8��"O,�B׊�$��ڃF:����"O�(����0<r�K.v4PX�a=�7�zH�lČ+�E�5.B��$�ϓ|7�`�Fl�3WbR��O� Eh=�I�mń8�?E��D�6��]'���$ӠH�ē7ZLF�`K�D1�nɧo��V0+����~� J+YB�)��M
Yv��p�(ҫ`���5�'Kڠ�u��'� ����f0T�9A�:h�Rġk�r�a�S�����ƈ!TB��	'�"jTm '{Դ�WG�;]��$� F�Dz�g�}t��U��П�Ґ���N1�q���/�����h��(-��\p\~��B�'�8D��Q>���O��iNU��)o�-�R�/��̂���:�(��ƝҦ���#}�r@#�����CC�<�L�;-��9���}8594D��0���}J|@��Q�&��	�]��܀��F-���O���ѕK��8�lІ��<�-cFˎ�$�r�"�Q	)�Xe�sK��f��,@"�(���"�5��0�b%^䔍��`��]t�Ĺ�cO3-'RU�Un��	�M�E�[<>��O��許 �9KyN��w��I,B̙A��
p����T���Z"�92a��_#t$�����v~�zC���1JW������@n�E���	�?7��>�2���;�
(�a�Ҽ82<���C����V%ypf��>�����6BM��H�e�V0JA�?D����֋?�x$C'��"z�:R�D0D���UkM1z�rt˗$�.sq�`�6� D�`���F.���L>��XA@:D�q0�U�gH蜲F���Y�p�8D�x�!Մ$KU�V�@�!�0t!�d�=V #s$��{��2����#�!�Ǯh$��r̖(AQh�C�M�!�#����F�%�-��ʕ$E�!�� i@��(1)G�5mHmҰ�Y��!���s�)�h�q1���ꗹ|!�$#*j �iŚL�^�X�K
�$!��I=!�����2.�����ϣX!�d��N���B�]��(��
0�!�G�EQ�`T1u҈{����|!�D��R��%� S�2���sǎ�!�� ���vJ�$[�jQH����G���"O���i�8�;WO��8$�"OT8B�5$B�+TÔ(�N��r"O���MG���#��9|���26"O�����0l[r� pD����"O<��G�C����_O�y�Q"Oq2�W�e���"r��4/�À"O�� *)��m��EK�cp��4"OP}�
_ww�1�o�
Pp`3"O�P �ҷu).)�e��&��D�"O�K��×3�fU�+Ww�J�Z�"ON����ݑzך	9�M�>2m2"OtQQ�7pA���֪��c;z��"OPa���O���f,��00�"O�XkBf��<E4�C�Kw���'"O�YcGK|g���]�^��!�"O,0���#i��8�M�n�bP"OP��OL�E+l�c3�U���"O��9S���n�����/>�T�$"O�� 
ёDtF�e�R�t"EPT"O��"�4Aޱ
�낓d.�9�"OJ��[��:D��&���"Ob�CD�e/Mh��L�
XN(X�"O@|8�/^���R�R�wT��2c"O؍ʦ�B�f}^�Ѷm������"O�< G�)!R"�X �
o+��J$"Oڝ�'@�9��I��⌵� �"O�$B�ȏ7b���6�*�Rˣ"O��S���%Ep�c���F�,x�"O���eo��<N:���R�1|�S�"Oʐʳ	�?��`�E�R�ul���"O�A�4"��]�tdz��1�:�27"O�42����Z�$�;Kҵ��"O�*�̌.`gZ��A�M*F"O`�K�%	�_`6��d��!L�m�U"OX@rDY	� �'A�޲x@�"OL�*�)�P� �/��X��e��"Oz={A�φ_.�1��V;I����g"OQz���@vRg��3v�f$�"O�U����H�E�k�|��li�"O:�Sq�E+H3��ӪD���r�"O`h���O����	�!|t(�y�"O����P�0u� ː!ocRI�""OTD����>Fģ��,(j��A"Oc �NWv�J�怵a�2� "OⰻV�Ӱ3�ҹ���*o@�=ۦ"OhtkτuްXk�F�*�{�"O ��eR,Z�)wf�bn4@"O��e�KQd܋%(�1I�V5��"Od��Ӌ0�v�*�H��m���x"O�t"�p7H j!Gـ1f�]"�"O�pXè��E�~E�t���'�j��|��'Ƹ����݆e��A�JVj-p�P�'{|0ٕ$�7+����3^����'%j@*̊kH� $��P���	�'���j���.��Ȑ0�K�n�0	�'-6$˗�!'��K ��z5����'�Z����΀WLjuH���q��{�'{:l�c"�9N3.L�FF^��P��'Þ�zd�tu��ud��Ap�B�'��q�NTeJ`т��`7V�P�'���(�g�d�wQ�RU����'���q�ǒEy[G���Aު�Y
�'���/�~)����\�2��$h	��� ��H���:OJ0ʖ�
gQ�YjA"O�(�
�0�G �CQе8"O~�۔�N8.��Zd�M�B1c�"OT[�`\?	�jQo��T\�'"ON��%�E(eH���@Ҡ=(�"O|���Z�80*��.H��܊"O��9�]�h���J_I��!�"O\��Ղ�%N`	�郒q�r���"O�y�U�X�=B�=��K?�n��t"O8 �&�F�A��:�ǣ\jC�"OF�Ġ��X���0��X2��"OzDQ$�.Oؐ(��EV��5i"O��AeI�G Z��&�(Ow���"O���šͶ4�d��%#PT���"O��G@�XC��i��εc����"O6�
䃊�}e$i�a"6#���a"O��t�=fS&�p��� ˵"O���6+�?������� )Hf"O�9ӓO�Zк�h ��8� �a�"O�+�iP�7 �F�ȩ�`К�"O����6Ąs���!�B%�t"O(�2��F�0���́}���7"Of 3b��9�@���,[��.�A"O-s2�]���"&�ӧv�x��"O��V��	��vI��[�p�"O��iDFE�&�p�?0<�a!�"Oi)��?|��`���9�t4"O�T+�Z�$K��QP���i���q�"O:�����v�q5̈�G�p)�"Or�HRaK!T�|)�"�F���T�"O䰙C/0�@MX�菹o��,&"O���/�&iZ�8t'����T�W"Op���D�E ������5���j�"O�X��!��.?�L��͕=���qt"O��a�Jd�p�K����+�`P�4"O �'���j�A�1G�)Q�rhR�"O������:fh��f�{�8��"O0p������Ã#̼\���"O6��ǡAqlcK��92e"Ot���m>PN���(�e�x��"O���7O�Y� 	W9Un�a��"O����P�#J�C`(8:R����"O�4�V$Y�D���G�On)��"O�@@�G�K����<H!D��6"O���R���$12�('gn	f�Q�"O�ʲC؁Mvf0�D(�S%�,��"O�e(#D8'o�AI��~�����"O�KV	Rw��[.�Y�fLJ""O���SK��[v�C���&����t"O�9ĂS�� ����#Y��Ab�"O�D+�B 9!̰▌�$'c���&"O~,�eI$9��� AЉr6d�2"OL8v#Pn �IP��ļ��@��"OƩ5m��@�F�kƮ �x6��`�"O�]��U/(zy�����dD	�3"O��I&�P�����%��aDԊS"O�x��,��$u1T&I�Z�r"O@u����%�	a�	�A�x!
s"OP��j$l���Ùd{�Aw"O��F(�O,�%����x��	"O$ ���&Dez��`	8��R"Ol:5�id*aAt�ț9���3"O����K0\��k�k_%E񞝘�"O
��A�(SEhՂT24��s�"O� �1�VA\�O�N�BlI0t���A"O�91w�OGtr���Zdj�)�"O�L�3kY�6��-����
Y(�&"O>�) IT�7�����	C/{XP��"OBU��*�$?�����.٢0(���"Ob��OE3�R��এ�K$
P��"O X��Ǣz^�xiÅU�|@,�"O��#�(�"C;��PC�D�� �"O>-�nͷ-p�c a�W�ܜ�p"ORdk"�Źw/��Y����"OΩ��!M+���C�ݢ2p,92"O,�ag��.F��#�+	-oL���"O�%�pǖ�E��y��KI�Gw�4�"O^��Gc� "���!���X��A&"OM��M�ZWJ��TGE�sNɐ�"Ohhd��j\��P�X�x��8�"OД� �Ў<�!��QMH��{�"Oq{�Ƌ�7����+,�4�)�"O��¥,I5=ȱ��X�W04i"O�I�S�%X�D���>Galu �"O�Q���EB��0rA0pZ�"O����Qx 2pEE,]T��"O�	JՌ�"u�%{�cʋD����"O�=ਕ�~˂��qB�C�"�"O& ��"J)MQ��Kဟ;~�鱣"O��B�B�x(�E�0�X.Qfm(�"O�xqhT�hq�g�:qB^�W"Ob+Ƭ3͈t#�&�:><�4"O�I����ڶ���D�-�fI��"O�%�2�Oli�3A�4Z U��"OZ9bG��A$��,�L��Y�"O �.����V Ap���ka��l�!��3d7*%@��_-H�	�CHƒ6�!�d1 Dف�Q(E'F���I��)$!�d@�1� 0Y#,�H�lp���Z�?!�d�0@\$�C˙�`�qB��|m!��1��P`L�/iy�x��JA�	X!�ߒ,�6��TiΥM�ds��ȱB!��Y=�t ��ӭH
�=����B!��W�<���J�� �=���,̀%�!��L<��Q�$ph���	�I�!��e��0A�ON�@�,ǝLP!�C�M��p1��$:�PXz��8P!��qE�c��H�.��,����2JpG:�t���B9�����	֤�I���3
�t�c��B��\L��,Ն<��I��{l�[�f�Z`h�ȓ3,2�hf�[��`�Յ�dr��èԃ�D��C�,%�ȓ;墀�k�o��Պ.�:~�P ��2\���lΡ�h�"p���|�bu�ȓVj���wh�Y+@iX  W�6=,�ȓKx�9`R&L���1���ȓZj�a��C9�����) <�-��+�qRf�_������C�g��܅�15�uV�Ā�ꭡ`C[*/����D2�p)��'wI�����$)��)����*R"qR"�&��чȓ	�R�8u�˘-�6��醡Ub ���]��=[�	�m�yжG�B��1�ȓbf ��-j������0��ȓM�Z�	��-�Dի���9q��ȓkm�51�[Q)LLZ���6+�Ņ��N�� @�?      Ĵ���	��Z��	�3V���C���NNT�D��e�2Tx��ƕ	#��4"�V����c��mZ�V�D3%K^�+$�ʡ�ښ�ePĩ�<w�����`#�Mc� Y!��n�]��i�;F�hxۀ�'���H��,�ڰ"�Ă18��pY�n� tR%�2�
dy-�!�dp� +}�VC>�*�#�SGt��֣M
K*��(�;`��X�'R�D�C����Y�*O!y"���`���_��[6��)*-��-���pۧd�m��=Q4+C���ɶv#�`	IE����n�ن�ȹ	���Ѓ#�'Q��<���A�'C�$�fl����f ��L�D?	 I�U �Y9pH�'*	�4�B.�e?�u��~�,PH<yË��|BH|���U�9����C��;taN�R��=[J��)Y*��I�'ɐ�@FΒ2��I�(�T!��Ϙ ���pː0tl�P�4@x�I1�?��[�kIH�$���`�oWtʓD�$�Geڡ:@	���6s��ɢ��i�G$7��ۂ�K��'F��"cB٤F����/� Gl� ��ɖ"�'���T!�
:��OPU:F��"�&
�#9J�Q�H�<��� AOʶ������ы�U���Xx	�g�w�P��4.&`UEˁr%�p�4��������)*(G��O�j�}�|	Y�a�J�	��?���"	��]�rgւ�$KW� �o�4�BF�:��`�ڵ�֚|b'�l���H�'\Ȫ�FC�ʌ0���D��*+O.�0�^��(OD3J<9W(�u��Q�G@�=U���a�Z?o=�
@O(�!�4-��ߕ+"�3GJ�k���/R�q�Q��`�apX���-� �'�)��`W�/{��dދ�4����.�6D �N&�qO��M<u�E*�D�M�<
fN��t���� �^=�LX�L�A׾S��0��ϡ>1�9�w�DУ~"�a�g��>s���Rb����U�,D��A��   �� 8�Q�Q"O|(���  �@ d  ��gb �  �4�[���.�Z(���;r���I+�Qf�'jnIa�[�?3��J���M:V���&V����;v�y� H�o�I��ß�ntd}��wIb�z���|��,I�ks|aG}C	u�O���p*�2E����c�MQ�:�r�'2��H���`��b)HP�0�h�'F��5	�YiJ2r�ZE. ��'�1�v��p�+"Y+ST"p*�   �  �  A  �  �+  �5  R@  XJ  �T  (]  ,h  t  �z  S�   �  X�  ��  ߚ  "�  g�  ��  �  2�  s�  ��  ��  =�  ��  ��  n�  ��  ��  }  �  | � v' �- �3 "8  Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�� |d��"O
`�(�;���8���-0��1%"Oj4��ND^[��"3/9�0|H�"OB���H��*�ʞRy=a"O�味V�!X��!&F�:J�$���"O,��a
���C�Ą�M�"O,$3%o�-���p���+Ն�:1"O��ݢ1����`���y14]2��i�<�6��{_���c�H�`�fX�$Kn�<��A̼VI�xR[�)�Ć�pඤ�ȓA5��('nߡ4�� �)˩%� ���,��r�؊b#`T�eT09���ȓ!�b��g��}�8�F��-? �ȓ
K|m�ș�VṔ���2�%�ȓ"R�X�j�4JN�1�˘X�i����̹	_�jZ��1!g��zܶ��ȓgil,*�J�
j�Ne��i�J%b���f	�(U��:���G��$Y^م�~r�� S�%T"���k\�jx�ȓ|4�1�îJb��@ӵ�ݩn�V��/[`�"�v4�R�!ʎ<��M�ȓ`:��z�ؚh�J�Z��$HY:	��H��p�m�C1��!��B:��0��EnjZA V;9����J[
2���	��4'J�EA�IVW&��~�(aZ��ӹ�>� o�Y�|�ȓ�f�A�
Ο7�H��M�$�����mޠP����/���ANXo*�ȓTv�����{ ��-7�*h��I��sB�8�8���3����ȓNe*M�悡;������X�o��!�ȓ'lj�#F�m�+R&;�|��2)n�C��0S4���T:
b���:�0!��e֊��)��ͷV��,�ȓ0�&�8#���� ع�L�����;�P�AFd���,w�6d��r�EQ�( �gVlɦ�M,H��,DP���|�I	$G#\���ȓ"�)���E�B	yt&B�^�LɅ�4�� ��eëF�ڙ��n��R�p�ȓp`@}bŇ�=�$�AUN��P����L��p���_�a�)�Y�!��-��u�5���o}�`iF�@A�p �'Cў"}�ɃJ��ӗ��GT��DKKv�<Qb�ʚ\���'$�QI���M�l8�xS�� 3�L]`#"��m�d���$�O"1��}t��qș�A"F�2�Q1�9��*Bh�4
�=#�����A��]�ȓ}�4t	$e� z�`��՗f:�ȓ\����!�U<Ed�`�!K�fVI�ȓp�Llk�%�$h-�(�e�}.Q�ȓ�@!xdOZ�Zn.��!�Z
�:�'Ua~�O=W� q# [ 9�r�������yRjK�U��ᄌ-2$,-����y�I�2�[k�!-\��"3�y�&�1��e�a��*r&qab�E>�y���
F�:�0���q�܄�!$ԻIj��=E���`0ze+S�h��$H�w&Y�ȓASN�5a޵�$��'��\����3[�)��G�מ0���r(Ȅȓ?5t����һm6�0ϝ�f*.��ȓ)����`E�	&��mBS�v`4��S�? *8G�#'��v�^15�\��w�|R�'��T;B�I�%�j���'��M��'0����*��0�0@ `%0�����'l�@�u�N�`|�}��n�%�X��'-���@��5�Ж�[#T	y�'�ư��!ȧh�J�����B0��'	f`H��GM����o�:¾1��'5^԰�%A;t�A��wZvi�
�'!l�iT�ݧ7?�i�	
6p��$���(O`E(A�V���+��ۂɊ'"O��e�@�P�X�S%�F)<D���"O���	a�-{D�[�Eέ���'I�	 Cd�!c��0"��ʀ�x��C�I8�h���ڏib��9sJY-~��#=1��T?��wo�+M�2�8�l\�2��%G&D��bӈ$�|����z���`/D����\1��A�*�|v��(Ԭ(D���5�Ɲ[d�)��ԩXE��Br�)�D9�S�'9�^����bk,�}�r��K�<!�$�92`h+�UjATa9���J�<��5s���I��I�R���)��|�<9�̆x�l�kf"�ν!Fy�<q�-�(
qI�I[�P�^xY2��Y�<Qt��3���V<X���҃�Q�<��$O4fm4��ON8ldzi`�.�N�']�x��%>
k��]�]��H\��yrl=n/LCw��8�Je�����y�ʞ�a"�@��Gy�I�Wi[�y��>��J�/D>]�\�('��7��d7�O�"�nL�[.��+�k��U�b����t�'���{��IjE�̭R��P��ʗ~8���ȓMc
{���>p�4�C�B������	v��?���.B��h�lG�P�����S�<A�m�8PHr(��@G-o������M?Y�4�hO>;��U�|�8��4N��`��ݛ��"�O�Oz��ㆈ5�&��hިBd���"Ol|�@O�kW\��!+6G��u�'/�'�xPp�X"}j�3P���,uz� 	�'�p�$ˈ5C�!�4d�@���(ORT
��@.���*�AQ�ؐ��'�"�I-�.�r��BXl����/� j���OJ�=�}�$e
�6�H��C��5;ڌ����o�'�?�b2�(o�"�h�-=�͢Pc:��gӾ��$ώ *h� FjF�YI�Y5@����=E��']����ˈkZ�|㑯�MY�!��'r��V���\�ڑ�̺v�jP`��i��~ҡO�{1�x#N^38�20ʙ6�yrj�3f�uRCnK!���`�,�N��<{T^��F{�����:%����(ċz�	I��yr�-���n�S�;l6$ 1AA��x(h�NOT��C�I(sAT�1R�Q�
L����<�㞈�D�)RL�,
e�qX�,#S�p�fF�#5&C䉙DgB���X�<UൂfI��>�E{��9Oܒ�EO�PZ��1�A�.d챲v"O�� ��$��,3ǏD)?<�V�|��)�	"! rFڞ4fz�� ØuI�6m �S���ě�&� �Bqh�%B��1`ϭ.!�u݄��wfY=�p���� 2M��w�'D�����̘�?^z�˕�G�,� fJ&�O��'��)S�^�\�I��*9_�%�	�'vf�{�@Ȃ=v�DV`V�<�^���'ԀmHd����ɒ�ގ#����'H��s��Bs�q2���Z�r� ��OJ5�
��3p�iuoJ:i��������Vx�� &�x�XQ������?9�dYs���:\O����O�IQ�x�����h��q"A�'�'�F0�טM�6P��3j�h=`�'���@:`�9cO���E��'*�tc0%Y�t�)���4�Px"AE�H�t0g,��b��G���M����?E�=i'I�.�|L�Ѩ�,'�Nh�!��U�<yR�ˬ4vnu�3��*R��Ak�a�v�<���D�<|	8e��'(y�9�a	Dt�<�SL�-�B���ϙ�U�b![Q-�r�<apD�|舘�BIE�2-688�HJ�<��ʙnx�5�F� �N���Hz�<��'ɴ'&Bi9!C;e7ҹC�M�x�<QЦ�7rr��͕4et\5�1���<��\-OD�A�/�2&T�����Zg�<�#��4%p�pR7f8��^�<�qꇔJ���kP̊?FzT����]�<��a�qsn5�MZ�98��W�^X�<�����n��5�$��Ep�<!��Ԡ%��l��\?l��a9�@�<I���*t���6eO!:¡z�i
.C䉸xࠥ:��O�9�p��$φ;1�*���O���b�O��D�\�@aFl
)e
�aF�!��P�@���W��ap��&��{��K}��)��IK�8&��D���z;J�4���hOj7�+�Z���i��v�!֭�3HbP�ȓ]��a�+аJ����hZ�h�ȓ6�V�pg�\~�����;L"����n�@Q�l	� �PH��/Y�.�<�ȓNF��'bѻ5�t��Q�I+g�fE��)��w�����B폣+c�%�ȓOa{�n�U��L���69FD�ȓy�l,Clks���"@ȝ����4�����K��I��*,{�хȓ5h��Q!(N.I���s�Y�?	\نȓeB!�%��;* ڡ��,�+,k���FoJ�����auOP)c��ȓ:TX	�'U1O��"Q*P��d]��X	�����Ъ�\���*؉4�؈��Ц}pb ղ{�>t����0{Q	�ȓ �v�+S){4TQRȂ�*q�ȓ��@h��  e�z���,D�b�$]�ȓZ���@:(>��f&�q���ȓj\�y�&˩a�T����8����qn�{�ȱ[u�J���/a�ȓ6���{g#�7����S*_ղM��U��A ���,V��*a)�>����y~�ͺĨ��csyj� Ԓ_R�ԅȓU�BD!�J`��e�v��@��ȓ�=�GQ��=��c� �����Y9R�s�E�fl��a�9D ��+B�I���O������N�9�^ͅ� :ƑC�T�<x��q�S?]\L��`�Ƙ�Wꆪ8��c�	:v�\L�ȓM��T�n,OZ�
�e��rWl(�ȓu`8��zr��!��kW���ȓc�J��џi2��2���"�t�ȓ8o Pc�	*/�)`�,�p������lZ�� <�p�͐u�<��2��qQ��%wK�ի֧�'?g���ȓdu�E�,]�6L�C^"&4Jh�ȓG���%�ؑK�T��ԡ�9���T0p$c��	#C@����n
'�X$�ȓ~;�I��"|�z�GT5����S�? ��+��8-x�@�GT	b��#P"O��Q1Ϛ�=!�]c�+#�p�ȗ"O��"������)��mw�)`�"ON<`u�(cȌ8yG�)f����"O��e@�L((i��w��Q��'��'���'���'_��'V��')��SK�QCTJu�''2-�V�'���'�2�'���'U��'��'�B�@�ᅶ^�hј`�V�ɜ5���'��'�"�'��'�r�'�R�'dNi����P�
���t�x����'�b�'e"�'q��'���'��'�JM*��݋1�L /ݗ\%����'V2�'�2�'r�'"�'c��'V�� +8�pL�'F�٠��'���'���'jB�'L��'<��'���˅I���*�hdD�6�'X"�'�"�'*2�'���'-r�'8 ���[�U�ZqiS���XA�X�#�'B�'�B�'5"�'�2�'K�wzTR����Y�FM��	s����6�'���'��'��'b�'���'�8DS�NY�}Z�-y����A'�QI��'�r�'�"�'�2�'L��'-B�'�$��ʉ�I7fa���M�5���'���'�B�'��'��'r�'��y2ċx�%@�ůQ�Ba�'�R�'�"�'�b�'nb�'���'�l)0�ς9ԴX�D,�xS�'���'���'r�'���d�\���O��
����| Y�)�����G%o��Iҟ8������Ѧ��#i�2�잹M-*4�U�ئ_�$�Wٛ��'�ɧ��'Z|7��s(,hb�,u��j7F�JҞ�mZ���d��Ҧ��'+�%_1\���ś~J%&W8� U:��>cV�!�`(	v̓�?�(O�}z`@�s��2��;8or� �"H�$C�v_���'�X�mz��[����"z��q"�P�0e$Y�MӢ�i0�d�>�|�g�	��M��'%BC��ϛ*��ȕ�O��*�'��<�R�Y�`��ea��i>��I[w���%�u�D����wb&�y�[��'���ܴEb*,�<�D
 l�tY�P+�t$h=ӣmK���'20���f�v���f}�K� ���#@m��>r`��q��-���߀3r\�pp��sp1��� ��i��	�X�\urAN�',;*����1xj��-O�ʓ�?E��']2A����d�n���oB?m,�d#�'�
6�ԍrW�I��M��O�yR�Nĭf��e(rZ�h@���'/F6�����Ɇb>(�mU~�Zo8�S@��3%dr�(g�ѩNp�-�q\��iV�|BX����I�T�Iޟ����=_�6!�,��B�&�Ay��l���:O�D�O����ą�2$�d�E
.Bʾu�@�	)����'�87�C�}�I<�'�z��4������^$#�L�JQ��.S]z9�" ϏF�2=r.Ou�Ԃ���ݣ�����|�.�x����p�P@Q �;=�8�d�O��d�OX�4�^ʓ>1����ybk�I��I�蘢x�*%	J��y��i��Tk�O��nZ��M+��iٖ�	�%
�[T�|3�c)��U���(L���:O�d��:��t�G�?�����V�A�2��� D	�\a篈�~��\� �P&j��qN�l��8	V��9d�5x��J�0���	�K�f�	'+/꡸U��0�*��^K�����F'*,���L� �䬊S��}���0*As����ˡ.	(�������uK�<��LJ���U�m��(m+X�"u&ӟrf�`���4�T��m .\{��'g�`�D����Ҏe�n0b�$ԑn^~�&��>����nK8qd�mk �Q�vXl� �U�Xgt�{w�n���$�Od�dX8a���%�����|��1W��Q/�0?!j]��.,5#���>Ip���?A��?A��ɔV��a�-��8!:5	��������'�����H$�I��h&���4h�xy1�Iǝ<�n`r��L=8��Rj�p�<����?�����$��l;��!��#\�1�O�"�&��Cy�IҟH��Ɵ8�'H2�'"m���8i���Ac�!�(��E�7Ϙ'�b�'h�X�X8%����t�k������*sVpA�)����O"���OJ��?��6��O�4䊇��d�����Eē�>�@�O��d�O��d�<��#k8�O��@�%�`��ek���6I��R�Mw�2���O�ʓ�?���E�V�~����g����Cɔ�Z���@�Ӧ���؟��'�pq��+���O@����Q��7#���Jяޓ7v�j��i�	ʟ��I�p"|z����ʌ�`�Јp Su"�B�h�\˓XnJP($�i����?i��6�	,i��ܚA��Smn0��1y�7m�O��dX����S����ēi�$���C,{�!� ��>}Z�l�(�@���4�?i���?��'�������i��@[��,a�q�� �%�7M�66h�ʓ�?I���<	�@u~l�t�g�zE���ܝ'(�y��i���'�r6�PO���O
���	�=�q�Z�q�v�D��'?��'.�e[�yr�'0��'��ڇ�X�8єΌudHX�4�p���DT*3��%������IYy��ͭ����G��1�Lq)ði{07�O��j���O����O �?80l2aEJ��  ���zn���"gU�'�b�'��P��������tb˕E��"��K�^aP%�',Y�b�L����I`yR�^�\v�擎y��i���,|�` ��QbV���?i��?�*O&��u���4X?��%�}I�=���A�>\���@!�>���?Q����䖉3"�<$>}�� :�b��{��d�S�#$��`7�i���'��I��0�	�K��b?	�`�4-�i�ݞ-_bxbb�|�h�D�Ob���O� S3�S����IΟX���?���B�Q>���쇍c����*��MK���d�O2�@�9�>��<��A@cf��+PF�����W�v�'�-оRk\6m�O��D�O��i�t�$�:H�1*�-0,� �s�ڠCk���'����s�R�|�O��'��s�)Fyő��\�[DN�mڴff��9�4�?y���?��������?1�[����,��%
�5s��R^��YѶi4l���'
bZ��R�ğ�zL���AƁF;<,�QӓNH��M���?)�h]�I���i:��'��'�Zw�A�WJK:}x��rm�/Z%P���4��d(Dt�h&=O�S�?��I۟D�g�,�\����~��� K�<�M���	�`�Q�i�R�'�"�':��'�~�l�]5���##��v�ibu����H1����Oj���O���O>���O�|�b�5c���D��v�@�>�m؟��	꟔�ɚ����<!� ���*��Q a㚴v,��
�<����?����?�����)�?Ӧ�n�v?�h�2�P�	�Ыq�D�"�R�4�?����?I��?�(O(��V)e2�i�5ꠉ<v"��CmÄ s���O���O�$�O��/�8�m�ğ��	����  +��O?��R�h@�b�n��4�?1��?�/O��	 6���O��IJ��)��˒�VY����O��6M�ON���O�$W����o���������뺛d��1��]�V"f91ԍӮ���<��VFP�ϧ�?�-O�i�h�+�'4-�u�ME����ڴ�?��`�N�!��i�r�'�B�O|�4�'��5AV�{M�`)��/�p�Ƴ>a�Y$�Q8��?�(O�� ��C=�����P&�:	�BK���MK��U��F�'�r�'��ԯ�>.O�i�'b�	N޽�(@�A:�A���˦�$K!���OUB.9E�`
�*��D���1��8�>6��OB�D�Op�@��Ǧ��՟��I֟��iݹj"�!+2�����v�>%�
gӴ�`��\�B�S�d�O��'S��2境 �
�Cwň%����UHy�L�䝈`�^mZ����˟8�ɯ������իQ�b=���w䐼w�^�GM{ӄ��#�/��d�O����j���O�˧h�Z]�Wn/Gf��􁅅]����R�б曶�'h�':���~�,Ov�d�"��		&#߰=*��ȁ] ^9j@:O�˓�?a��?���?QD�#���Lȃk����@��	r*�#a&��zZ7-�O�d�O��d�Ol��?��&��|���V@� A� � �P#�Cɡ)��IӟT���H�'<f���=�I�`C�,����R��!�B���,@lZϟ'�\�	ϟ(�q���O����H3G=����l�,*H�ŵih��'�割puJ$[O|�����ΐ��l݀��;����`�dP�'v��'*���'rɧ�i�2����ëOլ��4 $I0��R��CO�MKS?i���?U�O ���
ih�p^h��1��i<2�'`B�2�'Eɧ�O���� �/L7�@���b���4�����i8��'nb�O�0O���ΆOW�(j@)ϐ��|��/;N~�mژ4-���	Q�)�'�?Ѣh��u���AQoR�n�R5��ؠ-d�f�')��'T���4�,��Oj�d��0��U)TMB�Dɕ�G}��t&nӔ�O*���L\�S����˟<C���%j�ЀoW����ia����M�������b�xb�'p�|Zc���a�B[+�llڀb��2>�1�O�@�0O��?9���?9,O��`�ꔼP�2��F�9`i��L����'���	��<%���I��@���+����V�r��=��NG��%�$�Iɟ$�	Zy�,��3�
�!:`�
�oŽ 6�!��n��$����?�����?���r*I��0�	�b*��WB9�CK��J�r���]����ӟ`�Iy���!o�n���Ҡ&��=&��d��#�p���a��z�I��d�	oƊ]��[����Y�Nyh`��4if���#ꋌ:E���'\2]�ܹ�����'�?���Q���NZ2[��q��P�� �%�x��'���ݖ�y"�|��D�p����A3���
 �Ⴒ�iO�		;v��40��ϟ �����'c��H;@�ԧh:p����#(ϛv�'BHB*�O���E��b�y�vۖ��J� ��ּi�:1�t�����O������&�D�I���d��M(MXA���6r/�-aٴm\\�����S�OL�+�+U�����s�t1X�j[#9�T6�O�D�O��P%�IJ�	�,��W?�PcQ�S��z�$�*J�ֹ�%�_��f�}&�8��ꟈ���V�=�wK�&'Z�`[够2@ne۴�?��O��'���'0ɧ5�A=!�f=C�`��{� x�Ę��$ć?t�D�<����?����Z+;x��s�I��b�Ȇ6ZKP���F�I̟��	I�	̟����r�^�`G����d��L#bwxX4�Zȟ��'�h� �.��WV�a��,��oX�ϕ-��]�5��rT)7�Ֆ$�99�
ƪh��v��_��	�"�Ԇ)����H���O��!�]�F�}�Ъ�>%"\ac�K����N�t�z
�艁_���a�I�̹�#K�ۊ���)�b��"��H�,K&4Y:���
.GZ�I"&F�*�Z��ĝ>���H2%�*~J�	b�Ji�^p�Sc��|4�Tk�Ŝ.?�  �kF2)�iGbֿs<.-c D[�p�gŎIJn��H�
c�	�!�t��P�­=`���6mR��'ՠ`��ƣ^���4�D�!��9�S��~�/��h���7�\Q;��q����e�>��B�;�j�J�i�:9B���+�uW��8s��!+�π j`k"D"2rl��j�7E"j�A�>���۟h�<��Qi��]Ba����&8�l����Y�<����!�($(���C� d��)�X�\c��D	8$윑G��;m�x�R�� {��oߟT�	�� �%��=J�8���ßp�	Ɵ�]&m��5���3E{Ĉ�D��&;ъ���V���0k��l+���ӫf�g�i�L�框� ��x��H�a����u�Qm�����<��	��̄�Y���Oʹ�1Yռc@5o�R����ߎ`�����E�&�'�����S�g�	�S����И;cz�H!�\>JV�B�ɆFќy�ሺD@�*Q#��i`��
v���Sn�� �r���!�e	�>H�N(В�
"���O���O��U̺���?A�O����_1SU�B$��3��+ƃ�.�x�/R�J@���فvٸ���\�`�r���'G�����<Q h�:'B�
�]Z%���?��'nTHj�˚��B �e���;I.��'��)@$��T�N ¤��?�tj�yR#"�	?a��O��X4�(��D
b��J0�D�bm2���OX��O�Ol�$>�����y��9K���8Rm.9l:�j���X�Kx���D��`�����Y ����*4@�Ѓ!ebӂ�HF#�`N5�Q�Ȱ_~̄��'uz����?�*O�aP-]2����"C�la�9����#�O�Ěr+ܴ"���g�;QG�1��'7�!pf�W"E�r�@��D�Y��D�<�s�����f�'��Q>m�2����l�S숐t����b@�s<��K䟈�I�>Cބ8��ܧxD����?�O��4&�2%P�����U8g��=�r�'xhu�sΒ�OyU���ڿ�d��ė�
��a ,�$q���_f�I���6TbL]� �>�"�ʟp�L>��g^���ِg��N\�3�B�<������-|�8�B�C������$H�X��e���Ʀs:��z�i� d�� oZ����I���3WFR�Q���	ϟ��I���s�����
�U�n�VݍvQP��N��,� �`��O�Mi�QA�g�ɁYp����|�z� ��C�HP��G	/�> �D.J�A���f�2+��O��ŉi¼[���)|�̂7 �5k�8����T�5�'�0���S�g�	�]t
�[�Cխe���8 �ˤ'4�C�	Nc�t di �]ҨCFM�9��Sԑ���z�	%�&P#-�2Z7
\�@�6A>��!焎K2(�I��0�IΟ_w���'��iN�%�y��ZLbGA��rb�`QOp@�=)l��PaѢmF�b�BSc!��<�H��XG��j�@�,Yנ����'^����-�1��l]�gޠl��o�p�!�X�}jX�0a�S�fü%�a���a�1OB��>٧����v�'��#JE���:��& i��l�) j��'���!"�'��0�D][���[A�|��C4R�\t0$��0c���7��&�p<I#�͉xP$�(��*ů,8�EY�$I�?�y���+O���V�'�PO�ᣡf��Ĥku�Y�jv�y��"O��"�{��� ��ae,���Oj-mں$|���Q�]�!Ly"`�E֩'� ���6�M��?�+�����.�O���`V�Ba��ሜ:k�hc.�O��$�'� ��'�C �(-z�����'��ID4�R q�l�:o���S�OD�(�V��aj_B�!�$ޕ~	xc5��}�<)zd����M_�;v�Q��/����P����0_2�D;�)�S�~В�H�ő�no��Y�. �3:B�2	� �#n$�ȹ��B8����a�'�v܋q�Ɛ{�1!W.�v��I�Ig�����OZ��L�%����Pc�O&���O��4�樛���=:bH�%n�m�`�#�gã^Y"3�Kݦ��!�Z�aW,ȕO0$b��ĉ�N4���� XzҰ�U��4N$D���5fP�	Q�[s� �|����i.杰b�6��q.�$;@�zr���;�H!�4&剓j4���O���L����=���-,K"���4
��4�T�I��hO�S�U��CV�݁
��H�������;�� hӸ�����I�?��E�t�'�,ዷ*7/��Q@����Y�~�ɑ��z���' �'�.ם���	�|�s�w���ɕ��6Z���J���E8���b�>pkAnD4�Z���3����Y���?-# �0MD��6|1�Q�F�
=��j�O�1m�;�Mk������O����;9�ԛ���s�Y�
9D��R�KU
5J�P���W�yA7�I'�M����d�6S"l�ҟ4��$'�N���'�R,�E��[EX}�I͟��Ƭ�ӟ����|�f��h예x���[)�EKٴ	*Q�0�	2�|,�c��+EZ���	� H�ݒS/FiD��y��aKE�G�k1�9�bȎ?&�y@���9�sM��W$���&D�O�%�� �-���JeV�s��� 8���"Of|r%M�18�JVU�#��)c��{����lӦm�j.�x�X�.
+`����A:�$]�+��n��L��e��eާ�r`,@��P�RD��ZLp�D�}B�'UJ����U7�ҟ?��)��S�T_>qK
� #P�dK� �0�X�;#�*}�(aD-zt$�Y��:cf�
[�t� ��7D`�̧���;F�l[�bI�T�h��O�E���'74�O񟮬"F�^�nl2��U�b�Pb"O��c%�մD��Б�2Z�T���'PX"=�##������ e��D�P�(83�V�'�r�'�|ى��U%��'����y��Ӣ	0b�C�'ַ$7$1ruAN�4oؓO��۶�C1��'�h m�:"�z����_w��$�� �^����(��!�3���
������G(d:����ڨ&��d+?A��[��>�D�O����Z��Ȕe^/T4p��g�/7BC�	�j��t��a��g�rt��O�p��80����$F�J�8j䩔0o��偲O<�k��?6�P���O����O& �;�?Q������ɮ�\ �U�#@U*=��́
)��M��K*l��s7㜫D����ɻ�<Ę&"@�ui�D	�&(�Ų�B�kg,��c�O/x4��������K�%��$�I>��K� FC4��a̜�dJ^�8t'G�Q���	(�M[��i#�O�-�~ڵě�P�$Q�B�Ԡ�qld�<��ێ5���I�)
�]*L�)���{�"F�'��I�.�(��4�?���7!��$��yG��ز�C�X�������?y2c��?���������3�|���G0o�nY��'?vC�0�G�?���R���=��X*�BZDFy2EH?&��u�1��^�[�DԴ�+gV(9� �@���P�(���O�UGyrg[5�?q&�x"#!�2�`H]#8^�1�ǜ8�yr�٧jR��QϏ�
PMi׫ŕ�x�f�iV@ͼk��"!�t�0!�1�$�<t�4mZ៌���D�b�� �C�A�Î�5p��<�2���:R�'���b,�;�7�t����|+�@�{�k�Z��Sr���Z'�t`��>�Ub ;��@�Ä�B����2�R)�ug�@-*��X�O�k�лz�t� �E�#�H��3�*}2����?I�|�����&d"ܡ���$O�.d�Q-�;�y�j˻&~F�ɒ"�2J��Uy�J���0<	��/G��Z���}@y���B�#�H���4�?y���?�U�1m*N���?���?�;9EP��c+"$}��
r�%@ұ��y����<	��c̒�k���L�T�yP��d�[���牀i��`JVd���	6䝃�R��N>1v��>�O��%N�O�:10bِ�R0i1"O�����W��]ӥaD`��P�V��x@��4�D�OY��$�0EK�Ě�Fr��8y���O<�Y��O����O��D����?!�Oƴ� �~��|9��դ+��8ZW'ޥcH4�A�N��3چ��!�'� hvL��jG�����U���l՜U���J
���B�)+xQeʙ�@(Lh�=	�̌� ~����G]1��z6M��v:P��ƓZ~�EQ�n�1"��p�s�ʁ9��	�ȓXo��ف��n���,ν-΂��<Ip�iZ"Z�dP$ ��M����?ad�J&!Cv\`�c]y��/�?��z� Y���?��O�Ј���w���@�
R]U��x�LU�Zt��I�xz��d�w#؟
v��Q�-D�S�T�ȓ�4O(����'�R�'��hةw���H����"�AB2C��I�x�?E���-28^�����;rȣR+��xB ~�,%�*N/��u���B�jj0�3r��O��v6�\9Ծi���'��L�&p�ɒ`�U�bf"9�� z�� h��I͟`�Ao��t��k�R����q�W<��)�|J�CN!H8�D��+��Lx��%)�~��)yC�LT�� m̴T �
�2:p��$�	5D��ڴ�i�őS�@�\<KF7'��SҠ���m<N��I���S��.q^�+� ��@-2��d��m��ȓ6���̚O�*����h������4��<Fz�O˧�	6��"u�0P�۽�6m�O���O2���g�?����O��$�O�NC:e`Q�!bݮz�4���	�wh�<Rw��(Li���A�o�R 
�d#��g�Ɍ����^�CoXD�GO�;!�p�#T�a0�I�k���#���?�*�O��V�Γ�ywN�=WHl%:�AS�#[�AaUပ}�2��(��j�Oq���'�RD	�xdDt����-#l���lގ&]���C貉K�O1�(�`l�$F/�I��HO�i�OT�`�L���U�n�+�d׵Db�q���RX��R���?���?����B�d�O.�� PP�'��Xb��<������� O24����M8A��Z �E`�'E�y�&��}=�6���"�4� J�[�$��%��^Dtة@]�R�џT�.ͨI��耀GctU;�M�Y"���'�O� j]�VnH(w3�Ux�̀@�v���"OX3g�[���#�S�������Φ�%�����M���?id�2$�N�1f�q���5ϩ�?��& A���?)�O��	�R�C��@���!t�`���	�(|H�����8񆕢cџ�3�\ R~���BG� `��C��T4 ��j��ᄑh�	n? �-���4�I�$�X�ɫ$6�2�����4�V=D��C�ɀ(�4�+
����y㈈.%Z�B�	?�MC��w*fy���V��g����Ba$U)��iC�'��Ӣ����D��k��i2�\0U2v�u�	���e�S[ЙrbE5%�1��T���)�|�c�Y�s�Pu��5q&��w`�m��f���)�<}P�
� :E�-�;q�`�F�55�դ`���RL�(u��E��(��R�ZQ�I^�S��Vm���#�b��Cт�D] E�ȓ�f5#�THZ���C�P�����HO¬��!@�rʆQ�ҌgG�E���ڦ-����|��%1pt�0�$�	��i��HF�V�鑆��ITd���M�j;���牻	�@� ����i_�H�Θ�"Z�8�J6<O�УAc �4v`	��U[}P�4BD}�Y}X���|�R1-Ք݁�O�Q��d�p�@��y��LQ\`�LP�[f�D��ş4���G_���t�|�iG9?`�@ì�|i�j��Y�QxѮ�76�B�' �'1bꧬ?�O��W��t|���wDZ<Xm����g�@m��0�.��� L9\)��Y%e�_m� �c�Ð=�j(���T5�):�A�;����cˈ-\H������O`���O��D�<�����'���d�[;_�.Hx��,42a0�'0��ǐ V>�/�B06E'ޘ'�듡��_l*|o֟��9T�l���bM0|��Rr�RZ�I���	韬�I�|�$�@2
�F {Q�>Q�K�1K� 5����H��% h8�0�@��8W�<!N2��<{�G��[�"��fE��E3�U)�����x2���?�C�x�C�f"��i���V��bB�yb�D�|�"1�w�$�ƍ[��� �x�{�^\CDL+� \[���"@@E�A�%��R-\Am�ʟP�II�D%�5x"�I��\�`l�p-�!
ʒyÁA��n���'Ǩ����'1O�3?A��ڛ;k��y�Rز� ��u��̯6���?a�Dƞk�0y��
)=,
�:��8}�8}�Iܟ@��̟X�r��\��0|	A�*�2}P-�W̓�?	�͘����ۙ���A� 3b���I��HOT
Z��	�@�D�2��w����m��џ��	��3�������柰���ߕsvM���ˡ&��:���	��"T�H%j�Ƌ(,��
ք@~
��|�q�>�Q��z����C�~n!�3�Ϥq�e��'�)]�6��/Rx�큔�����ʧ,�Hu�7�~���e������)R�ۢ]�R�6n�3��^�R��)�3��և'��#�;�*�8dB�4u�!�$�+Y��ȰT��b[�q��C��_n�I�HO�I:�$K�8u�2������=@G���r��%Q�ka�'���'g�p�u���$�'9yL��ǭ��q3�,�A �4UN9�A_�|��U)4��-h�A�Ø3��O|u��l����
fc�%#l�]��ϡ#���P�+�:zC�3�U�q�6�&���t���P ���cX<,E6����jB�,pA�'`������I�X�D�͌PWִ��i��0�!�W(l8 �zg�X&6��(g�E>nP1OhoZK�Ic@ؘ޴�?a�57J�B �Uͨ����֒$atU8��?���ƌ�?����4���?�M>Q�J��B�­q�J��
ư� D
P~8��st@=��
"�}���X+0��QS�@���'98K��+k�'��[�1蜽�t�OIH$S�'���M'X�$h�4B�?{j���'�6-B�8�͹B�+~0��k%�C
J	 �Oz�!1 ʦi����ܔO���i��'M�ٓ� %!@r}) f����?I�(�`�!�J�	jd�!��i�2d􍀲\?�O|ڕ;g��A��{g��G^�<�M�34H@%?�b�x5/A�DǶ��%n���`? ��'�������4N�f�:�C�#1�p�O�ݨ5�'YH�O�\)۷��M!�@�J�9&p����"Oj��AY#W-�x�*]�|y���'5�"=y�����Lq�'Lo��)J�0I�&�'�"�'���7�G�B�'����y��K2������G�\}p���R�<�v��7 ���rGo1��U ��)=�DVgO�G�V3����MH�LZ��q���2F������ ;��蹗�^<駸M3���޼�0���9r�Ϙ�:>&4j�Q�i2�'9.4J�S�g�lx��@`D��[Ȭ�g�ۂh�B�)� � ����2��ݱ���*���j��t@��4��c��c�Օ}���$-S�2�: �FV�+���� N�OJ���OD�$�պ���?��O�h�c�)\�YfxT�z��xP#�q�����4K3�P%)�%Bџ�rwH�2zَ��G'�2{��dI���:�Tä��,VA��O�RR �oZS���M&�I�M��`"��w�p	cN�z6,�*M�O��m���M�B�+�ӱ8A��W���mx0����B�	�
)���*�d�ɣQ��0�jb�4�޴�?+OR��uk��Q�I��쯘OE P�t��*��鳠�Âd�R�'�`��'�;���ǩ(�"�"FΙt�����*T�����(�=+(��@W���?Ye�P;&�.@���4Y����
 m�h�l�
v�7+R�`pڴ-ސ���VN�n��A�	��M;пi��F�nJQ��ǰy��s���	�D�?E�����z�Y���Jb�S�o��xRds� �KI�D����Ea$f
�e!�OZ�D48��оi���'2��)LA$(�i!0�ݯ*���gձQ7�4�����|���,�4*��x%qW��3I4�y��V?1�Oq���թW�&�_����FK��ڄM��:�Hυ5l��ۄ3������\�S�k>�"p��,9��wO&W�)��!}ro��?ɒ�|���*ߨ!��`Fŗ 0���v���yb���`�P K�B0�b`�ůG�0<Ir�I2X���x����	�ޮ)��4�?9���?M��|N�uh��?���?ͻBRh҅�ķ5*�i��! ��-�C"�gԔ�3���>+찁)�*��OY�'�Rp�� W���b����)��I$<��q�mG�f:ly2��w���K?�mZ�b�8睆\�L
���5A|FY���ƒ^�2��M>���ӟ�>�O�q�Aآ�.�gぼ:M�T`"O����锻 �bb�׿jT@("��Ȼ��4�x�O���s��=�R�2I��zM �W�Qj�.����O���O<�d�ǺS���?�O2L�kFʛc�,-1�醬x���p��9F��E�R�)�H�u��g�џH�dү�8Pc��ϧ0[��EGj �j@4?��k�V060t,m��eN��ŀ7�I2�� ��E�o&J�Q#�Ǵs$����+�OֱnZ�M�����OT⟜���%@��E/_�Q
���2#�!�dƭ �\uhւR�0QP<!��n1O�n��Ė'i���-v�(���O�[eƝ�w�]�f��� =+Gd�O��$Έ9d��D�O��S@�*����D$;¾�b�%e
��Á�E/E^��2�*�9�p�Q�eҧ��O���U�a�fקC���`#EA�*$�1�E��-(�� �el "7��d	n��	��"��n�r�|2M��\x �d˚���Ct�V��yB������Ȋ�CO���t�0�Oޣ=ͧU�!�>F��*cJ�f�I���f�'L�0��q�6���O��'~�$��@� YsI�4|��1,E�z]&�R���?��%
+Î�ڴcF�w���p�o��>w��1���?��	�/��q�f+�+^U����̎A\�t�r@���Ճ.��J���(y��&�
 K��'�u:F�DC���{&"JLoZ(�O�����'�ڒO��B��j��T��+N|���"O
= �	X�N�r����7qlU��'?�#=IA;֐�B�!Ѷ,ڼ�Ӡ�R'C���'���''f0�W��:}"�'9r�yGO@�\�����u��h��E�n�<t�f�(2�6]�$�č`����T�	I�`�\�'.t��f�m���y��Fl}�Q{�K�Qb�`5,��]�8��FU:ĸOs���0̐�<)fY�'r��jƄE�:�4Y�ߴpb�'�<Y��S�g��+�����W�`ú����E�g��C�	�ir�49$@��n��HҨE\�L�Vޑ���I�I(���dnK�|25��*�G���C�&T�w�0��ן��	����\w�B�'��镀f3@=k��ơf�F�s$&�5j�4�XqO΁
�BN�p�P���9Ѣ-C��	�!�dBN�4r@B'K��������. �� [��NՐ�C���ΤaC�\�ɇ�q�.���Vi�J��*�n����<Qa�i��'cBTxB�jӮ���O ��cT�{!�5(�ֿeU:���Of��N�(v���O��LM �I��Z�u�y��ĀAD��Rg� B���E�SU�lH�� Z�'4޸($�x����+Z�ᒊ)���ɧL�T���hE	Y}�B��V���{�J��?�J>9�iO�V�vI��� +�����^�<Q�nY4J��]1⌛�P�$1�M�W<�U�i��TPb)Q,���	�"3+����|�#̥
%�7��O��|��i�?�U�K0��-c�������͎�?��b}��������g��m� 0Z� G7ߺ!�U+3}�$��O� �b'F�.Y��A��>�0`:ט>	�F����L>�
U��M�^�UK�F���oP��y�f�#���y��������0<���)� �풰�S-c*��H��03�pJᄝ�i�����I�i}�8�#��`��؟��i�e�N��4�V1����8IrQ�<���K�o�Zܘ1B��Y)�v`�|2N<a�+�-�k���^-�ob�(ic2`��M�x=(�/b���}�L<!�Ù4,����㇒0��8ZD \ ;=�� �<�7�Qǟ�>���Ol��4���A���(B�����9�C�	�
SB�A��٧E��=:!)ي���0t����O`剆n��4�����s�hm˥�ѥQ�yk��{(b��I������\w���'��Ў��ժ�E;��]�$l�?�V��U��1y���c�'�dq"%�^�4Iѳ@��S�R5����h�)Ґ�ئ�0>)VH8BH��@���  "�'��t�~�	=�M�g�i��X���	u��s�9�MBc1tu��_�&_ܩ��pul � ��Q�#iʸ��<������'��x"�m���I���9�,��O-Mq�b�u1����П���;}��<��ퟌ�'lB�-��C�P}<p�f�1�|�WA=-���񄖃CH�OD�x��K�0#B\ڪ>�Y ��'�ʌ(��n��'�d��R�2��qĝ9F!�J�'�T���I�Ф�fc�'U) 	�'#�7�!E��HA����Bׁ�!or1O
XP@��ᦑ�I����O���S�'��X�E犏>�*e����;��M���'N�-n_�T>�=?:���H]!~���qŊ�$�΀�O~AH��)��=;���5��<X�H�2��D�/�h�'������^ɧ�O�|Ṱ�5n{�:u$&}B ��'�r��U��v�r�a�o�i,����=Ñ���p��=6*��gGB�*�������M���?Q�P�v��?!���?�Ӽ��az.�gŏ�$B��c�4��'�<�ϓ0�6�yD�)j6
pSQ�(UR� �=�ęsx��B��З4#h:q�S�@���h����C���)�3���J<p�S�=�.�Q�ݢ`�!�dR�f,Z�0C���Pzs,��8Z����HO>Q�FH�d{���Cd��7�rM8DJ',�L��i�ٟ`��ӟ4��4�u��'�2�>�R2�<o[��Y��	!{z�;�e^�"7lx�Gc��6�F�3�1:�G~'��!�Y�A���lm3D�W�[*"!9�'�7|�RsN�>g��%�F�>�<�l�#�
_'sP!Yf�#E�I`�(��� ;��.H	��@M:���
gd�7)p��ȓl��MYgjj- \�(�:WS��<C� ���mZ��I� ��ؠ6�-x/B���nL����ɟ  ��������|��۟�'��kA3ˤ�9P!��z��cG�<O�����X�;��p@�i��gF�Q���(J��x��Q��?��xrj\9D�t�9� �? l�Y��+M�y��B {��0W�+��<�ծ��xr}Ӭ	"��	6��1	w�+5�,̉�"O��Hb��e��Mq�a�8.�J(�B"O���ښ]��Q��с0I���"O�  ���8J�¥Xv��}�B��"O��#Ն ���ȑ�A$D���c"O~(e�݂`9d���i�)�v H�"O���W��|���JCK}���!�DǱ'�44	��{��SA&Tx�!�DXL&FҒE�^�>Xx��B"�!�J�p��C�zE����#�!��V����B��0^Q��m�wz!��W8X�^(h���:'{n��g�ɣg!�$�,�X���G%��CU�ׄF_!�0L*D�#��B�0�!�^�L=��Y	V��P�B@!�$E'b ���0D�t�F�B�d]~0!�d>AK��"l�<�{�C��n!!�O�Re�d�۰��%ya�H�:=!�Ӣ:'���K���c�a�4!�$,Y�L�ZƦĦ9������y)!��!n�i1�	�.�����3�!��E5P�����)F�rUp��UL�!�$Ьt,�� �T&A�F����)e�!�d�>X}R���L�Є���ǋ{�!�� x���FƲ�x�B!���jsaS�"O����-EdP}xѨD$2n^4�&"O�\r���[�ݐ�) _���2"Ox��1�U�K$.y��yJ 5ٱ"O����4fѴd�D/-�HPq�"O`)c�&P������&`,���O��x�=�)ڧi��$���Z�MH2�넀�`�|��5C�Ik��A&�!�72¬�O\�c�B#lOV2���38�\�:���)�(bV�ɛ�MS������4D��p`��C\���c`ԖQ��mHQ�ӪO�V�9�-��|��^2�lJU��Jx�@K#�z�H��&v�,S��>��P��4�)�hɸz���SÀ_��tb$�F=J�)z���4�a�C[���=I��i�t7-8u���"�˕:-��[VjFp$�|����	8L���� �i�i�� ͒�Z�!��C����D��!�a3�@"Q �ɁNED�'�Ш�ԁJ�K���blӈE�0���I�Ţ�!����	'ۦq}&�Iy~F�c�Mh2�H�r�:�a�Ǉ����������p���J͆��L0�,�P�&Q)*�mڥ���'aɧ��B*'���� ̫@���
U���p6�\�M{@0u#�����Y�E�ģ\'Cv�ɩ��4#D�͂��JT}�E>�?�Ɂ���ëM�h��V���8T�ݢr�_�U�<���	567���f�/6@��fȧ ��8�0n�k�F~r�|�>A��;�,�ض�K�a�����Y<[<��s2)W
Cl~�b�� �?Xċ��V6'ql����ل��'#D��
�Xri�ås#�}����ēgF=�o��w#P@ �
[M��a&�@����3p�ݨ-�a�(I�d
�:�.=��˭QR��曲԰<!U��(l�@4�+u@���@��65���"T`� �P�X�J�ay��R N"N��Ф�6��	�4��(�,B�Ɉl�:`�P�ߠgj�����Vj���:$z�0'��#���$�W��ZqS����O�&X2薳�0=Q���(�,	p��$<���%���~��Wbʿ	bs-�d�AD�]�2��,v�d����N�i&�'� ��oC2�m��B�K�Ld3�e �Ʌr��6m 6%aZ�D�e�D�?�V!�`��u��,��J�4���q�eU0B���Ys�ނ+)D D~�w�∘a��7?zR؂�D�#�H��O��ӗ�4GR���I
z��X����R��P3��V�~������E��*� 3���_:�M�� �:g�Bԁ@�A~4��F��f؞<J��&_(ذ��51�������#z�)gT*�q��O��^ Rz�[�X���$ֲSV�A�WmK�uf�I�r��%3���
`��܀!6�k!N�m�֘k")�5w�'��ҥ�^�f�I����AB��ͯ�M��/�|�n���3�D�Pp.�X�H�mP�2Ua�J�@�����9�����F|B�eމ	)ĞS�N���aW�UFp�$�<9q�η=��L��Rbrl��J^����=��X#��������k���nT�-:�=�DFDx�@`i���+o8�ж�ߧ\�����ɑCZ�6-G
#��l �m�4#	BD�����P`2J�D� �>��c�O�f � `�$+c�	CF���@�I� )�F�ke��kz���`�~Y*e���)�I��y���YV�:e�Ѭg|�7�ZghB��2t�T�B������K��1��@i��@������O(��T���j�1��DϦq�� � �R� ��%�ը��.|�	$QZ��&���t�oØ� O:�BG��[�뚩[j�r��]�07H��<�%�,n9שFz���h�j&@�L�����DM߫&)6` ��ԑ[���BM��؟`18T��o�t�k�f˸*�PC������÷fؾI�O�Ts��&+Rt�D&�*g���Sv�@�>��$UNl2���{�Z6��k�t�F"�
'��Q��~Kl!i�jE�4X�Aeȩr�!Kt�Tg��xbA�a'�ڂ$��霐Y씤~kx����	�x�@ e�G*Z�P�鳾i^�0 rFL(��JAc��M�5ϓ#f�n�+�{r��4" , SF�@#�p�����Y FI�	�f����B�%@���#����4(ɪ	�X�9��Պ!�U�L�R(����i7:���D�;�N�9��/tv��V���J�T��E�D�{`�PE�i���s�H���>i�dR¥�s�ֈ �K�q������)Es�N�4H�8�1�i�}� в��8�$�Φ)D�OT�	��M�`�Ol�02čERB�(v�n �"Kڧ"UUs��GQ�'dT�1q�R>ojc�$����Ү�;��tc�,R#�๲�O^�͓�?�i����֦�Z�ua�$B:��DP����jCG!������� i9F\�v��ƱiP� %��r��^�y��D�[5�ࠄ$z�p�a��%��|�Q�!N�8�C��7a�6�Z&�'h��1Sf�!.�ޡsn�G�4r��\?s���'���I�����<E�,W��0u�V]�g�ա2��Q��'p�8P�p�7�B���� ��TZ8�x�o��(%	��'�t=�3�-�y'��7@�@�SW��e�b%�C�߻�HO�<������C�d����Ӻ�wKN(tfPA��G�$
��p�Oa�EatH:� ��B�1'��M��$�{�� >b`��2��#��Վ+pKq�i�L��U� �!$�".��|��u�i�Z���|��H���bG)R�?KJ���Z�Jp��nl(dwoX+�@	Q�|8�� �>%D��W������P��A�'�>���?��R"���'F��(�V1�rf&���Z���>J'�H��)W F�z���)y�p���	�:phGl�fJ��9���,(,�"Ö1Q���f6M���*P��M�3Z$E�&E��)�4W��	�FЮ��%��D��t"��L).�����,�#B�<Q���!@��`'�H;8����wDQ��Ms�����ޕ?y�6-U�G� h��q���>�o��0ZAq���p2���o���3I[8F-Z�p0���//��	4W���~R����0i���6Yv���"�:5y�BU�44s
L�a�.or\���	=�F8i窒�B�\|P7��%<�r��M>Q+O�O��,"�	γ��dkDo6d�W"�8�q8�ϋ&B6F��
�1�d�tB�7l��G�D��pJ���9p�-��b��=���#�S��gɶVs<��+F�u��NE4-.I���Z5^�3�}B�F�Wp�ya��U�е� �V����'���)t�$�^8Q�cZ
DT�&��ΓN������6t�u� ��g*tM�OT�z)Ŏ3���h��R3�fJ�7R�nڼ]m��EbV�:CL�sqɧ��)m�t,HaMx14r���9b��Bע����QG�L���ֹ&�rdѰF� 5p�T��n(�l�irW���O��kv��٦i��@	Q���e��j<�ir�����=�Q������1G��C��K"4��FO��m	�!��8O�%@�����-�� ��@_tM������0dy4�Z�3�~i����M;8lk!��'H��`��`^�d�ʓ^O�e�$'��'W\�0�i�Q�B���O���-OLxx'�y9�<�����HR���A�Bd�b�ˀʋ�]b81�B�X�,eC&�L(��!�S0C�.#<���`JEb«/5�@�jI0=kJc`r�HMz�XțDߺ����!%�L�p�m�}�j�hIOb1�ap��.���<�{��M���a>��q-ݿM���"��|�&�x�M�YW����	&iyLJ�d����ñ!H�?����q�E�::�AJ�W�'�@���kS���.;�	�bN��Y1��>|��"- ,�'�	�@0t!I��38�VM���$!6��'��ܛm�){�$���MiȄI��ܝQ�̒��x��>Q�`4;(6�#^�8I�D�j�bP���O�a2�A��tpN��"&5�h,��&	���V5��)�>���C�<F*�a'�EY��0WJ�y��&���2SBř,����o�;���"��^�I���Z�����m����>!�M
n���2Q�D����Z�\�� G�(ip*$�5�H�)�<P��<m#����l�$�y���.@�]R�+ZN�nxɓ���'�~Y���>-�J#>�`�1j`��f��>�L���I�tc�Or�q$͸YF��C7Ȋ�0��1$��<��:I(�:q�t0�)eH�eF�L����S��T��"~%�`�ĸ>����4Xجk� �(n�����:�
	H��ݚf������O��?ɷ#�~ZA-��|��t�uO�hق����T�(Q�Y#�ѿi��"?���Ѷ[��q����D�0�D��Ц5؊�$�z��GvP ��O*$���ڸPHi�`A:5I	7�R"H����Ei�i: -�ȼ[�nʞ���Yg���2݊����<�L�d��ѕ+1O\�6���٢l<��1&�t�J(W�"�I�RJ��o��Qpl����J��Ov���I֥>�l�C6&M t��	q'aG�N�ȸЯ��1Hƥ�&����źv|��KM-y�e!�f�W�\��d�W�A8�Ր�A6R�VG|�a��qaV'���D� ��]i�M+?w�
,�p����6t���t[�%�9FH����-V<*Ĕ���FG��hO�q�`6O�e�����C�6^�,j���'	�ѺbmW�]>�i�M=O�%JC㚕=v@�;[�:���� �@�� ����$	Γi9@�4;O���ʴD�@�gyb�G�S$�|؂!��`�k�j:}e|�Z�}�FO9:�j��iq����Ms�I�O۞Ir�B� ��JaC{z8���G��D��T�4!����s}"H ��Lqq�eҹ\yNP`0B�=
.����7W�&��)O(�ğ>�w��Q��6��r��;l�j�iQ}�6-�/@p���O��򨀐)9�}���|Fy�m�M2�H��	֭p��&���XFO�8PE��9�n�Y��P� �Fغק���D�u�̀>Kę�օ�5���B �'��-c
J7���Q�w�Y���Q���B��	�O�t払]@���d��!��O�Woݍ�"��8�U�M� L����R���Y�m�]�����}�LG3�1#�'�J���n]�=O���~�Ȱ�K1 �Lqy%
/R�������M+��	�M�ƃ�R?��5���|�I,Y���}�R)ˁAԔOٰBTl�֦���K
%�0��N<���}̓�X� ��M/@Oʄ;����(�e����)�M��Y�0'���/,O��"���$p <R悲U~�T�G�䒒��U�C�i�����c���3o[V;���ѭ�%Q�R�j���@�����΂�2�n��Zc��<2s�^�)��Y�
��JE��6��sG����'�Ey��ʜ�ħ�<U(6�?�	���.?f$%{�����K�c��O�lт�}A���Ϝ�$�б�'�>��.V�*��H�1؃G�L��c�ʼkbԩք�ZC�<z�4U��]���I�i�<g���C˨d��ۄ�HYZ��u�1l���H�e��H܀��O1����S�? 	r�rd�HFE*�&�{�J��`'�a"C.@�$Ԅ���c�[X��r�k�
I��iԩR�T��$+��MS#��&�?锢�� d$�;��)�:�T&��?�x��獹G8�"ӓ6��q���̣ckLW1OUȍ�ǈZ�1,�a�h��bJ���P�̘>��'E�M٫����[h�O+xC�[1An
(�wj�#��s�}B�#>f���EY,E�+�l߉��	}X�a��)b9.����)5�8Ӈ�ϡ�M;A�im�|`cB]�q��'�a��8=�vjV�M�	�N�i��;v~����O��֧�O��P���z ���A�D��s"S�n�C��K1H�Vl�t�Ǐ�H(�m�[�@H<��G��Ey��$I�������,�`�L7�y�5)���Xq���"zE!Ћ3�yb��b����2w���ʆ,��y"�����%
97D\l�U��yr��E���hF�"14�܈UM��yr�Z�:3����`�M�l�-^�ybB��=�2�k�J_8�!b�U��y�A (��c͂/�~lY�"��y�f��j����(�"%FUF����y�Ҿnz�]�HK�U�Mc���y�׬w�v%&�ߔ ��k��ycՊ-3Q�KRz6��/-�yBo�"�K��Sg��i���yR��\;����E+WH��;$����y�������ۧ咬#o2���B�0�yB �$�Ԣ�5�hUsJV'�y��݇	�v��R�M�J5�r �;�y��α)O�PÔ�M�|M�1�R���y�cV
Y�P�#��!e�A�q-F��y�eA�'���'L��M��%K��yA�Z�(!c@�˹���ڥ�қ�y��UWy#�Ϝ����(�7�y!ѽF�|=B�D�?���f�'�y2(��"�tYk%+U�/5�u5�y�j!l��J@�Y�j�����F��y��"6���(gɴ|���R��y���4I�pѰ���X�$U�A���y��ɳp7��Q�	5@X�BX8�y�#�{1�u;e�܏{ْ`��bC$�y�N^�Jx�R6
�JA���'�y�^�w��@!Ǭ�)4��k���y��,+���ƈVL����
�y�����Q�`
�z������yr.^�	+��@F��u�r�z2���y2�đP���g�΁rAh���隝�y�NA r��� ry��Lp�j���yR�¢)���RU(�0y��
�yR��?1B,�v�>|J���"N,�yB���w���:���<�vŋT)�y��C:2HD�1�̯��x����y҅E�^�
1�v�C�
���ӏ��yApd���ꦸ�˖;�y���J����2%G��L�d�θ�y���*ﬠ������2�d����y�ϒh�5��lN9Ψ�ȓ�H�y��T��9z��'b9����y"S�5V,������m�A˛�y¯I��A�$�0r� IJ3����ybbE� �`ApH�a�Hc!)�yR�ʈ~�pLҥ#�	Z��=y����y�$Ũ�����,��C�02��ў�y�G��$3l�H7#J$"�2�D]��yX�g9�(�tሰ�,���]��yB��w�DP*9m,��A���y�oG )p�����4)��-ܢ�y
� �<���ےk^���2 O`�D���"O2,a�n��F�"/��Q��b�"O&�����v�(�f���Up�"O|���,U2W�V���'�*�x5�C"O4ٳ���1�@$Y7��^8��"O�a"����4�#ԥ��6��=Hp"O��g"GS�Xq2%B��:�Ұ"�"O�AS5G��;V�9:����1"O`١m�U� E�# ��@T�""OB��A��=U��8�!<8|���"Op3p#B&3�> *�)X�0�a5"O&��-ږ�p�c.��)
�"O�u�F�\�1m�p�bź*S|rE"O�d�� *��P���1oN~MI�"O�y�FP<������i>v��D"O�$5� T�Dx��݀t<r�"O6ɠ� ��gt�z�τy.�}�F"O��K%���_Ͷ���ķH(T1Q�"O�0q0��vH��)�'\6�)�"O��(��]A�����D����"O0q&�ٺ�dL+%B���b@3�"O�MY��ȶ~/���&��&[�r�Z"O�\3�e=���۔iؙ }f��t"O�pQ��՚t,~��h�j�!�"Oy� �LI�!Bç�S,\Qu�'X�R�-@ZT�D�+���?[_f���'��"��.$\�9B���Y������$;�!��l˘r�F��rb�Aю�ȓ#�BdY��R"8��l	6mQ=�zt�ȓ7D��@��:x�(����&�|��F>D�B��vb:����üR`>��ȓ_����--� �j��igd��IG~R����T���΂un� �]��y�뚪x6�a�`�t9P��P��HOj�=�O!���a-	�yy�I(g�!SaPm+�'t��z��B2R��a�� �DՄ�'�,��3�		n�	�uʀ�h�.Ŋ�'9��%��1t�̄�uϙ4]�6A�'j��ƭՠ~�ѣ����h��'��1I�I<Qʘ���7�L���'
H z�'��{��1�JӮb20��'�Nh
gEJ�y5�!X����'�&�Y#m�vs���e��>��d�
�'Irh�G ��= ��' &t�
�'��y��@O�o�ؽ�pI��yt��'����� 0�:0I0+�#.��0��'ג��u��C�F5���ė i�1I�'��)�̍lm�J�jN>���J>	���)Y�+g���pN8��1��5F�	Gx�t�c�ٚ{�|�	��6�� T%9D���(y���
]����6D�x�2�V)o��� |��ٚ�I�}��W�V%h�&Rut$�`v��GW -�ȓ�p��`�*4mz�*'�Y�Z�`�ȓ~��䫅䛬$�L=*6�NV3�(��}���XRLX���`@Ti��P}��/ntk��ߴ}Ql���
�(�tU͓��'*�?q�t���4�2�O�?����=D�����W�B$cb��1.�K�N7D�hQ,L�|�.�rf �K�D"0�4D�<:��Y!-̠Lcp��P^h	c�4�Dr����xT���������W7C"C�	U��a�煚)~�^����S0\�JC�I ~��<b`
6~�pY�eCR�kitC�)� TI��q� h�� �ptm�#"O���,�_m��if
R4D	ve(�"O���Ms��� �*n��d�"O�X�0�΋fv(�K���d���
"O Yв I�Y�e*q����`�"O�4��o߿��EkЎ �z	!�"O
����������o�U�2���Y��G{��)�ù9�M�`�Q�v)P7$�!�DO!Y�Hey�!T<hkG(��qj��4�戟8[S��|�\h�q�L�TppL��"Or�24��&<�%�G��d���;O��x����w,Y�%,*�#e#-*ʐH �� D���IB7zx�͡��Fb��XsO!?I`�*�O����`��lH�@&b��,�u�'=��D�4bP κ����`D�����Z�hS�Ά>��r����^�L��ȓBEtu3��ƫ|��Q�\t4F|��S5��İD�ڸ%�~]��"�TO��=�~��j��0�(N��r�Z^�<QV�T�ݲ1s5�Y�?�p�r��<�5
q�>-j�M]�v���9��}}�)ҧ1�M$���K|`@5�D$&��Մ�'�����ch��*���b�>8���Ol�\J6�m���M�
@ިB��#D��Cq��it�99 ��&���cF�!D� �&φ:W2L0�͍�;�(��U�=D�<�%Gѩ����̜O����G'D��2 Q�o��]�%��_��CT�/�L���O�00Ó
��C��h�N�z���������5H���`�@I�0x��ӮĈ+m!�F�"$��ap Rw'(0��كgP!�DOQ�8�V�C		$�љgcҊ;�!�_�l)d�ɔ�v�8�{�O��a{���N��X��5�J.�*X���ٱO��D��Q��h�k�p��RLƵ]�!�č�S,T����>����!aW�"��}�<A���F�����uG�tCt�:}��)��3ql5��ʝZ�X!���	 42�C��^.���O�?8�h}��h�%~C�I%|�z��M�&�8����i=PUZ��-�S��?��n�7z�0�c�#^i�}��g�<��$E<�x��C�k7
9���_�<�t	Ҕy��Ʌ��:nvDK�m�Z�<�cM��.U`r�ߗ>4Pؒ`�}�'g�'�O�=���V9��pH�b�6���O�|{��Z�dɬX���#{H�y��*��*�S�'^T�]����0Kε�w�7�\%��Fz���#�!'�ʌO����b�$�!��8v�-xV͐Tļ�b�:E�qOԢ=%?ys����f��|8���?D��y�cY)$��[��A�9V�X�"D���1+�ZR�¨ �x��C�%D��&�H����v�]�d@Ԉ7ci�	�\��Q���J�A& �kbǚl����	`�=+TYx5��+�{!���o�^,��8��e��w�p�B�I�('ح�'��~"�J�F�`�e,S�dt%p� ���y�Ҡ=̆���ŋ�X���q����yr%����&X� xW#O�yb�I-4�Fa�噚H1�s厊��yRK
�*��c��?sQ*}˵�0�y��Q�rÖDڶ��x1���ҧ�yb"I�3
���MDpXn��F'�y���,w<�JDoEל� ����y
� �Uӕ-O�,	�6�JM��1#�j���	D�*���,Orj��� q!��:=������u<x8�4����hO�|�@��	&Tx�'��!\���'���Ey���ܵV<����oZ3|��@I�g�:7m-��r��\B!���A���PCJ�;0)1D�8�G#�o!�`��b�8i�r�h10D�������2�q�tJ7]�n�@�1D�� C\��>��J-x�0��
$D�tj����0��CL�#
���d!D��0cCJ�s\���%�,�T-�>D�,�g��3�V��D�&Y�n�0$?D�\i�ʎ�5��H�v�I�Lۂ�XP�8D���4c�!�&YzGO܄acV	2D�8�'a��
�@����]�t6�"D�,�A#�1wrl��b��m�,�� e D�8��MXzV�帒�58���D?D�H�u�l8����i�CB�u��*;D���Sh�Se������ s�-���3D��e�B9"��@!@b.<Ⱝ@�.D��q�雋|��x[�(�LԤ��*,D�x��� �u��h �wHČvF(D��K��Tlhu�W쒥)���ń;D�� O����Æ-~�l��i:D�Ģ@�I�C�`"MЃ^�v@�DK,D��KPMʉ1"�i �?���->D�dٗ̩MhbѺ�#H ��5�<D�h�!��i�R��v��'Þt�4�:D���C��K4�����]�P�*��8D�`AB$��ʎ���P9~�W�6D�p�g/�+}x�9���K���� �5D�XX���!�<���������'D�d�&(W"pq�H�������a��:D� ���Nw`��F�@6]@�L+D�pQ��N,R��1�@�GE��8A$%D�\���C�4�NQ��Z:�lӑ�#D�ܣ��Wi�,
1�Y�9�l4r�;D���t�P]0i�q�K�v�~�.4D��ə�UXD��(��E�\hi��2D��[EI	93��(
��m.�IP�0D�8H�GT�[����p�
.c?��h��)D�({��{~8����1wn�Za�:D�dK��'��l)U�wqU 8D���l�>�}9�n�5M�ɶ�6D�pC��Z0Q�X��d�Y<q�f����5D����)P��=X��قBCZ����3D�l�U�
w�&���)܌x�f�0D���so��^T�H6c����H�,D�8 7J��?Ѐ a��5 U�y���)D�0(�"HA�D"�P�.@��3D��q&D��*$:d
/*�S �.D��:�d�a��pA���t��ڗ�.D���C+_�z]���Ǒ��Y�R�8D� jr��Yx:CwD�?a}���3�7D�P!gBߟb�P���	 KCd9gk9D�P�����q��kڣK�@���%D� !FQ�| ��dU�Ui{!�$D���&��N@&��r'A1#��p�'D�p{�m�5=^š7��t�x�8�	%D��K4��?�q!G��+yYB�qs�#D�lH�%:G�,ϛ�rZѳ)!D��O���b$Y�X;T��CE>D��ɵ�S�B�|4b�cB�p�:�i��8D�@�v��=��|[�	�_i.�Ň,D�� ��;ƀ�%pr��`͓.����"Of�Q(�,~
�����L��#"O�P���-:fi��D�}-Z��&"O���PEDj��v��B*��� "Ot���!KI���J�Դ:�1��"Ou��	/Q�(6.�8+H��"Oh��Q#Sg�8�Y�"	�o#<�R�"O4ls�n��g��t�u *�<� �"O�� ����4�ʯ��i9C"O��h��H�6���'˼����r"O �à�91��Q3���Wg@0rV"O*!��"X�>�2�%����,´"O�ܺB$
#,����#�cEh�x"O�]�2 ��=����,ߕp��"O(1 �X�H;�ϐ[;����"O��"GÙ3`H�� 
�0 �y�"O�eA3�ݖ~J����$)ϴ�"O~,�$�Iǚ��A��\�"�a"O��H���RM�%�$��;@��99p"Oj=Jg�}j*����N����"O�%�%�سd� �$΅L��L)C"O0Ѷb߸"�T��M��0�S"O0S�mC}Ҧ��R�y�anY�!��z��t�BkS�Jo�-k`h��`!�D��41:D�3↨GU���6(J*�!�� ���)���O�L+ӧ?�!��\�D^��h�ʂF�i���7�!��!E&P�K�����3k\�[!�DM�A�8���nݶ��-��J�"O��;�*�gz�Q��
)y"E�4"O� S�d )n���#�Nh(D#"O�qT���b!�%�^3\H�"O̭ʆ �>A0ƇN0��k�"O��r��$7�ցZr�	@#���"O�7͛w�f�3v��pALA�,3D�$���$@��T�@(C�<���+D�0j�lR��.��s��D:h��&D���EX�.	�g��&o�Bi��	#D�X������]93��	Pu��C?D��"W�W�S;�A���	5�}�P�;D���.��JhR���?O|I�3$D�� ���R�j����F�ر( D��QRU_��J�j�XDn���L=D�4��(3VvAHs*C<*���(��'D�����\!�(p�oD)��i3� D��Q�)�dJ�*0Dչ*r�p9p.=D�$�ဩ%V�˦N��t���6D�|q�'�&_�T�7[�����4D�xzVN�7�fu
5�ՑH����B�0D�xHAo�&ʆ��`��z�<��3d*D�����"/.(���Z�P�[4>D���1d֋@d ���WI�^xᡩ>D��C"N!��ж��hS�s6�<D���A�0\�)!KY/$<{�n5D�l1��j��!�`�L����9q
4D�H�
7T�Th��̙{A4�вO2D� �wC �yR���8
���m.D���d܄=dȵ�D�W��q��+D��ȇ�� �Xj�&�.���!��$D��4��J�����j�����4�!D�˳�P�bb��U��.�|�*1@3D��ؓ��=*�á�?/���D�;D�Ԣ`�Im�@@HLؕ`�C6D������O�a�s+��}���2D�� �@�&U�p�%٠R�
���v"O�����V0�Ȣe�
�V�L�"O��S+�l	���F;Y`�@��"O�ۢ�����d���V&6-B�S"OV����.ns �w
��j pܰ�"O�;�� ��akW�^! 6��Җ"O0���:��dS2FY�d�S�"ONx�A/J�:�~�A�∉_6h$"O�Ut)�U����Y�(0�"O����h̲6  3�a��"@Ҭ�t"O�!��H	.�Tg�%׺XӴ"O�%X�KO�Q+�<���˺'@�"O�a�'+�KXHX1A�M1���"O`SCۢ:�&���E��Z
q"O����)ѝ$�ܠ*'K��wtȈB�"O6�PS��@[�XC",9`�I4`�!��˹S:�Ha��R�c�T�3�!�d���
i ��N�Ʃ�'��2�!�Dҧ@V��*B}z y�Ã\�I!�db[��1��БFmv��2��;R7!��Z�l��0iQ�pE�%����-:!���>1 ��a"	�=�I�0Xx!��2i@}���;!�<y�E�``!򄚡36XQfկ.�2`���nY!��0N^fq�% "F�@�j`m�T!�$��i���$�Ջ0n,��̉�Q!�$�5]Z�R� �0]�
1��5A@!��'�$��H�i���w@ӲR!�د,Ɖ�P)P?W��41���#s!�D�wTF(�R(%W�=��n_�ld!�D���m�K 
������� 6!��B"``�	�6�R���UP��ߵq!��
 ��\���D��,x���P�)!�DH�V[�d��+�8~5Up��D�!�D4��q�O�:'�p5˒�Tz!��R�h^E#R A��u�C��2�!��K�=����N\c�
Bf!�ĉ�<ݺ��P�ذ6��-`!�׷(�첰c�	J��Q"F�K7`!��;U\���IH�5�`���a�b�!�D�".m�M+A��HqĠ�AG�j�!��\�5?�3#��'Tz��LU�a!򄈢�r��[��t%��eQ!�$�8"T��B�&F�>p)tF�6;!��+P�ԉ҈Ƭk9MC�*��v2!�$��Vb9Rb�+ �c�ǉ�|!�σb�$�թ��,���f�ר"!�-h��,R
�Z������!�Y T1�̹1���5����FbT�s�!�غ~F�(� �jG愫ѣ��!�D�,Vf
ѻd�����H�9n�!�d@�Bǎ��U-@��̞c�!�Ҩm�l���"�U7�T��T*�!�D_�������F�X]�nʟ\�!�DHQ�Ι���(b�*�+�l�%J]!�$�@d.BF�P�U�@L#fl��!�P�:Y�x�$���~7ʁ�ᡔ.:�!�D��
�phf�/*����!��Ƶd���	���.*,L�F�U6�!���7�]���A%`��B f�:O�!�d k=�x! j��	j��O�6�!�D�� .
h�.�	pU꠨G���9*!��:Bz ��@���c=�Ei3jF5!򤜟|$c��Q$i�*=�2�đ !�� L03��
����D�]�b�>��"O�j�$N��� ��x�n�I�"O��=�}k�I�k����E"O<����Y-a�A�2n�Ap�̊�"O�Sw
�)E����۽UÆ\�"O���0M�>nJQ�ǟ}�bEp�"O�s5��- e�֎�)�����"OZ�S�j� ���@�n��s��8��"O���q�[(8䜌��❔����"O��P��(j��[� U?u��y&"OA���!�: h/J"6lH	�B"O
�Cq��`��1L��lBġ�"Od���G�Im���ƈ�y�ʨ�"O.d�0�Z��Ԁ�`�M�l<)�"O�	�ѡſR*�y��Ão`�"O�@��`U ��Q��̂(����"O���e�O7~O��qc]*�Ac"OB�r"�ٿH>:���^,Y���
�"O��"bz�T��
~��<�Q"O�%
�L��N�t�Xc\
zɶ
�"O��e��;�B9qa��4���,�y�KI#�0Q��>kh��ٍ�y"�xS��qG�+Ři�p��8�!�Ȳx@��3�/�j��2NK5�!���&b���" dP���zG���X�!�d�}����qL��]�fu�"�Ca!��
�xi6��2BL�p�x1��F��yD!�7%!Bᱲȅ�&�8�;5�(;!�е9H)���H8w�����)�:O3!�$S�ewHe1)�%=l��cH�:!��=��Բ����SXH���	2E
!�$�<ΐ�bs��IL@A�Cu�!���]���� �.Pq��1X!�$
Z; �96-�.,|��c�73!�R�eϐ<"�ëg�4l�*!��Œ"r��D+H*! �����ɓet!� -�l[��O;
�Ғ+�\!��!���;g���S��d�S�S!�P�Z�J�Y�Q�7Vк�*Ì"/!�DQ��|kePvu�U��L!��0H��8
�����p��(
!�ČL�h�Q��TRH�j�&p!�QyNlK���Td8P7
X4C#!�C��0)�슪r>��e) {!��M�uiH�PB�Ҏ.Ƙ4�t $:!�$H��"I{fBF�$
.(�W��+y�!�dLY�u�n�7�̔�e�hZ!�d_�d��maă
 �Tě����!��(������th ga�17�!�0z~���c�T�)�����9K!�d֭c��;D�F���MC�T!���-��q�
v����L!�!�L�<?�2��ԭD�-yR��=a�!�$� V���c3��<��Z��V=_!�$���҃�I�s�J�02*W�	�!��3�=�A/��-H
��HL>X!���h1��bd̅��%G�~!�۶l�% gO�/:.N�椗^!�D_P>��r��O~��26��:�!�5}���@�ϵ8�����W��!�dM�W9�$ß8�EҢ���!�$��c� ��T><�~�X�,\�!��8���Ub&m�hAE!�+L!��d��<��K�2u����.G4;!�� �\�ꅆ}��]�#!�mt��"O�1��S�(���:"AD2BH�St"O�1p�
J?XkbX�'@��}�"5�4"O��jd��,�
 ���Ua�=��"Oε�B��\E$t(�NY�q%�pj�"O�����3�>�Ra��o,��It"O ��-O n�1�j�&
?���"O(��ujAJ]��Ѯ>�"O��"f֜4\sbH�G3�h��"O�����6�Pl�h�	F1�9F"O&M��C�\@�	��1��0"Om�� ��� ��"�8�ld+�"O�����,�0� ��s�p�8"O*�YWM �X���
A���i�<�!"OV�!G�.O)��ÂW8t�:W"OF�3`	җu�0iz�c��o��a�"Ob����#;Ix�"�ݯc$֘Y%"O2x7�N�	�\���#z49�"O�e��+џ6g��c6,}[̌�"Ot�XR�J��
��j�%V��i�"O�"�
ѼvfF�*;*P>��"O�x�q�	�=ؚE�1��	<�+�"O���A��i�����l2Ƈ
4�y�
�^���5I��*3��A����y2΋�.���2�_$%�Hae"Q%�y�
L0~��a %Pr�) �²�y�K�-	�D�3a�*.��`@�۫�y��O�( �p�1�����F�y��=vp&В���,,�p��Kˋ�y�1g	��XqNJ-'��G@��y�ރ)V�0���/9,�:5fV0�y�MD4| ��d�C� zJظ�h��y�-�I ��R�˦'f��ڄ��y�(ǵ{a �J���:k�������y�$�3C�:@SE�>a� �S�L�yrI($\}�%U�R[��̕��y)��VȽ	s`K�3T4�#�*�yR�%le�F.&?x�R��«�y�&��0*X� )Wq��� 	��yj��h�}#��82y�Ma�� �yBd��fl{pB��-���1��G1�y�C˺��WH��p`��k�/К�Py2%�=(���z�D74�x����y�<�"A!�6�zGĵ'��a��L�<�V�e�`jd��8/C~�^d��&n�X��C��-�L!i���n� �����@�ۿo���lT�ԇ�i�X���	s�v-a��!B��ȓDhx �Q�~8�㥋�x#���T<9R� ���.G8�RF�U�<Q"�ֈE1:ـ���1gV���g��l�<A�n�b+ΰ���"��,)�*�l�<�� �3k�D<���Fr��(oe�<���
 ��`q���,�@�W�]�<y$�	�G��LJ�
�2J+ `^�<�O���Л'K���i�Clf�<I3`��j���E20���:���e�<Y�'԰p� �T�\�i*�"b&�e�<aD�4LT��6�	:{�ڝ�0�l�<1�*9/�x���4{��貍Se�<qp ��j"X5´�Ǖw����-e�<�@B�O9z1��-�y�+_d�<Q�(E�p���#�&<������MW�<y#�=0V�QG��!��p���IV�<� y5
�xrv��1�Z�h]z"O�����7zJtb&�D�R�~�"ON(�T�]�7иCՇ85����"Ox ��Ľ7����Aǜ0F0��W"O�=A�Ɗ~�X	 �%�:@�8F*O�T`���Q�N��#�8̂Y�
�'ڔiG��K@��K!ϯc:i�
�'��SŖ~�b�x����c�z9�'��*!��	S�<A 2UO���'{(�S��չw�d�P�I#.�8�'��:��(a,%� ��I����'��X� �Cq�����H�oÐ��
�'\�ي�/�X':aL�m>�i��'P�Gn�.C�T\K�aé6�%8�'�^|�U�WK�`�YѪǵ&�����'>�U%��ba�J��N	H���'�2mK���#W`F�P�� P���'Xj5q�:Y���ÀZ�qM҄P�'8�a���ʃP�<��E�y��:�'�Μ{� �/��8�@C�w:��'���p�eO,o�Tj#Î�q�<�'w����m�T�"bb��1
�'�ř��\+J��X�AN A>Q�'���c��E�45���r�"�;�'�>5��f��P�>��,÷j*"�"�'7�Pr�g�;,Ϛ� �f�����'���2���?E.��,WV1Lؠ�'�\aE��f��)eL
<B��H�'?�!��E^�qdBH��1�'N@M��E��!�4LO���b	�'�R�	$��c&ذv�Үa�����'*M s!�$�]�T��3]�xݒ�'B����}��� J.|X�<D�P3�K�5��1�P�Y�i�����$D�PPMG?Q��
�6D�r`"D�,�GA:W&4i���[�+�.�� D�X�D%�����Z���! D�03�՝#GJ��s�R q���p��#D�S�Y6<$����b��LIE�6D���d$7��ē1�J�δj�5D���d �+J��!F1Zc�ѩGG1D���BC�.oLءqiB0�D�0�/D�4h�H��"����+�6���a�:D��ՀI=�޼Z�a �AI�1�$B2D�����`�jUpv���I�C;D�<�֟t�v��v�bO�i��3D���#�M�.e��-ff�u�R�2D�L����$`���w�ټ
fXi.D�|#a-2�i���'y�P�;� +D�r3��\�染M.0�۱�)D��uV^��1z�ˈ5Mp�P��3D�D��.h�1��:P#�����/D��÷�W�6
d��RJP���*D���휵rK� +�m��S4���'D�tA��#	^h<�W핈4R8l@��;D��FɆ ꢙ�$+I�b]ބ�C&D��*�.ʄ=,�GG�)o�@Z�$D���#C�G<��0���Bl@�`��!D��:���65n�y�O�+e@����9D�����t�B��KB w<�!1��;D�h�`���lhã�*B��m�D�6D�Dy��L@��)�`c�'�Xxc!.9D���5W7:�2�04�ϟJ�$:5 "D���g�܀>�\�UIϮc��8�S�2D�� 81@#�o��q�#FaL�tj�"O>����NDP��T [*p��a��"O�y�f �����_(E�@�"O�0A�`�26��2R�oY7"O�,��#��M9�G�)_:�2C�8D����G{2�Uc���1�<Az*D��cl�*)x�����z�B�&,D��8��)h��3��I��G�*D�ī��P<%�@$��@Sx�� �$'D���	y�4�a�c������%D�(�c*�B��`g	U�Ps֙���$D��@U)�/�ƭaB�M�p�0F�"D�t�O��*�}�n�4�t��E&D� +u=_d� 錑r���j��&D�c��O'X4=��iλ֘��h$D�H�%Ǒ�`�j�K2��s�#D��#�*ŝE P��O$e�4;�=D����e
#e��K�%K:X���'D��8���7O8M���S���$D��X�B�2Ek�T�1�F�8���Sd"D�h��-B�zܼp�2)�X��d(R;D�(�HB�L�d�1�aY
�+��8D� ���~�Q�uHJ�J�H�c�7D����n�x��hQ�&V� Fi+D����.L8Oc$ĺ�dB*=Q��z�#&D�|C����Ҍ܌ O��˗�&D��p���l#�@�%`[�=��D��j)D��)q؄de�5	P`T�4�j�`�&<T�H��쁝:Ɛ����3G���u"O�D��4�
��"G}=(}��"O*5h�C7 2Jp$K���tX!�$��і��t(ڼa����$ЍpB!��1R�P�
���ᲀ"��RH!��4;/���&�H	�J�	��E�4-!�D�nH���Ƙ[�^�c5�ć"!�^�S�82v�b-5A�l�m!�W�u}z��`���8@xjq�E�9�!�$M;�BMj�]�*n � �X�j>!���|���0陊B��Y5dޡ;!�D�>M(r��.�->E���!��W3!�DV8���@V��J$L�(!�DH�U{&"�j@�	lXiR���&R!�DD+A[� p����d0i��ؤL�!�$�X�,	*#�G�Ҁ P/�!�$�&eA(ɹ���6{�M1�MZ4c R�)� 
��Q�D(�Q��_ڔkt�<D�������f��4�ʛ{I� 8��0D����*νz�LuSVe�^j6�zF/-D��{BM�-u�С��Ą0&�E�ҁ+D���PH@�/�J���EX lDa�u�&D� S�F��~߮�7Eđ-�:Y{$D��a��!pm��宖�w8�7�'D�0Y@)��z:V1��#S�f�21�r`$D��S"2V��!�2G5)��;1C7D��S�@�Nf����P.3C�(�DC5D��s'��!��DIm��8�o5D��X$��;U�&-�2I�5
D� 26�6D���,�Y��u���t����M4D�ܻ�'�}>*2�!��ti�m*�H1D��c��_�!gX�[�o�(���+�4D��2�A[V7VQ�0�a~���2D�$���B	�8�wB�#M��r�a1D���J��HF��4Dٰ?��N5D��:�o/����&W��̒׍7D�� z�A��~A�YU�ϬX�Aj�"O
a��D�	�2�+�)Ы�:t�4"O��6�9�N�k�O»0{�b2"O�-Ӕ��a�}3vM>̼�*g"Ovx��K�d|:�AB�0���"O�pB� 5�5�q��u�f��%"O��Y�	�4a�,���!L�C���1�"O�u�TL�T�ؔ��1��XR"O鈶�G?;HՀ%�P;1��4:2"O�3$@��]d�A�&J���$��"O9�W��;����+�:�> XT"O���
1UQ>iS)�:Y�A"O�m�奟�Cv�=3R�� yJ�"OT��a@��|rZ��'��q���"O�d&b1x�hR(���J�"O,=��#�,`4n� }�0��"O�]oT%$�@$�ګR���a�0D� �$�T.Q5���T}�����<D��P�J#-���+R
9� �W�;D����¹D��* Ɲ�udz4@�:D��A7��Ah�Y!p,�:Md����7D�<!��(�j�[2!�"Ģ" 1D���.Y�b�J8#���2'���x��.D�h��L�}/�sTl��l����*D�80qk��R�ī	���)��$=!��׷����Ř",
���M�&L+!�9���� �ZG B!�/f!�d�8���v	"���fJ�.�!�d��.*�%��	�z|���7V�!�ױF&��D��q܅��k�!��а���Ȟ�s
.aa#�P�@�!�D�ch۱�	qj@�� /�$X�!��*	.�]�3M՟jX�Y�C�2�!��_�� �K`X�`v2�
�"��Ag!���ڼ��'!�$E�C�7P!�F���J��ۖ4\N��U�I!l!��w�<8�f�3p>�C��5d!����N��3��L2�$rŢ��D^!��wc493�FO�~b�A!�R�M!�d���Ԉ^�A���`ˏ�j<��
�'�x����ZW��*Q�]5U�l�	�'�8�¶f�<��(��� ����'���	wn˴i�Ɛ���.uL9��'k�Ac�C��C}n�3�,�S(�Y�'�p�B�&T	N�ҽ؆��y�����'�`
B!��U��S�N�$�� �'���[R��#t��gE�M�6|*�'��!�5f/�t9zDe3W�u	�'�8� ��S�S�ݹK	�*�����'B����2�ܰr���Kڭb�'��M�$_DR aS�I��� �'b�)��L� �R�����0M5d5��'���.	�N� r#E��{�"�8�'�d�[2�V�4!��F$oѺ@ �'3��9Bɔ-A󮬃U�h��4"�'U8p̖7.�x�X�Y�4��''% EΝ�d�\u�%��X��Q�'o���B���3~���\&M�@��'8��ӆ@I�m�]�³=�uZ�',�10W��� �饨���8�@"O*��A/�� �깊u�U=С#t"Op���G�jJ\4h7��q����"O�{5�فS��\` K�h�@<�w"Ov�Ui^1}©����6&<�sA"O� ��8A�^�7O��j�B�45��cW"O�=� #f�Ж��55vx0Jw"O��q$�(i�����/�=�W"O��+w�/kwNQ����y��p�"O�AH�n�(((�X�G uxx#�"O����LZ�dV�4�GǤψd��'�t��'�U��&����D�f�5��'gh�X�ׂ?.��2"�Zph���'GBe�7( pg6`������'�&E@�E�̝G?���	�'̄P�� }�]�$`�9� ���'h��B1I��#]���^ò�"�'Pbh�%��/w��D�!"Q�Hu	�'�dI�M[�l}t� ���KWvb�'Q�u���+w:�@�	3A��I��',��y��Y�V0Ha�̃-ࠤ��'Uv=�qHK�%[��
�W<�"+�'�z���g	M-.�R�g�$KW:���'��X��-�PC��1%�/8м|�
�')-X�gˊ>�V�s���6��){
�'�l��D�O�D{#'�>��hI
�'�����?��])��G�K��4��'ώ:�JN���-P�>��Y��'�>Yi5B��w�T�q �A�i�X�'�>Q�b��8i;�d�5h�\)��']�؃b�9'4����Z��,�'=�Ђ7�B���H�IƕX�=i	�'L� ��{��ų���f��1	�'~�]� k_"O�I���O43Ju��'�R�٣�6")��94�ۆ=/J�'2��S��٨] p4�@�	3��C
�'��ypi4S��#0N��5I.)j
�'�
�aqM̽5����� ��dԆ��
�']�<�9g�*D�Y��"OX��(��8~��#"ږ=!2���"OԜz�Hٻ�Na T!͍f\�@R"O� ��&@�1ʤ 	u��7"OVHbྲ�٘ej̀4����C�G�<Qp�r2����^�t$�KP@L�<���[aw:!(@D�5�&P��d�<)��<���(¨�.:�$�r5�Wx�<iSI��(A"�����;FzDS��Vw�<�d���4c.�B�R�����y�<1�(�'[M�	i��D1e�9	CSx�<��_)`������'#�ְY� FY�<y2�̷2�z�(���ά"��S�<��G�5V1A-�#\~8��H�c�<q�J�&`�4��F�R�Q��	�!�U�<g���Xc�X c,4f�*�8��x�<A�e%6Z���H+I�`�[�+D]�<���P�4�ᘤh��Ȇ�BZ�<��a�6Z'��#OE�8@��KR�<�� <ۨ�9τ�~�B	P!lx�<1Wʂ�DǄ(F�<M�x�% P�<7� _�H��X �fp�G*�O�<	uo۷2lv�VEl�L�&��d�<a��S8>�8p�/A�C>�p�a#b�<QWL�'⦵��ܷo
��m�e�<�1��:a�BϷՐ�*��e�<ᵀ@�-�Jy�V��;P9���d�E�<�oC�"�|�Q��b� �s�	�1�y���bT���M��j��=�Ő�yB��7~���'�۷J�f��I܄�y�&�mF��s�(ƵVy�e[5��(�y
� �$��L�^KV9 �_�ʐZ"O>�� f�tL�Raw��""O����W؊Z��04���a�!�b�<92��<I�E�pn)z6 QF�[�<a������XPj�$��$R'YP�<��0<�Ƽ)�灣�^<	�CP�<� �5��H�d�X_j��0��M�<)��B�E�A���9}L�K#DCH�<9d(�)O8F�0�	�53x|��(Xy�<�s�/���+��\���\�ΐv�<QաWf���X������Ǉ�u�<�Ǝ�x)���7�%B,����p�<��)�*�xۣ�Z5q�\��D�<wg��xQ������.���� �Y�<y�@�D���`��Q"S���*OOS�<AI�a��4�D�Lb�r��C�[L�<�Gޝf�-ӱ�c��"�(F]�<!נ#y���P3�C�a��|�4(O_�<�V:e�M�LZI�2���CU�<�ڸVQ<���dgf��"	�J�<���!+h)[Q��0则aC��H�<��M��6::��R<F���a0,Ap�<٢�^�q# h����5o[�Y�Hl�<1�l	�<�\��@T��J��P�<5��#,�^���Ȯ�p�L�<�2�L�:�
�Fӭ�X�w�H�<a���>=�
&���W V!��(�K�<A���s��JQ�'nz� �fO�<Q�%���M���%^2�;��v�<��"�2(0�	�-%vi����r�<iN�$}6��	,�a��_o�<�� �K���T��m�f MB�<a��_"Q0��
�[|(űG�XS�<��(B$T]T��WÅ))�����	�x�<A! �=�Z��צV� �1Aq�<AWbʬs��@��: ��0W-�i�<��bK$u"�Bqa�;4�����MK�<��KŴ%4�;�l�74�f���M�G�<�昦�F<�6dG�E�DIT@SG�<�4�����ԉe�J�Pm(i�!���+4����Êo�=Z���*	�!���.�N�sV�_��h�F�^��!�6�-�,��D׬��C�d�!�D��_Yr��6-W�!�P	���-�!�d��u�$%*�I��lz��$)E10.!���q�xA�"��`a��b�F }!�ߤ)D@�aeJ>O�D�����$zk!�ХI�RbŁ�4��0	 
�I�!�]�=9h&N��F�V�0wI�y�!�dX �FTa`
N�B�H��S*@�!�Ԋ6����Ś�M��v� p�!�DM{�1u��M�d"�ŀ'N�!�҈j��`�P'5PbT%E!��Um��{C���(z������!�)o`�FM�tr<݀�U�@�!��+O�.����ԗ}T><�4�Xw�!��YwcԤ؆L�i����&�Id!�$B�^���+F��.?��9���R!�D�9Qd�)#u!��1=L���c�`<!�D�btf��ǉ��/3ހط%fQ!��X�!b&��x�aa�+�!���Z�R���O�&l��h��;�!�Ę!F��JƮJ2p�d�){�!򄃋~�JP@�'L �8�A@hn!�� �l;��ȢDNr�cB�W��L�B"O6)�p�ӵ9�x��l^�{<%�"O�����^q��m�9jm��Ip"O2�xC���yb'_�iЌ92"O���<&��
�/ߏD"�	p�"O~P
o]� t�������
`��e"O���wf [� ��M����̡�"O$<�d�5**��b����#"O,�C ˖�v*�uJ�օj�8��@"O����/��]H�(N�B�eH�"O�@�",��H�W莚݄LAr"OHh���w���2)�\�2"O��˓��rȨs`��M'�P�7"O�i�1,�>N�³/W�"p�t��"O|�(a,ϑtT�=1s/�4���@"OZ�pC큨R�P�b�C+A�$(�"O�����a�T��ņ��_���"OX�jF&Ib,���ˊ�k��$[�"O�5ՠP/� a�K
�**)�5"OTt���[�7S�hP�IU)��Rv"O�T8-)\LjD��̵=�d@A�"O
�
�
�$f�3F�c���cr"OE���̙:���! �<�90�"O���EɖC�̅�����;�fq0"O�!sf��;yo��ӱ �6��ճ"O��S��QNX�Q2 Y��@0"O�<�bꊰ8���B�0g�$ܲ�"O���Ǐ&8ή�a�������"O�T���
�qGr�a��×$��x�"O.����881� ��g�����"O�Hw�ӭ}���@f 	 n���"O�@�� ��(B6]J���F�yٗ"Of�A�N�'r��`aBO@I3����"O.t{��.'.��!V��'m87"O&H ì\JB%f.?�$��"Ot��6Lu��Y�,�!F�@��"O$�ȂH�H) ��F��Nb��"Oܺ��\[�n��'A��[A��d"OaA!ꊠJ��03T�y�t"O�%���B�_u����dV�9�"OE oޗT�eX%���>�,4��"O��)ӭĔw�:��;|��4q�"O���e�)+����!�Y�s"O*��˛�*�@�/S�עp@�"O��y���8'���
(şe�,�	�'GεrcD�h�@3pdF2^���k
�'�zM�&���&<��K7	�A���A�'x��#rDɮ+ٞ��f��(dM�u��'��hz�$ʇ4Fɺ��
W��q	�'x$��կ�����W�S��h�'X�X���>C>Ƶ�C�<{%�YP�'��)��_)K���n�~�f���'Pq��	+"�@��剱w#�j�'˄����U�Q=\8R���o�``�'�&#�Φ>L���Ő7r�\��'Պ]rb��8���"ap���']��P5�>|��"��hi"�A
�'��\��E&~�X�f1]=N���'~��Z�ύ V��
E7\O�\��'�H��g��Z4��cd۟U�����'���	V�	:w{��20�¿��uY�'��q[�o�1�|�ȄJ�Ĉ�'~�{�ΫX�nX��aM,{:�� �'��-�E5t�u �.��l�Ԍc	��� `�����	#��\�B��72�|��"O��3 ���@I+&����"O��:�D�c5�8��Q���RW"O�T�H�:>0Ab뜬a_h��&"O^�0@��5-F!{7kG�p�2l��"Ox�`�.J;hBi�6����"O��2/F�`~����	�).�H��"O�i���O"�Q�'v����$"O�=��aF�Q�� �O�Z��P"O2xq��ש}R~�AH��r"���"OH�A�@봉��-��)\����"O���&�<P��m���=��0�R"O��8v����I�a�J���"O�)�c��
��0AS�Xb�ī�"O�5��۲�Hܒ ЂD�9�a"O�1�lɤv^�噧�;,<y��"Op1�����Թ�P`��t(h�"OX��L����V����v5pW"O��;�n+s*t��Q�	�����"O*�YFbރ8��*f��:z�JͰ�"O�4��D�p����ۜB����"O�j"�]^�aa�IA2GP�ٱ"Ove���j�#kI�f28|�"O��L�=>�U��l��A���"O�Mr��/���ʗk]�թ�"O�٥ろ`�����
� {�	�"O�sV艁 N��p��3a�r�"O�Iz�o\<u�ЊC�JU_QIt"O���w��5�&�����YZRD�"O(p��`)���Y�D\�trdt "O^%����)[�FY�r�N�` 
��d"OJ��`B5�M���V�O�8E�q"O�e�uϊ%L�!`c�:+�H ��"O~ݩ��H�����~�jj5"O�D ���gZ�����!#n���"O����k"�I2�� <�A�"O�|c	��uWN�PNM����1"O>)��ԋ.d��-&G:*	k2"O�tR�/�&aA�xq�J�|9�s"O�d#�օ�e ���ucDJ�"O����+��ԃE&I�:M�=�"O����Ɏ�"�0УQnI�x0"� ""O�����X$G~f���C�o#��*6"Oz��M�~�mN&><H�"W"O���� #�����*i�8Y�"O�� �F0\L�ArF`���s"OH "���KvB�+Rc�mL9i�"O��b�� ���rd/��n<*h��"O
y�3�%*�ɫWL@8f+����"O2e�1��i8v���k���l,P�"O�0i4��	h�Hk�mV�k��A"O�-��Ú.?�����+_�B���"O&�R�gK_�Xt��9Ϙ���"O1��!*)�>%Ɔ�>��� "O�x��ac�(�Gќ.��YR"O����~���%��7�����l�y�A�7����1j 0+S�a��?�yRAE�$�zt*rg #,�2$[�g��y���9hK�ǥ˺����B%�y2FΎ�B����M�|)�d��m֩�y��V�X��a���9l��m�cNZ��y�Έ1L&	�GV�xD U�����yR���(E��q��t�0R���y�J�f�f9X�� �,q1BȘ<�y
� b)�W�
�&L3��͛D9���"OZ�
��?L��ؑ�<E|��r"OP5 D%�,|,�[LûoN� "O�hq
�<���:pD�(gĜ<0 "O�QxF�J�
���XPD�&�P�PS"Ol��C�R�cڀQH&i��>��)"O��
8:���1�1c���"O���2-I;�:��G�U�^��D�6"OzR��9h��K�Ϙ"=���Ц"O��&&�l:Q�	k���k�"O2�@�jʿ<8�5("��#�T R�"OvD�2,<0�XT��g�aϾy�S"O&Q��(�I\����F�B%t��"O8�t�Nz�z�r7ǈ�H͉�"O�ѓe
خ�4=�B�F�i�Ե��"O`�{��W�R���g�����"O�x�R&�Qb`M�1+D�j�����"OP�3�]5Vd���#6��ē&"O���IĆ^3@8�ew�b�b"O�F !I�6T�Vn+ �pXqt"O<�2�f^�3ܨĻT��� 	�C"O�A;����"�����Sa�Jh�c"O�|9QjO�% �!f�4.b��%"O��QB��4���Pu�4�j�a"O�9$^�H��@4��K&mТ"O�e���=�l18�c�	$�Ma "OpŸ���RX����!�
;���p"O43t,��s�����劷e�)0"O6��0L��I�������@%"O>���?Mr�U�-�/����B"O ��7Dׇo�J�	�6���!�"O�!K�)�r���{�O���$�R"O8�Z��ޱ5^��S�֘/��|��"O> �A�8s�����l�<p��*W"O�+i����a������Q"O��)Q�N�l���r@jJ6v�I�"Ob1��8�2ջ6Z$tb.i�6"O�t��I?:���r�C	&i�"O�����B�t�V�XWL��@g0���"O�9���5�1���Q8(��"O�lrr�fٞ��I�*��=�t"O�I�K�]��"��S�G�4$cT"O���������b�AI5/���e"O!B���5���gK�^T�v"O�����Z�y�I��M�����"O8@���ײ�v���f�}���"O���(�}��W�q^�-�"O"|"� �Cx�\�e�^�XU��q"O�t� J�$:н�T�Š8T��x�"O���H>l�BՋR�7J1["O�B��'`: �� �����"O�	�ʜ"=�,����ۏC�0�2�"O| �cMM�P �UaT�Bـ���"O�`2�G�Eq�T!�%E�x���"O��آ׆2d��Q2��K� �f"O��� ��4W�Sf/��K����"Op1!��>{�ahg ¸�*�"O�����ޥ���O�W�z�ڠ"O�t2�+ҙF?�4B$�۷]�H��"O��� :}�h1�'�Gr��@�"O�<Q�aF�.��� ��n9��F"O �IF��������ԅn���"O�@r���o�:��rM�/���z"O��8r"�>,|���͏�{��)��"O� .�hP�� <� ȀQ��K��]J`"OH2���?*�ȪvG�: ��l�"O���vo�_ކ����_(q4��Q"O���D�`�<[r�J�`$B0�"O��S��ʅ	��yAmT%}�P�2"O�x���.�2�9�N�m]p5:�"O�HZ��N�b�S��\�<���q"O�������3�Ȅ�֮��g"O2\�,طYP��aH��Ӯ���"O��h#��<��,��î�����"O2�b���a��D�0t��$Q"O\A��Ɋ'*q�0�I�#Fhe�&"O��K��]%B��%h'��n��8��y��H4u�0&����qԢڐ�y���+	l�����y��q��D_��yr��b>V8k��БA�JX�mY��yB&�>B�̴�%��H� �b�S�y2�f�D��A,�?>v���R��yR��%�Xݢ���%�����/
�yR�?t������-d(�4	��yҪ�*O�,�S��I����dl�
�y�I�w9��`MRD�Q�0�y�Q����N���� ���-�y�)�%O�	��N��tހ]����	�y��\���9h������yRd��
9b�aY>fX]�t(Q��y�3}�0�Ѥ��eڌ����6�y�*u�rUZ�*�&b`� �#�y�,Lg`i� ܱ~���S�B��y��O�gR�@����@���4�y(I��\�p/� ݪ�;!]��y�ƅ����(dN�/q��:G���y"�N�c��k��7��KΗ�y�!Zr�0�$(�-����L�ygF)���"�dX���G��yK�F����wGߘN�Q0�	�?�yr# �B�M�p���#C�Д��'���EyJ|2��ԫ<����%��Xi�A�7Ä`�<S-Έ(SZtHd����P��σ��HO �}�G�z��`ZM��ځ�K�?��ȓ)LҥA�/�'(�49�]�(|�͓��?�u�Ժ?�}x*�_�:u*�+@W�<At��P~�He�+d�}زcVJ�<Qg��~:�@��A�N����uwў"~�	�JMzQ�� 12����_����#�ɑ|K�l �M�p����[6U/B�ɰt��ӋV�w�L�80)�$>�C�I M� ��pL,s>�:qKT/+_tB��<�"��A�V�d��7"��B�	p*u1�)ȸQ��y�D�N�gf�B�I��-�5�Y8f4�lr�	�d�Z��d:�&K2ٳ����d��8�&[?���ȓZ8ɛ��G7.�<���djf���'1j�Gy��ɜ���a��&�3]c�Qi&)�:|�!��L�
��R���t��i���z��'�8��dQ�a�64�C-����0�R��}!����W�9<���  �<�ȓ��2ю�!B�D����Ee�����
��܈&�l�x��@<;R�ȓ*��3E�6�����	ٞz��P�'�ў"}�%da�`p;�ܛN�\��C.�{�<)�B�� lp��A^���K�t�<�T�\n�"f��"�Z)G$Ct�<����87��@���<
�d�t�<� ���'�N-���^u��HÌ+4��P�B.A�5� +ډ=��Cv�9D�dҶ��C��;ǈԓ	0���Q�*D�hPAI�'*&�@��U��uRp�*D�x��I�Z�� ��O�(Lr-3�B*D�4��:$ʁ8�D��T�4%�W�"���<��!�N�PPn�;A������h�<�`��;1�̹j�ő�cR�����O�<���D���mk��K	�¹�NM�<�FP�|cB�'�X0tݪ��K�<�5GD�zM�N�;w��I�R�D�<� ���z�{�f�4��� #Q|�<����fL��⚯X�R�Z�o|�<��	z�
���,-HT��гa�t�<��bٙ&Db���L¥��q��)DG?����.]������-~`
!s��ͩW*4B�ɭe���2C�A�V���͍G��C䉷z
m���X��L�-H�ͲC�.*��`�	%�"�?�C�	95��1�@ˇ��: r0
#?R�B�I/-�ڸU�C��:u��[�B�	�sƞ�8'���@o��B7,^�"<9�'��?A"��V���`-ߪY8`o=D�d�f�������e�Q�l;D��CЁ��%�� ц�";Ar<�o9򓥨�Bq�NN�u����"��,�"OYS�/�2[���!�` +,Ќ�"OX�ק��5j�Y�b�Z�@A3�"O�Рp'�N�vIV+2'���"O2q�b�� �Az���m_�t2�"Oz����e�� �$!U��"O&	���*^��`smτDܬ��g"OTiZ��H*(����M՜�r�8���!lO��)�ʉpP��{&��P�"Qi��	��<a�P�Bx��!��<	��y�)�{�<9�������Ȕ8q���-�����'n��P���Z $H����5��;�'�(�l؎i�}����)��2
�'�ll!�E%��;$�V�N�v=c	�'�x|�b�N�|2(���0E6^%*
�'�ZYH�@�bAp�9+�����O���&<�& Z���]`:�[V�UW!򄌻i	r������\���L�!�d�!�e��m@�+�F�#@i�F�{R�$�4.�XH􀌫�vd{��(�"�$/<O�C��|(K`,sv�;�"Ob5�Pƀh2X��
Liʁ�"O���pD_6���	�44� 40��0���i�VUi�� ��ǬA+zPB�I�+�dH�k��J .\��*J�c�B�� [.\qQ��Zq�q"��1P���T�I�e�q	�H?�2�)�i�rB�Ip<Z ��)����QFG�c���|y���~*��B�5[w�OR�!��K�R�<% Z���Q��]e��y�TʒK�<���.�@��1l&{p�Q�.�]�< .�]�(b��N�ŰlA�@u�<	��V�9?Dt��C^���� �Be�'nў�'#qĕ�$hV�Q�T��#�U}z%��F�p�;a�A�S�$�1��ڿ&�>Ʌȓ�,AcT�آ3�l���oο;M9��q6 �o�Zl�Uف�ֻ0�:��<���	8$!���5)�8U�|Q'�0:�!�$O�aĝ`Q���R�Zu&B�C�!�� ؑ�!�ߝ1��X�j]Pơ���'1OD��&�eDY)U�� #S��#n�˓�hOQ>=��b09�)c
$�FeBc�<D�D��/A|O����J��a�	8D���T�<+X�hrLe����@�v�`����G�fe�UI����9��
8x%�B�	����@)�e,�كD	ȈSI�C�	�4V�`a�:z���ɒB�PB�I����Ђ��3(V ����e���&��P��R�N���u�֨��7	)D��[PJD0�(��j@^�`c�(D��Y�(ڣA�\)o��	V6<��İ�����?xD����1�����n�B�əHir�೨�S���8'�@�`�B�	�}j.LH�M@	?���B�D���B�
>-�2�e�(6�Q�7��O�d��hOQ>QЃ`$���$Bͪ�.t���9D�x�bΞ"U�X�l��H9p�g=D�̊�&,:4�PS��
����";D�����=���[����|":D�t�v"�<KѦV�	Ҽ����9D�(BE�=WT�w�2z?tY�-*���^<8FNU�q��D�P��<�ЄiQ"O�xzf*V���թG����z�O�<t��,��@�` bA�52�J ��'D�Q�3��?)r�� �)2DE+�''8��N,��� G��&�^( �'�d(F�'<1�LHŎݫ.��1�	�'�0\��,8c(��$�M�8F،��'.�����&N6� �oP=,�^p�'�f�a�F�a�����#�"GBt�'�����F�z������,*8k�'��b��Cx�K��^%�r�'V  �O�3U�z2�։���+�'��}�0D��̔ͩ��E�.8�
�'�z)3�R+buԸ�F*�5g�.�2
�'| ��X�)�
��C�%g�ʔ;	�'r��k	Ю
�N���=dc\X	�'+N)�fNF;4�2Yq&�X�����'�\1���}��T��	Y�>���'J�
����0�D��JK(W�uK�'3�y@ �����i���G4@��'	 �q��9$ҽ��gO�G,p��'�D�s� �,�v}����<���'W�%CJ�Q bQ���x@�0�'[ę
�N�*�%�I2��s0��z�<���Q8H��ĩ�)ZL��ѻ�J@�<�DЦ-��) ���nҢA���}�<A�!�$GSa,\ip�9S/
{�<���z�j��f��~�p1H6f�w�<��B�?�ڵ"6%��w�؀p��Lp�<�c ڍF��	b!єs���pƭ�m�<���1)\(#e<fZL C��i�<�ʊ�R�t�U��<��dk���b�<��KL�e���
N���e�[�<��(^��*�~0��82� m�<p��9Aʵ���N�ͨB Mm�<�S	��V(�#��:�pZ���o�<)��K�y2���( _�4��h�h�<A�8=�4<�IK�<x*e�L�<�Amô+�x\�s)O�k�a����F�<��I�lNY�� !h����]DC�I4n�(��(�-O��6A��x�@C�+���2T�E�D�5ᒛd�ZB�)� �y�F�Q�{Wty�%sZYXD"O:����%j�}��c�Wh�d�V"O��+#��6.%��'�:e����"O����,�vm�Ɵ�xdDM�'"OF�av�D�}o�,��U�F�{�D�+R�X���U�a�R����HW1O
U:�A�;�.�84C��\i�"O$�9�E�,��h0��&���S�"O���`O!}���5n��=ZVD��"O�� B/KZPR�`�o\)EC�+�"OH��$l^:	 Gj�ҭb�g6D��i�#?
¨��f��!����*O���֫lD�\Ǎϗ�ܙ��"O\�xGN�l3>УcLX�*ƨh�5"OL�s�<uҬh�)�)e�"�"O� ����8[�9��hB1y���:d"O�	�Q��{��ӑ�Z����k"O��3��{��pƅ&K�t�0"OL���7 *��p���\�	"O4�!B �`ml� ���}4��u"O�T0�#����%b��eS�"ON������p��L_LDx�Q�"O�|��JP2�\ D*Q�ANvH6"O�]�� ^7�xE�����#����"O6���]:i�\�ۖH�Y֬��"O���(
z{|�R��o��y�d"O���n[���\�����bH�u"O�� w����*΃2�B-��"O&��0G�I2!Z#�H�q"O�EQR�F?m�8	��ǋ�}�0h!�"OX8X�
��D�|`����lNP!�"O�9��j[��<�s��Z\���`"O�g�R��;���2V���V�'g(m���
�"%s��\mטG�������퉡t���z�J$�rU �8D�@��'�		��b�	&�<�)��ل<z��0�`N�E��pK��(��wb!���$�^e`�%�5��]@G�w��|RaA�cP�%��Bט��5B�S0�ց���ְtPmJ�,�F�<�0���)8nd[� 5O�����̙obJ$���p�����ቼX%��O0�ʈpT�U�7�v�+�%q�����-5�HV"��a�E�61�@�v�6��4�M�w(h����W�1AtĠ6���TM	s!z���45Hd��I��H̐8�BV�I�xm�Ok�	N�%���6�� ��?�!򄜇ex��i4F��x&�;��	��U &��@`V`@��8w*tȀ�Oy��Q�Ts0�c0��G}�A�\����T2�<P)�LI���=1c	�F��P�3&S�Gvv�)�k �;���=?�����'�ҳ���>���˚?{l�E}ŕ&���k�C�� ���i���'�8��F˨J!qQ'�F�'�50���$m���T�� ,���	di)U
v��*Z�o�^ ��M��p?!w��!.<|m��yǲ�`��[8paD<�#�F�m⇌Z�c�[�FE�(1fYs��Ѥzö�������Y�D����.B�<����t�<)!��9p��D�� QՐlz�/�3��K'��?<5��$�L�S9r��`�3 ңW؎PQ����@�h�8Zy ��@�6-t ��g"�d�6,v��'E�b���GR [�d�2�|r0�(d�W O%rA�	:]'�|�t�N�2 ��B��R�������J�`��ȃ�H(Q�DI�*K�}�86�X�\Ƙp�"B�&����JP�a��E�lɦ,&d"J�3{�!P�əZˀH��!"����G��]ɐ�
a ��u߮\��)�2;t�`���'t�!a		�(�;s&2;���4m����0�!S=6l`��ɀ�J��dc��H:�c��V2;���D�����Ȉ��ִ2�Z�s5�%W>���fJl���]*:�&�ʑm� Wl��$��+f,�"�Uz�q��h�� G�	p0bGY"&�a��'���Q�ě�.j0ɵB�Pq�M��JH�5��ơ
��:�l��@���.�R1���
)�ÊR:(Z��� `��0
Q1?�(���!�h�L0��C
ƭ��錼i6EÈO�^�(�� ��9N����F�7������	ؑ��-��!؎0��VY-�up��:��I2���& |I�e�Xp�����
 �&א9HB@��^"�E W�
:�
���{Tp@��C	��c1Lbb���ǅA�f�6�,-^ȹÓxw�m)0,�S���Kө�&��lx5�_�q�<P0����5�^�z�nO�Vq��W̃V���k�	�-#��D(��^	u�,xXU+�}q���e��	�����O��a 
�g�ht�H�3hH����^�}j�IqDT�<�@Ԡu \�*=��"�R�)��/�TI�qNӼ1F��p�ʅA-t�B�N��$�+3�ȑX�>̺��[�D����fĒ�剓m�i`秞D,dS���5�p�f�ux�m��y2N0��L�gn2�ʩ�R�L�-�~�a��x��	�i.��®ֳ��p��@����� �!ɤC
K��I��ʹjv �Ĥ_J'*��/�5�����BL��d�i��-�c��w��\�qȈ=&�^�#�b�2I���vD�f�'�	�1!��x#Y=n�N�	�/@�'NΙ1!�S;�� �L�
?���u��$"��	�Ý�Mc�'W�C�fE�D�D�8�n���ػ|x5#�VJJ��j�2O�T��ř�)�L1�P�� '��(G~���.�Di���^=�%g�%p]ɇɁ����q�$��f��}�Ļ���2�iBLA�iTE��� ?������S�#���E�{�l��3
������I��`�6���96eS�8>���F,{H�k�؛dX$U�C��p��1���m����ի"X��*�m7%A��
��^�:�aU>i�8���Qb���A��)!P�'�P�6�N0u�q0�C�4_�<A�m�4k��S0G� ?a�%���a��l���2 x�MHp���[�4A�͍�i�� A�ѓ9	����Хsj�a�2��3^
�s�λ A�_V8�p1d�vt���*��8[�Mi�!�;��1�G
u�@��#���H�3��uq��תԞ?V�]A��:�˒:T�����l�D�Jc�
=6�T�I˓R�0�2�`T{n�2�]�pډ�W���6A����n_�o���%�x�x���X=Z���f-O�^ޅlZ/`��k=uи�Qf끹���zWH�?�*��ѫ[� !����ɭu�괡�Ø��Á�fy�R��"Eu�<����_#F�`��>b�Ԅa�~�"��5B����&�M�Bz� �G�Ҹ\'B�<��F��Nr��&я+��%sdCY?�C���5�d`y��X���x)s��?M�`{SHƖu��!����`K�$�-W̓��u�ə%CZO�����><u�(��0=11�Ѽy�Ƒ0"n�3��dI����|���	݋&���Zs�̗&�x��ĝBN/3��L�L�?�2�1G��ai��A#�D���#ba��o(��P3��[��ә(�r���AR�;-�ᣎ��e�a��y�����扰x��`9��&	��! ��F��;b	�K�؝�F����O|��[��N�α��쑉>7v�Y��k�mq� ���NyhVHI74Z>ݩ� �T��	3BH���iN4º�R �DCh��r%*G�x�PE̽Ho�$�)n@����/k�a2��ċ"2L|����Q6|�V>5S�f� v^�bgk�6�h(�sAH�Uj�xׅ!w�����x?: Ѕ˔縘j��ɳtDα��C�^�D��q�K�@u��~:C�֒��1pL��ګ9j��[B���sv�䑓�Z�/1a�E��Tt�X�cA�%Z�#
ʺS�����Ŕ;j@�U+�)9���+�nM/qJ^D��	hL�r�j 1����u��*((�?!�KU�6����n� 0謬��O����+�]��EI2��(E�0��'OT�#jB��~ ��f�"g�9��O2�X��ͅ+GȐc��Ɋ����y��n�mu��2e h% �B&"O�I��T5	�|�
0��Fs����:��Fq������|��J
)�!YCǍ/B����P�y���3>D)��͞$�Ρ{�Ɍ��y��qAxՙ  �m�ɒSb3�y2���@I~}�iV��k���y��pd�5A���=V���X?�yr� �hL�0�`d7*x��q�ń�yrJ8Lp\ʇ+BQP`�!����yriHycE ��D��Ԛ��à�y"a�089����2Z����
��y��	) ��p�I�"4��m���yb�D�_7*�c��krh
�GP��y���dMA���Z&�YT�O��yR!�#L�\:c@��<��t ���y�&X�(�F�Z��-?0
�
��P��y�lJ!na���g[�\���w#Z��y�,U�h@p@��H���CP&�y�`�T�:5q@�4d\�9�j:�yB��S�L���]~�JS/ۚ�y�a�^��Bm� b����u�Έ�y��5X�p�Ѣ�?f�P���AF��y�풣QL��
�b�а�;���y����j��	�r`B0)�-*tO��y�N���x��62�Q��Y��y��=2���S	Є�B���=�y��J�dR�<;��B�����0�$�yRJ�"�� a�o�,Ѯ �gʊ��y�l�L������TD�h�G���y2NG�-l�ɺ���	|�&=kW��yȋ^ļ-�g˰|��YceW1�y��0!X�p8���r��2i���yR�ϋ&�~��g�G+s�h
�*Ő�yb�E)�^�;".�+$x� �*3�yBD[���@��%Vx��1'N}�<� �Ps���	`�xs� 2/f|�q"O�ųao�W�x�
��/4��"On�r�ߌm�*���]�=T���"O�D���/%�̵�gN�1�͑�"Obȣ���
�#a���Ĩ�%"Ob�R��^3:���g��`�*"O!	��%L(�	��#s�tK�"OE�������u#�q��Z�"O�JAfU��X93��@M�҈a�"O�A����-���{@�$w�e#"OJ�W�t+���`͈8YP�
�"O@8���8� i�j3B�؃�"O�CBO��~�8D�E+A�G�<��"OXq@���7*�L�)B,�f��q"O�t�`%��ChM��z���K_�<a���6,���۹ho|�`Ca�T�<�ӣ� �PqISDޏN�a��R�<%��:�*�w���u�|IBƓg�<��CE*��@ S ��&(ϓW�<���*������R|�}HЏ�P�<ɴD¢5�v�`�o^r��=���S�<���@�Uc����N�EÆ�d�P�<�fW�S6�=ӯ�Df�"��k�<��P3,Ryp���S�0�j�<�1+�h�<aR�
><<���ԥK}�<��)��B� -J &V�Y�T]
��e�<�㦀�Tj)c��1���C�Ņf�<af㍒FtR鈖�y�ӆb�<���<-d�t�ʝ��蒵ir�<A�/_�}�&�ŨA�.�*�e��K�<Q���D� I�"�J6{Ba	"DX�<Y��w�IZ���#���Zl�<!0�6�mQ��R�p�H�P��i�<!��^������G0O�2�9`�m�<��+3[��b��JJ��+�B�<�%���F���@�;=�TX���P�<�N��V��q��Q��H���j�<Iv@�6���%f��l���XChUh�<��K�FV@Pp��(B1�D�Bh�<i�k����EP������
#BXd�<�Dk	 p_ZՒ�皓7}�*t�<�%J:?� ���h`�3b�H�<�&����Ag1I2�l��ȃ~�<Y�m�	���mL
�%��_]�<qF�ų8�����5!��g�<�6�ȍe�ZҭݠG2���hv�<� �H�JZ�7��A#��foY�<�&V��}��c�:v��oI�mB!�W���z��3t��8a�N5t?!�d@쪭�U萑S]�*`O�1!�$�+g�8��� XD38�
�ُn!�$�1h���OH�q"��	����!�$��C�|�UI�- �ء���p�!��V�V��$�ϋ�a��4��S�!�H�T��������@{�F�l�!�9e�x���	z�pi��fѲM�!�$E�h�jp��Zn�:U�Q/tI!���#�f%��h���q�ʹO!��N�h�n`z��EB���Z��|�!��;V�-��cN:8x0I�s���Pw!�ċ�Ia`�@�g��-g(����;^!�D!v�C�V�T��A��:!�D�`���R!7��â�O#'!����:e�5*��tF �13��,~�!�� ��⣉_��>��r�'m��+ "O��2fiS�z�>���,ʷ{���"O@�bk�4�n9j]�_�����"O���FF�)ۃ*�#`�	��"O�Qp��_�2�񀙱*X�x0�"O���]�X�9yP��{+�X�"Op@������س
��7f��V"O��u�G���5CC�:@ ��3"Odq����;dZ�qIr'`��q"O�ɒHۮ���B�W�*��4"O་����[`�����(a���"O�u@thR��+�6\ј�"OjY����p����j��:�#�"O��@v�$Q��Y')9IHu"O4{d쎉r��U
憛���q"OX4�"��*u�|��"� +h �I"Oh=kM��}BZT��CP<S�$��"O���7��2�ꠊ��n"��"O�`�+���q��Sxy��b"OL%���w~~�b���Bh8�"O�5Z���V�T8V�)e� �"O�iaQ���PLr!(�4iR�a t"O�5���^,�f����)y���"O���H�k��H�S����"Oh��"�J�"IT������]?!�D�2��(#�H�IP5+���r!�$�%̦�����$�ܡ�bh�+c�!�b׶@�e��,�@�xC��2^�!��U<y��B��W�a��ؠ��+}A!��ì��([X�����y�����'H�Q" �������5vdea�'����Dg�f��XR����8�N��
�'Œ���gV"��'F�>B����'�|c$���Rɀ���D�-��'���pq&FRX�d
� �+N���I�'쨘��O;��k %&w��
��a+��锃Z�R�i*aG��q���X�O�"l	&W.56���l�"O$�sGV�)l��:�`ۈNtA��,=sl媲fX*	��ȴ�x��S�7�T�X�yBn\�W��T*� Oqc����-�?�p>9Ç˶3�L�+�(U�=�d;����A�V���.}�m�@�`x{���i�,����'fB��P��(�$2x�+�]�'�fՂ���3��{�5�nي۴P2=��N��r霡 �6a�}�3
�!�\�&��%KԙIR��`R�G� ���a kX�V�Ѵe��"mj�@���4��E���KQ��'�y��I�1�4��ЈY�"k�Qc���yҷ�D]�h��a�$��,�m"Zܩ��7)����C3O����FQ�bh )d�2(�DLH����φ1kdx����s��۴����{��:N���1K�7f�d�C DrH�;	� g�����i��G�(4*�'�?e��!8f���~��$p��38���Ǆ2�~���d�$��O����Ҁi>LHBAJh�*��IF 8�fú1<V���G�=P*���u��KC�8|�~2�(K�.D8vkG ;HX}��dT%���4N�d�h8�sd��8E\iZ�k��L�4pP��8NPu�'�yg�Řt{j](��(��Dk2��+�y�g�E���"��Z�{0H��IT�;tl�2ċ^/Q��=� �Ry���D���juo }=t�!�W?���R�7�ܤ�c�N�h�`�(�Z�I N�l�p�h�i�*-jc��*1:��do�C�4��v
����Dڗ�MJ!�X����8�4����&xDĸ���J����so�)
���>aG�οv�6;GM�!u:y�tJ� t���K��S�q���0gSN�b"ת=s�()S���$x I��jעp������2L!�� ���3R_Ɓ��aF~��4�T�<�OR=I�j��E���uO�W�� ��B5p��!UXl��/�)c|x��i�RnB�E/~�^�jV��L�(,@ՁG��b�Ȅ^���s&X}TI��ɖ:@*8��0�n��Ӫ�<q�nї_�i�G�-�
Di���3�U�U���uy�ђq�sE I���[�1g�\��xw�O�H���"<;^�*u�A>t�,�^��`�k4��q :>�$(�S�Xy; o\&�����O�;�Y���S#D@�R��"j;���3�Q�H�k���T��uu�{��\k��dL�Z�4��� �c�~��҆�,�и�U,��c��+n*�B��
]�*��1��0d�f葢f�-���)әX
(�օS��>}�B���$��@��0>ei�/�x<��*VN([d� ����mG�A��0�B��Dd�,����mǲD��(�"E0@o�h�L��W�`s� ]I#4\�U$��(���z!�Ɍfj�T���Q5�F���
D�FX��5� @��ZR*�&L����E��~}(֐V� A�d������b��A#w�lQE��%JP`�کO� ���{0�9
T���ZH�l2w_��8��_kt�B)�>��ٸ�%�f�����WѦ�ӟ'�v�w �S*L@F��	%���)���x(�Bu��g �`�H�s�џ�b��ֶ@=|�
s͞)��i���tYcc�+6jn�Q,
��Qow�d�j�M�!;�-kB�S�Z(������k�Ȣs�O/XaV�z�M	�.���I/�4!��BB��34�#�"xre��A�"\d��
�B�\M��0 P�.�T�S�(A�C�i�TjO��$qВ�E�L����ҟD�|�C%U(��OmEbڱOv ���OP�J��g�O�"H�`ň���d��L�4�b����^�D!K�h���2���I�<t��%I�qO:����
D8�&J(WX�5�Q���0.�S��$S�C�^�>eZSC���xq�J0A1\X�%�ҝT/P��+q�h+ cϺC��1�@�]
�*�H���=�Q�߆d�8T;�BU�~����Jї��uxVMô -Z�G�ȯE�Y��Ka�"`C@��x��
�
������CP0��0�ԡ��-�Y���YH<$,	�|:�qyAE�!\2�q���>PI�đc�]�8��C5OY��U�	<�aY�� ^6�m�dE]�UB����CX#z;��cG4-!X�:w��'o��yrg�4,#\�*W�B�n���CB#d�y�%ض&0u3$�9;(4���ZQQ�Q�⒴D=��ˣ ��o�5��Ď��2��M�- ���aD-VQ����Ƀ�)�>�� �8Xب�%O9�4�#aBD��B���"�t�I�t�ҿ)^�����9�p>�s��3یŘv�e.v�s��SU?�&�5fbA�\�3���ѷ��k�xx�&��2ڡc�ٟ� ӦE�2UL�}��Eb�2�3�"O��Q���"}�D@%�]5��mH 噘BD`�yb�	�S/�]�̞X��Y��&�"��[=`�(��w3N��"$@��p�	i��3�'�OH��As���Yo�� E� P��2SO҃Ȑ-�`&މd]r(JuK�7�6��b�Dy"����� Vi�Mw�p��
�ݨO�9k`�f�L��� �2����Um]3i\�a�<T�9���(�(\i�&��5�s>�O`��#�_q�� a'ع bf�`��O`���ي>��)A�#G1���!���YZ���sL\�01�S�xΐ�T�
o��I��2�zB��1I�x��d\�L����s��>s�d��\/N���ҳl�=y�O� ����%y�(�TԤ����3� a�l��gޔe��	2��UKWIR�+��uAĠK�J�:퉆�K�W�(}��h�G
�$���S�i��i%��w�'�J<d�L�a�-��&kv�Y��P�04�@����A���1$e>��l�H���� ��Hjz!b��<D� "���*�>\a3(A�s:xT�$�7?��P�N�|���	�/%C�~r� T� X��t��=���p�G]l�<��,�?f�f���#��g	�(����͘'� �ըR`�g�I�$X��m�%t� �Ȑj��*��B�	��:��m�N���F��U�C��(�{���=s � J�6��B�ɟ���j��ZR�ʝ�Ï
l��B�	$&\�9Idnx��8��%�B䉦v��Cǟ)����4�ȾV��B�ɴ(�ȁ���M9l�p�C�bӨ@P�B��0����v����iqsM��lX!��"@k޹�âU>p\� I�j�Q-!��f+PP�F^�a:�eh�*�(!�d��(�
4�DP(N�F�kw(VY!�$
���%P�Q�4h�Fȟ[!�D�?}���@�J�u(������t�!���;.�RIp�A�2�XU�O�o�!��La��:�	�\
x��C�D�C�!�:W��v�5U㦰�&A�  �!��.�0[ӍS�r{��0'�ܝ7n!��O�\E�Ν.����o�<h!�d��k"��٤*�o��ED
�G!�ر	�V�cW	�,7R$�r�7�!�$W�/�,�[d�HoD@�b�Oɂk�!�$�
�򭈵)IgC����-�8}�!�D�-Qp8�GMG+'X(Ң� �,�!򤒵,�>�5F��&�}�1�O�!�ĚH�x�F�-�ѩ�R!�I�4z�5�U�4�!����!򄝢t�8�s	L�("^��t�q$!�Ӟ6F�8򄕺
~-�T��= �!�$�!U�L��Ę+�P�0��_�!�� hp�a��>��i"���
P���"O� ��
�P��Q	�o���"O���
�J��as���H�|4�"O�<��
�.f:`��(گUH�;"O�)��!�;��܋�U�W&����"O��p6��9�iKSd�C*��"O�l�4��xY��G�+oZ�,!��<� ���+82��N�,$�!���h)x]��* -}�r����!�5Y��%���E�<�q��{�!�d9��SN�0�XZU'��{�!�$��F~鷠ܲu�l�U�4�!�Q $7]�"��N�HuZ�%�c#!��a���  ��<�RQ#RD��u!�C+;b���	�V�H�(BԘx�!�D��kbP����g��-�A��T�!�D��$�|�+A�T�8w�@�!� 
!��U�/��L�ײj{�!`d�̾!��R�r�|��Wj��=��`�"�!�$ӳ,��(*Au����N�u]!����Q�ħR#[m.ԉ�� X!����xx���E��Б�F�I�<�!�^�挚uūb�Ы	�n�!�$B�`��%�V����R�i��S�B;!�!�(\X�G؂Z@��g�
d<!��Z�pFjY� �ɏKAʡ"�K�<!���f�H��U+ԭs��Q�e��2�!�$=���7����`�!��`!��}�
�*�S5G:���L��!�ǂcҜ�dD��1n:ac�Μ�-�!�W:@�L�"sG��`����� 	�!�ĈW��Y#����UztEK!�;a�9QY��c�K��y9Լ{V"O��Ib�ޮ*�x �H�>'�0q*Ox�[b�_'��$���H�=�hݲ	�'{X�S�+���X��!
%/hЉ�	�'" b�@�1�, ����S���
�'w.(VJ4o$�y�F�,IBZ�9
�'*���&Ā'0j�#��ݻU.DPh�'֢X��l*�VL9A8NBx9�'��8�򂟖e�t��T�t��'����F.A�U��(��F�#g�
<i�'Hh5�䎂�c��LIp�����xy
�'����u��c��Tv
pX�',�E��@�B��aEF�c�����'h~)�#�ڲA	�آ��7]�8���'��UI���"Fz��p�&��H� )��'	6aÌ#h=2.�4�*d��'($yZB#�;4@^5��ս$7l�I�'�m���м4������&)�ܹ�'!&�X���hдXpBiO��2�
�'$�z�H��d��J�N�$��'_�1���C�q��ؓՊ���'�~�C���2��<B�6iH��q�'���D�u/n���1��1	�'�j���STt��#�[�	 �'"��H �҈e ɳ��opҔ��'���R��n�8�H��Ϭ��`�
�'E،2W%ŒD�ݫҡ�/�c
�'�� �#�ѝW�֌0�#�����	�'�Td����eݲ�O��})��s	�'�f��@]�/c�+ܔP�Z	�'Ǌ0U�n��H��+��S8�$�''&��͙�pؠ2i��R=3��� ��`���1زc���2�@"O�%Ӆh�fz ȤL�7{"�R�"O��@6�P1<ڕ� �";��x�"O��r�P�B h�K"�G�;��ib7"O��K5�ؿ�}�j��pJô>P0)��q�^0�TK�45IL�`' =s弸�ȓV�&����O����Fm�c�<u��6�h��`T,u�r$�A�K)}���  z�܎PX �qœ�(�n����m���]�:�~U��e�k2|,�ȓ���ٳa���0@K�B�B��a�ȓ5�����(�a�أ+ud��[��-Y�b��S�X�Âh��n,�̜T��M�c�Ԑ���G�8������	����2h���	H���;���� ���l����p!� z��'�vd6�����7|�q�Q��8@@�B���:>�y�����0|�V˘(�����S�4A15`�R�~����l)��(����|و��3K��9� ��>	sGր}r2b��z�NJ>2�,��*­k�d`x��Q�<�3��Z� �nڌ�v=����:��H������֬m`��$��?:��c
*-]n���&֊���?ɮ�ؘO��9���	ti;Bi����X����~�[�@2�C}>�cd�GB��E��]P�c�%�ص�T�%mb�R������!K�[�C8��)�ӷR}L��&��:�ҡF��W���'8p��c͢E�1O��0lC�FHn/�����>����+��ts��_<J����蟸Apɕ4D,���/D"�>�:��i ����8��O�Y�''���A��=��%� ��E{�_}}"X���'~����E	��i��ub�J��4�>���Ҵ5���*7F�()W�� @(ȘoOaq�΁H�	1ޜ0���ԟ�	�`�0f��S���rOU_�X˓|[L��J~r�:O �A�kڧi���L�/�@�f�'��y�&�O|= -O�i/��&r�P�!���&�J�E�e�Hh*g.����&Q��$?�SR0A��?������\�h��H
G��B?qD��LW������$6m1 !�5C�H-"tTL�#?tv�O꬐&gN�~�
� N��>M��Ct�����	"�ʐY���<A��K�#&RF9}J?�A���&�����0v@Γ�b����<Q�y*�qO���#|�̌��J�=: ��G��y��0|z�a��Sn����NC� �N�!�w�'�L��S�2�^�|�'Ԭ��a^<i�
đm?��qE,��H!�D߷	'�Cj_�l#@�`2�Z T!�$���T1afY6������7d�!��]�7���QV�S�,��٫�P?Q�!�d��)k�QB!&�(���©�h!��2_0M��0vK�L����'I��!��lî9�郣@-b!`�'�B�#�#ԅYݐA#5�ّ>l� �'{�I�b#�UfL�`ބ�I��'C��"�(P%!�$��'�* ��'�n�ɑ��`o�	1��7N5+�'9�vkD�M�2M�FٳEi�;�'��$YR.E� y�Ó�Q ؉��'a����d���Oxp�(G��y��8}L�G~}�<�v�b�<���RE7�Q,�:k���di�I�<	�����Nj#���1D��j�B�<i�nK�]��|R���,Ʈ�m�<��.T�!����J�&g�n8��a�<q�&ѴbJt�eO�!0�t���CE�<�Fó`s��B��pI�|y֣�D�<I�͇�a�r�02l�se�I!�KB�<ɢ�I�_�آr��7+��dF�A�<Q0͊�!Z�쩐�:�X8)�o�}�<f�.k��
�b #a2���i�w�<�@ͽ5�I��G�3|�x��Hm�<9���h�t��ؗnHx���r�<�4��x�x�:���Lz�L�7�E�<� ���&�a�R(a�M�j\�aq"O�=q��?x�ȥ�PD�ZnQ�V"O8�����L��(� F�3Q���"O��`3�
���$��\*>��#"Of��3�_�Tʠx#���ڰ`7"Ol8����S��pR1�T()��+�"O"PRD�G�[.��j��I+5"O�M��
My\UjS����h��"O�e*C`� m��C�o��?��8�"O�p�Fc\,�<a��O�nx��)D"OV����@�8YfL�tAE
p�*S"O���I��3 �ü]@R"O�ua��Ǣ3O(�a��9��}��"O�*f�ٰ
ԡ'�o�^Qd"O��C��N��� ׄ���v��"O�̨��M�MnvA0Ɓ�f4���;D�Pʄ-E	|�bYr&�K]~����c9D�P���+ِ$�Q� R^p��i;D���0��%���Ӣ,v�1�c"9D�|j����U!0B� 'T��8�(:D��p�
�B��R�ޡ%18�s�o7D���Ѓ��ڡb��RL92�$8D�����ۊn�f�
���T 5D����x|N%���X�I(88rDg%D��д�̐�q3R ��^ �SE�'D���`iTO�Q� l@;%p�	C�.(D�$�U��/x��RO]%\ D2��+D�8J-�#=��`�f�;ƚ���(D���$a�.�iz�_�%.3B)%D��".�2����E��}���7D�8a�$#B-B�� 7L��`���5D��;�l�$TR��ؿq@�d��� D��@����O�q��QLr�U{��"D��꠬;|渁K�LN�o�|��3D��b&pf�@�*@*Y�}�$?D���ҋ)<Z͘G!A4��%Ʌ�9D�@���T�3n]�>[��V
8D�@��+�]�zp[���w����(6D�D�@,ԄV�S2�ܘA�����3D�l(Ї�69x8����(KYB!��P>\�<��F�3_��Ż�-?6�!�:K*�Q1L��8� �X�T[�!�$��9�da(A͒	�����ғ3�!��	>�`�yT��9���1�*�?Z�!�$tth�Rh�$谅�o��!�D�p�
Ȩ �
_�KJ�hB��y�'sJ�B2��"c�8*W���`J	�'j�$�B�՘C��)��:����'��J5�(E��4�Frm �'���Q���:�Гj� ��4��'C�� ��I|&er�MX>l� )��'�4x 6��?���"�Ǐf&���'$"�:�D�R����5��:�'��u��1Q�u��K�4��M��'�� H�f�":t���$\	�*a*�'-C�aN�=���â-��\q�'���AF���؅ϙ6)S���'g���!
�[�`��U�&�\x�	�'�]zcN�2_�$�[u���3&����'p����Z8 B	[�J�0%�h��'Y�07�^<~Y���B�
$� m��'��iq#��֌Â��10p `�
�'M�$�UE����
B/E0r:1�
�'�X�c���T��6���l�]���� �L�@�?g2�D�"� �xi�a�g"O<��]7n�J���� ,2^�0�"O~�J6��^L���W� 'C���"Of-IP�K������*� Qj)x�"O�M����ht>�8"i�T1��a"O��Q�Ý��ř�
��?����"O Ie�[(���/��"��l)3')D� JӅQSw��{�+[�8�DE1D��h���l�(|�GD>N��͊�d,D��臂@�w���#�3W8��E+/D�����&j�HD�%څHr����J,D��c��'��ir�4y�`�25M=D�,qfN5�28�&LK:R@��&&=D���Il*$M#a�֚8f��d/D��3�M�(]�	-��z�4�D,D��@@�9Hܠx6l;*����E�4D�x)7EI�m�j�hǞ3n�:��2D��y0�[d4ܑ"��F�e�vx��'=D���WB��Q ��[�D^bzL�b:D�X;�^b��p'̓*��I�F3D���a�B�t��.<(��/D�h��	��f��)�f>
<0@�/D�T 5��/]��@P�/j-�!�R�2D�(�����s�8��s��o�1F>D���k��u��x�W�\7Iy�B�1D��iS�RWL�-Sgh��ہ�#D�pi���`�Tm\����,'D�,�ш��tW�m�g˰F��Uo/D��`q�?j�@t�J1E8���d-D�X��d����&-�@f����(D�4��+L�U$��7
@;�<	�)$D����&ؙ9�x4j5���i�LR��!D��YD)_Y��rfG8F�Tx
 �2D��
p���(3�a.\��볡>D�X�C���T�Q���6j��l��;D����f!:m�89E-^`�05�5D��R)]�H�h�D��1���&D���h�1��f�_�u	!�I%D���j��N~)�1���O����1�$D�dh��ū�F�Yfo�(pؤA6�7D�����22���� װ\c�L;D�p�/ .3���H�@&NQ��RJ9D����#�
6�n�K�F��Gd0��a-D�4B��/��m��L�x��\��#=D��cA�x`�t�dn�S�&<�G;D������}In4�4&�&N�\���;D���1���"`��h6Ö�Y(�*,7D�����j�r�AG��w
�I��?D�`�`]�t b4'�����A�=D�T�s�J�e�`"��Xrߺ�!��:D�8'�2{�n�a�fW�3�ˁ�<D��B���'4����`GڷJ:�PC� 'D�HС	I�k�H� �V�G�l�A��$D��n�#T��ą׎o�.�K�b	@�<��! �N�B�B�mE/Maf5�«Az�<	���z^�ꆧV���bЏ�x�<�E�Z
:,m�!��2�&����Jo�<qdo��*s2�S���v�<	�b%=�6����ܬ+J��$I�o�<�E�� ]"ֽ#�DI�A�<ARb��Sq:�0���"�`E��!Uz�<1��ǳ2�<8�G�@4l$��S��t�<���?�q�sh� �*IiƎZm�<��"�%�x�X��N�V?``��i�<� ��{Oé2G�Ÿt�=4A�H+!"Ol�Q�-[�t;�5�Q�J3)�Y�"O�U��$�dւ ���L�#$>�d"O$� �F ,t�j�+SmزF���1"O�|a%�Ɍ��,�Vp�x"O�Y�A��$n��9���W~s�!a�"O 
��G
c���4x��$�2��y"���O�ՁO�}�5�"�G��y�E�$6�����x���_��ya�>���	4��g�QA�B��y�
�]��p��& �ڐKAf�4�y"� �F]<Yz���q�P��-\�y��� 3���%�V��P��ϐ�y�!BY�l{��>^�uyOB��y�HT#1�$��/�pL��B�5�yB���d!���S1t�������y�!g��|Ia%� >Ԝe,���y��2W/��a���Au���t&��yb��6����;,
qz�I6�y!��N+���/�ʉ�$'���y2�K8c�P4xv�޾&7raT�V��y�l�fیQr�!�&J�\ )`�4�y���!z,�a�Z�7s�:1m��y2�ŁAa��0�OF f��pЭH��ybH�:*ڀ��7Κ�Y�(|�����y�e�+��������!2s	��y��[�!���2�pd�ɸ����y� 9&��j"iD�9U�D�1K=�yr"� `
e
c��{���k�!�yr�~>|m��� �d1�a�� �yk��a Ĺ�CJ�m"����5�yk݂rY̬�d&c��)��M��yBLN`������y�cr�J��yR�]�c�$!�&ʲR�h����y"DJW�x��Š�Q]q�s�%�y2.��N_�hd/P0}��T�b!P�y�@
H���qK��pX���y�oH�1�H�j�hBut�!QW����yb��!*����o�H$S�M��y��U�T�j�c͛o����K��yR#T�/����Ɯ'rem1$�F�y���g`�}����/ L"�J�;�y"��5 @  �   =   Ĵ���	��ZlctɅ<C���C���NNT�D��e�2Tx��ƕ	#��4"�V���$W�6�o"=L��@�▜i��w��/+5P4�A$�&p,jM�/N��M˥Ň2�N���"q��FR�r��']v�'��{u�D�	1,K�ɪ �U�s�>���VHy�#�� ���0dg$}�l�-~�qU�ΈQtb�����L�@���.7T8�'���p��:�ش(O��X1��1�N/��	*@֡���PS {#mS�Ǎ5��a�f*t�(F�<YB�|)�����>i(��K���#�'X,��1U)g<�9IG�>v�˓��h�Ň��ē|H��X�������4qj,���&1�B���!���~rC%5��@F�xR'^�Vv8q���`եn��9p)Z� P#2��pbg�0S�2b~�J0E�1c�T�B\�v@ʝP�=ŀ@�p0�����,H$�'�.��4�Ќ*��	�?��'8<
�.�]���;f_��s��-P�jxWi�r�pe�ɌP��]��)��'[��bo�o0�}�'�?)u�ϲV�  �@\��i�ӧ����e-O`�@��jP�08gY�T[U�'/ ��A���LX�B�zZ��(�O�*-j�iw�2]̓E����Sl�<�'����� �yRNq�hH!!n��!*���S�{.QiӊF�N-`����7Mݥ�?�d.>IE*6�m���R���B5-ڡy@t�qf%��`�A���^ʒ�O��s�b�S��'��9�� ^7�y�H̟;_�����s~��[��$I�5��Î�����If��9ph(x��e������<#�"<���;�D�n.����� �B�pH��a�aŴY�l��N��x����$ED� y�T�\�Pl��h*\H�Y� �$�jE#��z�	��o
��X���2#��Ֆ'�z'*խ��eǨ�&��k�7�l�d�W3G1~H�" �:b,M񔎜�D�D�O��;��*J�1O,���靦A�ؤ�!ÃuE
UB"d�H�hC�I�L�� �  ������3#�\ M��a��Ѐ$�B�^i!�$�(!_�T�2.�
$oL�BGY�\!�$D�C��,���
b$���1@Y!�$��A�� cV�QT�=�F 1G!�dL�I/�a�BoܪE���e�!�\�=�؃�U�8dp������!��E	0�2A��D��jS�[,[�!�\ >��6��&]J��A�!!�䇎]��0   k
    	  �)  �2  =9  �?  �E  ,L  �R  �W   Ĵ���	����ZvI�$��P����@_zX�B�׾S���A�A�8K��$�.?�����ɐ8���]]� �Ț�g'ʜj �A�a\6�0e�(�4�$�O�,z��1H� )�� ϷH]Ƅ�	O �
$�\[XP�a��P�?��0bS	B��f��ņ(�r�Y�( �x�;Рg����f˅Y
�TX�F�3W{�׋��0��;$�A$�t�.%	��]�?6�X�^�F�!�L��n�R����C��Pa�c�{����?6�y肤�7�H%���?q���?������D k��i0ǌOeEܘ��G�f�
�Չ�F�|X�$�y �,iW�[���T�27:�%�4)���%�N\�B�Cf&��F�(�fF��
X�B�AI�]7,�|�'�k�%q4*��yB-߱<���ȃ&�0�jY����X#��`$LOH-2���yx���xR�aO�����TQN���PJ�palX�Tg��a��4�ޓO:��u%?L8� K�U��Y'bѝ;Hl�	���O����O6�D	ﺳ���?q�O00�p�|_l�6�M&�HTcK�h��D�?S�2��#��pZjD(冒U�')��G�d� �jAi�e2��i�,ЋV�9�䎚���sť�޽��'�O�@�C�|����?���Y���-�(a���S���=i�!�d�B���+�Ѝ�6�)M�ay��	�o�\y3���6r�H��F�����P��6�|��[ ��7-�O���?�%��=���Sf�4�ZHj0�a���@�`�O��d�Of!!�L�>�v�ђ\Iv1Gg�"�\"��=(J�BC.�x�1��̝��Q�dK�=7�	C)K�h�ֵ9�
Pۺ�i�&���k参l ���o�-h�o��L� �O&��g�'J#|���S�w����?!<�,��BE{�<!v�ڲ2[*��"�v�"��W�GL�IP����&8?��C�"R�����<,��OJG}2c�k��6��O��$�|�wk��?��)����n\���X��߳r"���i�d�!f�� �xxۤ�J�+�5�Ш�~R����M1��k'��L�Xb�!VY�"F"A��Ȣ���n�u7�:}]�MT��(L��V>Ř&c�8g�B�k&Ζ�_P�M �Ğ���k��O��� ?%?e�I|?�D�$����u��FA����}�<���]nX%H��̘~>����Kz��?e�i>}����?=��� ��\�(��%�M����?�G�@b������?	���?�A��:�dşrW�K��̞h�>�p�Ő��~��'<|-���,)�C�f��)�ԪD�\8ܗ'�D���0�p�@<�*�s��̤���'S����w�az���7d޹�c$B<hS��ƕ�yr�R��`a����#Q���� ���M�g�i>e'�<kG�ׁ�&�zs膕 7�cU�6����B쟘�	����ɔ�u��'lB8�T �t�'�ޤH�ß�M�`-bWI��9w���;�O�-�Q�O ��S�S�j���:v!ӋXw���'p����~�<�s@=�֥k�/�wդ�X�"O���RA�-"���⍀���H��"O�;3E�;V�U�⍆���[r[� J�4��F��-1��?Q���TmJ8ya 5Ѫ(c�*�3!j��M��S%�?Q���?��O׏�?9�y�O������	
|����_4�p�Ê�䃭[Q?=`�=�� w��1S� x
ǭ<�q�0�	��������	!8|��/��w^���"O��������$eK앚e�HuYb�'4�A�"��@l90�*�i����$�'�B�a�'�2�'R�95�:a��؟�)@��1���#&�$�!���M{RB��?Ɍy*��O8��q!�#ix*,Æ�B2.(܌��'P������c�l�#���YI�M3W�ƽP[�m�	�<��$p�)�-'��svḣj'����.̡!⸬	�'�&��3�[�,hHUz�m@�N��]Ez"5�'I�j�x�*75"�	U.Vձ�i��'P&Q��8�R�'�'����5����Q�Х��غH��=�լě���+T��|��ÅA����w�K�D6ȑ �����q�|��X�_E��)f+6�t�D����D��Z�0=�P�7�����<߀u��I�`�<IVJ"`hP��G5:�"H0�@Zצ����4�j�O<��c	�p���A��P<a�8��Fh��0��Of�D�Od��������?Q�O#��a�jv��r��SL�h�6"T%Zq��
w�'6T+�'�\g��v"lu��e�_�0H�\�(�ɷxЎQ��-D�y$e��k�!�XŹ�'�l��`,KV0�u�!`U�: �e��'<��A	�U/>����A�`�OVPmN��?��ը�4�?)����,ơ	��yv�#Z�`�@�$=�Mۣ�
��?!���?!�HT��?��y�O�ވ��ƖJz�V�h�� ���д�Q?� :H�C��p4��
MUR\H��	�����UA�OfUz4�7}������!C��`�'�X��wJ�)�$*/=�H�@���ɷ��ũdiD86l�䭂�~���9�v���?Q����)�?)���d�O�����Fh�S㺐(�i��}���џd�<���'�ҵ	u�3\(T��f��C��k�s(v�Fx��)Ԉ��8c��s�`�g(��r8���2*�b4���B+�L��. J��00ǣW�{z����Cp| 1�'#�ջfC^:��Gzr�'�T��Ń�.Pv�H��J�o�����i�2�'��pI�C�����'���'�f�]�֘�`� q�(ڛfc�{�+	�UH�K B��	}�F�˳�E i�� �wAT� '�ʓ4�|݇�I;9������ú �i��f��˓I�v�I�0=��a+gkU���.��H�d��Q�<٣$�:@s�u���(H�\�SsfS榹���4���O�1����(�< ��G��y"b,�G�Q3q�Ip���Of�d�O8�$���������|r��C۟T �	MT�1�"��8@X����F���>�5@Kr?yfc�$]`�s�!rn�Eٖ�Ox�X����O�$�t�H+GKxD�S�ϟ^c��3��G�<���۹@
���6AIW����u�B�<���Ѱ}�q��UaT�,�`�c}Ral�R�O>(z��ئ��	ٟ\��:�R��ֆ��{H~�b��?�V�mZ5P$М�I͟���.R���y�S2��F*h=�$N��.��QGQO�'z�ۉ�iB�X\F� �_$7%�(ƨ՛H<ў���O�E��ቜ;w�I���� 	������y�H�\D=[��F�R ���%_(��>	И>�#��?l����n�3�v�)�é>!�'�x����'Z>A#�����K|=�%��\�P��c�R�҄�ٴ�����������DVdS< 3#	F�f�Ӆ�&�B!)�O?M	���%
.0Q�G�BOJ!�BD��@"� �Oj�%�"~���ܘ_>�Ń1`c�*�b�
��yre�a�$�)Bl�X�<�Q�ŏ�HO��D��A�-�B�	��8�Ĉ�̏�H86��O��d
�<�V�*� �OV��O����ߺ���֏S�v�6�ʠCD�jMR�Qe�P@y2Ύ�p>��˅�J�R`�I�[Ќ���xyd	�p>�vLֹ{���`�iɦ��ui���ly����?��'��Z���5�Ѱ��ءp��	�'I�tQ���?�A���ڣj�"E2�4QՑ��S�	�'M�Y1��Sr��gf�6(�@� �g|���	����	ݟ�2Xw���'��B���G,X	t$P<S�ȃ;c�R�Za/�&d6��D�.n��<���H����3���&eR�����/s��;R
�5}T�`(����V��!�����r�C��B�z5;Bh�'Z~n�Ot%;"�'�H��Ɓ'�	�M�<	�(D��ybjV�W�Ĺ0f�+\48Э%,O��<��X�c���
:B��s���D}��xӂ�O$�����-�Iޟ�'a�Q���lP9H �϶1*lڇ������x�I"����	y�S����K�pع��=[� {�+b�'ϰ�S��	
�G�x�C�d�,=��󓺂`������+�'_z.с�T�2C@	�$(���Q��]`Ҍ���υ+G�mQD�E�R�T����4��$����՚0(�_qz��se��M�I�%V��4�?i����i.a�����O����a_�n��h��d�q^rH��QȦ�s$�Z �д@#��9p�3b�� S�tE�ɄP̧d�$a�E�\��j���<�~�+��z�պq�B$Y��]����%A�����O��>��#�_�3���VDH�b�0I�B������O�'�"~J���Q�0(�$��,քt�Q W��y��	�05J�M�8$�@��+�HO��F��D��(F���&'"{%���r�A'Q7�6-�O`��S�s��O��D�O�$�ú����Ї�)E��P��21�����oT2B%[�(�q�n�3�ԁ8����O����Ao�I=e8�����#��Y���=�����L'k�J[2cT�ER@ҫ�|R�j�e��B.���~.�,���V1$��lQ.�Qyr�܂�?���'���v��p1�K��Ф�н��'h���Q�] .������gv���*x�tADz�O/�'��R��1-�Q��H؟h]��8�i>WM��"�'�b�'�v�������'@����J�� ��Hz�()%F`�~��#��<(�d����h��?a׉A����r&W�"����A��C�r9!u���3!
2�+�"�Xߴ��L�e�H;}2�'��L��2� �����а;����W��m/�����i���?�禩��A��Eq!�t�K�B�$X �/D���Rɂ*�5c˓/C�`�
�>�w�i��Q��K����O
�S�`ڼ1U�Q�gB.%��=�6���7�����O0�Daq&I ���j�@�;#ɍ"�ͧ2�L)�fڨ+����F��"�*G{bɀ�d�b,�U�Ϋ�>-�Q�4:�ʤ���)��	��"¯zMԭ�À�6�@QS�-Tl�H��-�I����}���L�
�D���F9A߀��r�V}r�'0�|��)҅M:n���jV)U8ubl�*
���M԰ړf�J(j�7�^�
�B�?,�t�A�i�r�'V�5>x�a�����Q`�b����h؇@FP\�W��M�2H�M����sΌ9���B-���!Xd/\+��O� �2O� �*�2�I�b���'�.$*n��$���	�h�<#��\B��B���3�·�U��Ӱ*��5B03���ϒ�<�j����\#8��Yc�)�rK XzΙBU��䟘݊X
�'# �
%EW7�Ѡ���
LY�}��'��#=ͧT�baZ�#�=[ظUH��VL�1�i���'�┺�dY63�'"�'��ß֘�I_��KW��7 �8r&�Ӊ^���%%H�(yc3�F%P�����|���/��O,�i�ᅡ���A�% � ��F$}���r��=�i{�+K�2��A���v�Z�R�7O`"��=��I��Nؐ�ҠawV� �&�On��鉅Q/h�cƎ5��1q�ȕ�f��B��	��M�7`E,����Q� A��4v	���F�	�]V�)�gŁN����� W�x��gV�Z�Iҟ������*[w2�'C�L�/�� @0f߉7���֍�9|F��'"	#7�HQ�W�z��1j���IV@�#���#S��I�j[�:e���Qf�9�����NN�L�m�R�7,8PN���6(���Q���'����L�^q	����6PhP��59bv��t"O��YU���PJIa"�mH�,�B"O2,�Ř9e�
�)C�c<�%�V�4��4��frJ0!�Y?��	Nr��	]�t삣*V�#L��5l��)�@��ʟ��I����ø8�|���|+��k�LԬ�����B25�6<~P�X�hO�AY�"�\�x󓇂D˄�#��x��h$G�hw�a�`ҟ&}Ե��@O�er�I�U .�	��~��'�q��,��	�uq��c� AR�b.O����
�\Zm�U Ȇy��!�F09a}�9?I�*���	��R$:�p1B(�F}b�@�;���'��]>�X� _���I<�4ó�N���CC��8�d�1شn(( ��c(�:ԁ�$g
��P?��|��.��f��T�6'˾'A�ys�:�?�D��]�PJfA����4���uw���\��I?53c+ڞ�\H�@C��'���EEΟ�A�'�������'��$��]�F�؃l�<�!i�'}R�!k
�Y�5��fe!����HOP�D�T@���"}����9i���1l�4E�*7��O��ҷS?��hu��OJ��O �D��|��V�I��@0�Wz�*�lS�y���w+�3�H(	� �E�荘��Pv���I/ ���h_�5��M��A�Sv�U����1	��Y���]�gf�4��|Zݴl����&Fx}2��a7LZ)Ox�u������d?Y���hO��I�ODu%G�H��3�����B�ɪ&�D}@I����VFI�6-BW���T�'�	w���k�N(�	�~*uR1���n����	˟��I㟨;_wq��'�IT��z��	^<�(3'�Q�� �e��73�Ѩ�B��">�qy%5��q�6h	��J0B�u�3!g�w-C�`}|`Y$��3m�p�`��M&�O� ��=���O�h��!�v�D���ۋj]��D��!E{��� z�B̡�ܱ/.Py�N��zC�I���U8ү֠
]�QY�G�S�J���'��I!I�,P������?%��L���	r�ٝc�R����s�ꠐc �O���OR835��&~a�F��!2%�|�I��%y��$s����Lx�'��l����\/^d��O�Oevp23����'�ָ �^��@������V�I6za�	�����}?���O$�̙D���/t4u�R��Fڋ�u}��'Y�� ��Kv�@�p󂛒C�.d��Zx��(b�*,+`�ME�l'��2{���oX<ub���?�����)��2����ObU����B:j19�� +Q��ȦQ���	�I:�����RI������):�ӘD���#�Rq��\*���	�GMPPQ���>:>*�iW�sr�9��HH�����B��3W��̓��X�\���⍳q��D|?1������d�>q'��
�Y{䩄�|�bq&�D~�<q��+l���h�5W�l�3'I�a�'��"jAG�]�L(�)X�e�P\bp�����'-� F�}������'R�'R�O?R��R:8:UI��m\��h�!�,�8c�`�zU�Fa�)��|��d.[��q�3/v�-!��0�t��i_�N��D�fI�E��5���z�4�i�H(�$���˦+G*�-�+!$Y	2�K���5�~r�'�ўd�S�? ��2	ܪ�68�G�U�]�"OD����YN���, -�l�뀵i�#=ͧ�?�,O�)0�i_�bO"8�5�B�]�@e0B
��%��]�%$�O~���OP��I������?9�OfH�*!h�?�����QI�B�c�Aϊ'�)G�I>C�����	%fhџ܁$��.ٚ�h��]��=Ҧo�!�lX�����/^2UY"�;Z�V�o��E�֢%�~��;M��H� 	N�d�<�A@��T7&ړ��O��p$O4c��Y��B��2(AP�"O��� �B=V��� !�t%�i%\�L��4�?�/OA�dLK�D�'��I����AJv���g�&�S��"���IU�N���'*B�_)E����e+^;��#v&Q�
T��ӌv��$Z�b�+�h�"҇���=��%5�i@"B.l���(b��u���!�݈�A݊"ϒ$����Kv|�S�T��'<����d�}�1�m�>��`�B�"M��s��F}��'y�t���	��X!d�2l.����'�ɼR���㜝�p�cIX�<��=���	���?I��򉊀`o���Odđ�D�`��(��Q���5g�¦I���)K|x�"h�7ئ�R�Å4��)6�3)�l��A ��7q>��7O�%Am�	(+p�d��l���&��l��%�XWa`�	�:�N�5��1~��1�'��	-T��?��������>y����o�RD���Y�m���+Ji�<�$@�=b���۳l� i��c��@�'b�#�w�
�c5,�X�č%�2D�'E��}��F�'��ň3.LА۰�'���'K�O���#g%���`�7��r2�5p� �s��Ҵ 
2�р�;7L��3E��|Z���V�>�ҍ1%��F�h�f�|�e��� SwA�����|�W&�=� @��OC�_�s���Ёd�	f�d�cP�4
�'Z2�	y?9���$s����'BR�����`�T�<��<c�ش�HX�n�NM��Ϧ�{��4�����<Y 擮�6�Еn��������>`����?9��?i�4�n�O.�k>�8��̖z�=�Y*FeL��g#6JHš�l��97zWdM%HWDbW.m�:\�6jѫ�%�Q	�!a�+�6f�5 �M�*X%Z�����MK5��<aV��=!S�Ox��䈖���L�3�ͽ[Sx��(�즕D{"�I�Z��pz7E�n!���E;f��C�ɪ.��9	%�Y�B�!��Ä5E���1�6�'!�	�k�d�������?H&d��lCC#�Y-����n���A��OH���O��`��.$�X��"J�� �p�[�|�1�
�k�h��aAx��"��V�'��Y�,�$��%|^��	�#)���3"C|<sF�#41��xb&�:Z|�"C�+.qOj��?9��4*B.~8�DY�9����f�_���*�OB��C�<H�R�K7A�Z��%�'}��,��c��bfP4ۖ�ҏc]fA�'BR颡�y�8���O��'jHp����?�Q�I4E����3�.1c4`B�U�7�C7_���i���_���Q����[Q�г�O�1�4�	f��,��4[�Һ���F�O�q�͉��da�ͧ,kL�5�5ޜ�r��'!��ʧ��)��(��AS�/��!$^��p��Ɵ��R��O$�"~rs�=K�ޡY��ιo�ёG���y�jJ>fs`��q�H�xD�Ѕ��'���8��|��L.1�(�n
��(,����!7.�6�'��"�% *$H��'0R�'=bm{ݑ�i���R�YG�)�g�څa*���E��A9�B�L�~Yha�tT����|�T� ky�Oj-��&\�h���j�kQ�;v�Q�X� ��I��>�� A��7S�?R��*מx���n�¤y�Q&*�p�A���A�F�B�$LO�R�� ���{�m��?)d�F"OfQ ��G�#�(�0g��,ѣ��in#=�'��C��p������VVw���0A˂i���3��?���?y���Z���O��ӕg�,lȥU�`�s�Á^���R�@�bM� Yt�Z�M����6HD��� P5�ɑbOB )wK�8�N���H;� g&\a7��  H%{,@̨��)Gf*1h��ɂTY��D�!i��)��L�@*�%��� �
x��=zXP�m�0Rˌ�E<"߮%�ȓo�,@(���35�\��(߂>E���'�`6�)�d�-c����O��֟�,��L�)>-kT��#�`ŁB�i�>(0��'�b�'@ȱj�Cs����N^�!v,	+w>��$iƍ,C�u��	Ѭ|~�[Em8�H�����%N=X���-[h���z�O ���v�B5<��{#� ����%4�S#���Iǟ��}:�'4�nusf!��<��bLY}"�'��|��9�|E�`�_9Q�)`�됡��>�7����VhЗ��� ��!v�%����>1#�а-��v�'��Z>5�㡈ޟ��I�Am�l����	����D.��t�viZݴ%K4ܩ�g�<O���J�i�&e�>HPAW?��|���R1"�=p�	=(Zq�Y^~��Ʌ]�@����
�f96�$'�H�D�DDחU6��[�y�ˉd��4[C�'R0�����?�O�O���ON�Be֦#��=aeJ+T%���"O� ���M� t�[ף%�~\{��	��ȟ��02�N�F��l�ŧp9��*į��Q��ޟt�!�<�����؟��IßP[]w<�&�
�h�S@��6&��`Y��46�A l!?Ֆ��-�UR����Ƕ|:���v<�9��"NZ�3G�3�t�െ�3p�lR!"X�
�h:�\>q���)�Is��+�k�P�����-O8�	��'�2�'��O����2l<�S�`\ m����ɱzg:C�I�)��� ��qE��yB(��&��7-H}���4�'^��6x[L�R���p�ޤigC��-ޒT�G������֟��Iџ@P^w��'��)�ct�ͨ��Ъ�D�W��b[�Df`�@�T-�BC�I[��բǟQr�x���A�T�����������h�3,w
�I����;��@ %�C��P� ���M�W7 1��_j��X`��>�^���kYm�)
	�'��Q)P,��H�=rE�I1NF�P�'�����Ó�x�(E�Y?JK�X�O"�oI�	=�&q�4�?9����ۡ/�`�`2��H�J�D*�4�M�c)M��?����?$ ��6Tz�b��?���r�Y�Ui p{�����܊f�Q"\��X�甈6� tEy��O(�\��d;ףƕ�D���S�>�"�ձ-!�(�d�4���w.>�~��������[�M޲[6r�!30[��e"Ofܸ�">���d%A-��9x��'� �G��t��&Y	Vߺ�3biS<{ц��'���A5l|�"���O~ʧ+rM����?��)7[�t��ቚD��IXd���@�f*Q�^<�2a.�2 ��f�T�BQ����.4�1���s4��0�SťUch��l�O�RC#E3��!b�K�W��Uҧ*���0"ƥ[�?��'C�rUB �D�X���ez� ���7R��I=��S�Oh*1��씭.�L� �Ȕ?+�:�"O�٨�	$VypU;BYE �I��D�O�YDz�O��D���n��5��xM����!i����O� �?7�&�D�O����O读I�dAf`ь/'�0��d��<�M;��,tX��d�Qj����$A>	cTi�a�>5����	F��,�@�.*U:Pɔ�
�Z]'X>�<!�F��kŒ���΀�/�^�vJ�٦��	�68����=�M�bW>��?A�'v$�3�ȝ|U���+�y&D�J<��J����.>l ��2vW60mZ�M�G�i�'���O��I7W�@q��5vu�a��<]� �զ��E��X��ܟ��	Ɵ�Zw���'��)��x��02KQAj��	+�D٥�3a�`�C�ٍ�@ٳ��mb�b����3`�`�вd��ۄ@S�����Kc嘳��'�t�z҃,/� DB �U��(OR��C�'6R`��� G��^�c�J�s.?D���ciZ�h�8�"�g^�T�xL�`�;D�4B%�F=e2�Hb4�O�q�n��`�>i�ib�'�L�4�q�����Oj�S7l��[�ʏ �ə��@�@�
6�������O2�ĖY���D)�?!31)�'��)9S��!]@��"!�'���G����=5�[�Q=[�Hy��Nɢ�hOpc�'k�#|j'D�(L�{��K$T���WO|�<9�EI>��!�R�R�FQ�q;�ύxX���OV�UW.jl.%�C���G]6;�_�Pbq-A*$�9밭Щ_k�ի�/?ғ<;=�7,ۓB:�I�`�71j��ȓd��0�͌;J�z�Vʁ�Me�P�ȓU�8i�ס�
��c�]0O�$���D����(}k�M@fM�%�j��b�D �iקf|j��D-Y�jt�,��rX��
��JZ6�@(�f�J���ʓJ��Ya�b�)��x�<C�I ~
,���0� ����^�C�I�5�BI[@�B���#�~t�C�	�xX���_$l	� 6Ez�C䉚F�-���� ������Qq�hB�	�d�2�І�V67��+u��f*C�	�T�AR�p �z��B5~i�B��)oa�!��LN�-T��C �c�B�	�r��AkУ(����&n�|C䉱,h�%pU��i�e3G �IDC�7F�mK�(V� 
��9c�B-��C�	�$���Q9o�$<jRH�"n|ZB�ɾ �ƀ1Fϝ�Ͼ�{�G�V�>B�I/��T��hG�B�����cU6��C䉪T,�բ̊%| ���02E�C�	wΌ���
��R�u��B�)� �0zfB��;Ybs� ҡ��(1"O�p2do^�\��S��ծ+��C�"O6Ac�B�0���1�H� rV$��"O�8� �V�R ��(����OR�1��"O6�8�JN7 �t��f�SwBTxS&"O�h�Ck�%#ޥ
�LD�T���Z�"O��Ol<F2R� #=��g"O�L����&}�y1�*�b�%y�"O�H��n�$}�0 ](Ck�C!�ϟx��wI="���a��05!��J6��x�	�}��X8�`��B�i�c)^*hC�eSG	G���p3�*D��t�î,Kƃ;E(�%G�=&!��C	*�I�9N�85j6$�7`|!��F:� J�oB�j��	�*I|d!��Ӌp��p�'#s���!ʒ�*�!�pD����h��7ƚ�p�!�d�.B��S�G�?u �����!�'&֔��Ƨ�3l�ʭ�$EI(5%!�2iF��ef�
Y�.��%.S"!�$M�I����1�g(l	n��:!�[�.Φœ�UQ��B�D�{!�Lk�=Ā�\�6ɢ���y|!�d��3��]3��GLv����Z \t!�Ă�����C� �c�V�Sp�*u]!�DT������=T�atH��!�4c�:�(d��/>�Rm�D�P�!��2�T�{���6����I+m<!�dP�RD���OT�C���rl� %*!�D���{�H�}��Y���2
!��ٰN�� v��6km�e��? |!�D�gj�J4ƛ�B^�����ɬYV!�H�{��yQ���vKx��#�*�!�D�~#��ÄI�Vd���LO@!�$E�;�ʸ��
y<!w�B��!�N>v�	�'�Xq�n�j�˛��!��Ȥ4b.с��Y�0��y�&�6\�!�����pÊ�7�:�fNX#�!�D_G�,�s��r����1��X�!�d��%�]IDA�#�(��W��_�!�ڦ2�@��@�e��X&��_K!�	�EeI���"'8�A��
�~K!��5"��zև�v浡À�	�!�)��s3eT(|Im�<2�!�M�^<nT��"N$=_&t2�L�-3!��>���:�"@�@QM�ぇ�aI!�G�q� Ϡ�����ʙF@!���"V��3���L�����A�!���
v�Xa�ي��a��V�F�!��\q���BW�����׌W��!��)}K���&.E��h�e�P�|.!�D�4)���ѕ��<D���C7��M!��9L���R�y�na� �3C}!�D''�Eh�*��(3P�B��)Gu!�Ă��&,3�'H,@2������hn!�SxTX�̑�!�@�kdfۆd�!����2C�C]���P�!��#h�Z���|����wi�B'!�$ޓjxb&��^�q!��!��0a��Ep���L��e2#OV�!�d:#��R��pW4�Ҁ���!�W�_����VD~Y2$�ʙ�{�!�d	2e��4�gTY��d TʎO!�dO�L�kAn�_��ɂ��R�!�!�� v�b�g���G��@��DBB"O���	�(����7��5bS"Ob��2O4���b�cБ �Nc0"O��C��\0&�lQ��w�R�ѓ"O@01��m�Ta���I��"O��"J��D�Aʩ^ �#A"O�[�5$5�h ���j#�t�Q"O�}Ʌ�K7M�!�`����9J�"On�Yt/T�Aj��63�Ȭ s"Ocà�(2Ђ�ˆG"i�B�KU"O�L���[�~�h���5ܑa3"O*�f+I�ഢ��p���"O�@�'�4\9q�F�J*T��"OZ�$b��W.2�D뇏qt@�v"O�8	�Y�%0b�k!�1a����"O����	UD��a�&G!h�"�A�"O �Q����Q;ZP@�dA&Gؔ���"O�`#���%�"�{%�$����g"On�� ̚<Sg��p��ڼJg�U�p"O���ŃL�ԙ!rB@?_�zT��"O"E"7��*RȔ����1�b�AF"O�����D�0T Ū�C��ye"O�8�a�����;0ʋxB�u�D"O0 ����&D���hV�%Ұ"O�+�O$2tB)����B56tr1"O4�:�Ձ|>� V��w4�k7"O�x&���+�JY���O  
�h�"OX�B� s��y�c�B�b)�E�"OD�{��U���u;� �?*:� ��"OnC��� gdA�RG�r���D"Oj�� �	n��ѦF��z����C"OF��n�:Q���(���A�rh�"On!�'ȒJf0�(�c6v�L�"O,9���231�"�Ŕ>M `��"O>�pB,�1n��!$�{J�P�"O�����=�&�YU��M@�0��"O�e�)"�rQY�
\!L��y��"OFdo1Ia�0@��ZD�yj'"O�mcSO�#V$R�.�~D��"O<1�2/�+p$��r�����Ģs"OFQaӏ� Mjvp�w�P�8Y�U8�"OΙ`�@.0�.,w� >��T�"O�i�i]=\���+�o��h�h1"O��1f�"�{�O��H�"Ohd�g�� zP
u6�˗"O���k�T|�bQ#ߐ ��"O�)�����Z#��0�J�f����*OBA����&ʊ9���$����'��y���N�6�e�G��<| �#�'� �ँ� ��;�bh�'�V�0�H)t�Ƶ�aT�g�T��	�'�v5P텧��p��Wt��t�
�'b͛����1�*�C����|�~�C
�'u�T9T�U�F��J1��&��1
�'�
eC�.,����nޕ���#
�'�^<�%�Q�Xr�d�hTd(*�'��-)���1�e*иT:�5��'�f�pT���j���¸�:ip�'��9����x���I��X���'��a���Q����A�@EI��'њ�x�ΟC��(�b�w����'��Sͥ"^��\�g�&E��'�t���l��l�����G��c���'�n	�����n�i&�іH����	��� �$�`�� >!���CA�U��E�e"Oܨr��@�#����"��9�V�"O�a�$ �4P�$�r�a�.����"O@� gV�3�I�S@��l$���C"O�܁�`�6����2��W���+�"O� r� ��;6`ѓ��+���"O̕XM���e��E��:�:"O�\�G�[785����� }��!!t"OT�0��@�`)b�yr�Ӯ2N�Pb"O�a� g��ؑ�m�J'r1R�"O&]:a#Ʊ*X���㎜���}(�"OP��CMڧ,z؈�6mO^��#"O��E�[�Y��D���kE�Ds�"O����@�+���Q
]��*]!�ȍ(�X�Fos���5l��!�d��nR~�9���/m{�ma�#�\�!�d�)F-���"n�zb�9����+�!��ׇm��EM�F��2��	*(6!�<Y�p�jL1i��8��i��w*!�$�*N8�I�DG�>#�A[��Z�{�!�D\��
MA4f� %~0�Ȑl�!��߬m}��l�������Z�!�d*@�EȆ��"B	Hԙ`�PL�!�Մ3n6��b������!�D�yw6%	�`I.|��̀ֈ��B3!�R��dQjGޱ� �(�51!�$�@��D�۪e����ϛ� !�\���Ԛ��= 8F���d�#1W!�$�:s�\���ݞ,�X%[`D�[!�Č�3�|}��C�	��EDK�7!�՗9��@�W�ԙ?�ΤAC��+{!�$�<%��K��'��h���ʁS!���%���[���ACo�q�!��T�jb�#� ��;�ձ��"9�!�$��"�c�\(:��a�fԚ#�!�Ĉ�
�.��C�8u&��z̂��!�dX�&��`��_x J��Go!���4K��b��F@� I,n!�D�N�zԨ+�x]�-�0T!�DL�%��%���*Y�z�!��Z*���!'U�)g�cʏ&V!�Ϝ_�D	��ߑaf��`" �!�N�gg> �p�0FhAh�	�g!�dB� ���Z����	�(\0��^b!�DCm���R@ �x�P03���`!��akZ�Y!�.y�>��˫Nc��)_�����/0�uQ�Ơm\"=��M�n��,W26��x׮�P�<9�n��/8��w�5�lh��p�<�)�5��Rpi�4x��\P� X�<�q�
�P@�LǪ�U�^ep���R�<I�d��p�H�Rfc��^q` �P�<� e�`�ڝb����`��
�K�<��B�M�%��!8���[F�F�<�%�����zt`�}8��+�B�I�<Qsn�
ps.�z�/Ǿs��9��mW�<��g������64�6(����b�<٢�F<y�Qq��
�%-�e�	v�<�`.���Yb�*���+m�#H!���L��-A�-X�����\0,!�d��dH����ˮ""�钇�#�!�D�%R�h*�(��	�����@I!�d
Z����B�q�|�DP�'f!��s��20��a�<����B"O�d*h�"������(>���"O� RAh2BJ��Ŋ�M>.	��Y�"O�q10O�F\T�aMڸ���z�"OJ嫐!�L����.��A���B"Ol���&L�"��01-�!@4~�!�"O����ש	}&�ZEF�%4lP��"OF!�2+A"��qz��Iέ�p"Oz�����Y�:=	����"O	�B&/-"r����@H���YA"Oz�8e�$L�!3E&[
l��3�"O,�C`-�z8P	�I�y�"O.�� ��m��4�ܺ%�(]�v"ON�0`�X�i��RbǘX�mp3"O�=ٗIP6���&a��`�a(�"Of9A�Hٽ �J�Hq-Ċ%� ��"O�E�vj^2[�FX`�A<o����"O�5��.Q)PE��/���4́"O��b��[�~��&��3��I@Q"O��	�	���I{7L�&�He�"O.��q�ʇr"ع�-�0v�h�@�"O����մ�$!"�A��`����"Of$b�ذZm�1b0F�{�ܭa�"O����W&941�&�K�i����"O�x�(��m�0� ��H�>���"O&�P�:8�aj��"xR���"Ov��D ��"����Jr�� "O����!W�M<d��L��U�W"Of�ꋆ��=�,	5
N�RG"O@yF�+���j�3C@]"OVP�`)݉O��ը��0��@"Ot �Đ3K8�CE�&~e�"O�@v�H	=!:�#f˙�ciP�2"O��W/1��{aj�0���Ka"O
,�f�Q9e���p�f��.�s"O��b�X�y��*e�>
)Z"O*M�q���b�� k	�,�*5��"O*�֊�(7H��'W�1�Nl�f"O���L�/y��ӣe�;�\��"O�<@gѬ]"A�wD:�ܜ��"Or�d	3`������`���"O�aY�V�GM΍+G �H���"OR��T�Z�2m
NA�ff��C�"O2�I֨&'�p��F�y^L�C�"O�Y��ĶM���L�1h/��u"O�$���^�(p;w
U5��QV"OlU�S��.���)�_�~-�"O��iD�S���0 �A��u1"O��"���~��pi��^,5��u��"O�hY��P:OT9�V$�;a\Y��"O�̉�f�a�z� V̻+u"4��"O ҧ�P�	 �}Z���#\q|1�a"O�R�F�TL���p�3bR��Js"O�=�"�
oސ	���O�٩�"Oڀ
���\pPdP��H�'��"O�ɃREۂ^�^4�#�7$yT�چ"O̙�X?<����`���vs�Q�V"O8� ��N�S��p�U�E>D 0�E"OZ�*�((��L �dE%4)�U�"O$��`�ݑ*��� ���OR4c��䚗�(O�Oͤu�@���s �8@���m���'V����Ţ=����V-�d�><a�剆�H��	�5��eˁm�4^�z� �N�� t�C�ɕZ���@�������0N�C�	8-qd�z���.I¥Z�8�C��\��	�m��y̕8�)iq�C�)� �$�R��l�v$�����}���4"Ox�va������_�p���"Of,�$$S"2����M�j��:�"O���3��+���7$ȵe�(�+"OF�x�*�xޞу�"��7j��"Oİ��/A� �H(�?O���"O��{$�я��a2 �(/��"OF�sW"F=H�5�D�D陇"Oڼ �j�?�
�bݜL-�L�"O0��'	6v���Wlݵu��$"O�L��F1R�5�Pn�Q�X��"O2i	Uc�N$!9��G,b|��"O
]x�Ϗ=�
�iw!N$y��e"Om�I�i���Kea�?m����"O���fI����`�G	�bV"OP�� �{����w��B���"Ol�+�7�^�
 ,O7V�<k�"O���W#{x��Q'*C�'A��"O�u��.��|�S��Y>C n	�"Opi� ����hN�'�ƕ�$"O(��$��8H�t�U��ڄurD"O쐡�D
=��9��B(��|�"O�x�5Eez�X��.	D)�"Oڵ�w�����p�᫖8<�T���"O.\A�H>�:�C���Ht-�!��#V���e�
qa�}����n_!�i�!0�OҼ0A�|�5 @.&����I��O�!� X�S��r�%c��\�"O����N."L��q*MB��`�C��*����"�Ɯ1o��ہ΍�;F��{"OR�xf�2NP�(
���K'@л����O
�}���D�4��0:00=[���Q�0�ȓ�`�i⠇�E�������2Y���{�h��D�<�xt!O�J�t��gI�B�|���	e"����>���^h�"��nxz��D@�<	�e�0W�J�7�O]�DzrCCq�F"���F0��eh�
��:@@@v�M� V�۔"O�=q������l�t� U�)�a�i�<#=E�ܴ5nYF�,&ߘ%Qf��2q╆ȓ�,$�$O������;��8��v���0��ٚ9�\H��K���ȓ��M3���+���`�G�9ꨅ�u&�+�Z�d��X��M��jK$��>AeE1�S�u����.N)B��[D�Ǭ!x�C�,n+(�@U���M܁sp� )"e3�"9�I�H��	�^���U;��@BK�.�B��5E}P��W�3e����gN� M�
6�C��M�	�`�Ѝ[�DS^��<9�HԮ�`9��I����Nv��XwaU�.,J���3�!�d!y2����9n'L�D�C� l!�%�bm+Ţs��0B�>7:!�Ο}G2��T�ۃMr�B�G*<�!�� j��)�C�2D���$c��u�!���r�xѲN��Z�����`l!�G,6��H��,,��� ��?Z!�A�����e�a^�����5R;!򄗯y�^�날˲�H�yT�$X!�D�?f|Š��R58Xuf�Mh�!��.]�v,�Ueɔ��p�O�:E�!�� �'�9��i�!sN�y�����!���(��/�1x֎�(��"O��g*��C��G-\�d��U��"O�}x�&Y'�b5)Ů(bL!s$"O>FI��Ɲ��
%j
,� �"O� ��z�/Z���A3W
�'A	��R"O�U�É� �8��iZ�gTM�B"Or1k��V�YH3�B�n}N4c�"O�AХ�#w*�A%�̌ p�0i�"O|\S*�	+�	3��1-Aޱ�"Oʩz��A�$Kb���ȟ!*R}��"O�!��lA!m ةfR(~�[�"O�т"F�3v�#S�߈/���G"OR�R@'�"n!����DP�-r���"Obt�%YhBġ$
�qٳ"O�"��<K�JMp�������"O@���=v0�' ��@�p�"O���׭��%φ����9"2��"O"��ф'L��+�nσ!<ĩ�"O�5�H�QXD����]2X�ݺ2"OȠ�5Cņ%Y4�zf���L���P"O���΍\B�����8�rx�6"O0�ӴA[�r����[�u��d{"Oi	�,|p��逹g��0"O*c�O5ʉI�A��/�0`�"O��	!�R�^�H� 
%|��A"O"S���C� ���+k.0�"O�Ě�C֩i�b��w�",�f���"O���HU�A0�usb3|�8Y�"OheA�G��G�lep'f�:���w"O@���E�MY"�8�$��#��5ɒ"O���Q^��U�c�aV���"O�Z�+E�{Qn��v�ĭGj6}��"O�8Ԏϰ���BBվ^�
�"OV,�Dk��#Ā��@��b�5"O6Y�޷��	S���EM���k1�s�·[,�;c��$��ȓ<hҵ�8��1� D�\����ȓY3N�Z��L	~ ����� ���uK����ԂSm��혂~\�Q�ȓH���	a� t���㑀 ��хȓ3��E� ��Ҡ�"S,&���T,��"��A�6�@h��4�����XU�]�H�0�H��a���:�ȓ8:P���V�8���� jת�ȓg�x�A�K�F"ܬrC����,�ȓ	<d9��6���h�C_�9g���t�Ԡcv��
yƼ���J	*8��ȓq�L�񗭒�<�(ԦG"T��ȓWiH!4��1K�<�M�B]N ��xI���� �39� $8'�-}2�(��]�\���,.��x�I&u�
��7SP��#�`�>�[��M�2���ȓ%hؤ��,�IҀ����(���j��t��K,{�����i��D��SH�� @�?   =   Ĵ���	��Z�3t�G�4=���C���NNT�D��e�2Tx��ƕ	#��4"�V���d��6�oZ<}�F`s�Q�9�)���Dp|Z�x��>c�G�@:�M����*��n�
7���3V ]#3-
��	(J�"� �-
�Is��*�Ś��ªj9V�j�\��ɱ��)=��@M��`�Eێ>�T=Ɂ��)� x�͋�z� %�n.��I�a�!�4_:Af�ʓG��a;�}��Q�'�\9qD��(�~����,|i�Ds�˘�Y@�s"K���d�'xh�U�Il��V	 �өO 1"��
U�B%!\���i9p��(K)O�mq�#�#J��O���2=j��5I�P�S���$S�r`�gՠK �	�GԢ��GQ|�I=g��5�"Ob�S�T�t|�Dj�l��Ь�(N8��;ӡȡ?�t�O���'��m�~��Oj=	�)ۈ,�L�� OT:3&���aҮ=" :�Q埄��E<�)У�����'v�p[孍F
��:���橔�vɎj�J	! ��Sa�'��t���Xa}��LΟx��O�3J�
!�d7����8Mm�1!�T �n��$C�� ���Q�<���O�`r��LyR���  $o�43)Z3���)��O$_�\q���ݴb��7�Y�<� �<���Sڇ�Չj�-x�'�>7��M�8E(�`��Obd�!�%�� *�E 5v|���y�v�d)�*h��4�yB��O� �&`�$����ęi��ݘwH�	�N>�#%���m&����'�M���	�i`!"���g�1	ƭD�}��˓,��� 7�$ʓ��O~H��i>�,���5+���f�O��i���ž��a;TW ���ԛ�/���8?�:5Jԍ�:�XI�aQ��b�C��@$C<�3(��W0=���97��ر����2���?P�V�1ҭ�4y���t��<�S��X�ԭ'�|`"���P��O�3K
.eq0��"7Mo]h7� �2aR��Ɩ|��Uzr�R�y2/	j�ъ M�<:̲�$��wk��3e"O�0��
�  ��k�cl���A�	J��b"O������������+�8$����"O8��$�Б%��!��x �Ѵ"O��!���9X���
�6��j"O���C��=��	��Q�DC�"O�a�4C9Pd��Z�[}�P�"O�@*%�I)dy�@�V��F���r""O�%#d@T�X@Ab#=�}��"Op	���&���0��ˡw�M��"O���sh� AAUm�� �G��A�<a`%��.�2�f�d���b@��V�<AA���z����A�=Pt�]M�<	Q� # :  �   "   Ĵ���	��Z��w)Ė;"���C���NNT�D��e�2Tx��ƕ	#��4"�V���d6�m"	��u�@ǃ.	M8��b�0J`iЂ*ۯ+p8l𤃢�M+����Z��W�>��;Eئl���'5��#F)�2�d��2�ǝe����H��9c�QGy��0t�|׆,}�]�y�VtB$�R'���
Ĳte��.L��(�' >#C�Ȩ� H+O����K��0l�S����V0Y>���i&��"����EǦ�MD˓�H�#H^O�I�+~�����\�� D
9�J��(V�8s�O��J�G�q,�OPQ�En�;t^��lZ% � 1	���e��>if��kU�� ��?�;O>����Kpf��?Q@S�х`/@"�@V�O�����J 9	�F)�b�d��BnJ����B�	�[���B�@�=�4%�RM]�/V.��P�A�'p,������	%\h���ay��{W����Cߎ ��S��?��	{.t��8���@\ќ�{�O���'����/�~ �t�.���Qg��$'��r��<�����$�@âb���6�mhp���Jz���&�B�&Nm�(�Ō���?���R�>]`��7R��^]�>t�C��&�bA�u���RQJ�)�C�8����-ErO?P(,m�<���'��mQ�Һs[���w��*�P%��~��'��шâ?�(�O:!�P	G3��-%*��H'�/E$��WK�?;��ɤ,BTi�剪6&�'X��b�d��dk� V>ڙ��'t�0Gxr��a��~"!F�yBy;.�5%�T��f����M+m�n�څ�F�T�GT��tKA�7��ʧT����B���o9"��P���q<��d�\���,E2�s!�QV�#L)�2��9��Q�7C!A[��"�X��ƵJ�i�p+�'�Ī�i���'�Zy��h�iq�Yx�˹.S�H�\��c�"O
`�p�  �  �� 2  � �Eƀ+���ȓ/�:pBҌU�";2�Ջ�
����'S�63��^���D�Oj��?)���5O�����E;p2�rucl��[���O���ON�(�)�O�c��S�f	Խ���A���4C��7:¢=1�"T[�O� 1Z���*�,�����P>
ۊ��?@�"b'�'((��6ѯ8����>puF�ȓe<@cOM16�dk#�Hjt4   
  �  E  )  .4  �<  >C  �I  �O   V  �\  a   Ĵ���	����Zv)���P��@_zX�B��S���A��
�8K��$�.?�����ɐ8��2��]gZ=�	^�4�tM��g�:d[D����ܡ�2�`q*?�Op���ΘqݎPp��w_<)a#F]���a�̊�Nn�)�7D�H$Jdp��J`���H%�cwl�!]"jr��Q����dɍ/�L�A�+Ո!ȱ��IRx����H�jɸb�}�Z�A�l�:� 	@)��=:�Qy�O�M*�ST��1�����z�|��3{(�L
��>�����꟠������[w�bj�JT�صN&}q�(�h^.\ Њ0��k�Y�ԡ��)�$5���o�-��:r��O�� EZ;^�* 95�S$y�2<"��PxXbe��U�>U�%���k���;;�ݺ�S�$�Jm�n�
��Vʃ�m[����&K���ė'y�m���x����#�d�OB�$����!e�Zm
���!>�L�kc�>Q��?QL>E���&8,�a�>CX��G��M;G�iH7�?��������<����P\�y�!֪!K����LBGR�l��E��?����?��?�ݟ���#�)8�僻%I�Q��'zڴ	�U� �c�G���S��'�����+��ڃ��/L�c�K'V2�m2�N1�`��!B�O`���Ig�����&X\n}J�͢s@t{d�cS��m��M[�����O��\��SO&�3�*�5U:m �N�"o>Y�ڴ�?��F^�!# "U�E�k��6	�'d�7�Y����'R�r��'�r�'��	N^�ɚ%�/n�XH���oP�dŊ[�b�'���:$��ԟH��J�:zP�3�ƜH����Ɋ%�̢~b �΍9���#Nܬ&�V�[��IX�'f���f�>m"����`�0��� \1,��M>D�H���	���Z��B{f$���I2�O2��'T���1"P	~�T,���xɫO�#f��O��D�O�˧�`����?��^�W+���kcIKáR�77@��ڴ_l�����������}�9�� �_N�|�p#ա x�c���O?�Go�q�t���Y�t�� �Ԋ֟l8��O��$�"~���YO�.U��SV$����E��y��3/l����Y$��S'�-�HO�D�T�̛o\��0Ƈ��uTna��[�t��7��O|�$
�	�\����O����O���������@O�^kl��0gB�|s��r6��SyR�·�p>���4-���7y�
 �P�uy2��%�p>���V&���:���+h�c�ʗoyRj@,�?�#�'�1���3B�@��v�בD��'P49AsnN�'� ��ʍ�uwܨX޴X����N�ɇtCdAC��@��v`TZi׊� K���	�`���HK^w%b�'8�ɔ0t�B��`-K@��8 ����F$�l��D�?8���,�Ե@'H�8t�jȲVĚ ��}"D� �?�v�г1(Z�� �週�p�A)�!�DņK��qZ�˄L�$���22!�d[�-3b�YS�
����A�Yw�	%�M{H>����?)��?��Ov��x�&J4"�V¾k栠VlӢ�DE�O����O
�� ��OVb��ӝ>=@����qL�� O�?v=A�!BV�O�页�x��aƪ��p �a���F�A|�i<�'f��s���q�>� �B�o���/��i)AO�zZ�-H�"�-�����dա^�K�bݲoʹH�B������b2�E��ԟh�	U�4�@�kS��'w2�`Uj3\]՘�/���`9;�-r�j1E-�O�c��g�;��(�'�	%o2���Q��(��I�I#O.T"<E���Q�CfN��`�5o�vh`�
5T�fĽ�?���|����x��m�KO�r�05�v�
�gSB�61��f�:>��bC�=OL#=����k�p��� �v�����'���ٴ�?���fۄ��?���?1��������,V�Hl��$�8���'.�Dy����p>i���m�v0���s�6���Yy$�p>q�jM�?8�ڐ�H>a���L\yR�C�?A6�'\���/tVEX`�F��t3
�'�t ri�Z�q��Ѱ7ǂ�4}����S�7Z��b�S6��I�h�l�벎ߧzI0a��̟�������Yw���'��I!H"�F�O�$���T7�r�s�j�,Yp�����=�D b�ճ��л_=`<��)�?B �}���?�?a�/�o}B\JD��"v5t�B3/� �!�$С%)���g��t#��0��W��!�Ğ9H��{ W,Z8��tb˽Q��	�M�M>�P��&7����'�ޟ��h�)J�	S�Aہ,�H%�EIB�i��"��'1�'Y��R�'1O�)�?��Qr�ݑ8����֎ܳIў8�`@#�g�? bE��(O�q�ލHCh�D� �퉆Z�.�d�j�Ol��Ӧ��o�(�)Z���j�'�P�°a�6N"��p��<D�%��^��I�[������\R!�$��.�����?9����@34/����O�(��
Uָ�3Z,�E)qG���]{S��ßp�<���':�j, -@Q��f�+��OԹ�A�)�V�X���	�L��s��M�D���h��3���I���S�O` L��nY�D\ ��'�[Z}x"Ov�� ��pi�!aܬb��鉈�ȟ6 qL�\����UhE�N<@ɛ��Ԧm�I�@�e	������ڟ��	����_w6Zc��s�#�-3��P�I�m�]`/O�py4�'�Z�௛� n�Ҁ�!_,�ei)O��f�'T�Q�f���O���8@���[1�|K.O0�2��'rH��d]Mqr�@m��I�
ܳq���!�$Q5~О<#u�W,S$�@��bK��6�%��|*M>i�
F1|Ѣ���=���h�z�Vt��;�?i���?)��o��.�ON��a>-"k�O`9X�kčf1\��ulC�G����pG�_x�ē��������ޏ6{p�+�<K�L%��;�OB5��'%�1A�FhX�V�&d�0�(�(;D���`��/���#%�ZE�Xk�9D�,q�V�*~��Q���	9 ���>	�i	�'��%�2�e����O�S�1Y�u8S�Ɠ$  ����/�47��qb��D�O��[7���=�?��	 �Ҽ��ދs��	G$ړ2(��G��,_�R)V$3H�=)���7���hOV(�w�'A�"|¦ɶ7�d��&A����f�E�<1v��@!����A�S�h�qU��|X�,s�O�ǤU�C� �$f7=H��_��e��M���?�-�ج�-�O���p���a#Dn
����d�"&�>4n�|�	[�S��}«�"��c%�(=d�����?�3j�X����d�B��0q��"��P:�c��O��'�T�O?19��$}�D[$�P*Pl	��"M�<qW�@d��6L��g���ƅN�'ъ#:Ė7C��i%)f��x�H�(p�f�'���W�2�'0��'p�*pݩ�i��8�h��s�jIҔ Ϳ����
�<���^[8�$���]਋�"Y�C��j%�<�Q��R8� �s Y da0����Qy�c�I�<� �����ӓI4����(�%^(���$	*DԱ�ȓ- Jh�4iɀP]K��L�)��n���HO�I)�$��UfZlZ&�4�ؙ��Y
eH�C�� �X�D�O����O�(���?����D�L%�?1��e���"�k���kd�I2`8�}'D)�~�Ɗ�vM��9�O:rX�P����>�ٟ8�7�hK��{& B%�b-�D\��y�	N�c��|	��(P��q0��^0�y���l����c���,��J���dKڦ�'�P�$T�M{��?��O�*��-�V�&Q Ak�u��ٴm�^�[��?�f����՘���� i�P+!�G�������)�hO��
E��`�Y�ʳQW��A�JL	Uvԣ=i�&Xş�"��i�����v��U�-���!�DD�,��l�FN^4H9��H�jTa}bK*?��%C�9��(�c�&M(�0AP}�H���
7��Od�$�|��D��?��<���!��K� �GK�q�����i���h�f�,�ic��M�\�a��|����\�'DqJ�i���'akf���E6p��P��%�D�v`�*��
�N�*q��O��>58�"J	 �U8�&�����'
ȟX� b�Oґ$�"~�� �7":����V���Y0s��:�yr�_qi�u9`H_��t��,�8�HO8�G�Aܻ,�`�B��qRi���O�Zd�7��Od�D�vܺ�
7+�O����OT�$�ߺ+��+���:�#r�<Z����e�^����ny��*,���O���:�Ǌe�"J�a���P�R�S����bJ��)̈́Y9��"�'K:@4��C�7؜��'N
�3�\�5�:թ5�F6��=#/O�H�D�'"�'F�O���&똕u���#vjU�#�r=�C�I@aH��靽NB����o&;�7��V�����'�	�~e�Tg8�Lh�QZH�j���pQ��AV�'(�'�Ҭd���Iɟ�ͧI�&�J����fL!C_�I�T�!'C�2T�@���*\�������O�	��#�fPy'	�� di�J]{�8��b� m���#�͊�7�'=�����C�ɦ=����C�? ���Z�\)d����PF2��@B�i��D"��=�g�K1#�2ҵ�;�(tjQ� D���ϣO��kw;"�H�b@�>���i�rZ��b��Ϗ����OT���+'H�[��	=v��0�]�I��7m�=}ml�$�Ob��W�|%�m���
j�|EXc �c�IΧ{�\�!�(t��#�݌f�]G{B�� ;�JdِX�����׿���	pr}R��N����*I4~���0��?L2qOFM��'����!\s̭X�)R�91�P�E͟F����Ѕ�܊�1E�B4��E���E����$t~k�}+4����}��]��=����$�oZןX��U�OFo\r�'v�ABŅ�EO���(,r�̽{emyӘzvn�Oc��g�'V��׍+s-$mc�Ő�R��I?I��#<E����J�ӅLL3(�l�G�?v��a�9�?�v�|��i
e\�c�F�bX����άK�C�	<z.a! �ʿ]��H&fM/צ"=A����K͈�	6mϯ@����͋�.<���I֟���d՘x��蟴�������
�u�����I�;az ���]{���S�ihr���p��Ox��ҩ������u�!o�Q���É��=��*�k*���7mD��g�'~)r��P�C3�K�%�}�pcٴ�?�`H��?ᗿi$z�gyr�'��wf�i�Z�;�v�su��1�'|�|��M5smFhC��LCצmʃ��2�MSQ�iB 7�#��������<9$�Af�Р����:�Uʧ�M�RB!�V�W��?���?������O��w>hG�ൢ�@� k��;啟.;z�{�-�ZN��k����v%�m��%�%P�Q�@{���mnPX�UC���#¤��kR(���ԥw �ā��$9���5̡-�@��4��Q�RN�!��+3�S#.:������X�C�	��
4K��K��q�Q�
V��C��++�1y���`�n�`��	,3�P�H��|"�ԫf�0��?Y�O�x�P1�(Q�|H
�LM�ܹ�ܴHz����?	�Ϊ!��g�o�
��n�&Wr=��>�`�`�Ɏ�r�D��g�c��!��ɲoIJ�àAQ�9�ZH��b��A���;_�L͐R,=}Ȫ�y�%�	��͓�����=IQ�O��$/�#B(����MФh�������<�O<b���~*�j1$Y�D�\s��'�v�'�q�N� aڥ`&
' ��|�'�ԩ�A�'P��'��S�	R� �	ԟ�"��|�Qw� ~��
��Ӂ�MÒʗ�~�r�P��K�n���RU1,��SA̧|]4�� T${��eJӏ�6�����'���˴���$� �h�J3��k[w�
�����Ӈ�|d��X n�u�ɒ.d������~r�'��)�))}��>�b��8{h}�o���yǈ�+����/��4�d�����HOn�F�t*� Z���¥e�(�V �#��3\IT6M�O&��_�q�y�U+�O��D�O��d韐�n��D#wk�/2>&�@T��y#.݁�
,E��qZ�D_s��VF�F���Ɂ_���[3i6EM�t)��X�����%����g�S�i�D"�M�|Z�4��wf�}}OK{U�M+�,	iʲ�{��<��D�s?q���hO����`���&�Ϲ`��LR��F�k`B�I:.;��pV�hѨ�� �� �6�\���d�'��I	|���x�A�P��܈U�E�b��@,Ka��Iǟ��˟�c]wQ��'e�)ɪJ��ő��ر����&�@�_��8��nV�-�|��
B~���i&��q�^���(�1;�EjW.ץr@��b��3:ZX���@�2i#�BM-�M�u@KQ�X��=��O��Pɑ9/��h)V�ԅ�4ȣ�G��}D{��I�u�B@��C���Rr@�Q�C�I5jW�@�2-�8���B�������'��ɗF�Ԕ�����?-
d�@�mA�ȉ�'�hq�e�o���5�?	��?���\�Q���@�*R��HUMN5�� B���������	��=
WўXp�]�P`�CB��:C� ��S�Bɺ��B�W����f��V�8(�EC�?,���K�P��d�Ov�>5c@"$�Љ;r��?.t�s�"�>�l�|���"�,FՂ�pv �D�NX�����������Y�Z2jv�`Ї����8�-�IßT�I_��J���'U(a0��:`�j��ʋ����C`�2�:Dk��DB��� z��S;�2�O�1��QB�O٪-&���SH��1��q�J�O4{�ä+�Y+�ʃ W�6�K�w�QЏ@�i� �O��	"F�XB�h�@���2�~����'���ǟ��䧱�	I{$���ӷmw2Ѻb(��C�ɬ-�^T�b��mp��0�^�b�#=y ���!�0�� ��d��h�m��-@�4�?������վ�?��?����R�)�^M��휍 �i�,�0��ӱc�<]�]�!�B�~�+�fϮ'W�T�'��Aq�Ĉu��UKנݩQ�f�!dK[�w&N�@�ˑ�zc|�"�@��B8�ehL3d�F��'�*E���/,�i�FY![h��.O�����?ً����� �4��Me(��2GQ� 	ӥ"O�i���4l9��,̆G���{6�i�|#=ͧ�?a.OrD���J�z���(V�	H[�Ę�%��8���O6�d�O�������?�O�H�˵�Ii�L�R���t� �zՌ�.m������_��#u��W�џ834�
tԠ�q��0�8��d���J%"r@�n털�s+�%: F�n�5}D�����3�I��~B͕�G��f��5K?P�#��Q�]��7�:ړ�O�����S�c�<��J=��t�$"OZ��cS!�8 �r���*��L��T��"�4�?Y*O����I���'V��FB�x�g��J��#.X�&O���'��A�+.L� '�(%X2�;E]�vLT��J�0y�Ch�15� q���+�֣=�E �{��t��/v0�0�a���u7l�.kT���!ٌ,E�k�	1i�b�*�͐Ÿ'6r�	�L�}"U�Hr�����9
&�Vn}2�'%:A�)'Z��w�C��:�{y��2k���)ߦr���4m�/=�h�j� ���?�����3(����O C�Lҳp6<�Rc!�}���13�Ԧ	��Hȝcl\C�m 
�l�a䕠��	7��3m�(Y3K
Q�X���ґD���'�r��!�� ��\�w�0���l��S�'%��!�$�h�:�1t�!?�Q��qI���O�S�D��#<�ʤc�����������!�d�5��0g�źfiZ�CCH�@ё��q��i�V�D��g��0=������]���nZ��\�	�,�N��C,���Iϟ����?i�	t?�xe��=���r�ٜ+� � 3E�g��C!�5��q���J��I+��,xr�[�����%$�� �x���l�?p`�M����i�%�0(ID��i� H�	E��D�2|p���2�9�a��X副�~R�' ў��#�(���2aH�k�*Ч�ڔ�ȓU"�,�� ���"$Dҥ:M	mZ+�HO���O��زh",�&�1 Q'
p`;�V4w�B��?����?AԴ��D�O��?m�����=M�"�"C�T&�B�12���
����%�L0���s�(@�'g�кA�������u�<A� z��SJdԁS�@7c+(I{�L���F-�h�q�{�#��@Y�F�e���eT�y2��5����M����:�7���B�*P�'1N0LI,w���ȓle�eM�?II aYp��_��d�'M 6-�O�4ڔ#P?���B�b�QB��I�@X�\	��%�ۦ�����������AC��^1:�D�38�>��G���D͒#��k!E pQ�i�A�hO,m� BH-�V�xC�Q׺hȇ�v��𲢛6<��1��E�i��5s�NQX+\�ʠo7��-�~��'bq��!�-Y��2�K��?����X�D���0p�l�s �-(��dG^84���$QC~2��Q��S���	��B�&���QO���o��@�	Z��Ȇ�%�"�'7D�i�䙾���nJm[��yu�uӲ �4D�5)��q�σ ��!kF������)w̘4I����J���
�*:�d��"D�M�;���� ^1M���H� �$��U��m�|b�kK<Qh	��@�� D�C��?�S�џ��H>E���͸S�4œ�O�Q�@�ʳ%%/!�� ar|��(vښd�EްbF�O�DGn���4L�6Voԩ�� ��.����smeӬ�D�O�-c!�$z����O����O�����?�18v~%2�O�i"����&ʪAAd�( `۹CL"��愋4'|45�Ѻ�O�x9A�+JR�	 |�H� �)s�@�E� ��q��ǌ6��R��Ez  ��!�|�L��#~4O2�@f�@=G �4#��Դ0Z8�7]�p�L�OZ����-%;���E�B6�s���s]�C�I�{H�@�Y�
�4 "&/J3�7��V����|F�5J)�E+?Fz�H� ��0EXA-^�B�'��'-�ם�����|���D�`$2A{DEؗT���aDӥ'ԝ��@�Ht �v*AqE���F�|dآ<�� �H`U)����KbZ�ەaS���D�5��?�8�wa�jx���C�I9n�T�<نMEԟr7fȗO�f�a�F��3#�T��.C>�y�H�H��5�ŉ3fLHB�e��y��OT�<!�W	�>&���y�f�2�������'� s ]����O��ӹM���c�G�������4"6M����$�O��DB銐����	K�ذ&A(:��ͧU�Z5�7!	�7Dh0z���  $G{�	�?a�$�0��	�-�� �cN�8��I�5\���C��V�<��ƿ
�ў�Jc-�OV�:�ӠIm�9��e�z�a�O	[�j��?!�}���Cq�T?^��0�ko��!��	�����2��)x� �6\���<I�	7"�6չٴ�?����iL91\���O��"W��C����1�6��� ������)�q0�K#��X��d)�����1��0ʉ� ���L�C�∭(8���I�: �@�b-Y'd|P��� !	{9D�$Ɖ8����F�����M�R����I��(���?��'���3�ϊ�-16d�g9~�,���� �L3 �; �41����	*!Z�"����ȟ��s��D��(8��9Xr�@�FVզ��	ӟ\{'��a����՟ ���l�Xw��ET#Ll����\�w� �P� ����U%ۦEz�Y��
Mƅ�2��|���d /x��M{�&�� �%-U|��pE)�)gT��q��6g���4Y>��c�(�	_����1�ؕ ٬h�v`�'�x�)���?1����'��Ɉ6}Yl���°��2ۛ)�!�$�cL��5���S(���Ԯ�#D��ƌ3��|�����q�~���팸T6�q��3��\3��R����O��$�OtE���?���)Q'o�l�@�5�= p�\�7f�����!e�y�'�5P��0`�'i�dDy�Ce��A�j-4�����Ab6pj�EW�(N����Ğ.��w�N�,7�=��C6�	�hO��$�j.���+�AED�p`O�i�JQ�ȓC��Ӆ��-=VN�q��Q%�M�ȓhr���jP�)5�aQ� Q%5��u�'|�7�:��C��m��������ڷ2�@��O��P��邌ꦩ� �ҟ���ڟ�y'���.���iV�^Ȧ��PY�c��y��`R*@'t�A*��/~4Q��<c��<�� R3@U4\p���Q!����uKG�]3;��ӳ$�0w�v� fW�!��<!�n��,I��)-E��␌���vMA�OA� !��?X�-������7a}r""?�f+9�����Y���X��Xt}r-$�7-�O����|��(�?A��,�$T�'�	XS�`o��x�ZFw�ȕ�"$�	2�^imڟn�=��4���|
���F��+LzSIR�$�v+�O��Y��M8���hV���Q����%@_Y�L�n�����'o��� �IB�L@e�C�D�����R�b�Dæ9��4�?.�lb>�P��%kb�x8���v�|��q�}R�'2�'[�	ȟL��ݟx{P	ƤK�z)&��b���%�Z�a�^���4�䓒?�\?��'$��OC��嬂.�F(�4Δ'3�Z��q���D�O0	�/<���$�O���Oh��;�?aR�]�=l9�a��4����$׮|ڑ#��i7����h�XT��/mݩ���M'Ke����0n���rj�+=�Ā@
> ��:̊#�$��U>����(0Xf]���cL�edʳ�ѷ)�2d�ʹ<(�����شpC�'
2�'����RO�ѓB	�>~�cw@W*
(��ݟ�Ir�)ҧr�p٢e�<G�lC5�
>�~�lZ��?��4�����'��$߰ �(t�@� *d�r@�I2\ 8�s`��q��D�O$��O�M���?A���� A�P
#�D�2Uع���
�v�<�爇�I���Ӳc�F$i��K禀Ey��{��T{���Z�|��	�0g�FW�.T����Z<%f �#�˙�fa�H;6�I�ac����5�j}�Ν;�>p��m�$[B��ȓ58֠��A�y����5gդ�����cI�d����h�`�)S��"ܞ��'Z�����0k�}���i�R�'p�	
p'F�FOˢ%Rxp�Vꋩ�?����?	��?����?Ɏy�O��� ��	�$u�����F*&�H���*3Q?����J< ���chB�C�ڰ�2ړK.(������l�	J�T��B�,c�1P�"O�H`�X��=��J!xw�ـ��'�(>��97��s�X	B����zL�'� u�&kp�����O��'Q�|��?��� �4�HE��)�1�KTSa�_>'�`գ̔	�1�`ρ0��'��O�h(;���Oږi�g���K�fx��'Xh�g딮N����g���2��2w��ڥZ���!���j 獍A�`�)0 �,N�Pj��ss��������'�?1�'k��k���py~d���լWS�q��'"�QǏ��v��2b��$<ZԠ��D�Z�Of��2�(��2�ˡ}
x��o�*���O���Џ]���'�2�'�a�����kyN�ċB9$zjA�@�2F�� ��t�ڔ�' H�`�T���A�lt��QN<�(��uh5���J�hАqBРH�Q����A[.O'��P��>.�H���:1#K)�MC���<����k�Țe�H\�chDMy/#�?aE�'�����*�>}p��N�݀�'c����B�-�Bp�'�N5а"ӀoӠuEz�O��'7��� j�)P��eX0��)��U��6�2��'r�'}Bi�U��ߟ@�'~Ʈl!��5��y7D�tƵkc��x7<U��MR<J-$Ѳc����ODQa��J,Y��ţ����D�'��'vVE��KC�`a&��QD�8@Ӳy*��]�*�4D5,�D��*��� �킡��:��@RBN�9�j6��O���E��4K(Bb�3�x�JT`�?�0����b�'�&l��)��e*U�v�PUZ�O�o�\�'�rx�<���O��S:V��h�"A�1�x@P2H�/~�b�R.R�'��L�b�j)��#4�6m�O���(q&�,�-J��d�揄�ʣ=�ul�=d���JK5��OⲰ�g�;z��0l߁���;��d�,��I��'_XТv�Y �2T�ǿ*vE�&�i�r�|R�'��R�h������E�� 	�މx���1�x��T"�Ms�Q�̉HI>���<�'j��I,�� �e��� X�g�C�]�>�C�U���V-���M����?����b� �?a�z~�ZSF�7�<+��F�b��E``�i{DtB� @�w˔]��P�3ipx&A'�`E󩌄A�q�F�C
��CѠ �C^��ć#.�j�:U��6=h�ԉ��ǜ{w,<�1���t
t9
"f�|�C-�#����og�#���?��ݟ��N>E�t���6\$3�O��g�٩ �C�N1!�dM�I<��
ĥf�h��cᐿ�O��D�y���$���L���02��M�,�H7E 1S�7m�O"��@9�b)vF�O��d�O(��������K���v� l��Aq�E�G� ~d	`4)ͬp����ӽlJ��O�"�1���M�I�e��!���7I�4'�4"��%H�zx���f>ɘ���|�G@�DqxgD��y��R6�x�퓴}����7�!����O�"�=LO*�[���ÁK� �l����A��x���<@r|��#�=�`d"v���zhڴ_Ƒ��O�	�:�dx�q#	�w0u��V�)R�Q�cȘ���ꟴ����qXwn�'M�ɀp%dI Q6\yj����G� ���hD���I.��S_�L3�m
�:�*Di�K��(O6h��D�%esrUq∐�
���nS? &t�FF�:� ���f��M ��<:a����=�D�=:g2��z�ū�'N6�ʽ���r�C�	D����f�@��q;v΅'&���d,ʓ8�N`�GQ11��z[����&�>���i[�'���fgӢ�D�OT�/~�	A�A�`���$.݉M}\7Mހ^�.�d�O��M�i�,��.�-��q����!#���ϐS�p-2wU��8t��`X�K�XJ��I4Sָ-Bt�ط��� ���&{e8�;���8B����"��Ls��H��=��Y�G�F|�'��y���Ol�G���ޣ(�(��
F�����&H��yR��+�[0N��Rl��ͷ���hO�x~���6������ynD�P �_��$�5o��oZɟ���M��FG�$��'ڜ�gJۂI�Li7��1�@)Z Oo�lu"�ϗ��Z!��bݱqh�M���V�2�\��1H8擶$.��%DժN<p���a��4��)f.��J7#��q
0��)�KPM�;o�����[>��O��][6��"H�4�R4LW6<���R��'d,���ɧ���X2E��8�L����x��d)V�&D�����_0q\ꑹ���!(����:�	ȟ<X��4�2�r�[�&y�"&,��AV@e�h��	̟T�`ɑh�
i�	��P�I���XwQZcePu�E�(A �@֏�,7��:*O��a��'_��"���1ƀ�pK��e���)O�xy@�'��ѩ�A�&(��Y�nu�(O
����'�B��DG�Hi�I �� ti�!�o!�$�\z��	��A�� ��#��f�0��|O>!�.�|:qY%̎'�P���2h�R9
�"O�T�CG���T��b� V�hd��"O����p�l�#pͪ�\D[�"O���Ü�'�N���ό���H(�"O��-��@�ܱ�ӏ�;b^(��F"O�6�G;'*�80.]=8��A"O�죄ƞQ��ix#ӬR�2er�"O��j$A�(�P90�g�W�^�H
�'b4��eJx����U�It�~�Z�'�mr�Y��p��G�n�� @�'+�����	IJ�
��4|�ژ�'[LZ���	Ud�.�.)��ͳ	�'����c!۬P,��F̢n�4A�'��-GaƸ7����A�żg�V���'vذ�G�D���#��b�V��'�0�����G`�8��l����'C�I��BR�v��ܒ������	�'d@y��"� �����k�JjL-�	�'�<��)ݲj,&�H�d�13�"��	�'	f�����C�$3e�=1<N�2�'5ܕ��g�`P�Q!#X���'Y���3������R�Y�Z=҈��'\.������c,��#�ݢ��y�'�*�[0k	��I���K�<)�'����^�|_��
S�Ռ̢Aa�'��9� ��.�
q�&�/o� ���'A��Ef��o�*�����&��'>]V� ,}h���6F`���'��ʓ�� jB�[fb�{+����� T����G�l�.��Ђ�Z�r�"O�}��@ /���i�a�&�.X�"O�̓�b�!f)�����<�"OhY���Y�3o0-�D ֵK� ���"O�C���#$�ԩ�w�$�� j""O\���-ɞ�r���d���ʑ"O�����g���С����q�"OP�)7�o����D���F	0�
E"O�͸�%�>�"���ڥi�՛�"O���R�ذ@c,�)e��I����"O���#G�=9���j���`0#"OxaIr����PE;P
P�� !2�'���˔f5c74�[�M�2����'�hq* ��M]Ztz�L 4�R���'�l-�T�K��&���aХ&����')�´H��s2�H��E*Hv�t�	�'p��C�Ab`1e5K�h��'0����,�y`����L��'�Į9�~�	F�O#G�8�
�o#D��Ц�I@4��fOw�Ȉ�p !D�|ـ�/g�1:wƙ?���Bo+D�H*b|x��X�E�X��a,D��1bO�;�^!䩚"T�hqvN8D� 0c+U�t�1�͂,k��1 t�&D�����	�@�u�@$�N��c�.D���&�L��<8 m�3RJ0�@R*D��I���IV���$���^�˔))D��EB�#[v.yQ@�O�T�Hܣ�M"D�Pi��I��t@XE�K:�*8!D���Ҭ׿>��%;@��,a�$� D�D��I,$�X��
D�m20`�1f"D��(Q�JV��̪��|$j�p��!D�T��f:h�&�P���G�P`)C%2D�ȀQ�F�E<�ӤۆBT<���%>D�8��Т
��1� 
�8�,��ǯ=D�|*�!G.g��D�SHB�.� {d�:D��2�mʰn$�L��T3|�֠:D�� G�?j�z�����!R�8�,8D��,�cR�psN�S|T
�M;D�$�ի�#�Xui%�@�+Z<�N.D�|x��Ah�)�댞=*��T�!D�XjV��W�rd��
˫1��؉sB%D���I {��l+�n�E�|�Dm!D��u���8��t�W�Bz���-D���0i�P�Ļd�K����p�1D�,!�cQ��Re�w�J�Ͳ�'0T���ݸ2o����1e�r���"O��!��OD�A��ߟU�:��"O,Uk�; �1P�
][���3"O�Lѵ��6<d�`�	��|��q�t"OH���Ԝ,WԌc����0�#"O4Y*B!��L��H��Ѳ4��"ODea��Q�R���Y.?S6�{�"O�xjDo��45b!K��B�Dq�"O�!h!��78��u�c) ����J2"O�U���B)���3�ٺ'�
	��"O$��F�5�6 �N
�:�~��"O�Ы���}�T�����L�B"O����A,N`���
!V{�\1�"O�@�d'��x.|��#���NR�L�"ON`�
^$�qq#�ԋ_�Ȱ��"O�%�4`�-d�$�(!�<3�$�j�"O�@�@U�0�.m�B��#�4L��'1̋�I<�f(2����\���
��� �M)@'�=(������G9\	P��"O�Q B$_���p4͟
u~.Ak"O<�:w螫I'�ĺ�̑ct���"Ot8pc��
4~�u�\�]��<��"Od�*&��11^�r�A�T�A�"O��x?v�qP��1^7nx�"O�i	G�Oh����#�*�"O��`��#������x�U�"O��Ö.�l;$� o i�>h��"Ob�f��5c��H�n�5#���xP"O�����Կ9Ӵ(�PNQr��4[S"Ora��F�*;H^)
&-� %+��C�"O��[m���L; Z�'�AI�"O&��@ RJi!1F�ڥ�R"O.$�������@�  "O5���έ;"F3��+�Yx�"O��1EC�R���A�+,%����"O��k�Ʈ/6Pb��y
 �"O��K�+�"cΰy���;1��l�b"O��������T�܈?�"�(b"OHL���@֊��m[> �L�Y6�Bk�<���F�h�Q+�.��(/l��!
Bs�<��8w�X}ӆƋ�C��Ҧa�v�<��gӎc��*t/�	�0
�t�<IǬ�#J3��h0�A}٬L��jAi�<Ase}|� �'�"��A�f�<�E�n����d��F]J6'�{�<�$���;��|{��Ǩ31����`�<�����L�B���vL�9*�Ay�<	1Aԇj���Z��� L�����t�<Q����Jy[WN��-�NHrt��V�<�@�X0(.����P'���n�Q�<�d��TO~�9ր�]q�	�jQB�<QD�σ~���#�:	Z4ep�o�d�<$
��:��@�Qe�3F�]x��WE�<�6AJ4���ܳeB�`aC�<�ª�3l�Xa��?�<8Ia�VJ�<��m�H�����G)74��mRC�<a6nn����l̑.���]�<q�iC�r?�h�3�݆:o>X���P�<1� �(��Ko�M1˖��n�<���M�Rj@�*@bN�I�jE���D�<�P
N�ґo��8Z��q�GX�<ie��.�� �,P>S�v)�焀P�<	�_(hS��pՀ7/��]Ӳ�Lt�<����bx�%oV�n���ҰXj�<�'^�n^5��l^"1�m���l�<���˕U(�x��%Q�uل��Tč}�<���G%\*�a���QK��[u(VP�<�7�§Ǭ��3C� h6Sm�<���4&����͘�L��PH��i�<	�/�b��X�����m� �k�<qN_�*x�����e�ʜ� Cs�<y��U8���-�z?Lۣ��J�<!'eش��1Xgā-�0A�T�z�<�Q �N�@��[k��� ��v�<!u�I�YB8�{�O/L
���Rw�<����,4@U���T�"�|�f@�O�<2K��)�j�Zdǉ�G�����WO�<I7'H+}���9��-渜FCN�<���VH��P t J�l�HHU�J�<i�3� ���B
Ǆ�3DH�<�5���[r�� � =Z��CKn�<�����V/́ж$�9�.pif�Q�<� l�Ar
��o���:��*7@.�""O�)7��&j���;SA�b����"O �I2.�iܺ�`q'��G�^\��"Ol��쒍o"�B	�~�.�`�"OH|����4u�����Y�O����"O�M�ւ�W�<� �C�%'J�R�"OX����"_�`����,u�8<��"O���i��ZFYX#�C7~�ZTP�"O0�Pl8]d�������c�"O�<��B��Rv��{�����]C4"O"ٛq�F�+�l�б��&Y�āZ�"On���Nq:,ˢ�H�;�2�H�"OP��R��3�|�� G�<�:z�"OH�o�4P����ٞJ�Ȼ�"O
MR�j�l�������:�B��"Ob��ML1V;��T`�+��Ū�"O��!Ƌ��T{3�8n�>�q�"O�E+ÏU�O�K�lQ-|�&)��"OZ��Q ��Y��\��e]�t�tʲ"O�h[R閼:B~���]���v"Oh�� �(A<\0G�i�TЉ�"O�A%�� b�9a"��ޢ�XG"O�����p�j � �_�x���"O�ͺ�X<1X�C�f�2D�t�"�"O���g��I�,9���-r��X�"O|�`r/ .��zR��.L�I�0"O��@ .�(�U���݂Xjhlr�"O�dQ��܈/�N�fM���l�T"O
T��Л%�<c#,����U�q"O���s��V�F�AfB��z�ڬ�"O| � D��-��ΝneD�8�"O��h�c�5v�p�ALS�F���"Ob\Q˖�~Xb��ި;��P�"O�E����Znx�q���ގO!�d�#V�>�ʁ��K��맡�?�!�Ȝ0��Ϟ:G��Y�%.�`�!�D�n�(�Æ�`�|�2V�;�!�$R�<�r�&L�Klh���!�D����a��a@&o��l��FZ�aB��4qI����ɢi��E�e�`,����.D����V /A���l��+FD�(P�?D��Ȅ��f�z�"�Y1*� a���#D�T �k
B����g�XE���%D��
�&�"�2���]'.���(��8D�����	�w�
LZ�Y�R�$�*7D�ȃqbз����N�e�$��5D���p�D��
�E?w3�L��'D�(�_<p_ ���# w�iq��%D�"�Ƌ 4��TG
����9D�t�ǰ'�l����t��q�P-3D�43��[$.,dRS���"�z��R3D�X藤�('���4*�kB�ꒂ1D�Q��`~|�2�4r1���ч/D� �q'?Ѵ�(p�ܨ.
(�.D��I�����~�hC^v�UQS�,D� Kg�A���آ��?Y��X�C�+D���7!�<�&1ks��0������=D��2�F�P�>=�Խl�������y�J2jX�B�!}E �p�nH�y�R>���ڤ�F�bE0U0r8�y��L�Q4rEp��)V|��"� F��y�'Y��X�"��%<�Xs䈌7�y�O�X�L��1�C��	i����y��R��UK���,E��:&�F�<� �����-T̕�e��7�\F"O<��#�#2�u��'؟�����"O�� R�|����霙P�F<�p"O���ủ5D���i`��!:��8r�"O�%y7�ߑK�1+6�\�.�8�ɕ"Op�q59Bm��#Fֿi|!�"O�9jE�S!^d��JŅ 6=�>�A"O��eᑡ8�0Ib`ՀN�Nɥ"O�q�b�WdD�rM�X#t�x"O� s�	� L*���b*���"O��X7�R�<�FIL�$�JŁ"OBIPÅ���R�5M�����:4�!�d�n��e��R�����P�!��|6��D
�,A����U@X�p!��46�BA����'A��ȑ�Μ�!��S�%Q�q�4��=x��d����!�J�(�:Ů�%S� a*DW:-�!�$ѐ~3��9�D�m�z��QC�5	!��$i�I��c�J�ڔ�����!�Ђi�|�R1^%���Q	>�!�ۃaA�8��Kx��� I�("�!�D3]��|kA��]x���ۥ`�!�D�?�u����<műp�ݠo!�"@tdz3n'k� ���A�
p!��@R�d0���X��p�Ptl�"L!��:1z,l�!aR93<�S��N�b�!�DF�R�:�	�29-lū��/x!�D	�Рi�+_�.-��СjO�k�!��)^/��:1�
j�4���g�!�Ĝ�H3ԘJ�i��1��%9[!�$S�v�&����^8�,�R���Hs!���!���S�K6s�d���ow!�DC�>¨Pط×�|�{��ߔ^!�DG��،q)jF�10���E`!��>3��IQu.�=eH�\a`��}!!��9S (��e�B=ɓ���+>�!�$���͑CK�!nݛ��@�,�!�$V�?u$�{��ӾVeك�L�C!��1N|ܐ��[�&��͓A!��
����#,�/�F(l
?Qr�B�ɚi��A�ІYtN!sŀܩ%vB�Ii�Z�{d ��C������[�
�>B䉵��(�bd��P��]��X2*�B�ɡw; �r�c�/<>�Ţ@b�$*� B䉼G2�I��G0s�R��FC�0C�	�Y�܉T��62�HS�J��$C�>7��ـ���)��AA�F3qC,C�Ʌ��=9g�Μ�XQ����HB��>�U��C�:+R�X�H9_
B��M7��j�ƆLp�$S@�-C��hE{��9Ox���ԜTب�rkI��)�g"O�e"QEW�tX�-�1EE�['�ACA�il8H��ɩ"��P3J��i�H}�t�',&���U0��}J#�\��F`A> a��3�­���Z9�$J�9/R��>Y����D�.5!��Ti�f�p�v���y2h��� ����5]h&yf���y����q���wf�/S	r˶o(�y"�ؘ+�����C�O�D��H�<�yҦ�.']�� d�Hz,Л��D��y
�����iB�UF�y�T,��yY�iBv��蕳R~ (���*�y����O���	B@SO��9s�g̀�y�H=Jk 0���@�X�����y
� &<��͛�yV2��A�3/aj,�"O�8 ���m��A
��W#W"j"OD����Ab�H�1GƠk7~�"�"O�y��j��qj�1դʷ�d*"O�dۄ<Zt�IҢ�&o��i#"Or�QAfQ.NqR�04T�sQ�Dh"O�2���%��eI`!��6VqAd"O�l�Q��Z�"�a��)�%�G"OT�c"<ILQ�Ο
A�x@$"O�����[�4V�dn�j��"O��h�L�y�ʙ2�۶L�Y��"O��[1�J�F hA�U8��:D"O�!�f!�F�=���`Ҕ�"OF)��U�1��p��
����"O��&��?o@�@� jF:w����"O��!S� �W��A��'ͅ*y6r_!��(K*���Շ]�gx��P'�@4�!�(r�9��=F�n�Q���$-N!�Y�	Dy�� �����B�IB!�R�F�
8 q�́e~0��E\5h1!��[�&Et�{`�^Y�`a�(pp�FxrK$�g}�lWI�NH�aC9M���@���yb������L��bZ�Q/�M�!e�H؟���i��,�0��A9��<lO�D�f-}�Ɲ�\����KԘch�A�O���y�eQ�HfA�0�
<nܽ2�M���'������d/]�/\�<�`��Qnh�(aD!�y�/��!rm#g��8]Nl�e ��o�čB���Pj���dғ-��c�$A�T~b%��dT�z!�$�-k���;�υ0p`���D�Ǚn���,C�t�����	ۦ!���.h��$[�/������$+���b�O���G�7�hɹ1��b�jt"OZL�1cM�G�0Z�ɘ9<�L���$g��ħ{NT���f�H������7}�������B㊎�d"
U@���uـ�G{B�'��@ `t�cS�D�L��'	��I��ķI{�Y7��8q���4ɬ��d�q���(��D-dJb��E��h�a{�j�u����4�Rb��]�Y{�JҦv7�a�ȓOb8A�J�L�l8�F	1��>�Ӥ`Ӵ��I]�}�"E���6����u�
g!�d��m�Tc��W��в�����8�S��M%�On���`�%I����c�d�<�4O�@U���P��n��1��� f�<�Η+;�����M��"��Wj�<����)Ha�g
ЇF/�HK��Q�<��)� ��x�%`p�����Js�<��V���l��%�t�z�B!��H�<!���,����m��+䄉A�<9��ЩW��4s5@�Z�^���O�d�<���9V\�����i�$�nN]�<q�h^,�<��A�t\܈��b�<�F`��J���$@S�@R�0铬�G�<y֨S"D�Sm�s�b��E�D�<�ơ�-$wTy��H;0���F�<��ˋ�DH��
�Ā�(�@}ɷ/�|�<1f�B'L*L�sb��?�y�/�y�<!%�Ր-+��'%u���
C[�<� KOW����S�.�7��W�<qQ*y��	���R�yk&��)�N�<I3ȖM�����L�j�8�eJ�<	���Lg�T��kS�4_�쪱�A�<���%:����a�\9�زa�d�<����R��CRi��?�6�Ҁ�Ya�<� @ � �K�7Yp�a�&~��H8V"O���-Y���[7�N�9�Z�	q"O�m�7��7 $�r��E�
zh��"O���P����x����u$<�6"O�%j"`Z�f����	>K����"O��Ej� "Q�h�ڈsԸ%"O`�X"���3�8x@�O_�w�2}��"Op 3%kQc㘘AD / �j,��"O�#
6&��uZ����L���"OVm�S��)I�~D[��L&:�ݓ2"O�$a�\�E.> 6"O|eR`�Y��,����B�q"O������R�� ��$&,d9�"O�+t�Ft��@ȓMt܃@"O�x��e��2�ǝ0aZ� a"O*X��غXR؜��!#��u��"O
��0D�!l�8��`�ΉX�(a�"ON�R��?h"|����),�����"O��� � � � �W/S�p��@"O��@�'e�ܣ3m���F { "Of�1�o�2R�i�`�H>C�|�� "Ov�ؖ �3c�0ّ�E��s���b�"O�$R6I� Mi�@���+(�x�"O�8�r̒�]�޸�e��ti"L"O��BgL�Yh��맦��RV�݂�"O����'���(�BF�Q�"OD�*�O�V��t*�'�x��"O�USD�T�1���R#*���"O�ps�ȥTc��`��I�xb�"O�aa�Bڒ ��]��ʌ#�09�"O�	:�$@�=$XYx�c�
c�c�"O��� 6���w"O��Б�"O�H:���)+Q�)�A��v�C�#�_�<QԀZ0{��I�עwA
E�rI�Y�<�φ�^v�$���\��2�"T��R�<�����n1)��&L��L�n�f�<�@Ї9U:ebE�P��X`��e�<	�̙�k��s�IK�;\�l�v�f�<����30�X���p D��p�\�<	foB�f����I�|rA�P�<	tj�4 �4t{�+��1��iӢ��q�<�%T3W��T�)�:oE��M�S�<d00��)�g�5s�&9��M�<���� :  �   $   Ĵ���	��Z��t	�;B���C���NNT�D��e�2Tx��ƕ	#��4"�V���$V��m"|`ѡ�,��Xb��`��ug�5�&�B����M+¬B���`�v)ccbL,�d4��7�Z�yu!U XO�Mƈ�+6���"B"T	b4W��)`R� �N�HM�p�@搥������e�"t#@�K�;����#L?L��T� ���K(��r�E���\ap��'H�Z]p�J5���VA��Z&Fm$y��
[���,O؀
b�jM�OJ�ˆÓ�C�j����=3I��E�Z1��&}�@�<-�L���x��ox"�h�1�0m;tL]�?������KaL@�Op(p
�9�PH�I(�y⮚�B�ι���O�iɜOPQ9ab�)tK X@b�88��eF%W#;%�'�kǄ�$�(�%>�Y�X^p���*O�S��ĳ�ú^~�j�:�$�1(d��U�|rbV!gD�(-O��A�:l�	�u%��:�+f�'>zU)�-���~R)~�4�g�Ρ`��CҞ?�A�n���@	����0O��WA	\tL���C�-
�I�j
z�I5� ���wU�ት�i�F9)�J/4�@����	��4;�ď#aK�8{(O��݃�܈q�%b�hݴZ[r�+��I��Q���!�0����L��%*�$�Onh
��	�(�cEozӒ�	��?)b�\�vQP����&�y�`�n�Δ��k4�d��a� �hQ�|��M�m�$���'v(���Fst��� ������(O�M��nA#�(O�5�K<��b��K�X�q,p��	�F?���0�4�O��gT� �pY�f�`u��IIq�H�!f�,��"ƌV�(��5B0OiT���O��HR/Uyk�iͺ��#�<}BU��[�h)*Ox�`w�a�'j��PTŀ�����BHx���p�_t�.������4%�0�'�E��b����E	 5��@� 0^��t���p�����b��d  @�?����  ����(�?k7�_�vߺ���(�,4�� ړ#��E���#��8f
?��z�[��hO�"��'��#|
��4)dġ&��u��)�w Ka�<ق ��X��L����*����pfIX���OF��2�.�*��b�ܪ��IpbP���A���MK��?�(�X���
�O��$�	X��دq�����g��%O�o�0�����u�c�ɹ&29���QfhhYc$N;擉�T!�E�;��8�����ɳ'3<��ᅖS��5����↝s��1Oq����G�4O��B�*���Ȭ1#��OrH��'!T�O?��C��$y�L���'��7�����G�<Y�$����bc`U\���\f�'�"B��^9y�pH���:oy�b�E�B|���'.��K��H����'�2�'���n��i��������C)Y�0v�xs6���Q�(y2ɗ�J�	��?M���'�O�z���i~ȼ���-~SL%��hV��n��;�`ěeD�w��S���BiRC:��R�Tjt�γqV�%q�
�#b=�'��Y1��?a���'y�I��	�m��� 8L3��b'�ۍ\�!�ĎuV@��؈e��i׬�(͛V!5��|����DM>76�\��虽W���0G�w��H��#ހ)�����OR���O�@�;�?�������~�	��V��@�)9b<u�x����gŠ٧hĊ��Or�r� /5R�hu��1�xy��֖)�j�S��Lڤ�2k�"�7R�M��y��UH�,L���LH�? ��{Wn�BJ����u��|�i2"��$�禕"RJo"��`Q��
�nQkc�4D��jscˉ+���J�(ȰIN��%ʳ>I�i��P�Ī6&F�����O��l� �rP � b�|��W���7�ʰX�D�O����y�v���3Q��%�ĭ�8qyܭϧd'X��R�ܢF0�%���)T �E{�BU�!�jT[Ԯ�S>,� ��0�B�-�e�b��)��1�9cў����O ��&���QPb�zM���i�1/#�ꓡ?Q
�H�B��,�$}�P�do�J8̈́�	���D��E,�D(ևY�N�6	@�.p*�I%|�
}Jܴ�?1����)L2A����Oֱ6cIK�2�rH��3��`����mQ�/Yߟ��<���'�hA�J��p	�s���bق��W�vTFx��	��E�� (0�V�$U��I�� tи�$��M8��,2r��fk�]��pFI%s P �ȓl��(Y�؏,zLrS-��?�@�Dz��8�?JtIE�¤:iBىEa_�I��BA�i��'_ٻ�nX�C!��'��'ߊ�]˟�X�����.��}���V�2��6��O�y;�(ס0���=�*Ģ2��*�挣u�Ϙݸ�������a�q΃!c�$��jFp�����kv�1I��ֱ&h-[tR�{��&�' ��:F�'��7�o�,O������J¤G1 pA�_�~�7��#�O��6�Ґ'�p� 
ȁ<7��i"�i>�7�঑&�����?��'P�@�MX)�e���<aS|�2m��1p�i�P�'�2�'�¨c���	��H�':����S=�!B�Ή�f)�D��/� �(�	�aR?r�ܐC5ũ�P]H�I/�7�,p3g�$AS<��G���R<����� t\[�`�J�Z1�g�5Zs��	4c�'-s���1�O�J�C�/m`�Ւ4F,C��5�bo�P�<1C�D�/4\3��Z�)E �'��W�<���5@�	�ɏ��&�@� �Z}��s���O�����g���'i�)�8����pю���	��Y�:Q���.0��'aR&�;0�RY&�>L��z�B�(zeF�S'm�A�PiQ�4xP|9'�;y�0�=A&�U�J�b�kW�E"3N��h�9�ug'7p�W�^|@Ab��
5�����[��t�=A��Of��;�S�'DaRn�?�^5RǤ��FP��p?��+p.|���!C����aF�MX����O���G�$ڂ�����.O%©+�S�$�.�ǟ|���\�O��h���'��O�9W����K�u(v�V/C�r�6�6EŘ��H�r� ՉU�ܛ���O)1��뒄ғ7_�q�"��b�l5@�D�O���`㑌;���O[&��|ݵ�ą��"n�O�p5*@��G��x���86�
���'3��I���䧵�I�O`�%˷��+޹X�Sq� B�I�1����G�1Qi)
��ж�#=Aw�S�|�l��g#��ԙ@�T<>"�Kݴ�?Y��5��"b���?y��?���b���� y��W_��#� |�|�X��!�qՇĢ�����C/���C�'k*0x���J�Ct�meҁ1r�F����,�;J��v�[��Ii�8�ˀ��"��	�D��A��<m*�$����>�Pʓ��D�Od�=��'�B����6Y#N�7���w[����'d� ���G[*f��!Ol_�ɀ۴;呞���'���H��0�;�ϗ9!��	�!X by�HB0�'���'RLk݉�I�ͧHn`��!�3?��=P�h8l!�LҗH�8a��Gϕ������$��O$����&G���b��%<$�����^_Udij5hD6���Ò���X�
7�D0M��	����Xf?)2���P������e���E Z'v����M�'�@Txsb�;$�
�u.tE��'�x�j񯆃�9�蚏��B�O�yo�ӟ��'��B�ϻ~2�����C�"#2���β:�R]��S��M���?����?�v��$f���W %ґIZ�l%��.��FB�:].a���o�ў0���0pSX	�%@�}�,��2�뺣��/N0�W�J�R��t���G��|� ��_�g����Of�>ŉ�KF����T\�#�6�(G��>��m<�J��hf�ЂE �����I�����*��+S��:l�h�R�^F��	�n2�E��ԟ��IG�DF�%C"�'5y��I�Lf��6���fx��%}��up6��!��L�&u�~%��+�O�$�	'Y'��X'5�Y���l�hY���T�ި���]9�l���6�X\w1��%�Γ��S�<�r��O�;��c䫀4(�0�I��~��'��)�I }RnX��dtӤ�Cw PلE��y�JE"��(��� �����m��HO0�F���D�v�A$���g��H�R�V27yt6m�O��dN�9:@0�5&�Of�D�O������d�S�6esW�,,�,]r2�O�2��LS��.@�,I���> L*rk�o��ɀ��u�S�
�"�jA�P!�Ed��Y�Ӭ5�l�A*�%����|"�4k����s�Ks}�]wà1��+�w��E�ۜ��o?9��hO��)� 6)[VL]\�^�0�nۢ6,u;�"On�����Yָ�AD���l!�־i�#=�'�?�,OD���e2"��(�*�C�=K��Ă;�4H��B�O���Oj��������?)�O[0T{vH��\.Aˣ�����l�ꇛ����%6R9�#��џ�:3mQ�l��@��1f� �t.
kˬ����9��Xz`�D�z�im�Z�m8$F?�	��~�Β�N؞��"�:y�@-�P�H$~9�6-)���O\m9�K��Z2�����+tLj1�"OȠy�K�:6�ȭȵ�[6EF�R�Lr�4�?�,O0��M�S�t�'t��w�~Q�ю�"R��Bs
�&�&�U�L+B�'r�N$;���Ud#f��\TĘ���z�,�p�ES�F;��Q+A[Z�=��Я|R\� ��'��{7lܖ�uG��ጰ*�d�/^ ��PјͨR�7��'�`�	�� �}�d�s��H���]���pe}��'�␰��
s̅��J����a�7���-q���v��K��C�!?���1�(�3���?I���i¾^���O���i=�HL�F&��N0�A�q#Ԧ-BR�Z^��ܡ���%^X.p�ю�"��	#�CDp�pQHݷl�,-��.ֲ
��H�I� ����/_+	�����o�<t%pl�;L����
Hf�)Yj�4]�!ܘ	�Ë2 �D�[?Q�������>9�����G�٘X�H��pR0�!�D��) ���H�� ��c(e��ӌ���s��p��P�?цT���܂a�2�o�4��eȦL��U�������?a�I�=8��GSJ
�3�MX�M{BXp��[�(T"��d���������>�xd(\�D��e��Y��ǥd��D$�z��!��˚*N@*b�q��i.0��2%ލ��E�1:��q�NU�?X���l��J��	��~B�'ў��p+:a���"i:�N�U��ɇ�&��f�2*�Ш�Pn��o�&EoZ��HO�I�O�ʓ��e`D��=�t$�E��2OT��s�N<�H-Y���?���?�E������O�瓯&��׏
��sӤI1�� "�I� !3����I�!B$y�,F8b�џ����=&���r�
)y	��U"Ǽ%�]	%��=�F �b�gDrn,�BͲ�'6���~RYIVh{���+��8l�"Urtnv�'�Q���$�ș?I2Yp���6�R�y�C0D��C��0G����׎J"US�h�>���i�BU�,ȳ"B,��)�O����\��U@sJ�mÈ@`6k�"s\�7-G�5el�d�O���ɣ͠x*PX�L���Γ�r���Χg:��X��+\f-�dʝ$�x$G{�	�[MJ�;�̀cg���`�D ��U�Ex"��	^�r�(�7�ڛ��Z��̠�qO~!��?��.1xx#2k�"s&x��G�[���$;�O����mϲr��M�d��K\x����'hF�=�$���+�)+f�񒆡�@��'p����w����OZ�'uZt0��?�#�O*�$)���:���9
K$�樍�����+�hib)������O*�U�t�O�ab���4��4$0���'�$�9%&�|>` �N>@��wKCSbLE�C�;G��-5�TyP� �i&�����(}��I7���PM�)�'I�QQ׀�$r"4�0&
(.b�k�'��2����bUHp��9U-���}��'�V"=�'C�(,�V��U��D"e�N�zջi���'����6^���'gr�'���]���P�X���<e+W.�t/.p�c�	#X~ �K^2F�n�x��H�uW0�fy�׫ܢ�ēp�^	�&J�F�BY��ʊ9����H^ֆ�ht+�/:�r����A��eܭb�6 &�T�+�(P�P�F�)S �h�D�<y�B�۟ Jӓi#~�T���%؜}a���u���ȓ#K|3�A��b@1tI<-��n=�HO�i3�$��}u�xp �P�&�)F��gW4���-~��$�O�D�O6����?Y����ͥڜ�T�ٝ�48���M'�� ���lRؕ����a����7� Dy��^R�H5ig\Y�����f tak�!ϚY����`�X#���<r,DyRGB��?��A� �,��B0;=���f�+1�!��c谋t�ȻZQ"�.�	�!��HB�}3�u��pR�Kf��I.�M[O>i@nM��������'r����'�Q�>�q�h�6Ì�nڗZ�� �I�����5y����V���M#Ԩ� �ծcn�j�O@&V�xS��#)�)T`�D ���ƈ0�^����Ҝ�*��u�p�2dYlѲ/��y����qa��=!�֟���]�'�܈�F�H*;8h0�"��;ȭ��'P2�'��-��J�6d�R"$�=s0aR��	_��ͫ&o��	�yD��P{�� C"���i���'��S��
��I۟�ڷ&O�c
jxb5#����.Q��M�A)͑x����R��t��J�#C.���Ļc�Ex���K4P !ȰL ��N8 ЗG�!(��#�4h���鉌Q�fI�b�Y�' $Ădg�����V)g��'��)�i�O\��
�*�
≎$ kP*j��B�)� �9�lB�	��P@�9d�Q����ȟ�!�u��D0�g�ip�t�������	͟�����'�z��������Ο��\w?�� 3�
�Ru�W�hP��G\$7����KM4o�yYr��Y��A��|r����"u �P��ϩ_B$�����<T���G�E�:ت���0xn^�S�T>)�P:�	/Ѐ�$�є;�(��E�� ���DP���	ן���u����$B��9�Lб�䔩	�F%�jւ�y��
8��j&��y��A�Ӌ�M��i>���Ly2�0D	Ʌ*�4�$k1�A5U���r��Y/^�R�'Mb�'W֝蟼�I�|�5M�.21�R
�nQ�	н2���6k�`�8#�݋v�� ��~<��/k� @	p�ٶ	��2b]�I�`�&ź5R������#<�g �2pd���'P i�a�Q��G�,��@�V [.69�x�&"O�E��(�T"b�C���8P� �d"O���1��)Hlj��p�L�^L��K�[���ܴ��Vv�3�ir�'���G�G��s�ʤ�\AIR�@$L��6'؀ByR�')�ؔ|��)u!�od���"�H��I�t U!XyxUK��#y�bE�'�䨓��F!eX�y���3�X{Ŝ=�:�R���e3�֓&Z�X�'��8�Uꕠ4�]J���������2ټ�^UQ�Γ�[�	0"O��6`ϓ(��)���A�05���'|��-`�T�$)K�E:8���'jd�Uy�X���O��'?[,����?!�`?W8,���ျ\�!J1��,6p����$�Ԝxe$gӘR�m�Ŧ��O>�S�?7m�0�I��c,F���.�u=R�WYB���!���Q����RI9�d�0"'u��Ѕ���Z2��p���,_�X�C�k�O�!a�'Z^6�����Ia����6݀����zD�'��(o����?����?-O��$�O���D�d�0ljl�F���[O�f� |c�^�=&���I��	�<����#X� X� ��EBh�rkХ����'���*�L�T�'?��'�Z�.�Od8`b�I�vS|�aю, 0�(K!kQ<&�@�m�/E2%�4�WE�-�\wN">�A��� a$��6h�`����=-`��x�M�Eь- �J6)&^H�O�E���@�@T�'�>\�c� q@�1�0 g�\a/O��A�'P�6�BX�IƟ���O?��a�>�	T�� d�`��w�TR}r�'YR�|��IZ�LV����h����l���Y/�&)�O6m%�d������<��ƨCW	�N��k	�@��J
Z.�0���^�?9��?!��6�n�O���w>�� &�<d�9�!b���T���K�j���E�Lf�)z�ہ�����N 
h�Q���eN@4F"�s� ] TC�fF�!AcHwT��sV$/~@�du�P��Q�����O��۵��(,���ߒfu|�3�
�i�<Y��_tPl� �br�`{$.�b�<1㚲`R�
D4k􄸛f�Y^}b�jӶ�O���[զE�Iޟ���s.�`J%�U�t��m��fݭ*�mZ�(V�����,�I�����Ii�S��d�9D�{�͘<Y���''�I�'`�������n���K"%�1F�Ҹ��h�ў(Df�O�(�'i`��K��%*�5�c�"D���	.�Cw��,���ڄ�\W���	���D��~�h�a#��a���V�@�y��	�8�����G�D����\�ttR"=q��'m�
��	Ҩ=���<��'L�V��=0d#��=�P�A�y�<	@��&8�XDR�0�
��t�<��Z�]Uh���D�cC�}k���q�<����5L-��+�S@^��aFe�<�&/�9 ���1#�Dg�d˰đI�<I�e�	l)6	H�I�
�4����C�<�'6����և�/�����A�<q4��<��E��@��\'�0Qu�C�<��ׅY}�e�d��=8D,ї)]�<Q�̳(�2U�ȯ$����o�O�<A�N�y��A�3a)z�Ht�c�<�CH �1���"1T��V��|�<q��͂QZ��X�c�fo��c��{�<�����|&����	��{s�w�<� J��Ơ��
ݽ1*ư�BRy�<1楈����X�<�r��4��8!�ON�qĮ�h����K)&�!�-=|�����|^%2�J�!�d����ۓ�KPRu0�JT�T�!�$CL4l��4m׎Cbz�ç�!��1��<�Vo�X�����0�!�� �5�g�f<P���R/]�P#0"OZMQcI�nK:q���T��h�"O`�Rg�L'y�P iue��� ��"O�EQ�)<i��v%/���C"O(�� ��N���K�h�����"O���X�~�iG�� i���"OPYp�ҙ�~0Q����"�>��"O�`ro�r)�$�2�O@���"O�8� �:	�4eل��Q��h"O�%õg���f��c�=�Ft��"OB [�i�,.W.%YZr2���"OZ�K�(��9�&K�z��k�"Ox�`��ʒeT�a�p�]5-=zE�G"O���'O �I]�LC���6	1�5"Q"OZh���s��Ia�O	@ t�*P"O�\ATeҹ1ИKӍQ�.um@e"O����È=S>4xCgG�b�����"O *)��jybmH�+ŧ�]�"O���7�Ղ*�5�� �!��*"O�<SR�JB��݉PD�(��m{E"O~���)�>w�("1�ʑV��Y��"O��t�CG4��d^7LD
Y��"OF٪@g˞-2��3c���c�:���"Ofx�	�&O%4����F�#�`u�"O�i�e/eU딡
�$|��"O2X)���W��$��I�m��	z"ODh[�� �O��Lp��Ć�y�[�b�'�o)�u�t&L4�y�؀&�z����;cx$Z�b�}�<q����F�$A:��3Yf:D��-�s�<����n��Y�ď]�x���K�<�  �8Ge�Ԋ��%��e�jD�<y��ܸ_���
s	
:tv$
r�Lv�<�J�˜�r� :̼�[�.�O�<A�
�7�
I��eN%���;f��H�<a�kİ]�O�r�z!1��_�<�4��7߾�8eD������X�<٤�C#h�;�`��Up���B��<�Q�CS���9(�RY���u�<�"� I�YVJ������Cs�<� �˧A�&0�S�V"��xJ���c�<��`�5�����Ɨ 2b��I�<!sȏ�R��� Xwa&��bG�l�<y�ȶB�P��L
�{:�H!� �`�<q�@9D��!�3��
�X�#�y�<� i�9ص��B��@�רOa�<�wl#.N�A�.��om�pjAy�<!a��1V���3�	�����@�<Y�Ì-��I�� \�� Y� K�Y�<�6ΐ�Y�i�4�Q�=������L�<��"T8]���(V␴B>�]�f�s�<��Ǔ�3�|U����^ꙙeG�<�JZ.f4I(db -sp�q$�CB�<iԋ�!HQHT����7Xh�`�w�<y� @�ԁ�`CH���B�z�<�����Dӣ��8xz�M�w�<i�U�O8��x�oӈVf0�A-�N�<I�)�(Pp��p��}1�6��p�<9%D,yPdx��ϠfeZX ��J�<@!�sBX�P��Z��=C-�G�<��N\�;p�a����X}�L֋�~�<!�.�0OI��a5�*��	H��v�<ٕ���s��g`ͱ>�
Mp��s�<A"$���p��G�|^�i��c�O�<� �<ZG�+>yhl��9�N)�s"OP�������������"O:6O�>B�Ȼ���f|&8kA&D�t���_m(F|�r$=G��t9 �$D���"�-w�n�f��LY�1h��.D�|�G�ҧ:���3
��^6�B�.D�X(E�g�D�J���{������-D���E�T	��<�֦HajҵiO(D�i��W0EЄ�,ՍU���G1D�@�)_�vo�Q:�X�i!~����$D��A����K�i�9�@���P�<���Ȏ79X�bJ!z�$��@n�<�f]w�0�`��\�1���a�<�C�C��R�2foDIlnAJr��~�<�E���8%� 5��1�����<�c�@"��4}�����*��<� ��k<z�26n�	|̬��*�x�<�Wf�!{�h8�$�a$xrmCI�<�T���0Ծi�m��>q^p�p�B�<9p��'q�ִ�#��)H\�HA��]�<�� eW������Z�P�c���c�<�R+	����0�Un��>�.H�"OR-3tfΒ�xc�#\�	�k�"O�a���B�L9��`��ɰ�f"O�L!�k�-Y��A� �^4HPq4"Otܱ���i�I�0)
�� �"OB����&n�:���P����"O���@Fg�F�Ћ�2dZ�i�"OR�PQؑjP���jT��� ��H�<�'�� VQ8cE��W2���UN�j�<I��t�A��Q�7�>�z1��i�<ᐣ�"�&��KəL:zm:eCWO�<A��A�\�va D��]�L����t�<��#T'Z͎1�6��t�J�"�N�M�<�#�0lqb��J�r 3���G�<Qh�#��HA�"U�'� ���F�<q����	�Jp*���	�ĊrFA�<!6AѦt21Q�#׏e�-��G�<9��X�5XQ�N�%�( �e�y�<��ѷF��0�U��
x���Z�<Q��T'Bc���.P� ~e�A!V�<��<�J���j�u>�<��o�<�e�M�Z�5q��FN�� r�<�a��x!��c1���6��.'!�L�[�2]��
�\&4L�#�3m!�I�6�����O��cĤ��W�!�dC�Μ��	9�$��U�{9!��&E7Z������$�$Te��}A!���<*!�,if��D1��c���~�!�J1h�L+�j��{2��P�M�!�!�dS������!k��J�o@�7!���x�ڑ�'�W�GLе��m�?*4!��Z�R���įGd	�鑺4�!�5q����`b���c�$Y�!�dܵH�Z��
62��b�3�!��&9�)3�D�� �0'l�!�Đ0U$����Ս�Fp)EO�BG!�d�'v,��"�GA����*�d�!}C!��OGA:�����{@"�"�9,O��d�;]"��f��QMF��O��y� 5!4�m�4kُH|��r�끇�y�H݅oy�Q�R\$yi�|��.�yn��w�ze�b�]���'LM��yòN��$J#]H���)�y
� �t{�`��;Tք˲	G'rN�eK"O�� ���n�^�%�@�~��|1�"O����׊*�Z�k5��#�����"O��їFW648j����4 �M��"O|�#Sk�>و *A$�$j(��"O.�$G��PA�`�)�d,I%"OZ����Nu�$h7��7G&�p"O�*�đ$1�Y0ϒ.dJ.��"O$5��N^Z0	�4��C����"ON�PaeŶ4p��s�^�4����"O���vn�(��C��4���`U"OF�9��"M��2'��LQ�"O��0V��||}��_�E}���F"O�APEA��q,2A���r`���f"O���� �L��3�ݼoYND�F"O
���	�W�vlɃ/��vO�`3�"OD����0�|X T�O6LHY��"O��;�'H9x�Q�vo��q��� @"Od�'��y�i�`�/~8H���"O���KCc����*���"O��Č�U���Ҷ+@j�P@r"O�|{�L�o��	�S��\e�إ"O�y��	=���$�/��1a6"OQYq��t����JC='�
�@v"O���/�� ���@�2L����D"O���!	&)DR(����#X��"1"OTu�  �!1 0(U,�lu\�H�*O&�S�`2H!.m	���,���P
�'O��
���<���{p#
�rq���'AD�#�I�G`N��$I�c��U9�'�Ҥ�S���3&`0�g@<�YB
�'���M�*&�U��%�|���'�ָ�pc�F ��"�X��!��'5�Q�u)�F(�ˡl	�(4�
�'��Ar�J�#c<�Y�ŵ랰[	�'�(4eE�q�f�r5&̽O	�X�'c�Yp��;�
LBF�K I8Ԅ�	�'�l���.Y�= <�"�&7�����'�ti�����Vl�`#�U-��x"�'�H�{�����u,��ƀ��'��D���n=�\��Hfٮ`�
�'��<e*G�,��5���I2
:%��'Т�*Ӌ_�<�^pSCiV�&<Nx�'�,��a���8�v�J���?.���b�'d����N����S���Q+����'�hA(7�։O�8Z��ɪfhYz}r��%� �K^%c�Rm����HO��A��ɿ~��킊E\mB"O�t8!
�,[�B-�"��
M@|��"O@���I�8Y��5�G�#�"OłF��4]�<y:�B2h��4"Oj@2� ��c���M?"�L"O`4��aU���!!ѦI)5"O�q:����&����+��A��"OD�¦�~z�tY� бr�z�""ORY��k<��HD�C1[�!��"O�Ux��@2G��aH
���"O����ȱP�6�3��&*��EkF"O|�A	���qWiÙ]�ș�Q"Ol]I!̉*o�XK
��d��"OV�9���")̐S 2[��dxR"Ox1�p��'t�Z�b��M7�]��"O�L���� `��(h�I�p��H�"O<�c��Ap�]s.X�k���s�"Or�pJނ.Zb� ����"O� ��{(\'M�,�sA ԟ6���"ONXQ�BZ�G���`@�Q*\\��"O���e�ѡ|p�y�N�G���"OT�gһ*�b `D�%A4�+F"O�1�5M�#w�Q���1���"O6)��hѨ7�Z)��S�ht�"ONb��_/Z,�P� �90��7"O�)�Tϵv�f�QA@�4.�� �"O� �,ޭ&�������"*�r�"O��[�$��� P���`hf��2"O��a2�G'8e.`�ƹva6(�"O�ٻAMj�y0!l�wL�d"O�]C�A���T�;�öK_tI"O�̳��CuVDYeW�:���"O� f�I+s',��qKE*�d�s�"O�,Au�U�f��Zg�S�v`�H��"O�z��ʳV{�|�6�]jV��a�"O2��"N�����`=L\R�"Ol�"scL��({�	�6]5Hț�"O��H�f�^Ny�&B ?��E�D"O,%����Kc�a����)6��D��"O8B��˪9HƼ3��� ��\��"OJa9��״3�J�xjT�"O���r����#	�qJ|�y#*O��{�Oǝt��ĨεrwpIk�'�<X�! ��V[��K�e��@`	�'-xp�����b��B�.��i�	�'������=8�؛�mǾ�bC	�'���S*Y4\�"��
���@	�'�``��-�0�:�2�9�8��'x������7oN�
�,�6Q��0��'�&����_�s�L��pC�P6X���' �"��g�l�2���5?�	�'�Z!#pdP	Έ<��Y�b!�ո�'� ���6^��)`�,)��Q��'x\� ����D�
�(؂3ߨ���'��)���Ѡ8�x�䋀%5���'3te���+C���Q�+��DPJ�'�:0��/Y���`*��.8�'�I�u,�h`ޭ M���h�
�',5��o�7^��zhC�	+��
�'&\�ᕍRR�a�E�F���
�'�n��`�N��P�weHl
��
�'�b�z2$OnS�Z2�+6�HM�	�'�j!ʠ�AF�xl{P�E-c�D0`�'�Y�F�['NL~i�@�iĩ��'�<�3�@˚jP�!O��_�r!;�'����V�&bѠ���"O'JPY��'��(A��Z��DT�Q�3I�yx
�'���P�Ě5`�8B�K�-b]z�a
�'�nܳS�Z=PX9����&L�}8	�'�̑s`E�`#�1��+E�PLXd�'��0`b�R :p$��%KJ����'CD�#v`�¨л��نr}.��'̒P�A��[پ��a��x�N�K�'�4�p�]0��hf�'8�瓪ē��ܫf'�%h&��F�ӏ2��}�ȓG���j�9p2�0��@�z�Fx��)"�k�O�(����.O�lHEJg�<elC�s�z�1�HT(Q���#c�=�(O,HF��O!����}�Au�U�r�4y�%"O�c�38�� �合Y�n�`�i?��^��]+%����XՃ
iO!�$Y�Jp����P5}�n\��c�"@�!�� �����4⌁�j�!PM�*�"O -�����T���Q@L�<b1�"Ov�[�d�56߈�P�(��	�X�@"Ol-�g���%�x�*�] �r�rA"O�1��B��b8X�h�<�*1:"O�Y�
��n���s�Q��d���"OBI�w)	q���jAG�\��"O�e�2�C+9v�pdʽlL�G"O~��e��1�VE*p�L���}��"O����p߮d04#�G�ĥx�"O���R���J&t��o�~��,�""O�����A��q�0�W!\��$��"O���� �r���4Wy��s�"OԠb���C� Ȓ��Y�!�"OJ��%��8�����[	0�1hS"O�$�B U�Y�2�Dlά�"OHeeE� ��0r�-�zx<t�p"O0e��jݤA���R`�	5yR5�"O ͚��V�^���F��h�Mbd"O����E�.�L�!��f�M"O䀒�*@�!O�(Zs
[�G. yW"OT1!��o��"#�+ܲA�"O�|I��~�~eZҢŁ.Ȓڔ"Ob�����`Fn�0P⍞����"O��v�C>i�p7��8wi^1Ja"O�������D
�d�S;:i�D"O[U���i�J�Ra䞓K;���0�'}(�&��" ����"F�h�x��/D��ʇ�ա!5�U"+��O\v䪁#.�I�1��"<%>����[5j�TD0���/�!��+D�TAGo�=I:��4B��0�QU��G��OT�G��O����� 9*0 �)ߞ<%�@K�"O�8S@���R�D���'���[��i}8t1��'�B��iY�}� S��Hq#dUp
�_�@H��"6�W�n����I�RyF�ۣ�%D���%L7|x�x�K��;؂غ��$�I�φ}�?%>� �Eu/��p��L\�z-$D�,���W�ؼ�V�CU� �!��DQ�'��D�,OL�#u�� AQ�,��.����E��"O�c2&��2�&0���ٞg� Q��iB�	�)�~IP�W�NLz��1ș�UT�C�Ʉ�0b�b�3j���B�+� �`B�I!W�-(ŧ܂P�\8y7��32�c�����)�	��mPe��^����P� �]�!�/lT`�PN�=cEj�@�oS)�����DF|�����6�����z�r؁�n@8�!��"�a����tX��"Ԏ��*��f���������
��rF���c؄?�l���g~�M `��	���F�8�yR..8CA�&�Ͱe�V4����y2 F��f���L R����,���y���+d��9r��MH�-��J���y��=���C
�I�`�t�J>�yBj�W�b��Q�қ1C<A�3�S3�y�m��|�>�#7%�d�g>�yrE�/4�6`u ���t #��y�k����h)d��,ƄK����y�@� $����F�W����"��$�y2 ��V���!G�Hv� �a�T��ye�PV�P`��5qQ6eʑk��y�O�%��KծG�kĔy[�$��y��/T1|Qz[���C�88�h��'� 9�F-�C��5���)�H�	�'!b�1��I$1�,�s`�ʨKXX��� �11�M1݂D�ރw#���"O
��.�!:8�'/L�c�^�p"O@�+�Q���0�`k�F��r"O̰��o2j&�x��L]����J`"O&t���M��z��B�*��I�"O[aօQ*.𬈦)�1����$"O�q%�:ۄ����.�ѣ�"O(u��a� 9���X��6B�� �"O�ӃaL�^ĥ���]8A]L�s"O� � ԟ����`�V`��PW"O\U�JJ)`�TfV�=^�K�"O$�� 
�$��U�$ݻ����"OB��FQ9�f�8������yR�"O�������8�8}[��E�\S��p0"OX��`�S�^�c�G*,6f���"O�r#�6���#���w%)Be"O\)[�/�Z��� #&ߏ^�d"O&� #�* i�l8���C�r�Y�"Op9 $L^��CJ �c|��"OVuѥ��7!���p�ŝa�r�""O��@��
�Q��=�Cً&+ �B"O��
7�[.V0Q�Õ.Qs��
�"O��$�+�H�6$@�X�Xb�"O\i�t&P��8D�#R	_���ڐ"O>�0N�i��11��	2}*ݺc"O�e���� }
l�p �e���"O�I��Ъ�Ґ�NhJ�S�"O��p�Ҥa�,吖n�B� ۴"O�#�,�:]�$A�-�<LhD��"OH$ �)��]�1LH���pU"O^| G	ؠ&�ہ�^�-*A��"Ota�$ID�S�R<��Hӻ7�n� a"OP����7N"�he��){}��˲"OI���H�&+���`�R*�G�<9p�L�I�7Iu�l�2AWl�<���0C� `���>X�*m�<ق�\��*0��;�X3��d�<�FIد��s1��[��%sG%H^�<�So�7�4"�)��d�aY�]�<I���E��	Al^#B���	�s�<ٳ�K�.0�*%Ŏ2�P&�R{�<�b,Jh�V�ڐu�F��q'MP�<�`��!��%I��ƘN�t� f�I�<y�� =.d,AwET�T�����HSa�<a�n�f|Ab�H��n$�A@a�<i�ԅm��%)ckN�u�V	ڢNc�<)PlM,�b	�&�[=3����`E`�<�w��7��4(�6]�v��ՇNZ�<	�����$��Ĩ�(j��C�J�@�<���u�V�(���5��@#Kt�<Qv��&   �   !   Ĵ���	��Z���)I x���C���NNT�D��e�2Tx��ƕ	#��4"�V���$U*��mZ�ar��C�.F�~͢�^�ew`X�g�:;�i��W��M�r����.��h��Hn�+a�'�
��dg��9\�����+D�� �skh���PyBB�/.��E`.}lȤBY�Q��J��q-��M��R9����'����  Dn�T�.Ob�-b�$�Z��F�����K�yQ��J\�؂�܅Hy<3�L�-����OZڇD��
�'���;�%)�P�
U��]����G#ڐ������>Yp�&�|9!�>!�!V�6Q��B�'�>=�0�
�L��m���e�	��'���	�OȤ#n��c/O�@��#K�,��'��A��k���k
�(�� ����l	��N<����
���P��M��â	�3�u���n�}��d4s�"O�I�4�Ƞ@��'m�Mȧ�H4��F-_ԣ�ʝ�,��`I���h{��Q�|���'��	mǦ�H�^�TΓE�v%Pw����(�Ӏ�9\ަ`3��C~xu���'!~�D_�<���hgU>�	#S0�QJ�~���x���چP�d�A�!p^�RV�~�N�����H$ ��<y5�'��,8V�I�8��$�˦�h��O4?���@�/N�B��4H�J
/� ��1��$��C�ß<�u��:ʛ�4O�U�I]���ж�Ԃ!��DcW��{��`�nԕa��'�ڥ!D����}��	��<��cؽNm����x��{D�	Tyr)W0`L8Dy2�A|≓k
�����o����ω|���ɓ�xzb�xP��A�M\�=��J&!ܟ[�� 
�`�g�0��s��.l��i�Q+�`�M�|��Џ(��$���'j^s2��3z�<y��X�A�.O�I��W���'S��:B�,�ēe��[#�, !��	�(6���EfS2^�&�T2�* �b��Y��(�d@baE
Y!�Ժ1MQ�z>&̆ȓ'�}   @�?��f�5bS��[����0� �ؤ"O��8֬�`N�
�	۫y�.D�q"O��3:�U�`+ ��I�"Ol��ɨNf����S�L�m��"O���	 �h�L�,��dW����"O8�a�N¹!����#��<�!�"O��Ɂ���
3����k��I4� ��*O�!��*Y$<����D`�����I�'0�m�Z+vcB\ztA�:R�(�'�� 8s
�z�t����ؼ���'�Yڡ&�=x�"�Ox�X�:
�'A��e��?\��ܙ&\7x_�X�'�
��A��P��}X�:vIn�C�'� tR6�QIN�Ӷf��l�L��	�'�|�1���j#䝣֮�3h����'}0|��ˆ`
h��Ԧ� `l��'�Ni	bW=!�f��+�^�R�'�
�i"��#2m|�SOٵaϚ�
�' �$	c�
(��K�V����	�'PZ�I7o]�h첣EM(9 ���	�'�W-�<��ACi�3%��R�'���b��5��Z�í2t2x�'5̐���S$����ʾX�Vic�'=*蘠G�5f��hEnN���p�'j96�� )" ��圔YV���'�j��aj���x<���ԡ@�8�Y�'���
�́t3*$:�GS6�^�Z�'�V!�%��3��i���L�X+>5S�'���P�жK���aR-` +�'ڴ��5i�U�����!�!G�<;�'�v��׈���(�*M.A8���'q�4HR�X�Ybd���l��9�Z	��'�`�8���	����r�߳"��L��Z��9#�Ȏ�����
/m^y��}f��v�Ģ]�aYc��_��؆�pn��6	��MLĻ� A�/�t��ȓM[<����<��,yB�ܾ,S����b�@ը�[�L�0���]�2��ȓ
�^�1�
	3XL����*�np�ȓ��y���ɰ!�U��������	�@����*1���l�8p��6�n ����oKn}���E�w��h�ȓu7ڰ2F��|���y!H͊0�ȆȓN52pR�c�n$�<˵m<DK����O�~`�h�8������d��,�ȓu� �� @�?      Ĵ���	��Z�zt	;A���C���NNT�D��e�2Tx��ƕ	#��4"�V���i��mZ8|l���Ҋk�Ĵ�����'�4�q��*�*-��i�#�M�2$'A8�.�s�i��GI�q!�'W�<������*H�$��FU�\�>��dyB+z��hA�C&}"
Z������e�|��RT��]�h�Z�x�'N�)J�`"8Y*O�P�c�٣��cV��
��	�Y�85��]Zʭ�1�
�U�V�!�0��Ъ&��9��|ri̤,���'�B 	�ƅ�g�Q&#��O�t�	�Z��@ゎ;�$�$4��i+�O�L��G�h��������
���~b	^�4<\t��x�g]XB�R���$ �[2���!
�;x����םTw�}�Ï���U��u{����P>� &�a�m(��0�!�5XRt�#�g��X�c|¡̑`²D�N>��m�cˎ<�'hB\��
�	RmA�-�p��2G��p�@R� ������tf�"�ē2�pp/[11F�-�OS!x�\)�!�E��O�k�i��|��w��Qܴ�������"4i��EJ�D��D�'��4�u(
���'x�s���(=�_Ħ��P	ΔF��P�q$^����D�;#��C֬%F��Fߟ(	�C�6Cԛ�3O����?�蘡J����剄�a���e���M>a�Eʢ���$� GGɫ_��牅X��(!�KH�]�4<�10]2�ʓ)N�!R �:ʓz0TOT���b��3��
�/Rs� �r��O��Y���Z?�ē�~�B1m��I��5w��q�e�֞Zn�\�4>� ��.�'D��c��S�s�j��N-;t�'J6"�.T�'E�P��-�Q�F!��I�=6�I�7�|��	44�)"O<�W�Xm�����aG�v	��(�GQ�R�ꁘ�Ϝj��	&���?�I2{� �C ߢw;9�"��E��Q �Up�<��& 2  ������:!��'
� �  �痨[�C���;�l���'��tz��ƭX��*���8�U��'��a2�o����h���3^A2�'ɖ<��NڃS�\�Q�Ę+�q!�'�P-���� VJ���Ƃ&D��`�4��D;�)��MY�j֨��@\�-�D����y�KL5`/L��v/э��2%��yR/X�F�F���ɾ�,)�Q�X��y��E1}V��/˨h�)hQ蒣�y
� �mÒ�j�����6���&"O��f�+$ҺA�%A0�Ԝp�"O����N+�}����7��I�"O�|J�d:ҔaVC���ig"OP@A���]o@x���B,b,��1"OF� ۡ:N���n44!p]�6"O�$a�&]�x��
�6z)v�"OV�r#ִ������\���y�"O�U#�j��W�l�D � c����6"O6A��L�'��U�w�-Q���j�"O��8��-_p���b���7�4!�0"O�i�h�p���!�v����p"O,5�1GٺO5�d�#ӓ"�����'��	N��O5����%��+0�^��!�D�/Z��!sSS�+�&9���՚``�d����=A��$��o�P�P4��3r琽Ô�ؙK�!�$W?8(Zu�<s��a���S�!�L78"
�i��I�gL���6K�c>!�d�DQ�,���(-"b�"e*�,4!�$�3	�Z �T���*L#��\�*!�ă�Y{d܈Ǧ�
s	�͉4'�o!��<���a�L�l������nayb��'h��0Q�5�����߯�C�	�l���ԁ0�%�B�|�xC䉋�&=9��o��M���X�DGl��$.�����-� �n��F�nU�0�ȓJĖP(�W7��q�k�&�����~"��J�X1�Ǭ�?3d2���y���	L�J �Ø^ޑ���L	�y"'�%`B@��� [;� �Ņ���yR�K�_D��Z����|��ٸCN�,�yk�"�V�3�c�3q�}*F'�	�y�Ő�<�*�"&�S�r7����j�8��'L�z��ɳ<��бa��9�X�s�jϝ�yRe��9[`��穂�[��j'����y2h^ -���Y�/ʖL��0�N�y�G?&͂�a���q����E!��yr�;�-I�"@�u��p���/�y��T+&Zڌ	f�� g��(�C��-��Ov➬�O��x�a	�C���vH�5,�	q�'�d�r �~��������h�����7}�;8�(PC5�p���1�E�y2Æ�[�)��ɏa��$�P���yR���7���:���0`栠'�P1�'��S&�<@4��R��bIxa�'�z�b K��4M�%�ȰaRn�Q�'|x���T�X�
�̔�]�f�X�'P��Y�B�$jA�-q��(� ��'�����"эB��u���)���r	�'m�����_�k�.@z��
8([:�	�'j�G \F�L �Cc�+/f�p	�'KT��cֶ"����ĪĖ#� ��'�$�ڂ��<JKL�j1(�"�����'�| ��Z
^��'�B2O��H�	�'B��jK�\d���j�Hr���	�'%���Ѫ�����3��#=��e2�'&��Y�J�P;P�`s��'ބ�0�'�f@��1��D�BC�	'u���'�n�k�mYR֢���il��h�'���3��K)V��2��"g/�p��'m�)��CߌXh���!���v�`���'%v�Z@�Ć~�Z\y�bA�]�
iZ�'0r���B�M�@��-��]@45�'(��iVl�b!�#��O<������ ����j�I�,hх�0Q�����"O�t
V2���� ���a�"O�	�s�
2y���z�(8P����0"O��G\[�%Q�菶C����"ON%�!#'�&�(� �g*lx�&"O�]	7� �V�pa1��o���"OF�k�i4���/������"O���Mֶ:� ,����%R�2��"O�yR��^W��`��+�7x�.`c�"O Pa��Kk>m�$IW��Ca"Oj���	(>��d����<	�"O��狨9��-�������r *O���G�X�j�$ �`�W�[ V��
�'l�)�"��.9�']�TX��	�'�b5�w,�S�V!2�a��S���	�'�Lxa�$mJ$0��/�� ��BU<���� ���\��)D��!��TG�y:�(ú}��)7�)D�X�âG����$�߷DuLY��(D�`�2d��g$���7��*��I��.!D��Ȓ�Ɗf�0��дR���HGH,D����ӏ@���� �U|H@�`-*D�������8���+S0�p�G;D����]�`��r��RD���B8D��ɄD(����DP����6D��j�E�k�(�c�L.��v,3D��P5�%�\a���fK �q�`<D��W-��}��2�O�H � ��8D������0)"�hqI�%2@�q+do8D���F=,W�A�Aȹz����%F6D���,O� �(�"j�3�pK�(D��sq@L�d4T�˲���@.d�d�&D��Q�N�jR��`�A�9��-s��:D���F�Y/d�����=9F���9D��9fg� -n��E@�e�:E�!�4D�4Kw햹iH�Q����0Nj�)��2D�������n�aD+Z4 s�a�D`1D���e�B�Z��4�
2H`�VN.D���sI�w�j�D�\U �R��-D���E _�R^*�`R�:g[�s�i8D�@g"Ŭ<����v_�D[�:D�h��l��3�Mb�@S�"�puh9D�4��FF�1H���#���/��ٻE�1D���"Yg��i抓�(" ����,D��+���no�!;g��7]��
�,D��P�=���QFa٘"Θ�0�+D����M�;����$�ջ#>��Y��(D�<�� ��
�j���^[��d8$�(D�T�F��3B�Ѐ�T�^@D��Hc�#D�h��h��vpn�3��]";��5�QN7D�<X�	�Y��i��/��h/����!D��R&�(��aHעC>��؁	?D��+��"�eysE�Aq:Y�A;D�P��J>B���M�RE� �6D�0�g�J-i������q��0D��z��E�Gt�8�!��j�Ű�j(D���P�[�h�"��*��V���(D�hH �){]�@�^ f�i�w�R�<1[
�.B�#\�0l�05m
w�<�W ůM%��"G����0��p�<	Ċd&��◈·^qH�)�HWi�<��9M��):�A�>����h�<�vƚ �2(z�,�32�,}�5jK_�<	#W�V�X�A���q�Pa���C�<� PY!���$�Zyb1��67"A��"OZ�R�mH�"��ȱ�Y*��p�"O\i$�g�]0�e�JrPa"O��Qׂz�(����1m�ēU"O�@��'֖z�ʙ��!�,D�e��"O��@�
/)��K�/ק@��c�"O�u��GO�-����� �	h�"O�$��&�i�~aD�S$HN�
r"O�q����U��sg�@��S"Om�͂:2���G&"_�P0�"O �Ȓ�n�X����@f|�D"OH	h&�E�l�
qCp	c�i5�A.�y�B�.�7�P�r������yR�J5MR�D�G���q�x�EJ��yb�?u> #�A�2(�i��ܑ�y�임D�x���śx�J�S��&�y����7�,�۵I�%m儰 'Y>�y�fS/�<���@���da�N��yr�D�j2D�!&>\��W!�&�y�f���L�5��;��2�H /�y"ċ�18Ms$�E!	�$%�f�˙�y��9xH|%iJ�j���A�'t��!��ݱU�q�v�R=4����'?0i6C�r��!���H28v�r�'@���Vj�ҐB�r�u��'��b$FV�z��P�Ş�N\��'F>\�,K'r�H�T%�5�X[�'����0'DO����;^D�1����?����]�9��7kI�2�����ؤq��?k��t �
 `!�$H�%��Z֢��#b��#	�b�!��q�h 2��/N���P��$7�!�Ϙq[�]��P�2A�>�!�D3<7�<��/�
d�PM�� �f�!�d5=tH�`N,��u��]�R�!�;1l�
�g��v�iwf�5�!��9xY��97n�}���F�4n�!��G϶H��o�pkHZ d�0DL!�Ӊ)��� �(V�8��G
ʘD!�ć27y���<u"eఫ�/[L!�D���)��F%'�@x���(4%!�Dͬ[ ����B�5� ��b�E(+!��[�Y�R����?wh�p� =!�$K�]*�U�@�a`mkVg�3k!�Q�TG�9R��7͐dgN�6�!�Dãw��is�,)p#V��@��;�!�Y�^U��ʥ̒3���v��g�!�͂@�@��t!�d�R�#���@�!�d��:(N �4ZV|蘗LE�8O!�D�pq����mN*~�����j\!�$^6rՔaq��ƴS�
Ձ��̴H%!�$]*9�];������2D׿/!��֧<��7
��)oB�# Ň�f!�$ۛr���0���C��1��W!���:�Y���-n� ��Ď.�!�Io� ccJ
I}r�f	ԥ�!�DZ�**Eq�G�l��M��W�Q�!�d�>z@�s�.�H�x QŚ�/�!��d_>$[p���	�T�ؗ�L��!��g�r����^? ���HӋ<�!�DQ���Au풜 <lɵfU�aA!�n�f5�È�*�.�UE	_(!��E!
�5;S�T#d���c$-�k3!��Y�By���eP�%��Tc�쟚^�!�D4��{B�R(b���w�ӔS�!�� ���J�-Js
xjGȈ=d�~�0�*O8�@�D�4���3 фH�J5)
�'?�eɲ�M�?���qCF��J�h
�'������73Ƙ{��CXYh,�	�'G,U�cL��+,�K�[Cֲ|;��Ą�K��Í��ݥ��uS����N�@�ȓW�!��	7���k���<J:�YŃ��!�$܂s����0�R��@�2d�!�d�#d�P��M;���=�RƋ�����IcH<i�3j�n��9U�T�����=���FQ��*���N[��>����Sµ?u�7��r ��!��]�^X�-D�'jï!�<��� �IY(a�rlK�p�>�2�k��\� ĳ���)��)J�>����K[*����%��!]8$����2@ʼz���f�'�r�3�-
�G:Hʑ��,V��������<%( �Ŧ#|�B�+<8I�i����'Y�vGx���1z�s'�S)$�0�Gπ�HOl�D��8��T��'�Oh�a�voμj*�	3���[��!Y�&F�n����f�߳&��ı����KY�b>)˲jJ#kَ��fʷs۪]���y�RYQĭ���X���j�1cUNeQ4m{݁ZC��:jٺQ��ٖTQ�tyq�=D��݋�D�7RÂ4Z7�Wybo���r
��G�D��d�pNH�J�9qD$���_G��$0�aE����c�D@�>��UT*�rF\�*ڻ�M��Y��T�AP�BҜ]��j�0��H�a��4�<�i���0=���E�ꜰ��C�^�%�H7I�r�3aK��,������pE�X��
w�n����P5��K�Hj�R��W��t�(��wĦ�B�pH<����O�S��c��:a�]qrO9�?y��ҫZ�vmPP�����o	�Z���'�ܟ
��ʚJ��$�UOO�wn������]k	�'���ї��:�y��U���-�r�ZǏN� �y	�i��� ĥ�[�����=.�l�7OBZ���b
�o�-G��ɩ��C�1`���̎�9�@\��`H�m�0�抾_�����ŧm�@��H�O�'�,�k��܋W���#���<��hʱ���©P%�\�\��ȳL��(�S@Q����eK>��t�!���{� �~�I��]"50��4�6%
ӓ���z'�X����[Y�ip���2������� �B�51�V@5
�A�56� P���]�˧q�xXIw$J+�J�[�aQ�a�X�ȓr����ԗ��ɳEŉ�\a�-"G�A�}hXUa�m�ZT���%�"����;z�����yW��)@A�l#/� <�	JT��	�p?�R�Ѩ��㶉M�)A���қl�\Z J�:n�܄�RdD�<�� ��& ���˖�x�'i�A�@]���O�<"��As����w�@Qʾ@�"�̟�be� 17!�x���0PɑCB)�e��JTh��OZ�4�y%�KPl�W`A�+��`�G�?D�9���~2F�:Ԝ�y"�M�(�n<0� ��v��3I!pڐ�*�����&ѦQJ<��3D_�K�Д���'"/�a�)�R?�U	P0�6QYw&��U-Q<O4rEY7� �:�x��_����pb�����0�n׵E�8��E�]�S�I��v�(C�MehX�deٱ9������l� m`�ǏH��$3��4��g��V����J�av6š�40�5��#H>{�䅁���T�R��s��?Y4��o<1�P�PJ��Qt���WK�~��=)5͟�m-T�)���}�Y7��S��y�vB�R�pA��,�r$��eM��M�J�/I�!�r��X���㠄��g��8�uf�2��	@�\C�I�N3ܰ<�C� ��8������`��n�;Xv����R)?�e�h�6n����@g��Y2�� 4�ɔj���#���?9�� ��Ւ�˝U>P��Oږq�vY3�#ғFda�reO�-P�$��N��%$A�%,X��� SFB�� �I�sI�ʱ��^�p!xŤ�?Ś(8��J�<镋UJV� l	qL���'�����/<?	�K�H�Ńߴ ��|�EgF��x�$\ {�l�{2�
��u�� 9Z6tJ7��<\���#��^:l�@$�<ġ�ػ2h���@q���c  �(Ղ�3��>�T�B�K�kƉzQ����aJ�P��[%�T�q�v��ץI	��I�JݲQ�H���#�ey�4U��"U�X+A��1�ц�L���i٩N1�L@��"n���u,�ا��5|��K�| ��i1k�X{� P�,��-��Gb��L��4��9�	�b�::(hӧ��R�:�8Y���$W��Da��t�'Ѫ��S#�+O��DT�*I��V�v�5p�+�(��� 0'yt�ӬZ�G�H��H\v(5�� 8���8�Tbb�xb���d�.8�U��;Ҷ�Wř�y2��X7��'t���o�p�Sǚ���0+����|�8�w޺�kw�͙qԍ����'�d<��~Ӕ<@�/͉�8��F�7n>�?��A� ��!i�Bߚ+u�����[�4�#�AФ����2(F�y�,Z$����G3/\��2��y��ӢH�8��ʚ6��b���y��߳�d�¿{=��Aƞ��y@�_�P�p`
LJ�+��y2 ؽ8����O�TaS�f��y�&϶�,�+���io���B���yb��,1��d�Y�8�dF'�y�W8M��Dh��>SP8�SD�M�y�[g�|c�C�H�؍`�Oќ�y
� ,�*��L*7}>HhC�@� �""OV��S��r8Z-�U����j�"O,X�������F>W�&�#R"O���Ai��]���S��� 7f�u��"O�͉��fƮ�
aA�M0n��'"O���A�4�ݙ%��5�H��"OH�ҵ�G���qȣˈ�N���Z�"O�I9�c$IA�����Pbv��0"O��3�D��e)浸�i$5a��BP"O����GVt�ad�>QH�*C"Oxa��,$k��SEB�#5N�`q$"O�`BQj_�lY<m����'"m{2"O�#��+z#�1�R���By~y!�"OD(�lç]v}��mʀK��#U"O���W�C�v@q�-0,���"Oh5V+��>T������0T�~��"ODiG)E�t��a�b�X`fL�2"Oqʗ D�@#�Ṕ��M
�ezQ"O�ei��Ú���*&ĝ&*R�%�3"O�Ӄ�2rv�\;�D<[@r�&"O�I�P'Ґk#(	2���=3��B"Ol��RK 6
:5	�h5R.���"O�0!	�1��}J&Be�x�p�"O6](��,:N阳��/fиq��"O���dA�l8~	��@C(5�ఢ"Ob�K���8��� nצ?�h��"OX�:u �`s���V�q��id"O��K$�[6��D#Ʈ�4���qe"O�d;��\Ryf�6��5:��iG"Op��E�ݿ.4*�Ӣ���])~%K%"Oۣ�ц �D�eׯGzL�Y"O��7 ��q��`���]�w��iy "O.!�s+�Yi�LUÇ�#R�i"O�4����QY��`��|�����"O>���m\:QR ��v����"O�(&�E�F�A�`�3.����"OΨQn b"\�	�b� l:���"O�p:t�W 8�Hx%�R�UE�T��"OT�����$_1����&��10E��"O�{A��Ю��e��>pP��"O�y `$�?�́r5���C4"O��c#K34 ���DǢe����3"O���4�<��`�a$��3��"O�=��
͓V�.�q�@ސ�&"Ob�!���	��nCO⺭4"OZA�ç0XSNtR5-�
 �l���"O���C ��6p��*ƌE;�"O��x�E��%f��+�[͊5P2"OD��b�;w \��HɭV���"O,X"G�K"'d>��ƕC~��"O��� �<;Z��c�#�{nPA3�"O�U�Ĕ12���a��|�f�Aa"Oh<��֥q" k�><��"OT��AF�s56�Q'�I2��=.�!�L���l�=Ip�S�ȞbJ!�dɈ!М,CD��P߾��ǜ�!�ګb:r�s���^h���S�!�ė0��xe��15��}���RY!�d��T�c���a1�I��n�*pI!�d߭4&,�ÁX�H�|�_�>m!��n?�0�P�V���¦,�&U�!���p�h��V�\�[�� �ҍ�"&F!��n�:%�r��q��a���J"!�ć�2�Х�P@Ws$<�s��ް[.!�� �y�f[�>²�¡��uv�0�A"O�P�0)ґ*p$D�G@C��$A�"O����Eؽx��鄏L���	�"OL�E(�Ak���!�u^��`"O �v��9e��0p`
K�M��"Od�W�W#i�����	
���0�"O~�[E� 't6tIwk�7�Z �#"ORԢC���x��+!
�pA��["O��25ѮBk���L3
���q`"O
�I!DX��ks��.0�d�p"O��Rȍ�X�V�@��؊.����"O�I����r�@haUG�x�,}�b"OxA��K��iJ#&���F\@D"O�胄�h��u�㦇�6��=��"O�\�`x�ˇ1rZZ�K����!�dS�S=�"ǅV	gD,������!�$�W	zM�4o��$ืg��a�!��U/m+���Z�\˷�
_;!�D��`a�"�<��dc�(�!��~��s4��6j= �"�W!�䞩*����l��1E<d� .�%,�!��>7")2p�A8`�2T#!]�J�!�D���y�.� �H�%�N�!��ݕ,���"f�4�a�Ƈ�)�!�D�*a�xؙW@
nd�We�>�!�dG|ݪ�H�!B^N,�"ŭJ]!��!�\�)���Q6�C�bV�X6!�$�. �h���םtlqua�,�Py�있7��р �P�	��a���y�㐝C*��0 �� F��S�	���y��u!^�(�'����)��]��yJQtɞ�Y2K(r�X|�v�L��y��W�T��m(l�d�@�A�y�\-q���qqo�+n���U���yr��>�\�:���W�$�R�\��yrɋ�;��x�A�Ę'",jV�@>�yb�822��� �p���d��y2�nz-H򯐅<�v���k��y2+2v2���K��|�xM8E���y�i�>�D�" 2�HŸ��_��y�%�yhV� "�z�"��&�K#�ygJ��*���D��ɡ��@6�y���0��ҤL��;6�p0����y�ŏ�e#|�ń��:�6-�2l�"�yB�.8�zݻ�,̂5��1+�	��y�*M�K/8��5��>����A��y�eQ"��Z���1�� ���y2b�2z�r��p�Ĕf�&�x�+̟�y"����q��#�A�\�2�H�y�/�y+�D�g��;e|`���y��N*2 �=z#�Ŋ*y.Ȼ�h��y2\��Ԡ�DD,-sz��fi��y�싵c��=:��U�L�����\&�y���0�"j̥���E��y"b��C� � �\\9�����yR�Kݤ��P�)Kj�� ͗��y��Ȭ�naP%�}�B0����7�y2E^�����KZ�r��; ��ybo��#�fM؅��"tk��!��\.�y�!̺'���Џ,s�@�J�mݟ�yR��$C����ߺqXah�K��y�+�@���G�^m�8�F��y�JA0%6,�E��g��<�f!�yb���QrI�d��S�5��o���y
� d`(�FQv�I0 	���@�{�"Oz�	U���"�Y��	2J����"O��#���L���{��N�p�l��"O�M��G��W�İ�r$�!����"Of�"s��+@j�����M�x�u"O���&J2k���jrEΦB����"O�aF���]Q&�qP�ҙb�L�K"Ot$SjE�\T-P��i�\j�"O,�wK8e��Q��A?r�^��$"O�pRs�c��&�ߗb��m�"O���6�Սg���v !!XhhW"O���r�A� )"�/P,N�lB%"OlXk������¨Ҕ{5�-!0�'*�1�+�yX�H���@�<���%Q�p���s�tt��[�8�hy��O�4M:��/@���6���c�	��01
�Ҵ9�!�d�J� �Ҋ\�T��)(6�Ɵ&��] �O3-��qbe�ۃb�f�Q��K���\�88&ٟw!�X**�&K�8Ț�j�F���>��(�$� <k4�C��p S"�Za�P��<{��aT/�2!��uƉ5�M�'�S�?%�f$I���zC������kp�Y9F�EFzR�R%V�F���I<���!w�2U�-<�<Dˢ�T>0(���1�ڿe�.�У)ö*FT�;�B<�O:�	t��'�QAE�ޑe�8��i���b�6/����	��&E�Ө��F'��J�i��sF셰M��*�ANxoZ=b�%͏�~�r6��B�I�NV�d����?�8XB�5�^��Lh��Ɂ�l�&p2.�1h�MS�t�v�Y�;͛&�$��;b4CB۔9a�I9�Ͼw|ju�����䊄�G�`O��C�D�)j�:m�  '<$ĽT$�=1A��V��'�������)ɽP�E��DOx�I<D/��)Ō��]��s�B�"p�#=�����ȴR��O��C!�:[��1j�X�zJ�i�Y҈.q��Q�@���C;��Ta�/aPQ�2���0<1&c�9<����HE;d�,�s�æ�CsGǙu{�x��'/��P�?6w|��ӊw��M(��i���g��Zu�ثШ����f��>z����uO�t�5�X0&����D�!*�,e�dG7]7�K"H�lE>���6It�|�E�Y�!����џ<���=���
(+������;%t���*�O���v�IUT����*H�e��D[�5�lۇ�OP�hr�& �\��L��ꡤ�KL���J���d��>����@Ϛ�x�T"O���/D�U1���B�^�b�0`��>��E��a�0(Q�9OxH �]�f�Q���y� ��'I���Q��5R)
���� 1�MM,�`��c�b<yP�ܓ��9��Gަ��aI��B�'�%Y1��N|�e�|��NF�D��B�A�B�j,yf �v��8#0[t3��U�S�̰�P���"��������4�Ԅ}����5�>1u����Z�%?	����8r��u���
D ���6��=�P�Ñ ��P0Ba��"��Į;9e��Rg��6}����k��^��e��,t4a��.����E��F���0��0[�Y�+>T\�x
׬l�$2���2mp����O㐍��� c�����*~�����41m |H�K��})С��&�%V�t��}�
�4�L��K(9�8���d��q�ty�g_��D�³
�hGB�S�@dx�U����I�5-�~����s��:x�d���C�~MsjX����d�-x"��sg�i��!˃��9ƒY�T��	&�������2;R(L�s�i�
}���Ha{6��*y�1���Hx"�яA
ұC�#��-���"ғ&*qhF����D�@��⡂P��t�A&oZL��	�j�Urq�ɧk�P���~l�Z�j�^����G�, '�	G�I�O1#&��(C� ��ѓ��@��B�,Dq`���,����~�!AFQ#R��3$�lI�(x�GS�&�����>$��HtH�,~<����*9Ѵ`Go^�F�D�`���h��#-�p���p$e��A���������9>=�0h�Ÿ�����
��'Ma}"!U=BH����g�Vb�+O�|,�C)��UM$A�FD�G/r��TL�8�>JŴi׀0X�'W���DxRF1l�~�kfǔ=;/�<�� I"�hO2�q��]��I�fu0a���ں`��+J�y�m\-�����/�`R|��'32�R#�T�uo�I)f%�?)��p�'sL�J��Ty�M������)Ǥ𫦧�?��D(B�Kl�*�o@&\�   �f�.�y�e\���� FVIh�z���'.��"̋x�O�Lq��P���YT��/�Ҡ8�'7~���mDXU3��I�@M��'�rS�A@�j,*� @�RM��[�'���I��ڜK@ޥ�˃U��s�'0�<�FNeZ pu��V�JH�'Ġ�B���
�����TWF2����� (��S�l�|�B�	�%�@�B�"O�����{�Pc�&\�Vu� �B"O�� l�z���e�P
\+%"O�	�e!�aI|q���#���`�"Ox!
Ƈ�+'G��3�ܣ"�ȑ�T"Onu��J�|`�2$)��%� �!�@��ɒ,�R�`SE[^�!�d�=1�`J�3_ٰ��4怮N�!�d� y� �P� �7�셨�ŀ~�!�ҳ"��L#��W�iʖ��l�`d!�$	 
��;D�/.�͂v��,d!��O9����i�;�e#�B�C~!���E<�i%Ğ�Q=R��,�!�5{2xa�ւЋH$��3�QH!�d2!���G�س
��V,.K!�9C�X2�)�\�Ǫ�?o$!�DW�k�$]���=, E蝷y{!򄎖,n䕂�����2�ǓD�!��-A}\��A��U�¡ ւ�!���^�	�f�#���{a��2q!�DV	]۰�0 ������X!��UL
�����!�4Pf��=_4!�d��UKB�:�^+����&-��y+!�Q2Ťc���.����6N��7!�D��!��S�g͇r6MC`m�&s	!� đ��&�����
�C�!��<=8�T�e]Y����k_7,�!�D	$Q�z�cI٤�y0����!򄍃WOXu2�IU�.�V��f)	!)�!�ۃ4S��*�%ܖ���RG\�	�!�$ղM;��+�o�-�aڧ��v�!�ި6+�A�BŘq ��A%���!�Q�e�|59�o-��1#� ��!�$�;J~�h�Ư�:IK�N��1�!�®T��z�	|T�SӮ׹`!򤊝/���nƿ
jZ�9B-��!�9����&I0����m2"�!򤙑a���2��+�~�ö͈�}�!��R</x��kV��Z
ի�F�b�!�/XH��zf�LIm�h���0K�!�䋑h�j�B��LbQP��ܗ+�!�D�-���ʗ�P0b�b��O/'�!�@V��A�cX*!XuKa.�K�!��'�.1���
8Nɒ0'ù>�!�$
�KӸ�q���%�Xy�T(׳	�!��M�wc��E�"c�Fu:�ʁ4�!�d�95evt�2(]�p�����^`!�D��`IH�(ڈ�h�"��e�!���=|��+�l[������g[0(O!�dAR�E���W�ན�c�?�!���%����a��.�ZX�e�Ώ+,!�d\�1nRP*���r>��B��f!�č�Җ1k4�_�✻CH�R�!�ğ�l�0[�6�l���[�G�!�ĕ</Ԃ��V��!d�ܥ[FŨ�!�dQ C� �	����j��1�*	f!�䂯&Мٓ`�� �X@�SF�!��~�ر!޶'pLLb Ȏ1�!��<BA� �&yC�Pi�H�!�$�Q-�pd�fN�8ɤH_�<!�M�5��&`��;�8�h1<�!���}t�g�(
�C$'	�q�!�dKE�6�(@䔶5����޴`!�B�<���S�B��A ��KWd<1!!�� �(�V&М��P��Ϟ$6B��"O�$�3Ɩ��$<�TCۭn����""O\���] ���Jl��1�5�"O�z��כld�A�w�D�v��`�"OZ��r�^)Z�Dͨ��I@Ľ)0"O޴ &,˒q8-��J	�h���;"O��cef
�P��v��8l�:L)�"Ozdk�9uh��P�s
a`0"O�K4n{�����N]Lu�!"O�x
���$�>PÂ�#d�@!V"O�ȑ�*]�d�xԂ^� |؝�"O�� W���E5|̀�� b����"O���!ӂ9B��ӯ
���"O�#����f(��NA�2���p�"O�p�
�(:de�RZ,%��,k�"O&�A�l
�\���U�d��=��"O�h[�e�a+P� �Ump��"OvA*F���H:�X���)@vP�U"O=�v�8�FY!t.��/O�l�B"O��s叔<@B8mݒE%�uJ�"O��qH�S9�	��I�Xx�V"OHP+�Dȵ7�҄Z���*z+��Y!"O�Հ���h�l��j��N�0R"O���P��V~0J�I�J�J�qB"O��tdQ�>0��B&W1�|i�"Ot�0���5?�����<�0�`"O�,3�-��|Ք��!e����P��"O�Q���N�*��eXV�I�&"OPP9�/P6xً1�ɉ)q�$��"OLISo�'O�I"A�>hf�1��"OV��V�ߤ*ؒ�8��͙S�b��%"O����Eg䠰��19��0X�"O��C����xj/�7����"OzmчB��k�lA����FX�4"O�� Ō�x�Zx;�-�UO��+ "OZ0$[��AJ kU=�\��F��Z�kԿOz�Cjƒ��=`�4O�~����Vv�ք
æS�m��i�'�ҩ�'�^O>�*�����tp���?N�,@a��z���@��W����L<E��f�v���b@|��V�7\o�%`�HH+!���jv���0$��L��� mX�� ��W
�K�Nl����-%��b�b�t�L<�O;vu��T�d�B@p�-n����y�D�n�ēç` �L ���Y��视0R
.��'9�8��oM�������XЂ��*��Fx�rٞ�yR`���*OC�S�O�� [�_#s�L ���! r�!f�H2!�1:�y
�'X|����(qyl���$=DPې�Wk̓=ER�ᓭ%��� (�aH�Y�T���c�\�D"����݂@��0c?7-B�?|:P8��a�<�Cj�	��C#����=���ԧ���d1ŧH<;+$}�!ʲi$  C "O��X�΃�zHX5�F��bPʨ�y�HDd ��DF�&6�e��'�?�yB�:o�l�Q���1uD9NA��yrϜ�x缨�1���j�0p��R��y�FF:>��s�a���1�C�HO�����i��x;EhE�|��,
�նm!�X Z�>�!��Q2@r�pE���!�$�)cN��*&
�Z�g&T\!�ŠA����ыF�@�hTYԤ��-@!�$N�8�|��nC%���CVH�w	!�?�F�c� W��6�:C�>=W!��ɋut�9#G_�^��݉b	3{�!���[�I�5V�M�t�����=�!�N>��0Ӧ#�Rᰳi��W�!�d���엃b�މ*��~|�)#�"O��re��<�C�lQ�>����G"O� �p�ኋ[f
����֝��\��"O�=X�_0i|��� Mi���3"O ��q��-��:dV�Gfh��"O`0��F Fc�TqW#G!aK�٥"O��j�b�-?��Z l !?�qP"O`i�2�����L�4˛�T8$���"O���;84q`U���|�F"O���I,s���CaR��@`@"O,`�1'�1d���	��K(�͂�"OB��[{�J�#��a�,I1"O<��)ׁml^�)SC�\��X�'"O���N�'K]����% o�`�"O:��Ad��}�ܥ`�$�g���"O��2c�%)���@��t�Ԉ�"Oh�R��[z���"#�)�"��"O�2H�>�M �B�E���pE"O:ࠠ�-�����"�:��%Yg"O��@��I>��d�%��T�"O��U�Ҋ8�lP�Ҿ-gH,��"O �!2���:� dȝF�����"O�D۔��?Hh����/x�ʁʗ"OJ�q���	l�U@B�>w'�;�"O0h�Sę,��=K�@�u��a�"O��*�hQ9[��E��Z%��"O�0(,WFR(��P�b�!�#"O^�o2 � HY�&�d=��"O��9҂K�5�3&%����"O��&�U��b�#�&����RQ"O�����&`��k�Պ3`��p�"OHa�`!Ιa��<AQJ)$Ji�`"OT�`���4����@5W�%j�"O��hBG�R�YX2����E;�"O�I�w@�HS4T�� K(8�"O<��3#رG
N�2���R4dx�"OVxU���X�
`�?z��s�"O �;ve�- �p(�"�6|T��"Ol�kw�F�6�p)!'��Q�%2"OJ��K�8^���c�6,Ģ�+"O�%���ÇE.� wO�"%�T�"O �
B+Ҭ_�x��M�:czX�4"O��a��Tqbi��,��V$��'κ�0!�"+R|c��,i����'�Pl�vwa��ڲf��$t~�S�'$`E��F�"�2g+5�6t��'e�4:�Gd�Z��4G���kMD�<��n�" ˠ"+X��m���i�<���=yQL$�oҋ7����n�<afCO7yV�j�.��q��I����B�<Q҇_0_��@�d�ƾ|��|���i�<�n��C��]��a;g� �0!�a�<�E�>6�3��7R��	*qR�<���{��5@�g ?_#!i���Y�<���<_l>|ʒ��>���ȧ�V�<	��C+|h�3���p��H�ƙI�<��U�
�UB!�t=С��HZl�<��+zhp��!J)%��x5��k�<��&N�h�J����=p����Řd�<���7uF*�@M��j�r쉐��t�<�1��WMf�Ƣ�7�9��Fr�<1G�H6q:$h@�?c1���o�<9q�'2��|Yq�â?�4��m�t�<Ѣ�V�8^��e�L߀�"W�Or�<9�I_V�Xݡ"���A�k�k�<����}�]��؅n�ډ��_�<� �4��
��:S��ic��%h�@��"OH�x�)��TZ�(P"��k����"ObQ)��,~�20IZ���"Op�c�P��z$IN�3�}��"Oj��VǛ0(|�8#g
�`��]�0"O����-��o�J�{%f�8�n9��"O�b#�,� �A���1�p��"O"5VH��"^�5�]�H=3�"O"E�tB��YE:�S#��$+���#"O2��2O�ocr��UE�2fڜ	�"O\pR�6�^ ��S0T���(b"O�4����N�`��Tƚ�Z��""Oj�ڣInq�!g�	$T�l�f"Oܴ�⦏�?��:d��>���"O =���� �D�[�ԫ�F�S"O�|��-�E"�5%-P�*��a�w"O�!�5C�i�@#Պ�-_��T��"OlIӥ�D�@5La�iX,��(�@"O"TS�N�8X>�u���-�r�h3"O� 	��K�0F��Ǉ�\SбC"O6�h�k�.	5�\�IQ<F���"O�(Ї.q�p$�����l=�x��"O�P `���9
��C�d3�`�"Ot(ՆJ
_{�c��]�#˚���"O�ՠ����V v��e�}���A"O�a���-��u�ԉ��F�j��&"O<��r'0D7��y��.{a���"O4T�Y�V�C��8"��2�H2�y�ʓ&G�<;󁇫m�Gg'�y"h�;U¨9ю�5h�\�(l�:�y��X�H����aK@����G�ybf�5bw�D�Կ0�\�����y"��q���s�+��54ԱJ��Y!�y��;{b(�
Ƙ4 <�э�%�yB@��c�I��*N@<���B6�yB���]�b�9A܈���pcѬ�y��@\����* 	�>�+U#
�y�И��@���U��3o'@B䉼xX`<���:"B�aD@��3�JB�%�,����G�	k ���&B��5e���F�K^��da��ܿN��B�I�r��1�C�^�&�+枺y��B�I�\MV�"'�6?ԑ���X�	��C�I Js�����?v�������}�C�9T������DL��)���?"QTC��a7�]�үO�`\���w��J�C�I#"��dا��Vi�C2j�$�C�I"X�h(pr�	&.�:h[��R�H��C䉆k��I4f��@��\@�iϐm��C�I�9��b�)P��9S�NH�C�|�"- �#{��F�د j�B�I��� #�(�/xB<2�d���B�	�V�Q�D�3*v6<�@�$�B�	��Ɉ�AƒS�>�;��kϖB�	�L=y�\�n=������[YlB�I\6��À  �Q}�JB䉘)�����}����,Y���B�I�%�0�C`�,[8�l�u���E�C�i�A%\}V�;�i��:�T���9D��wk#-ж<�禊:M�>Yp�,D��Ѡ���Kn���J�01���+D��qB�-�8�C�Ɔ ��3D�d2Æ}���( �!��'D���Ҁ_/4��x �j�L'�$D�� L���Ã�]�*��cnCa�&���"O�Y�'aX����5-�#Q�UQ�"O��)�C@��N$�P�\:�@I�"Oй`�MY	�<���^'B���"O� cn͜/�ڙSi�,
)�"O��X��b^
[�Q�I����v"OLq��Ϝy��8uϊ��.�B"O�4Q�ʠ<\�afa��F���"O�[@�� O��(�/�U��st"Od��o����5���7�t�`"O�P@��$e� ��N_���]��"O���mҲ�*ȢB-M�>�
���"Ol�b܉;�&�	eӗ`�p�Q"O�i&��)\�|�7��16Yp��1"O���I�����iJ75&&��"O0�QCƛ=����G	6l�v*A"O^����t7>5JQ2�bM�#"O:���L��ň�1�p	�"O^x{�`�+?e�h�D_�"����"O ��e�^@)�xf㏟i	taA "OH�8�	F��!��3X�t9�"Oz���3�Q��`��y��@��"O�T��r�L���^=�D��"O��/ۅ-Z�������D"O|�tޟ:<� ��?e��m�W"O�q�"T&TY��V k�^���"O�ِ��u}����W&�x�"OΑ3�/�FKrW��2z�8P�H[�<���96f�� g�+�1Q�X�ȓQUT@���ڦ7��E��D��T��4��4���B�L�%Ǻ����µA�l����(X�T�X�B�D@޳/"�%�ȓ� <��.�&1�w`

{��p��\Dt�HWg� I��씄<K�E�ȓ?Y��3tg�5�$�ƍ>����j�\0@�H�c~�;'g���ؼ�ȓ���ǬT�n�����Lȹn�V]��Y8�ś�,ǸdlE�T
ڊdU�ȓ2����bA�N�F�R���|�hp��C�t��� 0��R�Ǿ@tY��H�Zc����] ���e/hH�ȓD������&Eߘ*��8uI:��ȓh݌��#,�|�	�+K�=.h�ȓa4R]�'�&Cv�hk%�N�[��h�ȓW[�a��"˕-B>����V7I�Pi��aݚ��U/O�v�j�Ө�:Ѱp�ȓdT��s���'TC$�x `�j���ȓ[�4�`��;7v���>.莕�ȓv�QA��B��m��kܶ&��s� q�u��6DUP�-�P������,A�FC�((UkQ�Y�.�ȓ=i0���L�D�����+�����?�<�cV�����ƊF�@1�ȓA��s��86�1S0cݻq��U�ȓbN�s�$�"D?��2DG�Q̖���~�v$y�g�c�Ek��	pϘ�������a,�8D�+�֬@ɠ���&G�0Q�U�X��
�V(v@����e�n��$�*G35r %U��ȓzQ�hr���@��R��š~e���6�B8�W��?S��Y3+�g�V���Y<85��<#�v��ؗ}0bu��?N���
�Cp�;�\�j}�`��2��xµ��*�S�b�z�h<��S�? ʍAp�H 4�vP�4���"O��1� 
  ��   r  P  �  ]   7,  �7  �C  "M  �V  �`  �j  `t  �}  Ɇ  f�  w�  ��  :�  Դ  .�  r�  ��  ��  ;�  �  ��  �  H�  ��  ��    R � � J �  i* 3 w9 C xJ �Q X R^ 	d  Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�� |d��"O
`�(�;���8���-0��1%"Oj4��ND^[��"3/9�0|H�"OB���H��*�ʞRy=a"O�味V�!X��!&F�:J�$���"O,��a
���C�Ą�M�"O,$3%o�-���p���+Ն�:1"O��ݢ1����`���y14]2��i�<�6��{_���c�H�`�fX�$Kn�<��A̼VI�xR[�)�Ć�pඤ�ȓA5��('nߡ4�� �)˩%� ���,��r�؊b#`T�eT09���ȓ!�b��g��}�8�F��-? �ȓ
K|m�ș�VṔ���2�%�ȓ"R�X�j�4JN�1�˘X�i����̹	_�jZ��1!g��zܶ��ȓgil,*�J�
j�Ne��i�J%b���f	�(U��:���G��$Y^م�~r�� S�%T"���k\�jx�ȓ|4�1�îJb��@ӵ�ݩn�V��/[`�"�v4�R�!ʎ<��M�ȓ`:��z�ؚh�J�Z��$HY:	��H��p�m�C1��!��B:��0��EnjZA V;9����J[
2���	��4'J�EA�IVW&��~�(aZ��ӹ�>� o�Y�|�ȓ�f�A�
Ο7�H��M�$�����mޠP����/���ANXo*�ȓTv������h ��-7�*h�'��}��zE�	H�N�g
�z���?��') e!�NѬ���C+D�/���	�'�������]���*QR|����u�OH�!:p��O���A1��>y�Ȁ����*��9`Ǥ���t}�ѠܔN48x�Q��t����S�'~&�P7�����KV��r�B��  ��J����*�S��6f��Oz7�2\O����GA\W�f)+�V!�5"O�X)e-��R�"��6Z����"O��hC�Z�Ph(di"f�d�"O�9���Z�w����AG�e������'�ў"~��/0m/�8������``�)�8��ȓ���h#�!� 5��F��j=�'�����0=i�ۮ�"��%	)Hl��ƪ�`?I���k�3�<x����w.P	�GDA&�����%��l�6��[l���  Rhx�ȓ3*^y�.�:gN	�2IA ��E�ȓxBɓg�_F�5�D3�x��ȓw������S�ܵ�S#e׾!�Ip����YȠ�9u��4zׅ��|F���0D�HȂ�^�Q�U:SC7\�:q�D,�=J�D�O��S�$���O����2#鰴H#+ ���p�'e��n?���%��sPz\X��#*��1�'��~����
��ɨ4bΝ2F̤BɅ�hO��O��f�I/v��0���@A�V�ߟ�y��؍<�x��i(^�5��l���y�lE'S*Y;� A2+��Ģ�!��yb��A��y��A$Yjɉ�Է��{Ө�?E�T!H�R��D��lC
��!��yBO�'Nl�
�B�9o���*2�۸'��CS���KϠA82Ɔ�N����G劍Z�F}r�#����	�]�H$rcF��6w�\�с�; � ��=��1,OX�c�`�H-
uP!(O3P��J��Sܓ��π �����}FE��b��R"O��8v��E��[T�l�˷Q���ŀب�y��Ć��g}ʟ�Ű�.�� ��x�udI)'A$a�Q"O������g�
��#
N'6��(1"O�ey7��7{ ;`��1���"Oq�F�
I%|��rHR5MPaA4"OP���O	�,0vy���, b�$�~��9�g?�dh���p�9t� �O�h����r�<��JM*�<�S׉y�L��CAs��	t8��X5���J����iG�(qh��6}R�?�O��:W
�-S���!�޾a(�C&�	XܓaN�I�9��`zE�E�7�4Q��V8R�!�dƐY�zx{�J�J0츊q
�~s�\R�ӛW��l;�.Ng�v �sG�B䉇	:Ep�
�P߆H���]��B�	�y�4 sw� &�rD�T$��`��B�I><]��ȯcـ���@eAzB䉼m�Ũ�I]��d�:�B[? ��C�I�`�Y{aI�E�P�SL�=N��B�I5Z��P�D+z�����.��={|B�I�b���ԀC�k2,i�GTL�j��9�	�CH�c�A��U�B���8�.B䉖(h��sv�O%4�v�C΅�"���D%ғK�P,�D!�
�A�G.U�y�P0�ȓ1���*�)��*� Y�o�8�ȓK((���"وh��0�?@(�(G}���-
>��N��S��@���]���#<�7�|*q�Y;]ib�t�ӎm���{�nW�<�㎀F�B�5-��Z�o���}E{���i�t���B�#J�����T���1�'����S"c��� ��$�p鲧Ɂo���L��I�h%f`��D�E����b�<@6����O��I^�'��6]���BeD���-҃e+rN0���&杩Q��+W�z�AF�&|M�YF" 
D�O�~L1GIO�>w,�R"΁7oD88I>i����@\�9q`���V�L�ڳF��^!�$F�?Al�Z� ��1�����
W����˓)ܼ��C�&Yz��~�ц���l��1�N�c��bR�ȓX���32�?]^lu����TC�`�ȓh���z!��	8(��#U�rD�ȓ>rl!��/ގ(�a��
{u��'��D{��d"�v��j�nF!kxxQ
B��y�!^Xߨ(�����\�.���B;���y��$7�,34A*��J�pb�Q���0'pцȓI�2YI��	+�L���fS�,Frm�ȓyt(኷H�$L�f|zP��M��p�ȓv�~\��D
��F#�)�=Y�����AZ|��t%�9�rPVB��y��(~J<��M	*:��%'ԡ�y��A�Q�P���� U��4o^��y2Ú�_������M�a��,���y���of2a��k�=BN����`[,�yB@�Q����H\���Kܘ�y�H(J+0x�6U��@��݁���T{����$��ߠ�`�5a��w��0t"O(����>;ʽ�p��^f����"O��aB�LqDD[�'�7.�Y(��T�'j��OP!�J]=�n��A&�hT"OZ�*�oZ�B\���gO����Q��a>����ē)�`��n@-Bg�x�)7LO2��/����r���p(�ЕEo�TQP�)�H��(d�S���sX����S̓e��b>e��% ��Dɀw�5��9}��>A�S�? 
�ò���V�r%3��1���IҔxr�:�O�{TŭZ@�w�C69�(��2O\��D��L���s���s �'2�Tѥ1D��1R�ٱR�$���M�O������0��?%(�[�>���� P�v?�D
�)j��G{����+~�* �(_����H�Di�	Z��(� ĀRe4(@b�bw�ۙDNE��"Of�a <,��`��τH*���R��Ip��Oڍ��W�#^浩���0",�H��"OҨs�Hъb����w~� ���>!w�'&N�� E�']�&9�HD9HԸc��~��ģ�l���	���1#�A�5��'�az��)Т, Cj����!��(��Px��B�9�`���ƍY����%4�ȓBT��@�k)��Ju!]�Ґ$����I�P��Ф❢Bfՙ��"B8�B�I�;��xQ2���+��q�g��;�'��)#1���.xD�{V`
I=�|3�'�^ hN�2V�xa�՗	����
�'&�1��%m�Bm�����
�'?j\��E/.{h��g��3
�'�괋a��U��4F�F� "<��	ߓ`�OD��Po�X�*����"O.h��"J�;���!¤ɽE�\M���D}���>�|b�BMq�.�E�3T�\ C�Bx�ܬ<��'���a�DZ�7F�:��2��}H��$&<Oإ���4D�<��(^ۜ1P�|�)N�|����^C������o�pC�	-Z��s��
 b���cŒtAX�|F{҇����D�5dJ|�X`��<�q7�A%"m!�d��%�y+�%�HP��[9ZA!���%��ܣab�	7����Ǒ�!�Dא@(�0)-]7Fh5m���!��DfE4��!�m\��f�B�!�$81Sh��Iʄ,�����`�!�$"[\�F�Ͼx����C�7�!�dQ G��� ��E+h�,عbb]��!��]�1#�>���Цǉ�z�5X�'g�<�7eL�"�r�g ~f����'g4r#/DL�"�!f	��p�.���'��!D(/i�E*�	��i���r�'��yPcfJ*�^,�� .�t	�'*re���|�*���-PN��'2�uT*[�f�|!�q�7����'9I�&2-*cq���Jb 9�'�
B�#\�cL]����`���'�8�`۟
�n��'Ԥ]�X��'`��B�x���
R*�0nZ�'�~��d����=ڦ	H�\s��'+�Eas��)���h���p <I�'�VU˥Eڃ	���&�2o�ddc�'����A[xX4�"P7���I�'��]��(����7�NF|�a��'�4���,��hJX�i��?9D��	�'Yb�(d���G˘5Bb��f�� �'��;�<X���R�� ]��C�'6\D*@���>�� �8M5���',�P�$��� \�g$B<D�d�+�'( Y�DcO.S!����f��<��A{�'��k���G�5��Y:3��-�	�'~~ !�哽0v�bG���<̲	�'��P�UHrn1s�+%����	�'$F�8wC^ �HU��i֠��'��I��+: �x�soS�Z����
��� �R��\Ĝ=0�'WTB&��v"O���B���k�����I�x<��#�"O�-"c���Q1P�z�#�(o4�[ "O}�T(ׯKR�!Z�c͠m�TY�"O��R�ܠU�8�����d��3'�'q��'���'}2�'}R�'��'�����kZ�I~v'_�`����U�'��'��'�b�'���'���'7�pHr@ޡ~6H#sEO�q۬e���'B�'K��'�B�':��'��w��d ���|j��ʁ�F�P�6͹�'<��'G"�'"��'"��'�"�'|\\����D��:h��ٱ�'2�'�B�'/��'�b�'v�'O�)�����`�1��P;��ڵ�'dB�'Q��''r�'"�'A��'".i����:iž��SA��.nT�;��'���'h��'oB�'B�'��'�,xP����b@q�WZs$e)�'���'�R�'|��'G��'�r�'N�%��	�'�����3;l�hۑ�'���'1�'c��'ZR�'.��'힙�C"��w|� 3�����s��'��'���'���'��'�r�'Lp�hqa��p�xZQ��!��@c�'XB�'��'_R�'���'^"�'ΨM`�G�J2	�Gb�@���'c��'?R�'mb�'$"�'J�'m�x(�M˷'Þ��e̃N/L��'���'m��'b�'}�*l����O�����Ƕ}آ����Fq�Q)�lyr�'s�)�3?4�i|"�����8(Oh)����l"���$��$�妵�?��<a�i�V5pՇ��4Jΐ�De���cWAu����"�z7�=?�ŉo\���-*�4C��N��Ia�/�e��f��'��V�<D�T��a�&���&+N�իg��;-07�ل�1Oh�?����[#/F.�>�����cG�x�w
M�U�f�x� �IQ}��D�_�b��0O �aT��;A�t5h�ϙ`�LA�>O+�`�#�N�a'ў�Sğ*����D�xl���A�pՙ��p�ؕ'Q�'G�7m-'�1O���2FՆ>+�RD��d@�Q:�I:�����D�Ʀ	iݴ�yr]���� �.c2�����2& ���"?���íCԂ��V�y̧ޖQ�^w����@}����놝<�f�#�o��5����D�O?�I�F���`b�1o�UaD�<x�\�	<�Mc0f�p~�y�����nY��	T+�;6pXA�p
E�<�I+�MsѶi��ߨ/�V����p�A���ۆ��I��Ô�8jHiw��z :4$����Ϙ'���5.�%�=�7�ҖUN���Ox�n�KI\1�	����IB�';i2�AE��(H)��c7�;_x�
�R�@�4ٛ�K/��˅t3�,!�k	�'��xuD�.�:ybQ �O&ʓ[T�_��9����䓅�8Ml�	(Jb,,�e��a|r�p�|����O$D�"����Y���3n��	g�O��l�{�@~����M#�i&7����nX��Ȃa����ӟp�u)&�׵:��ɮ?W��A�B\h �p$?���ܡt~�8�/M�r���%��`�$m�'F�i�xH�e���%i
����ի`V�p���!Q�8�R'��t�tk�C�:V�M;�)��'�xx
�͚�(C�؃� ߱���
��Z���أ�J4K*�����U�>��z�'L�QJ��_*M2؀F�H>dᎱ8�	>N���2Ġ�bX�T#Wm�YV���Z Y B8@ǤO0x��x%4Z�r��Fł�q;�y3hк ��������22���b�2i�^k��]�&�	�b���e���k״<��E� ßj���7�*ci���D���P�>���ӳ ���'�B�'P��&R�h�	�D��@?a0�ɨ��Ԯ��@j����C_�Bg<q�<i���?y�&� �zc�i���!fk�GLX��a�iJ�,5���ϟ8��ߟ'��X81����w"��n�0ɫ��G�c�����3����D�O���OH�7���IB�Y���GIё�4���j�����O:���O��O8���O��{ ���p�yP��%i\�J1f�%1f�O<���O���<�d
��dC�M�|��NL�I��
e���M����?�����?��*�(���'pF�(UO��p=<���$KB���O����O���<�B�H����OL�j���[�nU{����7�P��Ҧ���e�I���0P=�c���F�^�(���{Bd@T��y� c�L���O��I�Y�,�����O|���=:j�h�kz*z<�3����l`$���Iş0�RbП$��G�	���S$lEsԁʷ�Jl�syr�=	�'���';��S��ػm훅�C�S��e��0�r�o��p�	�q9��?�~Rf�"X�N�K南91�)�����I�,ٟ��� ���?�'B�'?}:bH�3�8�w��in�[Ef����V�8�)�'�?A%I�f�(�:�MS'G�����N�>'�F�'C��'�4���V������IS?QsŁ�O���z�L3_@�)7��Y�M�,�<���?��bX����W���J��!Ȍ�ⷷi5"��]��I�������('���u�*u�S�ϲ>@�
���	^�W���I>9��?�����d�qT���4iY:�ao�$;*���'�<����?������?���]�r�2�� �Ov�8����oS%�רB��?/O���O,�$�<Q�̟!	��)ڡdER�r�guPx��d̻'s�I˟d��ݟ8�',��'6�94�'��÷EZm|���k׆jE~4i�C+��O���<QCL�*��O_�� �|�l�u��r�B�AW:�s�i���'o�	ߟ����td��k�i�A	H
�1D\�#�/⛦�'~�X���3#��ħ�?���ۅJ ����R@?F�-�D'ͦ��'"�'�X)C��'���<�s����z�l5��6�n$Ѵ�f�|�\�P� B�iKn�'�?a�'T7�Ix	���'�,{�t��E��t�X6�O��X0_���K��?}��M�k�1"��V�?r���IǦ��7!���M���?A�����x�O(���6�/q�DB�� n�m���bӢ\�P��Or���O�$����g~�Q
���;�l�%r�:��2��7�O����O<�����}�i>}�	ӟDRS�J�:��E����mR:�K��M3��?��03@�R_?���X�	ٟ0�sL
/cl�`0�H�_j.E��]��M��&��u�כx�OB�'��I/c��
V�
C(<�.ۜ,��A�4�?�an[��?�*OB��O�$�<���ܔ_"��t�V9P����L$*q��xb�'kR�'���͟��Ɋ1g�� ĀL:Gg����wl\�@���'92�';�����h��u��eV;	[���k&j�UÔ��ئ��Iԟ(�?����?�W��q��n�s?<��̀*D���g�׻~��O��Ģ<���k���,�&�Ą'_0.	�4&B�(Ő�����.7�V�m�u��?���g4���u��D�	�Mj����QL�(��N�2��6M�Ov��?a�������O����kM�xgf�ڐ �%,��*Q��V�'JB�'<�� 3�����]g�h�ǘ5	�j@��gP/-%�	֟8�b�ɟ��	��H���?���u'���o�t[`O��=_��(�#��M���$��cV���!J���i4m:�f�!E^a���<d���iP��'��Op�O���ձ�ֽ������-5�ŀ%�i��';��'��	O��'�R�5<�0��4�hbRd�V��0�P6��OD���O"��u��J�i>A�I���ÐGW�X��5铋�.�Rp���:�Mc��?�-O�����D�O��L,F�8h���ũ U5 �Jʆ	5�@n�ǟ��G����|����?�*O:hKu�S-p��Q��6p�<,0u��˦)�'�R�|��'�BS�p�4M��4��	�#�\u^��wݱ��RK<��?!����d�O�������g��f� 6F�;;��7��O�ʓ�?i������O�D�G�?��r��B[(:Q�F!5���[�Bo���D�Oh��IMy"�7�M�Rˈ���a�c/A4�'�L^}��'���'f�	� 	�%�H|*"��$\/���!Ñ]��8�����<K���'��[���	~�t�'��`�ءʓ)C��a3��F�M�!m���I}y�,Z,fV�b�D�k�-D5*\��%\P�2�z�`�a^��X����������&?�i���P��;Z�$����C�%�TH磩>��H��	��?���?a�'���fy���	'$�Ts" N�W!T�3�i��T�@�V�!�S�x�̼:r�&p��t��!�7��nH�oZ̟��	��D�S����<�e�Ň$x�p�JƷ!�F���eDr֛�����<Q����'H@S�T�3�JD�t�W,k��D�&�w��$�O�������'��Iϟ��z2i9!C_���Tjr�l�Z�n�f�I�L���)���?a�LZ��� �\�0t�9�&�2�Ӕ�iR/ʯ Z�6��O��d�O(�D�[�4�ONt��㔜G��i#���J�@�q�Y��[��s�@�'/"�'��'".
D���	T�]˲�G�;�*m9��jӈ���O����OPT�O���l�1A�j.�t�UG�-*�J�Z�S*RiT��֟�����|�I�h�ON\��t��U����~p@]Q�]�!,�$p�G���I�8��ޟ��	Cy��'e�a��OV����y�ڍ#�H�8�m𑦳>1���?���?��TL��QE�i2�'��@Y���Wn8�2��'��x�ouӜ���O��Ĥ<y��~`Χ�?��'Q� �􉏵0}B�bנпsO��Jܴ�?9��?��9�D�A�i��'�b�O$I�"�ﺩ�.ܜ(\��*�,y�^��<��3芕�'���|n��|v9���͔ހ�pC�A�N7��O0�dB9"��n����	ğ�S�?-�	�]�d����//�6a�ek:(d\$y�Oz���j�����OP��|JO?}��Ǘ��H!��S
".z���n�fmJ2I֦���ɟ����?��S�@�	ڟ��ˊݰ�( ���Ua1�!�M�6oɏ�?QN>ͧ���?y��l��x��E�D���RSK���'��'KV���i���$�O�D�O����� vdH���S�.��Q����i�rR���Lj��'�?A��?v�#W�R��0��m9Z�
� �%?̛V�'k�Q* BgӀ�d�O^�D�Od��Ot�D	�d�Buo͵U'�A�n@G���8��I<�	���	{�Sv�<�����>
H�k c �iD�z�.��M����?I��?BW?�'�rMGY�ڥp��̂m�E@D��D����'��I��Θ�2��?a��"r��i��i	��Y�0Q��l��Hg�l�x���O<�$�O��d�<��E��8�'c�tE�R3C����b�(&�T����i"��'/B�'�2�'r�Vl-���'���(/��)m��!XP|I��B��7m�O��$�O|��?9!��|���~J��I���	�ǟ{6�irT��!�MS���?����?A+Z	A����'u�'���g����Qr��t�r�b�/ e/�7�Ol��?���|�I>����(IR��I3b�ƻ4]�e������O�E�d�R�����������?���ݟ�I
� X`S�韼 ��Y��ŉCԔQb_� �ɭ>*���П��I`���~�d;�
�h��_��
�)���H�E3�Mc��?I������?q��?��ڲ%�Vq�R6R��צ�=q�V#_,���'��+�~zN~
�*�L8 ��L'=K6A�O �WB~H�C�i""�' ���N�7m�O�$�O����O�]��l�`ً+��HaU.�k����'�I+���)r��?��]��L�g��B��IABiQŷi4���4e�:7��O����O��DWg�4�O�Ģ�n� S�qNI9=*Ш�U���a��'�R�''��'��7;Ԕ�ƌ�&�f�Ń��P�3,mӚ�D�O����O���O��	�4!hKo�T��d��fT廀k�?Q���	yy�'��'���'d,�a!t��x�Ѫ�
=~�7D�K�0��6m�Ol�d�O����O���?-�`���ّ���ܨ��mQ|����m�>���?!��?��K�i���i�b��%*3S�4�v�ބD� �����?9��?A������Ola��0������$�d�6G�0�;�Î�9�~y҆t���$�Ox��O@�����-�	͟��	�?���e�5�hK�\56���b�'[�M�����D�O�h��ɺ<�.O�i5l��1��iBB�i��^9c�9hߴ���A���m������O$��\~��Q�g�%�@I�Wfщ�b��Mc��?1�)��?�I>�~��PJa�ū#�|���Q=ꈙoZ���$�ߴ�?y��?)��x�'�B��A*P=abo�/���H���r��7m�5c�8������A�}�y!i��0��}Ȑ�K�M����?)���@	՝xr�'b�OJ ���}�$�/�.R߸�x�d[�bT1O��D�Ov�$X�.���1���84���Ϸx��l֟��gă<���?����#G��Y�"��#��?td�a&}}� ئ78�S����͟��	Oy��N�B��hFQ)ëW�.Yn��w-�c�NO����O֓O����O��.̽+�u
Q�T�3>"W��J��$�<���?����d�&KJ���'g���x¯�|	�3A�u�DP�'7��'��'6��'Ú@07�'�L�;E�A�b ñ�S',:\C���>���?�����d_]7�t&>�B�%��e��|�C�UG�0�����9�M������?������I?B���頊C�8��!�ջch6M�O>�$�<I�Ѣ;��OR�O���p���|c�E[��	 �>���'���OB�$$M�$,�T?]�0k��N��m+(X�<� - �@e�d����i0�i.T�'�?1��z��	�q�� �!��.\x1ᰦMJKJ6�O"��M�YP��D)���Y�3��㥎�)���fNn�֬^y�7��O���O�I�z�I����T�n vh��n܉v^�j",��Mۂ)S�'C�v���D����́-r�}{K�P���nҟ<�I���CRb���ē�?y��~�Γ:l_.aioūfE<���ʁ�MCO>�Q����O���'�۪r��l��r�V�B�?��7��O�x�n j�i>qDy]oQ������µ*ъ�M#��A� �������O&�D�O<˓x��zg��L*�y#HS'
��!��J���'�����1th�:�H�Y�+��=��`�K%[�b��	՟��Ɵ����T�'�Z(�ҧv> Em����P{$cG�k-`x�'�>����hO��4[S���� ^��IY�F�7A��eE�Hjj�n�����	����	����.uN��$�Ob�䟔 �x�'��)��p־lZ��<$�x�	���j��Į��O��R�&LS���G	Td�hԾiy�'��I�>I��2������Ob��O	�f0���ߑ4+��%>Ho�L�J�qG�T��M#h?c����%O Tż�3�R�i��ן0��B�ޟ0��ןt�	�?���5����,'�1`CɎu��HiwK�M���?��"�V��<�~W�D����i��K�@��$�t�٦I���S�����ҟ0���?��Iߟ8�O/��A��G� h��EfX/�2�˔�kӌ\�P��+H1O>�����h]趥�5L)$sg�1t��`��4�?	���?ѵ�YH^��u���'�r�;�l�CÁT�aS"�Y�f�Hb�|zrac�֟��럨���ӣ2j>�(TK˭�hU[2�:���,UJ���$�Oj�O�!�/�_�>P�ɏ�G H���Sh}�e�K�����O����O@�$�O8��_�w�lub⏞ V�[�`M�!"T�QS��O���<Y����?Q�2�bM`e�.=���`������9�׎)�@�'
B�'r�W�D�� ̳��4CD'�nq��Ty�\��Ȩ����Oj���OD�\#�ǥ~�AgԜ,���`�A�;��ʡg�G}b�'Jr�'�"�'����P>�	�9xɳփ�RP&����_'D�Aش�?�O>��?��j�!o  $����B�-}H�h���F���}�����O���x����D�'@��CO���
J:���>b��r�=���O4�d_-[���'����P�DaF�,Q�)7n�oZVyBC�֦Qگ�L�m�'C�`3��8&�<�(7�\5t�H�޴�?	��d���Fx��b�Xt�	q*_>>rP�� =�Mc��3W ���'�r�'`�de$��O�j#��V�p`S!���9��[4����I��3�S�O�"�!&��q�D�R�B�*P�JY.+ej7��O����O΍ӑ��m����Ic?� J��0��Nb�t�֏�wz����Y�1O����O4���D��ۑfɾ����dd 6w��n�ӟ�����M���?)��?��_?���^���f��1�0!%�G0iL�'�,q�'8B�'���'j��'%�@b�LՕGs�ŀ�=ܪ]��qӂ���O����O9�Oz�	H�!�rb��nU`�5�u�Ԍt`n!ϓ�?A��?Q��?���Zl�9�x۴0�x��̀0�%f�0%���2�&	��M���?���?	����d�O�,2U4��!�Co��A4�AZ� X�_�Dd�&���E�	�������P�	ԟ䨅� 
�M��?�b�a@T�9�L�
2DP1���p�6�'�B�'���c`'p>���x?A����y�ʭ 0	�2.Dk�l����	�$��ş�[��Z��M#���?���*`��]��k���\��C2.��8����'R�Iҟ,S"Kx>Q��ny��MK@C +1�Zdk4
�%} �<ۀ����	˟����E#�M����?!�������?���A"*�(9X�xj��$��*�X��I	@�$���X�����~5(ݹ ��H#�/�(z����1��Ʀ�&g���M���?y��r�'�?���?�v� ^K��c�M�kxH��f�,ܛV��(~B�|�O~�Ob�n	$6-�
g�5e#�$Pb�H�,T�6��O���OD��e��ܦ��	Ο������i�e��,�}�p����],Th�2ejӔ�OJ�	�9O�S����Ɵ0��e�H�:�е�O(q�M�i(�M3�Q�P���i�b�'/2�'I���~���%�@}�A�֔52�	Io�-���@4Z��<a��?���?��A��P@J��\h���%_䰕�qD�6|����'B�'\��~�/O���E Fc^��T�D�����cX� 9�q�7O����O���O��$�O���6	m�5�h`#��ʋ>�h�r�ҭm��Y�ش�?)��?9���?�.O���`��1�BL��n�����SO5v����'�2�'q�' ���J(�6m�O��d�5k�гFKG�N��`$�_��Um�ş��Iٟx�'Ҏ������'����/v`|��D�w���J3_�v@���'|��'h2,ܹ{��6��O��d�On���,u���
����a���-Z�|o�埤�'VE����'C�\>7m�)4��Bc��*�D�8����?I���?�t/u˛�'a��'�$�O�r���S�XHM�;@իd-فb���?A�B ��?���?)���O]F���-��Ô�̖X�~��ܴw��\���i�2�'���O����'���'呂C�="t��!"m�������}�LB���O��d�<ͧ���?�#�Y��~��!&�5�0P��'Kٛ��'?�'����F{Ӽ�D�O����O�����Q�0���LL�;lJdv	*p�i�Y��₇s��?y���?�0M�J��Ɂd����I�vE�P����'M�iHv vӤ���O(���O.��O��dؼz�`�͋�}�����c��	.	��Ο�����I��O������Zs�ZEwa��d�"4lF�Ԯ7-�O��$�OD���u��Q�����p�"���.
?��Ys@�'M�kA�OB���O�d�OH��|J��W�.���|Eƌ��"q �����!�(6�O��$�Ob���O���?����|B2f^#M��Ԩq�h� �jGg����'��'v��'��^�79�7��O��D�9@*Px�6F�~H��"��A�{j�oZҟ��I����'H"#����d�'7����x�B�q��8t���3�E�f����'U��'��ҟ >7��O����O*�)�'b��&gO�0��r�QE(�m�؟�'����+���'	�i>7��g�r-���5V�h�@&�M�IG��ٮM�Z�d�� j-�d3��څH���r*�J�x� ��K�T}��(�@.�֘�0(Q��v�R��?��0�郤(��e"1� �7�X�I�
�^�Fz�ρ+r��|jF��(W<�W\��R׊��s2�(2�^|R�aE��#c���Zp���<D�H�$PC�tl��$H6+��}s3����Ftۃ�D�f0n��h�,��h�mO03�$T�F"C�
�~-�����ϞԛZ<��CР�~��BM���Đ�K�����&1].�i�ɀ�Q��-����?����?�Ĵ�:�d�O:Ta�&�" 圅Z�H@0-��*�O��I�*�O8�|wi��# i���T��~P`"Q�a�t)z!�Ӷh�b�m?���&�|�{�L�um�0cufӇ$�Y;G���K#�O�!�퉯+��lk!�*g��0�A9z�B�I+=���PD�=G�D	�J ,D"�I��4���O�H�轢�'�E�
ŭ��
8��vM��x�I����0�n���ß�ϧ"W:��c�3,[�1��,_�Y���#f�2��C��V�Y��ń�	?=�CIP5G�%#'$��+0�V0P6P�S
ܩB����D�(<"�'~x�ÔkO����V�wgx����	S�'ݎ�ӃoO,R� RBB�c��+	�'�\(�ê�"U��r!�J�)�H�'S����QO�,o�ן��A�4F�M�Ht�#�H=�1NL_���`�'m"�'�J�����(T�K������T>���9\�@��V�F�V0���"%$�
=�0�S	�"o��9����e0rU�B
 �ڵJ��Ĝj�V��bD��A=4�K�NM#}��0M>q�NM⟼;���X�t ���>S�b�S@�?K!�d�+��(B�[\�zt;�.�}�a|"L$��%S��ID1`�B0q�	*p����Lo�ʟ��	Y���*G*R�''R�� �8��AS8.�J8v&O%��cB�'1O�3�>��(!��=SV��ʏ����㍄	�O?�� ��JQN�>%
а@��7c ݉%	
��\�$6�)��|�q	V��@�0r�L�H��B�N0D�0�6ȉ%|������y�t@��.wޑ��z\�5Z�_Z��2ʙ�8����?���U=�JM����?Y���?1"����4�j�+G�@�D`N��'&^Аb�O��c0�s8�L����=)K"q�Hˠ�ѻЄ�}�^�@��n���K"� 1?��3ړbɼ@��I]�}���11��� t�O�
���u��T� *X0S-hq��?6�Xp � D���`Z�L�>���/��.@�e��HO>���B�.�MS�i��#������R{���d����?��?���Vs�m���?q�O<RIJ���?�p��Z��#�B�<py"L�Q��X8����<Q��(wY:��A�M�00^��
MU8��X��O:�m�0Fw�h� MK�2�v����`P�B�	7�����ӄؤ ��m�vWB䉾gK>i1��|�u�_�gt�I���'�4m�$
o����Of˧H�� ��ꍆ}���QL:O
�Ai�FF��?����?qԄ�dn$�aL�*nX�!���<z�.$�H�0�ʬ�Ħ4mQ�\�E<L�n���Ը:��|����(Wy��gϸK?�8��A�	��������*���_q�!ҧg�]��eP�-��l
(3�6I	�'�$�aB-�
v5K�e�#��I3	�Qĉ'y`<5��'��ɱ�f��p�'	�Hҳo�"���O�ʧD8l����?���O^x��oUw.��W��Y�2ey��	����DC�p՛T��
~~��{���e�ҥJ?"�~ah�P% ����aJ>NHB��ӝ���{CM��>SD�����wj�2Հ��y,=Qs ��:K\��A-Sb�r�N̖�䧈*OD�A�M����!��r\~}!�"O4��6�݌+Ahd�a.A�9A�	��HO���'ı@���9 
^U�G��E�(!D�'b�&�s^bu9�'q��'y"�n�-��ޟě��J��0D�>3�R�31̭�(�%5�O$<"�(G��
x '���l�W�O<�Y�'�����&�M��X�""�+L�D�'�h�E�a{�;a��;p'�'q��r���Py�PU)i�-�<�'.M��Dz��X�\��mZ�{����$]��d42d .T'2���ݟ@�I矐X���۟��	�|*vMП��	�X턝��hI*�8!���!E����D�G��I3w�^d��Cn@�H��r����De���'��
J#Ҍ��k��9܈:r���4��'<"�'��O��_�P��W�'T`�G�2��B䉙v	�!s�u�dq����MQ��ɍ��D�<id˜�0��'�BY>�)I$Kr��5#�9�.�˓�����h�i9m�͟��a	���V��<�O��:!�ԎD/j���G�|�\9��$]8t�C��ӶЦ��àL�&�8 A(]P�<������F�l	�8-R�)��od*'��y¬��{'����������`�M��0>9�xҍݍrr|���GָrRb��"�y�F�|f6-�O���|2r:�?9���?�$�ל^f�U�v�U�. �k��DU�}�f&%T�ɧ�	:��OH4�vQ�O��P*�L��nD�����Y�����,@|�)��@�Ō-�����`i��w`�]^���I���S��?)��"fB\� S$O?Y<Fm����R�<�B�O��1���S4��|�RLCN�'�t"=�O�HM��/�!_K.��&���^���j��'���ȆX8ā��'����e�i�����t�E*��Z�e��u��ϊ|
n��X����_V�XͲ0�v��q�^R��^x��}�G�B�xMsA��$|�>a��@��~���?1	ߓ49�0"���w9Ĝ�Qh�8����A��eY�(Z/6�ܪƄH6-	H}�S�)�'iw�9!��ip��+���v�I�!�:d]���'���'	F�zr�'���!RD��AAԴx��	вm��L"���^�\@���=�(�h�$��i�Us�Æ=lL\���O�?Z#X��Dn�=c�(Jq�K(�̃��IS�'��m���w(���k��KefZ't�m��@ �y��ͲE�T�sfɀ�*��������yBa�.bM���痌pS���t+R0�y"�&�	5s�Ѣ�4�?����	�����j΄Xyu	^$f��2n�O��D�O�Y��O�c�ʧ~I%�A�o�.�ʑ�Y=^��mFy2lѽ��6E��C�]�J��[���2��I/!�>���M�π :���+�Fl�$�ڠH��"O��iT#5<T�ʕ����^X�f�'�BO:��G��`�
|t&�K�h�04O�a1bj������ߟ�ϕ�N���I�<q�k@
2����l_�1�{ui�N��	��X�2%a�e�+`�^t��b>��+j_`5�1Ǘ6T>�4�TM�J��#ec�/S����E��|�$]��p�Ͽ�	ǯh�
�� +I�6���%L��1�r�����?���?)���'�^�ҷL<�"�«3*�}r�'���'���� Fb��A���Kg����m�'u�6z�N @'�ơK�6���d��,XdM��ş���}1 ���O���Oh����c��?�4F�0�e�ƞ6W�.�
��B?�Ҫ�x� ��I�7��5�3Iڌ'��bO��,9�(=�O�=��j� @C�@p���#`4)��O
��'����3H���Ó8؎�Q��X!�NO��0bt!�8c�p����ÚQA�Gz��I�>�@nZ�t*YrE�T#�p���@1U�RP���������{C��ǟd���|��M�7������)(>R��=~P�̨tlݺ2Wz��˞X���D�C��T�"�L����q`-�qS��� ��l�;���<�@E�C޲Y��%�MC�.��{v���GC׃Jb�Ұ��C�<E�F"kd4����SE����D�<�A�5��}XJýEM�	���I�<�d�$�$`$�oȟl�	R���Nh��Z&���	-x}
w��2����4�'��'g�2C�'b1O� �N��G�W(c�
t�GmF�Z� �<����Y�O\v����E�������[���uX��+q�8�OC�b�*(e�ó>�C�I�BH���\�����4b�#����$�X�	�3�6�r�в>�ք0��@�h�T�I;�r5�O �Ĵ|:熞�?���?eb�2�JC-�s�z݃!��<YdȌ3���4$��J�%.�*��b>�
�=ۜ�sI�-x��<��:7Ơ�@��8��˴��+�0�)��H���L�X �$� �>�n�#*�|��(�	<�M�V�����I�<����Q�H8�S*YW��Iڄ�m�<oTwD������G�xD�&X^�'&#=wW�;W`�:p���O�'~�I����x�I�|����A�ݟ����T�	��u��'��IX�� XqR�.6l�����~r%����>Y$`U7���qa�?~��D9E%g?!�΀Vx���AiG������'��������8��O�<��>R�H��ԇL0��=`��.e��B��R�0�G`�\p�V��G� ����\�E�ش	�v�A-ɈJ�J�S�M`\Б��?	��?�Q�H��?�����$f@�?�� >p��`��g�P�(sk�!��o�˓�ȜWg�[��U��"����Ɋ"2 ���O����k�#r ��*q函aRBS"O�5#2M�	M���+Ճ\#���"Oh`����w�Π[���>�<%�>OP��>��h\����'�r[>�+Y8�\rrHV�H��q�#�2ڈI���d���TZ���D�S�t�V�|��g���U�`)���(Or}2�Ӿv���G�μ_�D1�1-\R�<�%���@G��Z���G'�4E��q��y2N��9�)� H9# E�Ug�0>���x���g1���pj����H�GE�yB��d7�O�D�|�d'��?���?�S���@�Ю�=OrX{B/�=7Rv}!�������	 �yy��Ѷ<�,�7N��:���9���N�������(�|�����T�Q/�_��"@�'�,�O?�bF���%>�6JQ�IuT!�d]�\9�p�2��?1n�	��hO��c���?�rCתZȄ�')C�D�\1:d��؟�ɼb�<dФkT������I!�u���y7��e�	��`8Iݦ�(�h�/�~�iԒ+��e*\O�`I��ูŎH�X�a�Oh�Iń�@)�8��I���%+�B٨��d)��P�2~��	0+�i�I��Mkr���,O��<���M<��@� �]�R<��EE�<��K�3^����@�rj8��h]�p@��ؔO��I3{n�|�I�BY��Cd �����n9��	�$�IޟL�v%�ӟ��Iڟ��rh�?Xwd��ߴl<l|�����"��J2����I�)0�|
@��)?��Y��F!@eࠥˢڂ|8�ÄB�h�y��Y_�'�Fh���?Q'Z�$p���ø������8x�'��'e�O�i�O� ����+5��ĩ�-�8X���"O:QQ7�Ǽ^�:y趮�0tFZ�0O��o��M{*O��0������ʟ �O�*�م*�=N��C&��6f\%"�
 [���'�b'�9T����&(&x�D�:�H�O�S�s:�Y�!�=hR�qw��g�L�<A4IY��I'��-*�Y�L|R���((�d��k�ك�	�b�'��-r��vƑ>�ȇ��t�6���E@J7����)D�#���_M6 Sƅ�6<���K�&�OJ&�`arUa�5h�eB�����-p�026ɔ�M����?�+�b���a�O���O&\x�&�#C
�;���#����@`  *mq��J�4����0��OԹ����N^Q����Ј��tH]�qd�ȧ�U�F��(�����[�R�v�	��m��`�4�	o�E*u�'_O?��J�la����z�"�.��9�!�D�)Ym
X�;ň��b(�����p�������f�zp<U�6FҚnq6��OTdXq���^n8�D�Ol�D�O0Q�;�?ͻ�9����,�d�`3�ʃ=�ZA�F�+j۸u`�X��*�a�.XX����U���#E��=�J['�D�xx16
@�@�L��%\�P�ɳ��?�8�Ŏ�`l-��ĂB}�b� �d[��@�|'t��K�F-���%��gg�ލl�?��?9.O����V>8�T�1��9 4 "O�8;��B�:�*dx҂��';�0�pATL�'I�Jw�'��I� ۦly^w�L)��$#�&�pAN9#d*MS��'��'�
����'��"<�P;���.��d�|z��S�W�ݰ�ʎ�4?���$��%3�m�b��a��B�ϵN\8sa�"��1�B�ŲP�6��#�Z�6�OU��!��
34�t X�?K!�d��[����Q#�9�Y$�҃|�!��5� ��G'�L�ao�2��V�.=�=�ſi���'��S��\a�jޯ �<�s���=N�>u�`nӟ��I⟜���:���`�h�50��K�S��և���p����<#6)���(O�i�7� �2Ǜ�)��౳ų[��a��e�-x�`;$`�����'&�0�lI�� �*��'���O��n���M����R���E��Ԃ��4:��!���'~�O?�	�PW}��j�'\t�Brf˻�����m��9�ĩEmW)G����6-M=Jo��I&]��	z�4�?Q���I�p�F�D�O��"���z�QR�y�W�*eG�<s��]��EHF��N<�=��|J���5�0+u�R�t�1�"�M�'�!c '�`7��2��W�DQb�S+1F���K�:����~�]�{��R��ĝؾ���#��n�lu���� �<E��g�ur�D�
fU���@�I;-m6m��x���S�^ ,����9P�huDx�-��|j��b!�̵n���Xׂ�5������?�%L�i�mK���?a���?yǲ��4�(�2&X�739��NB\J<��B����Ŝq]���7�ʪkB��ɴ7��k�cۚ;^�`(�b�x�@�j@F�",3n�!�"�2�$�?��r��J��Ñ��dK,s�h2���7���@*��\����O���d�JX� �r��$b�*��S&�N�!�+�h�"��)W�ɔD�'m�EEz�O5�'�t���u�%�F��`X���ʴOC
���M�O����O��$
��d�Oh�%x/�����Vu��e�V�:�y#�%¥#2�n�>eS
�A�J�����A�g�	^�AG�	T�f�fi��{�T���g�tQٖ�Y� �pk�O@�o�F"lr �C�,�v@��[�O��C�IE��,��#�NHY�n���B�ɽru¨z�#�_

����ԃH��I�MK>�\�)�������O��Uq��� ���M7����N��A3"�'	�3V��\�E�>��t[vfA� �T�&��[v�?~� ��W`��H�Gy"�%��#�+J���$f׎*���}�U�0�F W/�q��j�?>`آ<�3��ğt�IR��Do=J��G�`x��n�<��H��?!�yްi9���%8��L�9
��؄��;����ɑ�Ć5C��X�U�V�4�x���]�$��@�$H���'@�Vbft�7�Ȱ3�Lʥ�\�Gl�i���K�m]D��1&8h� �T>��|��HBx��#)�N�~H���v+������-ه�M�\�P�S��?���n����N0��i�$�2J�X���?A�O�Our^�p��F�XCZ��	�m8c�+D�H��N�:x1F���/��r>���u�*�DG���	�O�D¶S.>fy�Am��|���Ot�Dְ!���	��OH��OD��[غ����?2��Ɣx�h�v$��WύR?!T"�Wܪ0cs+'N Z���w��AP6���X�F�z�U�H�DJ)N�x35@�"MĈ�y	Ó-D ��@,�	s��9B*ҡA�U��arL��	(�M�C�iY�O��O7ȱ���הNY.�RDF�Wn����� ƬJs�B�*$
"F��"�\[��U�'c�듿�D�Ψn�EzT5�wj+J�PS'i�"G� ��ퟠ�	�x�g�
ӟ��	�|�eNOFp�P�cاm\,daT��`iR��g 'b���#O��<��@�5�,���~ `�h�J�;���E��O�Xp�$����<�E ݟ`��4	dy袍W�.~ T{eR��� ���?����?���?����䧉?�D�[�f��g��X[��l�<�2A��g ���� Wrp#�oM�<�_�P�'��B��v���ODʧQ� �Sfd�$U/p=��a0r� }��b��?���?���݌}-*�y*�6�e�9�a2�0l����F�I�X(��'�/ڧ]u�y�$`I	W\uH稈[�HEy�Đ�?�2��*�>��� J&3	, 2&��\�>B䉯aD�%�G��`!�L��
޵NN~����Z��)4c�<��bZ[YeÉkvv牓J���4�?���	O	���O��<��ȣ��������Ҹ9�PܚSJ��q��H�c�??�O41�ҏ]*����/q�:��J֔A�V���!�
���k$��"~�I�T�P��i�Q/^L�B���ӥ��{(V�D�h�)��8
 !�jP���E>T�,�&�*D�����J�R�ѧ~sh���HV�'D`"=�OF��Ǌ�Wj�4��P�U2����'���ZC��Lq�'K��'Kb�p�u�iޅ��Z9�J���
2c����lֳ�?�H"	�`ReI����3ړg0E8�(v��U��I�X=��
��'�Tk�oU�^ԡ��PuF{� � k PhK�Si9~��O��~�[*�?IV�i	�OR���O��M��@[��\�||�t���P���2Ɛ`R.Y5�h�$KG�Wx`���	A�U��:�m���MӅ��A��µ)�e�9Jc�Ԅ�?y���?���*��y����?��O�Ή����?��H���HąG��"To�B8�0A��<c�M2]Dy�p�[1q�0�t�]|8��Y���O�\o�
u���r`^�u�t�#�M�8QIdB�	5J�lR�X�'���1/K>�zC�9(1ǆ'�v�J���I���'Xa(1g�j��O6�'E��&%{2P�Օ2<}�uŃ�?���?���,�?A�y*��1@�C�xw�8�sF�H�ཹE�	
l�Z��I�j���;Pʑ������F�|�'kl�{��f��>�@w�܇0�a�6�N=1Ȥ %m'D�в�f��~�v9�5��}�dHa�-$�ON$��BkD�lT��L
J D�鵌`��Rw��MK���?,�"0u��O��$�O��1lU�Ap���3"&	7~�ca�����!�g/�|Fx���f�0�߂���Z�]�y��Ye�_�S��?)�(:0�����
�a�a��	�����?����?	���'/�Tz��J
��@"�Y6p	��'e��'Ě�
 ?J�}"�Y)Xbpti���q���iP:miRh@=+Āz�#�I��$�O�`;5eR6 ��O��D�O΄���?��6(nT�G��:Jb=�6jE�F	�(��'sDɀ��[*x��@��	��O$���&�JA�Xw����)���|�<�ׂM	B849��i $�?�����\a49� K9�� Ti�B?1��	ޟ���I Y���uÓ,�z�r��%	N�C�I� ���K�Cvr,{f�����-�6ڴ^Y����^�5(T}��j��?�r�����?���?A���?������~���]�x;2/ͧW�Ij�M>�����˖�p>��7[J,b�I�[_���Úwe� "d������tt�v�l�ʥ �,;j�5��;&�v���"O,ei��ـ��e\��d�'"O���福9z5M�5d�4��G6Oe�>��]C���'��_>U�p �S��-��q������Tol���I� ����5��DUj�^��-O�(~�@�Ȣ�D�,��\�e�W�\��<�׮1~��Y���O��1+e���8��*�e�X$viK�򄗷D��9�''��aSC��8�`�W���"	��&�h S0��e��\��i[�1����I:��wv�(#󫈣l)j��"�Ȁ��:/�$ꆲiR��'��S9v^BL�IΟ8��=Z�p����a`�c�B�����W�J֟��<��OhX�tO� \��pk.[�չu�F�|��#<E��*��u��	�G�^��$��,"�Ģ��]��?�|���'�F���aR(t壣�@$��I�'"ebFD8;��x�@K�3�i�����K���� ~��G�>a[Z���M@ K|p���ON���h�t�'�Oj�D�O��� ຓ�Ӽ�q�Ľyx�Sv�]5f�@�Y�*E?2Œ�k���e, LO�L��o �l�U��N������E�Դ�&
S�X�,4kco��5�i��h��O��3S�]� �<!
uL��$�Xj��O����'����Y9^��Ex&�ư�j�B̳7̉�ȓb�*��x)h����O.~�fL��)�'O�L�iHN��UKZ�#�x! q�ՒSo�tJ��'�B�'g2��=bBb�'��i�e7*a"�"�z���@��G���Ѳ�F�:x
���*��p3���J!Nn=�q윙T���e�3L�=���A`jŘ�CI0<�G�J�'��"��U�Fe�"(���ͦQ�|�&(�y���$%htp�
P����fț�yBbɜH����c��{>���Y��y��1�I�T\�yܴ�?�����i5m��)��˛{�"1��̇5TD^D�%��O��$�O\D:�bI�HRl���JH�*��2J�h�4a_���IGoΚr�n���$��(O��rg�����iΎD׆p���~2b�Z�}2�i��	6!0Fqj�CI�'�6����h���g�={t|a)T.���BC�"O8Hi��ՌX�n�p�K�*dݡ��'�4O|T	aψ�#;��*ԬW7n����1O2�2�������ߟ��O���'L��'�	��@T,_DYuJľ	�^�`�(+k����L�vҜ\��M�9fcB��'��Ͽ��LJ"�#�Oݣ&�B5 f��x��|�g��U��%�q�YFS���T�+���M�Ft&l���œ^M:i�b�h����ٟ���֟\E���*V�Ј���A�~̪S�%&Q����?��g���6nQ�$�|� +�^��9Gx"�'�S��'D'n�2����ժxԸr�]'�'g��
��'V�'�r�'Һ�]ן(�I 	�4��קL,��a��=;�^�I,		���dN�FB��w!4=�����ȋ�����=}�}2��L���i�lVYwRؑ�E�~2MO��?���'���$�#JXA�" ��-��'���qw-�e6���|g��PCF7�S�O�Pܫ�hӆ<�0��:��L�d��W<���gb�O���OJ�DH/K+����O(�S�aUtP#��E��T)�#��ŜmI��<8/��B4��	 Ulx�
˓Z����oB� ` ˴o��"���)N8�8�,8l�Z5�'U�p�c��E��04���H�K����	�2#=���Dd�K���'u�����^!��1����a��a�� ��F9V��B}�P�z%���M����?�)�b0����X@�W�7h& `��A�ddf���O��d��Q��$HG�˞2��S�DKR�)��5����mX� `�I2�(O��MR��b前�	�JHd�H�+C�6�@Y�B�Y�BQ��
��O��}z�:=�>��w'N� U��D�W�<���H��m�@�����cW�[H<�d��J��i�:��8��_�<�c ��c����'$�\>�˂�˟��	��H�C�O�`�!v�ͬ}�Z��ւ� �"4�	Y�S����\�D����PoMP[��HP̐c�i2G	7�S��?��$��n(0�ݛTf8 �	C�nJj��bɧ���l֦3��saQ$.k���DY��yB!��2�@��#� R���2�Ȁ�O��Fzʟhc `��9��A:��C�N� �j���O��!z8���Or�d�O��$�Ӽ�5 �U؈��Ɔ �,�q�� {?1@�A"J��g�D����͑����Գ|G�8U$��9����4x�<Tە�-�x3�?�=����5\N��*��	@����?����?)��i��7ݟ�	���'� �8B eaρ����GF�.�y2�ǻ|"ȠR���b[aK�d�t|�#=�#Հ�?�-O��!��Ϻ+���>���j�$��T����:�?���?���6��{��?1�O�H�I��?!�$�/X��s���hH��9�A�t8�<�`�<AF�5�,ɂ�����p1Ge�m8���D�O
�l�%V�,��6F��8�ؑ�D(ORC�	�0�\��a�&$Z��Q��ƁzC0C��;ojz�Bv�$k�c�#�,�I���'Ȅ�tŦ>y���Ϩ$Q\��1�T�����êw��9�E�OD�D�O�c��%|�d�@�Jm��U��t�ԮF)Y�D�����G�nl��/���(O��9 (K2I�����u��Ԧ���i�)���d�K�ĭ�&Ax���\���G��0���@�)T&���mRC�xp�B���y"�'��}R+�M���{f�؀4(�pv���0>���xBΫ���p!�+-��r�Y��y�E
%�7M�OL���|Z��ؕ�?)��?� ��h�뎼Ķu�2�A*bֈLA��Q�&�C�֮;� C�KD�N�k�&1��c>����n���O.*͓�ի ����o
(�&|� Ɯ$��!§K.�������w1�8�T���E�DmC��]�n3�U��Nq�a4���O|ѡ��59&t	#&�W����B"O�qX"+�X#q�gBW�`T2���3�HO��MB֠�2���1��H#���6�u�	�\���H:P��5�	ן ��џT+[w�wT=i��<;+`E(� Wnx�q�'Q8ix
� B�d!�Q��x��%���4��t��	�~�v�2���
(�Ja:`l�e���I�u^�D�A؞��#�\X0$�6ƒt�J�h�<D�`�k�
��e�O3j�2t��Ǚ�HO>��%��M�D+�L����I$%�U��ʂ�?��?���u�~���?��Obr�y���?�UVq�9��Lp�"]("BT{8���'�<9�N�!�H@ʍ''�H���~8�����O�l�,k�m��m�2$Т)��&׆B�Ɋ �X!�͓�"��q��]��C䉪(Yx� e�~8 �eT9<9��I���'�>����kӎ��O��'T��2�&`�i�ŢQ&/��@��`��?Q��?q���?a�y*�leW�X
dZ�(cW�V�}FQ����B:�']�hI�F��=er��0�ؿ&x�MDy����?���)�:�����EL:C��R��#A�!�D����E�>��vT��0p���'_O�Zw����H0񵯀)Viܰ��3O4�HElDӦ9��џ�OU���'d��'��ᡤ�	Z�$�br.��B!���j�(.��T>#<�S+1R��r��Bm�֫X�;�������O��[���'r�S����Z!�4F�'�f�d�)�� �ꎇZmT����/h��酂)D�t��$��m��Q,E
h��I�dF�̲���?�A�T-����¤krR�zV��џ(��>&�TT ǁ�꟨�Iן��I$��9����d�}������I�zw�u�OV`��Q7<�{"��+rDp0��C��L4�<�c�'k^Y���I��=�cCza(���b�s�ԁ�� 
�?��R�?q���?�gyb�'剕M�F�we�?�d��)�5>B�<9sf({3�.�,F�">n�4h�����~"S��Ʉ����ugZ�v��p���t�Ȅ�(���'���'��e���'W<�fȉ$m\���%��[�lX�D�գ�s`$M��H�5y�fA���'��;Y�:ݚ�IZ�j��	@�D5Uz��0��y̌0�EPY��T����Of�nZ��$��F�X�x���g�$9�B�I 2L��%n�q񘸣��Y��^B�[3(�0q�78��#��� �4扷��'.����>	��򉖉"�*'�Ł4�6�kFN
H`[���OB�d�Od�W盪#/�y+V����T>�����2zMRB��՝+�PBĪ=ʓm�>��)Imܠ#�n8�S�~N��#C����͒��<i0l韠�۴*8���۵d�ZG�X��O�D `7OZ��)�Ot�EeI9=��	�3"O1�F���'�tO(��&d)OJ�<��̾)�2�3�?O�PգKߦ�����D�Ogrm���'�B�'w`I �af$(kw�шu�H��v�^der�T>#<y����/�d,�v��5'����	�g�Ҽى���O8��2jӕ>~�x�և>x�+7���/�>�d�O�)���ЂFGtAXR��.c�𙨶�5D�� ��/!�xBdd�'�"$� �%�{㑞�' ĸqj��T�v(�5�X�%�������?)B�	�A^�S��?i���?�%���4�b�'�5h.\��ګ�Є���O ���>)�,��u���Hб7�>�rG}?!�i�Vx� � �O�mc��2фýO�`�-��p;��O�x��ɝC���h�6uz
8�GӦj\lB�I+*�~]�qeV����d��_<HY���8EN���4],tp"�$R:�,�z��ؙCXʘ����?����?����*�?������*Ղ�?��h
����FT�9�0�gkQv0��I<r@�˓g�fHK��5�Tx��ąs��I��č�E�v�Cg��$*��_6n"��!�2D���!��?<ZB�����]*q�/D�|0�!T�W�^�w.[�7[���$b����}R�w,�6�O��d�|2�)6}6�Q���2RE����)-]�T���?!�$f�-������� ���)�L
�	��y?���f前[�~��Ǯ��h� Q�ǗJa@	+���d�'��L��;i�>I�á��SM�u���M�GN�9�e.D�`��)2��%��J:.=�|�Ҧ-�O,�&�`�#�^3�8�����uݪP3�m��(���>�M��?-�Z����O���O�yV�&J��A�!j��>���CW�
,w.�}�IF�t���'�n!k��]�E���t�	"lR�D�R�/v��c�}�P��u��*���F���f�B9� ��X>�%j��2inX�h�	���?a��i��7M�O��O�i��?aWM
�SbX��*\�$X�H�����<�����>�&#�!�R�z��9 i��Uk�'��6�@ͦ!$���Of:! S��-_����S�ҡlhԼc�'�RhL�������'�R�'�r�r݉�	�����I�)Q���q�+E$9��i������[��"�O^���4d�6�! �+� �u�O*�2��'���T�ě|U�`��I�#䙈�'!����FOa{�扣"�nRf��v��� �U��y��G$��4"Ypb�W�Z&��"=E�tj�	\h7m��>n��p�Eڬ`��q�TcݙU7����O6��O~D(��O��d>=G%˝rUɩ�͕LZ�;3ß't� HG�E#. ��@����<	t���-f��q�$�"mpXHJ��%iƌ��J�;q�ޙ��DO�"�ayr����?ѡ�i��#�e��q�Mۣ��3i�BR�'A"�'���'���'��O����5�JXb�-�7�^�٧&�y����U9B��+�$)[�o�.�y� �>�)O�I��ɦ}��쟰�O�t�$'����Q*\0n3@�3b�_:Ly��'�2��$���T>i�х<C�`���@'%��D·�<ʓ_4�G�$�D�wY��r *G�⡒����(O���f�'�"}��VqFNɖ!��&n|iYc�X�<a��V�Q��� ��l`���`��H<��㓱C�8�
D�gZYHc���<�g�)��F�'prX>�)��A�����Գ��D�bc�`�.�#o�qz��T�x��T*� Dz� ���f��ʧ���?Ie���>����+V1(�JAY7�ӋTdx���i�����n�M?E���r�2�jg�Q.�ȴc�S�T(��S��?���|���'X0ᑖ%��~��kI�6��	�'��yUO�F�ځ ��ɘ}6��ۈ�$Yh����@�{
�(��?|WΕh��@s>���OH�B&[8����O����Oʑ���?�;U�:�x�bM�o�,���z�T�5J��	��T��S�P�Ue*�#&�P6S;@�	e����8o$���sh�)q�칓@(���$L�CO"�=lO�tqkL�^���	X8(ur�;G"O��n�S���t�E�P0\x��Nf���\���k�Ovy��h�iFN L��u��R�i�O���O����t���O�B�LMXr��
�xyJ�J�)��hG�ڤi�����<$�l(��i͘z7��*Y�Ј�aB	y^6��%�M5�r|��D,HV ��'�t|���?Ѣ$��T��l؀
�f�舉v�D�hOТ?i5�	��0DY oʶz�Ĩ"Q
�\�<��9ph4��$��2|�4h2��<�p�i�^�X��$'��)�O,˧
hJ,pT�5@-ecc��q��,��J���?���?����<�H��7�R�xC��S�4E�*l�[�,�=O}�p���(�(O(0��M1`�3���e�'"�HbF���E��&���GyR�Y��?�����O�4	�Uo�!Ѱ���d�j(	 �'���K+�%S�ǎB�5������0>!p�x�nX:dXx9�!ќm�FQ�f��1�yZWc�lBܴ�?�����~���O�d�3Vv�Irm�V�¥Ѓ×�r��y6F����`�	Б��T>I�|����M�GTP���t�P�S@,��#��O�1fǷ|��)��X� ��	�ȡ� ˋ`V��QP����� �	Пt�䧔��J<9�����=	A�(e�Ƞ�ȓj�Ҽ(pbЦ�ڤ2�mۋ�t�Dx�O ��|���A��xBF׫n��}��JVd<x��'�X���FY�_�:x��A	���!�'���"'(Wi	D+��\}�}��'�$�wbտb��c S�#��U�'���+�	��5Sr�G'��q��'�dKǏ�?��ámT	{��Q0	�'���0/�)/��%1�/"yX�'G�p���W�(� H���LL���� ,�S��ƋEPX5���g~�QQ"O�4�O�K!��r �ǉ5w�mx#"OyqX3y٨���x_"O6�@���D�iڥe@� �f �F"Oz@�T�>��b��8�0á"O�}0���0��]��l�	6ż��"O~E����R
B���mQ9f��|@�"O�Ѓ.��C���)Q�P}���5"O���R`[6]qzyxj�3��`��"O\�Q�G�V�r��T5$���"O����O�;�x)��� 
~��I�"O\	���m�H,�a�ߔih��"O���0K',�ȅ"g�[#lK.M�"O8���  k% �!r���Z5v�a�"OH#7ڝ[50�����V���2"OpiN�5�$;A�yƈ���"O:�{�(���ViH$���k�z\�%"O�Qe�N,��4�Ĉ@"��$�5"O�i�!E�,Q���p����"O\�)��gת1f��N��#B"O�!�_�~���Dʛ_C�x���Ob��,]^�����FX���'&ҧp/��)M�+�ڍj�M��+�썅�^}��䪍�"9F�tI	�YW�]�я�.���� ��q��U�T,�hܓuCع�p�M�fRT��[(]�q���Ji8����'x�p�S�φ�!���[��}�C�a�	�{6P�����+�oӟ,�q ��?��D�F Ұבs�%� `�/	%@8G|���( �6�8v�M�� ��!�(�?�G�8S%��ĕ+��(r��%���1QjOQ�H]����W/ڰZ^�~"�+�i�=�͟���s��U0B�D�3(d�h�tG^!@FY�zB=���O�g~b�9��=j3��Ut� ��Ô�f.(��Į����{�ݨ{hq�D):�M˹[!��[#���hTH��Z����'���t�N�ɧ��`��8�3w��� ��i��0�(��QR:8 ���Q�d�s�ȷ��%�m%�l96�/:�}�4�xrd��tc?O�9� ��[.\ Y6*_�<����ǊC��uwI\?I6\�B����4  � ���+02���߯l�L�
�(0џ|�`̊�>?���;3�Pr7fU<�
ᚁ)J��.��7�V�U� �Y���yJ?����!u
E����SF��Hr�55��P�A��B7*�� Í'��Õ� �+��O <{�	��Gd�Hv�Z=�n�'P�b3FòSU�Ⱥq#0ڧ �z"DӶJ��DI0"F��P��7e�=8�4l�P�Y�D�bT�8�f�EzZw���'v��!��ɇ"0�rJE[}�'�	 P�	�J
���!vU��K���'�
(�0LǤ~��%�οZ'*��!��b�'
4�5!���,eH"	��L/^ �',?L���R& 	���E 0@�q��˔p�S���B#f�kl����ŦIY^�-�$Y�O���v���Vf���~"&Ԥ/p|�+.O�T�P`�غ+�C�$�����1��{r��E�(i�]rs��.1����KPN�&���e�)2-��R�d>#�n4�+W���`W�1C��ϓz�b��m�	r���P+��3���zG���9k�$N�BNQ��M�3�88C���?)�� ����:�E�jX���P�a�Ԙ���'JtPd��\�<� �X�@��}Pn�hfj��(q��*cݩk�
T1J�!di�}�18�M�Z�'+@� f
"�ћ�4F/��Wh�',hDs�4�V��^�'�u9�O �ӱ
��K��x!��<������@�̣SZ�cE+J6^�`8�AQ-5��Q�HI�#nz��N
j�ヅZ- �*oZ��AzBI@�<�@Y�c�zdᱨ."$�[��<u�PatNR�3�p��B�v��W�5g$4y�g5n�$�Y�剚L��u �R�L�hX����)^D���['T�:�ċ��<�bE���t�"��a[���	
`�h:�3#삄X�e�8;��N�d�c,Բ�5��+*	�%y�JR� J$�m��Y(���[�3.4UHРE *��T?�1!�|�':v���ꙜF^��P�'B���gO�/�O��y�@���M[d��1���4!Z*^7|)03�5zx��ܟ���Ö 7+��&��,���)9x&����x��HԯZ�p��CȘ�QD�($-7�égx9s�'�� �C��>�£��[64�80fW�m4�����y�dͬ�xDKW��?2��!�wÖ&R���(4�W�4����EZJܑe� ���k�8;~@ ��ߦ�B`�ӑ~e�d�l���'�
+��O� �JaË�OE��
G	1z�(�ӕC���	�PH�0d��3��I0�J�{*�l�p��Wn�b��	4fX5`7,S�nU���G	F�ȱ �T�<�O7Zc����4�¡ �E1^�8m�a�ם=���K'$*����	�&4NP���c���N	;< �W�Fl���(xu��� d7Ja:��'hD����O���GHѯ(w�ׁV0�����?��0�'�J(b�C�!}�gB�#���O
]��B�!?���/��n��tjb(ɷw����c�T�zxb	�ɾ��p�����S�:4�O�Ht�S�? R�����~`�y�&�"��@�+�>[%�F�G���[���ju
O_?�b�أ=����;��]Qg?J*K�/Dv����5E�V�0���TzB%e�I	S!��ʧ+Yrx��yr�)�J4f%�LД%�s�l"�/�<�7IC��� q��d�ڕK! 
����\),��0��=N!C��"Δ���X�θ��'5^Q�?M10�M#���@�E�'�zIB��;�I�g9zH@���4C�5�4��8KT\��~$@�*'e|���
9��	����<qV��),���w�xJ?# �P[ҵ��.&��w��$bJ� D�ʧ"��'�ĕ�E�\�O�B���l�@~��"*�>�qUX�rF����c�&ݱ�5�'�u�J]��?i4��N蘠��IBG��(�)#9��5��@ D$Us�'��c��Q�&�!�̟��|�@�ف#���N��a��(���?9&�AnD�Ct��X�(诟�y2�B�?˓c�x�kf�ɀ=��y�OC&��0I����&֞�=�O��Z��ċ�q�ҡcb�E�=�=�ԇ�6U<��f�Z��G��!�hhQ)O�����UD����
�,��Ax���Zl���	(�A�F�J�P�������<�փ\|#���eԎ'�N���\�j���%�hUV�8b�O�UiG�*ݵ�ڊY�̜%��ٺkO�
���J�ޮ�C� �,�J� ���S�����$ L��,b{�[�ZV��2�(�Z����uߴ�H���U�Xt\�����U|�h���[�\$�A�ѕk���T��F>X�ʧc(�My\<z���E�"��e�e��<-,jղCE�0fX�D��
ǟ<�{?YF��L0�ɣl�X��ƉY{�!�!e@��҃�+(��'V2�52�K^D�ʁ��i�Laäa��}y#�޿vO��r���@S�K޵s:��)sl��r�'P�ɽrG�ͻi{���q�XG�t���D��2M�p͓^G��s�CG�:�T�)��)����<iW�ms���`��y���СU�1��q a�3I^,}����o>��d$�N-��`�#HS�2Ui�ؒFh߆m�D2r�!� !Q�Θ)1O0Ɖ/m��L�T�Jf��0	���oWL%��@���?{���rMЄ��
@�+p�qO哃h01@�!��Eq(�3��W8e\�0���S�n�S�V�"~��`�%`�E����6������-�\ r�.�)����vn������<��DP�S�z�s'Z6�Q��l=-@��9؋K�/\.�Ǘ?�n���#��dTj�@�_�䠋0��g�漈�'P���A�c@z�cޫ�j�,O"�Ɍ}�2q�A�C�E��]�BC&*1c�����cڗ��'��kʷ5�4e�&	;��O����L�x��8�GU)o�(�{����`�%�CU��͓v��Iz,����Z��S�E8P0�� '�I��V�Z�Z@�%3|N ���'�X�h�;N X��!T�X	�!�LR�bq�'R�!���Z�إc�+�>%?WJ.
+@�b�)����&��q����/X�G��3�ˑ�"W������z�O��Y"�O��	��	{�X�a�F��?u��7���#��?�M������Q��?�$��C:�z�p��N�.w�L�v�L:D�0 R9O��vO؄�MK��&B�*����}��S��@b��C�_f��:��(v|�5�F�ʄf��D�w	BK+t�LZd��!O���x���
2��"<9Td �h��ᢑB.|��냊�����Ο��Cǯ�<h�F�p`��<~����g>�ʳEZ�M
V�FD+7Bl]����|ۤdڠh�X�T���[�5޴2f��z��+j�|� 	�f �? i�,�?��x�@ӆ�?Yb#P%)ڸ��ğ���tAM �az��ܡG{\ ��. �*H�֬J3L8�@�qA��S���DO�zM�5����d m���K����g��杼^f�d)�#��>4|ů�P/�b�|	���(����a�Z�B�Q��q�A2����d��"�H@�8gP��9�DX�$��P ��/�qO��i7�Ơ O�
p��<�	NO��k3�ր@�����0����y�|P�^y��P&�w��V��S_���]J���r�4\O$P��cܪA����˚
h�H#Ir���^���(�ĺ�՛�,Oz���(�8?��Xʐ��	�^�A`eb��d�Í�$(��!�6=iƱ�!��ɒP�@��7���%+ �XB��"����Oʍ��$	5kĈ�yD�)2�2M'��2��B�;��t�g.�2l�˓J������HK�h��Dé}:̡��`�&A��s�&l �A+���p&�=i�t�@T�0H�Jҙ0w8��ց�I��sϺ?c��k���Y�r�5G��K�� �&��ɒ�A`'�Qq�IO�T�
�i���<9���4����0�`S�m]^xH��)�Щkէ�A�6t��핧d��� ���E���@$=Yn�K��E�2s�Y��dIK�BAӓឬ$���(1#�˖�S��O���+Lp�`��O��½�%*��}8"?���=Jx]���4������9��[]�X{ @R�0�R�Î#�~��� �
8)�弟��RL�#e��R�YlgT�λ%Y�x�T��/>�JE��x��i��Bmny���E
��ũ�Dòl�<P�Od�q�Qc��E�Xy�ԇŅ
o���JL)$�H�%�i=��q���!5$�8���bw�һg�f��{ϔL�ppB��\ڎ0��阷p�M� t�ʔ����y*פ,�qA��TI�T8�F�9!F�.>�����!��m' "n��~"\H�6LE}�0��� &��K���~>l�;��L�p�D� �p���ެ�y�'��/s�A��``��,ѨH(x�D�M�5~�1�$6�t�$A%/赋���O$�̓=��p�k:o�Q�b씃����j���$���9��f��=��P�o
�p�dଟ�#Q�j��	DN*Lؐ��̙6g���	� dԠ����QJ�hq��'��'��`��%f��Z�ȌR�#pↆRM&t���84���%�D�I����O$��C��-��'*&�P7)GN�hP��-@X
�j�쟰s�O���J�}"�`�ā-��S�?�� j	b�B�P�.|�W���Z���u�� ���^�z�G|"&H��k#�G;MB4�� [�\�#�Y����&%M4�l��].�y*�@��;�u��d�dH��F��~j�����jg*��K\!z#>��G�4�@�P�\�3�x�+@g��<���Hup��4��}Od��f��꟤Pc�k�|��@�N&�����X*�V �2��'���`��������;�u�����5V�h� ��KN�_`8|d�L %��å������0+' (S�>ET��+T��N�cPj9�@���bUNQ����F%��K�(tA*�(��D�#J/��&�Ln�H�Q�T�݄8���]�-R�$�
5���$�	�w��l�@�+��+ ��	Xç!4��]��g=cG�� �@��u������y�/L~�.�@SDY4�>P�5N��r�BD�e�?TE���O�8+��|��O5�(sR�O�h|<!�rH�Q�d<��Gτ8����'��`
�������8�2�%�1C�
�)��>�(��.K�x���T�G�EȔ�z�-G!qRཟ��N�b��퍦<*,%2�*�}��ȃ�Jܼ9��ҒK��$F�T�E��,&�!Ef�0��l��)�;��I1�f����(��A��Qf���>�ǋƭq�j	P&�_-)��W��<#�� %B�Ԑ6��:<%���ޝb�'e��Ã֍_��Kf��&��<�D�G�<���Iٚ$�X���u����'�
��#T��iR#c�O��z��(�)���d����u���G}���"��F���i��7�Ӣ%�A?&f��kC�� h��8�fsӲ�˴��(H�M3G��77T�UpU�I�l}2,!��+S̐c���$�\�I�kJDB3�m����s�[?Z*\�!�$i E�k]��P��I�"�Gz�eXI�8���Y	.}��r��M�&�1p4)ŭ�5�\Pa���P�'�B���B��d dh���
 O}��{s#��$JH6\O��H5��51%���5W�r��6`T�t��}Q��'E�|S�b�'�ڭ;���<�p��blC)
Wf�?i��Y(��P�aΚ�M%(]�5�ك62P�QM.�����D�$b��$Э*p����%TE�%�t-Y(�v�
��(��d߁�8�+�����DO�y*���Q~�����
��4�s��	i
�
^�ዳOZ08$�SP�A�?Q^y�.ImcT�_4+.*y3�'��(O(5����}x\	���8��qi�B�X�(qك�ѵ�M��/jE����N�33�P�|�Y�D[*��h)Fm	S�,bńB�����F�O�T��hN�r"���e $�k#�F�4�i �5�l�'��0t1�LX�Eg:�ї�;B
A�ޤ� pSp��?=�0l����w�\!U@X!�B�* oBK����'&�LC0M@2sW#{���P�L�1�yr [#
���p�E�I� i�`,�*�y�ΚR.�рB_
E��t�u�2�yRK��xGTAە�Co����R$G&�yҧT�m��132��(a$��2�
��y�&��K1��Yum_�\;���/��yBjث���jc�=M�ha��L$�y2�G3C����,��L�Թ2�f���y��C�TE�|�ȥA^*������y2m^u�Y�⌇A�>�;� ��y����4��ĩ����6|��N-�yb�[4j�x� �,�~0��f�y�o"��U��ڕLÀ�q��х�y2��7V�z Gș�r?�$�e��y��;3�P��H�3�@���`��y�n^?b��s�DX�'����2�y�dõ&���u$ډ�eb6�]&�y��T �!�_9Tz(�����y2eR��r�E���\P�W��y�
�L�� ��'����C��yb�~��P;A��)?�Ę�y��8S�p 1���>��ń��y��|�<@�ac�< �F��A/�3�yR��#�&X�3̑-ou
� ����yREֽ`-�ur���~�*p#n���yb��*!���mͲJ �|Iԋ���y��IY�� � ��~J�@ ��y�ET�@6��AʻT'�|���y��B;B����وSt����
9�y�FF0�X�O�yh���6�yB��� �f|�"\F<�w.���yDA:}������}���R���yR��{'\�*�)kԳ���y
� Թ�e �X
�X��^4̊���"O��:0��!A�t��0ѧ��`RQ"O"ݫY%b���%��rv�WaW�<)1+�U�1U���Jh��6�Er�<9�c]�}�a����l�)�Km�<	��?-�ұ0����X��'Yp�<�R*Ø;[4� �2!�"�RHOm�<1��
ˀ="0�(���2�HE�<)��ɏI����f�\=dJ���G���<Q���pe6L�� <	DYtÕx�<�R@(K�>\�.[�W����fi�l�<a1M
6?I�,0���(O��3Ah�<a�k*p�X���\<�B%�1)d�<ɱ�L�2&��:��OPy�d�
At�<���ۥ��		A&W�.؂�!�v�<�Q.�7OWD4��A��x{r=*!��q�<�3�&h%S�
����k�<����`�2P�7��$�
���]�<YS��u#&�����I�@��R�a�<y��?uK&���κfzR]�qn0D������;B׺���(1��q1e9D�@����W�"���@t��x��7D�d�q�ʏ����2���ST�4D��)�E^�dud��m�R4vifJ>D�H¶ϑ�B��j%j@��:�
P�:D�9�K�:�Pڑ�P2q���5D�܈�B�d�|�Q�,�N8��P�1���<Q��8bg��pF��.}��`c�\H<I#N�.(o(���O�<9��
�{�6
O6M)�B�/Uyf���F��RY7"O�#A�</媵��S�m�,�e"O ���?@<�M9RD�=Pu(eS�"OT��ńQ�g�r0���X�Uh�Q�"O�j�� m$��j'IPA*u"O����1	V�$����:ZN���"ON���ͫ��=�Cʝ�86��$O��AD�%wn�i˓*�#�bySVI�L!�¦@� �2�T!-,aCY44ѱOZ�@���䜴7�P�q��W@�%f��yR�� i-�e��E��h�b�zW'O����?�ӓV�z}���<�����'{V��ēn_l�3�*@	9�5D�ܫ(�be��"Oꤢ�C�G���R�f��칤"O"x	�l_�-V�E�T�J+y��aA"O��e�RxR���W"Z�~�tTd"O�i�#�V�wST�Â�<ˠ�2"O�_�`
P��c����"O63�Z�-�,�ۓgH�J��P�6�|r�)�� �l�R%JS#��h�S��=�4�D�O�5j
�0x�;�/˯.�ft10A�)f*<nz쓚y*�V	�gBp*�	�(,a@f	ϐ"���N��S��B�7*���+L�Y��c���M�>��=������@E�ta߇�����J�:��9�2 ���p=9�}ҩ]�P��9�c��I��DkbA�
�yb-]���5S�Ά3�ĵR
O;��Ob#�tlĉܴB�sCF�lR��yr̊�J%�@�P #@�@�.�p�ў�_�'�T9B�/8Bv����-vμ�k�'��`�&&��QiԎ_�i�(��N��nm�'ݱO8�P!��<R5#"ȋh_�Y��O��U��� ��'w�D-B��=�$$�O\4�o��5�,���PB+�l����B���Ɍ1�&�;�jT�@�V)S�B�>�qO@��J�H���J���6̣��������,�~֧� ��1��z�.8B�� �)jV"ON��q��/b.=��'ť(������'�!��5V(�ģ��L
np��3@+]�r<�򤉜�����KS$a(	b&���y�a���v834��"o�u*qΣ��'��{�՝�������c��rȟ�M��{r�$,Op��U�"P���Tf>�X�6"OV�A�F�K�(ܙ���A�&�Q�J��Px2��O�~�XU�$hK�8�&g��y�.��}ܽ��C^�TxK�.ď�y�9:	6�c�R>ZU+�.�y�#�y8�!��K�d�Y(Ǥñ�yB��7v��=��VX|(y�R�y2l�m�<�q��|���Q�����y��Z%�����@Cg��u�!���y���<0i�REk�(jlh������?��e?,O���0�\�D^�"�N)Z���xD"O��DE-X�A�'�	�VkwmKmH<�q�S-y&-����'Ì�cΊt�<����D.�����A2c��J¡�s�<a�	��'~��#��2v���%�Bh�<� N;;�"�KB���C��(��|�<a�&V>s��A�RL��$$���c�<!C��4XX�2E�&���Ӂ�^�<y�c�GFec��N:[���(�q�'Uў�P�>�A�!Zk`V���E��w���ȓ 6‫!�֬�u	R҄)�O����jZ�i,,$Y�ŅXgJ^�0`�U���?E�,O�]iW��~ڞ�q���&?�E�'A�	�]�-{��Ύ�4��E��W1�B�	��f�:���	��t���o��">)�j�,�7��yV�D��A�ppB�	#X.&�Q��ce����M_�QM���T��h�^p��ÒX��P�D��ݸ��"O�Y��ͷM��Db�"��"r����'��	0;���(�-Z��\TCՂ�u�bB�	(N9��CVX�<����ճK� C�Iq͔��s(��D����T7G*����<�F�?|���r�j�,�V�b�jc�<Q�d
�t�L����v����P���G{��	�
	�A҂N7Mp	���� ��B�<W�,9Ģ��4�
'�W�m�fC�	�xh׃��px���3J�hC�ɳB����V�ЁPv$�4o۪&�>C�	�k�X��$�� bD��R�@ 5C�+��})�%�`���ȇ�05�B�	7E�|-�	X��|e`Q� 3Y��B�Ik�:�b�ǚI8�!��vv�B�&Jo�0��ՊW���2�!8C�I(J
0���R ��2C��5g+���3�	r	�8"'��|��@����m��B�	�GV���c�B�*N�h	1�ѝ]֚B�n=pD&ѕ��`p�!P�6��=
ÓW�(a�`�U7M�Š� Y�SCE�'�ў"}:#�)��M�bDO)� �S_�<)�m�&(�W�߱_!z��U\yb�	p�h��Ph6�ޱ
f�4f�<Z
P�� hFq�g�Z�y�ݢSM�2�,�E��S0=4�R�n��!�4� ��U,T��B�I�I�$�ƣ�3T2i0�D�3Q͈�<�c���v*Q
P�:-2Fa�*R4Fy�'�d)�-�G�<�ó�M�x����'��4¤���
܈��H�[F�T��'�2�&J�����'\Y;���  S�	 ::�b9�&�^k8`aCT"O�!�ӉMP�`���#90�@�g"OV�CĮWT�B�r������5"O���,��Cv A9�!Ƞ<���"O��FE��B8��#�Q)H4�U1"O���qa�:6�	H�o�"�0��"O,���@.F�Xt:�~���Rh�<�g+J�`,@4���.y:B]��-�i�<9Wo	�c;r�J��	�%��@�e�<��H�^Lm�r�d`�9Y�#[^�<y$�Dk�`�,ɖ\'�0�4&�s�<aE��+#����s��+"���V�<�&���s6<�i�D-k��w�P�<yDkO�6�Z�Aǭ��]\���TONV�<QT�(8c�}
tN͎_�,���|�<)�a�;��8�C�$f�`U`У�t�<	���N����GY��[�ɇ��=�����8p�&�Q8��-�N�<����*�(���+��5�B����G�<�E��
ѫ�U���8��MP�_�'m1O|�=�� �@�A��7c����O��y��ƍX)�qc�DڷbG�Kg'K�yH��L��E���5m�xM;�"��O�O������Ct�R����F�ti�L��_�����&�����0�Za;�˟w�C�	�$}��)C�4�&Y�#D T�a�
�'�n�C�菷E���D��x�1
�'�ȨY�S��H,��l��Oo4\�	�'��M��F/"��{G��7��iY
�'f�(�玷[3ȀS⬐�܄@��'�}h0��Y�2Q�C���LJ�'�䄡2o�K夠1�4 � |0���O$��G	=/��� *^�S��؆ȓm�����g24���%a����.�@�1��2U\�`��R�:0p��f��i2e�!=d0��GO�h��@��u�v���y�XBL¿z�Ω���JXR��I�,���$��ȓ}e����.��* ��-��܆ȓ��t�DC��'>��5A��i�(�ȓ&��-���G*!�$S�ċ�R��ȓ+C@X����txZ���*� 2m浇ȓ\���:#�� ��X
Uk�8f-�L��3Y�A���	ބe��H�PJX��\G�U�� �2 ��Ƅ���)�ȓN>BȪ5��*�r�`$@/&�>A�ȓl[�� f蔠+�>��6$�+&T��y�pDxq%L��� 3�]&O��u�ȓOO��6�� dlB(�"gI���ȓoF <A
j?����C���0�ȓH�^�@�?�$��!�I>O������ѕ&��k d* iV.uy�ȓ{���@h4n��U"�i�1}_\t��m�dA�g��L�R�yIN�*"���L�@�{�h��gM��@�C��0�Q��*��%AoC�����n�fņ�"s0:T��?�h�S�R�C�=8~�HЁ�Ao�����I�>�C��7�x��ՇuK���lM�q�C�?gb9���)l�h%���r+LB��7�i��[
{2 l�-y��B�`5�1���_�e��}�2L@f�B䉥>�0�	pH"����B ة:�|B䉰}oV�"�b��Q��C�:vZB�)� |���d�D`b  ��;����"O��8�(:"�li��,ºR�ܹ��"O���v�R�M�8DYE0�E�w"O>D8A��[���Ѧ�	!u���"O^�
Vř�9�85yKnr\h�"Od����NE�f�iFb��E�%0p"O� ȉ`5��ե^ Y� �7�Y�<a�뉖[@��ab�9$��$Sd�y�<���[��r��6:e&�2���|�<��(��cW�`p��J1g�0�B�JS|�<���W]����E�X�z)���ŮNq�<�/M�[+ ��'�*u���ISp�<��Df~)x�d.��� Qk�<QQ�U�J53pLR�l8��0�f�<1u��p�H�7(�"j�}����V�<1T�C�O�����"g�
i��S�<�b�+d��s��ǝ/�5	d�L�<i���?4�
�����$I�<Qv�Ԩu.H��%�d�x���C�<Aň�(�~(:��	h�ڠ kMd�<yE�
gJ�*�)[@2��F�a�<�W�^�Y�nܻ�I_?+�(����Ba�<)�"�6)���)-��B\���Z�<Ad�P�S�pl�@<5��u�P�EW�<���;��t�W��:�x���n�<yըn:F$��ЪM`��v*�P�<������#�ԠO���[c�Qw�<aU!��Y�X�[2��B.nHs�/v�<�дer��(D�[���Th�L�<Y�� D\X��ek;>�*��LF�<�cP�ݩG(�-'��bU~�<���>�v-p�hDzj!�`��`�<DmY�1ʁk�V=kw�Q;��_�<	iX�|q:�%�CM����`�<�Af�(��*u��� �� F�<Qb��+Jl4�� 	�&3�VP��f@�<9�� g�|��6�H�\̈�k���z�<�Cʋ���`ыH����A�Pa�<A��Oj#ι[�_��P쒁L][�<��"A�iC�b���^�0��U�<1!ܪ7�Lr ջQ5y+�&Ff�<�V�<q�b)��j����	s'�H�<��#�	�L�X0v�vX�W��B�<���d�u1�U6p��En�}�<��i�ǀI����i��/QB�<�@�/p�j4h�%�T���<1�$
�dM�&���d1��`}�<��d
�T#�;-:����]�<���/I/h`�sQv��xPǤSR�<iT�3x �8R��.]���S��S�<)H!��u@s�ͪP���N�<�0�ב�ȕ%B�x�P���kG�<9%���<��hD�Ϣ zR؀an�]�<l���&a{��%S��Pb�GX�<�Ã��o���K�8� -�S�I�<�7�V�h�޹�r�V+�@���'�n�<Y�*I�nL�����ӯ>��m���m�<�ǭQd�,�"$��w���
�f�<ɗNG��e��eQ'7�&%��o�h�<�m�0y�&�\�y@X�i�*Sh�<�rE�9����٢AI���N�<�4BL�~���J���\�\�G��G�<qG�ҁA��fo��	�@LA2$�h�<iumH�o��ڶ+��QSȔ{���{�<� ��S��/x��� C�(��0"O>d �j�H]�g+�U҈@CC"Od-� g�d�"��&���&<*G�$D��A�I�v�� ��'�u��X��('D����B��AOV��E�v�)D�`���nu�`L�F���H�e=D�L`�%T�.Lٰ�

�)��t� �=D�p��@6i�q��ƨ,ؤp�A=D��kәy9����.�j�l��D0D�x�G=Y&�ip@�5�\{g�,D����I�!�FՂ��J�i-(Ö)D�,�U-[>�x��hɾD�
xywB'D�����C�F�;�� 6��K%D�@�th�\N(�dI�����1'1D��"5�\�[K8���*�2Pw����D/D��R��E�~AɁ�V�zh)�-D�$�P��	F�v�8��(�bs�*D��b +?�u�mN�*�U)�C(D�8�"6p ��!@��R�\�E3D����$ /(��P��@(,��,0D���1�V\��:��s�>x��a-D�p�6/��6ΤQ��K&�(���l)D��Ycˊ�{�(A��-o# X)��*D��G��#,���եΗf�L�')D���b�8w�ݹ���._���r�'D��"��x�>i��D��x@pGl"D��xAό7/rdb�A��[Zl�Q�' D���=| ʘ�$��`L`�,=D��-�t�R�W��6��:1�-D� �F.�f��kF
�>\�W�+D��h��^l)~%`��ǹO�lڰN*D��H&I�@��Q��=�L�bց%D�� �W�1�x�E��:"��I2&#D�,��XpV�R�cC\��\h&�"D����q�VDqς�G���yC� D�8y��R�N�v��#Q\��0e�;D��ֆ4Q^A0���z����Q@9D���Eh��(6d!���{��D��L$D��ҀԳ/0� �G���!�&?D�pe<�R$��B(�I!�f?D� �re�+��z4� �X����֢>D��:�kZ a]6يC���3��ʤ�:D�T�v˅KD�ԣwk�
4��;D� K ��0�}k���5WL�#�a9D�<��A�'}�	�Fm�4Hy�ā!G6D��"�̆�k�ZL��'��VZ��X��.D���ҍ<@"��j%I�X�a�7?D��Ѧ�|�ډbR�#`n�لE9D�ذ���X�H��S�J�LJ�<D������.������߭ 1����:D�H��eA�0�T�@���2(�
v 7D��2��� �蔹�n¦?N����3D�H�c*^?>2p ��@Tథ�!�'D�p��i\�i��M��%ROI�T��&D��aN_+`���Q�6���/D��Av�^�,wR���Ǆ�ְ]�J/D����%
W��<�p��=:�e�Fi,D�h�E�ח� �0h�������/?D�Ԁ!cˊe�`�0�::�m� =D�̠v錹iF�$c�Q���q�<D� �㬙0�T�'��d�TŊ��-D�hb��
�05�Ap�	H�^"zb.-D��q�@-'��@2��/3��J6D��c��J7����BBßJ��# �8D�� �Y(�ضA��!N�~D��[�"O�ĸ���D@v<C�ҦZ'��v"O���DO�+����"���.1��"O�]��,�8:M�`G�0����2"O00����wXH�!�]u�"O��"SôqZ��'��@���"Op�8S-Q8�1P�Ѣ�a@f"O(�I��/w^�����ߖ�NQ"O���d)I�\�������$�8t�"O�����|�	��n�c�<)k#"O�����3
���SDʑ3�P�"O
I���պ%������j��0J�"O:q����	��I��R�� ���"O��qw�F7V�e0%H>/Ih�e"O�M��ȓ�=B�S����C�PJ�"O�iу
���l�t�\��a��"O6��V��s:*tp \�;(H��"O`���C)���/�lv��"O4�X�)��5�� �O,^�;A"O�(�"�^�W�t�+p�.V�݈7"OF���P�8Rr��!���z"OD�Cv�D/5%�� ���,�#"O|�[!eP.-ڠ�vŒ11��de"O2�dj�Oq��r�C�{�@\k�"O2 q��� ���KU"�%��T�w"O���3n�:V���s�@0cP����"Ox���*�9H(0���`�Di�T"O��S���)G��X����U9Ƚ0�"OK2�������j.ͻ��S6�y�����CH�a4贸"��!�y�J֟m�\��GE\h.���b���y�g�`}�a�N�Ȕ�-R��y���$B.t�a`9 ��� Q��yR'͘H��#��B���!s�-Q4�y�gݡov	��k�.� ��� �ybC[�-�jd�cJ!����&W3�y�N�
s���RP�����Ǣ^��y�o-�F #ᄜ8W��7)���y2�\�]d,y�/X��x`J]��y�i�P?�9!���.X<�AfD��y�-��)��8��	S� T@#��L��y�!ԅ4�4x�%�o`��2�����y�E�G��Y��#���s��b��'Q�E���G�OW�<ˀA���F�C�' ����d��M���ٲ�J	�'��	�f 1�y@̜�h׾�[�'n�ڐf]1����	��5bV,3�'��ur��_!`��NI�d���'�4�(7�
�}"��xg� Ul��2�'����L�u9̡���4Q,���'����ֱZ�TI��G)BX�	�
�'vD\p�DX�&��%�2&E'?��i8
�'����F�
6\-c�̍�Wll 
�'Lp	�#�9x�ĥB��^<� ��
�'nEq����^���#�o��2��':zh��U=��y���8(�����'7F�r��X�X����F�=#�*x��'J�§<
���Uo�"'�f-��'��ɕM�<
 )M�T���:�'�"��N�$b���(�S8J	�'� jwK�s��D��)��[[hYp�'���c`�ڍ,�0�'��+O����'!��U���+�B$cgHW�S�R��'��T��/R����Ǖ��PZ��� \T�Ӿ~� ��ǌ
�:��"O���$�.e$��+*s��� &"O��r���1����G�^�@L�"O�<��H2���c�H�h�����"OJ]�ąڷI����C��	7U��a�"O œ��S�Jl��%/
�$���"O��"b+Y6vadU�.<i�Tif"O��׆�"h8��J�G���Hu"O����Θ��d0�V	Q�x%"ȡ "OxI����Fu:�� �~�@"O4���Aj�|�"���-H��ԁ"O8�'"�RA������Nh���2"O��	���>��i  �#f�D��"O���k'"'�ف���<\eZ$�A"O���Ɓɬu-���,����U"O8� ���"�2��"#ܵj��D��"O���5H��_H����"��82 ���"O�`��G>1L<1@[�k���e"O�����=J�$��c9
�%:�"Oz��ό'~��4!`�ו-�D�"A"O����@�8���@�bҔ�g"O�p�䔂Q���ρ_ΖQJ�"O�iP���A�j	8�C�(~hX�A"O<!@D۳5.�M�6d�;kV	bG"O�� ���`�a�\6�"O,��gU -�ܡK"O�1�*!��"Ol�;q���Y=@a�1�٥]����e"O��!�F�:SƩ��H��L���"OLp8E�U�7�ڜz��R�i��2�"O�]▉�0v�Ӆ&��\UD 4"O��DJ6!7�8{��7��k"OJ1���-r��	+�P�3ϰh�E"OޝH��R1q\N�*a�ɇ��Uڲ*OV�k�.ö�:� �lQ�d��'���0�#X(n�̴`P�I�z�޹[�'��|R����B0j��S�)�H��'�ܨS�[ KXn�a7�E-&�fĉ
�'e�Q��dr��e��:ܱ�	�'y��c�7 }4L�fkV:h��	�'0N�a��L�D��`A8`�k	�'�$�q����Y�@�)	�'ߒ�{U
=�ƕ��*��hڽ+�'C�yqQ�d�,�Ie��
�q�'l�1�i̯:xJuPd$J�� 
�'B8�ٲ�X�h��"�ÿGc��
�' ��b�+G4z�yq2�@�=k�p�'(� �#�$(4��1�ӞB�V��
�'x�Di bU%cQ�I0��>��I	�'T��QMA���s
X2���;	�'h�k�Ey��tH�$+�
� 	�'ߜ����@5pj�c$f�=pT��'�jmSgΛ8�&ѓ�X��J�p	�'�>�S�^v�ʓ���4�R���'-�S���d�BC)�3'���0�'���S���rвh��3�T�'Rv�c�ʕ~|�1Z8aV����'DN	ڣ�L�b��e��OP.�ơ�
�'���m��E0\�B@��#��8

�''�]�F.��9a1���	ID�	�'��y�Фǳ ���̬����	�' RA�"�F4~B�4RpᅗF\4��'�"\�bCP��v����
i�'#4�Q�����������N��ȓv7$�Q��ǰ;{@�)N5?(�̆�S�? ^��BB�<7�}��������A"Ox)���/��؈��Ԣcx^�B0"O%+��K�.�b�)Ff��Q�"O��5O�Vq0� ��E59 3"O�t�d�>.��R�.,'���6"O�@�F� |�]��#� E޽ʂ"Or"��C�qެ8%-W{�IA5"O�L�SjƖ^<8h�Ҧv���3"O�	��/��z�>ฅ�\Sjup'"O����J��W2Fxq��֪��5sb"O�l��g'���3KOZ�g"O�X@#W�K���P�SY=����"OΡK��];q�H������f"O�+������@Xw :i4��c"O�	6�S�eB���O�n�Us"O~�Y��	�"W ���O�#m�T��"O ��4�ά/q����Ζ�@k�Y�"O<2`-յ;u$�i��_�$n�T�c"O4�#%e�������@[�D'"OƀbGhW`���e+\x�qG"OV8����M�r�z#$[�=��Q(�"O.��G
�;��}���#K�`�"O���H]� Ң���w@"Y��"O�59&�S�r�X3
�32<T�"O%�֮�6i>�B�k�0	2��P�"O�qb�.��;�.���	�*^�qQ�"O2l� %EZY���=�� "O4�&熊}䆰2����hAS"OR9�u$�=�
<X��԰kѰm�#"O>)Y��^B:x!��H';¾�г"OD�Z�# �|�d�J1q���A�"Onc�΋'&\P�KAD�G:��y�"O��{e9b�1R�&VNBh "O2�!M�
�& ) -fmZ �B"O���S�3}�>K���"W����"O�(�Ƭ[��5RR��j�4[�"O$����åZz4�֫��liF�"O��B�9T��U�J�1��q�"O���%��bn@�5��/���Jb"OnEh�)��ZO�郧mŮ;��R�"OL��B^�߾�uc9T04Mӓ"O� S'J�,8lx"@��~%"( "O:3�B
��:w�yql��"O6Lh�_�g#�l{c��+S���"O|�E^  ��R� �e�Ι��"O���v)�c�t�jѬ��S��		E"O̵`�g�6d��kG
I78���"O��:b��l�� ��	˯y��Q"Oxl;���;*�F��q��/a�-Ѱ"O�l�����I��g�S���k�)WS�<��$����3c��'������Jg�<aËπP-�q��َ7�������f�<1ro�:�:U�!�I.���3"aTZ�<�0��=�zx��L_�r���{�<�!"� �a�g#�
P�d�T��t�<��@�<fN
���2��8���Z�<A�P�Y��Y~���AL�R�<	b�NE ���G�|�����R�<�c�k!��b� �"W1L�@�H�<�G��H����ÇVx,D���#�G�<�2�܋\|�)jcKO*>�-�fE@�<	��G�X�����[5z&���� Q�<�oY#�l9���׈W4p���\c�<����!^Jd ���ejЉ��`�[�<� ��ҡ���a0(p���%9ʩ g"Od�� %~���"��r_hȗ"O 9C
�%w� B�:PD�H��"O�Ļ1e�D��p�ᘻ'�""OX4�2��<.gB�3"5e�D0(q"O�ٛ�C^#H��z�鞸O�A�"Oy����p��8*�i��zTTY4"ODE�FDA�P_�tb��f%���"O�M3"���?�LX�l?>�-p"Oڹ�h��e�p��6b 4G�����"O��چ�F ��3p

1j�J���"O�Թ��Q&+B,� @AAo0�KP"O�<�Wn�a�\�TO��h���9�"O��S"a�-K����$M��l*�"O<���0u��Iy5��.�4ls�"Ot|��H.O�uc*܇B��8
F"O(xVʀ�e.0y�C����|�!"O�����jδ��b]<)����"O&Hthڱ����'�h�T�X�"O��C$F�PQ�=x�*�8"OZ�ia�؛@w�QgR5+�F���"O�9���!8ZlY�thK�I�`TBg"OzR�c"z�qAg����"O��q �Wr��eR�rt�X`"O=�t*٫A�XM��Ajtr�Iu"O��ĥ�7!X�7D��z^�\H "O��A'���-�@<S!#GI_���"O��H/I�,�6����V�3,Dm��"O�4�E-�CP�X7F��m �)@%"O�(0��K/J�Ή	&EI<=���"OXiQ !��z�t=񃎅�h�hlz"O�$(v�&���N�Z��Ai�"O�Ts�G�`sB8�4�V�!��E�"O���Ŕ��l}#dLܷ �"���"Oz�����M�zT�O7(��"O������2���:U�'���XW"O0�c�S���z�*��f����"OtRmq�@%����5s��ps�"ONi��V�LD)g��b��]
"Ox��aH��t��p)de4���j6"O�ef+Çm���C��Ax"d�"O��[�-����s��UgH`'"O���.̕W�
i���Ë��z"O� ��ˍ'gڐ(��A�/N)�"O�,R%�I�~�	�� �$����"O*�H2$a�=@"��?�$U�a"O�X���U0좠#��A�k*��5"O��:0BN�LH�䢒�M� 0�Q"O��h�TA��e@d�@�V��F"On���BE�<�,�qw�J�b�k"O�-!Ņ�&?v�ϑ^�irF"O u�a-0���I��ϴv���v"O4 b���Z�z�Q����l����"On�X�V�&"L���H]�`�0�"OJ��G1�|%�g�#u�� ��"OH����W! ~�c�f���q2�"O^`)��Ƥ�0	�@�9���	�"O�	"�Ʉ�^��	��$ɂ?b��H0"O4ju�U+ �s��lN��"O� �!E���0�u�ǀ*OF��P"Ot��JӃzF��At�ۉ0n���"O\]�a(D+h�̹��cK�m[D A�"O���'��8@�QD �v��i�5"O���sE�	�^U�"#Z����"O� �
�-�#C/�i���W�C����"O@��6�\����� �*�"Oz�Z5
Q	2Wx��W�H��,u�"OY"�"/�䌁��C7R��iB"O�� Ẕ�t�EH%��y#��W��[T�� h������4�y��� J�����b�R��s���y2态 �LMH��TU3j�H��+�y��8���〛������$��y�*�B��JQ�=%YrPb�����y�a�,���EF	r�x���H��yB����aB��8�Z-�J�5�yb��t����4N�=0P�`P4���y2C�8��0��P�"��dYS�_<�yb��7"�{�H�*�I�U-�?�y�*��0nX�RkɈ@�*�P`�N��y慶Q)@�A���&:�(���d���y�
�/����v�F1-M���R���yR�F�{�T�'��w�6�)����y�)M��B��P��!8�>X)&8�y�)�tW~�2�].��ԡ%h<�y�N�%2J.�sf��J5YJ�<9"�N�N4xuH�k��7�j�<At^�.��2�լ>���VF�p�<A�A�N��-� ��h�<��n�<��Ɯ4+z��&�E&F=���)�`�<��m��i��U;���߈l	��A\�<����+^*@�!C߶-Wx}�&J\Z�<	$�	N<��A��2=�(�0�X�<�Vh^���X��\�=u
���L�L�<���_�>g����Q�e�
��A�o�<���߫UR��BI�Ex�f�F�<Q�`�R%��`����Ap5�VC�<����<_�"�ր�L��	��B�<Yrͅ�M/���\ 
�nyZ$×g�<AG�(爠�� >B
�a
gJTZ�<��(M���|�'6'��!��+�U�<Q`o 6ؐ=��M����%���W�<Y�e��g�
T�E@.�"&h�]�<�1��"�΁8�'C�p��b�D�<I"$����V��:r]��2�cWC�<��`��n�@y�`R�vA̽
a��v�<Qdh�"R���aZ��Nq��E[s�<��DƢi:���AI["F��3+�e�<��'F�$b�b�O�%�شᣋW`�<� C,7rM�7 f��D�Y�<�fcD�cQ���#�*X&��b7LYm�<b�A���Q���%�6Ҥ�3D���S/nت��5ۺ*ul}B�C6D�x� !�~J *�j_��(A@6D���ը�3i46}��k�Ad��1�L3D�X�a�G�\ov�IX�zF���"3D�P��NA2/�P��iT)ܪ�H�)/D�\I۳P.Aqਇ�fQ��N.D�L�����J�"���!7l�*q�+D��� �M-���  Z�a6:�J�5D�P�m�H�0�ڵmV*a��H��4D��H%�ϸ7����+W�<��8�q�3D�k�$ZK��R�ӥ��Ⰻ.D�hrc�1T��E��E��)�&D��q �P!K�,�zE�V;l�ɉ�e:D��G̞?���af�S�8J��AQ�9D�ī��ؽ:'�|�r&��j���d7D��a�΂$�耫��&:�PՎ4D�� Ti7��;I�j%Ti����=��"OP�P3%
)�,�Eh�8T�~��"OD:�O����uG�aI�и�"Ov�XE�- <�]�sHEM����"OA@��Q�r�f%Q�ʎ.?�(�'"O�1�0aƜk����������F"O�ؒ�ǲE?0A��f� \B�"O���6Ã���0�W)H�l��1�C"O�9�E�W.Yba�N�;d"OJ�S���.0p5+/U�~P:�"O�����dI،�T/�"�x��"Ov��F��:��c�W�?��E F"OJ�R��
�^�pq[#g@�.Ԩ�"O"�Е�MTq�-�Q'�.A����F"O����W�F�H��f�I~:d�f"O�h�c��6D�����*�b���"O0�1��D>����z�IJ�"OXL��Y�!�����%��d]ܜ��"O��*$�&-;�`�Pd�+;M,m�"OT�H�Mқ�X���T(j��b�"O�䈅��h�u#��*`��8v"OVݚ�,��`Ch)��N��"O� �0h�h�V����`�"OڸJ��ּ)���(��d/$RA"O��@O�~%xT�LY�4.A!�"Oz8r�jծlV����T�7=be��"Ob��`�ʹrv��GO�>v�\��"O�)������1�h&P�8$@�"O&��a䎿A��#���<�˗"O2���{�ҁ��Z�}�T"O�hh �^3d������V\U��T"O��g�.�,���B5~J�ps"On1��L�z�CL� g��"O�%��B��Dh��_�/WP�#�"O��+$��y�D���YjI�JG"O������x.�y�E�&����"O*� ]/45�,�7ENi�8i�4"O��i&"׉_4��A�Ƽ0�"OĩӴE��(��`�̱RT�J"O� {U��*Xp�b0Bp	R]�v"O"y"�p3� �C��#�"O�X`u/@�=Ƒ� ʥ&05��"O@$��D�S�9*t�@;9�$R�*O�ܸ�&��U\��V���f�z���'vZɢ�d7d~1�A�ُY�(�P�'��K��
=��T�Uk�1KZ@=��' ��w�^2R���&GI,=�:9��'n��Wʙ	_�(�E@������'>�f)�fM�l!5GL��$�
�'��p���>'ڀ�%�v�La�
�'+VD����1��s�iƧ&��	�'l���_< z�8�TȠ���'<
���XJ��)�Đ��Ƚ��'j<1'�?�X�Aė�x�Z���'��P�)�<w��x�PZ�
\i�'������la�t�R
?~���'���-�Y� cw��E4(X�'ɖi�V� .7��r%�	E���'=��8d厈	��tb�$H�D7,���'�x���S�>���pt	ب@Qz\+�'��5��bJ�	����g���M��'l��Ȍ�G:���F�̀�$Dr�'{:!c� �!�Сv�
j��2�' `�q�#�'L��MӶ�G~��
��� xD��_9}qX���i	�ҝ�F"O���O�.�.%针�x ��f"O�a����0$\���	�-�4���"OR��
�?_���yߜ�""O|X{"!�b���c��Ej0! B"OZ�Zu��$T2hq�Ae�@��d�"OF��DB�~�N�VU�~��}Z�"O���]+Dz�hkW�Ү{�,Y 3"OL�G��7E֮�
V�Ċ�I27"O�i�d�F�J��2t#J:��XKb"O�� ���/z���C�1XG�YXR"O\��e-X7�� 2+ř52��:@"OX�ySa�WX�4l��4�zM�"O4�(�HW
*��D�A���qA�'� ���gB�(�:��I���ɀ�'����!�6t�*-��D ��Ժ�'w��J�f�)G�����N��c�'�n�1dmn�(����O%V4�C�'i&�j�OLEϼp�b�z��5��'�`���6�~�y �E�X|�'s�e�W�--��p�r,�&;����
�'�� ÌM������^�L�
	�'��C2�A9+ޭX� P,[��3�'^p�1L��8\aQR%�6$@ ���'
�32�=9�``p!o�*��c�k�<Q��4��RӊB��n1���g�<��G�iZ��y�΄L��U9㠂M�<�q&'J6��D�=v����"��q�<e�ĸh�L���[�qa.����k�<�V��
u�q��ƺD���Wk�<��!��X�����`��B�K�_z��ȓ7�๒�C՛p����Kňx'Z��ȓ?�T%23�,Iu����`Q���	�ȓ�<\!��U�t��k�5N�^���w�x���1& X��W����D˂�H1�U����1qo���ȓeZ�a���6��aS�Wx��	����Փ����PS��) -E6�|��H?4�᪑�Yaa���Z3�n��ȓ_�u�-�>��0���u���ȓm�VYF�^�1��0�/?�	��|<�hj&��H8L����Q}�v����yW�(C@�C�����c�<�`
�8�ChP�G\D�c�]�<iqc_"�Z���/�?Y����d�\�<1EKؗ���#Qŏ��N�	�W\�<�`E |�k�K
�^�z��2��Z�<	R@KM(jh��%�<�>�5�MT�<q���*,��P┦OEM���jXN�<��Õ�$���j�/f�@��3��N�<A�E�"��1	�:�,��Do�<qt�E5b�t1���Ă���I�g�<�0�L��*��G�jx���j�<��ވ�:h۷��{S:�:���e�<�B�̾T���	�G�/j�X��$X^�<�Sǚf�$���]�;��٨��IZ�<)��4s��,�W��A�PT��G�Y�<9�b�=M1��%�3^!�tJ��T�<)҉Y�My@�P�R�xd��ԁMN�<9�
[�V6r銷@V�7����'�C�<ɒ�

J�x���M# �`�#E�B�<�V٬5�4)���":Pr��d�u�<�!B�2B_nuJ'c�q��"��Nj�<a��(iΠQJ��4c�d� 'he�<� �z7�˳:���T)�7f)�H�"ODp��fҟ`C4|�!no���S"Oܔ��,mÚA��O��dӂ1�"OrU�`�Z�lZY�E�׍X��I��"O���(�H�X�3�mݣ;�`��5"O���E+��~�uRrꚷd��$�"Oj�p""O%4�(�8��H��v"O����X
I]#��͸Y�`p�"Oʐ�Q
�<3�$D�p��K0���"O�8+��5u:D�9�eoBBG"O6�St�)]t��r��ͯIdDd��"O��:Si
�� ��Ǩ�H�L�3"O,C��q��2���@�R"O)ٷjR�'��\SA� t �0"O�ɂ�/��*
���&�җn,ʸC�"Ov,*�*��^N,�4jD�#��Xt"OZ���ӃM�VP2 ��>%\	�'"O����؜*�����*kT��"O������d�N��"o�&S�䐓"Ou�6h�+_�lŹ�k��^��S"OK��,�-CGaY�*ID ��y���P6�ArbB�%Ҿ�i7����y2,V�p\�5�U�P��FL��y2İG��	XU+�`a$�塐�y"dV�%���3[����dm�	�y�ǀP���rg�5O^rE`��L5�yb�N�L��T��FϾ�j�]�y2��*5���@ș�E� �Qea�9�y�葩!*6���煔B8F��$�	�y�ܯ"RX�:F�S�F�8$nʑvr!��H:�����2\�V���_�5Y!�	t��BA��5p�ȣ��
�6!�H'E�:�Z��8u�f��"f�D!��+@�D��쌻1Z(��@DE!�D
Qߢ��!�Hx��P%5R�!���.u0�����C�Lhb<��#��!�>D��9rg�"�@=ڀ��'P�!�D\�8�jS�1~4� ���	�j!�D�=;���9th�#'�M#V�ܧ!�~�(�#� ?-h�ʑ�8!�U)��dS�"I�>����̈�w�!�DK8e�l�LR�,bL��nCZ�!�dXC�>�H�ؘ5�dQj��X,�!�D�.qq6�k F�>Ɉ}YL�>?�!��M�&L����*�/�� �ǋ��y�!�D�'@�J�,G�����4%X3T�!�d$��(��U.^����PcM�b$!��ȗJ�<Y�\�i�<X�E�֗E!���$c!�k�c�/������3!���q��K�/���g#_�!�Ċ=Eop)�0cI� n|h��X	�!��_7RRjdk�K*z���E�t|!�D�&���V��.K <���#�+ !�dip�)�B�7'��u�UB��!�$^��%Q�m��b�� "ly�T"O���u��M���c`C�?��I1"O����F����(H$|���"O�M��Em���90k ?�Vi�2"OJ5۷�1$ $k'��,Tl��"O�H���Y �T��(X{u�!3"O��he$� 8�܅jv�Aso�dS$"ON,ا���E�4=�`�|G�"O�� ď�t�J�����?6MiD"O�� ��Ȗ�Ps�G�q0F��"O� ��8E�^6)�N,C�㘋3*^U�D"O��T,��5��ł�LxUq�"O�Б���D�*�!��q�v)�U"O ���$e��ɗ�ә�Di�"O����"�50d�e^�*���"OИ�QkQ�PAp�AID�M�"O���%P�q�6�u��'�Vrb"O�s�/_�{?�f��z�)��"O�	x�!�F�����%�)}��8�r"O�]��Qc`�;N1e���)b"OҨ��L��{>��,�<h*%ô"O�Ő��>���{1���9S�Sr"O��I���}��8#g�*v;� Hu"O�y�Ǧ[�;*���R<y��'-̵��J�Q@h؉����P��@�'}���eݎ,�°/��:��)�'��SD,`3LK�Oب4Д0Z�'�)����yW�mJ�M=5Kb�@�'���r�P�/l��W	K�~)����'�JЀí��(��U�)��D� J�'�.�����%9ZX��'P�D�th	�'��x��߱��ѐ��m�d��'N���'ʌ:_6��	�����Z���'	^\��ۇl�,XI�GĈB
�'P,�0"��i���ϤH�
�'�BD4	N�@����Ŋ��P��	�'}*�Pf��$F�X(�s�V2v�0��	�'�DYc�HΫkը��$��m��\��'�Hأ��:����B��U= ��'�\���g��<��!ڱ�Z�T.����']�4c!�)���� _6����' v�J7�I������30B���'�"I����<0�|�2�ʖ0
��`�'*d��)��0�!  ]�(���'(P���]��A�A� y$���'��uK�C�0:>��*TGǳޑ
�'B��eM�ii0ࣄ��(���
�'�R�ʀ��`�|<��/^��P�'�1s�OZ'c�������]3�Lb�'Z`=:WDbnܡ�s'�)H,9�	�'�$%�.�0f��y�'�,�	�'"VA���]�>n�P��U�T�1�'��X�u��H�@#d)�j��'t��"�!I 	 A��BK�M�l`��'A�@�tS�Gy�]�v��=w��'�����	�'kp@�ߚi��@`�'2U�A�̄�h� Z�� pP
�'�V�0�K��9ćӎ:^��Q�'I�`r%�8%�A`Pg��|qB1k�'�>��&J�I�Ha�GCM�v�D��'�<i���[�2�*LC�@Tt�V��'m�h��LN�4�؅iw�������'~��m̨R��!0�C7x�P`�'C��av��4
\���k�֜��'>���u�W���`�Ȥm����'!�T�6rjy����8c�����'���	�*V�4�jt@�#��+��iJ�'�4ԋ`Ɯ)\r�U��;�F= �'_��@
�!]�D� V5聠
�'c��	���sj0��p�]�s.���'ȫ��$UΘPѥ�2y7���'2š���*t_��a�&�-lԪ��	�'�8*��J�u^-�!-��k�	�'�v�9�i��{�QCQDد_y4i���� �(tbA>�lh�4!��� �c2"O\�Y���"�(�[�b��R�x�"OB ���˦Gr��'��"6���"O� �D}� �B��X�O�|�R"O�h���	�.|�B�7jl���"OT4�2e��
,۠!E%n_�%�"O��Y��P%\�~��IbT� ��"Ou"�J�%~�dmhZ�L��%�g"O~�`�ƌ�+�\�3��W <� ,��"O\x�殜 �q��d��`(�	X0"O0����� x��Q�L�Y�|�3�"O`-��D�LH1�	��Q��æ"O(k1���!Au'߄RGX;r"O~���:�ҙ"�K]Z�6iq�"O.0I�@�?ptp;d
 3àI�"O�Ӈ�MT�4�[%���ڴ��"O�z4L�;|���	B�3Xt��"Ol����ӋG]���ejH�]���R@"O �:R,����P�H\,rd|AG"O�L[�ƾdQ���F"K&w?0]X"O��A�jK���3X�7'����"OtQ4�d�0�
6��{C>uI�"O���d��V��9Ip[�>7�$KA"O�1zW�)�UqqNɇ.~��a"O���E�'��z�J�EF���w"O.��`�϶^�|� �D�2�%"O��&)ۯ3��Ѧ#ff4!�"O��!�		h#,}@�(��DG"O(�Q�A
0J�)�eA҆b�J�05"O�IbG��Zz��t��0]m
h�"O���g�#no�%��oѿl��2"Oll���φ�� �nԫ)�=0s"O��kèQ,"8��ת��̰"O�����%T�@B�AӅ�b0 �"OD�Y�I�xdبw! �H���"O���0G�8�� �JIh��1"O̝:�P :�s�� F[P��"O����]�x�&�G ,x\yS�"O�)� �Ls��l�E�,	�Rh��"O8�  h�5^&�`�d�y���(�"O$�2��8� ��BI7	�\89$"O���O^88��a�GR��D�7"Oy�P	V"��J�OŦ$��%�3"O��A�3w-Q����^j���"Ojp�A�Y̚��ń_U���p"Ox\����VA.�(ƨR ���"O�]h����mYF��p�\`�$��&"Ob	���ըqC��2ш�;
9L�"O��@�� Y~8Q�f���X�"O�A��Х7���b���/�B�zT"Otِ�BN(hm���Ug1VP+�"O&�2�9��՛ue0^��P�"O��P�	$-��D[cE46���"O
M���	T;R��7d�E~��a"O���O[n���1ڑu>z5a�"O`j$�\+�l�`�Ȑp��1��"Of����d `b2H�'���""O�Ɋ!G[��>�!ǁY�r�P��%"O<�G�C�7YP�BFa��� �05"O*[�aE�Pۤ��0�	{#�bW"O�S-�t�����1&)ؕ�Q"O�@���:��� � �6& - �"O������
��h#%®PIj�"O�=3�'óPT��Q%Ɇ�J<s�"O� �\K���[���g��i$4�0"Ox��f&Z$O�҅#gf�bF��c�"O����J�K��iQ/�5�}ht"O �bB�P�H���N5wy��1�"O���(�"Ѡ��v���3gRL��"O���/�8!�x{d@
L���"O�p�r��� R��1q< "O�!��TW���!�&$5,��"O���;uz�@fV+3�QbT"O(0"kL���̛AK�<>
h�"O~��CI�Q���ۢl+��
�"O�ܣ����&��R�щB?4�Z�"O����Hls�Ю���"O�ẀM��
{��R!h�(��I�"Or'�MXS@�W�{"O�:vC�1+�t�*�Lrް�"O|���.	vف�A�:�T��"ONػ���4g����d�ē8&�a�"O��H�(�`z���Vر6"O���#&W@x��&�<|U)�"Ol]��C�$<�����%��|ҵ"O TY2JO)*
�H���_
h��|�w"O��*v`�$�b�	����S��iD"O`�� B�OLʲd�A��I��"O���D,H�6c����12�`��"O���V�˯	ZH�Ju�l��$"O�$3я�jQȈH��ǒG����v"Ol`�1	
`��ٱ�U�#ϰay�"OV�)A	2�yCeύ9��y�!"OF�{Wn�zPb����Q�K��"O\�x ]	*q��6�ӷH3@���"O\U"a��0�B���6A�$TCW"OX��R#�S�V�؁n˸�5`�"O.-`�Ϯɬy3g�6 ���a"O��X��"c���%`A�N���@�"Oօ4%�='cf$��(S2$�=�Q"O6��U�\��Į�/$��q"O���pl����䉠핋@ib"O�X%�����Am��.�����"O�sRh\�(�T��+��o��ȓm�����dm�՚�-ї%��ȓA��aA l�HP`��Pl��O�� ���̳D>��S�P�3DB���q	CזSA�e"F�� x>���n�"|*��h��0�V�ݛBO)�ȓ;\p�INS�p�+M� R|���02(��mK7;�O�Uw���?�a�'Lz�V6w�l[��߄�P��	�'���+dG��*�� B�&�ܥ��O�taBoD�7Uθ�Q#ݙ�n�2��'����x���BŤO�4h��:D��3e�]�vD�9`���p�.����7D��H����C�Lc���Fɩ��6D�L(���t$�!˄��#d�aO6lO��|����~݉�P(1�|���n7D��Y�.���+D��G�8C��¦���00Ѭ��f�L1+�N�2�N0D�\�'%F�t�ԥz�`�v� P�0D��;׬�3Y\n�91�T��ےA2<O#<��$Y�r�Z�
u-+\�� r�շ�hO?�*f��`�BZ�9N`�p�B,Uk��H�<%>y��>H�,(���6E��C��u2�)�ȓ4�P;�lU�bĚX&�Dlb���h0&�"���)
w2E�a��F�!��S�? ��U��f��Izg�	����"O�� �G�1��0kP�V�"O\0YGi*A�h��gJ�2�<q2��O��=E�D+�|d�
�%�L��$�����y��S2lD� �N!Ѽ�&���yBf�^P�@7��
�`��A��x�,��dQ�ީ8��@ZD��F�B�I ߂��AP�-��r!J��S ȇ�|��Ō�!���ZaX�W� ��=I������	�J<���(N(HX�,+�GZ �?9���S%C� �%T\���2W<z�DyB�ɢ�"�;K�����أ@5��ro����?�'��j��M�xO
���#B�* � �'�I}�Z�'`ࡪ��@�
����		��i��'O�7��/����C͘�L6	����AR�d��&���"~��K ,�%��.̾.�|!jS�
Q�'�?a �fD$�M[6�]�9���gD"�	f��$Swz��@4o�6�h0(��<�	ռ��'�Q>�@0H�b7�ap�
��Zu�IQE>�IJ��8c�ܐ��]�@�B�!=�ա��c�������
A8j���A��|Y+���0h�!�$� ���K�L�U�h��Əξ_����G&,&�ґő3(K��	�)܀�yRJ,A,� H�&�z(#��?�hO���.r�8PR��*���'�ME�	@y��'͐�Z�B��F�R �*c1��C���xrڟGp���`�._�����ڞ�yG�S'%��O�&<V<��ʋ<�y�i�p��xDɎ�.K�%�Dņ7�y�ԏx� x��#��3)�i��	�y�
�([�~iۀ�-@��f����y����G����*\�*��m�&��9��'��{R�ߚc�|�8�O�0Y�Tኟ�y�NX<u,�8���'%��`����yr"K5W8�0�R ,a�a̖�yb��$mm�B׆en5А���y2dJ���� ��ª	�d`a��ǨO�"��+ǟy��Ke,Q�,�;�\~B\��%�"|��d����b��ɺA��C��L�'kax�OX��܊u٘sq����<�y���� S|P̝�!�@$�W�1҈Of�zP�]��تnn �C���d�<IC`G'p�x=�U# ���D�x�'da�&�-5�>1 ���!<@T����2�yB�G |���!`ĲX���[⊉"�?��Ǡ>�M<E��Bߑ;b�t,��u�P��v䘄d��D{���'O���
�04FЌ�i��'0\$�ش�Px�+�.C�n��%픣F>����)��7ў���P�$x�����O�)8�C�I�4g*�p���zd�$S�ګG}��	<ў"}�2eB%��)��a���!`l\�<g ԭ)VH���b^qdd�QI�W�<!B�4o� �"O�o����`�PT�<� � 4�^����J9"�ř�FS�<!���-R�~���K�DM�Y��^Q��:�O,ճQ�ł9��8�4N8�Z�"OR�c� ^'����_9��c'"O<E�p Π]֜8�alʬ�|��"OZ�ؓ&G�_���H�?���"O���'n��'e��y���/2�9�"O"�fFSEО���1��m�W����	�R�}��o �>���b�FP-��B䉗e��	a5b�m־�� ΍�t�C�,0�`�V��'C~�"����~C�)� �u��N+hį���\�B�����O
��ۯj􀠤���`ѱ#�N.Q�!�dC)@��q7�-,��H�c.԰@������o�l�O�H����Ŵh�x� ��_f�8���'��E�6�'�R���I_�	t��H>9���)�� �1A�M��O�*��~�R��Ȓ/��F�T�Uσ�&9�M�2e%D��J��1p!��b&O'w^�E�(6�	E}R�S�VVr((����X� �q�[��2C�	�I�:�Q@	�Kl�����ŭ?RC��:W&�X�`�ˀ$�N,��Мy�C䉭4V��2ퟞ{�lT�4�l���'�a}��[�,��x��2&�ތB0�ˑ��>�R�>є�,xo�iP��%[�4�t`�m��k���O֝r�ԎW�<	8Ӂ���4(��$��ȟ�k���ة�� ��Q[cX��E{��I3e�p�5G��o�^����;<��d=�S�O=^)���M�NS�����D�j>~U�M>���!lO^��e$�PD�,��)�S��h�E�'c^1l�g#J��d`^��N�iŮ�7~�xB�I�q=~�[P�]�Lt�y�Gӛ�T�>1�cw�O��A#�΂W�e�F��-E��h�'��hh�A��rMTy[��X�"b�Ȱ&?D�t�U	��f�0i*R��+�T a�0�O$˓\�J�� G�Ь�0n�\х� ]�1k���>�T�Un�&t��Ex��'9�?=�DmG��>JE,�U�A��+�O��sB;'J�9[4�JG�7dZ,ь��s�l�%�Ϣ.jʈ[s�˛�f��@�%��ȟ��V&�(Қ\��W'�!�CQ�D��I���kD�P�_�@<(�@�c��I��HO駹�Pʨ���4	�`�H�
!H�C�	4~(��^$s� <��!Kv�C�I7V=���S��;��`
�"O^��Q�
'~d�d���R�0%"O��C�R�V�8��Ho�qE"On�8a��lS�Ȋ�mT�fm�d�Q"OTţဈ�+�lUʠ��&��
�"Ot� �i�:E�U҂LT���p"OH г�5-��Ҋ��$��[�"O�H�w�ڭ��d�i�hB�"O�m�q㙒3/8<�3i�$��SQX�,��|���(O`P��i�����'�fR���W�'�B�Op�ؖ!�;p�6U0C�U>�����-LO(I��kI+:p�b#f	A
O�t�$�!6ԪU!V'�	Ӯ�3c���y��U	2���` �R>ȹ�J]���d-��u�����V�P��;��ɹ"�îM!�$/Bټ�R0J�b%x;W,ޚ��'�J�Ȏ��)��Q�����2x������[�!�d���`��3L��r�x�P���&`�!�׾$�� 9	W�e�>I��ȇ�&P!��0b¶Xi��b���3��I�^C!��aj@	�	�- �:x�e]��!�	1}C�@���
 >�|IH���!�����MD�E�"�4���j��/�!��U*I�!g� �b��	�Ts!�D�X�v�	�Yv��pc�B1a!�C�+��Z1mYx�JC3P!��̙X��`��B�R;qc  R�"�!�f��z'!�([���؄�!T�!򤄲`@A�`��#��:��{~!��V�sn�꠆<{ѢT�Cˈ�:t!��@��Kd���Ɲ���T<!�� rH��-Y#4[�jV! ���r�"Oz�S�ϑu�x�kaLZ�*ܘ�a"O6���˞|~�\� N@�p��(x"O�Mzqa��h5��iV��D�0{v"O!���$'����,U�c]��2�"O(� ��?�2���6 ��p"O*@�cP0wO�!��;.y�eq"OL�$�.|
n��ȨG ��"O�@ɶ˙����S�c>XY*f"O��q�m�4W�P	'b��M#f`� "O�L�Iգt����K Ufa�D"O� b���x�"%�#�V3N���"O��K�21��h�d/H @b��"O�y���R��jD�#�\I���"O��t�ٗs���+P�oC
-�4"OP�է
9-t�t�!��+Y�B�ӑ"O^�"�(ݹodaCJ� ���s�"OH�����-A��I�i�	�Tp�B"O$�� DJ	}<Z�#gݚݘ	�"O���b�DE`��hS=%gV� 0"O�1��şj8U�R�_G��U2�	� j~@��&�'d�%kaO	�J� ����)&`��'��ԣ�*A�{��%� �B�&�4Й�'t��õ ����X������Q�'4�(8��U�\ ����H���'"�5��O=Dj]�w�ݱp�x��'\�ԁs��QiZ�H��(i�"���'L<��lE�5U��N,d��) �'��l��k^8|-( �SmI-A<���'v�)�c��-d0P��q��}��'��zBd�=b@d4�-BxB��'I��ضe��T�pp`�G��s�����'�d=�及CmlI7+�	o�Ik�'��!���m8�-�f�,A
�'3v|��BTd5�efL+Cff��'����V�O��R��m���'�╀�;:<q��2j��c�'��d�
�N�|��)îI�D��'�V�K�cN�/(&9���C"���'A욱.*P*���Y�0n�ա
�'2`=��l�7*����	g^}{
�'��$X4n��1�5�C�Ъ�#E��y�O�-[�6�ȧ`�2G`TS&�յ�yRdJ�0�(�UD\�/�|8�m��y�c۔m�Y�4虿!�d�#W�S2�yB`ړ"��UA��oL�<"'CĢ�y�o��&�<��9.6��kVg���y򄁆|�,���4#��E!b�؊�yb˃�Ma�9zc��7]���!�$�y���	���z7h��xm@�����yr)��a�,t��X�p
�q��&���y��4�y�n r�6��֠�y"�Õ ��hiC�n�l��G��y���\��u�D���t �݁'�ċ�y���v`2X5� u�R�sDj��y�p�`(EB��1L���ĩ�,��O�	�A��S&b?�p�\�2�\�WH��Gn���%D�t�e.,1�@��
L��(ca���`PD�Є�>E�4+��;#��� Z�_R6����yҨ�u Vh"H\��&��BO�����s�l�����SZd��ē�Gr���D-ײ(Z��@1�K�;��})˞?�(�)�T�E������d)U�1=�PMy�O���B�A�� �E%�H� �%�	$<�P��7�Q (�dY�|� ��xP�q�uFB�8n�KB̓h�<� ��Z1/A�=ߊ�����9 ����p�'���3M��L�+pX�"~��O�Tߖ=�@m�v�^� �	%�y��ްVd�c5KƶZ�r��M���ĕ��r)3�H��4�
���#Z֙�6ӄ	�>�sg��%tay"-��~yle���e*�`B�Y��Hy	�@^;���!RH<)g�̅����nT�oH93g��_�\��$�RF��?熉��A�>Sȅ���T��p�bp�@É�xN�`ȯ��ă& �)E+3LO.m�R�!_��(Ԏ��@e��DR+|�E�@����79K1����hԶ;N$y�r�
QI�͎�T���S��:u/����Yhy�.��%w�-04M��\�up7���~XI�4��A#�KT������@�(O�[(O8�'&-F`C	�6&rH���d����I�H��QQ��z�Wa�\a����8���	��N�-�X8z5I"#�ۣʝ���)��<�'LȨ�+�ώ f:l�֮.?�*ǝ�\�t�=}��)��o�r�Q�OYjQ�Q�@�'n���y��H���y ���DH��u�P���g�
4��c9M��L�@�	t<�b>PV�Fr3��A�)ذS*�����V����2nĠ.jP�	�b:�|p�Z�:�q�a	@�5q�Q��]1��QYhO<�����5&f��b�2�?�̴�&�	4�\s2œ9o�����4V�)F�ؒ��	;ubLu{w���PY Q�R00X��CgT�rݎ�Z�$����Ov@qs#@�V�@���!��a����@EB��F���>E�D'�I��9j!��1C9D��#��>�~��
J9��Q�]play­��}ٶ%��0��#DL~�>E�O,hH��H9�1���
O0w�e�D�A�F������ C�:d����'\��A��F���C���.u`p���#�K����`�Z�6���Z�{r�ܛg�v���Z߫M:Z���q�-�R��P�t�L�K�l;��O��Q㓀�_�eۡȉ/�!���/Y!*}x%�U�Z�8����jS!��Sj B͊$eͽe�~Y��"�]S!�	�SD$)q啔�&�#�]V!�d
�g�d�1��+6�m)���!N!�D�+�:�S�	G��`M�R	I; !�$ �2� ��fעE��"#F�V!�d0)=�x��%���� ��3�Q���#qM�A�(ɪ'�@-�O�4`'Ȉ�{|��y���D�0��'�d8�v�T�j=ڔz���!��Ĳ�'vHu��M�F^�,9"+H-Z��?Yb��
� ��2m��z�J�
.�O��1k���ybN�E�*=0�LݜZ� X"�		�<��qyԏ҃c��Ց�� ���H�+�Q��
R�����8�)�g�(`�-l`���E$@�����X9�kI�`����)F��)�䈮���c/�5�$�R�*.�O��E� �r^)+㤍5&��}�ֈ�Z� \8q��r���_��-ఢ��fo���f��N��]�i�(}� �[0
L�ѐ,� ��B�ɏC�$EJq%��h�� Tk�7D�6�	$U�����@�^A#���B� Uz�e�m��0L?A�e1q�H5�f����slTk��@��6�R��E�iS�Lq&��c�<��$�D��U�eM�dW~�0`�K�C
Ax4kڷ��剎g(���sf{��d� �K
�
�|aV��D@9��x���0���
�xm<l�ayfa�o�<V)���L�Lu���+F㐠���_�T���#I����Z�����YM�$`��ܓ70l�S��:~(}�C¼�e37�� )V�9�4����p�<�e�9!�"�P�
_H+���J���;���"���T��s̨���#�2� 
�J)�O�$���R�/��X��(H82���	�)�����?�6�8EP�̪nB;4���@O2.݄�C�O�ɰ��4t�Y�N?�h�Ѝ�;�ư'hG	J��C <rz ��B!�)��O�\��Q�$)��7	ƾ�i'�D�
¡ Q؟�wK�
f�~}� �ֳ��h��\�q���p&�7�i�C��.L��j�>��W�%���ʦ��W�ZиѢ���y�E�X����A�ZLCt�sT��$�����.���2ǈ4��*_���K=w��$��(��;�TC䉪+&�l�4��;x(�<3�A��~➜c�`X�u>axrKE:xl,}�&Z>s�:aY4'O��y��'(�b��b��s�@�ʳ.��y�G�H	�4�b'F�p B�S��yb�M�/-dxZ��� �\�iᦈ��yrMi��oں|�zH*EΎ�y�öt��цK��CF�L�y
� ���.L��T��`S,Z�|"O�`�LI�cq"�zդV7VM����"OV�#A�]����bԢ��Uc�"O��,� �Dd��`	�	��ر "Ot ���WP
h|�V��dVܙ�"O�E�u�Im�H�2r�WE��]{P"O�"�嚫�D��uŚ�I��"OJ���M8Q�*�Ҥ�";�"O��z���(Q� ��G9k�Z9��`�/Q���=E�ܴt�����1d�Ԡ���@M҄��6�R�x�.[�.�j}����*���y����*����$�nb�#�.��xM�ؑ�lS��a{�	�:q�}�⛌3�@����x9g��!���WIEDh<�J��4	�X��D���8P�G�K�f��aÁV�&�i������Otl���^+rm���!�^-�<b�'���qD��?l���	t�ۖ^��+�hJD�"��6j��B4��d���(��	2V��T�$
\Ǯ���OY�XlrC�I|��ᕀ*w$��u�oZ��з̑]8�2�X*S�D�-�p<q'e�3e��$�\�)Z�kw����X%�٢���*5��iE��`B8H"�M=Z��m��[W�����àm��،W�r�Jc�ߊ^�'�v�bh�T~�!�,ۤ/��h����n�:KӲSa�4��9z3!��"I*�hx� �;�]Z��7x'�⎅4dAC[�w��h��	0?�媔9r���b���uO��h' svdH�vC�.T֤�H��t�1a���7k:,����̈M�p��D� (�M���T�������6E��y��T:��͚6�5B��8�NK�e���wa��h�N��D$а 砸svOj��A� e��qB(3aL�,�|H�cK�J#�R=0f-ަ�1��E$D�4j-�H��_$X!�$r�"O�9¨��X�||:@�/=)
5��"ޓ&�r��e�F�
����P�H(�P�mrpk�-܅3Є�!.��R�Ɠnr��K$���y;����:y�֤����G�j��PtQj�����*�0<)�]� �j�4Oŷ������x����B[�LT��$m]�$� �O[�"���1Ũ���a����[����|��=�wE�/~�V��M8i
1OT鳡픹j,��'(\yS��������K��J��ϱM�d@��OZ��yr�V��v�
2�M8����K%C`��ьW�#���È�O�X��Y�(Rg!�/`Ū�[�e�S��a(>D����®f4 `��0��3���<&�J�C�t\�s�+A�ð<�� ��w�t�#J���[�h�h�'QBy`0P�Dhd)�x�]1��io�lz��jO ik㷌l��� �T��d�@���A"ib�\٧��\&q(T���I;�@�0� 3�:��ﬨ�E��0X�0�Ŭ �~�|�"O��ȷ�XN~�cVk��y�v�d�i�t��"Hw�h)�O��a��&>7��v141��W�^���%+�;A�|�T.g�
q�T�vсrG�����_/sT��'�  @/K2��5��	 樈rE�8X�ba�VD��d��<!0��"ᮒO�H���"�e��_1P��D?r��xP�9ݐx�/�"n��A�ܷA喡A�F��֔�������H"��8�ȓ�g$��FR�%�@� ̬�ؒ`��Py��$p��u��i�9=�6��B۟D*�(��j����>��6�>%�|�t�E�.0ԃ2"��o���8��ܰ�y��Jp�Tu�N\=fD�8B'Q��F�r��p�H�Ű<��Z'�((aG���\Bѡ"nx� ��"����mW�+*2�G�Ǻzf�f��7r�!�ɤ(b>�"R�K�B� �Ə�3�ў�zb�JL��@2��	��W�b�0b��h�µc!��>�!�;txs�N��p�ڹ�P�?��$�1E�|+g�=��Ӕ%��M�&�ܣ%��5���	��C��p}z%"��0T(���WRV�'�i�p��E���QD]&Ie�yɀM_2��h D��[���}�����2D��#>D�$cr� ��2��Z 
a�08�k=D�\���S?8��͕�h�srk;D�� E�e��!� �d�1M����1"O�����m���b�
�I��%"Ot�) �OT'6�y�5���"O�X���D�&� D�����XB"O耍��?qH�T!����e"O.�#�O �@�G��4)�A�w"O̜c�Q�ն����5{	�'�8�z�Ô+?@�C3�\sK�L:�'�y�i��^@|qC	�wRU��'����0�*��w� u^̱�'�lٰqÃ�$���
|��'�x�!E���Q� ��&����>�y�
�K���!�A/+0i��E�y"��iQm���U�Sf��u�H0�y� Ww�\ˢNR:^��U����yr��K�˔�J#-��2j��yr)[� !�4)���6�0"�Џ�yҠ�8���[��Ԅ꼁z"�S��y�l�8k�2�H���_&���L�7�y�d�0avj!�_)|+D��n̬�y"g�� �8 *��\!��H!#*Ԗ�y��O?J��d9 o$�"E��� �y2';|��i��'��l�2�֩�y��[�X� S��T���ց�yBh$��0��	Q�y}X�p�M��y��Q\@+�a v�.d��f��y�WP@@s��c]*a�5�[��yB^1]�����F�=P����F��y�+)�Y��/ٽHv�i��f��yB��0�����ؤ��<�)���y�̍��8�� 	�0ūp�D�yML��l∫�24CIA�y�M�2*�d��.f�H!���y,	�j��it�	!nM3�@��y��Đo��1���%�x�Pl�y2�X,P��-`�	�'��0�	��y��-+r5�d�Y�-ˎ��$ ��y"�4pڰ��ǫ���ك-D��yR��RV"	:2��&
�e��OX��yR\B-f�"C�J�zXM��%��y��%E�D�@�����	�(˳[;!��[
kV�p�-Z�_����7H�?�Py�Ř�Jc�`S88ߐ�X孒�y""��$Xd��:;n�0i��yb�\-"�9���>����l��y��:и����&(	��j%���y��YO��#��#,�"�#GE���y��33[� A�,�(�k��y��\��ŋa����q�iI	�y2a�'�D�c��"Ir9�K ��y�l� ���s�a��#����� � �y"�V0QĄ�@��f����*�y�F�y��Q2��WtjQ���y�NWD�Ѕ0؊�·�L��y�$�0������(����Mݺ�y��Z
��8"���$�u�1�[��yB`�K殉�g�ر1�)N�y�K�?G.�����X) P��%o��y�P(PIxL�Re�x2�i����y���8,G�HT�G�i��F����O���Rd�Egxb?��ϗ,�\K&��0�n�e�+D�t�Q��n!���֕VwtA*�`g�/O����#k�+��)�'B�&L��y�B@�+=G
I�ȓpB��+��S��Ե1� �"Y�6ŗ'�Jc�&�S�h����� ���k���5��EYf���Bp�'���Р�E����WC�(�IХ�A�]Q�`[!B!�䃇E} �H���0W=���1a�G�ў�Ӑ!PN1
�El�O̧b�V�"mЎ~H��#��|�(��V+\S*˲`@e����J�4��I�w��s��U�y*������AClI��VU���A(s��i�0�6D�ᱮeI҄� ���y�lw�剢 �f��f��H�ن�I6 _�\�e� P�Dň�\�����=A�X��4gZ|�r4MI;R&���ϻL� 8p7c�P1�����9�x���_�����g�¨��J��I�4��y#��(6-�dÅ��^��TI��\fI��	�):NB��;T�ɂ7�ɦ	�<��a������$�n�X����;�*�Icc^�9O�H��NVW�0=�cm�71�c>-�c-Қ54ॣ��jI
}
V"ٞx$�IŒP8Մ��hOY25�L-u`�-����M#ZX��'V���r'�i^8P�)ċ KҴʛZ���K�U�(�Oy����DsI8$�7�N�~��q��?%İ+��=jsn�'[�r`NNM���:��M/\��a��� ��l�Tڬ ���S��?�B,�*��e����1?$tt!6n�X~r��frVظ2�\h���uÞ�co	�<��iS_>_�t��zL��t͚�����	�X~p����^6�j�pf�.E `]�ŗ>!�,Z7[���|"���6^���ЋΏC�h��������F�.)�2���'�T��n&�n�9���8 ����HL�X�1�LFZ�	�6�܁�����1���~j���[6z���*�p�{�K]�Ԛ�K��*�IY��>�D�S(���cG4i����͘O�0�Q�=<|$Y��X�"~�	�\��Y��K���iv���4�u�s�M&ҧ��^� �c�m2 4�(�~�EH�<�q��!@�x�ay����RX ���ca��8��Wm�>�O��{�.�1���b�^������"Sw������$z;� ���Q/?*�)���Su���e��j�~u�ѣ�?F>�:1cپZ�HA��{�,߭h�$Y���"��u���D/32�<IM�{\��$ω_d`<qJ>Y5��v�����@M�E�d�A��e�<�`%�[�R����<肜�ćf�<Qe���4�,}�A��4p6�y���h�<��G�+^z�𴧜�o�BDiE'@d�<���*,�Ɓ����u@�����c�<Y�����a��±yVi�4�d�<1E�E���bC�|N	�f�y�<�F� 8\u+!͂%c�֬rN�p�'a ����(P"V*�j���[�M���2��&5b)�t���yz��R�UX,@���G\B�8� Q3E�T�D�R������xXaQ��[�(�����ł��'�V,j4KR�<A�o�6��Xx��� el2��GӒW�j$yC�ͅf�&j��C -z81��(O��i� �ep�@f�*�X];��I�j�ds�AN�	?T���h$y�-?�f���%57�ZȠ�@��r�"���'�8��e)�+�Z�i2Ca��0.Ì\��Й��5}R�܆�4u����3A~x�B���'��Y�Ƞg�]%'Ml�UEN#A�!���r��%��T�wDH#���	X�j��qaU�tK�R����z�ЅL�\ɤ�&�{�g�-m���S�'���4�Y�o#|O�����#�8�k�4 �^��L��t.y�`�:6��bb�M����1���7�[-�h���$�=O0l������b��y�L�	.��O�]a��}�n��I<�����,����!L4%��B�fh�u�I�.�KbD�3M,a}��ߦ�j���iE���0t�8#��E ,WK�R�'E��`��0�"��� �E���G4Qbmۄc͈��V��?}�.4h�"ON�7���\!֝cV%+-�����'�b��傜:g_���bHK�Y�L��X+µ#6��k�S�^���څ��$P�Z0�tjN�?������N�������:�M����t��*��I��iࠢPL���PXYr������'�"��l-V�ꤨB"Pvv����N.[��Q��9���}�X��
ֆ�v=� ��'5�a@�&:�puP�'��	B��:-��o-I� ̛�� u�D���{Zw�֕�1à&z�i�O��� EDЁy��-���J/D�{AfQ�-��*�p���q>?)U���E�I>E�d#���sƇ�%�����f̣�y"��p��ްmJ���c�ɀt�qODġ�$�:�0<�W>0V�kF���� �W�<��)S� �X�&�P�.`��CI�<� ��2D�Y�01�$��G�-H;�ѹ�"ObXzPϑ�"�U���^�''93 "O6��#��c�~��TmE�da�`� "O��x'�/..��H�I�(Q���"O\1�[�f����*Ͷm\X�'"O8�vM�2�����\N�ih"Oݛ%�ڡ;����{����s"O8��Bɖ<@�>x��fY
B!��J"O��`.̰F&�c���Ց�"OT�8��L�02,pbƌ�x_����"OL�����k�\	psLYG�
��"O�V�8m%�%�5�ݗP�\��"�V�<���]�=�z��ЌJd{ pC6�C^�<1c"L;&c2�k3�Y�@ђ�T�<i���x.|���\�D�؅�0��R�<�d��+�
p����vǜhzע
B�<��lA?�j0K#��<��dR�.[y�<)�-�)�$��OT�������L|�<�r���O��5kΜ=!+�� c{�<�����JW�]�M?����U�{�<!�*b��C7�9-|�òK�q�<q�@� 8�Ap��AuqL��m�	tsH���'�@h �����tä�̄J��	��;��@ՔC@���pK�q�N��u��-'\E1�'����!�V�S�b��7�X@�4���d��Tfy�����O�ԀK�lR�o�ʜ��g߰@q��P	�'x^���Űؘ�@,0��|h�'Eh&�G�bj��O�>)�f  �jAޥ)*M�y�b9��H4D��I�w#��Q#��+�F5��� }���2[B�:t�A��I�&�k�����g0�}��<�O�l'�ԙ�z��ǺI�UC�c\=xXIa�
��xr���v`��J$~~Qw���O��P�FX�R���Q���MMJ�ԑH��<���`7Ӗ�yrJH�2���	�:\|(�&���~�<DEL����Qt��+vT0C5,��NS�4S'n0
�B䉇�nH�P���=l썢F�X2$8��'z��+5mL�gMt���I.�h�'��vu�5�u��\z���d�^+d�@wOV�n�Dmu�F,en	���&v�fC�IGx�m��(D� �h�&
�%䤣?!�-��? b?���J�:2\�xQDKe��#�9D���׊W$h8�b�#=b(��*D�Py��F�n�� ,S�j�p�x4g$D��k)o0Ձ�WR~t�B)D� �u��:Z|H(��Œ�+Z����5D��j0gG�o(vm�e	d�ZB0D����B%?�@�����_�H�(��-�1�*\�.$§����HY�6]~��AC�	K�)��*CZV�Մy�f09�MB�&o�e�PY�7���S�O�z��w�͝a�Nh�qi��,M*1c
�'�&�J���$��zQΏ5����)O ����<�r�C
�g�|�� �!/�b@����d�Е��	f��� �F*I�*UH�,�R�#��}C.���%ΐxҫ��ge��q��_0�=��	��hOx�R�kX6q��1����Z5b������A����x�mV��y�鍭w58Xo��%�	�diB��?ic�#�~ � B9}���g<6I��E��3��i���Ӭf<B�ɊMe�E� �ef���ӨQ�c��ʓ;��&&�!E ���$��S���v�W �N�%d��|[�}��xQF {5�A�h�N�EY�f9� �����ēa80Miw�P<Z�1�T3��<F{�(XOTԁD�V�Dܞ�0B&{rPM"#H)t�$���R`��"#�������5&:�̓&��4rOO��S�OB�2$�)�&��B�\"�T	�'4R�*ýJ��qaÃ'$w���H����Ƈ;OIaz
� �xk`��g~����5$>l1"O���c����D�����t"Op��J<���dcM�����"Ol�Cb'�x��%!�$n:ucD"O�	Q�Y��8�KI�!�6"O�p#U�0Zx���ׁ�y����G"O ����#�r���B�OG��G"O�a�L3R伕�#'��#����"O\�ԍS2���*5��p��"Oʔ�`��D%4lE�T��#"O���c��.��["Kq�|��"Op���FG2 �Đ'*N'/�>���"OQ@�i��`1�@F�`�r�"O�ZD%Rx�P�P>d��"O�@'�۔+�FQ	`��3:|=B�"O��H��ƃR�T�E�R�+t!�"O4��w�����\�d�Xi�W"O�=�)ن$,�8�D0h#�}��"O&h���vmZa"�:�:ձ�"Ob�1v��[̤��E6<0� Ѳ"O��
��:L��a��!��?GTI+5"O&y�F�Q�j�NT8E��&V��A�"O�%�c<�H�i$�?I ��"O,�jb���m�$�\�{(f�#"Od�#����N<�v�}��ȓ�"O\�Y�M�g��d!����~x�"OXy�5G�6S���8DH]!~��"O\̚$�8C:������"���"Ob(c��p�I`�-뎙���5>��z�P�lQg윰^��mZ/w>��m��2�6���H��X�ƥ{DǓ� ���GK���$��:����ԟ ֝�ScJ�p�.� 3�<(*��<�㞐��}��	:���$qF��w����ABX�9R�ZG�DE��ħ/�0���G��D�1c�U�
j��%��ʋ��ɗ_^��#��#l�P�%B/E���i,�̅�I�m��,)�\��mc�l�e�<B�I�q�R<c��h��d��nC�]�H���4и'�j�x�l�q�"����p�ƌ'�de�?E�$�	l8FP�ʃ�긄����|�B�ɖCDEܓ�?E���u�U>T:<���.�%6$���B��\pQ�,�Y�X���ɥO�`�T�DWe��"�M6�dM,�}"ӍR�|fj%#ЋLp傶����(O���6����j��X�2l��&�@�4��dQҠ�'�j�XW�P����A�%� S�N��'2�ܞ�������!(�~v��V,Co�J���O ��w�����)�<ͧۄ9a�?�0�2�*������m�s�����O~��a�(U�jl� �H�71)��H��d�O��@��)��iD�"L�䡴�E���Ƣ�C�D��%�@E�t�J(�-`Tq��,�je��O�Ġ��)§ꊍT�,��C	\'I����(A���<��S<s]��2f.�Q��c�@S!Wɞ�;ǅ/�	�WȜ��i�:v��e�+����&�M�;f1O���6�;ga���_\��y2kM�E����ǧ��D�(��M;4�xb�)�'hS����9V���h�_�?= �lw��*׊U7�����G Ѥ��Y�(���ُ&�5��C0IWp3��&D����%YT^���������h&D��@�LO�Պ�҅e�KP��#*D�t�a����%�Ĥ��#�T�<D���B��b!��D;����O=D�xIF�NL��8&E�Tj~ 04J0D��Qb!�����lĺ��P�$"D����i�(t�B�%+�0�P0H!D�X�2`Ŋ&�2���o̱GͶmB%%#D������b��=��!_�)҄-���?D�ds�%ޖ+;�d�d��p$Fa��M)D�� �l����}s(�!M�)�����"OxaR6A'�8��U!X:vyR���"O�5�(ڜ4�R��V2*k�U��"O�D���Z)p*0'�6$pe"O�p�0O�':U��!B�#r���"O��+�Z!g�R�!�J��HA"O^�#�� .Uvi���,��s�"O�pI����~��Ӷ�Q�P���R"O�d�D'��~���a_�P���"�"Oౡ�Ѵ��m���@/Iߴ4�3"Op�e�7/��x�Н?c��:G"Oz�{� T>�R͹Q�>O�@B�"O�ѩ�*����<�W�	2�u��"O�$��,5|����P��"O�K����&��
LF�+ �t��"O�t����a0�5qrk_�B�d�Kc"O\�r�??�8$��Ē�[<�y�"OT�)sCH�BI`�I���34�m�V"Om!��T�M89S�b��T"�	d"O@�y����,�6�D!�t���"O^9�m��_�J��e �U�z�t"O��˕��"cc�0���P3~:Bpy5"O��y%@G��Y�K�'8��r'"O�� �h�9=tD%`�	_ Dp�"O��
E���\�\dy��G�p҅"O1@��d��1jߗ|`�9l�(�y2�ʅ=yX��a�&C�,��C��/�y��XI���s4MJ�I�v�b����y������貈�*�Za�gÃ)�y�"B���0��\zj���yRM"|�AC��Z�JE�%֓�y��Y�7n�1�IA\?���`Ĉ�yB�͐69b�d�O�&��N�1�y2%��&6�X�&��F��4�A��%�yb߱Fͦ�W��,��t��#K��ybF�M8���C�P�dݒf�!�yrcU*o�|ؕT/0���cG���y�⏤tD̨pV��XI�Q �yR˚�4��!�h�L;:��e`X�y��#A�.8B�U�E,�)]C��茌s�6;/ڔӃJ^_ULC�I�*���ڕd�.!'���6�$�C�I57����Q�%98�$�ʸ��B�	�/��e@#s}��k��H�WTB䉹T�P�&��2J���W�q�B�ɖN�H$R�ᓘ\"�|X¤�)8>B��@�(���I�"��R䎅�B��1/;h�����q@0St�&��C�ɋ&?�QC���5 �H1�P�YlzB�7C�I���WbJM8���C�I�h���8w��_zu���+g8B䉦9ǔe)�^5�f�@�)_B�	'b���+B�;:_�%���>Wo4B�I�I��S�L���K����b�B�	20�p�铏q��0����:��B�I� �,�{�n���&!�ƃ Y*�B�Gc�t��X*L64再0�nB�	�%~������S��y��(�EۘB䉧;ӊ)�JI%+�*��U�nB� �r8:�jR�����E@�^B�	�(i|�S���z��i��6h�DB�	2q��Ѩ5C�JP=�圉:m(B�	�X����f�8X��A4�
|��C�;�N)�s�C�y �3Q�6�:B�)� -Q��
,(h`�h��*����"O��󄋇x.)"p(M�zE�|�"Ov�xr�H-=�J� &�/U�\*�"O��F #8D�q�FH����R"OV�K�N�w*�(F%7y����"O�3S�X�o���)�$^�Fnœ�"O(Y���A@.��9��181���"Oޥ�4+�%�*�9g(M�$�jq"O!Ӳ�
H�Ĩ!���xI�Y��"O )Zv��>p�$c$g5n6�x�"O\�j�e�<S:�Y�c�
2�ey�"O����j��.<��$"r�,�y�G
	odV� F�R�P&@��/�C�	��؁eȜ�P��&�V#L)�B�	�G	0q+\�<�>ȁ�-U�nF�C�	�Ff��J")�1�:�šȝfC�	a��h�`��n q6���jB�	���!��D�0fB/c�JB䉲T��e�E�@3>ha%�ٜpClB��"H �sjژDdxr��	�<B�ɐ )��TB�C�"u� ��>	&B��1�\e��#��_2"�@�mX� �FC��?C��4"v�_�ڼr0ke�fB��6C����L(^���'��.oC�	*N�ڢ�J�v��+�)p/.B�Im�D���h�;Z(�m�l�Z�C�	�\��
�E�*<,IF�Z�d�C�ɰi	f�d�ѣ^b���e��^C��R�Vq�b�03����U�u��B�#Nˠ,���4��-C7.��a��B�	�<@�a�ȕ-eӞ%P �X�xM�C�I�/W�0��/\�F���t8�B�I	3��h��]�D���TNB�I���K�F�2=��@dP0� C䉋�F����אQt�h�0B䉕9�"D)��D�bGh�B@��!d~�B䉜jb�܊0��+4L�����(P�B�I:1�\��_�4��{"&+�^B�7�H����U<J`t��P�Ց�C�I�Dh�� �d�8U�T�pj�B䉭M�@�VK��`4#��E��B�	�Q�2�!f�.�*��g�4j�vB�I�x~�d�'��Jn��Q1���r�nB�Ig6���W�2���(� ��3�pC�	�&�(T2�Ƌ|�N��A��)�B䉵`n\2D��Y_ҡkaG4:*C�$y=�ugF!�`		6M����C�I�t["�@�� �
������C�ɏ:vL��ԩ4M��ZR`K;5ZB�I>AZ^-��)���ia���6B�ɯq� ɠn�$���"D�)<�C�0 �Q�уہEJl#��&qJ�C�I9d��xx`�J��Q�X�rC��	`hE2�˛f`�����#h0$B䉮)n�9�ML0<)���N(\�6C�	{F��˘�B�䘘����e�$C�Ʌ2x�\b�Mg(���P'�;BC�	�>�X��W�˴
���C����4�C�	)+,�m!�g�%_X�͠���z�C�ɏh�D�C�:c�­S���!��C�(oq�QI�va�A�$�d�C�ɔ[-x�$�lN|dK��m��C�ɛ\XLS�T4k{X( "��>�VC�I��j�@��0M:��҂ٲk��C�)� ><��A�Z�>����W)E�vhc"O�lg�<fZ�Up1o")��p"O�j��12�0�S+D�]�S"O��eB�.��,��@�q�R'"Oƌ��瘅w:V�0p���(�Z"O�D���sO��c5�I�X��"O�3rL�#!�h,X(_�y��k�"Ov����U��1�e H-m�Z5W"O��tl�^���̟8�p���"O=±o� >n�J�Ǐ`��5��"O�8���_���i�����|��v"O.<ap�0�8���S�
���[�"O|%cQ璓�D�!e��Y��(�"O�m�TC�*E��3C��9��y�"O0PD&��� ���w���� "O"�Y�b�=gpz�yB�N��� �"O ����H=p�a���tU�B"Od9W�X�	��9@�Ō��rѢ`"Or���9�8<���
O����"Op�SŢ�Jp(p�F�_�T����"O��Ke�"M	ޅ���(�VH��"OL�S�T�GƸ �/�V�"O�)zRnUW
�X��;��=H"O� ���� E���K��]�p�@�"OH����:wj(�e�/?A�a"O0����
�Rx��B��V.��"Ol�m�>�0�ʢ��.���c"O�<�A���}C�iro�8+����"O�5�e�
Z�r��֋Mk�"Oj����	�������-���"OJU9�Ҕv�,�JJ#YM,��$"O�Q�mG&JȤ�ר�/ր�iq"O"	��,J��XV�0�\��"O�1Y��T"����
��taB"O��r�W>+�͡A�@l�[F"O�P8��[e�0Z�ɡw5��G"O�M�t%�wy����n� *�3�"OF�+ %	�v�F`gM�  iH#g"Ox(�Q��2���!�IǺxZ��i"O�p�� 8�Y����8a|�P"OlEؖ�L�M�4�c2���!��jV"O���5k�!�A0��/���v"O�%Ċ	r��$����'���g"O��AY"#�M2D�|Ȳh��"O|\�&��<y������H�#�Z�@�"O�ɑ�F�k���
�XEaS"O��w�ގ)�0㤡\�
�dl�"O\������/Z�y�F�E2&�dٹ�"OP�Ϩ?\����	Z
��sB"O>��T���r T�e�i�w"OX�h�d��8�֔��	�<˲"O��x�j�?\,�y��ſz�P��"O�d�5��~��"a�F?�6Y"C"ON���h�Yit�(Ge�.&Iҵ"O*��LT
lB1B�#^�x���G"O��Q`�v8u���ˣq�|���"O�}�7hG�]�b27��Z�j}C�"O"��,@+{c($s��� @���  "Oܱ��   ��     r  �  O  �)  4  7<  ZF  �L  �R  nY  �_  �e  4l  vr  �x  �~  A�  ��  Ǒ  �  N�  ��  Ӫ  �  v�  ɽ  !�  ��  ��  ��  ��  ,�  n�  r�  ��  � p	  Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�� |d��"O
`�(�;���8���-0��1%"Oj4��ND^[��"3/9�0|H�"OB���H��*�ʞRy=a"O�味V�!X��!&F�:J�$���"O,��a
���C�Ą�M�"O,$3%o�-���p���+Ն�:1"O��ݢ1����`���y14]2��i�<�6��{_���c�H�`�fX�$Kn�<��A̼VI�xR[�)�Ć�pඤ�ȓA5��('nߡ4�� �)˩%� ���,��r�؊b#`T�eT09���ȓ!�b��g��}�8�F��-? �ȓ
K|m�ș�VṔ���2�%�ȓ"R�X�j�4JN�1�˘X�i����̹	_�jZ��1!g��zܶ��ȓgil,*�J�
j�Ne��i�J%b���f	�(U��:���G��$Y^م�~r�� S�%T"���k\�jx�ȓ|4�1�îJb��@ӵ�ݩn�V��/[`�"�v4�R�!ʎ<��M�ȓ`:��z�ؚh�J�Z��$HY:	��H��p�m�C1��!��B:��0��EnjZA V;9����J[
2���	��4'J�EA�IVW&��~�(aZ��ӹ�>� o�Y�|�ȓ�f�A�
Ο7�H��M�$�����mޠP����/���ANXo*�ȓTv�����{ ��-7�*h��I��sB�8�8���3����ȓNe*M�悡;������X�o��!�ȓ'lj�#F�m�+R&;�|��2)n�C��0S4���T:
b���:�0!��e֊��)��ͷV��,�ȓ0�&�8#���� ع�L�����;�P�AFd���,w�6d��r�EQ�( �gVlɦ�M,H��,DP���|�I	$G#\���ȓ"�)���E�B	yt&B�^�LɅ���?��6Y�[�K	� H𑌊Y�<��)QeV�xJ�&=M:0�(���X8��Dz�!Q.]�0�kPg�j�j��;�y�C֡ #����*�e
Z��W�X��y��27�� ڇVG�	�ʩ�y��r��Ј!�|[�Qɷ�ۍZў"~�i���CiZ#6̹�E�M|Bpąȓ<+�<�4"KH��0���I���n��<��/"�͑?DS~i����5}sZ��鉚)�qO�P�+.�iHW��.���e"Oީc�늴*�Yp#�4,���J"O������lx��[!n��aq�"O��C�d��Y���N���� "O	i�A�Nw� b��&f0���"OxiY!GO&Q��\��!c]�4��"O��;�f޽l��<� ��l�P��7"O&A�î��(��%��n�C���w6O>�ZX�@JF��\'��W��<(�̜8�=\OlOf�X�;�պ��O�f�Pƥ	#���>O����וA;��:P���|4*����$�S�'X�0X�@ R.rjZ�2�J
Nt6E�ȓy���c������CpD��Z|�I��`��RHr{�{!��8�mE|��3� ���6urp0�.��_h"Ol$I5�UM��1(өW�AX�$ �S��I�d�@icv��Xx��Xd�_����4+@��nO�p�!��7~�*�<�`�.OΌC�N�6-�l:6�ΚG��)
��'�ўl�Vj��n֑�2g�,UM�ib�F'D�l˥BM}8.0y$�8;����,$��\��ħw%<5KV��6'��=��.�6��ȓG`�,x�H���L�3�\�,�ȓ�J	I5i7��=�S�Q>jw.��0�LА���<�,���P�w�Y*��$�Ic���Y��h�c1vW�ic��<w�}����~�L;P�j\r2��(I�xE+W�:�Ms���s�*�"wW�4��!��7Q�LE��c��AZHXSF�O!����ɘ-�y��B�F���{��TOh9y��M��y���;q�uڐ�V 4p�e�ǻ�yR��?W,�eP�DS�	��i��y����TS`��m�"^�Sp��ybB��� �0�ۘ1�4�$���yJG�s��5�Qc٘,oFE{��Y%�y��R�!\���$�*<����yBkҊ6�T�1��L���)cF��y��	=)Wh�7�I�A��HQUm���yB�D4&}����HN=�N0	%K2�y�Sg��� �j�F	(�j���yD��[Bt���.Ԙ(nΘXD�R��y�&��	�AP&m��&��(��K���y2�,2�N|�bh�/�t��G���yB�md��+`^�}���qB��yb��$���a�4E詊�!���y�K �T���L
����P����yBǀ0<������(Tڠ�\��yr*�`� 䡢��#2�#`���yҌB�"���Un�B ��$��y���&pL��$!,n=���ytC��(v,��94�3�y�dޤ;f�����ȹoJDk�?�y"	�t;��
&��FаV/��y� X���`�@߷	�x]Ia��+�y&�%�*�ʡ
W(} 舃D<�yrƙ 
�y 6�� q�nd�a��y�dY�+�<Q�GN'lj�!hf��7�yBiO1 Ėyɳe ]�i�"���y)�9/v��3$�M�ԡ���yr� 6by^0���E���1���yb)X�/�p ����Yv�[!�];�y��Q#H�jR�<%�Ѩ�V�y�)߈v4�ǧ˖;�N��� �y�M�#
�t+oE�GRD���T��y�A��mɞ� �E�@�;�ʟ�yB�Z0����d�4Od�y�勜��yR�h:\`aS`X+uG�-RE�D��y"��-)�"LH��ȊfE|�b�.�0�y��*Hg~@�+[q*MQf��)�yD������$�b$ˆ�'�*!�ȓ��-����@c�%��W>e@���x�{�kS�xk` {/7[�"��{>����E �Y0g(H�}#Z��ȓnW��éT�`HsY�~(Q�ȓaDv5�3LL8�H B����ȹ�ȓ;ޠ�B�䎊�����&)Ku�ȓ+��[#l܃W	��u�7:r ��j��8��%�a_��C���6zǐȆ�S�? &���V(u��,�7A�I���""Ob�BeE�
s!����%�ʐ+2"O��G���<��qg��0>h��"OZ�Z��),�L 8�@� L"�+�"O�t*�Ȝ0���&�εL_�m��"O\U�I�2,����K�jKuh"O ,a�&
}ZM�65�Ih�"OT�����PFb	Za.�.FXb"O�;5��h�8��KQ��"O̰�N�	x*��Ӫ�C�`�*b"O ���h�Q��<`�J�?jĄmz�"O`��Ț'`���r���2�2�"O���"'M .| �jC�@$)�`"OL0���L|B2W�I�>CJ!�""Op呄�s�IsE�X[T9`�"ON���t���qF��F=����"O$ES��N1)%`��Q߭r׊X9W"O�d�2L�sA��f'X���8�"OH!�.^a�q�� �w�j��A"O�"�����aK�+!H���JH��y��Vl``t��(ըH�G�B�y�$��5����}M��۞�yR�}�"[���5��8�#�H�y"����(��A���J�ÏW��yr`S�����+Ї���c����ybn��yL�#�B�:xc����A���y��p��J3��n��e�']��y��������J�<;���Zw��3�y�
ґ_�-��n��"B�@p�Ӄ�y��M�_B(Tb������Bi\��y��� *b>Pc���M"d:�yҠ�"JKfUzƊ��2ī�^9�y��'s0����8�(�[�CJ��y �7^�8���n;&TB��IZ��y��T�za[�U�U
XĚ�'N��yB�B�PD�aF=b`]R��8�y�iǲl��n��s@�s���#�!�Պb�l��"�zݰ�G[��̆ȓG�H������'�M)x��`"OL����nLdr�bM�8B�"O�����ָC�A�cӐ�c�"O8z�ELoOr԰3��$��]ɠ"O*yh�HΊ��r�$[��x��1"OJ(+�Ȅ�)P��B׉�3����"O��3�����t����8\��b�"O���
Z�EQ(�B(ˡR،�"O��YR̒Z;"�� ߓA5����'B���gZ�Ђ��|�԰�'���Z�ڎ:j���(�[�L���'�HM�a�b��' �Z��	�'��;!� ��v(��^d|9�'(�a[g�'A��	S����_f�4�
�'���I� ��]�b�2V>$�c
�'�H*1%&��IťO�!
�'4L�G��<ocRx��GOzrH�
�'6X�y��O�8� i�9x�ll1�'��r��d8�5��AS!g*�1I�'�6�h�/D�'xȹ�D�49�9x�'�uP�=娕)vL"-���'�@���|6n)�KK�5����'̖��pM�>�,IS�k�����'1"�BWYF����R�j�a	�'	����[�w�\�!�(r&���'Ζ�8�J�37"$@� ǖ�qiz����� �a2�X�(�̳�''ކ�+"O�$���ծ#�z+3�,aż��v"O������+1����R9|��Q��"O<RC�_'�����P� �"O�]p�hIGʠ��ݛ|���z�'���'e��'R��'R�'�r�'�J��sB@�*'d ��J��@��'�'�r�'"�'tR�'���'\��ե#l�qÂ�N+ĚA{��'��'�B�'f��'kr�'�B�'�8�p���dǊ�Ҥ/Y�v@��'B�'���'���'���'���'��H�7%�H�DlIξY�b�'�b�'���'��'eB�'���'�:%��ϖ�:����FC� whv����'���'-2�'�B�'��'<2�'�E+� Tv��c12Z(z��&�'4��'���'��'@R�'"��':��mƔL4���Fh\�$�jp�C�'���'���'���'""�'���'��ՙ��P!w���$�ɊWNB<�S�'D��'Y��'�'�B�'D��'J�*5D�?4��8��ز(Q�S��'\��'%B�'��'���'["�'R��KAˋz#�ua�c�e��I��'���'"�'���'��'��'� �j���!�h���ȿ �X����'B2�'%��')r�'���'�B�'L��q&�8n=TqD�A�$�$�y1�']�'O��'D��'���aӶ�D�O>Q���D�;&T��b���~|*Ney"�'��)�3?�V�i�=��@F+��i�P狘�
irb������Ц��?��<	��iq��Xn��JO����c�J�hko����
�6"?�H�����Ѧ?�4����BFj��iͩǘ'k�Y�(G�� ��4[�}pvHŉF����AEL�6m�5M�1O�?y������LC�kh�
u�:�@h��I˛vAa�h�e}��m@?���2OZ铣�)3��h��@�.
U�i�?O�2VJ�[u��*R�=��|b��p 	I�o�P��d��X8����>�Ĝ�x��:扔:�wU�#�j����	9tS�O�H�'�v6MBȦ����R]��(hF
g*�Iw��t;�I�nJ�Ô
�34�xb>a�4
����'�j�s/���.ݱs'1K�d�_�ȗ'��9O�D	�O�RC1�匲Ofڐ�7OJ�o�#c��kL�F�4�2��6=M��hi�IzD��4O0�o���M��'�Q �4��dVF�d���F��+�J,M+�Th�ZSߺ$ ��#HF�'7��21�e�g��� ��k��u7<�Bt�\�)�C�I��a����<x�ՊGjEgy�8��P�����W�r�nt�VF��R嚀�5k�u��h@sQ�����
fZA bhUE,r��7�@� [�QI�!�%0��=r�6��r��>�!��m^it"(ö�E�4s���"">��m�/T=Z�
(���G�S5^UP����!R�"���|6-�O���O���JO~�I��,F8a� /�6w?��x�J#�M����?15���?AL>�'���C����%J8)��X2��.D7M�"MImZϟ�I��X�Ӟ���?���U5}Ԗu	�,ڃLĠ9"�9j��HR�ҙ|��	�O�QۣD��@y�`��1]]Z�	F���I�|�I$x!P�L<���?!�'&�YJ&+�s�ش�Pm�J��ݚ�O���O`؛˴<����?���~/��c~z�2��T8�)���<�Mk��d�ܨ�.O���Oiʟ��ɱA�^�(���ur	8C��?T���'n*�`������O��$�O~�$�Ot;�ˑ�0�Z�:'�;or�ًj�|�8���OT��?aL>����?�v:n���C�,֦����_�YԐ�!�F~��'���'���'Q��'"<�*n�&gH(��o</����"`��˓�?�M>I��?qJ�k��hn��iSx����u���s��'27�듺?I��?���?��g��?1���?��[;`��x"���� A��ͦg���'4�'��'���!�F����41q6m˰gB�H�� �,nZ���	Xy2�1`r�����1I���N����aa��#7��W�ݟ���	xU�"<�O�xi�@���/���S,h��ڴ�?��*
]*���?���?����?!��K�H`�S����K����Z6$�86m�O8��χ"@�0q����������J3H�=q��T�g)���y���'+��'D���'��R>��u���b�`L��C��v��E��Ś�M�V ��<E�$�'�E04�����'��R���b.}Ӟ�$�O��MT����OJ˧�?!�'7r1鲠Q�7�4իt��t0����(�IN|O|J��?A��&]�9�#�°7p}��7#�8���iu�h�O��D�OP�OkL��iQ�	 B�R1Q $�ћ�'hބ��X�$��˟��iy��'�R�[(�uz�����
�~\`(����2��ܟT�����<�*O�@z�B<��`#o��R�PP�Tc��6�����4�	]yB�7Ml�S�nc��
�	&r8�҅�1�b��?����?�/OZ�d�O����W?=J��T;R�\l �A�>�|D�gH�>��'rh-�eĔ�zf��g�ID� ҀU�V\`Q�O���@�E�0�4���L�m���'�MQV���Zs�uy%�T��r��'*܂SK�z��T�T�%y��`�f�(2و�J�O F�����;d�)�J��1[6�zb�;��Ģf�'ZǬ)y��M�]]QY oB1PzX��6M��3�ͩ$����ƃ#'��� �Á�"$���x��A;5xlR�`��4��$�P?��d� ���	t���`瞹�V51J�O���OL|Ҕ��R��4 �˅x]P��F�y��*4*:鰀�G��ȟʧ���?���H�&�j���6H`I��{^ ��ϴ�`��D�<޴��BD�v,��O��w��0���yU�H���+��-�G��S���lӌ��
���'��)83��bI�IB�@7'(2�s�'4��'_�=JV��%C����j����1����c�'����'�>Q�ph�*�Q�Sm����
�'��lZ*�ȉ��'�r�'��Mg�I�I���Y����D���G˅�H��H�/�B}��Y���-�P�Q�"�p�g�'G��R2�@<u���CM��	�BE��5� 9r=�x��S��ɾ5��E�TN�)�I�T�^�ɐ/:�����=AM<9���?9+O�$ɉsP��#��^$jz�ir"OD��4u��tB��"����`�K���ɫ<���� Л�"�d���!޺n@R�j�/@�*��'l�'D�0�'��0��|�OΑ"�D	�b��VJ�44Z��U���	����D�4i�n5Af�/=�H� $��eX�irD�����xåü.,�󤊟���c���	"�eJ'NS=�l�2"O��aHy7�`{�l�n�:�"O6����Bn�U�ӭ��Z��)��7O�=�>!���|���'��_>a*�k^�)K�H�� ?T�L:ĩ
�(����	֟��� `�r ����kT�B&���?�O��,�&Z71�`J6�Q�{l.� ����ؔA�V?f��=�< �jP�ÂL#z�� i�#�59Q�l{��O,UG�D����fN����"�yb��r����eN�ś�'�*�0>��x�@\.(����A�\N��a��&�y�lǫ]�6��O��$�|���-�?���?�W��f�BP[q�S/p��5��![u�.�He�	�"�z�+�m^x*�Tb>��D�O����?����4N�+iJ����+g.����V�x�<(���*���q��B#@����M�}a�ʞ4�>8�I�S��?�����H;��Þ��k ��|�< �߭"B�@4@ԗ��4���R�'~�"=�O�^%s ��!#���H�6)�\x�D�'9�L�)}� �R�'�"�'��-f�e�i�:b��Do>��%�r?8��D:�?Y@N�n"����H�7I&�3ړo��u��:}���4螧l�����lR�+��FW�M�J��el�c�4��	���3w�;?i�*E)�2�xS\�{sT#�?�W���?A�i7j7ݟ���h�'�D1���B�b��"3[�|�'����%p[갑p�jdH0�o"ғ�(�y���A<i�����"ȉ4���f�c���	�*��C�'���'O$L</"�'��	ϣ?$��'=����UF��9E�O)}#d����,�'��غ�����Z��$���v��p�9r��Iџ�p��:B�}����}�ٕ�:D�|!V���<o����������J�<13��lY���|�>Ɇ�C�<��i��'#�����}Ӣ���O��'k�F�ٖM�4z����Ō�j!�4�3	ߚ�?���?!�f��1)݄^��Iq�d ֯zi�p��g�#nf(������(O,�Qd�[�jԢ����W((У �Lu��]�ƄÒ#N�\_t�3,@3^>ƣ<��c�ݟ��ڴV����'��ӆ�T� �Q}��3G@�]�aN�D�Ӻ3��9O��5@��Q�0��(�w�l���'�D6���	)#Β�V��)W��<��O� �f�	�J@x�zUlNџ���c��@�'?DR�'�B����;ԡԵ�Nq[4J��$�Nź��'1O�3!����g*J�L���P#��'-�(BUM�|�ȕHW�<Y�)��h�A���tP�$O^�Y�ơ������I ��S��?yPb�,i�M��,�1 ~%��QE�<�F_�`$a�f��#��:���D�'�"=�'�?Y��Ys
i��V�+��b�o��?��K��07�?	��?1�-����O�NTM�P���/@I�"�E���M	+�~�#�F�k��L�B	�6M���i�xL�PsP��4ZOp�R!��*�,���Į<�j�3�4��Q��C���	!>)�������1�=!�(�.����W�E� ��Ĝ~�<��*�5I��)��Y!n�D���뒒S����d�5�lk�4�����(\V@�ive?��Ԩ���?y���?Ѵ��?������$��p�phϒ/�L�s*�q��'��;58�i��T*�l��ԂA��%���cOS�B�F��''���&D{r,����)P�k� JRh��r�	�і�d��=*$��	�%67�X��e�׸�y��O<f!����+q��A��Р�y�Z<+X�2���O�ҜI����yBmz�ؒO4�t���������π ������)�� �%s<�4 a.�&���O��d�&��DaRLE=�
��N����Oo�D�uIt��\��I.��m+���/B6�路Z�A� GB$�
��{��/��ic1/��X�Q�����O���m���tX��.X|ȕ3�S'Ah�xQ��Ɵ��?E��'� $�V`��6�T�hS�e���'��6�F�M���d�J�!c� ���ᓠ�\�"�Ɇr�!	�4�?	����	^~{��$�O��Ʉ*Dt�+�gK�8`8�3Si^�u�������|�U>#<�" LN�����g�*�,rcɑ�)PHy�Ɓo�<�ph;����'�Ũf�3�b���=0tȱ�܌j2�'#���?	F��������G����	�b�~�Γ�?Iϓ��I�j%�`� �]_� �ܜ�J#<a$�i�7�1��?��A˖\�(�7��=�����ʟ �I�[���0��$��Ο��	$�u��'R�9Hl��(Qc��`��Ŭ�y���ε@���0=��a�>yj��[��K#�+C?Y��ӪP& �[�_���$F�!��LK�K��U��0��˵Tj�$O4t�$�$	Φ!��t�'Q�^���,N,|
tz�I!�@u(D+�xy���ߴ�?��O�A� )�' N��j�`�=#0҅�4K��nv���?��kyB�ػ�"7�G�LA��!��TX"��bA~���Of�D�Ozh�Ą�On�dz>Eb�$�ul�Ё�BA+x�^Ա�a��Gm����P�|�MK�q#���S�R��M�,�)�2�'L�`��}�ԉT_���"��O�qn���м�%��}=N����x��C�	��
��Ї6VF�9ק?Z�C��_��KT�E�slи8�^�=_�	�M�O>S�Bw�f�'"T>!�c�Ң%���%#�XE�L�uk=2�Iʟ��ɀyؚ-����j@$����l,4�ٮ�y�jF.4���r��U8�e�*f�Дi��H3��h�0'0�	�O���`GIC7p�X0����2#� ����D��K��'c��l��D�O�.yc_~\�@I	H$p����?����9O
`q�h�]�܌#B��DH@�ٱ�'��OL��͏6P����`߁up�7O���j�p��d�Oʧ;]t���?1�) ش��PN!���u�`Y���!G9�D�}G���&m"1�7]>u�|�	�>G��Z���2��aʷ߉p�\PӁ��u|j�c N�F;99�%�������> �蔅D-�I�M�>�J��I ��S��?ѷlۀm��x'�[�4z�t��K�<����\��je�A.e�Բq�C��?I��i>���DR�t��KI?��y�V$�3���	� z�$��VX9�	ޟ��	�X�^w��wL�ʲ�4��Y�mԁN�x\��'b��$���3nY'8��� e��=4��m�R��Q��	9�v(��J<2Jr`b����I�"W���<|OH`��	�d����gI�4�"O���-Au �:��\A�B��T/�f���>ف�K٦Y���r��0�cI�%�*��	����IП��� ��P��۟��	qBE�3��)��T��n�50X�葫ơ[!�E+� ��6���
)�j���D7ʓF:��J�b��<��*E�G���e�Y!]��Z�`�;϶�h�kP n#1� 0	�	!�M /�p�Z��v�]1�j���~ћF�'���,�'��&�:��H� �M��g�|�C"O~�d�%,vt�
%Vx�(�p6Op��@QƦU�'ʞ�3m��Iܟ��O�b�/�]����5�1f�8�u��x���'�b�D8iC��T>)3� o��SC¨^�X��'6�m��D�dk5n}���FF,�мҎ^�(O��%�'�"}*Pʆ�7�(���HM;o<�@SJg�<)3 e�����l�h�{� f���I<�+iC`gL����D�N�<����	rw�6�'�RV>A0 ��h��ȟ`1�)B�k+@#�
��\�⍲�!���ĺ��!$����S��?�O�1���,:��Rɵu���)T�37� ���ė;�H�JthI�q��Z����H �!*E)�����R�A�.%>*!y�M�,Mx�B��!L�ĐR�)��0ь��vT��) �4C����� D��h��9��)@J��Ji`xk�I>����Ο<9����<3إ��e/C��Фߟ��"Ж!�w�O���h�	��u���yW��4��e2rʊ$������im��(��Y$ì01�$�4-�R̐�O��<	�3]�x�ᣀ�>�v���E��dZډ.�hl�@֚��,�sĒ@B7e�LصA����9yƜ+�)@~>��aϋ$Z��\ M��'�>���(#b�6�8gGE�}��i�'����`��=O��fD*�T(��n$��|bH>yT��ݛ�.�5����O�'Y�f�v�F��'��'�&�4�'�=��L��i��r2� <HD/�Ip�I��F�|��ʴ'��D�^х�8K�"��!ڍ}����A�&	�� �VJJ+08���lí)k��ۓ��[�@X�2�U�qO"H��'Kl7��v���3ȗe�H��c#'2�!�$%h�L�S�,	�%������A�!�D��i��8��>_"��єE�0#m�$���9'��Pq"T��MS��?�,��%��b��R�qU����<Y(�
&.���O���RYC�B	4〕�fQƟ�'lw�93W�/�=��ҹRv<Gy��	�Y�2�N�4%���F��e}�N�p�RP`V�K�lKT#C�;��B�K_FqO����'������'��#��U	7��� C��lKJ�;��'��O?�I?5�+0�G�.&^Y*���y�T��$�f�Iq��i��I�*6�hK;9\:扝��`�ش�?�����\;�����O���U�t�����a��2h��Д||�1��O$�O~�g�'s� #���C���S&\ O85@0gA(D�8���F� ��Ç�^�6S`�R����ֵ#i� Ii�yB�fS�sl�ɉ�n�;3�$���O�������'&V�1�L�
z`��zbN.x��d��'��|bR���?1�DH�t��IHŁƷ >*D��LX�'s�7M_Ӧ��I�MJ~�s��2	N�PQ��֑L�)�Ő��?���z�<�p�ֱ�?9��?)�I���O���vOʈ�Q(�'>U��R2�ʕ���ԕt-�}'Y�i�^�CA�2�pL�-�~��	��>A�� #D1l������R*�\�sKC_?�!��ş�[	�T�t� ��КU��Tqv��;xn8���8�8�@��ѓ��tlƣU��y��)�'6�l��i���� 9 �mѶ��p����3�'B�'��;���'�)Fxx�b��9Ȇ�HV��@��p��'��r���c���]�����B�D�	��l�ypN�[5�1x
� R��Bm���F֦l-�G���ؙ	ׄ�0��O։	��'�7V�n��Zr�G�k.nh���	>G!���0��pB���V8:�!d/�"!��R*L�2�P�NڃI~zlPq��y!�����M'�@9��[;�M����?)�R�aeg�o�����
&�,�����{{����On���K���$:�|J0�X2��!��D�o�J${"g�'��k��I@,ٰYX��VH�F�˥*�&�Q�K"��O̢}j�G_�g	~��b.��� �c�b�<Q�L��;V��&G�:(�v媖,�y���H<�IR�{�ъ�͡&�Jǯ�J�<�-
� ^`ܒ`�G���4�b��a�<!��;4�� ȣ�
S��Q��a�<��o��0�Y'�ıa@��όW�<Y���:c"�I��L�/puy�&DQ�<�djJ�3N]���):ێ�+��O�<y��
z&�032Aʟ?��p�H�`�<#Y:ofڈ���G�l8s��[^�<�$�M�5���@���Z�X��E��]�<�%�������$Sd�P�"�V�<�1��!<���5��1jQع�*Gh�<9��K��D��`-�`�v�[�<1'"��z1"IV��R���A�DY�<C�KfY&���AԘ�X�!��U�<��P'� ��&eq�vYA�O�<���I�|����j� t:Vˀo�<�1�Z(C8x��w�t�yK�g�`�<�NQ,b&�JCF�''�J3 �PT�<�Gk�+p|��Kɹ:Hɒb��Q�<9G�#S� ���W�d��D�I�<iDk٦2o�&�]�*�,T@�j�<�1��2#Zz��l���0��f�<)� �;R9E�2��xopW(?�B�I�{N�᪦���6P���G�\
�B�	a`L(��b"���WA�B�J���gTw�4<���UH��B�	�����	��{QD0�j�:|�PC�	�N���A`؛;���iV�C�ɭz�`܁w��,�*��2�X!�Ě q��P�m�*Q�Jt���];!�D�n)&1�f˓5���ï��."!�� �\����db�t����.	F�1�"O�iUM�4�B�j� ���fD��ˬ�"M֪�<X麄J��d����j2��Jj�F�� E��yB�Y�"mF������'� mĚ$*�n�+ހ8ce&ʟ Ҋ�Y����m֝�Z��ߝwupf(*D����Yl�`|bSN;�Q3�i�z!����j�k�P*���*i�,��k�2Af�iAg� $Ga{B.�~����?R�4\� J�-(���g
�vhI�
O��1s �0b�#�I;Dж���0��, ��ܡ|CTm�ud>�S<"͚�ɣ"C�"��u���JB�Ip�Ĵ�
W�[��a`�j��V)r5sB\+/)p��!&V+�*'�g}I�8A�=�Q�ɥf���I��yb�YLVm)bm� "�)r�d���M녁ЊmŬ�@,������Ѡ͎�b�<�*5�>!�B�퉇%F�#LG@��;ƈS0f�� �ϖ8Q���wdP�O8�;����0䄁3L�ڄ�H�U���'��13G`�c=JU����?).;�S�i�T���H�G�":�Y2
44̆�~���x���2k�Fp"x�@�jJ�"��O��Ń0�i� ���'\Z�!E�Э3sǹ&�Z8k׀9�b縵 G�Ւ+�F�P孚�d@Z1`�˧Y`^,�g-^�xJ�A��}�	Ǔ7�J���.@(T��J�DRݞPE~R
7�B���`G�P�Z���ڻ�M;��^�"^.�/QY\9B���@��zu
O��6�]�q���C�c{�9 ���!��TShJ���OH��g�>�S�˓N���B��.O2��u��
ye�=�@�'�V�]?g�$l�b�2 ��Dy�@I!�D�(+��}�|��L���ł51d�i[ճZ<"?�P���0@"�d�-+zW��&��6fTF��2�C�-�Q��M��Fb�h��n��}[af�&�ZE;�HS��~"�ݴd(���F�-N�шCa��DG�wBlp���V<Js�	�fJT^�����i�XO�) �̨�A��Z���,ܰBp΍��h�*,�����������8�ZaےsURt(� 
(
��ד�yR	��]LF !�A>��X���) ���h`����V	��}TL��ŕ�I54\�����jq�'��}�I-���C�I�+�P3EG�9s�T����Z/3:N�GfP�Ek�"?I�
��oWz��u*�r�,X��٦��]3�
�!A�X �a���>�T��O��3D�t\�K�	�)�Α"��DP��1K�'9�`���ڹ{e��C�OړG0
ْ�O��)G��=R�=�U���\�0Ubu鉴m�h1��4�2�ؗe��)#DI�d�V0#K@��&˾���4N��-vQ��p�`�Dt�b�0�{���.5�N9q�Oz��0�鉊{�8�$���JN�G#��(�l�R�X!}r��Yn���#���jq$������o
��E�;t޶ܱ��$ߟF�>)�@�1��x�v�B<I}rp;�� 5��a�6N�$_jz��f�?�. �3 S�1�&�P��|��n�!Zl���Z�*���o�%���$��[V\s�iiO�P���Ht�X�PQ�3낦�~�"�Fh�!��O��2҃������-��5B�)�><&�jB�/c��� �f�m�l�O��'�
���#� /�x��i1�y����B��	��j�
��	�"�q[�AS�.q�u�Ɖl�!�דk��ݩã�¬8�L1��Qg�R��!��'�z���*��9��="�eA&�
T�� �v���I��FL^�'`p�_"
S�{3�]�+��(S���>����g�'l\�#MQ�:� �r�	�>7<��ٴ
�����ZS�Q2��I6XѨ$�	���;�c�[4�Q�2l \l���2`b�K��{���VAJ'�P��'tܹ��J�:@��BU9p1ޤ��$��A�JQ�$� �P�S�]I���q��q2��P�n
I@M�@�'��Di�6'�t]���<�&�ѿ�hq�@�u�'C~0�K�$��.kƀ�a��D>J!2�jX2Q.�����n�b��pď;�A��q�����!�(N��)r��O�yЎ7�	��X�'�R�BņǮm�>mAU�ݞc���1�v&��x��X<���x#%@3_3Z��_�F1)e$�>�v�����Y-z�-o#����	�eΤ؀�o���ΐp�m-y���,q"��?#���p���,3h�q�{�dH���mT�\����=d,�PC�4�PxRDǯ}��1����:"�Q���%���>" ꉂC��"K���cO"���t�T�Ԫt`�*�7/��jХ-�y�(�uy�l+�D"��Ȕ��y����2��:�p8��6�8�ȓ&H����T�@�60H'A�Bz���ȓ:�n�!2��.1u���q.V�'�ć�f��,���4��K�*+����S�? ��+�7K,x B����z""O�@��-�n���q��ۢ=!*s"O���N=MҾ�ڲ�
U	���"O�)i&-؂#����%R��h��"O���E?`ȹ�B	)8�X���"O���5�Ӡ?T���^�S~xH�t"O�5I1�E�:)*��U�F��l�"O��2�Ŕ=�J4��>�*� "OV�X$I��(�!R�G�x��g"O�-+� ���ë�	4A��"O�a�U�ֵn�$	VZ
�}��"O�j�	M}<���Y$v謡�S"O�poL)$�]�$��殉�"O�ic ��!>��ٰ����u�Ԁ9�"O ��Vf�p��\��"E�3��1�t"OX�@M!C �x��
05��Q"O�)굍�"DDvE��!*O#���@"O"��#&�1CJ�YZ$ .|�a+B"O�a���	x$�Б��Â ?���"O<��i��Hr���$��i>"���"O6`{p��4�ͩB��d�
Q)�-6D��Z�KK"js��a�b��Sɨ��l5D��+ff":���"@�/Wd���@i'D�D���$�p��r��+z���Icl1D��me8
�B�L�5)��i�cC/D���C䉨A82%a�B�apg,D�\�#�EaZ�(���T%~Ux*-D�C�
�-D��Z$k];u�D5���=D�di3*^[�j���䜏?�>b�,6D�åˁ�c��0X���'n�Zx�&�2D������N���2
��V4H�r�0D�h�	�s���҂$�!1���S�O)D���P�G�P�J)�b��/o����,D�h���<J��������lA�c�<D��(B��%~lvģ�I�65�Z�u�&D���▸\J+�)G_e��I�!D��a!��9�0��F�uߐ��o4D������	+d!J�cG�F8�$�P�0D� " I��u�ܨ�5K��71��p�!1D�\�4OSW@��AaU#�F��#1D�pY��]�g3�tÆثd�B��&K<D�\ba�ȍ+�P����=s�0t�8D��[S�٫�V�Cq�8�|��-)D�����B�h8>��ɜ=��Px�+D�\`�B![u��I7�I`܈$D���e'�/S��u��<����4D���b�:5˰\��/��0���'b8D�0�� w4B�3%� 5x����j*D�����m5�!��A8W�t���K>D� K"m�����Im`���=D��ZuN�6D�� lѰEg��q��;D�|�W�W��i *R)IA��<D���E\&�"��6��	>'< �#�6D�@�f`F�y����J`M:�9D��a��]�d	;Ì�#����n#D��B���
4ힰbv/����*�-D��&�P�*��b6H۬����P*D���a�"z�PUꃑX�����5D��p���l p(��IC��v��&*2D�[�͐2���KD�i�r�T#2D�����d��V��s8�!H�D5D����G�$��(�S8,��*q�1D�@��h֞e37ID-+yt��է0D����ǆ�]g`9&B��X�( �3D�� ��B#�]�:B�I����=H|ٶ"Oq���> 6�y�O�2H/����"O,0`�H�%O��Dؔm6|q�g"O��m��d"�չ���\,LI�"OP,	�ȓ�z�azǦ��z�vx�W"O�Ř�-�]�.��ȅ$��X+�"O�08����7,X�"#��~�a��"O6�bUD37hN�3c�2�I"O�M�F�܏C�~�����2#ʸ�"Ov!�'���H�)��˪	��
�"O�-hЂ@��ȕ��ס %T-@"O�u�t>d�����=���"OF8i�����p�F�h�x���"Ol1Q���T���b�L!v��a�s"OH1�� sF�,�Q#p,���"O����wU��`��ʹ�Ĵ�!"O�.OP��u�d#�r�޴�U"O8
� ��deaR�" $�!�"O@����8t�D1"�ؿ㔨�"O�����[�fA<YpD�U�ܔX3"O�)�䈇.�l�q�(�F:y�"O.Q�ADP�_=�	��EZ1��Z�"Ot:�o�*�1a�Ŏ�x,�Kp"O������?���s��!P��Tҳ"O�0��æN�ı��枸9���"O���Ƅ�x�!Sc��j.N�QF"O�!2��_�pA ���uq�a��"O T����Ft�9�&%�7tnDQ�"O�]���1�@��[�m��"O�zg��V%V� `?$
!�D�Oz�ѳ��'떤	 �>D!!�䚖m�T� �ȍ�ʹ��Fb��8!�d�8��x e@,I�H	p`��!�D���]`)Ѭs�~��W�=V�!�݀���I��@5<������6r!�Ď�N���V�Ԋr2���
N�up!�|\������s�<c&��1b!�DI�Jq�P�C��d��1��(�{D!�d�5c:���.f�ĔɜO!���)`
9��撧�F,Q�k
�'�*$F)���D
�0�|�@
�'�F��t�Ǫ]i��������'�E�ͺxtT�j@���v򊜨�'3p5;��޿Sx����vW�Qj�'9`���	�Qh�⒇e:�!�	�'�� �aG&bo�x�%�eGD���'nnYC5@_6z�4��Hqty	�'��sU-Շ��}�1�2Y����'Ĩ¦S�U�m$�Nyz	�'N�4d��7�A٦���",&|A�'f���G�Ґ<�6Y5JS���'��fCV�q[�U)�D̒h�}��'jXi�Q�֫r�*����KMz 1�'A���D��`P���8,�1
�'����iȋ0lLܒ��G609p({	�'�@��\��ƍ�<��1B	�'B����Z����Z7&���'��sQNC�)4�b�%z�V��'��3C �|�V!C��Y�ed*`2�'��`H��ġ|��|Dh�a�*!��'"Z�2ԠG���X+�f�R���'�����_J�Y(Ǝ}Ɂ�W�<��B�@�ޡrq'W0I� y��c�{�<ّힶ=�d �`�]���IVmAA�<� L�!�#D�.�T!�xiLC�"O�t�/amre �1M�T��"O>��K�-kBDL�s_�C88x�"Ol�N&�Dl�&�
*Z *��s"OT��et�$��k�:i�Q*�"O(R�o@�pZ���ܘ6֜[$"O�x�\�>��X$�X�
T"O��Y2͏
��=�w��$�1���0?�M<E��'��93,�.8D8:��T0� tQ�'���G_�]�� ��5&����	�'��J�\�!��r�E�  :�	�s�d�#E�P+GL�(#.�D�T�(xe��;�BT���`�Jh�A�Y�=��;�VA�1�މX) cH�	�q�ȓaQ�d��I�:FA! �˥^�:�D{B�'x��)V��?~�jX�qD��C�B5j	�'0@d�/����;S
�;;'8�H>��R�> �3*��S�и��nO1$�\ه���<ɆnH81��PEH
}���� f�O�<y$�F��U��L�����N�<�r�(��BgB��6F�M�-H�<9�ɟ=r��&� 5����l�Dy�ZZ��(�R��Iڐ2Ҏ�(��1	�$t�"OVu3��N��eذ�
�D(Ի��*LOe�Ѝ�N�ڜ;�
�A=�\��"O�x#b̄0��|{��\	ZM�2"O�Ƞ��T%a�ұr�� ?�:a�"O���s*R'd"x�2�JUJ�7"O�q��擩t⨙�:�#7"O�Y�%*ƯZ���g%E#4 �"O� �P#ڥu��9��k��� ��'�I[���)�!q��tD�d���:�B��!��
-�֐s�c̭s��-;cK˜��	Gx����k�&���[u�Xq	�2D����W:D& ���"�2x�#w�6D�h��G�:(HB��Y[���)qG�IX��(��u����BÈ���e�Y'�X�#"O,X�矕}㌹���ˋO��j&Q�:ݴ�0>9�'��F���ʯ�hI�aLz��lJ��i�>���/~U���,�=<�	��'<�c�dG�1�5XU�ϺAbƙ�Ó�hO�8y �M9*�+1)]��F�"OP��K�s����%�O�i�5Oޜ0,1�)�dS��co����x��FߌT����ȓmH���EO�yT�)r�	{c4�'��#�q�ݪ&��`I���l:;]����l������)]�v�z�����(�CuK�J������ȓ.	`x(���Q�
xZ�E� Q���^d6���n�P����
�VdDx¦VW8�<�慑�X���K.@�� � D���uf���b�z����)j�ȪTD;D�l2��W�89���O9!��ãB9D��߆b��1lM�#�\�� c)D��c�P11��1�$
��E�8�iǆ'D�ĢÂ�:�D|��ԒQ�(���g#D�,�b��/)���N��H�x�O,D�\bp.عK\吕m��t�
Y��l*D�����~߀ ��΋	���k�N*D�, E�M�R9�2�
�B��x)D�88�B�r��Q!G�<��T8��(D��7CݒoךpZp��4j
a��'D�h�p�]�I^��A��1g(% o$D�ȣc�W	����#�-^ܴ�5h'D�� ��Y�ˋa���A��!L�6���"O>��'�R0�"Ip����k�8uqc"O�L�GT E�	��	 K�2���"O�H;�(E@�M��`�-OQe�$"O�ᡣ�~�� +��E<TX[$"O�� C‭'���J�F��Ԑl��"O�LH��.r`�Ae�J�]�
q"O����nL;Y��!��"@�*=�"OdH�Ի)}���"Cs��Ɇ"OV5ц�D-%ÌScd[0�h�zG"O e�ӃF	`�0\�w�,y�M"Op]�B%��_��2C��0j�KF��y*�`��u� #��(r����y�!F#U� �J�܆}:���W��y�e��,���"�7x�X�E"�yb@��`w�	�mI�o[���'��6�y��Á�=HB�\���`����yB��{5� �% �Ɖ���P%�y�Jý,����N_
z&�5R���y��3+}�q��ā�pO]!@�Z�y�� �ֆ�r�gV�X
l�n��y"�R���%��J�#U�� gIB<�y2F�%�$�S\i&��R�AܺG�B��`҄I�sM� 	�Q���n��B�	��dAڠ
�Wd�a��ݱ#C�B�	9EĆ�X��F�}$����e�B�I��R�[s/�x��"kN�QFC�ɻvo
1��â6r�!� #!�(C��%/���XY���)��6\B䉪�  8  �Ϻ�
�$ı�ȓA���H�	S�Bp���EP��(��.n�9ۣ�܋l��Ȉu��e�X�����0�R�<oX��Z�k׮���O������/W': ��f�?����v���7�%Oz�����
P�5D�ibn'k��u�Ý��{6�5D��'B�Oq�� �;����G4D�X	���V��\��NLV!H�"7D�t $�����0nH$��i��6D�P�wO� B���#��#���R�5D��jT�?G�$Ȗ� �*�$X���4D�d8u��%�<	C���7��%u�4D�,� �Ⱦq���A�v'�uZa�2D�8���EV'��H��G@U��/D�x����e-"�pŕ�M~X ��./D�L��i�V}���A�X�)�(�AЩ+D��⫋�KY��2�"RA��A#7D� �q�J4qo���ԡ0{ ��j$m!D���,
�UL�`�N��p�0��C%D��eOA�� �p��"�I�#D��!���\x��	B�G�v]��lo�<Y�$%e:�h\�=�x���i�<����?�~ cƇ6?���@5�P�<a�,бpHL�b�m��t���GJ�<y�/J,NC<�Ǩ��~e�X`$��G�<1��5q����@�A7P�H�)�J�<1�eǥt�8-��,��&�$3���A�<����c�,�x7�	�+	��ڷ��R�<QE�@5'����NG���T
fčh�<��e!'�(� A��nH�I�/�c�<I��ʽ	 y�E����e�?`!�z$v3�j�5�E�D%`H!��E"����v�]���7o�!�D�.�<̫�+S,J��`b�^�{!�� �@I��ָtn�CG��J\"I��"O%(e#�`� ��rU�KX@Z�"O�P���2��� i΁a�H���"O����*�"�8k��]���H�"OX|2N�(]�:�ys�vh�#`"O4��w`@�k���(A��0M��Z�"O��q���,��g-�.X�c�"O��A���Co���LF�qT,bg"Onx	L�X_p h��t��6"Olk&)��n�6BD��6O�y��"O���Ŕ�(X���CS�>��"O�$�B
_.A`a�Vd˙��@"ON���`�3CX�<�F.R=aH�y�"O���C�Y�6���ʠC_p�|��"O�M��ŉ�MЄ�@H��:�Xa"Ov0��K�"~p���g"<��e�"O@C���=�t@�I.a�\\A�"OV��W�Ɗ�eKd�ܿc��`"Oy�@���E��h�(J�<q!�A"Op�V�֣&���rNĕ�l�1U"O��S̀]C�ֹ�N���"Oh;�m�E^�A��ݥ'�d+V"O�1����O ,�����Ck���"O�@Q �@5�P�Th�H[9H"O�i���^�~����M*K��B�"Ox�@� ���S���&IF	�"O�4�e�G.���]	!0�Ԛ�"O�]��A4G��4��K��+��-��"O�b'AG# . u��ەW�["O������g�*��D�a"j�"O:L�w��AT���B�2}k"O�(����}�ĉU+�w�b�"O���tㄟ.��5�"*ä�H��"O`�: �_/O^�؈`��/ ��ؘ�"O��
V�R7RI���Ŗ�4ĺԹ�"OR��#�E�����) 4��Z�"O L�f���BJ\��TN��<���"O�1[׬��Sts�̢%V���"Oz�Dbޘx����*�<k &i�"O���� Ԃ9F.�&�ҙU��X%"OR�s��AN�`�"I�/����"O��#�		H.*"�HN�?T�"O(5*Qn��M�l�Ҧ��.�v"O�����	�bJ3�[*\X0`8�"O�qcV�W[,�8'�V"FP���"Ob�3�B`��b Ѫ���"Of�ҥ��Pk�a��\��*�"O�I�T�@n��h�ĭ�\��J�"O���j������,N�J�x��"O�	(�
Y ���'K�.f���f"O.���� �x��7�҅;�ةQ�"O̠ �JZkh��ZH�ژ
$"OF��D�>`�d| �h��n�"�b�"O�D��ɥs��!��<^�^�e"Oޅ�GM�?�v��6��/'��+r"O� k�1�F	��	�_:���"O�ɲ�-�^�tq&�۔d����"O���/CCh`q�j��=�JYZ7"O*5�`�*��`r��@��i�"O����m�X�M���6(�>�J"O��i�*�
8���C���?̘�h�"O���d��)�]�Ǌߨ|Ȃm�@"O�TiR�,�Z�!��+w�\�c"Oj48��ԏd`�1�
�I�t���"O� B�r��6�\����O�O㒡��"O��@��J�8�"���h"O�k3�ǐmd�qXs��7��p"O]Ѕ+Ӹ	gT���12�ȩ��"OHԡ�-_�p�z��E)U�i�N98�"O���LO>r�z������:��M��"O�|�u�{��p�Յ@�J�Z0"Ox)y�d�DI6a��G�\���R�"OH�u	�Fː��c}���"Odmӕ�%$\*��ө��CkzD"O�� ��P�vt[pi�as HJ�"O����]>�>�K���j��<y�"OB�HѤ��$�l�bV�T���a�"Oh�xg ׮�4: ��l�={�"Of��a�$4�,�hh��_���Rp"O�4x���A?<�X�L!��ّ�"O�t{��N-f�pA�$��"7���"O��p`��3�9r�c�&S��q�"O��;���K�`��@U�2��"O����Ų'(ST��x5�"O��c���5Y�}A�ƈ`�,9r"O$��B��[�@�(#�J{��2�"Op�J�1yo� ��V��|��"Oέ�,Y0/9y����*3"OŻb���B=�a�]� ,LUK�"O�h`qM�&��hz傍N$��Q�"OD(�B�l�z%鶧]J#0`�"OR�b�,�+@�WE@2�"O���F� !�V�؉T�!�"O�d����b��\�CK�h\e�a"Oh��tOI�p����P�_�t��"O��s�����n��E�^���"O���LDL,Y��ݝ/��P"O�}� G93n���`hz4PSf"O�E�"���n�a�'W�H���!U"OR��e�H/s�(9�ƍ^�l��"O�tx%�
K�4`�g$⒜�"O�̪�</�� � �_z�dܣ"OR(���K9d>���F�#g���a"O�������%7�	�qeɞr�P��"O��EN::�0��I W�0A 	�'g��t�Ш�-ɫ�Ę�H|��
�'	
C�P8Қ�vO�4��Ua�'~�L`�	����(��	�����'[R���턇�x@"��U� ڜ	�'G
ݙ/
�,X,*קQ�{~���'�d|C,�6Yj~��6lMu�.�x�'��(�E���go���F,��pkp9Y�'P�1�$Ł�? t�LT�i�P�'�P$��@>��BI�Oܠ1	�'�~ɠ6��\"0�'�W)y���'�^�2�3�"������LD��'�8P��d=>�.����O��]��'z@A��C��8|p r@�	����'F]qG��8>.���!+�.L���
�'r,s1J�
�Ç��	�ڐ�
�'�f=Q��@<hb������'?�e���,e��e�Æ�-�x��'�ظsuΝ�O�>D��)�p���	�'�Q�bj�Og��b��@I\X	�'�°�ɄD>B�;5P2e�`��'Txpk��b�jlԴ�( �'��;7!ҜMúI��C�3��k�'�4yW�D�M�0ɉ i�,�T���� ��$�>d���)N�1z�iإ"Ori1�J�~��Ã��l�H�"&"O��)AZ�?�>8�w(�&#��+�"OL�d@ v*�j�%B<Y,��b"O��yRDC�%���@�Y�"�j��"Op-H�h�vϬ`�s��!�`�2"OtI�#3E���@��!����"O�X�!E�WGRqcՅR�)��h�"O\�3�eLf���o��pt t"O^��a�Q6��B�S�s@s�"OF��6n�
�e�#F��	Q�xc�"O6�Ƀ$�5Y���Wok,lAA"Oli7M%r�N�V��ln�"O�MbwA}B>`�'(�hLi�6"O T�c���j�͍i��58"O��s��;]
I����p���h"O�@�S��@��r�tиM�"O�y����p�8X��E�V��\PF"O 8PF[&BY��ڔ%�3(���"O��*��p��b2�� �2E�"O�Q�'5f2��q*ǀF�*�[G"O�(�-ݧU�*�+�ϬmBΉ*"O� �f�AHI,!�na�S"O�B�Q�q�Q�!J%2��"Oh����8YY��T�խ>�����"O<hS����PjU6]�(�H�"O����$V4_��]X��/{�v���' >��&K�>��:���H����'�3K疕�c���Q%�|4kՑ�y����k,<UP�i8F�|� ���y2��%5<�j����^�����yN� �b�#ׄϬl�5��Փ�y��M;V�n�Љd$��xt��7�y��/Y��=H��e!�
 /�y�'�`�P����DhT|��W7�PX
�'x�pEa�2~���"U2�T��	�'�䑲 ��E2R	0��K5Z���'��a�EFП���A��Y�X��'��Ȓ��\��ج����(a�j��
�'�4��w�@�n`8�1��#����	�'���#��H�"�p���	�'�fIp��W�y����,
V�-y	�'|Vl�p���Z�S#A1Mݠ�	�'�t8r
ݓs`��y3E��Lp����'��Ly�SR��XG�H��"
�'����.��h���
�@�D�!�'`��/]%_�>i$!�8����
�'2:)���m�~����G76�Ԕ3	�'���{eKX�CF�W��T��'����g��5ё��R�`��'1�i��!S���`�5�GDܤ`��'��L���+��H� �M��x�'�b]� �@�p�%�t�ˉp�aH�'��a��-Ȉwe��ٕG�g��3�'������=?dr0�压=Z�d	�'��A��0j��p�$�"SϪ0��' ����%rD�$��	�Y����'vX,�B�oS^��LS�C스��'8M�Ҩ�`�0}8�kQ�83<h�'����"��JK���U�ͨ.�P��'��!8q��Z��@��$���'ܡ��C6r8l g��s	��2�'i<c%ЉpOq��C�l�|% �'������F��7	�j������ �%A�
�!"l���`cHXg�`8�"O�æ�D�d64�9��K$9T�-Q"Oz�9�O�_~�M�������"Ol@��]�~x�h(r�Ԙa�|���"O1�dg�tV^y�
�+&�V�zc"O��K�-?Ÿ�c��[r걛u"O�B�m@D@�P�l��}nM��"O��h��%S�H\#���0^
�� "O��9���X�ƭ�����/�Ȃb"Ol����8���#)R:,B�P�"O��C�lF;p<(�Ԣ]90>d�"O�5����bH��2f�׮~�r�"O�|���0��Å��9�V�"O��:t@X�fI4iK �1]� iS"O�J�!�D�r}�Ӯ+l�-P�"Ot��D�,�H=)gEJ�M1��H�"O>�꧌"�\����)
��"O�����CG����8�s"O}��I�z�U1�g�O�)p"O$\H1nQ�آpfüc�80b"O�4P@�<.3>�£T�@ð��w"O���s�ǧΖ��gƯ�`�A�"O�5!􍚋.A\թb��X�tՋ�"ON�DP�s&����[�"V�a�"O���X�*f�y��\h]�Q"O~P�IҦy�<�`�!P�b���
r"OA��
� �0��q (B,p�7"OPR�Å�q7B+r�X�"���U"O2PK1a^+9� 5ǐ�O<l��"O��h���:�8i�W&˗P1(��"O��㠪�$!�2����.E'��t"OL�q3N��u���%���w"�+T"O�}���A�m=�h3�AHT��p�"O�,�oĦ"c���ĉ�q�"Ova���E?�|"%/|ܼasC"O^ҵ�ζm-���n��Rے�z�"OٻS��|��؃��I��TJ�"O�<	����R`*F�O�o���5"O:4`��!�|��L�-�JQ"OZ��S�B�d��˞XJ$	ٵ"OJ���9ޜa&GI8b)ۤ"O��x&��rKn�1eJ�iӠ��v"O&)ɔ'Ō5^���Ѣ2Ɛ�t"OTU;2(��_�IsV➍I�X�`p"O������0�� �!09���W"O6��-�h�*$$�\
�"O��kq��;�
��G�K
L���"O��s)K�&8��%Tw^8� �"O�p�E���Vn�H2@$�#R&� B"OHAgF��D-�,|PCͶg�!���m��lb��*$0���3�!��ۿV�t���M  }@��� &�!�dKK��D �b��P:�yI�mۤEX!�$\A���11�H)P(x!A�0O!��EV���&i�o�,`kH).K!��Q�;I��"#S~5J��JA�!(!�P�gnD@@��"=%���U'��D!�$�IJL�����8AhA�C�n>!�d�!R��*p@R�k]��I���!��A�V���$	w�=Y�L!(!�$I�6�ƌ�`ݎ._�C�� %!�D�97 �t����w��Ţ�R�E�!�� D3XI��-�l	�l�7Q!�Ԛm@
\����Z�n�+��џ(j!�� ��ЅK�N!��(�+|��"O�e����/>��3��Ґjx����"O�����P+�!*���0t<�	�"OX<��"Y �]i1h�:��	�"Oj��G�B@4�pݲzN�:�"Oz�z%���~�(�%!���,���"OzPst&۟6��8щA�{��}iu"O@�b�C;Rq@�8�M��u`"ONU���ۭ4�h��ۿ!nN�"O.�qr�����X�'� )��T�"O.��n�#g�p���M���w"O�`q�(�/K$�`�A���aE"O�CAK�,�	�AM }J�Hc"OP)�U�ܩ�ް E�"O;��3�"O��3F�ƳVU�F�K<Y�p$�"O�n˫���J�܆!^(��"O$<���F$d��h
�"R�`b&t�"O�!x����Q ` �C,-�"OJ�2�L�J�K㯀3��]�F"O��K4 Z�)�|l��lG�x!�y�"O�͠�!��~��$��
��"O��!2��|4����2����"O֔Z �̩<�U�l�i �9S"O���E���ۨѱ��X��D`"O�YPtm[��!	��ӡ)���"O��"�2\Oԍ��D�8�ZT�%"Oȍ���4x�r�l7.A1r"O�M�A�7��p! [.^L0�"O�5���B�ev\��\�.��Ŗ��yRGJW�1'
Bt,��S�D4�y�Jƞ+�H�"@@M�}
��a�!�y⭙2V�Fy������#Jt�!����+#kG1MF��G��
Wu!��:�@���
�<v�g��6s!�ğ�~�lE鶬E%���Ȕh!�d��`N0����N!D����\R!�Z� ͑�q� 9GoR5'M!�D
.\ܹu�Z�B�6�)�'��!�d�3i�9@��R�i�H��Z�\}!��O�sMf!� @u��	���|d!�$�>&X��u"�':�`��T��V�!�]�cr�8��쌧)9�U#��U;FV!�|������)\MM�G�6X/!��u�����\�,��@��!}!�$R'A�PE���
m�ҹ�b@��pg!�2sl�m{���N�� 薏�\!��&# eB��?y��S�#I)!��_H�V}bjĆudX
���(up!�D	&=´��-�Vl��8�L
�\S!�DX��>�dh�	*6�!sB�	�!��2ai\t�iJU�M�Aʏ�8�!�dF��M"Un�l/�X�`��}�!�d��#ҙ�CJ�<i�X`i�߽}�!�dT'��(�%��~�22D�& �!�d�?� bb��;|�,`!�S��!�� ����r��� ��|�@-R�Ji!��לG�&@!��	CMU�-Pgo!�Ⱥ� <�Dj��H2����l�#�!�dR�dN��z�������"���b�!�$�)
�4�a m�%ʰ	R��!�d�0Q�Dß#ҍ@�(\�!��ȹ8�p���Q1�����y�!��$�Q���
2�:���e�?�!�$J�B$�x�Tu����jE�!�� t��c׻y� %JC(�T<��H4"O�U��Н��
�G��:D��"O~Q�f$U<J����FY��ZH�$"Oؔ���2�m"sK�3*�VUҤ"O��r�U��Jܣ��S�B��"Oʠ�C.Ϛ�P�$p�6l�"O�iAE��/l���#&U�(����"Od\��*B�O��īA �<�2��"ON4��J4�ڭ��C��>�l��"O�鲄C$Xl�  E��B{���D"OeK�3QW"�b��<ij���"O����D�xuI�Cޗc��J�"O<!#hǩ0Iz��6uP4�S�"OJU!7$�,�<�w$��I[b��"O�58��,0�i.K-B?D�#"O� e�Y�vx��p�,=��"OBÍ�R��!�2KۅJ!��f"O<m��_�mx���iX�@��K"O�L�S�D�}:�E���O�PU"OJ�QB\�0��?L�ܵ��"O���� �9=7�Y3G%�N�t���"O�d��H26tv�HTcÇ{��;s"OT�����!{�Q�(x
԰r"O���'��th&u��%Y�I\���"O�����2f�p���VkEZu"O�1�#�!2�1��CB�~a�+�"O�����+k�ܡ�B���uT0�U"O��3��>@� ��g��}^X�(&"O�0�7"L'} �hf@Z/P(0��"O���@�_e��Jr���S2�3"O�1*��4H�ࣧJ�2Q�@�"O�|��
�A�����2D��"O��Rǧo^�D��@הJ��	�"O�HSF��9|k:4�.(���q�"O6!a��C(�Zy�P/�����#"O��ʠF_�e&�}����:0*l�a"Ol�� �l� ]A���7��"OVY�0bĘ]r��Q�IP��w"O�� �Q4+[��2Ô��hI��"On<��Ð�Ĩ`�↯F�~%`"ONA�$|��$�@H�0ZG		��=D��{���6;44�͕#X��Rh=D���u�
�l�ʴCDҡj ���A.D���P�.���	��+~��`©+D�0���)]�ls�gğx�����-D�8��(�!O �m�@Hà��!�-!D�X"�K@��y���Rْ�>D��QUi،j��Ys&��x	�(�s<D�<҄��@*Q��)�lc��f�9D�<c�A�a��Ð�0*��H�*D��v���h�C���7�`��ê(D�l��l_(P0�R"�6uG��1w�'D���ǋ�v
,cC"_�
Į,�q`&D�0ڔ`��TSĠ�0Q�=��ъ�%D�T�f��pJ�-���w�E�"D��kd�!-��)�&�^�� ':D��X��s�=�@Dܲ�U$�"D��JΗP~�Yy���gV5���;D��!Tc�;r�8�1�V�h@
R�,D�H�ᆁL�lD��O��A�r�2�6D��Y���sv`���
(�Z�{��8D���B�v�0l"�	�D���7c8D��3d�S"5B�h��ǘS[�DZ��7D�ءGlϯv�z�#AJ=|�����I+D�� �]�E ��+H� Ae�$a�Ɣ$"O��� ȏf����q-s.��u"O^H����=b��x�l+>��U"Ov� �ֆ.5�ur��lXp�"OF4�T�	�A���GO
5�R��6"OL�	� �d�}��K�8���"O���uk�6qz��B�1e{��HV"Ot0�KB�8��%�N�aa��"O��HL��!�b�2�a�"OL�jB#�6����A����4�4"O(���.-I~X�A!�M�=��"O|�q�AV�3}���fnZp�D�qr"O^̪rB�b^�1�oԖ{~u"O�0x�(QMI���S's�l2"OP4i�&�&��U��J\f�u��"OtI�!��V��w��<Ib����"Of���.E�nL d0�ָ=WJ0�"O�\:G�M "#@Y�%BI�\;�q��"On����u�F��
;�y0�"O2Qb��֊v�.��pƏ"5dȧ"O�R��.������X/Ι�$"O��c"�FE˒IxT�q7h4`"O&� ���Dپĺ�
m���"O6Hs��P#|��	�v��0/����"O\\Q��V�$ 4����=^tX�"O�y �#q�(H���Ψ�Yq"O&�E�y�D1c����+��)�"O��%Q�F�H�*@S�b��r"O��tK	n���Đ.���H�"O4����7m����$Y�z&��S�"OF) ������y�BD�m
"O�q"�	�R$B��P�N�f�6`�v"O:}SeD�X"DB�,#��`�"O��۴GC{A��b���J���r�"O��!���`pf=�0�R"<�7"Oz�e���uu6I!Ǩ�?iTa�"O@d{ �R	{�PD��RZ �`�"O�5
��W5Z���e�57@�Z@"Ob=)ţ@z�ڥx�%��[4� ��"O�T� �H�'u���S��{ 2MV"O�I�u�đ2� q(NC��0T"O<�uI؟\����(ߜWT+��y� ��$4��q�TN���D��y�$��@8��ߠ{�H@�%���y��Y����5�Gu�^ �L$�y�BX�(i"�77���T�,�y2KG#�����J�1A����hޖ�yB�8x�t rĄ�~��� �Bڨ�y�h�;}e��OH2M} ���ȁ�y����l���Z�ӓ@�rIc����y�L�5"�U�!�D{D�DB��y"
�j�x��g��B�����Џ�y��,�,`���9�����yb��ln��a��ɆɣS��;�y�&�"LK�dL�oL,X�+T,�yB�M?8��݁�)�*�b��ᇨ�ybJہ3d�Pr�Î�n�i��yB���x��M��F�4C�kɆ�y'"T�X���Q�=�8���ݨ�y�@ԫz�.s��>L����%B��y�a�"stZ�b��D������y�F�^<j�S#�;Fl�Z����y�DL5R+�ܳEIǊ0Z���D�ȁ�y��D�>��[3쐉/\�RǨ/�y
� �E   ���$��*K��õ"O*I�6�J��ma7���:�t:�"Od K�덼��œ�܏2P���"O�C���S(�E��<���"OTQ�c�C��^���M:���"OViQd��y��쩅%��+�p��"Ot��ѬV�2s�D��9�%"O"���M̓$2�ydbG8cl�(�"O����cϪm���p���3jRJ��&"O� xs#G�	4��O��M �I"O$c�E<8����̯^>��8Q"O�5���hԐ���e.��Z"O̙y㈅hu68P`m�{J���`"O�uK A���;%�Ƕ0[ 	�"O�p�B�17*q� ��<i��"OJ�KIO�X]���'	
,�"Of����F���Ua-5fVi2�"O>�&G6y��H�nNsI�8�t"Oj]�f��Un��L�r8`q�"O.��f��J$��� ��-4rd��"O��Z��Ѡ��Z]���p)\��yB.1��ٱ���$�-���F��y�B��H�H�,.�[���y�N�?*]P8pgLӄx��00k��y`�1i��0C��gt���īE0�y�iDjq�m�0�"	$��!�����yr�͹UQ��ц���Ш����y��M1n�*�H�F0ֱ����y��>;R�۰�9C�t��2��2�yYx�0��z	�$���yB���V�PxQ"��8�<I䈕?�y"�H#qf�yP�U|�c�A�y��8_�����$Z���� �O��yR*��pa<S�=m�>(�$]+�y"��Ԏ�0��T+n��TA��ymD-V���OH�JC��Fs�B��j��̫��L�Nu܍�K�A�B�	f*&���,���@�H1�"Ofy�q�ǐAԄ	�Tn�g$��"C"O��[���	@�6��R������#"O�L�c���89B�M@� "OtۦɏP� @ǐ+
欁�"OƥB�k�t��ٹ6	�
���"O
�z+Ąi��|�`�ߨ ׼M��"O
(����(��a�`�*	�P�&"O� ���ӪIf�$ 	3�10�"O~�W��cSX�S3�ÑF��|�r"O`��o-���-L�X��#!"O,��I�V`LA(�� >���"OZ�ZgO*o�L0��.)�dܺ�"O���B@3!��5���=B9�q�"O6��w�Y,b�BX	��'���%"O褂�J�������gS7m"�4"O�	;w ��8��"�퉐"ĥ;�"O����-�s��a��jߏB�6�s"O@�'�\�ҥ�W��^��)��"O���%ܱ
G��[��k��p{c"O:��Wj��R���h@�a���#"OB��r�Ϲy|��ʓ�O{��!�S"O�aj�J�R\�A[偏D�<)ce"O@H�`�2;��q��9�lm�c"O�	 %GX-|c`��L$�	 "O��CM;H��L8����=��S"OL8�q W�:��9P���$�`�"O� <��� ���z���9L/X�z�"O��:�,�)���p��Sf����P"O����]9z�ܴ�Z�V�J��v"O��2�Z2+�$�����~��+�"O�Ț����x�:(�,q���� "O�*'�Z Vv��h�M�	�:d�"O��"��"��Y��,Z��Е"O��*bc��� :Iz�=�e/�!�I$V%�U�mV1h��V�\�Gk!�$�M0��B$�[(:��*�%ѲHS!�B��8��G�
M�|���P�!��sx�����EZYr2�I�7�!�ͥ4�x�!�#V 4D�T;�'OI!�dA�RH�X�oL�Z�B)����"?!���X$�Б����x���&�!�$,N������@��1!wJ!N[!��ݸ^� �1ő�S7V�Bd�O	�!�מ/8H��u��!x�Ԅ±�F�5-!�$T P�-���1N�� !��6!�D �R�)QP��w9xLs/�A�!�"`U���C��%1��@7G��!�dH�|A\�j�@F��`c 
J%"T!�d�	a8A�w��QZ贲@�I�(!�M�tz6�Aץ��I��}��9d!!��{Ҁ�ZI�3uy~0�《�!�$#R�D��dc�	�*�*ABָco!�� B�{� 
:)J�QZLT!򄊻X�j=0�jX�b�V�0Ц՟S=!�D����-��,*�L��DB�y�!򄕣h�ĳ�-X�a���R��>5�!�CO�0i�ł�N��E�à�;]!�$��m�R(3���c��!�1�a�!��c�}h���S�9ؗ�U��!�D��$cZ$���΢H�2��v�B�%�!�$ٍdT:����m$8- B�]�T|!�D:b} ����78���C&H!��-Cɂ�z�/�.#)<3�Y��!򄛪a��ᚄ@S��Xiӈ5�!��'/d�1�)$0����
;$�!��(s
�I��a��,�.Q�����$!�d��4�Xp�`�$p�4���U�v{!�Š=��h���>hr}r���f�!�d�h˜��ՀT�ybP৮T.Y|!�$B/%v\R��=o8%����;�!�Ϫ
v�:"�L�KU��s����F�!�Dԯ%��tZ�I�yS��(��3_Q!���!&9P#i�řCK�}K!��Ur�a��½s�=���aB!�D �|Ų�t���>�` T�[%!�d��$u�i� �'�������t?!��."���U��Cp��J�o�/�!�>pޔru��8J>½����c!�
�C�`["�<	�DM!�B?
�����Xw.��XWf��}6!��Ίw�y���,u|�bN��z�!��")T�ː�ϙi�D8�%2�!����0��V�wRа��ߛ#�!�$�+2D ��Б2g�ˤ8z!�d�H�(��K3E��a��Q7;!������6�����O�"�!�Ϲ7�\TH&8hu����5#�!��	ތXWk\2'p�����8s�!��1s%��17�$:\�P�hӉ9�!��. v �h�!"O���f�"�!�� XP�8Dj"���vW¹�"OJ�� ;,Kx��Vl��K5ެ�F"O��+�
5|���
�Ꙫ#"O�u���T:/�#�*81��"O�-3Z��{���?��av K(�!��ťAs�ԡ��_�\�+�$�.T!��m�b s�ˎ+5~n����8�!���E��8��#W=9g�����6a�!��  G���W��2@��)8�!��Y�fNp��ǔo!v-���E�!��H�aCP��^q���Eh!�A
yi9�d�]�#�5���.vL!��'� �(�B8F��0�g=!��5|*F��Q�I2O�*1!a�	� !�Ĕ5<�z%-?&wTe1$�n<!�DL�>�x9*�,	�9fD=Ks&L�1)!�@�r4���CL޺Z�#�,'!�ߌ��)p�l��FLi P�P!�䊏hqm ��'
,m��)�!�$ J !Z$�Q"�����!�!򄟒k�Pp(��<E���f@�D�!�ѰE��σ� �� 4� .Q!�$�9j�}�aKϰB��ܨ���`a!�ށ~�@�ƛ�D���6-פ[(!�ĝ�|@��c�[�j�v�	qAP�_�!�Dڤ2_tXr�l5K���EA_�"��Dw:j�HĢ2
�|�Z��6�yr)$�����mH2V���w'��yr�tCT)���:x��'�P�yr�f��P6a��f�2�f/��y"���hl��(���'e�,��Q*�y�*�-=%���@�,L�^eJ��� �y�� &�A�S� 5O<�i��K�yb�E�PN�<��M8>єK�匿�y��1+�X��6�!��6�S��y"ga��a��ŕ7DI�����-�yb(�^y����I�"D$�`Έ��y2�W
ǲ��@��@�v� ����yb��~�=�a�7��|X��^6�yr�ĢW�Lr��_?-*�):�.��y�| ��lUS��[��"�y2��96 �w�N�E���)��yRA	�D�ј�� lR�,�F	���y���p�(�Do���Mp�`�2�y��X�,b��{���a\Xz0�*�y�
V�tP'���TՐ!� �ŵ�y"L�'U�*��O���� �B��y2)X�AK��$�U$W��W���y�M!)w@�L�AW��+�yr�<D�Kn\�`����&�y�(�4ǼT��m�1a�������y�jS�T&X���G�J��Bj�&�y�L	)j�r+ ��=��1����y򥁦&ָ�C�lX2��<A�����y�l"5�f�sc\&] ��D���y�d�'���sU�
$d�~��i�2�y��D�4���G�V=��j�n��y�J56-�a ����PF-%�y"fس=O�x�Şg"`��҄��y�j^��O i`p�q�L�y"j�e���ZE��2�A�yҪМ ��ͨ��� ����$����y���S�aY��W�e�ġ�4�y�G�/z���b�"њ�M�M�$�y
� "!����@��6����"O:�QC�Zn"|����5-�l��'en܀1nA�CNt9��A�HZ�P�'KL,АC��`�j�Е��S�����',D�2��u��r%BZ�d��'1�Y��e�-oV��b�/�O�Xq	�'�����%�3D�r���!�6M��l	�'��	�2(G�Sz(�)T"�?\���'`���"l9ۣ�7u0��	�'bl0�T+	,EvLi���,����'�4�*�+L�z��!!���u.4Q��'M\�Q@��]��%k'b��i�\)�'UT���C�-pdE3� �>[^�)�'�h}���Ѱkc�	��)X9}Hqi�'��HW|n�q��	w���'Q��!�e�	Kj&HD��#T,<��'^�`#m��`�~؈p����8@�'6Q�!��!G� H�7	- ܩ�'���q��B����{��)$^���
�'{r0(��2{>��ۢF���yp
�':-2BHcb,�C �5f�����'
t��u�2=�J�ZYla�'��,H �����;����O�jeB�'����0O��d:���F��A��H[�'��!JR�¹KSF	����Y`�'�5Ѐ%�8̽u����;�'�pt"Q�	R����fyn
dY�'�[*G��
S�Q�kͺ��'IH�����z:���F�i��1Q�':Fk�GH{�
��´]�ʹ��''�Z�
�;/RI��BЪd`�=��'�6<�B�[��9�Sc��U-:Ԑ�'=D�f�-�������`����']���� �%(��B`kˡVf&ܳ�'��x�n�2Ti���w*O���'&�{7�Q�M�p��B��}�f!1�'��`�OG�V>�H�Fn��{�]a�'�,T{��	58)���uB	���'��)�T�Ms�ԝ���I�g%PP)�'�^����sw��#�方q�@Q�'��J��> f�E`�,@��~���'ӂ����BB#��Hv�L%�Ȑ9�''aIaB�;l��ɖ%{@p��'��k���MK$Ó2�>(c
�'�Ɂ��9=Z�c�;0Z���	�'B�h�E
 �,lt�D-"-���	�'x�Pk�h͞R�,5��`K	�'(,��7KT(�ޱ�2�%�P��'k��Y׋�nҰѸ��1儘��'R�P�Ȉ!$n��A)U83�,�	�'r<y�@/"��'�л5C�0�'���!�!�/58vG�+9�4��'�0��&�]t��*v
�(_~l���'KB�J��(�<H5�����k�'�x���-��*� ���_�F	�
�'f�����=m�`���n���
�'�YZ7�ܓ@i�⃺�x��	�'�&8i�h|�v`YP� �3`
�"O�aE�hal5��E�7X���r"O�т �/��Ec�3Q��#�"O��C�e�
J~����� �jK��cf"O�����}Bǩ��,9(D�`"O�	0FÛ\� �S4ɀ�P.�=�"O����~.�5h�]	t-�"O� T8 ��(Pkr��S,��3"O�؆g2G6.4fIF2u��]�"O�%�p�ޭbR��{�hN�>궀��"OHAfԤNg�=(�U�Ol
0"O24��RF3T��℉MtD V"Opb���dt�剆D�8zS8X�"O�q�"ŻQ#Ƒjh���"O�x��Ӕw���@Q�L
iT�i-�y���4~�<P�3d�(y�~u��F��y҉@59�d�	D�Nn�`��᠗�y2�]��^��� � c��(�dj�6�yb��,,�d�:ҋ��1a&�E`[	�yB�'z�����扯  �C����yr=��#�ft�fdYDl��y"  #{�n�D,��:L\T#eM�*�y��J  ���EE0��IPaa���y��O�M�$� Q#a��:�yr��0Ւ��"���A��0�y2Ct���oG� �L����9�yb睋AP����_*# �سD�W �y��(b���D���#[��y��L�dW2�Jd�Q�
��h���ˌ�y�N��t
j�	i��@��B�y�A\;_ό�!"H�8τ�b!��5�y�ƙ�`��8SB�
��zp �X!�yr�O=1-�
D�����c���1�yr��5�< B7���� ����yB*�J�Q�C�(N9�� ��y�Oʹ^����E��~��M�2Ε1�yb�C#xPC�K�5��Q�K��y"��2uN�D�u��oQ\u���)�y�

��Hh��R�11�4 ���9�yb�H"TY�EM�O��8��[�y��T��A��n���ѳ��6�yr�9��1�uč���/�y�mՆ3�t|��"]�y�A�IA��yr���`��j�
�p�zi��)�-�y�@��%���&Ś�Pq�"?����|䮥���F�'8R�o�!IھȆ�8�����Ƙ�n{d��#�Ffq��mO�r��EADh	�e$s�q�ȓ"\���oC�H9FF�_��=��^�\j䚳j��`U��@p9�ȓw�6����Q{vmHA��A�*��_C�|�V��B��Ѧ��},�e��&�X�p��N�pƖ�Ү'��e�ȓR�~��f�1�4[��ۋ9
�ȓ#β��$�K�X�(�J傇�#�t��S��9�B�y�$�2A�R�,�tI��f/�5�P�6s�l�Ȕ��[���ȓW�z,+�,�1J���!� �Ox �ȓW�h	jQ&7~�0(��k�!J���Q�2�щN��X�)�,l�*Ʉȓ4�P#�A�=�X�s'*�� [X��`�Bl+�iq��a�q�ͨ3mh-��lw��{6�[/<�rY��EU0G��P��Ks�9�^�J�N�3���N1F(��z�dQH�Ɲ	c��Y�T@+	in=�ȓ54^Y��ҹc6�\�`�Y'�D �ȓ�Y����k��A�g�?)��ȓ8�BeSE>oN4y����;��A�ȓ2�|H�W�ބ>)�@���,gr���u�%���`b|cQĎ(W�~t���B]P#���f��i� ��$���S�? tA��BB�X�|Y�AH�|t>͸�"O�wc�7a|����%����"OV4т��?;�&yJ$�'6���"O���g��
<ջ�Λ>۴�	u"O��B#B�7��-��,Z-���G"Op���@��Ne$����	w\*Q"O|1􆓠�&$�@��w�"�q�"OTlK#Kq�D�i��Y,��=��"O�cPd
?P�X4��@��x�"O*����OL: �1\k&-1�"O�|���:ؚe[����U4�-�!�䄹g� �pFV�l9�ab��K!�$B�U8���g"A�,~,��v�S�!�DL 7!�iꤊL�p��"��*�!�$�#^0���K�w"\�j�	[!�$�6]!�E�a�d#�c]j!�$F�O�Y�ڡ5��eaVC?xb!�$��!_R��W������Ă�0J!��[�ٛ6'	^�F0�g$-!F!�O�o�
8�R넃"�V}aS�ҹ@�!�� �V`D��	9!�@Iz�#P"Q!�ߝ!��	�^,����(Ȓ@!�$A	!�(m�#�P�(�࢔�3h!�d�Zt%���c�"LPק,tK!�K:��K���ȴ�1g�7wA!�j�f���"f؂����Z�S0!�$qP�aWk_�[��!R��P!��� ��D��xC6XK�DƥWe!�9}�yJ�I:O�p�PD]#5�!�Č�<,�Uc"��A�C�J<!�D����	x�O;��6M6�!��-y�~)� ��.]�ɉ-ׯ+W!��2x<�KĪ�E������=?�!�\�^.؁31@
>NqJ��U�X�!�D�dnLS�D�aԠ8����K�!��$}`L؊⊁�"Ѕ
)R+-�!򄝫z'����(~����N�!�d�	 V�d��&���W���!�dYdh�۲��q��EK�F�<~!�D@17�*IFʄ"@���!��X�t1NAY�ft�t�`�)�36!�$Ѐs�*2�M�B=�A��2,��C�,s�~D�A��	t"�Ą��d�C��%8qJ����!�䤰�`�)LpB䉝@����� �i&�(�w���aEdB�	\�, 3�f�f~�̃�.[�	�*B�	W�މ*U�M(<�`@��8B�I>XM��6�˹}�`���-�6B��?J޸=���9u�6GD��B�Iy?Bl��,�q�4��Q�5ڮB䉧V"Z;�l$J� �X.��(�B�I�!d�-���i�čE(\��B䉼n�R�U$"�R&�8A��B�I*GH���e�?���C���^��B�	�9tZc�`j��(%��݊B�ɫZ�5��(R�+��{G�
�Q�rB�ɍ��İ��Yx}i��I>~C�ɔ
�tkfL�!'8~�C#IG�G]�C��	1�p@B�$���f7!��C����
�H�Yč��0Z1(C�	�$�00���K�B���g�l�DB�	�(�"<�q�w�t!VM�[�C�I�y��5�c	��/\�j��?	7�C�Ʌq��+t��0��ʀ�$M��C�)�  D� ,ƺ_����O߾"U���"OJA�P"�b6�J�n�0rSB@�"Ov=�,ω���"��9c����"O�Ƀg�K3�0��|��Rq"O�	q�!�`�P��kH�Y�"O4Cv��	����7h6�4��"O����G�ft�9��:/:)��"O�`###K1O�RCwo��,+h}+�"OZ��E��W�ndiu.Y�t�;�"Oj���ե$����T�֓ "�`e"O*K�E��W;VT���Ƈ1/�R2"O��;��X�d���
TER(1�"Ox����|a�dىK��Ș�"O��A�"����0s��kP��Z�"O���LD )|B���� jg�g"O��xc י&	�'Z�dL��'"Ot���`R�M�X�(v˩N:��[f"OdoH�AZ:���E�M�Ձ�"OʔB�&ϭFf�$0����G���C�"O^Q�ꖪ"�2D�@��v,�I"OF�äҫ@�=b�9
.8�"OUX�MM�0@��� S���bT"Of��C=m���;W
W�B!�T"O,Q���r5沅c�"��K�!�$^����q!�j�bI��.��TK!�䝤R�&�1 �I"ԁW�!򄊂I8��#��<�N��1��0!�՜4KP��.S (��՚#�N�O�!��΋���̓!olZ R���c�!�ĝ!�̛`��HhT�B� ҡ���L}��'O�h��ʝs�Fp�C�&1�5Q�'G�����2�8��"BM��V�	�'����*Z�F=��Z�%G�	�'A�#rg�$^��9�m�-PUj��'W���
+*H|�a�éI�J	Y�'A��ʢC\n���a��':8��	�'�������$1'>�����&�F��'�VA�F(u=��a��$#�:���'�  �f�<5u��0E�#�:���'�hI�򤑻!�>�{ dZ%|\���'�X�&k�c����CJ�bQ���'�@�0�Y������D���pc	�'�`�kc'\�T1���Q%� ���
	�'�����J��)��z��
.]��'�x��Mx���}�f��'�P�o�
�t ����p�Ĺy�'��=2��}�Zq)O�bT]�N�L�'*���O���k�AD�Y� ҂ 0p������y���;6}���4��k::�����I]X�Ԙ�Ƅ�M�h U�X ��]h��!D�d��.G;Q�8�� CF7lq�g?D��h���<u؈U��+T#{5����&;D���r�.��g��>����g4T���cA: ��Ҧ�<p��u�"Of�"! w�D�j!��3���"O(0(�!�,�i䫘�^l�Ýxr�)�SZ:��j����R�«8����'�D��FKƜ ���P2�ޔ�8��'��K���g q�Έ&yr���M>ь���P��H����Z:=�-b�Mg�!�č�\[<�iƨ�>�|��#�����(G��AE�gƁ�i6�8=3��ɦ�y�CԐC9�;1�䩪5!S�yB	ĕGeHEU$�
����d�;�y
� �8�7�V�6���HN��y��p��"O��wg R�X�F�A��`��5O �y�W'zD¬���.R30��FG�q�<�!�@L5�5f�pꈼs�m�h�<�׬���D��@7 X�z5&цȓ28.�20�ğNr�|�v(]�lsF��Dv ���F��6����lѪ*1b<���ְ�d��%��M)SIɧf4�ȓis�Ɂ�+�>&!LP���Y*�I�'�qO
"��N����72�°Y$��Q�<��/��0 IS��l���pc��u��,?�O<��% ±&�)�W�}h�9�`r�<��G	&G�0�ĨW�=���Z���k�<�A�L�3��e��A�	���Z��	e�<�3,1#x0M���ڒ	�e�S�h�<	e#
�dR�DN�rD`�#&�Bz�<����p��3m��&^"e;KL�<����DR�@�ejځhp�]G�<�cID0��`���h�E�A�<I��P^�d1�ѕ
��y#A�@�<� ��)E�Ё#"F,���Nq�<�D�8Uآe�Q��A5 E!u��m�<B��1֨�B�1#���؁Cf�<�q��$�6C�Gݴo�d�HQ�@e�<�W(̽S��J�g�*a�B%LE]�<i#�T<:ILq�?GŨ�����U�<� �
I؈��	E�n�huA�F�<IeCR<E���B)�7aT��aG�NG�<	U�	>����gL�3 (�`DE�<Y7��%W������e�B5�Jz�<ɗ �m�fu� ��vZ(Ec��A�<a5��+>��
 X��1E�RB�<�I��	f�J��L�`l S�'�y�<�B���C�*V�]C"q؃p�<I�`Վ2_� �'�ٮW��֣�o�<���ӓ/ɠ�YG#m,N��g!�o�<y���(�	��?O��]���@i�<��ɗ�$D�����7d�Z�y��a�<P� �"���A㉓6Zz�V��Y�<� .S&�6(JAg��H��X8�OX�<yph��8����ūuT��Ӥ	�P�<��@><..�� ��4��[Q��N�<�`��9Xl��+�87�����Hv�<�����Y��m��K�e:w�Rq�<AG�]-)m����S6~j�Lb�hJp�<���TZ�!��� �$��KE�<�b�
��Mhq�1r���pVj�z�<����G�j �⏉i�L��&A�<�a���x32���A{w�ȳ��|�<y`�
,�`�3G$¤����_�<q�b�M� E GV�Au�9QBh�`�<�GՃPd���Ě!*-��"d�<9�L'��8C���
Ț�@�%�w�<Q�G(!�a�P��?	0�)
��LZ�<aP��:h�]���<U�&=XDC�L�<I�̚8b#NX��kU4/
d�sL�]�<�T���!���w	�,S$J�e�<)��(a)Dt Td0{*�d2��c�<9�T+4g�1B'nX*V˞��bG�<!��С6��u��%M�T�;t���<Y�E	�,���7���z�*��W�]y�<Ѣ�/R@�2�J�y��mc.�_�<�Dl�/��A׏O��(��t�@Z�<�����0dȑ�ՒY�DB��|�<� ���4G�x��w�(��"O uCr�Q9#�T B����w8-jP"O�i��Jd��'`P�#��p�*O��u�8_�ͩ�L�	�Ru��'�<e"4!_:"l���×){�p<z�'!b)�T�N������X�zFp@�'f����FG�Cׄ�r�C5r?����'A2 ��ʞ%f����Ϯ�`Q�'�K��@A�V�W(�T�$�RM�<!�,`)�X	�B�*qPѮL�<10��,L.���	�m["�{qC�b�<���;Y֒�P ̘sSfiA'�_�<b�_�m�X� f�
V�L�Cj�E�<aT
S�e��IVC�q j�X�jUA�<!㗡b��a�Sn�Y�|(X��F�<Vi�#U� iy�IF�\�R�k% ]E�<�g^�慓�@�`�;�,5Y�>a�ȓg0X��T��l���{G�+j�4��;�>Q�UEѣ@����V�G.:��~/���B� @�+�f֋u��T�ȓ�| ��b ����Jċ!9ʑ�ȓx��eAp�NҴl9Mڞ<L�ȓR�>� �Z�e��d��Ċ�qu�Q��?f�*�W><́V��-n�D�ȓx�E�瘧W��18U%�x�e�ȓKKV�S`�T�bgH��&
�p�.��I�J�B�۩^+�t��3M(<�ȓJ�����B �w�z�ۢ�Cw�Ňȓ0�&Г$΂=�4�#�͈,(&��Z>0%r3�Щ`�dEÒ�S�MB�T�ȓI������,�.eڶKW��Δ�ȓ)�p�qpDG �	ZH@�],�,��}��9v$�,���VD�����ȓ; pIU?����f !R��P�ȓh�� ���ԛ&�"��f�@3W���ȓ`W&dr�>��eH���O��a�ȓi�� F$A;���'"� ���@J`�ע��H|0į /
�����8M�E�f���~�"6�L/6�~��ȓT��,���#�r���./3���4�,�Qm�3TKڐ�˛_��(�ȓg^���6�[4�8�J�(H�UP~	�ȓ!t�`b�_�:UJ�y1b	8ry�ȓbjA���F�-$rrث  R�<�A�Y��`����Z��u�F�<�V������ړx_4�[e(NA�<��O�	> �{&��6E;��C{�<iV�Q��j��O��(����x�<!2���SۈP�F��^
AZ"B�^�<	�k�xk�l��j�zq��W�<�眭E�,�9!�OuSF�h�V�<���%U�|ȑt�ņ`6,�-KS�<7G��V���6���g�Q�<� D0&���P� �ƌI�Md�<��̮
�-��M~{p$a���H�<aã,YR@����V����G�<����� sL1����>9x��GOm�<yGb�I��x5L0Q
�s�aKO�<�6I��Wf�0�e֨@z��K��K�<!$O]�8�dT�0!�<y��I��'�F�<YEl�gR�qj��8�'�w�<)�(U��P$��E Q��m�<)�,�B���!� �H���Rv��W�'w�(�D���		Nֿr�D$��'1H|�FgR=;:��S�X
x9Ʊ�
��� n����ĞhlH��0딇>��d03"Oj�0C�/	��̂��@8r��Cd"OH�ǂu�d�wB��ny��j0"O8�`#��v,D�&���Y{�%��"O����i�*ZFd�����Yȼ
�"O@�0 .A9�p�ZAa�VT�D��"OF�r4�#Y��Ͳ�aS�*�
���"OT��B�,GԮm�N�"�l=R"Oh�Ǣ�_�<E�R����"O`�S�G6�p-X���4.�T�"O4x��4���K�a�3��l��"O�;�&&��=#��>����"O\4�'���Nq0�!��Ɋ6"O �hD �J�5��Þ	e�Q��"ON�8˒
��[���!U���w�)D�@��튼a��5y"�/e�h�٣�:D��s���i%$��e〒�be�0�,D� ���|���b��`���<D��*d ;t
��O�Ԡ�J�#:D�8�j�{��x�GH��7��L�<D�`*��*&<05ӠÏ4c���<D�t�g�
P+zQ�JR�5�Ey$=D�@�Cg�*e¹��I�&�"�$;D�t��M�/,���G�T(Tu˦�'D��hPlS�\H�9�G�: ��L&�1D���"ӲR�4LdK�J��@�t�,D�P*���J��� Qʺ_T��P�/D�|'FGp#��ɂcD��.��I*D�(C�QR���g�"{�����(D��#�Gýr��)Í�O��pA�$D� ��팁	dXM��G�Ð(��E"D�t����:H�4h�%�K=.B�pC� D����ǈu ���7��v�PDP5�!D�l���[0p��BB�%�P����"D������`x�b�׼�DM@Ҍ D�D`�A��8��I�p-�\ ����>D����(
�qB��P�I�0�B��D�?D��!GkO�&��eӗ�S�=V=:��=D�����;w�x!��\�1X����8D�F�p���Ф�O��8���4D�����]����֏A���0D�T�c�#�ZՈ��-��,�� "|O,���+H����q����uc�
0���E�
%o!����L�S)Ή Zt�Ҥ��f��b[�hr.�)1�ËT�Dۀ��,-�	��T��5�aұ
l�}(W�ÿ�V4��BX��>����n.��BQ�BL�߀~�Xѡ�(�f,�Ad�4R���g��Op�@�O��Fx�����c���l4��V��HOZp`%h��9���6�E�eV�*ܘ��� Z���7��?-�P��Ə	|��.A�ł���I6$�佃ƅ��N����+��( T6M��tجx��5�?�Pŀ�iB�KG�k��XB�]Z-0X)�2�}X�F�gj���j���i�|�JR����I�V^f��$��,�>AkF��k'��@�%GH�A��o�c �ن"�U[b��$IQ)��v��>�J���=|l�RA����'�f����F؞,K��W6[/j��0 �Wm:����j\z�2%�-z0U�8^x��EW�m����A��p�+��ܴ䂝']�n9W�F��1ȃ�a�&�j�ͶjG��\�Ν�Q/H�0��'�@)Y�Z�&�±z��᎑�p�PM��1���X��jTk�Ι�	zQ�4iأy����4j�5sc�O��,[���~BN\
_g^��UIՄJ���'`�M[�+�)1�>��I�O <R����¬R[w�"@rd�^?�@b�4Z�4�cB�n�`s�D?i����) ��MBA��n����W�{�4	H��d��pU����3P���1V˝�#s!#7E?OE�!3��Ka���b�qӤ\�W�I�f�}��vӂ�$,]�&��$+��=\���Q!�.z�)�(
�p3�݇�I.p��hJ�|Ni#&H��6-C`�B���G�Đ7a�(��,�0 @*p�$~@$!�&ɱy�2%{0db��m�%C�9.)�� %�W0���É��	��yA)O�9�$m��ڃC
�v+��J b����5�L=:��Y�B9E9�4"눹^��6�?ɘb��'�v��1��Q#P&�̠!�)ܐ�)��'e��#���^�8����6� uHW$S�	`�͙���Jܢy�+�qI*����ڞZ�0���� d�P�טw���+f���[X*���	
�t�AOȽc��T��E�ZP��O�8N$�c�BC6Vhčx���R1�q�c��=.6��
!=�H���f_$}r��%8E���^����)�
}�.�r�rN���%oα+�4��g[>1�G��Gr�M�d��J�K�$8�f��A�h�<i0�ؒ'Ú��	4,�a���W�@.��B͸�`��$c� E�	��!Č+�*]�5���yޭ"�d["{���BOڌn���YU/�O�-��A=.�����{�\a�m�}�㛯jqR�s
��kL�"க�=��y�G0X����T��\�R�#؞b�b4�U�ЋIB�2��I�u�X D�>Bw"�kBGՍ=��I�`K�QG���¾%pT���	_Цiည	3z��PЗDN+|$�{΀�g��	�⛢�h`�ɸ-�:]+F@�#(�!	�%�����bp��ʋ��n5�6��
V���������i�vӢ	I�jQ�_�,�!U<�zr�ۓ��6��ǿK���^"��9�H�1T���!P�Y�'G�8��GK,f����[�� H�č#=r��:�R8�$Xj��ע#�|�u��,B{*���샥q�b:�.@��?)��R:�0xZ�)W# �d�U�x���"v�]�Z~�!C��?Ǜ���s�m�ܟ������&&�}I׼�,���4:��)���bAN\S�EJ������+$FdIi�d�@����(x��z�֕dEJXF}B�T)(�nU�VLT�/��p��8X�D�Ҳm�i�ZM�1�����	()�jU�,U����"�"s�"�U%T�J9�F���$.4Y���Q<lKx5`E����<��Q>iAlP.ؾ�QK�$6&8:���.KL�݋���5FF�0㠂��M�5I��|&��� ȉePX�'K��N�y�5�Ю新�a�Z8������ ?ۖlxG�'J�]���,�ȣ�5GF�h����Y��p�)��'�$�a���B𠴐�k���I*��Mq�	��O���E�~�X�g�_=O3r�8#ZN ���O�q���&	}�����]�����'�y���,^p�:Cj�8�L(e����8�H u�/,O�@%��?uʀ$�&�� �#�i� ��a�G�O�LSЄӑbzn��ڟ �	S�\c�uH���6df<�Q@	�EgZEQ�'�&)E$ǒh|�)Q$IÃ@T$��%.��SFp��F��'n�e+�嘆P�.}�OR$=��h�	�'�BВ��Jh�ap 
�=�-p�'H�ak"%�B���,� 0$�0�'o,qaᤉ�Sͪ�� �:����'�\0�B��]�������x3LP��'�t�w�܅?�؅JUҳp�p�Y�'	hh���o�
Ƀu(\�k>4{�'!n�2��V��A:�ό1Έ��'�8IqDM� Wt��0�"9����'	V����TB�$<�$MƲ?��{�'�$�����AJ�$���X�n�j�'�`��uٸA*BN�l�&�r�'F
�"��Ӂ#��%Qu��J�vE��'d�t��j	P �55MBEp
�'�XSUh�'a�,I���3s��K	�'c}C7d�7r�B9B�!ҍu~�MQ�'�\�A�F.��h�#� t�P��'U���� 0)�4�£_�u�X��
�'���
��-.���d��d8
�'p��+W[�B=Wo��Z�:��;�@q���K&Ds��ɫx<���;B�,Pg�քZm��b.�%+���ȓP>y�5�\�<@��g �(U���ȓv:�TW�Z�^Z�<�# �)�8��ȓ/���XN��I�H!����^켄�^�(���-Ah����ӣ}���ȓ"~�9�@4�b�bZ	0,�� 爜����+xu:U�GcT�(�ȓX��aP���yNX��i�l��ȓ<�q/�4�Tbj�<�\�ȓ,��C1,P
?jl2�+E��lL��i���	�уC���!���gxA�� d.,��f@
`��DAs������0�z	aV�+<@��.��V�b��ȓg���j�	�-�a�OB�Y�)��<��bG�->D�edG�>ڄ��7�&ș�#3H�$���H(	(�M��b��� B�3�PMK`�Q�����ȓX�dPZ�X�=�
�l�䉄�%�>,�r'�E��J�K�)�� ��S�? ���V��R���Tkٴc�<\�4"O�;t��y��uq&�D�%¼�C"O,}iV�8qH�@�p��/�(�"O������M��J
*PhlȖ"Oͨ�"�u��`��'L�J��"O�� ��=���Ɖ{ u"O�k�&j-RtW.pZ\��"O估geY�U9�})C�1����"O�8�π*��Hn�* �	�"O�Öʀ!~JnX��-IF��h�"O4�{5e�9e5j�g�٪]��p�1"OzŨƃU�oF�UѴo]-Yh���"O.�S�Ğ�=4P�(�1rH2�3�"O:A�A\�<���CF 0jH��"O(�x]
!4J��2e��[�H��"O���5�ɝB��� ��>�x5`g"O6��-��#�HQ�F	ܚyk�"O�I�S4!���(�W���Q�7"Op�q n̎Bz4a5�ʕ'����"O�L�%�ΩU��-�aˎ*��h*F"Ox��T愘�Z�B#�[�[��@�"Ob	+G
�?*�(�c|W���"O���f��!`Yx��f�ǹh�H�v"OzE�(F�RЅi� G�LH(�"OJ�`E��$Y��툄��H�93"O�l�ԩ��h�:�s��:q�~(�f"O�`�WL�V��<x��5<��)!"O�Q��= ]>!��Y�%�� `1"O��Csˁ�T(����.��9�"O.Ȑu"�k�<m�P�U�!�r��"Oz�8��¶,(����L���I�7"O�iP�
V�6d�؄퀈��4"OH�(tG��
�T\��L�,"ߴ��r"Ot�9f�lU��z���"O��J"O�Y+1퐾9��t�2�H�J�hr"O�9)g��4�bѺWM�*9�hq��"Odl i�"���t��R��dHv"O~�{���h��0�� ��%6�"d"OF�@6�	�8Ό`���A+*8#�"O�T'!���qG�"� �@"OPAR��P��d��m�!p���"O��0�֎wmHs���;��S�"O��JY_�T5�E��)J|!�T"O�H3%
�L���� ��  �"O�M(qnY�D�L��lV�S��9�"O���M.p�Pcr+ƣuΎ�k"Ov�JB-��G�1G���r�"O�TSץ't��a��[���"O�9�w �.yMJ��t�P�gP+"O�I 7�<a"�@�Zfp� "Op��m�^��k�I
;&���C�"O<���B6M���A��@S�@AP"Of��!�E�ym�D�2�
�T[�]J�"O6������fH�AΙ^�)ؑ"O�҃(�?r���S�V>j)� s"O���KA�r����	�.	8 "Ol(@��,K�����&S;P���"O�u0u�1
i�4!��͢zH�	�"O�w`���
�a��"?Ht"O����P�V^�Q��I;A��Y�"Ol�y���;r A ��X\X��"O��w̏>m	�E��06��,�C"OR�sҪ��TRB�[F&̾�YJ6"O��A�[�r0>M¤�3:�v�I�"O� �ѳcA��n�.d�'�.G����"O��'X��j���Ӵhھ@0"OfZwf�*L��V�� �"؉1"O�pb1��#�J�c��P��"O������f�ȴ�4�\�n���(�"O��b�A�P�Qj�n�L����"On�؇`�#/5R��1˾c� �)R"O����(ſ"��xW)ٷQ�fPC�"O�msU��=Ѿ̫ӈˁs�1I"O�p� 9~���4��#m��8	�"O"<p�^5������ߑ�VD��"O4�p�B�H'�=��kGAp����"O$��`�Q�TbQ1"d��E�*�1�"O�Y�fPb����c^�k� œ�"Oia�Jߡp�~���!Ŭr�
y`"O�Pȅ�=hyL��1O������"O�Y ����'��d@&�^U��"On��S7���G,J��$��"OX5���iu� b��"+L(�"Oꅓ�	[5���˂�͢N~u1�"OT��P�R�;K�u�� \-$p��D"O�]�r�	�K*0t­�S�H	Q"OF��H���zIb�6tS<f"Ojd�4	Ӈ�0�⡒
_����"Oд��e�]�*x�-�y<( "O� `&A��D�,��4fE�^�1"O�h�嬏;80���T?Ze{�"O�I��':��8�At�L��"O��0��ݿ}`���ҟ/Q xE"Onuq��iց*� �seh�e"O�)�֪���E@MFt�ɑ"O��;�E��-�4Qp�Ţ[4TM�E"O�v�9�n��I�#>܀�r"O��;�F�(�BX0q�.?�X@�"O`8���H�cч�Zǐt!"O A	�	��<�����޿x���i�"O&]���JLf,����ʭ�e"OJX3��H�"9��Z���<a ���"O��a+�:W�TPȣ��Y[F"Ob{��_,�Z�����K�h�B"O:=�'$ݳ=i�S�!���8R"O��d�	�d���FMXj���r�"O��[cHյDF� E�)�\�$"OL��#D�,M֡�p睿a�n9+"On4p�
X�����B�(�j�"Oh$YS` X��� ��g������'!�ii���X}"�=B*DA�$ŗl�0y�!�:�yr1��Pjֽ��-ʛ�M+&��+�@Ū�V4C@�QQ#f�����O��6H�Z].ɢ �M?~nD1R�Mx�!��b�@�(�J��;�"DZ@�Z�׈T ,َ�����-%q���`�'�����o*#<qĢ�'Z%�mK�e�+B��qgK�'"\,R!Ӭò��I!h�~ĀCB�"�>�[�E���8 �N�$�Jt�U�ٽ[-q��� &����B���ȣ�-�]i�h�"Fڛ�C�}���ԫ�ݟ̈�CZ�Q3L��g��,�r��B�;����wn�T�Ea� E����r%Z�j����'��ЦK�d~İc�%E��R�s��K h�59槍8PPB�Q��8Q�����Ѝ ���C��󮉕~ӴU��c��nQ�+э�a}"9���NG��S��C\��q�Ԣl��쀴�<�,T�NܗC=���ژ���b��ȝ�R�'}Ҏ��a�N�+�i�8�Рx�둻�HO�qQgKֳd-����Gm^��5H�u�x4o	b:�x�2'N����v/S%@�~�`c*u�PȇG�l�6Q��I#D��!���,�2�7�� ��7�)u4���e^�?�S@׸C:0�R�j�a�ǁT9���ծp�P�����EȤ�R�gxPؖ��<hjB��>3��A�Ǝ<��x��1z��#���h�����N6:K��������Cb�~;�m�}���w�x�K����N,�����:J�y�:H�m+�
>04��YR#���B���.�# �(0R�)9��-\ƕ�������	({�X�Bޟ�� :��J��f�p���L#qp�V�	��R��\��K���3�T�]�!�hd�ehG*�����/���ISa�%���FYax�%,��`�â�i�4"�M���p?��hO����m�>�$@��lǔ�l	цj�+��C�����(9w���I��j�`���>�Ѫ
p`�I�`�1�5K��p��X��հa�Ƭu- B��77zq*QjÛS2Z�� E�m��ɉPδ�qBѴ+�S�Oڂ�����N3D��ɦ���;��d�]"�Z+O4���,^��zv�W��퀐̓�O[�8# o�d٦��4C���0<1��ߑB�Ν9T��<��b
�9L�A>���+R0�o�!��tG�z�P���-yK��q�_� h�8��C�N��Q����5!���6Vh����=[��T��_���eK�F��[�����������޼���z�F7m�0�λ\��QH0e�?�Bȋ���%I����	\M��K3�W<�6h뷄S�,�p�&$�z�t�(%�C7}O:ݨ�iژ��a�׮���)	�3L��H����>�~=1�A� hר!�E��,3z#=����W����p!�O�d���j���Ț)V�Y�&��ؒt(���.����%�o� ����!����i�0�bg& h�p���!eD,)��p��x�$��ĐL+�d�|1�EO�O�3%�C�	X6^�X��E7P}�a���'(;�-�"'ȍ]~R|�'�y���	g+�J&���mzN���a_�x� ����b�z �&gվ	�m�7˓�d.�(nڏ&���9���1'��{V�R%��'��:G�'>.��Ο�x5��A�=���q���Bc�86�6)�@.<���!��%T��F'���g�W�'>������n����4b��n�ΰ����V�iR��߷�?�k�6t`V�!e^'V�^PX�f��6�m�S,׷o��@a5o��A`��)S�YF��y׭��7�4�q�J%<��r�%�O��!����ɓ.�ܨÖ� �?ɨ5e�Q�-�>�qQG��
3vX���D�Vk���V"O4̺\�8j�"]*>1&y�fH7+��fI>F�^�[�gF$NѨ�6嗇X��	��@��5�@�h��Mq�ׁaOL��g�'�y2K�1��A��+2C7�ۍ1��QA1#+�X��~�,H	FY\|�G��-��<�b���y�AċQ9|qz!J)g�a�@��y҃D�%�LibL�4SR��Do�
�y/�N5ʡ���H�g>)s$V�y�5��cri�tI�C,��yb��#@L�$����b�i�-�y����v�𸤅��J(*�
�yb�WE��P;��ش{Z�Ac�ֿ�y"�Çp��9`��J�h�������yBnY7hs\哵K�f�<Y�@�A��y"�՛q�-`քE-��eX�C��yb�� ��%�f
�0�0��J��y��o~�=��I�.'>���y��̻q����!��!"S�;�y"��7yHL�4��	�HTscV�y2g7:y��9��
�;�B�c��)�y�	�
��I�s��<�0�XWfW/�y���5��`W�+�UX��1�yb�g�Y�ț._�0���=�y2�Ż7҈�U!�M̰��!�y"#ɋdRXh��8F�� �R�yҌԇz���Y��(�"���%�yRCS3)�pQ�k�0'�T ��2�yҤ��V���,i� ��gaQ��y£��S.̰�(څoT�Q�7����y�N��ٱ`�΢dOJpI���	�y�Œ^ݠ�ˆ B)D�͛�ND��yB��;��u�QB6~�0 fe��y��]W|xRQo�T��F,�$�yr�ȵ	��,E.�L(��a� @��yr̮p[�R�-08D�r(�[�<t
0���V%�z쫆.
M�<�¬��`��!Y���k�,�/E�<y⦒�	�(]pSa����^�<����B��EP����Z�����$@U�<����F��q�Vh��m�tXbOS�<� ���ÏB$!6��kcg ��"O�4��p�9ږ�F�Q�Vt�"O���uN��,N�	*����ɪD"Ō:�G�1%�$�E�!z����"O��H�ټ�-y��#��$:�"O�y��Ä`yB�����^D�"O���1\��؃A!�?Z9;�"O��y�)�cP=yo�eԑ"O~( ��ɶ��P�H
@�8�"O���dN0&֌(1�Lb��:$"O�=!ˍ
iZi�a�WR^^)��"Oz`�ڤZ�l�P'I�tep��"O6�cC���&u���h�t�/*D��wo»#"��	u-��P5*O�r�Q)D� A�娕�=9��u"O�Eis 	$(�Qb���c����f"OL�+` �$�V|I�_�(��a"O�YjQ@�%|�<r��.�nP"O:�5b/u��#�0~n:` Q"OH�:Sb�)Sc�0Z͊�U`�(�#"O����Q!���t��.e� zv"OHI	r���� U�R)X1rHr�;�"ON���'!x��#HͮxP��#"O�B���t��ѷf
='����0"Ov0��	�	�X�s�N$h�v��"O2�&	�)Wq��Ô"q�^�zW"O�u�3�L&GİS�Yn��Y�c"O���r�_�#BrAz���8{
��T"On,`��T���8�H�h���*�"O �!�l�P�t9 żC��<�"O�5�2Ɋ+5�����^�\a �"O��j֨T`�)��읍l��u+�"O����Xߜ�(�JJ $��*�"O��x�NX�&Ƚr�H� c�~Pi�"O��	������s��,{��HB"O<1�'LY j_,Qh�L- ��TW"O��	1D��j9a�Nԝ]LV���"Odh �\y+�X��2u *�"Oz0�T�@�8���aK��[�N�Z�"O���d�5U��bE(ԖT? r�"Oj�Z@/Y�%V�RG~!��"O��a�8^���/�E7(w"O A�f�H�q���nP! �<`�q"Oڥ`��9.-�D��s<=+ "O�p�ىN��dlA���$"O�(��W��.M�R�e�<��"O�M��f֪Z�eB��y�Y��"O(1�cI�54�.0c��4Wtq��"O>����;[�~����]�N��"Oj�bFa�>*�(���	� &H#"On%�dH?�q�4�H�d�%"O�9�֚jd$p$��9q���k�"Ob�(�AyH� @Ƅ-�l��"O�,�(�}L�q`�� ��� �"O�5H#���2Ԍ{'!O�>�3"O��s&���Y� _m�$(	r"O�I���* �(��B���I�"O��x�E<K�r��1�ݡT���t"O4�R�ïr�n8� n��6Ą@ye"Ov �R���f0�(7�ס8�p��"OZ!`ǻ����cKt�F��"O>�z0KҼgj<��➧(jC"OH���e�-g2��B��3�P��"O>Ź���
zp�@b� �+3�p��"O� <���c��BD5��[��Ti3"O
��wG��.���f��VG�I�"OPP2��p���)�L���kP"O�m�sfM�CTД�FIղ���"Oj������|�����/�.��1Q"O��c��E`��h��$y��Q@t8O>=!�
rq�/�C���6ΓS�	��uc7L�2/ҙ�`ƛ�|���pL�7�(�J<�7��4o/�)��S9Z�irb�Aı�`�Өj���@� �k���'Qԉ��UH���$hM���V��3X- [�P@�∤hL���F�]D}
ç9n��������Y��F�*V����V)�"]�<��ӏo�ZԠ���%`��z�(��
0���v�%��-
1���)�C�@ҡl�	0L�6��Ik1O2H�&㐜Ija�d*�">.��H6 �t��QIO���$њl��H���Ӵ	|!�Ս��<��%ɢ��\��I�^�j|�c�<�)�'Xl��v-G�|0H{5�1^�4Y�զ��m�p0�<��S�04�x��;����Da�S#�B�8�c}��V�~�'���ɟP���!�dA{`�K4�]#�Au}2+�� B$\�A�Z���	�)M0Ȑ/O2f��PB����B�	�>=R��	�65���L��HH�B�	%b�yZ�< \����� ?i2C�ɡ3X����%)�mȜ��W���yb���(
�fW�^~P�bG�ת�y"+ЃeL�v%�Zp������Ms�'
J`���&�Lc��
��&A��'?�$��ݥp�f�rǂ�:2v���'X���4�G��
&���B�'$<|kp�­�ɢf醚0�<"�'��y�TE�12R��.��$�9
�'�ԉ�3�� T�|<[��t��t��'�dbMUn�ؓ&};�Z�
�'m�� �MZ6s^�r�(C����'O85p��
$+�ٱ��[@j^�*�'��q�ȋS�����9B�9a
�'���0Ƈ�H��s�$?~�Z
�'�J���%`�D8c�"9�E;	�'�@��D�:��B�f�,"s�9	�'e`���M����C%L��Ĵ��' L��Q-�"F4dr����8� ��'^�b�D�Q�	_: �%K�'%������/��D Uϔ�~�du��'�Α1���_!V��DBN�j�Q
�'��ěS��$[:*�)gG$1\�9	�'F�A����! ���5bW#.¹��'��x�e]�2��%&�x�	�'� P;ǒ�Zl��r�ܨhd�1q
�'�nQ�Fm�f����*�;\� �
�'~p���
I�_<>q/��M(��	�'�ppq�*$��Y�d�C��@	�'��L8�耮IIF\S4�G�B�1�'��1��a@@�B�S�ؙ#m*!a
�'^La��h�4*�Ne!�GQ=i*q��'�HTk�.H�2�0}j�*��m:1�	�'=f�h$
K�1_R�b�'bjj�#	�'���v��.o�PYC��X�l���'Ͱ���d�-1Y��{3����<��'���2�(|S��s��>�9��'<VD3cI�0N��z#�+M���'�J1@aŃ`
�Hj`� W���'��D����s�2�`q�TO6d�'!����,�F0����J��	 �'��\���D@��C�E���
�'���%E�o�h�S毅�K�m��'E���bk��w�4!#�*F� RQ	�'�F�3�T}w^����5������ L��h� �|\�����Z@�S"O��I�ʑ�~�Ρ'��t�d��"O������ĹڕKU9w&iR�"O"�J�DC�0��JK
P��"Oft��MG�3�am�����(c"O�񑴱J��sO:tJ�!�INe�<��-�e��3�@�r-R���C`�<1�냮��ܫף�s�4�GTE�<��o
=�n��ć�n�<��K�F�<Q0�V5_��|Y����@�!�K�<�����Ds\Z�cZ=N�4x�S�F�<����Q�(��	�;Ca�\C�@�<�7�ˬ �8�U�V0HH.�!P�S�<�A�dʸx{�`�5x0	wB�N�<AB�^#�L����_�H�MM�<�-E \����#T�;��Pr�jJ�<A@��q*�L`U�'�2�+G�<�@���?OT@�����^<�"WC�<���B�xb��ػgCd���NX�<��V�bK�5 fC̷c�8@F�K�<��,�6ᚈz���4r�`�10�XF�<�ĩ4�.��˂0��)�!�\�<��J�CnACѪX6��hR�@�<IϢUfJ�`c(�{�s��|�<W/�.q^T����L�f��R�K@�<	��E
~Xa��n��T�l�A��r�<ٷ�1?��4�U�a�X���I�<�o_J&|�(���3E��$YĐG�<�U�7ԑʶR3V�z��7�m�<�႓�Yٞ���2bĢI��a�<�SV�#V��0l��޴s���Q�<�v�K������,/*�E�i�<Y&K��>��Pz�����0�o f�<����K��4c�$F"-�:��V�^^�<i%
%+�@A؀b� fJ���g�@�<FN�>e��A���P!fqsU��@�<�B��#��K%����Pv��f!�ƹUxh�1s ��y��0�P�0"_!��
�,̊wȐR���E��"LD!򤇪7�~]�lK!)�������F!�� )hT�抎)`��G��\6!�$�Aۊ�Amͤ\Q��x�+ö&!�DT-����2B�R �8*!򤕿Ig�h���	�pǻ=�!�D:a��5�Ɉ�c�=�G�
�&�!򄕼;FX�%!�B��Q�L�(�!�B�M�8��Ć�4o���	"��2F�!�B|���SA�Ƴgx����عK~!�d�#eM(���CQn0��f��P�!�D����p$�*Pzl�0$X!�!��M�d
h=S�ڬ
:x�:Q��\!�D�/����'�@?;���#5B�!�d^�v�i(p(
�yЩ�gI�{�!�I�.'jIc��'gi ��`0F�!�dX0(bu���>t��JP�˂:�!�d͈]��4�'	�J�l�v��P�!�d��z�+���:,���N %�!��I1JT$y���FFT=��ē�#�!�$�)]*`�C��ܰa>�M�T�S�s�!�O3t9�b��vQ�vD�L�!�$3RL�p;7h�����W-cc!�dI�ּ�q��
d�|�rQ"�
c!�$@FX��s��e��� P�5Q!�D��3�`�#��C�k3��%k�!�� �(��HWJ`A��P4D���"Oޠ���*H��Ѩ��� F�˦"O�!���Ǝ9/�m�	��enx)��"O,��f��'b0��J�nRD"O|S �����⢇"@��QY�"O��u�bk�V<C�@]+2?�]��"O8E��-�`1��ȥŉ*N��{V"O���el��d*ܚnNa
�"ONM#P�V�(3�x!vKL1�X��"O|HPcN��1�l��
�Lr��)�"OhA+B��$<����� hZ��!�"Ox��EԤmt��"���@���"O`$``��	s��`r��
1<2 �"O�|�c��fN�q�NR%���9D�8�i��Yƀ��bHir�J�8D��#���"��Ep#B�'!��`��6D���f酶~�<��ԅ�2����B�6D�8Z�M�W����C�,��a���5D�x2�(J�M	�t��OD-�	Y�e!D��sq�W#��x�D��t�8�R�*>D���dێR}�PxC���M(��&2D���b�tXq3�ʻa�dYX%�.D�Xʥ��T|MJA���b!`�pT1D���'/�,��
;h��U�"D���#D�zv m(�薰e���C��$D�X	�ၧAeXl�4U�JĞP�C@$D���ѷ	��� f
��e�|�R�A'D����@�tlv�k@��]�H�D9D��86A\ -t��EoOE>|�;��4D���t牀*kX�ADD�VJtt`�.D�i�N��8�.Iy6��4�12��?D��"��_,k*���qFF�a =D�P���
�(�Ks�L5K�,m�� D���R'VL��6N�"�Q6N"D��Qdb��,n>@�.�m���+j>D�X�@����Td�ѧΎXW�����=D��s���1�*U���+�B�q�?D�
�-��$� �רC�0,���;D�h��F�:3j�A�N
hL��5�$D� p��֒0�20Ju�GAN��rq'"D�����v��Bt��?*8j���?D�x�ƫC$&�@A�cb\c� D����2E�n$�ѵal����>D�`b����{Q��提�T�q�9D�����ߝFr.�����5}���pn6D��;����rQ����l�r��*6D�ر蔬]�j�ӱ�Ci��P�0D�@XVN��D��l���=TZ���l/D��#
-,u�q��m�38Z��!D����oG�h��QIV��))g��8C�$D��rG�/���3�#W�Ē��$D��Y֦ 4�
CRE�%l�,��p�$D�lj ������#OK.m���H>D�P�S�4�<����EU�a�s�9D���4#�1s�d`e�u4����&7D��+%��.�>�1�0-��0A
)D�����:%[2!�c)b���#��1D��A0��)4U
�Pw��=��3�#D��`',P?����e�ݧq��T���!D��`n��\���H�f&l��K D������%�d�v#��$�ݛ�(=D�L�eS<2���X�����A�$<D�(�p�'��Qr ��1�e�$D��;�K�5Z����v��qV`;� $D�� ��YD��ЙG�ʐ(�*5�"O���&���(���>7՜ȩ�"O���6� �T$�Փ����zä<Y6"O�xC�C�9nݫ�i�++���RA"OrԊ����	������c��$Q"O�����I�D�`dP��J=^<a#"O`9R �X�$� U�t��<S�M�"O6	�c�V�iO8����:'(��"O|q�`�  ��hBU!J�e��Ec"O�ؑ�N$4H�����c!BG�\�!���S��C�(�W~(�1��tv!�����A�F��h��ss�[�x�!���L�W���fV"�	�'B`�!�"s�l����d�v�1�f�xD!���5I �Ȓ�C�k�E�X9!���^z�S�9V�p	Cce��C7!� uz�����X���Sj8@(!�ĉ�^�\̘7i�7�F� @�ܫz!�0^��"v�Ҳ.(BWa�a�!�ُ>�*e��b�q蠴SաѠi�!�C*�� ��K�00E��h�* o�!򤊰��2G�<�ظ�'J�%I�!�DG�\���C`�O��%�NY.bg!���7�d]��)�>{�c�.Z�\�!�D7;���_�K]*I��M�*E!�D��X2ʹY�ꚓa�8��u�C@!���5M�NY�`�#��� ŋUM!�d �Ls���CI�-�V�2��ìM2!��L8o���ڵ..�T(���8-!�DF#X����2��-�Г®�*[%!�$�-�^ �ꐅA���,��7!��]c0X8���#���R	8>!�$\��(�IR/	�x/�V�B<�!�S	lxs"Ǐ*��}�l+N�!�^�u��ܪ���*f�J8�vEǙ8�!�$��c `  ��     �  -  �  -+  �6  NA  K  U  �\  �h  �t  {  u�  �  3�  v�  ��  ��  >�  ��  ĳ  �  J�  ��  ��  �  P�  ��  ��  �  ��  S _ m �+ 7 J? �E �K �N  Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�� |d��"O
`�(�;���8���-0��1%"Oj4��ND^[��"3/9�0|H�"OB���H��*�ʞRy=a"O�味V�!X��!&F�:J�$���"O,��a
���C�Ą�M�"O,$3%o�-���p���+Ն�:1"O��ݢ1����`���y14]2��i�<�6��{_���c�H�`�fX�$Kn�<��A̼VI�xR[�)�Ć�pඤ�ȓA5��('nߡ4�� �)˩%� ���,��r�؊b#`T�eT09���ȓ!�b��g��}�8�F��-? �ȓ
K|m�ș�VṔ���2�%�ȓ"R�X�j�4JN�1�˘X�i����̹	_�jZ��1!g��zܶ��ȓgil,*�J�
j�Ne��i�J%b���f	�(U��:���G��$Y^م�~r�� S�%T"���k\�jx�ȓ|4�1�îJb��@ӵ�ݩn�V��/[`�"�v4�R�!ʎ<��M�ȓ`:��z�ؚh�J�Z��$HY:	��H��p�m�C1��!��B:��0��EnjZA V;9����J[
2���	��4'J�EA�IVW&��~�(aZ��ӹ�>� o�Y�|�ȓ�f�A�
Ο7�H��M�$�����mޠP����/���ANXo*�ȓTv�����{ ��-7�*h��I��sB�8�8���3����ȓNe*M�悡;������X�o��!�ȓ'lj�#F�m�+R&;�|��2)n�C��0S4���T:
b���:�0!��e֊��)��ͷV��,�ȓ0�&�8#���� ع�L�����;�P�AFd���,w�6d��r�EQ�( �gVlɦ�M,H��,DP���|�I	$G#\���ȓ"�)���E�B	yt&B�^�LɅ�4�� ��eëF�ڙ��n��R�p�ȓp`@}bŇ�=�$�AUN��P����L��p���_�a�)�Y�!��-��u�5���o}�`iF�@A�p ��F�\�0��[���IF/5���k>bTؖ�;K'DT`�^��@��fnV���Y�b�lI��	����ȓ,nٛ��Ć3���kC��8�m�ȓ'� I ���x<=���޳{��	��6��(� N�����
�y2<��ȓx;6q��I�
=  yG�O�,�!�ȓW�>���.؜ɰB��;�����`9"�ˁl�$@��- G��Dm�U������H:�\#�*�i��BW���y�H�{��Z��P�Q����E���=�O�ܩv�ټH�T�B����.�(��'I,#=��"�R��ǣr���@@i-Ȕ��G!DY!�W� XJ03`aDj'n����:F�O��	��M���� ���9w�V��ȉ���?!�d�?]�J�N�<\��a[��	s1���|�.�J?E��4&��􊰢	G���g�P02�ȓm�hk� S=PH����;�bu���'�0�3�y��I ɲ�S᭏�B�	Q�f]�e�����!?� ����QC,�����i�"�ӣ�'F!��߄WH�'戒q��gh޵㑞+��S0#Q&��7,�)7 PP�͚>9g�C�ɥX�`�А ��P���c�ڰ} �B����kU2.�<��K��0B�	����;��_�Q|�����Z�b�f�I@؟�2�FF��	w%�I!�(jn$?����S�<�.�E�B�71x��VM�=�DB��b��4�f͛�f�PyS�D^��0b�h���<q�.ޜM����!�� mf�+ւ�C���Q��xr� r�F$ cr����X=:]ذ��lF{��tk��33��E�҉;�8a�6��0<��40F(b�DS�	�0XBَD�KN>D����E��$�����%���*O*;�B�A);Tl!���"O �Q�Ѿ/�&Y+��DB
�%R�'ޑ�p;�B�G�j����܉k��X@*O6�i��L�9��h�G�mE<��!"O�����37�$�0���p<�`�a"O��3��	"���@�T2�%1�"O�4h�I�X/P|�ե�@��`p�"O�Mp�lB�J�NȈQήL�!"O�q�Χ)�z���Ѫ��1�D"O�[2iF�>��e�Ҫ�!AƄ�ђ"O������mq x S��;��H�F�'�ўxbC7:v��D�Q�P<#e+D�xyG�B'���[�ϳ@�4���=�	٦���I��Y��$��īu�3��B䉙l6� �ڮO�Y o�
9|*C䉐H!�x0�]�?t32���B�	�Dl37ᚭ\:��h�<��B�
dߴɻSmi�ޜB�%�v%|C䉄B�N�ZBC�Tr�����#�xC�ɺ;(�x'�[Ȑ��&��'c5vC�ə8<���a�nD��JU0O�N˓�hOQ>�X�x���E� �"���l4D�8�e�%��əٯ
�Q�֭=�D5�	��Q��mq�h!)�MYJ��t-Y'YA@$�2�<D�(��mφLe��9�ËYJ2��&�:��Ig�OK�5�"I"�Z	xr�ѵtbU��'�(��0n�6X㒁x�$�A���'�pm�U��6.�E!�MP��6z
�\�Υ@,O��1�cڊs���`C�2���C"Oh�Rc�A9' 5(Eo��+&Z�A�"Oȩ�UE�!j����ҭ< X8q�"O��C�S��PY�d#Q1M����!"O؀�럢B|��0���8XZm����w�O��`
f��']H��`�IT&�Ҋ}��)�)\<Y� �aD�[�d��굉йYF!��_G~�]���5_ՠ�I�g�=6!�D׎{����g�$�ȅ!&m�&;5!�@���$s��Θ<�R��D��@�!�Ĕ�T%��a)�+Qo2h�3��=M�!�䍍Q��0�.�/9S�yx���!�6�.�T�J<�]�vƋ�D�!��8�`���<: $����;�!����
�Q�&]6G�lt ��J�~�!�d�8��7����"pa�#l���N��P��J�t0�!A�A o�\�:qN-�OJ��ܨ;�ԅ]mBxhG�J�o�5��Z��
Tӌd�����@�dܔ��)����a(��9�\Yp�#Y�`�(����]�Wm��	/P�[�W�4n���xpi��G�F2�0+�/?;lE��S�? �� ���F�l��VC��V�t9�V"O����O�
g`D��>H�N�3"Oxh�2�G-9� ��&��m+��2"OU�2#����+��t�x���'D�X(̛�OE����ܚ9-�l!�$D��C,3A�M�FΛ�*;�����.D�@a�IEeJ4�ZAZ�r^�((@
+�I ]�azr)^�>��!a���b���������x�+�+�*��k�v0�Q�	��}6���ē7��͓��?im�y+Ǚ#hQ�ȓ)Xڔ(�����}al����ȓD�,�ȇ�]�(=�,AgJ��q� X�ȓf�,AXTg�x
<��E�1�DY��9{|ͫ��@59�f
s+��p��e�ȓu�VX�#�P�3�v��'��p��MGy��'�?�� �£w��ѺhY�� �9D�@KF�Ӡ~�`�f֛�����2}��)�""���C+L�)��Ѐ�d�~K8���:�$��V��Js@�0){�|z�Y�,!�D�5o�8� ��?D� )���s��������	�L���Gj�ZVs��S=Hx�C�i�6�P5Y�εvj��*/D����l�"���g��p*2tQ(#D�L2�d?�.�;sI��]I�������t���EՐ���EO�'��+w.�"u���D1���3�� ��B�w�6Hak�F�!�U�&}�%��MV�B<���H'M��G{ʟ6�00
S��!�,z<H���"O�	�tǔ�9��q�W Ã&"�}�4��P}"�~/d�BO
4I����Z�B�I�]�d��/�24�� �c��O�BC�IA��Թ�� �/��-��F�{g�C�I�y�v�%KV���HD�G�C�	K�`���_/mҠ� ��w|�C�I=d� ���M�@zFpw�-s�C��(m�b���*;Z&�b�ϯ<֬C�h����Ř
R� "����$�2y�|��M�Nc���ջK�!����d�!smZ;Z]�nE5�!�ˣ��]Q�Dκ���4bB�n!���[�8B`�V�`
� �P��\T!��b������=0^r���=@!��*d��!ؿQ�9o[�),!򄝖I`���BH�lⶀ0ՃG
!�ć&~�I�Q��Z�B�
 w!�j�v�:Ef�^��B3��V!�3�!	1#��BH"��NӸM!�
kZ���`�4ra�X�T��6J!�$ޤ[V���@Iv���޼1H!��\�BqꇤŰ^C"D�@�Ҫx!�Ɠ=I��mN7
-z@�T�3+!�d��&-h�!
2uˊ�Y�"G�6�!�$�*�fq���j��xK���@�!�� O���˔$�-	O�	�b��/�!�Đ$�p�%	�2�	�C��&�!��/����
��h���˃�od!��4E�Ѓ�G�j]���1K۬5v!��C'kT�;B6脔)4`Pa!�$�'���	��Fir41��rM!���\%P����$Y�1১�[M!�d�,9|yS�Wk�`'(�K@!�$o'��"St���0`Ξi!�Déw?N�ʶ�LS����rH�!��P'���w��l��i��EE�<�!�� ��8�L��=t�w�O� w��c�"O�{�@�'��`�U�� d>5Y�"O�eP�C�10tdX�rq��{�"O���U[Bya@	��h5"O���.4�,2��+�|�D�'���'1R�'b�'�b�'���'�ȥ��k���ր�(L�� J1�'��'92�'�'���'���'c�A�E�<}G4�k`�Ƙc��'j��'�R�'��'3��'r�'68\��щ~R����j�%��,Q�'��'�b�'4b�'B��'���' h�q��I�Pֶ(JV郎ewt�)U�'Tb�'��'}R�'��'Vr�'���D+�=�\���0D,��'�b�'��'cB�'��'b�'Ԯ�Q���RS�C�*pJ�ćU��?1���?����?����?q��?!��?���Ku�<���$C�a!�J���?I���?��?���?��?����?9T#Q�-���s��!o�j��d�%�?!���?)��?����?���?���?Q�l<q���1�! $�F�	��P	�?����?���?���?���?Y��?��E.f�[T�\��YՃ�?���?��?Y���?���?	��?�e>Hh�CEB!	��&�j����?I���?A��?1��?!���?���6�L��7 �XWQRf� �B����?i���?!��?y��?��i���'H�p!T��=)�V}��IB'�� ��ƨ<Q�����t�ش�V	;t�ծG2�1��,r=�`9�kp~�k|����s���4	&�+BB _�hк���,Un���v�iP���a.�&���!��1f>�EhP�~��
#J�Q8G�ت��e�qA�c��?�)O*�}�d��MT�.�&W=��G�P ��i�h��y�����݌F�By2B$w��ɓ��#��c�4BN�V8O��Ş`W�Q�4�yLc��4pPBxT��Ϛ��y2KL� ]@�@$�Օ:�ў�S؟�X��)ol����O)k }�a�a���'��'�&7m�g~1OLY�����d� �S�B7M�n4a$�4��������%
�4�y�P�p1B�#�����f�:\�|u'�=?9`E-�VEn�c�'%�B�2]w�:�dֱ5|��`��	�
a��$[2�d����O?牜$�
�D��Z��/l���	>�M����k~�.a�����k��8҄ұW����WhN> +��1�M;�i3�MA "ț6��d�W�O !Rȋ�m\�z�)��ڒ#���s�z�JI�FP�Y�L�H�Ƈ�5Ӡ�@�(��Kz,U�TI�\��n���eEׅ0H��H0 A�����U�F����@��>w���'@8/vU�EK�V�yZ:���B����O^h
�F]�"E���
dq�EHQ��%vtY�M�Q��Р��Y�Q`�&�B�O�l}�4� pY���Ї��32��dFR��
t�R���26�Y�v̕JS.M�'��iɣB[�/[��CY�.Ѻԙӯ��&K͜;���#!-�	-���ń�-C6��X��
&)��yq��/c�BtI��h�����O����"�'#V�h�+ٲ�D�!@���0��!�4�?Q�,S2%j��?I���?A����S�U&����U�kX�QaQ��a�\6аK�½nޟ����0�S���|j0(] .����E�C��I*�͓�v���j��	џ����?c��	Z�ֈ�0���1��X�D%  �4�?Q��?����#w㉧��'�rE�-'88�g�A�
	ѣa����?���̜�<���?1��
��Q�O�NQ�C捯]J�80�i2EY���O�I�O"�D�<���=9� i���]f@��v���?��'��Yh�y��'���'�剿Y�.�H��.&�|�zgB�Y��@%6���?���?�-O����O}@��=�Hӧǒok0����_M-1Of�D�O���<��N�9>���!=)b�S�h#�I"��@s��П@������'B�'�Q��iYVA�Cޚ$kQÙJ�^�h5^���IƟ��	ky���)c�l��U���&�,u�@�I���ȴf�����	�\�'���':N@���J1WaD��UBɋ[:
HÕ!�&d�7m�O6�d�<�E�D��O���5v��VW��a��0v�^�3���'�M�+O��d�O�!�1�S�?7��) 
L�fGޠu��%)�5-@�T�`�1����M� T?M�	�?���OB���OM�V�fM��fKg�,�ӳi���'CJ���\��&��Q5�/F�|�����	�N`�J �2(BϦM������I�?��I<�'T�r=����~�$�/N3���)�i��h��_���	��`�3��y2�R$���6�JB�,�I�dU�Mk��?���X�F��+O��O�����Th�iĵ��Z%��9Ⲹ�C��:ɘ'�&A9�m-��O@�也p��
N��lyD�J�/v���FDh�\���Z�*ʓ�?Y���?)�{b��6WͶ�bj�_���3�/����ߨ\�邓�������'?��#(�v1�&�_�&�9b�ɨ~�(��Y����ܟ`�I`���?ytE�u��D�E-��B���x1�˧D�E����k~�'�rS��ɖ5� !��F"�8B����\j��P�$�o���I͟\�?���D��Xj�@N���fA��WL*�ͦ(�L�2Ż>����?Q(O.�d�<0�b�'�?� o*Hx��@J���P6>r�*��i�R��O��J�k]'<&�'J�%�w�5W�
\22�k��ٴ�?�/OZ��RȐ�'�?y���ʲӋ}�)��k��|c������+i�O���_�I��Q�T?� ���6�ZR�P�G�.3U�Id^���I+V�h��I�@�����MyZw[�/�eE��V��')����OR���´" ���Y�e���^�!��r3��:<��F���b�'g�	�?m���D�')�PC��F1'Y��sv�R��>� �Ff��P)��ԉ11O>��J���c�|F�)t�V5�
t��4�?����?i"c���4����O8�	�0�bmA���H�� �,62���y"c�����F���O����%Ҿ���P"]2�Ԩf-@��$�O�a;Sk�<)���?�����'O�u:���!r���F<�TI	�O�}����"J����8��{y2�'!z �JZ	b�i$�+ �D�9E����ڟ,�I����?!�]Q���q��4
 ��r�R�j-�W&,fHf��'��'���ԟ�R�@�4�  �����F��kE�P�U�	۟t�	��?�Sf�+<R�pn�=_�h�	T;'s&�R����ZS���?�����D�O�=kD�|��'�02g舱H�N,��$k�i�ݴ�?���^���pA9���n�FЅ
U�!�Dd96Û�@����'���H8��w���'���Ò1����$R<E���öU�2 v	1��}yi�O��A�� �D
)���1W��R��Iȟ��O�L��by��O��i��:5dڕc�0U�F��<i�`b�>1-O,):��)�+t�}��|����$-��&K�-B�'�2�'���S���֟�Dau�<E3���0Y����I����E.��b>Q�	u z��W�ð P8=�"Ń7`�\��4�?Q.O�+0Ű<�'�?��~��A3{oH���^�Y>�݃��'��#<�����'�2�O^��ٴI�V�:g��0�H���'���e_�X�������y�(6b�
���4��XӍTG�&��J�I$?���?�,O��A&1i*1aŌ1�P�sT�X�w������<	���?Q���'���K�3Jd���2s�4q�ӊ�=o
���V���D�O���<9�������Od8��e
>�����?Q˒`�4�?���?y�2P��ilӀ�����/>2p��� � ��Z�H�Iȟ$�'~�@��I4���A���1%$\�Z��N��X��د�M3����'��ɾ1CvOp�{���~i���7KB�Ϥ%�@�i�[����V���O�2�'Z���?V�XQ!��c�x5b�)člr�b�h�I�<]��j'�~z(M:u\)@�.��;�Dpq)�X}��'�8e���'��'�b�OO�iݹ¥o��	3��@���*=w��O�>���Y|aA�o�S�S�J��tK���T :�CQ9�Z�oڃBGjh�	ԟ�'��P�����F��"+ͼX��F�C9Hb��L �M��LD��"u�<E���'����Bo�6)Ჵ)��ͩ.��E�R�|�H��OD��M�XH��|R��?��'&��[�m�'�JI(��N>x������$扂J� N|���?��'-t��v�V<t|V��v��/q��4��4�?)K)���O����O��,AG��0�}V��~���:ͳ>�%�;]���'X"�'��I����Ƈ�vY��$���b�Pl:b�!M��ԗ'��'�R���OB�&�R6eB@؈���#)3Z�
� <+�Ҙ�ћ���̟��'�!ҳ���9�8�s�ƍ8f�f��[�01���'f��'E�OX� ,Y<9�2�'nʱ����>9��p��!�~��'1��'��	���a2�R�d�'��1�c)��t�� saݏw=V���ia���5�����!r&:
� O�t!G��r�j@�4�ܚl�ӿi�"[���ɶT����O�B�'?�D���B�1�2�Vk����)/}�c�t�	�Dĝ�0�5�~�dX�}��0�&�̻a�4����Z}��' ����'��'~��O^�i�%��Jލꎑa�EP^"bx�o�>Y�<����,\O�S�'�$s���:�IQ) ��Ȧ���
��M���?���"���?9��?����(s�vl!���'f�1a�H-k����$4��|�O��O�r�K�lP�"��4on>ā%V�=c�7�O����Oz�AgS��%�	㟼�	ן,�iݭ	P㑱�d�3B@ޣ7K�	Bk�h��<�q��<�O=R�'����)����:K�ڜ����:?�v�'p�I(�y�.�D�O�$�O�4�O}�DR96Hܡ���#J&��R&�C�l	�6�V�?
 3�'���'U���'�2\>�����Zܡ�HЖu�x�6��~_�h1ٴ�?i���?I�%&��Ty��'��	�ڲ2��a6eYQ)>�Q闩�y�S���O��<��Ny��b}x�ӵȤ�]��bԏ�0&	�Xc�s�<��?�(O>�d�O:����^Q�� AdI���α�D����r��-�'�p��q�'�_�z⣆���)�OfIY��@
�PM(b�ې%nh��b榕��nyb�'B�'YhA��'1�T����I��AJ��nZğD��[y�d�C�^�'�?�������Իz?�2���m2�	IS)X�&���ٟh�	ڟ�R�}��%�8��vM��}��ka�m�>��w�i���'���t�p�d�O����2�)�O�L�# JZ$�{��I�lv���F�S}2�'~����'2�'l�!�O��4�V<Q� �$A����ӄ	0 ���l��ȃܴ�?!��?��'�R��?���	OJ�[�&�r	r�)5eC10GJe@�il��"P�'�ɧ�T��$�'�� ��ۧ.��t�بk�NU�,(b�s�i�"�'&R ��rV:6M�O.���O����O�A7��9��a�P1���]ޛ&�'�剦�Z�)����?����h�K�۟Z�*�â�G���i��-�2y�26M�Oj��Op�VF���O�(S�n�1�L��!�P�$�ҥ�U� ��(?����?!��?A*��}�$
/#�"��r��;A�̡���	� �P�nğ�������	�����<y��K, �aw���D�����Bl��	@��<���?����?�/�b�� �mZ�]���ϐ
yV�Z��?�pi�4�?���?����?)O���K4�i`Y��W�/�v�#c΃0�mY޴�?A���?��-��SJh8۴�?��(�bTiG��f� �����lLl��w�i���'VbR�4���^V��ȟ���<D0Q��bU�}� �t��H��n����۟�I�`�����4�?9���?��'D�$� l�'0�����,/V,B�i[�`�	�Vv���m�i>7�B�R�z}���o4(����3%��FZ�0R�Ѝ�Mc�Z?����?=S�O�4@��]�X�F @(L���i���'I�0�'��'�q�`pz�k	U��5�PNO�0	D�{ �i��Qz��u��t�����OT��k�ß,�.S�����	S�3�މ@��M�Ʈ���?�H>E���'�L	
�b�:��0�Ld�d�q�{�����O����<\�`l�>!���~RA C'zQH�"�@��3g*A��M+H>	��U,��O&r�'A��hRЕ���X�x9�h�<V�@7��O�Y�� �Z��ԟ��Il�i���j��q����-�c0�ݹ�/�>�b���<�)OH���O��d�<�ȟ��4�EŊ�YW��[wm�B�!&�x��'�B�|��'�"`�0)y&BʲGhd)K��	M*���'&��L�	����'G^=�P�b>1/C�MI�Z�V�GǸ�rW�>Y��?�N>Q���?����?�?���� ;���SF�[0z��BFQ������ܟ��'J p�!4��N�9��%s���><����d�g��lZ�|$���	埸�$�u���O���C.�Vt0�&��b�e�ic"�'�剦h��@:O|2��BC��J��0Q��U4^��r�0`��'i"�'���h�'�ɧ�IW�3C����ɱ&F�-�$ _rF�fV�P:p�ؔ�M�fT?��	�?��O����f�*8yLmj������,���i0�'f�H����=� ޜ��E�l�|l��ś�S�@6MN*ά�l��t��៘����ē�?9��Y�?4,�NÍ0ؔu��L
�@�f��%�R�|����O�,���*cr^�`t��B1�Cˇ٦���˟���$e�v+K<���?��'�<�Bc�)[ݰP�
�8%<�cڴ��m͚Prǔ��'�bݟDLp-��Yx
A
@ir��]�c�irʗ���%����'���'f*D�3�@w�A ��"RwT�"Ԁͳ�����O��$�O�	ӾL%�^˴es��'��}����LS�'	�'��'�'�JDB����]���ʌʤ�3�! ��y"]�0����@��ty⋂�d��S�#9�؀v�P#�tĈ@c�'��?��䓀?��c���yy��܃w^L5᷄ɨSK�D
$R���	���7�<��B�
H�O�i�,6}1��sT&#Nd*��t�c�R�$$���OP�������,}�F6d�XS ���~�@�ڀ�M{���?�+O0�I�#FI��ϟ��S2�`H��d�4L�&�1l_L�2UzO<9��?�g��?�N>��O�����CgۦE3p�V�EDvac�4��DY�Y��!nZ:��)�Ol�)�b~�e�#I�P����(y��a��C���Ms��?��.�4��'�q�ģc�͐"Vh�b���c�,�"�io�!b��j�D��O��d⟄X%�D��Cs6\:S��H1�ǀ�"S�(3�4F28�Γ����O����~J�� 2@�u����Bj+U�86��O���OPٸS*�G�i>��O�!ڦ�S�D�@�X��Ѧ0l���i��ꟴ�D�-��'�?����?Ѧ��:R�>8��aڢ ��M�bM�V�'��! tA �4�*�<���V0O��ժ ��Y��*�Ӧ��	����՟���������\�	Ο@óJ�-J2�e+"Cվ�f��T�uJ��	������l��m���h���K��qcCR1~�"��PNT&�� �"�	Ο��IПP����Y�e�,���	� �5O,��cW�٦	���� ��R����$��Q�P�ˤ$q��y���b7	���	v2���DU����ßt��fy.�f�z�'�?����U��D�(�f�����LM��3���'P�O�Hz��+�	IF2u�D"�#/�F��`(���6M�O*���O�$��i�����Op���O���J�hx)q��G�z�c6�̵3'.%���ٟ01Q�ƐZb��'`��$�t��$���;#�߲n>x�lZП|�ɤ��x�	ܟ�I矜����i�i��@�&�x��C$�v\��Cy��D�OD�"P)_!1O��Re���W�4�fx�Γ%[�^���iЎ�
v�����O<��埰�&���u�TD*͸��sv���Ox�0��47����Ϙ'�Rb��~�btg�6.H��e�6a��7��O��d�OJaЬ�<�+������x�M�]W�$�R�L'���cJN(��'7D����1��O.���O�1�.�=d�d�a T���F�⦩���-�ZX�J<A���?1L>��Ґ�zG��A52��n��%3�!�'�$�*�y��'���'�	�ʀ �	�6a�$E�H�]%C����-@��'���'?�'���'и�  5�L��%�M�oOb����'�'S�]�lR�f���t�I�|�$L!5�Q2PXā� ߫��$�O8�$,��O:�D#����5'�px��֏�v���D(
U.��?����?�*O�l���N�	0�Ia�� �c���2�a	W~d)Aߴ�?�K>Y��?�GZ�/.�Ġ�	>��%(\�o�ퟤ�	`y2�-�������!�Ȭl�V��ZZO�(z��t�I��������"<�ON�R��'0��j�"�AҀ�a۴��d�bƾn����O���`~b!T�K\���j=��OC$�M���?��G���OX0m�t �DT(k����8�W��~0h��C�h��)�ʎ��u�_.����#fV��5UoAH?q"�h�ؠq6ʟ�YWJ�8R�h�<y�I5W*~����$~t�8(� ���ecE|�B����d:jA�L?C.��*bL���f"
�褣���)Z����J�3C^]`�!:��	�#�x)�TA�$9�v�kх(T��s-��I9��2S��A�A %A��ܒ�a�2i0DHȳd�2���G�CBl=�IɟP��ԟ��_wD��'��S)�^8*�b)����r�Q��z ��"BZ�l�"?/�Q	2hX�'h���Mٯ݄��%�C�n�(�Zӧ�?٘�Â�B�_=�4�t�N4��ۓ��'<�İj�|�ԧC�
-Q�9+�v��tGٳ|�X%��c�a��_�vQ�U1��Ȕ=*��
��+�y"�
(��[!Ä"/�vժ�kQ���'!�6�7�d�+r Zm�ퟴ��!�X�Ԫ��Z�P�v�ɝJ�!��៘x�����	�|�&,��7e�t�%�Ezhh��4D�5h���9Dfh�P��9w�Z���	A�ؙ�R�K�<��	�&rh��^Of(		�ȋ%,��C�Nm7H��V�R��"��=� )F̟�iI<ɐ�Q
��3aV�-m��	@D�<I�!O:|�ڄ�p%�|%��i�@<�T�i�V�Yë�m:
����	r<T�g�| ��s>6=�"�Ĥ|&�?�?�uO#h-taY��&_{LP�0���?���]KX��vA	=85���f�H:Hz���.�>�'M�(yF�Q�%A����/!l�O$���=1�X����&��"�	5�Ouf��&�Á\xqb��h�kI�0����O��oڿ�H����j+��-Ǚ#X���2��#~�"C��#Ju��F!P�5�vȠ�H�9RĠ��DI�'����bǴ/��� ��U���!㑈�>����?����1;�P1���?���?yD����vG�����b@�kՖ�zp��6x?.՚3LBßD�Jĵ0��b>�Ox� w���$"�[�� �3��xk�bor}���_��B i��P�q��'��QXg�.��%��ޜIm(x+��'t��<8���4���=��J�n\�H�����4��J�<��-Q�F%r��������I~�&�S�tX�d���p0��,�!P�,dXt���'��з� ǟh�	џx����u��'�B2�>\B�E��^0 +t!J���u2S�L�7*1��Ŝ�fr`�SK1<O��H��� �ny2�ǪM���Q+(���
#+��v�����(Vaxr�U�i����)D�m34��4-ɓ�\���?Q��$=�����)��a�<R�!���G�C�B��;4Ύ���-ݰg6�e*� Ejc��ѨO��;Ԛ8c��i��'fp���	Z�����#X�&��#��'-f3��'J�i�b����T�6+h�kF�j���"��9BH�y��C򌀛��'�ʩ	��ȋ(r�izQ��z�d8AD���{�����.׊B����Dv��\+�3��a�=�'�
��T�Ify¢ܱ]H�YHQ� v��;$b�y��'0"��S�HܦA����1jd��:>lB���M@�Z.�ԙ�&�(��A[=�?Q+O֤��Ħ)��џL�O�·�'p0 j�T�_���XC��`9B�ɦ�'bː����T>�P�*�QA\9;xNc��#)+~�O~ {��)��+��!۔+��V_�����P���'��\��]ɧ�O��p�o�%R��2�3Ĝ���'Ԫ�Q�H��B3`�ZC�>u��]KÓ;푞pS��F\T��Ae��R��=�	��M����?Q�f���"�?���?��Ӽ��� &w�P���	�~�4����'����ϓtp�u&ǝ�(d�q@(\�WH�=��rx���d��9�R����f{ ���AT��e ��)�3��U�<Mr����!����/�4.8!��6~�㦈 T�����E�Y�ɐ�HO�	0��{��%h��7Q��ɂ�g�H_���
7[� ���O����O�!�O�21���yv A�yx������S|�]C��-_~�h�a�ŀ\�
�`���-p��-`T�8[�|1�G�G{�)������/�
d��z$!���*��oh��`�hPq���h7H?Yp��D�Ȧ�ڴ�?q/O`��,��"Itj<ö�9r�t@eǋ�
�B�)� "]�#� ��d��%�`�y���ܦ��	yy��6a7�6m�On���*S���j��D�^�mR�S��D�O2�3���O2�D}>�C�_9cX�$�4�%�Q'����4�	�C$O�!9c@ϓ:#�O��q2a>!�}�#��+�n���'�l�����'1
p��oT���L�%�	�d��'<��kק IH��I�9����'�t7�<s�8�faU�I7 �ЦєQL��O�چ��ԦQ��Ο��O1N�R�'&D�b4��@Ϧ�@ ��*�+��'���=`2�T>�EFTkC���т`�F�:/!Ҵ�O,���M=F~� �%%�q�e�l�!xa&�� 〴�O�\PS�'�1O��"�/$iJ�y��$�#��"O�0P��epTL�dp��#�'��#=�'�p��(R�����.M�B�y����'�r�'4�H�uG��R�'EB�yG�O�[����Δ<D�t@����8p�N��7#�"�b>�Or�9�@J-��X:�M�ge��zw��Wd�4�0���>�3�d�;D� �@��"����@I$o�,��d�B����?���?�3M He��Ьou�v�ǽ��xb�E fiA"�ه J���bL̀���L�'����'��	�*�"�C� ׵�>e���5_3<�뇖^SjY�������ǟ�K^w���'�󉎷)n*��E�	I�f�b�jL�w�\�9�O�=�F�TR � 1i��.���sA˳q�!�$TR��5������Qa��=7h�9#�'�����C�'X4����_�Y!JYBP�\(tM!��?@(�gK٪.uV���V�F01O�o�m�I�1mx)�4�?A�=z��+@K��j�֨����8�d����?I3ƙ�?����4�������(9Yt��ѱi�P����%b�!��ؚf+��	�a7N���T�QK
91���Mq �x���#��P�����LVu8�X
G�Or�&�8�dF�v�M�$B�-Xe����
4D�|Te�R��8#(�\Z�h�n&����4P?�5`�K �
16��`ϼx�dM>'��y���'��S>b�������*p`P3$"�������,�	�`M��!�V��̤�w��)�?�O5�ӂ)X�ٵ��v��%����'`�]�r��=\�-r��O�	ב>e���@�ıQ���UhRm�d%+}���	�?�C�|�����0�l1�d�N:QaN�%�y��ȦG�`�GN��4E�$���0<y��"�r ��L�+URD �_m�Zq(�4�?����?Yg* Y!�� ��?����?�;JJ�H�ƞG�|��c��tڸ��C�)�ȅ>����I�ʘOh�'��t�&�
^��/��Pb!�!�A/@���Q�
�<8q����Oz�'�b4�d�X4�>X6`�8^��ǃf�to��,�1�ß�>��?I@h�7l��� Ɯ/���B ��;��x��(�j���Ʋb7H���� ���
r�'�n4*f�'p�ɓ$�X8� F\�Q`@�HU�)$�i�&�5;����ǟ�����XwsB�'��R�)[�hHf��8	�J$#d�K�W�\�ÈTई�"�)x/t@��I� �P���;� ��JʖNl ��5/M�B&	L�v��˓iZ�0�b$��: �Ҭ�=���T��dz��8@$���<M`�
t�,�����In�ɴ{N���a,��<G"��� |c� �ڴ��=)�Sµi{�'i<�t�3�y�v,�lN�2��''B*R�o�B�'H�)��Ҝ|�/E49���7����q$	��p<����U�M��E`�#Q��l��jK.a*8���I�Fyn��j�I�(=�+S�0hl��I��c�rB䉍g]���;+!�Y�I�ϮB�I2�M�&m�;EH�r�	������_��h�֬�ŷi�R�'1�S���|�	$T�p��M؛Rf�Z$)�T8h��ӟ����˴E�"8�B�ʿd���ص͖H<f��Kx��nнFn%16�R�}a�ܱӀԂ��	4w�
h�`E��_��D.�$�4�{����}���ø �މB���9���'t�3��rɧ�O���0eH$X�<���m�.+�<0��'�@��N�4th�hcnڊ!P�0:Ó
����"
Ҙڼ����P�n��peL��MK���?�4<�G"_'�?A��?��Ӽ�c��[�QRf#��H�ђ.����'R\��	�E ��%C\��<9��a'5�=Q��ix� 0G��58��VfF�1�!U�A���5��)�3�DQ����ԛB�>��B�,X�!򄉈��`�i�qO����/C�	��HO>� �c�n�@zpѸ)��2���i���7g�v]�v'�O���O*���Ⱥ����?�O�B�3J�?!lPٷlQ�.��9�r��2q��|�s�BM���I	�sf	4f>7��Yٷ8gDba`5��A]B�)эJ
�P��I���j"a^� �8�hF��d4F�Y ��O�х�	�pxV`�4ɔ�r�n���D9`R�B��'5Ԅ���"_�N6M�3d3Xt�b��i�}RK��^`7��O����r�u�p$Y�!?���%���[>���O�P� ��O0��o>y���Î5[BE��^�2"��	��
E:!�/"��dX�M*/=�x"��n��gŐ޼P7�������LǵuKv�fiB"iZ|@®B*v�t���"I\�_;Hi�� �MC��iK��J�Jx�-�e�I,B=ZsCa�n��՟@�?E��� �b�y��'A�0Xa�˕/�xbH{ӂyxP�	^4@E�� ��Z���E�OV�>�������?�����)\a��牻*Z|��u#WjN0�㝈|����OR�	u�,cZ��YA�*3`P��|r/�ʈ��b��P�z���%"�Ւ��>ѧE
�q��t���h3��i�fD9bAvX#�/J"j P�S3z�Xy���O�4�3riG� n��'�Bi���?)H~RO~�c��-˸�I�쏼[�42�d�o��?�ϓk�f��Э�5Z>5x2O��x���:�HO��"��&d<�i�tO�%����i�ߦm�Iퟐ�ɲKU,�����ğ���l�i�!P..zc*����ޕ �4 +d�V�4��q����#�?��j�t��%�|&�h���37J"�)���6Q��"&��e^P�r�&�2�"��&����Ű$���M�2C���#D��0��X�"U����`���7�?��OV��1����?)���?	6l�	~�"A{�-��l�h�#���xQ?jx��oR�!�bq�I���D [�'����'��	�,�Ԙ�J[�hV�$Q�|��K��J!�A��ß������Zw�B�'Y��Y��v�;�D�h��t��傽, $̓�hG�i"��5,@5��󄏿7�1k�mB(G�DH��I�mکIR��L٤ R���\$�8�"���$g��R�j����'�x�#�Qz 
gc۱%�����?Q	�v�X�B��{v*U Ջa"���D���Ҕ �[��m[� K_�d]�<�a�i��'��U���>��O:D�B�W o|*1k���>"|�<Y���?��Y��?I����d)83͜�{��׬F�����h_d��IR 7�~]KA�Y9 �B����7` �uψw�\4���`��q�ኒ$D�Q�b�ۅ��=Sv��Ħ�ȑ�ơ,J��@r��O�Yl�2�M��D����F�ݰV�LEڃ�V�#�L� ,O|��,�)§A&��7�Q�'z����T�^EL��>ٛ&�T�Q4(�k�S)�l����\*�"T�8�ɞ�s��ß@�On0�K��'��X��eU�r�@X)�K˭+�\�Y�'>�lN�K�ll�CA�B�2��O��n�kK�o��a*�Du�ZE�Q�Į��I�-�h��A	�M����ҪS#L�t�R�i[�|Y
Ty&jʺ��-�� �1�P&V(���V��k�D��:Q��'��>��,8� ��
ְ#*C�I�*���p��\ o]"?���K0k�x]�X��ɮ�HO~���MK8Q�HqgO�2WԓqjަA�Iß�I�d�"h� Zԟ������ɯ�u���vɠP��f���`1�ȅ:�1O8r�'<�����>1����%X�,��2�{b�P��<��MƤ3��LX�J)d�``�Hj��'�h`0�S�g�ɍW?�!Iיo�*Q�v�}�C䉢�t`#牤-U�h`Q眃S�V�6���"|�D��Mv�p����[���ZV.�O�9{1�@��?��?y��Iw��O�|>1�%�X�?�*�A�%בI��@h��؁#�DC����0KQ 
"�;d�͵ u��s#g"�,kQ ;(��qR�c�8`�`Wfڹ}(��Kg؟D�HG�m���cn�
��L�u�-D�����G�U�̫4"Ηo�P��
+�	(��'	�)R��yӾ�D�O��5dˎ��X�,ɍqH鋴��O���<�����O^�!�h�d(�$�n=l�pc/$�>���o�3 ��x�ϖ��'b��q�+B���%]w���cǓKD���f��$I�jU"�ʕb�^=q�!-�C�I+%�xt2�dT|���$WPѮC����MK�@A�ky^�9�W��(��Oj�s���B׺i���'/�l%H��I:fZX��'ۇQk��k憄�4���	��< G ��,�<����؊_��%y���"J���?/�f���Ex���/R�0MRp�`�u��L���U���	;�F���k�)����)�-~ɶ�{@H��e;�C�I�XZ���B�'
,ʐ��gJ:X����G�' t�GL�L���"`ڒ<H1S�!`�����OT�D�3?�Z�1��O@�D�O��4�� �	�͙� |�51���!7�����B?�	� �X��$��X������>�,�9�OT�8qOz��d�'Vp	�.��3{���d�����*7������L>�"�G�^����M	<w���3Ly�<�B��Q�ΉuHA9r �C��[~�/�S�O�^`@V�ߦ���q���XI��Ηws30�'�r�'����a����\Χ|1��s�LH����k�*V�.T!FKU<ɁkA�C��;{��8�p�ˬgtm��$2� � D�x��͙w��v��qR�S�^8H��\؟���P�H!N�zTb�qd�`��7D�,g���!Spm@T�I)Z�,mjV#)扖��'^�x:bEi�<���O�r�iA8p�J�xs��(V��d)�O6�$��R���O��ӨJ��ం
%��C#�@�b��1B�J�*&�D��xbDE�[����<��DO.^h���)AX����e_G8��h��O8�D�<Yc��7��]HR*��*L�AB �<i���?I���)  k(ͩB�;^���
MA!���ߦ�!Ն�x�����S!���"g�D�'�L���'r"�'��S�3vh��I(43�����nS �a�A��6�0��	�d��#��M+O���|�'Q�a�t���0M:��Eڏ
�<��K�Tk6ŪW|���!�'����B�E�n�v��^(ٓ�܃'=��� N���AJR�>!� ҟ܋ܴA�f�'��<�Z����i�d�H�nquD�!�N5�d�O������{,��!Pf�;Gޑ�F�F��0<qA�i�7M�O0�l����g M�_�<D)�*M�JT���	�{�0�	Οd�	*|p$�32�Lџ��IΟ��	�ugn�($,�a��������;0�0��a�fa��d�'S� :p�|BOH=%{xe��c��dȉ2��=�"Z��.)Q��$U3@Ni���L>�%�Ǳ2�XP �k��#��I{3J��NC���p�J��ɫ~Ҡ��Y���I ~3$|�g�Q$UL�vÌ�'����Ɠ+��U�nK ��(S)B,{7�,�'�R"=�(��ʓf�|�`���%L��s↩5f^̆ȓ6��p-�xa�ћK��S���b�<�G(n�
t���f^qÐ�b�<��iJ�8?�8��hC�8���m X�<ɱ+ƚ.��i��ֵl7Ԙ�	�Q�<Y�!� =�������@d�OM�<)@�
�dovt��(�h���Ad�<afRJy��@U�H$hcBLc�<�D�ھ&Q�D�r���qE�s"�]�<�A)B�}sMb��E���c��Km�<����~բa돩_t9Sj]B�<1��ϛQ@N�"E`Q��-�g-X}�<��#D�` ���ņVXJI�2$Vx�<��Hh,�c2��V�bpiʏX�<b�\���R��v�$X�)�L�<91�ݤyHR���/��cӒ=�%\H�<�D靁"N�{En�gq&x3�(�^�<	�@�:.��)�dؗ\&T�&��D�<���	#gJ��c��j�d�z���j�<�a�Ĭ,p`G$_�k��2�@�e�<3���7�]�5N�{��ˁI`�<I��"oҡ�ŧ	�F�ܥk�-^�<�3D �!�:�`��F�2��(�UL�W�<��W �$:�R��&��P�YQ�<)�炭o}�9Cƌ�vXl:`�BK�<ɇ!Q:R\QС^5�b��o�<g�V�@��T����j�`���g�<i��C&<%X@�"OT$l����"#�M�<�p��.��M�� ac�)i�DH�<��3�x��oQ�+",d�f��C�<�b�'=���+��O�7��DRb�U�<�زe��8���$-� <z�]l�<q���B�li�,ң]�ND��(Oi�<!g��{h��rw N�7#x���M�<��jj�D�����,��KL�<��K &8�Q���W��,�� ���@e�C8Eސ{��"Z�Z��'���X� (y�""�,d��(��oW�(b2"O�|��v}B��`������؇i�X�Dy��O�B�� # ����8��8R��V	2�8��柢�94�'̒�f؁y�(A�DF�qjؔhd�K�k�@�ku�򤁕o��t ���%��%��g�:v�����C>1�<��a́=K��	a��W���@�BE�<��x����C��[���D�� 7p�ש5}� y``�)t5d�
v�0�P�c�'�p=I�V$��0���ؒ���쌅Taj�Vd1��X%�	O�Y���!k���=�`��'��Tc�!f�p\ ��ɮG��9��ɞO�!�dQ��hb��ld�%�a��=t�$�Ʀ�� ���`7����'2���%(���减V��N
�� � �̺=ㄉ����\ta|"D\=$U��্& ��ԯ� hn`q������i����@q��4Ox<�tM]D��Q�SK����P2b�9,��EB"��""cV�3)!�3�"$����7�r0� L������i�Yx��\�yIAS��դ��}�UF�.K����L%�^LX��g���p�ǈ�>7���ͳ-X��$�('��	��k�-|I����E�y���}Ӕ��5�� �l���.6�>�����I�.(؂�ߩ@J`̅ȓ;�*�q���>����RML*Sd]���B��V�V;_����e�����z7����E]/n�d\�;�f�i��)Qǀ,2��SM@݄�1g�h�(��."��-;��� G)(]
E��L�b���/���~B�BO�a8��=��<�Cg���"�'�p��'<�;Q�Y�]8tt2� �e�(����y4Y2�ˑ63`��lD!�n�$OnN� R)�a����4�
���9pb�O2Y�`,3��R%�'���V�ɕ�TL[�Ě�RҎȳ�Ċ4`�\�DCՖaż(h��_ͬ�B��TMY�̊�R�ɱ�O�֮\��gh� �iKQ��<2h���mJ >!
b�V؞�1bH�n֤ .!%�e��K��6�t�5,Q+�D�ҊL$o��X��Bܼ�"�'C��/�n܃dȊ�8P���'�,�Z@��s��Ј#OȫNO�ڱ�[�=J>��s��[���.��)��ޡ��ɮ���;z������'Gh�i�H*�x��,�?�O����Ĉ	Ǟ�Wb�~���|�@�W��@�	�8��@ʤ!;Ld��$���AS<�u�ܡkpd�� �$[�!"ԈX iG�T���"#-L3Q��d&J��Af�
���rR�5�"+��B���O���H�ꜥ\�D��!�;�j�AE�O�$.�Xȡ�Q�{��뉹*��� th((bXcR��}�R��6�H���*�b���/O��
�ވ�'������O(B�Hɒ���9�%d��0>�v^�T�Tr��ûw.Q���2)���0S�]+T�P��O4�?�Dzݍ2W�M�b�B̟{(u�f+5��՛���':\���4V!����ft�3���t�jZ�dĭ8��d3�培#!F}P�MU6\Z���[���9j�'%\�x p�+��&>(\��p�L�!B$G�b!*i���Hg����!��?�a#���ˀ;:����B�U��F���'0�3��H-CD" �P��n.L2 K�3��=�O�ju3�eХ	��� )�P�[��B�"$ q!2%BSwa|��i�:��wE�4���B��N��MO�Y\+�<}28O���^��PPB]�2�8�@d��TvVxz��V�"Iu�K� �ExH��b(���*�{,�D�4�P����X���2A���^��Ç�ź5�m��;}�ϫ5��y�[�h΄�0+I�m�&�YS�CQ��R�\�M3����g��u%:��;}��$��W`�Q藔]e���!� Q���D��2�O+��E���J��cD"O���c$�O-0a��6}�קew<���l;0��eHA8�0>yp$S:H��x���*=��hZ	+�	�*��ա֋p�D��
k�@�xk2�Dr�	�H>���D�ar���č�f�R�+v�\�'E�A�7iér������;eM.��ST>Qy�M�8���� J!G��t@b�+�Ig�u�牍I B(��	�0J���s!�/�xٚ *� , �H�,�:y���e��m�O���� [�8i�X���,�d�Aѫ[��D��Ν5Z.]�VD6,O�<9�V� ��#��Cg��w�ݳsY`%{�ܲ�"�;p0���%�fD�K|b���h�2��(D�%T��ӳ�z������2j��ț�1"�H�V́�<�j|Pd�R%O��$��HB<!E�ʗ���*T�CY�y$��M�}��E9=ղi�6� <��T@B�'j Jd۩6�d�eZ7 �x%hEQ>YJ2#'G�n����>�"����d��pp`��_�>�$�Z�b>�T�>�%eMݦ�nm�BD�P��/V$9���g�BF�y"@�iybD ��)���x9����bp ê���"�Λ�CI�X+b	� q�2�h���
�p<��`��C���7n���E���<9�⟱<	�Q���
$z�?Y�脿Z��!TCި6����(�N���n�y�B���fh[���;,&����ط���s,�5��c�	��On�	���/#_%>IB3G�g`u�A	�%�L�"� �ä� n�:$����r�"�S�56r5c� cH��i�B��[g+Gf@�h6.�x&�+��,��<!���c.\��8a���	�/�"���9�ʕ�J��2���"~�<��{Cn�:.���H�!Y��ߴ1�Ȭ[�m=C �1 c� x�$F}
� �����ѵ�J!Xe�.m�u�3O\Y���u�fq���J���)�	֖W��Ųd%\�{���N��L��H�D��4�s�'R2`Bv+A��y'M/u=����)r8F����C2ў�?�P��z��Q�����7�@��X��g�'k��� ��Z�p��ggFb����'�jX�e��A�,y�	I�R:���Lݕ�hO"��O��@@��.�"8Qs�O���ڽwY�pK��>��L1o���9M�$�`�ad	-?�ʝ7���8C @P�'�0��c��S���
��ODy�}V�9�� ��8A�	*��i�&�>�����g?p��u q��#�M�x��0wHX�"zgA�+l�u.�d0s@H�?��x�K����E�wL�9R���PB�(7��& �x�c� Y� ��c���a%����sS�Ɇp���z6��?O&��GBE/[�4�A�޳Man�	�,D��-�O�r�v��+�`T٠L�>i\I�!�.��d�{�cW&Y� ��<����r�f�� [�7��arp�T$+J
Y#�f�>P��D{��
GwHD�ቻ60¤����T�A'�];
��k+<�D�6�~�q����P���=�~������hP��dK����(� <������G=�����8R����JQ���dFK�c�����5E� `>`��%��D{�/Y�+���R��*f^0Y�Ub^�W~��F��EQ�)񙟨0̿W�р(B!$�8�I)�S�6(Se�	�?/4� �Sh&���TXa h���#CwxO�� ����*��iXa����`	�HP���p.��"b��N���e�t��S��y�x¤a5���e�W�ZR����#�>�򧖕F$���'� tx�c�$��CE�*B�P�B�'��I��	���!�J�'�|��đ�V䬄B�A�;)�B�s�e�';��kA�ZH�'.$!����5��Y����r�!K��u��P�<�&�{5�I�l�x�y�mG�剃YN�"�HZAM�MK���� #<���
G����A.��zB�>��Bӈg3bcZo�ti��3��֔X^�P��F���D ;�F�@E��C&�T�s5�Ţ�I�C���P
���8QK?�I#1P���qf؅$�j�3�,��M�44�IS�h��OX��vŸT��!$
n��+���/(�ЌHcM�9r�"��`�X�B��	=ړd�̉������6��.J�QΓX�>�#����P�:)CB!�f���I�h�C���qW�Q��92�S�4�92��8��~��Y"@�q`d>}SBAۘ@XZ���K¥sF�ȓ5�w�� ���UA0�7A��g�=p͟T �H*�٧ ��Q�B��O�AP�o�E���hj�q�*���63|�- b�0_݈\��H���,`0�k�0d���S��Nd�+E�*�缓0+ARf��cfǝ���DK I3�{nD��#,J�@���)	sa�0�?A� G�*��j�`I�Lb�pU��C�r�ţGą�dN�pϧ�~2 b��%q��k>Y��ψP�!&I^�g!$2 C��X�����9"�G{�A8�էO��8f��"��ЇT=�L�qE�&/�!�&'|J��$_��l�	�0��bv�q�Հ���79�eB���(��t,Q�/���1e�rZ^9%��OD�'�A�|�R�����ql��p4B�|�+�21�|X;#�π4Y����͐>02-����sR�-
e�<%D�,��#���)]�-z�1{7<��b���
$��`#�Q�Jo��z�F�h�C$mE>R
D�p��'��$4�VὟ�`���A�b� ���>_� �qLO5l��pZ4,�'l����]O�u����Kb�"��6��0��	�A*ܽ)̼邒��+����dBܘ���H� 1"���!��F��A�	�<A��6:+,t��ɨ_�<���`�&�Z@�7�S�������#�o7�=�c�Q�v�h� �
ԏb����^p�@C�t2°�ꦟ��+:J�p����<��b��[�r��Di���i�2���ս]��
r�Hn��#<)��T�d)�؉?3�<씱��I�3tHz��dmv𸴁3T�(���<	Vf�O��N�0;��(�I���ua?&(�֘�Y���s'Ʊz�t[f�ȩ^��9�ֈ^���qGς!����	�SP�!K,;�O���So~%)��!)6e0LS�(>�pu�Vвw͝�T�)Z"!�P�@�x�#Y��'Ȭ����S2����ߚlbTɂĚ�-N�4#�bU�O�z���Fԓ�~�		V+�}x��'"�DݔwUMKq��h��Zw'�{���:���PO�@�A���hO��A�eNu ��L�y��$��!��)r��,�#�
ESW��?�M3W8Of!I�dY�l⚽�G(�3���s�޲f�
���(B��5o�e�'!�� �̍�h��"�iR>����V0vM��A�ǀ�|�ԁ��q���6O�8�r��~j���Я`l��ˇD�!���<��e@�!��ua'I��+�R�����<��pcN76�X��#���3���W���k5;����E��!��h8��Q�O7�P��aʫ,Z�Z� 9�����9��:�ϑ�w��"���rD���a��cz8x��l�'�$Q�'� 8�5@K� �@�9D%�29|�� M�����J6E��2)E|"�߼x��1�k�9����Q��(8�Ⱥ��#�@D{I�<!���}:>M���*b�@��Kjϰ!ا�Ϯb�D�`��.|!�D�($�d�2PLq��T��+�`���"B�	a�˧YP5B'g�2�>�z�$$�X-{�c��ms�hA�4D�����	~X��TB�}UtiR��C9!�����O E�SM�5>��qOx��b��p�f�@PȒV�:�"O� �����O&a���w�	/8cb��1"O��'��1^�z��P%K4f���pG"O
5�榞1հ��P��U�a�"O�\x�`O�*|�aⶃ��z�4`{�"O�A!���<\r����un�(�"O���FT�~�^�F �]R�h�"ON��I��@m��nҗZ���xg"O���-��b�"q���3&�X;�"Of�h2�Y�?�$0B��5p�y`"OJ81�
�C�ܴ���y;`x1'"O��8��`{�i;!Hќ%]��"O�I��ć�m�d�R�FE���i�"O
� D�V�U~t��hY�m&�<i�"O�}�0	R�D�tԙ'�]!�d	�"O� z@M$D��p�ӧF�C1 "O�0�����l���#.$���6"O^�����$4�l��O�Œ�"O��6��N�zhs�$T���"O�[�
t��隠��d�x<;�"O��{�KA=6����:.+���E"O ��0��6,��7���I�*�"�"ODm��`�,bi,`��E��lV���"O�|#�!�2�z����e:���"O"��'��
|U��

�\�Ԭ{�"O��r�X36%n�x6)1,z8{0"O`��4-�4M� S���.<�(eS�"O��хmM!� �Ҁ,G/����0"O�y�u��>ϖ�k�K�>l�%"Oz�B�M�J��ۇ(X!,���6"O`����@#dF����G�\��3"O� P�K�H!�Eʠ�-Dx@"O��Pu��b��l3@�R�+w"O漠�,@� �<؈��D>2�&(xv"On��c,�%���R�I��pS"Oj�W�D2�j�*6�C2{|i"Oa��]?��)s�F$jmhcr"O<uR �$F|H���g��,O*ܸ"O�S�$T4���0��:	A�<B�"O�9����%ݴu�/I�*3j�H "O��(5�F,=�6���Z��M�E"O,Aj�3��}��DQ� "O*��R���Z�y�*��T�b頣"OR�����u��2�h��(�"OT�uK��+ �"�Ǚ
㪴C�"O6B-˩MM�D1�ӈg��
�"Ob]9�m�_cr�jgo�Xm+%W�<�*�	++t$ Rc��2�h\	�gWP�<%��R4v���o՟gD�X�K�<�0cڄ88��	 a��+���2�D�<iC�e�Xup���WJl	J���B�<��y(�`{��(iڦ��'�Fe�<���&x)� BЃ��J9��p��d�<��ϋj�T��NϪmD����f�<ك��K���3�i�-/M(�9�Jl�<�2$Z��N�"�B�$~��Y��Xf�<�'W�E���$�(P��s��]�<�Q��=�d�r�L��UNZ0���VO�<�s�\�8���3Qa^�~��d��GCL�<I���nS�d1��2I�n)�FP�<��MTX$ -s�j�-_lP���D�<1��1O�]���[RZD۠��h�<�EL7 p����
�k?`�q�m�d�<9��=K��SO��W*�	,�b�<)e�0�DG�͒A��Lw�<� ��z����`���$��Psf"O6���o����bE�K����"O)�*
	Ytn�8u�Δ��T��"Odi�"��]MJ����/
�vD��"O�� P�cL ���Z�
��Y� "O����Fݏ>Ί��@��]�,a��"O����Q��؀)��Z�~@��"OH-qI]
,��$kq�L�X��`"O� ͕�\��I�J��_2z@["OR �'��G��0�Lwf]�&"O�ivL�!Se-��ìto&�"O�y����-:�NY1���(e0d�W"OT'kԽ@
j���Ȓ 88�"O�,��� y69��--����D"Oh������R�0�Ԅo�r�c"O"e���TzĶ��CO�#ל�j�
O�7m�B<0����"�̑1�M� 	C!�d�%�X�e�%E�XU�e���m��xr�ɪ`a,�J�B�2-�O�0��B�ɌB�ā�#�6^{0Q&�_��C��+f�t��B�8#���bD�yA�C�ɻmtr��Q�E2�tճ#M��f2�C�F��D�B�Ʋ!���[)+n���6�	�h�����0{�U�0�Z�N��C�I��Z4��&1������/T�R��F{J~�R�?U��9��a�M+H(�w��L�<тo�W�T�ء�U("di��DR�'&1O�O`0;����1+g�Z�i�~L�3"O��T��	p�$ÂM���P��"O�h� SL�"���5�n`�"OB��G��#�)�v��`��Ucc"O��k��=���P�	A�0�S2"O�-j���W�`��J�)1�*��q"O�`�sCoub��V	�-����"O@���+��h(�GN9/�z	x�"O���&̣����@f�If"O���&ِe֊9�e@�'�l�b�"Oܢ�!�9o!���E̎G��ܱ�"Ot���6]���4bM(T�2$���$#�S���c� ��a�<��M1�
�b�Q
r"Oʁ!�FI�G��9��!�Y�di��'�Q��1�5H�HdƀE�+}r��o:4��BEbw�1����")t��W�X4('!�D��8��|�w�Q�W]��A�N�y!򤁠[R4�K���(0�Lq�`X�g2qO`�A�$�0���m�=߂�X�� ��P$��D{���/��9�t�T��-&�����%�C�I�F�����:��9
`A�)�ў��	�a�lq��MR�I�B�A���&M�C�	�b0���ư�M��`b�B��/cp��`�""���1vɁ��zB�	���m�e�h�mS�]f�C�	�ϔ�Jז5K��~��B�&(�A��R�TD�c-�)�B��;T��X�c�}^MR�2:�C�Ɋ>#\�U�M�'�,����%�bC�I	s+t�MԀ#�\��	��%PC�	�J�q:1d	�7�(ⷉ
:��C�I�q#K��>�����R�O��C�	Sp�m`�Mǎc̐���N��C�	
l�>����)ofP�S����^C��-B�,�t�����S�9�B䉽�m����66��]�j�4>�B��;~�6�0��o6�ʕ�J)C��B�)� ��� 	¸&J$0�Ε�.�J��"O�ţb�J�t�*&Sm�z� �x��)�S����ѢҢe��ءU��G�B�&c�Щ��*M̼��-�\z�B�ɍP@ҩYcc]v�,��l��1'�B��9%�<�؅
����1��%>C�ɿ-�ԕ�eO�dVb�C%U�_��|�x�"Smv�k��ߚEr<�Q�۩�y�� HW����t��2MS1�~��'a 4(P�S߆�� �rf�qB"O��
v�u*I�&:s�YK�"O\!@e g�,$�aeB;q��
Ot6M��n��aXt.��M6�S��.{p!�և�2��ˑY,�UQ/��]!�D�fL�Qy�h�'D6
@��T�!�@/c0|�@/�4�`s��S�!�$��H�0�x���1r�8��#�E��'�ў�>q�$k�9d�|5l�f�P�*�}�<9U-��t�2Q��G�$i�Q��M�<��K�y;8��H�-s9iP �Ȧ���V�}Svj��gT���+RAK���8V�I'�$�z�ʇ��1��)��Zp�Bo�/f ���kзt�=Dzr�~rv��8u�Ւ�m'RR؃tb��<ICcƙj��I3��5=�ڃ+"D�8b����:G���#
E�D��w��<�	�l3✫4n-N��} b�ǼTB�4���D?��k߁��qpd�=�\{�IL�<I���)�8i�LҶL=(��	�K�<Y@�٥!=��P��;��}���D�<	 +Ã%��Y��L�|��zsDv�<�VKޠ��3퉞��<��M�<	6�5s�@4�え�y�BtB�n�K�<I��']B4P��"�?M@L�1L�a�<��f^t��X:���9m�Bp���w�<A�H#�4m�Ŧ��r�qA�l@w�<�P�ɤH�`�7fÛ���Ei�<ACͯ4�@���J�r��a�y�<A�\d���r-ݰt�N�;�DQ�<��:�u� k^L�uZX�<�2�Bz�5cWɑ�#�fU�6a�U�<i��̓X�L���˴t/XJb��u����?��� ?&���!KH4g ��2s�<QdO�5 ����19&�)��d�<ydΛ�0��̛Te�)qG���K^b�<���=d���&��/w���A�b�<Y��=z8C�Z
 m� Y�ox�'�Q?%c�+"K�\��(ĽKB��55D�4s� Qj��B��m�l�ʴ���	�a�|1�`��#���V��G^���d.}�Ƨ@x�q�gJ��N�N�ɐ*A��yrMB�-���c�YR�9���yR�|Q$,��/D�$1`�N�y���D��P���<4ޭ�ǡG�G�ўx���O[>	{����_>�Kf�_�z����'HL0�Ǜ@D��2��~�H�O0���&2\<����Sq�$@��D �%z!�D��,�~�idOZ��z�eE.9m铨hO�,�z�U��l�I�[�E�陕�����(O�'E�EP2o� '	V��Á$,ؘ�ȓm.��R��Q�o6����H��S'�ȓD\h��kG	@�HpfH�^dL���6B�ÑD�9@��� @'ˊ��ȓ�i
��0�>�c(���Y��S�? �<�#J�3(H�Q�#�3�~���"OȘ���=;�L(�сX�N�~��"O��S�G��:���G�1S��0�'"O��1 �k���7���t�S"O\a���j�6��fD'ی� �"O�  eAʨ�����R]0T�"O��aw�\*D��؅��5N8Y�"O��c"�K�A��1�@#V/D ��"OԨA��E�7��2tb)"*�y��"O�5� 
�>P� `pbɱH� x�"O9�,��"� �V�L ��ex#"O6e(��� z���!�@\p�B��"Op Dǎ�~8�@���$"O� )6�DJ��=Ӡ,�/7D���"O�M�hK�4T��r���:Jx"�;�"O��+����R��R���%fĲD�$"Oz�����'gچ쓣h�'�|�"O�\��aK'd�e(G�;7>�Qg"O�P#ǟ l�>hS�h�_��%i�"Oh#5
DRH"&�Kv��pH!"O�py��D+XH��lH���h��"Of�1�Ȍ�h��iLP2Gf�y�"O��5Eԉ[���q
ߎY���7"O8����W-?I�1��T#O&)1�"O�B̓*m��Z L��E0����"O��8��3�$1˓KX�2�p�*�"O�� �О3�U	��K� к�hT"O�5�f⃹vx��FKZ�Q�x:�"On�C^n����ŨK�x����b"O�)`��P�:.2}Xs韫n��u�4"OX�A��v�R�0G�ߒb~��p%"O�=�V�@�B� 	�f�6
��a"OX�
!��j���@�ӢRx;�"OT�c$ �P��4-�6e�$���"O�0���)ߺm0'�2I�і"O�<z���8e�bm���jo`=�q"O�L��Y����%�	@o��T"Oİh�mR%so�#e��q�Х�g"OX�`,N�>>K$q*�+��6����m=���l7k�:�dnϱ$��ȓZAȝ0e�z;�$Täf�$*�p��z8��K% haXaĹe�4Նȓt����@�$kd�q�t�E�w蔆�1C~��C���л�r�܄�x��5X��o9�`��&4-�ȓ3J����-�)3�� ��8E�)��k�2������|̬�`�*_1[+؅�ȓS�%�d,�AR����˯>t֥��T0�yTDS;4����Fʗ��ȓ>�����
T�|!HJ���ȓJO��궅�� ���qc�Նȓ<>�1 a�6L��r�.��Ge�0��P+|���ٝ+&]jG�ҬI$��ȓu~n=(�B���؆
�5AB�ȓqLE1�⎳p�4D�7ѮX�F���T¹��U�bx��\�k�<���0 �m���gp0;ac&䅄�_|Dy���0B]��&� �9縍��C�� 3Tơ
Q"@P��*`�rD�ȓ9�,A��2k
qJ�o���ȓvv=ʦ����и�a@JtU��m�,�(vd�E�rW�9kh	k�"O�ha�?����=N���"Ox�0�j��Q�Q��/�PCH��t"O� ����*���x�Z��](.�`�rQ"OB��� �P�I��k/v�4�"O���,?>J�B��JuB��"O��o����0{wi�BA�q"Oв4kH�^!x�{��:"�}9r"O���B\!v�`� .Y�@
ڕZ�"O�\�ħ�'mڽx���b��@"O*u�U&!��V"��rGءx"O��˖(�u@�H�$�Ͻdf`Dy�*O���ګ���%���|���'b�����<$𱁡��f*ݐ�' ũE�X�����O��i.�ԣ�'��h�G���-����-Z	�z�'c��q&�EB�X;����`���	�'&���UdpuPcꌤeØ!�'^��Xw�ϟ|Yj����V�p�H���'���ѝ*�2,���D�a�����'~D�cpf�|X,��% �;V�V�9�'��(���}&��p�.]hY��'���Ru�сK�h�	�#@ ��P�
�'6� �!@�@�@���D-q�'��%/���L�نi��U�D�c�'6"AR�W��b�dޭI�ց��'M!JCa�#)��e0��Ӽxb�p�'}�Y�e�Ӳb��K��·s���'�y�%OܝY��P1e�K�AZ���'�B�`��;�`)e����J�'�r%���2<�}ٗ�&����'R�����e?&��7n[��ڡ+�'�:Y�r�J�4����5ܸR���
�'��9ᧅ?]�,�eB�E�|Ւ	�'c:@憁�J�N�Eǅ�
��0#�'�<x�ՈU�G� EN�>
�
e��'d1
��L�Im�����(��*�'��h�����HS� '˻f9��
�'9�-��$[>0h�4��BV�P���a
�'?��d�U?9��qQfǄ ]��'�B`HvN_��:�)��ضv�D���'Π�����-}. �����"r�'[�%YQ(K/[3���'fLx�i�'9~Iea��[�}��ჂY�Vh��'�<�a��*D��z��g�`��
�'�\�HW�զ:6�@wi�
e��
�'X���F��bV$�J��đ`s%�	�'�*�[V	�i- `%C�R9@���'y y
4�	�Z����#Y�G/vz�'�fy2�J�j�Z�{�O>C���s	�'�8�"�@fK���F!�AW�M��'#���h�?6����![�&�4	�'`���a�00)\Ȃg R)$�X���'�<8 ጟ)&^�*�\�ۯ�yi�>H{L@��UK�q�����yb��bN��ӢW��"�yrk�hh�I��G���&�pׯ��yb�U�?��GmƔn�l<�G���y�[2f�,�Ц�n�:���چ�y��)�.�r�m#��+�E��y�)�W�2�q��d��R����yM�!P���Ѐ�¨�1)^*�y"gQ�TPbEZ�d�2/�L��k�'�y�F2x�ɋ!J��1�l���薄�y�b�����c�y��q#Q��yr��R1�)�����zU��p��F��y�gS���ǆ�#R��#��Ŧ�y
�  �1� �I�@���-n�U"O�)�3ݛXŨU�'�BQz.yb"Oy:�i�V1-k�⟸0oP��D"Oz���K*o+~l3�9ĺ@��"O����&.E~<rS�١p؆q�"O�5qD,+���e��0hb"O��*ӳ->�40�jӫ	o��{�"Oey�J?�J��jR�S�ѫ�"ON������d^���ũ��>4Ҭ"O�!)��@/�n�[�H̄Z<�ܠ�"O< (��cF��M�}9���!"Obȳb�ez�PS3l�<l�zP��"O
��`�7V�� ��[���%"O�%�	������k�lu
�"O����*Yw�D@ �{ڠ��"Ov]"%�x�V�(�OʌvњUR"O�\Cf!Q�
*�۶��S����"O�(&����� TQ#R@��"O$0�vm�4ߜ�"�(ҡ:A~yr�"O
H�d(�+e�� �C��<���`0"O��*�G&��Uٗf�	8rL(I7"O��Y�Ǜl�̚�e	"�r�[t"O�p �U�G��i���1�� @"O� ��/���lCW�n��"OX�5C�([�Ԩ�5+�P���"O94��64�Հ	+?;�p��"O
Xȣ���[?`���Qt"O�d0�C�
;U�0D�3j�g"OI�� Z
1�%�P/�"O�Ұ-R!z/nDڀ/VQ�z��"O4E#����u�^��b�V?]��[#"O��Г�����g�"vs^ݚ�"O�X"#���
��c�*}?T#%"OL���B�)�T�q��?K7�� �"Ojx�7jGq�-�� 04ِ"Or��v��1M���5�1k+L��C"OL5�5A܍��	���(�,0��"O����vM�<�6�[�&���"O��9��5�J�rc�3�v�i�"OL@[�ϒ)Q�OV;W�b5i1"Or�x�LE�a"�$�� �8�"O:[!���e��$���5Wʼ���"O����"�7V��i��+{�2` �"Op��g��R��xU�C('?B��F"O 1D��+l�Hpc얰o.b�3"OB�*7��[�$�U�C	[�Ш%"O�-
���(z��	2&���T�9�d"Op|#���,���Kt.	�:=Ӓ"Op}:��'I��E��k}����"On�B�oF$Uq�,`"��0 y���"O譸�cɥ.���ӗ,уFQ��+�"Ov�SR&��qzf��UNG�I�ݑ�"O
 �4�>~���:��L,t��"O,JB&ΉM5��"E�t@�"Op�9���b.6��E4.����"O���S�!�e����"��"E"Ob4���
�X.΄�a'0&�3"Ot�9��]�N���G�O3s���0F"O��t�ܐ D'-��}��"Otdפ%�<@PE���e��\��"O:�6ʈ�xDLy�.�p��˖"O�h4Ռ
�fDl4'��D"O^L!��ў#���jP��Ivz�x"Ox��W��Y���!��%rV�Ż�"O� ���HJ,mE��1�1odp�a�"OL�ZF��+4��)�↊f`��ҷ*O<��v�?�)�Ύ<ap�`�'�r����+i!�]��V��R8c�'��JC)�79�rp��=kⴝ2�'��4s"��\��E!�3]�Z%��'�r%�k�#Z��ԣ��g�L#�'���"��)t�āDg��d8Ph��'ȄA�2�_QJ�[�*R�0��A��'Â8R��0 ��T5*�~�Z�+�';<�[S
F�%_p=fD�Ie@Y��'���Y�I�UI"�;B$�L�����'��As�-ƺ7�"\㡩^KN��q�'�����͚�_O�	�q��$~Q�'���@4l�3MC�ظp�ԅ��@�'�I�p)[Ka@ �Y�Ҟ��'��`7��k�J�{�L�,dlH�'?�����^"r&~�t�Y�s1Q�' �D࡯Q"@�<1���E4a�q:�'K�q�#��6��*�ʔ;w8,��'�����F�@}t��ck�]���	�'_B�i��F$+V��g�Q�]`�'�
Y��U�_"�(Xs�=P���
�'r�2��Ԧs��i��<�0]@�'�T�aC�R0C!rݨ�K �~�����'�<Ș@��:c�J��b��$�y	�'� �+�f��Z�IPb�����'�t�R�5"�LR�k�ɑF�*D�X"�L%�xP�`�:��F$D�|9���=�R�8��{��D�f.D���&r�x&��08<��RC:D��2�b#r��[�HI+{��9):D�t�3.Ř\�4�����6XS���GF9D�)�ԧb�:m3P`Ƴ]8��ȰF2D���$��k�V���@�O�p()��0D�cG�4q���C��qiZ;B2D�(�֦P��� ����X���,D��#��9rEH0�Sl^�B��#�$/D�Pa�CZ�d2�s���(7����4�-D�\a���bC LH����j9�����9D���ŋ�(.@^���eօkJ��CJ"D����Cc�E���� �8��>D��H�$"]ɤ%�EaWP���,0D���D��Jh�'� �;�/D�� W!��
�}�ӊKcy2��9D�|�@Ɋ�{�b���*�G/6e��4D�h�lɳZ�Xٴ��.�a�W?D�L*���,B���gi�<__�\�u�/D��cv��7�LL
�-��0��lǊ,D��r+ܭ
���"� P�����(D�Ltc�&{@�����-^�◣:D�8[�-^��0[�&I�7���ٲ�-D�P��cY,0J-إ(A9D���*D�LK�B*/Z|�%ۉO_�e8F�'D��� �Gz���μE ��%D���N���5QыL �HE�V$D��p7掑d;����ʪ��$�F�"D��!"Ck� L�7#Jlv��j&5D�̂1��j�<4Bg��!F:���>D�(;h�#)�]��H'_��A�j=D�p ���?^^P�qk�$͈���6D��1G�r��5Ã�U�3�b0j62D�`a&	�X.V��״kV���,0D�<���� ��#t��,S��/D�� B�1��Ɗ@�.�(5�[��(�Q"O���2AրVƈA��I�}.��أ"O�X��Q�/d��ì_Â�s"O�Y��L�95��{T�ږI��EK�"O���V���p��A���
�>� V"O�������*�سI"��S"O¹a�Çu�]��/2~!�M"O�t
ug�+�и���vh�"O� �ƌ�q��|�&��|-:8I "O.tp\�_�p��EN�R*챠"ON�z�&�P����ıA��Y#��,D� !����@�b@l08�d�=D�|B�Ԗ?J�8�l%X��H(�J!D��rAD�>$r�Kg��_Z�n�r�<���=0DJ%ۃG�;4�iC� e�<����2�A���3�r	�s
Y�<��d�-���`��S:>��"�HS�<�$�Dy�@��"�B!L/�P��c�L�<YqN�pj��B ;���t
�L�<���3d��0#@�B�	�2��"�I�<�c ��AA���矴yp���qk�E�<��e�RZ�h��N/q�bU��g��<Yv� �ƅI����0�MD�`�<	aDQn�J�ص��K����f�W�<�L�1�~TyG�.2Q��U�<!3�0"��)��	�-���0`�CT�<��W�н)C"څE�,��Fe�<�J�.M�0�$O�LS
����Xa�<1�R'7V�뇄�:cM���D�f�<�7�צ@����(� C�IHa��c�<����N_,�a�LWL�[�.�W�<���	.~�	Ň��X�C��S�<1�KL6�t�Wh	v����ҥX�<��?���a��Əf��ؓ�EDT�<���X�^,ڄK�"y<����R�<�BM�jSn��D�s�� @Q�<y��d΀���o���8��U�<��O�YRBD{s/�b: ��%^U�<��'�� �dٗ4���%[�<��b� 
�aBW	G!��B�OY�<y�!T�Va0�1BP5Bb̉��) X�<��A]#k^�*֫���[Q���j�<) ��#1�z8�F�%8�����!Za�<i�A��ciZdk��i8�-A�a�<Ѣ�,�nКP�Կ�؀ȱ̗e�<�w)<8hsR�	�J���A�F`�<I0Ǖ,�9�U��%L�I8g��u�<�T�^����q #8f0�S�H�r�<`���]��EFB��Au�x�<�(�d3��"��Ș&�Y���u�<�VmS���3��?g��%�Clp�<��AE8_��)����=e��@�F�o�<Iѭ	w6�y2C+�<K垍�Li�<Q����TB�RF'Ō��T ���e�<	�J�. >h�k2Bڏ	�|�C"�P`�<It��@��KX�}���C�j�Z�<���ݷ$���ԣN�Yg 5P���R�<�≎JN(��kK�PV��~JrB�	��f�:�`I�zM�v$�06�B�I��p��R�GRɳ$H�5H�C��T�����4�P����/4NhB䉐# yr"(0�(A#%l���4B�ɘF�t���.գHn�\
��1N�PB�I&~t��D�	�ۚd�q3v��B�)� �c�m	�1N��I5�@�(�%"ON�:�cB�6��QQ-�H�h��"O��%��h�"����k�l	�e"Or=C
�.l��MsA�xx�P"On}PRj�RV��a����Q�O/�yR�Ps��c�,	,b��bЩ��yb�ĉ@i� E/^��Ӗ#�L�<�&�\ t���Q��2t��Pk�o�c�<Yw�UY�mh�&ظQ�^k��Ke�<A��X�D T���b��x���G/�y�<� #F�8��xԩI� R�!�4c�x�<)p�Ǣ%n@Qj�۫&+n�CQ��w�<�J��0�4�h�'ox��r�	NH�<��AH�+Y�Q�"��z���r��^�<��,�^;�jD�:���91�NE�<��ɐe$�I'ǃZ�`8�
�A�<����̰��QӲmQ��r�<	�&C�L��L8R�2Vx�EEBq�<��ǍH?`Dh��ؙE��A��Io�<�r�c�As��\nb��ul��<�Q`
;:I'.���ʘ�A�w�<9qJ�뮩!�YB��"�nJK�<�$/U%_.r��nۋ/�ub &EI�<	U(D4"(�AS�F�NxhA��B�<�W��)0f�{V�V�<��5��lw�<�IԄM;���&��TU��14Vu�<�!+cF�@CVC��w� i�ÍRs�<���э9�T�#�V�,P�vǍh�<Y�кo#�|��$Mv����.�`�<�ѭ^Q��HZ��\� �J��v�	q�<Qi��)���#'h��d��kF�o�<A�k�-wyx��t�\�w-UT�<	�(A�K�R\��O�
J�-�w�XY�<�f���'�x�� �>M2Ha!RN�<��4�L��K� ���L�^�<!Gϕ ��i���[�d�d���DX�<�s�P�~�hd{0҅�@Y�a�V�<9�AR"�>10׆GhyDmS@��n�<��ȪArI�@��L�V�Ym�<Y�C�[��!�q�s�<�wj�N�<a'Y3Q����3�4����M�M�<�Q΂ ʠ\�"�6�"y)Kq�<�a*���b�q�X�pv�����ȓg�H5 d`J�)$<H���t�X�ȓ���k��<H2T\�@�\��ȓ-\쁲�@:��Y�b L�I������Ȳ�DQ=<�@2`�y��l�ȓ?�D�1�!�����4��ذ�ȓ!_��2��U1GZt�#듻e�z��t����ۛjOF�*���}�Ѝ��<[�h#��	�h�f���wÄȆȓa ��X�JZ�:avԩ�m��hZq�ȓ���kT'YAN���BB�x[��ȓW�Y�a@�
b��+O�b3`��4��D�b(�	�n}{��N��N	�ȓ^5�@X�G�Y���yw6���"z����~�ZR/�6D��i�ȓ_.�A�lGr�
��!�а,0Q��Rc��#v�ݶ$4�9��S��)��o��d� 藉M��x��͕�l��ȓ(�l��+À7�R��cG?f�ȭ��";(��q�C�f�؀"�h8tގ!��g$��(2%]�l� ����1 \��ȓ%,�4k2EU�"yp+��ذ(�<a��S�? �P���L�e�T(�aU�b��D"O��%j��V�akT�k$:�"Oڵ"@W,�z���\�S���"OL��[��@�)�30��˱"O��� �Ī.1�A����8r��a+�"O���03�|9(��p�<�"�"O�CVOź�y`�`���4t"O�=��BRj�4Y{�M7%����"O�9��LG�\9�l�/^�0��"O����[$�ak�Z/p�X��"O�h6��p�BDJ���i���y�"O�D`�N��֜��>�� ��"O:������$/�X��eA�)��u0�"O8ԡ�.ю0�\#@B�-}VҖ"O�xВF÷6���tI�F\��`"O$tud68�.�ȱ�\(օ�F"O��X���-_��;'�8 ���"O.��1#�*4��+���~r�9�`"O }[f.A�&X��ૈ1h�u*�"O�IB$8n�I���Ub`��C"Ob�`�6	��Ysfgܛ(t��"O2l���
�����$"��9SA�TZ�<so�?F�L]�I "z���n�|�<��C�)�U��E2��X��`XC�<�D�4�	2� V������F�<y5��2f%�h��$��ON����(�D�<	2��`hlb���^��#Vh�G�<�g�37� ���ǃ*do�sG�<qa�LF?:���b�L�L���N�<��֍���Q'틅�
��1�L�<�&E�1�"��B
?5 \�#C�FI�<�ҥ��c�`	�h��'�Hh���J^�<�u�G�aQRIQ"�Y�>#��o�<1l�"/���q@���R k�<�,%|��`��d��Pi|�`�C{�<�t%��=�a�Ӣ�4�jгҧN@�<Iǡ��7� �c!��R���z��q�<Yw�R�A� p�� ��$礅����m�<!�Å9U�*%B�ʹS��k�<q��A�>t��:q��L3��ǟ@�<i��0�`	��T�4_�u9�O\|�<Y�-��+e����&\4JK�9F��P�<� �	���I�F۶��a�t�Nu�<��"J��r��vjȝ�N��n�|�<���W4 0�k��H�
u�Ĩ�IN�<���n��`#&��|FZ����d�<)�fUp�ؑP�OO\� ����Pk�<��/o�1pV��_?��な�a�<��4�,!h��^�.:����&�^�<q@�_/>L�I�@N<&E� Y�<0��$E�
���LS8~��QŇ|�<��:�'�.{}�}�&MGx�<�碞90y��*L���_v�<��B�a��mz�aV�s�.Ġ�p�<��gR�-Ř0)�,�	/5TD�cFg�<Yf���;�~e҂����caCc�<qq�x�E8ī��kg�^y�<q��́T��!�J������Cv�<A���HNp� 	��D��!c�F�<�D�1T��z��.R��!bB�L�<9d�H<�R}�������vF�R�<��aɫᲵ�A�^%	�~4�A&�j�<�Gh��B��@�R-���Gp�<�v��6:�z��G�
4SѴ�2�i�<� ���� ����{��Cf��Q�"O��I��^ܘ�ɣ 9Hz8�J "Oz]3#��5�
�����X��"O  ��ɞ�&��x��lI�m�.@��"O��@E��p�q1lA�J��"Ox�3��,�E�7���W����"O ��0�J,��@E�Ĕ���bc"O�X�	ߔĔ�`փ�W�0��f"O´{E�ӱϤ�L��f�x��b"O��𥟅4>��䥟�Z�*���"O6 ����Hu!���/y���[	�'��a�n�b㾙���H�>4�
�'vZ�7�T�"x�0i4&Y�5ư��'{쭂�	��" 
�adH�:O����'7@�h�	��E�f�^��#�'�6�0
X�Xؒ�ȉY��4q�'
>�Ulˢ;�h�G&$�z�A
�'�T���'R
�srK�h�e�'��!4��T!�`Q�%T����
�'n���f*K#y��C�����:�'s���4�N�Y
��D�ͥ�����'�>���6B?|@
W#���2�'>��0�K�W�b��	�t���
�'��ej��ˌ�@���E�hb���'��Q4�?������.h� �x�'!�%�ԈK�&��1��-�p�ؘ�'A�q�Zv\L4Sp���]亵��'�n,��$�E����(T R p���'+ҁ���6 �Bc��532�2	�'�(�c3*]|�s%	{�z�X�'E�3S"�lJ���s���
���'�-)b��;��4�PO�~����'1p�Zg�E��6�+�̆{�x��'7�*����pt���KE�����'�p���ȚS�0�KJ�1
�U�	�'PLhc*ɒzb�b�$S�%H�i�'�h���Lo!�{��lJ����'���`���gt<a�g�7e�y8�';1�'��c��j�d+X+ <�'ʂAJ$a�Vk>��VjެH�H�'�>a�A�C/�1��`�~�8�h
�'z.ݹ�/��c&�d����	Hq�	�'ƴ{6�#'��F*̾E��	�' �ґeֳ1���DkވI�@ Z
�'�f�3���-olz��æ=ux}��'w�`�#I�"j��T F.4�.�#�'�	���֜��RJ��+uzM��'F�i�`*�j,���"�7,��{�'�p�V%B56R���`ㄌ*Z��(�'_J$�ެ!�urp��}��'q�Q�vA�6S^F0PO�.2Vٱ	�'`�]p���r?|ЭX�}%���'�~�q'��-+Y �@Įt��ū�'���0���XM	bU&�?e�4�
�'�@��H�&�E�4MW/d"�c�'h��:A��?P<�S����i�����'�q��m��v, /N���'�¼�q��&�>��B�� @2�a�	�'�l<E�ބ��IAjY�-I����'� 8i��C0j����8wAhI:�'���x`'q�D����j,>e��'�6 �DR�5�T�)/���42�'C�N�?����h��
5B�J�'��x���?�p�Oֹz������� >9b�BՇ!x<$��E�	>h9�"O�Հbg��TV��j�&� �"OTɓKJ.b_�1`e��o��("�"O��)a��|�9��ÕJ��Е"O1���G�-���B�fm��"Oz�����j-��V�2ډ�"OFX���P1
K��Rk˪q�"O"uYF�82�h�kƬ��.� �(e"OB�1�E5u�L�zU2��5"O|8��L\��88��׏Eۂ��C"O<ф��y�Ȫb�E�M�<MBu"O����&K�Z��8��׉b���"O�(d��H���E�(UY
!§"O�1����A���G-M�)�R"O��hܧ]�MK�!*�z "O��8���g[����M1@�C�"OR�G�(b<d
$��x�A�u"O�5YF��%�^��D˟�b�C"O���m�,6�l Bd]���p%"O�����*V>q�A�0���S"O��8�c$��p��@�jY��"O�UaĪO�(06MÝ���c"Ot�0�JуrT�ѓ�
�3��q"O�h2� S�,��b@�&S���r"O���Ū�3,qj�$[���kc"O0yb���>s��aC̈́�E��5"ORA�b�	(y;A��͎�R�d �W"O�rU��j����Q$��"O���e
�&Xz�2V�ֳ(�8"Od`�ƃ� ��͒d�ܯ5:J"OdcV�V/��"'b�n�f�A�"O�H�N�,eC���1*�+ �XͲ7"O,=*E�(xh)1�&ն|2�Q "O\#��[�zg`��C��{:��"O�i��X� �� ��1��=I�"O��S6g�ey�$��C�.T��D�"O��@�'*#�1	�##D�&�;"O�$ӓ�;/�J��%C���<��"O�PJF��q#��Y��Y�(�, 
D"O��SUH��<"}�F���lHQG"O�%�g�Dtpx� �2�Hf"O��'�Ҏ5bN$�fĐ�9� ]{�"O~��s�̦?��$ٖ ؗS��"O��I�`C�k�9�B�����"O�˓��!IQ0l�G.
�ơ{�"O�Aq��X�6I`�jEG�'���"O,$���	3�����+�|�#�"O��Ԣ^��3�%YN�����"O����>48<���C"j�"��"OB�bA���x���q�
J���r"O K�*
tڨs�N�+	
�0��"O�U�炚��\��LU�#��C�"O�p�V�Q�W��lJ2k��)�~x!�"O��P1`�3F��af�@�g7�p�Q"O�=¤ϒBz����(
#3 ��"O��h'T�Dl0��"{�BM��"O�e�Q�T"�la����hbt`��"O@94�^�X��i� l���)f"O��9�� �{�<�
�h�_�i7"O���UfN7/}N G��u"
��U"O������,T����d\):�*9
�"O���R% C((GMV�U��d�"On�0p�e
4\�"�H-2�"O��;�`P�>���c䡆=�(�s"O� V�CC�Аr��p����?μ�"O��p�	7�
���
�V#���"O��P�f�sEh�
�Pl��W"O�y��N,Sі��	^z`R��"O���jͪ&���+��MW�x�p"Ov����| ������&�"On�w��AA��-� :�.�A`"O��Pw@5(Z�Ւq��{ʠ��"O��bG�;1^�`� g��avlz�"O�eA"F�r��iCA��0����"O��I�@/3���#�ml�� g
1D�,��d�1�ncq��3#.T0�.D�h�"�P^:4لC��_���Aĩ*D��C̜!E'�0�&��8��a�uC(D��sք^4ZLjq�6(xK�&D����%L��xQ�Ů����w�?D��Ǜ�T��*K>
���C5#�!�DG$�Č����J"Jy�M��Py�!�/jtы"��Z�Ppav%���y��M�4���f�RfJu�E �yR���^����I��N��}�D#Z8�y2���L
�!T�B����R�ޤ�yb�H�-������\':��(�b����y���UI�� �T?v�� bE��y��¢ 2x�f�D�-��#1�@�y�C��Ye�}�G��.!k>(yP�Æ�y�&^T.�H�ʆ���N�)�ȓGϔ�#&D�<l0�q�W�lØ��ȓA
��iUl� ��@�IT��Ԅȓ!��qq�d�?6������1�,ЄȓJX0щe��?Y��q��^}ƅ�ȓl^��r� /n% �I�J|�ȓi���)vjZ� ���rCA�[�pń�����U��"�`A�cG>*T�ȓ,+��sIۀ0�Dm����1\.����|	��Q�rȒE��jV|��ȓ?V4%Pc-F��:y h�/T@�ȓS�	c��.l��	��*v�=�ȓ3��L�Q��5��Ńo[������B;-�Q(G"J P�;�蘟���|�dMj��W������C> �a�� 圔��C܀�Z�rvk�P��ņȓ'��*�*�
�fhrΉ� �u��-<��e��lh�K ���1�0���)U&H0��`9�a��ۧy��ȅȓq��i�E�� �a��	`
-��U���:�o�8��J�'��~��ԅȓ,0v��b%X�(S&9��*	U���ȓB&�09W��>2�z�A#וNIȄ�ȓ � �����J��uy C�^�"��ȓ\ª��_����^�&,��c-L!��כ.,���8�����^����S��.P$hXD+[=k�(]�ȓArp�QO� @ D�A-�C=���99�H�Xl���K��;Lr�t��9:�ʆ�F>��"�� m��Cڠ��X�Z|��B�_
ȥpP1D�ts�HD(��zA*B�	�p���o-D�t��fó|t�Y�*��+"^���-'D��i���!��� Gݒ �T���%D� �0�/7�H�Xpm���IՎ D�@Jء��ݣ����,� �1D�adH�%!1�I�w�01��jS�0T�ȠB�
6\܎�3���#)�@�5"O� ,�r��of*hY�M�!c�*���"O��p �;v��*�+O�9�V��"O}���z�h�+D��:��A�"O�<�6��o�$#:l���G"O�����W6Br��X1�»9Z��S�"O��۰O��l,me��/{W����"O�P�q���G�9���}=X�yg"O�ɒ5�Ȇ13�1d�86���"OF] �莾6s�<�WL�).� h�"O iD�\?2�� �ؼRI�T"OF4�	�j��$!-�=,J ��"O($J��T &�,���?r����"Ox��d"v��X�%�,d���*OH���Y7W  �bII�_4��';��GPxn��bO�0�V�8�'��u� +Ӊ�rm�!���2�+�'rN� �t7��H�.h���'��H�D�&�N�q��/W�|�'�6HB@$�)^zt���ٶVPՙ�'�&8��a���V+G�!�2���'����,� �P�JF_:���
�'��pi��3ņT
6��C��l�	�'ɺ��7���9�Q�"���6ԉX
�'V0c@�#3r�,z)�##�\��'Z��J��ܒku�<i3nʍ�
L��'�ZIz��J@�銢��*dw<��
�'����ǹ 8(%�$�?-?h��'���7o(h�Z�
7�C�"�(��'Hd��u-�3@����ѣ��1��'IP!�3L0.k��b@�l���':�aY�Ñ4��"'�3��1P
�'W�� tH�������J2��	�'��k�O�v�{�%R -��TQ
�'1t-٧�ZqLv��@�'�v�+
�'���E�� �<����Uۂѱ�'�A�֣_�ebI���ӥ=���c�'|����iN�,�Bɚ�E�.����'�`d�"�	r�@� ��Ϻ9}4i{�'�$m Wk_96������2����
�'B,��Wg�.�~	�2��. ����'�~lz#T ��E��K��o����'��Ƀf�*O�vH��ů_����'v�T�!�V�JI`��i̦n(����'�J��8c̈́ �%`�����'��0Ң�)#Z`
�.�s.	i�'Ŧ� ��ނ
*d���!ª��
�'�� b��\�=f��Ԃ�#|_2�h
�'h��$�Ԫu�2=1kԥ{	���'&ҡծ�#�tҦ�)AD��!�'j*���ڵM��ͩ��K$����
�'�rT�p�>X0�	�J�x�
�'�q0� �,c�.\3/� n��	�'Y�����H����0�ǐj���	�'�.ŋ#��190q:A(�)cP$) �'�T�S@&+�`S�]~��Q�'. 4�`HI���8�&˺A����vk���$��U��ZQ
B�@�(t���"`鑫K� EP�X�bL���ȓ9�<�+V�S,�t��g�ןv(�e�ȓ7(�i`�Ş.p�������U���ȓ#��H���Q7��4�A
�0�.��ȓw�n嫒���P��@��9����4��Sh�7�<�g��}����ȓ��h�e�&
��'�[��8��S�? ̜��D`������zv�\*"O:huǒ&*���3k��`6"Od�� o���`�*�I�1T���"On1���ʬ#�Jy�I I%�"Ob�c�C!x��Y�&h�{>�ӑ"O����U��K�<*�u��,��yR�߭4	T��G���2q� h��y�&T�b��I����(��)�,��y�E�,x�1�$���0�+ i��yRǟ$`J�D2w��=0���6Y+�yB	W:f"r��C�.� �׎�y�F^;-�j��Ň�#�d�:U@��y���
Nҙ�e&�&T|i3�g ��y�i�����Q�mn��4�C>�y��a�T%�����:���d$³�yB)�^5v�0gZ1 ��4���yO�`��Ӣ��Z�j]JdK���y�E_J�ܭ;�ΕS��14i޹�y��N<s>�9bk>EZ
Q�#�=�yR��
tp�4r�V�7t��C@`�
�y�e�)e� q�W�5���`���y����@_5���S�ED���œ1�yyo	�V��'t�1jG�W��y�B� }��
p�� �����n��y�W<��Y1��:h�0X�k�y��]>�E�c�\6��!@���y�`XE��S�U�"����fO+�yb��Z�;F�[%9LI����y�JQ�(�,M�U��aB�10K�)�yB.7	Eޡ�cM
R�~u��]�y��̥�R������D��hЦH��y�Ćb��	ehK�E����4aK��ye\�[�����ĠF8�`0��˓�y2"� qn�2&f@�8N|�o�2�y��;"*JMAkj	�͝It��ȓ5X�Ea�t:��歜�l�
��ȓ)��R�ϊ�t���$h�3{J�Ȇ�A:�����O��3h�S\4��/�(: �ї"\����iT"6Q����9�*\�DJ�<�`�h�e�3�4�ȓ]".�K�F�#&���c�?��0��Xv\�b�
6Ι��㎵Y�Ąȓ+.� ��5֮<�7n._pnu�ȓwVN��B� 9�@8HbJ�2NꘇȓA��]Y �¯d5�u��@J=r��ԇȓт��+�a�)���E3�t��ȓ�,E(O�;��)վ|�px��/: Ṓ�>Vh`H� @�Z��i��
U
qх!_�V4RTx�`Y�<���ȓ=�*A "E��DjE2I��p��ȓ_�LVB>3��ܻg(UqۦL��~6(�g���c�34l�WCN��ȓ8�}�6�ikZ`�v끅I���ȓ�6�
���<y���s�e�.H2��H�kf$T9_�X'���n�ȓo���J�c��M�֨0�n�E�����p��yB�Ta�Y�7��5#ŰL�ȓ0XD�r�H�h�F RKE��(��P�Ű��>ഉTY:�����N�
P�Vh�%��)T�	h����ȓe�����AHMd)���>,���ȓ}���g	�Mn
�c̾W/^T��f��ڷ&_�H�v�1�ꗼ}��fd���BE�R���yP��&T��S�? hd�ƬY�OR�E1�#C�¥��"Ox5�,�+�8H)AD�fr��"O�t��k�1���6F��sfX�"O`]�2��9��P��֩'qpAp "O�X��G.@	�HK`o��!`��"O�5�W�[0L�y N��QL�qd"O*�A��0*�,Y��F,D?��"OLQ�-�s�B�{@�ƱP	�D� "O E�D��&[l\9�CS����"OB}��mS�=�� �B�k���"O�Y��C�-Ij$i�l]�u��q�"O�j���B�� &aS�/��a(�"Oؔ�E+P�T��B�I'Ң<�"OZ����k}���u*Ю\���s"O�����lX	���ژ̛�"OZp(F�İ3~ +��;q9���"O�h &솁&'���I_�2�@E�"OvE���m��]�DB-m��!��"O2"�#E�MYz����*?�
��d"O|h���P�h�k�.çj�XI�"O��a�+�C+ty��Aerq;t"O�Ȳ�@��`gxD�q#(F)s"OT}jVJP81��s�U{>DHh�"O� �0�ڔ;��AA�a���s�"O ��KW���1��OU���T"O�����a�䁒�LM)]W���$"O�����=�p��H�?�̹0"O��R�M�kִ�YKU�@C4�z�"O&]��X2�Q��jI�%��I�"OZi�+&F�H��S� !�|�6"O8ԓG�¶Y���RS�&j$�sw"Oj��Q�8θИvg�\�|���"O-�J�)fÀ$Zt^uI@�/fB!�$E3-��G	�RJ��I»�!�DM��|� Ǫ��ELdSH�?N�!�JY���Q�1�h3�Ǌ�+�!�$׃^��]y�j�8��0��Ɓ-!�d6Q'8��C��t@�(��%�!�D�)�v)�m(8{�E�b�S�u�!�dG3:��rgL�zt��A3G<Gf!� �c�>=���6U�t[P��7ER!��T+�*$c1��7���Ve�!�dVX����n�!&|���0�̜3�!���J�L�j$�A�$���AB�.�!�䀈s|�8���^��`�1�B''6!���6,,CU��+}��cH&!�$��:	���͑NdTpqBj�6T$!�DE�(�aJa��!;0��0�_�K�!�C�^n�ɥ�Pz�VP)b��Mk!�`�h�Yu(�7W��1��aN5%~!��8M*�D3C�R�0��c�X%t!��� � M�Æ�8(|��b�@@�!\!�$�G�JX� ��5\r4;�/��Q!��[�]E��+5o�,<��6L!���>]�㨋�B��W��l�"O2h�q_!,�B��@�>z"���"O����0,Q
26PZ�
U"O�<�.�'�>|��Ɖ"C��"O꩓r&�f���3� Z��&"O1�m�2����U��R�`"O���D�	OZ	�Ê�D��;"O��QrE*wWf8�׏J�aǘ ��"OD�"Bl�5����/͇$L�B�"O`��b��/��X!N� ��
U"O� �i�������ӐN�-_o��KS"O¤H�D�48qr�*C�\dty�6"O��roJ�8lTU@C�"O:��㕫"��X5\�e����"Op���,�($���c���R̀1��"O�Y�E)�5<���I�B�2�"�`b"O�%��a��z�����L.��e"O^M����"GGn,V.ҹm���"O@t��(7���	cGJe���P�"O|�󢆀��Ts�9d��!�"Ol�)o"���e[�ko����"O�p�$I�7��17bL�9l��H�"O
�)�g�@�f˱ˇ~�|A�#"Oni�B��88���3t���i�)�P"O(=�J�P�xq�v`O�J���"O�I��	5�h�Qq�5cF�\P�<���	t�"	�o�0vfn�L�<�wF�;O���%� ʈY�XL�<���P�:��⢁�=�rX)�m�s�<!�f"���I�(�8Q-*qq�(�E�<	����Y2H�N��+6�KI�<1B�. YX�g˥�j��a+�E�<���׳7<�EgL͞J��%��w�<!&��i+R�iR� .XQ���GX����IJ�	  CDX��*��p��#�jV�B�ɡj(\��xK�\����6h�B��*%��%:�!ْ�0����YDl����3�*lD�}��._E���&���!�Ēm��C�%��T�Aah^��!�|U����	��V�h��}�!��]�2�1��T��Z��#��x�!�R  8�D�� 
�$���U�!�X�!Ũ�
1"#�h1`�
�S��	Y���qb' �!?x���*�H)МR��5D���Gӟ.Mr�"���&D�	���5�	q��$ag���*��̛%:Y�~���)5��O��O���i1J�Z�V�x�%�M�!�Z�6в��.^�r���e�1Q�џh����M!�(��ͺ"|xʇN�g�!�Dق<�T ��c� ���e���jn����ل�)Tά���8U]�sE5�B�I���f��(<������9��C�	����r��W����a�
���C�I�ܱ�&�Ƣ|�L�kf����C�ɨ  �Z0�V�j�,�I cK&�Tc�4E{J|J�mE�v!ta8Մ]�Q��@e�<y�Z-8m9UO�|Q�r W�<�#�I)ZԱ�jE�*���ӂ�Q�<�Ԭ�% =h��ѪM]JT��˦����d+�S�Ӟd�Dl�b"B�tU>��!L2)�DB�I�YB6@P�`(Z��"�RB�	6>6a!"`	���}X@�F����4�	�/K���B�ܥ��	���7m'��f���01�3��4��H0�8�O���0�f�	�)NN��A�TX@ن�.��t��Ǌ�o(\ReDW�B� e��ki��8��n�n`�!�C�J|�i��j�f�z�D�$s���EJ��&�(�ȓ%��1��2b� ��+5��F~��~b�-�ŧ����ጎ9+R�C�ɧn䊦��	$��)��Ə�x�B䉺
�P<��ܰwIJ(�B��B�I4�j����%t$�dLC�,A��3L<!�����LǢ-
�ִDG�H(bJ��R�!�� �!2�摫&Z��R�)\�~a��"O�Ȱ��B}��݈��\!?�H��&��t}��9O�Ic�G�!�����.¹؄"O�\�#l���Qs�HZ$6��&��Wx��� ���3&[#.� ��֨/�On�er�㒤��>���"B�9��YfO@�f� ��JN�A��q{�"O��� -�<�8��F�Z� �
-I�'��0�ӧơA�Аxsi�>a�����4�S����:���#
4|?�Ĩ����On��d��3�6�ʀ�/b��4R֯�Ö�'�$啧�g���	��M�G��� �X�+���ȓ\����B�3)�>T�H��Rd���=�2��Ǌ"+��� ?�����M�>B��E{���	3�(vJT3�(۬8i,�i��5�S��y�1[���`�N�D���+�Z��y�M�t��0�eɔ3l�0R�-�'�y"l�%Jn�q�O�:Y+b�M��y���;���²&�I�@� ��ԃ�y�`�1p�c�DGҘ�ˋ'�HO��ĵ���J��%t:�+`�_�@����ȗ{�<�G@�<ѨX[5 �X�>%���HO�<A�h�mF(�[��S=g�60H�iX��hO?�	%X��˴�C�#�z�MضN�����鉭u? �P6:5�i�R̟O"8C�@�h�p�P�l��CQ���
C�I�|�<<xU��v��	�(�̆t�'�IR�)�'\���s��=l�HP��:`�h��%Fօũ��~N�� G$	7k�~Յ�>�=�g`S�=_�m��([�cGP���Ic��"U,���zB�*B/
+\��i����Pk^2D�A���?(b��=D�X@�q�� �H�ar�s�i D�t��aC;b�ٚ���,�xe�� LO�M��{�V/�>���!�xDq�S,�(O��Gz*����3@�*c��t�s�cl�:��4\O�,��D=A��ɱ�@�*�n����v�'���~�	%b҈-�e��]�Q3DB܌4�C�I�z.�1� �
&q��T�sN��.Y�"<��r�T���&Q�Woz�)%�1~,em��xr�ġ_��)��a��&�� #c����=� �B�����;K�P�O�	8U!�Ԭ'��-⠍��<8:�ڵ���?�!��جQtشK��:�#�!�D5���QC�v "KыSd���)��y{Sk
�$U�VNܩI*m�@!,�d4�O�آbg l��b!�� '.$��"O���/*N��P�H�Y���M44�Јa#V8a�]9�ϔP�6Բ��&ړ�y��S�7���t	Ť{�8�p@�*�@B�I+tk���QTFj&��ꟐT5�=G{��9O��$DbV�3�H[j�P���"O����#׬1&(��%@�%�rt�w"O��c�I1?L�0@��s��H�"O���4���4�6�8��#:���s�'�W�8҆.�Ni�Жo=!����ȓ�6���K�&
:@�u�Ͷb�����J���*��A+D��9!�׮??P����s�t[G��?�56a����Xr+$D�d%,�/0UJa�b�K#�ɩQL'�!���DT%,҄д��;�6$BPb�}!��R��X� P�.�P��CA�:W�'=ўb?Q�b�G�!n�"�g�"��[�4LO�`t#��m�@�ږ Єd��P��B(D�� 8!t�ތBx��J�ǅ&=� ��$L��M��'zt8g%�\�V8���@�P���� ���y���vX�ٱ�ny����ȓ.d��y�#8M��	���Ts��ȓsw
49BH �w璠8pU��0�cv祟`�OZӧ�g}"1g��,�OUVY���8�y2�N�~f��C[�U$A�DH׉�yb'\:lH�ۅ��a �R�,��y��%��"|Z��3�� �d`�"KU�9iu��7�'�ў�|*���*'ET��f�h�jLk��B�<)��J
��%�sd]�cR{�<!��ޗ
�@L@�k܆���E������?1��Dw�F0�(���`� �aF.ɶ-�B�/2�Pl)���uE�J�.ElܦB��	"��1`W◟<���!�A�$ԢB�	�T�R},Ш�!�EI�T�b�<�yh6� �&Q�y�K^$�C�I�טYJ E��D�~�
�(܌MU�C�I��v�睙 f�̉��:PC�	�+>�<����.�T8{�ؘu6C�Ɍ�.%��ˀUJ��� �v� #<y���?53��	�uR�J�-@��`�3D������T���{b��/2��F6D��� �<LL��P�_�!
Zm@U*OT�(���U��a#!@A�3���P"O���b]�A�D\pao�#/�"O���C�`�v.��,'��{�"OL�:�NYS�)a�-ɂ5�n�Ad"OfM����A_:�P��~��H`"OD���!�`@`�4u�e��"OzxO
�HK0=�SI�X�Z|�"O��g���x��ܸ�'�9�V�""OD������l��fЮ�@u"O"��Ua^�O����Q�ɒH�p���"O⬁傀-M�������/�Dؤ"OU�0k�7����I"O�D�aC	����b�\!r�n�ɧ"O�)1o�R|<�+U�t#�Mb�"O���pE��m=9H��� =�H��"O�h�qaZ�1Y�Ua�D��v��"O��gmN�c�
���g�<�j�"O��H$F�lfX@�sf��N�(��%"O ���5,v�qP��!S|j��"O*\S ��/i�0��D 1S:G"O*I�V� LD�qU��e@���
�'~0�z@#���L3PH�h�'jL;�B���i)E�Z�:�	�'�����P�&��`�C�Ch��
�'�H��D��!a@�Ct�M���,i	�'��	��/�u�2���[�<x���'�" 3�eH���#���F���'g<�tb��}�rD�2B�
V�	�'���``ʇ�Z���.�Ψ*
�'���6��w��|
Qe�)C��C
�'��-a4�$�y���#��ɳ	�'�<��A ױB."{��
�D�
�'\�����	|L�F%>a\$���&~����AI�"��a	J�PEl��ȓt��I��f�>�p�q��
E\a�ȓi��hjF�
�a9��af��ocPA��)�t
�H
=��iR� �\1,Y��v{��aDA6!D�3���a��Ȅ�:	`)�!(G�IK�OBZ���zqB�������8 'Vo��D��S�? ����ʂX���aG�pt���'"O�Pgp�Z�����4KhxXy�"O̝�e��%OCP��H>]S��;B"O��²-�"�f�!%d�63�����"O�w%ˁ v�Q`2��~��Ѕ"O���f��_�21H�F�	�JayP"O0M��g��3G�lX�d�p��	�B"O����K�4�8� �E=��T"O6����#�-��bL�`�ڭ�f"OV(���U3d<������f�{
���ˬM��X�#�0I[qbtԶ���1��0�O��j���ڐl����_��D�W����S1��`�ԅȓ>1����$@z�z#
���@��I�t`�������I3���C�+���@MS� �lB䉕�4�(�mل@&�Z�j� ��e��C
�*0U��F�'�'Mpl��C� 6U�>�aăCZ$�A���?h������*���3�����Ό���D�N)PY�=+�' ���Q��?O1���OP�Ī�6	�
��G��$�|�GW�F���Au�� ��,��i�_Ǆ2��c
EA�����p���� I����0�O�����d~�"�mc��8	��L.:��iC.O��+��H�1��s�-��"��Y���1N�<�;u�D{�.E�.�8��m2,(��_�E`��R�N�`�j�&3p�qXq�Q�0�@��D��pAb�G��>
I@�4Q�D�x�J6�S�N3�ѱ�!5+¶MѦV�c���񄊆JҢ(��AEY��飛'&F��dԭz�&�^�Qc��+�ՌFJɲw���b���@��:��� �	�S2*0�G�ֺZS���A��q�r�u��+ţ�1k�Ř$�ƅ��'o����*�^�(�)G�X[R���!��J�F!X�>�A���_U���	ߓXI�PC3fޚ)�8��s��0��%O70e졑�9D�@@�NJ�YJ�L��.� �꓄�0�(���M�F��6e��j�B�+��@�6x���L�L�&îL�����n�<��'L�j$ز$�A.=`�y�F�>{�� ��B-K�����ٴ��' |���N�v3�A׻
�.؇ችv�"��pCY"��u8$��П���S�Zd��iS��YG�=L*�e�E�\�zAyUKN0z��'��':н0���q�H�@��"&~����O
�
����@A��AM�;��������8���UK��m����$��-@MB�kN�^��1�i��N .����zo6��ʏ�:�6.�o��m�gf�Y����c�r��f��${k:�ʎ�>	�q&�ǋk��ҝ	q�����������ϗ^!�$R�t𰃡�*}&:��t��-1�4�����J����ӘN���"C��m-�����y.4��T�(�ӱD�N\�E휾N٢�A�G�~�xR��p�*E˂pY���O�5آ��X*�p�@ܟ]��r��[.��钕���n���5�̡EJ�1Ȃ�Y.X(Q��H�d�5=��a0)[�(�`��x� ��8T6h���
�*�h!���8 i�#Ń�X�<˱�	�`wv�{�%P�!�4�;�����5F�8fZ��'.���V�j�`8ж&�9M����"K,l����IFonX���x���v.Q�k�d0��fչN�Չ��n�6L�I�Wm���6d�@mnyh�)C��f���=����D�ʼ#kNpIF�SR�R��c��>O��#��D�d�6A	��<����T���"hJtA&NS�P��Ɔ<a�U���R�/^�I�K�.4�z��E�y� ��������]=��Q�QO�d�( �2�֏^d�����'��HLB�)rb��5��?z��q�ѯ f�.0�bG�\`��[iٟB�d����S�`�:�.W�'���VCލ��!3vIٺq�����L��V�f�Ѳ&��k�1�Ҡ��tHz�-ܦɒB�M7gY ��C^J��Ѫ�ō�(&���A��]�K֎���*��4�9��>�F���R�p�)M�q��U�$h@@�*��	�h�дy� ^���*'`�&�JYB��A�H���Yb�L�v
&p� KT$y����'2���%S�h9�zv�):(:�:��	�VR$M��� b�6���Ӯ=��!����l0�=2�*);+0�jA�QIHY�GE"�@ X��6��ݣ��z���«Z� 8�!�Gɴ���CU���Epb�7s�d�@��O2T�o��%.�i#�ȷ�������aSЂY�B�D�`Y�ze��a^�Y"������fK
�4�2�LU�vE~Y� ��W��C���E�VW�B	��Eh`�(����@<nٜ����6���e�ɧ��ۿ08�Հ�
�v��� �Ь|Ѿ�oZ<�u�u�S6~	=�]��K����
ǩ<���G�Z=UPĨf�Y����v�6"X�2�%�l��A�H�k`�l3
˓��ax���s��iؐ�J�4�BhJ�o[#�ldz�ڄ	���ac)&R�ex�hǦw��Y�`(�6�LpJ����'�|h▤`��y�@E�&k޽4�'5�*�)C�3�x�i�b<�����	�0Jm8�)�À�W�8��dШ�\9�DƂD>h��Á:J
���I԰M`,�qd�S�*4�Q*	�PAbr�E/M},��[�s�^p�:}B�Ƕz�����4JO���)�F�r|��Q�C:m�d�	v�
�A<-�Sg�L�(nc�))2��!�w�T�2��r�ֽBS�]=/�sO>Y ���p�d�%��ð ��:��@g͆XЎ��A�k�6Mԁ�f$��.m���0�E@�%�T!��.�#��)�#.�3f)��$aU"��8Ar��P@ǮF\)�0fe�'��$*� V��#�;����<)�4�''q9���C�I�9�������2}r\�P'#O<=̀��	#��gGňt0�{�	I}��T¦��"&:��B  ?F���Ez��ͿM|8I��$���z5 �i�-Y���#V�ۅ�Y�Wq�	ЀQU�X�{�E=Zg�5%�i�)r�
Y
zJ��'�1%��t;�_�$����2gY�< �\s�O�W�q*Bk'?�֊T��09���W|P� {�O���PEiQ�'�b��BǙ1Y�8]`��ʉc�����
QP�5OS�5O��LL!^{>�@E��X�>Qp��?��	�
)+��Ы�&���h��'U�iA��X��1mC�:�RPiB%^�*F��G�zDo�G(�v�(@��w��!K@��\�V��DEӏ'��8�L���l=���OP8�8�'��)Spቻd@�xu�5P�4uI�)��*�K�SH�}SE�҂P��б�HZ঍�Q�	�l��Ir :�Yt&������V��)Y���iݟؑ�	��jj���	���'�<ҵR8:&�k��ӯP���XU"�)*G�)`ō2V
QEm�'�6�H���� �
!#���ɲc�QR��0 �
h�*��|��HBy6�Ňʱ ؁���Ys~��a�S����b�T1��hΤ ���)�;q04sfI.8�eC,�ҕ�l�{���0X>��G��[dF�����Q��\��VH��y��ʩr�졣�_����#�-R����H9L�} �b<�j��J�s��˧�~ºi��(�k3���J�.Y�$=�A߂R�Xh��A��Z��E��x�	h%+� ��'�`�4S�}X���0=��B�<��q��v9S�@"3y��
�<�(��� ���� #f��5+[���JU(O������'Mt〡)��(W��Gx�JP�a4��iϘ:��1#��,h��1�l��/����7�ٜv�����S���O:{����l�/z`��y%��"(�G(���	�|��V�V�/5���V*�0��]l��M��og򁨢���&�Z��Dc<cd��ׁ�x�u1��Dg;��c�&ظt���`gYE�J�1v#�?��`휄=ư"�"��vdL�N�����>������K*eO�ٴ�ڑ����ON/o���}�7�N�5RHbF��Nך���2�i��-x �*�擶"��}�K�d씁2���f.qbk;�əJ؊�Q�/Ҧg �xS���M�0�Aq�6E*� N�R�Y��߁S��9W��%a�D3QA�D�1X��t�$�t-�D��\Zr*��`�p	��דM݀�x��M%��'2�Z�iH+A�i��d�]M2}�,,�R���>��+����P1T�ꢂ�"�>��S�߻gV�cգ�-* ��	�J��ÚϿ�fAP�ʮ`���\G��t	f~b�G��l��I�I�"��퓙r���9`�0��|�� 7���A�lNo�1� +��i��i3��?�) &�1��T�v���4�����h�21h�)��<
�c۾q0���Q���`��I#19��K�#)��Ӷ�!�x��e���8:�L
+M�iy��Kl:rA�ࡋ f:ڔ�r䜔d<����C���Ox���كb'������+=�y��k!j�p���δ���O2-8Җ~*���7j}fI�̳�ZCe҆3��+_w;z�0�H�wV,}  1�g
8j����$�b�ZP���?���	K J��2�4�"��*%J�څ�"��(��h#l�=�Ft�$�O'Z���͵7�$��缃օ�
\5�h�W)
i�Z�La~��R���KlE�Fװ�H��	=��)����e��m�@�!����JY�L�I� ���d��BR�](2�~����	#,H�iͻ$=��# V�!��@�H��H	RC��<f���q ]�tD+�St,}��$J�X�sx�� ���z4����ɥ��A����i��㝼��|����Z�'t�Y�pCI�{�r)Y��/-̈́䣁���2�Ȁ��דW�<�Γ�r,���}�f)��+�����G�8��`���\�<�@�;�I��� *��j��(O4� /A�>�Y��.��,���ݑC7�Ya�#Q�x��dǒJ��;zⰥ�\Bd��aݓF;��1�CǡT�p�����'/:H6!�F�E�l���#��"��Ňm�Ƹ;ጂ<�ȟ��yn��P]� ��J\U�\o�#�,1����4�%E�66��擓Q^�@Qn�[X�tK�?��I�N�.H�1�ю4&��RN�$IqO�x9����5VڍaB�H�Ƭ52���.+���#O�
殉x��!���2�8D0���Λ�μFz�툚�ԉ����?U"l�Z��Qʊ� /]�O���'��q�`�8���'�D�\m�Lxa�0	��ӑ��>�P��B�\��`��Y<�����O�'�>�p� ^��l ��O��z��D>�y�!�JD�S"�i������=
�(`�0)��pO,����t>Գ�*Å�����D-6�"u�'(�O��P��f�dІ�N�IqAOG:��զ>�'Oj�.S��Yz�o��[�,tkb��&�Vq ��_$�M+�kӆhI�̕O�*��GOܯN�)"7O�I�TB�$v��l�/Դx��H"�\zw���F��p���sXq��f�M�q]�U�$�R�LԕI��5���Xu��(�"�� �Dy��斜�� P��$8�Q�L�����9�Ȁ��f�/^������>Ht�3͍�YfuآeKx���4.y��yek�#_�d��O|mZi$��B�EK�/�)�!.�o��i�vBX*E]��,._߮kG�!*�5����c����a�
0�t��
��L�|�����MS!�X.S�XM�r�)�$L1\�F��|�v�d�1©R�[����$�6o���� ��)U�j�Bի��<@2E�@�2�ӠD�F�Kr�:��}@��	���'?��ͭ! a��	�x����#�jô}YդR�0\�Wh��1R�V�[�UJ 0�&x��.��H" @P�N�1°斢:Ң�q/��h�����U�oh!��lb=�@�$/JrX���@�'v� ��D�?
m�q�B�']R�1�'�#=O^����*@jl�u"�D7�>�0`��	s����	5E5�%�6O�A���\�D���mX�q�|<p�ȋB�𐶫	b2�A獆�3Z�hqN�h�`�@�cKw�n0��"sr\�+�S��OERl�ǄM2���I1�&K:��<>�3#�K�J�`���șm��@AR�5.���4ɇ�l��8�E��%c�|#*��<v�i9��"Z5����3����ߔG_*�g�'�Ҽ dG��=��ȅĄi�t��ӊ̈Ez^ �CI@�Zf^h���8� 0$'aR3��5X���A%����r��tx�	X#R�Bm�"�)K�P�3(	��')��}2vj�ޤy�/��qܚ�ÑK�#
�,�'oӲ��'˕:k��ѐ�M�e���-ۮ}�H�æ,_�X����
j٦� <Q��(f�ޤ@�8�i;�T�4s�F�q���ٰ_���U�ҡB�½kɌH���	�T�
�̓Z e��'n%\�(����&n� �ebД�6`�V�
�L�Rb��_)}!��C�m"R��Ԙ
P�d��ʥg�ج`5���aC����O,5��)M %SrO.w$��ץS�WaL����$��D���<!��T6�0�p��˭�L ��HSlByc�k�q���a�D�,�F��~B��i#�|Pg!��=d� RP�T��a��\"H��ɠ �hy��@�rl����9c�,r M��V��S.,���E������n�$0�$#Fb��U�y衋�T�XU�1���ܰ"�Ydq�n\���"}ԬX2�$"M��рK�	8�獋�5N����Φ� ���%C��mٴ�I E�4�a˖� Dr�o�0���c��$���������H9I���\�fH !l�>��(D��GCe���po^^�p�p� �����勾#�&ĉ5列ph1�,zZ��{�l��[U�\��瑂��֝/�����WT,���T�y��<���RT���a!�By� �J^X�"#�D��UC�!5���tE��4�NLp!`��a @��@@��sS��8C� T��&�j	$�YD�N92-\�#�
�'fL���D��+��A�P��;7�"2n��2��͓�<7�PP�A�� ]A�9p &U8}�>�(c
D~ ��� oH�Ç�S�4�Fd��GǂZ����R��7������&:�hZ��J�(��� ��	˲�q�CH&����r��Ĕ���ԋ+��0��!��J S�/J�t�"
I�J>�p�K�6�6ܡd��� �����^,;S�c���q�٠qp�(��F*�c�$�)54�2WGK�d|q�=L(�B�{���'N����;y�Dؚ�Ц&}N����:K�ɓ���K=]"2'EM�Ҵ�c��?�Z�.�>1�SbD%Lk��Q�޼N'f)r�H H:�Q��¡Yb��ר[�e� �pc���C>�\Js�XF�Ԝ �7D�i ���XZF��NZ�9�=��:GER,�e��"�(A�ك|�Ȅ+��lm	!NH9lF� v =6���Ip!�	3Ů$@�"�Z��ɩw� I2�R�0 ���J8̈�*�o�%�n�I%� kF��3��#����J�ib��s��� _��a���#LR�p�Vf�:E�x)�u ��i�?t���Z�����}J�M��F���&��uj@�A����䝇b�HI��ӉX��!a�>|I�]��Fla�,��[� �� ��n��$Ҁ�a+P�����#u�Q"fM��@�H�'Ě[��<F{�(~�6�b���bT�D�I3��#f�,Q%�U�0�ŞC,��2Vi&�"☔aB�I��y���ר�Y�C��o�ZI�0��c0�����e�'y������*��@L��QPV��^=[NjM�R%Ge�����9aJ�ɋ�d��+Vr av�@����s���hA�"Gd����K�y���ĩo[�)(��rB��'�0��䝡-���a,2�D��a���@)��
�B	S���үˍ?�����PM�0ʒ��8*����C�C�
A#�d�!)1�E'�|b!�� d,d�R@�p�ER��'P�ɺ���cv(Ҋwtq��=#$)E�:�^\Q��Ўf"|�i���ZL�A���4��0�"S�H���4M�ayrl�(%$N@	0bۼ� ��&%��uL��Bb�DT�����s�t�NL)`��>�4�ض�K�vL��Jb��-D@����[{����e@�"�!��;�2쀣%P�PT1�0�o�C0��Z�a��<��Qg:�Xt9Έ�n���x'��ȇȓA�\�B!�[�$�>��U�ր#�-����u���@��<�3��	vn��!�݂
b4�3�X1A�!��i8��❻����aD�]���r�&�|,ԩc!�O֙:���60��2�Q�\$	���'1��đ^ �'�`I���)��=p�慕>	�]��'�Z��ψ�n�h{�ˉ�:DԊ�{�d[ hA�ᓨ*
��P�Y#V�~p����!d|(C�	 #:�b��ȡ�8H��A05xnC�%�V�#��P
rR�ڇ�¯FFzC�I�
 yؐa?�pd����k�&C������%gM6#�nY��O�':(pC�I��h �f
8�p��w�s@hC�I�h�p����E�6�~��PC�&� C�I��"SR�:�4�� �1�C�	�_t����[((�Tk�C��B��yJ�l��E�:x���+P��B�ɬRD4a����\:��aVBܗG��B䉟f�@�QM�� l���� �FB�I;E�Y;5N gg(ī�_��B�ɡB?�"$'�DrVh�+p4�C�ɄB�c� X�~1#ǒO�C� k��E��I�j����E�/h�C��<v�:��gGX#2�ا� KV�C�	4&���bL�s[8��td�8/�lC�I?,	����Y"(��A"��XdnC�I-v�li��D�d*�d*�Ϙq�C�	7Z����C�:��\����
h��C��;~n�� �ݝ>z�
A�65�C�	�<�jm˓)ʝfY"��*�zC�Ɏ`W��RΛ�3Fm(A�)	�B�ɌF�nZ�!��0�>����W�+�B�)� � ٱI�J�4CT(���F"O�9
��P+���"��F�1Rt�w"O�� ���-X��3�K�5l��YY�"O¹��#6b��a#L(�m�͏t�<q��E�(Ma���	{RX�3�p�<y)5T�5
 ��1x�L�m�<EL�?s������կ �aQ�i�<�7Gʠ
rH��R�ݤ|�F�;WmN\�<9cÂC���7A��q�}��k�_�<��H�}��0����8$.��*V@�<�3�ʵT��`0��=F(����-[C�<y  X"$�b�˻����w��y�<1WA�T*���j	�"�x�3��Z}�<� �'uA��� �L/~�%�r��t�<����K�z	���(_��T��q�<	� �qYp2t*���'έO��C�I�x�t��m�$aIT��Ck�+�JC䉝U�\yxc��'|�x�8�*f��������!��;��� �K���*�ɉ"
��Ф�-3�!�ܷ:0l��gN�<`���d 剟,n>5���U"JK��0����&n"x0�([� ����� ͱa���Ȯ~�z5H�Ox0��nBP�Pr�o��~GL�'+G�z� �	��g��i�'d��s����'���jG/�2h�0��)�96��O>	�i�7��ת9�S�=�V%�n��&��-9�hX���7Έ\p��Y�/�p�����'nn ��NS�	hF���-��l��5Q�FF.�0!�'�����䙛���`�U�rYKs�[�xK��!~>�!�NQdt�Ba��Z4�C�I?x��@F�*]	�_�Iډ�e�Cl�aA�r�)uo��!������M� 6Ġ��ʸטO׼ɘ�,ز)R|�j�m��	Ǔa�r�pqW�y<x�A��f�`���i�21���$	�Q�I�c�����O�~���	2@�Yʆ��'�5*RG���DP�r.$ZO&���OL���\�L��d(S�^�DG蒟�@H�I�6CH&P��&J='���
Ĕ������C�Le��+R/�)BBH��D�M8<�@%��i�䉶FO�z�E�Â�vS���jm�P�G [�O?,� ��آd���vF�}��.��\�9хkJ#S<L�s$P!�d_^�Q"!G>0xIT�݇
�ё6Ě��Y00ÔCK�I� [�lI�eR��\�4 dad�=�)зM�~A!T�Ʀ@	���
�I�ax�kJ 9>"uh2��k^^X�6�'�����A
��ʑ#ʌa-L��%i؃z%й .Q�1��@���)<���L�:@�iV��oV&u*���P�G�/J�B���W���'L�\ �bOK��db�i	8&������Fִ��(�$s���[2�X��=�f�S�oQb��A�z6�����h}.��v��(�?�Wc�+���F�S�lVr�Z A~=��� ,P��܄�4�Ab�`��/�G<	6��	O��r'e�Ib`9�$�Zibţp$I*rYP��$�@�PL�=���=D��"�EJg h1M~JI�<��(���%&�ح ��x��"����"O.����ɼ@5b��\�cnJ��l�ȟt+$��1Ai��+��T	0��4��l6@7f��<ʓ,�l�O"c�ZM��̆m,, �O�����V@hV�-B��YT�+������e3\|����E�B�j�,�=���`8_n�@�OD�7�P��d^�)�Z�LQi�i�c��"W@�1����1=��9�ڇ8�3O��zAL�0D{L����Nb�V�]+@ ��nYDܪ<K���&��
ABL��~F�h�xa;d��0@�t/��f��\��	W�@@�,��I�Bf	I�i�~i3dĎ1 D��ڠ�~B눣_�d�H�̛-�\xR���p=1�&�6��dԭ!�p�eI�/G+��2:��cqD� I�xu�W��?\=󱃎�G��kwӌXm� V�t��s��s.���I^7]7�X0�	��8=(Đ㙔dy#?�qG�8L�����6Ű ���p�]bѦ�$��t��e��h^%o��B�a�HvT�P��'
��AZ�fH�&���{B O;t�5�d�Ʌ6bli��������aH>�A�˚�}�`�y0�8іxrf�C5��u��h�}ֽ���$c�i�@Y���#�`%
�m�@^l�d�KH~����Y�{m~,��(�,����#P�q�w���������0��EYyjn� ��+�� �O��^���V��V��JpY%,T(��.�O��qc��f��1��j0D��т'��֙Q�ݑ/��0d._�~�U`���e��%�BJJ3B���G��ε��\�!""5�2�_�7�:B"4p�(�F~2��z�.� �����������p�H��|����"ko�tKE��)I�f�L>�(��f�5Q���
1dЯg�`���I����zК]u�p-J�f�*4����G���n,A��\%��:EH����;�P�2T̴Vm>�+4!U_����A��\'&xQ�-�L��0��	��������C0�����':Y8t ڧu\Ȱ1�F(�6��	QG�YG�M�'gjТ(S�[�]0t��&pTڀQ�ƀ-�:��)ф@�l���)[	~];�dP#d�.On-�5M�CX�h����9߾�Q�͝� h w�҈-���������+�w�&��B�X>J��ex�oM��@@�k�(����4n���� YU�y��e�Q�L<6�(�e�>���zj�M�Uj֢j���za�5o=D��G��'[�vⶪ�1��(�i$~�P�[�ȕ�O�LKPJ�3��q�w)�?�L��ԏ�3 ��h��%�T�'�t2�P6]�H�Cw�(��`��b_%7�}�%��?ut�
�h�֦勴FX�j��� U�钫D<Ob���ဉM�.�A0�^H��/�O���σ)���ep��}E|�)K\D@d�͚.�
��@.ɰp��0 �$D�Ҽ�2JQ��#Wo�PNN`��(���I�u�� �DĆ@*�e�I�zܵ{��mHk��&n�"=Q��Ѽ
�ΑcCψ�"�9@ٴn?��hsˈ��F)`ނq�����6���LU�a>���4�r�ӱ��a5��0�>?�8���G8n8��6'��O�r=Y�Ᏺ:/�Ms����b��`~D��VJ%��,�'5�<�s"\6RB*��fG\{�0�P�?M���� ��7A3�)��g͂0P�㔯��	e�xÜ�x�8�@ӟ�T �[ �y¬>� I���q�bD�L�-à��@�ҥ ��'���D��܋B�
<�M�d�w��M �k#6���BHm&@�̘�\3�!�ȓL�\��F�$Ê5��ߘQ�,9�t+�In "<)iͅ0�j�*V�۷xϸ�Br�اĄ�Z�N*g�I�׬��'s�u"�4Yi��j��k���S�L���ܭS�&�k�Bܮw���F잁=��k )�*��j��d9]�
�!?r|���'{ �l�"�� �r�!��HZ��A2�֦Ձ3�B5@�4 y@�1N,�҅T�<	>dS
��L�O?�L��C�-\\�UY%�V���a��O�T��B/�����F�~f���K�?�:P�޻mx�P燢2.���N�,X�L5�e��,T�nj��>3���un� ^�*���b�Ӄ[��;�y�U-Z�O1�XTlJH����AJ��YҶ��ԣ�&D¬d�įK��q�ul���OX7�4e��ΞCp��!ET�P�pt���G�z���9WJ�Y����J<�4;�W���'��WF��~�B�AS�hD�ؓL�x`(��@.G/*��F�?����s<v���I���T�aV	
>5��Kr�مTÈ����Ĝ4��E�ň="��uE,��O��ᥓ;l-���}H 	���k�1�մ~C�@�C��$w,����^E�gD	�=/@|
���?jW���+�7yN�h�3E$���H��a@#NڃZX<X�!��m���"�P�d�*��5���>	`�Yk��D%Å7�L26�T�������i[(l(��@�f�X�
Ш/[$�ve�?G�	�V�\Q�"����� ��*]����.��T�5%*ڰ�%��?=o����M_T��}��fB/(��`8�ը-���`Kʅ8����@����R����tp0��=U�`�Ȫ(� ���}�jʭB���`��#z���v��'I�T����*���g�hr�`i�Dɵ� �ʰk }����M C�`�q����b��"��M�P�ؕ[�.8-Q�k�(Jf��$+5��w0�%V�ig���$�\>��X����*�Z)'M�+R�x��o��tY� �⨔t�j�b%�F�]�<�0W���~���w?^���ԁ�c4��aу�(~-�C��(B	$)J�2FǍ9u|�E��ℋ>�z1�F�Y�Y �׎ }#T��sKV1kx���Հ;w�L���O�~!�6��r)X�����4����d:z F]����M(�l_H0��I�p���1�ź��$�!B�8Çȓ#�.ya��!�.�R�@�O�4�����|Ib�+V�)�(���Oidկ!B�c�D�	$H"���N�+�@�B�$��D4�h�d�O��R�~JA$H9y����Q�^O�lZ!)����H)@�k�� }�pbA�±�#<1��8*�F��gh7$����H�)���0'�6=�	�1(��8��lP��p9��R1%�1�*�!L�	�g��2#�&!#�iQ�|λ���5*�(��/6.���' 0* Ȉ[fH��C�V��>�٤	�u�z�C���l���K��$q�0���V�6���S�t�t�@� �x��!#i޹)P���*�����e�2m�8�@�&���F��"(��`c�i�1	1��mK�i�4�8x�*��D�x�F����H�G
N.��)c�D�j.�<1ql�������I�"<i�@I�*� ��֋]�$�V4�ԄT,3۸E��蒜l��EQ�Ne��"�-�%,�:�vK� �N �d�U�0޶e�2HS�|q�M"u>�Ԛ����R�"֋==[9z�+�w?�Ĳ�LF< �T�*�'��|�D�ֿbˆ�T��.s����N�d�{̉�I�9����#��h����<dĜ<�� [ /q��w�� ���	:���Ā��Y��(H>���MZ��800��l���Ԫ2Վ�y�`Ɲy6�+ �׎<%D�B��G
n����ҹ���*0Ҟ�t���$��;n��e�@��(*�	֠�2�h�֎f�e�c?]K���i���/� l��Kg�vA�
_k2yC4A�bX�cK�5O��5�Ab�cf@��;�����*0a���Е�ȼT����"��`�$ƯO\��	�$�RiP��^�5��
�:Wb�zr�Ԇd��1��H=s64ճr#�&h$ఊ����#w�	<s4<��,ݒ���O�ԡ��=�8Q��M�R��A�i�V����"��I�_9 d-"�T��s��a���wQ?�ؿ^��UQGL�xV��Ȇꁪ=���'�t{���V|rq��x�Oߒ���7�8#���z~J��M�<a�q� n��)2�ON�|G�St��T?;"��`�H�#à�)H�^����ߺJ��@6��;1|��l��Qx�>7�]'Urc7��]���pB-�8� )�Y�d��eo&�`6-G�!��(c�,�=��<9�k��]�bh*�(�.>���%bP,f�j����� �z�����W���dK�����Mr"o���@�ҤJAb�1��	�&���G�	�{�\I����D9��ӟ��!IJ,y�)�RD��04�p�觟�K0,�#���єx�`�-D6b>�H�B[%/j���zyb�1we$?ɧ��=*����K
Td�����|�գuŔ�L���Kƈ�@�=������9� ��$[m�T%Í�	@��!��7t�!��L�3s3؜k� Tg�`.�6"��'Q7p��`��n@����ʮ~�j��,M�u���y��ƝK����	H��bsg
%7�m�b�Q�Xi:|�1�<0~�h����4.�Y��&����3��=�Y�B�qݩ��zd�`Ʉƚ�C����SNT�x3��d:�0<�D�ןv������V�$���Q3 +غ��q 
i&�i	�L�z��M(�8���_�%���1�OD�@%ɵ��IN?��bLx�3�Da�)_P��'~�t� h̓0�8 	%؍8"�zb'���X#7Z��`	� "�!VBܒ4X֭���N��A0��B��?A��x �Lqk�p��3ғ]ʺ���*E~��ש��&�j�u,ʳz�z����x��$y�(��Y´��G�?����C���
��.BT��wƃ�b������[�0de���U}d80 F��>��O[�<Y��>[���Z���]�`X�.N�P. 싵H(fx������c�� q�A�X���b�FV�]�@���V$��Ղ��e \�ɴ&�<9�Ԛ���1���ͦ4��ő �V���$D�4�¬ۧ�C�^��V�,Ǵ�g�*8��:��r�����ڒYD��!� D�AyG��;K�)���T�=��r�Dږr ����`ړZ�E
�f
Ld
@i��M����d}B@J:*�H�Ə��h�*xsE $7���!��h�J����7�*Yʜ6�0�B�3a�M���t��a[�a�/O�{�/&?� 	yWJ\����|�6�Qf�����ZA���0��DD��u��`��nA�/A�OL�. 
���b�52��$ԟM(�W�s��Daa�/XwJ8D.	,;��i�+ϔ36��g��@��d��_�����4�]/>� ����S�h���E#�=6�-p#�)&&e�f�_�^0�c��3���BR&o���%��5��P/�ZIӠZ��@5��Q3;T�K����BQ)Ց/J���0����
K��hyX)τ�ɖ��7�\P�CiخP�4AGI�=7)y�MD�=���"s�����c��3�H|��	�-Z�i_w|��@���fԨrN �l<m!7cL�3�6��@�+�剌0����`"��1��3���KQ��H3��,$��Q�I�5�k,`�D��e����%��1���:��x)6o�XJ�)��Y�g�Z,kA�ע`�����{���#&j5E�Q���UN�T;����N2����4h? ��%�ȑl̢��q	��2W�-�V�Y���l���~�q�E�'I0��D"�V�Z"�j�.&B �����S�T�Z`�1Y�d�X�D3�4?9��4?����J��e��p"P�9&Z0�r�cI�y�|)�*�&"z�{�e�+22���Ǫ�f��Xz����� �(U��hk�.��=��\IݼZ�^�zU��7E�T�SI4��ٳ��	�_�F��g�7.�n�{�h��6���1�<pX`/4�	ԊЙv��<�&�_ >&�E!�cߚD���!k��9��B[!;���XB\=�@$J ��L�4k@tr#=���c�!E�C.���cIR, @r�jL 4�PZ�
��+�bI��o 1s��0(S� '6�d �b�פ:� c�lݡc`��� ��۵��>�ȩ��"*C�x�.Z&;�и�3eH�\ݪ�v�8�����/H���6��!n�)�mR�kc���R䏯j�qY��	� ���MF8cZ��cF�C����,��r�{&%[ ?h$r$A	����7%|�z����N�fH�(�&gR �H��ț|�& A�$�j}<� OHx��ч��dK�$�v�R�$��`��itZt��l�<haSh��t����焵i�"ĻW�3�ft`^Z�'k��	�(8G6d�tfD�V�4՘צígM���6LfJ@eI�zj*�:V� *<O"t�DES�(��֟@�I�.��܈T!�M�漑r�/#
,�E|ҥ���&8���5Q��uA%7Y������M�ѐ��L�m[�Es��
|x���\*��P�F�X7Q7���O1J�р���lY�A�Ox��7h	*N(���G($	�UK�OR��/�J:�����O%Y����S�U�!C8j+���/��5y�2 ���)��C�H�S�N�U�4#����Pi��Z��`�zA�C�>*�Q0��ގp��P�����@Q��V�v�C��鄫z8ĩ�ce�]}i��lMB�\vd]��&�S�� i����`D�݊A�'2��4���f>�@�#i�**�@K#S	Oъ��OV���J&�M#�#�<X�`���0�^��T�S4[�4h[��H&��d܄?�<U��LH�s#%�F\9���~�I�O����'�8���C	���J���W!\zm:)@j.~���"Oj���N�'2������}�E� MV�z�|p23�O��p�����r��#�fÖ�I�dlJǮM�!�ι@v�����.-��1�c�^>3�
$$g��d��b�<�O�}��C�[:@I��&|���'~>HQ���"'x��'�`MR�OI K�N\����~�Z�
�'�]�r@�/�ؙP֭֫$
V9�{B���u�ᓎw���*ߪu蘽�'(���C�	 �Mj��L�e�@͂��L	=hC�I�G�� 
a+�?�h4a��8H$C�Ʉ~r�۰e�z�N�qcIO�W7DB�ɉH��\ʤ�W���@��>dZfB�	_�p9��.�n�怰u��$<nB䉫i�B�rf2]�01��h,hB�I�m&�b�T5�L���^�{&jB�I�6��e��Iυ�6`A,Z��TB�I�4s���)4�4ؒ���W�\B�	H���K$9�D�`�o*<B�=sV�X�̉-�&�B��$B�I�p�C�B?N�& ť`�hB�	�E�zx�+_.�r%�"OrB�	,,�L� ��d�Ye�
4#>C�	�D�48�gb��-Rr�&k�,C䉖P��E!�*��y��BA@D<5�B�	g� �K�dXM�i�*D
��C�	*�X��`L�(N�T��E�LȦC�I�k���4�ܫE�]��C�	�{�bHh�^2�����	�>��B�)� P��3��p��DĀKй����;2�U)�(8 HF0�$݋`R�$����C�؟g\FyQE�I��dIP��>Ō�q�EԗU%���O� ���B=?�L�xu,ԗ[���yw-�H�(����TW�����0|��Gη$��A��*T���
x�xC�-���?IU�ЎA1HT���#HT�E�Q&H�&LeZ��Q�W�p9�T�ty�IQ�F\ʍ�����E!J�4���p <	s�N�m�X�O>{�(m�q�ʟ�ԓ�+J�A���y��ٟxu��ә����@�3?��%�"|*T�T�{<���t͈�O�������<��cػI֎,�L>�~�)R>�z�"ܬ3���*U��..��)����,7-��2�)��t��o���0|
������uCF
*��K7bL~前(�@'�1t�g�T?A�RɎ>��:�
!;�tU���!��]���T�pJ�ڸx�X��P��(!�܅�O�=Ԣ4�ɑP,��0 Ə`��l����E�7���c���XqO| ��F#����9��;!�	qN!5#ȝq��]1s��"~:�?S�Ћ���ShV�#��8#.:�;�
ç�ʀ�BM6CxH��K�?xPx�O��(O� ����i�Ȅ���G�+*��S댖&�\��n��_�x����R�?��la�'����"_L���DZh���2CaϚ� ��+�N0�,2f��9��<�B.S�ҕS�@�V��Ң-�0Q	�}ӀĪL��ڢI�Y�0'�$/���@��-��b�x�d�'Of�}�U,�̭1K�Rɸ)
@k��ژ'Ⱥ-��f>����cɖ�ҡ��Q��T��/}�c�ӟ���y��$MI�Ip��u�رR����XC}��ퟐj�yJ|����yB
�B��pX��7FN��ը	��	)�eY���	 v��?q��'X��P�O|�!r�V��x���( C����^b���1Q�<����D	}��X�"�}�B9�7��i�!�d
|��Q���¢� Ig��J!!�$��4���n�,�d�
RFb!�䅓i28D��~)�EN������'wl��d��G�Di�n � �F���'�T�9���\%�l�2cG(zL�lR�'�x���L���쩲G���Ġ�'vKw��w�)�f��������'46,���֯o����璻|kz|��'��a�6���#-b��>yȘ�9�'eP��6�W�l�0#�\�pE����'T�r�C��Qc(yb�œb�P��'HT	C���`��%*�d��a&(<!�'����$^=~9,y�Cw~�s
�'��1`���<y���Be�ΎL����'$�٫`k�o�[����2Q٢]8�'�J`�cX`����dPUhx��'��{"i
}SRm��e�M�F���'��E��C[�2���H�CJ��'��\k�&��1��D�EƮ7�*!��'l$�8'c͎qn�����8̢��
�'R�1��sT4�(��[�nM��'�Ƞ����2���c!*ؾ� ĩ�'l``xwb���u�q��O���	�'B���eF�S��36!C5Y���'���˧$�	��A"Fm�(	K��
�'u	C�NľI��a�A�m�T��	�'��U[�ώP�b]�Td�/2U�9�	�'�L����:[��<�u�T#�p�Q
�'�����їzX~�����m4�z�'$�@Aq�� I��xbMߜJ*=��'Q����T�+6P2�.�$���'U����"�<?X��'��6�赒�'9�qV��&:����Jֲ����'�����R�&l����CHc�'NJ$�0��(X:=�#�]���ER�',�w�\/H��� zL�	�'�DHPg��5�4M��*��Q,x�	�'R�=1��:�ꡪ��7E( �R	��� �4��fR�D8�q����~ Z�
�"O x��� �|��)ñ �C"O�H�&�4M>|�5�ɳb<�Ԃ"O��2)�OV*�V�F5e-�(�"O����^&x�V�x��S?� �"O��2 bV>h7�9���X�ޥ("OP���U]H����̕�
�(�"O"u�!ψ�bTL��@��RQM#'"Opa��I�k�4}����;|3x�E"Ol��Z9��
ԡY�"1����z�<�v����̳�oOG(�`��R�<��nU�Lb FP�R�ˠbTT�<�4�H�&s2l�- �;�)Xdm�h�<�mӝY��(��*�R���,U�<i�D�q��sA�ՊH�X@���@�<I��S��1u���"Y"� }�<���c��|���T�|Ң�h��w�<q�^9g�^D�+~��Y�Nv�<Q-Ɇ!p��VGZ�u��͙���K�<��Z ��9寅 �vU�EȎJ�<!'
#F X6�ߢs�����I�<)`-��<9���A�2��d�D�<�fX^�����ޏ6��E��J�}�<	�#�+ݖ�Ĥ�w�b���NU�<i�oװ���i 	 -�A��Z�<�!�'mJ�I�V#MF��^}�<)bi�y��P@�3R�d�� aWq�<��<P��P��O�#�D����o�<�`�Y��D8��{Өd�S�v�<Aq��0�`#�=:���q�<�5,J�j ��r�J�}�<��f��j�<)�E�<M�hP�Q�A4alxu��Hg�<)0e��>���k�:>f4bt`�_�<Q��9�(�עO��RT�<���+0�P� u�J1mFM�<�E]�R�9�c
g�2t�aLE�<q����u��8g�*!��D�VJ�<y�gY��F-H�*:D�0��H�<`Ȉ<	��]r�b�;.?��cƅE�<A����!|`���W[�<qD�B�<��fW�RR���GQ�!<�E:�	A�<1�� _��D�"f�t���0��|�<��k�>$��� ��,q��r�_s�<�rB"�4�R�b�e��u���i�<)���?�*]{� �Vp5��&�d�<A��S9�4+���,��l�w�<�pn�A�h���0\ƞ9�Ŭs�<1��:!��M�a�H��p`�#A�D�<��FV�DC�X�q���6AH3LU}�<qP�t���̼����. O�<1�D
KÀ-��lZ4i�I5o�I�<��H\�#��8S��/OϠ$�^�<i B��t�=reJ׀#��0����Q�<I�/7/�H�Y�eK�V����!�ON�<���ٲx�	)�P
�`C��H�< CR�O��iC���K40��iYD�<�J�JJn<[P@]�(E���VNJC�<��(�T��������M��A�<�e�B6w����vQҀ�`,�-(=�C�	1p�i•B-� �ס��θC�I0^���PP�_h��\qw��WɪC䉹`�F�����IQ���)H�C�ɰd����3~2�����?��C䉅/�F<)e�:f��b�o��B�)� ���]!�
	��W�al��g"OʄXBՉz���0#Q&e9�"O&�rT��.��l���(FC�
D"O>��1�ڦx+Pݢ��_�OG�q"O0�BW��:'��)���*5�4��"O� �����Hhl��c+�(Y�|�#�"O�5`!�� i�$h���I�z��"OF�9`B~TXta�I�!t��� "Ovxz"�Nu��HuKCj���0"O���R%���v$(w���U��"OF��P��è����9x��T�b"O䜡�i�s�b,����;�z 	�"O�)��#�\L����|-9W"O�d�EcM9<u1&���f�H�"O�@S�56���o��>����e"O��8���A�y ��k¢a��"O�S�&Յ�,��q�YYf�0"O`E{ªG�l�v,S�m�i�^�
�"O�H�4�W�*G�`@�J
L�4|��"O~T��ު�R���oU��"O���I:
�8�nZ'\v���"OJ����.1@B7 ۸7�z8�@"Ov쒡�>%�7"�*;m�=�ѧ'D���V%S��Rm�ϑ+b�� �� D���a� Z��z� P�Nä����1D� ӒFL�KDpQA��P}N}P.#D�S�m�%ґ��U�Z~.�Y�O"D��)ԉ�2){���S�Ւw�����?D�T��j� .�j��&j�_�\؈PK"D��aĎ�2=�|�,�7�&8ʒ"D�����ҥ�����i��&�j#"D��RD@�aŞ���LL3[��@s�*D�LSg�^ ��{&�WW3(��$#>D��DkG���'�&pI��':D�ܘ�H�K�M;��]��Q4�4D��3��76��YU��?N�d}h�D3D��uJ��>,5zcΚ�s5v���5D��Z ��*F��	Q��ZN�����7D�īpb؀w����	dB�ı� 7D���AS )��I S��<���#�  D�( �϶2���3 ЍHb*�:�b>D��j׆��e[�����z�� A�/(D���#���VA(s����e�&D���Ùc7nt���1T�ʼ�"`)D��AF�X�ت�O�B�ĤPCA)D�ĩ�G�$t���b�|��'D�����X�a��Y��ʜ-c��<)DD&D���F�/k0�f(Y[���b/D�h�����{����լX�$�x@s��7D���sΎ�2A�`g�҃���q.0D�Pct�R�xX!eDE�����d'<D��0#�͝0�p�+bH^v��-�C�;D����Q&Y���۹I6i�@:D��2���6�,��N�b���R��$D���1×z�4��ĉ8�d 	��"D�,ұ
H�eO��ӉU�\�F@1	"D��2�[��b&^�I�� 'J%D�Pʧ�ĸY�Xa;�'����i�e*8D��xS�@tKJ��g�/Vߦ�J�5D���G%NL�^䪗���S�2Ҋ3D������a�=�t�@(M��}kSb0D���I��pŜ)37�r�N�ڄl:D����W0[/�@�q��)D�t��@9D��2 ���&�iE�LhN�k8D�� ��z�ʒ�* �x�WDb���"OV]#g�SL��}(Gč�=~q˔"O�8��[�$F՛�B�F���+�"O�����0�,�WK��Vꄌ��"O���`�4a�.T�� m�εˑ"O>� &��=d%йP)��t��Lx�"O~�����,n��1N�;\�\�r�"O꼩���Tܔ�2�ҽ�vD��"O~M����6M�֕��E��<��q��"O&4���N!PP���:P�5*OPaPׂ��Z�<�A�H�  ����'��}�!m13����04f8�!�'ybiB�(̓Q���PNHvwr�!
�'�м�b���~L���#��}p�J	�'�NmC�(ǹ�lXH�&�(~���'�,����B~��襈���L\��'7$	�n�sP���OŋpT !�'�h��OиV��)c۾J!$�B�'�=�CM$���C�?�03�'P�
�.�s�\h�ֶ3`��C�'Xʱ�Ȭ?"�LHvΝ�3B���'��6;zg�ɣš��_nN��'�h�0�C��"��$�s!��o�v�x�'��X(s�Nm����̟�t��]�
�':����!߲}mL�X���d��2
�'Ďܺ�hT��sb�.W��9�'��)��,�*18h	"N�+O��T�	�'s� "A�;��m�!A�KyPh��'���8�샘+	ꤱ�+=F#��r�'��5  ���   �  �  �#  b.  �6  B  N  LY  d  =o  y  |�  ��  ؘ  �  C�  8�  ��  ��  ��  P�  ��  ��  �  x�  �  ��  � (
 l � � 6# x) �/  6 C< �B �H 	O �U �\ �b �i np �v !} � �� Ɠ � W� �� � 9� ��  `� u�	����Zv�B�'ld\�0"Iz+�D��g�2T����	#Ĵ�de�8�?Y���y�FJ%L+h�˧�Z�`<�!#�	�kw�=�F!��)X���&Q���S#��(V�N�_�x��H<J0>�	ۙ�Hay%�874��$0s́D	�$	�UYb��;t��a��e&�ݯ;/6�-��'�?���/[ �*�J��X��հ����_����� �J*��d�� �%��F�
6M[�N����O��D�O����|�^	��C�A>P��K�"z�����O����O$˓�?���?����?1�Kκ'L�JT쐎���{$-O�?���?!���?)��?1�O��/Q�<%����.˰#׶�Z�D��Z7�Ȗj�/�+RMk���']�	&�ɫ_JJm�d���_ zU!6F�\1�i���u}�;O �P!�F�0hTF�tm��<�DGԔn�a�N_�Y���!�gǟ���4�?���?i���
����)nލ27`�>)iH)��H�@G���S�O��o��MK��i�X6��O�o� fX)K�4x6Ԁ�)�#H����m�Pu�(I�d��!r\�Y� �F�릧(:x��A��y�^����u�K�Q���(Ń['?��QQ┬?� 䘱i��2<�@�I�$���w�Fhn��?�	�O�z��ƈs��P���0t(P�&ȵXp��3�4ZUF���.� n[25y+4�>̡EeX �5���ib7P���jC�T�[N����Q�OЪa�Գ6�V�����k���ܴDN�v�m�j�"񈇵r��}�V-^�X�~�q��݇$�ȡ3�ʞ^u��C"�G�i�Bx����:��	R���՛ڴ,�K#��\�/�7.��(��i�2����D4D�!��#��d�����
s�X�����0�	�,��5�rerqI�O~��*`G-E�d<kW��"�UPgݫrSlQt��ߟh�I��4�S�?A�dd�5�	QG��������~\̑��R��\e�R��蟬�'��'��I��A������K#W}p$iҊx�v]���Ԟ8�Nl���CPO�	P�`#OP@P���`>:KD4;�U�g(Đ_B�p 
ī\��a�B�����KՂtS�{�å�?�t�i��ʓ���R≠6�� ���޷ �0������	O����$��P�	�|b�Aڛ{��x��E?n,���B��0��4cc�mZ���&;�6er'ȗ4Db���ib)t�����ئ���Iy�O����''6�ya�E�P�����6���{��'�b�ǚ��+��D�W/�40�ji���?;$��� �C���H�X揝r~���]t� K�钠V�� C4���)�&��.�}��3�<GB�5;�Y���
g���'op��`͛�G'ҧ��Tᆙ(_�|y%�֊p�ZY���6��>1�O4���e<GB���.��n��*��	�M;��i�1���r�JSh'�C�@?8����'�[��AC��ٟ��I� �I^y�J�x+�!���J�n����Q+J HM����l�n��%/Y�;Y��V>}���S.�'�y-�O�;�ƟH�|�����Y��l�`��0i^nB����E�|�%��yer�ͻ3����eߦ
�"�A5N�bش'��	�����L�g�ɯ3H�U�R�_�#�b�í�����̕'���>Ah�q��I �ӧU��r�Jy��kӾto�o�i>y��MyBZ�.#����bL�
<�\��n�,r$�ë>����?�(OD�'����T*xI !*�0d����n�N��v�� Ψ�#P�S"��yb�ԙ_hLr�@�:i�J�c�8^����Z
P��U�4��v�i�t �l�ϸ'<��bW#� k�H��uI��1�v��?1Ӽi�j"=��&�2Ć�j`FB����� �Ps��'h��'0t1� �:Ү�q�LǤ0��e�J>�G�i�7m�<�R�Dt���֟�S��[�d������U6a��`[�h�ܟT�ɬ$�FU�I��L�	�E�>C��H�Z�z�H����WKM7�����I�P�\)��B��8��C�-i����T�u,�T3���B��h�bM2x`d5P���"��!G�@xR>�4�M<)&��a�$Dl���\0Q��~���bh¨^C���u'CDyR�'���'3a��N�M�nmI��ֲM�PM�w�����?�w�i�����Љ9��$*WI�>V
30.hӰ�/���
��i���'��5H� ���+�N�����1R4�A���e����I�d���� ����T�����'K�a�i�|b$A�G��Wޣ����F_����*?af��_���f��(��˴��)p{��%.F:g���`��rc4���۽\rj�1|Eͻw����S��O2�n��ħ��O%H��G��E�4)Z	�A�t�K>�����'H1O�0H��ыT�,�Y�fy�DS���G����nϟ܃ܴ0ћ^�M+�i6",�4a�x�#�9�+A�s�6-�Or�@i�II���?����?�,O� ��f��o$A!�F�+�^r�MzL|2��˦��&��Q^`��O���aWe�Y�40��鐦+Ԉ(&�
�Du�ĐTMN��楂R�G�~�*,�D#I��L��!*9��w��h����}T ;�I�5`�脻iۢ��'�@X������?Y���?���#j��l��K�oI8�����?���?A��?i��L��8!�ݱ:�`J��D�ʵ��<y2�i�6m�O8%l��t�S�?A�O��0�ǴXn�t�����^���',L�%�'��' ��~���?���9��౤✁RO~is خ^M��y(� ��/UB]s�9�[G��@��^D��ׂԼ�$@N�3s*�@a�sJ�͋3� �@e��8���Me��L>1��ZE��p"�܅e�J�˴�	�ll��I2"��qx۴�?i)O�1����<ɶ�PfypM����Nd��eʫ��d�O `3�{�i��'-�d�:W��bq���m����J�$����ݴ�?�)OL��i�O@�d�O�Yaᜋ\|,E��϶r�ZE g��O��D7-��D�O���hz��������� ��� �����g���7d݂
��]�q�'}��:���1���Y�ȟ&��Ҷ,BP���F�ǂ�̍�C���.��Ԑ��T5���=�׵b��yӘɔ'֪IƎHG(�5�bĂ7�%���?	�����(���ċ�Vt\tA#�s�����v�'� 7��)i�b����$}� @� K
�w� n�Ay��V��I(�OW��[G�'5���
�P���X�~�8�'�'B�FLhy���Y�F0:��6�f��˧��	d�X�b��3B��a��$?�	�V�K�	�?�h��2OZ����nX�	�XR�I��uW��8]�� 0��^�Rѹ U'��D�	L��/v��@lǟ<�O��<l������Q,�t���v�j�OR�d"��d�E�L�{��'F9(�:��P�4/<�E�k�4o�$�ڴ�?)��/ ���-BQ�h�k���#Z���'�"�']��3�yR�'�B�'^�N�s�*\1�`�4�HdiH�tC�ß*CO�ay��ےop����CwL�h���:�񰥀��z,�6�Ʋ$���a&��\-&�"��U�e"\Ȅn����7-�Wy��B��?�����|���.M����K4g�)�EpXў��"T+��Y� �~|�{�!��|�'U��|��O�)���˓P	��[0툇etP�JE��&> �
1ظ?�6LP��?	���?� �����O��D�T������C9��@7�^�tװ��f�:.�̐�-�B�0�K�'-V�'O�^�Ӎ�*&4�E��M;�|��i߬3��ɑ���^3^ly�e�x�I�0�$�<u�&L!�� �|�q�¤r�xq�4��u�4w����Gx�b4v���o�;�pPH���'az�c�5����)�z�Y�M�����ƀz��]>�`P�i�9O�aY.���� ���=@�z#�'��I۟|���|�<:j�	����&О�2eCI�1֝�Ek؋M":�A�kK�rV�t+c�ɸj���[��w2���N����2��YpfjT\����7G�n�)���_]Ǣ�$�<��M�Or�l���D������B97�bi�.G�K��'�a|���1~L��2��X(�t/��?9�]��6��oͺĩ5�ŗ�t�8�!Sc�v7�<�a����'�R\>���J���V�*4�� Ȑ�<�� PvF� �I$����c��VW�`C�)��u��ΐ9�6$�O��0	C�U�z��-zq��G�r���/rC�u3b.�"?�1�q!�0��Y*�b�=��u�N 8��	:UJE"6Q9�ZU�'q�����;�F�8�'���Ǎ6m��Bq�ڥ=�0������?1���3�M��K�?0&����	M���I�YP�4��'M|�iP	�1,�a ��jҨ����i��'��ϗ<��c�'���'	�2�P@J���X⸸����G�0����DM�q�az$�S9Py�PaFv�a{�����'���Z
ӓ0� �d��<[?��i���8.�BK>Q��X՟4�|�<��"ӓ�e@cA�2���A��RX�<aC�̖!<���@�ӠV��]�&n�WyBM=��|L>9�L^�'��5�RO�$:�d��'�"*�������?���?!��)���O����O����#NF�x����:Njt��˂�tݢd1�`�Rx�`�f_��@����$�f�j�M�#Y���Kc�� �h�1-54��������*%C�)/�\��`^7XuJ=Ps�'ܐ7�צ-�IYy"�'��O��`$%�d��\sऀ�+#��B��OvC�	�B*����1lS.$;��
Nǒ�O�qo��M�)O�p�L��I�	ß����&P�u�4d7q{n=qWn���,�I�%C�A��П\ΧyyX�9�/B[ƵȴhǱ8���i�6,hИb!��>@�p����O|<1�凞|�6���&�#J"�;�]�2�)�j��Bê�:�Κ�t]�6휚<����e���K���'$��X����	K�M�D��w��O��d:LOJ��A���N�E�֣A�DQ�U�'*���G�y�Hrq��	��قz���Xy���yH6��O����|z�%�?�s�U+h�I���ep�pB�.��?�����i��f��a1h2XqV�"N�?��OV!�S��
:^ ��ٺG���O�ys�]�F���gf2>T�ZG� ���r��.pr��闾�r@��Ψ%�,�K�(B���IPKn��Ħ9����r>��1+�$r��!T�ֹ\�j!n0��0|����I̤�f��XB����m�]�'~2Fg�2�lF�	'�8HVŚ�F�`h����#
+ٴ�?�.Oֹ�
���D�O��D�<y�� 䪩/�QxjF?���85�ހ,�rr2�i�i��P=����'��A�E \�+]D�SP�%�n�����o$ ]��c��1}Na����1�
���$$��BX�*�N�9�b؇ʑ%{�-�`�	\��6�yy��?A�����|��SB�A`F�V���W!@*.�2�'s�O�">���3 ��8Ò��&�E0�Ȁu~�i��6�O(mlZr���O��b0�����}�h�"B��6^X����!J������p�I�l����OxmkQ�=\��%�DbP�S8Db��+d� L��I�_iĝ2ۓh���� ��;�=.r���i��Y����6$N��1�S��azRc;���Ja��%������D�|�l���כ�nr�$�$�<�����'1v1g�� W&�,X0��#���s���:�S�iH��K��A��a�D	:�'!f�"jӒʓ�?������O�jGě0Cr�{c	��r�YVl�O���p=����O���ۡu�9 ��?�\XƪU�߁�rF8TV.x���	tJ*��:OJ3ᆍ ��Z���;����M�t<�҈ܦ^��3�m��H�IԠ��
�s�{����?ıi�h�#v���D�ָKh��R%�1h����O֐��'�R�'��QGn��Te��.6���P.O����Şr¯�3nDV �R�LJ�"mr�
�?�.O�YIG�O����O����D�K�G�O���	��L����P	S�J���o�O@��V)(
�1)�^Z�L7���M�-�H�Eb �`������Cܢ+F"��'K���`��m;N���H�faD���Z��k���	�A���p�T8ie�$H���|��ɩq������%(H|����N�g턅�ĝ�5���R�!G�䓥?qK>���̲f�x��CX>L�5 5��5���'��7͆��5$����n�i��HD&��O#���E%���M���?!����y��]9�?)��?���yFK6k��՚�O��I�<Y"EG FR����i��xؗ�JR�4!I~�t&�ڨ3T�
�)w-�u�^>�@;R�	�Z��٘"!Z�ju��K n�5*A�ʧhb�A�f���s�`�;7`\�B���y�v!����M{�R�����Oh��>&���4%�*s��y�e ӿJV�k���F{��IU�`�0�+O)�D�0%r���O��n�<�McJ>�'��.O@���F1X8�a�I+C���
�b�T��~B�X2/'��K!LD=o��� G�i �)H-#��ZEl�YQ�������hH^lGy�ȫ�l�0'��*�PVbU�<fh���D���k���L@�Q8��˞`ذHDy�m�T2��S
Z7�|�{T�!n? ����V�6��O��9�	5f���(��y��A "OR<$��we�S'�n�917�|��y��$�<�$&D�?i���?y�T��$���ޗJ�6��g���?���>kh���?	��̜Ѱ�Ȏyś��ßgϐ�n�"i��y�O��a���*�ax�끡H:���	�\����AѮENfL���0u:a�D4B��� �"�4(�hŒC��ZܓE�b���1�M��^����5�^q�U���xu�\S���O^��O8⟢|z�O["O�l!�N��,~4a�\l��f���8�ߴL��ȣ.X=�x��	[;t|�$�iN�	�*Yp̕'A�P>͊�#����`�-�"|i��A���5�G�P�������T�U��Mۤ@��M{*��I�*�cТ�1.<�#��U�)��'C��K�,�7H��Y�U-Aj,0��˽E����d%�K�r�ݪ}}4H�pGT�\ܥk%��Z���b�\�ɵ�M+�iҚ?A�O�tL�G�6�Z�  D�]��I>1����'<1ORQ��	G%��e̚]��ű4�I��M�iT�Ax�@�ĕ�N*������d�IslX3X��m��,���)ա�qb d����H��۟`�;bWH��Ӈ�	o� �=/�}M<9�ꛗ1L:M~�=����0�̰����XiIq��_iF͘ Ό�u�}�!\#!X<�|�<)��4z���%h�~������M��ib��$a��Y���	>�|);W��+!(&��+mTp�E{R�'Z�%A�(,��l��RZN�j+O��l��MM>i����.O.p@�9�`�a!��@YLe{%I�GZ$٩7��OV���O���������?���5�ܡ�P/��a\=)F��4�H���*���B�'�b���Eͯa&�ī���;=5P�ń�w0|����$Ȫ�C`e���0<�����?*��5A��dɠ)�1�j�6,��#�M�ԾiL]�@�	m�GRP<c�D�������c�켣��xb��<CPxŰ�	N���(�E���>ߛ�}�Z�*�|�`�ia��'�r�Z�	��u�ă63o��y��'��գnR��'o�	C�O�������Dlx��O�;4CϢQ��	0bQ�: ^)2��'*���AB&�b�l��M� ��`��g�����R���� Э��F%B<�K@&Cj�	�=� S�d��L~��Þ>��A��.l�^y؄&�0��	*7u@��6L&80�� |p�������W�opT\!��2/���p0��OJ˓�����?q����x�8����'U���"[E��J�]�0���O�a�c����0��ߣ<����|jϟ`ġSA
R�Xk��Y��@�u���ȕ-Ш6�M��OB��ԀЌ�Y�Х�1�;��ِ\�V�*wD]�{V:�ru��\~"����?	���h���ɺMs&��@���=8�Dځ��D�B������V�V��vp���"Q���?Q��S<c�<;s�_CAQ�A"%T���Od�D�O�0X&��6c��d�O����Ot��$2����� �;/�$ӳ�D*}h��#���5iV�m�L><1F		N�g�$�`c2�_-�� �G��>S䂥r�NH�,}�ٴ˲QӇ�\8ZH~��%R>�ZkR2E��=� ��t )�C����q p�'�ɸ���Od�=�Q��*:����l� pv	�d*=�yr�H>{��;!އZG��K&�?��\�ퟘ�'dD[r�Ɨ,����L
�[d��
�,�<|�"�'��'�Ҍf���	�Dͧ	�j�JK��:Q�0�so� 3W�:���p����C+�`z0b)$�ITL5�g��P�EJ�o��Ш���;F��{���!@8�˅��̢��4�n�/�6��.��'-V��W�Z�{�2��5��#aV��QB���?y��'�� i��Y/��Xٕ!	�	B���ߓ٘'.�yH4��T��8#�	}~Y�L>�Լi�'!�A����~J�eqx1�4�j���@΂�B����?A&�M�?q���4�΁P�t�#��%}����}i��b� �0=ȼh��$�U�c U/|c�Fy2#�	m<f�W��f���&Y�HɄ��ڝU
]���ăq�vi�b���F�~elZ<_�"�O~��`�'����@����7�HYᡎ�+����+��2�OJ�
G6u~L�����������=��|��'�(p��YK0�b�j��A�N�0���$%�Un˟0��w��ʱ*gˑ��}PriT�	wL,y��	��'��Y�3�D�G�����&��*�Z���م	��^>m��h^��f!���"`i0|cg{~b��v����Ȍ�D��Q&б0^���ʀ]�i8�lI��G
�xO�h11l^�{�Id����|�)�'K�T��s,
�'�0a���4{��Ň�dؐsF^mۼ���[�M�"E��1�'l�ޥH@���"rY$�2-��8�޴�?y���?���vL�+���?)��?�w����0ꐣ|�ʰ�� �7#�ȣs͛<����D� 6/&`�R�����	>%�6����D�Dt}1��%�HİT#KIb(��
(T���}%`����i�}Q�\��'b�̸�հѦx`��ϼ+~"Lz �|�gϼ�?!���yr&V���b��rQn���<�y���o*��RT/��k\��C1����B���d�|�(G�s���5�
�G��Y�rR�0������_e��'O2�'���]ڟ���|$���?hxk�-މN��e�5  ep�CO�U�F	�g��k�(�R�Q(�<�O�G}��ʔ@�2҄$ Q�Ze�0�gU�)�s�%dD�h��A�G��<At��	t�<�`�\�/߮�9���(�N��	���?��Î1��p!��a���H�<��םng&���@�vǐ���d�C�$�MK>�pG��L��ϟ���]9l�"ĸ����09a��ٟ��I�9?��IП�'D�����L�f�0��@�M�@�P"|ɒhT904\+��
��M+�/ړ~V�0׬X+:>�s���-5*d���(NI��/��(u�(�b���i�΁�1`�_�'1 ,���?��OLq$/K� �\���'0�\�!g�|��'Z�e���A�\x$Pp���_/��	��o�2�ÒM��d�6���id8KU�N��?,O��t�O��O*˧"jZ����Ep�yB��	�F����O->�t���?���4<C$T��N[6�3f�V�:��+Sd¶��	�
!���a/��̘��H�B��I�e�$@삈�J�2���AW�!��� S��cߟ��`�a:x@p� �
kܼ"������O���S�<uGƱhJ6��/N��ء��QP�<�'�� �r+�-@`�FEȠ-�r�'�~�}��Q,z����"R)���a㮒�M����?Q��!ā�%ŏ �?����?y���y'/ɝ&@r��X�@�j]��M�<���Ђ$�>��m\?w�X�|�<�FӲP�ف5�� 
,��jA���S�@(#�'�b>c�:EH�6(���[s��	'��5�s��O@�M.�����PD{"���n��
E
ҵ$���E'M��!�d�#A7�� ���4����&;=���g���ğܕ'�Ա�Ǉ�m�b���B,g�L���h��d�����'���'��g�������'X�vEbk�A�+ԥ���Ȑ�S! �v� 7ȋ*y3���T����O&�J���?c0��z�ÙT��d��¦L�L2��W���$H���*zh�l�'�	H漸����w��h�E��.�<겥�O����O
�(G��!��B���Q*�?y@�R�-�y��L��>����U���a8��l��6�'��	� m�$SM~:�#ɀ�i��b3c�L�:3c�ƟH�'�b�'z" �T�4Y5T"w�|QE�OZXHF�J<Dg,)�-�)+�4�XG�'<�s �D!ZGyh�� J���'.aθj�+�2dH���-L��0<1C�Uӟ\�Ik~�b^?MĔ��ЙA��x�K����0>-E|��!f�3t�<��)B�����$���l�ϊ���X�`����I��O�ʓV	���(O�So��'Wbce'L'
4�Y���kR�:�'B�S+9F�����W���*���O>U���A8,?4R@��%��A��k;?�VV�I%Ny��Ǟ/p,�1��I�!CS���cY��
d� �.m(�	35x�D�O4�}Z��� V���Ht�D·�Ѡ}��Ĳ�"O���p��	�e��/a*�*r�ɑ�h��D"�㗠<����fڣq�hP��'���1��4�Q�d9V�M2	�\<s�cL�j�~�! `-D�`z�ʕ�;$����I1'A:I�e=D�|���,m��g�:w[ˑb&D�4��L	�ƅk�Pt�jZ�w�VB�Ic�8�c�F0CD,����ObC�\��rB	�h� �	��8SZ˓�^���:��Abr�W�L��S3oU67'4C�	|��P4
Y�z�-so�'�B�9$:�[r�!�����.�!ZfC�	�&�����ү6|m&!J�AC�	�z�:����>�X�і��
3���d�u��d -K��"r��I��i�so<RT!�� e��a�F� >�,
"��6D!�$�-Oz���",YȘPF"O���2bΩF�V��5��l��Pv"O� Ňw�(�9�B���VER�"O`SV��HJ�i:�aP-�����퉸'8j�~����HT"˝9�iLC�<�W��4H:~�5�8C���S�<!`�ϱH�x	�ի"�ȡ���g�<�eA�&ː%���L? ��7�`�<c'�n�B�cU�ٌ�u��R�<	5(P�b��)�G�H�UVĉ3�̟���D"�S�O	r<`C�E�W��ЊeK�v;��p"O �ɦ��?>|@x�tj�8l:TQ�"O�-�S	.wy0�'�0���"O� 8 #��29�т%���9-½��"O�4J1`ˊ�pm� bO�;�)�O�xЍT�az12l�!���S��1ڴ�K&\=&z��E���(-�����%C�w{�$���H��]ע�	�B��?(�͚�(�2f\e`A힏�<b���n����r����ᕂ6Px�@Z1M����P�'��ܒ�L��&hP��F��LKAHm��0'��t�j'��-��9��d&��Ĕ���8�|*$��k�VX���(~�Z}�d�byB�'J�@T-�,|(��4KV`,�������[��H#	6T�0���>H��ʓt��}��?���L�$�F@ �t�r�2h�3��0�`nb��1�
3T��p1�퇉6���g͗�H�T�K!�������a�Ч\]B5r1O�d��N��i��Z�c>\u�t�kV�O��
YҨ�	�v~��3ɓ��y�E���?������D��d�!Q�H �	��_�p)1��h8D�42�J��$�����I����6ړ$r�?-6B֤���E�ԱEYP�[��]�ܚ�'"DIҟ'�����R׺���cE�f}��*��T(sn�&k�aP(��EW����Ֆ?��}2�Ԝ
�V�ᐯ^2�J�����t9��sKف:��i�jY�m>n�h̟Ri�>�
�)�M����^$�������I
r�'gў��%�$��be+`���TOK�׆�����A� hM#c���o����;�HO�)�O˓r�`��Ň8l��0 ��`ec����?9!�v���Y�N@(tP��N�R7��h��%�h��}�j����(�|yF~�ܙ ��hGE�)@��$�Y�"o��ёL�1�����^%c`5�g�����L�6���eЕb`
�z��IF�`�IQ�'W�D�!�Y�Z�V䁗k�$
71�e)D����2w8�\��%õ j�ys�&�<م�i�X��E�m��>�B��MO_ Q����C�B��č1�y�����?Y��-��ќn�R�3fL�zj,�ك ��i��E��#�*>��d�T ?ʓfj�`G�Z�<��V%�����&�s2��s&	�@.���(��da��{�e,�D^�T�	��M�՗�$���t���1ZwJшC����&�O� bR�D�O������
6�����'��4_�U�UB]�S���#��	ZF��'q֐9�'&2��>�7h��l��D���"���٦O��<IJ6�^q
��[����^��QS*,�Ӌ%�������]܂ ��l �mxd�I(K�P��υ�.�쐸����,P��e��j�q��4�R̋�8Q��2�WU�x�'0O�4��'�t7͔OyJ~jϟ� b�q햵di<�䆎�?`��p"O�D�E*!7������'+�͉2�	�ȟ�d�e�	#M���d��;S,-��i�O:ʓ&���ɘ!���b�ዃ\��;�� �H>�=x��7SiR���j	0��x��5�b�ُTi��'�"�`S��P�l�r`��>���� ��<���ƮY�hc�헟��i[m��ԠM��W��좀zbS2<t.|)b	�Oyr����?yҵi3�3�d���A˖t�@��Hɜ�V1��#6D�`���Bh�.�I#��2E�>�y�L�O�	Fz�ORW�,��L�}<�d����� �D$��gZ/)�d�0lLҟ �I۟��I�u��'��0�܉���#6�pb 9Y�L�ZШ�Dެ�[�F	tU� ��o6?��eH����(O�̋C��d:���$\
k�̉B�)�T��a2Ř2;�'h�>�C�J�=TPPu�>�DUܟ��4��@1j� P�!lTҀF���MK��N�'J���2
4�C���R�1��*�Q� �@�{Ɛ<� O�-'�BД'V6��O�˓A�4`@��?������#�!$�`98B7�ᘳ� ;�?!��ـ�?����?��ǚ<V�Z���d*�M�҇m�,��Y�LR��6vO�)�΅�Y��#>�&�{~�!��h�$1�r	�p��>u��ىօ�,���%�K=Z��%PQ��=Q]�kS�'�I�/g������HN|���۩OG��o{��h��J2ƌ�O~�$?�)§�y2C)�P�`�SyN>�Zf
����,�S�4,w�VMlZB�$�� �ۍQ�5�RM�3МT�'1��'=��'Gr�'�b�'��Ι5<Y��o�1Ӷ��"s� b�:c�d����)
0ɺ�*�C����}�Tѓ�<��K��?����,�`A��+B�\\g��Y�j)kU�ia�H܋k���eR��'����'��$
�h��d��9"�2T@��M%n���+RmhӺ�dX�����z�,)�)�?7��,!�'�y�A]�*��X�cN<:�(Q����ҥ�Iܟ����X�<�Yw��'����'fv���E�`hgD2N<�(×&_f���'mϳpf�0O�xp�۟�^wS�=�>�d�=*���H�	RV(i��s66��I����P�D�?_w�b�'d��O�͒�i�D=����&� ���L�OXY$�'�������O�%��ҟ��L�._���w�1g�<\�0�*{9 �#C!zӦ�	�.���O6D��?���ןX�D�� �H�b)<fUR,��T扥.��OP���?�'��L���O����� ȈP�&Tm}0ii`��=&"9jP�h�؀���+\�d�O�	�P h���'@r�H�P.6Y�����T/�,h���k��e�Bd�e�8�5-T����4���x�����tS�T-I��%�PcGzD��%F�L���</h6M�^}"��b7���?������А|�q!%/Ubx�JF�O��!�䞈VŚq�c��a���3��D17����'d�	؟��	�h�I�����ܟt*Fj	�|��YhCj��<�8�Zчѝ�M���?a(O���?y���?���)��lIǯ˿Tf๐��V�,�{R�i���'r�'"X������)~��*@�ȓ_Y@t�#�=r; �X޴�?���?����?Q�����O~�	�A�btb�
�74Ҷ��}�*���<1/O��x��zE:e�d�ߝ06,���h2���?y-O�ʓ"��D�C��H��J�4)��P���'��	���'��'Y{jY�!�
J�y��U�w�9����h�ǁŒ"�ؐ**�3%ՂC�	�iz��3Q�ͥ�P�C V[@B�I�uP`�4�ğ	��4��k�0:B�ɣK��eCDZ01D��P�O�-�6B�4%�
P�T�t֚��Ut�p#?!���?���?���U,%aV�^�8��M�-T%o�fm��i�R�'�r�']��'j��'�b�'Ȫ��q,�$D���Ȅ$؏5w���/u���$�O��$�Ob���O�$�O:��O*���	��G fd�g3�l|�$N���	ܟ ��ɟ����l�I����џ�����l�����@6���5���M����?1���?	��?����?q���?�M_N������4a�=[ʗ�k՛�'���'�b�'�r�'`�'�r͔�Wv���"jw�pɑ266�O�d�O>���O����O��d�O��˜m3�qآcA`>����@�$9�]l������������	ڟ��	ܟH�I4ء���2�D� ��ئ�V͡�4�?���?���?����?����?i��䵸sMQ�V��2���<f'j��R�i|��'���'E�'���'��'f�m��*0o1\�����nYj�(�b�H���O����O��$�O�$�O����O<����M	R���A�� :�\�������	ݟ\��؟��Iޟ������	Ο�)�Ă���-�W�
-HƨЯ��6��O��d�O��D�O �$�O��D�O^���uFN�2'K˾c�P�F쇝!��hox~R�'w�m�O	~Kq!�3��� -e�`MF�i.�i�y��O(�O{n7-}�=� E�;OXQK&g�(�<�K�Ϝ㟌mZ�<	-O�O�V��V�]��~B���#P>��!ǷB�V�ZD)T2�?��Y�`~(
$)�hO��y�d#�	��r��k[
n��хO�Or���I����ܘ'�� ��E@.\�� 8՜L�����Iy2�'��V6OHʓ>S���d�L�Od$PFf�y5��'�|�q �.xg��O�I�^��īo�� ��Y�Լ#s�
�fU`Q�vN�<Y+Ob�d,�g?�rg�� �*����L�lE`�А&���aڴ+�r��'E~6�.�i>Չ�#Q��X3�L�4�f����<��M��1�<� /�U~r"�Zdd���º�!'еF���RkǇh~��ҏ�Q�'Fb]�x�|�@D �@��h	.T� @�'�Ly��{���R�$2��[��㦡E�k*�j�9�
�.O���j���Iw�O�F����5%AZ郙z&��rRa�EۦL"�Oz�I�H/o޾]���S�[t0,�1��w;���C	q�!�g�1�&#C�M:� Z�c�1ODI*���`��]���΃�-�E��H���ܠx��a�O 7va����%ֹY�Tِ���!!��fP�M:&˚W��2	D�F���ۣm��yѥ%Xj�i#��^�^z�[���&xN�E �1\j���"C"B(��ԙ[���f��O����O�7MSJ ���4W��X��Ft4ݔ'�RA��' �'r�O?B�'�v��%�H胰�^����"���:�{�'��	ܟ�'�¿i����\0έ��S�5���P�����CQ�^��Z�Xibh��)1rlx�Kd�Y��U�ѥ��~�����:u4�
�bY(�$`�o��@X��vF��b�́(�a��m	1����ާ�R�S��.����	����I@�Ö4��/])���c1*
�<Y���	'���0+�7 �� q1�Ɯ@M�S,Z 5<�Q�6���C6(�;�T0�CF�.^*���`J�&R�
�3�4p�Be�Z��\���*�/����E� BM�Yez�7H1[�$DK!hѴ~9H���*Ց0�z��Æͷ��v�'�2�'i�tC�<s�P�AHt "�gD2��Ў��p�'���x��4��'��q Lv���$�M'x��	&h��|z�4�?���?!��+�'�B&�}�,R��$��m�C�,6~�>I�O��$�O�Ӣ�wb��
��2w���&c�O����O���H5R<����O`�'�?ɛ'�U�����y!`b̙TX�|*���8*1O���h2���Od���Ojl c!Hh��p��5d�O��Y	nw��$�<�	ҟ`%�8��I
R�8!�BR�|�T��� �Yyr'/̘'��'��Z����gT�b�X�y�o�.
�ȔXn��ת�q��?iO>!-O8)j�� 8���S�!���8e���G8�1O���On�D�O�FFz�S����ЪH�2\2D
Vv}|�d�O��D�O@�Ok�ic��'�L��3�N�lq�Ԣ�7>R����36#��ßH������'iFm���,�i�<O����<o|�_�-e(�$�O�O*�9�n�=�uM!-�$9���_�b�mc�L�ӟ���� ����s����<�I�d�I�?Qb��Le�Ʃ3u��u����[�I�p��,:W�[v'+�?a;un��g�}�)>�v8[s�O��A��s׼iR����	��Q�"h�Lk�oM�,d.Ғ�F 'G�V���2l&�Sܧm�t�vIH�R,B�a��f�޹��U��ɟ<�	˟��ܟ���B����D.�y���T*�m���[d*�E]�n��X�y��	�O�$YCHz��3
ވ��X��Ҧ������I�<���ڟ��I��@�	˟��@✔u&j]C��;gO4�r�h�ƟL%��[`��F�����I�|2��З~����n�	sҤ*׭�ğ\�ɏw�z}+�4�?)��?���g����<���֧fY��`�X3.�z��tMy����y"�'�b�'c��'���0WNv�3Q�V�	����4��L��A��F��M���?)���?)PR?��'��.(Sƭs��/6���4B��娝't�Iҟ��	џ���͟��Jс�M# OOt\ܪ#�Y#����,�*�?���?9��?�������O�$�;�T\���,���ӥD�m�:�)N�OB���O����Of�'U':Li�i��'(�IQ%��8d16�I�E"^��d*R�'c�'RV���I�`b�X~b�U���*K��0��HB���$�?����?���?�&%�m̛F�'h�'��$bޑf�0�Άu����O�(1qR�'�I��IA@>U�	ly�O����q
�$;��q�����Tt
����'���'��:u�`�����OH�D��^�	�O� �S��*"b�CW%�@�BЂ�)�<	���������|ɟ�`���;\�	[�*�+Q�4�X�'r@�U�p�&�$�O�����I�O~��O��sa�zxY�S@]�xa�� p��O��RT��O����<ͧ��'�?���S�)�|�y C#�������L�V�'b�'�jũ�Ot�'���'�RC
E�tiP�-�N��X�䗹��	vyr�W���4�d��O��d�7"C���$&"m:҅�;GFl���Oh�� ���	П0�I������~�I![H$
#�V- d��ʐ����<˓G���?����?���?I/��|J0ND�N0h�mW��eK�޲;�	o���4����X��2��I�<�����dc��ڊ�� ��I��q�d��c��$�<!��?Q��?���@�=�T�ib� ��o]5y~�������d��*W�'r�'��'"_�`�I�%���<--�Y2d�!>�=�%.`��U�	џ�����D�	����6���ݴ�?���&N@�	��԰}vX��Շ>���`��?Y��?,O����e��0?ICN�-��`Vk���`�ѡ�៼��ڟ���ݟ�롉ޗ�M+���?����:�.�']�Z2E��U�Yh�Z��?q����O��p5�d�D�<ͧ�� xy3�>{�P�1���D9��#��'�2�'�d8��h�����O��D���I�O�QBkIm�h�r����<���c��<��Ej���?Q*O�)>��D_��=�BR\\�{�ɏП�Q��\��M���?Q��*�'�?i���?)�@M�a�"����E�F9�h3�G��?��	�?a����4�������,jɜ��T�J0U"����H��n���p��ܟ�) ���?������Ɵ����-'k6��@��8:Tj�\ ��������I<ZHq���L��?��Iʟ�3C,٘@B(�e��v��8� �ȟ����J `�qߴ�?���?��>��S�<9��#F���%L�Qx�n)Nd�'w�Ё�O0���O��d�O��'h9�|���,G�����0��&ET,���'-�'���~�.O��Q\�8��nY�c����b��)����1O��D�OJ���O�ʧ�?"P���f��4?AJ���
]�=�D|�t�N�,�r�'��'b�'H�I������o>!�≲^���h� M/?bܥ�'��� �I:	�,���L�I��!S��MC��?�]�M��\�W��G�К����?����?q���d�O���72���}�Pu1�,,ȞQ3c/�.H�Fm��؟��I�����?W�L�*ܴ�?���?��&��0�&�Ԡg�F��u!�),l$����?�)O����6���&�4���� V�<Ha��耨��!�n�Ob���O5��ۦ����8�I�?���̟<A� ��X��4ذ�oRm�&JPoy��'�:�:��'�ɧ���?Q��2<��4�ݿ�\)��O�q2���9���� �I�?a�����Iҟ�j��=(�RWd̯@-И+W-��,'�J��������E�v>�&?����[ �x�c�%��!'Bu��4�?����?��'˫�����?���?��L���uu0�J���#n[h�����?��k��9����䧉���?Ʌ�'�H��ŭN�rӞēB�O�?)�4��M� �iSr�'O��'��'�y��߭Q�L���'���{��ӂ���B[1O4���ON���O���_��@�r�>P3ҎT�k�L�뢎�Ԧ��I�����񟰚��,��?�`/V	x�bq��t"z��C�PVP(��'��'���'-�8C�&��'p5�����A�����eDh�Y�'���' �'��	�?}��IDr2u� �$=4�i�щ��tBl��?a��?�-O�Ir��Ff�S'�����-������4F����I��%���'�n=3�{�/3~L�����S:��51e!�?9���?�+O��k'��S���$��>�����e��>�M�bd�e M%�H�'Q�i��ԟ �$%�>zD�K�6NF�1���'S�l�$��4��	�O<��py���m.D q�O��J�;1�\3�?�.O����)�����1O��^��A�lm����0%�4�l�ޟ�Iܟ�����O�\2&�Yg�H�N���8���ON����)�'�?y����Q�!V	A/r�	2�BS��'b�'UB��*�d�O���m�p����]���U͌�>И@�B�7����6c��I�P�ɇiQ<�B�-H:������q�"u�����焜��'���|"�מZ��Z��g8t<QE�ƍ&���.,�c�����X�IAyb���RZ�q��R�/�n� �,���[%�?�d�OB�D6�D�<Y׃��kU�N�0	Qw��^2@�<a���?�����O}��,̧G�>�X'�+l[.<�P�XHt��?����䓟�
K'��Y_��[��X��f`cLV"$��	���������'��U8 &���/HJyj2A�h�)��#1�l���OD�OnʓZ��9�=)be��.E�x�q�W%1-�Z����	��P�'����g�+�i�OF��A�a� �"�8m�RY9lʣt�X�OP�@Zz�Dx�O")9�lܯ���%삜p9������$�1|z�lK���'�T/�<��IH�'�*�Fo(@�d�
wiݟ �'j&�*�����"F�6�`�qԄ5X⩐���"�!{�6��O>���O~�i]�����:���>����%�����G�U�R�^�O>���w�j���}�� ��� #��`ߴ�?���?�Dd߀s�'b�'��$2d�%H��][��Ա�L�2!��O�})��$�O^�d�O.�yǈD M9� ⅮǗF�v�y��ON���"d��q%���	��T'���`��42j�#B�ȬC����a��Ry҂����'�b�'��[����?CV���Ɍ�]�N�rAæI���(�}��'�'��I%��8�$cU���̫�˰@���B�&�����I֟�'?�#���00
�'\�cv$r���n�f%r��|��'��'w�	����	4L�:�����!5��QV�4�J˓�?	��?!-O��Y�Z��d]{����|�d�r����T
x9��՟�&�<�'2<� �{ro��btĐ���W�fd�&dW��?)��?q-O QPG�_�S����S9CO�Pi`Ƅ21�4��(�4g4�%�0�'��1��ԟ��*� ��Fp����{�� q�'�I'��ߴ��)�OZ��]|y⁞*&�Y1�9O,���6��?i*O���C�)�9k�Լ�ThV,��l�pڝ!6^�����n�ΟD��˟ЗϘ't.aZ�gT�9���ZЁQu+��S�'�H*`�4�1Ov��'� v�����y;�1س!�=,�N��fwӄ�D�O0�d�Q՜�&�h��ʟ��ɐjj��#��1ϖ-x���?r�1�?�ӥ�s̓�?a��?!v�قB��]���
q��d�����?9�e��P��xB�'J��'y�I!�LY(tؖh��1���T>d��Q�'e�EÎy��'M2�'�剺u�ry�e���N\�eK�>FԺ4@@ᖥ�ē�?i�����K4�Y�%Y�*�6LBgcIQ;#��OV��O�˓[�2}y�O�����J���A���0q>�:.O.��O��O,˓v���i'�z�L�?]�>�x�U�=�:q�'���'�U��� R2��'Y�Y�X�>1f��#��v�5Q���?�J>Y*O81��D�%�|ز��ڧKa
���n]�Md��'�V�������ħ�?!�'s�^	�� 
,e��� g���Z�O>)/OtT�U�?=y���!����u��4<b����O˓0�@�i)�S��<����D�]��thW-��y����6���%sX��iAB<�SܧL����Oւx�����ajf���".zx��ߴ�?���?q�'<�O��iu�=u�d]8Re����D�O�`q1�)§�?�Ue�<T,A���+� �(�hV��'�r�'A��3��*�I��̓x��EQ�ރ\d���'�v��]�?���l̓�?����?�2N̲O|��iAN�6KnTx	ŭO=�?���t��T���$�O��O>=�R�@^��	���#M%�Zs�<ySj̓�?����?I,O� �DǕKW�0�DϨi����鈅#F�Q�>9�����P�����Aƕz��ʅ�%~\�-�d�$�O��O^���Hq��O(���u��|���:4���M>������L���8��	H����c�XtR���dz�	柀�Iڟ�'�&�I�%��ކW�.��`cI.��Qy�Ǫr�����O֒O��1�<��=y�aT9UhSb铚����Bԟ�������'6b`.P��+t���)��$)qw�נ5�~!�b�Ɠ6r �O|��~�Gx�Oe$y(�I�+�$��ː�H!X����lM�o�v�D�'9�t`�<�c�δVqx����!M�(}� �C۟H�'�Z�X���IJ�`4�a�YwID���μoJ2�R1|�7-�O4�$�O.��Vs��ҟ\���\kHB�X5B�C�=�WmΟ�bU�(�S�O���(j�l�kbѼD�&�K�_9:��6-�O@���O����W�I����I�<�
 �Go�`�9y/�0��y�u�l�<)��?���.~��;sDގKb*�BHt�Ѳ��?����v-�'f2�'��'g�]IP�غ0�����@�~�0B�[�x��"�ş|�I����'q��pd$�7� �A�e˜<9
qJ",@�DOv�D�O\�Ot�/>�)b��?�:� �@�e�Z�r�r̓�?���?�+O܅�2ʈ�?�dDN]�L���`�tE���<����?Y�����O�J���i���`I5I��
ӌ���\�<q�	��T�I���'��(ٰ�(�i�?�2@�5@mn���%d)���O�Ķ<����?��D�^��'Eԩ��M��u��H������?I����Od�e'>M�I�?�eۧ'h�@s]�1bD!G8&���gy��'���������ӧT�<�9��N#�T��Ck��Ʃ��Zy���JnX6�|z����R��c�[�HNX��@e�lyp��O����O�� �.�i>�'瞝���(r`=csg�62"���ق���iR��'�"�O�O��d�!V�6)�qA������̷x���$׸k���3�I�����)�D��c�W�ʬkࣃ;�M����?���/��L�p���O
�"��-;S�L
&베����J�@�-2�I��	۟��$�{�F�:�'�"r�b$�M�����Ƀ ~�9�}��'a�'8�2����/�2 �fdJ�J��6X���wG4������֟,�''J�0�̋0;:���%��~3�yS"M47�Ol���OL�On���O<�'K%�< �Q.��7aLp)ԨJb��<���?a���D�x�z�S�I1��:B�%�P5 V���u@���?I����?A����h��� �H�'�]�l肃� v#���*O|�$�O����<�NȃZ;�O�$8����"*���˙<L��q#�'���|2�'���R��y����(���$&�tRg
׉I�bt�p��Oj���Or˓~b����t�'���`��)ͶU(t�7�s� 7T��'~��'@����' ɧ��)���h{��	0u��e�)�?�)OR��L�ԦU�O�R�O��Y��%`�喂pu�R`N\���	,���J�d�	Y�)��.Th{d��lmh8���`����}خ�o�ǟ��Iڟ���+�ē�?)���Z�`�M�d3��G'�?11�̩�?�O>E�D�'=�)MV�z��LN�
Q !�q�F���O���ȐJ*t1&����ɟ�ΓoJ@@2/ѡ	H%�ȋ�� ��@�	&�$&?=��՟��'u�|�1Po�DY��2�j�Y����Iޟ�s�-ݐ�ē�?1����=��h� Si�A��AQ�=4��)Ot�ȵ��OPʓ�?��䧨� �\�u'���A8���*CĄpd��_�O����O<�O����O�|�vJծ3�d� �ż.u�Љ���p��<	��?����d�,X����S�"IxԫA�l�P��Ĝi����?���䓀?��������м��݋XVԄp�� V̵�,On���O�Ĳ<ii�s��O��E)��X�M],e�GO<�\��f�'�Ҕ|r�'����'_\����%kd�_ �� ���?���䛫VH��%>���?�@�#K)g���K��p��3��KP��⟀���@�?�'I���k��8��L��ùphD8�DJ�<+��I�#*̐�̫�ǆ�E�,��^�?y�����	�4�}P�ͦJ�L����\�h�T�|�'���'o�'�b�'J��q����hJ"�y(��'y�6�yӐ��Iן,�	�?9'?����q�����W1�������2`ĉ� T35W���P&����QZ�gK�24A���
 pX�b`	�I�l�BB�8�nqcpMĢKU���E�K uƾ<1��ܤ �� ����}a2Au�'��$����0:,��f�=
R ��mO#,��0���1zb(��A��D"��	.�����,��0oJ)8���9w���ri�&i����q��I����C��+R�ޅc�;�@x���7��Z�l�<[^y��n�]��:�O�~:���7��,;h ـ��N5K+ C�D��D�=[`��d�$uH�"�O���O���5K`�dY�M7tUP8`&A���0DD�V�B��Hڟ�h��T`�b>O��Ae�Ӆ˨\�a�T)L)3b_��鲬G>(��QdFD�
M�fcY��Έe:�]#�h�q�g�r�e���ǡ�j5
e�|�Lǡ�?�}&�L3w���	���`��
$�$�8D��2� �<�9+�Δ6s�4�!}�"�S��!�F��T��13�x�J�B[(\n�¯�nF����'r�'���yݡ��ß�ͧ!��uLS�L5���L\u|�x���;n�t�W�Y��xRG�� ���02ֆq̸dȠ`�+%SUтf[�6i�'hƃ&+b�2�C�-
P�����F�f��!��s�	�GN�|yǅͅT�"V�F�!���#���O��d6���'�eF	Z/#Br�)PJ��a�h���DN�3b�2���d���;.e�=�1�i:�U���e�����bӲ�z��Ϲ�v��4�͘f�i3 /����+#������ϧ.��K1L�U���B39O>6낢��Fa>h�� �g�=,O����kO5l�^Uir	O�<�d��=�~����^4=x\p��OX��1��O���>�W���b���O�m\�ݸŁ�V���=9s-@6P�d������ (z(<A�/ۀ|�z�� ���W.�Œ���� �?Y(O�ԑB�\¦���ȟL�O�-30�i*�0�t�G� �~�ە��?#FE#���O����/jt-P0�X�$*4���(���'��	��-��C0�֖�ta	�30�'D�Y���QN�P惕�Ei�L���TH vW�:3���V����SV`cFh���5����ɦ��S�'>�A���`�aJ�j��a�����T**Ta����U���b�3 �X��I�(O��Z&�O3�R��Ǝ�:�$ᩇa�.�M[��?i��2�$��"�A�?���?������ ��hǰ��ˍG��}"�����'��	�z̰٪`�Ε/�<<y�N\�3٦��>)%bAoX��x��L�B��5�F�zj�رe�	.��'m���S�g�I*{C��*ѦC*O6 �&.ܭq6�C�ɴ B1Z�ת7(d���-���*����?I`&�	�5��YPC(ȍ-���z��t�
����?���?���:���O>�Da>U� nY�;�f�ʁ&�9��-!��%�^���IZ�(\���	۰<I�%�3S�Jp"����
r�l�X�$+�2�H?8��1��7�ayR�8f�~�D �1)D��Ѽ(	)a��)�4P(�'���'��O�Py��] I�\��6`���,�ڂ"Ot�!@e&p(�Ʉ�|nf�S���A}�T� ��.�MC���M�$ʓ�� �1E(E	'��A��%N���'x�i[�'��8��P���u`4@񫙾z��y(n�����W+7f�)SyX�y�k��2.��f�_&E#���0��
	Fr���-����@B�nf`-x�L���֏/qO(�K�'*�'�D�j�O�:Ix�2���j#
���'��ܠ�&U8>���4�H	^LRU��'��Q��N"a��36�;kX�Z0����'�BI��y�����Oʧg���ߴH�nuBRFҒ*,��FT*;PN��T�'�#�5YD��#��k���C�d^	#:�}������"|XJ���� �H�YA�A��'�!˰bߚ&ke[%�F�A2x6�5RV�Cӄͧn�a�'+�@�`�OO�(b���x≞<�d�d�}�)�S�>�T����ڜH�ܜ*t�W9�C��
�t���	R�{A�l3E�C1%Ӓ��dX�'����G0��-�R��T,�
G�ߦ�������9����-�͟�	�8���Zx���+�b)��D��`��׮�JX%���?ѣ��$|�Z|�|&��[�JҼ{lQq� �8=�B��2�d����@�upcj�!� a��`��z�`���wg2����߶]����c�++���zt��I�I*)�����x
� �J��=��T����: �*�"O�d�㭎 �fъ��&m@�`�Ք>Y��i>m&�L
%a�07uH<!�A	*�J 
c�Ǥs�x)J�k���?)���?���:t���O���i>e�)}~<xq�	�\�c�#I���a�$AO�^ �iɅ�6U@\Ì��>b�ޔ(���6��0x�C��?4�C�f|�p�2J�9�Z F�!T��(I�%*�2�O�8)��R4=�E�q�P�`+��nϳ\��8�O�ܙW�R�b�'O6��؃��'}�'K�=cv�������J�6Q��ʋ{R�d��O�����Yɦ�	����7h'��PCX1u�Zy0����?��z ��?��O`,D����$D���A�o�[�0�PAK՝VMܽr�J�K�( ד!ښ#?Qh��WVn��"R�@���J����$�Σ>g,2gXK��%�$*B�6<j0�9���6,��E�	�%���4�D>쵉5�J�VC�I�1B�1b1@ǕMxx���%,��<��4�8�Z'B�c���Y����f$�A�V;p �OhY����M��ܟ�OY�,�ñiM~\0��@:�|��	\g�Ⱥ�D�O��ĕYbV��d��m��yQ����'����#>f-���U��
�i�we�'�F��FJ��%��:�ñ�21!��\��y��)�1}4|0�&"	7l�4A��Ɉ�!�pf�)�D���l�r�l�����~"`�D��d��`�c���R��X��?i	�K�`��I�@�r�B�BY�� ��I��(O�[��QPs��@��؏s�� :D;�M;��?y��'2�S 
�"�?q���?���5v��hB(H�	�Nnl�b��g}�;�y�n���<	���A*��)��$Q'0Q��ZM�o{���>^��V��c:T��p�C#^h���|C�?�}&�t"`A<%堠k�� 8h�,��'"D�D���1
�J[�L^�$*n; �-}B�&��|BJ<��[8I"}���<��Y�QOd�y��/"�r�'�B�' ����4���|j��<p�[���I�n��g�.��Y���8$����??dd����˟vf
� ��b<�DC�BP؆g#�p2�*^�4��	&�p?��iЋcT`X��I�0q��J�w�<�7�G(*.<���f�Hơ�Wܓr�֑|,�$l�6��O\6-Q�`�+J_�j�h�e��D]�	��4@WiJğ����|��Rڟ@$�� ʈ>Ѵ�* nЦ1�F�0�$,O,���$
"
G�E#�"�}�L�R�+�4>ay2E��?��>�w	��q� �;A �[.����PW�<i�GD�:/� �CF�c��y���\(<	ԭ������\<z���[��ʄrĚ��H>��'Iś�'�B\>eh �Ħ��J�[�bHp�oń��i���?��_���I�֘��Y���� F4�8T��BDw����%�DM�J�b?I8�jX;"���ȗ�D�R�� ���8� 3��)C5i��@�N�ir�iq�\$�!�91w �ɗڛ����[�7�xR� ʓ*�.	Q�*�M����J��dxb�r�^��O�����(U`�F�O����O���w�R�E��7S��q�Ё��zZ��C�X@�@����O�YBʚR�1��'�{�螀bŦ!q��ʒuبMA�,ͨw�6����O0 R��A�g�I.P�P(c�T
U�T!�e͍DL��B�i���,hn �i>���k�T,�(�L
?x���z�F�W!L��ȓW��c�-�X�zu����Y�f��OEzuӐ���>@��1/7@E�&L\�\}�U9A�R��q���n�2�'��'-B��$�I�|�4�]=��A����b�+���dP���~R�l�5�<z���S,ڽa�q�O�o<�u��K0� �pk�8�L��1,�S���	%�p?YiKu� �g,�)c}ƀ��`�<�m�gT��ěBnT���KYܓHU��|2(Fi��6m�O�7��;��4���F;V�V9���6OZLM�IןD(��Uџ@���|�w,K�26���N�6�u�Pi�+2ӄ����� >(���X�HHN[�K� �r�<���� Rh|��x$��b���!h��d;v�B����a���;�t��E�'Ƣ<�aL��'���u@ȳM?f(��Y�]�.�;ң9D����]/�t��M+.Z}�B�7���R$��@� ��ŀ	L�m� �$�x�WD�2����Ofʧf�Y��4S*�P�0,N98\ �UgY��nh0u�'� �n~E�b
���|������ �;6Ą��De�Qt�xgD���hSP�NK�O��� ���a����+fp�`�A^T�Ƀ%W���T���aش�?�����7�֙B'���-B	�ԃ��'���� &���c} =H��u����'�r�<)$e�8i/6|I�K $'izSkK,X6��O��$�O(1Q��0�H�D�O�$�O2�ح-{����,�,e����k 5��kA�V�d#vک���x"�E?8^��h��&���z��_q�8`��>Yʆ����'�T=�(�(+��R�4*Ơ�B��;N�'-Π��S�g�-}����Y�ʮ쀔c�:�B�	'l�&T(v�,y�jaK�`t��'0"=�'��IJ�X�O(rX@Ar��#��m1`��(E�n|	'�'=2�'�Bnx�y�	̟�Χ1�<�����",�X�)��H�0�dn�00X���1�ņ,\Ճ�+ߐ��ON��PNOd���se�QԩT˖�8������I"�=$cp��7���>����0�D��v����5FL��MG����'�26��I���p��z�(w�xh�H|���O�0�x|�o�<� c�%;��hÞ�`j�B��`�YJ���'�3N�lmZ��2޴�M��dR)/0�c�D�9���U�`���'?��;���'o�i��ީ�ėt0���߈��,A�m�V3�$@�>(`��2��Oh�v�
�R��[Rf�/���Hf+$&����'��
�[�^�
�?�w˟ߟ41J���ލB.�l	���i(=���7D���PGǬeq@��a���i��2��5��S��Fp|��p׉��^��-#j%�\�0fܫ�Ms���?	*��<�i��p���|��t��eT�tݖݒ�h�ȟ��IO1��I7k]6:�jYq�B	L�f4Y��l�'J01Ä%[�G��TIT!Q�a�<'��Q.N�Y��\x'�=P�*����̺;���?z��S�M���=#�ٕ�V�u�.t'�:���O�X$�b?��^0(�lP-�x!dEN�B�ɚBGȤ[�f�$%� �$MEx���Zd�'4��z���A���;g�U���x�H�������	#�h�����X�I�p����!T#ؑ~�X�`����:}��"[
q*�P�ǌ>��ls�/�.|C��|J������& �0�#J��:{�D��l0q���`�c�J*gKl=��@L�S��Z�=��HAn�+q����]r�&!k&K����q�&1�)�3��Q����TNK?�	bd��M�!���S�@q0%�H�C�\�Ŭ���;x���e�I�{��A×�L���91זx"�#'@�,u���J��?1��?1���0�D�O���s͒a�$$AsK�Yn ]�C*V�rb,xU��A#�T��M+���V�'A�|0��V�f��i���0{_2�1�DO�JdmA���.ed�n�ڦ�H��\�i)6�8p�N�7]>0	�e��3JJ�ai��^+3�j�B��A���#��7��y� � ���j���B�	x9*L(+6V�8��a�r�4�޴�?1-O�9����%����qu�ɲC�����8,�;"���?���F8������?��OT(H�����0��]k蚄`]ʸ���=,OR����D�]��D�F��bLљ ʔo�ay���?�$�>�(�"��L�r�ku'
-ή؇�/Z�!�2"�^�I1l#q�(�sR��(á�*�<Б!���;�~!����o�LH�Ÿin��'�"?f�m�<a�$D��ȝ�9� �3���L�&�C��?se��rɺ�j��S���&��5|�f�t�I�踹�	Y�!�t��V�����,y[W�F:	&����� ҥ������0<ƎJ�-Ì ���Z���5��Ef��C�S�'jB��� �+xd|X[T�\��1�ȓPcFX�n|��T뷫V/ln���	�(O�PaS���
Ͻ��$���T.�28i�4�?i���?��W�v�����?I���?���L�)3�藃{�ћ��\C8�MI��0�D��p��A�x�Y�!b��������3/�x��m�2����P�8��8`��0�3�$�}
��!bR�R�v�ZW��3~�¹�O>a����>O���p��U*���J1B
�$�"ON����b�ͨ�`�k�R��&�>a��i>�$��B1G�-%���C6�S�Uj# �(D��b�����?���?��(��N�O~�Dn>��p$�t]s��[�7a��d���+J �CE\,7�T�ƹx�ErDâ��4凈T�+I$N5���ʹMlR  Qb��I��q)�'y?���C�9P�$*�{������ĉq�F톑�W˘(o�~�)��%�~�	�Q��SE�L;Sؔ�&�yR��HBu�FK�Q���*����'��6�!�d$(�vm���n��P�c��o<���� ��*m��`��?Qχ��?����o�#��x؀&
;X1����c���5l0 "����Pi��(�	!F\ ��!Z'3��0� �\u�Џ�ygB��֡P�"��0������2�B5&�@�G!�O^�O�\ ��Xik�kЕX��x�"O�D�q&��~�*�دVvpP�&
O�,;� Y9V�̆�^5����
Z*��%I�U�	3,�~��%ٟ��|��F��M��e�XY��C�0�dԛ%�W�iL�'.����K�I̴�D�ڏQ�lX��d�~��t�aSa��:nB�s���B�l|zr�x�E��>��Y���:̈�%�M5Db��=HEֹ(��O�Z���lH H��Bs��[J1�K<��@ٟ��Iy�O8���7��̢���,l�b!Q�:MJB�ɧ\���0��L�8A`!l�K����o�'��]��̍=5=@���%{=�M����������	�Q8�Yٟ(�I��(�	:g6D(��K
���r�B��RYP]�F �}�(�{��7@�i�d��,aD,�|O���6 ����y�C�;�ļr���Ye@qP�k����P�s��0\"�A%F^J��pӔEY�w�z�b_2�a��Z�
N�3fǊ9y�B�O@�3&����ē
��MR��8QPt�6˔�n�v��s�2�y�C���X��gϮw���O�LEz�O{�'L�-�D9H�ꆅ�M��Qx�dJ(k�hS�#�O����O��$[º+���?��O�j]b�o��i��=��(�5,W�eaf�A�1�����-��<��r��Qxџ� �MD�,�C��4fS mz �ʬ	R�X wD
�^���%Ü<>�vto�2�h�h��%s��02Ҏ��#%Hʫ4W�ݐu��O�9o��Mۊ"�8�)#uD����!F�8qkE�q~�B�ɤ3�6y���H���'��  ���ش�?�)O"��æ-��ߦ��(`��˲��@́ҵ�ğ�?��Rb�|Y��?I�O'
A
&�ßrg������cVxD�҄��H�\�%��g�R���<)?џ��Κ�Q?B�K0B$�x`!��=F(��6·�[k0ը0�Y`�n��E� )9V#�	�l���D$�䁍kw(��ME4�U�VI
�!�d��< ��
UЌ��!��3Q���״ݸi���Mw��9f�@�	�D`Э;�D%�@l�����Ia�t�<l֛v�˖u�DA;f�W]B��x���O���D�OXi��"�O�c��gy�׳X�Ұ�0]:QY�� c ����W�j�Fx������ɨ�珚B�Jx�"�_��ē6�2�����S�'�t|! �	E���0ŭ�9}��0��W-����.)��a�f�g�
i���9�(O ���:��920X�o��-s���9�M���?����A
�`X-�?!���?q��ߥx6e�n+TհEh�h�Jw�X
�'/*0k˓i�tUif�Ŧ�f<c�#��C)�	�>�V`]SX�\���ʤ!���8D�=4�<���.�p�'�4���S�g�=Juαkƅز9�`*�V�/e�B�ɽB�"L�!	I�p�����H�vҠ�'�"=�r����@��5�J#�,��U��+G�T���_b��'�2�'�B�]ڟ@���|j�&��ZԦ������&݂5a�:���EoS%~6���I_���<��i�"�P��#� l��4y#o��!A���1OD.����hB��,(�Q�"��qg2�ɐ{�u³�I���&�yUΐ;�`�O~��	�#�>x�Ň�PQ[�e��%��B�5@�v$X���K���)�oڝxq���!�4��&D�!S�i��iZLIf��|8�)q�	6hㄅ���On�L(m����O���Kp��(�\�s|�EXA���^M����I�ay��1��'���1��( T��h���s9p�	˓S����$��U��C�T"�Q)�ېb�ZC��7}�Tن��^G���f	�a9�C��8Aa��3AȮ&|��j5�2�D[��$}�)lZ����I{��Ba䛆��qD���* h��q0gK�L�n�D�O"��B��=s~���I�GaXe��|Ҫ��maG�0M� ��i.	;B�x2�W6`���j�B�ɠ(0�R5�����l�0b�O�&�J��%+�h�熉z��I!L<�R�̟T�<�~b�C\�,�T��g�	0H��3�n
S�<����dm�-���-Av2b�mOP8�H��������4K��XS�[F�VQ�ٴ�?i���?��I�y��$����?���?�ݗk�^a#�ֽ`5���(�L|��y��3��<�J�n��Iѹw�D�B"�CD�2�H؇剎�$DIRO�`�v�����#sK蘑�|�&�#�?�}&��I�����xC� �)R|�h�,>D��0�ջ~�Х��u ����:}"�4�S�'n�I!4�ƺ
њ�:��~��v��?W�Q���'�r�'���f�M����\ͧd�`@P&M�^M⨪QI�c�;g��u�v ���C�y��0��ݸD����RG֋�����Ŵ�a)ϟ�d=` ̆	K�V�R�g���M�`EӵdJY�"�T���e(�'L`r���B�-?���ƄRܟ�;޴z��F�'2��$�>yc"N,K�|x�ҮQ�q����R��F�<�U(յSQ�P�BA15�#Ao}ܓ1(�����ҁX/����?q�t�? %1���6����D�q����Qٟ,���o������̧<�hh����B<&\k��њ0�\�P��B �A3��6k8P#2�'Þ�e���[�|D��BV�;eZ��\�2 �ce�- a*D��)��� Q�� \0"�=1BhK����F7C��a!�Q&"��*,D�|�ŨP??t���fǊ!8�칻G*,� �SH�u��r��E9[���o�2-Kt�$�܈�.��M{��?i-�nL���e��P��bU�Lx4�
Ƽ��`K�,�ן��I�(θ\*�+��G�b��D��t�cܟ��x���b��P�2�H����0�#��=r�6�:f�R�\�r1+�Oz�CDo�,A9 ���n(?�B�*eFU�-(Ҵ�ݱJ��&�q���O2b�b?���əJ��i	��8R����d�6D�̈q�R ��I�.��+���(�c"O�iDy��*y�`�h�4��L�v	�~�b�n�����ܟ�	�/�41,��������ٟ�N�..�s_�aH�9C�I6b�T��Qc���ua�C֫a���"�O�U̧��ɠNQRiQ&B.��z��ұB�֍҂B����D5gA�)���� /����Z�[n�Ἃ��..�@U�/Ȁ����([��OƐ��������q��u4ȣ��4�t ��k���2�C�/dM��+}��x�O6�Ez�O��'���p2���`Z�m�Pt�0��̒7H�"<k��OT�D�O��Ay�t�'*�S<'���kаdA���D��|��щ��3���25� h#��3
�d�'��u�G!�#.$���ծY&��@ӕ��zX�s�JP��3r���2���:C��#ɳ��:B��1U�@&W�ZQj�%1D�9��ן�i�4>.�&�'{�	؟ �>y� �J���X�j�Pd@F��]8�x$�8� *�0#�%�'ME*?�jT��n+�ɬ�M����D
�8�4ymZ��`m�rhs����eB{�O�R��1��?�!/ı�?y��?y�f��-���3�ۗ-:xT02�X�B���xbb�\�h]���&b���P��əx�������~�l��aeR�G�<9�CB@�f	V�Z1T��x "**K�Q�w.�	R7Zc�\�wN�O"oڈ�~B�Ú�����
4�Nh�#��&�~��'���4�lO^P���!uo�p(*/W�Ԉf�IO�����P�yN6]ʶnnCfe���A&1t�נrӢ�9Z��h�i��'��:c��lڑ�<��䢌;���R�j\d�����?��+�7'��1%��(��r䂦=��Sr���̞[�@�-��#�|�,E �ē,(Di9��s��,`��Z�?�H��s�tSx�r��n%�A<9L�q��cE�;DPЏ)�ǋ2��	۵:��L�Ê
�8q��P����V2!򄀷
������c0�a��[)X�XG{�OE��<g
��d��4c�e?4E0�m l��6�O|���Oxl+6N��̼�$�O����O��9|Q���㇡ h����.J��â< BK�5O��K~&����YM��[��!lL$���R��Fɘ�Ā�u^�Q$��+�c?��O���ae��Q R�{R�ˬ>4��
V�>�M�G�i���Ou������<!�43B�g`�� ��!K.�>3�O�}@��Q�,9���	�t�)C�]Fy�jӨ�l�ߟ�Q~~�{}rȽb�w�Ш3���"E"�	Qw"���cMR�$�O��$�O.���?Y����4��,hV�x��,Sf4�NQY�A�f�E���f��~��y�\�("֤yW�.L����*A�s:���]L�����O�°:��O�"@x�uܓ\�r�%DW��9��c�A^hd�Ǖ��z�$�*p�)?8*�X�*�t=�ȓ 8ub/A�6��bEM�G�F��=IU�i��'6h��2�rӘ�n� ��P��s�k
ժA@ƞ@���'��`���'l�;�T���
�/��qIa��zɛFB�^� �񡁘pX��ԥ��<)f�1�x3q�Y7{��o�fO~��q�ߕ`J�k�G�7�����J�+�R�'�¼i}����.R�Kƪ0�S�v��cЇ�<	�����OM,Yy&HPt0J��Ϙ`�4�ē4���;D�A#dw�lj�%V	}!8���ở,�'D|�iĩc��D�O0ʧ1�@�Sܴ2��I��7t܂]
�JV�nud�)3�'��L�?یuST��RIR&�aӘ�'��iQ3�j𙃡#J`X�$R�Of�'c�D���D���kFF��p���e5���K��?����мy����� wQb0c�)+�dU6K�s�,�o�����~bEL�#�W�Q�T�F��s�[?�(O���<���J��6h��3¡O#]�� Sm>,O.7̀¦]$�0`�I�zI�mʡ(�����
j�X@���?a��#��1�!eZ5�?����?���g�X�*4���!��1�Jz���bM�ue��1�">|̡4%ڴs/
�"����6?�T�!)�<�ĉ�J����J�%x����� }��Dm��w|RɃ4��3x3�4�O+3y��.�8��`��d� '#���Ɣ�d��D�<فƔ���>O8L+���~��I0��5)g ��"Ot��S0r@`�c�3P	c��>�0�i>%�$3�ϘR��Q� M�Ar4�(R�K2����"@A�?1��?���_���O���b>�� d��ĒO�e�#-��B`!vd��Y@��@�!"쀧�A����r4��'X�
cj�J���2
�K���e*�H�� cK[7u	X��������4tf���'���ݟ �>��kI�@����2��2K�.�,�u�<��I��6���G2b��(�r�Loܓ;���xy�+�[rf7��O�7M��A�2��xR\� EL�<5�4P��ԟ���j�ϟ��	�|"�
����$�`J��E�t��2!ӡ4�8�)R6,OUC ��I\�i��@
uުM �S�ay����?�"�>����e�V�����7�,��[C�<Id�Q�-����,Z���2��v(<��e�#9�	IP,�VOtIQ�)нx��3p`���Mc��?�/�[P�i��@� ���i��I9���N�ß�����, 1nX�M�ԭIq&��?�O����B�I��
��p+
M��&�4�hOب�E�M�H�E�BG*:9�a�K<Y�>+�A�����L� �:ș����$�aXQN�b�"GI(�d+�)��9;Taq�$)�0��5��B�I���YH�ϕ�[)�؂#��(e ����A�'}���G�|�� co�>��2g Ϧ��	ğ��	2;��W��̟X����`���9+ੑ�r�H�D�.	j5ے���4��#��isR� �T[�0z��L<�	ӎW�4�zcTg�[��0��I	�K���Y�C>#8ڹz�._��SF'�xr�wN�K%8yr\8a$�mʆ=Z��<�ɷoʎ���x"� 5��A��&E aZEbv�,�y��ؤ�:U��P��0)���ξ���HO�)3�ˇ)px�Z��
�ye���ÉǌɸlRFے1ի�'���'�rKu��I���ͧL���)�/gf�c �q��mi�LI�I��A�t��J@���ЖA���P�t�(3Z�@c�*�e�w,��$�܀
3�U02١(��Mc�b�P	�4r�'ʺ��Sx!j#�>��DŎ�]�<H�v��\��I�e��q�JӖ���H�f�"�VC�i��d�/F�@�O�g��S��4�I��M[H>���j��'g�F��Y�"�[J@�&*Ehd
 �?t��$�O�A����O��p>�"�Lc��g�M�	���	�s��YvkO	�h�z��Ձ�<�AjۇHm��&�11��U���ݛW��C�ȉ�PC��c�$�7Z�޴J���,Fh�^�z��Ƀ��I9��H�m�&YE��rFF�4��B� 9�Zd2&M�}
&�S"��#�C�I#2-<9�PH�S���9�/U,�h�Q��s�	��ٴ�?q�����\>]��7-޿�1��ɷK����{���	��<����{ �t�&�7�b��ǅ��|��)�~���À.hQ[��8	��	�B*�B�<F~޽k��<:��!C��Z�6�"$��;7����ɛ��[���`oL1ۆ��q��O<Y�U� �O>�~j'Ħ3���J)~)#�E�v�<���V� N�96�8�� �K�4�ў�9�(O�A� :v�4�ZT��kU�噰.U��M���?���}q<؛"\��?���?Y����p�#E$g��� Ó�`aZ\��!_�DR���?W<�A���.]pL�x��dB(?���[�%eR�8d�"b�8!�!T��S����zf���E��L	�QȀ�U>
�ʧ--��	�7�|5�$a��A���bs�ѻx�Y��̗��{�I�)�3�d���@;����&�� @B,e!��&�Sb��0	��\��U9M����Ox�Gz�OV�'0 ���H�V��d��bB� ���C��-�4L�OL�D�O��$\Ӻs���?��h��=Q��Ņ|z���D�ܼ{���	��_Uv����)i�ԍ[ t0#?١"T1��$Q��`up1�j�\J� 3쌚9�(���5��V����ШO����}���*rT�;6 G�|<QqG����ڴ���'F�⟼�'�ɷG{(��LT9>���0b����$6��#br�DXa��/@�0T�X��Ct�`�I��M�q�i
�ɰ\c�,Q�4�?�޴n0�{�*�n;Z�Y��ի �]�&�'�r�� W���'��ϮX��xb��;u���aK"H��
�ð<�@�}�Vє�Pu�1-G�{g�SkH���	2aZ����g���e p�g!]�6�h����`_!�Jq�`��&h�D�j�۲�``W
O�u(B*m��|b����'�]Pꈺ�'�, udu>e���/vذ�rH�"C��qx�B����'�ɧ��OR��Pm��sSD�5��H��垼Q���t����D~
�3$^%-���'�;��0(�l����7DU���(��%�!�>B_��B�܅z�����d]��'��z�a� :�LAw
�H9�'� �Z�
�uz�)K��]�b}����'��|IWo�3��A�IYR��`���� �xC%D�t�������mK�"O4y;0�J�D&��@�� I����"O��h�%�?E�5K`����"OD�R4���VF��t�!QB�i"O!�QbU�o:pq�K�V�A"O���b� � �\\���f��=r�"O�j"�ϔ
��E$L�����"O��!��.��cº��{�"O�`�� �P�-`u�XwA����"O`�Qv[��ԅH f՝&8���"O4��@�??�ٗ��)}-�H�"Ou�#��S�8��J�s<%Hp"O�L��J;f1����	�&�h@"O��!� �b���~���3"O*�q��8D�If/̼r�"�#"O�q	��'	�౳��"���)�"O�C�c��tdH�*�E�$�0|1�"Or1�'�E5"x��b �3J�<iB4"Ot}jp��0<@CgNĴx�Q�%"O>��򨑭7RD��͙�Dx1R"Ox�a:U�~���*ؗ��(Z�"O �S��H����	�s�!6"O���`�?7B<H��IQ`VM�E"O`���@�%[�a[ ��ؘA�"O��.%Z�l�Q�
����u�"O0�[R�Лv����*I ��M	"O~��1��'�48����_�4a�5"O�D��͏*�8��� �%x��%"OV=��l��HЩ����q4��0"O��PV��fL�`���=h���"O�X�@cӿF'�|��f��
�ڕٓ"O:�T'��x�ͳ�C��𩑳"O���ͥ�ة@�#'v���`�"Or��1��mn�!����:p��!�"O@Pك%�H�6R�
�� ��DZ�"O�q�&M����)���}H@�'��	{��� 2꟣u�j C�9"^C�ɟ))���G@��d��t
��*Q,#>����D�$��e�(��m鴀�1#!��	j�n�;$��`��y�CA��#&��&�S�O� A	1�Mx��f�1�$0Q	�'�d�C�Gc��1��PϦ	B�O���D^#$��Y�h?-�\E8퓻�a~�Y��3��G3�$�KP�]Ԍ�@�3D���aʢ}
H��u��v����qH0����D#�*�t�`�%���!�"OP@A%�/�$�ځ�~#�	��7O��=E��g[ ծl����v���u ��y���&�@�J��N�i7��H�Oۆ�y®c(�A�V'Ull�{`�0�ybV�nb��r� �3m��;�%��yB�)q�"`��LֹN�2�1���y�Q�s#^T"�##I:�`
1�y�,5)�ʩ�PʔI�*!�tN�yB�A�WCj�[q���q�}	�5�y2�@���	c��mk��y�Ÿ�y��٨ R2]*4GP�^أQ	�	�y�LH#T���a��_��%ZP&1�yҊ^(U�ݡf��Z\�W^�y2�"����y�Ft#!�)q��B�;u��x�Aņ�5鐍8����B�	9T�\б&g�?Z8l����nk�B䉭m%8���'��f���E�,{ZB�$(��Q%!6æA�2D�tEB�)� |����Jt�PB�5~J�E3"OD8` �^-k���j2
N"4��c�"O<=��BW,d F,H���4dxa"OXY�ч��Y+�1ഇ�4y, �u"O��c��[?!�@�*3�^�R\��"OലR�9�R�fF��/�6��"O�L!���)H�b�gEΓ/��bU"O�e�T�$�2�z�eC�v��h�"O.�i�"^��H��@�%�"Oz��P�]D�>a��M��K)�8��"O
ER!�M�g�2����M�M-URR"O^(��4O��`)P��:PHC�"O*�p�	�9v��������c"O�ˢ�X�x��tjD$����"O��P�k��V��C�K�t�X�"OB���I.d���5��.��͒�"O�Y�G�q��}YOA�T�F��A"O���BcE���Hg�|�r�)f"Ov,b�.��Q-l�x�����F�8$"Ov���OA�z���ȓ�V��$0a"O�x����h����ї����"O�!#��,N���#�K�e�l�"OND�%�<.������z�9!"O��⧝�He�Pv�΅b��
�"Ox N7(�`Ր2fC�
�N�9P"O�st�ͬ6S:����;��I[A"OJ�KU`�.���&Q^�z}A"O�Cg�۪a?��U�3	�f;!"O� ;��G�0�����"�<id"O�3WH[�\]���F�+oW��p"O�=Jp��97�%J�f%w4���g"O�(�Lե]�9��&�1CX�hSP"O��ԫI8K"ma��9qEB�"O \qw���1;����Pf��7"O�ŢC'��h�v b3�Z8'��X�!"O�X(C��b\�B&ŭ�k�"ODx�#
2�`�2�<_~����"Op�W�
R���j��ZV��"ONh����F��m����	!0���"O��[���>i����H!b;�ܙ�I�)��%�w(_�O{���PK�3�`�c�	�l��'�(�bD�7��)�æɜ~"t���'ex8��FE���Qt���p��S�'����rlB�)4�1S4�>�����'hI�a��XBB�d�'�-�F�D�H��ӳ�D%6T�ߓ=�L\rs ��~�!�6Θ1\@�����0�<yJb�3i���':,�3rɛ�7P�l"����r�}R���(�����N�$mf�L�M�T�S	b��lH��I�?y:��	\85�LC�I�#
*�1��Q2'�X��!�VWd�"� R�1h1[r�=��XU���>��t�}��(�*4�Dm���ΓN�*=d#�s�P�Id�0�4�#B2�YHQ�@8#�5���#N�.�>�rL
$�*�p4I�90#d�����c�'b�Q�(�Ș�AZ�8���"�����(�%b����/gG`\� *�s\�	��~1��p�����0���)�b��ga��(כ�Ș-��Iv�I�w���bEZ3���1�"��?�iPgX���Q�&�/Z�H��N&��÷�;�0i��I�f�,k��#8{�ȊvH��Ζ�*�̃�r��%��GO�h��5�;'�����\��u��O�j���v�x���j��٪@��n�f���_,;�Pt�~:�� �IP�TF�9��a.F"���#Y� M{E���J4A}=��hi6PO��'���ͦE��֩��#��%k����,,l2!2gl5M]\8��n�l�X�:��޿@(�
�nS�!�F�Pӆ��'`���Q�1�6%/C,n�9��$O>�0���%�:���s3^ur�_�$a� V1^�ր���ґxX4�e&L�råo�8�89���E3]3r]� k�;!XD��ɓ�"�L��G×4�xb�F�F�)��C3��<��䌰j.�81��d3"�y3�L� �V�D�P�qF�޺k� �1Ĥ�]B�t�
i�bԌ�
O�R����\����� L�0��: |��zF3L�D�+į��	 
�SB�ˮ4g&(�4��F�F�@8%w��ÆC0J��	=K�ԹŻ	Fr�W1\΢#?�N�A,�mp@bQ�>����m&V9c�� -&���Cw?�X�-�12�n�"�B�*�:XIW��;�ax��ݟI/ԁb���2�6�.��8�'w��!̷N�(�P��X	qq8�x�gZ�t�D��u���J� ��"��@t^�1�N�(����肽�x&X�MfhU\��bC�4P�as��7Hjrmb� Ϭ-<�`�&b��ӥ@��b
4R�}K�w��u)�,<<���� �Ϣ�Q
��2H"����5Iبu:�A�_(��eP�'�Y��훥F�l�U�+V=�� "4J߸QFz2j�rBt\�A���4ԩ0hP���O����B0Ä��4��D�ʕxu��;4
���������z�ϴ ��3 ؞�HH@�'0�-���8w܉TȐ�Ft�ѨO�㠎�@�h�"���yBC�?�X.e6x٭��I�		��l#�΍j~3�"O������H6=��Nβdl����@�#��&��T2�G�4T�(y��,��N��eo�@q�0�XLb�F����ЦȖ;��y��'�XHr�FZ�v\d��&�
6b �a���Y��V�5b��(�&
&�!*ZtZh�Dz�؜r��јT��&�(Izţ��հ<���|HBI���F%�R<�#nV2t��(x�)�N��r���>weh=sg�V�P��E?�U;�`�U�`�A�m�'� ��ȂG1Լ��g!i �Q��� �<�O�b���$��a��aśnW&I��'Lx��@C\v�����6؛RI.Pdp��cK<�<Q�VK�=)P�be�%j��{�oϾ`��B�Ÿ2j�d�B�(D��2)�0R�0i墀�%1���F(3�t%��7S(�kB���l�"#�I�$k
�k��Te�-��Y4;��$ՙzH*�cV-�B��	�UW�p`��	-w��xW-V�E�Z9a/'�Oh:R
[mN���L�C�Pm����P5U�hta�iH(nM�5a�㏰��Th��JSkG,i��٢gLڬ$Vj��ȓ\�x��g�p�:�]K�\��u�G|ڌGa��R�����]��~�
׬���ۅ(�X���!;yC���i+��Y�bl��pFV�'���	E�, C�Մ2�`9��ɗV���! cH��I��׀%�C��#
zuЖ&ڙ���*AfP�u��C�I4M�D��b�� ��('�C��C�I�Uu�%`D&M�F���c���"OҤ��@J�m��HbUE�-jS����"O�:���4 ly���*e���"O̰A���%S�|���)�4Q��� "OtZtC�k;�K�(BbR^V"O�yc���t:����'NX_Y "OZ��5m����)�gPt�f��7"OȱI2F֭N�J+�@�g+l��c"O-�!V�(4*���_!CΨ�Q@"O<`У�:O�{FA���jP�g"O.X���Ԋ��PI�QP����W"O$s�
E��͉�B�;�Fa"O���b@�/Y��AJ�L�	�P�XQ"O�q(�H�h\�œE��aISC0�y��я0$�] ♧V�L)�B���y2,��(hf���Rhj�,]*�y"d�Q��m�2@Ug��r�@А�y�J��-����AM�"v��Ѐ��y��#T����4*_Ĺ 錫�y�(ȭ2U̽����9�WO[��yb,��k�69#`D��z�&��7�ٶ�yr�ϐb^���*Яu��P�i۔�y��S>c�;q��T�ʸC��y���I���=:`(��E�y�.&��	���61X��ݹ�y��{����%��2;Q�X	�$P�y���!D��� �l�(���j'���y�*�"���1q,%$�4xWnP��y�,�)�B���;aHfl(�y��YZ� hfV�Z��$R!��y�Z4@�j`#fZ�C��u:&Z��'�$!y��O�r߼=���6�� �L>����|�^�7��*r��hpe]�<� p� gj�!�z���l,4<��"O��C� Dy��D���R�U%��"O>I3�^)pIؘ����	'Bɡ"O�i*�ʉ��H��&B��#W"O|GF�r���A�5@%~��"Or������0e-+�0F"O�8�7A��)�(à;�l#R"O:�[v�)sZԸ���Ԃ+�l
�"O�U{p��n�.(��Мg|�z%"OrL��I1�b)��!_�u�)8'"OVa�S+�%c<�d�go�4X<�%"O�غ�g��99�-�QnP*&}��t"Ojy �ԥ+��z#K�exȬx"O	���`ͮiR���e�L)2a"O
8Y��K�-x�ð���,u��w"O���E�Ň� ���شU��`"O�0���W�~���B�*����"O�������g����m͓v��ڶ"O
�!v�א>{&��-�3p��1�e"O�|�� 8Cن�����5��,�e"O�i�@kE'T�����˫l�~�˕"O��C�F�	�do�$��� A"O2tf������-V.����"Ox����;|W�eQ��^&N�b�2�"O�TH��N�Dd<���fvq8x�C"O ���b���������_��|"�"O��$l�Z?(,Avo��\���"OB�*���%:H�x��ך���"O���E۶���I&ߌ+�I
5"O�$�RO�8hT�A�:* <\!�"O�$�,ؒ�.��f��4x��� LoI�,��㒿.��1J��{�"~���l������4�ؓTB�9?��ʒgJ	o����	������*�3�I�n^(b I���X�S%G��&�6���FT�)��E��ha�?c���%�diH�#�%9�N	[%�Α@"`�c�G���bY��ℐ���ݽcD���w�FM��Ù&h�)��h�0�j�l�[���<����'��.E�C�^�*cD�v~*�7�f%���ĤT�V@��QΘ*rm�U:Do(?�cf��H@D "�߄�X@t*	jy�$�O�i� ,
!8�=s3\�9"M����Y�Ъk�F͑sEC�s�҅��Bߺ; ���a�<y�4c�����
�@�*���F�H�D�0�X!kx$����ɠ�
B%b�O
��2��n�   x%q{�Dߢ1��>ѳ��������F�i4O�'G���Q�K v�L��g��sԜsv�~�'��}�&n�u��O�!1ƽ�� �T��%��Bl���r%,6��~:g�@���nݹۦgŚ�JFmW�"���֨9��U�b�)q(���M���J�&n��[E�6Z�����P&���A�Iۉ���տ?21UL�K�N5��;m{���&��}ЪOJD
��6A�@�k/1rT�ףT�`�>mA�!T<v�'O�0��O��OIq�cJ�F0R��Gl�3F��| �J1?���Ƞ'����j� i�pM+� Vj�a�8L�r_mm<��b��4`ژҀ3�I;�0|
&B��W����$�$k�2�aǭ�$�T:!��RI����2�cå
�d*TX)�5(HYӣ�h9��K�d�Ǧ�'�e�S�4�F�;��O>���+��(ĪdjJ�G9D���� �wr$}#IG�K��P�Q��t�84/�p�I�i���̝{FM�<�Q/G���4K�/f�<��M$A�ʼ��C*�Z!��cR
���c���;�������&���c�X���'j�@��7* =_�0��/�L.�e&�0��'���d�r�9?#����d��U�T�+�웠13��y3^!L�viDx��!�'�ZMZ-�5��<(�Lj�(ޱ �����K�=P@ˇ
�D��j� ΑU����)EB�|�щڡ)Ɛ#F^b}��@Xv�'Y��Fy�JV^�x�#��@*���5�]��':����L��\<���C&d��.���&�gI��k�k�,�p��	�&:F�ʆ�7K#.����UKu���в%���bp��h� [�,@�/�,Yf�'9 ���p���%�:9�I\25pD,_Ba��>�d�D+fx�(Q�B�hx��Lҟ�D{�����pD W.��n"�!�3Kdt@ktW$2e�b)��HO�N#&��λ�t���
H���v���h���� �'�qO�o�~Rli1p!D�	�|8:W+��(O0:�g �>�lh3,O�Ԕ�� xH5+|��*��;Q�	��|�"1��ey��^49BB�C�)Ű�I�� �~����R�Ƕ'��(�Ɍ$n_
��cB\n�xmy����Ѹ���'��r��8C�n���	�� 
d{�O��8#�2M�������cቧL�Z�K�@'� P�E�z��y(�,AN�#g����]8���8��e��c�h�b!E��S�,���N��Q����#P��NI)\��\�5�Xy��,ps�,\���ŷ+9�O�>)+Yw��t9���2C^pp%
[�袉�D�ZQ�u;���r�^qr!K2^�剗��!���O\0����=�n�\�ny��{���?aJ��#:�&��JƜ��P�J�l��؉�	�}d�y�'�*U(1�ₚ���!��O�Ǹ���'FX@�G����� O\�.�d1��OHUI��D���`���(K���js�	����9Bʅ3U� �	��<�Q���x�KP����,0� �>'���`#����R!� �q�	��Q�0��ݑ��Р��A��t�"�� -ء����� ��O�>XwH�E���اlX��p���p������D���ȇ,���r���_��		t<:��M*9�nt 3��: �f�w)�a�=	�ןnu"7��`Sf�Bë,��H=���V%�ֺ"��X��>z)��Z2�uEl,0џpJ��^�-��I�"�V�j�8�A�*?�@M��dU>p��5)v�ɶ��X�'>
U��g�][h�؇��Q6rt�@%[��Bn�#X8#ѧT�h2��`��>Kd��4��R�Jd����G$3��X̻�(� #�5�Z�4 ������	�AH(��"	�P��%�쀡 ��֍ U�'ԦI 5z	�-9d`�%@d�t!�'���`��Q��i�D�X�'"ʩЌ}[���h��=�h�@�H�g�ʨ�`Ij��Kj��t���`p�@�3�Ȭ8�' Js.�
�:��ܪS1�I)O㞀�c�Q�[�)ppL�g�ȣ@`�>ٶD��#�=q�L%���3��[n�'u�	hr��<��s�&�6f;mQQ/��fg(ɕ'Z�z�GF�uBTt�%:[�����B�P�d�;U/T� �L��W7K�B���![b�鑳p��{��7h!,���|y���b-
��P�gMǳk>� *0� ��=Q� ��G]�"}��k�N���Dٿ< �P���_�_*~1�W�'�l̆�JB��<���A�2��]�ɍd�J�����-ib��zҍ��v��o[�(񦙓"�܍g]qO̢}�
k�=jd��6T��0Шn_�t�'��QK��PC؞d�A��4�詨EI�%B���F��O��C�����p<�Vgk�l7��F�v�R�H)N� A ���	vQ�{2$b:^��'2b ��g�&f�}A.VfT���ċ�X@�雏�	<
,�!BD�H�t��)��G5�O<�p�<�ȟ�=8�K	��X#�"������'9��D�ѦQB �34���yt\�q�y2�1_:�X�NV0��X��������242���΂%�M{2��:#=�g�;�:�9���b�>Uh�����W��<�ד�$�K�"ηjxjs*��Y:�p[$ER���}���'f�"�5�b�#��$��Tq�C� 	�T�[��'���2^����M�"f��s�&N��+�E��hOtт�����݀���4D�Ep��O��2��
@&`�V�R�Z�.�Cc���<1��* �a�R�B�7.�Ag��Ȧ��a�ƅNm2z��\J�Piՠn�lպԡ]&���G��b-գ���*,�>X4C1Dt���Щ1��D\�EOC'�e:�ۉO��Fy�kO(�@�#�Eƞh� �4g9����'�����3I�89GΎ0d�r���M0�0=��)����O�	A�&W��y'៑Ro��&gT� lL�q�EG��x"鏱��\���͙=t+��PY�:��$��3,�]���ݹ}�t)������r۔͑e�F���e�3-��tǖ��=!�џF��m�mo���!G���I�3�����/�~~ujd�{Z|beG�>9}"���GG�S��~�A�J
��&H .N�	�'Y�7D�> ܜy©�^U4� ���bL<҃k˳xp�R��D��xr%���6<�-O���O�>��G�ע3���8���<���Qc �:;tx,8�BY�X�>�c�9u���]3x�����E_�j}��f��-�6�ľ4r�h�_��^����	ܺs����I<i��iȂd���I���y�'��qă��	�<h��aآ$?��J���	g|�ᕮN�V����"������~�j�� ���➴��O�
�(�fH�J����iY�L �¶%�<H���W�r���3��$B!(mY�Ɠ4lxd+Ca.c�M#�چ�?�'
s���B�?C�!$$��r��7�����DX�C�0�0�gR;%�<]��oز`��j��)���	C.٦T=���kōv����pO���mKׇ �X<V��N�O,>��K�93�X�f�Kbr�RV��A:D�7+��+FQ�4�%.%��*_��ZՆ}c����I�;� ��Q��ep�m�5V,�D ��X>�@SYw�h��%�_�M:LRDK>:q�8���A�C h��!�O���V,'���cϮytd�H�!��4"�CW8j�T��7�f�l�I��z6�	/a��Q�n�Z�� �S#GD�?�f,� ���2���cFk�u�D���a�Jp
�#��%��/.�P�Q̾>ͧ<U���eoW�\rZ��HA�$� ��O��d2 ��W��?vv�ˉҏ	}y��s ʫ`RZ8�*��?ѓÃ�G"�$��39�R�)�'}��xF�G0�\ɵ�]2L8��"	��'�|Q�۵ޢ<�S����w@�cs8fP��B�K�	#�hd�4��0�`�(y��8��'�t���đ�R8Ψ�3�>�
A���mX�O0s��U%p�SoZ�~B���	���k�آYƚ�;4h#�yp���{��g�Qo8��Z��	�O��x0d��kp�T@�4�r����+M����!u W%M+��a%�z��] �j=�&m���ħ&c:@GGۛ�l��u"C';i x�<�q*S{� yh6�� 4���[��ݹp�,䱄�F��t4Y�hݕ{�М	w�Jo���BHN�q�V]�S���?�9��a6 �pg��;��0'��Qb A�f�5�0��?�9���y7$L�W��%3��u$�bf�Z�AB�yA�L2l�1�D>B�<5�S�?%Ex��Mh�����M��
pS��P	8�O�(%W�c��Q��.����őv��uz$84I���E��^Ů�ٲ��dܢ��@��(]�Q�i>]�m�9I�DA*�o[��� �B���B���`d"�����|�pQ)�Ɋ�n�j
B.��,����&�<��D��t`�%��-bG��s����2�9��g����m2hM���lhQ�>1W�+:&�H� HV�>��i	��93N���惖/��Ū�k�� ��E��
�7VtZ����ߨ#�z�s�
0g��yaA�Չ���8���]��u� N��]�o���0��[v�`1�P�6wx7�X�y�CJN� �Q�����k�e���,Z�lmI��V��8s�+��R3h谱-�J�Z49��"K��jw�*N�M�ѩ��>q2v���e����^�8�'ޖ<�������d��F���'�.U0u��s���@�DS%L0B�B%S��M23��.4�4T��l41�T3s��4SJ�?��[w&�|h��`��=���N�,�pm��>y�U�ٰ��P�ǲOm���DV���
,)С�H�ȊȀ�Oq�*ĥТ"]Z0)� �|}bo䟖�}Zf��D6d·��'Rx�Iֈԉֈ��ElS<;Z z&�'��?�KҀĩ�y�BQ4-\���M�(Fu#L���M������M�,���T>�֝v4�����c�(X�%U��鲬7qlh=�3 H�a�:$�Ôx���?o��XS.��?y�1���d]�XV��Ӣ_���G���d�+s��A�8�l5�eFR �>г6ϟ:������F���O�O/@�;t]42� �;�E I�B�	N� �w@� �"��7.��Bn`�j�Fu{
X&P}\I-FUD��с�M{H�\H/F�D��Չq>��iD��%�g���a��%q�9
<�E �I�9f����L2w�ў@�p�/<��NJ9%P
 �s�<t�D�q5�]�}g��Q�0ړ@�a 	Q�\�yh�9�?I��ɽV��E�te͐m�@�蔏WX�<�M�`����ڊBB�Ya�f�R�<a��-��Ds��� �R ��d�<)#���k���+"�́S��x���x�<�GL  v�J�3$c�>?�^��J�<���7@�>Q��
 �q���ѷ�TA�<)��G��L� '�'c��q�Q�~�<���U��x1ߣH82(��N~�<�i�.7���u�)��x1�w�<!�)=S�R�K�"�DB�nTN�<i񅏧K�X�	�C� ��H�� �B�<��-<�0$��w�����YB�<��)�V���B�S�GDx0�e�}�<���Z�P��C��
D��I2�e�<�&*�6;���t�ƚc[��K�/�|�<���� EX<s�΍@1*�cF��S�<�F&�*f$6��΅	|/�(�z�<�4�[��,#ǂ9�hM��{�<ٓ�G�Fќ1����2U
�r�p�<��RZM��6!�8��@  ��k�<)!�D(m�9�B
V�n��ce,�B�<�V���d�2��_$=��ǅV�<��nN�%��!�bQ�x�B�9�@�R�<YP�S�x��Ё�R87�I��D�V�<�2�� C`��P��@/^U�(`1��O�<9%�P3�ti �AV�,���TK�<�0o	�l�@A8��Vjv���M�J�<QD���� ��wRV]����C�<��,���伛��m��ز���@�<���,#yxkF?
�2��z�<aVn�+nWnT��P#�z(���w�<� f�u(�C��#����	vމ#u"O�ay�eCi�F�;�H�#���G"O�����T�#�h��U��p��"OޘP�+&�UK5���hB�:q"O�-��ݰ�c�ډwO(�a"O��A%�ۏNp�Y��CT���"OB�cf k'�Mʱa�x�!p�"O�Y�PnK^�.Й`g��/DIa�"O�$a2�>e|
`��#ϥ�dhc"O�aqU*��t%;R�zŲ�"O�� �@�v˜Tk�.��=�`�@T"OƵ�0bV�'��	`��N)3��i"O���Vh�'#x8H#c��� �"O4<��/�H�ѧA�)sH��D"O��C�G�^X���:gY��[A"O���w�^\�(�� 42t"O���dN$����`ͅc�:$��"O���O�4 X�%n�2#��q�F"O���RAG���� ΆxB�� G"O΄p��	�[,(��0l��;�i��"Oҵ�nԺvr�����Be"O*�pi�[Z�qQ�č=�|�q"Oތ����9`����M�.�L�Q�"O,��B욇A~V�z�D4z"��'"O~4��D�A��i7-M">��s"OC-��LK����*7���(c"OܽXCh�@{���El�? �"Or]��M�'4�`r	X,B0���"OR��"E֩1w\5x�	�%�HC"Ol���N4J����@Y"�h�"O�X��-ܙ�x��܆)��"O~1iw�\i1�'!�4b�z$k�"Od��@	�3P���7S͔�P"O0���H� ��]8"�ĐH�<�2�"O&�Jk�-�(��PFP�m��$�e"O�h �OG*g��U��<r<np;2"O@�h�
Yr���1�4X�ő�"Opa VN^',��M��#��yL4��"OlmK���?84(8�b�+~�B"O�]��'��&٪��Zxl�3#"O�5#M�g�v��tL:~g^�k�"O(�F��X�M�P	D�hIةy�"OT�p�N� b��)p��4ZC^$��"O��KpF41��9�7��&?�кu"O0�u(E��z8��dʂ���E"O� Z�,J�zJ��Q��L �d`��"O|�2��@�t4Z!)�N��P#"OH֡�;�H���Q�;�&�X�"Oll� �(s* ���ѭ	����"O�Zo�Aa����		�v�"l�0"O����6�\Y���\$&�;�"O:�x$%�*����$ɾ͎��"O�L 4AZ=+�D���DE6�V$�"O�)hu)�5w����V'C��P "O�}�A�+�RP�	��p�b"O��3w��7d_R��l�Ju��*�"O�@���|�,����<Uk�8�"OL��u��M��1K��۬�L,P"O�yiNBm�fh�#�j`�"O"���J��%U�x��D�O�P�w"O��`�� <B��-�'����2G"O�l�G���^`�A��Y����"O&%��ޫ{ڒ�C�m -@D�Z�"OD�"�<l�4�!W���TF��"O� dZ!���Bn�u
ȏ%Q��"O =�p+�'� ��ƩJ7,��"Oj�����M	d�p�H��<��%	�"O���4!Ț3�1R�fF}P��"O�=��3E�$%hV$[U�����"O�Aq�3 �<��T��>jX!�$���rx��i�6n0�@�lF4P�!�d��\�A@�M60��v.v*!�ݚq"L��j�hD��ѱ'!�d�9q������#V��Y�R윊-n!��H1��蔗:Z�H��OQ�!�䈗4���1'H?�0���\�uF!�d����D��ް�Ρ0@kD�=!�D�=��4O�$t���ĊI�m7!�D\�9����Ul݇(���7�D�R�!�E";OIǅ+�$���G^�&!�"o���R�
K�^�8��%]!�d�2G�����L�)�,9��G�:!�D������Ê_�DD�q6�\�!�$��)�U틔P0\��+K�!�D�%���QRD�,B�q�R0*�!��>�y��-P?Za�|ze�F�~�!�(h6t��1΋8�*����AG�!�ai ��C "��k�&)!�T�TK�%O#�t��B�x!��8F�eR5n�K�� +� a�!�^�/%�yp"b�p��Y�d��R}!�$C�b"�t)P�ޠP���j�9z!����RY��P�4�t�ˢ$��gm!�$S�3�aa ]�o�Ќ���rc!�U�O�nŪ��^�}�@�	b��*</!�D�e�r0���AIt�#��L/(!򤚜zl�!��i N����f>T�!�dH�.� �*�I�I�أE�B69�!�$�(���cT��d� I!��?5���b.�H�j��s
�p�!�M�8�H�e�Ϗo��H)��3X!�Ƚk��L��
l���a��z5!�d�;D4���Oߎ�\�t@��J!�ġ�҈�"=l���ዛ(�!�$�"*i�Tx&N�r9r�#e��0!�E0���+70�mp���>�!�ܮE�t��L0�jl �ܑX�!�d� fۤySR,�=6��R�L;L�!�d��;\:�sfϺy90i��_�!�͎:�����g�8r ���֧�!���x"h܀s.����;K!�DO( ؂L�e ^�\
|4���$!�ĉ Dt��:u�R.m�"��ï7T1!��/V�
�.��(�ݡd��fy!�;p�`��e�/#�}���E)[�!�����;����� R��
S�!��e��P��7v��8Ucܘ;9!�dV���I�Ӥ�A�VU�Ç_/a,!�d���p��!(�R��fޭ^~!���5;�а����� q��Ǘ��!��!M�P���+^>S���%Nm!�d�.���K'�W�>�ġ�P@ƙ1\!� E�^�ˁ���.���
կ��p�!�D[)y'8��'ߏY��t� �!�ĕ�h��p2%�TH8҄C=!h�Q0�'J�m�F��s� m�����ԙ�'M4�Cw-�0s�XE�AA&z���
�'�,(;�`9^8��nY	u�L�
��� ,,����O"p�[��D�)���9�"Oҵ8s�Z�x�������>n�>y�"O����A�g.D
v"ȸ��H:�"O:-A��^��U�ӯʬ�0-�"O�4���tHv|��O�C}�ґ"O aG��=����>\�u"O�ar`�2K��qq���Ob�ȹ�"O�x�a�N�+Ԝ!�iSR��R"O����	��o/^�y��S97��#�"O�e0�#�3�fM���7%�q�O���U�{��E���Γ.z��RQkG�~u!�$��:�����T�-R>}��)[!�$�0<���+��,kJ��KU m9!�T- �`IPE� |1�=:5�A�W6!�d��Tg�if��HA@� ��W!!�C+�
���-W-0�� � �{!�d��k��I�B���,,��ܖ!򤗽`�։RP�"4& ��K÷�!�c�Fi��U�(�u	����lc!��Ϛ$蕘���0(�J��u9!�8'�*�y�@�\�A��J"	 !��-a�@�8� �!3u 񻰠��j�!�DF�;��1i1�;�H�q	
9t!�$@7.���T��P���(&�	�\z!�D�/����( 4l�6�S�H�)Y!�$v���tI�I�bT��!�Y�!�L������L�Nx��s'AQ�k�!��Ve, ���Jzd��rG�*�!�DT9	J\0:��5D����k�@�!�D�f�j�aD���Fj�)�A��Z�!�ʙQp����)0 V�J�m.�!�$C�^\2��c�	�q���0�~�!��.?�Tq��ҿkÈYJ�'P�!�$�!�v��fa����ӐiE	T+!�Ğ9 ���T%_�c��U�奏6!�Ē<Y��IH�e�>vt�[��=[!�d��,]��h%	:ai����P!�D�aN�Z�0 	N5x����M�t#�_�X�+u�L2�yB�R�?��0B]]� e�T/�y�K�f�^IBF�b�>��4>�yR0&�PK�M�$`�4q�sB�y�eN<��`��Y�d��h�y���&~@!�.N7~�Q���y�*"D��0z!�%5\QR���y2ƕ1$�(��gJ�M>�	�yb0�6���FJY� �P ���y�+I3%�ȡHҠ�:\8`y0#�:�yrbA�#6��`�%Npl��v`M��y"��:��) ��'}z>\�%�] �y2oց{��!�$�r����o��y�"V�� � ��?_�18QN�5�y�ÛRs~����:�L�h�@-�y+R�l�� ��>2�x*�3�y�C�$�����Ϟ7wD�Z�%���y��'60<I����$,��P�f���y��ǺU��9������l�v����ybl^"Y��ɐ �MJ���D���y��G
E�2���Y�L�n�X����y��7g���P�nīK��d`ԡL��yҧ��Q��l��
C�2bHk�G���y�O��*��[6� e1ȟ��y��P,M
��/$��5��L�ybL#4�9Aa�V�\���R3�y
� rܩ��L��u��+A	Z���06"O�Չ���=K,����	R!�b� S"Oi�5Eҡ]Md�	����)�<Z�"O�p���Õf���`�ƋD���@"O,���i DS��`_�c � �!��͉=�f�� �Ůch�x�,�7cC!�IU��Zc�R�.M�əH!�dΪF� �i���)8w���0>!���?Q����o��7�H�� ���!�$\�B�zU2G�Z�Ӓ�� '�4!��>
9��X���o�r�b��Z#	�!�D��!�D(� K�w�6���U $$!��^s�0��y��25��[!��%#`R�`�HϯC��`Zv�U1R!��--�1�ר4����f���E�!��^��
rH�?�X�d�X1x�!���B'�6��C����gN#T��C�!5�U:��+̄�3�^(to$B�I�ܹ��0Cj9"�,ޣd��C�ɇ����R��3,D��	���B�ɓI�jMC6D��D�%(3�V�F�zB�Ʉ{���AE�(��Dx2֭kFB�	�BABqN�e�`�p�L�G�@B�I�,ʨ����n6�j��L�!@B�	�3Z�a�AKY F�4\�����hB�I�?��aᴤ�����`�K�'�fB�ɱXA��
��qCq)G.-Y�C�I�X���W�H<.ٲ�1�*îo�C�4>��صl��d���E�%�jC�2f�����.�pTJC�փKM,C�I���(�B��*k�P2����C�_��E7��s���E��C�ɿN������9���c�11p�C䉓f|�"�*���t	`�߮z	(C䉄>s8��p�@�ۀ͙1�t��C��-!J��BpFN�rq�cl�^�vC�	)	�4ac�19�4Q�� D�i!�C�OȻu�K�/qD��(�#:B��rFip�Δ�a��hҁ�����C�I8_��9[3�T�N���(8e^�C�I�P+�Q���ͱ �!W��:�B�	=Z6� @�¶�&@���+�B�I�!��W��%'ĀsGoRE�"C�IjCR$���=*gԙ���a�B�ɨ��0y�)g���`�M'-�B�ɷu (e1�mߗQ��m
���z�B䉗~�Dx�<Z��y��˞1�bB�I�cX:�6�ߊJ�^G��>�x˓��d �I�'
n���j�Mڒ��q�Z�n��:�'��pK�+y�Ra�K�4/���#O4@�(-;$��Dk����"O�;��M"7V.�(�!΀btQڡ"O�HY�����c7� �qQQ�"O����x������Z8��85"Oޜ�,S=e�ҙIѧ �..�@���'����@㄁��94e�zX`�@4D�(y��M����4�8��`�-D�8)��܁�=���>y&���-D�z�X��P��䞵4 \ �)D�|I�`�
�=���O"��6#�<9��員V$��Bǥ���� ���
�zC��=��AD`J=_>�q��H�D�TO����^UH��M��q�4��C�8=�!򄗘`�}P3�
���S(N�A呞�C�S�? <Ph���.f�0�gÇX��W�I\�OC���kկ|�d��S�C!4����'1^)Jբ��h�J�I՗�>}�
�'�Q�w��Q� u��F�Y���'�ў�}bEfM�W
by��LS�<��C���x�<��Ǐ"T�\�s�@��p{�M�<iPj%S@�
bd�"Vz,{!��o�	9Va{�a���ܫ���敳���1�yr
U$Pn0�Sq�����j���=E��< ީ�H((�H�+�I�2H5�ȓx���бNO�0���=P�x�IX����D(�'��$s`ԑA�gY�X�asb��3��)�t��}��M�BMBP����!RvQ�� <$|��%��
B�|����/a*��	�'�<�6g�<R��T��\�����'�8��7Q�8�8�cĦ��*���'ʆ�@CV��(8ŊX-%��4��'�D@2�m�7=�����M�E:B1��'s�8Q���Us�)��'���ۓ�yr�����c	�
P=�dC՝I)n\�.D��ʲ��TG����*�qǦ�C�,?Q&��>�H<E����0( L�shZ#9oxQ���yB$O�v����#�4.]���6
̋�y��J�q��!+�*ز+Ȗ��E@��<э򤂯�BA	B�=PC���8F!�ď�$D��I�*�'.TP#ǯ��=��O(�=%>ys@o]Al���A+�dQ2)��n�`CቔSZ�s�MO�EF w_�p�0�4�Q��Z�蛕�6l܄,�^XK �Q M{��?Ɏ���/b���I����h�]8C�U�%D�$ �O����J8E̭��ϊ
n[�����O�=E�g_��*�aa��L��i�B�Q��yb�xEhv�̻v�J\�a�M	�y2+�$t��!��H� u�
��yb*�qt,����\� h�ϋ��yr�f}�%dC�N�ҽ�)�9�y�] A�T{�ۢI��	y��&�yb�P�_�4��A�y�7!��y�ለ��a(�78��r� ��y"ƌ�1a0��U�+�Ʃ"c �yR�9XSB�Bl�%M:�$,I��y�eD�MX��s��e����v���y¥�?0m��7.K-m��h8��Y:�yR�-!�Y���e��8T.ŋ�yJ��Eh�#Ƭ\����Tk��y��o� �p�R�#��	��c[��y�˄o.V1ćD 
kU��˒�(O���d��XF�itBX3pN�*�`ߏ7�!��<7��5
$LCY��]т���9�����㉴Kႌ�'��F1$�Qd�[�P<C�	7*��T	�EC�:��0x̘;5e*C�I**D:A��3�HDi��!����D.�kj9�&�w��(��X0<�̅ȓ`#�Őe��x9"
�.d�rt�ȓs����aJR�",Hm8׫�#2�L9�ȓew�9���N#J ��$g�Z���ȓ����U 8��f�2����=�N]��J�	/.��5F��)잔G{R�'�<p�f�͸J�p��E-L�Ј��'�T��ƑI=��n
G?�\��'farE�!Ȱ��M~:�\C�C�)��x� �CQl��q.��)���E�5D��IN��<��� ��"�ǢsE-�"b��HOt�=�O1�i�/�0'�0�'�д%������� ��� �)Qz)hV�1,�h� "O��c/U�#	�趍�;:`l���"O\���Ů=*�h�́�PR�;�"On��Ťg���mM� �)�"O�h�a��jA��p����h��b"O��XB�X:E�R+���su��,\O�(���PF����D_rA�"Oj�1AX��^�3���.@�<�D"O:i�1��&v�!���.�@��dU�0F{���]/�beC܁k�> ��D�Fp!�d��Ng �d�ۯN�f��0j�T�!��".���w�ʼI��@9��:%!�d��,��}paI�)�p�yVݚ�1O���$4&�Za��+\k����HK�e{!��,b&��v͋��*[6(�/qDQ��G�DM�)>Y�|S�ʄT��9�6ƒ��d���(O�>�c�j��je��n�x�#D��ue�0(��0��Z*Htr�qw#D�����ٚVxP�!F�	� x��?D��Rv�X�H!�J��m6T��!D�x�6�&(���K�3	��=��><O"<Ib�	�|����.ӓ{��H�wƆM�<a$�S&�$;g)������<��9�'�v�I�/�:E���C�i�[^��oZ(<��/S#J�נF0+���u'Jx���O4�c��u:�w�3J�uS6�ӣ:u̄���?�%�X� ��]�&�L�Q�� �'�F�'��!�'x���#&dޚ/�bA�[�hҨ�ȓ"b�x;��;�Ҩ���0��,�'Yў�|b�-ܝg�H�y��G�<�����I�<�s��O:�z��Y�})2�.TJ~R�'َ�'�۟Z�*�V�ߊ4��DX�'uXh�0�� �&���H�Yٴ{�'�ɨd�+\5�10�i�!E�\�'=�p��Ɨ�6�����L������'!.)�TOT�r�� D�
0��K�<x����Gƒ1�1��q�tr�Z:	!�$�I�4d�G�/64��8VL!���1	��fψ)F2���� k!�DE�a%j��B��)���(�,�/q�\�O�`�S����N�
|�^ j䋂��yA��D�vQ�� w�*��#�:�y�F�)k��ܑ�i	�f��U��+�#�y2�^����ǒ�Y9���2!�>�yrmK�\��)-Lǜ�)B鎡�yrD�ac�e���C6I�L���aY
�yR�H1�U��Gh��<)J�)<�C�	;O�|�:��H5Ԟ������l�rC�Ʉ
�hQf��N6�)b��!*FC�	�^�:h��F$u�0�gM��C��(�� uϓ p�H`
���"b�B�	樜�*�ma�TѰ�ǭknB�	*miP�
��Xnओ%k�3�4B�	.r
-K�Lųp\�*1�C�iBB�ɍv�Li�IH��ˡ.��7��C�I�
]�s���Sq��J̚�dߞC�>�$-f�1zRl���:ЖC�I6+G8$A��D8+�*0yc׈M+�C�I��Y�U�S6,�"�B
Y	|�B�ɜo6Ա$��<�J����֛LM�C�I�Y����v	���ř3LU4-��C�	L��С�F��rW�}s���k^�B�Iq���f�(�����(��B�ɣH��Ax񥚄%}͡e�@�!�|C�)� ���ӫ��Zl���U� z�"O.xIb��B���D�FY����"O4\�k݊a�r����ՇuT��"O¨ ��M \��I��� :d�y�"ORD+i�7x&���!�h4�Q�d"O��%e�� ��T;��m/�e��"O���Æ�{����'@��ʕW"O=)��3��FF�"/�q�D"O�P�0�*��C�Ś3
��ɨ@"O8P�-}�ueZ�Fa~��1"O�⁡J{�M�.ۯYY�h�"O��bФw�zT�AC �8O��(�"OLLZ$CG�5 \�C�^-6i���a"O� �(O�/��4�*��Z�Q��"O��$I�i�DH��
W�k�"Oέ�$�Im���ǅF X��"O)Q�b�)~�\!sv$��@J!"O�U�����CE�B���"O�"u�%oY�"$�)}� !�d"O�  �&���CɆs��}j"O�ar���\PU��|̴��"O�LZӁ�\���	N�$����"O&��% ۙp�T�aFȷ��ѣ3"O�YQ��i��d[�YRx���"O�� KO�Q���	Tu�ȑ�"O@�h�2r�}��t��a6"O�$�&�� ǂ!1I�^��"ON@#JK8t�Q@'�%^���"OD�a�Ʉ�-a�,�f�[�XV�7"O���:}�D[�#��J0�Q"O���V�X�=B���%V��8a"ODo�7>F"t�ͰG���Z�"O����-]�$��L�� 6��\�"O�hУυ,�@p�*_����%"OR����t���Z"�Lh��"O !RE��IaSi�$� �"O���4�֣N��?K��	S�"Ol�;gK�z�j����_�h�~H8"O���oҿX��Т��?��-�!"O�	@Uȍ=}`�CQ� #Q��8	�"O����\�8�p��"�Ƒ9x~�;�"OF�rr����Ľ�D��jf]��"O�=H�D7YGL�b\���`b0"O2st-��+L��5���y��(����(Vݢ�I�k���yF���8 jI?M��ɉ�nY��yR���7N`�aڷK������!�D	�oij�ذN� l͉�ӷ2�!�DS><��0�N�/�����	&r!��%4��0+J�޵�So�1W!�dO�}��-�c/L=7غ| ��U0U!���Y��/Y��d�*�o3Q!��ы+RBAamS�`�YӣcU15�!��B�5
uWG�Hx���ٵ�!���fNε�����^¸d�6_�!�dSK���̙�	x�&
���!�d�9A}�u�ǥ��i ��:��XD~!�K�R��:�.C~P$�k��o!��hL��aڐ|R���ͶA2!�N�����PE
<�l�p��P(b.!�d�>�<���u�b$qe极"!��C�)�4� ��=�n��4��!���z���C�A/�XE���U�3�!�D�x��!;���/^�������4�!�� �XC�Ί9�i�$��]��R"OT٫�k�O��Tbǡ�$V1l� "O0	3E�&�T@kᔖo�ab�"O��Q� X�>2��"�ɓ"O"�"�����U'`�� ��"O��kZ)�z��&�ޒN�T�{�<	�ć:f�堅̐�`�\�땮Jv�<�uIONaJ|`VDT7/�H<{�n�<9�H�C;V�au��6\�@�⃧�a�<���j:��	��E�.��bt-�c�<��Ңz9h��!��%? ��sw+�c�<���J/G��H�nӞHY� PQ�^�<�!�>N����P��T��C�<Ѱ�7Ahp���cU�3n�D�H�<�"@�8s8���U��2�a�	�n�<���D��I����M 䰲�k�<)��=MZY�d�2QT� ��KK�<�$����5ɒ�"��n�<!��<u�QS�հDi� �DAEl�<a�I&f��r1j�z4Ey��Sr�<��扝E���A�i,&�WD�<)&�=E���C�J�z�n�ؕ�I�<�&�:������M�B�@���C�<�eb8(�53CoZ�{�4�$eH|�<���EB���P��Ҵ+��z�<ǡګa�-��� :R\���u�<�s �!���Xp�̦u��Ik�΁f�<��Ñ*xh��� $A�t���ف��[�<�aT
?Q\�2��(-��i�gQY�<����!A��%e�U�����*�V�<��`L^����g�x��&'�T�<!�������Ä�
�TDC��OO�<1��h�&\ഄ˿`�BFjBH�<��j�R�Jٛ'�D3E�;��E�<q �#JN�U��(Os����FW�<�tq�$L['�Q��(��RN�<��ǌh'R��FH��h�B}Z���s�<A�ᖼH����K�`�`Gΐl�<Qg�	-DȘ9��+�.�&@�h�e�<�qm�87�8+%�a�������x�<�3��y��ÒFU J��{R
�L�<��E
^�u�W�Ylι��Nm�<9�N��jB��A�ȎH�lKW�W]�<aP�
"KU((iCOC ;!��P��J]�<��I�*s6Z����O�l���C�<Y �D����˖�_�U�X�`d�v�<ah��2�r}Y�K!|׮�� �v�<a��"~RMH�JW;�<��NTs�<�`�q:�XöBq?���&�h�<I�N�B���Еm���nLe�<��1?����iDP�k �d�<��V�B�R!�MD�cvl8c���e�<���=�J1"�׍a�����JU^�<��� �QtL�����-���-�b�<yd��np�B!m��!&�՘b�b�<�`�YWa%ň1�ʬ�@&�`�<9�
�Dk������=<�a��C�<��mð��(�UjD�d��(�D�d�<yU�އm^���)�%�Ƥ8S�\�<�q�V�(	���ؒe�xlXP!IY�<�t�Y&��Pw)�z7����H�]�<�b)"[��Q@d-R�}�t=�pa�N�<�4�� A\����	a��iH�G�<���&[�R�����E���x�<� \]	�n��*"���CΝ�����G"O�%�'P�9`���"oۺM��"O49Y@��؝se�4JhL��"OZ�
���Jd� �|W�q9�"O�e@� d�N�A�HޭOz�1"Ob(�r��@�*(�%�@�cB�=��"O`�jf�&q+\�Q��D�[2�UB�"O6��R	M���ţb�'�VTò"O )	ĥJb-b�NB"s��S�"OP�"�<
���A޶*X��pq"O�����(1�����-P?b��q�"O�pA�H�P@@�M��4�лe"O8@����>?�:p�c-���d{P"OΝ#5$E1'zذP��7*���"O��2ꌳO@f<����3.�8UA�"OlRq ����,�#7�1�$"O�L���ܘ\���ؖ�U���Ԋ�"Od-X`o��t�^9pAj����}aQ"O�!�'��3R�B�^�<�"Oh��v�R�6P���GK��J9R�"O�X�7L{+rq*�(��M�T��"Od5Ȓ � ~������#a���8"O�Ah"�ӥǨ�@G͜w�)�"OL
cd)6 ��F��)v��8�"O`��W�_PqFPz@}��"O����F�?�H��pC��L�p�"OtU�' Q+E`��v�C ���
�"O��FΝZb�����ɏ���"O���灠=�0$(�OբV���D"O<L1%�(�:Y��$��6ʐ٢5"O��B�]��b�#�B ϛ-!�;Vd��yA�B�-L�r5mV�!���6l��IH�gX�%;B|��Kh�!�D�0��d�t �;[�Hm�ѩ� _�!�D�9o�� ���v��<r%#^4!!�T6<�0YU�W�L��*2"݅y�!�ñ�X����4[�M �C��]�!�E3T|#��<^6D��#2�!�d���0��A�[��[�A�Q�!�ԬA��٢#¶F�b��a'\~�!�R3f��ȗԦ5�4�O<!��ɏ^��T`E�H�mߔ�`q�̋;�!��
�!���>��m!-�9U�!�ĘJ���fǨI�K��C9b!!�D��~�L'oN&�b�gT�{!�!��T����&R�!��X�S!��XQ�����ؠv�9I���r�!���1>w�$ڣ�N� ����0f��!���=I�>1M��jU�u��.B!��Y-�b}�ta�t�25�@�{!��EN�В��H;D���C @�8$P!�DL?}�H�dJ֢z�~4�׮חJ�!��*{�
�bFT99�`��e���!��*�F�
�
$?:�X�,�!���!YP0݋��Μ���9���!���m�@c��X�O��-0W�2�!�[�S�f%��F7DJք�P.?_�!��4t�`C���i�,tyōP6g�!�ğ�5�v(�*ݷ ���C��F1q!��a�8��>K]*�q��*v�!�d��fXb5炪$*���E�!<�!�	'J=6�C�]|�`.0h�!��B�Y$�yu�L*F� @����h�!�І$f�,!�U�,�JvG�-X�!�� �L��杪O|�2"KV�&c|Q��"O�c�e .a�d���_ 0����"Of!Hv���6!��/�.��г�"O.����K�z+Z��-]�E��1"ObɛR-�gF�����`IХ"O�#�)��K}$R�
,�\3�"O&���$�J����D�z�ف�"OL@i� �,H+�)�#c�+V��$"O�i0�ۙ_��raA^� �S�"O�����R5�`���*v9�3"O��+@"�|�� ��ދ[T���"O°0 "�{X-1uȁ�]�^	b"Ob1ye�9sS���^��I�"O�� c���R_:T"�G�+*�vP�!"O��!EKy4�4P4�����{t"O�iYa�'G�h�Z�e����XxT"O�x��\2�K֊�7}3&��"O�,kfA��p�E`���1��Au"O��#���8Y2����ӾV����"OF���H����b��I�Rg"O@J��EP��|�Dj��P2�aG"O�M{��>6z���fƼ)!�Z�!�� M���C�,ΧJO\e�Q`Գ\!�K�@`����X�<�{�ܞsw!�$_8ּL���H5���!��=�!�$M�0�l��B�t�n�Pc�ߗi�!���M�VQ���p�H� d/q!��L�N��x�I�1��Ը`��1#R!�ɪ$��P ����&,C `�m>!�Р)��i�Q�J���PϚ:�!�Dѷ98\�`Z�=����n�!�D��9"��}O,Q�3�@1U�!�[���0��:[d<��+�?�!�d�8�&��^8G`��d$_RI!�Ė5�%9 �VFp��"�7f)!�$�X��8e�@/یx)a��K{!��"&Bd��q@�_��}p��7�!�h�y5��h��@:q��Z}!�N9�tH��8>�d0r� ��IB!��Nd�"u&;nIs��GR7!��2? l0��M�h��aX%!�B��8��I�~�J�1�_#!�d�ꔬ{��ΗP�"ȱ�K!F#!�� ���!Ћ��,���g*�2!�d��.<��"M�V���a�߆.P!�x۸T8B���+�>�Rr�ÑN!�D��g�a"���O��D9�k��o�!�R�*�BlQ�c��Y۔P��+Kv�!��µ<���/�T�xB��:#�!�$�46a�}��%�Q,��Rj ��!�d@U�&�¦W, �;4d��p�!�dD�0��p�v��U��R�9!�D��%�l�Z�Y2F��)����G*!�D��Z�=k��ܴb��P�s �)!�ɀ��aٗ,�S�T�#��A�!���F�~8S�-�1���Lۆw%!��Ҩ R��SM�i�8*'�U�h!�D
<Y;L�	X��RY�3h�7�!�P������d2x��[��R�N�!�İf�K�LDA�P�kd`��!�$�pU~�����R�k�/�)3�!���)�إ���(�����̏I�!�dL,n��C��0�������~�!����n�x�J�[���: L1!�� ,���%
8j��aJ�7�z,��"O�!s"@E�S͌�s���Ĭ��"O��03��=쳴� �@Y�"O���W�OUd��ӷ.U)8�6"OH�c��e��a���p� 9�"O����(��z9 ��#�zH�f"O����L�	�`՘12=
Ӕ"O��H�l�=2x����)��+.�)�D"O^4�藕$[��@#i
)�h1�"O!��ӑx4�-��(�-un4z�"O���w��;�J����ݓ	a��Pr"O��ꅊVA��Y���Xdj�k�"O���R��&~i�ڦ#C$z� m�4"OD� �"�'�,	b��!lt���"O�8�'n�3]d�&�H~eXu�2"OL�6%��`\�)�D+A&~�2���"O�	�pg#/hZ�8�d��A����V"O����P#0��1mX�1y���G"O��K�]�v��b��DY���V"O*�t����������;�"OFU�𧍟��q��υ�b����u"O���-1���/@<��`��"O�DhF
V�s���t�+uD9c"O��>i�$�a�(^�=�&"O�T��h�(\�D0�̆�O6m"OH!!�&�3-�9R��\>�p�#"O}�Q��,r.8͢�F^��"U��"Ot�-��}'&��Ţ���߅K5!��]��ᡢdHPR����hV&�!�d�2i>y(�.�\�F�=t!���h<$�*O4
U��5-*fs!��,�R��W`�F9�а�FY!��%Jh,}�1H�q+��Z�F�!�!򤕍�BlQq��+K�F�y'��!�N�P�؀�rFڂju���%b�!��X�69䁡��Z�6����P(!�D :j�MidCD�E�P�b�=}!��2M��1�!@M)~��Ժ:!�D�3�t,*4�&�4���Đi�!��ƅ*�UR�J�,���d��!�$=�%`��C����7�!�d͸�N�2#�f�`P��,�!�dK:^�;�mVz H ��؏c�!��5	�(A���
��%Ƣh��'\!۵g�8��=��"�!qO|yQ�'�@@r�ۘm<H���R�d��Q
�'Ԧ� %��7^�j��B�_	v�3
�'<2���� 螁�`�1S�H��'��{��mښu�'GB�{����'��+2h���1D�m�|`��'`��4ይ7{0�L�mdʨR�'B"�����Z�L�GL�l,���'3 ,���Hp/�,����f>���'=���'LQ!� }�wj\��0Eq�'�(�$��^�|��Gf�>���2�'~X\����1�RD����:~���'ߘ�RB,_�AΆ4!L
�'ٰHsgy�T �/�(oc|x��	/D�x@���.�01�O��tQH��U�:D�8rE1z������x��u".D���1K!'lp!��Q�EN��Y��'D�T���X�[��q�@ϐ6r���$D��I�k\N�����1s�hw*6D������yFi�聒J/�q�i&D�� ����#�%8�b������B"O\5�r�C�8�0[f�������"O(�i�l�)-4�Z���1p�]9v"O�qXѬŲ>�p�b�i}f4��"ONp�E���{��	��(�o{����"Ov�D.��[��x�gJ�bcha�a"O����G�����@��/U��"O�
�C�;a�ƽ���G6K�|:"O���4̋*��!@!��<6����"ON4�0E�gx]����|s�"O!��΃�H��c�L�s�& ��"OL�[1�	/�A�Ud��Z���#'"OZe�2F�kz2(���U�z� �"O��*�o��&X �ƦO �@��"O 3�
�0(��(�2�K�$�=XG"O,�F��&�FPҗ*9JA��"O�d�1d�LȘ�!�904��"O���GܢL���Aצ0H�Y"OtY�A§s�b����1[�"O�Yفk�	'F�1��3=��,K"O:�a0�M,`����^9��S�"O<Ps㔡��0��˿1��%Q�"O�� ��f�$���.\l`p�"OL 1h�*>t�t�Ŕ:�|��"Ov�@��ؓ0�ޭ�R
D.g�^�#�"O���%�%!V� ��Ë�>��"Ob��#9�x�jrH]�	z��"O|�B`nF @L8���h�Y`�"O���0O��I��鴃�I�D�s"Op��mh��ѡ�^2���"O�(���_���X�5���S�"Oʅ�k��H�B��:i���#"O�����f�53��V�|���PS"O�|;, ~�F��r���t`["OLaq�{Y�1�k�f\��"O�E��>-�<��K�7���z!"O�X@�挽2 h�jU>1���c"OP��Q�ڃsG|	0#���Y�V�Җ"Or��vi�/dp�w�Q�^:|Q��"Om���܀�D�5b0���"O�A;hN4��x�q��Z��"O�M��D;G� ]���I 	���2"OV!�Ƅ8@W�5�7l�+N�@�"O �'��H�R1�$��u��9x!�DFmd�1!ֲ �{U̜7nl!�d@���u�D��)CA��3S!� ���ـ`Z0.��ʄ7E!�dP�l�*�B"�35�40�7ʉ�qH!�Ę8�l��EP� ��I��fG!�Ju.,�g���(m�C��W*!��{���S@h�KJp����!򤆵H݆��1�Y�r5`��u���3~!��Y�)�t�Q�k4a5�|`6�C�!�DT�Q��""ѬV5�Dᥧ�&2i!�$�,G<H�
�
<k5ӏ(8!�D�*k�E8֥(L���+�*�65!�df��Y Z�Um*�P���!4!�䒖2Wސ�7��	a�x�0�#!�DG�$<�2��ݕ$Wj8x�R6!�D�63����ǅ5����a[+/�!�dC�=fUۥ�n�����'ɓ$�!�d� !���L��~��Ҧ̉�!��5�T}+.Q�0�s�H?g�!�d�U$lЬA"�Z�����!�� z`AG�J"��i1�Ȏ>fް	p"O��*�b���%��\�D�@"O��������B���d"O
+	��v�P�!w��b��Q�w"O����m�nv�X�!�.C�h"O�L3 N4b/�]��%�/m���$"O�0S�#ٲNРD�@��9In�s&"O�`�C�0#L����T<#Ԉ�"O\�K0�8(�D�U0��"O�Q!�A�[�E�ݝWh���t"O��0�W�=�� 塛.I~�6"OFlX����f]�AA�RA� 4"O2�h�'ɪ�����M�)J�l�"Oh x���8m:��ÌʵD�AAp"OZIpe��f9�%�;#���{�"O$�3읆~j��� �
z.�"O��7�!(�\��B�.]�G"O��	�*y�r|�1ס���$"O���@E1p��2(��VZ6�8�"O����]b��mT�� ?�|��"O*U�4	�#[:@!z�.�_ V�K"O�u�f
W7o��L�ׯS���A"O��I&}N#��h��9�"Ot��H�{���Z!�ɑ`UNA��"O��E:^���M��a0����"O���`�ȾK����K�
��`HV"O� ��(D:{�>���(@~��y�"O>�؇l��U���W�H�O�"O$]�¦H4I!~Q#�� �<i�"O�Ȃ��p�Z3"���tެt$"O����+2���t� !Ъ�b�"O  G�>~�PsT�W8aÀ��D"OJ,����`z0���:{�$P"""O������"�\׍̡qxZ-��"O<�2QD'"T����؀IQ6"O����@�tdty�Q�h^��b"O�Yk�'�W��A��!��D8|�	q"O�a n�4u�L*Q�A�r�q!"Of�B��n��T��)ĝ {�"�"O�����J?V��I*6
G6c0���"O�����92<U�R� #���"OVi��f��)P��6��tq"O��"tf�C��"NҰ!�ح�!"OU2sf�eǞ�(����ls�"O��;�$��ob� �dj�9-F0p�"OV�ɒ���Ty�⑞C
�c"O�Dpr� �dlK�.}�j!u"O0�c�ȼX8��D&�;/��;�"O�:��)|���$^՚��t"O��f�����hk$ǀ� �Z�J0"O�УAYg%t��F���a࠘؁"OJ,	�AQ�|��pن͆.}|��"O�8�������B� |Y�tq"O½��M�We�ԺPlV+R��	�'�(%r���+����t&\/w���'Y���2�&2�����	�"M�<H�'�I���o�<��� �i��Xq�'�Je��D��\���T
���'�����E�#3ʤ0�C�[�b28��'�ެ�f�!P���@,�T���"O�X���W$��Dy�șV��("O�-�7�O�/P�+�� g�x	{a"O
X�����V���cK�Y,�P�"ON�0�US�@��q㝡"c���"O� �X�b��*ٔp`uK_�t�ĵ� "O���7�[� E�#��֊U�L��"OJ40gU*L��Bσ7Gv� 1�"O4���M�g�6�S�<,>��A"O���$���D4.Ó_6�,f"O�` �H�n8����+l;'"O�!au�I���+�� S��(F"OBp�łc�0��O=��E�""O��X@�*X�-�pA�
NY�"O����'w�aH�`H�0 �"O��4$\Kݼ�X3�Y��0L��"OX��Ktcd��LR>��xd"O:t�U��%N�l�3�Nݦ���u"O���b�8^�T����R�N��YG"O:�8��]�{U��#"R�-����"OtmJ@��x�:����$1=��)`"O܁�bd�+Z�z�����A'M�"O~�J��=Y@�O۳~�<���"O\�Bf�ڸ��0���,�d��"Or�٦g-,�	�G=�2�Yv"O�����jj��$���$P[q"OtUSwk�B�1��$��(�0\�"O<��Ҁ�$CO����b�ܰ��"O^��2M� F��R+\����"O�0����\��l�3��5C��1q#"O�0���k��+���76�Q"O���Dmɥ4|�	G�	�U.x)�"O��NU�F�� ��I�D:�"O����Ύ�2��p�DJJ� ��y�4"Ol�y"�Y!�~�:��^D�����"O�����2uGuk��X����"O��(�@_�z��t�	+t��"O�a��#Yp,Z@�,zU#e"O$�(��	Q*�Њ�.
T�h�C�"O�4YV\�*�����L��z��0�"O����ȓ�	�"|�`� p����"O6�)� ��f�> Y�古{���r"O����N�?h����Sdظ_���	�"O֍z�(N�7���@�v���  "O����\�\�� {U�">��qI"O|����2O�p��ϓ�6e��zc"O*<{E
gX��I�.Ͷke�Ě4"O>0�F͓�i?�h�-[�^F8� �"O�+�.Θ�쨒��?Ǯm3�"O�Ea�*ҵ|m�h�v�	�"�5ja"O4���b�&@�E����0���"OTa!t@��d�\h��*�Ub亶"O�x2�-�W�H�VI��4nU!g"OP���Ƥ��G�x�N�I""O��JP.	=^�Z|r���K�X�!@"O�D{��U�i��e"A�h�(�JA"O^���ã*�}���W�M�0qv"O@��
4@���k���25�Vq�$"Oq5�&y�|`x��J�u��"OL��t�ٜH�Z݂�X
6l�Iq"O2ѱB�Q�@��P��A�T�!�$S�2xr�#�,�&Z�̈83��$4�!�D]&j�Vi��
�����*;F{!��`��<�5�Hx#�IC�!�f8�P���&��3��u�!�K/lȘ+�e��ɗ�@�!!�,Jy0"�	#C���נ9`!��Ԫ9թD�"nGQ��lE�v!�S)������f��`��̦F�!�� �U�D΍�U`@�AOz�\�"O�h��O�$S>�	������1'"O�	�tb�/P�9�*�:��	"O��W�g4�:gꌾ��q0U"OD���KĿ`M�fi
�*ip�"O6!�@	K(29�Er�4�`X��"Oޭ����$"+J]!CD
�q%��G"O�D�Ռ�-�fUQ��� C4��"O��FI9̔��HėS����"O��9�/�
d�x�2�#	��	�E"O�u�F�M�ibfE��h�&\�sd"O]���	�䥀u��]j�٠"Ol�q2*	jR*�
�
UfK�	��"OB�q7@��R�z���iKzayf"Oؼ��yGH4�(L0`1"O$�	0cʀ!iR�*�M���5"OfIq� 4M��Hx��N���'"O�}��%�2�^�X��^�N��5��"O~��2��##�pD�$��E�|��"O@y�B��Ɯ ��Ė�_����c"O��2�ڡzm�5���O��UC�"O 9u�U�$�JDⷉX�p�yH�"OX��&D��g�4	"hҨC��dxC"O:�A��F�9@a����`�VP9�"OV�b&ʌ� ��vŎ�sB���"O����@� ��EU��;xtm�c"O�B�ʪ b8|��� �^,�"OJl��^Gh���%3�T"OJa����3_��I�g�
N��͂�"OD4����"4�#���{����"ODd��	BlMU�%\	a��ph�"OPa(�*ע|����C,e��"O�h�4�L�$R�`�X�d
a��"O�J �	gA�5����1Vi���"O���� ��OR�806G��&0x�"OY�+[
�;È���01)�"O||���P$A�ɰ��4-q��0�"OJ�1f��wtA� 1ZƖ�r�"OD�)��P���A�����#"O��ѶcL�]{�����öK��\xw"O�b�������mH�
 �"O���/\���Q�kF�7�x�R�"Ot����p5ƔPW����U��"OT��'dI��h�)p�� "O��ө��B(0e��w�f� �"O���vO��XwL ��-$��=�7"O6|;vMӉlH�#PR C�9��"OJ� ��o��F��F8�"OdTR��'C�E)�DS�`���"O���g�F�M6 �#	�K�ar�"O��┯�axv@��M^1xa2�@�"O�H�B��W.�եVK8$;�"O\ H�$N�G�D��b�:\is�"O>is�D�/+\m����38����"O,����X�hҘ{�%�8�"OH2��PZ&~��wa�!_����$"O��GHG9SMnLa �U�5���5"O2� �"�/Y����寞� �&%g"Oؕ�3�H�]�ر�-Z�}��l��"O�uSp"�D���� %v4x�e"O���!���KbP�3�_���{�"O�XjEfZ�2��PR��U��YC"O
\#�"�p `�X����"Ov�C��^wF������n��"O� $8¢#K8��y�iL+w� ݣ�"O��oҏ'�V�����J���t"O0�el�#�����"T1	f"O��P�/�p��#q �bv�F"O��84D�$2����,G��<�"O~�cu�{J���kS�M�||r"O�@-� J�㵩���l�V"O�PVaǬA��� �
�27c���"OJ��i��,u��+b��7uF��"O�\�4�'r�Li���G�
/z�IP"O<A�qA�-�m�B� 8^!,��"O�M ��V7��	!<���"O� ���#u�6 ���a���:�"OjA�+BI�蜣`�
Y6R1�"O�P1a�$�(��vF[9j()�2"O�����6�Ȁ�U���'���"Opಬ+V��Ps�W\:�KU"O��K���m'X�2u�VT���z�"O��"�ل��AB�H�l���"O�IG#��\�LL �5�(a�"OF���b �4��a&ƦX?�%� "OdP��F�W)���G��,Fa�"O�x"̄�d�Ac�/Q��1BV"O ��*�څ��_?S���"O8�B���|�d��+�H�F��6"O�TYCSw�D��	�.>��,��"Or�����2I\��g�v���"O\]��㈣<���E�8K��t��"O�y�7LA�HⰒ�#H�uݤ(��"O]Y3��{ �	@� �:��)c�"OJm�磓%nd�aQ#
�L�;�"O�h��P"L�V�S1���(�p�"Oް���/����n�8�`�"O��o~T��dH!�p��"O^�)��J�D���U(��Tu��"OҌ3䤐�D� ��FW�5n@ �w"O�r�۴/�Xmb��@�N���"O�yc2�>�ِ�#�!{�r�qf"Of�QGıa�5���-G�J4y�"O�x�c�Qk� �3N�� ��B"O��C���gq���b�>�8�BC�	1%��sP$W,}�b!w��!-�fB�	�x|f��jɲ�~$��AKD�&C�I�E����"+_
�Bl�t�ޥ,��B�I�XΦ�����
��V͘�C䉉v��<���'b>F1��E7�C�I�_��h0r_0X$ I����B��C�I�b��X��ĉ'�$�@_2_vC�I���4.^1 UL�Y����TC�I�w'����-��I��]C�	uRDCSn�5?3��zu#�dc
C�=���C�R��z�G\�[B�I�,\TQ�"7�rT+%O�$=�C�7qR��ԜuN�p��]	-�B�I�F\p����N6*|�䊚>�C�		.q[���:;�ܘ�tj�$E$�B�		^,��㫕�[N��B#O05�XB�*o��� H�/}*��B�s�0B��	_q
MV�
Ik��"T�4B�I����`��W�����:)LFB�h�R��(W��`��>
B�
Ǝ�B��Q
x<���h��k'�C䉪l�����z�G	Yc9�C�I15*X��ä�0x��"�>Zo^C�)� ���P���T����Z���`Bs"O�P*C��m�{��%r�b���"ORD�R.L�P��S�h�6�r��"Ox͢�0I�;��t�� 4"O�(a�E�="�e�C�߄�j�K�"O(+G@�!��E� J��k���"Ỏ� M��XH̐m� ��"O�ɲAϽd�*�F� )�|{%"O:Y���<&�cB������"OLc���
CQ��X;"� Â"O4���!8X���@cQ��q#'"OMCD]8���!?c��`E"O�x)�K��kҠip�ͥ#�����"O咳jP�?~TY;�)V�J�6��"O�0�ZU�btO֕!���"O�]C`c]�5�m��� ��@��v"OpA��d��qz} "l��.~�ۀ"O0l���?�ڼ��îT��SC"O�E�f�$\B����<;c� pv"OjI%� "{��tӄ!�:]G�8�"O��KTB_:ZX��6BN	9BL�P"O�}��h��>����!����"O����N�1f�p!񁀈*x�U�4"OL�
B�Z�<��ؼpm�IH�"O ��'C�6;�`��H�R\Q !"OzTa�B|<&ȳp���'&�Ei�"O"x�UkX�Ay�ekf�i���+d"O���$B��F{��z�K30���ir"OdirC��Jl���rP��x0"OB��Ɣ1bπ��tːxl�;�"O�XW):[V�-��
�k�^��"O�՘f�H{�l	"�*[�6�0�"Or1��������IՈs�0��"O�)�㬆>|U�1�U�"��e��"O2���AR�r
:� 0b_�;�"O���ũ�I`����3h��3"O�4�S�ؑ#��B�����H�:D�d8Ԫ�-"�!�I�=��9���9D��2Dˊ<Ǥ�Y�PD1��*a�7D�l�g��!p�<"gǘ&'9lIP�g7D���~��o��ne��E9D��է�2\�)Bă�=1�b�8V�;D�p9a&5��*����w\!���4D�๑F  w��x����8�[�h(D�`�D�$eG�=B��2���$D���N76�KӧI�q$� D��3E��	nb��3��V�{���2b2D���%̏�F�\]0�`6°u2R�"D���p��3Mݔ�0��%q����q�+D���&m�".hA�
��1r��S�<ɴEF	[D����M��9N���v�<9�(G;+:NmJM�_v���
Cs�<i�d��n�h 8�d�֞�H���E�<A@��c6�(hb�[�1��A\Z�<рF}��dC��_��89E�U�<�����R��uk
�F�>l#q�WP�<��C��9XĴ�v��3-��]ۡ��L�<����+'^<�F��MfQ��SG�<����8�
�Q��7��Ү�C�<Yf�3`Y��p���.	�0�R�AEA�<9w���>o���uꏫ#�>������<�G���>�ȗ�$p��1�f�{�<�ՂN� zd���lH�ʕ�u�<I�E�U"  �_--�d82i0T�� �tb��ђlt�(�M�� �"O��z�DP?6���"��:'JF y�"O����M)�}�ʌ�:��y�p"O0�x��Ȫ@>h�L�6	�"O�XD�l�yC���:l�,���[D�<��[1�>;�G�7`4�ZC*�|�<irǫf�,#��5#⺵��|�<��ݖLJi��'����4�v��~�<)��G`�Ե �A0s�=��jo�<�ԥ;>2(q��-�,�d�#�!�b�<��ܮgr��#n�K5^��2` D�<�c��8�$I�n w0���A�<�p
У���Жl�*��X;&�~�<�E�ӗ� �hH�PG��aQ�Q�<���Z
.�F�W��7�8-���O�<a3�\ 0���� .�a��-ȥ�W�<JW#��5����]p��Q�<q�	'���jQ���jZDp��K�<���^�?�85����(@�h���R�<�`T#���C��W�\����LG�<�����>���RC��<��� �-n�<I����-W�<�G��X%����C�<���E0/�m@#�ǐ4θX��E Z�<a��@Hb+��^Y��=;fDX�<�F��$tr�bKK��6s_'!�\0(E���@�Z�|���kY�t!򄚋r�D��Q��5 ����򊂔a�!�/aj<��aο4�l�a��R"Yv!�G,&�����E/�K
�|S!��^?���;�K�-8%�s��;�!�@;zӠK]�F��*g©:p!�$,`A�İu>��lR�2i!�xxA�#-��h��hĪ�$�!���7q�T�ĕ��h��(�!�d��}Ȁ�1R�ґ͐(Rp�J�
��Ā��vc��c�V���� �y"\�K��D�¯�1�8�8ӣL��yRf�KN��B�~�����J�yb�Mb���I�
f�)�U�yran�&�ل���#bj�4�yҩF� ���ram�4Y�&��r`ń�y���<���Ц �)B��yr`�C�j�S4l_�s6	*N�=�yr�ޜ-_h)CT L?�i $�yb�гb�:�[�A�ˤI�e$�7�y��'j���;�8C�h$!ތ�y��H�����P h�L�p��>�y�	,5���qf��X�s�؛�yKԜA}�=� ͝2N�L`����y���Y^<��b�.֠Iqp(K��y�.�+"��e�	<*l,B��:�y��9F�Y��g�E.\j�lƕ�y��ϖV������:�KQ�_���ȓ��TI��Ұn��l"�42���:�Ae�1=��Qԡ�9"�ȓ3��Y��J�@KnU9��^:;��ȓe��@�eꅘȦ����Z� `����h�J�,8��	���եq�"�����-EƇ�4��&I $`�d�ȓ7��HcS�K,Z皬��=W���� ��]f��e]rp.�5CƄ��7�����%�����S05�	�ȓk�荢 �F.A�d=����x"1D� ���մ �ԁs���>�H��d-D�� ��)u
@�5A�@3�ƝMtnP�4"O`����¸l�q'�%��P"O.�5��r��<�C��G(X�"O��8E��	iT>�Y@��ZP�w"OԌA��V�[��=;O�|�~ub"O��P��<lZ$ԩ�Ζ�k�~Q��"O���Ɖ)< j�s�K��^tA#"Oؼ�W�J�5
��PV�`0ѳ"O���%��k4EӑGB�e��"O�s��C-G��k�5nʰ"O��P"��O��i �� ?V���"O��kЁ	 ���``Y=��yRe"O2`��EC\��3D)�� �e"O2DBqC��c�ұX��"O�yHp�	��d9A5��)V��E�"O��#��4Y���V(��$T:5��"Oj�����fC�Y����V"��HD"O���sdT�zG"�� ��&hε�S"O�I;�M����B��->�
���"O���Fa�#�tH;��)HL*�10"OR���!1�&̙q��e/��ST"O�T�L��+��R8& e��"O�5��Z�R��`���81�8��t"O�������H."/�
�"O�b6c��A��n8`r�z�"O��H`��\��ԃ1��p*��"O^�ce�E�d���q�;(2��*%"O����V�\�"��".�_ LQ["O��L2��,q1��7>�ha�W"O�(s�6Sbfx�H�h�6)*�"OҖ>$2�)E��� ��LK��y�I�f"UA`-Y�zx�R㚀�y���\��<p��ˇL���Ri];�yR�ǈF���@0.L8��1�AG��y2\Z_��3�bM�b�xe��y򈌦A�0���F�oaR�*��ԯ�yȚ�X2z�#&�ѿQԐ`���#�yҮؤm�𹩆��N���u�P7�yR�nf�yCW��rnd9���-�yZJ�u{�n[�W�JE���B�9e�D� s����cMը(�vC�	�)=\�J�56AH�6���dzPC䉵m�N4��рqTܐ�da�-#FC�I���0*uΚ,\^|���Η[4C䉧#��|2�ꉅ{�e �m|O�B�	86KJ������H �!�9e�C�ɜ^\���OKC`�]�2�	���C�	0a���A$e�G$��Xa��|0�C�I�|����ʾ_�V�j��<n�C�	 $B�ٲ�"'�	#|zC�I�X�V�YAI��f��@hSΆ7�tC�	�'�̹c���lC�T�UNF�U�B�Iw@<�[@N� q�h�� ĳqJbB�	��B���E%��`�3���fnPB�	;?�u�E�+?@��)��B�ɪ9�6�!$b&~H�l�"��!�C䉩m�P]p���A�D�Qc��zC�.=��NK�Y�f�� DL�V{�C��#5t!h�i��kZ�iEȏ>B�C�I�����Ue�m^���uA'{��C��X���Rv�бT\���q�T-M�bB�	�[��t�ᮛB���;jN
L�<B�	 7����q!�&c��1���m�B�	�?��4��C�BlxUb�
�"ng�B�)� ���B�Ӫ	��x2�B1����u�'�ў"~�j�)md�@$�M�t��d8T��=�0<y��dY�Ep��P��7�:5Y��Rz!�D<b�E)J^�A���������D�<ɣ�xJ?iy�O�����Ҡt�;C-�MN(�p"ON)q�ֲ�8
`�ˤ1?@�C��$Xa�$���\g�rw΂>U"tA�1Hޫ�0=)����<�ZFA��T��A�Ф�y��ϊ�0���"1;����@)�¸'�ў��(��$�u���y�E]�z#P�A"O �D4f(2I) b�4��S��IYX�t��HR+ksr��Bg·"������5D�4C�I� �f�0��.L�]An5\OJb�|a�����6T�5A�/�pA O7D���� �$�2$s�����Sf)D��!�B*(�hx[e���d|�����+D���b�� _Z^1r�+�';hx"pb-D�	���#�
�㔃_ "�B� s
9�d;�O����,8m��lŷX���'��}t��R�O"t�<�kdd�W�!�\�R�4�ĥy�n�xD��m����E��*ʘi��2�b�N���Z6�Y�U��B�ɵ[��m�$��s.���!�kTt��hO�>m"�B��Ql����=��d���"D�8�A�:�9��ѐ^E��0���XE{��i��=�ni��"X`a�%�?�!����&Y��Ҥ7��� Do4!�dAh�����ٰx(9�e��D%���lӴ�����,�� ��!���8w"OF�T��X٪u�v�^6-�D�
��	(�Q?�	�MżOÌ@`g�>5�����3D��Р�Bna$�Y�^C��J'\O��=�0,�Tk��N�Q� �	gNJ�<�Q�A*�Ek��K
_�P1s��E�<�&�J,6�B5���2����CC�<1EZ�2B����H��z�R�.�|�<��)�H��b�D��;E�v�<I##% =>]
��U�sѶ�(�+:D���q叺/�����FR�<m��#��2lOZ��J>���ϫ<���;��I�7>j��FAM`�<��˦�ЁAů�L`LMI E�T��7�S��'4<ȀB��;�FA�3�K�B����_��f�;�}������=��O��蹗`S�4&2����ˌe��Y�ȓ:+FuR2D[]N�1��$޽yD�EϓԸ'%�x򈋲P�Z	���" Q�Q9R��9��Q�`P)�}�����'=��3&!��t�P�"��P "O��s�Bڕ�j�ر�@((uk���OD��O����d
�#.����H�G���1�	4���u���F�GŚ���C�_�2����t����I;O��rbc׶G_
��M{=��hO�>�X�K@�	$Y�㊞:�p�6�/D��R4τ#|��,��?�d x�,?I�4�0>i������ШŔ*��a��X�<�&K�g��I���	~�%�e�R�<�&�ܸ]o�4�^*TZv��nN�<1�*	�¡��G�&�����T�<��J"3�z�q#
k.�.PS�<�'#V#Y� d+�� U���9)�K�<�S�פU:� �A�27�8}!0�LD�<1�(A{a�sa"��L�^����@�<1GHO;j�X�H���:_k�����d�<q��I�n��&D4v^)�O^�<quo!�4CS.(�Xۤ)Ca�'�ў�g�? �NO�.�b���J�6V��q�"O|q*e`H?�d$H�8Y����2D�`X��1.k:3�g��k�,�@)/�	ey�X��O���7��и�̄7A^�A��B�]�C��8����)3TS"MV��,�	l}r�O�X�ᓕT!��"e��Ta8Zb,���2}�ʛ' ^��t�I:&�,� �G��y"g�6`����
�;iҨ�q
 �yr�� .����P�3�� !]�eġ�E�V4�|�G��H�4)ز��%%�}���q�I�/��C �I*U�P�į>D�l�F��j����� �6l a�(D�,)�(�?��<RT��+�ℌ'D��# �NQ8�:���_ޥ�"Ɔ`�$?}��9O��Zg؟A�����^�@���h"O�9ȑ. �@^���U$ŵ�(�c�i�֓Ot,��I����"��|1�j���"[, �8F{x��B6�b@ȵF�!ɦ�5�yB�M��@BL��D�(�(O@�=�O��S��IV�BP��8D#\qK�'u�e�2�ھ.+����˜;��d����&�S�Tm�42<���
1�%H���M�w�)�禕C%N�S�0L�ϞGZ��)D���7K�*�����^�P�x��A#}B�)�S1��}#�MB9_���r�������/?y'�Ck��@�bQ����;v��x�<a��A�Ly
%L	4���$�_O�'O��D�O(���F'6i��wX��
�'̠!���[�U@ȸ�%
�8%��Z��d5�'3�Z�K3�ڀ���i��E�ȓq�xB  �:0�@�mC�8�ؤ�O^�=��D��Ib(0a�3�.�zagf�<AŀA�(��}JSd:z���ъb�<���"I��k%J��7؝���i<���%��̨��	J	N�{�eF8FT�����v�˴��8�,�h� ��}44�ȓ/��!�W ����8W�Kx�ȓ"��p���2�69���ک���%�4��I�|i�H���E�Qnф��C�I�hJ| ���5c����Ǡ�%1�hC�	��@p�ͧ��к��ޒ^4��?a��)�7�¹�R�K�I�L34��!�$�9L�X��ʃA<�X�h.K�'��斢~Z�ܯ#����K�Æyh��XU�<1ю�w��}jU�W7��{Ef�M쓃�'6�I(�y�	�
=�z�J�.H�z�V��Fh�$��x�$_37I�%{I�O��2V��N�*"?Y���kr�s��^�!	��C��nw$B�2)� ��Ĭ�4��st�E�7Rb�i�7H�8�' �%��i�&n]�h �̇ȓ7�H2�����2h��>ռ��Oz��D��Y��3���"=J�zg��.d�!򤏳:��8Ĥ�:9��KDØ*�!���Ff$�ٴ(�;X(��pRᐯ^�!���
MG�H�C,'6�&*	�M+!�C?�.����9K$r���nۘG���hO�j�_X<���U�q��b��'�!��V�J�I���Y��`�uN�V,qO����Y�6�J�J����x`RNMX5��Dl�D�p���7:�, b֨ )��1�d"OT���`�r�ʭA�5?�Q�"O���FeL�A]*IQ�Y )�	�"O��Kc���GH�X�fY�Z�D�"OL	���R,v��X����"�x�1"O� �m�E8&�x��]���$ZV"O*ل�	y,�x7fF�6��}"O�@�⡗$kY�)��":Gz7I"D��s�	7iR��jC5��M��B;D�4��>F�#ï�d��]�q8D���.:���bm_�/&�9���+D��k�G�;���7L���L?D�����79�@]�4Ϙ 7_��2�"D�B� �Y	���� C���r & D����gƪR��ApB5	�Ѻ�>D�`�R�-�DP�F�[�t��y� �=D�(��z���g �^�R)P�c;D�2��%v�M�A��J<bA��8D���
v7�S�A��p��&6D����m+n��E���W)�P8��7D�X����rB�ÕB�?����4D�L���ڏM��x1I��;	4 �3D�34c�#m�$""��9��YCg0D�H�����.ê@��E��`נ�s�a.D� YV$��Y�(<(׫%�Ψ蒊*D�H�P��m<����S��4eJ-D����&U:4��I��Dm0�d=D���`&j���h�#G��lڱ,;D�h�aN�,.��(4E��s�v] ��9D�@�˷{���IGO��N
\qqL2D���7�A�b�����匦[3,��R�1D��#���R�"4���,���-D�8�o�CE
y�X��#�'D����F��p���]�	ݔ��L$D�P���ո5���kf�/`\J�r�,D����(�9)
�5��[��(f�*D��X��ڻs���D����,�@l$D��KUI�2��1�mSs����#D��Y�@�&h�0Z`�L�k�4���"D����W�Q!J����:xR��r&!D��pD�,�b%#%�ƏN�a�rD D�� ���"=D4�����4̩˔�>D���V�l�d{0)�5s��P�,)D�d�WbT�;��ۦ��!��p��#D�Hڅi��=,t��.�d�Tp��'D�dR�+M5����W�[�dTd2��?D�h �C)���GcO<�: �!E+D�PY�� ��i��!�1��0z�j3D��T�֮&5���K-�´��0D�H:e ���F(�6;�~�{T"D�Ԩv�	�P�H4i�!ڳ�*��>D��r6ȓD=H)�QHR&�8D��&D�4����+L��x��L[
�**D���L0Nؔ ����,"FlȄc'D�xi�섞�����噐e�4|���&D���և��T�2���\��> öh1D�L��P/]�a�S��3uĀ�g0D�h; (�!��;q(Į'f�t[��.D�PbT��Zh�q$���{�Cw�-D�40�eH�m��o[LU�I�D(D��-�Ed�L��*[3B�@&G+D��R��GgZ�Y�p���i��P0G-D��j @M�Hv|�K��#لL�� /D�h���<YN�87.�e�`��V�-D��Q"�N�ݖ�Av�Ɨay "��*D�p[�<m�432�g	(D����	f�|�!�"0$�@��$D��2�ɨ)���'E7/�ޜ��c6D��xH��3Y&X���f���%�6D�� Z|H%�S(]�L(#V�b/&	W"OFa��Dd��C@F�2tް�3"O�͘���w��0�ҽ7�$���|R[����	�?�& UhN�C��[@.T0_�tB�ɒ ��E����5 ֨��(�W�^B�	*E��p]�1�:	��>!X�'H�'��>���9&�x95I)���DY+ojhC�I�3ʼkdO )ظ�D�FH�􄧟(�Oh��Ŕt���j��Ô[����"OK��
�I�m�H<��U�{�<�3��䦨!&	��*R����R�y�ܾ�-�JR3SgnU��˩�y"��d�\���D�k�� bDM�ېx�ḵ�᧐,�J��q��%7�8q��'��P�p�ǎ�6��+�<u�:��˓,W���W��� ����ҠZkl<an?D�(��KB
d��M�5ϟ=�b���K?��O*�b?!�sQ��i�6l�Dpەg;D��衮W1`�ڵyP1
���K�O"�=E����_X�`��g��ZՃsm�5e�!�Ă-G�0Ð�����:&�N'M�!�d:Q� ��L�n�}R��'t���)�S�O�l!Q��QSX�o�[�*
���rD!�6�v��!ԃ�f̄ȓp��#�.!+��5�p�p<H�ȓ*����ĎP�o,^T��ϖQv��oڄ�x2���60���
:ȉq��X��p=�P�$k ����/��Ԩ�G�D��$*�S�OV�ᅮ�(*d�)vA��f� �}��)񩊧]z�-�q�@9]��TlG�db!�$�"ǒ�	W�h��}aCL�1O����P����V)O{o� �dB� E!�d̛]����o�2ka@H���ܚc4!�d��:����RY���"ܪ%HqO���tC�	+Xha���'��c�G�	7�6�&���O<��q$OH&�Bm�tV�c��	eX���ؠ>����t��'o��ƅ)D����WM,�h����`�vHz���<�H��E{J?]@�B�!��$�rІ8spd`w�8OP��%X��8��-
��g�8��	x��(��tA!�߭4P�ЛlгN���ɑ�IF�OW�}i�I�U��Q��*[!�:��ަ	�>�����6H ���ϒ6G��Չ̥!h!���Z������>�,�8�0B"O��K2��1� ��4��	^����)��aAȕ�x\QjDL�T�zE0"O��6m�3%� �J�BZJ���"O��,� �'٨H���`�;O�=�'��'����a�#<t|S�L��RjƐ(�o $�p��&��p`g��$�D���9}��)���4��0���߁����MѠs;���$����$W�93�p2ϝ�r�F\����OC�	�x&��4�D#C�r�Ң8n�f��D,��4I`!#s*�tA�0�5�Aj��'�ўb?q�p���B?�����/'Y�-��h$D�蚡�U�F� U��@�V���/D����#Xx1q�aD)�c�#D��K��җl:�k�kq��Y�+!�O`�?8�t����.B��s�(B�?��ȓ_������aE䜳�(S�����	rI�U�����')�%(�z��J~��g�3�Z�k���|gP�ȓE���"����`�&ƛ�o"���ȓ=����&-oE��ꥭ�ڠ��S�? �k%a� ;�8���� A%�!��"O�R�F6\Ӧ����D�c!���6"O�|�P;�E:V��@���"Oh��@�Z9VLz�B(y�eX�"O�RR�ش,�u) Nф<��%��	a�d(�#B愄�2K�Jkl�"���5�!�.����5�՗>i �9@f���6�)���H' U=7y��U�L,&Bz�:��1D�l ��
�}��#�+.H�!k�	0D�����xN�'�-S��٢�)-D�zJ׸s{��y�l�?־*��)D�Њq�����iR'��6��9�7�1,OpOl�U*�����4��i#�/+X@���^����|����l�l8�g�:)�^a�I-D�H�)
<C��f ېTj<���+D���* %h�'��5(�	�3F*��G?��$�~J��ҽIk.����E�DJeIRN�z����>)D�փL���b�.�Ҥ9��t~RD�M���Z�����)0�t��"Y��B�'H��L�����̬a��:=ۄ��4�ē,��*$�I�U��z�u�H�%8��C������f��>&|��ք�:o�܁���7D�ʑA�=}�T�H��ۊ��e�gj7D�x��4( xM��5:��0��m4D��:ed�A�<L{ㅌ�K���b.2D��a��ʸ~~��)FD�i7
0lO�㞨)�e��@�C���BQ2�)�d�TB��$ZJ�q����Q<N8(�"O��bᗟ��]�C�:�xp"O����I9'�pda�����|B�U���O+�m�6hC"�"�Ã�]n.8���'�P�Kci�=�d�s��%b��|����=\O�����>�Dp���-��}��O��R�-=٠��wmיgԀ��%�g�<�&����� iؐ#(r�+���`X�pFy���ƥ�ndp�˜�y�c[�4n���g�� �  �֝��1���<�}
�nU�Y� ���"B:���Au��w�<a��&B'F�:?��ԭ2�lL����x�O�puQ&=%ՖA�E	2sA��'�x��0��-R�}{�k��j@����O��=E��I XE������6�p9�ԩ�y��_:���	
�\�����E���INX�\���
3�p8���٧P��Fc2T��Bu�Sq��]��k�@�"�"OtT3tbP�QbZ�y��ĶU�⹁w��{�O�B��1�ժg�P��uI�}����/O£=E��gY,F�`�(L�ژX�掷�yB�gϲ�ÐI.G�f,��Ԙ�y��|a��S���5�>Q[f抱�y�cE�SZ����K�2d����EK�)�y�hǝU�HM[�U�he�ȹ,��p<9��ā$#�vd��JK�*�$�*�	��JcўL��ɬSN,���Q B�|����*�@C�I%I�� �@H�-�>��;/�v�Iz��h���x�ۮs���O�fz��W�'qO��0E͋,iw�܀2
��'�HL
O6�@9 ��3��8+���:��N!�D%{J`	�I�Fy2�� �H4	!��1v���uĉ�c�@�KgG�5��'�ў�>E�f��bk���ABA���ԃ1��o���~,8��N*_��P�L5�6L�<�
�70�@�R�˲,�=��JP�*	���WJp,Q'��8E���4a��bp��S�? |���(����m�3h��"O�%!*����H��O ���"O޵;2K�0�zH�F��: �t�U"O�X�JΔ�~ТR	�+Grx��"O���#=����U^aPmy�"O4�0"�@���Q�F
a�>�y�"O��g��&���FK[%U\���"O�t�Bۋ�����ʋ�~Q�h��"O�$���_�?ɸ�r���80s�"O�APV�C7y��p��#O�	|��
�"O^|�&��:19Vy���ud��2�"O��*M�:��lX"l��bh���"ON�X6B�`��P#G`T���"OPAK}�htH�L.%B�5�3"Ob�����b>͈Q��i�R��"O��ƅT�S��p"��M�>��D!u"Oā{���~Wdl���,3� ���"ON���OAH�b0���K7�H��"O~Ԫ��>��=	a��=%4ͺs"On��'�Q�K�H��o�8L���
"O�ٓ�Ͻ�p���%-���w"O�b�_"fBZ,�Y�5KnIт"O�r6f�/h�lK�$Ѽ49���"O��R�BZKZ(83�O�KJr��"O�bg�����t�ӐJ
 Q�"OT�" n]>x��hF��q D"O����36e0���̒$x�Y��"O�M�T-�k�����&�+�lpp"O�x��S7EX<!�N��~��a"O�����ȥi����L�)="\1�Q"O��A���p�AF�)M!n���"O��Q�타C��yHV�Ǩ=v��c"ON4��Jȹ,T�p�1g2;��u�E"O��#�gD1^&���ǁ&u��l�"O0U���3dy*�ȊK� Ԃ�$N&Wt}rrI[>p
�Y(�AY�'�~�BI�(!O(���[���(	�'kn]���@�+�U;�� �'�"}�d�Ѹ��� L�S`\x	�'#n���A�q��H�E��%,�i�'I�5i��5gRҘ�����`6
�'�0%�"D���(�`JV>)��'P�X�M\�h�G)��n��m����"�;zʥ�3��#��J���j�<��o��K�4LP���y���\d�<ф"ހ^b���F&|9JU��>P�ZB�I��Z!�a�!\��t�С#'6B�Ƀ?�L� �kW,���r��X5G�B�ɜvN�=J��ѿT?ԌK��Bae�B�ɛv��p!JQ{M�+�A(~i.B��3fF�xR�}��Dd�>c�<B�_m�lCB��/(�t��W�ط
g2B��4TZ�����[>@6���K�vzB�ɮ{�y�"h-9� yFFKs��C�	6F$���C�ǈ�Co���C�+ZV
�ZVņ/�Fa��LD5dKC�!!����ǎ�X��Вb�?s��B�	�E�`h��ӣo��P-(@�BB䉺S-�(w�-L��D5(�	[�B�	��U��.�/wV2-��ď� ��B�ɦ�����_#QD��pj	o%fC�I�	Tt�2��.v�V��U�̠�bB��]y���e����4�4�M�'�pB��9*M�Y�� � �X	�˖' �8C�I�)�ܩa1f�9et9ig�֔T�B�)� >�#Ê>&\!�G!1���R&"OhrQ?B\��a.̭zh.�"3"O���fr����I�z9�v"OHA&�ؕl,!
&� Ьܢ"O�����ήvZPt;qGؤNǔ��U"OܸB�h@#���ÌGf�>��"O֡�ΞNE#�F�2P@�"O���*%�����H��@�p�"O�j�/��wɜ��6
�!9R�a�"O��c�؝s'Z�g߂m��P9�"O�iH���$s��P���HlK5"O�`TLB�U���*޻Z&P�2�')�ɄS��E�UO�G(���9w��B��"�!�/ֻ]�<=�7HOI�">y��i[z�.t�5bD���l1凄3s�!��*
��Q-�o��(���
q�$(�S�O�� � ���5� M�d�#9͐�s�'֬3E@�X�ꉲdgӱo�d��O����U6Ci�m@���b��B��2Ca~RQ��!QO<�2�bD`?R�V���G$D��#蓣����'b� ���(&���*i��5-!iH7_�Ġ�"O
�˄/C�������:%���S44O0�=E����71|�(�`�� 3�H��C%W�y��H�R1�W/��NlyFcܠ�y���d�<I3Va�	p7h%��`��y� �2b�p��+Y�>%�&Y��yGݑ�JR�$�V�\��O$�y���4�X����D�N3e��>�y"�U?skri�aM�<�z�R�O���y��_�Q��=b�A.f6���C��y"�j�؂���mYp�ӆ,��y�FI'�J�So3w�e�(�y£�U����t�ĺ�b�?�y�.�1��AjG�S&?~�qR��%�y�nկ
V"��w��4)e�����y2"ߠ\���ٔ��� x�@�����y2������Z����ځ[��Z��y�����q������ H%���yZ� S��hbȩ���̍,b��'^(4	UC������ �Nr��':�tJ�#զN,���������'��`KUC;Kl�Qg䔳4PP��'��適n��:1��zJ����'�`���6P�T9#�$��,bz5��'7�űF�!tH���\�J�`9k�'� ��פKl|���CX�i��'!�}��a�!G`x7A�3Hz�y�'M` yC�\�@�C��h!����'�����G�_&8[��;��a	�'b2z��]
���@b
����'W����&�d����^�HX3�'V|�/����Чp'����ɍA�<a���/�nh�f� jiӢB]p�<1���V��(`�� '�زr��K�<�3�"�͢�JM�x,����Z�n�!�E�D`[��M<ʩ��!�!��$pnThe �����"6�%!�!�?1 @�v̜#W:�a��",v!�䝳h[x؁W%�d|���U-�!�$B�rQ�)���R�z�MI�!��OztI 5�z譸"�ȓ��P�D
Z�Y��%!�Ճl\t��>��ݒHٿV�`��� +�T��S�? �,ؐB��u��i@�	u�v��"O�ɱU�XU�ʁ���T}��"OH4�7,�W�X|�"g	7bѾy�E"O�ա�!�%P��#��ʄX��5��"OD�:��כ}�d�iV�2�� �g"O�I��V/b蔩��A�v��"Obu�@bҤ&a4H(U&^�L��H��"O�u�H�'A����Ł/�n$�C"O���b"�G��Xz�cE42�"H�"O�}��<i���0�ǉ|���d"O��kr��?q�Z	���-kj*���"O"t�=Tv�:�ϰy���"O��zb+�XOL�f,�KM�ܺ"O��V(46)"��/ ?�DQ�"O  �u�[�:bh� ��YQ�|H��"O���+�� ��̋
z�0(��ɱ|��pZG��B�OQ�m�������\[�i��'	���44e>Li���Zs�X��'�F	���O��*D�K�\1R�i�'��y!v�԰��4�##�P��4b�'��Ѱ��;�JF�'2�!���R�!h0Р	.M
��P���@܎T1�-��F�P��`�*T
!�,ٷ!KiPE�'8�zs�L5?rDE�R��B��Yً}2Ð�eU��p�k�,0���5	
]�Ӹx�:���Ͼ(�� &'H#�B�Mp�=��5%�̥��7J/�$�D��2"��D{�L\�1Z�p��b,ʧ��D��?���Bc���v���R�r6�r3O��{t�W�n�R=)6-@@�k$+�:Fp��v�U�a�N�8P�ԹD���k��d	7q:u�$Ϝ�h��T�O�m�џ���<r���r`�� =��""�6d��
����C[|���挽i�B`JFY.1�<��'e�]�7�'.p�["D$\ș����{�*)�Ob(mډ�,؛Wn�)~�cR�ύ'Zč8���z���b�8&���@"$N�W�8l�Wgp�@�K�x"ł#�X�CGI�i�0�`�(U57T $��ꀷ?|� ���Éu�RIK3��h�B�� O��]w�ZE[�w`�YTi�Z@����рe��a�	��:��1���:����U	gr~��'��6�$�� �gF�`'ǋyN�5Qc뒻��A��c{l�����$�uGR:0N��j��L5oW@ɂ�6�:�҅a�
/`�Y��"�����iL�OKh0�WDU�Pq�Z�M��4��$F2~FPQU�M#h��t�'�z�!f����	"Ҫۋ]t��Ox�xVБT�R� C�%g6�H��c�
Y�m.;�}v��3��F��*3��� �'�+.Ca�<��_���x����hqU���N��ƥ��z�~
qD���Ša�bZ��[�Nq�7�lZ�W�6FL܂`b�.6$�K��'�Ȅ��(cZt�oI*�N�$A�D�4�r ƅ�z���",�:BKL���)eTT��H,�T�{�D ?I�
� H{�90�JAK���/�E�' A�S��2S<(g~�2�+� Q�)4���5_�AI��:rB��£�3E�Q�U�^'΁s'A$Ox�uǙ�yqX��&�E$ٔ=�gR�ēÊ�4s+�<�&��0���l�?=�^`+��H�nɚם�<����g�HcI:p`��["L�骱HB/|C�B��,(�ٳ�K�U��`��h���"B;Š�!��ڍ��E�&�@����KU��p O�k��
	*�RWK:v�P ��HY)�,��D%D�� 4S.���Bz����O�Q_
LkUbA8m0 ȧ�ʭo��*��5W'��Pk���<zS�hd,Ch��yɣ�"�u�ك "`Jd�J+����ΡZЫ���Y���,�;R�8j�`E�X/>����]gR�sa�G�n���Ar��	"��C=:půO��rl�"�؈
W�Q
�H���d�*�S;�$M�Wgбk��)�S� t�C�	�X����dĹ �]��_4|��=���"\FR�[���'+Z�A�篛���K^����O���c� MX��0��a((�C��q��c�`�	܀�ɃEv@N�7�љ|�*$���Ț>^$ )���u����i³؊����I
k���2��ȝ5���R� ��
���K:on�K�.��#�5
��J�@TKw`N'%PU[�%֖4N�����v�|z���D���Ng�J|�v����(�%���F�R>7�I@�"ۜ�Q���m�(�C�P>Uj�V' ���C�@�
7��r0C=D��Je��,#xXYT�גa� �0��X,V3��BbG�FSr91�����?�A��<�Q/�bl�2䋥y��ѻ�#Pq�<y�������Q�Q!z��L���v��q�-�3������`pׯ9�*Q$P8�㉗1� �)U��n�0����#AtLQ$�n�P� A2cܮ��0�ȼES�}��#,aR-+��]؟� ����N
�x�#���\�,H��$ %	p��;8  ��T��pu�8;%Bv���J`ϋ
���l��DN˺9�Iғ�؛dP��6�ЀO粠��$<����I}��~��0����%F[�@���y"KDh�r�I12�4  §
��~R��vO���A@�>Tay�Œ��H��#�>"��abGB�y��K{�H��B�9U�=�Q"L�ybC�S�xh*3��V*(���,�y�Ҩ �*9�m	�b�5��Ѵ�y�엔<�f���Ȕi)�yt+@��y��	?vً�䎵b!��&�U��yr�ɽi��Ha�ȄU�0�i��y2�]M	��� ]�=0Npɡ��y2l��N9cC�S�-�j5Z�i\�y�O�6�@%�dU4����U��y�Ȭ_H�sf�7d%�0��-�y���5����� �jV�;����y���>>������ВI���y�aL������_#�TC�,��y��B�( y�S4����N���y�&Im�Z�& ��Q���yr�ܗR�4�[�	' �F�+��م�yB#��y��9� O�9~�&����y2�P��r���y(�Hq�
K5�yroO�<�ڍ��`��(�ӷ"���y⁎�(�HR�c!o���#D��yr��� ���I>s�I�u ޥ�y��ÜX!̋���Rr!�Ŧ�
�y��I��`��%
/Ndnu�ČU��yB�(oEv}��	�rh�c/��y��N�)�"���H�~Պ�H@�R�yҊ�`(�q��r}�ap�׏�yB4�> I�hE{0�t���
�yRmأ���A�h;6a�5L��y�*�fϴP��b��;��q�Uc	��yBL��a0�c�c�1��Xc6A�8�y2����S+�/���nD�y2	X�u4<M�3	��,��ĉF���y"�Ѱ(��h�L9"�VAӕGٸ�yr�K>E�X� &)��؁*Ej���y�j�!7�p������|���d���y� YaHp��	M\T��f��y�z�`��@��<�L�����y��W:D_H!��^���b�[��y�b�����ppd����5�y�B����� `������C܇�y���e���câ}
b�҆��y��/�|=����u�H�ń��y�¯�������lm���o?�y��%N����A�/y���p!��y�K�`Q^9����U�A9�CJ��y2(�6Nt�81�AW�����y�Iङk�NV>=7N|��$�y�	�&a�r����:5����f*�yJF�R���I),d��b�Q?�yBJ�G	�is�I�w��x����yR�ˤ ������b%�F����y2	ك
Ƭa`Q�P ��3&���yb��+vNK4 �&dj��.2�̆�"�(�jZw|T`r�N�|�8Ԇȓ1�|i�i����aV�86��n��a`���m��@���߂hr"X�ȓM�(T;1�W0_�B�2��Z�g���ȓ/:J]�����G~J���jݱ�f-��S�? 0�y�ŝ�}�d4�5�ϛ/�h� �"OrDzeJ�cD�c�j-D�t�@�"O�P�C(�� �B�N��y�u"OV�"fK�vŤ y�NV�&aJ�,D�<���
6�IA���x����%M7D�|��J�&I�*�:�&V#v�F�2D��(#$��o�M�<�,���5D���W� ;���a�<n�͠�i7D�T �mؔh6:�G�L;cw��Ifi6D���`Ɠ,^�x���cF)��`��!D�4j��?��X	2��9o�T�ph+D������@�J �l�2>�j���b$D����C#aC(��0胨bb\�x1�/D�P2dݨs�8%
r�^�#�zq#q�,D�`��U o�VX��⊼:�괱�g-D�D��L��3�
��3�D�w#��ۥ�7D�����P�q�V="f(� F����5D��1,��x��A��FgV�#W'1D��4�ނm���g��
M���.D��3Eŕ?R��ᗂG.��p(��*D��j�\*0$�c燼1mΔq�=D�@��
�S�v,j@�5_J0Q�:D��+3��n�����D�0H���q�$D�T����o�"H'� ��P�h%D� *�C_�Nxd� #�� �dlB,#D�@sC>onЫ�O�p�{��*D�D���7~�$x�G�2U�pXȠ�6D��ʧ��c�`z�ƅ�,a��2D�TZF�+צxz�N@�^Q��ED6D�DS� �!��pQu�"��!�ց4D��u��8Xgd���PJjف�2D�0�'�9+Qb	#�	�++<٫�0D�<+�`D;~qZ8d�
�ꌉ�g.D�8��ɂ0�
�ze D���*bA9D��*d��)����aM�%A�8�Ю:D����ؘcy�(�rf�	�Ԙ�-D��z����Q��51�g��]K���'*D� ��+�>f�h�&;5Fl�!)D�����^�ln�c�
��j-}��E D����Űu~�S�@� I��Ӡ<D��c��H7N�p��ͧ1��p#� 4D�P���Z3'�P�@����z�yB4D��!rl�c���a�i^`Px��O9D� �Ν�/��̩���%_ *|�S
0D� B�9�F@c���ސ��0D��R�D�_t�l��]�7�|uJ��%D�(�tmų{�D		W!]
dL,�5!D�<tfJ�M���@��5��8�7!!D�HC� K�:d����&��pf�5D��#�	�3��-��Y�|K�-5D�`Y����vd&�'�:�ơi�>D�@:��8$x�cv�ՙ�~�ٰ:D�L1����H�c���,�j�0f�;D�X�U��y�X��Y�2̀�X�D%D�Ta�#1&�� S��݇z2t�T>D��9�.�0�S�����>D� 8V�Gsr}��6a@�\'(D���eA�8P^F ������D�$D���"E�.-\��/fP(�/D�4�SC]"�X�#E V,�s,9D� 	�	§lgTE�uIQ�
��9(3�9D�\�f�ٯo|@@��
[����2D� ���B����S�-t"4D�����OE~�򄃚X�N�!@G/D��  t
%�%P�����D�=��1�"O2i���Qev�Q�1bA�*��iq"O��kRN/0O��;�aǳu����""O`̂4E3S��ͩ��I�[<٣"OLթ�(�:2�1��gtc"O�	��/4����,hI�#����y�'[�nf�����0	��+�����y�)�.�`����ڪ{Y��( �A��y���M�t��o ΂�#
N��yҩ܅q�� V�\-x$^*7b��y"lK)/G>=���v�<x�6��/�y����8�ʝk�Mj�����y��YlViK �ܶ��he�,�y�E^2T����_�M�̓�\��yr�)b?�)1\"�@�Z� K��y��L9m��C͟�q��5`�`�y��\	�B`[ -�lf�i�5E��y"�24X��c�SZ^t����\�yBG93�RL�U]v�p6�� �y�ˌ(T%���F#WQ6d��O��ybO?=Y�`2!nE
z�Re������y"�8�Y!C��*{��!���y�g�F<y��W� ��ۆ���y�_�U�
}��b��L1lm��T��y�GE���R���I��i%�^��y��6��LJ��xڔ��$�yr.C�D�����ۭLP��ig��
�y� K�X���ƋDD	V��6M��y� T�&Z�hʡ��3m�4��م�y2#Q�4@�e �q1J�����y�iA�g
Ruj�Gt�A�m��yg\�� �sڛc��"dԎ�y�j^ e�B��Sv|Y�e�R��'xɩ��'˴$��Ǘ�ZR5+�6U)f0��'ɲ0!W�֙B��M����%|�4PLދ~�d�9�'�8��A�^8^X��CQ�?���a��$F�Ul�(�:�Ӭk�*(S��7@���B��zB�O)n��	V�hz�s���ʓY6���ؑ��S�O�L���
�xI�8HB��7?��yy�'�(���(�$@C+�7G�P@J>a3K�2L�LX
�;̵��̑�1�ȰR��=>���I�8ڝ��IҐ�V3�ŝ<#ꈣT�^�x�.��|M��:��*Y������cϘD�
�9t�r�#�߸��iTe��]rP���Tc�!򤛌���s��Ũ}��Q�E��H��I������t�)ʧ>Q�	WFV`ks�ݬ\<l���5���ҖF,%�r!���,!�H4'�(���$�F8��	,28��G"�1VL����W��@C���	760HE)��'��E�4b��x�.i��c�W��C��Q,i  ��?	_9����"��Dޅ}�➨�tk�@�Z�����6���T*$D��*0C��@9*sa�A��A+��$D��Rg��
�Nm���,N����q�9D�P�d�ɲ�&�X.)�ܙ18D�����Y��@��i2Z�8�C5D��Ǣ��h��D�O,Xw���+'D��iQm�=�8�5�٫~�h}��$D�l1��
�XM�9���Ҩ;)Ly"��"D�\)��	tX ΅@���ٔ$5D��Q� �<�\u��N�t���?D��#�x �ѐ@"t�Zy���!D�� �M�e��[�!��Qdzy�"�<D�P�cJ�%%��ȧ�09�:��(/D��WaHo��@F�C���ë-D�� 8��VF�������Q81fP��"O���@�W&Dd"�I'��ZV(�ڃ"O�[����q���pǨB��{@"O:b	�G@Z� ���.�X�+"O4i6lG��J4��J���"Ol�p�יC}ܝ[��Ӏ5$̈!�'�V9@'� ;�l0�����$��'o �Iө{K��)�'ʽV���3�'������Vb�V�ʑ:�'̜T��� ���E�4\J�}�'�`�rE��X��-f��� �$�K�'ƺ���,_����2GO��|��'xHu�r�\�����Q#�5iX:Ls	�'{nT(%��*t<�mT(��%N�M�<itc�"6FlP���ۣ>L8�vj�}�<��
�$�Uț[�!��J	~�<�AD�+ l�� +p���g�<Y7&�� 0�5��F���P�b�<�� �+Yg�9@CK K��ѫ�
�_�<����#�}ۓ��Rp"�+���q�<A�ER�q�Q�I	��y�`w�<��&8��#O�M��쀠�h�<T. �����sOX�Yp���Ùd�<Q��"�@���T�)Ѻ�$N�N�<i3��f�D��#E�g�	Q\H�<YC�A����R�œ���(�G�D�<E��t=,\�ӄ&"s���U�[�<ّ�B;!�*���G̎�!W�<���S�1ubPQ�M� P��Y�M�<ᣎ�;� y�kѝi$���CGH�<1�a��8`�ȳì�7�i"��\�<r(1kԦ�Ñ��|�R�It�_s�<�WƂ{����) &���q�n�<���Jeu��J	�*��i��M�<9s�ٺzl��ca_��Dї�w�<��n�pr����!��|U�b$j�<IF���Dm��Z��V�yv��i'��\�<1��-�R�wlķ@����E�_�<9vC��6�bMk�Jԕs&�i2B�[�<I� Ë_�v�JF�T�Āi��QS�<�b9.Xg��K<�}�s��{�<Q#l�pY;4,�]�DԈ��t�<��ǋmU�Y�P �+Vb�ňA�tܓ6�~�P%��;0@P�B-�B�n��F|�ڴ�6鐀���+�pW(٭ xf�0N�0@��%�S��Ԋ �ǴѺ��'�ؼH&4���j�P0�R�]�G�V�kԡ�q���ȓF$��aʂ�"b<�[3�ű<���E(�pa�nJ�&ڬ`�HU��	��#�T7p�̃veA�W8�܆�I\~b�Oܳv#����X�PnY�{�I���O>�=E�dc��A�ְ[�nL оM+�DS�Aa6�Gy�O����H�8L>�$��V�o�(_�o�*�<���<B0��=�j�єf��bx��|�FP�Oq�f!�����P]F�^�'��<3vP��KeI8�	B�O�ƙqj݄�2����Ã~A���ش3@���'*<8��������@�~]�S��%8�~���M5.�d�G`�� ��U�?�OO(b���#_���"��=h��}�� ��O�OX��З���򂘱,>H��f���,?J�<�}┍�3k?��y�a�7&���UfPOy��F��(�`9;K�/��@x���W�|M�D�'���Fy����	�dꢄ̥C!��:p�ԢFYў`%��}"�B�3����CW�R����)�P}B�'�|i�HA��M�GA�Xv�0Q	�'�v<P!׻$�^A��Y�_������ �E�S�L+xM��V��<��l8g"O��Ņ3�M�%Od���9B
Oz6�\'!Bhs oC�t~$<���ۓ���X��Lp4m�Ob��� ���~r$P99�`Ԣ���7AHq��>�yBf��g���r��;FN�
l؈�yb�T</�@�!͜[��5���ʁ�yj�u�p��-��R��u� P��yB�B,]��q��猿N�����)�=�yB�J�S	i�qnzz����A��yb�ǭz��8@[1f���$ ��y���F}�|..̘��:��=J�'����g��([vѓȔ
-�Α �'�~�h��ٛ
�PӲL��'�LqH�'�A��$(NPf�2G�&#��a	�'c��C���0p�����iH	�'<*���@Q�J8���`I�]-�{�'9��bEc��-�F�g'E�Y<�0�'(<�t� sɨ�(���Q�4�c�'f��ǮR��T���ʅJ)�4�	�'h�Ԓ���"~���uG�k�-H	�'�4����*B��U.T�c�L�	�'Q���ʓ~����Q�Z,G�X#	�'���R�,:�l���2�t�		�'�(y�tID�z��S)�,w�.*�'��wi0C�6�"6��_!p�P�'G���
� 6A�B?Oc��#�'�� ��������l�/c�yS�'%��0�DԳ!<�I!��?st� ��'��`���:$`0A���h��-X�'%�ػtH�&�"��� e��H�'Z�=����>b@�@(�"_!��0�'�4t�W��^\n�X�'��Ge���'zT�#"��I"�,l�u��'�m*���1@Nu[aBٚf����'�5"�͎�u^.l�-�_�J�y�'�<��W��Y��Y�P��;"�Fա�'5����"�����"�l�;F6>���'{:g��c�yٓ��<<�P���]�F	��dԌ6mP���H�%	�Ԇȓh<�MY�Ǐ >�\��gGQ�g����ȓ
֞m�P)F1\x�`�Aѭ,]�A��:��G�L0)�E�R�X����ȓ9	١VO�k�����ł"*��b�ڝ�K�dX@���*�88��DH��0�@C�JB���02&2نʓ	S�-�ˎ5 )[�.InwvC�I�=�>�����g��+�gGd��C䉍)u"xj�EX,n�쩡��F ��C�	�N"Δ�E�:���`@}�bB�I�;4�M��)%n`R`��ʑ7/J8B��:�.dR�Mq���A���?g,B�	�V�&m9�N^*�d��G�N�X�B��
:>�*@j�b�J,��B��B��C��H�` ��.�h	��H��@�C䉰
��	Y�a�5���� ��BhC��-0�H� 4�X+��%�* �J��B䉚r��@G�:�ɥC�� ��B��u��i�-�78�D���Z*;iB�ɥk\�`3�	NH�m
�˜55�B�l$�|{rhD �d���/�S">B�	+A�� G� �`K�82��B�	�w���2�O�Ib��x��R�vB��l���1�mLuߌ��pDXB�I��갬�%<�PE�!���p�&B�)� :<Jv�#�� ��A4���cd"O�iAAC�M�p���ei�٢"OT��N���� � נұ"O�mr���>3�%+��H�2��"OP�*�
�<(xْ!Ѡ��Ѓ�"OLDe˱0�b@�v��E���""O>E!��G}P8�V��x�bըR"O\�IѢ�>�ri�b����T��"OHB�!P Uq.d�4�Y����"O�eS�@�?e���dA��Yۓ"Ob��i�*�$e3�Ă:��ͺ�"O0��D%�$I�aB�}��Yk "O*(��LVs�>Y��$s��k�"O����a��3�~�����o��� E"O��R�O\<�xq�$���>D�"O�xHf�Mm_����L�<~�y��"O�+1����0y��^�X�!�"Or���ڤ3�kW,E�Y��1 f"O�D�)ʣna�aƪЄcK0�rS"O��"i�l��q#��V2 AP��"O:�s�ρ4q2p1:�,R
u4�)�"O���M(1�m���_N`,3s"O`��L�p�%�ڂ=�1�"OBb"K�>C
PcC�ݕf1��"O�
ba7:䨛�� !"Ec�"O�8�"�S�pB`��〨b��p"O�h�t�G_nP� S2xF��[P"O��p7���z�2�� �K6+-|,�"Ox��p�����p�&���yT"Ob�c��)���s6.�o�F��"O�lIW�I'�rջ����4��)��"Or �3�w���WLB9/Ɔ�S"O���%ڢ?�j���l��F�!"O�]�KC�	�PyK�F(,, ``"O��jBe��
����W+�$#�P�"O���3�F�t	˂5����Q"O������l�L��G؞@Ů���"O�l�á�Pז$!���^�>8�"O. ����9>�zl*�P"6>����"O8ѳ`��b�(0�]�n6V���"O�����+\��:$�u"�"O�,����fhf�#���a�=Á"O��E�';�X+V�Ɨ?M4�`2"O>Р�
�l܂�jN�1Bz`(*O�@+�B�*<ΰ�D�]*<p��'��H�tHRg<�%��M?�t͑�'��,RcՒ|D�q���K�my����'�Tx�c�^ȡb��Ҟ2���
�'�1 ���1�B���"v �	�'�ܑ�1���T�(�/aVv�I�'8���Q!S0g�0����<RzЌ��'B���eU(!4�����_��e�'1>h�Ţ�?7A
i/%x�m�5�q�<�g�_�/����:0��@B�Lk�<��/���j��Ă �[X��f�\�<�p/T�,ٳg�|���(Ph�A�<��kT���V�̺a� ��H~�<qP�J4f��`q�͚#�<��j�}�<��`��-����L�
w�S�<�A�M"&�J���Z�`xZ��d�Q�<��%ځ$����"h�R@���J�<���m|p�e"S�F`i�@E�<�6�;W��kV��K|���[�<9�L�`��IS!����a1�L�<� 	���?���·
ՇMU�k"O�a �J@2T�LP
��s�ĩ;Q"O��� �I\@ؒd�A��D��"O�ڥA�y��iHB�4%_^̨�"Ox�9�%�DOR����5W�h�"OƉ��&�p�R�a@�] NF4�q"O"tL/?~�u*d��L�b���"Oʘ��/�,~���wC�<\��K�"Om����V����A �v`�R�"O��th �7�������m��C�"O�i��X�g�( 7M��h�VX�7"O�X�U�'H�H���Z'i���"OLu�%���C���f�"^\�}�r��D�O۰��1�X�"U���e�qN���'״l�#�щpV4)��8h�@��'������H��X�-�Q���
�'����s��Bh��A)�5FV0��
�'�" 	o�_�Ƹ����*��!(
�'3�pbBC�&:�Lmq��x]"=(
�'�ڈ#�C۰&���+\�jDI�	�'I�u�RL_=
�,1�Q�=b%����'P��@�nO�Tis"�X�Z~�"�'0���fX�zʪA�Y���C�'®1���c&�)y��Ʊy��M��'�
�	�mW8丩�0�Az�^��'�͙�X<I��$���	�dl�ٙ�'��%��B�N�ʩ1e�F�&l��'��L��A9�P�E"Ģ(]έ��'�0�0�� mкH����%��'d���Y��,�sDE��X�*�'&ġ��!1[#��
�	[�e��'�*�ꢫΉ�f�2��=.-���'Lv���I +Z:^eҔ%A.<���'���9d��(�!O��	��'����#�ׄhτ@C�N�f�`	�'@T1��[!j�9�q�	n�81�'X��Ō�-e|�Ja'��z#�'���U�z;*�����%¦z�'e�9`�$<j���	�Zzc�'�F0�C�|�	BGF�cFH�	�'���y$�Sv�|҄����m�	�'��1�I�
;���d�=	��<��'�f����"��1�T��(�@C	�' �z!F� 	��%G�����'��lJ垱1@h�A.	�d�+�'�n�7fS?%�8ai2�C{�� ��'��5�U�_�����cɩw�n�*�')!��K�u�ڄ"q�U%x��mi�'֞�AЁ�?l���ַ��|��'��9� �#n`6�Z[��1M� �y���o�
���/��F���5C1�y�γp��%
��L�,t�&>�y2B�k��h���h`�q���yBm�8 ��9rw	k�X����J=�yRA�1&�1�%��\���K�n��y¥O���Vղ?jЊG�C�y�ꃕuL���=;���i���y2�Z����1��J�3���{�,^��yrF��^����lDR�$Y�y2�5<=�bTKA�b0��Μ��y�	�:r��EbPꗅ} HȠ���yB"�/�1�ίB�Q���:�y�lJ�JUrW	\q�V4z!D��yb�S��QE�h��̛����y
� 2��HQ�R@�%�7,@mp���"OB������Y�jX�EO|Tb"O>��q�}
H�G"��u6"O���$��L�rEP�
5L'"O��A�`%N�&��d�6�|�2"OZ�1u�S:z@� F<O#(B"O0�s�Ѝj|H) �4~xmJ�"O��µ���~\���A ޟ
���[����D���b��F��˩k���Ic�]�f�R�"�AD=w�qOd��^�T+��*&�K�i��j�eR�7O4q��i���X �" 5�d%ܧ����@R�'N0� ��9" ̑�����,��Gى6bP�@	D4��ؗm��W�̸�p�[;����=!��EǟH�ߴ��Oy�v��z9N�z���S��x��(Jnw��D!�I}�Ͽ��]=0uRp����6H��r�n8��r۴xu���i >�"���+<S����E�l���'���dl�B���O��'\$r���?�ߴ7�٨ �
H�Y��&ؠx�ڗ=7�<�����I#�g
��a�C�F?I��?)������g�$t�P4�s��&
P�o��	�2,��(Bႁc�L=0��R�1�zir�,#� �s����\�@)<�{eK� 
6vH��${�v�K��'Gj7�Z\yJ~jȟ�v�ߘB`�)�1�J&	�$�'�ў���*e�I<0 �և]�z���	��M�Q�i��],t��l
��e�Ę5��(_�Ă+O�DX����݆�	9F�r�J�+|�DBdȆ	Y?RHBg�$���{��+r��U���qnV��'� �0욇&=����ޥ&	E�?���A��=P�r��bS0S���6�07��A�	�l��i eR��|�tG� ~���)��A����M�qM;}��'z�V��0��
�Z:�	:�F�-�V1y&C&�����y����=�lY#��1����"�Z��Mc5�iP�'��$�O�I�M��*�(��뵂�t;l��!�Fo>�������9�&S����蟸:��B�iO��3��H�|L׬R�C���k<ű��14���2��ޭ`ԣ<-@=��@__�tuC���p�4Q"�dJt���ק��hTJ���M�ۦ�o,����7�F�r=���XӾL�SNL$G��+��3���Ot�$*�0�	�44��Ѭ�3_�đ�vn������9ғ0�؍�T�]-ԶJP%�g�֥��@�Vk��ʓj��i�R�'����)%��R�U�X �0�ӭG�n�9��F���?	��?a�+�mJ�(�ĀX�PR������]�̽Y6�΃ 
�1�uJ)n"��H�
D�B� �Ey2fD��
N4ZG�a�h1Qw���VpC!T]{eK�E?P��A�*���xѧب��$�"�B�eӐ�'>�nڍ2*][w�ќ8�L�@$ʆ�j�Z�h�������"��#< �`w̎�P<^�3ƥ֊�ē��O��o���M�ش~�0����wx�Zp���v����
�R���i���'���l�I̟�oZ�oˬ�3��X�8�ʨ����?u��p��W�PZfu�p�ȹh�pZ���g�p��5�<��i����X+5���1�ɒc�c��� 9��6mH�[��hq�%HO>Y�''�d��M"J�]�EC(���BP�d>�8��^�}6����_̦2�L�O��o
�����?7M	(5��|"�K&��P�3��v�铍hO�0<#���u�D�U�����h�����OʀlZ��M#J>�'�uGCI�`�V�; �F�[JuȖ2:4��O.��dٌ� 8  ��   +  �  �  7   �+  �6  �A  �K  �U  4`  k  �u  o~  �  <�  ��  5�  ��  ��  C�  ��  ȿ  
�  M�  ��  ��  �  X�  ��  ��  �  ��  �  d ^ �" 	) �/ �6 �< :C �I &J  Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�� |d��"O
`�(�;���8���-0��1%"Oj4��ND^[��"3/9�0|H�"OB���H��*�ʞRy=a"O�味V�!X��!&F�:J�$���"O,��a
���C�Ą�M�"O,$3%o�-���p���+Ն�:1"O��ݢ1����`���y14]2��i�<�6��{_���c�H�`�fX�$Kn�<��A̼VI�xR[�)�Ć�pඤ�ȓA5��('nߡ4�� �)˩%� ���,��r�؊b#`T�eT09���ȓ!�b��g��}�8�F��-? �ȓ
K|m�ș�VṔ���2�%�ȓ"R�X�j�4JN�1�˘X�i����̹	_�jZ��1!g��zܶ��ȓgil,*�J�
j�Ne��i�J%b���f	�(U��:���G��$Y^م�~r�� S�%T"���k\�jx�ȓ|4�1�îJb��@ӵ�ݩn�V��/[`�"�v4�R�!ʎ<��M�ȓ`:��z�ؚh�J�Z��$HY:	��H��p�m�C1��!��B:��0��EnjZA V;9����J[
2���	��4'J�EA�IVW&��~�(aZ��ӹ�>� o�Y�|�ȓ�f�A�
Ο7�H��M�$�����mޠP����/���ANXo*�ȓTv�����{ ��-7�*h��I��sB�8�8���3����ȓNe*M�悡;������X�o��!�ȓ'lj�#F�m�+R&;�|��2)n�C��0S4���T:
b���:�0!��e֊��)��ͷV��,�ȓ0�&�8#���� ع�L�����;�P�AFd���,w�6d��	M�$F�K��#&���lF�� �R�!��	����6Lm.�0��-'��'La|���2z[.��W�_i>bX�����0<�T�x�S��i�,[�^>�$���K�V�飣H�NQ�"~ΓED��H[bxpp��J{] |�0�$D�xK�!J��J5;�*��|��e.o�8��'n\�*�m��M�r��5�Ǝ�-B���'b�h�f�A#N���-���Q�K�<iGF<��t��M�*c:)cɜ���x�FĄ�2}�V�-��Y0*X��0=��B&��
#\]�e	]}��Q�bB�yb�]x�;���|��6m�%�y҆T+&�8�E	�sל:�Ԁ�OD��WS���d� ��!Zq��
�!�8U2~D��ĤU�.�aŢ��,�!��%"Y���Ï�L�d�ՠM�;�!�$��]TR�qJJ%K)[3	ۨ>�Q�0D�dI+xSl2�
�$��R%��ybn��X�ʘ���/t��>�~r�)�':��� �=y����(ʐ JB��ȓ���8G����D@��3{��O66m%�ŞBK�y�t�N[c��s(��n�()���Y}�a�L��穈1d�z��U����yM����HB�M�`�]
�����0?�+Ob �4��	���P���5i��ð"Ol ��.Y%KjUa�n�"}>�˶"O� �t9��ݽ���xT�W
�V��"O:(*N�VَXҤ�:k�������D{��)1<ŖY�iE:�"b���4+�!�DО5�D��P=g ���!6�ɤS�a}2� n�����*���!�!�yRF6�li Bؙ
��r��)�Oĝ��I�
i^a@��>�:H �ِF)�B�":�p;	�5��e���9bP�B�	�gJ`�ђiC���+���8B��^��p�	�u��̶o�@C�5[��ܹQ�0m�HC
�:��C�	*`l*�"�i�U��n�4:�C�	���H�Z ??���(��$�z�<Y��7O���KM��Y���5�1sUOr�D]�E� � ß<~�.�ñɁ�$!�d��q��E:c��*'��؂B	�(ax�Ɍ]9�ţ6�T�%�$�cs&��|W�B�ɺ`��<��_S�;"d�"A5�� �=!��ta�; .�aZ��W�C=��Z�����x�@ԧT(��C/�$U�Ux֢	�"�0xK���Գm}џК�N�^|D�q����4�� ,8\O�U�=�����U���_�<�H�a䅯/�!�dS@�zE�4��40��0 �9	��I��V�Ih�S�' ;8�5�J5bQ�m	a�ֱ!|RE���})Ճ]�8���	n�x=�%�ҧ�y��+$�!ugB�2M��7�hOH6-5�'?u\1�=6����#F���ȓV*ͩG�ـT��ꔂ������#����SF�.$!n�IE獚GY:هȓ>nPAz�^�p0�5iËm
X�ȓ$�<�9�%�^�&��1ۀm���zң#� [
�������i� Їȓ#0ܑ�JÞ8�Rm��%��]f�ȓ)�� �AM�2rh���B�?�h�ȓ$t�B�=��j�&ۃ}�����$�(�K�$*�U�Bӿ?����,����G�I�ع���S�]^�ȓ�4��d-��>/V����5?��IC<y�*Cu��x£��WxӤ�}�<�*\�8n|ʴ�Ε<�`�j�u�<Yֆ��4gZ�W�R��.�8�M��'��	G}b�3�"���c�����db�����$�>�1H1>�RU�Z�7z�4�G���~2�'s6�1�\<x��8�O��{ڴ�0#�S��?����#g��Ps����;�(U�F{�<�#O1��%��-�'�����ϛw�	c���O%��$K�3=����	x�&IZ�']��4⏕9�t!S�gZ8��S޴�hO?7͍�d�|��r^�Im��š� 0�!�����A�MX^�(9e@R�R�!�Z$=���V�	P#���O�6,�{�>��4�,�RM�t�@�a�%ǓWHH�ȓNlq�T�_	�0u�s�Z�Nќ��=!R�|��4�'(�dx0�F�Vv���T�W8���Ia�'�\��[*v~x�s���;5�f�)��<��� P5� ʱe� B[`+s�Kh�<��IF"���
! %��!���<q��5y"X���ޮZ�D\�� ��N�.ąȓj�ppk����n�ܭ�F�)G�����_��IO����&M��h��:OCQ�4.<D��1ä��@��I�);t���[�@<���	�2� �!�39�p�'mM�d��C��A5���!ý+������@?@��7�6�S��MC���1J�� S/UG`��Ka��r�<� dЇ��97���c⁕XV��bc;O�7�X���hOD�
'�\�a��0@�+̫J��g"O�#����e13��n;�X�>�	�`����]�F�L=��bׇ&8@���?yP�9z���p���������Z�<9��� ,�@���b�C����L�Y�<y�-4?�v�S�IC�|�d�m�Y�<��EP��	kF"��]g~k��Goy�)ʧ"��Ƌ�]�T����8r��'�:��p�θG�<U	w,�a��d��'AT;!��fZP��Ma��d���0�'l�h�3��.Y��"A�UH���Yp��+���?5�da6@�|Ҵ̅�!�ع %cʦbτ���
|�I�ȓ?���z��e80A��ML�
�&�l��I�Hi��zm��`!#A=n�DC�䦽�W"�	���B�H�}B���+�<��j5�O&1���E[$���?6���k��'Q���(r��a�:)H#��bPi��R��bL����g~­WQ\�"u�B�rz�J/Ċ����HO�J�M Wt}�w�@02��9㗙>�`�' ��'Q?;���婝�:�p`��~Q��'`3n��x���֨�2D���Q��:6�T
�#V�Ψ�#`3�����SA��6|�	��*�28����"O��Q���Q7j�F ��d͘8�"Or(R��wIJC�+��sU"O�$���5[`:��pM�$!��X�P"O^,jD�ŶC! M�#mN&L�Lq��O�����VO>�氘�8n!��9w��eIV��^˨Y;󌋚|�ax�I V�hi�wIN$>�B�
5}�&B�I�O���ӅE�0� ��̟;{c��hO>���ʖv[�Q9�fK�A�����<D�h; �#>P,�A6�	�9�H�v�9D��3G%/!ڝi�� >�>%J��!D��K�=n�ʱ ��C�q� �3v%D�T�4�W�p�8�HA�	`�A�.D����X L�J��80(��&�y�H�\��=�Ҫ�>i��\�R�2�y����6��(i�H��Rv�ɔ�:�y�I��,x4�� K�x.��k��(�yr�ܧx^�칔l�/s�x�����2�yB���g
୒�#� 6娸8��Z$�yB�	�T98h��B�2/a2����^��y���D�z98���x�P ����1�y�B� s@���ĳ|nj	�Ui���y�Bҹ$�����Ȇ�a�*�u�A��y�G֬ i i����.��t�Ǫ��y�L��07��*'E�0�>�&J���y�O�w�t4�c�Q�44�Y��M�y�hS�N݌ �k�C��X�*��y��X�]�| i#gP)4v�YV��(�y���(<�`��B,X(1���X1�yR��*�0de��/�} �&)�ybf�<O�j�S%�߶|�$���)C��yA��c�)z���J���S��y"'C�� �c�N�0��xZ�,�#�y��.Wf�(RW��z�Rm�Eۂ�y)�9(ق��R'
5>�U��k]�y�%�*d��(����&g��b���yRCM0��-����39b�"�6�yB�I�W�Bl�j��]�d�Җ�/D�����i�|���ݥ]PtA�N(D�� �hkc�ޡ%B5 ���#4��q"Oڅ��,]��q*hпe�И�"O�p��s7B@	6���&�J�cg"O�PF���j�jEږ�Ak��T�"O��[�� B�x��C��d��y@��'�r�'K��'f2�'	2�'�B�'����6��P-��eF�(�
��'2�'��'�R�'?��'���'X��C-�'o&y�s�P�����'�"�'K��'w��'?b�'���'�"aQ�"ڀpx�cT� ��'"�'a��'��'Zr�'.��'}P	�FC�K.�y�d�(|�.�;��'F�'h��'	"�'��'��'_���%��?}�x�f�ۇ"��y�S�'zR�'���'$��'{��'�b�',,�����63���7	�q�(���'�r�'���'���'G��'���'�0�`���8O�9��	4�l �r�'�'��'F"�']��'���'Nvad�?5���)��0v�y`%�'���'�2�'���'��'|��'�|M�RU<[Nz ҋ?@�~E�'Z2�'���'���'X��'���'T�)�B��~�tJA��<|�@�hw�'�2�'���' ��'H"�'���'��䫖� lE�(�͞�x��:�'���'�2�'�2�'S��'���'��H�AGYt��sN�n8���'eB�'���'��'��edӴ���ON9J��-�V8!鉐Q�JE��cy��'C�)�3?��ij��C��Kx��A�`��C����%����Ц	��V�i>�	����AּF-:�qF�X&I�1�v�
�M3��/�|H��R~үQ?M.�I����i��*m袆^�tu����I�1Ov�ĳ<i���*k ����t�`���q::�ؐ�i0z�؈yr���Ԧ�ݤ��Y"BX�L��԰�c�9�LB��M��'T�)��ͦruh�QD<O���2�\�"��th`��>7���>O�U���ņ�f��,��|b��0�̨ڣƏ�Ҥ�!ׂ>#3*����<���Φ���,�	�2`>4�P��|T���t`
�_�Hu�?qb]�\�	������D��<�L]KTj�,.Ly���5EU�	6�R�ꔂF�h�<c>���"L�j�<��	�i�����΄ue��;��E��8%�'�	ß"~Γ/K���BK� ^N�[�h[H0�5�;�����$�Ȧ��?�'\N����	`�<�g��� j|\��?	۴�?�F�
*_N��'��U
@��Px�c�>`���p c�+�Q4��4#K�<���?_J8�kRO�9��%�&P�(���&��^����>7s��b�i�x���k `���|�f��
�>0j$	�<n~�xS��"f���Jpo�L�t�J$҆!�؈"׌Z��R��L/%"���aQ�bJ�y���_���2�22�p�!�iaT�Z�ʏ(5Й����y&A9W��C��8��b�>Hv���S�Wp�}�wohQ�"' -���E�ڂs�� Vd�$d.:a� �X�CX�ݘ�mti�����V�;R��z���� ��DE �`�(J��d;2���M���?9���z����h�S��x����N���BNk�T�@n�����>Q�,ҁ�9�Tn��&_�8�զ�!'����M����?����R�xB�'��s�jآhx�aX(�4�9`bt��5�w$-�i>c�����a-p��fA�o�	�u,��=`r	sߴ�?����?% �-��|��~�G��xF��E9>�>IhUo^��jc�X���(��'�?���?yY _��ݪ�o88�GJ)b5���'�����-���O���9���*4��s|@�o*,"�h�uR�|��J+��ȟ��I͟d�'F  �Df�T�j2
�=-cH����M�Pb�<�	c�Xy�oY'+	S��V��U�`�ҮR$ʀҊy�'B�'�B�'J�[e�'�A'��2(f��.@]�@�i����?YH>I���?����-�8o��Qܮ}B�䅸~6Q��*'(<듶?i��?I)O�03�f⓷k]�Ё�g�O�3���$F���4�?1I>�+O����D�=o�<PIr �.$R�e"b�Z&?q�6�' ��'ER��|��Sy��O�\��@Y
sg.�?�ۃE ���O�����았��T?%QG sC e�E̝��$��|��ʓQ��P�i���'�?9�'A��ɀI���#���� ��R�9��7��<qT�Ob���OTV�������J�N ⓩ���M�V-��?I���?����r/O�'�И�EU�T��5QU�\^��d�5�i��$z`E�٘���ē(�I$ �5x��$bE*T;F��m��	ן���!�M���?���?��Ӻ{�o�'Z�8�Ӏ@���y[)I֦�%���E�z��?9�����o��P�J\f��휴�Ms�?~xɶ�i>B�'���'�v��~�AA`�t����%Rm4���"����
Kw��O���O$���O�ʧ�ܝ�i�[��,��(λw;�dC�R�D��f�'�b�'��i�~�(O�$�V�8A�ř�Hk|�DQ��U��<O�˓�?y���?Y���?�V�O�V�V�I,9�Dq��N� a�Cr�MM�\7��O���O����Ov˓�?i���|�%��c6�c� a5r�a�ُ6��f�'u��'�¦�~�@e�6���'d�̆B
:i���/7+�� !�"om7m�O��D�O���?	4��|RO�APjM=@�: r�,Mf��H+R%o�����O��$�O`��a�	ڦ}�	�d�	�?�Zs/��W��h`Љ�2�EӱgT��M������O���4���D�<��� �AK6��^ ����F��.-Z���i���':r���eӤ��Oh�����i�Ol�˃� V���ra�AT&T���YY}��'*���'�ɧ���~jf����m�q	���0۶bNۦ��v�	�M����?��������?	��?�ǈ=n ��!�O��:H2�"v��}6����	E"�'��i>%?	�	? Fx%��A�6�L��K�,�T��ٴ�?����?�� )$0���''��'6���u��
>{�`A�=P���R)P���<a�E�{~�O�2�'�D�
E�����9]6m��i�p�6��O�-pק�u����	��¬���CO�5!R�_�]�d��� ��2 <�O@t�Γ�?	��?��?A(�&�*�/	a��Ys�(��LS�}N�mZ����ߟ��ɭ��ɸ<��&���x�iO�V����BD�:���Ҡ�<Q-O|�D�O�d�O�d��~9l��O�FY��D�'I��a����Fs����4�?����?����?�.O��d��/Y�i�n���� \����BG"<�����4�?����?���?y�9D����i���''�5z0�O.�tmC��^�	�m+��{����O6�ľ<�1�T�'��I�,_h����8֑@6kY�U��7��O��$�Od�Z�iWn�l�������a�t��KL;e�HUg%��j��T��4�?�(O��D�'%;��O���|n�x�(@�G�	<^�)Ӷ�SH6�O��dG&Z�t�n�џ���ݟ���?��
��p���A6&ȱը��U��>�~"�$J��?)(O�)=��O�BIr���Z��SF��?�M��'�+m�6�'�r�'.���OB��'��Ř.cb�u�� ��|�Q�Z���ܴ���3���?�/O��,���Op��e�D[�4ٻ��ֺnw�p��ͦ�������d�x�ٴ�?!���?y��?�;}�r�H$��u��HC��´`lZ̟ ����>X�5"s��Z��?��"�� ��p��iXr���Ҟd����'(%Рbk�B���O �d�Otl�O��$	�Y[����O.wQ����ߟ ��##�F��?Q���?�������;h(�� eZ$$J���`	I�u��tC`�]�I�	ϟ��ß�K�����?���)YP���W��)44"��ݠU� �ϓ�?!���?�����Op���h��͂��~�8� ���!�ᑱ���M3��?1��?�������O(Y�63�kLV.o� 컧hPU�ܼ��'o����'2��w�'@��'��K�>|B�7M�O���Z8xO6�*�$f�}[R��9��En�ޟ �I��L�'{KY���d�>r$��vΐYdO��%�ߖ	Z7��O��$�Or��M�I�dl�ٟ��I̟@�S.Ԯ}Â��-'�ư���Ț|I����4�?A*O�����`���)�4��ơʶ/��!3�b������d���M����?����y��&�'�"�'M���OsB�K�CC��ԣ�q��*v��)����?�Ů�*�?�M>�'�������"��)���( .P>��7�@V�nZ韨�	����?��	ǟ�I :���85�̋td���"��Oؘ�ߴDX��p���?	��B	���'�䧡�p�I1��%� O�i�xd�D*\{K��'��'��}�� iӀ�$�O����O<������,�,2���ͩ1&��Ჲi2b�'\�@c .�yʟ2�)�O��D�0�LG�˲?$���J\�r��mZӟ$"�OE�M��?9��?ia^?e����4b���VC��� ��%�n��'z��;�y"�'HB�'�b�'7�)i3�������EɁ�vd��PU��1�\7��O����O��d�k��Y���c4!�EDX��*���!9�d1���1?9��?1��?�+O$��Ƌ��|�"���S&�l��ɲ#��A@�'C}r�'���|bT�09��>��+ˤ`�D��m֬x��t��
{}R�'���'�剭a�m�M|�2IB x� ��eI�|f�q�&��-��'��'Z前=��b����)
&l��+��9W�t� |�L�D�Oʓ^�Ш���$�'���+ѳ�&m�tc�1\"�y� '� O��a��!Ex����!�R�y�
ݠr�=̘���i7�I�2��z�4=��S����S����R�XT��1t�X�읈&C�VZ�����7�S�,3&�lB����BCbT #�ܐ�4, �	±i��'3BS>��?�傅�;L��`L@�O8�WÐ�m�����=�O>���ԁ�v��h�D
;7IV���"AqΛ��'���''Z�٠�9���ON�D��@0��A�Z����ۻR��!��6�	)��b�<������I3`_��[7�ڥuO�3�m��)a�4�?�n�űO��%���,ID&�,�2��U����X�iw!�����I��'�x	��� JpU`���c�N�h6���ZO��d�O��O�˓Of����M|�\��Q���d�����c̓�?���?�/O�<�KS�|"�	�	p,@�A�$H��$��DHO}�'�R�|P�б!K�>Y�b��v���!w&V�z9�we�E}��'���'z�I�:��d�H|2&�\�����I,��5z�L��!���'\�'B�ɲJfVb��ĢF �q��)�Xus#KcӖ�D�O�˓ �9K4����'�D4pJV���c݃H��A#�nS�O�� �^DGx���i&G;rD�
�H]�*'0����i��G�%"ٴ'�����S����Ē4;J��5��y��D��!� 	��V���� �S�@��!�C$0=�)�䢏$�8�o�70�p�ܴ�?����?��'
��'�B�͊s�tct��:�!W$��6�Q���"|:�*b� �\�u�R�*��4��{�(<�i�B�'�"n�`��O2�D�O���"�"3�,5Z,p2�,�.b`�b��cT�;�	ߟ���͟H�`/ܮt�6⅃�/�y�Ԣ���M��H���Ӑx��'b�|Zc� ��gJ�P���HD�Dh�O�D����O^�d�O��NT��� CҸx���B�Ǜm��ٓ5+�m1�Od�d?�D�<�s'��"m u���M������V:<�<	��?������@(���'U�b�AN;+��D(Ɂ1sr�'�4��K��by��H��$�4A,$H��4#,j5�	�|�	꟬�'u����J"�)C�7��+��q��⋁)~�z8l��%��'�^ !�}H�7)U
@��<�vt�t#_$�M���?�/O�
@�FT��0��?)/F��U8(�����OM�J�ݒK<�)O��8P�~�`�
P��+1�X�S �R�R𦩗'&���u�~�O���OdZ�}=�� �)K��E[E�ǦN��MmZpyB�R��O���و�)�%P$�x�@lH�>{�TKb�i��`Ȅ�dӼ���O���|�<y����@��,� @3P���0o��%���?�g��?!�-N�/<�i`
S�6��H��+��1_�V�'��'��ೊ+��O�d�OH��c��#;B�k!G�C�5�to�i�s��d�<a��?)���y+u��0��2�I!\����i��A\7[�$OH���O��$�<�1sj����	�*8Yƍ7S����'p�)��y��'X2�'o�I2C~�x��#�	$E�Ɓyᘭ��������?Y��䓳�ۈ`C����%��l�2���eD�=J����ON���O�˓o��C0�n���B� ;���O�:b���U]������8$�ԕ'g���O���a��'0��"n˚+F�y�\���E�Iğ�'��)#+<�	�?�z�!Q�A6$i�C�5d��nZϟ�$�L�'� q*�}riM�?,�7�V�y��%�T�Æ�MK��?A)O�a�P&E�Sß��S����C@���V���@Ğ�<�I<�/O>�t�~�E�Af���W�E.�j����MϦ9�'�l��Fu�R��O[��O�R�L�f��,����r��&2��l�lyb�Ȱ�O��.Qr��{�VQ�D��D�h�P��i��d�¤}�d�$�O������>y�$�y�`�Cաѕ\�a���/A��f��O>��I�KgR8k��L�M{z��5cSj6 u�ܴ�?����?i�L��J��O��������j��1�@lX�U4$5�!:"�+�I�dcb���I����I�!�D𒐠^[�L��
F�@�Cݴ�?�%�۔m��Ox�d?����(x������ă��q����bP��P�7��8��⟈�'����	�l;L�)���5��I��Uvb���I]�	hyr�&�r��v��?FT�#6ġ,��9��y"�'���'���!��OOХ�g�mn�0`�����$�O<Q�����DX�pp���4��w"�,/�}a�bƃ(��듂?���?9-O�<�q�z�06H��Qe�
Tv��3wKH�+�|��4�?YH>�(Op�U��L:��l�B-��W.��s.ګ\���'q�Z�|3n��ħ�?��'*ʔ!�v�ͮ_ � w�W5"�@)`��x2^��a`�9�S��"F�
8��@�̤D�6�%�
1�M�/O�]�P������������'$�Y���?�(zЈ�W��T+޴���.4��b?Y"���HpEGB��ӖAz��w�z������Q���� �I�?Y�M<Q��<�N����]�! p�BWR�aҔ�S�i������Sڟ�Q`�ٸr�$�9��O�c
@���ű�Mk���?��j㰄x��x�'T��O^�v��>�ȸ��i��G� 0����=Um1O��$�O~�d�%���'EYx��P�n9<K0n���8�Ag۩���?q�������˕�l�G��	�N�E��]}r.���'b�'�bZ�`Hb@�"F�� �B�2�T��kK2� 0J<9���?AI>1-O����c��zȢW)T��B'�sx1O����OD��<��ן4X��ZjRצ�)��YAd�C�I�����Ο�'�2�'�`���p3�.�7Wi䅹��+k[�XcQ���I����Zy�h��7?�����ç��b�Rt�*c�aaC�Ǧ1�Iȟ��'k��'�B�ʟ��+a�X<�h�E�-���>q�,6��OP���<	Dc�/�OR�O�X�H�
ӼJ�d咆#Y�m�R5J�G`�T˓�?Y�oUJ����4����.EF�C���c-B�	���M�-ON�/�B,n������O��)b~�A[�t�Ę;b�Ɓ.x�[���MC���?i�+P�����L<�'F?!`0{�	b'*-�0�������E��M���?����j��x�'�`\[�A�U*:�r��<2lUC`�i�� j%�i>c���I��}Fk\���ݕJ��� �oΦ5�	�����8\���؉}2�'(�$(/�2���X�n)X�g7�O���r��O��$�O���3�Զx��U�>pd�����Ǧ��	�#���ۏ}��'�ɧ56��2ߴA�'/-"�j	��Y�����b�1O��D�OR���<��� ���Eb����#��ζ�Z�e�� '�'��'P�'��'rZ(�Ꮥ�|�\���kO+�~������y�Z���������ky�g��[���+�Ne��� �I�bf˗�u|ꓬ?�����?���S?���Q�m q��(1	`��=$C��QU�d�I՟���Zy�8!�J�L�{�aYNi�S=-����	禩�	e�I꟬�ɰgV��t�$͂8��I�KM�D����h�$���'�X��ҡ@��ħ�?i��0�b��.ޖP����!�4� �!�xB�'ib��-Cb�|��P�1sKJ47'��+����](QG�ig�	CyI��4[t�S۟�������@f2�L��I5<�y�����3ʛ��'Br���yB�|���G�	�8*���/�U���M������'��'��D�4�D�OjM`�䃞e����^��s���u���b D}R�|����Of����g\4�'�٠%� 3a������Ɵ$�	.��8H<q���?1�'��}:��-6��{��N0U����4��U֘�	џ��'�rП�К�l8J���SE=��\��i0��H�|R�Od�$�O��Ok,ʪ���H�ʆwb2�i2�_'��ICW¼�	Sy2�'����`���s��Q�&���ӥ�]��sF�<��O��� �$�O���]��<�QTK�7Y�\���]~<ht{P;O�ʓ�?A���?!*Of�#���|JCn\�%��=#rLC�%�9 'Yr}2�'{��|"�'zb�� �.	��Y����JB�Z&�َ+\��?��?Q)O,l95B�H�S5;�Z@��� Bv|��%ŧt��Ȃݴ�?�L>���?�$��K�K��ʤ�"JB5(�b^�O
�n�ş`�	hy"�KW�@�����6����T�����e.��!i�	ϟX���&�6��?�O/��B�E�p��i�B`B�go`@j���6%��z�-��$R �6��|OR��� ��]�*���"�.ZF2����8ö�k���@��tb m��Y���h��%y���'����W���X<t�ꦈ�O��lθy��L��ݬd�`i��.WԾ<�f	˙K�=�'��[5�]�oɶe� �#��	�R�XPq$�pD��kD�L!X�DK��� S�L�ݸL����T��~����&�dl�5�Ō�/D��)�U(ɾ-�bt2�A7	�hӜf�j*�C)+w�	�a�'���'J��a���I�4��lL�]X  ����<5Kf�3d��8�?�w�%.�2 ���3�ןўdJA��2;�>�:�(	�	H����='�$��rm�-#��`�H���S�{� ��ʟ(�����
q�B�O[V����L�@zm�I���=a��R��(�����r���bB�IQ�<1��|�2�R䓵_Ӿ	���\���"|U���$ʛvG\'R��Ɂ��I�d�S��Kg2�'�B�'��ɛa�'�2=�L,���	�b�n��rmqa��`��!+�	���ɉr��'~Z%D~��T�{����KJy��C�H� �NM�0LP?(��'�]�����(6��M��̀K��'��M����?Q���[^m���,1��qP�aچ�hO�?9�E�ꆑ��f	+odƱ�ā�B��D{rA� 3cz���*��8�,t)a�y�Ix�R�D�<)�g�IB������O�:tDC�O�ु#��"MDh���WQR�'��EN�;0@5q�O<i�<!ԧ�8SQ`�0(ߤ5�V�Z� �/B�Q��[W�L#dq����S?��O$�T���ǘ	�i�c�x�|*��$	�B��'5�Ւύ6*x���Lӝ��0u=O�����_�p{&o�$~$��iސZta|23�d�Q6�����A��c��_� ��Dاa�*�o�\��M�$/x���'kbHӷ<�$ŀ�)Dq*�SvD������NRh����ā�Q)J�T>e�|�I*�����/1���Kو�L$���И{U�A#�#r�DA�jȉ�uW�P�J��L?��̌'� 1 �.6�(�숺k#��X��O�d'�"~�I�c�b����38�,�p�#��RB�	0>���9AkJ#?�
��K�aq"<���i>��]1:v� �/�LyY�>F+L0��埤3�@�A����	Ο��I�� QZw��w��9P����vm��y�6#�R���'�
J�4����D��<d��	f'��Q`���!3<���ɢx	�`�s��Q�	Xg��j��I�y���$�z؞xʕ �Rް�����:p�J�`=D������Yr�`�R�5
��HO>����7�M��^;)�hC&EM%`�=X '@'�?����?����l���?i�O(V��R��?k8q�7�G I�����@�`,�)Z4�Ϝr��X�9~� {��0�{�Ē�(�=��gX�q5dh1��N$�Q��	�u���U�U��`��)8`�KY�Z��MI����?y�������02)x�ځg_4N�)�,�YJ!�$�2ӄm�@M9WI�IS�S#2�i}R^�,7�ވ�M��?�-��l# 	�B��#
�S��ȋ����N��d�Ob��J-O&�I����;ٜ)Ö����'8�
(C��K� �pX��E)o�<�Dy�,�
�ָB���43p�Y��0��X��@��4�5s�T Ҫ�L�x
�l��f,�IN�π ^\�A�I7�����Y�1nlY�v"OX�����/
��	4�*d���'�^O��*��ҿk�^��DD�!��A:�9O�ȃG������I�d�OSv�q��'�R�'><��t��0�����"Ԧ%K|(�"��y����Š8_��[c�� .�	����Ͽ��#�<X���tɊ�x��a?}�	��E�1Y�@8)@kJ�(��7��?7��(&�%Wz��߹P�GӏP�BZ�ĊX}(q�C��6x4���#��S��?F����L
�*-M�L�a&�`�<�	rώ�!C����(��Pb�'z�"=�'�?��E��zDa�7\I�AML��?�7���/ʅ�?����?���6��O�|����Ð:Fg��*�0�f��	]ĩ�w�?�X�j�ܟў���P�Wz,���7"�B�l�&@?����#J'��{ �ȺF���Ц����,7j��ԣ���<K��2Pa��1��m��g@��	<��=!��k"n�x��'H%�pR��o�<��g��R�1D�~��;�EEf����i�I�IM����4f.�ðϖ�S�:D�l�9X�:�[���?Y��?a�C�?�?�������"?L*�ܰi��zK�-͢qiA�;0����&Ĵ7Ֆ͘1�6�[ 1��A�<'R�p�!8�`���H�)�R���R�|x�#B�X������٢)��QL>����[�4�
dj���%3������sJ���ȓ����bF�!a�xQ�AO�
0����V�'�����Z�}���@���\è���'@P6�?���) ���l���d��{��@йy�����},��u�S$�`���'e��'g��Sri	�R�0���I"̱�� �}�သ7�9��B�<r1�P�P��G�'�̩� �������D^'A���Û"g6)U"Y#iھ�Rö�����ͳKXx��ҋ\/��H\x���S�S���\?,�L�sMԍ.[z�1�=�y�.�0 "e��,�l�� �����D+��|R��x%�n���gM��)h:0��9�y�ZZ��6��O�$�|�1����?q���?�6OP�:j� ��IX7dl,�b�Eۧe�ƍ�� M���+���2=*��b>�D@�N�l)ʡ�֜OҖI�I�Y/T�(ڻ+�Y�$��@�Y����w�l�����u�r��Ͽ�qj�+���S1 2U��h��΄���p��bQ�F�wӢ��$�矐+g�˲G�&�	&
�����d�d�	[x����Z^�����SA���",�������X�0kװe@ e�'���`�AƟ����8lZh�'���������>�u��')�M_\n����<� � �0�~ݷ��>�l]�A�9A��6���d�|?1KKx�(�R+�Gn��
�m�>��YTK�� R���O���I1D#r飉�H����&��=�~C�("RP���ۄck�1��	�!�6t���4�*�O�TqUWʦ-Kਊ�'�z延f��0U4ɫ���H�I�h��N t�	֟$�':��	�y� E�n.�%(3C�D8R�5�O��1PW���bC���v��?e�P0q@2�O�]�'��6MO�b���yÑ& �z�:W	Y�0t!�W 3�"����F|��	R�=U!���I#v��v���FL2�Hަq$�X+����M����?1*����b�����`��\>�Qs��	Q+@�$�OP�$٤0@$�$$�|B'lN?h�д�
5�p�E�I�',a���^�6�e����0�Ѐ�ӷgQ�`[!�Op`E�a�M�f�*$�#��`�%ƪ�yҀ�1{M^h���On�(i
��0>���x��G�5E�I�0jŬ?�.� ԉC/�y��3(�T6-�Od��|�"���?���?i恇% �, �\0H�g#Q�[�HL�e�>�?��y*��x�t+��+i�H�#�_;R�`�2Ől��iFx���'���
2��Q�"�X
� �	�B9���O�s�&���L��-'\���"OJ�  �� l셲�g�CsNL���	6�HO��O|8� ��_8t�iG�$B�p����O��(��,$D��d�O0���O脭��?�;=��{3��<���ra	)�α�x$Y,���χI����$V�g��H����6f���䐄B��$H�~3n��������$%:�W�^����fυ�4�i����ɋ�M�F�iL�O�Q�Od`��S��$0Wd[�W�SL���'qf)��ƈn_DZ'����s��)ғ8���'剌C���4O�` 9�Ь*k�b�8W��-����?!��?�b#��?������#�?��8v��P'��<WՒ��͔1����I�d��ʓ6�����hk�,R�:h��JdH��Ʀ�ٲ�]9�ƔPA�D
Z~��w�=D�� `1��@�44�A��Q�aڨ�1�"O2��53��e�f*ęi����5O�l�~�J`P�Kٴ�?Y����iS#��H�!�h���rF��r��ʥ��O6�d�O�-"�a �j��1I0�_�^�5s�Ѩ"r&d�F��	5�*�eĀ�Qu&�{��(aQ��[�@�	���`̬g�)z��@3�2 o��rh�L:����6Z<� U+�$y=Q�T����O��}��A ~N�I;X�a�K�<	69k�j����<�~����En�I<W�%8Kz<��bZ~�x'.��<��.]+����O* L�"�'��'�� �d�/�zcw�ݢ�D9pI��S).�`PJ�,���|����jJH�@	^�a��(}:t! )��ņ
�|�y���>E���>~&!�V���bb���A�o����G"�?银iO*7��O�"~��IȊ��Q$ �8y�2�O�Q�������I�6����önP �d�4LD"<yq���?A�IA�H�!
Y<_9|y�%���#|���$y�j=-���ϟ��I֟ �]w�R�'��@�o�:������K?���s�'
�Q��Z1fh�鉽C] �$���Ȁ�ׅ�'q�,�ɴ.��@(t�B��az��L9}P�p+����Q�7�~�[)�?A��'>�`]�Y!p82Eh�D:@��'��lŨkH=���,z� �V�?��|
N>�-�h ��n�84���t�:���k�3d�R�'���'���h��'�r>�$��oR���#4jB���	��[�`�ӰE� z&�(0��ٶ���L8��^q"���P�2�i�H� K4TA�����"ؕf�p��<��e4�MK1D�8:�6 �=9�O�şP�46��*IP�Q%έ��G3f%���7�x��'���?}Bg�D�m�H�ేѱ5z MC��?D���0�+��A�-�e00bB	}���޴�?�+O(�	 	��5��ڟ��Ov��`���:�&�L��4�Ï"FW
������Ij^$�c���0x�&�ŪH:1�������M��H���-K5�+?�NQk���$1<M質�X`�:6���í��R 
I��i g�K��4�G�2yT�$S�O�ZqڂI�F�,��Y3D �
�'Ԯ(z��[���\J�'\%J�4��
�A�' l�!DT�_��@�Q�ļ��؞'��!�jmӞ��O�'$�^�p���?�=�2��P�	������V��W){��T
A'5h�Y�B	�C��D�O61��b	���r�̞�
�qԊ˙.�P��7'� 9���W�z$@�"g�!����K���Ͽ��i֝��� �پZ���S� ݽ:�n�)��c�ɧ��bN�UjDh�f-��~zJEiVÅ��yr��,8�� !�m��Ԡ�
��O��Fz�O���	�dt�h�E�NrƝK�aN2�'�V �Fir�'�'h��]ş�]�S���gc.�:��MU$}�
D@V(�kY.��2��+���k䩤?�Fz��מ"B�F�.s�T�3�Nnɤ%hCG�;2m��%�W�YE�l��O֛�@�5c��u�v�>�1c�H�@�w�G�C~(�M�~?QF
����ۓ
P+`�K���R�j��M�fD����-�2K6S���� i��i>i%�4��A�M;�Ȋh�}�A�Z�v��i�烚�?���?y��0�1���?1�O3qȀj�4�������`H��E��wÎ\A!Ȕ�8hX�@Ń`�L�?1���uԴyp���
���aL>L���5"Ш�R5��G�ti���i4���w�-�'�@�C��"r�V��D2��X�`#]���K��o ~#=i��dҾ�(T0ӫK��]�B�V&Z�!�ċ"0��HSc�Y��;���q������`y�/Ӛ}�7�O����|��#�,N":�!�-)\�T����X? �<ݺ��?��DHRE"�˘��ƿ���xV�Ħ�U�0�A!G�Q�G*��0v9�Vl�9C��:�g�q�hGyb����?�A铿\�J��Q��^��h�.��	��C�ɤ%���HQI��{@�檊�9Ɩ��WO≦T����T.��D�(0�e�7�:�	C�\�C�4�?1����Iz~���O���ϔ^U"�I�Q�g�Hx�"� =��P����2��Mh0�D�0ҴA ��O����w�8K/�>����煘:�I�+I�2�2��LC�0�!E΄�Ģ}���-;He���˂pr��cV?)����Tǟ��<E��TvXa��N���(��Z�*��E�ȓ]
)�fT�h�H@�A�1c�*�Fx��)��|���=�����40 b��JS.w�
���?q@�^�ig��z���?���?y����4��m�5"ٲY�Ad랄o��}��OqӃ.M�m���,�5��� ��w�)`�V$π�xE��#(	��YR�@TF{�b] zQ�Q�a�	:Q�u�s*̋�~�Z��?���'�ѡ�BD5W�V��͏�`�Jm�	��� v�K�/ِjf��r��,H��;V�XA�����|��O !�7�Y)m��vG�%e<}iE$�V!����OJ���O�͚B��O���x>a�"׬R�'��̼��-�4u(�K���St��*�n)�B�FB�@�Dp�Q�����, �(�S�;��V��y��P`����`����i�,Uba�^���'�"��N�F/ցS���''Ù(ҰY� ����y��5|"��)�!��
Xp�7��yb$\�	tڈK���\ �yT���y�HrӶ�On-x����E��П��O�J���Đ?�.H3��%/�A���JF��'�R�Zع������2S������C>�,c�?T5�kΝq�D�Dy���q>�a	�>S��j����q��^�4�j�ڃ%])>���͕���*$H�+qOT�	R�'vH#}��bɨE��`AE#ъ"g0�C��AK�<�DE�xf�-:��]�"��D�J<!�����U71U��IP��<)V�E&*�6�'b[>q�_���	�����7,\�ݻ���L�|��!,�=[�c�M��e�g��=
j`��1��+���.����tA��� T�P�K�e�1X�* ���eN¼#��X�v�zC��&(Ĭ;>�P���h�K��wt"$�B��5@�����0&�z��Aǂ2(e��'��)�	�OJ˓9�d3���	W8��$��PJ\x��I������rY]�a���w��Fx�1ғn���'b�5)!�ƈ7�L�@#�
N�Qф�'#�'[֢T{��'"�'�s��������!��s0 �L��H�a׍�j�g�"mPM�7ř(w6��S�'�r�Q��o�(��˜�32�qcۅe�t����s���r�,����i���������q��e�5�>m��`�@k�)p�ċ�YX"F;lOJ��V튢;�&x�׈���5"O�,���R&-S����E��(k��5�}���d�|�I6M^㸭�� ǕnA2Tc���%In���O8�$�O�PS�d�O���o>z��.o�Hᤪ��2ƀ݊�ᇝL��8�,ƶ?a61�pʖ7aw�`Dҡ�,/�&���;zy&�ɂcd����!�_MN���!L�[Gv�A��ie�d���E���'o4�R�a�vNf�x�5�W"X���dMٷ*��6�3��/�H���4.�ÓF�&��s(�+9!�dE0t���hƯ�6J@=bٝW�������y�
�*F�7��Or�$�|��l]�B.�=I��
]cP0`g�D�w(�s���?��~Q��[@7pH�0�/�ZP��GV?MS֪y��M���ЁG'����1�;P��R6��J�4ٙu�]t'j�Zw�r��7	Q�o>����D�=��Q2o��F���`�{��V��?���)	t�戡��7va��y��
*D�!�X	�8��E1%.n4�e$�ha|�L&��mm.�@X1gŬ��sC�pJ�d֙J�o����Z��A`�"�'D���
y�Z�JP�$ �|k���+%����'�1O�3�G�4�)�j��=���3�����.�p�����O?��
aN��4J��j������<�H�0���O�$�"~���_91h�]��H�9��@�/�C�	�-�`H�cӝ0:D��ChT0
B"<��)ڧO��T4C�oZ�$�b�f�?�?��.mDAre���?����?i�)���O�΅�b(��jƉ��ij�I��0����(xh�}�J*5F�*�'O�$�ЀJ6#'�~B�X��>�7��[�~ ;�f-䘊��c?	��ȟ  �|��)J� �6���3�J�+A�6ͅ�c��I�ţ�^�z��g���̈́���)�'W����i~6s��Ŗ7{X�&�L�f1��'?��'B�AϯQtR�')�	Pz}�|Z�+7Šb��zn�x�WA�J�����]�����|���/�pD�؊wt4���.R��:����)�^5y@΃O�ʑ{©�K�,5�=ٔ	��ЊߴH�^L��\�n?T��g��+)�����T�,�p���j�i�˫=�xP��V��y�G�A12q�Y�e.=Z��;�V�|r�J�t6��O���|z��~�6p�S��=�hQ�C�߈yv���?���4c$=�������@�D��1��C��	c�% �q�Q�cDM,��M��`��I�=�:����m<�5Gy��Y��?���iF��;���%]}z=�nK�llC�ɛAƺd����F5gΙN����Dw�I�����,+4��Q猿Tt��ɋaH
�zٴ�?)������9j�T���O:��Y�e����5�2#����B�o�)#5�E�f�6�Z1	-���|���B-��v��tF�D�2K��@x� ��V�S�I2�H��D�"�G�u^�.1x�:�� �~�]0R>T鐭��BI�۔mq�tT9c�Cԟ|�<E��d{bԲՅ���*w.��H�ȓRFԑU*J�T@�U�$������4�H�� �!�F#<��)����PCXDHRA�O��$��^}���b��O����O��d���3�Ӽ㖡 �}t�u`�n�b�0�~?�a)Zx��;g�J1��Uk��6h3j9�Χ���(6�O��c�!~�@��>��`��O ����'����d�,���B� M�||���&S!�E- ���m�e�@� �7OӦ�Fz��ͤ�n mں�&� "����.��f�L�����I����3fD������|�Q�L�+4�hJ���<O�4�8��r(>�9���
5D`�HWsSB[��Ɋk��(�͞�d�����K2d��Xq��@j�rI�,ߥyzj�Z�4����k\�P��<�dJ�q��e|�DhC�
�x��2g�,c���'I^�����Lyr�'��O��
��ѱc��pȜ���ژ6��B��'nʈ�T��<�|�����o����5�����_y"�� e�����	~�DI�&ͩ��#�0u�82h&<���'+2�'�4B�`Bs�M��$K�-T�T>�b6�	?g֮�0fm@ve���I ʓ_��`c���$T�4DAuk@L�Y�n��_�z@�rOE���Q���D~<�s�K���$���O��G����
<�1(��quf���y"*'�$�6�ӎ�X((���0>a2�x�/Q�7���Z6��0�4Q�O���y�P�7�O���|zg�ǉ�?���?�&I�J6ڑ��K�1q���()Ld�gc��Y�E]�N�=���?Y�|�'[-��$j
�`����k�,Lyfq�'DW A���:�5A�Dp��lJ���?Y��,�7E]�TT����=�t�b.X�iSڅH�'�1O?�d@X�V�+a͘Mz�5eŖ8"!򤋊T�F܊f;jgL����\8��4����:1q5��D�3i(�a#�/���F�D�O*h�F� �=�����O����O�e���?ͻG���`¡��$<@�bCˍ(�]�fN��7T�k��٢Ҝ�;Ҧ�}ڊ�ׇ@i�e�W�A��`(�E�������<M8<<9#ȹ)��� Gޟ<i�Ǚ04���O�X��m]��R�+T���9��|�d�Od� ��'�.��d�<nH�0�@Jܥ^��i�G隳F!��L3d:�1���{���!��H��0�Dz�O�'���Sԇy���Y��W(�����ԧ0�I��F�O����On��>/j�	�O�S7 ��eb���.��|��BL0�t-дI�f�(���.xA��p"��O"ɫtDɭV�r�ڸf,T\�r��)_D~0��33���D��T�Us�ʈi�L��%6�䊈i�BKv�@]��N@�t����2Pcz��a	��IAy��'t�O�S�"��3n͆�TQzU�T8���<ړ=��1��kӴ1f�P#X��\d�L@�&�'y�	6'��
ڴ�?9����)@*S q����_A��n�\j�0Հ�OF���O!�"��aiZA���
m38Cƈ\J�D@ܩ��9���9��Tqf��.�(O~ k��!%آL@��� +�������b�QS�`�}�CeoY�f>)�Ʈ�
 }�%�C��
 �+n� �'>����ԑuP
[Q�ӦÅ/"��	V��|"����k�
܀T��b>�c`��6���A����|��m�̟��� ��,C7�'�L2P�y�̻"eE��M����?I-�F�`���OH���O����TW����"�cꎤQ��.xC����A�?u�-K��\��@�Ob1���(2h"���'
�p�EՏ�0C� N����<L�5Y��Ũ쀐�!�:r��ߝR��6y����p@>�, �7@ͩ&��q�It�S��?q���2,��S/	�E�v�C�`n�<����^�S��;r�f�C��i��?��i>��	0 ���J�,U��@��B�ȟ$��5vZ�	6�����	ʟ�ɣ�u���yW���v)��1�G�0p�d`&�^��y����T
�I�Q��y�
P}����B�W�\1;�٦!��y����4��pd��(���+�O��XiB/
$k��+fΧ<���'�՟x"����<�c��M�gy2�iw��r�ah��Gk��<i�nךG5HX�ȓQ��x1�n٬I$��`a��BW��¿i��7�OT�G�B��@yR� 8/���<1
`"r�\眬(�˂Rx$��I�����Ο�cs���l�	�|�$6��x2å����쀵Y�V�B�Տw�Ĉi�3��<y�oؖw�6)A![]_���W&��"?�xJ2N -xB��#S�A�L��d;��١@*�I�C�����-��LL�]w�H���*5�(]��2D���.��Ҵ�U�x��C�E�;c!��$޶u�5E��e����1�Ȧm'���'����M����?a+��UZe�����We�#rΘ�2/ۤU ����O��κ�xMZ� �:d��'C):`�'&�Y7ň�<�|1Fy�ۻq)z�+�YGF��L~���	�/c�BS	��K���Xc^�'�2�Y���?��?+�ȵ&'�	�8���$ʚ���O�"~Γ�̀hn�4M��U�ō<͖���	���n�@��Æ��o,���	T�f}ϓc��8���i�'���
P�I��ɟ��)� �h1E(B>C>n	[�OJ�<P�JLg��42���5���4Bڦ��O���y"��%�h�a'U3s����Q
B�Nf��ψ@�ԉ���D�4�Ą��&1���d,ٯ����l$���_ �Z���l�����"mD�$@�qaش�?���'-�d�C�C4��;�aDP�0(�'t2P����I�*&L�C#֜nB������y2|�<iش>C��|�E<��� <�����X�S�]�m���'
��s�%S�<��'���'��������wu&�b@�	b[t1��S_��x�Aί,!VC�(Ip������?�y��<f�`������V-�Dz�4t�(Ydݗ`J(=x',�?bEi� /����Q�g}���HYv\����<G{�=��-V��~�cJ<�?I�����DR�L)<
���O�����\%2G,3hP��h���F�i>�$�������M{!^3����(�A�Аrc^�?����?�_���\���|j`�H�a,rԨ۴U)2�I�
��X�`a�G����&Jƈ��bӦ9�5�C��fL��H��C�D���,�O
%�' n7�ա+!d��t/U�<0Ԉǁ�v��n͟�'1���?����r ���gA&�
@Z��4D�8q�c��W/@�[��@ iN�sw�x��O�˓G�����i�b�'��%� :D�G��1��A2B	$������ğTXӥ���,�<�O��%��O |u3��-�3�� ��?i���0>WƠˤ��(5�)H�7�W~py�	2�H�(��L�tP$Ȕ�Bd� �d"ON�XV�ܡ�=���>D;�'HrO2�J�ǩm����T* �Kq�r2O.��Bmۦ)�	��O4H���'���'���K1�61%2T�-�>���rwE�� �Z�n۔cx*�Hb>�$�"�֨õ��3qM����:��P1�:jBXJ�ܼOL���P-ۄ�2d�+?���MzuRZ9XE蓤G�-h��T�P����'�1O?��ܲ2ҁI�E7V+�A�b��5�!�D[�p|@�!o9%���� ܶ��| ��4����B�*�
c��aa$�V�[
���O`�¡] ��D�O���O( ���?ͻ`�eH���U�x|�A�=MB�Yr�'���x��Å)�����	@F{K\�~\���*ɮL�L�('�N0s�,���gO�x�tTs���|���O�@r��Z�O��,�'7.��G�#�&�pw��:B�ڼ��'?B����0>I��Qka�+�0-�U
"�-D��f�V�vN@�آ�Ӕv-�����HO�	#��w`���A��f5���.04�4m��
Iޟ��I�@�ɩ~W���Iڟ�Χ��뗣'�4�1Vj�^���0���$?Tj'O U�f\���t���� c�\�NT@xeś,L�N���.Q�+1bN]|���	"�M��#�:pM�L1㬃?��sI�\�Iҟ�%.�?8��+�E(�PXyS�?D��R#�Д"!>�R�c+xڵ�;D��p��I�E	�(j�F6� �,z���۴��O^��(U�i���'�ө �^�q
�w�)�_"
'�lAtGEٟD��ʟd����DT��G��)�S���A��&�H��Jn��'肱�(O��ڴ�A���<�c`FZ}h��Ďl����
M�I�Hq�G��Cw������6. U��)%�������K�O��,K��Ď(�h��C�9|�̍b�'�ʼqR4zY� ��7r��:�/A�'<<{� ]&A�����^ 4����'i�����q�h���O�ʧ$D�����?1��z�Z��A�ժ���{�W���*M�.$���6ud��h���2F���A���-���2��9�T",p,�M���Ѣ:ﶼP��*\V��#�D֤]~�q�+�H�c�����wEy��?7L�5mK�lBq�S��+�!���OR�b� ڸ56�!Eƌ|�5��"O�� �/�`�HH$
�=�4����O�IDz�O@��Yo��yA�e�D�5F ���'��]�㙛_bR�'�2�'��]ڟ�����V�W��*(�&-T�A1�Ÿ3�-�%��ϩZ�B���?AR��䙠c�PԑW	��	�$hgɵ/ٞ��
E�w��Ls0�E�h^�Pӱڟdt��@W�6/R��QB�>Af�@�&��a��4gl�@6%�j?	1n��1ۓ�>�볫ԉu�������|=����?�����o٢��'�ϯ\ֺѩ֎C�đ��w�I>`d���4_��<�%D+`ئ��J��ٹ���?q���?����?���?�։R@�nu�6��J&�A��&�PP���L�\���g�
3�p�"A�)�Pqs�o�$��@�e�wE\YBOœt��Q����rjFi�����T�՞y� x��:�䕞y�R�z�6�ЧE	?H����M�N��%�0d�ڦ=�IQy2�'A�@��}���r�.Fk�PO�6��I��IV�'?D�Z'��5�>0����<���H�'Zt7�	��ї'B6�P�fwӎ�$�O�'ZD���V��	�h�!�CH�|A��9�?���?��@��?��y*�� ��t�[�Z�� (��Մ}Z(08���t F�*VM�4z�B�
��]�Kt�� "ZK�''����*ۑ>��6�Q�D��D�V��~+-1�c$D�Qb��9AY6ؗ�(D��	Rc%�O��%�ʅ U`D�k�,bq �N$D�08rA�0s�1�Fe��ZR�"#D�|�ড়�W)(�� B�P �aY� D����]�@��Uà�[L���h<D�d�O�U0z�JXpՀ! �?D�0��@�d�B=��b�J�~�Cw�>D��s�аj#�����-_�����<D�h�cԇXI�R�P �%
po;D��g�'B������=L�ʄ��8D��'I2ݘ��0�7��K�d6D����3@`m�i	�Ȉ����3D����l��'ϚpkW�ǎK������2D���b)�'X杣։�w:L�9�0D��st��>����DE�>� ���/D��lH�V2�ư`��axp"D��򒤉q�n�çM� +E�2��?D����剠
�J�z'��+yh�I�F<D��4$Q�I��� �=)4�[��&D�D�����T��w��>+?x�r�/D���B��rs�Yi3�\0E Uڳl!D��ꅛm9�e���F8@���1�#D�(���T��
R��iU ɺ�$D���p"<v�l�T`�ɢKk�<�T'���T(��a�>i<,�7-�c�<	!L��3�b,����tK0��pf�`�<	��ӯO�us�O	 L�89��G�<��8f`�t�����k���CF�<�$��6L�Sg���hڔK�M�<���j'd�S2���G�QM�<i�!ԆG�B�PG��_
�d�r�Ma�<�'��4e 
��2I�7���Z��D�<1àY�����^!%�̄2�v�<��K��J���3r@HyȔ�M�h?��hħT�<!�����%�|�<���G��]'l4��� �AZ��0r� �1B�C. ���E|��̨�a��">�Qӑf �O� �Zń<Vi�!��]�Q��i�6 �X�w� )!1F��tH8 @��~3�8�c �2R㑞֝Ei�qB� �	z}f�s���OΙ������w�pu���#��'��)��d�~�sƜ�/?����1��1�5�Bc�@�*O�AQ�`�<Jь -�~uf(�ا�&ٖc���!"�d�)��/��/R�$�ZwH�y᧕(Q���"WD�ty��IE�u"�'�E���"EÂN�:ؓP�Mb�RP�>�g�mW��y��'p�A
Q�ޏ_�*��vM��W��x��P����!���HO��O����N]�o�0���I�?�h�'_f` G��ɖ�y��I������]��jE#l�cB(�I�XQ�D(��kvV�
fs�e�qj��ǧ�:����t�$�"s"0�I.x�;�(�W���K: �[4���ݢW�B�
!m�0,������[~�"-���6^�	�"��yB���=x����q�𱚲8�Ḅ'�X��i� �!u�11���٢������>7J�A7+��Ķ�qV�N�"N��w��<43b��>�g�;��y�3�ߖ\a�Xv��< ���C�7|C�L���ߨ%�j���Bk��u�w���)C�b:�񲗌�+$�4��H�d�a'	E�S��$}�Dͦ����%��P[f���KD�E��m���*��?��!��5�f���CT��n�%A�9�$��?Į���@͍#�qOFHr���{>)"��t�Ϧ�<RЉ͊N��q9d���A��mS�ƭ>���K����g�2w�(��n5��?}��ֺy������D����F�ٗ�OH9�;V0��)A���H�<%hP�<a�k��;&�}4�����!��0&8�H�g�ˇ�O�>��B��J��cu�/I���$k{ӈ�tK�>,��a+�dl����O�k[=n�ѥ�Vs��Q3e�W-M��vf��Ey�'�ē�Ra��/��t�0Hi��	h�0�(�'��(O��'м40Ik�
)(0��jA�&$J/1�l�Zq�͊pY �?Y&;��?1BF�PHgx��r�@�j za�̼����O��T�+;��\�GL���OX�W��8.j$\ZC�J0\� p�	�r��pS'��:���_�� �5�o�*Si�"C�E��+H#q���D٫�����H�K��Ċg��m���8_�B\��.F[_mQ���^�ʑ��e�Ƚ"5"*j��q�����'\�z"���~(S�D��`�|��%P:��i��R��AA6��GQ���>W.�}���Ab`�r��%?rJ#=��{�R�����6��:����]�̡*&B��)4� �';��AQD�8)�h	�'�O���X�21"B)�\���CBJǤ{��7�FF򉮉�1
	f��r�2��/+��Pe�=|הJ�'�%0�����)ʮI����sE)�?c����0o2]�lš�jaâ�ܻ�`|�.�HVh�l�Q��ݛG����M�@*��LЛ^��'Ur����ñ=b�R �Rz(�����r�8ُ�_�`�0`(��B�Y�I#3�w�9�d�J�N r�Ӏq������d��J���O�p���u��S�H,��i�(��}���N0�DA{�p{�fѠW�*�=�S�k�������lDy�K�3nW����{��	�kV���W|ڼ��꒭h�~�'�`UA�.n���[�D�)d���� F54@����C�������}FP_� i�'JI�=�V���� �&:"��r�%��/�� E}�wC����@%��LB0�:ռ9�L�d��hz�S�'=tb2J����H���9c���I'�f#�h�Ud�]N��A5.���(�I݌�	r!k��'D�c���X�bg��ʌ{��?�Wă�Ywr����� *9\��
���`��Or��g�M5�b@��^�V�T@��Oa�0�� BΙ�E	P�Sԑx�9�ɯi�H=�;F��| H�>( �N�\Vk�)!���d�<W�R�bW��5!5��pj͟ �V��D�M���� ^ �p���S<��ڀ 
N �T�1m~<��4頻�-$\|�#�۹2Ѻ�{A^�<y����'���Eі0��Yp
�w��"?�d-D=h
��� �آ� ��Y�$���ףs;�)�*��s"F��dWe\�0pFԨ`�pT��l�*�(	�� ��H@� P�G}�Ik��E��:[�L!Ua�˓��$�FM���ͨH��q�f*-J�d�<���D"��%�hш	�AT�ɲ'�������t�t"�U�L̬-y�È�ZH-C��P����9�8`�Lâ
4�Xp�$F֣M�H܀��l��A%�7�d<����0�B3�Ry	�{�!��'@�B��+|OZ�[�80� ճj!=k0�Q��ZĲ	ǓO���q�ebX�,p2�
�1cb&F�$�^E���ʴ��OR �'�$#�"��4֦�m�qU��ya�:zb�S���mT�m�J<i#�%[��b?���E#"3�
#Y��	Z��>ugܼ��"}�V�~�f���!B*O�N��- ��''��Ғ0�3�D�7�$
�F��\�����K��W�'9��9'#�f8���T-[��]��+Q�x$`���9��Ѱ��'d�)6�􀩔��&h��#��D���I�>��Hf�|�O@�/� Q�M^�A�U����OB|� �����Oz�!�C� v�����˔*�\�K<�aO÷iՄ�b?��C);���8���~+�����>��D�|ݘ�"}�#ؑ0��* ��{�*X��hS�M;n���a�t��<��ɓY[���D�)euF�Sr�T/�=��M@
��6�ި?��(���"��|�l���vP��HR?�����HG�<�֋I40�g�����DJf���Z�k�=$�d�8RH�1I:��Tl5a���B��c�v@E}�\��b�b��p��P�N��J�d.�v����]p��xbLk�0-��D�2��M��h����>�fk��? <�0嗗�����R?),O0����eWl����g����|rLB	[��0��ieجp�KV�2G$e���N/��R�'���B� Hi1R� �)�z������%�+�/q��6�7�ӼP��e�0��%� -®�Hf�KT�<�B+��XS·�x_����DQ:l4B�>a��%a|y���m�����/�
viñf��eQ��<]��IP�~�����K��p�a�,`��#�ۜPD�P`o�U~2O �y!��#���k6-�A��׸�JBjI�[�*��A%��Cr e����d$qO�aÀhi�-+t�C%7����u@@�Ę�9S��` �����ł6V ���7--Fr܀(��ԟ�O��	�n��>8�!͞L;|Y�T��� n�[��A���˰ˇ���O��U �65zUhŁN��r�ܯ��ɪC<=�?���!(���SaF��h�ƥ�K� p�x�>�&c�U����eL*1t	��T�d�a��+��e�U�yWP=�=1�"՜�'�j��)� �lP�n�u!�B���|�����D�B�2���)1;{���eP�n�qO�TK��jٓ/�&ƺ`1dE5T���ºӕiQ`��x��H7��'ě&��(���
0�	xg�xf�Q�)2���,�?c�� �����^�ob8(r��2����Ch�+k�j�.��b�H,� ���O�NI�=D�{ �u��1'ԂM���A�Oԩ)�L��XG��'���j��P(L�� �E�[�e�𩲀�M�'��pe����[b�
˿kf�h��0Pg�%	|l���X�T�.!�d�	#56���6|��(J�O�RX��B��L);�OA�H{쐹��R�X�����#wOͅ1�ʓ=ʚD�e��-W��	!#�O���c��Q�h2��=�i!t�i��O$U�'W0�8A��9|��Ox�	a�!�<�B�ֿ`[�hǌ��PV��5�~�`H+F�L���S��>�IQH�Ca\T�����&�Xq l�~}�R�L�|�2u͚# ;��֝�T��j�J�N<	0g�םP��@���&� ����P?�dP���'OH(02әm�idOZ�Fpj�"c�Q��	ùV��k`_$o�D��X�(�2�*ґG'6��K��,���w�=�=8�f[��p<i�'�.tJ�)���$0��+Puġj�V�$��hM�M�X��'E�u%�$<`#jL�EM/`Z�*��;H����:
�(B���3M�
�E~BJ^�L��S4O"~E�h�'Dq��(W���@�̏�W�0؆H	�h�pٴ<���s�V"����"<ڧ%�ؽc�� �V<Bwm�"p��V�܁
$d�4W) S)L��(O�D��;f�D<rfE�qd:eoFYD� �J�1C��,Q�2��7'�><��O��d�xbi�]4~aӥ#y�h�DE�
�I�A��~`ѡ+49Rj�LU�J��I�g��2.�|HB��6fr��Gg�x����Ύ6 ��ac"=?��"<�'xq��@��)	�bp��F�*	ef�[�ѣ5k�ɗw*VH*7ΪM�[w�$ ���J�m���7ȑU�.�	';;���׎ӒDr8��_�BG�'L�֝�]K��i�a�*b��x�W�Ђ�LY% rA��Zh�
�hL�T d(�_� �0"���`���@AU�Oł�b'H����B�CeX�)T,Ha�q0D�D�\.�;P�U�EQ���w�rݠ�hC4S �ɒ�e�ou��)�n¦D2ƍi�������O��'��x�悚	qL�Iw��uP�W>�<iq���Cɔ�4�PX��O�Mp�9���{�Qd_i�`�h����J�A�U��0���r&�Iaz�W#���%�ةm_�EJ���-��$f���|	��:���,g6|B�%�w�	�d�����f�3O���c��,{���m�i��Ȳ�+fNH�i��n�����j�2{ɶ��F	�,����2��>,�(��d�-����	cZ���f�	�i�K?Ͱ������<1�Rg�B���$�,[��X�$F�3P�(4r�$T�[�b�=��wR�q�R�ȃ��2��H!�$�HX'V,p: rR(%�l��Q�(p���T9+���������'a(�<��i(L����!	{:�J����]m_�T��� 0O
�舳�Ӆ�veH].@s��?�'H��銷G�.{f`! A��;,��)��ۮz�� I*��cuG^�__v�ҧe�s0�&M��[�n�*��Þy����\�F1:�C��}D�1�0\�ΤFx��l�5���� ]����'���!p�Ic6� @FK҂#��j��
�e3b� $4$,Γy�11�DP&�MG���77�]s��9d��b0B�Z=yqg'�w�J�A��	F�t����i�=��ڀ0��L1/<u���5J�x��!3��q��C�(O���
���;E�01I� g�� ��-�(J���QP��hOR1��I{�lt�0�q��đ�@2��b�N3
;&-���+_�Op�s�G:eb��F�&�vc>�'؈���.���IIEbޞXX!�dI�;A�͗b檘+aû);!�\�C(]�t=$̓��Vf$!��1R�8�fE�,VՉ�� �1!��Z�5��AI��@�
\���J�^-!�Bi���?8���g�!�dE�p¥v�Ap)�\��X�!�d�)B�BLy Gv�Ka$�!�\�.��xbS���)��-���M�?�!�d)b��c��&�}#&bW��!���,���6Pf����ċR{!���5ZȰ��@�\�ը���Ul!��P�7��\۱aL���R�J<=R!�D�=7aЉ��!D��`�C���X�!������f�ɯ:��%+6�Р@�!�M�),E����Eq�2���
�!���1{�K��0꘤a�`�z��`�	�'2������b�����X�Id�
�'��Yq&͆�I|��#���O�4��	�'��I�C�^�6u!B�_e*�J
�'�NEb������F��d�	�	�'2r\��a��
�ڴ�3a��g	�	�'(J�kI:e+�YPT镩a����'C-��2`$^-s���,b�h��'�X<[�ԙ����U��p���� �9r��	a朘­�,�|i��"OҐ�a��jX�葑���}��"O\%��R�3J�$a��� .~��c�"O� ��
�zi�p�ޟ"tvP
�"ObH l]�@�9D��^M��Ad"O�a��Vcz�q�4���e=��
@"O~xʰJ�0�Z`�F�D:�a��"O����Np`��e�-5 ��BP"O�,JS�(c{z|�Ҡ�35�V� �"O\�G�\�Eֹ�_�t�z1x�"Oܘ��`M�k$�u�W��HH"O6���lF�5ij���I2Q~� xr"O�EI��&���CM�x�(�y�"O��P@ջg�@��QkǱ
���(�"O��e�x��ԡ�'�At���"OVX)4�˝:b����*Jz%��"Od�Q���h)��ފ�%"O9T��L�(*��_�Z��M��"O&D�@���I��5�u�P60��"O@Ad�Q����C̐A�xY�#"OT8Ƀ��t�~]P�/��Y�� �"O� ����%,�$�^���c"O���!�Ffi��D8�z��W"O���@'��~n�6��8�ҕKs"OBtA��]�ԥ$~�ҭ��͍�y5�|J�e�*e���E���y��X�,������ � �P��y��B�w�0�[,�i �8W�I��y����n(��Kg��br����ך�yRN�:�4p[���@��
E.�%�y")�[����"ޝ��31�J��y�E\�Dh�yS�j�7�Z�`���yH�(ԑ�coM�Y���)�I��y2g�6�(��+~%|Ā��(�y�FH����h�&s��\;vm��y�Ei�Dbu��<]��Y"�BѦ�ybl�"yn�T��FC�W�&�K�.��y����A��@p�� ��IM�yr��MT�����/d�ÁL�y�a���.,@�cԮά�QB�2�yr 6Y� QAQ!ĨP��ub����y��"K�"�Pa}(r�IX��y"#�`np|�R�]1%�ȹ� �y���:YĴ8��ttS �Q<�y"��\�z���*��T%���y�nM	1N�O&hײq+���y��#�4��d��/e��	�B�T�y2�	4�h�r�(��F;�{"+ܔ�y�O��Wg��Z$�L2k��!��I�yҩ�8�{��Y9f8jI�&���~��D.O��斈O�i�ak-�ڸ���'��I�h���)C5�j�h���W#RB�ɰrsI*��S
N�a�Y�{��C�ɧ[�V1�� �j��=�E�c1�B�	�f':Y`�@�]m��ˇΐ;1ydB䉏V���"M�L� @����$B�r����5NÃ[d�qRI�,��#=A��T?1���I�HXHU���J�X5���-D��;q�.D�Bc������%'*D�<BF�#�����'ةC�@	�&)D������ x���ևV��MCu�%D��r�Ǔ2���3�IՒ%Ҷ���$��p<9�G�4�(�1ƩM��)T��L�<a�gJ� 
 cA�$�~��u��F!�� �x#�Ɉx���G�\�U��"OPH@�c� K1`�����.!��H��>P�'���+��=w���p�G�
Lx-z�y��)�� ?���-�<ӎ�p�,��j`�C��!9a��Fƕ(�+E�/!ќC�I|:��K����h�'/Y41�z#<��%g����NG'�Ёa�.)�&�ȓDE�u2a��B/�P��'1pB��ȓ;����F�1Zf���$�ܯ_
�nڈ|p���J ��F_%�����F��y��
��*9It��<
�r�����'��{�'���S݁	� lze?�yo�FN�(�O�{7�Ǿ��'��z�$��O�M�&n�|ϖ��B���'����剿6e.uه�M 0p�eb�PDF���<?q�	@+daP<��ؔ}	t�J�<	f��*I!0���hTw[����L�<��#��f�UQ�k�k���)E�|�<�U�A��c&�`ؑ��s�<��g�X3Z|�R�HV{�}z��Tn�<q�	�� �
��O�)rSF�
&�C�'��/ʧ~�v�2G�;|�� 2FA��?S����_���CḶ�r���u���\��%�TF��'s�!��K7 >�D��ŀ�@��yb�L7^��dj��I��8K�BT��y
Ĳ\z��FiH<_�1��
ҝ�(Oģ=�O�ݹ2���U�9@C�W)O����'&2�����j ̨�"σ�YH�'�ўb>��'�٨�L�QA �+U=<XDU�'��DRĵp)��MiQѡ����D�Mݸ���쮨j�떼C�D|���N8�O��=�O�BE�?�J[��5T2\؇j�2�yR��4U#\AkE��*N�t9rj[�O����ױ0K	ox*��f�T��'� ӣ+�^X��#�Z�Oz1��'�j��S���LH��E�I�f%��'��0h�J�nB�	ڕi�	bLH�'y�zU�D)]#�����Q\�`1�'F, *1�R�"|��B$AZ�Hi��!�'���uߨrzn��D�4�h��'R����8M+>�Z�����"���'&`�#��#��Z�k��rZ�'�vp�G�{L��k�*<
�'��僌�;��, 3�̤
Nj���'ܞaz3�v����k����'.Ё�g��x�
uϘ(uN[��'O&�#U�]O�!��l؀uC����'�̐C�@��[Z^=�� �z 4�@�'Ƭ�9��?�)��kU,z5��O���DԼY?�aZb*�1F{��B !F1�!�ċ0Fpvp��̕r�l��/�6����>��Іk�DlP�ʑ� s��t��k�<���')�z�ʔh@+Ib�����j�<���� �P�&���J� ȈW��n�'�ў�'fP�Ub2`[�e����ƛG�X͆�~�Ƞ���S�����LI-ZDa���:��sn�7��8+��[�=4��ȓ��Иd�I�?��!ٶEr-��h3z�S� ��X�d�0X��Їȓ q��Qr���?>�]�s��*1�4$����%U(,�h"��D0����� *�B�����)�!e2�#�����a3�j"D�0��_�O>j�Sg�掁2n>�O���?9T�	�N]�zU�H�+�=���z8��%�� �ԋ�'8�P�]��a��>����i]�z��pxdTp੸1GS��!�d#ܞ�Y���7]g�tre��?8!�d�� �4-3�Q��,��$�2K4!�$�)�l�%��X���ӣ�,F!�$��aʩ��dP�	rNj􃓷|�!�䖞z��C�.C*aF1����=�!�Dȏ{�ǌ/X��+�KƐn���'�O��f�dD������n��m� "O0�r�ڽDny W#�g�L��"O�h�1F��k�!C�/A�,�"����AX����h��gZf�ۦg7K��99E1D�4�Vj}�p��pC�'Q���`�i-D� c�c�4E7XU�����:N�
��*D�\��OS�(]P��Ș9@Q`W��OVB�	%w������%�&Ց��S?�C�I8��D`٦n�"A���M�zc�TD{��O�a�%*��lLL���.��(O��D�,O��S���0�,š7mC0)t��U"O8T��ON d��)ua����W"O�x�aEK9N¾�1�ϘK�9XA"OT5�f��P����R��w��]��"O�����3ER�����1)8ݲu�	{����ˮs���f��N���'��d!�ۊk[ȼV/lԼ�1)�4@�O�6-1��?=�'��$:łB0}� �䈪<"�H��'32��"��)�u!8"��O�"?�`>��6,���梃�5;�'K�*����+�I*7�CڸZ��5ic� ����y"��Si'��N\�fGx�8dF@'P��B�*(�J��F�r�X�R�jr�"=�	Ǔ�J ���_�O�t��,H�jC����e�XP�ϗ�:Eb$�<_.�,s	�'����妆T'�����f��i
�'ӄ��d�3K)����)X�($`��	�'������+\�b1���#!��	�'w�Y�p�U cs)21J�3�p�A�'Z�@ ��K��M�P"�	����'!&�S��y�j�I��I�$	G:1@����y�� `���%=���!d��l�<	cI�3*,8�o3!M�4����]8�l�by2&��(��9���9'M���1�y��H�� P	�� Y���4A��yB�˜c�m�a��n�Zbdb��y®Fg>��1�	C�m��Q�Gӆ�y�,� R�y �`��p��.��y"Co^�����F���rh �yB�ñ��A��P&��s��Y�y�ꘗ	6hI��(��&��IO��y�`LbL�v�ȗz��X��ۿ�y�ңl�)�tH�B��V�y�'�f,���2��C@C�E�	��'�~�Q��S�b���P�)~"��'\lHׂ^�]x�Μ��%��'��8XTb �HG0��s@݁%%�Ii�'�<Ӵ�@5x�ܕ#s/
θ�C�'��]3�'&���L�n��'��yFaU)�h	z�4��'7��j�a�J��؛��C^b5�	�'��˫n�,���P0 ��B	�'��� ��J�e��f�J�0���'>�]��E�Zn ܑa��Hg�:�'����B4$e,U� ��G��z�'�D2s��77az�0�H[�0��1
��� hHq��ܳ[ .��v��vI�a0!"Ox��Qꙟi���2UO֑J@ %��"Ot����6�v]*U�W�_@�Q�"O����&�q$���h� "�P�"O�X�A��L!fIS��+Q��j@"O&Yp!%L�{!��r������"Odhՠ�7L��b�-���	ڐ"OhP0���
7��X��C%^�0��"Oh�0Z�4��]׀�i�"Oȭy�)W,Z�>�#у��N�""O�����0H�L�7�C��0�RT"O����G�!^$`���.���"OpP� ]����A%�4�p��#"O����	�'KΦ�����/���A"O�����$ӌ��f
�j�
Ao"O�q@�"z�p���X'����"OF-[t놾6C@�q��6$f�Aq"O:@�bԶz���IUcU�[��0h#"OP�m��z�|�x2�8f����"O��r��$!�q��U//��2"Or��FP;X��jGHĿD��\{"O�9�d�AU'��eB*�МJ�"O���2���w�`��ǭ{�4��"O�d���'uy����b��V��4��"O>Ix���8R$���wn��s"Ov����'Y��Q "Đti:�8�"OH8ST���}Z&�]�rnJՓQ"O�q���Qq�M�ԌI�z��� "O�����S�P)aƓfuP�YE"O�PJ��ń+� ݈�#Bf7Zxi"O̔L'9�l]�Â��e�$���"O�ȘsM���b4B	X���y�"O��ap��C[T���R2{:�Yq"O�L�rl�)��9"�gQd(�"OFY���Z.@�
V�+IP̐7"O�ղ�գj�ꨀGGJ�CJ�Q"O������b�D	�^�M6�S�"O2��"�\+�mX�j��N
6�I�"O�H�+Hf*u���!r)kq"O}yҩP�\��=CEʅ!h�0�"OΌ�`��+:�#b���#�LX�"O|�s��'yq6�**�YBF"OIu�X��@� ��sݜ���"O^�35eY.��`(�+`$�k4"O�y�Ү�29>x Cf$�
vM�i�"O
��Qk�M��00�ʱ_��s"Oh�{�F٦ΰ	�g���Y�쑢U"Oܘ� hŀ.��!7��Rȶ�ɲ"O<�����/jLs�$ҝ\�jр"O
]x�癓\���B���1��a�"O�|����UV�
&�A4rԀ �"O������ ���b�d'ek6]�T"O@��Ǝ�ze"�8C�юdT@�"Oj�Z%j]�<��(�H��G)N��"OZ��'U�a
E؂ϡd�pir"Ov0��N�)e�Hx�A'�HpX`�c"On���hL�]6 @;Đ&��4��"O�%A�*&B,U@&�)6�n`P�"O��%%�+�b�����-���H�"OЩ�Q��,9��*�/ ?jp݊�"O�=B�gJP�4�R�"(�����"O��`᭛�d`
�����j����"O�xvH�,%{��z�NJ~��	�"O&�(S#�&T��`�£ծy�z�z�"O� ��ɗ�.H��q�ٵ`E�4�t"O�!�a�W(Lh�o�(�,�v"O�e�$,�
~��%n�;�D��"O.��d���-��<l����;�"O��SIM�R�Q(�F�.1(�"O�@��I�e�,\���ۮo"�pz�"O<-����6^r`��Kݭt�1�"O��$L��H�4�2"dGj��p"Oh���	��n���"%A �"OH��t�;���"�Lofdy"OX�����*y�b��й.l��b�"O��	T���;�l��ƨޡEh�"O����H�hs����e[8e)(1
V"O�xZA��QI\��Aŗ�~"� �"O��ӥyâ:�F�y��=��"O��kY08m"-x�i�$Թ�"Ov�RW���8(3"����&u� "O�����d*T��-��e�"O�����̘{��śIɫHA�0"O��y��UT'i������F�Q�"O�p��q������\�<p9"O\1P���iJ�r�H��R� ]��"O�P�@,ٰ0�#1G�3�5�e"O��CQ I$y5B��af�!:��2�"O�ɋ�/O�U�PB0��w��ɶ"O�����Ƚ ɓ6	�]���"O,�HU��DJ� ȁ,
DZ�"O��p�u�D���S�.Y� [3"Ox)�"�/+��<ڧ$�>Y���"O<��td��5�p��I-= �!�"O(���
N�%�^�-e�"O��BJ߹ib�b3�	�m^@�"Ot���3Sq��PgnR�,� =ZV"O�����(,��p�#GN[��jE"O�T��_|�E����1jt�b"O���T��8P,���֮Z >кV"OJ���	��c�:}�G�ڽB�4��"O��[bl�F�2.�>r��)��"O��9�mN�l\��kQ�A�6�XF"O�(RE�ى�xX�G�N���q�"Oj̘��)+BV��%9:I:q`"O���� \D�9K eF�t��A#7"O��E0F
��td#*� "OZ��H'a���i���j�^�A"O��aa�H~��0���-!� ��"O�Q����3V�ۢ��T�*�B�"OX�aV�e��DXDŜ�h�|�u"OL��%{����B���ڃ"O�YXVLfZ��*r��#��Z�"Oa9QK_�l����Mϣh�$*�"O^Ƈ�� �ƙ���A����"OR�ذA[������&PT&�@�"O��22H�9"�K,7@���"O>lY�� ����Q�(���"O��b����d���[���̦B�"O�Y#�؄N�@�S,.?����"OzD�o� �i����+�p]
"Ol�hᚕbR�h�(Z*a�>H�"O���`ݹ�b�*�#�Ba£"O����B�]��2���2~���r"Oz���F�hݜ���P^�~%�""OJ���Eɓm3���bn�!W�$��S"O
�j�D	&"$�v�7�|� "O��A	�@��!�ʃ4w��Au"O� B�(�[dUnɉ�)Ar椣'"O� NX�{�y�c�R�Ya�}�$"OA�*�	R@&�y�&ϒ;P�J�"O<��f�E����ve_�&?t��"O����H�ps~a �ިX1xL��"O͂��D-?Y���ۊ8x^p�"OrT��ۙt�l�B��m^ ���"O�"���2WmR�zɅz� �F"O�Xŕ�(X�з�;��С�"O�����;��As�$�2	�x`�d"O�8�0�O�'sVP�"�: �lB�"O���c�.|�D 0��8;D��F"O<��5-�|��h�˚s�l���"O��)�oJb=����g��$�\��P"O$��*A��|�wEb���Q�"Om�v킹O�ez�C��7�*D�3"O� ��]�]��a�%�]�Wv>8)"O�����ԏz�8�*�͹J��5"O��9dFR�6=X!("FF+W�i�F"O2`٦o��-��8¥��K�X�G"O�m��&�a߲���D�L��7"O�8��� $q֥��CT�Hڢ� �"O���`#ҐA�%� A�b�"O"�0�N �ݐ�B�͂�0�"O�}�E%�
L�j�j��r�a��"O�L��?nJ)q���"*h�B "O�Ra� <�������{��eJ�"O�����nx|�@��8�~źu"O�ӵ��}�|YC1@H�"E�"O�%�c��9~>ec���1�-r�"O�@8�'�w��z-�0[��m�4"O:@���I�Y�R����¤||�\;V"O6�2B͉Si>��B���^Sl��""O�$ib�E:f�ȼk�c�`Jl��"O�Q�q�ƉN�FL����5�4(�"O�[T M�EȖ=("��h(ܑ�3"O��b!�(2�b�k�((�%��"Oy�ȳ�
�ʣj�9��5�v"O���!AC����B
_�9�~��1"O�i�a�m���v
�,>�X��"O꤉�FRn�@�.D� .`r�"O��kS�R�2S��X2OW�fr(\�"O>�@o�"��m����h �u!�"Ovࡅ�E�j@�{���$aպx�T"O	�bNH7lm@�PT��$�,x"O�l��Z|wF`��"4f�*5�5"O�QR�K9x#��"��B2��#�"O|�A5��*���YTA���ħ\�!�$L�t�2=�pq��S�[U"���'~�q0�k��O6��b@`�\��@�'����W"0����'#K >���'�TC.?p�}�UB�3F 4��'پ��c�(�nQ�ЊH�*Cn���'�8�ە�F���q����.��iZ�'_(��.1o`$��n�$Rr��
�'��L�B�(L`��ݭN3Ԕ3�'�t�2��O|L��!L�����'���f�+W���e
7yJq��'ʆ(Z�a��?�Bm�&�x�\�P�'����0OI9*d�ec@X�^���'&����MX�P��Ӕ�7X��X�'-`Y��O�
���H ϑR����'QK�>ol%3ed0⊼(#ώD�<1��T<t�j��m�"�Z�<� �%@G��+.!80�m���å"O:�����`�PIX�39�򉊒"O��롣�\�����Y�Ft ���"OJ�"�5dV"�� �oQ "Od�R�/��P�և65`}z�"O� +��@4sRa�A�q��"O�p�Ag����eYV�Ueh^5��"Ox�	C��+�)�����4��"O^�He�$��R�M�V�2��"O�I���O/Pռ�R��U�@��"OK�7x�+ͅ�v�����%�>"?\C�Ii�t:�L
�~j����7<xB�IW֍x��;�I��"ͼ|��B�I,d�b ��+�=q�VM�1,I�~n�B䉨s��}k��	��x\c��S�_T~B䉬�Ք�ŵE��e�Q?Xp��Y�'NN�	G��]�`MQU�L���'���yg��}��9�g�FZ4{�'P�����KR��"P�H�DY��'x.H$#&M��9;���`��'a�	Cs,�7(;������w����':�UãѤn�����آt�<1�'f��� ��,���)liV�B�'8����Z��H@�$��Z�jA�'�� f�~X$ As�8W�ꜛ�'�y���"E�2d�glQ�w�~X��'��e5m��v�RyiשFztfa�
�')�dHî$Y���!�~:z���'pl䉱T�|4���`��,�$e��'m��j3$�2T���@�L� g���'rD��Efʼ9zB��!���*�{�'(!�jB�zJ��[���u���
�'�KO*RGt ّ	�#�r���i~�<��aC�,��5;w�8�l�:���R�<Y��
5cH�$�D�ıh�"M�6�g�<ф�Ӷ2��Q6t;؁#r��b�<�1LG��2�����#Bus�
�_�<�ժ�����G��Ok���@W_�<��I�|(�$��n4"D�Y�<ICMңrl��0�N�5��!�!R�<��K�^�R B!�3���a�KK�<�rȃ\�������1������D�<V
�1F�*$ �=�pa�7�F�<��3K��uCń216"UP�&�B�<I�	��v�y�`N.^k�1�ɋI�<9��ԏa���এ߃R�n�+w��B�<4F�#a[�Ik1Aƽ
׀��Ǧ�}�<I�+ȿJ��� �ǋ�`2, ����z�<� �_2 H�@���.`Q���AUu�<Ysd��Uʜ��C�� �+m�w�<��#��[U8��s�$#tt�6��v�<A���2_�������k�*���	�p�<��CR?p����&F�P�a (�o�<��ok�ˆ� g�6��l�<q�H�{�T���&��f��:7h�e�<9&U�@�����΀//�����`�<9�8V��1A�p�0�Q�+e�<�%���V�~�6�K�v��M��_�<ɒN'Lh��mݬk]��aG�[�<	�D��{�������&�v���AX�<Y�c�8M4(�� �$�4���'{�<1�� �GbM&��}50��E�a�<��W�`�T<S�Q?}rXb6��Z�<Q4'G�dV�� cI�#��]`
PS�<� ̀A'p� ���IE�I$����"OJH�l�rP^lIuj?���s"OМJ��$Rk��C�'&h}��"O @���wPp	�Ņ�n���"O��Y�J4�|�4s°"OV$ː�]<S�,IV�
�HVm��"O����I��L�{@d�+J����"O@���9�K�"	H�\�3"OZ�6��T�A���W9EʨЃ"O�$K��K�ef �i�M�XE�0T"O��	4�)�Vʖ�8��S"O��bo�p�ʌ�F��5�d���"O��'ݤ8��0��b�ڜQ�"Oh����N�J���T�iT|�"ODm���P�qe�h�&͟:����"O|¥��k3���f%\�g� ]��"O@ArN��4�飂�J�.�~�J6"OJq��ǁ�v>`�S*�	��E{�"On��c^�5k
 D*��9(&"Om)���D�Y����1IZ�ȳ "O��&e� Ӵ%�)�W�-��'���PQ�1Bu�ƃ�%&!�t�	�'����W���iM��^�� ���yOւ�\z��B�b�bt)�
U �yraC�K�ZŲƁC�r�>�(A	H��y�o�#	�zu@Il���#a���y"�(�8�:v���2LZ!1'�#�y�� (,�YqB� `<��&J��y��A)c܀qq����"-�B����y�c�]�A�ӂ@6<"vT�!���yb�	��ɧ�ڕG!���a�P��y��8i�,�S�E�PD�$�y��%J���cPL�*9��P#�Q#�yd��IG���e-K�KJ��A�o�1�y�T����B�L�H�^��2f��Pyb*�
�X�P��A��e�q�<���c���r�Ȣ �&��e�<Agl]z��!B��I	���(��c�<�2g�]�l��2���} �n�Z�<Qs�KQRv�����?9D�a��-P�<	6O�*Jq���X>d-�y�(K�<16* ��\9O��{�	+�DAF�<�E)�"]�����^�S����N�<�T$�1Q��󡁐�AN攊W��I�<�B�%-�ICU��pgd��Q�Al�<Ig�1g�{���Tv�k��e�<�ꏌ�6 �6��G����rDX}�<y�P�n�Y�SP�\=z�beFYq�<�c�t��QYM���d�@b�<1��R?>BT(bJ��M*q(C_�<���Q	z�(�r����:�	UHs�<����$e@������q/�����n�<�g�Q1`��(d��#*��� k�<مÂ����?,�e��~�<ad�7���KpJ@5�n���Sn�<�CN��rk�`"��B�!Qj��jm�<���T��ع�O1&��iD_i�<y�MB�k�!�֮�@�X�����f�<1U+��H|B��î�!!]�÷��^�<� ؈\y����Y�<YV�"2-8�	�U�eZr���ĝW�<q��)|��ӑ`�txBy�Fh�<y��-p���Sr¶��Dd�<�iO ��iq���>W,|�����G�<� ��j�R�#�>��S��Eو!�"O&��f'�nuB-� X�'�
���"O(�0�W�P�P(a�5� ��"Od嘳�ɺ%J�)�uI�wd�Qr6"O����15�n��<o/���"O���׸z��ؔ{�F� �;D�``���>5�91Jwo����#D���)�'���	�.1(4�4�/D��9$/Z�3a���a�	d���-D��u�)�:��	Ȗ[����1D���j���H����2�X�k�
0D��Ж��qq�EA`��Z�$��! "D� �%�� h���#���~7b�A"D����0a��P!"Ŋ<.HH�fE?D��Yw$�^�t�p,�'&n<�`'D�(£
҅H���K$��+�X����(D� �WG�E���qX$a6��
34D��j6-G:��H1�ԜDPƭ�6�6D��#��b\`A��E�\פY �+:D���C��3k�Dx�EN�h�ᶪ#D��2 ��"��eK���FcDtbb	 D� 3V��28���P����%8D��q�CY�2s|Ah��H��e�1'"D�P#f�Ѣ�WN09�Mjs�>D���J	m�,$�U(�K�p90��>D�<P�E�@A��3>_l}SC D� �R�[�eеH�+[�y�)�3k*D��a1掹x����g�%9!ے/)D���fh�D�R �pKٞ1 �t�1c$D��b#��3쬑rbW9\����
$D�����<�8����+�m��*$D�X��(P&�\�ӂ��g��P#U�#D��0`��1`xDkB���Ij�ȩV 7D� � �J:E�hV��,�����(^��y��P+s�$��]-dX�A���y��R�<�H	0cV5��|R$�T��y�a��6���+�+r�vh�R��yb�!F� )J�+� Y��Ua�y�Gs~U�'��%Zۄ������y¥ P,�Öˌ&�����/���y�5I�v8��� ��1�P*�=�y��-�K�*��(�Bm�7�K�y£�ft���!萊%�,m���Y��y���J&"M��΄����d��y�.B 4J��#Z�Z�������y¤�T/�m[�@�/��S��]��yb��7=�F�Q♚}<�L�SO_��y��&Y:�AG�Lub�Y;S��,�y�,I"=�qS`I,fv��K����y���1fAJ�#��_�e,�aS�m]��yrM��$�[�EV�8�aD�$�yr�� ��%��fרc�@�������y�gƨR�����N#Z � ��:�y�3t੓�� � ��
�y�B�,
6�9J�ƞ J؝�b���y¡:d�����E_�A�bY(�&�y� B��E2U�N�&T"��q����y¥��vh�qSʞ?�ƕр/�y҉�
:�$tMɸj�)���о�y��O*R��`�l�
^�����yB�O {|��@�T`��I���y���og�[����>L�fG�yB�!}�1;�HZ���]B��ޛ�y".܇�"2��s�R�Ç �y
� �mSJP�0�v���m�+��w"OT�ǊE
]�L�tGN0�*i�"O��i�A0�2T fKy��(&"O��r�m�,�QrƄW�t��m��"O�4h����Q>b��qɈ�_��d"OlP��+��U�A���OY�-�b"O�i��Ȑ�;�6�����/PS�4Y�"O���U����8�bf޶k?R9a"O��8�훎:�^�ˆ/�"��l:P"Oz$���(g���Q���Y��1r"O�ڕ�I�R�G�u�PC4"O,�۷��|�d�S�`y�	q"O�$u���Z�
5�A��3z�Ri�@"O�8�BAʬ,2�A�*��\�PTД"O8�$�N��@���Sp�І"O�d��LƬY��`l�D"�-�V"O ����ӌ�|�5냐[��HP"O<C�O��&��4�V�r`�0 '"Oj���A
�:�$�S�@�7j䜅��"OPp�%�-f1����/�u����"O��A5���T�kQN�Od�@�"OHx@�P�Dd� �U��j�]s"OT=(��Z��u�B"�20��"O��{���	�L8��KC�;�a'"O� �KO5p��E��T�~��"O�eyƆ	�9���Kv*I�5rĉj6"O�����Z\���$˅�\2��p"OlA��n�*M^��blB�?	���"O�=(�jY�y �� �[a�-� "O��I�ߒ�i3On�{"O�1�C��v6�'��.P@�ɒ"O�11f���}r�3ś:2@|=q�"OV��C'�=�p��'惖.�)w"OJ�W��'~D��37��V"�MCg"O��H��[�*����D�r��٣"O�!�A/�	}Fd)��Y#J�,<�S"O~i�$�Wm�0s�(]�
�P��'"O�AQ ��Y�a�S�A�f����c"OV ��ɝ�:0)�r��U��@�"O�@)�#'�*�GJ�=(L�f"O@LB��Y�6Ǫa5<)�6"Ox��g�m�Ѱ����#!��!w"O�5!��]��9��̅��	�"Ođ�
��g���	�C���� "O
�2b�P%�4���a_1S��`C"Ouc3��Dvr��'BT�"����`"O�EAgB�2QraS*[� 52�"O��ѣ��CM8 �P�i� X�p"O�4�b!����PGND !"O��B��_1j-Ex�)�l޽�yB�NlA��:��xs� �1K��y��Y$�"�H��[nH:Y��Y �y��YB���C�F4\��t ��
��y�  !�D����ψW9~a�'�[��y��Ѯ`�42P��X#`HI��Q�yR��e~p-�i�W�v��̕�yR��=$-h�����\HJ3lL$�yB����������.�C��U�y��"�[f�*�0${@�P/�yR�
	k�p��$!��99UFC7�yB�f'<�GE��v�����y�%��,�� �
����#LΊ�yR�K4^��p2NO�y��@�$��y�#L�R> �-� ʅ��+�y
� �2��	)&|R�NAZ���S"O��rK�sތY����o�0P`�"O>$�N)�̓FdUc�6Q`"O����"7Mӣ�	P�4�"O�	��kM:Vs\��D�p���"On�&���Nm��P0�L�H�yp�"O�c�
K����u���~eQ�"OF����\��T{����A�"Of�ӂ Ȱ	Ʉ�����!"O�jf�6`�$�k��1�r٢u"O6�9�+J	6�ً�d�Ka
h��"O�(%��N�n��q#ձxz��"O���`iUKa�qrtB�?u� �"O�(ۇ���w̚��� �����d"OV0�`�K���f�Y��(��.D�1Fb�};���w-ՎeS� ��8D�4��% l��g�H1Rx�B��6D��%OZ�:w\���Aft	C'D��`���G��u��e_�k,���U/*D���ID=d�MAW�I,� z�)D�XjPWyŜ�cΑLh%�#D�l8��7]�j��E�E�D^.9��-D�@��Tm
��h�D���'D��c�8	tlR�dG�o�Pp@Î+D��I�xA����`�=)�6��'D� �����YR$W`�9o�xCG%D��@` SvW�xd ��F�&D�$���[;`�&��s��g)؉�q�'D��� �+�ث�$6���R�$D��h��@ayr#�7�]��!D�H�c,��;���� ��)T)��<D� ���8.���OԈn4R�(d&;D���Ϛ#r}�����	)�Y�p/4D��3�G֛&��|��N��,�1�
1D�p��Bt����.^~��j/D���P���!����9��: *D�L��q��Z�\����'D�[C�+�,01��W��%@
>&!��޼��w`őQ�� ��o�$4!�$�m"`Z2jP�M�m"��#L!��Ɋ`���Á�'5j�аF���`�!�D>y�h1$ ը_b�	���X�!�$��:܊���li��@b�Qb;tB�	�FAHYy��S�N'� ��jO�4ުB��3�|�d�f�FX���̠4�|B�I~&�Z��/.��4p5���U�B�I�9!��p�`.5͘���u�C䉻qJ,ˀ�]	ly4��!�Z"u��C�	�H��Akr�5[: ��N��vC�	&���s���X-��0&4r
B�I=�8 c���C0BB�s��C�I!c|���t�уFi�$�A*v�C�	2ՊPx�ٌތ��^�.��C�!�V�� L
u�`X�)�&7�xC�Ʉ������"[��=c�*U6C�	C�| �a���U���"��C�ɑ9�zf%��:��< 2��8-p�'�Yh�'چ�v���i�2G]�h�'T2�+@���>@� �e�<I���C�'e���� �N�$1��%��<�t,��'F֙#��L�(n��iB۱6w�}��'����KVh��瓖32n���'>XE�m��Cv�ycK�z<��{�'�N	K6$Ў>���ӂϛ�\��L�
��� ��XA������:L}�"OtaTlÙ�M�"dB�iȠ8G"O�,�@㎱Gk:��"N�tI���"OisQ��<\Q&��2E%*���"Olyc�%X=_*����o
���"O&u����8s�vMX�b�3t�ȝ��"O�qB�$Z�i4���Ȋ�.]��"O���S�����L�-VDiC"Oj�#w ��A�t�Ҷ����2�s�"O�M����x|�BH$�!p"O�����-b�X�`�Ļ@�`��3"O���ھd���i���.��0��"O�i8��C�P�QC3�օ ��tZs"O�=I�)�*�h2aA�X(b�#"OP��C�&[�r���Y��S"O��	�)��q�x�R��DL2�!iW"O�+pM��\�u
��� B:���"Oh36�J�_��ԢĔ�46"=��"O(\�։ȹN�n�rMJ�N �]��"O�h"�Gu� �3)�+�X8�"O䈋�!1.��ƒ1���"O���a��x_H[KB4�p�@�"O�)%	�G�����X +в�H'"O���0S�>��#`�)�K�<��خU4$�"f߳4��H��{�<�v�Z�>=D��gM�8T������r�<�A �?	�DZqf�Y�PmP�c�<i�� o ��yf�ޙhBB��C�Z�<9�/B�	���C�mTcx�H�)W�<)�`�X@T�zT㒑:�dX@�D�h�<i3�/��t�I� ��Zj�<�vD	��Y2���<lx�Mi�<Q�k���p���ǗA��}	�cJK�<��Ț�(w�AKs D�LZ���fR�<�0�$e��	W��	g�LU� )Q�<��EH��bY.���Q��T�<��e�8�J0`�n�;>:�Y�M�<)Q�O�(��rv�8T]�8'~�<��d�*:������K�u eeDy�<9���~��1�	�4	'�H���Kl�<AeZ7XU���`#�- ����C_�<90f�I� /�=ުQ! ^�<�M�u_�ݩ�b�24m��Xs��`�<��A۠ �9Cc�-� `�RBU^�<a�#V�I޴���'\A�i�FϞX�<a�hɕ".(�4)����İX���ȓ[�n���@\>rz����N8�b��h�"���	=jP��㄰��ȓi�:���a!3LT��ܨP;D�ȓv{�YnQ�˾m9G���Єȓ:~섙"i��Z1)� ������P�h򍔹)ݨ=P4fB-Xхȓ+;!��J�#T,����U�A��>g���y�4�##��3�e�ȓi�v)!�/�0���$�f�L��+�\Y#"�� �kq�E�d��ȓz.��ˤ�a�jd��I�;{(���6dZ�SuF#P�8[�
�]z�Q��y�1f%��m���k��s����ȓ6�$��i$��J�a�?�^��ȓ�J8� �уv��т��>��u�ȓ[������IN<#ք�r�F��ȓI
�a@��׽x��x� WBђ8��:)�Q%"�4V l������t��S�? �����N)jN�3%/	�Q��"O: @�n��i&6R���ⶹ�v"OH�'��XH� ��#Y|�y0�"O�	2(�I�� �\Є���"O(����_ 5}��ұ�¨n�z=
v"OĘG��1���jV�A�,#"O<`�V�֪d~�a����v�ѩ�"O\�h�T�v8����u����"O�l[F���G� -�m�&"O�)�HA 1E4i���kX��"O�d�l@�#7:|�ނ^1��"O|['��x��ТC݅5)F|��"O4 �w�F��ĂN�	'd,�"O2�x%�/}t�|�aҸ0$�-s�"Ol�Kq&�$�dDŠ�!�pi3�"O��
7����ⅸ�I ���$"O�pK��F
XY��BG\�
�*�"O:-5�0�ȉ�ՂϔL�̀��"Ol��0.�8�z�3%��%�#�ژ�y�jO�#��5k4@QZ���oG��y��+%������h0��A��yr˝�-� �ٕi�9����y���
\�l8��JŃu� �*t�8�yÞ�(|�c�K�6�&i�R�"�y�R7"����-,��)�)�y��<�F�����'���f���y��A9oPl���* A&�Q��y�
�L�1�V�k����J�y����Kx��c�M���"7��y��P�C-�L����	D�вG¶�y�"] 3�@92���s$)V7�yb�E-Uk
�
u�׭9��A#�◒�yB-[i��8W�ѣ6�l�t����y�dU�F�a��ȕ�clTj�(ע�yB-�+|<�})E�o�xQ3��ڸ�y��%gT��`���4g.`I�d��yB
˅^���GG�k�8e����yr�؆������f��ieLY��y���D.][��ǣhT`L�!�Ǎ�yB�N�>��
\R��,��蜌�y¥\�U�
�����-3����yR�	�I������פ�9���4�yB����Fa1�=gR����G��y��	E�l��ЈH*_2�J`�K��y�ܺw	H��b�a"w�^9ڰC��$��鸃��(��"�ǐa�vC�I�(�e�w�������XC�I��`�b	�M@:-!i��|y�C�0|V�����I*�8�`H�#�B�ɰH�����,uH��Jҫ=^vB��-��)��N�
�2�C�fO�B䉡q|�İ��Xa3���׍�(nk�C�v�>ܒ��\��T�pn�9�C��Y���!gh��)fj,p���B�ID�F��?c,:�����;�tB�	 9������k��6�w`B�	!���)őJ�P0�s+�|LB�	�N\,�� ��gT�jQ�TRl�C��*S}Αy&�I2o��Pe�SC䉳R�D����ޕ`,J��d	� 7C��*J�~�IBK�#s�1�����C�I�V� x!�J�D���DͶlC��q�<�Hʷj�}��-�� �B�ɋ���H�O >�`��� �Qb�B�)� �-�F�Q�_g
���AѸ5��A "O�%<X)�X���ώH�����"O���$(��V�h°�)]�V1�a"O����>4��h��N�0���ؕ"OR@s�-�L�6�L�#�N�"O�4�d_Wr@2�I��q�Fd"�"O�	��t��*��X�=0t!"O����*G�C�H0M7b ��"O(� s�˔
���K��D�&���"O��I�H��Oq����MB�i�.��"Oz-��[E�H��������"O����h&$P��a)�l��x"�"O$s�Ա?x]�G�Bd�f"O�| ���",��tl��c%�yX$"ON�
��� 8��R�9}5�|��"O��k%��l�p��X�V��0HP"O�]B3�N�I�)���>��ħ�H�<qr(��D#֥�i�(y�^I	V�M�<��CKi��Q�ńsS>t�T#�m�<9/͙Fy,�3�
]��x5�m�<a���E��xٖ��bE�HX�/�r�<�C/��/�(:e�gr=4nVu�<I�%�?u���`� �m��K�
�Z�<�g�N4f���a*��;�]+CHL�<�gU�^h�U� LŖH�����'@E�<9�J��;� �ig�Fw8���gBK�<����%�R�(��*F�Ƅ�Bm�G�<	�a�����(v�S�c<�t���B�<�U+��)F0`��I�&���2��{�<12B^ʁ;@o��b��u�-T��Cv���sԸ( ��M7���!?D�複WB�
I�A�߯o�T����>D��F����8���&�*��sm>D�`j�	�'wE�Pi��2p�Nd�n(D�ܳA�#��yր�4G�B�ʶN'D����H�Fu�Ik����f���%D��@Q�ņ&�l12��U>(���#D��Ӥ�;�j)(Pc^�`���dI%D��[�ᓱu�*�ՇF�+ p�jgf"D��0��A�BL�����k4D�(p�ةa��q��/��t���/D�� b��;��m*7eB�3ug D�`@E�dpx�i-�z�*��Ȋ�!�$ҽ��l`0��?d���Ȗ�R+q�!����#@��,g�Tݣ�M�0u@!�P�1
:4Z�?�,<�%�F�!��4*�$��
+5���Q5j�7�!�."qB�TE��츢��҅'!�
x�4�Q��*w�t����Om!�d�,��y�T
9fB���H�GM!�
�����¸�Qb����!�5M�0B1ir�ܘ%o�B"O�� �K�N��������@Y�"O�pQ�E��H}@��ݑ(�V%�B"Oى��
/���@H��|93"OT�������yk�%J-���"OH�
��_�N^رt��|J�i�"O�u���t�ƔhA%Ո20��"O"e�`,D7[�~a�F�@I����"O�| �/^
�J�8�B�-,9n��W"O�P�N3+V�DەA�9V)�G"O�ɂ��L7rk��yqF�9/ju�"O��Q��nlh�e/úw)��3"Ot�k�N �u'7kH�� p"O� �̀��1?�B���(EP��"O���i�g���� C|q:�"O�hY�E�#����(
3̤A"O�zq�%~1$,�r0hr�"O�;5�^ :���A��ƪb�q#�"O��h�醦?Q�8��
0z�誅"O��e�Z�>L:���Y*#l�q�"O��;w� �)Z��T�C.z�
��"O�( d��8Y��J�,�Lo���"O\h�@"`]�L�!R�\\����"O�����6"nXk`��_��x"O�uY #�nV��
 ΃=�N�K1"Ot��v�\K慉сA>s��9�"O̼�B�� I�di�b@T	Ӗ�P�"O����l�'S�p� �U�D��T��"Ov%!��X9�lr ��@��lc"O�4@�"qa��h���zaYE"O��zr�B7s�t�r���*����"OR!a�e9m��Ր�i������0"Oh(څ��� q8�cK�!�T໓"OEZ�L�~^*X�v��<Дi1�"O�-K0NQ�=����g�.����"O�P`�.�$�i  �Ԥ@��hs�"O��RUJ�l��Q:u(��"O��'�Ef���[�o�XxM��"O���Q(��� M�#A^L��"O��f/m�:}z�+¡58�a�"O.�37̌.T��PS
G�:�"O�H��+͈a ݁�.�EHs"OR@xV��wt���M�[d�1�"OД��EѩB�Bѩ��
5Wd��"Oz� 5�\Y���%9b�e"OfV�J%��tX"G�~�Ԛ�"OPtq@�,VaTumH$?t��G"Oڭ���)~.���-W�	����7D�t�vjU�LzD@v�V�*�,yс1D�LPa������w@S�	Z�Tx.0D��B7Bi���"�M�������"D�����
#t�P�&h�*`ˤ� D�<���(���K��n8�q2 ,D�4�V����a�FǊ ��i�!J)D��"�C){7V� �C�Q��%D��x�J�I\8�Kӈ�$= ���#D�`"O�,���jZ[����T�,D�dQ��<+�����+ˆkߠ� �7D�(�pO�,^1�Tp��4dЉeh!D���D�\�v�PfH��D<|��<D��S'���%�Bjܧ	s��T*O��#����� GLV�gz)�"O��UHT,ʡ!�)�9y�yg"O�J�D�"	pTo]�=��"O6��CK�>c��H�c�5��+E"O��"���re�qAa�Pz"OZU�!���n=ܹ�R����̸"O�<��'$�#c��<�jL�"O�J�aQ+$�H-:d����|`�@"O�����8*,��C���*�*h�"O�y1��*�Q�B�\�JM2�J�"O	�5"T��z�/u�l�i#�
�y�;G/8myA�?|��T��!T;�y��1��p)�l�u�8��-�y��I{0@��zJ�AP�d:�y��׀zV��R��!!v��W/��y2����HfG�>h���G%�y
� |��K�L�l2�ڹ*D��	�"O@�S���}�d8�a�2_�nU1"O^�B n��5�R��P�+S"Ol�b�g�9���Q|��9@�"O2t�hŦa�y��́��V$�E"Op����"�L(תD�s3
|x�Wa�<���].W'p�	'�Y�~�yQ�Z�<)���8L���D���ԠFȟ{�<�B(��v\���  2F{�1�j�}�<�%�
:Y Q�J�>KF�A��Qc�<��c�0IAVDƣb!P1Sb-�Z�<` �}�д�q*���2��X�<q��Y�B���a��I�n��j�O�<i��\#��F$ëgU� ����G�<)F��H��%�@Γ[S�y��QD�<B�:[(m��)gL�8�wn�Z�<�VA΃ET�u�4(ΧM�\壆��p�<ĉ�}>8���-D�IĚq+���V�<	&���b��R�H��aK��O�<1p�ı/��i+�M�m(9��ĘK�<�凋�����
�3h´=��MXI�<���X�v�K��@9(�d�bT��D�<tnE��@���ۺx��Q�"��x�<���7&�7,:>�x�I�<qã�!w{P\��F�5R
l����K�<��N�H?Hz�O���KU�I|�<�щ߈@Q\H94�Y��0�Q�@�<���T��4¡�=0�)�c�<�`0t�����D��Cg�tx(�H�<���E����ʟ8B6�*�!Gl�<TEϢ�Z<�G���k+~�R��C�<QecT��Xi�@��v��m�"B�~�<Q��*� i��ڰ��F�R�<�f� "b��sq�M� �輘e�LM�<��[f������ՠi1�i�GeI�<�Sxz2e�
�~o`I�1DFD�<�!���vI��6�D!H�J�H�<y�-I*2��m���V�jiB�
�m�<ir���4#׭DW60�����h�<�E�Q 42 ���<�rГ�b�<��n��&μ��G����D��^�<�q�vz��2�dBp�uBFD�<�%@Ee(��7�F��5R�%�u�<qE�=�.�!�>��Q�Ğu�<�@I�oT���aй��)���p�<9�J�.���թβ-o:ih�j�V�<�u�_ z����Q�t�1D�M�<��AW*P�T�1ɔ�
~�x�IL�<Sb��|s��Q��:��u��"	r�<��៛Z��!����;J�X�go�<��蘧�:�`���Xy�Ix���<i���4L���r���k����a�<��O��;�4Q��j�:\X��C[�<���#������2�AT�LW�<���
�)�� hc�ɢiu�=a�V�<y�	m��TA��֌-�1C�T�<y@��pC� ��k�Z݀bl�R�<)�O�K�6����W�%��,�Z�ȓn�nU��E��P���݃J�,�ȓ_mh��$�Š!�ƽR6L��"��yc�G��7��A��ԼI��t�ȓ#=2	r�̒��-���ݿ<�Z���hFޅ��)��%�t)��
Q=+���ȓl�"��ݖ~��0��OU�B���S�? vlv钿	��D���z��P���i��Ip8��z��ĴCX�4r�iQ-��	��n+D�X`*��1zB�ԪI�����<D��{*<;s������b���rP��q�	JyJ~�Ο���b��aɓ sR���j6!�;�E�p�؁o��T���1ў���H�R��!��L�J��E ֫r�~ �"O|�	� �@��ը3oI->�F�"O��`B
�jV<����2�ҭ+�"O��J�FÆhv�	8$��5��m�"OX���,̟<>h�I�`$<c�f�'�2�*OX����N//�`$Hd �BEP�Pa"O\E񂡖����-~' ������HO哤h(�u1��M]�����	+TC�I�a�x�AHG+�y�qȐ.Q��������!*6f08�Ňt���ق�\��y0�n5�5a˙i��MxB��'?�z����<԰�P�B޼].N\hU��y���I�*����N+< ڴ��yҏq�ܩr�R�ALRe�����O��� HL�zAA3Q}�|;a�G7#�џ@D�$�K$n$P�4`�!<�50®�y�l��L�	"D7/T� ��'�p?�!�Ot8D�P�0%d�r�F����"O���ԇ5Vf���֒<�y[��	��ȟv��KeLt��b�5O4 ���� LO���Ԭ�;��ix S,���A��O��=E�$�T�	�eQ4��4���f��yB�B� �d���8�A����?�	�'wlL��C�+[J�A�$�9N
T�
�'a���f>d(r�(7�ް�Y�
�'!��3��u�P���͐7���2�'.`�Dy��46O�M��ʹa�Yc��W3���$�2|O,�tς?��\)�@G�a���Q��$��I&o��p��Y�T�IA�D)Ya���di���	� ����G>rS*�(�郬����hO�>���/
��U�'	B��6)v�,��v�<�O�����
��D��[� J�SJl����$OH�{M�(~I@�n�<uP�}�3�|��~��4�?A�ë}��H�@��i�I]u�IN��[�bNqP�Ij��8Φ�Ǐ<D��)�`�B^�r�E��I���*�*O`<PCK�k�v���@9.��E�x�)���N�Tp������|"AB2��B�ɫM"V�0�ᗧ4����i�$]jB�	��U�wK�9-W��BQB*&GH�0���'��!Y�<�1�H�tZب�n�+��C��%wX�	֋���Ɣ ����i��F{���O�ܰ)���R�S<2$	S	ד��������+?.@0���]]�Co#D�\0��R�xZ������3:���&l>O��=I�k_0\���(Q�X�?8�S`@��ў"~�ɿ`��@��f8'}T=�\�K.B��3ݒ��%@N6�!���?<Y C�@H�0��8k&��ʴ�Z��B�I=Uе�"��IĠה����'�i�<i�GT=��]�%�).q���|CH�X�)V6/�!�P/� c�݆ȓ5�
P�7���)�%8�	=*�=�ȓ	2B��R&�"6�椻@�ϟ\pՇ�PTC��"J��a3$��u�ȓdn8�t/M�][�ٰ3�J��ȓZ��I�І�!}-~P���t~H�ȓV���z��6:�XӢ��
,gE��S�? �I*�gC;e��A:��.Fo����"O�� b%��Sˬ���B�if���G"O����5m���ڃ�A:
PPxP���(}��#>7�tzF��-=N�$	�0jC�ɠF(�=C�l�2��5D!J�jL㞰��	&)$"A��œ�d<l���C���C��7$�R��� �N���OW/�C�	�D0^�r�;�<�����	Sf^B�	�b���Hb��><�K��`���"O4���^; ��\׈�>",���Iu�	B��T<���h�\��J���
�x�>Y
ד6���Ҫ� ʁ� a��
����'�4�J���J�P��P$��WF�%�c`2F��d�'�RP6|��~b�	j��G�q��@
:�� %e��I`T0E|���"oJ��E "ܔa�R'F&�f�S��$(�g?�W�ē+"�Q�(M9f�8k�k�G�'ўؕ'd��QS���4fBX�v]h�#��1��ɽ>��aZ��� =>�ƒ�#����/�I%[&�yQ-L�[��)�te��BUBB�ɳD���	�5���c��9W�B䉏x�D��oޱXB�3jG���C�	$�q3���.Hb`��١-��C�<g2�;��	%j���'0UH�>q��	޷B����4�v��@��˅B��O5"$�M� i���:`dy�"O01ctdR?�T��D7Bq� +"Ob�[Ǫ��id����8c>e
�i��]Dy���ih1�q�EI6�E�F�!��R�����^Ȅ����'�6������E��/�O��薢��(ӵ)�0)����'���'��2��3�ތ�dj[�(J���'�Ԉ�h^�t�MZci(6�D�ы�*�S�DI<���� �I/>n���W��y2 ïI�zT�C��"HUHŊ9�M�6�S��M�G	[�v�ۅ��&,1�GYH�<!a��LO\�[2�T"\��}z�kVC�M������Ï_�7�R�+B�Ȇa�fB�"OX9*Ě�}�4ye ������-,O|�س�	�z����Z�h�q�"O���S�%��y�wNFU��l'4�xYs���Ff��a�A*��D�6D�Jt
ڄ1���Q�#�=%L�(�'�1D�t!F�	T�1P#��+����*�	P���OOJ�(���n<*�X�]4M����=O�59���B�j���8��a��"O0���%��RwF�yb�V�e��8H�*OF�@�Ȇ�NDe���+&l���
�'�0�qޚ��Ri�)2^d�
�'��6K�1M��ؑ�)Ƕ/9\E!��D#�S��oʢjP���'"���������p>��K<�n�����Nَ��I�@�<��h��q�Ľ(�M��8J�pҥ�~�'�ynO�:�u��7I�}���	ިO�"w���y�L)7jX�N���g��$�pigoB�m���`7)���Bx��g7D�d:[9�(D���\00��0�E��y��ڭbϐ �/� -��	�Ճ�4�M���s����".��� F!YDJ�9OB�=E�$AA�l�u�E(D�,���)��?��'��u��n˓7;IP�(۽>�̩��'Ř-�
'L%���֋�6��	�'8D�3 �N?ZАf�#cr6�*�'OvyYd턒��P�u�]�)�2���� &|� ۧ��3�K+�i�"Ov������E�>���i��	�5 �"O:<pw�аZg+&��}Jg"O2�J��L��!�*V	+�Zi�<9slɓ~@fdREY"W�����Ap�<��.O�υS;3+���d�"��Ćȓ2E e9�'��"�$��kҳD��x��w/�,��2�8M�C�4N�4���s��򤛝4疉�BOӱ+S��ȓ2�$xѮ�1�5��'P0(ɤ���`rܠ���0��$��mB2	����?6|a�T!��h�歟�F8���ȓ[�n�1!Ij��m��A�h��zCf$bM5_�D�[!j��F\25��9�`4Q6�\�6e�⣞1uJ͇�(�
���xu��AC���C�	1��a�`J'�;sEΎ�B�ɒ]v���b�ԐT���7�V;O�B��
����2⋞��`�@+�uQpB��#�[v�"I\:�0'u}�	�'�s�2A���G�3G`�H�	�'��x�Ί.o�.$;'�����5�	�'�Ш��؈0�6�0.�� 	�'��`ƕ�t`��+<2,�	�'z���&��^]L��D�Ʋ�f���'��0	�7�:���G����'�ZS'c
-3��52���>@d$`�'	re(֣�gؤZ�fB0�,q�'؈����.lh��)0 ^���'�D��'�R�\��	jb`ۦ_�潓�'$�<8�-�!�����ԉ$�����'t�Z­Gzq���&�1��#
�'�B�:�	 I��H�%㊆qdl)�'��<�-O�^=�T`g��\�B����o�2:R-W/V�H1�m��	!�� 'z)<�q��\*����]^.!�&f ℉���<��iba�I!�T�L%`��&��^���PGH�=u!���ZȾ�ѷ�׋�V ���!���8�&P�}{@��b��
f!��Rm���El��|�	�s�\�!�͋���s���L��썁F�!�d8:O���o{,<pal��Uq!��?4	X�Q��8F2`ɶ�A�b!��H�H�2��%E�t �S�^j!�$��9.��[�H.�r�{���,FE!�d;`�H\:H(e�Z���(�Py�I hDșp/�pX�)�y�$�+�>�0�%Bse@���N��y�l�5:�Y�����;���Q����y�h�8E��,��"٣g7L�{���y2���k�=�wbB�X)\;d�A7�y�
�Z_,H��)	���҄Z7�y�J�6��5���.���D��y"��*=���Gϣ"x&���Ȫ�y�/�[�b��*�AmH`a㕝�y� ܍/��Y�s.[�Rr��3�O7�y�!L� �!�$�B	߁7~B�+
�'�b )ń�
;�ݺR�/�m�
�'�v�[&�ێ@C�|�
K4�
�'?8Ia���R!	HA��2bI�!R�'� �6��;�p����y�S�'�l��8%3����@�4��9 �'��țЯ¼:��C0J?,v��+�'�:X����4wjlS��B��b��� �̑vo�� �R���5�q�E"O�l���9$x��Ӥ��@8�|z"O�YiT��lcx�AÊ�@�eyg"O���֫�?��x6Á�[
��S�"O�qJc� S
 t.Y�Y���U
�y�K�" ���Y *�m���0����y�HT�QA]�Z8@������
�yOѧ$�8�ybI�:b|��w-@��y�g[�#|�s��ޠgt1W[�y�}0�TP���>j$D�
����<Y��+` !���Qx�H���	�!�����3 AŴK��[�j�[�'Jў�>��sl��(��r��	NF<�P�'!D�ܺd���N�C��B�7xAѓ�?��a��,��kN�c��I�q�0b7�|�d:4��9% 
���C�Y�5.�(�"F�v�<�eF69y�C �:m��A��ITx�|Ex���8�FM��OбjJP��l��yB���AII	;�H��q�"�䓻hOq����'LEgr��w��=����"O�ˠ��0a�V!��%��-a��"LO(�y4� w���f�W d�"O�����$��mK4�L5/�VB�"O�Ѱ�"KG���)��	��#�"O���kD�9��}�@�D�Z��"O�= ��8?͔x#A�U0����"OER�+M+T�04�$��4K)��AB"O�I1��[Z��K�|d��ӆ"O�2��<rZB�㑢�J�B�"O(���j[-"�a�!`ԡln���"O��8�l*.:k`M�X[0��"O�=�B�����@�2Q\Lda�"OZ!��K�:��	y挐"&D�\�"O,�ɰ�L%Yu$ 芀S6v�q�"OؼRD�`|ш�m�o-�,�"O.�ٗ��}�T�S�j��a�,0�"OP����$� �H$i�B�V�i�"OFU�'c���]{f
�>w�<xYR"O����A�M��B���`K~��"O��i2�ιpW!��|n
�A�"O����,�)R,3�
	=k�$�yf"O�:���9k�ʃ7��@�"O�!�&���{&�7B�P�9�"O���+P�(��֦�E~��Y�"O�+��#�x��;Y��1�"Of�xr�ͭ�080a�MB���"O&c�#J�$�d|���κ{%@ �"O ���c��A"��8t|�`�"OΔ���S� �u��!�Z�a�C"O���l�(1���ӄ�+%l\�#C"O0J� S�|�h������;�"O"�6�Ɖ'Ҭm��'xeE���@�<���ݽ/��Ԡr��"���Q�� I�<�D���dV�Ȃ�̦zmXDQ����<�1LP4�DH¹J��!Ny�<�F�I��ຐ���(1�A���	v�<�G��5�M���(Ӝ=*"f�r�<	g�)o��aC�	M��|��+�n�<)�J��� ڲ{>�ꥥNW�<��L zM�r󌅨r�-����Ga�U���Q�x�
qjDk]V�b���H(�R@C2&쬡f�
�M�<Ԅȓ������W� i��COԻ2�����$�vm0D��/��p��M
DO,���S�? ��D�,aB9r���/�(�"O`�W͖?�H�ð�FU����Q"O�25KQ����aB[y9��"O��(��cʤ��Oc��Q"O�l���4.��V�.t w"Oh�S��A�^ɠ���K���"O&�J�j�)A�� k� v@ }��"O�r僐-�nQ�#JK�{�1��"O��1�aNz�v͚2�Ϣq�X��"O61S�cҨ����6���E"O�Mb�Ɠ�i�f=��f���"O }Q�H��1p��#�|<� {r"O� � Hk�L�`!��c�Xh"OzX1lE�f�NX��T'O�TJ�>�te��O��m�L>��5���:�r��P� 0nRT$�o�o�<YEi�u����P�M�|���j�<!�
<k��裃�cnA��e<)�*��:�&A�/��#B�!!��'Z���/�E�P2
�/�,diw Odpz��4�F~r˻��t��3!:(��WП���Ǫ	.�&}�`G�F�F�84"Ol��3-��b�d���D�es]�F�O����%��=��h��3�b����i��8�����U�>0ļ�ǦV6Kl!��ɔ�����DǵO ��	5��?C�\�P(�.|NtT�4�J�RGr�c�?��?����s�(DJ5&�H�(0�Dt؞L�����S���ءp�{a~9�T�l�L	&�	��T�WfG�R|B��D[�A`���"�&�<�t��B��O.��,l~��H�3]�`
��0 ���Gӊy;2���T�����F& �z���4���@#�l��X�(.r!�B&:bM$�K[E�����׳>&j|���V%C&�|�5��?)�C�'���
/��W�4zvə��\�5b&$�"O
m�!�%��,C�T�������$O>�`���g^�h�/ݞu�\w9�����צ���� �4e�@�Z$<a2=k�,�O]���4��p=A��}1<ݓ�A� n�’�.��4Y��q�C�E��!�t�Ø(��:SŌ$V0$Aĩ[K�2��r�#0QQ� �q 2g�e!Sɔ�N�X�1@�<�ɧy������ ��q�n��O��]�G*L I�� 0��4���p�T�(v�ۗiA8���`�)ȈrJX	�
�FN���u�K1Ųyą��-Dt�`�ď�]q��P�l�BW^���dƈBI���5�ˈ1Ŵ)t�E	.Cv���r��Y�Q:NE��Ň�/}4�B�;�:e��f�b�sj�5_������,V%�{�J�=b�>E��k��u����xŖ��A��*L�d��㇎G�ƀ����C�n�P lF7T���[דZ  �����g���K��tSli����)`� (Ō�Zb�PpW�V����r&�PU� ����r^vY�q��.&R j��ȅ�*b͌*0~��8�f�=jz-a"ѱ K4,����mlF�Ƀ�W�*�	3��Ѫ;�`��Ǯ��p2��0����O׉�p>q'�\97Bx��F�l�&Ժ��	v�q�Ä%LaL����.=�:�8�A�:2Jt�\w��� �!
&�^�f���
Wf>b1��ޢQ5!��Gg�x��DJB^	�	pV�x�d�	�I�$\�%��bI$��G�G�f�|�����]��	�~�mZ<': ���Gc���G�I�lFr���Q3}�H��[�X��|�PN}���$gM�S�J�Y`O��J�� �ǁ͟Ky�d���yR.Дi��sㄑU�f�P�כŸ'����k�#p���cmџ+�����_��0W�
?5w���w��a~�[���(cg"t@�'uf��4U<���^�=���B'	?l\kE\#zP�ɺ��/*~r��S��4T=�S�YX�.իg�p�Ȕ�m�d�&6z%!��&�x�b.&(���kEE�:VB���+�d��:R^P�3E���Q��8���O>�eԤM08��U�fyzh8�KD؞�J�lϏvm���*Mb���p��J����U��>�0h*���,
��=�iZ�\�����'bD�9�OS1Q@��fI�$[�+��D9fL�	���0UP���	� S�a&�Vt ��N�w�$�3�A�$.h�Q�'��\��D����{Gb�3Hx�)JjM�`��J?t#�{d�[��H�����ϿsP�[jl�����kX��8W�e�<鴯��)Q0�CEl�pl���O�*T:��E�n�� c!Fj����.qOVqCl�"S�X�%�++ �� �'*��@�U63�Ȉ��J��舳�[.6�)%B	?�P�A	�9����	�5���f�5e�*���a(f��#>��FZ8ǄГ��$p4�����B��Q.ID�#eB�V�����x�<ɵ�
Lr��Rdߟ_��i��w?�C�!���T�˵jc���s%+�r��i���j|��BD@�8�����S�? tl:��ƺŊ؛Q��R0����$�R]h���4z�95��JJ���'���S�V�k��X!���Ԓ4��' ���#.���@2
��%���@�:�FIy��$��}���qt̒�%],	�Z��N���y�ډBL2A�A��!<d"��6�� �y	�}���U�W���@��Ũ�y�D�	Y���c5� ����-��y̉
I�,<��L�s�&��m�7�y2N	l��UJ��@S&�qH�yBd�%X��Y�+��C4�p����yr�I�$^>��'�[0��R���y2HےGS���q�ƛ-,"uspƒ#�y���	;��ڴ`H���W�ِ�y�T%q0���7��3	�p�F`[�y���q
���oӞZ:6�0����y/޲�*RW.Q,:���oF �y�fH�z�~�zva�":2E���\��y�/�/r֨��a�,O��<�@
�,�yb� ���h�"�	�� 9��ٲ�y�T�rD�e�
<�
Ia��F�y��B��aJA�ш|�����Q��yے�L�f��f��C���yB	"�� ��j֪؂B��y��aƸE��%�H8�hR���ybf.�h�7��+K�.}��.�%�y"ܑ^���t�9�t�8�Э�y�H�7
	<ԉ'���0�BuB#��y��Y8@D|��$NV�#^��ۑ��y�Ō�gSj����'�b��Pj
�y�KT nQD��a�:$Q�m�L��y��=�>0j�/á$E�h
� �5�y�D�)N�BI"�O�m^�"�X�y�"O51����*��}�)"��6�y�#�?Ux��T�ϡ0!"uq"����y��H/T��pi�!��JB��y�`+��iن�7v�n�@���y=O-��sn��a9|L20o^��y�ϗ�h�3���N�������y�%��u�>�[����S��	�6��yrFĺo�D�K�L`�)8���yri
ml�(�$%ң;+�%dU��y2n� �` �ŀ=<����,���yb��/Dt�mÐfG�g� ^��y�h[(F'�atMG�m�T��F ��y�mZ?;���n�f�ԄrJЍ�y2F#}�Rtk���Y~^����R
�yR'�Eшaɠ(��9x��J�E��yr(�=>�|�����2qz��fB<�yҮ�nw���a+ ���Bj]��yҪW|�.��+H
$�l(;��P��y����6�"�AV".N���E�J0�y��[� !�)��6%.�xp.+�yB�IL2$��GV�;M�hg�X��y�);����Y���SKҀ�yB#�[���6��r	<�J�����y2eEb�L�QC�;rL��/��yRB4aú���	(Y��`��Ƶ�y���#����ѺB�(I � .�y��U+x��k%�D ;��R܀��	�'�@pa�Ǟ�S��ंk�|���'�4���� �T-�Ӆ��b�p���'V��%C�7� ��BiO�_���'�d��&�ϯA��I8�+�+Ubnx�'�$IP�j�;mO�"�&K�PƨI���� ��{'��+ AqE*�,�"O8I��OM$}�D@����u��h�"O�F�+q�qq��XR"O*����Ŧ�Rxq���q�3"O,�!�kM���a�3+� ���"O"%�傈|�:T	��¦w��Д"OʡY�
��w�����_7����6"O���6�T�;���9� �).L����"O�����W��qu��1&��"O��JB�^�!��Iҳ��$��"OL�	�̅x����d�5^���"O*Y3t&�?{�1�jʀ��Q�"O���ũM�ʀ#�oӠ��(�"O���%\<I�b���5�� "O�$X6�F}	 |�%�.��Y0q"Or����<{6MH"�
s�� @!"O�EK7ΆlY���r���&���)�"Oz���O%8T�귋�>A���!�"O�X���=c�����Q�޼�u"O4a)��1�`��Y�V�l(�t"O<АR!��i���:S/A�ez���"O4 P��
�n}:���QlN�qP"O^�RE�"��85HEZ�
�H�"O�kń*�h�i�b)��`�"O���b� Uci���E���1"O�1àʧP����f��~Hr��$"O�*'&ιD �0K��O�$6XP�"O�XB�O	Cr�x[E&� d"OL"�F�Q&4�	�$C�[X����"O�LY�%\�G �X; ��� 1$�Q"O,Hi�=�X�0P�]"��(�"OpHp��,"���Uf9@L(Y"O�� ��V�/�F�#1c�:jM����"O��z��P�L��;S:D�HU"O��1 .ڦF�^�0�`M<12((�"Ox����6Ng�9:nǵ''�tç"OҰ�2��[�T#t��>�,BV"OLy���M!P%�q��Q�@0"O\BEnԉ,
.[�A�(z�\V"O�(�����D;fi��/��A� "ON|�����Z�A(U�p��1W"O����F�%�<���K�1~�0�Q"O��:2�Wk�;T�B|�¥"O����$*|��H�+�E8��"OHeH:x����CI$�"O���b◄E�yb�GL6P���"O4ɓ� �i�e�L0'#~�Sj�<�t�CW��gH4K�=���WI�<I�B�h`d,1bL�5U ���&��<	�Q9h\�)T1o�M�ס�a�<�1F�)��$5�ES��b�<9�"�$,bfb���Ҙa��Z�<�C8}��Q��o�xؖ���[�<�f�Ee�-��Y,�H�F��Q�<y�%��:�|���%	�m���lA�<QpE̫'	F@��Nf.��vE[|�<�����9��M�JU�8R�"e�<aFւYa�Y���
ci���LH�<���D���Aėt��)GE�<)!`�&�U0"H?c���
 @�<Ĕ0u��l��A ;?-����BA�<a��Pe|��7��*(֦���}�<�h�]��B�E	�C���� G
{�<i���u�>)��!��4��S�~�<� ��cѯ9~d\�w��3,�,��!"O5��,5Ό��'�����"OܤӧGV28�\p1��'s��p�"O<uڅōT�����@+&���X�"O2�Y�

�j����;%���#"O��%�d� ]2�f�:pG 4hT"O+���}���/JD�B����Vq�<���(
P��*�V�18!-�e�<��哤)i��1*��!",Ap�c�<I �A��am���k^_�<� �0�D��G�.tծR_�<��l�9��Ჰ
��U�
�s�<�4�	i+d���&M�i����̊a�<�b����a:/�=@�J�A�]_�<1d(ҟK�X)ˣ�
95�$Q����X�<����-�����KISN���F�U�<��N�nh��
$�Z�"��'�L�<I�7A;�ـׯ�*a׮���!�C�<�"�ȯI\0��[�n]�;��V�<q$�_ ���
��"��ѳb�V�<��d[�0\l	��!Z�Z��AcF_P�<I&N������Z�0S��E�<	CCU�+�
$�d���]&��IN�<I(O�k����"o`đ��P�<���H7F����7���yFd�T�<Y���0-�\�猔�6 2i�V�<�P˔�Vy�Ԡ��V�F�9A���Q�<�)Ar��a��#	8�&}�"�MN�<	���Y�HAB!�@ 9$����g�<�U�UMP�@��J�e����I�c�<)�b�`��EZ�?p(�TJ�[?I0+T���>Q��	U�t��	�	��-�W�ZQ��H��L~���	�9 ���c��|B��z��� ;o�C�I7 ���	�ː�Y��ҥ*�#|�c��"W%��h׎(G������^�js�݀���J���yR۸SLZ��p?}�|$Ⴋ	!_��CuDEk�ɉ�H��	�3�N8(��E������� �PB�!�BYkâB�X���x�I�<,6-��nbNxXf�7�Ox��c���$Kbk�t0<0JW�'Jb�7�F�D�����(,\��/ңH4� {�D�0�!�KuT � �Ӻ0�xd(Xy�Oqa�{w*�~J�UC��EA7�[8) �+��@^�<�`N�(ͪ�Pd�@9D�5kS�U0��XӢ,:�ĕq���D�cؑ��ۿ81�lCĊU6�!��Q��yK��U�L�8hih�7���R�lâ�R��'�8��3L� zl����=A�i��~���+��F?!��X�B�pJ�a�=ظ�!��Ij�<�6 �&��0���,�`�Y�EK_�'X������ݜ��d�`�jY[��΅	2pB�	cA�Ls���;vaF�%-�z�tB�I�R�BS��/L�@irß�UzB�I�\nT� ��i���#�\"g�rC�I�n�����!<K�!"oڡf"XC�I�|_�$`���`�j��Z	�~B�Ig:\ب�H�<�|$DNL�WM�C�I�9Шa�gG�
�&,�4囬P�!��K�N�<d*��p]I�';D�!��\;�J�CӤ$n5t��Gѣ-�!�/Q2Px���)U/��#�FI3�!�D��2�=Z�"9M���`�b��O�!�<���cD+�-�n��#Ӄ�!�DG ����Ł�qC-ᓢ��!�;?�����D۲�&�!�-��"t�,�,��H+�!�� b0ce�Fp�5�6���j�#�"OX�Z�kĊ&��d��B�X.jq؃"O.|�m�а�l��P�r9��"O�H��┷},�I
�+��S��"O����N�>V�1�$jC�"��q�P"O*<xwm�+i�����^��P��"O�9z -)� $����0K�̼(G"O�QpD��1�����\,�>�m*D���DGS&��	J�F�t]Sp�!D���`��m�r`jv/�q��E�� 3D�H�cN	XD=p�-�*�m0 .D���Ҩ"+zٛw� 8�N���-D�l�ޞ7p���k-\Dy�v((D������V
"m�/h�v��S�)D��r��ҫL�p�y�I�+��6'%D�x7.¶H�(əU�ǫ2�B!D�(;Wa��p-��h�E#�t�/?D��aҬ^����	�T"�퉧/<D����P0qU�(1��1�:D����-�VL ��"?4�ע;D�	�!�7c�~�i�J� ���#�**D��#����,+j@0��F�3ڈ�$c*D���w%ʤ6������g~���C�-D���TiJ$���`N�!�� ��<D��{�j�B��R��ߡT���i;D�0�g�@: ���� ^���1b$D�8c����}^���Qaѕ#%b�"�/"D�ЖÑ�/�����HX�1N7D��*`%J�;+��pbj��(���4D�(��B%$�^�q �G��};Ќ5D�|����~�f	YQE��8Y�eh0D��Y�$R�!Nn�jA$ЈV�q��0D��h�A$/���E��D����7�,D�Ly�K?#�<%@"N)X��_a!�d�H�b�RB�8!(�i(b�;$I!�d΢^0M0���W���x%�
5!�D�)��<���»W� �;��\���$ʠ>��1��kp(��G��y2��F�FY�墓_�@ࠤ)Ď�y�W�&�L��'�Y P���W�yB픣'�(2�8[*<���Y��yiS�&�ָcPe�<&��±U �MC����w��	a�rhKݴwV���m	"*x	�c	�{�8�pw�Ig8�,��f��m	*�Q!�N�D6�0�&h$D���
5)zU���?/����)�y�^,NŘ�2/<�tz��=�y�n?��p�="�"<���y�h�9H�dX�n^��<��@��/��O���OO�Ep@�δ��0� f�������3ʓ�����@c��C�<�pWŃUrO*y���ɐ�}8����E�n�4��������8\-Q�"}���v����%�Z�vU���O��Ѯ6�S�OӬu���K� %��2�EJ�B.]�'�:��%�a�$	�S�@4⒅��Vuj��p엽�?9u*�.X�lbE�O�ћ�B���?��F ��Xٺ�(T�R�rjl�Mw��^%V� ��?��t�N1$l�b��Vڡ+g��$a�@;�S�O�	���\#YF�L���am��0۴a���<E�tgP�jܤ�����%*��-vQ�\�
ç;^��P�j�������U�F<�>y�1���ɣs����F�HJ��� � ��O.Ọ}�I��0���E=HK~�;!G�3=RC�	q>��	U��Tr��DG�w�dB�I�o�>h�V�:{�x�kfƏ�.�B䉆,p�pUEU�#m
9jo�`�B�5�.�*Rƚ�^�+eEL��R��d=�� �ڷ�ǐGr�j!ݶX�l�C	_*}Z~��V�i���v�*��I�����
���"H1`�R�KR�y��Z(v*P�x��� t�T Y����y҅�
d�(�i��ޛj�����0�y�$�R���1aY,q��ر�h�#�y"�[%3�Q��d�2j��P�#��yR�Ʌo%rm@eECe 쨻�D�y�*�-hAz$��0a>`-�D��y"��$ft���dO�L�jŹ�&�$�y��N�*��}d�^�?�h1�V���y�I\�%^�y���8�L��%�!�y⏏.r��tgA�nHäKN��yB+��w��ͮp�4ف�h٥(xy�ȓU/
��tl�%T8;T�ݡA�$��ȓ:D��CnS4����	?�6}�ȓGt�|S�e���5�[�O8���{!�t1��Ǵ*� �ҧ�� 7`���^f��G�KBiʗ Om�(�ȓ��=��R�-�E
�H�MWޱ��py�E���Z�t���#�A��8	�ݨ�恡1΀�Ɗ�
n!֜��?�d�83��8v�l��W->#�VT�ȓQ�Ls&��/&�\��@�Y�&�ȓ=�\���J
�j��FX�=�ȓMip�6)��\�bu�[�q�ȓW(#S͛�삱��?J�.P��4��|�e�՘&���ԇ=~�f��ȓ/D� %M�J��q���@7s���ȓ.�!#$��,NA�@��
pȅȓ}��xS��8\���Y�	�p�ȓy��<�gD�.�ҡ�1�Ǽ	x���~y�{FB�:���!b�:t�݄ȓ'����A�$%	�K���ff|�ȓ/��iVU�3؄r��;E��Y��_z���!��R~���r�C�\���zN��u/BTd0��)2��R�$��k�-L~�z�ƁE|็�H��Y�r�G:��kU�:/�������JEa  !�	P!
�E��a���5Z�e� j�hD6wZ��`ڤ�����H����e�nu䡆ȓR��)bא���-(S}�0���A�H�/P��(�R�$_�܅ȓZ�h����8��\2�E�Z$�H��>����� ؚHb�V�G$m�ȓ+F�� ���.P��`r��.;��R�2�a��7dkD"C�ʢ�T���F��9J�KT�i���9��˸<�C�/��p#�Ĕ(Ӭ4��:s��B��:Q��C9W�M؂�]0XG�B�I�*g2E̙�%:1=��MqPG,D��k����G�F��DmMcR�H��+D���Ti��X�V4�ą%)��D�+D��Sp$��p��5���ӹY��*�+5D�t�pbAL��[�g�����1D�x�b�W�KN� L���x,J��+D�칖���3UH��4���L�e���+D���q�K�>Z���
��
y���+D�����w�1hBi�ZT����%D�L����jh�8;�剃E��l�ì%D�p��Js� Kg�	�%�Ģs!�$\�%c���H�} 0�XBNO�Y!�
�$0��cת�{ᖍ�/K!�DܫZ�E"4C�y|m2 �Љ|O!�� �*R/?,�8�.�W��p��"O��QW�C�	�xd���c��yP5"O��� L��dQX��1��Ic"O��:ƨ	�zq�h�!�$M'h�<���[�p50�U��C(�<)�ت)n(�E��2�w�<�F*/�T��S���0j|���q�<�%�B�0TaEI��M�����p�<��o��]�����D�I��1���C�<���\6��@�����'�HV�<�aBq,}��)c�R��&K�<1��M~4���SAZ�j_���s!�K�<i��ɗ(�:ٳfu��@1��C�<-��Ũ7�KF�t��u�1�*��ȓN@�;��I��`���(�9��H�0Q�`�\� �H!�^s<��ȓ{+��:���_v��P��|[0��	��Eh�i3m��y7ǜ��8��X��!�`%Ob���Qf�m����j��[�a �a����w�T0���t��\S��% 4[ ���'��8�ȓP���,�	��d���Q�����}2���U?[��7fW�����ȓ6̋�l��J_ t1#mJ�~�X�ȓ	G�ɓģK��u�B8 6����j0���K!-#���o�$�ȓO[8��U �{8��a�
pr���ȓ"�,���E� ���î���g���GM`�&��í@(F�h�ȓ0�l �q�[�7�P
%� s����\�<E[��M�8�^P�Sd�~��P��H��h;��G�!�x� ,@B�~��IC��O�+��|��%�Aw�u�ȓ^�Wd�3}S�@�e����u�<	���g���"�= v�12!�d^����J!�k�*,�L܊{�!�L�y!�L�c�Z�p���f�[�8�!� (���LIF2b�C&��!�;%7rY+�g� �-9F�ޟ�!��19T��
,i��&k�:z�!�ɣX��A*�)�.0����#�W|!��9��-z�ã	�
���޹h}!�D�:
���FJ�.�~L{��^a!�G��"�ABIHuN�c�LO!�$E�@ց�uV��iK��DC!�D�?y�"m��E�Ef�`���^
2!�D��^E��:����p|t���M*E!�D̓cu����I/%�ɸ
P R!�Q������%���`6I��5W!�d	%'zBhz�G\-z��`�� PP!�d�b�F�x�h�C-����)m!��R��=Yr�Y6�yv��.R!�D	Q�ph(� G�X�B}��$�!�$�*%�8b3j�}r䝒�*�`�!���0Mu�`�z
z��F�0 �!��&Y��TML�@��e�A~V!����hp��!Z� 1'�� Q!�D��p��ԃ�&W<4�,�!�#Y0!���&y�(�a��5�1�LR<!򄏕��A��@	�T�@�ppe��
;!�d�	G��$��������B)!��<�&�Af�
b��:��!�dǮBZ�Tp���'O�j|�$H�!�$G�t�ڸ襪��8��rh*7!!��  �@uE�(��aS
3\�x��W"OsK�)X�`T�!!�(��"O�p3#l`-F�I�Rr���"O�t����$��L�b�n
j��4"O���D 3�����>o
X�v"OT��pL"{�d����$Z�l"Opa2��;�ڔ'A��uR Y�"OM�3�+<�dy� #�48D�8��"O�u��DѸKr�z��р%��""O�Hq-шe�
�D.�&@r�I��"O <��M��,H�<q��H��$/�SⓂ�r��5�I��4ْ.=JgC䉧��9�F��O�  t�C���B��z�
}x�ɗD����NC�+�nB� E!�	�7�����d��@ 5��C䉵!�6����L (��0��_;PHC�7ql��C�R8Ȩ; � LnC�1���pwm�!��\:��Z�m��C�9��� �T�tyǚ%<\|C䉶bj�&��&|�a�Pb�"˜B�I�:*`�3��)�����B��B�	�]��� +G�B�ܐ�lۤQ� C�I�)��Yhpɛ�G���d��>|:.C�	!XeV����5h��Q��n~C�	�3D&!Z�$ԲYw�Ic�G�r��B�ɮSkx��nŲ7�|h�E˂�rB�I��v�[��Өg(�;���9hC�I�0M"��������\<j�B��X8�ۏ"�H�{�.���ZB��\�&D˷�3:t������C�	�a�ڕQ�${��)�#ܒKB�C��4'�H���k�;}=�ɨ�[�.`�C���V9)!#S�P?���aN�P�B�	�v
�,��G�R��yd
=PB䉁��u�S��U���"J�4m��C�Ida����R�=_��9#`�c�B�I$
JxPT�EVN��ׂʺ0�dB�ɜ����v�G7T2���kS�,�8B�ɎƔ�H#DΉk[�l�r��6y�B�	�2r��c! (@�h��ѾkB�	�<��0J��e�N�K���%��C䉣x�X!�FM�:>Z�`����+H�B䉶`��sԍ<�vX8�f�hB�	�/��� MC
�8���D�v�RB�I4�<8��ǈ>�0�"JC�/&B�	�s��%�Ц�n?b�(F/�38F�C�ɜNI@5�A<{�͕h�nC�I�v���sp�ۢ���q6ʓ�KB�,'��ı�D"�`y꒸"C䉖 �"��*2~ ��d�O��^C�I*~R����	[�"�PՄL�Cq&C䉓4"|� .m��(�Fo��p�C䉤,_��ك�����QfR�^C��6k=��P�BΗw�~u�B�ϯ9�FB�	.�0л�B�=@�["��$B<B�		dR�:�!D/T���[@!$_)�C�ɹs2� �?(�x�Bb�_5�C�"\�"�h K��/�~pC�Ģ?��C�	8F.0��I�V�x����;��C䉚�ZlpB� M2�m�$`�C�I"Q�T��+��4Hէ^%�C��'���#K�(�J����C�I��t�� 暡;ΰ$sr�!O��C䉅w�LcЫمj�t��l���C�)� �����|��@h#h�-y�.[@"O��4�ωv�,��cML�x�@�3"O؍yUȐu8�Y�->l�$��"O �0���tbH�ˉ<f��}ɢ"Ofh�hZ5$8�Y3g��@āX�"O�b�.M^H�p'�
<
�P�d"O���w   �d�vq#2a�`GJ��f�Ђ(�!�$�"��H'�\'i=:�LӀ=�!�@�8���q6�ҏcD~A���E!��5�~�+#&� 6'j��	K!�d)M�&�abO�Ej|�֧�4Y�!�	�+��!�� �(j���rE�"m�!�D�/��1�ʀe���{�C�3m"!򤇶�0] o׷i�43���(!�� }@�G��HBi�&���"O�-A�
<*�����0.�� e"O\�pꀱ/u�a�b���ڀ�"O`�aE_�v5��p�bT2"Ol����&0��3_���Y�"Ol-S���
Ӡ����7)R�!�f"O�QJ&LJK�8[�D	�g�ư#"O��p%/T:�b��G�Dۘ}*�"Oؠӭ���l�[4�B1d�X�5"ON2�DAu��pĆ�]F�5�D"O�ɕ�zs^ةuEW�jT�;�"O�D"���S�0�u�H6�S�"O���@D�L�8�&㊸h	TĹS"O(y��	˙[��-P����b"Ov5�q*8^O�s�l���
�"O��C[�9�9!B�S��T��U"O`���O�DA��.�r���Y�"Ov��#O�#Y3�尶�R�lW&�b6"O2EJ�"�9	O�Uˇ����C"OBQ*�Ɓ �� * LɦF��e"OV �C�H�ul�	�1�,C�E�D"OBDcìY_��P�l6#x8�0"O�4c)��dBѠ+��	��Z�"O"i{W�X$�z|Y�ɒ�J�$�S"Od��7��^�8� giK�<	��s�"O@�"ch*.��Df�!ڄ0"O��o�67HɃ�呴j����"OD�0j�:�RP_��h9"O�����ƒ|�6��ģ)j12r"Ore�ϊK�ԓ#��2��@"OެK�\��:TE�|���"O�R�# + H��d�-ּ�k�"Ox���$.����C�#��"O�����6��v� 1��#"O��6 ,�0��.����U"O:�
���O^��`(�wG�\�u"O��o��6�TA�S�ܠl8��h"O�z�MI�d�*2�X!��:�"O�)) ���vOJܩЉ(��	Yq"O�%�E n� (+���C���@""O��VO\?�@��RǛ�Zd�"O�)Ą�3F�x�@P r֘��"O~M�p)Z.T���PÆ��gx^��2"OP�"Sk�2�C�Os��{""O��pc��w&z��3I�o�B��"O�P1&Z+&~h�#q�F�� �"O�$[����<���I��G�e)�$j3"O�}s�I@��Z�FF$I \�P""O��*�a^�R�4�c�5K	<�i�"O`�ƒ�v��sg�L.Q���B"O�\���� _������d�D��"O�8��E�6O$�h&�V�3�a�"O�a(�.�W%`�B�g΁y����"O�yS�g��W�UQuA��+��̹f"O�x!"�_� �]�F�W}��5u"O���I	1rr�ICB�^�Lnn4��"O81ɤ�T%ؑ��
O�@�"O��p�N�7X�t�C���O�ڭ��"O ir#M��̅S �T�y��$"O���#�9C����ݕ,��!�"O��Cv�]jGF\���B:@S\��"O
�)gؗM�@�����2OX�B�"O�P�稈c'l�sC�U�3�� ` "Oz��V�.7�p����O�����"O� ~��ʘ�'L� `��+�TI4"O&1+#Nf��	_>8=X1a�"Oh�rflR�Z�aj	%,;䁒"O�Q"����� z��%!&��c"Ov��R�4|z	1�4Yp1"O�!��b�qC�@H)�e"O
���ᄒ_'�<���J%"O>���$� ��a1A[�A����"O�T��]�@T0�� �&1��]��"O�)r�e3���FE�R����U"O`�P�+O7-t���Dܝ/�`Q!b"O<�Ί�{�E�Ҥ�.&��hX�"O�4`� �YG&�˱�B3J�I{�"O~x0 ��Nj��6nǵf���&"OL8I��Q%�>)RQkΟ=����"O�(�C8~h��S�	�.|�f8�V"O��{�#�
b�t��BÞe3�x�"O��{Cg�-������}zx��"O(�I�J�,	����J�&?]�qe"O�q{6G��p�bdȅ]�H�[F"O���.ߤpҎ12a��`�,���"O�"�7S���CD'=��q��"O4�Y��i3Q�M�"�M����$�ybC�$ V���h�C��
q��9�y��ӂLPʑ�,� �i!p'I��y�Ĉn.� �Pe�e��1B����y��nKN���E�e�hD�/��y�EYi�4eiчƌ%X�A��
:�y2��%+���ꍳW��|��e@��yR�̩>ݖ��FaX'ezaa�:�y��H 7������v�,�Z5L���y"�9A�yt�$ R|����ϱ�yş���%��0H�HX[�W��y�E�o�,��S�J-G�&AX)Ī�y� �J�X	q7�
 P��9�1�%�y�0;j��jU��;@��4�����y�cb!��ӕ�H>2R$"n%�yb't��DB+��1I���y2�d�lQB`��qz�!�a����y2��R����3;d�"oʔ�yªX
I��R�E�1���0d-�yr��%�j=ٗ�K�1�N
qlH�y�iI�_�h�Vl	4`�(�l��yr#�qmv��",(�L*�U;�yr��##kn@����\���$�yRN�O>�"T���.�FTA�C��yf��Q�6���+Ӊ&����t*�	�yr#߹t0X���^�9�=�qπ��y�HG�,��(P�D�LT2��	&�y�b�$p`d8Tj;K-�����7�y�뛶'@�1e��u�6Ԛ0+Ņ�y��LC:�5��[eC�!JufM��y�d$_�,`�ں^�0�����y��^�p����3]�$Ђd���y҇Q;�j�eʳk�6�$���ybi@�E�<��U0oF
�����y��/���!�ͩ��ظI\��y"'� ^��p���
=���M��y�i��D*p��H�;
%à���y��� u�f�ZP�]�r��c��ӧ�y+�3	�1��!�#�0�ҡ��
�y򤈀1J�B" ߡyx���!��y��\�v����o�
sA�AJi�y�>7�]����q�4ۄA��y
� ���.�Psp�ۃ�n� �"OB)�P,W�@dX�I���0�4"Oԝ2Gh@�x�!�s.�/A����"O��S�C�1f�QAgE 8�fS4"OV��5-]�b�8�2P,��+��"ON���.� �$���k8s�t��"OV���ת?��3�+��N�И��"ON�c.ǔ3��)��)0ʺ��E"O��d
nq�]�u�ӥG� 䚐"Ohqq�L�?����'G�o���Q�"OEɍ ؈�I�D�2���9%"O�@��K�^{D�Jǚg���"O4���� A���S��4&�б�"O�Q��V4#~԰� <2~��0�"O<9@��I�?�N�b�c�Y{��i"O��2��+z�`��A�5z��"O���	�&c�a	��ߌcp%x3"O��#�-KՒL��� �p51D"O�Eh1h��}}(����Q?�E8�"O>��΄]��A�/	 c�Q�"O|�&��o�:,�u.�S
̄�"Oԥb��ً]���ǘ�a�@)`"Op��r�Y  �NE:��A�{�t���"O�U�V`.N��a��#
����"Ov�zE`O�Z�#P�V9��"O,C�BK�蒱*���� �p= �"O�8�΁:���5 \�K���)A"O������Z"��3eޏ&��$�B"O&-(��5?�0�H��ԚtA��9"ON����V� w����'@�X���{�"O�q8C��v��i���$�`��P"O�L1J�4L��X���J���"O�p��H墔I�*y�P`�"O�P�a!�p���H1+t�z9��"O�`K�+ίj>���G�Y�L��"O�A��V��2����0�Ҩ�2"O��4�E�N����JC����"O0M�����qt]0	N�K_�""OXh1��3	��� 2�S�yPVae"O��B��� k�A��Ѵz����2"O��[�&?��!R�J�i�fT�"O"h�Qe�=��Ȩ��	�N��1Z3"O@�"ѥ�"��$�G��5	g~l��"O�K#��3R䚵K^29�>L��"OV��W��:�<1F��;G��S"O�	�6,Evh���ݪ�:�"O������ig|ر%-55��C"O�}��*Ȳ0<�ܰN���� q"O�8��n�Q�|	��앒ev��"Of�f��r1fx�pXH��y�	T{�-k���g��ຕ	��y�oB�O�pŘ�F��bb�0��I��y�$
�Ԑ��G6aeB���Sn�<)#��	(+z`BP��-��TZ�<�g"Sgu�tx��@&c|d�"&�]�<�d��@q��+U/�aۆ]k���\�<3�4q�$ ��nN"A8n	{�D\�<����-bLB�FJ��Qk�^�<�l[3Ҡ0G@ L�I֢WE�<���04��di�L�bO�%�`JKm�<��ٕe8�Y �{��1#�h�C�<IG�G�Y��"�Õ�0jk]�B�	�H�� ��=�"�J�+�/n�B�4 W��F�.�8�N��{d�B�)� T�S0�ʞY�|dZE��,�$��"O�I���W0 >�@ʤdͳ|_�1�@"OҼ����UQ����ϠH�U�u"Ol\(��P�z��� ��ѱ"ObF�IK��xWDO�+*���"O����Ҽ`]~lCc�]���"O�(0����c�pU�Sc�:����"Ob ���&X�t�`Ҭ0���kR"O|�[A픹*����/W�	`�`�!"Oh�8`/�;�\���Ǩ-N^��P"O֕Je�	�O��Z�ǐ31���"Oڭ*cF1+0�Dp0eћE+�-S�"O  ������;��,T"��"O=� ��Z�([�c�S��u:�"O�DA���)��1s��0RՒ�"Ol��dC�
��K��K�G���+�"Ojq;qC\�MɌm�6KD�C�fhI�"O��˲̈	%0�\z����Sn.���"O0���( \<�j�Y�"O��ʖ�P��fE(]\�T8�"O1:!͈/8�v%zB�ؘ)Q(���"O,��v���*�W�]�A;�(I!�R�<��a�&�A�����b�=\-!��ҟV�`ԫ���R�:� f�	,�!�P�pFD��k����䝙;�!�$��$����Ah@� ��Q�Z/�F�ȓ!�r���b��rW�y�da�-[��	��.az�j(  6ޤ� � {�"�ȓK\f�`D�mE���DI�=D� ��>��Y�����`_����;�%�ȓuF�A�ǈ�
&���n 2�(�ȓ;������t����M�{�t�ȓHNy��*��$��0�aM� !p��ȓOTBH���K�ÆMR%��(R4���i	��:@Ԭ<��"3��&v�r��ȓzH(l��K_�\�2uz��Q���D{�O~D������atP��ԂQ%�du�	�'Ⱥ�:�����u+s�J�tT 4��'����+��V�n�!��k�L���'��]Q��]H���kG-��e>hБ�'n�L1���a�+\KPl��'Z`�KD�ȸb��a+G�	��0�'��c����~��q$�sIZ��'�DĚ��,C�rTP!��r1
�@
�'����L[�
}��*I��2z��
�'�	�vK 6K�Q1�U�/�Э�	�'���a]��Q�)f���'��d��K����)0�X�k�����'���R�GR�1zu/�,�� �ȓ0}FM �@�o`��dl��MG��v+�ۀH��~��d�㌚�k�hC䉅 ����`?e��h�#'�1)�0C�ɚ.N<#�i�i,��st��aC�0�L!X�k^�0MNL�	�l�<C�ɷY���kG��S�O�>"aC�	?n
�������{��M3k7B�I�M��*�cܔV�92�N�5w)PB䉘R��ܰ���v"�uCShח+�jC�I>w��	Ʌ`��;�R)�!hV��B䉺>{���2-I�{�&0��U�7�C�I>3'���iK�p4��M��C�I-I�<u�#*�0*��X5��6G�B䉬C`��aBK!��ġ�gQ�*�B��	�*��͘�.����P*I/BC�)� ���u��Vc�Lx���kTiZ�"Oc�G.4�,��cA�A��x"O���G�.w(�`�!�,f�lja"O��[�	�!Pz�Ђc��3���i"O�8Tɀ�R�����L�}�y�"O$�ȡ�W�-ǘy�6_Kb�Y"O�e��뜛6�HE����%29����Ie>i�a�@6Y2a'�Zf �G� D����T�"H������&Dz�?D����n�,���ǋP/t1���>D�����&ZTjC�d���qT >D��#���"Hg�=�KMtX�pA� D�Ăw�R'����HO)��X��)D��1�.��0E�D�eD�w�ڐ�3
"<Od�d'�P�dZ��ې"i���f�/�C䉫:C6x�G#ƭu=Vx�DEQGOrB�I�J�Q�VN�5�@�"(�< ��C�튑8�\�L�.<��N����C�ɂY?����a|l��Տ
�th�C�I��9���ݹ}m�0����;"��B�I�YԄ��B��#�|����G�6�2B��5@� ��Ø�u|������@
B�I�&���w�C�xW�|���Ȕ�<C�	8K��؋�A	M��<���G0O�C�� 1�6�F� }2 	��R0"wC�4,��MҔ
C�8x(���x��C�I	9M�p1p�U���d�P�ǠC�	A�P�Q��ˌ8�iz�:P�C䉛#L%�t(�YH�2���F3�C�	�[v��bch��F���`'�4��C�I�xi8����P��u�0-��TM�C䉨]H"� L��9-�ihw��T^C�	08o��h�R����1�oT"TFC�I�=r]#s�I1s��	��P�%�ZB�=�2���Yp�`LY U��B�	7f��l�nE=U\�0�m�u
�B�I
��|�4�S�*�r�#�{�B�ɹD�0%	Ø#j���ji�|�RB�	�pIL�{�Nˀ7���S��ͪ�FB�	 d�Q��i]z}9���>Kx@B�	srJ�
3ܝ �)X�
�%?��C�	�4�B	HA�
{��{�k�3*/�C�	�m���2��	�$I�*�2�C�I,.�L�Ց=\U�G�X�ts�B� \���+�͊�/<��T	ۡdL�B�I���"B��S�N9���=F�hB�I[�2��L�ND�	�&�%O�B�I�xV�����črI\L���Yp�C�	36 Xi��Ԡwġ��2c�bC䉼	X�X�KWC�L�i`��Z�>C�	�Y�:D�n�j�8�%�-�B�ɪIj %�V�&p��bO�,|�B�I�	�xF���u�L��q-ŻqB�	�6aB��3#%�00a*�
B�I7	$�6"ץ.W�Q�BϞU�B�Ʌtl����AɆ)�޵��ʝc%�C�I>E�xAC���_�¹K��B�rC䉭F�XI0o��]d���|�(B�	\)@C �M93����
J� ��C䉏u|Ճu�M$E�\`G&���B��0:8��"iS-O�ؒ��E"~yC�	3F���N/#��!	ŷ!��C�	�sxz��͇+��P!֓rh�C�I:"r���"�~H�P+�H!��C�)� J���- <��ر��d �=� "O�͉���GФy���3弁�$"O�a	}�P�� �҉C�0(ك"Oth@B��piK�	!����e"O�4��$h%NT�EꙂ��:�"O�8:'A69R Y�f.�$Հa�Q"O��m�v�Ÿ��W�k����"OjX13j�b�T�I#�m|�(r�"O����\�;R4�	C�0n��2�"O!��<,�9��@vZ�䳔"O����+]4=���wO�\@���"O�i��E��U�ӈ®Z0���f"Of��F��,6ap�+s-Q6W � `F"O&�ڢ,��A0�lF�x� Dk�"O���	ʻU#ByIWꔆ�� *�"O��ȴ���{K���b���_���A"O�Z��т|jq ���uju�"O�ͱP�ԦQ������/Mm��[�"O(��7@
+ev�9h�J�3z��ʳ"O H�#I�Cm[�A+S�J��a"O���p�B�&�,��8�H��yΞ�j��J7�-R��|�����y"!O���)۷�RCT�����yr���HF�^NA[�̩i��Q�'F$�c1":��Y[�G�7_�����'���*�dI�X1�(# ���F^���'�|�ǩ/A�jw@�y�x�[�'`& � ����9��癆n�te�
�'*d�A�C�O!�AS�烑`2��Z	�'-@���	� ޑ[�Q��D��'��<�$ʭ7�� ��MI�NQ(1c
�'����lC�J��#PcDz]��r�'�6�@b�ʬiZ��y���wU�(p	�'�ܢUʛ�\n2�%�ƎCVx��'�t�:��J8 ��x{��ӿE8�c�'�Fy�C�1S���dI
J�lP��'G���J���l\`�=&���'�N�"��>S������dXvU��'��Yz
/d�(%"���<*���'I��j�NP��t�'2�0�� �<}x�!Z�#���1�'���A�D�c�&G,G|�$ �'��cn	�.���`P�*0�}�
����͟	<���P��Fɺ�h$D��2�K�� )��1��3txՙN(D��aAL��@�_�h�c����4xB��7eT({Vk،�~�ɂ�S�]˰B��2/�zlAcJӮF��%�f�KF�rB�ɀP3���$���V�d�j�čwNB�	 ����G���$�Ä��I��C䉫Q8p�Ճ�Jݲ,
�D�5m�C�ɝ^��d)Ŕq���`�A.R�nC�
vl� ^*P,�z�"ڈC�ɑ�:���k�#+��A�%�5�B�I�k��<�$)^M���iE	F�jB䉜W��i�7⑀+n�E��z�DB�I!Q�P9k�%T�d8q�Z2Q@�C�I)-L��J�<F�:����
�mB�-iz�J
��#H�ECPL�U�C�ɮ8"��&�ֺ2�H5j���yB�C�+T6�CWL�4�LEI�m��t�C䉹0|�-l��'U���kG:D���4�V��T<��d���	e�2D�\
�E��ܱP=c�|�c�k+D�� �X��EH`�}!���+�F0+�"O*����'2�,��@�:�H�*�"O� ��ˠ^F�x����{,�xA"O�ٛ���TA�ĉ�T �$"O�lP���
�B!�p-
k>�3�"O�i����7_�}I�̘�,[����"O��cV��:j�kZ)t���@a"OP1;�[�&*���U�F�|� ��"O��R��C��`"�C}��sR"O`,bvI�6�$%B�ѡ0Զ�P�"O�R�NR�/�R	9 $X#�T{�"Oܨ(!敡ce,th�@ى�fe��"OD<2we���@�e��xuɷ"O�p��/e��P���0���"OvP"��qNĄ�%Ci��e{�"O*y��!§����c
�x~��"O҈��ES>a�*l���=\C��"Ob@Z�MԲ��cC���_"
�ye"Oޡ��,N>W���&��i���9&"OpLӄ��"j��*Ǣ�%2<Z��p"O�|B���q�B`���I!	�&"OH�V�S#yj�t*v�-r8�%"Oܙ��_�Z� ��P�
y��8�"O"5+$��<`�0e�B����jUx"O�%q��PQCR�Zs�S�j}0��c"O ې��6(�~d��IbFU�"O��&�]d�◨�W=^��S"O��7L»��!
�hC�c�uB"O���w"G�&�����E�_�f�#B"O�]�`"U�L���$��(��A"O�ɲ�b�&oϸAPe�-��I	�"O��YѦ��m��9�I���9e"OHɲ��SzF�u�?�Te��"Od��-�y4	0F�N���U��"O� ���ޝj�d|
r��1:�\��"O�8�h� �0����R���"O����n�=(ڪuqЪ��ݠ(��"O���1ۺ�pR�H�|�i$"Of�`E.D��ƢկR�u��"O�L硇1��$�G"�����"OpPC��k � ��%�`#5"OP(�W�6!b�ɒjː p��X"O"����[���V�ޮ_Uِ�"O$i14+��L�@�N��I��t�"O����6�"e �J��]��"O|�����J>�L�BW?� i�7"OZ��W��m	޹ ��ĸa�>�rE"OJp�ǅ	>��ق���Jt���R"OI� .T<Y#��kb�`�D"O�|�a�T�)�d�ۙU��L�T"O���%�"&! %��⌈@ݤ��d"Oz�je�̕Z�H�H��&�m87"O.Y���P`ˠ;��4��"O�9�c ܤA��u�ƭ|����"O(<Pt'��Q�$YZ��,nua��"Oj�rƊN�6��7�Xl`�*4"O���g�g��1ň%R���#*OHm� (]�=pġ���2m�UR�'^�,"���!WJ���-����'M��[䋛 �1i$�R<
�lE��'�Li���טhM%I$�L�6���'rA�$�*Z�L`�THІ:�h0I�'���W�J��� ��˞1�"1��'ȸ����6)�\tR���:@������ |4����}�x��G@���*Xy%"O��q��\PIF���oV=
��-��"O�D��ɑ�5@�aS-�=h�Jx�"O���c�X�(��P��9�RH�f"O�(G�� .X<�#-¸U���A"OL��%%ͺ�|�bˁ2Y۸�t"O�8��/�J�p�)��7�Y�"O0@�($)�QC��/.��,��"OV}Ƥ��A.����F�d�b%"OV=�!Ǜ-J񃄦D0h(����"O`d��I�l�V`��Ж~? �b�"OH�S�� H�Dp��,�x��"O���7H���mR�!+z��#R"O:�:���9؞@�Vo�e��H�"O���7��R]&�� O�^��t"O�1R��M4]&�@�$/�>>����"O�fNӹ	�E�7��j��"O�� 7&ۛC�(I�@ߩ3��	�"O���f/�6	%��Kb��'2����"Ox$a'%�oצ���ޔH����3"OVAh��N6�PE�W+�H�Pu��"Ov5;Q��N�;�/ܬ	x ���"O&�h� ў(�jI��hI1H��;"O
����L�f$st��%GX���"O$-��nN� �1�DHW�.���s"O��q������0�˔>����"O��!VNF�|yXc@�K�l�"O,(�Ӥj:�0tE�Q�P耄"Op�#�.^�?E8hr�E�5W~ra"�"O�	{��T/{	���ӣ"=q��
�"Ojp��[�7Cd�c- y��1�F"O��q/J�>�1���GC�ֽ��"O��y��8v-�����ޤ.�p-�$"O���B��f�p
EM	/6��$)@"O��J���(��%���«C�
8�"O*Q��l
gߪMp(>���Yt"O�����ɞd�d��F�8,��i;�"O�y)E����I�=/s|�;6"O�9�6���h�	 ��̧N^�k"O>q�@%O?I_�(q֤�P�4��"O\��N��:F����A�P�\u�q"O|�G���	NĻwv��$"O�rC�V��t�3I (f���"Od�L�2��r�A0cjyQ"O>�痎���!.���� F"O� ��)�p�� �g�8]�U"Op��`�Hv+��ZP煤g�t�C"O��
M'fG�yA&��d@�A"O6�Rw��&H4x�C��&���t"O�\��8 ��애�v�"O�T;�!t�P��m��<��B"O�3�ʘ)���.�5f�(d��"O���g�cq<���#А.I���d"O<�8�-f|�9 �Z9C�=q"Oh�PW��?C�h`�C@� X��"O�S����/�D��o9=��(�"O���lE�����uߘ!`�"O���0�ջ��D�O�\�P]�"O@D3�΂P�hm�Q���wQ>pч"OV �D�gp��!�N��BJ�qk�"O��b�b�����T��w�4蚓"O��@�H�NyV4򂍖?�R��g"OI9B�S�u�(y�'�Z J����D"O���V���&�f���+���ȁ8"O� r��ŀ�Z$� kK����q"O"�X,�y���ÉQ k���e"O���TA�-�ꆦ�N�lѻU�'<�'� t b��1i��K%���|�x
�'܎PAEË3<F͉T�FQ�L�	�'��YӉעHTT�B��E$�4A
�'KR��A��1I�A�B��H�ڵPH<		�_�t��"	�  z譚&O�"!�9��	@����<I��'i�4ͳ��[���iA[r�<�tÂ�y�L�6�� Pm P�&.Wl�'xQ?�YB� �E7��u��i�<`RG�?�Iq����ªR�&+>�[$!�?�������D{��)�3=���靹5r���4萇L!�̻rd�tP$-2Gt�:u拺n��-?�ӓQdX���*��u9��	�oc�ap�<4�4�6W�F� 5��gk�p�G�?D�,�vlHOL�����c/�<A�!2}�)�ӭ?$2����,+xi5��3U��B�ɭc��Y�ō@~R��Fj:0��B�		C�ԑe�=kf۳��#1C�B�m��`LS�:�G	ưb�B��3B����]9�]��C�rb�B�I�P��0��NΘnDx�����+��p	�'+(H��H�iȔ��a��9|��'���遧�x�ݑqk�#���-O\7k�J����@��3�Ǽ*�~E��	V�P!�J���d�5�K�t� ��eIS�Em!�DS���S�Sl�i#�;7h�|�xr�T� �� ,��%X�o���y�ՒN��� %��
�<c�gR�yA� Qg��,]�gԋG���y�E���H6��,?��9�����hO�>Q���:�z���Yl��K��#D� �����0���^?)�����'D�����ۺ�~]���Z�fn��@��tF}��Z�
����o~<T�vǝI�0���6��5Y���'�T� �9H�0F�yrቍy��E%�]yV��:�̂�d�'��T�)��I�p�)�'��P(��>@����ɵ?,.u����gQ�gOCUqZB��8'8x2��98E��;D,b�Ԇ�	%p�a`cY�nk��+#'�+%��C��9J��h��
K�p @A����-�I0l�� �5�@V�X [�	�%t����by��|ZwQ>��'�M`�$@4Fī$'���)D��y����rEb�i@,��`�ĸr�l2D�X*�]
&eC��C 8��t��#D�@I珟�h���Z���L���!�.4D� �ѫ�%lp4�ku�M�d	��� ���hO�4˓L���Z��.c,���
����ȓ3�4�	�'E,��#F9E�p��G���"*ޏJ�˧J�
M񸉅�NC�:�̜�0g�[�(J�W�$�Fz��'��{�KH� P����*��'��p�RO��	�ף|��	�'���AV�X�`|�gɽv�J�r�'����� dlT�bh��$�Ь��'Z�iB�@5{,�C��X�d�,y��'�M T�AE�=)Ճ__�T�"�'bx9[�ÖHN�.Ik�zV�]�<�sl�H� �P�#�6|,�a�V�<�U���k��e`TdQ�(G\8��AT�<���p�~���-<�D�WR�<9�f��}Wx�dD[$vyv8�SN�V�<� : �7�ͮY��u��&1d��"O�)�w�8�"D�FY����!�"OHE����_��i�f,�@�j@�'"O���a@:O&p�L��1<�MH�xb�)��	T|Й�Q��S�,�Z���6�6�)�(�f���+�\m���Rb�i8��!D��ہ�;gyd��g�u����Վ �OO:\�d	�Z��-�#9� ��6"OH ��D>\`P �Z0q�!C&"O�-P0jA&
�搡oڊk�:Fn9�S��y��O�t|����i(6�*p��"5��'��S��?	�� vD
����u �Yd�V�<���,^��u
"G-P��X�NǨ�~r�$3��1�z��G,�{��"�Ҥm�����F�<�R����T�:�BQ�6C�	��><J�덁�ԕ81e�6!hb�Dy��a�5#րR�'� o���vJC��~"S�Ї�ɱ?9��$��20���`E�1FB�	zz�TU�W!"���6�E�M!�@i�'�܋ AB�XDЩ���>Ǯyb��Ov�O`�=�O#"��	���II�[�`A{�' ���'�ֿjC��o�\��'������U��h`8ZfT�����0��<(���Z��$R���� ��	$$��2�oB�j���ƅ�O�l#<y����<�&7���L�>t<�1��F�N�<��oQ\vسk�=�24
��I�<�P��l�ޜ��'���aU���<���U!!E��`5mғ&��0��g?	K<��O�>���M�u��T���E���p��2D�(	�%���(ȳC.�� �:T��0��6�Sܧ�L	�kD�;^����T& �ȓ
	*\�� A�f�f,�AI��=85���?���D�4=��`H�m�	�&J�Ȧ$�Ȗ����ev�0 `OU�)���`�R�!��Ʌ�VE�u���Ծ8B|�el��2d��Y�'V�X0$�և(��;��[��@�'������(R��e{���Y ���'ў�}"���5SԄ����3�P��U�Ii�<�SnJ�Tg���&�09&=�6j_{�<��h���}2F%T�f�2����u����I�{�fQ�f�6�D�2_vEXvM^3���<%u!���OL�:Ǭu��L
��}�|�Ӗ>	�������O���vD��TkTբ"��U��hO1��4�V��5�BT�'�Q���}�����O�L��I�-�zq��
��}�0@bLa�fB��#V>�#g]�l��uH@cK}h�<��'��U����J��ɠv���(0ۓ&���O&T�`��m^|a���+a�
�'J�I2����`���	��r�'���(1K>)ph*Ku�D)�'{5I$邾[En	�M�$i��AB�'X���QK^�著��h��"�'�Lș���z%΄�7�I�Za`$��'aX�#U��3j�� �e�{T��'���-�O�y�`�ـMa�$�&��#&%���W�'�	�xM��z�'[���F�K.C�	(EU�PP'i_N���#�	�
3^���>}���;��y�j۠+5"d�CK��y��CR�lF�<�6�c�/˚w�Q�(�Oiz����%!���C.p8���'�=�m�[qHX�6mP�Y�'d���-��#���r˟d�ltk�'��5��bޒ����G���2e�h�<� ē�J_=D�\{e�[����B�'�ў4��N�)5߄����H�X	���>��'	a|��&7�|̙��ުv��B���y��R�](�Ho�L�����y�&Bb��H��AW������yR	�9Z6y�hF([�`�����y�.�3]�踣����W��Uq��Ϩ�yr��枭[�B
e�rL�ŝ�y�%R&S�@���V�6P��<�yblإHZD ÅT�c�\y��"���y��xT�8��6a)
L ��M��ybK�1�P���P&L-�B��y���ZD�D2늛��Ȗ����yBj�
L� ��b�1<G����y�'�L�\��S��7,1p&	���yRd��-1Z�j���\7\Ivi��y"�µ>{	�wl��M��` �����y��6���4�MP���U(���y��]wP2����C2�+E�M��y��XG�D���ϪE�>�*����yR��x(�q�W�T|�#�_��yR��vI� h�@�#M6��� $�yh�#�4"����x-��y����B9�Dh��N�F6��#s�ۛ�yR��?K"�=�Ā)@L d���\��y�"ÇeXv<C�!*0�Qx��6�yr�C3->���0Eآ\�L$�����y"���->i����~�(
�b���y�E��LLș[�GB�d���HA�y�'�/A���!�Z56�8��A#K�y�aP�)��Qm�*g�4$�Է�yRÃ�$ ��uܳm�r[����y2M�v m
u/j[��'É��y՞{5T����ê9�z)�@홄�y��ʕ4�R�ʱoɽ6X�īQE���y�ʀ�h�D�!(�/�Ľ����yR(GI`fš3`��({��ȱ�Q�y�!6� ��tɜ*JlL����X(�yr��	_�$=@*Np�ν�3�T�ވOpLH�S' '\��:pp���!;Op�#n����&D�Bb~�)�"O\��&"�M�Vi�A C� $< �"O8���*�a�@!��ҭ*��Uw"Oȁ�%Dm�Iyfꀕ� ���"OBL��Ù�>�!s�OדY)�`�"O�@ɕ��"mg��Aq�O�n>~ȉ!"Ot�� ��<QH�g-"@X��"ONPA��j^.���˛0=2A"O<���쒖9�n@��
�+6?.��2"O�|Q�Y	<���C����H�"O&%x��ğ p��+f��8�"O>!�pǓ&s��&�a�	��"O8�KT�$>z؀�e��4�x���"O�a�CҲ�T����I�ȴ�9�"O"Q%G�����3K�+*���"O�����3@Z-KS��g��W"Oؽ�	����E�a�9x��d s"Or���4e�`��� g.vl�"O���S.B.T�ɡ�T4qFl"�"OV��
5mlP�l��Ts��K�"ON}Ss�Q��:���.Zx� "O�|{�)ʺ	26hbR
�j\��XA"O�9Qso+:{P2�Q7NC�A�"On�R.�>�J�r"�*A��k�"OЁQ�g��h�� ]� k�up�"O� ��b�2."�R���ufbY�"O�(��b�|���	n~1�S"O�˖�s%֩K��S5
`q"O��U�U� ꪴ�B�[+]�\$`U"O�hQ�V�[���`EX�����"O�Lxa剦L�8�UDYQt�2�	.Q?ͳ�/�:M��@A�C	ZhFK5D�$zp��'9�HCT�M����W��O�m�ӡ-�)�r� 94�U�\�(�cَ+�~=��'x��*��	41�ƌ V#گ!*|�ɮO���f����=)�Mգx�0���17�<����oX�hRc�\!ɕ]?�#'Ղ_�
�hBZ'�y"� )#��k��F/@d�A���HOJ�`I��h���w�� �.�JF�]"t8Y�"O�L��D3l&ظ�Ě�V(.�`�i���0�fD�S��M���jG葊��L06h �S|�<ao�0x�BEЗ���fl
�cPHl}2�B?wKn=��2o=�[��(�����&��9n���d]�;m���/���V�>m<8c����xM"B�	�n&f��rpҕ����|B��.���2HsĀ�b�dɇBB�ɇ~�^�[w��43��EJv �,. C�+X40�/Ɉ �<r��Q�8%�B�I8iHR�8�a��d�1~82""O�d0O!{�z�˕�_(f���3Of�'ꗾ]���pf=<O|`�ߞB$4�b�O��z�z���'���u/�/�����	��\�HP ��`�>�eOD9P4��
O��;����oE�T���#���*t]b�1��4j��T���M���O�nE)���3
(d2�F!mv8	�'(���O�>;]���gF�ه�/�.���Ф,��kf� ���ʓj}���&��E���瓳6F���Ɠx�\0�a�[���
�� ���i�f-����,xgl��& ��*���p��	�S�ʩ��� �S�"Lk�l��pո��	G�>U��"Y7�msJ8l���pOH)0�.�I�.�1S�N��V+� ����$]]���Q�k �dh~	 ��+Z�����2���T���3�Kһ;�vЌ/@��Sq���1
�>`���UC�)<��i�ȓv�p��DȲ?[,̳�n_%��Z�@
�B��3%=H��<�%lܧuy�
Amv�0�τ�kuf �GN�)Ks�鰡k7� į�;����̘$�+���*����Y�.�ܨ��]2F���A���9���G{� �
�l�@�_��  ���0<�GK�8���h���lM�P*�d��Hͣ�χ�]>�1b.@�y�5*!H��8�z�P��$�1u�ͫc 0asp�ؕfn���'�l� �0(��̫�Q�1���1���'o���\>�*W�^Lhc�ʝ
��3�m,D�JB't�e��[�c�ذ�-̢!~��gY��bv��� &?�"
M��杷Һi�`�;����Eg�D��B�	7ְ1�N̺\��Q.��z|i��#�Ҁ��A�<�xA�`B^�)�`N���HO�� r��>}�� htj�k>����'.��C�怢Wʜ��-�Y9f�I�aJr�Qb�
^�:a�R�Q��	Q&��$^}���'�RHQ�H)uh �JтE� �O�L��bż7�:ҁ�މ..�)q.^.V�c�Ȃ#����W�-�j�Y��鎘Z%�U�yǕ	��Q�$h<�y[p˴	yH�,>شPz�_s֤%8�9�N�O�is���y7o�}'��O�<
E����*�x��"�qB�L�}�t`��c�:N�0���A��"�؜�G�FZ2*��4NR�z.�1�ɍi�'$`��+�� Q���vD�x#U�	ÓY�����4'���{q(?�d��@�i�i8ai��ۦ��<4��[��������\{\H�?/qd� �F�I<]�ܒG�֝�؊!��N\��g��-x d���؟���(j��PPf�$3]� p�"Ov��b��$1&�S3�B�qKj��hV+�8eB�B33�:�B���-�t��J?]��	,X�]Q+�xণ�&�����G�+��B�	P)�\�S�	-\�$`;E	
�<D=��͋%<��Ț�jC4W��<��d�+ذL�3L�,X�Q�<�"a�"�P���l̿>1�4��f:On\ZE^�2����S��m�`5�*cf�����)�"���K6��wF),����^(�}rV��6qhqw!G�]�:�'m���n�)��iȣ�E�K�Z㢆,!�*ਂ��?a�-(_��g���
X�� � D�� k��~xT�Ò�G�8�N|)���5�������/�p���̄�{K~�Ӭ���]!�Ƽ��aд|�3��x-���]�����dQ�,	�\��ӎ5tx�*ڞ*K���M4M/:�xӁ��?���}�$��SJ�m�brF�����d	6R�
�)�FŇF�.�#d�J�RL���d�+G6�p��:}ƪ8�d}�Ȱ
�Oy,���mF{�XHR�o�+0�؁�=闩�l�Hm�#I��m0���b�?ek�O�D��ff��^����Ą�Hg^P��'6�� ϔ�T��IJC�qT-JCÞ;�JUQ�
�E�6P��"46�#|���>�x��G^ƨ�1�U�~��ģ�"Or�F)6��̳%OڲDD�(�#?O��ihK<Z�%CTD/?i��䕩0v6eb�
,@��pk�H�/�!�d�Z�	��,^Ѱ�U��N��I���>iS����V�iw�,_����eUvx���O^�xq�"^�)���]�18�!�'���M�>/��p�V`6��=���{�<���O�jn�ys/ܳ�H����%�T� ��_�n�"��-HBB�I=	�.(Z#�ʜY�j�{�k^4%�ܛ���4���/�5��I+p��Q����b߳o:��p�K )f�q�a)�O L!CNHH��@���~ L9�a�6'AD��'�.(�5P�'"�O��pD�9c��@3�#&Vl��S�I
Mf02&�1Vg���}Jǉ2NwХ�eυL8R!�У�G�<Y��Y�s=�-����wن T�F�<)�ĈQ�j����<� }��C�<a7b� a���WIL� �Z�۳)Cy�<a�LB'��8�cSQ�����n�p�<) ��4E�e�ĉf���(��l�<��t�Fl�Ո��T�+��@�<�D�֪2�����Nn���R^~�<P@�<r6t�M�7�E�4��t�<q���L���Bc�[�J�R~�<�1IF ~��"Ƌ� >�����@�<y@�(���� �8����x�<vg8;ExPؔm	>�t�:QO�x�<ïUL�0����׋ ���� ]^�<��D�D�HC�$�5��_�<	AKՁ;�\2����Hp��G�<Y�U�V%{ Ə~���v��J�<�5._9vA�A���
k��[�Eo�<��		Ӏ�!�L������Kf�<��)�u�,	�+�$WhF�!w�Q_�5�Ԝ+�J~����U:��jM�Nk�� t�Yr�<���X�[��}WIK	c�hL{�.�KZ1Ol@S��9�3}�c�X�nM�׏�3Ȭ(A�O�Őx�V/L�j$�B�.�ȳ� �TV����ǀ+W�~2A�y�8�Z�
�G�.Axgܵ��<��j԰%�FA�H�8q�#�k��l!ǍEۜ=�H>D�4��J55��r� ��o���)T�!�ā�j�r5�#�&��i��,�삕E"Y�0�(Ӎ0�!�d/=P����˷B^-��^�H��K>��M�����'pC�H>S�n��&�`���'������P+v�C�X,�&tKt�-hp
t9��'#X��#�H@$@Va�q�&��?	�p�����+8���(	+1)��q��AYbB�I�Y�X�;dC�-�����PdOv!T��6s�6�O��p�B`ղ#����A-ޙX�R�z"O
��FJ�Ta�I� �O�a�HEO�!��'�p5��>�इ�S�4��ԪY�;��\K�*�b�<�gGAx���S�͐/.�!�qLB�xt�7�'o�l8�*Ĕ,���� ��@��'�^`X퀯�tMqSM7�j�3�'�JUH'��RZ��Տ��Zd�
�')ZH!�Ɩ�c��a�U�ՆZ(��	�'�&��1-�K�ք*E`���	�'���:MSc~y�18�f����� �43�J\�7�V|���Ϲt���� "O�����̡DY�U!1�dj}�"O�����
�$�r��Vα�"O�� �!0;n:XБF��]�nDH�"O�}9�B�r�Z8���ZLC"O��I��\�t@.`��&A�^�~�8�"O�p�ő�y��la0�98R�Zv"O��kb ��>w��������;Zz��3�>4Pl
�`@�z�BQ�ȓ)sT �Q�� UR����Y�"���ȓ1R�zT�0���"e��� ��ȓ]�
u�s���i���٣e�=M D�ȓB�6������(�3B
?~vd�ȓ+�h�����Pk�!��x7�	�ȓ?ޠ ��ϜL9��r �L�6��ȓT�4Ԁ�iЉep\m
���\����F�du#���7E�(Zv�]$�ޡ�ȓ@�Y�0���\lt����z�Ԅ�/�R���ą'y��`��2�@h��wD����!g�)!�
V�Zq�ȓ:5`�i��O�-��Ęv��/��$��v��E���o�D)��<)�T��ȓ1{��,j��aY�P3�蹆�n�`�b3F��I]�	�*�(k�$���qX|��E� ����X�X�ȓ}�\���aW�BJ�+�0�p�ȓ%%Z��.W7]�����o����p�� b�C(�M����'�A)�'LV���L�	~�X� $l1Bx�'��XJ @�8?���;��0���'�i�ċ
�S���ѣڇ1a���
�'�ܣУ����[�i�"�>�+
�'�DyK�8s�o�P�'����G*�0�0S���e��s�'���1KTu��i{%��Q�dy
�'\�T�T��/2��Q�JB�I�8�J�'~&��GX)/
f<�f��(�=X�']`�y�L�H8��b K#2F��'j��EHv��x�S.�%��P�'���:u.9;N��zn���<�	�'���r$���_肈�"B���̥��'T�L�E�2AG�p�A�%��$@�']\��Î7�pȡ�X�-Y&��
�'���ٗ"ƛC!]yb.Ԡ��h��'6�M3����~uX�ۗ
/����'�I�e:,̎mz#����'Mux�hA�4��!�H
�q,�X�'���s��,
{���솆!NBU�'�|��"��)�T��P���&-Ѕ��'�aAE�ܥ
�F�"FK
7�H�"�'G�|�@"A# �}b�Ɲ3P��t��'h��sG��(G��-��� P�: K	�'?X���+V�)
�,�E�GV6$�R	�'���
�j
k��Q: �	{�>ȣ�'z8�$@@�QƂ	8��+_��y�'3鱢�kɨĻ�hV�qN@���'�`�;ÍT�&��3dT�g��I�' �!���0�0x�E&HHt�b�'���c�Xh��P!�>L #�'���Fm�\n=�Qe��+� ��'V� 1ƍH�?J�ɁK�!&F|)(�'���s�!Źo�؁�٫'~��A�'�阣��<U�8���`Oa�)	�'�>���8 F>���~i� ���� D��'��S��0���q|Z�"Or�G�U�fp�:ԫ��$���[�"O2��ᇝ3jșB�I�8/��iB"O*8{0D�|��t��g��6�~�I�"O�,qs����^Q��Ç���x�"O��+$�L ^��������	�"O��ر炥I�pV� b�:��""Oj�S�Zg(Y˧�R�\`�"Otp��Ǟ"m )�W��:1�p�0"OV%�F	�e6��Lƚ*���@"O�H��"Hm�1p�MM�"܆��R"O��T�Z�tؔĊd+�����"O8���&�*!ڬK���$��mKF"Ot����#
@�Hh�x�>���"O�`���ы2��	ȃ��&m8q��"O(���
B�4���`CϦ6qt�YE"O@�w��,R�]s�B�6S��<�"O��Jh�;�`[#��2Q�� �"O\��DW�6=��T�}�v�R"O�qz *Q'	'>��A-�rj"ɓ%"O�L����_�J\�E��	W��ZB"Of����B��YX#iʩ~A���"Oh�;'a��C�}�s���C�If"O�E󥂎�Pu����+=��`"Oj�S6���Z��Qa���?Z�9�"O2�PAKrr4Dpׂ�k\ ��"OdU2$
�y$�̩e�؟W��}Ӏ"On���c�5��x
��Z����"O�Y�#�@�}�D�S��D%JkdXj$"O"�r�O</ez�ࠬ�Q�xX3�"O�%Ҋ�FZ< �:2e�a F"O��!DBخ8
"��!FCBa�!"O�!9pn^ 	�:X�����+I�4pT"O�=���lJ�2ul.u���2"O2`0b�
�-t����U�&�ZE�5"O`����'1R�!�(A�s��k�"O�3Ն�st��Љ�:&�X%��"OP�3!D�8XY���Q,M(�p�"O��F�H1�	W�8�B@
�"O�P�Ă$@Ad��CL�`a��A"O\�p���f�p`a+� (��ЂV"O����iF��B�$��[� �f"O`<�g`(����(�=�
��P"O2�",��2���7mT�RD10"O 5�%����Q�0u����"O��Gɟ[����l���	��"O*�1�CְE�F�@���� ����"O�trgߒJ͊tkc�Қ6ŉ�"O&�q�!�CG��)o�H���[G"O��pq A1P�ٔ�g�>h�6"O%�"n���RU��\n,3�"O@��f,kW�|hq@�<~~��"O��@0��L���1e�I*��ئ"O�����]�%� ��%
�L���"O2�xaD:a�n�Z���. ����"O�p!;<7����L�g�H�au"O��cN��[U����M�H��,Sg"O�{���% ��胀�=����w"O��3�N�|�؜� ���8�6"OЌ@f,R�m�č���$?lb�°"Ol;ƌH�i��C�,��u38I��"Or��c��w�L��!Q���-�y�rMx��f�@zl,5� k�:�y��1q�ip*Ѵ~_��c��(�y
� ؔ2'熺#WP@�(���$!��"O�D!�c�fD0H��U7-��B0"OX4pe��j���Cf�F�{�"OB��4m��3=F}q4gH�d�)Q"O�UD	9c�b��W'ۋB���3@"O�(Qf��/R��q�Z+p:5:u"O����G�Q��q@""�'nuL�B"O����ײ@�\ 2@�@�[~�9��"O�����A�S����@P;g_��s�"O`]�B/��[��ٺP��/<_�4)@"OU��
!O�v�4��-1���Qc"Op��5���#`*��7:@��"O(�a&o�1��H�KS�.�l�z�"OB�ӵaT�7��x�v�P�'�B"O����#R	?I�(����>O-��CV"O�����u����K9k�ܹI�"O�ͺq-�Y�$�����)��zD"OM���R:�`�`-(
�ʰ#6"O�僛�cy����M�O�R �t"O`<Z�D]X@d��aAɣZ�t�J�"O&�J��dA�]�@K�j���k�"O��e�O]i�-2�-ǠS|@���"Op���h���j�t8"O��w��UTD(ൎ�u�����"Ov���晪t��HF�ֈo��P�"O y@WME�\꺹���_L�n���"Ov���;j���r"ɢ_��l(�"OT����>V���h��B�)P49�"O��Y�L%p�b/�r�2�jq"O|��ӣ�(J`2e�ƢA��0��"O|ŋ��I��(V)�a����"O��Yf�Љ<��rc�N��ʳ"O�	  ,:3
�J��[+-
m;"O�`I���*�. ����6
�A�E"O�8�2@7�D8*��
!-���"O�$@��
�W4Լ+�ND5�]i�"O�d�QbD0`���g�g蠔*$"OD��ĨB�2)�����م_ �9��"Or�� CN�Z=�� �L)*� �"Or,�M�$�̌@Kט&,��I�"O�+6h�l��P(a���-?���"O~=pq��.H���3'�óh 	��"O�h��Ӓ%��5���_�5���"O@ sRi�8IX\H)W &^����D�ЏJ~a�#�tt���%���@�̚x�<�m\��0�����S���As	���c��Y#�U_�g��"ebƀ��P�0���t�!��q�}�Z� ]pO��7@Y*�j����d����"Ғ5c����Cتy�ay��& `�X�ם>i�lV5�DA�bʙk��8��`_{�<��G˛�n�@�H	�R�;cH≓1����v�)�V�H��fNְsK����K)YN�C�ɳ,�n �E M$�<Q��)[4�!�қ|bI�^>�c?OT�K���$V	�"�	�;L���O�!9��	G˂�T�[�R�ҙ�gg�%�� �L8�O�P{&�2`J �0)Q: ��E+��'μ��� w�'�&u�qַ;�I���
� ����(R����bא7���Sa��+g���&�4)�"
R�b�'�b?��1��7vt���ۯYR��c!D� Rg�Q�o=�e�V��U$>1���Уwt1O:=ȓ0�3}�+6&x�C�n�]���$���yb�J
3�jm�f@ؓ_-^�����21���c�6�On�ɵa��;X"�P�wEb�"O<�p���8b�|��i�m[��k�"O� n�æ(ϥli��h�/x����"Oq�i	
c]Ƚ�V"�>H��kb"O@]�`DK��t�E�[���xP"Oj��ҏE	w����k�9H� 4+B"O���Qb*��+���
oW�Z "O��Ԏ�c�$a��L¨TF�k�"O�� G��`��+ƞg#2�a"O��Br �E"4<ي""O�h��'^=#�Ja�u,Z	���F"O��)��-?.�q3*ED�H�¢"O�;4��Yr`)V�ɢ��@+b"O� ��(RE����ʗ�x��j!"O29� ��,f��)��zJ"���"O� �Y���R��R�6�@���"Oڌʐ��((m���3�l�@�"O��`��>_����:��Og�<)�)֡=P�q0��]�TE(v�c�<��VV�r��C"-1(�L�c�<Q��D�v^�r"+�9bf��e�^V�<)Wa�$x5$Qip!� ~1�e$�R�<&)|��	�o�	(g:�	�'�S�<�ŌH�t:A�.�2't(<A�"�k�<�R/@ ���"1N#�iA��c�<q7`��
n�X�It8`�hWe�<�A�5
|���mۉd1fܒ���b�<)��E�$��JC�
�0��H�j�<�S �!�-����=L��u��aa�<q�L]�Q送�0OW)�9xDW�<A ���L�
��Rc�QriA���V�<)%Đ�;
��R�J�(Dhb�i�<9��)�Zp`�ـ`B�P���i�<1@�5Q����g�5.�R��P�BN�<�j�%w� (pI�+/��#���Q�<�wk�o���ȷ��H�ްa,XN�<	��]�D�p45H���AK�<1,�P��AU*�fՆ �FDLA�<�ӁR�t{�١��L'����x�<Fg+JJ�B�g+�:��d�r�<�WJ�@&��']�: r`J��B�<�J��]�r4*�"�54D�y2K�p�������nb܂�J
#�y��rT�p�h�Yg����G��y��P*2�pY��'B��U�ըƟ�y"��I�$x�͂<4
� uJ��y"'��:� yUIJ$!�<a�E���y�n�P�h@B��0W!�D������y�J�x�n�wE�U���NV6وO\l��Q.}�p�Cj�s����֦�)���'5y�1�t�S+D�u��"9�	�D�q������^�u�&�ȹb�Hj����M��sľ�Dx��4.���)�H�7jC���#^���D9�(O�>I�Tb
	4�a�g��98l�7��������P����n�%P:��3,�k�� ����<�����'�� 3e�+�t➌��U�S�Ӭ"ܬ訑�g]��R��\��'�"���ȤL:U	wi� �xL�!Ξ;!~���O⟢}� 
�;^�hI�F �����`��!��2����!*F�Q�N�J�_��!��u������,L�8����\%c�!�M�L�@P�5��XCf0�&Fքs��.���ۘ��)�'v�:8 ��s9
�8��
��Ral��������|�ܴ= �"��0)�^�x��YxV�����<E�ĳi�4I�쓽�mҐ㇩/� pr@�'@���N�^2�2d�O�E���C)\��OA�	�\���E�tb]/w�6����:���c���� �X5��7��)�g�? f��q�DFT���ʒF��y#Ծi9�����b� TQ�O�?��TF�V���pWB^�FU(p(ݪ�?a������z>���A!l����=���Oy��8 T��|cW�O�b?��9�B�f�P�U:f�<�#�̋�Ao�'�a{b�E;3cb�t�T�r���łώ��|��<�~"�0C6�Kņ�:.�*1.�O}�a�O�>��V�6M�����JN��)��+�+l�dۄ��S�kl����Ӝ'U<�h0�âv� B䉵|ܮ��|f(M����"a��C�<F6�X�nĨ��|�0�Ap��C�2�t�
3�>�ܐ��N_�O4fC�Ɇ=�4{ 	�$�-1({c`C�;��H�pH��R{d}�(4>~$C�ɩf�~1j��k�꽠1ID�H��B�*2�����?un��i��h�B��/1�-3���:����܌�B�	&�8��Ɇ�+����7�U7z#�B�	�
���%�H��x��%!4�C�ɗfn�����Ԭa�$�s�2e�,C�Ɂ4/^�s�3ss���W�N$g�C�I�4S��I�"[���s���C�	�$�,(@�pL�4O1C�B�	�wU�y���pX`+uYB�I�GJ���dE�c��L��E�a,(B���9" юD���)�+P�:B�	�j�\���(>z,e9v�YB䉞k�q�AK^�@�D=���׺Xg�C䉸l�ph�o�'6� iP��� �C�3cʖ�y���VD�����o�fC�ɉ0�(�C �؝]҂M�F�P2C䉒#A��Ӈ���x@G�(C�':n��B��g��|�N(h<�B�	\�}�R`�&lQ����Ȕ1;T�B�	;7]>��`\�H��L��`-{�jC�	�U��t�3X�%����bĞmQ|C�	 F@K�灶�lp!�,\C䉐I�!�B@�HX��@�BC8C䉫l�P�dʑLڬ��j� �:B�I(tMЅ:��*�H���bOXB䉱[��	���q���h` Y(w} B�	�QI(`q����c%��!��L�B� jxԙp%D'� M+�@8�B�	����& D0T����$�6i��B�I�s���s�Hq�u@́uC�I�`�������rrA�?��B�I�&��%"S-L"U�ʼ�$��^/�B�	#;�����.�B�R��q�U�e�C�Ʉ8U>X�� ��&}����M�8B�	��$Ԡ�05�֑H�gR1�B�Ɉ!�x�G�	0��y1i��M�BC�Ʉv	�3���:0������5zh܉r �wT��[��ڹ9��Y��V#��	bㄬ���ð/V ^Ȅȓm(�! ɢ#���A�G�_
ń�M	���W�LE L�Nd0�ȓ=i ��U��"���W**�ƴ����x�V�S+T�QjV�ȟ�T��~ޕ�(ȡ8�0�ن�\�Ƞ��dI�e��.�ݰ��9@Ԇȓe�1�Ӂ��wc�pxdH��)~Ri�ȓ<ZLjD��5~ ��%Gϵ5�����h����P�s�´�S/�����h]Α���o�eZ���p��ȓ��@j0H���1�!���t��y��S�? ��%��8�������9�L�E"O�"�A��Q��䠢��16�X��"O(�H� �$&�B�hΝ k8�"O)w�/�L� �m�
l�
G"Ol�, `"P��s+߯5�dk�"OT�1�%R�ȸб��0LxС@"OxRv&�0l����V�{�D�"O}��
ȿF��mZ`lO,�8t:�"O� �� �6#�d
e�����@�"ObL�'�P"�H �! ³~��U�1"O.�Z�aF,�S7@��A�,��0"O�m�@���lL�c��Om����'��Uk"��H.�F y�љ�'
ɲ��I��&�+谬3�'�T̰�,�u�xd�U�U#y����	�'bJ�pI��tM2�̅�v/ 9�'�t\{�싿�����>	���'����CeĽZn�!�W�SeR����D<�V ��{t/S+M�$xC�O-ٴĄ�]ǀ�U��Qsf�iC��%*%D�h���0y����3#�yA0��#D��Q§\�v���0��S�\�A[��4D�\����6G6��D�22����4D�ȨudɅ3�V8HCa�;Wl��U�0D�l!B�#Ku��zv��M@ĸ�A$D��q募�|{�;���� d+��4D��ըT�0t%��L@�i����6�2D�x��;��ȓ����ê�ʧ�,D�(bMLd�L2%�!{՜�`�8D��#�b������j^��`�b5D����W�����@��(��7D��Z�Eէa��h���|7`-��l)D����S�Am���
JYf�Ab�!D�`Y)Ե> ���-ɩ{ʔݢR�?D� 8AiT�W�z��DB=&��]�/>D�|v
� �N%��턡%&p}IpA(D��1�_�<�� s�O֫�(���$D�l��@��i��gO��96 #D�����Լ9���7�9
���-D��rG��	�	A�∜I�����1D���d(8��)��X�oP���R�/D���RfP�
�����IZ%�T̙��*D�x��"�
�0�!�K#z����V�'D�i7�@� "s�K�4��t`6&D�x*�Ȼ3�d]�,� z��|�e !D��&�)L����A�EN4�;w�>D���E[�l�B��!g.A�-:D�lcP�)c���a+^�g�F�!w�9D�����4,����k[�(3��9D��u"��u�zt:�H �S���B�f#D��`��	�	+(�Wƞ�%�t���@/D�l��eO�������\5[lF�Y0h7D��� �	Ar�L�!�\�@�4D� �ǘ�����N�cp��q3D����� I�!�A耞����/D�|zMZ6���!%�@Q�)�s�'D��a�#������x"���I%D� zu�Ld��Wb�P%�F�#D���N P]�+V�/!�Ju�v#%D���%MV�`Ң��%O+5��Y��!D����,�9�2��1� Q�3D�(�U��&p�,�[DO�D�Ĉ�0D��/߄S���B;?��3�j:D�HhՇ�+�JŁ��:(��!qW�9D�� �9�@�/�b�ӑ��2���2�"OX�cQˏ�S�b	h�MӬ>6e!Q"O���8O�i8��L&����"O�D�j��h�z�K�,��
� �B"O�L��*J|Й�[(O���"O��2� Ȇ%����I>x�"���"OFua��fmr�!��D�wz�ĐW"O64�Ņ�) J�1K�0/v0I)�"O
5�g�	�Tp�d�����"O��z�(K��ͩUJ�4E|�u"O�T�a�TC�N��E@�
Gt@�8"O&!��+90ͫg�a���Pw"O��C�Ӓ4ۺ�B2�ĐG���"O�q���F�����Ã��`��a"O����Ƀ.�����#VVq��S"O����)F�j4R�b_�a�pٖ"Oh��fdx2����O�*@�"Oh�j�aJp�F���&B&H�B��"O�,CV�Q-)|\tʥ��6}Y�2�"ON-P�o��j/��D���w��9�"O^��GDX-���#��+-Y���%"O]���ƙ�X��c�<�͈�"O��F+��U��K��G/^��8��"OX�9@�i��h�2C��,��yAE"O�����"d��)���o���"O��b�G�q	� F+8Hd�J�"Oe�m+Y-��!�O_��)�"O���6�4��Ed�;
@�]q�"O̍В��\���j�֛<�4�"O��p,׎_ x���s$6]PC"O��"��N }3b�ҢCB�a��"O��҇��Ae�0�ҁ��!TT2"O��V��7[��
Y�K���"O����8Z�蘁1��8�2�"O�,"�F�0�f ��]=K�|��B"O�+���iW�!R%�>��zT"O�O�Q�U(S'W�N}����Z!�_o����+�S�d��f�
q!�XpƆE��.
�R��9C�%І$~!�$[p�.`��Þ�V�q"��K�w!�T�[��eh 
��x�,	Qү��+�!���k!h�&�"�b��n=B�!�dG���z"L�R#Ve���"�!�D_�*��m�%C�ԮP4�
�/[�<!B2f%d��T��f)x7��T�<�q/�/�<�O-V��\�T�x�<�*�<;��8p�@�+3a��[r�<����a2��U�L#8�y֪�m�<�����-3���A	0���u�<���H��a��Z,j�y�`�t�<I�凿<��S�MӱmȐu��F�<���	7I\:4�U�T�2��`yw�]�<��Ht���j��ސA�La�W�<�@LR@��Y`K�"r ��o�S�<90��/ӈ���B��Ab�xP�VN�<as���y��z���Xf	���G�<!�ID?����&O¯!PP����i�<	F���W�h�;���BF\U�&n�h�<��j��"�,�#��=*6̀` �P�<!3��i\��`�[=,��C��L�<�&�أL��I��"KQ� PU�F�<���"fje�T%ɕ4l19��m�<�g�q�Q�#X�8F��5�	j�<)�/��}��g�����f�<� еSs�ў�l���㙕E�fU��"O��svBN�%��a�ld>h�"Op���
0F�4@�%���|tL�v"O�ᡑ�*�6D��G�v_<	bV"O��*ԧ!J".,�0�A l^�[�"O䙲u�ț/��i�怀B2B�7"O����a�%�8�����.,�h�"Ona
r��.���sl� m�>��"OYӃ��8F.�ۣj�#�<�"O�T���$OF�@Bk�?����s"O�y �܎ApN鰪�	 �z�{w"OZ]�W ՕIe8���:3��R�"O�1� 
  ��   r  P  �  X   1,  �7  �C  !M  �V  �`  �j  ^t  �}  ǆ  a�  L�  �  ��  .�  ��  ��  �  R�  ��  ��  �  ]�  ��  ��  %�  i�  �  � � <  �* }2 �8 �B �I >Q �W �] vc  Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�� |d��"O
`�(�;���8���-0��1%"Oj4��ND^[��"3/9�0|H�"OB���H��*�ʞRy=a"O�味V�!X��!&F�:J�$���"O,��a
���C�Ą�M�"O,$3%o�-���p���+Ն�:1"O��ݢ1����`���y14]2��i�<�6��{_���c�H�`�fX�$Kn�<��A̼VI�xR[�)�Ć�pඤ�ȓA5��('nߡ4�� �)˩%� ���,��r�؊b#`T�eT09���ȓ!�b��g��}�8�F��-? �ȓ
K|m�ș�VṔ���2�%�ȓ"R�X�j�4JN�1�˘X�i����̹	_�jZ��1!g��zܶ��ȓgil,*�J�
j�Ne��i�J%b���f	�(U��:���G��$Y^م�~r�� S�%T"���k\�jx�ȓ|4�1�îJb��@ӵ�ݩn�V��/[`�"�v4�R�!ʎ<��M�ȓ`:��z�ؚh�J�Z��$HY:	��H��p�m�C1��!��B:��0��EnjZA V;9����J[
2���	��4'J�EA�IVW&��~�(aZ��ӹ�>� o�Y�|�ȓ�f�A�
Ο7�H��M�$�����mޠP����/���ANXo*�ȓTv������h ��-7�*h�'��}��zE�	H�N�g
�z���?��') e!�NѬ���C+D�/���	�'�������]���*QR|����u�OH�!:p��O���A1��>y�Ȁ����*��9`Ǥ���t}�ѠܔN48x�Q��t����S�'~&�P7�����KV��r�B��  ��J����*�S��6f��Oz7�2\O����GA\W�f)+�V!�5"O�X)e-��R�"��6Z����"O��hC�Z�Ph(di"f�d�"O�9���Z�w����AG�e������'�ў"~��/0m/�8������``�)�8��ȓ���h#�!� 5��F��j=�'�����0=i�ۮ�"��%	)Hl��ƪ�`?I���k�3�<x����w.P	�GDA&�����%��l�6��[l���  Rhx�ȓ3*^y�.�:gN	�2IA ��E�ȓxBɓg�_F�5�D3�x��ȓw������S�ܵ�S#e׾!�Ip����YȠ�9u��4zׅ��|F���0D�HȂ�^�Q�U:SC7\�:q�D,�=J�D�O��S�$���O����2#鰴H#+ ���p�'e��n?���%��sPz\X��#*��1�'��~����
��ɨ4bΝ2F̤BɅ�hO��O��f�I/v��0���@A�V�ߟ�y��؍<�x��i(^�5��l���y�lE'S*Y;� A2+��Ģ�!��yb��A��y��A$Yjɉ�Է��{Ө�?E�T!H�R��D��lC
��!��yBO�'Nl�
�B�9o���*2�۸'��CS���KϠA82Ɔ�N����G劍Z�F}r�#����	�]�H$rcF��6w�\�с�; � ��=��1,OX�c�`�H-
uP!(O3P��J��Sܓ��π �����}FE��b��R"O��8v��E��[T�l�˷Q���ŀب�y��Ć��g}ʟ�Ű�.�� ��x�udI)'A$a�Q"O������g�
��#
N'6��(1"O�ey7��7{ ;`��1���"Oq�F�
I%|��rHR5MPaA4"OP���O	�,0vy���, b�$�~��9�g?�dh���p�9t� �O�h����r�<��JM*�<�S׉y�L��CAs��	t8��X5���J����iG�(qh��6}R�?�O��:W
�-S���!�޾a(�C&�	XܓaN�I�9��`zE�E�7�4Q��V8R�!�dƐY�zx{�J�J0츊q
�~s�\R�ӛW��l;�.Ng�v �sG�B䉇	:Ep�
�P߆H���]��B�	�y�4 sw� &�rD�T$��`��B�I><]��ȯcـ���@eAzB䉼m�Ũ�I]��d�:�B[? ��C�I�`�Y{aI�E�P�SL�=N��B�I5Z��P�D+z�����.��={|B�I�b���ԀC�k2,i�GTL�j��9�	�CH�c�A��U�B���8�.B䉖(h��sv�O%4�v�C΅�"���D%ғK�P,�D!�
�A�G.U�y�P0�ȓ1���*�)��*� Y�o�8�ȓK((���"وh��0�?@(�(G}���-
>��N��S��@���]���#<�7�|*q�Y;]ib�t�ӎm���{�nW�<�㎀F�B�5-��Z�o���}E{���i�t���B�#J�����T���1�'����S"c��� ��$�p鲧Ɂo���L��I�h%f`��D�E����b�<@6����O��I^�'��6]���BeD���-҃e+rN0���&杩Q��+W�z�AF�&|M�YF" 
D�O�~L1GIO�>w,�R"΁7oD88I>i����@\�9q`���V�L�ڳF��^!�$F�?Al�Z� ��1�����
W����˓)ܼ��C�&Yz��~�ц���l��1�N�c��bR�ȓX���32�?]^lu����TC�`�ȓh���z!��	8(��#U�rD�ȓ>rl!��/ގ(�a��
{u��'��D{��d"�v��j�nF!kxxQ
B��y�!^Xߨ(�����\�.���B;���y��$7�,34A*��J�pb�Q���0'pцȓI�2YI��	+�L���fS�,Frm�ȓyt(኷H�$L�f|zP��M��p�ȓv�~\��D
��F#�)�=Y�����AZ|��t%�9�rPVB��y��(~J<��M	*:��%'ԡ�y��A�Q�P���� U��4o^��y2Ú�_������M�a��,���y���of2a��k�=BN����`[,�yB@�Q����H\���Kܘ�y�H(J+0x�6U��@��݁���T{����$��ߠ�`�5a��w��0t"O(����>;ʽ�p��^f����"O��aB�LqDD[�'�7.�Y(��T�'j��OP!�J]=�n��A&�hT"OZ�*�oZ�B\���gO����Q��a>����ē)�`��n@-Bg�x�)7LO2��/����r���p(�ЕEo�TQP�)�H��(d�S���sX����S̓e��b>e��% ��Dɀw�5��9}��>A�S�? 
�ò���V�r%3��1���IҔxr�:�O�{TŭZ@�w�C69�(��2O\��D��L���s���s �'2�Tѥ1D��1R�ٱR�$���M�O������0��?%(�[�>���� P�v?�D
�)j��G{����+~�* �(_����H�Di�	Z��(� ĀRe4(@b�bw�ۙDNE��"Of�a <,��`��τH*���R��Ip��Oڍ��W�#^浩���0",�H��"OҨs�Hъb����w~� ���>!w�'&N�� E�']�&9�HD9HԸc��~��ģ�l���	���1#�A�5��'�az��)Т, Cj����!��(��Px��B�9�`���ƍY����%4�ȓBT��@�k)��Ju!]�Ґ$����I�P��Ф❢Bfՙ��"B8�B�I�;��xQ2���+��q�g��;�'��)#1���.xD�{V`
I=�|3�'�^ hN�2V�xa�՗	����
�'&�1��%m�Bm�����
�'?j\��E/.{h��g��3
�'�괋a��U��4F�F� "<��	ߓ`�OD��Po�X�*����"O.h��"J�;���!¤ɽE�\M���D}���>�|b�BMq�.�E�3T�\ C�Bx�ܬ<��'���a�DZ�7F�:��2��}H��$&<Oإ���4D�<��(^ۜ1P�|�)N�|����^C������o�pC�	-Z��s��
 b���cŒtAX�|F{҇����D�5dJ|�X`��<�q7�A%"m!�d��%�y+�%�HP��[9ZA!���%��ܣab�	7����Ǒ�!�Dא@(�0)-]7Fh5m���!��DfE4��!�m\��f�B�!�$81Sh��Iʄ,�����`�!�$"[\�F�Ͼx����C�7�!�dQ G��� ��E+h�,عbb]��!��]�1#�>���Цǉ�z�5X�'g�<�7eL�"�r�g ~f����'g4r#/DL�"�!f	��p�.���'��!D(/i�E*�	��i���r�'��yPcfJ*�^,�� .�t	�'*re���|�*���-PN��'2�uT*[�f�|!�q�7����'9I�&2-*cq���Jb 9�'�
B�#\�cL]����`���'�8�`۟
�n��'Ԥ]�X��'`��B�x���
R*�0nZ�'�~��d����=ڦ	H�\s��'+�Eas��)���h���p <I�'�VU˥Eڃ	���&�2o�ddc�'����A[xX4�"P7���I�'��]��(����7�NF|�a��'�4���,��hJX�i��?9D��	�'Yb�(d���G˘5Bb��f�� �'��;�<X���R�� ]��C�'6\D*@���>�� �8M5���',�P�$��� \�g$B<D�d�+�'( Y�DcO.S!����f��<��A{�'��k���G�5��Y:3��-�	�'~~ !�哽0v�bG���<̲	�'��P�UHrn1s�+%����	�'$F�8wC^ �HU��i֠��'��I��+: �x�soS�Z����
��� �R��\Ĝ=0�'WTB&��v"O���B���k�����I�x<��#�"O�-"c���Q1P�z�#�(o4�[ "O}�T(ׯKR�!Z�c͠m�TY�"O��R�ܠU�8�����d��3'�'q��'���'}2�'}R�'��'�����kZ�I~v'_�`����U�'��'��'�b�'���'���'7�pHr@ޡ~6H#sEO�q۬e���'B�'K��'�B�':��'��w��d ���|j��ʁ�F�P�6͹�'<��'G"�'"��'"��'�"�'|\\����D��:h��ٱ�'2�'�B�'/��'�b�'v�'O�)�����`�1��P;��ڵ�'dB�'Q��''r�'"�'A��'".i����:iž��SA��.nT�;��'���'h��'oB�'B�'��'�,xP����b@q�WZs$e)�'���'�R�'|��'G��'�r�'N�%��	�'�����3;l�hۑ�'���'1�'c��'ZR�'.��'힙�C"��w|� 3�����s��'��'���'���'��'�r�'Lp�hqa��p�xZQ��!��@c�'XB�'��'_R�'���'^"�'ΨM`�G�J2	�Gb�@���'c��'?R�'mb�'$"�'J�'m�x(�M˷'Þ��e̃N/L��'���'m��'b�'}�*l����O�����Ƕ}آ����Fq�Q)�lyr�'s�)�3?i��i_����1sB �:�b4l�<�3���������?��<yU�i-��a�P8c�V�Κ7T:��|��$M�_��6/?Ie(ȍ`�G'��'_��zA�量j1��wj�%٘'0bZ��F���8.����N:=�]�֨�6W@�6̓;�1O��?=i���S������<��.sĀi�2�N%���-���q}��T���`�f5O>�B�p�!X�m2�6�+�1Od��a��@�zȨY�ў�� ���K��:��%��h��(�"@g��'��'@p6� �1O�@A!˽EV��6�aX@uGE+�����$���2�4�y�Q��JQ���?O����*9ᶄi�A*?����9
��8�.IQ�'6�|	]wEb�$R�rIS���+�L8j�$a ˓���O?�I�byÒ#�$D�����L;��I��M��Yu~r�p����Ӹ<>N���`����q΄�V�~牻�MӀ�iIR�."����$��RΎ�/�t��ץ~�V��U�2���N����������8/�u��$�5��i�"�'2��I��M#�!ɥ����O��?]�웕'D�]��O՚0]��MV�����榭Z�4A􉧘O(��Z��� ��D����;��DK����nv�ݲb^����K�J��'��o�	[y��Y�1LT��ҋP0)z�u���0>1�i�ꉈ��'O~l��6 ���:	1x([�'
7-!�ɵ��$Zަ���4&=�f�"�"�ۗ�֍!~H�w.�00��8�	B8��DX*Iu`���Z���LI��R�g	��H!%�:zM3���,5�V��F���b��9�F�{ �W�s!�x��&�	&BR�sa���UZԤ�uO�\�D+�,E8���z�r�7� %�2�KT	u����s9�3'Ěf>��맟�D*ڜ#rQ�R��1m4(R��2j��2�$᢭�Ć/_I(؃a�X�77"�!Ӭ�?UD�U�8B�����q�(qB�k �,���
��'Fh8m��
"n�. ��+�j�Ȍ�Eԛe�x��7h�0��QJ	�-R@�0U��\���a䍡%�>��&ɺ61lٟ���Ɵ�����jy��'B�'����}�FQ����sdI��N�.��OBY�B���O>���O��
�.��E`�D�>Z��#)J�5�I$ɂd�'T��'���|Zc�D�x���9^�:�pL�a��٪O����k�O���?����?�/O����բ?��3o�����O���?A��?yM>I���?���,M@C$�F)Y��!�*�%E�x�J>����?������<R���<Pʘ\x$ F�%N����3/$b6��O�d�OԒO�D�O41�$��(�lI�pq��a�4�����G�>	��?����� 0�$ʧ�?a�dN,D9��	���3�0�8%զ���'��'$��'�P�ӏ}�/'vd�:��ܑjl�px�J��Ms��&6ͨ<Qp�����I�O2����89��ߟ(wTԹ���|v&��C	�P�	ϟH�������	U�~
M�msx8����UǢ�C�&�����')D<C��'�r�'9R�O>���\�)� �r�d��#�
'o��+޴�?�J������Ĥ̸0��p�U�O�=݆h:eGԀ�M��㖛�?���?1����-O6�D�O�"���%��A�*פ;^�P��'ɗ�MT.�-�������ڒ0�*P{@�_��68bfL	5"F��lZӟ���ǟ�j"�]y��'r�'V�DF2Z�c�L�8(�����N�@��O�h���O����OFh�co��KZD�k��"R	��耯Ħ9���T��L�'���'O2�|Zc:� 2�˞�߬؛�C�� �Lp�O`�E>��O��d�O��v�����07v�0qTkP1�@`ʱ�U���d�O���O��O��$�O���𭜰+�\(�䬇'lW���E^����$�<a��?����$_�K^4�'E*���d@�/{��r&&�k�x�'�'{�P��I�0���ȟī��I)�����g\ �j0IC�ē�?����d��'� 0'>Ea	� 6q����]4kI�\������i�R�'���̟��ɞ&�¹�	e��G�dJрe�Kn����.�&9��'��]��S��@��ħ�?�����-��3���s�L��W���Eæ��'3��'**����'��<�s���E �<aҊ��7gMu���Ƃu�
ʓrBT�ƽiX�'�?��'��ɰwf
xh��ʯt�(5#6��;=�r7��O^���=#ظ�DSn��?ɗ�M�f�P0�ꉉw�Ũ@��s�J��A� d���Ms���?����&�x�O����A	6�؍�6�a~,e�g)u��Iv��O����O.�d���g~�EIi^6���$D�&�0����X3"7��O����O�� �k�d�i>��I���ل��.�hY�F�fi&��t쑉�M;���?�� r�S�^?�I՟���˟�)᭏�i�ε��Ba炬�&����M���\ �d��x�O���'��ɽi�$�Ѕm�:�0��(@�m۠�2۴�?qA$�	�?1,O\���O��<ٵ�W�iIZIbt�>ɞ$���}L��ڡ�x��'���'������g�L ��J�,�h� đfZ��2A'�ϟ(�'�'����q`JmjFE^�q���O�@l��Ц������?q��?�����d�nZ{��U�eX�U8��l�~��O�s��˓�?!��
)���O4��dDG >Һ���J�c��P��
HѦ��?	��?���j�p�%�س�£u��Ao[�o1޽�tFa� �Ļ<���	�Ve�*�����ON���ȈB��,������	P��2�x��'��gU� �vI:�y���WR�4)�'E͑U7�DQvBG��d�OfQ#�O����O<�����Ӻ#S�&%�RĐ�%? �ԼB�%Q¦E�	JyR	ʅ�O�O|�B ˜�	H�it�S�O��=��4٤���ir�'L��O|&O�ƄJuJ����)#iA��2�j�i��'Nb�',�IK��'/��ԍx�l�ć�:O�{�̠!�6�O��d�OV���]W�i>��	�����V�V�2e�N@�>:d3��M!�M���?+OV�����O,��J�!*�"7��b9�ɑb-_�M]m��,�Rʆ����|R��?�/O(����!�p ���J�h��6��ɦ9�'��|��'��Y�`HĔH�p�x�EZ�Q5����Jݒ> RɚL<���?�����O����xX���d�8=±gȏ'?&6�O�ʓ�?I���$�O�ħ~�2�QyI�`�aO�?ߒYPW�~�����O��8��Wy�IA��M;1,B�
�fݏB�ށk��y}R�'���'��	�{���I|����7�����++U�h���T�xћ��'XrU����K���'�'\b$�h�kU���yB��W%���1�2�'�創���aI|����1o��ȩ�7 ��\JDGLd�R�n\y�'c��'_2����5"U�WT�@p�ʁ==�i��ڮ��$�O�PcM�O��d�O2�����Ӻ�Tɞ4ՠ	���}�t0c�(�����ItyRlƬ�O�O�Ё�I�G�B�b
�Y���޴4B�5�Ƹi���'���O&���	�x��(�@޽�!i�$!��,oZ1,�r����1�S֟�B��8<�l��&�
3���S�U��M���?)��:�j��CR���'b�OH���"�y�.�Y�aA�nt�8yf�i_�'7J5a���I�O���O���5��!�l3��>�]������]����<���4�?���?���7���s?�6�-�zcrD�7]*��0��}}B��(�y�]���	�������x��(A���1��TĎ<���3<��Ig��Mk���?)���?�T\?�'��d>��u@ �V�i���qe�H�'��'�2�'P>i�ƈ]#�M��ǒ�F��5�ƀr(ݺ`��6����'���'G��'���ןd�VFy>�w&��t�`4ɖ/�17�:�S�B^,����O����O`���OB,�d�Eۦ����PJ�	�i إ�4qb�^�MK���?9�����O���b4���d���qA�0Zl������=8��o���d�O����O�=
��Ԧm�	՟�	�?сrb�& )���PeU�,��eB��M������O�u<���O�i�R�����_R��ꠣ3*=H���4�?q��]��(p�i�"�'f��O����'T�#!��p,��I��_2t0,<Ӆ��>i��M]T���?�/O�)&��Q5��VCj
U�����MC�oY#Л��']��'���O}��'bҎA���� L].3�<�h�G�3��6���Qe���8�4������Xn�;��'� ��O���n�՟���ß�X���?�M���?9���?q�Ӻ�%M�8I���I��'u���Ze�Dꦕ��[y"m�'�yʟ$��O��d�8���% �&$���tK�'\&T%�ݴ�?��)�0����'�2�'��`�~�'x���䔇�Ԁ�TݎX(S�O~��6Ot�$�O���ON��&9�P�G^�hBm�j{�\�%ʱ9��m�ߟ��	՟���5��I�<��!$������mnZ��"��w@ݑ�-��<�.O �d�O,�d�O��Q!`x4io�e�<$"&NE)^H�W� �+�B��ݴ�?a���?!��?,Od��	}��S�Hh(�Q��q�.0�n�ɟ���՟��IƟ��	.Wh��ش�?���Ԑ�G���t*�����	R��}QU�i���'W�U�D�ɇ�`�S֟���7�d2P�L!$�����r�\%n�䟸����	�-
xi�4�?A��?��'Q�\p
׮C��f0Ӷd۫*D�c�i��\�P�	��r�i>7��S�r�)��4AgR�0
��w��v�'d�R�Q�@7��O^���O��	�N�$�t�? P���OrB��� ��D@"_���	�Q?Vu�	П��	Y�ԑ~���.�@������i�h]CȂҦ���cX:�Mc��?��������?Q���?�����H���R���^d����Y0����XkB�'�"��~ZK~��G��%J��Ɉq<��
��C�`���D�i���')R(!'gn6��O:��O����O뎊�:+ְ�RL�$dI��"g�@u4�v�'Q�I�`��)���?a�:+L��N�#1_�=����4\��(2�iZb��/ �6-�Of�d�O��$�C���O<��S	)/�ι�F�u�N���W��X1Cd���'F�'���'���rs��[6C#t�ोS����ĨX�Hm�d���O~���O6��O��I��8̇vPz��ʼeДE��/,`�b�	dy��'�r�'�"�'�Lp�ex�� ��+w�6�����pz:���	���E��ğ$�Iß$��Ky��'���M�@� ��ȣ�9,
<��Fo}r�' ��'72�'Z�e��|�>���Ov]�i�(�����"�8&n�;��B��	ܟ`�	Ry��'�I��OKB�OBUR�
�s%����̃�=�X��3�i�R�'���'e��$�u�����O��$�t�ZEبAF0;���3m�(��DC����YyR�';*0�!\������451<� 4�@(?� ���)Z�po�Gy���;)UJ7� w�t�'e���4?�E�Q�k^�ݳ���"?`�*�C]��1����$��D̟�'�b?�q#�m"���Ң�	����� i�<��G-ߦ=���,���?��K<a��)���tG	�4?vM�	2K��B�iO|8�'�ɧ����i�H��&��/报�f�ӑ`�o�������D1�)_����?����~R�=/���{wi��y7�yFo^���'����yr�'N�'��t(��U|��4��k�4�<��`�4�Dʹ
��@$�`��X%��غ#��1Z��p�'/�(�1�O�C5��O�ʓ�?���?�+OTIa�S�qr��Rc�<���e�_+
 �H$�����%� ���ăCn�)0���tӀ�0��R�TJ��IPy"�'a��'@�ɢCS2S�O�h�dLO&	��V�ߞ����O6�$�O֒O4��OD\����O>}���\3�,x+�� ��^�cΌ{}2�'"�'g剮/�d�I|�,�a6Lk�S!fg�ȑg���&�'��'2�'��r�'?�|�ɋ�J,��FUUjD�oן���Ty@��9� �R��蟢�5i�3��M�%��4s����g�y�����I+$���	~�~���1KfL�P�7uBH�p�A����'>��S.b�T��O ��O$�W`Ő�C�m� d��L�S FoZ���	^�&���h�)���a;�x�ge�F��͙�]��7-C�`��!n����I�t�����?�q���N��5j�	��V5E��toZYG.#<�����'�-��W)z 8۰-�>G��##o�l�$�O��dѺK���%�h����`��"���H�8 �{��{u�m�D�	�rz�T)J|2���?i� �8��,�<O���@�Ў�$`Ƴi�"�#��O�i4�o <(27�
6Ld̻�i;PE��l�ǟ�kRkBşD�'+�'<Y���q�LF�T]Q2�E!Iz���'��D{L<����hO��$�v.
��JԘv���"> � B����'&R�'��'��ɇRW4(K�OD�첧ȟ�zJ K#_Șl@�O���8ړ�?��%�?	d�6X素��],g0�4�����A[쟨�	ßl�	����G�Tʧ�?�u���@	_�d[�}1��0M���'1�'���'���f���ēityp�g!5�H��e�V���o����RyB,�3R:�'�?y����A�3�*�p��D =r�9��J�f��H=16>Y�s�@��㌏�CJq�r�	,�L�Pӻiub�'���e�'r�'��O2��5��� *XL�g��U�����,�M���?y�ā����<�~z`��:��+� Ϻ?��� E.���%�@!�ğd��П��I�?�'G�-V���ɠE̔agn�g�iM�	q"|�T�#g�LH1O>q���w�4x��3)�"&"�3!z���4�?���?Y����R��Is���'���	�}T����҆U�X�/__x11��$ H*��OX��O��D�*'8 PT�[8�t�2���I���l�ǟ�2��4����i�Op�O: x�E=`�8�EJ�N���Z'I}�-�?T2��O����OX���O ���g�zm����w����Ѣ]/i�R�pu�<!���?A�����?I��7�>I�*�`]���y�Xq��i��W\�'�R�'<�S�92o����T��%u�L��7!U�b ��sS�����D�OZ���O⟐���~R���-R�t��"ɗ#��L�1��[}�'��'��'�Pi��'~2�'	����ӏ8�����ĒbqR�D�j� ��9���O"��\90� i���x���0�Q���ã (�{��ܓ�M���?q,Ov�[��E�������\*��U� 6��)w)�!0��icI<���?�C�a���iߝ*�`���G O29�*�:O&�FU����-:�M�eR?e���?AX�O�DZf�*T>ޤ��׍>�Z]rb�i���'?��8�����: �xr@�Z�����B�#3�F��H�.6�Ov���O@�IE�џa��
*Iz��gl�w�����MSR��s���T���}z�1�EhF�`"1��|�xHo������̟�H���ē�?���~
� @X���u������X�v���d�Ą��1O��D�Ov��,TdQ�@ܗ
"�$�F�zʴImZk�C�M����?����?�V?A��/���h��'[�r��7I��-�]�'U�L��']r�'��'��'��OX�]��mZ��i�dԨP�D��t���z�����Ox�D�OPP�O���؟0�ģߢr�VL2�'��
��m ��е(�8��`��ȟ����\�I�����a��MSTn����y5d��0��\�*����'���'B�'$��ߟ��"o>�8�#J�.��g�{c>��5�?�Ms��?Y��?����?i���-0��&�'�r��f`����S)Y��5���7��O4���O�ʓ�?q�%��|Z���~��)���2뒀��D3��ۓ�M���?��?�2'V�V�'��'�D��(o��H����*_\쫁&%}86m�O�ʓ�?9��|�����4����7a�<�X�PS�dDgSxKݴ�?q��d�P�Pռi�r�'���OR��'!�eY7��2���H�)�cȨHa�>���h��K��?�.O�)9��	ܸxH�\X�JA1#4$�s����M�7 EVH���'���'��D�O���'��-5y�V��vb�I��c'����6m�!�L�D7�4�L������*f8j�b�&Ɯ�B�ݬ�B�m�� �I��X��M����?y���?I�Ӻ�D�Z-U�*���I�m:�"��A'����-f��?!���?�V�k@�E��ó!��)��R����'Q��Kt�6�D�O���OV��O���R_����e{�y������ɮ͞�	AyB�'��'B�'�-���^�֘@��ҵ`��d�\�66�O����ON���F�Q�������q�c�Y ��C%=]n� `�}�����8��ݟ\��Ο�	&4up9;شH��`��5m�"xttQAr,|����O����O��D�<���nj�ͧz��ҦX'��$��hwYs�#Ŋ���O����OT��O��`��u�Iȟli�ϓ�E�d]�����r<<�AG!�M����?������O ؙ"0�n�䰟(Pv�0m��\�l�3! ��y�&�D�O����ORixS�������<�I�?]Ae��8��5��-嶸���^��M������O��hE3�4���O`��vj�)�� rV�Q�,>�лa�r�L���O��I`e�Цy���\�	�?���ǟ`�t��e�`�BYyl��Ď�V���'R���t��'Fr[>������eƀG���Ru�> �����i�ZMa�u����O<�����i�O����O�}9�+j̰=�������"��=1�jZ�� �	qy�O��O�b�H5�h�ՂY%Z�P]`)+��6��OL�d�OX(	�E�٦�����D�Iӟ(�i�٫f�KB����� �|'kk�`�$�<)����<�O�2�'�rˋ<=}r�93�Q@�JMY��#�6��O�x�������ğ���ß�1����ɷC�8QhP�R�|W�`+��@�p�`^6���?����?I���?�-��9ِ�5;��s��k<��(V?F�-m�֟��	ş@�	���I�<��}�}r��T/���kDϋ���њ`����	�p�I՟��	O���M�]�6�]���U) �<j���Sd0L�0l�ğ��I៬��۟��'���D�����
�t ��AD:g��Dˇx�6M�OJ��O����O6�d<F��YmZ��	[z$�3j/P���)���$$��(��4�?a��?i+O����(��i�O��	�m@Ձ�nU& �H��cK�!<�7-�Oh���On���X�P=n���p�����F1�i#%Bȣ a��zu ��X�ٴ�?�+O��� �h���Oz��|nZ� 
��A�ܕ1:�}��FW)b�������'k�x@�	#qJ��&�0D�����]�SD�%v��H{��lݜ�q���	��1�N�N吠g)m��z�c��߀�*!��	�q�XP"�- �4��U+q��-z�O�&:8(��S��o1dŲ'+ݧa��� D�#�d�XW�P!o��ͺL���@�(I >��q���%�)�s�Gr�J�CS��(L�e��)I���-B6*���b��Y�9G��0҅ ,����
���\`A��,�c"X�aDE�$P6)#�Fԟ4��˟�����u��'GB���'�ԝV{�qvl�S�t-���6$۳�'�\D��,��Q��|����91���Cr��,�.�aE�k~�Hr0���d/����'�f�� ��-��hA���pX�'nll9��E�a{"i�%��ȶ�݆�<�i�\��yrkġd��s@�O���M���F$UH�#=�'��F��)�5�i�ܲĘcРP���q�d��c��O����O����(���O�"�l��J�K�� �k�?>�A2ԭ�!���R�&��a����	p�sb��x$�������(�x:�.�,�teaRDB�
azb�Y��?��n��t�R���B|�eQ5h����@���=��5d�����+>!*�Z��^:ؼ��ʜ�Y��T%7�*Q��b
9o� ����	hy"˟� 6�7��O��ĸ|�R.��p8΁��-˜d<DK�1 �R��?I��<��@1 ��(B^�������cz*��AD�%A�E���HX�����	iAܑ!G  <Q�H��3
�H+Z)y�EpA\�е�����x�ү&>��°��g�\%���B�O�E���	U��
��"�R�P����yB��'
;J��GՅ!7���,��0>A��x�m����h����+L��w�K3�y�B.
Y,6��O��Ŀ|
#ǖ�?i���?i򫐂|]�t�Cq�U3Q/��.�ԙ��Ș����9h������#���R�M���朻Mu����
� ����
�}%ޑ�3�ìM��h2�뚊C��d+�)���4�BɌ0��I�gNp��4D�숶
�-vD= ��ߟG$�X��7jt���'08V��HT*;i�͚3W�A�*�[���?��*�$w�a��?����?�#���4�̘a��S}2�`���8��*�Oj ��ǅO8�|�Β	� ��٠��٢F��Z��U���Mڱ{#j��P���3�n ��$@TR�3��X'A�b}�%�@��u��|�p(ÞY6F�HE@\�k,�أ�6D��&@�!L�8��s�ک,����I��HO>%�r�Z��M�6���z?�xw��gT���7�?���?���B�VH����?�O ��	��?	�(C\�����ڒW� �@c�{8���cȬ<�"�B�kM4LÓ͈u������{8��*��O��o�D !;)�?-�q�"څA�fC䉽�\dQq���#"�}�혷d��B䉾6Βmc�j̢���i�p�"�	���'�pxS6Bn� �d�O�ʧi�|��T���b,`@r�-K%�x�
�?y���?1$��Ea���UM��j���I�O����5GڻXU�pQ��)Q��8RĈy������3o3ƠI�.H�������0k���',Hk�������5H�	<ҧ/������KOƲ���E
�U+��ȓU�p<*�̊�l0LX��nK�b���I��r��um��>V��  �S$��͓^n�m��ir�'��S�O��T�����_|PɄ,ʵ?#�D��K7o��8i�AK�z����0�G�l/v��4,@����:���"ʡBV/V�A���ܐv�^Q�!�5-X�E�c�+�&�D�хRbąG��;�Y�k��3>���5Wf���A���?9ҳi8d�S��?��'Hqт�ej�Qƫc�tL*
�'DDL`�a��A��P���&��Y�����F�'���{0�d��"D�6PI��[T�@����?Y'�A��j�H��?����?yг�D�D�O=#5�{�0�@T�ªh�"��O�d���'�*�@��K��`��5 P�-��'��Mz	�+b�#ơҟ_2<A�D�-�����������=�f�Q��8��'�?%�B @���`�<�w�K!12� ���?A/ �b〚ȑ�"|ʓ�����f�0j��0��G�z,5�e.��#e��'Cr�'zT�S��'�22���!��'h"��-k]4]S%�P!pyB���U�p>���Fy�!&JPT8qv*�3f�IY����p>ae�۟@�� >C2���݈\�^�zvjD)!q�$$���	��?�ONX�����e�G%��!�f�
�')֔;���+�XYRRl�ީ8�'5~ꓹ�DDf�nZ�$�	s�Tj�0/C,ts��&I�>(i! B�q������'��'��y��_0'1O��0M(�XP#�>;zLuyF���b�Q�tP��<"��}▅�0;Ԡy�'�c����Ef�']�`����h�.��]%��$%ӕ��R"Or;d��C��0��U�]\���`�'R�O.D�&� !j5�ƣ'D�*B8O�)�c�����(�O��͊��'�r�'�$uӐ�G֖���'�'@� ׬�,;�z䱁�<�T>A�|��)E`�Ȱ��yx�Ti+L�j����[H@�L>E��R����Pf�S�y�G.��Mbxd"��?�Ƒ|���'�� ���J\��G�e(P�
�'�� J�DM�$�Y1�Y��_C���i���liqM��<�ƹ�����$i����Oarv(�/v:�$�O��z�V�u�Y�i�m�׉��0*��A��a�� S����(� 4�O�,Bh�B��U�4�/Ura���O ����'W0��K��% 4g�"t�a�';�\�����=Ia�C�Y�H�� aG����1T��iv�I�$��I�s�"�J���$�HO>����M�т�>3`�����&g�P�Iš�?)���?��KX�(����?	�O�`�����*+KX���B�#Pf,	���>5!�1	�i[hL��#�@�џ�)G��$+z��p�� y���R�	y��v�H�[ ���D*1��!�7i,�!Ҏ	�ɯ�M��G� � B�%*lᒳK�s�<����$U&ҭ��Q>+����f�n�<���R�D	p�pP��&J��\��F��<�c�$�/��mZ��|��A��b��XZ(��)�?@3�='-C,���'�2�'¼8�c�'1O�ӆU�4AA��N���gI[� �P�<1���_�O��0�1ă�{ߊUrkK�g�*����D�
�R�#�g�? �+R��'����˴U�D"OV�F�56><�FbZ�c�z耆�',OP]��#� `�����l� 6O�d�M���IϟؖO�4���'z��'4$�(%��H8p
��C��ٛB"�fy�@�N�0�� 9�O�E�링�Ͽ�pi�BJ^�K4̸,�D���Ć�
�&�r�bY5e/*�҈ٓG%�������1��C�PL m���w+X ?�p`������؟D��x�xuY��(�lu�g�֞G`�A̓�?)
�O<�5���+c�4ey��ڕ�0�Dx�-,ғ����n蜑b���{D��RS%L�`��$�O��0�ܺ X���O\�d�O�����?Q�]�@T8c�U�bP
I,��z��%��@�R����8;��!0j�!��Ĩ}
��I1k���]�=e�Q��
N�1#��I�˖�J��d�-Wt2j,lOI۷lXJ�4� �p�R��"O
����1,��U�5�N0\���X4J�S����H�o̦UR�F��5��U����)��I���������F�}�I�(Χ<�0�`d$�:/>s��Ѧj���BC��|���+�86u�m���2O|�A���?0�0d� ��5J��曚�X�s�L&~ �4�p��'�p<�#�����ڴ:o<|S1f <���#$Ɨ�J���T"P5�w�Ŕ. �A�b+��\�ȓt ��烍#(��1$��*�ϓ��O�d�.Цm������O�t�j+͞�� {g��Nޞ8���_00���'�A(~���T>�Y��0K.>��bm�pTe��,ʓp@D�$�̹�t��ŬD�7 d$2�!&�(O,q�g�'Y�>m�7o�>^\2�..N�D3��>D��� $_@μ S�K+�* +'�O�&�|�"oEB�]#iI�$��D!#{����%Y����O�˧}�����?���x�<bé:`�\`cR�T]��
.��9
�눪e�����)8��O�$�ХQ�h���g��,F�a���82�WǢ90.��K�g���'�pi�퓺wT��6�ևK\�gꗑ�B�x����䧵j*OV��CjG\��V
�9���`�"O&@@gP-��-AE�2x�Hp�P�ɶ�HOH�'�� �Ǖ���l�uk�
V��Hv�'M�iI1r��	��'l��'�Kg���ٟT g�diL�)��Y�ŔQ��M��<2�"�O$M�`^P
ND��k��uǈ8T�OD<33�'8��Su<a~��F�Р`�91�'��)��I�a{��ƍfb|$��im��ȣ�ł�yRo�7b(����^ J��j^�g
X"=E�d� c�7-ѯ:��*��#QV���"C(N����O��d�OJ��k�O��dc>��b$�O��N0�Y2q唶y"qy��	*a��|���ĥ8�8���J=t�h	��O��|R䗯�?���r�4]�&�!�L�7���0"O ��κq#�a�?ttIxd"O^�bw"0�zW�[�b� 1F5O��>!��
!ƛ��'��W>E�b�U��}�U�=�B��TL}@��I�����4l��%��]�S�4Ɠ�yb����$SgN8h�O�(O�<`w�6[\�QVhW�O\�(y�)�s�ڢ<�����D���>c�r�PQJK�GM �E���y���,xi��(�(3�����1�0>g�x�D�t�N���i�?[3t	�î��y2M��s��7�Oh�d�|"e�Ү�?1���?q��Q�FFr���MM�l*�����[??��uK������I�j1��+�,J5�$��'}�����`�����+��G���r�f��]��L: �̘{��'�d�O?����ctIy��1��]�1��.-!�dD��<��'�����l��N,�P���?i���.5���ib��}������ПH���(M�A����\�	�����6�u��y7IE0
#"��C�V$@�� �����~b$�j��CA7\Op�%f��~���ۅ�զ ��t1��OBp����z��ͅ뉘 �ʈH�(ّ.�����K�;�0���
t������M�R���,Oh��<u���4� x9��
Q;��{2�i�<���:i��`%L�_�V�;JС$���x�O�剿l���I>���ʐ�:|<�D�\�r���I՟��������A���`��ӟ���HR�;<R|�4�J�qC&�?7�"��3j�S�����	8aG5���2`^��cԃѿ?q�Ġ"`��]"L1ȡ� &qY}��a@U�'�r����?��%C�,�k!�f"2@ތQ�RO����O���S��� ���tkI6Q���g��R��EkB"O�}`��
�1�&5U��5��0� 6ORn��M#/OȔ����!�	��T�O;����~9��)�MI�k8̰Yr��l�2�'��"Ācx��U�HJ��Pp��O�S�5r��O(_lT@��%]\8�<�7N�P�2!6O.��N|2�E� Yu0E���1Z�"��D�'��I�X�>�����P�D��n̮v�d�q��<D���q��H��\�w��36H1���6�Oe&��{� ��0AL�eC
T#F�j!Gs�,)����M���?�.� ��Va�Or�d�O� &���em<��bڃ0��(�B�U~�xq���=9Gx�����#��OZ(�e��!i�IRBG4ߎ-;ѩE�nj��9Ѡ�4M�L����2��˔a���ϯ��o�-ӄ�i��'n��O?��TZ�f�1�B�%
���ҽ�
�!�DP� y��ů���� 
!�Lc�`2���?��$�C		;<m�$(��5$��!�ʟ����}]����������IџH�	�uw��y�]Na�U��h,QՔ�ks��-M�&ܱJ��	+dJ�/��`��O�@�<��M�h7f�ʑ��J�1t�R�.�C�'�3�((�so��Ad���?F�5a���B�6Ļ�O^�2jƜv��@"���pT��ө�Ol�aw�O�l=�M�gyr�'��Ɉ�d�����~luQ�	 ��B䉔8V"务˘J~]H��Z�^���r���H�:�p�$�<�G�*p�6��՛wI�u[2�i�$O����O|�$�O(�!��O*��k>�b^�'b61jR�B�O�j=�U �
Fu�Ȣ ��5���kzx����&�3:����g�9�%�ާh�D+׌=2J-fUjx�X��O�)n YB��WE�3_`��#wHęk6B��i��	iq�2#�5*­�=J\�B�	<L��A<D����j��f���I���'��)�3h�p�d�Oʧ8Q��횠b�|�� �R	�r��w���?A��?A0�JF
qI�ힲV��5�P���$ ��	uLX$�h�cJW�-LQ�X�Ѣܿ~
�	���|��Sm��L܅��	:q��u�7,��au~�ö��i�t$�T����p{R�s�F}m�ϟ �O!��IE�Z6	�R�K�,���#'�'t�O?�I�"T�H�@��=5A��A�I�,p���$�E�=1������8TYƸ#�i� J�0�	�NK�4�?�����l�pS�'|��'����ՀM~*���	6Y?����oiش���T-���e�O��J��8*�o͌^��i�RbXN�6b�#A�\�\�.����PU|��]wA�՚���������!�ت�pӱ,5L�gO�6(2�q(������R��#O�����L�Z��aRcH���y2@��	Hf9�ш�+QJ60 �/��OEz�O�В}�q�%Bޣf��,
��*y�'��p58v���'x��'��֝���"d�fɁ�M0Q7.�@�B�<V5:�{����Udއ[zBV��?�=� ��&KGB�H�"�RU����B�:�z��'GU�/^�QED;��' ��E�s��H��Ov��3�-7b���M�@�����Of�#�'��{��D����cS	 tf � �ˁ��y�Z ��`#ǚ�1R���� �Hf"=ͧ��!�AC׼i:|a�D��+U�6x�K�2p|��'	��'�r�G02�'��)'C�iH�+{Q��&I�dY�B����4�i��5���;QZX o@��Цi�Ekh,jäV1uz��d� [��)yw ʢL��R� D3x�qOb�KP�'} 6힅8���r�盛,�Te�o�{�!�D�&Ԉ�3�g��$��Mި]�!�V �2Ͱv�G�3d΁RbMڋ?�����$��K�����O��'(qP<g�ߓ<�p����J�p��Ɉ��?����?)�i˳�T�	����Ԙ� W�t����R���.Y�������<0���	t�
qղM`�hE7I�@zW%%0�j5�O "��Q�Ȏ�B��Pd^(	�!H��$ڂD��'�����j�>�f;�@C
D2��p�9O��$'�O�(�d�%^��$��OT�4ɠ�']FO�i���>�*���K$
6�3�;O�LX�m�n}"�'��S$-ЦE��ڟ����O/����G�d���Dx`Ƅ�h�>�AW�F�*X�̹�S�t��'v�y3���%Ar֔�b���6l��b�T/*C��
p�'����'��h*$��w^�)�%]�)d���QKH�Bcb�'��)���O�ʓKͺ�f���?����	�1ܤ��ȓH |[3��Y�b1���Q����Dx��)ғ���#n"�j�䉑�����I��$�P !���̟�IƟ��Zw���'���yBa�.!Lh�ІU{	� +�'���Qb�F�&�`\*�Õh��a�M������4/�ƉS2⤟d��A�ph�Y�'�ш&@ax���c6��)���16cl�s����~��M��?YT�i�87M5��4��i�i���T�&u
u�4R�e�!�� tU��� Cv&U#^03�tݲ���j�'�J�����Z�|Qm�?��i0aE���@S�%�m���	ȟ@�	�Pk�G�ϟ��	�|����e\Z`�R)P"lds��؆"��Xq���7}�\��c'K-��<�ĥ.N�t���X�2�2��5,�z���'�_��a�&�޻��<��'��p��4�J��V �0�������J1c��?���?���?���䧍?�w$���f���U�j�БB'ǀc�<3OI� ��i�6@
��iBd���<�Q���'"@�x��cӦ���O\˧���𳄗�GCp�;vO!;h�ݺ�����?)���?1�BѶ9	�0��y*�4([V��F4(�X�m�7j( S��ɣR#�(#u" ڧd F'\�V�
��B�8EyR
C��?9P�S�Z���H��6�M��!i+tB��5"��ԣ$�}X�йE'��Z�<��dR�	
���U�u�|!(e���Ɉ|��Sߴ�?�����J3��D�O�a^d�Q�M�];�Ԣ�o�L`h%�J�n�ҩ�G�&?�O�1��b �D$�q��hި��H��@�+-��+�ڒ���â��"~�	�'��!`DW�I(q�Y,F��C2��П0KL>E��v��$�@H�9κ��cA�.z�8���2�v1��n	�*��!�5Q�\@Dxl4�S�4S�$���N�><0<�˦�Ɵ,	B�'�4-*�/�&j���'���'7>ם���4Q~��e�^���*ԨlS��N"�Yir�A̪��C�?�=9�l�)@���u��A��c�DшD�"��1mD@}����M�)�g�'�Dсv�L"aK��a&ٽWt�X�'g	;�KÛ�&�D�OF���<���JVՊ��F�)/��e�E�<����/&�� F��7+f%�5A�Б�p�O��Ɉ���s�4���h��	�_�8�C�FK+����?���?Q�M�?1���dmK�?��d�B��s��n�ZL����|��ɪ_���P��d�X�
*�[s�ӛbӮ|��	Mo��d����q���'��T��?t�Y��%D��"5�t�y�Ȝ ��a1D��CQ�w���4[����ǁp�x��}2"�W�"6��O����|2�J��&�q#���&�}�]mn�0��?���h�U��������gg�����'A~��ag�˙*�Q��Сn<���JT�3hY�y �(WIMB"�EyR����?-̑>mP��%W��t��K�r~]Ȃ�+D�l��C�4i0�2S*�%޴t��d+�O��&�h3u��$����F�z�H�1Bu�$r��ҍ�M���?�/�l)���O��D�O �����8mT���M�,�Z��E	��Y�&BE�,�|Fx��w�tq�HΩL�<8T 8E���I�K�S��?���L�**���I�"duPlBTV�|^�40���?����?���'�B��A@�.�H���
@@��r�'��' �AJ�Ɇ'I�m�Ed�5F�D����o������J����m��+&�)���]�v�d�O��2����r���O:�D�O�-�;�?���r2B$â�1�J��!U27��'k��0�OY�W��Zp'����O��ec
�"�2i����)p��XCdq�<RQ��Nݘ�K�*�(��?a1CG�Ue�W�	�=�b5
��JD?a�(������D����%��� �0 �hC{C�B�	�C8�����5#�ܘ����_���Ë�ᓽ	�p0�4�H���C�$�T<�� ��yН���?���?yfm��?�����䗤U�F���De�ɻ� ǯ{�� �<P��\��I����bb o�  ;�Eg�
�W�D�-7���'�����h��ƭZ�\uhm�q�[O_�|��8�y�*Iq�"`1�F����j����yRO
A�<�4 �-F�r�¶�y�%<�I�n:�e�4�?Q����)ʒ"���Ҡ�CW����f���8r�L�O��d�O��8�,�#�TY���|�a ۑ<+����O9N_t5�_�'�@�b Y����iƠnF�D��	ko�`C7�)�Q��"��O>AG�t�A*��s�M,���ՈZ.�y�?H�x|�%XIVU��D4�0>�E�x"dW Ǵ%�u��8SBm��F���yrM	_s�7��O��D�|Z�*�?9��?A��ěL��U*V�^��Z�)�D�;���☧�ቪ=ƞ�Y @�p�D���
�ȩ�j�F����b�3I"\�J3i#:y���іj6>)�d�'���O?���:��HcC�4HM�0�@�߭�!��J�F+B�з)�<^ּ�Av	Ӿj���!���?� ��gA�3]�J�D/Gyzň1
�O~��� �P+G��O
�D�O���Fĺ��Ӽ%�Ӛ ��� �lS��p�K���P?)7�d��D�2LOR����ߤc�.)�� �&��5@S�A�(�jv
��=�p�!)W� ;��*j��O���e
%8��  `�`�|�#��O&��'b���G$\2�(�댵�DFUT`!��A�gHHA+EU�>�l�������Ez��	�.!� nT�!��/t�:͛e���m@���I���������ɟ����|��!�E�!q�����v�˂�Τ�<��PE�tg���CI
$��<ɢ��t	�A�@K��<(��L�u���HQ�A���@DL��
CD�I�B���$EƦ�A��E�3�1���5m� �#D��3�ө!] �b��~��r� "D�@�A$�60�,��̚>c�(�6kb����}�A
7&<7-�O����|�sI*s"����a]w�L�  ��$R��j��?��GNxh!%L=@Clӷ�qM]���]�T�.}�x��+G��t�*�K��(OJ0���7m��4��-G�,��y+b͢~"6�S`����H]�_�Aa��Av�'jd��h��	p�>>���`%8
�*�"OHɁ��D�b);`O�&o7���'�'��ON��i�� 3JԈ��)6#���t3O�� d�ͦ���ݟ��O�����'Dr�'�p�M��f$
0�F�>� B�=�D�1�J�#V��q�M��Wiv��'�Ͽ��${L@��dN&�Ɖ�E��{�-H�
;+�|�쑀y�����9���a�
��"��5p��O#h��Q�����U�I̟���ޟE���p��YёL��<���ʋ=U RM̓�?��?D\�˰e$NEFU���C;*��Dx��%�S���+-\)�t����*ț1�~R�'�(y�,Z&�2�'M��'�(�]����HX!�3�;�J1Z�C!'=���^��dh���m�13��X��A�!m�����['�}���SL�<a�	G�7��}ұ�J��~�g	3�?)��'6h�ʷ,�(e�81j҈��e�Plr�'�`lP-�<x)R������4�S�OG��[VOk�h��b�]
:<B�i�m��C�(��&��O��$�O����]�j���O��ӗu��]H�l�;�L��@�F��#5-K	kݪA��@J�?�P� �0�h��nE�__��(g`���Z����V�p�ґKc:͋c�'0�2��g���b 0G���4o��ox��7HǡH� "=����Ow��pbG´� h�Bgܓ �!�Q� �h��ˆN�.��5=&��'�J����X�YIX�n�՟���Z�T�У}<̠�u(P�Y��+�Bܦ89���w�'���':J���%1SZp�N��'u(�T�U�	�J8	w'؋\.-Dy��G(��FJ\P�O-@���AZ�n-68W�G8�9��dC�)��ӯ{�N��V#I�</(p��7G4B�	"��L��L�mB����9`���
p�	7P�`��c[;�����
�nT�	�z�E��4�?���)�,:���D�Ox�$��V��qA�`��D5�Pe�"<F��O�b��g�'�y�G(���B!����#[��� �Y�I��"~�	9��k�iϜ�(8�)œj2Pi�����H>E�����0cR�B"HaÐ��g�켇�gD�i��	�*�����猀R���Gx��.�S�4�� |��Y��<#�,���w���'�(H�2��|��'R�''����]�?U�#Vm�Vِ��6�!O��ɥ^\�d��i��Y�֥sg�'�R%*�{��3��4P�IR�.X��Y�ɏ�c�T4�'��,I���7OR�UD�d���;��^7@��=�ɏPDd����MP���,ON�Ħ<�ą�	'nd�p��� �F���c�<���VܒC��\��;שZ�H�������^xq���<)3@[�h�N	"`r��a�9O�P��r
�kN����ON��Ox��5�O���x>�±�O���$+��A����w��0�� �P-�|������D�܌i��t���%� ^(�|r`��?�!�i��h^�t�s��*tC`@1�D0�y"�[�����B=d�ZU[�f�5�yҫ��.+l�����[;����٢�yB-)���h��XC�O��ħ|JG��#]ZV=�f
E�<�(��D�v	����?��B���(l<!RuLK48yT6]>�á��
�l�P�`ȞX,��2Q�:ʓ:�L�b�=��qY��hB�'i�h��A�F�9��� �-(7~�5Gy��X��?qt�i�Zc?�k�*�9=a�pؕ��#�
����d���IDx��q�EK�	��y�s���2x�V� �O@�'�DA="(M��F�:h�2����{���F�٥�M��?i.�^�:��O����O� ��&�N� ��59�K�0�N�3`MH�_�&ty��Ҋc����R)Y$�V��%h ��c>�Ή�I?H��\$5��0�rO�.+����7X?�7'݆7<��f��h�~@+�5����ȟ����EHX�TC���f��)y����\J�)��d	�nXK�Li��@Ο#t�2��%D�d�%o�>���#��o�n#< �)��aȉ?�p3$oʔY岐�ǡ̏�?���aFp�ABF��?����?��Z��N�O�n�"f��r�B�g\����;j2�\(r�}�����)qT��1����"ۿ�~�����>����Cb��#
_�N�|P�	j?!R�ߟ���_�dx��,�U�AcK99�$e��7}�qPLeN�Aw�6(!��$�)§�V5S÷i��TX HKUt���iGt<�MK�'"�'��.2��'�Bd��'��a6!V�EtD��G�֝lh���
�xj1�'��	R�M�"� ����t{�\B
�����I��M�D�]^<���	�%��U��b�<�g�I�|�6�В�S0��Ac�K�^�<��.Z�'ں0�S�܏&��hd�Q�<�U��(;�n�l�ߟ��Il��J���������_��UC7�n����'�2�'!z��r�'�1O�ӆm�p0�f��;HH[��'e6`�<i���_�O������ɤFy�Mr��֍�d0����
����``Ȟ	8
��2,ŖHC�	(]b�L���߽G��(�*�:f/"����`�I��č0�Cͥ5�Ԍc⪌$Q�8��S��@R�4�?�����i��Cg���O���D�#��(�D��L��|�# �<i�nHBqm�Ob��g�'��M�� ���%��w��;�j�	n�"~��/e�ؕN�$Tд ��+|��Z�A͟�IM>E��H�� c�ŕ�$앳���!p�����)0ȝ#dw����)^!4	��Gxr�>�S�D�3V�j �1���J�}���U�rt2�'�ҘH��^�,���'���'���K6 ��G�L�BW�z쀽�a�r?�Vd[- �8��I�B":���/}����Ȯ%<j���tɤMb�i>|O���f�Q�h��Ai��ta�M�sj�O���OF���O�Y���INyB�F�"v,����.�"��5�E��y�iԛ-���0@���
R%ʛ�>`�"=A4
��Е'Vv@ѠIt��� O�/0x�6n�*)B��WL�P��֟�����������̧	F�ɺ����@X�Q"D�VA� |�ֹ�v��'bXه�ɯo�D;!��� L{�\�|($4k�b_�p+��a#*�/ ��DA����wӜ��raݱ%F��&��5	�j�"Of�#�'�|8���i�P+\��y�U�m6� ���ݜ�����D6�y�5��	�-K�OB���|bw����U���ۚL� �8�gMt7�(����?���[.�8�ń>��I�3#�A?�O�d)�'ɘf�����^�f5щ��$���(&��E�����*��\ ��W����Ą�(OF@x��'�T6��n�'j�P6>|sQg�)
��Zh�<y����>t��8\z
,���1���(�BQ{��[I<Y�`Cfd����<�Y[!S�<�Wǁ�)ϛf�'��\>�Y����� �����S`L��{�v䳠cF\Y�]q�й&�<9�	~�S����$���T��|v�l��Y�?#�8�G#�S��?a��":pJ��P�,���&�&���Iɧ��Bo� 4E�8�&*T.#��!c�aA8�yB��a�L�=���bÒ�O��Gzʟ��Dγiƈ$S��K
N9�T��Oh�$n ��w��O�D�Or��Vߺk�ӼK�o�*C� �R>Etp�sn�?!��ix���p��0�p(�d��%�B��"�����C/�O:<�F�:IdC�Ð+m�LUʰ�O�aHb�'^���� 0J@Ώ�)��/�7;3!��x����3:0��O�h1�<Gz��	��`:�lڧ9{�u!M��Z�z cׂ6ߘy��㟸����@E+X����|B���ԟP�IF�	R7���QXfT�Q�8����Tr���1v?��"ѮV�ptJtZ�a��Pf����A"b�}Ә�i��WPj�'T��t��3"O$T�b�7}�!�#�&]��ȓ6h����Y؄��&��X�@ıO�Q��P������O�q5M�
	�pX�C �Ɂ
�-W���'�cW���T>� y���"� ���.��WG��#��I��ƣH%[@z�r��;1��LU�'�Q���zA�>E��&1==�x2��H�l�8�e�-D�C���2,hJp�3��+u�xt3�J6�O�T$�p�Ш�{\XJ��N��]p�u��E�%�MS���?!-��|*3��O4���On�Y�둥A���!%5 �v���ʔE�^�7n�c��i�T���'�D����� mg`A�,��K���-"X�&������������N��<F��;b�azσ.��ԙj���(�b�a��Jm��HaӠ��:�t�E����-�$��br�C�V7����?��@��lbV�ו��gL��[Ҕ�Dx�}Ӣn�s�Ij��蛚Ai�hS�T�"��ZW�b>�'�x����3sDR�'	��'���ӟ|�	� ��Y��nR��k��{���/z��D(T�̼z�F)j��:���	<���Qa~��Ȼ<��=�q�E5x���#pA^^?I��Qϟ�;��sլ�N�����[;t��مȓ �Ztyb�ˈ,����b!�5Y�q��)�'6X��i}�pY�ȉ�_m@�ن�d~~���'�B�'��*I�\v��'D�i��T�^$��b�r�ф�]�C���Q���W�D�Xl'��	�l	����`�"�ŵf�8�32K�[��Qh��G9�����c�"U��8�M@FY4e��KB*«<�Z�sA�ś�?����?Y���?���?)J~��@
2��%P�|�'�10��ȓf��MPQ�U�HH��"�/u8�ϓ`��	Py`��+�7�O����|��R0~���#,��"<fNԐey�1���?Y�i���x�������1��9S#_����*75@Q�l*�b6�\ �Gn��>0LAr��Q^��UTbE;ҧ[��2��(I�XD�ͣV	@���?����C� ;��L� Ȇ)Kj�a��I��ē_��dKʯ5�1z��"]W�� C�Kӱi2�'��ӕl��	�|��"&���ð(K�z��`7�>��iZ�̐'�~��E����|"����8c�A3�j]S��a��YJhNĈC�/Q��0t� pF��S��?Yg�GcLty"�ț)s�U9�'^�uav���;Kɧ��rKH"�hQ�w��.j�%��b#�yb�U;M�FF�#���;�Ɣ��O eEzʟ�(aG�Y�7��ѣ�.ݍP��hGl�O���PW߮�Sf��O����O,�d�ͺc�Ӽ[�(��L�ƵE�l�B�c�V?q�dMIx����m���0'�,8#d����C�'�O�,H�gX�Z�Xpǃ�8Pd<���O,�2G�'�����JO�b��ܛHU@���ØQ�!�$�@h	�ebJP�X��c➗2��Ez��)ؚ���$Zl�nc�$ޞ7��#E��?���?��b��P���?q�O��h�	-_K�]�1D�g�B)�bK]�jx˃CV�-�����'����p�[/���i�AI�A�"+3��;MC"� &qVTzg�'M{��?��ރj��Ձ�݋'ꂹzҡ	��hO£?��/�%��swH׽���!Iw�<q�mA�Dα��T�\Թ��V�<���i�[��t�F��	�ON�'��	׈�G�z��� 0h\u@P��?���?��#X�0:񴎎����S���5�����Z�yt;���;�(O�2C�.�$q��'P�'G���ݼ ga'�p�~5Dyr�W��?�����O��(D��9)��C�Ğ�c�֍q�'���Dݦh��!�4h�;����C��0>�ғx��B=y`�y�j7"���3h��yr�ژ)#�6m�OF���|*�jϘ�?Q���?Aՠ��'F���Ë�2���Ǎ+\]$0��ɷ}Y�l��e�>�O�1���i/n�+����j�ͣbIO�!+��1e[�R��2���d}���'�L=b3BG�i��i
M�U���(#6��'��)��4�dEN�f�
f��@��C?�!��\�X.�¥3u P]� ���8���K��4�����md��	$�r���)�3�(B�'!v��2��M���� �б?�(C�
 ���B��KC�	����"2��B�I>:��iZ�(�Dʜ�7n�
72B�	�Q��b �W���aَF@>B��.@�쨒T�\�`�I6z2�B�ɳO=|�K����	����`�۝A��C�	�n�&����nBPXG�N�8�C�)� �=�VꛅH���	�x�ēc"O��J�^�S��
���.�(U"Oz1��M�)��Tv����a"O�!ؤ㝠0�(klا�\�R"O�L���5� ��q�N(��HA�"O<A+�%M]&�ˀ-̎h��h(�"OĀa� .I���N�fF�R�"O��[sNΝ]9�p��="��8�B"O �a�=������	���
�"O�|� ��7�*� �h�r	�dص"O����Y`t�ɕ�P���1�"O�����L�z	�	�!HՉ?�zɩ"O����씱'�fՃ��U�`�2�"OF0��k>;�t��n̼|�lpy6"Od�CEJZ �ˇLT�)�ܼ��"O��8�h��f�RhR�")<��)H�"O�,K��2R�D"�R�d�""O|�"q��&�t�V@��F�:�"O<��gAζi nQ�nϤmż�J�"O^9"�jG0�b(ӣ�|�F�s"Ob��q�� ���,n3F1x�����ti1M��5�ы-���u��@�Oa���b
19 �Ш/��W�٩
�'$U���6)F��C��co�SF�Ax�ph���{4,8��^���ء��'Ԓ���*H�!2��0"����	�'�����L�ؐ�Lɴ��̂�g�V�`a���ē[,���X�?	�lJ-�f��7>�ZcM �1�O.��4��G� "������C�f����Ƽ5�iC�	P9�B�h��4�VKZ�b�R$��hH.��	�B�\#+��$)R U<���ն����t����ML�fX(�s�O�?������<i��w������!j�ܠ��E\П����M}�$`(��F�UF���/�J�uҳDf?1&��Ŀ[�V�>-�a�^;	{�ѻ`H�,�Ԕ���ҢZ촑���O��VF]);�(�O�żCI��Htء`�z�����A�� u�$2�ɼ��
�,���&U�����-����@�	Zc"��0]��~&����Q�D:L���ƥx�,�3�d]�HO뮛�.	t�ȡ�=�<otX����kj�R�M�2	��X��N�o��?�CUK$�H�w�hCq��_t.(kPʆw�`��'����AF%l��'��~�U�F@PɩD@��n�z�s��Ϥ&<d�QM:���#��H�W��m]�� ��׿	�x�'�a�7@J!i�p!h�� B���O
h�@�9��Y�dw�O\�,��G
�[��� v�ٓk�%9���w�Q�q�
+"�<�"�J�3]��*������x����7���)8� ٣I�0��O����@�C��i��kl�A��b�1Oܳ�C�z:�zf�(0�����hO���Χ��	�c����O�a���"��)�$-��AS4_�� \kr���FC²�����ICs���^CvE��L�~i���[�1$^�%���Ig�X<G\��ǰ�`��_�TG��0�u�(�5E����f�*T�N����Y���'q�5{R$�PW� g+غ+P�8M<qCFR�wɐ��T.�� ��D�R�@�?yX+m�J�'�qGNB�7I���PV>7-x�U�FOI8��L�:g��4��V�*�г�D�XS�'nT���+d�5��B��6Mz�&�Bn�X�[!U\(� o¦#d���'\
�$?12#͚������y ,2�"��k�xu1'���O��C	�3������ifttb%MqU
a�:��Y���'�� )�P���#ǒ O�cEI3�:�����?����̀aԠB�F�����0K>�ۤ�ގ[�~���&?�X��n�	}f��ٴ����T���y��ή0~�j0	��9��Y��*���(s&�"hC8�s�jb�1��`��r��)��L��y/�X��=ғ�BђV �2zh\2���i�Q��!-��Pj#���<�vi�NBАR*�S�j����C��Cy,A2��ODv���J:y�(:��f�| �D��5�aެ�������9Z���B�єR��j��lhx��'*�T?AC�|��v��Q�T�]9#K�@x�B�,� }hD	��O�S�2Ɔ��t.��Mp�2i�84�� ��!�����͉�2��6�B�XZɋ;.Ռ&��1:3e�&�e�%�7

��ҧVn���$K}�|����9l�jD�2EͲ	:�7-Z�+��y�'\���A��lբeXu�	 0�]�JB�.��Y���o���@U�-󂣄/+N< ֙+�Ph
P�o�J��r@���6IB;��I��On�b�b��JަI*�c 9A�DU�Td�u��e����O�ܡ���-	�0��Jgұ4����� �H?�*A�p.̀�{*�"AAE�3�dmB��W�jX1(� Dz3M�t��1����<�O2&c��i̶n]2)w�J=U��)U���J��K����ʧ3��0�^��y�nJ�jԁIB"�����ծ�P�\(��'q4:̟���Z��>)�wH�d�6P�Ԏ��2Py�?n5��'m9��'�gj�����G����O���w�F�9x6QДeɁ{_���M�!��T	F�E�ٖ�n�{��ZП<�ӝou���O�ZE�S�? 2���;h�L\�m�%-MT���*���ԥ9Q��S�x�r�T?�aA[3d8�̻oN�b�������aR�Ȇf���If���	e��;fU�m�e�J�\�N�ʧZ�hd�R�!��9��H[D����G�p0�Y�#�<a�
�^���Pni�yy����i��F��e
��^8m�61�&�Y�F�6�j`CH�����'i�&���?��0
@��x���`�K!�/��(?��I%���J# ���ߠW����~���"��2@P�Jt�歍�<)6�hK��z��xJ?)�e��v�z��@���Si���'�?n}G�Z���'\%�"��n�8��v"]X����+���?K58#	��p�
��d0@h��'a����>�?q�o�F�$�ҏ�Q$c��TQ�%��9*��cO	j*D0�'�<m�Ui�?;�HQQ͟��|
�خC(�@�B��!b�p4IA��?9�ʛ!��&��I�� !ȵ?˓�0㖠�	5~X �A��23t4�d�.�:��=�O������⟪jԦ ���J��	�큻����Bi�K��8�̘"?Q�����g?ͻr12���ȟ�[Zf$ �h&h̓Y�x��mV"0^��S�n��2���y"�&ImrEH� ��Zz����Vx'�I7��2x�%�x�݋��5�֠�V�P&o=�!0m���uG`]�u���	���EI���Id��pK� �(�x�EN�4ʼ��@�J7��	�CV�d#�
�Ml���pK� �(�}�(�,_��,�#�L!C��1ǆS�@�91��zRȅ6LJ93�8�c�~�S�t��%��B0M9\�.�f��e��$. �4��U�C�$�� YR��50c��OZ\H�V$KJ�S"��st�
M�PEK�#�4#v��wqO��?Ub���*(�x�(d+Թ��fТw�R�k��Z.VĦ� �N��;*:G+D�"W�� �d$���<����y�[t^�ÓH�A'T4K�N�y��|	� pJU�$Y�U2�K0��'Q�ur��Zp��p���:�.��G�Њ1�U��G�t:��b�
M~�͟
iuR���5ZhX�)֒�~�ٓ��|���{�(�Tc��'�<��`ݗȘ'��h̵c:�̈"ouF��1�4��oH�a�&���`E�j�^=�I�[}�ue�VU�"�ųq'�ʧ�d
f��|��@A�m��B��8��'i&����6@S��kf��#8O~db�m�Oq�	��nżoq�<�cjαrz�i��ooV��=�O��=�gbޑ2�z�k�'�f��%�N�2��Xi�n�s�.(qQn�~�h*�ꅇrg�x�������y��a�Z�@��_�I�nMGB��5`�`�R�X�s���Ƥ0�Y�o��8��O�	u�	�<iR��{e6�����Wn�x��:I�ݣ@�ҏ�((�ឞ����F%�O,�ڄ���B���{��)�BܡDT�X��� 9,�&�Y� ��0���A�eˊ��ɢ<y�'��k�H�Oɰ("#��W�. �'wD،j���5FTAr� �H0rC�݈Fh��L$O�� ��w#������/��H�d�ʗG��Q���ONܒ@f�~�];�`��8����ĸiw�psE雃sqPq����g,~�0ӎ��3/�#>qt&
nrT�I/sm(y8�ڟT1cC�4�0.���X�J����� �N)�����a%�Xk��y����%ݠ5��7��6+-tͻ_�|:�F	�6a������Nf�4̓3�QhN{�5���\�F?�\��t�$�'��+t�̷���A��\,h�S�2'�0�f ۟h�S͚�9U�)qV�#-���aI���O��tE@�@B�9��;h�hţ�L��U��']~���'j�x����.d�ڼ�v�4�bQP�O7�����4�&���X]a��sr��n��gd�2�p<y��y�7�N�o5tTӒ�\�]��Y�U��.5K�O
]ءn���j�&�4�0C���RKѫ6��M+�`V2_&X� ���E-az2#�S,B��DC��V
^��W����|���ض?4t]��I�L�:y���_/����f}2����3��-�4��Hqs/V=N�P���Iٚ-
� �Dɺm��!
��4wwb���ĀL���[���o��z�!�;S�ð�����S$7&���5(x,b�{�_�eV��!͉9+f4��$�>��Un=\R��E|b͜�C��?O���ɕ.����SL�'�"T�ܭ�~��޿":�̆�	�p4,`u,�ؼ��b%4!���>�E��u�I3ғ�t9s&n[..MP�5C.�jh �'(�̘����4��Éq�$0I�O�[U$$�T�߶$4�b�Fs�'���f���dJ��҉�����ޞ9���%M ����	�1:��ɓk4 ���F��2���'ή�����7`����0�>��i�i���<z@5���7�xa�&�"�3扑J�p �)II_��'cU�9
��@ �����>�V��(,�4��,�j�*!4
�x�q&j &%��Ȇ�V�"�2A����<'"֢?��;�� �aQ���0�ϙB���L�/r��'�4�'�I��}�1*��p��4d^0r����)�H�'Y��ڃkM�as���@D�0QF���`��uRbe�j,^���"I�B�!	��	�ʬ�8F�ի|XP%KR@���s��N�,�ƕ���>�AZ���c?�0��$���� ºL��KQ�\v�L>!��E�C�L0��@,z��ӡ
�k�ɡ��MɣK.�ֽj�j��I��=Y�	�gpŋS�
l��S`o�U�uG�8%�Qb�n�_�S��<��!�'6y��A�,ڨH���:��IIJE���ɴ<0@��C�Y�x��@��%}��S�YJ���ƫ
���O�����$�f����D+͒P�	YVdT4#���`P<���[B�aK���b��!���l��Y@�Y�ABX�A
�X����(�<I�K�?��F�lkp8V�E�P^�e҆.FO?Y���H��i�(J�(���+#K��`�͓f
�e�F���r2�R�O�'�<��:��KS=v�J����À��	����{>4�aC��::�,,
a���}� ��'�����iPJ�*4��3�Z>isd�j���"N)h��J�O��%�H�%J�
|�qO��i$� J٣���Tu����L BQ��T�����4�eE|������7�G�vj�� 	 �=J�h�B�?��(M�O�I�O�7�T�W��ј��ɬx2���(YK��M�Ƃ�^j,�E|�Q&$ifL�I��Y��C���y���%/����6H�G/�����hO�d�v�[�3������+)�}���O�AL��r�aѠ�+���j�>Od�d#�:V��� EEO�f��C�Dm���fC�	K��O�;�>H�L�O�}��L�>1|�'�!K���b��Jք`q�n�t'1	�K�)QmHɢ`E6n�G|�o�=@���rSkXO^�Ń�(��s~��P��L؞$�v6���(����ILL0f5bI�J�^��Jϓd�t$RCfWDa� JFiA�j��TH�/��p�	�ɸ�
A [���V��[���kq�����aF{�жfm����svZ�+�#��~�(
��Ȇ�ɚ#yشCpL ��O$AE˂[Y�4[w,�6���%8O��!��C�8i�h�|њ�P �'� �;�c��F����	)E���#��$̜^��`A���%��	%�R�f���64�AXֈ޿�,�kr$ܼp��(��?Y�QI5�Ŀ66 �����R� ��A�'��N�5lC<�pN@<����S.Y*v�}R&I
V�4]�2�����׫�R$����:$ڑ��tf�%vɒ&�L�d�� �R�n�H��+٠FW�ti'm��*Q��:���'R��H2���q��HY4�Z4&*��I/*�8����^�49Y�D420�o%��X��٢���!�7U��Ezb�ܽ2n|�R����1�t��>�M�SΝ�ܪ�@�H�&n�ң�DY�'���5D� ��z�"D.I��AA��41��<\OdQPƬFf	�ś��Q�*�"ubڧI���#�'��!`8/[�}s4�B�[��ŕ�B�X�?a���:=rLY��6�
�`��66z��Ei�8+��5Q���=]ne���D�
��XC�����h�v#[K=�'�/�����Z "����n&��$��&0m�){m�a�/�[=����J b]���O��vKӢ
����¨֓k��,C�Z��02K�Ϯ P��g4��а�2ʓ�f�`�VS����Ã	؜���g�H�l�2!`p��X:�	���0<Ib�CeШ�8ř�Ur6�Љ�g�'�:�����XJ�P�u
�	+�m��?Q�QЊV �x1�/N�]
��ޜNm�(�'���`�7n�ix���<L"�T��J�0H�vy�r���g���� �\+�}�݂ss�����_�]	�����R���B�`3r]��bY7�1Kc��B䉑p�-���YZ����#xz�B�	�^��%�D�O�6)BÀM�d�C䉷3M���g�O�EN)0f�L�m��C�>@W�|HfoEMHF�[7/	�2�B��-v�
��U *3"��4�>�B䉽�@�R�Q1H��x �DƎH�C�I�+��PS�Ɂ�;��K�A:#�TC�	%N�\��JnZ6����^	|DC�I��@`��ԅC�hY�W�#C�	8~��TӰ��1X��#��Ք0)>C�Ie����ღ��@�fɈ6P�C�Ir^���A�<F��ЪH�E�B�I\00 ���^*��u�(.B�>*�|͒b%/i��}�q؂,��B�	� wt�r�K'ᜍ�uǖ>	��B��)R\&���X?�DQ��'�>0jB�Iz���t�۰0�M�o���jB�3X�&�@p�V���D S�F�C�I$�.����S�5���I�P)0J�C�I�f�ޅ#�DA�x�g�>�!�D��� �6�Г/ ��j�E[�B�!��]=.M:���ʴ+>-��>l�!��םtS`�I��'v6���E�,a�!�X��A��D!�� Q"�V�!�d�#�,�avB�0EX\2U�@�!�dY�]��L /R�@�&�	f�!�� ��� ����~'�	��8�B�'���Z��'���I�Wx-s�'�~����% �h�P�,��]	�'p@1���ê`�и��U~�$���'� �1�E� �V�·Đz]^H@�'�6]�L8a�ԁb6�֙qM��0��� ��(�jI�2��lӜ?��L�"OHEj'��$d����:BE��A�"O����80l�RI�T)*�	�'A=B\�5��pX������'�Q�$�5<z�9��"ս@W�q8�' FYJC*� av�!T���H��a	�'�L|@�ߵK�xtbD'I�'rL� ��4��E�&OG�,�.�r�'2�thf��&U�`HC�nXB
1��'�&�2�ßm
��т�@�L����'",H�����I��Q��k�p�"�'[���K�欢Ac/o��@�'g
�B� V#2�R�j��n�(D+�'��Q��d�`z���ͼN&(�	�']x ��rDn����~�ƅ3
�'I�1j��A#|��!/��qȔ��
�'�Ȝ��ԸbOx�!�$v"��:
�'�0�{GF��]걐���eZ��x�'���R�T��~M2�ŋ$'�����'V��A$]�_�z0�Q��##��	�'�x���О{��1Q��ѠGP ��'��%	��B�spy�"���8�^���'���A��Y~�����$��3�T�yR*�Ee�E�5�IR��"�K��y")�):��8�F�Y��8�h�E���y2AP���u���P�V.)�yB�?��@��%�~8��&k���(O>��D
��b��o�0Y�V���u~!���7/�(*vh��M�Xt;��_�F5�)mZ[(<qW�K�
F��a�	�D�4͚0	K�<��ښ8z�X����_|�C!D�<��$��H���������!�u�<���M�/����+�dS�,�n�<I��ݿ=7��Ђ��VN8$EH�m�<�gh[b6<ӰgL�(�2,I�A�<I�a�X�T�C�Ve���Z0B{<Q�!Γ1���b1b~!��i�OJB�ȓtA $�Ì��RϤ��$���t��>A'�)�SⓙwU�U	@(#K�(���1�B䉏4�~��mV�C�։:wƀ#ian�Oj�$+LO&�3�!�*/���ᓊ��QT�Z�O�i W蘻]���Q3m7��y�V�FG�<�!I/3D��l�0H3��S�.Un�<!�n^�+X�����0�3r��m�<Q�-��m"R�O?9@��[q��S�<�����(��ҹ�xQ�`d�f�<��D�%�`�p�Aڦ�8�I�f�<���C�	��)���ڌ��Zn�i���O�4�#�E���K6 I����?���"�O"E�� _�|�|LXc� �*�)%�iűO|�|:�A�
$;���'6%����	+T�ĪaOΟG)���
�'.8Pj��P�sd\>�h%�R�DV�rX�!�Ӫt8F���L�T03�Ξ����$9�	!0���3���*�&����|�C�	$dr�A�+t����P$�UX�>���I.ɂx��&�� y�L�vbۜa%!��j�A`v�o2\2AO7�`�=ͧ�hOR�R� �U���ZѦ�7KZA��"O0�X0/�qYjG��XD�s4�>Aߴ�O,c��;��Q�$Tޕ���Z;GlL���"4�H0Iֲ�Z$�'eG�"�h���C�	j�����=Dl���)���Bٸ��:��hO�Ө#� �w�@�[K�h��x���	�ΞIA0$�2�HF�S�W���'�	b�)��O� ��@� n�r@ХB������"Od8�d�J�U�LIx� ɇMԢ!z��'1!�Đ�u���bf�$fy���
W6!�d�*U�̅�����.u�`AU,h2!��01�l���a�<����	!1O���dٟw�P�72J�y寏�!���DXX���f��x�<@d��7I|̡�4�"D���6��$}8���Y��k�灣kK��dZ�^u��cM�b/��`I'!��K|^�9��C?(��RҤ��!�Ć�*���PdiE�d,�4�G**�!��[_�;EaZ��Z�j�K�!�D�+��q[�M�8Q�%�͐OF!��؏k��٣��"�e!f�BD!�Ę�!*���1Z�0[Alȍ8�LB�I�l����Ɂ^l���2gO�[2D�OF�$I��<Q���&iJ҂Pl89�C�<���K�*�� e!�)w���Dߴ�!�DR���lY1�R<V��d�îޒg�!��J
4]��ț,w�'��"O����	�y��Q���H���h�"O�Zbi�(�
E1��֐T����@"O��X
����6"��,�K&"OPx�l�l���� ]�9�9�"O� {�.��`�% �m���v`���	T����[�s��4��o���1��ٲr�!��H�8>�X��_6c�&���IۏKp�ڰ>��ߵ�d9�(�+��p2�"@�9��O���<�u6`T(K���w޼@RŚN����'F���F�'nۂ��^)G�&PX	�'TD�
�M6s��%#�	Ƶ@��$����MG�Ob�<@D�h���B�eϜ3�`��'���T$�$��U���+�Y�'�ў�}�b�?q���+S,����e��T�<Iw��j�܅
�KY>�F�c�K����'/��2q,�"Ieܸ��+z2�	�'�(1�5Ě��}碑��[8�"B�5w��9�㐷ky(Q��m[> ��d�<)#Q�N4�2H�9H�~$��/�B�<�p�F�!*@�+K��!�����D{��)�)I�
ՉBo��z	B,�wUC�%&���(�:ew>iZKT2R��B�I")�x�E�l;����\|C䉣S],��@Dҿ>�ִ	b�)�C䉺+a��d`�.WEޕ+%f�<M�B�	�=���Ά�^�qg�W=�B�ɴb#��2���-K���j�ѣfk�B�	�g�2��J�&l�8�P v�B䉔W�L��50�L������C�	4�|��!Lm>��*�\0 c��<�I�i�x��po^'�)�v���b�B�I�?J��𲂆���P�Bgv��B�	�W �"�$f�����E�:�΢=	Ó1�^�J��n��T	�aވ-����'�ў"}jBN�U�jC�Y�,\��Cz�<�T�X-x8U��C
5���*��ry���_�11byʢEpF�ɕgY�^$�ȓ6�x]���S�Rd�G_�<� GB�u)�Io_�=�Sl�1e��B䉄KF�IPG�?�(d80��D�z�<I˓=�����Cİ	��l	��d��Dy��'K��#�@�	��YȢ+F�N��,z�'��-G>`-ڱ!!�3/����'�j�' L�%�䀨����'�
��� &�Ci��G�N}�kخ!0(̓�"O۠���9�߬q(��:�"Or�!`.L2�(��k�}U��"O쨘A��?����/)��j6"O�):�o�~�b=Q�lM%7�l Z�"OD���k��Z�2���jͰt��8�F"O��[�ɛ:� T��dU�3cJx	@"O�1�f��o�� 
�0�а�"O$X#��מQ.�a� 윉Ff"O�Dp����9^.�����O��@�"O��e蔰[�4ܱ��T9 ���g"O�a@6!�����iW�C�~�$"OΑs��!0��hǦ��Y<e��"O>�P�C"p��<����0iv����"O����֎0d1�dՃ7��Ř"O4Y�įn�H8A"��(��l�!"OH}�C@E&8�D��NE"Dj ���|��-|On��BU/0��@�_1Vz��$"OZ�yrD<ͮ�8d�G�T"OԹ[ A�/R��ųB�\C쩠�x��D+�	$��`&Nʐ��˅�\�����',,��eK�y�E���CS�@��'�j�ؤg�,;m�i���?�$����,�d6�)G#��*��	*���Cd�5`m��C���B�&Dj�c$:@�
�,D�l��iX�>�m���$%��i�6�x����a�6,�G��8��b���y2KԬLW 1��ͰiE�Ӏܮ�y���2Oμ��	�O��l�1kT�y2ք$�K7�y�TL1���yR�]/1?H�:pA@�r�|��p&�,�y�@�?uM޸y���!3a�`IZ �p>1H<�w.�=m���)�
f�Ш��MET�<��'˶Q׎Ѱ��
<��st�Aj�<I��%�� �D�9���T.SM�<�U ��s��=!�7`,@�Vc�<�"dZ2�TݓA�6��Cc*f�<)��56���ŋ�1$�Ũ�^�<�$,5,�t	d��%�9��KY�<ѨR1R	$�S�����e���^�<Y#���%�f��;K��]��B�X�<�cK�8�rY�W�WҼբG�j�<�5\�|T,�cώ	9������]�<�OB9�v��\�pR��<>!�D�A����Sx��p����4!�$�$±�fC6M��e�X�E"!�d��P�phht�K=5�h�r��$>g!�dݎN�QȒ*+z�丂�K�9X!�S�F(r����̂��EΟK;!��tl
YjQ+�9Y"�9*"e�{�!�17�,IB҅� U�h�i�*+-�!�\l��0����8���o�"1�!�$�R3b5�$��5׌(��J�!�$ڵ4�Z�X�r_�X"��?%�!�DZ"_��L[��O�$
�n�=[u!���:�ЌS��!��ѳFh��we!�dQ��CQFM�|wfa�#fR!�)��%��c�}v�ň�R�?!��Nn��h�o`ĵ���P;!�dR�t6���B�ƃW``񵡐)�!��&#4m)�Iya�e����$-�!��ݺZq�QK��� sB���$j�-#�!��ʭ;y����1!T �1����!�d	&$敉EK�<C@�phצ϶Y�!�� l=���Ӏ�(M!���
L��\��"OҌhw���j�&U�m!�"OmbCF՞>��z�HD+W����g"O8���Ɋ8	̠�� )%�
�jd"O�{�ʌ<�L���D����
�"O��HW/Q��
*�U�*`�"O4�)d��9�����$@�~���W"O�B��:"�^��0�Ƭl����"OV5h�'�-o�9҆!���0��"O*d����e��p�&��,|���U"OTl� �6*	�8A4OȴE�RLY�"O��I�H�9(�`1��L�Oz���"O�8�B�Zmt����ʇ9x�# "OzŹ��8D��Q�*U�S��p��"O2ػ�EE�
�!B��_�A2P�k�"O��AS@G�?��kI�D$*�C�"O��Qt�[��z��d'Hl���"OZ V���=�����G�"<���s"OڤI�!X�O��I��]_�8}q�"O��B��Y 7,���Z�
Ku2�"O��Ā<'HIg�@�?���q"O ��fE�)<�Z�۲�(}����"O���!�t�ZG�_?�@�p"O\9�mD�B������$�eZf"OX��C�2���`w��p�"O�9���#b���9�L^�f�5�S"O�UYd*��>S��0!�ٰy%�0j�"O��!c;.ȎqAu�]�$���"O6h���&N�����,).M��"O4���L���Y���p@K!"O옑��B�B���hw�!��eB�"Otd��`ұx�Ese� �cۂBv"O��Q�&&9�68�j�<k�P��"O,X����>�Z�ه���%��"OJE�6��<��DC,�6����"O�T�0ɅkPJI� +G�Hj�ibw"O�ͫ0�ƒk6D�xCJ^aNp���"O���+M���� G��e6^�Q�"O�e��l<HgL��ԆN^	��)"Ony2c�˂HC���u�����"O�BU�ɓ��D""�~�&F��yR!C�t��0�A`����y�BA��y��J�5�5��5�j����y"��I�(9S ޿p�5�Ƈ���yr��<�u�B�����.��y���#������{�jY�͍��y�jC/jt��T`��m��� Z��yBO�06L 0ϟ97D.�VH��y�B״G'��FGĖYث���yL��}j�U�a�A]����NR��y%V,.�<0�6a	9&%�쪧"L��y�I�L,�����6k��H`" �"�y�'�N��U���q3������%�y2Eؗ1=�`�F4a���⬔�yf�,6�4\���ƣ]ψ� ����yR��!b�օ�t\�[�Ai'@���y��%:���۔Qj��I�A�?�yr�8VF�ɡ�W.MqB ̠�y�	�[fP��l����X����y�ǌ�j�H�RWT'F*tcaK��ybf[ e�>�� ��@��j5�ʮ�y�V�95~(a ��'3��lqA�Q��y�ӤF<tXI7�Y!8���+1.�;�ybE�z�b�%�?(��u��b��y
� $]u�	-R�h�0C�P���"O^����^X@�a�E'�$Xr"O�֣� ���S%jB�S"Opl�N	�����N��{�Đ�"Or�$�ʟS4�uӎi�:Љ�"O��
��+I����G)4t�Mr�"O�Y�&�2?r����I)<��Mr�"Ol]�ꗢ5s�� �- 3g�&�XB"O��:7�^�P!T!)-J�wVq"O@t@1
Z:G�
��V��{�R�"Op]@��q�!��@<c�ʌ�b"OH�D̷����E Db��@�/D���#X�ERR���8�}�#�.D���a-�.$�TCǢݍl ��bA(D� 2Ai@Sa�p9���0D�A�H"D�@B��Q��u�Y
#Q����!D��)��L�l�*L��NC)G�`��K*D���Sgm�0lP��^�܀�n(D�
�D�Nn 9�3�F5<��D&D�����,a�ޕ��j��;��p��O0D��p�)wQ���S/ֵs�H�W� D��H�i²餙��B�F�Xі*?D�����>p&5b6O_s�����)D��Y"���T#��'�O2!�f�;�#D��C^9��T�F2I��t���"D��{c�؇.��[EB%-�T��!!D��dM�&*�-�SgF>mi�9uE2D��PU��Yn��`*�!eF���$=D�|J���d�r9+�M���
�[�)'D��4x�x��0c�/k�u;f�:D��	�G@�L, �i�N�]����V�$D�������P1��l�1b��fe7D���fL6DD���d��-�Lœ��5D��C��� f
���^�O�����)D���u㟔0)R�I�C`�41�g)D�\)���3<�,��D+I��Hڣ�%D���ߢW��R3�M��,1&"D�T�Ʉ�hk��j� �=	b`rf>D���B�dl�S���a�n����6D�D��X�}�"�R �ȉ#P��H5D��2�\�7��r�1��R�L-D� ��勐Rb�jEʅ	F�� ` d&D�<R�䛯`��X�e��&uʄ���&D��j�`��qfI	OM�l��"D��Y��M".�D�� I	�h���+D�0L�6#�q���ȟDh��i�D)D�Ly �ҟ"SB�O�iԱ"�"D�VCL~� �A�; ����c\��y2�V�T8�MSfA�"cFb�`�OU�y�,մ=�x�ka��+W��dX��y'��L�+�.J�P6��(�Iֻ�y� �0<��/�J�|�1b֊�y���A�2���
.��+���:�y��-)JԈ���Q#�pZQ�ƍ�yR���.�֬P��[�Ex���	�yb�D6qPD��e�=��}����y2�������1�4�J�	BH�<A1�`��02�r��l�$��D�<�$a�JhkG�|c�����u�<T-�J>"A ���#�(`��w�<��)�R��ʕ�E��-a3	l�<�*ґ#�Xɰt�X�y��A3��f�<i���+��8��i��Z5�p��@h�<Q��UYWJH��R�b��`y��V\�<� Ȩ�pG�j�°I̢]����"O��#��[�.B�]���ʽ\�����"O���p���G	���+�"O�P��nL�A�Ȁ�Ŕ���v"Oz�!i��	��,�5S�\��}��"O�IG��KN`C�@�Fj|5��"O��!�(�>Yl��(��S�y+"O�0�`� 2>�c�kU?2�@��"O�0'���A���0{Д�{�"OI��F�[��9R���Y��PB"Od��a	�0�MI��L�`����7"OZ����	"GM����
YQ��)'"O.�؄��%�&���i��,�pD�F"O�\@�'�#z@��{�(��_��@"D"O���5fK!�҅�6��2�N`CG"Op4A�.I��`j�iÓ2�����"OH�FL�pNz�QK ,<�@\qE"O*m@V��0�RD���5\̺P�"O�c�FO�"����
���+�"Ot|�7�A��G��;l� �q"O��K���z�jL�Ć�%���f"O<�! (E�K��qpHX�J����\�<�sI�v�|���S��(%�RN�<���Ip�cj��:�@� -CL�<��FC8_�Z�`��S������O�<Y�����t��K����� &NE�<y��*^�^���HN,;�	Q���V�<�ӣ�(I�J�����}���b�^�<	�E��FR�@2,N�m�p��@Y�<	�_0H�H�4OG�#�=0�Z�<apG¸%cp��$��7����2D�K�<YVʛK=��ɑ��6[k�P�v��p�<q�JKڶD��%�q~:�Z���U�<ɣǟ��^�� ƁQ�va�sǊ|�<��Gӂf7X�k�Ν������y�<y4�� [���A�9�!R�O�<�P�p]Ҩ3M�����ZL�<������0��,�Dq"��<�_����#S�.�~��*F���Y�ȓ`=�������}v�x:)R�F�\8�ȓ?\N�˔څ%�i�4D&�`���}:�$h�M_&��aj�Y�h������u��m�*�Ru�Q��	z��0��zS�ɉB���/t<!V�I�Ts����h��!��˖h��8цk�v>�ȓAY@$�ѠI!8Prh� V4TBȇȓG������!H.ؘV#X/=���$/���W��%w�$�&I�v��@��|�r%J��_�mw`�H�!?u}�=�ȓ=t��q�%�r@�HP�԰V�ڴ�ȓw�b|�Ԁt3&ʦ.Z#v�D��r�Z�@R+\�XD\�Q#@�SU���5�40΀�'���*���	���[�r2r���}�ށǫT�DښE�ȓI����i�b�,x��ʼd����ȓR�a��d�*
�JUZ�)�`@�a�ȓz����lW$~����mʐA\D�ȓs ]#�`�<�45�G�2e���ȓN������W�x��B�6Q,���ȓ�B��.��L�X�Q�0g��\���6�b��x.4A��S12|���d�|	Q��1(і���猆/�*��ȓ,8�Ш�̝� R
�PkJe.���+<�e���]�w����iʯKqfH��S�? �-i�N)��R�&\&-�x�v"Oڹv
��h K�F�3B�4��"O>��AT�S��1%M�.�<�y�"O�`8��\�QWeT1o�@��3"Oz���ښiH��c��.�j��"O�����8�b�prG��d{F��6"O�R[8�b�Yakr�����N�!�=R�d����
BF@��N��=�!�D�n�4��5�ر 8��9e��9{�!��҄{#�q�",Z�@K�H�v�D��!�ǯ`�ȥY�+X�tUL)b/��A7!�DL ����B	�5� ir��M�!��A�a���b����-��)r!�X4qL�+�図<�t��abʕu�!�.�H�uE�2g�)1�J�8B�!���n-b��	�,g�N���'3m�!�Dٿ���b�o����a'f^?A�!�$��8B̫a�.As��se	;}!�N_�TQ�!���L��D�?d!�dB:Mu�1����RU��YUFδ3!���4d�x�.Y`R��$¼j�!�_<Vr�QZ��.|Tf8�Ď�|�!�d�$s�4lxr�X 4J<��`��S[!�+2'�@�3ɏ"6X�Y�_�jT!��@�e���+��5Jц
�d`!�d��2�f9b� &z��s)�8 A!�DǮ�VMܡji��+�iR�G)!�$�.�aѧ��#�\�Іo� !�X 5U
��P�RG�~�!DN=P�!�dRo"B���`@�<� �g�\�!���7Ro��	X�4�ԢݟM�!�d�'�x�a�A,icf��2�پ{�!�dμz�VtQt�C�y�8�E�S�!�$׽>{�|���kd��a�j��!�Ć�rLr����4�j�V'��!��eƠ� C��E�2%���C�U�!�$^�\x���բ#��&�� �!�	k�P�h�N����XQ�%ʖb/!�N �@�a�@�.-�s�"[(!�dA/x��dvMEn�L8+���I!�D۝Z`0�+�`]�<��`�L
I�!�$I�2�|�dmW�J����,K�,!�$	
ZQ�UX�g�+q�.�B�§<�!�
�g���uK�d"��y�
V�O�!�F4cY��[d���S c��!�d�f���'r��Ad�I�!�ė #���eC�p]8#�M�!��:C� j���9��%�a�Ku�!��{��y�4f��DIPP���{�!�DX�#�L��k5F�L`�ǈ�l?!�d?S`$�B(���(�-~�!�D!"�FA��ցA��Xr�_�!�DŹ9�$McL��$�<0�d��9�!�$�+-��qIW� zؤ@d�.!�d̜�$h` �+H��pS�#_|
!���*5�A��+�@�� Z� !�D��	-��aQ? �&�9BP/^�!��N�
ђI! n��B�,�7�݇*F!�D/Ƭm���5u�)cC�W1!�_�s�u���U8��=�̒�!���5�RdSb'�X0\!�0))���:w�)퇪$/!򄙶$��i&�	/M���cQ"ӞI@!���*�������Y�S�ۂK7!�� ���#/ ��)��4z��Y�"O�	Y�
ҶE��� <6�9�"O2�� ��Ϩ�q�H" -
��"O��9�A�q�⁁q���Hf�+ "OB`B%���;Q�����&#�Hm��"OZɺd�,/llx���8m�"H��"Ov�Bb�/2�	p�I�>�j�H�"O4����;o��
���2d��3�"O� �%�H���e
�X}.�Kw"O]�ǋn�L��%\�<?`��"Ot��Qj[�Fm$e�+5m����"O�P��C&c�@��7�Js�:!H3"Oft�T�B+C{���X�d�Ƞ+�"O���Xh�)�uCۃ^���!�"Of����� >b��:�L�{�"Ot0�Ǜ{�ܵ	� ��^��P�v"O�"d�ܖQy*��ރJZ�`"O�u�t�L�6Q v�"r!,�"O�M(F�Y�@bЏ�-��H�"O�dZ�l�����eNǹD�� ۆ"O8+U� 42����r���"O��YM��|�n6��Z�5!#�>D�\�%g�>�eSqS�	�"D�8Ё���;ҁ��GȌg�`A���?D�Liw�ˈyN�)�Y#�>e��)D���d�ѝU#�Ը���]2X�@�N&D�På��<X��h�	<8�8 �P�$D���E���(��F�LX
0�
#D�P��HH�
��sΗ�Vء w�%D����9f9�A�x�f��&J(D���Ţ�=udȀ�p%@�fs�s�'D��#��ۍp����n�73�i�Vf9D��Q�����%�1��+�� �2D��
��O�2�8Bʛ)< �1eF/D�l!���
�ЕoT�g��P�r#!D�s��	
(à�M�Z��h��>D�@�w"ֻfe�
� ��@Qc�&D�T��j��Tq8�h@�	(4���� D�`ᴠZ�5H��-�HΌ ¥�;D���%�ڲ�`$e;l�R�C�;D�h�Ԥ�!T
�h#Q#A�J��U�7D��9GG
{8�aӉ�
(�ޕ�q.(D��*pT"}�iSuˏ7f�|1�"D�piG	����'��*� �{p�5D��##��7M�I)���+Vg@3��4D���g��l�*��󯈎v/���.4D�8:2n�����;Y�`Ӌ0D��)��N�8�p�тM��Q�`�.D���J?(�L�� �Y�$M��+D���n�%R�"�HVe��`:"�#�4D�d��H�o\~A+P�Y���`Y��1D�d��T�W�H����6���7�<D�t2qK�d)Xu�A��bڮ5��i9D�p��������㋧qx��'�<D�xI���/V$�����3�ܣ��<D�ؙ�M�2k3z��Bh��8.��C��<U��dJ	+>�� ��$�B䉹}�R9p��@9P�zQ9��6]�B�	�@�8���5RTq�V��&4xB�I�. J$P5
�KB>!Y���mPvB��?�  �hG6pt8Y�MЛ"E`B�I�YR�q�tK.U���qq !"O�U�uo�3�"��W�E��v"OZP�$�w�B��^9�^U��"O� *%�1f�n����⌒msX��P"OL��u��#�����"3b 
Q"O"����*#���5�H,-
�"Ox��6��q���",��2�"O�HX���02zA���I� +<��s"Oh�@�Kf�(Y�O͎Wh��"O:�)#���H�/��W�>Y��"Ob�k@f��}+�1饎׆���"OZA8(�*f�ȱ;5�ߎ4��<�q"OJ(��j9%����A�6攭�"O8�XB���M<,yk��Y���=h#"O0@gEV�B���y�/ì�r�p"O�L�W��07^쉳ػF���d"OH-��(V�m|$#!��m���"O*t!��PV�l@#��60�����'��%�b�FM��[��C�:���2�'ǚic&��"�>h��V�2LTu��'���D�ͤ>F�Ӣ	 %��9h�'Dfy;r$V�ms�cBΓs��j�'�E�s��h�X��Ǜp�� ��'&���gL<|و1��cR�I�'����p&�I�,pkao�"p�dR�'v�pp��ۤ��u�E=bف
�'��x�j�H�T=���W%r �	�'�<y���1�i+RL�
��Z�'b���AS	c�9�n8Xp��
�'���G� maRL�q/·Q$:��
�'(<�U��z!b���$9�4���'��� ږ_g�����6���'_N�C1G�$N���jw'A�B�����'�\�Q,�P��LVB�:t��'�^MIħαJ,�kέN"܀�'�X���n/
�1`C�A
nd�	�'$�BSD�cE>���M�΄�	�'�N9�Ãbb�`��� F*M�	�'ټ���
�:Wx)�(�+Έ��	�'�|�HtҠM�"�%(�d�X�'jpi+��!ʦ� �]�*lzDz�'�N�R�(?�`�0 ��&"����'��1X$M�z9S�L3F-�'!�)2��9�Ԝ8��Z xZ&�
�'��L��Ѱ
B�(�q���
�'.m����&d� �	/�k��Г	�'��l���%<�K4��\�8#�'/��n�z��Ah�	���	�"O�,bᆈ$&�4i�S�~�T�G"O�-`Ј� v!� 2�Aʜn`H�r"O��)� ˰=L�+vk�?B8A�R"OL��t�šEH�I���Z
^0�d�"OҌ�҅X�3�i�E$ �$�(X�"O>����Wְ�	�"[6 ��Q�"O>Y(�&�*##���%"��gFL�E"O�TsB铯8H�(e�""a�@�C"O�Y�(K�as�i��*�i��H��"O���b�Nf��P)j�pհ�"Ol�F��ö�(
�
	�S"O<L�wG�����&��90�� ��"OP��p�J.Sb�P���H�"᱅"O��4&/�2aX#�"F�(}� "Oj�抏(��ܒ9x��8S"O�U��/Y���P��/�w�ԃ�"O���w��L< 	u�,|�\yʴ"OR�� ��)7��8��E�{i&��@"O�H�Q������3"W��h�"O� X�Ya厃\
h�H�,"�����"O�l(�c	��At��'J��iA�"OH�����3��В�C���h�"Op\�&AC�����K���|&"O4%�e��SjzT*/����ʠ"Ox����U9��w.��{�n��"O��4��<^gJ�9u�_7��]�"Od BW�F@J��A	-��4��"O`ВDY2[6��JW)٧$�0�a"O\�s�oB�j�p�GIr��!�q"O.�U���@��J�zf�upc"O<Թ`b�0]TΉ:�o',z ��"Ox倂��eiQ�ĭOU�2"O�4��_�z;�ř��E�y:qk�"O�)���W''���e��T,6�Ȥ"Oށ*��Q�aJÊ��nL"OZ��@�;��9�^;��ɉ�"O�9P���z�*�b/��E8:�Ҕ"OĘcgٶawB3�-�yF�=Zb"O&��@��ST�{��#H�R�rE"O �F��eUص�R��
V|��Ad"O:x����A�(��"�.3nt�Ӓ"O���@�@1���s"��$dD�"Oh	���f$��K%a�\�-
B"O(A��S(y�D9±��.e�\�+�"O8�WmK�cc���L�����"O�KPDձ*D�
�^�
�d��"O�I"���	@�L��c���h}�"O|�p�"�|���SkNd�3"O�`K,<������q���g"O^��3oW�
xX���r/jĈ"OVT���Ʀh�R�� ��*���:�"O	�� �"�����kj%;"O���Ӣ�#_�����B�|����2"O4A�����H��r�1d�:�qD"O@\ael�$,�d�C��>�S"O�	L�tm4���*S� A6"OR�@u�5�!�Ԇ�/8ۦH��"OX�*6�� !`��tG ��xk "O�P���ed�6Z�ʹ(P�"OH���'Zz�Qڱ�_I��AQ�"O
y��-ۖ8
ظ�MXsK��"O�s�a�@��Xс�ջ
8��	"O��e ʂH��x4LK4sp|��"O�Lz�B�$�N���G48�8���"Ohyį��Vr5x���y�40�"Otu��P�x��0����3�J�z�"OL�ڂ,�%d:�3fd��>D�����ͺdɎ �3i�C��	p/<D� K�8,��uځ
��9��!%D���r�իGR��P�@]C���"�!D�8hѮ��iB@��pگB]҅�5',D�X0 �*'�<�תX2	iV5c�$,D�(ڂgBQ"��k$�]j��>D���=^0$v!��-� J�6D�4 5#�"N��Uk.��ĪS�4D��9�oQ=uu���W��#b�T��O1D�4�B�	L�`Ѩ����t@�;D���6N["`y�4
(�nP�m:D� Jw��M�=C�>�P�B��7D�`+��y�J����!>B�0��(D��@����<}�؏B���'j2D�td;�9���3eQG�1D�<Ș�ͺ���-��Y���H�<� �%���7T�����[�=>$p��"Ox��k�
=u`�'��'���"O���P+�,h}��P���S"O��I�l�)��{F�ؼ#v��@�"O�([��U&
��H�'��> F2�f"O����NV�n�����'Vb�8�$"OR�(�N۠<���Ӈ��	=�IH�"O��/�=6�a�Ą��1@���"O,KvD��2�Tec�����"O�T��A O��#�AŐ?m"�0�"OĕK����m{b� ��؂��	g"OD��.�=vV�B�[
8�D���"O�Q���I$"�3�+נ�p�D"O܁��G��U]�@�`lH�W?�ҁ"O6�9�
����M LF+X�q�"O��ID��$Ip*#k�'��9
�"Oމ������IZ�`�~M`&"O�58�E�Tp�`M�I5Jt��"Or4�ר�A���!u-	�#{\�j"Ol�!�-W�a|��K�:_��Q"O̍�ʆ�_�Z}:0j]�c T�x@"O }��b ez=�	���X�"O������N�Ј�C���3����"OZ4����63�|��FF� �Pa"Of�*�W K���W'�{�|(�"O�U�71���y�TG����u"OT�Q*�0)k�R��3P+�|Kc"O�}W�B�ai��"C��:%�1P5"Oy����6�Q�)Y�fQ�"O��R0����HXyD���@��y�䉚D#�$���U�}!4�Џ�yr���X|�a�U%P����\��y�K�2o�s��L��E��:�yB�E818���#�B(�X�š
#�y���Jt��'�$�����O��yB�L^n�	���)s��*�X��y�E�������h@;�m�?�y�,�2A���J�#�8~X�4�y��ݦ ���L h@ެ��M	,�y��@�s�-�d��&g��p�U(͏�y�c\!������ J���"����yFM̭�2���K��Y'Kü�y��:�ּ�c(�?�������y	T�2�5k�/B�nD\r�.T��yb�^�vF��3�h�	d2��JԢ�9�y��8D�=Pe䜌%��A�ɻ�'�ڍ�'I��yzd�h!5D4�'Ƽd�4�
<P	���݉-�>E��'N����Q�T�t�Y����%,H��'��1D�=]���%���ȉ�'zFj�.�9�Fi���7&9�p�'�8H�t��# 1N���ÜE�e�
�'3�[C�Ps���!ך��y
�'��\���F~ᎁ6K�9Y��a��'�R�{��݂L`�0��
KRf���'��]���@�])fJzK�T�'s�e�E(�n���F�,u:���'���ʆ�͉Yj���Js�\��
�'�:IB������e��W�<��'���5m�<*f8]����+U�2\��':e�wJF�b����\�S"�j�'^��۔��v��T�O�L�Vd��'�J}r�%��s<�J��5G����'
t��Fʅ�k��Dl�Cd�(��� X�c�J�T�z�Hp�rp��{ "O���$GH*x66(�@����<���"Oʼ���+~�����i�޴��"O��ӳ�V5DY�hH� F0�"O��례 �7L�h��R�Y��Y�"O����]�_�$�pSf�-���6"O��:��A��dE�Վ�emZٺ�*O�(;穊�.��˥,�4b2	�'�h]���4sb�)ӕ�а?����';����\�C��#���2��]��'|�	�B�����hS��v�J	�ȓj� �x�L0�@�8Q�J�,��ͅȓ'�8���9���\-Gf`���x��ԅ��1Ϝ)S��V�X�(I�ȓ~�b�j`��g�:�1k�/T\��v�B���-�|����-�y�ȓ�B�
a���M�Zb�Sb�(`��5�rhk�/^��$����)�ȓs�,�9��J��B���ĉZ���ȓAU
��s�M�q�N��A?,�q�ȓ�<��D3L�UЖ��c�`|��%��	�eKN�WP�Q� C1c��M��4Ȏ�k�d�^
��1��-����Z_ڥ�Ν��(�BCJ&(� ɇ�1NR�Uo�}.޹w�ZX����ȓV��i3���I�ba���j�L�ȓ;Ɩ�#��y`kfǗ\���A��b��P�0ٞq#���b�\�ȓ4��aq�CF�J��0Q���#����\��m�j�<l������j�-�ȓ~������ϒ)�b��1/دU��x��p�~��CC�1��as�/6����ȓ7N�*�CC{;�P(>����ȓhЪ���Q�'��"#.��$�<8�ce�=Y޼�5��(����ys���-�BUP$*%��0����ȓ[��P�J�����ǅC�K4���jAN����X�<=��k
ژn�*݆�_l���6��9[�Ѵ��E�؆ȓe��Y0#']�\�$��U�\��݇ȓ��]�t-�!*�\كN�"6��ԇȓ��h�j�qP YE&dB���G�ȭ�q˘0{op�`�I6\ň ��5�ࡒ7�Q�^�Vi�M�
{����4�T <���ꞖO��U�ȓ*��y�N�5"�i�KAj�"���~a� WEy�t;�9FM��c)���� W
Thc�'\e%ࠅȓ'�0�)akβ(��P�	f:���Y.1�D�G)^re�d�L�oE����Q��E
DAC#z�Hl�����y|�ц�6p���$�|ʮ��'�]�,���U�
��$���gΘ��B�=~�P�ȓ��X0s(�(3�t��U����U��90���`HfI<�"����Ʉ�|jݹ6 U�?ѢyQƋ[�;a����S�`e��R�OX��T/;m�^4�ȓ[�I�ǀO
��Z��I����ȓ\5�P���\ ���X�Gf�ȓi4i9 $Y,��Hp��T���ʓ{=B%��%϶]|�
2% 4=�B�	$�ީ�b+�qTVA�!�8G��C�ɼ�j`��ѠJXR��u����C�	r|Ґy4�O�c��jQ%�<��C�)� j۳�И?kt9���
[RDZ�"O��R@�R�~zJ,���H)��P�"O� �A�{��z0���!�J����X�<Ac��'�j$�r&�PE�=RQBR�<	un��M���,�t�1.YI�<�C�OE*�wkH�o��I:�A�{�<���ɦ`.�i��T�|��Sg\�<A6�B��l�x2�י]����[�<I��ō]J.%�'kD�R��-��$�M�<y�OD��Ⳮ�Iݶ�	�g�G�<dL�j|�k\ ��ѡn@G�<9�LR�i^=�r���\!��'��B�<I1 L�*r�I{T+Ne.u�׬�z�<� aA!)��L�dk�<E@�*q��q�<q �B�U'X�3��"b ؑZ� I�<���J����VoC�a�
9���_�<�&>Q|�z�⇚R�<Z�.�_�<��aU�,W>]ap
.)F����^�<��!		�%H�I[8��i5�b�<�bL\�]$�5�6z���Tj�<y$*�P_�9���� f+�i�<���/v�~|���:�܍���b�<�$/����Ƨ����`�w��h�<��W��H��o
1I
�9u��I�<�C��n��I"��M9�J%Ac��I�<�DJJ&N
�E�󊗀Y����`�D�<�U���E�	�]7a��S��B�<9j��H�Ș�����v̳1	u�<��F��D���E�6��#�lKr�<j��J��-�F�oL��d	z�<�҉ܴ����IC�k?8�AhK�<�e`V�Y�쵰u�ʚM����G�<��hC�F���ï\2Jl][P�GX�<�6�`�H�B`�2�HF�U�<���	hL��"�9 $zP"��h�<������UBq�ҵ�d��D�b�<�#��I���Õ#M/C�p�@7e�f�<�,5�yC �-9Ƙx���H�<9��94-$��U#�:J���'�@�<!͉�?4��3�N<_��Qf�<�@]	�j�kH�Bu�@C͈a�<IS.�7��[1��zDZ-��O�S�<!C�� ��,�rc��Z��
�f W�<�Q������F�^!� A�T�w�<���	6�H���!>[vt҇�]�<��k�d8�dI�K�4�Z�@�Q�<Iө��o��-����=w��pi�iO�<! Eդi�4 Ǵs���6�Ic�<qC�u�B�����3u.�t1�`�T�<)bg� �(0Sg)��}q��ځG�<Y�k�4D�Ƚj�-2�J��@D�<9e��s�(��E�A)V�� 1h�@�<��	ݎ-*��do��N��}�ƣ�b�<�a��!^>ؙ�E��'{/�=	��u�<�eF�x�\d�SNкXFR�2��}�<��埫@,L�sHL�~��`����}�<Y�킉o�9a�
R��5���|�<��^m��h�ȋ3c:��u�m�<�r���F�����~
�0���h�<Q
��;�L����*2&6�� 
g�<A0�5AW���Q��0��\٣��X�<��G֎P���УR��`"'G�K�<�w��ȴ c`V*M�IZV��O�<ag�Vh�V=�����ؑ`K�<� �[�K<g2��sph�*�}�t"O PQ'aR���X��ĝ͖�R�"O$�blǆ%�(�2`�D����	�"OJY£���e�PbCT�rn�]�"O6-pq���v���xf��c~���"OHL�S��"+�0����Qo�,{�"O$<B�EA��m�v��򺈛!"OB����]z0�[�A\:6��%"O��X)JPހ2�G̛)2|�#d"Oʁ@�bPfk�I�씙&����a"O�l*���>z|,���˖L�#"O�ui���4�mE. QŮ!��"O �a��!,�ƠZ�m#]��d �"O~5ڠN��]��L�k\���"O(�UEU�s �Y����`����"OY#⌀�A���K�8W�<z�"O������ A�1��N�=�"OW�=Bh�H�)��L���@"Oֽ��Μk��q�eh����Q"O@ѫGi�%c�|���d�$q��"O��` `��H$d�	�f�TS#"O^�b��m����刂!
����"O�ꄯK4U�R�X�i%D�x�P�"O~�@��+�>1h�菟?����"O�1�a��. ��)�t�2˺��A"O�a3�+�.�Q����sR�@��"O�������_{�����N|��"OZ��+D-el ���uFrM�t"Ov\�e;k�aT!�1dH��"OJQ�B�2dL�"�T'sKf�!�"O�!O[�<�����M�H$�1�"Ol� ��! �:�
�kC 9��Y��"Op�Y�㕥PN0�Rd�<�vXyq"O"y�wH��n�+U��BJ�"ObY1逧R���@���;{�}�"O����o�0ؘ��M�Irjp�"O�U;�A��64-`VI�<Wbd���"O<I�T$�%��K�O�x��T"OTU 2o8���ʒ�B$��Tc"O�<�Bb�V>�G��ur��!"O0� $�\6�T��'��8rq.� �"O^�ڲ�ϓ��WD.iy�˧"OB���N/��T�d�J�Gi���a"O <PVO!���Aa�-*d&Ӄ"OV]X/Rt�8���e�'1`0z�"O�0��� 9dT�W�P1�i�5"O�eH_�g�~l�p`O�آ�"O���uY�$�0M(FT
�"O����-��1����h�����"O4�8c�QJ��|�p"��d��2"O����\{�mq��3n[`5`�"O�(�:�L�k�	Bb���"OҰQ�H�(p�m!���uA��r�"O��9�@�(�P�)��H9@�4�D"O�� 4�հui�E�&o�;Y*,�"O�y���S5?�\�f��s���B"OP�*�g�1#ۤ��3Lچ<���E"OA0.��P�+0��g���v"OX�!�d�6Y#2�cKB�6X:��&"O<�9Wg��e�x-ـ)T;,A�ȣU"O��IO��a�rP���R4G0$�Qb"O޵UEƞl#,Բ�f�(a7"Ov�0���c��|@t�E�<�j��"ON���ę(#��E��([d��Q�$"O� �� �
�M>i��$�p<6"O=�7M�6Q^���P���Ku�x�q"O��A2-��E��*G�as:���"O��Pc�X�0��!qoh��.J��y�G=���#-zgL�"��q�<)�H�?$��
E䎲Z-�5��u�<Y�Է.�|�B��P���p� q�<�$�3+4�� �}�F���Hl�<�ݑI�ܰ�l�8�U FHe�<Y��X�&��P��Ӷz��}�ȅz�<q��]����"�]�K;V�Jg
�l�<i�@��E�Sa��G�-�S�Dr�<����G�� �W�ү�F���cAk�<��✨o������K ��he�d�<I�KLD�q�A���b�X�<����@��=R�T�F�Z�h�<i5b� �0��4�+`��p�d�<!�OV�:  ]"Ў�#1,��0*�a�<���K>F/l���CJo����7�[`�<	 �3q>$�B�� w:��)�Y�<�)F�#,� ��
<$vp��fX{�<���	t�H�w-[���a"R��<����h�Pv��4m�u�Abb�<IQ$�-�f��3M�)0@8��r�<a�ƨW�xR��
oYv1(�TH�<	 �Y�F�.4�0e�-�<����l�<�e�
VbJE�e�-5a�;���c�<�gMP�kZ�$X��p!�G�H�<	%�E�X������ &ܵAA}�<�S�0	l��B,��3>�QY���`�<����:.�X%�
�F���E_�<Sk�[^�YK�&��5���8�	_�<�g�0Y����FD�Jd�p��Y�<�pLS�=������F8���'Bj�<���]�~tDCe�ׁT�p�Sc�q�<���5
R4C�Ǎ<�Xu���c�<�$`�X\	rR��W�H�ڑ"�_�<Fl�+p�����ց�m��)D�<3��B*a�����V�G���Z��"D�ܱ��.fa^�I��T�U���$D��[�@�?>N1XK��~���C�>D�Hf
��n�d!��qEޭ� =D���$�ɐ`Ș[�E�X| ���m<D�l2��K�R�Hk���&��-@�E6D�է��N�y)1�Շ<>�uC$�2D�|���Y�����S&^���bd+D���5�����y
�)Q,;�qh0�(D��&�s�!Z�L�^Ak�e)D�`kֈ��:��=�4P�Xu��/2D������O��AS!A�g�&��5D�ܰ�D�"�z�����Q�,42�)/D�����YL�-�#O,&��.D��rfEяX� )7�33l`H���1D���恭b���.ˣT"@1"�!D�Lkr@�� ���%ɜ�L��01�+ D��ɤh��qPL0TB��^v�Xr`N<D�TS���53x�Q�L��>�X��B�;D��iG'� �1��AQ3)�Ȑ�"9D�h�gh�?}�^�h��,O?�j�';D�B� �s�,����MJj��"�7D����Nĝj����Oh+>�e4D�LhB�]2E�BJ�-f
Ta�l6D����'�9g�ٳ$K�tD���g8D�t ��)�Шv��7\XdXSB6D�� ��	�k� EX0�EK��]���f"OL���d�Ϙ8�d��`� �1�"O�qč0.��H 錐?�0�H�"O��Р�Ɯ�8(�"�+1]�0
�"O�)p!�)a*i ��D!e!��P�"O�*�z`J4���S�T�r3"O<�t�ߐS���JV�o1���1"O�ISh�j��r 
Q"K�FlB"O��aD��/!���O��b=�Q"O̝��v�(k���tx�}1"O�E*,�z1�&#C�J���"O�@&�W�Eq����1G��x�"Oli+rHC�F��|Q�=�:���"O�ЈRS�>i��ߗ=b�2�"O2��`�V�M`>��+$Nm��"O�e��V}
`#CT�E����"O ��A/�dTXQ"�̇��X��"O8hAG�ug��u �.}0��6"O4, ��H�s5.001a�?d�"O�5h�*y���4 �'�=XF"O���7��W9���OB90z�0�"O�5����m���p��BЀcT"O��z�E��H5*�O�^�p�
"O� �����~��V�޵>վ��"O��Sr���G�$JSe�1_ ɑ#"O*���l�i�:�k�F+FTdi�a"O��2$	V�a�F|c��4\�ݲ"O��0A��V��!�W�J9L(aӠ"O���ϊ�E�V�C E�H<�ܐ�"O����� �\s҄3��ܵ{NF��Q"O�e0r�!�|����ֽD�M��"O�����G�X�����f�8O&]��"O�kcc �]:$3r���_���"O��#�IJz�ۧ��c
H���"OXْ���l��%1'��7<��"O�p`��̨�����!��z徑��"O�)``��p�"|��+�9�&<�G"O��CG`�0Q����U C��%��"O��#:_%PA��Z�.���z�"O@usNK6VU#�F<s�H8�"OL�{҆�%6h���W䗊+��"O�]��"^>g[�l���5�$)�1"O�١����h�C��0��a'"O�@�#�H� ���H�?�6�ʳ"OXj������5���\�g���� "OBx��>H�&̓5�6�F�j&"O���$O��Ik�B�Q��]����Ymx�<Q7m�V�*y!��,Z3��$d:D�\���U	�e�!g�>�@�P.Nfh<9��UT�@���&О�xW!px�lDxRi�GH�!��K�
��� �ۣ�yBF�]~��C��Tp�  ��/�y�)��uh���
���a�c���yR(�|�������>y'@��3���=�{R�U�c��	Z����wt��r���y���;wR!j��s������Px�i��m��[�� 	t�ܤlL���'�������l�:]r��Y��Zu��'.Ѝ@d��+�|X�"	!Ƙ��
��O�(	 	Jq��W��,8<XP$�S��yb���~��u�d�կG��Ę�G���D���(O�O���D)D'!q��Qp@�z��ή5!�$�2i�8 ���_%-m��	Ƌ�v�!�$�d�ԩ:�@
!1ڴY�j�#l{!�� �H��D5���qBL7P�f!I'"O*P�#.@�W��aWa��4���ʦ"O�a�vυ>+�đ�@HzQ����O�=E�LI0���'�^ ��͸D���y���:N'�y
�ߓv�DI���^��y�D~�ᅯi�VD2����x�ѩ,	��Bb�u�N�s�@'3PB�	�A�\h�L��i�|paDo��wg6L��S]����E�(��i`u ��L_���=����T�f�6�x�卌�b$�`�$�?����S35�|��%="A��c�.	�V�rhFy��ɃW^�K]�?(�{�bԊF�@-JAǒ���?��'�0�����x�4B�#E�p�[V�5��~��w�'�R��cP6Y��A&�s�V�H�'�702��@ʰJm��;��E!����F�"~�W�ߡU/N���Ϳy��d$I`�'�?��WK��n%JK�-�R���G.�	d���ӵn�@3j"�Z[�09a�*�<AȌ��'\Q>i����c�p�	S`�R�:��p�(�	d���F�� y��Թahۈ	1�eJi������$�(~� ��e,�8q� baE�K*!�d��d�+�OI�cd��qp�N?*!�D<ng �8�ʏ)�j��I�00�!�Af�t� *}���y�ǀ+F�ў��	-.��⁉h�X���)����D/<Opّ�A׊S�"�!G�¶x{�}��'i!�$�-�>�b�LP�D&��	q�1?]!���	kg��2�T�/�`��n@!�$��cT��Nt��Ak�E"!�E�<3V
�+k��X�`�1V2!�d_�@���a�]9aeRp�/ݲF!���z��"�a�+2�$u3�LJG91O���DK>Gp�`����>��P�k) !�DG�#A����oR�X�8�p��;p
!��Ϋ/���T�(k�@�1I	��!�$D"��g�'l����$��!�DEf����� X�A���q	ǚN�Q��E�d�Q�P��3@�)5Ԗ�z$��$�<�I>E�D��0�1+R�!*R�X�%/���hO����E63N͑�բ*:�[�Jɋ�!�$D�$�`��_ɞe�/K<n��D�tF��Lo>�j�I��rMr�[/���yJ�J#�a�b�����a��hO����<^e�4�ȁ*��l�R ƽW!�D_�8��u)�����R(͂R"�P}�x��	Gc5��I$)̹S HYҡg�e�t(����O�L �[���h7
R�ZU PԹif����'G|R��$_�.�N��7$G^�\�=%>��=a¤�=\���z!��(�1��c�<��hB,C����V|��dh���<�� 5�S�O��x��j֓��8�� �y���
�'T��g��=m��*�r����' �L�&��l"���T���'@x�:^�.$c���MX��3�'`jJ��M�TH�@���U�u�K�0���������G�:v��z�l��F ,B�	��U�6h�4h�p@����O��C�	�G3L��E*���PH�åf\�C䉈l���慃1(����l�'��C�)
��CWn�eH�ƥ**YnC�I)T����!`U�]��|ɕ�
�Wi6듲p?��#Đ���SE��2���k�	�H�<	�m�_*��B+9��y���Ol�<9@c�*�	��S�w���2��k�<� ��b!�DZ���iGD�lH>M`ON�DW)S�!s��h�
���b�!'%!�ܗF��Xȇ��p��iH�aE�j����W%	i�OFFyw��$�ةy�d� �|��'0ڝyPc��f�ҳuI�0O>���������!���MYzT��M�6��~^�l�ҫ�Thv�I�8-���
+D�\�T�-Mu8Y�%
6�y 2�=��V}B�Pެ}��cF P�v(�W,\��C�	 	��8�&�@� 5S��z�RB��+/;�!!�O�Nڬ��ϙ8:�B�	�S^�\zY��.G�n�hC�#}2�'Y�\�l L��ڀ�Y a�)�,7z�,�t��Q��<%��ɨ"�A�N��'��F{���ME_b1��	�:��p֌&�hO@%ڋ��tr�ۅ�]$�������<g��K��(�ι1P�Y�4����Z�uf	 e4O:�=E� ��P�6�YU��Tiy��V���@iB��DE��	�FOɻ}T\���e="��rH�Ŧe��� fƝPa ��Ų�1D��3T�V n��� HƪN�hX��ɨ2�L�}��4��D��O��=�|R._~H<�4-�	R��ƯC�se�A�g]j�!��%�x�U��=lب1%܋U�a~bV�T��X't�&qP�%=3P��!)D�@y`f�8X��A�G�21�h� ��;�?I��ɞ\6@��i���EJ�a���~�W����	T�v�f��J��8nLu�����D�}��dP�䉸�>�pŗ/HQ�E��M�>C�0�0�>N^2�05oЉ���1�O
)J��^-CN�\
�ԮC��ʠ�O�EGzJ?�O�T���МʕI4�\7/���is"O�`"F��=tUZv�UE��h�F"ONM3脄~�<S��CC0��v"O����"jʔ�k�2A(UZ�"Od̙73���Cq���
���"O,x��$��$e��s�i
�Br�-(f"Ox]�2�î|��z�E�U�� #"Of�S�[��s�䜟0|,�)�"O6�L�&^���������"OIRK̄a>��X�@ĀK��2�"O��1"&��g��8�ƛ,�z��_����h���(O�mA'�&�F�(��Z�M�t�JQ�'�"�O"(x��^"a�??�Y	��$:LOJ$�kB�Y)TP35���O���
O���4h�)�B�
����$uI՜�y��Z����R"�:^���ԡ�����(��u���W�8��]!��&3��Y�@�1WG!��BV��$�D�\�1�Vd��i�'Z�'~2������0k$��`)?q�l�ʱ
��8H!����R��� �,��1*��75!�� ,w|��/u��#N��,1	�'��t�]H�@�f"��>RtmC�'�y���r�@=C1Dھ��
�' �zl�.��	�P�ܗ� R�'�E� �"��pc�O���I�	�'�`����,C��	h��Z+2$�'sB҅��g���b"�Qw�P�'K��b�*ϢK��0�-�(I@`@��'� $��h�h�x%�!-�xP�	�'Q|��ġ,K_���G �!hx��*�'��1x0G�6�\@�k�_����'n+4Wo@�+WW1\8��'����L�~�j8 䁅��a[
��� ���^>2Uxk��5%&X۲"O$є�X�(D�	�z<J3"Oh���a�?��˱I�Z򂝈�"Oz�:���
�z�s#ؕ%��P��"O���W#E(��sg �%!�p9��"O�j�lڷU�r	K��H�t��Q"OjѠ�+d��m��h�5�╘�"Olau썼Ak���朲?�X�"O����O�|:�E�1�Ե>�Ҍв"O�p��+���%�RL��jG"Or`CC�"f.�]��^��N�"O�T�C��^(`I�qEݮix6$��"O4] �ʮ'@���0�	H�t��"O��b�(w(�`#�<�f��"O$�cIU�p�΄1%E�-����U"O~����v�,H�wκN&�]Ғ"O �U�S�

ڀ�4ǈ�h���"O�=�57T^&�� �76^D���"O�)06�3x��;vgB�qG�,��"O���#�C*|�*}2f�]�����"O>�����/3|$�r�B�<������J3�'�����L�W'H%����*��4�	�'I��� �ُ�"�	6'��/���:�'�.T��L	R[Di�EB���~,��'����M&`� ����	R����'��e��EP$q�Z1y���t�DY�'��(�(�Q��}�VI���R	�'���m�2q�]:3)C2t�����']z(V�G3�ڸbK�,]��Xh�'b>*M�9��00�O9Y��Q
�'���h�
4Q)��p��
*)A�er
�'��%�`A�/|;����`�)T��8	�'�a2��G�6�h�ց�$2�)�'��$Ν?.}�-�UK�#@�x�'~�PA��[.ܦq�PB�$\�:�'��I[`��6�"����U6D��	�'xr BfP�n���2�[�8��0	�'��mX��Ԍ$ �H%e�>
��x3�'=���`(�o��|�sA���@$�
�'�<P���(s>P�cD��ܜ[
�'�ܕ�`o�	�q�� D|�b�'�@��a�|�����}���h
�'�q���
+zp��#U�7h	�	�'���8B���k7�U��끶t���y	�'�AA���E8�tDPܑs�'&�����!UP�$aB=Qʱ�	�'����i�!3RR!�nY`��,*�'��Y�$aQ�@� 	2C��X���'���P�O�:vp��Ǒ)<�D��']^�3�%)��	�N}�r� �'jp��/G�R�+rM	�\��|��'��*3+X	e�`Yc�S�����'2	g�͝u�~q���O�*��'�H9D"�/+�(�s�D^"�Z�'�Vi�4ɗ	A�8�8S�Ƞ,E2
�'����ԁ��U����̊&�,`{���MM,0H��*��}ޔ8bp��s��yS�>S�B�
��E��@[Ů-�UA�����	�m�u�L�[�S�O�R�'.��3���B�C�pՂ�
�'�j�� ÙsV�`�������)O�Q��I18�2w'O`��k�>kI:b���'\F�2��'^N�rE4�v���X=����Ĩ���d��]h!�$_�[���@f�R�2��}���®Enў��'�� &����Lf�'fꌻ��)H��RgR&B:h��S�? Z��JDP����@5��,��'�N(Q���h4,xCY�"~BUnN�I��"V�#8�%�IH��yb����`[F��Fop���f����$Y|*��G�
���M<���2D�	$z!�g͈�|ay�%�J0�n5!�>�3AN�X
-�g'��(��!q�X84;����`PB<�fP�X�)�bbؤ�u��R��E:"��]b��%���K�f�P����g�fF����،-\i��D��Z.c1b�`�%*LO�񱀛P��\��a��OR�5�w����� ���4j�X�D��}1��P�d���ё�J����hQ�'��a�K5�*���
I�.4�-�R	��,,��q��D�p�ڴA��	����a �m ��]�^��,O��: 4�T�\���s'�(\�Fq���$p����4 \�C��DM[Eƚ���<�"�(��0��T�Qn����	J�/p�)���zVCE�*ˠ|qA*�5mƚ�+�,-?�bԒmՔ��9}����)r��:��NCf�@���(,��ė�5}��{��jB��$h�0��s�� #J��gGі)�\�N��2ŏ��+_�c>�"�o�-Pڙb�mт]n�!��ɿa�Z�� (�zh�9����4㣍*\��F�mBfq�F�8Ր���%��F�z�q5���B��b?)"�&|�D��n��V&���n?O2���p	⠺H���t�f�l��5͜V�y��J�Ns\-1���Y��iq-O?�d��OݎoXH��$;�h�{3����rG�*M|��*ז>E�D��-B6��&��q!(O���Ri8�04��C{(��$!d� Gef}�H'ko�(J���t�Q�M��b>7�P�D���!����A���f�M�$w-1�N��6��'���cٲa���S��:T�Qx1柒.5�=�dɗ̚$g?§h��qi�폏z�P����(�2������|rf�6_rAQ���=_&XiӇC�2�y���Y8��A畉f�fD,g��ȓp�-)�U	0���d3�2t��rbd�1�A^�$(����-�3}tF��ȓl}���r��T)��s!/t�Ն�+?�a�g���Q6d���@�dC�܆�Nx�ɳ��
�����ޱ� y���tkʌ~ũ�!F�<1��E}�@�'p�����ל;f �O��H�@���i������T�'6�r�'�,z��,^\�-���C?�jh#�'���ʕe߃z:�{��7#�?Q�4����X�D��;��qV�<\O.�0�C�~�] �'X��毀6��L�7�nql4R�E*c��i�I}�T��6gƢ���I�bP�����2)m��D
*uSx�Oe��$ʪtWr  qaFe�V��x�b�l&HWʐM���b�qژ(���q�����'���Ċ�?K��Sh�<dh%�֨Q�L��ѓ�O���s�Vl���
�<N����>bj5ўw���je=�2c#gK\H��'���r�ج%B� �,*�P$ɉ�W��b"�1"
�Ū�!�C���Ba�-'G9CR`�.)��ON* ���2��YB��}HT	T�'��ѐ�Z�q2�X��"�"97�T冂��V1)��n� Ё�Ql"�{P��wn4�� V>�<��
J����`:�� ��KVyR̖�#�8xZ�d	*U~�7 �a�I�1V��΁�Ӎ�D����b=��j��MW셃��QM���� �'�"�Yi�=��s���6戭��jS�c����A�N;۶�Y��>�(�av�M?���[���7㚉�w6v�d˰D�� �G
y��
��`Zj�zC䁣1`@��f��TKMM6II���A$�Yp�o�6q��p����OLB��Yb�\CO?���� �T8��Eb�:U[��	:�w��B���Ι���N:s���{g@�:�h��eI'@|��	��>$�3�O8��cL
K^��N?��ېGH�f�.�B�F�H�r����>QG�W[=h�F��@S�M�s��3��OZ�u��䛚5W�0K���ͩ��>E���s؟8Y�� ���Q`�N_'Y�D�Ơ[��( �����X���j ������MX�����	�dS�$Z"�"����L��0���I>ͬ�	4-�}$��D�<l\f���-�.��h1�O����֥F;��'����FL���KR��	�b��S�&գ�A�,t���\����!�@��)i���� .I�#Ȩm�( ���)8������sܓF��jXtax�\�t
̈���Ll��������DƤ<a�|"C��>h�`�:#n��;d�|Zu&[ +�ع��^
�y�⢆F�<9�眹h�|]�L����` UK�fwܹ�Vl״@�t`@ꊇS��\%?������N��a��C!��qf�:�O����B�T5jr�ŕ��}�B䝒"N�x�cѣ"OVDA*^'��=E�[���z  ��(�Kv��h�܊G��֙�'��1B��)� ��!��^4�� �0݌d"O\�jDN�:@��E̜%`*�☟h�Q�;N�@�e�*W��D�T�ܕ�D�g�Be�Z{�
B�I�ݶ]��eK&_���lB�}���O\���d,�S`��|"�E�BTjȩw+Zj���҇��xB��)CΒ�&m�y� �(�հK∔*�L	`�����I�y&�����/�	�Q��SԲ���īCCtP��O��Aa-I�"��(JV�_l���:�"OPEa�i���I�u�U�9�$قf"OZ�ġǺ`������!�B"Of���ǆ� >�)�7m�*q� �� "Oh(5-X
���lS��u٦"Ov���N�]���AS�|�.!��"O�����Eid�G�����m� "On,�/֨b���W��9K�|��"OTq5-ްv肩[&[�#�l�F"O0�!!F�b�UO�H�f	yg"O"�"Fj	�k�� N/_�(�ib�|�/^�,܅�	5ހ�h��A�C��xy+	 \�a��ߓh�E�@�ܨ~G,�:�g�)�p���Iա�D�9� ����G�r(ذ��0(Q�����J���`��)є:-|�����D�(IlٗI�!���ZD6J@aуo���P�&R�q�dP	�
T�do���)ڧ?����@C��_��C���:l:��ȓ�"P��
�ᚔ�3HČMq,�O�!�瑋��L0Ó[?�u8um�Ex�%+Q��}4B���RAz�X�·-p����bՔ=ʲ�(C�k;<`�"OX�P���-�!H��ÄT�җ��Ҍx�h�J1�DU{��J� �Pa1$�"���ku"O�� !��f���Ք}@��x��O�4�k�r���J��}�7}�q�N�=f����g�u�<Q�-��_�Ʊ�%�B�n����4evTI䋕65�ax��Q�ؤ`�"D� `��������?	t�Y�
�$�P�`؜����.ؗ]�4�T��Px�
؝6_�\���S�o/�5Hp�W���O�t�S�ڦ��O�X�q��� ���%'��r�]�
�'kޕp�	��C��f�Ǝe82${�'($a���Ҽ ��=�F#%R�f|s�'�t1)�NX��	C`��M�M��'�J����ǒA���'ε:�\����ט{&��~R��?{�1��$
�F�x��T�<!w@L-Y~L`�%KE�����.r�Ȫ�g�V�`n��C"+������g\�P�� ��Y�� ˷"Or%�e��o�qp�o_��2MH%8O���v�ل���O���&a���1��tj�,�����l���"R+.�OX)�"鉬�yR����P�fOܳP��I�%�
���s�LHr�U��<qD P-Y�$�����]�@�G�^�'}
�)���m�IFx�!� �,'J�H ���:����Ո`��P�OpK!E�G��(`��3tH ��1U�MP��|����^�a(��B�����@\��YdR}��9"O$���׬a��qk��ܥ
�hh{#�'�p�ZVkߴ�U�O�,�o/1�"��o�B���a'3lH�b�,D��;G`P�&�deJG.��y�D��G
�<��ɝ�NR��*�?,O������ m�pP(���"z�j	���'�b�&ʨoK�ɓS�ݞTs�IpDH+y�Fi
0�|H<����6g
�A�CFQ� ��% ���S�'Nb��-Y�p����~R�Z��c�z�.L��ES�<AB ��S�C���4��p�,N�<1�a��&��	AK>E����&#_�Ey�����2R���yr��� �2MM-Y7��j�����ɚ[�j�)��'�j��DE�xV��%d�3,��'2<Y`��9y���K�|^8�'-��#��+�"�b�'gR�2�'��P��9dF-2���$������� z�9��Ñn׶9�qə ;|J�"O4,J3�޺S����h�� D�qS�"O��3��7n������	W��4
�"O\�S�&+-��RDJ�b�T���"O,]��j�&��Ɇ�+X �"OZ̪�H��*�zv!�T�l�q"O<@KS)Z'N��-7`A'z�-��"OF�pT)����a�c~���"O^�(�n]+L�-�⣁�"��U�"O�y�f���sP��9" �z��D"Ot��r�&fi��� ��/���H"O���^�����Xi�]�a"Oh�;�AI�9���83��>|�!�"O,��O�&-��$!�g�<���"On�ɔ垭0��<iRf����(v"Ox!�'����|UD	^)���f"O�uy�e�z����'"ИP�! "O.y�C�އv�zT�%�X7&&��;�"OJL9E('N�J����1O�ͩp"O�Ç�I$x�Ā�I�E��01s"O�d��K��2����@�	)f�(���"O���l%N����$I#<U��"O��8u)��M�P��r��%�y
�"O�I@A�=!.ĻîQ&|��"O���P?/:��Gk��Vq�"Otx�׉�o� r��\�6h���5"O����%j�Z=��q:P�a"O�
Ӄ�>�\�	b�2?o�urB"O� �����B}pQ�UG�=9A���2"O�x�3'7 �u���G/(�h�"OpI���8)�&AЃKY�Aj(:0"O�� ��<I�F���	Tv|�"OL{&�_�6k��z��3.|X���"O�e�WaT�X�T�i2��	@�X�C"Oz����Y#�LE�_.l��k&"O�Iɴ)�81�2Ua0����$�"Oe(����t� �Ƌ�)��y�"O� `�_�Y�  {�S3b|p�0Q"OA�E!:��["�ܙU�`!�"O̽s.��t)���.;��-HF"O\{t��A�f��b���v�b}�6"Ob����T!�p͗-`����"O�Щ��$^��!"��*f�by�"O�ـ�đ4G@0�$/F��\G"OJ�
a?6�� @NE�Q��ܒ"OZ1H�#�;EN�(�3k�&}�c"O��ҷm�5nNȐ AЮ"�\�(3"O��qg�:܄�����u��"O�%JAG���q�Ǐ�yD��"Oj#�3�8�S党KM@���"O(�S��Y�8�\) ����G0���#"OA�M	V�"�Gk�8M30�"O�@F�>,~W�+v�����N�`�<1�Di��)s�����`�N�e�<�eeBE�����
�L���`r�	\�<��R�}O��y%�A�^y��č[�<�Ɗ^�ea5��A������%�V�<��Nܐ��]��MN�]B� "H�<�bb��#ļ��/�:f3�N~�<�E��?C;�|�s��8m8�#�iPv�'�h�#�CO�<V��� �2�U�k���1DO�,�B$"O���=|�5�ʶv�����0O*�sA���X��dcO�"~"��֑�l�3GP�7��S5�y�<��]$}Ϝ�Ve��|�R^qyb��r� ��u�
y�ax
� $��F��<j&i;�dG:�4�6�'8�,˖	S-l�>@UۉlV����0e"�M��R Vg!�D�ax�d�bÐ6X*����!MQtўع0)(���`ԭJ̧�����h2,4X!�il~݅�a���IWؾW�<��̉�*�H<�Iv����@� I͖𖧈���I��й[qX�c��k�p�[L,D�Ă��? ?����(ۻf����C�<IJ��j��:B
�0<A�k��LL#��J5 �x�b$�FoX���f�O�kA����D�
���-VR��QHS�*��i�lV>~�L�BO�1��#�.ߊ�b�[h�0���>ID�6��iB!M�$�t�� ۰v@�c>m�'�H�Y{m�����j��|8剠L32X���Gj����3OF!�]i����b�4� ��G�;�d��Q"�$O �)����qMvb>�9�͓sH|��s�#C6������@��ī�T8��	#A0��+�L�b0�9BT��t:�+��7�ڜ��i�D P�*��O�z� ���8�t8sZ��O���)�b٧|:t��
�3"tdx�Ó�0u�!ʾU՘�'����b��n2L��Gg��Zxw�݀l ����)}p"�S��?���8�"8��
<J*\���[t~R��}�J���v��}M�(��Iϑt������w.��I�L}����l�#����I=���zT�N�%e�N,��[��>�J.L�@��|��/I�^��' VU�|��"R.��aꑋW�3��xu�'�d��NIF�Qȇ��LD�IUF�����1��E�	�I �%飨 ����~��XO�1��" "~��q��Lx��Rb�ش�Sp�>���J�-���zJ����+x8�hP0j̸��Q�"~��1 �j���0B����KQCn�Oe�P�Ugѕ+��ҧ� �Ǐ�>tVdX��K ���D�O������uy�@*��&,OP<S�'*nܲ����ש2��1���E���R`@�[@�-�s�"� ښʜ�0�êx�R�����Ѐ��W�Ҿ�x"�ëglԌb�흈%=��@a��v�S���)7�qO�![Ӧo�F"|�"��\\h�@����5���wX��(b���'��"��oۼm���N�,�
��'Y�Iʴ�@ru���ǟ]�<LS�'Ah)�"�Y$["ha�JV:I����	�'�jt`�C�X
eӑ��"B+ja�'6,	`@'�$
��`�e�/0��=��'rl8��h[hl8cp�Z�?A�	�'��%ѵg5"���Hf�@?�	�'E��x�MѠ 6�<�N�4&�=ю���v�`#M�
� Akʟ�ԨUb@7��QSboW��T��b"O��b!O?:��d�
�QÈyc<OHѤ�O���;e,�5�ģ�3L�Kh�I4�",�L�e�^n8�<B!z���(S� �*�1qi�1*,���M����� cGQ��d��rZ>�<ٴI������À�V8V�0���l�'<Ͱ�ɓ;��'2h��+R$q(����F�I��$���^>rR�ȢFjY�ex��Dj�RX����o÷v4x��%��h���a&���Z�8`S'#����ɩZ��]��ǎ�0��m�;Τ�λy�57K�HpB��c'	)����O��i��/�s�6Q0�� :'��͓l�6P�*S�#�ٳ�]�Mîa�/v�&I��~��AW�]H���G[ 7tH�f��=� ���2fN�8�w�|�� �2Z�H��W�� h�`�CF+�%�%/�zRAZ�F
#2�3�k�V��D�6����I�� �6��?�B ^ل��U�9� �	0���
,�hhl��'�ᢠFK38g0t������j
�H�p��'F�>A�.������,��KF�{n��;�>A ɗ�ʀ���U'�V��a���ywR>�ִ�!E�<�%3t�Ɂ�y�@X2N�� ��f��+�d��OO�?�TH1x`| �҈G����1��'�� �W&��(�`�:Q�W"� 0�E�6��h��'[p|�@o�%�>Uoڻip��(1� Y�|��n�Q�Ȩ�&ǻ��R�kX�s�p��5�~�?��+�9T��мI�����K�U�'�v��aW�r5���@���#Lr�4`��g�Эږ��9S���H���?�cm�+$�Qt�:{#4��$��?�"E�b��_�Ӻ�B%�<���iGO$}2��=>ä��kͶ%��ru�F�-!�䋯3� ��!%��B�0�c���M��	&��u��S�)�'d#n����ȗp�ڱ� Z�p��G�����MF�E*g��@�	�=9C�ˠ����
�d�����d7��a�Ì!�T$��(��g�w=�99u���>�!�� ������vb4��"ܞ2�M��"OĜ1���#d��
u���>��sv"O�Ka\�nB���p��;^�.�1�"Ob%�����飒'�x��'"ON`q�&
�h��81�)Ͷ.���5"OHp�2
�o�5¶G�`#��e"O~�2�\�h��,��å	|RA!��2�`�P���% <�B��
.5 !�d��!ϺAq�� ~!��#Ȅ!v!��'e�>ܢ� �^*���EHK�/!򄂊fK6 ��L�L$��@gɲ �!��<&�)�!OӨ;cfE�g�x5!�����ER>v=^X���\v�!�Z��̑Æ�.(k���$�!�d�0A����φ�f�� �AΘ�C�!�d�p���b��*O�^�c�/K�D!�׀��]��핏s� �� ��'�!�?=E�}ےd����K-�!�dV�0L𩣋��c�����L�Yu!�$G�R�xI�e'�ϴ�+�m�z !���=����%G2z�$�Q0l,A�!��-HI�� C�LcH��L?Z��'bL��HX�h;��5.Z��ŋ�[@����=�O`��&�4<�H1%�K�EbVTaҺ'@2!��B�'�4pɐL�#ok��(bF��{Rˈ�d��!��&��Oeެ�G&ŗI� ��-WA��x�'�P��#�E2_��Y�&C=�h4��'/��
��K%4�)�O�>��!OŪ,�9r���T1 ?D�0sG�� C�pS'�cjJ(��c:}�+i�̤ ��Gt�(��j��u�$�w,�o.ܓ�*�O ��,��ࠊ"��=�n ����B���N��x��/o  �� �_�A�x$�gG�ܨO
�ʦ�����	�����q����GL��>S�jb́�y�B�#^1���V�,��̊0�&�~�
 �M�T��D��S�*$<�����q�¬q����BB�I�����tL�8X�ƬX$kQ�oP�'���i����$���I`І��E�;GD�IX_�"��$҄&Ū���Ү���	� %�n}��c�i�,C�	���9Sv�z���j����z���?!�Y�S.�c?�X��n��iϊ\����qF D� ��Ǐ�lݓ�NM"G:x�Y�3D�T
RG���H�d�	Z]�`0D�Tj�j�>��[4B�����2D��P"ד �F�#䪍�V]Ԡ��`,D����ǬAV��<v;���a�0D��Sk�|Q.�qO�Z���c�l.�9�RH�7�2§fFԑI�l�J�Z�wN� ������h�J��U�fİ�d��Oܖ��D�V1Bf�����S�OZ�B�X�g`U(V��/ ,<���'&"������=3��՛Uy\$�*O8�r�,P
Ti\�y	�P���iĖ@��U��'�/�f�����-�vȠ�吉����Μ�t�\�����
QO6�b`H otJAB�M�:~�m{����(r ��P���p�	P�U�=�Re3�A�T���"O\���n�*�0�!Cȷv2�����'����	05�t�O?�;�n�,�~�`���.�hi�GY�<��L�P�1�U?W}�ͲD�_SybES�D�9Fk�EX���LN#�(D�2	��[�n	)�
&�OjVJ��N��pr!,�Uڈ!
���iz�i��&��x�g��Q��	�@�
�K� ���$�hO�ÈT�s�<�������c��p)A���0��r.֑�y«�r���&�B�,��)ч%�3�y­Nng&��|��	X���{p�Ag^z�;L��+M!�B�F`4�"�(�	4��঩CU�� l��m3LO� ~�J1�[�S��z�#�c�V���"O$��Mϧt>����aŋO�^�"O���E	���;E �O�ZM"OV��W�5a�}z�]�.�b�!�"O�a���Ufa���֓Q�tI@�"OV��3]=��3C�M�h`R"O8�z��� �!�TĆ 4 (j�"O�Q��,k8y�"�����Y.�y�]�L���H(TI���[�y��&_�p��V̍��dzr�ԭ�y�N�<�ɚ��	$�<11����y��M�3U��A�(z<:�#7�I$�yb��k�1�!p��1 ǣK��yR�� :l�ds< i3ˋ��yR�O�Gnu���Z��l����!�y2Κ�l�R	�3d�^��ݢ �Y�y�`�D<��J����\uʃ�y�f�hB�ܫ��N,���t��yBB@�Vt�@R�GR.R�l�"���yc܏y��,�Ð&`��#dϗ�y���%�Jy�"�>�^����[��y2��/jȞP�*M��h�c���yr��A�0`��Z�=X��!�y"i�3	�.��Vk�+�z�K�.�ybN���n����˼�^E���y��S�n_>y#��v�X�#���y���]�����l��e������y��(j%�[��4Q
�RH��y�ƛ^=���AS(�Ȳ�܈"a�E�5cK���DE�DjӴࢉ�)�85X��թ��	�%	!JKR̉CS� ��n�-H
UZJ|֧�$���8�l�[�H�8�A&�I���Mğ ʮOl�G�T�.���o�,y���_����>	5�)�)����'T�uM���52��'�"=�~Z6Gߴ8�<�Q� B)o*����o��ga~�ќ2�䬐���F�C���yRi�	-��{�S����Q ˗�0=�	7�I(f ȝJ���2�&���/�2T�>�j��)$��O?('LН~e�a�t��]P��#A��!0���O>�i�Ӵ�ޫk��q��o����NZq�'�#}�'�>�3�F�zΨ��� ��zjh�Ӎ���)�h���k�dJ!����
�sPT a;�a�����ذ��cX�|a�*R�H��=��_D�	�@���TgH�h��Q���G����ޟ0��D�S�OT\��`��x,�����n@�V�'d�W��p��?c��6oX�,H&eګ)D�i���[��'m�ɟ0�?�"� B4�PC	5�� (�Iş�0,(�S��bM�~â����H��SÞ7�'��K<��lt�)1�	�:)\Qq�l��I�2tP"<E�T"� X�,�.P]��a�O$$@ ���혧0|REǎVa�!K�&�H��&���!Tv��<�6��P>�!CHhώMJ�������W�+�I:����G�+����,�9���B��>��	�d����5�?}�O��F�䍇�O�� iaջ.��ɄkN��M{�i��$,�r��S#0�r�a��[ϟ�>�	",؋ī�z����Q<�"��ȓ&��dɔ�i��4��KޅyV����-���*���!x���Ū�RY�ȓ(�)�c\0!F�	��	�X4|��ȓp7�H�"�5-R��c��	䘆�>����D�8'�B}ۦ���s��ȓCPaP��.M6����,�ܠ��~����gf�FX��!W��{^2q��q	"@)�%՗3^Dp�d�\�z���S�>��%��2mn�v#�=�|��ȓpc�CG��Hg<�H��@�?�t���S�? �)@ʏ��B�q�㓢f��(K�"O�%:P*��/"l�CD�-���9�"O��;�kטV�`�'�����mR�"O��k���� Xɢ���o�<ѓ��-X���"��y��+��Ne�<�@�&:�F���e	�'Ξ�#�c�<�VE^&&a�IY��@<"���n�]�<Y��^X���	b�9x`����S�<yhW�Eb�l�H��^v"�b@!�L�<4O�!^߈��P�C�TT���T�<��m�@� *@#�y4t-�DMM�<aC.��$�#FѼcꚴ��hH�<��Aʵ2��M�#�Àn	"����M�<��GP�[��I�"��WC�<��.^����R�o�3<萸���S�<�UgЉ]xᙵ�	�E	�����o�<�̚�,N�Ч�R�y.���o�<�D�	vmN�Z��|�D����i�<���:�8�چOX�w�*ի�L�<���[/	���HD.�%^����I�<�!�A�Htc�(�3NdI7�U[�<Q1��} �-��IG� $`�"�L�S�<��5��xF,2>��D*��G�<�$L�^0�SR��������HD�<��CD8x��'�Ȩh�����P}�<I6�̒y�Nq;!��X┝Ra�u�<����.P?����N�pA��4C
W�<�F�՝T�у���t� ��T�<���Ӽ��C:rH��DI�<��F�S�zEYB����Y;�B�I�k9���B2��I�%^�xB�IT����b�V#�1�(`z�C䉼%C�ћ�J��ZЈ��${3:B�	�{��A a蓯?�BȁA��.B�ɖ<Ҙ��@�T�FP�Ŧ-M!�C�	�hY�X�!�^�=����GrC��0&���E`2O1�i�" C��B�4[�L�$�;<��1�`�&~��C�	�l���HA���4H�e�!;z�C�	�q�A0@j�/&^���[��C�ɂhO��B�Drj$up��>�C�[�rp����#[�2�BT"�B�I:]^F��EK,�� �'��tB�I^^f��0`ڈB'c&R{LB�	�V��H&W�Z�n��&M^�uN@B�	�L@vf$;MdQ3�jT�B�I�g;F�I0�D����cFߢT@C�Ib����ҩ�+T.���pM��mlC�	-?���
�u؎X��)]�C�ɷ; r���P�sS��Z��B�ɟ
�X '+S ���`ΤC�B䉄*��b�/G�,���7l]JB�I 6��<pvɎ��H�ې�Kw16B�	�-\�����ә)a
5�6���m��C�	�x���Y1a�\���A���C�Ʌ�pٺ�.�8H���Rd�*x�nC��3��P�N�'/b��H�|�&B��<[�D�s!T�w�P#V=bq�C�ɗk'D�Q�ϗ!�Z`����"�C�T���
��>���Ȓ�0��B�ɗ)�rS�̈́��.D�I!|ʹB�&8� �o�F^�cë�N�BC�I�\"���)�'5�<�y�a ;Q*C�I=�Ƒ:B勼j#(��3ҖS��B�)� |�Hv�"t6��be��9'��iY�"O����/��t�g�A�X���"O�3S�T{�<2E�U�}2X�`"O�4#�n�5*�|[5)E���"Ob�23a@%ƅ<(�B]�F.+�!�d
�`3~�h�h2�2��$OO�
�!�Y�[̖P@3d��>��	�p���2�!�D�%I��]{s��#E�4���/��@�!��u����Ҭ�	Ū��c0t�!�D�}�8L� ��h�xj�Dȡ\�!��Ӌv��q�F,yYr� ���8(^!���E�R�$�˷��Á���\!�$ &��!�A�yq���E(5?!��/�T�ԫ?`ĈrN�(_�!򄗩NL왹U@�!:j=����V�!�î6�I���+������R�!��.놄�	�4Z�*D�JI7:W!�^�_mXQ�05� !�r�1NN!��I�kT����+Nh��{��<6�!�[�EP�H�j��O�2�سre!�$B¤�ꌽy^~�:pBˣ{k!�GD�vl��� WQ0b�]X!�d17�hy�J8;8����ը;*!�0c}Xm�t
�+�lx&$J6A!�DE�h�9��%������m!򄅓o�ܝa��F	��=yV�:�!�$НZ�* cЮ$�tt��7�!���M��b6�6�B����G*�!򄐩j��1�DP�\��d�u�F$V�!��	R��T�S��I��\C0C_�I�!�D�ț��v+��a���:l�!����	
l�PWi��PpҲ�݀�!򤑼0Qv����#T1�A�8�!�G�'��D�e�\	r)�v�J��!�d�'�~%2��߉MN�r6b҂.�!��r�n4B��Q6"T �kH�Tw!�d^�T�(��$���b��_<i!�$�M� ��k¨js�]ɰ#�8QY!�D�e��A�pe�:Y P�$#!2M!��^:�"�˔b�
_T�=��'�!��X�I�5 F�@GB�cd��(W!�d
�J���S%(�A���y!�$������ː�|��U���=j!�䟺}�t�A��V�e��� ޠ4Q!�D��@����%I�4�U�n�5!�$_<�ΰ�.N�"di�Β;\�!�DL�	�fM���Z�Mx��玅P!� �B:�K�ʌ�MT�=['G��M�!�d�>��{v�W�!�l��ī�n�!��ѻ(�P�`����N����)ηA�!��T;?H,��j	�u~�B�\�l�!�d[�MW���w �����G�`�!�$D�l�N����e��[3���!��S;���#�X�h��ナ"�!�$�)@" � ��A!4���Z�sw!�Y8z킢��Y�>�
H/go!�$:v��6�(~�.)r���;2h!�T�+WX(��\��`K�I+!���M�ӅTq��ǣ����ȓI����� =� �� ��X�ȓL�J�k��I<;����^����@ā��.͊pp�q��J̧g��	���z�+�˖\��2�,<��OVY�<�5O�R�Xc�͚cl���[�<� ����v�����C"0��#"O�}
���m��@���M�a��"O�@��.ݏ+B&�2eɀ:0I�"O�U��c��%y�����  ��f"O�(�2��67��d"Eș�̸�$"Om�O?�	� .�,	��p�b"Oڤ� "N����K��œ�d	0"O�-3Ş ��m�!��h�#""O�H����/l��q��+t
�P�"O�AKDm�i����DK��;���
W"OTY��K�L׎��J�<B��"OX�*�U\��Tѱ�@�K���"�"O0U�j�~������x{�qi�"O�Rp�N�lL,I�A� d����'d�t[����aUr�<k�&	�'�0�J Aցt�&�� d-V����	�'C��a�Ŷ�JM@��U~�)�	�'�F �$��p�
@(@r�4Z	�'��ȡ���ve�P�o�?f�		�'�FEhcD�	��%c�脈�'Lx�1Pi]�(��
ȳ_X�,
�'�4�Bv�ˤ� ��b��T"�ĳ�'Z�����OR�e�1�WR5����'�^����!D����@� <P��'A@ԡ�-�{ͮ��4�	s"��
�'&mP �;�dQQ�5o�6	
	�'i���·j��A[PgT*d�<�)	�'ewH��ZـA÷N��c[�l3	�'�Hq�>_ޤ#��TyD��!e%D�\��X�
�� h	�/d�P�(D�<�6lY�Q��5��������+&D�`�b��|垼p��&f�l�G�%D�(��^�U5��"��H[.V�4�$D���s�I�b%��!��0w��{�j&D�h#P��2V�� X�Ç!�N]Ї)D��+w�J�B�Z�I`��{\Yz�o4D�ؑGE�Y ���t���Լ@��=D����*��Ab"�r���6�0D��q+^'��mPbf�����G'*D��A`�ψY=�ʂf�����y�f'D�,� 	K�W���1�+�V�3��!D�t�E
�79� �q2�żH``�i D�Թ0����ذ�,^�D�Kզ(D���8�0T�ǡֶ�*�*4D�\��jR���\���f�F(*��1D�����X�>�T���m��IE;D��ALS!%��8 a��#2�鰂-9D�؋�Mԩ�0ădNLz��_�!�$2�0��Gf߭a�L%�A�$k�!�D�6�6-)q��!�Ɣ�#	Fi�!�Њ\s�]#�B:|�����b�j�!�8@+�(p/@*%J9z���,v!��<Mhp��<���A;!�̠	"tK'X�g���2��:!�D-4��T��g��X��[3�[1-M!��:o�$(�T2;��q�'�K:!�D��c(́�S�9�P;1�V�"!���=�N(��N��	&}�V`��o:!�;7߇l ��     �    �  �)  �3  �=  �F  Q  �W  "^  �d  k  Oq  �w  �}  �  \�  ��  �  #�  g�  ��  �  .�  q�  ��  6�  ��  ��  ��  ��  +�  o�  ��  ��  C � |  Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�� |d��"O
`�(�;���8���-0��1%"Oj4��ND^[��"3/9�0|H�"OB���H��*�ʞRy=a"O�味V�!X��!&F�:J�$���"O,��a
���C�Ą�M�"O,$3%o�-���p���+Ն�:1"O��ݢ1����`���y14]2��i�<�6��{_���c�H�`�fX�$Kn�<��A̼VI�xR[�)�Ć�pඤ�ȓA5��('nߡ4�� �)˩%� ���,��r�؊b#`T�eT09���ȓ!�b��g��}�8�F��-? �ȓ
K|m�ș�VṔ���2�%�ȓ"R�X�j�4JN�1�˘X�i����̹	_�jZ��1!g��zܶ��ȓgil,*�J�
j�Ne��i�J%b���f	�(U��:���G��$Y^م�~r�� S�%T"���k\�jx�ȓ|4�1�îJb��@ӵ�ݩn�V��/[`�"�v4�R�!ʎ<��M�ȓ`:��z�ؚh�J�Z��$HY:	��H��p�m�C1��!��B:��0��EnjZA V;9����J[
2���	��4'J�EA�IVW&��~�(aZ��ӹ�>� o�Y�|�ȓ�f�A�
Ο7�H��M�$�����mޠP����/���ANXo*�ȓTv�����{ ��-7�*h��I��sB�8�8���3����ȓNe*M�悡;������X�o��!�ȓ'lj�#F�m�+R&;�|��2)n�C��0S4���T:
b���:�0!��e֊��)��ͷV��,�ȓ0�&�8#���� ع�L�����;�P�AFd���,w�6d��r�EQ�( �gVlɦ�M,H��,DP���|�I	$G#\���ȓ"�)���E�B	yt&B�^�LɅ�	xy=Oѱ��Z��|X!Â=�x�8�"OF-���З[bP
4��
/�ȨPE"O��p�ɂ�{��]� 'Ч=y�l�"O��#�h�8)S��K�K �[h�TX��z� �G��*�=����4:Z�X���;D���C�۷F�Ƀ�^��Ӈ@=�D3�O�yōF�uu$��0��,�T�F�'����g��) !��<�� ��P�Lg�B䉖>}��R�I�b�����
O8�=�ç8���Y��ʟvd�HRQI�<�Ѕ�J��\C�ѭI��jXu\���  �s!]�p(�aqF�SrXP�ȓ2 ƙr���|�#�o�BlH�'2a~B��#!��l��M7w[��`V���y���)h���eE�sv%�f`��O��dE��ʌuH���Bݽ\�;�"O���уO�%d@03�J�7�PxT"O����"�a��1�ubI#sZ}��"O�Ys&O՗4�d����q�~���"O�!r��^s�pz˚:�J��6�|"�)7r��a�W5P�"��$\S@B�ɗ#�P�[-�?4���&E��7m>�t�siUЌ��GO�eܜa�!?9N�(i��3� f��� �IyԙI�(�h�j%!"Oεsv�4S��a�ͳC~f�;��i-ў"~n��L+���F�)?Y���DN�:�B�ɯ.Z�h��ߧ�=p ��
��B��s����B�Hh<���%����:�� 6�a���/Vq��5@+y-T�<���'��U��ʒ�F��T��,���{"�)�)�y��L:��/uh��%L}�!�C7���Eb��P�:�����I<@������k��:ZuVC��0.�4�� �KA��1f/+��O���<b)J�.(YT�4�P�N�=����Yyr��`أ$���㣢�5y��L"��,��;�O
����+A޶����0R�>Tۖ"On���p�t��eDH�yI,%ळi���D!���!w*O�G<�#�O;'1O�7-����'��i�|0�W)Q{ҕÕ�H�Ѳ���\]�<)'�<��)��QL�j�6��V?����O��O�Z�f��(�j���aŵ�� ��'�'֦tR3IG�9� ��C��k�A��DP>��wӺ�O��7��2>�������X� �2�M�B䉵P=*!�7Ɯn�]Y�j��E=�C�	�5��H�@ݙD��1{1�B�����6�0��͜|�f@���:.���+�O0�'@\ͣ���-~1�'�%G�8�'��d�D�ۮ=��4��!Ǧ7�n�0ǓXQ�(��a+��VB�~�㕨����'�z"�\��IɷVȶ�`k]�5t@F2�Df�2�ȁ��)'-p����ݺ+�!H�b�<��W.��%���U�u���[�"E\�'ɖ����\~�"�<(�h����!Y!�^<'�<v`��e!l�'�z!������hO�O�&��S�._�$B�@�|�d�B
�'�J��ƫ ܬm���C3�� ��	��<a�I=Xy�d*у�0C9�Ѳ�lYu�<1@�H���R%)�|.��Z�o��!񄆨k�������73�U+U)%1O��E{J~Z��0.5f(ab![�e�2�2`z�<١��W�~��B^*4�b�ᆈ�t�<1�bA�]}�`r���xP���G*p�<�vM��Z�0E"5R#h˶!�6�k�<�g� w6��@%@�}_�1KdbJr�<�4&�0 �@}�&��&�r���J�W�<�-�KYdmjd@�E�\�2d�IW�<	SgY> ��!�0m!��(W\�<�d͒Y�����˴�0��A�\�<��Z����6r�Q0��ۻj]!���	b�N�a�7�(K4�+y!�$(�Ȁ��?&��吶]�!��.?�&�(FMSe���3�O�*�!�D��E���& ����e."`!���|���6���B�J���l� ?	!�dL��*��XP��J %�!�'%���cX84�1ɢ�Z�t�!��'[K��Q-֖hs�%P��\/�!�� �G�%9��qwVuP�!9�!�L��4���_�e�م�6�!�d¼w�F9�0gR-IQʨ����^v!򄞄^��e���س[��ec��K.f!�$�!]e��zF�φ~¨phg�ɄQf!��;cN452g�*��Gf9g\!�D��&<���c�ӟ�f��w�4T!�$йCor]c�!B鶁�$DC�Q4!�D�t���T�ۯ-�Xt�BDO6}!�� b���mgj���L�C�<���"Oz�P��&ne�8R4kA�(�p�jD"OJ���H*@xIg�Y�9 ���"O�YPOI�K�Dlӱo	%i	� h�"O,�Y�!�f8��a���> �� �Q"O$<��l��Ik$���2�"O�mAŦ-*yĬ{&Jz���#"O6� ��v,}jdfC�1�u��"O�arbC�� her�cX1F�Z"OB�K��C�R��c�B�(\�ơx�"OH�1��W�&e���E�].�L��"O0Q�'K�7hH�YK@B,���"6"O���`J����D�����"O6�y���gŚ���G #��ٗ"OeS@ � Q@@��BĉwY�J�"O���d��U�����n>�cU"O���JF�#Ҋ�� ږ|��`�"O΄�M�#)��P��m�z�~���"O4��҆��$f �w&���=�p"O ��D�?yN�4�PD�PJx)�"O$�1U.Z�O�\��IͅC���JT"O�1��:L��C.��u��"O�X�W�U+\O`��@�X#U � �"OШ�&�ʉ`� �&ʀ8K2U��"O����O�V-Y��ڨ?<Mɶ"Ov�8�e��P^
h
%�tq�"O2���C�55��q�Ń���%!1"O�H�i
���:�F�'�Ne��"O�;�O����e�!�Ht�T"O�Hb"�� m͞m02B��L��у�"O���&�ųK�d�1��M���d�3"O� (�L u�40�Bؑ��9Q"O���HUWzH��+��1�
 "OZq��h�4BfAS��ޚP�`
�"OB�����&]�~��s�[����"O���0�;�� ���φF
da�"On�c7�X�����ӛr�p�"O6a(W��P]z���ݬ��!h�"O>$(b!xd ��`�[{�i�v"O��f
$��Ȳ�%�2Oؖ�T"O��"l��:z�) kևC��]�!"O~��r�1JJ0�{ī��-��"ON9i�C	-�QA�ɼ(ID �'|zњBc��_� "�ݘ#��\9�'�y���Ɖoҙ@���=m���'k|�pF��c�t�b�1jE�	��'��H�K�r��dy����/)(8[�'�d2�枎��!P����o�J �'�#�Fܐ��C��|C�'ȝ�rHݠd25��V5_Q�E�':��
�@J�/��`��.	 R-dL��'�����h��t��a�)	�L�����'*0@wɛ
��0p��*o��!�'����3j͌e�� �H�0UXTDH�''-���G*��4A#�A�M0��I�'T䬉��K�=��ċ��ښAʲ�ʓ	����UE���t�)A7#�h9�ȓ	<�Mk�g��eC�͚7|'��ȓw2���@�ULkGXH��Q��7�@�rFK��z�)C�#Y6�Ň��ؙj�cܢ	�P�Z��93�ȓR�(����*j�$��Č2z��\�ȓkP��e��1^<��R��	�w�D��EJ8�F	s{��JD�ǧ2ظd��S�? ����n�N���IĵE�"AY�"O�Mʷ@N����
�>u*г�"O� Y��.a(�J��Ɂ!Xp���"O�m9�N�|��hZ�}9�5��"O ё0l;���t�Թ����'�2�'r�']R�'R�'�"�'���p�R�s��b'��>i�$�t�'�"�'/2�'e��'�B�'��'�x%��-��ȉ�`�3P�{q�'���'V��'	��'�B�'D��'�8)��T�wjq�Ae�l!xf�'�b�'C�'��'E��'��'� �0a
6�)Tˇ�7T��T�'r��'���'�'"�'�'��y1�F����p�ҷ.�h���'�b�',2�'���'��'���'�����Ĳ=���堍�q��u�T�'�'5R�'b"�'��'���'	�#d�!S5ha��B�`�5���'9��'7B�'���'#��'b�'7���+���"DrƊ�*3�pm��'@�'W�'fR�'��'���'N���o�8[��iq��{�R�2��'�b�'���'�R�'M�'�"�'�.�R3�F��Ls�+M#^��-`��'��'�"�'?��'���'�"�'�d�EC~Խ"5��i��K!�'�2�'��'U��'hR�'���'�2�R2��2f)C��4C��ػd�'���'���'q��'�"�y����O�`J`HғT!p�h�R4�HhTfy��'�)�3?Q6�i=D����Z{�����"]=�`X��@���F���?��<i6�ie�jp*̽''2�j����B\�Rjq�d�d�3\�7M>?��
�/�05 ��O(�@�+��@��̇��8�B�y��'��{�OV��kS��v�I��s�B�	B j�����*���M�;�l@�-I�Z$0�X�TƂ1���iȰ7�`��ק�O�t}��iZ���6X����C�:x��6��<&Z�1ą�@ުDӼ�=ͧ�?�7C�;s�
�F����,��-��<9/O4�OjaoZ:��c��S4u�fGњV��1���	2|��?��R�T"ڴU���9OT�c���V��/R ��o԰c�L��'��zvj�+j+������-)V-�����
8��|�򈖠2�<EP��Sy�Q�@�)��<)%DD�)�vFC�	�^���@��<��i�ΈH�Or�m�\��|�t�M"1@ΨC BW�1��p���<�i�F6��OV����nӾ�1�ٰ�ʉ�Mq~$�B��n���7*^\�����jǾ%\~�r%�V�K�85��.�5Є�}&�@��D�
<�f�i�O5x"��m,D����/d����6�T-Xp��:���2&��|����օk�hS�J'u�Dl���"�����&����a��m��1c�aD���C�5m��yM(vn�pq�^~�T��g��A�\Q� dA	+�EA��D�)Uޤ��H�A��k"MU�x&y" #
7R�����.�����Wr�T�d�O�����zL�'�
`x��Zt�M��(B��ٴ�?���E�}����S�]A�ek�h,Z�`�H]�W~�al�?x� ���4�?Y��?��'O��'�"-��O{fu�BaFY��Tp@�
�MX6��/q*��0��ן��I��҄g\�	w����G07�o���ٟ(��=�ē�?Y��~�L�5o�r�{�@�"p�L�Չٜ�M�N>ɢeA�8ωO���'Sb��|�4y� B(0���/aC�7m�O�I���s}"�'�R�'�ɧ5fݹ ��yj��[7X��X�Į��Mk�7u2	K���?���?��?�(O����
�X$�`ʗ�y&*!N߯+�*TlZ˟8�I�l�IAy�'���'Q�x(S��)tuJ8��$Ǵ{)�3qH��B�'GB�'��Z>���R�	�4F��$D"G����b�4�=⓹i��'��S���I����	�/������ [�� &�?q�2P��
���4�?����?���?��l˞Xp��i��b�`!�#.�� ���x]�F�'<�'�R�'_�@r��'A��Ș7�Ӑ;�� F�{�,Dm�ݟ��	|yB���k�J�f���z!�����)�l;xx�E�IZ�Ο��	�FՊl��W�~Js��>g���M8;־�X���ʦ1�'E���FBf� ��O���O�b�Ll ����^�Iz`���ϠY�^�mZ���ɑk����j�)��=�$�V�
oA��Y���-��6˕{�,uoZݟ��������?���E�TM�<�h!1��y��HSh�6-�,?"��O��R�'�?�m4��ۣ��{@�CEjP�tP�iO��'�Bl�)�l6��Oʧ�?Y�'�`���O���b��!��t�ش�?���?aC���*��՟��	˟���(���P��}`�H:F��M9�ml��Рr�M�����O���O
�Ok,��O�h4+T�D�iS����� &,���'���r�'���'��'���'Y��	<#�H����"[��ȋd�	�g�>J�O-�D�O����OVʓ�?��Yߘ�f!��r�|<�E)f6��;E�Z��?A.O��$�O�˓�?���P8��$�$yԉ����1Vʡ�0�� �M���?)���'��DyZ�i�'F/M2���-�k�F�&���IQy��'� ��A]>��	"M-���P���af��$$X�vH��4��'"�'�@qz�yr�N`j��D�štJVl)g���x��7��O�ʓ�?�m����	�O����k�A�͘Djt�߸
	:la��#7�'��'����D�|Ҙ~� hX��팪31h��/aִ��1\����'s�`��	��ڟ�yZw>@H$]�ioX���`��|1ݴ�?A��E�>��<a���I-GH*\�O��ZJHщ�lZ6t��&�Nler�'2�'��DV��GH���@0�����n&,��i�d��|�9ҧ�?I� ��hG�	3�[.X �sȄ��&�'2�'�T��/6�4�x�D�O��*���d(h��� 87���T�	��̟|�	�f�%꬟f�'�?��'��TXd�Q�^�L����B�x�ޙsܴ�?i(Y���c�����".��@�g��3R8��#a7��m�ԟX{�� �i>]��ʟ��'�&�A *�TL~|�B�Ļ |���T��HdO����O����<����?�t�S9F�r��4��Xdb���>to=����M�T�&U�w��'f�(FN#��5�Qw��zf8i`� #��YGZO�;e�]a�i՝	�x(J5f�% � ��.�ڸ'K��HW�N��d0��)6�ID ϊ~9��
tKM�c��T5��5��4Xf.��0\@ZGK�[o�-3��N�o���
*�>!#�c�C����Pg����AɺA�`��!��w�|mÇ���k� �T�f����O�1r4 i���*q�N�(#�e�����! ,�����?!�-@X)��V�]�uo���?��c" �{�&�2*�@Xԫ_N��z� P�O0�+�:4�a��7��ۢg��F�De	3�>D��)�5�dvS�IX�fT>U5��N;�֤>XN�xk�cBt�(4S�KM��ǅ8��6���^G�9��M"b��]���1
�'�r�R�,�#y��Z虠�����0<�a�89�t���蜞i3���U�=^j��۴�?���?A`,�o�Z�0��?���?ͻ6k�ږ�"H.@��DV�nn����>]�R("�'�%��f�����~% ��ӁD
c�����Ϛr���4F�s����'<$��f�g�Ɏ<K,�S�
9~�}ܜV=�L�K>1V�ݟ�>�OJ��H�;�������Z�.Y%"O����a
K��D0��Կ9���iW���r������0F,����dd�J)PC�O�x�:|��ԟ������8�����q>=��!�wI�(���G#*@v�S��%o���z�A�`�~�;��Zfx�����I�n�l���.�$,��6�M,�\$��*�7���S�FGx�,���I|!���Fʙ,#��xB�D�	|F��DN̦��ݴ�?1(O��D"���\W�M�sH"�td���H�o�nB�	��t�yBlϒsKF���OY�"{<b�,	�O(�f� @! �iF��'��q�I�T��D`�!Q�%�J�Z��'�2���@�'��Eb�(9%���J#r��!�çJ8V�P���k�(����'+�Qyv�M�>�l���˼O�!F���G���1�v�i$��p<�fbğ�%�ls�E�*.p��E��5)���)D�����<E��J�S�w��0&:��Z޴F���H^?'# �q'΄^mT�<	��Y]l�f�'��W>B�ៜ��@Vd�V�b�cͿ��E���N۟��I�UVl��T�S��On��SH�Onj�#�Ԍ,�(D{��>i���+���(Ő,�Mh���Q�'4᎔2�GF0* .u"uc��> ĤONL��'M~�O�0A@`��69`�t��#� �"O^1�% ʆ,ܡR�W���K��'��#=1�
z���I�`�#�<9�� �2r���'k��'u�h!�����2�'\R��y�mT1w �@��(A|��n��=�1O�p`��'�\�S�@�G��9�@/P�mop\�{b�ĭ��<�"�ԉqAH��� 9��*�aS�-��'��
�����z�� 6��K�����c@� �~t�ȓA�L� b\�X#"r,�(vy�'N�#=E���ޏ=z��w���C�^d�Gg�(G�,Db\���'�"�'W��w�Q�I��Hͧ"U�4K�.N0'��ax%��qd��Fr�
Eq�R�>Μ��Q�'�ш��D')�t	�g"�c2*�D��)��#�&e������*<O�-�Ez���΁)��҃A�a���hӰ�m���P�'���@���$��A?e�����E<�!�dX�<��.�1(�����N�L�1OPm�'�剺(���ش�?���`8�k�S�^�ZH�ƌ�6%����?	��ȧ�?9������^�rT�*��H�	J�	V%�Jgl�W���Q-1
3��s`�2'���Yʎ�@��A)z$��B�X�![������}+��d�
�@<�=�r*_w�'A��(���� ���c�b@�!���&㏊;�j��9q�A����;eu���oH
0\5���F����Q꼄�1V�X�E1.��'+l�iRbӴ���O�ʧoԸ����-"0pB�<~,�#��ۃDG����?��#�&�?A�y*����Mʅ	V>�$�I)��{V�';4�3�����m����A�v���K�#!]��o�J]�	���S���M(wb�	J$�$�Xܺ�
��� �� �H,VKT�9�%� �$���'��"=�T���>�B�b�(ߋ/$���<M$�f�'���'��+
|wb�'?���yW�W���)2�N,[9`T�%X�1O���f�'��J��Q�V�,�D*F�&tȘ:�{b�A��<!��ЅVo2%K�������0 �ˀޘ'����S�g�I5;SH���Ƚc��mѢL�,c�:C�I*(��
�@�p��	Hp儾��z��"|�`fA�\��M�4$��`֊u+۩l^���'�?����?I�����O��$�O�1�Z�.(XeyL��)�Ѩ��O�j��qD8�O�m)�I�?'AN���b�95F��C���<��ABf�09DN��$�$yPȂ��#9)Ԡ����==���p�'��*-��O���6�I:4ǖ��F
��g#�"��˵B}���%ړcͪ4i��7�$���ڌu�x�H>9ƻi��6�<q��a��F�';�d��;2���p%cq�	r�f÷+ "�'khlX��'a6����'{�'�	ӣ�� ~��V^�7�|A9
�% Z��?�$��9�������S�d(����K8�L��+�O��'���o�&!�V�kU��)�b����$D�頃�o �C�����i�An!��ߴN^U��-�\���i�b��B۔��<�#n��@ڛf�'�"Y>�����4���C�:���
<^�t`,�័�ɸ`rP��K�ވ�`��ʧ��IHf�.(���*99��:Z�:��s0�ƛQ��"�>�'>��, $���Ӥ��(�4l�Oj�q�'A��O��EZ雳^�����~pi��"O�!���R�iU�����L�8j�ш��'i"=�b$��ĔIzb*Ϻ\3�`1���.G���'vr�'�Irf��mR�'����yw�F��$����oY����#��T)�t��5�T�Q�Ï�(YbKd�I"�\(�Ɲr��hn��J�㐮6�#�4`���W!33�b�)�(��I�StpׯD;E�óe��Q#0�aH>��e����>�O~�"V聩U����6'ŭ"�E$"OP��>;CA�c��#������y��ᓄX5r9�-�"Oo�(@@����!��b� ���I͟��	֟ ���p�dz>�yW��@���	c�a��g�<��qx�,Z�Sɐ�m�H��EE�~i���E���'�a�d��[t��s`�	*U�R'�cfP� ��?A��?.Ot�/�	�1t�8��iֆ�༉v�ɛ'jB�ɬ6��티㎣q���q'"�0Kefb���O�˓E���i�2�'��p�Pc��>�n��h�'⊼��'%�H΀6���'��H���|�+�S5"-���bh4��`����5R؞�L����*R��-�3+'Y8!�"OF=R��'�fO*���H�p֌Lp@ Ǯ&*��"O���FUq�-YgO��1X�{�OTXn�����(�$� +C���"�-w��c��B��Mk��?�-�����O6D��L\�����g]�fx,*'-�O��ގI��e��@򤌘��]�:�(A�O=�ӭ:� ��Ԅ#��`� K�p�'|�����*��a�w��9J�P�s�Ʌ=��,���,%F� ��15��,\J���D�S��{S|Eh`�Ň���qo�33�����A,Dp�Cʓ�#I�IY�,i�p��4�mEz���oഥ��T�Z�{���?X6m�O:�d�OAk�� ����D�Ot�D�O󮀃�� i0$R���&C��{?"ف�gϺ=
�ЈD��u�̚�c�����\�
}ʡHƮ
��h*A=�"lb.��Ⱥ0��O�6��d��l�~�g�If0ݳeA��Q�d��i�Ta�!kN>)�i��>�O�ظ�L����\��ޓ)���P"O�p��C�R��q$ ?6'j!ju���ʌ��ӝ6ҵ�@-�8lG�8`bl_�I�@`H�h%l�����͟��	��Xw���'Y��]�c�$�.��9�WEΫ/.��4�ū���2�[0&�DƘ{ڄہJ3�(O��"i��Z+��Y�H�I��A[U��+�z�0w#Z��T�Dݨo@3Qo��JDR=F�D(}�6A�'ԬT���28�Q��8#^�Q�7` ��?���'�(���1U޼*��/��8�'�iBP8Z�8�p �͹Oȴ� �y�!rӒ�O�4��d���˟P�d��2f�!��a��t�4�S��l�	=MK6���ş�ΧE��A�	n�ɐ_yȭS�aêj2,`b��K��$�񤑝;��O>1�hx<��R�R=M���3D�'Ox����'7E���^�Z6����O��MZ�'bV1��I#+��Q����#N����'��6� 5�'���[�$�ӱΓ-{�:!h�1�$X"0�2%l����IC����^��9p��\c�H
%t�N���C�N���'�*�#D�T"A������D�D\�d��>t��)b�_>�Zǩ�M�z�B��vp$��k,}��� �4`0�
m��QP�oX�kg,�IS�4iZ�|��Q *S�at�p!1Q���`���$Gb�)�S�����Vo�<a��CGH�8�C�I��ֵ+GE�*f�hٓ.E�XON��D�F�'��A�a��I�$��lM����*��O��DW?&��@Q��O��OT�4�Jp�O�:?O���e�( %�4�$��+o���d�"�BM�G�Яv� 1�� vqO�<��'��ͻ&fӑ8��@N�K�H�C"8���K���L>�N��`L%#�H�ig�����Q�<�VhH0C�Ӌ5+�8Z�mXx~r�#��|RK>�QeJ�X��H�dܬz�Pt�we�@�������?����?��Y�n�O���}>�2����`I�ji����@!��v���r�ˉ�]�U�P�7`P�Gr�ƶ]H��k�/DUpB�)5*܍B���$4!��)v�ɓz�&��ɓ�ڄr��,�>�	ф��r���.�O ��	�.��jPe	'y<�ش��J�C䉰b�`� )�NH. (���w��c���ڴ��`��U���i��'����&\��h�נ�Z�,���'h���B�'��E�m@�Ek`�p��k�����I�T��1I'�T�a�^��'��!=O(����ԯk�`��b �:pm.8
t��$L�ƙ� պc����z�'�J���?�S\�8���H+�ֱ؂aG�t%�Նf����ʟ��?�O��I� ěB��2H�31��$J�ZB����M��
����˲�t�"�S$ݟL��W���4@��M���?*�J�8$��O��
�>	��% f�@�R�� KL�l�	�I��������c�?	�H�a���ʧq�΀�A�vb�ɋ��D��ܴ�ObX�T+S!z ��&�Y  ��h��M�6� �b�f����O�*p���1 ���UlJ�G��'Bdq����6KsӼ�d8�	��ذ��͵=�t ����(@0tq��O��d�O�$ Oj���NbH����U��A����0<y�i��6m4�DK}jb�����H��u#f��,Hw�l�Ο����|�uA��`����	����ӟh!Xw)�9C���>�x-uh؄2��tH�����yb�<�p�ڵ�Y,D)����FR��'=]J�t��0)B*,��Hhс%h���a�y�%�?�}&�d��-�(#ƞ�|�D���=D��ؐ�K���-��P	_�Zc�
&?�w�)�'IsTY���ЩzH��ʋ�+�
�(�mɔ4�ة���?)���?��������O��&?P	�N4{2�(
bg���m���� :�ր��I��0yi����/A~U� ��������%���FhdrApkRB�'Y�l��Ɇ Ch�=�bō�ց�!�?!��']b\hP C����b�^�G2)k�'8m����A��]YB�L"D�ı��y�as�0�O~,Pg���u�����J�25 �V�Ȓ>씛�B���h�	�`���	��H�ɲ T���Ʌ'L6
�Oک+��>+He��C f��]!�'E: 	�c*R�,O���kՏ7q��Z?{>���'>�����?y2�ik�D�<aS8�C��p"��f�M�
G�ʟ�?�|�{��YHĻP���,`���� �w<I�i�2uQ�K�`ð)2C���.���s�p�Ie:x�d�i�B�'��S+)Z��	�&�|�����5��	TI�9%cV���ٟ�b�%��@�t	2�`���$��S�t^>����ڎ� ��˅t�u�5�4}r��9������M�IC�D�(���(����t�B\�'IN`��N*ĜM97k^�D���O�)�2�'T6�O�6]�'�B�O4e�E^��n@��"O6u�v� ti;��1'�Lmb��'��#=Ia��+� �)6����DB�����'2�'�}�Qaʻ'��'R��y�I==��7�^�t p��s,�܊�D[5i��i ������Y�����Y��DDt���k@�Ih(,Q�̔M�D	�����<Y@��.�F��O����g�Ӽ˥	L�(�Ήے#Ǫ>i�t���8��'n�t��S�g�I%Tߌ\��z$�\���W,I_ B䉄{���#M�Ga$e#�����up���F�I����d Pi��#�-�3j�%�	����	���]w��'�i��N�l
�C�!^ḠY�
,6Ǩ�҆��	Yd��'�@Ŏ��d��?�T| ��4{�r!b$E�	��1��+�pmN	jV�r<Ꜩ�n��m�T�-���{҂�$W8��2��1���@�G�e��S����?y�&?��q��-Q;v9)UE�{�<y��Kc �C��IjiXw)@R�6����|� i(7��O6�� ���E��R�U8���0|���D�O��$K�4���O��S)bv�ց��W�@�%�M+���It�X�e R�h�mNC��x����aDH�UH�B$_�ztp=Xu�!\���"de�u�XL�ay��l:�,�k�qO>Z&�'Y�Y� �5fF)[`��C�=��{Iw���	���?E��&��᪹��b�A�LH��D��xR�~Ӗ�s`�@�1�X"?"�$;�O�Ojʓ{�H���iA�'�哥_���ɷED�т@��]��A�(v�I�	���Bg獑-D`U�C(w&b�"�4��i�|Fߵw1&�
�m׿-����IIO���2K?ڤ8t�W�$�$y���,{HXy�D��P���p�O�P��h���-�H�ԁI��S��OޑmZ�Ms����'���/��x��r1ˠ7�8gh�-�?���?��0<�ߴQ�bY�# +����Ȟ�Y�Ԇ�ɕ�MD�i�1O@$��BH�O�1�&*���S�e�V�$�O��d�:�1:��O��$�Of���˺1-֏z �� ��k��@{��� ��y9�4(�V6�ڶ��M��-$��D;����$�Ȋ]��ႇ�=e^�p( �Ӧzf��*�>|�ֽS'�I��}�Ne�.f�=�7aG>	�T)����=J���'�ɟD�(O�d(��?���?A�laN'Z3f���.���'��ybJ�?s�~֔�2�	ˣ��/���|v��io�z�O�i��˓3����*��Ex��9�GA�SG~8/N�1��g���������	��u��'sb�'�	�%��Aa��%Ȕ�U��9�q��^��� �%{玙�2<O�-� |��X)�I�mA��B��jk����iˑ�p��%#��0�9�&�O�P� �o)��OXZ	�'I��'��k�@�?p�$�3�'Zd�Ip�~���<i����'v�:��Պ7DZ`�$c�4�ޘ��'�%��! !e�\�`��"�;6�|�}ӠXl�Xy".�,s�7��O��d�b��p7�	M�� ;d }u4����?�u���?!���?G�`�0�z��F����C�lE>���K4h�l��!�;�R��I�]'6 ��KV���T��vz���n
& ��bumٜh��8 j]g�'�8 ���?�,O�H3���?t�9�mA5%�.��9O����O�"|:W�U�L�Ya!��87�J�J�nMf<�`�i���gj�	Z�´a� ΛUhH��t�'�ў�F{�&M1�fd�K	��h���%�y{� �	wi
�ҡa���y�/�vxиcf�uD ���L��yb�Xm��Y �O�2��r�.�yEA�V���&ϺΞy;�ȴ�y��h�� z�ː9;�(;2���yb�V�j�b�G�W���̅#�yBe�	O�$����h��&��yr��)n&`(2��?��C��H��y2 Ϯ)�U��㔶;tf\0V���y���
�pm�o��>{|h��+�4�y2OĎ��8{FH;/T1!���y2
G9W8,h���b�\x@	��y�6;�`p)�	�T�F��g� �y�(�����K��ɹA#X��GH��y�g�R�`S\�� \�y2G3`�k��ѝQe����e� �y��O�B�`ȧ��6KX|8���^��yr��m�<�Q�+,h�)��ԫ�y�+q
bH�eDP�;���gB�)�y���<n�J�I!��7��H�a���y��	�7�}P�y��xa��߹�y�n�,>����Z9i$�䑠&��yR�Ͳ1^�zg/5��� g^��y�j�:W6h��Č"y��)T�@��yҬ�-7>�=Cp��"o�b����y�nL�V>0�K"EP����n���y��W�s�}9'R�8��	�筋 �y+��MC�!�H6�L+ ��>�yb+ۺ:HF�s��'ʀ�iG�Q!�y���;@ Ա��/	�0]:���yB�ϻI���;G�N#{��mx��ݙǸ'i6=y���*��L��$b$��bg!Y�T��Ձ�/��;a�B�I�x��K����e��8�'�H�e�t��&��S֖t�:��5F��O��S6��|<���@�:e��"O� �Ig�6~| 0�5�E w�,���'�$q�6i���^pד=�(�I!�
&@��I2�G@![^���	�D$�'��o��CI0
ź|��߹l��	��Е*�>C�H!@��pFA�O�����N�a�8c����^�!8��
�L�Q>	А)�H:se�
U��BX6C䉂3�J i"Û'��Ԉ�+	=n$r):���f��s&�O�p!��3?���L�W/~��C% �:�?T���3{(@=r��u�����Áq�0��
�a7*�X��'���0I�_�6]aՏ�EH��hӓ:�����d�n5
2�9MH��`�$H�̑��̡vbt���TH|��E�ܐXop��&KY A�"L�<�"CI >"MC��׈D̢|VF�J.���c�#+$��s!FM�<i�ȕ	�襉���k��P�t�X�V\H���N�xLN�ɅG�#|�'c��6��v5�e�@��}B"�2�'yb�s�]��R���>~��+�'�1�ޔ��&E� ;X�����M&��癆�l]9lM�v�a|b��9 �2��f�\X�E߼�4�eK+l���ȓ	S⤳q�\�v�xi#Ve[%i�bFx"�C,����~��8ir�z��@T���z�"�p��x�t'ǈ7�!��_�S�\�qu���0Q�*;�T8��<��O�8Fy�w=.�:�&�#j�>U��$F�i/����'��b�n�1u^���dL�Z�h��K>�`D�?Z�	�=F�x���S�	� Ȑ�a�3Kz��JQ	F/ra|�E�
�z8�`}\I	RdH�Dߎ�aI*e[��*O|9�	(�lS�?#<y�e��;ڴ�K �͘���Zy�&��J��4mZh��=ٶ�iZ��i>�3��S i��IKb�R!��u�UPÀ]E�rǏ�>��h�����P��@����sϟ�~/�i����<3����� @ʟ杮(A@`r����0[0E�{M�����=т��Un���T42%�R�Th�T�D�H;Xe&�y�O
�	cm`�	UL��P(:pU*ʓ;'�0j�l�5� �IUL�`� �E~��A�%# �3iN�"�h�Y_�N7�FGĈ��GL�X�Э�"K�}�n�s@�(}�M�(V{��F#K{&X[ ͓�9��� �9����")����&I��h��-�}��)�ܴawHu;RIϼ_�t�Y0���;�& r�D���?���D(M�X])��g:Qr��+I�H��`�ŵrm�	L/��<9ׁ�Kyb�ǪU:�0��ڌN�r��G#T��?�ό�+Lt�E蕭S��#Q�	gb�3�D�^�8�{bZ����T�f���K����<�lo�`�Y���'"���t��J�'�&}9��*^�>{@Ǎ��V�ڴPx1I=Y�4Y�'f��1&�h�4G�0b�� ap�*o��!�IK܄�����9/[���C 3�.˓zg�m�w�@Lt����a~���S��O�ԩf ��.4x'B9.i*蓳4O���u�>IWI��E��U1���1OZ}��-���h3�߾d�.Q��ŷyYrњ5Ú�p���I����'��,Oh��$@��IV�9�K���2ɣ��9(�4(�bI9�O�	�6�L$%��!�E�M��&�����iX��B��<{ Mck��PF����X'G"�.ڭ$�����Px��&ʍd4���티Hx�t�JɅ"��H1OغNC �Ū���dv�t�>v��XX��R�Avx��#dM�a���`�Ŗ��?A�V�Z*�2f�׌>���-+Dm`��q8Ox���k+\ʓ
;�X�>�EJ\n���Ȑ�^��x��[�nt@����X�8��#���8�M4�hOL �d�}���+ը;��@t�P�DG��0<Av��x t�K�F�����*ʡ>�8���@��$�T�CWA4�a,��W�ì.���J���W
X��T" a�ო�q�����R��"U䒉��?���9Pl��J���q����IO,�k3�Y0U�bT��}DńX�.�G�	F&<�d��<��e((}K���L3ډ�q.�ڂX�'��.F�� �)�E�(|IĠ
��ڈ�u&�0RZ�YR�� KN��p��@3�	���-q�$��D�Nw�P0k�0|����'��[�i�A��A�`99�n�i5e�5�V�P1$˦��5��6���Y��	?Z,�q�Rh��Q'X��o�w��I>�g�7~�|�6��ܪ�G/Sx�t(��[��pP��՝*��1�o;����ɕ��Pܫ�ɉ�:�t;��˝h�^e���
)������_W��~r�Ѥ���5�z擄!&Z�a��U*F�I��V�U=Fb����lE�Q���j5�ņ)�s$.1�d�i�`��$%EI�%b �Q9��

��I�H�2
欀2� �Tl
���k�8��r�y yФIՆ`(P�B�Cl�~I��	 �)��ĥ6�L�:!��T����`�&L]h��ďc�a~r��XP�!�eַH �\)#��@��QU8r�fʓ0�Z�gy2�Z��$m� ��Gaתs'@����͂!�a2�	+	Z� c�A��U�$h )�h2%
S�2��xX��Q���$\�.H��Aɔ!�<� <��r �I�@KfO	�)>y�G�ɴCh�M(�HR�ēȦ����"(���1a[-~�AgҀY����O>�#4�ބ��O�ݱ��G�E�� 3���bU�,`��n����OzE�����L�f<�c�a�<�J�o�@e"�e�|V�¥/e�H+W�H1y[� �(�<���qym�<�R�O��P�0��䏴	�:�[�f�7q|��WC:�O�0���줐�7(˴n�����
I<�r��O<q�'��&��I�
dq前i�h�h@m�j�Z,��+	:N@ B��<t�ݠ0Z$(-<��QA�F��=A� � 2����'�����[5V�4���H�QeJ���'�$�(�);��C�ת'~b�Ia�Ёa	�����
J�8�3G�(��t�p%W�|l���$��L�N>QD�܏n�Z�i��BXlr�RY�<�ȰlTi�q�k������W�	7+,���?�}�5] q'���dj�:A�Ӆc�T�<Y�W�a����Q\��U��l�<�W.��0�J=�&�\�:�P`Ջ�k�<�H�^�<�ǁŊ�-�Wbh�<���5U�� �uhKp�1#�W`�<3� /DJ1AA�\p�i��`s�<�E@�
K3��Pd�׌!�4p��C�e�<Y��8:"&b� nd���}�<���=���v��h��!u�Pv�<� ��@��
v���o\Rb5�؄�px6h�%�q��xA�Ҧ�`Ȅȓ7r�G�0�����
��#*����� �AGA�	��x���N�15t���q� ��$Z�Y0����]�>f^1��f'��@�Z9q#�����I,d�Q���ݩ�&΂`~rY�&(^+"e��ȓ��R���@X)��_�
�Tąȓ
�j��u���o���Gn���ȓe�J��7'��B.)[J�������,���4OZ���L��MK��io�-I��&h��Y
� ߓ(�Ň�+0���� �(*3���&�f@�ȓ0ZP��?C%�m\ŪE��y���0�Ή�L�Y�ݼQzʉ�ȓd��C��T�XC=���� ��ȓt�����F����@U*6SF2l��(�܁P*Ey��-�vm^.�>P�����2�S�wQ�!A�fĪ?l�P��ip��ŭC(>1�3��$q�"��ʓ���aˎ(1�.��DD;o�C�I
R6A֍�L�Aņ*Y\C䉞A,t*��Z�pi�Uۀ��:JC䉇ɖ1(K�.]ҭ��Y�#98C䉇b<�Z�(����I&�X)�4C�ɔ&I��Ч� ��ig�9P"C�	�3��l9�웦!uv|����� C�	�������Y�d P��'��C�I�u�^��3gֺe<Pe���L�JB�I�K,������"�f�"�*�0B��18�ʑJvi��4a���MM'n�:C�<M(�Y��ĖU@�У�V�C�	�#PP�Jp��2�s ɐ%�B䉎P���@����Q`��鳁�@C��%�0��pf�o�|!�K%,�ZC�	;<t��;��R���9#"���B䉐=Šd	��
L-p}��'۟Z�^B�,!aFa�"YN����غ�C�I�]���x����%�����/T�B䉔5��]@��ʺs��0i�΂HC�ɞB��H�af$Ar�RTA��tC�)� 9�)E���BcR�NE�R"O��O:��	�኶�ȅ�"Od��҄ϟ%��Z����"O ���؞C�pM[��\1V� (�a"O�Mk��2{�ex4�E �Z):�"O MQ��@A����0$�x�^��"O:ma�T�E �"n_9>��Q�v"OܨJl �N���c�Ε��i��"Oz$Q�H��Vzb��g�/� A!�"O��إd�|h���!�~�zMS "OE�7AP<��1��%מƴ`�&"O��{E�]�M>��4G��ap���"OX�j���>]��)��e�	���C"O⥊�\�p6 �e�p	 1H2"O(%�GEL!7t�a�g�f(��!"O�$��n����c�"��G���r"O�\���B&�te��׵-VTi:t"OrR�Z�[�q�&F��u0�"O��h2N֬!�L���>��"O,HQ�IJ�7L�U��-���+�"ORѫPNB�x:d�c}W<�>M�ȓ�K�5e�\z1LB�|l����$=D��z��M DL<���Y�`�':D��ң����̥!sbC��b����$T��R���>	-B���[
z��b"Oƀ�Bb�K��`�΋nLp�&"OH)ceI̭2 ��Q�I�DA��"Oh�
TG�}й�P-�
g�P��"OX T����n=d�Sʴ�k`"O%�rN��T4��`:b��#�"O8a��H�	HB�5	�1κE��"O 	�*A�
4"
���*4���"O|��3���\N�㫍�i�t���"O��H4(�F �0�	.*��=�d"O��Y����\���M}�
�"Ov�1Tkܐ|�అ�D��`t"O�!�P�A�|�F�x��M,��DH�"O�x��֭֨Z��%"���"O�8E(&m�x�XV�AT:�j@"O�Y2k�8*����pS����"O�@	#��(7=%ɒ�O튖<�y�
�?�F�j�K�&?�z�g����yR�׫oK<�;3-۴"�!���G��y"�O�E~�u��c��d��@��y"�lW�誰�ƶ~��)� �)�yB6�><��!΢o����0���y��5%3�di��o�N�Rp�۠�y�g��F����a���:IR�Ka���y"o�(r��8ׄ��4
�M����yB�G�{\,R$���t�l�(��O�y"��l�^A����@v�	�oޝ�y�!I�웴`�������M��y2	�_���y��v'����yb� �&,Lɹ6d�6o~޹AV�E'�y��7��	���k�����/�y��0Bl�⣂6R��s�*��y2���u����w��5M֨q@`��y�C�+6���� ��<z�0[���"�y ��x1ܕ0��$����H8�y"��/�DEɁJ4;�!	����y"�ٙj��ۯVI�傓Cʑ�y"��	rdѲ7	ĺO�@� �5�y���>�t[P��5O��5�jQ��ybC,\��ЬK�{�(=2t�O	�y
� �q�uJO6B�6�B1�� ����u"On��[�u��h!�DĉWy:  "O�=��I�Dل �I�]܅��"OF�x�#S�9o��Q��QV"O�R֩V�C�LPh4��I �R"Ol\�&�_1��Af���l�.8"O�L;� hL���g"02� �"Ot�{f�L;zT�1q'�=F<���q�'ўh;������D�çB7'aPx@��;D�T��%D�Y�h�p���6bҰɖe$D�(x�W�:h���#b�f㚘K@@'D�x9c�P�j�N�I��R�v֮= �+*D�А&�O�{��$
��Q�.v�9�>\O�b�8���M�� �Ǭ͓!�ι�uC;D�(p����j؊f���m���	.D����ECe5� ��GW�W����f,D��d@I�9���wN2f|� f.�ON��@�S�OJ؅�3l�9�t�S��b��X�"O��jRm��H���h�jJ�i�΄�d"O�x s�F]�t�$�(�ы�"O�7O~Wʰ�0f�x�@S�!D�\�A'>8(�Ƭ� � 9���+D�kA�̫Q4H�1%-ѻN�V�f�%D�D�%U���O"B���P�M��<q���S02�ĕ��	5?Rz dC6p"�C䉋���i�6e��i)�d�6T�ԣL>���	�:��t�	�9l�4�jC/�&I�!����l�3J�]y���D��8=��O���9i�&�{���*O^Bh	��āVPa��O����ZPh �R�B�Qm�`�"O6�Z5Qc�x���D;,����'������.��r�֪I#>�1w�"D�p��,ކ1�#U�_a� %y��5��p<���K�n�6q&.��8La�Ok�� �'<�@A1 �%a/t9Q��Z��Ț�'���y�.�"N/�U" �ֶ_<��K�'c�X�gn�hj��GO\)L@�5�DK(<�'cיL�����	�\ f$I]�<1��N�zr�g�p�bIKc/�p�<9��K4��QV� a������d�<���ۖ�8Ls5I�9xMY�W_؟(�?�p�9�'W�n�&���	�����;
��z�̧G$$|9��ƽc�>����?��J9"�h:��$2�L�I�<�e-R���g)]� e����H�d<ړ��'5Jqem�~��X #�P`���'�����q��yy0�?Z�Πȋ�/����EH*�ny��.�'�����"O��ԏ�)c-hqJ�Ǜ7Uӵi��$IC�H�'�۬b��pJ�B-A��~r\����N�?,?j`���T�ZJȨ�%5D���&+C:P��,�,0�'�r�$��	��H��vQ�ge~x§C�r�J��,��X�P� D���!��B���g!��
��`��gآ.�L�p��Y��,�'Sa���	�.	�����@Q0�*(8ub�'W�!�D	�(�BTY��l�8Q "
~�*O`�S�OJ�7��uoXE���x��5C7`�!��%h� H����1'��I�BO	�d�qOn��J����Q��;���!s�o���'	�'�*%�H�n��Hi�|���"O���!RHey��|Ղ�1�"O�{�dӨ)�^`1E�ξ r�"O&�a��6:u�V��R����1"O� �rW�������=R���QD"OМ���S�Y�
q�oE�U�4�"��'�qO��I׈Z?r����Ʈ��1�rl�"OLB�
,7R��wn�~��)�A��1\Oj�[�@v���n��#YB}�d��?�p<9���\2oh�� 18fѓ��V.!��&��i�D�V�*<6%��Uazr�Ĕc��X��셄>$&����@!�Ċ�\F����$v����3;=!�dM�A8⨋V�O�f]&�����;;!�L�C����e��4l����ʁ�k0!�ܰ{��!�<%ZR��*^�|!��8w��%��^�o��HP�Z�!��L�R��5�1%Ƴ/D�۵��)8�!�@�`��+"'W�	f�K�\�!򄒉m&����ˠi�Ep`Huk!�G�x�B��#)ll�镖m_!��ǹU&\jP��<^�i(	�2I!�D[�a4Ł"E��O����ЧI!�D�w��!�C��/��0q7���p�!�DB(=a�к©V�l�^8	� �9�!�M��B )�X^�.�JBI�M�!��,��`� �
I���s3��$�!�X�	��[�5�9����6Z�!�˸!miv�#N|�ذl��!�J�w}�̢VΟ6��S�i[�s�!��ͷy�h��b�� 6N�a�!�Ēq���s��Z�Z���2T���6y!�؈/־١1!�c���2��<k!�״qth�G�P����#�U!�WGPH�p�IG�nP�%)�-<8!��?j�H��7c��Hx��_0J!!��l(����L�n�q5捄	%!��ۛb��8���O���`c�dH&$!�dJ�`K�����pd�6�L�!i!���	��-�1���/�BixT�B�Y!򄛠B�����2R2L鹗 &I!��� �Z%7&B� ��HP.\�~[!��{��*��Z:�a
U��/W`!�ł}?*ҕKӫ�@]b��G�R!��unQ27C$]�h@���_N!�^,jb�9vB�.����7E&�!�$?��hE�@"�8�r!��u|!�J18[�s�k^�/�1�EE5!�$ɿ|[b���h5)Lm���E��!�8H��,�� K/8Ԉ e�i�!�$@4"&d��H�;F�e��L!�DإG2Rm�e4L\�6�W N,!�$L:� D2���*��AĮt�!���!{V���� V`�*HU�!�$��B����g΃>�z���+L�!�^>h$�qjG�2��T��$|0!�dGZ�-�@����D�m&!�D)r@n��$��	bz b�+@!���g�ț �E�Cf�x���-!�Dî7�t`3�E7f4<�r��x�!�dX�9 �ۇm��bԨ�ej���'��\yA9��$C%�&�,��'M(Ly%�LL(P7��l��<K	�'��t�炅(�H��o	�qf����'7�H�@i�S�L����Y�����'D^Y�H�d-���dM��p�y�'���W�����:�n��Θb�'�L`q�E�}\��i�hց+�>%���� &��.Q�$��!�ٖBIbQa�"O�C-C�(�@�B n�t��$"ON�@��
ilP��
�G��#E"O�8��텪#�֐ Ԋ��_�&T�""O� ���S2JIZ�Oډo�qh�"O^X�d��.� ��ǢQ|B��"Ox�JeF�.5�%�0׸!��"Or��l]5+�\�GMк�ܜY�"OB�yD!��4���8p���0\��"O�Pk�&zk�ek���
r�P&"O� RG����0U�`��,}�"O쭹g�ŗG��-!F( �,:rp�"O��C���6���j!m��b��9r�"O6��e��PҶ��!�)(����"OP��S� {cL���D�N�z�+"O��b@�,)¦�C0Č.B ��%"Odдl %ĸu�ƍV��a�f"Oz�@A��c�(,�J-(�Ҩ!t!���þ��c����d���$5!�ؔ�e�"�� ~:ѷ��{H!��<u>y ���$>J|x��>h�����r�0���85:�eˉ��yb�
!_Z��A!�8�T�Ҫ�yn�)�tQA�Ą��	)�%�8�y獎z7��G�\E!BE('��y�1Pw�=ccᙜO�v��FZ��y�,�Jg����※D����`���y�i��du{THC�T��H���@�y��Y�E� ���!�F.�D���ͣ�y�!7ex�BՊg������(�yrJ��.����!&D��e�T6�y@��+�q�!b��[04�@G��yR���́t�ѡp�ؑ�����y��ϩFp��;��Y�g�j=�ы��y �+F�	�.
�*��(��yk�:e�\��֨C�U�Ĭ�G��y2/��y�����~�f���7�y���M��q����~�� DL��y��T��,�R��т#�n����M5�y���@KvL�SC;%n��%FD�yҬ�D6�����h,�@�)�y	Y,T.�X�r���HMJ��׃���y��xW�$�H�2?��`AGj�4�y��U$%y�X�T��7����y��^M��;��Λ ��z�˟�yҁ��p���5+��
ؚ�V��y"�oX.=s#U�zjH<z�,�y�@�.����V��"p���\��yB�D�b�R�C���gHhpBIֵ�y��O�B�^0cA���5{ �B�̓�yR��wmj�J�$#y��"���2�ybK�6h�25�B�=D�c����y��ي�� g)	�
"m"��*�yR�E�y�v���ězq�TIԋ�y"O�7�\�[�M�l���t��/�y�$�}�9
��H0\��K:�y��&`�� [D�'SCFyjdBP�y"�ޛ$�����=F�TQ��l̗�yBnH/p0�Q2�A�`xSL��yr�g�|A+� ѧ.�b	�R��,�yb�Q([�\��Q[�~BH�*���3�y�>V��<*�Ԟ!�4��fH��y�&ÿ+_H!�kT���z�
�y��	j��9'��GI��2Vi���y
� v��6��-����F�\^�2�"O\���^6�Z��N�u\��c"O����п ����b�^EV�as"O��[��S*x|��4fh&���"O� ��Ԯ0�LLZ �0Y�\��"O���E��0/�Q��	l�)��"O.�`!D�"�,��E� $Ol �p"OTȋ�cK7���s��JG��3"O����ǰ8�.=�P�Y�g��j"O�IzG�� b�I���F��WCN�<����	%�[$@kf���tU�<��`ƙ7�-2�Jh�t�A�VP�<�#�0#Fqi�^�W_�!�c�I�<����2�h�Å)jQ�LZ��Qa�<�1ƨ7�H�2�C?���9�]�<q"HM7
���%�U"x���r%hY�<i�'6�5�3�S���C���O�<����5���B���D(0h ��M�<I�돌X<5�`�K�`���ju'VH�<�% ,�8-�RcN?K�2�$��[�<y� )����k�&�2l�e�QV�<y�
Xjd,�B��(L��HA��y�<�����$�dlDI��(�w�<��a^�@Z�0i�mI�C�2�(��Ok�<!�"�;X�0�b)�*�
T��e�R�<� &��b�!v�����В�PO�<�%��.%JZ��U�Nd�v��o�<I�/ķZ� &�$7:�r6gVl�<х��,;�bI�>h�(X ��g�<�Ҡ d/4x�Q(��s"��ku��d�<Q#�$S�q�@��x��_�<Q���:Ю�P�ݾ$�~��TX�<���� �"��eF5`Z�\pb���<�B����fR�#\a.��G�s�<��ֆ[7�����1��`�ԩ�G�<� Y7;���c�F�du`��@�<a��!(��ǒ�G���j'��y�<�ů�f�b�"�
�����Ȓx�<Y�&k�Bl��$�4��z�<IaC[*t���O��r�X����r�<A@f�1S�T�bE�9^D����Z�<YEƳ`q�*��E>H��� �m�Z�<)V�Δ%-��Ӯ= BP�[��V�<qы���`dE:qhiRx�<A��#6X���&A�]�`���s�<��aM�B�C��K#/�2˰/Lz�<)�K%qJ��tCMI~<Q���v�<q�[��
Hie��1��-�gCs�<)k� �f��&n�xu�x�o�n�<�a�J&^�!��L�va�ը�KDm�<)`e�#�m��%�����[_�<�׎� ?�
}�V�F��|�X�e�Z�<�K��qЂI�A�H|���T�<	�K�J	I���>D��1���w�<���
]�ant"�t����l�<��ONΐ� `$ܒ��}Ag��B�<!�E]p�d{1`ߑ9&�f��V�<���:1�T#��^(��dg�O�<qGm׀�Vp���U�I��I;k�I�<IB�ɿ>��i�ǈ�>8$$��A�<�3�B��]E�����d�}�<YGLHq�:����1n��J��T�<��N�E���Sn9co� ���Ue�<Qcf�+r`2%��i�\H�%���I_�<� |@h���(=� ����9_�D|��"O�i�����\��q�DE%^��U!V"Op�	wG�a��r��	�m	H�"O�q*���U��,YL��e��20"O:�K��S�4��P�@ߞN��C�"O�=i񦗋�HX�&�(Xƒ�"O�UyE�F�V��tP�	4+X�"O�`sBj��{��(AéRJ��[�"O�$b��01���#_."�)""O�Pr��=x�m�.��,�hc�"O�x�c\�1�&=s�͋�o*m´"O>p��; �@b�N=@P���"O����G�����D@E%:?D��e"O��RO-��eΖ ,E�"OZU�w��t3j٨��[�xZe"C"Ox�H�b��^�"@#��G� �Qq"O�j���t ��\T��ƞi!�D�P����E�.U$�IA�E�(�!�$�2[	�dQ�']�~�9*�DU!z|!�$M�y���c� �QD�!�DC'%�HۤC�4�2�59!���xdɳK�%�Ħ��"H!�[	�*�Cb����3e�"-!��U-4�dE!5G�V�U�#_|!�d�M�\�x4�u0�`��G?�!�X�ll��iڮ8>�"�MHi!�-QcP�r�9-��CܜBF!��\m�n�����>Hp٤��j.!�d�Yx�d*�5y��C@��>^2!��B������{�(�[� �!��J>�����µP���#�'-�!�db�8A§��'�V=�b!����(	��/
 y��;bG�<)�!�D�n>�W@S���zGƋ\5!�ΉY�!!S�	�4�kC�P\�!�� �i�I����4�:�d20!�d@�K�h)����v�p�Sa�!��� �N,��UJ����0�T/{!���\ِ���Ѓmy�U��ȋT!�Y�PTjy����crv0C�AO��!�S�g;DY,h{	��X�L�!�VE���ũ�^V��O�:l�!�Ĝ� ��@Pg�=,(���ܱ�!�ğ�>����AA�=�򸣂��V�!�DT�rs�]:�ĥ)m�Igф`!�$��Z�Jd�ʖ
'SМ�d9!�d��F�� (f�#:4�
��G�!�dI#0�.�c2D�)|���X�-.�!�[><-�@�ƄM�&�$�O2Pi!�D�*4>�P�G�����Nݑ67!�$�Z}�#O�3����NջS2!��"@�p{�BD�ƈ��f^�`B!��|��̑"��+r�����5)!�D�*���b�B*��A���Tv!�D�4u��1�_0W#`����/=!�F�N�4v�Ի3N����g:!�7*��MsV��EԦ�Q�ή+!��L='���xw,Ue)� c
J)�!�$�f���h`C�Z��P���N|!�$Ie��LK�O���)Y�g�?s!�$C:~�����C�PC�m��́l!�D��$�Z��S��8��4�3"Ȓy�!򤇡QjHa�e�5gw�9ySg�-<!�ؤ�H�y(4Ô����F'!�� �]H�)8P�,D��JX%P����"O̻�遢+rJP������!iI�<�gd̈'� �3�(#4�̃�!Z�<�U���H�r|S�#����m#/�K�<AϠ�
H.V�j1l��W�Tp�<'�,�~��C��	ne�!B!mWo�<��/�$ti)R>w�Dq�!�k�<a4nR*��)q��o�١M�o�<	pL_>�(9Pv�O�(���E��b�<a�n�,t����^	0#���`��a�<��/ǔ$[�q�⤔�V;��Fc�<Y��Xl0|��S�@���[�<9gXH��<JǬO�L�n��
n�<�P� �?+~��3{9�9�*Ih�<���Kߪ�)���djP� �g�<��Q6+�����_�H�4�H1#@`�<�R	���p�ա�0!�<ᡷ�R�<ɣB� n��J��#�%�T�JH�<)�L�uZA�'�N�)�^5�w�^F�<���ʤ8S4��}���w�\�<���,�p�@NWf�+s$�c�<��Ɣ	�%Cv#�a��8!`M�b�<a��
��hٳ'��Ef��F��Y�<�coP�q��1�#cƻ#|(�FO�T�<Q��_��1�3�Tk\T3�JF�<ٴ��)�T���$��H��8���I�<Y���i�dQ2��*��9��(�B�<)'&B'<2�	p��x�`���F�<ᄇ��W&t����ֽ1\���w�y�<!뛷��U�/��QJ�`�o�j�<9�&�S��2S�ͯr��Bi�p�<����7~�ʘ
���'&/��#��i�<!��p�ؐ���9��%��Tp�<yrˇ{��<�d��GG��;�]i�<	�Ρ4����^��;%�h�<��FʍP�y��טl^��i���}�<I�MVrxA�g��f�h���{�<�v�ߊݪ�`�l؟j�����r�<��K0�x���^��u`��So�<�ƁP�^$Z곫�_.Ah��s�<	�D�>���*���8�a$�]r�<�g�M�DP�E�Ch��r�*x���W�<1�(�8:j��/� ��@�x�<d�МS���B/� }YhTA�t�<	p�[�D��sc��{���$B�r�<a�N�-(u�0�CMz�����Lr�<	�������M�N� 񚧊�j�<!$@�e���h���~�J�f�i�<yd_��3�AO�;�,d��dAc�<A*4�ܜ�'	sƌ@�V�]�<�Фŏ%�H�s�N�n4L��Aj@Y�<� Ĕ)�^,sbޛ$��I{@�T�<������3偑���  E�S�<Itl�@1�u"3��`��c�+�T�<���4�4m����h��)E�WL�<�u�
O���S�G!N]!�D�E�<�C�B��Uo�	5V��r�#�l�<ё�	����BB!@/�{g��l�<Y�F/H��� �Ȳv�����]�<t`)���e���1�
�\c�C��(���j2	M�E`�|%� 2hC�I�I�r�+G���L�|(�	#i�C��P��Dp ���V]P�cS+��C�Ip��p��,�pRJ�2��*Wf�B�)� ��Yu/��6��p�	��V{(���"O�A�ʥH$L{ ���A��ݚ�"O�=���H�M%�M�F͗�D��[�"O-b�ɚ�u�j�h�*S.���"Oh�@��8W�,8��26|0B�"OF 33N%^ij,x"�Įzږձ�"OT�*p�I�\J.]��M�^��(@"O�@�1��!=i�E��$ƅ��"Od� 7��Ed��$K��5�a"O���D߈�pR�ۑA��f"O$}���W^ht��
��"OF��G�w�f�q(T��\��t"O��kvM�>Xb��*���d��i�"O�19�oI�|��X:�`׽��e�R"OXI�qE[q�8s��Jg>@Ř�"O�Y㦂�D��(5�\h��U"O��{!�(r="���眎p���"O�a��
l�`�����!0��ջd"O��a�?M���唅&�j� �"O�-��)L�z���8�F�K�"OH��3�͌}n3$M�/�=Ѵ*O�A�P!�B�3L��s,��'hT�0�o�ΠXeb�oIJ�h�'��phr�$FG�i���_9�US�'B H��O�9�1�c(ɭL��!�
�'��]8Wj�)�v�
&�Iΐ��ʓJ`��ܵ3��U@G�؞&|:t�ȓ/�di;	R�H��ٛP�Q榜��P�����ŏ�^�⼻��Mw*=�ȓx ]�m��%��Ή>Y��dQ�x�3�ДRKB`�S��A��Y�ȓ8�2@Ŝ�kU�,����#.�"1��{�S�eC�b�p�j�j$?e�=�ȓjz�rEΏ����!t��a��-��!5��4h�9jY4Pu��5U(���i�8fe�Y�2L{CO$|�ȓ1�N���I6 kx=��jLY��r�Xp��Z�K�K��ЄȓBdI!�#B"7L�J���4��A+$��Q�$R��T�QF�m�ȓb��ȓ�V�$(^��ܐ#��؅ȓS�n娐�ֵe,�7�	K_��ȓ<6<���+��+>�}��ʃ,M ��	���Qi��|M�Lxp�⑆�o*��hj'*Dx��DW}6��ȓZF
I�Y�Y�p�3B��3,����H6PMC��$\�@��b��n��m�ȓ'���$���d���P��H1����ȓ�`�
��"Yꨘ�!P䭆�j��$s@���%�d-�AeUB-�ȓ( 
���o�
�����*2�b���b�����9tDT��$(��Y��mQ:y`E�&���"�*\�g��نȓ��Գ���go�u���7�vQ�ȓ\Pd��-����ڢ�4#Z�܆ȓs�>xuiTp�ar�X/j��H��p���V�4ɰ�y��-G�b��X��lk` Y0p�B܉�u�
��ȓ5�4�!4'P�SA^P���$���ȓW�4 �Ј�#=���7mȗB����ȓg�E*6M�����0�?9��-�X�ra��aBX���ғiE�|�ȓߺ�ӔG��t�0�r����1d�t�ȓ��ɋ!n�g���@D t�q��S�? �$k	���a�GǇ7A$ �`"O\�`���H��3p��3>@D}
�"O$`�p	מ}c��seQ�7:zM;�"O�Q���ȱK����[��r̒�"O�Z�o�, r�A��כF�`%"OdE��$Z���7�܉^vE0"O��kre�j�����)	�6�0"O�Y1�O?U�tɁ�[�ىu"O�����0=� Yd#�"G����"O��5�[�3Ux��+ܴ-z���u"O�B�DH,h)�ڂ�Ԇ!x.a��"O`Ь����+c̑�p�:��s�^@�<�.e�D��9W��Lq�ӫM��+vB��UJ�.&p�r��=EMV ���R�Ѥ�?B�mQ����1�Є�`EJ����2�Э8&ˎ��,���`�(XQA��~xht�A♈SR؇ȓ1T0�j��з�V�bk�ͨ�ȓ���	r�O'ht8K���CV�h����x�ըg�{�c� 9��$��n .|�%�S6$Ѳ%�ٽ�Y�ȓ@�LH��a�J��R��L�*8�ȓ6-�ؓC�"]�QJ����~���ȓS6��.l��%#214�z2��<��L�N
��9B�
IP�j�'�o�<	BƩiǄ}��� tv !JA�<I���D��;���h���sf�{�<�� ���<�4%@�	��{�b^�<i�FH\u���=lF�Q�T_�<��*P,#Q����:K��U;7��U�<�`�H��r4�2jZ��n�M�<���ºZy,i�<��Qa�j�TB�I!T�9#"X�O*Jc���/��B��53V�aR��D�V�x����لC�}�@�z����n#&DC��E�zC�5W� eY�g�fo"hB4a�a�xC�	]ɠL���D$��iЩ���B�IDΤ��B����#�R�SBB�	1q��CaA�`�S�1P��C�	�{�b�c��h�L�0�+�;��C�I�kG~����ضu��f��%P��B䉗� P���1xה�f�C�)/�B�I�x"xi��H")!`�蔫�0�~B�I�9�:p�ULQ!�2}R�o] UzB��bB�L��N� ��'��C䉭-�v��bD�(#��baF@u�C�	��^A�B!�$T���T��2jC�Iy1r�Z�.�8{אQ�U-B9;�\C�	t1Z`���.`8�|����|q�B�	j�D`�H'A�P��	��C�	�h�s��[%l�j��[�D��C�	=!����;�:(���M;�C䉧
h���х=$� �l�!M��B�	D:�Y!�U-j�蘻!��X\tB�I�J	"@q��G�`B�SN<IP�C䉣p��b��F2qI@-
S��r`�C�IX�蹆B�<P:̓vˈ4s�B� ���S�X k�LU� ~۬B�I�c���˴랷�JCDc��d �B�	�(�(�إG��*�07LE4<R�C�.&b*p���K��\y�ϩ ��C��36@J���6o&�dC���s��C�I�mSR����(P�up$�&�8C䉦)1C��Ȯ���ThЇ&c*C�)� �@K\w�d|�$�ϛ5��AG"O�)�e�&Fm��S2e!����7"ON�S�Q�LB>yAcE�7��5��"O��z�I� "$%�Ԃ�	��l{0"O0�RAeL*��hpWg"K����1"O������Je\�8gK+҈4�&"O�tu/�2<��p�ET����"Oƥ�l
[y*�f�ҍq� A�"O���4��1`����$�O(f����%"O��IuE�>�tH@�	6Xd��"O"�	҇B�A����6��T����"OdZ!�D&>�R���DT�=:  �"O�y�pΎ�o�I��">,$�"O;��/��8"�7Y#�T�C"O��pcj�������/�x��"O>%�IA��z]x �v�԰��"O��{�˖43�v$�M�t��QJ�"O�}hä%��㤌�7{� tZ""OBx�Ń�`�V-R����`D �"O��
AL^-v��� b��j�U��"Oh��)J�[�͢F14�6a"OBa��c�d�i�4�<w���"O�a� M
���x�eN�-Y���V"O��u�D�m��|CqoK9?F��s�"O��[@�V&�FҐ��S*�`F"O���lD/~�숫��%��\9E"O�-3j�	o��9�b��^�4�`e"Oj�x�)�,F����ر.��S&"O(��f
 �Qvb*Z���ˇ"O�A��U�Ht��4
7���"Ojq��� {�n�b��9��@2"OtEK�G^�)��RRENh��0ɷ"O��hߩ^~\0�>I��{�"O�⊌�&�zh���78��"O��j���X��p�$F����W"O��:�	�-�@8��ʳ2�l��F"O�P��J�*:YŤ FH(2"O��(�(M�!C$��":��
�"O���䪘�tن$+B�X�h4z���"Oؐ	#J��K6�� EQ,�"O�[�@I�)Y�L��
�?x�r�(q"O4��wʑa��� �	�,�~��@"O�����/�����[�B���"O����@	�6`�dK6��'�>L2q"O`���*%��thV'�?g'V�ya"O��֖
�~�(�fR�.�TZ"O�\k�#\ﾉ����>(p%�2"Ox��%Y�.b,2v��K�qK'"O�Q#�)X#�.)x�O�64���a"O��)4�S)%�-Sw�)�@�K��6D��薍��R���[6�M"}���M6D�����0;�;���*SL(�`�3D�8���:>�H=�$��)���m1D��#��)�
�J�Ĵ3���ٓ`/D���� �J���	�)� z+�`�m?D��P"�I"X�) da���pЪ�;D�D��$��	(J5�'_%f�G�<D���P��>���(�jA9w%���6D��#@#M;Rz�%"�@�E�%��c3D��P�+�)N2�U����G���Q(1D���`�Ʌ9B>`y�

/$>�V�3D�D3��$�s���~�0]Y�,0D�T�`/<��A��(�==��tH�(-D�����""�f�k!�K�1ɶ�℉*D�� �������j8�=�!	�(�y�"O^])ҥ�o���Q����ظ6"O�I@�";V�jq�\�u��Iq"O^�rGN�.\���y�(�-p*���"Ob1 "��4纥����4hx ���"Oh����ln� �4\���JV|�<i��4T$�4{� 岡$�v�<�B���)�J)J�mO98fX�i�c[^�<AB�B�F�4�7,����[�!�D�8
�FĢ��";s�<;B�5�!�$R>]�HcP(�VJ\�X2wm!��_id���gA@=�%bt��.im!��H5Tlz )dm]�~'` ����&bO!�M:��UP&
D�J�P�"�L�39!�d�7]��I7J���P�-#!�dG>K�����G�+U�b��!��3I� ٛ�EC�C�������B"O|�pC	O#��7�=@g��zc"O�����;K�`�nL��6��"O�5s�=W��M�#�����"On��%��h��шJ��D��"O�,S�J�%��Z�!H<�fX�e"O�C$��Ux, a�A�<O�XŒa"O`Lkրفj؄`xWFU�bt��"OZ��Ï�ZdPа-n�R�S"O�I��E (w��%k�1�z�P1"O�dB�⃿/Ĕ�U���1p"Ov=j�l�'���K�*G�rR�
%"Oj��N�iN��q���3"��a"Oz���ϱz�D ��G�0&[�H��"O8p �/L&�͈�kZ�VQ^Ls "O8�ҥ�0������W.�"O�H`�R�0!�Tɀ�<Pr��E"O���Cύ)���B��a�bX(s"O�ѳ��M�L5�����Zt%"ON|��"�;*��)#�׭k�\��"O���/��K�,�
fFV�q�"OH=*�"��'�`�9��arEc�"O ��TB ����В�M��r�"O�ْb����qJ��Pp��"Or��ҧK���@T���,�d���"O(�[`���]b���j���"O��2�6
E��x��\��P@"�"Op<;pJ�{-f9�a �\�FM��'W�`�ܩv�qX��A %
H9��'<c�J��TB��"���h;\P��'(�9�6M�Xu���A��`B֌!�'�����O�N�^9��b�&/�$��'ޚ]Y�Ơ&D	�gѣyK$�S�'A��ඏ��o���Ď ����'�p!�!���,ꖤH�H@:$!�'j�0`gA�3-fL��A��,U�� �'��Q�IF�r�z��sOV���	�'>��`̅�^)�e�h� "?�8�'�"��I���)������A�'�����G&t~T*A�P����8	�'�2y�al-?�h��[{�M��'C* 97���+O�9�A��;ʶ���'��c�ɛ�8��pa�%ۣ>E2�*�'����S������ ��>4���'ܠ�ir��%Yޝ�# �5��1K�'�^�*�5E�H�)t���1�l��'�f���@�/�� a�L^7��K�'��<"���_�:̑��-`:pA���� �$�BdU�v��4�%��Q��4�"Op�J+Ѯl>��`�?6��)�"O���D�t�n5Y�n�s�pa"O��� F�=�P��p�˴��K!"O� �s��V�}�/��p�`�P"O�}���T�9�N2S�NPr1�t"O�$���D15��t�� S��RD"O�)ȵ�v��h����`'"O��2Rǀ#���3w�ڛai�蛔"OJ����L�ԭ����5O]8�b1"Oܓ֠S�
�ڴ�L�ETFܡ4"O��8e
	pB.��Nf`Y�"O�E� H�8Q�p	P��D�-:�,I'"OT,��ÀI�0��fV�'24�""O�1{��V�A��h#�� �|ɲ"OF``H�w�DmX�$L9=��왡"O��zp��8�xI���V�4-��"O��#AM]A�	��!T�u��M!�"O,�Z��$�x<a�@�)�(}�r"Oj�D��VF@!�O�� p.��g"O����+M/R��$/�1m��s"O�Hcuh�iE����C҈IO���@"O��:U��vY�����+5�"O6P!�Uѣ�(1�ӷ"O�0y������b�R7b(
e"'"OTA:r
[�\0�ڠ%C=&�f�I�"O@�	�n˭䌱æ�I�}D�-1!"O��zu���O���zB�8	a���6"OR�"FA�Mt~�	��J�c��[�"O�SF�(w�$���o�,5��KT"Ob�[
/hA�(�t��J2��e"O�`�4�|��dni����"O�4z�A&@ $�un��5��q��"O�LB1�Ч^����mƻ��P	p"O*M	�/ñWS��ْL�3^b����"OXI�Ё���J����΀-E
��s"Oea��ܓ���b5y:���"O@I��^B��Q(G���:��B"OV��I�I�h� �/7��i{�"OZ𛰧 �C;NᠴOF�r�Τ+�"O@�s��OhLi����%�@"O����K�a�0e�,.�6���"O1J�֢g,u2D�(a�$�6"O�%�'Y=W�޵ss�Y=?�:���"OԹh�u��݉3ȁ�by4���"OʐA�y椲Eiα^`�x"O���fK��q���\�U��:�"OL=�eO8o)�	��	�qQ��"O��"�5~!�g
:���"O���`�C'k����2i�1 ,��"O���#� =�91�2J���6"OVl
�̚ ��=2M�4#�=Z5"ON����<Z#�e�f�Lώ�!�"O:����r��ˑ�V�t�p"O�[�-�?|�l�� �@"O5�W�z�L�DQ�X�h+�"O��ӷCC��b�;��Z5z?�@`"O��r�$ ���p"� �i	6"O�ԁF��1��!
"!4F,���"ObE��m�(X���"�)���D
/D��2��i}>���G�aq��9��+D�42��E.-����+>3�u��c+D�ڵ�%��8�nʾ!����5D�h(�oʒw���H�@�5H��p�4D�� vP��¥6qPĢA_D�q"OZ�ʤ�ϭ��P;$` �LʉH�"O>J�D�Pf����96:X ��"ON�H�j�	0(:�� �U*:Ɉ"O����$��a1
�����9vL�YW"O��3�N��Q���h�)��t"�"OH5P�Ȟ�-.^�k%H�0g/N���'V�qJe�d���F
��^
|{�'!t�@��W'$i�����b�v-��'!P�b�p��*P�\
`�4�'�DD��&[)I�ƽz ���$��'�����d����3J����'�h��&���z��y���́
<<��'x�XC�lE�>]��g���*��
�'����'�T�1!�����
�{�l1k
�'^|�`�ś>���	S��4��'bf(ɄN݅`�2����0�d��'�|�@A�`����@$���	�'�D���>A���VH�77�B��	�'�.�C�KǒZ�|�2�ݶF�� `	�'�F1���*���娛>��AC	�'_�h�R�!
��,q%aʞ����'�@�ȳ�ݵ]���eD���%��'�$�pAш~圠��R
k���'���tl�X0``�Er)��'�ڐ����$G�̼�a.I�X�l���'RZE�V��/p��a�Y�U��E�
�' �:�@�t�DP�A�A#N��k�'~V�(U"�E���JV�T[z0��'�tA�&㎼U�>\�t����\1�'p��ۡM�\��i�3��´S�'�(�f�Pfr���|�����'���01	�^m���Qƌ�r�=��'�dh�&���d�����6g�B�
�'r��DH�	�����Q9e��h��'vT���+K�5%��C�NSà���'���ڧ��pf�e)#L�JT����'A����/�)g�������!	��'󄼸sL�
�|����%}V���'�R���$�2 �q/�������'�����Z,�P��	�n�x�'�x ���� 	�F��!'֫v�b-��'*l��ß�������g ���'����rAƳ��|�E!_�h)C
�'r����O�!T8�0Z��Rh� `�'=��� cCe	�婕�� ����'�b�H5O�	7��@(Vg z?~t��'h5��EWl��u�4IO6�
)s�'���,�3[����kM9O��	�'��}�1��2괴4�I�X�}	�'�\�c�,U(4�-�W<r��ȓ`Nb���Vr��a����IW�E�ȓb`�Aӥ�'�zё���oI�M��:Z��q���|%f��`��y�ȓ��`����,r�"��bD�
�9��G�����`ߋW������vjU��R ���
(+")�0�׮V�2���Z�����_:�<=�e(D:����C�|ڤ^46�6�A�����ȓjYT�c��3�<{�J�i����AzjY�Cvc��7�ޑp�&���@4Hg�y
i(�őU ����#@vu��LۄS�4L���\^�<�ȓI�M���K  ��=Pѧ�g�f��S�? "�Bd�N%L��`d�։%ލ*E"OX����-�\���E����"O�-hg@E!rL����؀1"Ov\�cY�*6�L�&���6�p)�"O�9�0@!N���`F�Z�Pՙ"O����%l�q�e�߂k>�4��"O"m`Q�]�}O�jMV� 4n��U"O��q'�F-�����9R `� "O��2e��1a:H�b+^�N�ۃ"O�8ۦ�F[�QCS�.�4���"O8��@톹1-���u,��Q�D��&"OԐZ��V�H�PT�D̍��T#�"Ox �3/xL���X�1},�`�"O����� w�9S
̹?s���"On �&��6Mc	A3-q�9��"O�\є!Ƽ�I�$�R.U�!@�"O���g+�p����#앪�l(��"O8������AY�Ĳe�Kcm�q8�"O"��HQ��Y��1eYb�cq"O`)s��"\��9�C��YA��x�"OLy���B%��ŰA���@�"O�IË3i�����­e��S"Od ���.bN|������"O^�X$&٪eoμ`��֌^(.(a"O4h�
Γ'?l͊2Έ�p�8�p"O�����(xD�� ��(Ws��{!"O8%�	#{��R�-<<H�"O�b��<x��yp.�)}1�h�<YBA-2I�\�i�;K8p�
r�<��A#i�ҭ&셵`��Ă��Yk�<Q �/���e,\�HL$a���g�<����&d~$����f��v�L�<��#	L\ZTe��G�5:�j�@�<ivj��2R���d��Q��!�A�<�R#݀{���� ��n�`U�R��|�<ye�Q73t�+!��*Ȭ�"�m�<�7�V'��y�A�غ+2��X���r�<�ď�?C |���Ϯ#v���Gk�<�!��#@z0r��,b�|�+HYh�<��H�8#.�4�EKue&x{F��a�<YaO�P�Fܙ�HMZ�u���\�<��Μ}�h\�BA��y�����m�<�4e]Fh�k���Aŕr�<٧�O(ڜU�FN��s60X��x�<I
�(�X	�#��,pC2���r�<�Ђ�t9�Ŋ /k+��;D� Z�<)��R5P���Ӄi"B�<�R�`�<��$�7�T�#s }��V��`�<Ҏ-8V�`!�O�|:� nIe�<I�$��>@��D+�2�2Q�HM�<�P�3oj� ���
�T��!+�%�q�<��.B���B��ڈrJ�ۆfEp�<ѕ(R�-�8pҕa�()R[a.t�<��X�4Z�.D>�<LI2@�p�<�ͮ|]�%3V�4#?tAE��i�<��JiR9;aKȯP��	c�f�<QW��uF��K,<s`�r�/R_�<	G,�T�&��u��,g���B��F�<��D
�v��`�@Ϫ*@���#�KA�<�GBػeyp�!b�:���Rgw�<i`�!X���D 
-�'�u�<9��@�.�p����Ww�쨧��J�<)�� �Y�8`�WI���hZ�'�^�<)� �$<h�B���	'����%�XQ�<� ��:��J+l)����{z}��"O^���������6EG nl�v"O~�Cj��%k RCN.T�)�"O�`q����c�� "d�*]����"OĸX��Y8S��#���|��[F"O|��IB�AjH��iC=��Q"O��{��ŏU���jDh�V���'R�l�u�T�	SB��#C�5+�j=J�'?�x��)L��`z���%#\��'��)�f 8tX��lJ1���#�'ǞړB-2���Â�4���FU�<	��ĳ�h��&�2�1�JW�<�k�7}�<��g^W��`��V�<���{�3g�(E�U�Z謅ȓH4v�(g�Ş6�!��iI->U����\��Zd���"�C�d��U�� ��/�\�F!C��#d6-��}�5h�/E�0^����ǣFCj��?�n�`*X�G�T1�u��f0��� \>�X�D
��F �"d-p�~��ȓJ�|9ÅD�\�`cV�,��ȓV�q�\\.( 6A�BlLx��5WV@��]���I/c��m��vE\!Z�-d@Z��ro����E��\RV�x��xʉR�ѫp�X ��h3�(��؛a7nY� �%#?"%��p���T��9T���Q���
1�be�ȓn���*��
�Lu|�92"�)���OVҴ�&�
1[g��7+ӏr����;
n�� ��'O�	@v��\�~@��7���!N�1b��׍B�_/	��B`j5��mc|A8�a��'��ȓ)G.D���>c��3f�˯u��\��|��9:DO>��u�P�L��q�YqE�
g�"�&=+��ʓf�9�C��|�8q�QO�B������e�+�*|�Q�9U�B��- ތ�+�AK�G��`!�9dޮB�	n_6�J�	\�_�D;Dk̔)��B�I�+dP{1b˴DVlK3FK���B䉂0�������~�J�3�m�=-�<B䉧7���դ	�T���֨fV�B�I�R��+"¶~��JCH�3�B�I�l]�a��*����pㄎ�nB�YEΐ�Uf��dc�D��B�� !��7'�.�`DH�%�-LC䉋s2�eJ�E+>�
QX@?*�BC�	�k��m�HT�p�xx�]5E��B�I�\o굲�h��t��lS����|�B�	�^�";F"��Q|�RmU��B�Ɏ�d�+�%��T����eV�O�B�I�`����Tȷ	Ĭ����F�L��B�I�R1Ҝ9C� 6s. 8��_`��B�ɻ�B��IƂ+�!�H�)�B�I.���O��u��u�%�� ,+�B䉇O�@�C,� C��#��Y��B�39<̈{�ȑ�BW�CL4�C�|ƂL�W��Pʙ��h,Ny�C�	�YQ�\��Ψ$֬�����7a�C��-Z};�J��hj��FO@�	cLB��.mؐ8W�_XH�C� 8qB�I,0�.Xɲ&�fa�	҃(�-4�
B�dA���G�4��:`��B�I��� �wD^dR\m��A ��hB�)� D��$�24��0� Ƽ���Zs"O�r�Ğ$d��Ӏ.�x��"O�ґ��C�&��N�>�ε��"O�y� dֿu��)�SM<�,ӱ"O�]���
�w�����0Z�4d#�"O2�ci��]� $˝?�Z9)�"O�WR{�n)h3!I)t��Qt�^P�<顅F�K쌃�ѡF��3#�Xu�<��f7v��)L�m��q����s�<���	
���<;��ī�y�<����9X<��H/�򆔚���y�ȵ�X\�2OA]�6x`6�1�y"dN�lv@�� b�>~f�P�S0�y�ȟ �~�a�)�p���A7�S�yRJE���IT��_j�!t�Ϊ�yr-�j��CX P����y�Ѷ/��D{"��w�������y�EA=�Tsg�\��Ȇ��$�y2h�
Eâ$T���]�(c���y�)8�d,P���s���R���y2���dh����oԅ���9�y���pop(�U��%|,�J����yҀޑe�"��W*�`�*�jSgA�y��+�ꩋ��H�T`��KCdG��y�a�3`l4�B��c߄@B�oJ�y�(��Ʋ�;e��M�b�k�-���yBA�y�܌���"i2!�����y2��Ȉ�f^'lN4b���y��@�j��㛑ܒɑ��5�yriּ�8�i�,�M8����yA��9َXx��v��dS�.J�y���ov����ǒv��8��Q�y�ϕ!��A�M�A��=�� � �y�� ��x:��%2i�Yŏ��ybL�G�Flb4�C1{) �����y���7G���e��W�)���y�啎b`�DC _,�H�PL�(�y��Ȣ1�Qh&Q*��"�m&�yBm,.e25��NP-p�JI�,�*�y2�=K�Ii�F}%4��D�(�y���n2�e�wO]�K���x�N��y�E��D��$F.G8�QV��y��,k�2�l�rT	��H��y	H�,�z<*�h�	 a(H
�����y��ͯq0���.�(�gi�8�y2�&t�-yC`� 1��I�6�� �y��B?<�b!hʚw>d���̏�y�E���R���#u��!eT��y�l����@��5�\l��ל�yX! �dEۅ�ݜ1jx��ri�;�y��i��]�m�t�|����"�y�f����9�F�b4�l�4K�yR*��܄�2gk�ZG�x9Q��yJ̗U6ړi�8Oe*)� B(�yR�
|��X��^�L���䉚�y�՝-r�� VI�:F��m��M(�yR�4+jڱa�E�r�jaX&'�4�y�*��~~��d���Z���y���8F&�2v��pP@����y��9p,�,�O��k4�������y"/2:p���MS�~�zA�TD���y2�����`��{�H|3.��yr@F�%B���+�z(��b��8�yB��F��d���2]���g�!�y
� �$;-�1$��V� !d�jѢ"Ob��a�^�G���$��'Z�Z�J"O���Y1pPp���b�����I�"O�aV(K39�B�a�|�,M��"ON\iu*�		���N��P��&"O�a�s�Z��r�oP�~��C2"O0�q cU$Nd{��FP���"Onavj��H�b�9t�+vV��"O�x��K�h��,�2n�x��W"O �J1$_/pqB}��͕�� �"OS�f�0&��U�u������"O��2��8��Xr�L+m�"��"O��ru��gҴ�YîF�x� ���"O@5�N78���u��Es���"O��H��=�ze��Z�HS���A"OΈj'�]`5q�B�5@I����"O���Ck&1Ӗ��N��2�t��`"O����/�e,���,����ı"O�-#"�N�G>�剧%Lk�AS�"O )�����.�"GAn��z�"O�@�QAӅ&��b$�"8d�"`"Oح�4�\���!S󤌮��L��"O�e ��@;���Td��o^���"O�٢�"�8h\*<頍@�qt^0ҁ"Oظ#�A�a�W��O�Dr"O������*ʆ��b"��B@z""O��"b� ?�&�x�n�j�� 0"O���bO6��4H	�p�.A4"O��0��V��,���>
�V�J�"Oĕ����@#�s4B�"O�����-��2*��S��ͱ�"O�Xz�'	�0�9XUF�4\��(��"O����!�$6���B�g>�$�$"O� Z��U�K�l�@Z-����"O>�SNAT�ٺ@�8�f)2��d-��&�'�� KB#!<�H��5�I�'�
-�ȓ)��I��Ŗ�pYXT�Ӌ-6n���Z�l����	")<��C���@�U��SJ`0���*!��{��-%��ȓEբBڮ9�R�2�'�w?��ȓH `D�#
~XQz@G?r�y�ȓM�L�VN
 o�s�`ޕf4<���idm8��I	<�p�;o�TH��T~�;F&��*�L�4�̝!"O�0�Ӫ�	.����5s���0p"O�Y:B̈́�ڸ�2*�yO��)U"On�3�.]�Jz�Y6�}D�[�"Oa�g<D�f��G��44-J��>!�P��Pۃ��<�Bo�5&:̄�w���*��4�&�2S�В�r��'�����ݸW�"��ǥ�22+�,�I<���	g�N��r#��j���AX!��Q���x���-�Y�S�L�|2!�$�	z�~���$�o��r��&iџ�F�4�C���D;�Γ#���Z����y2��"q�|rcG�8tL$m�����y2�غev�SF �6e�V<h ���y���	[vP8��dDd(�z�o3�y"H	#1טQ�I�Q�<E81��yRJ��J��'E�^�੪a�+��'�ў����s6.ŌH7p���^;}y��˖"O��"�$�pKCj\,�A�"O,�!�*E~���ă�&Wq�{��	_�����"f�t��"bB
E$�-�#��1�!�� ��Cd�ۜx��T3��oY��"O�Ȳ�N�%j� hb� @Q�X�"O�2B�>d��{ũ�*P*|�s�x��O��b?���Z�[.�˦.�F[p���-D�@ړ��Z�
�X��Q�eAjM7D�,��e��I�,л�ۮs�����?D�4�Bf0p��I+��v@%�h=D�p�S!�a� Hh���.�D���OVC�I6�:�q��M.��[�_4��C�I�E������10"�S�M�$`R2C�I;3ޞձ�ƚ�'�N��C��X�C�	�
���W4��� ��@�+��C䉝2N!�2f�L=�x[7���'��=����Ǣ����5OA�g���N@�1�FΓ��?q�Z)5��3M/�� ��GR��p=��!ʣs�0�SnP��:)�ťBP��D�<1��&1����;�z��ʏN}��'"RDɧ����Dj�(C_0�����1�'�V� 3+��8��ɤU��|� O`���Ú�	�niZ�.։'2J�'"O��J7�<�㷬A�S1a�F�vH<9���R�R&�-?/�i����h�<�&��.O"y�D��:D% �n�<�4�B6���ѣ��ax�UصD@�<���"={`�3��3p]�գz�<9V* HxXq!
�$J�C~�<�GA)�@�#n�dVt�yB��w�<av�XH�"8��d��˖��s�<�F��=�^�a����z�� ��k����?��	=WU�G�#9L*5� *	^�<�O¼5^fH#wDϜQ�,���X�<�FޠK�t�r�WM-��xGB^�<�4O݄`�4���6��d�V�_�<���L�g����EkEw�\(h� R^�<�B"1'�f#7�E?�tX��W�<���'c)R�cV
��%���R�<�F�m���P�����c�J�J�<1�k�Js�4V�:��b XF�<��-�$(J��b���DǄ�� X�<��X*CC&d!����,�p'.	L�<���=`�.$I���E A,Q!,B䉙Y���΍.���	' "3� B�6s�V� $}�<@ ��RN��C�	�qࢠ�NɳD���:��ՃC�	6B�F�������!��Q4q��B䉛]�\AtdJ�Jl|��V�M�4��B�I86��fH�<F����&we
C�T�& �1�*d��	�f��nהC��1jl�ڥꂸX��}��
Ȗ4�C��&}��X����>�)s��l4pC�;� �3Dڥ8�([���>��B�I<4~�¥��5J$���$� bIfB�IY %QU�����@��S^pC�ɓ*�6��c遱 ��45k�B�	��� �h��j@�eDM�W�rB䉶3A�=�1īj6}ᦫ�J��B�I�aI�d��9��<!1NM���B�lh��`�i�7y�� �F��1v��C�	�,ﶽ�1d6"��cŎL�V�C�+"��XUdJ2��"�Ň5B��C�I�gN|�H�R�5`� �ƱT|C�X1�\0ԉ�}�&d�׫G0JC��|����}���Se��&�`B�Ɋa�����B�����V n1�B�)� i�b!��d�=PRl_&Z>�m�5"O.�#�hH)T[a���^/��pc"Oha���N-A������ʃ*�8W"O�hx%K�-��]v��p�;�'�2L0Ƒ��pY�KϸS��q	�'y��0F�'G�>��%�רJ�HH:�'��l����*�������A�f��'�ȱ �!�Y<��ԍG����s�'����U�N�C�~�i��{�F��
�'��)A�ܝ<ˬ��3�5=Z&X
�'BLeD�فmL&D[$C)n 3
�'@�Y'd�
�N�ْE7��#	�'P@ݰ�E�k�x�����9/�(��'k�Iw� i�,˴	�=�� �'ض$�6E��x��}+D�0x@��'��E�c V�Dd��H�+�p���'T,x�����<���X�����'���ڠ.��Ą[c���:�'f������J<��a�&.ܱ	�'[� �1o;M�L��O�!X�]�	�'|�u�u�L�~�,BP�E6(�r	c	�'��-	�@@�+�j���@M�ި��'��]�؀g�(Y�A�4C'd�z�'����ƂO�Ju�bI��$���'vMa�ZT^`ka����<��'�(P0s�ӧD�V���G�6"����'�f�� �I.
9p3��..%���'�|�Bf�O�'D8a�"��6/9�m;�';�A�n�^�J����Ҡ*����'�,��ǧF�b�<��-�7�1��'�4��4���8���A�.	��j�'oX�5�E/X�tD�GA�9{�Dq��'�P(�X:z���ZdD��Hv�D�'F�x���ùt�f���Y�<��'�b��u(Ȼ��@��^!&���'�&�2��.yĞ���g�4@��'�̙�T�Z-(Ƹb��M� y�'=��zBeͧ�V��4�̉4m
T��'E<͉������d�.m:�S
�'Ī�B���54tB<!ЕO���	�'A���NB0*:��v�RD?�E��'[
�kp$�%ܺ 9uJQ�Kl�T��'eX�K���|4�5�� ZV��5��'��0��K�<9�d(�4@��([�'�����O؀��i�4� I
�'h>�z6�&4
�`�~]✒	�'���q��f��:ӤRr�F��'u|)��F�6#���"�Ѩ7-��'��كr�Md� ����Bq����'���;��� �H�x���P¶h��'_b��f�0�	���5B�x%��'G@�`�P�b�c�ď)X�ȳ�'_��!����X8��b��_7�m0�'����>O�]�����ULh�'�uR@�:�bX��Fʸ��=��'N�@��B�g�la��ǻy�2�A�'[RI7I��zn=�aHY*x�S�y����	�+C�T7w�jd�Q��'�ݺ7�/ �a#� 9��+�'o|8;��X3���5� :"ΐ
�'I���(E ��I`u�n	��N�<�e&A��6DP��1�ܑ"�AK�<A
G1D�p�SVO��b]��Y3L�K�<� ���V������A7a�����#	{�<)&n�:�t���zA���0�_r�<� . ����|�³��+o<�8��"O�:��ܒr)��#Gg�j�Խ��"O0�K���
tSb�R�E����j�"OTyZl3v�J4r�����ʶ"Oh��5��BN4U:��W�NɖM�U"O�������(�S��Ϛm�Լ�&"O0p�_7��ق4��<H��Ya"Of��嬍�cLA��$T2c����"O�9P#�(lxQ#A� ���)G"O�� 
>kB)� �`dj�@"O�d@�@]X���6東xf��qS"OD�q��G/8_�A���N�`I��E"O�|�sm�J��"�䈃9
�{2"O�%��
>�䬋��Hw2�ɣ"O�9wCa����o�3,��<[�"O��K�#Z�딘R"Μ�q+��)u"O2�k�-��k�f�9wn�-<�(�A"O��Z/� ;BX0dKƇ�>�P�"O��I��6��cU��.�Н�"O���
-,y�C
�Xi�"O����H�>Lz�pd��,X�}� "O8n�f� ��D�̚%�%�"O��B�N�9'�
9���8s-���"O�Qc�/Z�:��OÜC�)0"O�D��t�29�s] �=c�"O`�d�ަ#P��2ՠY���G"Oz(d\h�t��89��I��"O��'�K&U��ТT�϶4���aR"O�y�L��8�l�g�&l��"O��r�A&5�T��A³4����P"O�\J�䀎m1�l� M�p���6"OX�Sl@�9�4���l���"OB�A�S���!�L�����H�"OF�PS���t��mӱ�R(N��!Ѱ"Ojp�ק�r.���H�=x�#""O�(�RF���1GK�%�t)��y"f�y[��:�b�6��@�$W;�yb�J�9Q<�q�e�yt��0�,S��y B3y�B-�`
 r'`}��E+�y��u�m �U�j�vҤ�ۍ�y�J>H:1�2ES;1�r��O��y�k�e:0XJ��ЧG��0�$S�y���?�.���ɩH�J������ye��!��1�!L�C	2Mi��ȝ�y�� (�B<[��żDO��:F�'�y�t=|�t=����K��y2��Gp�j�
�x��ȡ��(D���%bX&1���ː��l��b&D�| �(/sn��b�G�_�X��G"D�t�w��3,)^5�䄋a'�<�c�'��Q
b�p��[oTL��+2<���\�h�C��:Y��A`��Q�!��#Ag��l���'B��/Ww�e�V(�z<����7U��IYc�U2hJŲ!�'�S��y�/T��Q�b �Y�L|C�ɞs*4���48K"K	nk� �3�E�^3��Gz��!��\2$��2Z�dI�"%M��?���! ?�ݲ+�(h����J��g�a]<UӀ�\��K ī*u~4	��3�j�'�x����0 d�v���F�<�I��򍆃Q��i ���O<j�X���/�b,ݴ��ɜ+"~�K1N�'"�,4@۔	�!��2j �E�'t�l�3ǫö�	����)R�\A2I8�h�1L�3k��x��PE�x��1��WYB����7r���a9��q"�Y�����ha:�I*[c�(�j�a$�tI�V��ą╆�Z��0vB/�������<�e:��a�E a���1�"�� ,S��D��$0I��Xt��	N^H;���#5K�L�,L�@���p�D� 	�0Z�j��� � �B�C�6) ɔ'�DX( ,�
�ΌȤc�>��$N�ʪ��lJ1��� �!#�!�,NZ*�S����kV���S"OИ�ش_�̽Bd�[
V7�@2�cL�+B�Q�U-ܩA_�� �É$9ތȂ$�?%��*B21��w�z%13/�"5X*y;C�H�b�@	�Di�X�.O ����n#�8)��U�jE����M�%NL�"jA�Pj����A�3>�R�d�� ��O���h�3�t��J���J5°�>�gU�b
0�[��)� ��%<�=�U����Eh�h,���$N�4@7�,�'�!k����ڊJ�JX#D�)|OlM�D��X8m��iբ\q�Xr\��؂�K�H�ɪCe �g��Q���
)����JЭ9] 9v�Ou��rkC<2 61�+�8-�(i�'�|u��%�U�DY�5	��b1���6e�	X� u�ԔZ�ҐX��mQE� �@����E��g4,�,p�b`�=
h5s�(SLl�!�O�_�H�񤕹�X-��OX�2��/���q`K
s~����d�R������x!�.M�=FkT+����+�H�'�hL�bƗP6>�C��!J�J��I�t8��W�@����*"ld1�����8��K���bT�����U.8"PU�䥳T%Q��z�{�� q��X�j&�$�0�>�>Q:4�I&5�|%�'��h����E,��tk 7A�}�3��G�&*��s���'(+������	M��a4�Μ.�<)��;�>�U �Y#�9�P ��lR�^t1@)�0R�$����:�<˧F��\� O.E�Nb��|�GfN�]��l��!�a"����nm���{c��p�HN<H&����DWI�F���#��ԛTb�K|E��.Ա�HO�,q�"\�^��LC�BI�F��+��2U
�h�(z�J�`g��J�A��J;���3c��p��-:V�]�eⴱ�c��0?A���-t��BF�j�)�C�V�T�(����2��#�܀�*Pj�܁+Y�+J\&>]���$��eGƇ>�F���=D�`b#�ڧH���� �3s]x�FKϤ3��]�d,ٙId0�e�e��� ��(�#�M��|�@�G�i̖�K�+2�O&���}�X|Kr��&J�ᗯI}4��7�D�!n���1"���=Q��Ƃ"48�Mh٠RdR�'
���H?HD�C
�K�!��f<�i �K�{z��E�HY�ȓn���&�@%jN�~2���'M��j����jE�¬#!�>���	�3oL�(� �\�m��2D�d�RLۼ�1Y�+�3��0�.����XH5�I�2��`(?�3扐w�t���\�q��ay4�Y$}>�C�;q��)�Sk����g�ύ^	���.�@�0�����|wa|��O'��m;��O�0+T�` F,��<1�Ï61(R�p f�>ْ!F�Z5P.�0��I���L�<�+��r�L���9����3��q�^FHّs�8����$�M�|�S4��k� �g"O���o�}z�)�Q��6�pē�"O��+-wi�q�l�f����"O�Y`gG�f��,�P+�&3�N͋�"O���bȖOl	Ұ$њ��Q"O4��P _�B�J��h9~�"O����$� ���ǈ�C�<��"O\�A���!gA���1�	�"�p�+b"O�I�F�<Z�`i����4��D�"O�yz4Hג}G���D	�Q��[v"O2	�F��=_�((b��I ���"O�t���ަ3\��a	�Av�Y�"OJ%�Љ�
|�Re�ꄣ_8�=�E"O��zF��	.j��gH
?Y! 0�"O@L���K f�~ȁ�'��Xȣ"OڐxG	,�TL
��%��@Q"O|T�2���yd��2$Pظ�"O�M��Ηr=�#�k� /v8G"O��� B�N>0H�GY� ���3"O�`���jO.	�2���l�\ˣ"O��Q���&tpK�'�*ں�R�"O�ep3M=orvd�#��4�^���"O�$��Ɵalkgd�*/��u"O�9��AN8+u�L�$!܌��<P�"O�2u��5,g��⁖�y�L���"O�
ˋ�C��-i􎌲����F"O��JG�T�+<J�yuL��od\]�"O�u+�`v�t��
�3cVPӂ"Od����6���cd��6xlb]Re"O� N��O��m�'A�
J�"Ox��d	A� sxX�@� a;J�"O�L��K![<���ʅa�~�j"OfPz%�O��=�c��4g�V�"O�-��D�8JT�x)�K+B��U�Q"O����ʍ�e�B`s����;��`�"Ola(���
�^L  )��v���&"O6eږ���\iG#ƿ�`
�"O�y��B��j�r��%f�>Q0�"O:�C�F�l��8e��M�~XW"Ox�2�׃z��yk��$��*7"O�az�^�˒`1���$j��A�"O� �'Ǆ'����C�5#�N��4"OZ�th� �Dm���H3��17"Oʁ��┕|��\*�#�4'~(� "O4i�h�>	J!��Px*Xjq"OD�I$�Z�g�&4iD��J	ll�$"Omk�L��n�R`а��OJ<��"On${1�޵y�H��X�V��i1"O���a"��u�Ո� � �x�"O�S�O������n��#"O.h�����7XZՍ:�d��C"O�z��;
�@����$��|�"OH�+b� n{��+F���`M�5"O���0�ͤ.uxq�@"u����%"OЩBDЈ7�
� �J�#:&��ч"O@�X��4'G^yb7)��{�x�B"O
 ��͟&39�  �^�\l�AT"O �`�3w�t �qI	0
-�%��"O�z"h�?f�+�鎐@։�f"On �6#\�'G�q�6�47 t��"OR`s��$/� �% \��T���"Oh��0G,����x�dyx0"O���E�2(X��c�Dϵ5�V�:�"O�!�"ڰQ�dX���Zv11"O4�gܙ��	feѷ ��{�"Ox w�� ;a��#�E%�� �"O��a��TqR��C,���3�"O��A�I��l����ǩM�^ѹ�"ODih�B�lYD@�`�=	���:�"O��S�ݬ2s��k�����ɂ�"O,�(ǩf�vIkR%�>tq����"O�H����G1�D#�e�z��܀�"ON9��F��!�Q����w@���"O�Ń#�3y��	��Mr��q"O`���	A�L�`q��5Kn��"O<ؘ"-^�e�<�+����p��"O������-�(zu H's�V)I�"O�l:��\��1`R�+9瘔��"O�̚1!�4Df��*¦S I�,	9q"O� ǩ��Ct-3a�Y�_��=��"O��#�ڐ1:Q�%������9P"O����͗;��#�Ʉ�	�2�Xq"Od��R싚X�h%���j��iyp"O�@�� �j#�K�<wqF�i'"OVx��2vI�QA��)?@��*v"O�����+N�	��P�\�L�"O��DBܮf�8�� :�1
v"O���&T2'�V5j�� C�֡ �"O��H2�����ٓ����[d"O��:��ײ&�Y���I$�ƌ�"O�Hh�˙ ��0hpl�;di�ذ�"OJ���]�6�UaWhD9(Tx�K"O����\|01��ǡvv$D�c"O� ��c�ѕ#��xB���@� }�"O���@�<+@.��׀&r�l#�"O�P��dV�(� c��	�w����"O��QV��i�xx	2%� �^@jc"ORdX���& & �󆥐�z&��A"O���Eߺzb4���$H6,,�"O`�H�cEc��}�g��aٶ�s�"O�E�q����JزE. �b���KP"O�3g/\DPr�Ñ%%ǂ<�C"O�\c1#��� �hq����)j"O�����@�|����D+C�d�4��"OM3�"Z�{%�y���8��Q9B"O����I�7����[�q��4{ "Oh u�����o�@�V��6"O�:O޾{��?��	�"O杳 �ݾ@�M2�
L%��br"O�8����k��q��*��ʹ�H$"O��7�C:BM�t(BN~���;�"O�|�'&��.� �E]�<k�"OlUa׮M(P:�`���
1�� "O2�0V,�49��[t��,���"O ���"ܔ`��-U�ct�8p#"O&�J4��6��p�b�.i`Py��"O�@sE�13�(K4��Sj��0 "O.�
#.FA^ �Ӯ�/k��M�S"O01����ӌ��e�Ƀ.��H�a"OH��u
�`��PS󣟝y�$(*�"O��5�7��@x5�Z5�,k�"O,[�"ԓVz�L�1�ޙ��۱"O�h�d�Ϸj��QأƉ| ��"O��b�@-cp�\��gj�5ز��m�<y��W�����cL�r~��Q͑n�<����L-�8 Q�вt�B���'e�<$����3aE&7������h�<1aJ�@d�1���6�Z-�3��d�<�	�	,��C��hA�!���V]�<��.��
�r$��e��X�jZ�<�PN�i��ث��C [ q��AT�<�#̈C= � ��jMd�3��L�<�A᜿/\Db�φ�'�΍S�,TL�<qR�0D�H�"A�4���Q��M�<)�d� !����O/_5~5�4cXN�<)�T�7�`�B`�O�7o�S�NI�<��Hl��-�g1�`�+ţ�G�<�
�v���h�/&#p8b�}�<� @԰J�nQ�I׻OSn�[�h�l�<1q/G"U��� s��q�\�����o�<��i�� �Q�M�n����`�]�<�d� ��A	Q�\5��i�M�G�<a�+_�\Fxh����v��S���C�<�7�*�� ���C�I�t��m�U�<)�A��G*��Ճ��X
P�S�<!���8���m��}���g�<�J�^� �k�!�&}�����y��PAbh�[f��W��|Ӳ���y�.�9�~�j��T7�9���y�E�S̨D��i��^��,��)��y��H�~.u��5�Lt��)��y�C\$��L)�AB�{D���&Ȉ$�y� �'N�"�O�-ZK�y�&���y�	�%a��X�W�� \;�<��lZ��y���2��=k�B�,�L��Ø �y�l3[xl�t�QI����b(A���^�+U��}��H�Ŀf*݅�S�? ��ԌðoR,����5c��,��"On���Ɛ=�R�#����k�8���"O�q)rfEo��9҂{8���"OA�mD�I�0M�����p�V��""O8�궣�>)��ӶBK� u�ZU"Ou�u-E9jTP�Ŗp~$��"O84&A*
�5;�Ί N��!"OƠ��ό�W����6.�4vQ4%	�"O�-rd�,UlL�2j�B����s"O�t�Ё6w>|�Fǐ�z��r6"O�]�b�6��U��f0O��sB"Oޡ��B Gg�I��]-6�-)�"O0��UKl(���ڃF*��u"O"��Ǚ�I�� 2QI��B��"Ol$�2h
�p(��3���9"�6	R�"O�M3���80��(��� p�6��"O����h�,#��Ip�0<=�B�"OP)�dȁ=T�+��G�"f"O`aj��D�F�JE�Q�o`u�"O�4+�"^-������|貽ɕ"O���ؾ}h��%◧��Q2"O>��k�8sI�=fкE�Q1"OBܱ���v8!���P��S�"O@cD�B/�� �O �e��#"O�P0�Ƞ��W�H�l����yb��)cwz�2�K�'���y�m��y�^�\�GP:(�½B(�'�yҠ�9����O<F��x���y�ʀ�u�(�&f�u��M��y��_0,�X��F�; ���S��J��yB�4%z���@�5��谷�	�ybn��6��x`3H0>*J�b"���y��6b5n�r�iF��f-�R��y�eH4m�H�����
��J5���ybGټ:��+�.�0�ɚd)D�y�
D4Wz���D��*^F��"_��yBh�8;���&W�@)Bk �y2/�EK��h�f�=>�A!��^��yr)�9W�F��c�ɚAt�	.M�yr$Q����4̗�hu4�b�+�y�j��SPɜ�^.�ڂ�C2�yb�_�]Ŗlc���0]"�A�V��yr��i�R��cU�H]�6�y��ٟ7�B�	��.AѾm!T���yR�l$#�$D⸱�#�٠�y�F��b���C#� >�F9R���y�͜/I���C��d�ԚR�X�y
B�Z��	���tѐs�m��yB� z�,�B��ȟt٠�KP�Ɖ�y�8'��Ĩ���X� ���y鋖:�*�ɧ�__v ;����y��8=B,�'.	5I}><K��P�y2�._��\��/Z�y��m�����y"��6F�F9��'�~!ԸkR+�y�DC�Vy�`�@��D&N����՚�yb��6W@9kA��4)n`�G+��y��Z5�\ѓ�R��`F��y� ɽA��'��T|� ����y���*\A�X��]6C�*�IBH��y�m�D��a�Ћ NG�Qc��y�d�7m��"
�l� ��#��y��e�B���^�������y�dӧqm�`!I�{L��ɗ=�y� DSn�t�F���j<ި�4�\��y
�  ���@�,rh��gE�3��i"OX�aqC����4�dF�A`�l� "O�Pi�̕0MeNX�E�$,o�#"Ot�[�R�y��=[���2$�"O�.E��42��+#��'b�y�O��;�Q�&N]�ml(:6
��yx9��s@�"H��"�JI��y��M2|t�C�:r@6��C���yZ��кs��79�8�E�M�f�<��f8M3u��@�.��a���OerĆ�Il`���RV������  ��F WD��6fU�*�ۄ�,�@X��I
L�5�֪u����Ye^p	F�	�cE|�c	>���ȓs������{S�m�s�UK���ȓ[�ȻЫ
�$�S�
h|ġ�ȓT�,�k�fB�`*�A�uK�9"���ȓo
� �U�C?S�Dc�`��^�]�ȓFGT˄]0UWxyS�j��,��h��Xev�B����>!橡�C�,
(H�ȓ�|�0�h�f'�Yٳ$�Q`��ȓ`kv��s="XY�@��wa��i� y�C�¬Al�����-l����**��a��՗ 4������b�ȅ��6��R�U����,aUD؅�P�<z���p�H8��iC	<H��ȓne(`�QH!�C�.�O'$���_�H!6��,xv-;Qf٨Z�0��8�D��fm��
�HȂOEa<���Hx�i�L߅O��0B��D����v�Ƹh�@�H��B6c�/�ꑇȓH�T�BS
:��{3E´:���!����¬�B�d��b7d� ��a��[!�5XT)J��� �a��pʌz0H�&R��I#BR�vS���=8:�G(*ل�X���s�-�ȓv�Bm����&k�Z�sS�l�4̆�P4`�0�O��g�*p��j˓K<r���\��ո���M�\iq�)Ґ'�4=�ȓb�1�����HN�a����z���-�:�If�(GD6��#�Ǘ-�Ɖ��_Dp	P��FHQDq�P�AK��ȓO�"$#Ċ� n�>0�v�W)��̈́ȓ)�p��NC,^��r�ڮ����>P�1�N3K爙r�Â�j��@��P�ر&�Ɲ8�"�j"�I9A���!�}�6�&���¨-4O��ȓ
�4��M�Wlb՛4�X)����ȓ'���@Q�w���&�.{ʐ��ȓW����v 3s�8����Wŀ9�ȓt:Y�nJ�+�h pC+ŏZ@����]��q�%Z�� ; �Ƈ2Z���ȓZ�\�Ч��}��`@�D<%���ȓlq�p��M4(�#l�? �(��ȓ�\!�Sa��-���"��h��y���� %FR~�-*&#����2�b����֒�6��C0��:�@�U,��6Î(U.�3^�^`�ȓvjMYFAU�8������)RsN��ȓR}�4���֢u��t���2����ȓ	�� �������Ӡ,	��ȓ~���Ʋ�x[d�MIp �ȓ"���B�J
D<�4���J<la���ȓm�j��0@���=��:�,,��S�? b9���
 �,�RD��	V;�x�D[�Q4�! ��n�6�pp/�BK��;_A�yb���?p�y�T�SJ�p#
��V+��'��x3*�u>Q�R�Ӭ0��!Q���>���8��D$?
���8���j�n�$R��{Bᚗ%�T�K�Q�Lɂ�Ik_��'��|ʵڭg�2��d�F~�tcŌܟ�r�
S:Lw��	�V͊���#:�[�2I[1��1Z�6 �6�44��\0��4Ҟ�I4Y�������d��:�q����Ǖ�&�*ys�K�Q8h���JN� ^�bb�ҷ7����<�a��f�P��1����Y@L�`��(Git��]��?��D�&XN�z�'���n�~B��)�8(��I
2�f����K���|����ۗ�h��SX�P� �P/R떔�F�D6�"�@+q�)�ɔ"!�:�zFOƐ	:np(BJ�#�!v�<�2� V�R�4���Hc-�@�F?�)�S�OEp��I�?(d�Y� ϵ�$T3P$�a�	^y��d̀�	��S>иYX!c�V�PA�A�Ӯ6-Z���K��Z
#�>l�pB�U��O�O c�5+O|4��l){�\�A���2���$��ɝ���<H��� >P�:�$�0(2�1�_�>��Oj�뇋/�)�ɌN���baOS�z?^Ar���[�!�
	"��]Xfk"RG���'��D3!��V�9by�ĠԀ'Ț;E�(+!��G�>��	V��<���F]j!�Nq`������B 6�rP��!�D��r�1PS��`�8�k^)�Q��D���7��!s��/���a��y��1vL���	ݾ-��b ��y�V$G��h�7�'l��2��N��y�H�VӦx`�A���fM��y��$J�tQ!��8}�ʙ�P�y�吆���g{mi�h���yb��
ӆ�ۓH�m�"a��y��Z4(1
�Ңd΁Zx=ӡX�y�
 ?���+d�/UX�kq����y"i��mK���zX�x@ �0�yB��]�0A��Ν�8\+`,�!�yR�5Uգ��G�^����
�yBU�#�����ýS��U���y�&̄8ƀ����R�������yB.WY�\�IÃ��L�z��m�!�y��:}�����u�$��tc�2�y�h�c��!&%�b�*d�٭�y�c
�p��q ��";Z�WN���yR��� %X)"��Z�m��yb矺V�Z��*�w�P]se-���y�/R݂D2`J�%r��DhF��yr6R���wJH��ȵaeC�5�y��\9H�X�W���b���#;�C�ɳ.�
��V�`}���!ɗ�R |C�	?F:Q�!"�.N��x���P�1��C�ؖL�+�ђ0�ʐ�G���pV�C��5S�ܙ���@�V��P����!VB�I�z�܌Aʙ�!x�A/����B��N<H�/�+VƉA��[9�B��(v���Rm]&QX9!Cݩ�nB�	�N�+Q4b�`��Y�1JB�ɶ[��(�Q�(��S=�B��;l��E��m��5�Ő�V��C�	�qH�=�P��?T������B�ɸb��іD8p�����n)TC䉿g?�p��ݏ!�J����LC�I,��
5eX'wC8U���F�tB�	�GXX�fjJ�09�`@�$9� C�	-zP���B��d��7�JC�	�Y��f �;��\�PCC[�"C䉫٢���/��Xqs��Po
C�I�Q�n�룊�'bJ��b
�+h�B�)� �S��D�k�
��R�4:�ˡ"O���ÁW�b��]�B�F�-m�$��"O�G�GJU�l���u��5 2"O��J�l�!ix�8��	��p���"Or�8&#�"K֕(��4ʴ�z"O�Q���N�N�,%1"�I�8�DI	W"O��c̙�.[T�-�+)��,bw"O�ԑN˓M ����[�1����"Ot�te	�5J<Y���Ҳp/��w"O0�KlAʔ���]���"`"O��i���I����f�V/� �P0"Ov4H���3�^�:�	Z�t����"O(��[�6�:��gt98K"O�u�5���Y��3�ܝ)���"O�Њ��SG�εʦ/=;���.�yr���0L����*H9p�9��*�y�%7i>�ˣE���U8"��2�y�%,f6D$�qM�lB�2 ���y�X6[I�����I�\� �S��	!�yRːG�B����<	�2�Ӗ�T��y��M�DҲ���`ԓs��F��ybLܓxpp,j��Cr��K����y�TZ����*o�T�E��y�)�	��� a&� R�d
1�yR,��3(���ܻY��H����y
+/"�,����I��16ˊ��y"+� y��8�b`�2:�@1P&�y�oե]�D8�bܯ]D�Z��Ӟ�yr�ݩ-�^,I� �0(�qq����y.
ȥ�΀�z.�h2����yRh	��0��(�f�$L���Y'�y�l]��aI�%4M���$\'�yB9R��`[u�)&>�ZW�Õ�yR���H ��%g��N�����y�Э .h��#�4]m��c�ʊ�y�@I��NQzC�k��a@¯[�y����+�t�E&Z�] ���9�y" B�;�D7N�V�ve��M��yb1L&�+7GY�p�ະD�#�yҢ��jo�=�d��Ɉ�/Z��yrj��kX��'��E�D�����:�y��V��
���h�r�H�����y�d��$�z��U�iI�̢����yRiS>:�d0%#=pr%2F��+�yr�������6J�o���褢W��yR�Y�|�k�.7j@��r����y�bL� WT��-`��c���y@�oGʹ��aۅn|�ŉ ��y2�I�t=q��Z4c�<)K���$�y���mQD�#D�
+E�������yR��;H,)�Qe���Xa� ��y2'[�M�\�*�@/ٺ��0�N$�y���[������)C�t�c7�<�y"�	�n�l� �Ɛ8��:WOL&�y��ߠ�h0�c����e␘�y�
�fz�!���:���U�H3�y��b��A��Α}� Z�	Ɋ�y҂I:�J ��Z��iڃ��=�y���1< ,1�(�vP��Y*�1�y"O�+{�䝪��[ $��У�k>�ybG��3����F`��f���0nG��y2&�<~���᝽+�PŹ�k���yB���e��,"u�#'�Q�A��yDÈnH^�J&r�0�&N�y
� �����ݫ*��e��$<���"O4�pB!��pB�A��T�I���@�"O�YrţV`}*YHQ���|Aa�"O��Ұ Q�+����L��sN pw"OyqE�p�LQ�UK�,a^�zR"O�%���μ"���(��[>�2,xT"O�l)��ݤ\��i�&�+��,�"O�5�ՄW�^���q!��w�Q��"O~)8�nƦIA���Q���P�(�#W"O��B����D��Ż�.�*_�@��&"O�\�4T����m4Gx��"O��AF�E�pi�Ȁ��.�����"On��.�&NhAA�+Nc��Є"O@D��k*�(��K�7u��0(�"O,����,b�lE�a!�tkN��c"O���!	��i��0����|tV��q"O�u�&�$����a�=i:��a"O�٠T!��%�=P"ʂ->cʬ	�"O֍������2]�8Y�$�&!���UސňӫB&�\����Ȅf�!�D��F.�3�C��^��1س��-�!�DZ�7#�<3Ĥ72�KZ�b�(q�'G���D�$.����C�N�\�,��'*�BD��LE������2R��i
�'�\y�cÞ`[@��>�D�J
�'K\��e�U�A���uiF@�`	�'.����m!J�� �E�E2kw�Y		�'gx0�+	b8�d2�ł#2� E��'��Ж�ԫx�]P%��7.�2�@�',�d�^���Č^�?�}�c�ϝ�y2���) ��Q֥ >}�")��ycD��D�!!ПMW�iX3���y�:.f�`& ��b�4Dj	�'LN�{�oEM�dI�A%�jh�'��$9��҈xIb0���0 ����'+�t��#�,QT���c�� ~t�up�'5 �ڔ�I�.����� ~�<��'>��9�/=}�pY[U�Qt��p*�'?X��Ԛ5��`@!�=C0hH�'y���dA�7����t�P�®���'�����cJ���Ȓ���SXP��'Jt����"T�9��Α6�FP��')l۶8�<�g���6�y��'��xBB��2�{G���*R�'^̹sUMV&L�m���@wg�T��'�VL2���$T�qᨍnJ�2
�'�.H�l5�&|��_��	�'��܈`�F6S~M�4��>	#	�'��A\�Oo��{�JW#�h)��'t=¥�̔D� г�JZ:G5$]C�'2>XB��
g�Z��W�2�n���'<dha�(d)d�s4 �+b���'�����Iiʠ�4'g��C�	��4��F6�.�z���<MS�C䉋SMΜRg�1BG8�D��DؘC�ɸx��C�o�&~��Y���;Y�B�I�~.�1��>�4[�"�*B�vB� 8���JDAq  rȄպ��'����&;� �Kc�:X��
�'�>�`t�	�l2p��V� �}��B��).��rt&�� ���P$)�@CrB�I3j�8�:w�-8ӈ��'�Q�FB�I4D4�� �4���ثY&B�	^x���C�F�n���I��&��B�)� H�$P6`���pW�Bۆy�"O�k3�#x�.%Q�O��W/�3"O6Q�@�8�	ba�ؕ'PxѶ"Ot���&1-���K�,k��]Xu"Od�@$��B�6m⢢^9F�qP"O�`�BJ&g08�@�F�lm2�#"O���w�Ǚ[X�2�d�1��k�"O60���>�М���&t�B(�g"O����-w�dq�&AK�T6�0�"O��kE� �F��O/>Cn�"OBMҨ@�T�p��-͕AXh�"OP��&�<�Q�Ƭ9	�w"O�u�W�A�nbT�킋 �R<��"OF���kZ�ed��zS��~�8�"O(���C(W'z{'IO�c�u"OtV��!�vy���! I� ��"O��c��z����H�(/hXha"O�݀���pYJ�(oţ���u"OHDra���G��4��g��=�@"O*���X��!�K)P�����"O6�¦0@�e`�& �)����"O���?b�VV
!�lt.�B�<)�@$U�e�&�ۍS�s6�DX�<����O5�"�T��Lk@8T�(A���@L|���	��X�a�#D��I���a>:غ DF�Ok��y�� D�D�Gn�U0d�
�JB������:D� 3��G��UtBݦ/" �C :D���&�،i�, p�%%0H�ib�7D�Tc��>���ِI�Vb�]{0�'D��
�   ��     �    �  +  �4  D?  �I  �S  D]  �h  �p  �v  {}  ك  �  ^�  ��  �  '�  j�  ��  �  2�  s�  ��  ��  J�  ��  �  ��  d�  ��  � � � { �%  , �1  Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�� |d��"O
`�(�;���8���-0��1%"Oj4��ND^[��"3/9�0|H�"OB���H��*�ʞRy=a"O�味V�!X��!&F�:J�$���"O,��a
���C�Ą�M�"O,$3%o�-���p���+Ն�:1"O��ݢ1����`���y14]2��i�<�6��{_���c�H�`�fX�$Kn�<��A̼VI�xR[�)�Ć�pඤ�ȓA5��('nߡ4�� �)˩%� ���,��r�؊b#`T�eT09���ȓ!�b��g��}�8�F��-? �ȓ
K|m�ș�VṔ���2�%�ȓ"R�X�j�4JN�1�˘X�i����̹	_�jZ��1!g��zܶ��ȓgil,*�J�
j�Ne��i�J%b���f	�(U��:���G��$Y^م�~r�� S�%T"���k\�jx�ȓ|4�1�îJb��@ӵ�ݩn�V��/[`�"�v4�R�!ʎ<��M�ȓ`:��z�ؚh�J�Z��$HY:	��H��p�m�C1��!��B:��0��EnjZA V;9����J[
2���	��4'J�EA�IVW&��~�(aZ��ӹ�>� o�Y�|�ȓ�f�A�
Ο7�H��M�$�����mޠP����/���ANXo*�ȓTv�����{ ��-7�*h��I��sB�8�8���3����ȓNe*M�悡;������X�o��!�ȓ'lj�#F�m�+R&;�|��2)n�C��0S4���T:
b���:�0!��e֊��)��ͷV��,�ȓ0�&�8#���� ع�L�����;�P�AFd���,w�6d��r�EQ�( �gVlɦ�M,H��,DP���|�I	$G#\���ȓ"�)���E�B	yt&B�^�LɅ�4�� ��eëF�ڙ��n��R�p��hO?� $�=t_����OĽU���Sѩ'D��
���B���9�߫�.�(�8?q
�iy�D�A�הS���g
�>���ɐ���ڮ!�P�*��1���2�h�)_eB�	(PԤ<覍B�%Q��A�K(܁t�I3P��>��
<?TR���Gш?A�A�����!�d��a���jK�Q6�Z��\%y���+Xaў"|��L���;�(��O���
�kXX�<�)�� ����@OP#v��Q�ڦ����%���M�rUST`�*qPz؆ȓac��e�Kx�2|�(��+��t���9��JI�k�&S�g��(��ȓ��#�
A�H�r`z�ǟg�Շȓ�@0���s��a�!İe�`p�ȓ9E́�+��0ha�h���d��GhŘ�k��\��IB�?󮐄ȓ(���mW�&ލaJr"Rq$�0G{�'�D�)p������BEѮW6���e�VA�<�V����̊�/ժ	�����d��0=i��C�Z�l�	3DU�N���K6�Z]�<��G��6�"yQ�ǨZ����c�^�<���R��\��(�+n��i�U*�W�<� �-��(K_�\�	�ꚶ����"O��ٲ"�:M �ൈޙd�� v"O$���d\�%��p�4�N�(YS�"O�D�W`	�d �����u?2"O�TPpE">`$��d㇯+7N����'�x��a�.� �	#H�d`�hY4ڀ�ȓq�Ic*ܡ��q�N�qz��E|��s�O�J��$N+#
XZ% J�z���'>Lm(Tj�W_�2�҇I�y�㓑�B!�Flڰ$kv��0�Їȓ�HDg��0�j�C g�܌��K��hW�-���&tȓ K����ΉZ��(ϖ�a���ȓ9�l�hC�ߘ7|�A��1����lE�ƌ>H����cd�4��ȓ6,f�Z�� Xrp����^�@І�W�n}�d�̬q�h��d�A���so4D�ܠ�O�H��}�F��~���4d/�����Z�'�H%Q4� �`qL0j7�Յj�n�`�'-������	)	���&cάn�B�ʓ+����/� J��h��M�1
�v���\���D�"�p����fL"�"O���vF��(��9��S0�\m�c"O�ӫC��mj!m�?9z51�"O^�j�͂�9l��匝�N"�m�D"OH���8_�=���{fp"O̴0�eC��2qI�;y��x�:O�=E����pZ��0p�fI��y"��o[�M�ÀK���Q0�����~rl�o���I�!���6��P6�n)�1�$D����N\#fB-h��Z�-r���$D���̙�
����pB
2vXR��"D��� �� ԉR��I+,��a!D�h��f�*G������Q����fi$D�\��+�����,�����g'&D����@ռ@p�\q��'u��gO?D��SCH��?�6�!�$ �b㐕��� �-�OH�Q�D�J�``aPNW�&�V�r�"O�#�������mL&�����"OX ��
v��m!,Z�c���ڃ"OX��� �Q9��$	S2D�2p�"O�hH��9*����t_�.Ԑ�P��E{���4i�X�����(��^�@�!�$ҐBfd���}K�f� ?y�!�DR*�,�;��ԍ0����ղ
L!�Ϭ!��b-6f�anŅ3Dax��I�YfQ������֣�.KpB䉤'4�驷��b<D�Q����JB�I� k��6���X��2g� 9LR���0��jUj�{Sh6z^�X`��_ ఆ�:?����W'O��I�p("�Gy��|Z!��#>��q�	Hn
��q�ń|�<�ҡY�� ����=Ά�*��,�ў"~�I�5z1��E�\��uP�/��C�(B�b��v������-�pB�	�:_2��HV6�|��u����C���4r�E��g�R��cV�-w�B�	�r����a�@�	�P��Fc�t"<����?-�s
��>T�j
 i��D�`�2D�t��eSFL���]Nr֨/ғ7�axB!�
-�^��q��%R�(�0�Ԉ�y2Ɯ_�.�1eǯEO,Rs����y�R�s��Cr�-8��X5�7�O�=�Ou.dR��>����RH�"v���	��� ^*��=p@*�Q��:��,Kr3O�=E�4	�ds��(!�Vp�\��SET��y�%_;P��y@�.m
����ȍ����ßt���/�"41�,Tj��bؚ�dB��֟��Ύ}RV�1���.���Jw9D�tᑭ��ur �+=�8��'4�g(�E����X�F���Jؒ
�L<yQ����y�F�z&ltY�l\W���iƀ�yR�)�'3b��;��O
(^�"ulW }_�-����t�� ,>�&-:s!� Ԍ�'��}��CO[�V�o�*a����~�B�>S�i�%���-t���F(�B(�B�%=��PA2BS�]�v�hҭU��B� UՐ�*�Q�q<�E�'��%�FC�I�Q�����X�.cuRN�9�DC�I�d����Ё"pV�8�B�	&`t����<i��.C��}���WQ�>q�%._�<���!:e�2-Io/�i����o�'��?A 7��=Q�$��!Z<j1:D�R��
2�6Q�6i�^U:Y���7D�;�P�[_�	1�Ͷ*R"�%�6D��e��QҒ���(G��sA5��)�OD�d�n&Ha��� n��W"O�,�Q��3�(����ݐ$�v�P.�Pxr��6V>,������ �p���M�>�y�B:��8a�{��{�@V��y�
G�_��!�E^�.B:VHO�y2ePKO �Ц�"$&��YL�&�y�FK�Mw��ࣩ�"܂�{�KW�y2ݍj�p�a��&��}�@f�3�ybk��P&SVmǹj�������y"&�V�z���e�">c�x�%i�y򫅒K�����Cf[��f�>�y"H\�>Z>�رAE�d	 ��`H_��y�Y��}R�ʓ�o4��r����y�)K2=�K���S@���hY��y�%�r8P�qC�D_�y(u/Z'�yr��.p�@�B�2L�|-�͐8�y�J�5H��Yp
6F� U���y2k2�|(���!V�>I 1��(�yB�P�ȁ \>]Ռ͂3�Y�y� �k9��"�£'��c�G��y��L��^Ż�c�V.m����!�y�E��'ZT���&U�=����p����y�F?1cp�R3j<䉰��ǿ�yb��[��:Ĥ/R�����ۓ�y�B�Td�Pg�޳J��3fۢ�yrEBt��B5@ָD���م�Z%�yʒ-@�8!z 
 <;�,�{e���y��J�~�R�Qv�X5;�X�UgU��y҇׳]��*��
�?{> Rv��y��^�͑�G�9Fa`H`�,Q��yR�Z	�A�T��4Eڼ�zq�۠�y�MR�6t��!O�5��%B���y�ƓW�A2�b��CA�H��D�yr�JFJ��	J�
$� �6�Ҧ�y��ʼvJ)��3ϐ���	*�yB�� �&(a�͘�+5��0�@B/�y�o��_����ņ�6����$�y�ǖ�h�F���6-���1�&S4�yb�]�bҶ��孏�W��pI7l�>�y���7 �`z l]�<)P�ge��y��2lr���t�29�]���X�y��&`�=c��%���A&�L4�y
� ��["@M�d����f5p�"OJ�S�.�%�R	�g�$�ip"O�,�Ο3n)����/�Rw�T�W"O,}�Q'L"o8�� ED�46�zQ"O����Y�}���i�BR%p�MKe�'GB�'��'iB�'��'~��'V�Y'@�:%�3x��IT�'b��'=B�' b�'��'B�'aDdZe
�@R�7��b��`��'��'8��'B�'Zb�'���'��<cQ'H��¢��NOZ4Be�'���'I��'b��'�b�'-�'��M�F�Ň^��[',�#~.����'I2�'���'=��'x2�' ��'n
�	�р�H 'L�'u��X��'���'���'�'�"�'���'�`I3c��0�FX����U<y��'�"�'E2�'���'���'B�'� bcD�9>��W�Ԙ1 0س`�'Y�'�R�'���'
2�'
��'Wn� �vxl�'��}��aK"�����������I����	͟����H�	���P�Վf(�0ᒄǎQƨj�����Iԟ����$�Iȟh�I˟��	��������2G6tMzd`A��4�������埸�	�$����d����҂�J��X�I2ʂ��B�B��X�x��ݟ�I�h�����	⟘���@�W��1gl��
A+�x]�G$�����IџX������I�����M����?ѣ$�$grd�&�Ǭ�P`�(@K�����������Ϧ�!���=�|�bM��0�
\�7.RR���-�f�'Hɧ��'�J7MF�fd\�q�D=#�ȁ�$C(��1m�Ο��w����'����s�L!���%���[UH���CH���D���d�O�ʓ�h���EU�z��#�A؁���H@̘�i* �/�It�'On��w
��!�F��hJצC�L0�,l�d�l��<��O1�&iCf�r��I�+o�}3@j\�_B<-��B6��I=�e���\�:�*`G{�O(2�T�%����� �dJ8`P���y"[�,%��R�4�<�<�B��\���Ō��@�Rp �@���'�<�<��F�y�(�	G}�n$�zU e�҈2�̨H3����ߥAj�ܩ���>B1� ��B�u�	A���4D^��!q̃�C����)O.��?E��'�$$�1�Bxb�d]o�Nh)�'56�X�KJ�	�M���O*~�p�cF")B�ҡ��f�F	I�'�d6-Ȧ!�	����mZk~"��1a�V!��"�G[Fْ���Ȱ�2M�7o`�]�â�0C��}��MA0��)S�g�38�]'>�%jC'�.W�B��l;4�?j_´��I��!򤂟z����ӿ
�<�Q3��8�qaG+x�30J�?���Z���#W6�ll��k�H0����'�$��n]21�x������ ���N�2��r@�<6󖑊�� ���DHkV$�(8�r���PZ`ɟ�m؂�klD�N�k�֘0��k
�'��,��A9c����'�"�'/��2?)�o�R��l���ޛ.Z��B�l���	ޟ���Qyʟ��I(}"�8\^���,�:{����d- �M�g�(G{���'�2�'�d/�4���!PAV;2����OE�[�B�tBK�9�%��]y�'[�Ϙ'¯]pae8�
�rD�׮�%/�27��O����OL���f�i>����ti��L���LkL�`�������D�Oh��%O�1O����O���A�r�1��Y�d�a��!V!DamZ�p������|���?).Opɹ��Bo�a+�
��Us<t�U�̦e�Ip7`c�L��ğ8��GyB/~v� 9t�24� h e��f�����-��O����O�˓�?�e҅aקMj�p8��3"�|IC�`SK̓�?��?�.O�m�� �|��K��-= f����hY���@}��'Z��'6��ßl��,�\��0D �.B�<�6dҵ��TȢl�'Y2�'�U��z��<�ħ`��g�?i,��V�I�&�%@v�i�B�'��I�\���	�c>U�#΃>n�������7�ڠ:0ǎ��MC��?i(O�-YA�w�T�'���O긹���ԅ"
���#^w�u`p�>Y���?��p"`1̓�?���D��#�O���P�ڱo�������>m���3۴�?1�h
�$���i�r�'���O���'�2(�AF�1�$�	-Qg����O�>��	��L2��?)+O��,�D��[�*��W��(�OR��M@(��t1�V�'BR�'.��O�B�'����m�@��D���X�d�"S�6-��}�j�$�<Q7�Y�|�M~b�'T�6�cB���}l8aņQ	(��d�is2�'���E�j�6M�O
���O��D�O��I�C�d�CCMVUh����A�S��O��p��d�OL��O�b��8G�t����k�� �ݦ���(	�Q��4�?����?��b���q?5bG(Yh�ݢ4��(Y�k�n}�g����'��'��X���F-�6h �O��f�x����B}�qs�Ojʓ�?y.Oh�$�O|��5{�����X b;spK%��ASp9O���Ov���O����O�ę�q�Lo�?t}�-#ӍĴML�=iu ��P�ݴ�?���?����?.O^��K(<]�i:�P09��]�D&�գ2lфrw�<o�ʟP����t�Iן����@ Rt��4�?��L�[4�L�Dh � ��	���[�i���'"�^����"^Vt��=Ӏ��]l�*����}�YJ ������Iȟ�������L ��M���?����"&Z:o�r8i1�W4Z��iy���?]��^�M�.O\��Vl����s�� ������'q�ĥ�$'�7KW����i�2�'� �օj�F���O��$��J�I�O �q���.2H[��8���A|}��'1f���'��U��B�i�Q]���MŃ U�9gI����PB�7-�O��D�O��It�	̟��R�N�d�h`�E�:!g"�9�	��M�����������Q�ZO������B�x�&ǽ#�To��\������%���?!��~r�ͽ6X������
`y��`��'�()p�Bg�П��I��k�H�)jn��4�Y��v/Iw����'��,2D#�$�O���(��ưUqQ	w��	  �J~$�X���!���D�'+2�'�Y��钪�$/��P��(�@B��9��}��'z�''��'q>|��eB<��D)D�!˨�p�H:W^b\�8���l��qyr�C�0b���!ZDl���5��# I�5B����?����䓪?��L�!b��#6>%�!T���Y��9QL�C�T��������Iry2J�7�v�p5͍�͘�K���9X�JM�C̦=�	w�IƟ8���~� ��h���&T�dXv���F;WU����i���'��(�(�L|j����ui�H_�z��R}� �#E԰<��'���'����'�ɧ�)�3(͢�����"�(���G��U�,�7�@4�M{�Y?q���?���O�1Pu�OΞPR�[� ���E�i���'����'�ɧ�O���Z6�ޖS2`ٛP�۶&l��4-��{D�i���'�b�OwNO����2MJ���v��4Q?"�;�-��2��n�Oͮ�	e�)�'�?i��ğ�К!b� �%�M� ]8�K�4�?���?)ѩ�j�'B�'�Di�H�� ��kĎ`"Qk�YX��|R������d�O�d�3B��鉗$��{��q�,��lZ�4���U����?a�������!6}�eo]�Dd�&�Xb}b��.i�rR����ϟD��Iy�A˗ڢ}Y� �J�(c��� B:��O��D&���O���J$I\�[�EI@���/F�q�u����O���?���?i*Oz����|�xڰdb� �@[�����z}��'g2�|��'f��G/�b�R,�zs�Χmg�����$c/���?����?q)O6<�A�QP�Sz�<cԦмw~q{��C�����4�?O>���?��Td�[BRtA�v� x0$[�4�@�[�C�	�
����3���\�C���
�0���)*m�q��1�e䁓%ۈ�{3K�>[���y�H@�2�y �
O|]���V�f��9���[R���ה~�`�#�e�V	05A�DtR=	W�U>h�(=17�I'I���Ҟj�&+RcQ���$�Q�J�x�^{班A�����@�'�~t�tjH4d֨j�e�7�Z�ӭ�T��;�e��h��(W"ɨ
����!f.R������JWb\�ѥ"����5A�-Z#�OB��Oj�d�кS���144bI� L�Yn��R��D	r,�ꀥ�<``���0gl�X����xR ݴCx1k!L�t�����=j�� ��f�A��JL�AQ(��S���fk�Y�%U��i(У@$X���[TFv̓[����)�3�Ğ�:N�ٴ�J���2�@Q+!�d��x�)�!Fʹc҈�ؕ�Fd��I+�HO�(���&m䈫f��?.�F��F�{�d#TG�
c~���O �d�Ǒ�;�?9����i]-T 83�͑�;�d���1^�pP�#��\���)M媰�@T��Gy2!� \�R[a�1�"�Rc�o��G�߯K���d�M}��$O5$q�w,x?@��N�'~4��⫗���� A�N���D
o؟X2��/���0���@'�Q��H.D�8:�FP�Cb��Ʉ)��M��1�A,0�I"�MkN>�Ǧ��A��S�L�I]4w�z�Ǝw2By���ӟ���2�5��ӟ��'_���S�'�Dҭ����yc�%@!R.d���މ�܀$Y,��O�1�d	hH�@2Q,��P�
|A�.�kD�`U��Za0D�n�?)U�I���ITyR@�:"���C������B�B��'�{��م<i�i�u��~K���aaJ��xrif�~9#�&<���*)�,C1O�ʓW�Ű�P���Ik��ŧ��'Y�L�!��bP<�;��Xp��'�~���#����	�W��m N�T>e�O�4��-F*|�LHA^�lyBN�`��-O�c?�@�H؞"T~YE���K6;�(����;F1�)�A� ��ɧv�"�$�O0�}J�6O�iH�CMHRQ�X?w�r]��7�F��f�_�X����8B��Є�
�HO�̨F��T�L���4k.xH��"�l}"�'0��<,����'���'��w�d� ��78��eh�P�7g�� �
 4���ʐ��O���� F"�1��'��E��(O�7�B�[�aۺo�� ��oQ�[�0d3���?!�����y�1�ZI�+�y��FJ��@�M�,����tÑ9>�B��Di���O�>ړS�04�Ǭ^�`�Wa(p��ȓ@n1����0WN�����ʯA����'Qb#=�O��I d	�e���
"OLV�a1L�U'�_���$��˟X�I�4�^w�B�'���TH������Z��g��4Q�h4Ȋ�� ㈉���I�>^��G��T���RÅH3[���Y G�(!�Wh�4��p���t�sD\
D�qO�)"� P`��ы
T��@�B����3���O�����dX�P���=�j�P)O�C�I�,�\d�`iQ� Z�AΙp��b��+�4��so��)O ������{��D���h�6f����Oƈ8!��O����O��r4 bv4�l� �tnZ�<���#��0��܈��	9IL����=�l�%¿�֕8�i�Z�� T<��m+���5]D�(���13�	�c(��;/qO��1��'nB�`��d\:}݆(�����}xF�zqeC�w���?q���)Z�����̣|j�����T���=E��`��|�A���-�}إ� ;D�"p�KŦ�'��`zѠtӲ���O�˧&#���:��)*Ue�w���X�x)����?�@�P2� L9�y*�`�DdPx;Sf�\-49s@D]	yʅ�Oܠ�G�:%o1O񟼽���R�lr.�3B�5�nlie�>�G�Z�����E�Sm��74J�$+�d�zP��3C�8	Zb����rx�����Lż)��Ĕ,�l[w�"OF�Ez� !3R��P�
�d�d�WFhS6�O��$�O�m���=c��D�O�d�O�Nˑ5Ӡ�:3�P�� �	ȩx�~��0�R5 V`]&FT�H��$o+擝��	��X��V �W���/r��Q��Zbh��a~($�X�,5�]-��=��d��ywg^�#��H��r4��'��iB�O��������E:�H4D҉lG�,��h����^�8Y�R%���ت��SM~ ��?�v�i>Q%��27,�t���ACGU2I�b���Y�]��(	a&�ޟ8���T��-�u�'�2<��A�0�>Odq3Wg=� ��u�N<i�!�D�%9�2L1���"$t\j@[���aO<\14��p�ZQ�E؁lЌ@��∭e��5�O��[c̗5���F�q,�U��'��{��G�W��uk�g�Z���y��`�J�O2�yeHK�������D��EK���9��K�
P,rM�& ������{AN��I���'$�,Y�IH�I�Q��p��wh4<)FkS�<Gl��$� �O0�H�I}�Hك'`K+.|α��'r�]����h���Yԁ�S����% ךB�����|�h�A�0���+�T�>������6IS�y��1�gԓFx�XW�����'�"�!�d�0�$�O�ʧ|�j(���'?΁9&��cH�An�5Nf�I(���?��e���?�y*��I�)B4x&��'g
����V9R���'�ʔ������W�(����i#�[���;w���F�I��S�'Lwjxa6�+:����"�)s���)dZA��"@",~��B��ɥUņ�
�HO�\�%,K2W�`c�ȡ&�ڤy+���M�	ş����;k$%���ԟD�	ɟH�iޭbGA�x�~���#/������j̓~ `��I�T��� S���.�8�(D�q�>➈paN+<Or�Xb؊\;�Tq�����)s��M�ɕ�����la�C��
|�5�7�ΠyxЇȓ��<2E��<b
(���^_��'�:#=�'��g���i�/=j��|����,�a�7<ī���?����?���$�O*�S��p��k��G�vY�eȡT`��S'�$�l� ͊�=�D�uIɏg}�SNG�dB�I�?��3��2�ֽsV�1Sܠ���m�Ox���P�>�b�C�|��-� X�!�$̬Y���pÖa�2L��	�1O̱nZV�ɭ[Z^�kݴ�?1�a��ءP����s4���������g/�0����IC0fA����8�ēG�D�KU�	[$�q�#
+t��ɾc�줐u#СZ��,H� g�r��� �m��)�`�R�X�r[�n���E�G��:�����ן�0ߴ�?����@��#��Q� qP�3�ǐ(���O���S�I�@�`�{Q���v &䨴C�� ���������	.�Mk��	>.�(��T:7�rD��h��V�']6mՄ7��o�����Iǟ��q�l�	�j����D�c���)f�tx����	���9(���Q%�M<Qߞ(s�������|a)V��n�Ai]4JF���M�d�^�<�V�'0L�}4�]1-B�c?2v
�2s���zi�jV���0}���,�?��y��t��9w����	P��y�5��*�y���
�L����(5�������0<���I��$X������<I�HT�J����4�?���?����n�0\���?y���?�;_&&�ɶa��zj�#6>��,��\*u��O��[!��K�1��' �����/h'�tP���8�6 X�&ч2H˕��OPM� n��Ÿ��$����%���%���7m	��h��yB�	��?�}&�� ,�BB��JC 0�e%�fhxmӲ"O�}���Ç!ŚŠԃ�뀙SU���p��4���O(z�"
\�rrEW�&�
��H�$'�A����O���O��d@ֺ#��?��O:L,aw�<Ǭ��󯜎*�� 3QJ�~~H�*ʞ+�M��h�'ʨ�@ta�t�'PH�ʲG��K�2}ٱ�G�:���Y�����M�o\�^tD����=b�����(O�h����y:f���JЇCA*$RT����'J&x��?%��Sh�p�r4��'����g�H	$f��Ҧ+m
^Yюy"I{��Op�������	���@▦b�
�C��(��e�X֟(�I�p�������'A�����a�	�
`
�#W	)���"�U�1R��d� �O�L�G�G=|�}X���v`I��'�h�����zJ������A� ���|T��^�D+v�#-D\H��ƌ�(��Ѕ��!���`rVJ.�,(Bף����'Wޱ���aӈ�d�O�ʧX�y��*Ԣ���-�4kN*�0��!������?1� �5 ��'@�
�p�����|�%GC%pb#��A�����U��N�9�.�0�
�;�&��a(
4qL�������|!�O�T�a0"Ȝ�zq�˸>�YJ�����O6xnڤ��'��'@��Ԁ�0@"�<ؒ�)C��<����<AS�i)�U�U09P!S�.�X�2��dQ�'�!�0GQ"A\�S$�\� 
�5@��q���d�OL�$�
`3���O �D�O��$���/(&O���MB�p�l���ҡ ��aL���pFǶ�c>�%�<�ħ��D�h� #���mf8�Pez\�@����0\�� ^8	;�>q&�Ds#�B
?�Z=�1��6q'��jo_���r#���)�3��$3D4�5��Ln>�s�KP�/�!�$��]RP8F��b�G�h����c������4�x�OX`�SKKx{�%�(g@n���,��Re{�'�OR�$�O���
ĺ����?��OO��{@f�$֜���;{DYȲiM�5d�lk2��9O^�"��'#hܢA�_92.	���&̀�@L�"�X��@���(_�qH�*��P��-�B�#1Un��=���"D�*O��fq
���5�1��(��?�f	~iX���+�R�����_�<�s�<�p���W�,X0���C�S��v�|��"@��7m�O��I�S���а�����gj�T��$�O��!K�O��dm>����0�v��L�b�L HvI�fadU�E
��M�~H�"?�D�Eb�[1.v	�Ɔ�<x�${�A�r0�]�7��,��qU%�p/M��M�āс_�l�=�����8��dyB�Z�	�f(���ߛӮ�U���y��'����/\v�����p��e)�_^<B�I��MCA+��cW+��z�)������?�-O�܃0\æ��	����O���&�'V4�Q��G�p���=f�����'�`�q��bVԖl9������O�D���N1���JD�:?����`	���C�IA#�&EB@h��ݬf��X��{!x����|�`͍�r��{t���}�L��D/S�Z8���>��)@/O[2��m۟L��a����/!���q���Eh��1��D ���;07ax�;�+ϲ�3��>Zm����Y8/�L��i�R�',B%���Z��'���'D�w�r@�1��9P6ؒUn��#l�u�N	�8�DBQC��m��h�V��O��'�d!i��S�����b�z���Ҏf:x�F	�ZOHIu�ǘ4��`�`�|JP#����0����"*"$|McIQ"ST�x�<YSIQ��>�O�1��O4g-pm��	ʍa��)V"O�;s�#mX���8?}T�74O���y���ԑ|�gH�f-F!�f�G0���0�6G5Ɂ�m�-Za��'�R�'"DםڟH���|rցW>Gm����L�a��ɨD+�x�4ur�D�]�\�1����<I�ɇvt݃�U�\U��P��&Y��%�U��fq�cT�a�B�u(ޞvj�e��8�:7۠��E3�B���c�*Z��('��O P��	�}�rI�঒?*��0K�Cզtj�C�I�$ɶ� Yl�4,�3
\b���۴��@l�8�շii��'��pB��� H���O�`�l��0�'�r$Y����'��)ٔ.#�}�B��>W��ț�n'-T��k��~
�baʜ�S��< �5�h(pi0cn���"�"�������*��C#�`wFm��˞<�ۉ��G�k@B"8�d��PH��N�~<U��4r�!���b
���ˎS�`D�gڊj�!��S��5�V�D�$QsM]!9*fA��Lc�h����4�?Q����E���d ��¬L0� bq�o]�I���?1@������,U	���*ү3��_�D�:L(�4��?]2�}��� ���	 H֬����T�v�1�	����LƦ����ϔۺk��6o[�%���	�8�kV�b��Ҽ2���	�.��t�fO�!1ԭC����>�!�� 2��Ɗ�v��($"ަ�!���'[�#=�É��]�<t���P��|����0���'���'P0����ʊ[���'C��y�#�@:�� ��"�2�z���RV�h$�x	6n�3�vb>�O�)])+ٞ)��ם@&��Q)@�I���Yh�p�`��N�x�q��'��ZA�V�L*l\�emK���s5�+��K���L>�'+�;�nq��� � ���\h�<�u��\Z=�$B{3��a'O^~2�7��|�O>I6e�Q36�����"Z�})4GW�.a,�[��L��?A��?i��[2��O��Dx>���h]�LЕX3���zf���b��0_z��А%5���4��7.L�G" M�h�"ɭ`���c� ��w@�@�#D�V'6���V�pl.�[Q�iz��З�H���'JJ��F�@�E֬ȁf���6���?�	�	t̵��_�K�JH�!��V�T��ȓ.���!���΅�3R��d�c�M̓-�f�|���&OO6��O���T!W��i"O���4m�E�74�D�O�L3.�O��D}>�I�4T����$
�,.N�F��+"(d��t�7Nx}c�-�-Q&�tG��ޚP�䅘���&jۜ�KE�|af�����;k�X�iI�x��D�7�i@���$ʍ���']�p2����~��,�Q`ݑku���A	� �V��d �zK�U����C�",Ԧ�����S�~�x�qO_�e>I�r
��^��'E0-�0+b��I�Ox˧�d����P�f�5i��%�U/|���*��?�$�oހu��>5xT� ���)�|r��E7d���C�;���J�j�dMMX�zdD�r!�8�&d�jf�\�t�T(eZ�"H#�� ɑ�[����ώ!>�'�M��8�Ʃ2ҧ���Y�JZ�Ѯn�J��g���xr"L�~�0	��]��t����.�0<	��I[��m�b��:X(�!��\�J�$pܴ�?����?��G�pF������?���?���X Q剓�8�,b��:�n��H�	E��M��$@��M���4\�\��|�J<�rh��ta� @����=z���j�:�f�kD � -�6͇4g%�����\���Ӧ]y�Ky�u��΄�z*ĩ7aO�*N��fj����)N��)�3�T?��<�0.��*lhx�R!A3_o!�$[ge.�zR+g������l�ɇ�HO��?�dG;d4�h��Se�j�P���&w��9'���\0�d�O����O�l�;�?���?9��]8���u�ɥ]�V�0T�[$r2��B�iۜDs��H�e�b�@�I�0�y�B����R�L"t���GS�mf^qˀ�F0e��8A�q��ef[�5�qOH�2c-b�ڑkp�R/s�H);�d]8-���}�,X'�p�	џ��?a2�ݩL@ ��� �����!��<y���1��)����g)��F ��b4��|)���'�"6-¦)�OBB@J�b����O̳A,�'p�F|R�j�8��ag�O��䛕z�����O`��G�vY���#��X d��$,�� r���v���A���9��: �~�'Y�;��4~<�"T��$�qCvɀ_�R��,I�M�@�zt��]��&�[�vX�=)F��� �O<�NW����a�v���ٵK�I�<Y�G�N$�����ЛHt�"�B<�q�i�T��G!΃h����Bhϭ]9�����|B��>@-�7M�O|�D�|*�X��?٢͊1x������I�y����r���?���dx@�4��6;����z�TI�?Y�O��5�B�*j�d�����Ej�+L�ԉ��R�v���%21��	v���r��n��I�.9�;Y&^\�Ǘ�_HB�z���l\��O��ҵ�'1ڒO���`��,��i�3_n�@2w"Ol5�V�O�H�F���U>,m��k��'�L"=��U3��`���	� �����I!����'���'*��
E0m��'I��y��A(>���[u�I9�$ق�Gw��aH �E�\�H�c��| �q��)$��3!$53��&��%i�#�a��(;r�\(5!�L�oPN�`%O�
R�'�M�&�U�3"'(�v	�We˟gj� �/�!�'m� 9�S�g��b�#��*�Ґ���ZyC�I� L��әJM� ���:%��Lj���Sr�I�Q�u���КVO �P+����5㍒+]����ş�I��H�[wa��'���D,|XiB�M.B��
���?8!f�=T�(a�p#G�p�81�p/��u����c��G�9�/f���bpn�UR��@$ޮ�b�a5j�/�M#�M�$�f�=�feD���ɇGU�n�����*X8L��|��d�AE@E�1lۗYJ�`S>D� ��)��U�PT�d�ٛ'"�}Ã�(�	$�M�N>�C甩O��F�'0b�D�$J����b�}�aa�)���'R�
��'R8��9�b�޺p������
�9ȊBш�aV��{%J�>$����@�����?!0h�1}��8Z��K$}|~ ;�`T�d���@�&K4SZN��FaA�G�hU�ݴ#�ڨ(uU�NiT�������Be�F��=9L�q�H��8Oz݆�Xo�4�VkЋ)�D<!d�Ϡ�Ƒ���'��� �Te�,xN4��j�1ǲ��Sh(�DPb���oZҟ0��C�TB!@H�;��ɡV�]�U!P��U�jRb�'�Py8V��k�Vܠw�â?�$M��,�E�,�RQ�%�׷jydŪQkZ��IY>��%ۭF�l���;8�n�E���XRjي$η?�l;[w5R�K�K]�j�>,�D��}bn@ N�`xp	�O�c��?�`�'�;Y���qt�Κ~��=�r�4D���%������#߽_�r�@KNj����>�]���Їd�!/��iC�](�-q��i�b�'*rhV�/Fb�:�'T��'��w�܀��7,F�р��И ���q�:dː��6"d�d��/�	1�F���y���$����x 4 �(a�2��0��3h�6����F��0XU�*��8rE�Ӗ3O�H�e$l���#��Tp#R�MA�	�\���|"�Ӡ@����aK>d�*X�g��y"��7/l���V�*�L�U�W�����R���ğ|�E�F�l�k��U=$#޸���t4�2�� D2�'+2�'�n����$���|�RL��]:3��1v�|䛷�ʖ~X�x���-ae�G�����ć�JI+��F_<)�G�=ts�	����%+ߪmr� ���6��	;��?ᇄR�?�eà�߰s}t)� �VG�<��"�>vF	Z!�(�DّA��K̓k�6�|B�h�$6-�O��$��k�b�8;;�T�;�FF)��$�O��H�)�Op�$e>�A��Ɖs��:ĢI23>���u�V,=�iRW�q����;�Q��ѼB�Q��Rw��?Qn!���� "�B��ߒ��J0�ˤRj͸7��_5�xBn�:3MQ���D�O��$�E�|��p0�ʱw�=�Q�$D�d���/k8���GT)p0�A"�n?����4S*�ik�C�:O�=rGG�=���;M>A�l�-:���'�V>���7��S�0�D-εLdR�@�ß@�I�b�:�ʄ ��b!��	ԥ d��@p���˧3;R�[v�ݹK@PQ"�S#^q&ͦO���BH�V�.�:��ɱh��}�d�e����2���~���s���$退`CON�~�'N�!��9�ɧ�O�����4�9Pdi��/�nɡ	�'�.1�2��lGP�{�ᑏ8:�*�Ñ��۔E�gb
Űԧ��Р�)�?�M���?���\C�j �ԋ�?���?I�Ӽ�P���c�BXXMI$����EV1F�U��*�Z6�J�6� �|���*�Nm!��?�(�@�k�����2�3r'ECK֔���� M:�I#0���C���H$Q%eTK>iee�>�Op�p�j�o�l�Y���9�^I��"OցO̧|8��(�7X�93"�����4���O��Qc K:��4���K����b�8CV����O����O���
��[���?��O(>� ���./��@a�0d�n�ӏ�x�e�5r4�q8p`Kg[V��D��x%�)�'3�qT�@<�.�9"HW�hW(�����?���'DXE"�/$(,Ж�љ,��
�'%�0��@��	�U��e;s0$��y2�7�I)yT���ݴ�?!��TN @��a7(In��Қw^�����?a�>�?)�����,�?YN>�ā3J�68�7��#1VB�
7��N8��#B3�	�abt<��S'86�4i��>z��V1O�҆=���D��Pq
ܬRpr���L�!��G<+����'(�
!ۃΛ�v�!�$�㦩xr�K *<��Y�!b)i�"�$�>]r�9�ڴ�?����ɜ�6#@��B�x�pH�#eY0%��J�&��^�:��O�*��Ob��g~"�C�d��2�牢��xP�����	�rw�#<�r�KE�q���&K>C��1	��z���-|����IJ�`4���Ċ@O8� ��	G!��Rq4� ���))UzPf�D1ax��'���u��� 	>0�C�o�^H��Q��i�r�'�BM�DL�2�'��'��w�BPI׀�8���b��,=Z����^b���l5CNPU�����0�1��O�t���<32p0:�_�_Gz���d�>Q��B ͸Ze>���"ˍJnq�O�p�I�;~�NurON���ceA� ����|�Y�L��\�֮�AИ�P J�6�yr#��.4J�Y�n -i�XL�����d���na��8�D ����C�D)y�"O�$�Ǣ���D�q�4Y��X�"Oҡ����<l�@ �.��Ԉ��"O�uzt�Ճ~Y\���oQ�)�x�S"OJ�؆h��I~�mP.DG]کy@"O��RAH*t��lZsm�+vx�ECX�<� fU���X 1�^	CLS���i�"Ox�AbY7?��R)�;d��A�"O��$�Jo:����=Ҋ@*�"O��BT�T~2܃ D#�v�W"OJT�Cǟ&@3�Xг�ʳ-��A��"O2Y(�	A�Z�0EJ�j|�"OI�
��+٠���Ƃ2��-#s"O�	vG$ˆu��*;7���
�"OD����n=��0LM�@.�!�Y�C�.�!sT�h���*����@w!�d^��4Z -Je�D��oJ[�!��!���옄���JG���!��[^�6�HP����	3,�!�\�t�ȃ�Fߩb�,T"R�U=a�!��\����D)
�8m��%@!�0:����+#z��l��H;!��$�
����bt��/&!�d�9o� ������qK�*�
B�!�dɰM������[/ Ҕ��R�^n!�d�$|��܈�G3a��� 3���D�}��l��G2`�M	����yB����-*��E:"�N��FHD��y�6�.�a N�����!;�?�űi��扽����UD�t�����x\��(�,ͅ�k����@K��z�NM��,]�'��Y�2�����d*`�*?��B'9>�@q��f +6m�R�V۰>�d���Zvh�#�K�
	!J&`��K^@���-͌&�T6-T�AB��_s����x�JR�y1BH(��Q3�,m�SGX�o�Dxr�Zg;⅓VH����Xآ���|_�04'V(IWx�K�TJ T!b� �1
H��O���{�D0�"f�0�.=t�ܙ�D�2��}83e�C�j����׭9�D)�F'Ƨs�6�8��}��ݛ�<��O~��#��4ɾM�3��.�����׍~�+��d_��`i����򤆣��*�"��@�0w��e��!KIH�
K��K�ę8p��S��ieݛ����w���CR����_�a{�CS�j���1	׍�`]�p�^��<��/��.���d����d;f�O�b��	
>8^�+���-:�P �)�5D����� &^���Q"O?���D�C+�@���*6@���� �5 ×��� L>�1ӷP�ם�F�Ĩ�E} �'�pȀL���t5���!y���4N�h��΍�f��a0`*1=48nMRR�]#�'j��K�dR?r���Q�P���(��ʙ�&���)מ��q�'�\�'�< rΐ2��ej
� Е=�� �9S��[������5@�����g�)v.ɫ��^�m�V]��#���%�M(�#�eR��w�Ƽ
w1O���֜J��'Ҟ�s?��U��([�z),&t���z��
�E|�xB�H�(ЌX��.j����++���n�x�L��.�*P������a�$��'~m�!��oڤ?i��'�d,d��\��`+4O�&�	hI<�R`��c�L	�Jl���#�r�EAxX���Ăq��,x�iH�p�>�@w���j	H-�ޢg�
��+4�ax"�˘SPT��$�D�Tɹ4�B�7���;Muӄ�ʠi�J}"�O\A�'#�+Y���VuH�];��L��@Y!�BFX���F��L'�l��F�=s�1�e�$vhl�7�'Zl�7/
s�S�m�?d�hm�3�ܖ`Z<��PO_�PE��ԉC�U�]�'�'�����:p�֩�Krd�?"*rx��E�3)Q�̉.%��'Ң5 h�S�J��CLU.ov���O��ɬheT;���<
EJ�	�lǠ�D��CA�Y;ū@�D� �rʌ(�qO�%44���+�$w�5V��n�rP@DK��,?2�IvoN�!���'7Oތ�7
ƀB@^Lh1m��6� 0e��|#`�>E��g;C�H�%�ɛN�!���-T�@�7�9lO^;��Z��3�@T)&m~y!DKk"]X����<a־ihb���o�$h]�K���b���:��xRm�-<@�:W��5����<]N|=����6^�P���L�Z���&B��hd��;H�ph� �ie��'X6풸;Ĥ�3����r�ز����'$�+�(۟D����Q��_�f�ٴ %d�������1��ʬc�H9�>����ƛffW�	U�8�5�Uļ�C���v�TM��p\S	��|i�6뗉 s*,�Eg���4��t�g�fO�Ӥ�+[R���|Ҥ6�(In[)%��Y���=��E+E�'�T�R�	X��n)3&�$CWZ��J�17�ka��p��J0��S2g�[4������<3�~�*e�}����+�,�&��z�Z"=�J�FC�Li�o��9���A]}�"2e�R��-�	;_�!�h��y�"��¸�wm0RV�*���%<�)� �%)R�X�{k�ؠ�	�����i�
�sg�0[���2�D�~��!IN<ͧ`�6��i/����[�	/q�1 ��{Wb�	��@�L������ �]��9oZ,�p<�j��5�Z,Ȁ���.�x	�N .)�ZW�>��� ����9X9d�BrOi92T �Ɯ8U4����K6lOڙ��V����'�.7�$y��S2R砜.x�"��?щ��JV*cc���G	9�c� �\	��	'���Fz��N��B�#.��� ��#���X�[�6�HB
���+ר3&�dӯd$p�#Ι2R�C勈#���L͢P���Anm�YСٹ	P.ynZ4
21�ĥ��:593	��O��>)3:G	*�۱�W�WX�hy!\�r���q����]�|z�m��W�����I?qmR=Y�k���F@yԤ��)A���.ų��ӂ��3�)Z�޳;�`@'c>lWĴ:��X���<�퉸g�)�w��1�IBX���$.�]��1��$U��}~�ގM�ę;r�� R� �	�!	�Re���v"�#b�N�FzrJ�6����M�rE�p9�����0B�ء@@ۅ�x!A�Aūd��	%BZ.�ói�T�JR�/p���o�?!CK��A�������,�UX5raIqӈ��)N���Ę����,(�'�T?��T��ٓ̅�j�y0ҥ��*o�6�Q?}���RQ%� Oƺ5zP�=O]� O�3I0�X[ ^6�P�2�O��LrT8�=���$�bg�	�$q�!L� �*�9��S$b�L��'�pȅL|�`�l�4a{BH
q�;y���(��xӒ��"d_(	�΁y#����VfM�H�bYw�෇иVc�}��[XT8������N���G`L�qf>���%j�ɚf�PL���T�m��Y1��ޱ�P�7'�l)�ƚ1�?�b]�����|�''���!x�BA�`��v�x
�4|�]0 �J�ch���0�N��<��?���.R`��MP����GH��j����&-�+aܥ�`x���Z�`"XH�aH
�8r�pv� �E�vaSL>qr�0��x0��r�L�Q���f�=�e�'�̑yD�B<B��	!ҋ��
�vu���L ��b=�I�dcG��S�ܴ �~)b&Q�}_����Y"J �OZ�� B��=Q������Q������� ��䇽>�t�>^�8�b��Z�{.Y�c��J}��3U:\�w��={�VI8C��|R�V�8���`s��E�∈����M�5S�X��`E<Q��pC�BM�S��' �04*^��* g�
:�)���-#����!0v����$v`*��
�b�0d���[7�Af��B
1O��g�S2�d�eI�}������Wȝ��>�1��K��{�K�
Q<��á		f�t��/��O�V)��_�85#��O��S�]9�����#l9�.\b~�Di�g]+XԒ�R !�j���R��5÷�*Ip(��>I �)}��h��B�<���pS��~�NK�V�����J`BOP�<� (E$H�l��R��K[`\�UL���� ���Q�*|�ua�+4�h�	 ����"�Q�N]�;2�
ɕ26z�R�;Ek���(C�p\(a'�7LOja���S�yx�!� �M�/��⢪�+�<D�<��~*� ��5C�����5%�!�.EX�F&MJ�Es���s<8e�a�P�M�b]{E(S �?1��T?���G�+/d��с[fpd1%� <5�Z��6��bvF�� ��%9����r��;-Fi�s�{#��;�^qJ� �4�d�� Aב �̠�'� 扎c��Cg����#Xw��i�L<!�o^����G�8��(�'����i�`����B#Q%��QC
o��o^y�W����[1�P<ȅ��1��5��-�-��Aeգ8�L��K�p<�s�1+��cc��%|X�*B��|�p7m�O��|~d�j�O@��@�@ݏ,���D��x� ž���B��'/����t����J��@ay�/̫��}���a���7½X����҄�`i��:��AKrcԬ��U;�orn�AA��E�'=.%�5bF�|��ó�w�ڡ"��M�G�@*���Q�16`������';������]Ŏad6}��o�n��w�MД �g�V�M��EέqN�f
�2z�؈�cU�|FxZw�X�A����J�ց�T���%@�щ5��998h�Pf(
�8Y�)�������j��m����F����A��<� ���+�	���O�H����d>\0���׿4,����'�Y�!)3^���Gդu-H��-Ă
.�8�SE �I%��Ʉ5�H��%�⺛�$_5A4��SjCi��Ǚ�Gټe����hO���TH
� ��s��A/�����O� �ՍK8Cfl B�!Ax��P����"�dÂ�ө�=@<�p�k8�� `����n��P$��ZL��ϓZ?n��i�YD�Y0>�� ¨O�Q�<��Ȁ7�ʄYCCxwL����N
�z��\�e�4���	d"��W
�&[�x�8�ψ8S��pC"j��:%�ə>�ę��4���λCr<�B�jA�)���ec�j�(��ɨaT�P:�'+���@G�BO��U��	^8����_!^�tc�����M�U�>7J12��G��j+{��qZ�l�2H������]&�hO��X�R�lR�49��9x�1O��d�4b�K֭[+a�=
�Hx��@؅.Șu��Z�1�<2$"�>��'�8,Z  4�\� \�����I�'�d��
�V���' :�)� 2	``�LN84x�k �T8v	�c � F6(����S�W;a|b�ŌM�����Y�e��I3�M��A��zxx �)�]y��$�-����ƤU`��T%uwL�B��s1ڝ��'�ڜ��'�uxu�ۢ)��L�ef�O�KCy:�$����lT��iǾ,�f ��V��?��Ea֚4N���n3�r��?��E���y���J�¹>�@�	�_R����%3<�VfD>Kd���',ZY0�4\�	��hO��i�]
~	� I_�\r4gؽF�ޤ�e�W�`��e�Af�����i~�1�@�Տ`v�CmۘV�}դ<D�D(�+�-���,�(|�%�J���'�rH�^w?R�05	��h�yʦ�2?A"O@��mҀ�H#u9rd5��s؞k�&W�, ��s�L �z�6����&#��Y��V-8V>�b�g�	�h0�"�%A�hԀg��0<�7���A�	�� əg.�q�SaWa�<\�U�Q��8b
2#�#d瞸&�̛�h���
E�ŀ}�Nۂ�ۜyFC�	�P� !k���5�2Pq/�<("j�	q  �6)�[�"5Pw"́��O�j�@=�E�	*F��JN=D_vC䉡�*�A���)y\��`��\Ƅ���Ĉ�[Q)
�`M���$K�N��' �\��Ϗ|�\m9��%�ލY
ۓmܽ���Ǜq� �� ��D��y�/S�>�<�Z7�=���@E/^�d���'k�������O��B0'�-oC����$]+褌"���Q�$��h^(^��˗�Y���V]��"�L�'����	�^SfDh�͊.��?yb��~�l}�0L��/JH@��@}b���M�����AT�zf��>���i8���R���Lltpʓƃ3�!�	�&�"u`b͗Q��-��H	��B�ubjݷS��	0i��ϸ'#����� w=��h��J<y��l��'����6n
:�JQ���G#�l�(�'ٸ�[3Ș�j=؂��+K�~��'c.�"$��f������=�t�H�'�$��W��. d.�I3�B/9��̛�'�!�$I��h%Cs��ܴ���'��p��$��QY㑨����'ɀ� �GX(+��Ӄ҂'��P��'خ�k� c�n(&��n@� �'~z�����J8�@��	
~�
�'a<(C���	r'9 æ_-��E��'/��p�\�1����4nf~���'�@eC� ^�8Pj�� գ}���s�'��=�J8{��c'� :@�Q�'�<�Ƞ��}hl�۳gZrD��'��K�F�j錰�C�(#�`�'&�\Z�j��z�"��.Fd0Q�'~`E���~
$�T��I���	�'R�Ub���\��a9���	�'v�0H��۠BD���V �╚�'��vH�=W�rIAuM��v��I�'����@�C7��b�� $ ��|�
�'iV��1�f�PUC$�Xn��a	�'Ȳ�[��Ą���Y}����'��1�%<e�t��Њq44��'j�� f&�$m�(�4dz�I	�'�^�k��Lk���o��T�b��'�$b���6T��3Mk�
�'L�^Z�hYC잙 ��azO
X�<�v�F��R&�p��D�d+T�<��Ȏ!U�,h��u%\5��D�<���̋q�L�5�HDM=y�#�{�<1���m.�0Ĩ�+mq���@#�A�<��l�/.tiRdN�<2�#!�b�<4ICq���� �)f@X@U�\�<����":�n��&HC!�j@1E�W�<1�
5^�Pi��fj�2g��X�<��ĵs��B��j�p&�}�<Y�B�!$�lu����/	|��d�<���:҅ڀKΎ	h��B&�Ny�<y ���ErR]�w瑎l:ΨJ�jw�<� H��D�V%�C���A�T��e"O�:c[�v?dD��`��w�B�0"O΍�O����2@�@�.���"O���F�C�;�:��Q�&a�t"O��b�����h��1|1��6"O4%�u�[:YXjE���O69HܙB�"OĴQ�oM�}��pɊ�;X^X��"O�)�Q��<b}�p�&��f9t�K�"O`�¤#�J+����C2��r"O��15K�}�x����
y � 8�"O���K�c�򹈂�א8	\TY"O$T8gIC��hawKl�L�"O���$�(o^�A#kK<GqF a�"Oh�t�V ���[�-w��h�"OvMR��V�qKJ��R(@[,��"O�@*�c�>�@QcQ���M&�,�y�M�4O����v�����n���y�획5�z1��e($�^}��Ӛ�y�.T(6
H�Q�.T�
h \���ܷ�yR��;����CB��/$A�b��y���� *󪙡x^>-;4-Ό�y+9���f�c�`��"!���yR���I��&��c͆%��ʙ�y�׊Bc dYt��&wZu2�]��yrc��8<<͸w��d��q�V��y��"q7�,H�OY<����	B�yr��3oW
���_
!g���Ћ��y"�a�l㦏�dx�|2wF��y�@�1y��� �J.X����֩��yr�߲��b��!��=B�c�6�yr�ͭ/�P���,I�dA�ǌ��yr�a��܊����\����p>�O<Y$jV�,�x��t�Ni�@argi�F�<��E��p��PM�UP�b��Y�<A� PbZ!�/͏W"d<���HR�<�V	�?ޑJ����ZL��5�L�<�L�V����0�ɝ|HjD
т�pH<���;���R& !z\�t�Qh��YE!������	��R�og���>�zB�$S��n��]&N}`�P#�W�"���hO�`2�#?<|�R��k��s""O&�VH֐�\�	�)�<|�8��W�d1lO�]��H�#P�*��S)@)&��|���R������*��eb%1��؀��՞/�!򤎮?#�9:�+ʚ���c��-����]�����bԌ��% ���7,��P��&�yً҅"��!lD$;��(���y2L�6�xQǖ�����D�Z�y�,K2oO��24gY �X���й�y"n^1R�|�����ފ\{��@$�y��X�i|��Q@��w!�:�(�yL�=1�Uٱ�Rm��T�EǠ�y2(߮3A�.Öl�.�a�����y�aٳ��Ȳ��N(`F�5�2n]��y��N�9������o�he8�j��yA̧�<&`�ms�isҦύ�y­�d4Ryt�ԞH��A��5�y⤂$H�f��OʔM(����y"�&U0�"#i��D��M3�F��O,�=�O�t����=a�� c��-/�����',��o�?���b��3o��l�dO*���_���hH���Kt&�CB"OvɃ���Q��(���|��%"O���E�6jӨ�[����P4�$"O� ���T�M4Krx#�l�0:�ȝ�"O�� �N3�����^4|8!�"OԵ�!�2�Dx�"�
�z�B4�'Vy�Oj�A�Ƌj������j�Q��/��6M���
��G�W�IΟ$E��K�;�:qxP���z)b�B� �M��'񬱈r�GDVDaw���`�0	�'� `Y��K2q'?�&F�A���'��I����OLʱP�惄�(D��'Z�l�CH�0�l���5$�
�'R,$�u�G�43�펂p�̈́ȓl��lj��0cb�2R��=?a`]��F��a8�F�U���q+Q)��,�=ۓ���Yg.H�/�j�0@"��pܤ`�� F��-�6�P[e�K�4��ɕO`ثS�V�'x�����C[6a��"O��H�k�V3��2KI�Ј�"O�H��ү&A� ��-ݞu.���'!�J���[5%�5���Rr�Όi!�DC<!�j��.�
�<q%��Q��O,���R�m4�I8'̑CS�����V5k�!�N �=��ˊC�����J=o�!�D�F���PQkH�^a��F�#�ay�剧Yz��P�i�`�t);�FC�I�l���Q��9Y�D[��&4��)��$7��`k6�@s��R�����&r� ��koh���"�}�(�N�����ȓN"�$�B�7Ud��a��x�^�ȓ]�֍�R���5�es���h|��ȓV%<Q3Pb	�4D��U��,�X̆�uvuM�q\}J���H����y}:} pd�I�E���n@��yR.��w�v�X4���M����B!�y2�m�p��1�1qy�M���y�&��EQ��e
R�a_H���ۈ��$3�S�O�.IH��ܾ)rNuӈ
P�"�c��y�+/ (a�oخ/	�����<�y�釯q�d򅉊�TuR���yBE�s�F\ඣH�dtk�n��yҫ]�?{���E]-w���c�'�y򅓵�ҙB��эg>¬�C���y���d��`�_x�\�3m͸��O�"~򓯔/��X�$ߠ ��]�O�]�<Q�OV�f~��adٜ)�DM1���T�<Y�ED�E�qZ�LK�6Q�-��I@N<���?G
����9&_���Ah��V��ȓ@tF|b׆�?M�(Ë�A&(���s��A�V�;�@��ґ[��l��<�	�Q  �&̓5X�,S�]�]�.1��r.�T:�?I�F����PfĄ�X�h\����"`�>d��i�83`� ��O���#�{
 U��6]��8�ȓh-�q�aD� ���5F������?��a���PiP%`��
�t�3�fTP���m^�	�Lh�{���
̎�@��7QFB�I�4�D�ib��<�`P9PGĔ+�"<����?�x3#��5��AW�C���x�f,D�� �b84bq�����0�(1���5��p<�Fm�7[<�}+Qk�I�b�)�iYjX�H�OTa+��A#We�)��8x�T�G9O���D@*�v�Q��"��)��=S�Q�@F{*�L=jR���O�l4jF�H-\��,�G"O���#�-� ����UHV�'_ў"~��W!T���x��e��� ���y
� ��(BE_��th��p� �B"O����Π]0���r.�#O�p
"�'����e��4�u���K�Խ�b��.�l8X�"O�(Q#
c�,��͏�Z�\��"O2��u'8M0�����%V��"Od��@@ٛ��U�e���^X���^�@��)�'q��H����;T@�b��V�^�!�ȓ_�<��F�1��C$ɟ�nC�4��}ڀ�c �1��1��`���W~ҦT.Q��\�ؙ<�V�q��Ȓ�y��]�0�9>�DK�Ô�y�V����9TJH�Z�o��4>C�	,<�v�3Viۍ=�h=��̀4�fC�I+W�5 ��
|�	`�����B�ɢ 2f�ۢ�ƹD��+�$�_R�B�	
)�����ռ'y� S�%�-X%�B���F��E�B����w�E<��B�ɬdOF9��IA1Y��h@�D�1��ʓ�hOQ>�� ��#0�(83�Q����3�0D������%��퓢�A=ɬ��$ғ�p<a`N�|�
x���U;��e:�[��,�<р��O�����4D2��U�W�<� AK�N"L�D��v�l鑆̔S����>�5��i\��̂�y\p9r��LY�<�@m_�l+�� ��,S5`�	`)^S�<�V�[(�ZɊ���&ގ��$I�z�<�oK�+'���/��%�h��,�x�<�BC�V�|�良NF�\",p�<�E�K.r/�x!���k�`�F)f�<1BM�cD]R -�G�V=Z��W�<�Ζ(,�&8���΄1�h�!��R�<9�-\,�T����Y��à�O�<�'��z洜;r��$��0�L�<i2�F7r)�d��7|P���A�<��� -A[sq`�CO��r�h�<�6ɇ�uq���dQ��u��g�<am��6[��B#	�T5���́e�<9�c\�\xrY�H��Q)0L�`I�E�<���>Ect�(� A�)���H�<Y�U(d,SF	��J��8ƮH�<�dϞ+)�f@viC�a��<B �h�<A3H� ��!��;$2�k��Yd�<�0H��p�@��&�'#��PaEg�<ib^0�\��� ��94q��e�<� ��<{<�����J�#,(x�b�<1'��ɶU
1�=04�u�
N]�<	E�8*���/�.K�PB@��B�<i��&H�Hu������Yy�/�B�<Y�DZ�*����B��(LA�k"�|�<I1LSqj�a�'CI�x�Q#XN�<��I$9���heJ�8^T��(P�<��8U�-�Fmke�1J�-�F�<���,�r��(ǖl�fL1��D�<�#kA�ݶ�!�fV�N���oCH�<�V*F:�ܽ��h�}@��8���M�<�q�8{αZv-FG�B��G�<3�b4��@�W��U�N�<Ac���1��4��3 )�@�N�<�F��� ���L��f�a���~�<�w� ,d�]�!m��K�xm�g�}�<1Sc�'�8�j��Y��8�TB�<��D@�f�L�)���z� ��f�<��%K����^�]���UD�2$d!��_�6А��O�6hjdۃB�!�� t%��hʂKC�8��ENڝH"O�(�Z�!c��󄈠�ͻ�"OnEK�J�)r��P�0�J9�"O�"Sɖ�a��DOs���"O�	��뚑]B5���t2����"O�5����Z�Be@4"�S�H��S"Oh���*�^5"�Jc��>�d�q�"O`sc+�'Z��eҕ��n����T"O,Iaq%¹O:^U�B��Es�a��"O\y �N
d'j�J���,�""O Ź��˴�.�Zш�QSH�Ig"O8���)A8({� �bQ���"O����)�VH�Ǉ�6��d��"O���U'_v�qsdI��^<�H��"Ox=9�K̂\�M��]_>i;$"O����M3LT1��Lѿqp�� "O�����6M�r�3��C�
��0"O�0�(D�bi�}�J@?*�n��"O�Ȳ#ϟOs�!Sg6o��A�"O�����X�538�K���"�Q�"Of�Q4c�2^�ƍ�'�X'Y���"O��^1��xs䘂�`�h�<��d��b��ĕ�*���rv��d�<�S�*s�4�`4�Х����f�<5F�ZU�%ː��%�,� mZ�<�U�T+^�9�)����x��k�<���\�o,@�����]}28��d�<ɴNֺ[pIv�K�|�!/
a�<q������I�->A]|�"��C[�<�s�̩,�9���T�8�~]
%(�S�<is�D�5�t����)O s��M�<)�e��:�t�ш�=��ɑ�T�<y@�K�TtI&
�.����T�<u�<-����F��802AZ�%�L�<qdD� cD��T�J��Rᭇr�<�B����ջvN�8 �P����t�<)�e#ܤ(s�d��y�-�m�<�>A���V+ZѲ��`Lk�<Y�A��;���y�Q�+^^�h�o�q�<�!�G�<�=	�GΡ'��U��LOE�<��ͣGrZD�g.��\N��ĎA�<!&��r��d�U�DXAB��<�$%�l�2 q�I�_8F�� �R�<�d(�>��Xӱ�i�m�to�N�<����R:T���N�SJ��P�<��H@� ��6�IJ�R10���y�+�/0��ᢁ�t)���P�y�K�-7�P���Cm�x��S��y��jc�� E"`�����	�y���"9�Z�G�P���J+�y�f^�o�L���B�u�0���D��yҠ
����̒=���
��@��'Y��ٕB�~g�u �O �Fx�'����X�,�dx��0
c���
�'�6$��ʾG7u�a�ˡw��P:
�'r���4b�9{l�~u��s�'�;�,D	p>z٣ �z�����'�СA� \6 }*ѻ�߅l�$1�'B��U	ӎ�ҝ*��D���'Nȉ�g3a��k���h�a�'W%���W!���`�:�I���$Q3J�$�ب���ʯ����ȓh"���ЎU�m(5��!5|]�ȓ2v���cC�z4p��NU�:���S�? �-A3�Y'A�x��gY���b"O�S����Z�px���9JFA�"O����@2.�@�K@�P.ja�"O0��B�w6�@�<
 �"O1�K�2��(ŢX-�!�F"O2pذ#�U4�E"��E� ��e"O�hZ���n$ Q)CO!x���"O�5C���^q����R�)�"9�R"O&	��N��9�l�Q�����Z!"O@���ŏ�Y���2�Ԝ����"O����׸{#��pv�*]
��	�"O���fڰmBB	:��E�j��-ڒ"OXa��̍�-�l`A�U�>����b"Ob@P���*T��+`�V�tyL��R"Ol��WH�R���3fְg�$� "O���a㙷&��P���w����"OzP���J���$X⇝06�q�'"O�!s�@X+dш�&F�4|)J$"OV������T����&FH&i�ġ�"ON����@oP%�"F;vn�b"Ol�ˑ��y+�����%,�0�S�"O̙g- 5�0(�NB}k�9`�"Ojq��;U�j����G;H �B"OƬ�I9kO�5A��'`��"OX�QU$������2`ԩ//J�x�"O��a�LS�vT|-JdoY�E!���"Oj��&)��8�x�'6���i"O�1��HI7�=rP&��6��E"O쑱	x�P�h���C�P�r�"O<�I������x�A�y�D��"O��f��d�)�G�	�/o^A+�"O�� HD�N��xC�%>n�	��"O�0��gؙL�ل&A	X[�˱"O1tj�7��2gFm,ԉP"O��C�F}��|ht�66l��5"O�`أ�I+D쐙&�$l4�Xc"O�M{��9+P��S �0o+F��5"ON}�FO�{���)��3$�䙤"O4����1-�`�e��/("]2q"OLY���ݷ|�P�U2=1���$"O�<	����=�b9S��s`3"Ox�*T�NޅK%� �.[x��v"O %%h1q�l�ӍK17R�y�"OL�c�_�a��PmMkPBD��"O��J�)��L-qQj%%H�B#"ORxgeƋa)�E9����T]8U"O�$���܈GT�\�B�Chd�Iv"O��0��Dz��� �%�L)A"OJ��o��TH��G�d��lp�"OuqpM�7:���g�;*���
"Od��ƫ�8K������9*�� t"O��
�@��+#R�Y��u�����"O�u��|��4c��,	(�hXu"Obݒ��_.1Z��a��:��p"O(4*hG�Z��4E�"0��;"O��Q��X!4{8a؆���!��#�"O�;��3!� a��,U�
Ѹ��P"OG�V�2芵�ö���`"O�{�F؁uU�q�I !{ӆ��"O���Sl�n��1qcś���#"O��c�o�%Â ��l �z}�"O�Q�s��3s��t�pL]�N� �"OX���M�$��+�N�YR0d��"O�2�C5#�값uDC�hP�l��"O� 2t�tBE2/���UI_,1��#"O�!�Ԧܯuu��I�_zx�W"OX,��3?�P2�h̜*�EC�"O���q+��g|<��3�R)�Fm#�"OzMqƉ�C���Z�O�"pD��٧"O������;
�\�HUOĹ�6�@C"OF�BM�)}��ف���j�Y�p"OR���ǋ�4�N%����!F�y�b"O�Tb�$JR|�P�><9��"O�( ��Ѭ\(2U��r�ʳ"O����F�[J������:,ҤK�"O8M�p�P�@ߞK��צ%R�W"O�)iN�1>�LpiX�e% �R"O�����;�&4�a�Y��"O�0��	�.n���%H�i��A1"O(�3�j�)o�d�u瓯0b��"O֕���F�&N�� "GA5d)��0�"O��sl�2U�tQ1f�� &�x1"OT�0�,�;e���
�/[�R���"O���*XYTp��-�R0��"OH���2L�nu�"lN*ǔ�K�"O4��ަtw�D@��W��d*�"O��S��ۅzT�] K.W�({""O���$��"��B���M|+JWt�<�1�ʗ8��QpƉ�6� �1֧I�<��N�RP�IЀ��]���s��B�<I�$�X�!$ ?|�2���{�<a5"Φd�@���&�7o ���@��@�<A�!~��ya6�ȵB:0��\~�<�*�,y���Ш��D���4FFa�<�k�0h�����Ni^{�^]�<�ƸP�D�P�p�TFV.�4T�ȓww���h˄v������%gB�q��h]Ӆ�)#z��*�$6A�d�ȓ-�xa׊W�B6� 9f�<����ȓ%/��b-V�?��c�ȹn�����y���PuM�@|�� �FH�)}d@��<��%��C�J`�)�d_�q}��wg�aKF�#CKJ�9%JK8�A�ȓF%��:��٥���9�.�^�<��7W��+¬�,w�؍iR� c ���x�x���ל}�h��Q�_~zV���zؐ{Tb�!Zi�'a��l��ȓf�:��S��.[�~���oz�ń�<_����!?N��`��^)�P��=�&0yt>h�iWDNc����\.�ۢ�0�T��Ə��^�����
�(%� ��R�lA�/�TF�X�ȓZ� ���5�]���.mQB����8=�V�A�>)бꆪ>���ȓa���ɷfά~�� ���%�n��ȓS��G�Е��92�)Sf4��ȓs�1qCbϝM������&9mn,��O@��we�H��L۲ˆ.xWL4��N�(�6�C���[&��`��4��E��di�
�9~*��R�f
�[\�B��,O>L�r-�[Q"��g#H<ʈB�I>X�q���:	)��,�y�hB䉦5o�L�rɞ/Y�ؐY��GB�	�!�4�%��c��@�Y?��C�	9	\@�&��:K�������S��C�2v�xd��H�)}�T� k@4
� B�	:N�YI�%��,j��]�k$,B�:_{D|��Ä��9ٶ��)mY B�)� >�ԁ��}T�X냪+�E�"O20�4fU5k���Aj׷h����"O09JD�[(H�D��dkV ���G"OJ���Qx�����I�K�`�r"O�<�%+5��:b��|�|��""OR,Y*=i�9h�>r�h��"O�a����)ˎ �%Ia�(�1�"Or��$
F�,k0�jG��\R�"O�lb����F�� �-���	"Ozaz�mP$���)�I��=�ѓ"O���fZ�&�=*�M�?\,YRf"O:Q2抅�#I:�
�O�=;�V"OL��w�,$<(EQ,_6;}qw"O `��Ͼj� ���!�%
a��¤"O|M	�Bµh�v�I χk<��"Od��ӬZ�*8A���=)3\8�W"ON�0Z�V�6H���/�qH�"O�yY���>M�Ҭ��!�=���e"OPM���ž5�ء8A�,b�xq��"O��aӠ�;>�����D%�0�"O����@�>P�.����@�"O��� �=gOh���wy�q"O��X)χ0�|�𱬙@^2��"O�=I"m�]^����gFD0("O�Dc6�[)6����J�+ĥ�"O�AaI�/(Ha�rD�*D)�5Jv"O<:p�ar��0&�ՃA9�ᙵ"OX�`��ѹRy�@`�� Y����b"O�%�4B�n?���&!�9U�X�c"On��c��v�������ф"O���5b"�% 1�S�d��"O���#�V�y� �GO\�ohf�r"O��9���=}@M���["g`�3"O��OE�P�Ơ��Eo�|��"Oj�i�˖��ř@%���
�K�"O�	5���L��A��tH�"O��6�Ĳk�|q�K"Km����"O�L1�j��.�b ��q<���"OV�ɴc�}��xg	��S6n�˥"O%0#bR�g|���hY�4�Pɵ"O���C p�jX˳Ŝ�;�nxH�"O^�b˘T�иBd&�,~�cD"O��f���h�
��R��
�K�"O��YG�D�|4�x�ܥ�1��"Ozh��C�E��T�dfכ2�|�Q"O��k��[X�Hf�?��c�"OR�ApB�[�,8ԄA�Z�a�"O�4hp ݃x��8K�C�&x4JS�"O�q�%�U��|"��o#v�4"O�=�ʆ�Y�"A˦A�?��K�"O�ԚѪ�%�Bi{5�F�M���$"O��3`�Ɏq#�a堁=?�`ّ"O���p���y�"�n�^��H0!"O�� �@�V�Z �d���~<۳"O ��`��	 Q ���Ј��"O�i� �X��  /2��Yq�"OT�����4v��4�Ҡ�����9�"OzP����/��)��mG	b���"Ol��\51L�d-R�����Q"O %Z ) �nM�-�P�!͚�A "OD�&�S#J�ݓp����豂"O^|j#���oJ�ՏK�a�^@�b"O�H�7g��$�R�#Q��^@#"O�����&�
�"#NY5Hm>\�c"O�  =������\�q"O�DH��L����A\~@�&"Or|��M^�������-I�4��"O ;󮆗\�ޜ�+:I0���`"OJ����8�@ ��\'�I"O�\ф�S޸q��QC���e"OA�6F�3�� h�H�7"CbK�"O�83��9.fy"3E	z'"O�����Sh�Pk�:$r�T�"O��B�Ó?��mPi�����"O޹(�i�!2ܔ,��*�oN�}!�"OPl#d��k�>��IH+Mj��s"Ov���"Z9\B�@b�.R?Nyæ"O���e]:�fX�t�3H�1��"O�l��ҡX,����I�]@�"Oh�{�-�{!܁xo��;�B��"O�`डR;_��5@RmU�}�D:�"OH� �oU�UǞ�!�	�~f��"O岠����x���҇4Y<��"O�<
��iO���M^$O: E�p"O��bi˂Hl]�MC�:G���"OHJR̋Z�8]J�v)�MU"ONdjB��5%� �'g���{q"O���pMT����#D��[��QU"OpDB�C�j�����8�FT"0"O�h�	��n�l����a
@���"O\��`���6<���Q���Ӣ"OPH3a��*}0�q�.]�h1ر"O�y��?TL�5�П��ȁ�"O����� V55'@P+g|�!au"O��3g�*fX�r�mY����"O��Y5랹�zE�4��}a��s"OdA��m�h��Q�"DP��P"OX麄a�{hd����6�,�i "O�t����,H�M .��@e"Oz`��*�S��$l��JA��"O
�Kg"�!��5I�j�)9t���"O
�����V��H�	�"&��06"O���`Ƒ�5C��S%(Ծ3�^H�"OVzD�L���u�ɥ����"O�x�5�ݴ}0�4Xd&��(��S�"O �z$
;G�a+�dڠ8�z�B1"O&IB)0�����
)S��=8"O��Xgȟ�0��!�񢔧p�� xD"O@��#)R�2�r�b� ���r"O��Eև2����%��'~��1�"O�i�Pga��E+��%Zj��"O��MHd_�9�#�+�B�ȵ"OxC��`��h�C��1�6��"O��wL�l!Ѕ[ "��,ň@S�"O���#ԍ:���q䎒����PG"O��`U�˳{*1r� �&��Y6"O��c랯RA��Q�ǎj���""O�[G� 	w�Q���*Y0�Is"O0�S�@<!4����K�{A�i��"O������'jh|Ã�EJ$�8"O�xӣ	��W�b��<0�>i�"O�| ��#$�ح;�͒Q���;�"O~�GlW>>��0sq,�bn���"O\ !Ug��nO�$��A�dRu`E"O�Hv��[m2��*A�$DVI��"Oz��&��:�ƀ��ʒ9k, �I0"O��Ht�;	�"�D�T�N9A�"O4���R4P�H�:�!�VXy��"O� �|�S͓j��-�V �3����"O���䔵{\�Gn�&Aw0��"O�Pƀ<q�5���2a�8�"O�}����UCJ�D��-Sh���#"O(���G#k�Yyw�D�yX��yQ"O��ӓ-�=�:��F�7AL(�"O��V�K�:N�t��b��#4�J4"O%qmS�kH*�`�,�8g*y�"On ����E���ȓk��Fi���"O@�{�Q=..kc��1]T\�@�"O�l��O�#8�"���:s�
��y"��l ~ԓ#��;$�}�w��yR���� �R�5]?��k�̟1�yb��"0B\�p��+|rb��yb��"U~�C��?$v�B�e��yү�O�F�Aq��hD��d�Ӯ�y���I@�܂ԡO&1BP�R�7�yRE�<l�����'@ґ��8�ygB�I�20�H-A��5AG��	�yB���=������G(=7�iӈU�y2��;)��:Sn� )��x�g���y���>G\��u!,���k�m�y��ƿ��q��X�-��<�����y"ЅQ��T�0��)��b� .�y�B Q�Fh�t�ƛ�
�rAL۸�y"��;�dl[��Ƀg�"<	��(�yKD�c4`(�c߅L$�� ��y���@�z� ��S9J��m�(�yڈIm� 7y/R��Ô$+�!��c;��'`�7i*��S�ǹW4!�d :%��a�[����҂��P2!�$�!M҄��wj@uj��"i|!�[;��a�5k�fZ�({U3G!�$Ԑ[�P!���/D��X�c�A !�C�oj��¤�V)�I(�/A�a�!�_�q�(���	n ��#ퟆL!�U�'�.p6�=��Dj@-4!�P�@n�b����Ҁ��/!��=S����)âD��q"���u !�/���ؔkS��pd�����!�dҿp�R"!�D�����F��\�!���>����G�)t��Iuo-�!���p�\���h��8UnY�.64~!�#2�����O�l�R7�K�X�!�^IH\�������u��!򤒷KVi���3 �9ꌭZ�!�$��'bB ;�-��iКmj��\�!�ď=�l��
Yf*<m��h�!���vj�ȀT��R`}��&Ѕd!��-��q!��1�^pE\3�!��E*G��<���<����D$T�r�!��2,�\���o�Z��ܥS�!��^5&&������:1.�r�A½=2!��3&��J�A�9rm��Ε
0!�$@'A�a�!e9M�\��-�s�!�DT�:)PEiߴ=��B�l�*�!��;��X���-7�DyvE*0'!򤟦-~5q�!�8v6l���s�!��;K?����8f, "��è�!�ȆI��Ồ�܅C��X�TH�!��O�eC�ޔRx��FU�Ki!�$�Ne��'�b?&��Vo�+c!�4��E��a'sθ�+� #r�!�d�4�f-PB��1�pA���!�� �@Q�J�x�`�9�h�2X�8��$"O��y��Z�>\q�`�L�{��q��"O��� �;JyB���� �X�3B"O�u��GZ#\�3�g��XzԨ�u"OJm�6�LY)��� I}m�T�"O~���mѭDfJ��Ş��<t�"O������(M���	d�)j�p�q�"O���&C6�R�J�ܧh��9 �"O �@��5f>F��JZ�n���ʰ"O�i�	�?H�`�CW�*ݙ�"OV@��&����d�W~�5(�"O^�cr��"|<�Q@)p&�c"O^]�c쇰[�Vm�`.,$[:I�"O�-;�WU���l��C;n�Jg"O�eQDF8]�(y��# z��"O����3َ��\��w"O.�Ir�H�B:hyA(��;�d�i�"OTH���+k5^tQ���s11F"Or\���d4~peE x��a�"O �3�j�7�@���	1h����"O(`�'d���-@��SgP���"O�%��
�e�f���c	�7S����"O�qb+C�I{6m8��-8�f1�"O0G�8t`F��cD��㠅�D"O؄����gA&��� �#R�8+�"O���G�s;"�IPɚ+ ȩ3""O����t�<�a�vfh�"Oj �S�/rȀ�m��$�V�6"O0��Ȉ�x��S�$�.̙�"O�y��(<�B�`O-Fj���"Oxq�㈃�NmԘ���R;� +"O,]�'�����$�e�~$�R�"O`�pĂ :g���%Q%Rkz�y6"OZm82�ҭc�ԩ�ߺ^�I��"O8 
bd��i>̬��Ɩ	-xT-�@"O�}���̃On~�Z,�� �䕢'"Ov�A@
$��LK�Ꚍa�։�"OD!�c��9Qf|3W�y�����y������ ���8w�l�����y�ŕ
J�����$���E��y����>����Jιn:��R� A<�y���Nd��!\n�����y�]B`]k�a�YzU��/��y�K��@��f�8�(����y"�ƹ$P�8ق�4���uqt8�ȓa"�f&�)��d	P�[� ��݅ȓ\@ZF̵P)��҆��%uL�ȓ@��ݸ4@�X,�&V�\hi��x��(0W�ٷs�ia���>ex��ȓuj�0vK�4	��E�eKڠl���ȓ$"X����Mx]B�/4_���ȓ^Zx�p(���dڤ,F7���=Ά�;V.��pUP���	�q��ȓW��PBP+s�Jy�d�6�܅���9׭ *�������մ���w�H����' ��Q���պ-�nu��Y4� j�,}OR�3S"3����KH�@C�_9���"#ĳNU�ȓU]�Ī�!�"/`���aG_�R<f�ȓVDn�1wWU���rՊ֨|E�ȓPy|���f�D�X�ˋ'<��ȓp�6������}g�H� %sт���boXx�LM��~$��$�65�b���~-h�f��i�H��]�I����S�? ��!E� ��Y�T�\0V�� �p"OvI�eПBf���A�᳠"Onq�D�T~uhA	�BТ��w"O�$
�'��'��e�/�.k��-��"OZ�	�$5��Af�ST�DiQ"O�AIC��@����l7A2b�bE"O��x� � ���$�S1*0�Q�"O<$J�(Ԙ�@�2`l�+/ �A"OΩkG�y$(�p,�A��(��"O�t���%e{�!@�^�	��I�C"O�X�!�u\[�&�2�=R�"O>1�w�T�#̄����>m�z��"O�=�7��&�ba1@�� 6�:5K�"O�=�a��TW�8�@"��B�f��"O<�+R��}1hI��O���#�"O��-�)}�HS֎�� �"O�A�gf��dX��&��hyv�p�"O$�� H9&�h�!
�wf����"O��h��w�>=AҠ�?P�AP"O��b� �
-NXXE!ޫB&���"O4��5'=!�|:���C?P0"O�
fNY�2Y����-[�4��r"O��iq�Y�`��7!Z��"O�U�F�@ƈ��g/�:`�xɺ�"O�Ih�Ċ�(+�����-���Q"O�5肀��>)ʅQ��<��� �"O��9w�B�T�!���Y�C���"O�9��-��:�����t�P�bc"Ou[R�ʪa�(��A�G.�D�0D"O�1P�!J���8�DD�]��aiu"O��рl\[��TD��{���"OȔx��K�n���ه�M�.i=0�"O� Q�M��#Q�hG�W0cW�$:`"Oj�Jd.ȯ%���c�"� J� ��Q"O�\�T�˵�H�����u��X��"Op��7#,�
��֩W�)�8���"OZDr�jϨ'�rCH�P4e��"O��if` nf��q&I1�P�C"O@�Vd[�ЂD�>><��"O<���0A��xB��о>@�2�"ON4a�e��_�Y� �R�$f���"O���r�+i���@ ^�4�@�"OZp��j�?D�ax��J�QV��H*OV�{��Ŭ�6)"H�8K��t�'��Q
@cR)[���:s��Da�=B�'��ti=K�x�Ѱ�ȵ�!��&p x�Qf��,pp�y"We_�!�$�,:��x�@(��tC )u�L�9�!�d����p$ݪsa����"K	!�G��P�sG�*7H6D���	�!�N�tl�����O ް�"�P�-�!��^6{5�p��M�m}�qw� �6�!�_�]aX@!f�]�X`t�K��V(4�!�D�H�	�4}A�����1:�!���(�eq��*A��1��[;�!�DNi��cA�=td8i`n(�!򄘠6(b�AӦ��
rL���F�9�!�d�d,� � �O]���3�ϯ%�!�F�%
(=+�Ɍ�Р����
~!�D�3F%<���=��܂E�&zw!�DM�*��I!��!c���@'@�;^W!�F���c�?1��2sO\�A8!�I��P��4�Z\��`F�O!�D�G� �,M&��<�p�Ҿ?!�� FA�1�3n���35M&/L,��"O��ï��m|�ZG���~?��Kd"O��f@>o�B�/����"Ox�����V��Pz���e�4�"Oʁ��$�!*��b�J)!�n�b�"O&�AU��]� Ip'Չ	l�3s"OR|���zƭ�1���6����"O�u)6��U(��� � �i��"O<��ai��"��6,O�o�R��V"O�t��]/=
�$�Z�7z��w"O��I�l �L� ȃu�Z�RA��"Oj���A�`�<t3�H=2���Q"O"(rp��NV%���"Q��%"OܑD��\����Ұ�"O����d�|� ��Gr�9�"O�u�冘L�@1�F�l�ڴ ""O�5��.��	����eM��6� �"Od����#���ЧI(i�lp�"O��gMã0�PfE�c�u�"Ofa:E�:hL�Y:ed�C�&�y6"O@D)���+CD̈��%۽b���I�"O\�!A�?g�8��ǣZ�C�T���"O�P���)���Rc��g�ʱ��"O�E���{"�D�Rb�%I��tR�"Ot�R�R.-��٘� �N���r�"O��طH�$s�YQ�NWK8���"O�� 3-Da/�)jg�LTH�Q"O �#��^�{��m�7Û5c0Ƹ�2"O�H� V�+�ya�H�EV��w"O��4M8)d�����4	
D�"O�h3咓ۈ��G�N�C��=b""O��B�D�H�Ŗ3S�P�#�"O��a�E������	�`��W"O6�0��ޱf��Ε�E�
%2"OI)�`��h�Y�DM��*� =�Q"O��#�4�z4�+:vx��"O����]5��z �@=6mB`�"O��)˭J]��e��.h���"O��ӒC"�b Ai�Eg���0"O^`���
	�ܨ�vAR�<i
|�!��c&5�VoA!Dk�9*V��"M�!��:q���yM��^c6��!ı5k!�R>!�v(�B��FlV���K<�!��!h��U�^�F|2%p�f���!���%H��j��o��yV���l�!�Y�A��A�&��
Ĝ�"��W�!򄚤*@2���O&o��]���	��!��8?�})T!D%����el�!�D	+uh�}��k�*8z�Y��E[�2�!�ē��� �M3E[d��"%��Pg!��|� ��i�]��E�8�!��ۺ�a`�ݠ!>>xbՂִ6�!�D
�@8��y7L٨R&���c��Z�!�X0j�V��O�%��k3#[�!�ė2,h8�	�ݧo�fhYb�+R`!򤋝g�N��c��@� �bamZ�!�68.�Ű�	�80�A� +L[�!���9Ӥ��d�%%l�E
T�>�!�dN�I�Ą�6&�
�@�`IT	��' b��0�A9.2���@��D��=��'LZ�i�FN�Dא��R
5�diq�'WĝhU�͚Pzd�C�߭3w���'��D)0OvX�U�4"\�&ϲ�B�'����É	f*��He�A�#��[��� �}�d#��7�m՘���"O�q��,��.'����&e�d�A "O�3�h@����)|8ޥ�"O�0c ���(Aމ��Ŏ{�s"O���"Ɂa��3���R�p��4"Or|�A*�C��8X'B��D{�i)�"O�ېE�,��Z�A��-yrT�5"O�4�$N�a�X�׏�Wdn�!�"OD�����)JX�&��|���Zq"O
��d��"9�仵-�#5�T	�"O�%�'��[��i�r\�6� �"O�\Q���4M��֠�%5~
	"O�%��0rU���D���"O�$�In� X9En�(9���s"O�%�
��|���37�49�8��"O�D�C�ӂMr镊�+kȔ$"Oj��1
Ƽ ېI�f�nD�`"O�=Kvg��h8H�e
\jII�"O�x���B�E��Q�D+=D�YD"Oj��b��
S�Uѥ�@�G7�ɰ�"O�T�B띒w��X��H�!����"O�y;C�ҙuRfY��W��W�b�<Yg��1C�U�����"g%G�<AGa[F�L�!�N�>|2��D��|�<W
�(l��Q�Ƨ�;wÜ�X�jJ{�<	4�+�������:"�� � E\�<���
m�N�zr�՘�.��~�<���!)n8`�I�5y(@�Ԃs�<��m�25����hM"T�#t(y�<���v5T+LtC�!�]�<�!����)��
� �B �s�<I�� M14TqEI�Q�B��I	E�<	�C�~7@��aiMA��Dh�-w�<Y � 1a@ȩ�X�1�,�$�M�<�_� ����w��d��l��V4(���N�.�r�A� Vud��ȓr��c̏�L�V�DL 3o䝄ȓ ���Ue���`ak;;�8�ȓ4�`�BB
�oZ�ԢGC��ȓ*
"�pD̖7,���΋�C�R�ȓ+(H,k2w?�Ǚ�
Y�mJP�<��k�1{�L�R�d Ĉ��M�<��)��i(�@�`�e����G�<�,�Q�(U9P� ��e #��D�<qbFSl�8}Q���Q�ThVΞE�<���Y�SU�`I��[2�pPfAD�<y���u��X9�iU)i
V�c�K�A�<��@�)�x`"	,f�Vy�S�E�<�^;� �i!.�\����m�<)�O?qLH(�%*:�]X�i�<	�ӬV-3��~����i�<�Bg[?�NY�CA�Pr|�@�]f�<�Q�� iSܤ��H׌u T�� `�<�%�,;�@�)W����e�G�^X�<q kFB��dS�R>��!���T�<i#�2^̍��JȼcOx!dJP�<��	Ƶd�:ys� �8[��i�H�<A���1} \�BNE�3��!�}�<����ME�����7@N�P�ȓf��}"%���(w��)�� ���9�ȓea��x!�:	&��ǣr�d��`{,|k'�Y)D�(	$	��)@�%�ȓp�d��'�0W
L�(v ���S"Lpɗj�8O�|�s�P:a����S�? Y��D��J0���EX,X`�"O4�A+dkD9x4�z�l� "O�@p�m([_�1����0"Ob�i���/��z�� �{t@��"O�-;�	q��d��=��pQ4"O��SC�8I�>Ժ� ��CT��E"O��P'
������'Ap$(ѡ"O�!5U�7:~ �5Έ���mQw"OppG���R��٫���8=�0<b�"O&�C�^5Jp�ІL����8"O��ԛ)(�ND�D	�a��"Ov�9e��PN^L�o�-3�J�#�"O:��%G����H �O5?��E��"O��A����((�-܆9��	8"O�1A��	6mD�
q�Dr��c�"OB�8�H�⠣ߑ3Z��8�"O��7z�`( ��.y��q��"O���у]s���"�,��~��]1g"O�͡#�N�@��@�4��@���"Oj�D�����ۆ+������"O�0���~:z�8#�ݝS��	`�"OVЙ�'�Bܦl� $� S��� "O$�'��t�T `�"��^E֕��"O"�A�5@�q��N�J(�%[v"Ot-j�Ǧwn� 9�@�)|�"�K�"O��1�Crli��d^!C�$�"O\�a£�"X�I�*Tc�Љ�"O@��a%_8U�Z��g(��Wm��"O�����T��[���d���R"O洰����a	^s�[�vx�"OZY�(� N&4����B�D�:A"OH!)Z�w��PEM�
���e"OXA���!Ȉ���k�#���"Oθb׀	8|4>�&����ܐa"OnX�欀�܍A`
��Gz��� "O�\"�ov�d���T�%r��{�"O���G��
G0Z���.Sc(m	q"O���㈉;q�0�p���	��M�"O �5.��*26�R�X�<U����"O-�pO�3k��:ÕQLhSS"O���Ag�=���7:�s"On큳'&0pt��?X���r"O3����I��� &�;+���94"O�ĸu�Npv��svb� "O�@�/�?5��3�Oڐ,e�aЖ"O�$ېhL96�͢�4gF6A�"O�頱�ş_@�a��\�X\��f"O�Y��Q<0J�Q�a�K!�� %"O����F�.ir��)_(O��x��"Oة�%�Ȼj8V�x�Jݷqмiҕ"O$��*[�q����CO\$[�!��"O��Oýmd"|Ʉ�XX��9�"O|`!� Ϸnm@��eGU9��}��]N90�K�q'���#��@��5��oQj��܀8Wr�� ��(SI�p��ch١С��F�N��ӊ~(P�ȓi�!���7uD8�d��	y�8��x�x�[�-��%�x(���H]�ȓ�^T����<d��s��sn ��r��[�GY�D0�0�FD�m0���ȓXa�Tk"@I�I�5hw���d2B9��SYPC�b��3t����%��ц�3T i`gP�3�t�t��	7'h��ȓ\�f�G�J2�r�ABz%���S�? �<Yn>$*1Z�RU�H:C"O�X��"4(ް1Et��Q`Q"O ���*K~��2�T>�$��"O]�� �?kL;�b�X����U"O��q�E���3!58����u"O$X��8/Z��5�K�8�&��F"O�Y��)� ��x��)[ \(�)�"O� �S	� W��Ɖ\/Q#"}�d"O�ۃI���q��$D�.�(r"O<��b	���Y��E-�&�1�"OՃ�吠{��	B���"C���"O�pʇ�,��t����Y"O����m.!���#ʎr��p�"Oɒ�����Yic?^�ȁ��"OƈK7nZ}���:B��l��r@"Ox=Q<izn͠ �,�����"O�(Ie�P�С3r!�X���	3"Ov-�7jE��m�Sx8�z�"O��'���xy���`Ǚ�:��"O \y��Z*k�8	����QX���"O��0�D��=�؁a��� D���"O�I:J��پ2��"T&���'�6j���1P10�{U	��9���H�'TX	�;h�
��w$�.z6�y�'AJ��t��2X�f����=��	�'�r�xPM�%W�D�6���l�
�'jZ��C'�!���g]�|�� 
�'`�|�T������S�tv�	�'{:���[K�*�dǖB � �'@�!�n;$P0$�� �9lU~=h�'08�!s�߆\�T��(
�R�\R�'C0�9�AٶP��V�]+EC���
�'�>�(p&K+�U�Q�u��as
�'K�8j7� aH`�`OD#i��LI
�'SzY���9H� ����[2W.:	H	�'���`4ŉ);t�E���L��q�'YD���㞰��M6l*����'R�]h�n��|QbMsP�k^V�`�'Z��Q�i@(7ڴai'�Gcfp0��'��*����P2��!`���M�Vuk�'�� ����P�$ȧ(��I2����'���c��טN�$Qr�:>�8�'��i���WP@85	N ?�`s�'x<LCQ�&]y���:?����'�Jp�`�U;e�P	�b��+���8�'i�ặ"�7w�2��)�&�����'Yt�y�c�0��t{Fe���U�	�'��u��iI+�\�"�&X-b�'`�RL�h�aۅjϣЋ�i�<I�I��>��u�U�rst)�Da�J�<� Y,kA
��ѧ؋%�D����E�<�7$� ���2�����;V�VK�<�c-P9d��e�-A�Z���#UE�<)b`��r��� e,2��K�iTK�<��C�G��4מ*���k�EDK�<) ��l�vչ�bw���V�^R�<�"�մ ��Ap&�������U�<4�\oaޅ@Qoߒ�����,�R�<9�D��	��B¨�-�Ih��M�<i1O=w5�E����'t�(�b�KL�<��B�����q����(�&@��UG�<�`	�(D��㔼S�B���`�A�<��#	>zm�*5�O�,�����t�<iRC@�k���`$�q�H�0hs�<� ����,�.:����a�+Tک��"O6uz�H_`]D�ŇXe�f"O@�s��x*���,֚jd��"�"O��k�@Ґt�4	!KE/��Z�"O��`��Xt��a�3�0�ib�"OJ��1���
+�}��jW66΁c"Oܕ{���5)�dq�n�Z���H�"O��f�I��:�-��"O�ð�OC\���j�}�X0BC"O(["Kқc�|�')T[��y�"O&�H�*� ���:���L��P��"O��g�L�9�|���è|PQD"O<`�1/�TXV�j&&�CĚ�;�"O^yp�*J7Ԍ��'f)8u,K��y��xV��b��0����w,��yk�^�����)�'��媔E�3�yr���a/���vOڏ3���t*�y�&���i3�(nJx�s���ybm@���Q���!����C���y�`w���A���$�#e�yRoީ��aH*����qn3�y�^:iG4@!� {!r�����yҏ�&���6mX.r���t��=�y")ǃQ߮ ����l$�݂�&_�yB(�u�VX���I's����M�y��.#ͺYpQ�
"�!d�b�<��$͠	Y�;rk��L����{�<���:y <b���K���Òu�<Qc�K
�Q�bb��H�ZqR��Kr�<�ub�(0g����d��V�s�Vj�<�e!T6X0� �c
�	��V�`�<A�M�3a��d,��&ʂ���U��+��֗U2a�K��D%��dU���4�Ӣ�ĺR��+�@H�ȓL���!�GE�L�z6,�9��a��F���{QC�y���C%� y�T�ȓ?��؉���`�i��C��z�ȓ�41ȣ�V��
�ᡊ��چ؄ȓ	��p���X�T�<<S�m�%6&�1��[m��*�*�+��d���H�y_��ȓP�08�[�8��L�T�1�ȓ0b`�8af���X�W�&S���ȓ�
�s���:���P�';%\��ȓᨡ ��El�1V�Q8'�Ȅȓ#�0�hc�G9'KFI�Z�H��,��N�����̠P������l��L�ȓWA$� bI���T�]�7.5��x�d���ʕ[��U��m�<���.v|TӅ�<1\���&�[U�<���Y�q]�$9"
K�i�$1��k�<a�k�$Wf�L�O ����`�e�<�F����P�A������c�<遅<	��$cM�8i�1��`�<�s��p��1S2H �[��L �CN_�'ў�'|��zt��iF�Ѵ'����c�<��!ۊ3Z�|q�C��g0�Q��@�\�<g%[�4Z�Ԙ�J�a�&I�$@Rch<a���+R�����ʛ]��ô���M��'G`�C��~lT�u��1K���9�1Ob��� �*w�"��)P9z2ܐw"O���v�������&uH��/�S�I[(?�阶��?g]H��[.u�!�D
w���2��� g� p�Re�D!�S:�&�q���T5` !����Sb!�� �4��i?]�X�zVB�����"O�aU���|5*1�@��	�6�)A"O�s�Ɂ<3�.h�G�4�p�Sc"Op�Ӣ�_=3c9*S�ŉ ��hT"O,iR�K׃#�P9j�͐�J��0���'��O����T-,�]#�N�cp�ҀV{!�� #��D{����j�.L�N�c!�Ĕ�k=zQ1�mЉ4�N	�
��r�!� G���x��bFx嫳G���!�ɺq+�� lS�H,��I��Vs!�D�&�(�R�']�/^�Q󈜜^b!�=ry���w�2
�Paأ�ۡ!N!��έ?��q�Z�4�Ȅ"��-��G{ʟRt��Z�Ut����y�T�!%"OllS� =+��Dѓ�]�����"O��*���3���s�f�8y���"O��lQ�(���EA�"d���"OxĚ��ԺM�����=j� ���"O.`G띥��y��탢H�8xAC"O,��T�W�J��	@l�>�(� "OD��i] /m�E:�職´���"O�C�h_�V�TPh�XKP�p"O�e!F��Gf���eA���IR"O���iսXFl��aJ�w�L� "O�Ã��:ep	��l�"O����k!T������P��H3U"O�Y{�Aӧ���3�ti��'�qO�ɠ��p�V����k���3�"O�,�ѣ׬|z�����P�8���"O
� 0dQ�_w&�K�oO�;��;�"O��kV'��^������L9k����e�'�R�����*m4�$�6)G�?��݄�,������@��r�B�]Ԕ�ȓq&4�J��}p`TO�'A��a�ȓ�9ۤ�Z�BֲMxT� }�J���^��C��
�]�D�y��M�P���ȓ�&�)��u� )`A\�{�D���o�6e%_*o�!�SRA.��ȓU�fdB僃 ���Gт����_4ĕ3�Yl�Yx�ּI�vh��>��x��

����Nߑl��I��Iay�.��2�@L 2�ր���F�O��C�	�L.�"d�1�μ�ҡ,��C�ɞ���;E��i˨�eV�ADB�I�E�L� �e߀+e�D��MR6HB�ɹ��C%�ǘ%x"t��ᏫU�4B�)5D�,jKU2NX�sT�͆e�pB䉎xT�H��]5U�* H ���|�4B�Il`L;$G�_Z* 2�#���(B䉮4\���պ`�6��w��!� B�	#|����@ɴL[F0���,S�B�ɯl�4@�����
D:u͢B�>�<Q�2�M�C�����H��>��O��>9s0E��h]�y�FR�RP�AW�,D��Bt%�.c(��i��e���#Q-+D����o��,��0-�7���x1D.D��#R�̕B~�}����J�`�H6D�ȋeew趗�EG�u�p�۫K�!�d�2*�x��d홥w'T��j�]�!�� L�Ā�oɛ��@�H�!�G�l�쀛ᇑ�n�<��P/U�Qz!�Q�crPɣi��=�r��	@oaz2$0�D�O���&�c�Yx�쓞 n���L�\�<���@��t�h�h%���1M�Y̓SP�lFx��� �� _�TKH<{��G	܂("O������<:�z��G���G��h�"O,D�'J�*D�x2/\�vԄ�0"O(ۤ.�$1r���d��WaV|�V"Of�@���#c��0�B���4���'�&�~�k��5�!�&��|��C�I�8}�f��0�"���H_5:,|B�	�e��ɅD�(L������7+��B�i����c��B>L��NO�7�~B䉠ՠP2��O
��ص�L�k� B�	� >��E%K)c���t�lؐB�I�j���kä
�@��1��`��d��Ī>�c敻#A� ��GW�
�*Iâ��G�<q�,��h�tqI��F)px��3ŤVY�'ax����{ ��2g�_��-���ܙ�y�	�}/ܙ($hǲO���Ar���y��	7~�e�աK�>��Dl��HO��=���?9 �=�!C���6L��kdg�<��Q:eɮ��b"�((�.��)�`�<Ac˄K:>L�cg�<o��@��u�<�"9��)�ק:{M���L�<��͒lXn���FO��jI�E�<��Ζ�tKU��g�xfj�(�]�<qU)R�n���oGll�I�)�t�'?A���	y�EZr"��$fMAV�:D���tʏ�~��h� A�$�V�Gg3D��hDO5[a���#�%@"C�4D��X�KN��%G�5>LJ%ȐH	 H�!��\�dM����h���vG�3/���"N�H R�ܔzT�8�B���y	ݦ_����r�f��K7�y�)�'����*�,Ը�'[%QtT�ȓN��p0AB� w�Z�O�rѢ��ȓ!�Z� Ԟ|�2 �4hŞ)�x��=����ӭK���w%l8�ȓ/�X�$�.�(-��m�&~�)G|R�S��D��'�N5Z4��qzC�	�}�Z�������� ��+F^$>C�I��n�P!�Ľ�hJv��cvB�I+x���d�B�Vݰ遴�1*�x�IB�����.ɫ.֚	�G��c�$w":D���u/�������[����rk7D���3�B-)��Xxr��6$D]��i)D��M�!i2\{�ŏE�J���()D�,P3˾ p��q�[�h5���9D��J�n��p�9�Ŧ��F/�l�D8D�`�3�04AV��ң�,|�"J7D�tY"d.Z�64�U�UZ-�wD(D��g�߄[��p7怈 aZ��#D��9�L��|�a���СZ�`!�"�;D��1O�"U��8'�6+Uj�"6�6D���Ɨ�S�41��&,[�� D�,�c&��԰�Ϝ03���+$D��c�'Ɣk$6�1�L�/��}�bG#D�8����_Z&�r䭚�e�v�;�.D�Xgϋ7�py���T7^�U�-D�8(%
#	Ѩ�"� Q�`}�D��C*D�iT
)Fv�P32j1fH��Ҭ-D�ġ�OH�M~�!��i_�l�(#��+D�X�ЉG:#i:�sC��"/�]j� +D�����נk����F��<F�p�a�)D��x���8 �PuN^�a������2D�8SGw�e���\*h�q�*D�(1@*&������El�
u�u�$D��  ��m��`�.��1��  u𥹐"O�q@��PI�lce/�z[����"O�\Ǥ^�nx*r��eRf��W"O���%ԧS�A���@�-�&"O|9�pIQ){��xJЈ��X�!V"O<Phd����eZ3�%!�Bu��"O�1Da��+,��q6'>".�k�"Oh���+�#F��1��%�<W
hL3�"O�ຕ�<iĪ-�e_/���"O���Q
�nlj|c�Â(J��P�"O��*��Ȏ�SA�/�fq��"OYCUGw��Mq����u>93"OT`��Ҟy2��T�-U��85"Ol��7� � ܩ��A*2BĲv"Oxh��χ2v����$҃M�d�j�"O��R��7}�����Q�.љt"O@�5a)�B�3�
���A"O2!p�T'��ذ��|X񓋎�yb&Ƭ4w*5t3Gj���n�$�y
�5U�����b>A2$xS����y�ᛶn���cU�7:�[�
#�y�jD 4.�TI@���y�����yrKZ<�S�oX�n���T��y2)��>��c�IY!z����b	��y"�ڴ��� `��n�(L��K^�yB���Q,b�g��hǈ��D�y∋'6�J��sC�n��m �h2�y�`ǘ���C���~�����1�y� 	� `��%�<@�d2��>�yB,� vN8�`�n	�P��&خ�y"�.'�Us��6e?� �!����yB��2��E��@eس!)U?�y�b,�콻�I$w_~���J�y����,��4bbI�%o)`����'�y_�l��)KW/�B�ř7��0�y�@����h���<0C��
�y%�@0A�R��E������;�y��2]^ţ�$=/�%� fA��y�_�wL!�'ؽ:�nXYe"[��y�E��j�RI�UOР7���qJ���y�hӚv^��E��6g~{�l_;�yRf�@I\�(���(�hq����'�v𩒁�z�OŞ�HFW5C�X��l�w�|���'V␘���n�B�����i��TE�	z.��N�H7�<�U�Ҍ�^�xV�U�>(åc�bh<��ΜkDB�ʁM�S_���E�4n!������Rp!�(lO~p�r%0���#�)U�
��b��'1r!��+Z0-��]��م�N�>Zn;�Ӛǲ90��9D�h�X�J��`�"��U3,�a�;�d�m�l@j�D�7$�kc	8�'?�R���5�Ψ�p�C�fd݆�!��zE#�]��h�c�C!�\���[�S3u�ŏΖ:�:2|�g�ɶrZU����9��陕��i�&B�ɹ�vd��k��f�.�`�#xG� �b����8�S���-�W�'��%�u)U>MŜ�c��#��I
�K��}���v#r0��N��i��RQ�=�c�D�Y�j��3g����x�o)\��ɫ)ǲ)�H�3�ˋ��$��g$^d���[��j��<{6"�?Qa�)ܠf��u)O�g�p�1�5D����ͫ@cj�C��ȗaC����>�R����v͎|v��0J�c>y%�Tb�"F�x��6��0'e�4��K,�Pz��F[c��x�Ɵ�(���O�9�&�b��9�I#{]�p��I`�V%�! !DXsb� !.����$��(� !X�B�]��K��p��,�� ��Ua�ޢ}sR(7�q�����ji�0��<B���yL%p�/��4��'�2�b�$&p�[�&؛C����#�IٙF��0�'P6ҁ	�hҨ���#JRz́Q��C�,��=���� hX���r��;���36�2%��Aa�)>���_=gj�ɘ����2A�8���c�'Z:�`���ZF��B,9=TP!�yҢ��<7Z\E~���?���%��dS�CPA�'Pi��I�#Y���eO��P��?��4�I�`[�k!K�|�) V�p	)������Z���8U�7�m��hT��H�ڼ����(k��h���؉Po�<�dY'>�~p���A����8�fJ�JC�e�S�6	:�	Se���D	�_X��a���U�>���^=F��'��m�Ö<y�1��^4�O�5b��Vk��HT0��	�(ʒv[<��!fʲK�V�PSAZ�B��➠�P͍��ħ`Ҁl���c8@q�`
\�h!v���x$�#�#�O��Վȗaшt����>f3V))G P�X冖��56�	�� E����`�[�bѪи'2�=a��'7ҩ�� �(�l�2��N9b�j�:���	��&�H��D�)`Eƅ�� �+�`�1b-ը�����Z�0L�ѣ�s늹!@��r����w�� �J>��ʦ�.�l|��Rr�,h�+�D����]} I7��S��3DP>��$�DI�G	..:V��@4T��';P�+r��P�����|��'Q��R��M�M̺|�pE?2����E0��I1L
�X���A B.�����ôh!Ȕ��'�DH2�ȡ(�(`a�� I㊝b@mӤdŗ�j.(�*`ɜ�WT��@�˓EQti�^c�D��נ�4_�8�k��T��ĭ��'�
�� ��}h�(�� ?L�d�/�ƙ��Ǝ��X ��2hH����\{e�b0!;H �6$@/�^��,d�>�e���H'~��R�'�6�!���O(`���͔ �<�˥�R �~�bt/$p0�a9Zw4) ��E��D8�F4���GR�v��>AV쓱�hI
�"@�3�����l�ɟ1��ݰR�D�c�$5#@I�C,�	h�-^��R�oQ��P���kiP�QU�0y�Ւ�eK�q������=�g�Ϡ$<���B��a䶐0�\+|J�822ß*�t�)6�K� �΍�$�"!1�ɑ�V�e㺀h��3(B71^�ڶ-��N�4�9��Qqh<�戙=@��р�Ś�q*>q0LO.V�����Z]�19�"2���
�H�<D���e%�t#,Ux�l�R���C� O�d�y�V��i	�a��$�4��<�fl�j�M�wę�S�x毘�����,L��!�I��{��͒A��>K��t��%���'�e�^{�'�Pq��F�l��Q �-!3�!�N>a�Y�";��f�Ԓq�pt�&���r�c]!n�J%	g�	�]|!��-�: �8hcb'@/\����A%�#l��}�6�v�Z�NZ�/5�
�g;8	Ë�+R�ᐢ�ЬG��Y�Ð�yr�[*<�"���y��ǡ�@�Y͔+u-�T
�	!��x��B�R����пj�n,�G�	F�:0�1�E�K�ƃM|J�0i�D�� <m�p�d��A�$�D[�Y��#����t����`��yC�ɀ@�'�f��)�u��#,FAc�ץ[+"L(��@�N�� շ`da�E�uW豄.
�*X�=a�@�IV5F�Ќ=x���ʔv�I�?v��A*U�N�Ya��0g;���!F����:[l���G�+��y����g$��cEW�v��
�c�]�P@�[�h�K�A��?'�)h�@��

~�5->�E���߃e�G�\�r����<!��;9��d�ن}�j���j\���^�f1
��?9Q<�p�MY�Eni��(�!bL���Iuڒu*�W�o�l-J�ٽ?^"�(W�$Ht]�6�'����ǹ�H�"6�[:M�r����@�����K�l����"H��Ɂ��e�څP��űK��t�����!�J��B ô�U��q퉙w�	 �a�{0�lRee�E��b�dJ%�N�A���уvH���#�RY��)�n�d1Zt��*�18f%�G�@�A�mB��2����>	��Nz���B߉k�4ВS�,������9o.���®?��r �ަ9 ߴ{,��� K�2��nW;ks��A�W�-���d
H�n���D�p��U��T
'{@T@!,�+2f�PW��/D7-�Ȧ���\1�)Z�%�V&��i��D3?��h�5�'Hf�G`Fa7<Là�ֵ"�� �ϓa46P� �7$��<�t��xN���o�#NV�(��]���������4�H�Y��e�I��h˘OA��is�I�%e�+3�_�!ԅ+�b��|��OЕ�BD�q� �&_95��Q࢜;5'L$�0�}�T�B�<>,� �Y�W����K��I$�=��CNx��j0]%}�$A
��y`w�L. �i��@2J:|�@i_�r����'6�C�:�à�ۼ��Ƃ�UZ�3h�m�����x�R$ ˖�ȳ��_.�����\�6aB����<�Ųi�0���K�#a�ژ:�F���aЏ�Q�	�ƽ�1dE�&l�k*Pj���ܘ���[�N�:���`�!(w-Αk�,�H�l=�0�f �q�[�L;��@�����=)v@6�hO�Ԃ����^f�ba� �T��٢�|r�@9W���r����@���3ua	*%��a$9q� J�%�q��($ڏI�XtʣG"WXń���*�x�g�9Z(�a��s�PH9�
�`t<�1AD�(��cwHĕ�47��u%*�h��C2r��̻
s��!�.��t�O�k�0I��c��/H�%�wS �Z�Ӄe��,���Ҧ��@��!Q��Q@L`*�#R_��8*E��%�y��S6�V!g�[j�H�KP���p=��@�V�h�7� �H�F�(��;i����ԃ> @E���RG����i�K2&��ӠU�L2 �P�	<�f�ҲȝVu0͹w%$4�Z�ԛ��Re �����WzO���s�?.�6�q&�i�p�����)U�ˑ�%�D��(F��̃��'�+��x��B�D�K `�`쁲4����7n���^��� 8�0C۴?���� ��u'#]��� $RdlP5��Vo���&T@"OjUQ�K�;m�L�"o(_v�y��`��m��'�����@�jQI���>f�`�ЪZh��'���0 ��V�A������:�u�f�ڥ���u�ܡ[fk<+���X�.�,$sLy���ʾIPb���J	@�<�
��յ ��DE��'S��;@��o��\�T��!� �X�}�
H94XP���X��j�E�)���;�O�����6@0x�zGA8(J҈9FY��!�\���匲({�0�&B�Laƕh`oٰ8[��rg_�Ua:x�D��	�y�eL���ilށ#�l��4�䀇��(��TsB�8D�(��I $��aJ����f��C�[�k��x�8O��9f`̽5�瓀%��qj� H���_.����##��񠰏�sΦ��J^�1����Ol�@�D�cQz�`"�ƈ:T���elL�L� v%G' h��S�/<ON��X�V����ү�Qja��	/�������}�v�r�H�~��d�/Sp�P{TH�[i��Ҵi�h�<�"� 8~����]�;��9��L�qy��Vu�⨻��S2�����6U)�����4�	�B�l�<Q��K�w�8�;%�������A7����'7@)9�����Ϙ'�a7�C(z��{E��`�
�'в�+������E�R�S#
cp�tM͟sy�p�!/=�Ou���=�d@)��^�T֔�Y"O:�C�[7�{B��l{�]�"O���tC�s����&�k�%Y�"O@A���s%Fdh�tY��؂"Oy �b/�Y���^�4ễ"O�,b�B�$v����cޏb�敻S"O�����>��-�#N����"OTI�ă�F\r���3�.)"�"O<8���>���y��7HŘ�q�"O�E�@ӜKH����')[�a`"OX@A�,pp<Xe��]�"8H"Oę0OT��=+��@��=K�"O��KF�b��|S�ӭ�I1�"O>�B�k��X���%߀C'T4B�"OT�h�@T2��cdoɑf4���"O���q& �r�P��X-n��ja"Of8�N�a0I���ōb��8 v"O>HY�b�0>�-H���2R.�z�"O��z��I�2ϐ���^ 5�ʡ��"O<�"ᯋ�4+� ��!�
���["O���Wo�=W�T�֯B��D�"O~�`�j�b��4Rr�]��$	i�"O6�R$hLǜȸ��F���Ԫd"O���D���fMK5����P#[�<�S(�QcLvd�.q ŀ��i�<QG+C?J���s�쁲B���Xs�<YQ�;NҊ`� ��^U0���"LA�<Yg�b⤣�V-yD>,�CA�<�ìX>��7�[�"f<=7��B�<9�$�,d4\��E:��UDm�<i�F����Ga�7E�R�S��v�< AETt�^(E������p�<�`ѣR�`PLгf����o�<���XH*f[.hC���tn�@�<��̛�b�,��b���0��8i��T�<�!oF�f�t=RҬ�?Z�d��XN�<�G �<.����^VR��3r$�J�<yD!ȡk��H � $~е��fLD�<Y���:_m�U�äƂe�t��]C�<a'H���l��D>;�Zgi
}�<y�@>`�����5B���h��y�<�EA�'��Qq1`ÿ=��(��u�<实�Jo2,A`���@��1tl�p�<ٵ�ȭ�^0 ֟Z[�%����W�<a��R�7,��ڙ^��;7i
v�<AĈ��.m�LY�iW-/�nQ�$Pz�<� P��b�5�2X#j_6p�9�"O�<�@	3f�С��U=:�䓅"Of��!i��o��%�݊t�FU��"Oȁ@7�%U(� �+ɤuf�is"O.Aɦi�)w�.y�3J�%w�4�"O u� f�3p8��P��K<��@d"O*=Z%��j@�̙ը
�T��Pq"O<$��K�G��5y�ƌ�yA�"O��T%�]��0sc�Q�`�ĩ�E"O���uI]�D��!�qeӫy=�"O�����&����2f,H���S�<	&��-:V��eR�0�\8�$-�E�<!��сet��Q�P6<0l�㲨GC�<y�ΓCl�rצ�'����G�<�b���FX�=�HD���PG�<!b#7�����*[p��t����B�<Ag�ۊ �&�85�*`_n���A�<����D��@�q,�/9���7��P�<-�(q�e�z;����F�J{f��=�Y�pF<^Fs�
�9��Ɇ�#��Ǫ�w�����+'N&(�� ��(��
�U��P�#GI0 ��h 6A�V�B�ȳ��J�\^�T�ȓ��h2"�0&\�C���
Gک�ȓC��A�bE�8��m��#Y)t�ȓ@�$��vDK�
��,��� $o���ȓ[S��l��lr��P����D��VR� 7
6��m������ȓ~��,SN�򨊁DCJ5`)��_u�yf�?���i�@��j�"Ot��qA��p�X�R�I@Ct���"O`#�6<�8�U�?F���"OHwI�N|!kwhۦ�F=Y$"OԜ"bO��Z$ ��aK����A�"O��0�B�T��B��E�U^��@"OF<�$�:P�0I�s'��ER�"O�HI5�J�^�:]��!&#�=�Q"OJظ�������4-AH�"OZ�8�H�

��O �6�N�9�"Od}2s`�A}%�Ύ�k�͛�"O�R��N�8!h8
f�3<|�Tkp"O�s�i����IwlS�T��
S"O����F�-j�9�
[�M@q�"O����Z�>
���HT���8�7"O��XBe�9�oҵ]1ΐy5#D�|�RKJ��T�Dν4.��7a5D���W��((��!��M	������#1D�����Y'B'Xm(�(ĥ��LP�,D��s��AT%�e�D3yIȤ3@�(D����@E�"�!��c� ���3`3D�$˓��O�̸)���<c��r�'/D���
*x�xHzL��q$1D���'��kֺ�S��J9NM�҃1D���C�F$x#�o�T�Lq�֬,D����[c 1qτ��� 
#�yo�u�F9���\�vb}(2Ǎ��yrO1�pWi]4J$�����y��	3i��Z���#кM���]��y,C1$�ɷ���>���カ�y"�[���B"�)\�A���y�iO O�����ν/
|R&�%�y2�ܔo�ړ䛾� C��["�y�Ε�W�RpQ�B�

vֈX#��<�y¤�'|��ZщգxĜLc`�M��y
� t���*F�BK�Dk��T�B�֥��"O�@�BG_"8�C1�2_��a�"Od1H���!����U��"y�dڧ
O ���
�ڄB��\�]��5�2��#��P���(%
���d��.�u���ҲN��cb	@�ax�'D��%P�.��N�&X [��Z2J	\����B�7c�Q�ȓ��a��Y� �`�✛*~��'�`���C��ph���GA>i?}	C�F#t�JU�֫X/6����#D��#b�39����+6S��8'O�.9%!�͟X�V�RC�	p����Oh{�O6`��`��`�dY����,J��$�� �~�'J��4�v ^�m��t
W.
a=
bJS�UG����a��D�bŚpF#��=A�dqƽ�f�)�P�QQ�H>@ Q�;Po���*�|�0"O:r��@����(< Z4���i�9:!GT�C�y��ڵ	:��%D�t!T�Y�K=��P�Fy�cAC��]���X��a��Q1Xy��I;��0E��D�S����yG@Β�`��`�I�<6�(��Ik4�h�D��QT��4@��A<V#Эґ���#O����n��C��+E�����cB>I��ʧt�~b�|��7&��!7�q��p�+)�$w��8r��%�mS`�]��g�\@�9��/V�F:P�c�!75`��$A(H=|y�A�69;^4J3ÀF؞H9'���;-
e��f�*3H��E�v���c�Q$8hPlZ	2��Y���RzD(����X|�xs��+�k���t�
���B�%�6�
ǨN$Y��D�~Zn@[�& ��Q��M�,�����Ƿpf
����Z �ʨA:�iف�\�\���-�5��Bc_y�]H�G��d%��፜(;x!Cϓe!��Q-]�/4f'X�2��(�1I3���ו �A�1��|�4�D�P�}�daqb�
:�ר�0K7c�4��/� �,� ���	KnL��"���
L|`rg��(�)��!��5��$F�rx:�"��;^P ����ՔP�p��T�AZ�N���e)[�TQ9%o�{��x(0�� ^�dM���'R|܍a�B��5�u,�/F�a�g�v�6d@�Y�X�zq���QzԉqW�c��A`.�~m���1 ֱ���44�`SAH��Xr�C�ӸT�]���O�xl��8&<�{�,Q� ��P!膔]y�س":P�y�q���jH�e�)<�ɩ�GV�8bbd;B�gx�̱����<ktPC�åUW��Ҵ���2$�T�N�8�T	3��
Lg����M��IN�8�3�T�tT����ޑ�L�,ё-�&`h�⒠,,p:D%��R�.*Pr���h�)���C`#4=�A$E�Jx����=odM�!cR�e�������6 �&4.=��	�/$��t�Zy˲t��A��=G�h���øNض�g���踉ӄ�'(	:�	�ǤP����?@���{�@�Z%(�dȅ�2�Q4�
C㉈sn�i21J��E� <{H^x��awf�'���͓F�(��
qh�Mj���B� ��C�Yw����a��x�H0(�p�@��W��ч��0*�~,��CJ�P���cցZ���5�4�<YX$�*@��2�P/ۀM\D��u�.e� �!L3	�Ќ��,�"�AuCC+{���I&
S"C��'���q�j�D�����̃�S8*����b�.Γ�p��B"�u֬�(f�X�v�`]A�>(/�<j'�:�Ol��C(J��� �X�)�,�R��ǝ-� ��ԫ݊v��«C-0�v�͓M�ޥhG,��*� �j>�̻�'��ܴk�*\10x��SO�ܒ� _�|)�b�*�.L����.Lk���'-�y��*}lٺd恛T�@Q&\,�4x�gA����·qrP�ظ.%���1<Opp�G�:*.��hо^R� a׋�&���+��<N����r�\z1�=%F@��DI�)�('k@e�'�XP��p^��h���GF�i�� �'@Q6�a�
ʻ(B��7yuȺS�b�2�1R+ٗ#�v�k�a�_@�\Yc
�$��Qq������>�e��i�Xљ�7s�Z��!��_Ϩ��f*TnLKI��>�(���馍�۴��aZ��F0E�nܜ8 ����(~�f�S�$��B\��$�.��0��-4' ��SKGMO>�[@?�7��Ħ��B�J6�P�f��`�Ψ�k��"*�D�'ΖxE��,=Z:D�.��K���<ٓ���tDR��+@��Dze'�{��k0�)-�����kD4pby`�N; r���	:m�Xp+���tў��!'�(�B	'ƑR�����!�dƐQ����3(@�}\����W| Qk�(8��I�VS�4���
/"|��!W���y��H(����I���9����6W$��YPLɇ���`I]�m"�Q�"
ʎP�@��?�y|�RT��`�VM�;{�<�D'b����l�P�A�ƓF^��j����e�\�!��H)�)TeݮU��I�M�W� 8����Ej >����A��L��H�O�H7���4hC��	�A����<�p�����=x��.�l�c��-��-��cT�A	R�8Ab�Qȩ�*�-6X�bd�
)LCa�*�ў��Uc\2?���e�
��ػ�N>�D�>����0��X8ܙY��-_��� �N>��7M;�eN�%�^���^�\p�PccLZ�v���c��Kx���.�BP��)]� l��h��{�h��9�̙����%M��-��yӚ��cR8W;(�T��;'�^4"ɔ��bm�����o�<9�,Kz��@P�FC	(�F�!e�+EǠ@�犎Ħa8!�Y�>�z�
UY�-�F��P��_��ҳ*W��yh��G=
8[��J�p�B �g���p=��6��e����# � �8�֝m�����탋�wn@%np�v�*� �� n�x�
�@�����8 �Oҏ0�JMzcm�_�qO"��F�O-uW(X�%�z�`�9�
nH��B�4fYecޞr; 5
 (�Fyx�U1��!�YW���Ь5�p�!����8���e�)
� d� ��UTb��q/B�\[��nZ�o���
�Ϻ㇁e�u#�Y��
!��$=̰m���,D�H����' �\��!����XX@c�	��L�=O D���;HȀN&�J�YRAA6
��d �O��GJDuI�z2�)O	N ��'��
2� � c]��&H��KǾ=��tUbM��0<��C'=�f��%U,Ĕ��3��O�q)u�+P�x2��8a�X�d�ظ(�0Œ�E�	�NtQ)=5閝�Y�p+��)�z1ܾ��	��`�nC�ɼC�,�!T`Ь�����͖�4�I�N�I�M�:c��c@�I�@ �T�a��SҼ�EcȎ�b��w ��}p6/r�<���&�Z���3�B�sG	�/�`�PLu���lE�ro�ͧ'�\1�lG.0ȉ'"h`ò�6Y愍0���vF�y�	�~�a�!�Тx���O�7�0��t���@���:#���� 8��J��d����Ē�8�� ��.P�`��HKRL��cf���aTę.t�\[%�ړ`q�u\q;ІͭE5*��2.J����O�Z�����fw4��I�2�0<�'Ҝ��(�'6�|����3��$.*�Aa�92�	Rw�)^�0��ȓ|��A`ɕ9M&\[0I"I�\��'ZX~� R F>�H����y�nO7�3`bďfL�	�"��Px��9$��qa�Uʌ:��+2F�8�,T���Y�^%��HEP�N�څ�&�M�~�!�D[�f�,�gT�M�Bı�(	6�!�$_8y����E�Zz��6��a�!�E1Q��%31�H/^u���©��V!�Dܧd�L9�HؙV���Z�BeY�'�0�{E��=Pk`�XB� ���0��'����F|aE�ف%�P�xu,X��yRf�AR��h��8'��� G�S��y��C:'X���c 8M|�Yx#���yR�_9=�����8����p�X��y"��+L��&Q%�DВ�*�ybiL�/kz��4* ����sG���y���l5�Si��{��tX�i��y��$8�Ah�Ό�g��i���y2.G�Y�h�Fk�f!�]��IZ��y����}[Rء��Ѿ
��X@�&�y��E�:��Q�nєt�T��/�?�y��8d��D�EBb_�]�T ���yB��\��[g.L�f_$ɪ�f��y���=|�`���K傔�Ʃǫ�y"�\�N�ڴ�6 �W<IW'�!�yr͋�!�nH)w	PL�~�a�J�yR�K�(��%��ÆO��1A�0�yR�A�����X�.��!��yR�MMR�P�g��Ԣ�J [��yrI��i@�PS!#�[X��AX��y�ܢ59�({G���H��J�����yBK_�=PTM��mߐr����_��y�°i�da��Ibq�᷀��y�ަdGf�򒈅�v���1ĂT�yRL�!�P �V�?�J��.^��yb��(�L٢3^1 ���g̹�y2d���\-:��4dmxUP3���y���pXU8T��Q r8Jb�9�y��Dz�iѣ�Q׼$���y�M��D���q2��%�y�q��6�y"�\0E�$�ǌ�5+[8,3A��0�y2�=f0��xP�V'0�X��$��yBIO�2Qi7$�zA���y��ׂ8�)�4m,bi��z��!�y�
ܱcH$��â�,�����
��ybC�����ɨ
��0�C�y
� ��S�
S��(@c4 ܾb����"O��
��9�lt�'�Z����B�"O�DI�Ռr��X�p�2Y�6x@�"O�#�%P��@$y�횽�9�"O(�sc�8���%Iæ�(T��"O�e����?.��0���O�BuJq"O|��s�ȥ0�.����7���*O<�`%�}#��8�?K-:�' Ը�B^�E3 �
�� �(��
�'鶀p�-9X�>�IQ`Η j�L�'ir��Ëp�#��
���l��'r�g-�*,�(˖�Q��.�		�'&88��Yf���;#B�Ie��I�'DRp$Z�� �҇�0F�|�k�'.���J��;R��j[v�!�'^@�A�, 4N��@Tr2�ȃ
�'gu�q��Za�ek�+�kq<�	�'��!2 iЃZ뜝�ҏ���q
�'�>|���HVX����
#�|�;	�'g����`Y�d��Ђpm۩�x�x	�'x~t��jB�A�4����y�J,�'vt(WKr\v���ٗ��yRG��s�^q�U-6@R �Q���%�y��WF��$�8n*X�H��yb�T"��5�Bn�E=d�@�i��yBL����(GBڢETR���k�yҤ�6�@؋��SjL�;U�Q��y�O9:`{׏ˤz��4E�y2B"y0�DaD�L0E���Z�y��T�\�0IRE[�	FH��`���y���8GBl*��=Ux4�Em�;,|\ȉc�f?�҃q��Ê�4�OY�i]� x��G�U<4;,L�R8zX�х�<Y��00�H��I>��SM�jI�dp� F{|�@�G[M?A�ó1��S�x����O��ۡCK���	X�B-z�J� �;;��"k� e�*�S��|Zw�$�W!�3����Bt"��Ip��`b��A��ا�	�4'���0UM4'�5eG�:�O@]����{>)�t�{y���ɔL`v�{�N/�$ҩ'���z疟�A�*�ӳ]�,�jB��2Y� %aT�ԷU���	�:���	Ic�)ڧ*
AZ֦�+o7 j4�(>2�m�H��6�M�S�OڸxXv˱H� (񓁝B�Y[���Ǧe�<���OʱO��&r��}�g .��S��#��6�X>��	�:ٌʊ���uW��T���eA�4Y6����۶mt�1i�h�ߴ�ēK��d�"�Η-6T*q3u`��}I2�!1<O~�jS�R��M�K<E��C3(8@1��u����@�a?ƅ8��C�c?:(X�Oa����#]��Y[�b��i��MQ�JL�<�%,?�Dժ�>��O�P���$���K�n����D(%�ɍ�����������CӠ�°O�j���1�I���ɞ%��i�C�S≾��O���� �?R�cvG C���ٴb{>h�G�s��L�ȟr�{ta��UQ3�͂y%��rv�9Gt7@>*k"�dӞY%>�D�<��	K�H���ئ���&��	:�6�5��S�~y&��X���4�ħ$8����ǜS`��HW��Cze@��޾P�~�1�t��Գ ���,Y#c��,Y��#��"�m���53�l��%X�r)�h("��6o>1�O� �:@(E��� a �L1V�`}Q�-)�Pp�IP}ˋZ�L�ʧ�Δ!t �e⠩�g���<ņȓs����Ƚ��H���ԊE�E���ڭٲ������'���0�|��ȓ�0�g��TN�Xa�C�+���ȓ2�(Kqe�F���!�KF)m��I��v.�e9��,���8"���z��ȓU0�H�ׄ�$@�� �,htm��*&�!�9�0
@�?려���� 6�K	,�R�^�����*�� �S���w^�9$ǀ\1⤇ȓv�*��Ec�~j���^R�E��S�? �U �CC�i������<{8�"O`���bW�7��u���&O�E�p"O���� �j�0<� ��g=fPi�"O�8f,ڌz�J԰�8c7n��u"O$5j�����Ph��	�'&h���"O� H�a�w��|9��.&�q�"OP��4�^�z����!�����zQ"O "N��rl� g
Dl��Mc�"O�L!�땑 �N�9�RBu̽�"O|��+�tr�Ň�=�$[�"O��`c�7Y���ȁG�KT�y�$"O||�Cj��_�vX�T�M4k5V��"OV����Q�j�֡v@�,AP���"O�i��h��n�4�j�PZ�V�:&"Of����
>T� H��O� 7�2l@�"O�d-ı)Q��ʔ �kV֔ku"O
�+�B9%`<Uq��Q[V��"Ot�q��JBH�:��*uV�� "O��rC�3ep���cC ���"O��P�
��508��F@��X�"O$щ��P R�k2�UF��B`"O-:��Z�5�֐�B�cҜ��"O,�ۅ�	8P�i�W� !w����"O��r#L53�>En�8D�А�w"O�(C��k�Z`�٪:�j�[�"O��q-ɔd���K��C�2q#�"O��t��<��`�ˀP��z""O��rF,S�Hthk0����yɱ"O�B��f&HdK��5�f���"O��vg�<BДZ�䞬l��ՙ�"O�e�#eIu���4/�8C"Oj���ț5T�xU%�(
��u��"OJ�ǩD'a���:�I[q��h8�"O�,�3⍖Y�=�Į� ���j$*O�L9R/�a��[-aL&iB�'w�io�4Q�n���B�	���k�'�Z��D_d���E����#�'`i�g,�~S�
Vf�l�}��'���f%Dz׌���N�2E`�'ܸ0�7N�6t�fiةH�6HR�'�TP��^(���fԒF�����'�\�Ӏ�pkn�����-�HT�
�'���:E��Y-:�dFU�,��m�
�'g�����P-jTD�أ*(U�t��'��P�K�ar�b�gI�K�Fl��'������`��J��@+�'����î��y��� �MۀNܐ���'L^ ��`P�Йv(_+Ka�tC�'|&i㤂�"n�,��j��5)���'e�d�Q� l�$+
'�,]��'3��۱e\'N�xX������ܱ�'f�\@Wn�<=����7�׋����'���ZS�M'W���aT���ra��' �J����FCx��fa��f�~DC�'ά��+֧[{���
�t%��'LZd����;p��I �&I�'&%@`�>Y3��doB0���y�'����׫�*'��%q��]�xv��'�	�T!��L~�D�,�1j��T9�'!J���/��0������{n`�'
���a�w����r( ZG�ظ�',Vt�!!f�L��С�a��!��'["DBQ��&���i��#C����'���R�ÐZ\-[SH5��![��� ��*��ʸi���b%��L�\��"O|Y��� R��Uj�"V��� ��"OD�	�'�&,�S�	�K.��q�"O����(�8J3�޷!j��"O:�ʐ����`!�u�ްBzr<��"O���צ�8(hݺDaS:K}:x�@"O��1�9�D@�n	|T�mCp"OF���9F6FU�"CO7cq�Ġ"O�� k5���!Z�m f"O ����ۂOR�l���-!O�`
�"Orlw���ؔ.�yP���&"OX��"�
�hTR�f�C�
��W"Ot�Sfǖ.F0������5hl.�S"O����	n|��X��>��a�"O$�c�%ϣ%�3c�ݒE�8�3"O �{��X����E_�f��x��"Ol9�u�>/��PQ$*]�+����D"O*�Ɣ�b�����Q�u�m�a"O�����JD��&m[`�{"O���L��;�Z��$MQ�E��u�"O��S!R�ސ�Cؒ&���a�"O�O����ɍ�
�T�z�"Oh$���K*�8�I�Ar�P�w"OPT�b���Dx���}3x��"O�A�2�_,r�b�����E&=R"O6y�*��Hf-#2��?u�H!�"Oa�uO��z���{@�={�B���"O(�xf!�/���+TcbxkQ"O�T�XN<�8���,��9f"O�� T/ƪ.AZ𰈖-�V�"O�8ڧ�ќ9�8X�p�ُ���I�"O��"�$ЅSjЍ�V�S!6��=ˤ"O6(��1���㰇��t�^�"O�T�T��?���j%��	h�"OP�rã/vb�{W,P�M���"O�d���6#N�P%j9D��K�"O �[�%�<\e�t#�.ƌ�����"O L�2��J�-�%EJ鰀i�"Oz�`$���&��Ч�I��s"O���kͶ��pa��O�c��P�"OQ6ԃ����֌,�	�"O���稇�^6��{�G�r��L��"OZ��`��wh�mB�P?�"�"O(�H!D�?�L��n�$����"O� � 9g�
4o�5_�=�c"O�l��	B�aq��t(��b"O�T(V̓���Ѝ_6.i�q"O�Đa�|V�Z0��pu"Od=J�%�3�Ԥ��+S<+$� ��"O���2�ʨ�:�B�̟6e7��"OL�3�h��Q���uˆ�~�D�{�"O�m����@�� ���u�8�r5"O��� �S��T�	fq<8s�"O�a Ō(���8���F� �{�"Ov�2b%Ĉ	JL�Z&I�0(_��(�"Od� s� �j�㩄'f\� F"O�MZv��qQ<���{�H��"OtYk&��FM��@�1>x`�) "O�� �̈}H��#���P���y�"O�ɀ��a&�(8��H�&WQ����#�y��̛�?�������DE�<�rM��\��̚�a�&`���Unk�<�T�] 1-| ��F�,M��Ջg�<a⯒�td���'�  ���`�<� ������c�A
[4q�"O���6�.x���c�1�ޅ��"Oh�rB�E��<06�H�z
�yw"O �3A��i�����̪5�:S"O:���8����U��'�"�b�"O$��W�K!^T�¤Rh�*�z�"On !Iܪ=E���!���W"O��a���0w�(t�0�F=20@�D"Ov�Z� E?2�K���P���7"O���#+g����ҿA�TQ�"O� �w��3J�H��l����y��A'L��`�`a՟���� i��y�8a��w/��0J|Ys� �yr� E`vš�-��-��C�E��yr"���pSrm��)��1�Q���y2�X27�>e�����)�|�����y�J�5$c��K@!����B�y"�86�ٳd��+k�F�H����y��C�J䬭I���sjz1�p�U-�yR��D)�F	�T�*qk�Mǯ�y����X@I���Q���w�̷�y�#��H���Æ�S<|gz�wAƑ�y�;0�A�� x��U������y�#��T�������1���H3�y�GJ	,�u9P����+�:�y��\� ��f�]?Ij��� ��yrLБQ*�qɴk�qf�y�ǖ=�y¡?w�x���ey�t&���y"!��6���Y�)�4Y7��i��#�y��ش|ft�ȇ�ר��1����yB˞�oDL1r��D.c@b�Awꞇ�y�-[^F`�"�O� �!�N�<�yB�P�[����G�H�0� ��+�yK�p&d����Kj$�������y" �I������qf�I6DF�y2R�i4t
шM~/(�P�����y�]>:�^(� Ji�X��,�y2�[ :�><"�� c�vL8��;�y�B�;�v-j%LE�G^��͋��y���EzU��ʌx_���$�C��yR�^��D�UbY(s�D���
��y��G�m��
��5t�$y���y�i��<���cc
4\LZy��)G>�y��R����"���
��e �	_��yr@���|��؟3&������y�!����\��I�71iv����5�y�B��
�Dz����퓶�y��,r�nS ��֙x��ս�y�ߑlk(����܆Fy����y"̇ ��W�v�R�Rۛr�C�IJBԐ���=N+ĳ+�P�Kt"O,� �ɖ+>_�4�2>.��	��"O�,�w�
\���#�N�N��"O�$�J�I���W�Ge��{G"O�����S��8�p�O����0"OڔH"�R����PAHW"o<U�"O:��P�̙ZJH�ҧ�"�,u*5"O�!�����ĸ�G�@���	�"O�=��O�1s/� �Ɠ�J�� @q"O�X˥   ��     �  9  �  �+  �6  �@  �K  �V  �_  �i  Ku  \|  Ԃ  i�  ��  ��  :�  |�  ��   �  B�  ��  ��  
�  N�  ��  ��  >�  ��  %�  *�  � � V � ( �/ 16 u< �@  Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�� |d��"O
`�(�;���8���-0��1%"Oj4��ND^[��"3/9�0|H�"OB���H��*�ʞRy=a"O�味V�!X��!&F�:J�$���"O,��a
���C�Ą�M�"O,$3%o�-���p���+Ն�:1"O��ݢ1����`���y14]2��i�<�6��{_���c�H�`�fX�$Kn�<��A̼VI�xR[�)�Ć�pඤ�ȓA5��('nߡ4�� �)˩%� ���,��r�؊b#`T�eT09���ȓ!�b��g��}�8�F��-? �ȓ
K|m�ș�VṔ���2�%�ȓ"R�X�j�4JN�1�˘X�i����̹	_�jZ��1!g��zܶ��ȓgil,*�J�
j�Ne��i�J%b���f	�(U��:���G��$Y^م�~r�� S�%T"���k\�jx�ȓ|4�1�îJb��@ӵ�ݩn�V��/[`�"�v4�R�!ʎ<��M�ȓ`:��z�ؚh�J�Z��$HY:	��H��p�m�C1��!��B:��0��EnjZA V;9����J[
2���	��4'J�EA�IVW&��~�(aZ��ӹ�>� o�Y�|�ȓ�f�A�
Ο7�H��M�$�����mޠP����/���ANXo*�ȓTv�����{ ��-7�*h��I��sB�8�8���3����ȓNe*M�悡;������X�o��!�ȓ'lj�#F�m�+R&;�|��2)n�C��0S4���T:
b���:�0!��e֊��)��ͷV��,�ȓ0�&�8#���� ع�L�����;�P�AFd���,w�6d��r�EQ�( �gVlɦ�M,H��,DP���|�I	$G#\���ȓ"�)���E�B	yt&B�^�LɅ�4�� ��eëF�ڙ��n��R�p�ȓp`@}bŇ�=�$�AUN��P�����xyB�1&0��5������yr+L1�����L�?�H�[ǃ�(O�=�O��<��hçc��xH2,S(�\D��'�X�+UʜP�> @Re��'�Iw�8h�E�R�*�Z#MT�r���"�7<On�J�}"F��^)��5��M8���5+D��yR��[�H�9�//x^u�ċ���=яy2��{T�(^DF8@��U�x��B䉪3�`a;�-��j�́q`MS�U��=��''�����Ț�f��[%FC�8���!n6���H���r���7� ���N�6��E�+��F݈js�}��%����c�Q���=�#Y�Q���4xQ�҄o��=��!��ل�3��l��j�B��]�kW�L����*��� ��O�o/$�rrKү@���Z 8���O�|j��C���=��a���X��!>�6)�䆉(J=dC�I�MT�����"�nh�'�U��B����,w
C�O�Far!���l�O���	
5�Q�ƣ~nd�1���L��䭟� <��Ȅ4f���i�aM3~�ea�"O64�(P,
�jعj�7�^%r�"O舳V@N�n�h� �n�a��<(�"O�т�����,�TG�-U^�xR��	æ%���JdH�4�8�T�+U�hC�I72Ԥt�b��n5�@CK�G�.�F{��9O���ުڈ�SQ��G+���"O
;��ǿШ�ԧ׺w'塢=Ov��D«)�Qb�6mf���џ��Ih�O>��pUB��jZԜ�"�ܟi��C�'y�	�bBX��I���:��'N@�i���X��A����'S24�
�'�pZ�-��Pp`��H�$2�p�<y�n�k܌T��eV���z�Jn�DQK�O�̒o��v��\�b h�e�	�'��Q1E"��*���� B�U/��{A� �S��?IL%Kv`q+w�J����I�<y.U7����֫ƗR�}Pq/�I�<�%A�
~��Ǒ�F1CH�<�FFF?XQXq1��@�)!$q�#j�<9#-Z�X#�㌷W�LɃ��h�<qt#=n����H�0%%��� �e�<	�GڀD)"Ma�`X�]Z���n	a�<)��6�j�SEk�(���a�SV�<96��u<E�@1m���e�k�<y!�1_����i��@T -��aTa�<A���q,�Q�{��	1cS�<	 M���� b��=��=Wj�P�<���S'�,�S���/��PP�<1P�	g� `dD�3�"tP�U�<i�F
;=�
7C��9"SS�<�%.(�H�Z恆�L~�H�r�LN�<�`�<Jȸ���D�ug���vLK�<��ʚ�T�pK@���s�\�<����n�i ���%�~�S���TX�(� ���	�Y�v'��D��NV6\?!��9S�Ē��Ξ3��b`�יL<�z������{��)%h2��(
�3�!�Db�B�C�X�H�&J:�!�&J��Ӓ1FRᩑˆ�0H�}���\[5�ޙG��$���&qr�S��%D���p� N_6�k���&���i�%%D���d��<C��C��{���>D�Lp6�ܯ]$���n�A�F�c3'�-�S�[|JyQ%hŧo��`y�$�*����ȓ17���6�>;L!�r��_^^h�'�B듌�$8ړQ�Y�4����a�fh��S����'��PI��*�X"�Ɋ�>�����)��<�@��<�v���"�7�́�ևA\�<��!��c��8��e�@b@��d�<aP
T��2�� V=z�didJ�v�<�'73����h��?��C�"L�<��Ɩ�{�8�+�bwC�<ӐJ=�!��	G�,ĲQ��	:�|�hKN(a{S��o���M	�+��~l֨K�g�*g��Cqc.�D�<�O>���D׀(Sꝑ2���o����iРZv��ܤ;J����GY��� ��B�}�Xh�'��P9��8f咡g�08��'�z$!s�ğ-~|x�E<x�0!�':��E�HN��|:%o�?�0��˓�(O���R@��;�hKH>%���'趘'�Ċ��5�|��S��@��6��p<�S _?i���ޥ�4�ˠ)�O�'}ў�'u���'ŦQ������4D!��PgO� �����O,W�A5�`�A��'��'װ%yf��)s��LQg�\�����'`n���ø_�`�!2�S�Ѻ�'��'�d>��?��G��0���C��E3�ܡ��):D�T�҆;���Y0��(e���	q̢��zH>g�>��O�BY��1d��A��5Sw��J�')(�A-+�GѺ ��'WV��0�72� ��	��hA��>�O^��u���y vL�@䊓l���*a��y����	"�pܐ�.O�b���'EM��y��N�]ڈ0�B�a4KƯ�.����d?��4��S�Oߔ�y7.�$�X%)Z�W'0�	�'ۂ)V&U�f�x��H%�B���5Oԕ�+�5�V����=o�E"O�dhv�C=xp���,�hj4ٖ"O�EY�Xwj�����<DVf
��'u��<Qf����"Gm�9�!ʷ�C䉵#���g�X �Q���Ճ+�B�	@����Y5U��PE��-�VB�:_Ďh�E��,Q�H��U u�*B�	6}�hu ٽR�؝�����^B�I�O�ա6�W*S��Ċ��;+/�����"�D
49�:ȹ��س1������j~BMD(Q�*�#���2��-@�ǝ��y�"��e�>%�"�K'U\Ψ�5o��y�Պ,&�U��ɟ
SP�DR5'J��y�����8�MP�L;��A	��?	���s�J�ul?3ܺ�(�@�){Ў���'�\�a�Ѱ<eOP$�,	3�'@ar��]�$��t���y���gbF��y�	�oT>y��i�#\t���k)�yReݨOx)r�OPo�^-�V�R��y"d�7¬��肝7'N�j����y"��pMҹ	q-L�_�,0TB
�ybſHX�-2���Ss�Ah�+��y�$(=�+�'�&z��4�2H��yb��?:P+d�O�}�Ԕ�\7�y��	%c1���c�s��T�$�y��;!�̫� Js�0!�f/ת�y��1p�����*o����DC��yB� l<nX0�p�-����y2��C�Ma��_hg(�pm�y�"J�0��<Q�f
gt�12nE��y���t*�L� �P�1.����<�y���&���\�#���C�&4�yr�4�$�R�)����� Γ�y�/��&��M���
��5эS��y�M�=j�:�"6�ң0٘@�ޏ�yr�96@~mX�	�0}jZ`����yR��.N��]3W�U�&�(�bi	�y����U���g�q���s�ά�y�Z�p��9�I�z����@#��y�@';���g�@9C�t���!�y�%�A�\�(����6���@B�>�yRN�p;��	�Rh��UkT��yb@��Dh�@ᘞY6���*
�yr�V1�d� F���������y↑$��FK^�r*��I�n�K�<Y�`�;K�� Xg7�``��JB]�<ٕ�=I��#�A24��]��.�a�<A�=�"بP#�D��0+
V�<A�_o"ĔH�D^�	F����"�F�<i�O	�
������u�@x����w�<Q���4SE;$��9�R�#Ӣ�r�<���ݻf���i���& '�(p!(�I�<� F�J���;���AӇ\J�5ʒ"O����F�/X�ȸ���Uq�8Ԉ"O@(lF�30���l��\��̚�"O D��U!��Ϻ\Z�9{�C���y"BW'%�*=8�ʬF֦���m1�?a���?����?����?	���?���?����Q��H��Y&KlT���T'�?����?����?���?1��?���?	$m� 2h�l@2J�(�����?i���?����?����?	��?����?��A�%o��A�U�b}��p�	=�?���?I��?���?9���?���?�gE
1�����Ԃ#v�,�#���?���?��?q���?��?!��?Y�T�D2���.؋X�V�iB�Y�?���?!��?)��?����?��?�d&�\��
慖�xqo���?���?)��?i��?����?��?	to�.jz$��,�"�$���C5�?Y���?����?���?A���?���?)�)V�QX|�Q$ha�iӊ,� ����?����?����?����?1���?��)-j40r�ʓ�L{ĬK�<�6�y���?��?���?����?����?)��+���$�U�B#��zp�Ͷ�
(x���?���?1��?Q���?����?)��P[���Ŷ�ҕ�a�`�T�y���?!��?!��?Q���?I���?)��p�L�Ȁ�B��� �&�;�\�x��?a��?���?���?3�i���'��u�4ـj��L��������%�<)����󙟘�޴JN��K�T�5ƌ�G&L?� �$L~~e�2��4�4���iӀ89E߈M7t�ya��j� �p�Ӧ��ɦ	�*m�Y~Bo�o�$!rKM�)�t��-bS�[(.59u�ο"�1O��<���	�*�K0 V�QB���Nܨa���m� 
b��r��y�
�+�r�pa㙍�Nģv#�0>Ψ�w�F�IIyJ~��bK��M��'�,�������A
�I>�!���m�������b`��`^B���D�'n�1!FT�	��}�7��mJ�ʝ'c�|�I��Ms��̓3�,�b1��S�P�!\�R�2�BG�<���M�'��Ɇ|z��Q$�1*vPb��s�^�}c��І̀�"��|z�ȍ��u7J�O�sE��v�Iɕ�%MF�����<!/O���s���&�W�n�6��⏆�FT����p���ܴi]���'%<7�/��?�Q��J�u� ���a�W��q�c�O �$~�l��6G�7�"?i��ϪQ�����'�CB�A���"�Bi�d$X�$�كGc�3
�SA��xR�E��a�:r n���!�3��	a�&]�0-�yCưƦxbq!E:&� S��?(��"O�<��$yp�'�̘Z��|:�"J�@���g e�Y0�N�sYm�Q$� 6`�D��A�O�t����	iz��Ӈ�/J���IE�Q	2�Ц��7P%L��4�ա�c��S��5f]8�b�LN�E!b=�'+9 ��vG �{ۦ�G�4or��@D���z$*E 6����`	��M+���?��"����!'X6?
F�C�aĞmM�a���d�OXб���O�e���$�O8�	)�ԧ��+0�0qF���#
��M�!�H��?�������ʓ���J�R��$�'X|t(����;�*�l�%��8X�4�)�'�?�D�O�-|]x"BT6���c�w(���'J��'gr1���'�T>�	{?!��Q>�舑� p�h�C�m�1O A��K��|�������F	�z���I����D&���M��-Z��J(O���O:��|B�'C�����c[��ٱ�D�2��f�t��� Qb~��'�R�'OB�'b����d��tw00�A�) E(k@m[b�'���'���|��'���ۙ.�H�♈)�������U���V�����O��d�OB���O����O�ق`�\5 �,�
r�� ԰;�b�O��d�O�D/�D�O��W�%y��i���C6&z	����bA�Zj}r�'���'�B�'��GX>E��N�����l�T�el߆�n '�p�I�SQ��%UBrO����S;P��߉����Ѳib�'��ɑ5��u�N|�����$`�M)�皭XD�ŠR�I�l�4�o�uyb�'ObBͥ��0��iZ|Q���:
�,ZpkJ84k�zӼ�zM�uq��iʨ�'�?�'ch�ɽSUP ��ݔR�F�!&3�7��O��ʿ����|B���&��D��j%zhP�O�*�܌ bny�|�R�M�Ϧ������?)�I<ͧ��9�t��{ꐘ�$�R�y
p�i7���c_�p����d�3�ҟ��SC�W��`G�*2f	S7��MK��?��[�V�QՕx�O���'�^�CG,�-Ҁ(�Uh�$ir�V��>����?�Q	�a��?����?)��BlE�����X�D@�(��?)���' |��e9�4���D�O�˓lE��@�H#U�l����	u�Aᖰi�҉ֳ�'���'�"�'��G�R�I2�LϣxUB	��v�μ;�
|Ӛ�d�O:���Ot��O\������0������"�����Y�$��AR2�0?����?���?Y/���WOҦ�ۖB`߀5"�a`k��@�d��f��d�O����O��$�<��$p��'~�Xc�������8�m!0�8�S���������џ4��2n��޴�?q��b����ՁRM3~�U���LԢ��i���'��_�x�ɹv�$�S��T�Iq.|����\;���u�@��l1�-� �IΟ��I(F��$�޴�?���?���X�l�@�.}Pȗȇ0<&$Q��iRP���	����S�������t�? ��{p���Mu�@`��	*隂�i��'A��Kob�"���O$�����	�O���U��
<��Ze�شd�$t %�W}��'"���7�'�ɧ�4�~z�h�6H��#h�0_����r�ϦyYr. �MK��?�����'�?��?Y��y�J\��cZ,�j��BJO�&�fa'��'X".ۗ��d��D�O�u�q�6>��h���O1X,���b�D���O����!m�2Yl�� ����4�I��]#=����NR>�	�D#F�V� b����1�I��	���Y�ժ-��	[�Z �8X{�4�?��:���' r�'~��~��'ׄ�{��@u�eA"~��O��5<O����O����O��d�|"���q��Db⨏�EfX��/��Z�(ذ�iM��'{B�'��'���O�uQǋ��Eܦ���Iԙ\�9�G�>��D�<i��2�?9���?�P`�{��i5,��1�W�D���ZB"tFn��Ž�pT����T��՟t��ZyB�������4+�:�+P�3��ݫ�	��x�n��D�����Iϟx�	�vM�ߴ�?��K�d�!w �z���p0�L`��}�!�i�R�'�S��ɉ;���Ο���\�@�"цB��Q���͟tj�eo�؟x�����$�!;ش�?���?��'���si��b��+G�6J�-r��it�S�t��	L��Ο�����4�* !��7F<lAҴ'�$	��dnş��ɖ �갋�4�?���?y�'���u��j�n�q�,�a��+պ\P^���I��FX�	A�i>Y���쓠�Ą��!:À+c��zq�i�vM���u�����ON�d���I�Op���OT�`&-I�uI̉��;!#��h��C�����D���	���0�e>$?��Ӛ2pA	� �IX��ғ�5���4�?���?�J�]���'�R�'���u��=e�8����$3�2��E�I��M������Nc�?���˟��I=e4���6��/����NZ2pJ��4�?��˰_���'R�'���~�'�L��y	�T��F٩�c}��V"�yrZ�������D�Io2���NT�f0��ɀ	�!K,��˃��M��?a���?q�]?��'���,����DΒ�j� 8�%�N7t�'���'��'�'���'��H�}�6M9(C�S�L�%+�)(��o��`��џ$�	��'F�%Ԏ��T` 
��Y-Ԏ+tKĬ�`� ��l���O����O���O&X���KȦu�I����ǔ4.�����F�j�/�M���?	����d�OHq�D0�v�䷟lH���=.�XhL��
��TIp���D�O���O�4as�Z������L���?�0�
=��x�&X[�Ɛr6&��M������O(���7�����<��e��!R��pcq��hd�yj�	n��i�����oȖ7M�O,�D�O��	柶�\�@��йT�R�eL�}1O��3���'��� �Ek�'^�i>����=Ad��oȐ��D
1
��ܨYN����
Μ�M;��?����Z�'�?Q��?�e�בYF�8ڸdL^\(Ճ�!ZЛ^@  "�'�rZ��h�S��3�lV�JPx,�(�S
(�{�ڕ�M����?�+~�y{�iR�'
r�'�Zw/d�A���N���dտG�����4�?y+OV	��;O�S����֟�Q.ڹ�pr�\+]/��C��5�M#��Bi`����xb�'�R�|Zc�lը�,L�n\p��Ͽ.Ѐ�'+�%� �'��	̟$�Iq�S4I�T�0�iƪu�^�h'��~��=s������?q��䓨?y�[�&�)���'03Dh�"/ޯ}������?9+O��D�O�Ĭ<��I��n���6\�@撺]�t�P�L@�w��I��h��f�	��l����.'���P'^<R��T���J�]��쉬O���O��D�<�0X�^��O14��s�� }��J�E�N:h{��p���$7�d�O��D§Xh�$'}R��� F���fF� ��P.��M+���?I+O�u����@�SΟ(�ӥ �]+����d~4y�����i�I<����?�D���<!L>�OF��@ ��kfЛ�>⼴;ܴ���.�\lھ����O"��A~���2$Jd�Ѐz&B��Mk��?i�n��?I>�~�!�Nt�A�w��� X���UĦU��F��M����?A�����x��'pjXj�}���En�wE`��q�sӖc11O̓O>I���=L�%Q�� :X�0���բv�Hm�4�?	���?y�����'��'3���rxh$vlK�tޢ|���V�6s�6�|��l����$�O����	J�ze�'p����--f5ڌm�ȟ��uɟ���?Q����[���-�(����sQ�bG�K}���hW�X���	���cy�ew�M�IV�:��lb@)_#�*�(9�d�O���3�D�O����1�j\�u�N�]��)�gF�G
� 0 ��O�ʓ�?���?�+O��G ��|�b�[_h8*NPP˖p���{}2�'���|"�'��e�9&��IaG��S��B^�R'\k����?��?�-OT,�Bk�-����a�-c ��D+T�5���ڴ�?�J>!��?I6j��<�N�\Ss%�?p �����&%� `v�d�����O�Z|@��%��d�'@�t$�)tp�T��o��^���ڐ�HP�fOV��O~ Ȓ=O��O�ӻ$�x3U(:�#�"H36��<I�-��xB�&�~����J��,s�F�V\��d�Ulv�F`�����O
�0���O֒O����ŀ�v���J�}R>uC��i�����r��D�O����(\&���	-P�"%eA/�qa`�N�^x�+�4m���̓��S�O������;� ۔�S�dp���UIY��(�G�7v��3��H$[����0l��hML��9]4(���T�&��(��N/v�����;/,�ӀmMz�q�U�'Wh�w(��rr�pc��	sJu��jÙ%�b=�g�2g�)�X:�9�tb˝k��4S��9�<�Ҩ�C3��ٕ�B(% Q)Q
U->���MYq��I����xm���.$������M�~�t���	Ңc�1��o\ Y�� ��6��}1K�PO�}��N�N�6������|����ɢh��U�I埘�'m��ٮ#�������<�h�Ij�=�@Q��.���� �J���O�H�@CխOst�����aCf�5iJ��C��el4I����T&�7m�p P3��$
9�bs�|#bR�O�F�JB&ZgO@���"Oy�T�F���k��B!a�Ȼ�"O*��BV8t��H�V�$�Dh�7O�xlP�L��a��4�?�����II$ˈ��sQ2v��i�em[�/l����O���O�I��F�m�BM�2��/A��`&JUn��'5�\�"C��|Hт�7�(O~�´!.����DJ��p���~a�ϽY��W#��(yL�
�ɑC�'�9 ��h�2ʄ��>@9P�$�+;��Ȅ"OL���������у�&d��'fO�9����fW0��B�2Q�b�	�9O8d��æ�����4�O.R(A1�'!��'Z\]�FM#��AӇ�@d� �y���S��x0�<Y��4	5�N#%��'ǘϿې�7��2�H:X xv�	���3P�]�t�ʄ�ʪVМt�s�����6�U�"6������mK t	T�m��$�O��S��w�I3�-"�. )��we�U=�B�	�Q$ޡ�!&շ~=�x�BK�0an#<���)B�J��a��
ՏA�Q	��j	�?��^��iQ���?����?a�[�N�O��D�*5�L������4���d�4�	�[1!Y��@�Q�Ѝ(eџў\��fI.W���ÁN5L�1�X>�?邃�98�p��W�8)�^�3ړ"Z�: $�jm�q�#�ח �,���"��E�	���=�#̓������
�^�\ͩ0�_Q�<�P�:o��L�~��ѧ�_5uJ��"|"���6 ��F�ؓD�H�	�(c� rR	�I��'�2�'irQ���'3r;�,�� �[`D�I��I#?�2�hV�'�,��a)C-KD^���i<<O�	�"/C6[+�x����9���vK�"D�+J8\���РG�^��@(�&���`Lj�{bM_��?YS�i�e�P�:�8��1FJ�Z�@�(�'�E�ԭ��b���4$^>a���2�'��t�glǲ#6PAį�#�(�J�'9�7� �˼s�\o�ßd�Ih�t���ҹ2�m�71p����O�;�`�'��'v��%#�"-3K*?��T>�XFC
r�1�b"�)Tϔ��!�N�(Y&�J�ȡ�b@ֵf�\@�W��A /\!\��]�Wk��r	fAbd�M�'E�L���P��>=:#F[��,�(�<[j`H�k2D��Bg���b��؈h"���͌E���N<1թyV��i� �2 B����<!B�ѐ*	�v�'�X>���K�ß�����Cҡ�2t�`,��F�%���Ж�9r�Ҵo�8	l�Y��Ɩ^��Ij1�ӯ@��(�|��(X.�80m».��U�E

�W5��"�̗:���lS�_�rX@VCǨle�d3��;��Ͽ���A�B�Q�%x"�����:�x�1�Y�&
�<��e��?Q�)2@b� Tm�5/�f`@���<����>d"Õpd��cH�0�l��l�H�'Mh"=q���?����hq"8��a��2�c�c_;�?��P|ʀy����?���?���	����O��ċ�^�J��4�C�=���3�P&(�`d�k��O~��E�	��e�ݟ����'K��'�zUYE �
��T�a(�+g��GI[g|��1�C�2�6G@���t��xx�q�o�h~R�Y����
�$&$�(��@>�~�Ն�?��,�f|Y�aޤ���О<���ȓOْ�2� P�V�|���#ݟ��Ec�i>�%��2���!�M�T,��f���D�|&�A����?Y���?A�Z�=����?��OS�(��4P��%Î-hu�W)|Ș���	:�p>���˦�j�|[D��ń(4����&�%�����I�@����֦�#��X,�pŅ�,eNH1�'D����Ō�GN��a��@�eF�+�.&D�TX�Y�{rT�qa��;��}{�Ff�hAش��T�p���iqb�'��S>@���"��X��9MW�F�NԪ�������ɟdPfiI�Z˺i���@�X�6��|zf�p�v%�ƛ�l���YB�'yD�Ye��X���:��Vn�'#(�1(0�̋ ��u2W�8�:Dy�,��?�����BL�bh�^�.����J��!�!.A8@��B�5Z��0���@�a|i&��Yb��X-T.Xj� ��2����)�r1m���	l�ԅШ.���'�R����L��ϑ9��m��$� #�4���'�1O�3$z@��vҸ�Z��c�<�K�j��O?�� ��� #�7s���RɈ%)��4K�-J�2��dm�)�� �0ő#�����PN�z�X�,:D�X!�j�1C왚���D�0��À5����'^׀p���Bjڍ�+W�l�l8R���?a�����r�����?��?)����4�,U[�SB^�[�`_:<`�&��d8BٹuB<�@�
1W���ɧv���	�=0�����>n�J�Z�!�$~��-�E�tY��h�?=ʷ+G�(a�x▜���,Nv�2Yp��V��ԊٟThG+S˟p��ޟ��<����$����,�C�Dظ��A	��S'!�P9�Ҩ�I�2�z�A���%1�HGzB�Oh�R�t�5�'�MkUJ�
9@v�P���3gG���G��?q���?�����9��?y�O qxӮB�d�T��%��4�PaX��0ѮU9g�C"b2�;��X�%��#?��+� t��r�L16�T�c䍖�2�(Q'E��`��O�v��y�b,Ӕ�yҫ��������� Z�o� U�T��S�S|\��P'#D�p��
�R��w�S�^�B<q�+D�)�,��!�9(�G�^����`�s�T�ݴ��}�LԻi��'�ӸH@�ճÍ̞}	x�҄հO��|������I؟Læ��,њA��O�Ke8��1�ٴx��ɘ�<��5YP�T�@H�����(@Q����B������/w,L��4fq���a��%�>4���!l�R̂B�Q�3�P�á����0�P��	��H��A��JJ.ԠaphԿ��lA�"O�,�ǁj�L,����c��"��'�NO2��T�Ď/9��16�P��N�=O@}��!�٦9�	ǟ��O�^���'-��'�h ��N�cf.� ��>K��RCnΫFo�9&`Re�X�W*�O��Y��P&DǟL�vx�����$ɛ�C-�l�DjC2-��sBL�%YW��]w�AC�b�����*��j�y�J1Ѕ���;m��@���L���WC�)��$�g���h��e�g̿#��C�!��dʡ�ı_ݬ�`w�N�#<7�i>�I,�@P�� ��+�)��C�
-�I��Ps'e��eX����	�H#^w�w��h�c ��1x�(P�O���q� ���oR)x�A�41�X���>��t�-ʓT3@��ƛ\��Yul�e|.iI�%X#b)��eO�'r����OJ� 7{����#��drPap�*P�Z��֯R1�䃂~���'� �S-K8fT R�A`/<Ar
�'�B�Y�Z�ț7S�a�FjT�i��#=�'��)5�b�i��q�Eߍ>f��P��`����'aB�'u��ّb���'�		VmR�'o�a`PN�+��u��l)l�\с�f�h�'�����!�>�ơ	ק��4S�H�6�\��/�M���	9�ޕ�F��;gnt�P2�O`�<��&�P7+ɬl(�u �)�Q�<1iˡw�
����?A��z��Q�<�P�iw�'���w�h���D�O�ʧGڰ�&�A�w�NQ1U�L�~)���HR��?)��?i�֔�?��y*�be�d��?V�^���.4i�4�	�w����Eڬj�>���jO;��MSi�'�<�"��h��p�O޽IkrQf����h��"O�dEĝ�X\1���$!�<��2�'��O Ha@![�=疥���J���%��>O�I�����y�	����O7@�s��'��'/�]c��L����� �|���.ul1:!� �*�8C�.�;VV�bR�ۣ4M1�'5[)�xٕ��Vl�D�zb����ď�MF��(BOɍ~.������?�x����g�L����������f�ǝE�h{�KĚ�?���|���'��w���|��	;�T��'����6q:�B�O-7��H���Ln�����'�zt�'��=���ɑς45[�j1�'��a����x��'�"�'��b�E�i�i�Q�+7FM)�jF��V-مk������&�O| ����:| 	T �6^�>���O�i���'�D%#Fd�� 
(1��oP)��P�'l�p����=�2��=}��R��?	�f�S�V�<!��Fۀ�9�SwH��&ɻ�Sc�	 �q�شj�!�{"!V�/z�����?	��?A�-ι�?�����$B46�>���T�t3��у�0_p�b�K�aM`��@$9X���#L�fDy��˛SM�����5e��QlS�_��1���&!�h�@�,��K��TBR���Fzܓ*���I��:ʊ.!M|d���l�Ỡ� D���U^B��� �$�^��#+D�\���U R/.0����dDy�Q*h���ڴ��M��3��i���'M�Sg[�)p�+��>��a��+S�,V�;@J[���	��3�H����A��\�װջ%_���I��lܬX��E52�+T�m��ԃ��&N6���ޅ�p!�G�]����^뇫J3x����%k���[�BI-N�L➰h�$�O��}� �Lu�]�%��H��R4{���T"O�����q#��J��
�'�.O�@���lHa�����n���g9Oڑ���W֦}��ٟx�OX"�P��'V�'���#%�i�V)�#k�)J��
D�V'di�g���פ(�L�v�<U���Ͽ䱵�|�#s�Â4���q�@Y��{�ڷ!~aЎ� >�(�!%7��i"Bc�����#fE�9t����ܭ]_�����;`V<��Dy�)��$IT΀�%:H�u@��q�ޝ�E&D��� Ki���p��(j�ޡ���6�	�\��4�T�dU��`ӣ�V���e��2u����O�u!�m�'\�,���O,�$�O��;�?�;Ix��mP��D�z� ��MPJ��B͏.��҄,7cm�	��#��|�RI=�8�,�4�ȡ<2,)�d�G�����+ߌ{H`:C�X�h,���DH�b�C�� ���������$��$MpMHT�Ԕ[ɚ��c&�3<�D¢z�ҥf�N�'�X�	ԟ<�'�����Q,$��Kڥ'�I��O��=��R.O�$�A���.������9\66m�y���M������'���D5�$l����܋�!�*�t�sJ��Q����	���Iß�I�x>����|⁌�T�n+b��('����2'��#R[X(���6[F ,�L�.|e�N��A����K�wv̤��q>�)�I��M[��D�4����dl����Z����'9���t�?�OS�E�g��7�8qC�)hN&�2�'Yhq5 S0�^D���¼t�T'��L�����b�֝�;�?�����D6���0�'Zx�Ъ��)B�AW��O��D�OJ�����a�RDY��E?l�L��|�3"A&T��Q�%+�]�*�r5̂M�'��h�0�8D�>��&�FM��lsK�P�[$h�$M�J�)�=7�@�3jZ����=!u-����`����M��tC�H��ZR$��
�(m!��/��jacZ_��5�̔	va|�A6�
�/�������0��3!*��Ě�5>�l���	A��ϝ�x���'0b�^X�)�S�*B$8-●��bi���:�"#�߹J���T>Q�|�Ʉ8l�E[��ð7L�4[�)��T�tL�1�Q�U���Q"���I�v���¦��->�ϿTW�����b @�q#$#�@rxeX�-ɧ����O	�Bic�_�4���{v*N��yB�������K�*T`�V���O��Gz�O!��T;[h(B��ŝ,��5�������'V��r�A�i��';b�'�����$u�$e�R�/u���T#�,<*&Az���0
8�$P�q�u{�¾?=h��$�2t	�T���j���]�
�����T�>a�D���Ų�,����d�W=Z~�Y���_��Ɉg�0e����Y��]R���h��I�n�8�ɒ�M�Բ��,O��d�<a�k\?Ag̔�WA7O�d����l<!�'�-�Bđ�5?��i��G�%L��3�I(��l��~y���C�:�ݿ2p`$�� ]���a!�I?nh�������ٟ�piO�� �I�|Z�(D�
��l �+	�|C�96�$`�(��#�4��K���<Y���#s���Ъm��P���Z�`t�Ы��L��	�%n�?M"�hH9� DDxR���?QF�i;4���hO�E��{1C�p5I�'�:����w�pz�,�l%���'���G�\�	� ��?[�X�@�';06!�D۲,�\dl����Io�t��xz��a ^�[��x5茌��q��'��'�@t���٣N�)�R:U8�T>��$�&3�)xc���}�,5x$�?�d= eD��6`t�Q�G�9I���yd�ߣyM��ق���`fT��
�B�8�o�J�㞀�7o�O�G�� ��L�ޡ�EY�4�Ah���y��Ú3�hl�n�OEB ������0>��x��3	����&��
CF aٕ�ű�y"�݌SJ�6��O����|rիڠ�?���?1���M�N4s!!�7or�n�K��X��N('f���� 
�`�*�^b>��ë:� �K�O�2�d�P��;Q1<��P�^�l��Q0-ƿ�Z($D��� 
�IѴ�X��Ͽ������'BM��<[P2",�|�� �Ovb�"~�	���M�5��/:%�E���V:~C�I�]�>lС뎦s�tM�f�T�E�"<qB�i>��ɱ1A`t)U��S����O���Iٟ����:\��p�I�����X�[wW�w��9�����%��l� X��|8+/�x�d:��M�qcNu�cK�����鉸F�L()�\:Z=.F�	<4�bg�H��;6�اc��E��e�?�oZ#ZSn�3E2?!4k����Xŀ�,>�q�G�Ak?1&��럠��I3���G�Ýu�QBqBW�<%NC��������=$�l�����T� ���4�J�O����æ5����2Mcp�� ��������L�I��z,�	㟬ϧ7��h��Ϻ�l��6�ӻ>��ƣ_?"_�4b��[x���l����O.Р��  ��}���U내��֚v�N�A1)I�O;RYd
� ,0�7��5[Ρ���J�-�"�'+J�23&�ga:�wm�o-���!�|B�'+b��?� "<��n�3s9&j��	-m��D��"O�A*�(�XqR��&�X�1�^J�5OLnʟܗ'������~�����iD�v�3�F�U�J�0e�C�5Q~�J���O>���O�B0��2(�,2��^�g�$lQ���f�td�� �
@��DDd���0�(O�ҁ➸0���1F�
T3�9��u��@�H�n�.@`�,�!m�<EK�.W@���,�I�!U�PӦY؎��l'�6��%IM�C�*镨���y��'��}��W:p�D��∘jL
I�E���0>���x�Ku}jE!�MW�[}�R��	�y�GI3N�T7��O*��|:!ƈ,�?���?W�Et@dçN�U_��z$�TyB���C�I>K��6#R#as���wW?��|��>�|��k�#�*Tj>`��a��k�ր�dY�t���%
��u׆�/�>Q�O?���Q�Y���˪w���*�6{��e�Oc�"~���d:���O��g-���&�0`6�C�ɪ1i�-xҥ�	�ti���##�#<���i>��ɕ�d���B#ъA ��X"e�v��I��*٢p�5��֟����(Yw��w�����(�hl0�C]0�<��h�.�������3k��`�×����I�t�ȸ��՟^�=��%?���C���C�����֪y>��ӊ�?�o�(*�}�=?!%bܢ��X�TK�� �$p4ɞ~?	TĂşīߴ8��'��'!� [�H�:c�*6@�����$s��C䉛){�c�h�u^�y�U3S�Eb��������<��ع<R�V��Fƀ[�	�t��O�>[��'���' F���'k�;��Ȼ@fęI�`H��Q�r1�RR+©c��/Q ��Ө�/��y���
 �DR�> 6$����	|�z��Ɔ"w&�+c�D6��A����>�n��a!\c�L3���I��M�B��
Ew6����P�-���\�<���=�`|Ac���z��0k[n�\E{���>>t(�F	�)t��nW��y�x�*�O�3u�q���'��Bd6��CC�5J%��Q���$��(�B����l�	Ɵ��`-B�z�@�ĭzVa��战����0	>�IC�$�.W��a�`�	\�Q���-�+?D�B��Ѷn�|�fպ#KB�5�B�	Taӓu��sa������j�Dܓ~Knx�I�M�P�	K�^r�{Q�K{����팁;T���O���X?�n�  j��3~z0�	Ca|�/�K/�P����T�t�AG��$�d�|%m���(��Y��%��b�'8R)�Tl����7S�` ��-I��� � �o4���!�B`�Wh�~ڊ���~5:-�kr_D�Z��L��,�'Gޙ�:qX�C�<�A��n��~G����yO ��f�~���HԺ��H y�i��)�&l�N؀��@쟼�<E��~̂��Dα�x z� �����ȓ���� �(F��2�#����Gx"%��|��N;B(�%�<[�(�x!n��[�J����?ag*R�ɖ!����?���?�1^?�:?�
�/a��5Y���C��� �R�uTm;�I^
v[��&�?�����s�Gՠ P�����J%QE� ��*P��PÁ�=^�*ҟP�����(.�=�!!�>٧��u��|����|6>ps�M(�?q7�˷�?)��?�gy��'��ɔM�d<#TN��"WX��ƍ��C��֟��)O�T ����&o�`,;���HO���Or�t�$E{�ir]�����(�\yƔJ �3�'�b�'Ab+� ;x��'f���8Ҳ��b��j�H���}M�A	�Ǉ�9Yj�`ř{ܐ�{D╏������8u�k�ɑR��� )ԐC�T8�0�I� e��ذ���x&b�"�6�2��-ʓ�ބ��՟����2�88�0
ær����
?D��a���-Y��	x`d��Qz�$�G>D��P���9�cS��4O��pr�@��4��Ajh@D_�����ĠD�M���S�#�uٖe�FJąJ���'7��'����gM	g�&rvc_�N�J�!խI�Jd̨�w��4�� �6;+�R5]�(OT-�e;�l�3�`�+ N,(���mS��:��N]I%�V,�*b_�;5/�(O���1�'�7m���m��{�4#��3"�YP���]x��(�O!��s�8��>�Qci��>����g=�Ob&��jf��)�X���,)�X[ы{�\3r$L��M����?�,�̵b��OD���Oh�p�
��Fer���M=�x�W�ě'Lb��iX;��9���@,�M�O�1�R���r����f�$���W�m%�� �/��B��H�LF&���؎��'�H��T�DF �p`�����Ň_ �
�B�F�<�|��?i�Ԗ<f�P(��@�WeC�<	���>Q�� 
�Z�@"M�u>��˃DN�'�n#=ͧ�?	�C�C���r���s�,�[�c��?!��2��`�'M=�?����?��x��.�O:�DПe��9�� ,�D��T�u�A�U�V9/��@��m͍:��Y+4ҟ#=YaHҞ5���҄�U�m�ڂj�=��=P - 4ȂU#�`4���'�HOX�%C�6}��(rEKS B�B�	a�O���f�'V�{2��&vJ �	ԥ:e�ڦA޳�y
� �
��oEjM�@��h�@�)T%W_���t�|���!9^7-Q�`�����!1�<�!	ȡfQ �d�Ol�D�Ox9�Ae�O2��j>!��� 0T���/��1X�m�:+��M[ �D�>>�h#��ư<�D�]�|]����V,'����ʚ�c��(����v�fPs��
	�|�;�kC�hO2���'��6m�e9���!�/c� �)�,1!򤛇[�^���Y-7ެt���V #!�d*;�N���
&��I�\�N���&�1������OB�'MJp�tL�n�����.�?�^@0t����?����?q���zS
$�
4h�di4h����S�nz����p�|5s D��<���֥TZe��	�K�<u
&�N5DV�K%!J�eH�M�^e�HB��	����
����̟4����<�O�����*��r�6Q1��@茡1��'��O?�I $�\}��ʙKe��R��b�
��d�i�	�L�lZ0�P+Ap����R=y��I
M���4�?����iD8�z�D�Oh���R�AIf��4��@��ʹq�:]`��RFDyI����f�F8�\M*�Ss���M)�n^9|��1����v*��Y���)���*�|�Y�%!Zr�X���w�.1H���<�̍�S��-JvS�
҃<��|�Z}���'�*O
��5'G�u[̊���MFfi��"OR3�#�Q�LJ���SL���ቪ�HO��oʟ��r,˭*
e�	��.'8a��������$f� �qBџ�������+�u��'��͞�̤sW!Ы6ƀc��,�~R�ӣ9�	�3��?����ĝ�fhH�T��%Vm�i�4�1��$�8Z
�1�KG�>�(��ɯK��d�!<N.����@����I$@�,��'�M)O���O$���O��[���"�	Xo f��Bl��Y�!�$�?=H6�p��(PT4i�0L�$�Dz��>a,O�|y�����a���Ѐ��j.�*����a�՟������	g��m��ɟ�ϧ*�,%얈�M��n�Y��'����ݘ\���D�,F�=�4jqӆA�����p�T|c֩պ8.>��B�'��x���?��ߑ/�8p�eB�_�@X�f�?����$�O���'a��)���$ p��Яɀx��p�ȓrP�Ǩ;E��r�Ѓ��Eϓs��Jyb�48�6-�O��$�|�⧝�S�Fl��i� ��;d.��S�$l`��?	��K�����֘���� 6�q �X �.%��]dQ�H9�@7�')|(`fN�d��qHL	:�)EyBo��?r��&,�P q�B�b%2��WP�zB�c����Ac�:|a�98"�R P���$n� (�r! w14�v��e���g���	8�lp���H�	r�B��r�'��,�j�pL�_�� QT�ϪO�J���� C�²V�|�O1��yB�%u�քP�h�c�i�j�)L$�����u��E!b 2�J�R'�=O�<�~��F��JÚn`�+�G����Pjq��ݟ���4I��6�'�?����@��[`��Z���Ѷ�J�zT���O��d8�S�'E��m!�mZ�h�KX9��̢U�'�&���MyӜ�O<�*�c���Bu�6�
'��^��B24��	��� �^��#��qc�L�g�%D�䣳��, X`9�`f�j!v�>D�@YSBYs z��@��$��x�� ;D�|�G��2�"i�R��Fg�\�66D���D�3�����׷e�\�
0D�����&����TI�)�<Hӣe,D��as�J�M�T`kgJ�l��Mb�F,D��`�V�OE�|p��,��}�S`+D�̰Q�Q4"9*�N�w"�ō>D� �똸&rA�.A�^)��=D�XR�	�*��K��6�P(x�=D���e߽lO��볬�";�D��f�:D���b�56_�%��-��<�&ث �8D�t�!);�j�§�Z�WB! 1.;D��@�
z�
�	�sjId�7D�H倠Q&r$Q��F�0FZ]Y%*D�p��R��`ˀ?�Da�6A(D�ԫ�)&I��$�Q��,��
��!D���o� ��qf��A�P���)D����ث�l�b/^��8D�+D��y��̀4�RGE�W���Y��5D��7��.\��I��3F�܁��2D�� ��in�=`�̄��
�6:jn	jb"O6!YC�^s��ITjߌkQ�M��"O`�S�_��p��fʤ+R����"Oz�B��F�p):��H2ZjJ-B "O��k���.n�*5ᗨW�/[�(r�"O�}����X����`Z�;�"O��Y�� /�%h��9PD��d"O����f�xI�Eܙ��f"O���ڨ.��1�2d���a"O��{cCD�9X}{e#�Tz����>���V�i(�]�7�iy�7-�|}J~Rf�4�Hj�m?�`9�HJh�<!Ra�� �H���K�K�Ib�����T�{�,ݲ�'�8c>Y(�LH����2a�d̩�όUBD����*T�!��!=�!�K�E��%hu�B�8��(g�i�|(ⱠB�D-nT�w
W[e�z���޾l����*α=�����Ꙣ��x���xG��Bn�'
�'ˠP��D�P�pe�X�&�%b�%�!a<a�
83�lI2E�vpm�&kL@�	�vm��EǺDLP@cn�	�����&yӵ&a>-a�E	�D1ĭx�ş�A�,"��14���
T�0�jT���ƶ�,�k�/�P���V��nm�0O�1�Uiⓥ<m��~�&��f��;)��x�)��6�h��=�0O��i2!֦��*��M�׎M?�"@I�$0�3j@� �8��IS��)�W�$f�Fjh�b�8h�"M0�_\6MN������n�tjd�n��BA��K�*��~�,Ù'>�'#���(CGP�=/��s�"ч	� �
ҪE�r�����!R�����Y؀�%��?`���?�Mָ'����.�a�������[%�l��#Ee�#U��HX�h��
ʁ9B�@#Q>�8��.�;(��ɇ~��f�� �(O�p�&�+{�(����<>���b��>q��J��QsE�+���.�o�䚘I�Z��L�.��q�H|��O�A�'ӨL+(h�c�0:��Y���i#�e�a%�L�B��T၎��
,/�(]@�!J�e���0W�ن\
������%T��Z��'�<���!V=7��4)�.!1��x��Ӟ/��}�wo&�A��[�WhzH��` ѐ�6��u���w��ñ��w��T�3ˊ�2��z�TP8� �VI�kN�� ��I8�p-9@DS��&��� =b�hܛ$a�	��:ei��6��L�E�0:D�к3A2?�H��[m̬؃��).��!�f��\U�GD��nZ;s��!�=Q7�S�g��0��<����#08$z"A�9��!cċ��ky�1 �g�ݪ�؞���Y�(�>�HIq������[� ʹ5a{�U����kէK�7���-�\�Zd����B�V2aN�s7-�:W��1�+TH�����!BU�u�\���cClI�ih�L�f'��,|��dY�)�M�b/��B�|��\<3�ْ�oXu�� ĺ_ud���$Ԛ�d�5��mi���E79��cu�� �.-�	+B�#%�^�'�)F�eD^�9R�.Pn�����O랟���Ŏ(ag�@$Gc�����+I��Y��B16�Ep0N]>qK�x�]�>됌�cA�3�ƭ�v�\�v�4�ٸy�49eb̪��?�sB���G�L�50���A�6�9#�Z<I�}�x�Y6/p���u�\8��it
�8����i$)��@�m�;�(�)�h�az2O��5�� �o6K �J���2I8Z�@Z�sl���H<�HO��ICK�\-J!�%˯y6J�	W\���%�I')o��K�s}v��Ў,�	63�v��Ԇu���ܦ��<��F'nb
)P"K0����jM��I��E\E�B��eV?\Z��=�I]�(8���v�
��6Ĉ\�d��Ѝ��3�h���,�@�Fz�>��W�p���0��<6B`���Klp��y�"�	5%�d�,��$ �8�i��$�~���O��ˍ����L�$8�"�NT)6��Td�y���Q��&~C0�p�ϲsZ�g���T|���#;�\��U�����>����;0f������P:���U}��ݍ*@�c+M�?���!��HO��[��֣G��ճ�.տ"���V��{��7�x�BF/8���(z��]��/H��A�UPDY��I���ɚ��FBδ+�� 
!k��䈌	���b �\�"����\�A��F{B�V?��9� �+x� ��R�]�4h�&.�O�M���4h]�@sцȽ5� c$�$/pM��-T���	�@���ݼEV^�8���1�ҥj�E�V����$�*f-" ����@?6��d�"{~T�V�m^��`��$[@}��&�F�ؾ_��F�-�^ �����&lQ�/�Vՙ0��!�0$Fz�)�+6n|i� շ+�M���0�M�������&���3o�'Ę�g��O~|bN<9ǈ�`��>�j��&���+'�, /�d�r���MQ���>e�Ճ��,�.���M��?�S�\� ^u8$�E�.� !P��>TX��E��X���'`,)(0��P�&�q��ΆN�*x΂�BJ�dr�l��� ��L>aVY���o8J,�v@ĕl7 �J0�:�O �l���?���V�]����#1*=�������h֫ہ��'x>�q<�<���3O�l�[� ��r�-�K]�zy['6ړ�~r�A �p����^=�R7��P��,�.w(��'a��{L"�p�R�P�q�B̈O�S�G�j,
��V��(s�:q�i�*��I!tP�0a�CN#b�O���A	ER�Lh­Ĥ;��,a�KI�V��R �ۤ�p?q"�!k��� �N�"��C@�gr,�B�i�EzZw�8��@K!I��N�~lPJN�?ݎ��S7a}���L�,ɘ��߀]̪��i[$i�Ȑ��O*Mbb�����b���
�o�D���|��Q�R����"�x�F�*C;�^�@�E3�n��zc#x�����/Z!nz�7-��qb�(�A�tc����3�	�K�Ќ;'d*O`�ge�8x
n�<!#k]:=������M*5jd�Cߦ�Iè�{?4�²�R�Lx�GNf���I 2��h:�`����QCnUpF& ����s���a9|O�X�3�K���9�׮��~��E��xC�~�;o�b�e���%��(ۆ�FU�ϓe�(ق���G!F ��fc](~Y�p� WG0��޴��D`�$�[kB��Ǝs�rdrtë+,�Ҍ�v��@%�xy�R���9G`�&���m��(�wƊ&�P�-��v��Z�	�v�FEۗm������@�e��jZ�m���O",�d��$�h#=�eL�c��2Ղ��I�L��CG��ƕ8�C��H����5,@�K��1���B	������I3^@����,���R�HMFHc`a�|zr�p#
�} �K��<�}/B�Q}���� =��a/޵J� m1
ӓH�ై�J� ��O�Jt����
�?�*Eڀ�Z��($�T��y"OE5���&$T��TLQ�B�V�i拈�\�Bl�b�D'}|�p�R.��T=��q�V��&>�I�1&�6o&qOa��S
��bU.��������s��L$#��H �L�u�F�)�Ig8�e�_)t5-D�X�(��p��f�t��JG3!Qa{�kJ�d&��W.M�l�B|A��G>��H�iB<eҕ�
�,a���Ǔ�G�J��Ǌ����'%��jM�q����FE%D�ɗÆ6�{RJ��<i0mjWi]�1+x�)t�DG�ԋ��[�\`�����$$��T1SՉ��K�����ǀǽ�0����M�bP�b���z}J�`B�I�Z̨a��'XFĢ"��1u��6&\��R�_%>�Ay���Bdb�'����hٝ�M�u��)Wb���S�I'
$��;Ԡ�qy�y=�pQY�%RF�hT֘|Y�\QpP[�#�2NZ��o�> �� ��W�(*�nZ����[��P8�����61͐$Q�B�$ �Ɲ�Ʌ�^��`�Y2�c��]r�)���El�GT1:��؜ZCf�h���X�̀Ն́?9��3G���hځY��c!ˡ���SL��;'�R���	)/��q�?i��Næ�;3�� �0�WjU,q(��	0�;�dE�"�
0΋�sc��	�C0?%V�������YV�0�˘�i��$�2hY���M��'F�M��.���5���ȴ�V�2��	�A��MѮ�'��D9&�<	����Qm�y ��X�'�����M�g�'�.TK$��,�I���Z���@E�R�r�0�F�'>u&��=�����G�D�ypS�H��80�aKcӺ����)�q,A+%��� �2���	1*��N"��#��N���$!W�1��u51|Xvu�d�ЙR��يt�`��j�	٠c���b�韜+a��q��Jc�?��5OhӃ�!|?H�:$G}ʰ��֓��*�@�v:`�4ZF��E �/-H��J�l ��ΧK����eO
u	x(���Թ6�� ���*���R����?L�i'��K4�D|��	R$�2kƤm��Y%�J�B�"Ml3fM�I
�q�,�(��X�?���р)�l�d�Փ�$�س�Q :�f��_X��n�Nd^���Gn�����]����F��. ��s��O��'��S8M�츱_RR���Ӆ��^� �����*#�)	Ón���� �߅gu�6�K�RҪ���:%�2����+���Ґ����'t����4En��[�C�p�=�d=��t�'�D���V*\&�څb � Hk�O�M��2 �@�֎���>�HA�OPU������W�T��T�^4c%U�HJ�M�􃚻z �݉b���*!Hˆ��O�'����㞩�0�2!�O��p������8e C�~�o4w���M3!�|҂M,a4�Y��H"4r�1�wbr���Bާy'�ˁ:��!g	I"ftzJ�bA7�M;R��O, K��^ �^-&��Y�t�&�۱Z�||�@��)��a��E��.	�JW^I�3S4Nb���q�X���uR��l��ic���R�֕9T�,5��F%&�)�O
@���F	(����c�&o:\ى��֊hn-c�؂��dۍU���X��E'|���E�{�����I��bG}�#O�}th R��3E��+r�i������"M���q���~Fz����Mb=07F�G+`�B�t�i� .�#3�4�{H<%>��E�~z'�|VЁKuZ�I�|"&���7��P�c��a{��� ��Sf�3P��P���{<�^����J���!�����H����#��Z�ˋ<z�	B�nM�&�\�h
�orH�#" �ua�p��"VtS�+��Y��;U�����A%�P�	��ܨ���Ǝn��i.\�c�I�0f0v<j��Y�[ 0�hP"�9{��Z7 a8ըT63v��֮��8���)�8
�*���C�- O�C�^-jnB����B����Y��(ЩA�=Fx�f�1#Y���Lέ]2�
7FL�_�1�MI O���L<%>u˴"����p�'�%q�I�1hq��1:Y�EFJ27����Ӽ�B�S /��PBӇG	O�V��NG`}����y�JO=6:H#�!�7�?�ë4�	�/XcT��&/���3r�`��A)k�er��9 ��	�|MJP�ꎔ���1��l�1fS��~rOZ�<)�)��r"�D�X�t�)����!�ē�04r9�%�4|�	�^.�!�$J�z�d�h񲰻"��?�XU�"Oz�
@G��qM��r�Ǟ :��P�"OdX�b�I ,yhgi� 9�p�"OP�;�/�C��A�g��@Hw"O �E�C�.� �s��ѫ����b"O�<�5��68��`[�6в�I�"OL ��F���+ �I*V�|�"O�"'�X�}2�j�-�"�҄�w"O�[q�y���я@�aܨyi7"O� �	��4�C�W<'��]�e"O����5/9�	q�'=�&��"O$�U �� ��L�E��S�"O��I$����Psq%�Ѧ��T"O�������Ij�mx�c�}܎��A"O|�@�	�x
}���`� ��"O�+�5{�B��J"=f�{�"O�Xu;Y��R�+ �H/���R"O��E�Eҝ2��Z�-.��"O\E౬��c�hʆi1|(�#"O(� c/�>EWx��hU7p֬��"OF,��%'`�[��\���D"O j4@��x��'	�~�h��"O�d�ϘG�Щ�R�6J$Q"OX����V��x�B�o��욶"OR�YUBP6.ۦ�R�*zPA"OvtZA��2+x�pp��9'Kl<2�*O 8�1AV�sA�uCB'� t��b�'�:Y(�̉��j��6�V�� �z�'���k�dØx�4��$��@��'vp�`�/ryX��Şr45��'7�|kW�N�)�v2g���`��'��phQ-0fkjEyq�0�1��'�f� �a�7&������Z����	�'��#�d.FS6P'嗛[���	�'�F1�\�le(���	�T�̜i�'g2�21LH�{��4u�ϦZ����'�f$���ؠ�ty�tM�5a*HT�'���(�.O��$� ��
$�eH
�''(�2���c�t��3��}�jDB�'�ŃC��9"DH��h]{S��Q
�'?^�z��10�+�=l���
�'\RL���P!0��8S%H'h��MB�'��H	�@�6@.:q��D��\x`e��'(ؔa�AʄR;,U��6U^8��'�(��g�wl`p��˶I�Vh�'����`�na�p�X&FB�5��'�� �����-sc���H:�
�'0�d�b�G�M�1p�bH	tW�U�
�'�ʘaGð3':���GU�t�t`�'4��i6h�5|��ㅌV�zs���'����D%F*)#b��s�H�	�'��0z�I�~�J4�1���vl ��� F!�ϩT���'ѦBA���"O��QD����r	�>&$Q��.P�ԩO�gb�ir1�6Z�p�ȓ;���[��l�r�q�f�$��ȓ�c���,\����`�꼇ȓ@�	�Ov9��b��yJ$H�ȓ<���c4ͅ55�L2'��(!�9�ȓL?8�R���8Uk��3,�x���0� }jb�\�/Ĺ`L�/$M����-�q(lcD�mi�m�%f?���ȓwT�$J�JF���S�ZG3$���BuIa��e�HA�d�&J��1��,l900i\ z���HA��C'��ȓn�����_�<O@)�dgK��
 �ȓ����+U�]Vp���"X�ݲ��ȓ[�����^$H1�� ��*��>Y�WK
D�0�G�b!���DJ��89
���͜l�Q��2aPQ�v��1��ȓB��%С�	D��1����n����?���I����&(ʝ�SJ5l	����1�Z$AۡM�@i�#��ڙ�?���~�d��a��L��4��ɂ�O�<	��/��hAե��;�|1F�I�<a�m�0a�~ �a�8[�|ի��GG�<�TG�6��R0MD3)�L���F�<��O,n�i3Zib��ȅM��~+!򤌈��y�mÓ�x��^!X�!�X��@�RoE@�,4iC+�'�!�D·-i�hB�V���IrC
�r7!�ḓP��1�w�O��<m�fE�s+!��>aN ���0BĤ��R���=���G�4��:L��H!��I� T�S,��y�EؒQ�j�q�#ʹvv�ys"�C?�y҈�W��僢��?�hHQ�G"�yr�O��J��Ш:$$�$���y�)Z�	o��1�.�3� )�t/Ǯ�y� T$ؙ��*�4Sܚ@�Nܛ�y"�խA��蓄C�:$���?�yB�P� $X��ʨ��_�� �6O$]�t�nct��DJ?�ؑe"O@1�K�@���(�i�?h�ĭ �"OL�1�
6-��X�T��2����+�S��y�c3P�ʕr�OҀoOVY	�K��y�k�0���˲�O?faiauÚ �hO���� H�zq�2�K6h^�9��C�azB����0������	�^]����Nul� �x�I��}9T�f��%XH��!����<	��ITPU���<1�lIE���:ЮC䉢z�����D�;8�[ l)[�B��4I
❲q�+��$mĕP4�B�Ɇi��H��ձS�eL�l��U�Т<E���X�;�~ p���h����4�K�y�_�#����d;B1����)�yb�Q6B\��fOD�Y�,���b³�0?9*O�u��CN7{���eI\<��,P"Ob�)cc^<~��X��1Z��M����OX��&DYoNe���2p(�7 ���p�'8��	�b���&x�4!@�|`B�ɢy�����s�ٹ���q�����/�/���qr͉	JŖT��Z Ms��ȓU����je���-M&�t��C�J�x�A�z"T�cI�*�.��ȓ_�؝�_$'��)sh�$o[Z؆�(�$�1DW��h=��D!ˤ���S�? �����?���2jD�,�8���8O����ٕo�PB��[��
�G�,�!�Ą�H���ؔm��6\!D%�
Z�!��	�H�$9
�M�ss�0�tj��/�!�$��
�p���#��=�����;,!�d��l�AㅒZ��-����'!�#1B�1k�]������e�!��
{NX0��hٲx��D�w�*+!�;�&�Q@"\#4�\L0��:p�!��qi��K�"ϛ|�
�3b�r�!��4kz�\R��ܤ=+�`��c�(+�!�DI�Ĭݑu
@���� =�!�$Wm���Ã�+ �,cSFX�p�r�	4�5�S��?��E�u���'�M��pE�1��c�<����KF�`�2�V0l�E��)�v~��'��Ձ0A��&��u*��kk\i��O�ʓw;���`�#���5F����,��q(D�͌2�p�H�OӲ#���Ez"�e��m)9w���6H˽A��[��y"-T�|ؙ��R�:�
��Ύ�y�4J/�����\u�.ӭ�y�@�[y�Lc�ϛ ^�X�B��y��S	���w-��tC�C�c� �yD���,x�hn^���M	+�y�O�j�~H��F�jE��#ŗ�y���K�
�����i����:�y��» ��]�"\�_V� &����'Zazr�EUo\�	��-	Tj�2B�7��x�C՘��;PG�R�B�j�K\�aꓑp?q@NF=A�|�e�ɺ$.t8S�+U~�<��L�	�*Y3C%�7.����"�N�<94b)����RHƗĸ���@c�<a�6h&�
�E�[�mb"*Zv�<��,�/�t�YDN����Bͅt�<yq�K�3���z�N~;p��B)l�<�Sf@�4��t{�Ĕ1kض$�)Jo}�'��|2-�U�ȁc,U�#tڽ[�e�۰=�{�j�4=���`CȎ4 �QG靖��' �z�*�_�\����Q�2�`A��L��~��)���>��$[.�pe!��W�I����J�<�&M�������
�L�ީ `I�J���=y�r覹Cw ̿J�$�Q�a�<���D0xN #`���S��;�#�`?q���ӹ]��
"l	�Tʽ����$�ܢ?u�S�T�\$�R������3���s�B�5REKI�Y3�ā�(�[���'��If]�����<	j�N�F/�B�	�AL��"��r�4�-��zU���B�ɱ����O����]�1�'o�%;�4,�c"O��ۓȁR���7D�%n� ���"Oh;��wZ��D���%�Y��y���!;������4_ �j�eM�y2i^�h�.t���82�J|9B�� �y���\n�e'Ȥ%'��a��8�y�"ߠg��5Y �̅!D>�j���'Ǡ�=%>��RF�%FR�����D�tL�4m?D�1c��R�5�S�Ϛog���9D��q�f?1v�EM��z�sӄ7D��S����-�dD��S�\+�@!�$/�O*��u���F�������>13�"O �L�x�湲׋�5��Be"O�kŎ�T��ݸ1� �� &"O�z��	�2����*ͩ}��Qh�"Ot� 3�֦F>���1i�C�ār�"O� �ui2iB�a�Rd�E'	�`��ّ""O�����A;r��Hׅ��> 	��d#\O�\+5�U%w���n�;1�	��"OR:6�NPLkv̝::��)�"O�e���qY>�����O���B��'<��"w/P�G_��*��ǂ�2iCү)D����G�|3���S����'�D*�S�'w>��w�\�g�����\�R��̈́�>L�]��N����0��@^(�ń�|�z�� ��� б4�ڎP�M�ȓVD�لč�DkP�Y ͦM��7@��Ҥ\9L�LiP ��9�.X�ȓ��bC�Ve]M3]K�`��i$v(��I/�'�^�ɶ�ȓVA�<R��	�h�V�9��/�� ��;�d��U�V
�Y���+����H�p�bo�M/�(x���5'�ȓd86Q���,��`3$�?NP��ȓ$Q�t��$eT�+QȌ:n�E��_��e#��`a�h�I��#>�1�/�.�`G���=+q��
�la� ¬Z�J�@��'����ȓa�����J��\ؐ=:�AH����O0r ;B*� ����4n���ȓMĜi���f��T�`�ʰI������^���LӉa���1C'>��̅�a0�+�eM�S�b���&(6���w��ę�G��_i~U�
W��ȓw���It㟫>������J�Fԇ�P��Y�!^�c��C�?n�ćȓ4'<`B7����¨
�E�"Q��X��tY ���:u�D+d�ǒfR]��UN$�CID�;W��)��]��D���7'@��4
T$��� �����=�;/�@���O P�<�$B:#\鰔%��I��)���N�<!���.%���I&R)a�]Q�<�-	~n�[�$�Hz�Qc%�O�<��^�m\A	���Y@�b(AM�<IU&|g�d0A�PE�b��`L�<q ���O�XamT>JF�sS��M�<	V-��q<�u ��2�04��K�<	�!͛��`�	�U��86*�E�<ѷ�ɢ!��lS�DC�Gmf���N�C�<i�M��H����Ȇ#�	��I
}�<qu��('/�XHT�k �N�v�<���K�|��$��mI~О|	 �t�<�5n�/�8���܂ ��4�Bo�<Y�̋c���&̤t�p YF�Xk�<��bӒ,[re��+V䀒�@�<�hS�}�|���V�%|\x��	}�<�@`ǘi��H�B�`�neh!c�u�<ц�\�fT�ˑ E#V#����C�p�<	T�ލ]��Pp�a\/��B�<a �P)=��[��D�1d\�3d+B{�<iw$��T���oF�:��S6Ow�< �.;<����*����"OZ(��WW�z�����%<B�+#"O>�:�
�+3Fi��!�}\S�"O�����6 hژ34�F�f���"OZ���D�*1xlS�S�FF��"O\(󲎝�I�\����xE����"OJf���L�%JL֦.��"OX�3Q�F)pj9P䚂/8m��"O� �,�oI:��!�e	����Cu"O)����u�򝰒g^�I ���"O�ʧ��I���w��"���ȓ;Ǻ�*�U�0�Ѐa`�A2T�����{f>��dGB�F�y�◔�4�ȓP��u8�ƕ97(Q�v@j�
���M���hag���$E3%$�$v~���X���0UdL�dzT�ڱdN��^̈́ȓ�.8`'c9&�� �3"�9d�m�ȓ_.@���F�;/t���cj��H0�ȓ�x�K��ˊ%�ى��
�A8%��g-l��Є�,8U!aJY�^��ȓY�a�hIO�d�l��>	L}c�'��P�a ��U~5�Тٔ7y�1�
�'xL��ei�4���Y���6䮡s
�'��9酣��F49P�&(�dђ�'D�h��/gt�x�w��+#��k	�'�t`:EM�)[�����J=	�T(z�'����#"�%u�*�2�k�: �q�'ad��u^r%2��]�n��y��'��r��_^)�Ds�nߋSu��Q�'?�ݢ��l�.9hE 	�z}����'�����,{��5�U��ts��Z�<c��2C\Rq��"_�%�PE�IJ�<i�O�mÐu#t`  ���[B�<��E����,��hډT=xICD�C�<��!��^u�����u��I��#k�<��M�[�n��F*A�
�)��c�<I��R�6	�!�oOH9��\^�<Iw���^��` �A�x�pɸ��u�<��ꁍ ���� �l��e�4�Xl�<A&)�7V���J���^��@��Om�<��A	V+bdk��E&Rb�pc�aDC�<i3I�5�d-s��+�	����}�<Y�H��a�p����>6�R��|�<�SjC8;U��ӄ�r�H	����s�<Yc�I�D�v�a���^���'��s�<�.�Bq�}Rf��:h,\kG�v�<QeDۂu�pp��<VFUSď�s�<�d��5�(��:d�,�ᶪ�e�<q��Ѡz���&BY2nt��dXm�<i�C�j�BA�P�D��0	1+�k�<y`eȝ	��iybK�6>��0�"\R�<�Bd]=g`jH��$�x˰�if��F�<yw(�"b�����$�\�y�B�~�<9�A�A��bK/:K�����}�<�rIӧ2�Xaw�ǢD��I���P�<!0��Y���@�"�}�	B��I�<飉S �ĩ�	L6.=X#ĀN�<(�&+t�L��d�+=���Cv�<тL�Z�ƨ���w�� ��v�<�&���X�|A{�GB��2��ab�s�<�g�@��~8�f-�+L�6���R{�<YQ)X����A�F%sk�P4B�t�<b��z�ʑ��	�y�EC^�\B䉠MG����ſ2�hb��2*F2B�I�,��h�L�(�d)���A.B�)�H#�>T}P}A���	c4B䉕6ڨ�6o�#p~@�����BqbB�I����� �_@�Ga�W�B�I~�E�B'i�R��cU�@�B䉳t˖�� �6yPzr4��D�C����[1�$S�68��1u��B�It�؉	�ŋ^}""��.	�B�)� ���.�o��y��L�M�R"O����.�0��e��; �y�T"OtzD�Sqx��G�4I��x�"O����p�iPmN�:��� "O�\�f�?/�������Liq"O*dapS��1�Cg�*a�r �c"ON�x�nM!yY�0!L!Tܘ�"O��z��A�v�<�V��
�P��"O��ȃAȉ3�Y�cG�k�!:"O�p��K;8�a�9ڞ\��"Oh R3&�*I��b�5���r%"O��*хϧx�(�@"��Z�R1��"ObɛQ��&;��p@�Y�ӜI�"O��y���)x�	� �k&�0	�"O����ұ|B�<㲡9�UT"OԨ��#4>Et�˷%ݱa��i�<���� �+�>q�lP&��]�<�s�	4h\ۂ�Ih�! ���Z�<����#8M�8f�S}6�����X�<��.R}�nM��C�:&��`�}�<�DL`@0�ɔ�{���@�A�<IO �r�� )ӄ{�2����U�<Qh�i�|0B��0J����VF�<��I�u�YYT���0�,��-�C�<I#��t
��k�aUEjZh+�͐d�<�V�Ћe��ۤ����千b�<�X�$�^)P��2"5r�Sd�^�<�Gf� $�T� 吵C�,{��r�<�r�O�!��F# �|l^+c�n�<i��5SUм���
܌q͍j�<q�����̃q�H�b�:�z�m�<C*I4
���i�W&4�^�O~�<i�@Y�<jI"���7$U,�0�d�D�<Y�����P�2EN�c=(��'�C�<��5~R䱪�$ˇ]<���API�<�&c_� ����g�Ӽ�%cIG�<��>D׎Q1̌7::�y���A�<q��E�T�օ�� �e:��:c��A�<���ƴ�8I��D؍k1�( ��@A�<���=w��p��Bɇf_��Sh~�<���11l��B�N>���V"Zq�<��!?V��Ū�vUZ��%�l�<��ʁ !ܨx����j$J�0'%La�<!s��ub)�V�_*B� 3B��x�<�e�J�!$�(�+R�Q�&8�R�x�<I`�D��4�H�n�:����MAs�<YV(Tj��KC��N���Ky�<�rcF�~qK�ۚ�P`Ȕ��v�<���8{�ґH'fٙ��I�5nCY�<iSI5E8����Ǫu0*tK��V�<1�N��Ǧ��B�ſ,��&��y�<	���\	Ȉ���8�N��A�L�<9�K3���GC܏f�H-(`F�<�F[z�>͐v(�>�l�s!PM�<q揇40�@�Ѡ`�=�$�6&E�<��ɕ,��y�JΛ}�N�d��C�<�Ш
�hѨ�#b�B#g�sb��Y�<�IL�V�����n�m�D��h�|�<���X�D9�0M3�L=#��c�<�R%��H�\�������P��a_\�<���Z0p/.�����H֩�@(�|�<!6��e��ыY�P��{ӭ�L�<92b�?��ѓ��Tf��+��S�<�V
:�D)t�ńJ��䉤��Q�<� N�b�+
�=KJ���L�[�4�P!"O�e��4P�d��"WV��2"O�Zsm
�M�j@�
�Z	�"O�x�e�)f���$8�0��"O>p���L-M�N���*�>��y+�"O�!��b��y�,�4d͹F��uے"O�`ۖ��G R�1WeZ�K���AE"OZ@�` ��|�zw$*K�^!a"O"�!����:�|҂�H�<���"O
9JCK�8����`@;M�1��"O2m���P�00!o=f4�`)"O� (���[��"�T8y2j(�"O8t�K�_�B�BI�q1*�p"O
ȃQD�$1Pn��!ǒ�DB5G"O��
����h���D��$Z�ʰYG"O���QS@-���ӈ|8v=�"O�9'(̦9f�eH�kI�j}0�sr"Of��iZ,
��l*c���4oH�q "O|pCsD>���F�-�Q"O���AJ�2>IH!�3�� N�����"O�X�g�ۻ/�6,ȡ��?r�"�
�"O��
��R$<�� d�;��] �"Ot�X�o@�������`���"O���(��"h�eA�KFlm�D"O&�1�k#Jԥ�!@�@z]�"O#A�T�P`� ^$l/�{"O�1�S�$���Z�M�'3D +�"O�!#�/� h�2��ʫC�V��V"OtQp%L.�Ш�V'�����r"O �H�DإW_4��ù9�H���"O@M�g����&����X�f8�9r"O�-���ъr��h�4�߂G�~%��"O��rP,@��=���ߩh�.4r�"OX�E�Ƭu���Q֮.�>!�"O��`����73$1��K.{hr<-�!򤀋�.E�`�ƍw��� ����!�D[�g�"ؙ�O�;�jdI�d�/Q!�D0_l��&�]+�����=�!�J�*�YJ�h��A�l��F��7�!��*X��<U���u��Ѫ!�ƍC\!�D��6�	���
G��]h @��Q]!�$��n�PYr��Z-�iY�!i>!�$K�N��$@A9
?,�����(`!�d�e(� �Ǐ�<I�Y�ņ?!�$	��j�a G�+���g<d!�d�+	��r�`Ï;#�A+�#�
!���c/ԄBs���-.��S�%K�!��+�ٹ�� &�(� 6/�!�I�~Y Äī"¥�w�t�!��/
̱�A�Q=(Q|�k�E�6o�!�T�T���C�̇|��rk�5k!�Ĉ��"�qq�� t��a��55^!�FL<S2���X
"U�s�ܠWI!�Đ�t�����X�A���P��T;M6!�ā�i�0M�)�o�X
��Y��!��ɪlȀ��j>>���S���]!���#sG��( �~�HBsn�jW����U�r)�SK-h���(��.�j��ȓ~TQcɲy�����OB�ȓ��p0��'���2��Э����������e	Jz����*Tв�ȓ	hx�)��1q��J����9�u�ȓG$��K�NZDF�M�� +[�p��ȓvXT����o>X����_$JI>H��S�? j��AI��&���q�"��\�p"O�E�/h�:u�G�9�|�
�"On bࠀ*��(���}����"OLY�$J
i�Q���\k�"O�ݫ����>��Eb"��lvp�[%"O�T���,h�Q�ul�9!b~0"�"O  ����sJ9�aI,��]#�"OԘ� �e[���#�I8A�ڴ��"OR*�e��X/^M��݋X�T@��"O�и��>0����Ȳq�R�"O��:jͶM����tF3?���z%"OH���*����	q�[�$$�1"O@�Q��	$)"j,;,"	T���"O����C�&(K����Jl��B7D��q�&v���# H*+V�ܙ �(D���ڼ�����n»^@D�X��%D���ǌ	A/f*���]�Z0��k0D�0ᵂ df��� �r�G�!D�$�!(\�V�OZ]���PFe5D�|B7j�,\�lպ#��>ٳu*3D�T� �jhtr�։s�&i
#O>D�lA�S5A	���t�rp<D�,��h��>\�����&���b�m'D���#����0X�p,d��d��#D���N��w�����	�0��u�"D�@X&�jas-��f���; �7	��C�	�$ ��j_0�~a�e@٪C�.B�ɱ~���b�	�[�^��׫�b)�C��$킍�Pf�)2�B�f�s��C�.D�t�����G�q�p�i��C��
���dM�a#��!~�B�I�
Z�Y��EMH܌Ѱi^(��B䉨����EФ������0��B�ɟ;�����ؽc�FE�B�	���h��%�ڸ��FL�T��B�I;|)�L�h�d��A�	��o��B��	��@g���k%����D� :}NB�	ff�q��)�A�6uzu��6Y�dC��E�<����?i	QY�)đR:C�	3V ۄ��B}��CVF,� C�I�m�ε+�͎`��E!�a��'�C�	,
ʨ@S��&6��LL�.\C䉨 +�tR2��+��UR�n̈KT�B�IS�d"��P����/0�B�	�,��隁ˊ�&zقf� <uh�B�ɥ�֥���*���A��Q�lB��RD� z4�C,]���RO�!��B�Fie�׍�%�p Ӂ&C��B�	|Z� sq�҃p�2c)�-@�B�I��L�'�O�54�B��8|�BC�I�S|2y��`�{Y<RDM^yC�Ii��-�%Ǔ	�@�؆�2�B剮nXX���AB�?����N��Zh!�%��9�䑎]�0L��!ST!�d�y��lirn��<�Z�*���o�!�Ę@�b4��ܟ��t�7���!�� 3��|���	;/�������!�O9G (�)��q��%Z�iяL#!��>KV$�vj��ʘ�h�1Z-!�I�4[R}�L*�ڑK���6Gx!�d�;n�fɃ��؝����x����ȓ�0�G�9L4d���׉VB͆ȓi��*D
�j��)��#$�%��\+f�IU�6�,�%�WS<p��S�? �Q P��@��[P �.{�4��"O�r��ժ|�Д{�!Т"U�l�!"O�c�E2J�qu�_?#C�#"O,�{�L/aB�#�II�/8� �"O�)P�
�� ��0�Œ�%��J"OVVː�V�>�ʓgͥ:�4��T"O��  �I-B�@L�@��3b�UH�"O��c0
R)|�t�&�ڪ3$j� "O��b���k?,���;L���"OX�Za�߱$*�T�K:| 8A"O� ů�{`�{��M�+Ds�"O8�G�J (�(�X�JN�Ԓ"O&���m��y���¢i�	ai��;"Ob�@� � p �"j
�\�*q�&"OtD���!h_�(�2k��~�X�2`"O@��ݝV5Z�@�j�>���"O��2h\�A�J���)%@��Ha"O>)�$�T�=�d�N&H���l"O�����00�D)��Y}ⅳ�"O�,B���
�,��煨Tvd+�"O�pÅ�J�`2��R��ֿK|@$�d"O������ Z�\W'�*ht�Y@"O�5	@Eڔ7�,d!�dZ#fPjH�"O �s�O�2����d>|?�9�c"O���MS���� eN:���"O `��#�R�P]�#�V"tL��r�"O�-*��8g���"mťX?D�"O������޴;D�߉
1:�"O|1Z mװ�va��%bE��qB"OD��B@&d",�Y�.yP��S"O� 2-޳��s�K�_M���"Op�Ԡ�#Y��iU+@�?7��c�"O���娔�"� �8R�#2�|cP"O^y� �̾,|�xض��1.%P�"O`T��V�k�6� G_�,�F"O�|�,�����{G��i�Fl�"O�����x#�AA�̎��h���"OlH�n�	�l �LT%���5"O@�����O��+�P
��"Ox����L�*-�\ T��\k�c�"O A�DU�k�<Q(���g8��"O8u[�JF�U�D��7>o�L:�"O`�ɴ�Fy
����(�=2k\��"OT�;��D�0�%�a�`@�z�"O�����q�:��G�LZ���"O,�u���%r֥I��Q�FV8��d"O�5S�+����� �)B�p���"O���&�%Y�1j���Q��#"O����`[���)3Цʍa��"OxBe�X�"�X�K_<[ӈ�8�"Oܕ�w�Vi������+�:-�"O,��mʪWlj�����D�n���"Ot�cB8d����Ţ_sJ}��"O�TZa�X�s�V����Hd���!"OvH��'AH�c�;� ѐ�"O~�i��hMFuȡ#�^�lP�"OF� �PCļ{Џ�7��@#�"O�$���o�J��@�F�^@��"O:�Aυ�\�:T�#��0&�0yi0"O��i�/A9zkx�p3E��B�Nqt"Or�KѦ�*P܆����U50"Obe�����
u�
P82l��"O�UAWcݜLՆ���2N+"O��nЫo��8聉5ܰd�6"O� <,�͚�t��)!)']V�b�"OVڇ�A�Zndъ0I�a���B"OVh��K�-��C��W�oF�ыv"Ozi���q! $h���:갱�"O4Å�ݫr9�ыp"׀���E"O޵�6kB9/�i��T�dY��"Ob12%٨?���f:z���"OT9{F�rp5�f�ƾ
Ը��"OX��U6�4��q(�jW�9�T"O��R��9ߌ=�!ɻJm���yR�I�Fcx�	�D���	���y�e�@�v�z�E�
S[�|����y2���0H��堙�`�ȕ3�g�yR�b}`B�i�;[98ŀ���y�L�h�z�s5*��d�T����3�y"ET�N&�@�ņ8�=9!D�5�yR��p�veJe�4pX�p�B
�y��.Jt�Dƽk&(��F��4�y�&�Z�"�{5��c h�0�C	��y��r�yf��U�xp�C�yrk_*�b9b��K����y�Xıb�q��UjW��$�y"
�u���hSm��:���!n��yR�A1X	T �H+G
ܽ���R��y2+U��
���.đ?��jҡ�y�("<�0�����[aȜ;�y2�������ߴm�X������y��T2XY��&��b�rТ `O��yr����}�f��]���!s�y(T2���� �^= Y�<9ҍY�y�GE1|�|QS*�NFxm8rb���yª�%N��]�B�Y�Y"5���#�yb+	�5�X��s�[9�6`�E���y2nݰ>dZH�t�H ֪"@�$�y�T�0ܶ1Z1Bϼj_0]R�R��yrd�+����!�^�Z ��D��y�H�n9�k�"[���b�	�y��D�0/�q��jǣ��0���̵�y2 �zn΄��+@�*Cc��yr�F�f��l+����y���c�+�y�풷:��$:áܿFХ��J;�y�K��2$X��C\#��qq�,���y���KмX`$D�'��r�'��y�ܕM��5[�m�V�����yb��;���жdT	@�x�L��y2䈟�D��R �*�PC	N�y�J�=a���g.	r8��!����yR��3;I9��\�ql���`�ڠ�yB�-*�yC���ذwaD��y")_�P�T�ە���*V0���y脎r��\:��<��eصlF�yR�U�JaE��ؔ9��@ⴭ��y�b?Ф���1c�Ũu���y"��s�,՚eŇ�V�0�S�$Y6�y�	��(�6�1�I�"��<��G�y�
M�4,2���N�-��L:�y��T�l~��P/��`QK�V%�ybD��}v�0�b�V0���g���y���6u6!�%ER�f�yb�_$?H��v���hZ%���ݲ�y���;v��B#c\<	���x���?�y"�ͱO�nT�\i���1��H.$v C��(TD�Ӥ��)bK���D!F�w��B�ɟG�r(2�"��`�����B�)� �hj&��=b�b!!GD�2��[�"O*�K�.�vN�1H��B��rXq"OT���JO��"�d�-n؁�"Oz�,�F�z��E�l]$���"O���G.Q�& ��E�f!h9z"OM��mM�RnL E � N��"O:Y���zX�E��N�
#�ư�"O@lٓ����U��L5/�v��R"OD�R&�	
/`�����MJU"OL�A��!d�xD`'���e�!��"O��W���Q)n) P�>6�6��"ON�A抍8D��4Ð�q�Ρ+T"O� ����IT 赢	n��(��"Ob(a��BQJЖ�@�U�p̑�"ORY!�ɫ`v��`Σ(�LP@�"Or8�U!TeM�=�
O	O���`�"On���NW��`�d�.\�x��"OEh��� ZJ��4 5! |��g"O�5A�FY���M���$�B"O��	`N�)Z��-���vDr�"O�A P\�X,rp�r̟% �.@xf"O�hj�)ٛ_ժ�!���=岠��"O�$ ���	|��q���T�1����"O�(0��:#������&�n�;"O6�!�j)�W�.�"�"OM �A
Y:�b��n�:�XU"OJ����X�<"��䕜2f�h��"O�
��ܠN�|��rd��s5;	�'���&ϙ�4�f���Ɉ*Ϯ��'���`�_�K9XU�7��́�'�^}r�F�*N��!�Ȍ�j��(�'���SΔ,�m!`����3�'���ұ�ĚcG^L�g��yGv)��'DBɈSS6a2�#P�
�n�>��	�'�(C�� $B*�|� �b�{	�'�&�1�a�lYd���*�=\JR���'���xr2�,�P��X0 _��8�'/
Q�u�Ԓ<��ݕb���'��t�ܖO;�I"'ԠNI,�Q	�'�}���@#�r,#�FX�JP-��'e ]�Ů�,�`az���o+���	�'>����ٰV�.1Q�E��tލ	�'�.ȋg��@!�sID�q���'���	̮g��c�L�}	D��' ��6ݤ"ZYP�_�a�h��
�'n֭X7m�")� h��ݨ]/����'f�SSH۬a�@#�`X�[�͠�'�Y��B!�8Б�f
;!�2E@�'�DI����u(�ٟ"�T��'1�x;�K\!?t1���I��4��'1���'@0�W��?��l��'��`7"�4N2x��U�=X9�'�8�B$���j��%`a�������IA��|�yTNQ!=хȓ>b(U�GhX�i[M�2Fߊ$Z����u�D)��
������1x��#��u(@ʑ� �D�ze�U�ڝ��G�2\2!*45�Z���<	d8,��u���vhE
|M��٠�Bq����N�"�jN��c�N�Z"��6�J���^��t���L*�"�/��e�A��JVj��wd���X�b�@��k�؄ȓ/�������G�2�z5�ly�ȓb��5�oS�W��@�a�x���S�? $q�m�8�āO��G Z�P"O���d�4tf�m�GN�<��9�"OƵBg�X3#⽓�G	S��� "Oy�V$[�<8�uz� �f���!"OJ�jU�W
H1���Teq"O�� �1v��r�Z�_���@G"O� !��ޒ9p���-���i7"O�!�g�.��kQ8f�BT"O�|Rb���H��ʁ�l�N<4"O�Px��+~�n0c��P>^��IH'"O������Z�x��(�&&�p48�"Ob9ϛd��P�w�^%u����"O�8�1��+V
�� '�	�~���"O�DP�D݌k8i�f%m��{F"O䜑� ��1`gÍ�`dꍩ�"O��BW
E=�ȜX��
l3H�[B"O��*T�%G7Ƽ�q�i�lq'"OH�����~|Mx��}�1��"Oֱ��/ϕu�\`FJ�g��18�"Of��D5wÔ���ܫv��4�"OHWk���,L`��V���!����{)�|J�-jt�8�7P��B�I6���W�B�i�J� u�B!�rB�	�)r&rg�@�<z�+`�<aPB�I�e'�Y�0M �o�)����'85jC�Ɇb2����M<:�2y��!�)�:C�ɠmI&�H�1H\�2G%^2�B�&H�d	0�ʜ&�R�i��"`�B�I'y�(,���($����&O�&X6C�	�4�N�����I�haE��&#�(C�	��x��$_�NG&eJ��O4C�	�o���4ES&$)x׎O4r) C��Q�ؤ�V.�p��{&�ϔ*��B�I�%���S�#�0���!D��B�I�Q���x��J�T�)��ܻS�B�I)@|⹲�
��C(��
U B�<B�	Y�RE�6A����d2B�WF��H��F,46��@�"��C�I�	�i�蓉Y��z��٧-L�C䉫#�*�se�"��#�c�!�C�(=��x��A��D�a>O�dB䉨/:�{��JWU(P2qT5<2B�(C�"�I炈%�TTpc�5�B�I�k�HHz6aO�H3v���&��q�B�	��lYӦ��	fx����m�TB�	�%�<Y�M�"[�^�9�h͎0lC�I�XMΈ��$�%<脸�b���2C�I�T�c�HÎ_ ^�q��á��B�I��@������`CT�I��B�ɢZ�6�( �Mm�4i�9��B�I$H^��8�G%I*,=�����$��B�	�|s��i�'L"�&�b���P�@B�	�L������P2	3AK�/.�rB䉷/:h�Cp*��J�� ���5O�rB�0^p�%�s��V(VIᷤ��nETB��yz��z���Z�H�!�z��C�	 m��Iq0��e�.���;ȢC�ɝ�L���;����΋�b�B�	�6�<�0B��07�@"�(L�B��Z����Ć�%ϼ4I��XƬB�ɲu١2�(3���2�Η�;��B�IR�|���J>�hP�
Խq�bB�ɊH����*ś����Q��f�8B�I�c&
�hA�O)��	 �-�DB�)� ��C6�V~8���F���9C@"OVT�T� ���D��&��QBU"O�@i���4�v|RN�	Bt�p�w"O�h�A�@�.�8�aAφ�[d��w"O�\�R�[8 t|�Ь�jo�U¥"O
(H"��HV�j�DFP��+�"O�݀c	Zw�ʪ?4X��b"O<����@�l�|;���G.��R"O,���l���^0Cs�Y.1�a "O��fAݫ*��5)T�{�Js"O�����Ǥ*��`��ߕR�`�Jb"O�8�r(&D�Ii�a���V"OԬz7���B6�
�Qo��{�"O����� d¦��(� wz(�C�"O|�q3g�n���]rٸW"O��J��@��х�z�n��"OJm�v��9�=��#q��-��"O�x#�.��h�vIʫI���Q�"OTŨq�1i�3Ȗ�*ɰԚ"O�ɐ�!�8�9z�d�F��5A"O�[�# %<Xyy4��ms�Q�"O����[��&�{c��`�0��"O~�����B�B�*���J�x|!�D\�q����ЬJ
x�$��'.!�D��`�Rg�@�V�C`B��!�D۫_��P�`�)&���%Z"aW!��\+�,�C';t�Y8 ��:LQ!�\�-9v{����}�����W�*C!�	61��P8�
$(ׄ�ǅ��)�!�O��=2�g���@�Ǣ��-�!�dе5F���*\6S2n��&Y!�DC=w2���+1ڌ2Ҋɣyb!�$�9[���TI�18K"xPW	A !�dJ�ux$yk���#�n�8rNľ�!��?Cn�Siϯ	TF�f�N�,�!�$5`��!C�6b8�a���Zn�!��J��H�c�KQ�-�5�Ik�!�䚐$��p���i4"��E!2�!�D�watЁ��r6�D)�B���!�d�.$��x2�E0d&"ȄbQ��!�D�x�t�م���+ V��&/�!�� �����5$ita"fd�!�D�B���"��+f��)4k��*2!�"\k��Cf��)X$l��A*}�!���3`r��f�e;2$� %ɳw�!�䜖L۪P�d�+��
��z\!��x��h �ɏ��p���Ԑd!�@<�,T��HGr�\Y!b�V�x�!�D̴q�����	�@V�,�2 0!��݈pQ�q`���;=䱰7E�G^!�D#;8�1��Y<�����	M!�$*~�xj�I��U��X��?~H!�D
�_{&���.�1m|`݊d�,}F!�ӄ)R򑐁��q^.�g�S�<!�D�~�0�����0⦄��2Y!�$��Z� ��j��2t��!�jBD!�$�--�(A�o]!M_t}�*U�!�d��t(㴮E�qi��X4��,�!�I�=�r��R"9POnc(u!�dG1H��7�W�'�xl0ŦC�E	�B�	�e+��p��ҳH�\,�ާ|۔B�I�*�L ꃻF]�}!'���ZB䉹<U�X�Ś�f�.͈���I�2B�	�1˦	�B��}��Q�	-*�6B�)� 6��'Q�.��@�0�è`=y�"O*85�O�4�&�r�u��YYR"O���Ĭ�%(,Vi ��U�;�-��"Od�Y D�x�CR������T"O�!x��UQ�}�C �Lօ��"Oġ��.�i�9r�P\�g"Op��3l���J$�pl�E?�=A�"O��B�*9�p���mQA��-j"O���OƵ17AtL����@v"O4��V�Z7q�\kw� -x�@��g"On���]'_��� �	Y�CA���"Ox�����ca�ű'IӀr,���"Od\���Ht4�{!�8i|���"O�xk�o[,l�&LH�E�"�����"O����Do��FFӳR���p"O�%� Efp� ��;�d�pR"O�c���!?��Lb�U�X���W"O���D��V�X�;���q"O �Kv�,v@�@B��z���"O��̐+>H��á*�:Z����"O$���N0l~�\P�ɘ(@�-!�"O2"�MT3P��r
��}%�9�"O��aF�P-�Q�ֈ��>n�Mz"OJ{Gt�"��`��
`B��"O�I�aF�A�\���ٻF"lp��"OBѲ7,� q���$D�@���g"O��%���X��A _���1�"O�5���O�a�ځ����P�æ"O �I֜q��7oV�!�Z��"Ot���E��8ޒ��1�ۉKǰ4��"O�����j�p$�"��G��3"O�X2t℔1�8�"畲Q��w"O��P��k���JTF�|gH�"O�	�')W�4�f�1�(����"O�	��?kb�(�⛢��� "OR)Y��9�*I1�gߢ#�Ā+�"O�p�s�P �t'�r�.iZ"O�%Wf3|s��QA�L�r�:|4"O8	���٣�\)���HG"O*��k T�����1{H�"O<�2���']�<(�
�u�|TC�"OHAa��X��(� ^�t!�dP�"O� ��	�-���;�>\��"OR�R%�9b| �{��j�Ej�"OL)jŉ�mWf�7L؆W�!R�"O��+GFϻz��Fh�'D���"O����/z����!<U���w"O�40�-�l��9G&��㔭st"O���D �L8ތc��M�*��=��"O��[����\����G��&i�|l��"O��)�H��/Q:8�ǋ/H����"O�<��'T&U�ʌ��!W�~]��"OF����`̴p"!7lҜcc"O:	r�JѶm � �4i��@B"OBT��aM�~O��eK�s�恙""O �BjF%*DX,�I�fQ(�r�"OP�t�ơ8��d`�ǒC��s�"O�Xp�i�F�blH��m&fI�e"O��z5銯�N�bA��1}"E9A"O�j�U?�:����5` 1�"O�Q���KH}����:G���&"OY�&)(�����Ғo/��*�"O����R�9d�s�'W@��B"O@i{��
i}@,(ڻ f-"O� �=HÊј}�*,rB�3���bE"O�X�A�	]Dv�%�6l��cA"OL�X$�C4E4�EKZ��&�8�"O��ᢎ�0Ud�0(�?'v$��"O�p��	\X!���<r�%��"OH�:���ek@��Hɗ>hl�"O�5��bE/d�~��
>
Df"O�hw���@-���M�i]xM�U"O�!���Wm8�@�M����R�"O\���,}�. �'��v�&�pC"O��c�?D��Ie$J�v|;U"O1���?|��`����Is"OHa�BG�F�I�l��H��A
�"Oʭ��^�F@H*��J1=�n��"O}"p.R�s��l{!ϕ�J�|��"O���j��H�gL�6�x%[�"O�(b���Z�v����),��q��"O���8��	0&T�V!v��"Oda�ԂI*�b�1�'=Ҭ�F"O���3�[�uNp �ţ��%�-��"O  p���v��# G�Zs"OpH�!�sF4rᡅ)sJ���'"OĘ�7@�0��)
@�E9�LZ�"O~0��
1��0�f���:-��R"Oj��ˁ�]�+���>j]��"OB틧�$)o�����}�&)�f"O��*Ĩ=<��)caP6#쐽
�"O���!k�Y%��"烪�����"O:�����A���1E�dX� â"O
ܛ�1B��ɸu��`��(U"O��ƣ,9|�Ja��W� a�e"O^�*Q�O��8p����y�>��g"O�L�cTM�%�r]�z!�Aڂ"O������&=�m�bƎ#P@��'"OY`S�\7w~�YR�"A�h��"O�5;"n�Q��i�4��&�F�Ɂ"O i;a�˾D��z!K[0d��t"OF`��������阗*�r�*�"Op���K2u��������-{v"O��{���'D@9����:5U"O*�ZC�4*H$��5o�FD~ԁ�"OƐX�'՟WU���'��:;$@�"O<U@�!��^�0���}�.�{$"O��K1)�~HX�s�5D�$��"O�
�Ù3�x���8wR(re"O��2d���� 2�@H�v���e"O.ݳ�g̠y���i�Y- ��I�"O�L���F��>%rb�E}&&��'"OV��lY*b�D���^:fz�ȃ4"O<Q�rl���A��F 0m"OV��Ro��$S�DD�_�T���g"O܅���/a�,�w�� [�s�"O�ȴb\ .�(�_�}��C�"O��QQ��0QHX� O�ܺ��"O ��6��?��ѻ�K�r0���"OBcK�DJ�hXf���$:�"O9���)�t�ٴ�E:Y����"O�&�^>p��ţ�	����� �b�<�p�
P�,���RD����+�j�<�� ,~$�5��=y��{��\M�<Dß�xdM��/Ģr�ڌ�T#�E�<��o��Y3��Q�D��:\���H�<y�"��x���`ۂ�-OV؇ȓ~=�+!E�+!b�����\��S�? P��.0lu����N/��C�"O��� FȈ3�t̑B
g ��2"O���t�Ƨ7�t�00
I=�Q"Od�Rm�'_��h�oܹ�N�K�"O� �D��0Qh���/7LBP��"O��y���R�ԓI	*y4>��"O�=���S�1*�:�BN�t����"OP%��M��{6:�"�l�d_>��"O�!pG�A�H��lA(;Y��Z�"O|�2 jߩ3�d,�Eѭo�e8�"ObU�G�I4x����f��{lZ�k�"O��ڗ�-z��[�b�?UX�A"O�\"E��;
PZ<0'���/F�U	"O����)�ԩ{���8��87"ORĂcE���T�*���6y:�"O��@��Ĩge<�@���/$ �a�f"O(QHoF��|�qD#.�� ��"O\���6%~`�yp��;�6��"OxW��"��Р���+3.vĉP"O<�*�@
,i�di��z�^�J"O���A4P���c�ħ��h��"O�bU�R8�f��)�3�$hS�"O ہ��5W�����K�r5�P"O&�� Ո9�P�c�U&&��T��"OeIG��+ʈ��V@)>�<��q"O6��
ב[�}��$I-#��2"O����%B�,z��`�y�F�qV"Oa:�R6zy�H��O�L��@"O �Sp�9R ��5O�m$"��V"O�<�rHH�jy�Y#%R�.*@@1"OX`�s���f4��p�DIR��Uʂ"O��)P<w���3B���P�"O���'TU��9��.7ޤr'"O�Ȳ읡a�xu��w~u�7"O�rp�2�ф�U�l�J�"OԪ��K�&�>IIu����C"O�`[��R��*�ȓyDX*F"O�uRƓ�f���#@�L�9ܠ�2"O�4�N�jdn[7c۞7U8 x7"O���e�ͯF��@4�5X`^���"O���bƒ�� i��C�Z����"O�Ms)
�h���TO)J�B8I`"OV�q�,-^$p��E����"O�5�'HK�
��q��.� S"O�A�S�\�rqXI��P�e��(��"O̥���K�0ɨ��0Ɲ�!��%!�"O�����M8��x*�EC�N��\b�"O�	�f� r�Dh����)l�@�"O�h�AK�6c��d� H� �ڥ"O.�V�S ����f!��Xk.8ZV"O%�k��Bz�IpG��5=Ľ�d"O$�UD�f�F`J���W��1ze"O�Q9��ѿԞ`e�Ү$I�M��"O\� بA��IUm�$=�L�"OY�dZ�@��4+�	ӳ#��� "O <{4�U+�t�S7)�v��!�"O��P�OG9U�P7�O&;t���&"O�Uj̚rZ6�Gnl�Hb"O���Rf���Vy-D�i��M�<��o]�5�^�ጻn���y d�I�<��"ĩ3�,E�G�6-�,X���YJ�<Y5�;U6X9����@���@n�<I��p�j��A��O�E
�Q�<����x��q{Ԭ�-��@2`�O�<�   �ǷIb&��`�*Ln��zU"Od����ױr�"@��j��m^��"O,����A5��t��H�[���b"Oؽ�NQ!tv�شHBC� �{"O,U*Q���� � 0���2!�L�<I��OA %�����D,]�<�(ǐa�I����gO`�P��Y�<Q���/(8���Ι7UVMP%�CR�<�$)h<t)��G'a�u���Q�<1��?\�b�k	'2�%�N�<	b!	?p��3Z �Nh���p�<��f�fo|��j��&��	2� �S�<a�Ύ?���V��$�(��*_N�<�r&Y�l����W����`b�<!��I!<��t	s��5Y��R�<�u�� t$V��K�F�Ĥ[�&P�<qFF�E[@�أ�_E�^T�ER�<Q��T9"~"�*�Đ.6�|�0-U�<I��\Qq �	?ll\��A�N�<!�0ɺuC��
�84����SH�<��,S^9dl����9zcdu��Yx�<y�N��[�I��X�R p�Z��t�<Y��\�3�^E��Y�G���Qb�D�<2D�
<yr���K�&)�
�\w�<1e@_�8���*��@�l�V�t�<)��_(�� Y�\_�(4jj�k�<q�G�%���"U.�Wb�A�!Wg�<�4�^�b�
|�eN��e�����n�<14��릐[1&��C�&�K-h�<a� �9W܌p��Ε"4�騆�\k�<�QjJ�FyC��	'�B�Q�j�<����>D���0M ��(����J�<���+�9�:Q|�ƅ\�<A��\ԵhU[29�J5`q�l�<��� �i�SJ\�$�`a��]�<)��Э,	|��܌V:@�Y��Y��0=��B�L����D��rL�g�XH<��Ƃ�=��X��@����Hfo�F[!�d> ia���`��tJ�NQ�b��yR�do�,Y�U!l\�dcq��zB#"O�(H��0;�]2q�Q�m�NDX���_?�4�H��:�L�i{f��a!�G�X*�"OyQ�۴[�U����+��%S��Or�=E��M��~]��)�,
��
��^��yR�mZ����,�L��m�5d��y�'m"��B�H���r���$�yrL
V��xp픩+fpK@J���yb$�q8R+ֳ9ŰcGnW��yb�� Z�Iy�"Z406�@g�3�yb$��y����%�
`[C ���y�N^�wDj �&iٺ"�ΙZ��]�yr攅�R�3c��k���DV��yBO�Q�0��L5'���r���$u�h�>E�o�mj��aq���"��C�͌�yrnJ=NlЬ@��8b0��%f��y2�]U^@ySm�
�@�`����yB&�>����4��qyCG��y�M���m*l�5}��D �����xr�0'�u�K��V�A{�
���hU�ē5�y����e�&�h�>��P���L�ᧉI�Jc�S�<K�̈́ȓ<��U�-U�v�^|����D]Ф��\.��QEVxm��J'�p���&�������x"�EF��	аgY<� �Qi��n����0��0�	M�O��I���r���R@3o�J݃"O����h2T�2�`����f�d$*!"O�8��F�+�ݸ3*^�/���q"O����P�J�̲�i��YԨ��B"O�,�ŋ�	r�a)�hݑrV���"OH9�����hʛ?���"O�衢�K�:���&��&��"OƘ���1ir���k�(uC.���"OZ�k�I�#b��9q�C.d����p"O�!pł�4A���j۸�d9��"O����@
.lJ�:�`�"�Q� "O��T��o4~!8��O8_�(���"O`�@e��F���`M�P�����$LOBِ��]9>i����f2N��s�'A����`c��г��)��ҕD%D�X�s�G(���3��
�H$�E�.D�8����l��F�F�qGRH�c.D����ِS��<�h��r:��Pr*&D����;[Sda1NTb����B)D�xk��)4e�rG]6O�tmcD���ԅ�I�K�J�ӱ��N_�ai#���B�I�7��sb$�D����Sk��NB�I5 �h 3��ĕF�h$ϗ!�hC䉃*(�Y)&#K��1 n�8G�C䉒*�1A���*4 8L8b�Wq*BB�	�l���i��� p#:E8����nB�I��Y��DO�_,�RTJ��hB�	<p\�S�a��s��
ƣ e�C�	 ���#@A1�����/d'pC�I X&1!�)؀��ls/V�F�fC�	;Ǌ�1@.ӍDI^P�AA�h�C�ɪd�8O�_� �õ�3i�C�%Y�d ��;���ޒ0�B�?2�\ �~bb�j� Y�P�x�If؟|�Ҧ@�rm�5dN%=�����%�ON�Q6j�Z���"N�,�U��6���ȓe�`8�V%�R��c��N�dF ��'�ў"}�E���b���e�
��@��
e�<A�P&}\@,��c�j��\H#_�'�Q?��Ν!^CPe�I�kD��[��2D����Ɇ"��e�5셛
��ъ�O2D�4"1��*f���5z�����ɵd\!�d�IޤxہU�J` ��T�fS!�$��[Ԥ�KJݏyJ�e��/K,n�!�6�^�����w� ��Α�,�!��R��`PdY��8��nպ9�'���E8�D�s��O�|P�)�!:Bڐb�'w�D�3SBT2R����b���N�!��S�` ��A��n�$="un��!���\�����d������<>!��Z0���W�3�,��D<ONa{��z�	 k��b@�8}��qG!�>B�I�o����� 6&ʨ���� �2➘x���Ny铠X�i˱�:f�����B3r�
��$^~��3'b��`n�"�t5�eg�F>������O>˓ӰQЗ��2��e0�J�lDyB� �S� H��;���\iE����$b��z�D��]�ꌚAm��3b��'���';ўb?�sߴ#�tq���&2������B(W%�i��{B�pӧ3*as,�t^����V�r��#o��:����T�GB(�ȓ+�(�j ���H�0�󃜝\V@��ȓ	P�lQ��
� ��u�g٘���S�? ~	c&�Cy(ΐY�閿(�T��"Ov�"�
ц �zˇ�����"O�M�c(4R0��rJ�H\���"O❚�g�o@��&�|J��[D"Od�t�Ϩ!u��a�ȏv ��"Od8�"��mw���!�E�b�E�T"O<dbQ ��9��4�	�I/T(��"Oԅ�BAU�VȂD� ���U�$�"O�q�d�--
��''@�1L&�Q�"O��*���J_T��cY7H-9q"Ob��F!�8".��ցٴ*����"O��b��W�#�!
��9m�1w"O(l���H�ab�yү_�X/��"OL�
���.P���HM�$*"�au"O�	 A4
d��;UEܒ5���"O�J�L�z�|B��,
��w"O��K��A����c��|Z�S�"OڐXe*��$������'a*��e"O�-��CӛZ?��lʷc](���'�Q����G�&��W�����(� 9}�)��8	`u;�L���`Bc��:dB��V�Wb�0�A�/_w�㞸��	E�Ez��/��q��
S��C�	)Ek�pC
˗:��2���2����'S�8��*R���l�5i�&*0��H>y�A��97f^,,�Z�,��["�̈́� ���aE�f]~�J�B�J)��Zn�k���*4��d
%싚r�쬆�� cDX��>���T�<����.;�u���]�x#�BO�f,2<��):���f�	�PHc%���es��ȓ�.�t�ޓ+���wɰWg+D���NS��P0�0/�D���`<D�4#q+��k7��WO�*��#q�9D�PP�2F�ᢩK>14�`�t/%D�Pf(��촋��լz�����*"D���%L�"�x�L��)l���h%D���p!֨7 ���E/���`&*!D�x�ᏑA�,DZ���"�~8h?D�� O^x� P%���y]�&�=D�D�5�ژ���f�� ns��:�n!D�� �B�l]��׬�#�*+ĥ D�DC���0�� � 0v=��zGd$D�h��&��%��C)N���M"D����*��R����2@����
6D��2G�u��S�J��r,��	1D������%��re��iAL\���"D���JF:	�L�d���2�;D��3�e��3n��+PMI���ՙ��&D�x�蒐T� �;���X�V�X�G%D��wk2V)���b�ł!��i��8D�@�v�V�Gt� ��_�Aq� C�9D�hF#.P�0��$
���N*D�|����:>�`�[c��(\�d 5G)D���um��D,���m�����Rn9D�� i�.W�FJO��2w���aN8D���Y�"!� ��.b�(`���8�y�@�:J�R�2� x�ı�%o!�$12Q:���9�L�{r�	�&�!�$ԫM��0`���-n��AV����!�$��FG��٦��?�A��`N�(�!�Dފo�
�k#�V�½@GOBs�!�Z�%J��Į	Xi�Q+K'5�!�D]1I3��1�.ßM�)bϋ4,m!�� B�[eM�t�����.�t�!a"O.Y�L�yONa�C�+6^d��"On�2ƩV�	°���h_>ގ�y�"O4�PC�8?��ȩq��^�:{�"O���Ǯ��)(�|x")N�!��KE"O@Y1%� :�(���� x�����U�T}�a�w���3�@'z%�a�LN����f$D�l$�$<�F�p#�t��-Q��%D���QF[�x�X���^*+6�}J� D����u'ba8�́�JS�ڢ!"D�X
�G �`	X]�R��s�Q�K"D�����${�j�S��C�(j��"D��R5!��Q��\�4I�~���y��5D�PQ��W>fBd�� &�#�"6D�@���י'�E��.��l�T��	2D���օ�)r�B8�ů��� �4--D�lK�d�t��(�*�2r�b���M(D� �d�<WK2�
�J�?�|�	G$$D�9��BX���W쀳��U�1D�p�!Dɡ�,i�2i^� �,�&'/D���a�؊mՄ"a��:�|ႂE+D�(*�J�˒�Xv̛�ږ��a�/D����Q��|z�LU'SU�q$,D�00C�	#X(�AӬ3��!��+4D�P��G�-�@����
I�M�d�.D�p'^�ʦ H��ف��� ��:D�@ i�zuI��"Dn|�C-D��Q��5)�]

T:_�eP�H=D��8f�9=�%�elXc�^ `!;D��J�n:R���闤W5ie:y�%�8D����e[�$��Iѿ^�"��Ħ+D�8��Z�dq[%c�#�.$;�k(D�$)�G�22��Q��GL*>�`��'D���S��$�P������%%D��&�_�?�PY��n��]��	��G?D��Ӵ�F�"m��n�5p^��AT{���DM\�D�t�'���S�ڏ#m�`
���3�=��'_R�C@"�7'�I�9
�P;�y�m�9�X�E�<���������Zr�n�m=���&"O6�j�f�l�ȂK ,;`Y��ӯum*,�昀-�6-�,I;�?�'
%���;ô�Q���E�x��'�F��b�*6G�1!�M� s�$�S� L�-�P�ZDےA�g)�<԰<�5�I9(��&�̀&3��V��s8�X�3Z7
��X�@[/d�h�HnG7)Ҙ5��,I6,M��Ff�~x�
�'1���k��9n�(�.W���H�0Z�] %�,Y#Aw�p�CM��1��:O��y�6�	Q�G����"O
ac�႓��i��l��X�2 �WQ�P6��H��x��5�C�xyq��Ԃ�Q�8�"B�B��qC��&݂�Z�`*�L1g�޾@-�E{E��q\
��B`��S��7P���G'%��=4f>���A��v̬ jqlJ-g;����I�`���H2.��وcF�cNj(7&%R�8�#G�#���`���qg���M+v�Bm�w�ȣhjj���
I�	U��F��ȸӁ�Q��5�+
��5At��M�b��d��	J�h*`O�(ojB�I�[�-q���s1�t�c͌]��91A��@���Bǃʅ0>���
>��38��'��%�p�F�*�!6(6 ���|��H��بr&���Ůڅr��l	��0b&��B��M,^�aP'��5�F�I��6�0����a�'��<�?���"g�
8(�d�1 �d�@?H������܎8ԍ�0���
(9�"�L�/��5�&�!E�xh������!'�a��@@,,F�I���p �-z�4��'u����V \F(&�	A'_�l�(�ȓB��s4�
7�`��b�;d��Dɿ@,"ӀIy v����W^�}(x�������XU�Vf��csJ_�^�����/�O��h%(�����3GZ������Խ��p`q	�-9|�9qQ�		L�X�k �L��Q��!��f�� "J��n6=��h?��>�S3(ݫI�i�l zkV��� ^���Z�aO�mp��	i�؁l�eK�%	�t؊���ܭ�8E��%���x�'�^ڄA��<$P��5%���A�˄�J�yYH?q�PÎ�@q\}��=	�R�M"D��&�ŬQ
�u � �=���1��l}F�bU ��'��@�M�4v:��ԛ�k͟6t�Ę�gA��S+{�j��B���ү��d�mS�L_2�B	��Q~0 Ѱ���q��qX�ͅv�ס	��I��ÀQT %A�,J�8�h����=�ax"I	�dV��`�Ҍpq�M�5��-�&A&��R����$.�Q�$�S&b0��	j�� ��"�.�"1��R�[���'_,UR��L&����m_�e~J��`��%%[�H�O���[�-L�s!� T�ҰD��=S�'�$�� ��8~
���o�;Ey�&*S�{��S�/�@`�cDQ'm�q���	�(S���./K&tU@�B�7�0�I�A�ph<�5(�d&��C	�'t�@Sb��9e�D�R� �1�D0�Ϸ"�̵��-g4"=�bV-hS��W����v��o�����L�HWrl�Ŗ��ty�`�H�Q�d��ѷ��u���Ӥ���XuMA�O�|���TO]s�`�*��i�0�����'�2p� �A!U@~�"2[� �zhqL��9^y*<j�AرS������,�C�	�}o��ᆪɲ9/�܉�a�2���f^m�� ���acࡃ�l�c?]Иw'%�%�3Al�Ɩ5e��,�
�'�,��p�[0����F`�  ��ÿ!�y�e#�D�He��σ��`�Z4�O��!��OAi�P�BS�+�j��u�'�l���i؟WԦ�q��/}�t=H� �rg�e��84՚'I�'����	�z�P��aC�@y���Sl@M�=��$ެ�f��4���'`�8 ��8K��1\�YI����
\�EK�@��C䉪N"Q�K[�}����`�&a���I��������I�]z�kX(J.A��	�7��b��ܮL pA�,G�m�!򤌗 ��щ��*g�j���ə���Dq�	]KvR�j�mF(?��ݓ@�~J�}�
R�)��i��R,n_�DYda���?�Õ%+Z�,S�`��&vp0!� �ƴ�4���b4�g�İ��&<]�LYUΛ5�X�`�4IV�?�r���ku�p�l��c�6ih�Io��B�*&z6��8���0R��C�@<\O�d�̔�#��	�OyZl�7	T�3�>���-�;PG��Q!��Ģ�5�^)	���#}�V)yUJ5�I�M:%q"��I̓
N<5QbA	i��?�:k��"����4Y�'��-E���(��*���؀nR'� ��qOȼi�"^o]T\ss,ՏDlp$: @L�-���E56�V�X�&�# �b?���H@�3j��$*�]S�1)��+;�,�z��M�T탅E��f]佢�T���i�%
lrĘ��ɘ/k�\���_z��V��_����J9Ch��QХ׊lrج�i٬m�Z��f{Ӹh�C	�?�:�"S�9g'褫��+O��ʐjL32펹��n�,�
�`ce��Y���C�Z
n��$�56��a��y�<�� ��)Lܠi#O�y���_�'D�$���fM(L ��bG��p' E�OB,c��Ǔm�Xl�R�2Pڰ1���3W�f�vnĤ��t�vw�mʰ�M��U�f*�+���I7'Yf}͊�Qo�D�}&�0���i�`鵦��+���3a!H�j��T�f�LZb�����;�,�F�MG�TP6s/:4�1im��v���P�+�Ǘw�x��fB_ l��(E�Ap؞�ĭ�i;`�:F卹����u� 8���֬g\ΰ�P��=�v�	kC�m0z�B��;
����M[yBi��=�i�� M���D)U��O�hz��K06j��R&Rt�d�q�Ρ|�^�8�%�l�&AdS�-�(��I�EUĤ��q��H�#H�<<�Je.2DY��ǲ<���U ��x��ÜL�p����L%�q���T_*�4�O��cŨ
?z� C� Pm�'�e��H���l��ӰD,��.�%+�ʤ0i	�a,-��ҺR�}��X?yp���'�̹�;]V�$Q�سD�ڔ1���	d*0���#_P�Ӳ��t*��=D.��(dB�.
:$<��(Ȧ&��+4b��E-���p�0��HR2����@���5��� IR�D%Y_�z����0Xџph�R5-zA)��5D}�P��S�k���,[�lA �K̚Uߔ�����7x�|V�T�2��e&mӐ���(�{�x">�7E�5NvX4&��#���*�e�Syb�Q__����Q
A�a���L���	><�m�$�r^ɨ���7!҈ZSʇk�,x��f�!@CbM�7�x����!Chp� ũD&�@�˥�+/��(Jt���V�T("iոX�v��� @lt��酃!�V��E*�)+���14A�|�$�P���퍍q�pX��	;���cvJ|�V�J�Jz�S bF�HXp�DW�e���$�Q<'�A���tOh�k�@�Mu
�+ЂߘA�VdW��#.�e8��I�}�$���0|ў�����F@T���k�(uP��͜��Pb��y�m����'��y���C�#�Kˋ>�ؚ4MSL�2ЈFA�|�֠��J���'� ���O�Jj8%�
ch)��4\��E�%�	�$�0qy �#T�u�%i^�Y������b�%$]�X� &ĬA�����P1���R��-gV�Jm������		l.�c���o�9%�ݸX)R��p����U����1U���B�
i(�c�jY�n�
=��w�~�8b�I�@.�(B����EO1C��)VH"�Oy{ ؠ
�0�K� �haU���%�6�r�f�:y����`�Qjƥ0rjB�2gډ�A�n�xy��!�$6��;s�6$C� �.�ļ��L\6Mr@u�B����p�qk ʓ����L4HxTQ�2FH���l��	�ک�(W�Ůy���gP�h�E�˹I�h���[�/يԄ��US�U����Ќ8���Q�x��@��4x��#��	~��G\�V[�y�W �> ߒ�'�P"}���ݱe3�9�2e�Y�)iF�ث �C䉧 ���#���du��I�� a���-*�5bs�YC٠��)J�7��Ԣ�2��Hd�˻O��!�w���X,�*��"�:yh!��*����K�rrn�����1]84��2Kp�)ї`P1�^Eh�Ń�")���'ޑ{)�QM�2X088���M>A�i 
�v���qr���O��c��˙/w��3�մ<���kӄ�W����r��<@A����#�Vü]�t��'��{���k7P�Qu�;|Odlz�n����$_) Ĥ��j�u�ȩ ��˟yM���i�b|J�n݊�����Ğ�ָ��*F�#u͙����b���+\VuR�b�<I^�92�"I����ꆆ*N��y�n��M[4	8�N��e	�>�7BljD��9�X���H=�y�*��|`�t�"غ'y���p��0>�CL��@�%)�<Z/���4B@�S�z7k��n��m���	�O,�ů!u�j���˟_&���d"�=S��0x�(m՜�����_����"�y($H�(Th߈���$�]���	V-z��@�>���!�`C4�̅"TI7Y�Ӌ؟t  y�L�h��lg	
�7���I���fx�����6p���PC+˙P3|qR�'�+0*^�)J�6���c�&aw��B"E�r��(r!���h��8�/�*<ɘIQb�"D��DB�/XZ���ן򄨣�   L%��� >x���ɸ$�ԢH��4:t��P�;� ��`;��D)+M�Mb�Fğ�����>\I+�!�f#����gL>E<��@*����;�b��nt��c�#`�L�����w�L0	�X�L>��'r�}�֦�s���2��Yv�'؂���I��b���1&�\k��f&�t���S;܅ЗG�;

y;�� WF��R�	~}����Q
ZQ-B@�~�h��
�^����k�����I!�,�Y�V 2�ܣ%Q~
8K2��'��9��:@,����{�<�F�V�<A�p� +R"Қ�kUM�\�DV%9B��7j�<�����GH�|�Sd���'Y�m�"B^�< q2���o��)��^JD�6��gV�L��ʃ�`��U�E�e���PV%m�Zi`R������f���VG�� ����EJ�����|F�����%8 ��%�N
 �Ah�;_3 l��@P���
��=Y��1tْ�KW�Qh � ��M8�lk�3&_Z���¹2�$�*��q����H HT=D�!�$�%�@��� 虚f֗:��A.�{��/(x$����h�O���E�H�6�.H���M���|��'�D�Pˈr=�����C��H �ս��0�3O8�!�+O�����84�u"S�Z[� �Vʸ+�^]���~��F$���!� 5��]X$�TUxp:�/˝� h��Y���"g���"�a�3~�&��\�82���E�h��y���'�fɫtE��w���)�Ιd�5s�'.�4���U/q�XX���r�@�J����"f촥��%Ř$Q�}j��Ć5`�\���iN�e�œU�<iU�^7Ͼ����:��|� �U��@��K}2��-'�b?O(��N�i����!դL�0� UO�L�"� 5.P��#�3\Q�� ').� H�b�X���|Z){�d�#�.��4�Y�Uw���AB��p:��Jj}R����H@
ǃ"E����S��y�*��;��%G��I4�ɹ�h����'���H��<H·+��D���R#�0�9��"ONTqG��>�4�T���=���"O�D��[c�)`��>���Q�"On����%4�^� ���b�؀�""O,@B�O�#q�H��f�Z�m��A�p"OnT��⚳O9����A��ZGB�{�"O���sMW ,6�"��#k��<s"O
Ib��0�\�!nĴS+n[�"O�]�#�K���ȍ�y�"O����U =�hA�FOq�Na�"O8��B�$ �f]��Ӻi2l""OfeА������!`���L��"O���Ă0u¸���p�u/^�2�!�ĕ=U��a�P��|�f.]�`�!�}v\��7�X� w��E"ƭa�!򤉃]G.����\�cl�ФO��C�!�� ���k�7hr�b#D�|�z��'"O������k�,���5h��t��"OLd�IR�1Z@#��Ƃ&��A)�"O��8��4Y��ҁܡJ��� a"O`@�g�؋tU����4su�ً"O�Au	@Z+.��F�E'	�d��"O~�1��$�Qqs�C
4��b"O�L��)�4�U�7��3F�%8�"OL��.D���9!v�H&rqč٦"O�HȔ�å'N|�r���0p���"O����KGJ9��Z�����PX�"O�²e�} ��s2�_�;�
-��"Ox�XG��5i�VT�Y�`�H9*�"O�q� �үV:���3F["S�^|�s"O"��-88䭠R��6XҐ(�"O��P��~�Fe�%��`�J�a�"O8p���.!㤘��	<z�|�"O���?h&�D�$	�j�İ�0"O�,zRB�*���QЂ��;���A5"O���O8�F���+P �X(ҵ"O> BL�~�I�7�1Pa��Ɇ"O�*b�A6P�䡲�dN�0x9{�"O �)�nb���8޼��"O��C��J�$n�z�Ȉ��=A$"Of]�Ao��s�PD�`�U���*�"O���q`W�M��Z�C�/2�le�b"O��h�	�4�,����PP�Q!"Ob5+\�h2g��e>}##�r!�D�>��,W�=Q@��Q�կZ!�D� m@x�zǅ�+Kތ0��)<!�Z��|H3��B1
�L�+�
!�V�3�2��V�4nŦ92$^;�!��9��Ju�����qBNݨq)!�d��=��墤�q��LQ6-Y�t!��xC�M:������@g�S�H!���>OZh��F)L��LjG\9'�!�8/���F,a��A�`J�|�!�!_�lX!eS�T���#/��>�!�־s��	��
]�Q�O�!��IG�ݛ֮Ȝ=��y��)k�z"G�v�*�RPj��Lr�-�d>���k$���)��9D�q��< ���l/)q%�4扯 *ʕQe!ԑ&��#~��� h���ĥ@9*���S0��o�<a[��NKr��9��sbΑ� ����iD�%�E�۴sM�-"��L����M�o�Љ(҃�kd�ϐx�-���pȘ���1LL=[�,�5:BN(�a�G
���)�DԲW�$T�˓�K6�ܨXv��ٲJ߄��؆�r�n�Y�G��y|��+�E�X�(����E�.iS��ʛ?��K3	���Px��U:4҆Mۥ'�c�Jl�w�K#��	�7�6��&��C���
��1j���{S�؞r^����C�\����V���b�!�X5� DO3T|��VD8�R�#��D��u!��l�L�����\�a'剕�4y�T�UHP��ʻ��C�I�N�-����j?t-��`�(i��QM��a�<��0���2&��W��?�*Z��4-��Inx�-�ƥRr8�0���6#��IG [L�p���%�m�xC��U�����`ڑN�@u��!�Op��C�B�}rf�٦9� �ҙ� �2Ix�=�D�0/bT��� L�$4'?���! 5NI��!G@#��ܨT'/D��qS/�?02�r�ª:=�8��Қ0���{�� � �>���C�$2��(���ÏayB�ȑ� )�u*ͻ)�������?�rj�(�k��6c�x��RE�#T�:����?@?dUKfl�)ZzEK�"џ�J���JO&A91��(Ɓ/��J&!Ѵe�YE>r�Bل9��p�'�k`�p#SB�?]Є �̀#+�1�&�'�Đ�ө��b"X�S���b_�M�,O��P�o@���A����6+�H�w�يU���H|R�JJ�[�0ՈP�=��V��J�<� �C�IO�F�r����k��4;�K�c����V���X�F�ΰ�O��x�&0�~�@��57�`����m9��i&��2��?��Z112��ЧS�-	@v-0I\T<���B,	r$١!"P�c؜5�tıO:(�F}��?g�I��Z�S|ƈZ1�D��O�5kT�޽nRP�aӊ;Z��0oX3[,"erTaR,�@ ���{���U��'E�~��8:�����m0$���S!�����6ǂ$02/�;�	C�nO�2�E��	'����C�扥q��$15Ƒ/�ʥ�ȓa��P�,O��Q9��O+}�8a&�у
*N��H��Dw戲G�S�SB|���겟h�v��$ݪ�+�!$sR�w%�ORd�jø&GŇ�wX=Y�^��b� "w[b�_���s"ϭl�����J�I����� �m|�Ta!A+y�ax2�%>XE��ˈuF�K�'8��M6j�=���"�02�C���c�~$��	�]�Vл�j��K=ĸ3���O��'�|�A�@�M��)`+��Bq���Ft"8�O�\�����)J+�l3`�	�'�b�� ܗ=����d�/G4�7H�+{�Q���G ��BD��}�q��t�A��S����,�e�|(`H�P��C�I
6Tnh�g����0�O�k��9s�Fx]NNO1j��LҦ�@�7Pbt���� @�+	6g�Ȳ��S����Dۃ1mj�C�ɉ��4y��$�<;T/�2]:��p�S�4�+�j�1@�J�"�|�֠��C�t�R}�t! c�m�=� �ΰx�:���&�M��[E�
�	��G؟Zi�b�! d�Ѓ89b�h��"O��'�iKP��D�k�(���[!m}���&dĊL�P��J ?�����N��{�(�U�4$�x����Z�<�L#zD�٥�1U��B������,r�Ĝ^�4������x@������wD��C`\ Q�L]�gdJ���>�WĊ�0)qEL4�6�R#*�M�AM�gE�iӠ$� i�8��b�f\�ۓ �5��N�[7j��DG^Y�J9D{�@@uJ0��"f�+2�ɧ�9Q`�;)C�5��ȋ;�l ���p���Bv�p�C��rx�/�	*?���=GU�1lFb�|��"��G�h�c�0Q�z�u��L=��k�b �`J>C�I�3F���b2pn$*4b��3G>�B��.Z0wa�#A+��P�2�$���=��YaT�� ��҅�v}a��@|�	8�L]�wN��#�_�x�,AT!KU��9�A��:�%�ۓ�X ���G�d��Ă�3��G��˅q��QNӈ<$�H&.��Ӓ�۝o��=B�N5�h�Q��u���m�;[3D�H4��s��o�Hu��瑲NJ�'X��EM�@�A�L�z�ZEE��DB�>xt�D��0o����U#��'������O "zuG�,/��]rj�@�~��gI�Qz|Ẳ�ݤv���(d	�)y�n�%?� k5J)Z�͋�l��N�6!
�ʐ�U�N�ڀ�X�����doS���~ʴ���@�P�R�MG�r��dL�+�RL��KP8u�b8�A@ƹL�ʨ�@�'n̐�FM�,J$��@)�@�����8j��BAĳr�4�2�T�z��ݠ�M -Jcw�/�X���.�ͦ�����nt��f
<&���׎�o8�(����-�^� fJ�:}��<r�A�u�H�S�&򰸡a(F��kGM�9FT�@YB�K��l�X�K�1w��˔��OI|�u�>T�tYK�e�$=�ՓL���n�
Lq2�)H�#�����\�h�ԇ�2{���S�����N�'c�0 ���!a*0���*��DX�?c��L>�2�_�X�V5+m0����ԅ,�yh ���hazq�b��]�JM�R@������=���Xc�,����ԡC�ty�l����� Ŏ_�F4(W'��=���])b0jqB��Jy*c/`�@&�֦7�Ha�A�U%G6-iFbW�a9|E:-��X]b�!���$�6A�l�C5r��ą.�џ���_�f�	7O���Hcw�ѽt��0��mǦss����FG���!�jI j�n@rG����=�S 9K�xf�P8�>pKg�hyb�ٰ@�  ��\�H��Q��@8�%K� 1	��E�D����c`�џj�I���K�\���2"Ol#�[+d<=�� �����(7*W�e���:� �?��!��r�~�H�~b���^�v�s�w�(q`�:vQ.d�R��3IT��#�C�49���U�#e�����Ϩu��<s�
�4d�� �Q��z��2�j�Q��Us�j�O�]�W+�~�K���q5��"JА�d�;��O(�s4��N}�PP���<�8�z�'C?"�D�Ԅ'0�46͟�	��pT���LI\i@b��Ӧ�[Eaң�`xF|�\+CC��� ��60P�1��L5����]�b�(�&ݽ5�tqgj"+*��U�Əj��3��r��qC�@ 斞4"�����"m����Ңv���d�~��=(gAJ�.��Ya��34\��7/� t�H��aM����+Cř}��=0k�hX��:&���̻�<881� Q+��)����D��Ʉ
�2�@%���� hYCv֑8���
VfLQQ���Ed�]�1��m�������Ј��Dyȭ@-��?Q�j݃00ё���zLh��|�'���'�VX�A�A��ʕ" F!O��鈖OՒB7�U1`<M�j�$h[n�F14�[�����χ�H���=� ���E��F�\�p$��� CS�|r Ó7�j��M&3Ai�LP$�$(!���g"����=2�Th���G����O�M�������S#J�h�cǊ�q��Q>~B�a��,��b�h��Y�rw
ћ���M���2� �g���yǇ�}E�q���g�)̻S�(l�@�%Nl��e��j����R� t���q����S��w9j�kF%�jčb�JH�:ب#ǿa]���faݪu�����4t�h��,K�yr�9ټ���*ӄw�B g�S,�p<�fj׫O�92q�\<J��%}Te��F�!rf��	�FF��-Q��\`4j��Blf���=a�,B���lS #lKp�'۠ Ƙ��� ���C�K�7k\8x�l��r|���'��4Rэ�K� �*^m!�D ���֋Y�u0�)2��ڹ1TN�!r��b���!��Y�$���kå�#���pU+�j��[2 �5Ĵ�ºB�V��%(D�����ʞK��]��EŖ}<�"�EF�mB�̑��]OZF@��ЪDVz�Ɋ�J��M�?!���?$b�*r��L�
�YIx���Y'f(�K �>>v�֫@'>�YX��m����V�h�T`
ߓg�<}�b�_R?��*g�w#�uD{Y(Lآ|�G�Ռ:��e�u��w���;3x�xc�&���2�Q 1>]�ȓ\�jI��=9����@� D[��ϓuk�)��ܟ�98De�=X�d	i��?�'�ֹ&aսC�=�Um^A��ȓ	2aHAl��$�	�P!?C?ެ�a����bZ�A�pn�#dL�O�㞼v��'g�&����ÎKʞ9��l.�O��asl�*oH�3��H�h5�M�*'��]`�E�dD�`����*Հ��d^�4�8 ���%.Hɦ��$�џ(�D�a�
D���Z�<`�l�WfͲ6�l�&lF��T5��D����ȓ[�� (C�Pe���]�qؤO�\�5�928�ȡ�P�c F�Ħ�K̢@�`+Q_����iS%�y`X!沀��E��Q2B���)��NJ�-4�l��8LH����|�T�sM)3�&:4E�uXQ�ӎ�Px"�Z��iZ�@� �A@��9qD	j�.1���U�"| ��'r�pBA��tM8�)�K�`�	�@V�)����'3�4!ۥ�D�.� D��:��1
�L�
�ʤ��$ D��[4놃n�z���/Q'/h�E�?}B��#MW�,s�*��|�v�X�>�'Q�2<xbB
t95z�,���ȓ>n�)
p��8��e
O�#����Y o֔��o~��B��Y����g�N �GH-����/+9��`�@#�� חdO(�� C-�lQ���0NhA1&�/4�"	ۓ3	��9b��C�0� �I�_2\��	=ld(���; �\`�0��Ot�3@O�"C�2�ɔ�>�ѩs"O� �anW	%s�K樋eST8���>��������	ڑc6��F�DM�ds�H�HGC/�)2�٥�y��V��QYT뙗=S�y:���\�b89u��G�󤟦������L>��L��	}�Ԅ���� �v(<q�[TM��
=j�t��ǤP�^\� Ŕ�S����a�g��0;���~�P0s�мU�0�A�L"O��30�MF�@�������2W�Nu�p/�1A� ��M+�yb��9hB):s�C�;P��y�/(��s�4�c �T��L0'-�'��<y�C�)2ܽA���8�T��ȓ �Ա�j�F\�5L�y3����P��'�q� /;�3��#,�
]�'%�G0^���c	*z{��$/�X8!�J<y|�`ŋw���җH��Ћ7�'�5��� �q( �0h$S7
5�
ӓ9U8t�R)���>߶�З�d��MU�S)�0C�'bq�(jR�	r	�]sC �-L㞼)����>�*U�0]�`� ᫃�)`�q�v�H\�<A��]�")�̕>�v}[���[�<�K�.(v�Xs���
5�Z�@�\�<�e��C�V�b��H���7g�Y�<���E��r����A-�X2w�EU�<��I�Xf0�)r ��~G�As��t�<Q�`���8 ��)�E91TM�<!��W��­K���r�va���O�<q�,6q� 9)b��`��*�jJ�<ԩ4/zY�S $p�d�`@ Qx�<�+�R<>e�ƨ�˚�8�$X�<�vȚ2KΜ������Lȶ�_�<� ��0D�ܞg� �y��,P�	�"OhҠ�K/C�@!��G�Hq8"O΍�"��Ak�}eGʛ;�( �"O��
W���.�Z��Ӟ�Vd2%"O��c� +垭��Cx�@���"O������E�ƹ��A�H��tR�"O��{�I�;�H��@�I� ;�"OT��� ��]���9 [��h��"Olȃd#��#�|\x"�>N���"O���BÊ" ��׋Q�#��-�'"O��!�¨:�9�ㅉX����"O�ي����:h ���6���q�"O�%K #�.r;@�c#�L�h�p�"O����V�"�~�1�2|�T,
q�N�j�t=X"̇��%�Gh�by�@�p�O�r� @/L�|��V1p��d�1Ǌb��ʔ�>~Zb��ȟp�����-��K��8�b"W��M��'������*'�>�}""�٬	��9xĚj���J�D�Hy��]�j����5���Sӈ0�0��9��_Б���O�4� �����O��}�V�Y�@�&	�SGŢW�>����q�M�:tV(�'��\�>YH�#�aHnh)��Û@Fx���T;��T��Oț�0|�DNJ"U6�=[��� cg�0N��z�:M�掠�0|��nب[꒺r-�}��%�qy�NI(K�ȱ �!�$�?Mٴn�T=��BܧkG"|ǆ:"��)��3|,�y�f��qm��+��O�Ḑg>P`���chj�:�DR�oNЙ��@�v�Q1���M֧0|�O�u8V��uD��:�V�wB��8��R�C�_F��=KF�����"|b�ĝ�c��ؓA6�&ԳB�Ú&M�]2�_��@�J�j�|J~�E,k�D���:v�JE`'̚T�I�u�T���n8�)�<L��E�Rl��0��}R`�@�,��	b�����B�)�'�r�`r"�&�d�Y�	Խ~�,o�ML�
�D6�)�uF1�Ɋ�\� �"�?y�� �vN��|�u�J2@/`��'><��铏sG�Q[e�eY!B�4{|���|2b���M��~����J��᠂I�C�3qm~�dE*&�`v�:�#�'�E�����zrjP��!�C;����'�(��7��Mɧh��p`gls0D(0�Ϸ #���\�6p4t��4�ē�0|�����rJZ�lL!�c����ܐRƇ�Z �Tb�|b#�Ǖ2�ui<k+����)6#|OT(��?O�?Y���(o`h*F�p�\l W�_a?	��i�`0�'�ms[r��&���>Q�J��h�:�r���A�f p PQ�<�ceϿj�JI9qF�u%�l���c�<I��ٴ-��%02�|ƺA��Jy�<Q��z.H�ۥ��<V)�A1w�x�<	eA��#��8Xbe�K@,iy�"�w�<i�ʐ�0T ⪃5;�D��n�|�<��)��n����l�0`�<����x�<���HVH��.�)uTy����t�<�%%�ri�3f��0欢E��e�<15�S������ɉ���beɒl�<af���9�7C��#P1S��~�<����n�%R�	m9��E��_�<ѴkOpĠ%�R�L�F��l�� �U�<�S�ƨj�" ����j�i�"�)D����u��e,H9R�U���(D��C�IC>+��dB%�?T�D��am,D���5H��YE�%/I6}�c�*D��
V303P$���� *���	w�+D�X7)��~ �d![(8B�)G�(D�\�����g^^��Z~�i-&D��3�@IR6yjwc�=p�p�c��9D�( w���_��h�uY����g4D��kp��!4�J05j �\0�AsW�&D�8ڃ�ڑ~Vh��[���xE�/D��"��$ ���l�Jn��#3D������=|MZ�1B��%�2ᒁ>D��"	Ŭ���q��0 �H�8�H<D�� �u��	�* +�����*���"O��K1�S"���suǀ�X��qiE"Ozd�nVv� ���k��H��"OP�2��_�E���f�]��`��F"O��w��;8>8�P�����zb"Ob�sWm�$b�L�3���<���"�"OXA��V�Ih&���h�!
���"O@%���2S3��h��_zL1�"O�Er%F]�d����f��%��"Ox���+G/
�tEE0{@\S�"O�9۶�
@���T�U�|`^\hT"Onq�t,B+hyh��V#�`{r���"O�9�B�M�6�p!@@LV��"O��9%��$+��X� �^	G`�q�"O�!�猐2�����ߓ`B"1x"O��˱/�#*��2���;!X��f"O�܁���*�y�fO�y��"O���ҪP�"��&�
e�s"O���+�1�0SJ\"r<<D�"O�tSr���7�$҉ҍ�4�	�"O�M�!�ٻ��x�3B�%
9p"O.�2%J�kHj0�'�5,��"O��{�׈d�p��V�R�*$"Ot1A�m835��J#�Ub؆e�e"O�]0�✱&
�3s�[�Q��,s�"O��Pw���a�(CK!o�T�v"O�  t[8���qM%o� Ȃb"O&��r�Ý .�cu
;_z�H�a"O̜ҡ�~�u�b�Oy�$��"OLp�$F'W�ڌ���=����"OVL���Ar�(���B�80P�5"O���r��r� 2c��*u`�3B"O�xk@��vq� �&q��@"OV,��L�D�H��¬i����"O"8�L�|iT5�P.P��>�ç"O6 :�$D<z�8�k�&:$���W"O�a*
�{��h�`�D.y�*@[�"O�[���|�
P���Ŧ }-h�"O��a�eU����j�$@�N�g"Oh1��88��}sE
�#z��"ONіoV�j�X��T�v]�Qk�"O��r*�/k����cM�b<Ij�"Oġ��oí�� R�C/!LP�9�"O��4 
�E,���zg|%V"OP	P��k�04V�K�&M��A"O�����P2_eɨbj�2vI�d��"O���IC)?�� �&�71��q�p"O���!��k>���ʞ,�\`U"O�r(ڞ)�8�$�B:
�I�"Oz�X�E����Iۗ@�9�"O�����!.�*4!��Bo�8�˳"O�mÂ�'���2* ��>�q"O�K4l��tU.����._ ���%"O&���*
���
���"OP�����RO|t! �X|� "O��� O$j Q�%�v�HQ�"Oa1�cZ>L��Y�V�� ��R"O��_����E%R�HA�'qށANw	 \�靾r����'�����,Cm���@�c��9Z�'7ؽh�K��a�8Q�DX2�k�'g���d��Y����3nѷ�pP#�'��U�D�
�G$pڑ�[�H�J�'�bp��U�w��5��-��1Nz�C
��� t ��F�#3��IL]�Z]bU"Oʁ�@����� �@@�Cg"O`E��,٣b4�,��A	�/��ɫ"O,�A�H!i���w�-A����"O~��PJ��A�؀��`�5l��5��"O�I�ס�.M�� �/��*��v"O��A���2Ą%	����(q��x2"O���^%c���ۋ)o^��"O�qae��k'�s2O\�,`��F"O���Q��V��$EkP5��"O��)d��N*���'�L�wK6� r"O�5����F	��sC�~M����"O@ ��)�� ��seH
F@�3�"O���3G�!���
P�S1Ux0"Ov��g�+D7t�#���0���"O�隡�&mx���7i��(�"O����!��m�d�u�[�W��"ONX(4N�h��y��͍�u��H�"O���5<��kM�!���8""OĹZ��Ӗx%�%�!N��r��%��"O��;�B��d�0X0��^���Q�"O~刷L]9,nt���M�XTѡe"O��s�ς!��]y��m��(y�"Ox���6v/�kgaC>0ځ�F"O�4�
��b�Ȃ	^
�P��"O�)���OG�m�U
O�g�^�9G"O��*F'0L�8�2
�h�X�6"O����R�����cAf��d��"O>������F�a3bH�5�8�g"Ot�a��'��<��ٗu�j�e"OJ|�FB�5;3��rs#Շp��·"Od����KL����{w��+v"O
H���1G\�@E�0Y��hE"O�\�d��tw�0S����5j�"O��R��Μ*�.�Y���z{ة�Q"Oz`@��<p��t`'�$bvM{`"O��W��G�ta4���.�,��"OJ�*Q�J���� ^�G�H�C�"O>e�1�Ii��3���T����"O�IQ˘�--�g��4j#"O��W�¢0 �2��
i�:��R"O��� J(e8b� |X-�p"O��7�]��0�H�~���*�"O������?�.�1e�0���"O�q�#Jސt=���C ;��@��"O���l�%q30!�sdLD���+�"O,�z�$�$]�\`z�ȃ|�n܉�"O�P�i!`RZPu�I�n�nP�U"O�����ЏJp�@���o�Z�Q�"O�r��^�VCP��u�W"|��4"O-�%,�]�J؃�%K�	�:�"OpV��xH`���Lra��jS�@�<�D�f��� F�?�B�z�JR�<�����-�0�v]�=��'�V�<1����u��|�,�E�T��J�<��0h\�c�+P��ŉ�C�<��$�WD	B��ET��w��W�<9Q�!ȼ�U��$gc�Cqg]y�<�h��:]h)�B)$"���#�%�x�<���P����K��P�Bi�<90Ȉ�"kDI�ŢOC��y��B�<��c U̚tqD� �0�M��N�y�<��ANq�����9 (Y\�<9@�ǚ0�6a;�耰T�|�@t#BC�<� ����� &� ���#X�(�"Oڬz��>��U��J<R�NTPp"O�Lس���@B�8� �2g��ճ�"Ov�K���`_|�@U/�e���$"O�0"3ꋹc�4,�Ʈ�(m�t��"Ot+�i���R�q0N��D�"O^1���'LV�j�̙�N�t�0"O�9J�n@8�F(;b�ڑ/|��"OrX*5�Z�v���_���i: "O�8�\~�t�d�NҠH��"O�yq�C�azr�1���2��	��"OL���J�Z��1hd�	E�� x�"O��*�eC�S.�8f�^1��b�"O^eo�8e�f���O�#�C"O q�� cR0�o�,YCE"O��q��U=Fg�y!B�W�]"9��"O~�c�H�Z��(�WMƹq+�Lja"O�=�w�+���`�l�]4�
�"O�g�b2�C�hXU,~H��"O9�5�X� `BaQ< �My�'qf�BT�A�A7��B�Ϋ	�
�'��Z���FѾ����R�Fѹ
�'-� �v�­u]��䎜&y�<��'��bcD�= ��	�y��:�'�`D���A�X����%=���' R\!��454�jq���;��%A
�'q���ʂA-�`��H.(�yR	�'.��$�JX8�Q�g�Y�6>���'=7'Ր)U峑�χ>O�L��'0� W�<�ư[��`H�]x�<�%mA[��؇�Yi�1�w@�i�<I"��1X�M�SB��w�Np�<Q��2o���r,��LE0̱���C�<� 7zQ���ȇ��q��}�<�sRYl �+
.��a��D�y�<&���nL\��pDEC$by�G%�q�<鱉L:��(W怍����0FFf�<��ş �lH�����5��H�<�%$�6���3v*ӭP<-c�JH�<�7���@]�`��,m"�9``	�D�<��\�I6���
ν��a!��}�<ٕ�Њ%�1�O�X��4�D�Bx�<����<�~�:@��VL�'�x�<)%C�    ��     U  �  :   �+  7  �@  �K  |V  a  ]i  ct  �  ��  z�   �  a�  ��  �  )�  j�  ��  �  :�  ��  ��  �  ]�  ��  ��  4�  ~�  ��  ?  ] � =! )( j. �4 �6  Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�� |d��"O
`�(�;���8���-0��1%"Oj4��ND^[��"3/9�0|H�"OB���H��*�ʞRy=a"O�味V�!X��!&F�:J�$���"O,��a
���C�Ą�M�"O,$3%o�-���p���+Ն�:1"O��ݢ1����`���y14]2��i�<�6��{_���c�H�`�fX�$Kn�<��A̼VI�xR[�)�Ć�pඤ�ȓA5��('nߡ4�� �)˩%� ���,��r�؊b#`T�eT09���ȓ!�b��g��}�8�F��-? �ȓ
K|m�ș�VṔ���2�%�ȓ"R�X�j�4JN�1�˘X�i����̹	_�jZ��1!g��zܶ��ȓgil,*�J�
j�Ne��i�J%b���f	�(U��:���G��$Y^م�~r�� S�%T"���k\�jx�ȓ|4�1�îJb��@ӵ�ݩn�V��/[`�"�v4�R�!ʎ<��M�ȓ`:��z�ؚh�J�Z��$HY:	��H��p�m�C1��!��B:��0��EnjZA V;9����J[
2���	��4'J�EA�IVW&��~�(aZ��ӹ�>� o�Y�|�ȓ�f�A�
Ο7�H��M�$�����mޠP����/���ANXo*�ȓTv�����{ ��-7�*h��I��sB�8�8���3����ȓNe*M�悡;������X�o��!�ȓ'lj�#F�m�+R&;�|��2)n�C��0S4���T:
b���:�0!��e֊��)��ͷV��,�ȓ0�&�8#���� ع�L�����;�P�AFd���,w�6d��r�EQ�( �gVlɦ�M,H��,DP���|�I	$G#\���ȓ"�)���E�B	yt&B�^�LɅ��wyr*\(u�@ UV$ED02�-Ə�M���sӀŃ��L%'�r|�f��52���5"O���BO�876A�%x�`J&"O��@��~�nW�8\0H�teE�<A/�6r^�=��OA1 D�k#AX�<�A6I�P�j��B�0�SJ]�<�t"�>{D$1�dȫK���b���bh<����d�n4�s�C6P�NT�T�E��y"�')��m�):T$X��䔗:,.mi��${��E��$�@�Xe��_�F�:#�_�yB"�	s�9�1䗿E����A���y�	Ǌ"�
!�حNn:tbqa��yr��ZCpܪ��Csld���W���=!�yb%�.��m����=1���*��yb�խD?fd	$HZ���h�E�a�\QEy��9O6y�D� CqX8!��A=	z�!#"O4l���	�/��]����n��DI�"O@��B^XX��V�m(=h��$�yҹi)�c���SJ�ODIi���.h�xsQ��E��B��~B�@���!���D4a��������(�xźgȒ�i�2I��cD,cĸiQ"Oиc`�A�*HV!���A7VԌ	��|��'K��*ͦ���"����� �m��	�վ��1EʓH�̒Q:O���d�w��� �D��(4z1ڴM��IZ8��$��Q&�,��P�$F-@�h(��j,D��Q�nE 7���F!Q�	�Z<���<�'/�{r� "�li4��*:��$�����p<aM<灵��Y2��
�d ըP[KF� �hO�S4U���a���?��;���P�C�;��$�RI�&"i�<�g��E��C�I!f���"��5I�d�ɋ `���hOQ>��I�}L�� Q���ը�O�B�I�E��+��I3|�b�nJ�1�P����p?����<8j�y�Hύp���Ɏg�<Q��KX�� 4/�$H��-�4.�a�<9��\�\�� S	�
t���`�Z�<qg��Z�����-<�@��Sܓ��=��$�FHUPơ�'Fa4-r��N��4oZ~)�f�΀.ל�rመ�wt��Ө����>��OH��<��L��Z<Pv�@���i���	
�a�m ���0	�xⶃaA!�dV=�=zv�ܼ(\a`�ۄ
,�	��HOQ>�PQ@Ъ��83Ff���*��$�IQ���'DŚagjP�a��:5���e��-�ȓC9�=a��ˈ.~��j�/��l�& ��Q9�-���
���Ĕ�T�l�ȓb�zT U�R�h�>X��O!\P��@���@����t��l`)ϨV߼����6�H�'t�i�#L�(���I�4C�^��.��S�O6�=a���6�`������?O��=���OyBK
/���@��$��t���O�x�3�'��v�i��x���<&æ�B�O'<����en�����؟��.�S��mܲ1�Y��悽9&�H#@��,+���Л#Ы�,֛F��"7�J;�!�آ@Ӕa�q��@L�K��P�!�d�Ȁ�[p�[�X�4����B��I��0?Q���rA�u�u`K�L��ܣ�m�h����'
j �S��}
 ���ć<sʞQH�'{�m��ꁨ%�v@i�m�Z,b��$ғ��)�O���?Bl	�p4�)x��2M1�tєǙmy��')����h0aCx����4.���Ì�dؖ�?����'�)!��T�n���N4(�2�럴�'S�OTi�礂�p,&0�	��	4����'����'�t�`����{�O7|~��;�O,�=E�T�I5O�r�2�H�r\�Pր26X�'���0,Or��e�_�<�����M�6���O��Ig�Ӻs���2��q �%�m��� 4�D&"9 -��P��\y�郂]�$:iY&1M���	f�T�d�����+�X�i�G�k)xyD}���)1���0�6{ؤ���(B��4%n0mS`��y�*��+"�D{J?�YU�Q M��yB.�a�*,��?D��`�2��ti�n� f�T�cq�>�y��O�f�ehG�~�q���=x���z��6-Bg��r�eܲ�r��E���r�ў���ɂ9,����0Bl�{uf8$��=�N<����8}���i��$M��٥���y" ��nD.���/��@��u��Ѧ��<��o�>+OV9��O�"�(���Aļ �v]��"O�̱6
H�W��)Q� �<9i�4Se"Ozl�1L"e�0�ڀKVj=`�'��d��d'8�!�3�!9�c@�(�}♟\��� 'pn���M�)'�<��W�/ړ��'���rB��b�F�ج
r'+,I��'�a}g��1�ŏ��(�&Ya�K;�?щ�4�8��'?��j'ҸP�ƻ�f4�Q�� iX�#=��S�? �PХEׅK�|�A��ԊQnm�Л|��)�ӨZ`>���ܽ|��U��_�C�I2�F1�$�ʤR��%�s/6�<u1
�'&�Ј���#�>d��g� _�D����O����S�Q��)e�9x�h���"O@�ц�Y��b�
�.�0u*��'UV��R�#���L�6L@��n5��"$D�`ZB+��N<Uk�)�VYc�<�ٴ�p>ѷn�@684��]c뒡���$��d9b�Q+Z ذ����,u���/i����򄏄���-�'�x,�KӈF��\�c��bӬ��	���:�:�	Y|�XP�n���Ę⁅(XN���'0	�!� X�H9C��.5��=�I��F{r�x̓!��-Z��Q ���DJ�X�̉�ȓk������$0�.	2�ŏ���u�'oB�i�1O��g�ɫi�,�7�E�E����&�������O��	T�� ����G)VR��碇;�M��'>�E�tK�1_�̹��W"
��F
��<��4ø'�V��AFH9�F�	�CsD�@r�y��'�X�
��6|M~���`N�c�T����4�S��m�=�,�qrڣ:F��uÕ�y�I�'�	iZ�������eKI��D{��$��9��DU*M�g�Y��*���yr�� 2�x�&���6��s� ���f��a��_��3�h��5kL�ȓ RdA���(��HAqB�֘��ȓT|�[ !��#�xiuݏ"J!�ȓWٸѰ ��X�����1����'�~}˕�%zeI����)�͇�=���� N �����pt�9�ȓrV2�`!͵M^6��ckݦƶ��ȓ��Jd�=oA�В��RU���'kP SMȸrւ���S�F�����>���-	�H�K�r��ąȓ�@h	�ŊC6�xSՇ�/�佅�*���*W����)��F���ȓt�ta���P�d�t�iŪ�\zH���{ FH	Q7�8yr�҇@�����XqF��<A���б����8�ȓ}T��e��
 *�����	LpdՅȓȈh���I'����L�=?�����*"�%��=.I*��?��9	�
�<��Lö���y }��w�L��1��8,�Yb�� e@U��9�@X�䚫Y��9Z�hO�i�j���*m�!�1�ͯp����W��F܈�ȓ_�\���ݤba��H���3r���n�X��6Jڽ�� 
�L0����5�hG�L}s������i\�Q�ȓ$zD���'�7ae�L�b��S��e�ȓ.�	��c��d�x� )���i��_c�*� �=���E�ŗf܄�4Ԕ����[�(��2��%nT=�ȓ���P����x_�!�	Mr��ȓ,�uc4�]�#֌��E�Ȟ+���ȓ92�I[�D�X�i��%t��L��K)n5
�)T(|SJ�r�J� n�rͅ�k3t��&և!�l�J�E�vi��ȓ)�~1��?Sq<�Z0�֘~7�p��;�}�Vi�<TW�6�LXo^��ȓ:̽1�Aϋe%�aQ��y`�ȓB)���g�<G`� eͼe����3�xtS�	�5Vd�]Ф��-�"q�����p����0����)�+|�$d��S�? �Mqg�;7�r����K8%����4"O��%&4�0����h����"OXLjgk :"��sJ��Z�v�a�"OD,��'S�#ԴT�Čc�Ό��"OLٹw!�r��� LVoӒ�:��'5�X�X��������I������&��;Ej>��E�Cx���	���	�������X����h�Iן���4<h.v2����,i���5@S�����͟��IΟ`�I�����������$J�ٱec4� dC�%q���ɟL���l�	��������	���I̟\�Ǡ�kC(t���A&���X�u������ğ���� �	՟\��ܟh���L���2�/�%��*��V &�2����0����x��ʟ��Iß��I��X�	,�x(�Vd ����ZZJh�I����	�����ڟ���ڟ8������ɶG�њ��_9{C�@� ��F~�u���`��@��˟���ß��	ß��	c���z@���.�	���I,>YBP��˟���՟��Iş��I�(��˟|�I)46��"�	t�Q��!	�B���ԟl�IƟ��I՟D��ş��ß��	*r��|j�O��8�D����H��͟��	˟����ҟ��Iɟ���RN���!&Ϟ,4\$��KLr���ʟ�	��d�I������ҟt�I/c���*Ԃ�4^ͻ�H�D�8�	ڟ��	�@�I����0�ڴ�?y�Uf�ܚ�?n���Q�ӗ'���wV���	ay���O�Ll��#�'�o���0C��q��=I�E1?�R�i��|��~��i�8 ��̅�l}�/��0���cӲ��Xb��5r$��sa
Y��kԛ~r$KX3�)$���vl�y�`�k��?q)O΢}b�gĿ:|P����0U]�uAEb��,>�VA���'m񟮝nzީHg-�"��9��OU0{���0ҁ�
�?!ڴ�yB_���I�b����F�:h0Ő0�0Z�<2��Ƽ��dPa4P�����z8j�=ͧ�?�G�	ce�)3Ѡ�� )
F�<9.O�O�l����c�p
 L9��0
��Z;:i�eBg��2���ܟtl��<��O:��F&ֱc��a���1"1�ŕ��S�#��0��b�(!�Ӕ3�PB�+ǟH;5͉�[��(㄄?b�{���ty�\���)��<����dR(���DM ,&�۶ ��<�W�i�H��ON�lZ��|R�a�F�f�0�eɹi�`h�z?����M3��h�p�a�H~�#�`F���*;�%��ѡi�)p懆�]�V�&�i>�'�O���ie	24R�q�� �<��O��n��rb�L�SG��/^��Sn��
"}�̓10U���<���M��'߉O}���'�4y0�� %:;���c��G�8�p�Ow
�
�O�=����i�,��R�hO�����$r��*��؈@Vyb�A�O����d!�$٦m�DOc�h���
�����"�ę��G���4�?IL>�g?���M{��#E\|C�f~�p1�� 1#ڑ;�K�=�<d̓� ���8	AP(2��?���ں+w�h�e��i�U����'��AD���c{�4��HyrS�"~2�#΢d�<��F��J���ŭ�|̓ �ƈ[��D��$�w/�1 Ϩ�˷�F;~�(�'�Q�<(O�7m��������H��l�胧��7q'��ԥOcn(pǣz����\��#amޤMPn,$�����U�����G�����
����C��&���	M�ɂ�M��(�]̓��	\|?��8�i�-nOj���J A��	���O6�x��$>�� �1�*�0�u��]�
�d	�ۭ7� #B2?�'qi$t�A&�$��x	�y��)6�A�����_�2(�/O���<�|�'Ĝ6��,��2�'�LzIr�&2�X�����;޴�����'1�v�e�&a4�I��}zJ��q�.6��O���׿O����O�M��� ��c��� #5H�xT���b�%\b�0V�|�(�'ZR�'���'��Q��S;�����
��,�+����-~��ٴ>�H͓�?������<I���yǆۖZ�x����8����4@æ��7���!����4����������MJ��YV~�&��L�.UXUi](eh�DҀ9���qElR�L� �=	���?��Ο/lE�)��@�
P�Qf���<�.O*�O�	l��<b�<�fF�,!S< �`eB�J��`s��ß�&��j,O���b���c}Ri�cǔI���P����S*���y��'���:%�K�p��O|���_�x��O��*�mW-�6��"ج}X��R��<�,O���s�tԮ�
x���dOB�b�+@�VI����1���"?�iҘ|��m��EJ.l�6`�רՔ}�����'Q��Jcӆ���?dz�>O��dP�A��!Y��I&�~i���%�:���n�@�H��7�D�<�'�?���?����?���TQ`t�]3�xs���7|˓G�v>u�7��OJ�$�����G2Ob���41� ���J�*0�v]�ƠŰl�D�'":7mCȦ� �S�S�?����#��5�C���$Od)CC,؅����s�%>�b��':�؇JJ�t��P�1�|�Z�<#Vo�"W�h�FCռ+�`�ʍ��<��ԟ���۟��qy�bӾ��6O يa��W#1㍷�PP�U��O�ylZc�i>I�O��o"�M�T�i�D��̈́�u>���7�EE-���w%�#,D��'��dK#naH�;�M�uT�I�?�2X� �]y@"� B6��!��^��:B;O*�$�O����Oh���O�c>������
�v�B�?��8���,y�^Y�'",m�z��w:O�d�ͦ'����m�:$p�Gɯ
m�*�7�M[�]�|�4;��OUN��E՟�yB�'�:���W#7�|Y���/e�m��ԛC"8�ڱnI�U2ў��	Yy2�'�A.�;�*X-�Xr���y2�|"Nx�||Cg�����I
�M<�B��-S���cF�2.o�	��D�Oj7s��&>9���W��!Z(H�f=�T�V5�\z%�A�����<?a�'#:�D)�9��X�5�ߓ<j��8��ɫ^65�(O��Ĵ<�|�',p6�շ7�^-��@Y�-����霑1�8}����4�?�L>�g?�޴5� �eJ��zD�[������A�i��A�x/>q�'�˔�$N������;��$GjjR���:��I
Ԁ�	1O����<A����%i�Tp+0��G�jC�%P0Do�n}�c����J�S��M�;<�R)�fgT3sU��  �GQ (���'w�6?O���?��S�
���!���,d���9$(37H�$�؋"o�牙CR|eB�D�0Bь�D{�O����S��񐥈��8��vc�)�y�]��'���4]t� �<�@J\5 �� �G��4�m���?	J>��U�@�Iئm�����'"ءD	Xh�Y��֤3?��O�� ��	K�(M�������jA�tFMߟ�g�[K��B�� wv�h��͟|�Iݟ��؟��|��h>��?����N����"��:/P<���/䛆kI�y��'s�6m+�4��Ή�!e09z"��<L�Tvj/������4
֛��];p����'-R��DN�I��_�2�\�(e�\ 
{,ͪD V�>r�񡖝|RP�`�	۟���ӟ����pd�9/�Xd!�K���8� �XQy�fhӒ9�7O���O�����d��'�h)S��:^���r�߻Y����'�7�_Ӧ�c����'���'S���W��!:M�|�UE7^�><�� Y��I�(O"m�&F��l�+&�.�'� �0gA�q�v���퍓\*�x����ħ<qJ>Y��i=��[�'e�0�5��ΆM�� yb�U�3O�m���$�泟D�	�����_{l����t!�ˋ?'����½ J���~�����1",��g�OJ���л�0y)���
��C%Z�B���:O����O.���O��$�O��?�A�ݤG��˄m<��ۅ%q�\�Iݟ���4T�V�'�6�$��Ơ���6O�JA���tn�)�Z nZ���ӧsY�� d�OqZ- &�[%�y2�'�(K��%�r�A���J����a@��?���� dVў\��gy�'���I�Q�Z҈4�H��Z(ɚ'��'#�6-���1O.�'u�l��s�ѵ7����MF�.�'�ʓ�?�4�y��d�OP�u0�˨j����`y=I�WDF|�
�q��:>Ĕ��r��8vx�)H>��� 4�B��媅�i� �����?�?���?����?�|�,Oڸn�:e���	�X�<�c��{������<?���i��O�1�'�\6��<X��6�?v��E��12ք�l���M�&gܐdF���?�w N�.x���B&���fi�Ѣ\	r:���˅3��D�<����?���?	��?�(����ņ��D@���֐1�8�ڦ9z�`u����ß(&?��I��Mϻ)ʹA�P4g�b�k��X�=�<�7�i��6��,ק�t�O��t4<(�y��'��LWi��jLfxH������a�'���(
nv�k�|X���	����dhF��e��(G�#�3k����I�t��ryBOퟰ��'�r�'(F��$nn�|;Q`�r������c}�`Ӝm�?a�Oĩ
WK��T)p�b�Ҫz��&<O��D?q��ڷ�K�w�˓��4���-��]2���Đ�� n����҇.�X9���?���?����h�d���B��(��I�j���WO�Qnd��MӦ�k��b���ɂ�MKK>�缫�@[z����bN��l���#��<���i��7���ICeJ��H�	��$�ei���~Dz�.2.a�p��Ɋ/s*P�&g�npƌ&�T�'�r�'`��'t��'; Y*�ț(*�|���oN�+"W��X�458�pR�ip2�'���#�y��'flȺ���^��v�<v��⃦>�U�i�07����$>����?��کH~�I�E�S�z��oU{\x��G�FyR���5٣aupўĉ��0jڊ��q�.hGB@�s�ܟ�'��I\�	��M!��<�IƁd��� wᄨky`X��	�<���i�b�|��~��'���'�	Q�J���b؈'��wk0-yG)�-^�	�'���&tA����P���d�(p��Z>�P˦C�
n�24�%�t|���?�.O��S�O6�y3DS�k��`��,*~�y"or�6��Ɠ��
ܴ�?�(O:��4�S�E����p'\\��a�̖'^���z�R���x��3O\�� '�n���;�*���H]�E�u�1A9M�FY(R�"��|Z/O��	�cK�X+CŊVo���� Dk���(���ǦM"��)�	H����2�Py�f/;Rhщ@�����Dy��'���=O$�`��AO�Q�0���`54�G`��!���Ͷ+ �ّ��d���Q,R���$�Z�����R�hB�D��L�!�ϥ���J�i� u#���%�&\�џ\�"K&ڭ�6�]�nqjS�Kxz����R-{�B��僇L�>[E$��"�De��;J(�l��_P*�Ia�Y;W��qQ`㎝x����#�Y�? 
U���q�=�b�_lC�Dڱ*W?)H��vո8�`��L��Z�IP$�N��E*a��]':��2ڀL�ͪו>�����j��&��3,T�&��'4��']�'5��'m�D����88��1��R=08�Rm����'\2�'���'?��'�����{Ӷq�'�>h�D�u�(aŲ�����t}�'>��|�'?B!Ι}q2 ~H���E�`����7,PY��7M�O��d�O��d�O���_�|���|z���'6!k%j�69�nQ3�Z���Ig������I&=,m�	���	�O�l�y��V�YX�,�VV(h�޴�?y��?�j�@�Ĕ��'8���I�U���"�</�dt�B�W�/$RO����O:0�j�O~���O��O�����)HGǐ��b��h~(W0f�s�	8U�>��qDP81�:�v@�0a�P��{l��k�;z+lPC���R0f�H��Ѿ/�y�i�'w�C�	 !���5#GH݂�yQ�^&;J,r"K	�T"V��������"�'1�̐�d���9Т[,:̲�H�-d��z�ȅ�R���u�H�:c�za��a�H�U�H�S˶x���>��'͎�F��h��&t�P��bq�����2?P�1� -�j8ДhE�?���j���3����˟����H�_w-2�'&H����ͲW�`��(�|��4�g��2c���ꖉ�p��S��Ƙ����I�d�P8��m��9T����E�qX�R�IK?s��%�s%�6j.�g�?�������'c}2���,��O�/���҃�~I.�?)%�iN6m7�I���	XG$�Pq��a
�!�.T�G�!��Ob-b�KX&F^	���=+��)y��	]�'�T7m�O�˓c6��{��i˸��K�Abz@c\K�<t��'���' ��8�2�'�}�1��JW�u���gB]��h�Q=d��;H� �@���ci�"?Y�� =!���C}}^5��L�*���rV��b�F����(J���,W�S��%LY���P���럨�A�֐wR�QoU�d��X��*D������#�H#S����I��)Ọ=��̍�g��L	D-�,Tܩ�׫��<�!�i��'����bj��d�O��'�։++V�Y�b�,��j6\��a��?���?)&��8p�;t-�*7��S�T�³AO��^$ V��� P4�(O��B�ϳQ �u���|�'v���&�Yw@�3D��M/UDy�bQ��?����'�?)��H"�D��U�'��(pI�>�?����9O^-	+��-�
�8��E�rv�)0�'ҤO4k�ʙw���7k�9XkZ��=O"	�G����E����̔O��1��'�b�'r���B�4%�r�i��0t���2bA���/5�m�G�t�v�T>��|�	�*�L��л��6��~�쐐�H�-�H���N
Q>t٤H Ɯl١.\ '����Ͽk��]@"��oQh� �-��&������ɧ��r&�-j�ޝ8�IF�}��1
A)�y��]<?td(_I�
|�Dķ\"<a�)�Q�X!x�E���D�`�lu�ի�?�?����L�&	�?���?)��o��n�O��+6&�0ud�:��5��Շi�
��44�V�҃Cҡ<)8p�!ɼ?�=&�-TV����3"z"Ѓ/W�d6m�f�PIU�A>2p�s��hO��b�ЂyÀ���]� TY�O�F�'iX���͒���(�aV)E�$ہ��)�!�84I�E�k�,�Ly�M��:C�|Dz��� XGL�oZ=��<isԞW�T₦=>p���۟��I� h��������|�p  ۟��ɺn�n�Ӡ(�(Pi��xrd�;�.���O��I=8;�%
Ù�Z��]KSH޲*����M y��Nn�N�� "
8Z�Jp)�/��/�y� "O���%�\T�x�Pd�ņ[ϼ\CT"OlmpJ�w�`E2�O27&l��b1Oz��>I�hϢQv���'e�Y>�P&��5Th���� �*`qG@�͂U�	����	�ܴ�.Q9h$q�J��?�O����^���B0�Ȼ1d\tY��$��3�A���*��s3A�!D��P�/Uv�T���@�Q
 �Q �#����'����G�td�:n��Xs�1t�L�鰦F9�y"��;�����hL&q�h����0>r�x���$0���m����V�y" �?E�.6�OP���|�����?����?I��S�fж ��	9l�i:t%��\�eI��8� i9 ��.e6~=�b�?y�|�݋' $�{2"�`��22+�<b$�@�<ar��jF��V�B��MqDҢ'K�����B����w:�=��E�q7$}�W�o��0�CۂLY�d2���O\�S���;V ����H3D+��D"O�S��ϥB�dP����y�&��	��HO��O����1�6�B���u��0)S��OL�n^٠�N�O��O�d����Ӽ��A<CL8x�����;�0pN���`�<j�PH����%����g�'���#m�CR���ޗ0 �q�ׂ�TPG��h��50����D�i6eҟ���Ϛ3$*����۴�|���:-���M�>���'戁ȥ�@�){q�sJ> Sف�'�X��5� Z@��Qā�#b�jE�f`*��|J>iĪֳs��� ֥�©J�8��I�b��p�J�O~�D�O���R�?�����OD�1U��U���i�<QP�	+Q,\�c�]1_�k�h�F�P$䈂��OE�4��p����6�OK
,!��#�h����Ř�.0ط$�
H�\\0�F =�\�b�,�dF!=�lӰ������< X`�S�Z��D0�"O�E��͔������J2Hڈ����'�ў��Lۻ6���'��~ݎy�� a�@��4��"Z�s0�i|�'�哛FT�ɲ�ı:�p���;GW�I"�
^�4�	��K������<�O� Ȉe�V+0���g A�~�hLÎ�d/Z��?�"��
�f�0�ƐN&�@c?ʓ7������H���
�D�%sh��e�+!���"O؜2��=ظ$�`n�����'�XOx�k#X������:"�����=O� ��	R����͟ �Orz��V�'z��'TV���	�u�6�� N�Q�[A��}���E�^o"�QV��O�Sl�矀��ß0�\��t���b-|T$�b��0mB�d0`Jݨ�8a���?��X�W�/��;wM��hf/K>es��LQ0ls��ʌ�?Y��|���'{�E�(�0l�rt{�D�rZ����'GҤ�R���2�"�s�>��� X���d�'غH�Ę%o�x��m�gI��v�'x���e?�PZ��'���'J2Lt��iޝ#%ǳU`��jT,.<�11R�������/�O�|��O$T��E ֊K�X0���O�C��'#Z" �]��E�aD�=41���'�P��1�a{rJ�  ��Րs��Pʩ�@���y�NW:�j�!��]�<)��0���m�"=ͧ��Tr����i�&��呠8 �
ӡ�-hJ���F�'r�'b5l���''�I6^���'\9�f�Q 
<t�j��T*O�U��p��M�'�j�;צR=5f9rBԐC�T9�RG}�	��M��ʏ�0��F�	��4[u*W�<#���VX���Y�&h]�B��Q�<� ��b�ҴKp ˈHl~��!��<�A�i�'T&!)P�b����O4�'
�0@�l�SΌ�P���hFi0�T��?i��?Ƅ��?�y*�PW�$Hw^�q�P�� �Z�'J|`��)���a#G�;͠L�F[.dQ���@��O�eE��T����T�ҏ2�6�Cb�[��y��h?dT+p�B#�}�H��0>�g�x2�3�P�9�@B�u@��2 ��y2���&6��O@�d�|2vD��?a���?u�{�K����|��@X����G��tFO�b��8�h�/O�(����4� �1��
����&ĊZ����R�GO:"Y�@�H�sD(Fq�x���'� 7�
ky����Ү�Vh��i	��3	nJ����y2�'��}��xX4�qBOG-��-����O@�Dz��O�L� )ZI�ۮmZJ��̛�/���'�´����Y�"�'b�'DH��<�ɶ"��	�뒰u,�=��O5y�p��x��j��R�z�d�
$��v�'7h��b\Yh��� J9�A�5O`���C�9w0L��U-7џqK��0o����Q�Q%2���џ��f����ش�?I��?q���?)�Ӽ{�C?U����I�|�$��
U�<qa��nt�p7�ϴT h̐v'��8��4�?�+O���EZĦA�)���:�:�)X4�
p�f�@ԟ��	����	9h��͟ Χ����֟�3��;8d��3��}В Q��1�Ox�*�R�LK��ip��B /7��Hء�0�OJ�b�'?2 [���������R.��{����ya��.T��25�x�R�-���yr����j���#y�q��+#�y��n���OxP�Ċݦ����T�Oؠxa#�����E,ʕ0��5=��'8�A�u�J�R0��Xt�e�,6v-1T�."$��paB��K�as�����@�Hq��!�L��Iu^<��-x����P���
G`�9B�R�q����'|B�0ҧ@H��#peG�rᐔ��/�Q�̄�$K,-�U�_�kN��b����,d��ɪ��}9���g&�1:48@1-�� ֞����SS�i,��'���~㪴��ҟh�	�.�h,��D�#P,,m��.kI��`�+'ą3� �����5�Ǫ��a��c���h�A�c��rt�ēm?fi;gO�Uv�:ƨM7tW��5e"A�.�Atg )W�F�zW�*��;���"�C�!BN���mV?w��q�h�/�?�6�|���'���oӐG�!�N{���'m�HrDm�rЁQ��qQ:���ĕX�����'>(�3V�r�u��IT�\���'&���%� �k��'4R�'*"i��i�� �HƯ����tpc̙���q4�O�!g�'� ��Ȋ�.���i��^�S��]�%,�ܦE�X!
��\����9�r���a�N�,�A&�)�	���N؞x�*ۖ@�0��2�$_X�b��-���I]�4-[6Ȁ�p�ȉ���3
+��4���O4t����a[W�h���p�왼g�i#k�����	ܟ����kM�i��ڟ@�';VI����+G�y�"��'�F4�"3&=��
^,b0�p1LH���OJ����LŒ� �g�P2�"W:P��h���ΡVo�lqW%��C)�7��Q���$ÆU	r�m�$!���.\\���ꚵ��}c���Ҧ1�ITy��'q�O��L�v�k�'�/v�"���S5-�LC�I�T_�P`G�CiR� 3#C�p�扼	>p�IQyR�_
�$֝ş���Z�T�A�y����v,�=b�X8�O�i�9���'���'���
Ӏ(k�R]B�j� Y����v���Z���h_&}�8��4���%��� ��(O~��n�=m�� f�б6@z�zr�R�$٣$
�z�p�(���W֐�`aaUx� ��*��Ux���*�'1U0pR� ��)�h�� L��-�ȓ���A�"[I�`�ѠA;l{\p�'�ў�0�ē��xcT.��T�V�Q�Ȑ���Yϓ(_�����i��'�S�#����Ο��4��)b%[�d����N"cܹy�M�;V>�-{bI�K������4���^qp���/\,���m�.yT��'�ՖpǢ���'O�O�����L0K�^���#��#�Yk��w�&��e��z\F�v�Y�9z��P�R\�B4���O���C��4s�P�����6"Od01���*�yzI�&�2�	;�HO�i�OB���&E�Xѷh�!� ���OZ����	�"@��/�OV���O���]���Ӽ3e�!F.b����	6� �Eǖ{�t�kW�� -oF��G�n�	���HO4
��K�Nd&�ȠlY�s�a@Ю��	x���@���!9c3���a��訣�Ԏ	'4��'r�ȧ�"CGlH�F�"�����cdh�O���I!k���'mG��M{���3BC��PłQ����!�`)��`Ǽjdq���4�*�O,$3f�O�ш�C!,2H�*D"�-��b��N͟4��������B������xΧ.���(�M
�k�$(�(�d��Ga
	��!�%�Gn�d��ʈLzfp��(3��� 2#܀tNx��R��;30 �2�Ň "�F�Ԍ/@r(B���D�X�AӄX��q�I>y��џ$��4G� 9 ���`�K�{z�U�ȓM�yw%�2�P�eoÐC~�����y�'�6�B�ٯ@8�<XpK�4m�*ܘ�'[`6-'����WK��l�̟��	t��� �2%[���8|4m#vD�)} 6�#�'�B�'Wj%�D�'�1O��1�� s�A�6+�YӤ�Ժ�~�<�j�h�O��`KA�c��bA.�:����D
���S�^��9���1@�8�W@ĔS�:B�I�eMX��AC�S6b��!�C:0Tt��$�q�ɯ4���y%3-/0��遈do~�	�;�I�ڴ�?�����	�$hl��O���gp|�R'��Y���j�
��A�,C����Te��9�����S�d��w��1a.m����v��-�:���gD%��q�'M2G�e�J��f�}�]�c����b�Ŧ@�Q����8�pU��ߟ�RH>E��k຤�c�b��JI�&%��2��L��oo�}�Q.�bhT8Fx��2��|*�~�,-�҆�"{� f�@-K�&�x��?9�g������?����?�v��8�4���3�T8>8x�yQ���?��4����NQ�@K� %d �R�!v��4ғU�|�x'��*b|��p`ۘkΖ3g	
�wwV��@��
�Y%�y*�4P|Tu	_I~bk��2�[�J��l(8���%�~R�ݒ�?yG�'�\��U��`	���fSo����'�j��A��Nޜٗ�ȩ%�	2�E)��|�K>� !��]���ǜ�tx��J�{v.(��QMzb�'�b�'�x��'��?�������_�L�.�x��p�m$Ob����6�
�FlP�'�¢?�7�S
P���Œ&�ֽ��	���
d �+�).kf�3�k�Z�X�۴5�pI��#P�h��]����M{�hٶl"=sqdD=_��ex@b]K�<�Bo�����;�6-��M�&-D�<	���$��#�C5gd�����<�F�i}�'-v�x��l�����O��'7=�7�U�^�"a����DFH�D�?���?�`	{�`����C�T>9V
KZ]��/^�]��[b�"����	�L^[S����/w	P�T����i�V�v���(�;�*�3���(O�Qy��'t#}�f(]�@u;���2���Ѡ	S@�<1�&�%_�<D�	�C����'V��I<As�ԸT��u�5�D�iU"��<)El�Q2�6�'�RR>����̟��	���S�3�����h��M���a��)F�9��ʶ����g͉v�Q9��hc>�� �)��"U�Dv�� +AJ�j5�\�KC�U:g�ڤ<G:��]�a�᭻m��yFi�\��w�l�* !ǚB���0-�8%�/��"':���O� i��:{.����q� �*�"O�	xG�M��"4I�� ,Aa��;�HO��OX����JU���� ��<>���T��O2�D��as��1���OL���O�������Ӽ�%D;S��u;��]�D�g�y#52��T�����H@�{���'�HO���%�+����/-4j�BBI�0z<�h*�g�&.LV�B X2��	}�R����6=r�I<h��E��]+82�
"�
�e��I.
�R�P؞\�e(\�,�����ɊBh��y��Q�,���S3��	<�F�V�ʏtV�"=�'��:~���i�^x��ɑ�m��1
f�<cIT���'�b�'FRK�*}���'��	M'Uфӆ/��I�ԉ��}�\q���Z��Ȑ#>\P�t�;��=h�����;p�t�[!��:��D��:Ix��Ґ��#^z�҆��M�ϩo{�=1�����p1ڴQtx�ஔ/�\��s͓�C��=�ȓ�5�`/�4����FAX�&��ȓm�<����'P��i��Q;I�(�͓g���|Rf�&�~7m�O����|:7o�)Y��u��?d�fo�:�����?i�b����CU%?��^u�@x�F�a���:�r@���5@yt�Gc��(O�dq�P*���p�i�.P4�̃D#l����� �sf�E��/�� %̄"g�G�&1D�6�����m�O�T,����Z��J��L!.�mQ�'t� G��*=���C�A�0Ů}���'LP0���L�L:�e	wӀ�P�'�摃��tӢ�$�O�'o�����?a�2���{7"��&ָ�����j�.Fq�%��[�#7:���}����åJ6M�I�֣�	��مǕ3r��TG[/Y��m�ɈXw��mHd������i����sr�җ�^=�L�iZ'I8T���h�)�� ;�.Z�� v��&�Dc��3D�|����$Z�4m��F��G#<qV�i>y�����u1s&��w�V�:%�
�f�����ğ8�V �7��4�	ݟ���ן�2]w�w_1SBڠmI�'���U9���$����ʱK���o�Ij��Ҕ��t�	��ty��Qf�CRM�p�ne�j{)�nKR�=9t'\#s���s�R�@b��z��6pa�c��A[2�0�@�M}��ɂ�����Y؞d��Q�	�4U�a� (�D+D�����[<j5 pG!x-������HO�),���z;��nZ"0���F�Ē�p����(K�!�	ҟ�����|��.����I�|��c��/�ҵsaB2��P`f��C��x��+p��bb,H�fTX����	�86�T�;�JϨX#ReB���f��Ϛ��ۮHn��K��p�(����-h8qO�܁��'�(6���"�*��g�o(����oϟ%!��H�1���gF�w6n��1�!!�Ud��  �k&{E�T�l�Y��$� @���4�M[���?�/����F�8ifHaBJ�rk�I� ��*!��$�OT��[�9�ШB�S!/�� A�E
���O�`���"B�;�2��O��DԸ�򤌖M�`m��N�����k�(����au�D����&5��|�a�J�2�{ѭ\�
�z㞠�V.�OL�E��*�cc��C�Ն8�V�j�Ú�y�&��[�����"Ե-ܩK��S��0>��x"D�S/6C���<|�;3١�y�f��\�7��O0�į|
p�A��?I��?)G��:���0H�L �	��!��z�� �:<�"��F�֙{x ��c�?q�|���"l^�Q��"G5�-�㝸���0`e�İKe��#	V����"^$Pm�~A:�*(��MϮ��I���Q�?�8�@�������'��O?�����lx�A�9\6u"���2!��)1�`��4�Cx�I�Dǭ�1Oh��R�����'ު�'����}��(S�-Ą g�'lrO_��d5��'�"�'�	�~�;pY��`�/�@�AQ+��=Bt�*t㐳5��<3�G�uH`B�w"��lR.b��w��IK�E{���S��4ȗK�FF���E�Q�S�.9��J��N�x�4�J9�����9��փ�:����.�$BT���ڼ`=:��ݦe��t�'�R^��j@��$�5D��n8	@+(D������u���R�j*@�B���$�HO��)�O��q<�=�c�i[:��gm����A��*0�����'���'.�KQ��'���H1+����c�W��A����N�T��aN���>����S�H����ڊ򄘵�>�7/_+`�I ��H���� 
�0"���V��Iմ� �n�4Բ�R���*���p��A�G�<.Z�qy� ��&���:�"O�hc `ٟ"�e����j7a�&"O�� ��@�
q
�@�K�!�d3O�	ma�	`��4�?����)�Z��+��84F����bQ���O��d�O|S�&]��4*���&=QbX��@�Uf�(q�V��-��9}��1v&�4<�Q�T��LZ�;�ڵ�B'8\��!�-ÄASc� "��@�F!�4(��+@`�i�P�I��*��@K�O��qqVjG~����l�8-�}��'�[���%�ha��)�Y�伹	�3.�'��ء�H$JG
�*��JM�%��'/v�0��`����O*˧]̤ Y���?�� ���(4e�0� £>�j�p��� 20���$|��jA�س:l�SZ����B���-�N�d��Y�с���G�f@�2�o`^%"��o��E#���w����	L�@뷤c�B��w�N�L�B�*���O�Ӧ�/1�Z� �o_+C^�/�y�G\0������)E��7���O��Gz�Oz���=C��B%."?�tͲ����e�2�'M�D��C�y�"�'���'�vם���	���qc��4TB���(J.D=R51�i)r����D�E��XƮ�qF{��R!�2�򂮉�dP�ʂ�ؤ9��P1�_�.�FH# ������Oސ�`���R���} �F�2oе($�,4�04��'��}��O�r�l��JW�5s�g�~�<�Wh�A=�l��b8�D1�똷z���`�I�O|l�#ܴ,,`��'H�C���H�)�g������?���?K�?���?A��@�b�D]���ΚaB�u�1d_�_�<���''�V��w�X$���?��#ҹ9���5(�v��F�!�$(��
�2ݢ�"��Ϫ`b�	s�,�覭Qf��F�zx�&�|B���?�&�i��	� OoNE(��M�
bp(�"��O��d�Oz���O��� �D�=y��Mp��8u[vx�o�3�1OB��$R�^��`i3�IdVB �r�?dC�čᦵ�ٴ����4y���n�ٟ4�IG�DB�����P-�:ym*I�ׁ� �6c��'���'&�k�kC+�����Mc�Ir�'�=���ƒ|�^�{��J���EX�U%�(O��C��Ɖl��h;��F	<�E�ԣپ"+����M�ҜA��ӹ ���
�&�ؒu�>��n��E�4A�"b�Y ��:zQV�8���'�rmCW.WD�<j���P��P�
�z��'������)И���H4Oè�{�'�:��y��D�O��'�A���?���\h~{S͊�p	tK�ES��EK�ګ����Ķi,r�#�&�O�x���y6	��hsDmA�!�E���F�D�؊ `v�p���8yvP(Qs��H�F/���]["أd`�)'\Z`�5ʂr��ť�=�?qו|���'�D�;�F�5�T�K�
����'X� ���-2���U��;O2E��y��'��"=�'�?�D��=lX��f-�6l�<����?��?P�Y��!���?���?q�c���O��(~�����(�LP�t ��5
�D�/p��}�S��N(�dL�P���y�!��~��<��>��	".�j% [�Z`I��	�����X	���4|O���$��B�(�!#�^�~m�"O:��S��k��!34�>�AqA�d�����|��2�6��� ���([ ��Drd�D
Q�D�O����O t�2@�O~��r>]ۧ�M�
f�h�F��2{B��O�4Ѷ!2a�(��$`�!�t�*�:�U�$�Q���AK�^�aP��N�����/��)2ՊD�U��-�W-�=}Pn���+׸d�Q��[6��O\��E��ZYE��X�X��P.	��OT�d�O���0� �GmA'
�� Y�M�=46���Bz��Q �1�|���U`+��Γs��&�'��I�\�Hi��4�?�����)W�3��*S G�I�ZPl�d����D�Of��Ov�0�,�e� 9KfF�Ih����|R5�E/�D��&D:6) ̺�$l�'�qs6�K
rF䃵�I#6@�|�ä,l�l����>#^�C� � 
�@��#!�)d��-�=�����	��	�k2<�����?�(�c`�z�!�$��Uu6\	D�<���B��{@a|�@"�L�x���J��)0� @�E	3��	,
R���4�?a���iT�gq�D�O
�$��;rT)�� +} 1R�B��oJ�� �K�$򐱓��>BDeh��b�d��w�,���>p|I 
��@�lP%*�F
*���˟.ͮ��)�	k���3���B/��;@��A{c�<K�,��7�N#8(d��?�d�|���'����썪�F����*na���'�����BE>e��Rp �h�������l���4�'���c�NR9y��\�tc��^n�y��'��S�I�u�'���'��B}ݭ�i�Q	!�8w���(�	\"
��ãf
dЉ��ʕ�d�\IA�G�`�S/`�����$Cf$�ᧀ�`�`�vA�-h)8�7��Fc�P6	=kz��ԟh6�P�Rݛ&�������i6�6��5';��T��Q%���Ca�`�D�O>�ԟ��ǟ,�'�Z��)�4C�8���O +��
�'�R*E+\��k�?J�8�֨+Z�#=����?�)O�Dcʦ� ��E�X<���Pf#RtsE�I럸����$�I�3���	��ΧEL����h�"�F�T���FT U2F�3R�;�O�uyX�8sD�X,�x)f�ЁU�L���-�OXY2A�'W7� ��R@矔1�"�y��N�=����"Op�����<;�m�1�ؒ�"Ofe��F�$D�����s���g2OJ��>`��]m��'��V>�`�@�3X����F�< �X�öR���	㟼�����*��*k�|�p@��n���~<Ҕ�_�A��A���Q3��r�	�@}�<��K҃Q�t�� QfR�U��&�4�2e�,�nIY��:Ke�F��22E�=�#�̟�i���~���s'0*�bp�.؅�PyB�46>b<a��/v�"�"�E\.�0>���x"��R��8*�˗fl�P��L�y��ݦi0���?�,�d����O��D�O�A���\C�X�)�"���y`�ۀ��7���A�ȝ@A���1��'���<	b�LS �rR���b��W� ��GgΥRP��9V뤭1�HL!���A�@��w?V���8+�~)��$1d����C�L&��'��6-�Op"~�I�vX�q�d��+@��뷣�$nv�Iԟ���ߟ|'���?�lK�|,�����rP�lI�\�'�6M[�U���M�a6���'$���fC'}���`g"P+!��?ig"���	��?���?�w��T���O�(�f'5�Tp�b�6ng���CC��l+@ϙ�.Y���uF((W��	�3�&�mK�#���P��Þ�@�Nʬ<�A���.��s�?M�u��zVl�0�����gn��.1얁/FJ<�%/<DK�DK;*��)lOF}rwIӅ~t���i��A��"O�!%��0?y�<��B
�!�b��1��a���d퉨+�����lX�R�"�@��Z�[LC�I2>��I��9�0H�5oT��@C�Ip��"��k0h1�c^��"C�I>w8�逄/[/A�\���	���C�
{�uC�-[%��ǅ\-�C�5"�xAH7�-�����5d~C�+%�z!���1Q�XZ��  �B�ɲ���B�b⺈YU�K.t�FB�I�%^��pq��/c���� E!(B�ɠ5��!�f/�O�l�	#�Z�n��C�� Br��4�X�7T5	RBӫ-5�B䉾u��	9��
^_���p�.��B�	���0S�#몡�VĕC(�B�	�!��0�	�iA��̔�DO�B�I�R���6�Q	 �1
v���R�0C�I�u��Q�	�r��HA�#̔j��B�I���@�8@g�,� �	 ib�B�I���K5��C�`��v���~B�I�j�:㋞�&.|	 �.I�nB�IO�l��,�l8ԵQb�A�{�B�Ie.���!R^��p�wb@8�bB�	8oD
A[�͘�i��p㇃�RB䉓F��`�u���Di��� /��sxxC�Id���:Q*ܝhC�D��$Z�C�I�\8�BߚC���#Ő�S4�C��2Q&���IuJҤ�#'�2V�pC�	0�,=�3���k8�$%P+3C�I�,�qҲfV:=o�����n�C䉛FI��ڠ_�O|�;RK>U��B��&H~\��7��(�ӆm�k^�C��)q�����1,�S���!�8C䉕L��@��!�?;��%ۀA�X�C�ɠ�lɋ`mOg�(�i ͅ
J�B�	�A�8�N�;,�:p �N� =��B�I�-ۨ� %�mY�z� E�g�C䉍K
�[�.![�,K#oA�!`����Ei����ْtr�S�Ol]`T�Q�|5�� P��}!�D�R��1;oD�S[-@Ua~Ҩ�:7���!@�w>��R�FL.o���O���%凲t�rx�;V�n$?�i�59Rg�V�3$��jK�� ��=�O���f�J� �u,�Y�#V�I�>�ZaGH�`�X���x�`D�p�C�U�Ա��H�|ɸ���f�(RD�������>d]q��/s�
+�����%Xw(���DКS��|@�!
���Y�q�O֝A��O���&>c�8�ǫЫci�p1B AA�̱C�H��9<
�8�N7c��@�'��(��Wu݄���.��Z��R��B*x�R�E�9hm�9���� ¥ju$܏K���'��3�t"OPzuI.~J�4b�	�T�"�3B�1O�(K׀EdLR ����^\��ףy�b���"�#訝�DȞf���J�@*�0��A�����W#����X%`�Ś�{`�x�BШE��4����Q{j:��L ��'iNʄi�+x���`
�/"��%Ќ{��TiHw�@#\�yB�%��!�2�k�lP53�	��B�j�6�%ÜO�R7���i�a{B�ݐ �j,@�� �tn��y�G��&��"��K�.��7��xZciX�s�QcG�Yx�m�n�J���E�}��3r���W_68��~�	�f��E��.!M��jfL��p<�m�x8�5����Q��E ��ќmњ}�%��
\/.�� ğ�����N����
ǫK�2	��$���D��`��:�� X'��rNY�-XE�	Gd<���GK�J��SU�<@kDc���!`,d��Z��MZ�h8��>}��'4&�r K5����k��N>��ϸWI�İ�kк@y���g���{��y�L_,;�	���E}R"	"`�0Hs��V	���B���#"��!  �7	j���$TJ�xZc���1�A4�����b� 8M����@�O^������;�f�ا�L�:�L���'��U��j��s��6���=�b��0��l#&q�g)��#��q���`�O�P�9�d�BE�,���Iu�&y�%@�$`:�0��oH�H�����&Yx�ɰ6�����]�04� D8F>��h85�ƪF��Dx�	ǿ�|�I� ��kx�h��'��'�D^�g�p��M>I�g[(�3��^��ң�
Q�s��#0h<�1��<���N?C`ߍW��]S��F�P������Ҙ&��z���M��ô2s����~)�T�\�m��)�1�r�z�s��|��v��D��䥟�8��w�F�k@/վPT~�[���:�>�zǓ{BP��g�R����0�]�c,-��a�?H�̄�U�GA��u�!�O��I���:V��K��S��|���H�Z�,,��	ڲ8�d��k�-�� ��� r�'����ɓv��AY/�uv�9�}2��=*5<D��&R!*l^Pk�@�'�~��'�J�GB<0C��Z���C� 5��QZ�@�/�{�R؊@��/
�Ѩ)d{���#��Hdџ��v�=�ƨޘXWa�@�F}�d�3(ꌋqmQ0V~����5��@"���1��/����#B���O%̓��X����b�{�m/u��:��Z
�x2��=���{��6|�h(j��H0,�i�T���	�]20�NQg���F?�r��`�O�7�� {�D�+ۿ:�5�T;2,h�*�ΣE6*�L<�Q��lU2���7��hC�m��$t١	�r#P�:�S�q.8���?�@�DT	I�v)@F��8ΓO���֍�<�B�1�D�Ƭ`�ꏪ*]8�ɗ!�8C�<�D�Z�@JqeA�D���{�X�N| @��T��H�A�W{�Ĺ��g8��ئM�6uyU'!���p5-@|�ڢ>و�W?�!Ny �CC�=��0�D��}8�pr��-)L����`5.vF�сF>=�8�z0����,�����~���|:���d��h$�Xy�U�4�h�Z`k��HSĚ$�TO%�ӱj&�4K���*����F+,ͱOVHq���M��`A��իx��a(��O�ml����#D�*VIs��{�&`Â(�K�I�y�L�A�!�5R�HI����^ԚS��9�rX!AH����OP	��Z(���<EsEфg�<�ա��^pj�m��(.�!����5� ��
aT�$,Z�+�4����_���O�N��B���G
��'	�r���c�
8����|�\���Pf�d)���_��q�J$y0q�R�Z��ē�d (srl�[Q�'q�,<[nV����Z�E�����A�N�D�gJ�83d4%� �VǄ1�
�j�`4_:)�!*�I�z�A���5zk�E.�_�t㞌 �ڏ::���$&.��Y ����2� ���3AF*h����N��*%˞(۞<`��f؞2e�]�� �W)g���`�]V8A�aA(a~�p��@8��غjd}A桞�Lw��E�I_�B䉲���%ϒ�>�<#֭Ħf�)��;��4zB�K��̅Qvh6>��X�²$�,q��LY�0�؅�I2	8tr�$U"X���򵧖�_)0�Y�N\� �p�ݨEr���D?Ra�窜;FyVDK��޵r����h�88.ʸa��,^.���?�VU+�F�=]�����ºA����fE��T������@�i�ʌP'�%ч�*7(8xk%�VΨ�
qJM2=�ayZc�)cT7\�I�%��Dz3�'L�����ϟ���y��ϳ�.����'�"e��َ~O��0�o��@0��?F���IC��	Ag �ѥG \O�QruJ�9�t���?���RDn��S��I�g��~?�]�K>�c��>��\ѧ�d�	:��tܓY"�(D+	_���a%��*�~a�=��EH5?0���W�@�����h�ɼ ˀ he��K��P��.	�	���	���������=�F��QF�I������=�cOЦ	�}a��o�]�D��p<��>�d+�%@4^�x9�F!��)u�l�'��)����3� �U���L؆�kaC�%wf����-Oda2��-yܘ�Cߺw�v1�"�R�u�w�E3.x�EeDq��ԛ&�\�"��ĻH��]�Ҩ"�DYH��	�B�p0
��P'���i����;!N�#���%��=�R��0N@@��L](����"�:���p������ƭW�֐�iY�ncH�I-5�n�p��̰Kr�$K��@��&��	&T�RT�c 
�ܝ:P*+��a@$U5|�������I?��� �*�2	T��~����|"�@�Wg4}����=MY8�;���2�T�z���<�ѐ����p<�1��|ن��\;`���o��EoZ���r�oL2�"���O2��N?e�CV?��6� �#"�8�����F�I�.��㉨@cL��B;=�&���n��m,��B0d]� �%y�HD��Q`�&r��0Y�W��T0�����'H�p"���=��a�"sXv�8�ĚNѼ8 �BK8`/�y%�xs,��0@^a�fێ_�@�Z�!j�h
�O&0��'NY=���go�<y��rR�F�s�D`�קE\}B䅳���!
��~���3A���L���iE�_7JR�܋��� �T��0����t� �ڝX
�䘺PX���Ն֏T$]�O	m�	�m�8�,�2�࠻�a@�^0�Ң��YA�#��K����D�0�"�<[�{5�����3gF3n�ɲg��w�ȹJK(Sf��CN��Eʽ?�̓XAJ �S�X�N��ܘ1�Ahl��	Ǔ"�:ܩwk�F٠����R���OM�^[�����d�zrI�I�Td���!|�3sLN�����O批#��<�" ���<�"�]K伔�v�D�o�=�I<)��Z_%yԋ��?�e�������!X�g�H�zi@�T�@�r@�1Zma[�ʑ"T�tI'܁G�k���4�[!`}:&��v�'=\8`@Dx�,hу���|p�(�˕#&�DՂĒ6}h��j���"��9cL\=�i҅������Ƙ��V�"���#���LMR�ɼ.U|�"�![=qb�B�$Okɗf�~Y!�ǟ%jр-;�ǪVϛ֨�?x��F)�E���Y��1���)g"؁������>���3C~8���gBc���A��,mxʘ
�"z3H5����;Exθ���Cq�(�I�zNL�R��+Px�0:��bʅ\�\��W���X��YP��0A䀉(�'#�V�(��MF�I*���U
�L��" �<p� �I�r8Xe[V�܀�z���ϙ�l"Z��pcۏ>��9���7MT+8nm��o�~����kY��|R�*&�L p�`�29��Q���H�,��`�� G�v-�WCh���P�F9�s�l�Yu��X���4��39<�ҷ�8lvNqAvl,-C�8���'����b�7$G�xZc���L���Q"��K�U�@���4X��p�'�+j��yh�N؟��ӕ~��f�~��b޶�j��	w*��!Ȱ)�H*
Ǔan&ݫ KS�`C.�"&���m|��q���"�Vd��N6vy� �[��Z�%�&�X�ȵ���$[��2�ȕc�?��9��F)X��&�	WXP2%͖,��j����`B��Љ �j�9X�=�3���Jw�!�π�Kݔ�5.�
G���2��Ij��!#
$��rs���c2ƒO�;�*
'p�1�g��/?�ڭ U`N�,�s	<����'���D�,LɧjT�@�T�p0�;U�tR��ÜU�K� @���T�_�p<�1 �EJ7߫_|ĕ�ϒ�&����'���U��Q�\b���0����l_�(�"8��� �hS�=�]�1���>�ĥ��CW�	@��`:\O~��bR�D��(�b�[8Z��aH��F0*�l}�M�<tdQ�J<�@�B��ɠBM�Li�
B͂M�\D�,�.��V���/�sk\��=�F��u.�� �nA4�-��
Ev�}	,�CPKW?1�(�k��O�(ړ�RD5t����"߰=��J��t�F�a��3�
�m.��Hb�>[6��;'���p<��w��$��۩ �h4yV���f���ޜȀ��-[�DZ�+��["���6����GW7D#%�лS���"c������i� bzR  ӓ���ɰH}�����D|����}t���(�Gz"�L~sv�ħ~��c>���K=qΒD��ЅB�xY��M�[����' .���R�/��ϸ'	RU����	�� GO��Ybߴ
�4�3�N�Td(��g��"|��&Qʺ�f͉[�	[���=%��(�c3-�Н�aɎ���>�wjYA2(�7c��z�`ã�~BI �Yթt� {��ݒFd����:&�w� ɑF��?��xj��'8�yhՉȊ#r�A@i�';:0SB��C����$d��e�|�3�[�n��)�'�@�S2�W w;�Q��$��w�Ԙ��2E�q�4)�� ��Ʊ*�(�ȓj�>T��J�9��0�/)mj9�ȓ�`�be���Z}��rfիT�Ɲ�ȓk�8Rm�"N�CE�e�\����W�0_��"	W-X�١�"Om�7"�]ˮlJ��ɿc����"OREF��d��92��%sZ�سb"O$���G��96&���ǇFPZ�1"O�̒��V�}I<U�ā�N98Mag"Op�F��3a\�˱���,�q �"O���a�7h�@�K/.�hX)�"O�@R`���+�@�Y�難SZ��XF"O� ����B�:R�rQ�CH@>$+R
u"O��ۅ�ޠ/�4��0�q&0	�"O~�p3�T�p8PL���J3v6����"O�5��)Y��r���a|<��*OR�k��t�6���W/j"P)2
�'�vCǌ	5�m�!K���	�'���6��B��y�d�.��'��|Vo'*�Tz���w���(�'���bcܲ[L�pAK^*u��P��'h�\C���#D����%��f�hD��'��QPq�ʎ-.b�6a�J���'�(9	D�:wRhbg#� WaH�'�F��1O�]�I�/[2Z��
�'���@e��UX"�� �1L��L��'U�a8�'=#����U7����'�J���&/�H��o�0
�\��'p�}J�UJ�-zU��3p�)h
�'9�4d$0Z��G"b�H��']P��c�&���ቖ�\}d���'5v��nWz��X�qO�)Uؚة�'��ij�A[�^�A&� ����y�
QG��i��̊�"�L10T�L8�y2lpǖyAAI6� ���6�y"�47��-#����su(���y���UI!d�ф1r �D$�y�D�
���+a�� k�4�8�����yZ��i��d�0��Lx#A��'H���!ܝ	�RQš&o`܁��'nԹ*��P��-!%C�+vt(<"�'0蘹%�~�<�˔OX�W���
�'8,9�DӝIE���Um��F1�(		�'.�uk$%4D�8��fR9k�L`�'�Z�	�M7�Q2�BZ=jB
��'���:�cM��C�S1`����' �,�sN6�\��7O��*5f���'�%�Q�Y�ax�l�r�\�'@���
�'C�4�@ga�D�1��	�F��y�G�^xR�2�M�"W�91�
��y�)�jJp:B")�SU)�yh�!Wu��C�֭`��t�X��y"��:��e��""d������y��V�6���Ӥ�b��YUM��y"ˆ�=f��EʢW9�Y)�b��y"�f�������Mi���)C-�y�&	z*U��C6wr��b���y��� �.,��i�C��聭I#�yE�2}4A�PnK��,p����y��L�J�(Ϣ>m��2����y���,��q�����z �Gm�x�<�M��K�C'��ax�ˢ��H�<�G�G&L(�0�	=��0��D�<	s
��"�J�Y$neѪ�i�<��GQ�u����~r�4S¦�n�<����+��#�m�6��@�i�u�<@��w�>�(�g��"���b�^j�<�֮47$V�� ��joV8�@�c�<Ifg�>��s��H#$��i[U(�`�<�m��@�!��!cw��J��A�<��ˊ=x-z	A��a��xi��GW�<i�h�)>�~�i'�K*�ʉ�g U�<1�.��	�dT�f*A�c��A�MN�<A��Cx�i����)�����E@V�<��œ�,ʙ�
�4+����cLUQ�<��ɮi`:���cҨ��"@�~�!�� T����՞\&�#��C�Z��`�""O����aт�ūd��d��]I�"O���%mV8s� �R%3u��"O��Cp+�O��k�-^�1	���"O" ���33��������b�B%"OVX�`�M�tpQ�4'<i?�9K"O.��OJ�^~�]�b��R�C"O*�ѣJ�!7�$��#�'�!"O��+IF��h����F�I`"O��ʲW�+F$��.ɴv��x�"O��"N{H3N�	q},%�Q"O��!ሞ$ .섉�M�Iu��H1�U8�X#�_hW�u����z�q9�!D����%2hr���V 8�B�$�=D�kTgB�cYp#%�S�S����<D��X��ܓRHb+T)�����ruf�<���ӗ:����0A�{jI��U5��#<!��$�O8��+�kP�����6��&;D� �(�*;x����SI(I��U��hO?�$8/�ZR
�=%���1�!�:"�2x�`i�"�4z�Ɛ�P�!�Ҍ}�����B�؃��s�!�?9��X�s�]�y�"� ��6�Py��Z�}��x[0�	uT�f/ڢ�y�g@�Y7	��J��~�m�vg��y�L�g��r�(.n�.����O�yR��=Po҈��,U�5^2i����y#������Uh]5۠if���yҨ
�`-�����bA Y�Ħ5�yb�3_6ܚ�^�P� �,�y�B�8�\�b���,V�����\,[��➈�S��?��%���b�G�؞R
Q�<�@nM06��1����
M����N�<��#Լ}`4��\�@��q�ªWs��l��Ц-�reV�m�r���3wx4	 �4D����	�nIX��2w�Fh���0D�̹WGҷC�,��M�F=�<�AB0D�lS6�O� "H�@�M.|\! �/D����J�-�$e���(XV� ��.1D� 6��Bb��2슨��ԫ�,#�O��'��BGb�	�p,3�d �y���cӓ��'�.5�k[,P�*xiPo�w␉K>�'qOq�$��u�F�-�h �_&�m0"OF�B��DP�� ��2;���9�"O
���-���t���n �R+.�S!"Ov,ȳg�W&�4�[�".Wb�<� ��:9��Àeت�tYH�aP^�<��/N=8�x�0����iz���<)ցU�i�%� iJ���!��mz�<aB��mf@	+���rQi�Ev<	��n�2�74�`@�����1Ϙ��ȓ��`p�E?eJ�*"(ŪR$r�Gy��'70,��	��2{����N12�z��C��8+�B}�rf�LR*yP�`ψN�\��D#?y�O\E�V,&���Q(�4;�X��"O�ywsOJ9W�ߪi�����"O�`�P�3>¬�R���o�p���"O��e`�2G�g��bx$�"O�r���n�jx�gCA}@���'��F��R/&��d2�оGʴ��g�.Z�!��G� Q��d�H����G8!�8�p�Ar�h
�9�@�j!���6-`��R����<d
̐�O!򄝯d|��%eR�%X�`Q�l�%!�!�� ^3��B�I�\��	4x�6MA�_��o�_�'�Q���d��!#�TMP���t�>�@b�0��O�6�r�(r��I�Qͳ�a^��壔�B�!�$ԝD$eZ�b֨^㬴QW�؁x<�{RX���'>��x�J�r���T��3�F���Io��V�X����{��T��׿K&��ȓv\`�/�"F�=a_9	?�%�ȓ3��={2EWG�傗A@����y������gx�(�,H1>.���5��J�IQ;��;!A߃N���/�PA�E��1'�=QUϨk� ����'�ay�H�'Y��Y� ��$� �S`ڶ�y���0ʤ,��4aA���y�ő4;H�up����C&C���O�#BF-շ%��9����))�TY�	�F�<i" ߿�
���$/��M� d�l�<a��P^�M��'� i��Ej�<YQ�	� �#�eM-^P�HU��i�<�㹊`k���"����-��z��D__��Tc��^���BG�G��̅�	�>b8���H� ���C6���pw`��Rn~j�< �(��c��%8a�&e��yB��8[�����g�$+�qb���yR`�4>Ҟ}����\8��g��tX�蓡a�V��x��&U�ѹ�'6D�`�O��z�Q��o;�(KT�1D��פ�$(!H�����|0��/?�
��P�!�MW�\,&��beP�H����ȓsӈ��&�lH��$Q-����.�ְ r
��|Lt@*V�JX\�ME|� ?�'�Z��tϷyT��!㉸p���2i@�a厓rw�(вG	1D��������Y�H��#�#f@��0ReB�<�h��p�/\O4,�=q3�)X4�-*]�vg
ԋ�o�<�����>���L�
�BQ�ŋ�$s�Gr��hO�Iu�
'�D���p#��G[Z	�@�>�����ba�6��p�7�_."
x�*���s���������a@�4lE�a9D�ܫ �\�^��Pp�#�/�d%�r�7ړ�0|�1j��nb(���>�B�:Ņ�Q���'���0i�E,҅�����P㲀�	�'��Ɂ�Q��b��C<_X| ����Ob�}� '����8�a\72�(kW�GK�<Y�@� �0�ar�7 K��z�Ïq�<� b A���C��m�ޡ� Li�<��M��T�v��p�Z,6�B<�Ea馁E{���i���9���4' A�$�
 :x�Qh�'7�5�AW&
�������:��'���ޱ$���Z���}[:T�	�'�2��a�ɜ3ΰZQA���`��'�*Y���j�F��H��
& ��'��h��a\�j\HA!�	:����'��C�ۊ]�]�Ι
��9��'�>�ⶅ�"z	&
ޤ�B���'�!Z�a�z�$`ՀB�z'4��
�'+�%P�A�s��#M:s�`�'��cLv��do�3r^i�
�'�d�`'��@J2E�4�K�g-��R
�'TMA'l�ʦ�d<^���'����Q��-��\�'� P�t���'���Y�&
�n�H�@B.Gۊ���'��-���
�7���:@ܠpӼ	��'uX�	ӓ~��<�#Q�6�0B�'5��R3�/~}:�	���7F9��k��� �H�a��.��͠ �,Zצ��!"O�����;7�T� ǆM�z��m�P"O ��ˁ<��`U�T����2"O�91���>�J��i�%j@�e�G"OJ�@�j7zua�Ɍ�bD�ؚ�"O�ii �Gm��i��9��9Y5"O��)� T�
������hɀ��6"O�%x�-�;��R�o�k�R�2R"O,�2는<����'��X��̛""O:	�5�L�L�d�6g�!A
j�"O�`��s]�4�U25
�u"O���&�h��:P���_�RQC"O��d�IJQ���"O(%��i�X��b���n]�"OL}�#���ęBL��&���"O��R� ��N%�d�����f"O��P��2���[�ǳ+{�e�"OR���@T	 �Q�f��p�ԃA"Od�cl�~A$ִTJ�
�"OI*f�ڮ?�f�S�HH?�$0�'�ĥ����h�ݲ"
��H�X�'���a�,eˁ�:WԜy�'[ 8s�gL�y:���ƅ�+>N���'���a�p˺��
��y�'2v��ʉ�v�,�b	L&����'D�!"�L����I��-3���!�'��DcD-�4�QRP�^<aΖ|��'����'+&�d����ņN�Y
�'<��׫|&�@2���#H�D��	�'�p "#,�z}4��&�W?I"Xy 
�'� #Ӥ�rB�8�6ď�Is	�':L��瀧0t�e�V7N��8	�'VB�rU��`E�HqO���'v~ѣJ߲�x���L+h���'�b��f�ýfХ#��)��0	�'��		$� �A�㇌��ɣ�'�*.н09h�����3A#����'<����M�K�vZ��\/j�`��'�4
��@�1 ��X���!�<�8d���O).��C�IÊ<N!�O�<W����M˃�ݠC��}!��ݱ6�q��·/����Z~	!�D�,I��fK���Dj#�I�!��cf����0�����*Iq!���o�jx A�
�\������C!�$Y�Oׂ�������0 W��!�$�&Qж!�.�+=Zpె�7l!�$�J8��E�:O>�yu�I	b!��9Z`D�!n�)��(s���]���!5Q`�J��b��Y1$�P�y�D�����1���.�8Phȓ�yB���Z�4` F�|`D����y��X�y�HR�@8G��ݪ��Հ�yČ=r��{ab�D֜`���yb	�m�
�����K��؀�
�y�I�1\��U���J��h�`�'�y"�	"�Фmէ��	�3���y2n>p^m"�hU?c�)�х�yr%�H�H�E�%�4���%�y�cS 6V�d�����0hL�yR�^�v�ň�X�N��w����y�IX���)��		7`�	���y2k�)cv�u薏[�z�N`8d��y�g��d��`Xä�<�dq/��y
� ���Ũ�r���f', P���"O�ap��
�n��j�CH{� (�"O||C���+b���E��&Mb�"O�$0�K
���*ឭE&X�"O�1`g/��eol����<6@<	z�"Ob���5+,�՚�e� X֨U�"Oʜ�r��4϶��u����6��F�<�LH�ad�b��:^�ěU�D�<�p�L�J&ʵ��LS\��V��B�<�ƍ��#��'N����`!�{�<��Né+�0�EK�-]�@T`CB�<��^"��t�\�e\aJ4��|�<�1��<H��B�Uz/6I���UM�<I0k�;1 E2�dЗ Z(Y@�L�O�<��Y9^"B�R�脖D�:}���BS�<��ШF;�P�6IO s�@P�<�`�Es�HQ�E;�IAt�LT�<��`�a��j�X6ؕА��I�<�P���4�USwȋ3O���eMD�<�E� .�\�F��B;� 	B��I�<a��H�Fc����,'L��˕E�<��/����������T�"�"�@�<Ad�ӞVZ؀� X�j�$Qy�<�a(^)i1Nty3KRT�T�D�k�<�5�\= G4+�"L�s�D��#M�n�<�p��]� 	bRa� �<e���g�<�@6e�8��w�h�jq+�F�c�<�Ɵ>}�ԃb�	D�D$GZ�<1O�0�����S�\ŪQ��Q�<a�/޺jZ~�VG�SzNT�CEYv�<���9#�x-�0�&�6��TA�n�<Q�-ʊ^�^�k��o&�����"O�P����x�
ѣ��p�QX"O�$PG�� u\���ʟ�+{�I��"O��"�@-��I��Ϻ#^��҅"O�����#@`M8�A�/H$y"O�P򆅗~K.���ʒ�s+FĪf"O��$�Y�qK� B�+�
>F���P"O&��F�P�,��h0��<4��Y"O�������d]��.e�p��"O��+�<�`�8�='����"O�{6!��/9�Q�+�O�����"O�bo-n$͛3�pm�=�"O>��-G�}����)pW��r�"O����pO�y��
L�8�"Oz`Aէ�:Ijz�'�O-@D�r"O���KE�*�0y�p�W�z^a��"O�p��(5��Zw�:WT(["Oꍡ�&�
���\B��"Od����n������Pvt�ɒ"Op�!�,�+)F<k�fwzH�j"O����ǆ#v��7k��]��dy5/-D�x9E�ڊQ���UO��ㄜ0r�)D����%V�Aް$b��F>pƈu{�&D��`�C%r�8��È6'Rݹ�`&D���g�%>ܞ9Y0�[��E�q�?D��t � j��{3˃�Vn�]K�&?D���@@��b l������|����"D��r�p���V�����b,D�Hz��Y�J�P3&,�����M6D����^*g����hB$T��a6�)D��JTE�.|D��#�� �#h`� �%D��30) J���A�G�0�\�Q��8D�`�U�]�m4�����RX̀�`"D�� ��wÞ8Co,+p��tKhDZ6"O6-�q
�9����G�̱`J<+�"O|�a�̀>Tn��j�Ҫ9()�5"Oҝ!"œ8&�*M#�"��+0	��"O0��_�qM,����ۺi����"Ov�X�Dߦ͞�ɗ �����xt"O �b����P�R ��RS�"O����.���GN�5���6"OV��eaR�a�4uy��BI��$��"O�@ꁭ�68n,��R�3u�0��"O8��C(  ��}cA�\�?�I�"O8Ļ��^�zqC�
�]&�W"O�|kO϶a�
�j7e�-\�0�"OB���g�kH�X2DE�P�"O<D��Ļ]���A�X%z�Ht��"O�
�kſv��y{��[p�V���"OLPQ�=a|�kG�ĥ*ٸ���"O6$��Ks
6���H Wil�"O�R�	2qxr�6葍-J����"O�����6��DA"�J(^�`�� "OQs��ʲ$�5igC�s�Rd;"Op]S��m!z�ӣ��"c�x�"O��)�O#@�l�Z�/d�xE�"O6�:�X�~�:�ra�B<~6��P"O�ݩB�I�>�N(���ȠT{ �!�"O<�1�J�h�P8a���gw*�v"O���b�N;)��"�"�jf:]�"O�m�'�>"-q�"ʡdt
��"O�tx�"��2�n!'���N�i�"O�A�M:r[V(I��V2�@e"O~Tb�U>����LV���"�"OʙB���h%�XI���<�v��@"OKݶT������B�P�@5c�
�ybm܎!ʜ�p�/F[�L��lʐ�yD�9#~Ȓ�N?-TxA�VE6�yB��?}h�5A%�F3k�p�F��y_�g]0��%I�<"�Ր�OW�y%P�E�X]�r �%h^!cP� ,�yiD���a1@]�� p����y�&ʓc�� �᜛�p-�gjО�y��O�cJҽI"��+,P�C�@��y�)�12�n��񌈅GLqr��y",�Vz�1�֋@	�� Zsl�;�y"�O�G3|Tb�b�2iqb�8�	Q�y�kY��<�z��=ƨB���y�JE� �1[��¿W�m��g�4�yb灨q��e�e`G���)C8�yE��bK�D	��ƣ@�ּ� ̗#�y�!�U��"u.�%����9�y�韸�T�PE��&+�	���y�#G. ����H�l,`��2�y2@�^V�,ۗ�π==�ᡶ����yB͜�U6,��ėC%���%/�y��޲U� ���	�;5��Y��g6�y�?(b�ݪe
<&`k�b���y� �:��,(D ���(U4�y��m8�Z3-O��(���+�yrF�I!�$X4h;�l��	�yb�ڀ&�R-���\�f����/�y��է!�d��#�)�J\j�'��y2m�J�،B��C� ����y��Η	S �`��HԀ�F��yB� {� @�]���YdEܙ�yR�b�m����F��PQ7 V#�y
� ��%�,�"����	րZ�"O��'l�eZ\ ��Z���@�"O�qC���8-ɃJǟ,
�0"O�pxf�_�>o �z1��G�t"OJ�Z�CZ�4�V��c�&�ac"O� z�

$0�jTؗ�D���"O���`HS�Ob JQ	�$�R�1"O�AYD�C=Aa�碘�"�ReY6"O�����%�H�bկԥV[z|�`"O2 y�*mi��F��*��;7"O���B�G)I�tY��ǠB�M�#"OBU��%͜~�h�4nΏit��"Oسg+�#*M�})�fϣ)�Vq��"OJ�
����8~�X �� �~�9�"Ola��d��!kç5k�1�"O� ���	3��UZ��d�fI�P"OX���d�"��p��[ämZ%"O!�%M��>�m:�9��C�"ODA*#H�-P�l�3��6v����"O(ɸ3(�<c��x���E'[�Aw"O�����[-?VB����NG���"O@��gMW�th�� wO�
�"O4�`�+�I�X��p�C4><���R"O���.\�
��d�A�95��"O�8I���Z'~e��0h9  �"O U�AdD�6�fe
�ט5��k�'J�{��K�P*����}x
�'��TCטV�j�)�YF�	�'�zفv#��b�fHRĉ�g�$��'`�l���F5I�-�D*̶���)�'�Ū�&�0Y��Z�Z�m�-��'rJ%M1t�^�T/εZ����'�ҡ�Q���5r$���Z���'�\�Iĥ##l�� ��V�Y��'"�T�G�ܛK��DX�[�w��k�'0�бc�Q����c�5�'mbh�G5�ɚ���8a'����'"���@I���+��%�$T��'5� `�.C�J�W�M;�`�Z�'�C��@�Q	tlc��� z����'z=
�c� ?���Ń��eMF��'������ �N��!�3Ұ�'���4Iɲ2�8���BI�B���k�'0�JV�
�b-7��e��!�
�'| -���K���kV�
� P�'���pŀѣ^XZ���?2|jH��'���$��)�jE�TH\-���:�'z@�ز�N:
�������
:|�ة	�'�������7�� Ą]�B��@�'$T�b"Q�
�:�(S�Ϧ�����'�"P��M�xn.)��˂K��i�'��,�k���a��(H�F�%��'cv!rH�4� je�K�r��i�'��AR��/�J�5�(dpd`8�'�`�h��u^P�D��k�.�k�'��j#f��7��MH���,a����
�'lfٱ姅fp��bf\�-�*5I	�'��%S�ņ2U��¯����L��'�6�D�ɵUDJhIVJY�(��'��i"gC$s���ť�(�Ę�'�`<�4*�2i�M�5&T��
��
�'�,�i�����TJ^p�&H�	�'Sr�r�����UD�%e����a:%��i��g��z0��5��8��S�? �C�蒄e�j�z��4)��0"Ot�{&M�; ܞ��+�,�@9�"O29�G���i'Ef�l�#�"OV�{P��������NZ��}{�"O,��tjM���Q�b�)C��a�c"O�  ظ\p~s��Ǚi�
dRP"O>�.D�́�!mM�UnH�R"Oz�F%ą]�lT����%z 戲�"Ox�"r≈G�� ����v�(��"Ov�SJ_%V��qB1d̊"���y�"O�y:4E�6�d��aC�#M�(0��"OliyC��
���z�
,2�UU"O��2�O�k�0 @Ԕ!�,4��*O�9��ޭ{8Ba�6<s��(`
�'�J`RAg[�p��6!�'7��)
�'Y �q[�gMv-�� j�9
�'���P��C�R��s�#��X�	�'���X'��D��E<
�qH	�'*�`SMGz�֘y��ڌm��	�'5�Q0�
��R5��8|�,��'R ��ܞ2�F�q�̀f���':8��;+P�hw
GI�d��'��i��F)n������?[ո�'�E��nd�H�2	�18�쑢�'
������5����I��}7�%s�'���խC�(,s�#ԍoB����'�"�{����վ3����A�y��3=g|(Y3��[�PtA/�y�I�n��Ӵ��Q������y�HIj�[��M�Ic��#���y��(�B�;uG%?�UJfI:�y��Rz�و2O�$A��pF@��y�MȚ\�X�*�@�p@ᒭ��y�d�;X�� q�\�?����n��y"'�?K̴�Z�AW�c��Y%h^��y�E�N}hSeU#e��@A��=�yC�Y<&-�@h��E�G�y[9S��m�(�V:�E+�Ꮸ�y�*�	/�D�b�̉�J�0�"w)�'�y2�L�|��ؾY �ٶj�y�K�sJN	�#�#_���K���yr	S_��5B`��[�z@A&P�yEK�VN�9W�6	��h��_=�y�"K��f�3dD��gD�ybcH�1s*Uȱ���5�吴�P�yǓ�^����,W��*1�"��y�c�k|B�
FHW�}�h0cB�y��V�v��/	zwxe�@���ybgٳ'�H|�aDR)<���^�<�F�q��I�1��ve~��(�e�<�`�܎;�����F�C��	��/^�<��&շj[��q��2��љ��M[�<�2��(��E��z���.
Y�<9�fʬ\��S�'�����q�L�<��U�
Ҟ��d(��5�.�؁��J�<��-0Xb�p����|�2�x�-FD�<�_Lak5D*6G���a�Sh�<����y^��ˉW��b1'�d�<a�唕���Nಝ��^�<���
K��z��ܞxܘ��BF�`�<��`��8�K�@�y�X���H Y�<!A��v�&Ѳ �՗��
��W�<-|�UK���@O���b�ԎD���o�4c���
��n	>�l͆�S�? ܩ�J�;5Δ۲��:.<��u"O�mٳ�W< �mrs��[-�a"Or���wN)�BJT'|�D��"O`�h��J81�B���c	,x2@@"O�1Z2��?��A#s��:0�y�"O2Q��)�������kF"O��S�"MB"0$�$m�P<�Ybc"O.�(��o��LS�U:0f�"O(|	p��?Pӊ����	V����"O�� ( �V��W*�z���"Ot:�?W���r]��9u"O���}�l�ʢ��1TJl\��"O� �!��8a��4Z�M�i:�,�"Oޙ��J=���䋃�{�b�cc"O\TAw@]	̼P�c�>!C���a"O�h�5RL�a.�?A-�9�"O�͛#H� �!8�#0{2���"O4���JŐOz�$�p�ʨa��d"O�����,k.�=���Q��D��"ON���4
�����-U�o�^ s�"O���P�[�P�0�(�_8(��"O��Y���z�Eb�U�@u�}�"O���c�r0^���ЋIr�'"O��)���q¤L�D��0zh���"OBW���,�p�D.̎M �| �"O��	�)Nq��q���zp"O�;A�X|���bK��y�R�c"O<�3���:*�謲�HWd��h�Q"Of$x���Rά�3!�������"O�qU�F�RPh�q�j���,��"O�hhdV%h-�S@g�� ��"O�w��5F�s��4^�@�J�"O�]�T�DJm�m���`��p��"O��ل��#�<�h3`�s��[�"OF3B+�pLh�	mb�M�1"Ot ho�"��P�r��5=n�"O�:4�R�"�#c����b%���yR $��jTBȌM4�h@R��y�ܰ*��xڵK�5u}Ba3r���y�@�(DX�C�8kr�	A�̑��y��V�hy�AH�U�|J�#��y�
I-/�b%瓂>p����o ,�y""N;*�@@�Î5��H!3� 7�y���XD��{v��/<���a�i��y�DL'3qV%ц���8o2�(���y���:�ޜn88�>��Q�0�y��S2�j��՗7��p ���y�	�Y�䬫&�˱3&������y�OE���(x�k�3�Z�XWoH��y£���	��j8>��+֨�y,�2��Y�D�%���æ/��y�hگ���hb"�;}�\|�J
��yb��#ԉR��ɾak�<�m��y���	Q���bQ��x���F�*D�����0<r��լXGt}��,D���#�Hu����$���z&Dܱ�*D���� _�W��)� J79��H0�-D���T)EJ��I�%��	��(D��B'�4R���.��,w�U��'D������ra�W��(p�`�� (D��)b�Q�8����ˣ7KZ��J D��X��<]�(x�nE�F�k�#D�D���A�}�2��WH4U�0M��)&D��:K
�p�+�`�yc����$D�� ��'�ҍzJ\��D���t:�"O�9F�����K��	�7��R�"O�x��2���$n�?q��
�"O�@�'��+8X�%r�/�5���A�"O$|�b�SI��M���#!u��ӧ"O�0M\)Rg$d(B��+~��M1%"OD�8d��tZ�i�IH���D��"O�8��\-^�`��T�\� ܺg"O����ֻjS�4�#�6�,�QA"OPM�G�k���R���E�����"O�9�&-W$!���zp�C8cb(�b"OrDr�BO<TU��b��.�8�y�b*p��1	�
��,�c�E �ykWI�����c�n��MY�N��y2�/;���Q��ʁg��H�' ��y��3j��������^$k���8�ybΊ2#�� 4��9�xq����,�y�⎎7L���!�"4�	�[��y�O^�RcT� 5�՚) ތ�g-���y��<-������~xZ�dX<�yNՐ}�����I���!�7�yaQ�-�Z����4�fY ���yr�	/Tf�5��vb���Α�y�hۍ|F�a���G!I���֕�y��D^L�4����`X�:�y�h�?�l��fB�θ�S̖��y2��s�P¦��u�[�H���y���]#���F6>' (;"#M��y"!�,/	P����,*:Ъ�#[)�y"&�s���9$'vE.�D*��y�֑~����.XK`x�&EV��y��D�^،Ԙ�(�?kvm�w,�>�y�%��M�������y	���v��y"�T"w� ��Ԣ�r�"�	���ybi�Q*\њ!��^��a!E`O��yOG�t�D��Ћ�W�l�{�'���yr.��_�H	���:�٣`+��y��.i�n�b��%��1�'��y��*;.5����` Q�N]��y���7oI=sq�-bN�h�v퉉�y���Irl��!��!��dp��4�yBlD-� �*G2Ϥ1��.C:�yB �&~)���c��oL�����!�y�k�9"�R��a�i�伒�cx��'K�bW�x��S�-);�*��a�%D����K;~�d�	aIV�*&��@%D��
w*R�pP. Y�`A/h�9:@!D���Hʱ�rw�^�r7�mc�� D�`���@�I7�T�Fi��
~)��f+D��G�K�0�Ж@[+[-���&D�T�%o�8�qa�ձ+��eT�(D��[Em�Hd<���:!����f�9D��j��71�I�#�R�Mf�He�7D�T����0��X�M#t�^iZ2o:D��� nCy̨}��L�W �h2A;D����٪n<$ͨ��C�M����6*O�՛&N9
0꘹a��6F4�F"O�p��*��m�`�K�==�1"OƵi�oLx�0X:�c�;{0ɋ"O��S��˩�2Ѹ��x���kE"O�k�(޲(����(���sg"O<X9 ���T+��za�E Mk�5@""O��:ԅVf>,,�@�����sF"O@M�p�ކm���cTiDZU�xi�"O� "�X�cB�"MP43�IR�5O~XcG"O��ۗeYZERQ��Gŭ38VI��"OPE�c�^�#��TP�&��W|���"O�8H���"Iب��B�cc��`B"O<!	1��.��D�C�)����F"O]J�Ǝ�,��i 7ȅ4�0%Ra"O��1q�[p�p��U}�fPB"O�ЁgԿr}@��C�� w� �	"O�abfԔm�KubCZ��	��"O��@F���B�qq��Q	.I9I�"O�إ�֙y�t}���?sG~��G"O\2�(P�H)�r������"O���e� �C�@�����!hN�T��"O���e&=��3��8D��Q"O>��$B��a���3b-נ�y��H,"���(0!Rq��ɇ��y$��N�L�j��Q�ڼ�򦒨�y��+�5�&
�>��HUK ��y�)ߊ;1��薃r��S4���y҅O8xJ	eA�h/�:Q-S��y��A:B�<���LK�*�0!�� �ybcA�D؜0��$M~�|rQ-Q��y�	 |yb����E/{켝 Q(��y��A�2�5�FL�"m�j<�G�;�yR��e�B�k%,	9���q���y�'�(&;��`QO.4?��	����yB`�]Z������=%�,�CE�B5�yBm�i�pC��Ô�^�"�L��yb�� �����.M�f9�yBo;}�`=@0������H���y2"���QY��D�{�VAbGH���yB�F��(��Ώ!��҆G��y��ՍO2 �cM�Qh�R&��y2X=_�н�7C���n�Е-X7�yb�wPQZqƞ�G`��#Ή�yB���QK da&��E��԰',V��y2��0:�Tq��G�%�HT�V	��yB�F�NDl�����!��[�&�y��zI��pǫP/M �pV-�y(���X4x�l���t�i�"P��yb��B�l�A����t�6J���y�)N��8��Ѣ}���0sM�-�y©�� �ti�K�(}��i�ыZ�y���55��C�W*xҨ-A��+�yB�Ό(��T)�D�̭���=�y2�A%220P�aŖ)�"=��!�y���r*�sr��wU&��u�Į�y"cͬ��*"��&"���) �L��yR�P	��`!�M�k�ǨI+�yſ 1 nL�{��R@+A��y�BvR�` o��z0�Ӓ`���y�lJ7f����p&�����Q��y� Eze,,4�B�lD�1��[#�y�O�Q-(�a"K�]�LiS��Y"�y���/mɖ �dL�dz�H��yҨ]'a��9B�O%y��x��ٸ�y�L��{�@���I��Hx�uP��̚�y�&"Tb��-C���a��ٞ�y��ƿ6!��5��d�����&ԟ�yR�S�<]��x�j=X��,�"� ��yBǟ7&~�Ee�F�Zɔ|�������$�<����h��ĝi\��ydG�"�)Q�+%'�!�dI/DT��3C˙I�>D+��ĄL^!���NqT�4��!o&��R�ˡm@!�� &��wE�9�̔�b/B�T��Z�"O>��U��g�|P�n��D�z�"O���a%�#�:���
�ND��"O�M�C;*iC��T�]~fP�"Oj�"�g��i*N�B+Ŧ!�����"Ob)y���{x���n� �I�"Od*`�\�o�а��Ix[�\y�"O���M�Rq�Q�W��>,D�bv"O����Βm2 �O��'% x�"O��B����=R��!D���D"O4Y��OU4\��	�s���h�^�P%��F��'̈ˠ�� �ܑT��\�x�8
�'\�%�#(x74�I!�L�	`�'6`�"Չ ��Iu�iI��	JH�<)pc�?s�
�'�Q�h�R�WG�<��n�2�fx��H�-sb�1@a�G�<�T��i�p�:����kz=9u��j�<qA��<f��u�V͛� �P��*Qyb[� $��|�5"����sŎ ,y<!֏�t�<��#�a�LВ�ܳ?��0����z�<�����D�F#@�=��=�hZt�<qa�-�1���.(���)��s�<q�J4j{B�b�
�+�� "rJJ�<�����g�Lpsb��#xo�4p�GZM�<1�M�6�"(�n�8Z��5�MIpy2�|�X��Fxң�*AϤ�3���Zy
"�II��y"��b��)CF�}Q��#���yBO
<�$@"F�ȴIlnW��HURB�	7v��T! 
��=� 85a>'`B�4ej�Z�ەaB�I�@+B��2B�I�$@�K$$�H�@yYXB�I/j.~6		� �G�� !�$
�h\�:1�ƟNƊ���I[�!�W42����&���T\�Ү�l�!���P��a�n��>�	n�+v�!�Ds^�`�52�vP5���[�!�D�'D�yC���%>V<1��J�0�!�']���[�;&a���.7�!��T�x�����!�1KT
uH�I�_�!�D�6
��p�V�L4[P3&�!�d�]�D����Ú�%J�T��'��� ��7N٨p:���=S�d	�'@�e�w���=U�ę�i�N*���'��%���T�rM���!D�	K���'��sB,,�t���^6
���'�4�����#e��!�(�/�ޤ�R�'�a�t#ԋt�q��'��.����կ��y)ԙ+������
-Se)���y§�#B�H��p��/z�0�XdDG�yR��+o1��Q�Z�~������J��y��K'��#"G�t�4Y
�B�y�$� �X�0��M<g"Vx����ybU�c���cq!�%M�$� ��ա�y�m͊gqFY"#ݜGx�S&%Ś�yb	��Z��	�1���z����y J3X`q(��Y|�5�ӯJ��y��ݑޚ�	@���N��`��-^��y��Q�%j�11�뜈e
� p!�$�o�h����TJLA��~�!�¯x
B������Rsl	q+�7h!�WX���p �YWڀ�U
0 �!���Ay\�8�BB�}�� ʦ��L�!�Z���"����4��2�A�#~'!��ۖM�������J��H#rl!�� d��G���B�R"�{�^���"O��V�����Z���=����"O\�C���2�3t.��l�T�b"ON]�O��38�Pm9}�DQ�"OmP,�+9��Њ!�Z n��t�"O�p�gbߚ{�N��2�LL_�"O9��언�L�ەQDC� T"O���C�_��H��!�7:΅��"O���tbٷ�P`v͜w�i{f"Or�IA� ю��4��H�d;�"O�ԃ s�tY��C�^���+4"O���E ��%�g�95 X  �"O�����ư&�.!7��=<�֩��"O�pHBń�M+D����-~F�� "O��X���?nT�!��	�H���e"O<Q�AIHDʔg�5GPE�"O�3	�tD���剀=j�|aX�"O<�G�R=0ɮh�Q��P "O �e�Fp��ȂFI:ݬ�f"O�d{��9R��x ��$�6(*5"O�q"�͙�Fǀ�l�0'�ܛ�"O8�B��;s :'쇃|�0Y�"O^1`իQ7ty��YgKHnd�q��"O�|@���[?����q���"O��ao٠PHLQ*���#_O^��"O����62�zɣ�c'��"O<M�%��
-�(d�ѢT8I�M1"O$M2�勳~�J�z�a�5����"O�ax�S�T�RFK�!3��$SW"OF(򧚸'���1�W;��(��"O�0�G�F�5�V���'�"\"�`B"OƝS�5(MzV��E�ۡ"O��!"�=hՠ\ C�?;���"Oj�W�Ŝ�B��	Pu�"OB9��!�= /vY��F%B69�"O�ԙ"��BP,,aÆ�Y1�q�"O�(p�
���&!� ,lt��"O�T��i�2~�:��2凄jr$��"O��C�Z=H��#�C����t"O�e�7չT����c �:_�0�i"Oz�S� �q�l\
v��&�^��5"O�(��@�<^��P0.�<lp�ؔ"Op}X���=���c�4����"O�0c��-{-���c2Vp�b�"O�)�)�/^�8��c��9��-��"O2�Q��Q+j�Z<�B�A�/�
	�"O�8 Sb�0j}r� +E��Cd"O
DC��|`PꐧGÊ-:q"O�c�%��0e~$h���P�*�0%"O$%B�9>�0�q��Eq��@e"O6�Æ���\1��9�Z�]����"O�P `�_j�^�˔'�]�4u;�"O0e�@OO]l�LYBe:Ax0pd"O,@��$A(F�QK���+J�cw"O�LC�DaQ<Iڀ�M���)�6"Of01���*�xP�aQ:L/b}�"O��G^q]�tBt`��$}�!"O�EX �Q�Kwpd�Do�;��p�"O�=bW�%k#�tmȲn��EY3"OB�u%��<���8�K�=pz����"O$x�6�Z�>�Ɖ�]k̘!B"Ot`�/�T�h�[��v�A"O��8��OkX� a��1?�D�S"O���r&�6^-rM����h���"O� ��xD�	{��A: �T0L�"O�#�Ŋ>b�vM@S.�ZΠ��"O�=�N�J�`	j�l�?sYb�@"O�Q�ns,�w�
2&\���p�ȓ�x%��J�;(d�"�6|�����%�a��N(bZ�0J爓���0�ȓH��#R�,K�Y���W�r��ȓzN����F�+'�T�k� dn���x��Ҥ�*��pcE��Ն�g`btQ�E,|�p���ԋY�)�ȓcyl �(:�H� 4BZ;����{~ez�-�-B4���?@[�I�ȓBD�����$:?����E�0`?�ȓc��P�E)J!��b�遳�݆ȓj�*�(��P,J�L�bgN_2wRĆȓ������P m�R!���_�आȓy|�PWl�s�ʜA�㖒/Rd̅ȓSŎ	"�wB��$J�p�ȓ>���v_r�,���]�1������M�Ňɋ]���"���B/���ȓ
Ւ���Z�Z�A�n��
����ȓV��H[ ��J��1SN��:慇ȓ?��`ۇ�Ϝ_k4�1�1$�b5��k�vpx�$D<Y����h�d5�ȓ�h��RM(�X��_�*���ȓdf��ӡ�Y�NH�e�2��p�ȓ{�0"T!}zmд�_�:��K�r��ͬ>@t�w@>"RQ��k��$�fI�)7���A�h0���7lpA
r��H�,��.*����ȓ\t�9ʠ-�<P��ab�ٜS�����G�TT���,S���!��x�6��ȓL��@���M֨�Ъ�B��ȓW���"LW�ʁe��Q��d�ȓ<�ܜQ�K��zH�� D�8
�Q��0S�a���߈3���4�B��Rф�$(��C�P�� �Ƕ}�����V��u8�O�&Vu���4��2}���ȓT{�i�#��@���� �,����󨹘'@םM�� DcF�=8��ȓ*�tas�Aϑ ��4�
�K�ه���k���6*�@��-O'&V��t8ꅩ��E�e��*�D�]�nC�	��f����Jy��GI�'URC��)�h�r�#��{�~�1T�-N�B�	f��RSj��%�FP"A���)˄B�I�BԆ����H�`nh���;I~\B��t�FX��
=SG�l���ekRB�	�X�
Q�̕%��I�k���jC�I�!��)��Q���
�Ú�9�\C䉠T%\ �`�ٟf��챣mX!J�PC�I�����J��n$����<�~C�	;u�麤B<V�;��� C�I.}���!��٠{����A_�|tC�9Z(�t�V�sS���<f��B�I9QX�fN��Y&�:�NQ�\B�	TI"�H�/���v�ȿ�\B�&`����b�ϚR�xL�!2�*B�	%!9�����Җ`�x�v �K��C䉩Mkܔ�d�C�Δx0wdI�;��C�3VsfY�󊉊`�@�jf��=XB䉾U}�{��<B�6IY7�B%E�xC�4I� �q�E��(;ٲti�f�lC�	�WC�pc�%ʍ2`���D��e��B�)� ����C�J��)IdHA�*�v=�%"O���/�p$6j��_�
Y�"O�X��-	F߲-���X�d�@쀆"O^��R�L�G$��Ҧ#�@ԓ�"O(�q4��,0t�3�%�����"Oи�C,ϏGd���z9TG{�<i��R:2���Փ6Q^p"cJQ[�<�#^�]D�t�׎/r��z��a�<��P�"�X�♕L�d��f!�\�<IrjY�-�`�D#�$^j�$�P�<��BU"Ib$xe��pR��DÌO�<	���qw��UO��*�r���`\O�<���[J�xEX&�EH��Y���L�<�6���vT����dZ�ȥʜM�<�օ
}nAҐN�.5Eh��G-NJ�<�&-����Ҭו:`��S�D�<y�cȏWӰ�ca@'[4��g�j�<�UN�u|��b�����b����@h�<���Q�8!l����F[���R�N�<�w� �����R5N#��z�͘_�<�D�Xl�P|�҈0G��q+ϛ\�<�QAE�>�.�A���snt��a��a�<!���/Z`M� l� �pኅEa�<����3|�9�U��G�H��o�u�<� ;r�ji2��H�s�*�K��0T�t�`�Ԅ'�����5[
�9ᆆ9D��s��ë
&��R똩'EP�0V$8D�xj�I��cĂH!L�IRD���3D�dk���.6��%��P�D�*$B&D�H�i�4Y���ҫ/0ޔ�@�7D�t��π)	f`��iһq��]� 6D�()׈����ɐ2K��1W�U���>D�|��ǀ%����Eړ�&����;D�X1a��u3J[ �[(G>��6�:D�<���=g 혗@��
0\�D#D��weI�} D�o�lB+"L)�y��́Pwr��w����S`��yB	�?���h�l���'���y�9.��y�W��
(8P�5a��y2)̠Ow\��e�#t>x���j�0�y�'J������		r���"�y�'��1]�\:�
� g���٣���y­���m�E�_�-���q,��y���d��d8��G� �^��#���y�F+)��q�7n�
H�,݉�?�y�O�Cp�$�ggS�l���y�(��y�iZ0,6�U��)A�a>�ȫH�yRHR�$��Y`�F*X��5�o݉�y�I�T�TQ�R�%�μ��j:�y2B�O�� �͒�J�x����y��@������ l�<ɲ��G0�y�R.L�L�aaʗ�Q��  
B��y�{�����2��yCi���yr ��P��-]�a��8E ��yr�Y%Bg��j�×���*%@�6�yB��3~���Q9����	�2�y��O5���%�R�/��`'G��yBi�7K���#�&$�,i�僋�y��?D�XM#PY<�h43�ܓ�y�Z�. �DJ[]�Ē��Q��y",Ǐl��j��D.�hvÒ5�y���\7�5˖��5+�]�uOZ��y"'�))�Dy�h���&L"����y)Z�qa��"faV;Nth!�߇�y
� dd`�nI0�:��
��3�B�"O��rb# �*aj�7��2�"O\�x�C�^��@� gƊkg��"O�I���6z�����'F��"2"Od�m�9ט��:8N��"O~�:�i��i��b�&)$��j�"O&}�W@̄T�B���S�X0j5�"OBA��W�F7,��Bmĺ('�I!"O��a�A�,�&���%>���"O��K��G]�ր�g�f$z"OR�F�<#z��!�`��lڒD��"O^QZ�Ů;���r���3�0�*�"O��24@.���f�N�A�خH�<a��BN��v�)�:�gWg�<�ɀg�(�Re�#�NB�.�e�<���Ҧ|H�i�\�-�4�+�c�<)"�M@9 m�AI�|�I�o�v�<S���w^�Ce��x�p��CBq�<���.J@�KP �ݡՆSk�<q�¾NV$}ٔ �A�������e�<ir�D�k�# �@i�@R�a�<)�+F���9C��>Y	Ę8e�^�<A��6��҂h��Z�`�"N�U�<����%c�V쑳*�>Hm����P�<�`�ݳ�̜Y�(6*��=�0�AI�<���ցhU�T B�0 p��i�E�<���ȨOVr����J�U'(�
���F�<�cş+��MB���Y�gH�<���o�1)Bϔ6PM�� ԡG�<����.E pY��yI�x 妋@�<a���!�ԳtG�it��v�]r�<�b�*�̥��̇�К��Jv�<��C�)\8�m�3�Ĺd3��C�
�w�<yԎ��\�P�I�+EQA� �]�<Q �]{��٢SgK�P4�V�<!F	�4ClpiA��������R�<�$�R=#��"ƗKk�t��Q�<�bN�u�����)�f����HDI�<9��.y�
����ҕs&$u� h�B�<���&H�!������p�|�<!tiF�]Dʐ��&�/EN�T"y�<ch�"/��Cܭpw��D��}�<1F�Õ9L�2A��'wL��h��}�<� @L�jԢ��)E��w�<10�˹��4�q�ˢ0̢���fUN�<�/Q-52��, "��L@-�Q�<9�)ˍȸ�ڒ Ѐ1O�͒��%D���- x�l�+0k�ULd Ra $D�Ԙ&� Ug~�ڧ�yFZ���i!D���(� )�yǃ��-SV0��4D��F�m�: ����<'����1D����� uf5"g�1V�H�p�<D��j��&"x��c�%R�xp���C�7D�Ȳ"f
$0�D�JA��
T ��!�B4D�`k5�˚<���v��D�����3D� 때X�)N-�`�XN�:2h1D����$��D�
TDL:��/D�:��� Y�����\�P6�3D�`z��g���mo�2�yD*0D�H
v��l� ��)X18�Fd*D�!D�p�$&�a��<�#Ղ)���s�$D����fF/s�:�B����� e�=D� �?[��2Ta��Q��	���9D����(��jr�eS�X����S'6D�� �;CI��C�6��e�׬Z#$��"Ov���T%eN4$i���8���q"OX9�e���YAlIt��0+��;�"O��[�R$PDT�$�PJ7P�Q""O0�r3�G33��da�̈́$g���"Oj�
�	@��<�5\�E$�0 "O�1��+ۺR�,x�jV�kr"O�� `�ɒz̲�zsI��r"O~L�l�6��(C��Q=$8�2"O��BdĚ'4NP�a��)���i�"O^s�[�4�6챒-
7A��E"O,i(�I�����K�A]�9��2�"On�´h��c�^� q��?$��"O\�1�5����e ��_b��3"Oz�
�FF�0����I�2\""O��!-QK��H��oK��l��"O�R JN��r��I�>햤�2"O���m3BB�3U
H>� 9f"O�ƬRl8�1fHŅ2��"O~y:2eQ�V�R��� �:E��"OZ9�>�ܹ)��m	@q�R"OD��e�O�6�V�V�����)�"Ov<
�+�8?��̀�O3��"O~�ð�0֐��G2K3����"O�� �W�8hx'�G�GS��s5"O `��'M�Y̜��^��:�ra"OJ@��y�8
KPɄ9y�"Ox���"j�(�B����"O^C��%�L4Y���	%�pUB'"O��X �޽gZ���J9����"O|]I�L_9vN̅��5	aF��"O��� 0w�(� �H���-zs"O��)�+T.8�IR�/ء��(+�"O�-hs.M9�&qQ���@hh�e"O���u�-}�8E��T�s �Pȷ"Oh�b���2T����b�|�Y�"Oh�x ���S��i:P�X z��DJ�"O����,�TP�	��D�;�޴0�"O�t��0��p FR>Xa���"O�����:�r�D��qOVT�v"O@-�t����������_:.��"O.E��B��K�h�3��0���""O�a��M��5H� L�Ut
t"OJŚFf��I5��ᯄ�

���t"O
����Áq>z�XP;���?�y�
U����L" ��pe��y��
62╲�K�{C��Pǫ�yr��;���O�B(d�L\!��'}ў�Oi���A��2) #O�.U|����HO���	�����7Zj��"Oɫçʍ��djA1YI���"O�a�2cS�0%sI�F^���"O�ؐC�?K�&�їm�
޹�t"O�awkP��Hb�[1R�ؼ�p"O ��A�M'u��t�ԉ*sּ �#"O$�`�DD�.a`t�vF��k�ք�w"O`d�J�']����R@	�2��1�"O�x�� GT)ن���8"t�q"O��	R�Z��5�j}���r�"OJqQ��Ѯ +b����D� A�%�y2�1Bd���JL�δ��iT��y�e�-l��xCa��2?ݸd#��ɣ�yRk�$&�R�1��էF8�zW*ܛ�y�MP��]1���Rz90�焀�y
� �,��#�#M����o9��[�"O2I� � �=8�x##�1����"O�a�C^Kzr�h0�ؠi~ *3"O��q�7I1���Yz�"O�}"diڀoi ��7o�&��"OT���-cp�d��KX�>|��b�"O�I��D���Ij�=�0�u"O<[ք�6���V�2Rj���r"Ova1EN~�L��1'�aPp�8P"O��Sf�<�u"2˔�"���0"Obx�A-t���C�?��E�"Oxe2���,t���V/�r� V"OSQDݵ^���d*�n�Z�@#"OZ�����>R�����
,���Q�"O�<(th��TC숞��p��"O@%����d5�Mb%d�>4��0�"OP�$c�m�ґ鷣6+��@E"O�@�C��ZU@u��7(l@�4"O��a�L�HGTS2B�-S$E�"O�����
a6z0��!��m3"Oڙq�EV'{���ӯ�d�Z\�"OH���nE�'��`�;�ht��"O�Z��	��L r�U,M�&DQ�"O`���*�'��;beߢG��]�R"OB8���M~��bw��j��'��$_W�	�f
��	�̎3w�!��"�1�(�@���g,G o�!�ǄIP���3�.7F,qkJ�z!�
�&�
<��Ț�K")���I�Zr!�DɌ&R�s�"@'�6M���ӼuZ!��7 h�]�F�
"P��@&��98V!�Ռp�́өG.ze�(�W���0T!�DC�;FB�)�A�~n%&��kF!��U�
���1��ȫwj�I���'HM!�d26:l��d�d�`A&�1hS!��2-�ዤ��WQ�T���(7�!�d�5R)�7�� (h���eb{!�DϠ`晙v`�	v�5��K3Nx!�ă�q�:ݰ���YĠ1�A�/?t!�˺^�~4�V"x�����  ~!��
&��u-�d�\�I��C6�!���H,�=)�H��T���BU�(!�Q�n:"�#è��W���@Ё�R^!�䌯LZ���ܘkX ��m&)t!�d�)(�BΎo�V�P.��HO!�ą�*HFU��	D��I%�ɽ`1a��O���A-_4(�������z�"O�̨��a���7�?`H�@"O�L�$ W��Qҁ�<B��"O��p�ET�s�P�s��Y-�h��"O�J`�B�Vs����m��nh(B"OB=��N�C�~]K0�3m����"OzEs/�� 0X����ĵ!��e1�"O�5KWCկ� Ѡ�!�c�S"O�@v̍�ݒ���JT.(��"O�M�FƞKG��ʷg(T�`��"OH2)�	Q�U���W<��2C"O�њ�,��c�:��0P��"O��k��	|�)#���j��"Ol<SW�D�  ��`ŏL�s��$5"O���G�-L���� د+|Z��%"O(0�����E'����(�g�����"O��Z��D0;~\;d(�!Sy $[c"O�X7+�70)0l:Ӥ6 �X��"O� ��J�b��)��d[���̩""O.���`�3{��]�%�9�~�[�"O�
#oC�>	�U�P�3<�|@ؔ"OA�G��:Yg��d�����"O�Q@6)^�MAjt��"�6]�*aq�"O�� Č~��4�a;U���(�"O.|@v�	�U���sBO._��u��"OfHAg�Ԣ0�j8(� �e7~t�"O�p3���3w���c��3F��U*w"O>p"V�O?L,�5p� �*|�hay"O|�� �M�Q���	���<ȡv"OL�(�(P�K��� �(�0]cn�s"OB�J%Y @���@6Aׁ�^]*�"OnE��aQ�Hu.�	��O�B��)��"O����D�_;���VM�0�N�B�"O�0µ�G+MqМ��M>�फ�"OT��ΣS%zS�nH0ێ�P "OxY��M��Zd<xV"O](��T�Ie���������"O\�HbmT�h_���hPv��LY�"OdV�1'���\"aҐ̊�o�B�<F%A&}ϤE�2@B�*�y��S�<I�cݗ	8%�a�4(ж%B!�P�<�5���bI,���#�\�5��$�M�<�c��)�|��!�5`"(�QJU�<Q�a؁?�$u{ŨG)e.,r�.:T�$�f�^�}v�����\�*���"B:D��1��\!u���J�*�Yr�d1��<D��	��� u�̺'ma�pBc0D��c�)Ҡ*���}���:�,D����X� ��軕H�k�^�V�(D�H3�O�,n�a J�8D��S�+D��s���^8r5�S�_����(D����b�?H`d�˒��уS2!�I� ��U쇐mx�ъ���2t�!��	�&���G(��[i�)�!`Fg�!���j�8�X4�X#����'�G|&!��4M2 ��ٔ+��[b�W�'!�J)w�&ҥ���d*�M
0K9!��P� \�t�[�*
-R�I�,!�d/zaʹ���(��)J)M(�!�$��E���a 8�V B�+�!�˖L��0a��]#��#�/�ct!�䔍 ��T�[�c�l=3����Py�
�
H��3@��=��b�iA��y��Y=�N�u��;6<Z'
 �y2bI8;�$�[0ǶF�M�$��y G�6z�h�� T*��8r�P��0?A�� 7\��u�WLXL�NJ�*g�Ik�,HU�<�u�-9�R(`S�S-z�8�Qi�V�<Y@5}�$s7B�|�6TB-�Z�<�FH� OU(�S69^X}["mP�<9�$��-��K̳\*|�` �P�<)��4w����d+q:�����R�<Qe'�&���CA�K :�h�r�N�<���4{e�\��d�l����D�<��F
��� 2�K�3�F)#ea�@�<Q���u�D�R��3C`
R��I�<	�/B��A�!���,j�!I@�<��h��q�ZQ�-C0D�ɠ�Gi�<Q&�wi�d�V�PI*L5�w)J`�<a�.��e��U����Y��`{W'�_�<��/w�=�ƥG�Fbp�B��LS�<I%��U:��p��<i&L-����J�<� Fp�v��
W���w�>:�2䋑"O���kM��H8c�H�N�^��"O~�1�kY5l 0�gJ�"���#T"O0�s�mQ!,�F<��)�%4�H�Q"OZP7\�-˲E:��ͬg����"O8U1!��q�	�W�:/w���"O��c�d�6-V��_e���"O���d?l50���h��B"OF�+������-�I�� G�U
f"O�3�%X�2(0W���2�p �v"O\Ywo��VjH (��[�X5��"O1i�k��Nzh�Fҭ/x�$��"O�l�o2p���"+Uc���E"OzԢ�c[;_&���/v@�(�"OĻ�ˇ*@^<���='��JV"O(}��BS<�D�A"Ɏt���*"O�ܑ���� �4ա���9A���S"O��j`列2�Ό	��ɐ+]bHX�"O2�ۓ��!w.|�4fO%TCT��"O�1h��B<nۖ��%�W�D���"O�Q�]4��jG��-/�`"Oh��DV�OSL�JE�E�Fl\�"OPx�!�Òk�&Uq�� :츥hA"O
	��H�uMr�3��2�t0yS"O~Tba�>]�(��J�7l��ȫF"Ob\[b����ѳ�HF�t���R�"O�y(��C�*�X�'��h�a a"O*��S���}�h��kְ=D��F"OD9jaA�B�ȅӆK(;NP�"O&�Y��ړ:���0(�=Z%�HY�"O�|#h�-2�ВAn��Ipx�q��'3�h"�뒼k���z�A-n�t�N/D�,����0�&
�.������,�*�S�'j ��n݇T@���J-XCɇ�{��ĸ�d@Yh�*��%H�zT�?��05���\3pq��s2`�:�����F��e*�ƳG;�$�ߴ=�ΡQ�'ڹ�ìZj� ��&��'���
�'�P��"��&[��5��HE/b��Y
�'

�K�tY�"f#}*T	�'�1c%j� 욶H'�Pd�'���!�J��TW�rf�J���j�'���4l�v�m���(H��]��'W`��S�7t���8C&J�2�X8��'Wf yG'��P�H�9�*�' �`�"�'�(�r�(��%�d�
!��;�'��z��,C`�꣄�"�r$��'9j��(�j�u[ �O�9!�'���`�dP�l��X���C�	��=��'�������t�FP1/���^�8�'60�� ��yh���i�M����'���7��	��0;h�q�y�)擡8"�Q���>$6	"!�
�#� C�ə.���B�lQ"DO�����2B��B��;
Z�\�$�P�e�pH" lB�I�)��!�"�'��3��C�2l�C䉭p%<8q�F��M)���?k��C�C �h�I�.B��0� ��|9\B䉺-J�ujQ%��>�d��×0tv�B�I&l���I ��*�f�Qw��F�`C�	?R�쑪�AK�r86�ܕ%�JC��\���P��҅AD��"��(��B�Ʉ/ńU�2M�'|݊ �V�2�B�	���DkW#��-)�X���r��C�)� 6�r�.O����d�u��=:�"O@�j��Z�Vf��E�&��e��"O����k��i��J|XI�"OZʑ�5[��|Sq�J�G����"O����J�'!�ܫԭX�flT���"O@� ���1pRZ���l��y��P "O`��� Q�j|���3J�lk6"OJ�j��,A8|d���7�h�"O�S"���K�2e@���(km*���"O���Al]�W���iɡco���"OP��"O6t���"R�,z"Of��	�S�v�!׆׶!%�r�"O� ��o�n�D�ֈ�ZfU��"OȔʗ苨k TX�ƨS6����"O���4k�o0d��ƅ��Hh�3"Ob��'Y�q�:X"�%�J�(h�"O�qu)�&;`�Ke�V��P�"O4�EU����`���]e8�J�"O�M����"&!�8T��QP�I�B�IZ� F�4.O)PpQaA�A�t�%��1�yrJ�em��G�8�~��lL�?Y�fA1	����W���2h)r��j�2`|=aK�?�v�ȓM&���%L_4)8L,+&$Hn",��t�'��M���gE�x���YF{��#$��"ѮY�K��8�����0>�g��\�.h��k~��${��JHa�x�f�,֠�w�̲������ �.�6����:W�@j{�O�8s:�u$�46$\�U�.j��˫ �ֵ�B���/9L�a�n�m�<� N_��]��A8k1\A�S.����9��$	X��Fc=�D���	���i��9~8[�P�J�y�D+I�<Ѷ'��X���ZF%�	�IIo�x�$=�}X$���s��PЦL��&���H���Ѓ\r����ǰ�@�S��/LO������s&�5頧��R0O
<R�P���ɁA�\q 	��+����se�iޚ��|��:S�7w��%¥��b�����$����w��7m�X���-_V(P��؟z�RI��\����F_�P��*�"O\S�(�E�������3���T%@4V�"�tȊ�v>�0-�JUTC՘�D�!HQ���=
�)[�Lk<��V&��iy��d�p�BWLܚT�ar�2*E�t ��v�֍q��$b[����t�r'L=v~�ɸ�o >/�~9�*�?j:x��I>.�v-��ʄ�;`.T1W�_�/�"�HF悚6��]���"��Bgc"�I3k�u�tS�k��OMv1�fM\B���ӓ`$��@����@�5��9���o��Et�;?
B�ӰWj݂��
�%@�QDe���m����ذ;Ѩ�;-$������%U�ժ�Һ�n����ڙi�DqU��-K�Ҡ#��āX,H�󮎆>��%pHɠ?n�A��N
+z���RX�r�JՅl�&��p�� ���a��b�P]��	�dTyrn�@�j��Uo�6��'��r'�)@󩉱6�$`2�K8����I�3�8X��ʎ=�!Y�<���	�ϒvr`I��T�r),��S�S� M0Qg���oZH���ɞ�&P���bH�_�L��䙽"i�'�\ӤY�&`�e���#����!5LJ��3�6� d�Eʞ,&�rw�S�4$������Gx���'<���PMîc�0��*�1�$�c�;�"�Z�A�=�5I�,�n9���H~3̂��y���7��*���m+��"��~r�iرO�42��H6��'mp A���p^�Uqm��ZQ�r��$�tSW�ߗb�����E�*�` BJ�tW��^yr$Sb����næf�>�#H����<�&�'d�0�c�IL$y� �#"����M5S��@�bؽD �PB	=N*�\;�O�=�'�T��BR?b����'^u'����i��%PUqD=*0�s�,�J�HP��|��L���U��jm��P���r�<aǪr�z�+�h�?|��(3��DF|�jw�F:��؋g	��0�Ax$D�j�S�3�Q�;qx������ IW���ʅ�y#�<�ȓiy�Y�'ʪw<,T[S�� � Q����Iv��B��C�1=��@R�i{�I�D�*ʓ����ñp!LM;�'?��,��	�������DR@�gg�6� Xrb�7Pc�U
Z�ʵ�pOM$�T���M�X8�,�I��eN���/�J����b m��aAƴ�T�E%�la�D/�
1�~m�G`�\T�i�O[(�P�ҜF��]k�n		#��k�'Z*�X��6\Zx6D�"N������I�P��I@���dEx5Ҥ��	l��	�-=�'4������k$`�A
�K��q2�h�)=�!�� P�dg_�E�0aJ 'pvl��j>@v�@4!
u�ZR�Ƿ
��t�ɖ#]2e�a�2��1�3y8j����n�����ː,�89ˑHH1Ѩ�yDF�-@��!�S3����Qm�wJٌl�J ��'ףv��Eyb�P
a�G*m�N�ח��*-�i����$���y5�J��yrG��n!^� �IؓJ8Pis����?��40krIG�#l�I7.\�4����Iv麦m�=�ZeA��K�?J
B䉆�J1Ť�n20r��$��C�ɍ(� Ԏ��p��$ۜ&@B�ɿP�(�  ��<<�đ�B�X�C��Y

)�����h0Y��*d̜�
 ��h��?�)�'�}j��`�+L!$W�\9P"Ov�
5F#Z]c����O@�a��.GNH#�I�e���n�B�<��*]6*���臏R�!����yX��Ey¡��X�*�G����cwd��y҇��~�t�j�Dڑ:t�BV��-���hO����ȶ�p���焍_��G"O�@�U�L;�
��R��Mȶ���"O�-J7��9V�u� F\�G�8���"O�(�$ 0��Gް���B4"Ot1��_ HX�M�F�\C��y����lc��?O��r�Q�I�����H��-���!eąeA[[:�d�?U�g@�8�r�@ՈDO~ԑ)�K-D��Xe�&O*$%�6�WB��KT)�<���[ ^G@ i%�0|�!��"`{�4�ō��QlT�#DVX�<i4,��~��mX��O��u#�@Y}�<Q�݅w�����	q��"E~�<����7`i!���Q� �z�&Gy�<1��ޡ=9.�ń�N�s���Q�<CT�n�~�+5'�0��|S��M�<)��U�W
uA�a%3  \)�f�s�<�W)��"R(�R��-X6I&�n�<1'"WPp!CGǒh� ���GMP�<A6�)"����e�"Mz&�0$��t�<Bh׾8�<yB���f'BH���m�<��)?J�h �Ʋ5>�"��Em�<q�����d�F�D�y\)֣o�<Q'n��4�@(΢Z�`��f"�e�<Q�k�!PM��@�,�bEN�g�<�b&�A���� �
hȱZ�LT�<��&D�.�@g
Ǉwd�`��S�<���ԧ~3����S)D렼�BaL�<�Q�F-1�t�ׯ*$G�����J�<��!Lh)*�c�L�DaK�Pw�B�ɛjF� S�o�7{*怋��QE4�B�I;>��� Bƺj��j�"��"�:B�I�[|�mwe
?H��mG5I��C�I�n�ԑ�I9h�����P�(C�	�}n�c�l�.�mq�-�omC��. �ڨ�h��s
�,30�A<C�I3�^���#@�bv`$��� ��B��Pkr�ʕǌ��U8p�P�!�C�>��c�A�%�������C�	�1��`�^*:s\�7�
�\L~C�ɛ-r����O`�)!�@$�C�	}-z���I۰@e�-c�i��S'zC��C@T�@�"�s��	��AȪH4��$&?�Ty@	كB�Fl�ք���!��\�V�sR�ݎ�H,E�ƛ&�!��B���5��$��+} �a�5D�dH��V6�����.�`C2D�8��зW�8aP��Q�>u��-D����]�4Lx�ِo��}A�*D�� �@�b�T��r�`��!~����b"O,h�d�\�_������dh���7"O�M*&/^�ZߤL�v䋸Fl�}��"O9�kA'Yb�ґ�ن�B��S"OL�P�b��=���ȇCDX�x�cB"O����OF�Y)�����{�"O\,1w��H~���U�:}�x�@"OF�)ED+4LX+�U�c��2"O|ل.�CW<��$#\j��"O�q0��{P�&㊐@"��5"O��P)���(x��W�"b�4{Q"O�[�O4h8Yq0�Ɍ@o<���"O6���iR*�a�Vᝃ]x\�$"O���b�;>��9�&L6M<��7"On���	W�p��DW:H��!�"O,��$��6����F+z���"O����s!����[�|�"��'"O������%�V����P,\���"OZ���5�а��k8
F�4+A"O^�	Qm���B�_?,5���p"O��j���+�V�1
��%�y��"OV��h��+����	��Ux�"O�dɧņ��q(9����"OҜk��]�'�@q!���!��U"O@�@j���i�m�3d�
4��"ObQ;�ʔ=���gl�## "��"OpD ���@ ���投�B,&G�!�X�u}bI�EDC��5  H\�kp!�d��E5P��er��2��7�PyƟ&�С�E�թD����y�ʛ6X��=���M�i8 L���Ə�y�_`-X�	���� �l��'����CR�h�H�� ̔#��:�':�q���,1{���ʉ!����
�'�0D�H����٨�g��5�0%0	�'�*�������I��\+3�2m��'�؄��KÿqUt���N!��ɰ�'b�,�o�z�`�/ �����'��b����3�ܤ�'�ļ�,���'�f�kD`��g���i͐�o�H�
�'�@`��FJ���jէ�
p:8u�	�'ۢ�S�Πg�>ʔ��_W��	�'��E81!�=(�0,�C�=d�X�'�u B~\Y��¼�l�+
�'&��01��{��a��0<��!	�'��ŕ)g[q��_�@�a��'NY�q+_�l�:��,(.]8���'�Z��e�z�X�"�з&1�ar�'Lp�p�Q�^���dO=nl}1�'����q�ں�N�2� 6	B�R�'pq�� ��P�V�Qi�J
()��'ϼ)�"$�UR�:���C|li�'h�ZQNϣ%Zz��h��V���ȓ9u��C���&���cK]�-A��ȓLs�B���ԍ{@
هwkvԅȓ-׸���H�c��m۱��n���ȓ3Dq)��`:�u3��$j�͆ȓ,�j��ӈٮ@jŭV���}�ȓ`��寖�{�Huڒ��?�ȅ�{2:,y��W&D��)���X����ȓM]i��V�(s�h4�\�7�
 �ȓ> �����-1���{��%�\��ȓn���3���z�d�El�>>�A��(�� ��7ްx#�K"��S�? 2y�^�EqI��H>Deh�E"O��A��=50�kRo"!�))�"O�����S�ΰ[�n�V9,��g"O���$D�Ik���Ϧ7��y"O�xAKT�oBZ-;1-��[����"O|��$�R�uP�쨵���(��"O�|rfE��c��PQA�O%X�"4Z�"Oz�S�� H���� ��|�L��"O���e�i!B�R �M�sr�}��"OL���˧DB]� �06qʕX"O(����1�6�6���Ju��"O�0K�� AD�Z���Odp�W"O�HI���%Z�
�j���T��"O��9s�g2}����Ol��Q"O.�B2H*pw�\k��ǢBR�:�"OF�n�q��KPIJ�ԃ6"O,�!LS�9��Ԋ��j5@5�u"O��B�9
I�抃�z�Zu�"O�@�ĶcQ�B�o�]6��""O�!��H#���Ã�SO��
�"ON�K7��3�$���4��"O�����[��I�E֡D�"��"O:Ԡ�B��hX��# �O�����"O"��UJP�	^@(���;5���"O�ɷc#/�蝳�bC%:F! b"O� Aa!-.�*�����.��u��"O�I��H�)R �Dq���B��%��"O��8v��)��yya�ɛ+`(��#"Ov<���*<6T�a!�H��B�"O��k�*B�'%2��!�2�~X�"O�M����d�}XBď/q��a�"O���B�T�v����U'�K��i"OHI �-ԅ
��[3�K�`�v���"O�t�_�|�"e�"b� �0�"Ox J��
����b��F(����"Oԕ��KG�G<�=I�hH:�,�Zf"O�-KE ֋xK��@�	ŦK��	�"O�$kc#yɊH�VgU�o{vu�"O�I��WoS� W�F�FH	*O,�
��;j�����Q �
 ��'X̘���_@Rr�	8�!i�'�f����(��D�A�Ϣ�f|p
�'klh;�$Qr�������� 1�'�$�3�O��zH�!��ʁq=���'}��YEO��77ڴ��j�*w^5��'f@#���%"j�H6h������',�s�ǅ=�3�Ǉ(A���'�h�Ӣ%�&�(kefK�d֤�b�'�H(i�FͲ_�( kd��d�pj�'��̱��G� \8@͈�l	�
�'P��e� 7lMe�	Z�
�'�\i@c��	�jT�w�4[Vdp�	�'�y�WoE�Fp����^Yz�'�������H{`p !�1|+0��'��ȱ��(�*Q�##�#r���'������ض)x��S ր~�"���'ή�������Ȩ�� ~b��2	�'�`L��L
�0�zwK�$*�x�'��E��ƞ�g�D�i\5�Z� �'"j��D#��$V�I�G�x����'P��+�h�P��$2�#��d��'a��8D�h�d�cek�"q�dh��'Hh��<t���t(_�v��x�'K蜱�AO����2���I,����� �E�FD۷!y�U��EZ_�Ll""O~X��$z��ҡO̍�0ă`"Ov1ɥ	ʏn�fUj��̛�|س�"O��J�NĐ��G�L?N �!	F"O�������J��'��B-�\h�"Ob��$� 8�� S��p̹��"OXP	�,G� 0��a�K%1tN5"O(x��F�5�"�aN	Lz��s�"O�)��IC%���8a�[�����"O(�;T�S�,���xlUys"Oz$1T��%I/�U��͘�E�2C"O�!`ʈT=p���Ũ3�H���"O`�a!�1i�rqB`Q�D�Ȝ��"Of���"2X�#afyۺ�p"O���!�D_zqD�Z0i����"Oڵ�G`  ����T����� �"O�hpCϵ}���q���4��da�*O��k�	N�ղ�	?{����'prI��M9*�Yx��@\(���'�h��A�8����N��JG0�i�'���� �[Z��a )0����'w�4�ƃ���Za��m̹�Q��'��<����uȖ%(�*����C�'�N��4�E5e���.I�}���"�'�dW�Z%>���1cB�i��{�'�:{`i��&�qȊ�[r:-�'��0FG�/s���6FT.I�T@�'�,��H��^�8Y�=�3�F��y2e�6}�Ƥ�.�\�R(33��y�D9C�~ᘕ囂L��]9�㛈�yN����CآI�'g���y"�
k��f&�(0�4)֏̫�y�l�N9������ $�|��Ь��y��}V:I�k�(펌��Dƾ�yҩ��!�t@+Ԁ֟@4�* /��y2�HV8�)��s�^8���ȴ�y�C�'1���MԺc���o]��yₑQu�={Ή�Pp� �h��y�o�&j}�չG�+U� �Z�ٜ�y��C�;��%0S �r�:����A��y���-Wqȭ��� �l��yR��D��y2+T��HH�PBӤ�ڍZ��נ�y"�L#cҙ!�FίZ�\T�`���y��	6��| C�B�^����7���yb ��[��#͑6V8��'����y�J�V��k&gP�>�B�ذ�@.�y����F��=[
��{<Dh�n��yR.��_8l��iK�ܠ�h��yr��>�+�!kv"�y�y2�v�q��XQNIy�g���y���9D"��\��X�uc'�yR��Y ��RGݳd��%H��yB��'�^��"gN>�E�,�y���bb��KM�8���?�yҋ���z���$-��	�yB��$i0��h�t�~<��N"�0?9��е�:u�bÛ5"����H71������o�'�|Y�����Zh�ɰo�4 �5��oɖ��5��0��	��>q[��OȔӧu�[�S-B���U�|]�P��`ݭO���3�TN�S�O���Ğ�0��S�&��.��l�����I���8E�On�U�G���s���0`n�qQ�@��������'9��ɣ�T=��LR`I�} �L�O𩑴�2�)���<��3
ӎ*q���S�N('����Q�tP�?E�ď�_� �FX =�&������=�u*!�)�g�? \<��el��(�m�	r��S��<@���É8U�|�A��Na6����7qO�Yc�'�)�鋼'�ΌRen�~t��jâH�6�����+���NΝ	���fb�L�5A�'%�~����O�>�2�ț�J9�<�����K�:ir�Y�s���������tL���F;e��qSi�H�܈�?�	6�R���P&$Eh�gH+X��KB�Õ,M�㟒�p��R�*c���W��JG:`��>��H��?�J>���ܠf[�	q	��(Z�0f�"-i�d�K	�㟢}*E�O6Q��e�3�^K'��`@�D�R%�`��O(\��g��n]�B��2��-��$s&`xk�͖u��oL���
_�2��A�p`�<O�F1XwW���'�������H
2@t��GN�{�&��G)�;���N��I�?����\0hR�ԣ`(E�L;�@ـ�CO?�2�^�������$@C�P�)2-����d�_@`X dN�y�p%�O� ���S�~�l���ڇ�	,)��"l�)�~�ζ>Y��xZw��0�51�D�k���U+
2�X����:d:!�_We&!i�ɬ+Q�:ç]�V�!�d�4w���F*�d�t�E��S�!���S��A�6��.D�&
Ȯ;�!�$��l��J֏�z�q�Ҩ��!�D��m�X	�`NY��C'�K.M�!�ѦM��L17��!p�%!��ʊU��T	%&E�0���)7�-h�!��X0A�ݸ�'2���C����!�d�9,o���iQ#s#�	�)j�!��T;;��	 �ͱ�H58��5�!�=S|&�r�M"��,R���-�!򄙓�e��(}���1nݡ�!�䄸ҐȺ�G��*T��NV�{�!�D��t�څ'���uod���n�l�!򄚒ByH��ʎ�uF���%Ծ �!�$ׂm����98��G�q�!�ϟU0ag&��w���֪� 1�!���^�U9�����f��'�!�D��=�KI�5�PC��ƽ!�!�K=4��0���er(!U`.k�!�	=-�hɲq�J�DW��pS�D�1z!��IպDh��ٜC��J��7t!�D1,/0H'
ߗl7�m��Ӷ2^!�$U�i.�b�M�E8
���ʂ�c'!��MlI���ŅI!R4s�'�o6!����H}���P�� ��F.!���Ehle@U�Q�T�HȅC�+9!�](n��8��FH��,���:Z�!�DI�C&�r��(F�`L�$b�3�!�Ĕ
3*��!F���}�p哧��1�!�������?:�8�� �&�!�d�?;��l��ĵ8�~̹���!E�!򤙙M�B� �'X!���s�I�=}�!�d�����h����芷U�!�$G��X���(�btA4�L�g�!�d��6�
�R���&^�Ez%���!��Z9�8�Ts&E�5c�J!�dQ$t��8��	h48:%��Q=!�D_���%��^<�B��1!�D���a���Na���2�̎�!�$�!hx`�A�d�(�z��K�.�!�^�YZ:�#�h����ãt�!�D�']��y�k_Vcf����&G!�$?m��A� ,|LP 2�	�a!�dľ1b���FD2Ja�y���_!�D�#��ŀ��!}�0eC�c��(U!��U�^��e�̃���0��'O!�� R0@eN�+�j�{���0'~݉f"O�cC�Ȟ[�K3ʖ='�,�"OnusuB_(� ��JX #�-{#"O\�����I ����[�w���і"O��#2能(�^���/9)P(+�"O����j�qbR,W�%@T��"O��ӭaz�����V#R�[�"O���Jۧ&L�Ԙ���	/(�YB"O��鱩	#Pc��#���"�9�"Oj�ʇH��$g�yH�i���~\�1"O�1�ҽ���iBy H�3"O�5@�nK-�% ##:T�6�	w"O�A��`)&�Ӣ��.[ళ�"OT����1ng�����I����"O�U���jt�'*�~,Ji#
�'��Xt��5s��{��
��
\!�'`"��T���:(�؊�ƾq��p�'hr�K�ҵ)̝���[&{r6u��A��0q�`L�C8��r&�7a.DY�ȓK�H�fC�H4챕`մ5�E��ltRY��X S��a�V�	�H��@�ȓ|$���64�!&��q����ȓ"!�}*3�� ���g
F�̍�ȓd/����eP�8p�ԠT�ȱ��7�8, wk�#(�fē�\����3�X*�'��k�B|p�*ߗG�xY��@6>���O���{��X�h�m��aR���hQk,����6 j���~��� �T��
�X��+����ȓ[�Nţ�J45̉�F��-y���ȓd�&��#�9}����ѫG&�ԇȓyv	�!� E�n�z1EP'S�f���7��8�B�`Y(a�>2?"��mm2�����QY��C�J/:͇ȓ7��B1A�>�<ĸQ��7t�����O�ȍ�C!��-�T��K8]�A�� �2����_9< � ��+f�Y�ȓ)D��I�E�-�`���U�<K�t�ȓ@ �S$EH&p�b���r�]��g{le�Dϐ�A�ĭ"�E<����ȓJ��b�ȇ$:}��k���:��ȓw��}:P�P�~��l�'�Q�0���6������]�I��H�dJL9N�Z��ȓ/�8��`/H�X�������ȇȓ}#�}{A̅�I^���$�5Y�0�ȓmq:�gH=`�J�Xa��1����ɥ�ܲs��I���3|R�(�h0D������ʀ ; jՉ����Vg!D��ɢ
������ꔚ-��m��3D��Ss��,c9>�1qeR���T`7D��@�ٚd�B0�gI<pbd�2wl!D��.�'e��З��TN�h�a D��rc"N�N��%���v$!w�9D�$X"����R�D�@�2D�(*pF�$u���@���
\��-S�i/D���+�%���Ů�
7�إ��,D�։�"/�`U�w ��c��ѪR-+D���0��WBt�V!��d@ƁIv�*D��;5�*���S �k�zm(D��ó����QCB�T�+lp1I"�$D���_�Ndc!�βgt��� �&D��[R�O�9EnM�P��N�kUK$D���V����(�`�J���&c D�� E�גi�02uK�8DXp�#=D�� �0`G6b����cf�x�l#�"Oh����;^���f�l�F@sp"O�D+f.��d�U �׾-�t`q�"O�i�p Y�lX`����	 ��"O\{V�_��w��	wȞ�ST"O���A�7l�d�;%BI���2"O�بt�7X��a��B�;}�l\��"OD$X`̘v�($��(�$I���v"O�$�M�C������o�rX�3"O4�8�h([G��+c!I+b�H	cR"O������z��a�O�	/t<r�"O�E�W��T��z'%3=a���3"O���@��-e��Á�ңE̐�S"O2�C�"�����z�K)p9Z��
O>7�A>|g,�SBS�"�2Q#ڥf!�I�1y�AWD�*A���b��5�!�$J�r�m
��͹P������ڈ<b!�Dӹs�$��#�$(�I�u��?`!�D\t����勃8Q�	�d�?W!�E&*֘Q��g��Y� �H�Mv�!��Ѕ)�� ��C�_Yn\�talx!���b ��3"Y!D R�9�!��.>-r����l~���O�!�H�k	@љ�� =:� �Oۤ&!�$��N�d��g��N�nhȁ���!���(��P��H�8-�R�d
��'k�|IeĮF��x@R��#J�
�'#��� ѣ4m@\���B8RC����'B8�9ƠK�*Y��� K���1�'SތXR䈷8�ؠ8��A{���
�'m���Όd<����=9���'�b)���<<��1 eM�bꙋ�'��a�r���Bi�HH��z|��'���į`�v�5J�4�Ji��'KFa����'�XPC�8�03�'�B40�K��]y�$���n�e��'�����U�:���D�Id�dA�'�f�T��]
�D�$B50�b��	�'�QY�� 1.,Y���x�|�
�'Snřă�2Xh�"�I�����'�L��rM�w(�y��~t����'�N��V���)3���n�Dљ�'C�-(aW25�8h&�ܨ|Y�u��''�)!Pi
#�����"��G��aP
�'/��	CĞ-nf
@Z�O�4jhz
�'�{���"���%枞_򲰠�'ٸ]bv��z��Y�-��P�}S�'@8��x�p�"�
�<�H���'/d��N��<MR��[�H\�'�����O�%֐p���%-6�H	�'��ajū�?7������@
>�l 	�'Ԍ�3���vP,�	� F�!L���'�Ĥi�"#wJD��%9 �x�'�5�b�<#+���#'đ|�f���'|�`q��Oe���A�
ͩ�'�zYP�D�4*��bA��~� {�'��Z�Kמ9=��H�u�d �'�5�F(��mT�,XeB��<т�'�Q���07��zD��z��8!�'עpI�ϗ�6̽P��̒"O���.�>�����4�����"O��j%G�s��e ��O�\}�"O��1E���E�ؠ2CH�\DέE"O����F/h�"$�/
j@D��"O� �3�Δ
�6|�îIM"�ј�"O�,rb�� ���۔�bd��)�"OzT��D.����L�ZOv���"O�0�b�H�H|���>=da�R"O��Yt�_���+�[��.��"O�p�6E�D���c�^�x��"Of�jW��Ḧe�F`J�+"O����L_��궁�$#��p�"OP�3�n]�=�h���|�W"O�l�6�-@+��r#��5u��$r�"O�Pہ`E�b����h��Q "O��b*��&�0UA4Rt䨽�"O��ãܢz�*�0������"O���k�<861�&�'W� ���"O�p갈Z�� �J�T�.mp'"O>�"eU#LA�};�i���A#w"O�Q�p��'v�<����*Er 4�S"O�Y;��#tHd����'}p��r�"O���+��Q��-�YS�"O�-�PA� s@�#�e�9i�j�"O� 񖱴X�3�ʋ91H�3��
	�y�(X0i p  ���ɓ�!D�d�i���0	Ae��.Ͼ� �>D�|��O�,&Qp���5����e� D�q�Ł�e����E�A����?D��p�e�+-D�PL��F��#i<D�HP��J�%C�ꐁHX��q�(D� �EN��T0���5� �c��%D���ԅ	= }�
� \�Hp'4D���2@T�P�t�q"�:���qD!!D���u���lU�P�Zo���aF�+D�� ��V�X���S��Y��&D��k�K�� ��yѠ ZF;j9��%D�4y��!x���a��K̀0G5D�(
���--�@�0�D�2F

4;�(2D��8 Z+������JH����2D� !��g�.]p��L&p 듪3D�Љ#(۹}�fUJFJF�U?�h�&*D�a��D�%|� IѦO�XE��!+D�T�TB@l�IiFI�,9�a(D��3��	,���&�L�h+�ܒ��'D��R�ԕ +J2C����ӆ:nB䉆N/�=��a/:��8��
,)?C�4��!s�4��l���]8B�ɑl��C�ڍ2g�a
�kW�)B�	���/B#�I��R	*Q��$������E�A��LK��ߺx�!�d�C�l���4mr�D�ҧ�,�!���P��/�/]kX)�F&�!�dץ@..l��$'O�81Pd��w!��"-���2be�����$�!�d�&06L��t�ԗ$����DƯ&�!�:n�P�"�.vtdR"%N.�!�$������g�zi�Q
3���!�D%'�f:�TYCl��
)w!�$� �6PH0��]��P���.sP!�L�R�y�0Oբx���k��3F!�Ė{]ı��(V;A�̔``\�^�!�<n����]�@�&�{�@��C�!��Y-Lĭ!5
\C:"ez&e�5s!�$�>$�B�ӛ}֌Y�$9!�TD�=�C@ȞE�hQBە6�!�� �\� e�3j�����͍�7'��D"O���%Q��0���n4q1"OP0���� ̈�R��="�$yRa"O��IC��*х 1	��B�"O~�Pu_�K���q-��8�"O��֧E�`�|�9uL�r�B�"O��x��M���$&�5I�1��'Sv4j�['w���&� ?�td �'��`��s%���M<a%�
�
���<�~������G办�� �AL}��P�*V���7W�\H�"1��G�|1D�o��"�Bu��7��	y ��TD\��®T�x�që�g "]�觨�ܵ�&&�-%�z����yd�q�A��lc��Z�G�����(����'p8DX��&�g�t��S��� �c�%In �s�'�.�'nKp>�3f,�0:��elV�^�MK�c�`��_�d�hu�E�1ж���G�c{Lp�pǒn�
��b�mM|`�I�v.M�v��?!�����O��q��-_ 0	�V� U�E��a�7����'|����蟢����ǥ*w�h��+5�M)��8�D�8Z�D
��0|Z1�ǯ*2�x��!(1q��x?Y���?�S��X�������0�}����>#M���u*�d���cK�G�S�O��|A#�P�dQ.xҶ�@� �at�+�I�1���+�'%cf䂗�Ρc���z�N�yn�["F�x��2���+�x���)�i�)��� 1� �D���5Չ'&%" �韉'�9`���Ci�!K'�C3EZ���'��	�,��9Bg�"mר͹�'�4��#����X?^��9�'�~(���S5(}��)���Ia�8S�'���3ǟg��!B�u��D	�'%D��'̽Q�-r0�M6hYą(�'�ȭQ��E�[���I�j�&*p�#�'>�8��K�(F��y�����~3d�
�'L�"���s�R 9G�p�h 
�'�}sNZ'�0��/JZɀ|
�''Ɖ`��/FݴĠu��K�>p�'$�#�˛W[PH��?�q;�'�8�" ��.v��!j��̏6H>���'{v��J�?
M�Ȱgc�`K֝�
�'؄�ӆ�p^0L{G-]&c�>
�'��k��N0(��(��*M�P��	�'��f*F��D��7=�85�	�'<P��\��(d���;���'�6���l��=� bF6L��'*Ф�\�6Բ$)�A �-X�1�	�'N4Q���XQ�����lSꤥ	�'������#sڵ��"ʙM�4�'��х��9y6!��J�7@��P�
�'�&�� !-n���u�X7>�d̢
�'T�L؄M�}\<�7䔕/%�T8
�'�n�{��@�:P%sV�%(Q�	�'��� cZ���������'����У	�)��@ϙ�~���Z�'~�\2��1f��`��R *�Z�
�'>H�0ɀ3
l��kD�/v��Tr
�'�8�3�mN���"�%�$�<"�'�މseU�u2�	!e`3�n��
�'p���4�4{Jv�����CU���
�'!
i�G-��V@ƀ�T7>2`� �'�����@&w<0[I�~�$X��'ߖ�sh�c"����§u�JA��'�~�S�MF ����y�h��'��0�0�]z���e�ϰ0�I�'�4b���]i:Y��L��%#^d��'�ԑ!�� ��ـd�IQ�(�'������+���c#7(�5 �'@��!�I.W�2���H�Z�'�H��3��.��2@�Cj��P��� ��1��Y�Bƒ��W��<&QHf"O�5cP�V4l��U�%k�)���:�"OjeI e�GH1i���{Y���"O
�i��9t��	EO�(X��BB"OV�i�bJ�?�
x�!A�e��,�Q"OL�Į���(`%�)b�P�3S"O��s���8�A�wd
(E�H��"Op���BT�H��05c*����V"O�샵��Fw� 2!��6mLt�R"O�|⢍�iż��'�[e��0�"O`<����z�r�E��^K�D)0"O����F���)v�)���R�"O �ˤ�R+!�p3�6�2$ʔ"O$�˃O�,�Sf�Sؚp�!"O���S"y"�Ax�ˌ`�&�ZW"O�p@�$�*�~�j��ǝr`�A "O4!���6z-e���J�#o|Y��"O�S�Gd}n��G��6[_
���"OF剔A?4�� \�_*��H"O�d���1�d`���)[
J��"OD	�
͉EVV��ÏH
f	��w"O��FN�N�H�٠ON74e&��T"O`�SiW�F����� *XU��"O��i���
3��Ѡ��OK>�c'"OmZk$�����T�-к�"O8������g����E�6Z%����"O��ҡ�^;!�T�uY�:�a�"O���'d�? hk%�s��8:`"Ot��U��6g �c�D��^>�"O�!�ѡ!tN���1��"z2�js"O�T��U6�楚�*̮D{�m��"O������_,�@)La���"O��
��
$-��I7 VJ�@�"Oh����Eh4ʧ�W�T��""O���k�&M��ȩs(�N4@�H2"O05hD�]:2{�Tq%��x�d��"O*�����H��,�n��S(��� "O�@c��W�=1�i�' �~���2"O��8v��(Xnh$ a�#z��"O����_>dVn s!N�ga8�x�"Ov�j٦P'��c$O�=@Fxz�"O�U��EX�"b^!R@L%&S���"O��C�R���a�B��&\��"Of@�T��9@�dIJ��f���"O�e�pB���P=`t�x�:�"O0�Yrd���`	Ҭ�#t�h�A"O*�I��ʷc�� r��<,�bL
f"O��D)��M_�8�Q�J�Dh�L&"Orܻ�g�Dj!v�Q�ytЍ��"O�)pE
�:���h�bE�]Y�M�"O���9{?0�� ,J�"!"O���e���h�p���+
_���H "O�`Q�O	>�EI�S~�ɸR"O� �#��lYʉ�hH�N�J�"O�\�­K�>it졆-�z!�A��"O0���^�L��]�L�1��#�"O0<�Uϒ�l�]�� �t�@ؠ�"Or�٦�Sm� b/C�n�����"O�d��	��"fl�HE�8����'�!�䄒'X�qG�����K�j�11!���[�,HK� <�,�P�j�"P7!�d��
��	y�$��Z����
�^ !�$Ҟ+�B`�1g��g�t���-[	!�$�&] �!���\�� -�';!�� Ri��Ь�����/ئ8$T���"Oz����٠ P4Y��X�CJ}bt"OT"cɘh>�;�f�)3-�4z�"O�(P&:&��cOC�C��[U"O\��R˄!6M����7&����"O�h����^��݋f�.���"O8bU�M	��b�c�]�0���"O���w�ٗ'ō����}}]x�"OD��&�D��%�6M*2���D"O���@_�n���E�
L����"O�L'��4_�.4��D�F:��"OR�㇅I1��Y�R�YB.�0��"Oz��0#��O��)�sBW3.��"O�� ��D��A�!#F�qޅ3"OJa���ЭM���	FbӖh�⨣D"O��aǤ������֢F��'"ODa�b�"*t�� ��W�(�"Of�s��ϸ]�ԁ��>-��)�"O��J�J�!I�t��)�
#J!��"O��9RH�))\N�~�%��"O|ႆ�#~�zUm�p�l�q�"O�t�f`L�sPd���l@�L���"O ����i̴��#��*�TI�@"O0%�����"i���ek��7jtIz�"O��x`��8��E{*ĔxA�UA""O��tbM�6���؛<���"O:`��D�H4 ��l!N��"O�1�E�LY����o�;�b=�D"OBQ0�E^%7�|(���{���j���y�J�`Pdh�&M� %�%D!Y��yBJ�qdXi�B��qFo҉�y2��LS��(ӥ��+,�L���y��קh���5��8/���5-Z��yA]l�Z����~fTE埲�y�	 -&�S�眉�"������yr�׭Y4�d#���#����y�]�";��Sem�x�8)�X�y� 	v�!:�o��+b���v�+�y2ƹ@2H��gc�u��0	�X��y��8hT�$�D}�Lu�k���y�*H�<�d���)D7���@�#�yҏ�2Q��D�"k¾F߆�x`�L��y�V<�� ��%Aa�%P���y2�:X��sp��,���b���'�y"�!4`����"ʺx9R�y�H�L��z�� �o���B+V��yB��7�p��a��"k���j�I�y®��"����GF6i��pB����y"!��,�Vm8�K��0fЋSL
�yR.��6l�Qx�`�/#�
(3)Y��yb�4\)�����6��®��yRǆ c$�`R��Y D�|Z�d0�'?6�A�y��Y�LL.H�(k�'ҩ��G����I�	Z!��K�'�&�d�F�P�l�k'�=#�T��'V�@UC�!K.x	dƌ��%�	�'B���v
5$�1$����	�'
,���Ŋ^7�Y��g�9p8�� �'/%���J�@ Z���ZO:x��'-x�I1K\�;��vKW�R� �'�,�I�ǲVıK5OƢ&��L)�'WR0C��2Tz�̀$gm'�0�'/(��t*�+�&z3��*`K�q
�'�΁�#�)3�v��rJ����h
��� 谬�R��M�F� N���"O.ѓ��E&W�t�R(��^N�]aq"O�É�u���+���Vڪi��"O�}ȣ}pr0cQ'zc�e��"O��{B$�41h&�q'C77W4�@�"O��cƀѝ1���h
~ݼ��%"O�P�t��H<�ahͧB�za�c"OD�0��ަ�ܸ�@�ͯ\v�Y!"O�P(����d�:5(o��b�"O������)=~09�����!"OVQh��֢?�%�Kr�K�"O4�A���1m�Đ�#ćc!�K "O���ЄK�C��0�� �K���"O�E��^!Ģ�� �L�ț�"O��r#��3w��t������Hsd"Od��jпN�(��,�3�2C"OFl!��E	?��p�'�1/r� �"O��f��/I ����pP"% �"O�P$���P>h\ɴ�T)#BV-b�"O܍8�$�����=;�B�"O�!+�������@A��:��,S�"O��6F��l��т�ηN���5"O����G�;�NH�����	��"O�)Jp%D	�&a95P?���"�"O.e��I�/Eh9�B&S�]����"O����f�4H���"����"O�A������}b���+����"Or��G�Ѵ[��<rV�|xެ0�"O$-qV�Ѱ[�Π�+�a",H "O�8���Ǐd�$�Q�رt[d�a"OvH#��O��jճ7��<��,��"Of��!�Ml��j�n�~�0\��"O=q�'up��3
���k"O�PC/  0�ĸmZ�n�=Za"O	:�ώ�JC�lB7 %C3"O^p�I�jP�E����K��F"O6�2��  �/znؑ"O�� �Q���BD%RvH�a"OH�+6O1��8hS�hXf�{s"O�&� � �
�wc�
d"O�dY��Q
j+x�����!kAV�� "O�=U��@��=�`��;�2��P"O�0��M�;��
�NT�����R"O�|��Q�W��Y8�+&ڀt��"O�Ҕ���#�8�S�,J �E"Oڈ�-�+	̪x�6�TN� � "O������&n��v�ԧ}����6"O�������.Y�D[5+�'�~�Qr"O�19%���5ҮT�� ;���X"O8Y�Wa؆U9H�G$J��Hµ"O��q���T��`� (��� �"O�xw�6^Kҵi$��4~6H��"O)�T���f�U�`L�Rj �� "O�#��>^�f�����4)EF�;"O.M��H�*�>�uJR�F�D�ː"Oƥ�+;H��1��@",\p�"OԵ�COܿnk��5��O �|�W"OX��`I���mӧ��z	#"O.�x�Iɾ?��	�Ř)�r%�"Ot��נ6'�4���6�>��V"O<!s��Nvx��b쏫p��"O�qg$R�(��i���=P�\&"OB���N��v0�eKG�?�8��"O��Kwj.�D�J�`�@!�"Or�3��T�T��*��6B���"O��C�c\���a:���b�"O�|b�BFdf�����W�B�"O�-B���9�
��@��TˈP3'"O����*�����¨~����"Oh��a�X�0l����ʈ��\J�"O��,Ωq�ک�����_=�$�"OJ�+�&?WPBG�H�\#����"OVas��Q�(�x��{���c"O��¡�Mp倅i��;Q�( 6"Ol�"�HY�m"��.��d���:7"O ��Ǫ��Υ@F�t���Ǣ'�y��"u�5@n�>e���7�S�y����{⮹+�g@��c6����y�C��-�M�7Kׅ �h��%B��y��X�BuP�b��ߋS�E� ����y�hP�b��m[qiS?joHu��Ƴ�y"�Z�)a"9�'@�P�Z����
!�p>a�C�
+��@��o��	��Ñ�>6 b1�aCX�J�zB�	.B?�I��U�,�^��s"�Cc�`qC� ^�vT�nAk�O6]c���=uN(9��KqJ	j�'���B�E�L��L�5xE*'l�1z+hda���%I�����4�"R"MZ��:}"�T>.�lCa)Y8a
#�۲�yb�,{�X�X��c�b0y��#1�8̪gO�&�Bq(�J��7�r4�O�����%k���O츩Q�̙*:�Be굀�'J� Rӓh�:�j����!c*G���Ȼ�]�g$,AV%�'�`*�I�JA�Q�PB�eQ(a�ρ���3�v���QlBr�0!c*Jp>�%�� �E�Ix*�9�A�Ϧ�	@�˺K���p�A��g�l���C�K6���@X�9PH��� s9�̠��'�$`Z�%@�F*�����r�uZ7näcQ dB��	�D�!g�Ѧt�(xj��@B#�� �ŝp�qrg�w���Y��j�m���!guҁ9�'sѓ�T�@����җL=d���o�>KN��w@�JO&e����:�`	����:z Z��T�I4j���V�?OB� )Ҁ�^YND���fڪ�2��@�'�����m��PfY�5a٢@B4�3Ę4��+��IP��k��?�^�)���w��0IE�Q>`MF�C�ę6��1c7���L�i�ѣ�<T!��HS�L��'�Dt����TP�c��h2l���W?��j A��˶F��x���|�� !Z�q-�P���	B�pA�'\O�`x�͑�O�nщ��S7z�,ijB�τa�Q�dKW^�&Y�w�R�&E�P&m�5I�p��UL4|�<Q�D�f�P �6��Y�"�ȶ�7S� 	"O�Azq\���Yr���Q)��1��ab�!�%����#����R��Q��+t�@���
	�"!@ D�Z�ܕF�M� �t�#,Op�gLV� �$(a�		����GQ�D�p@OL��i�`�_�v�15�˧Ċ[�=�U���U��`ꠠ.��1+<�����@%� 9�J$+�"OHY"�ϕL_(i`���������!��lѴ%�dYD���3kn���+	I$�)�7��v�v �F W�Y� ��bR�������B�x(W��S�p�:P�|�Gt�T@�,�8T�n�rЮ��~��Q�J�y"�*�0����A�B�&l��m�-M$d��-�<�B��	���p���+s>b0�C�g Jh!o�rǔ��rgS <�k�4/�]��0VX�Xrt Ap��X �7��H���$ш�	C?f͒�Q�'�n���ޱ`�ʜ���f/���!�0:>�#^�X�H��ش9�>,���s���#�ҪR@ �CO�!f!j@���?��I:zFs�?.T���o�5o�b�����k��۷��"2ŋ����f�`�v�O ���ЭJ���ƍ/jENq�FI@mD��4��la���&$6l�ax�f�0z�(��W�Y�<�&��K-6mD$��n�+{�a���W�>�*S��s}2L��T�\�nZ�3f@,��l�Jjl�'��/:��H���-|Ț���'$ư�4���Q���S@�?g��:��M)Lp���p<��'�4%�e�T�9�$�3~�Б����S��͑��S4���kϘ������5�VԮ>���Qu��P�DL�T���f`��a!�
�O���CO�=���m_j@ʴ씫m-�LB$��6S��<��
�Mm��e�9T@5��k�sܓ*���ѵ�X�S�b\�Ј.(^���
HY��e(ݴY�����F*FF\�q�싍@�R�)��Gt��$ğƤ�@��U1��O(��e ��U[6%�Q�8zt
�0-W�eyb�6b\�=AU`O!C�6)���֦���4gKX�H��A��l��S�j�z��G���%@w�O�Sè1�'��u�Af�pB#	�rMZ�(�(�5F��@���'2��;�$ŉQ��I{a�g�T���>u@L�`�;@y.L�c���Y�Bݰ1DK?9�D�s�G�����ŽPv0p���Җ00�xa�� v�Dx��V�$uI���$-�IB�@)��	��37�P9"b�%}�h �R�����/������E�}\�9+0L2��6e�mZ�mB�9SbY9C�ƊA��D;�@٦t�.���˷N��\X�6  x;��_�-E�L�Ԫb:DӀC5'_�%ʊ�ě�F��`R��d��$��˥me�-RT@ڈ#lF�lǲD�6&["E
��X"@��M#���L��T+d�@�R��=*�
`zT���	���c��|v޽\vm�e�3&�9! �c���ەAW�X9^��a��Hx�N_?ZhQ��C��
4�yQ����Iه�F�^6�S��L<�JTe&�O@l:�	�#)4��{ C
7u�����+	a�eɹɾ@�G�:~G�J����UX�����6q����$*A����>�|�`BP�p�YF%��9�Q���3L1�p�P"��r �] fe�8�: A/}����uZ$�|��e�5-Ӕ�᧩�	ZβA	�/G0<Y�P�
Ǔ9^��$�&Z��Q�ߌL�BUoZY�,e��#3,���O��-`�������S����BV�y:���	
�ZuXM�(_`���'}���FƂ�w���ԇ�9y��{-O�mxf�&��u��/�i`���@����I9x���'XT,���ԺXH���`J�kB��ȓH
P�'��9h��3#�4���a�$ �}�������Y�Z�L^�r.�d��ƈ�
�.-��/D�|���������W��|�|����OX<H �W�4��I2Z�ёC�0��Г��%hB䉧���AK�M�zx��� �xC�h�V)S�k[��Z��F��(3����D�H��hI>�c-�&Pr,)���#`h���W�<�4HәD(h#��K8s���#B*Y�D�s�|i��4��I��B�n� ��&�Х�QN 4!�V��ѓ��K�^׌i����&V�fw��طsZE:���͛L�\��@հy�Ds o�&cN!���I����C�^�i�=��ђD���ؚ8�٢��4(��_�Y���Rl�"L�L���5'�4��ea�bx��1c!Y�M��apG� c{�!��/�8�`5��N��F��U)��''� h�	M��\ȥO>% ���[��j�'�N�VЫ�;D�ԢTd�3$� 	�']-aDMF̯IF�[9֤�tBMZ�g̓^� /	����.!4w����_ Yt*-xQ*�)�1vZ��'F�>�:��7�O2��
�=;�Q+�B �m�8tR&�'�r��g̀� F�'\rq�+��Q���@炚q������ <ĸw�ô">b��OU�'v>B�"O�`�J�Y��)�7"	��"On<����	��A)��"O �ϟ�?��yZs��X�P0"ONi)T�$Ŝ���
αZ�ihB"O����ܼC�n� �H�,D�S�"O��( )O�3F�5{�"ːo�*�R�"O����Dmqc�"�z�lPw"O�P #]���`�je����"O�4b��+�zL��T#[�U)s"O��a��53rDI$Ú�05����"OT��IO5�d�;"a�� �"O΀�EfO�Oy6�p���67�r�R�"Oj|8�C�^�2�+��5y�*D
4"OL�7.K�*��(je��#�j�[w"OXuZ��^�R����D���"O0X�HF| +�)�hPʇ"OFBD �0k�@0�!T���e��"OJY��h�z�|�s�O��>�ڴ�b"O�Hb��,ΑCw.�:����F"O��s��]�
-& BC���)>���"O֙˷cL�&0���%O����"O�K0)Q�ot4�GI��au"Ol�9K�"J������$?�@A�P"O�T+r���1��f	�S}"	�"O�(�0�%���[�gU�8j"8iu"O�Tz�/�tUP9��Z�c_NM:�"Ol���+W��#&�I1TQCE"O�t��	;
���:�Ɣ�g�B	ZD"O^��GjK�!��5S򪌷��!б"O4�)�DS+-}����iO��֜��"O�|��!^�{�B)S��ԆiUF9Yt"O��8e�W�1�:xCfE;Y8i�f"O��れ�8�@邆��&1�`P�"O(��H4V�����S�Z���r"O�t��ܢ
F��X� )"OFTTa@;~C̭sRȇ$.|L}�"O���`fؑ9B��h��R�j
��{�"O�4���ߋf���xºB����y��̟n�Z�c֠�?���Svc��y�d��f��t�ޯZ&T��E�y��<YN�p(�%RD���L2�y�Ξ�il�gȌ'Tzs`a�y��Kb����U<��@W�
�y��M�k�����*I�s��̕�y���..�j�h��4um֌	#�ֱ�y�蘂.q(�����dph�$�N?�y2��4#^x{��Swn�KC���y��BTu�5RƌI+<&� �'/  �yb� 5��|C���L�&$�&�\�y����Ue%3pM[A� $1��"�y¢O$ ��98We�*Ic����-��y��@�$����ϞI��PH`#�)�y*O$D��&��M�)� O��ybDN�@qRH�S	�]���n���yb$�qۆ�[$��4��%�FV�y#�&�P���L�W�٢�y⃂��x�n��xBW�A$�y��MŬ�I�I� xr ���hQ��y2I�����bi����i��yb*,и�f@e���Q�	Y��y2��/D�p0Idi,T�F��y�,�6t�(�Kۑk	��s�*�y���(.����@L5o�&hC���y
� @��a �*�6�sn�2.�`��"OH]X0�����0�.���\1K "O �!�<����1�� �"O���5mV�1κ1(�i�.#�P��`"O�P��
 w䀠#sn)]�Vm��"O$p�@c��,+B�SC�M|���"O~�<X���P#\<�B���"O�J�Α�o�Ph�Aa�.4`�lB�"O1�vj�6)PQK  [�Ih���g"O��;7���G���uoW�k�)�u"Ot��-BH�`���6Wb��""Oޘ��ı iQ��DD����"O�R"��f�Q��S?&;�8�"O&LҐ�ٟX�E�@(Ś~�.- "O�!+t�yh�MȢGȺV�X��#"O.�j b��Mu�Tڧ�߹J|����"Op�O�8�`|0�Kr�%"O�):`���
5�H��K�x+ԁ�Q"O�e0����� (�ҩ���"Or<�4�=����τ�p��Rt"O:Չe`*^z��b��J#(Ѐ�u"O���[��"5Z��D*M.6���"Oh峀NU�A���9�f��i��"O8���j8~p�t꒜L�$Q5"O\y�D �v�ź�hJ���`�"O�e�4��8kH���	�@��"O�=RA��$�V�䣋�~�j�� "On%"��t�>�P�%� ��"�"O���J�DP��1��!(^��2�"O��Ҷ�T(u�x�0�c�d4�l�q"O<�*�� ���RW$^^�IH�"O��ir#�h��a�Em'pM��"O�PZ6��3g��9�3�%^�j9�"O8�9F�ӽIz���'T0t����"O�h�AJX?f=J0ғ��7İ���"O�m���OC��ܓC��X�`]ۆ"O~U�E�0���p�ƷkR�3�"O�e��FƖH�D���MݱEG�6"O��5햏5�D��.��,#��0�"O xz�)Q7W=z� 6l�',�l�7"O\�ӈF+���IUkZ�
LtRf"O�����Іg0��hEI��X7"O���e�ӯ3�1�!.�O"�"O,��6�X&xF�0��K�O�L�	�"O�`��O+ؤ� �R+��h�"O��"�
�m��
��<}l��d"O0��#%�6��41��?.6TҀ"O��:V�%UÚEBb+��m@��u"O���WT��+R�dIZ��q"O&�r��
4MZ��K3<�(�"O�����>��
G�։:�١"O���իA/.��4*@�>,�TQ�"O@|�v+E���\�4Q�q"O�@�v�Z�V���B@��-�lP�"O���T�X�'���cDO� "<Ȗ�'܀8��`ێe�6Պ�H�g�[�l����h���G�<	v/�V����Oώ>3�y!CI�v�'f.E��ym|��<�'"���xVĝ1ބ���V�K݆�=�$���l���ZC���iM��C�?}���f팮����?���C[�0��TxM�h�@� � %~��ӎ�������0D�ĨG�0wt14[)|Fb�#��s��SbN,��m3��H,sE�p�'Z��&��Z��'4��1��d�*Ō|3E�ү:��Y��	�"�@�d�%a_�lʦU+�А�Ώ	\�$DH�L���T��O�)���е,BF�X���������D�M��"��j�,ě拊01�qO�A�5EhA�DB& ŒRx�\�]w�z]1f曓>��� ��J�F�z9l5���4���cL�(wh���C�#Z�a|bi�x�D!�JӦY�R�����X��A� 	��"I����J+>̙5�]{�dipj�$]�B��Z�'띵�,\���^^���&!��y҆A:1%�}��)<M@(ۦ��:n�d�4K����d�k��T��&�:0!�Q��ϿJM��+J8m�#�΀C���Z��˟�����p=�'��C7l��S$عWؑ;b��;�k\"�~x�S�� g���1[����`hƴ8(V=���:d��s@�d��=O�9�u �t5�,q���I�{Rb�$Ay�2��lE`1P��y"�uz�Ǐ P]�f�G�j����W�l�F\��i�f	f��V�Y�z_���FM$\O^<j@-S�9?����3WD9�š�$��#�j18�y󥄐ACH��<?2��6�Ü5Z\<i�$Ţ��fD�� �B� 3k�{�"O`���#P�.�{��FSPMyUǸ0�9Uj�~}���*=����*U�聱�)� .���� ���bR`Bq �F� ��7ެ��'�p��2�ژ�tB{֠M��KJ�q�]����~�`�'�Z��pq`��`\���W}ݲi�Q+��''���7n�"/�$��E�!�����}b
,-#��@��;��,�k]�|�����b�%���
�m��/_��SW`\����t��.g�8��˾p����(LO�}�	6X6����a�0u�c6��L�0�&���qF�R�y9�I{�εW(��f�*]��C]6��Y֢�j��}2S�P�P���:4����J�A�BIc���uJE� N���!L��!c��N�
���`��j���aɕ�b#�1���V��/�����M
�-�������U?��S�,\O�mS�f�=���[fN�/tlY�B�*����F�8C
��۴,�R���Öxz�� ⇉"pv8ԠB�D�5~i��'���I�@m�f�K;4���0�
�&�➐q�S�m�tz��B�R��!�FD�Rg(M��'�2��j͍�)5�.��j�0�(8�A��<�
��ӽ"�~��,�ʍ!���!vΡ	fgJ(����b͝�5���x�G]f{���B�޻+���=��8���e�B��{��:1�o�F��J$�E���+��?�nٵ"�lQ� ��5C�8���8�qk����	2M�>��3[R `�!��oP�p�ϸgў=�ӤE�S���1�Q��8Q��'�`�[�%$C�&�G��q@�	fr���Ūšq\���'L48���-S$����O B�&��6�°>WF�
%{y�EJ�(g��Y'N	� E ���	��'�$��3�ž*_$yQ�n�w�Z|�֩C�;�P�ҵi��qу�r$-�`�p!ݝD��h�� �l�p��2��id�I�A���4��	C=�,�K�R��ja�ɞI�d�X$㌑:���p%�-N����4��F$�!).TYh�4&LxL{����AUV�ӄ�(yMf|���$^��d"7�B��#�/;�(���Á_@$*���[>~��#	�8�e�ҡ0�T���c�+0��Ph[IG�V e;���A��B0@jQ��(:�{R��%l\��RC��b4��UᔏAxHD�oZ�W�Η�����*�!> ���-,UdPAQ�-	�l$��B�*x���rU���߳������aH��C� #�	5w�D��B=a<<���0Ā|�@�xU$�C�-�iX88����	m�^uQ�mN�a��P�VeB /DV��Vm����D���P�7b�\��TE8�xs��S	�
�C�&	7�Z)	4
5SN0�ؐ,�<4e�@3�,T�M�ʈ$�5�G&]~�=x���(�T@q`��>�<A�g�C��h	���t����y�F��+��rj���@ǁ�*o6<�Gm�8|��]a7F{ ̪���% �^����fz�A
�"	�t�Q�\�/�a|�ێy�\`�鄲>��y�ID�R�2�K��ފx��4c�� �TXuO�<�'�2r��Y�)��P�:�k�hދ��ę�B9(h�T�Ėt����E�2�Q��9o�A?$p�4B��v����eMI3���8��B�d�{�����l���BY0��B�g�&�GJN�� hp�T�p<q���eP���fB�q���P�զݺ����\�t.���T?M`sa�^fe� h
��T����*&��¤��"N�������xo\�l��@����6��12A�����2WP�l���8LD�+7���;�>O�9"aΓF&#���5����m_����Id�<�����l��))�0ؒhĘ\� AHP�	&)��I�H���8;$൳�蔙"E>-��M�R��C䉟"7�I��܄sR����2�����4O��E(�Qy��P��C��s��P���N�cZX���2D�<IBc�.{3�2�A
�*G�ړ,3D��X�C�'j=2��bI�2��d�Q�2,O~hh������jA��q�6]��KGY�N��6�U� 5��*���	r�4u�O  �%�	(��O�q9�3:��t��3b��0D"O*X�F��� �$�a�cD��ɮ~��hvJ)�3�I��%��ᝈ6zj��%�XNB��$�iK�&J�&�0i�~�xd�F�B5Ac��!Q�'dr\S�.� 9(���m�'�"
Ót��Q$��j��'��a:1 �Sn`�6���T	c�'I,q;�쀌i>����$V �X�1�Otxie��-ƭ�K�"|jՈ�)Vh��:񋝎>4�`�r&M�<Y��F$R(��JՄ-���3�؈`:h�'X&)a �3��Ϙ�� �����+hr����~�Z�qTO������I��l{��L�G�~e���r��ţdH���p?�U���9�>�zp�M�V���b�L8��ⴊA�6�\&�DB�+Y5^Pc�]$j�D�a'D���U�=X�i���aJM���$D�<�p�^�t�.'�2]s ',D��	��C�F�p�7*�w6�B%C+D�$:%N�5��xr��yc���=D���d�ʒj;Z�v��fµ�ƫ:D��q�(��&m���H�Pc�pVb6D�xh5n� N�I!$d��y�9�-)D��1r+F)`�4q�n� r���� !D�`j���>*��DJ�LE*��CƄ?D���K�f�p�B�D�(c�0��h1D����B�Ss�(7���5��[��,D��ɕCȬ�h��f�k.�h�c+<D������>�@X��Q� E�> 0!���!r���"ӭ^�*~\m�"�L! !�Ā�ab�����Q��\Q-�27!�D�(%�i �M�T���ɇ��q�!�$�
�Q�G�!%�ı�FX,&�!�dEi�t���@X�c��P�J�?^!�D�?̸}C��J�|g�%��$�G!��1@�|�ж�C�m�J���r�!�Ą�%W���w	�6bS���#ގN�!��_�r�H����� jؘ�u���Pr!��澱3E
�0V0�q/Z�nm!��:_�\ZE�΁�����@�Li!���HB��7�]��٠���"H!�D$i&�%��H(���)w̘`!򄟅l�4��`Υ�.8��L�=L,!�$�+f��У��d�T�0��;+
!�S��a`�m�R�Q���>�!�$#X�bi�cL��6��-�*m�!��3Ox�JB΀�0�΅��$���!�F�?�0�a��7-��q�J$B�!�ξ	�$�y��#g�����l8q	!�d��Gi@��q!�Q��J 
��oV!��Yc��5�H>�`�1����M!�$�=H�x8g�?4"ܐ�2�ۤq!�dQ�Q�B�Ҧ�7>�t;Gܻw�!�Xo�����(xdp{��w�!�dA�
����]	*Pε`�ÏY�!�D�@x a�K�<l�9��!
�:�az�f��1�|��e�d��9��m��[�<�"O�%C1��M'��'V��EyJ?-��C��+T��!DƿA��x� �<Y�*Ɛ�U�<�;����|�SBD�@A����ȆJۄ�1U�9$F���ʂh�'/a�����_��8�u�$`���J��(-���Y|�W�B	��
Z�@ؒ(����`T��v�����EJ�~b�D#
�>�3F��)�riYrLD#s7�`` cX�okn��\����&C���xSc+�~>M��������I<al�a�4gw�l��H�(�����ZV}���+�v��Uc,K��Y`A�]eu(���J��_4�ŦO�T��
'�2�QU��a;v��8w�Py���	4��q�6��'fJ���&�j���5|\��*J�Vӊ����ḭ������M��4"��h$>�O$Ԯ�/Kt��@^,f�2vϯ:�F��d���7��P����E�����9��U�KA�_16M1�O��a85R�+�0D6e�Cs��%,Gc�')�O���[��њ;�ܨ�@�E"���̎=E���3��
���Y4B���0|J�F��"u�űW˕�`L�I1�-�tiv�"BG�{�^��DؔC���~N?e�R䇠g	d���(hXS��+D|r�`ƉN�|���Ƶ���)D�8��M��n�X��B'�+P@��)�y��؉�iΪt3,�U��|b'=0��r[q�8�cF�ٟ�(A�w ��7�#�T>c�0x1��
b��� ʎ�D������)D����5��	��B� �(��r
,D�����"?�Р#ѻ�����+D�� ����)Ĳ<nn�§L0spl=��"O���A�>W���!��(9�px%"O���w��.[ m:��h�l�:�"O�{ �Vw6�;1��3X�*4R"O��j��1� �+���(Y�"O�x�C��>��\�� �E�v���"O�H'�Ck��=�#*�3$���H�"O���J]�\H����)�h��"O���'_j���gɓ>Ҵ��"OB�[�J�9D�0����=L@��"O�0���)k}>x(�#Zv�U"O�(���`l��r��<R��"O6��
��6�P0ۀ�Ul��"O����2$u"	ZB��XW�#�"Opm9 J��5�ʘ��^�K=�d��"O�\ჃQ.:0�А�.O6���!"O%;s � ��|�s%��2��Eȳ"O�:��[�l�tD��E�>�k"O��
#(�a�ڍ��%���if"O�U�r�:4 �I���3�b���"Ob�c -��8vX
�E�|_n�(�"O�푔$��E񔤒�D�z��@&"OԸ�`�"*H��WC�%�RE˦"O2��/G8nЉ��&J>�s"O�0����(��,��	,&��!"O\�QQ�O����JX�y�y�#"O�3���vT,M �ğQ�v���"O��r���8=��ɒu ��\��d"OH���%B�K������+(�a�"O(w
S���C���+%`	�d"Oft�#��~�&�D
݋k�V���"OV�t)لV�T	��rҪ#"O�����Է&�v�21f���("Or� Ƌ(Z٘��FD¨&��M�g"O�Pj ��C�"p�q� �"Ox-�ȮH�ܨr�"�6���"O�s"aٳUi��� Ō����"O� �IG�	������<�Q��"O����/Z�;[�̫��
	��m;d"OF��� Lb< ���� �e�q"O�i��Y�84��Ѥk|ӔQ�s"O�%���4s��buA��~o��"O�Ǌ�8��L�tc�g�0��"O��cpH�Tt�4�CI�m�0�b�"O�t{��Z�Y����8�Ⅎ�"O ����Z�4��Ʊ|��a�"O(��HܘDl��v� zݻ�"O��`B1o&����� J�)�"O���&��� ��m��B��4��"O*txQC��4ٙ�k��X7J��"O$���ϱ'�,��g�Z�)N�ѧ"ON�I��?I�h��T6zI��"O�$���+*�B@*���4�H��"O�	�D#�!_�JhzE�W�(�r"O�ĨC�ۨ�����s����"O�<	3��!=��(s�C�Z�ȈyF"Ob��C�%�h�Wh�0�( 5"O�����ωcs� ��U�Pu�$"O"�ɄJ@�-����''�0H��"OH�9w��1^�=)���68�����"O4�;��
TQ��BF���3��`"O-gk3xb��E� �ـ7V!��b������6<i|͠���^�!�$�'/��<���&3R>pB��2p!�� ���B���Pћ`#�/��q�2"O*h{�CR?%�0��1��8�G"Ot��m�rZ$i(��jܬ��Q"O�!�ѩ��/�� fQ7����"O�m��`�1@�t%	�Õ�7^x�"O���ݘ"�Xt ��7�XI�B"O`�h >$Μ S'�Zi�~q�"O���4cB���(��֭��H�1"O>Ls7�B1�X�w�ѹ4���a"O�T�EO��-D `�\F8%!�"O������q"ܙY�G	=}�t�c"O�H
�ϔT��Q3�%R1��"Oj��ǃ_/���*7%���Bt"OV�ĈFZ~,hنjSdߠ<xc"O�q���l�\3���"��i�"Of� �ڜϚU����&7��Ȅ"Ob�!�IR�f�C�@�[��%�p"O���1�H�;�800�X�#�*�z%"O,���ViK���lt@��"O�Pa���p��a��(
|$��"O�j�	���M	�aY,3�u	�"Or�CQ���PpS a,��j�"OX����'���� >gvX5r�"OUQak��b�z �$�����"O>���J؏P�J�S������"O��0�K���@�oFd}@��E"O$ɘ�d>+��,�AE��Esv��"O6�!wkn�Z��dLH�`"Oj�Q�I�JS�ݡF�+LR!��"O�(Dß�m��љ��2H.�(�G"OP����χ{���,P+4':�Y'"O2��a�.Fd�+ I�?�6���"O"	�n�+���4-ӧ%�q�"O��s1+�Z:� �}��HP�"Op)۠@B�XKr�X��ǝ,%��C�"O^��3dH�v@�E�Œ�x��Z�"O|�q�n��Jb�����ߤ1.ʑ)�"O�e�w�F�0�j�q�#~N9��"O�)�P�P�9�X�q�mN"#�*�HP"Ob�1���<�4�j�
ג�T�r4"O� �%`��	'n���r�"O܈j`E�)T(�\ʞ�.����"Oθ�BKÕ���ab��-e.l��"O �$�b!~ђsL��]��eB�"OT<A���j>��T�I�c��ق�"OJ��өT�30���i��Ȣ9��"O�9
��Ѣt<$�Z���-J���"O|e[�΋�iZ���`�t�V� S"O\���Ÿj�U���Q���(�"OB�ۢ�t�N�ip��*�ĩ�F"O�R�I�I�ʐ3��I邙�"O��B#bP�c��q�!̗y�&�[�"O$I	�n�gl%�v`F�@�b�ٰ"O�A���,���x�Κ3I��q�u"O�л�)�&QZD��x�jD��"O"��V��"�|�XӋN�(�R��"O������J3~��+�"5}X�i�"O���B+;,f �L�TU�a�$"O�9rp�����X �NB�D"O�p:�	�ox8���VM�$Q"Ox�0�
D�����īZ8����"Otk�CN�!I*s��>/�r�+�"O1r�E��%/��`�V ���y���mu��. �E��Z4�y
� 0�H�OW�4x����" M�dhQ�"O
�P&L>4���5�¥،0�b"O��K@�_�1���aF]+H�0P�T"OP�r��-+�,�p��ǬF���A�"O�,����$f��w ��k�8�A"O`��p䓡RBhU8���c���r"O$ �rL�[�.��o=�["O��q�'�V�>y8!a� m��	�S"O��1q�ٕP;�k�����AR"O�l��Ɔ�M���g�ǈL����"O�	g呔B�>���&�&��쪦"O��J��_=�^����2�(5��"O�����F�>Z���g�E=b�4�q"O�Xb�̄4�TcC�ߝrq��:5"O�}��,��[���Ã ��Ra��"O�q�$O
U80l:���+�1+r"Obd��l�%n�<	1"_�Xa��y�"O~��% ʺY�����AחM\V4�F"O&�Gh�J_��� B!t�thS"O�xp
�z�}z�ܧ>�v�`"O��P�lM�/xj�#�kV�{X$���"O��P�<F�D%K5«x@|YP�"O�تЬӔb(�6M�$T&��"Oݐ1E�&��T{PI�-Pm���"O�e�R	N�X�E{�f���-�ӏ)D���ك2���%_�:�
*D� ��-��-��Q���G$ ��&D��*�@}��t���=>��Z��9D���@��m�^��B&�+�I��%D����_�	�tL�(�tqa��$D�<��������&�%�=i�%5D���S�lؐ�Z��R@��cF�>D�DR�F/$"M	df��)n�B��;D�8���Ŏ8bb�SE�ھI�����8D�hJ��o��p;�Y�-�~H+�9D�r �8'�\mQ��Q�DbB$6D�����I)G���DҠGe& �L'D����&���DTB�fQ�t��[�%D���� �K0�cA��4m�N�<������-`\T��Y�B��	�ȓ.h��$��X� 1�V�K�Y4�5����90�aM>,�����,O5>� �ȓBn�$��:��	�`��&[��l��l	Z�z0!�3�@��0���S �/D��b�䆜Z��y2�C'�N��/D�4��`�=�x�@^�zz�y!�,D��1�*�<V�F���"G��LS�K+D�0�w��	E����@O�\d>A{d�'D���A�KbE*c�N�*��B`!D����H�|�% ��_��"Ak ;D�ċ��v�0�P���0�J�%D��7�:a��ӱ��8L�}��0D�D�a�� ?�F���BM�z�~�Q�)D����  ��0�NK�3�<��,D�i��l8 �*��LO8���+D�L���P .��Q�ӡF�"gh�ʖ�(D��1�����ع;V'�0�>!H�K&D�$3�ɞ!j2 ���؎ef��'d#D�,	AKY�uZ�A���X��XLҵg!D���eKR��1�ƌY�n�ٶ!#D��� 	ۼ@ tiy��*�Xp�U�,D��ijV�`�����Q7.��1��*D�< ����12�T��Z�?�`���=D��K�~L^L���~����<D�� �E��Nϥ1�,�S�ȁ��R���"O�,�*�~�t��5�L�s�nP�"O�%�v����� u��Le�"O��jr"���XqqjfJ��"O�l���{̨E��E�n���BU"O������e��-���@�"O�I���[�܈�ūSDg�t�p"O$A���Js�h�����RN� "e"O.U[ccV�,9H,:���98 ��"O�y*   ��   a  <  d#  .  �6  �A  (N  Z  %e   o  �y  ?�  ��  �  c�  �  ��  ��  ��  G�  ��  ��  a�  ��  
�  L�  ��  ��  �  ^ �  D � �$ + k1 �7 `> �D 9K �Q wY Ne �k 8s �}  � � J� �� :� ��  `� u�	����ZvIB�'lj\�0"Nz+��D��b�2TH���	#Ĵ��@��?Y���y�FJ%L+p���ؽo7��g���|~�tz"��)b�y�cFٵH�h*���A�N��WJD�i�A`��I�"H�YP�ԋ><�`�T��������]�mN1҇��7��쩀�	�0j���;P"�����?A���<	��)��K��p�"a�łS&��dJ��ν]���͹"��X��ėn�6mC�:����O���O���`j�%��V@~\:�J�8c����Ol���LU�ʓ�?���E��*��?9�DP�cV6�(Q+.y�U�����?����V�':B�'��L���ug��f�(�p"(@�Jm�r����c��{w�Yx��&�<�O�Ԁq	-ʓo���(T�	VdRd:��I
c�R0� �����ds���}b���x1Y�\{��J	}��Q���z� �!�&2l`Ӵ���O^���O��)�O<ʧ�y�B  ��)���ʍu4�Sdސ�?As�'B�6,lӔ�oZ˟� �4f���S�i���;B`�%����(�n��	�a����$��/�P|hj��E�I��d~��k�Ik�_�`F�|�G"�<e��(ڶip���b�H�~4�7^ݦ-R�4��4���G'�EV�����3Wv�P��=D����v�i���s�(<��m�^S�D��!8���sӐ�n�.�M#�c
�05P���3�(��năM=l�1e�߀9�8�&�i��7m�Ϧ�:&o��t�T��FY�v,��Îp&�d�`^�)D�(t#W�t��
�mJ�
����BO<�M���i��7���E��B�P�J�{��F�![R����l�tm�g�(��p#������e����,���"n�n������(�?ס֑S���֊�L���BYh1�ᜒ+��Q���?���|:��B��()B�?����rBȒ���}�|D�S.��<l���������O��D{>���IS>$ba�C�jUlڼC�*�U�)5��}I��U�O%����82֔y0V�O _���Rr�м^�E���2�QQi�,=  �L�(�d���	,�qON�"�'3f7-[Wy��
i���a�� �^��&$Ŏ�?���?�K>I���?Y��?�O|؉`��Z.?����Oƍ_/�@i��5g�VJ޼@$ ��Z3`�B<	_�7�O �oڞ_�V���4�?i*O��������I3���"���~�I�	J�����O<8���ݝsADX���D( ӖES��͸O�@	�L�<'����4��nW�� S���z�n	/�d�{�`ّ A���]���1���Ϋ$�M��)���
�JB=��k�$ Iv�j���ɰ�M�c��|R��[�j$f�
�(����Ԉ㪙@��d�<Á]�/�D��@ˈr`���N@�'�@7�ܦ��|���$;uʄ�ӦՀU��ڳ͍ӟ|��MybBʪ9���'72�'7�ɤ+$p�A�������I9ܰ۲�J:.��9�3˂�c�h� q��`�4�O�R�'�\s��#��ѷ	݊��i5ר" 1C��U��M�"�2���"u�����)��h�+�9�d��/�֙��LY���paaӢ��'�h����͟�'�V�2B-�lC���w���z�I��'�U����S�g���8XDl@��!o�(����JJ�I��M���iɧ�$�O��	���w��y�c@ƌ,H��D���k����'3��'�	}��0�F���_�Ճ�pp4�{�ς�)�6uP�(�*PX�B�?<O���"�H�Yf��4m��^h,dH�f�$�GO(B��)���r�7��$�l�v�Ą�I$���o�:M��Mz��_��H���'H�6�ZQ�'��O�hQ%D?'ĝ���S�<�����O^���O"����%��M�TnU="��\q䀼�'s�6��Цm�'���>��{��L���ɪH��T)�ፘp������?i�Lϔ�?a��?����0�*�`����TlDp�0��t�
�)_�D��l�3hG�e�Э�!0�m���CT�RH�8����8;��[�N2Vߜ�6&�p�����U�buk�4Y �K>iek������4Wӛ��'����PB7&m8�u�Z��[�\�\� �KyB]���	G�'y��q�h˄C��9�����^��+����3�C�ퟌ�'����$����n��cBA�((�:`p �0�?.OT���ʦ!�����I�?�1����@��/�)s�8�3"�z����A ޟ�ɷJ����Tyt������M�.� �'c:�ಓ��a�~��$L�I���Ou�Ԫ~�l�B�	nv�izb�ضy�b	{w�N���t�C�F�	7(��Yߘ�:�����D�*-�rCe� i%>��|�$c�"��$gX�>�6��G�LG�	џ$&�t�I؟��'�U� 
V=L#�(PQ��*x ,K��d�ן�n�K�\4�W�R"� fe�h�a�ݴ�?q(O��"WI�����O���<a�$�������� X��S"�	'v>H(r2�B�K���F&Dx��X>E`���
%�U���ʺH�0�C�B=8Zd��B�\�.��`*�bK� PX���eD=#q��n� �)bމ�dC�?�b�@�ǐ(�������	��W���K�O�c>���OH�T�{�!� �K��
	���߶���O��D�Oz�$:�3}�hM"r����/U�Fi���A�G���D���q�4�?��iK�O��4W>�;'g�#k���2�� C�fUrS�26�	���x�I�� �I�?�������I�_̹@�ә-F$�Q��#,�� � ���bN�/up)0Ĝr�@F	�V	��2�K�-7z����*I�ƌ5G�$�c�ɓnL�����7j�	����3Yɰ�i�d�(�
pJe�'w|6a�'1�O��5�0;��1�D�6U�x���-�ON���O�����ne"�"p��6ax��`K�l��'�N6���'�( ���dӬ���O�����\��}���P�D�b�!A�OX�W�1���O��Ӂm��5xP�܁Tڦ}PCS�Rm�� T�"qi�A����EH6���q��8�di�-���Ip$CP�ſTߠ�{DGZ�B&o�q/��1�1AB�D|��O��?A���J������P(zz�(�S�I:>F�'o"�'j�3҆�"�0��1+���@
��[�k� l� 	Qp�Ž�&�
Ԯ0�?.Or��O��d�O�ʧ6�l5��d�~Q�Ɣ�̌��Z���?��)�= �� C�[���� ٽ���C�$�*4��� F9u��A��Iߌ��F7H�x���:�|�ATBSp$�&P�Ʃ���?}ʀl�q
��4N�_��mì5?q��O��d'�'�y�.\6�I��Y�D�&T�Ǌ�(�y�D>s��!�e���=h�C�B\���O2�D��雊ZQ ʌGjr@;WFS�X����'���'�R�B����'�R�'��}V��a��[e|E�͞
��H�3ቫ(9�7��>^�Nz�Ǵ|�B�$�	��"3e ���X�^CҔ	 )�zRĖ#Ђ�y�E���S1'D�"íe�Aysl��r�I�$^�,YԂ�Ӧ�j/O.��E�',�<��?ӧ�wH
�>����B7Q �ԹU��ɟ��	~yr�'$���':ل@իߖ;���a؄6�����?AT^���'����'�!Q���T�e���ڥQ�������"��'��'��`�E�	��ϧ$cμ����+� t�ǳ(�l(�e!A}<�G,��>-�r���XF9��jD�{� ���=)���J_�5��P��S;	�4="�m�ݟ����R@�hҨ{��6�JW�|`��O}&|�QA[�pEG�"�V�%�`�ڴ��iXđU?E�I�w�DŹ�e��r_Xs���+L5���I؟��E����|"�#S%-3�B�AF�w[�	 t�V�8��7#�*c'@��C'�*Xj�(����m�T-�jŎ@����tLʏ1�>D����M<�(z��V��џ��A�O���(?�$�ݱQ����ԥߥr�V�Q�MH������h��E�1��&,@�y�+�$������ �D�3A�� H���&�x1#��Orʓ�l5��i�r�'/�<��M��$��X��� ���A+�x�d��͟�"&����d�%?�L��FN*5e�%P��M�d�Ӡ9Qb��	Fs:|J¤)H�ɡ�.�hB�(R��ԳW�ƗB��r�� x'�'>l:����t�����A$�\�'68� �}��f@*�'��.Y)͌0	d͘6_����wbP,�?q���:�j���F�'�x5��k�~�����ݱ�4�'S쥣#i��^,&�J�*͢S�f�[&�iu"�'�R�B#I�Z\h��')��'�=�r��p�;��u���O��p9��˴*��q��m�,��x:R'�c11�Z�Oΐ���+g8=�B,�92F��. 	tq{Ŧ���e���/�1�$�O�l
�
�r6L�B.�!|��R7Ml�H�'�����Z�'��'^���a��$s��-ـ�Lm��8#�"O��b&4P`(��es}���\�|Z����y��Hyb�^�`����C)U�*�3Uß:Q �E��8���'�'��T�'�"7��i��ХX4�xY�
/O���cF�6M�勴Ń�%t@��KL�fУ?�e��K�� x1�
�
��M(�d�^��hRL�a�4�3��"#��q�4t���9�dD��`P�n��Q���-��r�kų�?Y���hO�#<����UDTp�����������Db�<A�H�'3�*�pB����>P��C�I�M���򄆢w��oF�t	M2D^İ�(�B~L�I�kο�?))O��O��#_"!JF���eb�l�`i�����hX5�f(K�"'�2���QZ�� $�	 ��p�uo �(!g�oh@uҴ� �l�c�Ӟ(:��Q�@�;M8�Z��d]&}�.gӦ��'�Y��v���;7��'Z)���J>��	6�4���ل:�`�kW��e��'*�{Ҥ}Ӗ�9 Ǝ�K��rH\`?&<�@�Hʦ��'?.�a1�yӒ���O"ʧ;��C�?�`��	F����r��Уz�,�����?AqֳT�ֽ�dʖ	*�� b�����|�g��Qy>��C�[���c�+؝��d���q��L�������'���aQlݼA���"�Ovf)�� ��i�M�%�Du� ���O"�P�'�7�Y�O��)��c�B1���5�� p��-��y�	[�nLr5�Z�0/j1�%܉sLax�mӢn�m̧E��m9B��;^��9a�nݟO���R�4�?�+O�M��������O\�D�<�b��<P��	Y�KI5�	ѵ�E�x*��+V��
2ۛ6��)�8(@Y>)���K��\ `3��T�rEze���s��Tx���Qx����W�\n���EB����~��ܸ�8�(�ѧ�1t����L0q��bӌ��'�����ϟ�'��(�5n�Rx��	�R0M������'���d<�O���i�Y�$����i���'��6cӼ��L��OH��\>�q5�N�G�T ��̖J�����s	�L�v�
Ɵ\�	֟,��#�uG�'�3�j� �ى8�\rŏR�SY��yD߅V�B-	p�-}��ơ�>�+@��<sp� ֽˡ/�
����K�4� ()�Р�>-P��5(���`�-�@�2P"��C;R�%=�"�f������͟<�?���;�B���D�� R%��-��_�!�dD,c��`ٔ�@�a�`�+�,Jg��'1�6-�O
˓e��4��T?��	�c�� f*�9I��a���G�@�F���ʟ�	��ş �I�|�TlA���鹥'�+{�DC5/�B`�%�0 �,M���z��A���%Mh�(�]7��␄Zh�I��M�d��2�*A�:���ær�rm�K�j�qO8�ӵ�'b"����T ��(6�z���)6<�G	6�$�O8�����db��CMq� @���*l�����Oḻs�[�U#�E�Q+�?���p�'�	%]�Xs�O���|Z����?��B�af�a�H�0d5rlh���#�?��hΖ��Ee�v*r��DN�f�]>1�O��53���0w�	!�킴Z���c��db�
�S8R��� ŤT檔Ke(�Z���ƅ/�iM`��7�[-�4�ٰ#�>0��7Z��d�䦙��4�?���,9NbA j��sҮ��T�>��V����ȟ�'?�8 ��V�x����a_�f�*"-;�Y��p�B�Om��+ݻ}h�H��e+��0%��Ʀ��	ȟ��	�N�@VW��0�	ԟ`��켛��C�$:P*f�@��x�a��zz�x�1�1U�� ��N<xuFP�|�K>���-t�r��7 Ío,bA3a'T�
�l��/S�Mq�X��/r�Ya�Ŏ���ѓa��hd7�dS�B�	g���!ƻ�P�ؗ�'���v?|�$�Ox�,�I
!v� Y��Q�;舐�⋶Ȭ9�ȓ9,h괪�x!� ��0S=n��'�"=ͧ�?�,O��4��N�5�g�}�����eʱ�$��O���O��$A�[���?���8-�D`�K�8&��wI�	�N5k���B,�d��1x�x��c�{��?�d�?h���(N�*Y���bd-��>���v�Xh����/C4�?yش�����\�Q�j� k�	,��Ci˚�peɦ&D��,�ش3y�'���'O�O��@CG��%�0��qg�=4���Q��"ړ�0<���Ŗ^a��F��	A��ML�I��M�A�iy��7e�d�۴�?��342P8����5���Q�I�g"(���?��FΛ�?������'L<<�2�M�Vc���[؀1�2��JW'&Naiu-ێ#џ`��A0k�� 9�@�[�0�%�ȐV(���V�]�8��Ӏ:�4�Dh���?�����$��``sI��Y0����i���'%��'��S�N&N�� �LE�����1��%��Ӈo��m��T�Y�?�*O��������ܟ��O$<=�'FF���`DI!�Lw� ���'�b*^}(�4�B�jH��� hg�N�'���<�،p�K,(D�����ˑ^#�y"Z@��TЬ����_!X��^w�2�Е��3���J6�R� �u�<�*��ɼ��ā>t�ROq�0�G�T?�P�{�Z��X��!�M(%�1�B�'���IrjɊ{�"8���?r��,�`4��!ԛf�pӞc>5(C��(�
�06���Z���yu˿<���?�R���'������?����?Y�O�Z1��ʒ� ��h0�9c�N`#���V��Ib��® |(*%�ɍ�� u�'�v�3d�L�
�"w�ܵq'�m�uq�*��&� K�&��Q��t���7-�lt���%�4�*�`�2�ܫ����L���⦽�I{T�I�	W�gyr�'�Qi�Oό|�ސ���7t���'��X���R�g�$Ƈ7�iH�W'	[9Uk5r��I��Mۗ�i��'4���O��I��)�n�;��xȂG�T1,��,�_��u�	՟����8�Zw���'��i�m!�)`f��8�,�B%%�Nݴ�S�'�9	*��Q螲`<���D^!(f�h�%�1q���*.ȀT3�E��38M�fF��k���x�+ĩj^�0��9[B�O� ��C�,
.C?Άe9�*�)a��'���D:§"�~x�ѡ�vm��!i�%%��P��]H��d�  9�(Y�e�wt��$�Ԣٴ�?Q+O���A�M�d�'��Ĥ�(:���W�m[��q�'\b턹y��'0��� ��g[�I..U8��OX�Q$?�V����B�dBДb�'yn(XD�X<Cr":� Y�?d�8Q�E�0h >$��&V��i����:y.�5僎"ּ�=��AGٟx�	I~����s{:dh�� O���+W����0>�V!�r�8;�(ˢ�v����SP���b���T�K��	�gHT:�噔ERV�	xy�mT�[[B�'��P>�"&�ş�#���&_$�a���
�^p��M�ß��	�e6=��\���)Q�'�O�SG���:gsЄ`w@�	1@�J`��>���J)�8#dY�X(
�+��X0��k}�H�O��<[wcB�����fƤ{�|���O8M��'�����<�%��;;c"�r���$a`Y�
I�<�ׄI�Nl��iQ��K��!��N�M�'�Ģ}�B��4JP��U�XH*�X�ʊ�M����?	��Wj"e8�dΗ�?����?����y'���E-X��W���O�H�A�� �lDL�P7�)_d��$jI�P��಍��|Ҫ(1V�-(�%�-H�0� /�!{˺����$:NX�t뎜�>Tk���t��x��|�`*s�� ��*�k 7�� �VG��4�'�'��I�0!&��Oz�=٥��Q2(��e�/�$��d��y�E�so
c��"��(jg�H����S^���D�'��I�I���`�NL�T�M[�=P�!'����	�|�I؟��Xw4�'�2��SvШ���4X敉�I�����$fGs,�9��R�O��u��It(�Vڙ�~AY�!˱$�B
�c@WC������px��ыH)&Q�lD{�Ր~T*�6�U+Mq�o&i�J��P^�鵑x�Z��!���C�#CHx��瑧-4\�րU)�ўP	�
7?���TP�p�di����b�zr��F����Ot�l���$�'�ʘ�6��~��b@@H�e逋U����7|[>����?�c�+�?A����d�5Wz9q�ޤD5�ə�B�)k�TdB��O�m��H��K�<���/�џ����Z���W��L��.����2a,�9jX4��BMN��-mZ�ANFţ*���BMFY����`�'��f�9,j}YV�D�/��1O>i�)�F@�4d�%~��MUB������?���۫`�ዐ&%J���"���ؖ'�j�2�Jc����O��''ߚ�r�Q6F��ȏ�:9��x��� �`�����?)�g��el��z�
R�O\�a�b�.VT��V�L>��z��4��6f��*	V����O>���	8]`����K z� �Fꖨw���I?� f����3#���_j$\㖮$?�'F�����N>E���Z�I3F�Ԧ6����ѩ�y�Ě F��ӈ ����D1��O��F�d)΀k����Z�����a�
h����'�'��P� CJ����'Y��'��.R�9)�y�no(<A��j�g�����:d��EP�v=��.Pd�>�����l���~�L4Zj�r�=]h$�&!��tǊ�i ،�
S�F	f{�p3���aK	\>���p늕�΂�K2��A���F� O>���՟��|�<!�$���L^<7!LY��d�<�T`KC�B�%h���|dyǍ�ty��(��|:O>q #^TS���%q�͘c�iϚ�QbI��?����?�sR���O��Dg>!�@�.�J���_�p�{'�W�+n�$��II��REXƪ$G�������Q������^����AĐk2Nc�ȍ����a�{O��ED���\`	S� �+~Q�L����F�nb!�� ���)R�;1���\`���Q&R*h�2u�G&9Ha�';D���E�.}B�D��b3��9i��<������'�L+�α����O��
�%%�1�I@�+˲a�d��O���!����O��/Q2�C�̫;�b���T���0M�6x����A_?Nz�[�h�צ�3�퉖(.@��M�>-L�)'!�i��J�k�1���Ї�]�L��K gK�2���7a�}������'�Xk�-pd�ꛄL�D�J>�T�
���15J����ğX6������?�$g^�4���#	�5"�����˟4�'��=�u�'/��'#� D���I�&�`h§��N��)Hw��5��\��؟Hk�,�Ci�Hi-���5P�)|�(��FO��N��G(�"v+O�|c xY4`,��䜅>���C��$|qY�I�cļa8��  ���O>�]�RM�"�Q�cV64��9!�O�IR��'Zb���<9�nʩE6�Z�)̜|-j��GA�<y�K
�Dv�)�&�������z�'3��}:%�̇P�� �w'�fx
���^�M����?i��;$2g���?��?9��y�Ġe*��0�Y�,�T�Rro�^ 8󴀾>!Vd�L]VL�|�<1b��;C�ၣ(O�t�Dx�f�4��	� R��d�-d~c>c�Tj�� D���H�B�L��O��!�Z�	ӟ�G{���2Ң�Y'�A#��*e
�U?!�$ݝO�a!v�U
���A+@$j-��DR������'�0�2̗0f��(��ĵ{�
0��!�?IG��j��'��'2�wݝ�	� �'a��� �k5Y��N�p�(a��*8���sO�w�:��i��q£?�X�0�Pj�6
����{nb]��F�3���h�eӴJ�!��>)	�#>�R&P��*LQ$l��_��� `��x����l��I���@�,��}�g@�6h=��!�!�DL�%�^8GI�y�~h[C!��o�'�7��O:ʓ+v�� ��4"՟(s�p;g*ۯrt�4�vP��?*O����O��ʈ�%��I��5E`�c� џ,����p�>���Eގ4=���R�9O�9*f?��$�C�X��)����,�	4�@���%J�r���Ԙe)�'R�T1�E��0E�� �5��O�����q��9�a �vK��8p�=�����O� c1�M!s!&�*�d���k��'�	:b�����	�|��Κ��ק�N�0BR-����̻���?y������!Cn�.	�BYȧ��.#ƃ�?F�$59��2�p����1#4eE4���W���F��+�9�B�`
�y��z�����"'��'u�>�S�? t�A�
��A�oS�i���V"O8ܺb�T<m����'>غ̂���7�h��`M tJ,hL�<��� ��'.�� �4�Q�@�b
�=���OW�͜M�c,D�4$�ۇBi����뗛q��ibW�+D�,�vb�F����"e��I��D�4*D��R� x�!��b����l;D�|:�C�
&	���qBr�@�8D��C�dA
y� �R��pڦ�z�)�<��C�~8����#��iw���"MS���3/2D�H	�@�a���Vn�b�h��"D��� @ 7�"U����oϜ�ې�>D���N�[tfLR�L����bb=D������:O���3"D�t�����M7�O~M	 �O��ѱ�]%_�@�aڌ3\pA3"OP��C/� 9$�Mb$ �-	�%�"Oʍ��H�6�J�� �4@J6e	�"O����+0��LhA�]:�69"O��FcJ�u����ӴG�� �"O�s㇆����"�ϑsy�Ɂ��ɴ8"�~u��K9�\�Ĺnd! ��m�<��)��.i��B /����W�f�<	E�pc�:��(�Cĝ�pn9��k��u�V��C�ۅ�J�Y��)��\Oj���@�Ne�qi��p|2���}C^��Cݸg�J��p�M 7נ�IS�*"<E��j��>�q�	�����D��!���+HP���,C%P��Ց�"_'\�!���'2ҡ�%B�9}�-�BK7@!���2@�hy��ˇ�;o8�*�*^;r!��RѾ�k!cЙ�~����]@����Zĩ��A�"�4���[��АЅ�M��nZcK�=Ӧ,����E�;�?9���=m�N@��_�|��s A�v�d��`M�$�֥��/my��I���I>wה]�u���7Vv��f�(�<=�f�2���6
DHZI�7�κM���y2�7ʓ��7� �z�;q鋕\�l!R���7 �8���4#�hu�&Hg���)H�'�Ԁ����v0�)Y5!d�� dh�w�ș��9��Ie�����睺)b���`f�"0���:�Obp�'S��ҋ�%MN��i"gZv�V|*(O�I���O����O�ʧ0�X ����?с�*Y6Yq�/�)>:�����?����3���끥�*^�������I*擐kU4�y�/�_�Z�Q��.M����	0� ,�L��l���@�k<�P�(M�d��c>�s$���c�H���	;z-�Nj���1��O���1?%?��'ܬ������	��I�'�@3�퍛Y��hEH�#5�a���E�O'X|�BFwb�a���7�v�I��'"�'.f�0r˓ F|��'��'����'8�Y���>�l�����0�K@�.{���܃`��X`|W�?#<�Ej(FZ��ɤN�,� ���i�T9[�%� .���4hJ8���O*���'�����\mYt9����i|��g��q(�ɆV����O2�=ј'$�=�����{�i�[�P���'�L�j��R�b�-J�tD��ow����4�H�d�<�
[�`E@�B�0:Ȳ���R
PQ���/�?!���?���J��?��O>l٣�ɦ͔��P�ͣa���(M�v��%#�J�
9t�k��MʦD~��P�6�,��+*Uc�Uh�eS-H-�)��<�r�{&��!<6e��DҨi��Fy�)
!�?�ׄ> rz���=$P
&�˃�?���D&�@�,�5l�?�2����)���ȓ3n���޸'@R���n��;gLQ�'`7��O��[��� [?���|�p�W���_l�y@'KW1	R:�$�"�
�D�O���Q|ɐ<XAj��O$^�!���(	'���ǭʤ]�8�P�j_�Ex�T�P瘜l���&剪]��|!҈҉U0Ј�!U�l��L���O�4^����$��sYp� ��ؿz��0K�0Q=qO����'���鞓R-��(\7�H8	i 2X
�Ib����0�]*+����FF��c�H���D?�O�p�'C�0����h}F����LYO��/O��ڲh����I~y]>��	�� ؇뛢$��yb	��|}��Q!"�ğh���T��E��%#N�i�mּ%C�>%�Qۊ~����#�@]�h�$�~������o�� ��-{�~���"V5~0���%z<0��O(�A�qkڼ�:04�Dt��'�������?��O�Oj�)� ���D�~���	0Ɋ��t��"O��y@ �)am(f���`X3���=�ȟ���E�M0���gڋ!�@c�OF���O�������"9���O~�$�O" �;�?A�$�8 X�@ȵ�S���]B�dӹ#*	C��h�(�/֭/v��˟���>�7$�����R ��T��%L�K/�Xy��fh¡��.�>?|N��O�b�8
w�I�-����p��c��q�??���ٟ��Z�'h��#Ub��L
SD���B%O�&O!��F��BE"�8/J����-R�!��|*����dƹ.����@��<���-���\��!�Ѧs�(���O����O@���O|��b>��b*Y;�֍J�"Dv�p���/�T"gdG�$a�  ���h����E2��:dŚ$t�-�قs�<�s�P��t4H�#�w0L�9��� N"�;)�4�d��{��#$�*�	�d=,����-ړ��OB|Bԋ��mq��t���e(69��"O�k�	Ӥ*����g_�aGޑ�v]���ٴ�?�*OJ��Cd�<a����		�N�āz-ȳc���C��K��?	tO���?Q��?��-4q�%c-L�_�ld+�	�y�����bR�|26c��'vz(�#���ȈO�`ˆx�&|S��x37e�ٚ��L>���&��F��Q �9p�,4Z��/�I8mf���O�al�ٟ�ϧLC�<SufL�	ʒuJ�O�|�Z��	��?)���?������&�~��	�n�dx�͆�xz���$Yʦ���4�LT�$��
.f�3��b^�)O4��O:�d�O ���O����<�t��8���"��A��Q�rͤ�?	s���'c��E�F�--`,Ж/Dh�.�x�BEh>�OV��xbC���O}ZT)�ҵ[��E���_HVT8!&`Ө�D�0���
&:�O����'J���r+,��_58�a����'Y$98�$�1�M{��&ߜ����yBD�������;`П���<|	��XD��(�B� �&��7�'���R9	��s�q�O���'�䚗U}��xgNA�`�3P.mQ%�'%B�� "5O��`�؟�^w4�D�)�N ��GW���d��O�t�z��zr��	��I�,� �?�Yw���?��0��p(Co[6j갊0J=c`X����1����I���2�&�x��4c�L�禹�O1g�5x�I�� rѡCb��!޴�y�i�?!��5��<�O���?-x�,��~��Rc�)=��D ̨R�p�'>�e�����+]w�20O�j0h��$7�?i�J�ȴ��BH�G� 
��1�F,TͦIk����������A�����|�W��%ji���
��4
*���Įx��`��6��ߦ!�S韘��4R��I�`rP�t��?؂}�!�+K��۴ ��a������?�n���)O�D�{X�|c�	�o� i��C jC�I���-,�a��·:�.�!��`���<���?Q���?q���?	��Uf���.�;P)�c��f4��0�i:��'G�Jy"�'��'<��9:H]�%��	{��z���2|�7�O����O,���OF��|����?9�HR��y���;)�l�s/�9$��f�'��՟$��X�ݟl��k������l�0Y"K�+���'T�yrY�pQ�l�?�z�F��c�V����P	��O��~R�C�i��$j�-^����G��'Q?�
*2�ҕD�K�01';D��B�kE=4�&a��̖"AtJ-��m3D��{C�
��P �Hz�+¡2D��E�<�F�����7�����*<D���QOٵ}�ѠW�?o��xА�<D��1��>�"ܢ� �;)ؚ���K=��?����?!���?)W�+�ԡe'�TNTj��s	�&�'�"�'�2�'b��'��'��~� l �� �H=1�ӡR��7m�O��d�OB���O��$�O ���O��ey���w�M�*������R��hlΟD�	����Ɵl��͟��I�(����E�Kd"��qKV68� i"W$F����	ϟ,�I㟼�Iɟ��I�p�	şx���V���0 S:���\V�o���IƟ��I����	ş��	ß��I�Y����W/�����>6�,���4�?���?����?���?����?1�nC�,���V:�,�q��	aQ��f�i�'	r�'�r�'nB�'���' �I*R��#s^��x�"��B�^�Aa��d�O^�d�O��d�OH�D�O���O��WGX8���1��-|!��ǚئ%�	ޟ��Iܟ4�	�����ޟ��	�L���?CF���|sJ$ r+��M#���?���?����?���?���?��gò|n~p(�(�0݈2��#͛&�'�b�'T��'���'K��'Y��.\\����=(��20$ 7��OV���O����O����O���O��䋋X*t+��ۜ5���ƅ<w�`n�t~R�'��	w�OJ�A�e�4�~A��eZ�r.�ķi�lX��y�O��O�N6pޕ9�l�J�Y���]i�i8��ٟ$l��<I/O�O�2,�r�i9�D�	$)����� �I���"�E "Ï�L(�3�['RNў��<���@�&��<��A�6�V� ����Е'K�'g�6�/�1O�� &�Ђbm�ȕ����ʀ�D�^yR�'Λ�0O��/��)�5��hH"��k;�q�W^�\z�̉�tb���!?ͧ� ��]w��	)e�p����z|<������q�����Oޣ}��@�t�pwM�q��DB�`)H�DU�	�M#6NPY~��t�Z��S�:����g��b���ZQ�� !�!��?!�4�yr�'�M#�Or��ʊ
���A\wM�y��j�4����L�tv�P��d�O:ʓ٘OY���0��%��,>V�ΑR�Ư<���i���y��)�aN�Y1����I�«�A<�'�2�i���-ҧ+VP���m�;�0��3MF�E�d�B�J�P��'��`��4���]�pybݽkG�d�'��6{!��srə�C�R�'�r�'���'v�	�M��[ �?�#�_�s%`�;�o�0w(��q���?�5�i��O֕�'.B6m�馕�=z`���`���A��i��05�V4O��$S0`g���R敭3�@˓����w�B���Ǟ%3�����!������?����?���?1������f�f���o��(K��'02�'�R6�t��$�O �l̓JgZ��R�E�(�*D�P��L�.����$�ͦ݋�4�?��J��M�O,U�cZ6D�x�B�BP�� Fʝf�4#W*sQ<�Oʓ�?Y��?��}�t0�LBtA���p�_�ax������?I-O�9m��^����|�I�?}̧wB��a�*k���X�e�F-�<q�Y���ٴÛ6O>����{RM3���,p0ـAK5�qa� ��,�ah�<�'Wjx�Xw��O^��A�@���b���W�z�����O����Ov���Of���֛��K�]b����:+�@�5��5�l��'�dӌ��&��A}B�n�B`Xpv�hթDQ$Mۥ��̦mڴ�
�bٴ�y��'���i�G��t�2[� t/A�ajEz�߮i�.�*W%�ş�'���'#"�'���'���?��Ԋ%!B�PĜd�cG_�8` o�Z�(L��ӟ��	J��R��62OL��s�>RIP1u-2�h�רaӎYoZ�<A�O�������d�i47�`���S��.��8�`��=zy������L��̘*}�0��埌�	ş��'���'Q��[G��!
Hv�j��V�n`�B�'mB�'O�X��Y�4�(-�*O����&����F8(�dze�F7c,�O~�D�s}"�{��Uo��<y.�9�s�37΂��AG U�b؋p�'��*�? ��[���so��?1qb��ߺ;g6ONq��Y�r�I jQ�Tٚh�I����I�� �IH�Od�䚬	��̐�!L0e����!�ߚkCR+m�D���O��B�����h���?�R�I1.o�A��)�1;�0y�T�W���K۴+.�&�'�D���i���O��1V(��L��9��]�&i�&
�i�\iG!���'��'�b�'���'b��'-�g�%X2:e`��*yG�@a�]��XݴE-t�#��?�����?I��,$�|KP��U'���e�G�I��MSR�i!���(���$����h��5�b��$i�)�f�֛L�m��O
 ��Ho�D�s@ �u�=��<yǪ)i��i\�B�3g�2m	�����������	���'Ƞ7M۶�����AsF��ؾr�<:�Z������?Y�Z�@��˦ѣ��0l�њ�"h��ԉ'FVC㰤;�#Sަy͓�?�a�S� ~���u�����R��݁^�l��C�N�p#V�{�~���O���O����O�d3�'z!����
A=w���V�0K<��	͟��	��M�g����I�Ϧ��<)��ę
K�U�a-V`?hP�"��<��O��o �MK��5(�ش�yB�'�J������)O�,�5FЎg����6M5e���@���t�}�EO��\�4��ԪL�?SwC^�P�x0;��O�"1�d_?O���Zd�T�����KC�A�!��і(d��& g�Lը֊*%�y��AG�l	
d6��c�,��"ʒ�%\�k�!Ev�A��H 1�D����?D�:�X�ǟ;v=l<��ꌆGzP)��-�[iD�8��8���(]𢑱�cT,^z�xs��όKY:�
�řT��u�7�� q �ʲ��BJ�4@v�Q�C��ɹS����X�Iʟl�?��4;����.,�ܳ��E<�����'>��'� � �'��[>�Iϟ�nڎA2hq�R�
c������ml�x,O��$�<E�4�I�
rI�ƄK�\�>}�#F�3x�lI`��3aX�dk�j֌-V�#vO��"��2�C�f�ڹ9Ѐ�(N����i��B
',Of�n�����OnE�'%�NY|���a�FlYBw�ϠZʰTDU�a��ءF�(nÆ�J�#
�Zquxb�~<���ʪN,z����B�.�j�͌	Fv,h;w&�J��BMC�lʔ( �E��iS��Ae�G�:�l��g΋ZN|�{�$�^���ـiؑ�F���O ��:�H�	}�7M�O��$�O� �ǡ�p�i>u���L�4�AI��Y᥌,�J�xR�ay��'�r Y��'���'��Z���2����Dي�.v�r�'N��$4�4�����O"ʓrTHIC�D��E�Z��<h0�ß��I._nb���	����Cyү	�-1���'�J;M�Y�mP�#�-)���O��d�O���?��q��T�b�;X���YЩ׃k�d��҈]̓�?����?�-O��	7K��?���[�V�I��z�~����Vy��'���'[�I�X�IS����6 �ӐO�8 �P�m��r���?9���?�*O^�����U�!���۰E�,�bi�PjׅcF��I��Vy��'�B�����O���[�N�#6�(��C�$H�����'�r�'>b�'�� 5 j�(���O|�����@���Lr��芜*�6�Qd�O��ĸ<�����\̧�?�*O��=� �)��`� q���	�O�in>�CR�'	�'���&�sӎ�$�O��t���O��cݎ
�*!��:���<��)2������OmM�#BǂC�j�d�S�Qb�0`T��ğ��`J��M����?����R�'�?����?�e�Z���z�E�X�L8��K6�?��#�8�?�����4�\��N��<���W#�	�e�i<t2
�oԟ�����YԣG�?E������ɟ��	�!�� ���o� X@��:L$.���ϟԕ'x�(Y����'`��'<Ќ���X���bҷSz�8!r�'�g@�� ����O�˓�yG(�d&(��a�^�q��*#J�����S t���O��d�O�d�O�ʧ"�iKA�&K���^��L	�	�բ�mӟ���ԟ��I���)�<��M�̀�D�|��`QN!&���"�_�<�/O����O�˧�?A�̐(ϛ�@)E͑��y���,%"�'���')B�'����x��k>}P%띔���hD��<< dş@�	�����ȟT�Iԟt�O���Ms���?�fD�*`bS��\f�%�ǉ��?���?������OP�z�6��D{��r2-E�z� ��	�<��m1��Oh�d�O��$�O�)��-��E�IП��I�?�0g�ܓ,�� �p�_O��	�@���8��}yR�'�8D	�O��Q���B�huz!@M_8cƟ8�y�	� ���S~$�ش�?���?������1�|yW�œ&�b�86dBT�d�/O���ɾn2R��O��d'��)5z����_��X+P�$ĕ���ПL"��	�M����?Q�������?����?������M*Ղ�N������?)���>�?�����4�H��D��I<_��a�Ђ�.�!�cE����oZ�0�	�kS��?q�IޟX���0�i�E���8��Ҷh��a$����'��'��`����$�'���'���j⊂:�8�i��z����!�'��A�=Dd�6��O����O���Z��0O4x��ؼ|��(n\��8���<�� �<����?����?9����I�jڪ�bΙ*3�=2�NL�$� P��=�Iϟ������`�����?I�F��e����L�	k�5C�"�;grN%��?����?!��?	���?aV�D8q���[����5��*t'�����ş���۟�I럤�'n2C¤���C�Hb���}`F)�ri�|�D�O����O��*$�CZ?���e=T��a�	���b��	�;9������'}B�'��n����~��A
γ�D��eI���)���O��D�O����O�e��
�������?�9`/�N�X�!g2o��,�5j�러�	oy��'Z�˧V�(����f��W�zV�D�l_�@aݦg���'$����7m�O���O
�i䟄�d��#���h��q?�D�
P�F"t˓�?�Vm���?�M>ͧ�����7��Pj�Ih�ܸt��D�B�
j7m�O��D�O��I��$�O6�$V=��곾�p�JBL�`n���	,H���d'�4�ܒ����K6>�̄2���F��0���`dioZן��ҟ`�Pa͟��ĩ<���y�C�
�ptA��E�/�(��U��?���򤑯Oʒ� �d�O���B/�
����gq��9�/��c�����O�m���W^}"U���	ky25��`;"�_�._���i�)j$ۃY����i�\�'+��'�b�'�b�.M	�H��6�ld�
V��Q���Iʟ<�	@��fy��'i�l���F����a��7BK:�2v%��y"�'��H�Dr�'�R�'8�@��Kt��M�Q�J �.���_�K7�ӥ)�O@���O<���Op��<���2���'/�Y Ȑ*o�e�K�Ky�����?a��?q���?9��x0X���i���'����4NÚL
Ǯp�D1�"Z��������ky2�'�
���O�r8O�Uq2M�z��Բ��	�a���'�r�'>��'�e
�#~ӂ���O��$���y�(�Vږ��2kE?��rA�O����<Y�b�,qϧ���|J"���b� ��7�N��,�����?!.OT���֦Q�O�b�O>�ʓ�T�
)�	@rP�[���
3���Ꟙ�I-�l�	i�)��"����7oے4_p�sdg��� ��� mZ������������?є�C�tP�h1G̽q�t񂵌�-�?AE��?)O>A/��˓�?�feeUy��8i�)�B�1��UmZ���	��c+R���?)���y�΂/r�l��p*�+h����;�?1O>�cn����?����?)g�F�&��p)�
)x<����?Q�q���Pe�x��'���|¨	5:�dU������I���0����`�zy�'c"�'��I��e#��6U���Te�8`pl� �Q���'��|2�'��ꑏ*F����lX�Lx�q�dG�1��p�'��	џ���\�S7�|d��'rެ����Z#.q���I:P��'�r�'A�'�b�'+��4�'4�M�%I�j�i�DcQ�=�U��Z� �	ٟ��ky�)[O���t��Q���бvG�N��8օ�O���,���O���Z�lsf��<qw�Мrˀ)�g���
O�)U �?����?�(OnѪ§r�S��,�S=H[��!S�Vt2�飰�I�6���$���	ʟ��G�؟`%��̧,T��C'�'�"�S�D��)En<�	yy㙦"�6�|z��B0U������
~$�99���w&�q���O��$�O�y(se�O��Oq�~�J`m��w)D�#�m��0ɑ��'l��(d����O|����$���I4"�R%'�	Cd�TkT�#C[���	2��:����� ܰ;�!z^�R�܏^L� x�m��d�O����i��%�0�I�XΓq	��au��Q�|�T �~X<�	^�Ɉ��8&?��۟��V;���&L&̀��цχL H8�����H��	4��'\�|2�QA.Y1%�^�D,	���W[��1~8�yyr�'��'��I!#}l�aHR�!��p�3[v��*G>��'G��|��'FB΂���p���^�Ҝے�>%9Z�H�|��'R�'@�I�i!�Ds�'V°]ap.�	g�N)2�X>m��=�'!��'��' ��'������'V4t���^�()z6Nׯ;��DZ�@�����Iiy"�P`r��8hf�
�Jc�TSOV;A�B�0X�B�'P�'@R�'��(q�'"�	�n�ĕID�Q�R�(���	o|�lZ�2��q�d�S [pF�P M�ض�S��I�!�eG�����7�
�)�d��q1�ɲO%d�����?aI>Y���?����R��	�'�\+6�:�Nj�P��0H����?I���9O����Op�$��`О�B������"ʀ/IA��4iG�֫�O���O,��(���O@��	gnB%��D�$�~�a��#M�쨹e��8R�!��`s�XrT��R
���0A�:
�ʌ�;��Ak�wJjš�$ �X
�M��Z9u��z�'�q��jH"b��x�p�˾{o��
 ����Jʌ� u�������$I0�K�r���dO�oG�yJ�����c(�0a��Qϓ�!�2�:Ai�"(��ܠPa�!)���2��.��}"���9��J�*��5�b8z���,4B����ܚ����VT��'ˡ*z9�cjŎt!��B`ȝFu����O���O~����M�p���7�Ȋ���`�����א"x�q�qF��^�k�o
j0��%>�=�Ĥ��J���G�8"��	;cf#�`Mɗ2�5B���#	Lp%>��=IR*��h9)�d��(u��-�.�T�	�S����X8��9�G�Qs��X���c�I�[x�B�	'~L���A
7���p��F8>b�����HO��-�dHs��mа�"|�ο@JE��F2&0��O����O�m���?A�������L��X�Tg��r��ۃ���F��ȅ-}�"4e��E�Zx�'x�	�ħ\�~a@mVt��<3g���Xsm�	ɤ7mV�]����è0KH}�F7�D�0l��ϧH�0��o�9{�������=�IU�'S�����ӆG;r䳕D��q����&\O|c��S��H� tJ�)2mY
���qS�&}��e�*��<�4LW�X��Sԟ,oځFR֙��IǛj�h=h5�2[d���(;��!���?q��FI�Ae�U�(�&b�(<d��c݅8�ҝ�p-ޠN3X�IPcL��"?gh�\�Fɫ��*Ph��Ǐn��XFH��^`%���,bE8 A%�	�C�\��O�J<�PD�d8��;��*+,�Z6�>Y� ���2 .U;;�6U���K��Ƽ��	�~�#ğ�N����9l�Xʕn��_=r�X�b��r�ixb�'��ӯ/F����ʦ��BLvΡ��	;~�~��/�	�?9�#xD0���,R�Z9�2���?�I�a���@�V0�$�V�l���>0�N��r�]9I�h��6�i�O"9:��Ȝ7?�铱��O!�z�O����'�1O�>U�TaD�>�]�4��
7 �̱5D�:��dP}r�%��/q:4bg.�>Q?��DOP<���T"]�"�i��M�?����?���c&����?����?١��07-<y���+�␍����CF�g�rT��m�$�?����V$8J���}R+�3�¥���X���I�쀵��]P��@DQ* 	ӝ�6�*H|f&	OС�'7��j�*��$;!�B3�
}H<q6B�ğĆ�I�U�*y�a��w�Dđd�N8BĈC�	�5c ��@o\���i7��<"������HO>qp��L�X�����I,	�cץ"J�I��!�4��ޟ����u��'�1���� �#SP�Ep��]�0Z�s�l��-`Z�0�Rtr�zC9<O�qQ��R�ln�F(N��dU9r��S�S��z� �)#j�3�( �԰|j�	3�{2�X>�M���M���K��R^�k�%	�`R!��x�u��E �����m(�!�d�9D���K3�6��)TM@?&�ћ��|b�W�a1�7-�O���x���@����8����#荧Yk�L��@_͟(��D��P��̟�xr)�+\"�Y� �D<iZt���є6�:�R6jg`���C���M�8ҵ�߳Q��<!7* g�-�@��#}�X�� �3e��m�%EI%'���S�Aڨ��p�mRHTz!.�I7+$"���eܧ�����L�q�-�0蝚Z�:�� �$���)$��ZbN�&�A��I6�~RkD�F�p%��[Nx��I��2�E�2�M����?�-�@�s��O�7���W�0(���V���� �h��	���
��m��*�^�*Be+V�*�t�p��i���K8����`&����,R<�@���Sxz���i),�Z�J�8�}CSQ>B��Ʈ=a�Tp,�o0�񲠷>1�꟔#H>E�4苋*�J$��"#,�)�F	Q��y�%pD[7�(���ha!J��ON�F�$�?_��E�U���1�-ź%��d�O�����&0����O����Oz�䇺�y� ���Q-����*��5gv�¡F�4.�t�	 X	��A���g��N��R�e���eŅ�M���H7�~R�Z7G�¤�;��DU.E�����mם#�`5��OT�R�T��,O����'ml7M6&��N��)�\1vm4J��11��̬C�!�dɉ(���0g��}��aRo̦���[F���4�'�,���/�7�b=�ua� %����
;	��h�	����	۟�	^w��'�i�0]ZM��76�YC
^�E�Tq�V-�@���&��%�"8ǓqZPDcI� k� 
�k@� ���B�IFe/t�1��E�)�FS�$O����i����OF'�� �)�;)x�������ܴ��'�8�|�!��5��|�d��1()�q9�M�D�<�T���q�C* o����w��˦���`yr��7�x6��O��$a��,{��O0 8���  _�T�"����ܳ�@�� �I͟,CCc�䦩��yZw-@s���d���0��Y	xM,lэ��P#���&���j����׋̚V���B�X�5V�"?������`��$�4Œx��A�n{���8�y�曔 M(��WB�e�l�:��V��p?I��O{qk�i��a��G�w��>�qo��G ��'��T>�ل(�ß�oZTt	%�O�i�<X���>�6�@��X*����K���p,���y*����و�J؃�dR�@A�����Q�8q�b�0r��6H�7-��"��/mY��"f#4���D��C}����?1B�iJ7M�O�"}�R��3�zl٢ჺ-{"��w���O�����B����aȅ�6� ��I(�Q�@ڋ�$!JЄ�!�5_;Dl���&�J��V@�Od���O6I��� ���O��d�O`��wW*AA�$3�!����{j�<�K<y��z؞��$,�e���h	˃�'fʴO�ms��'�Fءi�8VxU���[�6G�y�M<�����4�
Ǔ"a�H;�f� ,�v8�C�33��t��]#� ��v�HA��:y��I����SC�	<�h�H(xT�Q:D!ɴP�XĪ�S�-N�������I蟤�\w�B�'��I҇y���H[�.�X[����>���^��?q�ʜ礪:��M����Bd��:%��yj�4�O�
5�i�6M2� 2]|��,^�+d0��5-�d(<�taO+���Ҥ�=A��4y�m�f�<���H����Ȕ�m޼�8��Y��O֦}'��b&)��M����?!�4N��l�7���!� 4Afe��>�()���'��0"�'\"�'�l����[��O�nת c��`��:�Li�@��+��a0�{�%9��F�4(���#M� ;��A��$kH�RLD$ݦ���E�;,z:�?I�EOƟH�~R�P>���։G4N|��&@_~�<�c�P$*���%�N(j�@��{��l�'\^���!N>v�a�q�TJ�%�K���5
,�MC���?	*���[�,�OJ6��=���!\�A�\�v-Ya�X�	?Et�A�S�!���?��u꩟��t�L�]�"��H�p^�u�tY��K�Se4��G�}`f�YD�u�OBh4a�iŧu����H.��ګO0�C �' ВO�>9���^��l��`8	�t��b�,D��#ޭ4#����ܪo�IAQ /��Q?U*�b�-��IG!�02VJ�j��W��?y���?	a�?r��@r���?I���?���w�Ɋ���e���hc��JY���>+��*��'Q����n��K����O��+�B���`�*����� ��K� ��N��|I��ѻ=@�Ok�5� �:����G|�Q��+��k�Z�։'P\e#�
�x2�$yi�$�=�i����6�y2�-8���॑9 B�Q���L>�~+1��|bL>� ����3�(�"&�Ĥ���$k��������I۟@�_w{��'��X�#t�!���V ���a�F5�lU�& ��qv,�*WDB*�����F�G,Q���^'^d�d3�8��W��#p$E�#�I�}����D�"t��-�2S<h�B� �0U����"�M[�'�z�p&"�y18$��㚌S���9�'*��b�cD� �&H!a�5��K��	��M�I>i�W>}����'j2�i3m��`TF�Ұ���+�� 0#�O��M�O
���Oq�tf��(�D\30q�Ep�L����&C��%X��ǭ0��j�#6Q�,��u��Y#���.k���8l�X���ܮ;i����K�&U.�z�)xQ�D��'�Ol��}�̈�1�P��G�I�G�sH�O�<��k�-�]�6OH!���pk�p��<��'
H��3�vW:d;��ڦ~���)J���QkJ0�M����?�-�VH���O\6M��`��m���Gx������aC��ɂY��T��y�S�L>� ��p���+0�6P����<݄ �R��t.�S�O�bׄ�_�h��Wa+fx�ʯO��j�'m1O�>1��`M<��a�J�K�PX:�*O�uYB�ܞ9&B��B�R&h ��(ڨ�b�P�]/OnHX���U� 	N�s#�ϟ���`"��R�]�h������	⟴�[w5���N������<I��K1˔�;v���֟��G��<ߎi1J|�>�2Ꞵ2o��Cb��&X�� �D��=�,�J�V�����Ϙm].5AI?ɪ�m��1�R���w\vP2�f�"2��f�U�<%�HH<q�͐��
Ǔ������/1�BЁ8�`���%�D�d�W� �&����V�
q��<C���w�	�JB�����%q�<��5�Y�O��а���:\��ӟ���ş̋^w�B�'��T��M!�ܲq- ��c->ʼX�hY����2�*��qeR�'�v�رkd�PM�A\�9�bʏ''6���N�j�"�CQYl�@q��+}��QS�r�	)}�6�9��!�t��0k�txz��K1L���'�4�w�U(�dI'��r@y
ד��'�1�4���w��E}D�C������I�MI>ѧ�о/��'���i��	����X���&��"�20V	�O@�b���O��$�O�E�vB�3v
na��?�8�He�j�6�jt�S'���{`L-2"=���]9�ʸA�B�#!lh�B�ײ|����pD�%\��Fo'[?� �j&"D��c�^�p�O@��3�'Zz7mߦ���ʺK�O�X� Ѡ��8g��S��[?	����h��d*"��v�D���M�1���'sZ���>�DAC�¢(A�i�G� 
c>��k,O�8#3�Y�!(���Ox�'[���P��M/��X*�	b� ���C�$@��ҟ<$�f��80�gD�o^xh(A.�;��I/��:f�x�J٨yb�DK��2�	o�����Ł(k��}��">VVYF
��<T����P���<uQ��� 
{a��۫"H��'E�Dx���?���i�R���U?�6N�6,����5J˃	��X �9}��'ў($�p��j�'<�0Q�"aNt���7�E��,b�Hb?��d�רNl�e�����q�0 ���?����?�oǭ|˼�����?����?)  t޵���#jXX�%�O�~-�w^�RȀ��5�'����mٲH;:��OXdρ%G��d0���3Жh��r��{���yn�@��ˊ�o���O��&�̯z|�;~�Pk��9)E���s�O� �@�%�y�g�O4����Nr\�	�ee��PI�K!�G�i{�(���A�;J^xr6c��{���y����|2�Ql�[�ED�ꨛ��F�KB����G�R�'���'Dn�����I�|2h�[����$�F'�ĸԌ�i���F'&S$Aw���<Ѵ�?SM\�Y=;b�h��-%D
��Ǘ��q�ࠄ&��aPR��89_���24�I�-O^6͓�nB̂ .AH}����%VJ<��'���j�C�$��� ���؀	�'���S󈍟w4��&
��v�I��9�4��K&��c�iZB�'����	;@`Ifb�V�T��A�1���[$#����O����>WpE���0)V��6�Vڟ֝�<�*�z�e�-�Nh���M!t"?I���-�<� w��gЬ�2��`{rM��Nמ$����ޜJ.ډ��"W&�=@��?�ɒt���&��y+�@c���>2_L�2����t�HB�!�<d�#eB6 r���B
|c��� g?9���"��S�!y��͸v,�d��E��o�x��w��J̌h�B�il�ȣҕl�Y�H��4�Z��O h%�<�Q�ȍ6wp�Yp�]I�����n�%����d���9��d�#�a�bƹn�-�4�MN�d�A!�ӗC&����8����GY��NMƥ��1�M���+�4��_CB*�@�/�<~ް�1��ZLL��?�
ۓp��x ����� KڑP�ҥE}b�0ғ�u���-����G �2fPK�nЬ[����O���Ĥ �������O��D�Oh�����y�����H��"���r�@��ēp*�Q
�BZD�ax�b�E2�����<�Бb&��'Y�Ir#)o\l�0�F�N_���'$T�U�5��1�i�"��}�K<Y���`��	9��`����:�,rvH�]@&C�� T��Lj'ƣ!���$��Z���,�HO�I(��8kU��z�L������q凖�F4 G"X�����O4�d�O���;�?�����d�T�B���I�@��Ԅ�e��E�)
���g�S6n,T�P��	�^��,
 Q3^
T�c�0	��R"oP�3&i��N.|��q�����vFι=F0�d#g|���W
	�O7��RFoH�S�T8�yH<Q �U9\Q��.1Fes̙Y�dC�	+����Ս�-F ) EG��f�4�'�r7�4�ܧ,0b�n�럨�	Ŧ��AB(_��D��&�0Fr�r�%θ�?�`�?1��?	��O3	�ѐ� 	�y|�M�ム@o$���� [�iRBɞtD=��9��e��3"����I��7S�����{�? ��)S�L�=|�ɔa�4����rf��.����6�I�@��d	fܧ��FCK >|��3�	��$Ȇ�2�� �q��e����5f�*9��I;�~2/K">�1���S<�}��'��p{�|�ڴ�?����%p�h�dj�P��e%�!J��S�(ߣ"VPP0П\����(5ⲅQ�M3�4���%���1�iLX�C$��\D�"���	���u���G:��.��LE�;zn"t)��C�!�a%�L��_��lP`԰���
�,��` ���d��Бi�R�8!�D���K�nC䉌7���$)h�����%G�R�0�>�t�S�	�ٶ@�5=٢cKR���	��?1�k�1pr��?���?1�Y���T|�)���fG8���ׂpY*�@����^�*6M�I^ح��G^�@ܓNN`�Ve�&��}`�)] �x���I_9���P�4���*<�����K�g�6$��ӳ���S�Q�
��Z�4k.2K<��,��ǓS��iön�U�ۤ��]�	�'L���Q�5D���5-Վ?�Ly��'rl#=�'���Lۅ���Ss���&`	:����C��&) T1��?��?q���Z���O��Ӽt������F/���{�iۄm_ %�gH��P;3)ӿ!�,ɩ��n�'N��A�H:i��z C��&o��q����.k$s�hC�52��� � ���C]�ԥю{�!�.�M�يG������!��D3����4!�D	�nLJ�%�*F􈰘�l6C�!��+@���$p������C�v���|b U��>6m�O��Ds�V�ʅ!��;�L� �+͎	�̹�cfU���Ed�̟���ӟ��w��&_	�iA]@���؀	��Z���G��Gʙ/Y
� WI��S��$��L8rبQj��Z��%��˽l���g$��Jb"���G�2>]��lD<DF�8��##	�/.�>y Ԕ	�+ݠE��m���̠s�FB䉶h��5h� �lіYI�1>A���d�o?�C�1_��8��'�h{���Pi�r�D_)��,m��X�Il�th���ix4��DK�
����O��k1R!����O�h�b���ɸv�)m8"���B�k�4���N�u9$!f�[�.֤M�uÐ����+����4K���H5J��".�����	k�� #*�:�� Bǀb�n5Aãݺ<�#�Y��w+�O�b�"}
%^;�>�#��V#q�z���o�J�<���F�"��Q��=�=х�b�'���~��/C�ZˮD�1�C�i��9�`ɩ�"�' B�j�a�p�'�2�'�BA��۰l��#�L��f�".3�!(#�K�.�:��țLh��q��"�p�'>��=���&*��x�n�/P,���e�3	D�ݣ�$�'�LAc֡�rCxp:I?Qo�KF.���w�i`��_"^$��"j`J<q�%D�T��&k�@`é^�}��xڒ�D�r�9��,T��Ak��Z����m�r���%l���Sy��� �#�Ӟz9��`��ºp�ByI�np ��������ӟP�[wzr�'�� �0@�`�
^�P���#x!�n��+���$�|נ%��U�b�R�?�e�J(x"16(�")]3�)X�/Ua�Fإc������]�g�p�jٴ���gjTC�Lnboڿ5��1����vI��z2�_�o��7�i��"=ɏ��J2s	�����G�H� yQ�#գ!��[�
 ��8�.	![�x�����=I���'Y��
��A��d�� z��-�v�1b�ď.�(O��=�O�樢��0Nj�2 C����k�O~"=��M��(��=D�D��SjG��zd�X��a�����'�C�	qlJ��	�pׂ<����C�I |�Nd���W�C4\`05�����C�Ɋ�˼Q����UG��}��9{��-D�d��hD.w�"�5e��C�e���.D���l�D��Jӱy�J��-D��@��2*D($��OΰF�X���)D���'��'7�1��@c ��ec&D�|�g�9�h�H�[vR̀C�� X�J@35��5'	p�Ӥ�8R��B�I(}~ZX���ӊ�L�!�i@8S}�B�	�!�T��LTO>,��4n_�Xv�B�I? ��5xa�=s�1c����HB�ɰx�.ЋH��e$�8*�LB�I5-ń�/$�|����v�l�ӓ�)D�h��4^�aU� "O D���ʘ�^]X	�I�4-3�?D��k��L@K����#��("p@U�?D�� ���$��]0b.<�"�"O�С�蕔��A)3OJ
�B�(�"O4����,F8��e �cx�e�"O�u��m�6/�.*f�Fx�ՑG"O��a���cʅ{����z�m�"O*�Z1�J#�0=�#��~��Ɵ�drb'x���1�xZwt��i 7?QGhӔ2�t��T� -u8YZ�$�y��4QC��OW� S�mp}l�R�Kp#8b���2��d��N4P�,�_�':�*����oʔ �/��������P@���CB�	+{0�"�M�=W.�/ �"����ݍ�� �C�2�O���"�xRq 7�[�(��'�V�W�ІqԠё%�m���b��/�yRmZ��I�B`���� �c>��H�D��:[�B�	���4���[${W���dފM��[�4f;vi��/KѦ)�W������J�0q�J��"�xϓ>�JN�،��1��A��P��	�i���`'�+%]r�8� }�R� �!G�V�0���d�чO��f�3uh³?Wb���ڒQd�8�f�.?���DOIr��@�c��*>B(N��]p\i����:ـ�b��F%.N���c�tn�,m6x���S�$�n ������0aY�`n��g�߀��6M�>!4 ��,��W�X�# �P	�k�1��8�O�\c�hA����5�v=�4�ӯv�0qa
�'�,ݑ�m��(���,�>V�xy����	��ӎ�v�CU�V���Z�lPf�^(q�*P�n��$�2�N:6��,�BY~�-�������C��d�� S$5V�{��z��A��뉥,>UBS0���gm�&^��Hڊ��
�%;��dSY�0Z N��+���T���Bt��(B+(_=g�[_f�a���O�F5J��ؼ%[ �:w�Q�W	���d�T��0?�Ƌ]dR01�^1 bfc�N���X�k�.��S��.d���E���ސ��]?fG����k��7�©��/�D���I�K"�!���)��!y�AG��TٰqꞤq�0������m�9�\���_&v����?�=���T�>�{�'Q�4�ԁ�S�XE �UN#2���>�N|
�K �����e<.5�!� y����L�+VR�{� ��,�'*Ь���@�I"& R+@n��E 5h-|�آ=q#
��r '�#pZ-��+^�3<�4��bE,<��CC%oF@єӁ" L�ïP��0?����
�PX�Uꍭ]��!"����<���E�X�����\�r8ĸ`���Nl����/^��)�O�� ��P���EF��F�œ	�'���*S��W��h�&͜;�T"H�,7y$�� ،Cn�Ё3�@�����3�ʈ�� mL��I�Q8ڽ�!�F�oҔ�Óg��PLa~Cǩ%G�����^R���@D%L�bH��{čJ�,��%PU�K�AY�XRvD�<A׺�BL��ՈOFL�̌ o�` �Ć�Ȅ�5�I����͘��-���Y
&ʥq��Nژ���H��Z�p������B��I��I�u�'|�)�3=B��kN���$����(�DP�(���#���#Gb�Q�̰;I�+�?�;>^�� �.�~4�!`G�FX��a=n�hW�����ˉh� h&C
s�~y�H�8\���֫Cº�u" XJ �&cO**��֧�$`�����+D�;���p=�Q�E�R���{�ƚ�xB"���h@�$l	h` _���Z�n�X��"W	<���{��������X�b	��$b��ˑ�C�1O�����ʉG��)��-�~�0�&�8���HTM^��PBFf��K���O6H��IGL �gaP��	�+����P�ع#<��;���%{�" ��)K	C2É=d�d�-�1,�������; :��3^w��}��w>� j�ʁ�Y�<#2�A�C2\��'�>�
�B�!��H�"c�g�QY_�r%iafI�HJ(H����0uͶ�/Q���HCĉ�#��`#zy��R-&f,�0��U ���֝�0=���L.�`���s�t�C&�7t��`B��w���@h�#<k�E;���!�=Gރ
��5��	����7.C4}�Nq9���[#�b�x���^.�,��Ɉ�y�,x�'�tb�5�Ųi6	��ܠ*|�9�	�(� )����"����4y թ�W�x\��/T�T ����R�U��`ui�&=�\I"!��*MHɎ�T�pTΧU,�ͻoR���Ç*�F�I���k�����*02����wyD�����/�ɲm�x�P��jF�X�O+4>��vjƌpvZ��6��e~bfYv:]��+1�T$jTgV��0=���CT!	����5�t��#]�}�M2�ǻ\�:1�nJ�f1�)���D�b����� ��IgB�x"�&ަ��y�4�ɺ	e�b�p�T&�8i� �DΤEd�Q���_�Nl���&��cE��BT^4^o��3��]�wg.Px��ܯEga��L�B/��$Y,b��[@n�7���cD�В,E�y���>�L ��[�D#1�r��.`�ӛP��r�H=mIvK	q����	��H�D�?	�f�-&¹s�"�i�}��j��łd�0��b�_�F�* �w�Q�w]^(0f
�=-]���JÁ��"g���`�&�'�����2�Bܺ@��J��԰�����6�@��@
��5>��
�21�$���hzp��F#�"��T��f�o�T�7 K q(NMx�
&ig~�i`FM�~��S�? ba�dgH�}��� ��ͩn7L�!G�֦Ot���ʈX҈���s�ny���~�`1EL�i9R�1gΖ'Lu��a�^��&�ЮȎQZ:�O�]zF��!�؛��M-t��z���u����Q���hy�6-ռUIڨy0��[9����w������W���Vu���9f�L�8'떀LӺ�=�&>W��h��P<�٢ �~�e�@�CVP�A�&*����Aπ�[��!�%Vd�B+ݯ�T�'CZH�P!%�	 r�.8�,���9A�mׄ����B�,̞!���!�fQ�L� �ħ&N�����;��Qh�,E�V�օ�Bʱ$�lH¤�ֻ4�^,ZլݩH%�CR�'��ӳ�J6\�@�c��Q�R�}����?بd�E���Uwr%`�'i�����3���@�T�v�{ޱpS`<5�Ё�aAк'��-
��8�OZ�{D�_�d|"S)G
|�~Dr��ge:��6�r�З�%5�(AsF惱��UH�Iƈx�r�)B��i�N�j�K	Tl�M;FΎ�e���P��DF
n"j��G)1��1s�'��B�d���6ξ!�U�\.�Ԑ(��V8�J牂\]�Ų��'ܨ��g�Q/M��b QUP��4�$,�%iÓZ�%����#��]qI|"�����\cF���࣊�2�1:�b0�p��'O�Y$Ċ�l�3��.dhtpcSD[CF��2`a�;w���*f�F43N�i6��ټ�׭�'�|��F�L4G�  �O
[X�D`2��Y��h�Q���
S�8x+��� #�Fuؖ���Iͪt��2ob(�bv�E%[$%�fD�"=�&�62�D�T�S�(��L:�g�"��tƁAd��A'O�d$P�Q�yA�T>�0�_�+���w���?	pecQ����="����P/�,���4�U?����ᨊ�Zz���,D���eB /I�f�HMת2�����L�]"���O%�~���
���g�'�ԍ`�0gKZm�4B�u*�H�
�s�i�Į�*z���1����1�MS6����'K9Wr���yW&$!R&��:fD8�3⍱q,$E|2�
%@��g̉ep@�!&^>��"V4C(pѕ��
S�I�S$D��AMң6�{V/ґE�^�����`��E�x��<��j�8�a�Ԍ�UUZ���烡��hte��y2��-�6\��*@�~�$�UEA��'�$�i'(L+��ϸ'�p�q� �I�ΌS�9���s�'9�<��0S��܁���WY��A�k�q�����{p�h�r�ڡ2�Q3v�Ca�	��D ��1df]	����rjM�$����ȓk�x�{eE��v�̭�#K�N���U�Jp #�ۍX�P�5L�=�����A�V5k ��RDh	�Z�(Td�ȓ��(��غD� �&F��j��h��^H��t�D����W`G�����ȓC�n\x�$47�t�dC�CD9��}�2]�4D�M�mCH�xЌ�ȓ;�z�r�C�")��t��MpR���o`|��g���)N&�ä�[A`�ȓ)�0	-�1X�`)��k��L��z9:l�d�@#8��@��]�G(��0hP �1"L:{/nTB�ϐxV�=�ȓ�U�.�7#��sA�b@����E6�M�se�M����t	�f�ġ��{v�頦R5dD1P5$�_���ȓAp�
�.�.Y��C��� *dԅ�"�h9�ƅ��#��x�5�8b���ȓ	��L"IL�xs�Q� ��u-`Q��a�V���ܶ{X���G e��ч�|/\���O~�<�de �^��ȓV���r�3;t�2�$5���ȓk[��8i���㤖$5�X�ȓ��̊a��<`�ƽ��&E☆��,�Is�~�9q���%Ӵy��M� -b�
%��B6
�E�����s�"�p&#�1\-Hr��5xJ~���}߮�2e����1(�@�@��L��z���z��%c�n�9Fa�D�ȓ�F��	^�B���2���1o�t���D+���#h��r8���,fz�݅ȓfh��D�V����(�-���S�? r�v�6Mz(��U@!OX��r"Ob�"��'`��7�W@}�<)"O|�,G-���(V��;Y�M"�"O�����+p��4�7�T)F�١�"O e�@��iy��XP��u�ЀJ�"O$���'a���qjų5�n�k&"Ozd���g��t�b��r޵��"O@���!B���j´y�Y�"Oh���b�"m���aϑv���h�"O�2����Dc���V�D�f"O����T'|��%
1.�X���"Of�22�?4�1�G`I�B�����"O�@S$H;:�P� B7>_p��"O,��ah7Ԥ�Y3.�v7*�KG"O���t/ܢ��٣`��4$py�"O�pX6��"gf��2_�A�q"O6���Y�'F�e��"����:�"O��P���m �b �4NI� "O EJ& [�Ne@,9#@�f:��C"Ob��F��<z��)�0M��N;"�"O��JɑIŢ����L�U��1�"O0�S�mE4g�~p������	�"O���V昣{\,щ����P���XU"O<8��Z�Jp#%K;,� �"ON�[�_�b�L%�U��K:"�
�"O�<&m��d�t���O)����#"O�mHa*��4@�`�n\9x|�(a�"OP�ӑ�H�V�TM��ĮJ���W"O�|ٱ&Ӝ<�LYt��`��+�"O89��]�E\x���S�]\0}�T"O��᳍��Ey(!Ф��!-4�1�$"O����l����µΆ ^+���"O����#�8(�p.ʕo��]��"O���N��|pU����>
rx٢A"O[3��
�v�i���L�ivp�� "O�=�A)����͚b��x����"OnY�J�8sb����؞H��x�Q"O4M邠�:IJe;'"݁dA�x��"O�-�Ӡ�*2Ԧ��OѧfL�9��"OB�U�3���S�g�죡"Odi�C��iǊ�Є�Ul �`"O"�P"lR=�^8�1�נ|M4Y�3"Oԡ��kZ	_O�P���"˺�1�"O�@c�#ʃfL��L�h�z�"O�aÕ)�yXe�Ӯq��9ô"O.�:�b�Q�`��jw̭�"OA;7i�.;RH�I&�����J�"O���"�P�~,0���,�.~o\9P"Oi��G�Z��X�W� ��|34"O����{�(�!�W)6�����'W��PHG�Y�ƴ��gڕ8-X8x!'mB`��턦{�lB ɉU�<��b*�@��Ѥ~����%O�M�<��þ?@İ�T)��h�e���p�<��"
�T2������z\@C���p�<q�&��S�̒�<���,�U�<����^��2���l�؁�Ƌ�z�<��A/�v��k	|��#���O�<��(��3��Q�
G��t���v�<)��az��h[�~��5����k�<���	6:#�`��g\�$�~��C�d�<�E�^9Eܚ�+w֣G���s��J�<�EJD�iR ��}0��qÓ70G!�;[<V�� nƪ.r��+3�N�s>!��"]���t!��
�2Q;4NY�}�!�� *e��Cu���$�Ҧ�"O$=���5^p���&X�d��"O�`�Ӌ8@���������y��"O��ċ�7N����/�!5���"O~�j�k�?�,����B�A"O�Q���c��3�!
�����"O�(yFn٥u�����X4?yP=[�"O�\� �;4�b�7l_�Q�Q"OD�
0�D`5�B��F�yN�X��"O����I�*��H�F/�@�"O�!cChd��g���9&D���"O��PD]�IC�9�2�%K"��2�"OHp{���!=Ȫ9�^�On*��e"OvPi�@Şe�tRr�V]0d���"O� �Z!Zn��JB/!�}A�"Ot�C"ߞU�%�OЦ~NjC"O��C�eO�]�y��.M#Kz�+F"O�i� �!A�X���ȡ[\6���I�$�\D��j܇v�!����%Ȃl0k��y�bنF�z��ah�(��<�q�Q
�M�PHN����(�8�I�SݼɁ«ڥ!
>\��Ex�B䉾��a�וbiD)�4�%���ݴ3�����,�Of�lZ������<Q�ih�ɤ|�-j���%�JaC���H��	�$%��	b�%�4��4dA�W�60���9���Ç�K(�$�	3��'��%z�esӠ1:�
�5"Tz��uQ���-ť:J؀�&6Q�T�;�䔵D�6P����;RR]����*b�I-/�DhIe��t�
iɁ��<�U؇�̣���H㥀�\�~a�g)N�=��=�d�Ʌ2C&�+#lU�On��� �0\*7lR�rBVT��n	!l�z�JZ?�nm���,S�:�����I-����$��1�,V	Ug1ȠED�c2yPߓL�D��5.�'E���3q��$	�!�%h����1�@�=�0=��&x��`$��� %�eEfR(�W@�$)�إ`0ěq��T��y1'ڪN�̥R`��	�>��OޘQ��K>T��
�C�.��'���h]�w�������eF�Ǧ��'�rdF��8��6�E<b ����L �$�Z��+*�X�$��0<透�,8�n�qAgL�G�J4K�朁Nx�Ȁ��V:W�ƕ{�T��ay�g�8�c�A�>$;ȴ��iY�#�H�r��'�Д�tF��H� 9�m��AJR]Y쓅�'��	*� B��I`!iϴkw�ᶅ̂'.^�����I��,z���fq;źS �� ��bkP����E�7�:$��I�$4 @2%I�eD֡nR?W�ޡ�'�@Y�(_53�JWҎu�^4h�}�k��W�ZP
mQ�<Uͺ�"M%�~Z�y��܆C�-��o�keU����F��l:��Ȣ<���R�A5n����$�5լQI +X,45�Y�b��
N��]�U�
�D0��@W+��nF�ӺGz")�.!"ɓ�΁�b}�r�Ob�ю�p�%b�e5`��3K|��帟�W�xJ|�0b���ҷ���]5cȅ+��ŚЬ��y��C�<<O�ĘԤ��9	�G����	g�ތl4�Xِo��;7�Xj�K���M�������Y��ލ���#`�-��dmS���O�U���kW���#,�:و��|�lg:؊�eH����rM/��Y����"�?�D�f��QLF�}��Is��Q
G�K,sP���dR#��3�
�x���
X.� #1�̡|Ӯ�u�'����Z>�	/7��6X2�	R�
{���G�ʏE��i�-3��dC��o�iQR_�\J�����������6e����pם`�T'��w0��>)�2!pToEwaʨ���A�'a ��$�ۦ����Q�g� 鑆'�W��a�B�ەL���zE��J�(q���m��\�pß���D�r��~ra�)�l ���9��L�AI�7��'SpQ��ե}�f�b�����O�D�b�ҒV� �h$�H�n|���4�QXւ�_�+�ȝ��p<��c��7�8��1%�:ر�k�_�V�y���8YӒ �Whp�~��N?�{���_�E(��2h��үL�'�@m��
O����"�:(�~�yv��+JB<�r�F�+�ҩ�f�Ǽ'��I{�ӱ#/(�tå?EJ�"��s0�u�ֆoKZ���	*<O0�q�Ʀ/�Z���Z�D���
$���Y����&��L���O|�D13R8yZ�e��˝)2�����>��CEk��Ѕ�â<��;����ɂ|i�9��f��aj�`]4R:q���j����ɠ�L��4,�t@B�t(�8K�,jL�1�SDӲ�$�򤞖Jܸ�ưNr�I(�{P�h�۴[W���A��u� d�q����=}ʟ��Cqd�#n�`y7�H�D��]��T�!�d�L�]aFI.n)Z= �I�M�M� ��5&�4�$�|��y�������� ^�Ðf�4��B�?J��i��'�Fl
���O� B���t���x�b�r	�)U�`P8���G��1$"�������8i`�'a 0��L�d+fg��!QL�2�oE�Nf���N,�"�V	�
S~��G���?��c�|ǚ����T+���H�>z�F�w�I���I�|����U	H��j��.#�Hd��c��ɿ�<6m�m?�r�֊D$��I��MK`���M�S?�\1��-�D9"��蕉,��D��'�1B	����I6�F����<c�M��h��?�%bD�~���wO� ���?F؁���^k���'L�dQde��]�!3��7OxD���[v?qt���y�+Z6&߲(�6I�N?᫟��蜤{��� ����(�6bCa|҇N����'��qK�����7�H9 �m�a/r�$��<���F�i��d���7>��e�bG�O�r���@����!Fy"��~�OIs�Y�d��n�1������;J�#�	ءk�`��]=` H�דE���G�~k��H�f͉�R�`�(=��J�d��$�O��SZwj�|nz��y��纐���׽)��
 �-Oܝ�D�w:�:�"��v웆���E����G�2�j�ʊ$�
��J�o��ӬU#�@e�9z�F�7hB* w�%Qa�TH��'�n�H��H�N&-#CGϨ!wLJ�^�d��i�i��j�x7jJ8� 0
�5}�fĴ0�0 b(�c�~]�EeQ��u�{&�M��n�
i_��H2	T*C�b�ҐA0`6���ğ���3.����O����9�D$C�)\����+�c*K��)��DTT��ߛ2����d��D\����J�sH��R��[�V���9�aV�/�,4;��i�4���)��7f��APu���rx�aǚ;q��1���-8������-.D�i	�2�r=@P�]�N=8cp��
̀���D�y��C/NAݪ��r݁�� �#DE���ŃX>�(���j��K�$p�d�>�ׁ�?WXH���ڦ63x�CK	�\]X,�q��$,mk1�����DW��5zrn�����tc�(��O��`s/�=8i�ٯ�>�"�)G�
]�C�
�Z���Ҁ��㍛�� i0ҥȍukXiB%X�}^89���
�X��|�=����y?�����N)%ܼ᱌�ɦY 1�2\�6�+���{���2#/?	ꙹ�B1L��e+`#�=���Ĩn�� AH�B�rٕ'�.���OY�?r��j楄�G1���s�TtF|��Ƀ��D��������y&T١�\����&Tn�8��iRu}���xe6�p�<�B&�,�yJ?Uj�n�7zZ���O�JN���j9O�h+f<O*L:��K�%�"ӭI��9�q��t Jl���2ܘŎ#]���Pi?�M?}[�{�cB�މ
�d�*?����h,����d{���"���Ӻ���)E$���r�I�F�bAJ��қj԰��*�*hG�uk��'�H��ɑ�
 аwiΊ;h@}���Y��L<�P�~J��χ}��Y�y�E��W��ȫ �ȱuu�ha`�V�y�CU��ꃡ@�Z��P'�>(?�`RQ�ˌ~�
��a�"H���;��)��M�Jp�Z�dx�nX��U�g:���K.�M��	�[V��qQቮ��#�.e�H�DlN1o�6���4*��T��������T��,O.�� ν#00� ��"t�ظ��'���9S)r�(@���; �.�X>��~Bp@	�z��}#-��T�p������rQB1��'��0��O�Kr�Qa6K֟JTNpp�^+(�u� 5&3d��Ӻϓnq�W��/1>!3cm�OK�jpJϣ�p?�� P�"?dY�7c�Own@���4i�̍��뭟|���W�H������-���̈/��Y�3k׿y�QiGlE�T+�j��
���>����6DV�H�(ܘ2.f��O��{��p���m�(C�ԓ��>���&цѫ#�<?��4�w�x�m��m ����x�HNKn���/������V
0�q1S��lQ���M�0h
L�$&�!�`�z,��Jg�F!��K&i�8�0>��i�%9�J���}��-��O&X�7�4��?�r�y�w<�bÓ�#�� �� �g� �p
�'s �rF�f(�L��P�aR���+E�s5d��(O� J�B��O�����ʙZ�`XB�n��&Z�I�=����$�;R(LPF{B��	Va�cGQ�!�0��ņ*�~G-C�N���M
żɒ@E�p|h�r�;OܥBQċi�TÏV<N����T�WW*MB�ڶi��@
f+�z�r��a�l�@� 6� �S�D���dʖ��'�0�+��c���N[XZecRӝb>��s5nZ)a�{Μ*hb�����<:���F�Z`̨�"��̡���9[h����U�Wk`��P��#{|�a $�O���I��0� 7N��73�\���d��	2}���<q��r>I��nְk��#�?z�]��
̘se�q&:Q�:�aŪ1^�4�F|r�s�x�K�F���X��F�G�<9�E�<~z��j��Z]R��y����y>D�'g�O��ϓwKx��K�:���h��i:�1+O<GK	�k �)b��,9|)�A�F�0�(
�"�N�`�ˇ2\�j� CC�<)����FX��8 B�\e�G%\ �r�ʮ3�"�2��E6=�20�HH8��pA��7O2� �8�B����-�M{��'���+�-� JjZx�7� ?}x��T 
\���G&H�ߕ� ���e/�>�1�<wTi��iSaz2�A�Th��I^�i����ԉ�]hTHWMX���d!��	?�$t �dG&�M�"$ȧ0����t�x�
)w��X��P[���?�g�Q�;i�$�4$�7T��	��&A���g���0�J�h��4�v̄/q:-�t�*O3����!].GL���#��"U�@ v�1F� 8 ��]F%)V�$">a��#�~�Ah$O����	Fj�ea�)Et�ǉA;y���D�B\�x��+5r�@E��_�(�Ժ���w�$�3"�	l:5sP*�:ʲ�!W�|R鉣���S���
���qC�4�� 10��Z�6�q�A�2�hO����*����M���9�,O�(`�Z�'�� b��!1���ӵf�>	$d�O��'�
�����O�Y�H>���4���x�</[XYZE���<IG���<�i+��Z�O�!�i,��G�eQЩ�y����kH�:t��A��>!�'��<��'vƌ��F�%"Z%B�����٤OD�H��+a�b�%��?�U)·Je��E�� mt8i$!&D��B�L�k�D� R.?$�q����'�$��t�g�I�3�@�������q�s>3� C�	 k6n��ro��x^����	��B�I�|�J-�'�\4}`p��̈P*C�&`�LXJ�`�$	q�)L	/\B�	%-��lӆBJ8n�����_���C�	�Y������t��[�b��dV�C�"o�����58J`�%ͱasXC�I�#C��{�(��X�D��g�&C�Ɏ;�q�*Ǎ=�����r�VB�	5:ѐ0ِ�?�|+�� o��C�I8_7� A�1	�����ro C�	��Z�mY�-dJ�s�N:D�C��L���`�(.x.�Q�C[xz�B�ɐ*L���� !�Eyp�Z� ��B�I�|���D�V��Em&zB��n̠b`��LT)h�nS�k;�B�I�,L��{u���.�,�q��X<B�ɓ�fr�_�GJ��c�'"B��+RaD�"�*-�e���o�C�	TXH����y���Jv�C�ɨ2+�s`(	8h]8(!'��?�C�=��,ffC,J�t��ʗ-[��E*b¡ ��:~��đ+�!��L6&��q���� oxb$!K+�!�ޟclr`ru���>�2�A���9�!�DD������	F�F9��/ŦD�!�D<mѨ [B,�?�T�E��&B�I�5�J��eË�q8� +�ሽx��C�		XP �3�X��d#c��;��C�	�g`($K_#i�v��,^�B	xC�D��kD�_�Y�LM�PHY�G�:C�	!Z"�\�Q�
�iR�ᣀ�ַ]<2C䉐K�Y�W/26�5�֥T&=��C�FUp��Y�݄�Z ��<��B�f�|����\@E��	 �hB�	�1n0`�'&[x��e�,�TX�B�I �޴��B�q��S�$���B��u�zE���z����¤�8V(�B�ia���r0਒3 b�Q�=D�(iC�ֻX*^h���ϣhuj\��<D�<��D�A�͐�@����df8D���͎�\)�Ɗۄw����6a6D��5l�/fj���F��nހlB�� D��(�l�3�@� �fG��Z0� D��	��p�b���`��'Dhj?D��� ǟ
B?���MDq8���C>D��%�X9*��5�C<�f��C;D�8��ǵb*�(gCF"�13f�9D���L&���	0-y��@aǅ%D�� pA����x�0�E���dI,�C"O�@�w��'O��K1W�=왛R"O��p���1ih12�`��f0(�0�"OH�ӣ
8��asC�_�h$Z<��"O��Pr�ɶU�rd��oV�gN]1�"O��:d�-#Ҙ��m�H
 �b�"O D+��@0V��UP���-&
p��"O��i -H#-Z*� �1Dhڔ"O���a��]�lX����2'9���"O �p�C$na`\�̚� /y��"O�)�WD�Ksz�`4f֑w$�%S"O�XQ�Đ$-r١q$H�
�t�t"O��i"R0x�2��LA9�d	"O�ո�W�������d�L���"OD�#��ݯ���Ѳ*/N0=C7"O�$�t�R	)	^%�J�,=����"Oޥq�E�!?^4�D �q/��p"OtP�s���Ir�1�OK�q"�"O^��d��b�Z� �0  1b�"O��P��ĒR6����ɽHBNls�"O\Dö��/_�=� ��e"��a�"OB9
� V�?��͸%&
�̘�#"O<�uiI�g"�ZREX�+�J���"O��Q�b�"}���$�5Z>��Q"O���!�8@�j(�#M��,'���"O¥�Rg�x6���q��+���r�"O�]���
.&J�1 D3.�jB�"O�y���&E&�R1�*s報�"O��*�K���0��E
N�*IJ�"O�i�!b�l��d8�!!Ɍ�2�"O�CЄ��F�.�2���M��"Ol�)B���G����ϓ���mhg"O��3!HN�7��my�.���S�"O�A�Bw��B�i��u&�Q 7"O�I�gM�v�\%R� 3t�6"O�бv"c��lD��88�y�"O�e�B��g����0[� �u"O�e�Ç]�n"$��p���W�~��"OR4K$-G�]Y����+�H�%"O$�Ie�ٔ �ȭ���1X*��"O�dZ��DO:(q����j"O�Q��ϕv�`TjB���Um�Z�"O���!#��W��d�0'F*l6�+u"O��P.J�g#̈��G�<T~<�Q"O��4��"Q4%hu��6M�Q�"ODt�@��#,��:%M�/5���Y�"O`�g-QdQ���aA1�Ak"O@4r7���,aaU�Y�g`V�K�"O���-��Allb��˺z)`�%"O^�[q ǝc�X�97L�ltIۖ"O�\��J�2|�|q�$V�Pp"O^��W����9�%���[1"O"�8�˭]b��¶N�#ۄ�e"O8�p�yG~��b.'qa� ��"O���ԪN=#�a��I�r��@"O�����Z0��a�+�	VǬ�ɷ"O@iHP����ZW��&�@T�6"OJ�b�CRC��|s�e�.*��5h�"O��(�>`��F/i�r��"O�Mb��u��Ţ�C�"3h�M�"O��E�:��P����1���U"O�Q�a���mf4m�0�,��Y�q"O��ir�49�T�b�	>2NZm�u"O��*VB<n:]	�Ɍ�g`1 g"O� �<{�#���*���V1;�Q�"O�	SE�9VNd÷�^z𹰰"O�4��`O�+
�;d��.s"x@%"O(U��o��L��t��C�?�����"O��Zd�Q5G��L�V7d��8�"O��� R(e]&DZ���?R0Ř "O�eZwn�T���H�O�yJęZ�"O�hЗC�)��Q!Ǵ/Dy�G"O$�؁��?U�0q��%�����Id"O�T�D�@��D
7�
(F���iS"O�بЩ�,�v}��-�0\!� b"Or��C�M�jmfg��so���"O��`Ӭ�\6�����8�4�@�"Op���A�6'����[�9|,d/D!�$WU�I�aL�P��i
�Г�!��Xp-�ڙ!x���c�#V!�Bu��H*�a�:d�&$�$T!�@hq���2i� m��^0r<!�'`ꢸR$G�(��EK�c5!��9�^m��o�=�ܥ�-D/G�!�Ē�uJA�C��yaL0 �1O�=�|J�!�=m�B���mӐ!�"�@�<�#��-�Ny�K'\�yӇ�g�<!k
����K�H �qJ��A,Wl�<�S��J�HQ���Y
=�9rt�j�<�!�(aE�ԃ!
͂t�4�I�hg�<I$��
�@���9M%��qff�<1��M/l�^|V�>��j�*V`�<yaH�'h�q8���U �`�<�k^� $��+զ�5<2����GF�<�ֈэov1!s�/�2Aac�QA�<�@�W"�X{��N�!|�as�EFE�<!���3���۱�R����&CE�<��.����Sg��X�"��G�<��רT�>H�n
$�5	U�}�<Ys�T�(E��
�ˈ�^+LtK w�<�b$2��*��� q��;3��|�<� *�.K�袥��i���
w-|�<)�e!z�̍҇;pw*��vƀx�<�ƒ�i�h�D�F�J�JcF�{�<�QJ��Y�P��T7@�����@�<��
=A����E{��TbC��<Ql�u�Ma`��)�K0��C�	j.J���P,}��x���W��C��E��K�k
�BS|UE�ܨ9��B��vԦ��S��7k�Jqk�j�<��B�ɷ^ahWǔ> ��[DÏ24�B��Xm�D��BCrT�7ˌ%H �B�I<\�p�Ō�;�0퉲�]�B䉥-�(;pd_�#d ���lG3�&C�I�Z�L2�擂b>�Q�g �0-,C��Q�d�7.
@��Z�#3@C䉨3����Ðc��I�$M0 C�ɤ`��0�j�$xEr$a¬����B��.9B��`B����!� �%- �B䉘lL�[�9M����h��B|B�k�XzJ�2	�A �')8�B�I�mҺ8bw��*=k <H�O�W�|B�	�s�6|����fY�YP�(G-pB�ɱU��<�UJ��q�ε[wÆ�+i.B��R>�u�C�Y����E��O�C�c)p��V��m�7���^B�IA`~��v*<n��u��.L� >�B�	
fz�GB6��1��׳�B�)� ��VNK��n	0dpx��"O�Y�_�x��`q�(�0P"O���"-���20��K�\|�"OL4��@(5��x��A�i `��"O�P!#��)���#�8�2t�R"OB5:C�*l��aۃ����"O�A��ye�x2B@�%gﮁ�"O� ���~[�t�Nӯ�J$�"OpAj���*�����ܤBu�؃�"O��I�=#�z����^-{����"O<����C� ?|9!�%V��P�"Op��A<i��Z�˓�
@�A "OFur'��	I�(�J�1 v��"O ��C@�q�ŤͲ7dX3�"O���v(6E����*��9@}�&"O@E;d�	�rq�R+ăs �-�!�D��T��]C��i<�!��\�i�!�݁y���*���N JԲ���+{!�d�.��aҪ�,c��ؖ�\�"U!�DP.}��)PG�1��(�)U;F�!���B�<HK7"h􂱩��V)N�!򤗾 �2�V&�4�}��GǨ4�!�ߥ��3�NN�f����<y!�]}�plǫ�	 ��E. !�ĕ��,aq���9}��(��9l�!��
�A�T���,���e˵N]!���=ᶉ+'�"���s�%W�!k!�I:d7�A��\[�Tl��)ĳ<�!�d�#M̜���u��=�Aȟ�f@!�d_�2�"%�dn�! |i%Ѷk8!򤙯g|lkr�!��A��ŎS$!�d�229���ŖN@���ǤV�O�!�	�B�j/�{��)�d��]�!����
��%+��R�2���#�!�$�!aJ;���2{�8�GA�"2�!�$��ZP;r
ޖ:��;�`�U�!򤟾C���ce�<�4R�@�<o�!�D��0�%ř$��UG-Kx�!��$!ݬ=:&�$��\ p.�7$�!�DF�}��@�ܱG�6�Bp��1 �!��G���.
�A���!WA�)w!�$�9o̐-L@Ĳ�I���A"O(��dMD�]��;$��H�"OLp�EN�qj�����0F_�9�a"O��A���3�n=�gb�$t꺔$"O,!�������	ԣ)S��X;s"O�����{ֲ}b��W�a�x�D"O��Nt�,e�&`Q�Y2��R"O@��
y�%+��ƊC^|yd"OjM���|t���ȘR\S&"O��E�J�d���I-;q��"O�|;�m��ʐ���ϙd-����"OH��F#��b���[Bt�x�<1��ߐ'�&,���i��a3�S^�<CG� q�؀��P�NkN�P��~�<�����EP�ș�"&���#[z�<C��V̕B���s��Ȋ@�A�<y�M��7�i
��14����N�y�<!�E��L~�FF�-4l0@�h�s�<��\�\����Dִ��]�s�<����:x����$IV.`6��C��g�<���^*D����GP�}�N�e�<a�,ȟ=Č�DhكA�b��a�<��@��|�-�VɄ=`�PRrK@V�<� n�91ƀ+bk�nP	Hvn8"OZAR�� I�5s�Ps\ #d"O���KZ**� ��׎��[Y=�B"OVD{b�(]��p��/^O�hHg"O�1�󧞣FT\�X�%֙I*­��"O�dQ'nݲA0^P����]�V(��"O���P㔲���i�aD���D"O�$�v�D;X��A����h+P��"O,���JF�I!��B�N��O&�a"O��Yrj��ȁ �O��c�f�zS"O�1�o�&a�3�EW?G?p��2"Ojh�WJԭ�!�JS�n3�R�"OP���*�UJ��B�P"O ب�����iG
\� ��
0"OP�3� �|9w؈�ܨD"Ot���S�F�<C5��� �p5"O~,��M�v����-j5DB�"O�|࡮�#PJ���nŌ��Yb"O��"I�\$���wj� 6"O"��+�)K�R9{p� ~�,�� "O ���(vh4���o�&͚"O��5"Q�\a�B�h�ɥ"O4L�t��:gꥫ�,HI0zW"Of�y��R*��(��n���yC"OX���fx��@�P�;*) �"OD `r�C�o�B�H�Ɗ? �]�%"O���&�'j�@���$%w�l!��"O`����:/��H��4.�^%Ҧ"On�y���!&�j��o�ki,�R"O����R�3��!�N�8*D�0"O��KR������pe,�P� �"O$����+͈d;� "�}�"O(h���ZD�s�ϓC�j�j�"OR#b�_�j����˟<����"O�X��Ș�׀l�A�̰ED�ѐ"OtL�a�-���K���]���"O6ŉE�C1���x���c�V5r�"O�1 FA�QQvm�����lI���'p���5 6��?m�,�K��2K�Dy��'	������ �8�K�ޞYg,��'v��R���Vd�
Q�ܴ[��8A�'pL$��:�R�p��Zz����2��|��4qM,�So�S_��MW�5_D���O~���G��$�-�Vd499֙&���?Q��ɋ/@mi�A��(I:�GA�!�D�<��,a���`���蕎A4��5�£<�j��N{4�(¤'
�S]F�s���Xh<�� �rBh�Ƈ݆f풤�"��y"� &�Օ^�� u���y�^�ܐe��,E?*�a1D��y��R|����!CX#@�t!�`��"�y*^-)xU�$�Q�g�0�`�W�y2d7�ju�܂0��j�fݜ�yB�Q�M�1w�.�w
L1�(O4��'p�-�⫑���5��'��x����ȓ�$�����"<�ܺ���2���ȓ��S��C�>n4���V?�����O�6E#�G&����AW��U�ȓtR����!^d&��2 ��H��ȓ}�P�0� �9!� )���ڴb�Q���ո ��=Fp�����soH��:�X5���߶c��� ����X¼��'�ХHt&T[+�|H�B�,�y��s���3CȾ5��rp�uVn��S�? *��c�G����}��;4"O�pX͊3v:��PQ��y����5"O��0$�W6a-�9{э�>fr�I�4"O�ls��H3N�SFL��Q��x��0�!��1h��4��*{$L�ȓu4��K���V'ґ��%Q�xD��/���7��.��v��x%@U����m�Ɗ����[䠕q���ȓ S�Q!�DYP����5��-�ȓ ����U��E�*иG��?�}�ȓd���j�[,%ȴ0g���@����ȓ���C6
δFg�	d��E�e��.Ĵc �sW��tBۿ(���ȓ
y�� !�"�N�xEǑ?� 4����$���W.,��h���q�F{"�O0*�\!!� #a�^�'�B�	�'@@���$
F� �"�+/��l��'���pWR�O��<���R��̡�'}���! ęX��h�'��O`
4�'߲y-4X8i��sk�4׊�HO�=�OA��a%V�6��Ȗ̳Ch��@�'�a�i�=9~�*&C0iϊ�C#F�y����Ȁ	 �ЉNR��1+��y"�	�$H�8���F�l�k"���y��ČX:p�5�Y\lPB���>!B�DG}��9pzc��� ��U��y��$�>�}�'#,u�F.V�}����.Y<f�t�A�bY��F�T���M|��
S�9o^>�H�Ϟ�y��ҡc%~hx��F%o�B	�M�'��d/�S�O�����g�5���'�M"���R�'�B�	�>]�`$i.%nȠ��'���e�	5���З �|y�'�J�QD)0S�PQwhG��Tk�'�1pr�N/W�j�G�0���'�N���H��.�|,'��H�P�'�:�Pᜲ��I��
���D��'"��C��F�J�5�E�w����'���R$H�i��pI}�,���'���"?e�,���6W��	�'�%C��X;M�D�G6�C�'��J8F��WmH���E>w:C�	�,8v��u��.�h�Q5qg�B�I�a<x|��#�
w$y�5QL9�B�I��&���F�:,�	�E� |YzB䉪uH�`����
��=��䛘�@��hO>	��B��C�ȭ)��7:�R��.�Ox�O4x���9R�"�+@�o�x���"OT|8S#W�5�u3w�H6[w�i�"O��J��
�~���\t��"O�hPjM�I��Pg^�.< ��s"O(�����?+b���k�
B��H#"O
��F��i�z�B�+ɴAD�� _�<���=]��xA����-�X}rՉ�6+��C�&�)B��6l�1�&M�C�I��5S�o��`�V:�k�Eo�B�	 �^=3�iF�2G8Z�A0T��B�?O�P���؅.����am�C�PC䉗8h�	�&D�)�'��.C�	�[���l�]~=���nO�B�I.����1�0rBI�4b�*�B�&l.��q�La>>i�PmB�nF"��p?Ѵ�Pe��Q���P*�v�3VCPC<)���Ra��k3��%��)����ȓ��qP��4��eM�<m���S�? 8��g�P;'.:�i��*	�H(s�"O@Aٰ�Oh��b���ijF��O0⟀F�U+l�z�"�!ٙDκ��U��yRj�;F�Dس�X�8|��B➚�y��'�Ա��+VT�j���b��;�S�4l�/���G�S(���0d�I@�<�!N�*�Fi�1��+m��4C3��c�<A�$X�^���r���\% IDH�<i�C��r,�DБ��fޭ:�@�<I���S�v�<�z�N'Jj� ��ʎi��ġ�ؓ�!N���#�
G�,a��.}��'Z�d�ƮU��=Y�#И$B8��
Ó�hO�KP��.�����M�Qn�ZA"O<��4+]<V>�� �ES��	a��h�
"<�Os�M��G��}��nI�!����W��yRHT�5�VyK�č:�d�5�Ģ�y��	Y��0xTN���ѡpdH��yb$R�v��Prp�R� ��p��1�y�ꞃC����M�sI^�S�.�y"�T�J:�I��$t�0�*D�"�y�F߈a��5 ����a·6�y���l�PU W'i�]@,�0�y��N��:��/��5I��:&L��y"��>w��IWOΥ4�2	bhS(�yҋ�6+��%
g�ɡ0@�����y�
�
O�)�.s�D�d��yb��N��a,,.$��$����yG���8D9UF�',�Äޠ�y���&����H�@E��I��ynip��N�.9�L�
f�؅�z%h����7&�)���M�-�ȓ>dfi��kҁQ�
Q鑃�q%�L��#.��t�9j�h�����̄ȓSݎ!�c�|�FE��GX�zrX��ȓ:<��b��>d�8����T��z̄ȓzM�4��ͺyc\8I'�3x�u�ȓ-�^M��םS��P�un=����'���C2eLv��,�4��p��w�x�����T�k��C����9����3fQ�V�(�
#N�G2���k =qU��)DF�B�bB�Ʉ�_:��@���"�H�n�Ԉ�ȓz��Q "�\��(�S��X��RQ�`B"Q�D���aF�]����D��t���D� 0�M�`�4'>2H��u�����[�U�I�	�F��ȓ|xb��M�j3�<�a��+�8�ȓ���S�#=gO��cN.��ȓ\ȽB���iT6�x�/Z5����P�
G�՝݆�� O�,4ه�G�H������G˼��񢜗oo��ȓk|L��cC2������g"~���XY`�����+o&���(�$?_���ȓ7_���-\ �Ơ��N1BL��:$A���	��yЧ-Z$f~�ЄȓGy����V{����h�X��ׂx����ֈ�r����(�y��C�b&R!	æJ/k�	��$A��y�B�)g��`E����t8�����ybM�[=��X�̞�<�!���y�	^:������lђ�#�/��ym�?/
�s�BB,Xp�Q��6�y��V� <�@	�nح,���'OU��y2cJ�@����n֔qZ��f�
�y
� Y��Լ]�&���)�p���"Oڷi��5	��ޱ>d���P"O`��K =R���u��1aY��{ "O�����,r���r�^3l9�I1�"O�p�����w�)����Y�:���"O(�Y��S# s ���݉��`��"OvU�a��P�D���,���X�x�"O�����5w���"櫖6[���p�"O%cr���H���+$/�, �"O�DG��dm�!�ڲj�X�r�"O< PuoX�t��s�	Ľ8��]�V"Oȱ���̤`���`B�&`�
�j�"O����U'?0ҭ�,��n�*�[c"O8�����G)�=��j�y���0"O�x�0Ő����q�k
J��j�"O�m��HJ�ޔ���՚�ر"O��`��q��0{3�֢W+bm(q"O~� ��g��ّ���� ��"O���5M%P%|��g��%;����"O�0����Ld^y��˂�/en�*�"O�� t\.Fu�q+�jٺ6H��"O�Up2FИ�@����z�"Oz�T挭���(U;)�ڭj�"O�aKW�N�5�(U���#R���"O
}22��;R#�Aw�J!�	@�"O�$C��=
L��rB��S"O`J �ƴ!)�w��P��AKA"O��K�튗?pE����/Q�L(B�"O$�$!�{Rtq��0�:�е"O~�iV���+24ِb��f��l v"O4���-؈u���f�5���0P"O�IPm��GȐ4�!�97jZR�"O:̠&٪Qb8ٻ�o��)XJ��"Oҙ�'=(X����8�"Њ�"O���&��&*if�r#�=$t�2�"O�k$
ΈQ�0<�#�"V#�Å"O,�PKӶ|B��i0��|�E2�"O6l⠀�R8r9`���* �Jճ!"OhE2���(��$8R��T�'"OR�ِeF�J.�e�3nO�<��2$"O����MF�:��D��mƥU�^4�4"OV�#N�2�,L�(l-��"O.|��,T�}i�hȡH!��t�"OP(s3��n=؀�W��.'�ʌ�D"O()S!�t2h �5����G"O4�,�
m�=�T��	_,hB"On<j��L�da2-BSĆ�g6Fp4"O.��!-Z(K����"j�d�@�"O8`�e8����G�d���`t"ON!9�����\���ݎQ⒡�1"O�sTk�57�QZA�t1�aۢ"O<)H�O��s`c�K�<��"O�lKt�� �t�9��އ(�Z�iA"O���F :~�3����w�X�a�"OЭ��X�Q�0�8p4P��V"OZdcaK�AZ�qD	�:Z}j]��"O���K���у�߻m6�"O�Xk�.�(#*Ȁ�EcP���I!�"O��9���5�^�@[�u�Ez1"Oh��%�b��6���3�B��"O>�#�� e�@|���I�(T�a4"O��5"�)<@���;-J3"O0���L�?3ւ��_����bۙk�!򄁡S��A��!�;+�@�$��3�!�� ,,b5�=u�f]�۝ 뎸��"OP���n)=Dћ�!D��:�b�"O��w,�@j ��P�D	�'"On�(�π?z�H��K�B����"O�hR�"|�4�F�^$:����"OLQ��g��;Ir�'�R�b���"OJ5qQjD�sHRu��(+y�5HS"Od�$�O��Mh`��~k�a�"O��8�������k��r"O�E!��,da�����eG2%""OFX C�m�Z�ˡ�:5*Ż�"O�Ev[-�$���z�J0"O�0KP�6t���w��'f���c"O�UYuI@��u �i�1U��)�Q"O��	�D�ƨ��H��A���4"O����"k�"؁�ͳ��"O\y�!G�3S�ԕ���mR"Œ&"Od�[Qf��BAL%:�������!���a��m���9!}�q�"V� ]!��(in���EY35k6I5b��zW!��8>����ቂ0Y$y�s�U8!�D_���G(V(W�y�s�@�!�� ��䫵��"Y��S�[�$�!�H�D��u��w66ܙU���!�$�N����ī�1z��שGy!�Ӏ)h�hu.DV�"-1�F�_!��a5@�Qp�Q'6�.�ˤ��/1&!�	'z�	8Ӫ'�F<[0i��C!���5TT*Ă�C�;�hE2�պ7�!�D��x�F�2��]�FDʱ���
!��S�7�r-܇)a�����_�!�	#?p�����2ppr,�=�!��C�W\IZ�O՜*��#V�ˤq?!��_.���M_&9�X@���/!���+s��k�)]%'tbI�cJ$h�!����ܓ�(\<_��
f/א�!�D�?�ey�����3�횺#�!�^�2���a�-Q�5�V�y��%cb!�$
O���z�h�O���խ*NO!��AfѰ�H �J���}����j/!�DW�t����c#�"� ��k²'!�H9AČ��A�g=$�闋@!�DK8}:����#3�p㑇��!�d�&�D����4V�m��OB;a!�]�ya3�Ρ.[�z��
�zf!�Đ�$�Q��L�nV��pbN30J!����w|ش�F���'7N��mE9!��7��`��ö<b4�'mH�!�$ڕ+�5�6�?�č�flْ�!�\_�n0�dfҞy�<��",�Y!��&\mఙ
�G�+�^'$(�	�': )���-��P��o^�Z1�U#	�'�+��
Y�x���6Qjp�� �&D���,U����Q4Jt(b�"!D�� 7Dי��,��N�arX�A?D��Ԁ�,,b��d�Ɋn`|I��f0D�d�A�ʘ(P��r�kƊK	���Da.D��HU��D������`t�4k,D��S�Tb���"���g��B�.X�|4��
>��4A��Q�!��B��5e�(�� K�C��L�!ϔ�q�B��DQ8�"Dտ=�������=|B�I�<�2����"F%�	���Q�zB�C�5�Rl�@Cˈ��!��Lј7zC�)� f�hF��E�v�(��6~���i"OTA	b��9�c3U�@"(1�"O�h��Ŭl�Zd1#�޽s}���"O\���H&I:�	Y�uq3�"O�m��GI��x0��;�Z11�"OD�3GK�u����%�H��"Op���`����ɥ�Y<r�j��"O���Ä�2F�x��v�pp�"O������`3���I[F�W"OZ	���*�f�q�\%Uc�
@"O��i��� ���V� ."XDI�e"O�	��b��N�B�^�#��aA"OD첰@����ѵoB����"O���	:S�|9J�!D�
�r�"O��G���p��aT"j&�,��"O@�z�-Q
n���Ǧ�d�� "O&������<hph?pyd�i�"O~E���P4U%��Ѡ@߷fe\��"O(!�
S�V�l=d��|����"O��k�?����d��jt�Q�"O�)B�K�%&lت�����"O�"pA�xO��i��W9Cx��"O�Q�D��l!�e��ʿ>x)H#"O2���X�h����-�80¹ �"O��#�A�'��Y�.V�Q-d]X0"O4d�� �;j0�0unO�"I��P"O�����^pj�q+�M�\&���w"O8a��1�0��Wj�'D��j�"O
1�.:
�,�(R{Q�v&�J�<��ƶjrpy���Q$/��؇c�J�<'��(YN�-p�$��%9��jt��M�<���Vn6Ȩɴ�ƖM�6D�Lr�<At.G��j%��a��u�p���l�<��耩�'Z�>����~�<�eK��jL�H�Y�<h#�K|�<�����%�%�D������y�<AьT/A�w]��M�b�L$��"O,4�����̐7�s*f�k�"O�]R"�P�C�����*�|[U"O��D�TrlA��n�#a�v��"Or��"Ɏ�b���a�L�gs�1��"OĩI�(}���s�Ѹe�PS�"OZ��Ǆ��8�
��V�R����b"O���v�v��r����&M�"Ojກ��&M�.��-���R�"O����]b��D�� �%4 6!�"O �H�C~�Z�@� �:d;"O4���Ӣg�6���5t���"O����S�p��D�e ��O%d���"O�8��״E��c&\=�8̣"O\$;���Q׀17���a�6�I�"O ݪP�3X�X]��d���Y�b"O>�3,S�҄�0C��<	"O���`���58&} `cM�g+\���"O��Y��FO�z _�T�a"ORe���1}i�Kק�q|�� "Oꄢ1 � a(EAd��-��"O�, ��m/1S��@^��"OB�֦@,dt0y�؛.��8�"O��j��b������_���Т"Oe�ή(tF�b�'B�6uX@3�"O�|h�*�@54r�f�'Qpz5`q"OX�؆nQV ��W��EZ�0�C"O�(��CU�#��@aA��;F"O� p�0����ȫ �*I_���"OL˗	۱DZ�e�6l(V?~��7"O���'�{<����n��5��"O$�)4�ۡ.��T�0Қ�"O����4D��;�C�R^���#"O��hF�1�bա���+xf0���"O�AY���4,�,ZS��r_D� w"O��I��Z��|1��'eV��"O�i�.�>"��X�W/Q�p:d�b"Oޕ���P�4��`SI�J���"OL�3pŝ<KO�yr���4Ozk!"O,�8�eR1+^��BIڞDy�5�T"O<l+���-7�f��Rȁ�b���"O�%����08�WF� xQ�I#g"OR)rSd�QB>IB�EV�!C��v"O\�K���iJA��e?d%D(2"Ol�:��4e��Y���Ĭ���"O$}��F�Z,�q�%|Ӑ��"O��9f͇���q����m�]H�"O��
�$��QTF��sKX�:��*�"OT�Cs+O+Q�4p	q�ABN`�q�"O�Dk�-B�s�@��vhF+=8��"O��Ӏ�7px��GL*�\"O0$30��	x����w�b��"OJy��o;,Ȃ���9v�,���"O�4q�'��`�kw��6�v�9F"O��8թ0M�d��b��N����"O$슄e��I����6*�<�Z�"OR���/C&Th�`R s�v���"OZD��eݛQ�Vt����>�3w"Od��%��A�\��)�8�P"O�y�s��i��ˎqX����"O�`B��5yT�{bJгE���"O��XQ#�	�Rx�I4rR��sB"Ox���ˊ%�l�&�J.`��\�U"Obx�
3Y�(!�@Е�@���"O }J���<H�r�"�����M7"O��IdI���H��1�(���"O\Ǫ�T���J�U�@`�!"O�Pb@� �X]hSWG �Q8��Y"O 	��]�rn=�5�@�l*"OؕA���h���^�Hk��7�yb���xfZ�f����+`���y��G�>Lk�%ͧL!H�g���yb��i\�#Ņ�Qb*iV��+�y"%�(pP�q��)�~��qՈ*�y�IH2S����f\{�̱k�)��yR�R�P��d�Nyx���yB�W"J% ��6_~�h�&���y�F��.���AԨK����%�y�"�6 �.��l��@�F&E!�yLM�(v���dA���q&˄��y"(�0G�1��܈g��0��.�y�M�pbn�4�کE��� ��5�y�-@�("�P1ě*?	�K��y�̝'Ԡ�cֈ3c�kp��y�(��s�*<�C ֜0�$ǧO��yΕ	���H��6�P�{��X��y�I-���2��35X|J�lY��yBg�Z��}��-fb������yr���a+�<�0tz�����y�,M*k�8�1gO,�"1�å�?�y���3�@\"�m�%
�����yr�%t� D��,��!��i�r �8�y
� ,Y"��%�( ��tR&�2b"OJ1���w���� E4(���"OTl!�ȋcy����Iؼ�fp� "Oz�C�f�?Ό��5��V�6�"O8{r͋!?�j���D7��<P"O�%��-�$]Ŝ�:�g�j��1�@"Oʍ�L� Ç�&�:)H "O��WK��9jD�p�ҥs�0�X�"O�M�K<�F�PB#�=#x�R3"Ol��C���P9s�C S8j�C"O��1Ã!c�8Ib��9̀h�Q"O %�v�H5���Ɓ޳��%k"O8!�#d��I#6�)BFX>�:(�"OL$Ӣ
�_�F�
�$&}X�P��"O�H�w�L��r��R )F��)�"O�h	+κ!H���ӭ�"�z�"OB0NX�x ��`�ěf���XU"O����b¨�J���IL�<��AW9'De�b�TQ��`���I�<A���=�8fL4RX��E�<��8mH�ӒHߙLz\)��D�<����-���;�#��X)��Rb�}�<IBO�9�F�ニ�;l�T���
�{�<���B-Rh�	��
;�-����x�<!'�S-����WH��	�H�i�$~�<���e�<,)F�V�xT	�/_y�<�r쐳vT�M�1�pi��x�<AD,G�T�0v�U�)��:1f�^�<��-( GD��#A�-A( �1�@�<I��0Z�,��㇗t��1e}�<����b�*���J��ie�_�<��RQ���02iۋjX8���Y_�<10�;\����0�݇X �dYrl�q�<A�dJ�eW����  ?b�D�9�jQn�<���p� ��cP%pṞ���s�<)�_��M�l���n�<)f�](:�X��NM�b��tIj�<vhó0t *]�t��$�b�<�C$��=|P�k�BO�S!��1[�<9Ge��,B��`�C�[t�``���U�<ْ��<z� ����$|B��a��N�<I���&S]��6.��v��
�-�J�<Yu�Z�la�Ս�h784�Ak�<1��;4�`�T�m�'}�<��\�b��'������v�<��D��%�n5����)[���b'r�<��ωR"�{���(����fE�<9�V�B�Ib�[���	�DU�<�f���&�,PB�߳.Z�!�D{�<��S�M�>������
��<(�A�u�<IU[�o��3A$޶ r���U^o�<Y���ɂ�ِr�����$S�y�c�:'P�`G`�n��i�O��y�%�Y���B��d������1�y����p�mqvJZOP(xq
��y"�  t�i{� К&�������y��&j��l��؁!�X��� �y���� X�3�(��%�E�D��!��h�Y���G4fҝ���t�^�ȓ:�テ�V���A��(Qj��� )H��`hƜ��*�)k�d��ʂ ��MKN
� �W�Zt�ȓ9��X`��2%��B@_������I�pbŊ� }:-��ˏ�`����S�? P,����"0��eO�d��A� "O�<`��ҽ	�H�K­��z��Ӷ"O�M��&Ěl�&���=u@. ��"OxL"CK�i.+��+.�0��Sv�<�T T�p���,dVP���u����F�d�G)��oOĠ#��+a�%�ȓU�4\h5 ލ;��x�A��t�y�ȓ|~��x@D�[�@��B�7�\%�ȓ 0�1�vɢdxH���!5歇�{���z�@�{J��!�%G�2q�ȓ{^I��bE�/6N�����i]zІȓK�R�:0�جH��e�
Og؆�ȓ!C�L(r��_�&����[�	:� ��J>b�ۣJL�2�$I�A�(w����A�n�!W�
��Q�ğ�
�f�ȓ^�D�AK#Z�T����w&���Zu��:rd@�%��,yg�.uD����H��/~�l@�v�]+$��ȓv����L?����N�P,�Ȅ�,������{ݔ���	��i�ȓzm�m�Ň@�L�m2�J�(iLب�ȓ(�q��g�S��Ļ�蔧C�����$��=� ��!+ĥ3�̡_�J0��:������ߨw�p���ZŜ���uG������U���8 Ϛ+�ȓ_��(ǁ� `����u���`hY�ȓAn�lD��Nkĵ�ԁC�U����Xj��"<�,]9V�ń}�V��ȓ
�^����֓;bb13�ܾN�Ȍ��'Q�rH���� űBW�-�ȓ ��%A��� ��7�H39����	Y�'�|MBU@K�n������k��z�'�jq91 �;Lr�غԠ�+R� �@�'|�pE���	6ܪՏA�M`���'"��y�N�)�*D���PAw� ��'Ħ*�%�"p��SI�%�B|		�'�y[�'X
���3M�*�P�'P�ZB�8Z��9 ��v�b��'舕��N�%�j�0���p� d��'�d��v��gV�{�H�e*,�#�'�P0S�o�4 �hc0�Ӫa�&4�'�V��2,t�|Y�G%%��C�'���0$���k�:�@���Tn����'��3s�Ȧ+� �*RشM��'uʭ0P͜r�HD{�J�>��
�'�z�a�
�})��A'���sW�	S�'�B�'��up��D�0=��Se��$
��'m�k��C@�ǋ�{m^���'�5�TBќy���Fy9@���'&� �gH�n�t��V��-�I��r�E��������5Vƒ���S����c��!eJ`݊ e�m���1݀��� ՓF�t�AnH�(܄�4�d���(�m�1��H��5Jbلȓ0�Q��-I��I���� dlنȓ]��CV�:Q�%;�@�(4�U�ȓ1*�Ñ� <7>i�"��U�2�ȓe����En�I��lKV�V,.�Ԇ�E� � uE��*Ƅ-�Ճ�A-6%�ȓ"�a�`�^�t,�5�m7�A���]�Bn	����8�A=wajM��SF��*w��;d<�e� m���ȓ�.F�`;#���)�,L��"l�<����X��k�ń����h�S�<� ��B�\7{"^L C&��/®tp"OA���O>�d��EN�H�T5��"O��&D�v�a��F��2�x��P�d$�S�',�h�k��ʚ�����nZ���,��6>0P��/^��q��(&x44�ȓ@�&������Jh* �"�� T�4��ȓ7���$�v>�����ԙ,�)��:�X3��~/��p�)ݩ v��� S�h��d�Y�D�*V-T�цȓdS� ���8(d�
҉�}Rҁ�<	�����?y��QCQE��t��G
L�!�YU<��ZG��>����!��!�	q����L�l⼬Ke�.Le!򤅹>���a��50�V�z0�ͦX�!��Ʈ45�M��/��l�Ɯ����-!򤀐e��만¿²�p��_>;!�M�B*�l"sl�����!*��!�D_�!���1�UY�<�j�{!�d��f���ĤQ�$Tq�D�m�!�5�lyP4 �3�` �צAb�!�dN�7���.a�h=HS �^W!�d6-�ji2�ͰU\J%��/MW!�T!��|�D�TiJ���%O!�$� 5,�`v>�y��!�D�@��CAW�.%�,�`!��!�D��;�f�:����_�Ċ��S�!��7J �8��.L�rI��L�)@!�D^�&���s�3s�&9hӭY
9!�dJ��	*���H��|��l��U"!򄚃k�B=z���i��X���Z.o�!�dI�{؄�H�ˉ�>���Q��F�J�!���P�ҩ��g�(X���O�!�dO�1�ͫO��B!��⣬Ӻ�PyR��!Ȩ���[';���L��y"	R\���pg�l���w�_��y2/շ*1�qĄ˹g�F%�wH��y�O��+(����ɕ%`�t�w�Z?�y�*_
0���Y��S[���R��y҅ϳh��R��8K|xA�gS�yB���~�8�"��կV3TA�aٱ�y��L�aR�ZS.�%���\�y�N�o��ApA�^w��p�〜��yr�݇%&ܰd�!nφ���Ϡ�y�j�}��t���ֶg�}됤\�y�����D5bA�y0a�u�Z��y��גU�����:tz0�C��y�DW"VH{b���^�s#�G��y� '/,�`Ћ��C����n���y�`�z���4���>��-:����y#�:�<���;4��"�
�y2�A#̑�t@F�ػ��ů�y2� �<i�Yj��0�֔�y�A��zYL�h697.$h	#$��yRi�D��94�׼&'� :���y2��XTVh��Nŉu�t����yRm̵H��86Aб���Q�H�3�y��|CڝHP��AC<���"�y��'X��,9�I�&8�3����y�� ,����������P:��'��{R�ڤ~�(����*��
 �yRjf�J ��C5zCJx���\��y�f�_?^	Ѧ�ؠo�Jmk!D��y��W2JY���j��=��ܽ�yj�a����f�\AY�T�y
� ,	������c��U��x�B"O���KW�s�v����$l�tE
�"OR �AE��v��0/^�R��@�"O��"G�\f���!ň<L�^��"OLM`�K�7d{L�Ѕ�OYD�"O��:b��&JW谲���c9<�I�"O2��6
D�y�α0�-�4.�5�%"O:p�Ȁ&h�P��[%�L�"O r�É+ZA���aTxe(�4O4�=E��A*ZG���O�����'�Z,�y2��zjp ���ũ�his�L�yb��
I�Ĺ �L�6s��Q@
�4�y"/�u|X!��gāy��P���2�y2i�-3 �H�$l~e�wiѓ�y2��"e!0e�d�6G�`�p��J��yn�r��}@�+6P�"9��^��	z�)��<Q%ǘy�j��gA�u��'iƪ�hO?��x�5ҳ�K����PI�56�C�I�W1\�R�U�I_�}�g�=z�
C�&�L���+/־M(AD�j��B�IX�:1$�яZ̘ݚ,S�b��C䉗A�ؽ�L��UJ�p��.�C�	E�`A��O��F�JػQ�Ι2��C�	[2�I�EI�|��t@�N^�C䉌��=�#���by�
�qZlC�	�#��<�����s.�����mC��
y��m�����ޮ��B�	a��QE#Kn��Q�,�nB�I�VĊ};s��w�eJ��9��C�I/ *��!�̏oF��b�pC��L��}Xc�Z�4����3�̉^iC�ɲ0��l����(c�4�j��L�+3�B� a9�L�� 	Z$X��f�,P|�B�03���)ID�8�hf� �K��B��#C6��e�8\Z4]����2�vB��-q�SD�/h	�a@�F�C�	�2�D+&nNKTai5m�:z�B�I�_|A��A��iആ���B�	3.�X�AA�W:C֮d�G��q�B�I�|��e��$:���ق��0f�B䉰E��p֥��n�BTy���nz�B� oʤ"%hT�v(��h �|B�ɕW^9�p�H&r�F���+
�n�bB�I.H�j�p�ɐL�&L�*�i6B��!e�:1��iK�B�D��F^�C�I� ��%2D��:*|��D7J��C�ɬ/ΐaåOn�P�NM�;�B�I�c�����0\e�3�(Y�tB�0�j�A��@�U�a� rdB�ɷE�Ziʶ��z䖥{C#C<12XB�	.�J�R�l��q;�b֠f"DB�I�e��1����&�N���(P�X��C�I��\Z4�q�D���N
�\C�	���)xB
0j*uRv
��iHC�	��`�M�P��S/��J"C䉣{~�}ґ.$�h���p<C�I�r�"!�&�V���""���;lC�	;�,�M�4I���r'���B�Q�u�"��3d�f��jҐ*>�B�I�;1������%fG��s���z�C�I/uF���f�79,�M)��!MlB��&��f��YWb�*�+ �D�.B� '�Z��H�M$
��d�X�p�B��[��8[���1{=�9�3d�0z(C�)� r-�B�G,I Q�NH�W��*"O6�vm�/UTlaH Ċ{�>�!"O.0¤��Iq�8�U��#^����'"O�p:L�x`��I���jE�<��k�&]\qկ�()K<-c��|�<�tB�7d��p�BK3�V��Zm�<�`�
�n]�� A�ݘ�oU�<�eD��Č�;&8pepD�{�<i#(�=u������<L��f,�w�<��l@�X6z��PD��r)�hZ���t�<SMN;r��;��1X�|��.h�<i��A[ִYBR�@$-(X�(�_�<	�?P\h��Q�tf�QA��a�<���*X��cN�k�P��0H�_�<�T�Ե2GϚ�~z��x'�G[�<Y�L��!d��6��E�}�ҁ�r�<a�݋$ɰdr$P�Q�<|�~���D���ʆ�$]��`GJ�U5����'�:+��Ҡp�$�X��6:Z�ȓ)6�y���Ze봱hbD�49��l�ȓ\�m���-oy��p'�*-&2t��7~,�)a�1p��*	�+~���k������7 .H# �ߣ)\x�ȓ�&�0�#ϧ�������4P=��ȓv�|H��ՅM$�5�,۔�n@��E�N��QM��K¥�ҊWs�$H�ȓm&����!� 8�I�۫D�z�\��Fe̥
i5��O'�����H3����{
)QB�"��Ї��ĩڔ��diN�1 �
7j:�|��]��H����4F<� K��/K��ȓ��u9�Gn~	���2��`��_3H�B�J�9N�#F�,Z�:�ȓ����
��Z*d�{�N'<Y���ȓWQ�\؀.S��4�k��%<��ȓ)���i��6�����]�q�����/��� ���-]Ǝ�(uK�q���ȓ8t ���e�(	5��BC�CP>���T�d���gF�$��"n�{a܄��0 ʇ�Ï&�ĝ����4-x���xo^��� �VQ�%��
7!����\t؍E��[ �XvIҋ����z�b�	��!��p���-[��̄�#O��5�ʹ Y��P�_�p����@������I��XȦ�C<p݅ȓ�B
�[�L"�TH���-��Cخ|�WډN��`��
���ȓK��3`�g��C�j�����q�f�$�ܒ�,�so�Q#l0D�D��n�=oFR��o`�7H.D��
3��&U�l���)CbTi��-D�|�Gꃂa2"���+ϕ��y��-D�|��-H#��;p$L�࠭�� D�<�,-h�f���͋������$1D��[aC�ll��`FK��~�P �-D�����K�Z7���,H�6p��۠&D����/��@$�"%�E�!ϲɢ�#D���=M����,��Q�~I+ !D�PA��M4{��h�L��V�p��=D�L��Cy֪А��U�N��0)D��z�a�6U�j��V��{6��'D�L�VFǒ5��,��(�!ye��$D� 5m�2)Ǡ���:s2�D��<D����Ԅ[�"-�E��<L���9D�� L�U�T�f�a�j� r�,��"O�l1U
��R�U�Ŋ�Cd�`�"O���,�<�V��HW�c~\bC"O� ���4W��Ht����q� "Oe��a	w�J���f�@m
�a�"O���
�<+��`2K�(	c�Ⱥ�"O6\P��ʕZ�|�J@�W9��$"O�;�Il��+u�N�(%TDa5�<D�̡�Eܼ(������0m�&d��8D����DF[q�܈5�	\�Vy�+D�P���ɳv����ʇ\X�ÓO$D��8�o�1Mώճm�&'�Lqaug D�����˾*T �P��J�3�	 #D��sod�ҵ@�!|���D"D�`���Q�����[�w�Έ���%D�$SeҾ%�9ʐd�)9p���i D�x`%N�Y杂e-s�MP�"!D���ƚ+1�g�TٞXcխ>D����oR�&H�����$Ɋ�x�J=D���U�R|%�J���d���:D�T)iX.�}�`�\���m0��5D��Aǂ�j\p���V�Ɍ�Pd3D��1���֙
Ɔ�&V�� $D�|���]*�f]j7_��r1�t�!D��Qr䝞7a �-Ȯ�6�6>D��j3��=�$���ӑ<�Z�Ȳ�9D��+�A-4.��ԗ.�^Y�L9D�tzT&�9I�pe{��YoDP���7D����B�$���*��.V,�p�6D� ��dÆ;�-c�Nn�!��8D��KP��@����4��2�u�A6D��Y��dn@ &G�/d\���4D�8 �"{+x��i�'q�i2��4D��"4@�6{�x��&\R���2D��cɐa3���� 8o�M��b<D�8q�@�d�(�d">㬱jq�8D��;R�4#*Z���/ҫ�j���6D�@�6/H-;'`c�(!�'2D��T��Ҁl G⏪Y�dj�C��I�&�Q��Π'"�d��Q�L0C�	�B\au@Ɨ|��)a��5��B�I)=rn#�l����O�1[�B��
X��DIV�P��� dӏL�nB��E|mie莸=���rt���:B�I,ҔYI5ʿ3���f@#)rB�=Qz��Sb�ŋ=�	3rn^(��B�ɀ<oر��J>x2�xq�C�B�I�v�f�jw ��A��XM@�O�:B�	�YV�<�@�Ԅ6� ���ݞX�&B�	�}�"XAA��76���)��i�B�ɢf�,T��H�lh*A!Ya,���"O�����T@��x;��D�����"O8�jY!o/���6H��Vq�1"O��v�в���N�L���A`#A�<����L��"�d\,�.��g�DV�<�A+˫Do���fY�Y�*���T�<)1�ֿ��8BW)������z�<Yg��~O�@�̀�4x��ACo�<E[�}$m�.�1;�<�R��n�<ɗ�ӻ9B�u�ă�	�tB䩉m�<Q�$�oΦ1�e�VdT��b�Kl�<�!�3���ၽZ<[�A�f�<����&���B�t��"���c�<�d*�1DP`������B}���`�<� ��k�<��8Q%�ŵ�|e��"O�xа"[p=�&�|�"O�\(r�C9p-Ce��J�Ȩu"O������i�$ ��< �B� `"O@�"c��B-Ne������e "Ovu�TO��o l�l�&5�^8*"O�@R�$�&�()���f��f"O�]`��ܦ5�*(�c�A�jC�"OFxK��R+n���5M%{�J��"O�}�篝����aˋ?*L�"c"O6%� �Fڱa��(Y�"O��	Po�{�JЃRk�m��E:�"O���l��@ʨ
1�[�?��L��"O�U��0}kp	ӏӺ`c���Q"O�,A�@�Y�@9�E@�e���"O�ի�j)���G�����"Oʘ����(E��ۆ�[��t�"O��p��N� 1Ģ�ʘ�LLPT"O�%#��L&`�6u���B��[�"Ot ����`�Y 7�/���y�'��M��g�5tc<�㒃S�@��t��'GX]
��{��U�Z�(����@�<�q��3�P* ��rH��O�d�<a�ʇ-*U`dΊH6v��/@V�<�!@׀U�f��4�E�`�r�2�O'D�̰��D�7(މڀ�G�'�D���0D��` �]4�|͈��ǳb��<J� /D��S�n��~�&��.lq���(D��J��N>A� ���l]�5(,D��"eL9b�T0�uE	�}�)+D���IʤL�c����6��`��O'D��	�!M��L��DйG�x��a1D�<����|�`p{3IMyVh�rbE/D����E�X�d]��nU�W���7�!D���T�J�_�$��.n���qP�1D��A�ˍV �	p�͈[�b�y��,D�t0�P�QX>Ȋ!�E�d:pu@ׅ%D�P�0b͉sd)k���h0P�d�-D�l�֏.{�,��Ɗ�,l�hL�gO&D��`�-n��Jeg�#��8��,&D��� ��)�x:b@��r�b��(D�@j�#�$vZ�R�e�<&Qs$4D���p��9sK�-K4��3:�<��2D�h�#D��+� t���D �،*bc;D�P����!�Z�2#�� i�͆݅�L���c����`GF�@�&���` �Q��O"���Q᫃8�ů9D�\	��;E�x4� ���8�E�Bk9D�̣�ϔr-t�s�G�i:���5D���rBQ�SP����G���uF4D����j�0+@q@�+��$3D���4-�3c2ar���O�BM���+D�HH�"B%Rv��9!O^� +��0�(D������=����SC�	��LSB+&D��Q�0�����Ɖ�2��dx��#D����K�	R�t�ӡ��' ^�k,D� ��"�:ɀ�9`�ǒ
�� C!/D���A��9��jD��<S�IK�a-D���S��l�@Sa)^�G*}��"+D��ѱ�G�~�L0�'Ǩ��<SD�)D��XW!$ Iʍʓg���ܚ�=D��x�N9$^�)�#�/�ԓ��=D�`�73!w\��mrh�b�g;D��)��Y6N��u���	1�V�7f;D�� Lt�B%ǈ&B����u�Ӧ"O�P�J��uǬ ����"O�Hh�(�)v��A�i�,�4"O���ץY$E����ĝu(09(�"O�	���*;7�s$f�t(`͒�"O<
��_&V/�QiF$&)l���"OHܛR�ȕf�|5 �L� ;����"O>呖"��=Z� 0 ,/���"O������!�A&�
�Ѹ�"Ob�B$��>�$ҖFP*k8p�b"O
�R��TZ�q�����x�A0"O�H��N�Y\V��f���UĠ �"O��c��)���Ja,��"Z�7"O�cP��XY�� 5<�sE"O���Іmd�UHF��:G	�<3�"O����ʧ����ӊ#���b"O�D�È0�ѩ��C=�J��A"Op����y#Z�Rg_���J�"O`��w��M� u���v�D��y���A�0aD�%B�Ph�+��yBj�,?�L]�%j��?sPA�v�S��y��O�3�P���Í�=�jи�&�-�yB)�,j�p������4�Fp�IՆ�y� �*4{���+AI���
�yb爠S�t�u�[.�T���1�y����|������Ŋ�sm܏.��B�ɻ9�>H�L��k�` ��#�l�B�I9G"�qgS�aJ�0x�M�
 ��B䉷7���3�{
Ƙ������B��!n��P�@�r�h�ä"�hB�;E�ƫOh���yѬ�&oK^B�I�3̸�G	���΍��BB䉚p9�h"��= <���2%�bB�,fmJ)"�m_�r4��/�XB�	�[:�HH��ƓoA���7�T�` B�Ibtp�(�Z�:p���U8B�ɗT"�
B�e�,��D�ވH��C�	%s�>h�ĉ��&�B9��G��/g�C�#��%cʘ+��I�dL�`V�C�I1q�r@���NؤɉdA� �xC䉤��s�^p��ӉV�%UbC�	!oH�IY	
� �!W���C�	�R BA�$��M����XKzC��!�1���ݫr���ʔמ�B�?&��a`*K3ằP��G3%<4B䉡.���3�9Q������$B�6�JA"$�[�F�|=�$��W�C�	Z��-0�P�&�0�c1j�4jC��l��1�)Ł.�kp�D6cG�C�	���b�l�
A��%:��O� nC�	,s�n� ņ[�2�6Q2%�o:JC�ɑ�� �����]�v�˥?<C�I�W�|H���2&� ��D�a��B�I�	q��"� �
+�ܨ�0�ÐO��C�ɹx��Uk�0��X1��*VB�	�W�������6%|�D�g��0�RB�	�_Xq��ǝ�\న��Q8i�C䉹I��,�ǖ�%�̔��j�6~�C�I7{��jEb �N��4y����C(C�I�k8�2R �ep��@�`� C�	�P8h�����Qy�nΌ!8C��=wܹ�%)�^k�Q1�̓N�C�Ik��Y���R�
�YZƯUFs*C�	!Tض-3"�E��Z4❻4�C�)� J)r!*��N��dؓ!�,�|��"OH�G�>=6q��@L7���"O��r�'_:lP^0{����ˢ�X�"O(9A�E�<	�1`�wL`*�"O��Ң� >QVUq3/�"�荋�"O�)�6�.�F�9Ү�� ����"O�0�B�%����$�V���r0"O���Vˆ!Fv��\�#/��c"OFi�R�֔nRB��Q#�(EL��q"O�]@���f�����ϙ�`0pM3"O�Ma�e_�����B+V�f"O���!�[��T9�L�n�*q(�"O ��D&��l��L[-Ծ�a"O �8�����) @�c��aa"O���5*R�l�:P��Z���z�"Ob9u��	k,�j6��x�PРp"O�S��F����J�B�|�*�"O.D��A]�}|"TJGS�t�8��F"O<����Qi*(���9:����g"O�Gk�;'1(��D�>��J�"O�p�$�u�:�(O��l�J "O,�Ӷ���F��JA�]u�7<`!�$ғ�ph�c�;(6xt(hN�{d!�ʔs�1o��?;j�+��M��PB�ILG�h�a�\�z�	� ��lC�'9˔�A@F�,)�"؈B"��YT�B�I `-��I1�úK� Jugٝx�B�rPt�15��1����7o�>����S�l(�����۔w��ܰp���dK!�䙮O�\��:}s�0��EP�^�!�d��hG��@��P<��a�C�X3@�!�ā(��� �K�d�P�N����'Y�X���|��,#�e�E�T��'t$#�	��s��8�ߒ=!:��'���Qt-����9(�d�h(|���'u�E����#{ht� Y`�����'�b��B&Z�Iq��ڽnI�i�
�'�X�P��3
�jCT�nN�M0
�'���"է�9%Ӟ@W��f�c	�'L�B��$l(49J���%:��(!	�'8�9�$�H�,�����T���'��͹v�$/C�����"�H��'�l5�7��'x9U���h����'��#0�WX��H�(��b�P��'�<����A<J��!!��K�`�� 3�'
L�3ML�~xb�s��V�p�'8�p�bP�Hh̲R��<�n�
�'~� �\1p��	3�E�����'S���լ��<nU�тA;%X��'�����Ƹsb(R�F��E<��'����K� !a���"�a 2�y�%V�p�&I!$��&�D�
7m����4�O�t�sdݱ݌l�s�7L�N�C��'��'��1oB��ᐕi�]i�hs�TB�I~��x�T�O�v�-�&��>U�,6�'�S��M�`N���h8s�K�Znz܀�	K�<�t/��(�EJAK'�8���oLJ�<q�H�5����i��[�p%�5�O�<qQ*U"@��27�ɲz��h�5#g�IR�4�f�P��u9�`[C"�E�o,ʓ�hO�.|��2ק\`�=��ً9C�4ᒭ�7x�i���i��MҚJ���XBj�'�y��i�eEyb���#�~�Y���:ePR&@��y�]���,X�ƞ2ȼ�Y�k���<A��� �T@�L��\8޽z�-�*Bæ0Zb"O����+T($[�2_�4T`q��'\On�rf�P�&��1
8�$A�"O4l�'o�B�9�D�u�<��f"O���C�+W*��1�<g��Iu"O�80׌[���"bA0l�Tks"Op��ci�V�v|ڥ��0n�!��"O�m�p0=R�+7i6�'��'�0YGkF0��AQF�+i����'}��"�#DH��4V�C$H����+��W��f�K�` `���fLL��ȓw܎AsO�0=D4K��O��h���hO�>�ks��,p�����9(�2u3��*D�H!��?���$D%Q�D��%H>D������p���3s��6��h�RG=D�T" ���p�t��e�\G����7�~���O��@���A����Y*>q���
�'�A@OD�PS l�f�^�hEk
�'N�Y��K��y����&m����
�'!�]���W�N�y�P�if�
�'�n%�S-���4 ��`@��{
�'G��Rq��^,�x����W��Q�'��I!`�Q�8�x0��G(%��H��'��l��,)^�8�X #"�u��'�vm���2>p(��G�����	�'�@���M3Y��8��0'3-��'^n����X�e���@C�%v��`2�'b�AkWܑ;�L�{e�I�=��Ai
�'����$ƓHQl��wH�.}���'��L�R��8��9�Dۢ/Ҡ[	�'!p�9!�''jh�b�)ĸ��'htz��T4[^]
qk� L����'��#�ba�,Ա���M:�r	�'(��ɒ��6t�F� �W�]�����'&r�`��@��{'nkpp#�'LT����(�>����UcG:���'��Y!��Ue��g�qP�=;ش�hO?7��l�E��T�X�PQ�"�?(]!�ċ�BF4;�i�e�V%��W:�!��	Q���z�.^���@"��2[sўTE���'4�<�'N�HT�Y�d�"!'�	�'���؀�,���
��H$A�AI��hO�)u��&����C7U,��f���xR28YQ�<D��QgL*P�&�����cl4�<��O£=%>m�F��/Oӊܐ��;P�D()t5lO�➠:��4z=ĕ{�;(.�Swa.D��3���$";���E@�l��ƃ/ʓ�hO��O�rU� �"]���d�O�C�I��~�W��>�ư�ԯד#��B�ɖ&�x��n��O��{e�T���B�	�3�X0�P��! X���UDT��B�I'7�0�V��#v � �!�Q4.)�">���)Ř���b��x����d�� 	S!�V8H�Ĕ󅞻8�|�#��)[�!�$YZ�5�����t �R��*a�!�DݞI��s�"1&��RmL!��8 ������$M�yZ�+N-�!�8/�����?���d����!򄏯k� P:Ħ�u�� ���0,!�F�s�Vŉf��	r�4�j��Ҡ!��P���ӥ����B����R�!�D_�A-���?�@���>�Py��ߜ���ƚRr.Q���1�yr��":��A���?{�� s�o���y
� ��p#ƕNt�8� Ό&�L�8c8O���dڵWא	{E,�2M���b��G8O��{��9���;V�P����_"���"���!�x�(Y��j"
�ĺtb��1�!�_�H���o�_�XEBU ]l!�d� r,��E�^�*uh��=O!�DԌ:1�|I���)��l0���?!��`�%�F�E<k��@�Ɛ9s��Ig��ЪԢۜ�X ,�;A�Y�,D�Tr��V�2'�!�r�Խk5Jx���,D��;C�X��qHz�9�.D��
u+G�Q��8��[`�x�J6J"D����l����- p�r8Ul?D��1R		�,�iԒl�@�!��(D�$:�L�'c�L�U�T:)�2���$D�(�*Ή.!��@$T����"O��=!�m�35��PjVH� ��G��w�<)���@��Q�P�ʘt�N�3TlEOx�@�'��3t�Ղ"�$�b��t9Z	�'��e#7$E�F����A�A�x�J�ߴ�hO?7�	�1��A�(&4��� ��'�!���n��1��)#N4SG+ �!���"Q�AS>\4������|�x����Q萐3$N�0ݤd��C�����O���$		�  E���* .
 \�!��ۿF� ���MJe���\�/!�B1iv�jC��.|�#���n����5���<H��eSQ&��z�#C����w�<ab�]iQ�"m�qxjd)p��wyb�'�a�@bB-}Ц��q���}��$@�R�*c�7����jPP���q��4����=�4��ҧK{X�ӆg8����\��<4�,�x6�J,x��ⰢW�G
&B��;c�URU�I�Pފ]i4ˀ�)�˓�hOQ>	RF�T?w�E���]��	9�e?D��c��S��L�1���_Y�q���=D��Y�mZ ^(8�DS���1b�0D��i�O�����јLi�u�D0D��CGIO�P@~:��[2\qx�/-D����h�[�Ћ�j�0Z&���P	*D�X8�O++����J�Bx�`��e)D�XB �G6|��yQ�
&*Ś���#D�@�m�H'�[��
��j#Ԍ D��gON�9�e�1�Ә5� 0�=D�\�q�'��%ƑSJ|�QG>D���[�H>�Xғ`Q�I(H�1�.D�8x��ʩt~��ɵ�I�{ ��zV�+D�0��,R?�@RCH�
�����-(D��Z�$�(q?~a�C�@�l�f�*T@$D�RJطӞ�H�n]$E=�;5�<D��	�K����a@�m�/���0 �>D���BP Z����$hK'�!�dޏg)��$Ɲ1�<���Ք.�!���2.L�s3$�f�fH�e�G-X�!�у?��9�E�[�8z���#�M73�!�
���I��&z�E{Z)����H�X����-zwtDj���>;d4�ȓH���� a;l�VmR���9��ȓB; d���P�q�v�7v `�ȓBhа�҃~�d%0@�8�P�ȓN�Z����mਥ�5��'z<tՆ�EhPy'F�J4|(�S�բct|��Ĺ����M� �����)�@(��:�)�΅,B�0�!�ϧ)����S�? ��Z�� Vͦ���GI�v}JiZ"O\��w"�u��!hFh�=zI��"O�����aF݊�	�;te&�J�"Op�1��C�p#V�2`#��V��S�"O�9��J�Wu���>JU�+E"O<�2@-ʺ~��{�@�#H��#�"O���t� ThJ��2���(/Fqy�"O��[��~{
qn,&y�@"O�8Sv��S���gfY�hj�ѱ"O\a�����b�i>��q�a	�_v!��'���$n�9(/(=8����Xk!�d_
�U�gI y�A#B �,_!��c6|��䠙�J�Lh�b�S�!�$B�S&y#� �\�܌����c�!�$7t��}����0\�"�O�fS!��,~���4�L�p��I���K�8�!�D��DJN�AƔL�����FWt!��F�?���1F�.m�q��cԾ1e!�X�iJ�j�;����[�EN!�̌�����eތ*�:�zH!E!��>0~�D�Yf(K�q�b��a"O~��g��;H���P��^�R��e"OZ
��eP <I򦐸
��1"O�y@���+C�̌�@E��a��@��"ONxұbDZ�A��2�^�І"Oֵ	fc�>g�R�j�d;s�"O��d 	7D��R!�S+_��)h�"O���m],|@	�+�C�`9�s"O��Nz�5��C�<�sa"OJmS�̛�.a�x�)\�g֠�S"O�-���G�E��m�H́/�͈"O$}bVɢ�|X��^���=3�"O�$)�F�Gc��`��%|�A�"O��#J�	@D����_�Rr�  "OF,��A�
:lD��O�T���"O^���	�h�\�Y2+-6��0a"O��
҉ҰjD�a��
_wЁG"O�ɐ�#���@�_.�.��1"Oҝb�  7����X_&��C"O�h+��C�P�8�a����j"O6�(�E]�m��#r�O�1�͋�"O�	F�Q�:f����s�8۷"O,t��H#tP\��"W-ɤTz&"Oj�ɒ��;���jaHS� ^2iH�"O��M~à�t�O0^�7"O&��tŃ/bT�� gf(,N�J�"O� ��ȑ"�P(`�8;��"O�@�.Χw
$(Q��75#���"O~C��Z�f/�a�(�8�ux�"Oj0�фE���A��[/%�&�B"O�8�C@����]/�|���
�u!�C�FSq��[@J(Y�j�j!��\�>�d����.�}V�B�h!���^+����F��D? �Bb�Q�!���^�� I�KLNŢ�dR$J!��Q�&���ɲ>�\�����f!�d�+U��ȥ
Ӗ�4ـUL�$�!�ձKh�Ȼ���7��
�̏F�!��ۜ�]��m�> ]:&R�H�!��;�1�=f�BP(Y�!�d�N�L��띮w~<���љe�!�$��d��9�![6>lܓ��E5/�!�$�;^y����� ֌{���4�!�DV�C�M��.f��Ѫ� &a|b�|
� ��r�!��yUN��� �Đj�"O&%YTBJr y�����r�"O�a��Z�v����3�j���x�"Oj�#��W�b��x6jB�y��Y9�"O9�)Y��E`�5����'C�'u�L�a�ߧwJ�Ȱ� ��'�tX��ET�2XQuoJ鴈K��D$�S�d��8H����߸c����(�	�yb�T� ���GK�3y��{�Û�y��J�(/j���eY:)!�(�g׾�y�l��{h�q� ��mffD�1�	��~��'V(��'!҅Zӆ�3�����X^o(\��*W.��Y	g�	2!�d/7ܞ� �ͫo��]�)�8G!�U�X��\��%�=Y��Ȧ���D!�D̍�0h�g��afʸ�2'��{�!�d��Z6�e�ȫkL�{lC�I�aV���qk�u�2|�@M��e]PC䉚h�t	���@�{~���%�{v�C��}���oڌY�$���� �N|C�	(C���:��(&nJi�F�H �C�I�9L�}c�#^���IiT���,:�C�	U}�h��^�H�����Ń�"L�	N�����9;$�X7Ё�׊�3'PA	�"O4��1b�2R#�h鵪ٗlO���s"O0��#�[�F4[V* 
=Ω[%"O$�DK��Q丧��9*Q�ȓO��9���+y��c5f���Rj�'ў�}�p cU/;9�|sp�ۦK С��~�b5�4�zZֱ)W/���^5�'�ў"}R%یL��ꁣ��Q�8ͩ�l�f�<�����P�8������:wt���k�	�0>�V#îl��@)���~Z�c`Vg���ϓZ�J�p�$ZVA8ْ��Ԋd�0���u��BfSa�N�2`�-C񒽅��� *	$�Y`��X��Zek�"O�E��9,)�k����%�n�!�"O��R��
a��H	�w����"O��Q)�jY�IB�Z1�~x�0"OR�w����R�@/�����"O���tFڐ\ �'$~�5:�"Oh�_�$�H�%�&BX������yb��-c��z�֓�Xd�a��y� ��s�6�IA���';�8�@H͐�y�,Y
2��H�)P�Ixe-O��y�a��<tP�#�!�Nl����y�	�<l�	j�	�3��Ҭ�y���?@��0z,M,G���`����>�	~����\�efj��o� I�H@�o�G�	Y�'�q���H7Y��L8���dS�w"O��h� �-�iȖ��b<~�s�ቖ°<b ��#���T�b=!���!�!���H�֘B�FƖƠ�&i��*����'��#}Γ����C�z�Ѓ���WϘq��2_6؋� ރ,2���M�P|<Γ�(O��=�;�l������f��D��'�
e���}�i)�N�A�Z�zU �@60��OT����/���Տ�'�����T�TK�OP�=��Ru��A�h8�(��f��v"O�yר
u\h�00�4AM�����r�X� ��B�������P�ܳ��5D��h����h��L�c���`hR�-0}��'�]9��(�t����������'��BL�6gv�������(Љ��� �ͺ!�^`���N�%D*���"O�1����Ha:@q�m�H��"O
���8�����D0o�Lء�"O�#�+g������jؒL�"O �����_�L=;�G�.@�b1� "O�并m�Fg�г�&�w̐5��"O�%A�=K�)��X�Z��w"Ot�`�?�Dp�5�ޫ���4"O(l�$9Zsh���!��RRYb�"O��H�\k.�X2K�&����"O��9��Gv��������"O��1�,yf hx��] r �H�"O��c3���T'���I8$鄉AS"O4%�V��b@8)A�J��H��"Oh�P&ㅭ�~��[�p��yS"O:DdO�0&��Kc��:����"O�U5�?3����B �g�`��1�R�����
2F<Y��o񁄧��y2����F�b�%I��������y­�eu�0 ���|�4�-�y2��'Rc�4��c��(��k�n��y�d��&�����M�+�2���y��F@��`'"��$A��-��ē�p>ya��2*�����&.*�S�ǀl�<QQ�ҴS�jIm*�aB���P�<��
�U�q��G�4^�l��2A�W�<I��G�i� ��J+U`�*�m�<A�(�Wg��c0e�A��Â'�O}r�'}>�"%�=r��댘|�NĀ	�'x�-ЉZ*@�z	)e�Tm�8`�'�tŋ�h��j�<yra�!^�{��)�i*{p��Y#�	�\�4����έ�!���	��(��Cz���%R;.v�D"�A�D��,n��	��Y�ZjhRoՁ
`!��/��d���r�B=w�$۴��'a����\�f�ڂ~H��҇g�8I��!6D�p����*b4yZ3���9p'Q)�y�ྟԅ�I�CF��*$N�6 ��]�@��
�B�	�I����S�A��u`J�$��B�	'`�x-���Y�x�(a������	Q��h��$�%J@`$��Q:)у*[�%h��$B<4T�!����t 8$k��8b�B�	x��t�7�{��g��x�B�I�Y2����%����/kъB��͎��ĦS
���R�IH�b{pB�I�$�Lu[�V[&R@
��
5+	�C�!�@��d,�	G(X2V��*x�PC�	&6h�AR�\�9�H�f㈾-�@C��1O�\ ���HP0�au��bs<C��XH����O0V2b�2c�B �B�I=c`\`!�&p�
�@ˮ<;�B��]�Z5C����LY�V���SFB䉟m�d��UoP�MɌ�r� T68�B�ɋa�DXt�Af���s�/�a��B�I_:��R
�v� �8ɬB�I1-F���M;��� �#��B��%ɼɳ���(S���.�[B�B�.����DdH�B�k�P��C� a�Ţw`��Jk��gڞB"�C䉳d�)z���:-Li��iL�C�ɒf��=a`EذxP -rN���PC�!;�M
�Ky���_�XO$C�ɮW�2�����k\��O=��B�ɧ�b ���3Z�T�؇훦�B�)� @���
�HR�"�2x��
�"O�u��
M5�f,K�"�
l�MpS"O��z�L�0r���@\�HO�=Ƞ"OT�En++k�̀��<X ��P"O�}��ҧ9K���"�J ��"O>�s��Ɲ4��1:�b&(!��"O�i)����`�X��r	 �"OH��֠����%�2)�&��9��"Olm�ǁ�60��t�S:�� 2"O�1�5�
I9�,xթ�*��5)�"OD�Q����V�*�>�Z	��"ON����V�o���0���N��=�"O�I� Z#|������R�����"O.��+3�aڃ��#~�Y�V"O�P'��* d�8Z�-�rD��#"O� B$�X�-'��JPm�51Z��7"O��@�K�O����G�J�h��"OF!�;m�i��S �^
"O�y��9����S��S��u��"Oź@�[3F|p!�G�@u��9�"Oh�f�ݍ;|���"�xn��7"OxpQ1� �m"�5a�!�8a��5��'���x&dL��+&�ѨSJ05*��i���J���"����@j�<A�Ý�s��=���\����ϕe�<�! �$vɮ͉���)f٠���F�a�<����,}�	P#ƞ<RD���L�a�<�c��F���E��>���jP�V`�<��J�{�N(1���\Z�H׬�d�< ��7!�m��M��W���3�`�<Ic�ӍA�A�g@и��䠇D�^�<y��:&��p(#b��-���p �Z�<ꉅ!�fQ+�OY�AtH�RMZ�<�4��9,Jp�ԇ~$ܴxө]�<���;b���c%��3XԀ��b�<IGmJ�䫢J�F3n�PeB]�<Q��R�AU�T"m"�iV�T�<ѷ�@B6(�!��H#[��� �T�<Q�f�	fn� 
�&�	�A��k�<1�
�}Q\D��@*����`�<AT)�Q���m�� �B�SX�<���B)�J`�K��K$DH���]�<���<؞��*T
u�(�ۣ��Y�<��K��q�6�$�@6����G��H�<�WPoN5%�$����r�F�<9�I.AI���?5G2M�ע�@�<!�ɖWO@� �Z�[�����}~2 5�M+�Bs�i�YCW����Ăx�J�R��)n
R��?��~�o�;	2����^�h`'S�C�Zu`Q�#R�A���ʀ"T�G<џ�����
[T�H�K�
$��8�;�e`K
� �D�'l����O�K3 �K�j����2�ȥz8>؈d�B���?�Q3����QA�7�xUh���h(�]��d��`���yrh0���	6
�'`�����=|�E
��@�Dk�'i(�[�i3B ���%o
+Z��H��r�>�Ih�<s���
n7��f�H�{Wk��R/�`��>O6[��j �6�"�Z'�G�7�a}�.�)gXAR����PXT���H�!f!�4d� |aťU��T}�@� LH�݈��ԍE|*N�qM�@ ���^)��Q`KB�HO�1e� w:�(�K��S�,�eaI�Tzڸ�@��3�N���J@��X��ۙ�:��m�M��|���f�e�6-�1V���[k��qJ���7J׸`v*Sy��e��'#��m�T `�.���5&��c�Zd�P�Fs���iK:�y2n�7w(pG��+l�Z Ӳ�å$��aS�p���n�f^�]�$T?y3'��i�D�b-'�y�F�6:�P]��x2j�Pw49��I>3��L*R�1	y���IU*V�7� �A�+jE�`���U�j�S�#N��ʔ�f�P5��O�$㊋^<rq�ŌՅW!졓��	�m�,ʡ%���"�*�*�*��U����Rbp8�-���ڔ���Q�!�Ѕ��N�	�S�? ���dܝmz�J���*�X�x��i4���#�C,Pd���E�*�T1`�:>�0�%� �8P���{�&C0rq�/V7 �$|�Lh�<��
�wSFh
��\T�x�1D�=o�4IGe�$4ıa�H���O"2�Q�n̨i��p�������T!�H�� �pj�=�O�i�� 8W����w�9��%FOy�`�%ķ
^�*�nX�xYpX�d'�5^OVX�pa�h�'��uR�
�9z�Ę�*�ej�������$�Z�Z�n߄9<���gDؘ::�u�'��	|��r��Q8F��P*��Y�o����G��.t�����2=�9%l]�89�U��
̆J��Q�P�ĉ�c㘆��@�ī�376�A��\9=0�M���?�"#�6��0�nG�C05��#D��-$�f�B���;;Hn5��
Z�0�R��䴑�#�V�Jf~���?][�/#���8�+r�<[M�[�@���"#�`!P�4�O�@'��n�q��G !��j���U��e��*�%>vd��-�t!���^��M�s�I�b=j�y�-ёSZ�Y@��n�#<��MߠO�p�jS� %�2�2c I�]��9��L.~������}k�dr�Nh٤��q�+)ɮ��D��)� ��`��? ��Zt�ڡ=>"$����(��[2�(C�!�3�C!.�>�ʰ�ؽ#���'�yW���lά�d�݌g�RY�LA��y ��I�H�Q@��\lN���MA�l����Z��妔?J�
p�^wL �
���8`�a�OR������)c��
k]�̰�o^(5��z��Z$4"�gJ̷L��`e�@��c��
Ѕ3I�[X�x4�^26)@�Ap�\�4��H���|�8}�K�)u�
QCX=YqO��AL	(=$�#wi�[�RУF��􍰲�B=s��1T-�)@�j�Z��	�S���J�!BЄ�����n=!�EE�x�|yQA�2#)(h���WWB �נ:S2�C��pIueD{�pqYwˊ���w@��[7@[`���)�.ԢV}6�H�' ��G]=y����G�7p��b�a�+T�كǍ�*{VӇ�q�:'\�����§�0�!z'���!��-��8�&�7R�����OV� c&I�.��CQ玥N�� �F""�KBe�-y��d�D�_��~��2!]X����' 
��F$���wd�#"T�a�yR�P� +B��@�#vx��*�8{HAHҢDۦP�����n	 ��q��!+^ k,A6��x��ԓ�<y��J(dZ���/N�g�Z	��(Rv��j�F���� ;.�$U��J)��į�1�y��3*tMZc"��X�x	��X��y�"^�|������z���4���eI�O.6t���\�1� p{����]�j��T�x��)�O��s�H:G�������4]]���'`��W )�4`�_(C �[��զeU�IA` �u.P���9r�FQ"�\��]i����0<�E��/ZṆ]�{*H!�`K�R̓z.D=��˟�Xl�R%�l'�	�Wbձ	����@WL�� �G�]/!���$�X��ܘ��).�O:�IFOT#/�4�I�X78�d�+�R�R,B�d�.��#9FhĘ���U�)�&�#F	�~:�&U�z�}rΜ,+V���!,pul0��-WB�'��@��Y���%>}[�a�2|;�P5~��Z6�_�C��3Ӈ0�u�ǩ�*`��yCġ۽6vn(sqN���ēm�.�`�ңML��df`q���x�azR`&1w���?��D�Ma�|9fGI<i�<���
Jtt
Xy�L[�±� '�}���)��B��`��
say�N�7����$&?qg΅RP�'�tC��'c6�7F�)4�ui�������&=uhҽ"��&�hKa�]P �y�é�hvD�Pg�2��}rn�3��M9�mY���"p�K8��t���ůd�����i `9�cWj����%��?�*`����1�^Yb#)">����U3N�f���	�V��\��Ϋ#�bI0��*�ӂ)�����(Jx��G'�Z�^0��/�,A�ʝ���]~p
ɒU	e>�"�/)H{qO$ 
Rfů'����5mY _�`�X��'gP�RbZ�_ق-���
W<"(&>!;pY�r@P4��> j�8�l�/�Qk�j܏��+��� �J����Z5��=�UO�0IFL�u ڿ8RPP��O�\�8��dD4_��˳EķY���%��D�]�i��|1���;L��ߝ�ҵ�$�J�f����!�ƎEa}�#D����C]0De.	�A�� L�;cB���%T��F�tʁ03$ ��
�Bn:-�!�O�S3�M�k�kI�q:��!`W��BБ����'܄���dF:�2��a""���V��I�5��@�� �<��jD<h�����Z" XHQ��!<2E8�Z�T u��`�h�"LۗFɄQ�ԽJ��4E�O��%0�k�	9M�ʠAB�a4pU����!��Śnh�x���O6C�l����4a�J����L�Hx�p�����x{�ʥ?A&�8C�w��E#�l#t%S1㔳`;���	�g�~��#�4m��1�$Č%{D�""�(Z��< �%�NH�x��Ǆ1�p>����`���S�
� ����`�V�'B��r�T�A��%%B�
vJ�{ ԟ�`#�X0;4YR�'�!I��<K$"Oz����K�v4@����ߣx�����'
�4A'�D;+���_T�����,�'J��0Ā*{�$]I���8Z��"
�'�
 �q��M�7O�2�n�ЁO+qr8�إy��	S�ꗌ���I�X��8B$�41�q��h���Dδ�0����<
��] o���R����X��� M������� ��d��~�J!�ҷG��g�Iv�j!���F��P��Ȁs�M�h�ĸ�cIި&�N�����yr�,SD��قӷ~r��Ul�~MN�=�����c,c9�<��ӊkw"��$��7�\X����.�C��",30U��`� ă��.Y�H%�J�D�'��+\��&?���#�"d� `���ɱ��)�ԙF�
�4�~���э_���z��K)L�AON�p-�>-�v��1��%ۺ�"O5��E;}PX���XT�(V"Ol y���+ e�hs_�x+"O>Q��O�	 �hb�C4��q"O�Pq���,��Ċ�Η;)�X���"Oh P�V�Y��[�� 'j�ٚ�"O����$�Rp���N]Y�T"OШ�F�F�UT����'&aQ��"O2�S4�N�'!�|z6.1(���"O~�K�C� ���V�<(��� "Oޤ�P�G��8�H�m���"O1���a��I3�ޠZDPR"O�l����O1��C�K�=G�캇"O�T8B@��:k=���
�?��p�"O`��J�@��y�(�!J:�b�"O��%ڙ@��j�br�9��5�y�`F6W�0 #�$<���;c�̬�y򈜔(8�8yD�{�J��B�9�y⦞-W�\At@�(~JV9�r�W��y2��
1ʐ㋶ls�t����?�y���:���$S2��Q5�y򪑬D�馈�+閑���4�y�-�%m��A���� �ղ1��yR��R�|�A��N&Rr`���L��ybk�$��������0ujO��y��׈h��d�ÃQ~PwdO,�yBԒJ@Q1CIW3Ux�9�c��yR�Y'��s����&f���&f��yb��L� ѣEC�`y��DW/�y�K�&�N��􇀰`&Ry�0k��yB�ׇG�(PsE��J��dsA޺�y����0�[�ݵ~��5 �O��y2�-p�]rG��5!�0T�5.��y�%�/I�t�	���� ���KP甌�yb`�i�L}�E� u�AS@앏�Pyҡ؆c�cc�qLV�K�ˇQ�<��E�L;�e��5QЅjW��L�<ia�Ef$ƴ�)�/m%L�5	|�<�Aj�26�� �f�R/	q���K~�<��aV9�&lᦏF7���� NK{�<���ɶ�@��	?Ox|�SG/v�<)�c��y}� ���.0�q���K�<Y�
Y�?WZ�3�-9K�(�O�F�<qD������Yi�Υ)7HQ(!�d�
n���WJ�?����jL�h�!򄛥:�I#'��8H�n�s�KS�!��);u�dC2��2R��0SP��	9!���g�4�
tK�<q����3-��nv!�Ĝ#QM�4���u�Ȣ��O�@�!�M*7�50�爱QRĽ:��\�.�!�$K1�sr���~�t����!��F�&O����N�n�޵�K[�!��)snSK��h��)�5���!����N��H&r�*	X�k��f!�D��#��P�g��/o}� �ꟕ�!�I�w޸J��ҩPK��q(Q8~g!���
�4�3� �=nf�J��V!�� h�S@�F�n��]9�6n��"O���N_�0}� b�H�'H����"O@a��U�x��� �ǁ�$��"O6*LH GV�����;\� ���"O@��F��o��Ո��i0(��"Oz��A�_�ncҴ��A�?\��"O��B�%PUÎ����ƪ��ݛp"OJ�ڃ�x��Tc�KZV��S�"O6d+5ȃi��YP��\qT �5"O�U�����CՄ�8�Ƙw
^�"O�,a3fT?/��ƅ�q����"O��c��ECI��_���D��"O�rBbD�U'�Qs�8_��E`�"O�k�[�=�V8�qD�5e���Qd"O��;��Q3w�ˇÇ�4�t�� "O&�q%"�r6"���Z/q� �+�"O2����۱M�80�k�	~��b%"O�ݚ�+D�+�l p��j�8ZW"O`maP�������&�����@�"OL0x6]t�&��q�A�$N�\@#"OV)� (�
iZ�A+СP�9�xZ�"OBP��J�u3xĪC������"O�BՇ��G"
�YE�Kl\��"Ol�f��A�G�2���G"O޹���ƁO��$��Gѥ����!"O�4�Pm:a�,�k`�X�؄�3"O|�����`������eꠥ`�"Oa��b�5t�~e3N�!1b�R"O�p"ͫ/�ҍ�4#�2j6�t	�"O{,P �8V��!it�F[�Ѕ��Ɲ���C�{c��X#B�q^L��ȓm/��B���)9��Q�ح�8ԅȓ�2�jq*�#���+.�t����j��E=H�� ��L�6�ȓ{�\5�eI �7�(�Z#n�ȓu��@�QOQ6	�npk���#
�b��
�d9�AC\��q����j�N���#��q&��$)���g���rm��\��L@�"�D�T⒎}[����FhV0z��Y�~ز-{rc!��H��IFթ�gڴ
>@�P�:B��(��KT���w@؁m��$b��,�hA�ȓi�b�)� �(i��s��B�p5"O�Ⓟ�#L�4e���S�/&tU��"O�TcM�n�-+P/ 8*���P"O2�%��K3�hCn�?�e��"O��E�Fe��1R��(���"O�h؃��aX�Z�)Q9���"O���8��x���F�K���2@"OJӊ�/z�J<A!An*��#𐟐p�bӾ����xZw#*,8�%?��Gͨq���@䑹v��C��T�ր�7���A�`C�?�2�!w�I����;q.
����G-f{G��T�'��Ấj�Z��ق�fF[[j������9^�Xu�0떳Z�������Ԡ� '"�9�̵~� <ن	O�P�`2�O՛djJ :��t�"c��m0�'����/��\}n9�~�܃$����y�"���S��4a�c���}J�&�I�C䉇9��HD)�;cơ�ߨw2Rt��4�"QbG�����׊������u<Ȭ�,V�U�h��6��@�U��H��(��FIVԇ�	�r����w&S vX���U�N�2��3%.������]���QE���h�ႃ�YfDэ�d�
C��@拙�rl�w(߻T����U�������c��-�!��}�^�RB�8o2F��DNA2\�D�{����C�0���U�M�,��ɉn���w�M��mZ�&]*2�7�����8H`ʄs�/���0mQPO�>(���f�z�\c�� XD�=eBb��`�c�`��'���J 	�+Q���@��I~�]��-^��Xܩ�Ѯ[ػD���)��+�l�"P���9����S�? �9�F�Bl(�أӡ��W����'��E˼ �V@��̈/Y�U�c��%�������B�%��?|��*�[��|�A�)�`pb�*�fK#p88�gc�Y�J�Ezrʏ�;�F!:CEл����q��-S��$���ԟ!�R$sČ�|���2�&E���q��3D�|��đ,2���e�� ݂��"ǟbm�fƜ7�:D{P@��Wv���͢Zl�M�!+������~��}��p؄@\��)P�H$<��6�&l[�(֥ro�|IRCKմp"S����r}bW�hfpYb�[���	%ph�T�㊐آTΓvb��`t�/t��XI$`�g��i�����xu�D.�<.��/�t޶ٲB��'� {���k�� y��ۯ,zD��B�0s4����DV�E���Be�x!H���E��,�ў�լѻ��la�_�W�*\����_������lIڀ�AL	m�� ���./����$�H��$�C�E��,�N�D��~��q�+�0u�J\c��\%�	��՚B��knķ@�'P�s�E!LºHx��'s�)���M?j	�C2�N���H���T���F ��#����K%~4���OJ��1C��N�b�'~l�� ��a��Z�F-;(�5��ܖ|��+S��D�CT"#�<�P������j�J�'l<R	Zr*�b�\`���U��xF|2Jߢ�����ڄd���+��Ox!��+T>G.<}C�M�7(����!�X�#D��^�X��]9s9� s$NE9��I��A%�p?)f�d��mV��`�aC��7cE�I`v�7d�h���fߵS��IS��_�c��Y[�Gb��{������3~��b�*S*+AX@xª;D���DmG�	t��&�
t,�!t�:I�n��'O�iȥ`�ÜE�T֝5	,ȱ����t"
��p'�>��J���F$&�Y)�6(�z2�	�Eш\���j��hp�@O�Q�\��ŀ�/+��=zf̋�R ��a�,T[f��"�� bϲ%�	�	�8����ȿ������x��c����O�|��e� ��(���Cp�<��t��+��.-�6 �8?�E���K�W���!B@ n8���9��}��%ܛEں�@���!Ѓ�%MRԑ1TM��#��A�p`�>��A�DE��Aݶ�X���.  �0Y�B�^wp���`�S]"X)�"O�|�n����v�l�I��eg�!"�	�Q@���S�,)�fۡu����p�r�1U��1�^4Z VA��ɇ�Hb\A�$*LO�@�c��7!��
��O�i���	Ƣ�}i����`/J�5��g#Լ�g�:L(��D��"=�ax�fдf�޽�DH�	uf�pu�����'wn�H���$}gq�(zN��᠇׎P�En�#l�r)��B�:��:A�u")�:�|1��O�|��sxDQ�
��`�T�Q�k�=��g��b���r�H�7m�@��a�zv\q�:�D�!6�ibdB߁�`P��ZxЅ�F"O"��h&�nJ��zh̤��S�-��qR1l�!�`��Gf�	H�&���Hۤ�pג�[h���'P��Q -2�R<Y@�޴p����ӓx-�0h�ϛ;HD�y�nގH3,�(D�ڥ/�d��saγW�^���#E��a����;� K���X�x�2����+�)J�~�,�$d����' �4����ਣ ���� �KM��Qa<Y�e��G_�6���p-�8
A���f(<q�+�>���&U'N�h�b/T2�$�{�)ܜoJA�t�A�/�V�������Q?A�G�y���Ք5U��Q�*�	.�I8D��2�!Ͷ��T�@�6j���A�#�/u�\��k�>�I�O�Q6��*���{��p�3 X��ē1G�����A�3���z1�}��ɿv��PWN�gW�8��F27��@�&���>u��̃'%�~snN�h�|���풦H�:|�剬a�RA��<$�̑�A۶\X�b�L�����!��Qru!��Pk�₆h�b}R��%Uߌt[U�\$9���׶XhVu��Ox�����]ʨ '��-��l�g�W?[��ڇe�24��YN$�kA+�>�|��J~"�w��"��*&Ȋ�P�l�Yd"��'��l�&^�`29CӃԧI�z���7Rk�:6ѳ59@m��KG ���ިa05�=���۠A]�-P���r|d*�e�|؟(��7@U�S��	%�z�bGO�H��A.2#f�`"(� > t���ݐ!R<�0��ߗh�jXr ї��y���j�bHR`n��~���;Kꎐr��� `3���D��yb���i�d�ή Z�s�/����'!X�c�o�aW#��C/���J�ዀ~��9&��p�<�e�X/��Ќ���ܚ�Bl�<A&iI9'���c[Y,�8$D߭o�!��.mj������t�k!Ù7{�!�d�9�+T��P�2��W�5�!��1s��UY3Fwx���ʡC�!�� :��۠���R����Үd�!�$��G��9��ܠ.;@��7�&}�!�$�1.lh@p�Ҭ8$��K�/m�!�D
�?��m1ǥ֘;vA�da��!�� �1��IK&;����$*@��U"O��Ӈ�O��ak�Cطi	���"O t��	ʈ��WO�<3���B�"Of-�2+S�$S�}5Rr���"Od-Á��3C�D�V�D<1�2"O�(:�O�;�a�B!U����*�"O�DZS�ؚ!���r��3:�*�ѥ"O�8�5��<&���6��m����"O`�`D�\�X���:5EW(/�|��""O
Q���ʝ�ir���@��@ "O�eTl�!#������ע5.�9��"ODq�ÁQ�W�ƱZ@o�،��"O�Ds��
�}�rm�w@�P	ri!f"On�CudL- �ɣ���\�TĚ�"O�e���1x������l�D��0"OֱKEAU�0�F(� J�˸�p�"O�}��l���@��A�}r�"O�1B��� T��k�L0셃b"O�<C�_v���s�I-����"O*�3�Ē7x�I��Ή)���"On\�Iȫz?�%�ň�=o/���G"O:���D�l��r@$M�J��hS"O�%Y�A@�U �!Iê:{4���6"O�Չ�Ŏ�A#V`a	ś*j� �"OT������q a
�,h)r"OU'�\#����˦�:Y�B"O�p!� �*t�v` C��o�,)�"OS�������bD�X�*XB�"O詪Ƭ����L@G&�u�� �"O����5$��'e��W�:ٙ�"O�ta� Q�LkT�`��:\�p���"O*!��+��@k6�N�2V4�J�"OLy����d|:��d�Okl����"Opd�T*� #5��Ƅ�[[��J"O���"�$�rX�3-H�>�,4+�"Ot�Y֤Ґ)�.�5�O��4r�"OX�r`�q��l��L0%�f	:r"OzQ%e�R������A/u��QS�"O60�-��cj�!�����*����"OJ�` �� ���h��р+����a"O�k����X�]�ӧ��p��q��"Oʠ{�!-J��˅�c� P �"O�9*r��[
��ӫE D�.��"O�x�1�ǳG�Dٙ"��;���"O�iX	�y亀)F��gɎX�Q"O��*�#R�2n�%x�E51_JE��"OUzUGLV�<�s&ӽvE6�:w"Ob(��,�\ hʲ�����0"Oli�a�6�pQ���8A�P�sR"O�M��M� H�����B%2T��"O�0A���%y5Rݪ�*W���u*""O|xR(D6j�LD���1�T�t"On�Z��H�%��rM˷_�5"O�x�%���c��a w�@�`L��"OV��n�9j��Y�T˦'�֠c�"O�ɄHխ? ��`M�|��a!B"O��D���D�aO�J�L�
s"O�b7R�E{�Y�å
�ƪ`��"O��"C؛>���3�_7��@`Q"O|�ZaMM!i)� P#V,a"O��:�l�� ��)��k(ʜb�"Of �C�F��� +u>�d�x"O4AA�&�`�C1��[�8u8"Ox���9Eipt�qf�?#�:���"O� ^��"ʝ��-�1�ӻA�����"OzT�&_�F~�!�^�"o&�J�"O@<�v F?䴘1C-]�8}0"O̰�6�I�]d��$�T�Z�r�"OF�C���*u��,���&b@Qj�"O��2�J[�1 ��Ql@:U�ma1"O�tP��D���52�'S��Hk�"OЄB���DJ�D
�1�J ��"O�22$�`W�l3&��)�n�c6"O
�zS!�)L� �1��N���ˆ"O��1�hL�8��1+���{Ԗ�v"O�P��z�8x9�s�dɊ�"O�m�bN��=[�	p�d��&��d�3"O��p�B ymd�� �� O��m�!"O���s%����!�A)t̤ �"OR`�jÏ"���Q�U�ni��"Ot��ǋ�g��XqSJ��"O"��&�]	�F�2�M�5H5�=d"O�A�/�(s�eP
*6�x�"O&� f��Ar0�ԯ[�Xĸ�8�"O�%bc�����YW���t�N��"O$|9�߿�R�*�%H�S���`S"O��C�S�]���#�툵H�"OL��1 ��CF��%�\�@����"O��ٱ���b.���'�	\D�Z"O,�`�CBd�v4Z�`Q,�zu:"OD��CF[�,�򱊅N��*
Pū�"ON�9c �?y�$�D�=1�!��"O��e���d1j���H�T+�"O���T�U�GE{`PY �ihE�'B Q`��FVz��VA�"s,)��,Gfv�iAS�� 6�*�p@iA�V6Q�P-��`2.8��\�"|�3"B�.R����I�02�H�V?�BM]8��@@r��Y~����4�pp�(%@OH�K��+I��I�)ǁg�T
�z}��	5����
9ʈ��� T�00�"�b�"�������:B�m.���	׃銨����9+�����J=Z�r9����<	��2*�jF�D�O��.WF����Y[H�	Ä�r��˓fn�r�Q?�m�(!RٹBF�#+�4Si��/�t��+ �	$u��f�S���~�D�+�p8b	R�k�!���P�W���[���	Z��8�{��#,10,��I�-*�<gY:5�'�nU� �� ���HY𠫐��Z٠c�̨��iA�vzE`�"te��̊���v��?�
���!� \�	\)8�^�3a ?���s�H�Q�b�I�i>�%?Mx��9^��d� �BƩ��j?�$@�����td�'�y2l�2ђY�$LN�5`���(� ��䚧as��a�{��ɏ'FT��rㅪn�`#���5՛֨J�0Rl�X�47��i>�ԟJ�O.|�,�;S3�D�rm��u� |i�P���q%�~�5�t�<�O��s���Lx�Q�	h�$`�'��%�M��=����Ӟ|&�a�G�N� �`}r�ꃿ9e��/O����4T��!�h/?ͧ�ħc�"��Q�����r�F�8WMМ�2�ji`5l�34�ӧh��e����;f��d�AlU�x�̘p"�:���kf��T�S��Ms�Bք��`AKL(,�����F@=(fI�!
O6�ɧ��4��r��V4��p�W��T�$��&nɠH1O&��6�O���['L2$�t�����O`��Za�|�猆Oa��Rq��O���G�?%�hsĉ�r������]�Tn��/QJ�=�ԭt������=�)��v���i�U�N�B����\�C�	�e
���.��+h��kDQ�R�B�	5' <��όX��<P�Ԍ>L�B�ɦ�������
P�S�d�B�	-b:��f�O�(a�M8t*O4_�^B�I7A�ސ��ϔ�C��I���˻m�.B�I%S�0a��͸<�=�A�N�d�B䉪4�}��#�$�ցJ7�-VJ�C�I�g����ek">�1Ũٻa��B�I����9�Z4uJ���P�Z�^�B�	>`H 6� m#���%Ջ"i�B�)� �5򤆂�}6�X���ߊC���r�"O*itjN�C���	��<{��""O�I�D(V�h�lòABg����"O>��D�ٽX$�#@�PK8]� "O�%+� QF��t��	7��#�"O؄�FM�Dp����O�[)p��"O�1� ,L�MD����dUD��qq"O�� `m��^M��ٗ�ʺrl$�:�"O�9IR� 'G�H�*��O�ZSr 0"O��H���h��|�.Z�>P+B"Oޘ�4�,O3�	�le�2�JW"O��N�Z�EQi;X�=��*O��g��sz��é^"Y	Na��'��:���3nm
	 \��!�'5^�	&��W��)CHT=s�MC�'����&xh����i,C8`��'Z�����B��4Q���|l��'i:�f�&(
J�m0j�*�
�'ڕXc@�&���c����P�	�'�bu�cH�?O�
tP���T¬��	�'�\ġ2:}��(�'W/�y��'*p䛷�ۙTGf�0�·;�����'d0��g	ͯ+�Հ#*�DC��
�'� ��-a��8���)=�x�	�'������7��M��N�:-����'G�|z�g�<��y(���?zU��'�\��"JK'q�I��� �̢�',�4Qqh�q�1}����'�h82.^�\y&Y+�	�L��Y�'j�1�R���!6������C�<�
�'_��s�O
v�dȪ��D@&{
�'Y���3I��R�d��i=6�Q��F�<A�&]�eH9c㗫a�i��*�M�<���/��4�`��[	4�QuJPR�<���B�P����_�/�|���s�<1�[�1� ����m ��rd�X�<9�J���u*�B��4���Wk�T�<)O�@�%�I�2!�fk�O�<��dɦ6ވ[���P��4�-�O�<��"��)B����F�Qq��v�T�<1և����8� P�Tڨ|��k�<���@��b�Fǚ����cH~�<�2�
~P�r^� ��Uj�$�P�<��ƅ�p��٨���:���V�<ASH�^s�i�-%I!b��K�<	 ʝW/2`*g!��0r�����NF�<�$�y"j	��GA�����ƀ�J�<�Y�\���鶆��(,���|�<i$ ��s�.�qS̄�J����c� u�<)F��1T�;糭L^�5�` �s�<���݀��u�^!�l���AZ�<if$��2h��	g�8a1��qw�\k�<�vD)lq��e��A^�p��p�<4+�:��5ya�\[�^� ��Px�<���
�}�H�i��ܐ@P��&�O�<q���$S_�)�� X�
��Q�N�<�t���p��`�J�1��t�<�`ӛi6b�1g��u7x1���n�<Q3�I+����4LN$6~Na��k�<Ѱ��5�t��џ]�a��e�m�<���͌d��$���V�vB)���o�<�ȗ4FO�,X���@�"@canl�<�q�F�>|�zq.�-g�M�t)h�<Q�lU���eP��U�#�x�y�Xa�<� &��ŉ^�ꔐa&DJ� q��"O"m"�1i>V0���&Ѭ���"O�Ue�=�J-�q+U���U��"Ov��A ǌ�1���Ӹ۲ xb"O��k��-�,B�k*C&�8jF"Ol P#)���4�I��,^yP�"O������"@V�\��ϋ��@�P�"O��!"z%`�� O�4R|�S"Ox�As�7l���.���
��"OBT+Dm֚x�`3�MK�4��"Oh�5l��~<��j2-5.#�L�"O|�������|l����#��Y�"O��ţ^/�ڸ"AKW`��$�"O������8z�	�WJ�:!�d���"O��q鋷X����+Z�ج��"O��s)Z�K��*�eMO�Xh��"O�y��02���r%B~Y~�٢"O$i)��$�%!v%�XQl4jB"OƄ{�'Үh�M��B�3�%��"O ����9J"t���*p�1�"O��A5hQ',�j`nP�dd>��C"OXoؽqGU"�݇Fy��$�|"�)�S!d�<M���*�h���kdC䉶^7�0 ��#)�չ��4*J~C䉨ԀYS��^$��(��ڨ.VC�	�!L �QL�U�@���� ��C�%X�B�k�h]�W<��qC��
�C�I�Ku�=�ᥚ�g]6�ф��<'��B����1���[�H%����B�X�@cO�C�1�Ǎ"`C�ɧ5<������6�0N�B�	>LN��ӣH&t��-���3{�B��+C��8����?�ҁ`���oP�C䉒g�ԠJ�eH5x��idC�`�B�	"�vuSOV$,�:-�u���	�C�ɍr��QT���|��vG��B䉹qX��R��ڌ(�$���k�Qv�B��5��DRq�Ôz,	�i��pk�C��Z� ˳&]9����6�]�J<RB�I��D ǅ�V:��b�I�3~�JB�	�;�n��%Ν<z�0�FE/FB�I�Twz�3��_",����C6m�C�>HL���<Q�� �A�X�Z�(B�	�O4��5�_&sĆ�[��2�B�I�f�Y��ā6�[��8w@�C�I�P���aI��JG(4���+~W\B�~7�%1	ۧ7���N�IvZB�	�"�"�����3���"fa��Z�NB�	1)�p���Ǳ<�`B+�4(�C䉧0���ke�o�=�3�\;k�lC��)�Ԋ3�7p��uSf�0U<DC�I�Q!A�B��0p�$hۇ�[!]�B��@��S
�]���+�n��ojrC䉨A�Z���BJ���E#p�^�#�FC�*K:�z�K{	����+�z�"C�Ɂ?+Ba�ǃL� �M�PoE1D�PB�I8N�-Q�)z0īQ��	,�6B�I�D3Nu��L��^A�ď3;�:C�ɹ�)�eO{P ы�Fe'�C�	�@e�1�5P���Ju�W�R�C䉜Pg@��&G�L��H�V�xʘC�ɪ�bud/	s�p!['@�� �JB�I�P����
�'wfPVGЯD��C�I��z��D��,a(��2��a=.C�)� ؀Z���
�GF�4g�<��"Ozp���ܝWV�]C�DY�aF�j�"O��S���*U�(h�b�E�zCb���"O�K��
���9G���"O�t:%���KJ�S�A߲Iepd9D�I`\1��j�G/S٪���4D�D�A�?o��Y��Rk�@er7M=D������c�6���A�3P!��%D�T�V��*YW���l�8��eK9D�(�v�(<��ڧ�ߔT���#�6D��Zb��>#X���2��j��6D��a+��Ӂ��>��!��"D��3E��.[��`ۖb��F�=aF.2D���`֮;��0w�C!&n\��S�$D��Kׁ�T��> ^�zu,E�<ѐ
��s�)�3@J06�B���	K�<�D.��Y��L
��,L��5lQH�<$�AF�l�VnE�=��B�CM�<9u�U�Lĸ�qGۥ{7�qգ\q�<ys���e�˰��璭��u�<����`���̷d�>i ��r�<Yr �?:8��3s�S8N����##�g�<��g��&TtUz�÷�ȩSU�I�<��!L�7�p*aG�0#>��+fjK�<��a��e����d�V����s�@OC�<���Tz{���TI��*�B����H�<��ʽ\�y�"[$k��$sdJSZ�<)�e��n�lM�ШdO5�!}�<�� mp, +���jw0�i �
~�<Q��P��pZ� :�0�!�f�E�<�D��8, >ŨUdڒ� �b��D�<	$
�Z�@�2��(x��U�~�<I3�mN^�2��_GX\��I�S�<��G�oX�$�=5�Ij!e\Z�<��D=|�6t@T�͵=�2�iVeSX�<)@J�
n��H�<E\i!E�p�<�1�n� �
UW8��%&d�<��IVՆ� ��Z�6��ՊUw�<I0MаoX|0'��T�싅a�M�<���3tM^lc�#�~rً� �@�<'�[�\Ȓ��w�6�:D���}�<��/F�u=�0x�bK�z�&8W�Ar�<)V�o�>]�̇�ds>�;4D�V�<��,�)JI�t����P7�5��%w�<1�8�|����AFE*!��u�<yegц�Hq��A_0�j��G�Lx�<QF²Y�%8�+�g �A�v�<!ci�	s���㔌�6g�H3s$�q�<Y�ɒ�D��$���q&d�)n�<y���%��"�*�x�l�ْ�PR�<9��,<,ȫ�ǁ5
�Pkg�P�<ITR�,!<�b�D�y�r1�lRJ�<q��^N�U�S
+�BVH�L�<�b)�!�	��4.�Pz0��y�Nـ.w���c�ֻ3��`$�<�y"�C�
��)pV(��&�V$.��9��x�=�$�O=c�b��E�o�8�ȓkB�%���PVMi�N�%�2A�ȓ�4�j�Q�K:&a"iJ�J��a��I䟼q"֬C�v�if��F)brN�s	�)���Ǔ�?1ek�{xԘ�sn��C�X���NZ�h����S^�	Ɇ�)`�z�EyB�� ����+C6|5���˷L��ba���O�BQ�&i�0�f�J0"B),�yEy" ���?��W�f�	Y�]�p%aWV�)��Zǁ }��'MR���`�)r�Sp�G!zC��r�)���GX�� $ȃAcĖ^�v��&HȤo;�89�A���M+�i���J�N�;�4�?IO~�_w��|*@��w
��1�m�
cn��I�����%gX�&�	}�DP��O�Z��g̐f]��)�1v��h�3
�2T�-� �S�J�O���WA� �]K��β(���l�7��TRS�O��	��	C�! ���QBܶ~��+�}����?Ѱ�i��7�O��O@�d��
�S�`C��9l��P�S�T���?E�,O�R����.y���??�Hp���'�j6�Ц1�'#���&]�J��Q#R�t��24��1c��An��L�����O��Oj��^�D�Řu�?,�Ā�G�-l E+&�T�mr�}� 道i�j9�bF3���� �ݰ7�Z<ht엷GJ,PdZ
C�� ����-wz��@ �t���J J�v�������ͻv�`�:@�.L>���.F�\�)kG�'��6M�ny�Y;���;?u,LxR��^;�x�a��$/&���'�O�"?I�)��!�*���;�Fd�DM�Xܓ0�&au�4�O�����@7m��
 �%K�Ќ�,'5���ɡu	�8�ƫ�ߟ���ǟ\���u��'��i"L9s7i��h���$�*^à8�w%Z�t� ��f.�p,`��G{"Nq:ԏ�Z��O�9��S�<5$�#�j>~��Q��8�:��qcS)���W��V��B=x�h��J�t�2�J�����ِJW��^���e��X���Fu�X�*6�'9�6i�'q�'��)`���+t*��\�Ikxt��{��'v��Ə�R��(��c�E�>�*a���%��Y�4�2/O��+����Ym&��� ���P���0��M����$�O@���E�&qℲӆ	�Q�f���T ��maH�<�X}А�
�}K��qqn��&�Q�����,���pl�K�����$C���!nǺ 3���el��oi�Ј��iM,�<���ן���4&��Q�b	��\Q��ό��lP�eo?}��'a2��� %b�|�Q'�-U�(4S���Mˌ��s��ݢ���yNv(���0Z��A��^��Mà�i��I&p�Y�4�?������%8"�YwÎp��Ĉ	y̙R�O���Oj���`��	]�e84A�py����OX<$=z�%p�A .�&,��ba��d�H-sK+�I$fbl����t�`R5�H�eڒ��&­?� J�(��lYY���1&�R��D���<��L�Oy��?��i)(���o5:M���h4z�Hр�$�����d�O>˓� �q�d��Ѐ�!7n���'K����ߴ�vV�D���=J����@�w]6��� }�'��'�����֡   ��     �  �  �  �+  �6  �@  WK  �T  �^  #j  /q  �w  ~  l�  ��  �  3�  v�  ��  ��  I�  ��  ڼ  �  `�  ��  ��  ��  ��  ��  1�  #�  n 9 | ` �# �) �.  Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�� |d��"O
`�(�;���8���-0��1%"Oj4��ND^[��"3/9�0|H�"OB���H��*�ʞRy=a"O�味V�!X��!&F�:J�$���"O,��a
���C�Ą�M�"O,$3%o�-���p���+Ն�:1"O��ݢ1����`���y14]2��i�<�6��{_���c�H�`�fX�$Kn�<��A̼VI�xR[�)�Ć�pඤ�ȓA5��('nߡ4�� �)˩%� ���,��r�؊b#`T�eT09���ȓ!�b��g��}�8�F��-? �ȓ
K|m�ș�VṔ���2�%�ȓ"R�X�j�4JN�1�˘X�i����̹	_�jZ��1!g��zܶ��ȓgil,*�J�
j�Ne��i�J%b���f	�(U��:���G��$Y^م�~r�� S�%T"���k\�jx�ȓ|4�1�îJb��@ӵ�ݩn�V��/[`�"�v4�R�!ʎ<��M�ȓ`:��z�ؚh�J�Z��$HY:	��H��p�m�C1��!��B:��0��EnjZA V;9����J[
2���	��4'J�EA�IVW&��~�(aZ��ӹ�>� o�Y�|�ȓ�f�A�
Ο7�H��M�$�����mޠP����/���ANXo*�ȓTv�����{ ��-7�*h��I��sB�8�8���3����ȓNe*M�悡;������X�o��!�ȓ'lj�#F�m�+R&;�|��2)n�C��0S4���T:
b���:�0!��e֊��)��ͷV��,�ȓ0�&�8#���� ع�L�����;�P�AFd���,w�6d�'ў"}"`FŪ��:w ٢Gy��نND^h<I6�Q�,�X8y�nC�x�z6����䓷0>A0�G�9ٲ̣S�ޔ$E|4ˢ˙}�'��?�˴�ܝ0�x�B��'i|��J:D����ȍ�x�z��jW�w�	р6D�̳�eN!���M.��z(���!�d�3�Qc\�O���&����'ўb?	�v�� ��-�"� 09-c�*<�ORʓJBJ\�,�+ �4�����xu��{�7O�c?O�	Jw	Ţh�|blR2Z̈��IE�O64�Gc�y(`�`%��&�d�� +$��Y2�)L��a\(G�z����0D�l#���?sz`�E���m�f��϶��xR�!/t�'c�{��ڠ�A���'Zў��Z�@�P0lH�"NJ>FTAR�"O�@�<�`	(�GA�~<V��E�}�<��_��ͨ�)
:|I
%�a�n�<�sΚ6g�u��a̸D\���G*P_�<����;|���թ����$N�@�<9C��!�"`�W��+NϮ�9��<)G�A�)� i��E�&�J���JQ~b�;�OD��)��Z}�l�*��e����'�󤂔d����*�5�zi��A�*�!��I) Kb<*&o�;$��XC���ax2�I�>�����ԅa��Q#��>-�C�I�Q����(�pC­�c�V�C�)� ��C��5:8؈��D���"O0��˛'<��Æ7`��*��'1OU�dAM�D��)�7*N5k~)�'"OL��c�C?|�#V�4E�JزA"O�[3��$�Jp�Sg.{���W"OZ����b]X�����,j�K�"ODXP�A��9t��3I��i��p{�"O��%L]7)��� GI�R��鉧"O���-���L ��"�@A"O�L ��
7��@�R�àYεpB"Oh,���	(<�@�u, �5qDŹr"Ot軠J��*���1�+�>QYb���"OD8X��.�삳ʃ:Z9�D�Q"O�ai�*S�@ԙԇI�9i�"O��S��1�̸U��97"O��`��z�2\[q� 
b��д"O(�Z#�	8#k�%��*�)I\:�"ON��������=GPTT�@"O�1�ۺx�T�&�۸6Vi۰"O2�j@(th*u1+O/�#7"O��jԯ�/9�B��� �FD��"O�E#6����B�s���4�B�"O��"��B�XC�`�l�-k�ʅ��	C�O�l����36�� ���\�"��']��k�`�K���FJ�np�8:���')&D'	N��05Qe��D�-���y2�3b��
qOJ;i�0��a��#{��b����	�
��xj%*S�d� y�'����#?�����a�����?^t����<B�B?O\��� R�^�#��y��: ,c��q���i,�dY��P����ť}��� �ҵAa!��Y�*M8p��&<�B��#l� X��;�O�X;'_+5h�Y�u�ā;�����' �IuE�]��/L�T)D$���B�@GȐ@F!Զ1��T���Xvs^B�	�# =H�[Sfl�1�GI!��C�I�u�0�Z�j��Fu ����B�I�Y�BZ�L�1]VPZ�
��L6����n�t�4�������D�O�B��&:D��`vC�R�3�E�0#4x{�n%D�`ˆ��{��źS!.!=\=1d*.D���ANY3M�����"�.,��c�/D�D�fEQ�V����%�M=D���&9D���KP���X���d~�A���8D�P@c�H�T��y�'6��="��6D�4��4�,4ZW�Q�B��	8��)D���J5��XH���q_�5�Ri(D�̢7F�-n�ޕ҇�v!D!9⧦��G{����&H���ф�L�pma��H �!�d� !����p�0+�&t&iG�M�!�D"rz����@N���	W���)�'9e��HR�r�K�'�\��M�'�L�1K�>���bSNU�=����O����	:#�$A[���*+Ҡ��b�=�NC�	 P�����%E��a[�H�u:�'(�4����6�!I�,Y�G3X���'��MYg	�6[�ܼ��ۗtK��	�'�u�-��a�� ��Xf �M�'�ў�}�Lʧ=�xah��խg��C䉦�|�$���0�&ܘ3�չcܖC��-J�\Di�o�/,J�p�T�{ĎC�IP���'O��e�v�өkVC�I?d�Pɨ�i�|�|5[6�:K2D��iդ�w����8]��DB�J<D�� <�KDHW5Z�����-ǰ+|x�0"O�|���-�fܚP�ds�$�O��c�X/�0�N�T c@5D��e��#'��%�^@���4D�\Pb��R�P�aՁƴx&���@"3��'�O�A5�L�g\ތ���	�C(l+V�	A�O��̊�˅)H����B�Kg~α�	�'��ђ"�.e���b�۴�k�'5�x����=!&Ҽ2Ra�ꄅʓ	#�L����>fY�!�@�nv���M�#��O~�xqg�\.Zgh�4��;'���"O^��k�	�D��S*YP��2a"O��
*��P�HQ�qh8pӒ�IX�';���i�HyxG*Rj~��SS+��G�!�8���!V6sw
L��	ԶVk�	H��H�r��$�߼8��IAdƦ{-d5B�"O�0�V��H��[�ދA�Fa��O6�Ig��HOv5�-]�M%��c��NZ�\O�ƅ�s;�	���Hv�p�%'`�;2�|��n�Co8�y"a����<���1	n��L�W���K��P�l!��\�$`�(�A0�B� �!򤈥H�J�S���CV ��$�� f!�D�Z,�HZ��N�eF�y+_��}�
�'z$��s�ԇS������
AT�x
�'�vMQ!B�K�֩I��*j���'ZԲ���,U<����� ��p@�'���(ӃK��0ň� �5��'=����R�(I�����9��h�'u�`JN�j{\� �	ߙm�I��'-�� ��=ye���Fo�9Y�ъ�'cd�E!�dzt���S5 \zM��'.��`���h�2�	���%�D��'V��
d����Qsp��5�82
�'�f��7�Q�wZ����3�H	�'���F�=-���p-�3FU�'�2���-T�?��Ѳ ϥ$08��'|jy�E͂8lu �s�f�Ʊ��'q���1H;{l��A��/�"Xa�'���dꂍ�ҥ�P��iv�V^�<�N�'bqN`Q��V6X{t�UGV[�<��A�l�3d��[�D�g.�T�<�b�,* �v��d�>�a ��X�<T�W9����cg�B.�`@T�<���[8|9lL��3T\<!V�
z�<�R!ߏOΖ�;f�Ӛ)�Ȱz���n�<�$��e´j��_�
`�$�Mh�<i��ՠ0�(�!�j����
E�b�<��H��f�2�PH��Nt�e�QEZ^�<qG�ׄW�|���}>�Q��Q�<	�E��d�ag�F�`Gb�<�vJ�P �!	�>&����^�<Q�HDT�
H(�œ81w�� �Fa�<� lJ<
�Δ�UmQ*o Io�V�<����#	*� 	���bx.��{�<��nB:0�� q�럧Q�LDo�v�<��*�C"�c���Ws�@��G�<�G�фJ)4I[�NO �����j�@�<A�J��#�(���F�M���K��|�<9L�3Þ��na ��IHy�<� !� ��X��J��,(���@�<p�P; ����c�~R!1���S�<�r��~�œ1�Q��`��RN�<�d�T8j7գ�L�,lNT��L�<� �)R��G�3�>1F�OB�J@1%"Ot�L\�~�teP�G�u��hR�"O���ƛ�a媄��D���	��"O�p��^=�� �U��%��"O.AB���j�|��a*9.^�F�'�B�'v��'!��'�2�'8��'���6�ٌf�L1�&�ҥK�����'���'8��'��'���'
��'�,�y��:zX*�I��f��]�W�'2�'���'P��'<r�'��'�0���a'��*W�Ʋ��B�'�'�b�'Ir�'H��'���'<�x�2.Q�а{�
�!FDtRd�'���'���'���'��'B��'�f,���ƨ8}t�ۡ��|��!�T�'n�'�"�'���'��'���'���� (`
��"�Y���'���'��'�B�'V��'S��'ߔ�ɂݞ	G�AF&�%M<BH���'���'��'^"�'Q"�'62�'�pr&훥1
��W
®@9��'-�'{r�'<��'�b�'��'#Z��2�5Jd�P��ܦHT-HT�',r�'�2�'2��'\��'��'"&��D��)0*b`� �1k��t�'�r�'���' ��'B�'a��'岴X�j�
�T&$�#x8h�P�'���'Y��'�B�'B�'r��'���J'j��UU�!H��J� �nj��'���'C��'���'�r�j�>�$�O>P�J��4!���$� h��dNUy��'U�)�3?��il�����g�ŠY~������N��I�	W�i>�I¦�P4� �YBԄ���Y�Ds��ɏ�M���1��K�4����,Im��y�����wT�+!�	��t�#��_���b���	Ay���?	愇��t���+�.U[`�ڴ:��<���mp��NCOXb�1���k�:a�t ȴP�4���ݦ������L�Ǜ�0O��s�
���!�����M; 1O�!Ʈ��ha1�9��|��/��4�#FB)�la"�#�'�����$���Ȧ�i��3�)f���Q���3� !�bnU�X���?Q�Y����ɦu����v!�$C�XV:��ןL�Ra����:W�����&"�*r�\�]�?	AB+k��@�_�@]�!c�C��d�<i�S��y���CiɧdŤt�|f����yB�x�������� ߴ����DG fՆI��瘪7�a
��~"�'ƛ6�'>���ǿi2�	�DH���d;��Pう='yF,�U@Ng�~)cPL�	Hy�O���'��'BgU4>�b��!#6L��/��_E�	�Mc���?���?�I~�ifp��H�V�j��V���Hu�T�4�޴����O������E8ǃ h�)��?Ųm(�I)es��*�<�a!]��MZw� �Op�9Pq���O]@{��4��M+���?	��?���|-O� n�;Lͪ��I)aV�0R��5H�\��f��[�L��I��Mӎ�¨>�G�i�<7��O贠D��$b���J�N\%c�h·Y$�6�3?Q�̊�m8p�	d����';,ǩ�^X��rS
ߔ<�$��U�Qs�d�O���Ol���O��D7�S�iF��g%�mQ>�
���=�	��x�I;�M{G"�|
��:���'���"�����(~�B�
�fN�!�LΓ��DK��iz�4�?)2��M��'��J�H� ���"a�)ீ�8�*x���	�#߄��|�Z��������lڐl��M��x��E��p��@�蟸��Oy�Af��m�V��<����nzL��cm�9(*��լV8�'7L�1|��	j��P�II��?��D�٢W�~���._9G4��@�OMJ����K֙_��'!�)�"	k�� y�ɪ+����jA�d���B,��'�D���\��ן��)�Gy��b����W�&2+�Ј�\$��o���D�O�nZA�u��	��M��Ć#\A#u�%)�R-��V�dy��'��M�i5��Od���l�4p���;�̢<�Q�T/?T�H�&� ��²:��	_y��'���'Eb�'�X>I�d' �I��S�r�ꝨI�M#�_"�?9���?�������O�pnz�ea���S�����$���E���\��M[1�it�Ģ>�'�
�B�ҬZ�4�yRˍ�=�٪���!;0t�ӊA,�yb+$�x�PCČ� ���b�ÖO
#�U?Xk��17А��q��Cn|�sfn�
X�Й��K7_^(��v��)L�>���_%��*�� )y{��l�<9�����Q��7s`�x�Ĉ�@;P���/��P򅓁-�zh.=�6�aT�M7���qᆗO!M�S��pI�br�Б"�uU����k�z],Ԃ�.#��0��۲&��A�S�V<<��Ǭ*P�<1�J�1a.u:#�C-A��p�f�r����Z]��n�۟��I/|B������^sxL���_b�� ٴ�?1����O����:/I����٠��s���IR�[5,#�tj�i1r�'H��f.����4��i�O���� l��MܩM0YpE��2.�,+��i����t�I.\�b>}���?7-^�DT���3��!�|����	w���X�pZЦ��M�[?��	�?m��O< 8� �,V ��sk	8�`I3�iF��'G��*W��Sʟ��3��S�=�43Vc��Z�8	𠋂�Cڛ��$ajl6M�O>���O6�IPM�i>i�!
5�xiw�_	fp�����%�M�'��(����O,���1O�۴j
}(`(_ A��ݣ���0J�p�W�iK2�'��[�ilO�)�O �Di97 C=J?`�)1���B��b6k�>����?�W�`��?����?�� x]����?�hMr"��Jp9�%�i��+SN��6��O��D�O���T\�t�OH�D���vɒ��7�TjeP�8�&eq��	럴����	@�㍷j_�y�VN�0*0t���C�>y��-�v�x�����On��On�O9�I����#��&��!&�F
C���9��o���XyR�d/R�'b��'0,:F�{�4ٰ��Lv����C���&���E�I̟���ǟ���[yR�'��h�Oi�����Ӹ2t���p$à;�����ItӼ���O��$�O4���O����Ʀ����\�d�L ߴp��fF�Tf���凁�M��?����$�O� �4�������p���m.Ԝ�T��GV4�RMv���d�O�˓1�� �P?}��ߟ<��P,q�r�Q+�P9
�-�xïO����Ol�͛'��D�|����ς�;D��hV&3_��e�w��&�M���?��K�t����'���'���O��N)OJik���y�{&� bn���?��Z��?yK>ͧ��Ӣ3����k
�p�將	]
(�D7��W�@m�̟@�	�d���?���ٟ$�	."D]S5/ڱGd }�6�Xh%�$��4p��l2���?�+O��8�	�O���D������3M��\󇠞�]�����	,V+4h�4�?����?����?��}{��ipDl`��Wo[�/��mПl�'�>9[���)�Oh���O���fV("�"��V�[�T�>��UFڦ��I�O���4�?1��?�����r�I&Yt,L)�ŗ|e"�z�*� ��x����?I���?q���?I-���y�@� Y���^5\�L��9]�l���	џ�����ɿ<�I�DPs�J��zrh����e:F�����<����?aP��%�?����)�����n�WSd�R��	��ej����X>q�ܴ�?q��?���?�)O��D��t����7lȸ�Q�D�~b����[�E>Vn�ٟp���4��Ƛ��� 1���ߴ�?	�6�J�xUg�C80R7�r���D�i�r�'��Q�<�	�)� �SF����7��
p���6A� �x��f�'S��'�F�f�7�O����OR��!^פ�9U�=o�P1(W�])sP�o�ԟ�'��L�����'��i>7mC�'2U�H�!V�s����`���'aJ�?yor6m�OL�$�O����$��	V`��+V�i}@w�D�!o�d�'���@?%�'��i>���ZHV)Us�`�����$��8��i^��C�vZ��	П����?�����I���4E�� ����DK�ĉ$�� �MB�ߏ�?	J>ͧ�䧜?0�A�5M����.`lf9�f�C�)B���'��'7LD��*�>�-O�����;C)�f�l&�J�7�2�k�>�,O:������ޟ��I�T�D(��M
N][dd҉v ��gF�MS��	�&q���ik"�'C"�'�tꧦ~��YwsJ9@a�$���B�o���d_>=�	ß<�	������4�I>w����e����d`�M�@ŲE;�Z�M[��?9��?I[?M�'�Ҍ^� �|��N�F:D�c�@/8���p�'[���<��Ɵh��џ���� �M��X�^�3hQ�7�i����=��f�'/B�'��'��IٟĐ0nb>�*�݄+�4�*��@f�X�	�<����Ot���O�˓	>|ͣ7X?����+e8y��͋W+��R�bV�p�cٴ�?�)Ob�D�O|��'Z����O����s��<�aX�Y��4sC2
��6M�OF�ĵ<A�c:6{���T�	�?Q�%Ӻ+�,���$0��0�mA$��D�O��d�O��9>O��O$��5���A��|���F��\�(��i�"�'Ţ�S7qӤ���O�$��V�i�O �� l��9�>2�8�AG�z}"�'1V̚��'h��'��4�:�O��Y#�Яug�dI�M968p�c�4nk\ "��io��'��O����'b�'Q֘�ӊ�a��`��ț(q�`vӾ�a��O��d�<�'�䧜?��eE*Sن�Y ��8���)`
T�q����'B�'��ձ��u�<���O:��O���RX�@�?nLh[��8��DR��i�]����`p���?����?�@l�L`h���^�8�B����Z���'�V吓(|ӄ��On�d�O2��O����8d�M���l�z]I#R
8��i�2O\˓�?y���?y-O�|82��+FY,���[?nv�����.J�ڵ&�0�Iߟ�'�4�	ߟ�R$����DQ&H>p��}�Ř�"�Uy��'���'W�ɰp���0�OJ�ͱF���	Ϛ����hǌ�i�O.���O���?���?�PDւ�?�cM�&r2��"��
k�
����ʣOn�	֟�����x�'���#�c0�M)�9��M�t6�DAƞ�2W��m��%�T�I�H��GFݟЧO�1PD���|�S�'ƫ��$��i�r�'+�	�~��I|*���D��5��Qr�b4Dy��G�Gˉ'���'K|��'Gɧ�)� >0I�#��J� �P��)�?	*O�vB����O��OB��Il^���A��L)���4^J�n��l�I$@b�}�	I��C�'�����W��wk���)n�4^��i�ڴ�?Q���?y�'qU�'����3];]b�, �|�>!�U̝?�6-J�v����=��埬Y�(��?,��ct��Af�{1ɞ/�M���?��<��3ҙx��'[b�O(ȰB��!����_G����F�iQ�	������6��'�?a��?�B%�}�z%b�˄�2���!��3^����'0\�k�)2�Iԟ0&��X�I����eуGbU�TX$�&�{Z����O��d+��I�(� T Cgb�9�w�/3K�����r�Iٟ���y�	ٟ��	�l �C�[+��X�Qɉ%O��,��hNٟ��'�b�'\�Z�H�6�Ɉ��� h��g�� ����&��IR���	��`$���I��� %�O��H�}4�y�GƝr���RO�Z}��'��'�剎M��h�K|2�C4ޢM("a)l��)HT�L U�6�'U�'A"�'��y���'��G����	6l4B�����S��l���	hyB)px�������'kY��2� ����b��Bb��G�	ϟT�I�|I:��g�	[
�g֝n��(!�w}L�Z�#���ɖ'+���#gu�(��O��O�P�8A�2E
8L�n0X��դ��!mZ�L�Ɏ[�\��?���� ��aQBQ#�޸���8gf��M� M�+Di���'#��'��G-���O��Ǆ�r�ҹ�C+Y!���V�Ŧ��$���� �'~("}������Q�I.2���0�C��Ô�iR�'2��#g`TO<�D�O��	<`t���TC�.j ~U�@�ĥ6��7�<	�9AxY�S�'
4	vs!h�!Z-��A�nȊ p�"ڦ _D��RF� BJ��5JD�uFn�+�H������_O�'R��Y�'-7xp8
�-�t�	�2J��&��<YgTd�G�\�n�9�D B(w#~����[�d�.�K�b��W8Xt�vaQ9��u�&kP�z5����G"[{Ε1`�P�P��E
���ܩ�W������v/��Q��`+a�)��fj��ƣ�?1�n8,11�ϏPfE�E$U" r�8�c�Xc&��}�jE�UL�.F"�'�@��G�'�b2�ֽs�T6oʦ�2���>v�x��/ɾ/U���U�y�r���nQ<&�J�?��Z�#���a] ~��0S�h"�P[��J�>>� Ⳍdx�A�����*�¨/���c�N�0���9@�R ��t�!���&`��[��
@(V�\�!�D�ݦMz���m�@��Z)&%(�;dk�d�*eD�;��|����IFd���՝"�J���M��z�Pdp����^�|���O��D+�`�t0�D�[�M[RM�8H����|�3��?��<�w�k�����j�����:��K�r�Po$;(ݐ�e�!Y�l%ɔ� к�m�%@�*'Mٻc좡b���z��Z�w���'Q�>��I `�n}�3��;><�=�� �4\��C�	$P�zP��]f>���bD<�aF{�Ok@"=�6��?M�:��¯� 7tP��nT$hS���'p�'ʺ�t��}���'`���yMC���#�,Z�ITN�`���-�Ap+A��l�ҷ#�<gf9���.�d,]����p�2���B���`d���@��a�J�Tlj�Z��i=���D��:N6-�udWk"�X�-�O��!����i>E{�؜_���À��.����O �yhǴ)�h�g#}�.�k�c_����U�����<���ϱ��e�D�O�V@V����'YQ�����?���?��7��O4��w>Y���<a�؃2a�����Cr�q37o�<9Al@��Ŏ�"<��I�-<����L�J����f́�Xb�$�&O,Z���Ս�[�����-X�(�+1'�=�8F�Z�L��XIR�O:��d���ީ�G,r��
�-h!�d��n z��Q�[]$$ȕ��-
~1O���>QWM��}w�V�'<�a� ~ �3�Ƨ'8	�B��<0Z�M����?����t̚�}���O��M��@�A�ib�)"c%R z�3z�)�
�k���!ɀ#s$x��d�C���W^W$�k@�G �����C�����b�'�J�q����)���a�Sr�h2�����H�ȓn��lP��A1wM�C!�^Wn)��i��$�=m�^P�;.����@T$�'a����atӀ�d�Opʧxk܌�x �2�!ǈ'ÜY�eğ,L����?�B(ԋ'^�|��� <�3����	�|r/F=zP+d�8RZT�qDhc�$G��{N�,e 	�d�\��g-�*�ʅ��O��X`@I78�F�q�@�-���cK�����O�b��?}
qB��8����	,i��hd�6D��	_��9Y�LRG����3Od�Gzb�&_z>�!���)P��y�1�N	j@�7�O$���Or���H��2����O��$�O��{<�t:�=�ǯ��s�F�9<%����	p�
�m�ȩ!� ű�ej�#�ރM5޴��+�!<$iE샚bx�ї�� ��Q��d��  �0������T��;qg6�I�*6JDi���t�B�hc�|����?�}&�L��:S��(�H֝L���@$D��j��5�D���)�cc�H[�#?�4�i>�%�L�5�R6kC��
t�щ@Ofd��B�|������
������ �ɳ�u��'=�;�|M�kR=\Tp�ks�Rw �@ %՛�i�c%d�r��yx�P�D�P� .�I�$�M0Đ����6E"�	#cX U���`��ڒ�ĸ a����$2A�aO:�� ��.R>r�U�5�O@���	�t�����n�,��[�T�`�ZB�I�;�2�DvZ�uTQ�J�c����4��9��}��W?E�ɳO4��;��5��xW�_y�������j`��̟��	�|3�12�XqITAS�lR�	&7ǀx��̜N��8F��M�p���O�豱�%)E���ڞ'��y�)�Nb��U�\_�:�(�Tx��I�M#�X�� ��PbF0@�8aRdР(��EC�d1|OLi�3�k]�cL�.ZᎡi�O��oڸv����v A�7���f�[�I���Ihy/�s$7=����|����?�蔌m�h`C��)��H#R�L��?���	e��!-�<ӌ�ѧO�vа��(���'�4����p���L�47��ԤO�m�V	�y����U�V�^@���X|4����J��]�`�H����h�OX�l��H����}�G�۳[�h��%KY �&B�	�����
M�$��ӑA	2����D�A�'�	Ըp�s�ۋ.��ӥr �7��O��D�Oe�q,]]����O���O*@�;hDt�1B���d���#�^�(3�y����M{�	!�����c�(vSv����l^=�<9�&���}&���W���:e\���,��e�0Q�ʕ���f� �)�3�d0n�a1@��(C�ޑhTl2`L!���/z��<�cm��o���J�IP�.h�	��HO�i(�DS*ͼUr%'�#3�v=�f��9>��ah���(w>�D�O��D�O�Q���?y�������3e�>�Q�j�;'��2��!5x��e5ڮ�p�A��0=)u�H�\봑�!�MS`�pTІ~Tmh�S�$oJ���W���L|6d{pȐ?f���r�/Z@� ���'i7-F�����eyR�'�O>�⋠tt�� �#[�6n�bW"O����]��i��BA�i}	w�d��i�Ġ<� -�pg��O����S��ui"4�mʷ��2��$�O��C�O��Da>�{�o�O��O6Lz��T�y9J�L�',��A8��T%(�I3@80��2���ha셨���ZE ���ʉ�R�&񄒭#�$`h�i9
liP`]wM!��T�r �0�dc �I�n�%r_!��ЦA�f�_��J��&&�N���#�Et�	++?�M�۴�?����IG�&(���Y-����)-@������$�O�����O*b��g~�� �w,�i����n��I��N/��ɠ5��#<�Z�#�8��e��A4`b��I��	u�d�h���3��酇U� ��aL
�a��̡U��Т�',�|�g�X��n��'mQ�"t� 	Ó9��<jS�*D�x���z5�ihТ�&�M���?Y��'�CJא�?I���?��ӼS��5)���+�]���
7�'���*��K�����d���+�����)Ǌ�x/��:J�Q
����A"Y���d��U��O7r�����3���	$Eӗb��)>|(�,8��'9t�S�g�
w�X��n�;`݊�"qM�A�B�ɛw��ԓ"��T+4�h�J��3\�tV���J�4�X���
=�(8�rbƳ!%�Xyfſ�����ߟ|��џ�_w�B�'��	��#j ���!�`���X1$�d2���,r,�P�*
7
rN��P�!�9Aj$�R��:l�d|�#͈W�Ȁ{�Q�-�8�UO�.] 4A�B���O����U2N�I���y�t���g�i�r�4�O6��>\�+D.��)q�"O�%hY)_A����(ܐ`���ߦU$�t2BN� �M����?a�߅2bi�D�4c���j��?Y�3�Tk��?јOu��ЍM�Q�����:��P�#�v�ʕ �*fj��Kۆ�p<ᣬZ�l��ٙ����]wh�:���33�ؑI���.	@�#��L�$�`E�/�Ex�e݁�?���x�Ȋ#[��;���2��=x�`���y�iЭ:��A ��T���Tψ��xr�oӤ���O4B���c��^�\���a*���7Z�p�mZ֟��	M�$��8X����~�0��l�8*D
� 4��'#�l�E�	�R���ח6���T>��OàLiGI��!e�8R�K��:o�@�N�g���6U T���T����E���>���[R$щ`~4`[s*ې�����	v�)��|^�U�7�3�TZ�n��[�B�I�B�0��N/i~���H�o:f��Z~�'ڹ������y8 �V/"��u)��}�
���O��	P摈@��O�D�O��4��x����_��`:g�^�'_��d�R�P���)¿sr:Ur2#_Kx�c>�1��|�d@+&�v�T
�E���d$��d��,cC�K�||�Z�&Q�L*Z7�2�?)%>On�LL�X�Ȱ{s�2G1�Xk�L�I3E1����|R��G���!���\��(�C����yr,�2/�H�t 	�ez6E��J����m�����|���wl9m��(|*��l�8p��g�)���'��'

֝������|��&�tv�%����[���y5�JC0Ȁ��WY�ek�@����%ET�E�0\ ���|<�%k[�=�n�ꧧ[�W�"!�w��8aA�t��Q��� Re��+�q��TR5�Y���u�"O��Q����x=�u �D�8\@���j�y�DI駺i��'O��H%��_&<4k�`.u�8����'b��$B�'�iDi���!q�_7e��P��AsӨh8�I sV��a����Z�G�'��ȥ�Ww�� �I*n���g��<Z=`	&CP�2?S�fO�lŤH2�V�ZS���=IB+V��I<�`��;pE�cM�9���"k�E�<ٗ��d��p�f�Y:M�fq�6�C<!`�i���S��<�1�E�E4�A�|��ٞI!�7��O���|B�B��?�YMI����/���87��:l���Oʑ��,�D�!8 c�8,J��1�Q����^>=p�M� @��������t�
��,}�B-�X�f`�%�p��n��8����IR��ӿ�>Y��nݶ`.Vu�A"��r�>�t���0J>��m��.��I�C��Jش5X��X�<i5�H��t!��ޞZ?2�:�fN��hO��Q�'�(�6!�����C�I(I�pD1ҭr�"���O��D�!J^��P��O����O��4�4�I��	�Y#�]*�ߡU_��Fφ@ܛ�$9vb��"#Ԝ;66b>QN�x�0j����jQ��<������2�B����1/�(����E�*a��(sM@���iξH�$H�w�谚vϏ�F=�̀a�
2�LM� #n�V�mZΟ���LCǟ�>��?y�!�^�J ���=V�\�pa�,��xG�6� H���<qN~A�a�����_|�'"���'��I�:�
�0��(�¥z �
�Ŏ���Y�=� ]�I������D�Xw��'�".��Q��A(��T�ZAj��	�u�2�˄l[��`�H��vK@��T�>�tD��!;r��t�ҫjdڀ�$ �,�ଳ2�_�G���Հ��zg���qk�#+v�)�W��p�	�+v4�pU�Q�z�����@H-
I��:���O$��H˦��sy2�'I�O�e�DI��1��X� ��m?8 �V6O���$��R�� 2\�y����pKZ�O��mZ��M�-OtM�v��6��O �� ��J�
�6i�)�739���OR��F�O<��l>�3 �Y sl<@�e�/P�m�"��0J�:]�P�gOO8a����3g/���AC֦*TH���$b�� M>Ah�Z�$3/��� Dh��h�M5h�qO:���'��'�Y���ƻ��]1$j$[��'H$Y3'G�PT�L���JO��*�'��7�ij@�0���}Sb@ H,[R�O�� �W즍�	Ɵ�OV�$1 �'D2(���4i����&@�::Xy���'����}x� %�N�(�U(�O��N����Xm"��D)ʹǦ��-ٺ��DIFM�kV:\�fm{@�>H��ET���R��$=��!&b�$/*�8B���4ªē��>91�Fԟ��O>���G\�i�1p��nGʴ�`�<	G*LY�I�CC��6i@Z�������/}ͻr!�A���� �ɱ{��n�៘�	���t��;������l�	���<���1t S��U�eJ �up�O�gέ�7�O���QF��A�1��'?����g��C4'ټ>]�ݪ�.�M�u���}�ɋ�dP�K9J?9�!�r|��W�lE�fI�o_}J��2Vz`b�`j�A�Oq��'Ԧ	��K>/@AQb��<�X{�'z����:m�z�[�jF\� a�OdGz�O��'*��!0�Ό�Xj��|�2]ar]�1R��(��'�2�'�b�n������Lϧ]�,H(���>�uJ�� 	!e$(0���p?VlsFQ�0��p�O��Od-�B�kaD���$E+(�9�ਟaQ4 ���=� S���zd���hO���+�p�l��
�Y�0���S;H���k�.H$�P�	����?I�a�b��+ő;���E��T�<�l�1H�<ࣴOLy��T
dZ̓{��'��	T�Xl��4�?I�31��C�AX+]}T�H$Β1�HPI��?1B���?A����ԥU0�hHqw�<}�D2@��(�L�JlV��2�F��p<��$�*mdhh��!��@��J^�*�3ŭ�fiyp&��X���$�
d"�|d�'T?T�c�� J�v�Ɗ��yާEz,�!+G�����E�x��aӲ%xf�R�h��Cҧ�6ۊ�c0;�dJ�n���o������n����<c�cO
��u �A�L���i��R�e:B�'
z-���Ȅv��ek��B�8�	� �~�/�8l�� �Z�xh�N����U�>��?h��}diR�[�t$ɴ͍��u�nT�Z3�Oa*j���4tӲ��T����I�tȦ��Olb��?��!G�R�J�r�I�>r�w�%D��1� =AY%��K��> )t, O�Ez¤R�dv�mb��'�лJZ�Y(7��O����O�A�5�����O��D�O��E�p~��xg��nfH�H��.w���
���A���u��3���$�%�S[�	+��b�3Ɣ8qn�Ac�#,��=M�<8�j��M�.i����1�h�O集bP��y�&��,t�J���&@�3��5c0�O(P�s�����qȰչU��_J��G�T*a Ն�S�? 0�0)�5?�tZ6�/G2h�R�����4�R�O���ɮZ�"��c��03�Q�d΋9dTD�Q�
�On���O��ċ�����?��O�N�NW��jm�D��.����9Y�U���Rk �}�(�,�џ�ڕ�NX0| �b�E%�ػ�f�3���6�ģ��R`ĥ|	�nZ�� Dqw0�mNQj�-��i˒�2�%B#�-��b�O0m���$N� 9% �&460���"�*B䉺�B�yG�X�yE�E��J�%W&�c���4��x��y��i�r�'꒑�U酥@H,9) �^ad�'�'�B�K, k��'��	M�vо�C3`RSn�i���U�]-j̲���0�*I��H^�F�����(��3��$G�9C�Za� R��Ms��L;���c��3>�!"w%38���2	.HK�{���?��xbE�T #���tH�SĊт�y�'S�`�)�B>��o�1�x�l�f`�R`��h�"!Qʶ��H&�d�<��mΟ���}�t�� D9rɎ�H�L[�)�
\��$�=�r�'��}Ƀc�f+򍰐ώ�X:j�R�h�~*��Ak�=f�L�Y��Ͼ�J�>�A
̆}	�5Qe�]+h�Ԩ$*���u� Q�zQDE��O��|�`J�WN2͈�B�@�J�`H�x�%�O�b��?�U��)RG�� b*\&b����1E;D��QA�:)e��#`����H�`��&O*�Fzb������qwj�	l�i�M��F�6��O���OP���K]�Rz���O���O�-�&E)���]r���o��(�*P�B�\�Ty �V&�[�.��P�/�SN��0�ܢ�O#RpH!clC4#�t�j�6Y���6!�.	�(@���έ"���Ok^ݩe��ݼ�'U�jMSE�&Z���ѵ���'�����S�g�I�<� �p�A�h���y�Z7�B�	*jX�0�x���x��SR��z���M�I�\抴�D�ռ�~�{�㟢,3�5(j1(�V����p�Iǟ��\w�R�'��I��?c���ǂjbb�� e�<HA>��v�X�P�,�t��4�q��=�AJ�iӀOӴr���TH�2pR^����64��k�N�{���CI7�&�Ҁ�,F�R�t�vK�44�x���ԕ(����%�W��D9�O$xr��@�&�O�VRD�a"O$��BB��j�4Cǖ8M��`U�馹%�`)���M#���?�w���E۳��6x� ��A��?y��C2e0��?I�OWt�'�]�8�aL'B�TdE�.���G�aH�����ªQ�џ�ʥ��UXZ���&�=��ݛ�M� HZ,�_`���0��t�m���1B �:��]��d^��Co���X_̖�X@�56��C�=t�j%B����\6��d��=�C�I��M�e�M�Gw���c$L��s��+���8�����'L哴T�F��ɟ(�p'4}+��R���Dz��	ҟ �u�G�Ar�!{�#���Z�8E 0���|�g�ʟX�l, ���9P�>$� n����G�8�I��:]����0L�9�0֝4C����q>u�&���@�rU#%/V7D�$�t`:}2*^��?	F�i՜#}���cSN\��_ n��[�/ٚI�R���m8�'łnL2�5����x��	&�HOB`�v����(�Ǖ��@��F榝���h�	�� u��B�ɟ�����i�5����>@҅����=�(�ŋ�8Z�4=��"/Uܛ�l�;_��0�|
K<��W�����SFUq���3*�ţ�b_�\�6}��Y\����5���OR�����y�L�6Q4�("T�	�(�[�"Y7R%1O&�[���� �L�0�LLh<���tNI�Dl���I��t��B<T�hz�銙_|��'W:"=�'��l4.�A���kLX�9�����M��d���r���H�d`�3j���>\�ȓ`��s@�M�@ƅ�i�O��4����I�*0L�H-C���5lO����:�չ�h��9-$l��H�&1%��ȓCe�AZB倊g�
��!חanZх�t��S�^� ���$�9C� �ȓ�	�!��I�d,�!�0l�q�ȓ�(�hCgB�2��d��	����ȓ)fР�#F�R�<uC��7vl��W�ؑ\7�d�a��	�����O��`&��� ��Q2��ǫ&|��ȓM�t�͐h�ޡY%��H:��(����	������V��ȓW��$�7N�`�.ݭ�bJ@Q�d"O`y�Ô,j�T�J�>6����"O�I��F׸wp,L��N
3�0Q"O� �=��![�n���U�,
��"O@R��C3"����m�)z0�Ik6"O^pK�F�% �P��N?��3�"O�A��_�2�P�s�D)|'�{�"On�0�T�D�9���>&�{�"O�)�A.�6jxxKD
��'��W"O�<z�� g�D��"J�8?V��"O~�s��Q�	�x|�Q# �4��"O40�"W�6RQQ!H�5��l��"OƤ�#�(b����[�#)V��P"O��pk�Z�©��eN�H'2s1"O�Qi䫊�a0x�Z��W�V�r��%"O\���͔@�dXb��D�y�|5�'"OR�X5Fݛ&�Y�p�Jy�"O(�t	� .b��-����IP�'k����ib�r���r�E ֩p惡C�'�2y�X����ǱW��	��$��%��#}��폜`B� PBD0ެBD�D��p=1�� �jRNXA`�W�fa.h���397M�+���G�&�.i���5�M#V��!2�Ӻoz��	$s��@�&��F�z���(�GR�A0��z��~a��a"�Y9i����Əß
�V�b���O4�<���_�o�;k@�R&��Xr�l�Gx�����3Μ�!t ^�3^����a�4��խ�:���i��X�'b�4�7��31��G�Ėp�>y�'�P�B㋬B�μ"f����h��}Bk�	jZ�(D��o2
$8���!�ē{(��z��O-=��s ݽf�q�����E��ˊ�x���i�i�;���>����$��S�<��Q�B��_ZP��G�~���q���n�ay��c�C���0\�t9�6���;~���ù����e��bp/�k�����M �QP�E1|O�E����	E����1���8����u��sT$�\֮�ـ�\�t�����%�"-0���Vˁ)i�2O`����ɢϷ@��8��KG&������["`R�-���z�j��[`>$Dy�S�Sn�Y&hB�mz��x�b����DI�n�i�p/�iy���7)P>��d�Mw�y����=<4�G@Y�.X��S�f���a�@I�#bk`��m�J�x��a �!�lj��d�<i5B�ub����"�����R��8�T/^��`��k�8;*2���iIHǦW�15h�4�>\O�'#��:SQ0-yc �D��L� ����|2)�,S�6�a��D���a+�p�ȲC�=M� �>�u�i� ��� ��H3�Ys�#W��u���>1@G�2s��}k��H�R�T�Șt�'#�b���%f0�������(O��C�K�&z�]�$�>1�8��Nt:40h�ɥ
������]nԑC��d��s�R�{V�Z�K:�i
7J4NN6�9�"ř'�亠���0�E��������|B��A���+u څO6x�A'�,dјm��'���2GG�{���)t Ɖ W��k�-3�nZ�6��'=���`�
t큽�5v�̿D�Dб=��ٸV��
+����� [W�RemI�?	�,c4fܭs`9� $�19s���D��<I5��O�2�7�J�la0n�M�g}�K �.	�9�R�Lf�xe�6�� ��'���p2��A�%Z��Z5s�q������)�D{�C�Vuh�ku�M�Y;��vA��W��hbQ��7����T��c#�D�2�@�C�oݻ$�4�Ku��v2H(��TyBC#��OּI���uǡ�,&ю�+#+�QW��r�>Y�j�`�8�O6Aa��O�}�<���@�'�,a�V�'�7M�51����]����YشT�'����D�0}Vu�6�/e~���ɜW<H�����D�n)r�-T�H�MX/��(��1�O"�BgҊ8	$牭97���~
��QZ}�c�	J�z��N'�����\��O���4�׆S��2!f��sς\��y�M�>Er>P�`��G�.�M#�i͇�X��"	�0u�����Z�'�&�ڣmӪ ����;d6e�` QΠ<�2�y�n�A"iC��?��O�d��r�F�-��H��
 �2�W��?�aKQ6^� �w ��q�edD�X�d�1��&��n2��JY�u�O��x��!_�Ee&��%`ʿ��=���ܤ2Mo$�Zqs�(����0́��8�ɣ*m� �e�[�KS�I>鸸[�W>9r�K����¬f�q��nӾ2s���hO=?ܱOr1�W�K3�����6������~nZO�4���'�;z�2��/ԶF 	�41���zC�O�b9���R� a�$hD~��L��pSF��~��A�f� �~x\�ӈ�Aԧ HXl�7���E)�T?A��zI��Ğ9,&�u!2$�\����`�s2/J�<���
�"�D��S�gs�����q�	L��'׈!*��܌E�2�h!��	:ݐ%DB2��A�;� F�a��.����6�0Gt��i��M��VY�c�'�<�J!��4�'�t�'�h���ɘ�"������T T!�#�j�n4�~r�'���f��f�0ErnC�d�d���O���9k�C4ag6H"@�O�F����u�<��&F_
D��(�抌�hO�-��l�ᤈӓ
�{�j��&�ORm�vR;jD�5H��2�@"O�0R��-UrU�D��! 趸���i�*غ�Z�
�9 �67���!��t�O��A�'�w��{4c
�9�H�hr!T��f�`�'5�Y;dZ�8X q�mȫ��ɓSkk�LA�'�^�+ .>�6-Q�$r���}4�1�W�F�:�"���茜����䜼[S��CK��6�ѧHA>L�I��G�(2�b��K��W�h����g�9=
���4�	�wU^<@��(/&����[�UV�lګGb��Ms�x)شU8�T�'�\ڝ'+��ə4����j��7 p +$'�O���;EڮN-�hx�������0J����q�Ĥq5�E�5B�'c�D�U̓�'���d�R�k!F%J넛fٺ@چ�:,OB�H�
�)wM�t����@X�uD�<�X�Y�!�";� �W��S~��<�K<��X�x�,O=6�v�'��'_5��b��:�P$����1OP%�� �1SL�y�Q�
V���A��=g8m��O���.�j��Fϛ��>�Ԣ��[�L=�O�9��� �Pʺ'���c�D���qkߦL�ƀ��Ș!h�B��<1�lȐg<�Il��ƛ�j�0?�%��O�6_^@ɶE�)���I~$�k���,{P��d�bu���CO܎/��<�L0 ��O� EzJ|�c���q���S�Еu깘���
��<Q���P�긚���*;&(8"1Ȅ%K*FA��ү�	�dYI�'KJ�'�,�h�I� ��� S����Nў1y����1��@��Ē8R�q�n�7
��ˇ�X?_�'���H��-;��)H����$@��߮��E�̈Kܴ�u��{>�(@/�K*����'��5bgЬ)0���6n��̓9�N]!rݺB#��S{����?�O�y 0�Ӽ N����R�7pM`Qd��<	�,�9nQ({��dX���� X�ʌ�b�@�_�����:K���i��H6��ΑY� ��>q��֯�ͭ;U֐���Q�j��`Ù�{�ĵ	#mR~�!�D%n�<�a��*�X���*�\�P���'��$�&�M��M5NHr=�g�iԘ��S�T�[�|���wD�)%��P"���p=Qe�O�x���H�["��͗T�Ԉ��C��c�'#H}J#BR�hP��:���Oq��'�ZL��5!�F|�p���z�N����D�[ZM�� U�O�n�1lH[�6J�c%�R\j�'Ȗ�a�T��`�뉁u��Ď=+�}*&%�:Z���	��ٱV�(?�|��LSh�t1���Jcx PbO�@�`1 �g��s^���I�
�x!���ö
�hڃꁟ-Q6�Ⴃ�M��AQ?�P<�-�vT`T��ES�M_����O��n�|a�����Ѫԉ��x-�#?)��,e�-�R�^�%O��i�e����FdM	a�"����R�h��,L)�F��*Z�A���~�&"�9O��Y�O&?����ɩ-���I�U���U� <M�Nl�,_�m�ꭊ�/�~jv�O��'�Ji�[	��a栀('rܬƦ��%�d-x1pVL�c�����
M�t��W ��5L�^�����,�񟀙����d�O����|7o�;����!�Y O"�@���܋��Em�e<�%�I Mр�G��*B|4�"i�KZ4��<�&aq?��,"�V���?]Ц!��(@p	Y��Ĳp�RD ��1d�!Ѩ�|�,	�&U$o+�\�`�T�#laӜ���+₨kD �3���(��OX@U3B�|�oڭ����2kb��i�{�b��Ti��E&��T
[���E"W }2�OC	,m�����O��:}px�1C�٣>h���m��\�ި��W?s��<8珞��p=��A����G\�s�x�K�M�E�d�аl����>�n�O���):����&S�6���$�'�A;C:m�����*��E��Ņ'����6��>�K��'������+o���I�eE?PJ�b�K3���#����D~R��r����� _)����+�M�-&DƉ)t��$>���F���<!�d��<�7Ǒ.t�}�%8b�֨+p��D�|~i�1�ߤUwrHp��֫M���'~&����t4^lp3D#~?����{�$���$?*ց)����ܝYnD�4Q b�&B�P!����Vd���Ё�D�(A��"�4���
Q*ɚ@�h�K����fj��])Z�Oj�����ƯP�� ��c����J�G�w�Z����ϦE�e�'"��FV�wW�#�>D�|5BI�\���i�`�dC<x�( ʑ�b�\c4�7ώ幡L&B!����
�q���zr$�-%�2�@@1N_ ���Ai|��&�5�bTp�'�� H<����[0�(��[Z�`���Nl}B!�@����6�� �F�����������	~�;3
�5����X�v�������
C��}:V��(C i���z�~]Ze@�G�= m��]q1��7� :E��(���,Q�@�|�PP�$|��M>ь��nQ�HYB O�.Y;S��^����t��p�w�������#|he �,]�x훚'� ��D�7<�L��n�? �����ڕ^�f����%6͡��XY��c�u8 ��҆y����X�(mz�ƅ���,`f��(<����e�@�!6<S�Jۨ�11�G�>)bj]j��(
�N�K6���<AԩV`
��"U�D�$3z�(fbMg�'�05Z��ȏ\�rq%�, 1��"ٴ����#F�b��E�(��6`D~��N+q��w�ɲ��m������`/^�=�Q�,�=���U*L�v�\,_��9	v
�h����NH�_��y�a��)*���e��5n�&�\�Ò;���w����>����`��M;G��aa�,͐��=�1�I+wm�	��MÐ�l?���!�a�@K��$i� �kF<p� �'4d�I�4@��	(0�I:�����]Cw���G{ꑳ��S3>�����σ}u�Xs�	}B�U�����uۡI�^�R5�[�y���?~0���Z9ni e����'4��ٴMZa����8lX��F:��HA�ME�<���Ӎ,����cj�9|S�"�B�<Y�BM{<��V����TT����<�E�xl$�pmߵN��[�@|�<�V B�F�٤$�/E�>أg�t�<a� V��C�@�ּ�Q��X�<����6SS����Z�m���CF��P�<�EB@���	�+�+)M%����F�<�`�O����@�Z/.A���L�<�Q�ִBYv�+�^�4�4�#���N�<i��<>���Rq`E,$��L�I�L�<Y�A�}�@�$�B�+v��
P+�L�<9��_�Z�~�1  Ar���B�.@�<��@�y�lk������%�@�<1Q�T�I���T�K�pE p�e�x�<1 �Y-�6m�q���"5��*@h�|�<�gH"9Ѐ�É̴y�h�7��|�<���b��Y� #[%Mײ\�A�{�<i�D\`x)�"�aTcu�<��#F8g
�E��e�&M)F)#'�Lh�<�SF�f~��,�l�ic6���<���Ӌ.^�p� G�*Խ�� x�<Q�'�c��(��N�U�q�6/�r�<��i�f� ��	8�N$A��Bd�<�4��c�r���3è�ô��^�<11��{��9�K��+ni+��\\�<�R�EX� �ޤ~%���t �Q�<���p-S4��Ȉ�2p��J�<���^�IJ��΃^�ڔږ	�E�<�@͖�]�V|�(ߌ�r��}�<��şj��A�T��!��rr)O�<�a@�b�+UC�/;�!� nW_�<�n�h�:�.]�C�,�
q�E�<!V(�Z{�����_�&$B� ��<Y�*Ճ*E�P�WKN�<yS`DDV�<Q��RiC�`X�� C�0�3�X�<��@��K|���Bţ~���1dQ�<��iݏQN��5�R"
2@DL�I�<eT�{~��:L]� ��KI�@�<��_4]� b%I�!�&T��Ma�<� �Z2e��i�"Ų��t�S�<��gԋz� ��MXqj�R���W�<qA�t����gɊ�����G�h�<Yq'ٜK�I���*fR~9��YP�<y���Q^T��̚&oN�Y�!UJ�<I'�F�PQ�<zƅ��#w)WG�<���K�vh�g�q�Y��G�<9#%O)zKj��DJ�XV���N�C�<��D�<WG�Գ1��|�6�:@��Z�<���(aŘQPǁ%D,�2UZ�<)RA�0b��A3��"Ik�PZ��Ok�<��؜h<TȰ�a�RW:����i�<� 왋S�2!|���%�H'adqK�"OP����7�4t�F�Y;?I!�A"O
a��E����k��RD�Ě�"O���`%�n�pl�1.	jA�AF"OX��7�ۘu�Y�OI�\L�A"O"p��0*���
�D�:Ozs'"O
� �9)YBMs�n��{�d��"O&���G�'�v��썖(H�m0#"O�1B��3���+��r"OZKA�-iɰ��U	5i��m��"O 1����\�b�R�G�hD��0"Oܡ	g#
.6ۢ�#@)� A�Up1"O�y���^�:�Y��ꂞm֚�8C"O��Z��0$���(� dl�K�"O����/f�F����]�j pِF"O�*�g��>,.�kC��~I���"O�͠g�Y��Jm{�c��%"��A"OX�2�ʯYL�ć>3�m�E"O���A��JQ�"�C�3��S�"O%�E%�8i'�dYs��G�ыR"O���2f��@ڢI�����"Ot�gDȟM�Te�!��5P�t,��"O`��H͠>y���'@((��"O�Q��Ny�= ��;�"O��x�oR.]�|����E�!�"O���J@�l;�qsE�� g���"O�E��!q�2|`��R�ZP0i"O�����-�Y�aW'U[Ta$"O��v�g<@׉ܨ>��0�"O�x��
?N,�akĀ0��a"O�L:S��|928��(E�b1�C"O�{v#ɏ����	��(�q�>9�OP�=�O�����\$|�8Lh��3^��(q�'xx����p�Ǆ��Na��'�X� gܰ`b�Rg%U�y"�����D�	{
��'&z��5��m�]j� �牥5�\�F���	V���GcڹD����%�pJp�y�h٠P��y�r�(Z��
O�E)���-R��x����<�&�'�|��=!F�s�� ���ns`�J�/O@�<�$B��p%�JY�c0���K~�'.�x��Oߪ�)���MsPʷ�	��y"͆���4a�8AXR�)�^��y���[fL�0ǂ�
4�X�x'�L��yr�׊VEZ!�Ɇ�3�8ȶ�Q�y2��Eh2��$�E�z�J���kH��y��^Z�6���V����%���0?AGꪟ\���@��P!B�R�YӐLYD�(D���v zxh�GIcN���'D��� ��5��{��@�>c0i�2�9D�, c`��8�l��,
8q 5I6D�<"���a����p��I,>�
�D4D� S�.��-Ԏ9i�DX)t���qh=D�����T��Kw��4]>|�`*:D��x�/�${�9�D� �����7D�����p�EI�96p�2s��7XC䉭kN�:�i�"o:�I�5$�@C�I�&�Zњ��W
oDj��#�<;>C�	�R��`�V�6un���낀X�(C�I��"p��.~�̃��u��C��$P^��u)��z����gH?�C䉋g���ļ��QMn	�"O���f��	1C�h8�A�;�*q!r"OlTq��})H,j�O��"����"O� :!���E�z�p�wtҙX"O� H�@���6�qNS$&eZxi@"O�q3�LOK��k��� }`hY��"Of��'I�"p0ʡ�ۺcN�R7"O�,�(C"��i����|c$��a"O��3�[ �2�G
H�x�U"OL�{�B ���m�����1q"O* �BH�*�� .��F��p��'~��ɌF��hj�� �:Ĵ �#✠M!!�dҢ+((�W��/��y��b�
a!���+J�4T1�m&D�2�b^�!��<O��d�و��=�!�I?N�
��A;+�ʄ��/���~�R���6�Еm�@1�`� ��m(5Nf��D{���ҬL�8�i�`D|:j��p�U�@|�y2�I�*��ػt#�]�J��٫�.B䉿a�([��N�1`A����B䉊ux8Y����$ms��sHB�I�X�zl�!fS�Y���(E���'�0r���D*�)� @� ݄����7%p��dĄ@X�d�'az	@r��N��a0�̒Xx��#@!*D� �� y��M㔌f�x8�H'O&#=���U6�H��甧ywl����H�<�J]dhJ��'��d�����<��Jbh0��(��5����~�<��^�8o�0r�KйD�޸2Q�D�<�2��ZP�X�CɺRGli� #�C�<���ԡ�n@�C�рl����p'I�<A�J��u�j�.ظ
-kSG�E�<�w@NvE	�$��O�Αx�DD�<�6�P#��q��*?��P"~�<!��/N�)�$F�38༱c@��y�<y���5(���#�&,H~�P�1�^�<�j�w���ʠ�ڤ�`����\�<�$Z
x�41�d��F�ā�F�X�<٧d{�5�W�ՕU<
7��^�<!`��rfl��_7S� :���W�<��̆�^5�1� �Ҍ2~<0J���wx��Fx⤓�+�(�`�����k_�y�jD$̎��BH� {�X��o� ��&�O�$X�!�;*�"����.y�ĩ�"O��U�S>��H��O�*tđpc"O�驑�I~]��
�/5�3�"O���c��J�G���v�DM�эQ�<a�����p@� �z@�ӭAu}B�)ҧ;s�q���'Kp	!��>�Ҕ�ȓOb�a�!�ֈS��<*/�4��m�D�B�L��W���jy�8��o�	@]1g�V��`�R��!��k�,i��RvO©(��M�#s�Ʌ�#��\@AH�&U�����K>��(��#(:=��_�Iֲ�I�	�;p���ȓD� 5�G��`�\A��m�7������`��a��>T[2dԳ3̭��hO�>�ӫ�#r���B�v�%��-D��p-��X1\qE'�\��j׬)�	C���(�`O�"�6-!�N�P��H1�%D����²y�y�n�.����u #D��h�݊g�L��`��
 ��{��O�dF����0s�^i*4-�fƌ�T[}!���$0qZY;�e 9� ��e�_�ew��)�8�4��I�#[<���l�K��!���D��+�v�93�	<U�T���W�zj!��U�<���v�>�` �.k�!�� >�8��/^��@>c���A"O�t(S���4��d��ۺ
X*P�Ib�O���x�E���dI�K��}��Q��'�,��6,ҫnne��B��v���H�O�IU���':6� ���!A���AA�Хt����'���"��#
�E���b�DQÆ"O� 9�f7Q�}80A-)횔z��'қVR��JTm�!����u���0���Y�� ��O�� ��ηr��M+�/^�+�^��s�+D�,9��ړ�X��%��	o���C�+D�$�R�N>Wv̡���Y�K�(�9�O(D�(#��N�?��� V�3�đÖh$D�L	bb̎wpl�@N�)g�VEP&H%D�0R�-<��Wd\�R��@�C%D���B
�Ф�P�ſ	����k$D�H2�G�Tm�C<<��@Q��%D�x���G6���I���Z!t����(D��� ��<�h��g��%u7nmq�3D����.׍>f�e	B���E�f-+/D���fI�'��-2pk�X�|��+D�����0"z$��.�{̀	0��3D�4�0bWx9 )R1�F6Bx��">D�0��gS�h��С�	��{�0�Zg�/D�t����<���b��q���鄢+D�d��K��%a�a�� W��0U�7D�H���2u.�`���	e͢d�g�5D�l���1$n$��&2,�B3D���$ɎVD���b _��u�2D�p ƅ�	!�Y�!��3m
�6�1D��13�ܔ9X�9�Mɐ+�q0K"D��(2.5��9�G�9D �i��( D��B��,i�e���=�$@�$D��"��!?����)�=Y�^�p�4D�����W
h�Yw���E="���B4D��j��՚��M�"I�%dL���4D����X4%��"
�+,�xh�f1D�8���3���p�_�DaB4ˇ�/D��0&�92��Ԉ�mS����(D������?7�Hd@񥚹O�`S�&D�����F$Ԉ�@�j��M��("D�pCJ��#��FHL�Ռ���c D�)��Y�~ �w��>o�T!Ul>D�ؙ�ߛ ,D� $�s3T\T�;D�XC �[�T��@���$�h�S/D��Q1L�	zR]�ȉ3H�l ׌-D��9Ƅ�Qh�<�rN��8W��HÂ-D�Hv(H�A
�!�@`��JD�Q*ch!D�|����q[�Q�G*bv���"3D�T�$�үt/�	���+TM4u���=D����hXu*����-oQ�ՠ=D�����ː\|��#P ƌS��0�-D���2�W�7]�Q%5(��.+D���g��P��P;�$A%E"�!�)*D�����.�zMB�-_���p!�:D�pq�/�k𶬜�R+��C�i7D��נ���*u!b�� fz�s��/D���C&�� �NM�N��&J@�-.D�dr�`�=�8Y#1��a���*p*O�e��� Ǻ��D#�a� "O`=��@� i�]�^(p "O&�C + u���C���b��Q3"O�����V:�	P'�e֎��"O깺�jB#U���LK���}2�"Ol�����#'����f��N��"O� �� �K���&�Ώe���C "Ox��ԏY/�,��F�p��,!0"O��2"�I�j�L����B��i��"O�ݡU�_�%2��h��5"O�葇�(n�h���CW�|\ൠ"Ot��AV,�[�cGPC�9�f"Op��D��֕�$-UBE�U"O��3�fG4�ܴq6��wQ�K�"OP\��)OEzj;�Bhcd��"OJ�	nґAS! ��H�-��"O���t(�7n8P�xU"�d4�A�"O��f�>T%��*q��P@�3 "O�̻��V-a򦸱��ם�P�"Or�yV)_j�J��E�L�h��"O(��˓��H��ջ��yp"Oؐ3h��t����_)u���{�"O����E��]̂0%Oj�0Lq�"O���U�QOPX�
�k�b�6"OF,C�h�$
0�UJs�Y1#+�Ř�"O�"��C��"찐a�X��!"O%���չ"�@˳n�:0���"Od�"��ҕ90�a��ͯ*�| �"O&���@*_*�x E/�bD�`W"Ozػ��H�z\<��a`��[�ˀ"O�]{b!��W�0{���9����v"O"D�r�ڈ2u��YU/�"7��q�"OB�R���hU "�F,т�9�"O�Sm�r�y���:��B�"O�l���Iq�q�A�,��) c"O�{R%]`���J�5VMf-�3"O2!�87Y�)�tD6�� "O,h+�E]��V�ـ�G30l�U"OLp���yu�-@j=���"OH��R�ce *2	@�f	H���"O��y!�»NΞD2�F��@�0"O H���3.D���(�_�"O:���:�ѳGʋyP*MX"O�a�֮�5f�*�0G��HP�ĩB"O��c���!���D�C�.�"O�J��'n1��1�D�?O���!�"ON�aLO+tT�Q�V���5t<�y�"O�� �N�.2�0��NM�k���"O�(�5�Dz�	d� ;u?�P��"Oa{TO�v�䁒B�@
��ȡ"O�E�& P�y��xL ؐ�"O�@_��(��N[Z��$��Y�y2jZ��R|���L�P\�P�% 5�y�G�?�n�)�hAh�%zD�"�B�ɺQ�N�KDGξzU��H;dC�	&j��$)��/:�����oI<axC�,�0����B�e��LL�)��B�i�D��y?6�*�J�Xg��"O��Z �-��!��	"|s� JG"O�H��bSHuS�B��8�(�"O��2c$\�n�θY��E}�@��"O��C��I�1��� /�%��"O���5��r4 �1�X=b��u#'"OJ��a��x���1�}���B�"O�l+��u�h1c�kY�y����"O��Q1���.rH�rFj�(��R"Ob��0�F�O�,yX@�˶>q��z�"O��I� �x46O��tM��"Ox	eЙO}tY� �(��A"O )�Ǳ`��"q�/�}pB"O� ��B�O)M�d�1(�,G}��a�"O�z�#ͭaB�IUf��NeJ��"O�y���i�^]��K�>\Gf�C�"O~��͉:���EkL��Hñ"ODȶ�W�W���+t��4���X�"O ��cS&M(���.�V̒1"O���0�VJ����.a9��{�"OX	��G��DP�ю�;)���"O��y� �`��� %@�|
@"OPѰEI�&Y	Da� b���j�"OFPU�fD̬�c��)�"�`s"Odԉ��ofPJ��]/xp�i�"O�	���E?���z�)��9r1A�"O�"
����3�	 P\��"O�Q��  5sJ:U��L���t���"OR�9�*�~̞�1M�;\���s"O<�f��!����mX�+�"O�ɉ�k�5d<������p��&"Oh�2���
m�83��r��,`�"O��Sț�G��+�l̓Sb>���"O��
@��u����P�+OG"O��0�ǰ����c׈v���"OdtJT�J2=h�@��3��}�B"O�y*�>tT�`»\�� �"O����Ǒ�m����	#���Rp"O4���M�C�Ui�IVB7���"OTX�b��A�*��e˵���"O*�r�!D�'�Z��+�A(�4�V"O  U'�3���&HU0f}P4�3"O�GL/L��2��+\ldH��"O����[f s�#��W��v"O�9ꗋ���4�&�9 ;h��"O>�[�AC�- !��/�V��"O�$��,*L�r�[4/�� c��b�"O�(���V�qR�)�3�,dG`W"OH��7��#k�0;3����A`�"O�u�r�� b���` ��pP�"O�}SB�ŉ+k��Z��I�p!�$�%#t69h��ؙ;S�89 �H�L!���I+�e����n0�"�"OT�z�gF�x���6���1��`"O(�7Lɛ!�pŉP/-g����"O��s��̠�=��N+�2xJf"O����1X^Y�'.Va�T� "OV�b0E�9l[�����F�6���9�"O֤�E�+#��r�����q�"O���G
�9?�AA�G}��`"OH�X����(��-��W:x��W"O���� ]�i��8��R>Tt@��`"O�aɵ���U��ib�@����S"O�Lʂ��
 ��P��۵n��{`"O��ӫ$ ��;���Jem�r"O�AZ𮉅uxV\��*��UD�a��"O�9�V�ّ&���	�4���Ⱦ�y�d��et�ӄc\�M4�x�%M)�yB�9r��&C/ Ek�LS'�y����OfVlc��?A����%���yB��)BϤ�p��E�>I�i�k�4�yb��]_&��$��5��u��욊�y��G�w.Hi �e!0=������2�yJ�93W��&�41լ��d�N9�y2��2XHY��Ɋ0W�0����y"�ґ%����*^)q��2�#�y2�Q�B�~� ȎS氢�͐��y
� qqFvB�P��AR}�BŲ�"O���ǎR�1��l�D��t�ٺ�"O��r�]b� P�@�u���!E"O8�J�ֻY�.L�פ�(�~ԓ�"OF�*���%j! �0��{���"O4��LV2VXne�1�J�'m��J�"O:a����< *VI�b`%wv�CQ"ON�;lR�7�����Y�,^�)S�"O\�@���8x,ؘ?��jW"O��ޡ�X�V�ޑ
-�y��"O���!X�W�j�p�]�2�	T"O����n��"���B�o�b�"O�5�4�!ȅ
XN8y��S��y�N�e����D`U�T�@�C?�y��� `R�ǎG������yRˏ�$`���f9���r����y���!+�f�8b�ڀ`����델�yO�@)*q�JʷRs6��a�O�y >v��X���Pʵk�#`ࠆ�=z�*�F�ԅ��Ͽsb�q�ȓO3��3�.}U�Y�.��X�~P�ȓd��H�՜u�ޘ���M�cI5�ȓ�<3 ¡l���"�ԩ��$�ȓ����τ6�x�E@��k����ȓOb)�3F�]�݀��.X��0�ȓ#��Ic�Ի0�
p��#A��؄ȓ^3�c�՜nn�2��!�"܆�l��4Q��V�:`��;H�9��S��@�闢uG6YZ�.��g�ąȓ)�`�u���:�Ե"�G Z� ȇ���Q�.�f�d�R�My� ��f/�݁s�ɉ9s��s�N5`��� �R�G�7�����b�K5Z`��;3�y�S4s"	��p6ɇȓ������-\����y"��ʸ�	��/Ҏdi���-S8.ȅȓr'�uU�ۃq>�
RH՞Y>���q��p�g#�M�"�Ӣ��,ͅ�ݨM9Qk�0��l��c�/M�نȓ-	~���.֥d\�`�S��,�����3&:9��L,"8�����?�`A�ȓ	G��9�I�O&ԭ�䪖;)x�ȓa�z�ДB"����E�ȓ�B���	�.'^ެ��#�rp��>hP��o��yE��1v �T*$H�ȓz�:�0��(6�:Q�3`�g��p��	�,�h��ܑ�,8p@��jI:i��q_TMe@̓% ��mtN�I�ȓK6�4b�C�%�������������@��8q��clw
�dE���ȓs� 96�!Y���t�#����ȓKa���JĨ?x�-��=�.i�ȓS���#�EL�a�ֱ1�� uJ������c�6L�B��>Dه�-�l�j��ͦ>�$D���ץ#���ȓ\b�5ϯAxNYA�H���Ć�=&Pq��^�* ��x$$�'�p���le���7HM4� ��`��p����d����B�$��#Ea]bU���e���G3��Ip��:�����]�T��!u�}���4����-�6�!V-��Q>����W5Q }�����ҥj�1��Y�R:<��ȓ:�>2�aΨn�p��eF�W�\A��S�? R��Hݱ0M�� �c�Kd&��1"O2$#QL	�H�h�KgB�WZҐq�"OL}���ڏt��e��aɫ=�z��"O����	��s��2Z�,��"O������7����% ��G�(̓7"O4�Y�*љ|���d�T�!�VT�"OV-�uo��m!�����W_,��"O<h���F��\��V<CIh��p"O�jd�ڼo�\CD���15<�8a"ON����[�O�>��$nǁ\$��;�"O�ʰ���3�X+�N�,�)w"OBȸ G�St��!�*�L�Ƞ�"Ov�����rLpU��A&qC<hC"O�!X�M�Z��2)IQ��)G"O|�j���$#��Q���U;$���"Oִ���'b�� i�&h�����*O2胂�!�dE �[�^i�'k:��"��$5�8���ԣW� ]��'K���f�ڱ�F%:b�W�p{�'�~h��@�d��t��J�A�	�'I��q��Q&�d$�vb˘8�J8��'8�e�R��#��m�5��5 \QA�'b^����*�H�Jtj��&��(�'D�У��#jh�A& S����'�!�s�9I|�s�����P�'[^���G�K��qr,9�$�	�'�Ā�6a�D��L��l�*-DE��'�l	w��Ok��P�f�&;0��'R��G�� y��Q��lE��'nDTc o��V�9R�Lۀ}~q!
�'?�[����")A%�T�WB.5Y	�'%�Ř�t��  5�)R���'�|����ԇx�
I�+��NP����'^P�AE�Z�I�4Uj�o��?�h���'S>��`�L<~����giٍ9�d��'FqS�㖃��<a�j7��,X�'=0���	Qk�5p��ړ:uh���'�j����=��I�mS�|�f�'�����+K�P��@��>|w@|��'L��CWlӔhf�q"0I�1 V䨲�'fr9�GI]<\�7�^A��
�'��P�F��~(�
��;3�!��'�z����Q�_n�u�������	�'�̃���m��U��hW�y��9��'�α�"MEqZ
	1��X�#��Qa�'DΔ��H�Ej�J�M&(��I��'��tr�e�Pc�x�C!Ї0�L�8�'"}�\$4P��8��&T ��'�t*�f�\㐌��o�8�i
�'�|3�DD6(��@�Iά'�P2
�'⤡W`N}�B⦋�0 �	�'���@Ԏ&�^<J6h	z/8@c	�']��d�F44t�%䗏F����'bq��;�M����1J%r!��'�48`"d�;a�-$� �H�y�S�w���Տ�9�뀫��y�n�v�qKSKĝ!��`���L��ybG��$���@�Ǿ0��h���y�_�%/���i�u�"����y�hX���\�K�0^�@�����yB%ږ��E��n[�~��k�����yb@��}�tSTO�n[����y��W4!`d�k!b_��
d!�5�y��� T{#��[I��
�M�y
� ʴc�e�8�B�D�3�F��f"O�  �,ճM��ZGF����"OԤ�3�p�����L.Ğ��V"Ob����8)�pI�)��mNꐅ�N]L1(�@��Ba�Qч�^++O�x���� �͹-�8qD�� R+N���(���ZG+ô!��4���3	�0��fU`@�'�ط[0�U���۰V!�m��06�@�E(�<���P�8n�x�ȓO��k�&I�f����C̈Ec�)��me�4Z�Vj�tF0}T�ȓ7���+�+� m�Ld#�"��]?�Ն�	�P��0)�$\HA��[����ȓ0�����,�6c:����]I����ȓ�n��D��0Z��͢pN�=L�l��#^�	�ӎ� `����$�p�a�ȓj?H R�ؕj��X�Q��.(�X���C���2�b��{� }�uS?7���f�i�E!�N����X#d˔��ȓY���R�Q[�5��M�3k�ȓW�x�h]�:�mJ��0#5d���3@��@�K��^���39	�L��Z�	aS��V}Nus!�ɫj��ȓ70�Y0CB�xy7����}��V���Qeh�m3V!Y�#�#'P��ȓ_mr��6�НI庠Bui�@��p��8�����B�IAx�1 O��L���ȓ'�eB�h��A�I�Ɵ�:b��ȓI����8��4�7&�T��G�z��"�Ċl��e�51v�0��D����5޺�x�P/W�ҡ����$!i�g������{����ȓo)��y�F@�M�����F.SC<��ȓ?c6�I`�L�W�x�y!ʚ"0���ȓF��m��a�4.�`�ԄK�R$�5��dlF0�f)5�U�C˗P4��N�&,kc�GY�	vF�	�詇ȓs�e�#a� 7Q(��Ɔ/}:�ȓ4f�s�!F�H��f��O�H��ȓeZ��ʤ�߂/�`����?P`C�ɀ7���l�7$q�(��o߆r�LB�	>=KH9�b�+sxhp��6:Q�B�I]X��À으H7�H��'o:�B�ɣ= =�R��(|~n0�eG��^�B�	I�̪@�_�Q��we�.24B��#2�M��/T�!�H��\<]��C�1�b�J�=��:t���zB�ɵTa�ͪŁF&]P��G�֖?�jB�+|�J�`�iCZ��@q �ƫan~C�I8|eA��'fb�)ը�(ݶC䉁'��Y��r�AWǜj`B�	Q��� k�-n?���À`
C�IY���p��:F���릪֑L��B�Iu���soN��v�s
���C䉰J������L�!M�ARl�C�Ig�`��ǆ ��0)Dн?ӖB䉊~p��	w�ژ�d`P)μ$�ZB�	�X:�! �!Qy �]H�N�aJB�5j ��G��%!��g��
LBB�IC8�.�}� ��!��/�^B�	%��4%`	
��Ԉ$A/0�B������/>'�h��s^�z�B�I9~�����:n�Nt9�)\�W�C�	���(0�G~�����4ny�C�)� F�Ô�F{��6�������"O� �	��jH�q)Z�g��H
�"O"�p� ˶/���DHY40�����"Ov8X'� 	B�EH&ʊ�8�hTH�"O��*���F��rh��Z�,`�"O��x��S!f�UKP�����b�"OJtC�(K~FL�z"�Է3l�"Ox�)�m �L�b����Y����"O����,{�|j�M:i<y�"O���+�v	�B�#
}�)��"Ohx&	A����	��\�Y�pR�"O��zs�ЗX� �%�ж-����"O��"����.��1��,�hp�"O�H(``L2�A� Z���hv"O�!Q�-� *(�t@B~7 Eٳ"O�Rs�66�
�U�8>�S5"Of9�$m�%�b���S�� v"O��r" _�I���0�̠lX��8�"OD1;d��6�DJ��ս-V�y�"O�|�ƃ'eUd�1��S�ޜs�"OK_��f� �#��(v�@ц��yR��@q�Yb��3%?2=�5e��yB�ǩY��Iˤ�ߎp�d�DB���y��&U�<�3W�N��ܥ�����yB �d�-"k!��@���y��FtX����!mQ(0�L*�y2o1WW24BE�0�q��L�yB��u�hP*��T�Ө�c*?�y"����zv�M�y<6�
6F �y���w��J�Η�z&�9Ū3�y�OmZAqP̙�H��$"����y�
4K"}� �ż=�jJ%̇)�y��&��i�%��"�"]Y�L��y��9~�d-!ǩ�6/�*��\��y�'�
�"�YS�&�I3�[��yB��?\HA��!S�rL���y�k��U�t�s�f�3�t=��ひ�y�=5�@�1A�@�'N�%�v����y^�R�⠧�
�����y�B�����b�
]��+5č�y�D�Z��BÉ�Od��X��	�y"��K6��2�Β$^���1T��*�y���>e�4�Ue�V���)w��y� �c�f}�4-�D&��*%��0�y�hď"h9i�I@�O��լB��y�؎.d �0�K�]{Ll�'
�y�����IYW��&Ut�5�Ɂ�yB�	�C$��L�wۄ��"J��y,Ŭ[�p�v�>v	6�P�L�8�yrkA�VS�9K$%m{vD�7*B!�yb�T�&[%��(O�c��КV`�y�$^,	/�<c�k,�� ��	ڝ�y�F�8������Yk�,�bO߭�y�C/ ��x��Jt���O���y�ϛ<@���և[�@�� �����y�CRv~\RC�^a~�Y�_5�y���6��s�JY���̑�y��
�:�e���V���1��yr@�x����f�Qq�Pi!�%�y�YT!x�2�BH�Ln�͐��
���=��y�FH��1X��E�H"Ԙ"G��yb`�3�`��D���.�a����y2��qJ���F���x:8�#2�y���`l`�
d�
T����0��S�? �9�r��Ԕ1C�͇�"uK�"OH�c6CC�!6>�N�Ѡ�C"O��fFX��!f��Y�
���'�1O� rq$�\B#E�}�&�C"O�	���X�bk0}�n�+�,䨓"O�I���R!�dЪ`�΀(�"O���E�W�EФz�a,���y�"OX�0�$��	�D���Ś�5 T���"OVt���ϕP^�r��1��D�"O��; -�t�v��aZk�Ɣ�"Oh�#Ëq;**�ƍ�_��q �"Or	��/H6J#�H!�'���<�Ђ"OtlC�L�O��0��Ǒ0�|1�W"Od�&Q�l���i�$ �tx!5"O�jf�!CK�p�����D"O��2ƙ5H&�Hq@c�/X4�+`"O��� ���0[�����"O.� �$R�t�\sHT5U*8b2"O�ԓ4��w��P��P�]��ۅ"O@�ȵ�.b�̴!b���S�&�+�"O��k�l�W��ł�E���F�Y5"OX�`&�W�7t0�B�e���;�"O�yb����p�p��1\%�"O�y��O�%7��iWjV����"O��ӫ׭t�\��f�%�z�b""O\Ɲh�;&��8 �fBa"O��\���I�E�j���"O}�����UBc��$�XT�f"O���b�Gu ��4&W�"<�Pe"O�Z�/�_P�E*Vd�_*E�"O�(@AљB�0�Xe`�)��k3"O����NY����Ȅ�t� xp"OlU�͇�h��!)蓝:�섒F"ORtб蝺6(� IuG[7�X��"O�xa$dȺ[�֔ud>�<�w"OS�N1*l����M0�����"ON�㣏�3���r��D[����"O�%cB圯y��1�f��~VH��"OPhF�=l"� ��<*D"O�{�lâ)�X�� (H#720�"OF�˂��*#� ��E/Jd0"OAp��Y�6�!+�䌆o�p�"O��хސY���k��X����3R"Oxd�ǎ�)L&��!��v,�"O����j\�TЊ�`U0Z��T�a"Ol��LP�q�~�b�N��g�l%Y�"O�P�m�+/~~,�/1D�y�"O@�����aX���x		G苪�yb�'I�ک�g��	DY�0�VB��y�lU�Q�p`p�)��5^,lsw�̧�yb��<���"�*z�@F�y�@" �"�8!H�u�D�E��<�䓯hOq����D��� H��-"��M�w"O.���M #[�@ExC�4�5"O"��A�W
02��5Ċʺm6"OD��Cj2_����5X��IQ"O��DDW6i��PmD��0�E"O��f��7��i���>~�H��%"O���@C�kB�U��i������"O���E���Ȥh��9��H�"O|�H��
!*��蚅4n��@�"O@Rs�Z$b1T8yeG��>h<�B"OƩ�&T�m��E��V�8E$���"O�9�΄��L"jA�GATy;w"O� 4��LAY�U�E�G�5x,�"OȤ�mتh<��q�痟 ��dT�	c�OgX��4�7 [�L)t �@��I	�'���7l�9��l :�����'{`�x��ڴ
/h�"*I2p�	�'��Ȼӊ]3B�Z)��N7er�'��$Q��Jh,)ѬH�w�M��'��d2�+K�6<Yy�
e@)��'d�u�Rb�z6�8��כZ��uʏ��<��	7\>�� ������I��<H!�$�Y�,�����8�8��7;*!�D���THk�'XU<	�7I�9`%!�F�;-��A�Y�:8��q��S9!�1��9ɥ�x�ޅ�e�W !�dD��`�1 �>{�04Q���2!��R�Y�b0%4:��D�%fL?V!�D��M�йÅ�˕R��Ũ�%�r!��?I�A�s)�M�Dx�Q���Ic!�D��D�� 3,�M���3PL%5U!�$�5��E���]��pL"�C�;=!��7Ϫ��%�M;�<I	��R�!�WD0��R%��J�t�<u�!�5i �s晚6�� ��ښW�!�$B�OXDId�I�#�2Qy��ʆ,�!�d�{�p�"i�H��1�T*r�!�d�� x��Eh��%��`��b�!��Ҡ
��p�D53���k�Fďg�!�dĊU�&�{���K�jِf�[y!򤘮Q*ܸ0w�Ҽi�PٰCo�'9�!�d[#OM"E��A�"s-h]��Gs�!��*�${q��	Cf�p��0	�!���`��@��i�/f.qڡFĬR�!���D����W�] ��Hf&�h!��1gs���C�"[��h+sD��Xa!�ܺJS @�Ei��|��a�=Z!�S B�N�q�G��lT+U`�1~N!��՜ʄ� �HѴdP �9=!�d�H�v0��/��s+~�фJ��f"!���-�� @A� �މJ���(�!��8r#�����#�	����!��!t���Uk	��l��ԣ�!��<^9H�@�Ĕ�u�|L�0�T#u!�D�#�4�g	U4w��=bqd7C�!�ED�]Q _�aL��;�"=�!�ɳe�p`�*�JR�c��5R�!򤍆{����E�+H6����,G!�ΖR�64C�$7A�H�c ^ !�$_�K�����2e���� ��!�d�h��`�1I�"t��xi�	��e!�[�.s����V�RÔ��ab!򤒆^A�8�S���`�2�j��V*=D!�D >~,��$�˶c6��D+
�,�!�]�1�y���h�*��KB)a�!�&�D�Ev�D���o_=�!���3%�d˓�էj�*-)�NZ%T�!���Mp�<R�Մ?:��aE8/�!�D�-�TȰ2A��v9�%̆�`!�ҫt��5P�$�l&�`�!�!������-�W��[��ɤTh!�D݊vѪ�b�)�`SH!e�!�� �� �n2{���f�62�!��F$�x�
=9p�H%��.�!�d� 1�|2��ȲhHܸ��DĔX�!򄆫:A����G,h�⟣�!�� �t"�J#a%� q���
#���"O�S�W�g�@��|��]:"Or���-݇q�>0��Ǎ����"O�\R�O7Z^�� ��L�|ݫ�"OPU��o˻�Z�2LǻGv���v"O���v�}��|���EM"�"O�M�0�F�~IBMzgM�<M�u;4"O�x0%��PSPQ��kZ!3�Hص"O6�(��IEtڈ��`\�v���"O������|�`�I���0`j)�$"O��H��L.Z`�Pɛ�`O` �"OH(b�O3K��Y�&��5J3�@0"O�9�%E��,��h2r� �"O���4�@���0����|j�!a"O��p�'2i2t1�A,c	܈"O����O��
L�@؞��@D"Oz��1���N�����y��*"OX�a���%�����Sk��Bc"OX��C-��%,� a���`)Z�"O��wg�r��pس��3��H"O���<<�R1
'%N�x����"O��B�hρ9:�@2D�#�� @"O�Ibk/FH���b$�B��"O��o��t�BAWa�<ȃ�"O�������l,X�j��^�8�B"ONpc�J[�Z��qc���p�ʼX6"O�yI��\���M��L�_��M�1"O`� ㌟0
̖�!��;A�Lq�"O���F�D��A�Ԭ�"}���q%"O8(R�JǢD��
0��
y�ɰ�"Oδ2�)ނH��-asg�n��!z"O��8�Ku�u:1'	9WĐ���"O.5�gȏ&~�t��rF2�H�"O6ؒ��D�B�C6{F�Җ�I'�!�ĉ�`&�@�B])Ww�U�C�94�!���v�`T#�dJ�HZ <�� ��i!�ĘB?����gИ-��q�aE!�D,>�Q
�,U�`�#�B	�!�DU�9v�|y��-�zT�dm8<�!�dŦ"�F0 �� Dj�1<�!�$B%C�F�1(Z�_�u)��[�!��w	����ᙱ3~��4A�$�!�$ń{d�����	]�mP�O��C�!�$	�~�xa�G�QR
l�+�HE!�Ĉ�JlT��D��B��e�e�U<l*!�DSY�ȳ�iI3 }�yj'�O@!��\u��҅A��DIp ��)rP!�$S#>^Y:��#!�r����
7!�$�"}Xt��5�B$��-i�	#I!��[2v�V�0f�\�Zw"��#J�.>-!��G"�]�T [°(5�օX*!�h"a��	Q�o�Hؐ�r�!��'L5����h�	rK��&FR�G!�䆗h{~D�E��&Z-�p���D�4=!򤚑?���� $Ͻ8ʝ�DD%H4!�D�p}�qk�@ϻI���cD;!��&"�] .�@��lx�/�&�!�$�1o������Q��ĕ`#��(&�!��X?i���KN�g|� �U�^+�!��A�0�t����j���xf^%[�!�܏lKZqx3 
�G�f ����
7!�Gr4đB� I�2���2H5!��8i!<Q
C�3h�{��/!��3}[����,]I��S��?F!�� �􁶬ќN�BD��B�T��	w"O����`ĪI��aR�w�ڠ)b"O܈q2
BO������w��}�"O�M���#2���i墒�xd�Ag"O�)҆L?a�Q�Db�?Fb" �"O2Л��K�|� �'O,=ґ"O�@H�+7!��àS42	@""O�M#D"f�x+`�T�a���XP"OD�婜41��4ȃ�wm�ઠ"O<��6�pMC�M�l⤪�"O�(�EKΕ9�(�%j	�kN��6"O�0��@�1<':ëS�+���J�"O\��7��B	�o�J������s�!�$\8[g�]P�Řh���JS�!��ʲi� њGc�1^�ꍗZ!�C>�,��xOT�%鈋s�!�� �0�ACN36'r��7@S�!��͟���8��e*�	����*M�!���M6՛�����kaB�0�!�DN=3�Q:Tj�O�Ƽ D�U�|�!�ѿ�|���ON �����4`�!��H/�H�P�¿h"(�ceII�T!�)V2
�%�'b�tl�ő2K!�;sv,d ӣWY���#í��=@!�Dn��t���آ�M�z�!��

<T�!0�ۑ~b���5L�4q�!�dŽfx�PC�Y�vM̍�L�)�!�\"w�EGEGKR͒����_�!�$+�ZpyP��+_H��a`G��6!��1�\�D�V�[�"���E��!�d��'�N��B��29��S���$<S!�׏m�� �:L�|����!�+���1�N
MIq�7j)�!���, -�G×6x!��J��[ !�\!��ͣŏ$
CQ�]�P�!�L�l,ܐc��;va
vhVe!򄍓U:��v��>k�}�󠆞�!�$��s��bp�1o�d@�N�)�!�d�=tZAKA�ksн ��R�d�!�_�Y�0�����w�I���Hr�!��QlM�0A�L�u��y�j�M�!�͂/�jqC�%]�6q���2d�6�!��ԋ��uҴ�&���iA�_�^h!��ՄT�x���B�\�Z5�f�V\!�d�&", �0�/G�x]wi��YE!�H�F��\�M
��M����5�!�dD�~�|�AWF֫:��r��!�D�6)R���V��:B1�&�!�d:ň�W�T�S�V�K��g!��'L�����If����5��2!�d�E�p���ǽ�n౐慽�!�DV�u����M_.>��� fWe�!�䊊i�
��I^�`��(�&�V}!��U�V��
 k(G����Eś&�!�d��V�4�6H~P�X1!�.�!��։w��Qf��i���,{�!���� �Ci�9B� 9E�@�y0!�DD�k�f�ap�_IyP��Qc�!�[)"p��Nؙ|eP��Lr�!�$Z�xO���"��-Z$l2�鐖]�!�>�2p�&�-mA�p{��ʧL�!���sҲq�E�n0TX�զڮq�!���t[<A�v�W�b�@�BS!��GS���0���S�B�q#���!�� 6�Uk9c[L��2"Ϛ���Y�"O��`r+�zX�2�a�2P�Bf"O���$�'H@!B�I�<6h
 "O�!��*��t��hT�c��y�"O�Q�T'rH�����*w�,̱%"O�dX'"ԯ��q� &@�h��"O tQ�ޖ*CԱ�
,W�h0�"O�dX�F��j@]
�
����Y%"O:\��$@�f4!R�h�/���"O ��7��=oi	3�ΌOޙ�a"O��{��ǰa總�$��
o04��"OLE��ázb-�劫?)�x��"O^��&p�0醃�xs�(j"Ob�2v��|�t�#�z?�T E"Od���LՒ:Ѹ�#�(q�-9"Of��&Ю,�9d�O�6<[�"Oֈ BI��x��l�Q$C�=�x9�2"O�p�T�Ϧ��0�
����6D���3�Y�_hFa ��8���Q�>D�8��!�%!F U����E� ���<D�����Y������(c�6�q�<D�l�!��X�^ �GB%�>p�<D�D��MD�jdᄄ�T�tjV'D���$M��`�n���
�4/���?D�H
q��%z>��I�l�.(�5��=D�0 ��Fo2�Cc %oI�0w;D���FػL��pd�G��U�c7D��A���s �1���4l�Q�6D�܂�
Й+2�Y5I�!�bi�O4D��-P�i��YX��)(F^�s�7D�(��Ȋ�Y> Q���� -����k8D�l;�c�5�@��f�R�N��!�;D�ԃ��Ӯ%�����CM��Y u ;D�DJ7%��@��T�@fP�M���`Ѡ8D�l�F��:[�%����%L��2��(D�,Q �]�.x�DG���R�<��YT�d���ꅰyA���a�K�<a�GA�����ج>��-����I�<IB@Q�	2�˦O�c�@ 1�L�B�<���S���i�1na�����s�<!@gO�v�F�J7ֱ&�+�k�[�<�`NQ���PҲ'I���PK�\]�<�O��+a�бS�m���2IUV�<���L�#��)P`*Bwx����A�O�<Y��������HY��X�ᩅH�<��¹KB��U,ɸ^���	 �L�<A������eJӳ]��9� �JI�<	V��:�pİ�n�7g��e�ĉB�<�gD����9Q��-wH7�S3�y�Q</=≃��@H:�" ��y"��9r�J=K�AK>2L�h�+D$�yҦ���ӡIT2$�p-XL	�yb���~^�R"������P�y�A=P۔Ջ��+e�TZvHث�y���],dIy���6!^@�3VfD��yr�ۼw����`�d�p2狑�y��2�8�P���E���1���yb�X�]�p�� �/ج�!���y򬆄�4�� H�,J��X��P1�y�ǰN]ذ�d�߭���zR�ؒ�y�MP�	1�yiâ�
t(���"1�y2�P��������c~�D���y" �R*t��OR�O���h���y����:�x��.O4ؐ1���5�y
� `�u��?.��3�Bn@X��!"Oځ�pD��Lp��NH����"O�u
Ga�O���Z����E��yC"Ofh�FC�I�
�`�mJ�G��z�"O�,Ȱ�F�V���j�	t
FJb"O��8��7P�9���=w���R"O谀�#]*=nH��'�Ԛ�V`��"O���j

\T���q�.  �"O�(j�$�=\�x���h��iY�"OhH(�Ѷ����P��t#u"O�)i�j^��R@ۤ'D��n@4"OJ�v�޶�s�EJ�s���Zb"Or���A��d	U��5�hC�"Oj8����*�r�B��P9(�0��`"O��� C�:11�@��݈BN�E�Q"O�Rƍ#�B1y�D
=Uf���"Od=���P���D/Q.!��"O���E.۪e����1N�,ä"O"QH"!4.@pDa�[>o߲��"O���VJ��\��P@O�z���)b"O4�kBf� {�H��ʉ^dx��"O�����ĕE�Z�	�e*wS���"Od(p��æ}g���v� !I�"O�92pH�*��� K*_yR�6"O��r��(i+���B�^pvI0�"O��"sX�70��D,��IZ�52w"O�)U*�� E�X�!E�Rxy"#"OPus7	N��Du(Q䐠6�H�b�"O ��do�T�$���!C_
T��"O�QA� ��]-2�`�/m>�d"O����e�	��-3P�0<� "O�aqE��Q�L����f�D�D"OL!�u�N8�5�&�[�D0�T92"OJ��g����i�M�9+�\��"OpЏ6�$)��-�3a3���t"OĜI�N	�z&L�%g��R+�QZ`"O�dɕ�L�XM���b��%;C��"O��0QGF `��)�a�"ʪ%�"O&(rg��4�r��I�Q��9��"O�͹c��0'���V��3+�	b"O�5��$(3��Wm��
��Ez�"Or9i%�O"����C'��0�2@"Ot �����#K�\�b&Q,;�\#A"O���.T����OD�Yr"O�8�P��O�t$��$ҘMK|��$"O܅����Z1�cF?=Kf���"O�ٸ��#I��@+����9���J�"O�L#��	����z��P8)�q"O��;�N#D�DXnJ�%s���"O<�(BKϕb�b}�T-�Sn�� "O�ի�V�^���쌞} F0�"O���%A	[�$Iɣ�Y� u�� �"O^��v�ң�b�W)��XA"O�� ЋͮZ���8���"ջD"OJih��]2Y��s3�H� ��"O�8@Tc(	ب�%P,#=��c"O"P��%|&H�E�R�B�&�y�"O4���#��Q�Vx�F�ԁ�F"O�[�l�b�TLn�� ]=�"O-�&���iD/S�*��p"OT �Q)�?Oe������/10,m�s"O��)�eX:��v�B�k([�"Oz1
���?@�Jԉ�����E(f"Oju����ym����$�H�0�"O� ޼��	ՉH��9Q`��*� �y�"O4b�J ׊ c��Z%*�2�q"O��1gA��cg!H�U����@"O�1����ڜh��H0m�(��e*ON`��
>B㆝�D�!�DB�'^�p ���$�@Jd�T�L:���'�H�z��$}YT ���?�J�
�'�f�Qu�� 
l�¯\*6!T%�
�'�P�[o
HZ|m�,Гg��C
�'*$�� ��>���c�BK�^o��`�'��ek©P�*Iz�e.O�}x���'�(˶��Fք ��/�PU��'�}Qr+P�<*�4�C� O��8�'��k/-ɐ))󠃽x��Hs�'���2�*������z�<�J�'ݺ�	��J��57��;+�QH�'X�D�>y������'۴Y��'
��R���"�ԃY8Ȝ!��'m�y���t1�����m��'��q��X�s;X�C�� vq�D��'�Hـ�N���Ju���Y�8�'�
��c�"@�$� ���	{̪�1�'���p��N���H����y��)��'e8���&��(	1�M;l��3�'�L\�
4�ā���[{Ͷ�s�'���:��.`��S���x�x5��'L �;AI_� �~�c�d\�{����'�b����Q���s� w �d��'�j�s`I�pv-�AöY&ԙ�'%�i�$$U,\�'��		GP�	�'d���Y�h�x೧�X+*N�!	�'�Hs�iF�}r�!Öȅy
h��'�~�X�f^	K,n�8E� r�tU��'NN��M�	z۞`#V!���HU��'����BDG�	p���[:�6�!�'�Љ�P�	*��D�5�U�c^���'�Mp���q	传0��+\�K�'9V�d_�`�*��v9�M��'+,0�� C&H�V�z�L�XK��J�'Z�QX�S�
�T����'Kx�:�'�-��/R.QO�C�JC�x��'�0��'�(�WH+B���K�'��@┫�;+�eJ�#�Y��'�
t�/���P����%Y|�	�'��Tɱi��"�9JC�_��̴��'� T0Ae;58j��BE
a8����'p���(�-}W z��Z�v,��'�l���ㅛa'�ث��X�}�,�s�'����Tf*`����tV�0�
�'��p7fC&dZ@����#lJZ�q�'D�3��\�E9�5��/qi��'�n�b��ڛ��<���Ϧ2+�'�u��X+`�����ÃyR$0#�'ͺH�gT�&�H٫� `Q�+O0����U�*-�P4���bk�6Z[!��� O�5
c�ږ-{�ȉČN&!�D�*޼��7�U����i��p!�ą	$��И�]W�.%f��x�!���"N����+M��e�#^���wx�����]&=�M��B:|(	�C:�O��K�:�b-�~��s"灹<s"d��)^��5�v��P������-�^��dMҚ5s���Ō1m�4��ȓ��4��`_�T�b�2B����(Γ�hO?� ��	��%��3l�&QJ��"OV��.	&C�`�C��0�QӐx�'�D웑��%*�vq膢��9��y
�'�f�u	�Zo��y��I �+�'�~qXe-_-VFDh���;��y��'d<�8SM(���`=08�u��'�tj0lV�dG>�Ō�,�<��'���@�ˑl�TĂ�(����'��`B'���b��9���ی":X��'��i w˜�ٕb�
�s���� 6D��J���H~�Z�	�\ �� DI4D�����\�$��� !lj��l2��ӈ��E���)%|��J�mW�v�p� "O�]�D�Ǵ[q���Ǭ԰0�u��"O�x�!*�7�P��0mo�(��"O*܋��_�z�x���
�\J1��"O����ɬ~�\b@kKK�4T!�'��I0ٞУ�$�)RLa�'"ѥv`C䉾d�a�Af׹.FJA�Fh܋r����)�%Ta`���R��K�~��ȓ#��X��*%����oסk�0�O��Dz����>�l8`6A��b���S�]<�yҨ[�d�X�1��^,0�lYhT6��'*�z""%S.�|�4�Ҏ-Rv �r-�7�y�$k�b6Mծ4�����%�y��'	sD�J��R51"��`����y��G�6(��ö���.i��r@����y����S+Ha��S�o}��9P���y"lҳ1wR�:3�ɿw���Z@�3�y���".��9u��=hj �R�k��y2�� 
�D�v��Y�����ybl\A��p�bʎ,�YdǾ�y�d:v
���F�@�V������y�.S�B��(�G�Ɯd����C��y�b�	[
��HۚQ�"賷+��y�̐2~K@as�DP&J!ԉZ���yb ��l���AF,��,����+�S짭?�fB�}�X�⇏՗JS��@�i[z؞(�=�u!Լ��|jeII	ع(b.y?1�l
JU2�/�����W��1^��?��)�t��$R��F'� qDTa��ljў"~ΓD��"��0S����JS�B��ت����~"���'-��rB9N'�� ��7 ���
�'�:4ʶˊ&>&�#�c�/�*�0���hO�>mړYFn�30&ٍ>�As$*߾d�B�I>3�|��h@�:D�'G[�3�J�IƦ�Exr�=X��	�� �TA!L��%�X��D5}r!ɜ"Ɣ����:����y�!˦f�l��ʭI�� ��HOj�=�O�T�!��)Nzl��A�P�~�.|�� 6�%�c�Bq�5���l��'�ў"|:�i[�iD`|ȥ��rT�p�Ec�<1d%V+*�X�K6*R!;6��Ĉ�J�<)��	+g�\�VF� *����_�<IS
t�&=0��:��쐵L�W�<�vCժ.�Pa��i����I�<���,.�����&E�hP�F�<�eꆢ\=�d�Q�&G.t��d�<9��3G�="�O�1�tX�{�<����]<�$�����|x�4�Uv�<QBN��JD`���I�yԩ�n�<q�l��S¤ڟC� 4�o�,�yr�ڟ`��ha�Å�#�:�������y�FF���L��C��+c��jDaܯ�y
� ����%"YjM����)u��d"OН�E�"N�9��NH��#"Oʁ�$'��5�cFT�f��3"O4��ϔ
b�~I�Uď���`ȁ"O�e:c��7�"��҂OYv����"O�����.oi�lh���
eT���g�OYD�90�U�#�*XU��7.K|�k�'�f�����"q�)d��;��q�'��| ����?�\��c��4��)�'*�`�$�8�(�ȁ�2��Q�'a6 ���?���3�"^_D�:
�'޺(+0��}�L#��S�ZE�N�lD{����P���B��e��@e)���y�&��M�,���-֍]�ީX4h���yb��=��U�t#NYd���rJ���yb�RQT@��GJ'�	:f��y�*I�^�U�J�1V��0�V�~R�)�'g���F	�pT�b�ٰ{z��"�f@[ddM�``J��`ܩ4N��M2��r��)y�	�DC��"��,���I1~���$F0k��8(�Zc$C��X���:�Q��C�)�9.���<�W?I���J��=��C�T��	@̞֟܄�o��ժ_.B���r�ج	xt%�?A�'k�?���Y�K{T�� l�73��5D�aTe�2�̂��W��3���<1��O ��h�������ʔ��s���{B$�,�!�� 
�(��9��@k��M!�DɄ2��$�WD��	��X�4�A�Б�d���h��!� �I�7�<��e�TI�L��"O���"E<��͕�j7�����Ir8��Ye�� ��I16c[�K�\�2&&+D�,��JD�)b�
�*M�e4 p$f;D���b��Z|8�`��8`��{��=D���#�4Ncl�{��X<P� D�|�J
5`u�*$Bͧn�:e� D��k��eO╫�G7h���G9D��*t�� "��6⋈t�y'�6D���d A)��
��I0e`��s%G6D��h1���a7F�[%"�����g�>D�x��к@1:����[�b���Ч*D�P��@�5z��ŁZ=?(9��A'D���Ӆ!}�V���"J��t�VD%D�`��2�Dh�kR���@��>D����jB�kt��[���*�ֈ�we)D���S�"K�h���xj�<��	)D��PU"� j�����&ٗ�쌣T	)D�L۶��,lx�A�dק	�p�8,&D����k��"ur,!�OV6s5R�E%D�1���Q8-a�gR<Zw:`Q')D�4��Q�a���*��\� �,` ҍ(D�4
u��:�*��:�$Q0�;D����#�.�8�ꥅZ�rP�9�O;D���q�;$����bʜ�F;�����7D�h� �u�z�ӣMP<�����0D� ��I�?xbp,�b*�RLt�aj0D�h� �9v��ؤ"'oKP���9D�4���?���B��f x��8D�H�0�K�}j���І�:I(4*g3D���ƪK)n<ڵe��]~�9&�6D��P��Qu4��P� &��k5D�4��������S-c��!�/D�����)jO�!��H��L9���P�-D���U��6��ɫ7)��ʁ
Al>D�� ~���C��$�q�G<?8��"O�L����S��P�-�'w��H�"O6�:"�X�L�P�Nɳxl�"O��Y��VG:�02/��rW�8!"O�Qb�$�V%�3K>N18�"OH8���Y?8�J�A2T���"O PɄ��'�\��a�3.�`q�"O ���CE�R�刐�E+?�����"Oz}H�j��@�Pg�_5%�̻�"OҔ@kK�n���� �,
�G"O�h��Z"_����΂��A�"O�I�Wa
�[��R��3*�ꬣr"O��`��0pd���Ok;��B�"O��
�a�?U����L�,���q"O�����(1�c'�údo��B�"O��B��M�ȝЂkE?d����"O�<xaO3P���ya�>=�0�9P"O�|��
��v"�f��J��RF"O�QY.��x��M Ed�8�h���"OD�1ȶ�b�˕䕄ٺ�)P"O����i�<^�DiQ��"��Q�F"Oz��&4
�`6�З�^�+�"O�a��+:r��C�ѵuxx!C�"OJx�G[�:��ͺ��V 0�E9"O�f$��3�����&S�*|)�"OL���ǈ�;�޴��Z�o+6���"O�@F�"81�@(�+�py��*O��ƍ�O�
���A�u����'�
=��Z�Z�r��aID�sC��	�'üY;�i��|6V�A�'CX�	�'\�}r�"��|rn�蔍E5����'_>}��J�1Z"��cGj�Ț�'yg,��C�|jdDK_�Y�!���,���A�K]�8A��K��!򤀑'[5:�B��_[8��q.��.����x!�|≊z7DL��ְq4�pa�F�h9TX8�m�F�!�3[�tɰe��L%ڍ�qɜ�o;8�'�L�#��i}�1�|z��$q~�9�ah�8k��N�|����MK%=�T���	�`l� ; �J�f 	�ň�/R�A�匯1��Ё.�>Ѡ�O�.ap�!N�'��-���[�8u��b�'�Ea��$ɿ}��"�I[�_b0͓c����VF��A	N���Nπ%����7$�nb�!� ĩH�a}�BO(.ε�B� �/�(�S���~b�Y xY��a��`�Xٴ(-ƭ���A�qh�"���T圗O�� a�̙ ޞ�)0�S7�y���1(�$)��%gb�y��r�^p;�`��J��3�FFަ9��.ي��	I1'`r�!���ycUjJH��˅���L��p?"�	kL-���'2���B��5e@���J�2*�LB3K��)�N�`#&ըl���r�I%6�Q�@�#E2%���2���[� �ё
"�9�\8��ȯT���u�Й�$P�S/D"h������ƫ���Q��??��)��B`��!�'_���2��L^8�E�J�w�@H�'İ}�R�A�%[8؃%��,��Q9l�*ܮ�\��O�:�`���!�Y2���lI��)	�'A(���R��J������K���H�f�9���*S�$|�� G �O�Z���Jrc�ͻh[��+Ɗ��+�������A��~Ő6kR���$�N-T����HS=q�<P�/I����*>�2�#'������`��R�
�<��NrY�e*3�>7�<PpE��P�'��EX%4�@����T`��ȏ����RH��,��CQ�F [�l�ؐ(�8*�V���N!�O���
l�	�.ϖUh�1�W�Or<H���:pr��:CFtpB�#�0v��#G��7������:'lԭm.�q�eF�$�|d�ȓ:��-�v��(|I:�dŎ|4>	�OX�i�����B�mAX��'#��9���'$pQs2B����-���(���� �§�k��$�X4Х� �I?s���HfI� X�v	b�	&��k��`��,�u֣A�����B��u�ڣ<i3i�)X��sv団s#�!�z�'�h�S㬘h�бH��!m��`����^�h�t%� w4� �= `��n�t���G8�S�%W�a�B9PW�O/��-�C�<����;&��:G,N�͂Y���(Vʡ�c�
�w��T��]W���R'�a�L��G��^]�9��S�? 4(��)zRh�"(40�:�K�Bn����e/��dS�꓿q%<$�ϟ ��vF�%{�F��p|��':,�X-#b��OXT���NZP�!�GO�q��X��.��W�υ"J�z�n��	�<�Ɂ ��v
�`����/t��d���d҉��H1�AX%lvbqF�H	��HR iĉvt������4=�@S��'�P�0gB�"I���qZ�+#�	�1@)*� �9u�}b`���D�MpD�p��
`�1�˥]��QI�dQ=z��x��N���x�u�_�uM �;P7�G	]�E�m%L<kc��F�Q�y���@^	�0���T�����<t=s4�P+�		u*��a��[��O\�@bXW���A�o��y��R?$�(��͞�A>`�Cu��,��=ԃ�W_��J��="cTM�c�R�=��Yô$͔G8�:bT8�4Y��OY�KD�pT��&nNq���1/n|Q��%[�p܉�k�l[��H�ҍK6fU����� L�0���,רxK%L,A��Af�Z��8�ƽD%4�x4lѝg ����k��1a%Ɵ{�������'.�L���]�Sn��'	ɒCUb��l���&^�}������?E̻j	�,��A�oʼ]H�K�.�H<��wB��� P�>��v�@D|����n8� ��i�f�@��ɬ�#���jAE�������Q�D��o�h�P�C��k�j�8RFT�H-V�^�*�C�#��`����uF �R%\&5N �pH��!�p"��ý'^�yQ�$�F�l�1r�N�/!$�r�g�3��l�?a Ɩi��ʓ�P\|Z�� i~ɡ6HѮ=�DD;�A1���e��7r��- -6 |���ɥ�`a�ա�8S�H�s&�'3�M*�-�4Y$�K��@�?jhD
��&�~]��:V�\�c6����/��H0o�GT|�ҭ��pC�	!D��uP҉[1~��|�0m-,+j-:dI��!����/�&٠��RB���e`����x��H���ڮ+$����%��܊&I⮥Z$��@��{n�+F&a�)O$ �2p)�sg��B�f?v(�3g�B�w�<�I��Sa�}�ӧ8p�,LF~2K�M��:ul�,6����N���'���a�'�m�b�J��_a$���]#{�U�)��p��X0 ���jI~h�B�;:o �8��)�OU9��ҭN�L��6cP���'�^@Q4�䋒�w��@d�^�k��a�EA�O�,�s����	l�M���衫�+q��!��0D��&N̮��m�ҡ�v��������n��Њ'�[,�!bgK]�i��S.~��q��A�#u���'
(�P������i�8�4�)�h���f	.�qC��=VJ�L�a��m���(ض&��;D6��y�VKY�`����[:Kð���ى�Ŧ"Kqfxj�􄓫o�$㶏ҹd!ڬ��*�'<:.�����"�K�	E--��I[H�/.�T
!!�� �˄���(QW�ǞD�j��`+�ON�)I��t&r�i$o�:���+���$A��d��)2hEF��+_H���B��w}!�ą78�:����dAZ�J�� TV`�3j�O��4 �DE-$\��U>q��@���rF�z��ơ{��Xc�d�7v�\��ɐ4}�p�iO q�E�IwRua�*�@��ٴ#ʹ8�viN�,�^��	�6|lp�!��,p%QL��(�=�0�L��p�I.$�8�U(�'MOL=���R�X%jE��%����x$��n	�N�������T��|��"��0�����?{�A��f8��q����1h����
�{u��?�L��6k˧?X�'|L����'+D`�ӂ��C��QFnڭ������e%<�I�v��Ah��Đ1�t12�a �T�6a'I^��'�>��!n�Pܫ��D�t)�8��M�B�`�0��7�����Tq�Ƒ;9��I	FL�} �嫀l-�O`%���9i�R8�s��ȰE���9L��SЋ�˶M���i�6���#S:܍[����D8�9��'��A�Q-�Ud�0�P�4���L<)AdV�Fl�Q����4
>�-H��IK�;�`��O��hа� 
��	r!�C\��M1v�I�x¸���I0(y48���Z�aÐȃ�=������x�ˌ����2' #�J0�t��Pxr�� %@q��<>"y@��ЪNL�Q�ʐ�������F����	8�f��ZC�<l�J��$����jh �� �*H�^�H2���X ��.�?l�p#��:��	�'��<;��
�4\��t��.0TlQ�O�<z#)�*Yi�4��S�c`�E���+���#�l=��#�.LN��%�X�(�rC�IZ���cK"(vl�e�Mk+:��ua��;9�<�"��P����&�2�SI�w��c%��0�H��H=GC��~s�8;��C4~����N�X�xPTOP�7,�)��)礵���@x�Г�B�=�,�����*�=�+O�X���/Po�mPl��5P��`$�ǘ$ ޻#B��"�.zC�C�	Vdہ,Ҩ'�})2*L�~(�QF��$��::�dp�@o>�I��� ��J$ �k�2X�"f�'@[�<�"O.��%�#*
%�!��Xa`�
���[>��"��a�ͫE�F.T@1���O�Hr�%(*b̲�O�q"Y��O�@j��^�d� �c���Jج�*���Z���6M��3�D���Z-cy���%K�ȲI�01�虃�U ��x��S�����NK�PI�SiD�rE��(�[����ؖ%����R��u���9^�<�� +;S4}�O,q����U~�H�Ċ\8LU�|(��)8@n�	SQ~�r����P"Oѡ��rk��0��.}�1�МII�	�fY�?����ڱ��'k��P�ωPmJ�
"A�z3>�	�'8Ќi��2�@|	F[�|��"�%@9��b@�Yۧ�'�q*��M!7����-#�$=�ϓ6�����,!�"1ې�p� �Ht��/-�$a:Ŧ�$��pv"O�)[G��%�,�룆>'�z]X��$�y�( qgY�����@zBd[�z����e_L����V"O��C�&,�DP�AW2|�F	�� �n8&i�=ш��O�H3&6F�*�[b���2�"O̸�-��2Z !E�>���"OvES����8��@k^8<�h "O%:eч:����WJ��?�4)w"O�)�S��5�	 T���z�ԁ��"O�����?�X�Sw�ڳs�R��G"O��߾8{��*Ƒ�v�$�r�"O��#A�>KK$�Kv%�Ƃ��"OH�YQ"���Zq����{���"O\��]Z8�"#θjo"OP �b���p�@��qC��C"O�mj�/�u~DQ���s�ά��"O��¶gC�*�V$e'�~��5("O��&n�$@�Ĺ��A�v�쑴"O�1��랊u+��s	hqh|#"O����ڌ0���N� �r���"O�5�Ůι+H. @��<1��	��"O�P+w�H�t�,��+QO^lM2s"O]��AL��D� b��hN��G"O����E�&Ě焥]0��@"O��&B�b$
g&�h�R�Y!"O^��K��x,������rz(��"O�$��@S�yκj�oJ�^3:���"Oz��"k\,�ԑ��L�!NQ[�"O�v��_�EQ���*�m+�"O"���Rg��C�':�@�"O�!�'��(|1p���-u(
<i�"O>E'��6��)�d�&nM��"O`x2��E�8�!mݺgȘ8e"Oި#7n�!�6l��c��.0E�`"OD(are��%mnUX��K�(90L�c"Ob�8a!U�}�lt"�J´07t��6"O8$�#���x�����B��y!�d-M�CF�,��	�FjK �!����yY�8c��L���n�!�$
cӴ�0���/�>e:�+���!�$�" ��I#�2�~)��I�P��DX.J	�U�.�i�Pp(�?�y"��eVĸ� M�tP�a�M�2�y�@�8Q|s"OG�_H��s���yb�^�6'<����2X0�P�ejɧ�y"(��/��0���R��8u`[��y�l ̸�A�ҰM�����Ț��yB��2�L�˒mT1Fu�͑�ǅ��yRaç1�x:%e@HB�!��\��Py�,^�ND����(�����J�j�<�@mқ	q����N&,ty�H�<!A"��X����#d �&	D�<� ���A��jIK�܇r�؆"O�C�o��؊ӯG1f�:+�"O,��P��/t�Q%�V�2�R-�"OX�*��N.s�`	Cg��@`$3�"O���)Y�(��e:i� :d"O>���'� O!Z��# "����"O�Q�]�wgx�yP"��v|��&"O����Ŏ�c󪈂�B[�o1v\�"O�dx#�L=\,PH��`�U�Q�"O�l�cL��.�0(��.Z�&�8�s"O�9��B�����^�!�6Q0�"O��fO[7d� ����SN,jq"O~�q��
!HK�Ko3����"O0�����F�x��T�?Y�\:B"O�Cuň}2��(�G�m,��H"OHU�Di��Z>�<�����!���o�(`�֕N;�b��N'c!�$� S����ԀO�ٛ6�@�A!�d?����d@�c�&F/�!�dX�'�6��-��ZԸԦˏ^�!�ϘZ0����8��!�T%��Rg!�$
�}J���գ��@�R/Aj!�D�$I�B�)C��U{�%	�D�!MF!�v�%B�I�����)#�F�63!��I�Ɣ�3��.7W��{�ƚa"!�dM-y`f|D�0XYV�P�'� 7!�D�ޤ�y7KE=DX�)��(�!�3]j9�T�1UL 2�c�'J�!���wfNm�A\�-����!��4�!�D�;gQL@���5w2��čN"i�!��; ܙghK��Դ"W��!�ˢ)�q����0�<�1����!�D߳rN��#2�d�|-�r��!�dK4�$U��/�;��5�� �&G!�B�C�8��s�F�V��	���֢P !�dR�Oz��@�f)� Xt����!��]c`4P��5ft!��jV�O�!�ߏ�:�"Q�3rH����}!�J����c
�e��d#�%�'l��±�f`|�ɩ|�7[A�i��ac�\c�oߺ�sԊK��!�L��p�1��x�.��4&��y��\�'�YS�i��9�|�p&ҙ"��1Γ�h�+5RIX�XA*�������b�C7!
�^x�����%X��\q�a�t����ŧ>�efʒe⸫p%�O�'nڬ�1��29i�m��M�*� �a��$Ռ{��q��[/h$\��F����O���������^��33�˽-=�ȡQ��,_���䉥Q)�A���$y�'Qd5�$�7~�>x��R<%�>0�Ѵi(�Q���P��M��#��IK�$y���1m@$[v�Q���þ'�!�d��RA�(��m��]s���cW���5U�+ـ��G�*�M��㕳D��� \v��a�>���B��lR�iS��ܸ!.��dF�H��<���-�����<H����0���6K]�}�X�'�>10��b@�]/�%ʏ�$�=/�.]�N� Q�����Q�����t�1x%h�Yְ�8@��,޴\��GXO
�`c��qW.�h�'癚K����P7ޖx����mCE۶���0��ػ��h�&��t �+sO��y�n�&��oY�i
�?,���T�W�k9�%�H�e�!�$���	���(*�ȵ�c��&�hs뚡o~���R]
9�^}�����	n�H�Y%�R�y�Z'=��#�Ǣ(A��Y5g�!�p?�"Ș9oj��P��*�����:�n�h� go�:��Z\��(���@��(fѩ�Q�Li��X~��)#u�^�f6K�a4�wh�����߱T�12��Q�VLQ)g��\�$xz�'ځi����R�B+j졵��$Rp����'� X�	؛L6�[�J=v+����'�� X2�0M[�3�\.G
�ڔ�L� ���ԅߺ���!)KŜ[".$;B�͚]�L5i0"O��35 ��Q�
sp��OĠ(R��
�V	�U UHP2�Xx�$�
#&p��#���57"��f[��ww����AE�"����k.! f=k��fn朡5�»/˞lrdb� r�vD����0A�$��2��$@-�(b�I6_2�4kD�8(ĄX��� 	�uA�h^�RG�C��#�I7ZP�!���amp
M:F	vi�b!�!��X����@@<�Fۯ+8-r�H\K
��^3(���:�K�B��2!��{��.�4,ac+E�C��i�gl=0�����B6�\�kTɾ?��b���:�����G4
�&Y+vk'D���eO!����)џ|�h(8CbC)_��0I�B�?>�с���1. ��u�?-���R� kRX�;qk^ I��~�d����lM�܄�IlO���3N���pԇ*W^1�  �LX*#�O*^A��ET 
��q�jE'6E�����I.Z⹘��fv��`#��&VR#=��J/�T��ȱ>]l�ih��,��L��	2Ys
%B�^$G*��r'K�C�����#:���d[�Dy�B�wr@<K�ڹ��Q�A�b.��1�g�0r�������CE`v�	�qyR {G�z>��6*��8#U��*-��1$�N%A�!�D]�O���n
��t�S��/_�ʉ� X���{��6=��պ��������?� T��ꚬX��N��W���fl�*���)Z���{��\�h����!m�0Rø08�h�`����U<�Ƞ�a,��&�*�q�� �F�;�(ͨ̢@r�"�w���Ee��+Mx����I����?��c��[�>Q{���wX�̒��Z;1�n��DړN�j���g݆(:�!�� �9.�0��'Z��'Nȼu��a@HŻS�l�a��}��3G���J�C�)G�6D��׮	?r��E: ����wX�r
R87� ��׬�dk�'�8���*�0�����3g$��Aea��"�Mc���ZF�MB��T�͖V�U���,a�$0�'���`�T�l(���Dh$=�ΰ3�L�:\��H͸t��i���4��$��,KC̢h��],w|;���~���I4�Ks��J @w�'��5��G��:�����̈�Q�Zl����
n؜���N�<z���X�t�����M�: ���:�o�5HB�Ȃ�L�J�X�('���J�.g�����'�D�IG��0��D���=_]��®�q�
�)h����e�"�T�a1g`>M̻�ܭ�II&/^Ċ�+fÚ��ȓh���͞�+ȝ*KN2�`q��)��1;��ܨDD<�$��?���-�0&֡B��D�LA,���cvX�9(٩��Q�cI�(Y���D�<�(�B%�.f}B9�"@%�$�F�D�h�R硊�(�h� ǎh���8t��v������
RF�  ��������P�N6�O^B��G'��4��X�rq9)�"Q�vh2��ɶs���Iԫ�(
F0t!�W~ H\������Q좀�䡌B
b��8\&�YUK�K�d��ā�'	T����S�T綠´��T�T2�6�8F�c!��
���:�Ҩ��"O�B¦ ������"a��D��C��"a�P *�/z#|%r��	n2�������"�#e��ʓ)j"���*ՆUvphxra*;B���I`��|8��
K<��+0앙W�H�s�o��p
�a>�J�!��O&8>}�v�	&Aax����`A��@��v[\$r4���HO�<X!�\�*`@@���)' R�l�@�,0����>䘲�Dr@���;n�BቁS}B�He���4�.3/����UԺ@�aOO3�N,k�BZ PzL�h%�K��O�l *�(�@��<z�3u�L�"O��҂�k�4�z��Mޘ1a�K�(+d���S�V����͙�w�q��'N�E�o� ��E
4$��X��+�'Ҡ�:�8Sq�a�ïMm�)�ݴ[��1;'�4Nx����	�L����ύ+SV�P ��1j�����L��mN�Xp�Z�)��� (�(}�(�1vj.D�L�A�РR"�l�HF�uc8�@�K D��!$O��J��1Ǜ�~mD[�h D���#�^�A1����fL�D�?D�$2��/45d���)���Ɇ$<D��C���U�ͻ�a˦{�D�#�<D�����(&�V=H��K<H�+�:D�L!J��,
���P�p�P�7D���7��#e�j�PL�/&�@�@'D��dk�;^�,�KC/ډ|��9��$D���AbI�(=~���75S����a>D����F�2�&}K���Eb�Z�h9D�|�����-XA���=��d�u$7D�,#v��']�8�r�@�: ��0Y��8D�83��Z�2�|�%��X���u!4D�)�*ʱ	�%�0E��  ���3D�x[�MW�U���)})�չ6..D��YE⎡��`�k1}����/D�� Fk�$rx�3�F�|ڡCN#D������J^�M��%��U��<D��smB&>�΀�`�Ҥؚ��fd<D�� �b�,�h��*Q,?��2�"O���iѫ�֔�j��*�i7"OP8R@�$mV��eI��"�"Ox�Df�6f�`��g-SϒR"O�j�C۲f�R�+t��uˢ"O��0U"Ϭ{�2x��j��L����"OrZsCY�@?D�pQ�Ɓit�)��"OH�s��ݔ+)T��K�Kmȕ"O������h����)UT@��"O d�X>'g��I��)@��`"O�\ʕ`��Yy���rn�jj�m(�"O�ъ�l� ���#G Ge.53�"OT�DļR���mâQ�!�r"O"���GK"�\���
J���"O�p!DI��j��v��p��Q�"O&��"IJ(���ʓ��_�  ��"O��W��*D*b����,b�J���"Ob�؃'�^AH ���
NV$��0"O����NVB��0Q2fEpQ��"O�m�#`3�����$��!�"O�d��AX2�院E����"O2�3s.�)V.5�1�޵$z(xt"ON�ģ^�U�J��u��-V��"O ��E��O��ȱ�(b��s"O����ȭ9���G�B�F�H���"O�16.;5}r�fY���s"O���ZJDk��:yvf��w�D:�y2�,:��1��җlzL	B�ݗ�y"��#&l���'k��W�x�%dU�yr����)�!�O��إ*��yB(ɱ]��L���1ld�Z%�[=�y��@5*:����FHZͻ�CU��y��	&���jR��)�~e��_#�y2R�Dݨm�3�A�H�g�r�<!��/�x'A|U��E��M�<�PKK%W�T��
\>eF�� �A_E�<��,
�p�������C60�� ,�B�<���ɩ�9�*�Ji��;F�g�<�n%�^LJ̽ZGh���i�a�<Q���P8����8rj����f�<�1��#;��<�7I�jf��Ѝ�`�<q �$?W"]qGI�HR諠��^�<iƌ�d)4�q��A�&���[��C�<�׫���|�[��ԡ!�ɹ��f�<!���F� �1-��R���
GE�<��E�}$m��A���Y�"�N�< ��P$�S�Zv|>!�0�HF�<yWgN�@QN�8�V�+=����ZI�<����c����@�"�4�p%H�h�<If�V!WٞTZ1h�v���@4�g�<Y���"H8��!cٛ�j q��e�<��>}v<J�MG��A��\�<�P��ys�E�4���`��X�<��ǹbS�} 2��/�aC�XW�<�ʋ�I�Lu*P��R��(f�J�<q�e��9�@��ϟZM0,��cO�<��W�J���`�jb���ԇDm�<)T$N'
�y�!,V	�D�%�i�<1�/�"h��D��
éZ7|q���S_�<��ˇ�+���L],뒈�W�KX�<�D��!<��y5�˰�:��f��Y�<�!
Q�L�F����-�:�S��c�<�f�>	F�`� F�`z��s@�Gu�<�蝒M��a%#x�� 3 ��J�<� d��#&�j�X�1	R�3��p"O���jO�!K�P�r�J�n��j�"OV��DM�?)�.M����1:���a"O R�}��`���f���"Orݲ�Y�r�e�'#F)&���1u"O���3�2�yU�
M��+"O�	��F:KA��&c�4:�Թ�S"O��V��*���v�3h<����"O|-�f ۮG&-�����!1�"O�m� �ݝHc̍��,�@��P��"O2���/3*ܾ ����>� q"O����.,֩��a_8*w$E�B"O6I�Ζ
�D���@Ȩv��d"O�0 �O�(w<CШH�PPS"O�H�!���K�.�b���<WK\e�u"OQ�M�(R����F�Ք%K ���"O^젓 Q���$.77&��#"O�����!3�T|��Ɓ&8D�J�"OE�� �{cVܩw��/�izd"OА�BC*s/�4�&aM�#��q�T�I��^l@u΅F�&�Ad�Լ.���Ɂ ߒ���X�J,"�*w ���$|q9��R����=?E��K��8מ)���ѡz��F'L[�V��c�����������|:ec�y��Q�����,S7T\9��_�U!���?ib�O!��R��D˕�˘ő��F�}�ޥ�
L����b�C�)4�	5�ӱD���6'�P��NV�W�Z�A�JE/кYM\�cM|���)��Be녧�;��t�a+����v}��S�[��)�<�&�Z�9[hI���"OD��J5��Eê��ɤ �)�,O�Sm�O?��t�ҽ
"���jH=NUx�#�H�,٣(O"�0E�-I~���
|��Y��E�y��b�G[�n��t��]E�Z�� 
�6{�1�FNW�$�	IL�,�<a�J�IrN,y�'	�N���S6A���4Ǆ7{�I��}����;h �$���T�i�CB~RiB��8�{���Wc'j����?����)Һ�~BK%y�xl�}�)�L<�A�]X�90��W�q�F�
�E�!ّ��C�S�t�i�ē�. �w)E�+�6A�W	Y�L�9���z�P��2L|��d�!�~�����x|�q�焘/L� P�L5��Q}r�G ���	Ěl�rCM�P���0�j�'yT�a{&������4�M���٬kF��D��'���
B h"]!�"��Ř�'!�6�"*��O�]>�'o* jE���6�晸�c��2E�49�B V5j�c3I�	���Oszx(a�|����[��rd�B/9<>��X�NO.�F�tџ2m	w������Y����u��'����e�OM� ���Fk��x ��D��`M>0�Y:D��h����Oʨ1���1>�"L�MW�(�%h �l����)��������YsO��M�g�I�::Y)�J�A���R�[E��B�I'|�Rm�WIG�@T�a�ق��B䉪�Z�Y�'�2 �X����~B䉞Fe�¢U>�JU� �1O�zB�I�%�(� �7,�0Y��� #�vB�I�&bR
����2��!{vbB��3+#
���c�;%����F�D#T4B��hn����Y& as�EbtHC��&T��)2�m�:�@(��mGdB�	�~ ����lʄ1��.Jo�2B�ɽ9�>�c�,�%S�XQ��O�l\C�	3J��m�A �
q�VA���T8C�4p�tQkr�5c�t��.�a�C�I4Vjh	#hܪƞ0�d�9p��B�I;YꙢ�`���H��E�\�B�	�?��Jp/I�[f�tE�G	X��B�	(n]&�8�IG&W�t	�dY	KlB�	�Z/ޝC�
�'��0�֬\n@B��+H]��)T�"�M���R.�B�I>H���#�˓:��' Q6��C�	�Ymd����93���"e�(;�tB�I�"0i���.5�KZ�i�P(T"O� �@��l	MÖ9�L�5Dr���"O�!ص��<�,BFƝ�]���p"O^<!��64^ ajWO�b�1R0"O�l�&S b�.�1�&�Bq"O����2���2t$�3v�L��v"OL���$At8i *
'h�Lu��"Ol���펩�k��,b%"Oڱ�����9Gj�X�ZP��"O�`2�ޑ%ŤTG�%r���"O��1m�$3��3f((^�U�%"O��a�.L�C@�I�D!�����"O�e`���&d�j @7��}��"Ox�{�+?gt�S�E�;tC"O�)X�e�5nZ<��C���E��"OP#�B��)���`%��#4�r�"O�p0�0�
���@�6$��r"O��S��)m��Iס��s���F"OF�ɣf��E��i��M��H<D�hic/�;^�
��"��`��D�#<D�t A��7a����-t�j� ;D�@�2��	O�$<:�KS"L���o&D�T(TɎ1.�N�Z���,@�F�P!�6D��kp��)���H`HG��FA�vd/D�DЗ�\>2Ш�W/��Ny}IWn-D��Y��'OL��ӔMؒd�yC��7D�\�Bŋ�\Hr���R�C��<��3D�x��0�(Vi݂[���z�+1D�t���%sdp
f$@95��,@��0D���@�w3:l�*˾N���j#D��'m��\ݐ���)V ����$D���%�⎁���	�U��=S���y�B1��lK`���62VAc�>�y�&Q�%�hit��E�ĵ�R�B�yra��)D���Qe\�5�*`#���y�H��E���S+.F|)����y"H̸t���d�Λ;�x��1�y��;k�-����+�Hx����y�>��|z�ԙ20�q�@(���y҅S<I�@T �i�0���z ����y"�5G�~��7Ň�u�0�W����y��@5d�tsf�H�q�L� ׄ���yBj�"��"�E
�p.(x)�d �yRE\>T�PH�Sƀ�~?�]�Bٝ�yrJ�%6���
�'�*.�Ψ��9�y � 5WH�,?*@i�f(���y���rz.�Ȃ��0P�����ܥ�y��x�0��g��]����hTjB�I�B�^��)G��ɉq#ֈO�,B��9\�Ω;��T�}����!H'+<4C�	!a� ,�D��%�)��nєcYC�ɖv&�:� ��� ��/� (ЮC�ɉA&5���;&Dt���(�!���p�r����;|n=�Al�&v�!�<��Ec�D��h��E��(�5:�!�䗌P�<�� �O��%[��22|!�$5 �<�aR�{�����N5D�!򄄹��Q���6m"�5�g!�D� JR]0� Βu6���l���!��;g�a%�� %�ź�H�@�!�$�r��x��
YY0��� H!��T; �,�!���WrD���ɠi;!�D�Y�jI(�웪6rj`����u!��P�B%�h�r�yt���h�u�!�@8\�ؕZd�C�c_���᠐��!�� d�*�d�`0���0�0uc!"OB�fjK�qU\��g��4u�f�"O��Q I�����5)�s�8P��"O�,(��/q�1B	B� �	3�"OrܪbB�V�Eb��oX��S�"OH�P��C�Nm��a]lJ���"O�P�Ί/X���e	�<��`b"O�1P��X�Y�B�c���~�e��"Oh��")�+�C#G�X�m�R"O2�xd��'p��Ъ��+�X��!"O� ��Ξ�|P� k5eGN�Xz�"Oꠠ�	[�b�dp����0E"OF��F]�9Ͱp"!��;XN�XÀ"O�jv%*+���I��d/�s�"O$����XɞA��Hw@�p�"O��w�҄N/|5X�&�jb�{W"O��R�Ղ/�h��G�+�h�A�"O"��cL?]���	D_�@��!K�"O����T�9��9s�]�.��5"O壑B�!'��0�UK�0n�@p�"O��3q��%?J~	듪H8\ʄh9�"OQ�0g�D�)�e
ٯP�2�b7"O a�g�S>
2���DXVu"O�y���2�����)MH�;�"O��V��
]���"tK.?΍Q"O �����VE�e�D7�X��"OMrtr�!�IE�:�9�w"OJ�t.6bF��VI�	%bPAP"O������dNj�s��J�>��p"ON)���I�th��� "/XD|�"OV����6"h�=���=9t�I�"O���$_�\�$R��-�yr�"Of�3�I6	gp%Z�� +f+*e��"O�i����9�(h{d�0$T٩�"OV��ɷ'<nh ��v��i0"Or%���Z7w
���)ؽX�"OX�{��F�Ne��1`�\(RN���"OZ ���3Sy�	�,�S<�4A�"O��R�9�6�B��E$�̨"O2PrD�_ި���h�*�0-�F"O^}�0$N�3`������ z����"O(-�ǃ�,v�~���?�V���"O�a���1鮼�B�޷rDq��"O��G�&0�^�0�o�&d��`%D���c�N�j�Z7IZ�����>D�8SN���~�P��\�4qT�1D��@�h�?1�n�&DN�"߀���j1D�T2B��/+t~�d��<��%.D���CD:�N�x�oI�0�3��(D�8��2̔��9��9�L*D��:���:6:
��3-�`\�q��=D�P�u�I�p�zX� ���C�c0D��y����FC�Λ3 ���'�-D�#W*�r)��Y�DO�2�X��+D� c�LD�n�T (�`BK/�lp�")D�@��cD���j$�2N��XR�e3D��q�V5>��if�W⌘�ס1D� ���ڴ?�`a�7	��j.EhC�1D�tP$�Mqx�I�ކA4�X.D���gh���\ F�Z`�Q� .D��"�]~��$�m\�&�P�2E�)D���p#N�>��0�����T*L���i&D��0�_17��T����D�"YF`&D��(�B��&�|$qQL��M����j(D�� ���$�N�@$|��D��l{� H�"O|�����C'*�i�Л*H�"O�����j�x�1�Y�Z�I�"OT��T�A�M�e���P8u,�}�S"Oq" ���b�<�҂a����qV"Ob����� Z���$�܁vfHL�s"O�uA��WJʩ�P�ZK�`�"OP����^�f�Ց�7g��ɕ"O�a1gHD��,� ̚�`x�p!"O�u!226���M��y[h�V"O��S"._/n��Ȳ�)��c[��"O�EIG�'Tq0���#o �]K�"O�D3���	q��H�A�8sz����"Od��獌�zd~�ibō2y���"O@5Y�D�R9�1�ń2�����"OR����w�A��֞.gQ02"O���U�[/;:�ѐdפM�
s"Oi��bX�l̚-�S�A�=��	�"O
(g��,�j���RH��A��"O��+��B2{�v�)o�d�^�#�"O�,e�o<�NI�[�<�P"O����&ie2Ѳ��Z6���ʁ"O����K�k78����؟B��q"O�����P���\2���;L��d��"O6��U���j����k'���Q�"O����ӵe��� t���R����s"O��
�Ɏ�^��s�H�""O�`���[�"�pH����F�*�x@"O�����y�����EzFv��W"O(p�`��![�	-J/SI�Z&"Oh�:�%�~ x�!M�	(��"O0�4߲n�Ȅ��邹_
ts�"O&P
�$ֆL�x�rʛ��t`G"O�l0�а&���("� ����"O$HqG��*+�T���LG1H�d�F"OHʦ)���(5�E
ˀ�ɷ"OT��ua[<�̊�,әVz$S�"O�١�)��D<-���,=�9k"O��ee�&;Z ͓f,�*����"OYЀ�V�b�����
#'>��"O$]Ц�[�}�^e�R�Յ`�"�["O80ڇi�>m�&|�$W���(�"O��˴�[�1$*���cƶ:�0�"O��;a꟨$lM*� �T�L�u"O�"T�Ç�0-`�.-���[�"O��93��g��K���8e�`��"OB}H�m3��ap7g�v�m;S"OZu��� J"�([�W���K"O�x!   ��   �    K#  �-  7  B  �N  �Y  }c  *n  !y  ۃ  `�  ��  !�  �  ��  ζ  �  V�  ��  ��  a�  �  V�  ��  ��   �  d�  � � 1 � � " a( �. 85 ~< �B 3I zO �U \ Zc �j 
q Mw �} �� �� 8� x� ɚ  `� u�	����Zv)A�'ld\�0�Hz+>�AI��m�2T����OĴ��f��?Y���?��FJ%L+�}�`�:b2y�4K�,#`��8��4]��)%ۉx�:��W���8<�n.XWr�iS7C��� �+�P���>"�i31��$��db�/�(X�Cd;h��2a�^LG�I���h�'}��6�K�o�$��&\�J���Ǒ�%��isPc��4�6��5D�x�5fA�xʘ�n�qG���Iȟ��	ş��6�A��&�����0��1;B��I���	�M�,O,�DY�^c0��'��-C� G���a1,U�⌁p��'Eb�'%2�'��KE�u���	2���gK�c��h �ɱk�z�ҡX�̀*���<��Or�IU�>�#��U� HT=4?�hKv$:0S������{���?Avd�9:2e!�"��y&	����f&ïY*4ɰ��		�?��i!B�'$��'.�$�'��S�c �ِP��5:Gg
4_U�m�ր����J�A�MKG�i[<7��OzY��L�8\Q�iUY�!���~!<ey�F8'���% x٨<*��"ғU��P3�E[��&P<lT�;�u��])f��cL��@�dD̪&�ڠ�u ��Z�P�8elP�AG��Gu�Tl��?�0�OyH�Ye�*K����q�A�&������?נP�ܴD<|<���Ͷ��@��n�8�K��K�pLTe�ip�6��Er�||���{��ϻ!���ˇ�@�����4�v)h����H�E�h�ǀ��9}>	i�3>l��D�T<h���礓!s��5�fN1�^�cQϚ��U!ܴMϛ�=M_���c� %��4�Y2;T}��Ip<���fC����A�nu�h�b��QҬ`T@��8n�v-�O�t��m�8\$���5BY&Q	j�����k��I�e��П$�	ԟp���?�J�W1U[pݓ�����d�� � ���	?*�����ן��'���'=�Ɉ��:��?j���3%�~�zɥ��6A��p��]r�%��'O�{��QȚ��.��cfD�d�k�^ѱ#�&.�~�� �:81����6*�{�{��N�?��iGN�d��Ъ�O�ysb�A"\�����IS������ޟ@�	�|b��:�TL�ǧ�p�ĕ���D@����4!���1d�ĲI�[����("�i�2�s���qG���%��埐�I�?!�,�*��ų`���K�匃y,��S- 럸���]4��p�����$#V�H0S�<��O-�ӫ�����~|����S�B터�'���e���X�ANgG��c�AAP���B�SLJ����6 &y1F��1h��P�oMb~2�^-�?A��i�6"}��O�D��½ad�s�%ܧU��M���O���Y�H\���&*ҭY�,]���ɕ�M�F�i�1�����ߘO�����8,<.��v�'ab]���E��������hy��V�� Yb�G"sh6HC���/}Ģ�QbH�5Z��;��7#�@ӶZ>]�S�$��'\j��F���8X;�I
���녢�$~�B,�R�o��c���u�^���|gb�k�uλ;,���HC�X�N����=X�(��4.��I)D�����j�g�	+vHN�ӡ��,":,�r��:Z�nm�	����'����>CiP97l�ˑ �0\Q�I�k�Ty�@d�8oC�i>	�SayR�܋��\B�ɔ\M�0�I�j���sɫ>a��?�-O.˧���DA�}ՠ)ɤ옂6�~	kT�줃��~�T)@`kڪ��y/�H��P�7%�<4Z��a�Z,"���
���wT���㏂T�FQSQ�isPu���F�ø'�<и�:"]��;T�ط�6m�`f��?���i�N"=�����6.F�P�W�]Âe��-B8O���'���'���$(�D� ���	�Y����L>YF�i#z7M�<F�j��������_�kO6��b��lS����mϟD�	�;�d�����t�	�M �,�R���U7�X�4K�������^WRM��j X막�R������	M�z�r&�#Dz4��A�%Wa�-�
5}B,�(Bp�*��@>aB�B�$߰	�de�Il���BU����,��HL�i����j�^y2�'"�'Ka�T�Ni4dz�m��Fp� ����?���i�FlS''6-]�MS�V�C쬼:�Eb�(�@gPMZw%֑�?!����ÓXA��$L7)�QK�h�VZ���G��"0�p�d�Ot-��lW�+ �K7!@��JwNZ����^>���ўLh�U���("dd�GGT~NӋ=�HP��D��+�:!�����	�l� l���O�����R�M�n��&Z^J��O<�d�'�6	s�p�'y����&؃<�Z02V@ƓK�h�$���I_��ǘ'��9��H[�A��@r`ǰ19�=*.O����Op6��O Dn���M[�E;��w%��S`cP�eԦ]ё�]�����}�|��<a�*������?������F9z�TǨ�.	�����#B�D����E��to��^��Ey�ǅN�DG7�I�S�A������3Aᄄ�pnJ(a�|��F�� 2���+oG-�$��Vh�h���ޠ��,��wM>@�FKdb����4+��;G�ip`�'�(A������?	���?� ɂvd^'�Dt��� o]��?1��?���?i��L�hZ��C�OZ�8��eY�\� �W�<�S�i<7��O��nZğ����?Y�O�|iɚ"!N>��w�.*�t�"�'��)""�'���'B"��~���?�B��x<0���l^Ĺ���2)>|:R'�i��A�	�K�>���/���#�<,k��㇌�$r���a2�K�E6��b�F��u�2LB�m&ĺ�X�å?���L>Q����4�x5)�)>�����	�O؁�ɬ�̼�޴�?�(O"��;��d�<%��PvXAb�"I�I�ڈ��"�����O�H�{²i����'��$�$`��8����>{���)i�}��Iǟ|��4�?q.Or�-�u�I��Ґ��\z��;3��5ϔΟ��	��<��	ܟl�I�%π�+�˓��D঩��9��� �\�b�Z�%^��'W��B�f@."zk���ݫB���E�/��U��F̃L��4�D9�8%;�AW�6�4�r�e��5�ñi�ءN>A���x�޴o7�bq��b��E�!o؄IУ�e�$�O�=1�y����;V��c�*�>{�*4��-�*��'�ў�S�M�%�!�� ����5COҽ�4�]�x#��]�,�
@ �M������|��"�>*S؃tp5��OO�A/t!��?�g$�[��d3_��6���Mˏ�T �>L>$���� QQ�DQ�	4�I6�j��dO
(i��R�nK�V���h#jČ(S�V_]���6�UfJڿ|l�|�\z��5~���$�����il>��5�
Z#,�{� ���XN�O��,E�dņ�r4L�a�b#H�,����=vax�i�66M�O^ynZ�<��. ����)-FlsBl�)�M��?�m���ԦX7�?���?Q��y��!F�"g/x"�űeM�
y���7<*6M^[��b��|�"�Ĝ�s�̘�F-�*|��e�)�r�NBU���Qǒ+HXJي��(���<n�TX�%Di��SJį4��`"Ҡ���~��hCݦ��ڴ�?ه��#�?y��,O(�$�(m4ٕ�L>��I��ǀD��D�OR��?����?aq�L���'�T=jbj0�Uт�A=�r��V�ia��yӬ��<�������ix�� �&fR.P˔�&n���Ve\$	�����O��D�O����?������UUĸ��"B�X��2���H�⌲1e�KNb,�B�%jI�)0G�0!:8Dy�f���D���hsΥȔ6%
{�hϷ��QgQ�e܄��g�-�(���ϐ�R�'�.��hE�h[b�c�E�h���b���?I��i�#=���D>����Qg�J����.;�{��$E�Pe�݉F,^�
3� �g��'� 7�O�˓>c����i=�-5��q�X(�L�Kԣ�V����<Y��?�O=�|��<"�R�I%�i՘P!�8d�\��b�B���-�H�c6�N�3��ӐJ]DERBFތ(݂��p���4�|��#cՀ�s�ٙ8@*�Ik&F�I(J>a3k��3�4f�	�kh��և]�bIc퍢>W��OP���[hJ�+E$�hԑw#��t��'�D6��<�^!`Hdʩ@���Y���nZOy�#�p�7��O����|ڠLʢ�?9��-f��]�ċ]	 �pP����?i�B�
-9c�
�
�����m@�d�p�c7MP	:����+�X%�H�#�B�rEڿB��j`�7?���o�F׀�1���q�2d@�����4�DBФu�����(u0��5�����$;��j�|)D�d;�X�s��
.f��"�ؙS�Z�P��'pў"~b����8�V�x�(���@�s���0<��4���$W�/�X��Q?,�:��b�n��7�Op���O��r��XY:��ON���O���1eMP|!��	J34+r���Y_ȄR���d��g�=""p`�a!�S$C�����O�Y!r���M�frv ĈE�I`�F��@��U�Z�]q*��d�A�h�J�|��䟤t|�̻~�rDd��\3���=[x�zٴy��I�wDd�D��p�g�ɪ ��!)=O��Ӎ�?oWl�ȓ.;.�����$-Ö�W;'!���I͟ܒ��4����<�AY1���1�H)v�B�S���?1�iD��?���?��5�n�O��d�O�(�`«�z ����ZVH&8�t�Ӈ�&�4�@�Tux�`�Р WilT3	�Ukn1R͞�F�xZ���(�L`X��>!��5��ȉ�e��!��2J>{�k߇�2ڗ%a�M�W�'���(Q�0�Ӻ��/d�T�'/�(V��HC���4�J���՟��	t�IUy��4��[ơ"I]�'��8r5Cۥ���O`�m��P�'��$��jn�D��{�x��L�.��xB��R�-׆A6C�O���?�����F��� ���ƵS1^i!��ig$Q	`e�81޴Y�H�oaLul�'���`�;T ��2`J��x��#�5M�x�B3��6�P��ᄚ�B׎�6�,%�=A�Kğ��4E�I�����v�	R�����QB�O���Г.�D)�
*J�iA���	z�����4f���ڴ{:B�P)C�_j�9g�i����\�Z۴�?�����iCr��Nt�t�� -�jĉ�"�S��d�O���.�"*p��?)+��#�`�7G�"5B�HP�|P�X�'W�PA�&�5����CN�"}BSo�tb~�PP$�;`�T1ЁFX~��H��?)'�i�N"}ڛO!v-��@t0�*�"E "��@ۍ��)��'ˎ	�`a�bm�(��C��\�?aǸi��7m+�S�|��#�h�C��QE�~ql��D��şp[���3���џP�	��;!�)�r*<;� 
��ۄQZ}*3���:�ꠥ�V`ѹ�#�~���O���$��ꓯʕ}}$��)N�X��ǖ4�f���`!Y�(����ű2lEK��I���Φ%�h��w��X�BN3<�Xe"2��8ȅSûi@��C�����?e���@,H�C��5�Jр�QD�`���hO?�K3�s��h�D�	��3B�	ݟ��I�M���i�ɧ�d�Ol��!1�ޕ.l^�Ywɍ�?��
���)��@f)ٟ<�I�� ����u��'�R8� T�WL;�aP%Eo����ㅘ�,q!A�����j��b\��?)���N�? ��B�~�dQ ���B�3&��:@6˖��a��I�Zr����"N�T���Oν���j��	x1a�Ov�xfюq	r�'���d;§�4�)I�t�r@���B
D��A��y8��G�^F�5�g�шB<�Y&��R�4�?Y.OZ(���¦��	��2�E�3�`��/.7�T�X�$���O�� @j�OD��v>Y��7��!��H�Bܠ!����x���E��b`lQ˖��)ΤM�Dΐo�Q�T�e���U@��ʷ��n����-Fud�!�F��e��z3k�w��aW�؂�����z�	����~��:k$��B�@\f8#��^2@��C�	#�8���`ا0�t�j!���|J�G{�OZ&�$��h�D-k��$T�Jԣu�'/��PsKu���d�O^ʧ"����rsޭ���\,`�����K�.\[~����?��m��?�rI��cJ%-�	�Ҷi��Sn�4#�=t>,�� lM8~b��kނ4<�	�A��cR��4,����ǟgxL�)����Iʣџx�T��l����cE$������3g�Ov�o3��'��Oݚ���/ͯ%��`�$ӻ
9<	I>!�����?	�����%tT(#���V���
#�
;P3џ�����M�L>12��2#1 ���%��P:U��m��'�r�'h���B��gM��'W�'��N�"���م�/X.V4R��Pl�1O؈3��'q�0�g��F ��3�ÆzG<�yB'Ν�0=q��ۘSĵZ&��Yp����N֏��Zt����m�g̓{�T�u�L?N�
�HP(Y����*���wIY�_���!'�I��䑩�O< Ez�O~�'�����5Q��	R��!&��BmN�2��'b��'��.�~z��?�e%ŽNt<�I�$�)E�n=Z7
���kP�M�D%÷B��y�E w��i)�	�5�H��)�05�l�㫗!Ҁ"`	��T�*�N
��z���g�t�f��<�A�na����X�~�d�s���ʟ���4Y&�6�'��	�8��ߟ(�O(@��қ~6^1��L��f^���'K�9 �0�F-���.�p�IK>�i�:7-�<���S	��6�'Kb`�N��YI��&84h��<��'�ꜩ��'��5�F�(�'	1O�T���ξie�P�2��R{�婱�'1(�
���@U) ���m6�W�A]�Ȑ	ÓF�d��/��i,�Qc� x8)�@`D�r�2܅�9�v9�f�-'� �*��2=~��I��?�$�ӊ7�:��d%��:Ѡ����Hb��nՙܴ�?1�����^�@
��D<S}�e)�M��ܠq���?Y��D�O�ű��]�fh�DDæi�� �jU�+�H���+2&����I�,,7�J!i1E~�hTjnj:�d��8�.�Y���/�De v��2$]��ڃ�O||���vm%PUC����|��O�$J��'�,�O>�r�E��*���E�� ��E",D�8��N;]=��b섖5h����h%ړ�?�3� #�<i� �MDt$����0�Z�+�4�?9���?!�`��l����?I��?!�w�z@Y������1�8}�L<b+I7ƛ��'r�Id�S�t��3ʓ2��)`N��PVP�ӕ�_�t%�Ѱ������J��)iE��$7C0�d���9o״�3k��#���<�/}y��?���O~���1��咑�C�<�c4 T�f��˓�?���?I��>A�ϧ�?q��8�%�GM�}���A�L��`�ؤ����?���1��gy�_>�	dyr@�;A�+Dj�k�����cR ���Q1�@�R�'�'O���'��7�.T0�⁪d��ɒR%^�gW�q!�I�R�<u�v�F� �y���6]��"�O2e�Nӧmh���˲~-�,+��_\."�OT��geXb�A�լPD2�Z"O^D���R�m`�ì�R��U�|2ClӦ�O�E���O����O8��t�Iw:u�CG¿=�����O����Bq2���O>擃@V$�#��3Ӆ�d��䨱��=�2QZ� O���	�I�b]����<���P�\�F����L��,�� ���1h,w<��Cq#P *XC䉭g��J�Έ'���Ӑ�	5uq&���Mҟh+'2z�T�2!� �4��e/�$\��0mZܟ��	S�d��-p"-F�Zh�����.�ZT�)�x��'�Q��'�1O�3}r��2l���	�N�0V���򄀛����U�W��"|�0g
j� 2�@#5�D��5�FX~2�ʁ�?ɣ�|��)��XH�G�'}�A�ȁ:6Q!�����=�b�ʳ@^����_���'a|"=�t�מHnv�D��qf°rP�
��?���?�.�r��ЂW��?i���?a���y��=>.~,ʠ�ǟc�^���G�P���d��;ݛ&j0b�|����$U�-t��5��C]�@0��L�'���`fn��7��p����Q�h2�P�O�Ȋ�`��y� ��W�
�q��Ɍ
���0�'w�I1T�$�O��=)2��+j"�	S��5K���ف�	��yB���s���5Kρ3�P��0��;�?y��"L���ٟ�'uV@S���n�ʂ@-"�L�p�[�9c�����'Q�'�Z��.�O��~>iR�aCjJPܳ��D�)���#r,;V�b�yF�H$[4���a.J&����HPJQ�hyfbģ;�=y�LY�(ʞ���!#��c�j\�՚��#J�p�b�l��G�7�/Q��'�;�fɜ������W�QpVmF4�?y��'�Zx�@��3�n�a�ۍc�t0�ߓ��'|�	�ԍ�2��v��[@d�N>��i��'�Bt:"�~:��m̞���X�o�t��@�ԝ9��H��?�H�:�?�����eU6U�(�#�P���ya&��);Z`��dR�Z~%�a��e�<`Ce�r ��Dyg�&5�����W���I�CF~.t:g�&C1 �XbW��!O�I/��o��ܓOP�7�'����	���r���J0i+�m8��0�Oj��&��Q��e�q��rj�pAs�D,��|§�'�H�[Ri~K��8#.|b�x���DܒhG$�mZ���	m�W4�b�R��c2m�#[��C��5�2�'��}Z�cх,چ�sZ�2��B�U�<y!���IF�!��<��R��t��^�[C@�)��%���=�";d�߉p��ۣLQ:�f�O�(�$�O�.�Q-`Z%q�f~��?���|��I#�	��@iFЬ�D-|�!��Q�#�FM*B��8)(��gB3�џh����"�v����Wm��8���?��7m�O����O6�W'E
4,j�$�O�d�O
�) ��:2�ֈnTliz�`?{�	�$�7%�5��,Ge�T:Qc�|��O������V?i�X�L�X%�q`�pz0K�K��u�,A��H�-f~uK���4P���|2U�Ωd���Ɂ6��˱���T��4��,mc
$��14
�O�b>c�x�q
I���Bb'V>�'�*D����m(x+"y0�l̢[� �[@j�<q�i>�%�`J�!�2����D���<#�T�#B�(:�^��W�ڟ�I���I��ug�'O�=�f,n�=�p�&�?�J%Pd���$܃3�?H-��j/)Hq{!i&�(OxܓsɄU��e:P��L�(ụ�	z��!�U�*@,�p�H_�as�!����(OB`P�����]�ёWir]��[�i���<�O0]�u/��7y���R3	�t�"O��f�=7xx�J⧊wb4��|Hu��O�!*A�j���'�$@�Ά��e� ��|��C�'���F>^��'D��(�\�c<��d��bl�h� �!�3���
ǩ
�7��e�%e��|����Lq��=�C�D�p��q$
9>�E�.�	2e�	�1ʬ$2e�R�A��@��I<R�d�O��p��|C"��Uq���)
.o�^�{��#%�k�M)*�	�RU[l9�Oh�I�Z�D�z@CC��sW�\�v�D�<��f��?����?i-���'I�Od	kBj��B�Re��W4=/e��Of�$W"�����ݟNyZ�
ѬK�B���j�(�
A�r}DŘw��6M����Gߜ:�^��'�z9��I	68�D(²/���6o%N�HX�C�WjT�B�SU��+uν[a������w~"���?����h���I�b��H!ڮA��j�g
�[�C�	d�Ҧ���Cؕ:G-ɀe�d�?Q���X��{f�QZܬ
%�	2i[*to�����IПl+�ͅ�P���	�8���X�;ٴYX�Mkt�҆R�n@b���ҝB�����p�rI2�3�+l�yc(�6���Q�ެ8Dʑ�S����$F	Z��} ��󤟳FXZ�˔2L��
4QK���$�O���"�	k���FA�R=��j/b|q�
�'(I���`'���AJ6#m�[�R�����4����<�VhѶ>u2�	 �P4 ;��@L��r����G��?!��?���t��O��Df>}��	(fȲC�T�T�.l��K�W������5+���96�'�rDFr炞T�!���]�Lk��K�'
����#:���S
̼.DX$ra晑�O~�B7�y.�pU��9�@,�61#�b�'(r��'�'[MP9X����@�:B.��
�A��F@rs��D� �2�РIrCr�&� +ߴ�?	-O,u�7Zy�S1�����Fֽt@�k��r?���<���?��k��u؆�Ѝo��%��.�f���[s�l����f��hq���0<i��H�7�6��&F�;�^�Z�)��t[t���� 
y��	!2 ����O|�e|a��H�6`U� ZSj�D���'���(����$�
��p�G�����E����%��)��E�O�   d��O�ʓT�±(O�Sn���'`P1���Tr<Tz��\��!RP�'I"Ɖ�M�>��TI*!���xub�O>s�bO�$���*��ns����'?	��F�4����ST0���R%2���2����5�Y���ϵ:����p1*���OP�}ʜ�� n��.��`@��U#�d4��"OƠ3�$O0n��p��	�2}z��I,�h�B=	F㕸n�2mё����t�3�'ˠt��4�Q�숐iR�B�B�ϝn�t� n'D�P*�'�Sa0���L/�p�P�o"D�ԃ����.�|d�A F2>r���-%D�`�#Ǌ\��H��ѥ|7�$+��#D�h�K �R�Y�T1�����?D�H�!( n~�T捊�F��q��<v �f8���0`۲^�vU���V�F�F$	�<D��:#�V�H���2 �v��e� �=D�(��Z�vM\L���״N)���7D�<��`@�]�4�p�.TN�pI�7D���FԊ9˴T�PF�jZtTSQ�4�O�����O���CA�����07<��4"O�A��/�ļ�!G��g5>���"O��!�5A�Ņ-Hm�`"O `{��>[~q�O�N9^1d"O��fE��$�.��I���g"O޴�U.>&��Eq �Q#y�yH2�	/HR��~�f�|��{1%�_�ܠP3�V�<�W�ׯNt����j�?9�)���!�^������![��f�<!�d��*�R��WJ���FR/�!�d�q���G��>�!��b�h�!�dFQv��cm^�=V�i%��)}��X��O?E���JX��J��Zy���G �i�<�%�N*S!$�;���CXn���G]�<�c=j��\ �E�=�4�a��S�<��fF�� |���Rxx�Y���S�<i�L�1���z9��[2kډ��B�I�q>���jL�2��u���A�Z��"T�,�a̸[��u�7�� x8tQ��d��Iعq�D���?<\������u,��e���T��-�	< 6�������S�ezg�-U�Y����=f�,ɀ�ŕ��؝���)5
�4��$b&����2L�p�k���a���8��ŀ)<c��P#<͆@ʥ���{���y2��2��5��l9h�O�9���'���i�6J ���j˿y�R�HCb����j���X �E�&m�����N�,<"#��4��/��|r�S�kvj�b�b)S�N7z�`�Qn�<�k�!�?i���?.��9���O��dP�x�&L�4m���̱TԹ<���d��d��A[���������O`1���y�c��`��Q�L�>IHP>O�Ы��U/ѓϟ0�"��̦XfF5 �B�-��˧%��2O��%�ܸ�K]�#��)�)�D�I�����'���حg�j	��@5%>�g��f�!��_�e��Z!)$p����Dƣ��O���E@����M�!.8��#Ao,1'� lf���O����58]�A����OZ���O�$�d��H%"��T����#F1n0^D�G���dq&Ҥ
Bj��G)��r���H��"���C�<=��m@#�'��q�¨2&�I��[>SǂE9E�4X��c�	���ϦvР ț�B�r���&?y ���,�I@�'�Kv�X4
�@1Tup�
��>���Ս�f�rT��%��B�R�ņ��IQ����'V��$�z��k�'r�$`R�M2�Fl3sL�:��Iʟ����d��͟��	�|���,F�v`�௄
U��	`C�jj�AG /<��<Y�.��?����;�.�j�;?C|���*�2���e*�D����$�N���䁱`�0 0G˟3&��O>,0G�'Ʊʲ�	�i{TY��-O�-�0�K��'Jў$E|҄@
Vb4�+QK_{h�(���'��<i��D�$a���y�'R�����@3��	 �M�����"k ��O��>�@d	7j����e�5·w�b�z6�'?�	��'��'��بd�� �L�·I�g��T�ωϺ+#mؿ�P]Q˃ V͐��р�K�'5zݲ��" a�,�R]؀1��ְE���I$�N� ���^���^5H$( )k�'�X5P��?���T�[�/e����ϛ}>��;�Ŋ����7�O  	C�Cld��ʳ �����|r�i>�3)OlX����T��Р�Z�b�q�_��k�-��H�	🨕O���'��Bâ|Fm8̊�V�.8�sŗ�\�"`�)�rpkT.��"����菺Jk���'ŘOl� �?rq`d���1)��Ai�'@!j��K��.	:!)�r	�I�'?H�ܑ�mX���"1P�E!λz� �;`�I�!En��X����O��S��S~
� Rᑆs�֜�7N�Ek�łv"O\	�#d�;|L���U�Sb:t���D�ODEz�OC�]sV�R�u�偀�	9H�3C�'5r�'��M�G�10�R�'f��'��T�'�]�e 
^\���4V
8����.LNjT�ry����c�+y������'�����:	�����&���1V�T�Ԙ�S��|xUQ(An��ӮGR�T��gD�>4f�)L����5)`�ȱj�H�"�i7RL�I��D{r0O�]�Wn"}��`ij̮9[,11 O�A�g�I�.�bFM�N���d�O`�Fz�O��Y���fJȗ9����䃘���i��Քt	U��۟(��Ɵ���?�����ͧ8c���	Kr��3A]E�d�Sx1��cP��Ex��\v1����2BB�/�<�1g!�6az<p'G2Z.LA�2b�Y9es%���'����BZM�<0��m�M��D�Fzak!o#z���a"U@4��$%ړ��O4�	Q�"�I��a��"4&#�'��h���\�H����R��è<�ԶiBS��ʤH%�Mc��?1�O�4@R3A��n8��2�	�� Qp���K�����?	������똧���R�F�م%^��0�䄷��O.M �S* b�S �� ����BI�~z�">1�͟`���T��1@ȡ	��C�^L�
2\��y���{/:�@ ,f_PEj������!�S�$��<��B[y�����Z	m�fR�#�|y2�'/��'���'��`�D��?���9��ȔH&j3`G���DK<\�1O��Fz��>�l%`��`�|�I���,E��O�x�U�x�j��l�OV�%��d�#f���`��h(�%Lq� �$����I�e�z�d�OH���Ov牣%Q�x��L�'�D�҅J��(�*�xG��Ӧ9�ɛ^�p��I�<9��fnz�I��ON�I�U�R �!猃eԾ��P?�����?!Fm��y�� ���O�)�OH���*ql�)󪄲U��h+H��`�9��O�$�6 �J���ܟ�J�?7���y��v'��z���~�RՁ3jݪ02⚫�?���?�؝2�'&��O6�D���)݉4�B�k�c	1��<C��#H�-�ɻ?h�d�Oj8�T��OJ��I� ��s�- �!�;V����Q���36��t�@���Am��<�����,�I9(���?����g��-�d̈ j�,g�]���B1]'� ��'�@Ɋ��?�w����b�+D���?Alڗk�DB6aܞ]���i`$H*L��'�M���'�	���?����=�����8��7e���TMދ&L(���E�=����4D��eX�'�(��6�i�7���H�ĉ��0��U�?a��˙�*��� �c��=�)Tܦ����M+�U�("�'�M[P�O]�韜]%&(Zhx�:7�8�2K��"��B�I�E$��ȁ&,��E,�2�H7M�O6��?���?)���?����?�#�#i?`x���0K�e���\��6�'K�[��'��'�B�'�~d����5q����_��R�́nџ������������'�2�A�7c��z��ܮ��js��.F
7��O����On���O`�D�<����~2b�9��H�ǈ�~��pB1*�'��d3<O"�b:�@��դ'�19��C.[v��G��ɟ��'���'k2��5���03$D�AZ4�DX���>-O*��?�-O��'f��C�� _G����C�.U�8Y�	�'Y`�����R�h�e�DX�Is	�'�=�d�~��I������	�'>x8��[�:5�e�y��U�	�'�\P��T�>%��"�GB�o�TyB	�'�|��V�0`�$1s�i��`��:��D�O����Ol�D�O�x�pe:Q��uP���_!��:�"�Ϧ5�I��ş������	�,�I��Cg���v���7h��1��LA-�M+���?��?q���?���?1��?q�N&���f��V��|�f�T�W(���'��'I2�'���'UR�'�Rj@�+�F`�'�H*�ԙ�PM��6��O�$�O��D�O>���Or���O
��ӈ�H@�Q�Gl�8{&d 1@Qm�ޟT�Iܟ���蟀�Iß��I���I/(e&9z���ЂO��J� E�޴�?I���?���?���?Q���?i�FG��j�j2y��6��?#�ڑ�s�i�2�'r�'~�'H��'��'�X��fh�-+�+�u)�4��y�$���Ox���O���OP���O����O:̛�ْ2��t�@1m"B����ۦi����@��⟔��ןH��͟�	џ�[bbX�KA��c����ҩ��MC���?���?����?����?y���?�v	�VH�a��$4��iV"���'���'���'u��'���'��Isl�=�P-S�+C"|)�gL� ��7��O����O����Ol���OD���Ov�$� d��ᅶ M�t���P��o�<���?����~*���(� �@j���#���M��OY~R�'�_>�ɞ�M��wE^��EV�����Aۆ]��M�G�'���;O:�S�3w��0b4���V�Ӝ7R�����յ�	����O��U.�\M��n:�	���<�Ѣ�Bxh�XR�!RʉC�`�'z�7-�C����\� �D'M����yP7&��q z����'��	ܟ��)O&�${���INyr��,0d��ʟHJM��-��$��Cx(��!�7]P�i>a�㜐m��dϓ2dV͘ �\����I�N� hE{��'T][�DЧ�rdy����ъ�C�F�î�y�'��7��Oj��|��'G!4Q[W�T����hGm��a(�j�'t�i��n��U�Jh��O�Q��
II�R�H]w��H�ģ�is�\
�%�9��,2�B�'�r퉥6ᠨj7�ϲ&u4m UE�:�0��'�:6�אk������F���'��z�&R)9�V*SA>Eb!C�<Q���M��' �>��!/�-��$Q6.9C�mJ�5�R=�2�;?��&�2m��k��7���?Y���RL`��	8:b>h��
	
�r��(O~�$�O��0& K����'<�7�4����L7e��[���@����`��ۆ�����1&�@�����ĕŦ-�ش$���";��$�C%�O��xcC^�<��4)H�<��i1�Lk�̟79��$�(O��)����ÈZ<���F�i�|�� ��?����?����?���?�����O @a���Q�>�ۤ���c`�����/�?��U��v.�	�y��'�7�7��I\"l)�����h ��џeI�	R}B�f�"$mZ�?M�� �i=X�˟�����3O�1�F�9(��dkU�D?�\"�g��^ &�X�	0��ퟴ���� ��(���(r�O��$� zU�P�p�IpyR��*��t<O����O(�]�2�'MҌWʁ�a���(U�Iڟ�P�Of�m��M��i+P�p�I>[c 	bA�4H.x�I��=����D
&/2L���<�'O:���p���$�O>���f�-H
:�(��I)3��B#�O\��O����Oz�S�7�:�lBy�An���ʱ�ń,ö qO�O��v�*���Of�l������d	�>1Źi��	@GV�U�eI�˽A�T���/|�N�nZ�{OX��r�q��	�Xe
	���K�-���'m!�CP*-T!"�͏!�$�8b�'%��'�R�'�2�'c��'����:��96����lM`��˻L��Io"���I���|��Lqߴ�yD�v:V��(*R�<�y�j�!v�Ƅa�!nZ)��d���������$ƫu|���h����X7Y8)��#�Mi��$ӫy6�C���#e=N�O��OF���O���gٯF���8&&��!�Q��O�$�O���<A��i�j@#�'���'�Πc��%FU�� �7r��U��|2�'���m�Vk��poZ���K�p}1���6�h\֠²���'�X�bL]�^s*�Q_���d��ŉ�,��4�r-N7VV�iI��_�:���D̙�0�	ߟ��	ҟ$'?iQd".6;bpΓ���t���P��] �Q�Z>	�I�M����<���?	�L�O����ܺ+�OX��1*�PN��ЖПA�D��9Op5 ��'b7��v�(�X�3O���à%|0�9�n�i4ڕ��lA�u-��c�	��8��X��)�$�O����O���O6��O��S�B���iB�Kxx{�GG���a�F���y"�'=r���'����@F��V��-O;;�ḍ�D�>aӹiy�6�Z̟ '>��S�?u3�ߜf�uA�#�!M�+��,y*��𢙲@7�ɨ�Ժ��H�d�q%����ʟt��+W|���S�GKcS�]�0n�џ �	러�	�r85�ڴ��ā���@�L�?4���Ҕ-�
;�pr�P��|�4���?!`R�,��4��u�Bk�$ (�L�W��?�����G� p0�b��<q�'�8=!A��1,�L�,O��	��3 @�>"�1+�`:	���@�?����?A��?!���?q��	ӽn��P�V��d�0�񂧞�S�Iڟ�B�4$�2�̓�?���i��'�08х�G8��"0 &�Ae�O(�D/�&�t��iT�!��a�%1O@�w�*�hJ��U����#͚i�����܄M� ��P�<)���?1���?���?q��'.�(C7��7v�v�ia���y�W�P"�fZ��(�4$/�0���?�������P�f|�1O� H~�A񆋪qР���?�T�1ߴǛ�O�� �I�[3�t�&n�T	<�0�N,1�!��a�0?��@�T��<A��;���
B!U���;��L`��O�	�|X�����'[�m����?���?A���dH��|�+O*in�H#vd8��_#w��Q�g����D�g�x�I��M�O>�'7
�I9�M�Ս�	;���Q��.�k����Fbr�69`��k��d�O�L�w�])A�X 7�<y�}�1�Q��!8ei��w�H@3i�/��uHr�Әj��U�.��?�>��ҹ<wd@�iA�?v��	"�U�<IDM #k�D��ᄛh��Ѵ�\�x�,`R��Z�I��oW��i�O)� q`��t�~Q�5�Y�l�|�2�	Sz\�(����E,/	�B�p�$Ē4�j��@��C�J!rq�@e*���C���|���;�e$�HM0�Pb�0��x�'���xrh��8+�m@Wd�1|��kbEƜ�x�O9�,Q[f-CLq��ڜC�ZM �H�uN`p�F�g���+��|��e1{<��v�ߖW�
�@`M�'�ƭs��؏n�nkD)����wO�*h+�PcӼlua�`�	�e���w �ծG�Ĉ�<�L�b���@��#�K�@r���/Լq��&�'2�'_vQ뷡7��O|�da�̨��B5���[�@L�^k��bRK�O ���O���J�Z���'�?����?�������J >�`@�Ú$e�9���?�
�H;�'q�'��'p�;�b�0q"�H2q��c��ݛ��'�83��'>�']��'���'���wˈ�+x�93����0� vO�O6�D�O��O4�d�O�XE���elF��gj���@���,0.���Ob���O���Oj�D�O�E
���?%���m6u���R&5n�aZ�<���?�O>��?Q�KӒ�?Y� ���O?I��i	���Q��9��'��iB��a��=_2�q��X<x�b5[�D[�ൣ����Q굈�����h�2�6G:ج���OX�d�O���O�Isf��y����O���e>��_:dTR�ۦ��[L��+�O��O��OX�$4��p���3�u�^��QG�/1���v��Ol�D���oZ��?Y��?��'��'J���1&�K�	�	���'B%h��EF�3��Kt���^��Xm8��F%1C"( ��ſ(�U�A

n��ӭ� Pu��J�R�h�e
�sc��c����pN����z�|�k�//۔!��#�0w�D]o�avЅ���`f�yΔ,c�쩸���SD�Y���D�q��'M��u4��#���Y��R4�@D����"'DsT���"ұl��$�oP�xLj!�t��01M��Mi�^�+�'-P{����I4w���yV"Tt#��*���!@�~��d��]S�E��eB6LtP����O�@�d�O��DeӜ��T)�i�iH+dThAg�ך\��{���;�L4ZtK
ou��1��n?цB�_�H���J��E�Wh�TG�Q C��1�p��B��C���Q�e@"_X��")�|BQ7�,�5fѭ�\)U�9z�L�(7M�\�ٴ;��8��S�?�'��O��|�^�K�6 �̕@)8D�̋P��+@Y�q���Pj�T(s�1}r�'^*#=	��idR�ib���Qn>3�Hqa>,�ny �O��a3k����Oz�d�O����?����A�l_�[7*Q���ii)T���vc=wK�H�2�֌��ם#ʈO��'҇["< 0��lެ��3��=Ue=�����&�1��؅~{jԈ��$Knr�'\�Bb�<}@p��I�d�@��޴[L�p��rX���e��34��J�s�IҀ�#�O$�{��U8C�H�6R��T&�18�Dy�o|�8�O` yw���mnڕeO�y@E���+�4};F�ĭA��\y��?9��ysL�z��?�O������D�p��h�T6�&ia�
G��j����������b�L ņYJW,�K�c��sR�����W`�]
ª_y؞��O�$bӸ̳I�zE.���b*2%ڃ�>���?ٌJ~�@��*3��yw�^V�A��k�m�<q�lJ&Scθc�A�����k�a�)W1X7M�OLʓ"'tQzѺih��'��S�2f�}��@�_�� ���+j��:�����	��$뜱C��Azf���f� 8��S�T��H�Ϗc�БF���'����3F�q $�6 Vj}0ԦK4��s��`�`ź��ڗ���T�)o�P$��\z1O�Pd�'o��~��\6k,�#�`ԹV�j	�Rg�g�<���6�Д�vEZ4GB��Ă�l���j�{b�O�o��*��� ��EÒh$����C릹��ʟ��i>�+���˟��ޟ�m
�T�
5o��Di��ɧb�j:h2�\�`��ٗ�FJE�7��V���Oj� �Y+��8$��N�H�)ˉ�P���S�.��i�#}�'����EF�lv��xU�&d����J�O�L%��ɏ�Y�L���K�Q�� ��64*xa�(8D�)`���l����1v��[5�Ʉ�HO�O$��HD�?>϶鰥�	we�LjD"�O��ɵ,��$_���Or��O����6��OǨ�6Qv�
ek[i\���l�"�M��Lx؟�#�B��X�^ъ2!@%}�I���l��4�V�'L`��͏��L�r��%C.�Z�4w���I��p>�!G�*>Jν˃cYY�����y�<���G��8�EnG.y�:A�Щ�u�'b�c�XZ�J��M�4J�v�
��}��Ӗ�͆� ����'�B�'�L����'�R>�.M��1.���TL5/^ȴ�6��*x�<K��_�*!J(�c <Of�*�߯��re� i�at�E;�I�u��5��E�傏�t��dj�$a�^�{�˒��?��O�����Aj��r�'ّ]�~��"O�u�2"��hQB@t�4@��,1&"O@Y��GHN���QHT}�	DT��M�I>���R�;��'#�R>UR(B��$`r!�tt$2�ȅ�RK(���� �I� �x+U��=ꨜ�R�Dt�dB�ޟ��]�P��vfp%0 GF��H��}2`�����+A(z�e(w�l�T�s�@�~%FȐ�mS�ys ���v<8�z�(C�y�ГO6�z�8Oң~:6$�6��e�+dz�����z�<q#��%�t���]�D��lJ��v�� ��{:��׃|�2I�D*�O/6�j����
�$E��4�?a���?ͧy0p���?����M�B�ЩR�`��C.˥k�ZQ V�P�M+ՍK":�p��L�O�i�'ܘ���ԟP�X+�%©Ar�H��eJ*1��mh@�J�!{�<3'��=z*l��T?P�"�B,�T�}޹�b��p�@Ǐʜ-�l"׋�;�?��y�6�g})�p�n����ЯO��@Gj�/�y�F�7+�X� ��(p "�@Ԡ�'�"=ͧ���ӝT3���6��h�.�g(3Zo:u��c��)ʐC���ş<���u��'��;a��r���	u�^�# ���^p%H�)A(!1�Q%�1�Nغc�	�0��x�J���9R@��l�#���'�*l���س>'ΰi��jݡ۰dE�>~����U�DȀKL�T�'nq����C�$�X��4HH�D���p>� ��i2/�NTٲ��>��9�5�'F�	�d=B9�w��6~�ǌĝzw��<Q��i��'L�B!qӄ7�%G���!���l56�xuOZ�qC�Q��ʟh��13�i����,�'OZ���f}�iY�,8���NK~�&]�ΈŰ=Q3��}�f�-�V�7s�%(W�!j��DW�����l 1$�N�|I�@ћd�VxG�-D���p��2N��	���:&�>���a D�4j$�95}�l��̛	��A�`�^#9=�OJ�qg�Ϧ��I����O��A�"Z�%�����H�TǲI�D'�3,"B�'+r�S/x⽃`��%�t`�U�O��Ⱥ��@�\ F�ĥ}�4�F`�r��p�d��,)��s��9(��tɐ��x��i��ʀ"�r�{�B��P8��A$ L��ɠ�OE�m�(`��)� ��+9���*e��y�
����B�)=dp��"���p=i���Os���8��]J,��!�R��TA���M���?���|b�F�:�?���?I�4/(��ǉS�P����4P���'�1O���g�'I�I��J-M��Bs-�	KR��KV�3�^��>�	�0Y����Ҝ�U/��TV -�0�'T�O.=F��O��b` �(��h�D҈��lI�"O�=Ɇ�:dMY�:3|����Bf���DX��0�]_�����î�Ҝ2i١�?�w"��+�������?����?Y��f���O�����(2㔂Y8�����M��F؟C4i�0o��h��A�yK��ڀ�tӨ�s��'>��1�
�&�i��ኌ� =��4>"Zq��'�p>��]��[VEٷ�I"fMy�<)6i��&<e��D��&�b,�c�	-�M�L>䃟U����i�
0��r&�z�B!GYX�RB	�O��d�O�1����O���f>��OL�l�@L��nц2|����<b�0��I� ��O�Pp,P9@�B���A)>y(I�s�'?8h��zr�D �O�\��O$�b)H�*!�$��)[��YaȄa�T� ��yl!�)4m��B��ĩ
%"DU�^S�pm��4��	�+b�i�B�'1��%a�2�����C ��'\7UqbD��S꟠���4�'J�hN�%�ěx*�Pם�C�4ap�U4�$	3�i��tb� /�3��ɉ�IX�2,`!9��]7M�z�Z���IW�O�,��'��6��K��w��%0@�, �E�5L|H�l�)]��`�)�gy2�+�"	2a-2��ի2�0�p=12�dH�J�&UP���?���B5nH5J��cA���M���?���|��O�?����?IݴU��uK��)^��Y�3�8]��P�-R?SZ�أ6�ӏ���U���OV���B(P��S��7�~�RB��M���� ԥ%��Γ Q�>�O$!)�H��ResFiG+@W.�$�']�7m�O"��K���Sџx��Ɵ�mZ�1H*L@Ġێ&��E��n7C���y��Ұ?�ܡ<vn9BIFn�2��O�ss��dX�4�?a�4�R8+�AP)�x��F�?���q�'��e��Q8m��'���'�ٟ֝����ƘJ0�
c�UC��ڔ>�!���iN�%b
��{T�:��O�R�a��Z?���nZd���dϹd��L�pg,��`p�Z�GM����?�
�[Hd��o�=$c�x2��q�ȓ�8�v�@�)G�l2��A���Ey�a��O�TJ�ăælڻ"�J���n��2�����C���?i�=$����?��O��Q� ���9���:-�X�ti��$7T��` �XmȈ�#K
RfH�У�g�'z��3c�o��9᥆�����ʊ~.��6��F��Pb-��
�p�dt�'�@��!��ć;Rf�U�f
�9j��"
1!���C۲uH��ز-j��*�/D*�!�7-�z���B	�)R uՅ
��(ݴ������A�ii��'0��76BT}1�#��y�2��g����eiw�՟�	��H�hS�vI� ��U�O�r	�ĥ9 �,� �$Xպ��)��R5�(h4�HO>6eB�,�^�X`Ƃ�Gj��`�U�r��гJ�	1g�tB�c�?g�>�Z���2�dX1K�+�P㞰����O�<G�D�P8Qv�x12g��TI��X��yl��'��|�E
�0	R&�b4�5�p=���$ACO��W�N�V����트x+�CUDE6�M[���?���|�aC��?I��?�۴fP̰���ۥ8�EZ�.�2<��E�'�1O,�g�'�8���gy�e	��X���C�*\��P\�P"v�4U��>��^�zs���4�&�t�.��A�'���O �G��O` �u,8Ru(m`Q Ƥu� ��c"O� N�)���/,D�S Y�nM��>	��aM���D}��F�}��� E�r�&���;R���]hX��@��OF���O���Rպ���?�"�|�w���S��S���]  U@1�,B8Ό�VG�R�,���݅E}�I�w�R������|
�Q�m�<��,�nE"��Z�#רo�M�\wy��E�:��eCJ>R�O�L�l���'ð��Q3�e S�����'%66���}�IUy��'��'mt�p�CAL���ee� p���b�'�N�3��PW4�(���kd�Z��ڐQ�L�$�<!s(�iB�u�:<a7��/lrxM�靯g���צߟ�����Q���ޟ����|��o�	u��T����CF�Zu�K�1���z��,+�H "f��bvR�c M0s�L�<	�H�5+��!!$͡W�4B����BƘ#�D�plj��:s��Q��٬'H��'
���#H���~�B�*�ĉ��oņ����� �y"�� P�#5�J-�$�rk�	��Oz#:3F�~߶Q G�M:=9� ��3�*6�;��ڂ$Ql���	N��۶>�I�e�4s�F�c��`�|�P�'Vr�'�.�h���*[�y3�/c�(jI�~�Yw��򩖌�,)p� TT��}��'ռ�1.N6`^¬ڶ�
��)Xrr�����
���B�7ٸ`/�N�qObL���'���~����7 ����Dc���tcWe�<Ʌ.\� �t�4I�0�hH�5�Q^�����{��*�З�М8X�逪E�7�-:�N���9�I��X�i>�qV��㟘�Iӟ�n��<h����w>N�U��	#�f� A��(Y�y�$�y*�I9�?��|�'z~m�'�¥.�"��l�  �t8�aa۶N����#�O2v�f��1lK9,z�m�t����4�O���ݧJ�,pȢ�����M)Ț�)�O�m%�+��Y����]�P1\�H���{�
��=D���Rn��<!@�jZ8�Q9�b!�I �HO�ɨ>1G�f��!\���gF�4Y)
�2��'��D��Dg�'42�'���۟������F@�!����ۿ!���1��Jh��Pq�7HiJa,ԗ/��N�7I��C���ܦ/���ߥ8���2�m��^���B��Aa&*!�I�Y�,��^w�`�݃I�,q�>�Q�ݪ\��;���L��i��KI���{���Oxu��H88UC�AR6� Rב�����>i���p�*|C�_�Cxl�20G�[�'�
7-;��ĔN$n������g�Qz�u�!�:c�����L;�?���?�����?����T,!�?��O�D���ТVĸ1y4�Io�<;1�'����J<���[�]��3��M�)g��Vd؞�i4e�O��S5���Q��/4��Lq�¿y����ȓ����5
Ƃ���%��y숆ȓ҄(��I�d&H6*����r�8�O�� ����Y��ԟ(�O�xs���u'�PZ7��}Z�Őa�S�1��'S��/"8EZ�e� _BZ�[6`��G+h�'�u倃�x-�6�;-R%a����'��@�L4h\��� '�
dAV�~��ƨj���� b�F�,)���@�HBt�	���6!�u(%@���	�̎���,q"O������������c�^���'_���kv�. \��B�*%o�B���<F��ҵiT��''�O�*R�'@��'ݛ�bݦd�.HH�G�2PA�������2Dm:,�d=��bf@4l�x|R�O1���I�0�ЭsG(��,�4��BG�r`.�)��в@�B�ca�^��U)W_�	��a�TnNw�����'��k�L��GBY#+.}��
�}�Ҋ4��D���đ�%���X���&:�0�H��"O6�Ɛ�)��t#R)B(᠌�&���t���$Z��`"��m�科��������?�/լ	�����?����?y���n���ODC�C�dˤ��9%�
�)P�� ]�5��ibf�9��#}��G}O�*n�)���!W�8�NȦH�d}�" _�\���� 憸]���_w훶HQ.G���H>iQ�Ö(X�j�M�"�Ԏ[��i�Ҁ�O\���ID] j�U�+Ԅ\�F	!:��C��q[��#��<Z�J�̆-Z�<Y&�i��'����Pmz��7m#~�2�P��D�~���Sa.F���Ɵ�I�qH\�	���']��%��p��D�(=��x�J�%c�ư�P�?�a{��$��� �8<z�ˣ�	�1q�Th��0��9B��.D�1 F?�A\���+�~�eƐ�|�b�GS��F�*�J��y��܎z�쌊�)��[L��y���L��S ���Z��W'a_��n~�	�z��$�4�?a���i3g�a� ̀;'��|Kg�Y�f�"��O���O �����B6��a(� ���:tBW�D���@Y���-�,���mX.�C.�O^�f�)?Z�� I.[����Ks݁��" 	U�:y"���E�6�����z�8�&�=�<jX��Uq�OPԬH�A�*�'`�8��'3�l�W��<u+���f�E*v9X��qO� 0����� �'��k�f�P���)-����4�?����?�'D�X�Y���?Y��Mcr
��+ggvr*�yPl����R�Q.�a��7�LU����O��K���c��>�t�H�%�$����L�0����I�t2P��	��r�e�,�� s�����._�p�	�g.qcR������?��|�h;�g}B�uy�#�jjv9���&�yB	>^a�BE���H�ZSC���'۲"=ͧ��d	vt�02N�%@'VP�bEl��k�ş\X0N$�\T�I⟐���� 
\w�2�������;<�@��G� _�-� �.�"�؀E��y���G�9}MbT���O��9n\�D����>s�v�	�$�i�=�C)�(M[�8R�m�`!�t��(�$�ھ1�';:UC�a5�^� Klu`� fӤ����'g����]��Ƶ�kQ�_ 0�k2C��?A!�䀗:b����i�ĥ���C�Q���۴��K��1Y��iU���ô�6`�֎��y�6��:����O@�d�V^���O��'ߎ\Qb'��*���*boK-7�
�I6��v� ��S#@)9�,P �PG�'Q��W�B7ä@����u�����	e��і�ߘ11��0&�#N���3�P=��{�?1�O���π������?d��Ʌ"O$ q���,{,�- �JɭB�6���"O����L�����lܖ%xJ%�ǎO��M�O>!�B]�	���'�BQ>�c6��!5��D��0�
��Y�F1��֟X�	�DՀ�k�8��`7Ԗ ��Qr����9n��f�\�JX��$��OG�b�<pchߑ C�|�p�M�cT�a[rG�κkG�!X�� �f̺Q@��ɤ`�d��Q�w��U�]�(��I���� U�C�����)�FA��z�1�"O�es�oH1������H�6��'ψ�����E<���U�(H�t��ΆIW҅��i��'��Ow��!��'["�'��H_����,�X��i1��KQ����20�����D{� i�OC1�t�	oFZZӁӅj��S�(�i즁�ed){xEab�R�S�����V5Z����Y�i��р�,Vt@�c"e��Q��B�(����'�B�O&�F��O:e
��Û�X C�U�=5��0�"O&)�p�
� b�)�!�!Kl�H��$OZ����R��@�o�d���[���V) "fN�?q�$�i���?A��?�ս�L���O��������4f���0GJ�/�4��.)�$�bG,ED:��ZwQ���m>-BG�0�����^='�0�q�\'R�3s*�"VV��z���87����&�|��ϖ.� �Г)ɥm��m��@-�M㒥� ����mؤ_9 J�%d�\����ȓy4�qt�Bp��Q�f
�y}EFy"Hn��O8=�$��ܦ�m�S������cĔ�1�ߗwo^�����?��m�h!���?I�O�JL�u��E	�q�̜q��q�N_�Az�S���8\AMq�OV�`�џ��ȉ�Dî�0Ua[$o4����,&bx����3^Њ�D� �[��o�f@6�r�l4��2"^��^?� �~(��V`�*k"�w�<�V�L/KmJٻ� "$KG?s�B�	98/@���A]+$U��T#W�{�i��'�m�)z�,���O˧9�4��%��_��4��l�$�<�h0���?���?��(^�4�����G�1x�"��J����պ�U�L6|)S��H~���D�S�|_��[4 >(�1�@l���u��
-'�U��#�' ��F�R[Z��'�O�.$9J>�g�O0��ɘ�D��!�ˌoN����A��!��^U���!��h��Ih���D���-��|�����fԱ��J,'����d�P����kŚ��d�O��4���c ��O|��O�6��_|��)v�
6���$n\������ SKPp�B�נv�.�C��.k&��|:<��\r�#��_��5���	<�В$���Hj�c�O�??��	�%@�_���;P�7���y�J�~7�!8�	�GhI�G�%Q�V�$�¦���4�?)vi4�g}�D������݌;R��R@X+LA��&�O��+�ϙl=�8#� ��<���y�'��'��F�x���@�K.@�!*�"�;����E�l�~�IW��O����Oz�d�s��?���V��#�+-Jh ��DL2r��RH�	Q�����&x .�
D�mݩ#���s��O�� v+�;��2`@�-�j�yaWt��1���P10&�i��o�� ����v��I�2�I�[���i�`�'����/�M5k�ҟ���<��]@R�O�]���a��!pO^i�ȓz�0-��Q�\��ѹ�E���,Gy�v�j�O�p0�]��nZB.�)!��;��,�C���p`����?��@͔|Q���?A�O�8� ��Bs ��f��/n/r	Pd��3{�l�Ab�Ǡ&��lse��ESĸT-�D�'�l�aa��(��|Z�#�&Kޑ�b��p=�%K���lF���!bS7@JJ�D��i�'SD�j�'G��|��e[���<�U�g�dj	�'=�Y1e�3w�KI�}�k�'���W��d��h�d�܆B�b�#f�QЦ�&�cP��$�M;��?I-�� B� ���vj@�+����dH�"xvf%��Z�����ğh���[}�m�u�
���G��>���~�рƊ��,r�0��ϩ`?�ęb�=�	n�D�2J�lй����@M���)aAiP�!b���ԉF�0t`0�DQ8��%���h�Şc!�-�U��3�v���u�<���AN�`Ͱ��n�0,B2�뉌Ӹ'�@E�!o�F�l {!�-a�zxy�遜r�
4oϟ|��ޟ�ӹr������t�	즭��P2m$p��DUN���s���w�	�#TJVx������䞳V�v���#/�X�n�6�j勚�8J"����G.	��5��S���Oy���x�Zp�t���XG�љ6�����]����'��#}�'�d S!�ӂ�9h��;�c��yr�1M�bLH��])2�"a����'nN"=ͧ���� ,1�L��.��.t9`�*���I�8UB�A��џ,��؟t�	5�u��'��;B�� ��Ўkn��a�Y��1�'/��P��m`��R,��Ql+�&�F}��_-2���Z�+q5�4��T_. AC 4]� m+b�Z�}3�H^�M;"���i�PŸ@J$}�g@�vl�Vj(�D��&�_xL�`�ON�n���M����?���?!��?�4P�nJ� ި�$�#��E�n�А���hO�>��	�����Վ�4���Q�>,����|bc�����<�0H�>ۛ�i����1� A$�;Fc�"
 $��s��O��D�O�	YW"�O��De>�B�e��C�(��MG�+�BY۠CI7I��p��B�o��u3�Y�Ox���/G�V�Q���lN�Y�P��O�;kD
<)��Ա�H r�q �W~��"��q^Lr�;�I�S��d�>�6�T!B����E�H�y�.h�<厚�^����W vb�yy�[I�<ц�A�^S�-�b5k�(�Ӌ-m��7M*����>�2�o֟��	U��g�� |����
o�xp��݌U+�x"p�'�"�'Rq9����"�7m�#�����|�[w��|`��Z��E��8a�}��}B�U�D_Q�q'@��kD�[9	�`e�Ģ5~<���]�4��ة��	9�00��W�_���ܨ������},"�NE��iD"O�q;�N[8z��hЂNX@iX��O��=ͧr�qO�E��b��x}�xb��P4�G�������/�M����?���|�CP��?����?	�4CRFm��iJ��:]@kN�|  Sg�'�1O���g�'���3��	E�Qk�A����86D��>� O �	s��#_��yI�#�s8i��'1O6yG��Ov�;b�ߤ!�ȬQ��6u
����"O,���V�_<��#T %�rM���Ym���$Q�h'['����`��t���[�)���?�0�������?���?y������O�� ���(A�f�q��Ä�Z�9�P�!|�`�KݞZ[L(�^w!�TJѠ]�s"��A�Ȇ�z5P�js�V3/X��2������.����e�����9
 ��Sdf�P�T��6�U?y��+��s��D;��'���|��'���xr�վ_z d3j�>�$�g�U:�y���-Av=� NL�u��6J[��(Oo�� �'���3�cx�*7M�>h�5!b%O�V����b�V�de�	۟�	9�\|����0�'u�:�����d��MӃI�-H|`g��s��t����Uq�'<O@=:��*dp�K�(��[�b��`ו|MeS�*N�y�*�V&?2p����^�,� ��{"�[��?9v�O�iPt,�i��%Ӧ
w���@"O� �i̷,���	��f����B"O�u��^j� `�7O�<bdVm�f��MCJ>9�n�'>m�&�'2[>y*���F	1���X�l���ڢ�t��	ҟX��O?v��H�;�R	�o��|���x��L	�d���ےg��BE�H�O�c��Z�͓UT콩��;Yk� Ѐ,����؁vh��ҥ�yz� 䊔|`�P�JVQܓ=4v��	����n��n�	ǐ�gj�<�q�"On�agԎL�|P��o���'<�㞠 �O�>oJ\�X�9&]�\����G:�i��i���'��O꘸Jq�'A"�'Л&���=ԕ%�76������߽랬��U�j�N�*`i0b �-/fP�i����ܼ��,Rs�,Yd]+&��ԁĭ,��U1�I�A5"q�Àz��p����uC�����׼[��M�fĝ5�1��#E���E�r�'���'��}F��Od$�4�B��:�jVL���P2K���	�A>A�wF^�&����� �>�'Er�4��
���M��lՎ,Ԉ4��8I���Ѧ$Z��yQHp�d�'5��'�Ҫ}ݵ��ϟ�.M�
Z&�Hu�\m���z�oL��&����?�1����m ��͹bs�!K�˦�zvE?�O:ph�m�/
TJ��2n΋f���X��iʾm��1^�|2Ó�w������ �f�^������y��C5>�r���Z֔�kv����(O���>ѓ�D�b0�f�i]�ٖi
Ljn�GW(�X���E�OP���O�@{%��O`�y>���`�h���H�ۀ ������	D�uLN�@&��(,K�R�����*�^����W�����P�(Rj� 4�K�7�!)��C��݃!�hӢ�(�!�8�qOT����'6>�I-j��	bfŝs��١$��/�.C�)/y��%*;'�=b��QKC��6MN� B�B9��.^�m�Di[��M+J>�q!P�=��I����Oy���W���^�B| aM��cf6)����,��'�rY
<�j�����z���i���4Pv�⺳�g^m�����&\	T"�HRk�!�T�����
/�%��F����is��"p��1� C� |ؖo�/XhA�r�&Z�|1j�O�DЦ���Eⓨ/PŊT��;���aU�`9�����?a���d�O��?���Z��@�֊&8�K��6\�B��'�87M��1�	��(��Ǒ�j�)��ƷM44m�m�t����g��L�Iǟ4�Sz���I���Iצ���- VN�@+Ӯ�=[�����.�T��#4 �|�'���Sk�g}b�L�r4,�!��&L|e����)Z��4��;��(@�$��2zH�Cr傖rG�e���~��3�E�a�?+��M+WK! �X՟P�J>���>QE"ɿ[n4�ÎT�wh	��Z�<Ʉ	'/d��ۤmՈ�XѨ�DKܓ%S���S\} ��0��m���L�"��H2���~rM�5gd��DyR�'��	ȦQU���!6�8��B<`�r-#�$=�S�'\����珤G�(�˖�E)JNE1�����?q��,��e�$��-�p8�"�O�<9'�<b�,�cU���:����E�<ဧ*Nj��g ʤNL��@Ԩ�^�<ْ��	.��bK�����)�G�<�\}�����]���kWa�J�<���0f�(=�&��g�T����y�<I�s��쪕�5(���y�_I�<����W��=࢙�s,~��&�J�<�feHz����!��3�0��_�<�A,�����/�0�'CJU�<a�)<$���(Z�N80�A�D�<��Ѥ_�IV[�;��#3��@�<q��N�VhJQ-^��B��E��}�<����EԎw��FUa��)Yw�<�蜭7�y��B�ex+���s�<M� �uU���X��r��AB�<�`�Y�y��4�U�uv��z���p�<1@�\�b�4E��M�;�z��G�<��� �^���u�X
W+p�A6��_�<��/�U~�<��Ƌ%�H�)��I^�<���څ��6j�����¡�M�<�q��ml�aapb|�됨CM�<���M�bРiR�H��4y��q�<qP�I>��Qy�˙�;�z]iom�<1� �Q��b��:z&�8P�W�<��e�Ӓ��"l�<BT�PV�D�<9�H̓z�Y�PN��Vo����H	�<т�;U��h�-/r&��ⷤ�z�<��N,|󀑻�#�(G�T ;`�t�<I�,���M 3�!~Ԕ� .L\�<1#�ıVZr�� @��ӰD�P�<i�LN?8�\����A&FdVd�KS�<�&������	RVN {�m r�<!A�\�h��4���C�Ae��R�h�u�<i�j�T�H�KS ��ZR�Qu�<�@�6"ęX�� x�
V�[u�<I�nUC�|ɰa���:Q�	 _�<A�G,�5(��F�%���C'/T����l�H�.���*Ԗ
���#�&D�X�f �&c�&�Yp�T�j���Q;D�x�@� �p�2m���65��U�b9D�H9��އ6ͣ5�P�v�x��5D�ة0EV�����`D"hFe
�$0D�h	�Æ_���oȆI\\D��P�<�UJ�XX�H�GŒ>d໶��g�<� �\Ӓ��[&h����%u��[�O��D#k�bp#�L�6P	�A ӍC�!�!�d�o�H�����?n�����4�axR�8e�i$����ALȳ`b�C�ɚtt�7D^cdrG�5>]~��hO>a+��W�(��qL�)JT1ec&D��r�FN�a����e�0�3��̘߯'��{2ᖄ	֔�8u��\�h������yre�%P1p+�i̎L��c`X�y"�Qp���2���N$��R8�y"�ʻi>�2b�ӬF�ȝ�AM���y��i	h�dF BЀ1:�T��y2�@�t�rW���9rj�*��^��y�K�<}��)�Bז1���7C�9�y�DN4
o�b� �-�`UQ�h���y�LQ�	M�e��K�'`��P�ɋ�y҈E� u�r`m���ͫ�E�.A]!��Y�Z
�0qU�Ed���&#ú?J!�]�^l��@[r��<"���N&!�d��m���Ѳ._ ��1P�ׂ[!�D��R��;��N"`�+��q�!��ٚ	9�.G& ]C��γB��x2�	�"��{���+Kv������&C�
da���Ě�r�pi�)��Z�C䉎9(T�O�0�~e1e'K�B�	�'{��S0�]�l�L!b��C�Ph~B� ~�`��Sm�[t�v�s_B��,6l>�j�� [�	1E��1(B�I�w�Nx�$7N#<�� oӼ)6B�I j2��Y3�	R,<��V	�	�B�i��6�E�ق�&` +�>�y��B�F�$�O_�1�R�@�����y��#�Űr,45*�`)B�<�y�LxV���RA�(�������y���-N"�8"f��\��lеD���y"%3p���CG��J�I���yB�i�|̻���`���F-6�yb�W��`I��Λ���w
D$�yRA��N�8��Z�ubpJW��3�y��0^���a�ȱ
�tŒ5��yB���	#�}ʴ�s�-cE�L��y"��
q��	�o��{@1��y���64>��ר
���!�`=�y2�Ă��l;"LO��LY�$���yrB�L8�
"�ɵtA4-R���$�y�Н�����"�7d��a����y"H>Jt
���,٪y�����y�d��Iv�iv�����2����yB�U
��Q�2��b���1�yrf@�+��X�3���.b��T,� �y"�MD��Yԃ������0�yB�֟_^�m�1��7j[q��5�y�\�. ��s�O�+kM\�A�Eɶ�>���K��~�k	!O�|���C;u�tٓ�
Ϋ�y�*yl ��!@/m�|��L�(Oΐip$E+�����'[5}O�AS�lR�^;��J�"OP�s�2NN�-���� ^&Bd)Ž$�	�����Oʍ)��yg��hd� f`F��"OM�Po�0o`p��B����a��O�� ��9�0>����|�����@R�^6hd���p8�Ԙ1�K ���^%|���G&�ٹ0/�Q!��O�����Dn֘/,����/cQ��B��?qP�BP�-Z��Ź*0be���-D�9q�̀��wKA�޺�Y�dh�
�9�#?�)��� d�s�Ąq���ύN��9�"OVt[2���-E.U���E�}�й3�"O�l�W��9Vp
"-�gΤ��"O�dr�,R	j���J�,�!=���	B"Oj�+���_�Έ+D�Թk���!g"O������Zl�1胧/>����r"O�X9G�g��	Za��%y��9�"ON � A�[���Ş�-2�Z�"O��S������w�r�8�"O���%�bg�y�Ň�#kRa�W"O~0��O9 O��E�E*����l�����.}o4����}�Za���$���ͦzb��=E�ܴgY4�x�H�9R�ؑף�}!t�{��)�矜 w	[�xU~�0!L3�@��A��Иw��q��!��'K��!��,\I�CM-g>��c�'�ax2�������V5z
�Y@�<A%R�X(d`j\��n�M�6;ָ%���L
���H2&��t�f� 	��M�D��͙����UfV,�~� ����520�,:Q�pBE�i쓫M����n֬<2����nt���jp�l�j�Ã�~�V0�v'�O��!��Y�0�&HU<2�P9���ٔ$,�:�M��O��G��O��a��?�|��T�_�M��䡖��y��V�H��-��ʞ�p<���HLQp�Z~*9�WR?i�� )i��tH�[@���#�N,J�K�/Ϻ,�^	�&��n���Rۓ��v���&���X�:��c�݆I]��%���SC]JU��9w��,hJ�0���m̧;H����BL�)��Bu��p��d�t��N=E|� F$U�>�04���_���Tg �b@T��C��R�'��L8\40�s�^16*͉T�[�ZR��DAa6h����sJJ�ql�G!�i0��|�IAw$Ռ�X$Z$B<OT�˦
�}�ba�h�(X�	��'�dI�hR�]�5k+�=h��!(��:[cL������6;�C�!Zs�!��b8��GF�7j_q����v��'^a٤�E�s��HI�!ҭxlzi���i2~z���o�7'+��a�D�4�!���O�RA"É�a0 ���,*�\�����4��@Hv�C*
ي�	"?�B��I`�K] Uΐ�kq�fh<���e��!�pJ�,�p�F*غ�na��X��2�A�5n���;	�r_4��F�
	��G,.G���	�g�̑%��༫2ɝs��	���4o:��&gCjǞP'� � ���M!t B��A�&x�FQ�A+�&y�NE�1
 +��<
��D�&�b>ii6E��Z R�z���$���B&D����!R�IӔ�i!��J��m9��Ƌ}.�۴M����a�D�i�t�D�,O��'��+�vԂ��w\pT
 "O� �@[�~�����U�2����ϙ1�%ç�=K^����p<a�j���Q!g�*�� l�t؞��a�\�a�y���չq�"�c�A���mqӕaά$��"$�d3΃�2�d�u��Vd��ł!��\<�Vh\�f����d"�>�cPO,,u�AhU��yRʗ�A�ƙò�L(:�����M;"ȓ8rZ���K>E�ܴ�z(�VH� M�$�����:&�%���ɦ �d�:t)�� `!l������l�4bd.&��Ĥ�<M��5�+D������/h�!%�it�}�C
2�ӈ��L�jN$4��d��9��Y�#"O��7�˰p��U��Q9d�l-��"O%�-Nns�t�U �i��4"Of`0UDĈ*2��� ޔ��Q1�"O\Hvရ%���3�؛p�@��d�8�ŞHT������2�׿9;L �ȓ;�����B���B��L�U�U��0�`�h���Y�@
���:���ȓ��y+ƢQ��}�R,A!�rɆ���h����vĠ�!���0����oN�Ě�.��}q"��
 c��� ^�:�h��Z|�b �7nDL��ȓ`d�b�8Ǌ���Pjl ��S�?  �ɓXL�P�YWm"s��b�"O����<���ȷ$�yp�"O$��#�1�r�;D"�[
�<��"O�)
�h��B�8v��	�\�b"O�y�s��^|�U� p�b-C"O�0h�GMB*ū��8al��I�"OF��'B�?t 2h�,a`�Ib"O>����O�~� ֿ[f�aaE"O�h1D�5�phIbʞ yEX��"O�׏�T�z��¨G�*?"�1s"OԜ2B� BL�i0�&]7k��h��"Oz�	�Ɍ2b�b,��kB�y��a��"O��`��,f��y
�k��Cr�0"O�QЊ��!�;f���Hɬ�6"O4��V��=/)R�/J^��	��"O��I�T� �h5S�o	�d�f���"O �R$�JLB ߔj3fM�B"ON�񕪒8h���I�O�I5�}�"O��`%��%���a.T"����"O��h3.I%{ R�s"�s��Z%"Op�5�:���I�h���Y:q"O�����}w敪u�p��2%"Ox-2Q��%ʭsI�3|��-I�d�����Ď�	�q[��*}��`�7�	M!�䐟����UOG�j�~������D!�D�:,��{�ו1��T���w�!�$�"d.샃�F�i$��F��� �!�$��S_�$x��G��sЋ�#!�D�.���a�
�}���Y��W
-!�cf]!��0�$l��V�.�!�$V�ʰJ1�@׼�!B&��x�!�׵t��+��B�Φ��EJ�!򄜻N�����/z�d�AΩg�!��ڞv�z��M�';GNx��iƂY����ٛO����E��׊`����yr!/f�4Ԓ�OY�F5yBL�yҠ��I��4�A�.T<�q+Dw�<yȑ;nAP�scHυ>�:�PV�Ld�<���X�~q��p$��U�И`��^�<��dǗ\���*1k��+h��K�Q�<��ŞhS�E�g叺+q���A�MP�<�,ol��CbH:�lZ��R�<�D��*&�\�����P B��4��O�<y��$= �C���DSr��I�<a�*��i��J˗J��EE�<ɄF�T	d�	�W�J{�� ���<IC�,;���C�ɂq�H	���F�<�w��1%�>��e8]�"=	�ODz�<�#���Y�� Aj��A�JPp�<��`�'r`�4�R��Y'��H�@e�<���n����+-v8�ѯ�c�<i%�W�P�̙���lI��C��^�<��	�d�Z�B�)��(�5�U�<�7��6f%�!&��A����[�<!�ɀ"pM����K	u����N��<Q�`A�~��d�*S�p�u"
z�<�W��Z�.�pQ�L�I�E{_H<��J��zS����1Q.�Fx"�х��	�$C��h��ŀ?_�:���2������<�
�>Ju�6k�k���$ԍ!OzL��)`�04���ֵ79B�.q�� BS�!���In�'u4���'K*� ���4�:��3��b�O��e�^	��<�pm`�!�.@����T�s�>��&��-�L��	�L�:���|p���ԟ�� 6�R�a�x4ر�v���ږ�'� �cC���-Y��2+	�:�����G: ڣ��0Ւ��� ʐ}1Ay��}
�S�O�� �qBTA���qC���(9���a�����.�(���S*ɰ��1�5��-#�@#C~%��c|�ĥO��H�FF����nŖ%� �f��T�� ��A+��I�Z�OeFL��3RZ4����WQ�����F��b�d�()q�-QZ(Yb� 	f��x�<���5M�^�pm��Џ�U+�OlLy�)\�f�05(���V���3'H�'��,�Ш�*�X����޼l�aS*��h��M&t�½�nR�A:ay��hr�y#�̈́~t�ۆ�G�l���2�\�s��Dx0g�e;Z˓3��(��Ѽq\��j�(K
)���DyB�L:g��uB�h]?i���6��ē>Rzt!�eB'x��K�(��>���7q�0�W`t%�| go̸L�\q�<�6�?��	��qc󮝎'���6��8CL�|�"#�G�ɔc0���'���zv�K�c �A��02�c�)\���X���H!>���J���#T$ء @�
}��G�#�'D�Q�d� y��ذS��~?�l�-VbI����-|�Z�S�i�ў�6k1$|�����(����$$���&�H�D	����5��A�/O !��cW����%m��ȃ��	�U��=����+���E���f����?���b��4ɒ�ǊZ��[b�c�f�l�QA��g�n+���y#�h"�ц[��h{��&��K���|���2M�6���"�̌!U*����;iS�i� �
�p<A�w�^�P��C!	g6TQ���~�����O�L�"b����O��|�2F����XE��=Z��F��m�'��a�ώSvXi��
N7�P"�+�tQ45Y/ S@V ꜆pP���O�3l(�h
U?��K>�O�h{��i�Y�gp�[�j��
N���(O.��af�1n*9#�Ӿd�Zz��d^0{%�0��KS�bo������*%��X�C��?)�Z����B�Bv�o}�����ĞM3�YK%h�$|�p�QfK/h!��0+��&L��{��K�ķ���	3���ʐ�.4ǀ�1����|�԰2g�X��Mہ�~��x�>�>ܲ�d�1;N�eՖ��!�p��h���h?��'C����
�� ����G.[
�D��� !���D��Z._9l(��^C��A�v�� i��Qjْ*�F�����F�(pS�i��d$}⮶~��aDilޱYd�"w5��U��m��3f$�7K� Yq��4剱<^,�l�n��	2�o%ia��<ѥ�T���A�3 �
�ؐ���Ǧ���ߟ �D!;R�6=��C�J�����o0�ɳ ֥�p��A��I�AX�1�<)jM�I�� ��'�y��'�6쁐�O�*JD��m� F.Tc�>H��%��LP�)Y��$`�x� 0!����t�LHKZ!�B�!��~D8?Y.� ��S�e���z% +;�Ѝ�p�CI�'i���W� 4,�	@3�ҥN����&�>�&��3$�% ��	D�T R����O��7P���i�To���@�D $���g��|
�u�G�/t��m���$�h^t6ʘm����G�N�Q���T�C�[ ��+�	�)vjhxIֆqӊ��O>�1�F-oI�1XC��7@X)S�D�8� ք�5�>�b��(C��┉�)"��8R���9}bA�QD���q��&d��K�'�P��\A,��\�m@�(-O@�ݼ'�� �fU�
D}�6��_�N#=�2^>9w��M���2M�.^��)�ɛ��O6dؓ��;xHp��d�:]��aC,
�y���E}��p�W�/�7m2����)^y
�����(ߛ�Ҥ$LB���a�4t�4Jf��7?xb��.O`��� �9G_�ዡ�
��r|5�I�3;4�˦�V6G���gބW'p�9��'�h6�Gq��͙����M�d&k�eq�}�CN�g	�����d�k�$��5{��(.��G��/��ݯC^��͊�ho�ؤJ64���k���k4j#O��8�mA�Vp��L��,�����[�dB�I�Dm�Ȳv�[Awz���-?�)S��������gCP����E��ɰr�#�>=3�a��ha� S�C]���<ybB�*Q¥C�D��0��Ad��W��E�#((05Fto�ؔ�剀` ���E�"�^�A'�e��<�3�@�`P�-Q䀸���R�	+"� s'	�9d�Fu� C�Jc��+�o�(f����#��P������Byֈ`���?x��|�b 1 ^r�W(b:�锯Y�)��-�1倁 �K+,O�nk�ʤ��'��@�tH��48ѡ��ؕ#hza��dD4'P��@+�0R45�	�'(�#�甲�`��h��l�&a�,ON�쟃E�ԙ˓W�l�Y��׈zR��OB�~E�'u �#�K�V&�����-z�:����_Qn@Kw��>&򎤠��K��=��KÉX���$ (i���?i�c�#YS�,�!H��1^��37G���<�1��\�����Q������N�_v���f��)49�A1"�8
����a��H8��λ2�%�Y\?���ɯx�t��u�YS!��:W�� ��Z77xp[Ǔ��]�&+]`���eE�:VTI@֮8v���if	ܟ~Y�@2AX������}�̓&lBHڔ�g�L�����&/@u�g�s~kh�^���C�'��mن!���(O� ��[eb��m���I�jA c/��ڧ�x��Ţ F^Qa�G�0;+L�S�e��'���ŀ?K��0�uL
yZ�A�H9p���P�C8�L�R��9v�q�л=�
�"��Ȅk5ڜ�e��QP
����yW��4*dQ�Q�6	�t|Q��ϧؐx"��D�(! I�s���a��	�s��?Q��m��H�׎	gP�tj)%u��p��B�s*��S�ힻe�C�4N3R�'n�T��|sF�=ʾ��	�1��\��U�p0T��c� ���l�'(�8�6�E��Z��+V�n�T����tڲ@�D�<$�Z��ѭ2(�	"f��!��ͯ.��d-��i.�I=Np]�Rf<rޑ@�S?B���ǵk��!%�������nQ2�EF{=��+c	�G�h�	s�d��K^8����?Y�M��h��`5���∨�O"9����8�QE�D$A�VΙe�'�<qZ��V59�t� -K'­"t(*md�8����f����'5+ayrABM:4���7�V�@��/p�Ȩ� W�(4jH�7�:#�.�բѪ%%�*h�Ѹ��r�%Fy���1A�ؔ��nϠC^��p2EE�ē�i��l��Z�|�8"��u���>���^�$+H)�Ӯ^�v�� �o�Z{�$���xm��$[E�I+xȲ��!z�B��P@=LĲ���{�<�3'Ԫ�p<1�w�t��tT��p�� �l]��'�x�����k�az�%��93�.�FXj��� z��?���̟#
�e�]��?�C�(�r�9�薘#� ��]�"_�`��q�� "�C�jžU� �@�t��� @m�T�r���6�<��^��Q�/0:�I���'�n-�IKHy"�i��8vo�c0
�B�p�`�3�/D4%�OZ�@cjO�(�8�tV���1��V���t;"OX=hOL%K4���맧W�C2ԁ��\⟰�S�F�^:�u9&GH��Y��c@	��Y�6��Q�"c����F�F����gC�\e`)0
��y�L��0u�MP��F�^��MR5*	Ʉ(
Q�i
R�Iֿi�ԍ	��:���!i�0ت�Ate�$[f�	��0�d�d�Дʕ`��N> r�Ǩ���0UF	�=�<ykO�5w�x�$�x���O�i	)�q��'q�]q���%�	�pX�0#���)dZDq�V�`�Ǆ�r&�h"��4��c�+fy��P47��	!k�"��P��[�;������s����}_z�S�ğ>F�Ė"QZF��'�I�l?��;f��9_�]#WO�$TN6d��ov������<ْ%˯)w��hd���?��"Q�������h)Hlj���c8���Vb���?���ԆZ�82
���� p$�<x��#2j�f@yЇ]��?�U)� �f8c�ݰ<��˭\1"<�oجh~�+�#�9.�џĊ�$�!36��7�\�d&8-�t'O�G'�m;6��=�ƨ��|�X��	1N���S#�	dy8=�����-@��@�E���L���X[�b��-O"	 7	�""�씈'.�^��y(�O0��F�X�b �
�6߾(�'8�������,9UOX��+�=����7%|�����R�	���s&ƌ;ǐ�q�(��WK��6`� Z��ͻuA7���B�IC�	�w.֬���O4����%0�`�S��g[Ƞ��L9N�NX �F5A�Q��IӼ+�ݓ<�:@���^�y���+�Z��<�1��l5��+��� �F~��>>������>�"A*!d,'��?�R�K6�y����yp�I��W
u���(˶�P����O�H`�Sc����O��y�'0�}�A
�Z��`J�0#�Q�������0a�xyB�C0^�� C۴#���5��8���rp4MZ3�	yC�i!A`�\`B�K�ʹaPЈ1�x���)C��jZm����\(��'�H9�v	DtĐ��=U�08%���	W��JBKX<I| ���sBH8�rҾ����� W���;l׳q�N��+rf(p� ��S@v<���KX���gcv&֙"�9�D�HVx����:J'�(pϘ�md�`���ɸ[z��b�G
}]�d�T p���a�U ���I=&������%C������C�~�e�Ȓ(��"��_�8�"��G����S�O=d�N�Җ������XTleÉ�������+	���,�~�qv2��D�c(x)�E��]��Ā�^��A�CIjD(�g�'��D@�KS�V$�#�'��ND:x�#_$x4D�I��2�����:y�'4�l@��I�1���zC��C���Z��?T��DF1]�� ��o�I�֮˿A��(�l �"莤*m��DV�gy�O=��uHG:tfx�V���J(x
�'D� �R��-N�M@,='.4�
�'*z��愑��%ц���r� 
�'���(�,�O�$�b�ې�=�
�'� ����Ԩ,&F�CU�L�B��B�'�Dd�4��w0�4)�'�6U��'���XAIT�B8б+������Z���TH�0��aH�q��I�ȓyPp�A�t���
�[�T	�����f�1c�4�)�+Q�������5�P��0X�+�cKV��S�? A�m݆Q��Ti�������T"Oĕb�N�rq�9�d`C>u��"Oj�C�+a[�퐅�6"+�5H�"O�x���1f3Z}� 	P�3~�=J�"O X8���3g����gYnG��"OQfkQ����y1	�)D��PG"O�y6&�4O����s(��i�ԉf"O��wi�8�0�qH�E����"O(��c:l�*��&����Z�"Ovx�b,�1!X��%�=<{�1�7"Ol���)YaGf��%Z<*����B"Ou!G���)���D� O�th%"O���w��n�2���+E"O�к��ݤ?��ѢC�Q�$*�"O�(�fHJ/6�Z��"�i2Z�"O�� Gg��$$�0g��x�"O�0Tʇ5UOX8�Ҕ�D�"O��
ԢǋJ�xyk�b�7=bIp"O�I{��Z85� ��+}��y�"Ol�2�)ٸc�ȭ�Q��T���{�"O�m0u��:Ad6��a.�-Z�Z�"O�T��*� C�t�&�Z���݂�"O��X2˗�肹3E�W�E�Bak�"O�Ff�?fF�-���]Zh�)�"O(%���i[��KSB���"O��%|sT\:�$,#tq"O��Z ��iu:,1D�^V�a�"O�=�-Z D��k6��1/Ry�W"OB�+��%-@��\�E,�<#�"O�usF�O �D��̀!l�H@"OrH����/3�l�g�	'ox���"O�Ի��A.��2�*��f荳�"Ot�R��"^6��S�KMW���"O�J�&�@}�,jf����"O.|3`m�,wo� 2�!:It�S�"Oԭ���´0��dZ��=/�=P#"O��0��c����Ъ�4'P�:�"O�!)Ѱd}p�2���'���"O�1B�l�
}~�`s�� �	��"Op�����lZVT��dq�Tp�s"O�U8�ɊtppAK'Ë�ܪ�p "OX`
��ؚ1;�yH#��$��C"O�Q��P��6��s��q1�*3D� rRm�,'���䂖 Gn�Q�0D��3n͓SOP!��B5� �97H#D��� ~&(�^�$�ql!D��������X���؅	-U>D��y/�6K����q H#xsJ��g�.D��p�۰[�z������l�X�B 0D��Z���D�Ҥ��hX#M1x�H�@.D������A�,���F��9ْ��)1D�P� _�vtЀb���4��u�u�.D�;P�I�9b��Ӏ7��!#-/D�Pz7��5AG��k�iQ �ܠ��.D��KB,�x�J)�G
N�}�4:h,D����G>+����r����t��0D��Idfƾu^�	K��D.|��@�(*D�@3�\) f�	8"蟆u�|X�bg(D���1�O7gz��_8rS\Y�A&D�@Xr�C�%B��I��x�p�1�"D�d�FDג���i�>g�,��U�?D�xa!�3D���XvKZ$t��i҄�1D���� �j�x��X>K��#�*1D��*��סA��\) �U�Eb�P�j4D�� JI�!��+]�H<3թ��VE��"O��F�#4���S��;[d�)"O�}�@o�;p�P����i��"O,�
1��-gl��r�F9�29+�"O*,�b�:\�Pmade��]�F1q1"O@5�F��	c�H���(N"!D"O�����;`fbPbq��-^(�"O-x���R��W���hqB�3�"O��f�;t��-�u�K0U�:�"O���v��/PU�`H)%����"O(,�Ug݁H{���1'�W�9�"O�� $�N���{�呷A����""O�I2a��93&	1%L�*���"O�� �N�N�)�<a8��"O�IA�;3�@(�[}[X$@�"O�ԫ@D
�=����bL!�(�P�"O@-s���qu�� "��0k@"O���F�7.�@|�eL �йQ�"O��x��05�`�U�5İy*�"O��j$iZ�����*K�{����"O8(�	E&u��12�)6)3.�c�"O�=��� �\]��ȃ�^$lu��"O,�{��œ?����>VrZ���"O�I��ޚ١B�MXj�"OŨ�@ӊ{����'AչVX�IB""O�-�ԧG�8)�R �u$P��V"O�����6a�����ó Pq7"O(!�5E�v�Vq#vnٽR2���V"O؍��e�4 ��dk�CY�F� �"O h(�.^$v�.�c��ȄI�� ;�"Ov�x�l�>E��)$Jօ�V���"O�t	Kѡ���[5���|�da"O�,  mR�!)���ew��1"O���#	D@$4��F��<h�r�"ON}�1�	�Wq^��0T[Nlq"O`��"fA�Svl"�&�<
h@)cr"O̍���Р?��	�FaYR��y�)ϱ�p����82�ȃ�e�9�y⮌�Y+p�DO��2Av�q�9�y"�ѦQAN� `� ��#��,�y���|E�SU�Z�|�`�RL�$�y@�55��`��ƃ�b��B�S��y
ց�9cd[�_�:� �m��y2蚣� ��%/ՐYgu��0�y"S4Q��@��E�0d	`yjcD���y�L���t��X�\�83hJ�y�Z�p�*�# A	�b>�#fn�-�y"-D'$;��H@�ݫX���X5����yR�M���%Д�L�ر��#���y�I�r��5��ў{`�b���y򇜹&(����"x�F��HŸ�y"I��	��i`��["&��C�Y"�y�ɕ�2!�Y+u�����Vk�yA�#J�F�r�L�dҼ]�5��!�y�-�U*�9y�fW��b�����y��r����� !m��s卼�y��o4I#�Iػ�Ju����y�i_�BJ�z��5���iTCS�yR�ƨ`��h��C#M�- t����y2��>K� � �r�<�`�y��E{Z��DY>n0�58b���yE���U��b=z��0���ybF�-|:���Q����T�y�?�,�z��� �����y
� jYiB�UƮ}K� (y8��@"O��rA�O�)3�0s�MB
E����g"O���7J�k>Ε�7O�%�^�ړ"OJ��W�z��;0n4<�H4{Q"OЙ8���?*�()���Ѳ" �b�"O��{��H�0H]�g�O�Cؙ�4"O>��$ٝn[�1֊V�l����"Oʭ2P�u���C���d�l$D��p�$��j�B�x �Ўw]���� D���c�
,��1���Їk�dA[f+D��jЪ�#b༅:EhI�'�*���-D��yg�U�lt��sb��i"�A� '%D��:��� ׼�с�J��"D�㕩(E&�d�r'�>P6���g D����`�%�(bW)�<&޲8¦f=D��r�C$��n�`-��,�zB䉆>2%����F;Fd0���B�I&4��Y�\�FLYB� �C�Pb.0Sv����M#�67'�C�I�d�Q6�_R���g�-}'�B�	��������m��-���60�B�� ^��A2wg<�|��UOZ)!B�IV`��ƻ^��0#��%�C�I ����9XL�Vɛ�ns�C�I3�Z�c���p�0$*DJ�8j��B��(]K�2&� � 2�FI�/O+BC�I?6�t����6a*�psb�7lJ8C�4+�hr��Z(d@�:Gڦs�ZC��7.yJ��f'��@{ԉ�y�XC�I�s���z��#	��b�fZBc�B�5y⁒g�XC���
���:(B�
|&r�K!�/f���q��Ȥ}�,B�ɲGdJ��#&hA�r��uO�C�I/%Q.��GT���i�1o4�C�ɲ*���f:y�4P3Ý-2��B�I�� �@�#��A+��B�	�d@�!W��28u�D�)X�B��5Q}$�b�A)Fr%��M8?�jB�IDފ�t�gIv��1�-U�D"?������f�F��X�8
ԍ�!��\X���#�b��)�M�w�!� $]~��Q�T��v�p�0"��C�I	O������(�B3VR�$��C�Z�ܑ'-K�~��b"��i�(B�I�w�����I_���|�RH�9k�B�ɺV>"�9QO ''B����|�B�	�w��cŤ�� 0ب�#��p�B�,�F0��]�QJ0"� �B䉯V���D �(B���)�J�}��B�I;@!U˶�Ɋ]�����m� ^��B�I�*V�r�)K�b|>)iC�V.v��B�Ʉp�*}�`���b!xƪ�0q�B�	T��A�U@^�/4�0�e��`%�B�ɶ�b]∜�v%�HG�E!o�XB�ɚ7�؜Qf�-Oʹv�^"RS�C�ɝ7��ّ�ע6�V4��H$+�C�!�Z��۠iH�]�!�׌
pC�ɿr��m��
��7�Ģ4X1I�DC�I�:"a�ܙn�Ʃ�$��.�rC�	 {r�ҁ�
�ą�wjX�j��C�I�;5�1�F͟�	�l�c(W3']�C�I-�p7 P&O� 0ZV��r^B�ɷ.LD�q��	?(�E�E�n�B䉷SN��D��p9�ҍ��3�0C�)� Q�wB�-L
�˄UJ�H*0"Oi���\ �'�(ED��$"ON���P�U�$�hPG��0 l�"O���*4�p�¥�(|��4"Oh� ��71��T��G�Q*��"OL�y�
�vq�j��\+!"���"O~��A�?����pѧ]� !"O����'7;����Y�`Y�$�e"O��bE�(2���M�Mdɘ�"O��y�c�#_9r�ꖿ <l%1U"O�AC��2��������Zd2T"OX3a��b=D��u_@x�s"OxU
".�?�B(��[�Q1�"OtԨ��I� �w��B���"O^�+��D�9u�1 J�X5��r"O"�8�,�P����B�'^$ d"O��)�Áx;|���	#p�B��A"OQ��/�,̻6߰6��M�"O89�H��+��)Wj95����<�� �+���&>$2
u�F(D�<��I.,
��C�L�7 6�I*D�X�<y!@( ��`Y'!�4.�LeBS�T�<yedt)�W��P\Ń����B�ɵ &h+��K�{Fũ6lو~��C䉹]4�@���ٓ%�z#	;
|B�I		o��y򫍀�(�`�`M�,:C�$MG�tRE��0����vC�	�/�P�
�eO���i  Kיh �C䉷��l��_�G�<�R-�VHdB�	Ĵ�@f#�Wd����&bRB�	u�
�����3�����c�z�0B�	�ŀDJt�:��"��M�JC�I�*�Pq��	.d�Di�4�LC�I�)U�5�%o�4���b^�C�Ik��S��3��Jbc��
C�I�?��\H��@�@�h3Ι�I��B�ɑ2�N@���Pbvջ��1��C�I'KI�ҍ�5:ގ�q->f�C�	'[�� �אS���֨�'l�C䉔vzLApˎ�a�:�b',��qYB䉤a�)&��	 >�!��@=-3�C�I|I�d���G�a�G�C�rn�I3s��']�L��aB�C䉛Z-��ZFfeT #K�A��C�ɻr�,Ii�޷$g:p���t�B�	��H�t��8�r!��*�(B��C�	6��8�N6>lј&H�D�6B�I�Ga.��2�IH"��A�*�0B�=o9� ���͈ OLj�� ifB䉄Dv��ف%�(9-��0t��/c�B�� *n�p+�!�5�؍���*U(C�I	���F�̓Y{^U1��S�C�(m��<�݃L�B��d.W�AK�C�ɛd�B�S �? �T�#�I�0B�Ƀ<]��*ŉM,rg8�+eG�^f�C䉳F��i3��ˆR
-)$cX0��C�'��)jA�C�F
���P�T)?��C��!t�D�*r�W�  ���gجZ�bC䉙8���A�I�iW���0�׻�ZC�ɥ|ߴ ����&	x$�s��4rzC�;b�څ�Q6�B:0�0g��B�	(-
p�!��W�a��鳎�w *B�I%6����ԡ�(M�*u�Ӣ_6B�*��m�VO�f����K��m�C�)� ��Jt�N=���nT�dӠ-*V"O�aP��-?H�ۆ��^,J��"O4Ӱ)Vp�%)�k�:���:�"O���&U.a<Ő�)Ǖ�HU�"OE�q�M2z�<�cB⎗Y�l��"O���a��
x���T�Y�X��,P4��9\OX9QŹGz"���.N��
u"O���rA�3f�����RM�d�V"OPQp�T> I��[��̉I;Rd3�"O�@HD�Ku�$��.�EJN�PW"O����1oq�%2FN�Vl	c�"O4�3h bA�T�"��=,�١4"O��#EM%4���
�4��"O�a��ҧ�0ɨ'�B+=Ԁ��"O�T�DU �IKs�C�E�P���"O*q;GɎ�!ǎ�E��K�^�:�"O�π�|�,;Q���S�d}Q�"O��(S��(5��%��V��T�� �|�)� {��6�X�-HD Dj;^��B�I�E�X�y��et��,�=|C��+{3 �����qP���H�"$ �C�I) = |���}��A�o� D�#>���	�B0�t,e��!�
 �/��$N�xF{���喩"�����V:r;R��%������O���ا�8mQԭ������,��O��=%>%�mD�g�:�	؂a�xW)0D�(��	G6���Þ j�@���)D�(c���0|�g�øiT�p�2�&D��:u	_(�|�1C��H�@�&�6D��q�a˸-|FŒ$DX!n�Lå.(D�pC���5�Aö/���	�W�#D�P��ݡEq6�W��9��c��#D��+�.֪Ib:��Ԣ�L���p�%D�����a��A挨O���T�(D������#`�ʷ���cDh<D��H0��!"FUC��%Ch����`<D���3k��3���E&D���,�f�8��mܓ��O���S� ��k�h)�m �3 �z�'\��`
׸=}Nt�l؛Y����'n��1����j��!���iY D��'�ح&�Q9n���p�.S�b�t���O$��)�O ���e�	3st�a�*Ƅ(]hݪ�"O��E��"�~ݒը�]L�+W"O�,�u�K�7��&�`GX���"O�eaRa�oa�|j� ,���C"O����I������6Y%j��"Oy�t��7C�8���J�%t��2�'w�~b�i�$,���rj|D��h��L�Ó�~����0I�nQ������ �`¯,?!�d�?`�T\(��3d�zh�l�3�!�Y$�C��Ȓ鸄+�f�!�d�2t�N5����$��ay�ڟ�!�DC�c�x�@_+A����(W��!�$	�$]��%i,���!&4
V!�Ğ#Xf��Q�D9b&>�Ȟ�!��"J
�ѩ�(�;7(�φ<!�$�.���3�ᐂfǪ�dP�F�铳�>�B�N�L;���� �,l��IacD{�Ik���O�ʵ��Y�|������#�*�YO>Q���0=Q#��en�8J�dE� ����u�����*5(�Ъ�4TQCԎF�'����M������z�8�I���>S�̳U�%D��
�
Ly"��:�H��S���x3�.D��{��A;]p�ɉ+q�҅���/D�� ���tΊ o3�$�qĞU�`���'!��\�Ii&�� ς�m-�L�5L۪u��B�>K�xM��g2��ţׄUx`B�	�o��yRTJB�J>�qXalU.u.B�	=G{��j�EH�`�U9u��QB��"+� ˤG�M������4C䉺A4S���{P�gN"(��7--�ȟ���(?���k	�V�ɲF�?��'�ўb>5 �$UO���[nA�H%��e⩟�onx��2ŋ"�j!i�\���� �n#D��z��X�"ò�!�
!Xв�
�s}2�'���gY>;3�T(��ա'Ƶ
qf�.�y�$�#_r�X�,[�$(��͛?�y2�U$hZ���ܤc\�Á`���yB�O�h�^���ș�o���0@*�y2O�v�ܼ���	`%n\A	��yb�/�@��"��5Y����U �����'�uܓ!S(T�J)t��@�W�Q�e�j���v�C�	�<��E����<B�:��2b�0���]�&��-H��.����	��E�1�BA�ԏ��_%��Ж��:&�!�e\5h@�
N4�/ݫ^t!�d��	���R�c֪X�N]�`G�?zT!�U�r_���G@�$�*�/���!�D�t�|i��a�T���C�V0c�!��ײ`�0 �.U�G> R% E��O�=���O��@��f�»YZ����j�<a�A��7x*��J@�^�a�c����	��]� ��u��u�Б���b�V��ȓv�]R�Ú;?r�H*RΔP�mZb�������]�8V����ڛ@����`���y����p�I̜1@��0�/��y�o�$0D�4�Ϛ=-�X����V�^�6�=E���\Ah����!G�UqG��MO\݆��"��0i�[XH�����$xÜ��ȓn�}�5�M-E����ҝc0؆�I���-\URA�Ü�M+��΍\�B䉕L����g�Q)��u �N��
O˓��S�'���j&KQ�3-.��@�y���ē\�a�N�3�p�KEK3<�B�(�iN��?E�,O��I/O��Q2��,�x	�E�'H�x35I �%��qN�-@���D�;?	H<��J�@!��M0�p�$�Nz�%�=������ě,V5�P�[�Jq��@"�ڣ�y�K>@n�)���!A�:a���R��0>�N>Y�Гg��9J��Α}y
Q#"�~�<�A��<7t)�E�&���$��C}�'��X�"Y$+�#R�λx��]���?y�O�ȣ���4>�TQE§A����"Od(��U�y�ZE�^V��IX�"O�A��L������3g��>�}�"O�xe	J�+��
��12�z�,�S�i�1."@�B�-�z8! '$�!�D�Q
p�&��I�Jy5��� !�d�hSL�3��J3B��!�o�.�!�D�\��PA�O�J��as���T!�d��i��!�bL�U"g��EJ!�R����CT@��UB��E;R*!�D�<;��{���,Jݺ�xwF�F!�X�xG�4ʵ�߁j٦����=!�D*z�������(�m��Q%�!�ڨ~�9٢�
К�qǌ�4)�!�?:�|h��?�"���;�!�Ĉ�-`XMK�d�S��A�G\ u�!�� ��1����o�=����Pk؍�G"O���3�޿fƸ����X��'"O�8c��ϙa��2g�Бd&�ձ�"O,���f��p�^yS�60f��"O��赥M�^,ƽ�(Q(����"O�T �`I.r�4|�`�	"=FfL0�"O��ٲ��J����`91�X�"Ob��<da��R#��h-b5��"O�����r[����/ջ9����"Oz�(A
�"B�<���[�3N���s"O� ˕�W[DXp��^�v��"O��ك�S�x��Azb���M����"O,��ɣ������:�j�9!"O:���O-vM��3�>�٘�"O2�Ҕ@Ou�9
`�Ȓ3����5"O��@"˼U��0������X�"O����3U��E�ʫ4��"O�=ؤCR�I�"���9jw�t �"O���t���dZV�c�ܘg�A��"O��� f�?!0�u�FL�F��T�"O���Ɔ͑d�DUJA�<a�xr"OR<k��z(�!����P�V"O�Ա�ԋ22�B��" o��"O�����"|u ��0�Y�RmY�"O�qZsfU�c�	�3��.	�
�9r"O�ʔ�͔PPZ�a��]�
�"Y҃"O�A��a^@h�#S�/s��8��"O.9�G�]e=�����
#�e(p"ORp@AiS�SJx-��O�'��E"O���2��4;_V���a�f� �U"O�%Z���y`�yQ�P<x�P]��"O^�"�k̹k��=b�N-'����R"O��@�,� tk��A,s�ҁ�p"O �b���G|9"r��]
h��"O����A�:�Z����
j�Z�R"O��aZD԰�P #ѩ<�&tZ"O"�1��ø[���#�#/w���t"O�y`v`X�H
@�v�&UZ�LA�"O�mP�M̪f��B��ڊ`3B=1�"O^��BF�G.^���L)nHph"O�\#���; -x@"�
;� )3"O���v.I�>/~���c]�<;
U"O攨#cۏ:F�)vbR�u%�a4"OH}8�*�[0�����jq`�0�"O����
�'�>�
SW-�T���"OX���0b��uR�׾8��<�4"O�5����H=��M
��R��"OF�#V.����!LC�u�X�"O$%k���/&|};�+�@_�a{3"O�Z��E�n}�͓�KۭgZ���"O�T1��(Qp$iT%�HB��3"O�x����Z ��ڴ"�.
'�M�"OVm�#L�c��3Qa�p�y��"O|$�Q![>�̩���ֺUb�8��"O>UҵF5 _�ч��$9U@m2�"O<�ʃ��rO�dpQnŀ?���"OƑ1��\ztD�!D�-w-��y"O I`D �Cz
yC�B�B�Y'"Oy0��.�@�9�Ƅ�,b�"O���&_ͤ1��!`rl�c"Or�Hf
lc��k��T	ZR	%"O�iG���N^8ɀN׵HMN��"O tA�֒:t��`ֳ9f��"O2D:�J��N5��OZ�O[����"O� "�;q�ϳ2�\�G����#�"On�a�47�v���V�f�(�E"O��;�O�]��ݪ�i�eҩ�"OP-�P�Y�Z�| �#NU>�+r"O�X�f Av�	��Z��|d	�"O�i�歓�
��*�aO�S����"O��;tN��L�4nR�A}bu7"O4��cϕC�¤��H7xj���"On0"t��)��]Â�&)X�]'"O҅h5M�	};+$�:Â�+!�dYa���� #�4rp���w"׎[!�D� ���p��NR��v �Z	!�$S A|��A��)E5ҥ�2	>�!�$�1���� ��ew���5�0u�!�Ě6Bbp��^�<q�i��Qi�!��?�$�1�eJ`a�p�'��4?�!��ڍn�D���@�LK��#gk�;�!���"S�"8�����<
�RU-��!�$� W�m"�͚h�|a����!��;ss� �`�K��1[��@(6!�Ğ*r$���d�P2�y��CN�F0!���(#��A/vӼ<k¢�[q!�D�7f�HQ�!J�]کʦ�;q^!�$AzG��8�
�>?�4 6�DWT!�ٗ$ a`����,;z�H$��� T!�
;g=bd=	&f����P�X�!��!�X�AE�]����I-w�!�$R�:PqĂA�>\�(��}�!�D
>I�q�%N�����eT6g�!���
�]K�P�7�M�����D�!�d�=��KJŌ|(!�mL�A!�$�l�␀R,�7@���S��_�!��R�=T�`hB��u�<�!��T5X#�ӄfj��A��+�!�$;M�� `A�	#@8ēT�!�D�0ts*�q��&�0�BH�@!�d
;cl��5�O�k��"���i/!���zY�	 ө�>xFк�b��\!�E�X�u�J}�85�Ɗ�)v�!�dD(\�@+ҿj$̥�u��5R�!��:�\9�M"r9ɖ���#i!�ďf�ّeX�ec��p�f/Y!򤕦%�1"sNM�s'6e�ᇜV!�U!D%3�۵9�\ِg �HJ!��Z�]Ъ�gcˠ�x9�&eJ�,�!�䐊K���c.F�I�{DV5w�!�$U,u����6��uɵ�_^�!�DL�Y�N��7�1�hdQf���e�!�I�xH1�&�O%v��E�&��WZ!�dе]ʱ���V=Pd��D^�RQ!�ȳrDL�Y�j�)M���[P�ά}�!���Lˀ���LԼxز\�� �1!�D�I-4��h�
G����X�I!�'�lᴣ'���#�/�L��4��')2!+B�9e�$D v)@G�RЈ
�'Pȅ¨�4��ő���9&,m�	�'�fi�Þ�Zx���Ğ�-~���'J�h�&��,H�Ŭq��'��q�h��LkJ����*y�
�'�1B���052t	0�
�'F��r
�'{�a���$���A$Gհ���'����L�<��)��'�+r���'5$h�rL��B`��8$Ֆ+����'�� �oʂźg������ �q�6�A�踀0]�j��0�"O*mxU�Y�q��z���^�q(�"O~���K� �``	�AK��M6"O�Cen�n�98 �<���""OB4��Y4v$}À�'h>h�"O<Ҧ�Y�\���Ɂ'�@�Q�p"O�Q �˕�qv�s@�G7(+�S2"O������2UJ�P��*z�A"OP4HT��2�� �Fa��U4�4(P"O�*�)�0Ϙ �s��/i�XU��"O��д�^�&d����v�4��"O6ur%��8��x�U�q�Ÿ�*Or9�%���p2�[']w"l�'J�Ղs�Xpw��j�)��Z
�'��\Ç�y���T���%A(���'ޚ)	$h3&9�4�7g�=$,�J�'.z���x���Aǭ#����';|(P�`MT.v�I�M��2�@��'J��*S �����2S���'����#��~��YTC�#lN!	�'�x���.�쎘c�d�(U�\��'q*q���.P�*�"`�%����'������.u�BG!��4�l��'a2(y�U����D��-��(�'�x�E��$&d��"��۴w�j�*	�'��̢�������2�V�t|P���'��铺l��̡D�F%mҔ��'Z��J%��12$�Ѥh�Y��'���ՠ�8#�,t�����
� q��'�XP*�I�$4T��iڰL�"�'U��% ��X5{�k�	�]c�':���Vb�^�� 	�8�Όz
�'�0���A�( A�44���
�'�V���j|,���p#O�$�(�	�'�,-�3�צSnE�@�=/zhP�'�B����"�&�����7p�	�'�~D
���s[:9�v,�ì��'&�[�RW8<�b��
�RŢ�'w�D[�N�I�hy(��tI����'עA2��*4�0=�J��o6HR�'��i�Fۧ '�(���ެm�Q�
�'��a2�ƃ�K� �a��v8��
�'�<�d,��6b�$C��	�'�B��b������ٵW?���'Ѻ��I��T��t� ��?���[�'�>$bVeF!,Ɩ90fԎ<�V�;�'�!�jH1qt���TN�	3]N5I�'�p��JP�o�@E�ߥ�����'$p ��΀X|1�d�ɨf,��'�2`f��"-Y�����}d�q��'),Bp��it܀g�y��qA�'����p��!My�0�7�ՌlOh5��'%<��u�+�
챗N�q�����'��h�cTXZ�18P�	=i��� �'!l!� ݂�H(@�D�)ih�D(�'S��`'o���x��J#gߺ�`
�'?L�˱�N�[[�l�t#��ID(	�'Ŧ�S�d�<i��U:	���(�'��9Pn�GW��+�	A3~���'�lYJp�͔��e���MG��@�'�<=���۱z��7j4xQ��'���yw#Z~:�hW�&\5
0�	�';ZIkE�� /�0��B��>u���'w\q�w�@'R0>i�5ϊ:�.�h��� ��ED�%�� ��۠,q8�z4"OV����z�y�
�R�&`�P"O:�[���o�H��#kX=*��3"O��¬;�,��꟮Z�E	""O� �D��:^�J�K�,�0RhI�u"O2�ҳ��U D��@)G�(��"O�U���@�;L`�7�	H�vM�u"O�)���L�e�����k��!"O�!4��:�5�@]�dJi;F"Oj8	����*�ڌXgaD!6<���"O
���@5q�
�률�d42�"O��RѤN�[��H[�写,Y�%S"O����@�pݲH���K_��=�W"O�p���??�A�$�
�u�.4z`"O�a�F�_*�te��J�P��}ӕ"O �#�7. D2�f
�y��!��"O��@�ˀ�Y�Дy"gŦ5�(�"O��񕁆�W�V5
geO>TiL���"O�P�4�&I���d�'cfj�r�"O��j��O1jSP%Y3m�2Uk��*�"O���M��%��R*��E�<��d"O*	��@�:\Al���S8�2��"O�is �E�dxGIײgъ)d"O&����3"�E�Hm�H%�'"O����M̚H�!3g��8�؂�"O ��"���Vw�Y����kh�i��"O����K{
.��
_Y��P�"O����HM�`Jɨ g�xSb��3"O:4�p��.�
�JDe�d�4H2"O����kx��	������c"O|�㰫����岧
��~��p"O��򠁐!W�l� hĢ)S��q"Ob�* ��fx���0R�Q��"OeKd�Фt�\l��'Żo9$��"O�a�#.}R,AS��E& j�"O����*A/��1���D��f"O��2�d�Y�&�sҢ�8��I�r"O�=�`��5�ةQB��Cu� {2"O���F£�X՚ fH N�XHc"O>�gG$s1���F �K���0�"O�����K�
胇cM�s�dĀp"O�X�Ol���㳤?fn�� %"O�P��퉁S	�y��ۊiƼAV"O��ҁD.=��!)C�C�L뮜�"O"d�R�L0��E�
L����"O�=3��R>�.�F$��_�.��"O�eR��ΝF}�9ô���X�&"O��Y�+A�v,*����� yC"O��ڤl\�U���r��j ��s"O�x�� !������X;|	C�"O
����L�~d�=ڕ ��5���1B"OPX� �κN�:�h�J$j�R0"O��g�J�2��ckF�m�D���"O��$0�����¼8�4(�5"O��kVd؆�i�7��Yv"O��B �g��[��XL�,e $"Op���h� ~A�m����+b��[#"OrB���W�4:���T�м�5"O��I��׶~kHm����$z춵�#"OR�S��J���ʲ#��&�I�"O�U�'g�6]*z�"�Hq��"O�LJ�_�ޭ�g��VY�M�$"Oh��C��u@v@�"uQ���U"O���ш�� ��E�ׯC�5��ST"O� ��Y�j�?Q\>LHf�A4�1r"O@�q�'c����-G�LAkr"O�<q�f� e���ij@I9�P�v"O�@������d*`�\�<F��4"O�2�/̬u�.	�!�42��U"O���N_2�y�t"Ĉ(��q�t"O~I��)ƗD�F��!$:��Ay7"O&˃I�6g��ċwC��
d! "O�x�	-���t`Z%!���P�"OD���i�2�|��O��Q�C�"O����ʬg��e)�M��>�.(a2"O䈡��9
�R�t��(�f�H�"O�4($N\ABЄ#�j�*i�8�c"On��q�C�W�`�y��ͩ�"Oڴ:�@Ðkl����I��B%��a�"O�13'���*�#�C���D`�"O�ȻB���fft4@w!�����7"O>�2具XyH5Ѵ���ʝ��"O��f�Y�p����R�z���e"O̩� dI�����-o��"O(�a᛿-!\
�
ћ*]2E�G"O�c���%.���
׊xnxț�"O�9@RV!j�l�sEO	)_&y#�"O@} �OQ!�F�2�nN M"��A�"O�+�/طEs����ʚ �h�"O\x��X�F����J�/*
�=2�"O283G��<6�T��9+���7"O��x0�W6C�z�0���h���"O��*w�X!A,4@�'M����"O����������+�a��H�"O��	��wA�$��)�@�F�p"Oh�2L�3�3B"����K�"O���r�Pc
��t-3�"O�iK�A�E8�!0e��gXTA�"ORI�P��,iZP�@rIUu?����"O��ЄN�Y5j$��}޲���"O����P���}sB�6a�L�"O�x��'�X�!����mM�t��"O,A��)�c�N�	@d~��E"O����N� h�p�����"O���ܗ{Z���'#�:T8]�C"ORLCf6k�~�Ip��*�"�A�"OP�a�坞K�4�C�����NĢ$"O��rP��0���z@H�w�DYD"Oڠ`⏓"G&&�� ��e�"O4���.�_�ڡ8T@�&���R"O�@JU+c����N͖H�d��%"O �����!���J�%���R�"O���/������J'� �ʓ"O���D�Ѱz�T�C�4&��c&"O:�G�Gr�Z�% ��ٛ"O"	Ab��0K�.�Em��<ђ"O�`���ӗg{T	sE$S�i�4��Q"OB$��&�6܄�4c-e�'"O�]�k�5 G@�sÔd���"Oج��^�;^%C@�̾5j���"O���K
�;��*�� �]37"O0P'��`}�M��d
m�t���"O���įϒ/�:%���:_���s"O���%U"�n	A���S�fH˃"O�����J���&!��u����s"O��!�.�3^��p;C�G [p��6"O��"CA�#+8(*���:Vr�l�%"OJ����7Ô�g��4��a�"O� 
dٕ��
܊��PC/3��)�C"O�pò��Y}�`���X����r�"OD9�����j�*�ǋ9��e�"O������O8��!���?h@��"O:��ɚ�	 ��%o��-�	K�"O^1,l�8��MY�L��%�E3XC!�>x��Z��l�8a��
1!򤑸E|�
S@Ԥ}S�����+!�$�41q�����'��"'��:(!�T
�h��5�ݠ`|
u
dn�!�D�5 P��u���p��xx1�)~!��&iw�h1�	q2@7χZv!򄃍Lw0�+Ӄ�-u�EYu���Xh!�dV�D"p��@�A�qmb'îv�!�=n��y9â`H1��e
�N!򤛅b~�D��^� C�\8a�?�!򤆡U���SB̖3~��@�"Q-!�=�" �U�V�l�i�M�0�!������2�ʙ^������E�z!��	%�ꄙALP� ��њ ʓ�}!��䰣�g�x� @�+�T���4a����h�ts༡Rj��y��)\�=
�$��5��R�GR6�y �i��M�5�͌w5H0���3�y�e�!*�4���ln~%9R

;�y�N۲Z[�Y���ݻdW�a ��^�y�F�H�N|�ƈ3r��H�a���y�b 
^�b�1�B�8s�l�>�y"����R�g���[�H��y��?h~��qcbC<q�pリM��yb쒟x2���"V�pr�q0E'�y��J���@��*9��js��yB
D�KZS�+���H[Fk ��y��ݤZL��8c��xMY����y�k��m68��w��"��t�ĭ�y҅ֺ��� D L�=
�!��y2N�"g�j|�ҏ���yK�%�-�y�[>/m��:b ݳ�t 6�V��y��D��cweF9<�Ed�y���2'b�c�	���k�����y�`Y�Aʬ�Do���bB���y"SiI�
4��Ӈ�H%�!����ꘊu�ʪ�����DI�G�!�DĥK_Z��0F�f����W��U!�dL`u�]���y�h蒢TE!��	�:�V,�GK�VO��٣�B�^!�� �lۢ��z����E<Y!�D;{3*�3�C�$�ؼ�DŮL!���wO`eSE��36�����n/!�B�/��f�Y�I^ ���W�!���
4�X��a��$��/�!�$��"��#�e��J"�,�$C�k�!�G�N��dB��T�0n�R .�!�d�aU|Q
��'�V���F�'�!�d��|G�tj��]y�t��3��	4�!��� �<Q���Bj�}��8�!�D�"|
m�!׾dJ�mBV�5F!�׻0�S�Ï#4=D-���Ն�!��)G �H6�Սm;��A �Z�!򤑿&�H�Qm��W"%�/
p<!�D��Y��i!0��+C����#m��e"!��&R\+��ҁ��Tے���!򄉠=[��0���%R�i���R�nl!��L�=���B��T�O�}�剈p�!�� �a�ǓXİ��9*V�4@s"O�񸤋C yu��9���3=ʘ��"O�=1���)����w�.~2!��"O��gA�L�"fS�85�Q"O��ѩ]d�x���V6(F)�"O!t'�m���!w�U.$*Ҍ��"OH���"X*H�.߿�Z"O�b���@T���F��%�5c"O��v�ڶ �ǎ�w"D1k�"OP|9�,]*Z�1A�|
��Jq"O����k�>����Րj!�"O�`ԍS�8�D�2�׹k���B�"O��¦L�������-�*m�c"OHݠP	�	d((������"R"Op��ܙn0��t��p��:A"O��C�ڿ_��8��[�ł"O��QNA�p��	A��(P&��C"O���nYD�,��n]>��p�"O0�����(��1��T��(c�"O
5��戶q�x��D�h��c"O��b����`.2�JSe�#V��a�"O����Z�T���*�7V,�z%"OuQ�+ߐk��x�W�3�ެ1�"O��r��_-3�t��D�I��0�"O�� Q��=&���v��
`�Ȓ"O>u8TmQ�<��TQHX�PE4٪�"O��
��[ch��X{5�D��"O�ظ�� ΂�i�&�q��h�"O�i�Ɨ��d�[��*		N��V"O��āɢ[?�$
�E��ʰ�@"OBD��D�`�m��3*��h�"O��;�ɪ~n\��FI���á"OV�`'���`�M4�T��A"O~Y����2�z��T%E4V���"O x�d�N�nizx ׍Q��v ��"Oޕ���I��r$�?����"O�q�FȄ�Wjδ�KG/k�~�7"O~i�s�޽b�4�K��ǎ��Á"O�`4OC�J��*'��<2����"O��F��Sp���ֵL�l)�"O�$� Թb��t����#Z2� P"Ol��L!N��U�6m
7<1�E�"Ot� �m߇FTç�š|L�x�"O�Y�S,ʨYz��+[pƘڣ"O�|b�G��x�����JG>hg���@"O
��6/�=E����I��O_�E�"O��AS�� 8����5,��A	"OX���L\x��B�*ns "O0��Ӊw������ =h�us%"O�mX�,��1-^�.J�=i�"Obh���ݰ�f��!�@��4"O&H��c/��T��	ċF��$P&"Oh���`Vt�2A0G�לV�
��"O�'/�g,\�{-�7{�E��"O2���@66~$a؆ʒrx:ܙ�"O�xs��V���%FҞ$��"OlŒ`�ҹpÆ�Z���}���I�"OB��Ř dZ�����
�"Uk0"O��jGY;6|rl�#]�%h6�"O��2�D6GA�A�a�)V�ap�"O jv�ѯ�~�0�Ɋ?1ԹZ�"O$ʧ�I#u��e��­uŨ}�"O��U%�V�@����M ,hd"O���3�ԃ���B���Wj��"O� ^��«�/�"�0�"
�2j���"O2���D�~0�щ����SUB�*�"O��`�*T�o\�kF�ʠHz�8�"O� "���|��!9$ѩ7"OV:GC�������.E'Q,�AH�"O��CHĔ5���ӲMKu�� �"OvA�m� S��*EL���R��"Ox%Z`��(l�%J1�^5�Z]�U"O���T+RY����'M�6�n<:b"O(`*@�Ɉ~,��z�낮�.�`7"O���N���y2WB 9���"O�}��ih2��srͶ�v��w"OK��\ ���5�ҭz���0"O�	�F�Q( m���	
:YzP"O
}�d��M����o3P)a"O~�c��=�ҁڅ"C�::�Х"O�9# &ɭP��0���F��VT�"O~tr���!e�0��-;��M�c"OH�3�珨{)J����ڌ���"O(��Q���1Gf�k�b�J�B=��"O�1�N����ɪ�a1*�X
�"O�@C�X�Z}���7�p����S"O�BwM�<��ui@��d��A�"O�I��Y$��yjsB��X�"O(q/�20��ܷ V���"O$�a"I�z��7��o	tD�s"O�d���� 	�T�� _���"Oč�@!�!���p!��vudpsC"O|p��ژP��ݛr�Qf��"O�h���+���"^f�H�jt"O��*�
s�@�ړ��*����"O�}0w��	��50KҚs�"O$���F��Eh�G*��]�����"O�L���R�HҲ�����u�dt`w"O�H��fʙ`���t�Щ
%��#t"O��S�� ĺ}�1��O�tQK!"O�A�nK�@�0�lڐ`, �r"O�4� NOA	H5ag���J]��Pd"O����F�M��a�� �N��Z�@�OZ4��"	�)`
�`�:$Z6�H�'�:��)��^�n����6#ߠ�	�'/�I2Œw� OP�O&���'f��!��5�5@���S��Q��'j��I�e_�VW��@FA]��|�<�&�<Zv5AAV$�l4)��o�<9�՜w�4�C��:!����oBh�<�d:�`���,:2�����&�_�<��J�?�L\:�e<���(�W�<���YT�YZJ9{��@� �T�<Q�hX�x�4��f�0q\��x'�R�<�ޅR/ބX4��/Rn�S�aQ�<	3�(?���"R �xd�x�<9B��?9ha�v���̭��'�u�<D�����3��N	�$�Q�L�w�<Y3*H(F�p3��R�R��mq"�Mq�<)�'��w� �(�ܿ!��T����o�<A-[�9/<	��T��H��*�i�<�͟:*qbH"��֌p��7��f�<��Ƈ�U��t��˿7o�����a�<��
2��$
�N�>r.Z�3O�a�<)EF� "��b��	�R���eZV�<�p�E)+H���WC7��i��H�<�%@�?�Je���2 ��a�FC�<Y0�Y6눥�V�C���0��u�<� ��iw
49rPX� c
	')8ɨ�"O�A
sE�n�̼�c�z�5Y�"Op�����(h2��T�Qa�d����'��O��b��O�U��do��7����"O��+�F���A��Z)<8�"OF�FfK�:�Q�dD�yg��(�"O��CJ*ʰ)�7!�2yP<@
�"Oz��AI �Fq��O��h�q@T"O��C
2%���WNW>���"O|��עS:>Yl���bY@Q�!�"O�v��6)���w��6,e��CF"O�i�F�{n�PX5&6+n�2e"O�ي�K�(%ܸ㥙��B"O���5
يX2zp�vgWc�*��"O�X���	Wh�c�睛{G�`[5"O^�#�6����D�%�L�"OL�HT�l�X�e��B��H���!�S�'~� Ыc��!b�y��	�,a�]�ȓ �	{���6(����)[�����Jq�[��@�"�D�2ptl�d"O�\`��:��5Aǣ��HDN<!�"ORk�,΢1ݢ� %Z�j����"O�L� �K�zڄ���˞.ݶ��"O� `��\|�4 �"�)���`�	p�O0bl{"�,XȜ8+�0,����'�����ҫ\��]�GM�!���3�'j���̋D-Q)'�ۙ(�$+�'��
D��!c�:3�� [���'�ZH���sh��qV
�!�'ܰi�!"Y�:�9�"�����!�'kv8��E�S[�%�ٜ0G<`�y�R��D�T�'��}��`��0�`.#�iZ�'4�0��,	���.�(w��8�'W�Ř�L��v6�x���7L��'m�$�S[FʘAu�1,���
�'��!�&�
G� =�͂#QB��	�'���92�W'�0�+��Q>M���	�'>���p�K�0��F%�1?�XHÓ�hO�9+Љ��S����v�ކ.g���y�G$@:�a���	(L�@�-K>�y��]!n5���A�%�֡�s�
��y�B�:M^��դZ ;������y�GۻQ�x #�*�Rh���ٞ�y��ϷD 82��4Y���դ��y�YS�z]q�eH�1��,��Ɯ��yr��9�4�"P�`�́���y��'m�l���Sd*���2�y����LQ2��C���Ӷ]��y��)Eʁ
'F����1FN��yΉ�<�$=�F��zm	ꆜ�yB� �;`֝��@��
�<�k �M��yr�r�6̒�G[��)�W���0=�����|OLp�g	��;Q����Ǆ����ȓH,��G^Di@�"K�N	�ȓ �R� ᎒�?K����U�'U����E�h}8�"˖s~8d�v��
 ݆ȓy��qc�A,� �D����ȓR��	�	NH�k��Pm�ʓl�� �+��\䪔(cC�ɵ �vxk�-��`A���'�E�B��$_��uR� g` sAD%'AnB�;\b��q��;WP@��[�t�4B�ɾ9�k� �B,J���Z�0B�	p6��C� ����J"^_�C�)� j��V
�Z͞i��% #a�rP"OX�K�G�B��A��Ip�j��� G{��I�+�p��)��f3���q��[�!��% �(I���ɔ"���i�H�!�0�dm���m���w�D#�!�$F-M����a��	^�*��\�!�̣��H׻zR~%�ӯ�"�!��2fd�P��:?5�ɊG�
�!�=t���h�fŭ�����k���!�$�!��e��dN/k�d�!�*r!�d�: �tܹ��G����2��8lq!�D�>G���	^�4`$&I1f!��b�(:�&P�$��dR;�!���$U��w G:4���1&Cƕa�!�$B�|���)v,D1p��<����45!�DO�y�")ʆ�V�<�M�.��S	!��U� ��ta�9"�B ��P�!���8N*�؂U����\���E-b!�T)��R�q�" 1@*� 6!��
�(+�`p�6,A
/�!��1`��Pˏ�od�Ql�"}�!�$��*|8p���ӷ90y�3� )2[!��T����' </��b��&cC!򄏚gw������u�1Ӯ��R!��}��5�SR�-�N �B��!�˜A&x��!5A�J!0g�P�!�D=l�b%b���.f���Ӥ�!i�!���D�; "��Rs�,�P��\�1O�=�|җ�^�-�wC��|+p�a֫�e�<�GF*��(T��N뢜b��v�<A�l'���b��[�DL�V��X�<9`�+��yȳ"��t`��Q�<����u^RTJ�S��p�&JL�<�A!C�I�,�۔.�=�)x� 
E�<ْ���q ��i��9I$���΍K�<�D�mJ ��ڱbO�����A�<�'bO
m�th��O�V�0YZQ̝|�<i���=��YD��)W���q�Oo�<Ad��<o��t�vf�(W�^���LR�<��.��`.����6;*ɩ��LX�<��Y�A��)"DT�L�3�bYI�<�4/I���:#�^�c�����F�<�g䆙d���M�O�iRm
E�<������8ʐ�T�7�������z�<	f��|��P���в,���+G�@v�<�D	O~,�=�bL7CX�{`��z�<�c��a�v=�s̓����a�����1��� �L��7/*��E̔2�DA��O���xt�]�f�V)�e�OR�$a��Q�<b��(+���x$�W�H��������d9;#�]��Ĝ�p|�̈́�k�Ea�Jí@�8�x�l�K��9��J$̠'��m��`U�),6D��K�|#� 7Ӥ!B H�&k�n`��W&m
�-����)���0��tt^�ktB� ��q�m��2�����,�j�':5w�X�𢄸/*���ȓI]�-X��RaQ�0!�Äe�<�ȓ!��M�R��+9�n1����uک��+
X@�a��% ĠjB���_}D\��)� �s�Mr�t��r��y�ȓ�,��w
T�7 �=�G�Ł|~А��'j�\8�!-`N� ���1�ȄȓR��	+�LC�up���!��.u��=��S�? h�s_�6�Ss*p�8�&"O04���Z�V1iQ% ���f"O�|���m�~�:��V�/��"O�Xf:y����ުhj&$�d"O\�_� Oj|*p�B�JI�H�u"O����M~‴Z�m��T3(��"OD�����y"T���ݮeD\�F"ON@�I�8a�E[����e֙#�"OT�Ӆ<%���A&ɯ"�V���"O�!�`т��W+e� i�A"OhI�N.�ƴ���[:7>����"OZh��oƈKKȹ��͂�O"�ئ"O`�r�M�>�.U��M>;B��p"O8��ٕ=T A�덃[�x��"O�uq�� Y��g�՜kR�{�"O��ˏ/�f���^2Bx��2"Op,y�&X;wm�dأ�ӵb5(�p"ON�ae�A�)Xb.�;2��xB"O�1��&W�@
`غ6MʹJ3R8�5"Oj�y�Oܵ7K� ���)t$,;6"O�9a�`�� ���A§/jJy�"O��Y�`�1U �8�[,tf ��"O���C�� VRV���ݭL�u�q"OR,�����'^��� �DFhK�"Ob,�Q�Q�*Lt�����oA��i"O`�
q��.��$`0,��6,����"O:9��5m���b��*s"�i�p"O$�h���t�@�15��؊��ɌH�<)fZ12O��ٜ� v˕{�<!��s��<ڐ	KyM��6G�\�<��^�z��딦�W
��&��M�<Q ��g�Ɲ'�Y�HG:d�� �^�<q��*����"�Ո(�h��1,�B�<�m� �$ ���ؘy�P�x�<iE�!-2��5mކd��Y��u�<�Wʂ-k�x4F�*T��!d��U�<����7-�d�%�7�Z���h�{�<ѕ.հP��Y�"�2Cz��y���p�<1�$�#kp����B�r����1/Km�<I䥌���؇������Zi�<1��^�N�ӥE]�Tp(���b�<��	��U	4*�;���"#B�B�I��yt LgS&%�F�ϣwC�9s�~�2�$�A��H���-n%�B�I4�ހ���ˁ5T�.ʤ2�g+D�|H1�*V�087�R7dd��C$!$D�La��ѹT9>HY�ƒ/?�z|�g�-D�lB��ZsB�q�q�Ե`����C,D���aJB	� �5��/y�����)D�܊������ $�F�<t�0�%D���W�k@@K׍��-:�S��#D��W��*(�������L���J<D�����#&����c/
�z��
�:D�������Y�\��a�L(�䬹@�6D��F�׌Z6%��P>x @6D���dEҷ{��]dꎧ(�qy��0D����T_�ZsN �1��uyBn2D��(W��/I0��S ۾eb��,0D�����G�_�]9Q���ypz�xsC D����l��$��Y��V�EmA�@c!D���aN�$\�|��e�{��d�F?D�4��^�	Dx@H��]�Su��iP#1D�8�t%�$� �(��QM�\CG0D����π�P�d1��I�1�@���-D�� ��%Սu����Ƒ`��t�E"O�@���J,�t�B�Ǎy]��5"OXE��N�>xn]s៍?4xaa"O\]R�
�>.!ۖΜ�eČ�kG"O(�1G��$�gKu���"O|xG蔧Z�n� ���
�p���"OR$�G�ū7f"%�T��;᪩��"O�MX��NV�2�ad�s�tur"Oh}���ܶ7r�1BL�>���;g"O9x��B�$:� ���r��k�"O�hㄈ�1[��b�:��!C�.D�l��ëm0���'C#F�U��'D�@�t כw�(�y4�ߕs ��@�a'D�4R�-M����H�2�N e3D�(���TCp�l���e>ڈP�g/D�0��,+K��ب�A��ظ��%;D�����<QT[��V�~�~�0 +D���֬X3*���ٍ�����'D��� �b�ָ���v��3d:D��9���;K}0Ёi�7�p���$D��CBF�a<HA��ʉ=�JL�V�/D��(�kD�eZƨ�)[Z��)ɷd/D���J�o(�2G-�pZ�Q��b"D���V$�H�r�x��W�w} @! D��J��U�H����A 
&|�`t�<D�8P���5nܲ�#�	V9p�8R�%D�t#c��v�D�C�X�L�Ft��1D��xp�C�u�
&���z$�5N0D��k5 Nn:�
�-¼|��d��";D��b�B�%3��B����h:D�,�Q
ȃA	l�`;v�@�Y��2D�H����*�̅��d�5
8>L�s
2D��x�BۄMB��1#$�'q��:�;D����V�{�D�a��F�H=Ȱ�We8D�$�m93`|Y
�ĲJ�JI��.3D���àЃ}�f:�� 2�|i�A�+D��
����4%�����<��v�7D��	�Y�E%,̈f�[�	BLр7D��!]T�$@�A�Fs B1�!D���G+A�Ҭ�5��X��Y���>D�����/Z�yz�k�0x��Y�G7D��x#̉N�Ʃ�r�8Z�Qs�5D�D�'(��u�"��r]Z �1D�@��к� ,x�!�0�X#/0D�0��͇�w�Je��&ϕ �.X[��.D�xs�%�t��$j�n
&<[f�'D�� ���.� 	B[����2D�����­19����ވ�{D�<D�|EĄ�RJ0���Q��E�J<D�h� f���ËP��v��d-D�$k�ϔ�h2<"�C�.��ph�`*D�ԫ�����٭EV�乆a];!|&B䉼�n��*b�´2FA	)B�2v6▋N�T�@���Bv�C䉹;��첣є{"�zF��=,�C�I�`�N���ײ,2�����	Y]�B䉁61F@h�Xn)����-5�C䉷BHJ�x�Bq%�(�E�&2�C�Is���JVN��"����3�_��C��bg�*���e��a�&����C䉪rBС�ꕄ	�14a��9+�C�	T���q��͊�P�ğ;X�C�	;$��P��+
m`Q��G�JjDB�	���$�
W R�ѳ3��y��C�)� ���G�P��F��[֢��F"O(K�V A�T���d�N�PS"O�dz�V���T���"OvasѤ**���D��.�����'�p���LP�u�dY*��It�^ ��'��y��ϔz��-�eŐ�g����'<̠���6�,U����^z.qz�'�p�"w!:k5ۤ��R7����''*�9�D�*I*z���?_�X���'
@�3s��Q5���#�D.B�B�@�'��P��s���3�V�?��C�'y���Ľ
�^���퇬z�8���'B|����u �Q���$hج���'h��0	�O�X�:!��W%�`�'A�H;�#s(��!qhJ=8H���'��Ḷ/ǓY0�Y�aB�9.)&�)�'��r¬�~��Ӑ�$-��Y�'|�(8Jԫs㺀ÅD��i%��'�p|�#�8.k���J�1g��!
�'90��FO��e��	5���e�5	�'�D���I�;�����¬Tm�`0�'r%"EJD�9� �Ѕ�҆O�\���'J�c��>^ܠ����#T=��' ��9�d�0/z���\��@��'���s�	#/x]:�N9FR`�'�t}x���lݰqs�nJy2�0�'��yS �=������ϋo�N��'Q�,ZҤ�"��t�W4Tv 8B�'�u���Y�~X|[��$}T� �'w� �I
C���^�Ajz���'� ��W��F�J]�q��$:u���'�~�x���05���B��H ��'�Y�儽B�@��Q�O�ˈp��'�D�����E�m��j�@�u��'a�M���G Kap� �枾
	����'T"�W��&s��!:��� _E��'����EѡU�t�Q�M%x4��
�'��7��'��Ya�8i(D���'���RʇNp*���#Ү\Jx���'O|�p3��Kc�;��Ȣ BF0I	�'��=�O�P%��8�!J7H��A��'�`�
1p��CkJ&R��'����G1B���Òi�P��	�'㸨��Zx�8ly�	C$FvBZ
�'�=�aCڬ�P��e�NDSX)i	�'������*�� �T'86�d���'�l%*��@�aR�V2��!#�'��+���/���抛C���'��)���{8Vp����qn�J�'H�H�
�8Q�� Fǉ�R���'Ȗ�
��\W�֍;�E?j�èO����3Q2�Q0���ZhD�Rq@��}`!�L� e�ϛ�
�t��4��SF!�dI'#�])d	E�:��H�O�K%!�d'��	`O�$n�`��$z�!��>���I�iX�1���].%�!��_	�HCq��r��Qx�
]�Z�!�9[��B'�u�����h./r!�DΖ>7&���*���[Fg]�!Y!�D�&f������4y (!q��Py�B�r��3��|,�js�ӌ�y"kΊN���r�-�mH���ŀ��y�ҷbX�v(͒<��Xg���yB �h��/lV�:�CS2zx,j��� $�*�m�7:���@Jޫ[¨l��"O��(W�T�N�EH7£1��Ԑ�"O|�&�˺Q���"/��p@�y+q"O�8c&�D�O F��/U�~$�U�"O���rgY�m����r	��z���"O<�)B��-�^6Ä�?��|A��&D�H���LNE���E>q��&$D���Ћ�����/c�M�.D�L��fX��+�W$r��1dJ0D�� ���0�TE��b6lY�k,D�X���U&(Q ��΁��C�(D�,�����j�Χ��Q�e":D��k�K[��D��
�rn�]���7D�dh��,P����
�1�����)D�X�aFLH\�N���t���b'D���B��~���#�=j�(9D���� n�ݲW��)P^�` M8D�T'�{�i�@��0yt�I��1D�LC'-�8B-\���EF.*4e+=D�trǦ��o"غЪ	~Q�L4�/D��
��B�g�!��랽|`�Lp�..D�D��Ő�.�~}���X������!D�����5��.���%q0�*D���! D<3<��@S}:��r��4D��j5�x�lH��HƓP��%��4D�\qg����x��E�G.ޜ�R�-D���0 �m_x8����".��@� ��mZ+	\,�zQ��t6�9q�_�+I2��hOQ>�'�ѻ)B���ʀ aN��[�D.D�h2���|]���+^/5@bh�/.D�tL	/���:U�Ȟ4H,Ԃ/D���5-A)](~ :���"+��:D�P�&��#?��di@�\�F���8D�4�j�>�X��pM*yQրsU�8D��"`GI�$�9��	6A�,x��v�,�°>yW(�9V�ZM��m_:U"܌�7�
i�'e�D&��5)n0zEoX-6�xAHB�R��C�ɋ5���H�4sl5` OQ�f��C䉓rCn��1,I4A6��#7#�\��B�>>����%�;R�d�6��d����<����@Y�0���~�2h���TP�<Y���# �|��1eX�#k�"ݨ�O4�r����d0Hu˅�R@���(�a}^C��DI$���L:NrR���ÙB�	˘œ�F؆)����e��p���'ћ��+�	�?)%?���'@ fȔs�_�m"ȡ��:4���х�"�byHt�Tj8���\�鑞b>-��)s܄���J��%Ҭ$벬'D�R2�E#��*#@ܑU�x��e;���<i@�H+Q9������q���PBUu�<��`A�[��( P�U.X%���\��8�OԁBg�7|ABW���ҵ#S��3O��I��� �I	.�Ha��RA�B�I9 F�i��%=Q�a�򂑷�xb��͓��<�7��"|�q���;OzR��C�Br؞<$� �a3@bpz#(�8��٩0�Q��G��æ��J�!	Pj@aD
�y"�ΓED��$mS��*��[��yr._�w���ҷh�����ľ��'ўb>���g�> �B�iDmX�[�¯&?�
�6Lʩj��B:c��]pf'c�`����~R�'���"������-\,n���	�'4$T�i�M1�e)Wl��l�<0�'8Ɋw���N�+�ϖ�8	�xk��� Ɓ��+� zT�sG'"%q�]Z��	Z8��*s*�meVa�r�M=
:��,�lZ4'\��I֒4��)t�Y�aB��X@�'�򏊃i,`��f8a���6��:�p<��}��':�J��V|a���m �1��'V�x�h�2Kt|uo��Pl�d@�yB1�S�'~��1SB̟&l�)�!ۙ!(�Ezb�~�Ub�$#eNx��y��B�Ām�<���<��B@it�s��Ch�<�3��g��DT�tL�i�  �d�<Q��ÅI�ڈ��-EL����Wy�<�4�F0Z�A�-L���YM�v�<I�"^�P� �pQA��Q����s~ҤBʦ}���d�)§)�6l��h�ڕ�F s�y�Ol�=����ɧw��q�LŦYs�h�`Ppbql�n}a �?�t�3�ɿF&�QS��.*(%z�̀E�D㞰CFV�G{Zw�$�qd��(��!�JͤR(��'Na�f�<�ͲUl����%*����<�!���+���b��WE5v!�P��4p̓d@LX��q�K�_-&�$�bߓ%��88��]�.�hJv�ɷpI��z���D��=yd��2�2�6"O�����M�p!@�H� ����Y�HGz�\?a�	kyR�"�q�;�F@AW뗫4�c�H��I�f$Z��Q��4[��4��I4h���z�'��D�'=�>�Q�� �D�1��_.���	ß��'���П
���@�֫	BQXiH�F�o��x�<��On�y*()a�4k��1I�Aqu�|��)�S�Q��J��I+R��`�B��?�6��O��'���<��B� �A�.@j8��* N�&�\����uן|�&��Kgo�$�"iP�����4�O��#��>	5@iN&i���2�'Q�w��Ⱥ���W��sDJ( �hԄ�	w�'^jXx +V��v�ah[5,��')����!X�0�<�� 3�Q��d!��#� �X����X��H2�%`?D���e��v� 33'��a�d}�6F<�d;�Q�O+^ ��AR;6��):tIA�=k��'����b�^�^�p�V��0�4���/4ў"~Җ'�����(	�'u�N�KTNOD��$�l�'���Y1 ���8���|�.X��'KЙ�/n����f^�w�=��g�>��M�@� :��#�Ņ9E���3��Lm�<�ag�'&�=Za4עjc%S�<�q��.J��r�/`�.=��MDh<ٰ��Z����D��6)-�������x��'�8����\:H{iq�Y*#V��Ó��'wk�>��AH�iĈ}�����̃���'��z�:u�n�k�P!��Κ���d8��|����,RW�?|_�PK'�N�`f س��!�?ً��> \�0嫁�@_��B��I�L �YFx��)�S��T���bg��Up�,�a�G�<!$+BR���<	�ԡ����E}��'A���6��h���).Ѿ�z���xL�\�+ @p4Q� ĕ�'���ȓIq4!��K;9![�mY�L��̆�	��x�c��	!��gJF5Sy"��ȓ��1f�ǩ3*B�2�@�ej��<!�4�0=i�nG3xG���W,Q���J@	�nh<qP�O}f�z�
O
K[̑۔ ���MS��'-���ayJ~"˟��$�U���F�H,Jeb� d.��=�N>��4W��fA�y�֥1@�J.ad���p?Aqk̶t� =�����F����HE��hO�l�*O�	�E�
����W�q�fI"O� ���ɘ"4�]6�ʈ��5�3�|�'����~�'LF�2u,R>\��8�A��'jLU�pGS�Y�Pa%G��E����0�q�hiش�~��Itܧ8�L\� �296����#S_�݅���1�'*`�XR�Ô�<�8��^�,qv]Y��;,Oh�bsiPO7LM��iR�i���w�OTU�u���L�Iץ�$�y�
�'M�  �38�����l�&�b�}��)�	
�� m^6r֦���g�!�r&�EA0%�Ns�X�k�^!�ܝW\�X��ߎ�`5�iũl!�D$5�b'��M�������)Y!��j�22��tyd� w�N66�!�ā/
R��שoo���V+��!��X�*�
aC�ۼ^ �c5�Ġ?�!�dG�<�v$Z�`�
+HΑ��*��_e!��M30M��*�F���M�G!�DT��`��AP
��]��E	�!��3{�ʜ*DC�o�J��c�$t!�d��j�T�c2D��w����VB�6{!�$ȯz���	u�[�a�z� �Av|!�Dߔt�,bp���/��|3�CA\!�ٻiG�{����a��}R�N,&!�B�Y�� ��aG1QUP�P �+e!�dR	��q��5JAR�r��/!��A���1�]�c�)V��)�!�d֩h��,Q�T�:o�H`X; �!�	&~��%1E��bnp�q�)�G�!�d@��b �M�e}�(+W)K4c!�̤�b����P�,V�ur�ׅ'�!��>	i�8j=h���p�0��ȓx��.Rb��ӱ�� >��Ň��tLh��$�び>��D�ȓxgzd��c�|��0@�.~8�Єȓsx�0�)n��pHv��rnĘ�ȓ&���c��ji�e�@*�qJV���0��n�W��嘰f^�d} ̆ȓ=�%bE�O�P��-�f˕3f�t��ȓ:`nuJb��%2n�i�P��/�l��WX\b�N*Xc�=J�j�$ �j|�ȓ=LP��@,/��1/�8 `�ȓ2�.���T0��(	��֖#�`�ȓ,pl�q��Ȇ%��h!���&b�X�ȓK��b@͂ �^�QI� M�$��P�Z�z2MA�m�0H����W�L�ȓP�f�h����J:ؓ�#gr,���'�I�eK@���!,apP��P�,"�H�7��% З|��A���"u�UF�0<AD��M���ȓ��l{"%�.�"p�F��	;r��),4Dm�0_����=怸��7���q�P�SAJ�6��+P4ԇȓ-3��Cѓ(��H'���6]�ȓLN���J7mF\��V�+��ȓU� a�V*�a��V�G��&���\q�U��[�ew�M���ì�d0�ȓ&�(0{��\)xr2��	1��!�ȓ/�ڐ(�*��
Wt�)C�ȁ�^ ��@�b�c���S�3� �e0��1�x��g�*)8�R��7��I�ȓ	��d���L�#���jb�Ƀ<��H�ȓ���0U,��P6<���?K(VX��\Z��i�+G9.Ҳ��D� yT��`�Z���Ҽq�ɪ�fωr�Ї�S�? I�m��W��0�p��l'~,+�"O��+���! ��*�٩I�q t"O�]��(Űu�P1��J -\PI�"OXq�Ԁ�iҔ�H3Ή�U�1�7"O(-���Y��M[�lHӖ�aS�"O ��LA
XˆI� ��9*b"O�S恏��Ƞ�%;�]0@"O��G�0D�|�#�'�b��P��"O����mA�=`1Qe�D)R^ ec"O^(Y�+P�TJ ��CS�a�ܕ�p"O��I�`ٗg��d��M�-�D�V"O�@{��ߌ7�֤z6�S5�0ɒ"Opɰ�H�Xhp�T�K�#�b�a�"O��C�1m�$����[0)nLa�"O�Y���P�j�(ĢW%Z��cb"Ol4ɒ炙J!��v��U�@�"O���5OT�nT�w �w��`��"O�(��fjh0�$O].K��,�"O�1�#�	ۥ�>l2����"���y�JD�e�1�$���b�Ƀ�y"n�-�DYq�'T�f�H����y".[�J�r���B6�|`��E�=�yr
��ll�|P�d��W��y⪟3 U�����T��cw���y��N�]V�R�Z~��pƃ���yB��	[P��c�1Q�"�R6�]��y��J	����چz0���ٚ�y�	�\���q�%�-H1$���NK��ybUjX~� �K�1��A��)��y2��Z�ތ��ލ*(�cU���y�a�,$0�P�/o��|��ID��y�eP�~�����'g�	X�.��y��,p�DxK���+�:Q� KI��y�7G��@�@aж���{�����y�#�PA2���6J:@u�'����yb�ű2�@�C��y;���i��yrȌf���(�I
�m��8�a�y��� p�C�&:h���&�׿�y̜�=μJ%��?1����0�H�yRi3�t��Bg��*ؐ]z��H��y�J2�64�v�F&3�b�B��yBŐ� F�aSR( �2�x� C�y�gѱQ�tl��T�5Y��[���y2h��U�Jxj�fى%�na≏�y"��16�Vh����$��x�1��6�y�dؓoA��f��>"Q<���. �y(�= � ��ǎY�#�"�J�ң�yB��:	5��Hd�P�"���F��y⦒�}�&����6��8Y� ��y�fʟ)i�Im��y�RF¢�yR ֹ��<�N�=���e���yR��=z���c�F�qAG(���y����r�2ɪ��j��5Cv�,�y2�۲y�<(�ҷl%�j�jO��ybɜ� ��(�0%&p����TD �y�A0<,�8���U������yB�r�0u�@#Μw��KO�<q��͉+�\�AE"6eɖ��Ѝ���\�?�KS	��&��TXQ�JV؟D��O�l� "#�(7>m��*֏3c@9��g��ѨP嗊v2J�BO��3_l���u�R�X��ѴR_����Ny��ȓu�0U�A�/fXЀ�EY�qƙ��"u�y���J
a�(3@eE"l/���S�? ����_i���l�?nN�d@u"O�Q��G��d�>TS�kş0�L��"O~|�����jF
rx��"O慢��Rv ̄ FcV�5j,<0�"O�-Js$���"=چ��_Kbl�"O��'a�#pf�����+)�d��"O�p����jBd1�Wlw��"O���*̔!@�LYЈ�6<�9w"O$qమ=j��`�Ʈ02�ʷ"O�u˂�I2k0B�D��=�|Ze"O���M\ s�X{RHF/A"1{t"O� �Yk���R���@�*�"O��ˤD� #�h�!t��Ԛ���"O���¬V7!��d0��08�
@�*O�	k�(E1 p� ŮXk�y��'?L��``�l���I�ȅ���y�->H1ޑ ��h��ۄF8�y�FD�Ϯ}�2j�X�����y����Vu�]��k��Ti.1a���y�O��P�B�FL�x��,��y�mEVV�窀Qנu�ӥ��y��و@��Q��Ȑ>d��S����y��Ŗ{ Na�	��)6�)���y��H;b|�R�LO� j��Z�,9�'��B���,�h�Ydk ;-���A�'i�`%k
���8dR�+�4��'N�b��S�7쀄�RK#\�I��'���K�΂C& z�f٘2��h�'��� ��B	DOv��RiU@�FP�'m @�gn��aw4�aR�DaN�
�'{8�M�1X��NP�0Ț�	�'e�+sꚰC#:���K-|4���'M�C��M�U�Ę��Ϻ)/�5��'6
���%�1
����nV$b����'J��Շ#%}ps7(¥�*���'��ps�d���$���yL ,O���DA$;C��۵b�.B��A��$l!򤋀$O<RPL_�H\j��JL_!�$U�"�+U⃩F]pQM��HC!�dr�h��f����֩0',7�!�dA�#�`���^�> q��G�D�!�d��XAYe]�)8�MJ��S�O8!�d͍|���B�ͺ(0��b�
�!�_��>q�4 ��(.�t�m��^M!򤈊vDKS�}舝�,Qd�f�@�'Xi�V<X�4�P��4=�9y	�'���� >,t�Qs�Y�/C�8��'��k���2��]�r�T.�D��'X,� GT����ӥ-�#-���A�'.�p+�Q&L[�A2�i��(>{�'��U�W+ ���H�$닟oR�\�
�'��4�X�V`�[��<�{
�'���
	,~:�����1�����'�0��bK�T���i��Q$%厉2�'��-��.��z��(�p����x
�'EF���t��5K�*�� x�	�'"L�B���+
�����,*�4Y,OT���&0�4MÖ��|0t<Qq�O�*i!��uԘŚ��`�5��@�WJ!�dЦ����$V�0�!�〣4�!��]�V�FH�.u����v��c+!�ĝ1! �kAh���N�q�,>�!�D�}�-SA��k�.pqp�L�6W!򤄩C��d:���3}��9�I��D!�� 4 �U�D�}�h�˒O�FMB�"O\h�A"��D��f�5v ~�JU"O�}e�J���|���%u1�"�"OJT����*k2V��#�I-n�d�;"Oj|�@*�6p>���DȻ�iQ�"O8i���;�jM�g�_�-�Dh92"O ���ҤcN����V.R�\��"O�Xk �O�4zpPW-�<�ڴ8%"O<p
��O�D����I�O�mH"O���$�-�T���a�U>�,1u"Of�S��OsuyٲNG+8�I"O��2D��h�:9���T�|���S"O��Qba��ہ혉�@�c0"O
�"&"(KDtd��-P&nJ��1"O$b�L^�0	D�(ʚg�rHY�"O���F�-|��bTQ��'"ODI�b�ӿ���wD--
eq�"Ox��5+G�cF�)�p�Q�	�|�R�"O.�ySm�=7��=� �OG��ź�"O�1���[oՊu�vl�s_�P"O�@�a^��th�K˂>S�y!Q"OƜ���ڤ["1�U�K��"O��p���.I��%X�C[�v(d!0V"Ouh6�JH���(ʙ�e�""O6)�&  +^���K��C�*z�h��"OtKL'X�L�k��ӷmtY�7"O�����4Ѫ1iF%�
N�16"O�Q��a�f�`P����D���"O�A�OGcE�l��"ع[d�̓1"O<��@�80K�
�4qLj3�"O� ���9a��-"s	P*t'�E1"Or���@	o�4`�'ƚ�7%Bm�"Ov|���0�l��:X�ڣ"ON��B��>���	Z�.���3�"O�����=��h��3Z���)�"O�D��Mt�<��6���|�vp�$"O��ö��6�Kq�T�yߠ��"O&��0B֯Rm܍�`٬q$hH�r"O�Ŋ��۟YW� ��={��`�"O�]rg��h��g�.�(��G"O��Q�cS�H�|�Y����ݮ�H�"Oy`� s�ށB���{�ƭ�@"OfU���'v���
� Ŭ1�"O�X�!!�,����`jK�2��Y*�"O�E�ԡ_".apt�JQ�b��Hё"Oz�8��&:��x�;H���ȳ"O`�K�ʩD��B��L�:�z��5"O�H��ɞ�BEҳ%��m��s"O64����#x>�*�	|C �	�"O�j��Ѿ�x�	��5)54��t"Ov	�@D/��z�oEX4�)!"O�)��_�;��b!��*n����"OX:dJԝp䚘2�J�<@��bu"O�+��0m��(0�x, �YU"Oz��3�V�2{�ȕ'A��"O�h�u�U09
,�.�Qx�@)$4!��@$����2O���3"L�^!�D�������1�j�"uKL�+!�d��t:^�ygD��&�(A��*D+O�0W$�O���戆W��jB	Ȕo���w"O���A�	8����4���"Oe	WkU�ck`�26c�4x�r"O�%���51����ҩ|��@2�"O
��N�&"�m�� �R�"O� >�Vg�:R�JЉV���_�µ�f"O$L�F�ۭH0P�d&�Qtإ0"O0`���iE���E��ksJS�"O��x�E1d�,95�NH����v"O� �Mb'�P� O�Cn> :b"OP�9&]�.D8��0#&Iv"OX����3&�p�q�Tj�ۆ"OL�z��P@PҲ�\��9��"O쌈��M�3��j����Z�� `�"O�4��e*zX�AgP.��)c"O�8I"�\#B1�ubpg<��c�"O��Ç��mŚ@��H�]���C"O
��Fl��d�=(��AFI�b"O�0k�!B6�B�`���t Ip�"O�1����+f��6L,��q"Ot4+�1|+��c'M�^ ���"O��š�8*6$�dKE��"O��vOł{�JQ#$,���2Q"Oh8q�	��㶪̗o�jAF"Oh$pE�̈EfI	b�)���R"Ob �O	--�l��A��_�=
v"O�Y����G��q�+S��D=��"O�4��~h��#/��D��"O$i�g&��3�ٯ�.����gFP�<�e�$_�ܚ��E�*F��pM�<1��4hҁ���ň=����Ob�<�!R�[���M�7���³ͅ\�<ه��"��A��Ғm�.�[�<I�:wV@⡅\U����i�<qqd�l�\��X�&QcEi�<a���gU�4c4$ďǦd�4�O�<�#$x E�#|�jU
KJ�<��ƞ@�,eh"��*���X2hGb�<��h��KG:$��^.-v�4K�l�z�<!T^�A�Z�� U�<SS��w�<1�ٿ5Ep� �iS�Urt]��
�m�<��H�1)kH�k�m�5GH�� E�R�<�r��]r��r����l;7$Z`�<q$FT������-����`��`�<iB��s �\��K̩N�L��
�v�<��nk ������%&�Ђ��w<���Dv�A� �<)�� 9p���^���
3�Ql\��CR�����	X�'���AR;b��-�Bl��y��'}P�aP�V�!Nܣc/�Zyb��O@�=E�B���4�@6J���Cte���yRO��.P��3���^����LU���'��{BÊ^N��;��݉�b�*Ca
��y2o��oN�('��o����5$݌�y�)($�ft�+�U <� g��y���&-�@(���ܠ��N�y��$E�<�a�l m��Hh�nF��ybG�FAjL�4e���p�Ѹ�y2���s�`]b&�0Q��MqeC#�y�L���L@&�(hu�U�yrd�(18v�a��7J���A�:�y2��m�h@�vJHv�,l�AEQ �yr�ܿ_�rA�t�e��1�0-]��y�!�7/�Z$Ȁ�^#rp�NO��y�Ͼ_TA۴���Kf�#�AY
�yIټ@�� �֣�v!q`�L��yr�I�:*'�>!^�7l���p<��D��l1��I��1?5а�$�<X�!�D�+*]���S�m¢�bR���h!�� �y�7�m�i�����Ap"O�D�7"�J�ڐ-�
yz�v"O�4���C�s����Wˆ�rip�9�"O�e�Q%� h%�]�S�>xF"O������,�4}�$
��`�$!1�"O�H5�V�*��Y�)W=�|Q"O"���C�-�@�qEK'h���d"Of��c�D�*�(*��E�G*Ea�"O,�җFI&^61�.N�;> � "O�M�>�����	RK��c"O��
�b.4�!C�J�eV����"O�=�CgI�^n�M�ŀ�9z�hl	�"O���uθ*�ִ���B59��Aó"O�	��J
4����%K�8���r�"O�p�mݢ@8I��#���t"ODu���r�0���k�����"O&��QfD2�I�&)�1v42u"O��ɳ�D�� +�)�y�6���"O�����^�%�qG�������"O��hQΌ	����1,B�8��I��"O`��Q���^�ɈfB2} �
�"O�L���	<��@p�_@�Qx�"O�yҡ�ʦ;�He��7{hp�)"O�UC�jӓ,�$A�;""O
�x�(�w��M÷N�'pk�!��"OV����:*�T s�/@9LP����"O��o�u�
�"�J����"O0H�P�E����ٔ�я$E���"O�!x����x�BU����2��۷�'g0�A��O.)z��00�,	"�_�S���C�"OƁi��U;?& �R�Mv����	
=�ȝA��S ��`��L�h���@ �	�s�C�I� �N��c����6ࢲ��J�j�ҪU:��"~��h��[��"0f
��8hB�ɓ�>����%8���jA�4��I�e�6���'�P�iɓ�r�$ÚPҩ�	�l*l�jf����n�
`5��1�����$D�y�,֎|7�L�5퓘kMXza�'ʓ�vA�l6�2��E� dSq	?0��	��۞D9s��>'����J:}G�oZ)cH��?E�ܴ���\}�l%ϟ(U��S4Cr�<��Ax'���E��5  ���u�<a��ё=�~�;5�>�̂Q$Wq�<�c�F����f�5�R���s�<�c Bt��#�L+P��Wc�l�<a�K�/u2�̋�IJ$1��ccJHd�<��T�
�^�iB�4D��KG�Y�<0A��h�
�@f��;T�t՘�c�<��d=?�|��i����p�+U\�<a0�׉Q�"�YWI�#?���)�̖e�<A*��I���@L��2���R�e�'Oў�'D���c̔�kM`x�(_�Am�[b���b��s�X�B��	09\�!B8K�����j�����@�T��e!BAZ�- }��F��y�Iۖ#��P�B�G����d��`H��:%z�Yr��|��	/�h�!��46�%Q5e� 2���Céܒs#rP+!G0ZR�z��i8�'�<4Qb���P��p8�mI{��a�{��N
<���ʴɓq�:��W���t�4��RM,TH6�W5v`�O�7�:�S��3?8y��Ƈ,�0�w���>{���CS=jp��Bʣ�?�g9�gy��Hw�iQ�e�0+�E�צeGx��>y6��ɘ�R -	�WOb`����+g�jQ��l*؂0C���:X���d@%�������}����R��?��D<�����s��?��X�:vi֖ݔeД��B_�;6H�a�b���+�DD(<�l��#��7�@4�"햬?�'�D8�B�.5R����׻<�`�a��� <t�ԁ���U��jP,"�Daa"O`%�r!�?`P]�WI@F�8 ��(j�c��7{�ty����2���{��YVÎ h7�l�R�]"����;�аhL�,�XT��bC2 �p�"�M
5Ȱ��J�&";� ʇ�0<q��Ư/|��0�@�U�ի%�]Ux��(��Q����d\�"�~�"@�P�L�D�`�/�7�N��L����y?��K�B3"?��P�I��<%��H��	 � ��[:b#��c�Ḩ	��E� >��j1�^8mq��\C��.�#[��	!�ʇ�a�h퀥���6�x�e���a�z�f)VO����Ĕ<�����ʘ\J�Ds��>~��$׸D�ʵ�O�-K�*�f�ԄS$k��*򠰉b�@-gb&|�
-O�]��
�>2��`�a�0 ��Z��'�j��P��}Vt���&r��i��;��a�P�2|��Q�'/^6�x�l��"$���[0��l��Np���<��3Lv��3�̩+�J�uA�|̧�
I1q �R��3 i�yxjՅȓ]R|��V��3Ǆ�'RrE���E�o� �J�8qO�6m���(��ɟ1B�
!H��6�a��hB���D��Ĉ�I��A �GQ'4b�̹!/čnE������a|yR3�'�Lh ���@��{A��2�|a��`.�If@֮n����0"�\ϼ�ƕ�E,PsA�Q^�戅�)`!ӡb��s���6�2ml�Dx��T�Z�#EL��	�3H��3ST}���&J��y��"Ot�锐;�M�m�y�z!�Ʊiu"�R'[")�ɧ����e�s6&!�e�W�`�.L��L����0>!��J�$�D�[�d��r�*�b��E��T�1���+G %��L���&M�������밂K.b��LE�1F��"+�ʜX���q1�Q2¦G�U$�B�+�����M\;}�~!bW�Ⱦ&CC�2Y2���S(32*��J7\R�B�ɲ@_��7j؛%����I��d�zB�68�ɘ(C	��(���"5�jc��D{���aىg�D���U4��<뒫��y"hS�Q���d�Q���AbO��yb�Ѿ3& 1S�]%#���&���y�@V35`=*�6w����Q�S��yb��E�x��h�oP��Ѐ	���yB ��2���+�
@�\��Ѧeܘ�y���(��۴���g�Hm��A��yBoԨqEfDKoTN������y�j��Z����ߘy�b=  ���y"L�_Al��D�+k),��eG��y�蟝��	�e��2�&���fԴ�y��=
/*�PI�!h���%�G��y2�Ԋ�2삱a�$&� �����ybBH�{L��b�1nV�T rŧ�yb
 
�A�G+B�>�H҇H��y��@1ݼ%�!�!f�m�B��y�kN�=CE!P�B�@t �3.Q��y�iK
W��ai���V���*��y�)BE Q����
�A@�"�!��L� �V��t��<"���p��O�U�!��+$ ��BS�I�B�k����0�!��2
XF|�Ɔ˽Lt�Q!U��G�!�OO���@]4�d@���nh!�[0!�d#�(E8C'��2���h!�G�t��[���������LLm!��:B��ykH� cAN �jл"V!�� :�2���C�@G^�i#��e�!��
5.�X�� \�R��rt�&�!���FW�h����1�<���
b@!�ұrN)�u!A./2ƕB�Lҙ[!�d�>��p@쏝Z �9�k�/_!�DS	{�娓�.:��@�WW!�� ܹXg�3�JlHցȞHpQ�"O���(��M^a*C�B���"Oz�T�RP�, ��(S%}H�+�"O^�����h��3ըǌEd�"O�$�6��4jH��(C96�R�S"O���6�S?h��0H��C�A�"O��N�so���AQ�d�H��"O|�Rh��^PxR�G�.� ��"O9��g�l�P�s�ߠ7_�y��"Ob����}(4�@X�%f��b"ON��&�٪)ݓѠ8#�T��w"O��9eF8
��E���� s���"O��9��Ę��\�d��&V�%�v"Oݠ蓖	(ʬ�s�O�#���T"O<�j�J�vil�G�G0yL@B"O,,��D��C��S�Fت �V5*"O�{ �U(!n�M�d@t���xr"O�ubÛ;����Fm	* ��r2"O�l
�f�2*�xH��"_�H2�"O����\&8`�1�ƴ���#�"O���ɯ"i��@wȌ,A�^��"O�8$�� P�>]����5y���"O�1�v�[�ce�I*T���180��"O�X:d�N�,�����o)��A"O��`��" �t��*;��j"O$	��I������nR�r"Or	j�ڏ"���Sl͆[���J�"Oh�W��JYjl��l��X���"Oza�d�J������t� ��"OJD��? �Ľ�1�ΨN&A"O��PE�C�Pʌ���	���I��"O�M�f��PU��(�%�F���"O"`CF�+�.(BEL�8��"OB� �E��������KY� ���"OP�'.N���K�E,]�p�3"Ofu�aI(~;�-��,�+l���"O@	�$i�='�QA��[��L�"O�a�(��!A��T����ݲ�"O�t귎�:�ؕС�?6w<耔"O��[�C˭l^I�C�nN�1�"O���iv��1#�_�`qV"O�1kb打aɁ���\HƑж"O���Ꮴ^n-���_`Yq"O`u�FT��+�-U*aN���"On<Zq �	�Fd0#@7+	����"O�����%ua�`0\p樀��"O��t��GmB%�A�'s���"O|��bŇ�[�f����_�F��hJf"O��2g�3�izd
��
�"O�$#�Þ����aȅ�rZ�<�"O�L�
ψI�b}��hL�#{����"OM����Qb� �p��-�}��"O���L�Q�`����ɺC�t��"O�P�f� /~�21�/I$e�r�IT"O��i�%�##��pK�I���&"O6�CX3٤����@"8�&1ړ"O��g�\:b���a� ֛%~ڌ�b"O�y)&�کXd����w1�l�U"O���G�ՙQ�B�G�J%r�@�"O�����.|X����U�."02�"O�3s���zu�`C�����,ك"O� �Q��X�҆�/���"O����� �ze�A$��|�
�A�"O0Ġf�ߘ`XD�v&\�	���S"O� :��KJ@읲�S0�4ɓ�"O�x�UP?=��T���V�~i�"O~�:po�z�\�$��*�
�3"O��a�4.��P�\�n�ı��"O�YC���A�x��H �&�§"OnE`��S������n\d��"O�M��F�;��1)GCH%��|Z1"Od��@�B0��E��լ/s�9e"O x�ѭ��0�@�W�cf �}�!��F�R����ɽ�*�+F�	�[�!�Dݣ7:P$��e�;�|���&W|!�$��GL-IsN?����M


Y!��\ے����7~�H,VQ�AA!�Đ�t�\�$KW�$�v���HV�,�!��#Y��5��j���;F�:=0!�dH�/��Zg"����X0��, !�ĕP�z�0J�& ��<[C�	|�!�$V�ؘ�C&��AlС���7v!��¼_ �U�C �+LKL$5&�3[!�D�:<K�ڗ *jhʁ��_!�Dy�\��c!�vO��"��!!��]�p�Ź���/5,�n�
�L�!�$ӓ~�P�Awd��-(�{V��#�!��v��Ფ(�/L��YkC�ɻd5!�D�GG�‬�;5��A�BՇ1�!��2@�
��`�
u:�@�oSO�!�$�%쨽�$��4�f��v'MS}!�0f�L�JdE
7}D�s��E3I!�D�#��|�P�2���6�O�	�!���f��@��/�'p�e0O�bW!�$Y𼨢��_
P]�H�$X�~S!�d�=�<!�N�nS��Jbm��r3!���	xմ��G!��/A��Rp��!g�!�$76
��7'��L���	�{�!��MQB�bO�4k�����)�Q�!�Pjb&��ԡ�)`z�L⇝s�!�dJ�`P�c� �^0���@�ނf�!򄅼OJ%�1��HK(�[��!򄐃QR1c�M��I���++c!�䃔I������ �{���W.�X�!�d�v�T=���I�h�L]�{�!��0o�`�V��$2�e���d�!�D[:�\,#����='� 8�Ϗ��!��,o|楘�D�^�<�@F�	!}!�@�]e��f$s�H�Y�5R!��}�j��D�Ɉ~c�$k�C�)GO!�$�7��%�&lpȔ��3^"!�$�;�R5�%�
=t�l��-��`!�_�?k؝zo�3qv��$,�'g!�d��D9F�L8j��ԸTE�>!�ē�f��B�Łj"zP���$�!�dU)I�μp��ӞS%�I��dX#]�!�9L?�@@iC�O
�e%��w�!�Ӏ찶��a�ȼ�pŊ�0W!�N
&��I�I-,��0��&��(!���P�H"ʍ�n�dA#��<e!��M$p,�US� }֜�DV!�d�e[��Z�$�3?��!�c��AI!�ą.49�tȀ��XʀU�#
k�!��P�]ZT��ɜ ����EA�1!��3U<~ظ�G6�.0� Z'(!��N,Q�6#�Z ������P�!�d^�W8tp�JǓa�FL�Ӡ�:�!�$ʣM0���S9a�:��e�V yQ!�� 칚w�
kC:x���̡i��ő$"OX��5��5j���*��Y���"O6�R��4X.�l���/��tQ�"O��j'-�ik,d���&0��"OM���YE�Y�
)60"O ]����(W���HPk���"O��r�J'@���Y8!W�,�"O$��e9l����+@(q��"O|���8*π�Q4�؉JEkU"O�ذ��'(r���t�ܺE"OBPrw�U�ov$[�֟ �B�@"O>\u-^�Wv�02�p�A�u"OF��v�2GM��@��wk(H�"OT��bձ ���Q��B&K���3�"O�hj"Q.L�p��23���c"O�����R��&	Qr"MI�"O^�(0�Y�N��PI֙ Ö0�B"O� c�,�id��2� �^Y1D"Of��mt��+�� �l���"O�P-�2�h���%�Th�O=}=!��3X����Ϥ��w�	&t>!��n�<p�B�b�~���^)^/!�ɔ�Es1,P��xBc$x�!��:��x+�Ƃ5B��y��S�!�D.6�6��P�C**� q��E�!��?po���� JTT�3C� �!�$�- �<H#��w7@K���.}�!�d�DP0�`2�ߥ>'5�5K^9�!�Ϩ�<��`��$��H�EJ�*!�d��?,�2u�֍B��ū�霓O�!�d��ࡧ��z���vz�"OXx
�R�*��UӠ�P�o���e"O���уԷ6�p�b��N��B�"O|e���?t�0�������"O�Q��ăv�6���fZg�z���"OΘb%�X�Q��E�L��ʰ"O.�x�I�+ �`R%��4<��"O��Д�Ǿ>T�h��7oo�|��"Od�C"�1t �
���4uN��#2"O*�����\������ O�H;�"O��6Or�b}��O�Z����"OZT�D�?m����C@�ܜ(Y�"O��賤� #��3R������"O�H���Ք-��k��T�I��Ā�"O^��ȝ�.��D ��/u��Q��"O�������Z�f�P��©!Ѥ�;g"O�,�k���t�ôh�5a�C�"OR�� ȉP	�'I$ҀC"OFDI	 �1t=���ҹ����"O�C�mB8ٖu;K��4�>��T"O�,j2a\8��%K��M�|�"O�1�t�,|M
�7+߭K�5"�"O
Vc��c�Kź+(���"O�(�EN-!?z���βR�Cp"O�Xh���O������<j��r"O�Y��gے^G�ay�SS��@ "O"Q!H\�B50�F,~�(�q"Ox�@�*���I��べ �((B"O�l(��T:�B�N��P�f"O�(
��R����BΕe���6"O���@yv� �"�4Xp0"O�`;d,G+T殥[�������"O�%�5��G�] `�0�@��"OZ�AEJ�c��!@�ЍS�!��"O� N� ���4AaR����i�"O�]x�\l���Z1�)
��M�A"Ox8����v��x��/t�(�nF0l� ��I�^��X0�Ov�u��b���;R�U�U1%u�O��'T��O�G���)M�}s�$˨w�؁p�B 7��D�F��ا�'u?��p��A#B�n���g� d��%��p���R�S�'m]���UM/4̒��%B�8"� �'�z�i���S�l!�Eڳ�ћ j,4h&���b��7�7Hzt�""!&��Hi�ə�?u�Q���c2�PXçyu\����>��0(A��T��>��C�����'t�Z;��.cl��s�E��%�{�*�e�S��d���I} ��a�L��'�rL��� ���d�Y�e�6��wK�
LS�6����n�"
b꟦����.�P։��(� ���`��'G�p*�N�h� b՟F~��>I�џ���ħc$�0㵁#� z�'��~��'��I�(f�S�'$�$��S[0q�w灯)Ԗ`�'�p�����l�P���e���0`�6;⛖�U
a�O�?��'H�Wd�M��铣,�<�磚1i{�O~P��S;:A��+D�'�PŢ�"�6Uc�b��@�m�X�S�S��f�
ĎđRڌḡ+�-N�O��ac7�)��0-���[R,F�Zu��F�@����b0Ѣ����K&t%<P��Ý"yBd5ˠ�ثDc���ćJ��O�?�#�I	ۀ��ׄ���L�r��O��E����W���L�3�@Li�+����OX��0���PO\�'!���?E)P=L�X�Ł=gn}�U�>�%�xB�/�'hA"���$�A�2�(��P�<���=T������*>��$�VW�<����Lfu��N��"2��n�R�<���ڏ&�؄ӀÆ &Wv�����z�<Q�џh����4b��i�S��o�<�a*|�n!d�'}�<ȈPe�i�<y�j����P�މ3^}��� c�<���ЧO}Ƽ�g�w�v=�0�!T�4�����X&��`^�Ty0C�	��1��
�R������\���?J9,Ta@g�􉢗g�/k!�dY�r� ���菈V\�b �Nq[!�d�{��Q^%!P�S��ȓ<��T�ȓֲ�Bf����1sr�͒�d4�ȓaz^�'NLm��"��ӅVX����@A,0�v�ԐL����ь�8���ȓ2�i"���C�>p"�I�,s±����l+�n�}�AR�gJ>��d��g�ՠ���'s �ᓨ	����ȓm�����
X���q��(!`p�ȓ[
"��a%�u@�#&�� �~��YT�-�G�Ԧo��3į��``�Q�ȓ!�\�(�	\�fֈ#�� .���5G���F�M[)����B�e����el�P!Ȑ,d��]A(���ivD�G�ؠ+���4w;�x��	7:��@d�&V�����Ӳ-��|�ȓ+�P�C���$��0K+��d�2]�ȓD�x� �@�{�|M�Wϙ 0( }��?�U8�H�u
��2fY9;%�؅ȓ1 �ax�;H�T[ЁI������U�\Y�Q�E9S[%� � b�4��ȓ[��aP�,�S�͂gm��Y�u��0<M3#�!U�U���_���i�ȓ"�(�umK�zd{�dO�_��y��+תT ��TYj����G�0���	�v���/{7H%�"C�*Y$|�ȓq�mףi$��y6��+Bj\�!�"O� ~�'[ ~�-�!k�;Q��q�"O\� �mX&��+�)-HM��"O�*���( �ە)�	����a"OTtP3~�"RcJ�#&�N�@"Ol[$L�U�v)!@�J�)@"O�P��
�u>�0�ǣ]���"O�R�(�HI�GF�U�^8��"O�%2���E�j�Bc)�1,���3�"O��Y�o�!\؜��`��-l�Y
W"O�0��N���ၭZ7a��@$"O���ǖO�\|x � J�.	8�"Ox�0���g� Y�bӕ.����"O���BH$nzdM����*�����"O4��#ʐ	D�@]8@jʓ0ݢX2"O�ѡ�4D�6Hj�ꌍb��=��"Op����Z&�:��H�҉��"O��@ꓩ)�t�v _���H�v"O"�(7#�[R���� wD��2�"O����:D��( ��-25�"OjĨPC^qC*�㌀�`�D#W"OfX@�բS��@x�EMM t���';��5eW�"�8ex0E��
�'d�U"f�я(J^��g�9|�(�	�'N�$y�
*Jr �c.2�`���'��X�V�hd����g	7T�d���'ܸ:vh˜	q$d��� E����'�����ާ}�-@�oW�%����'���IU��� +r+��h��-��{��=�'!W�K����!e9.0������� �8� �RѪ�'V��]��C��+��ε&QD�u�
�,��؆ȓd9�1��_\li:'`R<����ȓ-���Rw�j�bn�4ڒx��3(t��*ܡH�R�0lHv�ȓF,
����q8!��ALLI�H����4	�'RK�]�b'ɿ|�\����zY����&vPl��(�� ��<��uN���7\/PFsu�:.� =�ȓD�}�Q)��e�)Q���0�ȓF�|����$�x�BQ-�h,V!�ȓ3<��R�@�j~�t�D�j�d�ȓ��h�E�ųk�a�ց[,+���0�H�IăV�6I��VfV08�t8��Z�B�Z`NQ?(Z*uk���K�r�ȓ�6h���Q�J���²�IP�Q��>70 ��EZV���<Q:�ȓY�����	��"кf*� "@ć�l������`=�xJc%B�Uu�\��!�ʹ`dA��U��=�Q ���ȓ|���S��w�l	
b������ȓJ�"\p�Aˎ-?npҶ�*��ȓ_b��8E`��j�Hi�R%�>4�Z�ȓz� �Z��U#�����$6~u$��-���rc.�8���W���z��F:�\i ����y��?j���ȓ_�R��B���2k�?,=x�� %D����ʝG��]�,�ԙ��'D�4�G�0k���2��B�"�M`�m"D���!G��.����1&���Bk!D��']3�x�¢/e��j2�>D��Pgˇ�>�np��$�92��*dj0D��ẅ	56�x�%��dM�`�q*.T��r��$�v�0��@*+�D��"Oĕ)ce�, ^�aB���E#��c""O� �0��O��[�#�� ���%"OdD��)B
�VL��o�o�X-a�"O��z�&ݚp��D�D��<I�nIk�"O��CGdҊ�b}XRmR6�4��"O�Pw��[ ����ѓ4"OZt�e�6M�%��,T�aYH��U"O\�!�ɫ&�2�j�A�o?�a"O��q1��>`+�	�	S&l |�;�"O���bH�'J�l�i���f�v�"O$p���ƥ+J
��6�D�;��]BE"O:�:1 V���v�Z�I�D`J!"O�D�,�4CX�S,�	sF����y2dU^�¥a.�M��(�@��yb�Bu� ��6�I+fTA���y��o`����쇓''V 0�\&�yR@ؾ����d�[�Ir�����y��	�O�઴O�#R
6\�"�P��yr(
3��%[c��Q��iQ�F�y�ό�hm�C�)Md�"�f_��y"=�V��a`�����Y��y��t�
ё��="�H��Ь��yrk�V��;�a��j2�e�gT�y"�0v}����ehd%�wLД�yBֽ,i���צ��[#����e�y��!���s#�¬^���&�"�y���-'��a J�'\�")�
�7�y�@�r�Z"�پ��!h�Ї�yb#��)� DФ���%fK�n���ȓG'tTA��_+7��kp�W�Nx�}��"���T.�=$�zx�qς�n�f�ȓT�����Ч0zEa�J	(vҖ0�ȓVU�D�W�~w���&V��d�ȓW�:dвG�z�Xpa�?=��D�ȓN�l��(��]fty�Nڻr����ȓ.Z� �C��}Z�=0A$ĭH@��ȓo<x�jK/��-H�Lɥ*0�ȓ yz����:��PbC�9�-��?��y��f��L�^�S�FJ�^ij܆�E�R8P���w�B�I5n��X�����A^�Pd�@�`6vȩ$V�`D Ԇ�U����Z9J�tH3��n#BԆ�P�1�Q��d�y�CaϽK��p��%�xK'��9lD�v�0N4���?�8@z����Z��m 0��iM�A�ȓs����%Iċ>������E�ȓxR�Q12�R�J��%����0*�h��*q��m�/>�����x���Xn¶�\�F��ܐ7])���q(�@�Lm,�����^'m���ȓ� ��'�9)s꼢WF�/����d	�H�f�x�d��d\.!X �ȓ���0��Z����"%��5�����r�T�r�F���ƪ'D��ȓ7��dhġմ��EȻz��@��gi�L�b�[0
�B�#��V�g��A���D�q���K�p���@6,o����m����f��[�|M��	1L�ʴ��T���{�) �@(@��R�&SU�A��C�i�����1�BD�kT�ȓ�b�Y�d[�B�
�a�R@:�Ն�|����կc!�x�p���!=~I��i�H)h��ܑK�4���Ŝ&�B��ȓ1�X$�a Έ��y�Ǣ�sgn��
5����`��0�
&�N�
# D�� 8\ӦF0\���Y��R.5��๠"O�a���G��H�w(�,q���D"O�q�2(��tf�T�������E"O\h����� к��5�4t���d"OX��%�M/5�����&\�]S"OF,@��D�6x	)`!��Pbm��"O�Qօ2IO.��ꋗ�4McC"O���� �1R�tɸ᫔�}�T�h�"O���a3��ؒk�" ���C "OVij���S���Gi�%QrX��"O��!Uǘ�7��{w�Z� �ps�"O�3C�3X���E�C�&��a�"O � I�5o�%p%D�O�|A�"O`����H vt�X�D5LI��B"O� `-)�\kVi�"F@$�W"O<�Ƣ6z;B��]#�|R"O���j	�$D8�M�¶�H5"O�����<|=�c��6��Y�"O ���K�/d(& � ����"O
AjWFÝ#'�1��/U7�t��`"O~��C.�:o�R|�����!8$"O������$-�2ܪǈ�6���"Ot��P���p�d�8
L��"O�H0��SHq���Sᙟ3�B}��"O��1��%��XC!�W�&d#�"O䍸�H��$��(�I�;Z���"O���T�|�ՁЅ�3c�I W"O q��ڐ�X���c�6
R%j3"Op�����F��(e��+�<��"O���@٬i�f���/L�1��ī"OR��E�
p��H�! ���ȓ"O`���ʱv�ؽ"��J
(����X}��'s��d�Č���/{fl*G�3 ���3���� �Q1�J:bU�r���!1������?��S �M���Uy�����Y�@�5y������.�b��g�����y	��y��~��� F���b�3��a����Oe����SMZ~���H'��D�Nq��Gr��O��d�O�6\�1cfY���k�r��En�qO���dR�doE����ۊ�ʴIW�a������u��4�����'��r����D�"�-x*0��C��u������?9���?1�����OL���)> �D+"��
W.�}E�G.(���L�7'^���6dSQ}�x�2k��6���
�I9$^4-�UkD�%�XrG�Fg
mC�)J#���s�m�'p�T�`s��/D�`�[3m@%���k͋UyRʹ�M�1 ߝ$�`}u��"K*��A�ń���7M�}�'��t��hJ&X�����G,��»K�'�a2��NC�AO?�����K���I!�M���i��ɍ0�lߴ�?��O���7�ǷdǜT���#@@X`p��ş��ˬV�<�����5��c�ǅJ�-� �֜��t�R�4��H`��oΣ<3���6�BH�5��	X>M9c�����%D'a��M�燇=��&Cײ�M�g剈y���Ěʦ�ȷ�?�`��t��#C�+W#�����?9�����h��I���S�`"����!ȵ��5�t��#�y���	
�Q���)ѭ](���E�4H
�U]� R �Mc���?�.���f��O87-�2��0[D
��k*�������E�I7f�:��@������FpU ����2|�|��R>A�;g_����e�>)�L�p5�S�Cl���'�.��W��Ԉ����!�U����=Q�@џ�u r!Dk)���&�׳��q� ^�H[���O�xl�駿�O�|m���(V���� ѪC,Yy�'��'��'���t���X�I��p13�՘m�I��J<ʓ�?�5�i�n7�-�$pݕhB�/�V�X���=R
�ɣoY��?!��?�#n�E� �����?Y��?9#oy�)�� ٥��!D��a�b`S�ə+.�����#l*ܒF���a�D��?�H�ǚ�~b`˓e�����ɡB$�����^ ���J�P�R��� ���퐷a!S��H���䟂�����Novλ8N�	��!��D��A�w.��Sʸ<Q3�R؟�������?���MKwC�z[*q�@Z��tO^X�(Dyb���F�-b�ЧUo��q`��~�rӼnv�I�?��fyr��1U����nP�L��@
@��p,�B�',��'K맴?i�?����� �h����S�G1�IK����
y��w�Ї��Y1FE�/ g�#?Q1jʠq��L��W�w~~��V�ӆg��9`�O�vo|q�w!��j7��9Ռ��4Ԭ�o��O����i?r�1�]��0��[2�D���#例�ڴ�?�.O��$*��� �QT��
k��ZF!̇t-
Pч"O��L�45Q�HW�_kh����O��������4��'�BV�D�w�    �"O�t����Q�=zw�U��f0�"O8��3#E�>-jTJf"F�3\�w"O����_�>��}��ו�:��7"O�M��� �b��0��Hb�"O��h5j�X�\#P)�+��p�"Ot���&��U7�L����\�xJG"O����mܠ�T�St�Q�$�� q"O8�;dO<��XB���&�HH�"O�L��Eԑ�48{#�٭O����"O8p��g�%	�TB�<$������2D���Q�?$��ɳK��v�!+2D��sQ�Ah�XI��.|tySW�/D�����r�މ���״r����.,D����g$C��
�iT��=[�./D�p8cN�,D��9#M.!��I	`�0D��x�&>�|��S�J�x\pɃ��.D�l������jG�GI�B��F�7D�L�0D ��W�E��89���5D�D�Af�XKM��#C�@B&e�v�5D��H��Ϻc�쉩�Bݥr���4D��2F�3n9 � ��Z�dd���VI4D��	K�o@z���F�-����g�&D��1aI#I)"E�5ءh_�p���'D��g+Ӭw�N��wB��u��Uɓ�(D��R��8X������w^�傤�)D��J�E�*f��V.�٨��"'D��F���p
	P��c�xeBb&D�P3�oV�,�2�9 ɘ+i�X}�h/D���p%�X1&����%">5S�0D�����I'������#v�q$+D���2
�5J���ڧJS�9�V��0�*D�(���	��t�� g��L'F�(�D*D��ʇ��-����QC�H�a�l&D�H*�g��c��HPBJ�v'�dy��0D�(��������ۂ4�D�@�/D�$9$�K#FZ��h�n[� L�t�.D�Г`�F&n�F�)۽:TȺ�1D�`��� ��p`��W;�\� �.�8�O4�@#k�Ń1����(1F�t�<��"Y*f����)E�2hT��"��k�<Yd�<�
(0�G�V����H]�<1���K���`T�)\}vT�$iN\�<'ܿn�m2a�^�4r��c�՛�hO?�ɭ�٧�O�G��8��DH-!~B�	�xd�d��A������mk�TB䉫b��[7�,�9�lS�~R*B�	�D�BuA��\���q���O b���W<��q��*E����GC"5!�T5��a���e*�fH1\|!�d\�j�b��cG��A*P$��]ѱO�����`�B䩓oůJ	"7�N�aB6Oh�B@̃�!?�ZǢԾ@7Zm:W�4D��ٱ�ϽPef��mE�����
6D�P�'�L��~H�TB$fz.�%h6D�`;&J��W�H��� �M!D��>t06R0oZ(1~�5�T*D�� &���-���<�Ɯ�0�v���"OpX���1Q��]�'X�#�љ�"Ofã��$: 413�	n�U�"O�B�����R F��[Y�x+�"OX��0�_l�8��+Y�Ò"O�舣L��2`l�)(I��"OX�1�DH��a6˒&yH���"O���C_�U{�p{D�M?H4u2�"O��Z��Ci������4I�N{q"O8yy1�Ҩ.vH����"��� �"O��F	����Fk�>��)�"O
My&h��C�*�4��i�L��"O�qȔa 	��aQQ�47�AyQ"O~��s���h�R�a��4��a�6"O"U�u�&�`������^�p�"O�d0Wkے�h��sj�v���"OL���	��DP��ıE�ZU"Ol��B����h҈R�x��"O��`�2,?��a'P�I��@i""O��tL��f��Y��4;�Z�*F"O��{�F�.�Ҹ���G�&�@�"Oh�rƂ[[j��C���Z�fi�"O�|�v��;�̪�ٹ!�.��7"O��:�nM>����++��q�E"O��x�̐����8�W61��9ks"O�Ͳ�*..��� s	�P���8�"O��C��[�b��q�HH�gѢP��"Ox�B&`	d�J�{�火W�"��$"O�aV�E�&4�Lp&�L
�l��"Oj1%J�: �n�� J@Y��D�"O��Y�ڼ���`��N�4�I�"O���֨P�0p�D!�x6T|�"O�%whG�j���9 �(T2� �"O�����V`e��+vb\���[f"Of��7�ݠ@���"E��:y��"O0����!�hH1W �1]�v�P�"OpX����R�h��`L�D���G"O ���R��Y0�O�v����"O�Ӏ��+;�䉥-�36"O��d*>B��x6�*2�"P�"OV�h%êQ��U!�N�(:�(l+�"O� ōF�J-6Q�ͣ;]���'2�kS 3o"�mZq}"F�z%�����"��"Ӄ���OF��ڝPP�KB�޺ \���A�C�$����62�Q:ц�'0}���ph������`>ʓyy<�3w@��_(�����
]'0�	�@�1�pܣU�7c#bM����9*��(�%m�Y��O�oZ�~��.�djU%�W�p: F��~2�'���D1�S�;�,��K>Xd8�rw@�|�:C�	"F֕a�dQu���C��3|(�qn���M*O���Pͦ��Iџ�Or��27�i��ɂ�T�U���@�g֤�.�Ks��O��d˘`�M��ƭzDX�i��U�XP1��>$�,�~;<����P�c��@e�f�*E%���b�ƾ������`��[s,N�	�`�� jS�(���q��(+��S!�N�Z�@8D��rT!�'�l*��p���1ҧ�u�ƈ�{����3��M� ` 'MɨO�":�ċIh	�B� v�nd���`8���4M:���xb���nq����&�R:�
':��n���Д'�pl���HO6���F9~���i���sl�5Ȇb�o���)��&�q��Pjg��'���@�0�杄!<z�)c˛�^[��B�;���)�!Y �d�V�� "6���Yܧ/�R6m|�Y���J��GI�.�Šf���!țFw}R+P��?�}����n�J�H����Y�d��nR�sNq����=�g�+���@�+V�v��9DPA������4��������� q�Y�ץ��5b�ƸU������P�	���	�ug�'��'�2)j�[�Y����-Rc@��e�%DU�p�t�׮Xx4};6&�1cF��C���(O�|��D�Dϐ��fK׹ �~�⡨=H��P�n��K�k�2�6�G�5���6��i�� �"�03}N5 Յ�6�j1rCmҟH9۴.��'C��'a�'-����[^�1��k��|L�F�9�p>�I<� ���$M�#���Pd�T�T�����X򉛫McB�i\�I{�.	��4�?�ڴm�@��
��R`a"�(.�8��f�'�b��g1�'��jєh��A0���3������X�Pm2���L��A��%�� S�y˶�����|��uk��T-B�x��&�_�C�|<%gS=hȍ�vCM�m��C2��HO��S��1]E԰ҒG����C�<Y�JڟH��4h ��^6z��޲�8SA�*S��O��D"�)�S�gU�Y��߀u�*��B"=����9�L�	�Bߧ/���K�
A m>�I���ܦ�'�kቩ��D�Or�'q�T��4o��� ��xʐ`a Ů���&�'q2�D�/r�${�L��X� ��^�Nk�����˖.���"f��g�8��߁{؉'��y2��0�t�@Q�e_ ��r�L-�i:A���."1{PK�!	7�����-Q@��h'N8�dY[�R |�-nş��~"&lװ_�!5�3\ЀD��jܓ�?A˓P�
�³ ͔j$���e� cP4F}��'��6�PӦi'>��d.	�T?d$s��.����H����	]�Ik�'
��B� �� 8  �9�75���0�]�Ȇha��Q �$*�ܕ^U���J>�ۓh�J� �  @�?AZѫf�&Th:��CFQl ��"�&Z��3N>��ŕ�܍��m[.UPu��[�g5��R�}�n�*��T�4�������z-���V7Ej��!`W˼�� �vXQ��P���w.�J}�����?�4�i�Oh�$�OH� �i(!g��L+��藫�/�P�D~��Ӊ��`���"cl����)9j���i�t7�)�d�4��<D�����r�U ��s&ݗ:��-��_=�?����?)�;� �SΟ��	��� J�;�]��r�cGY�
Ԓ�Q�>5�� �˥B�^#?9�+�XV.1h�!�4&��	��Ӥdab����d�󄕃 �������o�`����o�`�	�O��c雝l�Х��dPj��"S��1�M�����O���'b��t���w���X������ȓyd&���d�V�Zd{�"M �T����'�d6m�Ȧi�?��ē{�h� @�?h-둸�l��t�?�N��l�RQ�֖�i��>1��ɚ3���G�A;41��jC[[�a��J
�X��)�Q>cS�Ό)�L]�eB�>P���>	E��� �ڴL���O���4��ҫJ�5����eݜ2�����>	���'R�O0�!�,D��$���%M!�e*���>�M���i�'���=k�y�5M�Tg��K!E�$yӮ�	Ɵ���>iT���H[����ȟ��	#}��΋�h��	X�M� xsPnZ)c�fD%�\��jYa%�C�3�:4ݟ��	D2v~r9 Z���*�!M>�"�!TMU<�a�
��<��ɛŜ(V.�i�������Ì\:wV��ٝ~u� `��|ޝ�o�J��5������ǉP���>r�f��Kަ���������ҒQO�n������c5��D{���'�Հb�b���Y�b�%k��k�'X�6�
զE&��S�?�'"��P�h�V��A�ۤ(��-�v�U�k�7M9<O���:>����ǯ�0��]q�Ő�fj�/�9�%�`k^�+�����H���z���Ʌ8�걨A���t�v��#g�1�F���iܹ2����Dț�
��#��+�`;�r��lZ�)�L˒��)����׊I�,�$�G�i���O��d�O����[�p\�q	����k �[3JҠ3��'�ўb?����y*���ub��+e~M�1}� gӲ1m�Ky"ŝ=V`6��O|�$n�X,�q��-#Z�9go�XA��֟�3bߟ$�	ɟ(�S$��`X�i�$�����ʒ,Y\�j�K�>/h1P���6
�Haxb��7"�x�<1�+�c���+�-
�����U��|`caD��7�(,@�� �Y  ���")�7-]2��'AVpc�z����4�����������C�X����w+�"p���O@�O�"�N߄aD��ї��,`l�̈́n��hO��Z��)�7�ѝE������Y���ڎ~�%�'���Ӡ}�~���O��'��aS��M����z�&\�u�����b�H�zXR��c�^�ٲG5T�nt�t#͖@���6��.�SֺkUM@�z�t��p��V7Dqj�!�Z}�&Yap�5�B�W�;�d�U��!dS���!��!�8������Pj2�s���V�d���*�CXTz�O�>��џ,�42��O9����:�h��F����p��'+(r��>Y���0=a�H�&�6���[+���R�Q�<��4O����|"���LދS8�Yv��&
}>�i3�O��D�O�d��&]�NCD��O��Oʔ�'`j��V�7�|0���G�t��<y'Z{(�7H�e�y9�����O����<i���F��p�� ���S��&O��Wρ�g.����+9�aℼ|�1�Ţs�.��3����"���̽�����k`�(�M��c: ��l��	ğpl�eo������,O`D���]1G�C䉛:�� 3o 'u��-#��x �����Mʛ�D~����|�����H<��
�g�Q�Y�.�x���x!�X!UR   �kӖ}�}cN��!��67���ՅѴ3��Z�j�a�!��J�!��J_���Y �cՔ#�!�V�B�8�!O�VQ�z���B�!�D��(�R�ф�M?(��JY~!�D��L k�bgA��܄Em!�$�#<+DA���N�/J�	���Z1C�!�*@g,�X�j��
2Z0ŝp�!�6	H����[�t )9t��5�!�$_�@X��p����un���#ӊ&�!��e<D,I���!���7F�����'���2ɗ;(,t
�l��b�8�' �ԱpMn�H�A#̀���	�'f��Ƞ�O N�K�d� ��Q��'[���Eלl��-�����t)��[�'Œ���k\,wНѰ)�W�J���'ly�p�0F�Z�� e�{gX��	�'�llX�k@(�~Uq�+ҢGg����'�]�׆Q�U+�%	�fGC�Z���'̄	�w΁V��`	L-D��̓�'8$�aCm�x���I�>��l��'���җ�y ��KZd��͸�'�~5�'�\�G��|�b��'۪���'�.�(��MkL�L2⇘�k�"�K�'���d臓����D\�(�
�'�~��vϔ�m�~P�"�OY���	�']��G��G���o%o(�b	�'np�-��a�
�Qf\�>���h�'��f!Q�+�d�aC�&;*�T��'$=��� �n��("�M�_��YI��� �4���4�%谣	'��i��"O�T�� �!��Tj�=;�j��d"Ojhz��Ӗ����3�Q�%�U�1"O,�	u��9<D|��`�?͜Q%"O4X�A� �(A�ToŔ"��i��"O�1 w�Q�7]�ɊQ�_��X�Q"O4U�CEצ$���b$ₐ`(2�"O���R���Lf ��)##"Oh`zA
�.�6�c�Ԩ,jR"O��X�Ό�(4YG��a�:�h�"O�a 5,ʂr�����Iy�E�S"O̥ɂA�CʭeL�	�=:�"OF8rѨ���*�SB���+�r$��"O�訄��zCp'����""O�pi��$W�A��kѶ*[�ɳ""OI�+Q'<&��(9y&���"O.�B��>�tvH�;PN0QQ�"O~A�s��A���ŉ7>E�k"O�T���7b�`���eP�zN֙+"O�в�f��Ш�d�%G*ڵ"O.`ѴOX-'8�*&��:�ֽC�"Oll��W�m@�a�e��:>��9"O.d��C�=Aԁ���Ўg�$���"O|P#��@�p�C��V%�B"OZ ���I�"Jr=8$���H�\XPS"O�]�s�ݫb `�s �+̴��%"O���œL#�ɲ�ׅ?�Ĺ�d"O���R#Ҙd�\8�k��xH�F"O
�P�$�9_Z����^'�d�0f"Ozh�N�頀9���`�T8�"O��O�X�phH�&�th�r"O^T)��Yu���#�%͑~�B,9�"OD�`ےAu��H���)��#W"O�0C��� %J���}n�A`"O`�r�O%<p-�'� Hy�y�R"O�C!�S!�.����V$\\�5i�"O�d;�DQ�C%̀Q��)J�0�W"O�59�>,
zpր	�Hn�B"O�u "Z-�<m�W��`-ʰ"O,�8b쏬-o�2ł^/����V"OD���ο/�����CP�H�e�I����F�pW���)�:Ri���R�O�����,���qO��dzD8��L_�'�Z��d!J/^Z�;C���4lއ����r,�S�a����Q�'���k�7�vQ���ҜSWj�ٶ��{�(E+�Ήs�8:F_�w�89���.r�t��=�B��X.5�Z%>�o!�ȁ�`,�S����cW�\�����'�>�n�H�E;�NM�a�R�+��Q=kZ�|��f�foΦ�ä��)e5(p���G�`���륊��4	�<�Mc���?�.��(�O ��(A��IͰ#�\}�"��/i�XA��R�s��:��!Y�Dh�&B�W��فo�-��y�OW��ư��-I�?�v\���T�cx��Y�i�j���%_�[��X� j�.�>aT�	J�Q�iC2�*�Z0��5�̎�T9��-Bz' ���G��Mۡ*G؟��4`4�)�)#n,���`Vhڳ}��x�*M>X��PF{J~��*�AqfK�0P[��4"Yb�'ܼ7-Cަ-�B]w��8	5$�()�@Z�Ø�]�Rʿ<�%�l.���'"��0��YL���k�v��FE�8'�ɩ�Ƈn&��nWU"���U�mi�|	�|r�C+[ƢaX������f"X;R>�s�B ��)̔L�:�rB�r���\ܦ�hO>	�j	�y�b��T�h���E�B}�����?)"�i�p,�O"���O��+�v ��J#x�v%�����Vx�UF~b�ӵi"U�vh�ݤ̙A$ɑ q]cѳiU\7m$�D����<	Uˁ�f*��F�bBm{��]
x�8P��?i��?����0����?i��M�ѳ
	.� KA$Pѐ���M�u���BR0$#Й!��ǂo��-�T�Rv�'����a�)4kY+��B�m0V5Z@�<�_\�~L;�F_\�5*s�i���ڴ%���'�l)qE�O���� �/	�� ��[�2(q̚8r�%�H����&��%>�Î.h`�Đ�H� ���8O�#=Q�^}�T�x2�8�^����x?aT�ib�7�<1��9P]�f�'��W?� �I�5����C�Y�hRl����?}XV<�I��P�I� HmҶ`ș>pF����[R�Y�q ��I7�0Â9V9�3��'\8F��p�=ʓ%���s�?���0)��o]�шJQ.q���g��!��)�2S*���:>�U�l/��D�0t�R`tӮx%>�o����8��\�7Z-����S'^�!�������"�ƛ"��N-D�Z=�p��ē��O�@n�8�M�ٴ|ਓ�J	�8a��� �7R�����F�i���'?�S0[�b��	ܟplZ�0��*�≌<
���o_7?�CIL2q*vȸp�-O�$�Za��8�ʜ�7��i���XL�h�(aΛ�0I-��,P�p0�6P�'B�ŢDG�\�P��.J�B�]�G��֝<Q�F���W��89� v�p<��@eզ�
'G�On����4�?7힍vd*	�I�g�`=�IV>:��hO�\��@"Н��h&%}�h���OJ�m���M�K>ͧ�u� �^������L�s/[8�0�O~����rv 8  �B�`Z���;�B�%�ܠ��ϥCb�HA�4_�:���*�"��'�%oڴDp��0S������F*_3����� 9&��5R����M�Đx��'�[�qOS:��P��]�,�5�;������c�)��]�rU�u�@ k���J�nK��M�s�i��'��4�O��	!��#�I�q���r��
FmD�a��Ab����	��$��ڟDp�M_����	ڟ��7!�w��]*4�O�'�������;9��'G9�b�@An �to�h�pEބe��<��'�  ��Pز�QIU��RS�ѐ&D5ᡴP��R�L'V�Z0j]�M�Q�D�U���>���XHb��ɲ化:��yPN�]R*T��ęR㑞�F{�i`r�)#��0g���`�k̑�Ǔ�HOޝ0�	�<YءS��Ҭt�{#�O��mڋ�McI>���?�M<�ԡ�5 .  �S�#�)� D�'U�b�I)��l����#B�4C>e"�K�c���?�w��R��U?8�ba"d��=F�(��^)a�u�kؾpd����>D<��Fx݉�vO�|r�4r�
C��x�TFP�|���5CI��ĠpӺi���I���i>��ē��t�m��t�Z���ʌLr2`9��)��l1P���������<^�#�§���ɺ�M���i�ɧ���O<���<�n�����&��(�b�/k����i؟�	g�   ��醧R�'b�pk"�٘eCL���ג` �@�|R�'^$^��I�;.G��
!�w�^�3�t�cԨs��4@��KK05�"  �" R���&�T�Oq �]Z��##(�%;��x�vn�*��e��z��fb�<�.�o��?��G=��eT�
G�]��X��kß4'����I>��ar��ʤۤ����� �'"�d��l�F��?��Sɦ�3'-�/h_�s��K�&�V� t�ȿ�?Qp�8N�
 ����?1��?�S���d�O�7��O�ƠQ�H�4L/ܝy�i�?`͊�N�����7DљN�DA��X1j�.4P�M"�I
F����E/Öq4�ZB.ڳA#�mad��<U� P��GG-!�8Q��u�}�e	�>{�\ЁmD�x���T�i;& T9.Pd�����3T�nZ;l����̦xJ<���?II<a�cդ~m��@�� ���:a�l�'�ў�'�ؙá(Y�9��D�FL��zx���W~��OjEo��?�'���){�$7-�d�%��hʟz��Ȗ-ĵY�Bu��ʟ��Ɇy�Nl�	�,���S�v���D�j���s�fNlu�TR�l��N�K�
�;� $��A�b��9 �1�H��J6�ҳ+�Ĩ�6g	�1���C�H)#e��"΂�`|d���C��M��BA¦Y���5�DE�5�u��@w�<zG*rf/{�F�����(O�=!�O��h�
�� �I�U%�-��X!���N�O'N�ڕ��+��Q��K;�bw�즥i�4���?A���Oh��@ ��-xC"G3�)p�����DAH�ga����O?��~���&��Y�O?~t�2q�	���O���.PB���N@V�8.
��b�f�'�|7͆Ǧ$���;d�A�
���ԙ����tL)Bv�'�2�'
��ր�"g��'���'\)�;L��pp ��TL�1 /v�����ßGh(�&�
�vHtl�?=��?� �D��<a`-��(g�u�	T�j���jF?��QCq��:�A�EJW��(��|��4h��Xm�ݼ�G��j�~h���|S�%rr�Ӛ}�6�H��}��7�MkΟɧ���8��}3�X�jH�a*A�'�ayB�)LX����C/A.x�6�Ĩn���$B٦mc�4���|����ē1�65���ƭ0���HS�*FФ�O�HR�   ����X��ܭ��ђOl.%o���P�'�b�'�©L��yҘ>��ͻ`��rI�94ج]�e����	ß�����dȖ�!�M����?������7�&�jun
�4�P�
����Vț��'R�	�����a>]��Zy��M ��w^�)A��S�EB��`���������L9��ɗ�M��?����:���?�B����F���E�	~f�p"��8��	şt�"j]����IHy�O�,Z<<�kA.���Vo�@��lڴp~���4�?����?9�'�Z���?�����PC�&;����3����Q��io�=�t�'v��'��9�Ow�OA��Ɵ"Gp���V�C� ��P)��a��7m�O���O�*�L��������0�	؟��i݅��B��%[*v��_����$�y�H�$�O����I�B�)j�'�?���r2\�d��;u�.��d&F�WxzY�i�b8`�6��On���O.�NY���O:�(�&Л]�,D����[$)��iz$��dL�?�y��'���O���'���'q�r�EL���|�a�B$(<��ǅ7P��6-�O��d�Oz�$VX��Y���I�<ɢ�:f��g�*�ĉ�+ 	n=b�,i������g��������	�H���yشT��Q2�f�@E^�XT�Q�x�3G�i���'�"�'��R���	?|6�S�79�%�u�˼j�x٥%��`�K޴�?I��?���?Q��y��p��i	��'�n�C4A�8砜!NA!2�b�u�����O��$�<���Cc��̧��<5)j q�C�7tJ%���8��7��O���Ot�$��Zf�i>��'1��O9j<Jp�ˈ)7�9�!�GuthIgokӬ��<����|��'�?�)O�i�čaW��N �`�`l�������4�?���
~b�ɧ�iu��'��O�D�'��Y���-(�������f�p����>��Xs�8����?I)O�)?��O�?����t�z{,���Ш�M���1`���'���'����O�'�rL@�]�����$��YQ��M8��6�N����O��I*[D��!���xz@�0+�~ �#�$|u����Ѧy������Y��#ڴ�?	��?Y���?�;4A�1qeD��h��R؂MmZ\�Y�b�)���?��;i� ~L	c�V/O���1��N�vNYS!�ii��\9��7��O���O�����4�O,� ⛹�̙d�s�%�\� �oa����ϟ���џ<�	Ο��	;G��,)Ub�	k$������,�I�%n�,�M3��?����?eZ?��'���Y�v�4�{���	�p�Gɛ�Y��P�'+��'���'��R>���W��M˥��vWxIH6�7A���K# =g����'�2�'y��'������S�w>�����.XgPjq!�-s���4���M��&���!���?�)O�|���Ky�S/X��eb��j�����W-I��8kڴ�?�M>y.Ou�g�DG�l*r�r��!e"<+IO�9�&�'p2T�(���I��ħ�?q��|*�@ʦ��wXP9ye�u���R�x�\�4@F8�S���K�oZ���Э!�ڠxd�3�M,Ov904�㦩S��`���:<�'�&�H#`@�[9��"�#F�.A�4��d]M!�b?!���>� �rIQ���ECc�4$;!A����	ǟ����?H<������U���0R�HT;��hd�i�x%0�����|�i؈N����`i׶+�v�(F��M����?���IȮ�� �x��'�O6��ңڗ>��Uؒ9X�R�����/�1O��$�O���J�=��B��� :��q�oJ6y�FIm���D�`������?������'�1Y���!Ȝf�ODj}O�-'���'��X�pR���"IsR��e�+���Ee\�\
�L<9���?K>1.O��s���3L䔱3���B6qk���5�1Oz���O��d�<�IS&[�	B�TD��hVb^� �����v#�����}�syB���$�9z83'��R��d"U�W�	�$�	����'�މQ�$>�)��c!����^6:��C�E�!��lZ��X'� �'&pIڊ}BÇ�aLp1��YAϸ���B��M��?�(O�$�p�ٟ����aО�bF�� L�uAd�]�VbhM:H<�*O"< ��~rr�� F�>}@C��Q�z���(���}�'�zQӖ����O���O1��D����v��/INČb�l�iҠyo�~y�gܪ�O���`�*��qn y*��:y��+ֻi?t��m�����O��dퟲ��>Y�ɣj$�يq�S�K�b�q�+9՛��
��O>��	2���@�"0�<��4�6`놔��4�?Y��?q��S�VЉ'a��'�r��ec:�;g��=��� =�c����$&�ş��Iğ���һx*�݂!��:<H���̏�Mk��q+J�Yu�x��'c��' �i�ZW�� �V����B-�U����>YS�W̓�?Q���?a)O"yQ1�*m���k[>��I�2��.]x�&������p�	by�^��Ha`\�#��t�P��3 ��"�#m��c���	蟼�	Gyr*K�=d���fM�g�_�2��Q�F�V�̬&�P��埜�'��	�L�Z�'�`qC��%�"5y�P(�'g��',�R�����ħF��qa��K+��#�b�(uY�i�b�|�Z�CK4�I=`��$��r�fL('��"�7��O����<aL�
x��Os��O8`-�HH?Xv� #�C�a:B�+VK:�d�<	�R���铷SW��'oW-L3t��D�F���fZ�LA����M{s[?���A��O�9�̈́���X;s"��W�� #��i��I�#<�~��@��yB�⅍Cb�֎�� q�M���?������x��'�v�Q���VA�cIƗ6��az�g�bȹ`�)§�?YR�	s��Jӏ�)x4HD�ãb8�F�'h��'��	�`'��O�����L2�K-4���B�X|�&.!�	�m��c�@�Iݟ ��?,+p*aN�T�I����'Q��	ش�?�$+95�'���':ɧ5���В �q�݊D����ÇLa1O����O��Ķ<�4�|x��:�kY*[u����-zT4)���x��'t�|�S�H��b�:d�𝁱�	�8f�ta��c����Ɵ\��YyRe�j�j�S�oc�Qv*�%����B�)�h��?)�����򤒨{�I
� �j��$��ZQh͕>p��?����?�)Oꀉq�Ec�'@Re�d芊t�Y�Ӄ'�z�ݴ�?QH>(O�T	U�?9D�x)�yz��P��U�+��v�'C"_�StD���ħ�?��')D�x����eP�ib�AHA�;A�x�T�D[s+�S�$X��A�/	+X�x����9�MK*Or2%K�צ�­����។u�'(8��6�3 ����+
=r���0ش��DV;#�b?y*��ٟg%B)���&q!�y��|��C��覽�	ȟ��I�?�M<	���X%��E�2� 2I�&���i�����ϟl	�D��VmI��?j� ��� �M���?��^���P��x��'<��O�=y�+P��p�+-}"��5�d��J1O����O���.A� !�F��U8�i"n�	Lf�n���z��F��ē�?��������^F�\�s��!]��c}��ݔ֘'6��'�BV���3� �.Վ����A�^�:�k�04��J<��?�L>-Ox��A���"d 1*��E��Ɉ�]�d51O����O���<)R��Z�� ��k5�:I U���,65(U�@�I�($�D�'�JDҨO�a��&2a�%bRm������Y���՟$��Ey�J�C���^a� C�NrA���n�l=��ݦ��IF�I@yB(�0��'���T E�+l�X�"ʈ9�f�b�4�?9����J�$e&>��	�?iє�V�GFZ@����d��H*�!+������+���D x1�Fפ2�x������U\�lZ@y��S�{fJ7-I���'����4?�aB�*w��z!�H�����l���'�2���	�s��}��H��5P��p�V3<���۠h;7��O��D�O��ib�Iޟ��7��I
XMC�$�5�~�iϙ��M�F�M:�����y�'$e �Z(R�i�v�F:�ܢ�s���d�O�����g�ly&��Iퟘ�	�k��1���%H�˞4&L���
g�!b�0�<���?��>�����"@]p|�DN�jU�Eؑ�i}B��hnNb�T��ߟP��5�g�"0uF]�`�2"d s�h������r�y��'���'�剁/#� �ǂ��xZ�@m��R	���Md�	͟��I`�IMy"ϗ0���r�P�K���ʔ���
�L	�ҙ|��'���'6�I�\ 6`(�O�u0��Y|�B�.F?n��a�'��'!�'��'grY��'�:�2�U��س�Cֺ&*�Y+D��>����?������H:@8��&>�`�_�>�A�g"�I�d�a�+U9�M�����?��?͚0;�{ҁ�X) �M�82j�<2��\��M���?/O@ Y��^K��p����M�3�Es2�t�I��^IjN<���?�`E�7�?�J>�O����@�&�H�C-�$v�~P��4��d�2Q/��oڒ��I�O��I{~@�J�F�#",�=c�MPBc���M����?�$���<�O>�~����yHpm� ��}
�U�!�զ��E�H�M;���?����j��x�':H	Ӎ�	�r�HI�	��}� �g�n��0O�O>�I;r���*�n��?�����U%�%�ٴ�?y��?��g��x6�'bR�'���<���5ᒵ	+|�I�4M�Ol�3c-���O���O>@R��՛.~�z0�Ҋ&����,�Ȧ��Ɍ5yڸA�}"�'ɧ5��H;^���# :�J�	w�\���]�Nr��d�<9���?a��򤉵�S�)YV��S@E��bXH�ODq�ʟ@��L��ʟD��:m����R�V������Q�]�7���ؖ'k�'�r[��3�ѯ��4+1J����CS�df����$�OJ�$9��OH����M��%�:]ӵ�K��"�Ywn��j�~��'ZR�'��[��F[���'Nג�S��L��E��F�V�`���i���|"�'��b�y��>醭�8,�%��]�Q�fuS&�_���I�'w����<��O6���8lMT�X�낲)�t��^� ���$���I����0c ʟP$��'l��6)_�����CJީ��l�ay"��UH7��@���'>�T�4?���U�IAt��J��a���������(��z��'�b?��̓s�l���N��rT��$*~Ӵ$ʑNNͦ��I՟����?)�I<��kf����D�V�{s�W5jn��+�i\���'nɧ�D��<z��(���u	J��D��B�PXo�ퟔ��ɟ�K4O����?���~2]�}E���^�J�kl��M�H>�u�����OI��s�5yP���&Q�K��TQP�G�O����ŘG"��م���t�T͙��<e�[�W�����Bq�8�¬ɀv}(�87�G�&�$�xW,���cM�l����$�J��h##Z�t҂H(�AF$c,BhLX)vZ�bh
8i5�����(��E2 $7���3BC.w�(�NS?5)���m"]]�4�$�ʃqGR��SMԑ5H�m�SD��[���6�'�����܍(i8���ωXoR(��Ó�5.�͂j�
x��MQh���m[� Q����0b���'��xKQ�'R>��Y�)���у����V��9d�w�j���ތ��e�%,N�?)��\�oZ�J0̋]"FM��zT��WŢ<#:��w%%j���D%בJ���Gx"	T�?y���d�5���hW�2D}�ㅪ7�1OB��$Q�e���"[��)Bt�+�PxbGz����A��:0�Ts>>��p9O,˓D��Ļi���'l��:�$�	�:����^!��+B�1VVh��֟l�� �"T�b�c�>t��0�S�t\>��i��/Ħ�3v�<�r�z��!}�K$#t��D���в���i��� t%�2h�0�ͧ<t�H���+%�D��1��
���O��W�']��O���pa[3*S^��ČT�jw�u�"O ��CY2֖� �+O���h��'5,#=�穂�D�����1�N�Ig&p���'���'�\Dq"�I@-B�'���y'��7����3w���#����f\l)Iq~����!;�2�k7�|E1�rU��k�m��83k�L��c	��m�$��Eh��
���S��ɭ��� )�� �;�V�Q�Vq6@8�-	�c�MhA������/Of3p���d�O�O�Q�_/W� k�W�~�4�#�"O�D[.9�)w�3�f,㳖�|������I[ybh]9( ���N�*,�X6M��+�2�P��590��'���'"��Ο�	�|���R�uC`�R��t+akX�$��b�I�,7x��o�+&�t�c��R�X�<�	8� �q�F���/�`�@`�!y�niC�_cZ���㩚>S*�3�ꆉ%qIE�ɖV4J��S���K�};UF��"��-P�/�O���d	.^t^�+ �|jHa��kL5^K!�D]#��Y�g%V�(f�bT$T�]�1O�mh�	"TJl��4�?A��LC$H�C�ڽ=��)�P�G������?9����?!����4צq耨S넀p�eyG�i�
	B�Ǐ#��y@�HU-�Q�	Ǔ������>EZ��C�q��������H%�a{E�)?��Ha��5k����7E�-nT"\�<�wE���ZH<14,��?�pgȁ7>^y@�@�<ᵋڥj5��bbaI+&���*_w<B�i��в�C�[Bp1���ܶ��4B֟|���0��6��O��ī|ON��?�a����$��'+�DJM�p�I.�?���u�RK�P48svT�b�X�y*�"�'u\e�׍��r<����<Nn��O>EW���t	��;����..�.�@�`�|�i��)뀧�(`��<��'�_�D�Qg��o�n�o��h���aS�!�<i��,&-D(i��e̓�?���rU����sZ���%V4*)�}��	�HO̡�"�8%�eXVf	�ی<q��\:5"H��O��$ Z��t��O��d�O����s�߫�@�����j��X� �ט'�*�yϓTeH��F>Լ�v@�%\�V�=RMwx���!�>4j�:���i�-����m�=�)�3����8r/� ��yX�,R�Py�K�/�d���W4ѻ�����JP����|BJ�,\\I�A���m�������%Bú����L��'�2�'B^םßT���|�p@��7&����;v�rexT�?>8���`��K�g�>1Zz���Mٺ$
�I`<q�g��~g6D@�"ڿCPrm�U�?(�Ƙ��|�����K+S�A��T�Yd���t*D�t�&� ���2��|x�4k�%'��-�McN>�gZ�T�f�'rn�<z|p7�)8{ �1rOF�R�'2`��'�R<�����'q�'��(���l�D�J�0g����]� �?AT�&'Ea�ѢǨs��eP`�Pv8�1�m�O�'��v�̇�b=IFi�<V?|1T�=D��!��B[�h Fj̼��)A$1��޴T3��3�S�Ue�Pq�&�ZpABM>IπV�I͟ �O�p�D�']@�1��o�4x�J���,b�'>b��/y�x@3�T>��'LA�	Ը6c�CMU'
�t}pJ� ��0z{�c��?e�` 	(KV~ �9�a��d5}" 
 �?���?!����O�t`�k�$&L�Iw#Ɇ_��4��y��'��yro�)1���c�p�2���/J��0<q��ɉ_Ğ��2��&�9�v�ӆ~\���4�?y���?�@��nv(����?q���?��; �d9����=D���*�k�=N;�L�M3K��	9w{�ɓ5���1O�Uz� �~8���E`���%wer�C���nW��{��Xo,�CT�i�p�DʱÖQb���-Tw��(�ݡp�	oZ �M��*8H�A�S�gyR�'������ Y��q�Ch�V�| 7S��G{����)J��� ��9|��t���.E|�	��M{ĸi��'������Og�?K�.��� �*Z��m�e�>9��2̝3~����Iȟ��I��ȨYw���'��� +A���r5Ĕ�>'�M�F�.< ʱ��ODp��.*<4H�hF�m��0�RdD*�!��/*nx�0
Ɨ8n.uK�D�!��t���'b��$�Nc�{���	%f̈$�B�,�!�D����2�W6 �[��Ȫ=�1O�4l�Q�	2e.�aش�?���]Ip��"+ׅ9*P�ˣGMZ�Z���?yDL]4�?)����T�ڞ�?YI>� *P�2�֥S��F,zB�$�^8��"T�)���+�����R&Po��!G�
vn����ԗJ�"�|bJR�*o��{F��1�>E�6k��y�*���H���>l��ȍ��xr�c�2��rdT]��q�#H֋\WVQ�V3�d�OdUl��$�I{�t�	8�B�B3i��p��7d�����.�b�'���"�&�
 �h��<�Oa�S�1s8�H�A�5�d�X*ƥ�Z�',Py��X�suJ9 A�<'iV衃�U0(���OA���á�){���C]�ĝL�HCѯ�O6�'��?X�@]�{�:Q���^#~&&�p��9D�3�N. @�P���:|�1cG9O��Fz��@�@�*��Ddo"ш�ܑo�6m�OL��O�x��M1T�4�D�O��O󮆸R<��s@�cf��eí�hb���G�/<Op�	�B ^2�eB`� rv�St��_�y
� ݻPcդs=8AŁ^�~|u��'扫|t���|��ߴY> ���\34"��@��y�G�=L�L)�n��* �I�q+����D]����|�-4�`]Zɓ�rެ���=!�< 1 g�B�'wR�'�b���d��ş��"&�c�*d�/\�u��&/4�� ZU�J���>Iw-D�f�d1� Jr�^�k��)6vڄb�HR�}m�� ��d���b$�J�NP�1��
�0��@�+J�:H���O�nZ��l�'5��'��',t�z"ώ�6�8�a�5\���R	�'�^��'���!�Uq̋�%x�Zg�|R,t���lZty�a�
�@7��O����?9Z��C,�)�� "��;;����OJ�k� �O^��u>�ʀ*�OO�9�B��tE24; O��(=�PR�'���jހ,:B�"��Y�'RP�`��=�p<1���xJM<�L��N���tL*X�)q�%b�<����:�ő���G��H�m�^<0�i}@a`��T�H���կv�N�يy�l^�U�L6��O��$�|��.���?qr���/�r��3�M�8X]��ϊ�?���2� �Cؽo��`��/� 9�)�
�?��O��}��-OEȈ"2�5yOr�I��h��\��4�f�#x1bAY�4ň����eͤh3\w���W�l��ӆ)E�fQ�H�$���O��|��D���v>A����8l���rU�L��yC_��lxbW�3�pd.X0,#
Ó���4�4�Ŝ=�< �&�_�5Xb@���M����?	��sM�Ɉ���
�?)��?��Ӽ�%�G�\�饯��UL\j��Ǐ=H!SWO��i��%ɾ4˒����L>�/C�g��1E�\+�EP#L�w�r8u΄a%$��Q
F*���i�@��m��Ԩ9�2dj�E!.K���#�Dv$�A�f� }v���|�IS#㒥#���s�֨����y���<�,.�6�y��'Bn��'w�"=�'��"2���De�7M5�yA@hZ4�f�H�Ɋ;��m����?���?YT�� ���O@擝Gq:��b�D5��Mt���p!�c�n�5�X#ThA�m̲��O����͗�D���Zr	�a׀�s�"�FͮU;H�#���h�%f^���˗�T�`s��3���ZYHEmC�:���y4O@!H�J �g.�O(Q��iUE	f��) �ȷ�5TN"������ѹ���� ���+|Қ��<��i��'�0����q���D�O~��7AK��'T$R��/� I���'���i��'��9�$h(��i��<+M�q��mڛY�p1��55�)���Q0o�:��$��Լ��j?|�V)J�!/O�!sH�qV��˄�N�4���ěI�H����^����h��O��Od0Ԇ��xs��8lx�H��~�<A�O*Eq�䗚Dk�=��)Tw<���i�>��c��L�*�B��A�{�� [v�|R�|��6��O��$�|���3�?��FF>�Ty�f���&��]�K�)�?���a!��Ia��.i�����
���Q�@�?ٖO9"غQ�?V��s*[�\��lM�1�aX6[ղUA�O�h�b�#�`Gq�e�ŭS�������5�)RW�,�qv*	�#e�Y�O�I ��'�ȒO�<�$O�/�$�6%�{]hLB"O���#�^�FϢ�2��F�U|�S�9��|B �	,����e��zt8�A"F&6Ȧ)�ڴ�?A���?�a'!t�.����?!��?�;t���3�Ol��Q�/B�)T8�2�l��
�"d�DNQx��T�AEN���O��'C�8��JB�`�B���E]'�a"�B�;h���9]�񎞽7
�*O?�nZ�C���]	\�͒�H +4=���D
-�\�M>1�D˟�>�O�]�n�1έC���:f2���"O�q���>-��[b��
�aJŝ��8��4���O�8�#�:���
,�Y�|h7�X"d@P�o�O`�d�O���_��C��?Y�O�� ��(�^8%z��U�`
�i���x���+Q��@�K�(�p�Q8���
�',Q��i��l�yU#G<���:�G+�?��0 ����D�JW Q��e�0`��
�H[d&B>G��m 
O7.��<��io�'. q�k����O�m"�h��=�(����N���x���O���f	����O��S9
���b¡�v�	��=+���X!+J7��YB@�>�l��p-�W�'z�A��&,���fAνh0��QMY�0���С�\�5ު���ř((��F "L◡5��"�5��D;{�+Ն۳)P��b�/[4�!򤞸QU��ń�c^�+�k�E!�DAǦzlU;R,x��U�ߕdٲ��b�La���ڴ�?a���)K�c�DA�7�Ht�"�ڔF㊔�0;X ���O�Q�(D�<S�H��N����1�XH��R>��"O�82��,
v����ɮ\�B�'��$K�-Bj�J��TÓW	X4��>�����{R�I��Sl�a$@�Q�8����J�M�va�ɸ��S�g�? L�E,T9vb�Y���D<��Q"Oq�- ]�L���-7`T��'�N#=I#g��SY�e0�%ϗ�y��ʇ:s���'eb�'t@��Pi�K���'WB��y�����!pG�֪;&-X�L�04�1O��9��'	Z�Y�:lϒD�EY
@9�q��{�����<���H�q}b	0�)�-�nLAA9�'�fL3�S�g�I�3n�x��ƪh<���DN�_I�B�ɐ|�b��v�L�)��(�j�=]���K����A�E�0��ǥ�;`(pK�<t\��S�iM��������I����_w�B�'�󩉽Į�"�LN]���bG��#3Fu@O YC$f��6�>�hv�݊B��*!�[!����6�����\6
ѐ�ˎk�p8��'�"M�D�7`KDe,P���<�yb�D�~�B"�Jc����,����'�Nc�����[!�M��?�6jՎ�,E���R8n�H�2��?Y�T0֐{��?A�O���`c	�54H�!��Cě���	+2�"�\!gyr5+��Ԧ�p<��p�ne��*A9B�Z����1<�\8q�b��\�:�ޒ���[��	�( �b��;��@��I�IEK�gB�1��2P�]�ꅆ�)�1��[%�|��P��3��Ň��Vg�f�J$o5�;"�A
[(�rM�.'g�'�p4P�ly����O�˧�,a����@Y'�ݷi�zA�&H�,T����?�KZ�#d"��W�� ��16��a���Sd����"��!`��愸�t����	�0h		��ܾ;e"|��ܥ�M���� !����&��ug��.�f)�tB��N^��Ҥ��I�y����Sd�)�OT:��t�Մb�0Q�4��{�C�	�O�zy+��Ь?sҼ���LN����$�v�'�N(!���5^��s�̞%� ���d�����O.�$D��>����O����Ob�4�����f�=��ᛵ:��E@ 7
��	���D�0W^`c>�O$4A��˓h��Y���_�jӄ��
dn����zj�6�([�6�a��#�ĳiъ�C�w��y�h�0>����W�̌2u��ȅ�̍2q��L>��׼Zp�@����6��xI�!EU�<�ͽT����h�8 �x1s��L~��.��|
J>��%��ْ꛶BE��VS�4-I%fƬ�?���?9��*���O&��p>�Iw�Pk"|�F�M1MF���Q-;���)��XPڐC��rx��P��9U�=+%j�0����O�T3�sF��{�F�A��3}���xf`��KU�:�I8e�Xh�"��C�}:��@
"m|` 1�O���IZ���@��\�`Y�@ō*{��B�	�@u�b��\Ȁ��r��d@�b�h ݴ����!�i���'<DzD��-Hb�p�f��$Q����'����d��'�iG6~��:�S�4N|;�爸qAR|�3��)hlq`��������~�'z��``k_8�|h�	+2��I_"g�5�a�6N�M�UD��:%zr���x�r�|��?��x.!B	��:dGȸY?�E{�eK=�y��4]�2��%�� UҊx�vKU�O~�=�'_�v"���:�
J�>rP!�O�&�'�&%P/o�X�d�O�˧��h�ä́T(�a_*�"�8��B[0�B���?!�ϖ�l8���:V�\�Y�g_�����m�D���k8@`E%P�㏓��	}D6�� ��c��S¦�xZ�9�eA��3�f���C�Z3��-Q.��g�u��)P|��\1�k3���T89�B���	�imNx�2d�/~�!�$��ZY��ĆnS�W�cfI��i>II���S,��'��=
M����B[G���m�<��ß,a�&W�X۬t�I韴��֟�t��,*�EP?(���W�@���S;%���pW'�O��911��'���P��1V��$a�<d��䃁- (Z4�ÖiC�_�\��(A��Īs�|z���>���]�0�����Hat����R3[z�K>��R��>�O0M�����k���X���|�-� "OlaY�$n߂M��1���W���`��4�,�O�H� �0j���.q~:�s����kan%���Y:��O����O�y�;�?����Y�7�H��B&\�8*X]Qq�O�LLY�O����!`؝3v&p��	���dЃLS8cl�:w���D� �0A.�
������E�R�8��Ѧ�@]�C�T�x��Ή�c�vI�0I�T��Q�,j˔���@؟�8�Lř%o�s�#�^M���'�8D�tB"k)-�T 
Ӫ��V��)�+�I9�M;J>�� �&~S���'�RnѼK�H��܋M;p8�̌)s���'�R@��'��=�r�U/�/_^��1K�2c��u�fY9#MT�C�'��1���A�⓹nkr�?i����pĆHb�ō�y�������#�(T�G>J�ⶃ<f���ٴ3"8�`���Uܓ�n ����ēD*|� pl� f�|b	< D�܅�S�? J�"���75�H���Q7*�6u�PO�\m�T��3�I�E�ĸXL�%b�%��tʙ��M;���?�,��4`0��Opi��*B�!�`�:bN(�-i�L�O��D?�<��c/>����ƈ��@ �OT���`�RH;&����/$E�'��j��R�~ʨ[��ۗ*0��a��,ȧ�\���)�i�D���or!�%�GKN(!J�3�B��I'��S�'"w�İ�ؗ]�`]H'�X%v�`q�ȓ.，jA��Cڠ�d�*J���ቴ�HO�D(!��0���!nQ:)��23FĦ���ڟ�IaWv�V�\Ο�����T�i����=g���eH=s��Q���2<���`@J�n�a� !AS�`�|�K<��mJ3_��\q�Fӣ
?"���J�� �V�ǝ~�˃�ܼlp�tq�+�o��m�V �2�&\Zf��::�<�p&��h�.i��d���x/O2Hcg�����Oj�O1�D�xF<4���ЦT!�D�/�l�8V�{�d�����2P��ɑ�HO�i�O�z�.,�5(T�+$h��_�{�u�T`	QB����?9���?1%�����ON�lVJ��"
?8�:tj�J�(, �D�$F��2~h��J�:�M;�������4�DE�2�l"��Lur1N�4�����G�Ⱥ�iBd �cJ�"5ӏ�`�'2����I$a��\�BN���� ���?)��iB�6�2����O��;��,D�f 	@g\6J��e��	_�	i��,�'b��z�AV&T*h��b��!�4�?�(O$�QlϦ��	ן�JÎ�,%6�c%a��`�\�F̞矌�	�2�L��	���ϧ$J��)3�зS��tJЦ�����⊒L  �SnU/-�*욣� ]E�����/ʓ[ $�h�4��x��Nj$Fh
�‷/o  Rb��+Nf����<GC���/ʓ���N�i��8�!� N�\$�ga�2" �	�'D̍��H��.� �q��D�S��:�'�26_3w���CG�����x��S7[�O�HxŪƦ��	֟(�O`�E�"�'b�j��G� $��� Q�|�0�!�'�B#Ћl���49w�-۠
�]R���'��K��S�d�eC���k>�hb��\(c�'����Ǥ
1gX�l�$B%>�`[�Jw%�(�OB�0�ϋ(tY��	ŧG:iK�@O�Dq
�O8�'��?E�H�z�PucQ�Q�1��X�#c0D�\#p`ċ'�P��I=�@��2O��Fz��]�-�F�B J��B*<�B�[�`�7��O����Oa����	Q^
��O����O��F�4&�$!HdݶT���>W��K"�Up �ѕJ��v��)�p�&�@�I7DXȀ�HN&����c�]$K���rO�C��Ah�,� ճ��+�M�I0᠈�1�� _H8��dM�8u�^��<�$M����>�OB��#ו��TFȘ�Ec��Q�"Ot�����7w�y b<*�K䘟��4�D�O�x����b��T��&�F�'nRI�X�wf�O����O���Ǻ���?�OB���w��!M�n���ԩ52��ǐ4N����'�R��9+ �'�>-��c
�N�س�Ϙ� �C4�T�۲��-}�ח�e/0@�+
?a�t��E_�1Oz�U�D�(��]vI��`a	%k�+A��'����W-<7�I�u"���:�	�' ~=㗈�d�(��1�O:A�届yZ�c�H2tE��M����?Q6,�cӮ5J@]�)�z��Δ�?���*�*����?��O�p�����<Ŕ]@R�NN�� �e���T,Hܩ�"O-�,��)g8��Y�!΃��5�1�N.���I'���P�-�a�>$�@ˇ< t����U�'P}+�C�'�x�E��6Qp,�����r�'0��MJ8+l�:׆�?}���2�'��6�;SqL	�IN�0߼��%���O��a��ͦ]���8�O��ђg�'�|8�7�Оu�T٩�o�����'C��]�\/ q�(FԒ��6A]�O���'��I��𒀃���z����(��6x`e�	�4iq&��`��i`�t0r�U��Ju:V�.�u�ԪDϰ���-�_eHX�u�ޑ�������}�)��5V@��&�Z�p91ŅG&�2C��,,7��Q�`��- I�0� F����$PU�'ЦA�vBέxN�u �ꅦ�<��Lz�Z��O���Q?0Xhx���O��$�O>�4���uB�$f�)jt ��mQ�E�Oon���]�Fr�)�M��$d�b>����
�<���q� /n�Z�s�����P� �q��l�h˷���a�C���']A�M`w�1�a�V�+4ʤ�&.��YD�J���-����)�3�d 
�^,��' m�a�u@I!T!��Y�K{�1�n�j�,x�ro�wS�	��HO��"�I�y42ź�K(20i��0 �Xճ�`�D�����OD���O��;�?���?i�+K��`�2��BִpPǚ�D,�BR�J�#���#� 0�yro��m��8���v��BB	)IhDΐ�)b"])LL�Jr�R�'ܜ}��%�2`IܓA�<�NX�T*�E�T�$D�F�y7�ޟqݴ@p�&�'u�I۟��?��˥'�<�j�&J` ��4�J�?	���?q��D<�� �Y�v�����0c�#0bw���%%>�d�6Jw��m]y"�03ϴ������	�c�&Ah��M��\b�HY_�h��	���P�� �l���|Rp@ҟt&��
p F�PL�B�.�h����)O��s�d�z�l1��CB�%���	�(^�x�̛�?q��x���@���-MP"�2�R��y�"�*|�xqsw�X�Hi��p�g���xR�p�^)z�F��7r�q��E6��L�S�5���^��Hl韘��]�tH# ��'ҏv���t�O�3��5�աu��'v�X0�I�挂P��=+�X	��τg����|b��:� }k@nN1#�D3V-�F�d�T"扈�jV�+-�B��od��~��OmqZgCZ+�2`��J+O��$�O�x����Ob��?��7L�:~���د7@�mxe�;D�L6!*Ϙ�FմP
V���;O�TGz��˗�L)Y�$It��;�d-e��6��O6�D�OByB�%P4<�D�O(�$�O�6�X��O'�zp��ʄ-<�&�co+?لŘ[/P��|&�X��o)=�s�߽vb���g�-��ĉ��WEz� E�Iuv�>�Z���~��A�|װ��1�]&>ɖ\��難Zq�O�Lã�����l��U;F�E,u���$Ewp�M0D�$P�e�X�y��jM=w\�\�a!?	��i>�'�@a�l�*`]U���8|�ʱ��I��z�f(A 
ş����������u��'�">�d!��HO�-mP��&͜3�P|uBȥk��D�#�	�E<t8��H;kF\�?����Q��
+���}�Dɔ"X7Td���+c㼽���ܳ}椭�޴5� ��v*RkܓR�LŒ-��!� ��n�4m�~a[u�O�<
����T�-��LYe
ʮH�x���X6�H$'&��t��J��u�$�<b�i2�'v�`1��j�p���Od���M��ɕ�΀"�}�� �O���G*#L��$�O���4!���/��L�q�!S��Y�6hT�u��t��x����'��J�J�8p�(�-�j&*	�Ǔ
��%�I3�ēE%�S��/IG��A��W�	�ȓD��E+o��K�F�(eN�=�����;��B�ܰ�k�"ԝ_����dNП��'7⥐�op��$�O��'K �S�����b#�L�N	T�R��F�4���?i�X5wz���Q��*��|�(���4.�+����M�)xࠀ�G�>)Ť�+S�$� �
��r��E ^-BEq� ���n�Z��$N@ ����>Q�I���d�<�:���
r��� �]:7l�l��C�s�<�G�3Z�*L�̠M��q�`Ws�,ي�d��� �(7�Օo�n4Ӆ��`<>�l�柀�I ��'¿w�ri���\�	���2�LI�daX�>�SrJE,�$,�<i��Hux�ѵ�ޅOC����S�NJ���`�?/���DB#��%�.B�bN��bEa��1&��2���Oq��'k$d���L��i�g�������'���q.D�!L�ᱵlKl���#�Of�Dz����3PДKs���U2��ݸc+�%�!QK2���O��d�O萯;�?Q���䌊�F�rp�I*���3gc��U �=X
�'[�sC�l{-(�WJ	6D�U b��?�x2h�_ޮ�J������X���BQa�$�]�D\f�	"V$S��A4�y§�)8�8��ՋĄ$Dd@��B�'��c�����)�M#��?���
�$UJ�@A�q\�q!�G8�?���J��!A��?1�O�������v��@[��ׁ>��dQ�,!�,��Ƀik2���a�%sZ�t����\���0�$O�y���'>rO޼��l�qN����H1FUbQ"O+FI����Q��'���	O��lڪk�����N@,vH��Q�����b�dz��8�M���?i,��,����OP5���)���4�;n�༢ģ�O �D5|f,�
�1��S�W>!��O� 4����a�#e�ldxԉ9}2.�}�n��c.>��	�>0v9��C�z.�:e"�rT�0���I��MC���d���B|����
�{E�Л�a
���'Q�'���Ad`я� �r��H<�P�
Ó|t��H�O6 � |���P�el<E��ͭ�M����?y��(n(������?����?	�׿��Z
ټ��0��DH�2�Ƽ��'D���	ϓr!���W!o�a����^�=y���\x���c�&}����#��Szp}Sfc�{�P~pm�)�3�d�2hv�E�7	�̦��gT\!�C�L\�\A�-�@id��#^'sH��!�HO>� �$�C!RI.Z�r�9o�$��-pQ��j���O��d�O(�ߺ;���?Y�O���&�ٝ6�Đ	q�C������fD��xR	ԆS�����N�8�� gҫB�$y�'�A R�F)M���0@�y�/�(�?I��'I0���ц&����Q�BP�j�'��lHU�קS@�1��:�f��y�+�ɹSuT ��4�?!��_Lpk1��<�B(�c��#+�d�����?!���?�����Dn�p`�� ���üY���,(�l(��`��?��I��N��X�&Fc�'L��ې+�3���0�H�/�l�Kg�O~X�A�Pˑ
�f��gÞD�џ|)!�OГO�9(��
�$�"����F��c"O� ���
:�Q�ф�G�jŊcO�oZ1	�>,)��9���*g�؁V�6b��c����Ms���?,�������O�����Ѵc+~���L\n��x+v �O��䕉O���)�|�'ol����gM�(���s�8I�J�(��`!�S�' ��7`�, s��\4>����OV< ��'`P�O�&iS��R0Wl�j3ˌZ�"���"OС�#b�:H��p靉1�j�P��'�*"=�W��2�,�'O
Y{���U�<�U꒑;���K�(�����O�<��)5N Ab䖷5yTx:�n�L�<�֣ 9�65*p�ȯ��X�$n�I�<��g����b7�Y�<,�a�&HA�<q4��t�,9��J�|��o�{�<��Ɲ  ^��W�֬n�:}�D't�<��e�}~̍
fD߫Q٠A)@�s�<�%��D~�m��I�Yg ����l�<4�ڴK4�M�!��Ix	*�No�<YU LD]r��D�Y�D����Rn�<��oOal	����.���B��h�<�"�V}�$�s����	0�a�<i���~`�Jq(QN�>)c�*D�tX���:T�����p).��''.D��1�G�;z�҄$�.*Ce�>D���\<gԕZ�L�L�\@d�<D� ��Č({����H�.Of�$M%D�DY@_W�l�"d����H�)9D��2�e�{1�Z��>	=Z�C�7D�{R ��4y�(�C�M<�<��8D������b�� ���
��K&�+D����; �*o�YP�4��)D�t��
���hZ�-���UE;D�`�a"��>�����8�z̸�B4D���qcX����e��`y�=2!�$D���$�V�q�>l{Q�_Ԕ%��.$D��CM+�*��cHQ؀��s�!D������8r;�M3�lia�K,D�`WD��y�^���O�.ouPu҃�)D�T��&�{��� c��G�6Q��'D�D ��"� ��%�\4�q�9D�p�����/;���s�@�H� )1+�O�Y����{w�D�R3��=	�%�6:J�;�&x�~�z���:�H������#�h�c���HO�H#�����3��h�(I�n�B�Hrϱ*oj訄����<�S�.B�Jv ߑj�j骀���H��@X?xa�8�Gָl:�XG�d�N���'��#!}�����=�uO�X�Go_�E�<�#���t��Z�A�>��ܸ'���vi<����Kw���m��:Π�0&�@�x�dH�����qZ�Ȩ��*#"Պ�B�4�O�Ol��"�u`����_h�#H<��G;(?8�`C��7bV%��<�	;eE�)`�a�Xq�H+�ϔ"!Ŗ�Q�"��R>��c��d��5�:D���"�H�A��I�C��à�Ey�'1�� �xޙHbdD�v���H�m��Z��礒�d�Fj���I�4��pH�*�|�@��o۔��O�l��Ȏ�)�*4�HE6y��v�>14�V[N����B�e|x#m�Y?q�Nȿv�c`�:?��O��-!���(��C#Y�FK���U�
<)3L�3�ORB��R��H�e��	'�j�V�X�ex�͔���O8p(�֞P�숹��cw�94���l��Ǟ���P3�ʳ8�?�!h_�{��$�v��n���i��Y�b�@j���O�SW�? \t��*�bQ~�j��^�����T�<&r+�ǉ&����]�w<��Aå��*�LɊ&�D�V�l@+c/B9R�phJ�Ǖ�(�Nui���|`k�/#�;	�~y�*[����� 7V4b���4��5Mn$����C�,���!�B2�[6D�����Q0K��c�\?8�D��E�X: �����?Yx���={d����%�	g��� �޻OP�$bMK��%�q��K��� �_P�p���)�	@6)�p�3 �"PB��!E
�5�' �Q�G�,��"�.8�@��?�%$ծ`�j�d�rv�l��J\��O^�����埄7-�3J���gO�xQB@G9�5��J���r�?��?ySJP/F��H�&�H0��#�R=:�� �>iӈjF�4��?1G�TE�t@��R��ڄ
��7!E.��'�LJ��\59�� ��CA�*�:c��@%j�:|�Î�'���b䈭<y��>��?�!��n48`
��}Ь�#�G��|R�+�1���S�ʞ{20�x�!�e8�{fпr[^D��H��bM�fn���'Ө�GiM��l{m
`�f@q�b��w��a
5��0N.H�ȓv� ,�TO�d@�e��8N܀i3҂��EĀ�(O�d��-x�܁ϻR���V�K�m"�=C��&3H��'��~B��6 �쥢�g�$��]a�)� ��'�4���-�<�IAU�\�Oh*d�L2>Q8�k�:�1���xr���>�1�W���C�HCCn�3Q�OpB�����e� #��S��#J^yR
<�$�b�ɹb`��j�Ğ�X�!G�1g��;��5q���)NN�v�Q�,s���/
����,[8Eqf�h��8
����O�S� �����@ҷ ��P�D�F6{R�	����?�$|	��	�jEc�/u�-�u��Q\�`F
�1$`�ȶ�����������?mI�N426R(��J"xF`�D�>�,��ٖ��(�l�R���p��'o��ځ��bO���Ѡ�2 R��'4�y�dzz5�Q�%�@�8�����]A�ϱU<d��]z������5$��Y�K�1x0�4�BL(�qO�Y��`�DJ&2��N��j�)��ͮ<�2G QJ2��� {�X ����l�'!�(��D	4U~��I���(eйA����'h�!�{�S����5C"��((8M@���j\1 j�	R�D}�a ,��w.lӶ��UI��f��>��}��V-+8�"}��O�t�K�%��ievD誏�Ğ(u����c��4(��D��I� �H!P�P��r�1�i(���'�h��bR���#@�e�I�=$�K5�I.�-��c�%76%��&ј��%��Ȃ{��]p�iCz�qO�Y���f��Uv�Y�f��y/�ӑκ<bś��2�GW+��[�i�}�' �|{��˪#$�]FF=��΁3@�<��_]&�C �^&Mp�a��@���m��m�D�d� O.�/5i4��Ƽ��W,Wں훅��+]1�9��,�D��L��G�QL�E-�U;Zd��V�z�
Fyb�@���A%�<�Ze��F���A$2�lxЅW8s��1)2)K�EX��@�Unӣn<�c�Y�	�J,��(b�,X��9'��F��e[�i˞#r�� "���q�`�,k�X ,O�c�� v]t4��cð�2����馫�?uP>���n�����	 ����S��<3�����ө䲩P�!�~���j؞���/�,l��� g�.iB�@A�(}~����.�O8��u
��y�eCj��-M5wTйh��$�p=I/O�M0�mS!L�h@�ƊmY����F�{���I��^
O�5�޴-٦���V�;%��B�����Hfl�ɒ$�^~:���<� T�l w��y��#�it*��UET��@ꔤ��3i�%06��,8�i��)tӒ�pv.�ĸ�����J���rA�$�n��)�6��-?/$�j��Ć���Dк���0tU�ah�YC��n����K(A'�'�Htp�LB"z5rY�FC^�9�4�޴NN�HJ@�6O�{���?A�.X�]��E��
�;ĆUɶM�g؞��p�ȐjY��)Z8c�O
��ƌ�����#=��`��T���}B���&��w]���C"�a�.����g =��׎<1�#��i� �q1��mڱgF@��t��s�<�`��sSv��0�1<��|����Lƀ�@ʊ�Y���K����#&�� K� �8�\�-OX���	8,��[�⑼'󐜚BD3Jֶ7"4�P=��b�P���� �#7)��J5�5{R�U��( �'M�	�B� �!3��|����&�T��q�"U������KY
xz�'3����d�>���ǩg{B1'K:{2��ğG���$��O�� j^�4vd)
�C�Ox2˔0�0M�f�Y�%'>� .��M3�	�)P�<���ԧw���c�b�Iy��$߃M�<��
�^��9ؔiJ�,���� ��P�ц��eK��Q�f�ў I�#޸�D�W��V2\(2Pe�T�⌅�	�5O�}�c$�W"m����-4�Y�ϧz��B��d�7D��j�9�� \�ѳ*�*m��#�T�,� ��'�\�ӷ�-Y��i�� 3�buӆa�g������/2���l�@���3?����gh>�i��_��*�K�[�'���� �I(�~�c�@�D,���yLH���F�(��)��NY�<�zቔϔ$�he����"^l��w�ԟ�	�/ې`K�~\�҂�3ʓm��!jte[+n��		���$�Fy�aV��֔�1�AR�X !��f$ٌ{҃��?�O�P�;T�[�hQ�UːJքB���% ՜��t�mHU�'2&8�G�̼#b�/V:u(tJX,dYTLr�	"F��`���)�Z�-ջ:8N��ҬS/	ܰ��l�'`V���nK�7�p��ѭI���c�OR��3�Y(���*����\�R��OB�R�'&��$��T�&�츠�HY�S�&����G:V�69pE�,E 4iO�:�x�a�`��C�t̠UP�fqT���>���߄l������´���_y��3;�|
׮S��`-�3���(OF�	V'��z�m�E`N�^>�&gԺ �qO� �_����	��'St�ȢjD~r����ƅ<� �y6MW�l*F�����o�\i6P�Y�$.��B�탵��X`��8A����'_,�q�4O���Ğ�?��E��<K�a�«�\J@��"�?��D�a�� -9�0�p�G)09��n�����B.�UA�];m�<����T��&D���i�H�i���F]2��%%&
��1)��<6�kժ(](L�HC��%:���h��-
�Ё�į��dH�%#ڴ)F:3�R�,O��G�)�H
EĒ>N��E�	&T�	1��>f�|5���ԁ�(O�8{rla�����Be�	�q�iώ��#H0�@�U�Ly���Okl�8'�&(�V'ڂve���ҩl@F�q�`�*��,jS�i�!�@�Y��]9x
u(�(Q�7�24�󣙄E������ ��Q�?��,�v�<�w!d�AI��h:;5��=}��m�>9uG�:�܄�%oz�ɹ:���"�<Y��xAG#;X^x�歖0-�R@�6O�Tt�x�͋�B��I��]�P� ��
E /�@B����H����*� QD-D?iU��vW�)���2J�����p�
�=ܴ�%LI!��r��U(s��06��
 v0qъ"�ڲbQ�u��o� ��YzQ�_��M[T(B�N�|���&ko*�i��s��I�ڴs7 D�9��6aY)Mt\ :sR4@�J���h���(O�4iI	�\̻~E��� ��01��Z>�����o@-/lh	�J<��
Ž����i�I*C�d<���P �X���%+�	V:~t�&�,I���L��0`��O�LZ�����Ey�AF�Ҍ �ZM��B�`7h�X�� �,"<ͧY�ִ��G�,An�B�D"P��}ӆ�4t�Р���3��  �"�q�hqKG�-*���7!.�*ŏS*Z��O{�dzb�{��&����I<a \]�F03�k_�oB��e�'�	3W˘TI�%Z�}��d��ê~sD0q��A�t"���E�o~���3O4��YI@	}��/	�����@鐵DĐ����^��Fy��T���D�`ޥK�i�;�I%�ԛF���#�H������q�ȝ(��	9����
2��.6fՋ��\�}�2e�F�]��,}ԩ�l@�G�lͨe�d{�d��C�*[���{� �!J"e;D��?3d\J�۝p�0� B�TJb�(�'?�ɺ���{a�c0�E.(�Hd��
%�1ʑ ������`�V)3��A�D���.$䲈
Tm�"c;���W9���fh�5w" cPbZ�v�~�R�mV\�t/F���kS��e.�ӊ�d�.+[6c
8Z�h3⋍1	h&����Es&�r�!�&�X���}nZ�h٤��)>c�X���&=���E�!r�1��5�ӺC��]$V�4y�;`)zb��%���qc��\�n �� 8`!XP� �j����^Q��}�O����R"~��4+T �!k�&��}b�J�I���!k��
	���֤@!�M�0������3��/�<]�+�TMfe.�6Q2��y<\��ԟ�!H�lF�I�6P0�$^-���7FI-h�� ]�_\�����
8�uӆ�	����>���1JQ'M����K~b��ȒG��!��I/SLf�a�*�y�	�&��`ǀE�3l�[���W�O�	�'�	r���T�B�bVnX�H���?�"cAMU��)d�| ��)��Zc�����Q�B�
��
�e���p�N,O;�*���; ����qJ(Q9��
 ���򕦌�~ �i��I�b����.�𑮜�>��k��8	�t���9�QLL�&�~����
1�OzX#��tQ#$)��_E�Ei�����='���	�e�0�P(Z)���$��aB@�@�`�8��qt�9��"�dc�Ai`Y@�7Ny���1��,��$,�pۂ�/N�|��qwʄ(sA��g��M+1F�v�(X��H�VDڦ&�j�R���-�
�\���_SHB����(��q�pȗz5���ȓ)��E[ǁ�2���1aَ�X��ȓe�� �.@�v��(Å�	6�Ʌ�K&��;���}��芐���+S&���v��S#*�6��q��N�������hA
��E?6!�*L�n�Q��)���;L�=w�}�ŭ�:�:͆�7�^e˵��f2J5� �g1v9��S�? ��h��*�T1����%�| �"O"42riT�r1
W���h�V�!7"O@�cf��7 xZ�*��@�s�.0��"O�HX�.�4\C�����]�z�^LAE"O���O�0al�iV閌JH�@�"O~ʃ��Q�V���;_BB�y�"OTK�`�J����B�Ǘ*�p�"O�9R�Ơx�\����%G8���r"O�Thn��xԤ���޺P#��q"ObP$�͚'̒�Ip�\��jd"O� �C'��)(
�K�ʊ��`'"OX��!K�e�E�)�Y��0�"O�3�N_	1��ը�gV+f�ԥ��"O�I��d�+�:��f[�;K�"O8�A��02�PA@Eݚ>���s"O�0܏e��	 �E�20���"O�!��X� $8l2$��6&
`�"O�qs*�4������x�"OP�t�N�LК��&`0���i�"O^k���Z�u���,L��у "O��r���S���B��ӝ	�
q��"O ص( 7�݉���9�`��"O�}r�+�_Z���D�޻a���Y�"O���ˏj��� �逆j���A"O�Qc��hk$Uyb�T,ps�9AT"O�<�N�z��}�Gg�q�f�S "O�� �s[�zׄѾS�n8�"O>����O�ulI�G��W�~P�"O�����F� ��$��Sx����"O��J��[�Z��b��=$�|8a�"O�(�*��>��Y�oP��*��"O@���/{�홱�F�-�>A&"O�%-Ĵyi@�!��ĉ~0^�"O�h;RcdLYK�$��/#���"O��I��ϛ�l���7�bs"O&�)�	I��
���@J�,��"O�� �A2& ����йA8j!# "O:�J���+_�V� �
��h	�"O��8��#V'^�ʅ��V!H8�"OR�H�#��~���r�EC$ ���"O�$��i�K�šq��9�U"O>����|�c�3F�x[p"O@� a����u�����`"O }�d�V.H����!��cbD5[�"O�� ��x\�p�Q҆|S>��`"O�t�g�'`�fD*��-Y@��E"O�!P�F͋-��X0�8k�  �w"O�h5"��4������{�"OV��� ��\:���#$��(��"O�x#$T%;�@k�dٖ���"O\ "`f�[����.ڂ:�P1"�"O�$'=y ���MAB�|ɨ4"O2���)C���2l��[��c"O*!���C4d$h�M�D����"Ol5��kK�k�9�7�N�f����"O�Ix�.���H����J�"O����e�g(����l�w�6h3"O��x��թ+�H��?~����"O*as�J׀H���@6�K;���7�I��YG��jŴOv`6��O�p�WG_V!��E��qz��� �ay���)<!�$�0�����䀂J�H����  i�!�dX:T*l�ei� ��]�ÃQ����u����+�G��#dN�4Q���'aVӧ� �(i��#@Y����!��X��IY8�4�lWhy��v���G�Y8T�+D�����Z=T���*�6f���G�'D��Q�]]��3d�U ��I���#��-�S�,�J����E�G������h�VՅ�+F�ٺ��)��:э�.nE���Si����HE?/ު\BwhC(7�|��ȓ^t;Q�+�`��&̜�7���'*�"=E���A[�4�2�ʧ#E�!ёU���$�Iv>-�w����Xd���u�\㟔��Imh�I"��RP 8r�ީ��B��9/�h �ԯT/D)4��
�l�vB䉎=c�T`a ��F�����d�#$���$M�Cf��C`��=���27�e�D���٠[� `p�7 �~y#��=�y��V3`�|{0���m~��R��M���sӴ�jQM��	6L,&2�m�"O����S�j���!��o�:@��'�Oh�H�#�b��D ���ԣu"OtݣW��TZ��ct�U�4F�"2"O:i*G��,.�U�F�z@�T"O���M�GŸ݋W���
����"O��˶�\c|�
��
�-�V���"O�)6�>Ҁъ��uq^Ik��Iz8��A����cq�!���ܶ4hf	ySm?D����G��xa*x�A&gL�Y a�vB�"B>=h��Ȁ/q�EW�΀H�C�	7^�`�r��܇Gt����M�T����$a�|���5��!!F꘼n�Rr�.D�h�Un��Ck ��v��I�<P��+��蟲M����9�y�j_P��"O���q� �V\'ȷ}�d���_��E{��I[1B&�1hV�,<S��i��P�����+���G��0�VU� �@�� Fxr�)���"ij̓E��3&?��XҭHb�<y�o�O#�e�`k1{9$]���]�<I�H�Va�]R�MN�9+F ��-�Y�<ɂ�8�� ���é�XtB��OX�<�TL�u��4��Y�4)�d��ă~�<I��P�&���U�=/|��V��a�<q�#�O�J)��IML[Zm�6˒I��y�~z"'	����;7o�0<��s`'D�*&,��ޕ�v�U-VYN���ؐx��C<،<�g�J�!������W��'��hEyJ~J��Ya)�6�� /�Ua�V;�y� ���t*��&φt#�����y���TA4$�"�UC�-�D�ֲ�yR�)!����7�ϵ>�Fdh$k���y��VJ5x����H9���u�Z��yB�̅>�-@ǉ�,��cT���y"�X����:�)S��yr���hB�Sf����C	�y�'��FF�m��7����H���%�OT%ӐND�9$��s1�&bVU "O| �E��/$�����CZ�P�"O8(#ÊƏ�}�d��WZx�!"O� %��g���f��7u��"O2�rCE��xFc\�[�)+'"O^ĩ��L�I��b'��N���G"O��X����fZ`-���9�t@T"O���D�=T�<���>Y-�h��'剃2{�Uj��#�~��vL�K�
B�	��dj'��3�}C'�_�f$C�I���aб$A�Z ���bܪ ��O:6-����� ��H�� j}��#�O);�����4�S��ެq�0�뚜+�~�ys�O�y�!��#'��=+���"vzn4Z���n��'���q~�>�d���E�2*���2��+>^95*O"�3 m��5_��NŘ�:�S�,�'����|%��k�X�Qqn�'c
��k��\�`)z@D}��O�#|�h��8v�ac��PbQ%��k~R�)§}@����*{[x���P�@̀�ڇ�)�� ���&�5Y�7:� B�9D�����^8'*���zo�aj e$���I]�'��-�7M[�B�ܭ9�鍼g.�h`���ΧB]���F�g���JE+<	!��Ķ�2����x`��P��!�R�z�4r�(�15s��B �#�!��AWoV���O/>���"���<f8D{���'`�Ci^*?���&���t2a
�4����=ѣ�еm��(xB-O4 ��@ ̃J}�'A�D�����i].�2�Jڊg�6\(�'�\A�QAǍ �p�9��/[sl4P��&<O.��rM�x~rd#bJâ) \��"Ol
�6pcV뚜��8jV@ �!!�$M4{�JM��^�)��)p�L�#!�սꒄ�4(���^A�5��?/!�D�3\�\d�U�f��!�!�܀�!�$��V��?�4���g�!򄜦s���8�.B������&>n!��N�Q°KT���h���S��!�DL����3�Y=[�VM
A�!�$�
��E���� >I��YV ϩBD{���'$ܔ)f��l��5��H�C���k�'#��rj�!W�����B9�����'e��
���%�6LaA�	�tS(O��D@���ER5��0D�O�wg�Iw����@�
�k>Jtc�O�k��Ö�	l���ͼl����uo9o��Em�1m둞XF{����hek[�}ZL��9P����U"O�H�BU�L���(ӕ7�DI�"O|��`�?��!���6t���'��OVD8+�SS�|�7J�|o�� "O"�`��DE�U�G�U�MKF��ԇ�	.jV ��Gl�z~����ȟq�C�	�E��\#�^5����B�x�0B�ɩiR����ԭ BZ@�+X�\�.B�IZ�:I"%�؆��m�`jV/B�TB䉦B3�1Qn̙��M��N�C4^��Dl� Aw����t��MZ�J���a�%D� �kY2q[�H�NW�e��pZ7M&D�cƬ�:"�~2�n(E�4+#�#D��!�Ä&1��cc�@.~��V�&D�X���	J vx����>Z2)3��!D�,{�FM1�|(լ�!���?D�#��^=~g����@���D�=D���Ee��;T�Er�	�Lŀ'�9D�����!ms�����ֽl)2�rb�:D���R/3� �2���#��p�g&7D�D��2hA���пM�􈚱 "D�l���nz�)"��`�X���%D���&A��_q�p��mU�]��� �#D��B�4P��c(�Q�4�uf>D���E��<�R �-h�Z`J2�=D������ `�6�Z�O��~m� !,<D�lq@��L���5ϊ+6@�PM:D��q�m�x���Ik�3:`�y dL;D���V+�o�8a[Po�
�~� �e-D�� h����,��@��O�B<��v"O�H�b�T1<��A�5�m*�',���p���e�Z�hՠyu���'xr] ��)=iV�:$W�r;P�	�'d�T�!)a�5ڃ�	kZj�0�'j���uJ�
�0�(�'j$��	�'������C0 ���x�(W�� j
�'�.�ħǷ;R��IE�˜S�|1�'2�hм! �r�'G4��]���y�ךo�唄}F|�H2��y���-v�1&����jF��y�n�5!"d�F�G�����Ĉ�y�P=2{��Wꓽ�5k�ˉ��yn(F�4��d�R&q���T�P��yB�� B�0Y ������MX�yҌ������O���F�!D��y�� P�Q ���$)��S�yH�9BjJ����Q6��8��L	�y�LU8m�v�3���ļ� a'؟�y�FÞK;�i����e����g ��y�7g����/�-x$�2R�ނ�y����`��"G��9����y�n�%g[�%HÌj/��x0&���y2�σ6�|�9��1�.�`�ۑ�y"B5$w�xj� [7	��'���y�*�U��T�F'��,�(�GG��y�Ɲ��M�����"�>d���1�'$J�6)��>�<�I2��:W��z
�'b��Rp�
-ex����&-rA	
�'�d<�d��Ul$� gM�W(H�
�'����cU�P+�M0GI�B�*
�'�Z�C!]�m����oY�O���s	�'�v\`3�	Yd�kIG�P����'*��K�͗U����N�6I�����'\H�q��ƒۣ͆�D!`��'����b�zp�`��[�Y�R��ȓ snq��G�6m,D%kѣ1E�(A��hʭhg�\9DЙyuNK*O�l�����	�ƈPm�,y$������	i���=bg�URfJ�1�X��E0�ٙ��ѩ|%FD2�D�EF�]����Aro4ikH�8S'��w�f���6+�A:u��eɎ������ȓf�iyS�
�b�N����ϗ��T��vk�Q�-SK6TX������ȓHjV-�'MѤ�iPV4b��0��j��1k�Lvz8�%Fky�%��b�^!�@mS^@h�K�So�e�ȓ׈-��M)A�>\�aK�!�u�ȓ ��!-Ț+%%#cC��$�,чȓ�D\����@W640��Cl�6i�d��	5Ć�{,S�aR͆�#���r�F[#[���ҏM	4����ȓA�����ӈh y�b �o>�ȓ�R��c�ȟP�" �M>$?¬��j��a&�b���ʠJҤm�.��k}�ҍ�t2�R��)p�9�ȓ��Pi�IY�:ʆq����dæA�ȓMS*4�1cC�4� A"�)S�d�ȓ!�Fͻm��9�pX�Bo�F�^4�ȓG��	2Ah�d)�)ʻ�Y�ȓ`�PE�P��&a����L,��|��\��`R���[v��FM�hT\��ȓ��i�e��D���j�V���S�? %!b��HZn�B�/"�a{u"Oa�W������%�G�S�v$*�"O���ʔ�/c*ԫ��[�LJ�X"O��qP�D���0B�W~Q�;�"O(EV�	�^�Tx#���n2�m�""O�(��Q�O�x�K!?+<aQ"O8dpS�E'	�X�����f�<���"OR��E�SJ<VѲ�kۚv�H �7"O� "�Y#C�dT��+��$�\e��"OJ�a��:S�21S'k� B�$+�"O>�2v���$��	���	 3$\��"O.��
� .��P��v����"O��8��W<�zЙ�c_!%fv-h0"O��+��͸U�;�kçev��{D"O�\���z����g���~i��"O���C͋+����7KK n�ZE��"O�p��Q�;T�yx�,1 t�[�"O��R��2+FRȒ�,\�kt��"O��S��I�
�dA��&F�l^�I""OiQb���x|SdC��>;����"O<��q�����:���3m�^D�"O���`H�E_� t���]�:�0�"O�}2���"0��Ti�+���"O
�XDJ�7g5�D�� +T�<�I�"OB\
�W�X�ʘ��Q�Ј�1q"O
]{��Q�@�H�֭�-Y�`��c"O�u7�(��tLX':�z᫃"O�U�OM�8.0u��aԅ#�"��0"O ����'`༺D!�.yԸL�#"O�1�D�E�s��e{�I���г"O�|�b3=���
>���"O,��Ū�<ϲ���ؒ �����"O"4r�	>k-�1`Hv��49�&D�4���>�z0B"��Rw�xJ��&D��21֎~�&��v�!I� �b1D���욐��R�G� q |)@�*D��Xbm�7[������/B�����)D��JW�O�5v�x��LB"��31�#D�D��L�
"]��$J�T����;D�,R�R�e�AA�?A� 0q`�9D�\a҅O�+�`Yw���i�\�4D�(r��^v,�L8"L��8�T�K�'D���ЯD�T<�u��'�ymp(;vj#D� ��G!����U*�z�\�a0�>D���b�Wq�	�4A�emp�1D�X�`��k�$�1�� ��}i�"-D��x"B	%ԑ��2`^��C�`,D�Y�$̦J҄���HR���S��*D�\	P�ɾR�b���F�Q�n${&l3D�4�Ud�m���p��Mv���/D� 	L-�ʱ�B�s���v#D�@��A�� ���]����y��$D�`���X{�Y�&)�ۊe���.D�\��%�/	��pv�_g�͢��?D�<��'��A��4ja�Y�.9C�=D�<21h��4����b�c�@<D�$��(]�!�@@��DN[vNm�'G:D�Ȃ����"PWd�1-�̠AB8D�T�dDɸ0�LtH�I� nHd��1."D����]�e�]z��PUn ��?D�� �
7W��h�sށw�"ᙗb*D�,��噉/_hA@b�Y�o����1�<D�9��.B($��D!G�x�`$7D��#�3AmƸv�Ҍ)��� o:D�� @�2��/O�Y�H_�~>$2�"O �p��;���i��@kA"O���� �:a,��_=��$y�"OV�r��!6��bvlW�T���"O�up�	ZT��e��l�w�6��"O�M�â�"Q�����-B�d����"O�CFE��6�,I"<0l��P�"O$XS�e�����2I��"O��#�@*G��x(�g�dei�"O`��	��"�df
�ilP���'҈�c�gSL�Q�,iT���'�D�{!�;Ѣq�䑰�JD��'o�i�������)�"K��l���'>0����	5�Mh��
�b���'���Um�&�� %ѨW��0��'��� V�$tw8���3G�f���']����c�Z�����CO�+E�I��'������̯intpKtaי'���'`���gZ?wߒu�$�-$�
|��'�$IS�ǽl\у�ܖ�@]Y�'�`	KR'�a�4��+�4�̍+�'��*��{.x��F�)B*%�'�\]S j	4���#$%	��b�'���5�ґu-�Y���P/ Ĵ���'��s�K[�
'�y�!jK�j��#�'���T�V���0��M�h�I�	�'�z�p�e��H�q2M�Y�'��S�/S�zzz-��e��[�4�X�'ۂ ��`�K�n�V0[`��9�'Հ]��AO6�wY �V�P�'v�4�]"�@g&�d��+�'�����K�!2�\421���͈`D3T���&�͝g ��)��K�P�^m�"O���dBR.��x��	6|�s5"Op�0C�[�(e�0�uLD5<�"O�����6��W�ë�ҁ)�"O�X2��ٯM�!@֊��4�LS"OPUsf	>X�p� JZ3��j�"O���%� �l���&�9p��MZ5"O�;wc�@Q�ȹc�E�r�"O�-C�"�%*�D"ȏ7B��@��"OH�	2�	?A
�-�0�	�"R"O�p��T
aG�E*��؛=p�ip�"O"�卒2 �0jW	�w| � "O����Ε*�y8t�	i2`c$"O����Lό
T:��R&T1Tu���d"OX�*�`�;.8�q�Rƅ�spƤi"OP1�ņ1V���%��K���q�"O�)c���S쾠𧦜�h�l$�$*O<�K���c��{�JA�Q]b	�'�D�A�d�x�hT�	=R����'G�A�
�d�ో/҃|p��'Dx@A c(N,q{c�s����'ST��� �F�Aqj~�����'��(��;FMH![�GݗB���'><���+
97}�г��7�HD�'�^U���?e슼AV�?�r�'A�����	�(�%&�[,��
�'Dh���*۹]T�35���v�5��'�$]�-�t@���	T�p�rhQ	�'�l���ڮN*�B�ۏa~��8	�'�"t�'�M6 Pڹy$�J5V�3	�'�h�����3zk���k�vR���'�zqp%ꌄm ���CV�Cm�Գ��� ���7@
$qp!s�k��A�f"O(IEI�3ol�PKմf� �
"O0�0Ҫ�C϶���K=m��y�"Ox ���>QF�h�L rF��#�"O���\ 8v����34��Z�"O�L����!s&A��C�#d=��"O�����N�͌�2��A�H�xD"O�EJ�'[M.�{�aɄy� �:�"O<�c��J�GL���"G_��%�"O,��D�$�zX����贕�f"Oz�1t��3 �b��aC%yA4i�"O��gKCii�`�U�#�x��"Ov�6CѮ|T���m�D�����"O4�i��^�|�Y�m��#��RF"O��{&�O�R88+�LD4�����"O�|p�]�Gs$��Ѥ�*�$ �"O�����8]ے#�Ev�g"O�-�Q�-{�ٹ��s.\]y�"O�Ej�iL\�
��֮�}- ���"OB���I��x�����Hi��"ORQ��mF
93
�e6Nz���"O dp���=���I�����f"O>��ީ0pL��l�d���5"OT�su�W.K�*��5a��%���@"OV<�A%�,G����э~Ċhҧ"ODQ���";H���G�D�NU8p"O��Fd�w��J�	��t:.��"O��i�G�NRt�bb/�.��"O<�hSPla�<��c��7͚@��"O���#� h�����dڨ* l|��"O4pؠ � Xpl� ���1;�"O��r��32���j�J0��d"OFPZ�	�\,�[O :��c�"O���d@�Y��Sԥ�[�: `"OPj��iNZ�
P��3W�P`t"O,�w'ڑt�i�׃������"O��RjQ�R+�컄�^{�dī�"O���'K�qBj��Cc�݋�+�y2�D!'�sW��(p���a�ޑ�yR�� ~.�:'�ރ�5@p�=�yK�0c6P���GH��W�(�y�NX�2�ճ�n�`���#�o��yr�Ҧ��Q��OH�A��d���y�*U�1r�9b�Aw���;�a ��y2�\٨؀t�CrOvU�p���yҭ��.�����IfwZ����E�yrL[�z�8X�f��,��=8W���y2��=}*��h_�(G2����y����Z�4@�b�� 2	*$�R�ƾ�yƗ�@=����G��yV��0O��y2�T:L���c"��V9�VC̒�y�=j�q��D�1�&m���G��y��ˮ}<4XȂ蜰#�`���yr җP<TQ���� tH!!S��yH6���  ��
n����y�8$�XB���A,����y�l_�C���+3�_t%vL��@.�y��Ϭm��d�di\��U���1�y� #v��cKؓ#z�c��5�y2�׍%���҄(�>.Tŉb���y��׫S-�X�v�Ń|�2��B�y��	n���B1�I�)�M(4����y�� "ČӢ�S� PT�)`�yB�^���A��k�|lAG�["�y
� $��%�JZ �)f�!:��x�"O�hXq��/1�p��IA®���"Ox�;����v��MX�Fߐ[���k"O����l֙��;ѓ^��\AE"O��cG��>b_h�A ��D�u��"O�%A��vZ	��I�@�$0a"OH��F�Q+<kd4�F)�r�VX�"O���Č��~��.	�xT�v/̼�yRI��T�xYx gŔq}�DHV�G��y����H�� KV��-�Tõ�S?�y�·�U�Ɲ�E���.,��
�%�y��FUƘ�7%F>P8n1h��G��y�݄#�"d2���,Kˢ<��FZ��y�`��l��v	�?��I���%�y"�S�Q��c�MB�F&R})FJY_�<��mQ��`vkf{p��g�r�<AD18V^ظ��Y?��M9cFF�<�q��?#��(���X61:v��
��<q	V�.D�����J�,:%�T�<	�e×>/��B@��o�HEh�NX�<1vA��� �bs'Ҵg�����m�<Qc�W"c�Щ&S�9AR)rEDUR�<��!�ZNL��@J|���ňd�<Y�H�OQ`�DG�ƈ���X`�<!C$��]c�#�h��O������C�<���R<�sBӜx�)�p��}�<���Z.���E�G?b��)!�m�y�<9�N��$���7
 t^��Ms�<	1��+g���I0/���� Ʃ�q�<���bn����I۵u�0���x�<�֤�>YYH`��̱XW��b�!���^���qQ�^1`�4���ɔK�!�N�0����!b�"<b�e	��59�!�[�Ob�[�GԊ>f@�Ao˱0�!��:�n���ؔ`�b���֘Y!��,gYf��-ԅ	��u#0c+G=!�$1_8蕱"��)1��v��!�$�(��TK��>L�%;eb��&�!�D�-
�t%��'Q4@Ԙ��� �!�q��AQ��t+֬�&%V�^�!�D�iH�NuD��R��q�!��&t�abʹn�@�a��N�!�DY�>�ف�������t*u�!�Ć�_0��
4�n,�����!�V:���Wf�-�e�U���!�D�>���y���|Un��0J!���L�PQ1k�
,T��IW�ȝ]�!��ē?�@�Z���*ԥ;�!�J�h�P��l�+�"1���L$7z!��\�@&����Rq�X�4 �:k�!����@	�"�$� ��̑l�!�����'���0O3s�!�DֶQ��`����ic`N�h(!�dW����b0�Ȭ9���	}6!�dO�r�ą�Qؖ'�@�G��R{!�䐽�(ؓ�N�J���q�&�g�!�䎖@�<��gT�h�H�9ťB1f!��Vld�m�0:�zi�d�!^!�'$`)��o׊d��q���)0E!�d�Y�ih 
	���1�@�YA!�d��̖�`�]�V�v0*��D�c*!�� 9��2�O�~RP� f�=R!� Q�NH�7�T�HFz`���۲!��YL����*��_׾qq���b�!�� ޽���Z�qMN�y��0t"O(�:��6x���a�z���"OZ�Q`$A�1�
��á {Z��"OZ�����
F(�Թ  � Y��"O��a@)C�{t��B��SI�٢�"O�be�K)b�
P�T��v���
�'�:y�埓��ȣϞF�B�a�'|�h��W��b���>82�'�<˲,B5"�@�E��?3��E)�'JD3�-��� 4*_�-}ƽ��'�4����H�sԭhӆ��KX��'�H�����%7� RLX�¾��	�'��M�"{����G�ƶuj���"O��B�4F���O�k�&��"O��w��G]��rnB
-�X�"OD��6�՚4�^]z�,@��VL��"O�UB�*(8�&X�l=�%"O��@�BI�f
%�r���XiW"O�Y( 

df�h�DPwꔃ�"O�p{T*�ud�܈q%�2H��Hg"O����MZ\  �U9#��I�D"O��т8,�r]�E ��d�z$c�"O�%1�Úl\k6 �15�� �f"O@hs�D�46F�0����lޘ��"Obu�a��=*rej�(��*u~(��"O
)тCG5O���H�. l�Lq0"O���J+���g�)]���!"O�d &�A%i�.�y�	�^����#"O�Y��+T����b	�8�X��"O١&��- ��9*�)f`bH�b"Ot}8s��3�Y�@
 0"Z���"O�Y{VeY�9MtᒳO�J��0��"O ������li�T����2�
��V"O69�"�-n�x�0f��q�p��"O�q� �����a��=!_��:�"OJq�Ю�,h��MHD�&/R�`Q"O>����~�<u�TB�T3�"O�;H��g/Ե{�#��j?BQa"O�Q���/]�a�����*��u"OpT�|�>��6�2
���qq"O��QU�Ҡfq���4�ˡ]-��"O6=acnK�S*uK���';���D"O�k�KJ�x�V����ɋɖd��"O��"#6#��*C�C�9�^a#"O�	�s�˧u�����M�D�<���"O�;T�^j���*vֱt���A�"O���jT�N��Fϛ!V�`��q"O�!�B�ך�*	"$����Q�p"O�!��`�U�,9PMT�j|�[�"O�횐���kW� �H�� �"Oƀy�#��P���nH�"Oxx3��P�r�p�bV4B�x�&"OHЂc�G�0�i�`�~ܼȪ�"OR`�s�ؤ{P��C��# �L%��"O�T��%�=A�q�#�!�H)�"O^IS�8X�7��1\�\Jw"O�a��-���NL%b@	6�%�'"OF����Y�lقTN^+�ݹ�"Oj�+�hߛ~x��@�ǝ\a���"O�	 �i�mplq�,�'�W"O���3+^Ǆ����βE�y3"O8�`������eK�!b[�����"O�D�j�͘ŮY0�1@ "O�x{$�����;a
Vha6�J��y
� �	����%� �`Ƥg��L�2"O����C��x	�׬��V�mZ"O����$����M�r	���"O��	EƉ~�<K�֤Y���S"O<�V$ɋJ���F�!.�`�"O�Ĺ���9_7T�HU��,K�"OLXrV'ŜQ�Rx�噚�.��"O���\6���8�֔D~d�&*O�(�C�A8E�!�Q��?���z�'�
9b/L�-@�I�q�� �l�	�'6M;�I۹"qp\zA�A&)�$	�'9liy�脳If
����(�	�'��%�d�	J�4�p�	_��)�'|^��E�F,6 �p �j��h�'5�x���=���` h��o?�e�'�b��@R),�R4��_c\<��'�(a�p�@	a�l��eI.'Zƈ	�'�l|�"�A�V�n�t"ˍA^���'���R������Qfn�4X<A
�'�ְ�1�[�:JZH#f�\�`h{
�'�Z��@���zBLs�5Q�
�	�'�T��2�X(x(��D�����'�P9:�����\�`�k�8����'�R�2���<'��Ae�նbה�p�'�I;����̠4�!b6���'�(d��W*�|9�(��\�>�r�'w�Y(��"��C��i6"a��'E���A��T�`���4^A�I�'��#S��yd��IJ!����'@��3��)=�hX�ѿ���'4,�*ף�0ҹj���xj�'T��U�NK�m�f�Cg&�a�'�(Du�A,����V&8�ux�'h�צ�8���Cƕ%:��Pp
�'L�A6�O�v����B,ۼ,�ā3�'��E�V�A����"X7x�b��'{��2�$�-
�3��3#j�I@�'�(�&�	��d�(��ާJT�U �''����,��=��$�ɻyH��;�'�.Z3�*I�fE���C�%��B�']z���$ؒ
(J�M�F�8��'V��`��=�(!��.҈w,��'M����~�ts	�kh���'C��zT�
�jXn%��
PY�y�
�'���lV�9��E{T%B!>s,p�
�'�*��ʫX>5���1�(A�'�`h�b�7SL5�wM�)�]�
�'��0`A0'+���V
��
&��	�'�\�9���f�x��"���Q��'Q �P���:n�h��0R�,A�$+�'>�-I�Y������s䙡�'FL�hv�0˼H�#�=m}d���'l�6�� �J����R�oF&���'��a��;��	t)K+V�^4�'�`;��G�S��]���ET} UA�'\�L�d�1m��`2D�!��L��'�R�!�ʇ?W��}���2��i�'�($�A�
	P�زir��'S�UP���r�%n�+P}�)��'������R�dZ|@��
�N�:e{�'l�H	��á3�B���,F�̤��'x$R�V$`Ȑ�X���L�B��'�-뛈.�`�!��>�N��'0r�Ȃe|m�g�5i$�(��� Y���+�D-ش �\�����"Ol��Pk~2@B`JB�"���"O�m��f݃1��5��T�@�rA�"O�\��  �txAK�`�xyѢ"O$���@0>��z�ǢϢű�"ON�� ą����+�Z�V���U"Oޝ�Ub�-�q	���(~ڢE8C"O�Xy�
��D_����l�2qC�"ON�q7���@�}�596�\�j�"O�ɫƥ=r�C���>�\�#�"O ���hɼz�l<���I���8�p"O<L�$��=�dق�G�x�x2f"ON]�n�e�LM���L�#^.�9�"OB�0��\(kLл2��%FJ��"O��J��T�L��(��ŝ=2�Ċ�"O������2`�N�9�#�g'N�T"O��r0���GJ�f�U�K��"Om@��)]����& ��d��H"O�p��C�h��viN�?~�)�"Oh�; H�<"���!���5�HXj�"OqY��6`���w��v����"OL=JC��*`��&�A f���V"O�	GʐS�����@�ro�u �"O�����20�A�*ĽQ(6"OH}�r�\�'���SU�o6��Z&"O ��T��)w7Ԝ:��K�5X���"O�q�U��_��5�����>�!�"Of1�N�;��5
f��l9w"OX��DH�&[*��6#�Pۄ�k1"O���װ"���c��ުid橈!"O"���"M!6B'�KJm�0"OVԊ�"�eU�p��`��c���"OB,���Ƶi�-���[�lu�"O���@� ;rH��zv/ʒ4��I)�'��4c%E�!6'@��wk��[����'���H�yn*�c�7'��}@�'����c�T�k���q`ӇN,�
�'`ޤЁZ��Lp�@F |��K
�'�ç�A�ܚ"a�u�b�(
�'�Mr��U�/O�p����lFؠ	�'2����&]����	�<h�����'�<�ƌ��?���;�E\�fUS
�'\J��Zr�Z82ÊQ$	;:�*
�'�*0�G��E�&���(��'����t�duz�/��~^��
�'�д�dC�0R����R#��h�����'�������;G-���.��� U"O��87Fx3�t[��M�:iZ�zU�,D��c����4Д�C6��*|�V�1�)D�h�ׇ���b�KM2��,� &D��ǃJQ��y�3#΀
�{GE%D���%��_Id�b���$	q��"D��@�g��e��Xj�*I7]��@�-$D�@p-͌�H�.0uӑ���~!�d]&:(�dEĠ�iCM�*/m!�!�4%wN[�m
¬XQkզoK!�d�*O�4qPƚl�s媕vV!�D�Xk�U��U1sT\���ϳ]!� ^�J	Ye��L�4��T�(~!� [�r����?
A�,Z��/!�Da����N+g7�0����K�!�䃖s&`0e8I#�\���!��%r&���]��ʹ�r �!�dC3Q�,���ș7jT�� D8v!�� ��"
��%� Q>O(�g"O.�',�8��H1&��{0���"O��xĎ�[5^��c�POF��"O���ѳ8��d8���6v��!P"Oz��u@$;�^d�NԶZ�d"O��b�.�:	BWT�s�AK0"O��Z��_�(}�ѧ�	<7�Y�"OHt[`���4�Z1�G��&=.H�	�"O��1i�iz��@��C��j "O�S�b3�lͱ�j� u�)[�"OqpMX>m���B遮 �����"OB!sa�W� �k��R
a�޼��"Od:�MRe	�;�F�+t���"O8�C ��+�z(XS@F�FcfHy#"O�t��㈫M�t �.�.%徕3�"Ob����S�J퐗.�$}f���t"O|`Q�*�.AH��sHΜ����"O��{���(Ip-�DG0^f��Be"O`�Aeٖp(��Y�L�r����b"O\���ܪZ8��%D�>&��Ā"O9�s��9;��d��bS�\�mR�"O�x%�ȳ�|H�& b��2�"Oj�*���e����O�-T[X��"O\�Wf��g~����A�\�
""O (�M�#@S�;�A�7T����"O�\I�V4hG��I���
�>��"OLXhpg�#ؼ��E�h��D��"O��C�eW]�6-r���YU"O�0`��.w��D䝆FH��"O��Ї9piv@���>h�.���"O�HI�o��7/�5D�h%��"O�`���ǣz�� ����0���"Oepv�T+:l�a�T���}���j�"O�)�[�0l5jGaU6�<a� "OXı�$��E�E���t�V�Y'"Of5ѱI�:|� (�*�$����r"Oh��a�!2�J�S���&�h�w"O��!�S��)����#�@Y�"OʐP��M���8��_3k&��d"O<�x /q}�GR*I���"O�tm��Oj�a�$썹�@��"OeR���Q"�4X�I�3�fAC�"Oz٣�T ,���f�4S�b�y�"Ov�Q��4I�V4��E��\�8R"Oj�2Q�7�ށ�â
U�����"O�h�A-'$ݑ��[��=��"O����I�1$��ģ�`Ķ\�(��"O�<9�!�9����!`�N�����"OX��jٵ(��=
���M��*�"Oԩ3��N6��� �D�^�
D�"OP�� E��x=,� m�!-���1"OB�1�[���}���Z q��"O��'�իn�^�j�'F�&~~,Q�"O�՛�L�������]��^t��"O���M[��L��5,�!gt$��"Ox��1�� �&qq���)f0pz"O�Ei�*,���|E2�{�"Or�qt�F�c`�\S�)�&�<M��"O�I�'�$@ʹ�k��U�����"O��S&.�H0���d�u���"O�%� ��qT
=�m��nܥk0"O�e�pO�3g�����ڀKN�y"�"O"$�2�Y�vd��*�*��W��]م"O6�p&�O�	x�а��β8�&�r�"O� 0��,H�1�	�`���E��H�"O����$7��d�.�/�<T �"O��s�c�,P�0E�n��M�kf"OT�s�o�1���B�+�5z��0�"O깑��U�==
�s �F���Q"O��t&�w8y��	��M�1��"O~-!�K�,^���
��7�@�( "OPQ�N:W�������mk "O)�F�W� ���2�C�Y�e�Q"O2i{�G��,pD���o��j�Ji��"O,����׃P������gݬu@%"O�a�U@7@I��g(ғäъ�"O���))A�D�ZGEH�]�:("F"Ov�Ƙi����R����j,St"O�����J��}#�%��к]�D"O��[��68=X�ÉbnVh�"O��bA	�.��H� ��\m�5+2"Oq�G�.��p��r��93"O*A�$'�a��	��V�wS��!�"O�(�&�ޖ���k�5E(Iˠ"O���b��<��c`ܬ��ʧ"O��j0��%����D��.�|��U"O��h��ߴ(;�<ـ�ײpƌ��"O��U�=	�\�H]�� �C"O8���BD#�!X�%��u�3Hѿ�yR8��ÕK��ڜ�VhϷ�y�K��)-���,������y��[� <��3
�~����C.���y�B�頑��f�ki�+Ŝ�y���1�R`;��R�l��}˷.�#�yA� @�6�x6�Ȉ<8�Qd�ʯ�yR�G�Z� 5��kC�e�b�RM�yr��^��X�F��[R ��Y
�ykVJ�@��'�?�Qh�'R��y��ɾNt���$o?��i�F��y���/��(�
�>D�,#���yB�N'*��3�Q>D�y0��;�y���0,&X۱#J�7�bH�����y�.�jz	Z�c-��hh���y"f�U�BTS�XO�œ� ��y���NLAS�L�.8��b�=�y�#�g�L-����=�(��Sb��y�ˍ*��tc&n�+�p�#��	�y��M0RUYp�  |$�Ӄ �y͏L��,�1�K6=�ÎL��y�"
��8d�Г{� p����y�Z'6F�R'o)\�"� ?�yr���*�����c:U�eI��y�&Z�J5��TaL���Q!�yB��a]�2_+E8>`;sƦ�y���l8uڄ�?q��@ZwE�yr��S�*�G^R1X�S��@%�y�ۈl�I�_6OM��O�yB�7F\�t�ި@�|�0#���y��Ĉ��� ��37ܜ9����y����rU�J�'�0�ab�i���y�A���b����%���%&�yª�=�F�C�`ކ/�t���A��y�ڥ`�g�T�(�bɰׄ��y!Яx�ab���!PHT���U<�y���	h�@m�"��J�.�p����yI
�;��Tх�Y�N�J�C�'��y2�[�4yÒ���Ay
x@wK��y�&]����j�4R�<��oQ9�y
� ����.K6ޱ�ƫ@��Hx1P"Oꬨe	G(���A�"�4�z�"O����N�0aR���T?y}��"O� ����2 ���֤�FgfD{1"O����O�"-�;�i��5U�<�W"O. #��J�-8���k]}�z-�"O�HȌ�w )(�K�u��Œ'"O�	ȥ�H;w�m�S�£g�t���"O~��7ME?V_&�K�I��ةq"O�Ujv�)P�;-Q�sKխ4�y"��:�����uB�!
]�vC��	O����*��WL<�ҡ�,C1hC�IN��doן�ʵS�i�<.C���L#5.٧[ȱC%3J^C��-I��8z���p�j1Pen@�t�DC�	?	�҆+;r�Pu���]#`C��p�dL��!3�	�hH�g��B��.G���a΅���P�B�II�@��rl҅W��k�fQ)\�C�	4{I�CՏ^�rm�KcQ�?�B��q%���%��*P�`�V"JfwtB�I5&�`؁,PK��4�sNF�ER�B�&M�|��CfR|����ն���y����,�Z�0t@��Ό�	!�/�y�(T�������^��$q�O��y��V;i����Q �Y)�=�D����yk�N 3$+ޓV�L��^��yR�B��d 	r�Z�K�>��S�/�y�Z�(�y�FF?���c��*�y��ʩL���	��Į.��`��) �y�HT�#X���E�*�Ti����y���-�����EA%���!�(�y�	�Ȍ8P���1Hߤ����V�yR C�ys��6��< �,:f�&�y�Ȋ��yY3˔�-<������yN��nAx�@�l@,)��p��K=�y"�/Y,�m�p�\"m�xEe�Y��y"-�-1��y��X�1���yZJи��"��(V�(P�`��8ϲ��ȓ'�JD0gbA�V��H��=^ ���-��8#(�':zY�gӹ����'���@��S��U�ϵuu@��@���C�S�'D|h�a�1�t��ȓ4(��S:<��̑V���E�A3��[$�D�O���X��=�b�����<E(��@�݆%�p,�ȓe�s�8 ������'���ȓ`|����ɦHMҰ�';DbpE�ȓj�\=ˁ�N)�
��D���@���o
�y�n�;��ruBR�\�`�ȓ֮l��&
1QtA�7o�1vʝ���ٓ"^ԵZU�\�FX���ѣ��y"�Y�\�x)�q�0>*(%H�f�-�yb��W��TXR\�:T�	!��ݢ�yra�2�V8x6 B�[SZ��7���y�jK�(�(d� X���jd� �y��+5�@����Z]R-��"��y򀝇LB�t����U��C���y� �-&i���K�������y��ҫL���k���Fq�e�]�yE�3p�X� �A�ҹ�!�&�yr�Ԁoh��1�Z62��"+���y�мpq��nӠ(C��)�y�H�?y>`���*�[���QE5�y
� d�G%�0���gфd)T"O�P��ǒ0p]�I�'���1���r�"O�m�)A�?`䈛�M�.J��Zu"O�����tJ�}�q�6�T�� "O���F�6�8�%oO 3���X5"O�5	u�I>F;��(��S3!ح�q"OZD[�cG44X�s����d$*P"O�1���#f��h�/Q�4ؑ�"Ob�z0h_�ሡ�6�X[�"O���'mŀ*z*pzC
�<e�͛�"O"Q����KXJd�t��q�-�"O���L=���Y���"��S "O ��Ѝ�<.���%'߁��M36"Oxܲ�̟c��q�K�~�YB"O�qQ� �,$ �v�V.>�"��""O`�+a߹eG���&E(2Q�g"O��@�?##�l�DB=+�:�J�"OZA#؛aH���ьW�N���7"O�p�l�+=L���W�r�XP "Oڵ��'T��C�K٘N>�)A�"Oիq�)&��k�
P�R)&`��"O�I�D��I7�}�d�ܪ`����"O�I�,E����R�+ ̙��"O��Z�j�*������ �HT��"O�Bm�fY1��E���k�"O�1�@��M�A;P@]4]�؈�"O��pU(�K�`�#��);�h���"OLhX�`˧($:A�t�:r��l�Q"O� �ϛ��X��*1��a�"O�3�C�3l����CȽq��Yk�"OIb���7<��"��\���"O�,0�)�(��|�D��P��p��"O�u�D��n�:� M������"OVAY�l��/ḭ���W�,����p"O�e�	)"�a!m^#&o���5"O�H�'΃A=t]�e���8L 4!"O�L'��uID�q�i^Z��ZR"O 0�`��k!����*��t�|;�"O����.��*x�*��5	[>��2"O���5�%uĹ�@���R!N�[�"O���'E��HJ���Ԍ�P�)G"O�p�������+�yc&"O �s)�t������)iJ̐ �"Oq�.O8Zt�}�����H���[&"O�l���d0N�P�e�������"O8�{4*Ϻ#\���?Ϥ``2"O�:"Vk�h�
udO��H ` "O�����vp��x��Q��(hd"O�$�6*΄Tc��b�#�:�Af"OD0 �4_�Y;& *w��2q"O>Pr&�R�����"0��"Ofq*��#�
͠ĎаF��TS6"O|��	�Z[j�#�L"�$#�"O���ƚ5�,������Y{"O��)G�����a{\���"O�t3K�7m�A�Ǌ��h��<�"O����ȩu*9�ЈH�j���"O�Ѓ�Q�2��4�N-n��H��"O`I��D�7�.2��A uB�R"O�D`��K��u� ʗm�ݺ�"OVaY���s��QQ$�=hF���"O>����&+�hFd�-c� E�"O촂��R�Vx8��r�ݡ8�(��C"O�Z�)a�A�1�{�T�B7"O� |sc���|mq����h�@�`w"O����c��`�~��E��S��D�"O��"�-BM�.�����ē\��"O��	�.�m�d�Fk	� F��&"O� � �O�2�j� �,P��P�"O�+%*Q7|�6���H��G�iQ�"O賠,C��LX�<9���"O��T�
rcP5�S���S�Pd��"O�h��G?\Ohipd��J<$��"O6e䉮U���갋�]��""Ol 0B��a6��c��7k��4"O�fMM�h1I����N]��"O����2v_�A���H�hjp]R�"O]�W�&J��`�.�/Nj�Ҁ"O�ђg�>w0�a7�#G(n��U"O�X�����eQs�2&�=��"OQP��:c����;��(��"OF8����I����5@��~��e0d"O��Um�Z���H���+����"Or��c�-8@-�$�>W��ӷ"O��h�ȕ�I��%��B���Q�"O�JV-��,<+#�?p�A "O���.S�G��-i��ч+k&���"O@P��@H�5L�W����"Od�����xjdE*�
��q#F�9"O"-Д̏�u�D*ϳ!�p*G"OT����ӢjD��qG�+w��ʷ"Of88 ǈ?(,�f�-B
���"O`�����"E
��胯d��"O
T���?�e���_�;��e�S"O�hZ.@_�����8�N�ِ"O�a1 .�=t.���L�B��$8c"O�9q�B
�E�Pj�	�
u�f0��"O����Ȓ=���4H��2g YjP"O�(����!"h�(Umׁ �(�Bv"O�D[E��L�"=��*�(����"O|��e�>-�tz�JF&E�i"O��˰d�&T<���IäW�R8��"O*BA�>s�͓�Ǖ<-�\J0"O��`��!��Ӣ'Պ@���Ap"ObDJG�� &�����կ����"O`�H���7A&�A��U))Z۩�"O�سc��ܨa�_j>����"O�Փ6`��:�h����v���"O��1
ʖ.9���!�hhR�"O �haN\�pԝ��Db^��!"O�҅"T3,P���ƚ?	�|��"O��;6N1K_��BP�)j�2��f"OJe��)Z1O]"X�Ԉ:�"Oz��gf�: Jh�qmYM����5"O4p��䈪J��0���^�ٌ}a'"O:�G�ȗ>���� k�0H��q��"O��P�U�.:�
Eꉢ]��B�"O��y"/X8b��ixvCH�4��zW"O$Ek��+�陆��}�6@�"Oƌ���ӹ%~ɒvl�c�.� "O�
/̄^��)#�Àe�h1a"O��8"Ȓ�Z����S0 �t�"O�9�E�8	zt蚗hBa����"O�&�)Bj����=iP���"O1r�$��u�2uz���+uk&�YB"O�Y�f	�<I(FYʖ�	�UB*ya�"O� ��ǧ+1�Xju�R�@'���"O%K���3,F���C��i��
`"O� � IZ�)�l�V��$�3q"O�	y�%�1K���� ���n�A%"O��4�.y���7��+vRE�"O��)�e�x{"� G�fn͓R"OJ,[�ѵ&�u	�ϊ'%n�m�"O���A"B�Y�T��c(��?��u�"O>U�B��>.mr0#���	H��7"Ob��ӄ7p�Y� �>����"O~��u`�	6'Pg ^4F��4"OfU�AL��@���(.n	�"O����"Ev9Fh���1=��@7�iy���Q�C��3�`�Y�R�����y�!�ǌ\��ԍ5Z@�g��S�Q��E��	�TI��sPc� )��Py�mS��y��T<3���m�i}�i�耒�y"i����m{�*�h��$m�.�y�)]D��#)���H=h�m���y�1O|6�3�ŞDWp#��������S�X?}��q�ȓJI���&�%^
(
t`�>T��I�=y�������{l�y *�
���T�#�y�f�8S�lۢ���Z,�C�ټ�y�S�^�N��1���{B���s!��y�jNl�&]��
��n�h�s��y�L�L��P �B4^�K�)����?ړOt��|���6TIFeb�ҫ��b�_��yR�4�6�2a+��������y��{3ԡ�%�O|jI��ƀ��y��̚!WN!���#t��Y �M�yRk�1-c���a�
��M���_�yr.Z�`��8�%�ko���b$��y2�A���m�2+I�^ϖ�:�lV��O�"~�'H�)|��'�׮'6ܥ��f�<�o^S0V���
��G<<C��TG~��'T��v�\39.��'_�F�@�'�ʀ�d��Z'H�2aBZ$����'P���a����-�PO�B.hhp�'WjT"�	G�0�	x!뙭�P��'�``,X�1�؇a�	����'��[B�˯7�B�"k̷6Q~�2�'aR ])s�Mi�#2-<.u��g��y2�.j�P���%�pY��9�yR*�%zօ�e�H�Đ�[F���y�l��h�:�H�MPGE[mC,�ye�F��A�'�Q�d�%�8�y��J:jHTS���1�BMEiY��~��'�ƔS��<\^��@��ޤPK�4��'KabMQ�1�}���Щ�ZK��)�y"��1bz�$ӆ�7`h���N)�0>�J>�%��Q��5�ӃN���c�w�<a���p�hXt�÷�QAuN�|�<IOVGh���$��;`�ڙk�j����G{���iJ�űf�;a�4|��jIl���'aeΆG�����\D�$y�)��y«�p��-jԜ`fʌ�����y�ʉl�X1٦YN>� #�
�y���?��QJ�D�<Q�i2��]�l�=E��l;$�;�FԳ1�Q��$��8��VTflr���sJ<Y� E]'|�D�ȓ)R(�DJK��@0��A�<�'���=E��$A�j���A�Kb��oް�y��z���cÍ;N�q&/U�yb�P2KQ:��
��*����pX���=��{��X~��%X)vβ��W��	�ē�hO����HaꜪ9%���nW&oȠ8� "O� ��ӊ��3�P�!6���r��f"OV����m)���S{~MSF�xb�''��Zt.�/i؜����R�2A8���'�-��!>˔p��j��t�`4���D��h��Hq���Z��`a�oѢE��"O" ��E|���Iq͜T��i�"O����;I�P���Ӿo��a!�"O�4�ʍpv����$4Py:dB'"O��p��:[����Ś�	p�2"O�����P���`3�[�=4�"OJ#�1|����1�R�U+�y��2�R��7%��1�\���yrl�J��qQN�)k<)�CR��y��έJ�� �� ("&z��E,:�y�`�?
��P�pl��E��y���^
y��t�,������<#��O>�g��,���k�(U��U&��ȓvh�$�Nِ$��Z���؂<�=���)�鎙"��3��?x��\a��� ���E�T/�T�V�B����ab�8҆`M��l��D#�|�']J!���mV����ݞ-���a���/ړ(�~�Z����uL�D*V�5���\���iAaz"��.�N8`�l�9e@M����ۈO@�r5ό5��M3�͔�i����ċf�<y"�Zw0�0"�<P��\��e8�,Dzr.�G���kpe��sF�X4����O�#<�'w	vP�5)U&/蔉�H /,D�lZW�����VL�r�S/ i�rQ�/���'�ўb>�x#���&���"m�^%���2D�,����o�l��t/��h���S��xb�i>U&�x�'##���#%Cݴc���kV�"D���FMY�Y*%
�t<���>�Is���O!,�D	G)�����W G49��'�H� �%�h�6�[*��}��$(�S�OԖU���'�*B����ƃ�yRJKKk� 3ႨkW���P�F���'�{bBǄJ1�K�M��Qt�}��C����'��6�	w�	&��Y���*�J��3l')$xB�I����9R)Z�(CX��a�T�"=���T?])�.P�l�����	@�й�W�3D��C�L�P�8Mg�V�3S��8��-D�H���G�0a䡔�y�a�-D�T�	H�Ga�h�2B)���J(+D�4�plI!�|�Z�oξjF��M�I<����ɔ�n:�ӕ���kYz �6d]>m���~��� 4�ھ}�<�Wo��/2�Xs&;D�,��쁦�������/��2SF%D��[s!L�d��L�íхP�*��5#%D����2����񊝔uN��5�6D�l�4�F,�l!KP��><(�`5D����k�*y��z�H "��b��4D�p1�*էW������ QJ���!4D��#HƓH�B���"�.ki��&lO���O~���k4 @8���7Jb@Ij��L
��O�~ڧ�\�I4����Οz�~@����k�<�S�W9>����V�� �r�<q6�@-,�Vb��	�-0���p�<Y��Q("H��� �N%����Mf�'ayrDKH��u�!ŏ�UV�!c���yrb[����Rq��,�:�+�H/�y���[9ؙ���Ο���b�ך�p<yL>ٯOR q�e!�L���-�;��B�"O
�{�I�v�nx�VG��Y��P��"O�@r7lT�`�v�Z�$�b�"O� ,�a�jL@�^Hz
I2-��:d��TE{���'����Íڛ�dX�$$��UQ�Yh
�'w���/ԛI�zCL�8G�d���y��'WR��=���w�*Asc	�' �7�R<v��DHZIf�1�	*!!��{\�����CnP8ds��H���<Y��I��� bÍ��?�~����
�y��B�>N�\Q�c#֟;�n\�E��b,�B�ޤ�ҥ�3.;@�r$�Z�T �B䉉<�蕲B�F R�����Ę�T-�B�:j�nuy¢ګ0�%�u�[�TSVB��l��-��鐞x��@�X��C�1���s-��=u�B�I�ff:]�&�H3�@#��
9�~B�ɣ���� �4i�x����>B���1�ab�b�j�R�l�j{�C�ɗ�]��C�f������B��8@°�b��Ig�����B�HɴB䉷/4@xі�	
�x8;ǈF�ۦB�IP^��!)�&�9�D
�jB��${N0�a�.��2��I�dD�D�dB�IS8R s AS"'���`�OD,'.B�I$r� �ɓ63�Ʊ�nB��C�	3H�:�ˀg��ZT�m�Ê3nC�Ʉ��)R�i��$� b�;[.B�I�S��8��"��Tv�����K0"��B��
A�X�H� �min̚�D�.d�B�	1^9��cޤsQ`�%fF�I{,C��Pf��pR ���ϸ,��B�I3op�{�JL�Q���.V��B�I g#́sԌI&��iGK�+]�~B�V�iB�� }���ء�� �,C��GP���ą#|����6LC�I+^��"��ȬT.�}z�iV��C�ɒ���
^G�� C�@���p"O�QS�شAN��j5E�˦
&"O,�e�<J�Q1iQ"�0$*�"O�e����
 ��h�'�2��"OAV+��7��#抏��F=с"OrQcth�6n�J����\ ��Xɠ"OX�@�7�n��רԜt~���"O.u[�'�dGH�Xpgƴ>�$ɒ�"O 0���$s�~� 쒅n���k�"O>D���� �����*\%"��!&"O�\����5m��k7 �#��[�*O>�qf�ݬH�l�0EPT|�X�'�`����D�
�\�9ӓ"��[���2=�<�b 	m:.ņȓ&�P蓶G�._D��ʡ�����D�Z�Ν,�l�+Ɖ|�������z�gԅ2��ImeP,A��|��h��ueݥH'���u�݂	F0���96qYv&E���0��)K<74��ȓG4��EL�:R�Z�AD�K D�LjT�K�uJDr��U(y��:3.D��q2 �z��� F�厽�a#D�������Q�^l��c+D��+�u�`ܠ#�i�&E�3�5D��"񆃻j����Sh	8N��ܻ��0D��0��#&�x8XaFK�4�ye1D���ӣ
�h�B� �{�Ļ��2D���w�,F��p ��w��(gd.D��"P	Q2[�R=��cF<d�btQ�o6D�d�&	�*i󮼓��ذ.r��1k0D�,S�˴��4yt��,�$�q*#D�� h� b�B�������P��e"O�س�C�r���!2L���@�'"O,y�WMӿ����� ��"OF�05.�k��)gFCłxR�"O$��(igZ4��ŉ4>E`�*�"Ob�s�L�<|l��P�0k�^���"Ov剁N�*:J،ʑÞ�e��hS"O�#��#P��/j^9�"O`����A�/��)�s�qS���>D� ��ڠ	$l������Tbl���3�4�HO1�t�唎@z��:T�;uY�<�"O����F¸8���`J�w��MIt�ĝ�oQay��LRv�]���"8|P�DK�:�Pxbf��yƥQ��S��X���3���gO����Q&qY�ah�A�
E�A�>D�+&��DXY��ե�$���?D���ЏA� ����R�O�xtk(6D�(� �0]�n%�B�ZV���1�^P���	>�B$x2���@��L9Dz�Oz��J��Ll"�ǒ�cM*%�a�5}Y��󦌉'��>���O*�����/-`�x$圐[6:�;v��?E��p���iZ!�B��D�h)b���#
&_Q�� ��	5s�}�I�b;xh�u��96o�I�&L������S�$�]��Ņ)pD,R)�0.�F扵*]Q�"~Ra�P&b��q�Հkb����"�E�	 hh�����'�꠨�`P�g�PB0/��&��-��O�T��y�伐g�X-Gƙ�!��%��x�ˈ�wӊ����~b��h�,���jsW>*`��0<�VA_���'+�Q����HV�dˣ!��.�f���$E=�����\�0��T&
b⾜��"O�0��.��r�l�`˞-"�8���9O�����W ,lRq����,-h���".C䉀����ݼ^�ҵ�a�<z��x�X���
"��!k��3��c3/�-a~2��C?��!F�*�.�&% 5c���@�i�<&���N[�\�C�-Y����#^�'���G�T�0��I�AZ'�T�S��yb��R*`�+t�ף`�R��G���y�b�z�����i�B 2=�peb�k�4�hW"O�p��N"�:���I��#�r�Zƚ�|:��'�\"E�ۼ��jQ�ޑg�L��J���I�Y���Ӕ3��}����6%4B�I)ZR�#S)M!Xʂ%[g͗<:)D#>a%+�?X�$��'G�*(V"��$_��$��W9�8˵���^v8X÷�O&T��P�\�n�<E��z�"9+ƭ�p��1�`��y�
+�.���Ŕ[��D��/W��I��p>٥d `� EL�5=}�dp�ʉv���b�'G��co���:����X�'l���H�}�Xs1hP!�Jlk���>�'/L���B�� �xX�f�g+^��ȓ�����9>2�E(6*����ȓv[�҈�$QJ���G�=h�r��ȓa�r��	+4��S� -9�X���uy��C�ᐔR��kk�6|e��ȓPH�u���]0"Ж��b���.����ȓ_6¬�+��1>މ1)b��ȓN���	�n�A8����A3���]4�QG��$�B��X�}��U:��K����N��`^ġ��sY��ǩ]!�Z���`��=�|T��y�*����9M\,�"�$�-6�ȓ+,6���=��(7+F�,��i�ȓ �v��eM�(��L"���Ks:��S�? ��āݫ*��$3�'&�{@"OD1�D2Nd���g-�3Ir%�'"On:f�ٞ^NZ��T.ՠyf��"OD+B�۩|��SGƮ{����a"ObYZj���C�l���+�"O@@���2� A�4`��:�"OD�A�ƉjP��Kb���Bgh`��"OD�bl�-m>�{5�߷o~��"O����&j�Z���&��cg�t�"O��S�O\�0d��)q�66tU-�y�� ~b��y���\5�d��(�6�y��°Z��,�^,]nl�k���y���H�h1�_HWL�2�'J;�yR���n^�i�a�	��t!w/���y�fC�Xz����ڨ�N����ь�y2�y;F9J ����`L�Ⅿ�y�.0�s��R7V6n�DF�y�"R]k^A��*�V�n����yB�.�<ݳ�.ߺZU�-�U�,�yR΅�H
�:DF��D����E��yϞP5�5�#Hɖ5���P����y�"��(��;�#�-%�h��A���y��U �"H�?5� ��*F��y��T�.��S7�:us����yR�B�B�ƽ���	#O�6�3&n�+�y�&�;�zu��$G:d2�@��ň�yB뗸o�Z2�׿)���HeK@ �y"X�%�&��c��?���\��y��[
x�>�p�c�,-�#���y��5{;
���Ε'p�[�]�y"�x ���B J�E���p���<�y�肺u�q���k�TY	�]��y��O��$�Rc���6X�1*�$�y�K��=,8��H$�b��2�7�y��ōkZic���<$\;���y�Ω<�YY��߼N�:}!ABN:�y�n�p�,j	K<�2�3Ή7�y�� ?y�Zu"a!�b�����Q��y@�_� ї��Y.�D��,��y�J�w6��8�	F��|Cэ�y�M�j3�>GQ~VB�S�XC�-��9`'���$�B,�@5^C�� ����� F�{6@Iȷ ˏI�0�OBM�� �ɰ<)(_�'�v��
݃1��mم��J��d`��� }r橊@G�(q��DZ�`Jj�����	u!�d�5eA���b���C���HD{2A�dB�Ѳ�dX��.�	�(��e��IԐ� Ur� �g�!���5bI�vO�,li{�b؋z�Vl	���g#Ŭo�^ kAo<�禡 ���g�ir3gM�?;^< �.D�̃�!�D�ن�W�d�̝�4Jؽ�)��o]v�q�,\�L���g�'
�PEC؛z󘱚aJ��w'���؍P�j��#D@���(yJ4�a*�M��ː�X��&���$�O,���L��9}����i�B���6�I o�&�#l�<w����C��S�qdu�7��s���%՝?�ZC�	�a ������I���W��fRj�
6bُ=�\H"!�(~��)A�Vm��y�D_�n�ʂ��.\B�Ӫ�y��B.�}p@�,v�U�"��=��|8�؆rX�27 X6/*�-��O/ўʄ���(���qgo�1Sh؊f�,�O|��#V6.mQ2�@?
$Pq�"��e��Q(�"- ����@U,`��O��>]b%B�G1�qb`T8y��g�ß �M��K5�r@�V��h�䤍�w�c���7~��@B�yr/؈(K�<��X�_[�Q
��F����Hu'��u%��dlf�Ya�s��AŜ(@�z)+�ޜ>,���I&D�p�N���=j�"
;�E�K�&C�iQQZ�"&��3�.�&-���V��� �h !b�;B"ГqF���=Qb�'�ĸ���ww"�HQj�2��$�p㔎3���k�`1�d3���6�}EJ�{��i!�c�Z��(�P�M�(O��B�����Aq1cKY��$�ȟ�d��(Ըh<^DS�Ke��"O�`��"��g���*
�*ؤe��lN�i,��J�/ϸ
����͚�Q?�d�	�9��G�+A��90�#a�!�
W��Jw!ѭn�d�k��q��x�t����7:�Z02�[?#=!�@$p�h�1ㇹG>
%��mX�ZЍ�X���D%�/+J:h�Mn�`�0W�C�lQ�쪒��F���h�_�OF�T
s��wFD��;ړn8�5��c��)��P��=�	>rg��eE߉>��]�����!���"%�V]�g�Q}^:����Z�"��Ċ="����M���)�'s�LYHtgV�xPl��A=B��ȓB7b�0�f��?�F��oY#T�e$���O�Tay���k�T)�OS4�~eb׫�-�yB��
�j���GT.$krd �T��y���1:�J�������s&EL��y����J* a�]0fS��A���(�y��Q��A��E������s�O��y��Z%lV��g�/t0Y�#&_��yR�F[�5��]%F�(%������yR�@9�8��V��9ǚ��gjX-�y�Cn�͙C�79,���ݹ�y��0|�hu¤��&�a�CkЖ�y�:c�Zy���%�Hx@*:�y�^�E����jg�M��'���y�_
p8Э
0I#fE���r	V��yrjX��}C���',"���lL��y���n��I��E߹1�P����%�y"@C�E��`�¨�Z�`cEN.�y��Qp��$�����H��5`V��y�D �z�Cr�~��Y �@E��y�/�8k9D%"'ʛ�`A�z�k�y�#zf�Ur�kޯ\,l\+�!���y�o��2����\H�	�@c�'d�ŒZ��]����
}<(���u�<�d'�q#�<��� �j�{��w�<ѠF��%��i9- ?<��I��/l�<a`G�s���%#'�.9�Vm�l�<y�@�=�"��_#j����A-�o�<f�
+�� � [4&x�5cG�e�<QD�L�^=H����њ M
`f��c�<��������6�ȑ(�};a-R�<I��I��|�V��4!���J�cIH�<�k�!Y������C�@@��YA�<�'�Ǡ(8��9WDG/6q�q�[x�<i�mœu�b����)&�*D�r�<	5G�=���rF�ҭ<C�E�Ar�<A�hþ � 8sri�w.n�b��q�<�w�Ȁ@L��+`��x�
�BԪ�i�<�F�ŠG����tJM�F�:咢M_N�<�OL2X����8k���k�Fm�<Q�-��.� ���Jh`|��&RP�<�c�_�g�,=��H�i�B�9�k�N�<���&N����X1��T�$l�D�<	)���S�����X�W��C�<�FHS8/t�.]�I3��jV	�C�<Y�L�B�z�(���>`n�\2��G~�<YtG�I!X9�b ;de���s�<1�J�6�Z��µ]?�Z���R�<Ѧϟ#U�������4����Ak�<1���`P�t��$ �q�m�e�<c��$S���z1k�+|z!A��b�<i��7+�d���`�@4yǈ^Z�<� �����D��l��K0X�q��"O�"fN^����[%J�6Ot��V"Od��B �<vh)�UI����+�y��P8&,�I9�ժ2��8�0A��y�M�� �jFF�=� ��H���y��G�J�Z�j�+�e��Ё*�y�!s�ʈ+���:���O�yb䝸|ʬ󃉀9}���ԣ��yBl��v��@�Zht�i!��S<�yB�o�v���$ɉVJ���EI�y"e�>(�X����?�R�I"�1�y�T�#d4E�P�DE�`X�(
�y�L�%>%8�Ђ��D8r`97��yR��>"����$Bz����ɷ�yrǅLٸ��h�u���E�4�yB�K�s=���M/]Y��q� ��y�b�tڵF^���� gU�y�+��=��u꓂]'r!r�0HD��y�H)cS�衪ѿ[�\�R�B��y�OԦ#Tv���b�<QC�TA�K%�y�ˆd��q���J��,Pg/�?�yR�F�`��c�GK��~MK7Ɇ�y�.D(T�KG�ӋyJ�Ջ�ʬ�y�i�#E
� Z5�$�@9�s�0�y��;Y�.�:k� b� C�\'�y"�	13\0�za�Dg,ԚW���yR�K�|XH��%U<�h50PJ��y" 2�b�ƣ�212�l��'Ħ�y"�(3R���jT;1�$1B��H��y2���A��	(��e����@���y�J�h�`���.>��X �M��y��`P-�bI�vR��b�S��y���r��0aT<r�Mb���
�y�N/�be1�aY{�I!�F3�y¡z3p�"�b��-$ra�GW�y"L��a����M�#M��Pf]��y���d���Gs�" GE��y���8P˜$�e�-��Fa˓�y�=#'�9Ȱ"��I00�:����yRL�GQҨ�S�$N.h)����y2C�*<zڬ�bL˯N�����CL�y�l�1|⹀GLő�����J�!�yR���9H�0�ES=y���*�h��yb#H"։raH�q��T�"�-�yr��r�L��!D;��k���y�m@�W70����zm�X�!�K��y�@*غx`���u=��:aƞ�y"��u�(�(G��$t���藺�y�:8a�8˴DQ�|�X�����&�y�*Q�~>��̘vN- �7�yBh��l��e���qΐ��7FS��y��>i���FF=ޠL:gQ��y��U�%,����*3��Q󑭅��y�N�*$V�k��O&5�t�ah���y��
��ၘ�/�~��v,���yr��+[[J�!e�]I1�%06hB��y���[b�$h��K(�ɩE����yrf֗L���pӃPA���E)ȹ�yC��>
�`��خ8���"R�V��y��5j\Z�!�dE�$A���y�{\\�9�)_�FBj|��Ğ�y��?;�ޱy�F��k��(j�g��y�C'u*�B��mu6��pB��y��g#�����Kf�QЅ';�y
� ��
���50����lP =�,��u"OY�"L+W�߷�f� #"O�$��O�%8@�c�:>cj�� "O0��e[�s����T"O�
6ܤ�e"O��x�)��
D�r���8s��#"O,ᣡ�S�TR���%m2�T�&"O0�����(����ՄO�yB���"O�t�HQ�|y�K�bC3( �yȢ"O��H���=t6��qNY��@a"O�<j�-÷e�2���l�tUr��%"OxE� �P6Bx��p'�ʗ{�Ts�"O�dCF��AB���DѼ^�X��"OzA�PfU ���;iS�W�� �F"O��䦙%94��´o�6!
�S�"O:T�WcM�?VZ��O�8P�#"OD��Q&��SҘ�a��p�*��T"O�$�V*� �Z�K��U*��²"O4u��% f4i�B�h`IC"O�� �هr'��ե�(Tl�8�"O����BM��ʀo��k5"Oޝ�⁇�fQl,냅�:l�U"OxQ������W�cV�!P�"O���$�Qz�
l�mމu6�݈�"O8`��,�7[�t�r��P";���"O�ݙ2ံK���)@��:�n�+6"OV�5�L�T�C�b�=k�bTA�"O8!V�#?�`��!�F��#"O����Y5�8(�\�Z�PX "OX$�3.��3��C�te�"O�  �F�5$QP���:�<p�"O� ��Aر�d�
�� h4�1t"O��x����"�I!���H��"Ot��3o��10 ;6�UVG<$H"O��Jdµ}+pH�F�0J���"O�Z�h��K�d�[c$D��z1��"O�sad�l�X�c�;z�(M�"Ov�A�Q�c���P�B�}s�}"O�p�@�� h�i��L� �d"O���`�>aM$12C-��-���"O���$C�%|r<��g�62�m{"O>��boV�Tc�H�Sŀ�V��"O�Rj��o9Zm�t"�KZ�-i!��6�����n�
��L$!�D	#�DHa.^� @F����?!�!�P�m��J�c�.X8v|&ʘ��!��_Έ� �$�@Ĺx#�

�!�D�*��0E)�!����!���ssH� #��x�:�,ޱc�!��?B�N�!��N�~�t@0���Z�!�D��0��l;� ��U��y��
f/!��4/:Hl"R�Q�~ʼ�5�G8E!��聢�`�/<�Mˀ��x!�d�1!������{Q�����L�!򤛻_2L���*T����!FB�@�!�Ĕ7	<	8G��>��8�!V2�!�N2K�޹�f��h�iB��x!�D�� P#X-;f. :h!�O�0��X���=�h0���Y!�$�3ZC`�)��B�|=L���k��vJ!�ï&��-AA�"8�h���;#K!�D�� �T��	ߵ?|*��.Ĥ�!򄍵���f�8n�9��F��P�!�$H$�(�P4��1e��}��T�!�D3r��0�Q(k��`�q� �!�� ���S��}jSɒ>3T���"O�HY�>c����V�K]<$��"OR];�c�W3�Ax��0v5�5*"O�h�݆�������.
l!"O*Y0���~�e�5y�"O��y!E��V�����O��A�%��"O���`n*��پO���1"O&PG�ݗ.b��c�C G�^B"O�� 6���4	𢈆Me�5 g"O� @r�22�^�iB��,T��I�A"OԨ!F�6x~���"�Y���}Xd"O�,���=w���8��ƴ#�$Q�&"O���#�#d��đ��'zp`�b"O
�Q���5w���C�	rծ���"O����h]�dV�#R�0U��"Ol ��/�5�$����*r��t�"O8��
F8�����!S�.��w"Oi�3h��(�pS�Z�4��"O�=�b�=w�4��nC�X�Dx"O��Cϴ���E#�%�t�r"O�X�v���r��y�N����"Ol9�3�]4Vd�k��5���Q"O���#cVEܬAq�M�}'@���"O�K&��_��AeI����"ON���h�?.ޒ��Å�\�Z�[Q"O�(9�-UQ�5a����� H�"O\�QP�Ƿ,�܅bBH+.����"O, ��� ��y�
�1�м�"O,yQ7�ǚӔ9k�ɂ����bf"O��1���:��SD����ĺ�"O��Q`�}������L�aA���"O��q�I�5�8�q�ՙ7h�b"O��ɴ胕e�H�A���^H��D"O�9�@��C�"���nB��6 ��"O`	rS!\�:h��F��3 �8�"O,m���t��]�
@#M5LH��"O��H���!����T�����"O�e;�ŰF��ȑ瑓R|<��g"O�5����c��u�f�|f. ��"Or<sV�]>?��@b�W9Kf:p@*O�hHRi�"�^�B##�*�	�'��]� H�_�e��,��	5�U@�'M� ȁ�G4K6��֨Ď�|�'�N�b��G5Y8��E��
MH�'��EY�l�<f�<b��C�	���'^�5)Vg��S���C�'4����'Ԟ񓱭ջ0f�;�i�#	x�q�'��܀g
�&���c�2
Ph�'꬀�J�@~��s�B,+�����'@uȢ�Y�%?t@�ҪY��4��	�'�������<�.e�!��6#��x��'�YZ%AY�Z�����A7TJM��'A�ݻe�ޞa��a�q��"[g�I�'��l����Jx�@
�ω�]b�N�H~t5�t��'g����5ߊ9��P��4&�����Ц�	p�1��숱z�4lj���=R�e%�l��I�
q��b�X����Av	�.(�B�ɓ3�lq0�ń$)z�c�A�9<�B�	07��|��D�<o`tJc���b4�B��*l�0��j '�|��ʝ�E)~B�	�j�6�[���!T:�"Q�5H�Zb���'��>��ǫ
%@<�*�71fL�GJS�F$�	p�'�Q>��M�{��hӔK�n,��s�gӲ�ъ��S0��٘1��;h.�����{�L Gy��$��h�e��6GM>H�.@�I�����DҾq��� ���qH��9������OߖlrA�>�U%������O$`�ss�HO�U[���c^P��R"V�7�����&���)���/)F@�M�t$8 ڼ[f�P���(��Tk1�O�?��W��HO�epekŌF��}����x�'T����W�P�K��ߋy{P�y���� tb�4y �)���b~(JA�Sr���b�Q�9��'��Ey����,c��d�#�9r$��� ^����%�(O��<.�P �a�'�3V�8x$��$����g�	11�D�ȴ�R#f��q(��S�U�C䉿5ƶ���ƲY���B�)��C�ɼ<�  �ff�Y���!��8y�|C�Ig�qK�ƅ� ��Q��p��-ʓ��� qN�=��࣬�	���II�'	�9��Q:1'�mZ`G���d`�ܴ'=@4B7�d��Yv	�Y�'�4�>I�a�W�J�Z��Ķ�vij��1D�,�TL�bh�DR��uF(� a�!D�D!@�\-p�P�Lؕ��1xC D�@y�ރQ2���$J�K�έ��c?D��#`�P����u����{bo'D��aNA1���G�^�Q���h*D�L3�&J���]0��}! �ʘ�~B� =��9����6��K�dNǰB䉉a�b}�`��&G����m�B�I�Xɬ(��+Mm@J!�\E$^C�	�:��(Ñ��j3JE;��[4J3�C�	=}Trl:�o)Gn�`&��)j���ćj�S����]��+ɏ�!�1{��QÕL��@��2kM"R�!��J�96�t��/�ybl �w
B
L�!��5� �y6�ƴ`X�\q\y�4��ȓg���ZQ埞RX��$ʄ�R�J��ȓN�h�i%��&gW�$b�C,3r�}�ȓ�zҖ�ٰRA�P[� E8^؇ȓc�)&���u��������y�Y[\0����#�`]�ȓ%����!M� ������V�ġ��m�Qh�b��)yq�C�u�>��ʓ"h$%�D��d^��@�Z���C��)@�E��g�4�v���ZO<�C䉊KZ)��m\~�v`1���m��B�I�=�Y��J]�w6�=��-�R2�B䉰!}2U���&���3�����B��,v������l-���#	J�bB��3^�2�B�?(-�U��#
NB�� �z�h���ij��6pVBB��J�8�QYĺ$)'��CB�l�D�##�Q4��$���?��B䉋qb8��6l�$;�X�eb��,��B�Y �"r�Q5+��$��@��B�2K^Ƙ�
[�x��9�A�˟|rB�!���+�Q쾑���2��B�ɲ4FD`�C�G��5;r�X��C�Ʌk�>)�ԇn z���;|1jC�	�s�4St��f1T���W�pK B�0a`��s�F�(H�`�iqʑ(s*,B䉜*�u�U�Փ:�TA`�	ѝ9RB��(���e�h�(ف��[DB�	9X!R)ؐ�1g&L���O�54B�/Ȣ�Х�ʢ�(���4Z|�C�:�L�{��!M�4��"+��+3�C�I)�n��#iؿG)��-��C�I�B�Zr���E�̹�蚕^ ^C�ɚ3䒭p�O�)CX���6�B�ɋNi@U��@A�7�ĩ0�C�)� ��q!N�9^�H�B�Wf�P�"OT�+��I�R�0��A��8���"O6-��fM_�Na:5�9f0�R "OJ)�3�R�*8�'Oˆ'��8 �"O� ;�*H\��aA阏tSH��"O�DH5O�8[a@��f��Q�ԍ��"O��r2ϖ<�����$N�^��"O�E��ƁI�����DN'�T�� "O�I�0�W�N5:�81Ě�16,�"O,)PD	59�4�YH�A���I!�$]-ED|�4�!`L=�����!��ލ��!+�ݔv ^� L�i!�7T���B �	v�	�X!�đ�z���0�F7bZ
��D�x�!�$ּd��Y�*��ҩ��Ē-p!�DֱQ���2D-[�)I�@"v�!�$A�-��Uc��,R����qm�yj!��?E�����Ωq֞�3 O�%j!�ė)C6q;&뜃r�P� �M�!D�!�d��H�����A�c�!�m^'H(!��^5x�GdZ�#���7�̤:!�@
+�:�7�C[Mq�툞!��Ӑ;38Y
�"X�-�u��c�!�d�Y��)0�$��uL41�5b3A{!��ԩ1�cV�N^0G`PNa!�DX�q���ےCY�?B��AG�X/�!��ƏD0����
�P�N�� ϛ3�!�Z(������Ꭱ)fl�� d!��R�I�Z��t���+��3�!�^�4	B����^��	�� 5"�!�����v�7��jP���z�!�%L��9�l�|5P@@Īg!�d�C�(�[�A
���8��ɟl!�\�N�x���m7b�BѧN<Ez!�$͙) �Y��n�`6�A���yc!�-��w�H�2'��Ж�
Q�!�H�4�B����(&�&=@�k���!򤏡.�6t tL��'���@QK.J�!�$�\X�����j��u�K<�!�@�qp�)�(�4L�v�jK��!��^�mĈ	R��I�6���H�i��!�Ej�3�i۠]��a"�4!�d�A}���N�}F� ��,�!�DԬd�h���ț @�Ze0ਊ1iE!����!ȇ��?ԈM�P(B+L!���^D���	80��ńK�7!�Dg�M�5�6Q7��{#ǰN5!�Ňy���Ҥ/[�\=
�+��O;2�!���ºp����-
ձ��=c�!��کi��mZ ��-**�i⠇X�b}!�$�5A��kc]�w봐ab�̑Dm!��ݝzr��Q ᆬ�x�(A�B!�psd+�3��7]�X8�"O����֤@F$Q�զZ��˃"O4�
gD�	8��8&ͯv�p�"O��
g��E�<��w�# t�%"O�9�*�p��i��E�mm�S�"O8��JOX a-;:	�̊�"ON,�d�*��QP���̜�D"O6ܙ��˲^��h��
��6e�Q�A"Onp��%��䋷	�W`:Kq"O��FL�?A�N��fꂑ4J��A"O��2��ʺ<�`����\E��;�"O�E�BND�Dt*��@�?P�X�"O� t�AB�I/P����gϸ�@"OT�P"�.muvm�	A;b�RY��"O�����̝O�%aw�:�Xe�"O��˱�X3�(�炣i�� ��"O��Ћ��BOFMR��Q��(��"Oh���	�['�|K2N�	�l�"OV���	 c5��r@̂�DK�y "O���מv�l(;2�]#y��}�"O�<+ƪ��!��@d
��0�"ONyp�.�IP����B��u�	�"OF�0��4�0�	�!R��Ұ"O����n��|�$���[$��y��"Ov�bVKF+!�p��K��4�xЀ�"O<��+B�b|�,:r䍹-q����"O��ɪ`�H��I�K]V�� "O�q	Bő�B@r��$�?3[`��"O��a)���r#�]+3�}x�"O:pS� ��M|��ufNg/*� �"OhЪp�J-��< ���-,�Xj�"O��A�U�<n>�q�cD���6"O��QB�g�,(yv�O�o���8"O�������t[V(Ȇ���"O�X�t�Ѡn"��Cցm|�р"OqӲI�C�v��a/�7�vՙB"OX��S%�62�u���D%bs<(G"O���a���%�uy�O،tr@(+d"O�r E,ai|�
�h�O�Q8d"O.x�ئ^ݶ�3gR�5D��27"O<er'�:�����bPX0"O6Q�J�b ����%�Q^��q"O>��/T�]������,}Gn��'"ORmk �G�4N�����(���"O�P��L<`�`�kG�F N�s"O�ՠ��0ڈ��2��&R,�#"O~�)�,t��v�E�-P"Oȹ��S�>$F@s%��d 8�"O,Y���R�B� ��w�W^�]h"O�	Yץ�\��uQ$�L�Zn	"�"O��Y��!)����RU>��V"O �c��12RD0`BH�i�h��"O��r�*�_����A^&�~���"O.���п%.|��t��m���:7"O��Y���>x B�1B�+�x�V"O���d�(��q�Nyߠ8#�"Or<��I�-t��@��b�W-�xa"O<���mN�i�Dq���3*���"O�!!4Ƈg�@�M<<t%�"O��F��av�D8c�!p.DÕ"O6D��I��'��p�B�Uf9��"O*H���!t��E3f��w�R� "OR�)�@��q♪R瓥�|��P"O6�+wJ�)UN��ƆN�&���"OB�t�@��Y�%Ǩ9Ȃ�jR"O��a	������y���"O�yYF� V�:5�7mV�;2����"O�X�"&�8+��(5�%7��H�"OZ�@�O�,L~,��M�U)D ��"O�%nI%m���wiɲq^	s"O8a��n��@P
�VRy2"O�- p�V<Y)@���(�138��9p"O�5�a�-^��'�g7N)�"OK1o��8˶�Һ�i*��Ɋ�ybG�YJ)�Â_��d
b��y�	�	+��R������A�S��y
� Z�y��3j��5sЎ�/��	�A"O )�p�߯�r��N�	N=�S"OF�k�¼l�<ˠ�N�8E"OlHy�nI4�
��g���)�^4��"O(�!KJ���}C�Ζr�h1Bb"ON��K	F�pRT��d��a"O>$�@EO�d�xf�®|���:�"Oޅ�v'���	pe+��G�VD��"OJ��W:�L��W*J'K��4�"O�dm�-� �6i�,��p�"O���Т͐d��mbFi�-� �p�"O�� rFƶ#Hp��4iY=B}lA��"O�0��B�<��S���I{F�"Oڜ�IS���K`!�?\l9��"O���EgW�r�d}�T�L��BC"O����#� w&>��b�K)S�\ͨ�"O���f���.�7DI]�*��U"O��#��O=v)�)���Ζ ���;T"O���aE�&�����B����"O.IV   ��   a  {  '#  �-  B6  ?A  ZM  X  dc  �l  0w  �  ��  	�  ��  ]�  `�  �  ��  ��  ��  �  e�  ��  y�  ��  1�  s�  � � ;  � ! F' �- �3 : T@ "G N OT �Z �a �g �n ,v ?} �� ŉ �� �� A� �� J�  `� u�	����Zv�B�'ld\�0�Oz+0�D��g�2T����OĴ����2�?Y���?��FJ%L+�a[6FΔc������)���2(�0A��3�	��LcF�����#��Y�t�i^\���	h-X��%C�f�%�_�VU�<zW�Y*@B�130Q�X�q$�M�(�*8��A����T�mZ�Qɬ��b�ޞ1cG�laP��F̼&Y�X���);>̀�銧.�:1Ѕ�i�B���P�������	�9��y3"'����9��3H������\��%(�4�?���?	��P�͓�?Q�esb�j�����j�#VR�RL���?i��?��?a��y���^FDJ�)����	�0+I �,��HƄ�6a��O ���I`~ri�6@Q���!X`^�Y��y��v��*��ӄ�>i�'��O���ve��$X��f{�#@bϿyv�`��@B�;弸sDH�O��o����	۟����?���]��;��US#!ؒ43�@3��{�Q��'��7m��Q*ٴ}��V�'��7�[l�lZ�R���:&n��zZ88W/ߝ~n�0�V�,���2�4�?IS�i�P(9 �'��u`��=|h���-�|�D|R��ON���c�)�8�!�ɛ%P�V�R��������S�4�Qh�MeӸ�n/�M��'A��IT	j��D�� �6sl��+ԁ袼!�0I�fj�B�v�(��1�"Yc��Ak��<Q�M�S�7� ��{�4_F8���*W_t�UAǟ:_�2��g$_�3��9Q��(q�f�x�m�Uӆ��3h8��90f�ߢ#�r�
SB���j�'@$=�r2��!09P 8���/W�$��4$$��Ol�X���+	^�r��[�n�Ʉl��)Z�-R�X����C ?u_zHlZE$����V�0td��W.K�	�X]�IH��!&�-��98�vfY	_���c��.����?q������{6xk�&�tӢ����<�d��E*Q+(ȀɄ�rlv�r���$�O���m>����"(ؑ��"P�k� �o��q��!���R!3��Y�����h��ɋ'��I`��.Z5�$�̥r�P� 6a͡]����0ȋL,"P"iZr2��刐%7�qO��rd�'��6�Byb�
��l���CѦo5�S�LҒ�?Y���?O>����?����?�O��yq�H�'Sz���L�"���{�v��.0�,�Q/F�-߼�@iB�u�(6M�O*|l5M�r�ش�?9-O�����|�Ĕ.WW��ue��m(�D�R��5l>�D�O���e@�?���2�F�6a>��o�V��U: �@
T>&��u���b���Oȍ����ZW@GW?�!��f�Ũ�H�X,��d�Z�D+H�q䦟Yl�eo�9��d�?;��~�4�G��4� �B(E���s*0w�z�r�'��IG� Q�c�8.�AS��v�<�?Ѵ�i�T7�1�ӏ>��
b�D�C2�k���c�X�d�Ob�llM���?���?I.OΥ�&��,�X�E�6�`��v��#}�|�Sȝk�q���]��˧�
'� �$��6"���uFˢ:��D�M$Pm��A �šov�oZ�s�l9�4��1���O ���ğ��y�
8s\r�Xm� 9�1�����j��f�<၏������L>1W�K2\�`()�)�z4�[���?Q����$�O��?�'�(1���Ǿ&�|�Q��Q�Vʴ	)Od�n���M�H>ͧ��,O��P����]�����@ϦWb0��4Aʮ��'{��'�	P��0�&�����C��i��Ka�'��H��9d�Ëf� �� <<O�e��
U�X�<褃�_Ţx6+�c�|ՠ2�KMR�A�
�S�D7\�'n�x��d���u���4� $ڀ�_�uj��'��7��l�'��O`Q�'�Z�[��-���t�l)XdO�O��d�O����T�XI���l\
�C)<��'�Z6���	�'�bΥ>	�)�B� ��>�ZQק�5WA�S��?��?���?1�8����Ŗ=s%�]R�&��u�2+A|6��ç�<CFV��0�z{4Z@��-.��L�^�R�(�(�"F�j=�6��`�AQ���r�c��TW�XHJ>i��ğ�[�4?��&�'��b���faXr��25kΠ1cV�` -�[y�W���	W̧b���xdM۸{^8��®��L��<��4F�dQ�����BM��p��[�P����o�x�X�R�'��"u�ajٴ�?!���?���65�QI��p� �*Bk��,��f�);������?�+�X4P���.�3:��\[2m/����]�T"��A�*)��LW��ErA����̺9*�B�.{dU�ƮZ�UTz<��"`"��q'��?M���ޒG�Z	��FU�XF�5ӗ�>?P��˟�r޴nO�O�1���A�%h2����J��'���#�|��'��Ovc�����U�9������-c�4�K�)�<y4h�q?�ߴ�?95�i�\7��O��o���HB��̝S��`�dͳY뎀������M�����$��@2��i�O����O �;0	Pԩ�5H��a�#����=ц���c�芄�i���R�۠��S���'��)���mZ��dx� ��h/Ȩh�
ʬ/�Q���ՙ"Jz԰����3ogb��R1�F���/�9#J�yRw)�,7�����Hgӌ} �O��rc�'�1���'�B�;}SN���+�ȵ�3k�(*���'���'�"��>aӄ��xkT8�' �brq�'�gyb,c�x	nџ�0ڴ�?����:(�ƙµIL&A�p<�3lPc 脳������49O����Ol�d溣��?)��S��4��(лT����D�'[��0 ���z����$&M��,�P-�6X!�4�%�Z,���g������;�D�d�H��� >3.� �FEm�y���&B{�q����OUl�?�HO�#<)�$����h��t�dܛ�	P�,���6x��W�!C'�U�B=�jT&��{޴xZ�FP��qs������<��k�
	��ic�a�f�L��H[b�1Di�8:�~�1"��5}��q��i(� %9�J�"�St+�'��eAqh�I�'���a�A�*lg�p�t��q���0��W�\I� �S���G�(�
A 5�#?q��՟��Ic~H�$O���zRA��8��Q�7 Ѩ�䓱0>�p�ǧ�LB��+icp���y��d �\r�*� �{e�q�2F���	{yҬ�+ۘ7��O���|:�"L��?i�'��{�zIH�ܐ>첵�u�8�?���|�ݠ0�V#m���zt���b���yDM���l�͟���Be��A߮٢P�
f�J�뀟����*#�Ӷ��)8 a/�,lu"�:"
ղ��iPph}����_L�@��T�O��ɏv9���Z馵
���|>A�l��|�W�. ո�E=D��1+�3p|��eL̯lQ��PY|џX���)(`7����m42z�顀f�:��7M�Oj�D�O���\g�v���O4�D�O���)`�
%�䐡,����2LV�t�o>_t�jS�`�D�2�I�#�t@+�i��aV-�")�,d)��
�r���XgQ'�ĵ�c���':�A� ��ۼ3q	�)�"`�����9֝)�\��M��T�0б��O�����$�O��VO�8h���$k�Vј Z��?�����$�OV�?E�O�Lp�`g�>h��J�;wC�YA�'t�"�>*O��'�?Y*OR;!�G�MX��v �~b*t�5�;J�Ȫ��O��D�O~�����?����A�mC�Z?8k0Dən�v|����Ж�G#4"L8�j~8�t:��֦L��i�s`l.��)VňJ��l��W�7��uD�b2�D wJ:{��!���]�~� �$nJn���P�)0r����'
�6mII�'R�P�D�1μ����@z�$%=��I���s�eHIBU8%"��<�<��Q'�$B�e�ٴ��áP oş�̓A���j��˫a�0���n@)}f����nyB�'�r9��\��l�&\��1+͒�8�ı
�jz�} S��3��(�C7�,D~���Bd�PX�G3r�ŢL=��#�ٔŎ�$#�Et����� �@��ak	wA�'�Fٸ�B�f��<ч�C�G�v�a�+F�V?��x"O�M�	z���F���e[�6��P�!�,�O.���ҦM� �:����N׭}���9���M�+O�@yqN��e��ꟼ�O9B��'�,Y��I K�T �)�d`11$�'?�e5��)I��jg����8*2<�!�ג#e�g�0�Po�byX�Q��>'���'�, ӠJ�J):��D*�y(�I��+�^-��$�t
�c� 5�!׵B�Ĕ�ӝ�r���OB�m3�H���Ӽa��p)���>>Ӏ)Jk����/�S�Ob<��o<8豩�9��@CU�'��V��2b��Y �X�XTK&I�34\}�,�^}��',�A,j䚔���'�"�'�6�^}Qa��#n��)!��}*4B���"h�s`d����H�,Pʧ7D�O�Arv�,�P��C� ~���(߰\�4���� �z�x����p��M?=��Fϵ'��]�<��ek�lػ/�n�����]�j�o�M+��S�|�������$�O�R֋�0^��T�Z%���i�O��-�O ��'�H����Cf.&�D��Q��3�4��|2�Oe�]�8:0�H.�
��@��.���r�7Y&��䇍3��L�$��,,J0K'E����q쎴j����%	�dp�����(�<�ڍ�ĉ�gԠ�g
�`V�|
b`�e��2���!]���:4�Ƽ0T�T��L�#y~�����:j�&-�bZ�b����� Mv���'p�7M�~�'���0&.�;��q#`[�����-,D�$����H�|q��nD�u��L�T�=���鈴�Ioy�c�oR~��?Y����>�H�,�2b��k�!�?���jB1C��?��O��1�e�;S`ހzu$	)B֮�X�Ć-1I�|q5̜�Sk��D�Xq!џhh�"�+E~�5H��޴UMd9!"l��Q��x���3�H���E��}l�$#�8�s�;�IF����O��mg <��du��85���h_}'���Id���ȵGz��\X񨂗O���.:�O\,���A*�s��I�h��ir0�C#u
��ı<�S��<���Ob�`������{`�H�/�����,h���m=��X��L)�Хs�ǖFnD��6�~����,2�yS�̷xg���CD	z~�CG[�D�ԁ�Nl1 ��
vX�	�g��L	1�8����W�R�B�2U�P�z<�I.�����ᦑ1���e>�2E���R����b��X��a��#D�`˵J�^�#�!)DJ���E#��6��>�3@��s���X���71g�yv`T�����KyR��#���'/��'d�I�&�+ HR<N���G�(;˄]!�^"2��Y��4�y"fg�"��	^��rϦY3�d�/!���#��K:tV^��,s:�l��%/d��E��>B�@�Oc��h�����y���,�DM
�&��Iԣ�f����<��L។�SG�L>!�`M�a� ���;$���?�?����'���X�
�\_�D2���6����=?1�4~ӛ6�'�l6M�|:�����K�d�(f�C���]Sƪ�"d���&���b�"�D�O2�D�OP��O������ՠhut,��oU�,OV` dE
��fP2��J>��UⰂIB3f� ��*�%4)� �8�"��o���W�D�Z�J��@�9  �H��Pmj�3ƋX�~oz�sq��T��Ox�sab�u�.YG��-RJ�@Ԧj��d��Aݴ�?q-O��>�ɀP�f�@v쀎AO@�HG���]�?��䓞��O���3d�#`�`��%�M�\�H���'��6m�OPAmZ��M{/�x	�5�@ԦQ�	�� ��/�:��Q �iC�#�P��U)�П��	�i�:������̧����ǆ��*�/��	�ū�,0Z`)D��cPt�c&���OL�r#6��,� �&��o�ʥ�K��r�		=�BX#�.h����u~�O����'����8)׮�u��̩�̽{!�� �c.��O����|�I��=B��H
 JW�=q�OP�=�'G�� Ε?B18��B�^��y�<�?A)O�!�Q5O����O�ʧA���������
T��#F6l�%�$=������?�TF�c$����LVr�D����i�<�'D�uk򢃰X�և"}Z���O"�ɡA��."��CF���I�?b�&+&vh�*q �.2����@/?�e�x��(�^[B,�-1Oąx�cEpȅ
�'A�5I�HE*t�4�3�N�]���1���^]�O~�-�C�FWd��A*���ip2�'Be�%g鈙p`�'�2�'D�0��|�pM�$�8E��9N'<)9bO¿-��8b�o丙�t�ޕ�1�r!�7���~�h�(o���I�Q�M��ƒ�~���q�9i�v�j1g��q���d�Џ(m����k*&ձ����v֜Pw�&�0N>i7V̟H�|�<����t�^HX�ʕ�zTՈ���F�<y�`F� "�HS0mVW�1�jFyҢ>��|�I>)��Y᪂B����Ʃ}R�d��� m�4�7gåF�l(�lqsje���x=��ke�ĝ�BAd`��Љ�4�x':Ta�"�G�8=�2�I��P��'�˔Vg�yz�(��:�ɒ�K1LT���I�`	�9��0+8H�����&e��D����O� oڻ�HO�#<�SQ�
��ev%;x�t�X��P�<A$ƃ�rL�����`(��p�&�J�I,�M����򄔌}�T�lϟ����J��{�	�?���S�$P#R
�h������U�������|B�c���<�$���\�2#�GӼ �B'�SD��[VG4dn-BbmC�`W�YK�����8���iZ�$R�I�[$���F�|�� K��İC�>!X��L)��1c,�I`���$A��� 4���o�������V�;���2�йn���L�	^���ϰ9�2D[`� �O'Vs�|kH�/D2�'�X���Ǭ6�8x�֥�KP2\�h�~̟��C�kC	D �Ь�瑟t�2 �8XP*��A���`����p��"�E�?�끭�,D�b��\=b�A��$׃hUB�'��>e��>1=�|�P�D%!g��Ѱ���q��H/d[੗�r	ؙ�# ?�N�Gb�>�'��a
FE��Z���v��($��ٴ�?����?����7��%���?���?��wOH� ��i�(�p���(VR@탕��+6E�a���7.E�ٶ�O}�'\�a�g�W�5�wdg��ؒ�c�HJq��(TOx \�v�@�T=R���(@���K��X33�Ġ�S�.4 ��������8C+�OX�$�O$㟐j�D����qcmʿ/�p�Ѓ�C�<�3K�"��sT'��!����Fy� .��|���������PΌ9t�82O��@�
	ޅ	��$�O���O���;�?����?�c�I9@b�ї�M�e/����ڞ-ښ9bS�H�JO�\�5�£x�ri�BK5�;$
��%�b#r��(�4tBF�h��M�d��9u�z���i/([m]���P���|b]/Ҳ���F�N��-���^�����!i��+=ғ�O�J���u	����Q+ɚ�� ��T�( H�(}�����~�XS��)��H���ܴ��$2A��n��H�I/�E�k2/>p���n��re�U�I��0`��ϟ��I�|ru�T�q.*D���ԳE�m��tH( "S�;t��9^����I�&��a��B^�u�p�!΃AT�0��E�!����/�x�\�	�Ʌ9Y�8���P�qOQ3�'��x*ʔ�D��	�hP�u*�°�"��0�O"�q��Tj��T�Q�E�Z�~4�T�'����R:J��u��H��J�&�b^��4J��I�ԗO���Jr�'�����i��C:B89�Ѱ$�~���'��"N�YQεJ�.{�$a�4��O�`��	wfبr���dI�)V5��dŻ9Gq���^�N���H ( �a�����;'��j�V����8+�`�9�'I$K�6�rUlA��ޟ�F��9O.�*�"`�1�,�&K��`h�w�<���� �[3^9GN��r��v�'�~�}b���(2�
<�RO:̀��嗴�M+��?���?A����?���?���yW�f,PPF!Q�nN��S� �q��HT�|��*��?o�'?��H��,y��,��ָp�(Q��mЛ.��p�'�}�Gc�јϘ�� �຤C�Ln ��J� ���3��'��4 ��'!��O����O!�h�?a����ɔ���aJ�+�<��?y���?Yd���|����?9�k��
��C�(`�Q�S&YS#�q���?q�Y���'Q��ݟ��'[����
	i��Ū�0[�p�s"/DԖ����'���'7�Od��'�bbB5s�s!���{h*	��E�`���� ���ѕ`�x؞ ����2<���ʐ!��z�hpK4 6Gj���B��88wLI�ۓU\�����:~ǐ���	A���9#F��ȟ��4o\��GxR*Ö�
�A���7�y{���"���2�S�Oʈ�0W��N5�1b5o$�9K>���i��6;<asB��<���?y���HS
]�w��]�!�DH�?	�m�����?�O ���H*}�h��y�j�<0�r��$�b�c��0<�rO�V !P/���Y$(@S��S ]�Z= A_�>]���IF�4"<�(�W�a'�?`"1q�	WM�<ٓ嗃@�4� M
�*8$�c�.L��<#�Dꑘ��X�	��%{R,ճw?J��IAy��u��7�O*�$�|��[�?I�ɏ!w��0�MB>	Y�z��*�?y���T����P�n�o�u�$��s�O>30�Xs.���L�i��Pñ�*bT3w*9?�t��:�	e��	�n��!�]V���!�Īo���w��%���g鍆��XK��2���iD�$�)�s��ƨ��^C�%"N��!�,J��a���ӱ{� �?�2� r�H0!�����㪕�*�~l�˟d�	��Iu�^7c���I�����۟��;�w��m������O���ۇM�q���ȴбg�U��7����S��~�"����	��<��@��(N�Y��.�%<�� B��bh���g&����ZƢ !�bP�� ��vI��P;�l�M>�6I�ϟ��|�<�7�E'��5���
P��h��}�<�UMP��`	����v��#��nyr�#��|�H>����r,.��'AU$7�`�QF)��?�` ;���.�?���?y��U-���O��dp>����ل$�4��`c-i>Z bFDߗg!h�A�N!d�x;���V0&�Ȅ�Q�PA2/B�r�Ivf�'7־(�'��-c@�q0���p5��� J�LVaC�P�$RQ��i"EU*M��i��Cb�Z�?�f���B��R�[�D9F�t���S�����ybN�!}���K�j]j�H��9������|��A�!D맭?�E"@�ʁj(�7,F<7'�>�?���DBh����?��O�QC��>(JS$��$mC�V���^�h��%� ~(|J�	��Fm�T�'>,ۥ��>r~��@�fDR���?SJ�J�O^.P��v���>c�i�@�T��Of�
V�'���g��� �P�E
gF�	�h-��%�OL(P��߶�5`Aǆgu<	���'w��D�;�(��'b�j��E�0�&#}�Y��C�c�ڟ����O�. [��'���w�	
�&�2@�гM��'�l�09�҅�1b4�L����0��;��8L�ӭ,ߺ!Y`� vL�m)�$��u���)�p�Y�PYV̈́��f�XQf��F"�(!"̔L��)������o�0�.
&��$#�	#:`���Or�}B�'ߐT�ǧ�-x�L����
8	P�y
�'6�9g���]_�Mx�M��*X���C^�O����T���(��$
�%��`���Q�i��'."���j�j���'Y�'�b;�x�(  ��8�6����LK$c���'�v9d��ӘϘ'~�u��H�s�[��0�	��Ov�%ӨO�i�G��w�1�1O$,���S8�$��-�8�z	���'���p����Ox�=�! @
G�2��v�`�d����;�y"��9|��\;�e�5mM�%����#S�	�HO�i�ON�I��&��2i\N�F�Ě9S0��K5+"���?	���?�2���$�O��ӄ�zhX���_�����C"��pB��3�r	�4��\�����џ� ��$n���!I](&T(h�(-�Z���JF"�
y �`����9��)�}�^͘��v�(�@&�͇]%PQ��BE՟��I��`�?��I\.1���$Ȑ,K�����=I!�dX�9̸��
�W�{�DN!:�'�6��OB�I
���Ր��ę�����"�\y�Ujbo.�?1)OP���OX��?Y�bt ��d�R\zM˟���MU�?;���e��nðn%OrAxҹ��CE�oRD�T��O� (��֓c�bц�D*E�I��'��+��?1�O@|��J��\���i�;�j �$�|��']e��ƒ*44�x�DI3l�
��>��Cދ#����!�=��ha�$ܞ�?�*O�X����<�O{�Sן�� Q�y��C�"�F�P��FΟ���:Ej|�ʞ#	�p�f��?E�tC�#nuC�Х4����I�����q ��)����A��˖/�'Q��Eb��J�Y�1�ѯcݺ��'������?���	d�� <8"%BT+��Ƌ�iWD���"Of��%M��(#��A$�쨡�����h�\����;,>��[�iS���\(R�'R@8e�4�Q��ِ��$V�.Q��t��
$�>D��;�>����b�nE�=���<D�t�"*nƴm�������%.;D��P��<����f�]vzX�7�3D�\�		�l�97�0�8n3D��8�L^�,��JXR��8�ϰ<)DcU8�D��'�[��zFa�p;�X�.D� ��]�*�̠�N�vT�-��7D�HIq�K?^���C�̗/u!đ�'�8D��8vD�?�RA��:0��]�G�7D�h ��C�d`:<��b(x��	4�O�|�F�O|s�B�`�uY�	-o�dpr"O�"GaKC�ļ��GA1<%|e"O���R�dԂ�ӷ&��|���"O�|y��	,⨰!˒������"O,`-D�ܕIe�ǝ8����"O~�AE��3׬|�2���L�"���	1`���~����7+�ba�TlF`�� �C�<��K����L[��`PbȂw�<i��^h�.�YKT�B ((���O|�<11T�$���C^@��]	���s�<!�bP�Uz����Ef,�[۴�yb*� }��ӕ�9�tr����?�&(B����@4��*�)����Ȁ�DU.��@2D��x�
ّ*C���ݎ$0.-(�/D���o-Pre/t�E�C���o�B�ɥU� PS�:Zru�6��4;,�B�+H皅I��6R\��g̔;�*C�	�)�U�p�I5R�Bi�h�'e�Z��ՎZ) ffU��&I�1uz6%O54Z�}��Ƃ-W�&"i�v���w��@[�ިj$�6	��e����	�_�|jv�@�T�쉻S�#ng��]w�\`�6e�V��j5@)墉���^v�xTy3,Mq�Ҽ3qc,+\���Bά���L	���qdƏj�X�D|"��5�?����O�݋S��Z��a���E��BH)OL����.U
�qS�B�U� ,��!+��'�ʓR4,e���e'�l�F)�� W��'�2���''���>�a�H�^9	I�C���$m �	�<ig��
sP4TC�E�,��rOiW�>ɢ���5j{d��QD�X�P�a�Oc���`�"(eZT�Ԯنl��p��^.�H�j������:�P6�
�a��)�B3O  y��';�����f�&��u�!��$}�Z �1F�%�2%��9�"��L��,t�4"� J���D{��1�!���n�3N<�ؘӬO�:�
������9[��z" �i������}��A%#�"h�Y��H��+���$�S�cT2�ɟ���>Qbc��PmD��C�/Cԅ�b��Cz�y��ʴ8,D��B��)�O��b������_����Ѣ��@��1?���Ɵ���x�'��d�Q�^+����@BhbػO�!�d��0�b��t���EX�*a�F�9��|2�����`4~}����x5����_<m���S&�O�A�^�L"���9u����IY�Q�����(��L��W3�J�D~� ��R��9Y=`9�6c�9y�@<ڑ�Ԥl!�Ѡ�AܚYF	�$��9*���x�-�O&���@Ҧ��u��� "E���{g��O�=Q���O�0e�H"&��;�j��&��w"!��gz `�#�Ɉ�K�K����I/�M�����d �{|����Z�}A�FQ�u�T�s�jĉ)�T�e�H�K��C�51r��:�u_ $1��%<�ĪHαL?�m���D�O�D�PB��q����/J���կ;\��q�R�j4�A���(~� lG|��B��?����O?쭪` BEƎ�
C�ݪ:ZU�-O0��ă� ��z"�!}�J�h���#7��}i�<�G�LDB`!��`J̤1O�zyOG�e��'�RP>� Skޟ��I�B��#a�
��d�Pv/���ɴ~��kի'~��h4�C�<���Z�'I�R����|:W�_��KD�5J�r%�ì�<q'l�+s�p�)�yT 
e�|�rGώ5}։OѦ���/� +� ib�k��h3�'�����?Y�O�O:�)� �JV���)�̋��>:�$"O��ؔ@�"r��Cj\0
�Y��	��ȟd+�nĺ<���r�֭C���ʷn�<A��I�d��6����?Y��?�x��N�Ov���@U;��qX�-n�*����W�(d�)"�N���}�eH�]���'��'ȼ�q ��f�)�l	�|X�*�J�0D�@�d�J,��O&���f�t�*��R���D�B�X����6�n��k ����Pm\���O��=Q�'Q⼃��^��p�`��A����'����a�x(�2�AA�G��i��㑞�S����'9�a�$�I�t�)�MX�Mf^mhC��O�P��@�'�"�'�B�a����⟈�'=�5�"ǆ`�@�A���{�XH@H^�T��5:���'�����)3�&5 vI1�H���C��m�}K����`�0C��(�r���蘪2��q!5IN��:q�A�
�^�O~���'�Ҍ{T�ȼ7�x�uk�4TL49c�jm�\Ez��	�����+��;�p�����=��'�B��@�Xh	ڰ��rT�)O��o�ƟT�'l���'�'m�[�)��=^�=��jO=*��A��'���� l��p�-��x`z������c�ou`�{f�C�l��]���	���K��Q�t'��ħj���3	�@QR=+ףB�-�G|�Z��?a%�ixF���HXbO�8M��� �,�evf� �]���Ic=A��I�fM)��ɊsϮ���<yC�iXt6͑�]��C�
�(�8�ӳ�ۈJ ��?���?����?�)���n)�iY`
 ��ٱ�E��WS�y;���*��1O8�n�z��� ���+čf���x눚Pe���B�L���[<���~��Ö�|Ԃ��T�� ��G#Q�c����'�*��50Oz "���~:�'�?	�'�hɛB͖7�<<H�BS
3ؘ��@�ӕ�-�O�����Oh�	�Zݖ�s����Eʙw���#�A� 
�@�wr�s!�	�P�	du�̓�u7S>��˟���99�X�S�Cn5zJT�(��C��I����	�W�v����<�3��wnz�٢>O����ެuYz�"R�X*?�~�j�@�O��B7�' b��JZ���u�P>M�S�?�����+�@��W ��Y�`�2��<Qam��l�I#(� ��I��?�� \LnZz�6�Z��7V�D%k�Z�Q�j({���M�'��X;���?��nK��Q>��6V ���WM!ʀ[d��9'C$tZ�D�<yR��ǟ��	��u��':���O����{����'�F �h�"���PC-�66}��m� �?iPb]���ɶ4�t Щ��'Gmf�����)R��T"��`L&�պi��b"1OD�h5c���oZ�?Q�	��?��)����f!	�1]1h�ƞ�TIYp�	޴Tf�xR����D�?�m��(O���L_���2��3=e����#GTC�Ʌ�����m!��a ��i�(7��O���?���?���?���?Ydh�6-
����U�Gռ}hq�7*���'8BZ���'br�'?��'Y(\A��3K8 JE��Ȕ�X�c�f�D�O��D�OD��<ͧ�?Q�j?`=jl��*Eh\�R��j@��Ӱi{B�'�B�'{��'F�I����`�x!�����y����M&�'�y�Q�|BF.R R�C�̖UG���@m���O\���<�/Ođj�	%yz�Lx�DѢۊ�K�"z}b���O�|jů�F�H衣E6_^�%���u�<�GcNg��DK6�RG����V��p�<	7��D����9e�
�i�i�h�<�v�!�����Ϟ&�zX��*�c�<�c�d���)�S�P�"B��]�<��f?g���ҧ!�%T�@�ǜV�'b��'��'�r��X<�0�̑{e%�b�:!�h7��M;��?y���?)��?���?���'mF��!F�	A=JD��ρ+�P���iB�'.��'R��'�r�'��'o�4Б�"(k����/�=*�!��e�B���O���OH��O��$�O����O�������wC|��'��{�؈��C�M�I������4�IğH������џ8�p�I%&���b)X"~
���M��M����?Q��?!���?q��?���?9�䛄:i��x%-�R���Y�+^:'��F�'�R�'Rr�'�'�B�'=r!ͿI��4 !��&u�8�%���>�T6M�O��$�O~�D�Ov�$�O���O��d��ݬi`p�� /�&
P�N�H��l��t�������ʟ���؟8�	⟸�I5"�B#�Ԇ:� `�I֕C"9�۴�?����?����?A���?���?���Wh�� �
�
/���Gn�Կi�'���'��'/��'�"�''$@I7g��C��j!P�·��6�O����O��D�O���O��d�O>�D̎%p��$�?Y�.`P'���P8\m��P�	ğ��I՟8��ꟴ���@�I��\䄟8q��H�g)Q|��"�4��d�O�˓����}*�.��.UF�1�FLE��X�nwӼE�����ޓ�$Al������p��5qg-��@'�`�gi��?	�4�y2X���b�2�?K����q
@�[�
_�XŮ-��,��&��#l>�ў�S�<9�G�U�z$ M+2y�l�Ŧ ˟��'��':�7�ΠHj1OJ� μ� ��{j�Z�IR;L�A
���`y��'��8O�a�:��ۡe�����=d!�'��%ɶԪ��\i�O�ɍ�Vt�!�$a�@i��F���@Ǒ���k��<����h��DJ��})��$U2���U�k�r,v�6����@x�4����d,�?wOtH#��E�jf���aI+V�d�O\6m�O^����ھ �	-f|�gg��~�뮟�+^
��.Zc&�����9;ў���Wy"󉕷�T�A�.�.+J��3L�5]/�	<�M���X̓��O&9"���q�1e���tyFO�<y��MӜ'Б>a0TnO |���p� O�b��դ��>��($?1S��5(��O7�45h�$g�*��z�F2$��f�ʀ�ѭmb\�&�	�~w���=��D>9�bK�fhs6X�3�P�+[f�s���^{~�0��o���h���0((9���ϔ��&)�L����e��8{PH�e��z�J�BQ��)nD.�(󆇜|��%C�F�4c8�[�M�Qʸ�i�	[5:R� pGA��x(!�L��u��u��G�5c<��Xڜ�96K	��U����2u�p �C���Bc�� �_0�|3T�
��q�"�#�r5�*��\��`���>ye�0� U ���;wt� ���@~��+v��0�"
#�4��$�t��g�8���� N�OӔj'cX�q�������Zp��̚�x&���G,4J��0�.
�b�D�+�dW�M�t�
-��Њvɑ�T]<�k��E>O�%i6 ӶO?�ADP�8�p$q1b�	tsҥ���o9�-R �ȍEP:�P�i�b�'������$[�(��k.@�҅�'M�[���I�0�	�s>��y��� 
9�7
�)�aq��<�?����?�*O��Qň�¦���֟<���? ����3l0�_	HS
�iyb�'P2�'�@�[�'��'��į�~A����/te��SW���=��'�LUr�7�O��Ox�i���DνE��I�SG�NN���C_�h��ʓ�?�(؂�?I���4���'E����#ɞ��(#
UA��	�%�ٴ�?����?a�������?Q��f�,ر�E�	�́P��$��xC��g�$����?�(O�i"�)�Or)C�'
�R-�h�9=�ĜЅiC���ܟ���'*<,��۟�I���������v�ƳJ��%�0�0e�`�A���	��AnU�mI"($?����������T��d�+D+^qA陷bX���I�H��*��M���?����?��V?�ϓ8H2My�� �i��11ui��eD��	+8���z����������h������ɻ~Ir� L S�`b�����F<r��M��M���?!��?i�R?I�'�c�
=��	��_4.�f�
 Ĥs��+���M3��c��`���?1���?�J�b�f ���
$�����|h�/ε_��'��'���'��	���H�t>�PjW��1�!Mٴ'f���ܟ���2b-j���ן���韼��j��M;���?q�i
	3�d1���Om�0�@`Q<�?9��?������Op�z�5����j�tń��~�~}Q� �$u��.�O����O�d�O�#!�C����������?����� 2\}"��ؠ���S����	Xyr�'�N1z�Odɧ�4������C�<N����BI"u���'8�,U�Y�6M�O��d�O(�i�F��B7U/��(�aO'R��L�Ci^&p
��?�4c:�?9����4���k����Q�k,�KQkJ� c���I%<	��4�?	��?I�'�Z���?��2A�aFZ�f|�xd,B9l�����H�����?�.O�I �I�O��v��bR�+����\���c2 G������I,G�������I˟@�I����d�	�"7�O�g�NMф� �I��h�!K�>�&?q�����I����r�ȅ�&�+��"�>������cR���M[���?���?Y`V?�Γx�p�	g����j$>,x�'�${�'���ןH�I�\����	�?"�6�3�&X�z��8C�8�4�?a���?��G��dy"�'1�2�-Y�:
0���.ns8E���y��'y��'1r�'��'��Yj��mӴ�Ѭ��X�bQ�c`v��0�U��O��d�O���O���<��F�r)ΧF ��)G�T�&LPH�0l�*���?���?1��򩆧J]�nǟ���Lļъ�%0'��l8r�K:E�\�I��@��ƟX�'�b������'4��˖Y*�����%��v�B�dD�b��'�2P���M�0�ħ�?��'e�����#��'���@�I>�/O����?�*UMO�[�YZу��Ym$�3�n�O�ʓj��	��i%�S㟄�S���RxR��6�^*��<�E+r�0�'y�,^��#<�}��Q�B����[i1JQ�����aL��M����?1�����x"�'	��I�^)>n�C�r�D���'p}����S���"��oﴉiER 6��B�����M����?���sE�x�'��8Oҁ��;dřC�%����Đ65y1O����Ov��O�WNd�8X�H�R6`�9�� ���'1� �0b� Of�D�O֓Od����@�"3ȸ@e]�_�KԇA��I��b���I͟H�I[y2#��hr!Kb*�b�����3�z�J J7��O��0���<!�n�7m�hr�"��fVYҀ	:���<)��?������N.j8���(30��!6lY�m ����(�T����?9�������M����F��t��a��Q�򬘣xl��ϟ��I����'-���B0�i�z�01T�S����BW�fk���O��O��W��4�=��O
=R�I �H,�0lb�Kߟ`��ԟ��'n
���4�	�O���:� ��ˋ/>�8p�P)�ܵ�E�|bY�P7�*�S"t�]�VU<�� "P�FR������0�'��8	c��˧�?���,�I3.Щ!F�?�|�3��ʲn���$�<��Fz���O��Ed X��t#��x���i�zܚ9�Ӱi��'��O�b���=$���WC(+�P�۠-���C��1�S�O���&m~����h�<i�W�0'�6M�O<���O�t���U��?y�'�ԘZ'N��}�&��U�� ,����b���'���'I�N��mREΤ��dR<.0
9�'��ߥ/� O:�$�OJ�$�<���\N�P�>A�P����ӆ2�1O�$�O\�D�<Ab���|�zL+�NJ�O��`Iӥ���A�x��'�'��Cy�P�W�Fػ!�8a�D�6C� �,A�y��'���'���@מ�i��v�m����=\�	à���B!�'�"�'��X�P�'02���O���iV�Pj�j�S�͓-5@
y�+O����O���<4a�:A܉O�~5*�� _���Bo�>ahF%�#�'|��'���py�ҍ���O c�ʙ F�F!�Ɵ[|Թ�$�'���'��I��	iN|����R�*���J��ίV9n!h2�W0����Ő>���8.G�����TY����0���'@�0�"$�4����O,�)�Xy�����e�A��v���s"�<)Op��U�)�ӑE�H4@�G� 8��� �L�-3p��M%{w�l�˟���Ο���$�Ov��aɃ[�|�0mÌ[�6��'�O�8��)§�?y ��	�� �T� �����rc���' ��'�@���,�d�O��a��veB�&q�Q��Bx��л�i �	�9��c�$�	ğT���1���6G��z�c��H'nt��I�5m��ē�?)���CFN@�Qk N��G쉞E��Q�.O�C#�$�O��D�O˓6^�ť�f�N	#צ�*|�bL�<_�'�'X�'剼��R ��Z��YKFm�Q��eQ�#�	��d������'�v,R+��D
�m ��c�d���={a_�P�I�P&�T�'���'h�aB"�%��a��@=s�.O����O��d�<��D��*?�OH~���iV� AҜô�+qeh]p��'�|�Q��K�6�	�t&��#\�s@�xU�4Y��D�O��$�<��R�=7�OX"�O�00d�\�<A< 	��>m8�;��|�Z��Ņ3�S��.(�>S���D��[���'!��b)t�Fʧ�?���,���>Ĵ�{�bԵ�*��2(�T �d�<��w���O������969)�HK)'#p����T���ie��'��OH0b�|�q�X���쀖NHPA8@���8a� �S�O�@K�4
9�!�N�ph�y��;^�6�O��D�OU�$�V�Iڟ8���<��;J�4}���
Yx4ђ�z��v���<I���?���wW�k�ü{�:4kQ��o^�M����?v"̰r&�'�2�'��'�t��%۷VE�2��@�xL�FR�	2 !�ܟ(����'��8e��|7ʼr���,0c��Ц�A�T��O��D�OܓO�ʓ<<\D�����9t�j��#~U��YW��F��?i���?�+O�@$f��?�0�-ۆ8�~8��m�0���A�<����?AO>�)O�Z��O4A-�;:K!*&�Z3�:��Y��������gy���e*�����4�ѷu�<Z�oI�J�va� "�O��(��<y�iK{ܓ0�J��B*��L����z>�e������dy�T;lT�.�D��H�:� ��%�J�q�)��g��x�$��<�%�B���$��"�Ԍ��P /9.x��ם�?!*O��[�𦍔O���O0�˓U: xa儕:�tI�� ,�p@��Wy�攳�Oq�������80nE��x���H��c�'�h7��O��d�O�I�m�I��,��`�J�@�ѕ��/-Ap�0BBӟ�"2�S�O��AD(�޵H�lD�6��)^�6��O�$�ON�!k@C����ğaF�[4HJX��E0q(����w��\�Υ�<���?��hb�Y鷂�<w�P⋍^��{���?a�	�\��'���'��[��q#��2�	�tϤS�����Pybf���'�b�'�[����*�$ >R�E�ީ8���&T,~��}B�'z�S���Iɟ�;2l�o�$����=N~�{t�PhZb���Iß8�I\yr�O!�IV:z�н���w�ȠQ��]��IǟL��C�	Gy�'T��$��VA&�s�@�0����X�2��H�I��̔'*ƈq�')�IH S7H��c��<}	�Oܾr ���O��O"���O*���O�����c�G��ᖣ]�8a�����]y��� q�������Y�A��&q��X{U� �9=�x���/���O��d�)/����Ӭv���x��%���ˁ��*>���d�<�Ǥ��K���P>����?�Y-O &L� �4��qL�ps�ŲU�'`��'M�q
'�'gɧ�O�1��gO?F�����,�1���m�ބ�³i���'~��O�~O���?� ��c�:'z����OA~��W�'H�p�'�ɧ� �d:8$-K�K�	c�܈hbF���m����I۟X�v�B�ē�?����y��,(��Ҋ 5l��`&�8�?�H>�GG>��'�?Q��?�0.Q&n��@4E�L��@1�?��� � }�s�x��'`"�|⣓:���y�'�_r��Ã;g�AȖx%����ʟ���~yR+�r��=�3BI3U6�
ட�k�4,Y'9�	��%���I��b�2�� �r��]�Ȑ'횼xkV(��pyB�'���'�剛XU�i���o�������7h�H���'l"�'�'m2�'�
@1��'@��#�
�)4c>@����Z���3[������t��ly��%^P��^��iN�M{�����%X���O$��9���O&�M�<�@�V�a �pFȫV���sW1�?����?a-O�\���X�ܟp�Ӊ<a݂&� �� ���9_�'���͟��V
v��$�ϧ4��ض�!w��L�5(��%�B���Ly߁+��6�|��²T�(`��]�4����6�lP��K�O*���Ov0č�Ob�Oq�T��ԁP�q՞�T9:$\10$�'>�Eh��i����Oh�D=%���ɆK��-�<�-�uOҟ@�I�j��s�)§�?�u���d ��Y9m�:-�2�G�9����'[��'��Z��4�d�O��ds��Z��	 F�Y`Wf<1$/�O:�O�D��n1�I�OX��v>�n	�'0����BE�9b�`��O��$��lZd�'�d�	���&�`�̇�h�25��*���CI}y�����xbC]�>'a`Q�/A�	C�%x����&p՘��E��m(���@�P_:��ʼT���D�Ol�d�O���U����:5Š@8�Q#�03��S�cǤ! ����OL���O���/��~��j�s$8�����Cܷ-������'��'h��|2�'D�r�n�&d-�i� F�U6F��� 9gD���ٸ1L�:$��]2�a{��<2��=c"A�I9"�y#<����ՠ Y��ۖK�*���`���~X؛��	ANa{"���z� ���Y.�SP��&
�1�m�7r4lp�K0!�H�#GM������Q��Q�ѣ�2$Z$�whқ*��&M*'Hb �1 ��?�is�#��DZ=X�a�7X���c�9Zz���&Ј
.�+��?��+C��;��E��G�!S���v�'جU��f��:����B�*�?���˨�#���?!�O�r��CJ�1���QBV0E �Q�7.J",�&T�5��p��9���X<M�џ��N;<TUghB6U�聋BG]�ؐl�����!jv�^.Xՙ�
�?uN�#<ɗ�	���q}�&X�Av��j��R,�<b�aԸ'ea{b��l�`!X�#�t� L�$�[*�PxlF�ZZ@� ��o���YsP������d�[1��mğ��Ih�b�³irNu��o�	U�N����o��R#��O���"x��p���r���f�П�'��i�5����fE#G�(b�ܜD�'cP�p�NH�)AB<k��^�C�8iue|�\\:���?�h���W��������.O �:"	'�"WY�`2��)�&z̚!ZH�7"�+����"O�A�j�1,@8<H�a �@��M[��'8N�<	�I�=f ���D]#R�6�Ò-��7��O����O*\d@{ ����O����O���09UpA�r�C�aڼ�)�1J╒2�Z�o:���	S�Ġ�3�3��,,x|�G���?Pvi`#e�Cd>|��+Ng�X�P㚟U��Ʉ�	�
��O?b$A�a޵b��C;__fm`F%���R�9� @+,��ī<���ٟ��?!�>ya�8Z��
�M��8���ĎE�<!�"&&��b� ����(TG��u�'!|6-�O��F�@S�ԙt"������b�A�(��`b��'�B�'
r�t�����PΧfd�a�R��-�8�	���2a��R���a#���,=��iPV���r�7ʓ���Uȋm6`��s��v�H��nK�h� $�e���#)���<�t�u�/ʓ_�@����δ�2���J�Jn�ٴ�����	,t�J�{Ҏ��8�Y��B�ɸd	�̛ᩞ>{���Hs�L	?\��X�޴��%���Q��iu��i��$��D� (��4�珁&��ec���O��!^x����O��S����va��6��e�+�$���L+L����
�Z�u]@�F
��7GČi��G�wV YK�D��d�RX�T���Q�l����/vh�C5�	r�&$�<yu�	ϟ�M��%��?�
�" V�bC(�qp#'D�p�@ب �M�R�U�.��ӆ�'��'�ˆXh�+kB�+ȢE���*�E#��^���nƟ��I]��J�,��焈q�`�PѨ��S'l�DC�0ryT��O�Ey�� Qv�قTቀP�N�|��΁rq`�sX�)[riͯ(���R��x���f%���ˢb�0�ٴ_�z�����+��I�4��2 �"%��m��Dًe�O^m� �'%�7����i�IS�'V����+R88�k�,
�L��,�=���۰<y�3H{�� �.+4ѨQԯBl8����P8��1�jG5D�.ك�M�-H�����@����(B0
Ѐk`��IԟX�������Öwu�uJ bˇ�2(K��758h�<qq��BX�0qt�E� kUBQ�a��|�f*���3���� TpD�X�h�x��Q'��w0���CE	��s0��)�3�3]6zU�V� � h4UC��<!�$c���*(R�Hځ�_+[�*�����d�	-s6���E!A�>�|ЂsOS
5��
�I^>(�������?I���?aU������O擷N��uRw�6�x�A#�Q��Ң�6�h+D�WL�Xs���	F,�w�p�C�����%e�YDHp��6t�a��O���D�2Z���K����W�C7�!�D d�m�$ĕT̀��1lɦf�qOo�f�ɴE<f]
�4�?޴,���/͛HvѨ���6"�X�I��'�BK�2(W��'���=�b�x2m��O]��pDD�e=�!�������<��g�<d5��ۓp�H�r��<a�X4��I�%�H�d�q��!����U��t�4�R�:h�!��U�[�,q��ح2�@rp�-�w
O�!�E�ڂ]�-��e<"@�Q/S�gĨ�O�8��|}��'+�S�mτao�?Nr����0-kt!��%�p�(�[���?Q�b6��x�y*���7~"e�'�O3QT�*F�	G5��%��˖�ڟ&�b�b?Iz��F !��D�G�@���g�(�֏���'�B�'����!�6nΊ�89r�ש:XDQ��$�O�����f8H�5a��b��x%�2!-�xҎ(ʓ8���F��.lp�+#���ti�1�C�s����Oz�$�9���Vc�O$�D�O��Dc�mۡ<:����2XL�d�-h ���\��B��:Y ��$?�OQR�H˸"�����Ŕ{�x��ɕ�q�jD*2��Y�����.��m���j}�'(M�A	\?8n�	�p�,͓�$V���x���DJ�K�.��Y�n�,]��q�A�62*�I`�یi�
�j,O��=�2R��V1"�[�����X�r'B��PȦ��4��,8h� ����d"o3N᠗�J4\D�V̎�E��B��[7f�@��Ο���埄�_w��'��鉀-F��1a�0Yjᒐ�@�m��O�<I� ҭ8%�,�� Y�2��HY��Ȝo!���,n���u��^.�Y�0��Q���?�c�'n|$��k��V�t+�&B*"�
�'�r!��U ����H�9�(�(�{R	c�*�O��iQƦ}�	�a` ��8w�d	�d��7w����2��?���1oti+��?�O���8���o���[!���BT�[�+Qx�剀=c>����](_>P�f)� M���)%�'�,|�����y2lX�j�8��׀��w���ȓ�
�{�NT�!_�0�i��)
��zƉ��'�'u��R�Rd�k�蜸��\h�m���i��'`�S�!��o�'�e�0�G�N��%G�S���+��?�
ɛ:[2(8v.�(��|2��b�ZC�J�t��H�aH�	5#��x�&΋3ި�e'�n�ؖN�$1J�� ��,�2�śG���#���_����bn�w�ɪ����h�)��&�x�`����h����N�C�	WV���ԯؙ5��x8�㑨R����č@�'����DN9�p<YQ ՜E���z5����ş���!\�@�MIޟ��	�h���vpy��" Z�	����lQEbGW̓-�����/�\�v��},�C�2� b����+ ,O"�0��ֺEF�x0�ɦ7q����/�f�4u���)�3�$��s��i�Ao\�N�BР�%E�s!��� ��Bi�f'r��!��3u��52���K��0z�\�#�}O����O��4C��`�B��-���?	���?A3������O��D�[�ju����]����(X>9��E�-[,��=���<#Yb�C���%QRU��G^�1@�t�¢�%"<(�r�X�,.��R�Q�U#P�24��'� ����0�'�b�b�����<A��?iI<�@IW��)�C5q�����F�E�<a��.a��H� t, ����'�7m���'e�p`��x� �dr�4�����od&�X�%�s�N��	5a�ft�I��'L���	g�� <��G�Q�	���F��\-���d��Dw�OD�ѤOX"L��4K�<g<�b��'�L������_�]z.2�Yb�� 4�6a�ȓ)s��d˞3|F�@�� �(���F�N��%�`T�r��,-�1*�I"�	�88�q�ܴ�?1���)וv}l7-Ro���@b����֜`�"=�I՟��n @(u8�Y��aH��/��I�~n�A!G^!q�	�bPPb��l�ɱ	�4����m�8��b��Ms��߁|^�xw���>1͐�,�b]��Sgӗ]�����xҪΦ�?�Q�|��� ���rɳyD��竛�w�����"O���H�z�4q�k��vV-��'��<��[(���.OdN�1���Y5�7M�O��$�O���6��u#F�d�O��O�%�.Zvh �R��D#z��8i_*X�f'J�L����v �3�.�3�dN]L��"��E���)��9�f��G� 8B\S�/��h������~/��O��&����G/z��m�Gb�B�"%FW+u~�OL�"e����ēq��ԊԦrv��B ���܆��j�Zs�C)�}:�Q l���O��Dz�O>�'h<|xSKȍF;���-I����F;�N���C�O��D�O��d�ͺ����?��O[2�BW�[��ҠY��2t���jR5Fe�	+���g�P0����#?!)	bb�x��	/r|D�`�;D���h�G@�}���rǥ��G�u:'�b�4Z$H4��a�I`�Y� jMbƃ@�V��̀�-�şX �q�L�+�
n$%t&�)L:�O�Ouk��vh$�i �9uBQJ�����U&��Z�$��M����M���¤;�R��P>$p��&ټf�l��I럘K��������|r�ȗ���5�	!L��قgR=	�܍��H�#UT�q^2��u�'�:�SRETQp�Y��X�3�������[��M�hH�P&�\�V�pӏP�A��=���Ɵ�%�(7�<:6t�UF��>�<�	��1D������?��YdO��T��.%�4���S�W���"U��\�ѐCĆs<�&��b�E�M3��?!(�ι���t���@��7��I7�[5, ���� �����IW,d����N�����pf`8Dҟ|�$�,�pe�Y=G����E�T#Z� �'� ��)q�:�p�&��"eC%}ɞ]��T�h��$B�Hh�0zdŏ�qB�@6/4g�E&�����O	'�b?�r�D�Bc�1fGBy��..D� ���ۼ]0��#	ã(�b!��� �hO��x�'8s�ǌj3��*�.߬S�US��R����۟��ɖg�p�im�͟�I�,���6�S�bZ�L_-Ԭ�.*W(�Wi� *!�7���q���
��6q�6��|�H<7��)@B&	�)N �qqƃԼFJ��R��B�L�T�lO���$�ND��h�T�P�w_(y�蝗LXf��G�(����DQ�	E� ���x/��Bj�:�� m�`�cV�y�%@I�����ɮ_�\�3����	,�HO��5�d_e��8S��P$L�@�T�%��Ekf� A"�t������I�@[Zw��'T�IQq��H2DdBI����l���sDOr��7�K�s>��7 t�N�� �F8L�!�dK���P�ǧ�3HH��a@��z%Ё���'�a��#q���A���:r�j���I��yRB2 ��ir���f�F}!� ��'\@7� ��S�;���nZßpmڿaXR$@4�#)�����ǧJ�|����?q�-�*�?�����D��8eݪ)����2x��}Ktc˴��h��JY�Y�nA�6��X��B��ɺR=�a��V�����q�9��Jc��>��bF�0(��T���E�a�VAZ�o7��M>�AZן��M�Hʕ)8r�ӣJ�E�J1�s
7D�������DA�g�?=����6�p	s��4:y������8u�л��Ƈ�I'�*� �M���?y+��Q�-{Ӱ]�%-�]�|��Б����E [ǟ��ɓ�؍x�� k$<���+��m�v<����'\����A�{��F��G��'�hh�Կ�A"f%n\8�f��˺���L?I�,����$��a� Z���<2�O����'"^�O��>�����?~�Jlʢڸh�!"O�rD.Բ���w`�0¤MA�'4�<w����3��̿\{���@�ءt~7��O��D�O�<�%n�Z�L���O6��Oa��v��@2
�6p���@�ȟ�c��9tN3,O"�h����.��YإK��+pࢴ�B*�ayR�Y6A6�DBF�[�J��C���y�~b��c�m�Oq��'�xU	�O>9B��׍�1���i�'1,1D��ad���v�]�u��=�O����4��O�}��g_:.�N��lA�Q��0v�>xd-��Eݟ���ޟ��ɽ�u��'��1�n-8�^,!��Mr�L�*7H`�B�U�!�D�7i����F�
"�m{���i,+IJC<y�O�nO�u"� M�K�hEPAoȓ~���I^؟dナ1��<`D�բ0�(8�� D��Kgˈw�&���mϓJ���f<���'�A(0�|��$~�z\SA��4��I`j�2%��Thf�����"_,��ǟ�ϧ"�()*��K)���a����&���+0�-��E�<�%�''�LzW�Ɩ~���f�[F�� P�Ş�:m3uI�`�����j���h�ê*i��L�=Y�	���h�M�����B4*���I�T��\��@7D�� 0 �ҲJ̨X���jة�
O�	 !��]H�DA��,a.����.}r�Oz(8A����	џДOP��#�i�l����D ���!�A
O�X�t��O��D�-�Ԥ�WL�Xђ��m0�$��O�S�l��YucW	,^pYvE�+A��O� ���J�d��!�����¬`o$\\]ѧL�;
0V���X��D]�ď�,I
�y����ēZ<��	���S�'vjyZa�I⽰���4��,H�|a�E�B���8��E2|���I��(Oh��`ˑq:YH��ӯ*���Њ���Mk���?��X��њT���?����?��߱�f�_�e8m�e�	/�$  +X: �qE�<l!��r X����L<Y\�1��Aʇ�]�ܹ�eI�U5�pM8,��`�vH[�XLp��G!���S��X�3�x	/l�%��BL.��PgF�9x��<�gF���>O�Y���x�U
!�HR��;V"O0�0��<B��b�8���P�>�2�i>e%�l�&e9r'LtiSe�|�C`¶Z] 2�.�?!��?)�}&���O���u>ih�R BB�[ ��Q�nI É_}���⑨3�pv,[]x��UJ�2L��iq�g�=7��U�X�%�8)�W�^>|FHr�i��8#��c��}�L	���!�I3|=֭C�"A� �����jЄ6������Ol���I�M*�P�&o\�ℸ�6%X�B�I�P�^���B���)q�Яl�`�hC�4��E�!��i���i^��@�D���X��
Y"p,�%��e�O���0�����OF�S<�h9r`̔�I��cD�D��$��1p3���e�S��6I��)É��O =���4%�di9��^�}���uGѠH�P��pa�	T�+Ӆܟ`�����87���c�>�䅢83��>}b�Q�cK�l�"K��W�±���E/�yB�G�U�l���U7L�`�ŎN�(O��=�'a�V!J'f?�V��1�ԥc_XiR5M"��/�b��%�i���'q���o�7�aU���D�Ȥj��B�`���?��Y����H�

�������G��*�O:�S��~dzS'��Z�vԩ&m�:#�rO�Q�Kگe�Ac���{	��g�X��v�*d�X3 \����)p�2��e'Rw�|�EUi≥����j�)�S�x`0���F�L��C�^�C��0|���cW�q5N�!ǮO#'����4�%Fyb��,h���+��5����=(�nZ����T2��@8=/2��ڟd�I��΃��pT����<��qfw�����,�8�����O� ��P-�1��'���z)ܢ/R<�`FDK8H$27n�5���cv7\li�H?o��A�o~��� �l�'M����F�òWH¼���5�xJ��|�e��?�}&��"M�)��q�N
=*l�1�d&D��p���0`"�ITi��E \ia&2}bG-��|bH<�7�հ,<-���r]��5m�{Dj����
�r���'�B�'0>�]�����|����9 ���,��DR�._;��d$k��5����0�Ê��F���z�
��G�,���.9�^�ӲJW3>�~ ��M�<�`)#�{Ӳ%k�@�=�qO�%�r(��s��Q��*8��� .�-�RG1�O0�cK	;^<�!�Q)G ;7"O��Ѩ�eK�E��鈴K<����ڦ�'�,��	��Mk��M��D/3��	�G&�O6��r�Ҽ9�B�'�T���'�B>�T�����]STu!�ߧ)��Lg�0�!�D�����}��d�/��1���+�N�-.x�1�(ԾVre�w�ϰfH`��1.�9۔��C[&�M��ɰAZ")�=��d�៤�K�t���NUr�9�b,uW�9���*D�H�o_�]D�|�B3����D'�x�O��&��Xǌ
"B�����xB��&�xb�aJ��M����?�-������w�,�;G���XU�7�[�Q�F��G�����I�Y|f�5o�"N�HZ��ԓ'Ӛ3����'a<ԉ3�)�����\�q댩$���g�q��R����Q��3�Qúk6��O��d�Ӝ)��@��(�PM�GI7"�Oر���'�F�O���G��;)�NA��⟇Z�J��u"O��y¨ٔD@%� 
P��M�t�'��<	���` �q�7���/�i������7-�O����O�,�������O���OL̥n��{���%��ITO٣,���g��&G���+�S�p�J��l,�S@��J'��Y��(J$j!$1S�`� ��XAAI�]�����o���@�D���OY���������7bD���̀-t :dy!!ݮ.oD7M�Iy�Aˋ�?ͧ���}​3=��v�J2D��|���#�yr!ԡ	�T���+ߘIJ��R�� ���HO�I�O��+|v�ʄJ��]�R� ��ˆ
$�RAN{-��u�'�"�'keݭ����HΧjv�j��_�"Br��'�	EY
�(gI� �M�1w��شw8��ڑ���A��x��O't����lʐQ&Lcv'˓E�f �U�M��M{a���i���x2~�
2*�O���F�(8�Ԥ��(�*Y�����J`r�m�Ql�R��Mq���㲎܁(�j}�6���0.�f�'>��� *E90dצq��CfA|�ɳ�$QѦ��INy��Ii��6M�O�6��7c�&���ʚ�e>�ҶE�1#FN���Ο8���4�	�|� L�*�څ�*3��C���DX=C��Z�tK����#�&��� ��ծ Br�<1ТZ�t%�y��a��DYq�D�(0J�Z"n6b7��Sg�5�\){��4���<)�����$���k!'SF�7��+tuN4��-8D�X�q �/���pf��t,�+r�7�8����
Ρ��j=a����u �%A�}$��t씃�M���?Q.���b�f0�T�\(�=�)I&P�l��i�џ�ɗ\�J��%��
);�tو�/I�d����O�cƋW5jr@�Ԣ�#m].��M<��/H�G���adI�W��e�����Z$3Wk�|��@Ћa��T��!n�(M��F!�$� n��c!�"0����8�pA�d\9/�d�u"OVl !�ZQh	JU�.�=i�'��<��K�`n�i&���r�N�����p�6M�O���O!`6��%i8���O"���O��{^�A�H�x��ÃJ�7a�l��� �Y�$���Ƕļxs�-;��m��@/!��HS��)��%k0�	%L�LH#�F�^>y��*,@��$�I)}��J���q�	4oL��E�'S�0c�:���Oq��'"�(���DI����̑?����'X՚#IS4w��0��ݒ
4�I����4��O&iQ�
�H��mO�u3�)S�mw�t��wk ۟�	��dӊج��?A����*"|5��C��?��a��ŗ0yl�sZ_]���P�ql�y�W�0#���T�S)rV��6�K�N�#���Hx�w#ՒVT ���P�#T|�7�W���'$\|H�'U2gS$l%@Ŕ�RyS�·�?���L��P�өI(�8@�/ۢ3�X��ȓs<��w㒋�"| ��Ld.J��=���ՀY�4anZɟ m�:rX`$�G/��W��0t�.������?�f���?�����4˙�`�aEN�5'r��e�J�t����&C� W@M8@�
�,�v��Ą�%� ���`<�Yse�2�"uc�#@1�"N��L�HQ�+�Uޢ=A�B���YK�����$i|L�ËϢ@I�p�+D��E�ӹ+�t(B1���pc�Y	��'�,Y�	��l�Ԅ ��D�`̚��bM�Ġ$��Z�_ �MK��?�,���QaӞ|B0�ō[kΔj�
�X��ت��I�\�I-e��1�%�	�io6�����l&P��n�TUT�	�I©@����a�N2\�n]$�(�@E�R�E��OG!���V�Y�;K�Ս�1�Nda���\�t��Q�6� �ܫ�ēgi4��3��S�'p�!1��#����J\8q"OX ��:.qʠd�5-�p���'o�<ٔ/S&P	(��s�J7��k�o��@�07m�OR���O.U��� 3����O����O�نK�R(+��߼�+��מD!B����ɪ$�\ఠ
�2R^IP��9�+ed��)�'����3��IϺU��	K�#2ޘv�A�-�R��gj���\<0���a�� �H|R�����	�,�2���@�nu
2��~��I>1r��ן�>O�X����%�T}���ʚG4.I��"O& `�*8oa�DAE�D2/3��Q�>qu�i>!'����nM�0s��P7 �F���":cI��8aV2�?y��?���aL��O�D�O���JP6S��S�!��62������;#� 74p�XêNxx��B�i^=Q�k2l�%�A�DL�L�J]�#��9-�扸2�/q����n�q�B1�F[�\L�7  � d0�붉� 4t�����'�6�ަi��^y��'��O���Κ#��I�Dn�no�٥̛����	�E{�x�-ze D2f�ϝk�B�.�1&|P�O�x�঵�'�l	v�k�I�	ߦ�{R�Y����.C	 h�f�S�����Oʱ�V��O(��c>!�%(�O|O��eV
7�|lk��/@�T,��')�I��}R�ҥ9y��Z+U�si��k$�<��&V���O�LP�iU�u~��@���xhW�6D��s�# m'�0�M�<���8��Dک'!��')}��cP_�.���&��IA��Mc��?�.�Q�r�u���l��Lq�cM׭N��[�����	���M�Gޠ6�t���
� E�L����0zdx��O^��Qf
�(�*��2we�QxM<Q�$3e����h��s[l��]?aKzqh�|�PO�-U�y��RGFiV)�j��
����/�)�S-�l��U
T�+RL�a��	DW0C�I
:B����Gկ�r�b�-b���@`�'u,�9��!}�H�r�~�x�����ۦi��˟���4th�;�o�柼�I����P؛E����k1���yc.I�I��'p��.v�P��|&��!R����*b��1y��K����Ƀ�N�:8�Ԣ�c�;"&zc?e��E��y.Τ�������)�T�C%�|�g)�?�}&�x�t�Z��fD����&_��R��4D�@6�]##��҇�J�,��a�<}R�,��|�I<� T���	'$<^�sD�S�NnȻA���g�*�4L����	����	��u��'"�;��J�-2(!����T�
9bD�ЫK����õ$Ӯ���˨3�b�?1����y;b���CB�R(H;=LF)���[1 DV���Ĕ�j0��4\)����v�Ȉ���H�>��ÔAz�8Y���<���N�y�ټ����V��	��q�ȓ�ʱ`̀�%�e�r�
@t��=At�iA�'��\KA�~Ӗ��}�NaY��s��0"�\�7/���ڟ��	�G��	��ݟ �'5���P�I9`�z�z�m�9�Zq�Ć�K�n���ER�O��ad�H:Cllc�(
s3T�H1�'�������t��-�J����	 �A��1��zɌ���� ��N�i�$�3����9X��m^(9,m��>�����d �ɳ>�DSڴ�?�����i� ~B06-�L|�[�EͅvJ`DZ#�3
N"��I�PU�K�5���;����T>=�O�p	)�"R=��TȁOD"vNRhPJ<�b���D�x0ёaY6cT���D��9_1���K �8����B�I�(�uAg�x�Ɠ�?1�y��TDʛc8�C�
��� ��yB��24�JeӀE��x�nQ	���:�p<�b剎���	����I��]���i���'B#��d�H��'2�'$��h���ǋ�lҴҔ���T�����$0ay�BX�f���GH��Ib�"�@���'閐q�.X�D@+ &����5�U	xu��-�$U��L<�WDz���*7c�<Wv�0 � �ȓ3dBE!Yb �P[e�`�O�9Gz��tf��<��!ـț�c�İ��	ngX�)!+  r����O����O�%�;�?Q���BɁP	�,ҥH�
j�, ڄEԓ)ۖ�)�'N|��"N:�2Ar�U s�H�q���x����b޺с�JH>�ޠ����'�p�	��:��~㖱Tt�IC.Ԋ#����P!�y���>L ��)TA��'۸'U^b�iv�E�M{���M��OД-�Q��^����*���-���'zH� �'�<�2�0�'�'UNm���d��թ)�Q?�\��.��m�>ѡ�@8��8���)`(8Zv�IaX�4�q��O�T�OԌY���(�~�YGǃ����x�"O��q�Ü�J��XG[% m:��r
O
E���M3[�A�g��0c.H� 6��'�@�A@!{����O�'B���4z�\��@�I�P����_�H�����'P���2E�
Ma�|
��(u(B�ۜ%Q��3c}Z �&�xbC�)��4!q�7��	��'ˑjG����a�mA�ɀ��xB�Î�?Q�i:��r��0q��=zG�Lђ�J�X`��kD�$�OZ��D�;(bʔY���<wL�����s8�x��&ʓ�dY @l�>d�T�m%�����lvӞ���O��$
�~R�IW��OZ�d�O���z���Qm��XV@��DO��މ!�H���'� 93
�G�0���K�?t���1�#UZ��D�>q�[sX�82t��5^#t]�rȎ�{����A#����'�����S�g�I'Of��`�Eگ'#��{ӡV�_[�B�	�$���D�ywx�y�ꕔ �z�'#=����Y0e��C���&c[
^^ҁ�G�	��'w��'2��ƟD���|r��
]���T�R�<{�8�-��awt���~�0I"�CQ	v�2������L�)Bq��}<��>oq�E!�@R�u!��K��G�;����I��p?!O��0����C��8�@�iE)Lb�<���N�����M:+��Q&�a�y�O����ަ%�	⦱���U�r�ѻ��E-����+�?���%V�����?��O�raza��,��9˦�V1�X튓ၻZ�d[�D��fgP��m�3uџTIQ�.�D@��[��Hxp�͇%s��YFd �lh�ǐg��E���?AM<�V�Ŏ]�=&)I	~u�T�@�n�<	!��!���H!'ɜ�z*ゑg(<q��D�6j
�c5�B�,�1���s0���w�[�M3��?�+���:�lӂ|��hT2*A˓�Ǚb�Dps�"H՟��	5Ơ�Iw�S�,O@m��c_���Ц��$Hm�h;�xҩ
6�O����2�|��5�#b�]�(9��x��Ą�?�b�|���EC�Ȼ!�+�(%#r����y"l�f���� L$~چ��)�p<!��I[~�딄ķ-S$C�q�ԁ@��7��8h�Q>�I¦� F�p�-��+� `篍�-�hQ��>	�y��i�9X�)_��ኀm�H����[ "�lm�H�-�����yx�Ԫ�I^r<�bE�=s�<�e�;D����X	:m���5�ݕ r�4��g9D��)!�ZB�\�:'-G}�Ҁp'n7D�����N�DrZ��`L�~�x�k�*3D�X0��MR�!���6/�ط�4D�@�u��2:�x��N�(ѐ�	�o9D�`hGn�H�Hi�@L�WBb!o4D�Ƞ��i�hxʠA��$g,U��3D��i�aV�MOx��1�ڌ�ue*D�xp����
�� �*ߙe�h4���+D�Xہg	$l�@�&0W�N0��a$D�hCvA&��ђ�K�����7D�l4P
5��h�V,�s:6�q`�;D��y�i�(�X��*g�LM�!E3D� ���d[Ʊ�KρB�\	p��0D�ܸ��t+��Pd�J4L�v��g�0D���������aH�_�8��i.D�c�J�E�f�ORAe��5+D���%F�$�$�A�%G��bE�z�!��+�pe�	�f ,� �$ң"O!���2�I�`Ʀ+��xf� 
!�$��x����C�L�6(O�!�ҳe���Y�-����&w�I:�"O^0�B�!�#J�E���g"O�8K1�]�
���Rv!��m� Ы$"Ox��������`ȩ!s\8q�"O�����؎% ��N�)!�QX�"O��#�CL�}��\e�
f.2a���$Es���.:��&�$4z�m �F`���ȓW��cA )R��{�%֕Y��i�?�"�_~8��y4���Ksġ0�� eP|���)$�H�&���d�b��F�/b̱�Ѭě&�Յg�xr��ىifɂ�dȑf�Ʉȓ4f���dN�F��R�%�(�"O��"��ZVzX �	[Fd�"O��#ס�!2�0��V���KU��Ct�����4%��b�7��Y�u�S�f2�'�az�������O�c�f`R�+Z�g���	�lx��' y�	&��Ń���hr��`	�Q�\��N>�I�P�<��D��)_�Y0v%[:F�h#?���3�DL[iK�\����a� <�n�F�Xi1�"�)§3��@؀
	
����%A�
d�Pe��RL�<E�dcI��s!�=I6 Xh0HN0��'5.p0���p8�8ǌ�G�^�#�g��q��+��/}R"`��03d'�&Mf Ac��i�����+��p�D�'7���g�4!2U�E:�rA�E�W5��ɝ�&��>��A.~y��/�f���hv�t�'Rv�D��+��y?tU�p�-Hk�8A!�+�yB�<u�p9�ĤG&CA<X�PK[�~��Qd��h��A�ӥI=t9�a�٥|�TI�"OR�(t�ò"R�5jSƚ1р����>y�&,�ON)i'IG�^-,pX��p�F챰�'y*��Sߪܩr� �Fz�����.͆ȓl����ʄ�H����I*K�XG}"�N[�O��1 ��1�b� �A�"���'UTXh��O�~���H�*F���'|�Dy��I��vhH�H�.!��42��ۙ�!�DE��4`�v�A!@� ���ɋ��C����$Q
S^2��u-I�q�\@��H~��~��_�<��n#l�T���A�!V��IAN�n�<�G�_ ���ӈɷ@�9p@.Jk�'{�TD�dFV+|A�9�B _mL��!<�y
� �J�*V�O�$���4�|!�1�O`u
���2HHn�p��"�̂��^q$�C�I�_�������}�sE�.7�.O�u��W.8Y�- ?c��)@�@]�0�<����<1dM�<E�$H�F���$�  c�<Y0K�S��W�\� b��P�'.?�Za�h�x�J��U�_L�zw�(D��bjK# �-���~�8��#D��he���
�9�LM}�P�q'�*D��ꀻ}�� a���8�*H���5D�P�p�φ"Z�с���,,�F�K�f3D�t�����6�P�J�ʄ�26��H+D�0j�jV0.���0GJ�[���O'D�ԸDGW>:��I�i��~�<Z�.)D�@qr �� �L��qo�@�|:k#D�H�2l��q��(Ĕ1 P���y�I�5�h��4�w!���P���'܎l��MZ�v:r�Y���_�ܻ�'�H}�š�7$�gNI�Mg�m��'����%W/��")đ^��P��'�y����7CS^{��M�oJD%��'�R\
D��!%�� Z5^��E�
�'��Q� hF�+ ȭ9���,#�>p�
�'撱�7L�4R�iX���aB���'���΅"9F%q�-K�,i����'�d`P0� �b�ꨃ�`�$��r	�'?v��ab��]$����Ι����'����̟\ڸ��å�7rf���'�F��e��&?�uZs�_����'b}���2��Y���
�) 6�	�'U��ǅ�\'%��Dׅ[��ܪ�'M����9��`�fa^�P��U��'|��eK4k���&�@� �F���'��`��<=Ρ��Á�4|r)��'b!*P�	 	<�3ɕ1/��A�'��� �ʅ3��Š2� !��{�'ˆ���FL&���J�L�+�����'l$����7h0�P&$��-ᤤ�'�����D�����H�/G���'���V@��Cw�''��aA�'���G�@,�i�:�H�
�'���
Pe��ԕ�0� b��+�'���!����[����i=��I�'��e	!�@I�h!�W�O/U�]s�'RB��ee�3i��9*@�0�\�[�'VĒ�J�
TR��)��E���'�&Ĳ7E�2�`�Y�k4A�hX�'s�1A�n��^�h��V )�| c�'����qÎ?`��hhe5j�'ц�j�=��-B��Gp�I�	�' et#��v[�GʪX���'.�fAKv��qC��Xx�' �I��\� �ؽ��Ɵ7G�~���'�ZP�I�6&Z�Uh��<62�
�'�V"�7wx�q��$���Q
�'��y�gg[���`���,�lX
�'�:1�sN�&	�v�
@�٣7�����'F��Z��)=��0#�(1����
�'f���k�-n��P�(��5�NY
�'�M�5C�os,h0�A^5#(�=�	�'\����<v5>u��R=b�����'nz	[U-ς:��|!!H(\��m�
�'g<9BB��5Bt ���J:J�I��y��
�J�M���7q�Tx�VoԶ=1�0%�S&LC�)� :�u�B�^�`��%c��j����U"O�TcQ��3� ���ء&�i;S"O�H�CI��J̣���&<�R���"O	�u.�C�fl�3w��*� ;D� �'�R�=.t�K��ƠR~�0QD�;��7�R���T����j���IF�r 1I	�'�F�i��F-_�2���n&/܉K��D̃7n�"��ŭ��'A��$��-̔q""�CO(e��Fhx�%� ;�IK��:��p�Q[��� ��6�H8��Y�"~z����Nv	�%��7=D(�&AH_�<���^6��*K2�z��e�	���I��e�	T�F�r�np���N�~ռ�ۤ,\1�lp��]��}Rh��_��1�7�o�L�;%"�l�zP��W�|�ѦIĸ"QQ��Gz�f��yx�`JB'[�mR<TK�N��HOx�js�C�?I ���I�+�-,����$cYO����k���t���>�;��ab��H�;6��bj]-�%���&�X�󣚭2���r���"����'�����OV�͠��Pۂѣ�'����$$�J�:��T��/T����rۈM@ ��j�(K|���
�)�����-yA�5ɜ9��)Qf�Q�p>���0Eev	��ӵ
���D�ܣ&Q��BgŖ3)9jl���H1�5b��ɜ��9eC��a����6c6l�<q�Q��(Y��άg����f㗂��)�?x�j(:vo	�|9���	@�#����>� C�S׌��dn��:�0,�v�"]4�
�N��#l��k�z=����V8hӥ��!Ȋ]1�QY���ˁ"O�PC[����L����qgc�43 ���O5�ք��HϜr?��(ғP��Q�,ȓG%,uk�� 43�D��	���س�A��sL<�� �j	F�C�-U#	ր�I�A��\���� �{X��a6��MA~�kӆ=�v�Җ�!ʓm��Q���HJh�;C��>�p�ڮ�<=�!�[�~}���Um�8v�A�';R$�GL���`�Hs*+��5J�Ţ��A)��1m2����X"%9?��݃3��}��J�kh<t�E�)!�D\9:���ڲ��&SZ��a$�E��΅����,��y���BKHT �]?#=I�o�6���:~4�\i���lX�h��ě�Z��څ藢m�v�2�܎>����ᣏ.U�p1�F� �0?aP�Mt5Fp�unFN: i�HZs�'�Rà݌�p����G�A�S-t�Rɳ�I�� ;��#V�J�HΘC䉖3�B�A�Ij�j� ���{D��E}��6+F	`��w@4���y�k(�P��[�2\��"O�8�T�1(���P���2��:��+?���b,�U*;����7
��0�cO���ɀ���?�L7b�M��B�DH���0��-�&��xB�t����E#�*yV��ӢoI�yr� 3a2� !��z,�m`"%.�y��Xc��z���n��Ak����y���R|+`?q,�p�$D��yH4�2�pஂ�e-0��K�yr��*s�j�)t�E������)T!�d�"	�jJ4"@&_�U��㏜u!�$͏0�m���Z���P+ߡv@!��ÓvC$��UHҕxX�)+OA!�'t��ӦIV1b���෉��<7!�D�ej�1���s�L�+��� 6=!�@���a0��:۴���M�0w!���C34lR4g��p�&G�!�d�6-ܶ� �Ƀ.��5Pd
R !�Yv�yQ�*G�7ҖUz�j԰!�!���|2�3І��v5�k��ӳ�!�Sp^i��"Մ.�B$��%I�s!��8N�e\�2�ąђ
y!��!���2���>��FVx!�ă�W�4�6��O>��c�H6e0!�d	�(�c��J�q��h�':!��6C����f]� ̻D'B=�!�D�!.��]���4D��`�c��T!�� �x��AX3J
FU��� =��@"OV�re��"Y��h�l �O/�H�"Ot � �25���C�fn�*�"O����j��[�����"Opr��CFUf�0�%��H��"O�Pu�J00]:���(z�R��)H�RضXI��&$ B�ڧ�$<O�l�"G.4�Ah G�^���"O�|1��߯v��A�N��͞P�P"O�aʲ(ߔ=R�K��'M�؍��"O����B�)&[��@����T	�"O�����,�� B�(',�@�"O:yd+ݰN0(| ��#"s7"O�U�ek0eZ���?��d�"O�hzge�*������m����"OR��V�� F�؜�p�1�v ��"OrX d��*R�L�^�o�%"O�Q��!Ψ5Zx�C9L[Z��"O���LJ'?��!�P㜘e�)e"O�=yci�
*&y��"1�����"O�R��%�H�Z�A�2�8ū�"O�   �
0x6���`Uz�r!"O�z�(3��]���1W�@�*O���Ѩ�<6���+6솓sV�	�'"�\C����L�V��dK� 6Z��	�'���I�q�<�$,�%t"L!	�'��0jA�YY�8
7�6fsrP3�'�:��a�xvl�3V���Z�4X�'a|�X�O��qldM㵸�p���y�V74��S�ʃ �Pn�9�y"�� ��0����8tҲtXw��y��W#�����1s��!����'�yR�]�|�s�e�*pGG��y/�M�d� M^���3քư�y⬃�D3���
�PZ��R9�y������c�O�2T���;�y2�2^~��⅃3(���@[��yBiP�ր���� �x�;�JȘ�y�KB�N��R��Ww|8o�w8Rㄮo�,�zqϗ1p��r��	I�\����D�b�8��ҫb<���LͯX�L5S$!Ưy,�DzZwEx5+c/���Cm�	��)xw� \�I2��P-TQf���韨(zs�#H0��@���,�Ȑ�梘�1�L �Ԫ���?�G��B�֐#q�UK㾘B��e��B��ȡmQ�y�b�2F�Z � @�'����D�~2B�J \= A(��A�T �yF$ǫ|���۳A=*�!J��'�r����	�}��ӧ�)��G��A��EW= ��|"�K����'v�} �C��ZdNPs '�:�t��>�`��r�H�Bp 
�:�j��۴O�p�
�'�~lb��7�d�&�q,D�5�׆q���z7F!�Q��	�%1�,E�;�ě�@�E�8�Z���#'�YnZ�8���?E�4[����lŏT��R���Oܕ�5f �<�^$(P/ɪ_��Ik����HC"I�vEc��	7$�)�"�>1�#
�MN��H(?I�Oθ ��@Y6Q�p�#���,φIx��ڲI��y��]�r��3+K&�`�!�34�ʴ1�&ۓ!���S��L"t�@�zA$�C�ɶdigh��H"t�B�jA$�S�HI�e+�`�����(�b�S�u� M6`W�@x����j�mF8b����g�S��*x�R�1�kF�R�Lո扅8&��#<s<fE+��iݙ�u�+�����# ����ؔ=׼�.�<T�|�o �x�?�Os�YiT���B�&�6� �LZJ2Z�@/R���'��D�t��bl����^d��M����
́[���j�'(rʍaŪ�>�6,#,a��n-}�O�<@�Wf\�r.�����$�hZ��eC�0n��X)���8Ȓ���E��ExJ|��������� �Jdz�E_�@Jex�	U�Q.|A��c�a��OTIړdώ>�xAS��'�F)*�H�D�'�"}*��}I��1%<h�,8	�A��v�\(CR��:3��������P��Dy��6`\)AV7� �6MM�Y��P�RgʸFr�r��i^�����O3Q>���sRa*�tB���&�6��2WX�Р��mf�!�P�A��#�NQSw E;�La!�,	/�D�'�"�Dy�'ld�$�!˓�hƦ��C̞D��h��̈́v�
}�!��$����C�v��Mj#� lO� �A��@ "����n���e�6�D�l_f�쓡 �
(��}����{��A/-�⼻�MR2�y��ϣ��|aa��w� �b�"Q)W��=HT��7Vެs�"��?�`�*A	�y���&ypA
�s�İp�����5�O��;�a�&�y�ǃ��
�0PG�	&*bH�s��>`�L�'e��V��HiG� ?MDջ��ʙf[j�OD➴�'u���v�ɶ�X� g�5�$
`�9�R��4�
q�RgGP�@�֜�,O,�'��HM<���H!&�f�	%�~Z��^_~.�<�V�_�'�
0K3�<�z�ݹ7K�U���f4<�ڝ��̽��'m���T?q�`L�	�����5c�կ�HF�����h�У>1"�J�}��]�_��#��C�]p��(W�:7$�6�ې:�X�"}j���l1�#?u�$Y��m�	kT!C��	D�m3�+	5}$X��e�)O�T�|'�Kg��)M����92���j&4,�{�Ƽ?��r���s�	�f<8{w�NK���@�K�_���h�둓7��u���A��U���ʭ�����'����ߤOhH&Ş�Y�<���O��D�U3�x���3"2���	A4�0��^Tm$I��&�F�@cܓ9A����F�Y�F�
C�V�b���!�ccԼU2�d�hQ���@ q����I3�#ʖI�ڀ��Z���h)�O�>�^w���aWA�d��jW�:o�
�Ɉ�мLX��cSI�"[伭hS�/R�	�^���^���ħ� U@�刑X���+ 4��	�O�:	P�L�X	 ���fv-�p3W�̍e�zB�*�F�Ac��3���ZR��T/B�j�f*�?���?f0�3c$ȅW\�!*���;T��K/��AP��-7(�,���7�Gx�]�0��8Da_9{���Yq��13I�4
��'w|���뇃;�ء�A/�Hd�0t�z?~9����ߨO���I�)�yGJوlr�x�b���H� lP��xBBɨW� *��\>?ǘ�Q���(ڰ�p��D��8���T&��#L���G4-��	�T��x ��:~�y����N��?1F葤GkpI���:V:�a *c-��,����
?�J�p/���V 4Ĉd����-�N��O�h��ܓr)�<��@"mЪ}z5C� ��'�h�R�ËY�v���]�T�I{����,\�T�+	�p��3�a�g���aGE����,\Oj9��-�G����JV�`8���3n]"A{@�\a8���Tڼ+�(ٝ�L1b<6�\!�bkNV؞��'�b�䞧+O�	���!M�$#��X�gT�=Q��ڳ/Bl6퀆6Ԓ�b$ϯ�~�.�%�8��n^k��J�H���'�ʓ�(�s4M͜NV6-�1 n��ݴf^�DW��n0���v�Z�����p���-w��J���T��$�gG�_����v�̌$�qO�}��D~jik��M�dP���A�E7cUb(�'E�@��i؞tc�IĠ1�4�k��E;m��y�&�OD�F���p<9��X]6�ĜBi�4�e�(F��ŉ3�Ӆ{#�{bDL�x3:\�')��j&&�(7�t[��ӀG-��)���P�#;�����)Ē2H�TІ���-�5�� ���'�e�M\h�O��R�Ý9���jQ�о8x-���i�:ݛ<�)�)Vؑ�eK��@A2�h��-�\u�a��6��F��'�~���,U48J�!�<=I��W�=N�Q�'�P���	�� ��@ ������Z}�7�<d��
�5�����r��#i�z�	X�,�9"�T{�+!lO����Փ��� Ͱ�Z�-��A�䕛0h�0�ў��6Vl+�y��h@9e&X-���)t�vGl�e��;+�eS�d"��jyr�96�l�a��({��dQ�l���M��q�
YSE$e�h\q%���S���"�RB��5�> ��<��{�/Y�	�6�˅ ݣ�5KƯƖ���LDh4�ԤI>��dɓ$��#�������{����U�&�j�$�O�l���*�M[��D��tXAàR�%/晪&�̔E�HUZuC7�F,{5�d��ya��US��GW�$���*>��{e�pѣ��!n�r�d��y�6�	7�	�0s��>u�py�K [��ɑ�Q�ع�ʌ� K���`��[^@5sf�+O|Z6��@3L��� 2���=�ڔ���մP��҅	\�c�M	j\L�MO��1��E;6����� ��I앑%M�_�tI�F"?)'C�?"���$d@��&��]�'��-cD��,�����4`1�!�&�qO�3��~�*�;]t6�s�)��@�>��(Ζ!���Ao�G2�G~��@����<q��1��5}���t'̨s^6-^>���"}����jt�V�JA���+_�K����剝1ju�R�Z0����#O�N�˓�P��̀-&Ű�@\�I����'���j5�$�V�eˑ�^T�1˄#Jt4�Cb�E J_P�ȯZ�<��@G�d�^��m� `���Aœ�L�qO��O�����գR�^�!�H֤O|@��󗟼G���	��(#�RRx�xP�+�S�? �ԉ$��1k�x�b�EwD���\�2�➈S�g�S�4�ο`�̹�f�Ю;�Ȉ�F#�*as��	�Ì�-f
츏���/����w*�����%V��̨C��X�Ѝr�4U��q��OP�7
u����*�u�%0:�dYᤠo�����
���(O@)k�-z%dX㠨1/����R����R0_G�@��	"_M���ю�>9��$߸'A|�2>�53U��S�@��j٢0͠�'A^��2�J�	=.�,�ڀ>��Q�'���Ox'�,�@�<|f�;ѧ޲C�l�Z�3?1rZ����a�&*f��17�I7+r�B4�F'�8��	Ĳ�<�$7�Ig8��(�MFWb�!JG��,d[̈����"Yd�r!.	�4���@����	��y�	�^�.%�4�<�@�d$I����#�ONt�3��+B��ɠƽn��jF���M����o�7D�4{�}򊛨��`�Ejؤ s��0�酸��=	6O�-c^�I����O�)�����u��x5�[V�t`1d���J�X(X�Ē�0�>b�(Y�����O�5�%��6`,�ۄ��>l+Z��T�dU+v�ivC؇}��Y�}�j��4��i�G)d���2]�i��'>$��A/�(T���g̓#��Q���vL<[�\�Ʃ��-4�S���<6�<ۨ]������TL%+X����
�Iv�c4�@�M q��ɚ�].�Y��D��e?�1M�N�'�0��}��W�LWJ����Z�^�|� g(B�g:�,)v�ԩ�~�'+gY E	kĳgf6�A���
���1SV?1��Z������J����5 C�P1�\(�%$Il!���0\��c�إR��A�"��o�^ ��M}��E> |��(�)Υr-�x�Ef�.&�8��I�y��'@8��Y�9[�](�J�����>�j	<��t���ٰW�����!iV��S��K��Ƙ\=n�z8Oz��b�7�ıC/=93 ��M�L��tk]<{t�Б7�@�Q���]��rgE=9��j��e��*��?_��Б��v���,E���'�Ե����xYe��7 uv��3OQ�Dv�L��ɱi\"E��j���k��,Il�'��3�aޏEm�4��E_=~��'X�,h�I\����MO4}�~��#��c������օ`T�X�Ϩ w��۲^�PBd�Z<\c�b�c�
Lu|��q)5dV(��7ҟ�`�Ie�\�C�M��C@4a��ꚿ)�7���1�(�w �lX\�3MI�~J��DZFO�1���bM�cu��G�4�}�'7�8�����̟��><�Б����W��(҃�O���W�P�n��Ix�b�}��Ÿ��i��%��t�����UУ� �4� U��|Bj�Q�BQ;]
�➨{���N��u���~,&q��d�`szػ�&���'wT����M3`=�M�b��&(f��qG]8KN^4�F�2z1B �0����*���1B�t�?�'X_
]P��J�/���U��%z�Ib���Pu���WC�j�jXa�K��@S+,�����V��H`�������bFÚ(K�V��C��) ����QG7���	`u���UOG&����``ſ��'��)�4�ҹx%XB,\U�y� ��M󨝊U��1d�B�qR)��?#<�$�I?&�2sE
WZJ\ю�z}t�b�k�	s�Ԡr���Qm8"=��E4z�Q���s&�x�����#Cv�#w陦bK��	qϖx�z�Ey����c�v�!sቆ"˼�uǆ���E/�i�\i��
�j�|x�A�d�'�>H�C#�=	6]j�����'A8��q���(7q敨h�1;� �'���)]0�1bj6 p����әG�<Mqu%��3(q�I��:n�C䉔N���P.F�z_Й۰C�'vE�B�22�����ǂvk�`R�ȳ��B�ɰ� ��eE��1��Uʚ wb�B�I%i�h%�!ζ2w�!�'�Xz52C�I/2+p
�P&�Q�֩� #�LB�	�B]e����)��#ʈa�vC�Ʌr�P�3��Ө�r�R(�B�&xڴP����u�F��.�G�BC䉗T��iP�+�a���y�'7Jd�C�ɼ,J��NV;n˾}�vN� 	�C��+(��5�������ҪC��|C�	�v|	��/޸Y�����J�?!4DC䉮jt<���DFJxjݨ��Q)BL&C��,%�z������#Pk�.��B��7UOH1s	� ʴY��	�+-�C�I)u7�-)��(vB4�!��*V2C䉷N�>��f _gU�p��.݉wV>B�I�F_/Y�6�Y��ʝ�	K�"O"��A 0R�6��U���D��"O�c�#�9��	��?���D"O�Ѳ!�_/xA`��`KP�x�q��"O^�3	�t�tp� ��6��h�U"OB
�/À\��ܠ�,
'm2��"O� ��x������dk��b���"O�A+��%o1^X��g�0y��d�`"Oʤ�P&��#1FG�G�) "O �$�W�#4���Z��:d��"O�P)�L��j�40�Pa��Y�,��"ODA{"M��\��U�b₴/�L$�"O�`�u�ذXFF|cC,�+YЌa"O�tȸ+�,N3D�(�31�G-�!��I/:��:�!��w��SR
'�!�5Z@��$�3v�l� �F�!�DژFN��94%P�*>\Q��x!� �-�ȡp6`��6#̜�u�W�!�$E�ycܨv�Ѿ �:�{b�6�!�d�;*�hP�,���hh�!p�!�DY'#�\��ӡ�͑vGԔz�vC�ɧ^�r1���BDYz��ש�>�jC䉯d��㯂�i�X��G�}f6C�I�.���m=<��y�-ڙ
V�B�	+�aI �\�|�	�P(F�C�C��_��D�v�zx��tiG��B�	�>� �c%Y��#���߾B�$(thAr�#�"@ᥣY7�B�	�}����攪"$���ӑ[�jB�A����H-F�Y��0�8B�	�)�f��&�0w���K�OL]bB䉦C~�E�C&��w��Y����DC�ɹO�3��L;i߬Y&*�hPC�+W
�Иe 3_~ q7IΗ8O8C�	A����'gO-Q�l�sĈџb1C�I4a����R�a�D0���(C�I�M�	;�h/k0\V	���FC��)� ,�U"�_�^$����+�C�I:\��@Bʌ-'��8��� i�C�	�#t(���<.jA�S��uB�C�(����ֵtd:��F��g*hB�	�$�2�EKBA�lU�ѯ�
��C�I�o���� M,@�T��9fTC�� \�BDr5∌H�Ը��i��5�C��d�0�T�΂-�����" ��B�ɯ<�� a�	]��D�u$T�d`�B��#�:���H�^<@ł� �ZC�I�L�hJFㄤw� �����6C�	�vq�y�Ӏ�"?j��wK_΂�-D�p;���3���j��ŐY�x�S�N!D�`�@^9Y�H,�C�I�k�x�vH;D��Z��=�5 �GC�`���%D���	�@K,���QD�hY�g(D�����Ħz�n����Ah%�@"�O'D�X[��՘H{�Κu��YE#'D�̂�4v'|<z�(Wb bU�Pi/D�k�
ͱ:�v���,ҫJ�|���.D���"l�b�Ju�O�F�xRF*D�(	�D_�L���%@9�ɒ%f;D�4QL�-�z����ϩi�~�3b8D�T �U\��ĠHK� ���5�7D��X��H3?yz8�4�J/3C��Tm6D��FM�`2�d�R!I�\���zDh(D���Ȝ	k�6�#���p������%D�	��^� �p	��D��T����#D���bͅ]�U�Λ�e�h��<D����m�	+�ኦ�[�P��.D�\#�
�<2V�G�Ĵ��y°�.D����G�L���t��;���3�-D�$���\a����8D��[Ak*D�� t���V��Xf��$�⸡�"O�1	�ĤKb����͗�}�z���"ORI �Է{�xb��?�V�U"ON���$:L�x�Ÿ[K]��"O�t�B��u�,�w)X?o3~� "O>q���ɷn�S��;c��q*'"O�	sE�	-�Xqg��/�(#g"O��&�M&P����(��z5�"O�!��1h�YBHؙ}c"�@F"O�Y�S/;BgJ��E&(IJ��p�"O�X�!ʒ�[���s��v����"O )R�'�*�j� T(<=1�1"OLxZ�����¯ר@�RJ�"O�պB�՗Q�5P��4�6�c"O�ui����R��A��}K�m� "O�m���Yw���B̈=ȼQ!"O�pS@�9\P�A�e:�Q�"O�hY�(�[����􈗄w�L	s"O$,��k�:e�h�$IПryh���"O��[T��,vw�9�AŃ�w2�Z�"OHE�����,�Q�D� &p�X�"O.�U��/)xT2�̀%,m��r�"O��2t"Ҝ;i�ҍ	c�t�"O��+��1;�D������C�p�q�"O�]��k��=��鲲j�m���IF"Op��w�O�r��<p�OO$����4"O\<*vCعW퐑�󮑫#��1�d"O©��-ƎxJ&EK�h�<��aG"O�x�OD;.���wHH�nj�(�V"Or����`ݒ���W|�!(F"O��8�ǌ���5ZPiܔ^�ܘ"O^���b�*�f-B��>sV|@r6"O����kQ�P����S�5E2,�s"O��1V+��B���K�L9d@�h�"Ov��w��:+E�p�d���a�PH�"O���eK�>�=����|�*�`�"O�1&L��pT�ٓ��\%:���"O�@3�o+�T=�G%M(.i�=�Q"O��`g�"�X�Q�ؐb^�5A"O��$ǒk�R8i6eݬ EF�3�"OxD���3rb��ʩ@f�x�"OZ-*�֠��S����%�R�x�"O�X�ǀؤ)�~�8�&�n5h!"O@��Nպ7(̐f�\��8�"O�@z�L�|����f���!���5"O<Tq����(B����)��i�"O�����K��)����4P,ja"O2�0��-��-"��%�@��"O����@����ώ�e�P�;�"Oh�:r+�=���tn�;B׶��"O.�+ ���k� I� .��zɜdBv"O����F+.9 �!�L8;&���@"O��pF��2�v��9p�p0"O��aF��+�$E
�'�2,u$dx�"Oq�1 "�&����_W_@��"ONX�"-ϼU��)ba,D�r���"O�A(5h��%��쨰ς7��mɣ"O����A��+����m�v{��"Od,8���3�|�j���7}Ԭ%��"Ox�*N�>�����
�8�0 "O4�[�Ӑ0,�q�Q�X)U�uBt"O9���v�r�k	�:2���+�"OmiP���!Aɇ�(�x�iu"O��b�S�q�6劲-]�V�X$"O� �pp�$Y�5!t������"�"O�]b� [u:@S!A��dfn5q�"O.HzA��D�L�j��J=NS>��"O^�@��d��0�W�M0��"O��P%OV�(O���i�`=�(�!"Odx0�
P3z�ԪpI�)�U��"O�	!�F� ��T��.d��Q"O�����=���(Y�Z���"OH��Z�g��U��3:�.(0B"O^-�aˏ�6��,"%ͪ'��x*"O� f'L�'8y�BE5M�>]�"O������	�3Xg����"Or!��A̟3��Q8Q�\W0PKC"O:���!ފ����R LU�i�e"O�jVJ�b��}��֜S���Kb"O��Q�@q'r�k�L#H�^ѹA"O����ς-�L)B��0B����"O�@5���9�D�v� R�:�!�"O� ÷HַfA���G��N�ڤR�"O���I0|�A �pfP�6"O��𫔬_�j-i�̈́�nfJ���"O0��� .���q�M43VZ��d"O�L8�Y&,�����lF��P�"O4��!�����+c�,<+6,{�"O���A�"�`x���^E4h"Ob�C0���q��9�Ε�B�ኂ"OlE�vWd�Q�0�B) ����"O�y9��T�u���9���Z�MP�"O�m�q����@��l�\e�t"O��c��0��	��$P�N�s "OȠ�cD�:f
��5&4;�
��u�|��)��(����pL���~s�o�M��C�I
l��oO12*6��b�˙H��c�$��	,�ݨ�	D*'��<b�*���B�ɓJ�nP��A�}a���g��36��C�	�Z:�i��Q}�.��@�,�
C�ɽADUHң0�e�bB��YsC�ɨS��A���6e)�L�UdXh�$B�	�">ƙ{6��:�Y����Q{B�I�JlY��&�
.0mh�M:}8B�3g|p ZdJ��0#�$9�B�I,G��̒"[��$BG��Q�B�6%ز�!�Ö�7[lH���L(�C�	���Mk��j�:P@2F�7A��C䉿k�%�K��O�ܼr� ��f��C�	�O@�p� S��$�b�R���C�	Ƙ19acהYh���e�..�B��0~�H��:S��S�E-i�B�	 nX�!#��ʋ7H��Q6(S�B�	��l-�2���Vp���e·��B�	-�bуtIZ�CJ�m(��X�\�PB�I�|��e����W0���0#\!_tC�I�z#\��E�J�b!�1i۠�~B�ɲ(��ѩ%��$I�s_*K*C�ɬd���5)C�{��A%P��B�64.��c��-��ŸH�(
B�I
d5d��v��-w<���p��o�*B�	"b14hD��;G<4[�FG��B�	
{B6A�`�b�3H$eB�	<Hy>	�� ?T�#6�B(O�C�1xrI�!ٹj,E� �]̐C�	L��0hR�#tLԊ��z^C�IEv�
�5 �2�P:�,C�	VoX|�vA�0@��GlQ�C-�B�)� NM����)kV������rh�z�"O@�"���l�ri�͋'�D,I&"O�pjޜP��qa펎-���(�"O*�JE,G3�!����^��(Q�"O��3s�?	�20�Sl�8����e"O\:g�d8ܘH�K;Z�¹�"O�Y��H�,9���ф�^��� �"Ov5�'j�P�蜀�ڠ���"O^=x��'%2�ʱ!��"�p"O�!�lE�8�:�Ԧلip"O�%1!�$qw�R�l��5u�yT"O�B����&�WkH�I3"O4���֥{�f`e �j�E"O$�Z`��4�|	��-�{�0�:4"O�����c��[U�ɑ	C���"O��Y��j��0ëޏU#�x�e"O�Jå�,�Nĩ�ۨ-�ȑ�"O*h���X-2̬��G�+-A��"O����K��C*��f�;B�#"O�%�d·�\��y�dŖE��<�P"O��W��12&Zd3���bB�%s"O6�b��T2F�D�bRSK|5��"O��q�$��ɂ���C/4�"OH� T�Y�{�qI�G�t(8�"O�K�GS�Y���Xb	P��[�"O)C�HW�$���c�G�P	
 Sw"O����L�z���[Ѧ̿S��铷"Ot���z"�]3��jB��d"O[����$%�F�/x 䐷"O�-�K�Tx�%CG�(�pa"O����Aϫx9X (ǨO����"O�y;�c��(�8��e�׌c�֨��"O4ҢȞ0�fHbJK��"ᘗ"O��ڧ|�J���*�\���"O����� <CU��)S�L겜8�"O�A(G�u ��Bvi��U/���"OV����H̄<c��P�OF$I�"O���K�ֲ�)e�P-Y(��`"O��bn�Z��8�#��6����"O�|��Ï2���u������a"O�A��,�<����%��z�"OM��C*f�Z����:'
|ڱ"O2�)'-+J�d�5+]�n3h9h0"O�ͩ��
#����g��H��"O�*)T�]��T���J m�(DqS"O���3c���<���T��pIy�"O�UGG�B}$��)�� �^!�"O���#
�B��=���5~ ��r"O�	��$y_tq�����[#"O�X� �2��9�&B���PYA"O�Hh���tup��S�?'�	x@��ߦ�F���!FH	�Ɇ�EFQQM��y��!P}���!B�b��P�y��ID}��##n		Bd=1bjĺ�y�E�4���4H�g���k������>�O���� P�J(�,O�"Jr��':��8T2h8g��R���rei�w&�F{��' ]�%H"��
C>5��X��'�����eղe"Z�1qi("x pc�'��(�Ǟ<i^�x aς$Y�1K>a���	Ɖj�l��C�1{#r�N�k�!��.o�h�B`K�i	�h���E,<!�d��P�HB�.�1i��'� '!���R9�,���BN�l"��ֈe
�I��HO>� �G@������I�x}�uV�H�<a���J�r�R`X&/_�?Ō$Sa&��(�����	�U�ʕ0b���V�� k��J��'A@�u ��:6�"e������a�'�|��o��������g��5��',I��l
� w`s��O)�\����?�_�"�b��K�ZpZ0^B\��i"�@'�*1$�M�Яd)�!�	U����t�pvNE�xc��vяK��P�L%D��eGyvv=��fЁi-�� @K&\Oc��X�F/:�0����%F$�"D� 1"�;Xh&`KWgϨ�6(�B, D�� C�	���S�B's�
��?D���.α}� ��5��:D����>D�L�f�*up �C��j��j&&?D���E���J�L�0"
Dbr �{fn3ړ�0<�ul3"Q>�#�Vx���eEX�<�@�դ������P!�������X���W2��Cɰ��������+�x���`��xz��_"q3`qI�h��1|؉����?���Q�=\ܩ@jc ��)���^�<I����9҈��k�eQ1�Y�'_�?
c�D�j�0�	���%?fm�"�+D�8���E,jgm
�]T�r �<�����2 ��$B��
Sր[�$�2cd7�(�r�K�4f� ��@`̉m	�5��hO�'u�]*d��2Ξ�'��=��B�	�H�ܒ�A82��<Y���QضB�I�s��E#W�ѽ-�����\R��B�I"nY�a �ݙu�X�0�F�"�"O�Y���;A֚xaSiW.!pe��"O�-Q�DY3 ?�U�#hN�S�:��"O���b�sN���|G.�iu��f��F{�Oz,Aiå�~�����\�
�'��� ���Z� ,�e��t��$*$��e(<9�i�J&�*fdٞXd���]�%�t�<%>M�����q遄&J�g�2�BG2D���#��+-6�d���S��*�!/D���V��-��񚀍%]�zC�	��q���6hڀ�/�
��C��;F0��f�ݫ���� �$io:C��p��t�Y-7���)uX�4�*C�IlP��hs�ă)�$�b�V(eC�L9^���` `������9
C��(42��,&K��[5AU Wo��')a}�N��w�bl�A�C7q�������yB��k���F�.p�8�I�O�5�y� E5�`�
�a@l��p���yB��:�صbׂCR�41 D�y�FI
�ah$C0Q���Aȶ�y2��L�� MћH�)�#�<�y�o�.6��XB���/��|A&a���y�-'�.Dk�b���ź���p?��O�d2��!�4]�aƌwU�I�"O�%�"��Q�v	2��_�;8���"O,,a��+�.5Q#�S}E����|R�i����<�㎣e�He�E�?}=�y�+�R�'Tў�3�Z�c�ñp$.��%!ݲP�BԄ�&N����ԓ�D��vON�P��Q�H<��O�Y_�'&
��vÑ�l�h]i��Z�x[vN�B�<�wbX�7�6�[bcmU����P|~�Q���Ic�����O}���%`L���=6�ɛ	͑�l���OԦ��'I �BL����a±��u�N�LD{�������દ�}:��0� ��MÏ��s�� �h��A��<6���a�p��T"O���DN�%	�.}�1�] C"�%����u�$>.=<`&7�bӃK;>��<��Ik}�a��VVغ��B�a�^�����<�yZ���pGM���r8A�?n��؆�W"��iC�E��x�����a&�ȓn�*��J�63g�H��
;�m�r�����vo��J����DĢy�4�BFΒ�?!N<1ד��)�Bf��庐����Ac���'Ia~�b�Qw��	�Ƃ�:@<���^�yb���B�^�U�����)B%pi�pZ��D$,O��Q�ȓ����Zph�*"�퓐"O,���IG�WK�8�"G��7~ ���"O����N���R�oˇ5Bn-i�"O0�ZTG�WAb+��Ԗs7�%c "O��A�T� h[�+L2DF��0"Op)"�f�~�(п�]�BH,���r]K�Y�b9RBL�44 �ȓ\y`y��{�laPf��`p��L� @�x�[ge�T4A��)D����~,pCAEZ8_�`%��-|Ӷ�=E��4d�� sꑔR��C䧆�^��ȓR��U"I��g�2��f�H�A����Pn�T�b�E1r��t�䦅6����'��}bA.b�y#u��+چ�
#�
��H���O�R`R�mN-	�^Djr)TSn�����D/�S�h
3a���B畨�4�P�!�hO���IV�v��h�@���<7:�Am]*@�!��56�~�Rsmɴa��� !,�#oy!�{^T,kS/�a�-h3�йm��zr��@+*0��E*s���%K�(�!�dΠR1  ̇�?d� ��(���铢�>i���$FK"EA�c�7J���)�V�<����^�����Y�+MD��c�VS�<)Gd׼@Blk�-�af�$�eKV�<�ぅ_�
q�_� p�̐��TN�<��m̺�"��^���u-D<���Wˎq�3�ǈkl#EK�N&R�ȓ Ϩ��T��p�|j��ֈG7|ه�|�|�X��Dr �������Їȓ>�
8Ae��BEb�cV#g"T��&�fH�Q�X� ��G"�h[����@���@�ق���iP�
�Ȅȓ$(��͚�i�x@$C"fe��]j�Pqȟ����H����0�ȓ����돁:dؓ�iU�/�Ԙ�ȓh���0M�=,� ��Z�$�ȓ�ɩ��B7�nY�Hݤp����ȓl��S҈Ǣ�"�@e�"@l��ȓ_�,t{S���DA�� #@#��i��o�j�󦫋�]
��S��/"���ȓL3��h J��UVuK�d�	'^̅ȓhR~�8%���| J���嘞L�Bx��M��|�C�K-{pr5�D��D��y��I7P�
At����Q6��!�ȓ1��q��
�6�8�B�A~RU�ȓ&|N����
i��	��u�8@�ȓR���� &|�� �ʃ]�p�ȓg^|��5B�sk���ƅ��$�ȓ
b����W*Zv9���Ɂ�6��ȓ�+dM�|�X���?r�M��br �c�+L�,�P5a�;w!�}�ȓ]�2�Q0���-!~̛���o1�D�ȓE� �����+M�a;s�2+�ę��S�? h����:�:�S���>���E"Ot�"��?x�a�X�P�,��2"O.\1E��I����������"O̱S�B���͹��9�쥡�"O\hᥡq���l��~��7"O�Q�j�9^��iaE ]�>ٓ�"O�}��Ȟ�>���Qt퉻&�(a�5"Oh��d~�(X��,�I�"Ov䚕ʒ�O���a�L۸p�D�Ȗ"O^��ӉC�&A����8�����"OJ�0��P:+@T�B�I08�<hx4"Or��p���'�.�1e	�
]>���"O��'.�/xG���Ȟ����	W"O�0h���o��\��f6Xk��`"O>HY����U��$�6 K�XK�P��"Oxt�O�= ��%;��/M����"OB]�u�F��xB2 [0h`��G"O�A91f��{��T���yk���"OuC��D�Lq"��q�J�whD��"Oι��Oɍ��\�"�8t��x��"O�P��H�
�j�b'�����"O�q���.`nI
��ÅK����p"O����3d� ��,��F���"OV z�O��;��y ��F�$L#�"O��AB!�5�r�#���T�1��"OEz�' ���x��>��*�"O���Z"Wg�+�JI�l��`�"O�}!��~��a"�OI'.f�"O�X6`�^��	�.�;ld����"OX�2���#u�*SmևdQr� �"O�y`����4]`�F-qBf�;�"O���a'��K.0ȷ�?1���"O8��V��P�(�eO�$��"O>ȓQ�^����0��7�ʴ"�"O��ģW�Y����l֓x��"O!�S��3W#��a6�ݏfjdػ1"O��⅁ٛ-��M��)ڨ����R"O4��u�7X^Mx&��[��l�A"ODH�w/�%|��X����\�2�""OP1E� ��ny�I$.Hн�u"OT R�	@�6:���c�-A�-8D��2F�F�)�is`�M�ypӥ7D��0vcʒz�i5�הH,va�r
6D��j�K�\4�c�Ea$q�k(D���1̂{ϊY8��Q:fm�TQ(D�8����4Wݔ�i���L=4��#1D� ��o4n�����ҚOT���
#D� a��ߔD�v���lQ!CeLq�f,%D�誗�C�oc��.Td>R]2��5D� �%�Ûe������uS�4D�T#O�L4��[�-L�M��zf�0D��!�
6#pH�b�ʼgx�-D�d�6��$FZ�X�킜:4�a"�?D����'���l�yD�@v^<��>D����� j0��w���rA8D��b��S?P�d�@D H2���a(8D�p9��T�r'����a޾:KJ3][!�d��Mp�3���8�ZU*s�JRP!�D�8�H��$/j[N�Ȑ�=*!�	���]�d��0���#u�E,zC!�B�6`�P� ��k��H8�AN�-5!�b��a��R���+��٧ �"]��'7�x�As����_�o���'��]��� �|��u��eY8�R��� ����kW�vs4���)G�=ņ$�C"Ov��0�
�x�[��7hî��Q"Oҭ�g�M��d��G��j�X�R"O8��3�\�/}DX�A$��&6ع "O a��J"2 �@��Me��Yc "Oĭr�.Y5�$�fD�M�Q"O�G��3Br�:�$Ͳr{����"O�i�0��;4�ŀB�?t[Uc"O�m�4g��kR�yР�=C�Q�G"O��R���,|�c/J�d)��B"O�-xgi,u�RKC/S!.���"O�\����Q���햷!����"O��2D�JI�|�Z �Au����"O8i��>V���T�A���C"OΉ2\�$"=�g�Ⱦ4x��4"O�d��I��*��ZUw� ��"O>Y���Ys�$�.� $\�[#"OP�*��S.�!0����s�"OB�s�
T?�ͱS����F"O>h�L�<��� ژH��a&"Od�+�͇�	�@œO�|O��p3"O����9���`4$T�#O��"�"O�Q���O�D+~�Qsh����"O��	v�ʲS2 k��*A�Ju�"O@D��h�u��m��O#] �a\C�IF `[��ՙ;2����ܿ B�I�)/6��f�+�����&�Q�C䉞kL<�2��Y\�����B�|�<B�	 ^�K�j۷��Z��5/o B�	-�� s�A�q�����s!�C�	�
��E�BP�����=v�B�I$�bV�˯,��ې��x��C�	r�\S���X����7��C�I�4��@��űf���oݔ��B�	�%:���QR�x���,k�jB�	23�&q���W.5��g{I�B�I�?�]�c&O*�:�+�M��/vB�	?�����߾
�&�����>*
C�C&��A5醟~S2{` �"B䉣fY���&3:�
#�XE�B�	(��AVN�h�U�bjlB�	5;v�Q���
�>�so�$U B�	�}e��F��=����!S�lڐC�ɝS��<I��#0�8��ѷw�xC��?a΄�*��[7Uݔ$��.�+B��B�	�4�D����=Bzj�*W�1T�B䉶k���@;"Y���3��Gl�B�N�|��vЄ{sAS&�B
2��B�!���j $B�{��A40ZB�*W��[a,H� O�5R����"OH]�Qh�,���RM�2�Tec�"O��#�J`�5�ƫ	�v�
��"O`���o�&4�E+'���k��Ѐ1"O���@��!��Ap��Ϊ�hIW"O�@D�
)������' R��A"O>�j�IH�Q2�!9E C|e� "OV�bv��4I�.=趌!��]�O !��9���������ʅf��'�!�dD = l�Ӎ��?F�xe.g!��_�ͪ��r9\%:��d[P!�d֋_X𘂤	��Y.�s��,4!�d�"[����#däL�<�tN�'!��\!Z�ꍰFdǞ(�pj�N��o!�dI�Z��:Ԍɢ�t� 0���W�!�� 6�������G6T��bu"O�Uq�#�&e����[�4�B)yT"O���'@�$���X�֢!��xK!"O��N˩P�M��Y�>�X��V"O�ꄢZ�/����#!QJ`�t"O\H:"� $k�6m�2cI����"O����s2.0A��"3��w"O����';��̉���c��(e"O����-�n[����σT댵H�"O��1`n�89���a�T��"O�Ĳ���*"V�����4F�Ѕ�4"O���5��{V�4f�81�ĳ#"Od� ��W("�I#�\�,-
�8�"O��Al &Y��5�i��	{p	�"O0�r�B[�(����ը��8g�	�e"O8�B f�l\K�=b����G2�y�%���A�GA<�b(@�-���yª^"v���!i�#�H��ъX�y2��l�X����,7>B cI��y"�9T6d��M��V�Z�P�@��y�!��s�9�-��}�~U��h^��y��c�˶엾x��5��F���PyB����1�d�Ϻ^T�0i�W�<I�4/��iђ P�@"0ńQ�<�c@Y�v�DlJ�C��B�&�z�/LL�<)'��
?�zJ6��b�<��g���(�t�B7cXFuQ�Ib�<9s�!Cq��լY5C��)ASȀZ�<٧��i��-[CB�֨+��NY�<	4�ۋ$
Iz�nH�0؃�F�S�<�Ө�'��}qB�,��BJ�<1�C"?�J����9Ƞ�
A��_�<��ZE;�*�`��L��X�<ه�'�R�S���H� b�}�<�&*˧T���1���
���Da�<��e>*c�4*�n�6���bXq�<!@ևi��H#14F���rU-H�<�g�ԶR�� �-C3Z眙�c�}�<�uI��.Z%QA����u�Az�<Ѡ)�~!�TB`@�:h��	T�r�<�È��/�0��ȳu���&�Yr�<ك N� S�\,���:cBp�<)G�,J�� �Q$U�(@G�<�A��2>�,D��U�')�h�D*�J�<��$ڱeò �Q.Ӭ�E�d�k�<	`ɯ1��p�M�"aez���F�l�<�K�E�,4��ጩ4s�;զXR�<��䏨?bm�w��'pR�T�t�<Q�#�k` 4��n�h��ɚ�JFm�<i*F>N#>uY��SEN̫aE�S�<�7!��#1��b�D�1�R@�U�<��q��#��Ն9	RE:�kz�<�u��I>���
9�eh�v�<��DL�f�nM��.#�rA�2+j�<���J�zV��k͐n�8���q�<�L��Y8����_&Z�t-[q�<���3~�����Ƀ{kX�����B�<��
�bd�)Ca1S�Q�g��}�<��J�5sX9�q��7+bT*7M�z�<�ԃκ���*Rd��j
*���\�<1âi���'e��q��0c|�<ih�,I�h�E�R�r��`�Uu�<ѓf�8| �����^��aFON}�<QWj�c������)J�,�)�d�<� ��C#�¾ �T8ǂ.tt0��"OĬI����.�:Ƭś"�zd�w"O�pc�Z�	� ���H�2U���R"O�d���}��wʚ=M���"O$��w/Ц5tuR��P��xi�"O] ���(|�f1!7L��� "O�����<x�8���Rn���"O���%i�|UrA�7A�.�S�"O���(�AɪX��Ѷ_ډ�&"O$����2���8`���"O4	a��E�a��X�(�"O0<2�O?$J��
Oٖ�:9q�"O~1!eŮr��<@p�ĕjpv��"O��P�Ǭy�
%�E��!)X�rG"Or��S�a���9Q��6��1"OF$+fY���d� MN��y� "O��P��Ʒ\� 0:���<N�bIh"O���"�!��T�6�S���B"Oj���K3\�9KP���k�5z�"O�IK4,]�%6�A@O��!YQ"O�i &(�=�E��.�6In�qC�"O
!�A#� \YQ.�?X���pu"Ox���
$��I�¬�k"�]x�"O��4
Ѝp�a�`�1��A�"O�x�.Ӯsm&=۰��պ��"OP�b�mU�~7���,k�A��"O���XwmR�r��E�j�Qg"OT��`��g� �S(B�t)�"O�4� F!D��ě��ɓbR4�'"O����ٳ[�����˪Ee����"O���ȸ1��`2�!�SPdQ�"Ov�Ǆ�R'4Xz�`��u5�1�"OhI �2�%���{���"Ou`�b���Q��!Ԭ��,�Q"O�%I3�54.�0���
��$�U"OΖ�Ae���2	ǡ]��D�Z�yb��,K֌��-�������A_��y�f+\���G��R��t��y2%^������N:�1"d�9�y�JY��슐É�dĂ8BR
�y"��y<%��h�N���r�]��y��Z'sh���-�:��� �#�y��"���q��D&2ъ�)��פ�y���5��U9N #�0�B���y�"+|q�`Bp�&(�q�ۓ�y� ׮\b� !R��%����'�0�₧�.m��13!�a{�'�8��E�~Qu�a�7�P�Q�'�D�a�FD����Ga�Y+�'T���d�5Y���I�E�h0��'�����.�!�td:�|���R�'��)cCE�{ @]�x;D��'Fܡ�ƍ�c�hh��O��o�����'bv��d��HL�$�Lh*]��'w��B��0o9��t�VRI��j�':�q�V���S��(4� ������yB�zv��q4� �]В������y )Pv�M�7�Y#^�F8���Z��yB���.�kU�*X��� ���y�932�q��!zK��X�-�y2f]&�,�C�äu��\�Y��y@��v_�MI���j���������y��9
�|M	�pv�;���6�y��ex�%bQl��o�Pqm���y
� f�k��E�%�@���݀!d��"O���&��N�v�`�5��<�"O�Pq�)Ͼ%(´z�H	�>��I�g"O��Qe�R�8� v'�w���r"Ox�
G��&l����FQ��"OP���O�):İuEL(�j\Ha"O@5�� h����"�v�\��B"O�dKQ'ċt&�Ҡ ުQZ���"O��g	�*3�^�Ĥ��f#"O�e%�}:�,h3C�1Vz��"O�JG�	�~cPH����bh���"O"U�w�Ie� ��E��_]�iG"OZ�0R���#�2��Q*lCM�C"OT�i�ۭ��Ш�d�Қ��"Od���']t�[�-{��xr"O�-`u��s�j#�/8�n��"OT\xCa��Ѝ��¯&�T�`�"O�� $�7�$I3i]�P�'"O$!�s�W�V>�h0�K.L�N ;�"O()��hG�:�n��!�ӌH�@�A"O�y�,'fI�y�G$����"O���aH��H�&����][�"O�5;g���`�^�SBD�$���"O�D��bE�K\j�R�H��\�\���"O:u@%S:Nr=��N!Z���"O��Iq �)!.�ᡶ�$��h�"Op�A"	��^@�����a��M�3"O0��`
,�Ѓ0�5 �֡�"OL�fo m�v(���*^�x"Ol��RJA��.��#mF�.�6�`�"O<��eQ�ztZce 	���A"Ot�@7�A8]7t�['獻	�U1�"O�A�ѩ�c��=҇�Q6u���"O�l�R�K�<�ҙs�唴��x�"O�t�ߩ^0���"��5�$$re"OF���a6�ɷ�Va���Cv"OX)�툩WH��B؍'���s�"ObՁf�>6i��YQ�]�xr�aS�"O�|(��HgX��aQ?!����1"OH�!a�#m$q��^�(��F"O�Bj̗U�)�AG���-�v"ON����׶�\��d�I�F�B�iP"O�8ڂ�ڨZ ΄PaΕ���i
B"OjXP�	����,��ޘ�!"O>9��E;q��1kΗX��%qG"O�iR��qC� ��1����"O��+�瞶*p���ʊ�}�tDh"O�8����~Cl�� �NC���"O���͡(T����R�F�zc"OD���p��U�&�ζ
�����"O���4j�)����t���r���2"O���,_�3�LS��;U��D��"O&M �j��7�p(�D��{���8�"Oθ�")ةخ�򥄉%/� 	d"O�D���
�r�Z��MpDҵ"O ���H�5�欚"�_!QY֠��"OVh�c��$�����0��uj"O���"j��wjq*���
���A�"O,���F��k�P8�0��5s9$��"Ov@S���J�ʅ��`҄.�n��f"O��$C1=�L5��\�U=P��C"Oxm˲j]@~v�Qs��"N<��ʠ"O�q���ܾ2�XA��U�MT�u"O&�R1��2z5�����LjD��+!"O� �1�ҀD�L)"� Q<$7v ��"O���P�W�->��Jf@�p*
9�"O꼺�A5Qj�#���3��ّ"OҌ�%/�)\���RgL:7"O�Ҥ��TH��9ԣda��p"O���5,N!]LR����]\00;p"O�	��®:XI���!5��0�"OD���J�9y�\e��/J!
n���"Ol!b�fإ"oHqx�`7�d �F"O�Q1��2r���Ӈϓ<&<�� "O�I���B�����=	�Tb3"OB��
�)1}v�;Ǎ��;���"O��r��G6. ���U�wta�Q"O^�����xSV9�'�+ޘ�4"O�5��N�$���gA�9�t��"O
Ո�� .�vPa��@�Wz��+"O�0g[t"F�c��4�� j�"OZ��ߔ]�5�҆Ѝ!ϔTې"Ovu���˵#��kV��n$�B"O�ѹ����b<�e�+%j�YI�"O��0jR;��݁��@;tT\���"O�����G^REI�Q�5G��3@"O~�R�᎜u�h�f��6~>�x	c"Op�W�ͪV�X��Dd�5S\�+T"O���3/�3Gn�a19z�H�U"O97Kǹ����1���+~X!�L�c�8p��&�?j���c�"�5HD!�dލQ��1�F�D�m3���AA��!�$�#~�.��2曵[⑨�oI��!�
�D�Ja����) �u��Λ(D�!�DƺM۔${�Y @�=���p!�=���aF�-[]`}��	J)7!��H�J��\81@Z:2r.��	M5!��H4]�f��%X��`�l�!�D��P�VCp�I+ �� ��U�!��X�#/ a�ǙR�8�R�g�y�!�����2�/Z�aؘ�6g��s�!�d�!w�\	��
N�� {QLb!򄕀w�>�{tDE�U����a��{/!��HX���;7E�-�r�pᮄ�!�.��!ف�
�s�:�@ 臵]�!��؊P�4ǽT�
�:!�	Z�!���-�~�[$�6�bD��鈣�!�d���2<���3��� ��=D!��l>@bc៧1��RA�Q�.(!��$�2��$r=����Q;=!���7�d+��83.��2bĝ�2!����aq��H�:(	eȟ;i�!�ĂZ\"��b�8G����g��(V�!�
P�IC"
������(L!�$�
qbdK 1"��z�Ͼ�!�DE�>d�ʳ*
�����%	? v!��O�,>u�%(A(|�܉W��4h!��C�b=҅���ŧ�����Ʀ�!�ר�h	p���
�"��"ɇ~!��M�p��$e]4/%LI�\g�!���tX����f�D��Y��!�d��O�� cQd�j�Z�8å�U�!��Ģ.yh��dK�5
݈�Ȣ_�&�!�Ňe��Pi�b[83��Q S+�m�!�$S�*=��ȰL� G�>�� �H7-�!��ՠ�(ڢ�ۄQ�h�j�� �!�ӵ&HH�3��`,>�ѳh	>$�!򄃧x���Z�Oݝ' �H�w�]i!�� ��ЖC~�i4�H$P�x���"OԅX�/��vZ�����"O
I"�
|5\�2��ÖH����"O�h���W�v�z����[J���"O�mYr�� htA������D"O�Yp7�/z��Pr6Ӛ8�"O����IE(R4�����H2�]�"OD��$C2d	ʍʇL�>N/r�ʳ"Ob(Xf`Ѡrv6Ms�%�	7z�B�"O���DGʵb�z0��D��@��C"O�FM�I<|����Ɣ5�5a�"Ol4�4�'/���Zp�	�+4B�p"OFz7$��)9��! y��"O,1��^4"&��b#���0챒"O�Y#Ɩ0,������6���#"O�!)eD�4&��Yze��:eG�Y�"O�y�P�b�T��CB2�&9*�"O�5����Ze���7�l� 5"O���Ph�8U�hl9Q�΋@f���"OdL�1`@�B6�NҬ9X�J"O
�1c	�w�|��׬ܒh���*O�5c��@v\`)��H(cؤ�	�'ne�^? ��@k��1^�$��'��*l�r�0�;2B�A8�(��']v�	�cN�t�Z,H�/ "@?0���'[���4��9�^(@AŦI.���'s�鴄Q�6�䴀��ίT�A�'�B��#�mVTḒ�����'7�$hG��%E>��b�]�����'���O�����J�k��	�
�',��KFmL����k��x��'�rP `S�S͢&CB2h�2��'�4tz�e�&H�r�ؘ](@��'UP�+��K&8��&+��Mq:$��'N��S#	��Nli��ӲC��-H�'s��Pb0]��PÔ�ʐ>�d��	�'�qC�I/g,f�24ݲ6G��	�'*����N��<W�I�}��93�';J���+D�/��9���S�p�
��'J�.����T
��y����'���N_�#%-��l-Ԍ�'�4�B͊.N���	]�oMb,J�'���X��"(0Y�@c��h~� ��'f��X�%�2Oyd"Pb��_Zޑ�
�'��s%_!A��b�s���1�y2.�=\����d�ٜp���re����y��>^���Q�)�/`�8�H�bR��yBF�{�(ɺދW!�LS�)C��y�U�o�Z�I2�ĩLu�ړ�L�y���!k���"3@Q2����y"��
,�<��/ѧ*�=A���/�y��1��d�����!�1�E��y���
)�����(�
л�i��y���I9N�;V�ՔZ&��I &���y��S� ���槞�M�1�V�
�yr�B7[���4�6A�l$C��ʾ�yB.׋tjZ�(2 8���r�\��y���I�F��Ҋ�e�N%�$�T��y�O��'c6�Iʭ`[\Ȼ#��1�y�[7B���"%D�
�������y"GY*bl�Q Q*�r�@�j��U �yb�I�|@��*V�Ѱq������̄�yK�a�.U�A��cfDA�ԥ��yRP�,�p�2�&�:O�^82��	��y
� �-�� �}5ȁ�eԖZ�[�"O`X#����8���@`ŏB�Ja�"OTeXa��ix*]s��Hx���F"O��wd�_�dٖNG3���ye"OrA�ɍ5��#�nѻ.��MɆ"O��:����B$:P�F�"�.Km�<I��_5K�<2�"��V���J�ϝP�<�0��Yf�*��K~(	`�B�<�����}��Q���Z\/����[Y�<�Ƅ��<��q`s�60���E�{�<AW�Պ"��V2ѡC�H�/>!�$Ѯ-ΰ���N'�j`*A';!��yϲ̳�=�(�(��5!�D�4t��UҤ㊣:�T<9hM)!򄄭\J<2cm*�B���$!��T+�`1��ƞ��Uˑ`�92�!�۠�8�Y�(P9d���$>��'��� ��U��H�c͍���1�'tD�%b����"�>
8x�{�'�n؁�'ydj�v/%��a�'�0���bV�Z�`���f��b�|���'�ੴ�B	T<����[&[^Vp�<�`���k>"��i�0!$i�UJ�p�<���H�:� ��,M* r��)�)LX�<)0M�jHʅ�l�&�x��s �Q�<���T��|j#�X�M&d����P�<�O^�3�$\ �( ����FDP�<q�k�]������4|�P#it�<��P��IB'��1`!�5�GǃK�<ф��`Y�\�Δ��J�k�r�<�e��,J;,<9�k7"Ur��6�z�<yr�5B4�	�3�X���Ln�<�� N8洔'�C�icr�C��f�<�! 7�����f��y�(�@�_�<�&�ک>V��X2̚g�����R[�<	���5�XmA��@�D��bD�U�<��Ȋ%uj0`�K�V��p�mXQ�<��p ���AB�[�d��׃Ys�<�g��u|�{�j�#j�@p��FU�<�6�R<@���t��O����!AS�<ɀZ�p�d��f�A���ɈM�<�5Ț�Y.�
�B��"��$����R�<)u��/lP��$�+���[��f�<�#�+n֌%㦬W�*�}�'�O{�<��D� 7�����dZl;E�o�<��,����B�iÀ	��CT�<�hK$�|�`۹*L��J�'�i�<!Q�+?��|���_�$���"��g�<鲊��بL(A��T��8\(��Y����3�o���I�&��B�HM��:�X�3�kˆJW6m��:'�����a�x�w	�Kp u9ኹ)>���`Z���蒌u��iY�@�~1,P�ȓ�*�R��Y�`���BM�*/D(d�ʓA��������jBY	U�7D�`p�c�Vd��C�HV��Q`V�5D� 0�Φ�Fp�C�ǰ~��-Qw	 D�<	����EH��1ƙ�-��"D� h��\�_�t
E*�I��c��!D��������T��)�,%�dmH!"!D��kf'.�jѠ2�F B�N�S`�=D�LQQ��-&bz1�#`R�;"a(�M0D���`��.���Ъ��9����F*D�@�񩈕!�^��+t�����)D�� �sFl����4y�&��q봥��"O,u�$�;+3V���ƈ�s���IR"OQ�t�ݍa�R��sg�� �z؂�"O�`Rq��W����f��Ez����"O���_�
�n��e@"mL���"O����.�:i�y�j�#$T�%"O��*2oܤ!G~Ա�Մ:�|DAw"O~��D@Ҥv�x4��T�[�b0�Q"O
8��=�ꅳC�ӟ4@`J�"O<�j
|�H)5� "<�e t�KS�<�2IC �*��RfÜհq3 nk�<�G�z/�z�e�k~��+3H�g�<�M�
S�<��M�j~��b`Hf�<	���g.6}+Ď�;DT��%�c�<a�bQ�dv��eE`<�[F@Lx�<�B`�J�`�uiA�E��A! .
x�<aF��98_�<z���� �b�i�<9�$�p���3K_��U�B�z�<��!�"��@�k
�q�6]1��x�<a'�
;���Hu�N���_�<�J��FԺ��� �X@xi`��G�<y��Y�kv8����+U�ځˠN�D�<1�2%i�$�eGMx;���YZ�<	���/L��5��`͑Vzpc�
^T�<���T�f	B�c�l�d,�O�<)@O3�����zi��R'�A�<a�ժ]���z4�V�9J8Z��V�<Y��Ǧ�l�Yf�;lndaH�H�<�J�n�Q�حB�Y�p�Ck�<a�"^�r��!���2<���}�<aƉI qBz|�t�{EHT/{�<��@ļN��\xBH*�:�{��z�<����q�pc��c��؁R��r�<q���Kz�YI��؍{fB��+�t�<i��\���S`�(�[�q�<y�Ft�i��K��̩���n�<���!	4��k� F"�hA�j�<�%��zyv���ZV6����	�i�<	���k��i�Qn�F*䨃f"�c�<�5@L��Z���~s�S��Ju�<�kЌ�I�� 9FYTE�d̞t�<1��*3��U����4[�L���k�Z�<Qs�ш5�B�0�ʊ2x	\���-�_�<)���c���Y��*XS�Ͳd(�q�<᠄�M,"�٢�ڢC�ʹ��\e�<�Ħ±OW*���'�#	҄x2'�@e�<A��A�O�x�"ㄠ-l��[J�<	à�+U���Nɖ���K��z�<yCfС_S�X)����V`_[�<����r��M����HTJ�iU QQ�<��2c����_�X-~�:`*�O�<�1G����hݙ	mtщ�cU�<��.�:�:��qF��H�@��WP�<��Wh3Ȥ�Ѣ��a�$9I5�M�<igǎ�pN0��f�h�5yקA�<yG���T�fh��� 636]p�LF�<6��-oq��f�ݸ!�xU���D�<��!2$�Ю�5�z�##�w�<9���Y,�`��įO"�D9T	]u�<��K�,�� )(P��-Au$�w�<�ҁ�9�e����(0v2	�(q�<�"�B�Ǧ���΀0�u�D!d�<AW��@ :�8�.�;�8Mӗɀ_�<)!ɍ G�\�b��)�d5��b�Q�<� f�I�C�/[��!�ў-�湓u"O�i���Z32�\�B��[un��"O,���KP�-�Jm+�!jD��e"O����	d4C��2=T1	�"O2���HQ�( h�_�$MF]P�"Ox|)��̮�,�!A^�$E�ɒ"O��ۗ�V�b�i"��$[���&"OU �θo�\V�.k��X��&�\�<)r�Z(0v4��+�+T����]�<��� �OHQ�GL�\T&�8�[�<����0N�B��q��<0w.�P�b[V�<�5�X܈��ϒ4oR ��õ�!�D��EFV��6D$�|yrdm�9C�!�6e�LtjO��;4*�y����n�!�D� p�b �֤ܹx��Q�G\�Y!��!#�F%@'�S�6g��ЁmL��!�$Ϻ����U�_��(�� 
�n!�ƭ�F��|?�9��N+8S!���E\�{���b����FH�*?!�d^)&:8�S�-9]�1����?7!���_n	h�[?i����^�Q#!�$�5*L��G�.���5�؏n!�䒞F��ȧ@�#���h5��4a!�$ױ((,�8V"\�6�v��e���t�!�DQ�@56�ҫ"��DK��g�!�d���Yc�z:�]���Z	F!�6^5�2�/V$|�7jʖH!��4c�b�#��/eP�ɳh��G(!�� e>D�o�Ne�����!�,|�F�Q��1R�!2"O�s�!��BH�����$<��A�φ$K�!�K�H�01� #�T��#R�!�̃H?J�sEk�)Zj���
�!�Ę�g6r�iթD�
��h����4!���kjx�زd��P0WgZ}!�dN'o!p��.�#W�pȠFP7y�!��ۨ���[�a��U� ��ex!���([wZ��"��0��jv䀑Q<!��P�\dԢT���Bu���!��'-�p�����@iV҄�&d!��>X�Tw�
H4�+� �4M!�Wuh���T�B�-�3�S�m!�$!�{�e�'+(cu�Nn!�Lul�3GM�*R �Qc�0�!��d��`�Ӏh��6���y�!��)S\A���;+��J��;�!��@��X�L^9��B�� ;�!�D�v⬘��	"������R�	�!�dI��\����W-�$����#,B!�J�z~�E�%
�x��0��'A!��O�Li�(��#�@�@�I�.!�dJ�N�v��&j[�u+ш�L.F!�N,Mf<3��?:]Uf��^2!�DT�U!���qO�J��|��X x!��n�6�J�.Ǐ�耺D�A	j�!�d�d� ڧ��;�� ���~�!�DE�E���u)��E�Ԩ�Q�!�Ą�����U41{��g"�!�dZ�G8�c *C�-i�q��G�!��v]��a�a_r1�6�y�!��KaM� �Y 2� ��Si�Gw!�$�%b���jWʁ�utX�v(�(Z{!�ā�-S��@�q\:-�����%�!�d�W���i�;Np� kP�O�!�� J�qE��4$�ju�P&n�Y�"OR�;�-<m�R�uEםP���"O�=����Ez�T���µ�����"O2��E�Q >0�f��cX�� "O^5�@ �`����' S>Yi(Yf"OR�����CwƁ�� F	9U��*"O�P��[�"�Q0��(/�Ax�"O�1A�f��1���'fL�J�X�"O0�h1K�5�$xC�*��I!�"O��I�bڝH������ߍ$�� �0"Ol͚��	|mlIbT�O��$��"O��puE\�t�7C��0Y�)"O�S'�՝- �H�cCV�+P�<�"OJt# 	�!l� �Ӷ�	Q10���"O�����~�D,�`�ӱ0Q�"O���MA�pS��h���*���1"O<���� byrE�T=@i(��"O��a��&{�ikpk�[a��c�"O�8Ks�M�Y�T� b�AWFl1�U"O
���Ο�V����d���I7���@"O�y�%K��4���#�ƥG'~�CQ"O����7�py�cd��2����"O���CB�B�T�P�J8Q`U"O��J�A�$z5�0h3��!�����"Ou��F^�a#�(P�H� M�죷"O�ݘ���9�H��D�
�D���"O yy�`�bT���ĮP�%���	�"O6��6�����NC�a�f3p"OHe{pF�6X����C��7:���"O��a�ժ��؃�L�O��`�W"Oj�K)�0�|��rl�$L���"OP|9u�͊z�:�:�jJ�0�81�"O�ā�,u��@©ȵ5wС��"O��Z�A
�<����(�:XV6��'"O�#sJY�t�xq�d皽h;Ɂf"O��֨KpC��BS$C�X<��r"OB�� 	�Bzi�! �!
�"Oz-٭Vylu�� �#�(x v"O^��bٿ/Ų$*R�Q;k�n8�C"O�(S��+p\�z��L�A����"O���G��K�0;`��%��\�u"O�KF�W�]���6��i|Ujb"O�ѻ����Q�#o�!
ٔ�AS"O�l8�dȍmmP5 E��/��0��"O�� �%U�e�Z��� N=]�<ۓ"O�]KClK N����*vZ��"O�\��ذ)��h�o�	aZzE��"Ob�	REɩ

"�@�L��;WF8P�"O��3�Àqs-��IX8"b�yR"O��[AJ^�����G����2�"O6�C�*3�8�@@�Bj��80"O5��lT���!-�`��;"O�8����8��P���#c�����"OȹI�-��nL|��T�q�,(`"O�H3%�@E�d��Z�����"O�	W�^�C=�|�F�CVx���"Of�2U'L8](T��$*�X̊�"O���3�	�+*H��$X�k���Q"OZMxvb�1Q�� �$l8�"O�l�'���V���*�k�t�"O|����8u�x�+sIʥU����"O(�S��\i�Ε�3�\Q�P%;�"O�tq"���9,N���Ɓ�/�<��"Od���nѭ*�(LPD%�4�`"O� �{UJ�HLT�aW�/�h	�"O؄+��ӑ��E8!��l����"O�9S�"lVFYy�Ϙ?Y�Ԕ˶"Ofl�Co�$gi�HQa�1Ơ��"O����˙�o�Z�s�.QR笽��"O�X�ħ��H�b�&Q?�F�!�"O��zf��Q�z�{��ْd���""OX0Xw��h��`�n)o� {�"O��c���*������|�y�"O����(S3�z���-ʼC#�i�p"O�k��(>�u��ۘi���� "O�j��V���$RD�ʄE����v"O!��
8\�9Y�j�>U``"O\�2Q��=:P5crkM�C��\0�"OP��e��m݄�3ר@�!e$;r"O�٨�eC(H�lU�և�[R��"O�1��C��c�$�r���GBTyR"O|X�PN����Y��#&}'"O���q*�
k
��Ӫ�ep�7"O05�a WkM�M
���$��Q�u"O4D�p��?c�����-� |�"O �3�&єK�E;���{ک�P"O����a�@�E�恒q`�5p6"O���u�ˬ&V���C��;L|=�"O()g
�"�����Ɵ� �#"O֡:%���P�d1蟢0�d���"O����b���9�0��$1�6q�q"O���d�V��`�H�3k�~p�r"OX�#�.�%[k�M�f[(q�ڑK�"O�|��һ>�n��� ����A"OzS��Q�!�*rӦ��B��<�0"OZY�#W��،��%�2��"O���	A�@S���/��(8b9�3"Ol�go��KKJ-C�F1x��"O�ڂ��)*��k��V�& �D"O��c	ɏ#�,��ň�X r���"O�� Ũ�<b�<]�E�
��u��"OD�I  Q�N眑����_�x�"O|�
�m���s%��?\��P"O|5����2o^��F��%-�&3E"OT��bE˲e|@��P;P��h'"Op��%���u���]�
,��"O�1"�m-Q�aCsm���$�#"O�x�u�S�q��-����+x*X r"O�Y�P���,&��33U��&i��"O��ZRN��Y��E�AB�^-�@"O����cƮvcp�	��V=V0���"O�5�`�A	5��
c��1y�!"Of �' ѡB�|�hCf��!g�|��"O��۹M�4�&_
f��ux�"OX�Aȓ8T \	�b�"w�D��"OF�P�,��|T���	>�8�"O~�۳d��@�,��dS蓡"O�a
QF
�M�E��D3gF4�yR�ۣ��؉�L	��M G���yBNǱ=�f ��?6�4	��LP:�yRȏ�c�x9W��>6����M�$�y�-�$[|k1)����xr���y��e��h�HT����ÂU>�yb�x���w���
� `�t�R�y���q&�1�E�<����y2��b��l�����p
B��Gʌ�y��B�?Vr��0d2a���R@N^�y�O��|���HqH `�����_��y
� ���,��v�����#�"O�YYr�A�Jl@ca��qL�8b"O���Ď�&AV<�7J�����H�"O��g��>\��d0�hC�
���"O��
�6fS������\ *�ZU"OH|����t�Є���j@"O��
2kÙ{-,��IQ�9�r�+"O��`�%�uCDxAbݢ@�<90�"O�M��nۙm/V�ʷA��l�z���"O�%a�)9�4�v*��&;b�w"Of]��N	;1!����T���"O
�rca2t��%)�ȏI��ȷ"Ol� �$¶v붽��FT�e���i�"O���9�`X�e哷e�����"O��� ;~bL���?5��Q9�"O�;��߶^�j�!��$���S"O�a�B딧Z|JmP*�x�.l�"O��,��I�i�EHJ�l|�k�"O&����<�2�+�hD�Qż���"OL�:�Ϥg �`Sr�B�K�hX��"O���#�ׂDNX)�b�@�q1
�"O��r�CC�O��xa&��O��sc"O
�Q���t��rp�B�[�eJ�"O��փ׵ r�3���Y��"O�
��0 �a�φ$d�H�0"O��9@eޞx{R�z�(�\W��+�"O�P���� ��8f�"Ot���/(./�	�E�F�7� �C"O��J7~�P)��j

ch�K�"O 4�-
�Ʀ���*��x� 5�"ON%���v������ ���"O@�K]�g�p��D%�d���"O�Q�bP;O�e��'ԾQ��b"O�c�@��@5��!ͅ���{"O쀓���9Ii�\K �Dn�EP"O��:u�a��� �H��p"O�(��$�9%bVlP��=
�D�XC"O�:��C�	>�ٙ6��<"\q/�y�޼Ts0�ar╆,h�k�`��y��'*S�!��G�,�7�ߖ�y��O�>����%'�, ���(�yR��y�z�J��ʳM������Y��y2�,�. 0��;�@IC�G�yRcU78���0�'��w���yB����� F���8����*�y£�#`b�H�U�A��F,{6����y�&X�V�r�-��0�%�J �y��EY����QlJ3}]���

��y�c�>>�aVf�r�&1���A��y�GJ�����d|���Ğ�y��׳���F	��_J ��%���y�.��{6R\
�I�L�h!��Eɟ�yn	�$�(L���N���L�P!��y���]�zy�r��|-��h@1�yr��BJ��cˇx�%qP/â�y��Y���{��=CY�j�C��y��Է�R,�!���68@}�lޡ�y�
I4f	�P��C�.^�d�yt��-�y�$�3#z�]#q��X�rG�\��y"7R�p��@��:TN��XS�)�y���4J)"w���M�`1c���y"��Hl�0u81��J��G-�y����"6^x>
`R�f��yb"��n � �f*��u��tj��@��y
� :��v��#m�!BTL�U��%"OD��ggP"��� ��NP��r�"O>ɢ��R.Y/����XH��"O.Q"��ͭT��P���0�T��"O8D�gc�"�P��G
�^�䵋"Ox�z�/ȓX&��� |l�i"O�Q�Dʐ�����Δ�|r���D>�'X��Yxu��hԤ�K7.�1jք��I�D���I:��,P�Y�]���ϓ�y"��%kzj�#`X�	u2�z�[.%�C��f�t��FH�t�� �$�S�v�h�	Ϧ�J��|�i�Ap�eG�}�`j'G˕/��uk��8D����c��	6��p�1ȖIHR+�>����n�| H'���YAD�E��8"=��Ar�����	N%�RӦ	�$y�� ږ�!�䅙_w8�#gԻ1e�UFNA�����I�8'���� �\L�$J# B�	�2����RPqL<cD�ջ����X~��'�f%Z�,T6f�@�٧#�1Gqذ ����$�lh�ae��{P���قzw�'2ў�>�It-�E(�i\�/�$/-?)?�de�O�,�x�!T+pBJ̒��e��M9�y��'�z0 �cO1b�~	xV�˪]���+ON�=�~��48X1�h�}�&%3�cM����ȓ H��2� �]=�� ��52�|�ȓ3?�@�5��#<:��b���d���D|R�i��Op�Ss���A���u�`���.
7�FB�I�2�`(qfX_vȒ���1����hO�>-��)�&ae���7MG�u~�9t�1D�L�EGK�=\T+7M:8E �5D�0�3.@~o6�"�Â-,ް�S�7D��pǎJ��b y9Ո�+#�	D���'19�ء��) b<�6/ԙ`����#n�l0���1g�:!Y<s̹�ȓo_*1r����h%��'^�F~8h�ȓ��dL��7є��ֵ����s��j$���0%����j���;U�;D�8!��^�.6�\S�,�,d�A�n����ɐ2+�d��N�YA�zcMx�O����ÚwR�#��\H�&ASCe�P�!��X�8=�ٙ�W�o���4/
P!�d�"3�xг��Ȩ�ޑ�n�l>џPF�D��!��(e.��:���QfƑ�Gў"~�rž���
K�T8���$]�m��A�ȓ*��U���B, �@��A�J@�<m��U<���L�(ƞ�a�E�r�d��#J�K��?��ĝa�:�,ap5������r�=�@B䉂T�*���)�	�R	��H�;)7�B�I0���dEC�R&��b�dڦw��B�	�,��)1Jբ���!eY�C�I�b���jV<\�`��$,�\~��y�*�<E�4�ʿ��-
��9W�����]��yb�'��l�TM
�<�x�Gʑ�f���R>O:�=�'�PM؇'G�z�$aHn��g��C�	QC.)+�&<s/& ����@6�	R�����=�1���Jm�7�[�M�P�'��O��WL��q�'�S�*���"O��#J��v���V��F��� "O$u��@O�J;�8	��"T���"Of�b�( �J,�peN7�}+�"O��`�2��$�n��TXА�"O��r��՛���4]�4�2"O`����r���-��%��X�"O�u���ۄ6%~�����$R��2"O� ���F���S��.��9��x2�'�� CƜ�i����҅ɓ.7F(��J��	�6��5`���s"�8K#��lB䉏.B��)�=W\������CB�I�#��X�I�&I�M���`:B�I�D�d@��� Z�f���l��'�VB�<~��0"��E�;�"�Zgl��9�2B�	3(�8y����S;@a�$Y�n�����>Y�e[	�"e�%?g<��hx�<�`�"u�)��;����� �����q�)ڧY ��G�na M��#�E����IF�I�Rz���6%*~L�с lH|��=?�ܴ��~�<ᤡ�5����'��o^���En�'�ў�Sd���W��)W$Zj��!Ƞ�@"D�BH<y����G��*@�)"elh1�ˀB�Ii��h�z #V͂;U�6�ªN>^2��'��I:�t�y�E���� ,��V�c�n�N�'!�'k�`b�蟴kyV�yf�׻@�$9��dp�f�'�1���@u愬&�T�ss&��k����"Ob�!Q�Z�?�.�9�&v.�xg��=�Şe.xp��B]�(�ʀ�L2o'�KpOr��"�ʔ6�x���6������'�B�O�b��T�
%S���#��(tVz��4)4D�ؒ$��?F-�Ek���u Bq1��-x���hO1�x�C��`H-�է�$�8���Z�O��S�K]PHɓ��g�X9(�y��)�3q�<�鴉ßi(�bEB��D����#�S�O���.
�c��H�E� :�z�"O�q�R�W2�M)���i !�'gqO.��b	Ӯ,�n�0�R.�eK#"O��#��c�qU�.I�e��X���iB�j�E� RDc�Y	��(�!��ýKG2@��Jw���Y��/�!��ΐGF����5��(��
�M�!��<|�hȑ��6Q���ĬE7!�D���C�h�d	�E�^�!򄜝i�2XQ�5BQ��D��c�!��A�[F�<1R�A�=
��D�zk!�
P�:��s�~d�0m��>[!�D\*K͔��AL�*d�Řo!��-�2�k�'F�x�����ˍ�#��T2��)��H�`�B�!�b\�E�Are=D��p�էvz��g�Q�#%��pGz��	�)��k�.
-?i ���,R  n��d5}��<�9��M��h��(Ѡ�yR�ҢLy�%���-@.��z��y&+��hȷ�5/�\IP��?�y�N�d��2�v��왒� �:���=E�G��d�Y1�_�Iޙ� E�P�0$HvOЩ+7���j���ɅV��b�"O>�ˢ*��g�4�zEZ;_M�{0"O��u�Wq����0��!YD�'�'�`���	�eK�uhH�;�����'R
�hQU�t�)"�^&i�"8CM�d���'��O�AbT�(q��T[5Ĉ�bp��O^����0��\8��Sh��2$UV��K�l0�
�_��@
�ヨ;P
%Z6�<D��c�̟0u���PBI\!���ƃ{�\C�	�?�Hx�D	ɱ|E^ *��,r-�C�	�v�I�`��A�(����L�_� ��$&�- (p���f��I�A�;`(��R����Ye|p�O���̓�?�c��%��,�7�;%���7gɲ!�C�I1b���ąQ�<��U*�g[/"�㞘��)� ��R%�7 ��b�ߌZ֎�"Oxe�B�
]�V-HE�d��9:�"Ob�J ��'�������D�u"Op�*���Fx���y�i��"O�v�O2',4p������@�"O�X+��^�+�����@�)i�D��'��L�c�yX@s�⌇/�����'����C���b)z�DH&w�J,[�'�v4���G*�k��Qq��'�du ����eD<�H�h�{�'�dCA�jdbx; �4a��9��'{�(GL\�E%6�K��1
�\<�
�'8��c���Y;
��#L6��,z�'���Z�,��uEnP�rD��=�*�'��1b��$'�` Y!��Ot�1�'�����ưv�4�0g�}�8Q�'l`ґm�^=ޙ�4@֯+O�r�'�P�㛜$��@��)�:D2�'p�-sT���A��D�O��'_�H�TI\7��*c�E&���{�'��KA��C2����R�'T��("�
$:��H�V�ΆLNM��'
x�Ω:㈄��M�6Z�4��'Lv�8��Nn�*���,҅�y���|�P����PY�t���y��NW�@��R���[��
6�y��Sָ�;��_DZ�%KP�ª�y҄�!f`��%���K&�Ӱn�&�y��Cql���3"�F�a�� �y�o�q16� W�P;yZ@ P�R��yb)L����v���+�8Y{�dڽ�y�o�-)��t��d� ��<!��y̌��84e�6��Wm&�y�$��s�騖/�~�X�S"�@��y2`É%g��y���� �0 �1�5�yrMӧq/�̛�ŀ�fݞ�z�� �ybZ�;%R��3jƑy���"̨�yoNpu��3񆂋 �;7��y�fY8�ؤ���;}�40���(�yrk· p���->�C51�y2ߛ1Y����,;�T=�Dfѻ�yrF�b�6�)��J��<"�FU:�ybύ�gH��Q$ȍ@���2�D"�y��[_�I!m�5o�������ybC��(T��/1d��ThAħ�ybb�K4d(Y��J��#��(�yc��!
�{C&4<�T:�OV��y�Ð"�6���.�:��P��*��y¬�"�2Xhc��;� �GO��y""G�R.�����>&�h%��A���y����b��Y�N ݹ�i���y�'0�������ژ�`�ϐ��y���1sA"ݐ����l�u��6�yR"ߨ*
 T��~H�;5F��yb��=(�䠳�V5��� �/Z��yR'T�5�P㒥z��Р'��y/\�9��A��B�kB�L����3�y�Fˮz�LX��ޗ9����FJ��yR�ߘ":��뱀5Ҭ�AHW2�y"�[3X��sBZ�
f5Id�ѩ�y���oj�o�7Z6@�Wj�	�!�*r�c@�D��P��-�!�d�6&b�Ȕl[7g@pe��=p�!���4�䉱A����B�N�|f!�� n-:D�A�)�f�Y��^7ITTjW"O�1R�@#iJ^��C'3E��\��"O��S��`��ZCG�1(���7"O��֮�0~�(ӄ�g����"O���*���UH3ރ)-n0�"OH�['Ǜ�7ofp"`�[%=2D"O�aN�-ar��O׸#��Ѳp�'�!�D\�z�F1Z��G;V:)#���c!�˓��,�;b�¹����9��Eӎ��#�u�(Θ�|��u�w��*��X���|�FK&���pf�#Ux�=��z�JC�,HY��]K�zl��\��|�
��y"��X��Н
�H)���y�i\ў��Z9+h#I�X!�X��i1"O8�P�(���Ø+�*=�S��*�S�S�c���S�a�P(D��:y��C�	�y���+ݫ{$@�`BW2B�If�e9�(�XK�pT��/{�B��A_Q��c��6�ҷ�.0��B�	's��]���ݝ��SB(N��'Cў� �4�ē_�Eb��b�z(B�V�^�*�ȓ�2��*��hT�i2*�pG�t���ƍ�r�O�@pV����T.�q��fl4l)�lת%}�0����%M2D�t�5c���(��;V�*�á�/D�|�D	��#tб���~T(#g�(D�x`�!̳sA`��#L�>S� ��1(OB�=I�F+ ���e@��c���r�<I'��Q:�(Q��j�x�a��T�-�O8��Pô������36���j"O2͓�@Y�.����ɆV���d"O&����0Ȣ�h��;���Rv"O�ahA��7�!��E
>��� ""OԴ���0��������m6�xx"O�Xj�gI; `U;"gD3�&y�T�h����R��|��F�2��4�3���ePpB�! N��J��Z�A�d��r�1ڤC�I�h�>��͒�riy�n��9�PB�	��5��D,n!N�i���%`tB䉿y�Ee��?� E2����XB�I�AipY�0 ��3����b���p?���lɲ���ŗK�� ��ƛZ}��'�aj��ő P4i�/�Q��H�'��L��K ��6�C��Q�l��ē֥C���D�v���#I�_�͆ȓ+�܄�uh@!E�,���SuX�ȓ!�pʶ�-0H�����d7��	r����ucU�Xo"�iCҭ ��إ`���>q
�R2�څE�,�8 �g�J�+T���M[(��sU�,�Tݹ�ILPF4��W�XI�I�$��`�!��9{�Y�ȓ(:���ۮ􆄀�lV�PDPn�������N�u�X����
�ГҬE��yb[�F��00tK�Kbe���y2�ͨc�D�ӥ�E&{�����&���R���OS�9C�K�-d�x|qW�Q�v�"�	
�'����BʼIV����K��T� 	�'p�����x�j��푤�F�	�Ø'�" R4��n/��H�o���Ľ�M>ُ��	B(w��v�����r��J<�!��B4e F c�aW(lc`���E6:6!�۪nȁ�5K��hf�L�� �;!�'5a|�M-OC�H���J}Ug9�y���:$J��anFB�x܈�G�*��O�(y��� ����	�&Kh :�D#U��"OX�a�)5�!�O*`��x{4"O~���o���� WHS!c�v��0"Ov������h�H�(��-v���RQ"O�!��:���QeFL�d�x�"O����	�
�2����ʀ=���T"O��֫F�t鶙`����v�QqT"OD��po���Ba���KT�%Zg"Oh��#(R�LuF ��+J~Ȅ�"O�8�NE�o�5�R��,�n���"O�����^��2c�F��Lh+�"O|����!@��$9d�n�^P��ėb?i,O����S���dD�j���@�чSl�<ר�5JF!��7��ʐ!�~^��� t��b�Hz������ռ�C��\�E�Ӣ���O�"~b���J�P����4��(���d��~b�T>�<=�}I�J��b1�Xi�D�F��}�'κ]a��
�͠�[!��5V~Q(�[�T�V��y�˃�W�T�0WH@"����Gd�%ͨO�"�4��(�~ѳR�Z�p�v��g�@e�<�t�M�L�dyc*�T(�	r�JX��Ey2�����ؕ,!/+ ������0<Q��$y��������Z֋;WdEbT�'ў"~ʃ�#z���Ti�+2
����'Nў���=��c��I5: Rk�:2-x7"O�˂�/Y�	�)�=)|���x��i>��O5������ԡE^�,�)�"O�1dEA9��3F �{�����$�S��'\۠�`Ą�)9��9PcF*kR�B䉃k�$B�d�'+���ADT�Dm��=a�'�b��N�m��VF�*��%�c"O�ٱ�NG%=Y`\9��+2⁬)�Io؞��A��iK�M�::�
}�p�(�	�ExҘ>A)��"\�U��[!/�4�Ae�I�<a�� RU�0�Vk� Q���B��L�'ba�$%��,d���5@�mt}Y#d��yb�ɆP74����N��H��GH��y��G�#}Jy �+�-���h	�yR�">|�[N($u�P-	�y2�ߟH&���H�6XBD�	s�����hOq��&M����	�JX؝i�W�������-� X�9��M�B�-Z5���sG��~'F,31	>7B��&�a1G�F�a$ta�#�[�.C�If�$�ar�C�$*Rq��+G��B��80-��š��a_�A�n�XV�B�	0[<��ɶO�>8M���O8:�B�	�c��B��8���璂k�ZC�	9t�yS�*��*團e�<��$r�x�'��́���Sgy�qm
/K�ͱ���;�']�%��)p��Xn���@���6�@ڥe��ZX���_^|P��:7��҆]�~O���"#�(x憈�ȓ��$�����9�w�Z�CFzb�'j^����ݎH�$�
c��73a�B�'P�q"�o�^8S�N�$`b��'�`��g�j@"�ѣ�k�btK˓���~b�j�����ˑ�S�����yR�EDT����BD7(�35���yb�Fx�$� Ѣ�A2����C��y�fO	y�D*�P��hݲ#���	���N>��	�l���z\��DaG�<Y�C
�O����@�m�*�z�-�D���=	L�:"xh��X�]��`�v�XE(<��I,� �h�6H�T;Qyvɹ�"O��z�.�$/�p���V(n���x��'Y$⟼1�B]��n����YX�0a��9D���k�F�~eѧ�����ht�%D���ï�	:��X�1f��B5���@�&D� �P���u�'$�!J�\��A�?D�;�	ݤt,-��D��~.HZ�0D����dW!'?ʭ:B��˃b,D����Ņ5k ��O�<E=��e5D���@$dN�〒�9�ȫ	 D����KF>�nH����.�p!�>D�S� ���& �Q�@PC*D��
�Ñ0D8ʤi�d�����d�&D��@�����K���2��h6�&D��y%�τW���Í]#|�e�0D�[U�ÔM!]i"��L.��#2D��#��M� �(�U�-a+��.D�����ʡy��%�O�Sb��E$.D��1_5�ty�Ŋ׮���c����yr�Z���
��1n	T���cL��y�I��W��5���	�^#)��br!�'�
�x�l[G��I"���r�.$��'�4�u&��ҹ�G+G�m5l1��'p2��V,Ł'�u��i��g�Ź�'i6�A )[�?+H��a.�2(����
�'N0	t�3l(�S&�#)���'s��{#)	1��$��b��٨�'�J(������a��@>[����
�'�`�v�n5hc0$�� ���X	�'8$0�b�W��� O�w � ;	�'��|Iq#� w�����B��7S�0z�'X~����Ͱm\��� G- ���'�y��%Tcn���S�ʭ+@�{�'d�Xuݱ#�Ƀ�!V$?<�I�'x&�򠊟E�4}�BI�E����'I\ݑAn���j@�2�S�o2��'>�a�� �>OJ�%[�#��li��j�'�`Ii'��4zn�A`�.pz�8"	�'B���!�ڠB&fɀ�|pt��'����D/��<��H[͜�zT�a�'����bl�:O)y���#���p�'�0��faF&TG�a���1v��0���?kxX:�D�1�` g�'��`T��"Yg��)��nG�51�'9n�6I�w>x�@`�a����'5���H�g�b���Dͬ�N��'�"����Џ/6�e��l�x��
�'��\c!���l��M��kE�sn��K
�'�l�
�C��gp���
5`�6)z	�']b sM2I,@xH愝3e�8m��'�"��*�GF �hfM)_���	�'�J;��&U:\�Jɰ=񀬱	�'��P�Vi&7���s�Rx� 
�'_ �H�儶V%"�	��A��
�'�N�!��CJ3H�[�)*!rօ�
�'�� �ڵv� |	C��2!q	�'�R��m�Cu�,�!�E�-b���'�h}�"��	��X�J(ݫ�'qH����~9ĈhQM����'ޤ<	�X,?e6�)s� r�t�z�'w`��µ]����"�o~��
�'��A�K�e��"b�:�*	�'�HrI1�8e���W�(�'���Y���,c�"�.�ܴ��'�T$kah����A�&ōd ������ $�r�՞���=#�.��"O4�����He��ߤ�����"O�j��]}�L)kV�B�:I9"OLR��Q�,�"|@�B.Hٺs"O��y���p]��;�f� �����"O<�3 d�tMIw�K4;��J���]���'a[�qRVB�<m����Z����QT~���-M�ը�
�EM�Dɑ�)O�a��	x�������7b[̐QOnɂ�G�A�!����%��I92�:y~�B��V�����$s�lb� I% �~C��,Wx�sEŏ,	d��q*��38C�i�qI�ęu�L��զ�=D\C����}��_"�P��
�	� 㞠Q"�JDX���,�nC��:����z\��R�0��"LOZ�1fEF[w*�g"I�j��I�-}-j@��}/��^�Xu����v����ň#a`ax�J��`�R��=Y�����m��叀o�4X�@iWl�'��"~�L���1rѣ?v���r��p~�B��y�l!�=E�Tnظ`|�A�b#]5}��E��+Ę�~"L�W��h��t��lոb�-2�S�L��8V�䓅G�� �5�QqD臮��Q���*h�O�I��0�M�  ^�_�,�x CG�?�������9���č?�y� �:�����j�;4�<}�gE��p<q�����'��@dLK�n��\`�*҅u<�5���Nƈ���p��W
��q�
�~3f���"O���ʛ�9,*M�M.	�����O��A����%�\
5� ��B3�! �
C�� Pgv��P�	`�@����!;���'�D���I�/;�S��C�S�(��î�aR���<)S�I�T�H����.,�:�E�R�<�̉^te��H�H�@}ڧ��D�'Ț�D���՛Y��*�C��vϼݳ�C��y��{��A@4�`�h�E���~�oc��h��	Sm�A��-�cI("{t�"O$�Ҏ�(�|$���8�@�%�>Y��1�O̊�gп^̈�Z憑pڒTz#�'��̓Y����&	̝i��`i!J�@��u�J1���μ�i! Ⴣ~���G}b��c�O�~�g
f)�v�ݓy���x�'�b�2� �.'�qjG��y�f\�'�p1Ey��)�&3�!�6)_	�d��6�	4�!��4X�ѓ��A�X��vES�P&�'�z�����^���g��DL��kg��0Fa�(b���k�4%\}����p#B>D�d��i�q=*���D�.���ô�2����&�+�L�{�����'Z�J�f"O�uۀj���(��P)��`�Q"O�5��%�)�$�ѻ����"Oąv��0FdԅE�UHѶ|��"O�M����):y�,�����"O��ij��;G ��9�V� �*O���珓�w&iY@ĕ�wdtxR
�'O�\���#j��@"C2e��		�'��9���}��!;7�+"��'*�(�L��<�
W`��H�	�'�.݁PN��[0�Uj୔f��;	�'G6���j�#�@9ve�E��%~�<���L7?I04�)��P�ș���Xx�<�'%K1)�޼B��7'�T�䧟v�<�T �*����b)D1�}q��u�<#j(�Fi2�-H5�������l�<�!��
�=���KK�bT��BC�<9�N�m� J�V8�p�"+�|�<� ^��DCL'Q��Y���{���;�"OT����Ȱ2l"I��KV�;�`��1"Oh8�PI�'��\�����+�D�U"O��B��EDD��a\��D��"Ox������p����V� P"OD�g�]�-���2��;{��졡"OXܨW��"3v�Ur�ڛ9X��"O�����ՄJ*�8WE��H�0-1"O�\����0�T�����]�l�0�"O���O�;oO�R��J{x�3"O�1rۡ�����?7��`�"Ord����o�V��k�#�t��"O��A"�@�J,(�Ѫ� �x�"OF��u$�c��e���N>#wF��"O��й��,s���8d�:�"O(��&Y�X�"[���'�  !�"O0ԋ�0`$)�g�`4�p"O����1d�p�E!	�ɲ"O่2��#̾�R��X;���
u"O��B�GY)H��w�ԫR��a@"O��v�V�.($@���+eτ�xt"O|��W �%�B䑗�[.�0��"O $Z��2V����g���;�"O��qM;b�Z�:E��$J���"O�:3l�E�Mz�!����B"O�ٹ�ƛiSF�s��^����"O�5�7��3`c��;o��'
B��"O<�To�( u��#H0K�*OT�(�	3�l$K�_�bb�da�'!Z�3�[�y���Q�5]4n,��'����sĎ�MY"����Ȃ;���'��3�@M�%|�H�3��#?�T1�'XZ	R�O֐v���{�g]4�:�'���1t��uU&6e,�)
�'�� j��m�0L�.f��YX
�'n|�����(EΥi���[.�+	�'�l���!	��u�rM]����'�Z�̈J�e��I!9hlU �'�m�7��@�`u��!�e�D��y���e�F���=h$�RO�)���G'��V��C�I�uP��%i
�(`$�9dC䉍j�Hi��b�}����
�)B�xC�I|�<!P���$�� ��l�d�vB䉳V��}�1i��s��H�T�G!i�B�I�	���sF�[]�tx&�\^PC�	����	�r�]8�Ћy�� #!���x��L �B��i˛u�>��lǀ��O � 4�W�IYڨcM~Jc��T�z��7�\��g��K�<aU�T	����S.)Q�!��<y��H h�6���"�t�)�1j B�䙉�A6�V�S�($�ȓ;����ވ*�H�9"���"��o���2鄟!w�$��KQ�:�"=�ݏz�,�P"��6[�a2G�����D�����7
B�8�!cKQ�OC&y9�C�+�j]�c��3��<9��� L��R#%� ����QC�0G]��<�ҍP%�t����@F\Ѹ1T>:���	mi�y�oX}l���)}2�'��\P�-È/�X`:�=S��arNM�T�8���D$���Q'�>��O�=�q��H�t
q�ع4��J�"Od�"r S��\q��M^+`���* 4a
an��J���貦��d��3��ߙp�,Ψ@��( ��L�k�0��c/�O�!����9,J냤 :5���ee&/_@�C��ِ3D���[T�Gz���$��(j��R�zE%�:�(O��C����!��@��)�^�Ze�~�0��#c� �A�LX�~�R }��<�O�嘅��69n������]��*$��X�0p�CfN�[6�ـ�i*@���D��;H|��SA�$W�̒sF��Z��M��S�? ������  �<���_�_��Q7��]De@�2~���EK��p��	3ғ3������6$����V�)�pt���2�`D�A�ͪ{y�9�Q�� u�����*A�uVu##LX��z'�jX���������ӧ`�^JK�H�Q�$��k�9%�������rR�WR�4��&EF h��$j�&h��̔.�yB�Q06�0��U�ܴݼ�1�,N�Ot{��CX|�e+q횚P��d�d��Oh��FE 4f*�� �×��Hi�"O��H��W�)�Ј�p�PSU2IR�G	E�(�؜� �Q�W\"ij�W?#=��[_��0X$�Cz�� PX�(�g�� #t�h�� [1Y	�+ F����l�,ذ�U��0?�7����A��a�5C�^�j�"�I�''�� qF�t�z`�%��V����!�����­ԼM$��;2�C�I@�L �a �=���J�nR�y��I�p  �3�ݮV� ���!)����p&����"��ה"�ڸ�w"OBdF����c��E1Jb&<?!��֑�d� �>����[7-:���5\8X���=��?����7,l�w��3�����`O�:ɠ�q���x��0%H�����/{b��F��y�j�,x�Xj�&�kӉ��y�,�~�0���J�	�F��� ��y���7x�� ��� rh�W�0�y��B�xǺ���iG�{�>d#���yR�];`w � �ң;p����	��y�Cq�Y"�ˁ>WD�
�`���y2h�r�D<Q�Y���S����yBf��8x�\���C��8�ÍN	�y�M̽%��	�C�9]�l��%� �y�F9[<�Řs�_G�pղ3jU��y��$U��pz� P�/�tA��i�ybB
bxq�FC�$X��2�դ�y"73�u��.�Z�B�HW��y���-�����9SL�v&K �y�J�H�TA� P<��BN
�y���7\S�Q��ny�z��S�ʾ�y$�i�.����qj�kc�y҃�c�6tSv�]>��������y��Z��5@�5�aӖ���y"L��H�,H��)�rg:�#&��yđ>W����XQ`�����y�$#K�f�`%�� �+O��y��I�Q2|4~� <5���yB�[tO
a�$��"�<h�5/��y2g�.�* ��j��,D����
�y"L^�	��x��̌'� Qq����y��R�0���hFI���Ǭ�'�y��ΊV��rt�E���b�����yb���i@���<i��ɓd���y�ԴF8(�R�+�8��
��F��y�Bǟ$jD ��@�1
�S�f���y� �<��T�
���Xƀ��yB�I~���iQ�E�5*,�����y�I�L��a���M6?�(iB.�=�y�.ؓM:P�@�kе"�n�b��y����N3((y���xas��y��N3tbҼ�R�K�U�p0�r���y�l�*t/Z8â��U�X �Q,	��y��W��0���C�p���j��y�3��k�*�)Ffb#�"۽�y�y�Z��#j�(?����Eч�y�g PZ.�JQ'�4\�EP5�"�yB��5>�д	�� K�lYe���y��̼oW���G��r9Yf	!�y�J�/���x�ᛑ���0�/�y����� �� �O��\��ECU�y
� ]3b%��8�����5�v@i3"O&�2�|��T��#80�Zuq�"O���'��Rt�ܙ#�9	�"O|�8�a�	���SvT
Y�P��"Odф�̜[��}�v��&]4���"O�	�T"��3;���!�e�4"O��  6z�@��/W;���"O�4�w��1���)�
��I�@���"ODe0�D�%wJ%k hլ}U��J�"Ox1C1'�Hx\�,Ǿ]��  �"OhD w�P U�G*U�����"OL$�r�ڛZ����*�-e���R"O:|�փ�� XrqK��_���ò"O萋���9��0r��B2P��g"O��� ��6;@<���=0��aQ"O°�2M��y��(AH�
D+��"O�� $a�>�A�M��t�"O4�2&�� T�帱ł*c�-zV"OL`�͏� �J����ؓ@�K�"O^li�c�Bi��T=���q�IP!�Ͻxa�l�!I��[�2x�����'K��2Έ7L�`�c'1�pa�	�'���ˇm�aw�	�Ӂö)�n��	�'Ӏ9! 1{��ic�;^�n���'B���̀,y�a�%b@"\#��1�'���cbR������
�-u�0:�'ּĢQ)��:~ �F�s��0��'�(@�[�K���@E��l<b�[�'��I��ʻF�&�R�E�!Y��`�'K\Li��cc@��'
�~�x���'�!�����h�bk>n���'4���N�d�M��LXnN�B�'�@P�G15�n�X3)>Tk<�k
�'ɘl�R�߈A7��(�%TANAP	�'�$e���z�(���̓RE0i
�'4�e�T��o��|@P���"(�K�'�<�@1��t����i�� ܚ���'�B��\,vf5[P�%�dB�'����#�S-O>��D/�<�#�'[��B���f���鲈f�P��	�'���F���c�9O�g7���	�'2���R&ޚ/>�&XPn"M	�'��� Ńk�9A��B��Ȩ	�'*8p����'�$�)�,����q	�'�PA үO (w�����y���)�'Qh-��ˑ&D�œ��*h����'�����3^ ޅ٢��;��R�'��D�O&ne��I������j�'m��`�IS
,Q*��S��+2��
�'�.��@�:U��$S�$ʄ�V��'�*hт#�+yz��ѱ͈*+�N�j�')�M�G��0���Q���Bu�	�'\&�v.�:^���"���B���'+���ӌ���)� '��|��'�NI U�,q2���L(x�p�'�N�e�Ϟm�Z�㴢 �%~�aI�'ZZᘒc�.̀P-�-�:��'��It�F>	>�b���9��ɹ�'a��*�£f�JT���&^�
�'�
�;��Կ81���Ņ�:5�ؑ��"ftURv�LI$p���3��фȓ%K��2@�UG.�y��Z�]���v��ܲ�J� ~��C�χKH����s��J !wI$V����S�? ��w���c�F�q&�rg`X0"O8%��Ոp�0�*	�k^���"O������ ��)L�P�ʱ"O6K�M�'n���ƞ�
v ��"O.��GN�Du�QD�;=D͹B"OjLi�R�� a�D�=$�#3"OpA��
U��hr�
1�!P'"O&�G"P("�\��c���"�t�"O��SA"�0=�����ȭ	����"O-ѦV>�x�6��$wbjS"O`�anKY��HևaQ���"Of�:rgݚN�Mk�G�'*-:�"Ox��ApbY ���*a�JQa"O���Uh[�rr�q��m���a"O�X� .J�Tn�a)�닗Z���E"OV�K�a��`S&uz�+V�I;���"O�Q#2~����%�s0B�"O�yڗJ����U2��K�~����u"Oj���*1i��p�g��S�(�f"O����|����ʈF�ΰ"�"O]DȒ�#ՠt��-�$	K�"O��9���+� ��o+�Ne2�"O�e�S k��4��E�xY"O�`9�I�+� ���
\�!g���R"O�Eҷ��54��@�v⎹��"O�x�kW�[~0�x�f�T�4S�"O�UƸR:,���P��Ӷ"ON�y�"�*���2b��O� �p'"O0xi  с,�p��`!�H �%"O|رt,[�{@b��NQ�v�$\�`"O�u���'nk̩�Q��t3U�%"O�p�cϗ���%��8b�@�"Oi���#��8*G
$��#"O��F�'p����V����Ex�<ٲ���p]@��̠e���1mPv�<)��&!Q	�Ub�,,�A3�#r�<�SO�
���sᢜ@���' �s�<Y�]ߖ}�wm��F�:�@���B�<�d:#V�a�
�;��:v��z�<ᕮ]16�p��
�=ؙ��L�c�<i�E�8{İC#�Ѯ���V$C�<a@��h��u��ŗ�z�2䛦`�R�<!���a7\�Ɂ�̭
o��v�]J�<���@�����! ��,;:����G�<Q �1,�zY���>t���p��d�<ٰ�ѻE:2(b��X"pa�o\�<��b�Dl��W!h�l��I�u�<�@IK���pKC�K�	�L9A�z�<�`��B:>��X2PU�x�t̗u�<A �Sp�T((o^�*��x���o�<yc�ΕW���c�2W$`�!��d�<�!Á�l|T)��-g.�i���k�<9� DF74La�^�x��$i%D�C�<I�� >f1>��f�h>��C�~�<	��6	��)�dރh�N�z�,HB�<ၫ�,=��{6�Ŗy���
�JK�<�:�0�d��=�J�p,�K�<�so�$Y�Py���=EN��F��z�<����+�2����ĽP\�h���x�<�Dۮ��c*ݻ-���w�M�<Y�P�(vF�"�A0M�͉��BH�<��_>�,���N��?��I��U\�<q��-^�%8w��5s���B�LD�<I�&��ud� 2`�]S�lJ�lYY�<� �*�I_&�x���勢6xV\R�"O�=�r��8XOB�$yI �3"OX�� E��.�}r�f:Lt�"OR��KY�Bh�C�P�"���"O��Z�&U�aN�`����#%����"OLp�M��op,�JPL�k�Y�e"O�{�o���I5�E��}"�"O,{��K�0銬
tm�Yp��F"O�PM�}j�諕lG�i� "O���D�i�xYe\a�6Q�"O���,��8���9��X�XC"O��zA�]�>�B�O�V\�4@C"O|Q����9�X�zR̒A6D��"O�\)���'q��e�����$"O~-�s-ݮi4"p"�&�!�,ȣ�"O.M:)�'f|.�h�f�$�J;"O8y�qI�	�ZȒ&�Ou�63�"O��Y��	��a�����&��L��"O�5�a�^����&�ϕCy�l�"O�]���B�k:tAB��7:�%k�"O�H1�� ��сeO}���P"O�[��$�x��'�(Za2��b"O���e��Q!j0&J.|��8�v"O�(��gV�F:��0q7Zd�0W"O��#A��H![���,�����"O�ݠa�Йm�
�C�����9�"O�uQ�BA�E+�� �̌*L��=K�"O�hb I/b�"<��B�=p��t"OpٓP�t��x�ʎbV�	#U"O��fS*cI�U0�)ߌT�4��"OBu+\�M���Ɲ��hX�"O���AܓX�P��̀:`bPS"O.ȩ����Q�(��$��.Q�d("O,�QPa\*���A&"�:|�%�C"O��IC
��L�h���(��� �"Oy���r���Р3���C�"O�d�G��U�x#��f��IV"O��*�-��7d�A#CY-!����"Oz��s@L�7����㑖�A
�"O�H� �N�H��D&b��c��U"O��"���FL�Dڱ��y3��y�"O��G�n�����C�tBT4�5"O,Ӏ�)���cS�ƈ{7��"OX�[��A`��#@@5,�!z�'�M�N�n�	�/]=��H�'�
���[yiP<Q��T:eg�\�'i�,� �.|�,=�F�h��P�
�'�2}ie�[�/����H X��lB
�'�����H�4RX�(a��B}�Ȳ�'�`�r� �F�Vek�_5O����G(  Lqt��5!5�i��@��~�
�i�앺6����M�O��(;�.�
r�R�X���
*��9H>Q	�|�ۆ�H3R��	bEl�w�X�ȓB�8
'��0�� ��Th�P�ȓLL���ĺA���)R�U`��ȓ�h|2RlWz[P��ǚ}�8��ȓ=`��y�s���@���=��Ob�}nZ5`��QA��ґ^}Dxh��G�^���'�Q�XF�$�R�a��jR�F�a�$,0�b��?1�)�S�O!�٨�N�?:�PX��M��#���c�8ʓ�0|"#�6J0 `آ�+3�� �h�O���iExJ?b#V�&rB���؞c.J��'�%�$1=�^�b?����٭vɴ�X�U�;M�{sdE�(Ϟ�b�'�x�a��O�й1�2�q���"(|�+ �m��jŰiPܤS��OoJ�R���/K��1)0M[/BV������
t>� ���a,O}T�l���G���	2�$T��(O�'lX!a)�8F�<���#FT'�8��)�5:�>��Я8p��,� �&L��J�£<�����K�L�BƐ�S3�Lk��D%_G2�x����'��݁��K�n	@PaՌi��
�'�j�����2]����H�*�l	��'�N,�䄜�90^Tp�JҖ(b��C�'�֬c�ؕPfR%��c�-I�i�
��O�iN��?pHZl��D|��e�'�����-_"�@��J����O��(�OP �Mk�� 	2�ޑ'�T*���&�71��i1r	9��
r �(�y� q���RW`L
�|�Q"�'�y2@ݑ/�.Ȉ3eJ�g��"���y��I`�1�dҤwe,H�؃�y�,�O��iH�H���
�'E��yRN�+; j�ʐ�"l��[b��+�yҬξ
�8��(֐TN�x��y�' J�D�IA�	�()�G��>�yb��]����y�,��0�K��y�EO<""��h�m�*0��%��yRƛ�n�p!��-�E"�T��y�틊#?X��c��!h�}���Ɂ�y���n�����(�� ^�&,k	�'F�dqE��D$�(Aȍ\L���	�'�j��`[�5�����R�X�j	���B!�( v��u���!��L$D� Z5`N1���@�n�	�TE���"D�x�I]:u��i��� � m�3�%D�Pz�'����؃#�nL<0�F/D�肂L@P\a�aڐ$Y"FG*D�l�Ӌ	�k=ܤ���X�j���N:D���6���D��H�%JKq�A�b*D��v���!�����}����'D��2g���%)F�겭�2u-�- k0D��h2�=D��"��N'��;U� D���aE�u.x`��'�M�v�	"=D������js�B +Δ	P�R�5D��zb�������N�-g�يi)D�`�5���r�P�Sc!T�x���B��%D���rF�D�hp�Q��%`hʨkg�%D��+�*�$1���[㪋�Pa�M3�#D�$*U�H0C�MA �\��և"D���֡�!n�USP�F�6�<m�`(,D�\Ё�H�E(@�H5�85*�g)D��se,ƫ5�V�y�d+83�(��#D�D��cY7���tg��W�����!D�l� f�y�J%Q7LF�gV�����=D��Kda��~�P�Z��+c�5{�/D�� U)�5��J5���r�I��2D� a�J:_��%�b3��/D�L�������ѷ+ �12�-D�Ȣ�k�:
 �l�)i�ѐ7'D���@ш�H���B���Z��&D�H8�L�.'&��0�
��R�����%D�4�p���XfXAh2N����J%D���"ѳEE���懈�a���7B%D��Bsi �x���h��$S�ذ�DG"D�p��
�	nޝ���ƶ
� ��!D�����`2���)O!F��"'�?D���A-�?����Uj�f�U85�>D��C�ڔG�j5���?=4MsPb9D�������M�x@hB��R�R�c�<D���3�M��d1W�˰Y�S&�<D��OA�9�9����̻��-D�� ꠰ �Y�C$�M	�j^:^��Y�"Oh0#c�(�@)r@�׋x鼱��"Oڜ9$L�*]N�,�,JԈ%8�"O�����TA��Y���/�M��"O 1�X�{�Z���"�,�U"O��XfO8u%Yb7��y���	"O��Ҫ�c�>(�1E�}�"�S"O�y[Հ�=*����d�=i�,�{�"O��q�M�T��8���~��(S4"O4���(�v?�|Kr,K$zV��b"O.���I�1� �w��$|b��"O��H�J��v�
ԭiO����"O��b�J�@�6jH+H�0�"Oh�zf�P�H`��j%E�YV ��"O�0����t��36��nA]�3"O��O*}j��Q�,3��q"O���'�еB�Ij�A��Q:"OX��`别U"ꬂ�^>s�H@ڣ"O�-J�j0H���@�l�m����"OR`)��)9�nm�lP5�p�QQ"ORDB�H��T2�� �}L��"Oxd��N_#�|���X�IwĐ"O$=k���%���⅃�?w�"Ov�뇡	�?���DP'9�R�Pu"O�@;E�؉hJmߊJ:A��"O���c
�3m�D�5Żh��"O@��� 7�C0��! 8X�a"O��� ű=�:8r�(���""OjH�OźZ*�U�@nк$"OX�y�K۠%�U��J�J�< )�"O$h�F��7K���Ԙ4t(H:�"O�r����.eK� �(Z�4�"O�t ����l�Hui�)�3�|(a�"O��;A��<!��2�H�L�ҥaP*O�M�b�&ĸ�x"ǃ_�HH�	�']���c���2$�(Y�C����	�'z6]b�΍:��ݸd(x����J�<QԄۿ3�"�h�C_�~ �t@R��E�<�L]27�2̡c ���E�s�@�<����sF�4���L Z�X'j�<�u�N��	�T�I�&ɋ ��w�<�e��;�B��$�]X뢅w�<��.�D���Ta1L�;���q�<� ��Qf]� �N7:Qv d%�b�<����A����3	 �PF��Bb�[�<����q+:���ET}��pY�<���׮4�F��fN�0~�{��SU�<�eH6U�­c��U?j�N0��)N�<Yм�\I��� 7��� .O�Q3RB�I>��U2�JN�P!��&K�z*B�	M{��j1�R>0� �"�R��C�	"K�V�Z�ƃ&��#��R��C�I! *��"L��F�~Px�0^%�C�ɂnrґj�&]#��D9&�C��)�tMS�kߎN%p0���Y�)��B�	?/�@����2��7�� n�XB�	4ظ���/$a����!;�B�I��ș��&,��@�O� Y�B�I_�B-�#�X$5��5hK+�B�	0U��u\*2�x�a�J�%jϞB�	!W$^��Wd�S�Zu�Sf�#prB�0'e�9R�F7Z2���E�K�hB�I(������H��p�2�%D|6B䉥_w:e���+�<��rE@�%��C�)� |@��C�#�,�2���^�`��"O�9sQj�^�)[t���| #�"O��*�,�0d�x����C�h�"O�!i2ջ���"Ӎ]�� ��"O����j�v�����,V�.��z "O����.�8c���#v��$���
q"O�Pg�R
g��ᢂ.�����,�y���s���Hc(J�ln!�#���y"��}ܜau@"b���C'C
�yB	��x ��҆� X_�XC�M6�y�&�8�Qy�.N*&�`+1E$�y"Đ�^_v�$�X)
�@:1N��y�D��g(�旰	�℘�kݾ�y��-d`	���̣4��5�T�
�y2NTw���*D��)��m	���y��Sr�T[�n�Oj�}[�3�y�Jџ$��iH�HG0�Q2��ݖ�yL��x!2�"ǔB�|E��N��y�o.P�zR�O7�慘�NS��yBI�����Js#��(o
�0�5�y��G�'�@y#�S
`N�i ���yb��7:aPGC\(�ٲw���y"N�2�pu"V&Q�C$�S��N��y��ܷngdp�`�TJY[fN���ybo�Z)�I��-�V�3�?�yb‼� ҥ]�$�@����P��y���wj��#T͛l<��d�)�y�B	4�
ͳhG��Z���y�̟��� p�(»��S&Ʌ��yB��"95�4`��I լZ�f	��Py��G) .H@tk�,�Z-�p�x�<��SZ�0�Ec�(�P5�3H�q�<�%�0��d���M� J�l��Xn�<�u���i����J5<R��j�<����d��=*"B�;1�:nҢ�y��H|������A��x��O+�y��=���#�Ц}���K�ȍ��yB��@i�aQ��)gx
p��n��y20a�~1ѯ�!Z�&ȢE��7�y���j|I�G�	��]8��
�y���}d(C�m�y�@Ti�
[��y�I�.�����*ϼby3Bl	��y��$c�ԝ���k�~�"��S>�yR��u�P�Zw���cv͉�y���+�@V
W��<Xs�S��y��5�x)9���i���׋�yd�>�h�Huk�6��m�ҩА�y�K�*��E���M�2��1
r��yb.ȵ�|qʰa	s�������yb�A�_��D��n�%b<���y� ��Yv"�A$.p힭��!�y��N�H��Cԛh���'�;�ybA�/l,�����U�2�JUgͳ�y�Lܪ2a<p�r�^�NV�}��b� �y�H�i;Ҏ�\(���t��)�yr��t�B���Q2" �DT*�y҂��]�n�b�oZ\���ش�y�a��N��`�WOCM�9��k��yrlǰ
����ᢌ{B�q��D��yBJt��q�͖+	�F��R��y���޺�;�@��<���휕�y�nC!i����ɍ3-��4��-0�yr&�
������˭Q�4������yªġr��E	%쇯\I���,��y
� �d�E�B<u�zHY�`�240*պS"O��� ��):�	�W�
/���R�"O.e""��@2�)JU+�)5����"OV(zafW���㑪�W�~��"O�P���&"̈́��4KӝAH 8��"O^��ъ��J�H�酽]:��n"O����	W��*@�֏u����"O̱ہ�� KPF� ~F��"O��+�ֲ>j���eX#hR$�"Ow.ܭ"D4K�C�|8"h�"O� `h�z���1�_�J1h��"O(�Q�>c�Ts�Ϙ-q$�{�"O�uٰ�q�p-� oժL��ؠ"O�9��f�8�(���Ɔ4�Ȕ�'"Om�5c�/g\q�ɱ+��*R �O��b1���M�O?�
*�T��F�7��	S���W�¨��lLnlh	���W@��Y�	����T)V� E���Ͽ���)N�i�U�5��(�ئQ1��,]� �ʅc֏7Crp �ѝd�4����Ƽ��/�6>�ৌ�g��X	�i�%���?A&\���-���2���(�'�2��Z0m�����f��HO`qA��	l�X-[B��0A��[��	:�M�i$�'��Ա�R�X �	�u�*18�5.���s�+EyR�R�Jʨ6�>,O���䅯s[�q�.�����8b��gGر�U��>2��"��?���m��O�-�V�#�j�(W�7Ya*���Q��� 41��ȢGE�~�B�3ƠYP4�8���$	�4��ĵ3���5o�Uc��ɤ.@`�	�[��̃3V?˓���>�ċCz| �VLX]�.�{C+�U�<Bm�.,�!�ׁW�+���x�!+B6���5$��S�?}�'��+�lg�d��$_�p�� a�$()�Lq�'�ɹM8�P���,�^E�Eb4<�h�x�2�B`�ct�P"��*�M#��QF�'.�����S�&�������x�$�C�uk���E�py����I�%T��YT`FWܓ+}����1(��iwj��y�~)%�|c��Q�G��ē�?)����'{�S�>SZ9�!(�瞭�� �*2.�B�	�S��qV�� �9I7�^�oh��I	�Ms�i��	�P[���ٴ�?�����HV��ə1��!R��lTވD��؟\��ٟ��wK��q�	�
 >k��$�̂�f�J�S�+��NRB��J�H�)��-]#��<A�$W�^=Ĉ�W*x DPV��ot݀��7$z��#�߾Z�m�f(�Mj���B
7�"=�.O<��v�'466�fܧn�\I��O���c��S�c�:�����O�c�Ȳ��������&/܎�iԍ.�OB-oZ��M��4/ʌ�!a�����
��^Z�^��AZ�ԼiPT���dP֥ӆ�TC���H#
�YA:�@��_$�5���0v�)Vb�^9�����	�����C'F�)2�!\^5�B
�M;��ȕe�2����69�ݰA/��]���5��ͬf���eOB-@)���aܹ�M�������4A�z��?�G��4a����ѫ�0#@�e��@�%����?�ӓ�~ۖq�l�!D!V�'�U�ǅD�(O��l��M�I>)���u��� G��&�	u*`Hp�,GX*"���O�9bCX�Z�X�D�O@�d�O\h���?Q�4(�B��<�^�q�'��n�.$�rD� �vb���$��%�L")�T�[���0I>I�)�pJh�2��%G��D
�������C*� |
VJ,|(�2�.���Ȉa�<W�pĪ�$���;�.D�|��@5Z����o}Rl��?	��i�DO��$�O��=F}x �/`7=���V�_��F~���	��H�A�P���X2�ޒQ��`W�i�06�%�$�`��-���2�D �  ��   F  '  �  �   t+  �6  �@  K  �U  Y`  �i  Hr  }  �  b�   �  ��  ϡ  �  U�  ��  غ  �  _�  ��  ��  *�  m�  ��  ��  z�  6�  �  �  � � 2" �( o/ �5 �; x=  Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�� |d��"O
`�(�;���8���-0��1%"Oj4��ND^[��"3/9�0|H�"OB���H��*�ʞRy=a"O�味V�!X��!&F�:J�$���"O,��a
���C�Ą�M�"O,$3%o�-���p���+Ն�:1"O��ݢ1����`���y14]2��i�<�6��{_���c�H�`�fX�$Kn�<��A̼VI�xR[�)�Ć�pඤ�ȓA5��('nߡ4�� �)˩%� ���,��r�؊b#`T�eT09���ȓ!�b��g��}�8�F��-? �ȓ
K|m�ș�VṔ���2�%�ȓ"R�X�j�4JN�1�˘X�i����̹	_�jZ��1!g��zܶ��ȓgil,*�J�
j�Ne��i�J%b���f	�(U��:���G��$Y^م�~r�� S�%T"���k\�jx�ȓ|4�1�îJb��@ӵ�ݩn�V��/[`�"�v4�R�!ʎ<��M�ȓ`:��z�ؚh�J�Z��$HY:	��H��p�m�C1��!��B:��0��EnjZA V;9����J[
2���	��4'J�EA�IVW&��~�(aZ��ӹ�>� o�Y�|�ȓ�f�A�
Ο7�H��M�$�����mޠP����/���ANXo*�ȓTv�����{ ��-7�*h��I��sB�8�8���3����ȓNe*M�悡;������X�o��!�ȓ'lj�#F�m�+R&;�|��2)n�C��0S4���T:
b���:�0!��e֊��)��ͷV��,�ȓ0�&�8#���� ع�L�����;�P�AFd���,w�6d���hO�>a�IH�8<��ǫS�<��d�,D�����#��qAv�E<fBu:��<��'��{�ʍ-7�(\"��0O��b�'��0>a�47z��l�Wg��9@��Z4d��Ȱ}���hO�>�3�L
�@�9RH��k�d]��=D�$�׭77TTjbL��gؠAѷ� }��'<����˅;b���!�*��qw��!�#Ќ�y�9���O%B�	�3U��s�H0i��	�"ON c ���J*��rc'ʈ�^Րf�JH<���P6W�舂��|��`[��Es����'�2�I�:��l� d�#�|tj7���yRF ~��#QŐ2J��C'߈O��r����|�"۲�	�&Ae.�l��p=لL�72��[#L�m� ��N�<1R�O,�L<���D|�@�EʭS��˷��G�>"�((D�к@�]��JCJ�zqB¯L�@O@�`D{"�B&B�~(��CDsy�w��5�yK�%�����ҙ �EW����y�)]�~�$���j�{C"$��c��?�ڴ��'�?��f��]��UB�Y�_��0;��j�<��N	7pAb���D��H\��%�OМ+@.� ֆ��g�ݒx���@"O�p@� N;z��T[j萃�"O��cA��q]>]㇃��XR��{0"OFՙ��
Y�b��x!��:��Iix�����8nfE�O��GE,D�� �)UĊ+7���9рH�"�.��&"O���l.k�6� ���cɨ�t"O������F�ވ����n!(* �'!��	�j�c@�W�Z����G��{"�S�v��/G-<��)N�F��~�V��xNހp",ڂGۙP�]�q�7D��4��b�ph�FԢj��S�K6D�����F��6}k��Ֆ1y*-j�o2D��[��=��=��W�H,�D�>����~��|�Aa[ &Y
��p���{���(�P�!n�U��<�����b�����?lO�➈
���Yox�x�DM5�,$��D1�O�牵��낡	+F���8F����Q�=��'l�>�ɄU�U��N�:+,������B�I9�� �ʐ�"� Y���(I:B�I'9z��÷I�ޠ��A��X��B�1_�T�iԂ0�܀*�"�j�B�0@CxT#�FӔx8��X����ad��O��H���<�	R������!6� �^2oz�B�z7qss�ɶr}���늅sm>8��hO?�YW狻w�PC&� D�(���cx�XDx��͏cd�Qv�Ǎk��-JG�ݏ��$(�OVI�DmQ�����Q�P�X������$�Ş3^*�b�"Q�{���F(�[nB��ȓz��Q��W����u H����ȓ �ʝ �-qnYǫ[�]�<4�ȓKT&-QEK�9a-�x"�fK��P��&T���f\�l^~ɋ�h�&
���ȓt $n�jP
;�j2�p܅�	 �����0�d0W���{dV��8�T! ���]�`@�E�*�,��IR}bi��PP̥х �$u����#�(�ybƂ��BRG͉���Ѩ�)�hO�G��D�).��y�n�;
�����f�<���Xz�L�`	&T�",Z[�<�.�&��P�>]Q�u	�h�o�<��F'�P(�!&W=#>,,�B��u�<�'Md��zP"C�6���rx�t�'zX�����Ī���<��'�ڔ�瑠��3��P
�
D���'2�I��d��P�[�O��c�O��dC�N���F�4i�ř�F8��OZ�=�'�M+׬U6*Y�]��畺<l,B�(��b�Im��|
)X�9�X��F�I=P����%��y�~�⟬"צ�c�J|Il����Q�(D�03�DQ�[����Dڮf��S4"�<I�ODc��GxB θU:5 ���9`�^u��.�hO�"�
־p|0� ��P$�PxKEOL,J�O���&u����R�;��p�֋!Y�lm�R�$�>E���8�*�c�H��Z��-�bN'+��=��t�*ec�+� �D�G�ь�?�yB�dtn�l9��G1�ɰR��&G��}rR�4y��Շs��)5fQ1;O��1��G����hO1�\� $��I�����ƨn	��'�0c���gռ_������i����E7��Z��0Xc'G�MШ�B3$_
v֐;fl�O��=E��C�[�>�b���,raLR ��O���܄t��HB��?)��)���ϑu���r���i��Emg|����ÞTr((`9D�0s�oV=;A�\) �H��RE�;��L���%��!�'�H�R����0�[���ȇ�MF����?6e�#ԫʄ,F{��'�bYe�WjhP`Fز7G���
�'�0m�T�1>�Gc�)(�FTB
��� ���k�::���SW�޼JF���"OƄ�̓]y��{Q���uCx��"O҅(pF���SD�%6+��Z�"O(�E.��>DR����ڱ1���"Oʸ8`�Ι0b�}�U�7g*<�f"O�4�?�N�ծ�
 ��8bd"O�(�ƨۙ�B��d�0+ ݹU"O��:�!K(@a����!=�6ث0O��WgJ���֡.kp�13��V�
��IQ�I��rٚuF10f���2�n�ʓ�hOQ>ɸw�X!�t���(I�9=����'��hO�Ӹ�Ra�f��cJ�;�F �DB�	�-�H�x��T:Q�D!ÊOB�	��v��3�5],}jWD�25��C�(-N`�%�U_E��^<"���^�'#�����#���p���xČ��p�!����R����}��*��.!�DBd�r@���֐��i( y!�_0;��G���jz4��C�ni�OD�=��R��K-+�n
O�t<C$
OF6̬�b= �EF�J9�1���I�r�1O0����9fi\�K�SѮzFG̋u8�xB����A >v�#��/?�$A�%�#D��B F|�Cė,)ž)%� \Ob�X�o@8a2qa¨S�s��b��=D�,A&�6>W~d�!	�*NV�Q�Fl<D��;E)�4�Z��RM�`����pm�<q���S8�*��@/R	q�V�k�烂t7JB�ɿ~6NDqq��X��h6������?a��'%�h��ȱ{����eۍJ�٫�'����+�@Q(�=� ���*�y���@�z����W�7���#Q'��y¨�B2"EcWX�$��W�F�y�́�+؉��k[eyΑ[@B��y�B5C�`"�IXVҚ�����6�y��̍2d�4t�W�yx���D^<�y"�͊oRzM� "{�l�*Sc��y2�SLt��.r^R�C"J�y��,�(u�V��.j�^���iF��y�G^�>`�����t��7�yG�s��E׊�6�P����Z��y���8��[��.\Hai��y�dM�ƽ�uhI�Y@��h!�yB@9M(��4F����F1�y2�G>Y�D2��R��d��I���y2#ڡiA4�fiҨv���X��H��y��\o��Xb5X�0�Q�A
��y�ӰE�xy4a��)�GE7q�!�X{���QȊ� �n��"��e�!��T�`rDFرh�- ��ʪ�!��V���ےCR+3�,%��G$�!�g�h̊7��:{r��1�A�=!��P�2�<qS��M��t�.�$�!�d׷C+I����:M��̖�+�!�ȥ}��Ÿg �.
0�!����!���E��A��D�K�P�蔩΍t!�d�2j�Jux�B��B��i���"O$]+�L�	;9@�Q��Y��1�v�)D�P��̵"��L���t����**D� �����a%���r��s!<D�����?	
}CGҁ�t#��,D�d �?@���h�kPT�X�d�)D�8�eO͈��y�EM�)�z��r(D�ȫ�#ڟf|�� ĨI/&G�0{�K&D�� �,��`������9$��$�`"Or����՝E�x��D!�*x5��"O����P^N�ipoT�73��+�"OZ�1FGӿ@Ph��Q��/21�e` "O\59Cb�!^$�ja&ȅ���'"��'�R�'<��'j"�'kR�'Ep����~��3��d��'=Z���'���'��'B2�'B��J�uhv���'@�O ���*�e��'��'�b�'z��'��'k"&�*�`��$��.{t�x%CF@��'h��'Z��'���'�'UR+@x�f-���4S����AF�z���'9"�'.B�'��'�R�'��LSc� *�N��h8� 6<�R�'���'<��'���'�B�'��I9���(W��; ����4W�2�'L�'!��'�b�'=2��ߴ|,>�3B�C��4q�U��(9�ʨ���?��?����?����?Y��?!�40�����Sk���j�W^�!���?����?Y��?y���?!��?��B�����"�5��Ly��;F%��k��?���?I��?I���?���?9�1nNx���#��I0�"�V��q��?���?A��?���?����?I��Ģ5�Al�� H6*�&v�����?)��?	���?q��?���?���R�6�`�gX�J7dY#G��#��@����?A���?��?����?�R�i�B�'�B��D�Ue4p��l�<y����<�ش�j��慘�9����2��i�A�Y~r�o����&�4���|��g�>8_ ��Ќh��!ST����ɗp�:?��b �tC<��#\���]�g��<j����'�Y��G����*,\*4
.���d��
�N7��1O��?=������ɝe�f����V
��)Bc�N�}�r�i��Ķ<%?i�i�:Zw�扱`�^H��OJ�-�(�@Or �I�Z/���2က=� E{�O��J�`�̝�G�;yRt!����yRX�L%����42w���<����^���A�A-1BQqa�:��'����?)ߴ�yRT�(c �&U�Z тF� *i��T�5?٢W)7�@(pɖş�	0����?A7�=���^jQL��]���$�<��S��y��}����!̾,_�e�'/�+�yR�s�X�A�����4������.%�����sE|u��V��~b�'���'�A�����d��FVźc��;\������<lH�NU��T�v.V�E;�(b� N2����Q	H�奬ЧiL�Q$�Y��(HE�߿g�R��&�"2@�ijdN�[Q�CV�ٗ^%&cq�зd� D��F�1zn��򤍯U
z�A2DD�t�������K���e ��#SfL�GNӘ%4�XT
(Z*8xYs��9g�L}�S�_��0��c]5�N[bgV��-��D�k�.�R"jZ�� ��eP�[6lP//��e��bzӸ��GF��^E�����.="Iq�'	�Y ��!a�q[Q�Jh����T��'#B�'A��>�;*��Ԉ��^�Y��= �޷-�x���O��Ĝ�>d��Uyb�O��'�T����C�h��2�,m�#m��I�ٴ�?���?��'u<�	by"!�G1l�LP
�8��ֈ'�7-��z��D*�D&��ǟ�q ˟�e�T��S��$�h�r�� 0�M����?A�(�!���i���'A�'(Zw7�� �M��|�aKݯ/����4�?q(Ov�[@=O������	�ѠmӞ��5��]�F^켹�	Ɵ�M���x!ܙ��in��'z�'��'�~��X�[�)���<�������dW�$�O����O`�d�|���4�.�s���"���&���~�9�#:K����'l��'�bȷ~�,O��^ ��I�'��/�����`+
h�s?O��$�Oj�zGm�O����|��-��v�6O�v����JR%�lE ��\q�7m�OH���O"��O8ʓ�?ɣ��|�0���'6�4�e��P�b"�(U֛��'}� �͟h���0��>G6a�ܴ�?��#6�RḖ�y�rD
$oS�����W�-�	��L��`y��'��O���'�� �ǎR�C�q¢�_��q���2�'-��'2�����U�IɟX���?�f�)��Z�a��.�b|x"�I2�M�������O*8k�1����O��j;��!^�!�Jd���CoA����Ȓ�Mc��?a��47\�&�'D�'0�d�O"kH<!Dt8�g�=Z�j��C_���?��/H��?�����4�z�O�
�A��1�V\S���y$u��4,10�i�R�'�"�O����'��'��T�щŦg=��&!�;">���qHx��}�Ռ�O,�O�'���Of��,�&A� Mc�ǅ{��8��d礪�����	�^����4�?q��?)���?�;_�d!�s�̯H���s�Bl~=l쟘�'�R�������O����Of!0��ː_<0(!�
�.̲]jp�B��]�	�B@���4�?��?)�p���G?9Q��^�<���I�V�����b�P}Rό�yB�'jR�'u"�'���KJmcs�M�J.�$���6>��e	�iՈ�M����?���?��V?�'9�[�zN4�m�>2��1�^�P�'���'IĔ�7�'>��'��.{�X6M��5��ʟ(\L��S��]F^�mzÛv�'6R�'��P���� y�^�Sybh��H�6ĜL��B�Xc����O��D�O����O6��H!@�AlZ����Ʉi:��0�퀫 �h3EH
Z$j��޴�?����?�,O��S�
w�i�O���Ol�h��K��z��!	� �0?h7��O�$�O��1f�um�����0�/`(�H�,Q5G�Nt�e�Tx����4�?Q)O�䞅0��	�O���|n:� V�[BGdT��PE̗�t��x�i���'n� 7d}�p�D�O��d��v�)�Oh�S��3u)����힢{B��'�h}��'qDH[`�'o��'��5�Of�X�
	�b�Nr,�׷*G8en�%�\D��4�?���?��Lt�'�"JP8��������bŜs�86-��~��"|:�lB��t�1.�г�&M�u(5���i���'��*��a>On���O<�I:e��i���@��9�B�V��c��9��?�	����	�0"��҇r�60H�*�V�׫��M��\}^�t�x��'8�|ZcKU
 �\Tإ�!,�l���٫O�9s���O��d�O�ʓP�d�z�O�y����2b��)m��qE�	�S��'P��'��'Q�ɥ;ڤ����B�t��Uz/���JX�G1�	ԟ���ş��'Bm[�~>��惇�.@PakT*�;c�Z`BK�>���?1L>*O���!R�`��OW�89��t�RI0o�>����?������%>��
F�z_���=O
�Y%/Ԍ�M��������LN�O�����	���B�'�Fl���i;��'?剠8��sL|r���ѨY/RX�QS���\�stD�2Q�'-�%H\#<�O���a¦6
EKuǑJ���4��dX�L6:)lڧ��	�O���JB~2O޸=� ��b��`OD�x碅�M/O��H��)�S�V(\L@��0�t�{��.K�d6M��6�Qo���`���8�S����?qࢇ��\X2��5lY�!�MZ-����4�O>M��zԥ�'Lԍ9���A��N�MK��?��@�~�뷗xb�'��O�i�dZ [�4iZO�v��P��$��az1O����OH�$[�	>�t�����M��}�l��^�ll�ԟ�sR���'ab�|Zc+��q��ݺT��h�� =�:l�O襻f�D�O����OZʓV��q��}���2n�M�\Z�$���O��$�d�<A��4�����h��s�����:F���<���?�����R�y8:�'^[,��1. ]n��zgeC9R��'jr�';�U���'M�}������CB�H3��.b����S�d�	˟���`y2�З� ��x+ ,� Y�(݊��

4	"�ͦ��	ퟐ�'0�	����g}��R�=�42a2O�Ib%�,�M���?�+O�I��)	M�埴�S��
qI�IB�#q\�B܉K�F�޴��ĥ<�W%�e��O�iuNm�� �
tݫ�j��-��5��4��Wh�`mڥ��I�O����V~2$\��BB�^�T0������Mk(O0໠�1�i>O�P��X�@�f�ޡ]����i!b�Z�c���D�O����Px$� �I�T�ε�VG@�Ii�c�!�R@�zشo�, Dx����O�E�O%P��kQ��Qȴ<`S�������������KV\�N<���?��'{���:.���V�� hM���}b��̘'|b�'����D���Fs��;c
+�6M�Opi��`�p�	����f�i���
 A�\����� ��>٥@L��?����?,O
1cƯ��?�4��O�s�Ĺ�P1Y�JT%���I��$���'k�œ���c{��ö�I�]���;"B��'�b�'��W�x+)����Thʷ^�(d��+U����Qm����O^��)�$�<іv}�K�?C̮����|R! �����O�D�O��1�>h������е$�i��1I�i��⁻��6m�OP�O �����>�!D[�d��1���ʪ U�@�Jۦi���P�'$�a"�)���O��I_O�6��6�Qr|�����ӸIݶ�'�0�'Y����T?1��B8N�8���aU�KL�ӆ�}�2˓53Fdb��i���?��'x��� T0:��%h�*����BQ�7-�<QkGe���O��À�$�ttQ���	|)P(y�4x��(
܂��?9��?!��$I�'KBJ�P���2Ѧ	H
т�
A0p�L7M]x<�"|���j�Py2VK��¬y�M�	�6�逹i���'�r�98�6c���I}?�c�8U�ْg&ĸ��A�N�a�Ϯ��<���?��a�����(����Fڶ��!Q�i��!~��b�`�Ij�i�a;j��Q�؀�ȘH<�҆ũ>i�{��?a���?�)O(���/��ɴP�'L�q���V��'���ߟ�&��'�};��H=]��:Q��.��9������'�r�'��]�pi!OS���de�`�����[��6�7��$�O���#��<� � p}���/q̐�"ɑY7�(�˳����O�$�O��h��y�����*�)�R1-$�c`b�#�7-�O��O �a��A�>1��J1p��-���]Rn�嚗���E���'&���8���OZ��N�a}������&���T'I-�'��'T��`��T?����:(<����N/r�2I���uӾ˓���령ij\만?���j���	7��1�!�M�-�uw��6�7M�<��}���O��)�sh�#[ۊA�̙�?�Qrشn����S�i@r�'���O�lO*�$M`y>!a&S4_�>�����(R�Hn��!��"<E���'��� ,��C�7j��t.�i8���׸i42�'�b�_8O:���O0�I
'2��	1D�!�\��A��>3Zb�� 7�,����	ߟ̨�&ٰ	l�Q�k��:PK� �6�M��U�t�x"�'��|ZcFP`4oF�z�@��O�a~|�OP����O����O>� f���L@�E��u,��H��N�n \jN<���?�����O���¢Bdl�6�P�9�9�wf��k8x���O����O˓`�ؠB?�8�{�B��;�z�8���<t$��]����ٟ���My2�'g��	����� �D����@�z�Hz�E�jw��ܟ���ßP�'$�	��./�	H;3eԔ��BJ;C������H�l��IPyR�'
��[���Y����A�eP�HV��$�t�A��d� ���O�˓=�x�`I~������ Ɨq`@���;�P��L"Z��'#�ɱF���?�O*iȗ.��̴��O��4��ڴ��T�@��l�/����O��)�J~�K�B>uk)��SԦ����M���?�3Ή��?�H>�~ra��`j$m�#�J�S*�צ%q�C��M���?����ꀙx��'l�����$�� ������X��l������6�)�'�?!� ��wS�r�T<e�5pE�X0����?y���?QW*�3F�'��'����3=j���g̕
eܠ��ޛf�|��)!	�� ���O,��@�j�z��pA�2-ġ[��X�=���m�ϟ�y�a�����?�����ӡ�%YWI8�l� )�-�pb@W}BgO��yr_���I̟$��}y��ĝO��iVe�9�����KE!�-�p)��O���4���O����K�\����ͧ�I��HW�eߎy+V?O���?���?a+O�	`�E�|dl0Dm+��| ��n�p}�'(�|�')��
$Z��O� a3b<�z���"��r�O����Oj��<�t�",�O���#�ŝp؜�"¨��8t�z�&�$9���O$�$��7��1}bn��Ia ���D�r�z0��M{��?�+O����d�S�����I�����جz�M�ri�%}�0�M<����?���[��?�M>�O^��EI�	�r$�kp%+ݴ��d�`��oڠ��)�ON���~BO֯DX�[�
г ��%1�*��M���?�0K��<y+O�>�!�K]�r~�:��S5H�rW�y�Υ������	�P���?���}�K��z^Mzc�=-c$���mC�#f7��+���,� �ɟ�x'R�X$�8 `b
�A��	�UE��M+���?q�#�����x��''��Od�"�o�'@P ���0E߀�	2�i��'F���1d4�i�O����OJ�3�	�"��� Q�2��/���ɑ1�
�QJ<	��?	K>���� �L&I�P�ࠅÃP�2e�'�-�'�Iڟ���ٟd�'J�\aVd��vŘ���<{6M�	녕xB�'�Қ|R�'���@(�< �k�>'��V��{�v�[��'���4�IE�S�L���O� M{�NE g\��xFN]'jN\��O���O�O���O�y���O�=:%$�� hH7�R�P��ѩ�P}2� k�za+�֑t�bX��B�
e��7o�ld@I�'��>x A��I< �"�ОE}�5{ƌ�9:��SEX>*��0f�C�E��C)�HOL,���0
���B헌q��9��O�A0�Fi�t����")�0�T�WPqFʅ�B�ȘBP��WA�<��a+~4&��  gS�%8�%˦gu���圌����V�))j�uf�BL���a�S;>E�S ��K�0(�V'R�~Z���p��L\�� (��`�K�C�55d�y�Π�ʌ����I�xC�';��'�z�b5e#J1b\+���#}U��)୍7l:����ʽ&�n�����0���'��ϿKt���@J�CD��n#wr�%:�K��L��"�$sE$�K$gR�)�*�(1m�L���ið�A9tivq���e��є�����Iܟh�䧵�v�Zi��O�F�h̡K� ����ȓD���Ɵ0J4��I+��d���Gxb�+�S��΄�hI��p���5�t:rȓ��B�'f���ү�!���')b�'��]���I"=>L�D����e�%�ܜ+�h�� 1�ɉo�^�X��?�=��
�Ԍ�Ge�($7��Yջ����G��!:w�*��1���Y��*]%*'���c� ?��=k' tj'I�5\��%����S?A�S����ۓL�>�Y�oV�7�{R�	|w>U��f�B �r�&�j%`̂5��٘��i>Q%��P戅4�M+���Xw Ƞ�ǧ5����!�2�?1���?��.��1#���?I�O�xP��;Li���ҍ.2�zc�� D|~jg�$��}�B�'/����̬8��eXq��q���@,OfVN @�aݖ#�<xG�9�:��U��y2��=AbNǟ�:�43�!��\�e��Da�B j) ľi �O$�G��'j��C���od�zщ[�*��e��'�ȱ�a��1��a'�){Hٱ�'y6��OPʓfn$��i��'D哶��Bq�J�HD�2TSv\��������	�X5c�hx́srI��ta��z!\�D2�I�U�?>��@��y�w�U�,V�<񐣂&>�V��Cmζ7�4��4�Z80(�p�Lp��̫�&�/�Y#�k�I��<��mN՟xD���٧N�Dmz���(RH$ Ĭ���y�C��L�Α�& ��~����3�0>)אx
� �l�4BI�nA;�M�}���@"4O����dR�����ϟ@�Os2��e�'v��'���R��*0�ȁ!pE��z麄�A*B6C�{��&2v��tH�O�`�矴��#-I �\i�Kˤ~�x���&D+ZTzA�D%
�v�Z�{���hO���!W�yV&��Ջx���,(�`A��2{l����+I_������?a��|���'�ވ� ���81ʹx�<�JT�
�'b51���b�%	6�ʌC��d�f���4�'�����܂8��R�BNȄ��'}��K&G�B���'��'�cc�1�i�%��ݺ~l��cE�ʴia�����<qE�"l�,�:U!�p>$Er��,JF0"��%��EY�リK0�ㅁ@�� ���S���@�ߟ��k6�����'�:��ƎX���U����L�L�r��'댁�`�'�Z6����<����d\1&�� �d�	�d�T��aI0�!�D'_Y��@c/��h`Ќ��G �3�ڍEz�,�r^��Z�l��u7��8�T"�9'L�E�m���'Y��'-���'s�3�n�z��'���K
/�i�ӽ"��8���p>��KyrɆ�`24K��mJ���vF��p>�#O�؟���4�tTm|T�[7�ȳ/[0����Ԑ�k'mЌ��&�O8l��`��:Z���g��{����̓R��|2�( � 6��O@�$�|�Ց,�Z��Ȉ��N�Y� �������?Y��MF��:�������@{��A# ��
&�߶(�4	R��[;S��?)�cK z�աrƞȸs
6ʓ�`9��{�O8�*Eh��<�ҡ�K��s��y��'{B���H�: P�SEҷp�4�1�Um�'�fegiՕd��+�
�c�����'W�ҥ	�H���O`�'<0& (���?��ZqNj����$|lY���G�=*r�!e��?A�y*��H@���(L�T�v̔44+H98���G��Gx���'9�	%˛ m�.żG��1�#��P��@!���Of��4a(*�P���R�DՊ�"Oz�W&�i��+ǅّ>}6�#��	��HO��Oȩ��c��f���2@J�(0u�O���^�Vpp��D�O��d�O���Tr��w�uP�A�N�i�Fo�$na�'N��Wn�.��=I4��0e��(��֟><�4a Q?�E�T�|� L��ɭp$��7&��6�\p�"�̴61���8|b2���ɟ���?��?�)Od;c֪vd���{>����"O�]´NIo���� 
�%��Ӆ�Z�'����'u�38Dسܴ1A4 0�	�\V�XS �y��i��?���?�6lǙ�?	��?Y��P�6�0C��?wPЫ�ćNH�AE=D� �']���"L63i�lQ늢�@Hc���	�hq��$)��+s�ʮu@�#?yU���8�ݴl��R�AA ?Ң��� ��T9g�i�bW�\�	t�S�t�^�9��X ��J������y��',: �B���)��yQ�Ɵ�~(��'�� ��Fx��˓˼�E����d�O˧}� �t�R�F��2؆7Q��8��V�?9���?�c�@��?��y*��%�r�ؠAm��pԩ�� U*��4U����)}�>��o]%S^ $�,�m�'�*ؒ�'Ǒ>E��Fı)���Z��6bzD��G'D�L1H���|!�:U�*r�.%�O*T%�t�JNֺD���Mex ���f��xČɃ�M��?i)����F�OR���O4ũ�G�#�&�#2%[q!A{�L�]���D"�|Fx�gW9�j��.R�Q���	!�^�,�)���)��4 �/K�C�M�w�խ+(
|KG�H�q����	e�S��?����=���	��@􆼓��P�<	�j��JG&�(W ���f�T�'o #=�'�?Qã����k	-C44"1N��?��nັ����?��?a��B���O�N�.�z�!1��-RҚ�Y㋶v��DƒwZn*�J�90Z��dڷ3�� �LT<k\<���CR2x�z}��	��^y��Ǎ�^_��ʄݟ��9e,lܓx��Mɗ	P
\eJL ���S�jA�O�R������=�vh�%�N���p+�����n�<ɂ�P�2%+p� �0�@�Ci_S瑞�Sh�	67��ش_RB�Z��ہ4ݢ�H!�8c(�����?1���?��N��?)���T%#�?��
LNu�B��TB�AK4"�p���@�p����n�,S���PLQ!���0Gmh�$�O�i�(�O��H&�Q�W�Θ�0"OҘ�eOމ$(*��t�
.	j�"O �a�ԓAb�	��G�.{ʵ(16O��n�|�I"����4�?I����� �`��?"y�0f��!$	��B�9/X�D�O��DS�* �T�⦊f��f���ŀ",dYa*�">p���o�6�(O���ɛ2L��X�,�[�O�. ��F8Y�p!���X�N��� �� ���'�h7-�O��'c��Z��p���Xu/���ބh���?�M>E��'�V̲PH�1*�dZDOU	g�b���{U��f�����;5�њ����NS�����Z�V��D]+m�4�m���I[��o�+��'$r��A�V��O�.xZ>tB�`͕Pg��y'�'�1O�3�}���"֤X�5ĸ\+7h/qJQ���w	Gx���'yB�3 �,��UV�GD�LB��T!9�0���O���� 8���pԪ��Q&h5��"O|�
1*���V
��?{*	0ቚ�HO���Y�p�"��J����tbR�E_`!����;@�	-�,��	ٟ�	��h�\w��w��:ԉE!P�h�Q�%k,�iR�͝7s�
4b�-��т�E�=���F=ʓG��<���&ʒ��V��;~�̝0'Nc��Թw@�30�D`R�JX����@�=1�L���p��O2�wDǣ(�8����s�.���OUY��'�����Έq��T"RAQ�U�D���N&!�$�4�>��*�v��c�ß1��Fz�O�'��St)j�J]��Hz�D�j��k��]���O����O��Ć'c�^���On��	\�x��iپn�RF*Nm�\`1`��&	d���fT��=��I$e��PՄٱx��%�C�7���DYg�=�!C�!A��@��A��X#��$wG�➰�E��O�n�!Zl� �G��Z���b!���pB�	�I;�3�`O��n���J?�^B䉢2�z��4��#K���xvj�	,�'�MsL>1b���Co�F�'2R>q�d��%�H!��S��DH!�Ԯ�<d�	֟��I 7ݒ};`�	$@^� 7���`�x�9Rݟ|m{��H����H6&<�pC��6ȴm��ƀ:-Rh� ��^n̋@M�,@�8z�V�z���;�hA8p8����K��y��&������O��F�Ɓ_.�0�0�X?9�"���+�"�y҄L̐���A�/d�I�&B�6���"��|ڄ�x�B�jI�1Ic郏�V�06�,�yR���<6M�Oj���|Rc-���?I���?���#L�nBJ�+�0-�R��)ff����4S�n��bU�e4��T>%�|�I�"JBx���#K��%SX�"�P������um@�9��V+R1>��Q��þ{��Ͽ�3j��e
m;u영2h�y�%ş:��x�������2�6>�����&�R2\a33,ͬ�y"�Dk?J��N�P��8q'���O:(Dz�OCr��!Pp����4D�x +���0���' p;��pm��'{B�'�zٟ֝��)t� �c!�� �Lz"�� F�I�ίS��0� �cnX��1�(O
T�w��a3n 4b�6[�>E17�@K��%Q���C*�9�E��@��)I�/S�{r�_�B�j�z���we$Y���T�� ��(� ��	�=y)M<U�ҝkX�lPwjԾ=2m����?�"�>Bm¸�&m�
Vpt�s�-AR����Sa�)cl۴SeBD�jǯAnb�HdgKK\�1��?����?Q#(
��?!�����~@6 ����H�҂��wJ�|�wFv������
LT\z��	�&P�UdB't�\!G���Z���85�C1=l�TB�DTۦNӦ����I���B��O@�lZ�:B��zGE?K�H�ve܁@��B�I�K]L��W�C�^=�I�2M�C䉴 ��H� A1$pDm�Řk���I�M#N>qc`��9����'0bW>!y���P0�;�,H��*�J1�-#$v�������*7,�A��A�S�tΏM���+� ���`�¨�(O�0K3���@@ 7�B2m��P�e�<:?�<��ÁӟG���� 4�9x���f��*� �y����
K���Ə:p��ӥdʲ�0>y��x���-gdT	G���x����yB��;j�6��O��d�|�W�Y��?1���?��"��`/.�BW/
?��p�sg��an\�)�b#C���b�?�yUT?��|��3@�
)�bߵ��(a��sN<;(�KL��r-)(>B�g�+�u��O��b�Ū|�6x`�qq%�ρY�4��t"?h�za�G�֟@�M>E���{X�R@�B8K�H�e���� ��64x��鑂n�j��1^�*42%Fx�j9��|���? L�d/�3`� �3��W7k�y���?��=CR��y���?����?ѳ����4�*FM������#)�@1��B�(��آ�B���<�Q�zi��aڟ�"=a��>k���ӄOb~�e��7��h�V(�&F�,x���J�j��y���M��B�UH��'��H�DS�i�B&�Q��r�'� ����a{�N3T�(��B�K���xӇR�y�K�$-D21��L	�D(T|I�e˄BJ"=ͧ��~ZP��iy�rFӌi@��s�FW:7N��'}�'���~sr�'q�!�"��� $|���8�ec�-X�x��'Sj�X)O
�J������0\�<��3"�'���j��?Q���Tߠ��M�k�3��~�<i�D��UM��@��� �*� �e�<Qd���r��揕u�F�b����<���ix�'-�Ț�Le���d�Ot˧?�Z��GI�,G*�1�>�~��A��?!���?1PZ��?��y*�6`��5�[5T���� ���J�Q45�����G�/�4}@�IH�'�|�h��h�B<�qa_�% ����عs7Xl��"O�k�
	����"�6z-\p��'�JOl(iE�ӪYZ�X��J����}��;O�����զ%�	��4�O�>1B��'�b�':����X�B��@��J��}�5A�58�ʷ��IdV��k�O�w��43`*E�)��GNΒ	;y��_� Ɋ4��M�Z�<��AE�uy6��#�6����d) ��;s�8�S�Y�E�u�NT�/fd"A�#�?�Ԟ|���'R$��-:k|�9SM�y����'�PM!6��#J6Y�%��/ ܼA���_d���$�',�X`��A�~�c)�l1���'A�e�Dt"����'&�'N�{��iީ
6�i���"�*�>�FY҇`�9P},qهI�0b��Р��8Kd&�S��(O�y��%ڜ
�`�"!MBY<�����l��f�`�!�L]��Ɇҟh1� �:Ir����>!�MA:X%1�*˘{�6����q?�*�ȟ,Z� ^�E�v/Z=5�l ���
)w� Ć�s\���`j�A��Ђ�^%#�u�0�i>Y$����ѿ�M{2��5���F��t��ى��'�?����?����tl*��?ٜO� iH��ɦ_����[�ZRF�kg��#.�x)��B�|da�V�'_
��%L4K$�1�� �MnJ��F�xa��C%7oJ���`��6�F��5Ŷ@8�{ך�?���s�Z�/��~�
�ä��?v�����B�aT+Q`��ӂ�g6����lL�x�J88v2D�$�$O����Û�|"kȻ2.�7m�O���|:�Q�KF*T�Q���!~�dە`��?��?��cG�o	@��r�K3Qv0��������?tA��C�ڧ:/�)�d�0�Q�tx�j�?Fa|a ◾*[�ʂc���
֝�S^�YAă6���
�'�N��f�F�H�N]�	��H�~��aD���
���Xc/!��"O�$ц"r��Ԣ�g��H*���t�',�O$@�7!�Q����dä'V,H�7O~m�!���E��̟D�O��9Z�'!"�''8�����6BF�X"K�oV�dpc�dl�
p��5�L��e� 6^� ����ϿC��1R���C�@�ju�3�[.�v���;���#�O.:���h�ᓱ`x�!k�y������'�����H0m�"��������'���O?�D��@UPK�;�"���K$?!�
Xo��[��шFv�d!2	2=�1O����M�����'LN����zcD�B"��j�T���'��щ7�����'F��'���y�]�i�ٳ�䍙o�P�{��G�iz1"k�hN<�'���G��D��'�	#�4���(O�y�@LҢu�\��	>�j�E!��<�r����B�>�k��@{���!.��R�h�4�d��8)�EV� �J#�
���X�.�2��հ=Y�ŃH�ܐ� 6� ��ի�K<�Z&�<"��ߝi��ɄI��=��%ّ��Si�`�:�4W���f��'@�B��� [�!2�x���?��?����?������V�m�l`!��רs��I	b��f;�A���%F7ePeM��PF�y���>t7��Y&ꞇpBz�r�
�v���R3C�����w��<��15GD��q�G$�'@L����n%�� �Z?
���+Y��`S!ڭ�y� Ǆ7�����ܝE"��	�G2�yb�M67�d�!���C���Js�I �yҥi���O�{S'Ӧ��	��\�O�p�0���9(��� ��(P�,� ��;"�'��~e�Pe��WN��ʀ @:�'A��q^��b���[9N��FyB��:s�h��49˺���!N���	1p�o�^�t�$S��@qH^~�qOF�8d�'��#}�F���Ax�8yƨ�#Xh����+	I�<�BeK��lya0��	��� �*��'�ēT�6�;&`��Cg 8�B�%-b̓No���d�i_��'���W�y�	ԟ$��>.i&����"L��Ό*O5,�{䍉f���(������:��i"���HU��
B�h]
��`�Vb\�����K����G] aH�h &d�l;H��;1ޢ��g R_��w|A�3��G!�p�.qq8ѩ2!�:���!���O��OX��tG�F��"OT1æ��q�F��4 M=5GB�
 ��HO�i�O��3�j��s�	p�o�|7V4�A��O����=d�q1 C�O��d�O�DN��Ӽ�UM�2fDs��βД] m���(%�q�K/5�4��bK]�:�ވ���HO� >��fGǤ>θ�A�Mĸ�X�3#NڃYt�� JC�r��R+#���z�p�1��I���I%��w��4����������Y���m؞��3F�iؼ�(���?3A��*�e*D�z�@���j�c��ك���HO�	7���=<�<9oڅU� i��*�O�>1��n�JK�i������	� 3�D�ş<�I�|R�(�+'��iV�Y��n�2�ٷ9�T̨��ҳ5��@Y��B4�Rͺ�����s�|"�A2-p�h�udע\x�ZnN��($�ŞJ��{�$���\��qOX�s�'�X6�u�*9Z�*U�:
(x(u�_�w�J�l�g�X+�>���ҥ�A�Ň [��
�#N9�0C�ɈY�P��kB�tȥ�C�KJT��:�MC���D	�z	�-�O<RV>	�6�ܳJ�����o�9��LRc%�7 3��	˟0�ɠ5��b�eX�y�jA¹i�PG �?�)�f�>Q�~�;�C2[�2�RS�&ʓ��`HB`%b����i�"���FP	% 
�*1:l�dL�w!<i��M�pߪ�2p�|�-4�?� �i��c?)b��	
2L�����*D�	s��j���Ixx��� jڒU�<��Μ!5v���K.?���4��T&�����R)f��5�U���@�q�!�v�PR�F_��M���?+�b5Q�/�O���O�����x̦��7],8�@J,x�&��ĮW3
���zff9�&`��mЅO��c>�.H�@�rE:��Ψ¦@z��I)���r��[�T�0[ Ɇ>�V̙���w���Cu��w�	��hN�2*`I�!��oER)���H�������2��$%C
i��F��/���6F��y��V�L��uvf�R.�O�O�Fz�O�Iםk�z����>#:}���\���'`Z��
8[;R�'��'8�̟�]�����a�7Vt��(�%?�3M�}�=+r��,/�ȣp'�?U�sm<1O�=!�kN�	$�9A@�Լ)��LS�b�4���߉j�U��e+v��I$���!�y���{�<pYӎ��lケ�D_�~�˚�?��'�rt����O
���:P�(�'�v� �'� �\;���[-d8p5�(��|�K>!v��z����P�i�(�E�� �dyA�L�H�2�'JR�'M\	��')�2��� �Z��U(c�@L��@3�J�r�&�Ӑ'Z�C	���U)�(	�p�?�F�N�h	N���������p�ΑJ�]0�K��<��=�cO<< �ȏ�$/*�'��\��
��@�~��%(_�d�y��'yL(���Q��lT(R�&�="�'� 9�	�:vp8���F�!�t4��'gN7-.�d�n���n�ޟx�	{�$��I�h�q�
l� H�@��I��5�!�'}��'�����(,`蠃!?>bz�T>MӤҡ#�s�� �>r��%�.�y=4��D�=�1zG��L>��&ǃ�}�EY�a�;'��㷈�P�x9�s��|Jt�<�3��Ο�D��,X>U+����k��CT\ൌ���y2	R[piP��u���2f��0>i�x��.4����aB�E�Q�ۇ�y�&��1y�6-�O|�$�|�d��1�?y��?��p`����"_���RI ��Q�@	/� �cmY�Q�^6]>I�|�	�"�8�+�,M���*E��x��2ӄL�C�<P�E�D�B��ʂ�G� O�(I����y��t�g�۳Y�<�:5D�&k������I'�?Qq�|���'��T�󂕽��yq$��,@��'�dzw���Ȍ@���o��hq��dEd�����'������	}�lY����p��aB�'���@�P�
%*w�'���'Yb�i�q�iޑ�Bn��D�L�[c�
�q�` ��n,UH	�5���kڼ3h���s�'�L����]�R���8�m�%Ls�Ԑ�.٠Uʈ��5��q�\k�����JT�IB����3��65=~يg�%����#X�SZ*��=a����~؞lP�d�7U�0#��]Z4�H�G<D����*�敐+��LS��Ȏ7ي�Ez�O��',
FJrӬ����;0���dk�'@L����O��$�O6�DK����$�O�S�wn|��Kց+h�����u���DU,�z���(���+�F�<a�]��#Ot�'{,�Z����
Vg͓F�.	���pJ�U[���/R�g�ҭT�4�Ѯl&b��X���OzTl0�Z`e [BAi�
�2JZ>C�	�A����)N"k��YbHב_LC�	^�@(X0  ?o��x�z}�H�'��7�?�1��o������_���h�x�a�!Ƈ�9�e��9]�4͡6�'R�'�T!��O�Z�8�s&�+7;|"����AH�$�E�֋m�~Q��i�'/�M#df��{ 0���Z_��Q�U�X1il���� �����"Z-hԱVM�n��=��
�՟8;ٴI��V�'�哀(Z�@E�+�@8;��N�zþ���E��?)��?.O��Z�m}\92�-��m����tc#��II���4)e�6!o��$���F�#6ti�N�%='�l٣�}���a)H�$t���l�O�����'���'r Ȩ��;a��0ه�� 7�J])$�J�l���T>#<i4��w9<�a ���B@�p��F�DY����O� �ta��X�!�#NIg)0��d���dn�)��l�E��	A�<�+C��7U�(�&D�T��:� �r�l8<f�08��%yX���������$
�����7(��
C�p���h��T H��������I��u���y7d^�;�)Ǩ��?8�����>9C�K!�ŝD�؍�qE���H��OC2$BW��W�/O�6hL��X@`��X�J~�#�^����*��ANȑ��y"ƠȘc^`b��s�KйԶ��$E_�Q�bpRF�������O���D�4�p5"V���x=���B �!�$�Ƥ "��X"%x��ハZ�,mEz�OS�'�v ��tӞLQ7�Ġ[̪��#���J"�l����O��d�OZ��4@�����O�S}N�I����TL����i�#ȨYJa��#?�:��e
4�O�E�G�7C�
�M�3c�$�	�Aǭ}�D��������zE��i�P{���C�'����2���-��/��U�$�Q2@#�� #�۴�yb!4t|��s�e���j�0�yrσu>8`"g�T��#V��y�|�ƓO����R����	̟̕O��ab����)������dƉ#M��'�b�-f,93b��6d�<(���/g�'�������`f4����uraEy"�.�Z=���Wʴ`u�Θ#�Nɽ`\$ Y���	F135��%�5{��L��qO�-�%6O\"}�c*� �(1+�/H�-9���n�<��k�	J.6,��ɑ�6w��K�͟C�HBL<�D�1��X�����[K��{�O��<��!M�vX���'2]>5�4j����� �VM�	AQ@W�U������/H�t��������I�$J��є�	��Z��թ$��pP"DC�����/.K���!O�bę8�AOj�|�R��'�֓O?�#��R#/��Sp���Pc!�$E�:��I҆䗳f�,"��E��<j���?E)� E�ZE\,x�ŝ��1��ǟ����+KN)X��N؟l�IƟH��=�u���y�a�+�V�Ғ��4t�m�a�]�~��Vllib���ay�$��b����m�|����˻K8R��#I��Pd�%1}|$��O�ԣ<Yt%�Z&�\�Р�'d,!�Hi?	���ş��I�29�`�%�x����X��M�"Ol|K5"@"bk�6̜l,�l"�(H������aJ���Yh��/WҠ��׈"� `4��ş���͟��	�"� p�i�n��|f�t�Ixy�P����y�X	�(��H����ƻ2��	++���c#�=���`�͟���d6>��j� �KW��k�Ԕ떡�M*���"ONe�f^0u��ABP �5C8m��"O�����3�L|� E׆cd]I�8O$�>��矆���'�"_>)���*�H�%-GF��ѡ�/6���8�IƟ��S"����<�O�<bS��-G6fU�bB�nMyَ�X�[��?šjN�J	���h�#Mk����	$l���e�Okab	�+R�Ԉq���m�4���'Wh�H�#THH^�hc�?9z�P�<G�'Ij�եH�R�f�����=��s�'�.Q�If����O�ʧ>�Ȁ��?I�	�6�ćj/DQ{�ȟ�/��� �^;�?��y*��H4��wd�Ց�gؑa��Hf���c|��Ex���'s`��Y�9�*R��v���2�K���2���O ��L �d��j�1Ӓ�"O,A	3ló:��l#a�4"��q�ቊ�HO��7<@EcW�̦7�
I����',�J@�I����0���5l�������˟8�Yw��w�<�����$v��� ��+ܑ"�'/�5�.K�7a����ݦ_�`$�@�[�I�0�0ǒ�1��$��z����'�B��akC�k5ڥcVjId��(���P����O�eo����?�����9��%��Mbt�v��!�DW[Y�GKhx�z�m��GzbX>��'g�L�6
gӊ��'A�1F8�08�%	{[�ԋƉ�Or���O2�����d�O��ӘL7����O��1�]�-��t�Q�
�fgt��%�'sD-�*O$k4CT!K�9+֤8V�m���'g�Xy���?)�f��PF~�Cr�l�F*Kc�<y��)=�0�v˗�B���@�M_�<��B�#bq�|8��Z�^�q����<���$C45�D<n럼�If���Y I�4b�%�
!�����]ݒU1 �')��'���'S1O�S�eH�i)�"ۚ x��E[� N�<�fYX�O���/�&�>����g�`�����:��/�g�? �!��A�$)�!;W����a�p"O�91�G��� 6�� R�
��'��O�t�s!�Q�\Iv�!o�g?O,@�D��զ�I�$�O�<�u�'���'Dҙ�n�`��1��	�,�M)G�U��� Wm�g�\��#DҔH5
�'ݘϿ�@�@IѲt�"@=p��/�6��d��F��@����ʧ{��������&�5�� "���E�M�%XoY�@�D.�)���yG�ҭ,3���@D�=
*uca D�D����@��P��b�yl$q�s�+Q����'<�X�ᄂ�Og�lK%.�l�$h��?��
ݴ$*�����?����?�5���4��C���M�ԕM�?o���v�Ob�k��'a�aёq�@��R� �p��'�P<��M/��8b��~�F���
�������p��ɨ԰=1�b�L��'��g]���@�K�<�Be���a�!*�=gD�F�I.V���"~Γ	�|�{Ą�"*�1�Fa�(h��E��-j�̉Ɗ �c2���tm��pv	�ȓa *���oҪX�İ�DN�����?�H#!W8UWT`��o	)�H$�ȓGl`�r�ִ�D����CiI�A��zIb�����<	橪���訇ȓ&y��&�D��4N�̌�ȓD:l%g������H
ft��PY^9�Цʮg` �ȕ���E���}���r���'�pY��k���\��s'��(_^�e�DH3(�q��jfvѸ� ��m�LY)�kF1H���ȓ_��cG�7VP A#n�,h����<Д�����?(�viҩ�m�Ն�}��u��i�+hrU�gJ[<�Ji�ȓ�@�tK�!X�F���l�0Y����՚ѮP�D]NIS�h�.fr���[����[5]�Y򐬀+.���k$He��r;n4� @�);�]��&赙�GP�S�l��K�?ˮl��1q��bf�Ç�>)'�[5la��I�\M�a��>�-)����%H!��o2�����'l~��2.���p ��b�َ*o���aC!�y��W��Y�q'Lszr��q��Ok�����mZ�O�F-�Tѩ_b58���Cx����-գR4��ٱ!ӘK�	�ȓS&᠃��`�b�Q�

�H3��ȓa�)a��T>K�*%��ȺΞ���p�~5hb�۠&�,p����<P
j\�����Z����qUA�����r�<X��p�B�3�D�4czM;�ɻuD�FR�2}R��1��:do�3�F��F!�	h�x��+�2�\ٹ����{�T�2�R�SPN�0R%'擀S�8�x��
r�A�!"_��`�P�T��� �/Qy�<� CЉ=d�}j�lÏbZ��pN�`�6�K�\�6J6��$�>Og�2e��Dh�DF��O$���C�99*�R��˛f��Y�O}�$x���B/Ÿ���$ަ� �
1D�eZ$DÁiL{��ltЍP�@UZ�MR\�u��$>��?m��x�2�ЅO̵ �"��S��)>w��O�Dh����O���S�O� ��5@�$`[:~�Z�<�$  ��u�A� 8�r-s��ؒ�*��
T�@A��d�H���:9�8i��O�$[DEK��D��t��w���$J2��}��cԜ���/G�m"�O��(ý+����&�5�N��ר�	2㟔ƺ��\�s��?t��CqBϞ��䋾 ��rC��0.��]�/�:4����wD��}���'��X`d���i mT�tc2ɑ��%��]3���ERF$J3.�<�0<)�F����bn�\�n)� ��)Ǒ@�C+��~�J@2�ވր��.W�5(�jP=p�fZ��O�][RdĀ�HB���)��5"⬛=>"ac��� |<<�r��C34���8��	�\���ِ�����D�����nS�Zs%�7{�Y��#:�ɺk��؉��\��q�E�N�i���	F�n�;��9�MR�!��`S c��ǿWd�%A����`a�<5^&(�W���S@�:z�`�cH�.��)薧�x�4��S�����h�� ��:w�Њ�TP�e��
O��MT)ڌ3��E@'���@&�4��<�����ж"X�X��� ,۴۔�ג>	�IHV���J<���RS��3�^�<1��ƼI.���Oӊ�1�掬c<3��֜�?�L	��IPB�
%Mn��XV.�_�"���Ex�O�����TE�6�k�&W;x4(��@46��u9����H�G����c(����"<��?,���1@��/�B�)���0�ь�V�c���A�<}��^!l_@˓����Ve?A��\҄傲�pMIԆϙ/�6�Ey��)��¢�!#D)�~8:�j�g1"$�9r´ �Fᗃs.��s+6��?��%��?���@C��S䦠+�I1A!��xChZ����.�x�a �0����3�&��?X���B.�z�i�<aC*�L���)3	Ɇ\��'�{؟|`ÎD0^4��aƤ�=4*�=�/Z"0G�]`�O�S�剆8Q�;6�;���	�ҬI��0F�.��gO��@��"?��n]g�0�s��;���z�\���HM�?Yl�k¯9L�����Ui}b�d"ړ8:&�p��$u4XK��B2k^e��O�!���J�/��Xq�"#�8�&�J`m�`����.�CQ�	�So�`y��#O��'��}��c �v>pq3d�|=Cb��g�'�ak��q��QC�����A�/	���ǢW�x�훵-�=�'n��ؒ�$~�c����Dhi�.T�!ʇ��ⷕ�|A�:H�<�Y�g�H�"��!�:�韄���[$4.�e�.C��P��JH[�2(h�zYw�<}���՗l5�d꒛>!&K��Lƭ0��UR�� a��+"2ĩ��l�*��=�=�g�=(Q�s�Hc��}X�I[2�\A�Ջ�}'��3Bͧu�$!�%�Ӽ�Q�J�
�+�eM h�� ��)[^�ۺ@PP��?])*Β�,l2��{�|�Kp۵R!Q�,{4��c� �3×�D���.���@�d%���
��vI��C��@� ��AܓB��	�0n��ץ�;���ul��1� �*�T~���b�!JE
i`���d�������C�3v��9��;�vɡ�%�/Z�qO�Q��g݉r�&�cg��xC��N�dN+����=bnn̫�D�:OA�p���0��!��ԟ�Oa���8�Q���Y�pA��S�K �?���1%i5;��4	lըO�N�J� �y���)E3I��lP3A3�
f-Dy�'���L��$����T%Rv�J�0�U�t�4�"���$AE%���
'�A���	a�,y*DX��瞷w ��J��y��xyꝍ$�>�	e��`�!��`��a	��@u?6(�'@����ˡNj~mRFKq�bxٍ���PbR�g��d��⠇�[�O��u��1!ĥr��B�ȹ���>ybȞ
%x۵�A/m�J]��Ô�g�H�Tꑗ���
�AL��th� .x	�C�q��]��Q�vq	�W�P�ԝ���5�7w"�3��F�����嫚��~�'U�Ɋd|���D H-�9�1�ėB�����	�`������<R�
 �"	?!_�}q���9cʲ�R��X�zY֠;��d�<�rB̓#��d[��ķ1�\����K(@b�&J��Y��d��c/�D�*o3���R�>r�p�S ]�IU}2�Gx�H��g������[��~]�(8�eE�|}��j4i[�̀2(&���	N,�����	U�TC�CѾ7͙p���5������d�'���ȶ�-:Z�T{�%��J����d"��,�.٠ߴ*����U!#Ok��(� ��#X�OI�����(z(��0�Ox��;0봨��ˈq��q��L�!�  Ǔo��D�v�-���綌�鑞uPL�P�'��p ���:�m���`�[%&æ?ʂ\0�iF�0H�ɢ3�xb�ìz���=�~�A�0Hj\��CM�~�lT�WB\^}�j�?:�:��=E�������3�,W9�z��qO<��_�g�ɀF����M�{�<��A
���Odz���4�p<YbHK"1֤pV���W�ν �,��(h�%gE:�O���;a�z��͓3?��u*�k*�z�
����5
7�)%�`	��c=s��ՁA!N� a�cgf³A#>�cV���s��`�iN�L���?AY��B݁N"��s;�$��C��EБ��iՒ}�# ��Ux�I~}dS�+��0,�C�ޙx�i���~�^��1�H�,ÀmHrm�;^&�D p &���J�z��d/ۛ4���Q/�{5�����v��KG��Iyb�I�;��t��ݤq�t�Ї^�!��E�W ]7M�L7�]'O����i��Z(?|4=[I) ��-������x}�)�{O��P�Bͻ%�sA�\�Pax�疒T��*�g�+jd�����ٝ]t���f�1��yiF
�/�����oM�A#�-�;�%)�+ e4lc��Y8U(Q��ρ��$�0*<R�(ſCgz����-����ۋu��<2"+%+,�L�+-�I�)0b�3!
�WkB{`LF"
�X�'�d�#"�*
�!$dҌ(�썛�Cb�n� �h�1�0>�1"�`���X?[��H&��\�#�&\�����E�$!��>�{�? Xx����Dr�x���(�: �"�>�Fk�U��I<�䑹O]\�{�l�~�.��1N5P��>���ՙGI&���エYcdQ��
��7 �b��³�s����=Y����'9��S�6�.eզo�p�:�Gը^:,1�7�T���=tY`0g��*����E�g�c���޻1O�dP�g9*����F���=�u�!�u7Lj�m cH�C��ӲA� 'W��e"�(G:��P�4%M�rD�TdOF�S�>A��&�|�2F��T�(�dI-$��|b��ڷk�ĸ��@U�R͖�>ͻ ʅ��	�y�V���������O`� %/*�)�S1<⺤!��T}�`[dJU��'�I�Q"�B���PP�P��	zB�=�����T��#��,A*���=�՟Ba��ГI��i;��	F]�5I��ػb��'�Ui��ۑ7�4��7!-g��!�'�<x�=O�4��a�0s�A�8cKZ6nR:r�|�3!ٺ�&D�!&�2�cdY+��Ir�d1�%g������k켵#�G��V`c5�i�2��v���V$r6ݟ��TS����qaҁt.4;6�//�0ju�ˈQ�&�E�R�#�*�D}�w���;5�*Of����H�W�`tR���ssz@��X�D��M�|���O���'��!��H� 	�,au�J�M�U`P%�y�'İ(�e,.Q�Z��!Ε�cX�XS�}M�(c�@K�g��i;�!�������O*�4�'OB��r��5�^��	L1gS��(�t�����8���T��(��D]?eU���]抅!D�7�?�oJ � #�OG�߰��b�F�'Ӫ��	�>��$���Py�S���qt	(}G��[VI�A1:�B��O��:��բ*"��%:�h�48"cI3K_�����.U�âV�X��(�t��@6u�Q����X��؄ M�;`���w�� C�5y���mHPT��O����[�g�ɡs���b��a��1��֦l��8��Zj��f��-!j�0��Ɔ,�6ۅbpN�B�
��.�ru�D@�(Vޚ�(�\?T���P+_�M��+��?5�U ֙>(L�0F��5�j=����
 ��0��O���S��O�V�@�AT&V����u|��j�,���A��!8��c�*SL��Ui&)l���-�u����XKXU�f��
�1�'"�`1����H
`�o� �� �"�63�(����h��	q2k0�(a2��*Jg�X�b�r��s��*-��6�\=+�L��E&5#�V}A�ͅ0�(O�D�Ɩh+TW�T(:�@��G�A�4QX4l��f�UK���-t�~�����?E&� ���ح Q�l3e�[�2����� 2Z��Dy��`Ѱm1a�K�r����p�93T��0d`���J��;��(>�q�E},�0�jО#\��~5p
��DOv�Y�1A��lX�]�G�����I�d���B�x" Ty`��[,�HIH���%H��J�h�8<������/�2=�DfH�$	�O��]w�&��e��(��}���E~򥜦P�b���%K���
a˚
8��hA �=��p�f��0�,��񩄖�����51�Z���3���&�ݬ:'��R˚��8���/"�̨w�'�P="0`�$�4S�ĕ��Z��"�3"C��I0Je�܈���͙P����T=�ң]r{�Kv �#!>�Hw 2��6��쳃&�!��RR(͡��ka儕M�cjS�5�.�1� �z�X�F%!ඕZ��;#� c���'bu,���e!�(sE[)<��	W+	!l���"XI�U�^��`!2� ����!�!�$~�l�������.��k��C��ݍ\��@cqM\�lbc�\�+w�)���$���ʁ���L�IX��5��!S�ThqAJ:G#�������lڎ*m�HH�lL�>��G�t,Q3?��ÈͿ~�
��'Z��D3��.q���c��
<b��(t���'�n�Xt�d�H@ ��V+r8"�d�Ml� @��'i�#M?A��b�	~�����OVV���ώ<?�1�sc�x����_9�V�� �߮|��0��m�̈#�	a��U�W�،7��xڴ91$A1!h��?��.�#ݸ'e�ӳA���ZtO?F!�0AOP� ��8�CIy�E��}��S.��Q!�'&MD�+Ǌ�
P!��[F.��yh. b�LT�2,H�
ڟ%d�٘��@�����(�x����U��pP��%@c:��5��?i��%n��Q 0���ɚF���yv(��ON�)p�@A�N"��'R(��̈"g����'�PP�)K:�5��F26�ƤX	�'�z�G�
�0߄ػÅ�.�����'&DhS�H�h��x0�쑑"@e��'}�Ej��FؐAL��q(D�̒�ֲ���V��
+@�Cd$D��K�D��P&���!�Z�}��@�� D�谴��x�$�K`iZ�?Bl��?D�(@�!Q�(z��e�� [�.Ċ�F1D�i��
-"9��:��R����C0D��iG�� VPdr�	��S��3cN*D�I�I	�$��y$��I�<8��<D�p(T�C8}���qSoS�b�h�:D�k�-�;ΖD�1�*�~y��:D�$b�*Ď#�T�Sb��Fn���7D�8`��N�n��� ��	��C�'7D�� "L���ߎ#@��	㍃�� Xq�"O�$�BJߓI��b�N2S�6��E"O��h�=�2Q �^�/t���"O����iJ>1l����<v�Mq�"Ox��ʓ�&�zh���>䬨z6"O�d��p'
	��.{3���"O�1�t�d�2��$�B)J)hH�"Oi�2�ڙy���&��GLKW"O
�����DҢ ȁ�٢|1����"O
m
Fe�
"�Rh $���4"Oh�E� �1���*$)d����6"O�TѓJ̬G���3���
7��c�"O��E�K�N6�T)�e��*ZY1D"OH1`gTt(L����%:r�"Oݑ �7<h԰A��]	F�u"OB��v�i�j�%D��<� �"Ov�S��:��-�C鑋1�f��"O��A�cQI�h��y�l�Z�"O&��1蔨s�d�wg�'? �)��"O�3��h�����-X5"O�p�dlH�
�t��#��	6�L��"O�iTU�����?$�4t��"OB]#���u%��xch�T�~	��"OB��W�]�<��FX�0�#D"O��5��!Qݘ�UF�8*hk�"Oxq��[�W8h���v?jH@�"O���U�R�C�~|zRc��S3���S"O�)'HZ:�j���Uw�s"O*�`��("�D��p�ԛ��)�"O�-	��#4���ϝ/P�$��6"O�X�e�٦f_�$�Ώ�∢�"O�E:ԃ��+b0�h LȮt�h�r"O��A�Mې6�R0���N�Ղd�4"O�pH�D\�Q�UY��ă:�<��"O�r�hC*jN*1��c
�Y��p"O����>�\)@u�F�e�l�R�"O@��H��峂�T�l����"O^`����;���9♃�6!��"O:����>@��*R%av����"O��֬�
A��|����F��a��"O@��̸T�Vl� �,~�Qd"Oaw���L���b�bY4Bk�8a"OJ�:�eZo��S"���3<8��"OXQ`%m��c�͘�a�V
T�G"O4�#�'�6l(�e�Q@�0L��ժ�"O�5�+�6MN��XV�I�"Of��P��->�z�9�Ñu�hPa"O,,�a�K!���2g��dmA�"O�EI��;1HŚg�� =w*���"O��x�Q���a�eɮTZr��"O��I���s&���f5EU`��"OZ� ��]�'�<�iVg�LL|�z�"O�xc�#�r�8-c�'.!�9�R"O�UYD�D�P�țv�F�x���"OXX���Q�#)]�F`��"O*a���&0��	Z��:�B�I����ቊҊ�0& �9o�֊B��l�\������$/��B�	&z&p`�Ӂ����c�
��'&Q�L1��\�<��B0/�.bX6����*D���������a��K:�!��H%}2O2�S�龟�c�1*2��)��805�,0 �#D��1o��DtK�;
����&D,D��Tǘd��TQ�g;&R	Ҁ�+D�� ��`�B�)~}	վ�"��_����ɾ}���3��X�Z��M�)Qw�B�	T^�xp����e����9Pc�B�U�x�2�V�p�1�h7,��B剖$f�+��ċ{�.��� S  ��A1�OJ��SHμ5��H�h�sH���i1ON�=��O �B�!��p2���-�5��X��"OPIs��7gKd�[��^����XA"O�(�����h�
�y�+�=
���'"O� yv���bT=*gJ�1Q�*\"O�MW��,�.�+W�^�*˾!!f�	mx�,��]W:�|x�B�̄Ѩ�i4$�p� 	0)�w�"�T��է�yR�h�1PS.�<~:`�"B�2�y��*��8�!o�	o�,� ���yR�)�'`7��^����sf�*!^�0Ӈ*O��Y�N 3L�Ԭ�lϔ� !"�' ����EP �s�ț>p��k�'�P�J шhŞ8J��֫4�P�
�'���oZ�`����ɝ{��t8
���~rH�&�p�C��D��QW���y�%n��jc�Z.K�`� VO����O��~B�ˈD����fߝq7�APr`�f�<�cE�G�x�a�gޒu/�@�#Μe�<�c�J�[���!��1}�Ý`��hO�?�ȑ��+��]���}j�ȓk<`���px�S�Λ}��qEx��'/�u8(ގ��zF&ב*�Τ��'~�<R�*W��$�ժJ2.n�=��4�HO^�=��z�6�[bLb��d�\�e�ZC�� *wz*�Q	7�T�[q��n��c�P�6�����Q�cR$��	����C�	�q��2&� !�P�윪L�PC�	�H��@oO�!l8@�}��C�{�Q���T"MG4�97Oِ:QC�I�I(�%갢�v4̚��[�B�I�U��S%��L,��������d"}��\(e0N�G�v�9��͜��'�azk^A�bȊm���)�D˖��O�F��b]Bri����E a��1�yb�~��D��;LV��&��O6���	Ȣ�aR�ًi<H9��C��l��P����ַ;À}ԁ\8:�T��ȓ3M�*��[�h�$hQ7W�6݅ȓv-���� �6[�%ڴ���Ix��ȓ�$���
��xu7X4)�ȓRöP+!l��vDk�C�Ne"���:\|�1��o?��� �ժN�]�ȓ/Q*IA�hC�"y	���.�v����W��A�=V�0eaS�2r?Rɇȓh1�0�G�ݖt�a�U@2'b�4��
���|��h 2�0P9���3^�HÖ��z Ɋ��-LdDU�ȓL�V �W����j���(b����ȓO)�BU�ׂ����"vA����pSn8,h(�sI�L�p��Ô|�G�� ����b�>?�ȓOX�4o��A��f�F��<����	ߔ8
 �k0�
� 8�B��/i�!�ŊO���zN�g�\�J�n��|R�x��I+��$����K霱��k�����)�O�i���N��A���}�鱥�|�'1�A���9p�b0"Q=M8s��yR��TGneKC"	�P�C�y"AY`��W[}Z��S�� B�H�F̵0�-�2�I�$�$+��'�=M"�� �^1'����`R������j��{��d)�IH� l!�ï��B�J�p��O>➌�S�gy!]`��2�k_�y���Уz��IJ���n� �$J�.�(jT�q!��۱e�"C�	+M��5k��s�V} C���j����<a��O�'��=�C��$SXɊR�	Ԧ�D{���i�f\� @�;9�}��@�*zҴt��y��)��0�Z�Bd� �BU�FB�f��C� h��f`X{hP��m��;DB䉻v1�!�G��R�"X�s�$B��)��iĄ"n)�(S���K��?��ē�ħO�fɚ@���0����C2݄A���I�'����l�; %���d��3e����'����N>c;����Ј�������\��Pr�e��h��q��+�!򤔲K�V�i��G�`�V ��!��OF➀��NI*i}nb� �1�!�Dَ:ո�g��)}��,��E�!򄈔B44���U!�lpu��!�
[��`�R�K*��q@W�!��8�.aA`��6�my�!I�!���9X,>l����XL�aD�� #!�d�d0|��KO� Eb$B���\�!��K��� +'K�R^�\Q�Z�ס��yӬ�xaMّ"�Z X� ���V"O�qX�/�,bOnhZ&jނ(�Ѝ��"Od�%���\[�C0IƸ��ij�'�����@V��YP��*#Ό���?D�T� �ϺHn�(�ᒠ5M���@m����ɞ4�l�r���<p�Q�y��d��	�S����.]�h4|f.$&G�c����	�K�
@{���x��h���"ϬC�7Z���{f� L��u@M��>+�C�$g��|��A�s��EsЀݺ"l��c����x��K����"bl�eۨL�'�O��96�G�=����e+�/v�\)�6"O��Xe���vj��'�%�˞!"�!�$
�D���v��?W�|mx�H��!��!�z���R�D��5+t	�P�!����h�W�؆��5���2�!�dޓ@l�x!��Z��Az�ѩh��O��=����p��x����i	���I�"O��r4�õy��X�"���f��"O�c穏�Hw�D�0E��>�<��"O�i�4jǓ2���x���2�(<�5"O��d��>Q��؃�-��,X�"O��3�%K�Z�8���͊�4�J	��"O�u�1��Zt���D9t�hY�@"OƑ�w!��B�nɈ2E�B�`a�"O����kjԥc�Ê�[�d�k�"O4��5삲3��ZQb^8����"O��S��	@L�*U��;���Z�"Of);��G&F�*@���S8g����"ORA:vi�W@�a"Y��洺�"Oĕ9�kQ�:�
�[5ϺP����"O@�1�(�z=�� �AB�q�"O����sɲ���]:00�-��"OZi@g �jSBA�Q;�D��"O
�I)�(-=
���W'j�J�"OԱ���Q:"��W�Y�c 6]��"O��#��� ��WlQ�,�:��"Of� M�H�����-�;P�4u�"O�у�L6n�n�!C�0z�l�z�"O� �8c��B)7����&�>*��x�"OhvF+4�:����׳E#a�"O�����_�X�K��C.$�i�`"O���͂#Ll�Rd�]�k@�P"O��i'��*u��i��Ϗ?��q�t"O �Ni��\2�Ƅ��bx;�"O���4����n�p�$�	���c"O��q@��*_�%r��8i�P��"OB��D,U�oj�A���!vl:���"O�K2FG�c�����H!�6��u"O����ƒ�xlC�bC	g�F%��"O�5B�IN�u|n8�oɉo���s "O����y�5cS��>K����"O�y{�b�w_����&&G�Th�b"Oؕj�!搥"E���z�8�"OHy`�Ɗ���y¶�Q+�n	�e"O�p�2@�.8�(�q�;�`��"O��􎅉!D0����ƀ|�te�c"O �!�@%X��S�&H�G�@U["O��D��Nk�q���N/J�a�"O1!E	�pK�-!��g5v�X"O�XӠj0x��8K���%l^ 2�"O���!���ǐG�h��A&T��
4�,A�� #I�pd���2D���i�6s�v=�+�_K��!�Dei1aq&��3e�}�aFS�!򄇃q���o�8~]�Xc��5�!�dZ�bw��6싁ZL�:!f�1�!�W�4L*�����%�����@�ck!�~[ԤsQ��H�ق�`ě9V!�d
��=j�h֡X�kpM[� A!��e��2 ]���؅-��I,!���4�F9�V(@(QV�Ma!��ֆO�&U4&#P���A�`�5J!�Dϐ8�D<;W�9�܀�ݥ\b!��Y�}	��!��jy����c�!�3K[}�AK;Vd	Ɇ��(-x!��'D_�;D�D)F	�����:!��Il�¡H�Oܪ��w$�v�!��:|�`���g�l}hTcN*�!�d\,p�٤���4��3b��}E!�D�P,L���Ϋ	!<�"�Z5!�d�%4~�x�Uĩ��ٳ��&!���$��}�����M�Q�/el!�ט;��l�w�ɛ8r�R"(ĥN!�$Z*<Q�M�Dc&cq�A���	u�!���;4W:��w��=f��5V.�!�d��w�z]y�J$"6�d���F4�!��=�(�4¯C���!q�!�DB�wX�@���Z0~(���N�!�dY�Q���ҰKܓ ���*�!�d�3[2��W��;QZ�cЏL/v{!��M� ���(���\)�O�5n!�
�-4��f@�s�<\�c��8Q!���O�����.���Q�@�,5!�I1"�<(P�F3%2(���??!�Ė0mDl�����a������T�G.!��y����%F��̃6'
�G�!�r�xm�s�ߨ�`	æeA�t�!�D_;Z�4���̅Ơ8+�%ؖ�!��eL)8	ӓ)��h���'%�!�D��f.�V� ~�`���׿O�!��/l�if�=9�j%	�P)!�̚�IXT�C���`(�5(!�� <����m��۰̗�r�Ɛ1"O���i^�>=t�p���p�	S"O�u¡-J�B��z6�*!�i!f"Oi� /��K��%3R�����"O*��"F"i�H��&kU�Y���r�"O��� $H *����	N�U�h��"Odڧ�L9_�
X!�E�
%Ȳ=:�"O�d`S�@6^"��k��Wt����"O8����o)r���jX)IH�0J�"O����$J�w�eڵj�,��p"O�P�A�׈M�K���D� "Ob�"э��cG$�2�L�R���P"O�X �^ (P�2�A��]�4IH�"O�Q�SJQ�L�c��9�R1�'"O�qJ�MU�����K��ٌ�&"OF��7��c�ڨ�e˘԰1�*O$@���k�!�Df.���"�'�*���/�v)i��\�-�H\��'2nT��;.�<X:ToCzaN���'t� �i2>��D�a�(�'� �c��X[�Q�͆TY&u!
�'u��	WM 5�Q��hZ+U�:��'��xʑ�0�$������Pؾ1�	�' �e���&�  ���7YsL�	�'j�3Q��f�Z�k�<?�p0a	�'��	�e)� Xg)1GBy��'�,(s�4q��!�@�!3:ٱ�')ȉ�e��VQJD3�ΣD���'`��a%L� �|����?�}��'�P�y4n@�p��#B��:�'ih8+��"!@����# �H`
�'-��!�)|E�aj���&rC"r
�'S|�qqJҴdȒPZ��Z�~t����Tl�&ō<\�D00��i��ȓ.8Z�q2	I66Ь�����.,����0m�dá+	nd���V7%X`���w�Ƞ00Z�k�.\S�
������ �0D�����h��=.�9�ȓ[�Xq*QF� 1��4�G�%g����ȓJ��	��ЅL��yʐb
�I�Q���<L��"D�0@����]�v������҃�A�*{S���:�@����^�S���"��xr�
�Q;���D.�x����U���c��Q�(:�	��}u|�!�-!�tl\�AlԆȓ=�|�8e*Ql��Ҁ�PO ݅��*��#�Ih䠓u)�	l#.���x��� �Ə �� �Ӂ:�x|��J��b��B�x#��)�P�	x���WyP%�Vo�TJ��)-=D��{5���d�f��ȋ��(F<���F�xQ���Cp����T%bD���z�tXi����WL.�I��"[eN��ȓK�l�ceKRD�H�!SP{`�ȓi((��V�^�8ʖ�i$�Lތ$�ȓ3A:i��_`3rS@O�G[��ȓ7z�
doW.�8U+"͗-4�ȓ愀Ce���F�n���M��J˔��7QtE���/|ެ�'�{���g�n���F������d[�A�ȓ_S��c��@�*�<�$�̇h6� ��C䜥��*�9� �@#�ż{Z�ȓzz����#JQ�UCɷS�
���d��Y�s$A#k����I����S�? ���SD��P�X-�A�l\�4"O��c���b�����P�F"O*9��G D\ue�E�)rv|�"O*�2��Ҟ$;\�I̋HH��'"Oz��f�'t��.ض(�B��"O���q���1fn䑡M�)%��E��"O�p��(������+@�<��"O�}���X]R���� �"O��+g��%r��:��ɥ�@h�r"O8ȃ`�M�R����q�l�8�"O��r7 Ic��̨$I^��j��"O�]���]\�᳴��2�&�R"O>p�b萢S�F��D</S<���"Or�C����X)[�`D��JV"O�]�ሚ$=*�yU(��T/�� "O���*��{>T���+6MY�"O����lh��e�K�N�1;�"O�yz�E��j�yA�D�Q�T�y�"O�}h��$a�6|���֋H���r"O����� Y�z���Ώ:N����"OzMk��ؑ}-�}��[=���"O&��!��>���ǆʺy���e"O��s��F�0`�cVf�n	�"O �Ď��
�r�G�
��S2"O ���ȓj��pD�����P"Od���OҐ_�q�L�4��Av"Ovas�� �`�pAlN�/�D<��"O��pENiд��b��x?*(��"OƘ�B�ʽ� �D*��yI���"O�y� ET�k�T�#RH��x��"OJQ�Uo�)���R�F)y4"O�!#`F���~A��ƿ��U "O\���-�4�F[��0�Y�"O�C�J� 1!�1����"�h� '"Ox�:#�.��I��D�FAZ��%"O*�`��U�1�����55�P��"O�q��	�n4���:���p�"O��IgnͲ.��#�>](�ly�"O 1�a$����4��,r��jf"O,���e�!��(P4%H�M)�X�B"O��@�g�)B���c��4̋"OpI*��c��X���y�bay�"O�,�G�ҏ�v����ڐ��"O����}��%ӧ:P^��"O"Q+wC�.����C4B.�"O�=�QeR��L��oXC/�(�"O:l�`0<��!7m�s$�( T"O6���'p��5%r��B"OT$����n�Rx����^8�&"O �i ��=��I���B�6��i�"OXe����(�nxC�n~\�B"O��t�jJ��[���
�}�"OXC� �"a��A`F��3�tjT"O*H�Ƒ>7� �ӄ���:UYS"O���0��SC�,O�`B"OB� �OY-{CtQ:B�h�be��"O�,��Ý�(��i��N/�.�SV"O<�1#-M�u��0SRF�#'r4y�d"O�l(ElSN��:S�`|� W"O:A)c��m1�4qGDI���Q"O�1ʴ��(�,�с(U=��0�"Ov�2�	��s�X�����>��	"O�й$،=ӌ��&G!�01˄"O�(D��f���bя�a;����"O� R�a,�M��eH!O�d��}""O�]�"�Z�N��#�&^\����"O���&L������?��r"Oԕ��IN�B�Qz隐"O�u8��µg�B�эD2Fn%
"O�9�ELV|�= �J�=AN�a"O�!��}�\����S8?(���"O��a��Ɛ �b]��M�r#~E1R"OzI�K�<�f���l�
_de7"Ox�	�]�G����C��#��h4"O�m�֥E�n(��,��|���R�"O�p���۴a�D)�E[d�*�`"OЭ�Pb��R�ڰc֜1���3"O�0�����0S��լZ��h�$"O@1���ɴ.���Ң*��9r"OH��S�
7�0M�V̒k���1"O���S��.EO �ФK@�N���"O����J�*.4xGˉ�gW�ɉC"O�L
B�hL�R��9P�9;f"OLDK$�"?�$��(_�6~�S"Ox�P+�/J���脧ii���"O8��E���%؊峤�ш@N��"O��Q&�9�.U�5�A�	=����"O�YXQ�	9G� 	�O��+1|{@"O&	[5O |���P�nȌە��QB�<���u�x��^7R����D�AA�<�q�܈(�:T�$)_6I�A����<�ϋd�]bcmȶSfbLp�ƙe�<1�F\� �A@"(ҷ:�)H�#f�<���H�F[`=b���3'�]�<Q�(��8*5rEl[4`�0 @�T�<QG�]
U�ԙ��ș-D�ĵ;�AAS�<f�Q�����"n�V�k�K�O�<y���|��4�˞2�XCt��_�<Y�lςD2�|@��
>�����U�<�7�F<����0ϖ�l��9��(�M�<Ѥ惧1�|,�A܍`Gv ���n�<�r��>w!�b�V�0�R����j�<��U�����gF�O��P���e�<�ED�5�y�E`�Z�N���yr�	�_��YQB��#`h��5�6�y���b��[v�87p@��Hɉ�y��ŊF�� �C�hw^
#�G��yF6/(�W��^��I)2���y��J��^v��KalȻ��C�I�4q�9�sOM�������F�IMC�	�(�V�q�V�X��΂�,/�C�k��Җ璹8d\q���B�Ɋ�@��C��L7��Sˏ/�B�	=V"Y�!�]��MX*I���B�	�'Ȗ-�r�z��at-G��0C䉁n���9瀜1\��Y�O�X:C�I5-�,�h�䖦`x3TAX�5��B�
; (
��MZ�uK��z��B�ɽ;Nd=)dg�#�����/֥<?JB�ff���n׿9���$����C�l��qpV�D�f���ӣ��l�lB䉿B��mR/��]�CTHR�JB�)ߖ��0����Q�fL�C䉖H8�`�4��s܂|@�kO���C�ɱ~�⧄ۻ_�TTR�̠Y�C�0YCd��pY�q��0R�/ˮ��C䉩 ��,�$��f�X����yH�C�	"�0(&D�$���cnY+eF�C�)� Fѣ����{|#��K6R ��"OP�����rY�	��3>���"OL��%���4����7���"On�Т�Ϣ4�:���%H!;�\�"O��C�F�7F�>��U���8�"O�	4��G�DY��D�!8���Sb"O8U��딠�葨�Ý�8�����"O��Z4$��J������%P��t�f"O|]x�Ə1?U����	"$Ԕ��b"O:�(g��<�E"U����P�P"O��:R	<)[d��&M������yr�\?-l�\ ��� ej�e��y"�[�_P���-V��r(�G��yBo_�n�����ص;w�I$�y2fF�X�r���|ɰ�#@��*�yBJ�~�}k��R|dH�H���y��@-^�����?r����%���y��;���X�l֊h�� �J���yB��Np�ȁ�>R=�<�.��ybǇ$uń�f�!=u�$�y�#R82O��A�D�ane2d�@��y�[��p9��֩X7\M8d,��y�*���v�T�`l+'���yr��8/:x̪���?}�ؽB�����y"hY�yx����k��ѳGo
�a�!��ܼk)� t�M��p��.�0E!�d
-	�e!�k.�"��E�w�!��&���ņ�0~�\|eƋX�!�D=9&-`r%��V���q#,Q�E1!�Ě ��i�5#G�
��[�剅4�!�χ|��a��MB�C:Mb�M�!��C1Egd
C!��k	���#�%!��ZeV1�)�<ea�5��N��!��L�u�a�,<O,0��F�T�!�$F�-p�ո���0v;X-:0̞�]8!�$�3�.5���K���T�� b
�'����BE'�F���T�9Z
�'h�$��j\�\����'��MCެ8
�'Ŧ�!�$�w�84�6LQ#EޠH�'ܒ���j6O��`���=m����'F&	�n�NX$YE�Y�g��0�'685 #fQ�A��슣A��[9�up
�'�N���'�P#%H-��[
�'!"x*�e��y,�1zƘ�m��@
�'D4��6��d>8�� ���(��'�$�Q����<p��ώ}b�A	�'pFH�MM4Af �Hmd���'��E�A"ץ:VfAs�ß�G����'����؞a�m�怌�>e�ȣ�'�r���	��p8ƅDc���'a�8�!k	9�a#�c�6%����'�J�	%���JM��� � �p���'���P���\E���������'B<5O�1��4!�Ƃ6 �����'��ՙ3o�!r���I�m����'���i���3r�� ^�i�RM��'.u:���^�(P��)/�t�R�'�.(`�ğ�6YY�"��)e�"�'D�\��(�.-K��헩l���'
D��aR�����d��+�u��>D�)���,�%G��
��ݳ#�t�!��amBXs3�H�	��$ڴz�!�$P'�H�c
"i��ɡ���>!!�$�;}X�d��X�U2'�O9�!�� d��'�)��$�� L*�2�"O,X�o��tn�5"����M�$\#"OVرU#�)�ȉ�$
)�"OF��̙� �vLA�`�d�� �"O\�2�#K�������	���ZB"O�x�Vʔ�$���AM��d"O�8����#2�4t����2st"O��5�� GϘ�Rb��݄\��"O�����Uw@�В��&]����"O���D.�/<?�	��E d�`T1�"O��*l=�FHyaȈ�R�S "OL����9w���c�c;x��4��"O65�vfT�>~��"��
�V���"O\1Э�;@1�D�٢�g"O`�Is��X
�N��d��xzE"O9S��F=^��8GH[��&���"O&���'P�Ji�F7O��`�"O��K��ޗ'`` k�ܒ86	� "O��;Ԅ.��xJb���lh�3W"O4�����53�V,��CInR�4
�"O*x�d�J�h���R�I�_�H�k3"Or�i���y c��0ժ�"O�1�'�\�=H�A˓`˸�(��"O��L�%���5��a�"��'"OF�8Q�1e�d�� �;��(h`"Oh��� �%��JM�4�(��b"O`���g�ҝ�q�4YoB�R%"O>Ucw$�%"술��<���"OBu����^�xU��j�p��Ey�"O�{�%9���`	�7�ѻ�"OݚGE�{��C����"4>0�4"O����E�`J0Q5R���`�"O\ qF�A��ꝺ�CR����"Oz�$
��p?�h8$	�<O�SB"O=r�%�;/�^x+�:n(H!�"O:|�(ρ9�L�b�g\dn��p"OH�z�A^�%�`����ڪ� "O$%�1�U�
��(�B6�.ic"O�ŻV�L&k���.F S�4Y0"OⱲ�P�i�
y����(4����"O�!@�gۆ=[�X	�3���
3"O�ڡ`��T���[�ϖ}Ѐ2�"O`A)����I�f��K�1��"OpP��c�%)��E��m@�F���"O�P��X�<�xHђ�����{&"O�MjC"�Z���J^9f%�(g"O�5cW肓O�Bq``ǚ��Jr"O����Zɰ2O�?U\��x�"Ox���8�t8m�[L� v"O���Æ� NQ���B�žsP���"OP�9w�ϒ�8rEތs��P"O�,�R�g�:��B��!�`\;�"O���㍑ھ�s�%��[�L��"O,!�@EG
3tPi��U:<l�'ZΜ ��H�y����Ԭ�f�p	�'P�i*s"_^^Ll��&�+L��'���B@�fN�d	%)N�t[$�"�'Nx��j��2�8(Uʗ3l��q��'����_�<J��3`@�fcL���'ZN��4���/Kk�n��L��Qb�' *q�%(����#�J$ \��'�R������`�B�NC�V�#�'O8�&�*/�����E]�3�M��'' ,
��[�1���v:*#MR��� ��X��:If�c��T�3T��"OH���זz�RDk��.���H�"O��q��1I�	�fJ?v�Z "O��+�/`����q�ٰ'��A2"OTԹU�ܦ0��U��I՟�� K�"O`A;���6�V��f�8�tDф"O��9&h�h��ܪ7(B�2�̢�"ON	�h�?��@Qf�.%v�e��"O()��ōP��䪦B�Is,�0�"O4 [ ��`ZR0�W���jO*�)�"O\�b�F�-ۨ��a�@<�i�"O 5��lɬ]��(Ga� �ՙ�"ON�q��� �d�XF�ݤ�V`�"O��i$`��py����B�ӥ"O� I��]�I�@��u�,��"O� R&�t��5*��uW� �"O|Y#U�L -Q��� =1б��"O~h-��|"R
0��"Oʨ@��R�R�����H�2�"O4 ta�R~|B�E�,V �p"O���f�~Y�)��DO�(�`1�R"O��)��1ew� �򢂑c�1�"O&(`B˕�$��7�@�։��"O���o�R�fY15��**�꘺�"O`%��M����ْE�:�P!"O����C_I��ٹ�J�a�X��v"OV�ā�3�
t��H�D��h��"O~YBsJR3x��qPFQh���v"O�p���q�����@0&"O�tbW�E�bö��aL�'���"Oxy�W!P��ԭQ� ��"O�1�B>.�n)Q$N�<Â���"O���s댭g����Y�?�V�*�"O��ؔ�?7:��I��L�RI�"O���jY�=@x%)`_"�i�"OP�AbJOx��j��GN��"O�1fE�D�:��į;
�Q"O�P@eI=5(B�����`J��r"O4!��[�pV�j� J�y<J)�%"O����ܐ]1 �g�0U����"O�hvjCm�5xB��31��x�R"O�e�l&J����U���3"O����M�0B��Cp�+��h��"OPxY��U��$� %�?c��8`"O�(�Ԋ����D:>�@D
�"O�)��,ӂ3�̢�T6 ����"O���t��0)8���tC��>��D"O. 	!h�_M*D#i
T�@�D"O�E��#ږ�̤�Q�+Ɗh�"O�<�G�@L1f�!���'�� �"Ol��W1���r!U1̎��B"O�u��b֚	*6)@`�"I��� "O: b�ᛡ �D(�s.A	B�<@�"O���R�7,P�����j�t"O6$ǆ\�~���"+��v,�	�"OJD�e@%p�X��	��k����"OB�31�A�7����#��5��:�"O�q;3m����+�I�1�t�w"O����2��ݫǪ@�dw��af"O�p1U.��*:��0��36]�m��"O6��!���l1u�_Hc��r"O�HԮդY����F/ea~YY"O� ��j^7M	�V#I�~G�lA�"O4I+�i��M��h!��[(T�1"O� ~d;Љ�e��+""�I���p"O"����f�!�¯٧�ix�"O��IF�
]n�zS��KҴ�4"O�G=l=|Sv�ʖ3�֑��"O�h�s�Mپ� V��>��HB"O"a��j�G~��`�-ۚ*ʤXP�"ON�S��2j+�]Q���>A��q[�"OΜ�������%���'K�U�"O�ۄf݁;��!J�D�2w7dp��"O$�w	�F�0d�S� (Φ̀D"O���`�1m dK����t�ZE"O:�!�-D4|���U8�l �"OhaD�$SX���u)�U)���'"O(��ĉT��)�I Qd-�"O�Y��<~j��q�ō��,��u"O2�䄽,:�90��b�԰�"OI����3��u�����e�"���"O�E��P.m��)���%����"O�4�s�Ќ��S�ׄ{��] 2"O�'mM)lf���U��!Vm�"OFX�AȶI41K�N�t{�q1"OT���MD>._��t��u�\ �"O�<�s�,6~�0%�U���*"O,��H=l����ߌuڣ"Or�e&�M�tE��ݔb� Q�"OX�[#/YDL]����H�pM�A"O�mPp�E�j$@,�f�I�%"O��Hp���Y����,%��"p"O��t�ýB�Jp��Ɂl�Z!c�"OT�rĜ�V9���S�9���"O��P��AF��W��(#����"OR��q�M�����>b�ܱ�"OtY@���ܼ�6�M@{��C�"O �B�`N�pBj_���W"O�D�C�Їg��!��2>��XG"O(���(�/<�v�z��OV,�!�d�5>}��D��S� 9h�υ[�!��?��\�`�Q��qX��1�!�d�+@N���I-1 UZa`O�8�C䉌��U�b��m�PC���. ��B�ɶC�����Y3L�̈�a�I6�C䉍l^&H� �� ���kG��?��C䉭?�NY�b�K�8#���S��.l��C�bc���B�ÁG9��ᶊ��Y��C��)if��n ?X�(:��f �C䉚>B�s���Xo���@�<i�B�yHE�MF%隈ҁ`ί7ĂB�	:r$Ty�A'T��H����u%
C�	E��j4*U\Qb�K2ML���B�39��X�D���x�R�0w��}=�C�7K7���D��`�H<��+3�C䉎-`�fV
*�0l	M�G�C�I�B���ũ��1�<u�C�OqD�C�ɶU��@e,3r��,���cTpC�I�
��"7�ءN���K���t�C�	�kP��d�\�����F(j%�C䉷�4!����W<��b���B�C�I�^B�I`��lT4�8E�߆[8pC�I-F0b����%_hl�r �Ct�C䉾C���̔V�T�S�ͷu�TB�I	 �vH��M]A�^�Y�)M��PB�ɪ>t9
���O.�!�d�/n�B�	t[����L�X�)��윢�B��rv��{F�՛P�(����?&��C�)� za�LI�$PX S�f^�dA�"O�����q)&9kE� /��K3"O���b�bqxI�W�ĕ�,`�"OeK5ϒ�91(� #(@&5fu�"O|y�֎p�z���U10�Mc�"OX�+d�ͬ�tIV�͆ p=�U"O�h���P�ܑ���]8B����"O6����+j S��ڠ��"O�H�bȼ.B�d��LD�F��a"O�I �mސX��q��d| Ĩ%"O�Xz`�K2*�����7vzB�0�"O�(�-։k�D�ɕ��(6,�)�"O�u����(��
ӉS�d����"OR8��.��a�Ï:a�b�ڒ"O&�3��ڤBPx� �AҪQ����p"O�1G�]ܺek��[
?yƙ�"O��Dn�~؈gL�?iw���"O�8G� ��&��RZ�b�PAr"ObL��ͨh0R��De� `��"O��Y�ǯW�����Ĉ&X3"��E"Ox�C��-vZ6-{�8h#���"O0���ϸ"|0"�Λl l��"OT��T+=
)����E ^�`C"O��`[/`��g�=�E�"Ot�����*G�<p��Scߚ\R1"O�D��(;ˮ�c� Ο���)'"O��(U&@
$��NX�>⢰��"OL���!�C�P��m��I��@w"Oʨ	��D4!~`���.Ǡ�r;"O�AÇ��v"��6 R�B�
�Xf"OL$���A;VS�lx �%$��1k�"ObD��i�P�ړn�r#�}��"O^s�	�CQT-�Ќ_�CD"O���qk�� p&��L��U��"OX�B �����iC���V�����"O2E�q*��j�nh����nB���"Om�cׂK����H0gkxA4"O�YtJ�$o�l���6��Q!b"O������!1<�+�c	"-��*�"O���j�X�U��Qp�	"O8�K�	߫)!HX�f��!KzZ�("O)FW�F�@���,^q���T"O�`���[
f0+$a�X��Jp"O�|����\� c�W�y�:}�&"O���PM�5x|Ĩ	B���Q�JcV"O`�c�l���ش�\(����$]�!��u�n�)ԃ��U�D�X��
=/!�D�,���EoY᜴���0#!�D1݈QCSc�K�~�bB�W!�!J�fhʡ��=?�0��" �!�O�%�#P����fI5:]!�D� ��\R� �|�x��S���LH!�D\�+9�H���U.b���h��jA!�D֫c�� �#�HG�	��K�dQ!�J�2)vi3Pd����8+�IS�(F!�D��MS���m8u�1�7)�	;?!�Đ�f�E�T��Y"-1r��4`7!�O�f>�+�&L(;�02��x!�d������,.��y�!!�� D��"S��4/.H	�oF��!��ΈqM�1���-G����5Y�!�d�-� �� ZV�� Q5m��s�!�$�-[̔Y�0.�y`r�L��_�!�DH� 6����	�U�5H��s�!��  �G��,b���@׌l+����"O^����75p���脣G bQ��"O�ڗD �B����Y;� 
w"O��b��H�@ ӱ S�|�8�u"Od���Y�8�nTx�4P&�Z�"O���s���s�-�!M6��K�"O�M�@�Ko��x9p�?2Z��u"O>�[䋛��p��ݺu$���"O@=�S��q���h3vt("O���@��>���!(Z��R"O�%��c��tƸ���8���z�"Oz S0��Sϲ���Ȓ�p�\�p�"O��'�/k(	ɑh���b�*G"O*��RgL	h�����5�u��"OpA��W-��Q�'�0�B��U"Oj}�Ɓ.7�~i���9.ע�ʥ"O��ٴ�ٗ@�j�0Ca��Y.b��"O�x�eZ	S��5����6#D�
""Ol�b�V�����T8z��i�"O�h"1k��Iת��l��"O��K3�D����R��M��"O�LK#̜t��i6���!�:Ab�"O�Y��m�x�Z=�@�B�=���"O���2M��I����g��):A"O�Y��WrLD���4r�T�"OlA2���(	�����,d�`س"Op����*&Ȟ��ch��h��4"Oԥs��]�l��C���Bb||Y�"O��F�E�m��F��W<p�˓"O�L����$�����8�!�"O^\��Ϣ6KZ�p/�-<X�{6"O �X��Y$Ղ<2��,O�,�z�"O��ч�|�T��M(I3��#�"OP�siɠ�~���FU#:-�5�"O>�WhT<s�L-*�d݁l>@h�"O����������!G�q�>��"O���X�lz-�FB�"�8��"O6�yt�/��+˕�C�b�q"O���q*�<1�~�u��'*Ғl�S"OȻ�Aĝ|}H����$��tI�"O���PDǟ64�9S2o�!;�Ti@Q"O��ҧ$֢.�$����p��R"O���3`ٿ�(�s�C�6� ��T"OPC�F$�Jf�;A�yЇ"O��{n��&���ۓ'��gȞ08D"O`$�B�l��9���6��p"O��u�X�#�LHxץH�w�0��Q"OԹ�wgGb<��t"�Q�)��"O�x�uF�#���2dB��RT��"O:�Bvl�9D�U5�n�^���"O�[pÐ��( �F)�.��{6"O��"p��BE@L��Q1��c�"O.pe ;����h.;�� �"O�K��&<_�a�FJX(�~��"O�Q1�cGo�2��G�V���XT"O��e�r����
��34"Oшj��I����Q�D�BjV+=;!��D^�2�\�h��z�Y?d!���Df� ;c"V��۴)<!�MM���[(|� \�3!�$WV����d�|�X\{���!a!�D�[�
ePV#M34�`!��յ�!�ݦ���r�dق��N�)�!��_��+�K#?���LIO=!�� P����k���q�	H�5ņ$�"O��8��.6�6ęt�Â� �B�"O��&�Bi0d[5@�7[X�&"Oh|K��6O�����U��DmU"O,p�����@�)�n�!�\�c"O�j��#|)�a�Go��em L��"OpPPƋR o�R��#Y0-��"O�p��-NPq<`��EN+E0�x�"O$�B dۜ�$,�]��!��6O�!�d�%Z�g��;:��J`�)�!���=j��ڿAU aA�Y� �!�D#F�h� ưcNv���K;1!��<]��1S"Ӧlgn�	�Ȋ�"l!�dS�
h�93o�,nUN��Ɯ�a
!�d�t�8����&��J��W�&�!�$ۺq�bI�DL (~������?P�!�d��\���ڡ�ږJ}�aSW Tu!��W�!]L�U�[�@}�Q��%�}�!򤓛$�`�����py�� '5`_!�D�"yV����V�k� 3���Z<!���d��W�4=M���An#w�!���art��AȷJf��)B��1!�҄8��h���/���K�	ŐI�!�d�e�[�m�=U�8bsV�<o!�3Qv��@Pb���`���ۺc!�R	_o����O�c�R�˔E�q5!�D�*q�:t��	_�:��V��M��ȓph�̃@l��J(I;�A����$��?V0M����W8U)��I�`���6��%�N�bJ���'o�j��ȓc�I���Ѣ6�8�Q�`]�x�,��Q2��s�L\�Y�$"_�Q�T��;3R�b��:S��%9�7¾���N�FUs�'� =�X�,\����ȓljl�Ӱm�#5����[/Q�R���~����c��/0��a��g�(H����II��Yi���F��(;$���!8��c�*.<�� �ǋ��5�ȓl�%B���>V4�1ͅ#H���ȓ!�����Y*DC��f��@�ȓH��Q����1V ��JB{��L��}�����S6(e��MB=��ȓ;Ld1 ː{�d���M�"d�ȓ3W���Ɵ�C4,X I@?c]�ȓj|����,S���"�/gZ��Q�,�h��X�fT	�ĖV-=�ȓ`d@�
���n��<�+ˆ;��)��$� !� �Qn������m:֘��hμ��F�V����C�]i�|)��n���h!�ZY}
�@�ڀb9��ȓ,�b������	84[fƿi�A��vmz���@�"�\0���5g���ȓ,�r�;#[�
��m8q��cڬ��b�"a
Q�ϽO�"���Z2@�1��lj����n+4��AL��BƉ�ȓ/|��ֳc��l³	�1{kf��邀�� I�	@�M�ɔ�9��1�ȓZ��,����c�)J��k-x-��fJ����R��A��,�/U-<}��fX���!ͥ`�<���-X�?�4��^Ș�[��h�.E$j���ȓE�*l�q�_�:��&O5����dzP8f/R�<�B̻3����ȓ�ڠ �E�	��;�^��-��S�? �ICfAؑN¢��E/
4> 8K�"O�)YB�
w HÂ��2:���*�"OаQ�W�=�M*P�ؗ"���r�"O��f@ lO�X��	�I{���"O`��O��|tSI��^�"�"O<��V��:bTx���G7z���&"Od,� ��- �������=�J��"O~y[c���
�ȕ[wkWkt��8�"O�kP�ƹr�Tl��	�iD[A"O�0���]��"ā��4h�@�G"O � %��&�P�{�kTJ>Ūf"O�l�i��c���HAj�)\�A�"O��j��O,N�@\��fQZ<�C�"O����KΨK�yx�g�52Ξ ��"O�@��A+p&|��� \�"�X�"O��s�B[�y����ơN|b��"O�����C	;��A��#\q�ea$"O�X�J�4��1��P�lY��x�"O���{=x�2�h�
6�P0�"O<DR�-�x�!1�y!D�x�"O�u≔+M�0|���M6��f"O�
�AE	��hÙ3T���W"O��c�#
<��E�̯���q�"O4iA�.v-�E���.�L�@"O~sDGY�`�^L�5���(x�y"O^��pX�E̜y��hoDk�"O�EۉP��'�n�&�"O�p��ˁ���g
:|88(�"O>Q��K�>?��2�E֮`� Mj"OJHC�ʢS6��J�f�-�ԅct"ON̚3ȑIa��u��8Q�L�ҕ"O�"���xd����!`�4�P"O*=¦��L%6m��e���:���"O ��M�N!,� D"z�<��"O��Y���~)(�k�c��|��"O�)�G-J��-�"���q��c"O���0��f&��aWa�0<i<��"O��sE���>�9����I~ؽ��"O�1₌8�E
�eE	Q��Q�"O����ֿ=�ʹkg���2a[S"OR�3��G�Al�@���f�2k'"O��)�Ӭ?�*=�7�%.�^�c�"O�a� �Q��]+�E���(""O��Qr��$�����,�vẗ"O���"���`�FN2�
�"OF��b�ӺH����M	�6�A%"O���M��2��8�L[�	��H`f"O��g�B� Y��A]6����"OƘ2�L �f���a˵f�&ɒ&"Oz
R�O�lI���֢i�XQ	�"O��"����\���S?���X"O��{��_ u�����֬=��b*O�i9����rh6����h��u8�'7|�%b��(�AS)F�J�D@
�'$-Ɂ�S�T�����ֳ?;6�
�'&��DF#S��с�=1����'9�ih$e8L�ɀF/I�)VDi�'>��	�`�%��Q�2-;a,q��'�
��H�=)jA"�9�"ɚ�'�!�ӀZ�Qɂ��1��3t��'����UG_]�~�
A�ԭ����'���Ѕ��/��K%J� Ğ9�
�' �T�����9��ڗh�{����	�'�>���&ܼ��v�[AX�]2��� ���b�UBPVES��Ñ?�x��"O�Hy�íR���C��m�:H�&"O�D�t�֌u�6��!��vvāY�"O��p��	�R	T��c%%p���"O�0	3��J�m�c��1"O�c��یp#��Js#!Vń�h�"OԼ��'�Rk������j@"O�"��*}���C��~	�7"O4�ۤ�����C��v�a�"O�p��$������㔇;u<X��"O��rK�x�9#C�D�y`f؈�"O 	�-1A��� �
�Sm!�T::��i� �U*,��0��&�!���b�"������T ��{���/ �!�A$b:���/�e&�(�KZ;l!��ՖP������h�i1jH�3Z!�CW��-1��t���)]!�d�PǼ��'BCv2(�b�!���&�`��1�'@ٌHKgS�!�$����ZC	ǓH���ɔ��%%!�$�0T��ə�B^(S� ��5�V�`	�'��(��R�^��<���02�TT	�'�������s�pǆ	)�r1�'}b};���ey�Y��ϲ��p�
�'h�ye�@09�)��H;Jb��9�'!ذہC��b_�9ɧ̓9>0��a�'}���pL@M�H�I�%a�T��
�'�z�(��އd%̹��T�v�	�'�콳1
t>���pF�FE�Y�'�ɠ��9"5���I7l`��'���p)�='9�!��2��y+�'���(�ܟi��i�N�+�x�'A<�B�'�`+���>lD�"�'V�=+��C�8����F@f�T���'�NmHנ�04��Q"�ZX� 
�'�`�&
X� K�E�0S�d���'�>lj��}�l��c�K� ���'��{/ڟ����W�\*�x�P�'��ɪ���A XJ�y@���'�tk�D�fx��ᱫ��U����'��}���_<��`	��Ce�	�'oZt�5+��C��R)�4��5��'�FUqLȗzK���s��/_�c�'N�xy�F�{��,ic�@%b���'�BhK��9B�����G�%#�ly��' (���E�
9�� ��ү(#���'
F)�6g"��4ᚠ�R�Q�'D�����(��T�G�K��� �'��k�@��|�!�d�J�^��'�`�h� H�I��eC抪>�'B�պ7d��v�U90�ۖ?Tx���'�xH�3�ߙ{��I���[�n�(Q�	�'ώy�1(�4`�`�&Na7���	�'f��Ã+M�c@�%���­^��M8�'���֤ƾ	�P��/@�?!b��'�*E+*�1V��#�^ 73���' U P�_�SWz�r*�� P��"�'a�dK%����4����P+ٸ�'F�M�Ң���P�X"��H E[�<!e��tX-�(ԗ�A�ЭVl�<����Mk� i2�+I�LذBi�<9U<k��䏽aF�qdS_�<A�پw�`�c�@ֶy�h5p'��S�<��σ65RPi����n���3���Y�<� �(�F"T�v
�S���'O��a�"O	9e�̎d$B�23�̎__1��"O�����y��Y:d"�$DO�0�C"O~ y�`Ѭ4�@I���I,,$��&"OS�B�Pa�$a�@�[��h8�"O�*� ;�ڱR�a�'� 9��"O`M��(��@0R� �n�j���F�O^��pM�<�j3*؉]m&���'�J�*���|C���a�W����'�@�q��߉xў�pa ^U9rUz��$=,O~�zb.M5`�.͊��v��	:C"O긱�#gb�.w~�y�b�>�y��U�u���8d(�aJp+�d ��0<ў'�O����4����G�Av� ������*,�����aF6��	Q�hB�+/�]y��X.�����E�<F�'a}2�DPA �E��v�.u�p*ن�y� �h�~u�U�ӠhͰ�b�f_��y��Z\^͹*������0���yB�B��W�ш
�\�������y��΅�\���ĝ@(�y�&S	�y��l� "<E���.��]2F��~�&��%���y��G�<a�u עE���Z��y2�ҷ~��
*?�(hZ�
ڭ�yR"�v<��bD�8�>��7��y�c�!b )�v�Ջ7_��g���y�iB3��\B��İ))���6���yR��(6P���F�"���Ş�hO����A`02�,[$w����竗�B�az����_�V�PV%Ӟ3���f��O�!��;ZL��'m� <�F�x!��
M�-��A "̺���˜�b!�d˘U|PPEg	 j�jmy+Ĥ7T!��G�J�
��(�py�ә&>!�Ш
������ݤ=ߌ
�OS8��Ez"�ǀT8 q��Dį� qЃ.�y��6��ѸG��v�%P��H��yb�"h�A���nS<)4d���yb��7$͘$�%��k�� ���yR��*E��ur��Z>oP�{�cҖ�yb�X�a���r�7d��b��B��p<��ڿn8�L 	�'{&"XaU��sW�xR�I�%���D�5<�2`�m�C�	�0�=Y��ك0����4M��:��C�6`�FR�I-D��� �ߝS/���hO>qo����I�-���[e3D�h�gA	�Q�~��M�?̎�j"�0$�tQbn�)�(�z�
͒h��� &�_�p<����	1�ep���=pT�b2)�i�!�ױi�h��2BC�U��a+�G��_�!����:��`d9��)G�!�ʮ@�TP0B�ێ�P��!D���${�>�C�+Aq;tr�	J'9�芴"O�%(���=,��b22�@D"O1ٷ@.	��'��[�r���'2�d�EcȷR���ٕ*�'QE���q�����S�����%a��t��_��B�	�XZ�q��o�����ۣGz��B�I*��h���9�Q���vΖꓧhO�>]� �����"��hR�`��>)�~
pcǨϡN$��P�M 1�ȓk&�"@��_����#B�t���INܓ��1�S	�W�t��j̽wm���6��K0m��J�8hA��l��l��S�? �Шe)��x�^-R��C5>y���g'�|f�>�:hp�p�H�(p�Th�c_�Y��i���F��H�H�pVԫF ��ȓG�l�DJ� If�8(�g�'a�N���2=R���F�QABxdc��%�vI�ȓTf���C�4F�����X �1��}|b%y�`T�4D�R�������A�* I�F�&phq�E�<2��Ȅȓ{�Q�E���mdΙ���	9+ZTy�ȓrP��RPgĂd�>u����3)]�ȓօ:��Wl��yZ�i�8;4"I�ȓb��4�E%a>�#��A-d���I̟���(6��0h^�1��q�N�f��7�<1�xrD�f��a�h�:BI�mD���:���sIH�!��ȑg)�}�O:���	!Oن-hw��:%�:�;�M-0�#=я�$�>aq�ŀ3f�� #pD (�F}g?�O.��ӯ	�\��9y��X�L�FɆ�	���d���K�����jћ+��TQF����
�y��ӓЖ)@P�Z�*�A���OL���:�8p`�T�.ZaY�!��])fsCaV";|l)�)y��E{���'~^`z��Q+,��Pa��#_֦�`��$v�2�}���W��Y�1g�5��u�V&S�R8tB�'�<�*w��4%�Z��%E-[W�}��O
���Ӳ����U.��6]SȎBv!�DF�K��x3�HV0!�B�	�*	7%Y���O
�=�jE(K
uޔ�uf�-a�\"�[�<QP���ZE�8nś�r���q~�'����ĆE�D�j�,.����T��p�<'��->;�Ș��f��P�Yn��p=�����8.α��N��N-x��BS�$%�l�Oȯ\XdU)�HT;(`��4,�Op��Z �U�K�6�`��qH��`��|�O����ض �Phq���e��pІo�`!���(f�|\�wh��*�M2��� S�O�����+����V�+n�J���;EC!�D��
�������~�v��e���&!��ƒ�ҨSJY�<2�Ap��U�f"!򄚰;�A�%D�E�r݂'�+j�!�dߨ:�(��RIP�|[�4"�AU	9��	F�'XQ�T�`��<
K�@ǫGD��q�%=D�����kt8�*�FE�?s��r%g<D��!Iթv>��[$�6������<D��x@�Ł-|�ĒeC�ĴMj��:D� ��I��(@���OCa�FYQ
5D�0R�l�#��c�VH%�ƀ%D��J�h�)t�m��((�H �8D��"@�(�H�Un8n?� q�"D���jN�Y�	Js�S.1��:ǅ�>a�'��O�>�6��5h�x�+�MF��!4g7��p<�D�?|4̹��քX�@��0n�<����UdQw���"�o�i�<�ѥA?u�\P N����Qp!�O���' ,S��>�J��*�Y��M�	�'n Y{"�
10 P�U��SV��	�'��+C�6 ��\��T���K
�'�H��d��g� 3�Z�g)�9J�(�d�<E����]�Þ
|ې	��o��\��d�r��j�;`�&-�rK<s��ȓcF��X�j�y"��BŨڼ�9��PE���"k^�T0,���UN�>���M��哫c 8�s��A�A�'�E�8�h��$=�DF�J���y�X��!�^��!�� ����X��E`٘m�lR��	��HO�S��С���ͥ���)�$4Y!�B䉕0���S�ㅯb��$�r�ޏZ�p6�N�����f�11�R��7m��$�U�V��y"I�=>,]�S���`lP��Я�yR��?)��8�F�:�({!��	RV�=��]�Gp�8Q�_-�!��&�������E�����ҾP�!�ݛl�H����
RHb�	�<�!�d�2)�fub�	>�ЀQgk8�!�D��G
���G����}(�� _r!��ϊ�0@�
��U�u��`�.Np!�$L/8{$]�O�>c�1���?]=!�\�w�l
"bX=�ɓE��:5!�Q�~�0��	:
���q-җ !���pb8���)'m�(!LM�!��X+F| �:��,i���!�!�$B2|���Hi���%G �:�!��ON��8A���nW���F_�A�!�d��K���bDCNN>jMz��\&L{!�DZ�b�&����Q2j.`<����{!�$�z���Q1E޺8�XӵmJR!��[+@si�G��3>tB��w�Δh�!򤀦#D���,�̸����.2�!�D�#ݶ�a.�M�F ��JҞ�!�^��HP�L��?nx0�I�+Y�!��X8Qv�|8u%[�-TMk��Z:�!򄍬4 (g�K���AԆ��I�!��M����E	��ㆅ���LI!�.�i���l�2�3��&9#!��h���T*N��me�R�h�!��D��sB�]#G��Ir���K�!�Đo��d0b�!TI
�D�!���=�\�A�I�Y��H��g��!�!���0$^)hrb��~�ޙsШQR!�D�&3dI�cj�:� @f�?]�!�"!/�\�`
���k6ȝ*u�!�d�x��#F0{t������[�!�7"+�aΈAh��M�?[�!�U<�)�Q��#C�p���ہ�!��J"|3Pi�W#�>:��{u�]�b�!�d�><b�����7.�YS����a~�L�ə����^�����ב"ED��Sb���y�BZ�L�RD��Ŏ�3������yr#�v�VypE�Y
Ӥ/�y�h��V5�犒�Z�$QÀ�-�y��ݣz��x�!N�V���a���y���D�±b��&K=,�eU�y��D�
ь����^4N��m;�J̚�y��B�-����cڒW0T��A��y�*�g네[d��}���+e���y��� �PCpN�p���@�I?�ybh�2Qx<m��9:�� ���y2fɖ0w����U=/���꠭�4�y2b@<�<q�4��<0q�pΒ?�y�↟}�^��$뙿F����WΒ*�y�M�$V��u�4�Y:>+B(�H��yf��q�4�ЦFG��tr &ݕ�y҈�,n�� (6���-ӧ���yb&7�R�:�$	�  ��Vȁ��y�E��d�5 ��zb�pz�dM��y2��$��!�t	�#�F%�G��y�c[�zD��'��:��7!M��yB	gI�pi�P�%D<~B���S�? �!C���,�U�f�	�8��@"O4�ҋR-h��w�#z�!b"On��A�٣1^��s��%Q���S"O\@`R��}�xh���%%�t�2"O�{C�Y�S/ �@�\|u�"OV!���e'$h��m�e��bE"OD5���ǰf]\q��ᄺ~N��xr�����p;�L�c�(r	��#�&	)��	�MV�K���H`A�9V�>� �A ��ć�2c� �V��5�"P�T�5'@-Fyb@T"3`�?Q�3��Mv<��K����H�� D��	4(�#Kf�-�RE(l
ZA�K<D����
�3rD���[�V�2a:A�=D�(�O^38�HcP�XE�@��R�9�O$�5��<I�g[�p	�Di2��,;Ѕ�3@UU؞P�=AE�'~������F��lҡb	~��L?Z0���(�_Q��d�F�3x�fA�[
���=���)��1p#QJ��y�p�©�iY�`�Cܓ�h����9D�ً1f�;7j޵�� +I�Q���Ǔ2�؉���0^� �VH�m�J���{t�$���'�$��$�S#r�ҽ�"hYG8��h��H)̋	 �����s0�W�4�x 5�>�h��Қ߸'|��#�&\�@hp�bP�lžaÍ��o��G�T���v�4�K�JU�X0dt)f��,ʘ'1`xEy��Dcјo"5�4(��^Ц�ڵ��	6����s��{�o�.�툅�Տ"�@��n �I�����M�H��xU&޼g؉����':�!�զ2z|��3J�0S
��#�A�#l\a
�'�zP)��P:1p�:GI�D.(U�
ӓ;z㞘�W%�m�0�FV�ئ�y o'D�X�NG���y ��XI����$�&YMQ�b>�:E���2R�Ő�$\	U�`I"l)D�@Kk"c��E@0K�$ؙ�h �:p��χ_���ī0��<�'���
!�F�<��!��T�N"�r��D|d��'	�xT��_�];PfQ�'MB�ӓ.���р�^�Ys�J�^$�S�0D�X��故|��,!a�+�˖�"�I*Q�b>q����\��ɕ�P�H&�H%�"D�DK��:K��R��*5�ր��� P���񤝈
�@C&�](c���1D�q�!��$�y*�M�	Pz�aA�AX��PQ
�'�������$�P�#�D�x�Q;דT�qO|Ib�nT)
��K�CU�@���6"OfH!��&��)�P�͠[��:�DPm���yx0:�(ղ'�@���/�[朆�i�v���,���
�ȍ9z�Dz��'��9��@�n�؈
��N�`�@	�'���'Ɛ�f�Pi� B�����'	��)�)��5.l�;�B�q�J!p�' v(w�G�n����U@wbPx�'��Aiq>f�`�Яh�b���'��=�E�B�;�*���	d�PZ
�'K2��4�C w��0�fƊ\V<��	�'.\�Bu��$,7X����di����'�6 ��+3D*��B4Qc��	�'h��!��;0�=�T#9��8�
�'�֕��m�-�ڴ��,�3���r
�'jJ����l��MxP������
�',�]���$�׌ҷ ��ݐ	�'q�5j��1+dn�牀?��|��'���扎�&.��OF���
�'g�ꁋ^�y������)}%�

�'�B�!D��-B1�5p��*c���� `��
 v�=kSb�q�b��!"OF݃ԅ"NV&�"���(���c�"OP�a��jkb�s��[|�Ƒۄ"O���V�"bt���i�	F���"O�E�B��?o�p�v(S(u�&u��"O�鴁�7�n������ ���c"O���EGN�0�f� *Dt�@�"O��E3�ڌ�玜�a��@��"O�`ɲ�����@@D��V�
]�"O�P�@eD�~�Ƚ�a�:�U�E"O���v�>����F˶�n2�"O���.�C!d����:c��}R0"O0`I�+Jg�Q��	E�<ب�"O�Q2r�-@����*RN�*`�"OFuR�D �(U�r�8K�T�i�"O�-�'�"O��T��P�A���Ie"O�)���"'P�9p�ձ?
f�)2"Op|��H�B̴�3��Ԩ�6U�'"O�ʑ�Ù1��j�P0�mP�"Oh���d�98�.�['D��G�p8"O�M
7��r��A4#A�^��a"O�Q�w̜v�H��BF�=f��"O�؛7�U�Z�m�/�n��"O�!c�P- ���U�A�B�Fe��"O銔H�F*ԁ��)�V�ơ�"O�x��g9~/��УzD�2�"OX	E�s��P�.uk^<K�"OZ�5C)z"����95M|}��"O�A�5�U��R`h��YUF�i"O4�#�G*��|��ϩ^x�S"O��򤀟8vy˷�
���Y�"O�p��(�k���R��b�,5�b"O = ��Dug�]3�&B�E�����"O~�"��%F3f�R%f\�(����"O8u
��ن0
fDs��L�(����"O��K3A�i�:% 0�����[�"O�Y��B�@��`(�<��r"O�U*R�M�V9�h��(t��<��"O,ѠQ���/sY3���4�na4�'%B��P}�*�F��	���/sH���$A��yR�?@�b�L
k����Gθ'܄���C�'#>�D��
�9l�,�AX���Rf(�yrnV�F)�G@�:���B4n�2&��j��L"z��qr�=y��L�,b��z�����r��]"�/>$���ǥ�=lڌ���܃T|�4`6d�_����mX!�-P��C����cə?����Nќ|�&��e�?,O<�A#��:��QX�kr��cIm��E�A�$�T͑E��D$B��9+��r���1'�vJ�j�4B�'O��"�F�m�x��\�TqG�Կ8�P����dh��5�R.a�P�ȓm��CtfL�77��c$�
�♓�._�@oȌR3��:FPL���ɞ{�g��l��6̗�=@���*F>�B���f�A4�H>�Fh� �!U�d��R�G�̻�	4Ȳ	z5
�nx�d����*� IQ���o�D0�3OY�W��(��Ms��@����#�V�^�^Ic_�I����J!O`hC�	�'rT�jwmM2y���T@ދ���d�r)w�A� ��E��Y覡A��	Y�M���1�*W�bB�=�����y��d8���a�ցA~1pQ��x��D:Fc�*1f �G��Xҏ���|FZ��9�Jt��%RW'R��x&�X���Pq@X,-m�5PM�bjH9�C�ύ���&zC�]Ppl-<OTaj�$EAjN�R�Q/����P�'(�z�ԈY�b��t�Ňf�:�a��a�(a[�ĠV�ı˓��+\���Ctpб��c#���"���z��>'E ���!�T  44t��BBM�{�"A�'��<0�1q�[�<�3�Ԍx��������g�2͒��؋>�^��wɊ�hN�{FIӭ+܄��}&�� �`�@_�u�\Z��ѷr�A�v
O�z�h��LA3��e3���d恂S�<u���67R�xv
)�0=���M+30zl��"�2;��6�
aX����fp�)�s��@U��iE+�8}P�ڑ.�.Ry������y�/�!W��XZt@W�F��R� ��8����BC��1�Jџ�(�.��E+ܵV��q���/��]�B"O�q��BƢ`�at��z�<u���}+l F�ZV?Y�������	?b�0�j��=q��`�MNKlB�10eb����͘	�AB��@�I�Vsf�X؀ɰ�:�O��Z�)\�n���E�Q�t�D�'�^�EO G}"�M/#�jX9�)G�b�N�9f#S��yR'K�Ĩ��O�\ad��E���y2ݑ!<� K�ȓ;@H�%j\0�y��^lZ�yq�T",9�3J���y���%+Ȱ��oQ9@<d�:����y�.E�(��ٱ��2M�Z�)��y�Q�Ug��Z��T�x�$�!����yb���~��h`�l�}tQ����y��6��ْ�J�F�����y�/��(��qB</Μ���5�y���'���	�$���q N�6�y��J�u�ڸQsJ�&�N%-���H�'�h$j���&�,��!hۚwx E�
�'-H���I-�4jP�Kx�V���'��y���9� ѧa��$���	�'+$��u"`B5qPK�6\���'Tb��2K�sP�h��Ύ����#
�'`(	�ˎ�m�.��*>"Re�ʓ4m�<u%��3�"	 5��k��@����;P�3$<��t�=��a��5�P�B ����yC�) 1�م�~b���֏� uz6���B#�|�ȓK����D �	 ��&��,X�d�ȓ*��U0�Aګa(4�:�f߄V�L���o� )V+�	H�B��q�ąT.���r��ǎ�$-��3���b�"`��숃�i/o�~0�����9�� �ȓ==g�F�~�s�\
Q���ȓg��Sӊ���ܕ�7�6Y��� ���OJ4dgV�[��R�>�e�ȓtЄB�E�o9څ���\f��A.Pոg��8x:H1�A�Yvr,�ȓF4�"Fr
t[wbA�8 |��ȓI�ݲcc=��z�j�gR�ą��d�b%M@�ڑK�2+�p�ȓI���J]���y�,	�u]����S�Ƶ��X&I3`:	�y2���ȓrvp���,��!��U"F�܅ȓQ� �b��H���h]*1��|!�9D� �cM̉vB�Q!dM�t�䓄�;D���񬀡_�h"�iͯN���U�7D�|�#ÑE����圲�܁�Ǯ/D�Ppro>̢� uR���A(D��"�FN>v�tQ��'�0���{�i&D��!@*2TP�`��YQf�pq@"D�(p��%E�Vxc���^A03q.>D��QW�.c��,#�Y�K��;D��B�-��_�@�CF�2q��y�G,D��	���7�:�x��S!/Cp��,<D��i�b^�F-$����9$�0�B*/D���������#�̚Q��#7D����#Z�|�r'
�m>�&g9D�T!G����t�ъ�>,P9 *O����[����ր��r�X�Q'"O� �����O�X�
�8E���`q� "O"\	��Pj�%au�čyΈ�b"O�Kv%�e�v��&$��5�\mٕ"O�`�3%C�/�EI�"^�]�Ih�"Oȭ[�E>���W��X�,��"O����0/�� a�=@фX��"O��8�ԵV�E���A�	�zU�g"O��6�Պ!T&�Q$���1���"O� {U��F6N�q%j��65�P@"O�e�3 ݯj梑X��C�@+vlIu"Of��'��OLq;�.Z�])�"O���2>8\����5S�HC�"Oʹ�ej�> |+0㞋"���"Op��a�*|�
�3!bU7$���pW"O~!¦���tX
�˒h�*����"OnH���w�(�̙V���P"O�	���S��}����:�QG"OX(�f�Qx��d�W�T�"O6�!F0p#���em��R�:�H1"O���"�X}��A���qհ ��"Ol@�C!ܛ.W����B=��"O\0*�O�`�v}p���9��X" "Oء3�F!G���1ϛ=N�����"O�ͪ��G0 ř@��9��3U"O|pq1IW�#J$� �F	�i��"O���eL�	3���4 �<cc�Mڲ"O�;$N/V�8�� E-bbm�E"Ovyr�.��|C��B6 Z
�Pb"OJ�
� _.6�Fu��2I\$H6"Oؤ�Oٝ-�d-вc�{A^P��"Oس���*7 �� ��HP}��"O��I���A2�M�W �2 [v�"O�)�a�	�H"�PK���9G�"�"O^��6��9'�4|�M�.EI�@��"O�Cǣ�a�vA�b�\�k��]�d"O ��K%	q��Ci�:�~!zB"O̤�n�8H��5:'A7�jԸw"O��Xz�P�Z&=�|��"O�u�����a� f���$��"OF�R'O�P�&4hĉ71�j��"O(���+Cn9`�Q��2	r!"Oz�g�˔2�L�c#�`{w"OZ��b�ת�����	V��@�0�"O��s��F�Jtc�H�*�
�"O`U�Gō_�XP��gö���P3"O��I�!��@��Ek�D�+]@x�"O2	{�珐g
����ˀ!%�AR�"O��
�םv挍I �Q�v�9��"O �g�9C4>T)�.B)��p�"O���k[�I����E��w�D3�"OF��D�5���Gn�~R�i�"O��zf�\;@n�p��|�
铒"O�C�Ř�\�č��)Td� ��R"O<ݐ�&l��$ڣ��/���K�"Onlz ��$��Z�!%�����"Ot����F78�:
��6gjph�"OD���'}�be8S�<y�a%"O8��Ĥ[2�~�2�M�2��5!�"OΙ����ꔃ��o��	s"O,)ɦ���2_vDy�nP�Du�`�"O�)���:&�b�C�D�]֥r�"O� j�+7��xO�7��E��"O��ceC�aM�Em;Y��#�"O��x���!/�1Z��ظ�r�"O� ����Q6
k��d��f�MT"O��%�]$v��l򱠜/:t0 +U"OX�:'皸~������ i��A#"O8�(rN�<Yz��p��41��q�"O$Tk%`,{F̑��WB$Ty�"O��Vm�*����	����S*O�e�L�7*�
d@G���'�~(K4́�&���#FK&.q8�;�'�x�P�N�7J%C�I�".��(�'���fN�O;��
��M#��}�'��Rq��+`MqR�Wފ�Y�'+z`3����ȁ&�A�\�'�^U�� ijl�5�����3�'m��##i�=I��=xU�Ҟ<����'9X� i^�p��
s�8V�Y�'M4)�Q��t�hQ�"$�e�i	�'Ƕ� ��[�'D��R,��r��p��'��]�4ûS�µ:��Ȉ\��@��'!��z���ŉ�J�ܼ:�'4 a(q)ŀn��`��<Cn"���'� ,A���<����ŀ=�R�	�'��;�n!Lv��5 1�����'벼9�cX)UB���Ɇ9|��A�'��A(�N��޽R�أGU4��'i�����M��ђ%��i3��x�'�Yf �ʉB�N�1�i`�'������A7Z����0�� �	�'=�Ty�Gԅ6bHQ�B�f<v0��'�B�ٱ����%��X��q��'l�9v�C �
՚׈O]�j��'�|`b`6DU��3�><'T���'-�|27� �%�@ xbn,L��J
�'�Í�(��Dn��t?��R�'�`,�6gW4����D�X�
�1�'�.xP��@-QE�գ֣J�<J�',�]�v�­$"�z%iZ�:p����'�@bES� ���S#ןE�� ��'��a�wg��@��|j�/[�.IXc�'6,�ړ�N�0qȃڵ=r%�
�'��(P4��4ھX
��=־%
�'ђɗ��"hȔE(q�.ik	�'5�кd�y�|��R>EԼU��'2Z,h��K�Pκ����;�M��'�#�/E�<�$�X�,�<�x���'Z\�0-�j*fLٓ��?3����'Z�����|�>��I	�#��q�
�'" ��@O?D���
2)�?.�� 9�'���E��N��Y�'��.��
�'9���Jݜ5-,]c�k�%c՛�'�A�wkS�S�F���������'���S��ٵrm�ñLP����'C0�I�+�&���r�i������'͚EQskYr<=Q�)��w��E
�'Wڬ�Ҋ�?6gf|��^�b���2�'U�Pt&Y=>B�4{���]�\�
�'e�芧���jc֠�'��@{�z�'\��� �G��|��c�q!@�P�'�^�bL�c9ZC H�w>^��'�ޤpO�(\>h�T�]:@�p��'�Ȩ���O3T���I�)\� �'m��%�~5�v�W�,T���
�'�ܨ�3��	Jv���f�
6S�x��	�'-��a����0�kf`�:G��B�'�Ja�0�:�!Bc�?7�*)"��� t��t��,5�~�r�#�.R���"O�9�"J9qj!!�Q�7��U�&"O�p����/Ll!�Lu8F\X"O�YG��w����d��L��(:B"O"9��B<����u�cd�tS"OD��Q�Ĺ����ڴR�%Д"O��7OB�aJ0�	e]�ؒW"Of�i@��i���3���_;�ѳ�"O���m���B�`b�T�H7�$��"O$�@"�X�E�q��.2M`"O��
@
U3�������� т"O�L ���7AE~p�@瀲&�pJ�"O��a �n���QV̀%I�Dx3�"O�����:G T�b,Z9 ����"O8���hRj�LŊ�4��"O��9�J�*�2|
����Gr�)"O�D��kq�m���ll�"O�$sg��]i�j��!����"O��i'@L y�҅҆��U��q�2"O 	���ܨC=��s�+��"�+�"Of �UMҶ{�� (�闋���r"O0��/�;6��Y��+\�[2N��5"O���Q�ǺLR��;,,�!�"O�\�HR�5�"�.�C��S�"O:�P��ǲ]�LT�u��u��"O$�b㑬)��z#+�(<p�0�5"O�	�@j�@f���jŚ`�� "O̩J�ʖ�AI�<� I�d�R���"O����X$@��R%�M�q� t��"O�qRTAW$g�X`S��Qr�"OV�q��G0tJ���R1^ڽ��"OL�����(�l0p��?U���C"Od�P���*Jآ�V��#]`@{�"O.�	�F8p�h�lë@VT2"O|�&��an�r׬�UFJ"OЍ�s��3�D%�A-�y��"O�h$�@@�ހ�FBD0Gp�"O(�%�
$�p��1�ЇV�|�"OL��d��J���Yr Z+"j�}�b"OJ���1+���bg/>?X�8B"OD1W��,�wαEA:���"ON��	X�Gm<��1|i�D2`"OB��6	۱�8А��2NBƤ�G"O��R���}��1֊�(�����"O(5(���9bR iSҤT� ��ai"Ov!����EM����m�Kq8���"O^EzS�W�t;��a��[�n~��"O��@a
�2�N�	�Z'GPZ�R"O���3��8(�����QAa�l�"O� �.�S���g蟐`��m�v�'�*y�5�;r��(�v�Ǖ?����$�VN�ũݴ%������%��lph��$^�\φDJ�*V�,X��f�!�!���bÂH���?hȘrE�9!�Ė
A�X�c�Fjbf���3!�$��`��!�(�률�'�(�	�'�̸i`�I*}1���8S]���,����������c�,&E���hO>�c���a�R�H�)P�s��Ca�l��J���S�-�6Q
F̃5�>�;f�B��Gy2�+�'�����^��,2D�?H�٩���)��'whiFy�'���ǧ+��#6!J��-
�韆6��'�,S���	J>t �X �$��<cd��1d��d��pY&��.�1��Y|��1���'���yTH,BO���G�_?��-�#Bsbr��Oi�W�)��h���FB4j����6\�|9��^�/f�Dx*�� dAj�F�#@G��W�*u>!�R�$�:�Q��@�G��[�Vi����x^ݲR�x"aQu�'c>�{�̙ EZ��C�|nZa p��>!�".�S�O*�����c
d��P&�G���P�4�hO�?i��α%��-��8)�����5\O@b��r��L���Z�����G2D��N�#��M��%׀Zb-���/D�d��-�: �r��'� )���-D���v�߼<��QY�M�U�.�qCg��=E�ܴ���Hd�G����x i�KNY���D5}b��$!-h(1�=(p���A�+ ��m{���~t}��O\QO�j1��I%j��A3�A�)���Cֆ�)Y�C�	>f[|��ՊB#V�aqU�a
B�	]�,R*�m�5k2�
�]rC�ɹZEB�xv�W"뾽�I�Hc<C����v�@�E�H,"C�I>%X�s7f�x1u��d�C�	T��Z��D�f�����%,FC䉠X�LѦl,��� �'�0C�	�ip}�1G�U�̰{����B�Q%��+�R�3��MY��B䉇;������ݷ�A�c��C�I�
>� �7ť\�peK�͊=��C��*5�xى�@Ԛ���ɦ$Y�B�	#^�>	2S�MQ5�ˆ:��B��i�$��,���>p�q�Q��B�	Ng�a�VYX��r/ó9��B�	Lkf��6
��d�$5s�bB�.|PC�ɮ�<� %GJ#B���`�
f�C�ILM�4	�~�ڌ0gW�}�&C�	�I��U�/��؁ �U�y��C�	�EM�1g�t�<ʢ���C�'8t�U�S:��0R�H��GHC�ɥ�n�Sp�ۧ\QV�� ޿8�fB�ɤi>�t��AǥF=\��B�#�\B�ɉ�4ܨ3M� �m���l[�xB䉎G��ڶg�|�jA�d�W�>��C�IG�1k�4-�����~dC��
 �.�Ej
�3�e�C肌^��B�ɪ\0 ���ʈ'�����T� H�B䉖E�g�Y�h�	��<��B�	|	��J�Q1
�bA����=~B䉯1Gp�آ��dJf$�clĦ�pB�	��xċR���}�B�y'�B�>~B䉦;4��`�׺��� :)�PB�	"bd ��d�  �L���Y��nB䉛[��Z����R���"�jB�	�l<"�I�)PWX"���� %�RB䉺z���"%C�@4�DX�MӋ1FB䉊b��0Ы�G2�\��Cu�C䉃S�D�����{��)V��B䉮YA�����N� �\k�kE.&C�ɐ�!8Fnӛ9���C�.�2!��C� k�B4�s�˥P��i�"S�B䉴U�x�B*�%��8�c��[�B�/^gTI�B�2g"�p�0��4~C�V�9 EB�s��R �{�VC�I	0���Dоn�pp�7e�1�2C�ɷ4N��j�V�p)bI��&lC�	!P�$:󃃹M�H$ �A�>pZC�əj�A���a(lS�b���nC�� R�d�� *C� IS�C�[ɐC�;(:��r�@�HX2�i��C6�B䉌 ���a�j�Qu�L� ��B�)� �p9u)!,j���U�N5ZZ����"O��z���΄��F���H��Ic"OT���CW��A-H�'�xԀ�"OJ\(1��9e����,�>T�̰�"OŪ%&�����,2t���2�"O��1d�E��9C �k�Iq�"OrE03嘇x=�1;D�$.+&d�E"O�}��ǷH�~L����0wBu��"Olբ��&1�Ve� Jï!����"On��fE����U	p P��"O�]1�޼[8~�x��B�\���"OD�!3�)b�R��G�I澸1C"O2��I[�'� �� ϟuv��0p"O<��� T|��	�oT�m�)��"OȠ��"
xM��֤@Z�IIv"O�1b��B�����IYQq�$"Ora#��? �zИ�"�}*(c�"ORy�G�F�pL(����f�`M�`"O�	h�OQ�e�p�/�?\f�7"O�� ǉ!�n�C!,� Q :�b"O������u�6}h��
@��X�"O44I��"+����pJC�P,œ�"O�%�����X`���;�,��"O¥��c�9C�`$𶋈�n�6=c"Or��bߙQ�L$x˖��m`�'�.a� �ݾv���4�H�Y�����'����D Q��Ʉ � ���`�'@���b�U�LA.e!�	9I,&���'�2	TlO|��t2`h�>���'��t��H�l�@g�� ?j���']N;ǁ12Ҽq�fd
b�LX��'j1f��`��qc��WX�5Z�'S��+'���Ij!�[+�4`�'�̹ғ�Q�$Y8�.�N�<� �'U����H��B���C_K�~5��'d�B+���k!@2����'݊x��lI�y��U��(�4�J�a�'64��`_�"���c�Ő+v88�'�6-�N�1�֘CE��n(��'M�ę�����*ƍ\�*�'Z�=��K�*�ങ�	 (^'|xI	�'��ep�ȋ9$P�xuoH�JD�u	�'rt�p뗶T�nY�#*=�6��'8�XqNQ+g�]X3O7&�Db�'r(ajGp�fq�ϛ�?JR�j�'�DIbd�y/"%�fn�7���C�'g����n�!�8M�5㘌AjrDX�',���Q�U�D��H�Ԫ��3@jث�'
^�C�.B��q�D`�,0KV@�
�'R>$"CeHX	���@(�����'�e��ͷH&~�4bU�=�V���'��x!A�+|�&K�b
�q�'� ���U�R,H{�HȞfkv ��'d.աce���J,�f�ΰ\�&���'�>r���#���Q[����'�^<��ܷ*΄�C�ŋQ��MB�'Y
�À��l�48�skH�u��l2�'�L���G9mª=rs+B�s5t�ʓ�Q!��ܲ+rT�	��24���ȓ2t����۱z�vлsO��"y�ȓZ*�D��ƁE��!𔤏��؆�1��j��I-t
�˰@� !o���c�|�k�KP:h�N���L����n�<y3I$�8������<#Ǥ�_�<� �j�G
�.�~���e�Y��4RR"O���t�̩C�V,B�ŉ�E���aB"OV%��K�p�����E��dRP"Od9�b�,�q�T   ~ ir�"O>�z�)%�^}`0 G���5+"OjI��KK�(m�R�X:Q8D��"O�=�W��9 ��`0c��
W�\��"O$b��B68I[��J#hh$E��"O�0�F�8X@̱�J	~@i� "O�t;��5��ࡆ�A)9xֵQ""O������CF�%�S��?4^bI�"O.=!s�N7t
(c',��Z�>�c"O��k����:X�x�dT϶I�"Oh����1�pYX��-��XF"OF,!�͖��$xc��S�d�ʐ"O��J���+5l�)i��4�"O�Y�E��?����3n�$~��H"O�aS��"F����n�2y�`"O�K�S0UEd�a��7��d)�"O����9Y�VX�u��# ��"O�Hˑ�ZT��e���Ψy�l��"Ob�s��V�bk�(�fsh�C�"O�� g(q���X�LH~�Ґ"O��t�'C ,S�/ŝKK�@25"O����a�J��u��+�18�$�@"O�0�DD�9j�u0ӧ�=( �"OH�ը��0t>�����_|�p"Oҹ�VȤa�V�7e�5"O� ��Kۓ~5�ԋd�W/r�nex`"O6�KQ/.`��[eěl2��"O��2��
1��ujF�"���v"O��8�\� �ZLq��7 �tH"O<h�1�\Fy*���+'���"O\m���?zV�����N6��2"O�(���A�ReƇ*M��t"Ox�bR�1�ƨ���\�#� �"O4�5ǁ�*�4�%iO �T��D"Or�Pg��7��	�Q�B���C"O�)��ں#�6I����MؽD"O�|	 �X6x<��j-�Ug,0��"O8lPv` /{.<���A˽0g@	Y�"OL\Y�Dl�v���ϗ�PN�X�"O�8�����@�@%�2���?t�K#"Oݩ#OE>A\h�``��c(��0"O։���ާ�� j`a�$Y8"�"O�|r���iW�x��oJ�c�h�d"O�a٢��7P�0C����e���T"O�hs�C>By�q��Z+cn���"O��bu`�$���4�Ҕ��	9A"Oԍ�Q��K(�ّ"ݟS���1p"O�=��̀Z�Ĺ��A@�`�R�c"Ol���ےL.� � N�<�𸒢"O��0q��>ew�D���IM��"O6!���sLr���S#,�*7"O��	Ī��i��B�$^L�$��"O�i����,�5ʅBT��"O���-`z	Z��١��R4"O�	ץ��h����FO�	k��r�"OڱKckP�>�6���헉 Ϝyc"Oh}q����q!lG�F���B�"O.�$�I'k�FM��F5�� �6"O0D�P��Rn��w�ԖD��-�"O�iR�fP0
#�I�Ҡ��4A���"O���Q"���}AB�9%(*����� z-X��2*Δ�B3���%�"O|��L@$_���J2. �<��4�"O��Х�|m���Xm��xKP"O(��a��c7>�:��FPZn�#�"O$���w�z�s3K�!ll�C"O��� ��RE����;<��@"O&8k�
Z��b�K J%�0"O�`�cFقJ$�±B4l���"O�9;���3�L�""��'vBd�"O�(��`W
�^x��@�\�-A"O�x�%���t��ѨR��up��"O�;��]�*�H��j�M�0��"O�����G�?�V���3N�bq�E"OX�!�؍>�fy����Q�B�9�"O�D�T�NiSpP�&J�&,�0�"OV�(�   �d   
  |  �"  q-  �6  �A  �J  AU  `  �j  �r  y  `  ��  ��  :�  ��  Ҟ  �  X�  ��  2�  b�  ��   `� u�	����Zv)C�'ll\�0�Jz+��D������b���$�y���y�FJ%L+�:B�o��e(s��!,y(��b��v&���@<!�G��뎈
$UD��L��"��J�+�4���ԌUe1jQ��1�\�`�.{�Ht�Db��mH�<{���baz쯻Q>d)�'�?Y�*\�1^\�"�pھ�	O�CG ���hZ�&I:M���ݵr{D7��s$�$�O���O��D�a�X�	��M.���iH0{��d�O�m�/�¤�'�jH�����'���@�<��p1��L�$�c �[8�B�'?�7��O ��?!��ٺ�w@@�p���'X$aJ��Y3�Ȭ(��fE�=Y� L�i���'��e�t剽v�p$���æSM��"S���7�x����D}"5O�㟈"�X)*R`�Pa��<Q��i�^�y��P!B�<��	RĘ޴�?���?��������l��Ѣ眺뺥���M�,�'�ON�nZ�?i�4yʛ6�'`@7m�!�:ml?h���a	�\����cFd�LhGKȔ2S`!���$�fy�!�H�w'6��5DJ)���a�i��,9L����l�4{^���4�����d/��M�3�������4����O��S#�4��Dc�9!��Q5m�=�|��@�$ä7-P�|��,J�G�/#��Qc�4��dj��tw��n9�M�i�Ҵ�VM�*r��+����jڸ=�)2om�iѲڡu��6M����[۴2ʪh��:]EjUS��'uh�y���	7L��â@�3��Ha�#\�w�"����(;/�5�E�i$r6�����p�Ε!o�e����x:|����)��<[üPɖJ	�'r��:���M˲f�.V�L1a򤏳*�y�'EӐ�?a��$�C�l
`�H�\}����1J���P� @2���'A��O��A�g!��g�P�L��ֵj�v��UKڼ{���H�Ww�X�\�I����'~��Q35헼G�P����M��
��\�;��͠F��8����0<A�LP�����A�oW4e)�#Épk��G��� ���!�aڌx\����CԬI Q�0�� k����\٦�+Of�!`L�2\l�@�ݮP�H$���'�r�'H�'��'b�'��O2j��aS�ڲ Z�4�	R.1��2�l�,H��"P�g��a��*Ɨݔm�p�Z�����MWG�3tڛ��'��'>�ĩ_e�hՆu��Ũ��}�X���o�?�"�'����ċ��/�Ѻ�L�A�2Ő�[>�O���C�-��k�ըtY�m���,;�O�.-e�P��ZEah���Ӿ �j�g��4�i�i��+�m[fi��A�4F����4���^��K��Iw>��@ۉ)�U�%��>}�La��e5<O�#<��Ɖ.&X�%��M�4��*�a�'�f7�����|��Q�8��4�p�
�j�|@����	uyM�n��'���'��	���-�U��F񴠹���/�������l�:�i�iG�ES����.w�4�Oi��$�pyf�C�P�lq��I:�)r��
�SCx|r����MK��2UI�Yy������*�T�`d7�D�A��B��H��%�V|C�)d�r�'X(�8����Ο�'ɮIT�E�e����\�_�� �'7RY�(��L�g��Ã�Niba
�#<*�gٴO0�;�M��ibɧ�$�O��I6_��A)vϤb�qf���鹢������O �d�<�,��擅K�N|3#��*pȊXPU�X�cs� 6��.	b�k��c,R��ɾ?:����A�'E8��Cߎe$|6�Ɯ2�*x� ���jW>i�D˦Pf]�_ob�0��ɵ�¨!�%U�	��8��T�4a��$�ۦ�[��$?��7ic6�أB�0%��с!*\�*}��ʟ4��^����I��c�$��`���M�E4����y�ܴ���4&�8�'����^�t��i�=k2�JM�Q�2�'�Bٓq�'�R�'����.P�"	ք��lAe� �N-�ʈSu�O�ijN���8�ax�bP�Q���ph�)of.�VO�l�QH!JH$�����?z�H0U�-ф�3҇�E�hC���I��M� �i�N�`#�qŋC�p�Z(��F����	埸�	ş<��3��]Q%�3d��$�0�"V���D[�uʢ�#"�q�%�eF���&�0�MC/O�q���4;���OʧH��x��N*j�0�`��m��N*1�t� ���?i�i�8���[ �R*� A�f��2����X�d(�35B��	/5�� ߍ'��ɂi()�F$/*�xW����4z��EDCLh{�'b�����	�f��[P�R��'��������3�)5�ӝZ��%풕P�2����)tx�OV��#��f̓	��� �Ҕ�/m��bЈ�<qEl�^?��4�?Y��i��7��O�n�۟����@�jd[��$ ���腀�M����d�,9`����O&�D�O��R\-Z��V/#�����j�=�t�ab�*cټE;�i��y�$��S����'o�m뒪R��Lqv��"����>�jux��+[T��1��1�z�]>��&��-n���/2G*���	ʹ1�!���<@۲�nZ+jX�Ic/\��'��O&���O�a��i� KZ�MҘM!6`�&@�O����OJ�$�O �?�'�4�pЫ���V@:����~��s.O2�nڻ�M��7���'K�d�O����:�Fݏ"[��sb�Z#z(���*m���I��I��"�����On�䁘F�QUH��ZeDL�/7�V5��Ԭh��\���C�*ZB�'J"��MY�
x"кp�
V�aփA�`��A���B=�n8a%�+R=�t"ժT�8_�P�2�|�N&�AD������K����#*5�?��(�32ӛ&�'s�	�u�T���'fx)٦ �sz��∁?�`К���ɽr�qOx6����t�,Q����
��`�Q9_'*��d�<!��-�F�'-�	(2Kܵ�ش�?1�������A�a�n���V�8XI����?�f��	�?���?��9\����a��l��٥���� �̑6`p��@%�gNX�E�Diw4�p���p�X��CGܟ^-�X�F�Ț[0���W�0�dp
EǗ(Lx��im��T�i�m�J>��A��̩�4�I�9��UY�gݡ)� ك��,	�b�O�=ьy���W>J��7A.=���F����'jў操�MKӌG�6Y����*k���Z��מiܛV�lA�(��M������|��|�29���+:���RcM�:�  ���?)3����� J���Թid��5��!�=l4��O�� �4�j�d;?Q4o�=S���JD�6��p�"��Q��!H`��b�|��m5��wlL�*��0�U>k�X�
V:���M���S�|҅gݦ"��0�@��=6W��a c�Ɵ0�?Q��iӳz�>q���W�0����vgR�7o��daӎ�n��D��4�y�bł��!;��`�㥌5j��ֲi,b�'>��Ų �|Qs0�'���'{��fU��'�-;��_|� 1�iG -��n�ʼbD�O}��''�D��(��D팤H���
`���H���r��5��	� ��Ǝ	@#J�Od��R���y�Ϻp�p牆�f�ˤ'��Bg��������D�t�$*�<Q�(X���K]��I�7S��R���?�,OJ���O4�Ă�]�Lb����9 Q0"�E�-����u���m����M���D�O��i�O��pDI��揑:�T�X�A�?��5��.��� ����?����?1�������O���.oK��`�a����%e$S� �7�
��`ԡ�r��,#���>0l��"l'ʓ���YE�յ,x�,  ��3[��3���V%��z¢K lR�cƦAW�� ���Xh�pK>��Q�]�bqz���	��� 5#
�	ň9�	��Mk��_�'z� ����>`���;�\y���'R0�3�B�kjj�iG�P�}�H>���i�U���7���M�ϟ�)SХ՘vFP����m���j7�'L���|���|��`���8�E��*HÚ��Dj���0RB�^"f�M;�F��?Et����I���b��֩K�`(�!�hm�W�	Hv�A��� f��BUI����7��(*ܚ�%�"����ܦ��(O`Ik�g�FѩI�)%z���'�d-�O��u�
 4�R4;�cT�P��e�'\�}�Cc�0A��e�C>����x�VǦŖ'�5c`�z�d�OZ�',$nD����ډPu+ƿ^ZB�E	?�*�����?a� Ik�Q�Ь�-)�0Qy��"b5��)���I�L��@!�k�D������%Eb�cBP�LʂDK.P�Î�Ő�x7�ȝ%���O�\ ���k4č����=,=h���Ob���'�|6���O�i�11jL�"�>TҼ�R�>k�r�)�"-;%c�e��0�h�!-�,�rÓ�M��i�1O~���h�.�d���S�(��5���D�OX�$��s�ޱ��C�Ot���O��dn�=Q�/��Zj~d���[�0~а�mG
��ʦ�?_�Vq�A��{��b>�p���L����/F����a� 6p �{�#�:>���0C�
H̡�`�8'����܉)P�'(��Lq`�JԼs�B�>���[F�˚
��X8��M�W�HX$��O��I)&�da�� v��<�f����Y����a(��/�H�>"q!O�Ov<��	ޟ�p��4��d�<ѳ��%i��Ѳ$��Ygf����.�?�����?	���?�m����O�D�O`9rn�0AeP��l��Jmz���K�>�:G�H�+�*x�D`�Sx��SD燯2)��[�ċb��eJ�Oٙ����C����,)�\� ��Q�#	3 H\|K�$� $<D��R�cPn�!N7�ΌP�'	�� %�Ӻ��rAK���t�EB4m될�%#@"�'�|[��>%y�J�;y�uf�Ǉ�p���<y�a����'剢L�xߴ�?�'l�L��@�"nP��'�7"@�(R�����O��d}>�J�BD�\�I��D��-lZ3P2�9BΖ0g�D��ƛj�dt��ɀF�^���#^���P�F��|�H���![�y{�Ř�h14�A�D8�����ׯ^*qO��@1�'.J7�Dy�bJ�E ��¦�WV������0>��B*a'��k�b� Fq��2�Fy��'�6�ݸO�Z�1%
O�@����!~�4�n�Oy���9�7��O���|�ҏ��<)%iütL01ŭ�+}sf�C��8�?A��[��m�d�Ⱦ��$�Ol�g�DD��	�'Jő8��d*%w��>UhW��#A<`AW�̭�H��Cn��m}���"�( z@�'��$`�vU��(�'���¤6�.��֮�:-�����,��'Cў�O(��)��E��y�G����Ë�DC��ݴOWH�WG
Q��-�T�A#v���`�i�2�'�r�I�k�X���'4B�'b0��tb@��1r��F��fL�}�0)�;1X�0��ہ=	��"<���?�A��x���
�<�&h� U�� NUj*T�c�͞_�
�r &�Z���B�3���7�� ��y�Gb�T)�灤��#���|�F��<Y�g�۟|�Sw�L>!&��g��U������p��?����ӳL`>a0���"��	1H�8�hH�	ğ<��4b�v�|�Ou�D]��kD�H_����'S ��!jd��
^CDXb3�ޟ��I������uG�'�R:�ށ�R&�SF���� [����_�n�J�1��&W�⵱�j�"� �?���_�? l���k�0y�L,J��R�kn�; �Ś�X:&OD�D��m� 8:p����8S���O� �m��4g����Ɨ��� !��6n��'����4§;N��恷9B�QjV)A����ȓx~Le1����z\X�U�#y�<�&��i�4�?A/O�r!�Ӧ���h0eČ6҈�Qӎ[bu��2�����	�Q�i�	۟(Χ�P��'QU�%�a+�;d'$A쎽>~�Q�dJK��`� '����'*ʓ)z4P!b�4ke����9��+�hK;?1��׫��f6�Yɂ˒!�d����FɨM>������$�M>���_�7"h�Ș�9�B<��H�<-}��@�P��JȤ�(��F�m�N��D{�OX��D̼:i⫘&���fBW�N��'��%Y�Cv�d��O��'e��l���'X��*8��|m�69�����?Y����c� ��`/�ZCXt�v�i*��\���^�~,��c@u����R�[<�ɓ�Թ�p��-;ߪHj����&d(�.^>�zػBܟL=�jޟIw�\�e�7V�D�3֔���R#�O��lZ��ħ��O�@�s���
4��|��$)sw�UQM>���䓦?�����S9k�|��s%�:%�,�Bb�?�џl
��MI>u ٨�,h1Fc�0
��Z�/K=7���'�B�'=ܤ����S,b�'t��'f�����I �/h��D�b�͖�1O@��!�')q���YA���A�F��y�$�0=�5�P�\��@I��ԍS�Hq{Eb���P�Hi��}�g�=�8���-��T�(��1)�1�Շ���Y�	W�A���*�H\��k�O��Gz�O��'�v<��&��$v���ilMR���8V���s��ޟ�I���	����OX�D��n� ㅤԑ+�(�i�(�QON��C$_(g,
Q ��L�&�^���:PE�}�2�p|��ƢU�#"�A�B1焔f ʠ_,�E�P吸��rA��YuqOl��� ޠ�L#��ڳ&�+!� ��t�\ImƟȕ'"�'u�?U���V�'_�4
@#B�q��u�Fi>D��x���;}I�|�"�%EF���>�D�ڦ�ڴ���27�D�m��T�ɟ3�D9����/���E/W�NU����0����̟��I�|�3/ڟ��<!6�DT�U��USB� �f��c�.6K��=0��F=Ry��:�@��@1v=��I�F7���E�3�z�Pl���`����C�ɺ%���@��*VB�`3, �70���$ş���2(�Р��%mP�US$#5��DǢ��z�F�$�Ojʧ4�(���V5 P&�=z�ND�'e	�qx����?!�I?JRJi�!�zϼ�)� ʠFǒD"�����)S����A @�b�<��LT�&����)	c/�@�#3�*jTڸ�W�0��I�F���?"���-7�(P�"��D�bmЇn9?i������@H>E�����c�h�I��C>7�\�؄"�y�C�i`�3W�3ݢE#d U��hO��Ęe�'9����N�P3���W �XRj~�����O0�d�O>�!�O����O�dw��2P�'�D��į�E����$,89��qo��\��nهM�HŖ�(O�Y���D,Wd�Zd��ra�:��8(>�ʓ�5�- f�g�j$4ḃ�ɟ~)�8Y"�b�H��	 ���	(f��H����?�v0|���d:dI��(ʬ��*OD���OV���O���=�j�$�OB%:�N .�` �`P�U�N X��ĕh�H���O���'&�A�d�')�I��=��?	��0ӊ�~��4!o[�8���I̟��Iǟ��������|"��V�;A�����m��d�Q���5��$��.r8��0h��FȊ�Xm�#͇W<�4385#@��;/��IxFD�+랄�I���?�2I�D�<%W�Y>x��7�͸�yr%��3Ĉ���<
%��aP���uڛ��|"%ݐ�"�'�RbH%/��qa`��ZgZPɦ�%��'�����'0�7�4� ��'m1O���v��'7@�P�͍BkS�'��	 ���V6a�V	���X v�H Pq�ax�H0�?A��|�G�,k���0r'�1)�N��y�⒘6j��f��q@�{7,�9��?%�'�����,�$�.��)�_x\d�J>iCa�^y���'��P>	��ןԪǢ�����YU,�l4�Z B�Пx��v�J���h�S�L��r�i	�z!������24ڐ�$?9��Gb�����J��n`Ui��(�2L����ܮ��?���|��[�l00r��,|� �vD��?!��W�d�Zv���M�&lj&�
�"�P�'O�#=���R�����6?�����+��?a���?��v8��w�Ғ�?���?����y�ĝ0W�ykr��=оʵH� A-��)`cЭ ��,z�ȱ���d��a����$Hx�$���k܎c�ڨ[d~��6��(x��q��_�˾|�M5FUΑ�{�? �����.e�L���H�'~���'y�I�$N��d�O��=Y��F�����eP-E�5�7�yb�;��Wl�BmD��VfM�?!��:���S��'��X"�$Ј��(�@W�
�"$ ���(KOT��@�'Wr�'z2p�a��֟��'l��� ��(�X�ҷ�B�C$LE�R(W�6Z53�)�N��q�[��r�!P�<ʓ!Z�*���3>H���Į@	�D�㣎7&�t�sF@�|��x��į�MSU���MX��2�D�"j��89҆s�$�� +�L9��'U|��$��;��kQ�ŇUl�q��V6&��{����B(�2C.d��0�V�2��'�f6M<��	7��O�reY�Yu���J�#� ,�.Э-�R�'&�4"�'�?�T�P�d0�̬�h���J19��	1rH��倀Nx���b�(c�	�(O:�uf^`h9�KBY�^���fA;<��X�慞�ca��$f��I���C�@��M3��A{�� }�����O4�w��r��� A��%�hm��$�����-+�lx8�N�.�������Ipv��G{�OĐ���v���"}R*=B��Z�\cc`ů�MK���?))��0Z���O�qQ�BG μ�4 �47��A��!�O����yoZL0��yO٢2fwt< �7��� ���';��9I
Gfȸ�JaO�j)Tq��O̀���/��(r�k�+̞e�P�^]>U�H?1zS'O,%�yYvC�;��u�8?���ɟX0H>E���.a�JL�A�½wo�� �c��yb�3��жN�r����`$$Fҍ9ڧM�H	觤�;)�m��K;u�T ��4�?����?��J@q_��r���?����?q�wΰa1`/��x��yF �6+�0-3�
��1���Dj� S,B�2r.S���	~>yfK�#{��DN�t3�Tj�o�?XÔ���$�]X(��e����|"�J�
]P͠w󩑣
)�q��'���0�	�7���j�P�` �0�|��P��?ُ��yщb�"A�!�&�T�wi��yr"�?a�@�U W#�5�%�
2��ċ~�����|I��3A�}�E��w��Tx�B$r~H�2�¯_���'�"�'�ם럄���|�ӫƚ� DKp�G�u�v�ɿ+��x Bω�7g�� W��X�tX�!ʌ��@�<QC��6lJ�
<1�����aD:(�f�+:TB �".��\a��
�<Y`���r�	�Š�-\�a�r�C�[h2�I��?��΂8G�m)E��(�8���	M�<0��g��x�R䉶X|A���I	�M�N>�3N�N�S󟀃���<�R0��� �#�0ˁO����	
)p�I�p�'>��$�s$��+��Bi���M��o����y@@H9ڤ��U�_��M{��0ړk�Ԅ���^�F@�'	[�M�01�"�^�f[nI+nY��c�ɗ%��=P�e�K�'��l{��?q�O���1�֕t䄩P�?���k֘|2�'MFq�"M;���7B� E�H�8�,�2��qA�mR2���{����dH��?�/O�%!�/�O�$�O�':ɂ(��yE(������
v�%�' X�=�dy���?)`�V/Mm^���N�$�Q���Į9n�:�������?pn���J=��}�ҋ��Ql���;NM�#G�,G�P�e��?�V-�C�U�<z��ݟ�}1U�A־�"�K�9kY�Y��`+E��O��D*ڧ�y2��\��H���&S+����#
��y�Z�"vD(Z���bW�u�DE:��Ot%F�d�X=���6��Y����%KfW��'���'-^QA��҄���'���'O��M�P��5�s,�5Hϊ\��P�bK{}RǸ�| r���ybF<(���t�ӑd`��-:U0 ��o�>1҅?[��|�<	���?3����D %��!������0�'M��{��?����߮b(����<.@$�P��.��C�I�,ߌ!I���{w�t��f�'2�"=�'�?i/O,��I��[B�\�DZnNzD�Uƚ�9�����O����O���ú����?y�O} d{G���x(�DEd�u�Ĭ�tȢ�B��I6�TA�@V
~�џl����l���d &�X`�҈�N ��)�-ؼ�C�J/8�=)qI(�#w2aۃj�/MƢ$Q�.̐# (�����	��?	����������:�Y�4 ���!�$��ԠR���w�^��/�WK�'2�6��O�ʓf����tǜ�/\���'�J��D��CГ�?q*O�D�OB���QCY�'e�45>yqg�	ğ���́�l��ꂯ͖n�1��'O4ؒ�"�lz|3Q�]qP �D�:/���Bh�_W�X��B,?>ax���?)���\��0��b��B�L�<�'��|�L��jQ���N���gFq���8�6Qe0�]w:|�Z���%9�0��I@y��%F��)R-�N�C!g2(˷��8�MJS!R�U�@�$�Oډ�PI�5�-Y�9>.��)§7��X�2/ �A��A��e��7��'��a�3�ƀx	�2���|>�>)*'�Uc �C�A*��*��3?���ʟp�	k�O��� ]c�E
�ʰi0/4LMx(�V"O�5����J�G�V	{D���I9�h�"H�D�k�\��0�޹gC4�
�'��K��4�Q�H����F�1HR鞴PBp;�7D��"�GB�r�t��	>!T[W�6D����0P�6�����B��!eO1D�T㗫�L'|:S�щR?0�[7�.D�P�Ѣ�<z�吔���� � D��� ,Vr`�c�UpE�<1v�CD8� 9��Ƶ9�$Q`cX�CRtIt*O`�K�B,U�*)�P���8��8�"O�@�f���Xd�0iS�TZ�Q�G"O@x�,S+]̰�ض�N8qIԔ�D"Of�0���9���eM��"�'�&��'/&t�ǿ9s�1顮�,o�H��'��e9�N�yr~�X��$D���'ힴ�V.ê[����J�
h� �	�'<Q����;#�|q4�L aWJ� 
�'���DO'u���SN9c���2�'����� �:3�8�� 	c���i��D��Q?��B@�3��zDI�-`%��(9D��b�@QZ��#�(f�D�ǭ7D����أ�Uf�ϜQ$�meAؤ�yr#�JW�-�
w�b	
�˟�yr�׌a��c	�*A��3��0�y��	�k��GK�}�'"���?)7��O����4 @a".Q�� �M�E��"5D� �%�%z�, ���ug����m?D��("��Hk2͢�E\
+����?D���q����˃e"�I�e��#d�C�IUW���āɠ���lX	y��C�	�J�jU9"��&bP����;� ��cN֪\��b�Iʛi
"L�D��<L�l��/��^����� C�Ew���*D?t8Qꀖ).a	FB@����,�X�I՟D�	9lP���,�?	��h�F�7z�52�E/R�|}�F*]� A�x��G�Qc0���dR6e6b)K��L�nAP�Ř :�ZE���<"U��a|I��8d&	�i��*��D�Ә|�	�
�?1���OG� h�ɣQ pi��׍@>��)OB����@��C��@�#o��b ̣)��'gў�S�����n�0�	aKх"hl%3t/����)|����������d�D�L2@��'�XH᫐��a)�D��v��p�E�'������2$8�)� ,l��$�~Z��l�?�PIQd�O��:q�V���yRq�$��Ҭ5Yt��Xs�'�P���l¹���õW>)�D#I$U<��H��
.|���~�XJ�C�O���1?%?��'D�|�S�yS��!v���Zc��
�'V�5腋P�"�8�Y%V�Z��m���'R#=�'^)�pHγz�&��E�5$D4���?���d���#�L�"�?!���?������r�`ೈ�<�~,��%�KEn�J6�E	��ʯ]2α�7�:��)2�	�/҅3���^��e Gf8�e�q�� QsJ��^H�L���E�DB�5���ĕ��`�;=�0$��9i�2%0�����k��TӖ)�Op�%ړ�y2��E�NU��M
*S��:��;��x2�JJa��'�'Ԡ��a��:$RK+��|����򄞇u�����N�O�č��ڿi����[������'��'���Ov��'����nҜXȄ�H!%�|�`�H�j��S���F���K�"@��$+��K/��b�L��\+}�Ab���$J�C첍z��TG���	ABTr7�֨o��K>I���� �֫Ϸi���˖F.��|1������G{��_�A��f�fUt �F�??���d?7��M��Dq��c��'��7�O�˓/_�_?5���|�������V��E'�0:�0�ɯMJ,���럌�	S�tX�G�0��l��!ں�������F҇"�B�r�� �
�S��TP���u����T
՗U��@t(�:&�5���(�f5���čs4�ȳ�4K�V)�shV��d%�4�s�O���<�S�:Y����@�hh8ӡ�.	���0?QP�DH0i:�G�-����{�IA����O�<i&.�+�*!��+�t쥳hS}y��_y^��'��R>I�F^����	]Rz�QnY9O4}�����2�~1�7FW<|;�X��ɒo3���"؟<c>ag�)�h�9w'ߡ{�2�u�}��+㯛�DW,��f�͋m�L��+�6��A@�!߽A�촔O�v(�q��}����.�_H)�'�����?��O�O/�)� fx ��,Z|x�-�0l���kd"OZ4��K >�8[g���V�<
4�d�O�IGz�O�~�s6���B؀(*�MɡG���q �'���'���#T�A�2�'���'��4�'����rcة`���L$.���T��<Lk��עp��G�3n��S4��'�6�����%)EHȑ!���V�#��N�	9l�۱���������5O��S�%��	��ήE����I�(�K�G�-����ʈ.c��s4Z����pG{�=OVr JF��qCCGA
!�<iIAOP!�".��;�1Sȋ�������OLGz�O�2T��2�\0c��!�c�&0ֲ�"_�䭘5&؟��	Ο$���?����`�'/�y{����f�p����.b��Q�+G�[Zz����f�ڼP�j��w�ɹ~�˄�ȩ�P����&zQ������>ĺ��.Z�����[��Ă��C�D2�%�ؚ���O�2�Ro�T��eP�VȠ�r���O�=���O'�rD�##MWR`�@�mڨu��y��I�]䌸���m��xBB��0u
����'��S%d(0ܴ�?1������U Y*���	�)�~���P��?q2�Ґ�?����?Y� X�?эy�O^�K��ȃ3��I���v�����d�F?�ɠ��"^(��θT�9hw�)�>t�����O���ƊG0<����8q�����'9p<:e�@�4Z��R���k�8�x�O��=�O(�ʓ8�ֈ����t�\���V�>1�t�'��'��'�rQ>��O��Z�l�8P~�J��ϐQ4A�-O��R��p�'K�i��X�O���ƁE?q1°B$��F�Ww�'پy�	L�d(݌@ V�U�̾M���8��߷D�H6��OԕѷA{���H�O�����������H�*3�����͠ ����D/�\5lП�4�MП�ΓeQ���]����0�Q)���;�����Ț1��ە�?�����)��'����O"��~�D��P�`N�0`�4qh`��St�hN��*�$�O��r���O� �I0c���s���/�y"����I�[�n���P�B2��<�?��V� ��0�'�.�O��$��4��Å9;
��"�O�L�& ��-�4D�l1�	�(���OL �O��	H���s�n1�s�@�M�n| 2�P���O�r9�)l��<�f�����?����v���'����2H
<
!k��^=�$�#G,��0O�P��'j�`����<a5d
����4�UIv�ϗ�jX6O4Pζh��b��v��O⽃��'���<3���?��C�4�+���]Ӿ���(�:ڍAF$v��`0P�w�8��Ζ�!ߴ���Z��Ҳ"��D�R��E��aà8���KS*qp����>766�N���nZ��B�4�TX?%��W	����5C�5Qr���Cؤ0�'x�$��ͧ*�$iA�"͈�F���4�?a,O
�d�O0�D�O��$�Ot�$�0ж�җ���"q@��Fm�M�@�m�����By�Q�|�	ҟ��Iß`;E��0���`����"�ǋ�M���?���?�����4�N���ON�)6.�G�P��P����h�1-��IƟH�	ʟ ����'	��O��i�MM�46٦��,`}�Z����	Uy���Z�Va�+P�d;P�J�'K�m�.#?������O��$֪<�F�y4��=���R���}���'��ky"�'���p�ɏD!��
ӏZ��:6
Յ�!�E- �|�)��µn�򑩑H!�!�D��"$b�Cc�jt�\���T�)!�M����[����q_��Xb�8!&!�ĝ>>'2��p
ۚz\��`���>�!�(2�&��@�9u@l�2�I�V��O�сA.��m�A)D�0K�^����Y�<]��� ����� B$u�e�gLC%Oo�{3ڜw�"��ؓJ���V"�(�6�(uEɲ;-
c�h���EL̼��
9⠰c��!�	�(�޴[@I�k� Y��
8��+�oO����F]�B,�4�E�	�;O��K����G�����MU��@��ԕس�	��a���c$�-���R�0uT�y�Y�r�D(�mV2L��8�t��$���y��M�|�FYK�쏆D� H3�B�>&4�y$h۫y����,Q����s�i[4Łg��O�:I�B͌�y%Z�a��O
��Q%���T`H�u�d�z����QK�NKX�r���hCB��C2Bдy�%� �D∠^,PR2j̨d��yO)���%� ��*�G�2ԌHCo�4j������ējД��	���S�'L�nt�r��(�Ĵ*5d�1gz洆�C�2�;�ώ/S5R�*'��H�2��i>H��
��La+��ceb!��"E%>x��4�?����?�%KҪ����?A��?��(>���c�ŶX�$�P��)v�Z��m����c�E?<M�-��U���O"B-C�i���Bb�-!_�PrT�S,*\�A��A�B֔;Q���u[��A�/rs�yB凷1�ӆA� i��w�����3
�����4�*�pB��H�ɣ6�&���xңY�I��q��6;��!�,���y2� [����$��+�R؉��6�~B�'�#=�'��!���2��<\UBer��;r���R�P /�<�E�'[��'%2�t�}�Iԟ(ΧaN�{tK:r\����Ő!��Q���4s�lTbK��QQ}'X�z4
+�d�� h̘�B�����ln^����]28`q��ͺ�~�ɅA	�M�2��ܦ�#@�(��Z���'%�}��IA�X@ �C��'����DU�,�6C�aX��$Z7?��|�x�ht��M�U]�۱��ڸ',6�0���YT]�Oߛf���=q�̛���P��eC�M�V֞���O=
���O���e>����ܸf��BṔ�a���I0��I��,���>IT�M�e��Y�LE��N|����T' 6ٺ��"7.��%����<��@�ͅ#v�V��A��?�:��0�O}��'�<����?!�O���U�RAlU���޺"Ƹ%����O����3j�R�!�
���� +�]mQ�PE{�O0���	�cQ���e���m @�jb���9��T��CBʍ�M����?!,���He�r��(,�	]���Ӯ��T�g�]ß��>�� �	E�S�,O*�+R���Y���m��g6���xB���O���"�m҄L���Y�͜�C�ˆ��6��A�I���S�V��hڀ�� �p="�h/��ȓ.hX(�$@"MCT �$���jY☄�I,�(Op�ɔ�O24���24
 :*Ti�$ܟ����ɫZ!p�b����	�����A�9aSN@�7��'x6�aYY��i��	�8�"4a6�� ,̠#4�K�$��c�P���%,O�q����S�^Dr�EW�$T�3�-Ѻ�� T��)�3�D�.Q���1b�; b]�v�@x!�YR���ʖ��m�u��ьeu�-$���g�I(v�����)գy�2ćW*!tƄ: דvW�(����?	���?����?�����T���m²�z҅T�"ظ˘!=����'�l|:� `"TѠ+���(Л �˼�xr.��J��4�ㆁ	Y��Y���27`Ț��x}�~R��r��xrVIW�i��Y����yb�Ks�L1C/]16512*B��'~v7"��K�Z4��D�O�6����+��<b@x�Ab�#L�PP����<h�Dş�	�|4��ڟP$�@������'�6Bp{�n-,OB�q���)��\�c���h@�5 	jIay�G@�?�Қ>a��	'�Fa"�/:ب%�0��G�<EIoт����,
X�=�(Pi(<Y�Fk�>��bK�$%��8���vL0�N>�"E6�?����?A(�":�{�"��4��t��@�I�q/���'/ݟ�Ɏg���	Z�S�,O�y��_�\ar���#�\�՜x���$�O���h�2n�iŊV�B�1�~L��xb-���?ٔ�|���I��)��U�"�/7m,݂7 <�y��9`����!L�qr�ˊ�p<a��	�9�4�aC�Q�]S� �C'��@��ifr�'��O���{s�'��'��;rt�P"�<������څ1��1�D��ayr��4��$��y�`���iY���'���{�#���)�?1Rm����bX�Ӱ�#�D�b��L<�@�B��qb m[= �Q�c��<��7o��U*�훻
�� �_�H�����x��I�2�j�l���r�le9Pa۟.i��@ �J9KH���O����OV����?y������:P?�,��$[d��15���xr��Q�yئ�/8l��xQNʐy�l:�'�5`�H�,y��Q@E4U�,�P�NA�?��'@���g ��r5���BK�=���'�j @��R
�ޥAQ,�e�Ĵ0�{b�}�ƒO���O���a�L��O'pw��J�D`ܔ���ɟ4�	 �Bx����ͧS���G�IX�����	�P�s�͉h������rw�O:dsFQ�1r�� ���B�J�K�ayb�F.�?�b�>����B)�$���f'��b��y�<��N~V&M�g('xi<%!FLu(<����oK���g$͆(�٢��7g֜i�N>y�� (hכF�'�"Q>r1>UoZ�~�2��W�ǝg�	���e�"D���?� ���?Y�y*��	**5�Eɨ~��ݻ�K�+�O^}�4�)�So`������!���$�ZF�O�4	��'���O��������r����#��a��D��"O�����Z�{y4���"��-��|���'��<ك���2�F�SV.rr��� �5\z7m�O���O�0
��T�V`d���O$��O��طn�d���p�z���K ʈc��z5d',O<!X��Z�9���UL̀I��5����&P)ay
� `��bXZغh#��P��H������P�)�3��o��d�p_
���1��,6Z!�dʱ_gd]��O:.-��+�b�������S}�	4u��]����. �< �F_4�PA�s�%bf�
��?I���?�����D�OR������1	U��ҭY �8^�h ���0�䐲�+~�`�EbN�7�I�E�<72B��*|׾�J+����IA�6����v-�OBD����D�W�Ѧ&�^]hb�L)27\C�I�kj!R�Aʣc\txitL@0$0���ٴ��X�.�p��iC�i�@��`B�}9� A���t�C�I�O$�$P�-���O��S�JU���0�Ď�р��gD���yʷ�
�ay���'B��gǀ�b"�E����X˓6�2\�I���c���{���~P�`ᆵ_�B�I�)>�1��Z�6r����C�=}pB�	�`���H$+����ha��/��m�bJ��1x�`5��4�?������\�F6mW�V���eT�-�IY�
v}��ԟd��(�����<���@"s��(���&V�2mPB��&��'������i��xA읡fmɷC�B

��'���D2ɧ�O�l�AcG�0f!�jV�ئu
 :�'A�u[Є�i0�كꘌEvlB	Ǔ9cQ��0Un�?$�89ӣX)7�x��\�f�'_b�'$�ۡ��}7��'dB󧿃��'z�2�k�,je�lx�C!X��2'�4޺L�`��A+�����A_t���N0<��a�'D���Cn\i���7C��׎�8wȼ�P����́*IʧXW�)pE?�uBc� �� �n��E��OD�w�����l�L���(4�U�N�$]����d���p)���:7"Weڈ}���?q��i>�$� ��@ҷ�9+V.s夠���Sx@̫����?���?�����O��v>�xrn�/���0T&�:N8s2"�!M�C��������8��a�721��r�4����hN*�y���w7�ŀA�$U�����\����JR�ka�ܽhP2D2׃.D�����I&e�m"3�X,�y&((�I��MsN>�瀘dқF�'l���^�0P@ ��7,�H���Ș1���O�Y8E��O���r>M9�瑅e�!Óe��-X�-�(�3�X��'�"b����a�ҚD����
[�M�Q��l�"T�p\����r��Ӭ��Rm�uO���F� �+���X�o�Q�p�6��OV��O��f��ܺ0���4i �"O�y���V(`�X��N�"�t
OB���!Y�eb�`�7���/ʿQ?��O�qj�������D�O�lp�Q�i�haR��?�d�B����t���O��DĹ|��ҍ
1@B��1(���<3 a�(�v����8T�
5�B��(ޯMIz�'����m]�h�Llc�eV�%�$J��3K��a�V/I3Lbr�F� F�*q�]�xZ�Ct�%��3� ��I���S�1�pH�&�&$�FT���Q{z��? A��)�������2�����i>M���DV;�)C"���I�9�H0o�T��ߴ�?����?y����8->52��?q���?�ݻ8!څ���T�	cD�H��űJȜ=�p�Y���� �Ԙ��GJ�;��O��r� j�ɀi	��A׉}��+���t���%��"uIT@�=@���c�̧|Z�40�>�݀"{��#`D�r������	'<h�����n�O"�$B4B2�r� 8f���C�X8[�!��W�BG�*��)_whQ�DZ1l�-A����֟x�'I��P��Ϭ�>m��](��h9�D'n�܄9QO�O���O�D������?�O�~[��/���sӉ@1a�DbbM�-2����I� �Ԕ��A��џT��;�dɱ��`�е���[*v=���.Uv��yE��gY|c�%� >��Q�R��Пv��		�	##�(�r'��t�>@k��'&��'��O�b?}���#����@�Xi�K"�5D��Bˋ�Xs�F�w�9ё'�I��M�����$f[�mZ̟�mZ�:�D(�"�� Cs��S5�N"E`D���?ѣR��?���T.���e{V�ʶrl���"i��q����dRK	^Pq�gJ�\�Rt��?#�DyBf�y	��	�a�>(}�p{��E���е.@�$<��z���\0g��g�ܜH�50&�'�Ԝx��i,�B�fUY��AƂ�����
H8\���eD���'��<z�p�-L91HFy��i>�*���E�*LfJ�|�֌� �(J�%�H+w-��M���?I*��e
n�L{``�m� S���	d|A��@@��,�	���� ��h+��B�͂Y�``+P�.=�E�O
٠$+Բp����sꏬ,?�IH<�aa�Y->P���)��Su�R��u�`���u�g�9�u'N1iq�R�#�P��B�	,-F����J�)�3� �-��@�-M{�=�N��c`"O@@c�Σ>�P��'N�[l 	�/ F���G0�]���2ī���+�b�%s�=���l�l���O���G�~���22��O@���O^��w$��[���$[g��k�	ջ	OȭD`ŧu,R��vdң#�5� ��@J�ʧ�����@+ޑ�I�$d���Ш&_.`��K�)x̅21FºtE����O�W�F���ܻ$d�x���5SFI��t���s����u)�'c���jAꉠN��O��j!����ē-�J�8�Z�����R���܅�v$ԉBa�V�~�lpa)�<��m�O��Gz�O��'���Q5Y�,�����U*^�hA�Mϕ$!��9AM�O���O��$������O���6B={������ԏA���p !�@ВH��y݂0�rI�[�'�܅�.#i����򥖤	�L�06�A�#��}K���&3����c��V��9V�yK�{�	q��H
�B��/�Nyۣ�[������8G{����_E��"!]�0��ܡaW�yE!���?�� �t��2u���#�Nߌ:�qOln�̟��'�X�@`�~J�4(�pI��9�h�hև�Bq���'M���`l�'��	�"!2�� '@�a�,��.G;���
�U�j�2B��~X�@{�#!��qӢ�̪pDv�(��4B���a���xdI���g^ �p�X��Mc�Fޓ(>��=i�O����>�g�X5t j�U�$	=h�G!a���=9��
"�=`#���ޤ���a(<q4bň86�����v��0�FN)������C$*�4�D���|1!���MK���M!�X�c�_�<,a�T)ڔ�'FZ�jP'�]�n�y�G�](��`�~���r���_�@��)I�-8�x��Ֆf��l#�ÿc����X����Z����c��O x%s�.;Z�V[�L��G��H<!��O>�D%ڧ�Ms�H�9pp��de�?���{.@k�<!Pf��Tb�@:�l�?�>�5��R8�tj��䝹/9�	����+5:��ҒD��eֽ����,����<��㝖2G�M�I�����NG�f�SA�<YƬk��^�	RT�@ש^!#}t�zrC��WE ���CQŖ��&g���H�	�0���9��˟,��
UO\^��h�-��cJ`,� #G:]�`��p6�̐�yG�Sh*�Хl�!�Ɛ�0�ǍD��d0?q�O�I"���p�#�)PѴ��(�	`�m�ȓQ@~`k�K�:�̴h�MZ	��a�O�dFz�O��Y��R��[�g���!���r�l=Y�� *Ab!�3jά�?i��?�������?a�O2��QAz�lt�ce�D�0�A��,zhp�T��:�!�����G�b� ʼ(A�Fo�L8�a߬H{L�٠a��@Y���5{*I���ii�,x�DV���'n�T�y�Ej��ʯ*�6 ��m��h�	G�'�O��z�%�x��8�Ã55��Ң"O��[E�H.H����Vc޺�1+������5�Iyy� <z��'�M[��Q�
n����Y�D�:��rn����'��= ��'�"7�`Li��SR��y� 蒨?�}��)��,���a!���s� ��]�f�?	�+j���ɞ�6A��OK�):ء(G%��n)r��n�+>�vd�4-����k�RܓHW�d�Op�?��Uړ���c*D���U42~v0�=I�R��|H���,s��
T&B3�����:�>\i3H��n�A#�_�s�1A����?a)O��;"�O�I�O@�'J� i��4P1��L��c����$D�#�F��'�RHŦJ �;c��%sT� ��n&S����ɚ:r���&&GbP�x�0*�|�'�~d�קY�]O�@����]�`�c��؅���c/����V2th؄$����%g���Oj�}"ݴ/��e�JD�S��@�0�F7s����qnt	p��*Bx�p��۴�Ʉ�	.�(Oj����ϸ?d0 �Q�FrP��퟈�	���I 95jHE&����IğD�����2,�rD�R�M�&2@%G�
��N�@�B
���i22�G����|�I�|���)�<4xp��+�� ���	(p 8qHN!Vd9#���S��H�BMO��{�ڀОw�@Yh�kҏn�j1�C�I��Չ6��O
�q��4�(#=�U��0%3 �f�`9r�`�s�<������H�,]���ve�l�ďJ�����'I��$	|#�蝆['����КfL*��"]8���?����?i�'�?I�����+��e�Z?�څ���G�0,��S�l��Xp(P�~��p��I�{e!i�O.*�tŋ@i=f3��q<��2��Y�>��ā�e��;1�Ʌot�㞀 �/ÇH�~��+�.<��	è�~��' ў�>���]H��	�gC�%P `�aJ�<6��./��kʊl��4�#n�$����'�?�x1��\6-��:T�@y��
_�t��&O6���	ПP"ß����|�vdB�&O��� ���:7����*�Rb�'E	YѢ���DȰR�����B�e���W���A�2�C��.wi:���P*x��Dgnm�>��թ�/�qOt���?�OT����K!2H�PI�e ���W��0lO� �$�E
J?}
�4�'Α0np~쳳
O�!%�٠r���%�]+q��H��kM(D�����<��$�,�?ͧ�?)-��m���{�(M�EX1y5��B�R �&������I�3G�|���:[R�٩��Il�u+���'A��FL�f0��p�'�`��L%�2�i��fm�C�N*��r�
�C G�,TB��y\d��d�w_~��6ɩl��O�����?Q��ic��d+�#H>W;N�Z£�Y;���"Oj�r��\�0��g;m2@�ä�'���<)&��	���r#�* �b���J��r���'"�'.l�+��B����'�����
[�CM�q��M��#�n�&P�?�|E
�C�]�&Q3Ѯ
V	�����,}ҬY�}�@ѩ�mD)T9�� ��DM�ƭ�<�� �aF�V�:P�+�D��'�M{s&h���D��R������M�YY>��c�
��?��O�p��|�����hxA�D��C� �:��:f�!��|Ѐ�"��q8����&ׇ.��2���Sȟ�'��T:c׺a1��*�I�>v�B�u�R,#D���O��$�O�D����$�O��S� r`Q�A\�Q�AcI��`�d`�9�T�/v�5�,�Z�'g�(׋E�'��BbW=VF�i����}����2�[�NM�U�s�����H�� ı��{R-H�s:A�� It8�0���7�>��ПD{B�D�.�Y���P|�LS!�$\)q{�����8H���+�1qO�n���'H����!tӚ��s�J}��D��T���d�Ϸ�"����Пx�I(Y�P��ʟ��'w�j��b�B,�b���	�;,f��C��<^Tpy����*��{��ˇC���c�8��I�
ւV:>��Ȝ�Ħ�ɦbҋ&)2�s2���J���B̖�XOfqɁd�`�I�ZOj�d\d�D��pR�P�D�b�R6����!�
<H�������.y[�b� �Q�|D{�O�(���O�;�B���
0d��j�	[	�'?"��N��d�O�ʧ.2���4EF��S�J'P��eAIovdP��'�b�:nr�L�Kl),���?j�Ь�%f�X��Zc���5���g�E7A�hO�|hT�ʐ~�FQ2��L)j|��G��p�~�-���Pq�G��H�#�Y�t�@	�f�xB�F��?Q&�|����+.%�6f��
R� ��%��y2�J�6(����� ���P��p<!W�ɰB2����M������nI��[6�i>��'A򈖽ay��@��'	��'��;N����`�C0�����X�N]��Q�Ij���G�'[����ə%y��S�|�U���S�8�DM"�!�0���;�E� s��m�bX$�tpp�B�Z�Lz�4�nΙ��w����L`�mr�����.C�jA�I��"���xB� 2�<����he#q�S�y�mтa�|5�"�]6v�����I�HO��/�$�,RqX�9!�PW��U��/ݚpR� M˛z2��Iȟ���ϟ�3Ywt��'G�)J�v� �$��/1P�$[�f��.��U���9]�y���ĩU8�qK!�5�#���اl��-�L��n;p����.��K�V����S���z�,Ն��O �2��(j+�<I�C�d�4��6�:S�2�'���D>��J�QP� 	��"�P�5��C��8^�ܫ��גLQ��e�ޕ>���I�4�?9-OTd��nJ�D�i�f�w��,,&�����&����O���Ѯh����O>��%^�]�e���������5C�|]zU�ЋCK�y`v"�6�ޑ�3��~�'|��%�s� 4�üG�������G|�ن�$���x�ʍ_�џ ��G�O���>���yVd��1�M�g7h-��}��?�˓L�0a����4�������	d�l��?g���Pᐭo��x�a���P�W��?!.O&��0 Y���T�'�哵y�FDlZ�l��G�&�RY�b.��q'0����?�BO�z�jW�+�!bt�����x�T��lF�Z�n��>S@P&�,�ēB<QcJj�!abkǼhY2I��FQ�3NF�j�!Y$"��P;Q,W)>�FOe�f�'�B�S�y�w-��
�B�iH�Y�`�EO�'��x��!�&@�'�cbj	 ��ֿ�p<a��	�p���&��7���QN I��hG�i	��'��*�,z̳��'~��'���3�P��D�ѕ@�vuc0��&	~&�8��	�kQ��@ǌ[�<��h��F��1�6��a�?�3$�<Dg�,Lt�����, ������4`�$�ĮR��j`k�C�\&>���F���y�0x��Ae�A�0�� @�+K�$,�E'�<`���Oq��'�F�Q��J=e�1r�F�<��'ㄘ�� H�\�L��s�]x�ͦO�dEz�O6�'�T�Y%�KP�鰐O8 ���2^��"@�O��$�O
�dJ��K��?��O�����+�>~w��	�g��W�h��wiUb�(њ0$x��/J����k�v�'�(	`�E�P�*���i�&���)F+�~4�tx��;��&�h�a��D]`�Ey����ݖ�R!$�k��UIc��j6���QQ�~���J��Q`���4���@5�y
� �ta�ߖ %��%
�+)�Q��ꦩ$�xv�D��M��M�3cK�<`��d/,��b�9B�'�t	q�'�7��I��MW� ILX��թj ��	Prk�$� a�|	9�!ωD!`(���(O.{�"Yq�����g��D��x&���v�rb��%D[�|����]�@�1�L�1F|�GC'���0@�+%}�̚$"^<�B�ļh��+��#�y��4v8:`X�FU�d�fIS�� �(O�=�'}-�������U�W�Vu���
��� ��m��j��ib�'��S=/N
HlZ.|��Yj�=KV=�BJ�B���?9�DY�!efPQRh��4��a�tR?%*�	� �T�?�t�8�2�1L�!��䄭|*�A�� '��O���T�U���t�V.c*�L<�!��4k�4?��&�'Ǳ���Q��0�mZ�?����v��O(㟬%����
��\�@�'�)�NA�g�&O�n��MsI<��Й=����b-�j^�)��g�7��O��D�O�Y���GL~L�$�O��$�O��؄P(Ƶs��:B,�9G/�����x�dX�UVb�;�B̂s�p�@�IИO�����ğ �c
Z6DZvXfʓ�D����
��uj'�ə\��� 1�a℘�}�%���E-�N��7�י*w�b� ���M:�!p�"�䙝M<��L<�@&�\�T���kԅ}x^X ��W�<��
?u�N�"I�uBh`IuE�R��Mu���4�xB��1Ekh��ǉ�Dl�S[h�A�B=V;�=8���O�$�O�D��#���?ɜO���Y�բ|�ZM���� ű�O��x��&~���Sǚ�T��Ǝ9s�H�@	�'y�m���5����F/Ȥ{>��㵍҆�?��'�n�#���yN��hq��`)ά��'��t�L
,�TL��//Ij�э{��q�h�OVH��Ϗ����%�FL���=�L�rb�L���?�-O�"�DA�?��tZ�A�!|-t�
C@�d��`8�$��Ř5����u�,A�R	�f�+D�pгn.[�2\�C��8-�L	1f*D���1F�& 4� '�$S?��Y��;D�(��冗��yi�m�&B���@7D��x�J�0N̄@��� @Q�`'�8D�p��K��ϒi�쑢Rn��ra�7D���"��g`�u�n�
yi�<[�,"D����I��9���Nǒp���A�B!D��Zf�?M��H��dĉd�p����2D�����/�Ȋ��ݛ[3�ᤦ1D�\ a$�,1%"|�t!�9e�,Ru�+D��sS�Đ+M�pEg�1�����	<D�$�"J��*�Lyф�|�D�7%%D�(����X��`�j��6=�<q��&D�4�&�R�&t"�.x8�`˳�$D�0�.D�G��8�ӂ͡d�X�8� D����� e��hr�	�q���wO;D�\�fC,�ᴥ�v�!��H9D�$zC��N!X��&F
�2Ҏ9D�0�v�&�&t1�*�-aK�`V�2D�H�0��c��Ds���$����4D� �E��''��hE�D�r%|����-D��" ��L�Ab� PL 9%-D�����u&��;���'0R�7�-D�0H𧏞er���s \�D�ܻ�0D��t�JH7�$c���;Ɣ� ��-D��bv�Qo\��
�.�F�"i*�-8D�@h��X++��m ���K7:Tp��(D��A�`Ҁ*�V�����
)8(�	%D��Bt��I��C@Ev��b�!D���&޷�>ɡ1Z
����ԯ$D���F��v[D��AK�t7,$���(D���t�YHY@\Ѳ�� CK����(D�@���L��L�qJ!*`��2�/"D�8"�
6m�6�K��F�i��%9D�,D�4��� V���#?:2��),D�8�&"�"bU#R�V%]�ѯ+D����`S�<��a�+�C�� ȁ�'D�� R�qb�π`��2!�}ĕ��"ON�J���*�>�"�o�x�x��"OjtB�l�/A��en:���@"O�x�T��P� K���$���4"OLHJ�#�C?��3C-��S�Z��P"O�"����9��F�+�h�0�"O洸ŁW>���ؒsVW"O�D1aK�aOh���(u0�9�"O.��'�Z.+����J?hB$�!"OƜ(�LI� U=���:\��C#"O,Xk1�O?)Xx��`���!N!#g"O�X2�醬t6hLA��TR*�#"O����T ��4ʞ�Vy�"O�����(@]�8��'DV��%aT"O"z4��"O������&D��*�"O<�rKP:&%8dh��M�n��d"O2T:`�_�@�Q冿#K���&D�H�Eɜ7+���rg+Ĳ4ĢD�!D�@dAG3h�t�"�gV �L�0DG?D���1�$ ׂ0ɗ`�C@��2�'D��b�ߢY��T*��i(��&�'D���'O�?,Bq�O�a�807,0D��17�ךD$)ɕ��m���`U-D� ۰�OD�\y)����e@؉��,D��A��U��h �W�pˤ���*D��; Ė�dx�9��V)�4d�3D�8�.��B���+����A#.D�Ȼ'�N.��9Ս���*Ԋ�L*D���U��9׶�AKЛ R�{1�*D�0*Tɓ�9K0@�D��,�z�8d�-D�4K�b> �&��F5��{@�,D�,#�Ξ	���"�T�DQ���+D����O�2���qL�.7�܉P*D�����@��5D���C�(D���S��bV�c�nX�l8��+D��K�  ��5(�ԲF�,�5�,D�<�SK�
���0�i�!-�:@@�/D�$	�cR�HnAʵL͐e��5 �'-D�X9qh¿"݈I��
�#	�� �C*D�h��چ*P�ხH�v�P�*D�d(ׅB
Zdȉ�ʘ9&E �g*D�`[�$��|���u�6O*�y%�(D���A煫)�r��-T"�����1D���f��C �1V	R9U�`�Rf�1D����H��b򭲔��C߄P��-D����؁~�b�u�L6HZ��9@�%D���fnD�=(�(�L�qvoC�y����;��pi儂� � kD��y"l�
q��E��1K6�<��MӃ�y��J�	A�L2@�n��)�yrӶj��LٱN�G���$N�y^�w��XЫY�O�ʑ��ȕ�y2d� / t��j�@�#'j��y�/Ă���7iB <�j ��E��yI�\��@p	�e�ZD �͂��yb�(���� �*l�>�C�d�1�yb�B�\U�U� 2j+&|3#��(�yB0�~Dr��'xF�Djs(O��yB�ݵ"�j|RPm޵]Ɇ=Ӓ섂�yퟓ9�[(���F?��A�
�y�H �v�RÄ�[�Oϼ�2�֜�y��9-��8�iH�5wv����M��yBi��`���K�0d��h�^��y +�Ͳ M�*g�D�g��2�y
� ̈ �N�a4͠EF��'}�a�%"O8La��A�jyv���>��ͨ'"O`�A �@1��Ƞ�^P9�"OF����ń`�;JF�A��yq#"O�P��T��b}!����8�2"O`x�Fg�n&��p�Lkt��Q""O����6@�(ɨRC�	J]�4�"O��!/��W�\�i�@��aB��I�"O޵�*-Q&��,3:�"O~P�� (�ĕ:5�H�m$�I2�"OP[bNC�{t�Sa'��@D���d"O"���)�n�����F�B&�h*�"O�2�ə��:@��$��PYh�"O�h��ŝ��*Y����E��JW"OPq#�&b�`�	�);5*�%*OĚ`'�'&Q��A���P;�'�*]��o�Aތ��&���'�`�su���#�౲a�>th
�'ͼ�S���1Mƞ���@�&� 
�'�`Y�*��P�2V��1}^��'S�`���J�&��#V#Z" ���'�JGO1K�98g�V&�5��'��(��G>+RD�����"���*�'���z�FܤF9�P��L�Q��i��'ST 1o�%gm�q�GiR�y���q�'%�	VRŐ5iG$H,a�vի�'�P�an��}"�AҜYȘ��'dȰAl�*=v�b���)Q�V�s�'�2�a���/t�&	��g��PՈ2�'���+��\�w�й�S�C�F\ƍ��'��J%Kͳs7n�X��F�?ܸ��
�'����⇳G{��鳭 �`��ɳ�'��X���?4ߪ�1t��-�*��	�'^�
aL�?p�޸��$+�J�P	�'{��SɆ�[.@�Su@��%O���'�d=��/7y��Ie׉��	��'#�8�@f
F��� M̀�n�*�'�X9��-0]��0�Ά�@��0	�'Cx@dj��%ӠHq��	)���	�'~�̟Mb��괭�)�A�	�'���Y�^1�t$ʰ ����	�'+����,Xđa�
R�`
�'$v�hvdG�o�b�� K	{t`��	�'L9BF+�B���1��Ӄ}iT�	�'�9���?Uu4�ڷ�Y�h)0�c
�'�B��7��Q��| E:A�	�'eb�˱�nc4ӡD�\��S	�'��� ��)^��`�G�~~�\b�',��.E":���c�FR�g�0C�'I`U���x���Y�#M\����'�>��lT��X�y6�Gf%P	��'P8����>/h�0�b&�X�tE��'�i �B�5V(�b(AÖ81�'J��F
�SF܁�� �3A�����'��Z�ȎQ�0	r ԙ4/�p�	�'��Y���X�`�!A��,���'{2�u��W��@��I��0��@q	�'�v�sG`ЋN�X\��΄�[�>��'i��$�_��t<���O� Ʈ�9�'�0�2R��Z��| �&�m� �H�'��(@WK�r��Yf$O�b5�y�	�'��U�A-��A�<��e�Z�(�T���'.(���X4���$̟76�lI�'�B4�%Eޜzsh����3"�r���� 
`���:QX`q�&���I>D`��"O��"�^�e-��@sƟ
}Qf�*"Oflb ږvB�U%fC�X�dQP&"O���SUbz�QĦ]�	�@"O����R�1��g�x�{7"O5c��֣g�\�U	�q7��i&"OAǮٗm?���ʓ_Ef�""Otpbq�^�	���� �4:.0Ɂ�"O �Ӱ+!�2Ap�)�_ \���"O,�aU�
4/�!�eV-1��x�"O�H�t��^�6�g��#T��xЂ"O��J�K  �f�r ��	�̉�"OzD��J�"\I�+�G��=s�"O~�h�l��a�4̰C�`!ԆL��!�d��L��l�Ц��|��t�4EH{�!�7S�<�c��`��bA��(sf!�DߊnpЁ�e(�XXbA�!��K�!�$N�D|�*��G\i���e+���!�đ
\X���FpA���6(.!�$�pт%�E�p=�H!�ղB�!��.T48�"��}��)t��+}!�Č�I(��HQ���a�¡�e��8
�!򤜁E��j��k�ތ;ҩ[�f�!�dڏU:��Q� lR�,�C#	�!��'��
�C1G#���#� !�dZ�n�"�z��6gw�| �`�(�!�Dׅ����F�0D�"E:�!�@62|�xkI3+�|y�@�Č�!���R�,��@��6��{��U��!�:D�<���D��Y�
���
E �z�n��"���Fj�����j�w�h|p�<V��a��h�<3@�l��8hd�7jg���~�<�' ��JT	��92a���Vw�<��90q���*�p�}��-Rs�<��G���P022q�t9G��q�<�f�G|@�[�L�nB�8!�O	O�<��Q6+#�D��aM�u����FM�<q�n[�Z���`�٠�Z�&�K�<�񍇫F��P�­�T��`��^�<A%����a�"k��?�RIr��[�<�S�x���(��}Z\��t�T�<A�k�6zD��9TDӤ%و���o�<�PA5��y�7���B�ǒ^B ���?����P��?Y�3�'x�<��>p�0��\ en4"�;]-�X��y�FI /L!��p���I@����<�X��e!ˉyFaPUMX)��u�<���22a�A��d̃r�J��T$j�<!�(��NF"LhW��'	� �a�h�<���7�(��@J�9aNqh��Of�<�t`ǡ2���dJ��R0�1�%`�Y�<��Q.`H���G�yF�D�.�R�<a�N3z���A ��j

 +EQ�<q����>VV0P�+��`�M�7Àf�<ɠ,�9-��Ո0茠:�FR���e�<�%͊8�-��,�}�$D�(Db�<�E	���-���^W ��h�G�<AG�ȢE㸴0��IQ�]zC�h�<�V�B:e4�,ZQeb$��b/\h�<�R���S�����6���r" d�<�e�ԇ7T���?3<l#�Nu�<�B�,M.1���M>�Yc@�q�<A�fג@��w�E�m�.�Y��Fs�<���ҳO̺��l�9�H��� M�<� �x�����T5�S3��	A"O�DN��*�IԀ�us��6"O*L15i�6Rʚ�[�Ĕ uI��r�"O�����	o�N�r��#��M6"O��"UgW�1�4���#;���"O�\2�ހ��E�& ��B�� �"O"�Ap��1%r���G��b�Z��b"O��3�B [TJ��G�%f���3�"O�"A��Zl��I�F�6Akp"O�1���0b�
��ʟ_��9Z�"O
8���ta�9�cnG0X�`�s"O�͹�[�n�L��׆ܖA�8�8"O��+�+
�>��Y��M�:�65�G"O�kv��#~!�Ɇ&%5׌�I"Op1ۖM�8l���#V+(�pG"Olq(�M]��4İ�
�v"hHx�"O�U� DC>-� 
 �^�8:�`@"O��jǎ>4��!�mE({�6"O �����o��i�	L�b��(�%"O	�2A=E�\Ö���.���"Oู���XuP8�'I�C|�	��"O�Xn�'g�ԀR�NZ%?���L'D�pz��>lk�աEe;JԘX��$D�����d�N���G��! �@#D��y5���o����d��!�c$D��ف�OQ�5B��ּ(&F���'D���p�Ix}&�SGY8(扨Ӏ$D��2@�6�2X�H�j�"�-%D��!��V&	b�HH5�E�Usȡ�0D��H��'a��P�q�5m�}ᶍ?D��Dj�r���PI�0������'D�dR���z��գP:b+P��$�$D�`Ǯ���)srr���"D�@`��P�)o�Q4�ɍaئDk��$D��2�F�C!Awǃ��~�(%�.D�,K6����@vfB.x���Ae7D��R ,��9�hE+h�d�9P6D��bJ$b�=H$�.F%´"6D��h��V�yF*Q�Ч���M���.D��y�,�i@�;�D����+D�H�ę4Tt	b�Y�c�=(��(D�@H��?��ԥ��NHu	�5D�8)��D7�Jԁ��C�J �B��y�$�<��e��Ǩ	"\H7k��y�'�~�BU������������yB�ɒt�2G�5���ȶ ��y�mђlq���y����X�}��-�ȓ%�a�LP1rl���Rh�&��ȓ3��#�L����)�W�Y�Ň�%J@�+��WCz1��I�\�����&&�4�C" N��a��3sj���6=�8���7n+��e��U��̅��$a���>3؄�V�Q(?ڂ݇�-ˎ�����~���0�#�E�ȓJ���0��g�d x�&P��r��B�zDp�ӓ	���	�@�a����O/B����E�zd��+28�ȓv_
�a���7�R�gE�_��q��Pl$d1���T����3π����6Q8B,Tt�(�*ÈsVt��ȓmQ�K#8;���@�u�}�ȓ(rl��E��(��ۗ"l��W�0���+1�p��L�y�LY��+��@�jP�x���"f@\h��S�? ��qu��T*lHe���Fp���"O.��D�PZ,~-�c�]
���"OM�2�ý4�9{��O>[�@��"OF��MF����qPO���+`"OlHq���?�������*�eٵ"O�D� �5EFج���Y:ij�q��"O����_�l��h���R�fj��
�"O�As5�(^� il��<���P"O|���[v*谫!��Y�R�yR"OTU��E�cT,Y�¨�oP���U"Or��-�4�|��o��+*T E"O���K� M��sD�-E4�	�"O6 �-��Y����#Ń.H�p�"O:H��%6M�O�U.E�"O*TI�E"�3�m˞y��)"O6�xqh�; �vi*�C���ɤ"O��r(Gq�R, qe�60 j�8�"Oj�sA��-N�̳�K��IN��"OL� ��FT�ht@��=bX��"O���������Ȣ ���H�"O�8z���� 
2��咛u�:�"O(ժ�Afp`���?o.��`d"O�hj�/;�{���98����"O���)
�!�� ˃~�Ոs"O:�s��(n��I2�ʞXzi C"O��y���>/��@���>o.�a"O,� ӄ�9XZ����剟Ŧ$B�"O��pA��P�@����/$�i�"O��Ђ˒(6L�+@Bx}�0��"O�x��L�q�@��$7aP��"O�3$�*p<�9��`�{ �tBe"O��p�c� �,1��j�(Ic"O6�(`K\3:Uv]�%@F�g\؀�"OR�¤��2�E`AF�HJ����"OЕ#�38'�EҝwG`��$"OLPfܾu��!�f�f���A�"O� �#J u�����rB�5��"O�P��"�9����	�!�d@"O^ �&��v"wA�<�:E�"O�9	j��<T�d�S�B*-��lRA"OpYW�����q���<���c�"O�����BqXe�Ղ�@q��"Oά0���mT���sM 7:*�g"O
<:3@ݰt��|9"O�(��@E"O���ہ2>B|A��]�4$��g"O8�d�?vxȡ!�I�|ܙx""O�hyB��*w }�wǐ�%�5x"O�h0&�߁It�i�hH>F
���"Oν�'��s�։s�/�;���pG"O�Ah�fQ�"}��hC������S$"O��rq&Ĝnp��j�,Q�5�0)Q�"O��E!�]��ꊝh�bٳT"O�A��	fQr�s�8=/�F"O��$H^����hޡ�����"O0x*ī_"Ц��3�I\��@"O�9ZG�̒3�^=0(���䵑�"O }(�%W%ļ�`B��2D��(�"O�=0��z���U%Z�C: �{B"O�<SĈ��_��)�Q���mFR��"O�B�ׂKZi����<��e"O�P9� Ğ�@�bԏ$���"OH%�#��8n�`PAA&v����"O���qaB!�v��}�>h�a"OҕJ�k_�-e��f Y���a�"O� �ܙu��![d԰`��.4��\1d"O�r�&�}7�Y�5�\�]Š|Q�"O6�A�OS5]
�|����6[�x3"O~!�6nE��@@���U�

"O��S�=�m*$��)i��` �"O4LC���k�@Ґ��;KL��"O8t�G�k��4�5	��Z2"Obd
���$K�����׵@��݉�"O�]#uK�5�� �&@7+��Uh2"Oh@+���%/Q;�-���p"Oj��$������m#5s�I�Q"O������$��D�X)\�!Yu"O�)t��\
�S�:�u�G"O pA����xjq�XGV�
1"O��z! �)������)\RA"�"Ob�˶F͘,3�e�)ʍpf̴��"Oδ��[�n���nY�2�J�"O���d�.2�2yY-֖VI�ȡ�"O:�*�	؋{9�ѐ��
O�@c�"O��Rd$� eܦ�J�����Y�"O��H&���*��0�E��.�8B"Ot��$mB q��9t�LB��8jC"O|�s5͜��z�
t�%� B�<�s@>X��A �(ŚQ��l��JD�<Q M�?s۶�)楐.r�<��ӥO]�<�U��V�&��ؒ%��A�C(�b�<1��F?APU�VJ�-A�)��g�~�<�b�̈u�N�u�U�>��q�נJC�<A-��A�\���Y�]���H�<)!��/W�R@w���f������B�<t@زW܄@�t�Ap�d�d\�<1��2B� j���='(HR��Q�<х��?+l�Ũ���@�uŝs�<Q!�R54�2%�\��B��p��LH���M��6HQ�O��0D�E9���h�照`��l�v"O�q��i��=���1��7�ܺ�"O
=J'��8�J4���4C�����"O.%�W��vLN!����W�ġ�W"OV�X@�(���s'�{��Y��"O
   JߙoZBH\�t�6�A3"O��X d�ꐉ\u<s"O"8SA�|gfy�h
�M(�"O���)�o�Ȥ��A���� "O�)Q�$��
�v|��j�Rix�"O�P@��ڣI6�\�G] �@� C"O%����'U�<i��$�*<(�(w"O�y�'B	m��u��#��]�&��E"O���v-B�r�ӀH�,��=��"O	���{�%�ʶ[B�!5"O��Aޒ �$XF��Q&&lC�"O�5�Ā�+��0�%.�jP"O4jD U}\�iFM>X�)�2"O^(:��������&=���ٶ"O"����@4(��4Y�V�(�~�"OT���h����qt�HW�Θb!"O���Ӏ��,�� ��9G��"OV1�c]$Sx��H�(C�mv��"O���#f�nuIcg�A� "O؁Q� ^�0�*�:�F�h>��;t"O@���U��0\��Rq��!�"O��"��D�<�w�ځ�
���"O�4҃��&"b]�U蒩#���"O�س`�"F�I��f-5|҈;�"O��y� .8�8XA#E72�433"O� ��1�1.��`0&h�Vh��z�"O���F� T��b���"
Y�U	G*O, ��N�iӕ˃�'�*L�	�'<�{qO�a�*H؞�3
�'r�H�ժ�2�j\	d+[�N� �k	�'=h}�bǔs�:0`&B���3
�'�V�b�ɀ
Qn�c2#��;@0<2�''<II�(U'zz\
b�*:�T��'e�-VFD%H
L���#�.E�'TXt�b#��,���pH�"F�d3�'��Dh����h�(Ur�M"Q"^��'��];�)Sg��u@��,F	�1C�'��a!KY5A�]�7��94�(u��'�@��Q L�h�(	ǂK�����'8��8��G,q�|��R$����
�'z�dq�M�f� �z������
�'tf����J ���f���0T�	�'��p˂&��r�\r傧a�%��'(�P���B��.zR��0��6�y��-��SG�R9s��@#�G�yb��m�^�PAE�fʚ��� H��Pyb/O<h�4h�-*� ���P�<��/�Ul��"dҬ5�L�p�PO�<�7�,�y�� ����4MO�<Y4��:	$da�쐍S�0�e(�u�<I��KJZTr��^+�`��v��|�<	m��@Ѳ��$�B��G��v�<	 �Iq��0���@<���)�A�z�<�NI�.gK�b��i`$�ǀ`��C�	'}�����%Abl��"%�E�]�C�IN�$��EIQi��
�V�^�C��Ct��J�i�*:v�3���x]C�
*D�"���l��bNO	P�$C�	�F�V=�S��LJ���<��C�3�P�H� ��DHrD!ї?�pC�Ia���b(�v��!xV��7�DC�3)��P���*fӢ��u�:HNxB��0_�Ar��`t(�J,x�2C�Ʉ?���ʇF4��ˇ��{�hC�ɺ�5���G��H%��:6�>C�	 x&iц�1[e��4�I.N:dC�ɝ?���aQ#0����
z��C�3"K��qti,��	������C�40x�􃊩c��9B�-� &��C�	5|���P�ٴe��� U���#3�C�I�G{�+a΃��u��D�4��C䉩l���r����x[PM�c�S�YvC��/MB�A�̂�-�|�tf�5FC䉌/�0�pE�d�J�1Ћ�/]�XC�I�~DB���^���S${T�B�	�l��x!�a�X�E�����DudB�ɂ!fR ��*V��%�D� $Y�^B䉩Q�x@��,Cy��;�`��K�z��d�<� ��xP4á�V�wՔ,���\M�<�`�	�F��SIC)i4R���J�<�Ӏ�Fl��+��R�C�(� D_G�<�(�/Yo�5z!�E7��7f[D�<�f
�@F�KPh�c&$�2�i_K�<)�B9X�r(��j�%+�|�BS�^G�<I�-')HbYᢣ�)D����KD}�<�pO�.9,�0s�.�=zR �I�y�<	�k�0OA��z�[���!�Eŗt�<�pY-���t�#S�,C�jn�<�NB=|��`�T�%63΀�$D�h�<� ��Z�(H:;�,��(ɹL�|!��"O*}��Q��l ��-�6Uq�"O�\+wB�I���CM�2H��"O���BA��
��M�bF�Q9"ON�@���$�d�ñ��|P��r"O6�)��]#6h���*{���"�"O쀂��(T���BJ=:��H!"O��:�+9�|��(ŝVo0l�C"Ox1�/_	y���v�Gb2!�c"O\i���;�� �H�
6%��P"O��/�f̱��17>R�J�"O�3-ج	�n�I'`��aP��zu"O��W-_�y3�ٔv5*0�"O"�ZŧX?����,%��:�"O��܂ zj�Lp�K�!u�@�C"O*M T*�*�`�D�/�h��"O�͋+�ń�J ��3}0�i�"O��0'�\���0 �5\�k�"O0��gh¦�X���3NX�ӄ"OlH���e�1F^�5$��"Odq�,�9/"ȃգ�5�Ҁ"O�18#W7IH��4��3����"O$���/6�䉐�����܀��"O�%���GEh��/�=I��<�"OV�1Ec.(�=;�n3nȒ�"O�(Ʌj@8w�@4�s퇐���"O�����`ب�X.���P�"On���Nֶ��uص]�5U&h`�"OV��b/�"����07���"O,)1�HR6H��K�i�.1��"O�����S�T�Ш�@��~�R���"O� sCM�6�1`�HS7b�*0"O&t��G��F�"G`�P�$"O&�h�@֍rfԸ���őC���2�"O�(����@�\!��ތ�a)�"O2��*Y(Q�钲Ǧ<��"O�u���O6%�&"�L�xTP�"O��c��x�N����%���Z3"O�q���Ś-�T���΁�a�<r�"OtɸF@*p�� ��B�fZ�"Ob,!F�8�ހ 1�B'bZ��*�"O\�Z �ZG̠���t_�Y�"OH|Ĥ�~��)�c�ID~��P"O�9���T�
W.\0&�Ek7����"OL�J�k�y7hUAՁK37p�e"OzԫR�K*7 <"��n�:qC"OD�Z��Ưd@����@ˇ �JH �"Ot0:����8V���2�ʼFx�C�"O�����6^xeHD�9}4���"O�P���O�	Jx�?_��00�"Ohp	� *�X�`5.[�I|:xٓ"O��A2CG�P]���D�_ն��"O�D�a!>����9��2�"OX�t�<�0���)\S�!��/K��ls��(%���HZ�X�!�$X�C��� �K�79 &���G��9�!��w] u
4Nt����%.!�D΅q�ʑʤ`�Y͸��A��!�ۛO�]�!��k)^H�#G�!��>�LL��C ��% c�P�P7!�CS0��X�K�� ��&ןh?!�d��[��%�ua�'_�H�'l�1S;!�d��	�%K�W��}��G�E�!��6 ���(�M@�^dIr7iQ�v�!�� *�1Q&�=6x0p�,����q"O�0�Z�"�g�%|�Z�"OIs �Sx���O_�D��P"O(hU%�/oϒ��(U�M���Pr"ON��G_�c�T�u���i���*"O��Ӏ/�=cڠ6�L��Eâ"OU��ldǸ����gkB���"O� ����6��aH`AޚkO��p�"O
�R�Q3*�"̘S��.%x��"Op-�&�'|1ѪVj��S��h��"O��S�ğ?���ң��P�1c�"O~�X��G�5 �"@M�����"O����b�=aTlT�&Mӆjy��S"Or��7$C��!z��3'D��`�"O���oцR�^����N&+��Y�"O�K�?�����#d�	"O�HSoҩuY��cU"Q7r�\YW"Of���"}N�zǠ�e��U�"O��@�f�ޕ��AƗ�@+�"O�I�˘ �ʤ��	�S��i�!"O�KcHC+�hs��B�3�t�`e"O�Af��O(̃4iK>EJT"O�ي�FC�~��2�Be�F��"O&���(؜ ���2Ђ8�
���"O$#pϜ�
�.X�"�M7 g���p"O�@9�O�F��P�$q�IS"O��aаo�^!!��-)9ri1"O"�!�,Ls�XՉ���8*�S�"O05˅k�>".z�b�����YK�"O>��U�D�&Ŕ`���Y����"O8 bV���Tn�`��! Y�|T�"OD��biĭ~�:�BFH�)t8b�"OH-�`��^0��c��(�^H�a"O�  J���eu���{F(��"O:�{BG+20E�4�I�z���"OQ0�f� 6
M�@�.L�L��"OB�B�ؕ��I��&,�$��"O8�!`�.QM�0Cf��Q�th�B"O H
�́�8yl�h��
^$�S"O��)*F�h��9B�˃`(��˵"OF0Iǌ�VS\q��<��"O�h��ԭJ�X��"��rU�"O4�H0/�vw�c�ۆB�H�"O��KO߃b`:)���1:��I�"O�+2�֬&�������G
4Qf"OȌ��NĎu�@�RvMX�T�^ջQ"O�EУU�V����²`r�"O
ݠ�3���Jaa� �j�"O���uȌ�wOfgeҁi�"O�XXb̓5�fIIٴ@���5;D���`#?A�2hBBg���Agc,D��BLw����Ɋ/:w��3`-D�౳LI�m8X@����?�u;b,&D�\��+.X�Z�$�3XvU��9D�k򀊐%F	GJ_�j�r%S�L8D�p�E�$�|�U��39�H)���7D�����,j� �@�Ki��i3"�7D�@��2,��p���gԥ�0b7D�[��6︹�Vc�v�A"��3D���G�'�(5��Ŗ�N�ԕ�P�/D��E��hLz03A��1b鬭��#D�d����:���2���/��O"D�hhd��� qb��,��b��!D�웖cP�\9@�Ч
��byX�!!D�� v�w �ۆ]�`lc�HP��"O���ţR��Z� p�_��R�"O���w���,�Yt+
�O.)I4"Ox���i���ص�3I
��@"O@\��.V�k��L;Q߀a��8Q"O�IA#!�~:�<i�M� ߂���"O|p`�C�Dy)�홍8�8�p�"Of0�%$�d�lSK�r�L�a"O Z&&�GC>@ZsKπv�ꁚ1"O(I�)A�7�����Y�@�T��"O��H��E}���8�X���3�"O��y$� ��mBpP�r�	�"O�-����|�җ��eν�"O�I�`�M�S3�@E*J��P "O�qP2(ە;�4��MMm͚��"OИʣ��&*`� ��7�(%�"Oڴ�t�Ԡl�ܱ��<P�@�ّ"O< �:1���r������"Or��%Eh�Z�!S�גx:���"O҅����[(<�0	,pxF%��"O�tq��p�P)��ι*xfU��"OZu���X�8{��8'K_l�0#"O�l�ӈ�n͢��Ѥ��>k�"O���H	]q�q:*�z[2P��"O�DH#	��P+��Z���xy�]h�"O}��)��m~,��Z�0\�""O �
&g_�%:PQ`G��+A�0 7"OZ�zW ˇP��xGҜ6��8I�"O��*6"��cQ6T��fI<N!��e"O���a��(c�|�i�o�!��=��"O�uh������C��U�|�q"O���d	ͺ9b:�k��H�L����G"O^A1���1�^I���ܽc
�mq�"O�ah���#�\�ɲ�Hf�L��w"Oh���K��\��U�H�dP�"OH���?\����.�p���8�"O
�s#j���+�O�$0*��W"O�=;r�B�eϨ�@��I$S�0��"Ot�8��'enA�e��Zc� 6"O��0��˗g}&�Q��o�!"O���1�"S�ԡ�D��6m�
$"O�p#�D�+87x!�[JZ��2�.�yR�M�ΰ��Mӭ��l�B���yRh?+-�013��
 2@i�Q-�yb�<Q|�<〦�z)��QɈ��y⢌d"���E�'$F]� �oɇȓY�U�C`K� ���bF���'�.t��E*YN���PkZ�)ݴm��'�P��"KJa�(ya �\�!$�aR�'J�#�/�#�2��Wl�7��Q�0��ɗ]eV�a�R���"%D�V<C��5nǮ h��D��=b6�Ԟ3 �>I$
%�'��8Xg���G
 �����0w%��@t&H��b�'?Z�`�Ʈ�-t:L�ȓL�T�`��
����%]-<cT9�ȓ0TQ�E�͔F��Kuf���*��ȓ��HpG��:\���5F.@؄����#r˚;��x�Ü�$kv]��~����Fo�?+���ZQǈ.rL0�ȓ_V�2!�&fB~����(L1�ȓt@�� ��s����#nY�%��t��yҁ	��D�x�i7ņ�L����ȓB�lm#S-�RB+-�:b��9�"O���cȤB�\� ����\�"�"O� *ћFk��Q�E@�
Ԩ�"O�,���I��ΰ�gE4���U"O�`Ң�C�"Tg9rT[6"OfxSc�#_<a@�A,h�b$�'"O�ȂC��f�Փ��\#����"O�pb�e�&vFd0uϧb�N�	�"OxXH�.͵E(�ā�.�ȴ@"O��R� A6&e���X:���`"O(��A�L�P�s&T@ b:!��=��#&�A�p]x�#_Y%!���&��
��D��04�c��Gq!�$�H�ݒ�hD� ��� ��[�s?!�d�y{*,!��J�{?D�1@gQ�o!�Ŭ�l�c�Զ!#�\��! �!�D��Y�1��ܗY������!�w����AF* )f��$�R�!�ě3BUT ��d�.E�S��_��!�i:px��ȋ}Y���2d�)�!�I"0��0 �4e!�wC��R�!�D^�	�9�kT�6Cp}
�特k��{?*Ї��8y��
ץ�5_ ��'�k�Z���<1�"႟T�l:.�*4w�!�'��yZ����S� K´J5	�Y џ�Rg�:�'͔}Ӥ!ݏN��Ւ�CxTv��ȓ[ޅ�S�ĭ+d>i�p��*��m�']����=�)�'.%�0䮉:p�,!J����5j�P��"欩�G�V9�"%@Sb�k˪M�O�����
8@��y���o�PI�0e��.�0�@ ��0?9�(zd}C�.֊�XkT�M�4�Q"�t�<y�(6%kDmY�D�`2��
�ˀp8��8���/Z����"�TF3Ƈ��k�!�$��\T�
g�gb�A1�L�P�!�I�H��HWAR>7V(y10�_��!��X�(Ln�CcfM�=>�ف��8/�!�dи[�($A�I/>�t�ȗn��~ң��<A�m2l.n��MD05 ��z�GA_�<��#'����)X#8����,�c�'�ޜ� �4ʧ�t�#��ռzt��4u�lŅ�|�z��g���|��נ�l4tl��Bu�6-*�)ڧy� ��խP� ����W͐��]�� i��{�Ε*	C(#�J�i���=I��'G�4VLB�~I�����7Q�Q��'�PͨF��7\�!�GɃ�Oͬ8�
�'�Z�r�C�y�%R��ɠL�$�+	�'���#�#Ř<��DcՆ׋I���1�'�n��a�i�*d·F 9�'���'`\u]����8���Q�'9&� 2 �.C���g�E�΁;�'<� /ߕ2��`ץ��d�A��'��M�V�4``6Ɖ@([��+�'�����%�2���pU�(\S ��'w��ق,�8�t�%�*C���+�'��TZ�M� `����>|μ@�' U�$�&j�(�
u����=��'�MX&���22��qG�3I�P)�'�d��,�7Ud�vM��[c*5@�'k��U`�0~Z�]J�I/k��ii�'��P�
S�ef���@�h7n���'#�I�e�V�l��,���!\cRū�'@���F�}�F�5g��Py$���'�>�[P�����1H䯔��pa��'5���!.R!2<x;�GL`���'��=����M�b8�@$����2"O�x0!�0	���P��4bڅ�D"O� T0Z��ث}�"���%=p�(s"Ob�Y�-K"�4�b�9��"O6yC���"uA�P�T��}�b�)�"O�D���H((�iSSb΁/���`�"O:`4c�&3Ꙣ�Ɔ4(�Nܡu"O,ʖ�;�^y��.z�l�Q�"O!��؜l�������Q�"O�M*p���J�VX06��&�� �"OD8��s!rX�CU=%�]`�"O�U����+�L����]%f�j�zT"OL9�B�!"�r��P�K�RȐV"O�E��'4,DJ���<#�Q�2"O(<��i�� �Xw$W/��u'"Oʸ#3`��{�&�� cO�H�� �g"Ox�#�j���dvd0�Br"O���%!Z�uJ��#wJ�[V"O�@'�=)Xh9[ �������"O@�c���0Y}Di���֯e��qJ"O,X��'ʑ_ꔘx�Ҩ,�Z<�"OT1���A])��B���U���"O"�ɱ���:D R���$�ի`"O��Jb�-�24`A�.à�j�"O�	3ň��U24��/�i��"Ox� 1*�|�6\�`�P,v�)��"O| �ӽ6ZHTYva]5a�ę�"O1ۦ#]�+&PIAG�,L���`5"O|�p�#�f��RfdА�>�C�"OMH�EД0���(WD§={Đ�"O(P�- zD*��E�*��"O�����Q�A��D�llX7"O�	MH�,$|��1bH)f�0%�7"O���	SL�ة�!ρm7�8��"O���ҏ�>8�	W�[./+i��"Od���7*_�dC�.־q��uȳ"O�򥉉Qt�8t��?.�P�"O���AG4!6d
6'!97^�`�"O �#��Μ-�T����*5�+�"O�\�t�-V� ���_FP���"O�R҉S�~[��2���1q�(�"O, �r
�lE:��q��5E�����"O2T��N f���E��^A�H�"O��*F�F��$0�)^3<(�ș��'�¥�}V5#f���y�Q�6`Yjx���4��D�Oh4{C* bt���,Lj���[����&X��ْ~�*ĈՌO�\D�oھ7�N�<qaM٨݌͉`m��� �(�!�j@�󏅡T��m[�o�
]*�qO�-.���;�M5��ME��L��u�Ԟ�ҭi�E&T7fH.GN�Iɟx�	E����C�J
��qV�-���+��M>!�$�V�2�ʛ5L�m1qk���$JŦEHܴ���s;�tlǟ��I`�tM�;6��ȸwfɩI�2ݣe��Z�����(�O���O�!�+()���)��F�I�.A�5�՟m�%���j�����,A�pL��K�k	�N>Q����/]�����A8zi:�kD�^S����BN*t�d�����P����T�ШBT���e� ���<1�C��ٴl�q���Z�OP
<v��� W�rubC�O`�?ً}bJ�P����c^���L�PK��p>�E�i�6Mk���!ݚ	on�3tɋ�/�p��O�����9�	Ayʟ�O�MAČ���8i�)V$�B��T�g�2h���E���Jy4�8'��7v\�'���~�ڵȎ�Y��lp�n_�d|6��k��Y�T�9�]bCD��`.��^w�>ט%+f<,B��De
��1��:G�b6��E�bn��ţ�O�$�s�|�ô�U��f�BGH��J���P�O���?LO �	7dO��:&�!{R �SL�UΤ�<��iG�6�9�d���ם�;�z%!���*�cU�@ʙ8��?9��sV�Z��?y���?�G���dfӚ����\�RmɳG'�z�)U�E*khN��Ԍ�24��¨�al���S����h�E4�D�CJ���O��c �4�7� ;F�$e�⢔���T�"M�_���X?�mZ(ZE6͚�@���|FT*A�J���W�L	y�It��$���1O<����?I�OZD�2�R�3�=�'�\Vq�\	��ON��$s�� � �d��}�H8��Ѓ']��A�a���M�F�i�'z�4�O'�I/��XQ���	�`Rf�@�b������B���	˟L��쟨����ȟ���̟���3(JN-��kK!-�n�@�(�O�� ����G~BQ�ېg�8(���-�L�<)��ٟq`>�sR�Q[LP�a�=�f�ɷ*M�Q�.!�5��zB!���ڃ|�[�O_�i.��i*O�3@�'���xb@<}��-:ע�=,H�E�ļ'�O:���O���'8�>l��"&��ّW�ր�'Tў"}J��� Zcj�2�L0!p�@��r?q��i�6M�<Y��p$R�D�	T��j�M��M���99�0j�����!W*�O����OnYR�m�	K��wL9Τc'�.��4�TM�"�f��
f�%;���HOF��T��._�F�:rJH�2�����N�r�c�?Z��y'�L�I_�As��4!� ��'&��؜4bIfӤ`mZ֟��O�0��1�͆YyF&Ei1r����O��"~�I%PW����T�\y�!X� Ȩ��d�O8�lZ��Mc�4`pFp t�I��*��P,t8!�=q�����'3��q� ��  �p=q�=��F,e��6�o�Z9۱W���y�(�_AqO���'�d/��'w$� �   ��?  �0g���&� �;uhQ&�&��%"O���`	ôR��8��f����dc�"Obm	�O�0�J���D@q����"OLx5oճ8����|�̼��"Ot��U&�>5w`���ZDo�="O�؂��',�JI���:Z�rCO2���6�u��O�)���DD�(b)!�dM
�\0��nR�G���c\Jl!�$R�_kй�co�LoƱ�u��)i!�DǾfe[9�V�Yh֐3$رJ2!��L��6�!�&��{���Q��IR%!���O���Ԏ��v��0��N�dA"O�憌(��H�Rfޗ}��QC�"O.� ���5p4h�A�X�:�v��D"O6\�b�}#��I`��4���<�y�Bϳ,�$ $�(j~�(�ˬ�y"&ɢ7<�E����T�H�*S&�+�y�
Ǡ)]��VB�]}N��%E��y2��&����X_2ɺr��yb�P�ya� �# J�Wi"��E�a����K!
�ɦ��i�\thRB�"A1Oܢ=�|��l�%Ln�v���R���p��@�<�wG	�g6�Uq���%P�i ��~�<�qҙY9jX����J�W��~�<�E���~$YBS���� k�B�<����S��P�#$ֿKg�[�K�{�<��J�ˤ�:J��h���s�<�4�҃}nqI���4S�\(+��Tm�<����t��-k�'�0��bu��f�<�TDL�����*�8�-�$�Fb�<Q�`�2�X���W�<�bs"��E�<�& D!"�za��/B�py��A�<���=ZXQLV�w�Ց�|�<Q�@O�z`����(����AA�'	џ,���� �r@S�9h��q�K�K�C�I��Q{��|��!�J��"�
B��2�w��8���aa�P:'q�C��L���G�:2���B��� 4p�B�ɗ� is��
�!��iw�oI�B�	 69�0��Q��#A �B䉑,���1$*W#P��(���.�4C�	�c/���"-߅i�M+�*E*MQ�B�Ɂ,BWbKA�J�T^=*�B�ɉL[�yK0lƻVm&UriH8YY�B�I3r4���%�O&���`ҕ%��B�I)�ux��A_/�ju�"S�dB�	�ˊ�Pr���&P�@hV�?�^B䉾#��!�D�:	�h
�
&	5����xx��1Nu���E@$B`\��iKy�|ʟ�$I������@�GܴU7�h�7i.D��褯��#p�;�5p�:�@1k,D�(��H�0j<�so��0���a'D��f2^}����% 2cU� D��xF �>��!��%�L��%?D���$�"����� ]K�HG�<D���R�_� ;��@�=���Q���0�IVy�U��F{
� "��3�ҰG��1��.�m�"Oċ3i�/��S��H6WX��)�"O�*�mO�(��a���#=bW"O�I���������څ*|K�"O�)�g�SW��k��(�֜�"O�ӳ/C��U��'B�Ḉ�"O���`N_��p�äQ!Cm:48՛�����5����	�E"vXR�W�;�C�	d�i���Se�I�#M�k��C�	��UQ�/��)H�q*1#+�|C�I�B`� �eß��p�k���>HjC䉑Uw|ж��:+�p�����2C�I7gmr��'كE�(��@b1W��?Q�����(Ytl��O�/(4$;Q�N��!��K�<�y�.������]w!�$��EjRŠ%��bPV0UK�	4�!�\:,|�TKv4��g)�&�!򄙟<C�E0�I�P#W	��p�!��� 32��"JHEX���'ʶC!�$ڐE��`cHכ2�Ѫ�fM��<J>E�$E0X��Tq6�Z{a�Y+��yb�)�U�d� 숣; �@9�(��|����C8^���ʹ7�vt�f��n>F��R�R��펲Ku ��WƎ�z"�i�ȓc`v���e�+8�m���]0XĆȓi��exG�Ai,��+��D����$<ιIwL�[��=�WKXB�>mΓ�?����S���|b$��>�R)2�ޱ�٣�k�y�B^�f���(C�,��N��y���>a:`5����s�9h�%��yRS;r��r���s�����%�5�y2KL�:H�\!���"o(ԕ��Y��yR.����y@"�yO�9�'�
�yB'�+	9�8Z�6a����y��'�R�'8l4)'�ݫ\� ��3��:��
�'\���g��Dʄ)y4�3h� �	�'ty2�Fli =X�B�����	�'_����''b�Lu+UF�!Aqd��'����9\��r���5��P�'���;��3iPv���e�;1��*�'u0��wKK
��ɘ�LS/-�&���'D� �-��]��dލ,�����'�``�$^�3�<��D�2�bA��'Uf<"VO&���RV�\���Y(	�'�.	��*��4� ��B�&=�
�8�'re�G�B �假1����'�d�[r�{$��k�η'�r�A�'Lў�'��/�j�RA挸!��#Kk��a��X<*PI�K(zC\�8�f��p��܆̚'�T-"�n�&�\��f�
�aնp�M��hO�(�@�ȓ/�p-�L�
 ����C�/����Z��캀A��b�*��'~�����Voq@q�Ƞ 6X���C�J{F���%��Ya��VY*�a�K����z�b�" J��%ab21�S���@"OĹ9���2R�A���h#H��"O&��a�"}_���Ӣ��N�݃&"OVe�5CK�xKW��b��Ͳ�"O�`�V���O�-�0��%e� �22"O~�t�Z3p���Y�A��0��! C"O���C �h%�Q���n�[�"O��yP(:g��r�(�L��"O�d���Fh"�:�	�(���"O� t�y4n�&Ti���AD�:m�̤�c"O��9 螯B��p��lÙW��-�"O4Q���cl��"�b+<L�q"OV=��̊]a��8a*D���@2"O̲rM�/}��4Q"�ڐ��ES"O����%\��rm_�,[����"O6�%����9iaF�@jD��"O����Z��  �d��\��E�D"O��X��������P_I8�B�"O�-��鞧x�`8��	)Ix��"O�P1�M�Ԡ��K�`?�{�"Ot�i�@܆�FѱŤ�f;�d� "O�tp��X+T�����,�;:,|��"O�y�DJo8z�ŋ!r2$�"O�E�#�5?Qt}����(eGt
�"OI1�K��g�<���̐5T�i��"Oi��B�h��E�3<��"O��[Ƥ݈d��H��*�8Q)V���"O�HБ��4;��d� /@��mq"O@��a'7d�Q����<yl���*O>����4k8�H�� ��
�<Q�'At,��I�6Ts�节@����'����H
l(�K�d�"�
�'x��b�y���HANX�؜��
�'����1��u:C�Ӵ2
�9��'���p@�"����2BŠ!���i
�'�؀`�@:#�0�a�i�*�){	�'*:d�Q+D��H��a+�%%j0}��'�ѥ 3O�,��� s3���'�|u�g,��b: <�Q�=mw^�J�'��k�C�<j�a�)�X��F"O i�'�B<(����4֚�I�"O��A'4G�=��ļV�� "OP4���׼E��p��G��t�"Oxmz���h麗�G���#����"O�8��ȶQ��0��H�B8
�"O�(s�,j� �	'%	3�b|�4"Ov�;�y�T C#�(H���F"OȬX��37b}k�"NEY~�z�"O�Y�� v�P��ELjMV�1�"O2�@�Hd�:!
�;Id�x�"O8�r�.������%��&"
�#w"O8e���P_ڠ�����)�]�G"O�3���:B�j��F/_4r��p!"Op����V��&1"�#�w�T%�6"O��ٔ$I�P-x:%#)z��d"O:� QƐmf�L��k�4r�.��R"O�u���[�\�0�0�N6 ���A�"O.��gϒ�Q`�!�%�)��ta�"O��s�A�(�YP�	I�ʩ�'"OTX��
�~+�l ė�+� 9�"O"%�����i|�qD�*/�qY7"O�a;#��J������J��Q�"O~�B���f�@0Z�a�a�\�"O��
đCFL��O�i�`���"O0��VoQ�o胑Ζ�<�0"OT� �J
�+Z �K��J�K�<ua"O��E%�<	]z��T$ɥE��p"Ob���*b=�5�bV@�b���"ONtꇄ�WY�cV�/Z���h�"O �`P�XL�r�j`��n�H��"OJ��B��<3��#�ġ'zxx��"O~�"�G��T�����'	�i 80�"O���K��q�	&@?d~`  �"O� �swF�6vu:��Ȝj����"Ol኱����R����B XUZ�1�"O|ڱ/�|�&��)�8KDaa�"O��0�9��|jBg�I�~ٚ�"O2 �ÃQ�M�(���&Ǿ;��XU"OH��E1�X��������Q"O���5��8ЂҦ�&ċ�"O|����X#f��x�%MW�QQxd�"Ol��&�P��I�"��\L�`�"O�y"s�Vv��1����2%��I��"O�37��:ki<�VJ��1�؛!"O
i1��Y�I�윲e�� (�8�"�"O�,y,N�G#*�dW�V��"O,YT���w����
���,s"O^��0 �(�z�r���4?��m�"O���B�	�=#�e��k�i�t�g"O$�EIݯ|�V����D�T#C�'�ў��'���6#��5Md�y�?D��:@*��G��򇤊Oh,��e�=D�(Qrdɚ?��9���ՏOҥÂ�8D�T��Û�v�Z����- Wd���K5D�`���|٦�b� p}z	9D�4
��0.����ܱ'�R��7D� IFg�843��y"��>��i��4D��3�F0L���Q]=L��!.D�R�Ę���gGD���-D�`��
TV�f�3��h��k��,D��h�h��:�)0.\4�tD`��*D���P 8[�M !֙%ȴ���&D��a��&'U������7���$2D���SnD��h��J�°f�2O��=�`�H!l�P��@�Hl½*��w�<$X�B�~!�@��@|�=��E�k�<�u$޸X����f����5)�|�<!ae<�d��Tm9=<��"��^u�<Q�"�	j���1RDR�Z�f�n�<���5<P=�2	׷~��r� �f�<)U��rB��
�_�:	y�*h~��'ͮh�.�kMf<#U�+�X�x�'�f ���ξI�8�b 	���2�'\�0�+�,r��sA�j:ֱ��'��)�s	�T��$��/v��-"�'��Pij�x�P��$ct��	�'�@�u�,s�ĥ:��@�s�&Q�	�'�N�bֺW�I˃f��a�'��rΕ�8B�����x��͐��^��y�L�}NE;�GYX�Aue_�y��|�X�pm��ƍE��y�=+�B� �2V%���-�>�y�ؓ+<�M��;*����"��y���iƌi��� I|�B�I��y�/��H��:�IL9����3�E��y��$(��E�AL������y�͋�<����_%|�4�DO
�yb���x�PUyJv�9�n�2�yrkQ8,��2���#n�ū�H��y	;(�F�ꗆZ�%Z@�H@��y�,iTa��'��0tH���y�&˲)i�E�$���B�)�(N!�ybCIL`�t�%"&���#�y"B��
�^��˔6��(V�V�<���#d�6)
A��)���D��X�<��ʘ2P,e���8q��D�R�<q�D(Q`]h��ť?`��d�%D�� ��H�,�8?4yAF(E
&���"O��3���D̐��5����� "O�90F�Q��$� ��.U�:��"O���ĭ��n�<�����G��:W"Ot�Q@F�ohR"l�Q�M2�"O�@��A0:�F@#�*\)62,��"Oc�A4TۨI��)�&j���"OT��Ȉ�p��C��v� 1�"O��k�"N�4<9��_�nS�"O���r��KV L�A�˳:�%"Ot�P"�b�8��#�V�z`q�"O���h�kLū�V˼Q��"O���nCe�x����L>��8"O4���,��L�#��:�n�pd"O�P[�툪GS��)ag��z!�3"O&�єjĎBF��
e��&l��"O̐!�	.3D��
�T��Q	R"O�ɚ�@CƔ����H�1���"O�@F`ֈ#�z�9w~mT"O��ð%E�h�p�f�]r����"O���L/b�̓��Z `�tЦ"ON���L%��4�#�>-���v"O*��胴�Q�aaV]Jd��"O�����N�H@�0A�5"�v�X�"O���S�Q!贙0�OJS���"O�� s�/B��dQ��Sh;�� P"O��Y�"��l�>a;W.ٕ&h�X�"O8Q���;���豌ۋh%�-j�"O����DD:��P!��`bp"O"���V��P�~�*�� "O�@ã���E�~��R�˴
��Zq"O�`�AY��l(�l�e �Ip�"ON]�@l�/]z|�MN�	�2xs"O��[udƶ~�bqJ�]�3��l��"OX�C�ʖ'�t�RR�X8Q�Ƙ0$"OИ0 �>+���B����yHg"O�Ѓ�j��>�@�����_�\i5"O��Ԩ�0s�dX��N6��q�"O|�s�S)����p��=v�A�"O�!���q��Y��F2E���E"O� �)R���A�����t"O.5K����D)�b��:���Qa"OΉ"�	��G�"kR'�E�&۠"O�� �i��.��e �^����o�<�&B�AP�Bk�3��$ $.�m�<�V$
)B�\-h��1_ة��Fm�<�� X���ٕL�Xgr!�f�<6G�`��di�m�
;�$X
0/�a�<a ��8�J s��M�4ܒ}����^�<���� ��h(5�58)
93!�Av�<9ҫ�Aa���C)|�x�Dr�<���ʙn�P Q� ɣ9G��6�Op�<�q��+;�]��OНt܀gRl�<A�aC�1uU��Z�}T�xFh�<1��2�L��=a�$x��c�<����F\̌zU��;FH�#b�[�<���S�$�%7x��U���m�<1�ޤ|g��rb�8V�"e���d�<�
��1�r�$+M�*}��W�Tw�<���V�@�[��9�D�~C�x�˓���wd��	�hVC�I�UX��w�ĺw@%h��?JC�ɯo�
Z��qj���	'��C䉖Y	�]:5��,3�`�Ƌg��C�)� 4i�U�Ғ�4��F�p/
��E"O:QX�K�P��q#(��
����"OB���O��v��c�Q�aT!��"O�cL�G��`�2g�YO�|)�"O���cٚSuh:�� ;�JlC"Op)����H�P�9ef՟zِ �W"O�M;�ɲ��l	�����"O>�I�f�Sxd���[@��9��"O��� ��s��݉��X�/����"O�������/��x�'OQ�Vz�Y[�"OV���W/�� *0��*[i��"OʩJ�E�D�rS��{��i�"Of����97�����P����h�"O��	�K��pRT�w��}�y"!"OL��DA�&�ӆ
�!x��b�"O�B�-�G,m�&E>�'�.D�82'��OF����УtY�@x�-'D�����<d�`�2m�!.�:U6E0D���A���¼��tjߛ"r�R�-D��b�,��=$Խ��m�$Ϊ؃�D,D�\PB-��%W�-�V`O���d��e'D�lZ��ۻ �� 1�N0!K0U�Qf%D��#�M�& .��Yu�Q3%k�G#D��Rt�r{:�c	�C]�ب��;D��j��մk�*D�����qk'/D�X1Ve��ho�t���P�}S0��l D��aTeI>k���7���V�B� U�#D�$P�(�&INx��d�s�B�f$D�l`��Vq��a���[y�$�(8D��!�˚YI�����(���#5D���EƵ6���*H�bJh����4D����.U�S����ڨ@*�UJ8D�� �o�w~i���	jN�r�L4D���R��l>��P�ɲ�1��3D���'�=�xq��I�6u��\�(%D�P���)z�rq�bh�
X�s�F8D�tVÜ�#L=�s/
H�"��f(D�����ˮB>p}IG�� ����"D�X	�`�(I�h@j�J�I4z�E?D���ǥ��"㐤���:����>D�܁2gŞ#@��y� �9*]�Lr�;D�P���ėf���2�JZ�I	/T��[
ߛ	~��wD�1K�h:�"O���(��Z�|�֥N��j!x�"OFX �KA�SqP��7fN�w��x@�"OV��oF4]�)q�ω�qU��ñ"O����.5w�Tt+3OZ3=�("Q"O��h2�
�l�K�2"(1��"OB�8� ��F�t)�R��7��}p�"O�He�Ѡ뢘x��^'aٔ�"OD�0�,��V� �%d�%��0�U"O�TS��2F�t�V�U�z���"O��
�`X���9%kF	s�����"O��rR��ZQ(��S��$U���Bg"O�;�`�!<�)����
hv��H
�'�xy��,R�Yʺ]شj��H����''�hó��1x�$ �$㒆D\V���'�H������� S4��9_�}��'�j�Pp䔧;���s4i�'do^E�'{��p��$S2%+�ϥ���[
�'�D�e��-TR6Z) X�
�'{z\QDE̺LTxiT���y����	�'��94Oҙ
Y|Q�cyx���'Mv�"���J춤;1덥f����� 
���&E,L9b��G+�;f�0u�7"O�{��.^�A�R�R"P��l�c"O�����8_��I�b� �\�p�"O@���V;){>���G�I°�YC"OJ,�P�:WY������!��1xQ"O4�2��$� ��o
�=�b���"O�� ��!.(�; N[3�e��"Ozy��_24ut�mI5us��"OL��g�F=b48 �gLW���G"O���$��]���7����"O�Dk�`�?nT��O7�"9:�"O���Q�G	*�����^/?��E�&"O>!z0�S,�|5	qɔ��$�"O��9aBה|���R7(�$v�~�R!"O,|����MA\)"��nϖ��U"O�ͩ����av܊"E�6D8P�B"OM����#��u궣�?
��(F"O�K�%*t�D��5�Ǫ
H1Q"O�� �A�q<�+MD,s�С�"O�`é��;�������rO
xR"O�񸁠������e42CY��"O�|Y%Y�0 �9��#a� "O*�7�/+���wcL;O��qr�"Oε�1F�LO�%8�CZ$�|��"O�m�B��9��4j��R�>n�H�2"O�%;䢈'OlHG�2H_"��%"O��)�-��/Z���OY;�o�X�<���Y�8j%�\�[|��40@!򤌁�`�`�.��>��l�2"ʿ0F!��t�����*@,H���C!�<�!���K��Y��@Ɨ@G���.D�!����S����Ć$zx�c�D�3�!��ߩF��k!M�i��YfN�2�!�F6s	�  (�O���0�ڑ�!�ċ�Bx�5q�E ~�Y�$�!�$�.(#��ʞ6�$-S���):P!�R-\�-:�n�p�0j�C�9%�!��	�F����= ��l�  ��!�%+x�}2'�N�p �$Ȧ��%W�!�$�#���j �v�|��'�I&{�!��/%���w�R9ǇNL�!�DY�xj��!2i_!=�P�1GY�p\!�D�"��EB`�;8��Qq���{3!��K�ٸ��زN��8I���A6!�U�WU�jΆ�9�"��ҩ�N2!�1G$vr�ݥF P��H�G�!�DM�A1�r�L�W�<%�t)
"Ej!��5L�:x�E;mlM�D.#bS!�:�.���>8g0p(_�R�!�$ܕlI�����6Px��F�i�!�$�8o��I��&�:1����E�&E�!���(#N.����2{-��c^ )!�ĉ�>q�]9DH�7�(�@��!�$CK�ȩc5�[,�k�N̞B!�$Y�uņlZ��I�`�(�E�?!��<}D����G�i�(`���n!�$L�E~��{$���G��4�bɋ�@�!�Tq�� �J}�q�g�ڬe�!�$_�J�� rSU?��Cp�I�#�!�d�P�P��D���'�d��H�G!�:(jv)����k��H	B*90!���3Z6�9�����9��ʗ�Q:!�d�->�M�G$ֶ0�<��W"��!� 7������c�d��`�<)�!�� ����@Y�(1�Gn�4%���R"O@��G~8�LBUŔ?�؀+V"O�(z3H�)����E'��9���kS"ORQ�7�R�o"~<b�N�P��x�p"O��z��٥o�td����9̨z�"O ��i^�W�ũ�KU�+�����"O�@3oG�a��T�˷c����"O|])DD��+C ���K��8��r"OJ�1���L��hS�G�1-�D��"O����i�?->��b�#���"���"O@��0ʕ���+IP4f�\�C"O�@J�N��C��9���M79VR�؁"O��L�}$�0zt��$Nr���"OLx{�e̓X�8YA�҅62�Q0�"O!hǋwKJ�-1*�Ѐl`�<��A0�qB��j���PօS�<�"j�?w�!R���B���0�ZN�<��bĺ�j 1U��w"���&�M�<GƎ�<�R����
�"=���n�<٢@��U���J��.�	�l�<q EK�bx�MC2h�'�~̸��PT�<���Ϻ]��9䆬H��]aQ�<قH��hK��B��%:�Xd�
�L�<A` 4�*�!�ڢ����
F�<YC"��?���#����1��ƼC�	�DITBΒ
��q1�ͥGj�C�3X��ʅ덒0�z�e�FB䉪I���%&�9F *�NMk��B�I�y+,�c�c�1%�Xȇ��S��B�
����	�zrt �T�R��B�ə �t�cUɗ ~w,���ƆO��B��A"h�
6�M�L�b=P�F��
�zB�ɐ E���(:P����״D�dB�"bc� Ic��v%U+7�Q�jB䉨a4�����Ӑ\cҩ`�F�5r�vC�	af~���'Ҋ]���B�A� '+lC�G+T�jg�
=���I /t(C�	4����Y2Z/����A�1etC�ɓl�h��&��U�&�Ц���T��B�	0+�a��b�+Q��d2�h_�W�C�	" M.�2I�<)��t�F��?*?C�	�ΐ�rǓ8����΋"qC�	�^{V���j9zE�$�'��;T��B�I�U��-���8->D��!m��C�ɪD0#$b�����X���	B�	4!�Ɛ2W��z�"�I��R)y�B�	��t�D�ŭ,n�uR�Su~`B�ɀ@� ���6"�v(��#��1&B�	*��5#�LEG 29(D4h$C�I'Y�H����>y�yI�C�8>��B�	-Ȫ�e�G��`���3�lC�	�8WΜx��T�z�$ fQ�}րC��&$��!��J�]{~�+��44FC�WtA�tE�0N>����ʾk?�C�	''�>�PP �&R%�GLfJ�C�ɭ 8%g�L�IX&a� K�*ТC�)c�:�"a"�i��`�`�/&BzC�IжyQԭ�Y>����&�a�C�	�P�� m���N�5M C��%T��$��С�@���B�	R��)��4����	F��RC�ɣ2���k��B4Jy��CʼE�C�k��QV/Ά/*���`�ڳm�B�	�J�&L���y��)�^ݖ�2��� .y�f�Ϣn�(�xf� \��=�7"On1q�2F����#��.�>�{�"O q�L��8\ݠqCI��r��"O��i�FL�Y�x�PQ	hH��2"O@�U�v\��[¡.2}�ͱ"O4�bB�B�x`\5iFT3eh� 
�"O�5UL�o�&]k��N�Q�4s"OD�x�wzVY��� M�X�Kd"O�郣�E�vw>���ޗ?�0"Oj��b�Ӱ�R�$���,H: �"Ol!;���8���B	54���"O~aZ�gX�&�\���΁!d��d"O���j�>�QF[����"O�L��!Tp��fLq-��X "Oz�ؖ�W H�Ԩ!!Sb�t�A"O����1s�d��7ʖ-|�i�"O�i[�`��}0��2P
;kd�9�D"O,,�0f��u�(��YI���1���]�<�4�ݡ�������ŰtY��_�<��q��)Q�ㄋ�[�g�W�<��� e�.�r���1�J9c�łY�<1F���l�~�cGS�V�VP�ȟK�<�JǼ:��W�T�n��$�b�<1 ��k�4��6�ٱ/!�K��]�<y�kC�}�^$J�fC�r�h�*Q+�C�<�%MN�`�����O)2��:�O�B�<!SJ���9B0̏*�W܃�!��3�f�{��\G������i�!���6P3![)N5<�jb�P7d}!��A 5Vj�0�*ϹI`� 4� �Cx!򄁞}����5Y��:��m!�č�*��-yĥ�C�Q�ѩʃz�!��.��!Zt�{1ve�e	�J�!�$��C��A����m}̸��@�K�!�$�8HO
���6;�N�Be�F�!��y���cՕ5��c���s�!��3sDPhA�
)�*x�S#F%@�!򄀁"�������/�B���"k!"O�uA��[�-2p�SH�z��X�"O�hpA	U;���h��&��@3"O�t�s��-"J!ק�s����"O^�:"N �n�`$�s�ݚ$����"ORt�� �)��2�dM/9�.�:�"O&�(����&�|͋��]貄"�"O��i-}Jt��!M&hE��BC"O@�u'.q�tu�3��3f�bd"�"OzQ;WL��Wю�@�ń5,|���"O���d��o1`��"�ЦU��rB"O���Ebͻ
͒X!�"��=S�(�a"Oҩ���J�}�rL�B��&N<��3Q"O|P��H6$�`-�v�L� 18�"O�+���`�,����K���JW"O@�Ш�&xp]Qpʛ)~�l��c"O,����+q�ܕ���B8P~����"O�|	s��>9gb-ש��	m��v"OzY9���K_�ʆ)W�#^^��"O�E
�*Y"ew�(H�)�>D�r��"O�0:��Z�P�N�i0g��9ɒ,�r"O E��C�?E��P�'QY��#"O*d���>�Z\�t#ԈJ=Hհ�"O�I����e�P8(.��"�"O�R#�����1�	�`��AS"OY��AT�fEr��Y�p�`�"Ov���C�z
��J��B���"O� ����h�]!�ϝc~j�ZS"O>��@d6%�P)q_���qҒ"O03�ƃ�r�~$Y挏4��T�1"OB	2BL�T�8�H�+���p�9 "O�}�7o�+Q7�A��gK[�0�C"O<p$��3U�;&�_7^81�"OZ0��$*D�avAOt*s"ODp��%i�N�b�G;BH���"O\0s��ۮS������r��(0"OĬ" ������&H�-�|j�"OZ̹�H�`�ƨ�e%G�p�h(R�"O0Y��%�
�Z�B�9T�eE"O.��CNB$0'�-�p�J	$��*C"O����	Ɍ-��XT�X+Tl�4"O1Qc됬����HJ+���s"O�U�F@��b�a�]�=��)�"O���d��
�0���ˌ�� Ik�"O�0��*�\�9�jCh�dm��"O��(��N� @`���&!���@F"O�x{b�_�G�a�@A/ ��x�"O��HRQ�v4VdJ'�H��(|A"OrpZ5�؀z�0�+�Lӷ*�N��"Ot)�m�0���+W�|���&"O��Z�b��p�$�Q����EG��D"O�r� 6d*H](8���"OD4Jc�Ϣ��]#��]�l+��z�"Oxx�	�G���)�ʌ�F+~��"OJ�@�h�����dg]�_FQ:t"O�� ��Q
E,��f�-<���"Ol�yp ֌C��d �υ,@ks"OTX��!޶ඤ��F�X�У"O���faY=}��)%$�0��g"Oµ�C�	uӖ1s��U�\z^Pʶ"O4H�@JC�b��8���4Rt�q(�"O�ATfOa(d�1��0\Y,%Q"OL�QF��?hLW�:�Na��"O̜���n�����#F�s��P�"O6ep�Ѫh[�Ȫadڽ�Z�X�"O4�+�� ���1�6+*�t$�"O�:rc�5T�@)�.��і"Ovpf�i� ����j2�4t"O�i�&��)�V� �Ǝ�O,��@"O<@�b�h�>���.t؈K�"O�!�%CۗI�PD��DˠhNTyt"OҜ��J�3~Л2������x�"O�5�T�ب{��|��҃G�|;�"O�8� 䓁zn�%2�i�μ�8�"O
Ź�K�<����Pd�<W�)!�$��L_.X �C4p���1O,M�!�$����H��oU� j�xS�L�7f!�$F�|  U+ �6gT�D�w�Ш~L!�$�:du��Wlכr�5��˄s!���*���S�#y&}"�);�!�d'.qʁ�e
�z���Q@�!򄋙bṰ����2
E�a$ɒn�!��R��ӆ�='���SÕ�!��]�t��L���ߞN�|US�H�x�!�Ě�"~<H�偍 c!��:Uȓ[!�$�R~F����`s�M�
 M`!�O4�J�ݟ#`��e+م@J!�� @ژ��P�=T���Հ�jE!�D�|A^]���[�x!4�ҡ���!��22΄t���9x�B� ��_�!�$\�-������4b�B�l�F�!�� 8�C1��]Ji�d���.�^�1'"O`š���z��#�ጐ-�i�"O�x�F�ݭq�VA��1y����"OH9
c���RԞ�ƀ	�[iV��E"O^�DGw��0��,Uz�r�"O��{2
ܲ*~;Ad	0R� g"O��:��@�s�i�$S�$�(ԸR"O��d��yQ�h�rcΖW��u"OP(����*ά��FB+V�8@{�"Oq��g$=���P���7�d ��"Or=z��[<1��a� k�|��{�"O�I��J@13���'B �|Hw"O�H*G���.a�s��ģd4�Røi�ў"~n)9r�-yQ��j� i���,g�C�ɢo\H!CB�	;6K��`�>t���>�#@ף[�\m�U�!<�<x�qk�u�<�̕"z\Ce
���!�EM w�<i"�������F�f�����v}��)�'`hX����	i�@Y�G�H�R�\��&�p�%K��g��r����9D��!� 'U (�B՚ʪ�8D� [��43� �BQ�'	�z��%nw�ć��!'�> ��C�
-����b4 HC�I:)��H0d	?^���jw���E�&C�	��B��R���W��Y4בp#�C�I�H�lP�Ϗ?��h�i� 4�\C�I�\�,ȹdHE�Z�����&JfC��:��Ħ)�Tj�$Wf�C�A9<���J�B0�&�բ(_zC�I	�<(�i��2�����#�8�bC�I%k��<q��-JS`��"π�&C�I�a�4 �-��$����<NC�	�9:�h��2���kZ*C䉫rS��2eC��>k�	�C7}'J6��5�(O?7�X�i%��#��ʾ��f��2	!�$SD�R`݊m��y���R�I{���a�O�?��(B��#Z��>D�x�6�8F�,Y���U����;D��+���sJ"Ha�I$|Ű$e;D�Ċψ���uk�l�8ӭ4D�Z&`B�%��|�VE+	VX ��0D����%��H��v`L3@��W/D�L�"�!Y�`�*Wd��@Dp�M-D�t�"�:���@\��x��.D���!�K.y� �ؕ� })�Eu�8D�Đ�$E�v5LzP�<Y��Q	Ї,?����<������ٍF�&U�W�[�m�B��&z�<��o������@]`�<xGz���#�F	��@ƍ	��a��&D�TyL	����%%�5l
t�bV�2D�ۃ�H�]G*�A�ќ};��[ң;D�(��V6���s�D���h#G>D��05`��O�΄�dׇ��@�gJ;D�IjN�Bg �fly��N�Q��C�I�<�8R�� nt0�bi�d	nC�ɾTm�i�4Ð�*�*�ar"O�_�C�xi��%�$L$��D�ɱ2ƒ��+O<��$�)�Xls�D����GW�yay"���e��x�4.B�8��uS&�ڻSͦ�1��!|O�c�8pP�?y;J�I&�}62��D�?�DPQ���Oen�z�!Ǡ�$��p|�P��'�h�Kd�X�dD��S�=�'p����Z$-Vr����I����'�U`'C V:�@Kb�L'���:�"O� �M��̜�J�uir�����'jqO�@��k��{� `J�,Z�\����"OHu��)bt�̀�	k<D!;�"O��!ƣ ���xu-�4 Jq��"O ���W4E�$�C�BL�+�E��"OZm#�B?t^`�B�a �hȠ�*��'@�O 0���OQ(�����I��A�"OV�����?���@LоR��S�R�pF{��)�*	<=��J�4#�^��c�7�!��]�Y��0�A����@�+T��hO񟴄h#*��!M�"C)]!p��-�`"O�q#CF(ԑ��2qM$�J4"O���hHV<tx1��}�t�'��OʥhÏ����m�C�ˀ�!"O�!#�;,d�т��
5h�V��v4O���DyrE+�S���I���A��(rj ye)L�y#t�Ҹ9��B�i��8���2�yb�9mU@�P�Ǩt<�=Bc��?�y���b�2 _���ugX#|o���'��)y�0<6y�Uq�8�A���-O�Xa1H+j�����M�P rǅOlH<�ň�w�ڈj4�ג�d����L���"�}�@E�H��1���B"�n��)�0>�K>�*��2�W�'H�X�L�<�ToՑ864+F"ք��H
�p�'�ў�'w�,Mf�H�  ��n�rlL(<��[6w��H����&s��u�t�:jgў��'�R4b��`tYSf��� �޴�Px�N@�S�"�nơ+&@qiD�B&�yZ����W�t��]��(ߞa�21���e�	Xy�`�&=��R����\$��	��yrׄ�<�0��L�4H�A��O06M7OBh�A�Q�KЄI�gRf���W�8LO$-��K��)�DF�<�Db�>y�XT4��djL)���q�D�x�Ĥ���J��2���S�<a9FcK;'�І�FY�d2�Cǥe���֣6a�>�ȓbA����P ȜP�Ɍ�,/v|�ȓ>�K!&�,k�E ���P��؆�dU�<���U�3���bҀ( a��Ne�4�"fT�i����m��u�m��w�嘓̐��1�o��a�ʤ�ȓ�¹�U&�\�HC��7 ̠�>)�m�p���'>D�cBBU�p�JŰ���l��݅ȓ��HNM`��c�4~-�q�)�矰�gό�Z�rŘ�N�H��@�;D�����,����Ͱu�xY#Nx��ᣟx��'(���.Ɖ\&���1-%6*b��'R�	����49N�%��+�'�`,��'���	Tܞ	
F���sϔ�@��OZ�ځ�Ȼ��Tz�$f;�"O ��D��"a���ʣn�AKQ�b8����C�o
,�����0V����B��`{���ӂb�����
�8a����m�C�ɸWt=��䂶G0���lX�'4�tϓ�p<���\8:Ei�K��r�,��� !�d�QB�ȡ�XWh��������!l����I��1�c�\㟐S��"U� QZ��ź���!�D�O��j����W�@��gO�5:"z��x��^n��u��|2�K�=����2m5)k�9�W8�?�'�
)h� D��:L�� -
�6l��'V�X�j/T� �8E�;X(T�e��<!I�lE��B�d���*�'�)7%������&F�bF�[6K��:UF?Q�>��S�? �H
Ḧ́D$�,�h,P���8��'��f�x"�]�<G�i����6�`�D,�'0ў���	R����M���K1&�}a�p��'r0�<�E�U��؉PF�3x�æE[a�<y��EiX��rgKV�\��D[�L\~��'C�Ub�Ɗ�^�t}�˃�^�4(s���ԏ;�V�G�
I�v��Wh{g�	ğ�?���D^9F�p��γ6^�9���Ӵ=�џ����$xݵ��c�G��wDI�_7���ɢ>цH8�hO���I�C�u�V�âʪ	H�=0�5OryI����It?Q��L=s	������>;B�X�!X$}@!�D�t8XC�C�)�����Q2��[쓊ȟ�-��b^a*�IBR�܎@I��`�"O�c���){�	pì�G�,I���O����'*����p�N�6��qF���;d	Uf<�������U��b�Ȅҵ���}�|�����q�<т.X�%X�p���".��zQ�k�<	� �h�ҹ����r�0Tss.CC�<t�J3A�\�r5�Ұ���0a�J�<���&�@�F�r�Vtȳ�H�<YЇE�w^�x���7<��	T�Sj�<�B�t�d#�cM��<�r��GkN�3g��,� �@�'L���ȓ:���U��*(�T�C	&GfX��(+�	�SH������ I�t<��^)���"�	\��,X���%4d���`�V!�a��d�s���G�jq�ȓ,��hR�C�1w��0�T�Q�!��ȓ|�$�rK\&A̤�䟗EP~h�ȓ$D>�9��@�xf�f�H��B��ȓn�hHAa���z9X�B05���WԉK��·v��sq��-m�h�ȓ�~�ʷ&��:���Gǩ?��ȓԞE��/�<<%�0�٣%����'���R�6�&P�e��~�����LR1�J!
r!�d,�����"O�EH�
Y�5��T��`U�4^���"Oly(���6k�)�O�;Sr���"O�� h�aZ&���ǳ4��B�"ON��L[2���
�0+�Y��"O�D�g@EUt ݣs�ˢ$���'eT!
b��%�Ԣ��{��l��'���䂡b3����NoD�[�'v"i ��,X�
O�!f�J�:�'Ju���{k���.�#o!��(�'`�(KF(\_����ȋ�i��Us�'4 ����E8�gE-hy���'��R�c�>�t���d�`yc�'H�i`l��p��U�F�P�'?"�(�D�-ye��5��V$����'� ��NQ�l9D8�Ӽn�L��'���H�Өu��ds�ς���y�'���HP=�I�nȮʊ<��'v@�)�[�aV�l��,�;"ܔh
�'�ܭ���ӀDd1	� �,�	�'���m�'M�TErF�8o^Ր	�'�����K�d� r�S�a%�� 
�'�|a��A��/�>�𑀀!O@j�j	�'�fl�퐊&��ٴΊ�R�H�'4�]�6��5q~i+w�� ^��	(�'eęm��D���#I�&i6"O�@V�
9�r�[G��.S�	p�"O���F�bw2ht*�^�J�9R"O��kO 4��ě1#�:����F"O� ���va�/r�굢�؀n�ɘ�"O^�A6���y���c�/���� f"O��JѨ�����9! ~9�"OT��*�?�����~�R�Q�"O��0/�'U,=��R�UL�"O@a����9j���E�P�f�B"O�$� �8pg�2P����L͙�"OZ���M��0`iv�L�cQ4��"ORLB��?:�	¡ދr�j��a"O��2���A�����^$k��"O�5#�P�U�N@8�M�>f�v)Q"O���G�R0m�� +��׎^'b�F"O/��XJƍ@!w����A��6B!�K�ZX���j�>|��4r���!�dӴ)��i:�!�����bLG.!�ZU.�&J�:)��Y��'R�&!��͡ID(�Pf�U�`%�o�!�䎖L3�}�a�(N��u����C��O��|�L�w��̓�(8Y؈	@Ɨ���d6LO
�y���2�($�DSś�f�V���dVr�� �;�ܘYg�͐m����@�'���S�M�k�"��g1n�J�'�v8�b!�#�<���˲]3��&��G{��t�ѫ*y��y��N ����@)�y�(�	�(�b��Ɛe����)�y�*Z�ܛ�!�(�n1��Y��D��a$|��$/�M ��S�DM�l{�d٢"O�� ��%0%��ئ}r�8ZS"O������X�<̳����J�Ȕ"O��I'"#��3�Y���A"ON����\�̀�Lţ<j�l�"O,����J�UR��"."6��R��i>�k��(/�[L��a-D��A�@�QP���T�!�@,ꥄ*D�l#P"C���|vm� V>��$�2D��pR�ղ^~x��@�JR��S �>��M��"i�H����Ĕk%���Ɠ[qH�ر�ߤ"�qK�#)���C
�'�� �B��0*Z2A#��4zp{�|r���� #a���Q �@K�a�"B��.���V蒷>>��W?q����<�����f	iȝ�{C�UB �,��
�O,����ܣ3 MT��<Q��Ih�!���\En"��̥����u.I>0|��K쓱���S�	`��d�[<x��l󕬙�QF�:�S�O�z������ɒ���b�bi1�\���	������D� �g��O�>��0@Ѓ.�t	8���$H��c����jӰ��a�v����%n\�fL���a�OP̻t�)ڧy�ȝ1@�;4B%3�����}Dzb�i�]�ɳr��$ju'�6�	4�
}O�c�d�_����D랣I���s�mǠUO�C䉺Ix��!�`!zPDcBS~tC�I6?�Ѝ{�\� T���AJC��,N�T��Ȅq���@���C�ɍ`�Z���!I!wƴ� ��	�O9�Q�Ɠ8����S �)E��( BL�3�U��OԠh `A(�Z�00���D�h�O"�	Nܓ��'v��P�C4-���Z�"�)f�h
�'�^�+@m�HJ��s)X�[�nY��4�hO?7��7e�&!��.m�>�0d�ƽ+r�}B�����.ؽa�n�@�U�Q���+4Mf�����Nx��� �m���/l.Qx1ƒzb���ɗ]A�'pԥ����AO:m$>؈�h� _Be+�"O��;�n�1(���� B0%I�h��Y��� t���%��m}n�#S�ܾ�<��"O�%�wi6`J0��CI���H�"ODX�.L�(��C�A�!Ui�}��[�D�O"<�I�t`G/˰�ӥ�3�حS��*D���Á�W�P�*�Ɍj������>AN<�,�i�<�O<����~��(�
9%�
�'j<�i�Z�49�iY-�
l�J>1b�'�4x���'4�� Μ)'ְ��	���~�.Ȝ*�	AV��`�`+�D]7�y��'g���q)_(e��}Q0�\�J��v(ړ7zў�]>�ޑK�nQ=	x��D��b�B䉶�2H����!�ā��b�j���hO�>��a�Þ%��IS	�$E���u-(�O�扣c�&X�T�T�����ьK{���O`��dG0iwb	IG����0!����!��y��O�O�U��CD={�L�'���Y�ΕЅA�v�I`؞���o�"vܺ#���.]^�B�n6�	s~r�'cn�=��C���~�P'ǟ�~��]j�M�$ݐx�,�7Sʠ3���xC����G�|�j˓���-���ӢRj�PA�"����-Bd�<C�ɗjΞӧ��k4`#D�;P|�$�)�矈8��^�p��y��㌴���-D�(��`_�.	�0�bM j�$X	�@8ғ�p<�Bk'
HА��X��}��B�n�<ї��$q|a����@"y�d�b�<Q��n�T�w���okr(0�Nb�<�e *V�@����t�v�#�l�I�<��@�V7�p0ӍS�j@{�PC�ܰ=Q4b��K���C���[�XB��A�<��m3D���S�v��i�'�Iy�<a"���D��`�#*ƛ.��)(@�<qE��.yș����^�� '^z�<���lu���є6�~���bU^�<�c�ݒpF|U�#�n�89�"\q�<I��*e�>aխ���9�/W�<1S��Sy�p�'*Q�P9P��U�'��x�MH�1c]74��P3����y��9a��L��xgԀ���X��MK�D�[|��bL�	xxm��P�ТC�Ɋe&l��Sǚ5v`\y*RM7�C�	�ێ�'�F5�� ��F��C�ɣgQ��P�����a00j��DþB��j���֧S�.��c�W;=��B��"s+��R�W�x@v!���w���p?T�D�:�F̛w�W$}ŞTjv�k��i��O֓O��K���]����[���*O��$�
�"H$,I/&�,Q(��Z-\�!�$ �v�B����Z6�M��ƍ�!�$O�<��p4�ЙD���#�C�Q�֢=E��'&Jt�F�D'GP�͐#nU�^�I��~B9O�|x#�6F�5�7Gݶ}�qs�"O0@*��	��ˆE�,o�ݹC�x���P�I"O.��዗wjhX�QŎ{��C�I]�=�bߡq��1j�'�<B�ɐt|	Q�k֢��=HJC?AM4B�
0���b�� ~4�����\:B�I���C�@F��x�r�,R��d���vw>��F��f;P�r�L6R(�Gy��'��5RP��z햹X5��gs6ఎ}��)�\,3��X�t�	?+8:Y��
�!�ąm����w�I�'.��#@O�o���J~�'Bj~J?�J#�ʞ�pU�@�c#��/נ��(y�i��̼G��ԩ#e�=l�Ș�����$ �O>���%
!9(̔97R�&�lԳ�'<b�� \��m�x7$�Iu��9� �	d"Oj]Rg��~������6<P�`�$�OtTG��ӟ��s�Y�o��X��y,lu�0"O�C��B1ujഊ�f
 L*�sӉ!?��g���)��$ͮ�\�9�N[�2���/��^�!���v���#@J�p)�C0��)�!��қo(����@̍&x����VY���L�	i�O�ԡqJ�`�f�s�g�؝#
�'�,� ���+
����"6]�AxI�XK�'�ܨ�� ;�NQ� #���'���Cv"��nkĨ#�%�����	˓�(Or)s��Bo�2H�i�]F)�"OVl��m��,�&�c�� �4r��>a���i��=��a���f҄1�n�c�!�G�Z�$ ���P@G�Q�a�!��H�����Ԯ��5w�8��*m%!��\̀�u�7g_�D�f�\O�!�WaKv����hU�<Iӄ�2w�!�$ںMց�$ ��fS̕�Y2�L��''Ⅹ�!׆7�*��&��@I��'���{Wlͥ�vj�(@�r�غ�'N~PDd�^��II��������'�Y�d�Z�!I��#1`J�f�`�'c\5񇊘�&�-)�h3u4�@�'�
�#�φ�ܩ;Z�JJ�'ܙ��=>7�9� ����Nh��'�8��D��/.�iSa�m(��;�'��)� ~X����1f'R�2�'�&��������2p	Ο^��a�	�'�b����h�1��NК�
�'�*�%�;~�p�t�]<2�హ
�'��82Lߛ;CL0 4Q�<�N�z�'.ʝ{BU�C|t+�,P�5t�c�'�
(!��N 6)ò`N;7~�{�'Gz��&k�p�R}��ɞ�%��)�'�*�a7��	fqP�����`D2�'��9s��074(
���>uRQ+
�'�6�I���PL�9;D����0
�'�j�JŊ0V8��T�"~/� �
�'F(���ږ%,l�
Ԋ�j�.8��'!n��I������O���;��3D�d:u"П<\L�8�ŜfM��U�4D��Yׇ��(Vd���[�JN��A2D���ߥ)$��c,������W�0D��{�$>_>���]Rड'�;D���p��.����q��4���);D�\�3͘  ��s䔗Z�t)h��9D��33�œ5>��!��ݬ4�N�i'�"D�� �Sl�d���%�Rh �!D�� �-��>�RV+�5q�� Ǫ=D���cGޟs����PU��Z�h6D��+����R�<E��OҜ*�։� M6}"G^'>Z�k��[�zjj�+��U$��'f�aٔ�	Sf�adʝ*wxRu�
�' b���/^�6}�#fސhMbI9
�'��1ƅ���D��G7(*Y��'�|c���5��)�H	�'�z���'����p#ҧN%���R���A�'�*�I�n�h�����LM�$�
�'@@��JРk>Z�Aǔ�~��
�'u��xg��8�$�*D:v���	�'ޒ�[w&F	�^��� �8rˢd��'(�A�˃�Ό ��S�vYT���'�k�`�(A��)���PX���J�'�H	��Jc8����:\m�t��� ��R�&��}�U
��O(0����"O��a��ܔشF@;D�̬B�"OY�eO\2�,���Ȥ7j��1"O��4D�&Rj<�P��6 �t��"O���l�1;�$��EL����"O>��V��r��:e�J�J��E�u"O�!:�%��m@biɣW�ʐ�g"O8qAF�-!<��iʪ�R�
�"Oڝ�I�P��$J�Oƅq�~�H�"O�#!煀#:vyQ�@�;��9(�"O� 
$��]N�pӉ��!�h�c"OTtAch�0O�4�kD�F�5�z�z"O�<���Ͳg)���f!]��@"O�Ղ�����0ɻ��ԙx�PUR�Y� �4�N�8hG�����#��R0�O�����0�#C�"^�0��omab O�O��"O1y@�'|���@�32�L�{6�$	t̠B���(N4�"|zM�'��L�C��
VB��0u�GV�<�t`�U#ޤ��	B��1���@�H��yeB.��(�'n"}�'���XW��)'�X��Q���		�'�8��Sn/����W�}�S�Ӎ?�u��KȐ4���Q?,Oԝ�#lȵ����؃h;t�.�az�핝�X�!�Զ>���1V��D��3��4��,�V�2>�����d�i8A�����'�Mz��-�ɇ&�UBV�L�6�&��M �q�8Uj1^� #P�j0Ð<æz�"O���@ʢlSpbʁ�*��B��J��@a��!�����8)�z�*�h��q螜yB&8�@*?Q>�Ɠt�rL��	�R)��i�Z��:�����#+�qU�YsӲIk,�!�0<���1\ \)ْ��4l:�Ku�THx�,�ҬG�0e,�#�JU\�k1燦Y��9��U!��L��Œ
wxl���\`I�v�0T��5c�U53d.�$�0#+�47n8��0ŗ�h��k�C�'�n��¢��Ha���=F1&q��z���d�<�\ Æ�ʸX�������I�4�{��ĳn����U\O�'��A@ArB�2�z�YԀ>&��*E�BTz��'2P�S��*?�r��D'SH��Թq���3� OT�B�LNUQ��4�,���'OEy�	L6�:�@7 �wG>f�A�.�����Ħ9k()�E� a�!�]>;�>dsPm	�L@Ph��h�/1�'ATd���+8�����B�О���I\�	u���Ř 42U�p!�ě)Z����&O/!�x�3��Ǌcm���u���de��"�	W�#z���3?	���5rx���L4&/�%@�'KP�'�U3�GQ`�Oڙ�d�U��^�ꖮ�H\�����]�JR-!A�,m����eZ\8���(�N���ʆ�
�}?�\���s���$�,n,��'��6U����&����*$B�u�d݋Ū�_&P��2a�����xK�Y���&#_��! �C��Q�'��ha�D�=���l~������|�W��~R����ٔ�v��"?^���I� 9N�V���l(c`;.��3�U5aHb`s!�3 ��2 �@y��d��~�]
4K2uu�"5�H��hO��z7�̑J�J�k��t	97�Ȁ1� L��0�����~�f��p�iR��'x��놩
�+%Pe0�\�D�h���o��Hڢ�Ԅ@��ӧ�O�j��T���yUg�g��u�d^�rg�,�ȓR�N��aIA ���Ha�Z4Z�Ė'C
X���o~�`��I� ���ɶjK	dS��B�A�c����k��[ ��(��(B��x��s�8G�20�
�'�Y���"F4�p��,B:�����Dh@!���Oq��p�B��z������F�H�'��
FmW��$i�e-(D��'�r�`�뒗P�ɧ���P�
u@���/�2p4�9Z���
A���%˔�yr);)��a{B ���ԃ�+Ǉ��I2r��G�W��$�J?D�O(�"s/2�Vf�#ʔ�9�Nһ3�L����n�<���[_>="��w@X�	1eP$m@��S� c����UY�~&�,��� �p�pR��Tx<ĺ�'$��A��%#SI��M�I|��СϪ'Inpb���%"Ȝؤ@�N����ƈ�.kK�p���:(Ϣ���8�$ϛtR�MyI�$	d��0� �"�
fk�9b� ��Y�\�1@�;��׃9�К�"O�4�3
_
R=���L+��q��s~��-:�@h��NawR�caZ?�����u��Q9�Z0�	��!)�� �`�!��ѹ}�Q�'�C�$�
�ñw-du�$o[{�(Р���?i���%O��M�G
���x�V�z�t�����3�X @.� �0<A�L� 5��	��<yO�_�:�9a ŐPb��H���Ǌ᠅�KhB8�d�81V����3}�hՓ�$�oQ~a�d�G"��ٶ̢�݅:���$&d:d��ˋ%p� "���>{��4�`�ڴ}.��9B*gFN�i
�'|<m���]�++�`��g�(��gSV~T=>�,}�3#�&/x>��O���!6i���yǉ��D�ЮOL��$
���x�)C�NL���9g�>ݠb� L|X�/�'%tO$�:��ߊO�N� ǌ<�əu,l�O,JX�԰Ci�ZҲ�?�!�=�<I�3cN�3�h�'��Ph3,��>�xG��T�O�<�U!Ǐ,ڊe	��.Z8�YÂ)�P}Bl��~��ڗO�̺��ӓE�@�
�B��[���
�����`B�I7w��:�̓ m)Zy�S#U�f�\#_����'+Ra��cԠ`���O���G�E%`X�psB�L �)Z��'��|�Q(ܴɚG��tQ (�Vg��
�t�Ѳ��?} ``7�'�qd̚	-pZ�j�-י#�� �����`�TT�s��j��4�tE�?�Q��W�2�H�R����U�d-�>B�I(MG>,*��.Q`�p�F P���~Ez�bS�&3`��%�ԧ����}��s���#��(�
q1"O�5��Ǳ77��p�bJ�7E���ܡ\�|k�+�+�$�r����'j`�����`|�y��Мk�P}�����㇝�w^�6iC�r7�8�r��=$��Q�h�<�!�k�d�Y7��x@��)��U��]D'�)`L�A�&b�R��O�v0I��w�z�I��@��)j�'�T�x!CJ ;�Z�F�3G��d��O �*��g���rM1�'}Lִr\?�BTCB�'`5Vd��/@@!�'F�-I�ɒ§Q#z)��/�(8WI�=m�:�"e�[�ڭ��IԂ4�J�[Z��@��o����ȓPb�!f(ԙ ��9{�^�%}�5�ȓ&#�	AFf�vM���Po԰��@�l�36�?M"���ץҬ@����mQ�̚���1H��Is�ٮi�&���'4��Þ�MH� �a�H����B��J�ˍ
@��%��iҡ)�vt�ȓG+��!�P�E�I�!Μ�:;�i��D��1�f�~� eء��u�^E�ȓhQ�e���`�g 	<p���G\!�3��@�ʱ��`��- ΰ��_^�m�1ɋL^x\cG�"����ȓ+q�ܢ��ɛ2/z4��A�T�<�=����*rC��i2x.��m4 X,	�T�ѻv�!�DU���kv�͗jS���a� v�^��@��g���q�q�;��=95���Hlj!M�Y� ���i\p��DX�Ė�
��l��C�\�#��Z�����@��BJ�a�D�SiF�X����dT�� &�b/X�����?m�1OZ���(�n��H�'bz�aV��{�T��OT�b�@�cN��K��]�?E�'�T�SJ�	-FL�)�G�*����k��?���̓Cx�A��I�W�b?]r�#u�19%�g<�x�c�%��A� 3D�X�F.��#�+LQ����gˆEb>5��A;R9��4e�Jw�P8��y�3��'Z8\�ܕf�N��F�	4���	�o"nD����^�Z牠W,pU	��AV�}&�_�k�@�BV�6<�9D�'c�Eq�FN
U+��L�#	�tS�:&�R Ĥ��b�"�ɀð�ۢ�%;��@�`�>-`��ʺ�u')�%���I3�O�d���{��/�l��e��7�� ��ɮP�~�p!+�� �e��=J<��Z��F��$� Z�$ͻ�cI.�uC�<�rdBd��J� �p�w�N�Z�8�
���)+�q���I�<��޴K�Y�b�2�ʗ�֭-*�]�N�&z�A�ɣ�b���^5�?�1B�?�[5�O��h���a�#�Z���C��'����`���>;���;��<Jr$Mk�0񓃪!a�(�I#&@�T��IҾ;�Q��@f܁~:z�cf�]+&M�h��&l�����:gw���{j��P&\���'?�0&]8b�L ���V�dQ��M3[`ִCfi5b�~
� t�����!Z���P�P�KD��X���q@B�0[[D�E�O�dm�%��b�������'$9q�b���:3�ل�I0uc�Qc�7>L�i�߬iM�4ˢ�	.0]�j��'<�Ѣ�$+�%[�}i��,� �	�_efE�1� 7�X��͋��.6�L�i4B�	�f�<�7A̭7���(�&�*D�V
��z�k��"�h-x��2)��-V.l;J<��- YЎ��)yY`��g��k�<�*@��h��˭G��(hVm^�[JAʲ��P���J��N a��m�)����Y^n8�G�:���Հ�2~(v��:���`Z�}.|P��M��ɖ��
S���6�C/f�d��i���h�AY�?Y�O�PäGD*��bJ*�8���I�t赮�;�4�FxR��R΀|(ц���V8�,�BD�
d � K,�,h �_�V� �����������apEM0�$ ��}P-ODz��N�(Ѯѡ6n��Xf�a  %$����m��i�2��32�ǧȕj��	����(P�`S�{�(H����+�D �֠�8�n,C�
B�	��x(s�I:�:�)Q��6z���
E�7�ԧ?&J�����N5��tFm�s��i��)O�&1����B�U�^x��_k��Y(��O��<�Rl�m��iH�Ƣ�B'�/����A��l�H,�az��R�o�%2��F�>�;~E����6��lr���K
�I�
2���!悹��C&`y�N���d�����.m���LQ>�ڸ�#m_���~��aeg:<O�Q8�%���EJFV'�����Z|����%Vbf�S��y"O�7 Ӡb�Ц3����Nɍ�y�QP'4����!J�h�w"��~��ǉY:y|���*��Ts,àe�P̑�)�O4�3#k��R���A�-@�1����l-�$4b�`YJ�<A���7��UQ�bۯ1�v��Lm�<كe4m�@�S�$u�j�Ԣc�<A�>LL�5G�;F��F�B�<a��G�j.�<�ĕ9�M[���|�<�S@7f���Q@j��%r����f�x�<�R#��a�����*D7V8�
|�<	W��g2,���ϜB��I*vD��<�7�5]��u:s-]�����^S�<��dG9$3v�8t*U��b�̊T�<�ʝ^���Z��%��T
��^�<�$J+SV��kQ�I�lJt,� �X�<2DT�#s�ȣA�̘MZ�1"��DU�<9���\�F�H�g���j�<9'���F'FT�S]?���&�e�<��<oV����9'(�#!$�o�<!��K=*'�%�
�-!d&�#�)�e�<A�`'�@`p���V�vE�0ADg�<��gX�V/��@#n� ��,�1��]�<��j�EV�@���zkR�S�_`�<�SE5tu�|�U\> ݸ��@_�<y2�ݒO�|�{�>S��M ΀C�<A�y���M8z�v��p�WA�<����S�j	�"&�;B��pHF�SB�<y7A��WĠS�ؿ9?r�cAV�<A�ވ�/ -R ��SS�<�׍To�X��
>ɬ zѧBN�<�w
�&T��՘t�ą+ά�_O�<AӭL&1��bL�AT�x0�b[W�<1f�H��Ub�f�� �� � 6!�DC2F�|�y�Ɛ:�`���D!�$��x}*쒳�_)[��	�/��!򤊈Y��1�'1�b��2o��0����P�i�M�� �H��Mq����yrH�;�N���^�C]x`R� +�y匄�LZ.нJ��A��<�yr�O�? ���ɠ7��"��y2�M~J�R�"�!�v���(�&�y���=)'���#`�5n��1���΄�y*� XG:I�ɖ�7�; �"�y�K{"�Y�(-zfy��l&�y��o�:I�jA�u1R �?�yB��g�=B��5K��k�k���y
� ��ـ(ƹ[�4�����b�"O<�5<d4���ޖ}��86"Oz�7��('��B�	����"O��rU�+N�:@�O�3��2`"O�4�W���藏���T���"Ov���	c5�d��m�.}�N��&"Ovx1��\�s�BizU��>@��k�"O�a:�����G��Z���"OT��#�ՠ)�J��§E

���9�"Of��@m�y_��1'��=��
�"Ob�xR
�1MҌˇ�@�9!l�s"O����ᜐKDF�S҃�f޵��"O4�r����<��-B���(��1K�"O6u�Ӣ[��Y@` @|���"O��R��|r�r����t��"Olx)��X��y�1ទ9�p@�""O$�[��?��4�ց�?m[��%"Oy�v��6���q��,.G�}�"Ot�7oR������5O<�! 0"O�qh2Ώ�=F���Q#��u(R"O�İS�'j� �	�w�"OpH���bT��P��4�^9��"O�mj��A�(�LS(H3@�hA�2"O�������:�gO;6���q�"O�L��ׄpa�a�E�P�[�Z��"Oh�⁀2D��7dˬ��d�"OX=���.f�~$���E$i)PQ�"Ot�# DPd��sR���1)"t#"O�\�$]�*��B�K��zl�
"O
�fGA(t^��QZ�ys"O��Z!�	S�����'YB<1x""Op���D\�w� ��FaM_����"Oa�d��:ZMxY��Aڔ�^�s�"O�����4& ��@S�4��Q"O� ���P t��S!̚��r`�T"O4�`f�Jj���KE?�>�B$"O򸣰M��;�T�i���/Z�AA"O@�C��I�Bh����*x��"O�h��
S�,�q{��сp[R"OޅQ��H74n���ȜA�QT"O��ŭҔ~���G�t���"O�!�ɹ'���g�c�hhI�"O�HH#0Ω#EH�Ut!1"O԰ǧS{6��@VD%	\,Rp"O�a��"�d��%P�� ���	�{ ;��S&$D��FÁ{��P�#ZWNC�I19�<d:r��M�b�R�5h���	�"�6���lh�)�'|:��<G>��2�]���Y��"O�� $>��X�I	r���X�U�tK��ѧ&o��C�'���J��M�ִ�DH8Hܠ=	�IجBэ_�+t�Ha�/̾�/�L͖�h�7$����x�9X&R9a�'ړ��m���ź`=c?]A1ʍ�D�Q1O����`/8D��X��� =��B��9`B �h��O�q�**Δ�N�"~�CmԬ���F�ja�iGJګ�y� � ��c4��gL��96�,��đ�a��I���<Ƀb�� LA2"&��A�f���nx�躇���9"� �hO)G���9f(BV�>���Ę�8�!���"+}�];�Y�W �)�.T�ў<���gЂ�QF�	�>\(��m���{���8N.!�DT�B�r�JE�Hd�K3	.6���V�J,�d�.�4�B0�d�84���r�a�O|	��ơV�Э��KM�f*2���'2��P!_�?�d�R��(X+�2H��,����"[!8��p�����Tl���E3^���k�"���ujN��y
� ���^�G4i��a�*��4���;��i���?�"�Ϣ����'�HM�g,@�y�I�py��b�'�y�GF��PVpˡ��1H���K7��{n �J��* �d�'"2�����f��dc�ka��bK<�7�F�*���'X<D�1���$P����L	��`B��ǚlV1*����d�2��*D��{u��4�2�ۥ��h�nE��GK;����+�L����q�֖���4U��]��5��³��;�j,�PgN
n�����O����E�*)��"��B�_��Tqt�݉r�r������$ 0��FrԵH7�F�*��**��'M \"�egK"W��Z�b	0Ck5O�|�a,�&,ހ�
-O*8B�&,T���!I/Pg*x��%��0(p�9B����25�"\O4�k�@�K��5��,D?���c��lC0OX�:r����Z�X��m��g&��I���*K��1i���t<$�`��&Y���3���>�y2HX�9�#��"�~y�$`_;����'D2��@i�x��`q��IW�H���w���b��`�Ai2-�O6`Q�'���2E(ɚ�PS�IV1��I�3	�(���9��5�D�"P9S [+b�<���TǞT|P!Ȧ	P�(���"o<��{`X�%`$Dר(2P"�~�#f�21|�6+�w$½D��t�<��F��5�f	��E�+��4s��[}"�9_(�@	�fY
t���[��S�4KB@���I$m"�=��e�+xd�B�	�M'~�СB�
�%�E!V��8����
�!ڣ[v���a*����O���`,�.瞵����fa�a�4��a�j��+�Tp��*Զ3f�EHD��hۂĖK��|b"S�Md��0��]�>��P��킃��O�y�.Fs�d�	Ӟm���8��<z3dX-j�P���P�i�C�|-`@��jP����:#j�+��W��m��V�Ry�l	P%F�����<�� b����@P�C��Xt"O����l�;�(��)� *�r�!+�Z���;��PY�"t���'���{&��#vB���t�@ }�P���J��I��C�-ج�)c�	/|����TN�0,��-a6���
�Scz� $L?b �i@��pDR�2��-^%92��O�6���E�^?(]�� �,h��'�Dh�Fʗ�<���A�H���ȉ�O��'�@&|�36��8
z����V��	 C��O�89��{�h<0w��^��a �!���G���aIU�#���Í�n��D�ȓ�j}@�g�1-gZ�K�A܍y,��0i�WI�a�4������i""Ot�x�͎dP��U�(v�����"O�Y��˄,� XUF�X�$��"O�Y�UD�>G��)����(�L�"O^	�J.s��f�0��Ј!"O&�jGoĭ_��yU� O�a�%"OJ�b�&���,�!2iZapB�µ"O�,+$4G��}[�)�gjx�0�"O�  ����-��*�b�R4֕#T"O�-�"�[�_���%�\Txq�"O�}�v�C�o�y�unՈP���"O���Dc�gΉ"4l�N�Vj��D�'i)�Q�'�FເA.Y��f��I�d������*�.G$��)D�M�C-�0�`
!]���z,O�В��ڍ��!mA�0!"nԅW�]Cs"ӿ��zb��`�ڌ���O�̻0ǈ�R�$���<�\�	Q�Y<	u���Ͱ>q���!��)��D��a�x`�E@�a�`X�CŁu}L�	YI�!H&ad<�ӳv���-؊C��K�B7�C�I7sĲ�y�ȍR.Q"���v�\c�,ژ�R�AR !�	6��OL�Qz�w�b�)�� %�DB7lF�P�S�'�����t��d9� 
��峣���'���b3��@�<=���I1�q�l�'��I�No��Z���q(�I�a� A��ā�ݖ���K��ybmǒ�8�&���(��0"�m��AXx4���dd�I#C�L�2��S�'ߚ�!v���s��|30��.t
�q�yo/q�(!�I�<)*�5���r�`k�y{�G��:��e���Z>E(�Y8c��7X���j�	�~�e2%䄱%�V�V�Ь���ϟ P�	s0���<a��M+;���a�E|ݝ�s�_OJ�c�*�<y���X����3�P
�* 5U��B�I�u���T��,�y��!,�P�`�hA>J����A��a*�ү�t���I�-�鐖�~
� ���q(hU
��VC!.~�i��'e�Ÿ(�l����b��=�O̠lMd��wiY����v(]�x���I�x��uR1�?b�Q��2��4e����Q�����O�!S箐��? ��6F��	T/�O���!����T�1 �q�����k�l�H�A�4�p?ycoÕ
D���	cJ�"��
t?� BTu��T0sB4?� ��+�p��X��Ia�!�5摘�����>%���߫&D��A,�:IV�1c�P�z�XP�n�#}+����z�Rh���)��I�
QT��b(�R���F�-yX�7

uS� �c�<�b�Y�- �eT�|�eϋ�a��H���C���sr��Q�r\ip��f��O�혂@B/wϨ#?���	*B����	4�����C��5I1��+k~<�GƲ�y�AX6����}�i�9qaH�>���3s�Ӥn�<P����(�0E��'�(`�fP?+�<Q�BH�i��8���.wC
���n -*�̲=�j�Z�D�98��i�1��L��pO��O�s��9�F]rb>^snD���I�j{J�IGL�';t��_v`l�
O�duڽQ�6Xk��6-޷)�)���<Af�[�~Ӿ(s�L.Or���˒I�lԈ�-�� ���ee�?B��4J�K�v�I,)?�%
GeH�U4�S���̀�h$�b�BĄ"��K�IW��X"Q
O�:�/�:"I\`��N�/������i��CG�H�hQ��ЄE^ߟ �%`�tD���VE�My�wQ�9��j�+Dxx
&-h�X���hl�h[��.��x�1��^8ּ�k��g�֘��Z<�y�#��L�L@-�y����p����2��:�N̚��*T��i�д9lX�Gx�
r~��ȕ-�V��7.��9fb��՚�(Dr[���g�F�]RO�`y����<au(��M�
Š�픉&��̹��N�V��P�DM��	�D�`*O?�	�Gو�K4�Y�!! ��I�I�>C䉬]P�qw�w�D��b�7"���ɻ��u�Z�azR(MRH0�3V�'{�i*��>6nR6UZ��CJ۩Tt�1�Q�J�.����)�!�$
�m��u��� ^	� �vx!�D�6pi��.ʃHT�O�0!򄁖x;,��"h�!ot���D�S!��
)�$��7_V]����%!��@�Sz�Q��3�\}8!/�i�!�Ěpʮ�sAo�&@��<Y�$	�!�$ϪIpҀQMD�e��l�HH�!򄂁9,UqF�Q�/b�#�U%l�!��ʣk��=X�NTd�;���+!��Ђf#�B���H\$Ⱥ�ꜙ[!��_"8��W��b^�� �%]+!�$@�o~`؇fK�UJ�Sd��6(!��K! �@	����qn��5�Cu!��&3Z�q�!KQ|�ԣ əu!�/l���e��ND��bG��!�T�5�@�$��#�YQP�Zqv!�FվH؇L�`
���T+x!�$�. ��wh�(6�ڄ䜈rr!�$���hqrAM�B�V�b	��VG!�$�!{��ð	';��E��	8J!�$�q��5�w)A3� �פ��5I!�B,|���Y�wu��q@T5!�D�=7~\j��߭i�(
�f��Pyr�5	<q�PE� (��-�"����y�B�D��c%��'J�,@���y���1�T9������`���y��§x�:p৮�|��	q�K���yr�F���v
Ll:��-�y(�3�����B�[:$Ъ���ygܘf*���d�0gJ ��+;�y���v�$�e�&P�x#��+�yR#�2Q�������f�+%'*!�d�
Ue�X��E��λ:6��qd"O�1��R�$�|�J��B���>�eN@��4��B#;)�aRa�[l~FwR[��h� \�Q�?;���&�=EBU�Ox�30BM��0|b�D�.�L"b�<7�e���Lx�䞻xo,�"����O����Ozܐ#EH ��
�킎R�M��O �@�N�mvp�����}��`�P��%G	]�U�T�p��	�5 u-2p��QS�O�?� L� 3��2�6�����'  $�)����2"X�)CI3?�C�!�Хӡ�\6/f��C+@�l�$!����0�i"���Rd-�n�ba`��51���#"�>��&;kc�e�Wd�<��I�-w�l�y�Q'��3d���>���;/�8�8�dء#����'�.ھ�Ms�đ�
�f����Y4�T+�ʝI̓Y5�P#���I��~��M��=���\63����.���C9lgB=���?��'$Z|Ȃ�"1�0آB�mp���E��,�X%��?e�~r��/?m��1�g�H� |�́�G�h��Ö|���D>��kz�]��eݲ!��uP�-p��'B���������'fy�f���ahr}�F��}'A�O���V�J�k�1O����+�Hm�`&=tܨ���_��~RJ��O�>�!�Q;�Խkr�B0+p�	JQ��?C�Ex��4��$�F8��=�g
�m�P˵��4c�'�R��Μ���l���
C�FG����ρ�:�F���[?.��	�~"b� .��u�O�h#|
��<�n�i�C��u���Y%�P�t����+��j}��,O:]P��L�sV�x3�&�p1G��А�j�q���R��-��$iu��P�*[6�i�$��*�H�F ��b�"R�i��h�<p�6 P/��	��D�E�4-�>	��ORM
DG�(ð�ӌ���h�3�䀊j6��O��ˊ��,�;k��W�Րs-��JW��rw�a��b��8|�ƨN�<S�A�'9+UN8J�*�X @]6�ȩn��c�ȭWI
���W>����+����q��j�<%S.C�ɂ�9�	ˬ
�m)֦��&H&C䉿#E��y��6�%�V!$�0�y6"O2�i3jJG��2eL��q�N1i"O�X�� �8*1p���q���["O���D�0���
E�(nrp�k"O�e��mE���f��F_���f"O6(`�O��8���Q֪����-3"O�1��g����V [0CJ,�0"O ;��W�e�����
`�t���"Oԉ�PK\s�<St��h@i3P"On�B�gO��^�	�Ȗ#@��:r"O���*�0̱��f��M�>X��"O��)!%áBЎH����[�\Ӂ"O����܅x��ة�i��n��eِ"O�x�D�G�Kp8!�)O��J�"O6�����6*�����G�c�F@��"O���A�rO<��싸�:q;�"O��@���k��Б,���M��B�	h�N�p�dޚwI`)��Q�;��B�ɚe;�t��g�1!\��7.��|�vB�	2,.�а'G�mq*���r?C�[8zx�`�9����1��B�IEX�XA�l�ʈz��D���B�I�i2�L�F���
4�-��B�?�RxXQ-Ƕ}���RaOA�]��B�	�|������\ 4�*-y�޾h!���v�J�	�x0�"-ֻS!�d�4׬ŀ��\�݁�Z<Y�!�F�h~mZ�c�1�� �+S�!�ċ"�R���d�/U�%1Ǎ�5�!�$ �+V�MH`n�8�Z}KwA��!���^���̀(��tX#K-v�!�DA�Nd�d�[%n��
��C[�!��".l�z�^���I0�T �!�$�8W�dq�v놎erB#H�!�̫�t�x��� a����X	!�
�WD�P*ڜyKb��@M��*!���6$=���U�H�Dbɂe!���'�
���86q�b�#f!�V<Y^���Y-T�x�Q�_PH!��O��h�Gl��V��⓭� Z�!��ـ)f�00h�:V����+a�!�� �%Y��×(x^�1d��8Vվ��"O�Q���}Ѽ��ӈб6%|E��"O�MauO�tG����M�AQ�"O`�0"a��:������;���#"Of�C���L�P� �ћ%َ�3�"O.�{P�gH�,����ٌ�d"OH��d$�;N�,Ju�+>��ᢔ"O�P(��^	9��m�#���/��TU"O����A�!�v�h��V9P����"O�]+J�)c��;!��:l���rB"OAt#F7����C�"%��"O�rDX3}dؒ���1J��P�"O���M��:��`N����c"O(��Z�	��� N6�U�C"ON�R&�F��ab��P��qRu"O�yB@���Q��,R0@���g"OT#�\&>�D tlT=$��x"On@Bw��5\1��B�R��pR�"O�"RÊ�(��҂�YP�L��"OXMs!�L#	]ƀ�C�D-9<�H8"OꝊǇ���@��O� E?��I�"O������*.
����2"4 A"O&��G�~��1�_�OrN�h�"OH	���{���*5(���*�"O8�z'�1l��Bb�O�v�V"O�ٙ̄O��B	L�S=��y�"O�����	��X�gMN��1"O�ܨvEГ5^.Z��O�S��A�@"OP�(�S��	1���4�*t�"O��xă�U�< 2��I�:ap�"O�YJ��
����D�O�(��h:e"Ob�1!�d��P�r���+�.mCb"OƘ#�,�u�:Y;�#ʶp��"ORӖm�
L("��I9l�X!P"Or ���O<���� �+Dڑ�"O�{��
H���D���3^����"O>MCuo\8��A��I+v�|q�"O���d��&��+�oX/����@"O&����_zۂT@r��%k}Hb"OJ�Q�@�6ߤQe�E?w^mr�"Ob����)u���*C�@0|i�"OJ�HpK�}A��S� �
LI��"O�1ZT�A�C�4�P¨X�yD\! "O���`�(@с��r5���"Oމ���ӏl� �C ]1
~��"O�3��'}_�)�(\X�"O�{!˜�M����$' ���b"O,"��E�^�$��C�����"O��@t�  fLqx5L���z�"O�%��@-L��,���R�RI�&"O	�'ϙ�cV����8j�y"O��@�>iJm�'8x<-@�"O��𡣔�p_�iI$�J�,�%��"O�]����mf��zp��lӮe;0"O�(u%yd��Fڽ1d��"O��:� H�pev��E�vW��;2"O�mp��!��(3u.�KP�{�"O��ti_8T�ΰ�2�#"F�IX�"O`��6רFr"��w��jh�@"O�eBe�	�F�y8k��ner!U"O8�c���)%�� 	�i�$iY&�j1"O��u��i@8����l�Pu�p"O�me��#ݸ�ܟ"Ӟ1{�'�u�cn(AJ�R%���M@ X
��� z���/��p�<�u/ȿ`����"O��l���F�:F��	&4-�r"O1B7���b3b�#�;���"O�����"R� � /T�I�"Oƽ;�m��g����שˁ_G2�H�"O��QƮ�XC��Ub��{ǔԨ�"Of�����J9�}9`��fqS"O��4�˧]�1D���S�T��"O�ē����@�z̰����
Q��"O�XsΜ�V���(�KN��v��"O�e��[Jv����q���r"O�[%�C�:4ޑ� [d<��"O�A�'@C=�uX� ZQ4L�"O�y���E�5�F$ifH�8>z�
�"O
hQ���?
.�0C2��lKʜ
p"O�	 @F�2.^�ݰ�N��O2.Qٖ"O���DĬ|Ք��e�B���,�S"OP�d ô\�d,;ߛt�Ё�"O���1c�Uc\{�(���V���"Oj�3�p��� �NX�!��%b"O�|ȶ�J1!~����F@*fі�[�"OX�i@A���<yE��(��X�"O�� Gm_���\ks��!�, �"O*���KT/nΌP����*\#N<)g"Ov[��S�2��b�ʹg
z<��"O��3u��g���A�u��!��"O��R��q�nͱP"G�kd�At"OV!8�)�6 <��\n��!�!"O2A�0�J7A��dab	ɷe����"O�pе��>Q���6G��Jb�ī"O���/ìB��1m�W���+�"OH(��H� (���b�ǳ�RI��"O8{v�Z��\XYf�t<�8�!"O� ��Th��[b�]*- ���"O�5yR�M2'���*f"Oy{%�ˈ]���uT�P(�"ObH����1j �"�ޗ :���c"O�A;2G��2�Y -U(!|���"O�@,T5M�B)��%�zbDJ�"Ol}�@=Y��a� Aifؚ�"Oes`'ҧ-�̩�*֑Z~!8R"O����g0lx�D�Ț,=� `"Or�h����F�l����֟��|3g"Oz�P� �R(�A��<\��$"O�%Zv�U�~�򕎟*TYڱ�"O�qX�`!m� EK��ZL��RB"O�Q�p�-�p��h��*>t)*�"OJm �RYV�	!'� �l.�5�"O�]�R��s��"vKM7֘)�"Oj �4%_�=ۊ���)<p�b"O:�sT�D$}�zԠ�"[��[a"Oz�24�iḓ9����E���"OT]�s K�����o��L��0�"O�`��ćCn��N
8���"W"O2qk2	O�=.ؖN����a��"O��WD\�qv9N�&,y���5"ON!hC��sr�Vm�w�XU{c"O$����'e����	a|M�"O�xX���5�>D@ !ϟkr�9�"O��P��/{��� ��BU�A"O����dInҼ��A��+�,;w"OXIe�@�lI���P/�|�M��"OD����C���.]�bi�I�"O�LxÁ
(��݀��~\^4�"O� ��{�@ o'�DZ@��(mL�E��"O�ٗL1N����H+ L�k"O��Ն�
e~��ș#8 4j7"OT�J�+H��Np��L'DU�F"O�X�S%�	]t����.U�=�z�@"O � ��0'���$�'i��|�"O��b�X&��(�2A�>sb�Y�"O�(u��n�8Ȓ�/�;&�֙��"Oؘ�1R cHv��e��� �"Ob0Hu �\���d
Ia��`�"OН�g�@$!94D釈X.v/�!�R"O�=s�l�$V������+����"O�<�$ ���j�ÝE���Ab"O~٠�M$n�(a��]�u�D"O�]t�����L�����J^3jX!�P�a3���)�0w�(mqC�_�+�!�͐6�Ȁ���
3�,@rB�2t.!�$$���%DM�|ʨ=�!�дq!�D=�(�ӧ3ʠ̈�
Ƨ"!�dɟ	�&�@sHKQhq�	U�i�!�d�1`^�2�^�Y~Y;&H��/�!�tpVb����x�FL\�,�!�������F�!w��|��̕0]�!�O�x����AV�m�`�
%���X�!�V�m�~k�MJ�ck(1�����~:1O$��Z$Pxݛ�4�H��5���0x��!E����>A��y{�H8�O4�N�9�`�fTf8�$�ϝO����-9Di�Mˆ!)�
Z*)n�e�>Tl�^y��� ��\��8 c�T�Q�z �V����A:
x�$b��<)k5�$�*O���f���$>��O��ѩ�[�v��zǌ�87>��C�h4�����r�'��A���?AFҘp�f����K1�f�oӲ�(�����׌;�`x�&����p��%JRl7M�OT��|j�'��'�b��3�ɚ{.x����[��ݫ�	�5,�\�4A2�I��.ն9��E�И?��0Z�N	I�$"u�Q
>4(V+�HpF@!aF�a�L����R�
l��G	%D�>q��wZ�p�Vo	96 �)F"6p5��E�OR�o����Y-h>��w)�u�Ō� }��I��^�$u��B�O���G~2�*9D!�I& Bf%[���:��'L�7����}'�����?�o�!{
`��Ë,88���حF,��	'08 ٴ��<�ߴ}B�D�������1P� xz�ƀ�zZ]Q�m��3I�Ĳ��Ͽ} Ґ�����'k��H��7�>E��c��6&�X���cн��M_9�	CpD���uWN�x��?r˔M0����a*Hd���Ц�"���O���J�I֟���~�ɩ-����&^�Vr04d�^1^�Io��h������*\�Ȋ�"�Q�$.����4��L����O8�I(	��x��4�Ms7�ܐ�U,�1�P�s�a�$���OĄ��͆>}t����2d�nł�֪!������&��`�OڷxU�kQN�=Q�LPZ���pT�ַLI�m��)�_�!pp��K ����M;m^/b�<Q0fҟP��4(���B��Ҷ4`�EkШ�"7?NI�q�-�?�+OJ��%/�i���Ok�(��-B�j&���BE�f�p��'�X(�#�Y�hP"�ϑ�W֘a��i����4��d�+���n�ퟐ$?M��ay�I���4��U��[}�T�O��$�j�2�w*���K�!��S�����6����_9�ԛ4�\�+����f� ?#c����.BW5�ex�I^�H����e��W�0H7��ϊ�B"�#"R�Y���U�'�HM���DVj��d�Ʃ&>��O�ʜ	gI\�H@� �㛺9
pѳ
)��Ο"|B�Or�[���ΠW�ݙ|)��k��'�7-����'�R���M�-Č���R�V��q ,G�X� �n�󟴖����OǱO�,��'�= ������	�)Ahŉ+]�1�P��J~�hi�������"�<��'9c��]8�Y0em��i��R��_5��� ��_`��)���2���0p��ͺ�%��μ�D�!Gx	@d���4��0��bO��Nu���z�O`�����Ow��}E��喰E�����.Dg��D+LOX�'�~u:����8�H�̡7ۢ���{�	sӼmm�I�?A������I�|�,������}�|���A3}B�'wܝ@ ���   H  $  �  N   �+  �7  �C  M  `V  e`  :j  t  Z}  I�  �  �  y�  �  ��  ٷ  �  \�  ��  ��  '�  k�  ��  ��  1�  s�  ��  � �	 �   * �0 �8 *B �I �P �V ] ,^  Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�� |d��"O
`�(�;���8���-0��1%"Oj4��ND^[��"3/9�0|H�"OB���H��*�ʞRy=a"O�味V�!X��!&F�:J�$���"O,��a
���C�Ą�M�"O,$3%o�-���p���+Ն�:1"O��ݢ1����`���y14]2��i�<�6��{_���c�H�`�fX�$Kn�<��A̼VI�xR[�)�Ć�pඤ�ȓA5��('nߡ4�� �)˩%� ���,��r�؊b#`T�eT09���ȓ!�b��g��}�8�F��-? �ȓ
K|m�ș�VṔ���2�%�ȓ"R�X�j�4JN�1�˘X�i����̹	_�jZ��1!g��zܶ��ȓgil,*�J�
j�Ne��i�J%b���f	�(U��:���G��$Y^م�~r�� S�%T"���k\�jx�ȓ|4�1�îJb��@ӵ�ݩn�V��/[`�"�v4�R�!ʎ<��M�ȓ`:��z�ؚh�J�Z��$HY:	��H��p�m�C1��!��B:��0��EnjZA V;9����J[
2���	��4'J�EA�IVW&��~�(aZ��ӹ�>� o�Y�|�ȓ�f�A�
Ο7�H��M�$�����mޠP����/���ANXo*�ȓTv�����{ ��-7�*hE}R��
I�91�A?b	�FW�Q�XB�ɸP3�)x`d�?�,a����~�S�pʴ� 5���r4�!8Du�j<D�01�gKazeȠ���I"j�(r#<�����[�Эp��r�n#l(Kd�'p�NS�iR�� ̺��D���C�ɝQL��F�E�D7Z-Q��IWuH#>����|�,}Q�H΀3����
�'F�ȁ��'������Ί_�p�
��iB�!�ȓz�@����,���&�A�m�+ D� ZU�Q�
ɾxQA�$1N`\Y2#6��0|Bp���9���� �4 V0�E�f�<�AQ�r��R���
k=�Uo�{�<1���!St�:�υ�~؈��!Cv�'`L�E���_�/�4a�1\�C-Rس�>��>��OT,낭@�?`���֦�e���C"OvI��j� ��Aٗƌv�Ҩ��"O�8���K��8Viگ�<���|"�'iڰ#�T�e������I54�q��T����I�y!A��9v��§i��yl�G����4$Fe�bܓ����O��(�J�O� �h�M_�WJ�t�R�}G�t	�'������c�*��SGɒ �����O���X2�y��l��
'���,�a�1��հ>�w���(�B�+C����@ k7�풡�%��ȟZ���i��P�a�' X�S�"O��#A�ǌ+>�9G၃o(�8r�+4��M�)5 �rF��SB���:�,�S�{�����Y)2ZXt9�b\�gdńȓ\�8��aB �n[�@QԀםd6�Gx��'��s��\�m6��T���/9Jx��'��<GԳu v��ԍSW�"���d5\O�YjW
�3Z��dHR8J����'h0�
� j�1�mQb�,\2�&m��%"O���� Y�S+t�� &W`XB@�'n���f�S�O+�E;A#_pP�ـc�>5UJ�p�"O����ȁ_�]�sb�+5Q�H��'O(�i��2pn�_��в`���퉦I6ʬ��OX��ٿB=�I�Iie���"O�,�q�^�wiX ��H�<s�b9�""OR���H�,r�Vx���d܄�1"O�j��҈|q ��J��$��]3�"O����Qb��oͨ?R ;��ZD�<�F@ȝ)c��9�C�Y�ڱJ�F�{�<���9&88��4�N=���y�<��Cu���
䏚�t��AzF'�wy�O���������j�/�`�IS���ze��"O4�TF.e�*@@���4���1OR�bJ<9A�#�gyO53�=h2G����E����M����s�FE�ҙ`,���􉂳3$���o�,�PxK��
D�$�q/F��ܣ���5�y�b�5��1hĕ79m:o��yLV�
������4�H !��$��'�ў��Ђ�
M�#��I�➑�� "O8D#R@�N�xp�֯ � ���}����B��|���(�/L&c���y�X/=*���t���K�$);�]�ȓ3@��2�U�?�H0�3C 9�`��X<U,Q2D��6�I?S<|�'`N�<� �ߔ/ڒ���a��c�
q�b��ɟ@�����D58y)�oZ��q�D�T���	���M�(S�Au*��n� Ў�aaIr�<����	�r噦�ϓAl�9Џm�<��fƩ*p ���V�L}R�x2�+��x�(2Q�@��Јo���8��O)�y� �)ST60Æ
	b�n���FX���=�y�pZAӁ�н#<Dʦ`���M[u�)���UF�|�2� �sa�	��G�<لg<}�=O�}���]�p�<xtdZ�#�Fm���~~��8�O�i
I�!X�P�jvGȽ�~�J�"O��b�ՔO|����ƉC Rq��'�@	^�d�=���)pĕS�'D��[&F�	0�6u���Vp��`����	%pf>�
g��[bp�:�@�l��"<y���?�)�&Q'��}"@��<4��l+D���a�5+OJ�Re@�7c����fI�\�'=�>�	��ѣ`'/�n};Bj�z�D%�S�O�^�@�`	�<bIp��w���"O
�A�AˊkҀ���LQ�v�[P����'Aўʧz�0@�%��V���A���k����ILy�g�S�p�ak���8r�1O���l:��<���K�N;^9�nƭL�����i�Z�<��DE�/LԩBǌP[��1t�b�<Ï�E��D����4Cwܹ�vD�Uy"S� '��g���K�����Ej��!s�,�l��{¹i��\��d�̆�A@<=���]��.��	N�;��i���L�R�jl�`��#J������~�'9����:hDZQ(.B�`�''X0��X�0K��`�H�6g����'�l1��^�Pߦ%z7DM�5��s�'M���E�E�nJ�њ�#�)��$S�'zX`#��N�&A���<V$pq�'s�q�3��gF\d��`�:Q%�<Y�'�A����0G~���&N�N�n�I�'`"I����/?��
�� N�X�'M��e�aoA�CңEq�6"O��6HUy�0����o"�s��Oި��ާ� &�;T׊,�h8".ϓhb�C�'�� ��!b��,\�}+�ØY0B�I?A���2��9$�~��t㊌QvQ��`g4�D3擯N� R��Ȕ�J�`0"�t2�C��9!�<��%U�D#U�!c�C�I�+�<��@&{{~�u�B�ZfC�.DA�*�k�A��U�1��4A
b#=a�\�^�jc�����r�$O`|8��z�	�_v� ֣+�D�k'��g7�B��,�M��H#�`y���S���0�FQ�<yGi�)��)�����Q��X��043O
b��a��# ��B,�����4�9�HO�O��)�`k��]��Q3��c�2�{�'B�iS�>�8BȎ�j�|QK�Q��d"��Z�'����d�Gc ��Qg@���.U}��'��O("|:7h��LbB�x��7B���b�gD�s%���#�����(w��Pv���w��O��=����!=U�P�7.T�Y���0�%TK���'%�E����9��'T���>I�b���#���%1;xU2���[���ȓY�xQ�D�}�T�s����"�����85������
��dk&�gY��c�i�"~���s��%i�aCu
fup��X�(�x���9g#�Vh���@� }Z8��/�U�ay�e,5��8�w�аDFP����O�"~Ҷ�Ζ!;2� ���78u@�jQ�<q��� J�lLc�$Ðk>�Y�V�]ey�	L�'p��I!��3��+���"}�"O^L��$�jV�i��qx��������֜��gy�'lQN���L�d�<҄�/c��M�&�'0�El�;!���s�Ǚ�_��� B����'W��I�'�1O�St�|)�bo��̄�I�
na�B�	��Ac 8��\K�+ʞ>���J(�G��t�eD�&��� �m�n��`�g%<OJc�����SL@��w#W��
���'��x) B��#�D0@�jМ����R@!P� �O��ю���$�S��r�笋:_NKcT��y2F�t��5I`�S�^��E�$Dޢ�y�ΐ?Ѽ![AeS�B����yR��j,�˷�h���r#c��yBBP ��+ ��&HD�"���yB�7h�D
&ą�BN 5j�����y�g���逼e��`��AD	f���	�'4�ɶ��	����(4%�
�'�l��cd�-���sa��(�x�	�'��yZC�1Tnh)Zk�/Fi���'�&-��� j���Z�mN()bꍘ�'�&�R��-��� O�� W6�	�'��8��)%*zŘ7	����	�'-�ͺ�Ҷ"�J�����+d�		�'�f�ȷ*bl ���|����'N�i�Q$|eT���-
F�
dc�'�~���韚R����c[p�Q�'#�AB�D�<,p����rR&U�
�'��,��F�6���m�l�.�*
�'\`�cT��TH��2`ZT
�'?d[��G�l�I��N�@o(P
�':�a0�Í�fR�f�2��
���W6D>����!�dt`���yr��.q2�"�n��r�(5i͸�y�`]{�M�o ,9*�
UC���yr��GznP�6&E���l��._��yr�H�A�*�'dʅh�8!��_(�y�l�(,H ��vٖH�.��y
� 8M�'�V�|��uY�N�1V��C0"O��JB*=��̸w^�"��"O��IEǍ~"20s��@� �"O��zD��n�s��O�hlP�"OTA&��&&<H�Hb�P�D��pb��'���'H"�'.b�'J"�'���'���qJ^�k^ 	Nc��=0P�'���',�'~b�'���'���'�	��G	�<c�ѡ�!%N�����'���'Jb�'R�'+��'���'���@VC�1V�,����>�r�B7�'W��'��'��'���'���''x���HI�&E;�̓�""ةV�'��'���'�b�'�r�'2"�'��z��Q��J��*{����O����OX�D�O��d�O��$�O��$�O.\�F�K�2μ��G!m�h�c��O����Ot���OX���OJ���O����O�0r&$�@��Q"d䍣^�R�Y�,�O��D�Ox�D�O���O����O����Ob�:1HP-��!���L�}�$ҧ��O����O����O����O��$�O��D�O0Q�MD�S��QB���KO֜y!m�O����O`���O<���O��D�O���O��R�F�!��1�L�Tx�z���O����O��$�O���Ox�D�Ol���O��%�]�,J��D�=
�F!��F�O���Or���O����Of���OR��O���qnM@<����ȅ9�p�����O(�d�Oz���O�$�O@�$�Ŧ��IџX;c�

i5x ���OR���	��$��d�OJ�S�g~b{��p�f�6e��)�E��`H���h�	.�M+���yrod�L�������\��cg"<�"�Lۦ�ɾL��Dm�]~�
^!S(>H����e��;ȸA*6�߿#>�Ҡkٰ�1O��D�<��i&t�va ����|�T�+'�ѹ��n�"nXc�������ygF�B���p�Ά,X�(�>F�6-O�������� -��7�s�`8�h�Zr)��MO�s6��aS!c�Рeʖ_��w��_�����'k� �e�0I��[�f	�y�yA�'��	[��M���{̓W�V�G	�>.��3�Nd�f r�RG�>�Q�i�^6mn���'F~q���O-"�㷮��R`��O �2��vx�HV�	�skt�]��?qGe�:_���2 'Y������K����<��S��yү�J2�s֏\>1&�{���0�y"`nӚ�;��� qݴ����4��`��P��hU��a�yR!f�*ynПX�#��̦Q�'j��� �<�+`/��j�DQ���rΰ�ve_5��'��)�3�ɒ9x��!��_'�̈hƕ?�B�&p�&��7UB��'xR�i�HRe�(�C��1�B)@n@���'1�6�CҦ	�I<�'����2x$��N�$PuZ���<�$ZVz�L�(O��[�IK�UX-z���n��I��� C�b�Ťҥ	�L��a,�nB֝	ԎB�%nu�EK!	�ڱKf�ޞN� 4��g]�j���3�)�Z*=HW�M����L;=�������l���!��C&��i��3M#Ԙ �,�z����CX�OD��tb�g�ؙ��f�@&��Y�%�6F3b��I؋nT�i��(����6�C6���H��F�8$"i!rԡ]w҄�0OՑZo�T(����hMz��N��Y��EO+<�3����Kaށ��e��I�YtC@;Mm2���@�D*d!��cN�~O�\
�!$O���iHz�ڃ"ÄRr�%	��<Va��#�$�O��O�� ����'/<%�fN|�����B�cǒ�{�O��D�O��D�<A�kC�O݉OJ��I�M�h�.Q�dkZ(_b=z��`Ӻ�D4�$�<�6�o�/�����=Y+|-��*GhP�o���oy���W��Z��៾�#�N��O�Z\�֩1i�R��!	�u�	iy�����O��, XD�F�O���Jƒ�G:�6͡<��D��_��F�~����c�� ��c�;��xR �˭tД�p�rʓY��Fx��tKِL�X;uΏ�{�P�����/�M��mڨ��f�')��'��t�4���O�d��^k&t��S�X�S��<��Fܦ#e'�S�O*B�
�}k|�S�I8���0*	7-�O(���O��Xa��?9�'��i!��;|�DU�9;���}�N�Ә'�r�'��E<Go����^�y�Xēa�ѹoc�7��O�E���K�۟ ��ݟ\��5��B �#KT�#5��x#�����Z�F�1O��$�O��D�<a#EU���a������:���I�r�S�xR�'"�|BP�tQVN]5kT�#IMFڡ0$�<�c� �����xyB���Hx��y�v��4�D�rh:��B73����?������dR�aK�I ,�p���_��8ʢ� �h V듷?!���?	)O�l�+�S�S5�lqSf=JҌ�6��R�(	�4�?AK>*O2����D�*ci��Pcf�!�|r��$F��6�':2T��������'�?q�'si6�1ǌ�/?�% Sk��5�z9� �xV�(��$�S�t��0v��@4J�TW"my�H��M.ORT:�㦝���N�����<�'�{3g�<%���LP$E����4��d�c��b?�i`aU-d��<I3�_?�h���}��)u��O$�d�O�����|��?q���h�Fڋ;���s`��%O ��i��%���'wɧ�����s=0�u)�ɾ���P�;��pl�������� r��Qy��'���'g�[m��jӂ��4L����׵_�OD<�=����?A��m� 4W�I��)�JC"#��|�s�i����0��	ܟ���ן�&�֘2Y#]X���2L0y�5�ҙ��e��HJ>����?Q���䝚Z ���@�1.�
�쉻	�T,(�`�<���?Y�����?Q��9 �d���Ǝ���
1�=����RM�0�?9*O��$�O��Ĩ<� ݏ���唔TD�pcd�t� G �M���?����䓐?���{t��h�'U��£�6,�n12��M4���p�O����O���<�@����i�Ol���H`zT@�W+.q&��u�	A�Iǟp�	||���=�H�(2��q�"fr�H����a�imZGy��B��SƟ��	�?�u�ƌ6s~D��(���TSv����ē�?��#?�����S��BI��*�bK%Ş8����;�Mc,Oҙ���O���O��������C����S&�>�`u:�cW��	����P��m�S�f�ġ0g�.]_�ԁPj�
{��nڿN����֟�������SUy"�'"#�(b��8[S�Sz˰�p7d@�4�7�mA �"|2��w{���6���4){��:�u�u�i���'���@0I���˟��	��� Q��JJ�xa���DkLl�>�A)����?y���?�De�<q�q���q6�,�A�C>Y���'l�aA��&�4�Z��Of�<q�-�aL�Dj�<�6(Y/L�X�(Ǿi=����Ԗ'>��'�B[��j1��<`�:di6)�7~�H��3s�mN<���?����$�O���$xCag]Hj���s㋆XT7��O��O���O��U$��:�ީ�aOǭf�^y�e�4w���Bu[�8��۟��Ijy��'o��H�A�o�93�Ө"lx	�4d�����O�D�O�ʓ)}�MZb��T��>��8@�j��I�A:'&��7\7��OP���<����I�O��O)��r(�Z��"21�]�ܴ�?����$���P%>1�I�?�ؠ@�Y��j��#{�@�04a�6�<���?���?)L~��k���� �FG�o�p�ia��æ��'��\k�l�8�Of�O��Y�pԅM�m���s��K���oZџ���ݟd������<�+��f�]92�8�ۖ�\�v�B��"�Γ�M����/؛v�'���'��dk;�4�̑٥B��kB��j�)��M�����g�����	ӟ0�I�h�'b�s�d��6��mI
�G�84���J$��xߴ�?1���?��5a쉧���'�"'�R4�@#�Z	~��yQ�V1�7-�O\��<��]?�?���[�h�EJ�5X���I�}�<��i�"b���Śx�Oc��'��I.R�p� �������b�F* EJݴ���O��?��?,O@mU�\tWL8�]QSƐ�󊝣T�$���I�<�ICyb�'��$�j��z��U��Q�n����џ�'���'h��ğ̰v NkZ��#�~�ӂ�92���r���ڦ)���t�?���?�dL�d��nZ7�X9��I� ��լ��O
���<��bI04@*����Ò1X^-Q����DC(�%/�čm�{���?y�=�N����^�I+Ss���"�"E
�U�� ��h��6��O�d�<�#�T�Mg�OR��5B�.�
L���/P��R�� �M�+OJ�$�O`��P@�Op�����=@�ň ^��DƪGI�xa�U���F:H��	����Iş���nyZw�X�����:i�Q���ߴ�?���x����7O�N�S�]�n�����`2Y��?v�oZ
{y.$�۴�?����?���P���D�0 rpHZ'�u���
	ٖ[�7��(�����O"���O��i�|�'7p��.�q��/�}u���lz�$�d�O��$��uUN@'�������G��m ���X%"a��#s"�s�4�?I��?�'�4w.�SB���'���ϸ\&��B�B[M�2�V�p���'��I�q[�컨����2��C�%	�W.Oz�b���DǔP,�%�D�O���?��D�,m��1A�L5 f��m����.O���O4�0���䊒���.���� ڄz�*`��Z~�'�B�'��	�Yux�O�T�"b�(�+@d	�+��ڮO��$�O|���<a��?�&.���?DD�,3H�]��ƣ*Ǵy+�!V9���� ��ǟ̕'],� ԋ8�I|��������-�b�����@�n���<�	ly�'"ҢM���~z�F.8�,��t'�4w��Xy�����	����'��M7��O����$��q���bb��JE�с��i���ПP�	�.�Ƹ��s��?��@�R8y�OK��($:����j��?�-��?���?����(O�L��"
ʷ ib��rY��lZ͟�	X6�){��4�)�p��eX3D�4S՞@i���1^Z7M�d,�d�O����O���<�O����D�-��!�HɄ蜬��Ct��ZQ�σ;�1O>���
)B��]�� |91� r�R�e�	ҟp�	,$�j�qL<ͧ�?��lH�%�����Fv���B�Z�T�zt���'���'�8�7��~b,�F�䮟��B�١5:}rT�N�A��<p %a��$R�K�(�%	�t��
����2.J�n�����恙5_\]��Y�D���+I�2c�D��~y��'�^ĳeD�51=���уQ�x醐���P�\G��ɟ���[���?y��Ot���(I�2р�2
X��5 �T���'(2�'�U�؊Bj��� �@��P�~��҇/�~Q4	��V��������oy��'�"ၥU�R��Yӈ�¤���]i��H�\ծ꓈?����?���?9'%��x훖�'����&�ph���ұ?J���Ⱥ��6m�O��d�O���?9bP�|j��~"� %P�t)F.��Sp�ޣ�MC���?����?Q�F�4tI���'�'��A	�}ܒ��q�/L�Di����<Vږ7��O���?��fQ�|����4��F�C<i��oT�ISz����џ�M����?��a��A�f�'Q2�'����OGr�G!R�L@K"�P�T���A1#Y�Dވ��?�`C�?���?�,�d�O�Dڶ�\�R7��P��V+'g��C�4ZRƩ�b�iR�'���O��t�'S��'��u(��'i������9Y����owӰA����O�O�3���O=a�(\=3+�ʑ��B#��ɣ&��������q��Kݴ�?���?9���?��)+zt$��$WX| ���J���'��ɂX��|:��?i���|�����>bd�Sjȴ'�-���i���VK�L7��O���OX���i���O@��uC;m�
�s�(L_���qW��C�z����Ο0�I矰��n��ʗk.� �#��Ad��i/�x81�b� �D�O����OQ�O���ӟ�E٠="��f0\���M��t�	��	���۟4�O�����fӚ�xE�H���b쒱Qհ炅�Y������柴�Ijyr�'��軘O��}��K����6�HGH,��m�V�$�O@��O��zN|[�Q?M��*/̌��'HH|�R���w�nؓߴ�?1+O����O�����d��|n&nQ��4i޹. ���fǛ36��7m�O��$�<��Ҵ\��S��	�?WB%F5�X�oA$k�$�!���a϶��?����?-klP���?��r��v.$�d/SM2`c2�z�����O�Ah�b�Ʀ]����T���?���ş �ciZ�%{d�>���A�����OZ(��Oz�O�	.��d�+�<�j��٧&�t��FML��MS4�Y0���'�R�'����O���'�rI�%Zr9W)�b�	b��y%�i�)�F�'R�'҄�'��'�?y�ϐ'Ƞ��b���,Yi3�X3*���'��'9��)e���D�Op��O����rd)�6HC̙C�~y�Ѻi��R��Z�%t��?a��?yd�M?3�!��OL�fԖ�3ūG�x��'��QQ�z�N���Oj���OJ\�O��$]�J�J����{ӒQ��iY�'�4I��'�2�'�r�'�X>%³�I�Il��*��,S�&���-
Æ�ܴ�?1���?���4��Snyr�'���P�ѷ0�zqr���7�`�!V����y�\���	��I�8�ɰz�u{�4
��l���^�ΐҶb-u�����i(B�'���'vr]�����Y���5%��Ԡ2��^�����d�X����۴�?1���?����?���15at�ir�'>���'�,4}�G'8w�$qLk�����O����<��]����'�?	�'�\�� jJ}�����e�A�ٴ�?1���?���z���B��it��'���O�0� ��U�/[*����Ν�0�B�a�^���<��<�'���|nZ%�J�q`e�Y��H�ǁ)`��7�O��$
��5l����	ן���?-���RP�Y
Q� lY�"��HI �O��dT�h���O.��|�J?����;@!�m��@ɲEXl-!��}Ө8�����u�	ԟ��	�?��ǟ��I۟$q��fr��J�j_VleJ��M�4k"�?���4������3"���`f�ukr��J�?u�H lZ�������۴��M����?����?a�Ӻ��n�0T=̄+�)|�@�N�צy��Yy_��yʟ��D�O��D�0 ��%Z$F�I��P޴k�V-m���Ҧ)���M����?����?9W?���]�fك��J�֌�c
%G��xoZ��	��y�`�'���'3��'G�*Y�T�f� /�J�J��V��xC��1%v�����O��D�Od��O���ȟ��"(ڟ-����4�ۚ�=��ּl<j�?����?1���?A��	�0�ڠ�i~���ѣL*2�p�$%) ~�p���zӖ���Of���O~���<��G`��'e�iGk9q�x��g��79?4={R�`�I����Cy�!P�
����b^�{���8��U;�����ȦI�I[��L�	}��t�$,i�<��2�8!YU�ϥR���'RS���藎��'�?�'a��E+6i]1I���f 0�N� 4�x�''Be��yr�|����y0/ڧ��]Ӥe�5k,�G�i��=�����4m����Ӣ����T\Z�Ǝg�AQa��/Z�o�H�I�f�
"<�~r�/V�,��1��?^]h``���h垉�Mk��?9���Ɯx"�'��5�'n�U�G�D�v�l�w$`Ӓ�8"2Od�O��?	�ɬ)� ��G�T+��jP�ߐDj�=�ܴ�?���?9�j��;��'�b�'g����P�EǏ�V��H�#�
�8����|�U�kp�P���OL�+P��@�
ڴ3T�aYgf��h�:7��O��ӆ��q�	蟔�	o�i��`� X�_KИ*I֓*�j��%i�>ق�_?���?����?Y.O���[u�h����� 	�W@�%�h�Iğ�$�l�	ğ��V�G鰤�� %r�t�@�?y�FT��jy��'�b�'��I0{��Q��O�B�b��(��h�-W#-(�J�Ol�d�O:�On�D�O�����O���(�~6��g@�G��ܫ6a}��'+��'���h����I|�2��Iyn��M '-�mY�L��K��&�'N�'�2�'�B<[��D�52�Kԝ����`m_�'` ��4�?a����D���'>����?�� `�D	V������L#R��đxb�'��g�l���|��d�CO=t������*��:��i��I�:T
�4}+����������	(89�ݠ)F%.zY�c���!0��'uB�8s|B�|��D�ɐXS��AK3����Q����M�B�b;��'���'$��'���O��b��6/���3�Eq`L���ϐæ��BJx��&�"|
�9�4��v�A�2uv�#�$]H�K�M��?!��9tH�U�x2�'R�O,����Wl�)*V���`H���i��'�Θ(���	~>�d�O�!*�/�9 1��A��2A1a榡�	;�,�IK<ͧ�(O
\y�KO�P@�NߛcKD� �in�	����'ZB�'��^�l¢�%B�|x�b�
y��\�am��9$�yH<����hO��$�>���
�mO�E�6	 �	�W���Q��O�ʓ�?���?�*O�Y9�a�|z��ո��s�mĹkN�iiT}��'bў��'��o�zUJ�e��xq�U�^Ė���Y�l��ןЖ'T¢�ޢ,���dJ�!M"�E��@���#��0�^yo��\%��զ���.��=@��.�V�	�~y��(���3GKP���'��S��K�>��'�?Y���j��5��y����`d�#�x��'*�m���O�S$�=:�١7���pi��4y`6͠<1�"E�+����~Z��z5���a�CBה]�A^Hr-�Pd�B���O�l���)��0C��h�7	�8��kĄSK�H6͊!�o̟4�I��H�+���?�E��n���1(��Y$���V����O>u��7�"�q�2I3P$��΄w	� ܴ�?���?yc& 9|��F�'5��'���u' Ҽa|��kAKp�n���	[��M�O>9�c��<�O+��'n"oX��u �4�t�B���l�6��OV�[qFIΦU�I�P���hɩ���	�tA 57oC�
�.�;3�"Kx�(�����<�	ޟ��	�ؗO] �l��TѲ��]�z�8�u�;8 7��O|���OL�`�T���I���� Z+P���f.��h_Ҥ�ib�x�	؟��I՟���ǟ���,W���4P8�.�TsV�z��zpS6�iL�'�R�'�2[�����b����-p�J@KG��V�� z����}��t)۴�?����?��.e�d�ƀa޴�?���m�Hш�O\�d�c�(Aܘ[�iH��'~r\�$�ɗ]C��S���l匉�R�U��X�Q�V��	m����IߟX�ɽe�Թߴ�?���?Y�'k�~�ok�;��ī0�гiC�X�l����c�i>7�גA���5�U*lLX�
@`��K
�&�'��"E�Z�6M�O���O���f��.@`n�`F-̥1:\���k�>6��'`��LK"�'��i>I���i��/X�N� �&��d���s��i\pQ�ufyӈ�$�O���>���On���O����,� :0ph��?ڀ��D���0��JƟ�Ipy�O�Oe�͉=>�]�������Z�ϖ$Hl7��O����O�L{sV�U�I���I͟��i��AF;{�.@2g1 N�؃(j�����<�P��<�OJ��'�RFݮ6o>���NtM��Z�s�\6��O�$P3i]����̟��	̟�˭���I��(���	�s^!�E>I��0a�̓���Ot��O���O��#':SGrdB���(A&�$��Q�j�oΟL��՟��I�����<A��)Q�U�P/Y�&<��rIK#� рB�<	��?����?����I>O�lZ�z�ƴ0�]�MC|�ڳǓ�7�J,R�4�?��?���?9)O��䎶5&�I��:M0�����0��D�����6�9�'W��'�r�'"�r��7��O�$��YJ�t�&�I�h����"�Bb���n�Ɵx��ٟ��'�Bۏ��4^�L��lE�o�jIp%�3FC^@����M���?q���?����6ܛ6�'���'�T難Fw������*0�`YQ��&g�*7�*�6[����3~���S�Ĕ���4�t	� b^�UY��5T�m����I��<[�4�?����?����:��""	q��G�/J���K�t��=K W�X���5����	��0�	g���~BvO�*��yз�ٹE(��g+��ua�ś��M��?������'�?Q��?RͥJL��҅L�(ta��D;/k�v.M�\�B�'4�i>�&?���3&��txgҌUU���ND b�Xش�?����?IV�l��'���'����u'mC)Pre��A
���VƁ���'�� �y��'���Ot��F�W�{v,�Y��m�}i%�i�2��1y��'���'�?IK>�F� 7-���åꐍ8��r�)�]�'���O����O���<���
t.���ʑ.{I&�r3�C +�|��p�x��'7�|��'62.��{�6���`��u+FY�E��YI��k�yb�'��'��/�x�ҞOk�p�u�Ι_ TD�
�H�(|�O���O8�O��$~��YCW��R�DZ�ly�P��>;�$!� �>����?a���?I��6c:H���?A��%Ҫ`�`@3Z)z�����*7s�33�izB�|r�'{��8S�O�3ROʤO\�� Sメ�Lƴi[��'e�Ʉ]����������O���L�a ��K�DE]����؆a���l�V��?����ƞ�B��֜{}b�;B�
U0��ĸi�b�'ZxYc�'���'���O����5�	�|Wȑ;��|��(
Q�
 �M{����7-���A�#�|PFpQ@��g��x(t.P�!��`���WӪa��hT��!��7{�����,/� �yƤ��IX*I��!m� ��Ƒ'~r`<��I�~�����;'TQ)�iQ471�!!a�r�l3��t�N��R@�..H���'$��GjV:#ܨa�c��[4�ϙ�|A�������pp|��ѥ��je�;Yc �@��O2d�Zq�\�`|�;ug�XxhZd�T/_�JE�O�I�^=Q�$���VP��U�8�N���ß��	��T�]w�R�'��I b'����
Xf�5SV(ڙX��P#4�7��!�w@+e�J���,'���AS��!s2�D>IV����$Z�i(�U*'O���D�$
�đ��O#;�<�v��Y�T5C��'����d��u�>	�P��, �̱+@�k/!򤅉�t���{���PO�%1O%�>�'mAț�'y���?4�R��7z4��5�L�\X��'������'��3��$3a�'>�',�$��ӌnV����L}���l\b��?����1��S
��㦈r8��Z�H�OI%��1��� ö�J��`ն�x�"O�A���@�L6��P���,�z���O�nZIo��[����Öv����b�ta%f܀�M���?A,�t����O~#�BN%���3�I�np�p릦�O$���P�D(�|�'fH\��C^�h	��4�
oh[M��h�� �S�'p���"s_��C[�i�]�O���'ВO񟪴Ȳl�1u�Uy��O/��H�"OhT*b����Z܋;�HI��'��#=Y4��D���1D��d�P
�Gr�&�'/�'���t�Ƒ$���'����y���Mz��I,o�u��+Y�,p�!���J���䓌kْʣ�|R� ���@摍_��u��K�5'���)�9
��䑌n���r��L>�E�C�N�*e	
+G�����bߖJU�'�����S�g�?G�l8ʀ��&r#"��ah�zB䉥&�`� ET�PF:}�'�1>̰�	^��"|�ĉ!.?��q���cިiT�^3"�
�"�'���?���?��,���O���r>S�ۏ*����ֱc)6MY�C�^�t�8	�<H��t�%vń�jw�O^�ԨQ�B2O%��ST.0L�4�*CF�d
�mB�-ط
z]KP� U���p�'@��J�� ��c	�#⦰S� ;�ybC
�/д�j�)�M�fq�����'T�b������M3��?��ZV���R���7U ������?!��6��="��?Y�OP=H����	K!���Z�e� �q��U�\"ȇ�I�\9^㟌c�^�^?��w�
ঐ0	 Ot�"�'?bO$=R��+�(����2@�L�"O���,��r�9��eݘ�#�O�ul@}�|���0�&lcN�<�lc��a�M[��?a+���·K�O,4�L �\�iQ�I��OF�����O���X����g�1)��i ��ԟʧ��)������@�A)QfH�C��W��q� {G����yrE_��H��(�c�c�L��Q��v=�S�>�գ�֟dsL>�
��#����<���
��h�<Ad��+L�x�A!B�x�Ĉ
�"�h������}�Zl����
�t�;u�V�|-��o�ɟ�Iȟ�1���[�ʝ��ԟh�Iޟ�=�>�Q�Cަ:����!C,�$��<���Jx�4y���������Y�g�LQ"�$�	�`kn��� �- �X��F��u���`�S*��c��0`,�Oq��'�:5*v��5z6Բ4��`���'���iD,
�|IHe%����O�Ez��I�&�8i���5r"E{Ra!#��X9e��7(��$�O ���O0m�;�?Y�����R8I��H�?haɣ䓀-�����'��T�y��D�ԒZ�| ����x" �Z~e��a��6�� e�@i�a�鐯ZB� ��%H%��A1���ybb�Z��u��e��Bĺ�N
%��'u�c��E��M��?!Ҍ�-dvh�Y���-
H�"�F;�?���KJ�����?��O1�����5�f!r��*	���.�1I*���	0 Ǡ�XA����V�P�d��ӇC:OR���'��OЙRt���E��[&F��jG"O��k��q����%�;,ˢ �'O�l��#hĸj��9ya���q�7i4b�4	dg��M����?�.���8pa�O�T��)B�Lu0��#~��Q�`�O(��֖C����D/1�|:/O��HĜ䔑c� O+Zl��薟>�j��b���<�������&��B)IB8�U�s�}����"�'�R�'Y�� 6�c���,�⤻w��2�|�y���OT���&�:ݠ�-�0Sڊ0P���ax"9�ۆѩ�c� :T"��!N�*	@��á�i���'"��C��ʃ�'
��'���w�z�R. �@|p�gȬl]2��p
+�$@0[<����|2b�xQ�Hd�� 7h.��R���[��O�q�A&�����:z!�fe�0 l�L9p�˃r�6,і�i;�6�O&��� �Oq��Iʟ�Jq�:#�dm�4F$v(�\)�m�fh<���F	|V� ��G��`���W~��!���<!d�+\]���$�8�Y��>�8�i׊�?���?a��^\�N�O��Du>���*K&v���% �܈q�=%�C�ɐ|J�u�&<Ήy�O��Bð��7�<���uK�D:��0��ҷu�@IHVJ��l����L؟tb0�d�r���]��D�+5.1D��s0�ٛ7h `:�c��N�~%r�:�I$��'p8�Vil����OR��V�Px��)��o���6P��O.���#z���$�O.據O��$8���O�Đ�"���W�����"sN�x2����'��ht%�z���!U�2jha�+gt���ēW���(o<h{�I�c�
���t�(d��mƀWI����#oF�D�������G��E�]'iu�1Y�#G	�'@��0�g�V�d�O��'��$S����J��Vli���ӮL"S^����?A���?�y*��I�F0����âc�6Mc0*�tG��'� ݻ���	� �P����T>�y���;R��%��l�I3��S����\��!�'!�M2wc�1��V�.5H�Oh�p���8q��%�HOlpxv� ����-iTp��FǦ������G�)�F���h�	���i�!`C(ś]<�B�b�#�N�D̓�� �2�׾[�+Al�7H�|$�|JJ<�Aq�F�ȗ�ӛ+��Bb둬�P$h����T6�m��V�$��I�}jE�Ky��������䙔2:��C�$̀�ޒO��C������D/+FmDV��u�Bd�(c�д��>v�ՓVF�.Ny�AoC�A�L�'�#=E���&�^��rg6x.nu:Ս҉1:�m�/v��'��'�\�]ߟ �	�|Җ�
#�ܶbO¾��u�͓�ud,81��	�%֌P�lX�F��m:��$�4_Rh�e4Y�l<�!'��2k�#�=O�l�3�+H�"���>��<���5h;�92 �CF�c�#������Vsrp�u��1�ȅLκC[�Ņȓ5�=x�&�"���#��[�+XJ��<�c���d��\n՟����	����r�ȕ����1*����	՟|�b+]ڟ(���|r9�q 3(�:�t�3fD
C��M{uM�2(p��-ʄ��d.��� t�,ZXؔ��✳F������7�t�	*T�XLs	�#�`l�I�M#��i�\�3��Qa �R�cɖMAGIƦ{�	����?E��-^�F��Y�A��L|�CA �xb�a��8�Y�A�~!	�@�=[���;O��Hڤ=!�E/�?�����#���ȟdE��蜷cZ^�a�D�?@�����O�eBec�Ob��g~b�α2��K� �	(���t Ӊ��ɍ$<�"<�jfȋ6�,u��¦༜�A�Rf�d��M%����ْq��t��&(��9	�C7P�!��3~H4���Y)3g1Aく�NaxR)�N��)v+���)��W�	Ȥ�i�r�'��*���hH��'��'��w	��[X`$��)§[#`�Ja���S��0=�q%T:f�xD0���!E�ܡ�&�Dܓm���dt�>��fG�6F������ZNb�mZ��Ms�j(�e(�S�gyB�'E\��-N�o,l����-p�:d0RO.�آ�@L����K�-'Ө��7��� ����|R-O<�����=j�r�x�*��(�:��Z�Wy�����O ���O��������?i�O�U����7�vE���N%*�Bƛ��x�J�,ڒT󇧉�&Q��cZ�_+�B
�'ݚTK��dN�p�#�K�Y�`��&���?Q��'G��@"��%{��r�ʖ+�>|��'< �3%��G.�8a�� w�|)�y(���PA$�	ڴ�?��VĐ��##8�9�G��*�"H����?!�/G�?����T�8�?iI>��)i�z�B�U�0�T�`�X8�����5�ɓG�����yFPDȰ`L�+k���LF" #�dD�[v��)[#j�랈U�!�� �����ϗH�����(��}��Ohpo���:�,�4��{l�8?ۺc��6����M���?I,��!���O�q4kS4h����L�<����׆�O��d<o�P��m��l/����I�|*񤕹W�2I��;~n�)��C���]\�AfU'Jp"Ҫ^�j����5��J�x�i'�c�$N�51�p�<�nZ���������Gg��3�W�lp�5NG\��?A�Z����955^�;�-�/�d��7�HOFX!G��a?\(�P�Âe*��!���qq����O����hNxLJ��Oh���O8��պ{�c��t�R�9�ʛ�?��F����'U(88�l���!j���A#k�f��=���\x�D0���}(]�1�Y1�Ʊ�#�P����ơ�)�3���;����|�2UP��S My!�,lƂ��B������[w_�I��HO>m1��V
oZV�[coF;t���PC֗`|�E��T��l�	ǟ<�I��ug�'��7�M�ƛ����H� �(ṡ��2U!�$S�8Zhٲ�b�&���M�2*
,`
�Ofɲt�8GWN ���װi\�t���J5���$�O�uA�O�_���!B#R�prV"O�Lr�� w����!�� ��^^�$�D���i�b�'ᄠ0E�ZT����,����#��'��Q^�R�'��	�b��|b�Q�D��� ��V������p<)�HK[�T����#�V�Kp�b�Ǉ���܅�I�Y�&�D�^�	#}+<e��Î���=x�́,��B�	>�J��g��;_���7G_���C�ɪ�M�� P�a�3�}��DٷKl�'����'��R���Ƨ�ԟ��� `��uS�݂Y�� ������ɳD��)��FL�Is��Oʘ;w�Ǩc�>8��.��@���>Ѷ�Q|�[s��J�hA1fJ���O�����AE(�A��XA_�j#}r.�=�?y�i��6m�O`������	\U cEΥk�2(��i��)�D�?�H>�e�� ���`�=G.�5��@���O��?����G�f��'�N�,���nѣK����'���'�����`����'9���y7��i���5�D�x�13�`۫lB^����<���ٙ�EC,�3�����!˔mJ.T����
�F�ZdkҊ�ny'I�h���}&�Đ4.Ӓs�AP�Ɯ+=<�YAKV���'y|X��S��\�IΟ�
��\3YWP�h�\�{�Vi�`I
mh<1�lݬN�i��M�!�\"D��T~�*$�S��[�ܚ���ՎAأ��;>&M�[�z�@�KYğ��������u��'tr>���aG�Y^"C�?.I�5�� �`tv�(�c�:2!�@�qB2<O�hI��3,��q�_�-�"�*l���r�%���+� ��sty˕�~�{�{��T�Ɖ�6LҪY���6��9B$�����aRdU�Q���)��<@3���JQ?�y2%Ď%�
C ��3,��P���'��7$��ge��o�ȟT�ɇIFhXR��S_��Dg��,���PA�_�t��ɟl8@���'~��G��:�l���FH!J7��2�hW�ᖃ�������-����F*,�(!􏜥��m�� hS<P��ޜ ���6�֖,���e��O�$���e�O�l��M������#bOt?�pSe��%OO,�+)O��D0�)�'h�p(���{ƶ@!�H�j풎����M��Q�O�~0Y�"A'��S&ȶ&�"^������M��?�/���$�O��XIľ;���xc�O�N���P��O��� �2dK7�D�3hzl9���ʧ����`Ol �����5�( k�a�$T���C%6h@8P�Ĕpe֨+Xwff5I�h����4��Q��<�E�1A��H�DA���	
`����1�)�S?;����g䕂T�6U9�(^�@��B�I3jS.Mxg�V#Ep��1II����D�'��h͜�A���"�k	�!e��YCHkӶ���O����BlzyzN�Oz���O��4���g 4C����Gh"�*��E�jN�D!�����	G���UX�b>�O�[2��1>�xx�f��3�� ˤO©��a
�.)��U��ʌ?6��J *d����Ӟw�m8@,��B@ԙ��W�~�h��1��W�~
��L>�F�%t5�,��g;�4�S''�K�<�D���]Fe���ҔmA�H��.�_~n2��|�N>1 CU�S��� �杊E�1�sd�O���ѡD"�O���O�DT�S���?��O�̘$��:�$}�f��(>-���@�{x���WR�)���'E�Q��3c�1GPo���nT�+�``#b�t�!�ē�H���(��:
C��=IGc�4������<zR�xP�N#�d��I��?QV#W05^�i�
�yu�����	I�<� ���#�J$!�0� 0$d��5���Ϧ�%���k�.�M����?QrF�L�|���T9H��ɪ�K��?I��=�����?9�O͢Q)Cԣ^�MS�4Di 6-� % �+r��?�YX��L�m��x�HE�r ��V�W�n�ʶ�*D�u1�L,B��\8w�X�a/�A�R
����/Y�ig�=��2�M{�i1"OR*<�$ˌ!",�Ђ��@'x��I��?E�ğ:-��q!E�����q�5�x�+`�z�y�͈>*��WCF�/���0��O��>yص���i;r�'p��3q|��I8t8���'f`�SV��K�@���؟�ap $eIZ�7]�6z�5 �S�$U>���a�	
vz H���okN����1}���a� D+1�hI2ǎ:�Z,1�j��g���[���8�Ja��k ��C�+�<i� � �>Y�������E�I�3-z��9"ǋ�i�TŚYPA�t�3���p��1�"�Q�Ƒ� ��Ҵ�C�����Ru�'�THj�a�7G����f8S��� wme�,���O���ו�p� �O�D�O\�4�tT�V�W7+g�K��K'��1�K�K���! V�e1d�b��Q)�vb>9'�䰤T;��c��(X�=�E��[	�! ��0 rx(�ÂV:k4��>	$�l;d�؋^W*\�H΀@�Ti�EcI��Ms���?Y0����?�'�?I��?���?�dY�o�r�)�`��~LjV���x��'�phdh�vгC�ݾ��$Q�'�D듃��2D|�D���0k+]�G�;YPJ���L�	͈�$�Ox���O�@���?����t�d��`������j5(g�΀8��\b�'�@�j$>��j�=#$�\�U���xr��G��p��eN8�`a3��$H�LX�3]a"�M��Ԉ"�g�^f;4� �yR*?L�bY ��Y�[�:���-�)��'D�b�T�Dj[��M����?C�!a�F�T�F�a���y�eE��?���
� z��?i�O����c�Pᄭ8��=$�L����ٜZE�I ���D��l�@#?9Pj!v$�lQ&�B�u�$���@"8��R3:T�h��ˋ�Gv�Xa��p��D����ش�?ib�͢<EfA���V&��3�i�����O��"|��#	�Fl���>��<�U)Yf<I5�id��H�@Qrsl0���*0L�ӛ'z剜w�ڠ8�NOٟ`��H��
��;ib`�����DI�"1H�"��)~��'��=(�$�5�1O�oyA�ah���b.N&O��  GGZ���z���8#)"�)�S?B?<����+���hA�5�t�')����ӂ�i?
7��O@�?�%E�,��M�V�Y*����2��ȟH��	�
���S��V���ha��,?���ğ`�'Y���F/ ���� HU�~����4�?!��?�SM2# �[���?I��?���?��(��s?(�jUa���Éy"�����<I��?�D��@��$�.��&ƙF�~x�ن�	�$�xQ��
��m�J�˷g�|�(lBJ>��gğ�>�O��P�L�2�xL�5L�N�\%)�"OD��EX�z�]�A
�!/����A��ᓲ9p�1�s�ݜ#)v�A���&|�Ğ���b4N�O\�$�Oj��ߺ���?I�O�,-�q��J|��G�&_�&�A�G�)��0�eH+�0>����H�vU�]�|À���!"���ׅR$V�Ntڅh%�O,���L����� m0މ����%u��'�2Q�tI�6-��a��
4<�'�$\�H��G�>��$G
l@R(r�yҨ5���yr1bݴ�?���S`��T���3��}b6D��e?������?�f���?	���$D���?1N>)`���t]8,�!^�+Xڜ"�	i8�h�s�(�	n��њlmW����aϣ~����U�m>�Q}Ԥ���yj��6 G�1o!�ΐ*PH�����q��y�Pa��{G!����-� |�2EEݩ)��e"o(�ɪJѪa*ߴ�?y���TMNd�dJ���pڐ(�?�P��V��4����O����O�b��g~��"$b�ru,�\9��mҦ�􉽻������	�x��'��b��S�G�K�"\��	t�S��[�Ւ��	�Jq�q�R:�����u4	��ۅ�y�ō=v=�<�቗�HO��Ґ�F�Lvr�bF3	�9�gK����I�����X�)���Ο���ԟ,�i���2�ɫX�и��V�k~d���AСSP�'�&L�ćǰ����|d��A�ݽ=s̠"s�X)M{,�+�AFf���*b�.�J��L>aQ�O`�x;�	G2�ܹ��B�?����?q#�+�?�}�'<�l���ů/?�ja����	С��;������C�`v�̳4�E�kV�	8�HO��Ty
� ~�r�ؔ}����� ����u%W�h���� �O��$�OR��Ժ���?ɝO�|����Jl$ a�*M�:-��Q;�p���b��t����Oׄ|�p*ې���Qj��o�Dp:t�
�~�)B4ή(��Ɍe�D�[��S/l( }:@�Q�m��@A��O��n�Mk���3��=GU4�H�G�Y\Ѣ���g�B�	x�*,��ɍ)6e�"���+�b����O�����xݴ�?���n�X��	�r�C
1 BY���?� ���?A����t�=��#�g��B��*��83�\��ۚRO�P8�˅xFp���)Y�=q!���e(�a��O��u��-��)��\�-�<����'����<�'[ ���D�5j���;'�ܱb�2M�'�f���j\7~9��QfI2��I
�'_�6M�{Upᄘ��Hp���Ӓ2:1O8�1un�Ҧ���ڟ��O�9��'C�u��aJ*N#�`V�Nu�L]x��'|2�PQ���e�ڍ&&:�S�t^>�a���7)8U�V�G�x�O!}�IS.,�ܭ+�"ۑ?U:Rj�D����>8����R!}R�Y7�?)%�|���iE9T���ӱ"�&d~��aI�:�y��ǩk�T�ұ-Ҕq1�E����/�0<�R�	���j+�#Z&�AzG�>3�Q�ߴ�?	��?��f8V:�����?���?ͻ0��
`�6l�F�ңm��Z|�`� 20���-\1����Ƨ�=��O��'�F�r��Q�b���f׺&G��To�;��bb �
1bZ	��O��'�YQćJ�9�Lt;�$ɀ��U�'��Ɂ���L>�3nT&9�b�y�"�D�X(�A�u�<�e��$[r��q&���?F0���m~�9�S�O� �!aÑ-}�0@!kɯ�p�C�H,+�����'���'$rAc���	���'ވ(s�  �;'�@�ІP�
.<S��+7O���$�(���$��t
u�ۘS6���H�5!�ԩ��MW�@u`Q8e� '�����Pw�'���d!��?H@�Ń��X4�1͘�?���'����L7:"$��E� �!��'�֡�N�"n����7KJ�	��A�y¤5�	�O��!aݴ�?��K+ `����d8xB�,Z�V��<���?� ��$�?���čޙ5��#�+ޮg����� ԥ%P"J�B�c�\���'�H�<���'�9�W�@%`$,�^m�$��+���[�j�5Q�)�"镑:�������?RǶ��у0�<���&�M��i��cF�x�^p8b"�&M8bl�)�6�	͟<�?E��Վ|� ��]�FK��Q�N̕�x�#j�8��t�6,�<=�g�Vۂ�(�6O ���$�c��?9����>$a,���t�L�3�fP�B\�۵b�"/���O&y��BI�Mx����>�O
��O�P����FnN�D	��H�'��,��zɳ���`���`#���'%r��2`���<��HY�cإO*y��'=�O��Q�ߛ'�2i�"���|B��ؖ"O|����]U B���)\�Qsf�'h#=9cB�6�Ja87Z� P��A��	3Ǜf�'�b�'c*�x�e�g��'a2��y����B�H�n �v�,��!(�83n1O��b�'��й7f��b���)_9���{�K����<9��Dq��M\(;HL�"�+����'OD��S�g�ɼq<��EY��� s���2	�~C�	�X
����#G��.SL�N�aq��"|��D""�j	Q��Ɵ��QRs�B�7����ۓ�?9��?�� ���O�i>��$,�,fRQTL�	.tB R(
C��
8����̬\,>1��&�=;c���?����b�u��<X׫zf*0cE嗼,�>��C؟\�s�J�v���!W�?n\3��7D����,ŏiJt9s���P�Z��%�:�I ��'n~X:F�k�V��O��1DE	k��T�zx���Ot����y�����O�擘\���S@~�ɭv��� �Q�^��˾jGr���J�I.DY�(Ī����:}�:�;� �%d��C���<��x�o���?�6�x�#�f���N ��q����y"�N�'C\�q�6P�@���׉�x�q��tq! �=z��Ex �źF�,�����A�&�m؟���v���W�(aB�C�i?t�X$lC*2�r���&���'ҸC�)G�+_�P^�(�+Fן�'��	F$]]H�XFĝf�}@T��H��&@8�`��5z�(U�g���"�*4@���D�
| ��sCUQPd���	�U(�:�������S�'Ql�h32lƝ|��|BdmE��%�ȓe~Xچ���B��DZg�3�nA��	��HO��@7G ;�bk�'�}��kqHO}�' ��n�����'<�'���� XMPc㟐3 tPi�c.���:�HX%q ���O�%q�+آT�1��'���
��
p���DO��WZnD[Ŭ%c��=i�')*u����b�g�ɣ|�
A��GPђ ׬�Z���4n?��9g���4��	 ��	e�͚��@�{g��=Zm��|�4h #㝆l��P��0��!�'&"=�&�irU�,S� )Zyr՛�ƃ>n���
��bݪt�#���|��ܟ��I��u��'�21���!#Bx�*�ᚳ6�^���a�Au!���8t�r	 T��` cl\6s��ձ3O| 4��C����!�#�|����+G��'<(�O��Q*�#� �mMBd�	�'8�
�	�#%�=��Ql�Y�yB.�ɍ��4�?��va�%�^'z". Y�ҵֺep���?Av�O�?i���TbS<�?	O>��oV�P#�L1r	V#zk`���\8��I�C$�ɒ1��8	g�G,"��\��Eؼ����Ĝ��"�|B�P�K>N�3�%Z�s�pU�e쓔�yr�\�K�Qu�٘?heb����x�Oc�J��f�A�QZ��J�G8��x���DE���|m���	v����y�Jě"��ђ,Ʒ%7=�d��7Y�2�'����E�O'�Пd���D�m],���:q�
L7D��A����HQX�����O,�"�1�^����)�T�Lr ����h�b�'�F<��V՛^ "|Z��\ERխݫ����aa�� �����$=�S�O������`'�P`�
�������M���i��dx�R���i�������U�ڼo⟐������D�b,$�	����Iȟ�]H���:�l�h�nO&1�L���؄�����i�]��������Ȁh(��]�4N�7�ȳ��
̔0����k�H����	����xe��r��=�,��G�/�4@G�|2��/�?�}&�0b�l.R�S��lb��g�3D�P�拦!^"|�����R]@f-?��)§P����)wT��F
"h���@�����z���?���?�����$�O��ӑ~^�]j�kGYV�`�)5XT�tk4�@r-�;K������ll����H��X��B�I:I�vI]�Wڀ�G�3����J�O �����v�@c#ߤ��)5�ڜ;�!�$YGRexB��m� �9���-�1O�D�>Q'�Y�5����'�҄��9���*���#w�	Q�	�G5��'Q��R��'�R5�\yKP�'}�'fB<;��7Fj$e���I(sY�� Ǔ)��9�?�ӬЏU�Jٻ�h[�5�X}c��c8��eo�OlM'���GK�gsVq�t�Ԙ[���kG.;D�Tb3OK�I�ɓ�_ $��T� �>����4z��Q�!	zz�A��UE"��<!U΂�WD���'�P>]�ǝ���)�k��0���ZRk�7C�ś��L۟x��*����	|�S��O�P�����2�HP{��ԙ����>�&�p���Oz ��C��K��l9��	��޹�H���r��O0�'��?�#閨m���tF��d	���<D�Y��)T�D��G�Dc�؅��.9O�\Ez­�\�`���`��{���F$D�8ب7��Oh���OH̲6����O
���O��A3^6�"&,��*ᜭ��ݓ@�b����-1<ONQ����J���M�p3t1��ģ/�az2N6A^ ��B(F��f�JW�5��'�n�j�S�g�`���Q-Z��y�g��4d��B�I���Ř)�P�$�k�������x_��"|�
�D�4�k� ޣ
6��D*I[�>��E ^?�?���?1��F����O6��p>q�'h.�U*���ւ諢"��>B�Ɉ;B�q)�c�Z�a
��W��Sl1�l	ǃ�1k���񅇨r�rx�0��0�P�d"�O|���-B���wM�|�����"O�<�q�޲3?dtiQb�!�����e�p,��`�iR�'眰 �EQ�8�
��(D�:�;��'�B+�5vj��'��)�gв�Ԁغv��hJ��'^�,��&Q�P�������?Kd%��g��er����G#6���OΟ�b�$	=Ol�JuM�~R�� O2� �'N<OȌai.v�|]I�fO�X+���D"O�!ar/��-S�\���+�\OV�n43J��EK��9�R(�)_��b�Lk��M����?*����E@�O�QW�H}(\YRB�,{� ����OL�� I�ɲf+_Q�|
,��  $8"e�7~����u��%��U:$�>ɧm�KrɂO>�J���&���m�է�QQ��t����O?�'��	� hт0ʵ!�"l�����L)[d!�d[C��� �&?!��˾�axb�8ғg�XT"�d޷ق}Ȑ�2�\�Zf�ior�'9��_5g�����'?��'�wKp\2d�G�cf	�W$I2]�\����ā)k��y�dD^�J��&��q�}ӓF�ڸ'�`Y��^�:��,��܁[�݉<v�ڋy��݉�?�}&�(;��N� !(Ҩ�"Ln�`E�'D�D1��+PҾ���U31%PuP�L%?���)�'x���(��ȹp5�Iz�F>)h܄�\����b�`u*�	�$��|�ȓyL��aVJ_� L4\R��W�Rڄ��EX&�"�ΘV箁HP�.���ȓZa<UiZ�`�)h1�P
T��ȓ^�Bu���s��Kf	Ɯ|�t�ȓ��U��	9c��C�-�?^��ԅȓ���&n8 [n`pK����̅�c#D(��)uI����j���J�5ӅÀ�?�$E���ۚ��4�ȓh�l�� �L�&�X�2&U�zM�d����U �֕��@ʳ�Wou�ȓ�dQ	��JF����-��H�b���vI�eC9&�|P�����`��-�ܘ��/C�N�j]����9a"���2eQ��#R�~�&�*�,�V9�ȓ[
6쨐1 Fe:q�*նt��&�$��U.���1���-c.��)�ͫ� ��3s����͏�.(��ȓ
�"�^.td; Cםdsr��ȓ9���"& ͕Q7��b�a��dX��ȓ����<SJ s�&	%wG����O��}���Y$��� �J�<��ȓF�`�1�g�&�� 	nK����"\��8�C�g�Вt��R3��2��C��]�H"�9R��Mg�$|��`��&�����(i3�La
GV�<9CIȳF���S�s2|I���Z�<I��#=z�%2��L
{	�-���V��d*�-M�w&���LȾVK�<[�C�V����jB�kH��i��'0<�i1Q��g��x�k�*؟3�9@��X%ޔF|��	�5�^��jVZy�d� k��[K�� ��;+֦����R?Y��~/�">�fe
;(�J k�ؖ"�d �)��DZH�r&�	�Q"O���ٴgnE����<I�'��XYl  Ǧ��!�m�F��N������8V�B�]/�Bu�$L�81b=O��+�	��
;<)��*"Xi`��R�9�'lqbq��erPi�e3X������ �}Ǧd�A송i�ԯ�<�p��sdZ�]Dnx�.�}:���hO������K��dH�	�mh�!�� ���p ]�t@0؂.Ql?-��O��A�&D�^
�TQ�/6Q�0A��>4���i>���Eġo����ݘ�w�A�Z��Y�'P4�`9��;��p��*�kv��n��0�%�)\E,]$B˞P](MX��B����LZ ���B]��Ҷ'Dw�$��d���bڷ���A�
�u`�Exr�,yI�"Ք/��@�w��5�?��'h4�%Uk!|xˆe�te��`�V�2Pʓy�Д�ƃ�?�g%�//Y��	oZT	�6i�dk����s�G�Epb��X�v�x �	�G���[P�֝�)x����B�$'���r�-5����Z�(�Iv꘺j��̓i�x�g�D�d=a��� �<34c]4x�`קL�}M�9nZ8k`I�@�36kX?���>��E�]�A���)xV!�CJť�?�1$�9ٸ-��o%ړU���a�7Ml��&�שv�@!�Z�`UJ7Č��'i�OQJ+���N!/f����	`����4��"=����5w�l�֌Jl�MCwi��9�x3���U���D�=cRрwƐ:O"j�YI<�缟�F%,Ѩ�H߸�?1�ƃ���gD�)!�����HL��,C�䟸Pv��,ĵ2�cْpD�I�cL�	a����?O��E(�������%��8�O\ղ����(`��'��� �۟|���˜�%&�<��K�*r�#�@�1:�(Xf*�5�$���'���'Z
���#W�s��ѣ-��ABUˣ�'�rD;S�<}Z���㉖B+~e��ӎ@�, �"*�q�IL��'�2O���/����#� Hd��I�54���I% O$-0D�'�¬�e؜.�* {&a�j�2�{��K�F���3	[��Hx"� �_ڼ�$�h���O��Cj�M���ٟ�:���?)BC�1j  ��KP�����$?�净v����3�(��p"�I���x���vvl͚Q@*w��I0�ʺ�~bcƬr�R��F�1�?Y�G����D��Hƶ���MH�\���G�Xsxً`d��k܄�1'��|T�$�O�K�cO2q�1�:��S,?*��I��N�Dp�0��xE��j�t��#>�� ^8Fc�tjQEϯr���w`�3i����N�y���$���	�q��.��P:��'�d��[c?��Qsɗ\#Z�BaOȌ>����=�@o��;��[�Q�t��#lV?"�H@���W��ypfߓA���P�iM�;Qd�N�%#h�6 �^j.���/�"��`�^Rwa���g�Vh�M���۱J�2B�~4oڪ@퀴�5j�!1�V�QB�ɯ&O��I�^��8R��~9�dT�'8 z�#�rI�M1p_6W�NeY���W��"�D�4C��dqq�D�E/�3��?�*���&"�(!��*-1�\��R��?!�B�&B����y���n��63��R���2�M�OG��!#��%�F�8#L(4v��\b��3�"H�/4Q��1ƌR�yG��N�d�@�^�d�h�+�nV�X�^���@ցl�������"Y�x�kUnW���ca~�*���0�o�
�X#=���ڑp�P��uΙ�IʘM�3L��<Iw�����EÖM�� Ux���c����X�%�}��ј�lC04pc�K�Dk�M���'��i�(7iZ�Y�
�<[ι���
�p1����5* ͱ��Tn�h% 
G�J�%?i8�+S�;>8MA�,EpS�S����;2�	�$�Z��&��*]%D�)�=_���?���>�d�`'��Q@&������M��/�쟄�
Ɇ4T\yyM|J�lp��ʓ5v	x �D̀?)vԠ��΋z-�`���D��fO:�p=�1]�r��a,�h&�m[���|c�y� ׹YNr@�b��OP(�3��w�Ӗ��i>�2��P������}�^\��',O$���_9Cz��"歟����"!!�Z�+B�A+�/�x8�!`� u����&�	�B������?RKk�4�ݣ�Y	R��\�J%@���^���w͛�j l2��w(�pV�$}�d�/4Bmع�:�c�(PfQT�ߓ�?)��:2wz��m�0u�<�FeșV2:�a��&�	�8��j��͊P^\���K�`��ъ��f�ܭ
I<��R9����$� P��m\�v�J�R���-iX�Ѓ`6OX�ͻNT�	1����0��jWV�͓��J~Z���<2� G	�C��8�"�]]D� �3Ή��O�p0�Y4l�� &��!�NE���iʹti�故j�F| ��9z�|�0���Ti�J�;a���Q�� u��_�L5�֭՛6,���B�S�8�*-�rO(��R���ID(yD�yF��)[��Fz��bT	X� ��I�8�0��A�?A%N��5��H�P�C/c�e���z�'����A��AR�ш%�����ˈl�$H �.|O��ܴK6��s'��;t�\�kī+s��L�`��Y���0�w���잏^����"N��R�q�
Ó w|��'��m��E`�~�b�"�-O����G�)4�2=��	3TIlx�a�U8~�L�S��(�b6��v7�}ˢ���%�<��A�"k`�2>�1�'EX��u�Kv?�D�!r����if{��L�H6n����,r�h�nƑw8Ε�`���ܡ�����*��}̓�:lj1�TDd�$jQ#!�H�ɆV�P0HAlP	"�3j��Y :�>)��ҎgM��Ê&d�z1���P�2��	;z������v�)���So4%&q.��q�cTv�H:�NCA�џ�2G�I���@P�w�|�Ă�#=8l��J <&Kҙ+V�ŧ��DV:!�,He�0�9O-Ja�@!v_:hE��#D0�m�głM��	@�=�I�/��c�iF�R�E�5K�x�	mc�0s��|�0$/[��O'q��J�e�w�	#g���H�mїI�0A�α{����W��x;R.؅Z䈃�7S�{����ce�\�A�Q�x��q1�'_<y8T"��:Ĝ勅�����d�p��͸|ڠ�s��Ѿ`�r >~Ѝɣ�]�	����O�x�6j��5��sM[K�� 6)�g?	�Ȗ#H�2X[�k�i��#:u��U�Pē'�D�r�X�M���h�Sq5Op%x���"-�D�]�\����Uʌ�@DX��#1( ڕ�'�G���D�?�A ���'9@֢D)��,S�Ś�NՌhk�Y��-���"oVDt�bLK�7M:���g�/H�(��L�]	��;�i	8_<�\k5��}_@�ڗDéCY���O����'���~��ەc�y�:�x��a��t,t (��Z�t��8�'�l�-t �ks�X
�лË�/h��� 'Y�
���i�dc�$F�\8"���C�v±b�
�Obuȁ+�z���	f+ea��	Zˢ\��$�S�L@!1��0uH ��$ڥ-��:�6[BR�":"�	�����u�A�	f�)��ӈ��lY�&@�j�T�b2�'��]#A�ʤ�K@�n�F- ���m�D4��D
\��	0_�Mj�֟��,Op��B]x�Vh�z�@h2,��tk�aH�+:���9J� �\�YGS�Q(��� ��E�p *b8t����yf�aJ��S�,G��!�_����!����]A�`A�h��(j! �*y��T;�I2T;��c�剂V�P����\�#~�%A�Kv��d��6�:<�Q(�}�`���0O�,A�N�)m8�LB�Y	VIx�'o��ЂK�$:������-C��$.A��!���o��� /ӎ8,�˓'<)$j��l{b���G8�']�����ZI�jI�%�?Z>�I�,�<o�����_�~`i��.Ҽ��F+Z��l���03^:$�و �촣gĵ����%٧@��ʧ��$ɇ �C`�	/�hK���!��d�L |5�c��3 O-1��1�A$Y>؆M���� �hBge�D0�d�á�!Wvq@#%�6T�aK�E�{�rm'4ҢiAai�$�Z����B�'���1�@�bu���H���P�"�;S���(R��ʎ�e��/���޳\j�I2�aQ->��(9� I�eC��ڢV��� ��#�R��'9�,hYw5Q�D�ף�Q��Q36 :����+S�{�Z�A#
#s ��jF�/��E���?�~���1.R�hr���HBH$��O�?~h<�&m9O�AF*��>����d��%��!ñ`��tP3�pkF�K�lQ":�2	b2O���bl>%��O�uR7�?���H�`I�#�������Z��oU�$����DK1�<�M>16��B�6DS_$b���Eώcێ�k�jB4pe�D�I�t�12�	�"#6�	�!��9O��۶�N��pD�po �F����T�T�ҝA�ԥOJ�nZh7��9KȈ�ٲeӕ	�T SI� ﾘ�t��f��6��*E�:h��|��r�$ÆkQ����0��Q�$��9��0U�%?� Q����*�$Tׄ���'5X�YąȊ>'�ŵ:��9���܁K5:9f�ɵv��(�h��dBͼk�
������oڈ<� �(�f,��d��P~����1a�rq(F��|�'BĠ��wi��`�`2��i�@�<[F��0��$3Fs�h2I>I��i����1D��z����A(v��L؈K�����ι��$��U����S7O8	 ��Ѯ�~�
�Bi��+��z}H��τ;��dM9x]���O>I�i����S���
t\�q��J9U@�Whl,ZǮ@/AN�R�'�� 9�׀�y�,E�8E}�(��3�攸�ѽ.��D�����$�æ�K�A6J��"❚y����[|}�7���27I�C �M�5mv�<�tK33��9ߓ7�N�'3�E�p)��j �̈,�\��#X�*4�	���dW�H�x�w�*����,9��{����N�l�93�,"�h8F~�ͳ,u�`߹i dCˁ<�M���5��]B6eP�U*�@b!Co�o�N~�\�eAD~/�o�I��'+TŃ�J�~?�MS�"����Ο�_d�0�au?Q��D7~T� G�7M#����![��0cG�v\P���k�D󗨏	��
IU����a�f�����tD�I>P�lE��I�,W|-b�N�#l$<+�� �j��v��jD�ɱvs� �Q�G�(�l�I��I��%EٓU�~]1!'�5p��1猎�Ҕ<[A�'\O�8�'2��S��X�O*��K<��y'��?12��P��9�'�d��1}R�&nv���e.\�p�@�ʞ�g	µA��f�'��M�	�YHRر�$Q�v(4���'���H$hU*#���`ɴ70r���^�V�0֤P�ēT��<O-��V.�~�@�`A��[s˔<�	�ܖ�y�_�u�M�ׇ� 1�l��P��y� ڶxu(Rs ʹ�y�E�"Ӏ�[��@�<����?1��%̾�`�ka0(�M���O��{e
Z+��t�LǹGW(�hr툛&���v5Od�;��"ߞ�9�R�(�u��D�����������͇d�XD%�1�az���s�b�=Gfh3M�j�	dG�,S&��3�PCy",�?5�>%�N�W[��r聦S��Z
����a��#?9pHN�R,������;JTm;��Z�:�1�*��B���xr�V���ѫ����hZ����OV�J�\����9��]A��埛�f"����j�dǐF����',Ta�&�+��5��g��I�����B��E	"�d^�=JRY��E�(�$���E#�,�5�\���C��?�d1��iN��Fz�M6mK(�A%I9Y3>�q"����D�r�v\JcD�V�v�ˢe�q(�c�E��)��gG��"J�a�G���p5)J�1�dy��I� �Ll�VÏ�k�ZP"�NV�}�8��	=외2�Rnd���O��Fx��'�z٭1,&A2�$j���E�B�<�E~2�l0K<��h�y!z�#D,�@:�%�����̙�Db 	��M2/>��<OtW������#�q b�s��Ɇ;6=;��*��N�|0:�h7A���3C��4״UwI�.`~<p�@"�q�X�sGK��PxB'�mp�H�X�
�����v;�,x� 
C<H�s�̈�M��ڢ�r��O*�XF�� �%�LZ,Qց 
�d�:�RM�0@->��a,�B��#��$]�Շ���YF�ӟ0�� ����J����8w�֨`g�Pu�aa���	.���D�?㘤�>q��!�Pd����7�СCCAl�<���&e��b�'y�����c�<!�H�C ���k��;��e�1�\�<��.�W�H02R��'ab8A��U�<��N� �lR)$,�P��@�P�<�'g�]E����C�o������S�<yD�&� +R��{7��a`��M�<��*�*N����R�G�C�� ���^F�<9�B>1� �S��U�X:�e��M�<��K\�4
r�{pl�-{Y(Y �"�@�<��	y����嘬�Xa�OH~�<)W�Ō[pby��@ը�R��c�~�<!��/�B`�a	!qB�\��@{�<��΀3!^!�7�MKܕM�o�<���Q�u)X(Qq�֖c$aJ4�B�<� 2�ѥ�g"����_���iH�"O<�{2K��m�\Xg`��Q�YD"O�ݑ��q1�$�R��j�r"O�Q�E�XFkvh�|��T��"OXR��}�x�:&��58�qBb"O����	0I��=;������3"O��#2)D�$�����cS3E[^LS�"O�����aDδ�VLO7GV���"O�Y��-�]���Z��K�N��)s5"O`s�A1L|v,�  D�i��"O>�c� �rAڼ�O�6�`�H�"ON��Go�,!����ڠ�Dt��"OP�Yn�/"^XP�v��W&�
u"O�-�!��	?3�4K�@ 'V��A"O���pß&L�����S���6"O��Vݜ?.4��DS*R�<	F"OtD�d�B�Z	���%��Hx��"O2���ێs~��[��7�H�8�"O�����I��G�Ѫq��"O����Ñ6A��#3�+,�H���"O z����E�Xx9&!����"O��H���(2���3��;"k`h "O�r"��Y<�DA��ށ-c��p�"OJ�k�eZ|����'ܽs��]z�"O%�T
 Gd�)6l 5y��C"O�D��K�	3 aXb�� �)�"O���҈Y�Ҽ���W�\�I�"O��Ȕ�� ��P�CI�nVU��"OXE��nR/WPb8��瑩i����"O��Y��X�F7��%�I�H���"O��E��ǾPB��:Ϡ��"O�`KGc�p�i���h朱�"Od��e�z�^�C�:�*�c"O��0%�>b�c�"��n��DB"O��CW�f����u[Z�F"ODxE��#����#-X�Mer��"O�32�P9l�<���WW�y��"O�	���H>n���K8X0��q"O`�#%��3͔���,]D
�k'"O�-rP���|��xq��<,(�@I`"OX����?�5iGѦ4�	�"O$�� �x��ɨf�Y�d ��k�"O�|��N�u�X�
A��v�buB�"O"���,V�.��L�bÆg��A�e"O�-;�N�8+�>p���T�A�&��0"O<uh%kE"&,z�а�
��P%"O�E��cx�8@�
GD�ŚvX�F{��Iوqh�Ydӝ��py��4j!��<2:.�K�n̪��$�uR!���D��B��:���$$jc!�D�*��V�h>KR��-Q:�O2���t4X�ܐ�@� B$�3H��O��D�U��`���M�A�P)�� !�d�6J�a�0b�MTt�����Aa~bZ�(H2(0S��)�h�����%D����;[���Y0x��i���%D��Z%eȹ	m�X��)����"�O��	%)����p���uB81� B�� �Y%
�s�z�I���&[`��E������xnj���/�u�)� �ޜMS!�d&c~����(}6��B�"_-f���Φ�Gx��	վ6��1i�瘯v���KB��S�ўd+'�"�m�Z�@@�4�б"�����X(&����I�nc�p����C��I���
�����dχ�~
� xug½>t��J&HH
o�z�QG"O�9��L�k����"�Pt*�"O8I5)ձpD|��$�!E|�\�@"O�A��l�n���゘atؙ���xb�)�S�v$JA"�lE��T(���˪u�\B�+�"Ը�-��5�2H�&쇨w��C�	�V���(��р%lcA�-�6B�I� �Ac�/��%� 
R0Fv26�5����A���@���V�V�c�-+��Q���O[���X _\����O2��*	�'}���g�L�S,�-]�h]0��D}"]�|���'3�D0r�00.�քE!'� X)�':��ĢFBvx��`�O�]��O"��S�M�	[|����j-i����p>u�U&�)9}*M57?V츦�-D�t�N<������n���7n?D�Cf�)6F���NQ�Rq��h`K D�̐�B��Q+��@�����0�O�O�C�I
�����D�|��q �-_'-����$�<���K�
�� ��Iƴ	6ܣ�l�M�<a�k#3�E��a�-P��<�E��I�<	�.ΝL���h�
�(S����D�<I��!a��dk� E�Z<��%�J�<i����T��jjr��u��{��Q��%w��g@XV��I �T�O_||��Z���P��МH{>Hᓉٜl��І�/�⑹��T��:%!�ŞK���>ы�����ߛs�2DĚ�n�P��0O�1�yB�#��L3�"X�T�p�'3�HOf���Ɖy
j��7��E����-�e�!�}?�x�Gه�Vl"G�ľF!���P��S)���	K#��X!�d��d݀���ۦP��\�D�*�!�N�	 	9q���}9ƅ�#gH��IV��H�ʽ�č2�2t�O�	��Y�TO$�R�s�R-�3K�;[ ����k?)�!��0O���eK��K�@�� %K�.�!�DB���1���B�v�*8D<�!�d^8�l��ɏA�H���T�!�d�P�4m�N�u��I)$�
:�!�d�?I�|�s!�H	\�PA@ $4!�d����D�0L�.4�q�ȣ*-!�dG�Nk�a�Fg�a��� �!Q�_!�I���>����F�r}30�[8M�`�G�F�<���P+��D��BƵX*�d�88�!�rZT���;q����'	�d�qO�����L���Q@�� �2���}�!�dU�A���C���2$@U9�cZ��!�d�3�p��D�
%�q���X"Ce�O��=%>��%K'xV�]��^Oj���>�	����pEEV�+�z�C���~l���G�6�F�P�&7X��W��c���ȓs�0�b@�
up���c�~+ʘ�ȓ��I��oR�>Y�EieK�8��	�ȓK]v�Cg�&Q�>���'�Tt��B��З�S	&���mص~�xD|�w�"���l�9�$��@�<�B䉂h	���?3+��b�-^�B�I!ad���S(i���Nް:X�6�'� �M�W�����;=����)}��'�f k��מh�Y�2ꍖ	�I��'��t4G�;r�p�L��6i�� �S��?Y�
]tD�Wf�H���v��J�<1`P	?ZYHrb��K��9�dI�<� ��kei��v�28)�@f�>`	�^�dF{���S�b��A��Ƅ[Ҭ ��G$z2!�dҼ#�(H�e����i7��:/!򤕸W��L���WR�!�`�ϱ!�ԥ(�2�����~��Q��뙆'!�M� |*�&y��yf�$t�!��ߙb��a�eNi����@;g�!�D�[(P8��~�r����]�!�Đ�(�c4-MŦA�3NH<!�d֓p< �	T�ͪ��ؕ#͕*!�D���Ds��~�T|��"%!�X����A&Ƙ2(c�A�/?]!�$�e_�]�4c���8Xsq�^H��M29�� ��*q�+Ȃ�y"�S�C\`j鄞B��V����>��4��$�bej�i7gq��A�T!�$Фze:�QA
�Ҭ3!9hM!�­&:�� �� `�24��[74<!��յ.S`�$��ɛ��<q�O`�=�����wm�99^
y�2�F�h� "O|�Puf��|��y�q��?��V"O�!dBf���B4�YE�`���1����0�����G�c�V=�ԣ�(9($B�	��&��g���>S,i�uC� !1XB�	�_�xH��\7q92ȱq(�1��B�	=hi$Xb�G�c�0P��"��"b�ȱ�����3�0
u��}�~mK��O`�=�O|���t��e��}�)p(�P+`�)��<A4�N15�$��hD�L4C�A�<��:��=��I��67�m '�Vp���*���\-��Ε�ܬ���A��<��M�hpP�ֺ9���gNׅ��`�ȓ1�Ը��
A�N4�4��L�!�.�O���dW�
���/�����L
!��>D�J���@��!P�h#�Ya!�d�K<,ѻ�T���X���9]�!���
Kܐ�Z�e�8*�RԆ���!��@s���de�8ä萓E�!�DB�&������\}��%��L�!��
/
�=�q�N:�^L���Ud!���~d6(��K]0>���U�,F'�y���d�0���Z����!5���)�~p���	��p<��#�%^^\��g!Ʒ+�������G�	�YW���?����v���C��TȚ��q+i�ARU���y�
�8�`��H)Bh���C��y� [�E6��v�^�(Ǿ ���^��y�dDZ�Ը�Ø1l��a$�$��'�a{�N��4��&ô\l�c��'�y���c�x��	F
�8b�F���yr��fz�<�$�7���еA���'��{R�N�F,D�	�J�(��X#�	�y��;>�������&�������y��V�5&�Be�E����cѹ�y���9F����!N��C'�B� D��y�
�%1:��p����*|��a�T�y���?b���a��YV�r�+F�y���"���'�´<�\�q����ybbF�4��	B�mB=*��Y�1�@��y"$Ž�2����/��e��G��y"%	m�Pr�h���ݙr���yb�#o�R�q�d�6�����J�.�y�Ө9g*m����70@�*!��7�y�kݥ$¸D�d)|�
�mR"�y2�ӛ{*V��5���f�(�@�y
� ,A���
����[��ʠ�G"O��ɴEE�B2��bA���0��"O�q<?�a��	ӹN� �1"O�}�F�j��mY$(�;MHڴF"O��v-=<��U�g��6<�e�#"O�ܘ��F�Y���&Ǟq;L��"Od9h2�\!9�­hp��6PR�mX�"O�Ll�/_6��R�EF�u��"O���a���K�;!��D�[�"OX�12a�8M�H	wN�-2>�d�$"O��QD�
I�R ���. d@�"O@����#g�a�_�-"Ol�"��+GV��+!�C�f�ɹ3"Oa#�%�v( �UiE�H�(�JT"O��(w��4�\ѡ���XZPq��"OX!G�ֱ	����Fb�jG���"Ol�҈�q��Eb�A�a36\+"Oޅjt�Q��n� ӎx��T��"O�`��)P=D��@�"ٞ$�A"O
��#��>?�*+#$-�
�Qr"Oڌ(�N��j�!�δ��"O(�ӂ�^�{��s�H@&�T���"O�9�7E0}��=�UG� *�0k�"Or���.P�#��&�d�<!r&"O��#���#t�)1��C��"Ods�G��|�zM9wT�^D ��g"OxX*"�˓њ�`��7�x�"ORXbV���:� ��i�dr�"O�myp�Z�HV��#(CK{dYpA"O�K��p���2eT�Aآ"Ot����O\���4�]
dJ��*b"O�D��CO�qd��[Gj�;5"�4"O�p:p�ީS��D�&D��h�"Oȼ�� U�"��}pq���N��"Oh���lS�j�$us2�_�Z��"Q"O�i+��x�<�K��^>=�Hs�"O��Rq#ǭb����R�^�҄#1"O0�� �Y_�8UJ�l�7�0�c"O��y��Ƥ]����j�8��ٛ�"O�!�.ŀ|�g�
F44�0"Op����P�x��ͲIš%,t��%"ONP����^�@0�� $J���C"OzA �|� ��F��f2^�x�"ON�yaV���$A�f�7&�ii�"O����	�k1�|�3GV���I��"O��!����w<���f��*C��"O.�#��GW��e8��P2[,�t+t"O�)�@Μ�H�cʫɾT��"O$�Z�oC�Ln��!aȻ@��� P"O4Аta����� A�N��i��D$D�$��,�<��e���
�<L����/D�Lȧ�]�ϊM�G	S=_F��#�A(D�A0B��
�@�o�~ ���u�)D��Za,��7ؘ��aa��6���%D�P�Sb�f���-�;N*��7M(D�D#G��o�l�K�a!�a2�j$D�h����!�,,��ډ1 ��a��-D�Rqn;��JG�S.���2!D��Ӏ�8"-!��<V}R1��?D��r�B<�L���d�w�I�C:D���B@W�p�V�%]E@ ��7D��{��f}��T#�>�D�*�!5D��H0�$�@dbD�N��)h=D�)A�5�ȓ$DB�D�}K�:D�� ��cG�C<4غ�&���`��s"OXhP��Ǎ]��d�æm1r}Q!"O�H�&��t9�|��n�/1,!b�"O�9�F�ܡ �`ec��Ƈw�u��"O�L��DK𰩳q"�&6����"O�<y�'ՄM��iR���Ce�0�"O:��Չ|}��ScN��Wh@�4"O�@��%>�ul�?hJ��"O�8���>Z7�u��ue�m2�"O^Mp���Y���V��(e\z"O�x;���,Ϫ񊂩� T&}�6"O���,F
~(&b2�N3�$�%"O\u��O�<e��%HBʖ�Z�"O
�r�*�5b�
q2r�(�X��"O����B��#'�׋	!|��"O��{CM-]ґKf�\+�Y��"O��st�ȇ&��8���H�F�nM
"O�-��21L��vG��g"O���	]�B<P)J��:wd"�R"O\�3�� H��hb�<V�d��0"O(�5lתs��+EFN,"�"O���FD�5#ǂA�g�|�`1b�"OT#ng�ڕ�p)K��tP��"O���H�Zl�Q
L�oi>8�e"OP��RE��B��f�1]�\h��"Ot�U�>b���0vDQ�Cl��q5"O�YR���1sPl̙�OIf^\J�"O���m�Y6����X>t��"O���d�J�_�~ut���RB���"O� �F�*4 ZyR��B��F���"OʱP�,�sl�ّCh��1�8�z�"O:�Ȧ�9J�� K���a��a�"O���$��q��V�<�X��h�z�<y&�*f2hס�Q��U�s@ y�<A�,�q=:����� �v�Q� �x�<	4@M�12` Nɒg5�`A���u�<�f�S�H���4)�%WM�4�רDt�<��_�8ayĨ�d�� ��p�<	ԦU8��dE>4�T+VF�T�<�s��!�>��w��:+	>Բ�U�<	6扫dp�pҡ}�zp�'�L�<q��3�@�g	S/KF1�u!�H�<9eʕ�t�&阀�J�j�d! D�<9��'3��Z�L�"\�id�t�<� ^C��7��%l�<%��n{�<�&B,')dX��ջ,�$�r�}�<��A	!�b}���س���҂�[z�<�Ԣ��E0e˥�J�I�P��t�<a͕ )9:(z��ЇE��z�HSk�<yغl`��Z3��i�^�VKTl�<y��ݡ#�*Y�F%��9Ѥ��d\f�<1�E�т�i�N`���� Df�<y@Ζ Zm*��5�E*P=�H�c�<�c
ŏF����}��@*��L]�<Y�d�g8a1�Jw��y��Xr�<�V��� �^1�2o��%�#r��q�<Qq�@�\�0l�T	�VdH]kd�^q�<ѦBQB���`�˔��,�Z��F�<	 �G�F�l��R���1㒘"�h
}�<�1'�F¹��]y ����w�<1���- �L�5�Q�FxZ�QO�~�<qK+Q����E"�	��M����z�<!�]+�����j�IT%Kv�<!���l#�ɓ��B%O㚥8�(>D�� J ����7h&�!`���J���p"OXC�h��H+Wf�
u�x�%"O����P3�,H	c̻Ob(���"O^ �Q�֧A�*��R#LJ֥��"O8�
uI�z� �Y�Q�mI⨋�"Of���)Ҩ�����Ji6�:5"O���c�H�t�$�ɓ�[)y�
��W"O��3�	I�L\v�� "��:�z�IR"O��(�ə�F)����1&\pq�"O:��EL�/�,��U쁩_^�+E"O���Ӆ�� �P�I#Nl[��a�"O�EB�b�+��y����(�lz
�'�嘐���8e��0a�B�P�<	���!Z`�)�G ?!��Q�N@C�<9��ϙ0:^��h�h:����Fx�<!���A����u��&�ه�v�<�����NX�S`*S��}��,�g�<�W�^�D��X�@�F,v�ܹ��f�<����&5[d��΀%zv�5��H`�<9'��F[���u��+#^�y�t�DF�<1�aVy�n���MY�u�Jt��mX�<����WP>�K�=�8a4�BV�<�3��0n�9 3i���d�hT+�m�<Q����;$��rD)��DK�a���q�<�@FŎZ���CD*ϖM�n�{���i�<a�h_!,����t͋�M�Ɛ��i�<y@�ѣm��A�Ĺ{�� ���{�<�&
J/V��|��dȚ��uP�#z�<�)X9>����&�O�?�༛�F�t�<�ds�&�÷j��br�}Cň�I�<�s���cX��˄'q� ��#�D�<�h�2� �qLՉ;LX,���}�<�r+�C\&ya���㶩�4N�|�<��ʉ&6&�� ߘ\�ڡz��Fw�<���=C�8c�k^�{T�#�v�<YC�R�	v��C��$N���b,[o�<Y�O�H�^d��샅Qِ!��WU�<��m��uM9x�Ia�f�T�<��/n�z�f��2"���8�h�d�<��$R�~]h��QI�����l�<A�	�x�ΰ�c�iJ�ЧKk�<��"��
op�ӂ�J����i�d�<IÓ��e�RM�I���wCd�<��B�T��ݡ�
�V�tU�bh�E�<�u��0aj�q0�V5PBq� ^v�<QD��a�x��%*�������q�<YU)�>W{t�f ʈ䣴*5D�\Ȕ�5T�j�R��7Cj4�a3D�<ؓ�L���w�y!.?2�u��'�d`�Td�6>���EɌE,�EZ�'���𴯆�jR.��gŖ�)ctP��'o�H�T�C?V��\�s�J� �a:�'DE*��/K(��/ׅ!p9��'Q�ͫ�*�+�xMB�����
�'z�piv�G�)n�h�}���;�'܁I���?a���戙{O����'H&�Ӷ .yP0�&AV�D���8�'��P����yتub��I)Ia.���'@��Ze�
--52�irm��Xq�'�Dp�G��b���Y�O[�$��'��(b�Y>%�w��)p95��'2fQS혔 ;� ��1^�j�	�'ǈ��T�_4Nrn�� [']$����'U���A�2�2tP�oZΰ�Q��� l�sF�;bp3 %P(��@P"O��!3J�.+< �Ve�5 �8=Js"Or���%
�,{ʜq����<��"O�1�R�(S��@ʄb�-��C"O�șc�H�ql$�JE2�N�d"OVA��2:�	RDb���R�x"Of]��d�P��bB�Z� �	�"O�[6�ٔI�`��CQ?1�}k�"OP̉�e��	S
(!&�
�k�P���"OX���([%��ɠm�5/����"O.<�׬�$K�%��KG��4ys"O����^��R݊�����1�"Oj�*]�y�L(��C� m�DS"O���A ֎��It��.ZY��"O���W�͠R	
8jT(L1wP��U"O$5��ިH3@-d�'U�X"O0��q'FN�LxB�S� @`"O�\K'!������3���D�(�1G"Ou�	��$�&y�UeW0�,4�0"O�Tk �[8a���ϚL� ��W"O�%�̘>9���P4�\b�^d�"OJdq��?)� 	��C��X�a�"Oh�ۡ�Ұ59���;�x���"O6���
���-QY#˞c_X@��"O6 cEM-i>H�Jo}
}:@"O��SkA zf��7��Vwh@J�"O�d[ g� jQ!��'�9v�t���"On �s� �o�`���#ݨt�S"O����Ѻ,rԁ0L�l����"O�	+Y�z�>d#��� R�C�"O�넨��C/��y��T6�L("O���B�4x��ͺ�g�R�TX�"O�@1�Ɠ:�PQ�v&ތAX��0"O����%j����e�f|��"O���lY�A�4�$��Y�> �!"O����,�6�A!�"G�K|�g"OF�"�Ie^uX�D84RI{p"Od@���,���!1/@
f�\�y�"O���t$�6D>��Ϝ*���"Oh���.�#/�u��lF����"O~T�1�� ]J��Ó���"c&�i�"O>PRԊӎ�n a�;9�ds�"O���E)B���1�G@A�m�T�s"O�y���2m��ł���p��D"O�Aa�T�]K�xDN�q�y��"OT�R'/�!u"6�`��� �[�"O�k��A\g�@��%V6q����"O�Ak5��7)cv��D٬�:h0"O�!a1�
\3�B�)���"O��l��C8�����Z��!�p"OLFƙ�1|�)��ɒ	K�=I�"O"]��.�M���B�P1�X��"O�lRg�8
n�l��.�Y=~T
E"O�T�0L.XSJ�:��I���*�"Ol����ј ��\Bb�*l��5��"O2� ��p�P�"����Ѕ�"O6�XN˼�(�fJA�F�~)��"O��F	ҐdGx�f��Z���(g"Ox J��Ջl].}P�G]��H�Q�"O�)��mJ�|���冔+5�|}!�"OP� eA$�<#4&�"°�Q�"Ol�u+�e|� %-M�LD��"O�гOJ�PH�u�QǈR�����"O6б N�}
���� ��y�c"O� Q��'�6�`�� �k��@(�"O��1��IFp���0L|��p�"O�"q��dXp꒓z�ݨ�"Oa�$�]�QXb���J�)p�у�"OD�{�ɚ��)��Ǜ�*X���"O�S�:_�u�S�ڪL$�s�"OB2��>��b��X�N6y��"O,�ۥ\�okh�ц��7_� Y��"OpL�f���%Lʱ�u#՛�\tS"O )`�(�2P�6Q�v�%y��2#"O�U�U�ظqA %�� ��P�"OH�P4�a�����l[�?��h�"Oz����/b�Z�Q���.Y�m �"OhlpW���l��rpJ�B�
�z�"O��F��E��ЉS���@"O dP�
�m�FAc ��M�>��r"O���KŐw<@���ȍ@�ҥ"O��f�W#	�'̏yb╳�"O��˂�z�*Iv��#-��e�B"O��#E#V�S��ە�C���c"OJHsdFY?yǆa���49�V�R�"O�1�K֬,��]���B��B�"O�S��I�<�\*c�Ț ���"O�  4�EQ,e&H�s�m*3"O��#!��5��0@m���ZG"O4}K�i��,�XrM� ���"O�Q�'NĮ�R�q�ȓH  1�"O�)��G(. Xq�!u)��"Oڈ7�܊-���R�
��
��Ȁ�"Oą���<q��Sj�z�bh��"O�Pz�I./��ԛ�ɇ&k�,� "OlU�E��h ԪP1*#:e�"OTq����YE��i�C�l��"O�<�����,�^艕�M�qX"]I�"O��S�XL�h���*V�""Ot5y�m�w<� sfX�	Qxq�"O��s&j\�%�r�� =R�
"O����#2y���& J���
�"O��"r��
�V����+ �� �"O��.GB�)df�&���"OX��q%9+p �;r
�qK@�"O����E�tQ���T�x��"O���	/�p� ��=~%ʉb�"O-�Ǌ0j�`93CN�r(�"O\]q�I�< ,l9R=4g���"O���Ԣ0]��lٲ(Z��n���"OB��lI��(!5
B�l���C"O��JF)ҕ-�<����� ��	��"Opݫ���!�:�q��R<!q�%�u"O���PC�,'
��4��7m�1٢"O�U����.צuPo��~��c�"O���!�Դ��DߥZ�!�"O$�'N�)7�<=�'MQ�:��I�"O:<+B���l�B��aB�f�tQ�"Oଓ%��;	�fAPp�!K;:M�"Ov�J���L�h���57!̵0"O�-X�#�xE�I{��I��4J"O�)��)�X���+�^~���q"O�D�f��&���ˆ�Q��xG"O�ԫE��[ ~�z�@�Q���0�"O�t�enE�A}B,�vo�#��ԳT"Ol��B�	�ёKG�n����"O�I:r	��&���R��`A�B"O5����6���A��C �2[F"O� ��&��1z${��;[��"ORP�#��3�֔���&�r�Z�"O҄�կ��\)^��v��4Lꥈ$"O��JeŒ�.�����L���6�a"O���w柋k�F�ؗJ��rs��0�"O<}��D�:���a��;#`�T��"Oh�I��8nҨ� ��:V��Z""O����E"Q�{b�ԯ|�����"ODd�r�C��z�qƍ+�h��"O��6&�j���e�8���R"O>��1nV�C}��"E}�\Y��"O��ӄ�2���vɇ9�%9�"O~��+س/~n��k�y����&"O�!3i/�2e(*ݺkѴٷ"O��;��-eߜ��	N/�69�"O���#���uz
�qqɕ�/��l2�"O� ��@?/T��`�Iڄ`�����"OzY�J��f�h���A�!:����"O6|���mj��q�����2"O�Kw��5R���y��wyP�j&"ODD�uC�-�l���)��&DB �"O�e�g/��i��h�HV�$�&"OT���*5Pp��C�G�Q!�u�"OtH�a��w�f�
s�X�Wr`S"O`,h�@2U��1!��]	f��"O� ���>b��[s�?���P"OdH!Ŝ�l|�k��6� ��7"O��#�H)'6\�@$�S�w�q)q"O��x�Ǆ�v�&�YF�>r^��"O�)B���L�ceᚽS��"O�@种*$HjLH����X�1"O�,;�F�*p�Z�-��1ÔI�"O`��p��:|2 �MǢ	�@�c�"OQ��dA�<f�jэ [�.d;3"Ot�pAĢrѤT�0*�A|�y�@"O.B���B�T$)�'_d!� "OX��g�ȑw��4�eeO=Hb�I�"O��C���N�>�Y񃁕V�"���"Or����nK�%Z��7z�<y+P"O��>���D��2�r��"OD�r5��l��8@bT-"*YbV"O�EP'F�i.z��d�d �U"O�0Q4�R6n�ة�d�Ol�j��"O��Ë����#��"?~���"O��e׌&R�X�!ի@-N5�R"O��s	��37Ji��ώ�� #�"O�x�[�xS�UZ�Oو7.���"O��X�*
�z�a�P�̰YM,��S"OB�Ah�i�(lQ�΂%�X��"Oބ��'W�O�zLZ�gĈ?n�6"OԠ'��sc~X�GG&Fd�x�"O4)��Ųw��Ps눋#%�ժ`"OJ���Q(Q�|a�	�>2t�Sd�<���-*y*0:��Z�`1���f/G]�<��m0GiБ��cc�N����M�<taH�O��ЇtF��0�H�<��G�[����ǂ��ћSLy�<qf,�-�֝ʒ�ݤ��ѯQv�<�d�Q�&�	#�"nm��(t�o�<�ЄP���㴉	�/��Hw Cq�<q�m��:�r���� p�����ΊV�<��Ɯ, DB0��,
9:�Čٳ�PP�<�v�ߍ�,t �@�Nr�m�fO�<!bM߯|�j�p�'N�3��24�M�<�  (���\�����)�-�fQñ"O�9��`"\~�0�P	� �P�p"O^��7	�-Ő��a�6)Ӂ"OƁq���!6в#bOQ�E""O��ă��z�1�N�7���""OR�����X��c��
:L��	��"O��{��#����U�ά5����"O��X66���"7M� hR 
�"O^�
�Z1f�8=��K��4��8"O0BN��=�\ {�+��1�m��"O����ˬw�b�ӂ��,�D�Q"O^���&L�"�L���ԖP��"O�ef�!���ŉ�{^Q��"O��E_,l�6�C(���A"O&ի�W ���$zFH{�"O�u`�f�n��g���{p<��"O�X� ���s��r4 ���Pq�"Oj=Ђ�<�qѢ�:�`��"O6��'�P�>�)�LC����""O� R)�#��m���3V~("O�=; �5	����b��-����"O���e��"���!��B)
���"O�}@�MO�-�` $�ޱ{+��*�"O��b�E�k8�0j�	ٽ�:<��"Or� dkY�Ca���c��%E"O,����2)�y𦕸}�<\�6"Oz-�a@�W�l�aѥ_�xM�D"O D��ɓ�B{.������@�;0"O���(�9����4��1P��9��"OVq��n^1(Պ�"�9B�����"O���aB�$yX�������"O
$;�������8R�H�C���"O�񀟺:V������5"O,i��a65���*t����z"O�E8#T(]�>�k�F+@���d"O
9V���d�L8��nL�U��(�"OQ�Ʌ�J�OH֎��"O,��5����S�B��3�"O���j�'!�lMZ� �Hr"O�-�q��4�����)�<wj,��"O� c��7gY�����l[��Z�"O��2ɎºI�ZitA)e�I@�<�q�I0=\L���
R(�Fm|�<�#�1tb5{`S�zJ�T逪�n�<�c��U�61
"��+U!Q��B�<�� (��1��"c�PDFA�<)�I�qH�E����c0X)~�<!uLB�yN6l�*�t�i���r�<���ѿ35�Q�u�Y�4�r��v�t�<G�,-���w��R��!���n�<�0��2Y���Y��r�hвf�[_�<q��O��b�Θ y�сA�\�<��g۞=��0�f�ŦCv����\�<a�E��z+��*�	�P1�хRZ�<���-<ęE���tp�@�/�R�<�W�7{Θ��ς�5z<����L�<�d�ӺJpX���5c�L�9��@�<��
�t���-F�0�Ո�Ty�<Af!8���ٴ��按���M�<�1o�
k�x��k��m�`�B�@�<1@덷@�B�����%ݩ��F�<Y�ʆ�B��l��aG""��)���j�<�jڣ�53쌞	�L��!�d�<) �K�9�%8ѩZO�^�*� Mb�<� �dч$į?���2�#��\� �i!"O���w�J��ld��V��r�"O���h	%��ƀ�X����"Oĕ�0�ҋ.F�KF�?c.��"O��B� Y�r$�a�T�L`�#�"O,���G�I$Q���f5zY�"O�0�a�-9��t���0HL ��"Oh��ũV�BW���@F;0��i;�"O�<���	V��ѱbONu����0"O�-�ׄB�*BDi��LUL )U"O���d��6��[w�98�H�"O��v@�=
�Z�[{İ8�"OTMA�g�bg�1!���\�&"O�-`�,2V�0�U\?D*){�"O09ag+@�IX5�N2#��d�"O�4�gZ$1(�H%K�\m�ip"O����A!R�\EjҀ$?�� e"OlҲ�H?E����i�:?N`ݛd"Oq��>qa��*���6�"O:����UHwB���
\�p�`"Oސ�a���DG�?�~d�0"O� �¬H)0Y*�N�����t"O�\�߈ �0	ҍ�d�<�"O�,!*ҙT_8T�p'�!
��Y	"OHe�%ǖ�=�H)�gR:Q�ք�G"O�p��$��H�B�%\�m����"O�$�3��BѪ���*>q>�8f"O�p�^e���ATĜ�B^���Q[�<)��Q�P����GG�7g��
�MX�<1���66�@��(r���@�P�<AS�է!Z,��C&l���cAF�<���R@&/�� �U��F�<�E*O5;��Y�Q♻LM  jUFg�<����'sLέ�C5�z��#Ue�<�*G,>䜼`��P@���G
�c�<��ů�	�-��[n�H#���a�<�c��5H�2Q@	ۉm�:�q�C�<�6��'�~X�Ef�E�����Vi�<aH�)A��q��@��sĠd�<y�-;޲-���I�*(�����N]�<q��Hz?������tbzi�U�EX�<AшKq6�I���ԙu*�e��S�<��D�/>��� �SZ�B5�AD�<�R�j#V�תT�\4쬨IZ|�<A���Q>F���j��D�RŐu�<A`�ȭ���C���o[vC�G� ��Q�Ϥ^)@�	���v,��ҥ+��2�oݵ+�P� GD�UE!򤚄a>Z�Y��T�Jfm��LE�1?!��é"��MYg&pe�YC�+!�!���A{�E�'�<BT�h��JU=f!��׀(�|9����E��A�МT�!��ݟb���,]3h;�{��?r�!�DF?�J��Pk2���fYw�!�$5ݶ�ѷ��|)H�)r��!���=����Z4%�군�iˢYe!�Ɩ$g
X�.rI8�X��ŃS�!�D²n=����̇NK&���'ŏg�!��4q,5ze�N�E-�P��ŏy!�d�(����-+ȶ�ه%�!!�� .ͤ=`f��)d������!�$��dk�8�"���!��<t�X�<!�W
��:Ei�&<��C�L�!��GB�(U��!D!;�J=Y#�S�!�� �c�l�w�Kp�X�`��d��"Ob(h�(���μA@g��Sn��$"O,��u.�$�r�t��{N��9�"Ofݢ���0!�\$
0#�mGl�"O�����L�7�
���bT{D��Y�"O�����p^aA8?�$:6"On��慂3J�hug�59܉@G"O|	;��Z�6�V��F��l/x��"O4U�P�L�XH s���.\-��"O�`D��X�"��dJ�0���P�"Ob���.G�X�`�G��k�J��""O ��e�!Y�RWF�eQL��!"O���P�O�<��e��6Y�8�V"O��� R8G������qm��"O���gw����36���"O���H66����N�=�(�T"O ᗮ
4$�k�nS:$ش"Ob��F� d��e���7�EP�"O���e!R�p
�pr�a2	v<w"O�@:��օJ<�iAP-o�r�0�"OF,�Q���~Ш���"9�j�3"O���c��2��!ȵ�
W^`�U"O�|(�����S摙Yubq�c"O�\�RD�D���e����D�2"OX�����T!�X)$"O.����F"O�9�D�V e7�qK��Z/N�"i�"O��;���L\����ܪ��T"O8�d�6tQ��	��R�D��y"O��3ƃ�
U1"��-��G�,��R"OF]"�ŵ�8��f��t0 �"O�a���V�*(f����3n��x�d"OU
 �/X�.l�&`�E��8j5"Ov����R95�9�gDhɸF"O�|��"�f�p���
�9�xi�E"O��IsG�V�mQ��(��8��"O\�Z�L�3���+�i�ֽ��"O"�;e恢m�I��d� Rrt�kp"O8d{�ŗ:xd��j'��i�ZQ"O��`Q֜q�fMjpC�,7<E"7"OP ����,Q�,��r�׏H"��p�"OJ(��h�;=tP��#��&A&��"O� ����'{� �!��Rx�J�"Ov�jS�-8�<y�b̘�*`� "O\����8
$�����=x*2��"O�ջ G�F�"�3�-��fI��B�"Oy�FG>*F���x6��J "O��%#�L��u��,ܜj, W"O���s
�I���z�֟ $d��"OF��uH��ND�@$�D7*�ȭ�4"O2̘S���=cV�AծH�\���"O��A�JÅ7'6l�%�L␨[�"O�A`�V� �c7-��L���"O��SҡR����y�*���	q"Oh�ʄ��?Pp �Ѷ$\G���3"O��d�)|A��̑'�L�*O���2�@�5�	#:M��'T�5`A�˜w�ҕH�L";	t���'��DCt`­���&��88a.���'耋�C��O�-���(עM��'��7+3-�ġ�3N(Һ���',�$�h��c{�)3.��QT|c�'w!��)!:�h#êB4QL��j�'5��c��4{#Z<0�-V�6e����'.=)�J%nL��R ���'RA��� �槂�?I�Ű!/P�?T=��"Op��cY�|7��*��P"w3ݢ"O��qPw��${�L��2@�Q�"O�;0��Fޔ����?�-¦"O`pS7+V��q@eI��l��%"OBE[ n�=.�
�H�H�97��%@0"O�d�D�E�m�$���ƛ�k`�%��"O�@@2��V� T��Gl�x�"OꠊV��5ߎ�{GLW0c�L嚰"OJ�X�&^��~�
!l��K��Q[4"O YpAM[jr>Q�v(Ix�"O^Y1���6t9�P蚫L�9�"Orp���b��P��$
* ~||��"O�ac�GT=O�9�R�?5�~y��"O�&�Q�$I�AJ�c�J��"OR����O�@֨�b$���S�z�B1"OF� �����"��L�G/�V �yB�M�s�t�)c�	�m͌к�.)�y�GWI�$"��ix�e���y��1w����CYs��	q�F
�yB�F�*��]���[�v$APb���y"�(��+3@J�_M����9�y�a�!USBAE3o�HX8�$��yb���F�h�aX�V(�&�yRl�0��t#ւ)oR\T�Վ�y2A�!#1���RF��b���X��yB��9~�z�R��-a�L�U�T/�y��L@�e�Ŗ,W���i���<�yҧCc0������vkO.ZW�Մȓ!���Z�X �>XsCĖ�H2���qd\��%�Aj�P��й}�d8�ȓ5�`[�"V�D�倊�;`�Ɇȓ8�2��@+�dݱ�a۳LD�P�ȓ�|��q�F^�(�a�)u�|��4	,�V�'��x�CV�n;�m�ȓ2ࠥK��(��x`��m��,��D�� �E�<Rw���LE8�VM�ȓ+���V�?(QR�H�[܂�����q���]���C��3G޸��oq��A7�O"l�T�14H�(M&�ȓk�
q�̋9>	P��,�����k�hm*�ɔ�l���dZ8X��0��:��E{D�Q�	���G�o�d]��DOd��o�85U^�(c.�lì,��y<"\ЇlIX�U�&�Xz^4���[
���ɋ�Cz��#�B�>�0��ZY����Z�ylD}@P�V<.���ȓu,30��?##$90�b�@�Նȓp�BA���NM$��4らy���ȓm��(���$^$)��-?b��NB��:qh�6?Gr��Iǂs�͆ȓWm���AK��)	�H"%�Y�;s�|�ȓr���	��Y��+�͸�p]���f!�C�OL��fH7L�<B�	��Pq7I� B��-�	�!�d»]@��L�AxZH�a��i�!�d�9j�C3��;gv�#�B��js!�dB�S*VT
�.S�(Bnh!� �:y�!�D?������R,>@�w�9�!�DP�SA�(9�+�2D\r��P.(�!�$_+�0����!<t���jU.�!�Do���R���'�<�C%�@�F!�c\�8R���⡁�)�7b!��5ut#J?$��\�qi��7�!�� �"�D��]���A,�l���
�"O��H2�E5O7Rx�hW�o�h8P�"OR�"�ʒN0�D`�f���|!{"O�!�-Ϝ^&S�G�3M�2TIR"OĂS��&*�Y�2��8�J�j�"O"Y1�e �`��F��gy�p�5"OJ���J8�:��H�z�t`�w"O�(���]�=���
<Z�x1�Q"OF��Í�U�0z��3@ag"O�1�t�\�D����d������S"O���e�1C�UY�}��@"O��3�f�����A@~5X�"O��pc�Q�V��3NS�T<��"O�s���$S ��A�3u)̬z3"O�X"� b.$Ł�ʓ�t�3�"O��9�BA3*�䉑 �BLU�"O"M!q�G�_�ը����%��8�y��ߔy�2�����4�������y��>�d@� ���b��a�P��y2-�*���z�L��i�&%a�#���y���	!.�#�ւ9�����J��y�Lb�
�[���]m����o"�y"L_/:Ь�T#��O���`-��yR-�,w��t"`o�E��Uy�cW>�y`�?|��Kp�ש	B̀!*�:�y�HF�&�
�X@l�"Z��0�H��yX��m;ӌc�6Ȑ���<�y���)A���r��]CB9k��D��y�E�|��PiV�f��钣ئ�y�J�b�����cߵe! $@P
R��y�(`l��O[8Fz���!��yB#�1�(�G��i�G���y� �n�Y��p��@�G�B�I�)� 82�H�N��U��"��B�|q~,�3��-.MP��C�c��B�ɄA~|�p�^#1������r�B�ɉyHp	fi
����ʝ���B�;� d�FL��!%N�x��B�9�p�w��0:R��G���nB��b����U#�T���N�*C�I���X)�f�&B�l!�Ѓ�f�B�ɠ�d��%�!`�r*Foƥ��B�I��
�*��F���H�ԣ��i��B�I35Qx�C�D8{�bl�g.�:=�bB�	�3��	�N��J+�@��'��-X^B��1$fRlX��C(d$��WQ�C�I�L�r��T�D�B�;Gꀞ)�,B�I�_����;m�xe���/]��C�	���Q:魌2Q�;'��B�	�M�r��V���D �5c���'rS�B�I�C6- ��7'։0�ےQ��B��*j,<���
S��­S	�	��B��0b�lu����`?r�Bi��R1�B�	�R���Zw��`�D�ܺg��B�I�1heRu�@#p��}2���w�`B�	�tPN]��n�o݀�7�[�6'.B�I�`H���ܐR�J	� ��<��B��RL~�%�]�
�d�H&�3+�B�I�E,0�6@ �K��U��sJC�	φ��r��%�Z�� �ZzVB�ɧ'Z��D)߱6�(UX$̗8\�B��&�v�k���Om$-`�kU�1��C�	C��@�� &-Ak�)�(�VB䉕�� �m�c��<���E�<;&B�)� �	��m�w�d@p�_�O�h@��"O�K��! ��P�g���� 3�"O��*�A`�VH�q#Y�c����"O� ��M��x��Z�~�"OΉ������C�-T@��"OIJ�M�_m��Fkޔ��A�"O:)4)\�vu^xy�*1
�5��"O�YR� QW֩h�F��f�ҕ�Q"O��0�,<IV�p!EIv@���"O��	%�^a:,���Z"�Ua�"OH�#aNXoI� W�W�X��;U"O|@�_��Z�E�2s9�УB"O��T �X�0M�r�+��Su"O8�2��^7U�#���1Ѷ"O`IbQbT*�(�`�[���d"O���"R>x�8zu@�%y{l�S!"O�tr`@�X�6X����<nw��q"O�ȋ2�79�0���k��?[���"Of��n�i���,ZM��y"O~�B�O�nJ�U�X,b֦��"O6�
���K+�Xs��:��H	"OlTF�(���r�"��w��4�"O0D��DH��|EHs/�	f8�!��"O�*�K\ D8�T��85xж"OV�	KG�tː�d�#\-"��a"O��@Q��d8�q9�e�+�yr���P��N�e��|�S���y��B�=깱vȈ
r�0E��j���y2��: `y�4-D�m@��"���y�o�Ry:��
&N:��1e-�yb'� "}���N�<Ab���� �y���u���Q�"T�o~e�@���y¥A�U(꘻e$X431dSG��+�yr	�B��b�*b����/�yҌ"L����'�Ţ'�H��7��5�y2-�5e|�	ʲ成$xu�f�D��y��ànQ����t�:)Ȗ��9�y�a��;j��f�6Y��A2�iZ��y�Ú�I��9 5�;x�X9����y����jl�z��������PK��y2���aIjtsхP�%ʰ�Ê�yRΙ)(¸���+ś�\Ѣ�Z�y2�L�.�v�ī\�������y�耵bbZ����޶o z�h��]��y��G�i��l���S\x$
����yr�ҏH�|;���O
ZQ�c�C-�yR!_�U����*G"4��B��yB���~ �Ȱg BĒ�ʲE���y⯊�H=����t��w�X1�y��%G�%�cJ%�,4��HM��y�N\q�6ѫ��2sYa�l�y�O<ad��@e�<y~���&��y���'�� `�vI5�Пpv-�ȓ�� q�mS�"?^�Pq�1�(݄�t�X�x�+�'kD�9q���!���E�B�Te#Tʐ�I�Z�JM��K���p�V%y����Nĺp�~���Cg֕���w�81�4�D�%[2H��|@&�9��� ժ�A�H�)Z�y��~Q� ����L����P�B&GQ���ȓ�����΄
����g��f�й��(�v<�-�#���� �Wm\4��Hz�k�%݀1t,��C �B1�ȓ<L�@7��9,��	r�i�/NX���S�? &��D9u]V-�Dك{̬( "OF�4�˥9�rE�E�W�H��ݫ�"O4!g�F�qa��砘�*È`�"O	�%(G>py��#ԁZ/4`��r1"O��#��7'��S �2`v��H3"O��A�IՂ!w0��%Ų%U�
a"O|�YD��)X���`��=M:�m��"O*e�ć�M��Y���%E�͒"O��YgƋa~��A�! �i/�1��"O,��OP��f �r�S�e�١"O��Ȗ#�D�:�Q��W9�xɹ�"O<��ˀ�7�tӠ �_�����"OPܸ��@_�^�x��қ4�<`��"O��@ҩ�,2[&�����o���3"O���#jK9mf�����-����"O���Č�:Z!ڠ����;`�k"O���p,��?(I��N%s6I"OZa��@���q�

t_P< s"O̅��۰~*��'Zg��X"O`@#bG]�a� ��ūWf)je"O���&��t���Յ\�
[��+b"O��p��۔���
F�|TY&"OBQ��%�q��Hg��$bb �"O�飔H�-o�6��5J�>F�$0�"O����bI9OR(��j�^4`b"Ou�En���d���*���iG"O�$�dII��\�a�e>ze`PQ
�'Y���+�f� ���M�/`z��'^F��0
�+J`���W�J.�Q	�'�T�1�˛'|Ȥy�eD���B �'�¥�w��(�����Β��lͣ
�'�)Qg�(pZE)eOS�t���'>n�� ��.T�l�cl��%fT@�'���-�AbЊ��9 �t�+�'���Ȕ"�^	�zE,u�' [b��"��p+b�2p �q�']��ڇ��/V*H5!҆Rq(,t��'��3a)�<���c1H�hl���',����́�&�ЅL�(�^�	�'!x��U��qD�貐L&��@��'���s.M3䦼A��GP�P80�'���  �Q"���I��O7���'W~�XeM�,�I��hB�\��	�'#�IZ���T�`[�	1�,8�'4Dm²E�$��	�Gx�$�'�ȡ	3C�{Τ�ѱ�9n:����'d6����\���֪��sxA{
�'9 �w�ٓc`�2FKC�|HVA��'G@� �̞;C� �EOy�^	s�'U�1������%���9��V.�y���,R��5/ǀ�꠳vn��yb�P	#�8�gSj�豂���y��Ք=i�a
ʱ7�挪qa�9�y�.�1�
}Ȱ�W�Ab,�"rF֣�ybn
�&�V�r�8)�� �!
ݶ�y�+;���"�/_�v���q�C��y�!��f�FPY�+��l��#��>�y���~�D@�P�i�^�3@@U��yIŠ a�ѩ�d��f�xp�#�?�y���d�B$�RWdR��y�B-_�5��d�8"�,p��A��y"�ֱj�^E�"��v ��"	�y«X�Dq&�I�h�����G�G#�y�jȮ q��ʇl٦����S�˩�y
� ����OO#8��*��ز,l���"O�۱!ϲ3)J��q咩i}I�p"O@`*T�U�Y�@PDD	x{(��"Ox�3R�N�E�@�%�N�^,t)��ɒ%I�>��če�|�bu�Ţ2��x��C#������`TH@	C����rA��V;�q՟��G{��)�'i���E�ǈ1�h���Ѷ0�!�䐵a*���G~i�8"���:y�Q�����mh���ɐB�`��祙-+�C��hΒ�"���#zt�x�9����'M ��M�r�V<�AoS� ���'�$!ӁH!�`	;Bc��G;����'�`��ޓ�:5)�ǋ1�"�+O���M�S�Ocrى��χǺ���]�qV:�
�'`�Jg�"�TK
,y�h
�'��G�S�U9�d�ӣR�	�j@c
�'}��J'M�/�PႫU$
4��!�'=Z�c��ΧQ\i�
��Y����';���F.P�ev�r"HQ�Tn dJ<���r  ��ҳ)�Ĺ���!c�Ą�Wt�� B �g0bӑɏz|ZU�ȓ.�iB�vN�W�U&�\D}����Jl�*��-in(��.G���C�	t�:�xRc��1�,\�a +.��b��E{J|*Պ�9�n��%�D�^���V�X؞0�=��OH�Q30�A��xCB	x�'��x�G�"�.L[�&o$4[V�Z��O:˓��Om*��#�ՒYE2��U���Y)�9��{��'�,��1��#�v52�%��Ky�P�M>����ՐJODx#V"��$��(R#�U ������\!�H�0 ��Ђ���"HȓO6�?��p�D"%��3�����)H��[�%<<O(��'��	�#,��9��&��F���o�r��<�g��m���I2K��e�x}9C
P�D��P���`�'c1O�Xiu�	�l�x$�B 0�hP��	�	�!�d�5	t䒔EČa�&H~����l�)#������ˮ(�h�zEL�
C�B�I�z��Y��������mܘ%B�I!3�^٫N����M���3*�C�x�3���6��r�,7lB�I	��h3����� �ٴSB⟰F{J?Ep�-\�%�2غ���(�A���+D�\q�|y���1�S�v�$lOr➀'*H
Zh�"R5:[��q2.�Ph<Yq�I�%�~�'-���@���~����'E%����)Y��h�ĩ�'a���`CP7vd$J�	]�>�2���O�b��c�@�O�Q���6z�#f���<5��'^h�s��h�܍�E��<�����<���IXۉ�Fz�	��*i��!2�ԝ9�n�@��
�y��L��y����=B��3���� Y3�|�l�3_G0�&�R�@\�ܱD�ܭ�y"1&�R���.@#�Ƹ˔(ӯ��O��'��O��������m�ae�LA�pY�'&ў�}R��F�a@��c�@½j��,R�G�}� �'�&DR'Z�v`#�C�HU�P)]9yB����S��r'�?��!�N�����O���<���I$_�by{UG��b�.�"W�8K:C�	�{w!����&��m����J3}��>	çG�x�X���Q' ��w)�F9l����hy��ݔ����CҲ9���B���'�a{���x�J| ����7c�b��Px�i��6�	�3"24Bď�c�)
�'�Z��FH�Vpp;�B��䙣L<i�R�3� �0�g,�Lx6�3��mz����"OTp0 ��U�>HPV듆
�� 8Ol�O��?����	#�N�8R��	6z�}(DeݱLe����?�	F�ZQ8��p0�jᚧ*��(�=)��fA���'����f��+Y�<9U��2\�x���{��)�4e��+ƮqjǆL�TPH1��Ŗ�y�P�/�a}r͞k��r�Ɠ�E��8BeO+�0?�pS�,�F�5U^x��@JQ�.�\D���.D�{�b�Q�Yt��x6���.�O�O0�x�D�'s�$q���͏km���"OJ}���#�x�@r��'
n��"Ot�u	�@�&�(�ʒ�[a"Oةy�/���Z�1!�$$1pc"O�@@�7'����w�P�D���7�'��O$!Ħ�K�Dp��ٷd�@yK�"O�ųrϞ/#�j͛4��A��"O�S�G�:�5�pIC1i{�t�4"O4�9c�� x�a�Eh2`�(!"On�i'䅀[G��v'�W6��9�"O�k0d��IX��f�/2����"O�}+��?]I�%�$�<o���b�"O�����.���P���?N�t{��'?�'�|�P��%d���) �#^��r	�'��B�	�!_��X���L�P���*}��S0%ʔ�`gHӊ�̕�#և{#6B�	b�=�cG�X��]37dƇ�RB�I;{ghM)V�8���`H��(�(B��
wA
�J�&D�n��� �?'�RB䉭BdʕQ�&7�`�0�
1$B��5Q�98W���2Tas�+L��>���i߆ 3�尳Z��,�k��-Pa{25��9'�h1�������n�_��)�S�OY�p)�	Տ(���� d�r��E@�|��)�SQ@pk�F�*#���sC"b�NB䉯[[��+�@a�F9��[�mT,���9?��%��S�AYqaҨ!XD]� Y~�<Q'̟6�`�i�ڸJ�5;���<��'�qO?ɒ�A�Fg&�AN�a����&�(Or#=��� (3(���_9\Z=��d
џ@F{��	"Ȩ��ŬvM���L2x�>C�	D����re_�xt���טX�C��3;�	�3�H�(FY�c���@.�B�ɞ5�l���M,5"�Œ"{˖C�I�T��t�sf^7y�Q�X�x%��$�S�b�O�6X� "��b���YW�
;a�B�I�S(H��b�m-`s��/K���IK؟\ʔf{=��a6Ɓ%o �����/|OXB�O�m' ��MW ��,
|�`I
 ��B�	/�V �7��?b���ebư5�#=i�[�\F�ԃ_^��Y3G�[:(@qQ�L1�yb)Q��Ъ��®F���S���s푞dF��'�|����$�,m���@LU���ēxI��C��5SGņ>42�!���y��'�<�a���!Bf�-���4K���c��y��'���:	���P�E<r̂`��*:,���O�U£�1~fİ���$O� �ȓ-�&I���5�y��@�V���訓aL�Hcf�c6��q�LJ>��m�qB1�$
i� �> ��ɉ�Q��ꇀ	�"v�����K�$�jH3��>D��	��)�>�bp�
:>�:Pb�*<D�lT��:|.h����"� "tQ���	�`���D�J���`@o;O.�B�lU�|x�D��X����R0���S�? �]�$8����o�-J��Q��"O���!��h��ɱ�����9J�"OB����Y�dT�@p-ģ!�ؼ��'b~�Y�յU&���l�8S��`�'����V��;��`��G�@���'ZfؙfA��z�����������'�:T�3�1���a�N��L�!�'�\��2&��w2T�BL�y�2���'��;gE
;qN�h@��v�$���'*\�����C�I�!�!8�^�[�'���CHY55���`ĕ��ڝ��'"���.ݟ��]��@S�}f�9�'�R�*�N�9��* ��r�:�'>ޘ;��[>/�̀�E'P�zx��'�F�@� I�P&�3��O�|�T0��'9���5FU6o�n��݄/���B�"O<(x���8o�ڼ9!��Үي�"O���6��nZ���"��Um�M��"O�\93�*kFm٥o/`��{"O4���	��:7r\��OS)DWZ��"OfL�D�P߼�$�N�H; A�"O�x�$L��	��<A��.?���CA"O �J�၌VY�(��O�_����"O��rs*�G�v+ �Т�Y"O��b6�
����;2��q"O޼i�	΄[�t�7���k�½j�"O��1G�Ik�-��K@$��R"O�@�l�,>�n�ە*\��D��"O���J�#���ԟ�mY"O�1#�E��/Z�Qto�+�����"OBQt�2x��a$V�r�|[�"O>�93��7|w�Z�"�VM�2"O�̐'n�(2lYhT!XyԜ�T"ON@)b��v�p�4��Te,�*f"Oh9I7�^�I0t���R<�pɫ2"O��h�#B�܂�����{���"O4Ur��Z)2�� �I":-�"O���	)&`]�V̋�_�$)6"ObdIj��|���cTʉ5�4�5"O���`�@*	g� hu@V�J��Y�"O��ɲ���a"���%�i��* �yJָtl�:gh�%iJ�Q�/G8�y$S��80�ꌓ[�!��U��y��W�	?�٢vˁ�Y)0�yK�yBfټW��#�J�BwR�pf�"�y�,v��FaZg�H	S^.$y!�ğ�T�V��W���+C���"�\W!�8����$�B�ekV�����nX!�da���%�.Q��)�bC��5>%r
�'�.qз �X�1k�z+�a	�'�4m���ذh<Q��G�G2d�1�'O,�����s1������6�H0�
�'��	Z%��%�C`\�l|�'>���!1�hЙ�ኄ
e�̓	�'���$M�'ժ���bׇ'�]��'�.U�R%]�s&-�r��~yx�8�'�<�â-X%b����A��i[��k�'���(��;���z�"B�(�c�'Q�Ug,�"��t3�E����
�'�L��V协^�|i�
����
�'u��"^�)�9HTn��vy.i��'%T�5▽��c�Ȳc�5�'�\��P��,3��2cF�)��Lj�'�����J�P<�r4L��,+D@z��� � �mޗ@�"�X0�G%l���Zw"O�,��L�'� �11MP	V�T���"O%x���7 zĭ�P�Yؖ"O�XF��y�")[�l
�#�@�2�"O䅙�i��|`^́��x��"OcR�V+K��iF�D*�V��"O��cw��7�|�a+I d�iA"O�`����,툤�-"\��ip"O65ABa��L�b��,SSV�1q"OlH�J|���z l~��i˨�y�	)e�$(f� X�X�3"��y��R"+��1R�Z0QA�yYb�-�y�*խ$�=���QQ��9QI
b�<� n
!z�����G�:��r�ou�<yÏ
#bh��6BF�vv��B�w�<	�Z+�΀�7�յHx:��Ix�<-����� �bE���0oO~���2Li��L��t붜`��3[�Ȇ�4���Э%��-c��ч4Dņȓw�P���TiJ�u��%nD���yFl#���i#�ɁrN�:J�JĆȓ[6��ˑ���*��E�R�������,ٹb-ф)21��L�-3T�X��^����Qg?��Qg�y莡�ȓQxe��'��)aU�*V���j���ԤݛJ�<�H��h��ل���Ԣ$�K|G^h�kx�x�ȓ�<�w�ܑ,���3�@�J����<9�E��K����D={��٩'�Q�S��T�/Ϫ��2	�y��!�⎗�O["����5V�`����/�!𤎯MM�(�%c7���%,Uߑ�hz�Q�Ԭ����?�z���@ŲMfb����y���o��(�G�8AS�l@$Y���DF�>r�!�B�#��)�'�
sF�D'�f(�y����ȓ@W�8��S���7�K�v���L�x��/�d�91M|�>9�FZn8�H��f��,�	V�a؟p`�75h��Ǌ�?��:�N7 @�3A&� }���ʍ�q�T�Zu�N�B'$Ā���O���ԩ]}�*I~�� 0̥�-ơ����D�<Ar �-Y|��s��T"k�=��f^}B�!�qۇh_��=I����4MɼA��0�?FaC�	��@�.A����,6��4HCAY�d[�ZjH�Q�&�B�3�	�#��1��R���4`�l:^����䞤!��-�Iߡ��T)W�S�8N\	z2"���B�ʕs�>�,�fLڏ��'��$���7
��񁆨 N�N}�	Ó?~�Y�t�/p�^A�3ƒN���4�N�>�l6-_+*x��x�遴t�n݁ϓOĲ�!k@�Ji�����K$����	#�zm�bÉ h.0��|F�ju(�,Pĸ�����!NԄ�ēv�,� jF�
̪����W�N��=��éc�f��%@T;=@��d׸?��
�L�[�,mjsL��yr!�;3$�d6��o���3R鑹x�C��H�g���ȦI�O��qF;2&�lN?˓$��4U4a�X!3��ҫ;�ș���0T��b��]~"k˒�F�Z��T�Xʇ�M�L��0�Q�թP�di8�� ~�ay���hi�J�s�&H�V�O���s�,P�&)�<���K����ۧ<����D�p�z�JYS�H	�(C^s$�e<$�ԃSJH�t���b��X�b!��R��?=���Y/O����,˙F��B�fܢ3��S�cS�λ+z�9�s�_�/�:�Ah:$�U��ް��f�!���0/�b����۾tg$��J���P� H۾�s��"�
�gy��O]�j��W���i�!Z���<yT��Q���Q�a�>	�j��=d�H�R(Ҏa�����f�ۦi��'̗\U�a�R5W�y����q�JK	r��Y����w��9m����i(O>���'�7/TH��R<��Ǜ[���Q��w�C�	�I?� ����(��r���i���tcO/xڴ�r�U#%��xi�(Q����[�_khe)�J���Px"�HU�? �$�e�Cn]�6��88�M{����\�4��Q �i�����	7.�`����ǎcP��f'S06��3�MU���Io�(��k�h��3��c�j�9H�7U��M9�"Ov	��V�3���q�BA!�.���Dؙ�}��j�6<n)Y�F�Y�OXh�O[}/B��� �b'��O�<1F�_�����ƀu���4h�fc�U��(O�.�h�a��H�(h$>c���6-��
��}9 ��8z�%[�+?�O���7��5C�1 d&��B����j	* ld��@ Fl0J��J#������Q], s� F,39�˲�<w�Q���EB34	r�b3C�(Q��3w
�����G��z�0���K��Y�"��R�<�FHy���PHF<�X��g�<�'��!�j�#1�D�L{J��6�x��>�R�-�?p�ћfBNM�<�,D��ULI�jV�#D԰F���[2�RÞ0q�&�ENS�J� I���'��(�-I6X�
t��Ɉ�1o����1m����΀%r�����Jm��E�<4	�I"��^�h�H����^��0>�3D�,oQ���>U�pa�Zb�'���U��f/@ 7T�ZRP��8�!
ϲx��E�e��"O�tض��:mJ
�A�����3U�'����v�E#UN@�j�>WR�d���Ӧ1���� @+z�f�ϓ'c8��ӂc�J�$�P�:G��&��ׂc�4H�$�A�;C��h�H�T����O��ٴA��F�t�	�
�Qm`��$Shnܠ����j���cC(Ғa|L�vi��E8|�&�	93�,99&�'�O�A8Ƀ7zR�BD"�1x�����xD\�p͟����_gd�-�'z&VQ�Z�u�iąk8b������<	F�ܟV�^�p��)�A���y�J0��1�!�6*��1 v��_�Ox�XA(�P����a�{�� "O�Pa�@^s:%z��	me�Цc�U�q1瓢u����fHh3�3����׏1�F�S�Ϟ�=�E�����*�hP�E�o���Z7��|D i��	;�.D�K�v��]���'�(�Q��Ӳ�:� H�8R\�R����g�05��K�:����~��^V��BᆏĮ]���#>OzQQ�K��p>��/Al��q壜Y���G�S\?i�-M+���R��>X����7��|Zku�t��O�l�:T�5L��x3#�e{��Z�'���
���T!*��Ù�`�.�1GJ�."ސ�P�?��9ƪ��r����ݟ�N�T��ϻTSF�x�F�'=�P� t�
���TQB��b�&+���s�
0��H��!�I�߿U�ds;O�a �&*���K�bΝ�C�<�P��
(X1cr�٩ް<qD��+R�"f�Q�W�ıo?�8Q��N/cZ,���-C�*7�[�)w�������=qWC2q����$�D2gNB��`�A�Tub$.�g�X�	f�
�zD��B����ʆ8v�#bEڑf0�2DhРB��d�!���0?�
w�����T�k>�m����<�T�W�Њ9;��9#�P���T	���c(i;�e�[wX�Ά���D�EE��<�(��ı~U!��!�N���*I6�L�4OZZ]A�ŏn���0c/��I��فŅQ!�D���h��؟O���Κ�x@�oׅ3�8�2�DZ,U9d����)`D������M����.S�p�,Z�U�8yp��6n��q�&nƨP�4n�P�Zw�r��d17t0���n�%�c�ď1��On��QF�-dd4��'o�5�3+Ď0��T#�c�xj�
�WS����%��@�F��s�:؇��MXȌ�$�ͼ�x�A�_=T�h\��%�9K�ȗ'�TͲAS�|rc��>X~\��Ou�睞v��H��
_U�48[]�!9�Cx���c�iL̼���-Ab����;>4��L�(�$X�B��H��#}�%,��\�p7���Kި%��(�Ջ�*!���z���Y�L9!�Ao?��k՟���"'��V�~*s,B�XF�<����u�BiHu�>itM�ᮥ�К�L��s��&`�CEe]<��qB���#Qkݫ)���G�'Hȥ0��>�Խ���L^��^�n̐�+�-t��Q) ��v��@�&̨���J�v��P�f<)q�A�j֒r֠��� ��dțg�*��I8m��-pp�p����ir�A����٠My���#�49ڶ��"�X1)�4􉏼AU|t�6W��9��أKu`�(s)�A��`i�,V=n*xU+�G0�2���l���7Ut�$�ȳfV�W��+k�6Tҥ(G�g�8,A�T�H�.$^�|�B�L�5���մw2�24Õ���%꒦
�Pq#'#Y�@��`к#��� �k6��
Pd/�d
n=����dK+�B��� g<-��H�&��db�)K�ɀ�@Z8�h�EU
N�|�xv)3��������J�&Ȁ)�luLf�q�	��e_�3rlɐ��<a���cS�8SjC�\���-ŷl�-˔nѨ_�8��E�O!J�ZL�v�P�J��ꝧ�\��"dR���$;fl0k�J�1?����N��ў0����K�Č�l�d?a�bѽu��D�կ�4~� 4�W8��smO�Z���_�NT��4>�h�OJ@�S,�5�y
� F9�&ܟ4�s�d�	^��Q�'h���!21B�<��U�|CSN�q����D1��F�7Ɋ4r�怉D?$��烑>r+v�A��(�9���E}�_������Ib����1�������%g����ǂ%���I7s���x≉��0mȘpƾ88S�,#�������!��i�
}�KѺ)�\�bb��	�@H�v�0���Ц�,�����L&�܀Re�$�0Ҡ��e�`p�>����߁��0fL�QLrq C& D��xG�CH	 �gǖ�d7LIKP'��DZ IX=:�� '��}�@ͫL�8�1��L<�4�c��M�<�@���mX�?Y��=��M�L�<�#� 8h�,��A4W��)a�W�<��*�3� �2�]*3�-r���v�<)��Sx�ݱ6lΏ�v���a�m�<��@Ľ`Vbٻ@�1*�,�2Ѕ�s�<� d�n[BW4Ţ�; 	��}�!��W�"-AV+Ũ�{e
�'�!���N��+��"ʂE9�L޳?!�L�1.���QI׻4�r�,v�!��i��S�Ӿ=^���ځ�!�$�~��q���xJ�*�k�!򄗜P��K�ҜCG�S �!�Ĕ�O.����J2u��-���K��!�d��S'�mp�I�* ��(�w�!�č�n�������A�$���3!�0|�t�,�0?�Xd��/��!���_# BFN��!��dS�?!�!�D� 
�(+�\+Q�f�#A���!�Dʜje���I��#s��"�!�dЛ ��=b��'2����B�^,p�!��N��^q2�&�,�4o׉W�!��D<I~(Ia�(U�|����(8!��_�2�X�`��f�D\�틯9!�#=r�3iF�
u���ծ@�Ry!���d�. ���9Tx�+c��k!򄕀't�s�O1rU줹 ��2�!��Hw3������4������&%�!�dȜ������D�L5��
�m�!���(� ��Cn��"��!��øCp!��F W���1Mk�P�ԁ2es!�䜜+�Ѓ��]�%����!�䅩U���Q��|������*No!��<M��L�"Qӂ8h���[&!�E�N�@�Z��[�$�<!�N=z
b���L��Q`P0��A=�!��ܞO�N�#���� e��-C7v!�dC�3�,��DݸJV�Dh$m�/!��Y>dx��-J�j�$�!*/�!�A?`AŌC9��	"��ŀP�!��%F���L��|; �ȃ�Pv!�d�T`iA�=$���L�y�!�$�3hRAr�!�/u4@U��f�!��'`�r��u�	�{� a ��{�!��}�N����F��R��(!�1*c&�#rj�~�	��@�!�$M0[OTI�*Ķv����e�[�W�!��Db�}�$�s�p���d�!�$<0��91R��1��YbWV�?!�dS�d�x��G��@�ak�)ֻQ�!�@$M#&@���/b�R��� �!�$�8�P�:��>@��`K��O2@B!��+8���U�3w*eyr�%s<!���[�r�rsnQA����1
3 �!��W*p⩣�"P���z �D�}�!���q�fgޕHl���/�60�!�� 8�� BɽY�8Mqf�����B�"O5����::p��wb�T��A�"O�X�o�7q���,�07wr��""OZݑ�+H=<�l����5Ѐ1"OX�C�*�'l�<	��"ǖd��0p"Or��� ׄ>�J� @�Z���"O�Q� AI9P[ԍh"��"v��"O�E��j.d�ܻ₈Aa"�q�"O@1�$��)��BS˗�Ff,�Ip"O��;���O���۠K+.W<\��"O�!�֪žso̝@��@A0�H`"O~���E&z
� �U�� :U�""O:|Q7Sg_!enK>8���Q�"O�$q ��g�*�*ԭO�I�D��"O�J��%_����,Of�S�"Ov�둬�3I[���1�t�aR"O�+@'P4xB�1�i̺����"O���O��AD���߳d�&t��"OJ
֮ �w���C����@�r�<1�E�(@)�,:��EH��i�<YrH�*Y�����Ɗ�U���-�c�<�jB�k��S���,���3��S�<��Ź=����YKH����HP�<���+Ɛ�A�K���\821��Q�<iwgͲ+�
4�Y6>�pQ����S�<q�۽TٖP�E��	�R�B�TN�<�uh����s��u�D⤌YD�<��#�WK&�2 �$ ���I��B�<�B�?%xԍs��U!\�����Qu�<I�%D"��D
��V0�����]�<1�#I3/�	�5�C�3x2�4CUC�<A�ه�&ق�EKxzX4�}̓z~H�;OLQDK�R�E��!K��h��'	HA3UT
/*h�x���)���я��kJ��O��y��>o݊d�bIV�9�b�@g��+]�e�&�[J��O�js3��ے�H�䙄_@%��'�h�V�,=���Q7��W�V�y�Od�I/�VĬ
M�"}��5khP�Ȓe�g8`��` q�<!&\�<�H�: oF��`���	�vʼ Qi��g�T�bi�T%�N[���`�a�����I7q������_Mx��ΈK���q�W�le�����'%y�d,6���A=S�-���d�"$�x���,L���'i��;�!_ D0��� �$��	�ȓC>�k���	��$�84[�-�'L�H@��"oΩ�O�>ASu�̝�l�ȗ�ȯ s��SR�*D�P	����P���ɰ{�����WU���c�'��o�3�	9]���Z��
@j��UĘ�h����9_��sc�F�v�t[a���jg&xHR�14Fh�c�˷�ZʓG������'�d�p����yrF��@H_�"�q�πă<�	1�f0��[**��1p��
�:ϊ6-QD�6ake�չ�T	ϓ.�W*���u�p�Ę*@L�뉢d�" AfJ� 0��ȟ
�t!���11j�E���65����Z{�ɒJL� ̪5ꗗ+-���=	�˗~���3.ɔQj�����P
�L�Q!*�_&�hb#�y"a�W|�e���J�VĘ�CΒl�
E'\4x􄤙�)�O�8Q A��V~�m�O?˓Ka�l�d$D��:�r㇮s����l�N-���yybMж&وL2�#��X't�"bH-B� yS2	'U4�@��$���$D'H<�K6��[��RH��'��bd���Fp�'dB��P#,jI\�ʉ٧�ۜK�n*afߠE,�\�O�E��'T�t�P:Fz� J��&}yJm�'��3�h�6m���Y5%;V����C��ݵh��!��Ӹ=�j�zE��-A+@B�	�3�2�{�	�3)1��/�6R��� �B�"��8���P�J�ˉ	1�&�2IH�+�<����-���ҧ�6�bh��RIx����D˵�vt�&[��B�Ւ7|�0�9>]|��D�h��z�&�N�
�'��<� ,Iв�Q��y(�J*:EKr�|�
�+	"uf,��ɫ+�4|�mI�?�'��^R��3�&<��H�Q�<����v0�G�A�.̨@���A�.�>q���~RE�O�b?ORx��lҮX�����T��q��
O�Dj�"D�l��̈́�
�-53��h����#k���ԍk�a{��߲f;@$+0 �0���*�p<�l�i�n8h@d��K����4��I�* E~Qp�n��>t��i:�y*ff��Y&Ҡ��n4�p�OH�y�l:�f����L��"}
5"��F���A�B{��d�<��Y�B~��Uhî*�1�&���mV��Q$�� ^��Bزo.VI�}&����6�e#�b��a�j5r�=�xZ��Z�.��Y`����Q��$p������� ����K_؞̲T���4������= �2��;O�ܣ�ʵZ��X����(l�(7mƜyyʈ��'���P&M��Y�!�d�5�ڥ�$ܑE���aʚ�6]�#��9��#�5k�0��&�;�H�ؑ	�A��/\r8������ё "O��ӡ�9�±l.X)ĥH�lP�;�]�#���Za������lXʌ�k�:��t3���t��Q�򙲷P��!Cv���N�&�X�j)z�R�)���0>1wf���P���`VpY�l�T�<�TP*x4�PD�P$d A�l�N�<��I�|Y��{���9O�6�@t_O�<�C�W m��-�a��."�0��'L�H�<� l�r��:�=+��%[�BG�<1H�"+�$<@��H�q�1�W�C�<ɢe�(!Mt .�-s@@5���Rx�<1��مa�,��č�r��m�Q�<Q��;/Z|(k���8���'�R�<�%�@�e#hD���6N� HV�OH�<9&NK�U��
�	Ҙ��ӱP^�<�p�͟%�e��уS��g�<i@nG ������yע�X��\�<!U��i~���O�:m0Ī�]�<�WCT{�dyn��t��ЩV��$�y�
m�����C1v�|M7O�yRO�;k-<��ɈM�=r��f�-�Q���tz��<A��H�L�˓lIz@P ����P�3�L1 �.o�(t�`ޛ�y�a̻?��ɩ���- -�HS¬Ӄo��k��DI�|BԄ�PF]���y7��$�����	�	��2�ȑ�y���(/L��*�	�� �r ��}\��B��/#}�� Nl�0���/N�����M*H�*�bd��K: [`��8L��{��@�L.��$n���#$m>�q3cE�cRP�U�~����M�>dh��ߓ9?@wC̷x�<l�e
�|\t��?��o,wf�d�f�p�P�;���:�ODH��q˄J�r�p��6U�A@���H`��18�,�׌�	�:�#��$	�<8�c�|�L̰�=OjY�0@ 72�8��'	�2�QeV��u�0���J��H@�NN�a)��:�"O.��GL(8z��ꀏn���.�8rڸ�cF�� ��&A�Y�*���)4b6�� ��T���\%�c��p:Tf�!��X�Ы>|O)��
��M�4ADb����P 6�*���M��	A���h�Z�R��M���X:�uM5�HO�,���GhT�1�:Q��������;Y8ad%E��~"K��S����O.(�	󌜥yR$Ly�Gv�<��� ��5��i�W�BTX�����P���H�`LPi�j!�BI��3 ��Ty���b$�Χ*W&0s$E�@�^�}�MKө�X*񚇣���Tjd�#�O:D[��F?C$�5�	'�v\�P��:&��;��Y��`"�����➾��+�AG��|�u���dZ�H�iN	a0U�r�Ny�'��5���ʱOr�Yu���"�f ����e@�t�Ю�N/�1��>��a]&�JSb��L�����<@�z}��j��[�t�p ��҅+[�TTh�
�S�ԈWȗ.l1PY�e�~��dS�F�����eM�2l:�A*�H<�R�J��]]���]J8�BD���Bg��ѧG�-�`h�`�� L�I�<9�]��m���'?��h?(X�X�xq��Y�Hٵ&�q,���2+�/Xl�d��+���/�P@BR=D֨-�e�Q�V�z�B[
Ao��k4ͺ<I�+]	j'����1��	k%���'88I�6��>: �ВQNv5x��h����s�ˬ�>�i�'�.\˖�޲�|j�cndJ���OT5uQ�-Ѱa'kbl��&�]�@��d
�	���z��D�0�h��-�B��$�)ޕ尬X�g%P��DrC����Ơ
 �uy2� ,�;g��j"bِ�O;�(3W�'9�4c�Hÿu
�D��R�>�k�<)�5��琭2C�nӹG����P�Y:}�i݅oe\>#�-�'�����`F'��!�D�0N����D^�356�!BH#o(��)������ ���D.Q��� ���G/��@@^�`rӠ��l��I�?HF��1g�8R| ��b�!���$��y~���E��*��$!��c�Ԝ���>LL��Iϰ#���H%��-7޹2��*8����ɜ>>y O�5DR����͔	�b˓`�a��5V(p��'A�	�	=_��'O8\�`G�z�j��fIֹW��`�W��X�d�g�K����tɼ �6+Q@R�@&N:�xB	�8'$�d�V��5p�̀"����O*I:�$������)�~�r��i\BpB�H�y����m��x�k&a͔�Z���0�~"��Y94{��|��iyMЌ�TK� ��}�0B!�V�
L��c
�c� u��E�)O�!�$�L:4I�6E��a��0t��S!���+v�x����^T	ĭ�ć��&�!�dȕL��)�&5~l�v咄A�!�dJ\���JGh��\ ��ӆCR�u�!�䝸](Bpj�
̵i% <�^�#�!��Y	�%��'�A,����!����TJ���8:�,��e\,i�!�$[N8�aeF>�IyS퇿M�!�$� ?��`gR6x���8�텞md!��p��u�A�˂8V��b<PW!�D^	C
Z�J�@���e 'N!��V�5��\ QE+��Ȫí�!)!�$C�R�2q�Ó-5G
�*P&�I!�dC�A:@B�	,&$$�1�%�=!�	;��s��4� !0�Cݸn!�$£Lt-qU�S(|��h
����.�!�$�#F���bŗ�c�.����3M!�R�:Q�tx�%$�Π��Š8Y!�D�8�&i�pN>/���ڴ`�C!�d�3Z �d�ࠈN�)��@Ģ]k!� �w$���@�)�ta:qn͛eS!��A�%�Ԭ��i�@�d�!�+f!�dZ�%�J��B��3_0}�!��]�!򄆤w/�4��ޔ*ր�Xa+ve!�$��}��Q��ʡf9�}�V�JP�!��R�mz���f�E`0ICBE�z�!�d�e��\Rf�B2���!�=w�!��u����*��*}�5���!����HH�J�}�|�a�4g�!�$J6�b�Rv���;A>�Z�*E��!�d�n��4K�# '�Ը􉃡w+!�D]��hWΞ`L��P面v��Є�[�q4@ g^�I
��֞ZF��'��	R?�	�'f�rYy#`W�;�h�x��O|�`Eo��~��O���S�OT�p�DZ`�I��g�-��i0�y�W����ӷj����E<r�ܝi"�ǯO���x���'�)�'	o�d�TC�;o���+���U,�I4����4򘧈��!�m�=�̡A�-ߙB�ua���Q?9�y
�'m�E
P$�k��E��9���	d≁s"��Mz̧����gbR�:��̑ô��,���'(�m���4�1�'X��Xe�Įd�6��`�\Fl�(O��� n#�)ʧ.��`)"fz��q��Z�=�Ĕ�I"ctT�?E�Tk�sMvH�T���YjP�1W�P�\��3�yB��O�S|O�:�J*>�<	K�`) �Rc�C�@-�S�'�21A( Giv�Ѵ��/g��'���b���S�q&��q��̼@��ػD �. 牞'��"<�'y�"��<����66���[��P �;?��hGx
�'u���k���nXh�8Q���0VZPGx�
��0|"F��"��"K�!HŮ�`�(Goy"��-�"���|��$�pK����_m\��+!��j�O�=����8p�)ڧ$�� ʉH�cZ�I*��3(���ĩ@��O�����\ 9��N��(��P� �8��ױ5�2�y3N�&�ʌ�SN1~˓�~
�'X�2�K��� C8ZyB�R�-�:<���<a�'Z�qp��)��<9j�Ȱ[4�d0�A �h`1`�$P�M5��>%?aq�<$�&���2a}ԨAc1}�	 e����=�*��#�,�i�->4
��ж���y���P��M����	�G���3�Q�s��m�� �1[r�y�.�1�fN��<9v�!� ��� I������y��B�"OnxC�Y��Ƞ�ס2
���"OL�1#h������Y�.)T(�s"OnQ�0�ā~������Qn�P�"Oj�K7�0�∪F�М	����"O�I 3�J�,얱A�	�*��u��"O,�rp�E�*�@
��q~��� "Ot�[��Y�R7�9z�%E7D��ؐH�$����TC�ҺdÄC6D�$�!�Y�M�Z���DXq�2D�D���P�I��^�Q�����-D���%b�$Nx���oG�0.�i��i+D��:'�����C�c�G�|���)D���r��QK�3�/�,�nu!H&D�� v���Q���#� \;EEJ�w� D�H�r������i�B�@�g�&}�C�ɆA����,,l�u����C�����RfB7]?|HF��1	�C�	>g�d� $�޽R������=r�C��!Nj� �dh�-a������$@��C䉆9�	b����!b6쒸��B��/&��x�Q��1d�iT��7X�B�I<g0�4�@�^�|�*��Z��C�*(pJ��a�T�=�:s���=j!��"����E� :�YB�\�!��C�E�HR �O�"�)��_"Ky!��ُPR0���	��_g����7<e!�^�<�`��5e�?g0D���؅uG!�ĆZ}X�1@��BM2h�e��71!�Ӻc7*�05��{�5�&oߒ\.!�$���AIS�K�d�%��g�`�ȓ};���ခ_(~q�Wb�0�����"0�=8�+\�l@�r�#�
\(�\�ȓ%����dS�b �]�go��gŨ!Z�cA5!��9�Bm��ȓ<�0�����
7��b�o�`����i�4�2ǔ	o���T�Ow6���W&Ҵ�DdJ�����b�%�쉄�-`��XFNT�c�v$jD��.��)�ȓH�A��l�b�%ǥ9�2݇ȓO�|�"&�	v��ܱ�^ =�����MrF�
�Cs�ajD�!7�$�S�'K��0 �H�t� ��,�0��'�����ڌ<��[v�I�>`}S�'X�1��ͺ�(�j�f�k�'.P�8G�ɺy�晁il��'���&��%PY\j���^��2�'$6����ap�M��BۅT���r�'��2C�-Y�B�y�� �p�'H��7hъg�D��k
��^ѐ�'Y������-x~���<���'���Q �,S��Z@K	��,h�
�'����W��"�84aF�9�@	`�'_��P��L�~��9�@�,��5�
�'#(�e	ʦ�;���S��s
�'WB���5(��V���M���'}Z	�%�V� $0P��@�Wir�J��� �I�$؂YN�
Bȅ(,I����"O���ǋ"8�����&H��<l�"OH�AFĶ(��E�A�� �����"Oz¡�զ�z�ɔ˚2x>�`"O����H[2���.e2���"Opړ2��(�#
ҿD��Q5"O�i��?GJy�$��	`����"O�"� H�,�҈�Xr1Y�"O���c�F�	O|Q%̸��!iu"ObY��,wlDQ�D�z��\�D"O�J ��b*�����)�6H��"O�T��#Hu+S��v���T"O���gMIo2�ģu)�I�����"O:$ �m^w[�� ��R 9>���"O��x�'һy�ڙ�P��=��4"O֙��F�JS1�vbF�HW� H�"OR�"��T���
�6J����"O<i&��4����,�� �C"O�X��5U�84�����1!@"O� mͬ:Q�H����L�v��2"O.P�eJ0&?�1b%h
?�� "Ol�0@^ [<��"cf ��.<�#"O���@� wĺl3fŠy�½q5"Of=��@�ip�{�Aڌ"�R! "O�� ì&jb��v���T���"OP����� ]�g�c�q"Ot��2��>T{�\� I߃8QN���"O�bUgB�)�0Ղ�	�3l-6���"OP��&�#^-����4}P��w"O�Е��3X���GH&Q� "Oxe �]Q��)p��y8�yh�"O��s%D�7P9z��I�H9�"O����&5�Q��F
7��,��"O�)Cs�ƏcF-9��ȋO��� '"OZ�r�ds�d�(�t5�W"O���fh'��������"OZ!��d9D��a�u�h��"O:�K3��#��p p+[5�6US�"OnQ��$�� "�3J�9T�h��7"Ojyp���$XH}y�F9�0h�"OفÁ�V�(Dp�&C4Wja��"O���A�	Q>|ɰ&�gYн�"O������M���f���9�`"O\�����zޖꦯ_)e|��r$"O�����O�I5�y�7a��\Z��U"Ol�aL$
`0KA��i�ɐV"O�u��/��i�̐+`<HRHj�"OX2��"`&E��؂�|�5"Oi���B����f��5\.h���"OBaC�����!H�#C5\4phh�"O0Y���תr�|��"AK�ܫ"O�5r��޳ � �J�1B��K�"O�PI5��=p-�Us2HѓG��q&"O$�sG
	0��X���s4�)cT"O�p2*��+B�ݸ����G6�LɆ"Of$9G$5
�ũs����S#"ORu(gJ� c�u�h4%r�"OB0#VdE,!�����AԟM��Q�"O��ӡ	hfHꔉ'F$ԘB"O��PO*[�2�!�ֹY:$���"Ov�6�h���� �ȭd�4['"OH�B�KZ�+���!@��r���(�"O���4�r�E����Q`�U"O�<K���a������
M�6"O� 2����|�duB��#=�D�"OX�+D�Tl��)9g�Sl~�	A"ORT����6ntqQ��]i���G"O�\2�"Sq؅����OS(��f"O��X��r8(!�_�F�ƅQ�"O=��R�P�lXb*G�?Z���"O�<
2�<GJ����H�I䊅"O��:�bo����z�,z�$\�A:!�Dáq�ʘɠV([���פ�='!��!u��<�f�*=���cA�!��Bʹ���S�J|°B&�P�I�!��^#�@���)f��)b��ʇ&�!�D�	V�IE�١� e�U���WF!�dܯ$��K�lXQ��� ���*�!�Ww�$�+W�?�D:�#
�8�!��5���6EU�>y>=�-"k�!�\/@�<��4���_ov�'.��M�!���'-�t��Jxf���D�7)�!�Ы3�5�d���bB�0�<7�!�d֝j�P���8EP��G�X2�!򤒅U����1`ߺn0�<R�d�e�!�V�)�����(#��9�T2Z!�;D�(뛾=�ʰ+uLѩ7!�$�0n`��� R�5��GKZ�#!�DŒ0+�%���`���0���" !�$0s�T)(��M���2�B�i!���;�xE*�J
&g��0�@m�]]!�$�R�$
B�Ͼd���x�ڤQM!�߭Y��aq`M�*b{���vE�%93!��h�
G+�l��9tD@:P!!�Ԇ~*ft ��Q*9kMz�#��J	!��	�D����$��TZDBJn�!�$�5cm�]�*J �"a��x�!��SK�8t����.����h�!�d�r*��&]/{ry����!���)a6��
ŠRL�v�=A5!�dǧ?�PZ��͑;T��c¡S�!�$��<	J���k�)r��C�ʬ]�!�O�'8z���� K�����K�!�dLku�Reߣ��aLM�!��н
Q��2�Ǫ'�*�z#����!�D��=��#b�O�%�0��(T�!���	7d�Qb`�?A'��h�C��!��R�Bu[�'��E&xy�C(�7p !���m���ƧJ��Ǉ5c�!��p��͊�}a�uI�J�G�!���Z��I�TA�sS�D; ��(!��[�DC�A(�S��e�<8�!�$V�LZ��t��aH������Q?!�d�%~�+��.�T���¦f:!�ɢk|,8[Fk�?����R,�)>,!���1�F��a�
����FL�%rn!�D��0����)ef�����V�!�D�1�M����{�A4$
�:�!�d��o�b5�"��S`��{��F7�!�d�s.���P@��%���#5-���!�d2si���qj̶��mҡ��#z!�D_.|s^�*��< 'v�@�M��9!�dά��Q��D&Y�|+fW�|�!򄛱_��H$D�x*�8
�E�/G7!򤞅_"��YRo	3f�Yq�D�g'!��yX�YK��^�g�Q%ɕa!�Ĥn��T���R�drm��ƃ�!!��#Y��`"k��Z��YWH+2!�� ���V�'�BQX�d��8p
L��"O�Y�d��~��am�fi��i�"Ojd����n���2t&�	u6�xt"O�qҮ�hvq1���G^0Ep�"O� Z���eP����k	%@,��d"O^K�	3)2�*�lRtF(���"O`A���4IO}�$�C3jl�a"O�Ѐb
ѥ*�����جQ	<EЕ"O�E�f���"~�z���:S�H���"Ozjc˂�)�ʱ�M�
���)�"O�	yQ��N���§N�Q���0s"Of��
   ��   y  �  -#  �-  G6  A  �M  pX  �c  Wm  �w  L�  �  h�  :�  ��  ��  2�  �  �  ��  :�  ��  ��  �  ��  D�  ��  �  O � � % X+ �1 �7 > bD �J PQ X ^^ &e �k r �x �� � V� �� g� �� � C� U�  `� u�	����Zv�B�'ld\�0BJz+�D��g�2Th���OĴa��ͬ�?Y���?��FJ%L+r|�L�ޅۄiQ-Y��+g�Ӥ��!U�6y�H��E
�I�NP1Q��	������\_Q����A�IOB("ۚ2MB�����,xmC����qI3�C�e�T寻�f��'o^��!UE� �&��f1�a��!UJ���Έ�Zv��	���R��VbmoZb3�y�I�0�������>�
�1���R�
���1���o�`�WƊ��M����?���9����?)��o,b�
#iA�\Q�I�㇋FrD�����?A��?A���?�+���;(=��BO�X���W�	�Y7�M�F��$J8i�R��yǚ�	U~�Ct�Q����'!$��5��9й�c�	�\ v��'|��%�I�3���0*��ei�5�~����r��,��ɡ�n�3tvL�I�M+���?����?1�'�?�(�X�f0�s�@?`�İ�W���KQ������n��M+�isR {��Q����UƩ��*s��Sa�
J޴�1!�>h�$���S���d^ͦ�Ra��ܟ�pAӊJ߶��!Ѯ�ug�W���T���/#�-�p N�����M,U�<{6��o��I��>���jӾ�lZ�?���Ot��R�7~dP��� �v�$S1!�
M�T���4?� ���*���釩u�:�2�cP
��x*��i�47m������I�5bÆ<K��N�dK7K�*m���)f��DMR��ܴ�&{��K��I"!��q"�&:^Z�m�G�WP�T'd�6�dpS![�x�����,��B�u��O]��E�޴:�V��"&8�ǀ�a���VG�b1L�C�O�S"qc�aYP)z:�t���rbP�iJ�-�a*[�EA��2���O���q�j�5l����
�[���"��.W�����D����џ`���?�h��_���#"*���\ѦL�i.Q��;B�ZM��b�,�'�"�'��)�y$�世	��V�x�'�wӶ�R�X�v�\a`��]-k��y���8O�0���s���zVȏ>6��� `nC�.�4�&gƞ_䘀�#�&E�����)��P�$`�{҆H(�?�Ӵi��nN&�Y�V�"ɢ���!Ѯt����ٟ��IF�ğh��˟����|���j�\���M;j�eң��R��0I�4]��]��iK.J������"W�����ioB'qӪm��d�զ���Vy�Ow��'[LQ����5kl� ��K��Lg Q�#�'��@]�t��&�_.9����&j���?q����X�̱�V+Ŭ�vd�ɉm~R�oT�}���h )#W�� &��!큅�ŗq=��ۏ(����WA��>�bP)@C���ɹ}���[��}��	a>�h��@'^�x���/�F,S&�+�O4�0��,2�3F&�trVBXɐ�E(g�of̧a=�Ƨ���nTr��p�����󟤕'k�C��'���'��W���-=rح�� \�O˨�� n��C����ٹjc!UL����O�����h≡��a�)��A؄��ĩ8Ɋ��/��1�`<�۴n��8dGY�z�-�)�f!
$䐇We�p��A�n"W����C�8r�6�gyR-\��?������|����|Ѓ�RJ�G^^�r�'Z�ɟ$��O�D ӈB�� ���ԓ:D:×P�YشFћ��|�OL�4]����Ǚ�nq����_\�ᨁB_7%�O@��O0���)g>�Ӣ�D�cRT<0QA3;��,⢡Т%g���%�ɘ%��Ҡ.{x���vbD�d8|�Q��L���)�k�t\굦�,,y
��i��lr�0D��+�8_�����mw�e� �.��`&J�OxmZ��HO�Ȳa�Ҡ8�$��AI=j�FI1 ��4�����?�01���/TpL�C��Z��O�!o��M{.O����r}��'�,��.א$B�Tl_�V��3�'��`сJ���'R��_���Ǌ��F^0t00eΙ[�Td�'��O� �S���Xn&8(Q��o�'��{w��^/ EZq'�"(���!�t$�D u.�
i2\���	!lQaDbB�)��|RB��?q��iK�7��O �I�h�w.�# �yҸ�a��<)V� ��<A���O9h�Pc�7��آ���', �鑈y�iP�i(4�'`���?����?�+T��t�p��&i&|�G��O"�y��)q�i�B�'���OordJ�'���Q� C:����=(�NQ��'m2�:8��1O��%�o���'���<RGH��@����gN=���`���<yf,�N��IC
�%d#H$����d� �׆$��i�0t��7 =	X���s���m��I {R�� �sO|���d�͞C^F��%DXBʑ���?K>����?1�O�	)�KJ�&��C�[��1p��	��?�ܴ��F�|u�����<��V 4=��`s���M�����[���I�Od���O�˓+�89��C
 	����b$@l�6� *��^Xv�� �i[ ��B�ے6�ӄ��'�n`�FCN)d|�15I�!z��b�L
�XR�D�Ǔi��Xj���&φ�auT>;P���+���ݲ �ZxK�Ke9�w�� ���Mz�*�Z�O� bP�'�1���'�r��f��Pd�#+~�`�'�N���'O��'s���>I�
�>M�ѳ�̛��́�a�Dy�&l�N�m�ݟ�ڴ�?��'��)���׊ŪM��hH�k�!t�bG�LS�"5ҳn�O��D�O�������D�O���̛g�$]�ㅅOG�D���r�b����ߕF\@�g�C�|Ś8R�(O
�����/���)�#2J��#"fR� ���� V�K�4�+��?axF�af$���W)-�hI��M��K%�r�\M���<���'���z1Jơ(�Z�� jU���B�'���'�a|Ro�
g�r��P!M�:|�Ű����Eg�v�q��ʓ}�8t�i�b�'�,D3�K�.N�	��i�(3,���'�b��.�2�'
�^5xB�8�S�֜Bⴱ�@L.s�� j�z�+U�Q�|�E�+	�԰WO۶Wɀ�����P�5Ҵ�K�/uZp�T�լW�~y:V�J;�(�s�J�@���c�xH���d���5��^u>>$�Ԍʦ	�� 9�� �4�!�Dl~�����;rfdp q� I��r��O��l\Aю Y��B�Ρ[��|+k��7��O��D�|��	]�<1��\��eAÐ4F�9� h��?�����(0"�3>���("S�[��S>e�O�&��#
'ipb���DJ6�"��������D[@�AQ���9��Pw˃к�"[Np��'d���z������f�3t�|��'�ũ��?��$;ҧ���Y"E�z��w�V����7��<��Fne�A��	խ��k@$��џ�yٴ��v�I�:j0��G����uQ��.*x�6��O����O^��O�)8l���O���O��)!ƘM����iz�!zt���ippJԭ]���lڳf�nтg+B[��*��a$DU� � b�lY�{�:�T�Y,T��c���3�F4���
XW�itE�1i�ܼS JƔ�4�iáߣUt�j�.���M��R������O�($)�O����l�0O=K�L��E�.�?����D�O��?i�O�Q�Co˸(\��c�OŚ"TA�ϟ��ɨ����<�/�N���<!vDW�L$���+�>t��r����J=`do���?I��?	�%�.�O��Dp>E2�珓K���Ū �i��Z���,@�b�ط-ƒA����ŏ
�,X�|GS*/!t%7*���p�-�8qz!�Ú�|�����o��Yӱi��XKӨX ȸ'J��a$n�"d��(S��ߕi=�tC�*���?���?��"�S&.%R��U�]�Rip����1+��B�	m�~U�G�� 97�h1���OEoZ�L�'"�Ѡ	zӘ�'
�:f�7pNp:��)81��oy�'��>�*��������h��C�Q�\D �*SV�rPT/Fx���"GjP+S��	D~����BY�"�&_#e�Z�d�M3R���a�Q<n�ޱ���_�J�@�Ck�*��Q�'hS#g,�'��Q��/���<�G�8�z���E�*(�~���a�d�l�0��%�)�����Ɍ
b�H���Od����ܦ�{���UD �H� E<�Dў�M.Oȭ�V�Q����ğ��O��rt�'ZL���(�q:u#��Wn�l���'��b�3gPr1y �>!�EK���KC 5Z�`o哺�F���PBѺ�iv�˱��'�|��Ю��T\T���Y�)/����W���Ĥ�JH	���4�hpp�F 4i��*������O��o���H���ӂib�����?X� ��-� {*��d"�S�O�����M����U�G�+b<�Z��'����a�b� ��+�3j����%)]�@^��A��^r}"�'��ݖj�݂��'u��'j�>��Ti�JܚnA�������88=�@�������aӐ� ���>wh�' i�O�`��l�:�tH�aV�,��d���Ϣa�Ґ.W����tcZ���C�q�	� � ���w�Tؒ��JJ$(��,]�{R�i��7m�OZ��a�ONc>˓�?9�"	,պ0@�ؿD!�����T��?���0?1�M����m׎� )x���eGXy�cӊ�mZX�I�?	�S@yB�^�Đ�h��hr��Eņ'6N �Y� >%+��ؕMYdb�#d��Q[3�Ï���#�wJ6qk�o�(}�,Q2�<��$EIT�F(S���3u���r��G��(�1gC�'�xJ�aB���1��"ʓp�(�8��r�y��EE�Fڀ|r��ԟ0;ߴj���Gx"�ϧ�!X"ԍQ�8!Wo��y��3��E`D�U;��cя�/��DF���'��I�V�@:�4�?!��8\`���98��X2�
�
	!8D���?��$�?����?��^�Y�&�"��?O��	�}t�qW��6<�>q�(^�y�+0Ox�Z��<e��dGӨ|(��AR`�)yG\�HO6;�=�G��
2L3�"�z�'D��a��i���M�<a�`�s0���j+�q-
G�IK�'�	��^Y����;X�<cE^�%R��������A�M�]��F�4A���̃�MK,O����צ	���� �O�Q3�'R1�G7g1���� p��v�'�B(����A�'E���Y�lK�T!�S\��B�X����1iD���&�[���ZgDi�a� ;ظU�f�8V�`���fCq>�hSܟ�h�eES������]Iiڱ0T�� Y��O�o�<�H�x�i��zg&T�?�x�І�I;i����D7�-�8!��A+h��(@�	�t��,G�dk�VhoB̧t�8" ,�D�d�E�mpP�Bߴ�?I.OY�q`����O��d�<y��]����Ƒ�]���E9~��@Y�c�m
�� �\t�8h�Y>�j���K�L�'��y����JW-L�@Ր��@�H��$؄LغB�н�H^J���u���f?�)`��H�|�8�hDe�@��
q� L�'g(��*͟�'���8E C�%���?&����'�B��6�'g�QrȈ�4M2�x4d~T$�'~���p�t�dAЦM�O ��Z>=�'摵+4�c�)+�hDǄ'@
���x�:�(�)�9��ey剝4Rn>Qs4H^���	q.�l�͂v �n�'�\��� ���F�ͥf���%���N"ĉ�#��~��T�4c�ƜK��c�'96�s�Ipl�8���g�42���?����hOJ"<��?f��"��*_N!a3�m�<�����j���pRn�q���i��#�M���čo��~J�A��~��@#Cc�a12�Yp��ٴLU0Ɓ�C�H�c��`'��2P���U�"��q��$��[��!�@\�#!���F³)+�h ���d��S��)h6l9	ү�Z�'[�$����?q�Oj�ꄀ�=���d�S.�͋��|��'(r�bJ�?�|��AG�I�9+�-��ř7�4�r�I~wU`F�'�?�)O
� �5O��}�=�=���9  Ƀ��99�zX�'#����ᜍE^��A�?5L���)�3�xYRDÀZ��]ؑ �D�x�1۞1�S%eQJ�.��	���[�M��O)���a�V� �֝qǤ҅3�\ȓ�Of�;��'���<q��7b�������k��AQmGh�<qх�q� ���U0
�r�$h�'�:�}�D�����"G��v-"93�-Y��\�	{y��Q$�p<�Oѳ#�5��AD `�p"�Bް�:b%�O������Or��|���x��H�k&���ł�%��̳�Fi�l�\�2�AKɡ�L����$���R���t�/"2N��zp���((D��O�(�)��D!�=�~	�`�ݭ^�F!�'l	H ���v4&+0m�V*+O$,Gz�O�_�4SŠB�2U�s�`\`t� �-AO����ǟ��ٟ����?A�I�I�g t�*LL0�b����l�D����\%�
���e�yf��z�����[,0x����y��H���1+�Nas�aA�n�}���M�����*V�����+�7Z���(���O:An��MC������Ox�t�K��I��h�wlځs��	�
Z��hO�'[���j�'I����@6:�l'�xܴ~�FT��G _ş����l��O�o=�i��O ��a��hL��$���>� �	�ΧGRD�E�3�4���n�;�?�*�/�d"r#C s��`r��`��2ފ,9� z!�V��iQ�Â[��q��q���RT�V"jL�0�6�\.W��"<�Պٟ<�	a~��X Ġ�2e�[zXZT�t�Q2���0>�KɾJ68�P��5�~�@Ac�N��+��� |)Bc^y_�u ���(�����QyB�շ*i�6�O(�$�|���[�<���� Y5�����2�1fȝ)�?��5���s���䓵�>y!��R�bҢ�>"Θ�CU �M~� 6K!t�K��#/U�uB �=ҧf�pG�{֍���S�� �'�s�.���I0�'���`�t*��1oC�q'A���'�ў�O]Ҝ0K�6(�H��iR�J�C��$O�qC�4�O�����^����c%:Jx�Rs�i�r�'^��=`#�(��'6��'�r>�V{�\�+�)�E�H�4��C�91a�'�}�2���Ϙ'F��aT�Ce�$j �8z��vK��y��,�2��n�g�oȽ8�&�g�>�3�:z^�|�IG~�Q��?i���hO^yq!K:|8���I)F�h�8$�2D����&ϭ_��=��E�,AR�:a��<�i>M�	lyBF�x�Ttb���8]"eñ�O�mg�(�_'%�"�'�r�'fV֝�|�	�|z�R(��pӠ�!py���-�,I�A��,>��������?X������͵�N�iB�ȁn�tt肅G~/\0�d��6�F�H��ɜ>��@�D(�f��-�-߾Y����S���O�ɟL��ҟ��?��	��0ģ���&!�(3�m��w!�$�$PE�5��7+jf]�\
+��'��6-�O�����aԴi���'�]���U�l�c�<S���J��' +2Z2�'���bƾ�!B�u�r}Kp���<x�c��64<)w�0]��!�1�'_�	�C獢H^f9c�h�;lv����7yN�u�Č� yZy��L)co@�����O^h�a�':rL�<���%�T}di	�0�\t9 �	�@������?E��k�:uF�󇂆 }[XlRaK����?!��i,y���G9N&���-|b)�`�rӲ�x��[6�i5��'d�<�.��	�L�qgV�z h��%ۀ/�T)���L�%'̮5~0��ٴW���av�i�@�dc	/� M��>f��P��X ����E��u����*tք���X99*=��ޛ:��ђ�O(`��E�*A�1[��@2\QVx#�O$�c��'|�6����A�	g���?��R"G8�V�S�Ê]�ؠ�(�d�O �D�Ox��?)���?���π45v��nL�V��Hc	��@�#�����?ɤ\?Y�'�bc��m�TP��I�	v�8�p�)�6�O|�D�O�P�4Ɨ�[ր���O<�$�O4督3��e�r�K�~��t{��Jr���;�ӝ'"��d��?p�z�Q�6�Sc�I�Lܶ�0b�A��t ��zM���I�0#,dkw�ɏgĚ���!�u�駦M��hS��y� �H� MS�Gɶ���]�S���h�'��I:E���d�O��=�6��s�� �H:K���{C�L�yR�M�7����� 2�6�x�E[����a���T�'v�ISi�ȒC��!�"��n�P�&n��]h$=��П��	џ(�\w��']beТm�X򵮛�08��_�6A���ȿh��Ep���7$���K����r�V�c��(귏�V�,(�E�-(�K%lG;L�b��F��
0�dG{�mF�L�H�a� ��u,|Ƞl\�x�����b
@�rx�S�����$�"E��S/�'�ޠBF�Z:?�ў���C7?����Ɉ�D��0$���n3t,O����Ϧq��Fy�O�,O�|�'�?au`A �hPfȤ2��R�! ��?���4xR��?y�OPp�rr��/"T����oh��I�'a<�L�"oRbzM�Ņ'B�џ��p�G�~iVq0�M�'���u�l� ��S��u"v��V&>� �E{Ӹ}�ǆ�t���%�`��f�O���"?i�1Zs5K�־d�s��S�\������=t2;R�K/#��ũs)�One�I�G��c��C�b��dӯ+Ŭ�Ĩ<��O�j����'nb_>��s+�֟HiaD��y�Q)�J٣c�T8���Rퟬ�	Q�L�;VK�^/�A;2�Σ V�PL�>W��<�O�̙*�!�-�����[�.rzĻv��<�4�Ϸ5}:l�VH�i��|����9O?��R3�~���O*��TQ��ЀG[���F�E~��O��?�ԝ|�𩄁\�]@^2�DJ �09�][�'��8��b��I!<��v)T�9�������t�O;B��ޢ5���3QN�-E��C��iw��'n���g*��'fb�'Hb8�-� G� �)a�V0�9ՋԊm� +B�֪+yf� �Đt��S�|�&,�ɂ"�]SCIJ������% ? �� GS��n�#	L=����-�
�p\r��ON�שN���!S��Jf h���$�$Jf$����A[��;�lH92�H���X�!�䜦CTXE䊪"H��G�/���.�HO�))�D�%W)��Ю[N�)\(*��={i�<�C�O6���Ol�D�ºc��?��O�20�$�62��1�m�Mp�H�PN�V�UZP�ۅ1�P���)9�Ȑ;���~�'�]zcm�7��k���s�� rW�� r�T 	��M+d;RAd��Cz��d��K�'т� �B�-,� ��W�^^<�Ӈׅ�?���'9���,ȝ6$-Y���#zd�!
�'T�r"�%�pYӀ)l9P��L>�$�i��'��{TI�~�`db1��.����J�R��Y���?��D�(�?A���4dL#�	��N�f�
�� �iIJ�� ���~WQ�tc=[n�m�@�iy��F{�.Z"�t��҆���n�Q!d��ʤ��ϬX�y0�+,�A�&A*X��|���՞o�B�'j���J����(V4)  ��剪Jn�O���E0L��ˇ%��X옢�I-w���@�O yC���
Sʈ�'X/,����'��I�r��O��O(�'4;�E���E0�|�� Q-N�	�"9SlIA��?���FN�PÒ�vQ~��&GbH�i� Ĕ���)K�{�*��4g[?{(0�f+ٷ/���"Id$�/۫����8�����CF�l�j�ҟ�l��#Ǝ���e�I�:��v�� �5/�O��8�'�y��#c.<<!fL�6*�t�K����y�����O�/�y�d�H���O�E�D��6xh��j&.�$�R]�� 4ś�'�b�'U�̰�@0k�R�')R�'��N� }�X ���U?�<���ϕr����OHh}���
Qr3���y���.
�EJ %
��V���L�X�Lث#N�>YE�	-
Rx�|�<Ib�_��F�`�	(p�:�l�����';V����?9��$��M �kJe�x����}�FC�ɦ#
0��4�	)XZ$��ՆU�N>i�'��"=ͧ�?�-O�lI�KV%F�I�`Q�9�(Ś�`��-�h����OX���O���C���?1�Op��R�X"K��<��!H�U�tu��l�*l�T�ʇ��Yk^$ۇ
Y�^�џ�K��*U��0��ƨ]�7�� �S 3=�P��監H'L�`��.�aq�.[������%?�a1шQ9���$�Of��;��I�O���T,K�o��G=P����
�'���34jK'<a�`!rnġ� 	)M>م�i2�[���E�*��'[�>�����3@�`���%���t�IKy��'���'=�
`�]*H�����I���d����x'Ä)�H���0T{ax��˦-I��Q$�C$B^���'<v�'�X�f��AX�M[�jH�h�
Ó
�Ҵ�IƟ��'tc%��
.�1y��=R�*]�J>a�B�͋ǣ�Q�a��:O������?yq
X({���c#�1T1>��G�ϟ�'מ=y�_������O@����W�q�|�!$+�z!�O��dʣ.6P�����Zz,�6��"|�fA5�ViC1L�1�P��h�S~�����L�%MՔ�������+X�xy�a��!��Ѹ����^bD�@x-����@D�2O� ��Z.U�X�X���\3��mq"O������3��I7f~������h�&� ���5:Xa�-�I�:��'��%��4�Q���e�,0M��e�$I�1�A�6D��	��E9N�l� 	4b#�x�8D� Z����f�>�椕>3��3�a8D��[��Q�`�c@G6����G�5D�|�&���"nP��р�*]�vIc-4D�\�AJ�'U�
F�� <ݠ%c�<����j8�@��' �%{^�g���*���%D�4P	!l%{Q�y�ڽ�G�6D���RB�7�j}J砟');����G?D��p���a��Z BvH)K"D�0@��.hht���R�I@Xkp�<�O�����O^�rӇ�� { (��
	�-mR�K3"O803��ظUdx�sʍ�|�9�"O�;����J��b*��7���"O�m�B'^	`�����#�G��\2"O��� �W6j���4?�ʭ��"OU�c@�c!�� E��B�2�AV�9*��~� ���|ڳH�.>� �U��Y�<!a��b�x�#��,tNƨxa��T�<���ǥ`���q��P&+=*h�tHS�<����.�B!ƥC�
yU�HI�<Y�a��HYP-E)c�p!ȟA�<)�ˆ�vx�����#�� 0��JҟD�ph7�S�O��=P�(�0Q�"�xA� ]vya"O>9C���`��9!t#�.����"O��֯Z^��y')P�sڲ��f"Ox)���U�v��$22�ؐ�p"OT�!��
�ZuVU�Uf� H���"SOرZӁ�$(x�4!Qo�c ��a(+0��q���O�|�Ōa��Ba4w�䈗6N�p��#��B-��a�>gr���,_���O�[�N�nO`�K���DHaJ�.���K4뙊y�,��1�2Y�BTV�'ٸ��i�fB\� һ�X�a�{ݍ,=�r�'	@
Ff�	RSD˪'���,*���'1��pbm�E�L�H��/"���^���I�)+�8�5�E�OMV��GHE ~B�����yb
�?,:�:@I�Y�> ���D���dE9|B��O��?�'Jai&dZ	0�a�'�M�L���'xEI�gMd��Bc<{x�� բ7ҧE扪R�;�"$K��	H&ҽϓ�J�+��g���7哢($-ӱ�S~k^��N�)�J�s$� =��牋 �����O�S�{~�i>܉p�Fڇ<�T�g�ʙ�y"iX�J�P!��~�������hOt�E�D���*nT�z�`L�ک�cN$+Q�S��#�%\Oj����HG ���g �<@:(@���{Oܜ)��՟Rظ��b�
]�����'���	��W4r�j�	#[%y h���b���j���^n�)����ɚV�pb�,p�~��!�e��\�� �'��%k��?Q��o��R�V7�4]ۢ\6��p�&.D�Tٖ$A4X������X&jT�AY6��O�Dz�OkrY����Cӭɸ�ҶI>��z��˱	����3�\%�E�)�\�k��/h��ś�'W?�~	� n�$��H�E�����OzD f��a$Ҹ{�L�>x76�K�J�o�<=`$遳>� 92$�Φ't�F~����?�F�ƃ)��9�S�4�z ��
.�?ɉ�d%�=�.1�T&c�*5h�N�)��\�ȓC����մAj6e`��E�{�x��',�6�OHʓ3���S�'%����&�^V��4�@�E�8E|�Aۊb�xY��l4rb�Qn�%�ם0)�D��Ⱦ4Z�bKh�#>1��N�2��"�A��s������C�J�NO�b���v��;�Q�AEM�#���TL�O�d(�S	
�Z�0Rdɇm2L��	�3��˓�0?Q��_�XĲ�e�]ÔT�&�Epx��)O�X0�bڍ��	����-H��)iqY� `�d����q�g�$^  P=!���i�Р(�H�%��xA �������X�Һy��(����޸O�i8����j��(�&'�&ZT��'�6��ɂ:[b��a�X 6�н��MәP�.��}��#�	8�@iH����0`���!Z�<���Ο���.O�O��3� U��IY>p�b��dl�%t�`�b�"Oδ'��&�B�"�$��y�%�I+�ȟf�cR�
O��Zu��0*Ab�(��O�˓r<܈��I'h��KeÔ�9"�A�W�E�(�d��D�aC���sc��+���CD#��ʩ���'@h`���
<n=Re�F�U�H�R��_�|\����[0n,"v������}ò`)O�T�uI��!8�Ys��O8ur���0A�Uy����?��iY�3�Di�5. <��`�
q\n  S�'D�80SIW,,�N�B)G8P$@AO�O�8Ez�O��V��1g��.H��p��2��x� !#ݸt���Y(h��d��M>N`qF�E���J'M�o�����F��mn`X_��E~�V �1i1Ƙ7;�� �J<T�,�f.��1� ��p�b
V/�p��x�ɚXhz!���;�LQт�^�K�\���x�'��da%Ê43��b��;�V1�h"D�����N��R��%��Xg�<��i&bR��X��ԩ�M��?ɛO��Ͳ%⍺9.z��^7�ѩ�q�ް{��?��"�(q���� _n)3�R7��V4����夗ޔ X!xg���F�ɣi�rL����9�p9CH��!ڂ�"���1D0)��O-	A"L�O�"����f=�S���������N|:砂�;���L�8U�|�dT��?Q��������)������b����;�O�oڼ�M�5��9'�^\�`�"*�9y�*���d�O����Oj���O�'���� *(D��"U�DX���LA'��d?*F�Ԙ�哌}J-�!�H7?Z޽� V�R�n �?�W�r�I�v��_?�[R���K���	��{_��y� ���M;��9���[�'�@�2R?�����͓G�`�tc�?Q��hR���t�B����MS��g*�]���yҁ������ڟ(�"?�\��,6
�ɕ�<0�s�'�B�@t��bݡ�OA���'�$�n��� 2`�+���净sa,��6�'VbdY-_26O��8�ߟ�^w��͓xG���5��lGP@�0�� %��A�Z����I�� ���?�]w�S�?��S*XD̣�l��8�J�� ��N�R��)������D�X��ě�:�Jq����ܼ)�t4� w�hp�%W3{w��ݴ�yB���?��^�`��OO�S�?-�C,�i�Z� ��� ��I8��B�i�	����џ-Ga���p�14o��?�n�i�(�;�k� �2M�Ðg���p����Ms�'#�a����?�5F ��E�T��*Y�y����y: q�`X|�r6�4(5��#�\n�?�MS�'�?���'�4�S��/��a��-?�2����Q�_z��z�iah��'�剎��4?���_���]Mݢ���5��)��A�>� ��T��(-����f� 9\I
e�IѦ}��Fy�'@��'%R�'��'x��#�ܬg��P���7)kԁ�s����O�ʓ����O�$�O��$��B�+�ƇR%r�T�+,yl�����I�h�	��T�����'��X�V��A�̄�jN���ϊ(�l7m�O��$�O����O��D�<����~��]�b��	B�q��D��̙���=<O8˓?����tm�8M�x-+��T�B*TX:B�Iퟠ�?�u-��j���`%������!�&'���A�ꨟ�%�R�݇ ����&l:V��"O�my�E �~yX�(qk��(N�f"O|Sf�����)��dԕe"O��򤣆2Yw�4���Q{&���"O���ƣ��[L�� �(�*8Uh4"O��)!K"B�8���ѸK/��.�������l���`��Y��R����4BXzO��ٴ�?����?1��?	���?y���?��G��\���l�@Xa��ԕ}")���i��'0��':��'���'���'�����&�8�P�s�X�a���Jc�����O����O0�d�O����On���O*$�쓍'�B5a��Z)H����(������D���0������I�I�|�1�'T����M���(ƣ��M��?��?���?���?����?��ڎ�R0ǂ����J�-B����'���'O��']��'IB�'��W�Z)�0�e�9_�(�QAF�".o�7��O����OD�$�O���O>���O0���@N���e,]����� ��)4Mo�ܟ4�Iҟ��Iݟ8��̟��Iҟ��I"8
�աËԷ<DƐ�gK��^0��4�?����?)���?���?���?��2t|�+q� ��-{}+&t��i.��'H��'�2�'2R�'�"�'n�b�\%.\2�!�\':hh�
z�(�$�O����Ol�$�O����OH�d�O��'#)`dL(�GLpIQ/�� 7M�OF���O��$�O����O����O��)%��� ��ח
2�YB	 eO�,n�i~��'��L�Oj0�)�劣6 ��3݃kk2�˅�iվ�P�y��O��O!Z6-q�uҕ��WJ������P�DX�Q	�tn��<�*O�O�^���~b咇{-�3�a�N/���A��?a�B�I
-��"M��hO�i~�$�qƟ�/���S�ŉY<n$ر��O����g�����'�� ��)dT,2��K�`��k%��@�d�My�'���1Oh�~t`�ǫN���x���"��'c8����U�o��P�O�	�UD���
d���ƃXf�\|��
���I�<y)O���"�g?��Բjk��B���Z �w
���ܴ,T��']l7m?�i>�H�;ʄ�r�߿F�.�(�$��<I��MS�	E�a{Q'Pk~�o5���캣rIU���ࢅZ5���X�M[�'mBZ�P�|�R��ae:U"�#��~-�BIPyR�`�,0��2���h{�ui"�ţ_׬i�ת�;�0��,O|�����Ie�O������1$����H	M�ؐ"�E%`�{�O1W%�/6��%�H'?%�M�o�F?�!���RM��ڳ@� X$���.���%�'D5Un��"`9�O����E��?	����V31��#���22���.ʞQ,̊c���h@��cB�<_���	Qdԋ<�T!��g>^R�mǪUn�hS�H,�d�Ѧb�;C��|�6gّ�`�`�[F��TJ��q\ĭ�kS��V�#k�,@xU�u%�s[*���E=X���b�=HL �k�$���Z��e��*r�c���lY*i+�̎�?&��2	��`!���F�x���. �hx
 /+�<P�Ã�z�Yc���*�b>Td*��ɍ�lT��n�'1Ψ!&���	�FMd�y#�N�2<�	�!�	B���ɔ�ğ9�҄����=����Z�Rw�04��(S��܁�͙	@l�Ŋ5F8wo�X�V	�6�dI���W�n�ӷ��2g�|�[���F#�zs��b�=$����-+F�K�&�#�Q���&vM6�xѥ#HA��
60D�mnZ՟t�� N�H�#��#bB�X�6*�`����|��ş��'��*H71O&�S�Ō����B����ZS�'�b�'*b�'�>H"gbe�0�D�O��������@JP�r<N�{G�A�+/�	�I�O��<���vZ���'���|d#��,�
�뇼u*��'�[��?���?qdJϿ����'P��'����O�b*C�`���r&�	�hc�D�hw�ٟG�����I؟dr0�}>��O$l��'G���j��V**�����g�i"B�'SB�O�4�'R��'e
E��^����k �y�T����'hR�*��'�R�'���H�O��O��OۘP��	�q��y�����\d�7m�O����O�Kb����$�OJ�D�O�d�$N��E�KS'�X� SF�Q�4����F��i>U����P�	�J�ıٳj�{����a
1u���	ٟ��C�A��M+���?i���?)U?��:��9z2��*tI�)�傔�4y�'G���'Q�	��I@��矨ӢMU�!���ϟ$^�pRDH�H��4�?���?���:@�Py�'��<znA;l��!B�Ԏ��<��ȗ����O`���O\���On���2�mZ8t��I�d��08���8�,%X�d��	�,��џ�	ڟl�'G�)���$EK>BNN�ȓ�˲;��v %*e��'�B�@4�'(BV>�k1Đ��M3��?1�&��.9��T�\)z�,1ɔb^��?���?�����O�X��=���kQܸR�Oݫ|�q��+1YI2��I����I���	5-&�I�4�?����?A�'_c|�Cw���`�a%"<���?�(O��d�(A��I�O8��|�%�Q��n�0���:�P{!T��?���?9s��6*���'(��'[���O��m�S#Bá��1H�( *ҷEp���L�������Hy�O��
ހ�e
B"I����ԁ�-�D`�X)nџ������?��П�ɕ���$��<s5:��W��kE:�I1~����	ɟt���$����'Q�aa"��U:��7#�.E�|D���}�~�D�Ov���,3�����O��D�O��D�O~H)���z���5����# �<�-O��@����SڟT�	ϟDPBN��J-R�@���N5�01b������B�� �ܴ�?����?1�����<Y�D�A��h�(ӌ��@��Iy���y"S��	Ο��O%2BȨ5?�b���['+��a��Z�c����'���'�r��~r)O|�����!��= ��2ƌ��(g@�cv:O����ObDq�	�O����O���ͦl���o�09~���B۰;,P �D� �������$�Iȟ��̟��' ��	���BW���%�b�W-%�|96j�HPb�'���'�U>)�!�H<�M���?�4��V7j]K�h�V~MP�*E7�?i���?������O��F3� �k����O� p����fʞ%``���ҁ�O���O��$�O�kOথ������I�?	��4}��+wWGǊ�c�@�ȟD�IAy"�'��Oɧ���D���r�I��[[\	',ı]�r�'��CČw2D6��O~�$�O�I��z�$�� B<-#3�>мh���0#0�ʓ�?pA_��?���?�r`��|�̟����#|&0��HE�V������'���gb�z�d�O��$�<���O����O��� =������u�"�(S�O�	����O:�d�<ͧ�䧬?����~_�dpHT�M��)�u��b���'&2�'��,��O��'���'-��L�qn��I���2r��&��rEr�'��P�Fq@��U����O!"�'o��ZV,_�X4�)00��Xy��s0�'���I{V6�O����O��d�J��1O
�A
�.rK�| ���(�*$P��8�m�����`�Iܟ�&?�SV��<.��s��J��Ѫ1L�!#��,h�4�?���?9���Swyb�'��)E+�dd�1�RR]*U.��y�'���'���'`��V5�ٴZ$"�(EM8h�;Ul�lt�����?���?����?a-O���P�_b�I��~���
�'�DX�P%¼J�"���O����O���|�Y@�SV�i��'4�\�E���U<�{�@
��4� �'���'�P����:�"���]1QR�
+O n���hH�������������
8F
�Iش�?A��?y�' �8;#�>K���S�G$5���[��'0�V���I2^LŔ'��i>��.�K��$���[�V$��2qB�����	@
1�؃�MC���?������?)�9�xE��ڲ^X9��/�����O~P����O��D�<ͧ��I"�~,��nY�=|����h#m"jn#�7M�O�$�O<�i����$�O ��_`��S@C�?Eܪ��B�.Z����o���<�')��|L~��� ̡���� G_@�Q'�Z���u�i8b�'2�H�pO���'p��'���'8F�ɐ�#~e���UΓV"H��'�'��<����'���'��!J����y���=3����'R/߂p��7M�O��d�O(��w�43Or�
$�ߧ1XP1�A�ɫ9�%�'���D/'�yb�'0��O�2�'��'�uۦ�L/ t����@C7HX$��'��jr�6��O����O:�D�Y�$P�p�	`t(���D�4מA.iԬA¦�F�k��d�O"�����B�d�O�˓R�l���O��r B�5�d@�@���z��(O��D�OR�O�ʓ%xm�,�^�KE�AK��)�����%���'B�'�V���L�8��'r�LX{e��f��9�*�0H�����?aO>�+O��B��؉l�:�`��%���SFBW#2�'�]�$z����'�?)��u�F���^,�`�&�'`�,SO>	.O0�&�?�!�I9
"��bP�Jn.����O�ʓ�āI��in�ğ��S����εPc���B�&�����T	�"V���:�SܧTARXgi�w� �W�G�rP���I�E�J�kߴ�?a��?����'}��wr�@��!�P܈1J�,i�"W��O>���a��@�bDyz��q�dϭG��Y
�4�?���?�U�</'f��'~�$��H>�9�%��^$��f�/-��O����d�O$�$�O~КS�@�w$`my�%W�Y�i���O
��W\W�&��	ϟD%�P�.�+{XL�S�&�X7V��s$�ry�C��'�B�'zr[���f�d6�5��F���s,\qR�zH<���?�L>�/Ot��h��a*�a���öB����聠g�1O���O����<�aݣs��$�?~<���7!�6`�,�7o���?�N>�/O��q��O~a"@��+2�u:�MXW��ѓ]�P������	vy�ˑ�1��.���BJ������W�T�H���O,��?���<	3n\e�i1⅀��#Y��ܑ�Z�~��4��͟���]y�
���&�`�������^%W� �Y��̸=����e"�Ĭ<ɣ�`���4	�$uҔ���� �¥�Q�L��?�(OJq�tƐ�-�O��ON��I�R,�0�"�ZuT�͙Y��By����Oq���Yţ��!�Od*��V�'�~ͱ�i����Ol�D�.8%����+O�1+�$�.=�l����"�5d��#<E���'��X9#j�s?�e��'T%]����Om�����O��$Yf�n��>I���y���V�N�p��D< 
B1��l���'+�9Ïy��'��'��q"$V$?�Jm#NɇC%��(��'C҆�6*�b����B�%�t�rh��_N�4����)@���'# !c�y�'?��'��I�#k\��L�b����ƚnS���Á�'��'2�|�V��X�"I�ꞥ24�̪ν���Y�b���I͟4�	jy2!@2�b��Z;+�� �N�n��r �29��'-�|�^�4�Cc�����H��:�$1��DD1��q�5N�<y���?Q�����U=E@�)$>��t�W6��`�f2��K �Vٟ��IT�	Yy�	N޸'1�htk��A�v��'lT.s�<����?������
���&>����?�BɆ)0��"�Ǜ7z��1cǤ�̟h�'��ɫQa��g~�O~�REi�
���M.^�na�G�'�剿-�d�ݴ��i�O����my�FD9�YS֌к-QĜ��K��?�+O��kу>�i>�'��T����b �Å�"&*(���.�$���iHR�'0�O=�b���c.9��dR��� dH��m���+F��|�<��(j-ࡪ9<��0X���Ax��i2�'2	'��O8�d�O��I�KE�s&��h�X钳)C-ܺ��d�O��D�O�]��	C�d��ƣ�c*�ش��O6��	Z2�`$�d�I�%�`0W�
�޽x���<@�S��Bs�'g��'�2^���'b��ԛeH�8��D�� ώS�FP9N<����?�K>��OT�T��O4� �d�� ��	6�D�O"�D�Ojʓx�<[��O��-(�\%�0X�"�d�.�+-O �d�OГO"<Ʉa��,��uZ�B
�ay��" ��dy��'�r�'��I(i]�@N|ra鏤v����3]x�4bV�X��?i�����0<��B�]V^�S�(t&LP��Rߟ���񟄖'aPpa2.7�	�O��i�Q*���%D[Q��@�M�>�O�����&Y*r柶yuƅ�g�/mB�X� �e��Mk+�������U�'����fmH�c��ŋ#CK(i������x�boJ�(JZ\mD�(ǀ�%�?ɧCZw��F�'��'e�d4�Iy�? �	��1MD��ɔΎ8p�0��'�RGܵ0��\%�[&*�Ay��Q���7��O���O�mӔ��x쓱?q�'��[�P�9q�թW�J�:2��y
ߓ�?q���?Q�/&?t�2�'΋��}�w�&�?��M)�xF�x��'�|�G��DJx�"g�Ŵ��m O�p�џ��	��I|yb�ٚP(�w��"8n�qL֒s2q(��"��O��7��8?A��ݾT��ٹ M��M�aP�"�N��?����?�+O��rg��?i���̪k�.xboM�w��{��<����?�K>���ā�=u������;�	��eH
Oj����	ڟ��'�z�*0=���AYE�c�T�1��DqQ��I��&����J�h�CED$+%"B��N���$�O ��<!�b\0.��O��O�j�J�/g�Ny(� �t�h����|��'����B��1U7�ԁ�\�:.�������݇KKZ�l�b���'s�TF�<i�FF�(��L�2�<vi�� ��
��@���M+�\H������`�VڰD�	
nX�E�4�?���?��� �'�B#6�B�Ӷ" 	GڞJ��"\���'���!X�i�b��=8B�2Sia��d�OX�d=eh� $�������͓���T`�80�N���g��6�T9���؟��	���ČI�M�Ó�P>j�0�b[�\�I���K<���?�����$ґNϸ(Zd%�
\]�MYFo�m^\��\��<���?�����X�J���F��pEc�E�[���A֪�Z�I��I󟌕'�"�'ľ�:5%͏Qt6M�c��U�$�Gf�Ƙ'���'aRW���G�_�|c����z5�OR1#\�y#ƔUy��'��|�P�T[��<	��#1]L��Q��#:�	#�JPy�'��'@�	)ʹ<&?1��		�Ov:�:s$�8M��� &H�� ��l�	vy��(�1O����̓.U��QG�:yV�F�'��'q�I|Һ��L|������Z����,�-6n�}�����䓶?��V�̩���SU��=l|��"�=[nҖ�����''`0D'{�N�'�?��'F��	�UX���f���2���L͠1JT�d�O��$�����>��l�fO	3�I�W�����`�Oĕ��I����ҟ����?�N<Q��2����Q9���3�'���'�Z�b2�'yɧ���dL�̢dS�ʐ��+5�؈A���l�ǟ\������TOT����?����y��÷
�	{��Wb��*ա�*�?!I>�"'�:��'�?���?� W$"8���"��v@�$D���?9�Z����xR�'�R�|BdEI�rѩG�_<� T�1�2uK��'�t)�A�'��	��	�@�'\,�p]c,:�а�߸A�H*SbN�A@���}��'����L�Iҟ0C����܂|+��O2帴��&R�' �`�'�R�'��]����S7���@�~*<�ǖ���C�;?i���?�K>a��?�����?��J
D�Z��E޾ry�]BS�����O���O˓[��k���Ĩ�A�Ԫӈ/C���s+*8��'��� �Iȟ\�#�W`��'C�0BLV���Q�3��*�j�����?A����%R'>]�	�?E邉�>vv*�
��������F�I���$p�����n�?Q[��Fp�Py�NT,���۲��On�`�\�;C�i��؟�ӧ���X\꜄�p��;*��*u������'F�̱HU�Oq�Pu��'�U��E+'��|Qx��'[
h(UfӘ��O����:�'�����M��A�6f�����6IR� �j��I�b2$�Il�)�'�?dg�7�Z}��$GS-�#�Z0Pu�V�'�'�Ҙz��.���OB�i���5N�!8����c���m���O�O�$���&���Od�$�O� Qs��Lb� XUl%k�xҰ��O���n�&\�>�����c��p�w���H�h�����M��?���T�¨�N>����?�����$	�l;t$���ۍ18����3�rUC�r�Ο���t��Ο��	5J��}�U�F�aj�BŧA��bw)ǟ�'BB�'T�W��2�n����on���C�B� 8��[>4˓�?a����?i�d�.%���$���	�C]�S�9q��X��L<a�.1 ��q��0-f�SuK��.�As���y�8M�AD5*�`ɗE�y������]�8W2�'���' �	�~������D�	�|bֈ��<(4��@Į��XCQe�՟�%�X�	Ӧ�ӆ�?���?i�w�Ȩ�G�FZ�)���.kR�O>���i^m��Ǆa�����nb2Y�S�FetX���M	� �*0��j�^}�1�>�� (�-8�`��=(�)�yӎ�/~�q�Kߒ2���h��B��ŢG;X��ǌ�>R(��>���OH"��s�K��������7I�a�CY=��x���L+YC���
Ԥ,B(�b���'x��r����hዱ"�)3Rp�A A�mZ�[Rۺ:����d@�0�(cE�R�=��t U
a�`b��9\ �{B��Fx}�Q�G�n+dxbV޷+X"Y��F�8,�@��禭� )<�izB�ͦs��ݣ%�a�?���/����ژ��Y�L����#F�l< ��	�1k�n=�� v�b?Q�1�T	r.b� �B4���E8��A"�+��� ��X���#:��%��3;�)�3"O��H���, :�zwd�w�����'�L�<���΄Ͳ�ِn2|��A���9�6��OR���O�@K�[�f����O��d�O�)\�Ѐ'��OGH�"�g�'ZP,H�A��H���ɼu>6N^�g�	�8�-L,�"��$B]8=aBӜ��i!�ޭp6�!�CY���O�$ ҅w�!�)�C�$��Ͻ7*�D!i�l��'-�D�S�g�I�3Aԩ3`�V�V��\ۢ��.=RC�	=9�>P��'A@)����*�F�0�'�#=�'��2~�����\͓
��'�H�p�%fI��k�B��?���?���x��n�O��n>9���;�:���Α�%�&c�� 햽3�J�,��	:!ɋ)Q;��G�*ŜgK��Sg�ͺqU�8�#m�8of}Ȇ#��x!~x��C����ѱi����VH�ָ'Lz���L�_W�(�_�H0�[!���?�
�VI�5K6�� H-���1�A�q��-��y"�%���A]�I�P���q@	�=Q7�ip�'H�4 O�>�۴iI����l b�����SLD�V�'�R���'U¬U8T� U��� w$��еCU�W�j���e�'z`����șJ�JȄ�	x��ʀCF�]���4A���#�L�
��Qr�O�!��X`l�&�.t��V%�b�p�O�O���C��nڗ L�l��"K�_��Y7�ļhE�}I*Ol���Or��<���?���M�шL?��Y[�I]4=�<��T(<I����A��Q3�C�DA�ł�3֒j԰iB�t��pX�b����Iɟ�	�?�`���H�b� � �j�ոD�s�J��?��>��=Z`	� ��1���*���D��ds0eDSr�I���ɭ0�%�DW?/J�3����(�r��Hi0�Ҳ�E0v��9'��M����^��qGJY�\��x򃏔�?ԗ|��$D[
�`t3�	�00\���D��y,����0i>*wQ�u)^8�p<I���I��J�$�?��%���r�I@TP���I�ؠ�ᆃk�~��ܟT��ɟ��ܴ �@3o����%H��@:���"�������RL�H� �t�'��	\~
!s��a
}��I�u�񸆡T���8���>JHV�aY��O,V`�Aw�Y9�I_7$�R�Pa)�OH�(T���[�����<Arb��S�?��>	#G�
���$Q ,�N�*#jRm�<�j���`�(Fa]'Idn}��&h�dE�����>�#K�+l�2LT,��LT(�ehC�8���"�C���'���'�0����I�|D��/���p���<$����3]�H����"�;�I�&}D}Ru.AS�zt3�`<�I��Q��^�\�r�	޿_X�a�IO؟���"	�?�h����G�M���&D�����I<�<���F�L�4�%�ɵ�M�L>��"�f���'b���NⅢ�͎x(�㗢]��@�$�O�{`��O��h>��e��O<O4A0P�)qP
�_��5��'�É}r����VFJ�3����D`��<���՟�K�8[�'J=�L%����i�j�f!D��3a!���H`���8Q���Xdn>�dK�N��:K�𲣟#Pۀ���M�M>���\-���'I�T>��c���1D�M�-��|I��PDZ ��?���m�H(�����Y��I�`G�Jr�N�*��8f$6�Ucb�b?�`'$á G�����,6��z9�XhR+,���� ���@qJV����p�H&_�!�Ĉ���A1�D�L�[0�¢ :�x�*'�u��R��K�7m���a���B��s'Ai�b���OT���+g��	���O����O���w���s�c��_?�I�ӥ�+�l:�k>�I�tB��$D�b<�����+e���a�P�O��O�dP��' <;U,oX\hLS |�qb�s�~����x�듎R(�Ӵ�
�:t$������yR,$|�e�W�. zi�K�����HO�7���EU��c��BD��CǑW�>=���C rV$0�Iܟ���ן�kYw��' �)�=*�� %�R?�L��D؄g��4#�O�}�UJC�l��x�EK�F���R��2j�!�CV^Бj`�R=~� ,��A��n�b��'3*����%l��e��J��"	 ,1�!�D2�6�����a&А���0�qO��nZM�I"�Dcݴ�?��4gT��0�F�XP�M��a��'�2s6�'c���Y��'�)��n�R�xB�H�Q9 ��v��lqB��1���۰<��kGN�Kc~��F�	�.Zly3�����T݆��]���.�ė�
q��ȶꕎ!�ʱY�͐D�!�� 8�H�#��:�0(sq��(|r�,��
O���!��(4�MJ�%:0ڝ���b�OP0���Mڦ)�����OB� 3�i"�#��^�\e��0x�B<x'��O���%��$�|�'F
ɒ��.-!ʳN�$}�P�xN<)��{���OѤ,�'��w%`qӆW;@d�QXN<����������	n�'#���Q�Б�*9y�]#8A�y�=�����<�q-)�H`10-�Ng�����x8��َ򤞱'�U���
B�ii��_�EQ~1sٴ�?A���?�$`Z=��	���?����?�^c1�ȳ�$
��M�a�F����d�U�,)���'��� ү����(�Z%��/��E��u���C�A�dȃ�++��,#�_�6�z,:�M�~�'/����B9O�DZ��W�t�vM�4a�X�.P!%�N�M4�iW"@�����,O7m��T����iŰ'� =2l 
��E�I\��h���rs�@=`�ޥ*r�S*OL��;>�"�io7�?�DQ�p�P�)�>���#E�P��T͚�	�D�k#׮A�L)J \ H���'���'�R����H���|
W.K�)Y��R�Ĉ]�H+�kAW�j���
6L�hq�C�0��PP��O�M���O�V<Q1�O��� A-X�q��qj�E��JP�	f؟����R��^�V�Х �4H��C�		bl���$�"�ΐ�'a��V�n�h�4��sXx����i�"�iRD�K�OM|�8��2B��'/�T�!�O����.%,���O��d�F��H�� NT��J�m����g�-H���P�nə&�2]� TG�'��Y�AE͡GR���KOjtpBW��=��(��*�>e�J$QV:thA�0���+�x`�O�I���w<"`����I*�hpr�U�������k����?�����OP�!�脄H�)����'K9�}��'�ڹY���ӵ<$@1�ԏ߸`�>���/\� u�	T��M�.OJI`S������Ouf�)%�i{�\�t�U0e�:�zG&�-�ڳ'�O���Q;@
�D>�|�' ���g��4�튶Ć�Bu�IL<���T���O4��q��L�p���fo� =Rp�L<�%��ɟD�<�~����2#4��F.��	e�`�<qD�9z��'�W� �J%�tǇ^8���$V�nW$q#��($�å+�V�da�޴�?���?� IN�vLP]R��?q��?�]-=����)�6!V0���%ά˜���x�'�`J\�����L>�#+
�,=a� �f�0"��K)�p\)b�R�"�ֈm�za^�x��L<1q�D:/X��#��Ys��F�� �N6���1�ɘ��)�)�<A۴7�X�#-D]���["@7s<���Q�|F{���=<�Bt�1�ږ%�`�!��	���
�M�ǶiH�'���O0��w"R؁#CH0�м ��V�^	���G�z�q��?����?Q3����$�O��S*d�8p֣��Mt&jpH�"8��4�wx	y��ި'�
��d�!2�p��g�q���yS`ǭiw�Z���"Zg`qp�̈ rv��3E����5���&�j�9�
�n������O��nڶ�M����D�O�c���ߚp|���j	�S���QF#D�t�7�ж1��ņ�^|bPI�` �	�A� �	]y�,W�fXם���nځ[����&��}�C�ן\?�x��?�w�?���������?�K<)�*���r� V�S�$�*�#tX���*:��!%9�XP�
S�B	��/�KW���d�8
r�?}��֛=�>  �!F�T��-���R:�y��Cx%\e�P B�7p�s��dH<	'�'8�D,!��!0��b��T)�x�K>1�mY+X(���'��W>Ugi�ަ����!����##
Z H��diK��?�4u,�@��|��� ri�8�0�p�R`i�!����a�6`��Eub��N�7�ap$�xB��<oı��NN��������EHc`�8�@��S�$�ْ2���gU�+s�Q7=��O��'[<�O��V1�2Jh�#�E�|��b"O����]$)�F�}l��� �'Ө�<�"87Y�y�W >~���b"D2j:�7m�O����O U��k����O���OǊG�TZ�؉�G'm}~��&�_�|��lI�ᇆ1���^�]^4�Ī'��H��� y�41�֋,7!@䒂lǝNI:���[Y�8�{�$H�3���qw�I���O�6��ɼ�4lZ�l�4��fܐJ��J���OҀJ�����ē{Y|i�eNQ�&HQ���-c.���i.��dmJY��R�կL���O��Ez�O��'� �I0)�L�1,�����y��)<t`	��B�O���O^��
޺���?A�O�.8r�&5g����so���i	�DJ���e�������#p�џ�d��:!�p�Ó�M�	{��V���6-��NY0V0�賅ۥT!��D���w������R̨XSfS��r������F�j���d�<���'L��f�['Fa¬˅kwZ����� ����*��̝���E K�����dJ�_N���<A� ��3h��Od7M�-kL���,Y�Py"���T����ܟL�d
�ן��I�|���-H���H!lC�bդ��%�i?8�2�\�\9�<�0�Z=��} ��$�D�r]�&ΐI����&%Xiβ�g�O�ލ�&Cw�~���lu�1�E玣�qO�3�'30�'�L�ґ��@���*�#��mQ�'Q�\(�g�p��Q�	&`�@k�'���`ۧ-݂��b�K�/��(��!�'����P&����O��'@1�ش�rܚf��(2$��B�=o��4{��'B�C�0`h�C�=Ĝd�gE4Ul�'��)ηT	��8!*ݸ�Bf���s��'P�`H�L�^�*����1H�u���!�@�`ZiK`(�HO�`���L�l����1���I���S�'	�t*ҦO=P�����/k���ȓ2l}�T� !>���P.P�n�J����(Or)i��v���2��Ԁm =��`�M����?q��C��EV��?����?���ߝ�%�F�>X���Fw^\�A�"k7�O` �煊�s�1��'Q���b��1_�m��\�.���"�G�8F��ڦ��X(���/,���ē`�����1f>1#����=�=	��d��=���L<�)�+m� ԂD:4ZRh�1.
P�<�Uʎ"J� �#�!/Y�>	�ѧ\e�D�S���ĝxb�&�&���A7V��RGσ�=v"�Q%�N�_=�$�OP�$�O����?����9RWܩ�'M�C��r����� �'	� �>R8�d�3�@�s�h��Fc�+�xҠ�-��xZ�	$T
p��R �������?نD�KU��	�"�G���S�k�y�<��a�5KW��p���e
T�+pcZܓzU�f�|B\1c�6-�O�6��C4b�hߒ%�^|�ݯq/H��	՟��v-�ԟ���џ	�.�n����W7JA\@g��?��4�aфy�<�B$,@1�홈�L�}c6�b�$7��`ං�0(sTxÆ%K�O�|�
#
ރ`�`E !�(�-�>��I��@��'F<ZC�J�L �l1 �E��'�R�'��O�%��IN6j�v\�r��r�H��O����!N�$�ug	}-�)@��:��ȒӦݕ'�h�:ul}�*�d�Ot˧{F5�ܴV5I2�D�3M+��2���N�ZAi��',�Ò4:Z���uM��3fD�};P���iK6�2	�#��q��5����+3�'���R����	3ft`E�[�g�E���~8���Í (�����j��Ɉ�;��qI�����,v����2�M��i
b��ϔupl�V���7cv�򅈅
D�qO`�D ,O���f	1���'E��hZ$)F�'�:�<)!� �q0i�휷�6��$�	e
6m�O���O�VP�I&����O����O�֘
no�#�,R>7�ɋ0��MJ)���Ī8��ŉa�פ��	�a���O��Wx���%��#���R�
��|st�T�y��;���#�2�3�@�n@=2N?�mZ<;��D�g_� #E+5I��B����F���|�(ݙ�?�}&��s����ja`�ޟ8�f�y� !D��ۣhݺB� 9��f�d̙3�3}2�.��|jN<i��A=lx����g��0�AţF,�����/���',��'vz�����	�|2�D"�ݸ�n		 ����1&[��l��g��Da1ʚ<*p5��$��3��؂省���U+���[p�c�QQ���"A���B(c�*���B �qO�P�p�&9[���`��uj�Q���̖3��'���x���h|���H�klvI[
�'{�9;�^hf��Ejѫb	:}�{Bj�8�O�� �MԦY�I��GG�>'�qp�O�c6�ʗ��?��9$b���?�O����@"(Qdv�3Tn�w��㕢��	G��qt�M}j�M;�)H$^[џ ��A� 5*1�VIҽ����D����л �|���xr˗�e\�mZ�C&�+��:�	�	���0�$Ez^8��֞v���N�#pC!�B#ZB���*
a<�DL�(C���D�4-�P�yT��,6�DJ�mZ�jD+5��Z;��n��X��D�����X����"a���{#e
=Sv:m9R�>��D�O��J�!ߖ�V��N9W��
0c�a�D\?y��ƍ`���8 �&F�Ijg,�z�$��%��.`���\!(�֝�p��e�a柤XQ,��.��uIv�([yF���x�lJ-�?��y��d �3��a2CQ�6�ސ�����y掍,���/V�o�yS�/)�p<��剄cPaK�*�$<�ޅ0�
�*�a��i�R�'/ZP���#Ӟn�"�'2�CSK�d���A���>�U*�`X$��Ax�G��e���%B3lژO��*�ҙ9�!_4�%�+R 	N���� n*��`
�) �H�����Q�K?Yo��%��ޔm6����T71�fm�wC�s"�y�N>�7C�ß�>O������R�, ���j�`�"O�mx!�W@u ���$^��3�>��i>I&�� �� �5M��CQa�X򐜨�n�	�i%k������ß���9�u��'9�6��@A J<C2�=ࢆ�� {��	7��7'`�|2��
ʈ�y ��������j� ���l��+[�|������6o|�� I�={�|��IoӰU��*�7gqO�|��o�5%����%Eռh��r��k�b�'�9X�'B+�,�˷K�a��'��Z5͐�*� �flŀ����{B����OZ����Y�����ʦ��&JC�:cV�@vER�hM,�R&�;�?)���P����?a�O$���i =Z+l#��г`���j(_s6�P�b�+H�a�I`�џР��U����xQ"�=[,�Wa��	.��z��·,��0 ��htVPoZ�io����3�	�5����4���z���G	

���I�!�!�ċ���!ӱ�9D����Ǆ� ʡ�$��H��iB6,CA
1�� �/�m�Ɗ<�$c�il���d��S��CZ�T�G/U��l�I�T�P����gq �D�O��P��	{�{w�4c���r�O�A�TV?�Q%@TAS��ӁA�-�VLâ�2��K%@?��w�U-��8k�L%F:��]�O+@�Xu.�j`�%�.5��������A!��1�xA�?��y���DE��|�gk�5Ym�D�C�L$�y"�S�j
x��a�&J�H8���p<��	�C^� @��R�$���W ����i�B�'�"*�&{.�*0�'��'��;`-�Z�bB�Ǵ䑄�սuHR� 7� 3O� ِ�G�}a:�"�`,1���'Mz���˒O�2�0f*�
O��m:�F
5L������c�|�WЦ��Om�<-��ꠈͬ _ԊG�C�3L���#�dC�3H��L<i �\�;1��1e���\�@��C�<A�L 7Wm<�a�ݓ4��k�e�{���D���OL��',@�$'�$���#ayz��!H�@��e�%�O����O����[��?i�Oz��Qf�E�G�\�%�	?O�5�'�W������k5:��"x@џka-6n=vh���ؖ9��萖i�f�����D�&�b��)�^��ioZl�:P���=��7[�l�D� }Z�d���̣�F�����O0��	�d��ز�_ks���FiNC�	���0J%`}��� ��[➸�ٴ��3n̼��i'��iI:��C+��4���o�3�mz���O2��ϙ%�����O��S5�4�!��W�
; �CĢِ
���H@H�S����`f�/U������O�!#VF�д��(C�G�`<PD�P-El�+�	A*�(�
gB�6a���F' ��d���<�$F& �b�<}�
۾P�i�|"��9�/S��yCK�Cb䕢�� '���p�K�(O��=ͧR��s�ǂ�	D(mI1�Tbv�j �����)�x�0�i���'d�S���n��2�iP��މIb�󀓶��z��?T��"�鋃�8f�y'��u.��`f-��ijl�l8���l^X��&)=�'�b ��_�?�e��+�?	P�p�D����O[40�AQ�AY�(���R�D@)+N<i���䟌YN>�~R�^*G/�5�%@5l\�4��Jo�<��튠"4+5H^+�d0��#w8��s���N�N 3�&x�$k��� ���ܴ�?����?���͝pT�`��?I���?��2W24@�U�0��4�R@���#ǗF:�-��E��y;�P���J���OTTP$�����UnP�գ>X(p���	�]ɥc_�mS0��?r�E�}������n�<?�0m����<Se,�s6��lq��K>Iv�؟�>O����Ā+Cpa3ԥ[0&��p9�"O")�ćXGh������{MHXy��>�i>�'�D:��J�=R��"1��c­]�4�J��Vϊ��?!���?��<�N�O\��b>�S6�ơ;M,=��'��0��Ϋ>O�B�	0/m����� ���(�l_�8����3D<�p�b  +����"F�NŬ�@C`C�B
�$#�O4 �%֪9��i"hC�%M�ec�"O ���%T�p�u�����]Pe��$ ��a&�����M���M�� 
Y����� *2)8ՙ��C{#�'@�]	#�'�24�x��F�َ L�U9�J�k\h��kݟ�v��o��[�`�+�%�s��?�Âߧ)R.��r-3}�9B�@�9�F���mO�5�X�Ďj,�����=��A0}���(��$*���;�][$C�yb��zܠ9x�gP�3bP�!Hպ�Px��+�B��2��U��ЃP�U�J�E��|�iըW�7-�O��D�|��!J�M���>V(�X�����ht�d�o��'
�����Kj�`�eF�>a!N�m�|R��ju�ǮT!A�� 1�!�:E�5�xr��)�ɻQ�V7�)SǮո |����~��o؞jF8����S�(��2C�F��=W���d�O�������1�)U{C<!��@�G���!�$�Ol��d6w��y�%�D;��|�0.��x)�l��h�c�Q��� K��W��:ߪ�Mc��?A��`kR����?���?I���� l:���y�qQl�>8Xq���E��v0(�'�izqh�|J�lb��+vk�T�`��N/��Q6�ЮQ�^��aD�ob�G@TWG �c�j�3O�Q\�@�w��j4�(K��9;��-E}vI�aNh��,G}~���x� πDl����Y-HX`�s�D%�yriG�L��u+]�<Q|5k��ҟ���HO��7�M��yH��^�Nb$�Sf��6�а���վ��������	ϟ@_w��'��,@��р
_G��p6'�	V9�;e�<bd�'BӔS����d'#$L����% �h �*K�L�� �#L�V�	1�@7Ø �6&�VW��-�d��0�G{�5r�cBF&�"��΋m��4#R��7�\J���Ke[�r;|����f����>D�`�@K^]N�kvn"t��(��?�Ʌ�MO>!VI0"��'�ɕ�) d��/	#�P�)c��w���D�OJu˅��O����O(��)Y�L�� lZ�"��i�2	I^�t�����D�l�ay��ĖCTaBq/�F�A)���,A�0�89����d�c��Ɂ���3��M2`�VB�a�&��	ݟ|C�4�M����f~��p�!V�\^�0�eY�T�	a�S��B�BɈ3	�<	��4FD*Z��($�'�bQ��E{�O����]%EI��;u�^6 T%��,�j7�<�� �4&p���'VY>��Ս���5��aV
�ļ��m	!h��M#�?Q��!�H�1Q���oȚ ˤG�5��S!�|�Ђ����殉3���x3��M�ʁ�x���|~����-2��p�gؗ% ��@�F[���RU:���V��"y�nN��)U��/��S�8` ��ፘ�N�
�����N��,vV@:��L�*�[�M9@"<�㉵�(O.����[�j�4xr��v�xPƘ�Mod�N���O4��pi7:ڼ���O �D�O�#CS�����ܛY����vX	P>0b�Ԃ��4,O�p�-�)
R�:D$C�oӼ]z�/Y�ay��Z�@�`)d*��m�Ι�D��*;^b���D�Oq��'C��x��D1B�8`�aƯ20h���'�H;�A�|��Ds���(�A�O�r���)OM�b��P�.��%�`Ci!$O1U��q��N۟��	ҟT�	�u��'"�2���c&�H���I�� gv�X��S�R�Z,�`����s�K�SU�9F~�朦U��e��b99��x���VJj̳�7~?�!��C?m�.PH�Dʼi����dU�	��'�%A0�%�0�Ju
��
��d9B�D�?aԻi*h#=	�}"��������ڈ��d/�p>)K<���#�jd	G^�R�rpjCjܓ'ƛ�'���`Y9�4�?��4�^�;�dΎBxN�@3	�1:<Rq�'[B�F�6�b�'��釖{��ca�%w��#M���B��|6Dms��
A�����	(������*熍��Bġ҈Q1 撔E���0���МJT�2��(���9K��n��o��P�vˀ�1�(~�^�1�N����O���?ͣP��*�������A���R� ��SA�0���QG�,}�8�,�(�10�O|�eQ�	Cs�i��'��6��]lZ����OD1K�^�H5J�$wU����?9�O[�m�n�KA�=>���a��P?��NN�^&J����kW<]bt�|�)�S?�Kw)��(zf�N1L��c>Q�r� 76$��ӽ7?��Ue-�d��{��j�plǟ�$?��`&1yG�2�����CӺ(Z���=�����')�'����V(*"�1���k0r 8�^^��$d�O�uX��V�{��E�er��t���M����?!�@Hx	�'����?q��?����5֥ 30�Q�،[K�ɋR�A	z<lP��-?��#�����|&�H#��#0sB݈���'`�����T�G��+ ��?�x�3%��.:^c?]9���y�Wl�rQ0����0Q(����a$��Q��Oq��'{�큥�كDMpDX��B���$�	�':��@�3������.��H�� ��4��Of���HVp20z�׿]윍3Ff�M��X�C�l�I�h�Ɂ�u��'�R<����3㈟I��@��� �~T�g�� _!�D��x0��p�K��)A��p0I!�O�"�EP%��t�t΂�Rp��L"am��Tl՟<�'�D��/^�����NU���U�^R!�$�����"˷5A���(��=�qO��'��ɣ2��Pٴ�?q�4&�fT��^�	 ,�T�S���a��'~���B�B�'��I��?��xb�ފc⌠�F��oF��l� ��<y'�F�p��uQ#�߅i� �(�,W�T.D,��I�	����n�ɥo\�a����-H�"ÓC!��&@�P�w�N
��2�/�&
0���̟j�EQr/��$��,��Z� ��ij�{�Lـl�67M�O��D�|*1Eƛ�M@�R�*�����b�P1�#(-���'�vmJ��'�1O�<� f�z�n�-%�`�a\ +�l첗�x��ϣ�O��=k��R�I�}��ϋ�O��mag�xBA��?�y�����_���$� ������D�<���$M6�j�j�hs��r�$�@8��#���]u�0˗�	�^�^���L�>���ݴ�?���?Q�I�-ssa1��?���?�]�JH|��_��faQ�i��_p���y�����<����"n@%!������Qb�t�NLH��N6|c�
rKA��$|32�NZ��$l�)�3�dW����j0i�	���G��[!�$_y|x��ԫx�j�U� =�(���?�^�mn�`���dp�5AS��!K��ajV��?q���?1��`o���O��h>1hc(��j��lRu%O7p�����m�
�C�I0]�9���'��(�G�b�*�z#g#���W�ر�@�Z*C�A��"�]���DF[���䪂`�V5���S�pu�Am9D�81�Et(����W_�2��e6�I���'�`���c���$m�|�AG���c�u�H�=���ȗ�Wȟ��IH�M��̟�'/J��_��4M���׋G4�Hy)�9Ah$���
�u|X\���'����������� 1�!+&#V�L"w�8o(�� ׊B�.�ج32����Oh�7�'�'�pV�P.#�j`J� �/R����'#�< �LH�k� ���ӓBD<9�'���uK#bi�t���x.v��6�W�X��'p�1��w�x��O�˧u<��ݴ^�4�*Bd
��`�q/ �5E��%�'$b��-/�B�T>˓xv)��N�s��5���DCj�&���*�S�';�L����b0!����Gb<�&�|bV!�O*c�b?���_d��0Ô�r�@,!��1D��z�׳f� c��Y[��yu�+Od$Dy"n\61ON�s�(��CK �х`�2��ao˟4�	ϟd�%E���������Iҟ����	:�h!!ܚm�4��-ƽ?GH|�<���dX�L+�e��x��鲁�+j8�X�e(�I�yO^��N8'hY�E�$P$�ha��~B��<Q!���>O��P�d��R0�H$M�΍��"O\5�&��&���Y�g�,u��醑>QD�)��U��*1��Y?؜zCE@*4^9����/`������?i���?�!��r���O��Ӄh�����CM�nT4��,�q7\ԫ��3���3GP�Gy��X*��#d��C���E��E`b��1���zG�Ս�����
�O>�����H��j�f�=$��"r�F���B䉂"$�����)yk@XS��	=�����}��<], 6-�O6-���0�N߼$v%	 @��g���Iϟ< tΗП����|
7��@�<�8��\��ȹoU�/I� 
�Fb��Y��ϋ,&��������3-)����B6�v\�G�ˎ#W��C��4���U!��|�2̛a#6��[�B��I��7P�"!B������ى��ӕG6�B�	��^ �g�A�A������v5�B�3;/|�G�C�2؁��hТq��+7��J>O��o��IP���/����R. �ڔ�R��,1LM!UdT�d�8���Oh�k�G�ee�=I�ߵ��T>��O��˳'�M<����Hw M<	6�?���(ԪM?�#BJ��~�ִr�ɔ
���q� 2�D�(��!���3~�rr#�L�J�ZB+�3!�$Q�f%|1iF�] �	*����
	ǓY2Q��ᤦD�^��H���*.�};��	Ck�f�'(R�'��f�672�'<��k�C�>?����.�lJ0����f[1O�Eȅ�'�
�`1�*�T@�4+�x�0l0�}���+��<�U�.m4U�B# :l�큂
�0X���O���������?t9���1#.�9R�FxR���e����A��P��
)bU�h�O�8Fz���K7�ش�T�I5*�ԺqE .���yc�k�'m�'���p�`<"���|�����+�>m��듴hO�>M�QnR�b��P��� +<hp�Gh<9�H�m����WJ�AC���Uv�<14�٬9�v��$��_��`81C�p�<)�ᚻc	`=!a��\� �GJ�<Asǝ���Uᢚ��\��PbQD�<1�Ėp*�iP�M��s>�S�
E@�<� ���n		\� �w�ȶŷɩ"O�)9�@wn�H��^�8ޞ�2"O�8��	��D�,e�dc�,͞�P"O.�L�$Pp�3�T#L���"Ol�ҢFW�p�����,d�^ly�"Oȍ��;HV�:C��`l*HA�"ON���H0Ɛ�J!Dĩ<r2�`"O�J��m9�X`L^	(}88G"OR\Y@.���YeW(Vކ�id�#D��2��I�N�y���Ū��S%?D�����n ���Y'8Z(� �:D����@���$A�lV�&S�1&;D��ʁ��$4��*98��x0V�,D����eJ�M���!��lךP��*D�At(�?�PUGI2��,r3�*D��8��
 8��T���R�m:�$D��8'�\,b������V^B�Ճ!D����넼�Xp��Z;_,=�f<D��З,�_������?j�ق��1D�����>B�l�������0D���@K Q+��J 
�(&�-(2�0D�`ڣ*���11Q�U���*�/D�0ڣ�A3k�B@�\�?� 0Ŧ;D�D$�k�"���Ί|�>0��;D����2V�p!gC��&�wC6D����A�4(��bkWw()�F�6D�4(4%΅F~")(IN�u-.i2��*D�,���T��@h��
4Lve�""D�XٱN�7i <B��U�j�M3��!D�<��l��4�́���O��U�B�#D�`��f��*�HuY��aR�9`��%D�� ���$d>xrE�ۓQ^���$!D����+��TZ��[�7�tx��@?D�,kQ$HI���r!̹4ǎ��6D�,�2���=(�[���". #�''(�1d�����B���/�܉��'�����&�zr����"9���'��`�hK�7!����\�}9@��N7�!���$\����)hZ\B�B�&Gay�
P��$���4��f(h`������A� *D��qb�8j�����mY��\�`+�d75����{��D�E�	�d2� �(`ђua#W��y2%Î@��Yf��tB`"�1WqO2=h�gY�g��N� ��.��3�.p��e��.�B≪K�4�{��<�T#І�,&�Y�r-B=t��R��$%ҽ)$�� v���@!���<i�醓O)3�@��@h�)G� �9�(p�"Or`w�?3�l嫝�$Yf\�Ғ|�˝%[�Oq�$l���ܥ2�����,U86�zv"OB��i�'r��2��X�;s:9"O�b��C���P�]��8��"OZ��SC;�R$��d�/�V Zq"O�yu�+6΢c�#�:m' E��"O
Hqo�d���&DA�W�`�"O��;����W�H �bf��_�FB�	�9NN�4÷rh6dQ��V%S�C�/3�T�����0�j��!��C�I�068�Y���-L9H�.��2B�ɧu~ 	�ѧ�+Q��j�IB�'�B�I��8��N��	��G�4zB�	"'1x<S�m��=���G�&!*�B�?x��� ��7r�0V�	�()�C䉒AF�	á-C%@:���iƭ�"C�	<�η�n�'*�f��g��%�C�)� ����IT�]Ie聃[,� ��"On�[�g�0Ă����#p�h� "ON���������+G��9 "O��F�ح�dĊկw hy�f"OZ�ک���AW��eٲ�k�"O�����P,��L��	�
����"O�=�"ң:V$�Id��.f���[�"O�H��n�!�X�Aq�]�A�
q�"O��D�����U�DE"_��{"O�QI�~��b�΅*�~��"O�A��1����E��?��8��"O"�bVj^�K]z��b���<�ɹ�*O�aZ�"�k���ňs��d��'C���&A���,����i% �s�'͒�cA�֗|=n4Su�@�iĨɇ�!JD��@��g��,sV`��;�����.7T��J�u��@��BP�`�ȓ��L�a#�<]���`d�\r{�ЇȓMO�b���7�$���
�f�TЇ�>Bu �+�cC���0�[��\�ȓb���0�%=��!D�d��ȓk�6���.ӅY�p�a��W:�،��J��!�i�/׆���NV?���a��% ��^��Q���C;H���6���xb
V�i��S� 6<#H8�ȓR���B-H�&_$\{èǻu������;��C-�𬀀ꉶ^�"�Ɠ{�eR�i�9>����w��q��ɀ���x��*F�	@��}v�]�F�A��0<��2.��3�"}b�(=�ʼ+e�ީa����!��y�
V/f�����nK�]�Iy�����C�,Jpd���r|���X�v>$�9�F�[�bUa�Ă!3*!���U@d=CGo	�;�����H��n$@%d��؁���E�~a�H|�>	�P��hh��N�,M�e��MEj��xC��غfjT�*�ɋaw0�p�A_�b$��f���QV��8FG�MX�P�gg�(���-J[���%*�1Q�T�_ ��G���j�p+�˔�0c�	L�+�]q��
T3K��HE H
�'2l�UɌr�(�8зp�ucĻ�yB���p�&�p@Ǆ2Z?H���A�f�O�����:/\�m�B0M�u��'5FhCgEïq�� ���^G�����cE7wR2�7�	3|;��!��(��I<*�#vgӝ_d���iSJ��h��	K��p���Ӻ*�D��A�P,˶坜���˂��T�2x0TO�r�,��B�|��iC�*>��0�Ek:�i�6��% ��#~�$3�N&>�rݒ�O\T� IB)MKTy��(��*�'�1���xl�A�K-<E�����%�G�QB>����i�=��i��+J�̈��	�?��Щ3$A���C�I:_��'�˒5$p݊��R�2҈�U(@9sѸ y�ׯM�4�[�|��$˿RҴ@��i����Q�Ô=��}B��?��ث��0F �pu�ȓ	��]	�f�3�D4�`�S�,���'�$4�י�� c�=s�Xi���D�<Hd�Ն�:=�N�H=TX���&X4�@[�'@�:�AR��G!f��C�	�S&Q G$��f0�,[V��8��D��s@�E)��O�`_bJ�CR$�}�����$��$�C�4�(�#���y�I	��"��u�,���C#��~��� M�[����\;=@��ϟ��� Ǟr���	�I�w��[U%+�O襲���;�h��M�Ct�~k"�9�� Ej��� ���p>��A�-hV8�r�LӅ[��=zъ�Q�'Т6%+T�8E�������
�(t��X}�"<94hH�DB�ɸw���װK�:,a�i����h��Q���I
L7N�P7G<�'�2Hf��8&��F�nr���ETp4�s�ΖHu��i�$�=5��=IdESyb�5�҈�ǔ��{bX�}�r��A�u���Q��Px�B�g�$��I�l��@8�U�&�kʢ=�a"d�9����QG]�Q�����E��0=��%�)� (XB�ˁ9��ЖIǢb���P�"OM���MX�p����2
m�Ay4"On��e쇸��${Qf�~I�qab"O�1�f"iVm�jA�|�HJc"Ot-j�m��$���S�6<䪼r"O��B���:j?�yӶn@?^۲���"O���7^�R9*5��h˞I�@! "O6�����6��A�o �9e"OV�B�!�Um�� ��Fna�t"Or��Љ��>XLd��	��&"O$� t�6u����%�E�W�4���"O� K/�%�۷�I�`�8 �f"Olf
�)V�,@C��0a���"O"� ��\1�Tx�	��l�'"O�,j�!X�c?���C�N�V�T�Y3"OHl���,�L%zpaF�h� ��"Ol fJ�+>RX�9E�G�^>����'�zH+#�O,9"ޏb ,`�d*+S����"Oؑ9��Ȫ\��,S��֖@�qQ�	��֍���;Y�n҂�\�1�ЀG^�'C�	?H�o	YV�y*�I���ڱ�c�����"~�I�mp�BAU�]Ǧ�A웲3��B�	b�����X0DE(٢�l������%G͜�'RT@�U�I)H��IU�MT`��T��M~��B+��"���'d�RJt��l3D���r�Q�RQ��(3*�x����0�0ʓ
���"�1�>���@�67�(� D�|���ȓs���͍ EY4e;C�уrATQmڃ>2���?E�ܴV��p�'�-%x\K��S�<	VK+h����v���}*4�w�S�<�᠚
t�0�To)B*�d`��q�<I�P����d�)9t�|X�#�P�<i�F�����3rи�k��T�<A2kЛi�8��I%&Pm�H�U�<�RH�aKT�(�%�GK�A��M�<�uG��a2�r	ˢ-�~�KӨ�G�<)��J�i|qiug������T~�<�צF�ir\�V'�#<���`I]�<��+D�_�(e�F�2[L�d��U�<�ӂV����2HB)����jZm�<�$��I��	^fd5T�Kh�<���Ān�S�� H�z|x�A�k�<�� $}<Ȉ�/�!2>�`���e�<9tM�)0Ty�X:i�8���m�Z�<Q3j�8:c
%1q�f�~i �&U�<�aK�_�0��e�S"мE�O�<Q��@��̘5( �L�l$H3 �H�<d�N�%H)Q���d���+ i�_�<9Ca׬i�n$�sd�\�б����X�<�'i��D�K�Ul��ȡ0�T�<a�)(mo4)U�K�f��`�B+D�x��F�w���Ȇ%Zpi33�)D�@'LF 7�x Hb������t'%D����fνh_�90���F��\�C!#D�dYq�1Jm�X��4*� 4Y��#D���/֙4����c��hs�uS�<D���&�%H�ܓT�Łb��ܩî<D���$�C
$"\xf���2VIU�1D�`P�ۏi4�ر��W�BTQ4K-D�8`f�5*jݻ��bm��h�+D�����V�=+$�N'q����5D����d��g�D;���: |tq4�,D�{�]�.�yS��s&8A�Mrh<�SLǆ"�qQaIK8H��ǠX�<� ��j�̝�tb�����Z�L�N8�r"ON�r�+ߕ1K���ah�4٘	ط"O�`z%��J�T���N��(�RU"O�cЁC�"3�0��Ql���"O� `-@#:$YѠ�.�YQ"OTM�H�;c�4��ƕ���Y�"O�՚�m�&Hf� f�U���cE"OvI�f��y��b�i�I�"O�钯Uq�����^֤h��"O�-�W,�a�v�����9E���"�*O��c?f�Th���Tk�h�	�'y:�X#�ʥu�V����J�H �	�'�>������D�����A�䙑�'�(xڳ%5�>��@��89����'��"RHGRJ�S��B�,ðk�'��#�(t]"t@P�3r�ы�'�����f�0����PɊX�	�'��g���mn���ܮ��l{�''ؠ9�#V��`yq��$Q;�'�J�0�K�zΤ�P�a��2v|��'��Hs�@�+Brv�xP˟um�1R�'���č��A��x�W�]�k�4�B�'�2ᙡL�p|pׇ]�ƁS�'~R5A�Ù�m�����@�0Y�*x)
�'�t=�E�̖v���
�ׂ^��X�'P���Id�p�`Pf��X)x���'zuB'�]z�MՂcL��'�U"U$B�i�>m��c &gwո�'R�$"��Y��9�wOJ�`��<
�'�R (.kIP�LB�[a ` �$���	!$� �G0HA�	P�5R��h2UeZ��T ���R���D�D�zLT����O�s3ȋ�"]`��l݋gN������	|��#�n�73ź�8�ɚ��']�"��R-�\�^`���7 �:��'\rxx��d_���tJ��H9�UE�T�SU^�miv.ηj��uk��9v%<�S�Mʶ&g�}��"N�&�P�c�{����9Dq4Y7��C �0��(6E�\�@�d̙=�a2� ��fkFÉ}RbG��<�]��r��q�>!�&"<�#��?�rDf��%�콓���:z�8�ˀ�LF��(Zf��)kJ��C�3��?�Ʉ�\>�y��+pV�x�d=t7:�h��K�MSgު���ȟ�@�B6�؁5&@�� �����7`��$�0��0\�<�c\�|��'c���VO�).
Aӓ�K�]��p�'BN�rU�ԟ��Kí��89�O�*2�Ps���j<Q5 7Xa��&K�P#���3� q�n/��?��pH!���d� 8�b�<�&\�'H�@r��k�<l��	�~�S��`̪%S��:�+��/
"�C�g�
�ƭX6͙�c=��'�(��T?��Ώ4K�:\��J<	6�)PF9Zc�i��8�6m
W��24�����KU,�@A��4��b�gR���q��E�S��E%`��ۺ��.[���44��1'��G�rfD��d�M���$Fa(���O����O�MV�xq�Ԧ@��x�V�l���ԫ#�&%*��>��c$6hϓ�ti��C��0w�-�'.T�\v^dr�K�Ԯ w�ς8bB��a�UG���?%>m�s㍽-Z̵"��M���2�D��d����'m�M�n���M���O�T�+I
�x��¨ђ3G�0Qd%_U�'
�#}R��?�b!JF��2G����f��&���u+�$�\<"wLʛ8���Gy��f8��q3�"��S�P*hƱ��R���p�i�H���O�Q>	@��y�X�N��\��n'�ɲk��� 18s�l��v�'D|ط�O2C���fH	�J	�֧<1 �[k���4ŀ2l�ā�B{� �C+�-?^�B�U�@B�re��~4"ٰ���d.X	�(4�S�S���{%����l�h�Ύ�vm�b��j�ƞ�6����Ð�":(y�}����E:�T�J''�|���Ά��yA
�'D���-��L2x9Cc� ���tJ�]\"� �0��?y;Gk��y�lY?�ɹV�U�EԺ$�$H��y�O��_?����.�{���Q����'*\��f��G?~�q�#MP��OX�#������(})Z (u�'�J�Г��gX�+!k٦��jˮ&ɚ���NWUb��eʱ?,��h���>��{xj�?!�53�)�.bJ"0�Fi�5��IB}Ba� �FfJS�Obd���*bU@��g���F� ]a��'�N�O \��G�? Ukl��T�*<x�L��IФ(���Q�fA6�K��ңWOQ�x� E����J���j_����E�/��mZ�<yL��?E��m�m����:4�bU�V�-��i�Pk9�J5�l��У^�4�`Q�F�m8�h�'�ܰvβ�b!�p�ӫ=�tX��O��!����t�܇������[V m�Ee�H��)"�*�7��Ph�
�&Զ`��ƌ(��r�V- ���� �c�xi�ʱc*Y��W �I�#G4U���9F.@�g�(k����@D�w$)���KQ)>l�Td�J�����rܻv������M��Bu"�i4'ם+g��;�M�9_Q��*P/����M�9������h|\h��mʎǛ6��Q��O1��]�2��1v��.ĪPc��yr��(�X4�Ƨ��Q�x�� Ԋ���{v��/h~X5�¯�<�5�&xe:d�?1�@Hr�E~}�#�C/���~-�0�i�$�(	."��scХI�F�GA� U�b�-Ը�0��h��>��P��� 6\B�YT�kqO��O>i�6�D���D&� ���i����4���^ȅ�,R�6~�|Дe���"<�䠌An�	k�O�m��	�@�	1��x����|�?�S9obl�d�-I-\�r���2-BY�!N�j����P�TרO�)�&l�%�y���,x	�\��Ò.7��@��Yϰ>	�(�Zx�G
U��*f�'� ����$Q�Q�H�F-
�(n�-ge����<���
^����[nN@����VV���cg $X�qq*�u4�E��L�rѨ2�&J����v��	��6-LZզ!�@!FRY�q8ũ7d�������0R]8Li��]�0���c��<�4��&6i����c�	.o�l�5�Dw�'��TC['S����/�f\A2QƑ� ��D�'L�z�́�l��刷%�l�zd��$VI)���K�8{���䁵cX��H�m���H6X0���2ns,��d�<�g��"dg҉� �۬G�ҭC"�f���ɛ4",��2��1F2�u销��Y���ɤO��D�`N[�.���@��hcc��'�E�dFK�n��B��(�L��4}�$:��2�P�� J�x��I�#�Q#G�i�A�3z2�'(�b����J<���KY�z�0� �>�%(U�Jz,�W�iӠ���B2�HOb���΍�>	|9�D�G�w�� �R�$��^�a{bCڀ���dk�(����JK��?ń�6V��m�2ْڴ�t�cCdηBj�9�n(t{j���I�cn�@�_�<`�'��h 	$f̛F�F+2�5ړ����4�'K�������u�Q�bjZ�ڀ�?�EcI;��#��=R����Iה*�B5�C���q$�,qO?ٳ�9%�I�uFAx�n]�W�E�fM^i��h��$�!���ԯ@��T�aקB��I��h�b�5��;��_h?r��ʘw�>�ɟS��4���'��� D�ߦ9�qL�H�}Rc�Y�T�L�٣���9$V�0ʓ�9{������'�J9�uD�5_�X���A�(�TLر��i8�=�w�G�ju�2U�v�z1J�[�t`�N )Cx��P��ɧ��(ae�$p���3��Q9��oyB����r�a׿3�JY#
�M$�0ol�pZuEW�V��Tz��E֟ ���t�h��^�g	Xe � �8qYsIO�6
jUy�'n�$@�n�V����g�IT��C��>���V���Rg2m'�h��FK�'�f8 ��A�P�r�D�v{�B�e�#  |0�
	���k�#�|�T?����A�r���eM��-?U5��J�A�,��Z�li���U�G��5��kv��֏�|�Ľ����\r��L>����|G��>�<��K�/��	����e\&\�|�u�O0�(O���'��I}���mLZ|�q�O|M�hѰ>���ҧAG�9%��ФC^1`͖�����,&�hҕh^�/�4�SH�%R {AF�8!Y|$��D�$V�����#�W�4���W�:�DI`���:(�R��A��%��H<?�S*%[~�K�� D��dC� 6�D�F�@�(����쀈H�lۯ>	z�Gx��1B�Jtz# �D#6	�6E�.a�\#�L�B8A6f��K$��'>q�t��N����f�?c<i�!D�`�2����=0�&p�7΃v�'�Bu
b'���!��ҍ���f���W�\�0Y�-�t$͘�L<a�V�X5NՔϸ'�2��	'R���*8!ɒ����F >,�<����I�R���"aI�����^|����v.#Y���G@��3XL&灠j�H0���� \�$�[5�dNb5M��G�� �D�O��U����
��E�D
9:N�*4(H�M�p�CK4_�����CT��	�jp4D�H�?��ql漫���@'<G�4>0�'N)z��%b�h}b6�ݼ7�T��d:)��I����D���2�4'*
$ e��0<[�pAƎ(�r��Ӝd�
��X ���[� �^իBj^�VH.ܠ����I�@k^ԩF2�VPK��]5*l�C�k�c$RM��e�$O�T�޴@���Bq�L�	�2���UT�n�|M��S�6�x+�n�LeQ�@�Pn�$<�L��C�v��y)�f�,��IáU�tҀR� ��?z�(%�;?>ЅK%%8�����{�
�?黧l�<ln��B&��:M��R7��*��} �G�a���L53�����AzE"dA��M�b΁��0� L�?�	`�>�Fo�O<�I"�~y���'x��L�?J|�1��Ƈ#W�옍�䐇H�̹9r!3>(�@��D�FNR�lӮda�� (Ò�kO��O��I5p^x�k�b۵3S�p�s�E�]4�� �w��j˕s��qF|b�ʫ;hU���� `���D@dd����K�p�e�a�k���g
�q?!�{�;q/8��Ӌx�����^v���?��&��Qb^q2t�Wq�gyb,
�o�Z%ڇ���)�TNP&r�"��t�'M�(�PF@2"��p�͙:�R���38X�F�6�ܝ��'�LA���5��e؞��A��r0����4%ZB�O;�� ��h1���[d`��'�D�3����f 5vn�*��Z6O���)���� �aM{M*#��o�@Eٖ��*��������rb��<��/t@DۚwI��9�BF!F����iH�/X��ٴqgX�=a!� ʓ�x4{���.Z|M�V�S8P��?����j򄇕kܴ��¥�<�C�H88��R���(���Z���2n����'�E���4���X���L���&i�
��L�	Ue^M
�߄Vrfh�B��nK$�RQ�ńpN�Lj)O���Jd�����d�"a*X��BڸzԼ�|�JʘU�Խ�ɏ!�f@)��e�P1P�2Р��;E(@��ڼ[�49  �<i��S�?�:��<��(��h�/�:t(SLЗ�<��7���Zf�0��3��?u*WD���yG�,�ԩ�rH��*}�Q�$�M�a	�����}��)��>�;z��E��@�AL|��*O6+>�9�?�b�WGt�̉"��X��E~}dO��T�U+UO�*ݚ���=Xv�qP8OR4�"��?ݘ�Ɇ�v�sT`Y���e#2�b$	Տ0ۜ��EP�R.�d!6�b ůp[���M@r�S��������A�W`ݏIj,��O��2�К_�YHw�ӜX�ba���	�@*�`���$,��#bؙ6S�����!N&��-O�M�3��~Z�Ղ3�-��$H�S�-�#)��X,�5�''DX�OB
�y���	G�<ɕ��6q\�� V(�M;�@�����h���ݸD�ܠ���!�vM�� ��DJ��1���E'Z����=}"&
�:q��)3Х&J24�A���$_�Q .��S�B%��q��գ�WeljY�aH��4w�<�4�z�zS®��\XKw��3c���P��T.,��%�F�_�1@�>IR�J�
�8!`��!*W�ȁ��X�7ǚe��*��W����¥<pCv�qw�ɮ�H�v��I�J�}[��R�08�f���m8�0HΗ5|,ԳU�(�Q�����-�9ͻsODP�>��!���![�T�8�LQA�Q���^ܓ�u''�i�$|c����1�8h��A1��'�8� �H^RS H��F	3U�fp&>٢#�'� 1쉔X2��vc�<هLԐg�b�r��˭96�����6�'��-�UQ��J�
E�
�@�ӕ�ʲU�jԤT��$���S��y",�'K!�4@c�z]�(V�<B�}�
Q!��Ǖ=b�ɏ��y�ʟŀp��W�
-�p���y��Mh�x�A0U��Q�W���y���gb�8�o�,M���g���y�B�!,���L�@PT���e���y��I?~��)�<.��rw�Ł�y��k��lr��2,���f��yRg�'S�䢡�vMv`���y�ռ�x�dN�z��X�U����y�� 51���/(,y
��\8�yrh_�E���QnѰM	����ybï;6�p�v�Ac�������y"��$FiJ���]B
U����y���In|���&�8-J@}�E��!�y¨L��V��)�#�dybU����y�e<=����F�ךF�X��Gʵ�yR�%�^L�1A��p8�����
�yf	�"�n� N��b3��t�A��y���~�����*�����Ū�y�	^�T��X��("�\s����yB��?rBvU4��8��HO��yI�:A:bبV�L������k
��y"��K�R��%,�p��f@H��yr�9=(��C��V7l�@�yRa-T��ԢUn�U�-�A�A��yb���^ea�	�HMX	!
�&�yB�	*��"��2xp���B�-�y��P��)��M�"�p�i����yRB�m�>���'�!z4��y2kL�E8�K�a	qE�pDS�yroƵ��$85Q�3�&(���yB+B/_��|cs��%'�b�J��X��y
� ĝ����7Q��G�$D�YA�"O��;��K�wڥ���4KZ6�/D��P$��`�>}"')�, �B9*s&1D�4�7�T�.S�4��jV�#�8Y`�L/D��q�:�ȁ�TH&Y_̥y��-D�H���Pؔ���&��[��yy�,D����Ǝ�G,���7l��	��&+D��1��{\\ Ja��kZ�q�	+D� �Ci�bb�H�4B��T4�X��*D��a �P�|�й��(.P�
��C$D���C$�5/�R�n͑&��9�F D��3���=t�(�C6 -X���N D����ǈ}
�hp�]�[�$�$?D�T	�O[]Ya���پ8���[4�;D��W�%}=�E�@Ėm�b��8D�8BǇ�a;�����(-	�i0�;D��jBg�|\D�d6`��9D��8�B־d�P�R�	�f�4�0d4D��!�,��]pC��-���$D�0�CO�\�2���M����0�
"D�8D�;?!��2�O�
<�e	+3D�h1�`[	T�!9A�
�쀚`�;D�h��g��o�ڽ���ƟJ�lR��7D�D��GЯx�ř�)[[8�G�0D���GF�}H�`g������0D���Ĵ:�d���� �+;D�9DG-D�P3bV<Y@XA&�ӷ].�ʑ�%D�b��˼!;��V�� 3�1i$D�t2$JN�|��m`a�J�~��09�#D�("qD�lI���AEǀ$V��G�!D�P�w�N�I�&t��9w4D�X0�ѐݚ!�rE�}��X���,D��a�$k1��CB\tar,��*D��bF �10�!�VP��+D��PЪҍ�P0㤕#@�<Ԫ��&D�,�,�T��B"��
&�d�5�?D�Ы�)I1Hj�M9���S��P˖C)D�(I�"[Z��駯 =/�|��&�(D��pՁ^2(�����\�~��cL'D����aȪ1�����[>G8��#&D���B��'I=�d��K�5U[t�E�#D��!�ňe8�����)t�:I�sD!D��Sg�ɲ5��(�+	8=j$Y��>D���"2tJ`I��� ft��y '1D��֥T6 T�s�A?S�a9��1D���e�7�DU
b)�� ���.D��m�Y���1�@ɣ+m>,I� \�<�@c:|��! ��PG xs��R�<)�c>�@1R���p� 봀�M�<iE_�q3�	���$=���F�<��CX0N�>ڦIB��1j @�<�'�:T:�I&�\%�r1�b|�<�b�1L(��`Q�`���z�<�e��jx����,P�J�����y�<� K7,^�L���]�Gg�	Y�B�y�<��HC4M�U9 N^G���#�t�<�e�������ˁ��<�
��n�<Y�lI��H;W�M�({��ʔ��^�<!�F�{����HJ`&��နO�<)� 9`n*)H�"�#4V��y��F�<��a�	<}f�
��Ȟ<�"Q��Cl�<	7���wǦcB��.�>�� $�k�<	Eh�?~i:=FS�zF�a[��j�<aS���b]DK�����d �a�<� ���a&�;\����犜O�U��"O�H)�
��3Gܒ�0�*�"Oꭩ��4qH�U�!�A2&��0�"O�����ԯ&�b���l��<� "O��#r���j��2�ˈO��,�"O�i`��L�7��=P3a�j��ұ"Ot0@ϿX[֌�q��.�JP�W"Oh(���xچ���o�>�����"O��n�*P�r�썛]�H1�"O���d	=�r zÊ9"��]!d"O�P��@�;���$) �O,�-S�"O��wnّR��`�B�L�s�m��"OLxSu��?�b}h�̟�N���"O���
�+͎i����Z�`y�b"O��K'Á<+���������R�"OfQ�6�I9K�D�ӣ҂[�RL�"O|�c��-nf$�j��^�~4���"O�"�L	*�<*�a��%���y2/j��lr��8	1���H���y�	�/F�X`/��yV� H楐�y���*��[��P.$�T�fU(�y�	[�d?,mb��R���7eY��y���>@a���
�TX�
��Z,�y���\?(�֦�,L߆���M	�y��=�Ι�$'A�l��STjH�y�S?K7� C1�� M��S�ß��y�mZk���O�Kj
M�R͟��y�O�^xhTsG@C�=�±S�jJ��yr�
�*�:��a	60�r�F��1�y2�V�6k:�১�0 ���'D�yb��)k�~,q�A�>/�(Ȁ�a��y��D���)�t������y�ιcȴ�v�E� �>�ת'�y�c�0���M��D�^Y�%Q��y�Ս�D!��#0����]��yd�<p
�Mq�j����ԳfJS��yr��2I�(���.�����0�ѓ�y ԓn\lQ!�Bv�(5�D\��y��� 8Rg�Z�k1���D�*�yb�ɴK3a �*K�o��	� ��y�ĳ�B��lСa�ƌ���:�y�͌*3�Y:f�B�m��L˓ ��yK^�x�$�� 	dh�K�눑�y2��,(��
E�׻Z�xb1�W�y��x�N��d(N�W�� A�ǀ�yªݗ=8�x�3�ɈO(Y�K^-�y�9E�$�!�rA��'�qR��2$��%(�
�r� �'��q����N� �k�/�=�h��'��u��u�-B0�H�	��h[�' �S�>:�� ��C�|��!��'�.4��D����+żP���'���Z0-G:G#�Ff�
fL4%��{��)��_�"4�������9�.0C!��E�L��d�҉T�
�\�Bk�e,Q�L���#��)���:�bG��eH�C��$!=٦,A1	��y0p�-u$C䉇tvz�1�>W����$N$ ��.2���Mj�jM�$'�q�!�d�Rؠu í����0�$��?;�!�$-E.��EC�=/��x�G9�!�$ׄ���SaF'
=Q���'Q!�$�
<>tq��N�o2@���qA!��
A�0!c�[�:�Y��E�e�!�� LJ�H��_�di�$f��BW����"O�Z����i�v�Q�II���R"O����F�HAX��'�GB@�6"OleQ���G�H}2���:D���"OX]3i�F���3Y<;1Z*�"Ob���C�)��2P�H!'�|�A�"O��D@J
/�B�bPHT e�R�"O�ѧG@Qh4�c%'ǐ4� �h�"O��A$���lᆈ�� ���7"Of���Y�t�	a��ϒ��@�"Oġ���6+teYaY7sz�Y�"O.����<md�P��E��|0e"O
E���,\�	�p��\N����"O� 5��'D���c"B&e�2 s�"O�42��73� ��"ÌBcb1aC"ON [�+X3# <���`/`9X�Y�"O&��e�ĵ5��$�u/τT(�"Ojd��F��_Dz5�!h;�IS"OF��ɘ?V��X���d�%I�"O*��h#�D4u�,�%H""O^�q���/i�̀��FA� ��T��"Op�U偭QI�X���H�x��:�"Ol�cd��EKҗ����d"OޥX�'�L�@��֊<WP�"O��k��Οi�YT
Ѿ/j�C�"O�Q"�J�JxR����_ CyT�"O�|#� ��[Bm�eΑ|nv�!"O���%ߴK�r��M;
]���"O� ��7<�JL3��^X��"On��@�6"������1;��q�"O\��4�"6Ř��e�27}��"Oy�P�דPLԈӳ�� *RC�"O�Ak�B� 5���̜		0j"O.(��J�&1߶2�D++�xL"O�i�U�ʺ��\���:L�čHC"OnP��+H���MV�z��a"O�MZ�ۅP�T@��K7i��m*�"O���T���M����C��^� 4"O��%��9k�||%�
�,�|0{�"Or1PEH�8r�i1�P0
��ܑ�"O8<	��C��!%+�:���"OVհ0�.p��z���x<d�0"O�0�`^�kR��� �p�DH"O�8a0ϟ5�8�#o[�E��AѴ"O��[��U�}�6�����	�"O���I@�\��ԸĎào�(Q�3"O��ӳ�#O�&�#`���\��%XF"OR	 �怣:���I��,l�<���"O:��n�yѴm�GH< x����"O(�`�o�f���Q´Hd"O�I�w;*0)���.��L�"OH��#���PX��]�[�E�e"O��s�+��%)ȚL�����b��yB툸t>�d��Fׅ=����6-ϵ�yB&�:J��`�/<tX�;G���yb�|�`�	��X�8b0)RV	߻�y'�5% `��2��7ez5��g�L�<ɲ��52V��`�/N;���j�z�<��;��=h3&N,j�d�� \w�<9VҼ^�@��R�����P�*�J�<a���So�ȩ�^e��=p�kSI�<�D�;&C条@C�2P�1���HD�<�v�8--`
CW��$���AX|�<��B� .���n�m��� K|�<� n�h��O!!(,��YS3��yq"O
@3��C�`\�}��(3REX1`e"O���b$C56�¬@q�ϱq��)*�"OJ��"2&�T}@%_�!q"O\��sO^<C�J�!ĸ\�*tE"O`��rDW�%�I�$/\�i��§"O(PIw*Z>:H�O,z:l��"O� !�o�q}(٘��H�TZ�d�"O���',Im�,يE�C�,9� '"O �*u� V�T	��(�8|1�zD"O`��k�>V�\���,f�����"O\��&K@��0���P�*eq�"O�mZ�Cمz�2�'@ d9�!��"O$�0tl�)��p��#�&�"O�q1QHM�g�B�[3Ǎ�r�θH�"O61�E�ժ>NĔ"�� z���"2"OvMQ���$b>`��,����i��"O�-񀆆W�Rc�D��"�5"O��7*F�6rL�����9�H��"O���닾)�Ĝp�fK>x�0��"OR1 c"�!3����²�0���"O����Iўm��e�
�����"O�-�JGX��@�%]3�RѲ"O�%ʄlW3m���� �()�a"O=u�M�-�,%�r�5�����'s�iY�A�$����h��9�'/9z�N\N�G@<dTQ�'�n��Ó�7�0�B]�n�<!�'S���$�*�(��-/�3�'��C���9~(ty�b�� T���'=�	�U.��&�BP����Ītq�'�<���k�	�Ȭ:B�A�qH�}9�'ѐhZ��V�?�����͔YrF a
�'ѾH{��ŋr{8=c6��<T��|	�'��E8·�X(Xt�E����TK�'�z�AO���I� � ��i�'ʰd ��,a��Xt��'e�Y��'c�p"�D� ���ؠ����h	�'+a���*OҘ�3����E��'~�Efm�����gFݣ �����'�v�J7H�r���ޘz� �(�'���%n�c�إ���~g0�h�'�F���J�c�����u?�l��'��`�Hr��)��fu�&��	�'�Nl����_�Zٹ�(�_��${���$Sh#���mݓr���Z��./�!��2�)E�xb����ː_axb�I:)<�Pgr�
%H�-X�q�͇ȓ-�8s��2�h��%Д��Y�ȓP�d�� ^2qc]Z����x� �ȓ�F�cc-y�p�S�`�&S��ņ�a�AL�����%T��`�Z'(h��M���+>!��i��ɇ>WLt�TFT�<Y�	SÄ]����]��	�iQ�<�(�8��}��cҼY/ @���WU�<�e.\	U�	����B���+���N�'i?�p��Z�i��%́k�L�O�=E��G��V�<��i�w��S7틭&�!�d�?,xB�)X�>i��@��D�!����8%��Dg=����=!�Ħ2��؁d��3;J}S��Q|!�d�OPU�c|wDp�S��`%�G"O���7g�
b\��� �X��$"O Y��&ݫ:� ��gB��ivU�"O� ���e��
%덗8c�c����G{Zw�qO(�c�CN�w�l��QyL,�t"O�-rc��pk&A+y��&"Op�i_�8S1�2��I+7"O=�&#�Z�^�w�S=
�9#	�'�(0"�@X8ф8�'ʉ�i�Hh�'�Fy�7FP� |Xr\��)C�Q�<��LɄDJȢU�"R�JI�s�Wt��'��ˢnʚoҢ�K$��D>�T�W�>y�hH�����NMV�X��|�&���4�j��ħd��9PJ�WiC���"z�z�������n�0z���q3��:i�L��C�0��JI$Y6���bQ7V/~��	u�'�$
d��c�b<��A��h/��p���*O\���G>o���s�M�v" ��T"O6� �a�/�-�$��,&�,p`O�h�EeԹJH�X��k��Cr��P��e�<��D�Q|=��1)�8��GC�K�<AEJ-0g�����&5�wCF�<����.#���aɧT�
��Fw�<ygŊ�K�P{��:U��Y"��MZ?a
������Ī"	�ahB)N����ȓk���#��?w4�0ҡb�r���OTf9b�L,D� �B�gAB)��TU��J ����Y�� �?|����Hf���D�6V�����6�ʵ�'��������ђ�'
[D��f�?{���D�����:V�m��N��a��A��&�����p>�U�Aey�iݨ v�8k�#Es����'d@L���m��3W�9k����'���"bC�$��"�b�f���'Y���Ak
,pf4
�.L[/f��'�(3��I2k���;D�W:�1r�'�����]�ճ#��SU�1�'�eT�a�ā+3�˰R�X��'HN��U�H�+� ���.��_�����'�9�%&�$������!6NQ��' H� ��c��k�o��|����'��٨&BN�kn�Z���K�1B�'�`��u�'s����Ӣ&c���ȓ~�4����56Q� .��1ͪ���x�p��F5DC���0��O��|�ȓ��0&�O���)�6N�,Z	�ȓ:�8BhƬ���p4�;� �ȓ+��E`�eK�/r�����L�~���ȓT�(�l�8p�� ц�����ȓv�P���Sn� [���33�Ԇ�2f��h�eQ/7��JԤ� wV"���1��3n�/Jϐ����8�`d�	`<Ƙ	ą`�%G�T�8��a�<yPٮYn�<�Ɂ 2=
P#b�Fc�<y�f�&o?�X��Ι]����w��]}b�)ҧL#2e�%(��G����EIi!���ȓ�⥉�"ݘ;��ĪS�ߕ����?i��0|�pj��cڄ�Um�!=��H�A�Vg��hO�Oy
�IWl�l�Z��P�Ɍ#��a�'���4F�P����P��"w}��'�&��2�D�.���� (_!���RO��*\������n5�-��AkH<)vg {�l��O�6��`$$XE�<I #�EyR$�e�gZ�%:V�	~�<i�%D�i�v%���`�\�9¢�|�<��F�0��G I�� ���w�<�#���o�F��!� �l��Ir�<� V�p�,D+bru��ęWҁ)�"OX�b"�V( V\�2%@�{�VH �"O���Fmq^�� bÝ:0��dr�"O���F�2J+���|xxL�����(O�OQ:�H+��a��-8���O�=E�Ԧ^� ��:!m�w&v=��N��y2��͚��I�0`�H��X	����O8�"}j��%T�@�9��ep���E�<�a�]7��a�Ǉ7�Ha@��}�<y�)�/>BPH��=�f4X�K�x؟��4��yV�I�!Jp���jF?�@�ȓQ����t;bh!=K�$@�ȓΐ����	>��0��&\�  R��ȓY�8[a$�z����a��(@���?�y��	7^��eK�'?|��8�E�-��doӄ���ݫE��-�A�ׯ ]b�B�Ιw!�d��y��
aa�A)��C@J�!�$[>��	�D]QCr��@mA+L�!�d�$����H��=!2G��i[1O�l�b�S�'zt{ׇ2�@i��fY'Q��ی��s�hT�Bˎ4�t�ڣ']X�zW`;D�����, ��Ǫ��+^�1��9D�DR�p^����M
���#��)LO�듆������u+󇃳^_Z�b��؝8�}2���5Q�Dz��˽Rf��@�#D��9���*g��Xp�$�<Q�@zs"D����R5��1�L;K� @H�=D�x�dO�f_N!���	�0��ѭ;D�8���߱dq~�`UOs� T5`չ�@)$��"ӢW�%�֭�E3$��ظCk;�"���0����OP	���:C?�p�F5RM��'łD1���< ʵY�'�y�(Q�O�d(���S ZIy� 	�&�,1�m��/�ʓ�hOQ>2�C2��]�A�!A)J�#0�I��p=���"�: $LB�z��i��_���<�Fڞ���PDCU�U��lJ�O&*ޚC��:�<5�&ټ��c"YV����5ړH�b�B�[���� ,߯|�jI�ȓ;I��sd�g�!J���0Ū)��;�T	�*ʴ8/��)�c@�(@���<8SedWA�t��_��lҳE%D����E�K�� ���� C�l�@qA>D�l��JV�bfA`�ߘ�
LR��=D���ݗe��M����<�u��O<D�$�F ��T��@��  vш�9D�8���-5�H:�F�o�r��4�4D���@��f��ذ���� ��*ւ2D��`�ʱx������(9��9;�+D��P&����A���G>U��q���(D�L#^,>���@œՈ� �#D�,·�ܪm���K�R%ȸ�$H/D���d��+��8㕯�h���ce�"D��R��]DQR�|�$b.D���� 5�I�g!ː+��Uc�%,D��K!���=��p
1ō���M�e=D�d��@�s�n��d(`Yą3@D&D���@>;DH��']���9��9D��QW&�K��̨�J]� CH4*�8D�H�KK�BI,�뷋Z�d����Ej!D���2i����pp'l�S��*2�2D�D����-:�.��Ш�'Lp�S�1D��p	�L'�D�$ �.>$L+��/D� @�c##���m�$Sj:P���)D��(gf�&2�1Ҵ�YX p�N2D�� �\�"�]ĈQc�O�J��LJ�"O@- �ۦK༨#	[ ~Z�H�"O��	�&�6Cg������a���"O|葑�Ԏ��':$t��"O0�����w���0&\��	�"O8�)W�T�6=@(4�
�oט��"ON�9`�@Wjd]�SdөTw���"O����x�ԕ�rhJ	��"O�!aLY2_�u`�3�n�a�"Oh�ia�¬f�8H0���X�Z��B"O�|�U9�.�`�S&��@�&"O�!aH�<S|<�S!�����V"O�x��+E=.�a�2g��d��"O�� ���!giL5Z��Z�i����A"O,aҦדa�N�,e�m�D�֮�y,���ʳhO2iJH��y�
�73P��4A��rxD�%,��yF�)����ρ�VS@H����yr��0E�Y!��OMv���_'�y����*hfaN-Nxv88���7�y�Ɗ�Y#�(����:�R��y2���5z����g�/.�EY���y�J�=u��P(�!(��"�����y�
A!W��As-��VH[�@�y�$�h��
����X��p� Ŝ��y���+tY�hҧO� �(�!A�ǣ�y����pU�qQr&޳v��yы�-�yRMN�	�4dI�Ȃc"����U��yR*�*\�Zl��ǿ/98(hg�U��y��ڒX���z��ȉ��q��­�y�f@�Y�Ą }8���&˒�y�D	T��+�+��|l�*���y҈YN(�Qg�	ܢ}������yH)@�F)��*D���ѡ���y�㏵3�H��RCC�`I��꛵�ybD6K[���ci吕8c�Z4�y"�E�7����MS].\�������yb�$�\qi�D�>Nf�����yRKܖ$U�9�*	�2��9��U�y"�׮]���6�T�#6��,~��ȓh�(�A���}�F.�*cj�l�ȓ-*�����,�Fx��C�	6ތ�ȓ&$v���-�: �X#4���&P��ȓ)S�� �.gv&(���>\����x �Ȅ Q~��a��K>lt
���k�j�����!>�^`�g!B�2�ȓў��Q��ku0�H'o�<{4�ȓXF`0�EJ-l�Щ(�N?: �M�ȓP\��j�3tb��vθViU��?)���J+.x�qդҳ0۸���/���s�d�0�l0�6�0$���ȓ@]�bm�J܎x!)�O:���l�H�1S��5'2��Y���8��u�ȓ WɁ��B5f�!R�D?/ֈĄȓ=���" ��|4� 9#ָ�l��Rs�!���)�V9ZfB�8�݆�y����Pƒ-!.�i��d���ȓ^�[�*��Set���B�u�N��8.؊À�Y`�i!��F�"�~i�ȓnD���Ɲ��,<Y�hT9��ф�*t��*WJ��=?r)�tb�(D��Є�f��b��d���H��)t�Zń�BT͘�cƷ3�pXé�#[�I�ȓLt�� ��Ӷ�ʜRt�ǛJs�M��S�? ��t�� ,�jE!�#�z;TE�s"O�!��Y��v� )�<��"O����)�`��� ��Y"O6�QF�\B24��ą^�w{�Cr"Ob-	�k���̍���=zeҬ��"O�p��$U�Rd�c�͘�����"OH��G��44���	�� ~v��"OT���LJ&.#�P�4蟉klT�R"OJ!*��?j�<�6lQ�Rg�\9�"O����Lí0�td�!�v)�c�"O��s��^�����]!��"OB��.ֈz�`�N�!��y[�"O�Թ�n�wM�y��Ȍ	?�I��"O��;G�ٷWl\��-k8��"Ox�T��Ho�I3���)J�"O���˛�K'�r��'^�yI�"Oh�0
X�K#%N����"O ���:�Ru'�X#�p��"O��ӣH��m^p�ːk�2y�~���"O5� �[�"���X�i�v���q"O�|X��K'���a	]�3- �(B"O����.,�A�s�ޅl5��ZR"O���jP0f��&�-# ��A"OnE�`��?@�EN�^��5"O�A���,ɞ�#cNa�"O���]�P����,��Q���9s"O�ű�a24��H� U�EF�!�"O܌[��6�Tл�,^}-��"O84��!m�ttRDLG8`vt
�"O��c�� 7��X�aP)N NA3"O�\ʶ�O- �Љu�	���"OJ}0$96��쫥f��	|��"O,����ǕG4F��hCLE��"O]��"i��%s��`-�d��"O���GL(W�$�j�@�!S(�d��"OH��� :�*��P��@��0r�"O��CA�G�zeޘر��/b|��"O�IH��ȯ-�jL �˺lXDI�"O0t;b�=4�X��Bi�w��]�e"O���#xZ2\ٕ� �w3F��3"OJ���)�0��2���D�:�ٵ"OR "F k�:��6�d��82"O��`��!����m_z�4�3"Oh|#G/]�&�
�P�j�Lk�e�R"ON "�Z�
�����9.� �"O��R�!6t������^"�dsC"O���F�f|5:�"覩Z"OL]�M^����� U�m�B��f"O��b!��	ytrA�����V�4"O��FO�*U�2ik�Μ!	�rԡ"O���0��^n� R�_�R�X�"O��3Rc�F+\$�Hf�py��"O���7꒼`"�Ką' D�u"O�9q�(��Y��u�P�?P�z5AC"OP�yPk_t�<`"CJ
T�)St"O&v���>EjI��K�WP���"O�\q�(G�{v8�1�0VeR�"O.���cÂ}�<TÌ��+�p)�S"O����۶�Z��j,6�޸q"O�u�@�ho�!AA�C��tx�P"O���s+	`� \C��.����t"O��`F)�Aॣ� ����"O��tn�]�������MԖ���"OTԡ4��'\ƺ�s�H� ���# "O� $0�G%��Av���׋J@�z�"ON1�@�G,IL���ӊ�: cR��A"Op�B&��>�`�`�5zЕ�#"O�QѶ��P�" ��l��m�\c"O�I`I�!1L 5���y�����"Ou��Δe��$IB�?C��*�"O0 ����?$��@���/6.4bR"O���я!r�Ґ.��>�`�c"O�$�C��6s�:���#٫
Zz�1�"OX�y�`�/�������S*tا"O2%�f��/[PY"�P+|?.���"O
	:v��:)b����($���"O����N��5���� ×(	�hI"O2u*�N�^�rh�Nް\�2�`�"O<8p���H����D�Y��9�"O�s3#� \F�1�� Ѵ���"ObxR����]
�O,m�R�q�"O6U!��H,E+B�3�XQ�=j"O��(sNA�$/���$�é �T��"O�I��I]	%�8�`��	�r�5"O��#a�#T��LҀ�<ks��ٳ"O$b���s��*4a�<	��%`%"O,4Z /_�c��� ���4y�p|x�"O��xF��i�����طPf~��V�<��S'��0��E,6LQ�ęT�<�C�
�FծiA�k�7옑�7�H�<)�P�V̖!;�a�%�|��aB�<ِ"��k���%�7��p�c�w�<����|���1��j��P�DL|�<)�ǉ�a|8H)��c�hp��<�b�^��z�kƮ�pv�<PS��P�<yPT�e�< 3C�(\TD�l�P�<�����14R�6�:(w�\�v��N�<�#���{��� P�N<%�ț��o�<ɔ�ȁ=�ɑ��w6Y2iOg�<� �=�����	nd]0���|�<9'k= ��UY/ԦL�/�|�<��+ޔ?�4(P5�п S�-(���v�<�K��r�d8{A-��mmRf��M�ȓx��3D�ͯ����Ӧ&^�L�����)a�_^�D�W!8A�~�ȓc��1D�݊>>h�[�}3n0��p
& �QL�X�������"k�Ї�'q�"敽{�¡�#�Z?�Շȓ{��cs�Y�����2�\��CP�ș�f�+c��y���C�$��ȓ4H@�!d] _nZt�!��<8P���O�H����EO8���)\!cRN5�ȓXvF�3��V����K���0�ȓ|s�t�T)�?Sܓ2�Y��v`��V<6!BWhS)���)����b�=�ȓ4H��T�U� u��	D.ȭ�tL�ȓ�L�bjV�|�+Ԫ�L��$�4D����yJ�cQ�=�Z�b%5D�@[%T5|����&�b;�%D��r�!	�p��!S��7)���ck?D�| ���/TA �;A�G�_��]q`h#D�D���o~~��D��(�v��?D���h�5v(�ۂ��,�@)�6,=D���,�*ʐ#�ʞX�1��N;D���#Ǭ�j1
���*{Ƣ��@9D����\�BAJ���G�&�F7D���E�4]&pP���_es�eس.4D��y#OU�j@���
=zm��GG6D�� �ᛤ�Ơ( ��QN_�P5���"O�"A�
4p�.wɤ�+�"O荸r�
l&2��c�&+��|��"O�iA�n�<[�*i!$�����dR!"OԜseŅ�&���q �|�$��"O�	y
/0�H�k��Z���B"O���g��x���Iv��4�6"O� � �	>C(��s�B�cq��"O�U����
m�y��Ō�z�"O�l(7M
-fDQ�Ed{�D=�"O�e�_���a��`����C�L+!�d�	�����B���=��Ϲy�!�dE�^�@C�`�,m��yç���P�!�d��I��x�b��{��ɴ�֙^�!�d��p����1M��r��bjʊ<�!���)���bW��.[��큵��/�!��G/"x�@cp�� rF�B����!��J\P��W�J7<p���f��9c@!��/Z�P}���[#-T��22Nر�!�DF�"���[>$X�<��-�-m!���ki��Ö��1A�\1fM3|!�$�iw\����=-�4ٰ׬27y!�DL/cp�+A�S�S���""��.Jc!��+F�+u���g�`�:2䒳Y!�$��8bT 9䖑Hs�@� �!�$�&��d w�ŭ%k��C�ݭ�!�$E�
$���S
L��� �
4e�!���oS
(∊?@�k4 �Z�!�D�n�0�A�`3@Z��V�ە�!��Q/nz��[�=H�ju�@�!�$��J&VP�)�*򲼡���%@!��׆WJ~ɐ6-��>�R��t���C�!��; M�칔+Ǘa�i����'�!�$[�!����Uz���*N)L�!�ă,qy�8���Κ~|�lztj�=I!�r��"$��x� �S)�'`�!��'�D�Q��?x���C⃧Y�ޔ��'�����&��٢�JB�v�B
�'�� ���ѣH�F�5�Z���'��+"Iӕ;T񳒴���Zc�<���'�ʵ	�HP����G�H]�<t���bfz}�Vٓ,"L%1�`�[�<!P$[?a�dt����!
��$[�<a���W�| ��
n��ey��QB�<�%�ڻ>��]@������� C�<�mO�8�x��ӥr�ջ�B�<�d�^�P�:r��n�dh���Sv�<�c��e��� ��( ��*��QZ�<Q@-��{˴u����̩�sFW�<�E��=L �	%�U�P6���O�<�C�Jɀ���TRzI��cBH�<����HZ���TN�����M�<��fd��-����s/h*#	H�<ɷ�L]Z���H�~tɚ�Nz�<�� �sh4�IG�~D �rȚs�<yRG�-	b�Y�����7�����e�<���qd@��U'�� M�p��$Ei�<IR�E�L�p R3L�?AY��f�<�G��?��Q� ��9�X�@G- ^�<� L���B$f��Ahc [�<A6��x���W�
2�H�A
\�<�`ˏ��5�ٲ+�ĸ��'[E!����@!cgσW����E)��!�d�& u��J^(P�h%h�(G,!�� n��ec�C!r�
9p��B�"O��K@�ߺ���xF��?�� �"O��	�2}Ό|�b%B�5٬��"OB�q-^0'%�\K��!��"O�ɒ����B:���P��� ,b�"O-@��Y	rf9Ӫ��viL���"O��"�,ĸU�
HSoJ D�Լ!B"O�(�����\��ct�5�<9v"Oց�G�r���Κ�>��t'"O�� �Ø+��ٱ�mб9y$�q'"O(u��O�2������7P=L)@"O��c��Ǹ���y'웂9�Xܩ"O�<T�O���21�_ %dޔ��"O��1���Г��2Ht�""O��򶫞����G�$)%�m;�"O�=�醍V�����O)K�@��"O��@M F�ʱ��L?"��"O0pѵ�3�v��E7�W �y�F�c�6i����,�,�[!���yR��2dv$���k'O��!�V��yb��&�֡���+}<�ءC���y��O @d��f�
�_a����y"�0p���rW����DE;z9�'�����EcG�	��&��9�6�1�'�-Ck�nA�}��3~��J	�'�����D )���F`����'�]�RA�MG�B�[ -M�U3�'!$��*�3׾�F�*G�$��',�pC� �ooDًDdS�"��X�'����Ba�7=Y�{�ML9�y_=c�.��v��6�]��)��y�dN�Q��ɉ�$]0'���¬�2�y�OU��E�Q�%V^�Y'��yR@�<q�L���S�����Ҁ�y�m�[����u̠K!z���yR� m��q�����h�`���y��	����,}:MC#�yB�?iW��SshʅWPJ4XA�M��y*/!�0A�(�9]��d��KP��y��<X�ç���C!� 1�ybL#I��]yd+T6 ܭ�ϓ�y��,x�u��#*<�u�P͒7�y��!N���� *�0%��Q F�y�힇V�`,�qA�/������&�y�f�!z����`�Îd�ⱙ���ygŃpvd�+��_���c�F���yBO�0
e��!��ºZ浺�/���y�@�,{�����F��VT��e��y�
�4�����S
R2�<B"�ć�y�*
� ��1D�Ft0á��y"�C..�*l{59:&��s���ybd�0_8
=���$q�MP�gU�y�N�-6������^�S�D �g�"�yҭV�Oz\��ve��Ly�`3G"��yrm�,5��D�Ё�ڤ�#� ��y�.��+o�٨��c�Թ#n�(�y-[6Kn��S��W=��(��y2�j��_�%oܩ��C�	J�n`&� K(E��/��~�B�I8\��;�g۰~�)�B&��PA�B�I+g#摓1��=l�,���A��LFC�I�,�PxCmەd�l(t囙'nC�	�F��P�U�_�N�;�hY�6�C�=.����)c����F1B�)� `b��&������;�4�s"O,X� �H#d<؉�吔
X���"O���j؂}.0i���p䰋�"O\���N��i@p0q��]/Ix�"O���"g�I #S�RD(�"O�D`֭oz��B��O�H�u"OvI{E��/1!X����'�*\�b"Obp�`)�	Hx���H�ؖ8�"O�I�b�E�mH��1]�#����"OB��G3M���t�ѪW��K�"O�".ϰ��ݚ��G.�(��"O@�g[���K�/�I�.�;�"Od�+@AQ$k#�X�G0�v�#"Ov�#$͠,5�A��,̿a�deyD"O�	��!�[��i��,2/�ah�"O�L�qϊ�.�5Ѡ�I�1"�\��"O�A�V1p����c�9U֠�U"O���&�νCV�SVM�$� �"O�PP�%
N��T���x����"O\�gj�A��B�`ƐI�����"O�i"ϤO����&	3id�b"O��&K�`D�(C�BF�p"O�ј�&M*��dd��A� a�"O�}AS��nZ���,nh�P2�"O�0ڀ�Z7. F�@FJ��`"O&�`U���m�򴢧ռ�$��"O�9�	DdM� ۼ�:��S"O�t	A_/#7D��,H�Y��mY�"OnK�L]��n�#�-&.�3�"O����M"XTBy�-��s��"O�r'�_T��
�Uo��qq"O�x��I�Xd�m:�nU�9tp<k"O����M�roz�Yc�6Y�h�"O���X�ڵ�l�2}C��"Oj�@! �Y�4p���L�{.J���"OJt��,��E�s����%hE"Ofxc��X4M�\ٲc�c ٚ�"O��R�	"7~b��1"�9L�@�"Oz)��䂡p���1���\"���"O��ѥ�� �^��D F:=g�:�"O��!膄gT�4/ʾsf<�p"O�Y�$U�u�_"!j��"O�)��bZ5$~Rt3��ɕ2L"Z�"Or���-@��JX��ň���d�C"O�9Z`�~� �cN["�l��"O��`�-����,x{b�" "O�l�viI/D�����{u$���"O�\"�.��xgO��(g"HB"O��H��6X@Ҙ�.T,9E8-p�"O̵�7%Dw�ʳ-�C��"O�%QGIU'}��FܫMB<d��"O���'�aX�)z�&�?B��PG"O~��$5�X��%ɣ?%Nyp1"O���c�K�
���S,'�4�!"O�,��K�^mĚ`͒�M8�"O�i�W	�K.9A'�V�m�*�y�"OZ�Ek�0M��ܳ"���&��"O�ыwd�#A����.^*T�\` �"Oz�P�̅/4���`-���Li�"O)8e��!Q#��9wA�.:�ܡ��"O���Vl��r��)C�ۻ;w��a"Oh�	ӭ�<2�^|	�D
�h�h��"Oe !T#A�j8Q��Ed(�q"O|���J$@�r�Gʦ|�4y1&"O� :�0c'�E����2��5����"OL�8��WQm��Ă�f�x�S"OĠ0����o��Hk��A&���s�"OL�)fd�-tŬ\���аS;�9u"O��3'ȇj��$(d�_�]h"O��x��L+IAlġ�Y�
�JLH�*O�e�2�Y/1`�1�`eʁH��8�	�'FvpX���'��8��A�A�$q�	�'!F�ʡ�ڏ}����fZ?x|4�	�'C��bB��#��p���!	R0��'}���ˁ��-p���zxH�	�'̸1C��) h��e��X,�	�'�D�M���I�I5��'�T)���+,G��1QfC3>����'��e˦I��jĬ�x0]�4��Ă�'YP�0R"�;N;��P��R2ܒ��'�.)(��?7r�0^&y8�:�'I����H^N������!�&�'D�Jv�G�,2�(�e��F��d��'�>8#%�%wAQ)���>�����'��y�!��W�l����<;��2�'<p�#S�;[:�m3�剩^T���
�'��	h��̄l�v��7-��*�uI
�'�4-D!��Jw42�[mcF���'�92�CήP=�p� n��QH�'m�p�b�3~h�FO6\*4��'|���V�Q�z􄡻'��f�Z�@
�'�VP52����^�8���'���b��/��������W���'�s�'�7f:`�+����6X��'��=�F�ö{8���k�8K�ޤ��'��X�'
O�r8"e9��M�Y�T���'l�{���" �8ҁ����k�'l�(��6q�Acǟ�}0T���'U\���ƴ¦-)�M�t�.%��'׮���܌
���f���e;ht;�'����O�o��а%��c�,D�'��(��P�8�}*F�F�a�tk�'��U!���<
.1�vΉ�X�b5H
�'��D8$�ތA>�X�.ʕV�.l	�'� ��G�����D1L�U����'�b� 1��('6!��H�,M�	�'�~4��+Κh ��¿C����'� �k��)r��Qd�W�@xj���'#�3cc�:#�,�t�!g��a�'�v�j >m�����C�&_����'~���0@
1Ǆ�3@���R����'�
���Gx�*m��
O�Mߔp`�'����� � x��F�|���'���!7$�tk4:�T���'c��� +^�N�{�!`�x��'�Bz3E^�!��h S@`�B*�'�=���n4Ip�L�?\���*�'HmB���������TZ�Ҩ�'g$��ƀa>����
($׼���'dzm����e���(ݲ���J�'�p8!1o��z��@h�I��'�X�<��@]yRC�m��q�:|�d��V�<q��ۧ%R�Q��ɇ^ �43�$CR�<	J�0��V)H�-!Ċ"�b�<���`�鰬��N��^_�<D�
A;(�V/����$�Rd�<!#�˷#=ΰ�f�m�d�x���b�<�U����𤈛�}���Q�E�<� nu2'�բ7��m�7�ތX�L5s�"O,(�`cPN)x����W� �h�X�"O�(i%(N�7��as���5�*�	$"OrE��eG�[�r��v'@�f�1�'"O��WM�th�z��!-�Ȣv"O��ƌGw�Kʚl�F�@
Գ�y"Jl�6ٳ'$�lLr�K�h���y2e��p���Y�ɘ54��8cC��yr�^}1za�`R�]��`񵦟0�y2 ��|�b�����9������y�` �/���W�VĂу�iK �y�d�L�B�0� �P��ѥK��yR�_XM�|��J�t�tG>�y��N�d4�d�Q͋���%�N@��y��Ó58��05����,��yCE����
6!�X@G��y���h���� '�2!-^�y�eG�ulΐs1\v���/��yR�яV�1���辀�@&Ϗ�yBG
�״�Q6�W1E�H�v�L��y�H��o�j�[��E�}Q.�����y�q�<�rХ�(:��U�Z��y���8L����F�&�@��꒍�y��Zc\00�
�$���lʕ�y��x��5�c(��F�������y铋a���S6�0�ܴ(��X'�y�̸&��{�h��r9��jI��yB�P�`���ڕ+��]E(��Ŝ'�yү�P4�R��
3N���@d�M�yb�����Q6�M^��|����yҥ�2��-T���4酪_��y�'ō3Wti�Ս��4�v���y��I��zsǧ{�fA���8�y2�ɪo��v�k��������yb��
�(��f4Z\����u�<���3v��H�#��W�n�XAM�<y�HC�e�f$�@cHN*m���F�<��L�b�\Hc%
R�$��%����B�<����?Q�]���Ө��ư�y¤	�T�`��I�;#vy('ML��y2
Q9pt�Г�	��Lڶ�F�y�DN0���V�":�mF	���y"hͺi͒�HF��*�,U��i�v�<�T�χi# A0E�(���@ª�s�<i��ʡ .���Y6�Q��Y�<�voE�XTfQ�ơq������S�<t���)(^=�G��=��,ZA�P�<i���3Yഀ��E22�F�@�<�4�ڢ2���K6,Җw��h1AAy�<�F%.gY� �0	��5���$�Yy�<Q���DZ��B����L����Zr�<���K6<KP#�`:�@'oH�<��#OA6���C	4J����@�C�<����.m��l��莆]OR +&���<�B�bZ��ƔҦ&�<�J�{3������uf\��@�y�<Ae�Ao�Ѹ����[3���t�Hj�<���G8��q�w%J��I�+]b�<�P�\
}��B�K�f�Bl�H�<A�`�Jk�AQr%�o��,�r�D�<����@����E� �iL~� �}�<�Α�x�0P6nJ8kQ.u�ƤYD�<q�+���A�w�2m���D,�i�<9B�F.h!�8�Õ9Mn� 	�Xc�<� �H+��&{>�Z�܃B^���"O���Kʿ#��l�WeP�.�e*�"OpP� �<���O�{�D��j�<Y��L�M�$M��΄�6J�� �m@�<A1Ŀ��8�(dp��U�<9��;L��$2J���x�%�Bx�<�BH��25�BNk�&I{ԣDj�<���Tt��ð��4��;GFh�<�/Ե���q�FL�k �鲁B`�<���Y8�.��vH�2X֩��)�q�<)a#�B�脁FL�7���W��k�<��?}]�T[��C��F�XS&Sd�<A��Ǉk|tTs6B�y<�Y���]�<��ʄ3�A���Jk�2���Q�<��+��'��'�SI�|�hw�<��!�y�~!����<j5�Y���	s�<�MB)4ڕI��9MJ�KDn�<9��=q��sU	2,����Qo�<!!OE(K4��/�[��C�<��՘0<�&K�g�dQ�r�t�<�T��C���S).l�P0��o�<�/�Y[�\¥K�����˖m�<���1Q�t���[��|#�
A�<)uCE�RRd �p�h �@�<a�DE��r	��F2���ʲ�}�<�Ζ7B_���B`�I��z�<�Gj�}� ��S��I�� S��{�<a�h�%y��ĝ�fp�H�Ujc�<���ϾP��Y�p�ć��l��$�t�<!fC�<ke����a��e��l�<����%Kl���W��p �҈�r�<��!B6�l�����Qִ���q�<�R�W��,�8ROт`�6����k�<�g,E;� Y�-Ā}�>I#B�k�<p,��;�h���X�J8�rF��}�<�����	��5�['-K�Ճ��Ed�<��S�.��	�4����d�<���_�(�����Mڪ0��"�`�<�7ԼrEN�ځLSA�L�o`�<I�C�A�z%�
�8Ǡ�`��p�<��_Cz��§D��#�����Οl�<�����P���Y���#lm"���Kk�<��H�"����0%��R$@$
g�f�<�gC�4=�qC5� d�qhD��e�<9慈p���I6�J�8�t�{�/�c�<�f�l�`@�mԽ	g�ID\�<���׵{���h$ 1*�ç	CU�<��C���+5���,9n�O�<��MQi�D�(����3`�V�<ioA�9ZV���Kk�u���j�<��2#��H�1IʗC5�-� jj�<	�3�T��$B�=같�6 Dp�<�g��FiҘ+`�ԻA�����nJS�<���J�8>�b�u�p�Z�m�M�<A��0;ְ��䙼[����]p�<IcM �k�@�H4�ԵE�����n�<a "��}{P�����@H�h�<����4B��#L�39��[��L�<�$��ee��}	�Eq"�^mx!������� �W"U��iF.*O!�Y��@d��WO���!�N�6e!�\,��]b�c�	/c�!�$�Z�u\!���@\�2Ee�%/��@P�0>!�DD:#9������6ވ�g�H�4!�� �4��?nC�M����`c��""OP�@�i?~�i�$��/R AA"OBͪ��	d�`,ѷL¼kQ8e��"O"����X���<��A�N?�d"�"O���F��tN�`�&�Q�m�"O>x$Aɿmܮ���$$��*�"O�$ؠ�Ⱥ����0c
���q(�"O��A�8{��T��� 2D1�S"O6,�S#���#t"�"r=N�
�"O��2 T-Q�H W�b,"�aP"O���Ԉ&d@h��D�>]�R��"O�)�K��E�;�e���K�<qe�R���ɵ�V�Pa�alJ�<� ��-�m�������+Gj�<1u�ɝ7/��2#��C�@Cy�!�[FZ�У��EVy�AM�Gv!��G�m*��ޝC���uY�9�!�d�otb�L�7�\r��+�!�$�u�"�r%��&�AĜ5�!�D�/:v�!ص�
(u�n��3D�!�d��bc
 ��%#G�}	$�ʾS�!��"Ӵ�[ �D'	����%��;qA!��~ZN�e�1~vf�C���Q!�D'�(�a���vO>�!��X�Z!��=�F�١��mD9nv��C1"O�b�%V}��m��Y�o��I�C"O~�(e���SE��nx�8H�"O�-Q2B�.Jmbu-�p2�P�"Ob䲷dȞ-� ��N�	f"�I�"O^�a^{�B�x���=W�jg"Ot{F#�T���a�B�J�b��`"O~��
 d����c�rt�Ip"O����ٜ��1�TN�.b�2�"O��ꖭ�!"%\]�'e�${���f"O��:��$jגd%DK3V�@��"O�D"�m����U���«F����"Oy+�b��E���H�4YИ�"O4p
�K�:g�n���jWIc�{�"OXx�g�Ȩ�`�:3*�`
��"O����C�}��nO�\�`��"O��QV��]%��{�(`V�pґ"O�D� �Q u6�e�N��  "O�I@ə�P�)��}��"O�j��B=Ǭ�	E>h�ʼ�R"O���� I1�5HŅ�9J�^��4"O�eh�KL4W6l0�J֞|}�0�B"Op�8'�:n�����	ډ{j���"O���Íty*�B�Ŵ}��"OF2� ',���i�&�]����"O�P1�OPPtQ!R%C�VJ�H4"O��s @E�O��҂Đ�|ޚ��"O"��ࢊ�ɒԑ��G��^�r�"Ov�'E�U	�P2A�"��%yU"O~����Z��*D��kU7"��u�F"O�W!O(N�a@`@.r�,5�F"On�y��[�r.�:I�'�(�0"O�г�(V�\�!{0hA$]s���"O��! w4�1���-F`���!"O�<��Q)9�&��e��!V��4"Od�Ў�s�t��E�Y�Uڳ"O����̓q-ۆ�%f�,[w"O�D�4E_,��u-5Bel���"O��T��,|�
�7�F*�\ #�"Of�ɡ#
qt\��t/Ms��Q""O� ���!ZSں�jo�;*-�hh�"O�p��F&��Um�/:1ِ*O� )�	f@�)vƙ���Ա
�'=l$I�(�����jUKP��>��	�',l2�ϗ)"�a�'+��Sg<�H	�'��L F�
���}ٷ)�~߂p��'�N�(��%q'��
�=0�'WL���6[@���cK<{��p
�'dJ�q��42�$p1bό�$���8	�'�:��i�&��hR�%�1�8��'t�LHFUso�����%,���'�0��Q�99�(���(���'�ޜ��@ڟG�6�%�WdPX�'�P�[�mD�`p�1僇�(p�'!<�z�_�t\i����B���'���W�~~>�C��P'z����'pF-��]��~�7�
 �QJ�'�Msg&P"����FB�%-x-Y�'�ԩ��GI�T]AV
B
SvK�'S�L�V' �w=L�� N:��;�'r���"
�H#$��ҿ p���'Ƹ�6��iF��A�wl>%H�'�VU���Y:=�$U��A�7���'ڌ��VIڲ0�V C�R!1�8�Y�'V�i�@�'L�4�p�C�'�p��'>��r��A�tIb�Lеj��k�'��ʅ@����p�c-ޟf;xtc�'E�1�'QRh���1ZM�@��'��3u�C&��uAq����j}�
�'	�0�e%��<�r��]%F�b&"O��:������b��.*��xR"OzQ��勧@����p��"OXD8��˦E�Ht�p'�i�D� "O�\�0�]1gqx�����Y���"O��Y%b��pPqg �&�4�x�"O� `q��X�~P�V��M��!`"O�i�0˅�b�("�����"O@g�)���ƈ�.(c�Y�"O~d;&�N�s�Xx7�@ ^J�!��"OXĀ��=e=>J�EW�]?D�X"OJ�Ud���p�N�&u^��g"O�h��&�����ϒ SV�`b"O.m#������W�B�N���"O�4c�˞a���!�W:4J���"OT傢�D,8�����.bM�$"O��17��� n�� �K�8y$���V"Of	�P�@����:`��f�!"O�Y�5�2�B�⁯�@Y�Q�T"O��)��3�x�'�M�}q$]Br"O�8���ұ~ڑp��ƊL^М�E"Ox�:�_ ������B+P�H7"O@�x�/��u�r`��C�L�4�"OtQ`�aˌ�~�92oI�C1��s"Or��w)F'*|9en�k <�SW"O�����^¶�	��5R�]3�"O��ac��'��eIJ0kA����"O���F蜍|9��P&UFd�Ʌ"O�z璣{����eҠ+�nI�""OlPQ0MU�:����f؋K�*���"O��9�i���|�
!F�;E�xYG"O��{�$Ӎ7n��c�{��� "O~����rZ�\Ie"]p�l+�"O���E��""���,1�.P(�"O�(㐉V�Ve�ԿI�pu�W"O� X1�D�g��=�I��];L��"Ol�)a��d�N|)Ө�w��<�7"O���Y(!a��"��ՆT|�25"O���B���w��1�[�h�"O�AC"I�0ti�򧀇OR��� "O��7e��)�p ZP�׻p��7"O�i�'_b߼P�P�E���0D"ODyv��4E����D� ~�lP�"O�Up��_"vhH1z�^�~�Ř�"O��Aᛵ;F�Z-�h�+g"O̙c��O��� E-�r� �#�"OP0�J׼)de�6#�;bZ��+v"O��Ks�F����:PK�$d�5�"Oj���J��(�*�*ERZkd"O>I���ēO��\����RR�Y9�"Or�+VN�o�]� �&5%�� 4"O\źS��o>0j��J7-�Ј�"O��3P�Ό%��081)��6 ��"O�8�ÏGH<��S��0�� q�"O0DcglI#-w��f�X5�섹"O����61��4���8X�n}K�"Oh�kg�J/ ��y��o�Z�"O�aq��bH�]��N�<����"O:��M¿9O�;�n����;`"OZ�T"����ㄮ��� ##"O2��KH�1����WΟ4�p�1"OBdR7�p�.�H�Aة}����*O�e ��ã^K|���D�N\� �'����-K�	`q;d�� �h���'/F�J�aN*ar�{�/�}�����'5(Vnʰ]�u�r�X����C�'O؅�ƠJ4v���C�L�1
��Q�'�� qO2�J�#�bZ-���s�'-�U	CƋC�[���- ���'��,q���mkbD�a���(���8�'���L
ad����! z`!�'G(9`գ^�#X6u�g
��h�'E���U����0mr���~�����'�Dy�ED�Zmv ��D�+���z�'�"�� �SC-t���OZ�#RҀ`
����c��Oz,��2'��_�b���:D������|��� �:U^̳�-D�0*4bN5=t�����=�\D�p.6D� x��C9&�,ो��"�LZ�i8D�̱6	ѩ_4ű�����	R�5D�QQ�� ��C�Юú��u�/D���g�޽gG62�c�� �Z!��,D�ػW�ݫa�z�R�,�T���K)D��Y�GL�<�l��#ѥm�)ڲ/5D� Y��U2u^�4��?�L�cTJ3D���$H�JTn���͵o����2D�P�E� �NQ�1�
L�7ؑKGe/D�Pq ��Q]�M��圇+�X��.D�4)����O_
Qs��etҩ�b�8D�T�Ca�)��@���
6^�͹�C6D��I���f|��� Z�v��03D�ly�Ō<ND����"\"�%Ð�5D���$��>�f���#l�$�i��5D�舳�M�7����V��>XƾAZ��>D��zg;|�r��1��,&R0`&�;D��hQ���<�$S8��B@�>D���M�ڭ�Vj/}�PZ�9D�0� �%�p�:���1�DJs�8D��h��Tc�e땅�*���yQ�2D�� ����_1W��E�7*�;0Z���"O��;���:@lAʃ��3͐h�4"O��s�k&qV���H�?(�KR"O�񰡛�?蔩a���.��#3"Oր�G\3q�L-𴣓�i�~�"O�#4HL�2b��(#����B"O�\�F�	�}R��[�
]�(�n�4"O�AE�C��P��蟡�X��"O����(Y � D������"O��K�ij��q�@�p��L�"O��1�W!U�Q�b�?&z
ݩ"OƼ���4.�N�*]�|a0Lk`"O����.y�D��CPH��
�"O
�:���Ed� �S	 g��ce"O�4j�,���b4�̶
�L*�"O&�b�iN0lŨ@/�'�8��g"Oԥ��_�"X��m؎1n�u�Q"O�Hʐ�E	�tǬR�B��$'"O�d2��� �6�C��*���Y"Ovl�L/?^	1��ǰc���ٱ"O���nB2eY a�(��hҊa�"O(�
d�Z:G�bA��6j��Z�"O^�3��I+pɚ��¶%�xy)�"O&`�g>D����X�Ss�'"O�H��A�%��A��F�Wj���"O8e	���VϾHʱ*��i3!"O,=
��Y7늘 �Z~�\��"Ot�)P�ܘ}E�	��aȸR�^��"O ��j��aB�!��oPx���$"O���c�0W�����%B�*+�$�"Oưӳi�&�14�%:�r�ST"O�H۰���86Qk�$�)�vX��"O��sS��y����#ܗ5����"O܀!P�4(���BR�Iu�@a�"O������
V� �Qb�rC9!�ɇ2&��iU%_3#�Y7蔑R!�M&Ѩ��dNI��)�']�;=!��ƺ{��qiF2opX �g� G1!�ġ@��k�ͷ9c�u8e�#!�!�$�s��Pۖ�L3ETpE�D��D�!�ݙ/�	3'�Ƅ��|uO��g�!�D�rc<�9����b�����^�!�d�oT�|��j���Jz�f�!�$^� �p�p����C
*_!��.(��;v�W�b�8��2'�!�#R�ȱ����:�P*���*�!���;)Pd�hA��<q@� 8�c�q�!�Ě�hq�s䊐:?��P���!<�!�D�1��H�,�v�b�E��e@!��H%v{2})����m� Ev�8H!��f�Kb�R:1u��ړ�&%>!�ٗ9b֑0",�,5o�9	���2B1!��S�&��D8sK��n]L` ��D+�!��M����p�b$�yd�ϳ,2���Ji�a��7_��E���ϰC�m�ȓ]M�����Ws����(Z�R��ȓjhp}B�Ɛs�
����m� �����i5b$;��y�1�qZ�0��EX�)s#\�I��#qBH
�h�ȓHT���FP.������דk��\�ȓO����Q�d�Pb���H%����[���� �[)҄�Q�]k2������j���<]rh� ��w[zz��ȓ=�j�K�<t*�*CeJl��S�? ��� �\C�������)c��XQ��'T-̓>tXB��=W#����K��,(z��ȓ�5`̋?R"!��
�+� �D|r���o�<�U��`a�VC�0�B䉱]�N�z%�!a������F�M�
�?!���X9e�@)���Ts��WAW9V�!�$�2P�򴁖EO�zi��.V=p���\��H���Xb@�<_ș��)��7��Q�"O��JT���9b��L�\(&�xR�'_���R�m�&����
���b��hOѰ�"�Ff��������A8�EX�p����I"��he�ځus�A+�e>D�8ԣ[�*� %"��M��jAp��<D���ډl+��7��7"B!Rv��<	���S�Pf� Bj҉~���J�eV�.��B�I�.�h�G�F�fS6%�u�S�d7��O���dB.nVb!+#�܋J�^�) "]�V��Dy2�z>y�&��*�j��a��/��+�(D���fƀ�jdj��V���0}��d�Oȣ=E�d`�`ܔ�S��/��]�Ɖ^,.!�O�1���[�&:���q'VK!�$�j�r�jd��V���s��.��~�]��{��΄jf����@�ȢŦ8�Ds���;.��f
L-�J��t¾�zc3D����V	(�XX9��W�r�!�+D�(#G��i��t��M�2Yhya�'D�,���,CѼ;f�9[��iv�y�D���(I�������|1�]�V��\���d �I;1�
����0ܰ����S�8�C䉝f0��H�Ae�L:��Ű-��c�hoZF���'HX�3�G�` d}�a��z�M�ȓNq��*�a��r0�!�iY�k����.�́SE�Ņ9���㊋\��Fx��)J2��	1��s�ˁ$/	Z bR��m�<yI0_�`���-�!*��r��cܓҰ=�� ^�N���+QQՌ�A��JX�<��Y��Zq�����r������m�<)���5�]Ȁ/A� ���*pM1T�x#bLJ�M̜�&iE�W� �CG�g���������1s)S�k@y�VJ� �!���RJ6Ƞ0!J�>���sSi��R��$/�O�$��&S�/��8rI�i��A"O!��C��P�h���\�P}+��y!®&�� @��T�lj�e���y��
U^�Уg�5e���8��Բ�y���;�NpAbL�[�^M{��_�m���G�Cc>ҧ�g�R��,a�&�H|	�t�V(|�q���|y2n�7"�*�(��'.<�P�B�ѯ�y�iFa~��X�`�D@�_����!���O�c���O`h$3ԝK�ݸ���3xX�c�'Jhy�҄4ft��VY`mX�J�'J
�yì���~mYgE�R�&!#�'��qz�&�b��1Z�
�` ��'����1O� t~{�N�Q�����O,�=E���p᤯Wf�B���X�SP8Ĉ�'�` ��3O��e@��!An^=��'�N���s�>DɤM��>��@��'v�85��1�� ��H>�2���'\��4J�5!�1���0��=:�'{l�b��&"�L�S#��4t�l�	�'�v���B��m�x��+�3O"8"�'{T\�f�����pDC�����'j�)H������fǼ<�\��'�j�d�\�p،U���;Ag"�+��� �#v�O�y�l�#��~q�(#"O�u"�.�S<�� ��W��i��"O�	���+zE���@�T$m�\;c�IMX�����.m 8� �'sjYScK9<O�#<�u���
�� K� ;�T���%���ZR&X-S��{�O�i�$4E~���L8��I�J��3�H�T��]QB�	/ ��&�2~��u�`���AB䉭_Wd� D\�h4�<��]��C������g�S�=�XX�L��#<َ��?�k��\��7�_��ۆ�9�T���O-��:��9}�h��H?"��a�'��Ԏ:��i��鑘�J�;�'s�0�/�T��sLN�NzN<������cZQ�`�{��_%N�ι��	��e�<9BH>4������J�.�NP*tA�o�<�@%E�s^�(��n�V���Dc�<�U㜨jG�j�ZvE"g-�\�<�p��K�4��CIW�)a@���U�<ɳHeZ�!5�@k��LS@#�F�<��N�8!|�{�']?_
(�I��W�<	6+������
Lxa��V�<1T��#)��W��?R�(�s`�~�<1A���tv̉"�[:
T�I��MN�<��f��R���Y�J5�u�RP�'3�?9��JJ�n}���I�+�@�	e�3D�\#cJ�mi��3h���p�r��Q�i�O���F*AH��ɓ�Y#zM��Eqea~�V���wN^�z������#i��8K��8D����`Čغ��p��-3�^���;�~�O:�mD9���G�'w�H���N�C� ��g�R%�w$�!xb`��#T�� �ȓ2*�mqp���N�21��3�ԑ2H�#=E��w���0č�U�!uh\y�B��I|�')��
d.�7���[���%�8�{�';a��	d~���Q�Ŋѹ�o���p>1p�>)����S�@�ՠD�~4E�2"Yh��|yߴ��HV�H���I�,UxsI
68��=!����$;C��ElJ&������ G�O&�=%>
U@C�[��G)�Na�#2D����nQ�ce���*^8X�T J�1D����dJ",�nx9"b�]����b)�ObC�ɱs��a���V�0J�x1��Ox����3����*�h;��Z�:=��Ӂ�$|\!��I�� ��BG�0�%�fS�ct�O*��(�)�	ɵ*��̙�ҍm���0�>a��|F{����e��a��� �-_��@�In8�t��;4�R���X��M(��<D��X�!�<Lזpwk��ԩ��.5D�pi���K�Z� �5��x9E�0�Ԩ�h� A�˂_;`x���2!t���"O t
�C�/c4�"�O�-1��Sr���0e�)�'GG@�ɕKӮe
pQ�l�,76��'YR"=E�4�^OL���1��U{P�b����'X�h�뉟f�s�����2�I��c���Ӧ��%�~��z6�џO9p��Wb9D��c�݆Fʺ��E�I#b0:x�6O�=QFA 	(\E�p��CTTk�5D��ѧ酲u��8����)vo�1Zŧ8D���%E!/���	���~Vh!��5D��F䎕5e�A[+��ԥ1D���L�&2�Ġ:3�7L�J9жb5D�x
Q�R�xe�1��M�v���(D�����D}8���NשT��Y�I3D�� ��H@&X)f��I�!D�(kv�"O�|���8
}B� � 5�n-��"O ���A��~ܼ�b�DT���"O�+���
&�+gğ�T�T�1"O� b
��<�TmUdܻ��5�"O0EⰢK�P�0�� =��7D.D�t�h�+�� ��ŧ|8*�b@�*D�P(��D�,�l��� 2���+�).D�xz�)Sq�6$��+��o��Q���-D�̑����f�Sr�M�x����l&D�ȊBN�?~��;�K�3M�޸�`�>D��*q��  ��%��ǘ�ш;D�T�u�
�C��I�R�����n<D��(���i�.����Y
,R8�Db;D��(��GJkT���C+
����V�:D�@{`эav&E��_1��%'8D�H"&���|��]�w��y���`�C"D�����E#`�aQ���,P���?D��3�ܦ?/�q宊�[<a��%;D�|�u£f� �"2nF#L����`E6D�Xc���M�F`l�_�p)q��b�<� ��d���J�d�
`��e�f�Y�<�$OF�`�P�C���|*f�A�U�<ya%��F-�q!���J��h p+�O�<�N��茳��O�%d�aдe�M�<�taE�o$>\ T^^�LyZg��J�<�We�x������d��A�p�<y$��F����GB\��E
f!Bi�<9��ݜ�x���Q���{��m�<���@;��I�Į� }Jrl3�Rl�<���j�b)B�4�ĳCd�<�u��>@Ơ!ħͳ%��9�$IGI�<��ҏp�
E�$��A(EφM�<�����g� ��Û'V�*%�g��D�<��6!���wJ]:^Ft�O�[�<@�S�G�>����t����(�{�<��a^K�q��.��-�RtH�H�m�<�`��dJ8}C��s�i��Ij�<�v,W�c|��H]�U������i�<���CU}�LkqP�tU�(j�b�^�<��/�X'����)�2�qS��R�<�7NЈ7>��!�+4@)Vk�P�<���G�9u����d�<Tx�i��$J�<a��J9Xø��ʞ5�>��AF�<i�,���0��Эي-R�騑,�<��m\�t(�&<qe�O�<��A�?E#$���11L(�f��E�<Q���%��eJrb�"{�Њ\C�<$��I����LK�AL�Uc��V�<i�C���ؘ�IM{P	�TO�< �ۜ6| ��gQ�����O�yB��4���lI #�`ѳ5Մ�y�h�%p`�ja�A��1� ��(�y��ݬJ\f̀�"��H@����yb�a�-
V��~��m�W��&�yB�[6�J�2��rM �� ��yM7Q���:`�@�q�^���ꌒ�y��L Y`����x�b��yb�͆y���KQ��Q�A��d��yBM�q\v]�A/�,�t��y
ՠF���0Cσu��p�M��yэ!ˢ� ӯ����hQ-�9�p>H<��Iϭ�\�a��Ӈ(p�f��^x�LDy��%�0q`�_�.���*_[�<� �����
GDD�"j�[Z��T"O�@�ק���	�FɎ�I��l�qT��D{��I�YX"��|� �Q+�6|�!�du�� ��C��0�@�k���S�!�$W
�����ԾWp�0@-V1e�ab�O�i=���rA��+&ll2S�$.\Op��.%�ļ*##gUp�@�O��$�oZ`�#F�ǽ4K2��v���|!�d�/��@8Avy�"g�!�Ē�K��!��9H|�:��?�!��M�\Z@�w͞;Z������|�!��x��	���@��E��!��	_�~^�l�晗Od��筇%&�bԃ��6�IN�'����^���j@bv�0(t��
TXk3D��J!(g�e@b��o�I)�O3D�,:�$���0Ӏ� �sꄙƮ0D�L�%�ނB�XcF���M�5��c���"~�I'�h�)'%�h�Ţ��-ycB�I%Z�0W�4��+"�7���'�4(��U:D�J
5g}�հw���/�J��mm�����:lҪ�X@ώ�d�ȓY]V�J!���U_D����2
mGy�|↧�o�X�	�N�0D��إb�w�'���S�|�V�AC���J�P�Խ2٤C䉞Y�vlqlƐkn�d�RL�/l��D(��&Vy\�Cc���ެ8V�N�w(:��.�$�6��x�`(IhQP�B���{�a}r�>ѣ��1x�B�PF���j��DY1`s�<iU�&8��d!��K�8�����EC�<iN[:m�	�å��<��s�VA(<a�4h��쳢
��z\���^6 j��R���	��Y�e~NM������,��l؅X�DU�uK���E'A�r�`���f9f�)�T�z���j��лa�P��	o�$�,6DD�%�����ҬT�&�z���gy�3O�Qh$��=	D�J0�Ɏh��� �"Op���`V�����p�<�p�d9�S�) e��&@K�9ȩ��C��O��C��w��ITpJ�"O
�*���K��+&���S����'�a{��O��Dʢ6�j��ջ1���Q�)�<#&��}x��0,B�xx�y���0�&A��%��ȟd(��@�(�������1�L:�"OJ�2a_�r�`l3���.�XY�"O�94�p�����F�ZM�"O`H��gM�[��l��Cʸ�"O&DIt�Аc?*��b���h���d�'�I0e��Ka�/<��+��S��D!}"�>%>�O���Q�ܟ`3�����V�D�2�S����G�4�70� -�զ_�IR�D��D�y2� �U
� 2-�/H삑cj^-�yR�=�R>ሔH 7X����u&C/gӆ̺�$�>��q(&Msp+�?�&��E�	Ss�0�O(��$�o:Y�G	�&U�JL���
�]�a~��i��ā�/��d����)�b]���r��Op�=%>���n�"�:��n��l�(#D�hBK�?�l��BAH�hK�@�4@>D�X� �6 Vha1ɚ00$�j����D{��i^ n�:%ӑ�+��4EKZ7#�!��)L9�bJ�',��@4�W�$�!�DQ,I�����=Jm�5*��_�!��ٕi�
%3��-ca`���/��}�!�d�$n(0͹P�^�8�C�ѿi!��F97/¼���!��P���7�!�� ڤX�Æ�eY��Au� ^^:e(�"O�%�a��8�*p��H�,"���'0�S��y"`�6�^Q"���oFlPw�=�y�I	�Kh ���h��%���*�y�!�)�2��R�X(Х N��~��'*QI��T�r��dp%�r].�;	�'�X!0�MS�6u0uǅ�^�����'�ː�7O\��AA-mE�Tz	�'�����FnT �bd�\���'g���6jϨH� �䊣UA�\�
����2 �Ei�.�BRb`��J�_Q!��zg��(�#8#4���IȈOQ��EyB����qd�5`�(D�:���'D�����uZ�!��P���iV	$D��3p�S�*��9�� �/^�ʓ�.D��"�� hF���`�ۄ]$�!X�
(D���T"�	a�.���%p9R� )ʓ��<y@��
 ���"�3H�B��jFGx�<�'�B���L���e�	�X�@�H�'~���JZ�Z�iiւƤ!�RI��'��)S��P���,O>����'�Tы��G��x5AO����3���:���� �v�M�)ˊ�* �Ć�
5��p���� ����[�f���s�nǴ�F%�-D�DiQM�6F�ʅS��R��?Ke!�d��`c0�95��,:��z�h�v�F~2�	�u�P8�!�;�T�y�L�mu C��+q|6�arf��'���
�Ë�`��B��TMT(�T@��[����$ߗH�!�D2X�� �H7b�*����ў��	6M�5Yqm]�uQ`d�5,�����d,�s�"L��ȟ_a!r��[�f�ҩ�ȓ�����R�h���1b��9�?��7|�;@�;�P�ɤ`¼�Z0��>$,�m��i�B%�p�T4d:���<'�8k`	�~�(���I�(F~��|
�d�n&x0�ӨH"=�4�j���`��I�t+�M��@.�@� рW5>NDc�TE{���A̜a��T�f̽;�؋�_*��xBdHL�
4�G���02f��'Z�c��q`I�Ӻ�'<Ԡ@K
>���H�F4R��'�d\x�ꌹ-$!{2�ЄV��1�O�䓏MK`�Q^ܓ�~�'��)��޴%�*9`iV�R`E�ȓDr�x��
l
ِ�Bض)��<�ȓrV4c�CC݋բ�pZ���ȓ�^���2)�kf�Tu��ȓy��w }<�};ֆǗA<��ȓm�ѡ��%z'��jAB�8Z�Y��&����q̆�Ҟ��$E7t����ȓľL�ҡ�+�X5 B&[�J��O��=�b$�	ef��ph�9��%�C�YY�<	$��/S��]Y�IK�u�p�`�*T_�<������}�FaM":��x��B�<	�F�J1���
��U��M��IB�<�'�n	�Hr�����%�QE�<�fbZ�,�"���螒(H��QD̓rH�Fx��!-}�JuV��.e�����S��y��
%tU֔zs�P�1�
U�q�R��O������Z*���Z-��AA/k!�d{��]�g�
2��B��tVB�	�V�lA�,��5�Ԍ��Y0gA����,��Pd�� �n�^�pǋ�4�81�ȓ~���XR��(i L��D4r7��$��D{��ԆQ2]�p��g��ܴ	� F��y
� �}R3˂�0�Z��'�0D0p""O��pW��=���p��N�X.��d"O�h2gN�D�r�0f��]��mP�"Ovy��]%N3V��2E�0���P�"O�I�7�I�L'԰����'@�qH"O��R�Z''�p(�+�"I	�=c"O��ŌQb+H��e�(�;�"O� +�Q� `n}�ǡ�H�Ft �"O��	�NT�@H����7br2J'"O�<�����=�&�2��+]4e3r"OzIbWf�a_tr�掼-pZp�"O6})��4:\0Q��mm�ى�"ORDR�@¨J	-��hC1P���"O�����ґ,�L�A�kz�c"O�E��M�_��dӠ���8��"O6��Ө̺_^��3�\ ��S�"O�ɧ��a8�A��͂�E���y�"O�U��i]?f�)P���-ɖ���"O���
���R5ѵ?ٖ �"O��r3�/)�f��6FY�5��� �"O6�0+I�"]f��% 9�LM"O������+Sf���Ƒ�� �"Od)�'�*��	�5�萝�"O���薿��Mz��͇P�h���"OYp�N�s�,�zХ��	�fT!�"O�)#×�?� ��F\�ހ��Q"O+�6�R�SCcH6��� �"O� I��:^L1sr�Q�70�U	&"Ol��Л�E�ঌ;U͞pQ�"O�!X�	�V�d�`��=_'BВ#"O\̻@	�*KX�JT�E�q�!�"O8�q�C�@�@<��۱q�Ti�"O ��IL�Q��� T�7RZ��"OT���F�mҤДN�dNr�""OP���J��QL;	=�7�44���L + �8��֍s5N�� �"D�@B�J,༩�q���fL��#� D���h	(u �T���V0x�8y!�"D�0`�F�:%�H�0���t<���� D��	�#���3�C�6o���� D�����o(����%Ab�|�U?D��`���' �B��D���k.D�S��Ғf�����0%^Xt�.D�$H�5����G�8��C&D��j1�������'f��<�̻p�'D�d�v+�+8D����b���D#D��P�Æ�bQHDAH�-5���"�:D�����];v���BiI�!��%��%:D��:�C��ZtP�2�?e*v�$j<D�43���L�r����?D$mxRh6D�d���>0l��Q�oB~z:��T1D���w,�
F�#r�B�Q�V�ʲo5D���)C�t�6Y�U`�S
�1�B�1D��s
���L1WnI&h��`�(D�(�ZȖ&Y�Ƈ�\`���7�'D�@�#T�̑�7b��-td8 Ƈ"D��CAD�=ne*����*�B�I#IR��!�(�!MH0�	ef]���'�"��EF�ML��LA �
�'�)����P��D����@@�$0�'�N驁�>t��m��f�r7l���'��uAqf�^ℜ���!u��'a���M֫A5ڱIJ92���'�<a$�ĬO�1R!gJ�,������ XT��!����y�c�׬"T��T"O.0fn��t8��@5`��L0�� "O��b�H�w����%*r��"O��	��X�*�c�ΤR�i�"OH̃�GݴBO�c�*l�2��w"O\(��"��7��H�6NI1S�
Cq"O؅IB�Y�kƢx �G�b��4"O(4'䚠E`�t��i�%~����"O��x���\j���0��X��0{�"ON��J��:�4!�]e<���"O�1 � �M�.�(���>�Zu�"O�����7��i���|�+�!���KK���F����֌ 䫉����$	�����maA��C�2#2B}ځ:�����@%x�`!�+P:5�f����.,O�t�2����
�6���$C�w�V�I��$7�����f��Z�E[�/Ӫ��LK�X5&�X��o��qO���@� �?ܸ �FŒ�>���"O�S2i :9!�$��E>� �%.�ɣ�\���L<y7�;x���ڗ�_��P8r��RH<Y�N
g�<y�D-�9�(zQgң8'@� v�3�O:�`�F���ub��͘F|R�b�'��ӴA[��?;�2����C�+մd*�ɄPB��,CC^�!�M]3c)� �Q!I���O��aa)�)��_���Vg@R,(ӧM�^��C��:�N�c �F�/�H�Y�ݬ%�C�:e�U�ꀀ
�	hv+��)%�C�	?Np�ۄ�_:=W��C����C�I�n�4�I�c4�BD�H�wԀC�	��C���/�4  �%ɗwYbC�ɄI'|Р��1�ޡ����Nj`B�I�>��-uo�'Q9j��a�N�uDB�<2VWaZ'�Dh���~�dC�IE�r|Y�↦nMղ!��r�LC�I=G���s��4}[.dJ"@�/ +�C�I�:-�ţ��;E�:xC��))/DC�ɓC�Z��GV�E�����-�sNC�I�r�V���|8�!��2+�jB�I�8R�m������p�e�XGhB�I��1'��>~3 h��,u�*C�	�b��k���r���P4j�-j�2C�I�dtȭ�s�W; ��[�7(-C���$r�A+��hD2c�B�� =������/*�Yy��D�xB�IBE�U	�ާnʔ���5�*B�I�@�<����U�iX�u�J�L~"C�Ʌ%�^tXR.��Ƶ{e�.�C�I�JVx����<7��B&B�Qe�C�	9��J�D�mP��z�D�<%�C�	�{]vM;Bj�;���[��I�6�C�I@�2�Jb*˩
��1��n[ g��C�I>+���hQlG�I>p%P�D�rlC�ɴm%��r"mő�����H�e��B�,� ��d�^��Tbc�#U��C䉣��4�5�(B�L:�Ё;��C䉓,.t4��፰9�b5��ɐ�͔C�I�k�B��El[�?/���F�9�B�I?J��\�B$V.���A`JO�TòB䉻&��l�C�z�L���ʆ5��B�+��!�7��\��%8��Փ/&8B䉢O�vḵ�+4e���"/M�fs�C�3|)�x��&wzztj�b�*??`B䉂S7~��Y�I�qX���,>HB�tT9���B�p.�q�(]�+D4B�)� ��[�f�[��=�o�qbڐ�'"OU�)S�14��8�m@�&id�"O���e�K�?_��%R�U2x|��O����[�3���ib�E�b�~��#�)M��C�I� .�%i
�f�sBe�M����dN(HQ�<S�ؓ��I.i�l�0��#[����B�Ca�C��=�b�,M�p��	�% �<n��4gƩ:g ��Q��çQ
P�c�$�U��r0v<�"O| c!o�[.ĳ��[���3�M���ɭe���*�� ��g�(dd}���Og���fd\�
&hh���	٪����#j-T�9�G�� �Na@� �	;�2(�����zö�'��#&bU:`$���
�s'�	����B9~�N�rw,�^�Y"�����A(?�h�Ц��!O�R7JB��y�/� 	�@�Z�Z�rՋV�P<vY�x#r9�p-J�8�zQK��ה|R�~�C��B,�� �!,��I�'�^L�<��G�R4L��`O�jQJ����lw*Eu��>-������$�ɔO���rv��)<��bn �(��@&�O*�!ǀF�c}*-1�ә_�((�s!K3����Tۑ.��5L�3:������h��KڣfB�ȋ%.�1}�ў����%^���&�=�r�#",��|҇ˊQ��:��<�.�*@(�h�<���� ����B�7��h3�埘O[}�>D	�
J3��M����Y�Og��i�gRY�>���!b��x�1"O�h�`�}`R�C�a���Dd��:��&�g( �C�،IH�SX�'ˠtrt/��9Z~1(`h��lB��@	�lA��x1,�%A7@�����Z(��6˚t�fh����E|��¿�0>���D�r�J��ms0�[|�'�,�M��@��i%�D�\�?�����M=yWl���ėæɨA"O&0+w���*��[�&N	�ԅ�6�'V�����=Ad�l��k\
i6.<;g�ӕ�"!�園t;<�x��,ĢɆȓK���r�K-c��hsF�(nz��įK.e��:�LN�5`���6G�l���.I�.�z��_�[��`��tDa~���: |Q*F�݋Er�
�V�X��+�aJ8'#С`�ᗮB�d���W���_9�|E�g[6F���>q`�n�M�#%|�mk���d�#+�@0�lQ*Ak��q"O"�Y֥�$�(��Z�&�Aq5P�DU ��.Ҹ!��hJ� ��?����P]�|�@/	2p.�̨� D�l+&�׶C��6�	9���l�c�z�'����F2��gܓ1���*#��3MG<��#T1_,�Q{v���@`�����KB�BJt��`h�	��#�!� ��K�BI�%�V�~�&���%Y�qO����պ$��@E�ʔ~�D�8�"O�Q��J���$;�b��y�(�R"O�Q�%�K�ۡa��I�� "O\���~��JՊǫ}eB��"O���(ťM� p�q�R�5g�@&"Oz�{"��P^l�C�O�yW>���"O�iƆ�"F�6�ko�D��#"O`�Zs�/*��IPN��H�`�"O��rw�R�eւe9�o�o�b��"O`�h&g�!B�hu����x���a3"O�b1@�IG�����3JF�8w"O����_���H#,ٲw5
<�"O���/M�|���n�d�#@"O,��r�K�X�
�<h�J��5
� �y��_c�-a�N�?�LE�ŕ��y��M-����,4�n%a�LG1�y��X�.]��Ǫ2'��u(3E
$��>�`�J�~��
�f��S� �FD�J�n��y�oVDg�l�eB�@7vt��� �(O���ň�Zܨ̼3�f �A��}��}��"O ��h�j[.��tg ��L{V�?��X�����OH����y�z���l�:\�dM�r"O$z�搵O��-�A��81�R����O�a����p>i�B]0lv�2��>9r���SL!�O��9����y
�  ��J�$)����МX\���"OƝqa$��r>L���\�0#��ɰ@
ȁYA�S�yQ�� �ȃZ��l�a޴-<C䉟o؆�����2���B��OA06M0��"~n�(��9:Ƌ�RUX���}FB䉁����Fډ/T �H�O�@���ݹ�h��6Cï`v�0`f�</�!�D��2L��Z5l
;RB1{���(�!�D�^/�]Ps��Ad�9ْ��!�!���!��Q���'+`pك��Y=�!���zIJ���Θjb,�Qッi!�D�7+GP@�mJ� �<!�@���PyD��%2y���˃Ɩ�97����yR�
��C�BkQq��;bf]m�<�UoZ=+5��J���a>��'Ia�<��j�!S²@B5 �?7����Åa�<a�I�����1	�.?Ɲ�B^b�<�aW����*�	�PR�&�c�<�F�=�|q�K�>��$c��Z�<�Ɍ����1M�qz����[�<����f�2�nY�z�h��S�<Apώ~
2Ap��	��<x ��u�<�REV�YȒaC���5�
��p�PO�<�G?@PaɅ�N��;��E�<ᴍ	�[��)рL)u�9�m�B�<��׽x�"f��dVdJG�\|�<i��M;r��ICE�t;rtj� P�<	��
�(Yy�_�F��m����L�<�BB���lC � �Q{ �r�<ѱ�\�`�l�z4�_�s
��2��T�<Qt�7�bIiuEݚ	ɺH�t�GS�<�¨A(UYS�͝d��8�	N�<�˅_b��C�@��0�⏝H�<QT.8l�>��Cҝ*$�kv@�]�<���M�P]f��V�ܘS(���0T�<Q��I�	��pc�.>�\aCg��l�<�1��m�NY����9��̪�D�G�<��`MF����lȉ;=��CT�<���E�t$j�
$pQB)�\�<!�,��(���ED�x�f�]�<'hCo�p�r���\�"ݺ���F�<�̜�a��YdD�jͮ�B�]G�<�E��p��%����8�%h�C�<��%'TT `#RC+}�h�r�<��Q?ZDK�E bR�Q5�s�<��,��$E��v��:l����Nl�<��&T�HF�;Z�HLi@�v�<1��?jF��:�m4IbMr�	s�<QЏ�Hp���DX(=�T���n�[�<Qv(��Z���Œi�������i�<�E���ॉB�L�jT��I�f�<)���oKz=���5+�p���^�<� �]H2�p� DԳD� ��X�<���T�TTp���?���맏�Z�<1�i�[��pf�iz`X[�<!&��sQ`*wÔ���t�Rύi�<��e�.3Kb�9seP�@ɖ�:w,i�<Q��Ǩ�����x��ܩ�NDN�<�����W��t𰍓�X�8�I�O�V�<Y#Q/;r\���	.Ѯt��IPd�<����dx�j�NN�!���u!�`�<1�S�1�����E2��D�6�PV�<1�m�$��p�M �`il�_�<�a��J�T�[.L���*�n�<� ��ӂ�-V�~����d�b�"O���Gمv���@�^5�F\��"O3�}�J�`%^*:��i�J3D�`��f��p��x"�j��>�j�A��=D��P���[�ʁ�ťI��($�7D�<�T-2�v!�p.z0{�mݨ(�!�*� s��9/����ñ^�!�d��)ĭ:@ D�j�P:ej��7�!�d��gkZ1�"�K*DX��8`�!���i\(S���:s�~�Z�k�-|�!��G����P�9F�`���5w!��u��P���(�-A�hI�Ov!��H��蕩	7[�y�&O�T!���d��q#4��,1�@��	
h!�$��h h뤏K#1��T�ǯĒ�!�x�uyp�بK���� .�!��J*3��4�Rܻ٘)Cfnۣ"!�䋣<����a#�9�ܽ� � �!����΀C�Dĝ[�^S�JE%�!�d5E���"��Җ�Z�A��k!�$��o�r���8���k�'� Q!���')���E�#s<�2Ƨب�!��uǬ�fٖKt��x� E�q�!�X9vj�,��K����3��>y�!�D�4��ȊU.��UpT� �)��z�!��K#\����ǔ� Ƅ�(�J�%�!��@58�V��H�� �Z!Bo�F'!�P��`@b�J�ĊX7�\�1!�d�D��=��á�ֳ7!��"d�~��G㑥R�P8�F)D�!��C"�`y�%�f�URb#j!�d�/���`b��c�  rcT�TT!�$@2b�eI@�#*d����A϶!V!򄜒j���1�?h>�t��B!�����E�b�6�.e!'�U� G!��
�.n�u@�9m��
�斊b8!�$G0I�zP�V,#h���ER}!�$2�&�P��5� CB�^�!�d��=�D�L�)(��Uc	.v�!�D 2#G�YQ��n��f��9!�$�2��CjL��樏�!�/ɘ�Y�gۅl�`�R��?�!�Ā���ɷߑ_0�1R�+h�!�DH4J�^�0��>� !��O!�d܏O�<�&f�2h��:v <!!�� �9�ǃ��)��M��ڐ�!���wWz�	��T)3(F��/�!�!�$�H�"y3��sH=��o&0�!�$�F��U��H�2����F�γZ<!�đUz���,�j�v,��*I1�!�d�nh.ظ0�Y�Z��ȏ�DO!�D��?���q�͕��,�b��D�w6!�Q�JjX������@IV)Dz!�$�&+�̨������ʅ��
�!�DLT%���ъ��Ϩ!�=�!�$��:^�����<C�(U�t�\��!�M�P?�y�L. ���0�^�e_!�A)rNVh����E��I�����E>!�$_�Wd|��JU��V�ʱ�P�94!�d8,�Z|raMir�T
�X!��? �H�W$�V@�ʴo�Y!�D�����z�(�6R�j.� F!�DIG��� ]/H?,���
#!��	V�p�agG�	?!lٓR��F+!�� ��{����7�Yx�	����ذ"O<	��@<:�qj��F�e�@�˶"O.ar$˖>*¦�=���3G"ORHb��IZ���@�r�jlQ"O$�;񧜚�V%�C4��"O����ε�:8�BҠF�[�"O|�#�@ӽ����Ԫ\x���"O��Z#��ص/E,�9�@"O]�0��R[�A��n����� "O���1 &6� (*��P�^i`�"ON�I匍0@B�4z�e�=�^<y"Oz�� �_�R�����T�^aY�"O���P�[(7��ɛ�	����D"O�H���&��ѩ���{�0��"Ot����5"�nT�`LaU�Ǿ�y�k��6���Y��̓$^�\�3����y�l\������ʖ4 �z	"�����yB��r0����8z�`D��#�y҇
1u
�i�/Œ1A�(K��yB�4>c�UC��"n��l�gǉ�y�HX�#���$���J�d2F&�y���~��Qa�hG H6>0I���y�#�L:X���ã8���Ȅ'ֿ�y�-[fet|`�	@0%�y�����y�'�wYRE��LC(�2p�f�ղ�y��Ԏon�%K�)G�,(� ����yI��j�T٣�)��>Vz�t`�5�y�f�
h��BA%(� ���A;�y�ݎU�:}#�(�$(̺��A��y���q��1�8�� �G&�y.�<?^�P�0�-�}`TBB��yr�
4<�RW�0f4�p�b�K8B��:V�B x oT�)��c�A�:+B�I���:t��01~����a�1��B��
Z������q����
�T�B䉱6��9dK�L;��I�M�++_�B�I=��@ �N�t���������B�I�\��Аn 6g�2���d��C�	�8������b3w23�rE�8D� 
rL_Z�:�y&�
4.t`�E�6D�4�`�8[���IBpsz���>D�,i���8[�,;�a��^��h�aJ=D�\����(;����]�1�h��DO?D����ő�m���i��ܴ)�t��rf3D���a��2͘�;V�8�jmi&4D�`��c�o*d3���]���؃�5D�L�Vb�6<��s2� }��YR�>D����N�-���
A�,O�P�j��(D��@�N--4A��#"H(����$D������>�LYp�G�
т�I#D�����M9[B��R�B�X��[Wo#D�P�Ќ�Px��J�G�X�� J>D�T��j�\��"���_;��	6
2D���C`Ә6O�\8�b��97j�a��5D������g�r]2��[�,T[�@0D�0�rN���^����4}B�9B�%D�x����9.Ph���e�R=��7D�[�+�5=z�3V�5w�6�y�'D�(*r,��7 ���ٴ5{!�%D��*���*S������Fۆx�@"D��0�h4B����ď,Z:)���!D�0�F~4�c�a�U{��	� ?D��B��=Y&pʁУrO�`�( D�H�@��e%)�N���P��>D�� Nu�%CK��:�K<kJH5j2"O�-�ve��N�`8Za�==6T�i�"O�q�r��
A�����|r���"O(����ZI�es"X?P�x�"OF)��	�a�$�HFa#)�Q�U"O���a�B2�(Ɂ�;t���"O`M�eBuX�8q�ЛL��f"O��`��*��B*�4�u�g"O:ͻ5E�*Q�V�C5)��~��r"O��2�,Ԣ�x��A+��<�"O��`B@��&y9�
˟|��h�"O��	��:b>x���	��G�D=�w"O�Y D��x]a@Gu��"O��X�OK�O�9��F�b���� "O�l��'D!n$a٦��$���7"OV\9���*H"�ď�1]�y�"O��7�	#?l��͌�AbjlB"O*5�����B�r��@� q`�Q`"O�k�MB\�M@	J�'}~��2"OB� ��D2�ݸB�E�>�W"O���pM�E{$���\�H`�Xh�"O���2�.tvd8�	"vPH蹷"O�e0HP&W�Q�ID,\�-�S"O��(�	��2������]���0"O��ѱ��'�����̖X��J�"O(�KHt*�����0>�:�"Oę(�c^�xF�UҦ��(a0B4��"O�x�m�8\M�Z���H8�c�"O	qD	�+dFā�
�6�%"�,�y�`KØ J'�	�D�֔�����y"��	'����ĤM�;� �"�O��yrI��$ ��C¬̷lt~a����yB�=_9��V��	Y��%��j�'�y2�O�7��y�%�G�Z�X`+����yrǣ��H��J-z�4���U��y��}�$�rJ��s��z���yr�HEr1 CCʮk!\A��y2`�J2��ԡ�v��3�gA�yD2M6���]�zV�Ð�yr�-G�LQE�_�GL*!����>�y�c (�,��\ 8�@��rI��yR�H�O�l)�2�=0�qp!IZ�y��,� q�W��5�"�y�	�Ʋ4�2,P7zt���$7>E��t�3�I�,0}P��B ��ᇃR94��C�	�ZƘ����v�.DjP&�`�C�Ɍq�<S勎/N�f�S��L'�C�!�>��b �"f��L�S-
�,�C�3@��
�B�(�4�8"	ȗk�(��5�ɐp�
�Q#��k'�@ҳ�ƈ�Bꓘ��hO�S:sW؉��ޝRH�UA�!�B�O�UI�����=l dӶ�Ϙc���g�M�2�>bQ��|�t�N=�t�	���M��P���P�C�)�![N�[�X�_���A	2���4��0|J !߸G��Iʀ�5�B�;���O�P�ti�J|�6MS�0�@�����[aM?y�	F�~BNUQ5�IH㴟Ę���w�D[�H�,���ĆJ��T���!��I�l'4P�?�g�Q�h����N(��k���5&�� nZ�|�"<E�D�ǇQ|X%��E�;)��E�S�ݘM��x��D.⧏����;%��{P�L�Rba{Q�TX��l/(�<���+(�dU %�\%b`�1r�|2�)�Ӡ [ؘ+��Ӎ0�Nq�@O�1q�V�ΰ=��'ۤ0"�J�tǢ�;�o�r�>mP�'�R����I� @����İgU�T��'A0�#qaY!!h0��Jܬe�Za���� �DJ��]8`���u��^�>U�"O��`$��piF%���N'�FѰ��>Aۓf?�3�L�7n�H�鱬æS'*	��d��#�V}'�P�����6D�y�1 �qR��� .���ɥ�?�j��`�I�x���+*D��H��A�{�����+ñ'p�q�)D�x���Ɇ�� "-A�T�d�xF2D�#���n$���4�&��'�$D���C�+q�� ���
��Y{7L$D��0D�!�H��J7ލ��!D��yT��!@R*�#vB�"��	8��?D���p��,����1`0�h}ӣ�"D�H�c+Z������y,9��K!D�<�AD4���C����@`
�0�+ D� ��RU���O��_a E�w�>D�Cp ؇Ps�� U�ܠJA��=D�Dh3銝)�Z	($+^�r 5ۓf=D�� ��^v�!�f�Z�����=D�\[���]���@�O��)܄�.D��[s���m�rAjr�ֵu�f��0k+D���u'��bڬJUK��mǤ`�T,>D��g��;�A7l�<Q_���6�<D�與(�#YV)��>�,`P�5D���/,�|L�2��/P`숧 0D�00�$�r�v�;���=:�D�:W�1D�D����I����co�2��ׇ/D��,�t��\8�+YH�$LӃI+D�@���X�N�h�&�5��j��%D�+B�R��qK���zl���67D���ӄҁ'(�PunܼJ6���4D�8����
u-el�|�8 *O��9�	�;q�8�A^!�i0t"O���4	�mAM':S�}�"OB�T�/ ����S,K/`Qz�"O��hY/�D�z�0v{a8�"Ox���˟ �:�H���5tZؐ�"O�@�@�^ Ox!��&P.x�!��"O8�ѧMH�B��$��Ç?\��@�"O@	9��H�t(&D=9Q`I�"O��Cp��ML���!wܴ�*'"O^lQg�A���"�3�f)� "O�y��M�O:4�ږ`ԧ�bQ�"O�H���^���+ �)�M	�"Oڑ��	aKPeq�dHsΒJ�"O�%B�����<��t��0hDc�"Ohׯ�`��-�C�v�J�"O"p��c�~�)�U���mL�� "OF]z%�G�ȥ&��`j�ar"O��$�]���g�	 p0��"O��c3NTt&���	��!�t"O��P��ҡ_��X��Đlɘ���"O�(�P�T!j�x�o̳bK���"O�`ÌUl�p��d��6U�J��"Oʅ��G��Z�{�π���9��"O��I��]
6�"����ޠD��8 "O"H��Z$[v@�2��M�i^��QT"O�p�Q�C�f�:4�,�aH�Qv"O�%j�4�&��dŔ�c7�l�3"OR�c4#6>��P��9{{!�U�\�u�0%��{1�Q"�_8h!�D��]�@�6�F�j�&�8#��*s3!�$;'B:�p��+���QD�;
!�1V��V�	\nv8���� !�'���1 KZ�o�	��-N�P�!�� ���W�\�}C��'&J9K\$i��"O1"勽m��=���܄P$yYa"O��1@�
�۶�ŋ/A�Щ$"O|�Cb��^'f�A���.-��p"O�U	U]�36�(y��5,6�Y�"O"��M9Y���;���E("O��`Z�;j�����L�+�"Oc��CY��a`�J:6t�!"Oބ"� �`��:��	Px�t"O>EaT��X"0�y2+�3,>�Q��"O�Ѷ�@�0 x�
��;@rY��"Op��*�5N ��x�*��TE"O��9g�Y��|��$��#t"��"O�i��C�-��@���UC^Ab'"O ��`�$�v�Ɂ�܎j���"O�A+w�:$bH���ފh�,���"OjIj���<A&�ЁMɼBOD���"Ot�1�o#;�|�� ,�O8���"O6�KD �8��({��@&7%�D�u"O���gK*����/1@�+�"O(��3;u���`c�;"N��"OVd���=����"��a ֔h�"Oڭ+bK�R
�P��J!qz��"O����X�U�ƽ�!�@�r �8��"O<`K�D��ܡ��D�d�Qr"O*L��햪\��|�#&__K4h�"O�)�4$:C	�.:�AG"ObP
�C\�B��p�W�J�="��E"O�T`EEݏ*�8�Xv�>u�p�q"O���)�0}֚��wㅼ2��ɃP"O"Q1�D(?��$�\�l�D,r0"OДj�LP�-�0�!ZRP\���V��y���\��a���o\Bm��O	5�y��		c���t술Yt����Z��y,΃hðU�m½A��t�v#1�y�S�O�铄`ĠB�D�p�F��y����?J�@�G�_0IN({���+�y҂H*4U�rA�6[N��	C�y�jV�kffU�p�L�n�ფeҹ�y2*�#n���Q�!<$���4��'�yB��#R�X�͗d&"��ÇI��y��Z���"U��c&D��O��y�'ס%���rRa���L*���y�$p��t�rK�\�\�G��y2���:����$N����V�T
�yB�8P �
t��A�h�Ō��y�b4�,��"e�4�%�A+�y�ϟ�#�ieH��Z$YDKQ�y����qnZ����ڈy�-�`���y��	�W�9�(� j n���/Ԫ�yr	 /6G�QY�Ld���!���#�y�G�ٔe�>]�0�" ;�y2%ж��bBĂ�Q�����1�yBGU#h��U"b��!��2ugH��yR��Iԡ��ß$�h1�X��y2!`�H��3����4r�aځ�y�W`���% ِWj��$I��y
��Cю�
�N�����d�ؤ�yo�0W
�|�
½2LX���yr�"S�� ��vx>��eO�y2c�#q2��.�Cr�k�m��y2ㅶ7~���d��c4�
t�K�y�J�)W�<�2��<��R㥑��yB�E����JS$t�+L:�T��S�? JH��)��J���- �fht�:�*O@��cOH7�Ha��ޝ ��8��'`�R�ؗw��qj�'Q6p���:�'�t��'g��|����޴a�\�	�'2��pL�(H1ĭ���(%��'j�a�2 �%E�,9�%�L֜���'�E�w��C���D���6�&�S�'��8���ӭ>������..)]�
�'��8��ҩFQ�􎀗(#h� �'@�!�
�354����S���(��',�Ytb�"dT�X�mΫ�P�P�'�~�i�'�GLVX s��)��
�'�8�`���f{V���K�H#F��
�'N�(7�p��Mc���..����'�Bhba��	�"歅������'j1 3˪h�A`DcК!����'S8��&��0���
�*LxQ�'S���]�����
ʬ�4"O�X#�[�@\YrE%�"J���F"O~+6����$z��K���x�"O����â&�hE�"J7
@͡�"OL]�@߿x쌠��@��`�8��0"O����%H�w�\� m�B�>���"OF�8�G	;J�[���(�T���"O�xD�("��ؓ&��
'����V"O��i"Q�1Ͱ��a�#a��ܘ�"Oȸ��G�h��<Pg�Xq|��Y"Oz��I�<}B��΂�uPHj�"O�9[C��K���U�K�),LL	�"O~@r�k��Gw� �f� j��qb"O�l��o�9�T:bI��$��u"O�����Ul�q�(�
d���3"O�3r�
�_�&����D�\���"O�T��ǁ,#Ҝ+��X䘔��"O�M��ϟ?.͊v+R�����"O��[d�+6���
��H�Faˇ"O�4"��ZW��� �(���p"O�X1p+Q z��8cG�S�HN�B�"O�8&�TQ��x5�?���z�"OZ�Z�,	.k��:a�&v|�ԃ�"O��a��W�0�h�H���>VH����"O�u��@I�v��9��ʟFX�"OD5�d�WϞ���� �.Pr"Ox��J�#�䥰��W><I�ԓ�"O��JÉ��O�H����i.F�5"O.XsIu	�i����;���@�"O��a�Ѳl����,Ө^p �&"O�p����jK@�b��͝;R]�"O�@Q�$W�TѴ��PW�ưk"O�4j�'N�@,�l����K^5�"On��Toԯ{6�0DlC��>qR�"O|���8�8z4,J�W��z"O@��(\��D�Kޭ9����"O��VDԢ �N�K��$ "ܴ�&"O�����e�(y iU:S�C"O�EbB�W����� 8:�87"O,���̝�d�����Yr���"O�m�F	��!�½y0FÒ��"�"ONe���=*<z��L�5��Re"O��"��Q# ��ۀD$�:��f"OXq��]1K@� �&"�2�0X"O�ab��7=����D��laq"O�������T�x�C�n]�*���E"O�"Ԃ	n�Ⱥ�_!�����"O� ʥz!�/��� W��,3R"OƁ�t�SV@�ZF�{��%�p"O�0�M��4,�(�C���i��"ORi
�b�a�@�������R"O:$)� I�q�D��'�IP�cD"O�p�nF2L�r܋��O"s�6��0"Ojp��NȾq��x3U�	�(�^��"O��A�J[�W�n�
� m�B��4O����99M�ّ޴��<qBe�-T����!��~��wI�0�]��
�(��T���W�@�qR�O�~H�򎃎��DF����F��"f*�
6���C�M�Ѓ~����7��6�F �O���Çgc��9M��!�@͇l���E�ǘp���h>8��䟸�O<Y���?��Opf�xu�yc�f��$�ވе�>���i f>tp�G"�9|o�00lR%]��ٴq��V�|R�O��T]�0J���b>8��p�Z�5��T�1;�R1�Szx���I�̘��2�[$<��T��@�Y�.=���	�,��V�\��@�vl��Z_�L�#/��:<�5��l���C�a�!���6��.]�,�$rdM�Ѹi�� ���x�'����+!�ʴOL=���DM�	��@2dש,!�&�'��ɀ!�NI�?�����*�p��C!�V�<�%.�+�y�3���ڳ�FW%�/һ�~R�s�h�mgy�i�![�*7m�O<��� P�̒;�8貳�޽Y�BL���O��#4	H��@�Ǚ����Ǆ��C�FӲ4,�(��a��U����1	�"T��FyR$2^Ȕ����e�v0�!M��cv�({�`��:�@4�pII�nS>i��BY8�$̠���ܓJf��ɩ�M�q����i.�I�3a�	1�1�tn΂Fl���b�O���G���}���̪vP��-�:��h���	�M�b�i����͜[̰;�mM�k�0L
Cf�$�~�'da�7��O��D�|�d�Q��?����Mc�B#s����1@? �%6=0�C����r���.gb����J%���S�Z���)�x��,���2�H$��mXA���A��6�.B=ơX�F]�4M�XQ�Z1��;�Õ
<���$�����ƌ١Q'�`���$̗�f���xt�i1�������M�<%?��Mcd�E	<R(;թ�-�n�����jܓ�hO�O�q{���'�9��]�?�R������A��4��O��u���N<��k��͸a.ɔ'DrLQ�d����tU`��ّX�� ����y�䑙nɞVYN����M#ׂt8�I��\��Y l�0����|��"�")����01E��@�	h�@+2��(�F�r�A86R ᭟��P�4!*�'�AB*<i��k��y�b��OV�I��'6�6�ޘ��ȟ���i}��Y"�x��G�M�^�9ەdS���O��~z�lT)F+�LHӬ�2�V��bnA�3x7�Tۦ'�4���?%�'<�� mU�	��i�t�Ùj-$��'[�TÌ��p�'l��'l�"��	���'kҷ&�)IAn��B6R��`za  �A�.{�v�8��S�	����Y~V=�d�*�f�x YE�`.���䋣?�z�)V��6qQpXPA��L���Vb֤��!�L(�f�9��d��+2���^9���E��t�HI	⌈����%�=�$�O��D?��|:���m~P��S��ʢw� j���h��H���#h['3��6-C��2��R�O�Em��M���'|�'\�J� ���   (  �  i  �   	,  �6  %A  �J  �U  $`  �j  t  �|  P�  Ƒ   �  ��  B�  ��  ȱ  
�  N�  ��  ��  �  U�  ��  ��   �  b�  ��  w�  % �
  � k �% �+ �2 9 _? �E vF  Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�� |d��"O
`�(�;���8���-0��1%"Oj4��ND^[��"3/9�0|H�"OB���H��*�ʞRy=a"O�味V�!X��!&F�:J�$���"O,��a
���C�Ą�M�"O,$3%o�-���p���+Ն�:1"O��ݢ1����`���y14]2��i�<�6��{_���c�H�`�fX�$Kn�<��A̼VI�xR[�)�Ć�pඤ�ȓA5��('nߡ4�� �)˩%� ���,��r�؊b#`T�eT09���ȓ!�b��g��}�8�F��-? �ȓ
K|m�ș�VṔ���2�%�ȓ"R�X�j�4JN�1�˘X�i����̹	_�jZ��1!g��zܶ��ȓgil,*�J�
j�Ne��i�J%b���f	�(U��:���G��$Y^م�~r�� S�%T"���k\�jx�ȓ|4�1�îJb��@ӵ�ݩn�V��/[`�"�v4�R�!ʎ<��M�ȓ`:��z�ؚh�J�Z��$HY:	��H��p�m�C1��!��B:��0��EnjZA V;9����J[
2���	��4'J�EA�IVW&��~�(aZ��ӹ�>� o�Y�|�ȓ�f�A�
Ο7�H��M�$�����mޠP����/���ANXo*�ȓTv�����{ ��-7�*h��I��sB�8�8���3����ȓNe*M�悡;������X�o��!�ȓ'lj�#F�m�+R&;�|��2)n�C��0S4���T:
b���:�0!��e֊��)��ͷV��,�ȓ0�&�8#���� ع�L�����;�P�AFd���,w�6d��r�EQ�( �gVlɦ�M,H��	&T�DCx�M� @���Z�!�Z�/�N5Fk	�9��gG� c�ў��Ӄr�b� ԮA�IV�/̡t�0C�ɃU߶l���ݵ3@*1i��fl"?���"P� �7�\E�h����!�d1�R��d�=#��y3�d�d���3�S�Obz�J�,T}���E�� 1�'�
e*T�*�� SF��5$h0�bI�`����VͬU��F Hu~�'�4"2L�?���)�
8�m��\�%l��CJ�X�X���]fId��0j��9D��C�ɓPۆ%�E�� d��p7�@�lB�ɦ<B��������`1hſ3����'ў"}���6�\ZwI��f�L0 ��H�<��j� [�(�q5��'L�S6��M��M8��0�ğ�,0RI:�AQC��d�*&��(O����'�Z�����X�� #8��ȓ=ʒ��Q	�T��H����}���l�J�����F��B�>`�O�!*|�F/ً�y�fC�e��3���	yG�.�y�dU��,h�� ���j� �8�0?I+O���#P +�J�;*��H���xRD$�OHC ��a<��S�A��6ư�a6"Ohm(���P�& �\�x�"OrIJ��+UH���T��\�� "O� ��N�3�($�l�;�ܪ��'�!��Ș&�n�i�OΤh��e0Ŏ�^�a{2���?��F��$L����4�!�Uv�a�F���u;^�RB,͗�qO47m%�S��E�8���-Nv�`'U [G�C�Iv�kR"oVp"foS�3w�C�	1�hk���(o��Qg'�?#^�G{J?�js�� .B@�MT�SL܁��4D�P��A�;���E��jL6x J&�IH��l��M+fRqB2��46�<T�5%D�d�&E�M��jCJ�'G~dꂅ5D��x4�ۥt�b�#��K&B%��4D���e�U��d|���kI��N/��0<!%N�1x�޼U��2G�$���M�c�<!��	P�fh����N|�1�L�����"�6���Q�	���J�eG"b)��UL�r�̏����6hf�B���<تc���$��挫��B�	 4P���:K�s�L��ms�B��&��t3E��94a�ԣ�
�;n��IC��)�O����'����F$U����=j�����nMF��6;\� l�Hf�ir�~ʉM�� [V��9������P���O�c���� Ȇl��H��)�R���/h��"O-BwG�~�Nh�JC� \�b�"O�٨DkY��d�[�H�

�,-��"O��B)N&\���<v�vH�S"O`�JqLĝ&���ȏ ����\��E{��ɒ�{�2���L�8IP�쀦��A�!�Y���3;nQ�b!5�!���f:��"��Z1*Ij`f��Wv!�9n˦	�=��E���{�!��DJ�na ������r0HʡU$!��?m��ij��-�(�C�I(k!�dĉKN^a�%���8$CeC�4`!��ܘrʺ�Xf�Z������ц*�!��I�^DX�W� �P��r#L5m�!�D	�P?~m!!�\5��P'b
�!��T0��Sc* 3����V�!�$,��Q�1䝖��l��?!� �H�Z�" ���0d�a��P�ԇ�	�T��L��BŠiY �	�	P	\�"��9ʓR������)9���;��ȖF���+�O����c�5r��ĀR�<k���@�O&���G�D!�q;�#�&.I�	�'Ү\AF�ThZ`���T0�q	�'X��[5���A��I�銀u~ձ�'����"��b��Z�yBhÉb�)��n�!.F&)ǡ �T�q �6�䓱hOq�T�4FQ$W����Y Z$pi�"O�K-ϣ%��QK0��%�$�"O�!kq�ٳyPT��uB�g���s�>A
�HE,����(R���S��;R�dt��	��q�=�j#I�̨"5�V�7�pU��Y�<IЪ�)~�Yh���,Ȳ��T�<�P��Z%������q|F�J��MU�<S����$���)7*t����G�<a�eZ�,:�����]gV�r�@�<Q!���|�U`�lU�qƪ�YG(�}�<�g��w�5���ƻf����"�t�<���ˀb�B%.��,���SW�ZE�<Q ���#��8�F@R�:�k�lM�<�Qo�$wt�e_L\-c�E�'4a�D�֕�4� �A
���p5�Ђ�y
� &������&�0�!�ƲA��+�'�%n�V�SFxo�2w@4�GJK����!G����>��Oi��;�L0�Nמf/��s"OxE�%�MζwdHy���I'��'%�-���u�ԣa� �Ip��1ͤC䉺} ����.X�*���)BR�C䉽��m��K")��@����ON�P*���s�xCB ~@ B���x��8U�*,O0�<�tJWsVԸ�ϝ�>k4��ӎ��<a
��[�np��`<Wc�ILH
����񉂱�,�p<��-N:V�tk�.F iU�)����M��y�DO��0t��"Q�.�*���N%��'ўb>I
��ՌL��a��^�.����e&�����'�p����$,Ң֪��!�ȓj\���돁 tt��R��$QL�L��3b@"����W������ȈB��An�t(<��DE�6�s�#�"|���ϊb����<��E�8e`$�b�O�r��[�@VW�<��J^V�i11��t�����Q��?��J~f꜓&w��2 �U��V9�JO�'Lў�'[3,�0�K]?"���
Q�DpP�$Dy"�'U���]���/Q�M�����1�y���,*�aR��7�h��*��yR@S&!ֲIڐ�
4��R�)�Or"�uc���,Ҷ�-(t&��q�k�<Y��l-V%���`U@�
Vjy���@��(������ݬ�r�1�бh�\��Z�����Swc*)bb*C�|��E'Q$3$ �O:���&%3�_0���kv[� ��%�̄���x�ЃQ�
`(��BAE���,D��hr���.e�$c�M�b��&+Oj�=��D[�|��e����9/T��aOO�<��
��&�P	��F,;KĔBPJVH�<G\ v�� �玥-&��c�]G�<�G��(�1n�%�P��A�<��Ƒ��4�bI%.��FE{�<��C0r������*jt���a�w�<�u@A)�x ��@��O�v�<y�b��6��i�E
JI�Y�DGZN�<Qc�M_�]��bO��)���Zn�<�v [�-�V�r�f�Z�zy�l�<DnBw�ޡqC�2�!ԂMS�<�`�E�� ��
��6A���G�<�T ����hVMS�u��B0�G�<���U�A�-�J��ԦFG�<���R��0�z�I]�x	��b�j{�<q�Բ6�*ӯ�"+^���c�<I�Zj��}IQI��ZN��t@�]�<���%{1z=@�S�������_�<�2�[��P�v��0��hI�#D�$�!�5!�v���A�6Cn�w�#D���u��!z�q�c��+>9{F�-D�����E�s#3g�=njޠ���)D�H[f�R)�A�e!�z���"�&D���dװh���c^C����:D��!#�T5�Yk&`�	g�����,D�(Ș;c&� �WgZ�>��y�Ԅ%D��KP̐1M ��@�?C��q��(D��!e�Z (���H��7@�T�w&D�Ph� M�Ԥ�g���V�H���'D����F�8Ҥ�`%��n_"$�2 $D���g�dd���K�4�*@�6D��	���&&�p��ȳ��)��5D���5�M�a����	�AR?D�� ι�#h�;DG�P�2>�S�"O��(#(RM
dp!O_�0�A�"ODu	�1h�fي�#����"OV���iH�!�F�1c��4�ը�"O\e@#lR8=��@p��x�5A��'���'+��'Y2�'�r�'�"�'�F��Ӌ�9�0�ɑ+!i�f�'�R�'V�'iB�'���'��'�����d��
Ҧ=�0�P&G7�,�q�'(��'�'x��'�B�'yr�' �Uke���{�&i&�I�p�\ِ��'�"�'8��'��'�2�'��'��]c4G�-���`ǁ�����Pe�'y�'h�'�2�'���'���'_�l�G�� v�F�@�)o��{�����	�����4��ԟ�	����I韸�� ƶ���o�s�޴ f�̟ �I㟐��՟D�����Iʟd�	ݟ�B� }w:�`PH�X[p	�ᢇП@�	ڟ|��ԟ���۟T��̟l��ǟ$9$�Hi_LQ��τ�a�:D:��E����Iڟ��	�x������	�l�����+1�ռh?flb�h�]øi
7O�����៴�����I��4�	؟@�������D5;�&�֯H1�ҔZ�)E䟨�I����	�X�������ߟ���某k"	�VK���Ūf.6IS�M����؟���џ8�Iܟ���ݟ$����	f��\$�R��vxD�O�П�������	������t�ɸ�M����?	�\F)�����ԓ >`���@�	ǟ������ć�{�إ�x+u !�<�B�뛷G���{o���'�ɧ��'�����)��-�B��2z���!���0Y�7-�O<�w ��3���,j[��	�&��iT�'y4B��v-�%K���3ՍI����<���;ڧR��P�!Ɖ.2��-'ԤCt�Y�i����yB���̦�h�(P��C'�l�K�Q�$��Y����MC�'��)�I�4Ǭ A�6O0�m�X�ɒ�!\�"vT	z6O  K�%-:Nʅ�cg5��|j�R�،��/�2��Q[7���~9���D=��Uه:��?�ܠBj�5Ҥ!�b�bx��?�W�T��ڦu͓��DC� x(U��ŵ;�Hh��o��ɍk�de�f�+�jb>1�A)�jl����x]��fVb2Ax�HW D ��'P�	��"~ΓnI�ɡҠ� ���!��Γ=\������æ��?�'
Q��uIS��p�'��\���?�޴�?Q�dO� P�i�'�Dx��e��\��'�saƠ�e��&;@���P^}�$!B�g�F��P��*s�8���a�C>z���0YY�F
U3.�P��ŪWȼ#�%�4N�q*�^2�\�v�&2
�¢E�X����R���sDD��a�$:q����O�h�Ц�BkB� b�@�R�@	t�$a@�Y���)�$ċ�G�N��rЄ�SO8��E�F��I��*Ybm�7�ʛ(Nd���ˍ7)�ċ��F�Bl(�gI����,��k�(�L��H��O�e��|8�H�<��}���Ijm�����ԯ�Z�EӍ5�tU��7��ӳ��HX�V�'�r�'F���O$¥�:yib���7��ʀ�Oxi�^�x�ɽK�x�?ͧ��	�nq@�!ŋӈ�Щ� �K-dn7���|n����	۟��S�?=�	㟔�IPc2Y�ƈ��U�n0�q���[7A�ܴX��Ax����|zK~J��S�v��a�VfT��peD暹�IQ���i�f�'�8��$�v����O>��O����*��S�\�>_���dZ�q����v�iq��'�`��TjQ�yʟ����O.�O�eC�Ҥ{�.UY�I]!Dm��l����� ���M[��?����?�cU?��I� ʀ�]S���R էj$tm��?�NU�2�s���	Ο|��ޟ8�I���I %FJl[�3V)��K;O���c��M���?9���?��^?=�'R�0�H�B��I��x%�;�@���O��d�Op�d�O���Oiؤ��Ȧ"1B�;������(�(���!�M���?����?1�����O�}:<�L�I�J[dM44)�*́Ie~�	C�F}�'(�'���'~��`�|�D�O��1e D�w�����ĺDv�a7ˉ����؟��	qy�'�kpR�0�bVb����'	�F���c���o��� ��蟤�	=��dyݴ�?Q���?���P���� hF�D�2��5,��}�нi_�d�	jT�S������@�s�n;p��|$�C���v ۀ�i��'pH���vӪ���O��D�����O�]p��*U�J��,|-@m�p�E}�'禈��'�ɧ��~�@&�?�|��Fƌ�R� ������@[�MC���?���j���?����?	�O��tB-�%H��5�X%��`�$B�'��i>	%?!�ɓmw2�Ȥ*]���҈�F�#�4�?���?� L��'�2�'=��u��R/y�����Ɯ�RLS$�G��M������h�?��	�@�	/y��x�ց
���)@�G¯{�|�B�4�?�3�T>y+���'B��'"n�~��'�Ҡk	�?"�XZd�� ܦQ��O�u��3O���O����O��|���x�pq�*St���U��$�I��i/�'�B�'4����O`e�E�̈́JL�I��ۮ-N�i���â7Y�I��@��ҟ���i�T�J��7��`��SAa�G�^���K(=lßH��ӟ��I�̗'O�&[7��$�޷$\�Dx��=�>͛�a�;��ꓨ?I���?)���?�1"�:����'�R�I+F�b�(����I���ӡh�P6��O6���O�˓�?I���|���?�슳h�dY��ɊZ�j��ٖj#P�H���?����?Y��ۏ����'���'����Ih��V�J5j�Q�e�4}�06-�O��?�p���|J���4��� Z �;��$��l�vj١c�i��'9�pa2�cӴ��Or������i�O���ऋ;e��x#G25"�p����}}�'x����'�U��[��V>�*!j�C�2�Bid!��=���A�8C�t6-�O
�d�OJ�I�@�d�O�����s`r5�V�^�}0<�cS�:�v�mڠB�����G�i>�'?	�I�&q@��,��[� s��	�FM����4�?���?@G�#Z���'$�'ArE�?=�#+U� �8ɋQ\�yGv�!�i}2�'Δ|��Jѕ�yʟ���O*����MkzQ�5C�/i��$�Ѥ$���mZ�ؘQ*z�ٴ�?)��?��L
��V?��U^�9�wo�t�d%�&�\}BǓ�y�'KB�'3�'���'�B	�fbT�`M�i+��E�c��A�B�M-i�@7��O��$�O
��h�TP�̧���z����^)#kQ�1���3Kr���	�\@��U�����ٟ$��"�@�۴Tob��b�J�.��5�5���ܤ��i�B�'���'3rU�t�	zQ��;��LcQ�S21
m� .�pf�i�4�?A��?���M��StF͠ش�?���m,(�cƄ�f7�$��@KR�@���i���'��U���I�4��ן��1�:�1 ��Z�3Ѥ��J~^yo�ԟ��	����2)|�3�4�?!��?���eH��2Qx� ��6�i��]�,�	/�$�S��8����4mV��҃�>Rl�i����q�o�����I-Hg��4�?���?��������ތɠ�ŋb��k�mˬu�:�Z�_���'ک�	ʟl�����~��P�p��k�¼Ƞɚ��e{diؗ�Mc���?����:���?q���?�Ud�h�~��)��Z9�]xH���B� ��sy���4���Ӽ#W��J�-܄YA��§��ev�l������r�K�0�MK���?���?��Ӻ{3�C�~h�5�����I5:ٸ҃ܦy��y��Ǳ�yʟ^���O���C�[�T�z4�K�gA��#�"Z~�Dm�蟀���ɯ�M���?Y���?y�_?�n%
9h�E�`=�h(�n�{�m��xrJ�(c�l�H�'��d�'P2�'�M��`@
�{��IA�B�K=$�i�`f�����O����O8��O��IןH�Er�ڼ�B��)w����o~��	[yr�'��'mb�'b��C��ʐ+&O��5���(Ƚ?`�r�#��1�Iៀ�	ǟ���|y�'�vx(�O��@*l�:b�<8����/+#DݱpOyӄ�dM�x-���O��d�Oj�04�Ӧ��I�� �$�m�2�㰂�;5F�Y9��M����?q�����O:EA�2�B���O�`V�˿zt�h�환#����Q�J���O�˓���ş��')���߂+5�-i�-�%C�D��O�(O�ʓzCj�Ex�����bDR^�F%�0\}��Q�i�	6�y��4%��韐������E<b�愂E���]��֋W�V\�8�%�-�S�'��T���V5�� �F�LmTlڻ(��޴�?����?�'FՉ'	2��"�,�XG��l�t�p7(��6-X�*��"|���rt���dmу-�mrH�J��i+��'yrôP!O����O�I) "�s�!L?V�m�!`ʝ��c�X�B@/�Iܟ8����0��V�$Y��&]�e�@��.��M;�M�0���x"�'�|Zc��ܠv�������I�0@āȭO|�0@���O2���O�˓]��E�L�AA�p�SK�;�D��	շ%ȉ'��'k�'�I�'٦42Df�r�y�%6��HA��?����?*O:<a�O�|� ��{��}�3��,P�բX}R�'��|B^���bˤ>1��SZ�!ȁ�>`�J�n�R}��'P��'���1Nl��O|�T��m_�܃d*Z{>�Hr�@�/,����'��'Y剆%�b���hJ/+k���4A95$�]���'��'r�ɡ3|��J|*���Z5�����k
%�
�a���bn�'K剱p�&"<�O:DL#�
Rl@��Ĕ�j�\��4��R��HYo����i�O2��Mu~"��D� t����S[аB�L�&�M�(O2�)���@�58uN�y�(���lJ;�B7��.=�0Dl���0�I���4�ē�?�M�'����E�-����G� f��F��O>��Ij��jL��ES�K�+��p#�4�?���?�ӣ�
g�'��'4�� �֜�g�K.S�b��� $>F�OH k���O ���OL��&N$-�<є��#1H�Z�/�������uhL<���?�I>�1iD���7��Q��: �C/X��H�'��p1�y2�'��'�ɒ#aj�2�� 2���]�TULY�caן��'V�|�V���!V)(���fŏ
L�e6�B�f:c��I՟��	jyRj��瓎&�̌#���n�>Q�E��&R�jO���>���<���r}�j�,,�6���I�@��$��'8��d�O����O��My<)!��4K�ihn��!��+:F�%�W�̌4l�7�Od�O�ʓR=��>�P�!�����m�w�Q��@�1�	򟨖'&����0��O4��!k�1X� K�}�ȹc��S�9'���'+�H��T?9ґZd��2̙�rȨ� ��}Ӱ�p�j�[p�i���?���aT�	+D��0����-�h�鶊�#%Ȝ7ͳ<qp��r���OQ:E���q*���G����!ߴ9d<�� �iB�'j��O��O���I)?���E��xyR���c��o�z��L�?�g̓�?��� ��k�S��06H� �b Y5�i�r�'��i�#c�c�x��П�B��ս8Z��te8d�4*"�L���'��5�y"�'�b�'��L
FaV���|`�_X��dq�*��4²��>����?�*Ok�8	��ș�Y�ngrX(�霉2p���c�4��П��	qy��)9��BrA#^`�8��N�C����o*��O��$:��=}���/}�>���� �3�@�	d؆��'}2�'�BZ�x���<���bքQt���#�ʌ5\īƧK"����Of�$:��?ʓ��G��X����q�8ı�'!R�'�2^��s�Ү��'hC�1�3OY_�:��1�_�B�� o���x&�4��	2I|�m8�O��J��X��#{:�6��OZ��<��'J��O�R�O\�M��A'-۰)�2�;Nf`	��*�D&�OY&aӅ�D�"dY:�I9F�i�剗=���z�4Gd��������8aX\u������8��6
O���\�>�
�AG��! PQ�idPDz��zӌ���O�����X'�,�	�K����04p���f�!��yA���?�r�� Q
�5��e�`O~\H���i����'��'�^h��A4�Iş���iN ����j��="�Y��E1lO����OP���*%�m $E*YGV�� $��En����W,�8��'42�|Zcz�XhC�E�� F�2�N�j����O��D�O��8�#i�pbm!�
�Pї���U��O��d1��%}""I���Q��1~* :�Bɥ��'���'BW�p�ׅ����aѺj�b�9��ޕ
A���U��D�O��(�d-ʓ��� R�G�nTj�+R��'�N��'2�'\bR�� �JK7�ħ>)�z�/�.b +E��lp�R�i|��'wj��.�|ؠ�h��`�4�?����C �X�&>�I`J�
	3 �tA0*� ^��J�a
J�	f8��i�E^�38�Y��<~<���pӺʓG�Nؙ�io�'�?���������֯��y������7�<73���ª�E[3h *�&�@�M�R��O����';��'��t7��O��#�*�X�A�`#͊0�<�bՋE؟��I$&(��h��ý3h�Qkek���}�����I�@�p�+H<���?�'�\��.���C`�F$~��ۓ�?���?!�E)���PN!0���z�m^;���'��X�
<�d�O�1���fdJ�N�^���X�g]
S���ʟ��I͟8�'|y�%��;�(!y��&�~\jB+J
W�DO����Ol�O��'�.�"I��0Pq
@�R��a�}��')��'��I�?*�Pz�O06(
��zHte��J@ؠ�O���O��<����?�5��[�$�e����K8|M�5".����OD���Oj˓g\��@���dmY5N���@���%�쭐�j�/��6��O��$�<����?���E��OeX�ꎞ0>�E���Cf\1x�i�2�'���6.�.('?���?mC�F��m��`!A�̚�)�`��I<I*O�ذG
/��~�4cց�Zl�6�/%c���ɦɖ'H��h��'�H�'�?a����ɋQ�JIc��/8`I��lE�7-�<鲪�5����Or���!����} #L�\�Z�p�4v���[Ŀi�'?��Os�Op�$�ty޹(�䟘6mL,��]�\w�anZ*xV��	H�)§�?���*	B !HK^��A1�bسr���'���'2.�
�A1��O�����\����V}�bǏ�W6�P���!���@�nb���	���	7`��`�H��+�0���k��I�4�?����c��'(2�'�ɧ5�N'y�Z�3���'$���a+���$5e�>�Ŀ<����?�����$Io���{7�-c��0��C���B�I���ǟP��H�ǟT��4H�ޜ؇㐢i
��a�(�+4l*!%�e�<�'��'k�X�蹦a����`ٮVRD�����*��C���d�O���2�D�O����.W
�$W�<Wh�yf�;얭jUKٻn���'��'�2U���G��ħZaVnܬ)�@}*k� �X�x�i�"T� ��۟��ɜ�D���Ay
Ob�#��Ul�Q�W��6�O*���<���
$|��OFR�O b�C�	��Qը%�bXh�&��)�$�O"�$�)�>�:�T?�ȁI�I��Z�כM`-�t�k�2˓>2T6�iǺ꧇?I�'��ɭjv" ٲ+�A�� @E�Q�6��Ot��	�*�*���|�'K~Y��,ז/�8�*J�&�A�4:�|ݚĵi�"�'i�Ok�O��$�E���k��E��Ja/أ}<)m�# qv��	v�)§�?)���/�.l
VI	�^�h@p�@�:.�f�'���'��Yը%��O������C�ˑ�U�pbZ�l�X m����'�H�:��|��'�b�'�A����$oM�8�e�J�(�FI9��~�^�$I+\�\]%���	ʟ�&���*'.X"�Ԫs�p�z�A��o���,LT�����$�O�d�O:ʓ!�� ��[��^(�b��G�� B�2�k�nW���'���'#�'���'���@��K�<�e��B�����E��m8�S�T�	ş���OyBA�l���ӧ#��2ށO��� ���O6�D�<���?���Q��Od,�a�X�T�P�Y �Y|��O����O�Ĵ<YT*�)F��Ou@���́n������O�&�4�krӜ�d6�d�O���)����"}"�N�J����d�0/i@	�nD9�M;���?.O,�)���e�՟�S�JI�y:7�����)R�	��	�V\�K<Y���?y�/�9�?�N>�O��D��3pu"�h�+���KT,�=xE
�j��� ��Ԓ���L�l����N,�I�C�I���A���3gDf�W�3=��"ȫ)�Ըy�`�:�p	2!��;`�{r�]��b��g�+^dN�ʰ�ޗe��q+ԫrլ�BgǮ��-�����*m�N!JL<�1�ٙy4��i�_BT�MS3�ĸe�@��!1F�i�"�/�h��v
Ϸ!����Tl*-�A	��q����b#?Y�dEAF�_�:��Ժ'��7�Y0`Z&^��r��D/���""H���'���'��]��	�j��)�B�@�0�z�`�,�>�B�	�%i����{�fҤKm�Xc��V���c��9���^ո�W��s�4h��R;���	� ���$�}؞��܅&��4�!�� � ��2�3D�T�"�[�XS�"�ل��HO>�:te��Mk��́(N� �1YN�mS���&�?��?�{��x:��?��O	Rݒ�4_�Q�DɎ4�I��ΐI"�[FE;Q+HhI3�<<O�|:E@E�fM�� ��
!�X�1���S�
��V�K�" �q�[��i��̅\����K�O�@l�iz�`!Q�3�\�`��p� C䉱'��:A��� DA֯ �B�ɱU:�0�p�F+
�P4
�ɼ�M�K>��^u��v�'�_>EhE-F�A���DnE4*��Dɢ�M;2+h���ݟ��I�$"S��r�2��h��DY��p�0�,G�t8��y�k :0��[R�	,��@��ʮd~m��G8Q��;%K���( �@��+!{P�0Ʌ� |*D�=���I���F��0���KReմb�t�1珲�y��B����*WBt�d�E*"=2<���ē�R��0�u�����:o�q�u�̀GX����@�d�2Z���'˂7$�t͋*����Zq�ַn���"qN�&o�"A���4!��7�|M~Γ%
��e��
gsV�w��T�8�[D�h�t1�5��G���0֊��oX�v�P V]�̟��ř2�^�Z�¨m\rD3���t�Z�)c�'�r$t��$8�矠�W�p�f5�����i
x�y�{�(������IWyR�'�b�'R�	�aנ�J[�e�����j�1�L"<�i�7��OnZ����S�?�"WAH����X�K?Obm��DF���;$�����h�I�������u�'�����C���'[P�⑬�0Kef���&b��ˆE!:�h����hO����GR0J !�Ʃ�M*.-B�E,��FBPi�PA6cQ�����>&���e�.��I!'�<�i�b�2|x�HK�?_���N���d�C؞���mX�24��%�Z��|'#:D��@vO\�n���Ň\:������HO>5��%A��M�!�H�h���,A=J�p!��!�?i��?Q�Y�X���?��OT���	(*�����R�̐sB��1���+1m��u��7�A �џ�aHɯJ�L`1*�#H����&�Gz��µK�1L2`�1���0oZ�y��7gނ#<���� �۴`�ht�gvP��n�2\4�$�i��O%D��'vl�+�g��t��n�-Xu��a	�'�.�A��AZ�\�ՏG7:�����'������K�QmZԟ��Ir��@\��ȭ�QG��[q�*"�Y�Vx��'�'�Y!R�'�1O�n�����־ctT���7j{�<�DL�OM^���E��_q<� q�˾n,���$ҟnI��5H� �� -B#]t�d���<C䉨&-�)��4����QB=����dp��w�vL#��'m���C% �H��Ʌ�� qڴ�?q���ɔ!I���D�ON�d�nJh���l^�IϋF�v,P# �O
c��g�'B�׊P D�2�J��v�ZYz%$��G��"~���w)�,�@�G)MRD0�7��)�HAע��8�L>E���>.��ks��Y�� �T��<L�B-�ȓi�J��e��(���Z N�P�Dx2�'��|���7�̍���"0�#w��*���?)��Ѻ �`X���?����?�g��@�4�j��e	"�$�3���6B�Pf�O�3�'���a0�KA���& 7$��u��'\���t�Y�� O�-,���Kn4���}�}�	�߰=�E�
TR¡�g�c?P@Q�a@W�<��-Q%N���Q�!l�2܈���$ ���Sg�I�Tٖ���4}v�(���$�����l�mJ���?����?)a �'�?9����d#��?�S�? ���FN*��lʖ�@
my>թc�'njU�/O��䗥%)�u�I�#k����'��-�/�����[!�웅��:6>�
t�V(�y�%4��Т����t
���y�oG%DB�3W�"�N|Pw@��y��k��Ox8�!�צ��	� �Og�h)ЇP:+��Y`�W�:|���Q) v��'�rLZ�r�T>�ɦ��f�X�@�B�*Y%��;��9�0�FyD�d(�6H������@�rT|�! �	��(O��)&�'��"}�`J_9�0H4o�1��`���f�<��B�0�P���T-nK��q��c���M<�U��.��U���E�H/�l{��<�U@]�0ޛ��'~�_>���柔�����k���vi~�� ��%Gz�A��=%Cb ��O�S�����u�bkJ�_�Y��[
J0��&6�S��?�N_Z��e�c(�e�y#�C ����������'D[��@�Ն�/��Q���y�A�*��������5r�nח�O(Ez�O�g�5���kG/��|���P�V*b�'1�]8 *Ǽf�'��'�~֝ڟ杛9�<�5W(9ݦ����U���	<Aۈ���:����G���p���	gj����}��*Ʉi�Q �6_���� "*lض>��'����D�O��w�j�i%٠<�Q�r-??����ȓD�� ��Lvj�J�V8�,m��I�?E��Fy"c�(3�6MF4ؑ��!�y�,Ӭ��J�x�D�O����Ob�P��O~���O�`Z j%������}N����ힽ�Ԑ��"� �p%�;^�8!َO-m��,0XO*�g!�*H��3g
.���NHe�����?I�e�� G$ W��IB�]�F�`�sG������I{yr�'��O�� xԢ*����p4�ćժO�@��+��k�N7�����*}��̓(�\��b�i��I|�&�I]wQb�'k�N�2��"��~iFpAa*�+-�b�C�`�	ϟ�� �� �<�O/�p��K�OXŨw(I/Io(IZ��dZ�K�?E���֎{����<	}�в�,ʓ./�T��d�O����s._TۆfNJ��:
�'�ܐ�6(��&���kf�MI\F(�	�T��'��aC^�-��Qa��V�C�ղ�'��h��~�~���O`�'zf�����?�8��c�߆%� �SK]0�ΐ����B4�QS��� � �B�h��R�����#ܖl	��zg��F3̤*�.A�nH�X��ԳgBag�@7V���q��Q�|mZ=4d�r\���㝨c(٠����7b� �e��	z1�ͦ��*O����OJ�B�)����q A�E�i�8O>��,�O�\�&/�YV�(V^6-?DX�e'�1O�!nZ��M�H>��'��������J�$��2����%՝�?	��HS:���Ҏ�?Q���?	�>���O@��?5 ��v�иW�9����\X�d�M��}�̈́4e�q��6]X;�`V��~�����>��� k՘a�T�H8<<�w�_P?����d�!f�)sc�^�t4�F�V�VB�I�>�V����3,�:P��C�:'�h��4�ГO�)�7�ߦ�@r�C���q<ԢФ�{'"�'��'�X퐷�'��'p�P3c,نYRZ6-M��t���¦P�����!L-L��|r؞ ��e��%�12��1LZ�~^����s3$�e��vRX���ɺN��Ѡ��D�!��|2�)HV����<�M;�����O���'V����b��#	1��hT�P�u������?�pL>FX��p��V�a����*R�<i�i��6m�<A�a�4@���'�RZ>-�G� 7��^"G�����!��1�Iß���<2GFt��#C �1h��<�Of�	��kS�{� 
��;fu�\������+l����]�M�`s�Gg���*��y(���i6~	iC,ŪY%Q���Ub�OFpl�2�M�����CN,aV�w�՛�k&	"~�d'�)��<���S��v�B�.Ų8Z��E{���I<Y��֬�|Tsf)F�W�½�v���<����.e��*���?�.�X|���O��d�O��C)LS`����K���!˃/�
� �|FxRKU�eH�)Y��X���T���5I���;��)�矌��$	�B����d�
C�@!
��ͨ9N�0�I6��S��?�2d	�tڝ�4�]��� Q�T�<�h̫���j�lȳ3�Hl���P�'�"=ͧ�?1s)ԽINtx2��uٺ��E
]�?Q��N��rA���?a���?i�y���O�.˻3�x�z��+;�~xa�j�A:(j NY&�n��
&� y�џ�4�ʘ�� �I�u�O=&P�(�T�H�Xv���`�l�\k���8O�T7�E2_!�I�;�+�bL$��$�B
���-,}n����\#_k���m�.<lO�lBw�
8lŔpp3f	gA��+�"O
�(�#ҵm��`2��D�$�p�C�q����|�d9.�r6MN�;x$���ͶP3xhiB"�;,��D�O����O�C��O��Dg>u�$]=s	,L��X
 �QgN�N�` R�`�F���ᦢ�B��`Dr����q�!����+���wL�m[����PJr�1d~�x�i��8Q%���'�t�����v�_��ţG[�U��uPP�A��y�f�1�\ xR
¤OT��g�ݺ�yr�D?]����e�BsL�P��JL?�y�`dӎ�O�)�L�Ȧ�I��ؗOMXѱŪ���h�ʿxk-*��¢Y���'����5�lp�6�9&x�i�nG�B��j���󣌯AuHL8���Ox�Ey�d�Y�*�	��D4zu�̸!� $i���i�����A�w+��(5��C��<)!Iğ��شE�F�'�哧L�l�^�j8ܡ��KŷF���A�S��y���9��S�p�	Y�I��0>�G�x��ˁK��A�S��x����y�a��p$�m1%�'q�_>@j����I��@+��#'�XS�FR%ʀ(tj�?/ۺ�:�d.N��@��Hr�T�[���c>�<S ʈ!Xh�a�A&!z��a��ۭdl�Q�H����s�e�!�	��4�"*Iu��w���+%k��e�� ���:8$���O��R��)1���OZ�2`U�@P��C+׿���s"OΡ�4�ZT�S��ER�����ቫ�HO���Od��Ƞ��k�E�$�a�O���B���#��Op��O �DEú+�Ӽ�bg�\*���O�-ШdH�}Br䑐��z��Q;�ҟ�"=)�g�;s�z�ꃦ�$�
5"2�]�Z"l:DHJ5>h�];�+�,���'�Mˀ&��3�Je[A^���ǀM |����3I��2뷟�3���O\L��I=��̓�b�=B�T�����t6C����]�I�f	�o��9�P�{��4���Of�+�@̦��	,x��ò�2`��ɋUF����`��<�N���㟨ΧC�v���Oٵ}Ꚉ��b*�[ѯ�V�l*dl4�Op���A͢a; c˧Qd�1 ���[?`��"�>_X�FfU�p<�!D�ʟP��p�qC�Y6VdB�A%����+D� *���2��u���9���dE)D��x�,�>�T̡g#��#�곦e���4��G:X�ixb�'��S-|e�R���&R2r�����n�����	��X��LL�L�<�OB�Q���
�"u��B�&(��Q��
#&�?�1��o< qQ��R�fzh��*7��r��Ic�O��؈�/h,Fճ�	��_�M��' ,�*��|0���^�(���Vy��M<���W�g�~�+�M�)z��c����<��F��_ܛF�'��V>ER�C�ן��	֟�{P�ӝ[�✪��J�Y0~̈d憻.j�I�5,J�i�8#����8��L����n��a�tk��@\��C�6%��tN�*23��z�I1i��¡O�H�ϿS�'ѓ[1�ɳ  W�E��p�d_E{=����?ٖP��)6��X`�K��~a� y#�Cf]pT؅(m���	T��hO���ʣk�Y�O�ax��4��M��iQ��)�)<R8���n�"'
��y�:���O�ũ�d*u����O��D�O>�;�?��2�~ui&��7'I�p�H�Z�K1(�f\��J��K�=��ƅxr��$
.Be�u�g��  ���I�5W�8dSG��8O�T� т�U���ޟ"7�^�9�����ؖ�E(H*hXx��`�t좝�I,I*=�I��Ms����,O�ļ<�'Mr��k����cD5#��v�<�Q.�={�5�E!�L���Nf������� �'��b��|���ӡ�#o��4A"DE�@��T���O4�D�Ot���5(��O�#w�q+���-[6!D�� 0����`�'Xeb��9v���z��R�'�@�A�Iܢ@����qM޹j�T+w�	?��<��V�%�<C�@�ru�&fZ>����{B-
�?٠�i������SO�B�ʖ	&6u
(Z�'��С�a��i61)6�	&$wP�#�'��D�1���� �֯��ia0��'��7m5�D�(<L�oZ����M��*X, \j��vmKU]|԰�hQ8)r�'���'��<AR�29����FEp�l��)�~�t�Z�{\p}���J�N�ވ"��H�'��=�w-WL:0e9CG$h�#1��̑�&��G�J1�pOӒ`�~�I�(�S�8�w��n���h��|a��2Q��g# �&���"Oz[�T�Y�����6/�i ��'�O�PRwg��D��Ļc��^���B>O�SA��������O�p �t�'���'�x1�GL;g��(�.A:ܼأm�L��	r(�*������Aڜ�'��Ͽ�$�c��T���Y#��)T�K%"�/@--�D8���f𞱸��h5zc�
$���� F���޹WgZ�+P��
QR���j�.z���>�)�矐#�ʀ-�
����c^����2D��� ��*������3�����,.��t�b��A�
��� 
'�p�Ċ՟@�	�X��83���\���������u��y7�ئ��&R�X&�	�� ��NJճS�J�W"=����8X~X��O%����#�]n"��T/T�ܹ:C	�Rqp \���zEj۶������#r��4g�P�'�$2D�B�mT���0Ŕ'c����I�}�Iu��t!��a�V<kV�WeeԜ�Q�2D�ؠ����0TF81`�0z��7oR��HO��-�$� �XTm�+۪�+Ro�
�B��焥jgƹ����t�	ޟ���\�p�I�|��a���-��o�xC�@Q�g���l�_W�5��K��%�����KJ|�`'b��t�b�յ!Zd!H�+��L��0!&�L�9˚��xӔis��_�qO��S��'��6���#Ġ����PdFI�+H?!��.s�X�(�����̒:>!�_�)��q����M50�{��ۂ-�$�Ȧ�&� ;!B� �M#���?�,����&ٿ"��A����?u�X�C�3pm����O��$LiW�=sԄU�2�"ų�J@�?�O�8�XB@؀x�� �5�jc��D*�8Y��Ԉ\�(�����/���]�7-p��P��	b��CՁ֨Q�,"��?w��1��O�}�g�	)9�>M�'k�v�i��QK�<�ed��s���?=�Ve��AVF�I<I''Ĩx�p�5�	�5P��!�<�R�ϵ\���'��[>}��؟��I�p�O��IaC��p����j�l�<�����'��j�O1�d1b���b>��ײt�(�C�#��)
M��D3x1�c��%ڠ1CM��V�M:'�W�Cv�D;oh����o*jl^����98� }#�	?�谢��''1O?�Ą|�.(x�
M+�݋�(^!�D°T�z��UDh�@ �H�@��r��4�&���z�H9�b/G�gH��XQG�)*���O���bB�8jpf���O����O���;�?�;n�0��Fӝ@�7�0�ʱ���^�)Y�m���M��Y��,CZ��ѣHrЂ�S�9M0�c�g�m9����"G�/����a�9_O<�џ�7M_�m�bƓ�X�T���MV�	���1��� ���p����O���T�7ޚ���Ae)ڍ��Ɛ5�!�� )�"����:Kltq�e^L��Gz�O�'���B`��p�Eh20^��h�
��R������O����O ��_ ���d�Oh�S7e�2�p�/��M�2c��G�J�&T�X�0�B3O�69��4��n�'K��_�]XքN�G�*��W�6~޽���G�c�|�	W��Hu�Ԓ��ǣu��'P��Ы�<10ִ�5mL�-���'�����7N���DI�4�����'��	��73b�Ă��	�V�ٞ'�~b�LBF�3�MK��?1(���b0���&7� �đP�W�=�,�I柈�I�*������N		������-�J����؊d)U�D�yrD�d6�3f�ɨT�T��g�؆TK�qq��SWY�;�"�;oYe�L��J�7�4���Y�)�r��=��,�՟�J����6>���1&lT� ����� >e�!�d<�P=TGW�{SЁ�ơ�i�a|r�#�$Y3w](�#TE˥oQr���Y.��DV�G�Xn�쟴�If�d�*�B�'�£ƪi"(=@�̈́�lؘ "�h̚W,��e�B����	Ż �(Vdsڎ��;*0���TC]�R�Ԅuі��*�;7ѫQ(ҩkk Yyd��F�Ā�]��0��&X���w�&���+��:�tp4�希�����o�Bj'���O� ٓ� /f��0REW1]4���"O 8��e��\PJe��$m�(b����OL�Ez�O�( �x�)`�G�a�	˧fȯ	�b�'�|�ׇI~kR�'{��'�
�؟�.9'���A� ��e��EU�,m}�`d��VAh�ꓽj�ᙁ�?�Y���c�1OZ]e�׫.j82�W_d��7	Y�`¬�b��+!�2xp���!C��	�����y��Uߦ�X�ɲ̙�G;�~B��:�?	v�'�f�Jl��/��sF�K�^li�'K�,x�eЉ^Ot��=4�)G�5��|�J>ɥ"�8)P�f��9�ԋ�`� A��(qT܎s��'1r�'R��'�5�L��'�*a�&��kC�u�Xp2�/�b=��P�#�k���$OH?9��(�D�(O��@�%��{�. z&� �LB��X�.��U�D�Z�Q;k��t{_l��dŪuK�Fy�Y!�?�Ƕi���5읊o�<P��o�,=���c�'�V�zUA=q/(5��H����'@N�[$H�	0ͱqמm �T��'}�6!��]7�Ȑm�����I^��%נo#:,�ŬS���`��jMx���ц�'���'�Xh�D�')1O�SP����&A04:b�r��<�+LQ�O�V�;у�6nz�Y7�����#��$�:���3� 0��Ձ�44f S�rW�e��"O�<x�"��%/�)p�`��zBιJ�'|�On���8{��%r�m,?(\[�9O���⦅�Iß��O����'r�')�)P7��\DЉ	E��=	���VCg�Qˤ�z��Eђ��%X:맢�Ͽ�OM'W��B����?�p�R�1�
�S&h��CY�c���
�Q@�����3�b
�yq���6N�}a� A�<C(��W�)�矄Ч^�ny1BU`,���g>D�t.\��p�?LL��4+�W""<� �i>q���  	p����5�Pa�b��3���П�h�A��c������Iɟ�Zw��w�Zycq� �,<r���"�ՈEhX�Qqs�]�G�>4y������I%XR�Q�#CW4?�F��#I�Z}���&�W�3t}ۃ��QHBP���?��RVE����eV+� �-�*xL\��,�Z��I���%���I����'&6�!!��ap��6�Ȝ!�(��'tl9����U,|lA'i۲y�����()��|����E���nZO����,|�qqoA%$������@��ܟ�	D��ß0�	�|J��L�@΅�'(�}�`MA��=y���d��(�cҀcZXX���[6|�<8��J]$bMz�G��d������h5 �X%�`�by�5�$�(�Uau"��O&��'��7-�7u�4�'�
"�=[���S !�$G6ND��!������NS�x�!�dX�MoJ�)�o@�;t@����9��D��	$��V�ɰ�MC���?Q/��\��c�km�l��ŉ7���a��7W:����O\��^�Q��y����{%R�H.�}.ݭ`T8�"P���i�D�r1�S5�Ω��I�1�BSj�y��L�"�,�"=r�M�5����a�:���%�x� ��7�6��'������a��>U!f׏T��y@�]�D4���9D��gbX�>�Ri[!%��N^�D�!�7�O
�%�P��n�~��`)����!�h9���b�Hq�F�M��?q,�hѨ���O���O�QB��%H7�TSS��/`�\t*�۱���eG�)��J�M�.�Ԓ��dK#H��@B��P^0�#�����F�����B u��k#�:"H^xAr�ɯ #��߽ �����D�*;0 ��� Q����Ȳش�?)���'�@E�v�\�P�\�kԨ�z�'b�|2�'����q�),�<	*&dS;��a�P���O��o�M�N>ͧ�*�g@�+��!5EՑAyD�C����?�4PfQ0�[��?����?��Mx�N�Op���> ��0�ξ�p���[\=B����C-�H��Z 1Ŭ\�fן¤k1aߟט'b�H�O�j�8A�ҥ�%�| �H�t�0Ʌ�^32��Z�Ƃ����CD.n�D��<UN�]v�q$�H��h�%�U?����lS�B��0kR��'���B�cN�26�p��pB�ŻIM<l��;S�D���i>�&��z5@��M#��R*9.Hy�*K�O�F+B����?���?y��\��q��?�O�������?��?�B��m��@�a��U8����<ٓ�Q�$�`�c�P�����bIP8��Ҧ��O�$�+�ɻ��6x�2�MZ=!�dɴf�P$Aw��,Y&t%c'oN�~�!�$A1N�\a�gʑ�P��g��w��$�i�J�@mCbZ���Ih��.A�;>�1קC�t^��C��j�޼��'m��'��]��@7-~�Y�@'E>ԥ��OW�$M�?rx��F@�@�\��f�m�'*�}#���m2L�`��'�������|����k�F9�)4gV��V@�u���͞M�|镒�?���i�b?���j��JN���I*`o�\ �f����9j��l��k�Q���x��ـ	m�hO��|�I;G�x٠�f�$�n����I��	'=|Aڴ�?y���	6<�d�$�O��܄re�@qt��d�^����$ �}!t�@W�ڤH��ٶ��T>U�|�ɟV��µ�R�`Yj1�g��v���	G'�n{�5!��;J�
�ԨSdv~�V��w��		�d�vk�R��4'��<���ېp�R�o�F�o��4F���"]�P��M\M�t)"Q���k�ϓ�?��eJ�I9bHI�����JBp�EFx��1���i�P=�t��	�	� ݛ�D�	�����O�H���9H��$�OT�D�O4ٯ��?��<�r�ze�8	<���f�8���W����ô|58��'��b�	V =(f�05@ ˄��l�=\�
R�eKj&@H�����4<ʓq�^Ez��]�n�6M�3AH�BR1+��1��%���N�&,�a�,O~�D�<�V��`�Iҷ�4)�*��Wg�r~��)§��4:r��4���r���%tR�Q �i�`7�-��|�/ÓS&���8D+*K�YKt��=%I�U�S�L̟d��矘�I�]z����ğ�ϧ&5��b@�S�l��e.ī{� ���ϚZ�W�'a|"�Ѭ8��qӍ������&��ܠÃ�:n����Ѡ. �k3���@#=�G
Ο ��4R7(qSdg 58��px��83�L��S�? �d�S�.�x��k�h��"O�Ib%lQ5`Z���b��Ld���5O�l�Y��K���Y�4�?���i�&P�U{��ݯ=�}�P�X%xc�q �O��D�O�a�da�O�c�ʧ0�A+ C\��G���U��eEy�-���HQ���(~��J��ָ9~:8à�	�J��D�ߦ�ݴ�?I(��\re$�	t�D��I�:in|��� �Of�"~ΓJi{���d
�*�I�3�ޠ���� �����է9'�q�g A�[��Γ�h�b�i�r�'p�.w02��	͟�����u%�Q�4��(	��%"0iP��VΟ��<��O�)B&�E�d��)'[��,!6(]�S>�"<E���K���@�0B<���G������1�?iב|���'=���U-Hb\ҙ������H���y�ؙW�*���FG�2(��%Ѡ�OB�Ezʟ8t{���1����N�@�X`c�	�O���K�M�x��s��O,���O���κ3�Ӽ[m��m ���e��>g�}S�H�j?9�A�vx�Ԡ�iU���`���S�|8�������7�O�9��n�1��x���Ǆ1<H�А�O���4�'��{r�87���)�GL���0��yBl�4Z�:y�Q�Ǹ[��h!��'i;�#=E���L�T6�K��c��p����������'���'"`��\TR�'_�)޳%fR�'�L �Ɠ�*���%�����[��ĕ'K+��-u
���瓌 �dӑ)<�O���'�r&�*���J�$�{� �Q�f	�y"�$����ΐ�%J��w.M�y���W�dHGe�!"����ȇ��yҠ5����]`ݴ�?����)�H�"�A�B[2 y�M >�ZYz�M�O���O$�ʣ.�O6b�ʧGx�����ѦDQ�*PBU�#"f\GyR�ˮ��:t�&��;[��}�'�5d���3��	9A�2�D�{�O<���b�K?V3�V&�q-�<��'�vH�G2����g�<e���'x|m���-�4���)6�蘚'٤q�cjs�h���O�ʧ!S�����?���Y��8p�ޤoJ肱	K�RR�%k�12�
����(�rYV���%��O���
��]
R��%2:T���B^�-=f�IcS�0���+��ȵB.1�"�J�(tc>��� ̀Hzg˒"D#��b-�q$ �)�O�b�"~����Jrt`W�K�%c��V�<KTB䉑(��PJ���x��-��bS�
 �#<Ѡ�i>�	g�:aSg�x6�1��b�%����x`�� "g����ҟ���ß�9Xw��w3u���
3f�J����=՘ 9�'F���_B���B)v�(�{Eo 1Y��#y�!���?yY^`9	ƛ(���kÎ�'���	�J0��d"|O��f�E���`kq,�?p<�b""O�(�wjМd�N�0+O&{�ƥA�DS}������s��¦@�B;DZ�5넌O 4z��;e���I��D��7�b,�IꟄϧD�����qU��S�d�0��q�p���$�OHu�R��$�	?}x00Q
�	_p�X��,�O"l���']�ʇB��+s��M��������y�bD�0k�u�a��!F�����Ą�y���E���+D�\�.�#s.�yb�$�	�5b�!ٴ�?������-k߾DA��ީOp*u��MF�I���O���O� �'��O�b�ʧ/z�@�%ЁE�x�.J�SW�XEy!����n��s쌬dn�c2�N]3�YT�I4B�f���l�O��+r�N�$bp	a�P�d��e��'�ν��E7[�9A𨉺f-�8��'�Nx*�/�5lԤ	�
DQ���1�'���Sgm�D�d�O��'H�,���?��P 4U#� 
�m�t�Q��(S3�)�u�^.p
z@��O�)&r�ǅ��hL��v��ߍȄSV�^��+'Ug|�Г��o��`%�A/�z���S�
{�	����wg����'��}�l���eӄ,?�lKt�ɹ/~"�6���O�5�%j���pl�OV�9�w"O�9�ъ�W�FHI��"YH�3��	 �HO��@5B�@�:�v��g J+�0��	�rc�_����	ߟ���埴�_w��wvAK��Q�Z*��J��N�k,:X�'ȴds��Y��hj2�,O�9r0���s�Z�7��632�"��O� ꔄܣqij0�GZa8�l�thZ�C��Y ���K�LˢM�� �wM�O��ɬ�TH��oѱ+�DU6�L�Mn
B�)� ��3ӊ"�����Aa$X��F@�����PVH���9x���ۚy�F@
���:g��ß��Ο�I����hͧ)�V��I��H���T�B�����tiPHQ"�O^ bS�����6*%�Aɗ�����e� �OT�S�'�~6͈�]8�]�$��n�b��f )�!�$[���Iv*�+��KfD�'�!��C�j��n�!Nq В��I>�Ɉ��?A��L#���+r�O�+����b�<y6�A�?��p���?���rÍY�<9� �i���g`���pc�-�Y�<	q���
�����=aa��C���R�<�kSX���KǙw|\h�&⎵�y�cё T�d��m��\c�&��y�>4\���lK�0)Z�{R ���yrB]D:&D����q#�Q�aHE��y΁:J�a{$B6 ���+ �ה�y'�2xo��#�7��l��)'�y#� OfP3�C�T%��h�n��yr$�#l����C�H�ѥ�>�y"ɶjL�T�p��Q�� H��)�y-\S�����]�$N�r�(��y�!���$S�`�+��#��yB�A�P.Na�c�2O����K'�y��|^43�MA�J�S&M��yR�ݸ˪P��NZ�1��I��U��y�B� r^�s���%
��cvM�a�<	r���T�d%@Z:�*ċ�A�<�R��j b�C�ο!��V�"8�!�±]���ۗ��*�H���I�!��M; ���+q���<�6e�M�df!��)B��2RE��4�r�b�>5K!�Ĝ5/vr��9��h"�A
1!�%W���Q��Ou �����9!�Kn���D�"ah��Z&�� !�DA�'�TQ%�\D�����.:g!�����KG5
9�ф���M2!�$�=Yf�"�/�Q�U�R�2s!�Dײc-
h�E^:��N��6`!�Dɦ.Ŵ����E6^�Ҵ �˔�FZ��+WYx�I�
�hS��[Q�Oh$�YV � ����Z�GoL� �NB�%��Pł��<�$x��h��$�c4%�r��A�B�� �̜KZ��5NC"l�h��#�O��ͻ����}BLω[#��-ɩ$Tx�hPI.D���1*ްaX��HF���Fd��F���ט
LИ���G�A�@rv)��<���ll�(���ON.�'X�h�\P0ҡHC*w�nH�áJa؄i����X1Х@S
7pnI�ǩZ2!X��L�]�(�BŬzzrh�����'��=q��4�a�w�R)i
��+�ڴ,�^�@W�ٕr����'U�dc���bM���.�Ex������h~D��K�)��5J6EںW�������Ű�u�+� �zM���A�iRּ�'��<��1!�풀Dψeq��PC�#j����*�)ڧ%�yzT΍�e���[�Э*i��Y2F��e�	[��ɜ5ܨ�nٽ�HO�����`���9�EXw��<j���'�*͉��T?���M�<��fZ�`�0��C.(��)����	6m\R$C&�yW����2`֍la����$ևθ'���Y�C�^D��蘵A3ne	�O��K�2���䇷2� ��� �`5�Fm�<��#hրԺSD�u�"(�奜M��?�I�'�};�� $ ��?Q�t�@�|��7�9?�d'��d��]Gx��ܿh���&}�<2M^�=E0�3�g�0&�6Xb�o�Q�Tۏ��iFj��(�&�ݘ:�p��W�J��f$�F��(ʬ�G�>���+�f6��?��g�q�	�����)z���4!���J�r�En�(�앐�����*��)Z��"+A^Gy��Y������js�(X������(�\(�쏬\���p�=�	7 �0#<ͧ#ortۆ腉$�ڨI#$j��ђ���h\�I:a� P� ��L��D���T�>���	�!���A��FL���g�ua�Dx�&|ݹ"��"04`�O�;w��(��EaF�;g%Zаf��)�Ȍ0�N4&�
�Ex��)�]j�C�h�J�a�f�<+I��kу�pipEA	}�M�c-Yj���_c��{�O�e N�$$I�X񲐋N���w��%aɉ�� < Y���K�ti!ƞ�b�m8T��Uz̢<��Bth#Ύ�"���bp��I)Y� �r4@�8;�І��<D$��@4"p��Ē.���)7P2��d���u��\�i ��h��d�C�H�GǱ]4*�ˁ�ԏ.����TO�x���U	O.l'�I�&��y�G��r]RZ�	�|^�k�D�|?������J_��O$>���D.2��� >�	"�!��g�r�CB�i�)��-�aԨ�`d.~� ��@�"��h8�\�O��AV���3Q�ϗ�@� ��H8$U�P����7����VX��X�H|��B�$ϼ�yt(^�����_���$�/�eP���.�Ir&�I�4u񖟜��D�h��݃L*v�B��5�韰<`$�
T,!�!V�tP���%�c�h���^w�%[e��D�"�薖>Q'*��Jz4p�'��*tQ�a�
5"ri��O�A���=�g�^P2SFΒ��Dk�/G��D����s��-[4�\�xr%��C4�Ӽ��Nl��k�:�x8KPM�89�
A�O��r��*�)��y�(a�
NF��Ȧ�!t��Й���2V)�P�`,�,Z�@�f��u������xSY#:JP�q.'�.]����=A�П����M��a���p���爱xb&�T���'��a��\u(0I��(2q�.�0�{��042��>�5
@NA�1�<��Y��KV(;������40��;~j�4DF1}��ZIJU(�%�|G�I7�D z�
 ���D�B�ʋ{��qO�`��'X,0BT@�+��N%@�`A��
��Ā+T%D=����
(֨O�ׇv�
u��b˩�$L2��(r���fH����t���n�.���6�x����%B�Ũ��2�no�`�c��? �-�$V�,�B��N�42�E�'I�؉6k4�I2g����'�$L)䌋��iD�Pdʣ������HVJ��ѹ�c"?)�ǁ�F�L�w�פ�� tK�A�'�%���O( �[a� 50@�K�`7��j� �f�J�D�VUX�5���J��b#e�x��X�N,8U��Ӳ�
v�&�ӈO�`�����O�:�� m�8l�ڬ"D�=S��9�`�9ORƉ�"��:a��1���w]�Q$a��C��S,�6�
�'� ���i�pع��oK
`�\Qe O>�	��=[Rф�����0@g9B��u`Tq���0CQ��'�ԀS1̙.
��+4�91�\2Ƥ +�����jR�>�"<$�AG�ń*��Ez$N��F�b�I�<Y�O2��d	JВD�`N��K�̰��O��_��Y�e�[V,@�FJ�H��$��Z`a�,,ƕr%,J4p�~�q5-���6���jL	B�E+O#?�q%�#o��Yu��:B����0X�"9����Lm�7),�p<��L�D�;�D�@��iF�J�����f��zR�>Is��+h��9$���U�b`¨�p<!'�#�8�OJ��t(Gz��8)V�G05��I���I����с��z�Q�b�`��dX��R
h�'@ڔ˴F�E�S�(�yv�]�@ߪ��ů��d���'l��R��M�S�O��a�6'X2�*����FZ��q����
t�d�~&��E���A�!���zc��x�D<�)Mt����R� �j�a^���EPjW*b�f��4@�V��������ː��*Kir�I��G,�n�Q`�̰<	�(����']�� ��c�Tu˄I�s$	��D 8��a��D��jm�I0 "��zI`@�/I���eu����o�����J� ��J/O����{TE�`T�ye~��EF0V��\̓*���6YAX��w��>Q�6"לr?�A&��H�
�R��V�֏^�i��+ŬT0���$ՙ/j��)OR"?yЁW�P��Q�b�7����w�¯G�x�a�A?E,��s�9�p<�1�|!���2*��!YT�Ϙv�\p����=�O�z`'��}�x�Kbl��'=څ���9O���&��)��j"W�'���2u
]�� A',x��Ҁ�q�'>�	�D���C�F�� �(;O�|:����{����r�Z�@D�Awh��1�N�\��e�Б�?!�P�w��aV��	v��)���T�#��$�&�T��h`�I"��'�Lx�韘h���V�tM�!:�.ӤW���B��!U����7M$}����b#�K����!^�r�L�[:~(2���T�*���4�!zE�
�R�`Va�=F��Q"O���a�惥r�5:wc1Z`���	*F�>Y(ӈM�3����[��ػ�� #BP���EM)�Z�[��.�	�u�㞨+�Oh�ٹ��֪��$q�L�PŲI�ǯԗ=��
!�d��O�o�zmY�KŲ$�Θ�=�Ө=���Pg��-`²�Έ��؏{Roԣ?����Z��퓷��ض�'~P��sJ��� 1��=L�@��8z'�}#u  Ѹ���}�̆f���k�I��&I�eLl9b�$�k;�P��b�!��E}�w��9GE�m(xk4�[�Gg�P�H�P��`BW�S��u����p��0��	�7W�@YZ#�.�+ؐ9�b�0}q1 ����� �9���\�v<Z��ìS`��I��d�	pA��x��O)Iq"��3ڎA��hFI�(�`FoN�O���lPP�ńμ2<�SuN�S��=�S�z#M�5���6̓��Q�`�쵨�{ҠDv�nԂI7���0kƦ92��']��뒝c��|�ãڊ?��%��m��>9.�;�۷�yB�Vh��ԟ�)��O�)jbjIj�
��b���I���=zz���"���,��)�L�$jX�>�;\�T	COQ
��c�H���(�M���7͐�?,��	�H����@;�	S��
V�l3W-�"5й	��ɰp�L��c��3U�Ɏ*��
�o�#(~��[B+6�FX�m��p��=��C����Ě@��"���&#aB�x�#i�^���g@/x܃U��yUB�A�T��ut}"E̻2�x˦��p ��	,X���,�'P�ȑ�V��6�3��p}�&�>����U����
mB���� � 19 f��=u����.D[?I��c$�a@��VaZ�}�dIf�H ���+msRL�2M}B
��^h��j��)�heDy�'
�U1�I@�hf�A4.����-B3�IC߄Ԋd"t}�j�!��i�t�Ѓ*�h��P<���D��(O�ԋ2j��i��&��iTVG�P�è�1f�|���H�6j��aw ��Jb4ȟ[8��c֎�!LI&���Բ3����dA�0�|qs�O��cb��K"��S����d��DlڂSL��bM�PJ�pp��O��� �%ZM��#���S��-2�� ��uw��#,h4[W��>�N��'@�=# �C�5V���w.YYz�2��BB<�ZgM��]�u�פ�:7�X< &�ӊ2�6��D�I!P��l
B��s�6MĆ3H4+ bA���ԣs���(O�T��4T��H�f��ܢ!(�4t���JJ�L�4�a�O�Z2MCUEٺ+�駛�J<gk�;(Rx�`�e�5,Ƶ����166�����O�x�b�m�F�ƴ����1�?�sbEa2h�H@�?���1)���P���΄�l�<X�&"<ͧ42��Z�+�F�`i���ɠ��y6�AO����DX&]�͹�)�`h��*^E��ӌkے�I
2:"b@퓔^�� '@T�{����?	v�`ݑ�! #*��h3A"��*XW��R�/]����d�/B�<��q��
{�$��F*l�^�cV��8�
�E����&��k���,Rй��iЂQ\�m �&��6�p�&��.,����ca�ԠH�����B��8"daN6���v삛�T���3bVf��}�J<y�bψ1(�ɗ'��F��1�/D������I�qighO�"���3	_�
O�p&��%e�T����"�p����BG��]S�H�!���K���sE�C�Gl
�~�࣓�K�~]��l��_���qA\���qe֓%~����Dx�%)F�J�?�=X���	��H��xp!��^�Pp�J�ƅ{'2���Ω�����d	�ЊT�\��'"���V8`:A�q������&*ʯq?j4��4;'z���A�K�"���S)-�� rE�9H j����?J"v��vAaפ�� ��)y~�� jGI���!�5ϗr����P-��Vv� �F��/I�p|�*5�:U��4"�qF��O�5��(�9
9ש�.h%fqx�OI�	���]L�p$�C3PJ�����4[Wo��,����	� �BX[R#Y�U�Vy�¦ *P_�
�&���O�V�+j��-��Tõѝ~65H.v}�*�-�����Q�0i���_��	�[=�mh�*D
���)�:(������p����f��*y���=1rg��?A3n �U,�I�]���/m)��Uf+D5����χZҎ�В��.�6�BP�Z!<[�}�!���}b�@�\�BЍ�|L�9�&P�]v��`�D]��Ʉ�3�T�a�i����1�J�R�$4�NLZr ��# 1��*GRC�'����C��\��6Mֶq�6D�%��-p��#Fl�h�`O�M�@��}�b�`OX	I�"�Zt"O�xA�쉪.o�Cь
=f?XB$"O�m�Dj��[�j����j��(Z�"O�y�aGD�%C%��
��+����"O��s�m�K|���E*xڀ�P�"Ox�g
�T��ɩҍ�F��%b�"O$$�G����"��F͎2ET^Hz�"O�y[�a_>'��$M�-1;:-q�"O��J�
N&�" ���k;ʹ�6"O���x��lr�jX�:0Dڷ"O�yi�	�h^�u�6��!f8]"g"O����q��@��ǿF�����"O�)"�lK�|���RV剤d�T��"O�AR@�*o��r��H'�q�%"O��5O��F�>\R� J�Q�"O��pt(ϙw6���gC�Z��8�"O�A� ,�;L�� ���I*8C"O6����+X�P#��%4D:���"Oʝ�C�(`n���E�1Tܮ�"O�ҳ�:3_ $�'{�l2�"O�A��%I�4�bG:L��"O�0$�<#���aB�DJ�#�"O� �x*�j�>kP,$z2�ї��]i�"O�@S��ZB�I aT�.倅�#"OPI��	#u4q�5OBv� ���"O�x���x��:Q�ޑ-�N�Ѥ"O�R$�!0S����G�|���`�"Ol-VD��$�)Zqg�&�"��"Of`r�G��[z��X P�|�� b�"O��!��	Wv�t"��a�� ��"O,$����&����&I�����"O�83�k\�P�����ϐu���A"Ola��d���`�ܺP�yZ�"O��+�G4K8�Ug� v�z|�"O�Xi#��q�(˴@˼'�vt��"O�]��V�K��d@�A�I���P�"Ot���cP��[%o�+&�#"O-q����s�� ��e�:l
�"O�X�aLZ�4㸥!$�d<" ��"O�pQ)X�CV�0���<(�թ�"O��k�V�P, ��C�%�8�u"O��A� {�Ei��7L�B�4"OP�*S�#}v�Ti1���t�<r�"ON���k��>GFlj",�"u{�HҖ"O<<��D�mB.=���<qF�)I�"O����O[���	�	E�m�m@"Ox�(�2��	3�gΏ]�j�"O|9q/E�L� [�&L�~���9P"O���jeҭ��M������"O����l�=_�
��+� 5"O�)���b�����5,r�"O8hZ0J�Q��Eq�`�"$�r�X�"O
���� ��t���Ət}ΈS�"OX��£�@Ӗ��>k��Yf"O����l�T�k&��\Đ8qU"O2q�EP8�Rk�J^ G#�@�"O�m�'�H�:5ƙ8�U ���)r"O���/������P �
P�"O(!v͙xW>HR�	O D��TI7"O��u!_8hϬmZwķw�P�X�"O�Q��Ș�n堥xCŞ�W��\�"O�uI@n�.oж`QQcC/=\P�"O�킕�Z ��Y��U�^O,��"O���4J�1��Z�m�6E�<"O6TDʀ<��� ��� <��1�"O�Un��M�5oC(T�$ZV"Oi3� A�k�V<s.�h+!Sf"Ov�!cN�JM�)I�
#[J�}��"O�P���,wMn�"D±D��x#�"O��1�EZ�\X�`C"ކچ�3Q"O%����";8J� K��va��"O���CÀLV"��"E��P��a��|"�)�ӵ{=RxБ�1A~8�2�Ռn�B��;�v�c��J�	�J4�0/�3��=�Ó�$��&A;������#t[�d��wir�I��N$#��,�s�Ͷ����c,����ߜx�X�e鞇3"D�ȓH�X���>P�Z h�c̆@nl����hO�>5⇫T�@-��
�%+�}P$D9��hO�Q��[n�@�c��1w�8B�	�(1���F��!*|���7&B��U�A�#	[&X'F\��ĘET�B�	D��I�+^�&>�}�u�*/�"=��D�6��CFȖ?o���tA�p�����e�B�)G _f \��Z\vy�ȓ���s��	���{�f��B���S�? nĲ� ޳�b��o 7
�\�b�"O��KĪ	PI���)M~�Ext�&�S��".�<���D�9���9~!�6?�Ryi7-���\�Yq� �nt!��EI���S$߈K��r5� K�!�dƈ8�Ε�"ǃ>JY8�L"�r�I��h�$y��	�0
Nr�9�b��@"�e "O�X(�/�e�&����=�l̪C"ONi"��H�f�(�ɰ \*I��
u"O����H�L�� �5 �:H�T�t"O�]*S� C��]a�E� E��P"O|Qh�g
742��!��+�j`{�"O.h�F$F�d4�Qq�ɬ]�ܙ��]�LEyB��������o�� �ꖢM�����)��'Z\���cC+]��hYfJ��N�(��	+�вH�1� �U�K���B䉋z���Ņ0P-�q �;B�B�ɴU=z�.P�XWA{�S��b�=E��W�@9G#��B".��F��2 ���w�,D��3ㅢl۲82@�ɚ{f�X��K0D��
�#ӝ{��Lx70���<ʓ�hO�S�|FTу�eI�<A�l+7��C�I�$�v�B���H�d��VW�C�	�i $�%��([.dB�ȽJ�bC�� 1j��� N�	�@E�RqB���9ړ$�Z�B@�5z��h���t<��6��8jAH��Q+�q�t�{����8v������R��AO�6����K����w��75!����IZN��o�|�3��.3Z�:���?h� �����1�r!�,o��2�#�M��as��]���?�$�ܺ���$	I�쓥K�Hܓ�ē�y��錻c�hxp��`i������"O��c�H�#@���\�Jt���|��)v ��2� T~P��8�OM� p�C�IF�d�b�(b:b݃�+Ld-dC䉰����CX�t���Yw�H� �C�	�k���Ic�EU��PS�e6+�JB�	�{4�J��p<X�!���
�"Oxtc�n�10�Ԑ�d��K%��k�"Oʵ�Eo	�Ip�d�S�ĕmj6	!D����#�"��ls�Ɓ�,,"�{2@=D���H\\�{ �'V&�dp�J%D� 9&�_�k�d�˱�]��c�f&D�L!�	�Z���°e�|:�b�"D��m\GL�a�O؄w؆�ch?D��vȞ;~U��K��2[<-��"D���F߀�����\+e	���_�<3L<Vkƍ8iE�
pv�$Ď{�<Q�D<#�[u�_(?��p�O�<aӡ��Gj�����Q�<�#=T�á���X#N��ѯĒrO�d;E�'D��R��P�W��P���î$��7�SI�'�Q?Y£�ܭ��T%&D�p\ҁa%$D��7�Td�$����\�Kުe�"D��i�DJ�9�}��D��<�~�x��"D����/Q��Y�-5B!�	 ��xr�3&EV��b��Y&05;�KC
�y2�J���@��L�����՚���?!�L�M*���%��)�Ҭڟb�P�'�}*�F8%z�B�9�0�Ò�y��<1`�
�,ԩ5*{��Y��hO����]π�R��@?=vDZ f���XD����u�m	��D���x���
�y
� ~��&
L�2�)��H�7�Y	C"O�T��%7!�'��^����u"O6Ċ��+(.�ce`����);�"O�I@חR�`���/U���p2"O(����^ܱ��/@�TrP��"O0��c�KC�>$)��� U���"O@ju,�Ĝ���ҀeM�lYC"O��1!�at,@���Wd<�:�"O�9���L5�F�IJ<�[g�>��M$�O��Z7���x�;c���8��`azH<�e(�k/f��i��q�$��	GE�<a#!��DM�U�Y2%�}�n*6Ob�'�L�K�/?7(�;�l�H�4�3�'0�@�T��A�E��>�s�'���O?nlt����~��r�{��)�	�b��hH[�f�tە�!j�!�� �{Qlu�.�f֦�6�O�!��	jX�%�Zl�a�*1]a}B�>�T��]�$��L[�1R��Nҟ�G{��i�`��������A�@U�	bqjP�<YT����0���
34p����g�<!��Q����s�_8��-B�fJb�<	��	'[���B႗F��X�!��]�<����\�5�(O���p��@yr�u�P��m� yv�].�ƅJ� S%�*�!�$ D��Z�
��m�>�qW�7�RT�	>D��q"�!nR �$#�=V$8�#�g;D��{�EM�%?�pJ�`�*p�lC��O������Դ�0��?6�V,3��A��8I�I7��+�S�'�lF���-i��_�j�v���jܢ�R���;>c��c7-??a�ȓu��̀��E�I���s��Z=ڨ��ȓh^�|���'_���@���'+��h�O�DA���M�f��
2IY����'~�yhd�����Tj]�Y����?qI>٥�8�gyr����9��r�D�{�
�y��?I�����*k��X{�����tO\0���ABƜ���e���Q�i	�z��$� �l�maC_.�La�1OփMa|�|��/��)P���X���"�/�O��Fzʟ�&KUp��-xpi��b 8$"O`X����1Ӵ�xe�(xV�`�It�0a�@��x��I�i��PSD�*D������Gr��X�	�$xSa�%D�{1��5]���SG�I�尲@6D�@�0�F�jD]�Pǀ@�ȸ@�&D�h($�R���gƖ߮��G�&D��I7��R��A��n֙:E�&D�$r�A���
Co]>3��Q�!D����P@hbP�f�,5�Z���=D�Т�mt�֍��(�/p4��l�b�<a���L#r�0��K���z�c�\�<�v�¾_F	�MӮN1�=c$c�<�vĝ0���*8K5+�H�a�<�Sdl 0B�+V�,�3��]�<Y$K�:!�H�S� �7OZuЁ/q�<1�,BpNt(Ɇ"�&Y&��[�ILi�<AU�ӟ1I4�A��v��heo�d�<)�Ȗ"�h�3U�ً~`��@�mM^�<�բ:�֬����	X(�$��i�]�<a� K�d�8%� e�6��BT�<)�f\s�-�����vP�4Ä��L�<Q��� f�h�g�Q�5�n�B�˒`�<��CC3B��h�2_�D����FZ�<� �9�a���`ڴ���Y�n�1�"OJX�,7Wa�l��a�l0��+�"Ops7�Ώo��(��!�#-;�"O���C��?���R�Y��N��"O� w&աi�<4��!�Xp�"O��B��ž'Hx��!��>���q�"O�er��TZ����k�q`p��"O���G�c�X���+�qpH�S�"O6�h�n�5%Fla���E]��t��"Or�BZ>4�<�0AذFA�"O>���nS7֝xnS�jL�`T"O^�K`
�ANj����[����"O�m��C	hY��iӋ:�޵;�"O��#$TEA@�����C�.-B�"O�bg� @f��rG��h4r�"O��r�ѨA_�$(��Y#e��X"O���1�W�Y!N$ȔδT	6"O����MK*fL,%�k�(�X@"ONi+ӊ$.�6)q� �1?�7M!D��poԎ4�p����~a�1��)D����m�5(��hRFΉK(��z�f'D�<#��Z�&d,ؚ0B�;IJ�Uõb)D���hOᒠa�j��{M��\�!�d�.Ŋ�i2�ڊ*iB��L�T[!�d�{���%`%YVP���̡<!��́!a\@r��U8 ����nM�K)!�G?3j��Ro�� �8�x�O�2!��;,�ɳ���*�h��"+�bA!�d<C	��C�)�2����i�!���9'"��s��q̠�ĮהW�!�$�/C4�ċ�o��Enx�k"�/Ev!�d�E�j�� �B�#i�`2��4u�!�ƫB*V|Ygk�����U�ܚD�!��B�Z�`Ѭٴ�2	��ܶt�!���)�����:��H���0y�!�6l ֘� �LB���#�6b�!�(�$��/	?N��YY�d�!�D޸(�j	��&T�jh�A�Q�o�!��!.�����"���10�(N!�d]�R fV�Mp-r���4�ɹ�'�.��P��u~>a9P �=�l��'`:��'M�|�:-8��6�0!��'���:S�� <�REsD��%9�9c�'���(�N��N�t8�,4~$p��'�t(��e
*�P!��H�&�6Yb
�',
�����lhr�$�&6��	�'� �q��V�x��*�؍;J���'p������,y�9"�t�hH#�' x�T�>
,`�j6	�}�8���'�<}���ݟR>� ��_8����'*�dcvB^=LQ&�t�C�0ʉ �'l��(�ʪ7]�����+y'jIq�''
���MJ�q�� U�I�p��8�'ĉ���1}0`���bQ2�Y	�'*���&�tW��D� `WVm�	�' ��ZU	"m�D@�4j��P	�'���2$�
@u�Q��
o�h���'��A��hlq�d�^�g�¸b�'�E���9�8���(8dTr�'��`���Ώ!���+0K����'������W��� �O�y@���'���c���sׄq��̠%���2
�'�v��W�tq6,�7�Y.�N��
�'i����랣d������ ^ ��	��� �ux +8�`�����(��"OzM��n�4!&�X�C$ς3�,��V"O��0W����I��� �@����"O؅�ůM�Z�� ���X�N���"O�}񶃇/aG&D�@��L��x%"O~�&�m}����Ūx�j�i6"OH��T�5�8����#Z�8��"O��q���=��M�T��(E����"O�������t�%�d<�mp�"O$��(@��F�k����n��b"Ot@�Ѫɟ\��
��X�p�"ODaJ��]$�$��X����"O��R�0u�
�R'�ޯ,6t�3�"O������uo܁�U�8� �A"O�)퀃~��Ѱ*`��Ұ"Op$2r�\*7ব�J�(3�8Z�"O��e,�2>-+��_��T���"O�@���_�NA0��B�Gq�q��"OXJ���?�D���Ɨ� 8I��"O`-`�,�%���������Q"O�pZ5�	=L��G%�~�ޥx"O*�#�ƵI��02��9�b�J"O.�$I��-���Qa$-V��xf"Ol� �.X� ���7��d9�HB"O�M)�+��a�0��=pȈ(�"O&�Ӗl�3?�<ф���l�M)�"O��RB�>Q^.R���_�1�6"O��ǌZ�]GR-�0�бӳ"OB�:g�#V@p�NK�,�f�y`"O��@aO-R���`uDޝb�h�@�"O�y����&V;x5�C��A��(#�"Oz6�V�wp�qƄ��zm����"O�����	T�C�bZfrA�"OP��DR�Pet�S� Q	���"O����-@�z��$@��E�+��JT"OHI�������B��#���%"O�\pW�ْfb�Ӕ�$~�ZX�"Of\q篗 yn�\��jW��U�'"O��RSMA'K���P��I?�<��"O~0�g���p��G�]�\d;�"O2QK�)ܬ4�dP��@�X�2��V"O��R��C9R�E v���q��"O�x�!V�uW��)�gI+%��"O.I�i�(W-���a�$��h�"O�ŃF��):������1�Hi�"O��֮�G���#��g�ppJ�"O�yX���eKr���(��V�Ĵ��"O�$��k̚+�<��GM�8��"O��)�Ҁͬ�kP��:*���e"O� ��o�:	p�œ4u�p�"O �26I��in(����rm�"O���6/_
D5T��3� R�p�W"O<`��ތ0�����mv�!ye"O�9�'�"&���K�Y��3�"O���B�$
����3�R5��t�"Op��4�ʸh~)�`��J���T"OD!���4�zP��@L+�.���"O\PHЃ�3
 h�+�N5G��=r�"O�� f+;\ɻ��R�K��( W"OB�kd�� @�ؔR/��wd�c�"Ot	A�lۣf�б�C���(֢8I�"O��q��9,:�(�.��d��"Od�Q���8lʴT	�Xu�xe�U"O�Ē��aצ!���D���}� "O� R��E��V�������*zCzC�"O*��J .y
ؒ6�W�9lԺ�"O�#2�Kd.0�+6�ϡ	�Yjv"O����ӦG�0
F
%-Z�� "O�d#@.�<	Q�X$!Ff$X�"O⅀R�L!{��#p
\�<�H4 5"OYs�I��"V=ꡎW�9<�	��"O򠻒$��J]A%���E,rp!#"OnL�S��6��! N
'!ƍz�"OJ)����J1j���H&$�g"OT9��蔉�2eƁo� ���F:D�L1$�D?2&������Qy����3D��OG6��i��ŉBDq��%D�4"��r��両�ƪ?j�`�(D�LB�+@�;��I*A#�DA�@��O&D���p�O*�iI#C>FB����%D���c�C�B�,��%}�d�g��|�<qb��<%�l�9�d�0-�Vё�F�}�<y��Y�,G�h�Am@0>HH��ԯ�C�<��"�1R���*��u/2!B�<�֫"w�Y����tς�d��y�<��Iw�:�8� L]Վu�Ddx�<�pkB�#K���5�J�	~�͉�M�s�<!�H N��膭ۣD~�Y�Ar�<!w�
�L���	�E�|)���#�V�<��Oˈ/$�`���t��Z,Vz�<q�c�7;�A�D�%�\]�so�<9�̖:(
��f�����%�%lk�<�`�͝E �%Qr@�<x�����b�<)��L'ͅZudi#
 <�f%�ȓ\�5�u�Ahh�㦔�@z��ȓ]�p�-F2pE�q%:,�:5��Y�H)iEdu�Ҭ��	��z���}����L,s�v��#�ج%�V���G��S��7�Jc��(0^H���3Od{���,�4a��c?F�Մȓv��S3*R{��9�����H�:��C�܁�r��:VF����u��[2�*e����c�
�.ҊІ�/X��㔭<�2�	�i��Zf�d���]yuH
* ���4iƇ-̄ȓY��$#��	�2 �"�H�\�(�ȓF��Ѥ�ApU:��U�/d�ȓ��DypK�^ �x2�޷u\̄ȓOtr�Vc�;��1�/�<d��M�ȓ�"q3��_�u`�.غ�2��ȓet�q4I_R(��C���`�8��F��̀'�!��K�훖,���ȓU���-כb��MAPi[�\�:����n`��自0��eS�-P�D�~Y�ȓn�0�����@f8�n�$P�f��A{8���bCXp��v#  h``�ȓ/;P+u�݀L���BßR,ͅ�_w�U��ԟ^�*�(փZ����pF�0U �7"Jd�q�^9p���[0��QP���4���4E��ȓx�T,#�杰5T�IE�ƲfQ��� H���3��8�ɗJ�Z~���] �E�e��:글�
S
_�`��+�����K e�)`�
��,��.ۆ� ����`���\G�1��x�i�P",��VNKЄ�ȓN5|���ro�uw�@d����1�f!���3p�2�(�?e tm��S�? ���$HB RL���� m�U#�"O��B��].#���պ&��,��"Oh�B�n�2~�^1��JcuD��"O$l��IB+���Ѧ��>mR|���"Ox1z��W8����P�C?l�!Q"Od1��K2E�����L�:'���"Oa�%O�81��q��a� 'j���"O�A�*�= �"��T��TUb)c�"O�`���4G��0�i�;VQ�Q"Op��p�� f�{���8e�v"O�tc"B�#LT�-˞~+n���"Oތhu���Z�Z�˹yx-�"O�!qai�5o��H@n�# �����"O4��q"Ҫ#+x��u��>:`X�"O�d�Ƃ=p�,���\�	�L�҅"O���E� m����#�Xb'"O�0�Z'�`z�B7	��Q�"O�}�5Fv�D
QH��P�J�"O0y�!Z�%0�����$|����"O������8�P���\'�e�"OL��w.�4w�.����F(��{5"OV���oN��X���K��a6"O؈�pƜ_f6X�bOآ��2"O��g`�X�|��0/Z�	k�ԑ&"O�����²}���t(�YhQR�"O����SILv�9��
C"� P"O	W� |`�������w0ؘ��"O��##(T�s,�e��+��P����"O�dHT�<<�����8m�
�"O�8Zf�%��RV��}�Xq&"O����ON; ����f��R�"Od!r��y��Dw��Q�=�"O�|��M�(����0j�g�ec!��w�>(#��M�ؘA�5��g!�P�@ub"ɜ/1��N�/e�!�޿-�1j��ק1�Nl"D���!�/�D�p���+��ԧʥ�!�$��&������2i��سTԕ�!��uB��8e��	����6S5�!���5iU�� CNo�|����Z�!��X�~���D�&Njh�! ��5�!�D�T�"Y�u��,^4p��b>.�!򄏳�� �$#�H�� Ѣȫ�!���.<�`��b14��&� A!�d�F�t�a�
'��cVk!�d�"aծ-p���2$��)�C�!�$�F� s��N�GH�܀�U�!�D_�o5��1ӌL	EJ��A�Hxa!�R���JN�}�T��@Y�Q!��(���R#9���x�,%?!�$E^�h�0�͙\Ϝ0҅hF�(!�$Z,�2���f�4ƺ�!hɮ9!��OFi��<`��iJ�'�$!�d�V�q��F�)�uQf��'�!������aP�/Vd��"gM�E�!��8aP����wKj}as���S�!�DL{l2T�1�!'9F�#K�|�!�$�<�"T��X1	Q��06C��K�!򤅔Sv��'Dt�pV�4q�!��S���G�2���4G���!�D[Ah
{�e)v%�Ȱ�Ȏ
x�!��P-*��%�Mmg������ o!����|���Qd��{P�$�� 	4Ve!���>G&d��� �`�L}qpi  O!�� ��� ���|��d	����C"OɁ�i��l$�`��,��;@"Od�J�H��l��hH ��Vp��+Q"OD�0gMF.�9��i	�"���;�"O�d���i�L���o��	�"O:�+�.�H:�lGX^<�+q"O�F%�[��k5L�o��r�"O��P��1_B�<"W�Փt╩�"O ����/ּ�Ӆ�U�Ss��"Ob5���$v� ѧ�\*eѐ"Of`���*@zH��¡زh�Dö"O"��ӭ�m�z�X��r�t��"O(��AY�l 
8J�OR���U�"O8ē�#�"*���®�' ���"O�q�Gס	��=)A�N�!����S"OZ�0���z��Ɵ�s����g"O,��'ˋh��"Si��L��"O`䁄� b0i�#�m6����"O�z��
c�X�f��J��d"O�񠕦O
C��x��=.����"O���#�E�Z����IZ���RR"O*�1aÜ �|�#CW�)�M��"OR��Ǚ�#�aA�h˖z����"O��i�ڡTҊ�0EJ�1,���c"O `�B�ٵH.�s2�+6Jb=g"Ovp��螛@i���'BE�SS�8*!"O���-�6cI�dC�@ݛ4>�y�"O� ���ig��*%�)q/<���"O���D�� �nX�!m[�X �"O,��_�Ms�4���,��e"O�Ic/RKy �'�� ��""Or�ؕŌ	V�.��T
T����g"O�D��M6$S���$��- P �0"O䈰�_�)���� �_@zz�"O�}K��&�3���4+��hK�"O���smQ�x0�m���1\�4��D"O�=���
t��ȢC4%���W"O�0;�a�6e �A@���4(��"O�"��E�^p��N�(��"O�E#2�&/�
�2N^�G
"O� �uDپF�F��$6�3�"O��!��j��p	3-ȪddՙE"ON�[�#�yj����ĠI0"ȎaU�,R�ru`D�(���"O�8ӿ�(�$�#	�EY4�M�y�j�W�r�b�F��|��0��W6�ybbSπ��1F!DtD��y��W� f� �=/֤48rEL��y�+˝L�n�Წݐ7�	i��1�yҨ\�@��	��^*��!�7hO��y�Ǝ�%M��@C�O��A�Ga��yba@)2"]���
����6Kޡ�y���.y�P�EM� � [sGO��yB�]�d�FMs��T6[3����y�%�4�<�����< L��B�ɕ�y���*Kxn����7�)u�D��yb�˓iz�Й�&��E� A�d��y��\=B��&��lԌ|`F�[��y��݁RF�����*:� ݺ�����yR���ΙJw$Z�6��U�����y"��D��HԬe~�)��$V��y�ӛE��(��Ƨl�,8�nI��y�.Ň#|�Ȥ��k��`����yr Ľ`�t���c�[JZ]��c�,�y
� �BP�C�[�>�qL^x?��B"OXPH�.(�!K��0Ј9�"O�`�"G�����Nc�&���"O��I\ M�@(�OF*y��0f"O �ѯƢ|0mp�N�J5��"O�ܣ�`�3[�h+B SD��`"O� �G�V�J\9���<~P�"O� iV$��=�QQ$ЕN7걐�"OT���K������L+�"O��زj�,fV6�V��l���"O�p��+G�is�eu�,9�"O�2�%��)R5n�3���"O��1^/�J�R-Р@Q"O�ib���R�)��N�/Q���e"OZ��탚t��}B�F��"�M��"OHЋ2��{O��I6F�(��C�"O�#�ɬ$����N�0���X�"O��8�d� ���q�h>1��$K�"OҔ�䊕5vO�AY����{"O��	�a��~t3�o�7_�JLb�"Ot;���#v�!J�CV�6�y4"O���%�� Ĳ�Ѡ��	�,}(E"O�����8��P���{x�4�"Oұ+���c�V��si j�U#�"Oڱ�c~��� v��%]^��5"OI �fE�@�h��f��yTx8��"OL4Q�S<D*��b��<�nd *ODq�`�1P�q���$s|N�i�'8d�SІ��>̅{e�ڴ3r4��')��z��Ӄ9��ik�X�8D�i��'OR��A/X))��d`U�.���'0��Q珂)�l�tn�!W?�J�'�<�öl��L��l�K�%U!t8i�'�n�J&g� *ԑ�bI	����'� �%�&����X�F3.��'���چ˟2!���"=Ӯ��'MpX�f��r�������kސ��'�� �a��77&=�`�_�|(��'>�p�@��9� LXE�c,%�	�'����"DQ�Dkģބ�^0;
�'���oՍ����P%�,@}Z�*
�'K�5���
w�fT��e�9No��'dȊǍg�4;4����e֣�yB�΁�t-�� Y�+����H��y� 7�( �/ ��4*
���ybg�	j�xr'_��i�E��Py2�@X� t���ԕZ~��&�}�<̒ L��VI�:8�>�ъr�<i������	!فa򸔚R��m�<Ig	E>Dvd����?=j�2�nl�<Y&7< �#"��EB�B��h�<��Am�Ѳ�.�� �ް�͙`�<��gD�j��"�P��%�Z[�<i���M�1�̘&J�N�CoXV�<!ր�m�b@K�ύ�*�ґ 2�	y�<�a	�:;u�9ȅ��dW� �ύ\�<����b��)@	��� (�ɓL�<�Ňɢ~5�WNP8^�
 �Zb�<	@�\C!�� ��Ȭ1��Ta�<�㨓�?�1����.L0< ��Z_�<��FT5R$MH�dt����`�<����X����q��
Ƥ;%�v�<a��ݮj�XHzE��
d]t�IA$Eu�<	�A�$7�����}1(� ��x�<� &�&lE#$ȼ�5�	&uV�(��"O�5YC�Ŋ@~�� ��
N=����"O<|�$�H�%8�GB�8v��e"O8���,M��pp�㒦�6"Ov�:1G�It�x����}��p�a"O�q��A^3*�r�ȁQ�dD9�"O�m���
DI��*p�E>_�T0K@"O����$99jxc�6�,aP�"Oj��4��&����W�ǘa~ ��""O�����
Q�T��FI�4e���F"Ol�����?i��G���Gtx}d"O4� ��L�9�F�A�eR\H���"O���-I�o�}��j�:Y�^źW"O�q��n��N��t3j���\)"O��i�-8�\����t
jY�s"O@���@�[��S�H�9.#�	��"O�XA&�Mn\9��G��!V4�e"O�(X�#��0&��M��&��"O�L1��P�0F�X�A�K�|p�B?!�d�)@�qӄC&� q��^!�ėv �%3R�,�:}�f��3�!�d��5�Ĝ�A����A�nC�\�!�NH����M¸Fsle�,r��C��/dS�%�U�����8w
�q�C�	#���Pg��"��L҄a+Z�C�|��G5[p��%���@0�B�I�E,�	�2��L���B�	4^{�p�.����tk�8~�C�ɒe΄*B�۪\$�4B6N�"rNFC�	T�����?-T|2�
��DC�	x��e@�
���i��s�C�ɶ=��%��m(��9���+��B�ɩq��mK	#܊tz�!�3F��B�ɷ�Z�A� �6`,�����C�I]x��
�"�(r�`�%@��X4XB�I�?�$�ceW-8��ě�o�q��d��U�xV��0E�.���"O^�
�Ə0:� uhA��}�$��"OL\X���A�+L�`�j�z�J�(�ybh�=���ᄕ$S`Zh�3��.�y���p�Vu��mْS.(k�J���yb��}���T� � �\��C��yR$�3/��\Sre>l2��]&�yN���U@�npx"eO�~/&���jpl��D�i�<ę�
Z�<�I�ȓ]{�h;�' �&���"���C�ԁ�ȓ4���r���
b��D�$�;��\��tL��G��A/|!���*4���GQ@<b�R+-j�1qk�
��ȓX�n����ۯr6YɁ���oǊ���-�-���ɇ:�����>D���ȓY	��"  $���b��.�]��	��dS��_�w�����.m�	�ȓY&�������gǅRK�)�%D�l������с3nؚ,�~���.&D��Z�ǟ7�p5�0E��o�.YJA1D��$��S�����:GjI���"D��#�ش,��@b�D�dS�,D���1��d��)�M!o���2h)D��;G�94����+�v�@&D���` L�g0)����/~\�R/:D�A�M"D��Q��i�)Y[�\c�8D��0�f̴"����`��5�}�%!D��Pd��
do�!�d��C��|`�H D�� ��cm�6��*�&�-nF�"�"O~܀ G�:&n����B�wi�,�w"O.@�dBI�P!P-k�×�5d�A�"OP�h&I���03"��U�jU"O��I'��:f�"M�AR���"O�9sQ��T����q�-!h��"Of�`�'�#b{��N�(np9��"O&!�2	�c��#5�H�d8�"O@�+�b.���r�Â?8��D�4"OfXP�
�1��պU,��j�*(�"O���/]���G��*Ѿ���"O1�Cˎ h(�$�."��P�5"O&�Pf�21f(�sǣ���s
�'6,=�Ȅ�n���BX+���	�'/��kc��MQЧ|�^���'Q�y.�\�D/�yt`�6Ÿ�y"��!LfjJ0E�ʑ�Bk��yBhB�W(�	9񂗪Oi$L[�	L��y�@i�}����L.-��d�.�ybS!�� c�*܁\xP�;��y�JI��q�֦�?WSd� �˪�yb" �Q&yHc�:A���1�ȝ�y�m�W&$�� ��0d͚�
���y���3���^�UY�ݐR���yb�V���h�	_�wjU����y�h��t,�0��KD�1hq�!Q��y2�	'��A��Ⱦ+�E����yR���X���
�u�n�1􆓝�y��`aW���Cp���·5�2���'��YE0�����R�-�س�'5�������WߜИP�m<%B�'�|�+��ݤ�鰡�7f�0y
�'
�h����m���@��=e��e��'����@	��?HFx�WoD�c@�l��'LD�8 ��+_�,�6�aָ+�'�"��.��-���"����{�'�"��s΄�j򦝫3a�{����'��䂎.8�d�J��wΐ!��'�~!�b��x����@��cnƩj
�'|�y��7-��%�(�����'*D��e RL�XH��gF8�y℔�/T�ɫ�%R����1i&�y�'@'g�\����$+�:	��\�y��B���D#N��(���,�y��?RײD	w�IH
��.�ybG�!R�
��7�
^٤0��/�7�yb ?STa+���*J|�]� M��yB@�K�љTI[���@@��&�y�.�����QJ� Xi���#�y"�m���%�+�tQ���]��y�E�7:x�
f������Sp"W��y��.'@6Q�!hQ�g�n�'#���y��Nڥ��
� I�'k)�y�N5�Eeή^��C�ϟ�y���j�f� ���U��3B�F��yb�+:���K@'�U�t�c���y�%ǆeF�p�Cx`<��F��y���^Ox��b(Ȥ>,"\s�M!�yb��k�\�w�98u�)�� JA�<Id��"IZ!�U����aѡ�q�<Y1i�
b����Uޕd���2���R�<i�ѱ/���2 ΋�8du2$C�y�<�v�0,E���4-��r|
xruu�<4E��U$��L̬�P��ʔZ�<� 2|�bo�,�pmR��K���Rc"O�b5j�a#,|J C&��`y@"O(-'G�)~K�bN�]��Ȱ�"O�)V���"�HÐ�� qw��c"O�-�L������i�ve�p*V"OHP��j�4�x�C�h\�u�J؛b"O�5�J�(�.H�U�{L	�"O��g�X� �<���H7#
��"OʌsVl�#��@1$�U�V�H�ئ"O��cR'��Y�H0��#���*�"O�$q�G�I0��g"ߣb���R�"O�E"cّDr� ����^�q"O4!9�"K�a 8]�W!��{�#v"OF�AE:G��@.4�}
䭋�{�!��K�T�Ȱr�˝"�44+�Y�}�!�dD65��9�dL��&���1�k�H�!�P:�,T�D�ͭp����ӋZ�_�!��Q�M��p��a}�m�*��M�!��36�����^*il�"!)�(e�!�*\S�h`T�1^`�a�ȗ(�!�d��T�"�#1E�@�GY�&�!�$M*�LH3c%{5�j��<1�!�-�`t�ʐ+,~����SV!�dg����S��4: ܈t�KO!�d����	7�1��[s�76!��3u�*ձ�	�{�H�(��B*8!�$��Kl\�!F�T�D�F�.w�!�$���M@�#δ-NL)����7<!���G�~Iâ%�9c��S�@�V�!�ɧg`�$���M-.tc1KO
�!�D �(�0,�S�X���W1O�!�d����BЬ	;Q�%t��Kc!���ohD��\�NL�Y���;Y_!�P$A6���W%�!�PW�[�`!򤔶p)�̐a����)�Õ�;�!�d�7W2����(�z�e��!��vք4bk����U�O�-t!���A���B�	��J��U!]l!�DөO�li8Ī*�Ń�D�U9!�$�� TV��1/K
|�H�֮5�!�ą:O9^ܣ�a�+8ePq!�O�!�$�2O�v-:��&ecR]��$M!�DF�+�R�p��U���͌�Q!�DJ�h��4(Eh�lZH'��5]!�A#Z��E�C�;S` ���W'?!��<?%��I�= S��zpÒ�
N!�d_���H��!�3}�0�3��o�!��&��t[�<�8tN�Q�!�� R�~����	/�x,I���r!��ִ9�Nh� Ys�@@��G�7p!�t	.h�r
[�c�n�ˢ��7^�!�$B*%��U�c�Ǝ~��� aN�W�!�d� �̔`&&�3;��[G@ !�V�(^�*���4Ux��ɧ�%NW!�䟵$��a�#h�x_L5@UM>0!��m��e�d�ǌco�e� M^�l,!�H�<`2-R��^lV(��!#!�DW�:�Bl���<Ha��IQ
̡uj!��B�:�	�� ��Pg�t�	�K8!�DGC
�P��U>�����, 5!���(�����I�,��I���1h�!��Gr��1��C��K��!�$��oY� �P&�	5��� ��!�� \�`��C�̔١Ġl!!�� ��B�Ȯ<ݮ����]=���"O���2X#y�X�Ѡ�S�V��"O�񃲯&H5bx�D쇈z�&e�#"Oi�/, ��s&�_/~T�[w"O�����DX�������7"O){��Q=`A�$�)�.8�"OJ�I�,�A#�MZG��8�Y"Oް����![#
��7���#�И �"O�T��)ѩ�ZI��`��A���s%"O�����-'a�36扻j��T�6"O&%@��(l]X� �\��&"O8�;Ц	M�(�v�V�F���"O�܈f�M�[$ٲv.��1��"OPX���|]x�v��+�����"O� ���M�V�P�sԭ�#}�N�1�"O�5 �B1�(����.(�|�s�"OL R�)\*B�䌕�|2�"7"OX0@4lţ0�f��!��Ov�E�"OX)�`��(���#�Y63R*䐆"Ov�Q��3�HV�Y�[2����"Orh���K�VŹ�)��!-xP"O���W*�o��أ�Tvt�{�"O�Q2�?zz�e�'	��X��"OD��Aó>A��PpF��@=��"OL��э����S�0q�@��"O´����#OH�Ա��ʶ2�"-�D"O�R��L��b%��ش0�h��D"O�1��U!�^�����JP��;"O�Ɂk�hd"��ܲu4b���"O8�S�&(;^�E��0u}8ix"O�MJ�E�f�L��ĮAq��z�"O�t��X%:\��FE:7�!y"O��!m*5+pd�
�&���"O�q�)
4�h��C^>B�X��S"O�d�\�m��|���5kڌ���"O$1�Z�TGgJ�h���D�
�!�KX�q�6��cN�D-§$�!�/!^$�
�k�f�$�����&D�!�[�M�d�C�1Ϛ�0t�s�!��	*G��c��O<:tJb��� o!�ߜ[n�
�㏄�M���37�!�d\��P��N#-�����ګ[z!�$����2��Ǩl�h,Z�'!�G9*B��u�_���\:�Hu!�� |��"�.��e�ԥZ�G��!�0.��i�Hs�2@u�P:Hc!�D�[p~�z!���S����W�`�!�,�����n�o��"�(xw!�$H��$����Q^$�z!��3
v!�$<jׂl�'M�>YF6����ܤZ!� %=���q��H�:ٰ��&�̻nT!�$��~�,K��9u��@�K�G!���\
�u��DD��>(A�L�!^6!�dۤz,��#�'9�T#�� *O!�$��C���beM�v�: ���#�!�D
�WR��$��}�-�PO�Z;!��:K�l9�Feڢ��!��h�e!�D5GD�`�N7uk�`�����W�!�D���97!W�rM�E�2����A�7xRm0��L�N �o��y�L�*��*�$A�?
�Q� >�y�疑_�8�J�(݊8�|u�@��y�gϳ)�|
��x2�)������yb� P���k��Ǉp��p�A�"�y
� D�s!)�E�a�,S�?�j���"O�3���"4	L�{�{g"O:��ӆ�
r��It��jfP�"O��[��@�h�RC���F�p�"O�5�V�%0��X���[;��"t"O�0�-��y�x�a��J��&"O&��p�%ˆy�E�D:H���E"O|I�G�*o����@
]�b`�"O���1.L����9�%#��ę"O$¶�Z�D:ڵ�T�]�p�Qxt"O"��ː�X)X1�D����8 �5"O�� �a�3�T���k�~"tY��"Ophs�霽0�����K�5�(��"O�iB�"�,���4!�_�JX��"O����#K�85�T��4��"O���ƣ��@,(��.�;�d�"O�����&��	�N�&~�����"O�K�/Ape3��-���)2"On,3�&@"`�b��#��02��Є"O�=�RN���Y8�ʓ�e�~9(A"O���t�؝M d�0@��9-�)�""O`�b�ü]^�#7@WB̜p"O�`ef��HT �@EOޑ-ڽ �"OR�K0�؉q�0�5�ͫ(��ب�"O���;�"��p ݙ����T"O2���hʏ3�ybB-��x`ɑ�"O��b%�ӱ���+�KĹs��Ĳ�"O�|Y$fOF� 1�U��m:�ɣV"O�`�F��_��A��-<���"OZqk�d��Z�4�P��Q!�8��"OT�{�@""�ZA�� T�J��"O��	%b�Z�fAr��t���"OX@QH�b������lx.0�"Ofb��e�����^65[D�+d"O��PƷ:�|�b��@��d�c�"O(,����2W�1S��H����%"O8�I�FZ���}b��Ӯ,�@�p "O�i+r���S�Zl<�-��( f?!�N�~�<!�a��2Z(�X'K�s#!�d�	Y�ʍJԧ��QI\�K�d�%s!�d��3���fk׺C8�Qy`"�(/!�ב|�T�@f�;L&U����G!򤉊v���9��P�^�c�΅g�!�d�g�fM�E�Ɏ����2�!�D�&SYrY�ֈ[ j�� ��!���;K~���_#X�s��/c�!��
d��x���_��`9�;j�!���&@�-�c�I�&�P�U,!�q�ڝ!��2�h�zU/B�.!�$O�,, F�<m5d8Ӕ��q!�$^+ �̙��ْ .DҀ읢r !�d�<P>(��c�6+�e!�D7g	!��T	h�,��$��
*��w�<%Y!�ڭJ�I[���>��Mh��6l"!��(Fμ
�3��8�^�5!�Dq���h6GC���Ä�-w!�dէwF���6�ٛx���b�B�r!򄗟n�,,��$�(�F`q��V!�� |[1%k�'Y�����Z��!�Z�+�PB��X��e�-Z�!򄝹|��%4c��]�T]+D��
�!�D��1�8�"�-&�nH�\�F�!��~�L���i��4�dl3!D��!�d��W��7��*��	1GAA ;�!�� L]zA��zk�	��'�g�AB�"O�! �AB8Y@��Q�[�Z�v��"O
H������!��EX�4���"O��;#G�Oۮ�P�D��{ĴyU"O�����Ϝ9Z�����1��@�U"O�t���جL�<��U*�a�>yS"O`yX��|�ɰS`�6���1"O���ÍY�k��,��ųY�R ��"O\��g��A����,T�n����g"Ot��W
�7+�HKAE��n��"O�H�e��bPűt�Y�N��Y�s"O�X��L��RX��F��D��t"O���\��jY"��Z3y�L�"Ol+����,�4�v�.C�pv"O�7�F6)��t1�L� -i�'�&D���n�H��Rҥ�E�ڽٰ�&D�@�PD�M.<+��S�k�h(D�l�i�)���kՅ�*�1#Q�%D�#'��¹�`�B�x��i�W�$D��8e���/Y��#�("i�Z��!D��(fn��`i Ɂ�N �R���z�>D��������X��ҫ�:1
��;D� ڷ�X�C͈�7+P%X0*q��8D� *��^���Yw���,�4���6D��qEK/7BDӦ`�	J�����4D�� K�>h8J�� H�-A .(D��yČؙ>*�q�%&�$A>a2��8D��BTm�)�@ʇ�,A��A$�7D��ڄ��(YDt:ES
��6D�`��dȏ9u��ǌ*4Ĵ��5D��F�KP���b�X�!�|��(D� 1�i� 8�XxZÎ�
���L:D�Īu�� m��36�ϡ.�X��0J9D�l7*�p��U(�NQ�ۗ*D����;�� "ц��P�3h�W�<i�+��Q���9���)TD,z���R�<Yvk��8��ܑQ`� ��I��c�i�<1���%�)�#�!+�"䉃h�<��FƬL���0`�*��|�<!Q�M��us!a�5��IĨEz�<�T��+f�I�E3�X���<����"k�le���P�a��@iv(�~�<ٷ/Ɔ?���� mSJY!�t�<��� ���iWX�8�`a�q�<�@ :=F���-K�6�0�f\j�<A��[��t!7#D�>E���b�<bB��a�Az��|40x�$KYb�<�C\�G���*᫜�cƲXA��]�<у�[�c#f�0�+B*"Q2�kpc]�<�7iD�k7^��rA�"|[�uKU�<���� x>q�� 5Zv��!.
N�<闈��ZѲ�X���30(.i	c�I�<Y�F:GTE���S�vr�%���M�<I�,ݚ�~��sʡ ����hIR�<�lQ�Jx)�L�gk^�(�N�<�f�bD�Ƀ�H?5*JPp�O�<q�fj1 c��ȣE���!�d0HB���F�t;VuÁ��2!��)?�^���B�t|8A��
S�L�!��x�̳��N)Bn*�j@��!�ί&n4Q3�
 SN��)^�O�!�͂���y櫒9R�@Y���!�d��\���+�2��Q�e	�X[!�$9m��K�C�=����@�M�c!�� ��� b��4^.���Mk�<���"O���CK��M��PYӉ�"���9"OЍ�n@�@>���sț%c�r0��"O`1yMQ-s��V)�/�X��"Ox���	�Y��|�P�D�d���"O��J���0�(
��0{���'"O�(���k���i����ju�}�w"O��Pwc�ZN�#)�-:�MzE"O�˔�U�#+�ؐ��8~�Y�"OP9C���,g�Y�r��/�n�Q�"OP�8��2>H�)'�M ]�"O��T��Mk���/�2.�b�"O:\�PG\�&��Țb/L�Q4MA�"O��)w�Z~q ��/+t8�#"OL)*$oҾ[��$2 �}4�J3"OةpA+={�m@��\?s�vC�"OH��@v���6aH�`�p5��"OZh`��xl���@a��f���""ON��C'�{�r�� ����t��"O���O\4n۬q�0�S<	�,�2�"O�0�F�0 ���H�MA�|���4"O�аwJ�?�R]�U�{�"�� "O�	�B�! j��S��`q"O���dń.�4��K�J��i�t"O�q�g��(��C� �u!u"O��:�K�xp�Y"��Qc�"O��� ٭jQ��KA�TU��PU"O@(ZE]0'�y���ĂD�493�"O&�S�nX�^~�:�ʛC�>q��"O���4�̺e��(���(:�0�S"ODA�`ǭr�-�e埤:v���5"O�!X�':0��!s����arʵ�""O4@S��гde�Ё��
�`���"O��k��Q�T�pia׭���<�z�"O����" _xn�ac��:z��B#"On2�nʍ�R�
��ܗ)�ލ��"O�Y��i��r4�m:��đ\:�h3�"O��m��F����tK��r*�m��"O"(���� �B�jJ��6<� "ON]ad$�6���Ssh�G����"O�U3�J����Ʋ�0�"Oj�Q���9d�0�E���8h�"Ot'�sIhWE��p���I �y�C���.Y�7)C;8ڱ�7Ɯ��yBj�&9��A#�,	N]+�d���y"*��G�{��́(?ex!&�>�yri� ���"B �7g`yѓ���y�)��P��)��#1N�h����y� T(�fC
^��`�&����y�i�KerL2G.�c�Ġ�i�?�y��ɭoy,�ٶV �9�Dڈ�y�,���,- �@��?sx��tO��y��F�;��5PC�?5��(CT'Z��y�� WÜ9�W$Y22�vĐS���yrJ�=9��X�U!t
@�S�W��y�F�oMX�AWM%Vv4C��CX�<�ak�ԥd��`��(��MԞS�B�	�-|�@����6��"�F8��C�	�n~v� -��{L�X@13DX�C��>��H	5&�=L��a��M�hʄC�iƆ�q@��n`8z�"
�9dC�ɶ3j>����ۡs�A+�G?RC�	,��� H~��Z�#�D�f�hO>��� S�B�8�����B�X���hc�Т=E��t�? ��󁎅;I��)�Dc� j)jDc�"OxA`J�6\<�[P��{�Ȃ0"O�|{�'7����4�ݛ2
��k3�IzH<��嚳E���k#��)a��(1�
�~�<!㓣W]�����)*��Q@�)�D�<!�i�:�b�b���;h�f�:���i��hOO�\ہκ.I�h3V$F�r���1"O0��2��1	r�ZG��d���Z��?�S�I_>-��Y����00���g҈a�!�$L("����ʏ$���p�t�!��F	�0��GֲF\k�&�0)�!�䘺I0<��W�䴠��K�!��ln����W_ ��hb�]+4�1O�=�H>���^	"�zq��Q�5bP���d~R&V�6Q�b?��G��)@L3��30l���0D�X�%�����ի�-p���PG/D��b�D�'��q2�5`�B�"�(�ܴq�6I+Â�,'��铅!��>��Ԇ�-:�E����v��C��S+I��tFy��O�0����{�����jZUӤ�S�3�8C�	+y9����@����KR?<FB�I�$��x�Iʾ)�= �F�L�hC�	Aͬ��C�� _���	Rn
tπc�؄�	*���Ī�)�l�`t�Lf,����Ig����*X�dG�}�U�_�l�&x��0D�0#B��As��s#��8�BP#��>I��铤(�����MT�s���������xʓ�hOQ>1�u�\�6Y�A���:2�	���!}��)��7?���ᧇ��ZDy3�U�3�C�ɦjXf��N]���������B�	:<��5�c�bN�y�bθB�~"<y���?��"	U_���gⅢh����#D�4��	��zhB� ��6U�a��!D��`o��];�(1�@�J���I��>D�ᐈ��n����09���P�<}��)�ӤL����1�A�G[�Q2A�J$e���I#*��G��&�<Ԁ���3䰛��ʀ+;�C��8z��@�ݪ��#��OȒO|�=��^�:\��S�&��	�
\�Z���=�^e��� I&��Q��X�(�֑F~2�S�>�+�(V�x)�tK��y*�'��$)�4�'\ꡨ�&/6�Q�×r�H���}�|��5�<rAn��K���BpDxb�'ΘɔG��Ē=�s�ٲg�&4R�'9D���CݔW���Wa�Xن���'E8�[����!v�Y
 S"$�
�'2Fq�4�=L���K�Mmti�'������(��E�c���S�,�yr�It���Q_ �Ӡ\�aѡ&n�2��ȓ)���V�U7)��ۖ�[�K$<��?��4�p<a��C�&Ka+��u�E&]�aB�/%	��	1�ҴZ6���G��0) �{ғx2�	=<��(��o�;�t�BvFی� ��d%�	!K��ㄤ@HF�)�`�.ҺB�	�t���1��֟r�}ypj�(\~�O7�3�Sܧ ��ͪ�&	.XV�L�R$�/?�,Q�O����Nz*�M�u▓��宊V�����t�dX��N�.[�(�dG6=����'�2�H�):�p0VmM�xo$��'����$A< ��9$n���V�`
�'P:�c��N`�,@�s�S�z�b�S
�'�,������ڡS�zl¬��L���)��6��Z��Y5�,x���Ԕ8�僀<���B����	�D��S�? ~%��ЦB�;��E����@"O2ł�#5b(��f�<�:��2�'U�dA��y)�C�FG ��5�D=�!��ѭ#�Иr� Ӹ:J"��jg�!� �3�F�0B�����Q�axB��!C\�4k_!P�d��c*T�jC��&O2j�K�=�&��rE�yuB�ɥM�D�sDo	eRx��'_5a�C�	�qbT!*�J[�� `;�"QԒU"OtTR4οB��KpE�7m�7#+D�xD�Ӟzrl�+T�E�k�8� �'��O���O�|�:SMf��Y���8Ҫt"	���D��n6��� f�xi(b�Ҷ&��'�ўb?�P1$ݗz�Lu0�2�rQL:D�H�i�x�59��U6U t�7D�8S���[��(���Z%0����R�2D��9� ��zS��:�L�;��Ȣ��0�O:�v@!6'�7Obz|	���9<����[
<��J��	� S)�.�%�$D{����!y�Z�2dֽD�V 	�A��y� -T����46򊜱����y���/tA�T	f�%6�rA�r���y"-Sj� �&ܡ:>���^���'Uayb�5=\��6","��p���E�"C䉮+�\��5%Ҩ�X,����0��B�I4Z��
6�޼)a�C��	s��">����ؠ%[��#⮜;7��Bvo��sў܄�I�qRQ)T#�ht������
�HB�9K�}q��@~ΥC���BB�*E�r���A�4��9�v�^-i����D��,Q@�T2���'��7x�r(��9D�hy0o�Zg \�T�_(Dr�d�cϗD�����dM-�L5���΄�-��@a}b�>A�a��o$L������3e,JD�<i��TŢ����-���z'��g�<�%FƈTe���o�D�ƀ`*�[�<�����Wr��1@l��b�G�q}��x��Of�>�;�P��`;*d�"E�N@ �'�4�x��HD]��LݯD���Y.O���$B< ��e�R��#o�f[0�Q�d�Q��Dy��]}��=�J��!�?D� C`�Ǭ��	��p>	ħD�:t:��#���~�S�
H�'Hb�DCs5����l��C$E �쁧����`�x�OX��v�h��7��/-�tAG%!�!�ش^�8ت��ɥ~��a�&L�!�R�F�4
��<N�J�Y�EC�sg!�0�����/�`s�4jW�V`~!�:ZD=3g��= �Xِ�Ƿ?!�d�9X� ����?w������R�!����i�m@��xa���ݥ"!���4�.�FN�k`�0*'c�>�8�O�%sE��%���;j��""O80�JF.']��Rni���c"O�@qեQ�Xd����l��T�vT�"OF���P'D%��r�L��=�p"OȔ u���;Se���A��"OH���Rc�%A$�+h�ִ��\�$�$4�Oh�V��`gD�˂a�-_�z��'x��A�hīpk\:6$�W��L+RC�ɀPj�8b�^"[�2��vg��c�6�=�çP5:�� ��1,4A�"O�n����D���T�E0|�S�<a���o�I�����棊c�n�0�jx"����)�y�HA�X��u�����\�����d7�O� dݑbc�90|8��A .�
ei�"O$}����}����+��?��tS�"O`0����nuRɁ&@�	"����"O^tcA�D+�Ire�h��Y�"O���UlH���<�$�p`�yXR"O��d���L�%�cN��+q"O���r·�+x @�S� �kA�%��"OT����v����r᜔,�	pF"O<�����Fm
t�Ǡ�
,����"O
�
A���PeO�6t\2�"O�P8�#�0l�m�D��`����"O�l�V�8�2���"Ǣn�fԒ�"Od�bQ���3A��A"B�6u$HX�"O"��p�R7.w:�g��*:cޭ�s"O���#U����Y���DD�託"O�i����&7F���.^#4��x˕"O�-���%*�2T��Àp|xe�"Of����P<yI�b̓	A{��Q"O���2���W,�Ej�	
of��3"OTtBa�$4�l�
��=Sd��"O,s��ӗD྅J`A�ZVD�ˑ"OV��R���k^���C�t92�85"Ob�Ƞi	o�abR�B&R���A"Of�z�C��h̠iQc�Β>�A�"O�Kv�Z��Z!��+J6A�ܠ��"O� q׃�j��Xb�����Y�"O\�èӯ)��<
� #F&�"O��zE�^�l�e
� 
\<��W"Ot��e|� ��/�2U�$P'"O:D(���"`$~\��@�&V�Tma�"O.�@K�Va�	CV��3����"O�!�(����b�˭�*Ĺ�"OF��D-[&q*����K��h�"O�E�7-ơ�� ��sq�ي"O��G�
�/����@C(Hx�mSV�\�d���;Tp��5j��	9>H�V�U�����6)u�C�I�d9v0 �	\6�bX�ȊA�bC�I�fQz��w��%�@$k#�H��C�ɞb"NJeE�  �h)#f�ˏ@{�C�<N�ً�$@�X9���?�2C�I�{�<�x�-'6\�����=&O�B�	�E�R�I��m��H4#�B�Ƀw�� *�����8��=\��C��S����&a��� �DJ�W�C�Ɉ\���*�cI�5���lޏ
NxC�I $L�3M�r�(�f�;D"�C�	�0v�� 3�A,x��pQ�9k0B��>#�+��(B����Y�:B�7m�t3��@,{�90��)H!�DC�F�|���tl�=�B
��!�dϩu�t�Y�G�T���xqg�7D�!��/Q�M��x|��a�E�2A!�$�(�H�JVI��^6�@�D}�!��C<Y��Zv`�>)�����)z�!�
�	6(ʗ.�{x��'�v�!�Q�LR8���Bw9bP²�+
�!���L���h*,�r���$M�!�$Я�����f���8p2@�!�dC�_l�I��,1|ѫ@C51�!��/?xe`�c�(g��ˣ��:!�$��<l�ص�F�P���I�АD4!��t�~��b�3[<0,A�̣1#!�$R9N� a��B�B�ZE��L��k!�[�?��4񦥃
WJ� ��S&!!��  ��q��w�D��@�[9Ô��e"O �1�Y�YB��'������"Oʹ��J�o��I�Gќ/[����"O��C��9��$Z�R���jB"Oҕc��ܩw�d��� a�'"O:��ιP�$4��_�xp���q"O&a��Q,di�q
7̑148�'"O��������L�-bfE�D"O�m9 �̈́=���gZ=L��Qۣ"O�q�tDG-;�1�0jF4T� �h�"O�%;w-O�a�^��3�L�4���W"O��{��?	�G�W�,��I"O>� Ӧ+'a*eK5�7���"O�mD�<���x�ā�Z��8�1�	eND���wg ���e� 
,+�ϭ�y�d��M[�H �ꊤl�$�b ��JI����ḧ����l���A�H�qR���Ô��y���T-xr)��uL�dʃ�~��AN�����K������	���'2�4�����(�'�\��f��0�,�J�֤ �8�'MLP9��*�dhŌ�<C	�E���Ğ5,FXL!���N�!�8�j�S���c��a2!���1.t�J�g��K�{֠&H4�2��)}qO?�D�?�T�����q�*TE��!�$ͱ|�]��R:��}�a�� ���7)�,؅�	�=5&�Z�^�B?��F�ׁ�C�	�c� irg��>O�8�FX�K~C�I�V٢x��I��l�p)���[>C�	*X\5�&̓G� 	:T'N(O�6B�I!}܌b$mZX�֑���R>�
B��_Ң��2�K�GK��x�Ł�B䉵R��YkFb��?��zFI��C�	X�����3
�YZ0��
NW�C�I!<&.�*Q��x$䠑�`L�C�	�F�|��u��)[�h�*B�ɓp��e��mH�\��t��c�+�
B�I9zF���oPrRĐ ��'0��C�I�+�H�����n�`���F �C䉪4�<���ɮ7�!�B2I��C�ɉ9O��G@�Nf�u�}�ZC��Vs����՞SR�d@�E]63H�C�	�>͚P{D��Z,p䁇�]��B��K�D)��Ƹ�|���eVBB䉧|3�-	w%	�9l�PF$Z�aNB�	2��$�w(�� �T�ؐG�<ZZB䉓\(��%��&t(�!�e�B�I�}tu�#�b�B��C�/La���ȓ�:����K5m�Y���^|��ȓR`�����V�8�T˰�� �L�ȓt��آFقP�wd��"oU�ȓU[�|"@A�
c@�,����Y�
!����+vp|�)��l���B@ֹ2�	��le�@�Y|�܋c-3D��r�*�����d�-e\��3�1D�`!!�.U��,�7AO�':M1p�/D���uNрg�ԐX�&�3�^�"֌?D��`c��	k��c�D��0l��c;D��*e�UBf�;���-O�*��R�'D� ;u�S�'�f,�
6rf@�HN D�Hz��8hXd�L\ q�H;D� �so:�
��P��kd�E���9D�؊5�R>de����h�����a�6D�(K��Z0u������[�ɨ�"2D�d���J��Y3PH��~��u�l1D�� m("G�"y$��&�VF��2D"O��q�K�D���aԫ�>�4B"O�h袍۠XE21#�$�0A�N���*O2�&ą,��@{�L�a��]	�' \P!�ۦG`�[�(\�\��`��'�:�c& N�C}
��HP��Z�'LUX�߸z�Fu���ÊH��r	�'\��N�F]��S�c�M.��	�'�����W��Љp��O�J��	�'��6.� ~�D��`
�O���'�^=���Pq���To�w ���'c,i�!ܜu���Z�`%V�A��'� ����Pvej���M\8B:���'�*|qvCʭ���ȧ5Z�%��'Zz���ǨY�H���-Y�-R�|��'	�)2wnO7���t�I�T�R���'�P!����9��\��2ՋD�5D���p��G��ْ��شN�%ʢ3D���dF�2WR���L���J6�3D�H��
���@��X�N&
8��.D�T0���e�X��W�Ijē�� D�����3�$i���?��5�=D�4C��ݶZ벐�SMU�L�lx{ 4D�D�#_�s �Iv(ѥs�H@Y�,D��s�Jw�]H7eȓA��
!�*D��xǠ[ ��Q�3��n=��aCA$D���A�n���!�l�#�0�'�"D�4�3%�:�P��H85����)!D�l�����T�	���-*����0�2D�4A���)8���g��~T�t�3D�t:��.4B�b��V.j�J�xV�3D�T� ��?�ld1qAa;��"��*�	1T��T�V���n�8|�d�w�<�`�kS/*�B�Ɍ_�֩�1i$�hІ�<�4��E]
���'x�aD�,O:���*�2n��$a�� ��1�OXu��
C����6BW&?�����
�6����>` pa�ۓ`e�mSE�UO�@Z�c�	LL����?�����̇�b��'쌽mp:����%xe��m�!U��u��'�*�� fז3��p�[�A�BL<yш7@�(
��߄Q��Ҋ�N�օY�L�^�8u��HD�[!򄝤]Rh�2�����A8%��L7�i����* ԭ:�j^�R�0E���|�Gf̌]bƈ�D̸}�Z��Px�C�+�B�D��w�@<&��+HJ�C�ȣ`D 00��D"c�LH�鉽dnJ�{eO@�l^(�0E�����]�z�y��a�,a���t�6'^E�D�5k'�d����$��q���54������^��2��}\浸wL8?��>W��3�o��t�R1����OM�IS�P�t��M�3���O��D
�'1��*��g�6Ii�As��Ӄ)d���9��CѺ���i��b>A&�L1 +Y3����gf��y��x�u� �H)@��.�5�
_�Q`s 6>�RAn9\Lb��%IЄ4�d��Ibg���&Eޮ��L�KM�`���d�7+�x5����_g�(KU@L�1�
��B'\7s}��(2@Y(Ex4��04����B�h�`�1IM:}Pq�3?ٶA4a��\�`b�W�H�Ѓ����OL Ps@,�}z�O����'��h��[�C=F�)�菽:�.�BsmL�yڨ5��D�S��ԃS����O��'z"�P�	�r�jm�����&���B�'�X0�LC�iI��:���aǪ#�'��a�:4�6�*'%ҙ26̚p��p��2Dl00�U��"Bd�TL>}2��G�'��l@@k� M��r�i�=[|e�կ�.�.�0vޘ<��y)0"�u�<9�m�D��q`Ŕ���1��u�ɩx-<�ssD��h�Y��yJ�a� }���#OM�y�j�=X�����O%�vB�I�LG��1
8u(�����'9W��3CD�:�{�"ޠnb�K�2�J�	!��L<D#��P����B�Y��5._��2 �4|1O�� �;36�8��d��9��P8�����R\*�I�S�? �E��(C�'����0~2���,b�@Ώb�qO���F�1�7O�� #
l�N�$eE�$��"O^����>���
AK�:0�.�V�Ի3�"�	F��ܓd� �'c֎܊���55�4�j@I*k��C�	5"�l��e߅=t�#0���&`Z��AFH<1���r���à�E�P��U1�^�<	P�Y#x��ݰ���a�T���Z�<Q"�6kD��L�!�4�+jLI�<�f!rб`#J�<;�hSdD�<!HW�h�+����rB�Z��G�<ig)�$��4��B�:���HEw�<ibds�P����5]����@#�q�<�W����aQ�G�>����E�J�<ᶅ� �6��aÂ�h�E��n�<�"i��]��IS0���$�i�<q�FK�K�ʂ/a���('QR�<ٶ�R�?\�u��ͧ s�!ؓC�N�<a��C�jH�a�!�`�Ny�N�l�<�p� ��1C�� #2P��j�<�vH +���Ku��"ZDd��AOm�<��	<pɘ! ��W�I�=`e�<!ªR!m���@d@FL��H�<QmU���{��əz �m���CJ�<I�풩\i��3c�!cD�q��H�<���S���k��݁=fV����ML�<!�D�:$Vh;t��i�5Ti�E�<a�bT4)j��r��`[�b^�<9B��N�����a��.�@����v�<qR�@-�r��TD6jX��$]l�<�&�\K`X"��`.$x�D��h�<�3�����!� �*"<|��a�<	�����@,2d'�	]y���*�_�<!�l�2��5:4,�|�45x'�T[�<��O���H١ �
�x��-㐏Ml�<�ť��IS�|��K��0<�,��c�m�<�� �
W�$�T*��LaIE�d�<q�d��g�N����@M2��Y�<!��W��k"��DR����,\�<F��!'T!��hȜ���1@�]�<��m'D�UjU�Ņ]����юX_�<Q�o�*VDiË��c�Y�<�����J�ƈ���Gu�D4rE
y�<��H٧O u� *�:��d�E��A�<��®Q�T�"O�{(���d�By�<�΀6,� FB T`�Â�Cl�<A��	U���y1��T���&k�c�<��D�!�x0��2�i�w�f�<!��D�gK��" �*��_�<Y�c�=%\��c�*3jy�g��V�<��!NFb�Q�i+m|J��A�V�<�#�]/*���`�	�F+��1GFI�<)tn�x	c��	�8�C E�<�U�~��I�p�� �Hڕ(�<�W��*&\d}𰭛:.J���d��C�<�R���\��EqPΎ1����j�;�y��:%�52��w\��2��˘�y҉_)^Z�B�,k�ޜ �Z��y�V�XQ��
s�.e4�`ڲ�yн��:�I>vDެ{" Y��y"Z�UIXX�FL�t�m3�.N��y2���lE������w�r$ �K���yr&F�u���4��e����Jʁ�ybe�������bU6�+v��y��I[F,{pdA�L�hFV	�y
� �!��B �T8'�^�N�Ze"O^9W��aedԺ�Hg%p� �"O^6��u����Vh
w�B�ٔ�=D���G���r���*�r�`ъ:D�v�ӢKG�t^jLh���O#��H�')|8��Θ�atJ=ZA)չw�u��'y�a�6�� _5�� c��b�Щ��'�hxȱhT4��APaݣvo��1�'!l11B"�'_@$ 萋Z����'��d�1���h�z�"V�S��Mi�'�Y�C��*k5pT�)&+�I��'=Tkd�;zM�'���C>l���,�a�
X�N��㑪ņ]��ą��z}*U�>��m8,@(�ȅ�*�V�Ta�o��\�#��9�|@��@�4С�ȿq°���V�F�d��:�e�fcR0̸�$�;(���ȓCʁ
!��HHj��Շ2y(b(�ȓ-��8d�K�lA&Hޤxu0��ȓo�����ݙ\�h(蔥�N��K=���Η�x|ԓ�!��h��M�ȓ~$���BA@�5���`	�2��)��C��T�Ӌͽ� YCK�)=�`�ȓ-4X��KW�l��G�4	�p�ȓSs��B�V(kR����׼F��4��dX6u1�)�.g����L���x��x��4;g�` �pA�r�h(�ȓli�-�s�ͣ%2��`
~�|؄ȓnof�y4M�w>���f����\�ȓr �e'X$i<��ꂪ/�U����d� ���R�Y#C�^"?�T�ȓH�)KEE�#v)Hzt��}��h�ȓ3V6� a��p2�(ↈ�5pt��@ª)	t��V�%K'��b��y��Btj0Hƒ6��1w̈~ �ȓ|q
��%��\�`L� XɅ�(���k��,���+�@�Va��<^���晠r�Z�I��H=�Ɇ��t����ψ+h�K6��%���ȓe�h��ĺ,����f�#* ��ȓ
X�
ڹ/e��3Ci�)������LQ�~K25�1����ȓY]�`����p�) �?f�`�ȓiEV�[!��|d&�P��P,�D�ȓd��rB�5 S�R;5Gp��ȓ�b5� �S�����S�?16p�ȓ]Ɋ(��W�TopP��ֽW��؆� c� �!B)|����5A&чȓ=�Xx�'T�=��X	q��60�0��*3fa�@Y�,�j�� [�D$�5��Hl9)�mɣLϦY���/�t��:������Ї`G�m���B�%�
m��*��} c#̔@?fq�r�K	�Մȓ��(��m(�pWaD(a|İ��>8t�)�'Ãuo�}�RH��V��x�ȓpo�`�g��V0�9�\<2�4��J�<��t��C� �i[rYm�ȓrjlp��a�)6��ɈB*�Y����w*�%�g�R;ح�ҋ�F�d�ȓ�~,ˁ�́q�Ȥ�A�ӎZ�0Ąȓb[x<�'�A�b��)6�
[�~	�ȓ ����l�&ת��p���Q�ȓk��a��/�VYh`�C� 8�Ą�ih)�,q�R}���߂`2Ȅ�S�? &ՙ��T5��5㐮[����"O��9Ơ�5�b�R
��(��K�"ODp�@Jю;�d��
���~�
"O�)[�/Z�D��00oߴl�*h�G"O��@���v�U�/ʩBz蘲"O�}9�"*jN���gH�p0"O�)��'H�NŚȨt'¹`"���"O*�{�	K �޸ۅ�D:� �"O� i���'��1RM�u�,-��"Ol��6U>f�d-H��|(�"O����K�B~���g6ڲ�p"O*Q�t
�)g�x-cefY<d/�<�p"O01Q�ơj&��S�<�mA%"O��P�*��p�|����a�0K""O,Ay检׸���Ċe\�q&"O�H9��Q����jQj��"O^�r�,�7�r���Z�E d�A"O&<�&�T��:	���Q"O�0Pό(w�:T�N�=�<b"O4Ѐ.45]��c�+[n��Q#"O�� Y=0"H��L���9+a"O���Ƈ�Ap�Q�lҖ\uny�"O^�3*��kʔ�q�R�!��q6"OdUJpL��8�N(CC�Tܘ{�"OơPCKE3j��CUe��3�"O�����?]m��{��h\ k�"O,݁dm�uC>�*� �&#�4}��"OP�х��bh�Mߦ|բ��"O�U)�K�2�>`�ӬW!Ĥ���"O��!G䌓P��)�R�ݟ|^"��w"OL ����!�p�@ �ܬ\���"O�u:2���tm�Ul�5i>�`qC"Oؙ���g����K�}�b�`"OR��#��;�����~B�mpc"O�u�q��3$��]CBH�d>�"O��@W�A�c�\E1R��X�u��"Oؤ@���Fa =;5D
3@-��"O,9��
}�hɊ��B�J�Rf"O��b��>`�Vds�J-��d"O@ Q�β5���a��=9њ�X6"O&�s�e�:�Yۓ��/vn  p"OI�P䎌/	�4H��R"Oر�-
��bD�2B��`�L�bd"OP���(_� raa��L��H "O.8��\��`��#;/<���"O4���*�f���v�۷
����"O�)�DL;��[(
�G�^5L	!��F3	W���F�,����0�!�Ě?��Y:b�]��� 3̈́�=�!�$�5����M������G�-�!�Ą1+5���	��x�i:A��f{!��ژ���p���r�Nun!�8l��Q��F� ���yE!�81�p�{���5���6,ܛ,:!�d�<j��YvJ�;��%Pa�I�!�D�>G.�y�?�E��"�5�!�$(U�L0��H�A��xqrO��Q�!�$UN���b�9�.4�#�
1�!���,*��!�u��t��#w�!�d��Ⱥt�:Op&8��!�)J�!�䁁+>$��b�kN���文%#!��W�E�x[ ���0�y3I�x'!�G�8��=����x^�bb�W=!��ޛ:���Z6�� Ye�,�bӬ;!!�� �qzc��)p�p�pj��xc"O�m�ʑ�U��PGe�4f
�H�"OT��)��chR$�@�_�"�`�z�"O.�J���(;�0���D��P���"OjzE猢{N��P�CٛϮl�"O�*�fߜt��u�`bF�>���"Očz��̆lX�����|��4Z%"O.�p�IJ-��UY��J�4E�"O(�4�!U��5a�lO�R�z�`""O@)`%��>B�ppsu,^2��}a"Oh��솓8P\��BגVE�<H�"Ov��WԘԳ�&l=�y`q"O&02�Ɉ��6��uÈ�f'H���"O����Ɗ/Fln]H��ȀT�|��"O(�1����H��މ���)�"O���W@�5q���°����49�"O�� �͇��N��403.�ʄ"O8�R��A��Ph��S� ?Zx�"O��b�* �`(�CPr�PK�"O踫�&�G�D,I'�ݱL��@"O`8+w'՗<�D�s].{����"O�u���+hd�}��bU)IR�I�T�<vូ>8]�+]-�0q��Px�<�Va_�F�����ɮ<�xi���b�<qԯ�9��:d �&)�4!��YP�<�[(n��ݓ6"�x~����I�R�<���8���"�ݛ�Z�!�KS�<)��A,0�*� ��LB�X�[�<qU�$��y�%IW�Zv�܃3� |�<�AD1�D��a�@���#�|�<ibײ|���צ�f���g�
d�<q�FI� ��,����Q��%�vÊd�<��BA�Z`��=<{(�B��f�<��GP����@�\�|t��G\�<��J\$�� �n$M\�xV�g�<!��U��"R/�x͙��`�<��e�	{|��u����f�[�<�wG�E���X��ȹF��-���U�<@53�"�Q��5	JNq��MBh�<��)ֿ�p��т�wO�l��F`�<٤�A�8^ɑa��L���PL[�<9���1N���R#�]��4j��JO�<�W�lb�p��I<$�a1jEF�'�غvM��@ �qgE�<#X�����-kH��`Q�J�������� �����=�K��ҥB�d}�<(%�ǥ��!`�?D��j�fӁA�T����� =s�\�p/>D��13�o�}c�i�u������?D��ȑ�2,Z�Yri.}��I�f>D����T�0�~�з���x�b0��f�����Isy�A�}�\Di���)M�~�R��֘'�ўb>��2�@9^]�V�[0Z���AF!�>���:�S�Op�J�LT	�)"%bߴc�ƅ�4T���<I��S /�V-��H�:�Q���0+�Fy��[��ȟ��K߼7�@��P'H�B
��AͱO6=��� ��O��Q��	
�>g�9`#��e��:|� {�'�:���]�h���I�qv�,��$�Aq�e�)f�h,!�́� M4`��,RL5S���I��i�H�m݆}J*�ѐl��(zT}�&�!�S�O�>�BÅU�A�����փc�@D���	��0|��b�k�ؑ�Ulס N��.�^�`Ą�<%>�i��B=��]��*5JN�=���+�U��(O��D�@�Z;5��vk�'�L�ұV��D{J~J�O�TrQ�q�t!+Ҋε���Ad��:lO�P�K+�vT�do[� ��A��"O0sP,�X.�(�~�hU"O� PJ`FH�z�|�k�X�Tg�"�"O��[v���{vF�+R�T.Y�N�*s"O&�J�h�4WS$��gW���̫����y�H���i�^I�D�ߵ��+�v��j܌钨�R�b�8R�2D��`��ԥP���,+H`��b�2D���B�M� ��pvj��H�$c�$#D���Š	F�� L�5|=�L��n#D����V�n��z��&.lt��G5D�X��i�JF����$qP��q�1D�H��a32Qa��	T�<�c�N:D���`C��p@��\�b4�9u�6D�����Tv֞4H��L�(j�』8D�lx�Gûg�P� ��\�Z��D8D������(!�A�V�$%c�n9D��)���d�n	jT�� oְm�A7D��@����f���U,Jr���$;D�\ M�' �}��e�|L |��'D�S�.�j.�%�R�:)p��H$D���C˝]�xM3���ڥ���k!�L�����q/�Ռ�R�O�oZ!�d�J��2&aB6��ei�J#NB!�&���¢C��t�B��L3;]!�dC\�<�ACe�<P���*%�.m!��C�p��I�)R�Qt�=	t�rf!��qp,��r&Kia��&J��v^!��T�ֲ	2�"QV��Q	��[��H�X8h�@�˰�ָ�O�y�	jm<�C�_5�5趀K��y��<#d�2e�?"��;����y�L	�(2�E
��b!A㍗�yn�?�ڝڠb��n���"���yK�t��`��^Mc�+r�A��y�k��b��]�[�Lm�M�J	��y� ٜ?��xC�F��5��eK��ӿ�ybg��i��q�'@�27��Y0B���y�D�j�EX��N�aN�)аI���ybe��%j��a̲\Č��6����y��8;r�{� �� �,s����y�M�1 ����{J�����y�_����K¸m��l���y$��d�^�ĮF�U?~ ��3�yr�	h�`94�=OB�����;�y&��n�HǢE�F���	p/��y�ŚY
T��Ê*:j�Y� L�y�ꑐ~�R�yc,�>4ب��ۥ�y�� {䴂�L��& ha��/X0�yb��]�LI:ah 
1��$�����yr&�u����$�d�!ʃ�yB%%��H��j�ۖ�����yR�F�Vt�HY}5�(����6�yBo8"� �[Do�r �ii.���ybHTxq�f�1cR,���Հ�y+��9�:�Y5'�V$<(`�^��y��KX�;�Ë�{\��Т�̞�y�bW�'S��{T�R9q�z� ����y��ؐm��Y�RkD�k� A�R��y���2R��l� ���uЄT�R����y¡û&�%��iT��He����yB���5R�d@�A ������ت�yrI
=%^���gH�2GB�0�y���K� �ٔdY5�F5��-���yf[(a5��Brf )�V4[��X��y�6E]����5x��ܢ�	Ԧ�yB��6w�yv��#ʠ�@����y
� �hq��͋m�
p���l��"O�d��f��Ti��lX?:�����"OF��K�'�*�P��Ɋ=��)#�"Op=H"!�H���0dئ^�[D"O��2$�ʬr�x ��$L�J4�`"O�觌��%�f��t�˒4�b��"O���@^z$*  ϹJ�h�t"O4	g�Ϳ �t��� ��
v"OD1��/![��S 䗥3
��$"O�Q�D �:P�A�#�
D^����"O|@����\1�B]�8I�%0�"O�=#�k\F�(���" � �a�"O脛@a�n���Pa�g�@T�R"O*��Bwp:8�@�@�>�p��"O֌B�`ċ1$���/�>!�����"O�v��;5v�xoP{���"O�d�O	�5�SI�*�LP"O`���S/�<���i�8	z��"O�X+bIՠ)]R�	%��x��@�p"O�|j���gZ�I�"P@�i��"OX`�A��516кu�A�Q��\At"OL0�EJ�6D�P{���!q��q{4"O�T�2@� @�������"O��3�̌.YL���	��Q��"O*d�M۫?r����G���Y83"O
Lu�޾Z�I@�U�$na�#"O$`�v΁�`˶cn�8b�"O��p�Q#hUB��!�k����"O�%���3���[G�V�Y�zI�A"O8��ƀ�;xdl����[0�v��"OLqÇʙ�Wݒ�cV��;P���"OޠiЧ�ԡ8 :�j�!"Ox��d�*zz�TI�؝dN��["OL$#*X#Iz�vIτ}��"O��IE木<WD�p(ތ@��I9"OԴ0�Ɂ��܊@��)h�"OH�#E`Z����B�U�a��!�c"Oj)��aϑ�>9����o�Re�V"OtH�@"P�t�-��Γ<x�eku"O� �$M!d����Z�m�(�r"O����Y$X�$X���o ����'6�]�w�Ɩ��|QS/K�deQ	�'MLl���<���3 �P2=!�=��'���%ނn��̊���h �z	�'NdX��J1� k����	G� B�	VL|c��ڼ 6ȸu)��[R.B䉪My��KS�K�n�*�;0$B��Ni`�B����f��"\.C�I+�I�D$)�`G�ύ	�B�ɑ �
P�#<ؽ��!n(|B�:d��0�1���db��y`B�ɕ�I*wG�5�h�Qte��4B�I=7P0�දSd���'v�4C�ɴF��J�O�dX��r�Ç?��B�y��)���/a� �CFD�	�B�4(;���%W4Qq���5:��C�ɂ)
���G甕|��@��˙<t-�C�I�C�X;%�k�l���Y�Q�jB�ɲ;���S�eדf���rш�%�RB�ɋh��q����._�Ջլؿ�(B�Ikj�#�I�SYx*ag.u��C�ɌB�^����T��b�`ܳpc�C��jF�(����8�wJ���<D� )p��>5���TC�yaf�Q7�*D�� �U� �$Fr���O9{�(�1"O}���$V�hs,�8#��#�"O����L�8\P�H�@�/b,Z,R"Od+Ʀ�_�])p�H�R����"O[��U��@1T�B�2��v"O�|��ă]������,m(�@e"Ol�+g	�������WJX�"O����Լg���r�jޡV*���"O�@�LRG�8t`Q������"O��K���9n��砘����`#"O���3O>�(ZA �"B�����y��F�{��A0c �v�P���?�yR�45�����j�-r�<4�t�§�yQ�7@�}���5qf`���M�yb�U2�a
�C�0'��k��A��y"k	.l ����/�.�
� C���y"��9h�����+�����yҨˉ�t�B@��:(Z�d1ǁ��y2�91\-�v�S�v|X� �A��y��D�k��;�-_,[IfA8��4�yb�_wF�X�X�vd�`/_�y򭋐, ��d����H`fJ:�y�L�U���L!�L�r�3�y2/��c����Ec�#K@��zՍV��y��>갓TB܏A�T|�� �yBh۹Q�]�� ʋ'�6��%:�y��$>x<� �.Н%՞��b�O	�y���
��(��I_�����qG��y�`nFu�a@<:�ܡIa-��y�.�'.p�&� ��zP��=�y��i ����S-�18W�Q��ybÚ����8c3^9jѠ.�(�'�|4�u�D��NK�FU$�r���y��ɐAd�ڑ�!1���q�ޗ�yb���N��4Q�%'Ȅ�c��ފ�yҥ�#T�$)G'O<	1B,KU6�y���t���U��%� �n�t�ȓ&�h�BiC�VH���M��H�m�ȓk:��I�6�>!b�)�7Nt��r�H� ��U�)�p�.�?`���[⽒��Ɗ")^�c!� �ZI��9���#��V�db�n��.Մ� TB�>O�Vy�fjW<@�f �ȓ L ����/��<r`5 ��ȓ\\�H���
3�| �q�'� �ȓz�Zx)��F�H�
�)1Ŏ�SW�-��I���c�
�'�FM�����>���@F���a��o)E��E��2�湅ȓ0������Z�x���E�!f����ck��2�̈�r�B�G�ۤ?����2�:���|�xqH#�ψe�lч�p4�B5Jj%B@!.^�w5$чȓS�&�h�%H&Ml���d�J�a�(х��6����&N�P%��K��"���C��6c
m�z������ȓ.�z �ҋ�"z���	*f�~�����u���~hJ@��-ʦ
����i'��� .k�U��eޤnj�@�ȓQ7�	�ǌ�0g�����ŉ	���ȓY��q���X�� @ǃ���P�ȓql:���΍~�$Y G�,9�J��ȓQ����/rTUH��*Q�����|�q������B�?s��H��R���2��?B<�C �={B�I��S�? �l� �H6	4����\��$X�"O��Ƀ(`�D<�C���b�D�"O��S&,С[�������J�"OX=	�#h
}��a���L���"O���fM���f����!"O��Ƥ�'a��#'&�)�v��p"O\�1Q6?2n�X7����"O���B�4�1��.)���"O����  
  ��   �  �  �    "*  �1  �:  3A  �G  �M  T  _Z  �`  �f  &m  js  �y  �  4�  w�  ��  ��  @�  ��  ��  :�  ��  A�  ��  �  W�  ��  �  R�  ��  ��  c�   Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�� |d��"O
`�(�;���8���-0��1%"Oj4��ND^[��"3/9�0|H�"OB���H��*�ʞRy=a"O�味V�!X��!&F�:J�$���"O,��a
���C�Ą�M�"O,$3%o�-���p���+Ն�:1"O��ݢ1����`���y14]2��i�<�6��{_���c�H�`�fX�$Kn�<��A̼VI�xR[�)�Ć�pඤ�ȓA5��('nߡ4�� �)˩%� ���,��r�؊b#`T�eT09���ȓ!�b��g��}�8�F��-? �ȓ
K|m�ș�VṔ���2�%�ȓ"R�X�j�4JN�1�˘X�i����̹	_�jZ��1!g��zܶ��ȓgil,*�J�
j�Ne��i�J%b���f	�(U��:���G��$Y^م�~r�� S�%T"���k\�jx�ȓ|4�1�îJb��@ӵ�ݩn�V��/[`�"�v4�R�!ʎ<��M�ȓ`:��z�ؚh�J�Z��$HY:	��H��p�m�C1��!��B:��0��EnjZA V;9����J[
2���	��4'J�EA�IVW&��~�(aZ��ӹ�>� o�Y�|�ȓ�f�A�
Ο7�H��M�$�����mޠP����/���ANXo*�ȓTv�����{ ��-7�*h��I��sB�8�8���3����ȓNe*M�悡;������X�o��!�ȓ'lj�#F�m�+R&;�|��2)n�C��0S4���T:
b���:�0!��e֊��)��ͷV��,�ȓ0�&�8#���� ع�L�����;�P�AFd���,w�6dz���s�<CMJ�(�� 2��3f`2� 0�1D��k�,�!V`��1��:_�
��AE/D����C�qÐ<[��)eî�X�-1D���a��#W`�Z����� .D�dI�j¤E�ɩ�C߃;�(Q�3�+D���k�
��1�`f�<�%5D���u���W�^��2I�:X� �H(1D�ܨ�Ƃ�/�Xm@T�ݎP��V�/D�����[�k���G蛥I7�PJ�-D��p�c90;t�R�X
N�$���9D�8�f�>Wkƙ �gV�$6:���(;D�``�G��\� ��F�R5�p6 8D��2����_Q���%M��X��!D�|gTCu�l���Ϙ^�+�m������ا��}R_.�xr��F:$�����y��g��� �	�;&c*$p���6�y��<#nx�&R��Ԡ{����hO87�=�vDd���E��6�q�"fT�&����ȓM����*<�h�G�~���ȓt(�5��'kg��!��<E8���,�l=�0�H�8|ɢ�JO��!��hO�>k���
O����#�z�T,�0#?�O|�r�����,Բ)ړ	�!%�0|�ȓ?�:�Y ���.RcU�����Ǧ�'������cQ&�8���列L���j��d�<i $;�@%sf
�I��ҀLGG�<� �����_�> ��DK�22S"O���떧$}��cI�+: a0"O>�`r�L:.NI;E&�m&i��"O< �W���9��˓E]���x "O�\�FΝ]w�m��dͼv� <Ju��T����|:��#vbC�,����]*!��V�O~X��P#M�s0�������{�d����eF?7J�h�`W v!�D�#l�e�6O�'V7
ȹ�	��o�!��I7�&�٧	�$"��2g���#�!򄞖k��9n;�� #�ƻz�!�ċm�h��Y�(e�@#�!��-Y\�0��䚥?�P�JQ�� 6���!�O��Q���Yʒ����O:E�^�R�"O(X�e�^*-��tS��VH܁6"Ob�����32���E�JzA�>y�O|c��?�a��w{nY�7 W�
C�P��!!D�Q#JX3C���BG	~1V,��!D����"t��m����w�*D�$ A�r9DX
���[��AB�3D�0��%���<��熣
�µ���2�OX�Ob��1"�~���4�b�"O�Zu�1��B���-�U���'u!�dļ|�RQ�]�����_�V�!�D��i�"}	�K�*��y�-9K�plZz�\8vG@%L2*vϒ�3�4,f�6��hO��/��t'�1:>��
��o�fC䉲a�~���E�o�8أA(8^���.�I16�T`w�*M�֩����B�I$z@�,{g���q}����D�,��O<�=�~Z��U�#~r<'"��.ڼ� j�C�<��O�B�4��_�ڭB���~�'���$��p$��Kqk��E���熌[��|R��!���[�t-�bf��m�sK��yR
^�iKb���K�1�4X#�A=��<	��d@*�bp{�@;V�Y C9�!�${
�e�����"$��k(����yr4O�c��O�]I1HоI�$��ӨE�L��'"O��;0���OT�VIB�H��3%��Pxb�>+�����v�����
�p=I�}R�:pg� ��
��p�ƅCbBȒ�yҮߘXG�D !f֧aGhࣱ`��y"*
�<��W�C9l����6�ynSYǲ��RϚ�B<D;���y���)%��'���8��%�����y�+�J�����"z}���NA��y�G�$x��e04eݠL��z#!���%�ʨ[�I��h��-�V_!�ǽUH�-b���H� h���%_P!��p���C�߇F�xcÂ��-K!��2y (1�peY�o��Q�ѫ^!�DM!] V�cXP�feq���/r�!�d�]<r �ڜ���B.[�67!��Q�O�X�Xrdb깫W�'X�!�߫)�F�a���?dJ�����P�!�d��=%v��f/ֈAN��R ��u�!�ǟn�d��'�ƫ� �S�7�!򄉇ga~��E�#�&�! �p�!�d�Lw6�+"fW��h*T��L�!���4X���d�fJ��!�@�Q�!��%��PZb=>�����+A�!�dU�N\�SC�#v��L��"e�!�dXn�"y���8-g��e"L�R�!��h��5�'ɑ{"h#��ց |!�� Ĺ�k��(�1ᖢ �xA�4"O�X8cd�7x�X�@A;3�>a�"O��*�[�U/���A"O�t�Ɓº�Xi��	��!��"O�H�1A�v� �S�E�G˔�G"O�%z͔=�z�ӵ���a*�X�V"O|͹� �%�̜;�N�-'��	�"O��[�莉�����%G�@8:�"O�ÉA�<��8Y�l@v�:�D"O>@R5IP�A��
�Bb�"O��4,˗s�Ȑ��q��S�"OH��4��)���bi �D��谆"O�#��w��JS�3$��y�@"O�J��O�p��(��}T�"OX!yǆ͛�&�(qG�'i8��"Ol��3�ڊ�� O��l�s�o�<�Bn������b:Dm.5C�I,%5aA�˗M7j��#����!����P��h08L;A�^!W!�AY��E�./�4Bd� r(!���8&P �z&���`�+c$9#!�d�Y8f��Ƃ�v�8��%X�
��Č����7�&H�E1�U��y���3!J��X���4mV�	�`�	"�y҄�X6���DE�-�y�#��y��;�l8�+�$:\Q�� _6�y��\�,H�pi�(��e���G�L�C��U;�A�+ոT�	+��-MՒC�ə#(���"Ȕ&'���K�,_>A�B�	�+)��'ۧ%�d�P� ��B�	�Yj"���-��r"� W�[�7 �B�I�tڠp����6���CN�|�vC�Im�މ����OR�#�+VrC�I�fӈLEMP�	���+%�0B�	��ycG)E
���1tm0B��/\C�mq�蔁.��E�E�=��C� n:��6��9
����t�B�Q�C�	Bv��cG*�64��C	�4I��C�ɺq������rケ�q��`�`C�	�?�V|At�ّssv�ia�Y5g[FC䉘k�|��� ء?!N�Sq�\�D>C�I���Ǥ��GfQ4�͛yeC䉫b������N�R�SQ�ʑGSRB��-~�
a���9��i9b/
�,&B�%>�X}+���'2~M���Ǚƅ<D��@�BŊ@h^���V*�>H[p�%D���,xԠ���/��W�!D��ɶ��K�����o�	B@� D� ��n2UĊ���`�=�;�D;D�`�HV'f�蔁��N�1+~��9D�,���m�HU��/�;U�P]��)7D��9�'_���;e�Ԭ#�(Ѣ��2D�L�0A.����&�Ә8�ijT�$D����-�[~큖��):�h��4D� J���4G�ҙЂ��|b�:�h(D�ĢC��uAn� I��ʥ,ӗ4!�d�&)��c���D��{c,K#'!�DO6;��=q��sC*�HblW3D��$�>+X	RO��9�x���=�yң��2t059ui�#�d�B��yBn�u+T�I�C�.�:Y{�a��y2�\'඼0�.���J��y��T�Jhh�Ù�	׎�H�3�y"�?�Đ�ӄ�.�P ��,�y
� fT��
��:�S��C�pa�"O�� ��+i�l���DB�6�Z���"O�q��1L��vmѲ1Ǆʱ"O �s��߈�f����]�m 6"O
�ۣE�8kz���gN'e�̤��'<2�'j��'���'H��'�r�'pAS�IW5��Z��E�}� ��#�'���'C��'���'
�'���'��)�І#�� ��$B��d�1�'L�'���'k��'��'���'A,�AsP�M��tʁk�40�fe:��'�b�'���'k��'���'�b�'��9pa�U�/�\A*C�ڦQ���!W�'IR�'��'��'�"�'���'GJ�f ��J�2�� U(�q&�'b�':�'��'�r�'_��'��(6�̭�"dbt�s��`J��'\R�'<��'/��'��'�"�'RT���^�o`��:u%�1��̳��'g��'L��'J"�'v�'�r�'ipp��OɢQ�@��DV��e�' b�'�2�'QR�'��'\��'n�Q1��sG�a�*U
S"p���'<��'�b��-6-�O��D�O��$�Od<��/�_/��� ћKZ��'D�O\�$�Of��Oz�d�O����ON��O@�y���*}��i ��W�~�~�Kӎ�O����OJ�D�Ov���O���Oj���O�|�R�N)1`n}�5��7����O�D�O����O����O������I$�����ba���w��E�� r!�7��$�O�S�g~Bm{�Π��� 	��l�$��FdVШ��O@�nZ؟\%�泟�m��?��hCfÎ^ ���"	4�����4�?Itl�;-Z��')����&��B x���W��ڔ)p*0L���T�Fr̓�?�,OD�}�r�B4\h�0\9��9� ��/o[�\o.�vb�t�����y���)N砍C7�W)H���P6���<�$z���TyJ~b"��w��͓ !,M����P���	`KS0B:��̓-�����]��R+��4����Y�)~��@��:��hS@��;�<�N>q�i4�8@�yR�ݨ#� ]ɠ��(jb�cb���O�)�'�ҽi��>A`e��;�c������D
o~��D�6ƺ�i�I���O��������|	Rn˯~�!�Ca�#3\ ���*k��IEy������**݁rI[P_�<��u}Γ[W��.����$����?�'�����x]� �W�D�ڌ���?ܴ�?�� B;��'$��­�,�Ǝ�q�B@$�*����F�d��DoZ�~"�I���}&�,a���@tĢ4 �s���9Ą'D����⇎{�H	�*E�zz�T�%~!f��7�քs����&JT���AW�Æj� ��v�M�nR���b��CB8,-~���c*	��X`UB_�DB�Tb�eJ0>P�2�	�X9�E�dEI. u��CBf ��� �@X�Xz���4F]�mv&(ж���H� ��q$
���R�H��Q�t�n���O���ڑ�'kV4�Co����{��<)�O����2���3�$�R���c� "L1ԝI�-Z�8A�FM&��7��OP��O �i�q�i>�K'�բ1�.q�rd�O�J%߶�M+�OS���'���y��'��h��-w:8jC+D�?U��zd�a�4��On�$N`�\1$��ğ���:厱�G/Ʊ51��͌�2B�"ش�?Q��?�fE�U��T�I��I�~JD��R�݌4<�x�p��)Pk@@�4�?9��S�'<b�'�ɧ5��C�PY
�a���D��w��M��/i04���?��?)����)�Oځ�TL�9XP��Boƈn.�i{vG�5s�4'�@���(�Ij���`@g��!c䂐>��Ư�r��b����ʟ���\ybT�e����_r�f!P���e-��k�On��>���Ol���(*��	�i�4M�P1('K`A8��?q��?*OH])E��jⓂG��|�!%֏zL(pAc�t����4�?y�����?�4_����7��{�I��M^:i#�j%mfӾ�$�O�˓�����d�'��$���M�J��N�XE|�󄩚�dAHO��$�O:�1��O���O&�OR0���b���tlW�S�&@�۴�?��Pd�bC�i?�꧝?!�'J���x*��f�
��8�S�3"ꓻ?�f�<��'��L<	ƥU��fV�zZX����[��6)��\� 6��O����O��	�D�i>�J%$��L)L�4�
�~��&�Mc�JA�?)��?����.���'�V��e]5a�س`��i"�'4�lOK��)rL�ܘΚ�K��I��'��'�fe���&���O�Y3+1�������蜼���_ Fr����O�*]��mן���pyr��~���M��D��
	df`q���=��6m�OJ��,�$�Ol�$�Oʓw
�K�@24�H��aZ"W���b��p��'���'��'��I�{�4�7�Ù5�2��s��W��u3"�ȟ��'.��'�R�@8�X���ta��^��x���O1;����ǂ�9��D�O���O�˓�?)��g��pH����m(ѧ�t�� �Cg����!%R���	ӟ��IiyR��	#���B�i��iI�Y�dD@7h���������I���'���'��L���'M�dJP���9��2#��Dc�oğD��by��I�������k,X�#�YJm`�s��7h��[�T��۟�3!��矤%?I�s�� �|¦oܳ}�e	į�4�����Ä�U�� G��XJ4S�3�(!�|�w�8}��
�Ĝ1pE8C�	>�0	�*&���q%�8;��A̒�H�֬i!hHY���!�B�9
�t�)��˗��1��$l-���-좈P���6����=BB0y���V�H�o��b��d���� ��"����7^9>ع0��\���"#�o�l���/�����F��O�Q9c���	 ���џ��	џ��^wp��'���(�ӢXĪ�BVS޽��P�t@b��ʖ|�bћ���<�lP|:s���BAh�IT*<7�P��#I?
��8��"�T�$؛	�e���G� �,��g����d��S��x�Fd�=풼�n�M.�$�7"o"�'�R��U��(r�����q���'���x=�)�s�^ Q࠴�F�1~�"=�'��a���jw�i�<��v�J�DPM�"���''r�'��m��c���'�4�f�;��5K^([��D�4;��I��v]�P�Ɖ)1�( ��E�'�ʑD�(�`��S-�tmȖn�7V�����:s"�qCrLWU�"����B6�JĔ|�CB6�?q����D3�GC�.����T���{ ����+���x�d[�v^ҩb-�h�����a�' ^�Q�O�N�H��$JD�:!�<;�' �6�6�DЪb�8m�\�	C�D!T S���'n�
<�|��a·x���5�'���'h����ccn��i��@�n�|zwb?p@����]cP�cWRn�'r�U[t�P�@x�(� �k��O%ġ���K�5W~�r��ox����$�P!2��$$~����CْXp�B�<�\C�I%Bi����Kglz`���Tu���z�	y���:;�r�ńg�
�	5=�h�ش�?1�����2b��$�O���72� �%�F�*ˤ�CA�G[�`Z���m��$�1k� 1}�T��|�����#�X��f�L��-�
�;R��>| �H���0O^�������w��+�QQ�LU#̟iB�;7�)��ФWI�B��L�k�(��3�'��O?�D]�V����ֲ7�B��m�%�!���8���A�)Kk����5�P�V������?!�So��:a�}�qBÙ����ğ@�I<�N���$��������I�u���yWG�)-ʩ�t)T�*�Tl1�#�~b+�}�*`�7䆉-�2��1�^��r]��X��o�&^.�ɬ��a��}�t�)>���2X�ʅn���p�]�9�|I�qT.��I����#�ē�?!�����	.ۈ��c�)��v��?|�!���jH,`.ْRh�y���\W�';��'��	�Xy4ݴ:��A$hת|�16 R�Ȣ\��?I��?�!J$�?�����e�-vwz�¥�$�IC�]0�V���B�h��r)�F��Ȼ��W$J�Z��%�o~�p�_����b%��gkP8*T�@+d~]���'��=S�����]�t�2�dJ�x5���-ΥO��7.�ɳ�H��d�H>���QA��7�tu�Jo�!�$?��C@F3���(3�Q�Wg��D}�X����D �M����?Q-��i�+K�`�r�!�I׈hA���U숵f�����O��$�k�DXkw��Vت(�'�哀pD�`��ՓM ;�&ª���<����Idt��@��~ ����0)�����XVxE[U�N9Nyty���/sVQ��"g��O��d�t�SΟӀ�ك@~2�Ȗ.̕i���E ��\�?E���'m����

�vlU�5-Cm����O��F~��`��1m�۟t��f�h��ac2!Y�Դj7�B:�M3e�"bM���'�r�'\�D��V���'�bE�}¶h�E����29&~PB]<|动`�\3>�<��`��BR���; �j(k� �0t�hQ[7�[7s�}BK��$ܐB��[�e�d�$�r�:IQ��A�S�p��	�|�]0	�4�����()���u�\#���p M�<E��
F�Z�f+aI�{W/ˮphN<�ȓ��麄l
f]V�!��W5��LEx��*��|���|�2����2��4��OXT���?���F0?���(���?����?������.�t�
v��i��	
�!Þ���O  ��;^�xb�ե�����W�B����P��69�T��'�K����G�5;Y��2�.V:F|R�5ٟH7}�ǩ"���?&䋡�J�(�8F$�5�2��WW���q؞Ĩ B���భ�@���P!D�(8�;7H��Ge�	d��Hr+_=�HO�=��Ϣ�,�n�: ` Y��ZUG���`'
��I˟���ʟ��&a����	�|ʒ��n|�92��0�*m+�Ș&Xj�0� �Ɇ+���i���%"�Ni���I� �\A�*IRД�B�'Y8h�	E�ۿ6\��J�ӭ#�ň�4�H��W �:b�v�#N>� ���|*�4	b튢a_I�X����C���ȓA�:�M��M�(��'B"Zb���o4�d��V�ν�^�hbe��<Y"�i!�'�N��qez�F���O6˧U��H�AIW�t�-~F(�x����?��?a�`_>�����*W�qs���N`)d�L4b�~�C�dQ�D3���eo��
�oB�U�>��@��^f����� ���sn�_�B��!(^�>q���U�qO<�ʗ�'�F6-N����Id����
�������Ж/��u����s���6��.e�����
i劅�B�?�O��$�|˰��t��I�҉ܬ;���:�3?��9�?�	�l�� �d��rM|��S
��-�f��ȓh:�b�<��:��4m��5��h��¢/)�d=
ơ�-j,�m�ȓ;7� ׈X(I�ʰJ��);+���ȓE� 1�v�ƫ[��@�aY:g�:9�� |�U0tgT
<� �����2"���>a`TӠ�L7D�tq���_'@d�ȓV�܀��J�v%	`d\�T�h�ȓY �ad�_ql�����ZY��~��0�瞚jA6H��c�1�"�ȓ�,�C��<Qb���vÄ8W眬��uҀ�C�̌�r�(��D��O׎}�ȓ!�v��C�+\�2��U�_r�؅�+t-�"ĸSLF�2����@����8��	��̉.�0к�FJZ�
��ȓ%&X|��K�M��2�N�N�*I�ȓAF���ef�@
�!ȁz	�ȓInI�śl��h��&�d�|�ȓv;<��3H�%��a��e��L��ȇȓi|�j��E�I�m�(͎T��l��m���j�B6/^ڙ�g���M`q�ȓvC�;t�%h\�:�c��xE�)�ȓp�U�FMܩ�`1ɣ�Q���}�ȓ:�)i%��<>p�`��׿	b\���
0
�
�ađ��I�0�h�ȓ����#�p��8*rIJ7aԬ�ȓKC�9��C�nQ@m����0'$.}��!��
�.S8&�P`α����'q�"] /tB�XsF��.>�ȓ4�>!���a�pH[��B4��ȓI��}R��͆V�f���g�v��(V53'S�k��{t� �O0Їȓy��ȫ!����m1�-UV�D!�ȓd2,��kB|��ݐ�ȗ�[;�݇ȓw���Q�t�^��U��*�)����6�B�o��:��7��-L�~��4����C�I|�PQ�HT�$29z@��e��#>�%�1j
�|*ga9�j(YtLF�#J���5��Y�<��I{��5���\�aX؉� D�<��$F�kK��"~��
�$e�#?��3B}�<!��m �fOY�KS�ipw�e~Ŏ�tW�Y��	�N���W�+7���F@-�$��DL�b����"�:A5L%�¨� k68���բ���P��.e�I�d���nX,8�*�O��aR� �R�``��l�ϚL󤘟�����&B��4��A�|�j�S�,�ԟ�ܐ,\6H�`-ԧ]��(��"Od(�a�
$i�tPR-E5S<�)�C��Y�A�`GuPɧ�S�*&x�W�w�15Ş�x5�P(7� MH �6�*� 31�N4u��0�޽@�iG�>a��� �:�*��e��e�b�^�_澣<���Jn��f��B�4��'��\�p�Bh�#@����d��r�ǌmX���N�'A*L&�3sl�ڂmN�and}��'eV�Ð�Z!q��� ��Xwo�tQ�O���EfA�`nލ릢��RQ(�{�OWD������9Ǭh3�K��<�B1
�'��a�FR:	�K/<�ʆD߄1i%%�����[�<�ȂL��-�=�N<���k�.���Bn<��%�M4*��c*#��I�B����(�'����B�����S��V�>�b�Dy�F\&$�2�)ƆT�X�؀aa���0<��i\v$�4�K�<�X%"�v���k�̓CZ6Țׅ.
���k����=;�m3�Otx���)����T�!��5�מ�b�ŉT�N�i���>�X��%�4�<0p!��3�z���	�U��XJ�"O�i���[�A�Ь�#� e�&�Ɏ�^�:T�ժ����)� %]&�1�� ���G�5[|�Z&F8Lq�O��� �\�I�9ڰhF0O�윪tC�=~{�ɼ ^r�:S�
;|��)U*��Q�l�3iˁ87�Z�KV6pI�7�(OŻ5�Ŋ�ȱl��#m�5eKh�̥��EUyrF40$V�o�4�R�L��TD�#�'��\��IK"�L�elN�c��8�O>���è<����-��ʧdG�ay�O[���bӾ*�0"&hD`����'FL�Rt��Rv���D]�I��'��y��o ���!�VMZ6c&b(8@ܟ�~���ˆal<�k�^�I0���'�N؟����߷MN0�S�`O��%��a]&neHX���u�����	JR�)��5���� \���[=:y���"�.�'P���>�.�`���,� Ӡ³��2�p�$���� ��p=	�I�N�ʨ������Z82f��c}RN�7܄t�=�O�1��A�:�	5l�\�
���7-�LA�D�%D���Q�L�Ґ�Ԍ�-DF���O���$��yBl�A0�;O�Ԅ��y�O�DI�ě�1azd���X��b@�'�(��d�-$�S���&M\�,/�͸���R�������$7�n�4��8ؠ�1��
C�(-�P�@�	�6�[d�� \��?���R%CY&��4���`��8.�i�ɠ"��y�N�Ys��C�B��MP,c��F�.�p=���R5E��*4C\- *i��n}GG�Ybj �TAێ&�pTHU!���~R�O��I(�R�cW��r#�"f�D ���ȓ+���ӂ���`�;��ݜ2F�����9{�8�y%�O��IR?��8g���W�X;�yg_���� bCڻ28p�p'f���?!r��N�DA�C����/�;E�����O��I�tn JS��A0D��yD8� Џ�< �J�/O�{]L=���:�>��x2`E<����f�$W�n?[�x�B]�-a�9*&�!A0n�ai��'������"b�z��8W&,R!8i�4m�3�N1��d�H�H��a�Av���wg�k��D�����B���~�PP
���5Dmb�`�'w(��d�,V�jACՐn�4� �4U=�M������yҥ�O�Q�SjEK��i�E8�Nxz@�qʑ�d�bV�_,\v!��T1��,jD�g�Q��X!W߂Fd�h��^�.Q�ũ�5�?i�''���I�JõXr�E���'	�rȐ4K*O�Đ�$�5�8HZ�K�����c�i%o������5�d9:�T4h�P��B��
�.Y�5F&|O ��G*��w�L�{�Fßh�� Hƕ��"�읦QLDC���>{H����,�韌��-�_��=��ظX���3�y�J��N/*D:�ӫ`���&�\)�h��R�c�8��{*��8!E�=~8���&<�4k�G�ލ�'$ƭ]�!��U&�b��CV�r�PxV��ဒ>����Hp����	ՄL~�Ci�j��$�9i�GC�1�0� �O1iA$���I�ڍ#�� ��H	&AD�	����̅a�,Щ��Xʠ���)X�]����^���II�6$�`�� xzNxCQ���*`��p��򂪤���bS�NF�S�fª����Og&�!R%[6,������ ���'# ��j�<I@ @�9R�޹��'*̑ LPᦩ1CB�W�FB�~֧�teތ�&���iÆ ̪i
�晤�y�$C�KB|m�0�ΰ(FX������d��!�$��דF: �� ��*�ܔ U�^U�����Ida�n��F^L� ���E�Ԑ#��']�C��=_�DH��*���Ƃ�)fC�;J�B���m�t���x��*C��|w�xQ0oIa�jDÎ&�C䉲#�x� �� *���G�Δ5�C�Iw��0�2"I;��q��?&m�B�	6r|�ɕ�C� u�uLۂ0XC�I1WK(�`a݄?�!��ÒVC��%�,�e�Z�%H~�"�L��ve�B�ɬ�
��.�j�d�k!�=�fB�	`򈉱$ճ�uʠd�-�6B�	.4v,Y�2ZI��y�j��c��C�a��mтܬ<���+rCoz�C�	�4�r����#N��(�G�*@o�B�	�$1��P�LR���C#�͏�B䉠�@����d�Z�HJN	��B��(��A�c�8�j�"C�I}� �F&�xP؜8eg:i�C�I
ֵؠ?��z0��M>B�)� n yC��H�B�@�5om2A2�"O���V���.Z�jFn͢F<V8y�"O&!�FK�:i҅��L�),6@�q"O2,���_�F����3*�H�^eAq"O�ܣ����i|\�;`�Y�N�)�B"OJ�@ J46�$z�G����!"O\��W�60��GZ9~���Jv"OL4z��1�P��e�ی�"O(T�� P�L���C�B%�� +`"O�u�m�7����uY ��y�u"O�d�!]/̞� %_��p��"ORTs&�Ӷ�`�O�x0�"O, ħ߼��!��O_����9!"O*�q�� m���go�� 햹�"O���5L�0i#�0�qɅ �=s�"O��Š�T��U�, ���B�"O�nƺȾ(�5�.a0q�"O�d�꟢����]�2�h�B���yB����d34DʽSPt
�iư�yR'H�Q� ��x_ƴ���_��yR �}3�qS2M�"�p���y��P:��M�`��!�G�y�)E�<%�M(6Lٛ' ������y�e�Sx�f\ �(�9 F��y��;iO�Th'l��L����
�8�y"dO:S�0��d�I���Dc���y��	���D��.D ��R����yr���Wwa+�E´q�������/�y���R:�	�"ܗg�t�V���Py(���j��ÉLȆ\��)�B�<����VG�Uy��� �M�|�<�����I����O�Pp,�#�MI^�<��cH�O�,L���d���A��<�SCЎi+ �ԩK�AS�	���<�s�H5�*�;d6<���#�g�<a@e�@!8E�͌�t�uH��Ce�<�P�hf����X7������u�<�Vk�`��(5�G4�*y�!/H�<1!o�u�<Q�`,Q�F� hG�<�*B���Hp �=fT�c�D�<���/�\s��H�d�t
��E�<��ùfdCr��2�n	:�I@j�<QJ )�r�i5#�(ޮ��fWa�<A+C�[{`�q$.ɕH�p6�H�<@*U�Оyq�^~�ё�/_�<11ʑ�\#�8��d[�%T�\AF��^�<pM� 梕���CU�$�Eh a�<ɖ��%/d��7�X�{�p�V�`�<I�Y+�@b��'��t)"��y��	�w,tS�䊽,���u�X?�y�B�5Xڵ�F���cu˙��yb�]�?����;���L��y��s��ɠ�C�7�!�f����yrI��I�ȤIMx���� ы�yRMO- Y,�J�%|4��k�'�yҮ�7Sx(��koTEѧ��&�y'G%s[��!LKb�Ab�ۼ�y��G�=>p4	�R9�1�F
'�y�琧N�Be(6�0Ms���6�O$�y2%^��ȩ�O�/Dgd襩!�y��B7LO�� � B;�r�� HY��yr�V�m���6'��1w�^�y�J�.���/N��R`�Qh��yb�ɝD3�eK���R�Rl�}�<� ����R������R	d;�q#Q"OF|2w(ѿj�e�g΅>Z5h	q1"O�����̓SZ�آTJ�$�Y2"O�����H�+�`�	���7xZ�{t"OFٸ��  U}l�Y���Ĩ�"O�� ������w��)���:�"O���QiRm�2��.Ϫ#�zDq�"O�ȊW�؈O�.U�	aD$��c"Oh�id�k�-�1+�')1.5�E"O���׬R�_�lEk�b� 9Jt"O�����#,J��:��[���Lˡ"O�HA�s�nkwMV��v,�@"OB� �)
�[�
�3��]�omD���"O��K��ġ+�θ�� 	0[��"OxԸ7�KU�A� �Z+J$�)�"O�i*C��Q�4쒦N�Tӆ	��"O�9z���*+���� �j�DhA"O,)kcg	�\�X��J��>�D�
�'u;q/Aa8�4�Ưy�Tb�'����e-7d���Æ�ǯx�B��'�
mB���d{�d�o �w�Ab�' }3#ت�Z�#�q��@�'��|PvܻV�l2D�:C�8�'��QC��m:@1�t��9�́Y�'�)A��[5�$�P˛01m4<H�'�J@���{�^%#�QVn=��'V�њ �"{�F� CFԻ�����'Ŵ�����=<s�i���ٌT��C�'1�A��3��dB`G3�b|�'a����ש2�({EL��:�����'o��QC��2��x��;�EP�'��4�U��0k���J�
�D=	�'9����X8�� ��ܣ/�<B�'T1��a
l̢K���q"�h�'�1rglT<0�(�b�ܨh�n���'*����mȈqv`�"�F�\�`(
�'�TY����^fXC\.b�|�(	�'���pj� ���0�
2���i�'�n�� /(E{�hd���~$��'xn$jf��@����FeJ��	��'T��ТZ'i�Jm�f�P�*��Y�'�Ja@MG�'������&hpĨ�'/�)�De�%9�xx85�

W�-x�'��Hq���7u,R�J@%Wv�(�'�	
�E+ib���Bʽ���	�'/ȱI�)Kl�(�e�Z?-�8`	�'���c�]d,T��W�Ͷ1�-Ot�=E�$b�l����1�I��V,�璇�yr��=rp��U�Q�/P �#@����y�/�<׌u���1/\�yΛ�y�왳U�rp�T��"s�Uئ�ڃ�y��yG"%�+A��x(��a��y"�A!�0�Ѕtt��ɀ��y���7e֢��c��#��SE�x��'��DX��*���m�Ht���'>�j�,�;v���h���?\d��'�4��o^&Fh�B� 8��8�'���[�
�k�pJPk�*�D��޴�PxB�U�W�RL�$j��b��!Y��yBM�sC��@C�&��g�B��y�"�'����2���GcF��W%�)�(O �BÓs�f�5l�a���)�W�o��\���*��TfJ��vt�UV� ���=�|��w[iɐ ���kܝ��S�? |����W�ዧZ�v|\�B�"O�8�eҢ1��q�� (f�t��"Oh�ҥ��y!XEUeR6(U�qXe"O����Г	���Y�i���@�"O�Qj���U�ɡ#�/lQ\ �v"O�A8r�^+3xp��Լu��xB�"Oh�c&�B%z�z�;��_6,���1G"O�ۇ-��y�ͣ��l��Hs"O�Ӗ����Q�BO�a��"O����bU�V����&2��q�"O��%兞a6�<C�Ã,�S"O$#N��reX�H��C(WS� ��'#��"��9�Q�˩2�FMx�@�VC!�P�$�Ӱ#-e N��W�1�!�d��1ؘQ��f�;���KT�-!�d\9(/꼱s��Y��i�w��jm!򄈋-�V�� �hI��B	u�!�d��SƮeZc���6Ś�rfoژ{�!�䍙<����Ľh��0��Ыg�!��&2���f��1)H̡��C�!��$`�j�)��ں]��� �*�1}!򤇇x��m9�9}�6 ��Ii!�dBg��LcG�m�Aq�����$h��-���D,��W%�6�Ơ#!"O������v� iӔ�λ"��D"Oڴ��)K�o TM(�*B�J�%�g"O���P�T#6���Ȇ��H�D`�"O���2��I��T���d_��S��	j�O~|���ҡ���HH	쒉{��'�p!BIՃ�����D�z`�	?�O��n��<���^r����e�9$�Շ�Q,��5o%l0���˷7�
P��7�"t���F�&N՚Rt��ȓ���Y��X��� +ҍz����xLh�ϚL�r`���B8-�ȓ̹÷��;k�,��Q�A-�0���>���@��R$ؑk�'{�<H��'�+O�5ʚ��+G"QC����V-�i@4͞�S�By� �7��iEx��'g���T�r1�}a�C�.8?<�Z
�'*���H,;M~�#!o�#bqr	���hO?]a	�%f� ���]���.APp�����ԏG~�֙����/ e�����cQ�ؠ}�J1�g�߮����ȓTcƸ[��+@�  P��6b�8�ȓ&D �X�N�3�Z, *�3MǶ���*����L�a���M� �Zi�ȓ,�b�aC!&���V�(V��x�4��Ӂb�,p
�e�����ȓ(����A'ݨ@j��	Wl�6>�Є�ȓ��<#�B�(��1A"Ӫ(�|�ȓv�1�$H@@��ĩŢ&{jԄ�B<��{��=q�])���E?�E��J�$�cW�Ɩ}B���2$U>˂��ȓ8�i�%���-��E ׀ӧK#1�ȓStv��C��u�����85|l��E�@3񋆈g�^ a��3q?XM��P� �aj�2!p�0�.R�O>1�����(�.�R�hqL9O�%�ȓx������{� u��R9j��L���x����=H>
�;5L�6S"��� ���2q,�gx&�CM�'�)��U���!�d���U�[�c\T���^MB�(��URi�V��],z���S�? d �c2�̍@7��ؘYB"O���/<�� �~�q�"Ox4)��K-; ���7üS�r�е"OL�b ]n̜A�L�&󠅋T"O>xC�D38Y�Rָ?{F��"O�s���6W�K�0Ҋ��,.�y��F��p(1�L�<��u8�y�Rfu����i��伪)\8�ya�#��A��\��T�rF!��y�]��"EE���K�Q��y���ш�:$Q�3�]�dB4�y"��e�b�B��w�e��#���y��@7P�([�	ƺs[Yj����yR+��&]�	�3␉  U�g#��y2(�8�V94�H	�jA9PM��y2b�e}�5�B�.|�x"M��y"���N�Ti����>ZpD�q�P��y2B�
.\�(��6���1�4�y�$M�"�fLH�O�aI�C����yR��(E\N�`dP2B)�xq���yC�\��	��:9�=C.��y�Γ/.(���癵D�a�̐��y�b��UE���*#tV�̓�U��y2,_�W����N�k܈ �r(ݏ�yb�
"�����0[�x�yR!��y��\�8�4�3�f<b
5�v않�yB	ʨWΙY2&R#I�Jp�����yB��+t0���l�I*�q v��y�R���+ �ݲD.�A���y�M�-i��]�W���g�}��.�y��50hm�3G��Q��)i�܀�y�H�%�"��c�Bf\U��Q.�y2�c�i	
#�| 4&Q5jId��ȓ"D��$$��p��Ԯ�x��t�씋f`��b��hlt��ȓ.����e`Ɍb��+A�X	�ȓ\Z$�{ �S:�2�jZ�U>ڀ�ȓ5 ���B�H�k�����F��ȓa�d����;�8��􆈱9�>	�ȓ 0�r��|�t(� \1q�b��<���V��ga�1@�S�@���q�L1#@��
:��l���K,.pʜ�ȓh�LJ0@�aG��kv
���ȓ|kT=�W���]�p
#*��w�TQ��5�b��b��K0@3����͆�R1hm؂��|���ٖ?C�P�ȓ_I�Y���oT�d��mV�LD}�ȓX����WS�$�:1C�8K�x%�ȓ],��P&�)*��y��Ý�Y�d��P�i��5N+�@�B$W�*B��"�ژj`d2tlP�W�ҡB����%���KRK+n�Tp�EJ�WU�ȓn� ��^�!a	��z�`�ȓM�~��p�U�M������:�݄�w!�**� <N6��E�k�@H��<���*k[�7W��h�.$��=��$єd�C��
bM��x@'ίh�~P��
��A%	�	:�` )V(
*M�ȓ0<�� ����Xh��R�8�LĆȓA�p����2m�P\�f���P��]��G_  �ӠǗl�`�Z��&��T��*��P�7fS�%���;d�;@�����T�u ��y��(SF��5���ȓ���BU&�Y�t�*���I����S�? �,U��	0fH����'V��X�"O�4��CY�|��F�ӕ	�]�"O����Q

'
�| ��+�"O�<0��2$n�E��jB�v�6!RP"O*��w٭N~T��ѮBm��t"O��D��sE� [���2`�"���"O,)!eh�S�@iٵ��?����W"OF����,E�qCJ�9D��3�<��ȓ}T�i�V"2�SiUj>q�ȓv��!3�%�]64�Тi�&�ȓh(�Ei�
�ڐ5�Q��rέ��x\nm!k�+o p�GJ�n:�ȓxN��D��'+i�"�QXd��'_��4�4>��Q����t{�Q�ȓV�(�9��NH!��E@�<;p��ȓ?U��I�&\��+��(2�Єȓ� -'��X���A�b�l�ȓQ
�+d�վ/aq�G��6|��@�ȓ�C2��75��p�t�B/:N
=��X	�1"��ʽ74��R!.' ���ȓ>NxRl#Y�q�&_�8l��C��p�Jk�f́����p��ȓ���v�a?��A@��H���ȓ<1Z�K��Z�k�b�K�<z4�ȓ�`Pd��*: �3��!��@"g\`���(���f.\��!�D��I\4
�À�S tx�f�4X�!�$
*{8T}�P�\-��|[�o]�Fs!�� ����n�+���᦯Jb!�V�:�� C��92�j����~J!�dK
sH.(ɇjJ�ˬ)�3M5?/!�w��e�2&�g�
Mq��ö}!�ýdԪ��U�ً=0��I�	e�!�#O�\����P�HȾ�X��7�!��yZ4%c�� +>��-�'��<�!�ǵ^�>\%a�,��Q
B�"R�!��5S�$��D+ǻ4��+`�6�!�d�W��R��+7�p�ѧ L�!R!�dς&�@��q�S2B�*��6M�[f!��ߊN�"D�wF�'pnm"��ZP!�$A�7��2�ɕC�dYF��7F!�D?e�$�d@v��5�r��)!�Ă�-��,8$��zV�X�K!�J�j^N����H{L�`$⛅VY!�$Ov�,�Vo��	���F,�!�D@�=��YC&2Kc�Y���
�!�O'e@e$V	&fԼ�!���
�L!�ϓ:)ST���%��|�!�d�OuN\J��7E���ۋ�!�D�$~�ݢu�X/x��p��L�]!�d�-7�(GC�q{h�z��%FS!�R�L{@���0B�<��N��Z!�d��j���D�
����R�B�!�dL�U�v���6b�ta��*�!�� ���FO:l��h ��/�!��R�K�ő�`��V�$ ����	/�!�ϣv�}���R9��"s��L-!��{P0����WX**��ĳ":!�D�cŚ�eK]�>�b�k���2D.!��)l,�gGA�C�����$;!�
�L�3C�J2�Tqh�![wk!�$6��e��p�6 �0b���!�$Ǫ!M���dG�+G�ȍ2���,�!򄊗
s��m����
�.t!�� r�	2��@F��6�G�I�a��"O�!!�@M|��GJ��%�h�X"O`H�g_�x���i���x�F�z�"O�L�fZP��ǋ�<��lQ4"O��X BM& ݨM�I� �z,:"Of9��	BJĥ��_6���I�"Oj!��Ս 66�+dg��kD�j@"O�C���@�Q���@&p>Щe"O|$9w㉹&�
�R�냊��y�u"O�(7f׫	�1��BwϨ4�v"O�K�J<��=b"���[�|y�"Ol@��	2z��;�L\�~|m�d"O�`��k�$�m��!��"O���F!נt��4`��'�(�B�"O������e5���$�-W�j�31"Ofy����9���@-G|��9�2"O���n'aC�m����]�qJ""O��BJM�DEt(��Y*`�	�"O��X��5%�ذ������b"Of<j�yD�<���"����"Oz��&�Ʒjp�(V�[%q��)`"O2]���T%#S�|RC�� Q�"O�U����4G�&��bE�� -�x2�"O����T8WJ�H2�пHRK""O�4�q�>-ziJ�đ�b18�r�"O4$���_���Rw�?P�p�#�"O�y	7��*+1d��]h�6���"O��;ō�j>�I��
I?�P�K�"O��pWG �.\KӉȈh���&"O�����@�����>|f$\� "Ob��",9���i� 7`�*s"O�l8�k�0�Tlz�1'9��P#"O����M�3.R��"�^�fT�p"O\� gL�Rؘ_&��'�}s!�$[�:��4á�	�\��*��V�[`!��X�U�)���/<:��$͠R]!�D�5V}:�!��=�L*�(G�CB!���n.�p��G4N|V�ç�
,!��~��
!Яaj�D�� �8�!�D@�M����I�%S���&&�!�d
�a�ug�2�v��ԃ�3j�!�$?�
m�E�V�J��ep�#���!�I���2���(V(
��f��0}z!���B�ny� ;}�t��A��gf!�߻]i84y� �H	�M8���PX!���#B^��$MR�_����re��!��)a��R+�<<���S���0_!��
͞��TICBx���ՁO�"G!�DV9Tp�)�� �@�A�B!��+g~*Ł��:u�5��T!��U�k>�2�HZ<!�&H�Ei�!��1�P!)E�-��RC	�+�!��Q+.�B����ś�4삕�
�!��.ph(�p��,�Е�"X!�����WJ��*�,�D�P�+U!�D+Enp�R��
��!��UX!��U
��9A��\���픎Y!��=��۳%I$TP@T�-{_!��42��Ӥe�/S�V�KPa��qT!�Z�/�� XV�|s��	�)0@!�D�1?"�r��Q�qi�iA%	U�Y�!��0�>��҈�:sC���'�j!�DFd-��kW�]>;¨"%��&DR!�䊏W����@�Cmh(�焼FK!�� ,AAJA-���H��XVL[�"O^l�!�+��Żv��CP"O��i�m	$�m#�L��9oDD��"OFs�MսG��#�Aђ$S��iA"O�h{ ��.h��k�i%m,�E! "O��c��/j�k�(�<^�(z�"O�5򦅃�+*��T"Ù-a��A"Ov�K�&��R�����>w{�0�"O����"�UKn]��A��^��B�"OTy�g�	��ԩ��		i�$�%"OP��f�ӕk��p")S K�X�!b"O�-�$(T�tc��P�0�"O<1˔�ԪnLde�3�M�@���:d"O�X��ٛ�\l�c���,w�Y��"O� K�$��\0QË��2��Ljp"O�Qb��VF1�E?��y��"O�8��Ǆd{��)����?e�%��"O�ݑE]*0jB�����ԕ�"O���aSΈ[Q#��<��3p"O@�i
�+q�pa�h�Ȥ�"OP��!^*��ƭڋpe@1cc"O�\�+У�J���-T�UKc"O&��reZU����E�S;Z1
�"Ot�xlA�}��a�n_$(S� h7"Oؐ�V�V5'@�%�S�4I�ȧ"O���NY�����YveD��p"OR�9G/�G#�qQ���TU��"O4-�/Ӓ���r�RM����"O�)pgFK�WI1�f��a�M�"O���'�;c�� �����%"O��!��݇Pf�[�	�bY���"O����ͩ`P�s �M0[N��1V"O�(Z�k��j�B0J�gk(ys"O���EA��Rᾘ�w��~a:"O��
�Ḧq��J�'/\D���"O�]��!Z���!��E�3��|#"OPT
N<aR�HTa�)�Ԁ�"O�����ښO�D�;A�Y w��$s"O �{��F�8�f�C#^T �!"O,����o*�z�j�`K�J!�$Y<q�r%�r+�S��D�2	ɪzh!�Z��$��"V ; �:�F��`]!�$�'n��JsP�5%��J���J%!�$�*w�l3��I5#���q�!�$.\r|`K������A��!����̹��6jo8E�2
W	N!�!��t��"8{��qcK�RJ!��H���L�B��3p4P$��-P0!��Y	�=H�x�4��5�V�P#!��7��y"�A�(<6%�¤W�@!�dZ�a��IFBd>8����2I!��-��	���7 d8�%����!�Dϱ�x�W%F��l��f�Hq�!�d>w\�Mya١|䀨�A�Nk�!�d:��iXdZ�$�:4���F�4�!��4 V��%-!E��� 敚�!���JY���ܯhT���E�ծD�!�س{mT�!����ab���QB�8B!�dG|�v�����\KVH�e�$O?!�Dک&�:'�Hw�NE����R!�A�^���#��WA��J�G��;!���Y$�	�B
�9,�����r�!�і ��8`ULB#[(0 �"�̽I�!�d\^�j��؝6`S����!�� ��8h��R_��hf�Sn�̂�"O�pr�i����1���!�:Yx'"Oh�6֎Qm��Pg�C�U��4��"OB�iUB�1g��3 V�AA6ew"O��k��ќ�(�p	#4΢�@�"O��2�+��W��ay�J�
c��p"O���EՖ�(Pҫ��t�� �"O4�k��F��y"+&AZ:=��"O�pi�R30��kN�ND���"O�dJ����|��K�1k1b<��"O�p��h�x�.��)L�^�6�!�"O�������҄�]�D���E���yҥ�5�Є8���������y2HO�[��0rb	�|�4��y�O	�H���h�Hm�0� �P6�y�fJ%41��!�`k�I�yba�$ �9


��!b K��y��R�m�=���&F�z��<�y�o��X�!���y{�0���yb���f����@��`�mѿ�yrlW=<�1��I@����	_��y��^�^�н�dʋ4x���׃�5�y�5(�܈@�(�ix����ybN�V���� �K�*}Y�(�(�yrgP�#|�( /f6�X�d,�%�y�`΢�D[̓b��t#�kɥ�yr�]�C߸S���V��!�y���	D%����NA�!�E�ǒ�y��ݎq��Y#�̹2�1)Fo���yrF{0����9q�:��UK�	�yB���L�䠁Q	id��+U➥�y�҂ �P�E�ڮZ�h�`QBC�y��߰	p��`c���!�8ZU!�G�k���9R�ǋ_D|���m��f!��1dX%sA-��\KT��q��M!��Dp����;>�*t *!�d�;+N@�g�P!L�{ga��\!�Ă'i�t���^49��zQ�ͯC�!�DĝM�2�rӧ�+G2�s5��^�!��"_~	��kI�e񎴬`����'�����F\�l�(���K��5�P	Z�'1��2�m�&,%��xr�=1�a�
�'Q��s5��5�N�:��۬X.r8Z
�'#��J � &>p�p���W��8�	�'��	�@��|w�@O-��J	�'��8�����	C�hzՄK�?Ɉ���'���[�H	y�=��(�:J&Q��'��Y�䜝an�k�l[�.�J�'2&��B�BN\1����1�l-��'�:�#j�P���!���L�	�'�YȤ� 2A!L93�hG6>9C	�'dpj&�M��A�I+{3����'��@�#eى+XnкG��%��}[�',@����"��q�8f���	�'C�ʰ&Lnit��%�I�Ƽ	�'��āg���q;B4�s�]o�$i�'���P'u�F���*��`?Fĩ�'����g	�H�؉94�H'`>�0K
�'O�e��ޔ_�E�6�ޫDPĔ�	�'��p����&��Z���Y$)	�'��a�+�J[�ì/�|x�Ф/D�TYb��!��:ѫ�X�!4�-D�d�`�D3�bTsq@لy�rEh�`+D������
Ym����VO�0s�f)D�� ����?6~*�r��S6X��X!"O<�9J%vq��)��}�c'"O@śf�� �lp�e��خ�g"O���G�7s��-83���>Y$�z&"O��P*]��(�B�
!U��"O�(R�`�Y�@XSaˎ1=��9r"O�T�^2,8�����k"��3R"Oԥh2��.ɮ��t@�U�,c�"Ov	Qwn
0'�}C`(�)J��a"O�Px0
�)55�%X�m�65�� q�"O�`3�@�.K�%��W�oN�r&"O<��`�:�����^�OGf e"O>��tF�.F($\ �㐚KT�6"O.QA�#�;[��5x�"R+`�dS"O���Th`��pY"O��*��l�Թ��fQ!Dڞ8"Op!KƗ�I���q��,F��a�"O�A����D�q�Ճ�}��
q"O`�a/ڸ����(J(ʢm�"O����L�2]�E(R���$9�"O~�Y����-�#$��,Zc"Oh0ㅁê/#>�K�K�!5H��i0"Oؓ��)]�b#L�/^���U"O@��@�� �EdM~�t�9�"O8<D�%8�I��"���	$"O(Y˶�C�J�x����Hz�Yw"O���c,�!M @�*P.U>��"Oy��I� O�
��[3 .)�E"O��£�߬G�a��)&lXC"O��Tɞ�;L��Rd�M�B�ʄ"O�@5fW�i(�t�e��4YB��U"OB�ǤN(T����.@lṖ"O��p�i�3������ �F���8G"O��b�U벹�(Z�w��b�"O�a���q��<ہQ�j��W"Or1R���T�@򠀗&���� "O�H���F����o4�.�a�"O����T`�҃?�j��"O�x��
��D�;CN*�<�S"O��`A�J3���Q
Q6_��0�"O�����?/Zڴsw<3
�"�"OZD�r,DMZ�,� B=x�"s"O�t�<f#B	yF&�9�4��4"O�������*�C��6N�l�#1"O�@["A4xe�%2��Q6i��	�"OH�K���7S�h�2�ɫKUĜ�A"Op��a	4~��5�3c��"��0G"OZ�˂"R�i%�ٓT��B�
\��"Of8�q���d�f�!CFt�b"Oh�WDՊ:0�a�m��O8���7"Ob���@̭m��Ih3,J�9�8[g"Ofh�W�"Y�>�(�k�9,�e�`"Ojш�B�*r�H{C��O�R,Q�"O�����{�
��U��]����e"O0�q'0h��H�
��
�,�`�"Oh�(�J>I�����6�4���"OF$ tH�i�����FH)�j`�B"ORe��!I*H"T�X�&�����c�"O�����s�	Qٴ$PƬ�2"Op8��'	"m��L�e���+<��b"O�$��� 	��I���X���3%"O0�bf��5���J�f�|���"O�<k���)��,+���(	�"Ov@� "M�M�X@��#d��b&"O� 
�ǭ�(�����ŗ.U �"O��16��Q7ny"�Q�;�n,V"O~����6�:�єn��J���ȇ"O����`�4)�G�S>b0}�7"O,��`%T�R��6��Fh!� "O�YS!�	M�� 8"`�5h_lK�"Ovɨ��WKD���DSlD �"Ol�����}':�!H�>85	��"O�+��Ί��YC"RL5��(�"O8 9��� ^�F���M����"OHQ:$��O��M����R=L��4"O��a��ʖT�� ��ヤ"��T��"Oހ� L�[ƤB��O��0 2�"O�Q�p��9U�*��L �w����"Od�!ǅ�Z�F
�ƚ:'9��;�"OR�����P���s��މUKv�1P"Or�hRE�)h׆ۖː8&1�xQW"OR��W��=<�9�Rjۀ���"O<�J��E���@���Q�. `�"OZ��U� *1,�0�3+��4җ"O� ��fH�(�x�CHB�A�L��"O�Q��/�$NŨM�C�G�2Ub6"O���Z~�QFf+��9K�"O԰��ʌ�oa���/��	�J��"O0m�&ٙ��ؓ����2"O�z�M�lt��'h�%J$BMӦ"O��bG+��f����R�Q""%+�"OJ��G��/�"�Hӹ��"O���2�ЧdYt���-o�v�X�"O	��o	�e�l!��D�&��lBr"Ofiy5M�(�f��$G�J�D�k$"O0���h�]"�D͆A��<j&"O�x�V쀳#�LQ;3A�0hԠ�k�"OHX���k�X��A�A�h�n�	c"O 8!b�{���Z��8N�p���"O�`�4ƉK�8pH� ֶ~fHD#�"O���$&�+kx���V��FS0Ŋ�"O"eIt�YЋ���9B�e��"O m��垩w�8�KS;�@�B�"O�yPs��y��U�c+�H��1Iw"O� ��F4\*a�=+�lsp"O$��NS�rZ�4��&��:��T3�"OْՂ@�Yb���W|���"O~����:SJ�qĥȱ/|b��D"O�x*r	fD�[tF�Pl��"O>d#�H�Y�D�3F�>��	0�"O^D�ʜ���@�dʧ�p�q"O�њ@���}K8�#`�6�5Q"O�AQw)�{�ꡫ#��
�X��"O pc���&W܍*bcУg��`�"O�L�1�ׄ5����_����	��yB�Ǣ1`��,�Z	�����y�,��|�Z=3e��g{�-��]�yBAЮz�Hx�o�,g��I�����y�����7 F;Z�f�����yr��E0h!c��`�"����1�yb���­͡� ��!C2z�H	��'��@���	�H�"e�!�ټFQڹ��'X4(�f�i)f`J�KįL���'L�4ȰA͋H��D��n�D���H�'� �����ع���(I��
�'0m�Ը{���4��-�	�	�'|"����ƐE�-�̜1����	�'�Ũß�(�:EC4�2*bԜ���� L48�ʛ�epR\��Đ�VA�`�"O>(��l�-Nl}Z#)���`"O~% ��A�.�0�x �^�Z��A"O�9��`�1��
��Q��r9�"O� ����_�A1&ޫX���8@"O��¶��)ޒ����(s�kC"Oxm�ӁH�M5F��L	n���!�"O��uk�6�B�����=�zia5"O��SL�4R�*<0�)�gx�"O�ٳe�#{\�ئڱ Ը�v"O��Ң$�m<� W��n�"O�؃"�.#�4,�Ц؋Y24��T"O�h��a��P%!���K$L���"O���W@�Y�Np(q�_){J=�r"Oj�JG'Y�]!2�
��"OVh�T��om�E��"�!)�}�"O��2D	J2m��4{���	{�930"O���G�$�v�(���<>n<��"O`QՉ�=hpvı��P(i �p�"O���ESB�f�PS����YR"O`l��*4R&����g�Xr�$"O���T�U67��p�8Z��!�"O2h��F۞U��YS'a�=KL"�:2"O�f��t�]i�ëj���"Ov��k�%z7D�1b3���7"O���s�I4.BZYy�m҇Z�4�x�"O@(�Q�
2h�a𫌟tŌ��"O�����B���{�+6m�NHsC"O�<����#ծ�xv*��[}T�F"O��-��m��<Av�'g���@�"O~��էȟ��cW)��Rz��:3"O�[`�B�}���0�mX�I`��&"OR�z6�E1��ʜ�iF�p(�"O8����12��2�.�
qJV���"OTȈBD����U�R �
[-�9[Q"O�1�F"�'4�\pҏ�/9�ty"O@��&�O��jb�P4:*V�"O�!����-;�����+
�&"��T"O<�j�
"+Φa�	��j��8�"O�u��(E
ph��T�؈z���jf"O���g�.���ǧX�(;&"OZ���h��Er�Ȑ-���x�`"OD����мnx�V��yή�2"OD)aFG�i�X5�AM��o����"O@�@�����(�6�bh!"O~a tō�
�B���-U�J��b"Or\	���~L^�r����0H�"O� ��B�a���A
-��Jw"O\��b��D��YKP�S3F�>��"O-z`K+4���)��ԫ<�Q �"O>icπ�lOI��N�9�bLBF"ON4P�Q)��x���	�X��B"O�8��q1T����˷̠0��"O���g(P77޶�zE��=�>�`�"O e3-g�X�҅:A�= "Ol���½cZ�˦��V@�1"O�}��`�#x�:}��i�rUP2"O*�`bD�HҨA�1���c��l�"O�A�@��A�4�����H{0k�"O�u �(K�f0,�R�g��Dp�%X�"O^e9RlX t��4�R	@ibhr�"O����w E����n��"O���琉{��\�Q��L�vթ�"Ot,{����4�@�{��]�d"O� �����=�����y~~ܒ�"Ojq�ܘX9j%��A�wydJ"OYA��$a����Xi��e"O�{)݀|}�� �?U���ز"O8�c����+�C#?�$�(e"OVT�a&�	~7,@Ӧ��,K<��چ"O�+�e�,U�ժ .��"Oz��C�/V6 �Z .�R0�q"O<TȒT:Y�ZU+Ya%�{u"O�P�_���U�T*V2q�3U"O���
��fTr��5Jɖ=ʆ�y�"O�TÖ��5n����HU=-�6u5"O���V@�0Rs�D���a�D a"O����f��^d�&�TF��"OZQf��/j\#_�;&L��"OF�C��3$Y���n� MJ"O�*gC�	�����A�6] �Y�"Oz)`��%S�����\�FN�j�"O,�Y���6��,����!TG`�&"O�lH5�&*�<���|a�z�"O��6W�6Py����vy�"O�$P�*�x���`�сXɸu"O���a�N=u!�H+2��=.��RE"O����"҆tA^pa�
,�)HU"O��C5�?hL1�Wb1�%p�"O���u�D�c�D�C�̹qP�a"O���3i��t^�t�ˋ�=��T��"O�!�_$(J�`BDj9��yA"O �'m˿9��R�IPO��1�'"OV	R�]?b��	qB���J&z�z�"O�� �/պ3��L�
��C�*OQ�����_<�T���ԍip���'Иa�u��A|E�d�J�\{�9��'�q�#�Q���¤�ʾ����'4�	���C��ذ�l��t��ł�'2z���	�6�
!���էs&�$A�'ƒ�xc*L�ti.�`3f�����'ٲ8�R�mߞI�r�%fUq�'��}c�@ < b(�j� Q���'Z������w�6�D���@�'P� 2�ħ]�f8Q��!7��t)�'�lCT.�[(�,��&H�zԴ�q	�'J�1R��8}�h�Pd 	Ҙ�{	�'F ���,�nz��gT,n�����'�V�`-U�xh`��qB�o� -�'O����4]Y�,�䊇g \	�'���Jqf��:��oY�OM�I�	�'���C3`��9ԩQ!朘r����'���d"I�TP��aX����'8�u+d'vr�ŉ���_�<P��'~�1�G�$ˎѠk�S�T��'�"���H��OI���M_K<�#�'�DL[e)V C��
��RB4��'�x��i�.:�4��dPR���'��
���2 1`���A��pZ�'p(a���F��2-��?D��'���;q��K����b'ΠH�P�	�'�ix4�h&e���K�O�>���'DA�pf�(P�>��Q�8Hj�H��'�j�Z₞0�����D�?�2�j�'��Bt���E�|q��l�9�.5��'��d�A@�k<�ȋ�N� 6��͘
�'�ri1/Ұ�f!�L�C7ؚ	�'6��[�D�/�&h�����R���	��� �Ub=t����cZ�6�>�Q#"O�T��G��|�`��!�vq��A�"O���T�I%7�
,ҳ�U/M2x��"O�ň`��)���{QA��Q1zT"OR�+�욺	{8�+G�Q� <��#"O4q���]bxt�Qay^�m��"O"�"�
A�(��5�E�0[V�)�"O�%)ه�r`�#��BLX�v"O�(�@MJ9f2<�1#��HӬ��"O��0��H��kF?ѐURT"O�i8����z&��Z�h�ڰ�Z�<a�m�)��BƢ�H���Z`V�<Q���8�q㖅I��$�#I�Z�<	Rf�f$�qؙxT$P�	WU�<��%��U"���J��4�h!�T�<y'\�yl�LI%m~���C�y�<�Gņ�M���v�^�T�z �c+a�<�G��t=���]5���)5��[�<��E0v������;�|����l�<ɴc�=Zkp �2��4S��@�@i�<ye��63����P�0=~� ��@{�<1v�U�|y8p��B �V��\�C�_v�<��/�13�h�3�'$Ϛ�P�Ȟq�<Yv!	�m�61z�m�7���)�x�<��D�̨�����WS�M9̍j�<	pN�)��1���Ƅ:�v���Aa�<������(C��G� ���(r��]�<�'�Xa�[#�=c������Z�<)��վ*nv��1oٟD�̒vBW�<QSMY:i���'AP���gEV�<Y�`ϒ8W�ΛQ�u;THR�<�@�Tq!z�h�� J%���P�<�����ET�����3�XI��KD�<	��Q	3��Q��
�F����f)MC�<1��� "�.	��E�c�DY���Q|�<1��9_�
٣��b_rU"���t�<�Q� �����yiĬ8��^p�<��KJ��\�㚀?3�Xh�Yl�<��Æe��lX�A�Mz=��A�d�<�� �p8�AX�\�a9���ȓ#X�A�+>���J��R�
��ȓq�Z��%��=)�ir�ܑ)Üن�f���s����
4h��4dx�ȓ$̔�0t뇴Ni�}0r�N8 ��ȓZ�8�
cC$(8�/,T����ȓJ��d�7@�xO�c0�(q��A��m�2�
�K�4;�yud����ȓ{�Ra ��i�6L�RI�<$�|��ȓ��M�ehK�y��q�<� ��1L>�c���2uر��`�z��ȓV}�)aeP���	2�y�ȓt�%��Y:kÀ���@�� �䁅ȓڜ˅�� _x�"p#D9u� i��U8p���i��`J�`PB�����qq��H�a�r�82��k��h�ȓe�Y����-H1(#�_/Ik����=n��R��u�� (��˿/.��ȓy��u��4e�N���e�p�&��ȓa�`��A>W0:�Ⅱ�{\汇�B*�h�R�R�l�2\�V$ݎu�d���E>�*a�M' ���ӑ�
�0��\��hF�,n&�Т5�Βn�n-�ȓ1&D����ٜT�炊����ȓYB,�+��'n��T7N��n�Q��S�? Dl9V�R�(��x6�5 nH��"Op���k�1�`��c�, J����"O�l�G���^=���@E�l�'"O�Z�ȑ���L��&��--�5��"O�q˃6+Q ��E�׏r2~�S�"O�!��W�ę�c�6�[E"O6ث��Th�a5限/R��"O����E�>	C��K�W;*484�c"O�uBTo9% >�[�
�-" ���"Oh;����:@��©3���a"O* P2aѐ=!$��v���6W�Xٕ"O��x$�¿���� %KU: �"O��"Eg�Q�"!B��~^�b�"O�m�mӖh�8�:�F���Ω3"O�Ճ�NM��&P[�%ɫY�f5y�"O:H���+tw�!BA��$)�j�d"O�4h�N	�P�@��P�C���@"O�Hb1�޸K�����E���R�"O��ڳ���X�(l�@iѐ{��ْ�"O����ԆQA�����@���"ObQ8b Gezg�άr��L'"O���2�v����1��p�"O�`� ��\@n]@��0�~���"Or*�-�x�Ȧ`C�d�"�Yc"O Y� #ѓ"�8��n�s�`;V"O.�q-P/<���՝��"O��s���i��|
�OĜ?Ԙ3"O�jBR�$^�R3�S�{^�Pf"O�!��E�_1��M��)�t"O�a�J��M���tG_�>#��p"O�����h�Zћ�F��Op�
�"O�lA���b\(�����J�� �t"O&�����Z��a���>Sz�Y�"O����J�qP�`���H.Q<�L�"OL�E�Dn�T�#+ˀ&Y��I�"O�qǤ'pP�!�����0�"O��e�ɵn�H��<N��a*�"O�H�rf̬4r���65�T�j�"O�1�H !+V��ة0u�r�"O���CB������f���T"OZ�� �8(��i�#`Tx.
���"O����*?J�3���!@� �"Oxȇ���c,��p"lL�c�,0�w"O$H����O:@��
� +���Q"O�@3�W�^n� �fg_9F���9�"O��q�������'T-^��<� "O|5���;�Ȁ�VIȮy���"O�t���֐.Վ�z�h��[Ą�X�"O�1��O\����Qaߺ&�.B�"O�(����9�bT����*y��!1"OXX�RB�8��2͑8��sS"O��3gL��B�D�� f8�V]�'"O�A�ĭX74<P�Ąoqj��d"Oh��Ӭ
�	�.�1cc�`<��Q"OFy#Ug]��"���ĊK�D��"Or���b ���	6>���"O��:�M�r�ν2r��Cd�C"O��0��.9�,`ci@��Rt"OP�Kw�/$��hB%��MF�[�"O��Z6�5�K���K2���F"O�`� ��#����ƛC1����"OF���n�8'���r%�Ƃ {T"Oy�+ؓ,�pa���Ia�xix"O��Y�gÍ|�L}3�����Ez�"O� �M���,y��L������Q"Oj ��*=\���0��"���1"O4�1�J/Q�P]��a��5�2iC�"O���)�(s���Ua��m�t5��"O��{�$Ћ-�iQWAք�Z�h"O
L	Pʖ>Y`�B�j��;��E#�"OV�9��Q�@�<%�	A�VD�B6"O �RUm�N-s�'�5Tt%�"O ��ޜ&�܄�`lE/8�����"O������a��}0�
a�f@�5"O���o��Hi
�	�	�|��-zf"O�AAu	��H�	�rA>aR"O���%@5AR{v��*49ƭB'"O��#N�v�4�2��Ҝ~,T��"O -2�Ȟ�wFص(&�(K� j�"O�]:�/�||&u�(F7�#�"O����BT&�H[� M.;��� "O9�S��K�,��LJ!$'��a"O��){�"e3��\���"O赻�N�*!��t��� B@�e"O|90F�o�\AA��<m�b��&"OR��w�[�h��J#N�=���T"O �[�·(5͎�j�*T5Юx�"O&���	��>�ؕz�C�JVX�"O��[^�z�P	�@��i"O�PY�	�s$��Z�N!<�L�"R"O1��a܅P�\�h*�?�Y�%"O@T�VW
��P�ѥ�Lr"O�X+��0�*Ī�n���!&V�<!r���j�H����#\fH`�lSG�<�ũْr�b�+U��*!���i�FAN�<1@�`=M�����j�����PK�<���hi�Q�L�l��3�	>i�B�	"6S����.C���mZ�[v2B��3���iN�c<�xg��"B䉮+8� �dɏp%�X��L3M��C�I(N����ާmU�)�����{z�C�I�`���g��(Av�����/ �C䉹�Rp;���&
Y��ز�VC�I�:�]� ,.<d�G�	�pC�I�,�v�3�� ��<�K W�BC䉙EQ�IP�$W$ �"�/;?"C��-]��`��C�
e�.iK��@� C�	(L�^qb�(�$��FH��C�ɢ#H�$���_#�	+�4N*B�	�j\D�6F�'u�6 f�����C�I�U2�\I ��\Fะ��G<C�	�P+� %O�%r�����T�B�"sѪ��s�Ӗ[����bM�=Ob�C�ɑ|�ٳ����j5���+¶4�
C�9&;ƅ��0ߎ�(��@#oWC�ɵ_���R'E�26�YK� B8g�
C䉽�H=�^�x�d�!^���B������o�=]0xX�ޣHo�B�	0�~蹆Յ2�
���4�B���m����<Tܲ �#� /+�C�9WDɘ���v��BЅ�`U�C�I#:��iC+FM@����׵
4�C䉱oz0	0�ˇ@> D@���@x�B�ɿ^�&	K�.������oקF�hB�I*����Q�`�؍��#o�C䉻6��|�QBߔRn ��`��}D�B�I�@ƽIp��  >�T�	<�B�I+d�&�1$���𺧪�b5TC�)� R�Rv�d38�H�_��b�"O8���EQ�ܰ����%gw�1�"O4\���h|��m�*,�8�+$"OiaC��"_i.ȹTOL7.�!�V"O�����tL�%�殆fc<}�"ODy�B̊g�!IW�0�r��"O>Qǆ�7{�����K�,ز\+�"O(��5��R�6�A����#�\,+�"O`l���7C
�	7
9��Ԁe"O$(�A��f�vQ�41՚Mc�"O��1�[0jQ��� L�t��15"Op0k�fѪ>Ps#���d�HT "O۴��� ��-�F�����"O43�Ě(W":�j �@�^��E3p"O:��R���6�s�A�E��!aV"O��	2/�(Vx���Ѝ<�ʄk#"O���%o+�T#���e�6��d"O^�'�F�*�X��ousܸ+'5D����Zd@ J�7H���.D�`+�E^�5`�Y���2��0��,D�D��L ��U�錖MXlhX e=D���-�7Q�Qq��ʁy~v�-��B䉙F�v��oϰNB��;p�Z0��C�ɝ
4�$:a���p\�sNٝ27�C�	1sTz�p�A�k������j��C�I�2�|����$�V��̕,��B䉷y*F|)��͸tI��ɭ`�B����i��HR�ހ��E�_�B�	�e�V�q	��
�0ph�5pϬB�I�q�z|	K�&yY�}вC�w�vB�ɅYeJ���
)��4�ۄW� C�	l�z��V�F,b�U�'oWN%�B䉕F��X�W��ZҾ���
�}(�B�I�g��jg�Y7u���y@O��B�I*v^� ���(��w@[?:m�B䉋g�4l��	׎H:dY�vę;'�C�I�˔DI���
?0yP��	�|C��He#��AM=�y��Հ\�,C䉝%��l�C���"h�ţ�b� &E"C�.>��@��b׊E���e��C�	6�2��B�ܛ�m���e�\B�7Or��H���-b&�Y��ߡ�xB��3�Xa+�NL;|=2�]d�B�	�O:����{Y��u����B�	7.r�r�Q�9��؂ �ib�B�	�q�@�ai�9l(��b"�� �C䉊Y�y�P��EZ�8z� [^B�ɘ��(�k��Iap4S"���|�JB�I�1�(�[�����e�Y�W|C�ɥ$}�T��(�0Lh;�o�6{XC�	2�2�sυ�oe��s�\*0�$C��
0��1�d��h�*B�6KFC�	/CWX�y��΅D��Y��G�qC䉥)�L�
U�E	s��y��)� "XC��;;��$x�C� ��=���=�C�I�Xu�Hys���zY�EcVE�B䉩	����$�%0R�!��@A2oC�B�	\�ܰ qC��2V����┧�B䉮(
��0�	����5��B�I�j"�X����(��weAYÀB䉨p���Fܤv���H��BFB�	W���&뀸��H��#(B�I�:�@1�Q�˿SPX�H�r��C�	-��)��Ik��C�R�^ `���"O� `X���J[�8��E��h��$��"Oh�j�ܢ	=���J��.��"O�$��
U�$�3�ٸP�fI;4"O)0eQK!����[�Vh���"O�mP�O7#BXqz�JU%IS̵� "O�T��H�cڸ�i:5�j�*q"O�Q��-�Cz"��U�ڨjJpI�"Ox@ⵌ�P֘�ł�541��"O�,��$���a�sc]Puq�"O�P[���C���5��/T��I�"O�����=������*���Jd"Oε
v.�:]��q����hL��"O��Q�N�2�����7��@�"O�,�%ʶ��	�B���$̬��"O�yC+�:��px`��0�T�[�"O�����Q�Ȳ��\c��@H�"O"��@�ɿU���[�	�K����"O�xp�h9}3�Y�V
��];Liq�"O�3�♿~(�u���(	/x�g"O�T�æ��T@!�U#��~�*1s�"O�d��eG�jp�u*S��@���"O�m��A	v�`�saR�d�`��"O�`���m*��O=Gj��Y�"O@�[- ���0�EfV��"O <�bkA�[�X"2�E�FV��P"OX�)%�/d IU/�>��V"Od�C	�"�`��rG�L#Α"O��c�
C�O�~РR`O�6~�-��"O�9��*��@�	�ff���"O�ţQ!�?�����A�IoƜ{"O�4)#���#�PXi�I�I��偣"OPpRb��/T�L�vǋ�Lh(!��"Oh���Ptй{�`�4��Գ6"O�����}�R	�R��)��٩�"O�ű@��HΒȢ���
i�^�I"On7�S�>t��f�6Eru��-5D�8s�
��9$H8Ҭ�, j�h-D�����ՏY��$ba��>.@]�4�5D�t�"���8'�!��i�e08�h?D�����q������R��Y��=D�D���EG< �&�-m��ђ<D����/� KFI�+G;�e��6D��H��@�d�Q@�Х+����5�7D��K��6�<��(�<j�PES)5D�8�p�ҕu�Qg�H�Gڀ�s�-1D�X[G�C?^J�5��:M^�H/D�4!���$�ʴ3��G+|?
R��+D�pH� �V/�\#�k�0}J$���(D�����lDL���֗g��р&D�+�k�9^R�tKԬ_���;��"D� Z��IC���Ȑ�R1j)�m0��+D����A�
�VH��)�����f)D��b�#J�s�����T6W� �y�(D�Hb�	��p�$��k:N�*�C&D�|���y�z��*���A�$T�x��eȆ"�f�1���ڨ��"OD4�',O#_� �s���?�0,9�"Oh\0j�4�L�R%G�_���"OB2�#^�~4��)�X����T"O:Q�&&ل>��Xr�%	,|z�W"OH�ᣄ������ jАȶ"O���ό
v0��A��Ou��!�"O2p��g[�j���IԢJ�Ok�{�"O��K�(&a4L�AcE'TX�ܡ�"O� �"��&)�t"R�VQ��"OH����+HP�94!'�ĘY$"OhpB@"ACRH'܇,ƀ@"Of�Y�hM�@h���ڛjy��"OnM+�[�k(p�����>s�X�"O~Lkb��iz c���z�`C"O<$J� �R�Y挻]�$l��"O���3ϑ0C�����NM�0��Rd"O�8���[)i���:�B!xz%j�"O�l��,QI	"�
�Mުv�d��W��E{��=C v��n��ư�GJ!�?i"�i�i+���X��Wq�!�Đ@gx(Xu�B�F�Δ�A
�s�!�dR�<&1U�L|8C�+�R�!�d@�y�"����]4MU�3�CB4s��O|⟨�|�GŁ:FC��ڐ8B<��Ї_�<I$�G�'^4�H��}`ٲ��o�<!ӂ=:Z��'��.}�L�RE�Q�<���\7Az�4K�O��AbD�:�$�I�<!�"�%/S�5���m�֍µ/{�<���7S��l����<q�1�-[N�<�Vfѧ��.��#J���p��A�<� n�+��[��(Y�b��d�<i���&#�!�P���n͐� ^y�<I�e��jw��JsD��-��a�e�v�<�f��y�dj�n�"c�`}3J^]�<�7^�1\LI�֓{3t�Qs���Γ.I����ه�Z��g�0�Ҕ�ȓ}��*P%G� �"5�,U�l���f�h��.S��{A*[�]�܆ȓt��dJ�#�Bdr!Z�"݌9�����f��ph�ha���U=����eW�Uу����4�S�� ow�-��37z�8�۷UJ�2K߻=:��IL�'�����.WGx�1��v����y��'
��*ׁ޲$�) @�$� y��'��=��D�_ �D(�%0#v&�I	�'L�aKT��L��bgY'e�\Q�'3���%	� �Cm͍'5<���'�8x�T�u�X�YC�!o���'�2TC��J�+�(L\|K�L7�y52"}�B�[�nP|ٷΘ�p:y��lNO�	�a{R'��~hZqb�f��L�����'�ў�D�)WhܪZ�t�
v�\�w��"�"O�����)
��Q2���$+��r��O�Q�N�<���>ч�n��=p�͕+s8[�#FN�<10a�:\�hՁ�@8'�N)/kў"~��)u� M	w�C�,�^%�%FɋRSB��d�Y���N�A�vp���B�J��C�	1Q���$EV>x��-��avvB�*{�I��ܬ��̪se_�hB�	%����m�7JU�1��뛱b-�C�)J������[6��ab�	"DHC�	^ܘ	�t�H&0�`��&�[!c*C�	. �~	)'���c�:)�r�˱{HC䉘R�d���p�a�$�=N�C�h�	��{
���eƗY�B�I�m��ٰ��X?ik�U2��=XB�S/x�L]m�6�RE-�97gJB䉒j���#�Y=#���	Q��%"O�01�`)@��+���.Qoz�kq"O� ��Ë?���h`K����"Ofa�"ʝ�A5�����90��"O>4(
� c�p+1�D;k�����"O� �sD�^�R� L����Z���u"O6y��)�?��%��!"m�����"OB�[��"%� ���W$>ypE��"O�!�I�hW�����>W�ٸc"Or��$
B(#Q��ǩ[�^<��0"O45��j�+����g˗�yB�w1 @���ݶC^�� ���yB"�#2���� q ��&���y�I(. �M2���RdJqd��y�����MB �`�Y�m%�yRK��B�<�( ɖ�bj�1`�\��y'ۉ!wP<�#�k��e��/L&�y2
�#{��ii
�m�SC��y2�֋MR�	���1=Q~yAtH ��y���c�ĈTm5 |x�cN��y�#B6Ƃ�q��+�9�]��y��(s�:�!�JZ�&ZM��� �y�E�"j���&#�>��C���y�ˏb[�<�1�ѤJ[�k@��y���L Z����7I��DJ�Q-�y�^j�Tba�7H+��gς��yRjI�'\p(����B΀idC0�y�X�����F�4�R,+D`&�ybd��)�`�`� )�^�s��:�y��T�hӂ�KF�P$'FD- #�
�y� �و�	��C�j@��E� �yRb���nx*bƓ[���X��y�E_��c���Zژ���'�y�+��)��y)vHGR�tt�fj��y�C�;��T8w
߽wV(��`.�y�@�'0BY���sPpa�dn���yr�جh�x�6�qؼ�AC \��y��$Ī�@5j�leP2�6�y"�$��0��;���qvk� �y�GJ��X�yC6
���c���y�(h�Ƞ��*��z�P8`�MZ��yr�?Y@p��G�8e��!�����y�!�-�M8�M�rU"����y�c��C�,)Y��::�.����C��y��ߓa�h��&�$��]��ǌ�y�Ɇ
MҦ�[�F	�$xp�ü�y"�;�+靔o��t
�L�@
B�Il��A"ac�qN�P� �|N�B�In�I�'q�n��"@�ƘB�	DNt`��3"�� "2pB�	60||Cbg�/�e�%m�5�C��;����������AZ#��B�I��욱���3y\����8[؀B� �킅�V,(� Cb	dʄB䉈n���[cNF/3�x��#R�vB����<�`�G4�E �ݥt^bB�I�0��j�B��V̖�pɚ9Z��B�ɓ3�=� �Y��}�si�$0��B�Hj�B� �2FM���u-�3.ҦB�I�d��;�)� ٪�01lW�Yh�B�/b�2�!-h�捚�MB0xP B�I$2B8c��0��Zǋ�-2��C�=HF�Ę}��-0���>��C�I�V��B�!7/`1��"YM��C�I�x<J �����c\aQg��o�rC�&s�]�k^�	�NAЀ��i�VC�I>���c�`�x2@m{!fZ4��C�ɧb�0�4zg�xwE�c�B��')�ttȥ@�O�%��!�%��B�)� T<æ�e㐄��͋'M�T��q"O�3P�BW���0C,����S"O���`'e^���O�hbnQ�"O&��daMx{�]s��0EN.P��"O���&3� xzх�?F�AH"O���F��7p@l�VD�d�����"O��2`�T�j���2ǃ��Yz����"O`��-m�l�B��Op��q"O�L�� #�����N^Y\�`:�"OؔQӤ�=X�>�pR�K�u�6Ȃ""O�x��V�=!��5b��"O�yd'N,ZN��@˝�xIf\�"O�!#fײ�:T����/���"O����M�C*:��/B�t���"O.Ix&��
���$��$"!>D�"Ohm(��� �d�e��!d�H�#"O@E"g��J�@�G'2|{ʔ�%"O�kmX}�J��C���J\⼐�"O�}�tl�;4�U��V�gJ�	D"O6� �Z�!��;���w�l�Z"O�:��\ �v����O����c"O�\��^2UIdm��G�Dx^�u"O0��m��`N��)�?sN�p'"O�2DfZK�}K�G �p[�%#G"OrYs�D�D�yǤY�M@�M1"Ovf`�_%>��䄓@�(}�"O�a�`��?D�L8�e]�*�7"O��hiN.\�Hqa��5�b"O� 2FWQ��}����[4ڍ�
�'ZZ8��L�d.Ĺ���>5-��'�<�+���13a���i� |bl��
�'��������e@a
�F�h��'�FE3�����l�H�.͞���DZ%([ʰ�$H.d.^"�hA�"�!�D��8��٢s�0^3 e�v&�B�!�DC&��X����(E�($��K|!��p�G�!�c��Z�!�Ğ<7�EەM�oI>hg 	q�!��1�4HW)b>�,� .L:���R#��	 �DJ�B�i�9�y
ybJ����Z
^��8��X��y�	�,�G%YH�x�q�:�y���*�\tx�#NNK��jf ۙ�PyrI�!2�|��d�Gȶ!���FZ�<i�O���U���|��;T�]�<	�a����ÏpX�5��Eu�<�ƃ���9�!=�J��t�l�<�$��`5���`I	�X�*@C�<�A�0L>([vP{��qPa�Tb�<!f	X(/���.��|w�h��]�<1b��&���k���.1���W"MU�<i���A�f\�g�ǔk��Ma�QM�<Cj�/Q���S��fJ�	�f��H�<�wm�"�
�p�휋s��:���]�<	�IT	^ڱ� ���2������[�<��OQ�;o8p�R!%E��b�{�<y�,ӗ|	���V��4"��q�<���Į-\��0�� �(�!@.Ht�<A�"��al4#a��N&pXRO�p�<!�Z�u���Uؔ(��bI�<��Ǖ(�ԙ��eٰ�cr�WD�<+���r��A._YrD�i�<��*�6Cr��f����F�g�<1�O�/V���:�H��q���d� T�<��'�����=�D=@��ߐq�t���Я?���Y�"~�)� ���'R�KR�괭؞o��;'"Oܨ8�eG$$
hs7K׈=�Hx���']t\Pb�@�v�r�����
-ax�̘xsh�:3�����r7 ���=�`�R�t�C��0�N��֩[�-�u�g� �g�XP#���l����d�=^t�������a����GTqO�8B�'�"(���"� �R bh�,.�銥x�8ź1_�y��� |W!򤐁o��B1 �9��@&�ȡr�	0�f�*L��c
N
f�2w�ӑB���۟u\t��ʰ,��L͏Oġ��a��`p���K�.��ME1i<��V��U_҈���y�X ���X`��">a�� s8^ #�iX�$`(&�HGX��Pf�ӱ3Q� �$"H*P� -muvY�2�P<uN��Wh�|� ���.�}�A�728��E�:d#Zl;F����ēt�@��&L��J(BpF���p��D
l�*�' Ӡ���ʎn���T��+Ak�\��4����#D�)�"<���5��s#l�X6P�Ђ	�1_���aC�[=5��O���I�����	�k?��)��^�1��1 jIz(<�$���8�YD��I&���&��d�7	� '�����P�aب�*���}�� x���5>�v����5{��퀓��%Y�xr+ӟ!��!Z6#ϐc�H!��Υ��!!ł(%)�ԩ��
In�`!��W$�B�֧���e����L�
j<؈�N���'G٭�h�A�G��a��>{q��z�[�`�-@2�*s�A�>m��&	Q(�ybLD�<T1D�G60����w�V�y�M�E�b�1�`R]� �aW��>P9D��6 4���y�A �찰�X�Y6тTCֹ��>�t9l����(�b�(4h�A&0I�ub�)���2H׉F�Z�x���7\-����@�.+�p�p�ȕ�F(*O`��7#ŷ|�S��=��8��ɳ-bf��w�Ŷ~�k���8������z8���.��3��&l��Be�rn���q�7��f쌥f��	 ��'��IY� ǅxhp��b!�) @9H#+Z$zH�צG-��*�"1��q)R��}bb����($J-`c��'jlyq"��f�019�&A������&�B��>m|����M'�j�K��T&�ċ�͹T�Ȍbn�9�H)xO�nzȰŏ�%�d�{�Kԃ�y�!�DrhF#�$\VT(�ח��=y�E 'r]�!ȞɨX����j<xг���uA��M��ɓ2&�~����J?1�>��Q�Y�05#��|��3���n}B��t���⁋?C,��@ ��'��+�c$%"&�bqEx�x�GoA�E5�LJ"bO�q�������z�RE��}�#'��:v��GO �Q̲8��ANq�'�0|ɶf 3�(T��J  M(�k0�Coc4)h��Ç�
��C;�$T�&��7�8H��ꀁN:�#�oBh΢Y)�� }ٰM;p琫2���g� ��	����%�v1#b%�*A�Bgj	�3���a"V0$Y ��1��q���S��ٝ �hk�e�*L�:�*H�7��ט"\��u�SDj��������=6�E���ֱ��b�k��L��T�DZ?'����K++:MȔk
&J~���A�����"�O��L�4[=/������*�~�k�
���U�9�`��w��9��'��MN-P�6�C$'֛������1�:�buKB�VXJ��ЛQ�U���H�w�0��$���E��L��;WAܱQ������V����ɒI����k��q��9}���.@	Odp	��GY�Z����K����f�ot��rh�U�L���k*)�풒bQ/C���H��'�ʴ�r �	f"R��M��8xs*L�-F�萦 �&�谘�o�1�ޜ��$A�f<j�kN
H�� P[c�pR�(�w�BY��B�)���A�(lOR�"5a�d>�5���R�4��#>��(S��?�l�P�n�8:.}�SM��#�Z�� ��V�8��3�<��<{�n�>�j�IH��ђ�_�(U��Q���P���BjR�$�=3W�H���Ǳ/�$�A�>^����գ=��Q�EE-h��m�5�B�^2o鬌�u��7x"?�Vŏ;�06�\�3���{�jאnV�\�#��g+��
�h̼�r�f�O�:� "�,6���/f)���N���@��Ϛ�1Tr9�����~@z���4�a��X�!g�4xC���X��o4A�AB&͂4��!aLΤy�(y3� �5"a�<hC����@�����ygjP�4V�q����G�@u��!��0>�%ʋ4�z�e�Qg*=���21pp`��9��	5&"Z�$<;S�G]�搙C�
Sd,5����O�����Z�=��	î�gT��剡!i��×hZ�>����)9sj*`�&EA�L����bɬD%��7nP��toй/��BD�'� ���*��$q�&L	D<��)c�q��l�vo�ҧ�O�p�
ڀ}Qn��1�

6
P��Lɢb�9�7�F|H<IaZ�Q�<��ځ�Dt��E�c�5 ���޴)��\��L�.������c�|se�:+��Oz!�]4�6�jP�/@�ؐ6�B-Λ�攤S�=E��4|�¹!wi�(ݘF��-^�Lq��K*+��
.]X��RO��#Y�Th�	0n�{B	:q�8�AA�0�R%	"�˰>ib$Q�e� �d�Z^�ha�L<�5���;`r!���M��08�M�;y$;��O0/S��p�f�$Rh�>A�U	>
��Ţ�D	5 �`���,D�� �@��Y$,K�0�� =wm�x�V�'X�Q���Ӗn��y(�I�:��i��`'8�����a#>��PuVL���$�T�5L��8���'J ��ɬ���bc�U�3�ĝ�Ņ��8#=ɖ���T�n�}"��rl���77���9b��b�<�"�!<�!QG�L��I)��AǦi
���'�qO?7mV�p�R��OL�h9�Hc�j�,�!�䉼Ph-�T�?a��萓���&!��%�P�'��1�S�""5F ���%\3b���I	H�p�u����MV�:N|kT�_��@��a5D�Ȁ�逦_J�0� �Q3V��O0ғ}�j\�$ 3ڧmY�M3ժ��E��y���#*:@��O��]����9:ȡ�τ�8��I�;��?E�tL�$�q�ǃ�$T��A+��&�!�I�|% @a��'n��C,D�u�!�^.Wz��)^x楺��U�[�!��]!d�ӂ'_`Z\�D�ܕ@�!�dH��������92�u�$�I�!��	6�~|���/U?��f!�kd!�$��*2Rh��&��<)���U U!�$z��*CX n�,0/ף|o!��M&g�("u;�=kvA�D!���oh����<���T��A�!�ܻ|>�Q����\p�ee��A9!���\�1苐Oʺ� �$E64�!�Ո.��y��M<P��-�E�K"#!�$��(��]���x3�EzЁ�&!�d�=5�)+��K�[\�8��2!�$��0p�N�19��'�,Z!�$�- �j�	1��J��!`$�\!�D��:�0��_ L��2�!�d¡b�t�(���5a��+�*���!�0/�j���ɦe�BTJrH���!�̫J	�8 ��$�)1gK3O�!���i�������Qr��"�!��?3V���� ��F"4��FK�Np!�$H��(���>5ļ-a�e̤�!�D�8<����K���
�߿a)!�d��T�����k�@��xVB�-$M!��V  {��B�˞�@���!�a��!���]7.�*�.ǻ���+�!Ѭ"�!�$�'~M.�xf/�[�~�9���Z!�T�wH�����[<d��H��!�Č�� �-F�� ��F�/�!��ر��Α
{���� "z!��P���;�c�b��S��0g!�'�Z�ZD�Uh5��Y��ݜ;�!�d�%X��!���8'܀9b, �!��
Sj5���:
:�ҳ�T0�!���
�0HK�� e�LX~!�D��\o��zs�Q }Rf�Ǡ~�!��L�Tl��nC'0�p��kI>8�!�U�]�cC_)ڱ�ܥ�!�dһ�Z<�A���3(#�U2�!��E��H
�X��J��ċK�C�!�Ā5_���*Q���&	�:�!�G�?An���ȝ�n�
�&#���!��&��d��kC#���� �O�-?!�o�B9�!�I�l�Լ�``ؿTB!�K�(Q{�� g��-)�.��]<!�YI��0��޿�p�0�<!�Ėn��\�s$�*y"�`�,�
1!�dΙ~N8ih���g�(`f��n#!���6��(7�C�h�n�
�mL�$!�� 
����^y�HS��(+׶���M@�8$�ɅZ���
ժ$&���ȓ\���Ó"��dE�������x��~���q�f��'_
y!��X�?��A��*��Ti����0tP�y�/��9���!h���BM-}0��"�Tؼ��k1ĤZ /!- ��.�0 ����TtU�c��d�)�˛:�*���;2��(uD�+F)x�BV'>>��l��f>P�J�KY�{S��ǈJ�F$.Y��Zb�s3�Z*~0P8��ڢR�&��R���yFBƉV��Ɖ�*�$a��6������x�6uaf韗@Bi�ȓ�H0�q��:���pE�֎c*����IY@%0���8�h��V`�<� &E4*a,�c��҈{�LlhAM_�<	DC�.�"�Y��#&��(�%Y�<A�N�
*!�ݲQ}J!����W�<1��}-�b�'U.c�������X�<Idf�.x���C�����=��DP�<��&�w��!wdғb��9K�g�<)DC,qGְ�e��T=3rn�a�<����;��d��>o�Ah��c�<٣$T�Q��%&��@���$D[�<�'�I�N��G�&�p��b�T�<�Dn��L^�}�ĺ�#R��&hڰ���}{.�"�H�U��$ �R8����`�i#�K�Y`�x�(�i�N���A�@Hx����(�	^�Q!0�ȓϪ����֘x<�5{Gǚ:��I�ȓ,��	�3�]*�Z���J�
5����>u�dJ6�%c�&�ʲ�L:��a��EBT �)V��h�c�L"�ȓE7�@��;Z-ZQ�qP�Մȓ?��H@NB8K�������I�R��ȓz��p��5�X���G<^R�X��4�N���բYsb�	�/և6$<��*��1t�>� ��)4'Xɇ�_�(�"��>UI�,�1�/Sy�ȓd0`mT��5��'^>�ńȓ!d�����ۢ�@0DƘ���ȓr�@Aq�N��}�Bt85���9��ȓkt�hE�CH����tF�%=>هȓ*jZl���D�8Y�(��q�T�ȓ�F@�"�O0Y�� ���<�t��ȓ<Q��B��6e��aۥ�A�^�$���gp̽IQ�Q0{rƤ0A�R�}���ȓ?ʺT�`�1��xr��<,-d��ȓ9��"O^ M�~�歚�D�r���8\��
Z�6Nt��N�/怨��5����L,e ���,�q����ȓ5X���yp]��/S�mk�"O�=`�p6��w�܃]�=Ҁ"O��Ȧ�+�P��]�F��"Or!s��jwt�F,� ���1"O�d�ecJ�Hݘ���2��4�w"OV�
�(���E�T�Q.(Y���"O�=�!`ܤ&��H�R	�&UG>M��"O������"�H�(��وX��Dj�"O6���� �b��H���۠"O�	�m׊d�j$�B�/\Ōa9a"O�]k�A^+28�jc�M�j�"O��t�Ȩ�@�#�$i��II�"O(�v��-MZ0JAb�$�Z,�q"O� ���S�ɢ!>V��W�H+���"O��c���\���k�"l� � "O���CG� *�4!A��_g���""O\j�Ϙ{����b�]�O[�<YQ"O�82��c���k�Tl��g"OZ���C��/�R�`�ŧ)m6հ�"O\Q��V�N8� �Q�u\��:�"Ob����]��|j��T>fT��#%'D�����!�4��ǫO��~-�VD8D���Ìi��!H�GJ8d���8D���A�!
\�@��/��H�i3D�����Hd�콳c�B0CS�9R1;D�l�E?r�9A�o�p����`,D�Բ��HvL�F@K3�$�u.9D�d��Ņ�0�`P��jx�\���4D��X� ,xЅ�#bٸo�PZt�4D��p*��#5H֥-V�5���0D��1� �$/�P����0�/D��c&!����'d,,4zA��L�Y�<����>%â�p0��.H����@W�<��A5f����ݷM��af��P�<9��&DY��#��C���2b��N�<�Q�_uOJ�J�����Y1,!��!:E���qDM5F�9�Q�ۧN!�d�4c^>��#��,1��G�J�8!�D��w9@�1@,�l)P�;q�Y7[�!�D�	Z����d~:���p!�$	*��uK��:]�('T�!�Ņi��m���© '�2��Ca!�$�y���"	3��jRI$1!��E�.x�"%ђ\��a�n�&�!�DƜv6i�� �a���4#��!�K -��e���TԠ=�ac� z�!�DћtJ���-����	�LT!�	 c���/$p�p�hU�#�VuC�"OtL��LQ�w��h�R���F�8���"On]:WK�%��+2�܇����"O��
��(R|�����2��M0"O0 �SEL6=�XAhW�$�z��3"O���/X7%�rE�'f�"]����d"O<@S� �3ͤ�FG�_-���v"O`�����8��@0��[�T��"O��+�`�zEl���G&6 ˷"O��#-B�[�^U��?_�8��"O )q'������Ԗ6�"O�pt��:c��t)�.���"O�hB�ÎJ.��B�X~�6Es�"O��CJQ�O�6���m˖(�p�Be"Ox�r.�E+P-���
�ܢC"O���6f�h�(s�׾ �
yJ�"O�X�U�]�c� �a�8#���QD"O��)0	�� �ѻǥ٪q����"O��#��z҈Da%M�9�N���"OP1a�[�C�2y�͓�e[�t3�"O��C�\�=3@����ӣE]`X��"O�M���0C��=P���=P"�Q"OqqF��b:����Q+2�K�"O<����]�	3�=�e-�r<�8�"O&,`ueA�%���t�*a#���"OH�cV��+Zx�+��,~���"O8�pEɆ�y�K	Z�i�w"OL�p�F��* �D٩�8���"O��)�dS�	�\��񄇯Gې� "O�E2NՉ�&x��LS�S���D"O� �u�'L�Xl|EA�+�l�B�Q�"O�,xQ%�;P������-/���#"O�)Y�+(�K�j�C�FHj�"O H�a�c�1	!ȟ�)�� ��"O@�H��Ie0�l�1�1�l(�4"Ob͋0%��RC�	#�^#n���R#"OH0A0�۬Q!����.���[�"O,���J��-�B�2��@�3h�H�3"O��P�BJv�� 	�_��Q"OȽ��'�/���I��9�F��"O�=�T��.7^"ic�(�=�v@k�"ON���*�'�$=H�\�p���"O��hc�ԯQ6�����ꌡ��"OH ƍ;{g�yF�Obe`��"O����*}˖�p�"O?,"V��"OB=�cƜ% `}���[���W"O�D��$�2�B)y &H0D�(�W"O�q2k�f�V!ce!xN��S"O*�RE
�>:! �`�咆e\�S"O:�Q�J�_2��r���T�a9�"OtxrKܚ<��+�CT�~I�MR"O���$Y;a�Z&��0
;�y�`"O��)��*G�X������$�80"O����ς�j|B��ߴi�jt"O����m;,j��p6�r��}3�"O ��S��,����W��zpإ�6"Ou0f͸1ӄ\�a 7{Ϊ1�U"O��9� �T�Щ@�e��v"Ox c��F�?�\��o_4:����V"O:t�0��6���I"�<:���"O����j5�fk�&E.��	c"O��&l��'A\كLV��6�`�"Ov�1��''�z���L�[�x��"Ot#�,�5~�� �4��B,��"O@%;C"Յ:��K�4(�`'"OZ�˄�͙/N\�穊-%�6���"Or���R�t�1H�H��\��"O�< %�9�,A� ԕpަ��"O�%"��, ��f� k�*�"O�W�ϊD���q��%=��|	�"O��&�%g�0�$*��TQ"O���ޢQ˴-��ȭ�
���"O�� �'X>V*��aխq��As"OL�S��00Y��R��Pv�q�"O�S�"ه}+@Š4,�ۅ�8�!�DB7Ue�@� F�5I���L�!򤀧��e��k9�ٛ6�TI�!�R�7���휨*�ڥ�����x�!�P�e������#M6���qg�(f�!�d�i�(�ѳJ�0(����ɓ�!�D�)AJLӅ��$��`1 ;{!�D͞��Y�&AS�Ҫ=YFI		S!�č�3��1Y2��p���Qn�!��] a}4Sp���/Δ�Q�-[��!�DX�ծ	زÁ�M�|(�K��2�!�DӀa��A�Sg�J�g������2eb��bA�R�C�@�
��\��wnܡ���8�2q�B��!!ے�ȓpUpm��'y9Kem�
d��$�ȓ?��%�2���6B#����C�T��5py[���U�S�p�&����f���J��{ �@�֙:R	�ȓd� A3�Qr,̠�H9z����W��cgh�XW�D���;Fw���S�? BXP'\+:ցS��\20Έ�aV"O�`�T{X��f���4��"O<���=7M���W/�H}�P"O�$P� ��H��&����%"O��q,�#j}�*% �G�ح!r"O>�i��[1RF�%{e�00%m֤k�!��CMD1s�Ӣ ��)�&��!�$[)�Ƒz��Ө�DP:��n\!��K�hD��E�'t��XA�>p3!�$�!���ȣAX�Qжb 6!�F�!��1�v�ԅP�5x��� �'N�X�4�@<&�R�xhѓ9̆��'(Hy
���4�10��:��a��'�����G�?>�E�M�K6|��' QŮ�)�� 3fk��NV�M �'eR�����m8`�(�o��:[FA��'Lh,�7@[�r�\���@�k�`X��'�<���� �z����B�lw��'ɨ�����V�>�㇚>ko|d#�'Z�}�'�^�8���P& 2� !{�'fPI���ۜJ�>#���*��0��'�Z�跂^#N�d�a��C+�:���'����ஏ�q�b)h�n^� �Tm0	�'�`�C�Ð�h�Z�QD�R!��'P5b��0Ca�0������i�'1ص��Ǥk��s���	�\)�'�$�dn:�P,b������	�'Y"�1��m����ҁxD
���'횙	� Ζ0���:&��UP�'��8��!�Xf��Ztg���z�'���C��Ǘ �xŠE�M��'�2�cb�[T�JT���J",OH���'�f�
�f�NЙa�"ØJ@��B�'&�e��^�lҵ������P �';�Q�Clz�X��>e����'1 ���ŀ�%�E	�-Z#?�	��'�~䋠͖�@\������z<�
�'F~i���7{�hqXr�����*	�'��Xj/�;'Rt�� �Gy�v4p�'&Ȕq3F��>�&��҄:}���"�'l
��c��-Bv��׮��)֨	����F6D�憟�=p"�{�OÝ'P�ɛ~����?E��O+���%n@�t��"T�#���j� \_� �h�O@��S���t��DF�1�]j<!�&�C���iMf��vq���H"�^a�t�]�i2��'K�Lh��U�N�������������a�F�$]��2c�
c�i�hQa��$߱)2��8��6 ���ç����`��Ėd� DT�6�L= L�W�H9PL	�AFqcS�iQ>�r�O�u�WeˁM��	�
�R[�D��i��h1��it���R��5��#��ϓ�C��myu�t����Rm���醡pƴ�2b��L�`iK)6qt\��B8tkE�xX8p�ѓjN8� ēA�T0���Á7�9���$�Rp�i�2��HAF��Z����� ��D)Q�ϔd5:���
��la�h�H��Hv掩f�}s���-�4Ձ�Kɴ`f��pf��G���l:�'Ci���3Q5��Ӆ";~�i9D��fNZ=E�O?1\�7���0|�s@��V�ډx��˷y�<��$�?6]`��L�6m�'4���h��MG��U 0��9�₴h|h�së9��'ozq(��'&�cs���3i��	�6+"���
�'I`�K"	�]�����q�1�
�'l����/�.:8h�	%�v`q
�'d^Ad�! ��&�.2�~��	�'�P�@�K��l��h�-º	!�'p�Y6	
 d�lJ�E74���'>�|����k䅀`̦+�Vٹ�'��¦\R��a�ůZ�S�\���'J�M��	^��-hD��D�X�
�'/\�⥤�S���� �C.h 	��� �ÆoŮ7�X
g��#@,�R�"O��3WhE	5a:%��ɟ�S~�Ƀ"O�E�aZ�D� �I�* �/RXeb!"O2P`UЩn��l�$�C�I0lв"O��$V'\?&YЇ�j��C�"O�h����!�p��P$�
���"O�}	��̓z](j�0y� "O���O^*6���Y$� jE�U��"O�4�茨
�i(��R$M(��"O�IDC��`4���+?`�i"O�����6&@�3���Zi�@�"O.XI�b��j��M��W�`lJ�	�"O�嘖�ٶf6�2���bO���1"O�x��"�ztA��-I\t�U"O�4�T�@+&�q�e�ٯ)��<�"O&�K�/;!�BU0�L��
��Zw"O��jA�J��th�a�D s��� "O:-j���2�V8���9i��"O�z"�E�qy��d	�O");�"O cJ�G��¶�U�A$��F"O,�Q����S4��
F"k!�E"O�1L-�ܹu(�>]`��"O�Ԙ�˄�5�2Y�%\�Y
���"Op1��σ3J����	�јd"O���G�M�ry��D%I�r�"OLtOӨ���$B�d��� "O�a2���F��%�a�2s�Z\4"O*E"埈`���C�eOB����"OL�c�ZR���e��l����"O�y0��P, |�S��{�*�"O,�{ �J�	� �Q���#(.,��"O�ᘁ*�
�
1��Y�E~"�Q"O�PC��#2�`�3TM׵K�x���"O�k�ꈂɰ1�A��pi��h�"O8*� Nn��0�Y.�^M�"O^����B[B����!O�$��"Ov��H]�`;��R�DXl:=W"O �2ւ0Y;�ҥ��07h\�R�"O��8Cm�9 pڈ��ɻv�T�в"Opxia��2a^Q��,J6Go�!�"Ov��RϚ( �d�+�?YRܙ��"O����h�	���R`� t�~���"O&�$��F�j=թºF#��*�"OD���0q�(����"O�B"k]]6��Ta�="T�R�"O,��'��-	����� J�ud|C�"O���֠��x�� V�:�x��r"O��[4$�%X��X��G�>�ba�"O�sÁI0.>ĳWe�I��`�v"O2���x��`�ȼ1�����"O:�� �� ;L\�%��t>�"O�� *z����cA� o$��b"O����>[Ub���o��<S^Y��"O�\y�n�N��"�ݜ���Ӷ"O�A��j�5�} ؑi�BI��"O�x�C+��D�Dq�%	6�JU#7"O(�2r)ـk�Υ��g��&���$�'��U�`�8�m��ij���sJޛ]!�D�p,��F]'2���fD�q!�dڍi�\�揭wz a��=^	!�ď\n�M�rl��,�Y����!���/��/�`���)zH��D"O�%sdL�=Wmv	���/d6�� "O��2�E��Y���G�&�]Xf"O� �e���X<P�S�(<)|Cb"OR�#gG��)�jU��
�Ń"OZ8��̔q̘Ljb�X�M��{e"O�H����pрhH�Ɲ�)Z�r�"O"X9�e������ڇa3RDXV"O<����-4\Qa��OC޴��"O,tq���M-� b�/B�.4�j"O8��c�A]� ��S8�̕��"OLСb@�1V�Y`��ì	��"O`Izv�>M1��#;�P�HQ"Oڙ��G�/D�N�S@�
���"�"O���ƀ_.ߊ���,S�{e8�"O ��"b��H�a섊x�}3F"O
]��`�ç��%[lP#c"O�k�������H�?jQ���T"Oj �fF�Ary�6(M?r@ ��"OD��FAo��u ��F�R'h�x�"O�Y���FX�-���jR	d"O�\���Z�h��l�׆I�-	����"O��pԯO9	��!���Q�:mr"O`P�8e�����i��"Ox�K��=- E��JR�?N�Tc2"O4���7A1Pi{��Q�����"O�ȋ7�)G�5���ɓS�e�p"O�ȷ�)r�d����"X�R�:'"O.䑲(�5	3�Y�e�]�.�@�"O �)�N^�Dc�(K�C�>:��33"O)(aU�d�����!R	I"Oh��DƏV7��8��9��,k�"O�Pk�\n�4	��� �3�pUb2"O�e�B'[Y�L	6���p�>�i�"O\)��0,��a�?3����"O�d ץK%s�e�"O^�B�,q"O��k��S'&&�TB��FZԐ&"OL��/_(1�� P�Ç5+
x��P"O<-����2��� �G��3"O���`��4�^���Ex�� "On���AP��`zsa%�j�"O�=�ु)*MN��f#B�O�x2�"Oڼ�NR&U����,Nb�d"%"O|x�Ĩ� d��5j�9X���"OB(H��B�$���	j�!3�6��"O{��°D�da�B*�d΢@:�"O8�#$_&'�q�i̦}�ZD�"O��!�5)j ��I߹��1��"Op���֩X���8 ��9�&�ڣ"OZI�'��l].9�!*�S(>!�U"OI�PaK�K�� ��Z�^��ku"O��ˠ,����s�ȮWXɋ&"Oؘh�F�3�N�Hr�͞_�`H!f"O��"iK�R�d�P��k�p�҃"O�q�#�Z�{�G�+M�U�"O��������TK�I�:uN܊6"Ob��!L�zQ��z�i:^�t�6"O�%�G�ÔX3G��31KJ)	�"O�DSd(��^U)���3P��x�"O����	�	Y�T�����nB<D��"O� �4l��u�v$вYQ<���q"OR�b�C&OJ0\�g��y-r|�B"O0�Ѳk�' 8�ͣ�X+G$�h%"O�����0fSlP��Θ;X�:��5"O��;�`Ea�xt�c� ��-S3"O*��BԁvXN�J7cܛ~R�:@"O�Ӷ���"�:�@�9�8)"O� �)3�j��D� ĉ��Y/}6���"OpF�<t+X\���Z��鳗"O�ic
�i���-�m�|��"Oܥ B,�:5�"_�M*�C�X�<�A?��=j��«\�����Q�<)B�(�Ib'��({M��:���P�<QD��\��L'd|��,\I�<I� �7I&� elF>'U@�2�cIn�<Q2�\�|���r���EL���LP�<��O��v�@�D�8K���hԠ�U�<�"l�8�.)Q��^�2,)��}�<c� ��u�卡8�0%�E��@�<�䏔�gY��%��$x���!J�@�<���h��!��G/@H�\���v�<)�OŊZXN5�I�'%^b$P`�}�<)�.�1k��5`�G"p�s��{�<�W�ؠbt�8C�&7sf�d�/P�<a��̋�Q�S���. ��C��J�<9�jӎN(��q4�A1q����F�p�<��'L�e�8��ŉ�����#@k�<QՏ�[NQ�u,_�|��V��f�<)�Ԍ�ޕA�Ipf��0��j�<�
�9��5aD�w�����JB�<� j�m`6y��LU�Y+�m����z�<��G]�9�@2@(�6$�Z&J�@�<9�[H�Y!��i�hb��@~�<��%��qi4��b_fy@ �C{�<�#o��s��m��)��~�:�0�u�<ick/Q�4BE�X6{���#$h�p�<QEϹ9xФ��<f��c'K�w�<)�Ɗ�:2��O"h� �V��t�<C�Y�5���y���!�$�z'e�<�"c@�b��]�`JB$���f�<� �0����/OZ8	&D#�y�<>��s���6A����y��p��%bdj��	pB�c��3�y���m$�q0��#����A����y�äBFR���&�D8��a�Ĵ�y�m>��l�pN\�U1J���\��y�#��3 >-�Ȋ�a���#"Ǉ�y��9eg25��KO?O��-9����y�a�$l�X"���B�6�	��M�y�
�:e��(q�#�!p���QaH<�y�	�&wU���2�ܹTɎ�aA��y�h�s	��BJ�F��{�K8�y�쓧}�ʑ{L�)s?l�[ ���y���C @��EiONH�ש�-�yB+�_�2�! Eۃ����K߼�y��,�X���)>	(JX���y�)Q,D�;�&��`�4�P�y�HM</�����m����7˕�y2fYَ8�Cf�eX�X���R�yb<a��Ps���s����&�y�E��jW!��f�)�Cg�0�yRk�8muΌ��Lϕe���ò$ܴ�yB*{�0ROƔY/��B$+�y�K�&����s���K�<��ҫ�8�y"�P']��P3D�̧L� =i�h��y�	S$M"���T�������!�yJ�C�(��'G��\�TQ$G��y��Ђr��ܩW
��}�������y�ś88̄IR*#e�|ɸ�T;�yr��)���/٠h��H��fǀ�y�Q%#՘!zaj2(T(��!?�y
� ^�Rņ7����'f6�($"O��x`NQ?(~�!9�F�� ����Q"ON�c����[�({��O"�x��"Or�۲��&aW`���Y�xr��"O%��<����)��BY�Hp�"O���v   ���.j�N��I���PF�{y�S>��)������g[!yq��
!m�O&$(O1��[Z��	ٟ��	yy�'��arD��s\h��c!�"��EZ�@�	̟��	���<Q/O�}#�M�%��u�'��+$��Y�R�#��`�%��@������~y�kG(��i�p� ����h4�E�d�.`��П��	����'BB�Js�8�˖��sl��bM].u_�I������x�'�<�JG�/�i�e⹒��ηC�Z!�nW���O����<i���h�fՂ����-��˓D�,�r�
|�t��"�5C2`i���\(N�#%l�k-"�4┠+�()��ߩ	V�V����s�ٙ4z�������IٟhB�Lء"���ğ��	Y��'A#ga��<���A�p��� [� �Iצ=��4���'���Os�S�U��Qx�(4o"�Йu��@���$�O�j�E��e.�I�WO�1m��7�Ϣ\HH���ܮr�6ȃ6�"�F����!j��1�o?m8B�I���Œ��J�GS��
2��l4��[T0��%��%t L�o�h�F��d�%AJi���1
�N� g��%h?>1!����i$�0�W�l0,"�bD� ����\-0/�e����?TG���$���2�A�� Q#6�H�4��[[1`A�$'B�c�#�:%4d�UO[�`�L�a��$MN����/n�H!�Ҧ��&�M����oz�)vA���Hi��N3-08��g��Axl���Q�S����׸|�84J������.\$�M#e�^������"F�9�p8�ΔMx��KR�I��M�t�۟t9K>E�ܴ0���c�ř�Y�+�\�J]�ȓM �����Q&Df&�	C��#���Gyrg$�S��J\_�JZ�bȟ4��l�Go�
r���D�O|}�f��-?�F�D�O����O�l�;�?�]�P�@���O�b݊`&_�<�z���'} �'��%? �q�p��~Fz"�!P;4�Dk��h%t�9��lr��	~�d��U���c���ȭ��� k��"{�>�;@��L�p���N�>��	ȟ��IZ�'o��=W$&��&FWV1��L��j8C�Ib�zE1�
��j�:}�'��6����A�)b.O��`���^dJ-xDo��N-�a��/���J���O���Oj�Ě3)d^��O����d9�|l�����_%!�Ј���O� ��2�A!_� ɇ���HA�O�vY֭+7�:5RR��*F.uh��хP�@�h,�Q�H,<����b �#.qOj`1@�'L��bߎk߬e�ʞڪ���i٘�y��&J�f�سMN� O�|�1���y�G�T�h��vg�i����~Jm�$�OVQs�ǔz��'P��m�59 ��Tc�Mp��6���O�?���?����cE�q�I(�?�O��J/���i�����p�ƺ�HOvɥ	W�����foǚ_�<�O�P�3��SQf��ǭA�O�P�j��D�f���'������iu��(��[��p�J��O&���
�JL������:� ��(z��|��3}R�7Iv���CKŗS�Żg�Q��~��0~#�6��OF��|���_��?����M#�ߧW\2�F�)`cT1B0t�V� 1w�)��r���T>��|n�3'���.ȬT����W�&o�7̤I�ԡ�v�
��D��@-9N`��,S`}j4xH?ט�B�
�J�HĿ<�8i�@�q�v7�_�WM�*1��s�TIۗJ�b��%�f�͕�f��"Oҭ��v�5�I0v��{�ڗ�Q�����4��6�P�v��xj3睞mP�kV��r�1�I���i/Y�f�	Ɵ��	ȟ�c^wM�{�? ��p���4�#�ዑ_y�	�O��?�]%dt��Ȗ	 ��3�-��,�5B�w�f�PCLLj�Xѓ�jG"���Ւ��<	���a��'Nߖ(YE��dyR�S>����"����H]���C���D�9l�b��Am�f�tP���L�4q�M9��p���g!�$H�j%�� @���a�U�J�(P�������Qy�-�"�����N&j"<�IƢ@'s{��1�����'g��'���'r0�(8P��'��vH�9��!y�Ș�{�*yЇ�ǻİ>�R�TV}b�>G����L�$��r�!°>�c�B�LnZxQȹʗi��DԺ��F�g�B��l���A
R�0�|Z��+$��B�=U�Xb@��&z���
%{
X�ɼ�MkI>!�[���v�'6�]?��K�8�DTQ�:��U�D��BD���?A�Y�m�������	��E��I]�4�q@�>O���dSGO+�p{d�V�R�@���kD�,,UDz�(B��?�E�s޼�����*�3R%�VB��BXd��7F �;O:�Z��Y2�����Vu�ĝC��"�F,Yj¬s���">���nz�n�����[���X6�B�'"��	�,MʖEH�G�4'�>�E����Ыg�U�3<�!L�j�2���|ڏ��4��0�$�C<�.D��Э6U�mڌ��|���Z(�¶�N�s��a�,�%�~�1#x��vk��j/ xq�h�6Sp�oZ��f��I@�)�禡pv��pE��IfMG=N�D��S�<D� d$K�k����L��	��q�h5ʓ(w���S�=q�J�m�"pB��-��h����?����M	���?!���?���,���O'
�2�V		D�_Gb�Ф^,y���B�j՚DH4� 'D]�
u�
�Gx�DƴHErأ���V�,	�U�z(�Ȓߴo|�§J��b����Y?��P/>a�l��T �S?/��%��m_�uF2�"�{}"��4�?���'�n��D����Ђ�5S����'t������9��p�RO�'0�Bs���Ԑ|r�[d�@WLU�E���P&ώ6%$�
��r�r�''R�'��@��'�r4���c�XP����F��!��I����l��XJWIM�n�܀S��=<OR�+O� Z� C�!�(Q~����n��rdAr��:x�L����12��`�  �Mb�8�{b�R��?QeZ�Fsp!��+ 0<���P�&�ZB�!:��I�H�0�.�f�5sC�y�f��Į�R"�` Aʴ*Δ����M+M>)Go�3���'A�W?9Q�Z�Nh-�$fC�� �Y�M!a���?a�jN�����S��>a$��Z���	�V����Nh=\ ���Ax����.�r!�*GJ��%�>v��qr4]Wh��FN��6=���7�D5���ɐ�(����'ʞ��,H{��7yt9�"OfAiN
�R��I��2:���'4�'#���叞�^	�L�G*��iY�'�L�b2Dj����O�˧x'P����?ݴ:�\��B�-$�X��#F�B���/� �"�T>㟌i����|bz��"G,�f`Ӻ3��)����c� �V<�a@[�r���"��|�||CV�'�1O?7�H�A.�0�!ɻnâ���FC!�䕻!�d}�FM5��XvŅ+/Q�D	��T>y0�@� 򨲷�)�f��R(��?	�H���]��?a��?�.��N�O� �1�2
���}J$;�����d��k�a}��P�d^F�ɱOܡӨ`[�������K�a}�o� r&d{�˛;�[f�����ۚ\�$<\O�ak �˻�%;�A��{i��R"O�\k�cE,^�mX��o�&�;�%
�HO�	6�Ď=(�1� ��Q�����Çf�4h��/����O��D�O� [�`�O��D`>ucg��)j�*�a�1� ��
\���(X@i[�)X��"�"B���S���	|�������X��a�c���M��0i]�h����ŋ�=:tlZ�&f�KC��-Ԝ=&��kC+�O$8�'��:F��4sUɋG��Y��L��y�)�87��%ia�ޤ(}��-ϔ�yB��s�EM5�Mcա�~a�֒O�p�AG^æ��I�\�OL���e�9�J�{QdB6����ۓfQP���O��$S;y t=i�����u¢�՟�us�t*���e���hUe�EY��Ez2i��D����)}ޢ|���>��p�Ӵ/��#�	,?�H�����V̨�Z��DlܓeP@���t�O��4*����4yA�eJ?�PB
�'�&��@4��D��f�� ��
�J�q
�R���s&�푤�A�*\f]�7Fr�Cq�i��'<�&A >���՟�mZb����7�\�<���q���B�^T����M# %��=.��Z�����"�s�� eXQ� r��������)U�il�d��@�J8 �pc%��	Ħ������̑c��!#��k�U� ,��kRf]3X �=��$Ŧ�* �Oީ'�"~n�)�aCe���"@����)�B�I0!&����	�yf���S�<���i>mZ+�m�$�4p��ȵAA'rަU����?U���n�@*��?���?�������w�j�I'�ƏcMHDq��=uĤ�0&lK�tF�\0��6nbDR��F��	�@� H>Y!�8B���#��ԣf�,I�&�!N��7.?Di��I<Y��E1��I�ɸ��}\u�1e�#9���
�*iʀ��'����r1�z�F�Ir���U!*ƨ�B��yB/4[p�SĂ����2o��Dz�O��'�f�{w(��5<Zl���N�Y�X�R��C ,��3S�'r�'�b.	�59��'��i
����i��\8!��������E2l�X�s�h�'��e��\ s��A0�P�CX����e�O�h����T����61g^��ɗ�
�4�?A/O8�$6��|җ�ӷQ���������XxPLGg�<qd?S���p�bT�6T�Cc�z?ӳi*�[��)������O���D�.�rX��xc�0>��5��/CM�R�'��N��1���%��T<DP-���ڰ^?�)l�>>6ұ����b�~��Ү)�_.$(huB�(����A�*C�
L�#�YKh!(�-��Z%�%��-�����r�D�D�v��O���;��1]� �b�e�lL�0�G0��I�$��IT��)#��.�4�4�À-���c��=ǼP+���+jE|+�k�g��d�)@DUo��|��i��(K��2�'�����&����E,K�E;�-�>OI !���o��`�����t�Pb׆�K���ưI	B�\/D�~���]?�|H	q�ipJ�������N
����s�1�C�8"��IJ.{��p t�q�NYW�'J 7́fy�������L)=��!�H�o*P��2��~��'a}B+�(4`}8P�:m��Dk��ڼ�(OR0Dz��O؛V��Y����aM���@�l�8� �D�O�d�t���Y�����O���O����?��4��)X� G,2�D���j͡I�\���O�xCpM�>I�>����D����ڽ r�tg��-������PD}"#�F�c��zhX8L<<�W?�J��Ֆt��5��Q?��ͱ!L�Ԫ� ҷ]j$!�Țr}�$V���47�zb���7��ae˲fs�P�H�y��܀�h�9�a�eZ�B�$�)^0�Gz�O��'��T�N@K�J����3H8�}�P�L*+_�l۴�'?B�'�2� K�R�'�i�1�Z��F*	�,�`x� E��
?-\�����*�:<���Ĕ�8�) �(ÕO��p#���"���rȋK%��,�䌫�ŵ5f� �ݼ��'4V���`|f������0l	��èz�m��!D��*�bR\Q��(/-��$D��J�"�Wؘ)�'fZ8.��xQ���D9ٴ��3-�I�bR�|�	@��O-�
�SR�	�2B�Q�bӯA�l�.�O��D�O�{��Y&7���;Q�D�+���~�4`Z� �����NQ;` �CT�'[x���K�G}�PJ���5S�	�s��8�깠N�%{!�UJD���� S`�Д�=a��K��� ٴ% ���'V���*Ir��痒Inͩ1Ϧ=y���������b��V�n�
%N�R�v����4�p>!&�>�R�}Ҕ�˔&�ę�CP?����N��v�'Y�X>�lF�L�I����E7�b�� �͢b��°��(d����@*�:��4���@)%�hX��(��8�H~J^c7v�kTH���)"�;cl�,_�p�F��l���Q�
����mP#J4ج��C��>��33�P;e{Xx�b'ze��2��F�b���O���ߦ%��i��M���U�1_�	��b�=^B��CV�X�Iҟ���S�����U:W �>B@H�5N�&m�8AGyrbq�,MoZ@���u�l�D�f�B��_�O�v0�f�?_�����O���mQ�e��d�O��d�On4���?	�4<(��t���E��QM8L�#e�O�8�H���<5r���k���D� ��ܫ"����~-H��hbEC�fd
�+
	%��`��A\v��ĦY�Q�mo"�5��m�u�YfaseJH��p�'�*����5Q�z�ϵ"�q���T&�6���HD��yr@O�y̱�7 �87��~�R��4�ΓO�P�6��oJ��!T�F�G�@�o�Ѕ�%��O����O,��J�po^���O��X�`T����=&i$�N��/��ԫO�n� 0Kc L�q������<Y��0�bB)X�>yӑ�)i�a� `�Z�K6+/��@�ҩ�# ��Zd�i���I,2�"͕�E�Ju�rF@�S�pac��%NS$<��qz !��o@5���PFM��p�ȓ��	����(=�F �t�F@����{0�F�|⤆��b6��O��D�|2���(O�
)RA|Ly��-`�]���?����pq�ў;,
_q���ڟ�h��}��8h��S0"��F�	�0m�4���#WZ�0A7�1/pX��;.� � �ോ��_T��b��$e�| [�O�n��� �'��O<�nڷ��'�M�i�6D:���6x���ʆ;Y�����O�M9"��19j(�0���N�
���')��'���J�`U",C���mI�M�����'@0�*3"lӘ���O�˧l!E;��?q�4}F�Z��7L��`��!c�x���̱=)�¥ORE���3��ˡ,m��ʘ�5��53S�L���'7��UY�F��M�t`ĎiΞ���$�� �AT,O-�u�(��q M?�X!Qf~�:V$�%)*q#eO�\�7�L�SQ��'d�韌#|n�+S�t�R��T�#��yvOL:?����,��	�P=8���$D�����AΒ�<��i>�nZ��:�PC�Y?S�*��bn.:�T�"��?�W,ͩs��Ԫ���?Q��?�r����df�XxQT+��z�,:v��-ll�G���?S���cuvYʳ!�ID�3ғK�IA��0DmXBFTuF��T
U�O�Z�c"ڛc��q'�f���*�ް� �@gy�Y-D[����F(*�voE����Ư@1"�8\O�E���W̀\����Yx>�g"O�����<p�,���M�zجKT���HO�I>�@�;�\�cQ�D�	�^u#`KC��(� �/�/�J�D�O����O�X)P��O0�df>�yP)��͔��	_'���M�A�V)����3C��Ր��dx�4�Q �3j�&I��h�4���I��Y�1��)aR��+�:���`�H�k��U&Ɛ�!a��cL��]8��M�l�^���3NP�S���ȓ��(�L�uˆG��8Q&��ȓ�p�k��L�1��T�r�	<W>!��#����|".P�fN07��Ob���~�х�_?0�z BB0(�45a�U��ȅ��'/"�'��9��+PQ�x{��O+8���b,��|Ґ!�#��!�'�A"cH�4�!ma�'���Í�F����bǜ�2�6��8|r0��?wo`@b$&R�@ւUXQ(V�q�v(z�a(�Dָq�ni�<e&>�oZ*AR���ƒ<#4tJ���?!�x��������bM�a���ӣȺ����"���p>1p�>�$�2`�� s"E��؃��o?�%ٓ8����'�i>��{"��p�N�s��҆�R�2M���(O���$�Avq1����j0z�T�,��d&�B���c�?��Y���'�ў𺗌p��=[�G���p5i1D�0#�ݵ>���L��Z�v��N,D��s��|���אy�(ôH?D�p	�C^�Im��h� R�D���.D�0�e��<P�p|p��W�pR=I��.D����`��Bt�-@EB֚C�h���G,D�s�X0+~~�8e�яdRX�!�*.D�`�����{�
H�K�#D'4\I*D��`�K�� ���C��z��H��7D����J�3L⩉p&Ӥ�ڽ��A3D��*�mX�&����oшp��as�C*D�X���B�P�)!��)=�J�"��*D�h��jЇxҶ���H�>s�x�`�+D����J�%#�b�34H�zI�2
(D��hI�R�EC�D!w�����'D�P��EH~�
�Aĸk�d�Ed$D�@��W�H-����,VgƜ�Ba&D���� ��*�F��r�r@���%D�xʌB��a������8f�,D��z@g"X^�Y�uD�$7>�qPB�1D����ԑ(ܤR���u����t�,D����~���ôk 	�`�-D�|0�H�U��P#QM5M����`-)D���OD�%BBق���T��B��-D�<Pfo��*��) K��\9��H��,D��� ��/�M��:RfF]�u�M|�<q4�ի$�����ES8x��d�<��\�j�ꝓ�ɏ�?�D�#͛g�<Y�`H }P=�	ZWq��&&�z�<����R����C�3*=�e�ӆ�S�<�h�2&���
E&��k6�H��u�<���/�4@˥a\�`K��`ՠ[	J���C4�~rŅ��Hb?OF@���o��|����-a�CODP���h+��s�k�!E@})�, �4�H����?F�p�`DT�p=	A�޵iP�f�M�$=8��"�N}�'�6�a�ڄ4@������8�J��g� L(cP�P�P<����*���9"OXl�.	X4Dm �D�#Np�ء�^�Ĳ�C�']m��FN�t+8bǄ�,��BA�'N4QƢ�;E� 'n ��"O:YP�I�Iͬ:QN3K�x���I�ֈ��T,J��)�$�F:��O%�y'�H�f���iD>�����)èt�aD�o���V�'X�1��
7BL�F���JX���_9��P����#$�D4� ��h�,��p�v�A!!�V�p�?����CA��0���~�U`�"Q
� !ء �iz��@%��_iT)�Pk�	t	��yB�f!ɶ��
\P�U&��*9W�R�9�*4[��ì/���Ӌ�pt�	������.�ݙD<Ȟ��`K�>/6���Oyތb��?�VKH�'����'�-�@ �7\O`H$:b\)�!߂���� �a1�d�B�BK5ڮ�ȵ	J���9S��G+��q��Z�]���H?m9�ƛ��8�6/����hQ�GKt ۔%�:�� S��+�+�D�HS��; A.��ɏc��	�7+��NJ
*�(�c_;�f�R��،j����#h6��j�.!���NK-�'@ $�1qQ��!�1{P\ IR�ӏ{�.�iU����
1�eD"�,݀���Y?�uY>.+�8!��>d�e��X����C�(��z� T�����T66��b�)��I�w�`L*��W�W�
�b����6�2�Q�J�.��U�2f�5w.�*p"�t���1�����ᕃ�J���MV�E�2HI#�ۍ=^1x�K�:���b50�\q��$�`�p���y��7]o��l:Mx e�!Ѽ�ɗ�V���~�Vα������+"�az�ME�o^�<S�I���T��_'D�Z���N1���I�� �vo�	i��t%!V*�8�*Q;�L!b�&��i�`�.��#��Gx�ʧ]K����W��	t�@��9S����	����wE�GY���%�:r�<���H2zX��(��:[���DE���m� +ZV�;	ˍH�@����S<��	1҅��P��ȸ��D�)�6��CZ������'J,hy9	��Q�4��*n�	�g�F�8���0fM�D��bQ�݃y�~�#�~B��1��t�buj ��
#s� �0�΁/���p��&+�"P@V�]9#���'�4I9��0>�V�Q�'�d�N�A	R�V2�sEsz���	���I�Q�l`b��89ze�ркi؈|K�N �$������6
��&��5�jB���~��9y�@���GK�[��-���I82����w�=Zt���Ul\�iۖ�#�*ظx����f�x�fd��Q���υ7G�p�k�O+c��dq��H�p�^|c�G;W3��J6ω�3b��2GoŶE�|�{U㎩f�L93&*p�T`��cj׌���Oب]vq�H�\?�I�^DFl�Wl�,	��T�b�-�0p�D�<� +�E$`���nB�U�&�wa�E�8����K*?�z�
�K�}̝HD��\鶸�s·�Q�,�W�\	D�:�����+?�r�"�+� ��|�G�c;Ua���&? P�팄x?���#��<��� ��|�'��d9Qq���'80<`�̓o��@����&��@{S��:.8,�f�i�4a�P�]nb�i�g�i
�E�r�'��KC��5���� [%,���k��< $�h�/��i{n�s�+�9$I��[���#��5����?���#B�K�$*�H���3js|�# +�;"y��S����2Qa5{��E�'��9A �q�	)�q��L�6zv��o�E8�1u���+N�8��ű��I�%�ڝ���Fa��@� ��*ɜ�hb�/�j� �͇l�"�H �ʡ��*Gg��phQ�A����ǂ޸s�D҈�a�"ĔT0a�W�vέmZ9�Z���J$H�Z��@��~���u���	~�xU��3�} �&�تL� �I�Vy*�@�n\���ʤ��p%��ȜStAA	`L���á&P���g�&	�o�g��"��6,{�-Q�Ή�B�")�'7�q�l��pF��W)3
�b���`��ȵ`CȑP�>v�PGJ��:6�]��;wd���gKv�l���C_�dD+0�F:~�pH�J֙>=�$;"1�V�S, 0��{S��Jכv $��`�u��ql��)pI�|R8
r�O�\Gj�����Qȱ';VHh0h&[}�-p A�d@�5�ǁk�q�� �I.Ruʅ�O�9P0^d��%��e-��a�K9a"h��m�1Z�q��3���k�"�ͦ��f� 2�L�cF�v�T���,(gj�<X���-l\��v.��tR��`�_�F:z����#?���s���m_�ؒ`Ǩi�n5�w��"
�9Js�,�`��6�B�E� ��1-����F)j�`-��ě�'�%r�	�VL#���*o�6����V2@n�Kq�I�,^Pq��O�Q"�Ň�X@!%�Z/$&�l��E�(�:p�&�P��"��ɵy?L��B��h�j�`��[�' �t�wD�,ŉ'�R�k�[ =-P ��G�"	�XQ���
�m-��Bm�<�9�Zy�4�߹G��8��@��]I��@�^�#��	��8���� 9��'�����P<n�3��E�-���|,ݣ6��352F��2.�1j���bP�j�
<{3�Ŀ+�0��@�~��rT ��3�ژ-�4<R�Ùn��B�I�`�x��gfB�>Bp�Cl��r^ҬK�-��xe$x��4|k���.Kv̠��/�Lz���7���)覈ͻN���y�kt(Z)���) �ֹ�����ؙ��눟1QF�16�N�z�2i���Z�Z��EIc�T�cg����S;��}�E� s���fk氱m�:��'j�D���vÚ�
�.@�Gݼ4����&�<��.Ρ,��/c��P�K�	h�T1�
L�T��%�QH(��C�@����b��\�K����A�v�'���XbpUAK��y�!O8h��U��F֗rٜ���o�����4yQf��uE�5"a>�GI�=>���Ǭ�Yd��������2m�\x��I�~ϼLP0��v@M�&��4]�|%�D�5�8Q��%k�e����J_^Xxp�	vL]�vo�6�M	ˊ		b,��\+z�6�����"z�P�b��T@�' :�#�*�'O���Q�(ޱV���u �<t��XF��=	���(���s�����F�b�:ћPk��x�`2�l=.h��j�<
���� ���7B�����(e����#�"Sm�7mH�t8�9�,�^|� rjM�*d�<!a�V�M��'
���\c��RC�;(
�MC�J�20��i`i@�7�d�� 5T��$�����T)	�A[�*)�ٌ(��g%���5!'�G.]�����S9{_�5ѐɝpPx���K��|�W�[���i�%�\����A֣bՠLA���Y��D��e�l12�J�7ࡸ�H�{H� P�}�"���e�6{d����+޶
���sm�uS���Wƛ)��Eːaڋ?���(���~g��b��5��ЃmwW������(�u+�D�T��`�&j93A�!�I[�@�3 ��.}� E,}]
�j@.b.�0`D�*UxН��MzmJ�Q �-Of�
E��9]�B�F	؜���*Tzҡ����zmH�	�L+/Jl�� ��
�	Ć/̺�34-%13�Pk�-a�NL�rʻEؖuB�#�7#A��jFIE�*���c��ijh��DI���'��X[r��7_���Apʘ)gwzI��a�!IVy��/ ���2��V&L{"$Ե[���	�O��Y&ܕd\���ѿWtY3r��c��e)V�
��K5a�5"���A6K�g_��C�F�Je�E�H,uq���@/�d���T���T�Tq2���\]�(��O�h"U�K�$v���=9��?��p�7��S`�C`C[�2����+BXڬ0�O�8�eis��i� (���L�Ra��[`�[�0�����B�Xެ]w6��L�	iT���@@zD������'��@q`���b]Vx��e�,�X��*L��8�6�H [����Pa�?@6t �'�Hk���5���*�K�cc� �v�� [����< �C�H7FKx��#ǯG[���7I�#S�'y=x�:$�Z�LcU#!D�4�P�GC�,A󤑴C�	cO@�z9b���_$8{̐�C�N IZs)�+9�]��G9���P���0�2��C��=q܌����a�OF�SD�� ���ZUI�Ǔ�^��Q��Z����'y8u�W���Dv�+����VUA�r�N��;?��I�TfZ�k@� ZGi	8��)�%Lm���d��p���г��$�Rf�d��8�)��	�'HS�=���_3LB���Ѣ�V=�%������������k"�Ӑ/Lfty�H�:T�(�X Q"��#Bݬ�AZqG�	��yYdŒ�='���A�>�H
�Zs^�õc!L"�,paOѵ,��h�E�(C`���JV%>�sa΃glLy�2�(_�zm�3� 1�vF�4��,O8�)@L+j[��Z'dB;�� �5*��8��8R"lӆDp�Ar�"u�Н�f<a�U�"�M�\S�R�C�G��@@�Q����hYɔ�@H]#��92�"Q�IMB�La��d�t3t�Ks���@	��U$DBE��0�$q��i����BDR�\�����nE��"q���o*N|h��T=d'V���d�.�����"D�Q�J�cF"(�uG�-{i�m�U��'&�D�@�/V� )�q���%Y�`B2�DP�v9h "1�N|�-���ē$`����K� P�΍)Я9� \*� ��*��up��]�� �,PB��-,��I05�\����Xw���bf�t+�x��Z�lׯIZ\`�`�/v���'�],�rOv����Y���ɋ�	I�إ�����a�˰#�2>��鈹~��!���
1!�7�� �(-Y��{�d��
���$�v��P2W&�����j�,ژ���G�~b_�lk�K�D����dɹ~��R���� ���a�8]L���5��T���%��6.��nZ:[Jʍ)%�я]��A��kﾁ��ݚV�ɰ��[�2&���N�8�M{�(;
IY*רԛEC�����5�\���'v�\����A�U3�U:J
]"��TDF�q��42�@�$1��U
�.Z�rd��	�a�b�����<^�����i��_���z�nW.8���M>q��Ot�	�Zzk�A{�<��@�|�АPE�32%�A'K�,	\��[`	k�B�}�0��O6`C�M�/�1��A<��lY�!�5���z�b0��D}"�̨F�ȱ%J8	>��ˡZo���H��	9Z}�u-�[�����۟r��7��((��Q��VU�O}j����
D���Cg�1h�\��OJ�qO*��W%�
f�N�x�L͝<F� C��{X�p��E RTDxr�;ư��1mi��B��#��ɳ�Դ ��lA��jBj�?̦Ѹ�� m��.+�v,�#g��Q8E�8�r���M��
_�U���SiƲe��ɢĬ!b��Iu��8�x[6�,I�2�E��_^P(�f �?5�
9��д<QЂe�D�i2���ёd�a��E��ZUH"=���)��,�GT�@��������‬ϒ~P���,�ͩ�������ԛC������r� ��6�*%K�V��B�!�T�1��.S�ў�ۂd�C�����EI>]��C�I�$=լ��舺,|d�B0޾�?�m
�����'* ;��+&�:��<|�2U����7��\:�!�4%�d��b'�I�o8�1!��3ֲ��4�ӓ�ʀy���0��Q�MM�� �TO�8�<8�`�]���`��/��L���S�B!Y��;���;�2 � �]��|m�ohT	2����#�(�/��1��!�Q�\["�I�W���n�!�����#K��	�*.��-��A�T�^���*HuB�11%�Bm�������
��`xg$ޓQ>�����/�X����(�9�ykA��G���`t��=/�踣X5� �	D��B�b�Pb�8�}k1�D��� �MF�'��̧M b���	A=u���)C�5"MȠ��b�I��Cw�I�3ǨL����N'h�bF��;NM�Pf�T1��y�PA�`N��ä�`�\�)�*7��ۺ�h���x�H9lV�d����	r��ap���<�T�q�P�tն�I��*���,A��E�W
 ������i㯝~?���]>�y(�Ù~�a�t�Rn���!D+#��#�H��M�b͔T:��u"E�u�!B�$'�X%���r��p�ۉf��9����dL�Ƨ*F剣:OD��aZ^�3�ɼ,x!�r�[�Z0e ��1��ۢ��2*u���� W�XTQC�~��-����?�RB�#��hw�S�b��XP��
�$W^xP!�'{*�b�V�/'4`��_�4��ԉȃ)k�p�sB�7o*��R� CH���"}���'e&9���C^`iiC"To�'���ᵉY�G����`��W�S�t�dz�G�$v=�!�@oT�uBC�I�d�0E�X�e��o�%(O,�;��s�@�f
I�,L�}y��)��i+���6DH�p�������Y�!�DI0�]Xw.��A��H{��S52��7�,y����kf��D��"�̍25i�����	B0vp�g�#�I�"Wa�c�,�;y�������TH<��B�0zhv��"�.1*�6��s�<�DGS2X��yJ�$�)#2��uYD�<1'ؼo�pG�M%� ��bG�<���B�2D�&�-��~�<����=BZ�)@��?�^�7e~�<�-��zhd�@=I��@�g�<aB瀔O����ʱR�>@1FJT�<Y�/T\����戎6/!��T�<� ���H�B�ArTL՛6�,m�F"O��ӆ��dg���vi��g(��"�'���Z5J�o�}A��N 'ߤC	�'�p��D.�T��3o��q�	�'{~�R��Щ�}{rg�<���	�'`�T��6��q,�!�$�	�'�B��p���C��F�8���'y�;�_/�HM ��G�n���'u$R�,¥'� 1$HQ?�����'� 㵊�r 92�c��M�E��I�rxI��R ��a�s�ޗ����M�5���?2��e�����^T��<CR�
���,Qe��͍�\�ȓp����2�)�|��3��FN���%�xP�&x���ؖ��te���ȓ,4ڳ쟅:V��"�*H> >x�ȓv*��:0A���Z�I�"~,��ȓDʲ鱤��kVy)��)4��ȓ>bXI��_�o�x�2C�6[,p�ȓM��p�d� c/&���FA^���a��q
rLP!g���xq�@��х�!"F�bS�&"l����ۗ/D\��+ɠ�;�6I�����+��,�P���\A[�#�|t8����� ��ȓ4$��+��c��PgQ4~M<��+D���˔m�.��BK�;��)K�)D��AA���f!S&�ـw����R�)D���a�eZ����)����a%D�p� $���-���F�}.�� $.D���
ė2?b�`*F�G�~��.D�4�1H�43L Y����`	N�p��/D� 3�(<y��1�F�< ��A�2)D�Db�,���I�g�-	r��8�(���TΏ!8�ru��
@.<����7ړJ�č[aK�kP�;��]���� ^��&E�$zn�1�,�
IM�ȓco�i�n��Gv��%�DW�Ѕȓ,Z���C��]�Д�H��M�ȓRw�,�a�P_�Yj$�[�.��ȓ6���r�"��4��%�$Х�=�ȓJ����'�(���f�-5�^T��rNl]��kU�^XXz���
��I�<Q�'Z<-.Ε�Ňʒ}�L��p�ZB�<I��O�tYB�ێ&,qZ���c�<Y�L�B�v��k��b7D)2�`�<��X.C��q�oω%�V��P��[�<A��١Syl� T���D)�[�<6K8)�9A���4�8�|�<iebO �z�`r�?���kZ�<	"��3CD�I��t�AISh T�<�� I�R�Z�A�B6L��M��EZ�<�u�%5&B�x��R�?W��d	T�<�U�Ѱ" �Ar�[����#c�I�<�E�βd���KFO����1i�H�<����^HLjV!��5,�rD�\�<�q&�~@��C��;2l��"+[N�<�ōҾ
��k���1j`}�Ђ_G�<9�NN�,�&M�g�M�b��T��
B�<�%�;[T��!bI�3�!���A�<A�Ç<P�*�(0fʙU�p�6.A�<2���$��]!lrR����Zy�<� n�[D�<:���~�D�D�j�<����16�r%2$&/zuj�Ln�<�da��;��JTg�6��(%ʀf�<AWaΧC�IF��2=>Du8���Y�<� V�1.�3j�� �hl��P"O^2K�
�h9�p���x��"O��e��L����fB�
 ĘA0�"OZ�00K*
��(���?1�4�S�"Ol8�/A3�����v�AT"O�!�G�A�@_�[�R�/F8�3"O,�QsF[2�@�Ks���f�a"O��a!��.�PG/D�Z�T(�"O%�d��Y�J�QpnKj;�!Q�"O��P�Y�o��(À�&��(�"O���E-~�HP �F���u"Or	X���3n�x����@� ��W&���z<�b�����xꋜ0��3�[���#
Z>��0��y>̅�ɰ'dZ��4φ�,�aUh�88�
�X���ĜR�;F����@iX���f�H�c�dM�Vf�> Y>�R�cʜ-&��8�A�(����J�'��	����b,�&5��I�fk͗I7�ݺ�dt(<1MCV�lx��/�CR�����J"��eGyDj�ѱ���h�H3n^�k	p��e�t`@���&Z�t�j�bFtվ��v�'h �e���Y��T���]�P|��l�kO��� f�-VA���_	j�F`��D	�M�� ��24����Oϑ�Tc�a_ x�x� C��}�b�xӈ7}�I�(Y{�� ���*�>�	 g"���'�
��B��hÆ ��%Ry�����$Kz�²d��"t���'����B�p�b�жl�����3�J�/�0%H�!V+-K���6O���'�JIJ|��O�(S,�1��&�Y���Q���|�6͒0XS�0j���<]�:����a��a��4(�D-}���ba��z�Ox�k��T���G:�(�g}�$Т[&(��b�r�z�FO��,صm2ړ	�t�kË�\9ΐ�ׯ����M"#�ΐHD������K�H^�!̓@<(����ʼz�D��=YPmN���E��!ؠ���Q�?��q�t�'B��(�O:�2�#���
�Vt�0������{?t`8�ʁ@\`�1F\�jް,[�`:��'ؖ,x��e@!fc�	pbU�O^�`%�+��)�㭊�0���:��(�0�`4��}^�Y��z��"�Oȳҝ?��L<wp�-�R��#�nX���C#c���3�oˠo�9rv旗kP.p"�]^�'���y�'͸i ������4V@�-C����y��>Al�g�ȼGxr��sr¬�1h��Y�>�)`��-<�60���3]FY���I��
Y�v��M��8CDƢ�2���'K�D�򣢃��0rv"�?��#<�wG^�V��m��
&v�AF�ȫLpk�Q�t~�	����^��-��h��<��=.\����s�&�P�ߍzar����p:�O��jfH	�C�h�O���}cU�O�=���\�|p��O�5��(�@�~h�	_�R|�\�'��������E� p�s	�81���
.7X� F wp`�:���v���'��Û���W�,t2څ �r��p+��l���/҂�"lbC��F`���Fy�'e�� 3dƢ PS����Y; f,�>���:]H��Gx"H9�����h�����������\�|�����"xaD�;�M�A� 3�F_kh�: ʖ�3Jȴ�c���8Z|��i�@�̓2p|0�pF�K߬���mo��m��>�j��Z;k솆���Re9[�̘
���6?i�26J�s�,B�)����4�΀֪M!�'�2T��/�-M���:����Z�2	�aF��^*�������5,�"ntXlZ'qh]�q聣5�d@˜,O��u�X�@�5���U��ı@�s�P�Y�%��YZaD\<K� E;�U|���IƮz��$r�F��e[����� �x��+H 3�82��yf>1J�蝕=��=	�\�QgF��0	��p��H�s
 E��Fy���?A�JK:fb4�y� Htz�z��<�c��S:τ-(A�_m�H��tɃX�'�X����!�J��O� Rl(\8�lֳQ!4��5,\��h���x��O����J"r��x��؎#�=�¸�
�&ĂQN9�1s^~����7��H��|���O|<�v/�-hx�$�c�ۯ{6�A��'�:6�b����;_D\Q!�@V,UȀ!�%יn������צ��%�{��1�XґC�>u(�#�Tk$Ϋ?cr��R��5*^�R��7.�1 {|A�}��|z�<.4ȕ4�1K�2���ҳHV�M{>8�'RN�<� h��hO��`G���&���1RE?�>�	%)�`D�ik�<c�P�O�	'@Բg�B�"�C��"
ڙ�6�R'lg�(˳�T�T�>�%���+�.�=��˹fJ�(�!��OCp(���Z��h�QB'b�x��k��h���'���Yp$����I;z`��4z���K4������,Y8I��dw:|RAo�o��uI�u���Π� q���Kɧ�4Ǟ�\�p�Y�k?T0z�$�1��(�A%^C抵�v�i��sB�O���I��M�2W~�"pX^}ҎL5'��Qb��."#��b�IҬ
-HUpVc	F� � 6Z��!WŹ|&���b̎�x��!�H�R<���U����q��?U�,Ð#ԑJGL�tǟ{�'n\�"r��*Np�!�CT�w��ܪê
6"_���e �B�D4zca;���5b�*p�Ӕ_}Hu���
7U֠ ���}�bHU���ڵx�K"0Ȏ�=9rIG�|�t(G�Ƅ2�N�]�@�n͠ �/G0�u�Sf8H����<1�� ����rᎲ?q�S�v�0��O
%��#":���J!�*��$ɴ�Q'����
ed��* ~;���)�@�%˰���
s��
ag[%@�~W�0aRI� �ͳ9�R���	Q��Mӂ&M�:�o@({�* H��'m���8|r,H�̞(8��u	��ԚF<�l�E+߰ E���� O�ds܍(F��$x�r-�O݂�1��i�Ћ5� d�·�H(WY��@F�$-.ajvG�*8㞥0M�- \<a�f��"�t�D{��v9�ҳ��*1��%�f$ǈ	��y#G�=sz�S�O)�b�ؐo�5�y���zܧ<J�Up��Yd� ��4)�*�K'c��DB���  �D9�A�.��d���c��xrײvoz!AA�FM� ���_�#O�I$�4��O�ӧ�4˃�D�h-�jǤ� ,*�[�e�t�U�>YR·|��5��!�R��0��-p\ɵ$��q#J��Z�.��QG,�.x"p�\�U@���O`�'���ҩ_����U�B��[�OҰ%B�d���!ʖN�D�1"�q�2���D�>j��M����3&�Q��ӧh�!;.Oj$������n��cY^�k�i��@�e��]Uڌ�p$�+8-b�J��$хU�ܺt�S7['r�+eK_4��=1��ýk��u��*F�>�dA��!�ɋX�Z����OB�d#*;p5	7'T�8��������0��Gs�'MB�
�(��^�� !���˼K2F��J*�i҅�I�vT�Ă���<��Z���,�,b>��O����"��ul%S`ǁ7OWzX�#h�u��^.���K� L+�0Ӧ��$��9���Z/���`>1ZdlW�?� �1�0y��rd�Ov���Xs�	�o �<Y ��K�a
$�U�] fQ�߫e����� ZT�f�5�x�[��p��'���M���qlN�Ps��)kM6uW����m8:�D�Ɗh\�2��L���6��+a��y��N%b��O^�}��dK:)s��B�ޚ�L
t����K7)�T	*��$ȍ~��p�#Ŕ��$���T�C�*�4`,B�1��� ���c�<��O@��'�T�ӵi!����?�I}�~�sb�J�4$�oКJ��'��K�	ƐU��H�Cݏ7�,\���СD��X�H��|bQ�R2vi�t
L�6m�E�Cݟ$a��[ןPðbÖ�ay�D]P]�T�oU%\�"�����N���ӹi������H�?��\����x 峟t�p�Op�Q0iN;xc�0�@*�=�����|H<¢��je��M,j�j�%8a�:9z��F֟�������Oby��`z�e�w�h�+4�S�B�Q�B��Y��'ph�)`��Ϥ�Q��ԋk�p�����y�D��'���%�H�SDS�t9��OE�uD16̏w�a����{�'��"����+�eJ'o��QO�|Ĕ���Jخ��P�d�P�a\������@�!ܤ|�CD	//,����	����-m���c � )��Y��]������`�U�cm�H�P�_�ӧ��t��M�Y�����ά_@x�aId&�.N�D��Do�K� =˴�'�ZdX ED�?ਰ��GX2{��Yy�U�E�D���k���(O�)_�y�2��Ī� ��ӓ�!���C�'{�Μ�9�R	PfV*:�� T��F�"U�����<���"P��/F�̨���֦'��a���4|E&�IУ���џ� ��R�CR���.Q�b�~������p�B�oN�$��u��J���0��E|�%Kf ��<��A6��K���t�ݘr��D��1�E�FFPn��[���@�;zf����(
h�S��<�T�S	ԅC*�5}��D���;�M3f"��0�BĹ��M�h�"�r�L��UcrDI�Ĕңe��a;2q�pN��D��UR����՟�)뗈�xܧ_���ɵ���-�||X��/�����a�~��`{a�[(��M�GG.jW�
!g�����+*���yp��6ŨQv�J1M޼�&����i�'L��������~����5vQ��S_�<`���L�~�j�+�~Zw-$<���A>��M#�-�����Jғ�5�!�2\�i���h��$%�"%x1n��m0^$��G�64��Q��'B�Wc�h��O����O�#�@�(�A�: 8L��.�3�?�Ɛ�Q�D���Dh8Q�%��]��� þ|뗎�1~�R��ȅ�~��K�4���i>ax6א��$�߱����q ̘�m��&Q���N"G�.Xדe���Q��a�Q�pK�h��DC1�IZ���S�%�>��.
�i�2���4%��Q�tC�1���'���'2N�����Kl�9q@U�zh>�Ey��S:r�N����fy���<�DO]�D�t	͛=���I���ʦ�ɓ��n��x�o��?Y%�.�g?�ÊVu�k�eGr0HîEQ����iE|1|�'�Dҧ���i���NOf��N�=f�ic�n�O����l<`h��aR`�o����\��I�n����ʆtU2� }�<��v��lP�؟�mJS�9c�y{�EŅ&��#@(��:g|�pm��w��z��96]�6 �6ŋ������I��p�t1"�V�Z �����lu�0l�a��|��%8�� �c;V�Z�RbƥҢ<yt)7e���Of]�'V�� a
;':�y�����yy�h%$���V�@*c��Q�d�@�)1t�9ڛV�P
#7qO�}��=�q�k���8����~�A�rΟ+� Q��'�v�a�DU�d�Ձ�U"z"Vt�'�J�	�n{���ø�^��q���y�.�xs�f[�9T�%�ò�y���. J2��&ER09��!%�7�y"�ζB"!�s�[0��d⇀M�y⊂��H ��.^#��E1 ��yB��(?�T-ZeE�+�ܩHsH���y
� �y��CL(��!�G,�xXp4"O8�i�-�$R�B��R^h��"OFq�e��>2�h�TZLFG"O����S�e��C����v�J�e"O�{Q`�;��D��/���%XC"O��Hu
�g^�	Pɇ	~�b)"OvP:�e�<X����\�?���W"O� q�E-s)��i$�˽z �P:�"OxpPr�N�&�)P�(�+^��H2"O@t��f�	������4;¬��"O0�㤟�Jծ�+-��@4f��"O�����"B86����S0p2�Y�"O��Q�H�=#JL�*�̻"O� �UG�>Y#����_!:���x�"Of��h�Z�Dm�+ϱ%�||�"O��xt$ł:~�5���H,D1�H�"OL���"�$x�|p�,��3&`���"OL����8C�P�@@E�>A.��"O����(�$������$�D}�"OX�!2	�Ui�Q��D�Gy��RP"OjPp���4s]�(xӉ�_A�1�"Ov��S�F/�\�8T	F�#�љ�"O੹s�U4%N�ᗇR�6ט�Q"O:ՠ5�C��l��&U�u�V�i�"O��3��l�<�3g���m�"O6�K��E�>rڤ���	�J�Lً&"OJYXP�˰b�0�Hs��_��h
�"O4A �o�3k�)
���$`�h�W"OX;1'Z�'h�&�68��A�u"Oh}p��)d,0�C���:YS��c�"O`$8�&K�oH*\�w��/p7��*O|�pr(%5m�dyb���� �'�y�5"?~�a3�EI�ܚ�'L�3�/^�l(`��V�Y�R��0�'\�M9���I"<8S�	�LY�<��'Q$Hp�)�%mr�xC�_�<AF��	�'S,�h���C>%���"ƀ��
�'Nx��f��SB�肠�m$u�	�'!����l#�����-ZMR
�'�0"F� ��X逇R0}���	�'�n�Ι�K����WmA�i��i	�'	��	ЕRV�%�w(ϒ MFe��'���+��� |z�vDܔs�*�R�'��!��ƏDv܀��Lh�y
�'jm�ǈ^��azF��e� ѩ�'F�m�#��U8�6IڃS��u��'�Ę���)ll��Eː�W풍�'���Q +!F�Z��� `J$s�'�ZeKvi�2	yd�S�_� ����'b�Ȱ�iJ<m�&P�V�O�p�ҥ)�'A@@{��� �2u��j�Z�
�'�(1j�(���t�!
ȑ�	�'��M�AgP3� ���D~�x���'JX�sv�]	w�%9a@�n��,3	�'���3�<[$P�$���p�hR�'�����E�T�>��aW�4f��'aX���(Q'�>�C��)! �#	�'ڤ�P�R�H�@ؤ)�#i�~�<QRi_0u���@�T����r%IC�<�d#�;h$x�dR�a0��2S���<qW'�>;_"��Eޚ�氡`�H�<)���Kwz ��o$��Bb�M{�<Y�
4Y����2���3��1S��v�<���]7t�6��`�B�mp��
�s�<� ��Y��{)��`�BĖr�n���"O�� a4W�0����H�	�^���"O�Xö��]���Жm�0{� j�"OH����\�n��u:��&J��A�&"OL(�ʇ�gU�Ac��Y�t|�T"Od���K'��`�Qh^93$"O������a��-d?&��E,�
�!���hEV`�%���#�1��K�!"�!�dG?/l�	���>(���	S�8l�!��8�X��@�O4�\���']�!��I/��D�q�2k�\�5��"V�!��8 ���vͽ[�!��(��b!���,\h�`�%5�潛 N��!�N �PԸ�h l~��C�쓥
�!�$���=e�E3 �����Oe�<�ލdf0PWm��z�1�Z�<	U�V6l�¦���<���`��U�<�EeI���	6�%P�� ��H�k�<)0K��P�ԁc��%���P F`�<��o T ����T�9S�� @^�<Y��ؾ��V��p"p�j\V�<�R�Mjw���IA.� Yqa'�Y�<Q���?N��+@���gK� ��N[}�<ف Vgm�;��A>s� !�,|�<���ʢ4�����_6y��P7MLx�<!Ӣ
�w�Ra��g@1K��8�C�O�<�t�J-o�8�Y+6�J�C�<)�{�ec�ޛ�Q*�EDu�<�c��%?�a�d�C�,z�gW�<�U�ݺB����l��+r\<GT�<	UI�?w�PP�ϛ���RR�<�7m�����D�{�1pW�Rv�<�@ن
x0����
d���r.N�<s�&G�@TKT 2a�5�DD�C�<�w`J���5P@F�Rh(�Ca}�<���Ep����B[ 1�PR��x�<�c�T�B�ΨUOێ�:���"Dx�<A�������0�&8`eϒ_�<�M]�	p���lN�A	�e�a���<�mV�WC<`��2-ߤ��7��x�<A�A]�+�̸To��8먥�Cw�<iV�
�F���G�ٚC�`iUoh�<��@�T~��$&V.2E�}�qz�<�1. O���!�����!bDu�<�!M�7BJD��B�(ےfO�Y�<)s�H�E�Wj߸6an���Y�<��X8��+e�J�Gb8�+QO�W�<����}A�,�:(��}�$�{�<A�)O)��:���
,f��4�`�<�`@V5 �ɒ5+Z\3HȲ�p�<��ʶN�,�z�K�I%@�����o�<y����w�V|�`K�F���"c��B�<�#�� D��bA	˵(��p�V�C�<��T����d���Kq��V�<)�w�Q3�B��CI��, ���_F����V#PTx��T``��ss�%Z�ć�u�,�;��1*�:��Z�.�#T�P$+5���2��m��ȓ
i3��۱-U25���
�2U�ȓ�08�-�!���GH^-4X��!S�,PE 7�^��������{�I�����I��Y��/ޒy����w7�y�Ù.c����&�@���ȓ`�T04*�<&��'�[L�d��S�? H
�*W7{!F�aa�T���""O���%�-6�B\� � N�P�d"O�!HFٳbt���cB|lN���"OL(!�a^-��]�ab�Ox��"O�!p�d�8�
� �ߋIV�Ap"ON�ؐ��-E�2� ��Nu*���"O�i0�0�0,���ڷ�j�`�"O8��)��G�
��a��;[����"O��C2��YJj��d�^�)J U�"O%��m��2��X1�_36���P"ON��`C)~VJ��e)��b�"O����m̫aHv��5�H�Jl�!�"O���c��	
�J���a�?���6O����Hu�J�"�JV%!^H-�� �@��|��x� �6LޜPӧG4HY#4��;�y�	"~:4����8�`a��
��y�D�6�8��C��z���2��y(@�!]���6�t$`������y�ۺb/�l��D��k^�Y7n�3�y��H��{2��b���6����y��^3��)�>0d� %���y��ݶte���1��=U@,2����y	��[U�� �E�;L�0q@cڍ�y��GPoPx��!��D?�t� Q��yB�7o��|#@f�p$��<�y�@@�}�JЀTeP.Z��P�����y2-C�g�	�CÂ�!u�UYuȼ�y2h�<a��d��"���F���y�J�<V��1J��q�@�b�yR,O�>���k��6Μ�"�Ί��y��_��HSjԤS�-2S�(�y��ݏ]3��q�u��e�Q���yr헚/��b�,�p'��3�]<�y�!\*r(��"�hEu���-Y��ȓM6�Ӏ��nT��z��8P�2��u�B-Bɀ((�N9�jǵ:�����j,bTA�O1@ZI
�2��G�<�"E�oT�jvi@�Bmɘ"�@�<�d��
:-���lЕ@�T`T�z�<���ōG�1#�8�0��7f^�<qR�B�5�,r�'E�$��[@ǆt�<Q�h�8*�t�f��P9l�3C]w�<����j����u��2����@�p�<&��yd��YY�2|j/Vp�<��Y�`�UR�#���;�Ti�<�Q�E��p�
â� 9 N�f�<����L����Ș�y�u(�eCK�<�"�<���j�%F�PE�"h�J�<)sg��J	�a�&Š�I��,!��7���s&��Y�`D�� ٝ=�!�d�i��Q��e�@{����
$`�!�Ď/X]|�a1HĘgH4E1���)v�!�d��I't"c�B�h/���*��!��N��x�  `'�hx��W�!���l�t��l�1X
���KA�i�!�׃Sx�Q{C�U�
 T0�Jn�!��v+�3� c���A�@�!���l�t!v�^�X{��!����J�!�$ޔT��30�[s�9RvM�w�!���-hBmy��	6�^�so]F�!��Pb�$@f
IB�h`�+h�!�� ��q���W�0�EL-�!���]���x���uq���<n!�d���zU��	�	&��Ңd!�� �D9�� O�I���T�/�����"Of$kC��*<�Fx�	�C*bH�&"O�X��0����#)���(�K7"O s!�լ0F�q�E�P3kIxt�&"O��@^�Z��YYP� jD���"O�����h�7��(7�-�4"O.���H��`��m�a�V"O� ���2؆HJԌ�&�j`Q�"O�,����Q��c�j0b�F\h�"O�AK���>fX�i�'(��A)�"OL!���(>8��v'� /k�G"O�\c@F҃l��X�s�uU*�I�"OF<�WG�>)��+�
�#I ų�"O���Qn�23�!X��y=�嘷"OvtJT���{�m����<~�,d��"O.E���㤽i�-оh�d]Z2"Ov����&NE����+	�=�Z=�"O�	ᑤ؂[::���jW3{��8��"O�1H�_�^BUb)B�n4 ӓ"O�$�c�D�x�H���p��#"O��Af�G+:"�����< k�"Ot���ĀP߂��l�>N���X�"O:�*A
��|��#3�
(�"O������ia��K!��(��"OP���ʌR�$��j�f��Ag"O�l�!��:m�@]����q���p%"OX���J�n�8�c�j� NZ�9�0"Oȝ����'�ȵ�b(�&h��Q��"O m����{��(���� ��YH"OK���J���J�C+x��1��-�y�R�9�n!�o�33����N	�yRZ h�ڍ���>[(���PL ��yr��B�4�顉�<Na�f�y�)��r�'ǎ�1��|�l��yR!�!+�l��Ā�5�� � ���y�kԜ|sl�� �C8�|=�͏��y���a
��BB�J
��a�5�R�y���U��Ѐ�*��.��l��y"��o T�� M"d%ʤ��&�y���acf��Q���D�PH{S�$�yB�@R�zH�����:�����@��yҢ��S���3��D�E->�1�F���y�m^�Xn��vm$>��=p&���yBI[�Fw��2Ri�<M&	:���yRnߖ#�z5��6n�+�nȎ�y2�?��`���[�dXW���y���?&h)H� E.b������y*�g�]	P"ٖU�l�V�F��y����Yq��E7T�dy�����y�&��B�+�^�4I��<�I2�'-�y�cG�~��*4C��8�ֹ
�'�P%�#,_"	P]�#�W)5�
�'Ѷ!0���~��(��Y�6K^)q�'L�b�._0hq��]�< H8A�'��T�to� 8֔��*�?+�ٙ�'�ܹ���P~T����O��e�$0
�'�f��̠G܀jc�M�)!p��	�'Y�1p@��~xq/"�����'��|�3FL�}��,P!��-NNI��'b`́��O9J��9oņ$C��K�'`$��|��$�3��H��'�b��˜t7zͲ�iV��Е�'8�$��0ez�D��ru��'}4(�dBA;
&���S�M�O�1��� �eq���\"�P�����r��Q"O*0j$FX!M~�)"#�zyT%��"O�Q��AJ�ԫ���;{U���"O��[��>�@�Cj�fg�P�0"O<ȓ�a��G7L�!��������"O<��V�
}D���a�"Q"O�m��Ѧ
�K@�K;c��� �"O��Z �7]^�!0�Ǹm�5I&"O��P�H�'�E���'n�fh0S"OJ����>�6��#��<�zݢR"O��7�V\��tТ���&X��# D�Л��C��v� ��77�m�<D�4I���&;.y3�̆3lZq &:D�����W�l�r��ɉ��0��%D��Y�� �Q�8���kG(���9d�"D�؛g١c�@�U�DXH=D��㒏���xP[��V�2�p��h0D��y�S
nOȠk�E��8�a�*O���NҀg4�P���]*Ą��"O����N�8	j�q��C�""O�<q�D t�&} �nL�9��"O��0D�T=U�ؐ��d:M9�"O\�Wk  ��x ��I�|�Mc"OܐȱjU�60�(��M�H��\`"OܵV� 
�,�h�
ҩ%��"O��p�@����#�C�h�ڰ�'u�`�w�8r�<��̆J	��0D�0JK�f�1b��Q��P�e-D�<�VeG�la���&bZ$���>D�T��F{��Z���7K��YJ��:��0|�c��"��li`͌�W dL���X�<�t�J(O����"Ű.���E-^h�'��y�B�R�8����'L ��7+ �yb(�A�=K�@FHQ^�3���?�y�Ɲ(��m�+
�j�ժv�yҌӕr20M�S��$^�9�6JH��y2�����S�#�a^�x��>�y"D	����3�gѺ��(��y�`[J�N���|b"u���ه�y������K9sK�`A��y2	M",���;��Sǰ�1a��'�y�A���50�ؓi�[ʎ%��OԢ1I�JDx��3+\�a9�4�UALt�<��ضZ�n�@��[/2�h���{�<Yq �A��:=V��f��0j��ȓ@z���,)����I�V��i�O��=���,Ԍ��"�͙,]���:��i�<AhH4"�~!J��,}(Jy:��	q�<Y�
����l�0��vp0�Ӄ��Th<1`�(r �r��R��L��hG�##�pG{���i��%Cu�.8�TĹ���)����L2�S��:�		?O�ա��'�}Ip�Μ<u~C�I6T\*�k��]SX�����4�dc����	2iED-B���P������KB�	��MSJȳ}@
�33�C<M�2
H�<��	��0�R���1=�4��%Sm8�xGz"(�(^ Z�H ��^A<8TjN#�yr��f��	YR�c0����j\�y2�H�rx0�� :�D����П�yb�6M�Y�o�[��]����M�'��O���=�I+t���R�LE'fL��R��l6FB�I;,z�B�	��z����0
�*xjC䉧1O�H�R	�HB�;1�H�XC�NN�M��P	0~�1sk�<lC�)� X��ĭ� b�}�� 5)ND��"O��	�7O��9�Ɏ�s	vܑp"O1�!Z�D�7KJ^ �"O��3��k��������&��Т"O�)�ᬒ�^�8=8�I)�$e�"O�q��27➡�F�/f��̨"O����J�>ZF^l@�*y����G"O��k��۫}0~[�+�t%�u"OjP�@�N4S��h�BLah	�"O@�ؔJX7\�r`9"L�~Rl�4�ı<ɏ�����R����qk��ӹ7D�4"Ox��R�q�A��v=t�'"OFh� ��ww��Y�!X�s�D�W"Oz��ML�vL��c@�7q���"O��a `�4��\mD�#"Op]��E\�v�~��vD�ZD�3"O��C`���=�t�JD��LW��q�"O֑8Gk��F����^OZ�W�'�!�dն���Z��M�P�0ujG�Z�(�V�F{���'��x��͹FVެ�e� At���'�N@`dD�It�TiRR~E��'��]�4�

���Μ�]f���0�0?E���sT��Q��8��\с�N��C剌5�v @�K^[��!�t��a��B�	� 覽"�*)8Pp<`N�f���d/��GA�@ԅ��%<9A�� g"O �z���b�����$etM��'����G�U��1h6�2��mj�d&D�(��g��U�>y&"M>X��U���%��)�S�L�z���k�7{:��K���5%��y��d�J����U�H]�d��5�����1Xv��נ-�;��9N�чȓ"Z��xlT<2A�XI1BĸL$��ȓ�xT*���;4i�0Mc����V���4CN�b���!h�&�̉Y���s����U�#좉p�.F)Q���C��.D�D�B'��K�J���o��N�����a�p��I�>QT�� J5�$�*�
����C��U\�	C�E�(^T,$�s%�2z�C�I���	���(B��b��͜-��'Da}�O]] �W�w��p����yb��,X<J�jd�ߖh������y� P@q��Kԟ/D6p�A���y�B7?~�1`c%%%Ɣ@a���y2n���@��/�i`�D��y�%�!,%	��V�p�)�d�˔�y���>Rg���p(βe���A��_�yr�I�\�i��)k�\1H���ybE��N�,pZw�3o欰�����y���R�XY��"l4��CmA��yb�N
Rٺ��8`�t�{��	�yBJ [�|Qg��O�q�q-�1�y��5�x�EC
*s�D���&&�y�@B�RޒT��	n=�Ñ�&�y�Gֈ���"�	��h�hijA��y"��;#8u���Z� ���kܦ�y�K(�$1��!S>�p2�ڃ��d$�S�Ol��ر��?��u,Y���q	�'��ب��L�gC����'.�k�'�F<�A ٧%��hFI�*�<U��' ���iC3\�,�uǘ��,u{�'@�hj�*E���b*�$<R$�C�'-��KaM%r�M�B�L�&^�P�'�^@s!E���$��,O:'WơH��� xңA)f$�C�<l��T�"Oj�Z��J�C��Z�n�`��"O⑚1�3�:A�/�QU�R�"O�H�J -M!�8�a��S��u"O� �1�$=��^V:%��"O���q��cq
 ���X�]���r"O�x��a��h�4�ZT,Ҡ����4"O�1���6Rm� y4, )V���u"O@� �בP��0��D�3}�)H3"O0�Dµo�8I TBC!k���"Oք�Ĭ����B�`�TK��h$"O��2@�M|�ɢ�OαK��!#"Oly��Q
��@�CNP�e�%+p"OV5(W�A��C�X�q�Uy�"Opx(�aX�.�~z�?W �e"O踐��\[��pǍނeI�\�!"O� a3�V�@���1E��b�"O�1ǭ\Q�fm�#�lx@k"O� `ЏʤC�����
L���"O6�"u�$9���A�M9�"O�ʗ��>T��I`��ə\�dm�"O�T��$/���ö�7�4ـ"OD2�6\����%ۑEk����"O�m�a͢@WDŃ�d�+_W�9�D"OX{��l�����ZV��mIB"O$�	R�_�Lv�d�v�L���*O8�a$)ڞ��g�*<����'�J���9ee�0��;FL ��'"�|k!B�J�0q�U!ێ4��%B�'y�А3k��2��� �%;,ܘ
�'��=A�n�'N@��E,���'И1�e�T�K3��PBG�\���'�\�;�h��LIx��R'�1j2���'���B�.�
vZx�!D?)L�	3�'*�@��E~n�����"P=��'"��g���j���)���^�
�'H����;��b,@�'����Q(+U�+��:�p��
�'ȆUI��\�L�NT;�aQ	��� �'�\�2��O2L�-��Hz(P�2�'	&�"�5�0���*vؚ� �'�X4xf�/e���G��|�h��'�x �'I�u����4q�.��'�\�鶡��)z�
���nt9��']�y�D� !_��ivG��f� 
�' @Գ�	�,�덂^yx�H	�' ���g��Rr&�%]����'���ʅ�S"������	5piY�'��u���J51;t��'�3f2�J�'���q�ںq�� ���*.�����'5de!���0"4X!B�09g I�
�'bT�y���W�jqRQ��4�U��'�D]B�خ�i��0 R���'��Bh#��	b�/�z����'_0�@�.O�B�hE����{Ś�'��5�CJZ�!��C��G�xyz�'V1S���U�&$FB8WR�	x�'Ķ�����&_���b�چ^���'�~4K���p���'�u�p�'>����ơ%e��T�U
2.�'����/$�.-IT t�؀B�'��Y�4\z����!�jUI	�'^xD�����8L�B�i��4���':`�x��ѓ&q����JT|���z��� �%�������:$kQ:�<��"O�1�b���Y��9c�
T����e"O�\Q��گH*B�{(�9}�"��"Ot5�jxt�9�1m��R�(�"O�D��	�\�v��C�e�V�Q�"Oxō�=E�Rl��,��9�"O*a�5�N�f�̦._pXK�"OZx,�m�r"G<e��%"��J$[t!�d��t�%�6'XE�؉i����!����b���k�"�*"�å=<!�@S7�As���&�l횴H�&c!�dU���	���T}��W�#G�!��"�pE��h�9XZ8˳ˊ�W�!��:X�Xf�ȷKP��M�*�!��/T��I	��0X( �`�c�!�dݏ"����*އ�|�z�.x�!�]� �x(0 M�3��a���}�!�$B�pAv��r�S�^Ҳ$Y-,�!�d�wV���'�>�r��')�!�d�/��Ya%��=ڒ@�i�!��ڐ
˴��c+,/��%`d��,E�!��4�8�e��9��(9��	Qz!�D�Z���{�	����J,���'��\XB� �87r���%F-���1
�'�Zu���эG��:���:p�UI	�'���Ry5�x��
�4 �'Άe��$.%�0L)�-8|PL��'*�s �ҽU�:�� -�8i����'��|�U��?�؄�p�öh��ݚ�'��šp*�7�Z=���ݨdc���'��c�BJ�kD�+ �Ϡjhʌ�
�'��a���O�<���#�a�`�	�'t��z
��9���k@*`���	�'�9��$�l"�2�ʝ�	#
,Y�'��X2ѭĒ9l��%G�#Xy
�'d��C��cT�E�Ȟ�9�xXa�'��p�y���q�eP(6<�Ix�'Z`(˔hV-
��A����d,��'��U�h��MTXۡ�P�zx|��'`@�Bgƕ�l<�AT�ˮh4Y8�'���S	�9tf���ϧÌ�`�'H�����4�4�k�KG:��	�'�xQ���?1"�u(#��:�J��
�'_4����#F>r�ÑM�;	�z���\g�a�P���i��#��u�ȓ&������=���`��*d�5��'2�Bu�U����p�!��5#6Ѕ�E�&����f'�\p��6ȅ�w:� ���\ݻ��B�D �l�ȓv��!�gȌ-ۜ49� L
v�(Q���2%�k-n�MYd��;� ��ȓ?: �ѩ!�����B>w���U���*K�a7:T����hx�ȓ]���R��F&:V�H6(�F��ȓ}mɰ -��t��8PQ�&g����`XA��1���ۢ��,iA�ȓF�,Z��-�U���A�$<�ȓG���Br ��SP,���
������`~"u�`fHE�⑹��δ)8���dƶPp�̒�R@4����S�~��ȓ:��<3�]=n<b��H�-!�nH�ȓ%vt��G���j�Du�%��g�r��U4�����N��'��me�!�ȓ7Ҥa �H�l��-ߧV�����S�? j�����'�i��@�<�b�[E"O^,���'V3Z��cFB�7�V�"�"O
 ��I�9��8c%�X�� "O ��Lm��4���Z%.Z���"O�͈���',ёǃw��m{B"O���1n!f�z�vA !Ÿ��"O<��F$��B��@�9U�d�W"Ox�i�h��"��\B��J�M:��"O�傔P����/PF�P"O8AIZ�&O6�%@ ��Mi0"Or�!�l�p�����Ә�npH6"OL4���"#�pd���(H�i��"O̜�@g��j
R\ㄆS�>G�%H&"O �	��
$0�F僙^Z���U"O��C�<��w��V��iz2"Oykf��-!�D8�5C��z(�e"O ��4��v���va�b�:퉂"OuB1�͡!R������pc�8@�"O�	PA��h � ���H%b p�"O�#��B(v@��̙�E�E�7"O�q#s � ��S��s@�kE"Oe;��%�(@ʓږbl�Q"O]�Sʕ!�ZD	��]2�YQ�"O�t���\"
����NWqj�k�'! 8B�(��R��X&�4i	�')<�Q���'�.�'!$z��',�K��a�s�̅���R
�'�]�p��� X0GK����y
�'V�T��\�Z��É���H�'��bF.Nъ6l�f�5��'a�$�r�K(~BLɄH��g?���
�'n
=P�"�=�B����ܓP�Xl��'����EMf����tf�A_jP3
�'�Hm��Dߠ`�6�۲)V*t��"OĹ�A�۵��Pf�99���T"O�آG��=�hrQI��Qe��"O� �
�iH�`���QG�e#""O�VY�W`��jBd��p`��2Ï^�<!��ܤI��5낁��%�rx�gO_Y�<��KF�Mvȣ���|/hh����R�<���A
M�$!t��Ki����W�<�R���"i���R�k��u�焝S�<q�c�M�v8��ԭ:&�j�S�<���q�ڠ�r�C��#e�y _����'�f�r�9b�\�y��� ��Z�[�XSRaߑ�yҬ����Sn�6��X!'�A��y��E!l��`Oi��6�L��y��|r�5��_�e/�� vbQ��y��	�3OD��C�]^m+5Aڴ�y2��4M 9�e%�?lv�4�� �y�'T�a �FN&2r�a������y�d�-|;�X��ȃ*N��i���(�y��)xnH��:z�"c+T��yB��_�v�� �|HF��"ME��y��O �Is�����6%��y���d@��d�v��ICfi�;�y���*�.����"9K�|��
��y.� :��B�ݛ,"��e���y�">4&�H f��X��ͣ�dG-�y�<k�~#VG��g*f	qC#M�yB!T�v�\|x&�f���%ؙ�y�ÊG�A��j�`6��8ry>B䉹���)�F��H@�G(J�c�nC�)� f��$��&�(
g�J�$%�RQ"O>!��U�����P�X���""O�,hQ"s���7���f�@�"O��b���>0�@bt����%"O��듇Q�?ٮ�Z��6<����0"ONh8N�1k�P�ч!A��P�"O�;��Ɍ'���#�#� "O��;M>W��躁A)��i��"O��q5�hc���S�D5X���3W"OT��K������d��v"O�Y���>b�	juEʠ}���!"O���a\�n�A��
9�،��"O�`�E�{�����;��lP"O�y�e��|)�%1%�E���x�"O�阖/G��r�
Fc�@�RbW"O~�)���2��a��)0�t"OLApqM�������D�y��Z�"O�Qy�A�8��,AF�̠ ��8�"O`,iU���e�$��S��	�T��"Od�Ɉ:�\ؗ�F+� ��C"O�qsCH?QB��Ǧ�(�j�JW"O�%�d�O�n:��%
8T�>��c"O>$Q炤��<
��	>X"O�e�ՄC$5�,R����>A y�t"OF�Y���dj^(�2�\6��� "O�բP�Z�_-Ƥ:afT��I��"O����*}nzg�=(��\B"O�	��˴8��}jE�݋t��"O�j��p	�8v зg�<Ò"O@�������L%Z�d�Vr�SP"O�����й�!a��z�iQ�"O�鸱��%����->ޞ�p "O�G+�0=�>��C���@�0�U"O�(F���c����ҫ}���"O:\(���1 n�9[�+[3[�<��q"OR=��f�1�iauL1=�v�R�"O>�P$��4Z�*�΀k"O�d����%-d��&��uSTp�P"O���,��FTr���+\�
k�a�"OJ��Sm������&�@�S=�D"O��{g�K+!xH���,�(pc"O�qʓ�^&&6�ܨ��p
uA�"O 2�5�hQ4��? "�"O����"�h��)�PH�3RX!Ȕ"O� ��T�	�x���a�;��dY�"O0�*�"�S��t��Š(�8z�"O~�j�o�-] .�h&�%t��4�D"O���'���
<h��"B����"O6���`�*Y2��J2vG4�ӗ"O �
VIX���#��o*r	��"O����ό�3 ,i"#ɢ-�Fɹ�"O�Udh�hpI��`�����"O`D�^
<y���&�| �ڵ�yR�hF�ᑈ � ��&�*�y�j��
P6�r�	���u�r�>�y��>��t��)�|�&�y�fG j�Rȳ�
"�B�k���y��� ht Ӌ�S�r@*����y�.[Zɶ�gi�&a 5�����y2fXܒף�5/�֡�R��1�y�`�E�^Ո�iގ*V������y��Ț/Ϣ�SfH��)���v�â�yB�X.g�@�A&�1ԴiG�y"@��"v��Dc���\����_�y
� Ё��B����;� _}�
��&"O������:�	�s�X
>�����"Oڐ��)��)"M��ї �0*!"O$1F)�]��=#5(�(7��A��"O
h!6�Z]�B�3M�LD�@"O�$�TmBz���Q3,P��0"OP�	��\�Q��L�&�{���"O�Yk� �W�0щ��eBAs$"O��z���!n��`�_A�f�
�"O~|�� A7q7��HfL_�.��:�"O��X�ę%��� 6��
o�J�"Ol�Cf1��|�bEX[B���"Ob�a�#�7� 50a#]�L@��"O�4`���n�HqXç�$����"O� ����h1v�!��ss�8�A"O� J�$
<�� ��U�"W��H�"OJ�ql؋V�"��F,T��r�"O�d�"ZA���e�扸�"OA��$�
�3VI]:?�4��"O�stcC�g,�тH1=��h�"O�q����!?pa{aAD�^vPh��"On<I��^1
az��̀��)c"O`�b�ŝq��S�%W	%�*��""O��jЁV�c�Z]�e^�n�P�"Oޔh�l���8t)e�	o��@J�"Ot���b��J�j<jJϓ+��9i"OP�@��/.t-�d�A�S$�,q%"O�LC0��9 �l��dB��@`4"O��"�S�o�V�����"O�%���ϕ|���{�����%�5"O�ԡvb]�ԝ�Ŋ�>|F�u"Od���+;�T���D	��P<�f"O�X%i��5.���c��.���XF"O>@K��+}6 ;ҡ�9^��Q�"O0�eĠy�hA���O1 �'"O�t��W<ܤ�3�*b�"OjD�W�U� ��`���"O��*B,9!�0�bGG�
��"OΜɁ ^�E��tF��)����`"O�|��悌k(���L5}�T�q�"O�|*�	�\�ا��j�J���"O�E��T��3����p���"O.���jZ�CkV+�H�u"OJ<Rq��*7lz ���K�pD�z�"O�ɗ��C�:@:Qk�1!��b"O�I�Q��_{R�����.� �q"O.l*E ��$'�UM9S@�zb"O���4���"$� s5��z4�"O��i!�)����d�� ��$"O��B�K�B���w����ٛ�"O荳4�&�8���{���"O� ���2�^����Hp�l�"O���mP-�����`5P��"O��;���=C�ؚF+	 d��"O�s7��B�هq�Z�a"OVm[��D��݊�Le6n@�"O�" -L|�dC�`C�&-�E*�"O �������؃T`�g"�#"O܍�䠂�.	ԩ &�9۴���"OvI`���s�D�b�d֬~�Ѝ
�"O�ʄ,D-B]���!G� Q��"O� �#
e�"m�#�� q�t}��"O6��VC$L�-X�B�j��U�"Ot�P��Fo.E�uK�'VvV��"O� �YI7�I��6\�'�G��"xbe"O*�z	ΆJ�bD�r&� z�uY�"Ov�󱃐/3���Qե#}\x�S�"O�|	�肟==����Ϸ ��)��"OV43�
	�u��P
�O[�uĈQ��"OHuJEc��S����I��@r�"O��A�������+}�:��"OZ��%�*->Ι�b
]3 N�)"O���qN�x` �!�� #�E"O2��&���N��!L�Mq�D��"O�����h��l{�,�*7���"O:���IÑ|f�J@��k}r Hu"Oڅ Ì��iH|+Qa[)^<�2"OL�8��L4R�Ρq3��' ��2"O.p�S͂.��q �1ߺ�q�"OdX�IF��%A��:vl�0�"ORmA�(Y'd�r��3{��t��"O~���$K�K�]i7��iW(�`�"O�p �.Ǔ�,��A��=�H�"O((�1D���(4�P��`%¶"O�g͂XQ���K�J��Z�"O�AȐ�]^�d<�c��|| ���"O�����9k6��c�;pgD��&"O��Qs◐15 $�v�D_ "OV	�s�Mcq4dB�	��QJz�"O�(�U���,����CG,^u��"O|���=X����. Ihdj�"O��!!��Yjl	@4K�?mΙ�"OV�(#g�
bUnPsŇ��!v9"#"O6H���3T�l;�HY�0"����"O�K M7yw�݂TX��"O8�6���U�f% 4�.�@5��"O�ň���dL�80�U�x�"O��@�g
-]���Ҋ|�:� �"Op���!ԏ?�2T[S
�e��a�"O2���#��-�X-2��%����"Ob�9��ݨV�Q�@��tQ*"O~`�ЃW-q����4Oƽ���@�"Od��7N]��y��M� em���E"OFd�	*o^��(�f
�\>���"O���E�0A%�8H��X'|Aȅ"OH�q�E�1{T�h���2B"^�#�"O�u:��8D�Vm"@IߺG��p�"OZ�����S�N�҆m���qRQ"O�H��kj$Y��k�}�x�"O����!�?H
���/x�J�RW"O��;d�?t�l�*@�?���"OH�(�&���e(ҫ�1D1:3"O�]��͆�*�,L��)ȿ
��C""O�����k�q�A�QQTPy��"O.�(��� ���i�M��vI�2�"ODH(7�	��-�DB�)�`��U"OH��԰+��c&Z'��l#�"O��vɁ�s�h�҇%��4"O�y#LS1 Z4�S�`y\9(S"O����O?��P��եKҎ�d"O�AJ��W)�a�4�֫<�F�	S"O��HE�E�<������A�Υ��"O�=��}0�K��5hX�J�"OU����D�X�	U���~0���*O���$��
����-<4u:
�'ɀ�� ��!�N؂�HW�NCT���'�����!�%�� ��o�@�(I@�'j"!�F-,x�	j��
��@h
��� J0���3Ǝ`�.R��B"Ov��5�ʷoL��� X� ��"O:�t�ˈ^_�$2��W
R�*	��"O.${��Ew�a!A׾p�x���"O�C3�?�Zz&.�5"�٠�"O0��QLώB�r�aq�21czT�v"Oz�#�E�,[>�"�a�B�J�"O$ܣ5�X�tR�y�@[���}ȶ"O�4[��Y�
�a��f�&�"�JQ"O�CbX���Q�'��&p�� �c"OT�"RaG{R5 �(��ޒ��!"O±≍�U^�����$Ʈ\á"O���"%s�� ���4WH�X�"O�YҴ���Sj�H��1+�h!"O�D��f��d�H�֦@,I(�5�t"OĠ"�*��Xf�84>=$��C"O��@e^�XI�PNgm4@�V"O�A&�x����6vD�`�"O�|��AO4�I#2,
�?e<��"O&�R�".�`!���[%J��
F"O.4{W�ٙ"o`�����;9,���"O�MH�')��8�#F�����"O$��-J/#Eb�u#�tk\��"O�����?>3`��#�	?@��c"O䚱f*p��\�� �+G���"O�̘p���:i�ҍ�F`���"OR�j���-0�~)I�댋0D|:�"O�`�d�N~��S�G�$?F\AA"O����'4���b�B'7��[�"O|����o8�@ �v4�[`�<���G� �脑�[3��%�p�]�<���ɖp%�yQ�K�C��	���V�<�Wm�X�h"�/U@����\O�<yQȒ�If�����)`���A��WO�<a@g��<�mA�;�Ե�@%@�<Q2_�:^i�B�`F45��B�<��뛻/�z�#�ǖn���̞Z�<��R��Xĩ���rFXt;�M|�<ْ)S�r�f��2F�m:~�h�t�<QX�jm:!�'@Y6����ӢJ�!��
6s�����@[�>`ٛ0���X!�ǜo:X5��`Q�T*6��2n��N!�� �v�5+�͏�$�����ՂH!�ۙnE*��5�
=R*p�S�R-#X!�Ҫ[	r����3��
IH!�T83�6�2'��U��Dk2jَO�!�d�#2� ��wAFE�ƹy�FДC�!�d<m6�k�
�?S�� �D抂&�!��w">�S��W�h��%D	�!�0c�(�ړ.ӕvjH���#�c�!�d^=:��r�m�!xFl�7Csc!�$���٘r�_+j�B���Yc!�H<<�T@	K�GV,h4��pF!�DL��p	Ɔ 5�t���OϚ&]!�d��y,T8�%b��{w`��1D!�y���1��r�$/��U?!��
8i����kX�DH���RЫg"!�$_�t��e��E�b�9h�JX�;!�D�1&���p �Jj&U��.`!�v�:|��7M�e(�B�>}!��*h�Ї��G:q��<Za!�Ę:>�T��a��Ɋ�{�	�WG!�U�n��W�B���E'��\A!���2������ԪQ�(���'!�� 2E���b�*�/�QYN	у"O`�:�N�%H철��:;|���"Or��2�Сq�D�탳=T��"ON��t�J�q�,yZ�ùaٖ@��"O�	��lO�\�RPlݩg��*e"Oҍ�L����KF��/fo���t"O���g���c(�@�2��+hZ�A�"O�	Z�bN=y+2�;¼&�����"O2I)�%�=;��8!���3�,u	B"O.-X�)ܮ~*���1 ۾ ����"O�yC���}���rga�'�zM@"OR��
�-{�l�B� ;^� ��"O���0�\�
�y��.a@2"O��`D�vr� �.R��uY'"O0��w�o��xÎə	غز�"ORY�g��0�4��L�B����2"O�uҗ�u��4�Z� �x!1�"O2�#�#օ@*�9��	��Z婇"O*�i
=*��a�Ǣ'@�"��"OzUh��Y���;��]A�Ҕ�"OP1
��N�{r:�8�I"^V�"�"O8|W�4�Q� ��� ���
Q"O�jGm�*�07���An.��XY�<q%oЉLwB@�e�Rif���K�I�<	�n��Dp��ĝx�)���B�<�f Wш����r���QhH~�<�$I_4]���B��{����p�<�ӆ��Q���k�]�cg�� &�GA�<Q��m�t�@Pm	EE�h FdAs�<q��QoZV��A�Ε5*�,�m�m�<9�D�&/�
QZr愫'N�5���Vj�<᧯��g�q���|�諶+�g�<��k�*!z*Y��iX2.��[�*�l�<�T�� ]V��B�+�*R"h��h�<�!F�;@f=A�C�k'F峴�Jc�<��*֟r�{�,ʟ(�	A��f�<1r��.��j�뇜%e�H`�`�<�Cʁ�j�,|���*��툖+�[�<1��dBV�ұ�z��(K���Y�<!��.r�afe��&��C�j�<�1)�'n����=����#L[�<�F��?���آΗ6�Vt�vN�|�<Au��\�t+RE�XL��Hy�<хI�^}��9�ߘc�<���u�<��F/�fX�����tC�H�<-�Q��A.��u�A,�f\p�ȓV����GB�}��q�fL ��<ȄȓJ�]Z���'3h��P��nt)�����h�h�,R�t�YPi�
spe�ȓp�!$l� |�Y2��8�O�Z�<6��H$iZ�Xq���V�<Yf�_�/��aHDFJ�.��|�<16��&C{�L@"/�<56��b��w�<i�(�O%,���N׹	��sU�N�<���q�� �&F�!j��ۂj�Q�<�XB@pk�� \�e��s�<)	ݧ(���Jގ/|+��F�<�%e@&?1��-P�N!��:D�D�<��MM?u�NɲRIYF���{�d�y�<�Q��p�@��,ي	�5���m�<�4D,YDPSq`��,�Zc��O�<I nG&'HV, @���tS�v�_p�<���M?����)l2�&�o�<�S�L�Y
�E�Cֈv���j�o�<� ꜫ�@Ć��ˀ [��4�"O!s��G���)�\��艀�"O��UdݧMp�؀A�<�V�a�"O��{��M�}��p�Q ]V�D��"O��AT���2^�������)B"Or�o�H4��K@����ȳ"O��"@$3Y�*�3QKγO�~(� "O(L�#�
�uUtX����0�֨k"O^-3�@�Nj���C����9�"O ��ؽv�&�%!G>	P�8w"O6��'�:4k��"O�o�d�F"O�����C�dF.����2~�%0""Ob�K��AR���^�I��x�#"Of˄+̉P��Qٴ�	vӆe`$"OT�˧L�K0�X(�N�1l�T
�"O���n\�tg�9{-T�,�&͘q"O��[����U�r"��\�����"O�����"%�N�ڡ������"O �B���0m��S$��7KXtaV"O����HS:T��7&��L�b"O�	y�Je< |�u�\
^��80A"O�ВG��>���8q�bűf"O�<�`C�5�����4s�Ɉ"O=��k�	5p��Ȑ��D[�8j�"OZ�"$��q�H��2�[�}A��u"OL�T�WVNp���-��@���)0"O�0 Y�2a څ
��zj��"O�tyI���+�J�d��Ę�"O�d�� �� �P	O���}�"O�e귨���I`A
T1�5S7"Ol"�
Ȇ<�Q�ċ�)oݖ\��"O���`׌j<��B����n���0d"O�e��	�X9��ᦊ�3.�,� "OJ�EG�|b�mq�ύ	���hR"OB��W�A9j��u��V�u�:}�"OH�AH��b�� ��MO�y���3"Od0��[�e&rS��E�^(^��S"O����^�#� � ܏s#� �"O���dC&[䐡S'��'t$��r"O 0k6@P�/D�=[�̈́Sd��[�"O�t�pl±d�N���dV�I*"O�0��Fld= Fҕ(M��C"O�
�αn�������B�$�"Op�c�m��1q��v<Z�r&"O�0��st� �(U���*r"Ov��"J���=Q�.�_x4E�"OJ)B��Y�Z0�J����nr��ж"O��8g�E�_6]Y�$�@k"i�"O�`�%
�����MT&O����"On|is�5]��)B&�=0����"O.T��	W��N��c嗴/,�Y�"O�-3"("�^i�F�јCwx�"O �Q��W9b��z0AF � ���"OP��ܒ1p�p��R��a� "O��I2E\"fz�pQv��u�ءc�"Oʄ�e�MԺ���= �P�E"O�|�4b�}R(�0dA�����"O
��d�!5�\Y���Q�`"O�����)O��{��ȶʕ@`"O�h�ևڨ9��2E$�%׋�y���^f`�B+�$����3*�9�y�坻F�p�t��QV���f��y2�ɷj�U������S�P��y��F�=�N���(���7.�	�y
� vͣ����NtYR��7Aڔ�c"O�hce!x��0�ƨW�;1؀��"O<e��d��u�Zi��F9~��l��"O UafM��iUX��G�"Y>}�7"Or	2U�>8�>�����)����"O�%!�*�)"e�VDH&m1\9ȶ"O8ԸX�g����#�Bǎ�i�"Oz�@���'nS�$Yҍ�4VY�Ej�"O�8:p ��7���p' �'Y�"F"O Ё,V�	�#�&
dL�ևP�<���U�<��a��`N`�8�]B�<�U�>R��̲]�����Bc�<I�@&�l��A�/Y�ĉ��@a�<�mC�:���e���Cc��y�W�c���f��*g�4�8�i��y�j�3>�-p����P�4s���yb�����aa&�M�Mh6I�7�yB$֛���*Į�F������+�y��K�lx���?S��Q�T�ك�y""�����; ��>B�z�e"!�yr�\r��s�L�"��	�"�yB��$<���E#�%Gb6�`.��y��A�g��@�DȶE�A�kD/�yb'�F#���@������^��yr�������5R��u�ƌ�8�yr*�6)>�	��e�1iڸ3�b��y�J��� 25�Z0@H��A$�yBd�7�vQ��"A�H]� �_��y� �/6�EC��ĺf�]�� ���yb��~8r=H�,Ff���B��y�-�o�e�w�X	����Ej���yҏ�g�P8�aD�qh�(�%��y"��17��y���4���B�;�y�o_��i �&�|��4��y��2*�Q('�þ��㒨�y��K�Xct�ʥ#��A��$$�yNF�zj�U�!Z����@V$�yb�ű^�v��@j����U�^��y�/c�Nl��O�|�켡�^>�y���A���j��%*�j�;d���y�b��q�:Y2E���u
#ơ�y�/Lxyx9  o��P�"�ٙ�y���@�$������0H���*�y��t�i$J�*��@�yrh��_����,8j$z��҄�yҩO�V�SV�>`~&I"�̘�y�e�o�L0#�f;��`e��1�y%S
+���(�:t�ָ�d 5�yR�L�3]�����WZ���s�۶�y��Ο
S Yh�3� }(���yb�B6�|�21���B�J�鈣�yb`�v*�y�.�X��rф��yrj�1���(�N�"���k!Aɇ�y�S9`����#� &Jp�g�̸�yR�*i�8�����x<fPH��^�y2�@52C��2Qねj�,�����y�!E�)a6��Vh��k$���y2��"|Ѳ`�m<���i�8�y�j��<���<c.��[�NJ#�yBn�[���-������=ĪEc	�'�CĆ�OS�!u��:�~]a	�'�l��Ao���i�3�R*^n`�b�'�ĝ $^+���+У]�A��@�'����$$)��	���?7�h���� �H��'�t�E*T�~g��96"O�}+��֥8�B%aϟ^U��
4"O��J3��2�- ���6G��Y�"O����v΄�a��r�N��"O���M��"� tZ��ʊ`ȂX�"O�Cq,��%��($]�eRd"Ot�U�פ^0u�eF���s"O,@#)=�&��_�1z���"O����(��)��A�8  @5SS"O�͒�"��:��m^��ta��"OĝР��I8,����_�x��Y�"O4M���Ć��F��3 ~�)P"O�zw��5�,�RA
��%�
�1&"Oڄ�M5#� I�!��/	���A"ON���أ6��Tm�/?'� ("O|lhV
�|�\B��ƤF�h��"OZ�sf�
Cy<i�v(?�(�"O�虄%�M�B���I��P� ��"O�u�VnS�~Eـ�L���#"Ol��ŏK�l���4�D�`��Z"O���H/Z���XR�C�G�!(�"O�H`�Q��3J�(6�r�"O�@"qc��]l�
�mjl�$"O�����>l����J�J�$A(R"OZ$RdN]2qv|��o��5�ҭ��"O��0<ch���I�eʲ0�1"O���fkF�D�^4����, y�"Oȝ#�n�2 �:�`M��m�8��"O�����C5#B����E
�9�49��"O~���E��u������T��"O0�@G��x��Ȁ
K#A�~�i�"O��
t�\Q��r�Χ}�,�(w"Oa�؁JG����'�=R����"O�q����*C7@�R2H����Ҥ"O����T6D���q��4]�^�s�"O��RUG������ЎS4��:�"OX�Z@���m�Ƥ�0�"O ��ΐ��E��M�#���K�"O�I�P'��i+�n)!�����"O��X��N�MҊ��6nĵ8:�՘�"O�� I�JL�d�6�:( r,�u"Od��*��o�Q� �W*R1C�'�-SW�5'�����+��u�
�'�Lc�� " �J)Q�gОF Lh
�'�*eq��a��"��8m(��	�'w�Ԑg��?^�q2���S����'q�� ���4�ޥY% Q!H0.��'�<qE�Q�P�>�Z$I�
�2 �
�'���#C�TD^��f�4|��Q
�'��e�7\��adC����!�'HHd��l�4 p�u4P�'��5Rv%�#�8��(��i��p9�'�4���V�7��;$.S-Px���ʓ+��a����/hMSC��/K�ԆȓQ��y6�ʑJ���z� ��x��i�ȓ!w�hs�'2'Ǣ��.�kf9��ɬ��V�CL,�H7@�Z��ȓt!���H��5����E������/��KD�8OTD��Y,3�ڸ��[W.h� �لL�(R��֩= @%��1��9�cX"4%CfkB.eޅ��~�)bM�16|��rr�-E����3i9
�J�i��R�䄴R�$��ȓL�kC�>r� �� �ѥ(�$ȅ�S�? z�z��ثM��;�n�!Sx���1"O"�i�*�s�^��K�c,�s"O��У��"VQ�l6Nڅnx�[e"O�k�T��	���8m�i�B"O�L����BF�R�(��~gR���"On��%J� �ځ2QG?iUh���"O)IE"ըN��}Z�臖W8BQ[�"Op�4�ހbBh�($M��$^��"OrU���4K�* �&�� J�"OP�b*�)=�#LM� @ aa�"O�8BRAY>]�$i M�$�w"O�@�uBG� $ �饢6?B�u3�"OY�2�P#�F�Y%�8&��s4"O�]z6�����w���$=��S"O�x�� "Up��5
�5��[�"O��{��Y�(���Nԑ~�,bB"O��qɝn�����M�.L�p"Op|b b�T������#O�"OBQ0s/��l�f$b�k�+|�~��Q"OX2��ҪB`N�Ȗ�S�l���sA"O0�@��,�<�
DHH>q���`"O>��+�+_����Q�/�rqR"O䙰�2W8��� 1W�H�2s"O��J�\��7����*�"O`�6��3�d4�p�Ɇ.�L�"O�t��G�*�4��DI��W�,y�U"O�M��K�����%��%Ԁ��V"O��	�`J�a�X�����+c�V��"O�11$��g�ɑ�n�?�t�
"OR����˔K��0v��o�NX�F"Ot��# ��Xk�0Y�]'����"O�e�W��	,��{�M�}��Q"Oމ�'`F+(��ˡ�ϲZ��	�"OΥ:��=|Fu�U/�2�z��4"O��qc�/��D��%$̊�Z7"O|!�a����Zw+P�~�dAs�"O�Ita[�n��x3W>[�h`V"O�YH0��=("�	��Ɋls"���"O�9a��!;
`Y��ߧ�D�""O� :�+ĉq��Qcɐ�i���p"O �P���p$9�.	W�x�"O̽���ڸb��s����CBU"O�2�AN�2�{6'6O&�E�"O` ���?9爠��%AS��!�"O�(�to�����P-\ԡ�"O`�A��I�>���dCQB4�A0"O�Y�@ͨf���tI�*(�Sb"O``yu�F�yE���ք:
�,9�"O�(9儛�|/���b�>R�x��"O�����2��m�#��.�"e9�"O��˄���zØ�*�Ɨ5.^�S�"O����ʾS��@rM�BJ�q7"O��2&d�9x��H�L��L
���"OJ}wʞ"6��0ʐ�7[���j�"O,�8���a�D��s��-Ռ9cq"O.h�g�ԛ(���ѳI��\�L�"O�qs��(�P0��v�b���"O.Y��]�n]�9��hҤ-��9�F"OP]:�#�4�)I�A��^�,C�ɱ=���Ɂ�%��0C`Џ �B�	�a�蹈�8j(�t�%��l��B�ɸ,.�z#�C7HPH����W����'9�E�AkˡcYR%s��V�^;�!�
�'htX��-G՜%��/�[і�	��� θY���%�*���]�H�:TR"O�؃�&�i�\l{�b �&D�u"O��Vހ�8p��ʊ((��"O�uB�.��/v.�f�
��6"OR͑c�;d-z���mX�I���hW"O^t��,U
sa�m�0�3�t�zG"O���ǆ�l�9�W�6��5�e"O��s�̉� k���Ԇ1^���+�"O�l��N���zY��<y�J%�y"�8I
�!��퀑�,UC!b���yb�.SO���§v����P���yB�G yuhu.�aP��SGV�yRO��CO�9W�7
]�A(�8�y��˨?m�B�S����)����y�bX��MbOX`�4�(þ�y�i��[D�X�5'.	�����y��!@��bT��H���!
(�y��K'$��&&�t��4#����yB�ϵ"����UjS�|O�ЃB�Ҩ�y��O�v��q�e�|~f0@g��(�y�*>^������>o��:�_��yr��!H�����rA��B���y2��"T��rU��Y�u $�H��y��+���R �U�Ty�靋�y�����S��^�E�n��l���yZ���CW�&,�:P($/̇V_d���Pk�|{Dc�0/��*��̄ȓ0��b#KA H�����o?B���PY6Ÿ���5Hfر@��'Z�X��F^<�ukč8�2�� [ٚهȓW��u��@�����zV�Ѳښ��ȓp]ؽ��"֭j�\����ګk	����17�[��ҌR�$�Tm�8B���L���ˑ��=Jv�r,�48�A��N�P9���&bm��1'	1~Z�ȓ+	��H ��cx�)ҭv�̆����rR�Y�J�9�$�Q�'�����<�u�#!��~�HE�RHK���J������7��@�%Iز|�&���r�d� OK)qQZ�N�yI��C�q� ��#��!������]�ȓ'�L�1S
Z1�����n=8��ȓg�2�9�ۏa���Qc�U�(�6u��m�P�BID�f®8#��V�<	FC�	�S�B���1#ؤ���
GPfB�I�H�x�f�/������@B�ɭ!BL��7��)B�&B�I/0d��C���H�Zq��/	FB䉯94Q8���=�Ѐ��ʧ�>B䉹h��5�J� �Ԩ�S1y�B�ɿ1
�-�E��E�v8�2!\>h��B�I�A���X2eR�sn��&ZB�I��X8�7b��@8�gIWf�B�	,�-���_"V>@ܙ7�¯g�C�I�m�|�a�CXT��5e�J-&C�	8���[�)��W9 ���ݩo��B�	/+lb]��@# ��x�A��C�I-:;�DkR��5w�����Si:B�9 ~���%E}�T�%���T�"B�I49��9 "L�	op@{���C�I�=i8�%�O�R̪s�� ��C�I�yn��M�80h�&E
�BT$C�	^�t�Ѓƀ1e��	 ŁH�B䉊H��!�����B�� m�o�dB�)� `y�g��(+�x���S���5"O�a�E��<�RyI���
x�i�0"O�PA��<6Ԍ-CSJ�0�l�Y�"O �BrgR�`\ˤ��NA9u"O�y����V:Z�K$fN5B�X�"OH8!ݖ3��H4D��Y/�Q�"O�1���҈Vt�%B�-&Lp{"O���ȜzUf�A&��^�Q�"Od$��
Y�7�.ey�!��t����"Or��֏ V��lce��#/:�"O<y��V�osN
@O�75�%"O�����n�p�p�M�>��"O���յp%�d;�,
 �TK�"O��{e��H�8U�W�(8&�R�"OF���,����$h��!V"Oȴ��C*?8pTi�>A�FՐ7"OT��#
6W�P�҈\)��1�"O�4`��ܚ �%k0ə9@�s6"O$�����H���`#	��Z� �A"O>�8�ڀsp=#`h� Pd��q"O� 3_Xu�#�8|Ϙ�v�\+!�լP{ ���������!�$n���s$H��i��8�ӄy�!�؊
��h��e�,���� �!�$������f�@�@�(�K��E�!�D���#����R,0p�d�%f!�Δmqf�%@7X�%F�&�!�ĉ5���0��Ża�zL�d� !�D¯z�j�P���K }�6�^�U!�D� �H�c�Z6�U�0
Й !��~���������!@j@�n�!�0�� "��e�$}�wB�/|�!�D��xT@qkDhZ0 ��	�!�ϨI�>y@��]�1�y��)M�!�DтCgf��#+\
~�00�	@0hN!���T�t�?Ю�9�MV!�D�E�H�����Y�rժ�J��t%!�V8D�q��(]��<	Gҟr!�d	M�ܐ��CQ)X�:�H擠!��Zx��#�K	D�I�D�0�!�9 SVt��b���4���͡}�a}R�;?	�&�nw\������HÖe@N|�<ɵf�*ɞ�	E_:0�Ě |�<Iש��A@�%��NA5'�м`,�Ah<1R�?w/�48�@��`�PyCEoϩ�y�"0u����E�S%�a��պ�0?�.Oty+ŭQ�2pX)֠2���������;z^��{�k�8L��B',�JUT���<����z�D��ҁu@��Y� �c�<qO)7�Ft��ǀ�a�qVh�i�<1U�&eXh�ުg9LQلHN�<Y��^��:�h[����P�l�o�'5p�𩗸P	��z��'3�΁��ڸ�!�۩VD,�VO�D��x2�"��	w~��;�S���RM�si��ey�Ѣ������>��O�H�F5X)4ɻV�1,�T�eЖQ�"~�	��X�#�H��z��@O#LEdB�	l��װ^g��2Gƛ�F�,B�I��P�jsF[�?v��zPؙd��C�I2]3�Y�G��3ň�vNԹ�\B�	*Rm���b�ɂV�`,`�Q�0nC�I�8�
1��n�).|q�j�7*:f���1}�bZ�$��E`
*�e(t�*���p>aԍ�: � �D,�=^��G�h?����4�i}
� ~X���)�:�Ѡ�ӫmbm�"O5��
�!Z��D�Rc��~0V��㝟��b�<�M<�~�Q�
H��ò#��$m�q��c�L�<�C�L&�l����B$�����Ŧ�q�x���<�}������K�_�jI��ʚ�Ysdˍ�y���%da}KS�I��E�Rj��h�х�h�P4r3Ȅ�"���%�W6���G}�5OH��5��
��Z�iƧT_�4��h�YC�C�	�s��3	�]Ԩ$P��R$?l�$��	�<5�ϯ�2#cK];BE"�it(<����a�
,�bgE�y�@�E�u�P�>)��	U$� ��J^�����݇�!��Ƅf`&��"��(�H�ze,�+?,!��z l]:S.��
�*��V�\:�O>��d	'�fd�1!�3]�x�	UD��n!򤙄8B��aہ8�$7M;{ay��ɟ 7��׈�+</$I�����~F,C�ɾz��9��X�0T@i��, :@����{�f#���[�R!�� ���$Xb%Pƅ]t��`�'qzqb@"��G��K1%D�;�' �`��	�,p5�g֩a*�@�H�K����>�ǚx���ⷥ	N��÷�G�@��d��I)�j�RQh�11�	��d��"���>����]�P��pP ��(
�$q��L-3 !�D�Kj� �rB��<tppa7���!��nP&�#�O A��@Sf�	' !�dX�$�0Py� 5�a��͋3�!� B!��C��4F%Jd�A�C�g��{����O��� �&bl���@3�Љ�IDq�!��8C�dc�o��){J��7��'@!���(�q��B`z���+�@�!�$���W'�3}�#� 2ԾI�<����'�DC;�2�B�KND- 6/f�x�'E�u�ԧ_�h��t��0�`h87�.�y��Գ��5��;)�成$�.�yR�O��m~��I��.�����c�%r9�$qQK�OO!�dD3y�P�+s�E�5O�hæ�\+@L�	r?٥�4��M,O�!*ŉ�dv<������@�ؤZ�3O ��$W�f%LEp���T@NX���`%!��.%x����ե83�y1L� �!���i�P2e�{p%r$�Pg�!�d���{���(��m�C(������)�禗�|>z)pK�Do�8���!�^0rQii�灀M�J��1F��Tq�$����d�O��(O 1�e�ݑ2�İzAk�?�0H$
O�7�ߣf>��5Ŷ�~�ӱ���G\!�dF�hƀ����"���ZH[T �\���(��%�I6y�T�)J�Wr�| �[�؆��?[��aD�к� ���M"!�JC�	p��%�0 	9o�M{��]v%C䉯O����B��a����3	WQ��C� 6���s�Ҹ6�8�`CA�\}rC䉾f#�%§G�|rĺW�]�.���c|a}"�F<Z*�H�Z��Å%U2�y�,Ow�Y��L.|>f��#jĮ&��b�����2b��'e���� �;Q� �E�'�D��y�$��M��DNV2k�ʠz������>a�r����s�L�+(<��&�~ �\���MpJ֐a�N��-�<AT�h�<�$-jɸp����X�<YD��=����W�W�o����(�o�<q�g�b�ji��!�4�GY`��4N�<E�ܴC�z���W!hF}�!hX���;�h8�v�+�rԹ2H�"W���'Xņ�)� � A1! �m��<����[v�0���'T�0b4@��D�V�G���R��j t�
�'0���˭g���@�½/x�J>��y��I�|G��R/L����Zj��'V1O��	�E�@��v�Q6n0�i��A�B�	�a��9�2+�T'��ڤ�ϖC-�B�I�%��E`3f�xϜ��eFO66�xB䉠vh���e��G���IҦ��g�2C䉝TH��O�Zgt��.ݰ4+�B�	�a�H��`[�-� h���������9�(O �J�) U��|*�,_�킳��J�'��NV�&��X� س��ҭo3!��(���r���N�<(֭�tF�I[��H��ע��E����� рlg�Y�f"Oe0�Û^XȘ��@�5kI꼢6"O��ඃ݉u�:��Љ�8G���{6"O�;�T�tW�0x@fOz���Q"Oh-���Z��
�	Pf� @8��"O��+5�Y�jEa��E�	#� �'"Ov��w/�M$v3IԟL	�\"O��1g�ןIy�x�N&0���:4"O�$�-��j�\�8�Z�k�bM��"O�����ynx���,s\l�U"Ob@�`ܪBp��ZQXbe�w"O���g��K��lئ)I�m2�\*E"O��t	K"Zk E�T��1"�1�"O�����@����#]�R�5��"O���1�@�x�(@��ۏ_��;"O��(2��2����bT�>Ce"Oh� F�C�eᚵ�T #Zq:b"OԨ[�D �F-6����՗*f��e"O�hٖ��*UK԰�����p!�"O�(�JH�\���Rn@?!�r���"O�3�ú2��:PǓHؾX��"O�@��[B`���D=|�$�ۡ"OFL��Y���ٓ�bB1o�`�i�"O�᥋��J�ZMАa�9[|ʁ�%"ORe��O�	*���B� �Fq�ء�"Otb�%Rv*eS0`,\�� �7"O� �d���a��O��,�<�"O� �ႏ�� cDLD![��5�"O���C�gލ�b��>�h��u"O,�&H�&v��a��Dq���"O(|�$jտ[İ,x���M�Ru�"O����JʓT�L8:@�>o����"Ot�+��7v�d= q`yl%£"O���bK�'MR
��ь ] 5(�"OH�ѨY�rrLQ�`H�)���"O�M��.34�r��R�]a"Oꭙ��Ċ|�ް@e�>�z���"O|J��3hW�,� �~�@���"O �3!�� &�%B�̀�)�D R�"OB�0с�#4b5¡������s"OX�F�1xG*!bQ��1��
�"O��+f�f��0ƊD4���w"OX%��(�Zu����D�""OhY� W�2��H���ɒv���"O�A��`O!֍�DLR�p�B�Ra"O�iq��2EI���1	u��"O(p�rኛY}��ؕ��(�z�,�!�$�*s���BR'�.)�$�nO�z�!��YD��`�l�l/��!��V�g%!��$E/�A�c ]#���#7�4
!�$O6n�t��J/~���L�T�!�� x�X�̱IZ�PC!�<*C���T"O��WlJ"R��KA�`MV���"O"t�Bn��\d�	Q�X!ZC��q�"O���L�{���2ď�3�1��"O�pb���E0����/����"Oʌ21MU�;�0���Bҽ'[,��"O|�b@�Ơ� ��G�-��bQ"O�yu`Ё1�|(a��D��"O�jC�^�Erށ@���:̾p��"O<<�3C@�kZ6A�ࣃ?%(14"O��
1�`}�i��9l��0�"O��A��/<D!&��^���6"O��Aơ�?:B�I�Rov�`�"O���i�$9��к�'�>�B 1T"O�y�`3T�R�p�ā�;S�x�"O��1�,L\[�| 	�oP�8�"OT�0߼A��3E#����0D�PC�	4rD�R D2)r�X!@0D�� d�Z��,Ȼ�B�N�b�CCm,D����6Z)v�{�'A�^^0\j��/D�����O�01dJBc*�V(8D�`�A�7V*�(��V��� 5D��8b�ԕ
<Q2�a�!��	�S�2D�D�ϰ,0��!f" ς�'�5D�4Cb�;zh�C�'VT���$4D����k�:PqjP-Y��$�ه!4D��2'h\2�69C��W(q��A��0D��
�	H8`}�C/S�7���e0D��Rs.+!���զξfz&�p%(-D��:�2!�����L�s��e�!� D���PfY�3$i�!F^W�p��S�=D�st��%vh�%�W%5�v�s+=D��i5K��m.�C���a�p��T�%D���	g�vl��/B�F�^��l%D���b%/w[<!��i�/�DM��#D�p�@gV֊@"=�&񚆫#D��X0'Bk^��i5BA�Cҭ)��-D��A NG�m��p���T9b�M3��*D��To�9S�|��͒2@���a(D��z��L��>l2S��&t�!e$D�Ԣ�j�֌z2M
;]>mx (D���&Ň :C�ex3�(G�<�X��'D�|Pө"@�Q�QOF����N0D�H 񡔥O����m(F�-����O �=E�T�ֱ?�`ؠ��7M�����8G^!򤖉$�i�!LčDLx7�7S!����vQҴ	'���!���5e���#���<%>)�'���-�Bܚ��g��y�"-y�'�\�v��o8���n�����'�17I�3C����eT�^v�-�
�'�0$z����k���BfĊ^� 	��'M�@�%����h�9@��u��']^��kO��N٨��T$e�� ��'��rd|���(���c�dTp	�'�:�F�Nܣ��	������IO?�Ó-��(�h�N�(\���i����
�'0D`˔�2�bQQ���&P!
�'^�:F�N}��t�nτH��1�
����0��O&1��4�U�yÐ�E~���(`�kP��8i˄�_��B�ɚ
��-1`�٘'
 UȔ�ybC�I�����B�2+8�R�&B�z G{��9O�����	<ؐ�J9Ӳ͓�"OP�3	�/j�f��牨XƂ%i��'ґ�� p�1G�rܰZ�E\�Y�j�@r"O��h�+C/��k��ŸS���"O8�r��C���ìlP�pKe�>1�K��P�$`S7� hBH J�<��I��?�G�^n�8� ��<'>L ���m�<�t�E&;Zn�Y�+�	F �ࣶON�'hQ?m�'��X���)A���u�(�Hn���� ���w=����l�L�+�v�A�'�O�Y��'{�R��d�P�U���*@(IE��%�"���I�a�,X����s���K�B�2�!�"���O_�hwJ�1�"@7�������GR?�}&� s��`��t�tLL%T�tX�QE D�P�Õ�v�{�	!!8J�
���H�\����q�S�9U�����c&4��a���Q�����3�$�HD��B�͒�xI �97!�/Q|x�#�ժ��(zo""/!�dt.�0���^�Rx&����e+!���7K����̋D�J��-Y�P��~2)T�<� jL5��)��27�d��F�<Y�E	w��{�@Q�4�4=��j
@�'*"~2V�B�5�B9є	�J;���$�e��|$�0�N���z��4-Ф��O��p��$,��d��*gf�'{2,��iUl4Y��kL^�<����a0�4�-Y�Q`�^�<9�L�j�r��B,G�Y�E�Y�'�ў�{1f�8s$�:<�135IU�!p��7��s.Mk��誵���8��͓��'�)�N�ؠ��`��5�d2�ۚ+ϔ��ȓ�V=��o˛v��=���R� ���ȓ	Ş��F�\ J+��c����D�Ȇȓ ؀�Rǘ	z��9�j�zT���ȓJ�(�����	x�\�VC�O<.��=!�����&V,�^�!��-G�P;U#R$�y"e��r6��;8���b�M���	hX�L�wd���*��`�J0K�����4D�H���v~��"'�H6p
�c�(D��ł),J���I�C�((�*:LO����C�+����P�`��7Ř�3ˑ�"~��$%N\b�$���چ���H�����7�Ix�'p�ZW��,�� �����࠮O�`�	�b��]#!BڋW��1�gI�HQ���hO�'�?Oڍ8׫�t�j�i��
W��%�'�O���m1d�<��tMJ�U��9�%�T���q��<E����8�HG V.�,�!C�A��y�& ���	��#���Bf�7�yRd_F;��h�(���(���V:���7��1�	*�ɾg5*�(���%��){��WO�C䉁a�������5$HQ�����v�C�ɕ&�}� ��$�P��5zpC�	�np�U`�u�T;#酘N��,1�"O� ��&E�=G��	���"O�)qD/�9+����sk��P�@M"�"O������(!���z�ߝ,�0��"Ox��֎!�E�-�H3"O�q*�$ݰ_��\�Q}\P"�,D�(zRoӟL������2�aZ�*��l� ?$�0�6g�8���oK&1�j��`��~��''��,K�I�5��\�T��3ar:��@"O����$� 	�D�l�܁�"O�(�%I��U&� ���_T�4�'�|����Ob�$����R��x��E�8��a��.�O���0>���"L�PpuG� ]��Y+V�D?A����
�X�΁�? 4����ZLEB�IiD�b�_�e#���G.j�,\�'8 ���OHY ϟ�S�� �])f`K|BR|�#	 ]�Ppb�"O"@S�E���Xf�,�՘S"O6��gL�"9���СfN�ww\U1'�O��=E����n�8D󀥚�[Z<I9S�G0�(O2��DW�}�R�C1'̱K�<��%ǆd�!�dT1U0,��ãT2�:� $яZ��~rQ�����¤	А�)`�S���PN4}r�L^��wb�(�!%G+���K�nЉY�L\��1D����� Mb�A�IK350{Ԍ<D��C0m�:M6�͏i[ \
W�8D�D���=zx@�S$���s������6D�h�H�M\Z�J�m˝-ܨy�S�5D�\�fН ��=D`E&&���/$���.F� W���� ��p,�âΐ�y���~�~� W�;�*M�U���yRCfh�d�b"��*��rE���y;; �XRA��v<�-XE�J����'�S�OJ@�J��&I���je˜"cٚ@�y��'�,��@��]{� Z�ҥ�
�	��6�[�QQ���d|*Ҕ	���6	�!���#����Ǉl"�yZ0޺!@!�d^y(�go[b�*F	"!�$Cl2�	;兒b���r�J�b�!򤊬a^�`��^������L.�!�ٓr����Q�2�Y��7AI`C��?� �1����x�)�혿~J.C�I:<|�(�'Ν7�� b�'�l�C䉼F�,`"��ܩW��4B�%&_C䉕z�(��#�|�d�Ɔ +��B�	?Z��0�S��4>��q&�#<rC�ɑDߴ-)��Q����"S��`�C�	�,+���I��	RN����k�B䉹�|�	�?݊0qBb��1�B��3>����'�ݝ%��	��]�B䉫{��`R(نV������P9�NB�	$_���W�$n|pe��B�B�	)`��U�@�iJZP���ˤS�8C�ɶ2ciٖ��P� �S�\'6��B䉫����\�f� |�Q��5=i�B䉲c̡��Ћv4D��AZ5�C�I<1��U �[�bB�0DF2>�TC�ɍ8�x:ǮC�o��[�m"O2���/�:�b��M�L��� "O��2P�4Z"��H�,�o�����"O���F�= j= � A������"O"9$�V�c�y�A鍅R|�M�"Or��6�Y4SJ�r��{r�5�3"O��#����i�0�]}�m�"O:8Y�'�$M����(9y<xpQ"Ob�Q0Y�L��1�1�	B�}�"O2�c�Y�l�Xz��B-A/�h;R*O9b�c]�f�<j�"	�<g���'�\h����-�<�.�.� ��'�$�z�е.�������'�P�#�c��4��ԃ�>9�q�'u����#< ��@*BϚ =0�E��'�0��0�I"��!QK�7Y�|!	�'(^Pj�L�/I��疙1֚e�	�'V��ZE��F� �X��^�^����'/�t{�J�1Hc�-����#J��'�Ha{3��>�0��*GB����'V�l�]#���I�ą=
�lZ�'J �k�,KL���#�.,��#
�'��	5H<U�&�醤KPe y:��� ��2�MÆ�\�y�JO�F�vy��"O�xjP�۬n���F�T�gۚ���"Oh�9@�Cu��h�I�m��"O�
� ~�)9�F�'t�v �"O�����T�E��qQ�jՑi�ZH.�~"��vS��"���$�6$��/�$�hO��Iݐ$ڐI��H��:f0�y�"O�H��={�TL	���Hf��"�"O�p���=�J���a.l��Z�"Of���%�2L����@T�TNJ���"Oz���45�H���	͟<��"O��v��f���#�Ο8L�z#"O��� ��8͸Ų��]�U�FA"�"O���s��6��CUΒ�S�"O�y3�f�H�0���L�&Ԙ�@"O-�C�2��aC��B2uP>��@"O6���CH�E���?\K
�!e"O |z#Y�%6>�Y7(A-P�"O�9(���h��-;$�R\e"MI�"O�U�`�(P|�;R%VT`r���"Oέ�@e���!ƙ�Q���	"OP���yĤ��Te�V�ȁC�"O�q���`�\eB�""����"OP�!�������{����*OؠPf��%��e�t�5L�ݐ�'�>F,�<ona��B�$O��s�'h�2�	E^�Z	���ZC+L	�'((	�+[�&�\-�܂��Ib�'����d���k��;uI�~`��C	�'ʤ��`
�& ��cf+C&YQ�5a�'����B�E�ԁ`Ĉ�8�ܜZ�'e8��1���&��'�J�9GR̐�'%��:�'�L�0�:0�N�1����'c�t�×�Gj�RN��c��,#�'����h�'!���"fcM�S�z1
�'��2�#{f|}�u�ΝDܜx��'�<��wfR4��reE��O��'�5���[v��戧-���� �9l��@��O>ax1��M�g�ER��2w u��)� gB3@(B��DP�u�1�P�O�ZQPv��9<D0�"���]�t�Յd��j��'{����ϭt�B1r�"ɚv�~h��d��>���#�h
%o�1��-�4Ƕ�b�Ş�T��xcd�)0�����!D�z6`�'z��ـ��K�Q�I	��>���$Y<�Z��Jf�!#P@<p�n�?��㌨�lR�ǰYG�l��=D��Y��,[��5�bE����P��f+���e+��M-V�
`ɝͨ�R�M>Y�eӯcX�܉��X[��:AJ�,4_0�*�%�O��`��J+���R�%3�i��z�%-BNyB��D-#>D��DW80ֽ��������0�H����ą)*,l衤׹3ұ���%�Ȭy 
O
P<��s�5]]��a���|��yr�L��T���B�<^y���´�5˪=o��XeR)]�����\r�	�H�|�#p��
Qv���ʏ�`2Q�ꗽav��O�νi� ݊b��l1�Û'!Y��X�'�P 36&J��&%��LZ�� �0ai���ݙ���$���r�͵/�<EX��_+��`�a�,��L�R�S�d8�ՑJ?���Eܦ�x�L5c���q� �2�^Pքa�aD�qWfuPQg�(���y��9�$B��S�	�H )Y[v���[#�*��������k��r��.k��=�ѡ�K��0H<i�c�q�`�����3�iQ�1΀ ǭ�P���  ��6�1CS�͉r�>�I Xyҩ��Ș�f^�ӆIF�Xrb$�'$Ye�xgG͈?���i�/�(x�i��ƀ
urЈ�O�������Aa�W�;��IR�N�O!�gn={�)��M��8��������a?�(0��ǫ���kwf	9��H �Í�%�h��'W\3�I�%#�\��B�<O�Γs�M�Ʉ(���Á��+RH,s���$"���Nm�2
�6?}�A ��G"D8�gI*��M�cg\�fRjLpdS8r�@y�*�~���&��Wn�Q���O&�)��鉎M L;��V�\���=����t`��7��ʧr�dR�S�����ur���h�cD+���r&~i�1&�Q��h��B��x�@MA�/�k��5�O��kDʊ�}��ģ�Qr����T	A���3Ɓ�B;1��{B�8�J[����H��H��ʅ�S��JC�"��x(�5w�8\ �"E�b��e�Qg1
d��q+T\��#�  �� �:S0�s�b��o�� �B�8��a
	k��XP���|]�$��>Q�ǃW�8HG��$u��Ӏ�D�0�dPoC�s��y
��Oz�3�E�>;���#�
kpr�"�W=a�R��Ù�?�ֵ�&gת#|�+6��(?9���S
jrt���d���֯ʳf�2��ekK)l�P��k��;�h\����v� �a���������E4e�-0��/� T!�"EմN���e�Y�W���d!U2+SPE�48]i��3ukY�I\5�r�յM���զX?R��1�4ղ)T45Ԅ�m�<ݑ0��L�j�:!A2BO�@�6
S�
[�8�t���:CT�ȕn�4�	I�t�
A�BN���r炾 ��ě��:�D�q*ɘ+v"�;`��XYn]���(����"�����̋��V;�H�n�3S�D� cҞbr|�`�j�=�P��aU&;<�A����u���ΓeZy�CҞctp���M�<�V��T$3,�+ֲ(���L�Xh(I�N��d�S���c�Ɋ)8��)+q��k�	1���F�5�z)�@ް��QQ�BgEpXsr'ƧF��P%
��t+z@!�ƶ!|v\R��
T��Mw�bL`D[2g�&D�� �J�p'��iF�Z;�p��� <k���C�N5g�͑�#T��,�3��9���a۴8�|(���q��IS&Ϟ[u��)��T��@�R���yQC�z�E�*�m�D�ԡ�)e<aۣ��6$���� L�O��bS6?���n�>K扸4h�8��!�"g�t�I���މJ��'�1ET�ԩN�<~��ai��,�"n�����*M�9?N6�S3�O}��c�҇d(�����ÿ6v���G��;�(Q�;k���@96�7��j�(������Ӧ$J,Fܺ�Ȉ�h�i�F��oN�٨�O0H��a�ε$�dXr���FN t[��5:�zx��9Y@�:�m�X�
���J���D"��`����7?�tl�G+��]H�1zm'
�	"eLdhŁS�"�<!f�+N��7�	�2h� �C%��yj�	жL޴� *b!�ă&��Q2u�Ѵ
Iдh�JʳL��Q�槃]W�s�A0c���4Ϙjv4d�% �04#6�>��k��7b��bϒ�G�I�e�r-K�.C� ƌ� y�\�NZ�.ԛ��ȶψs�c�(��M���ە;V�l;0l�2N�e�G�ˣpf��D$�l�5�`Vܓ�y�ʖ��N�i��H8]��Q��aK��P���ܪ^F���e���L��ذ�I��څ���	:Y��Q��a

��t��\+\B��[�������f��_�9�h�e�'�r�X�w?y�@�!���:㑎QV.��Gh�")l6L�6�U/?��0UeCy�J)��6l�B��s鐌U^ ��'�� -d&l'��b��%����˳
̸��%�0ғQ�x�Jrg�^@T�g嘄d�t�*%�"z,���OCh�kF�ƀ���g��mw��h4&�2`�~,�Q�yX��h�cȓ%ޤe�Hڦon�Ja�O�0q�M���AJ@�W����@�È&ֶMX h[�ev�2����2;��A�k
/$V�!�$B�����,���xrD��i4Y��*4�V����oM4��&S%	��6�*q9*�)�Mɧw,�H�D!�W`ځR�C���N�t���y� )$�m��Vd#�}���g+�I� �N����7�D
G���z R�
T�\��A[q
� sd���qK�!�P���޶�@w&?�5.V��$`�3φ�it$��O�����µ	mL�
��/a!�%�H��(*,X��f�Xr�H�o�$7Tl�H��Pn��ՀW	g��d"���w\}��y<ܰ�^�4�H*t�S�V�1��C��� �ȕ"F�.�)��x���{.�2UhФMtHq0�d�4���Ȓ4�}s#`0<g�<J��+�O�4Z��K����i��̄.*ж/�0R����j�U�D���*�&�K�%���I�a�.,�0�r�����T1�4Ds��ҼHR��1�V�0��$ړ��5�d�ҕ'~�I�!!��a�\O_���sd�	]% m���a!q��?E�Y����2 ������V���3�Y�	^�O%�s�甸+UD�	��ҿ������'.�f�J(3PA/伄��D+t]��"c�Ԧy�*Y�!N�i��-\���=P�i��(T����`�-3���3�&i�R5�L�|��޽Q�e�֐x�'[�<�>���J�vt��E,|~��o^���pP����{>�����s~��X��}|���s�N�~�ٰ�?c\Nș�&ǉ3q��(�����%ĝ{iv��>Qg.`�d%�RG�Ru����D�ؐ<^�- �$�P�Z,��<��1���SJ�!"�o��
��D�Oؑ>Z�P�dسoN@� �B�7��"�晒;l<-����ΛMͨQ%�	0\�(��јbF���4��V��x�RI��S�͓���B�f��j-�X�J�Q>m��� ��	;��x�riT-S�͛��]�C�l��C��,ۚ�a�^0n�B	�֢/`V�*��Y�To�-���ճi'H�*���7т�%F�2h�Z!��4Z)ʼZEF{ݡ:E�O�a
!�#MM�/�,���G�U���x�a<�� ��!Ȁ�r�%h�b 1�SM�*��'V0x��C��T�ڕ'\�H8��q����-3(	��]xĭ���P:t��c��u7�sg6�`GA
��h'���ذ�'�Y$r-��HʉrU�R�!L�x�q���^�����3h	�C[T��b�-C� ҆-�&Z²�@GL�^Y��b�� j�bHꕌ��u�d�5e��-E�,��-��_Ƽ� G�^[���1���pꄗ)�P��cT�"cH�Nܓ0�^�q���0W*�t�&w�t@H�T�D�l`YUmT4��!+1��Z�`d0���W�Hm�`���������s��ayU-T���	�d8 ��
)l�`�V˄9%�bp[с�*'
(�rM�n�B���G4������-�D��kź�y!K(/<�R-@l���+R� ���Ȣ��s4�2�f̽!���`
X-	��HwA�(`g��C�L���� Ju �
�'A���'/�u�8tp�0����-{���#�÷�? ��{G����;s�0d#��>񩧴��
��[dG�{� 4�$%�<�,��!��>A|0��W� �MWh����2}��؀���*���=��Q��kK�q��T��M:9x��so^&��HI�hEy�N�y��I\� >d{����k��af"�8RoL6HT�0�%]�#�l. ,�̖��	�C��D��$�)j��B�l
�z@�`�ͦ�\�y�bN�U4`�11���{��9[��w!��Y�����x�Gʭ?�~��;cOT�sY��ZF/*<���1Q�B�~E�8!�4]��5j���? �@Р���$C���5̟�Ruj�������Yd=_� ��$�.C# �{%ߕ}<H���<H�2�2���>Pm�i�!gw٫��C,G$*�SE�{6 P����qQ�b�)3���P�8���!��&.z�
Q�<:θ���F�T���7����cL�����;.Y�����Z�t:Q0g�-����� ��HG!S�q ���R��-C6�PZv0O�d����5��x��
:Z%��'e��b:�%;���CҲ��U��/yQ��@v�1T��`��:Z$���j8����\?��ց�<^�DӖ�K`Ux�a��j��%��4���"��gh�y�A,��-;��C�Ýq�*�Ag �=�U!#���E���rWlÂs ��4+cl��v(�9^���������Q�h���A��Z�M	5n<������@�Iz}�Bʸ[�r�3�Ƽ"��E⭚�-!���%�F�R�b�R)�%H� ������Q%���	C�`y�T�:\r%�[���QD	�I�����T/��G��G�t7M��^�4��GC�vK,y�b�C2���O(v&�1w��(�*tis`��]�<��gC�wI*m���6��� ��X�aT �������w���
�	rV�Y��	l �� ��^.5䊠GUZ�	.�~b��Gr�Q��Nޠ���h����'ۦY���hq�L){p�d�Ǝ�<Cz�Y�%Ҡ����U�iߡ?h����|�t��tB]�d��9
�#� H�1O���z�7������/�(��g����*K�7��e��W*��YFN�	�M��9K��]��ᓴN]P��%�	�����Y�]�lT��rܓn5�E9g!��2``g&�=z������r���Q��:j�e{ ��|������%3��Æ�4A ���
��I�^m)�iSt  	y����4��!9���޴VSi�aQ:9xH%) ꖸZ�R�Q���w��#�U�|���oS_AZG��8yH!1P*�:^�B�1�e��C3<E�0jM�_L�-�F�V;/"��@4#�����E$�j\|����_�@;.m���I$aLQ�dɛ�B�9D뗐k^XB���J��UԠڱE�h)Ѧ�E�hRe�DI��G�9D��lNh�S�}��8 �0g	���4�C�5I�A�G+Q��c�����?->i� �tY��
D�����"�'��-�-+g�W�Ep�� P���b-�2tMj�a�$��8�tcI�K^1x2/�3�÷�X��qO��{0L�SA>tR`�@�|�D�/�< ��� �$��X�f@�9N�ʄIP�N)H6t�R�OI�l���k�������V���t 9L�Ƙq (J5|�b�i��lHA��$U�d\�Վ�:�*��fO|�m�'Y�L��i;h�\���&V�bX��:�"��pF��w�@���@�V��*MG�?�Qbf�Ζ~�AE�_!S�xD���c��L٧ \�'�J�)��Is���s%�0F��.\D�qR��t����&\�@�ؚ#�T"l�H��Sj�9$,@���Ԏ�;žr�͔;�VP�C���+�̐���!u�N�>�C$8A���n�:�8�S�-�7zV�&Kϰ{=RdҢ�B��L� GD�o����cŦ-�,�s���|���L�w0|11��"s�$"<YD.T�TyGF�|�"�ܼF�HQp��A6V���W�҈{p�ن\��'���Ɔ �<���"���j2��H����΄h�u�v�iL�AS�I�18Lȱ���7/���!��X��dc?� W =Y�\G�Z�#޺/i�h%�<�Qz	O~�=��o!#��8�uC]3m�B�;�ܷ_��*�,̃Z0���h�<w��i�Obܒў>��'9nyö��y�F�
�$Ͽo��MX��V7m)�����f�(����J����ELt����ھ{�hA���@Ȋ�A�d�N�S�Oш! C��W&) +͗b��ʌ�Ӵc��(K��BK|�3f�#����t�[?r�� �.�u�<���N�O4Tx�g(A3I��L�&��<�d#�� �tkN���So�UZ#�je�]{�I;4�B�I�w���uBޝG`h�S��3l�t�'����jA�gڮ��I�:	�㌕-a9(��g`��%H����>ɨp� ��`95G�eI�������x2��^��Q��K���T�Vɍ��y�kC�V�\1yq�� m{�Y�� ��y��U����F�V���'$���y�!	8a��A�����tP��>�yR���l�@mXŞ�wq�����y��]E����W�Sr�!����y�F�`s��BTO7E�UC�aT��y�b�l(����
j�ӧN'�y�kG CM@p*Q�\�
���3D��y�Xjj�������KPCȺ�yR��;�`� Ơ23%H2G
]��y2l�3WF����R*)�;���y�Y.�ey��#�qA�;�y�&W�i�
��g��I��!��S��y�DÃw~8��$����5pJҁ�y���~�a��"��v�Q���y�;;���$oD�s� ��e�^��y�L�D�l�b�ɡj��(R��Ӝ�yb�ΩB�6�r(\�kZ\���E��y�j֬?\ܱ���
e=P[��5�y�"U/W����M��[^��ڲ!��y�C5VN��@n�.B�p�؂��y�U>���M�B�hq�lɣ�y"�1JZ��F<|p�ED,�y򪌟qL�zw�,6�!K�G��y"ESO��e�wǷ$Y����.�y�LN"VK:�Rf�����Bc闌�ybm�2T`��f66��z�	ӵ�ybb�K�5�$S�$�I�c�W�y2��>i�F��g.��⣧	�y2�j��b#T�]<y Cf���ybi�O�d��N�	.��
Wi��y
� F)i֪=G�|�����+[G���"O�%�$e��2�����&����"Oj�����'a��U�$nK+��"O�AA��ZK����X<�RF"O2����#���Q�@��o9m1�"O�}!0�0+�Z�E�(����"O�ɺ��17�¸B0 Y��"O|UzW �	C~�d9��z���10"O\�Ifo��k6���U�����F"O�>$I�����?bX�1�"Ox�3�ʊ%4�2�_O^6��"O� ����t";U���a"O*�ƭ��cIڕ�2��;��W"O�a�����PaVW-yR<Hb�"O���M�LhV`���z�|,r"Oh��ĉV�n�PpJ1 �!C�v�*�"OBPS
��r�*����^�9Ԁ�t"O��S3&��=�I��.Z�P4��"O���w�R��DA�ǌ���X��"O���%'�/*�Ym��Mv�@""OH���E�\H��̒�/���w"O��R�h�<Ü)*!��K�,�9�"O�x�˾"0���햌l�6}C�"OJp�!Ƃ�9�vP����"O�ް"O|@�����3��(k���g��&"O��XdB�wN���A�\�5��"OΌ�'��!ZR�ԫ���?����"O"���o���q�S9Y����"O����mMЩ��ȱB�j��"O
�A��'l`���2�H�ɲ"OR���h�&E[v昗@횵"O@=2gkX�+熭Yv�F���D@"O��X7��?��]�1KC�yRJ���"O
U��I�[&V8CJ�uD�,�"O��ـ���*y�ȢB�O# !a"OL	xBL�"V���9w��&t�0�"O�e�'-� 7�<y�G%D����A"O�X�3)D2���@�0��q�"Oj�SF#�*������SrD���"Ob��*��4���0�/�y��|8�"O�	{waŗal� W-��:�,u�3�0wRt	fඟйF�����/M�1SbƄ1T��q���~�P���/O�=�ވ(S6�r "}�ЄضaxEM�bJ�L�س��p=gfȬ7�Q�CH�sr^=��u�'��|`MN�+g��Y�h;a�̕	"�<;4a��H�<�Xq	��!��cC��3d[0VVl���\���Ɂ!؊��K_�K�z (���"����)Q<��9����KN�zg~�!�Iy������B�V�%b���}:��Ϗo� t	] 2cNa'>Q�2�|�˄00.�h�w�;�Z�i�G׼p�LÂ����+�EF|v���p�Ӻ;��5I�Y�pk�;P�Th蠠�)7���;7��
�H�KU
$�R��-?1��ވ	D �f�~��`�+�8�1%�D��e�B'D�k��̩��R�Hb�ȱ�+�V�^�@��X4.~T���͞)� Xj�Gf<��Y`m��I��-Vl�ey"'A�,I笘��(��!YcvL��5r��S1���rt�� '�Ƹ�_'4�t��'��!d��Q�����4o|q�e@L���T��ˈ$��0��f����R���$9��X����2oN���*���]�I�~���j�>��D�@���[Q�g�·X��	�S N6���ե��yF�T��_�;	�=�Ĺ�O�H� �?C�\T��*�19X��4\�C���KL��L�:�"��L[�%z�)=G�Lt�L<Y��s�j��'p�p9�b��be�76,E`�oҺh��0�O:^�XiC�O�M��d�{HL��r'
��0���I\�Ŝ9[U�V���p��D"z��%���1Qmd�0��/}�Y0a���ڡ"� ��O]9 ���7<���FOO� ����18����7|�\ҷ�E���A���N�N)'K%}��(d�x>-�C�
7eG@M���Vʨ"t�tCV���'nQ�����a�R���fBHE���dnʌe?�d����\a�r��9Q����δm�&�q
�4.�<�;�ʍd>���V��E�VA���QG�T6�(B���K�����W�sz��#͠<�耔;p`E�O�� �C�>�Գp��-U�@�@A7k	
����s��
H�R��Qɗq����ɩ94��$�;M�hG�OL�q�iD����>�d�s	�!�@H��N&c���۠�8�L
!�@�f��`�'E>ԩ�b��W
0��3Go�Y8�� ���C�?3RZ�X�2~��ц�?� �k��T7��I7X��	�)_(�N���� �:��@��\t�P�"��-�Z����T�o� �+�^�l��U9�@IS�!]�v�QI�&�z&DA����TʙJ�'Q��t1�&�hţC/�(>��mM�4nL� �>>󨝒��\�P��x
�G&�j�	Z(	=���.J�c$+�y�(�q�*S�zDbx�qB�E�P���`�&1�W$�*L��O��([�)?';(�xQ�\!b&�RDUU{v��(�$8��2&ҭF�V�1E���N��m�c!�#g,�bDL��Pp`4�d�&;��1ZE8�઒,�4[~йgbF&W�"�փ��*�]C��.vD2%�әf0����5�y��P�.��]v�+���X�<� ��08����G��i�uk
�i�Љ��0��k�h��X�0�� -�48�IA>E�����T�n_*]���<|�1㡝:*�T��F�Ӈ8����2е��T�oY&UȣN<	z������$ꖠMn��q���Ux�i�m�f��4Z%��+@a^;B*��4Y�6��3+�u8�+g�I&F<���E�S�F1�M@6�V- ��X.^.�	T�	�H{1� e����šR��V�4�\=��/Z:-�)U�*Hn(`�&%�X���(#����FdnlI�aJ�;������(-Jl6��H:J�Z_w�I(WgU�'2ԃ�'�?k�,:�ϗ.h��r���Hz��.â�|�Q捯A?���$��m�2$:aO��d��������Rx#~��@?��|+���2� ��w�j���g�l� �&�ۥ�D���>��p��2�0\�k�\]N�����_�A�5/�2��UŅ�h�T�(5�["��m�rKS(�ug�ۢ"\%���zӶ��tʗ�=�M��O�\A`�أF[ pf��������5$�>!���k�88�7G�#�H�I��:6Q���(�1�Z���R�*�,�$6���#Q�$�uR��(�&e�c��4�j�ᛦV�:,�Ҧ�~­�@�F��K>�t�!���M�!C��J�Ơ`io�4,��b[;;8<����	6�z�Ѷ*� )&���#B'�T �ƭ��ت�
a�4�	��L6zz�����J���	6^���Y�T��O^Ht�"�ϩ
�88RG �冸��K	o[�q�Є@���4tX�]qaMJ"9�>�p���xa*g[ٺ�pw V#&��`����m^}&��
vb�t'%��`��hG`$�Ly���y$Ι1S%��N��\R�.T�#�]�gB\�1R�=���&�^5I�їz,ܱa�� M��Hr�Δ�8*�ې��
!�ܜ�@B�@�"?YA�]�-�T���0N��!��~�H��#B�dQ��K�3}r��"(Կ<.@�(�E\?":���	�.�XɓS��gV��B�3�A�ū�JR�'>rD�%�#P�����A���	��F�1�e�§O�+�H�b�/ܭp��N#���e���6$��AB�r�� �Q!Z<^���]�ao�Ui����d��@���	Y�f�5 l��.	�i��%4cj�I)��a���`XU�u#��T'r�&$�-Q$�dq&��	5J}��lp�	���Jv|���׫X86��钆'ܡ}���Y��i�|#�F�<]���K$�3����3�2va�ዝw�X�æ\lv�DP4���ʰ���+ȬH ֵ����q��537aI�u�D5P���x�0hG��0v�HX7�Ԃv<�x�/�t��!+!�t��'��I�1�\�K�1�U�"{�ɋ�d�q�b$i�D2Ax}�5#�x@�D*g�X��<��%�D��@M�1&ը��
��=W`qP`�Ѽk
˓Gv�H�*-9�^Z2E��,F=mZH�J}ⵧT)EB�	�B)%��֝.Q�n�aժP�+O�A���"8l"e1�Ń!H(��e�3 ����Vx�����b�V���@Fd=��X��?>���I�l�@��'	�Y�c#��>������f<��p� ^�M;�S6?;k,T!|'�S�BX�>4�3��G�ў�e��C��0��χ�Ȕ��$)S�འR��.dx� CTڌ|�E"�,.̤��rf3��I��H'\'D��¬
,a|�H|��噕7�j�K��<|�đ9�$P�=���4wK�H���Z�1A�r�G֓C��(��{�C�$	����K����V i�LPIJX����	2i�����E7�d	��Dj�>�ϧ�R,q$���QJ�'��:� x�[rhǖ�:-�'N�f�p9ʱ�@�$�x|Y!��O�擠}��H��0-�WN�!a%V��6�	R�����ӱU�t�Uhb��oN�HG6	�`�G�M�"L�C�~����Er����H��	�l1�Ѷ>�@�lZ�� �J�!�/-��6	�J�#!�Ш�b�M�oy���a�T�)�hz&��5˨��Ł��y�T#��D�6�X�@iX�&�4�֊�3��UӍE7��Qkq�� I��(P�Kà. �EO�6��� 1�:ʂa��[��Q{Q�@�I��(X�kC /4�<"�aE�>,�pr��ߚ���c�Q�ě¬�2%��T��-��H6:�y�O<*�h0[Ҭ��ڒ��Գ�N4f 
�'_d�I1(�!�LpoQ g
��E�ڂ &�\40o"b��I��V�0Jb�%?�pF�,��@�%�7|)D$ۋe����J]}K��BF��� &_�-����E�x��$�k >���ꈇm��u)��Ӳ2����"�J��pb�[0yV�Y�M�b�����bKܓRS��N�M�;�v�ɤ�Ҋ-�4�� 3Q�ܡ�O�&���+��'�,3��N�;�jر$Mӊ/�<� ��Q�ܙ[w�����GЎ}:�ᳫ�1�|�z��X��'<J����;�l<�S!O\_��9E��z��x�n�Eޕ��Vf��Ϩ4!R�k�U���kh䈱�L
!�`��Q?uSG�b_�<�Ջ��-*|EC������L����4Y �Xɒb�5P�^�#��M�]��@�5�H�) jq+E9O���P�5H/-l5;�	8L�J��T'L&��h��ō3s�BwI�1z��{")�3��Ij�nR�*$�Q�'>&��m�k(H��ƽ ���,����ݨ�b��C�x�cA �؟@�w͜h-@�M������x����Fb f͸ܰ�F%|��%ÂfA^�fK_	~� R� �T"0@FD��bŴ��O�L@�l��ϞAɱj3A٬��e��
+*;
U��j�m�?_P��(O���Q�.�jm�@�	Ƅ�Z�.�*Z� �R����R��[bn�U9� �V���	�q�����öhF�JȀ5�E�6Ƣ�JMU(i���������}x}2�j�I�n�O� ̈W�W'Uf��f��R�'�6Ժ�-X &�  )o�CgK��p41dFZ9/Û6 ����pѤ Z�$��L+�%X�"4́�,�K��8��6q[��!r��&u���j3��9���W��0��X2w��1S��#hZ�H�<��O
$q���"�e�8���'D�1��H�4:���%��X�M L�f�m��$Q�ib��җ �t�Y c�^� �0e���0Mqp�֙?��(�#z�6h�F僠:��ԡ1v��$ߢq���dO<E0�%D�^a�U&�|�@&���仃��r3J$�Ǣ a�h|�U�=<DzxgcD2~*5h�/�X�����$��p4D���f�pH𭟾x���IxɜaG��3�Ԑ��Oʴ���Ǭ�A����׌y��`�4ޛPw�U�v�5� �9KP�B�i�x�"m�'iB����ٰ�:(Q�kӢq�t-�"1y(=�O]�q�&��5"�����؀d�<d{`�i���P�MI0��ɋ}B��!o������4t���"��#8J�p҆�*�XÇ�ٙ,{�d+6ɉ�'/챑�n��x����BG�`��$Y�BߘN�]˷��.~�Dc��#'⥩dN��M�FDCY�T��@�Փ7��1�c�ԬoB:t�eL�	
�H!�l�8J^�Ƅ[�P��P�U6�����/hN&tp�M�:�K1c��#� �h�ɀ �H��<;4ak�c��$@��̕푞, BΏzB�[�I��❕0�,a7�=8.��w�X�m#�aaS/��uw4���I}N�Q��]����I]�;��;�k���� �Yw�����K�A���=�F�,b.��'v������u�*�;��u[�ˀ�a���B���#��ԙ��iej%h��6]Q�#|�+˴R��	V+P/^�����J:~����{BE]>W�Tk����_�`Ţ��I�tQ��u��5t�CD&��\r�ͯ���䮘�/��B�`�?�����
A�5��m���.h���3�D���팢�M�L��B�$�Еǖ~��LC,[c��xCd�SXszٹ7��6g˦iQv,6F�(�ȅ�֞��l�,e��hk1Ȑe8D��"IC^[&�Ȅ�@��0V#E+�8 �5EI$�Y�+I`4���)�K�,��+��S+�x �������"K<`� ���2m���q�j������.N�~��!,����4h�u� ���0��<!!,� M��e�+͋<=��=�L�4F\$� �!gQ�1��=;���3�˃C�
�4M�1����>��H�2I��� �0�'bL�1�Wk�|��J ���C�Ι[ܓGK�{g�L�D��|[W���Sx04�_�r���X��N�N@��h�CV;W�*�ȔK~���t䞎u?f��*�
Ia�Ёwh>�x��:T�$��Ć�|�����4H&M�t��*�� jҨA�pc���K/,	�K�6�*�j�D0e����+�*�C�~k���k�P0أ������ cT�y2����H�>��d�hێ8T���#�j�X$���Ɂx���1�_	9�؀!T�m�	����੐c�A�XiA�Yy���	am߈;��`��g��S�a�����K�e����
k�,-J�J��~�,TY��DZ$��֋�!b�����(���X�P����ȷ9v��!JN�GҪ��U�U�>J�t�s���>�(AEm���Ek7A�� ��0 º!��+�b�c4��l���;p� !��H�A��}���r�Ҏ8<�M�1!�)�~"͈�Y�z�ف�ڎ�H��IОE:��Ȣ"׎���U�GX3��(QF̂1AWP���@��!?�~$ٱe%�s���� ��1�����-v,���Jت}�ʓ�ޡ���L���g�C��|
��%9���+î�
���'_�U��i�=6��@)!�p��͒�Lz���j��|P� #D5�H�A7,�P����a�'LO��;��J�PhN�
�
�+3��q�AO_�W8���
*���"�ɘ�����=E�t���7n,�6A^�}�p8{P���hOP��@�H��U��
ߩ��'2)؀P��D�9~�Y37cȼmtq�ȓ �<��81f�-�ϓ]5p�ϓqrܘ;3ƛ3Id�4�-O?�Ѣ�y��8*w#@�֍�� Jx�<Q��+Fȝ:PL�%D��#�v���"I�H�wb��0<Q#��9�N��Tę�IQ�D�T�Xe��PZ�L�����c��w�=�B�^�+Z`z0Or	�R�~)�):��ޥ>�ȡ`�"O��r7���4Y��hðx;�l��"O����K��&�F�q#`۷ *&Z�"O�A�� �E����@c�A"O��3 �D���HFE�.DVrk�"O��:�C�N�N���'�gU�Y��"O�����M�C�H�F�9$�2Y��"O¸�a��5�@ q�����A�"O�h�2�\�X�R�C>
��"Of� Rn��`��!R:V�z�"O��q�ȏ"h���zdNo��R�"Ozђ�&��gEL����Q�B"�[Q"O�A�a�Տe�x��Ͽm@���"O�)'�W������	9�h!�"O�d�,:*V������P0c�"O�,k��](X���bo\ �"O�1���r��HcB\�F.̭!e"O>�j@�G�-I�!iv����e	�"O�Q�s��6Ũ)��bL!L��L	�"O29pgdP9.�\��@R>;�V��"O(QV��SV�U,��J��"O��C��.oKp!P�Kװ1�й�S"OZ\C�[�0��Uo�t�.�k�"O���Q�&+z�  �`̬Lþ���"O�0�?E����� �D(��"O��#��H>+�0P�IO1	��x�"O�(Ƨ��d"E�J�0��A	�"O�qQ�7�<c�GE�e2��Q"O� �QP�� r0.���fK�kZ��"O��
S#�����OM/*�La"O���d�.4�|�qMS��Zp��"Ob0���9([��[F�ڋ(���q�"Ol��#)�$s�^,�nL�e"O4I�q%�'$�����NK��Sa"OB(�D�\�����j��
&�-�y-���3�môx�^Iˁ�yr��)?)�m�w���L��yb�ˡ�>�{%���cDf8��&Q��y¯ݣUVyqPK�7,9�6���yr�?g冑+�,Y�W� �r@Y�yr��9H*H,ã�N�mr�GQ�~��؝*{LQ�P@Q�;�ܼ@&(ݧ�hO�����9e]@-�aN�+}="��"O�] �h�n{h�Q6�է(Q,XI��x�L�+OP�\��L�>���$�<�쁉����mQ���
Ώ5�*���^x	\\��J���B|>�3Wϋ�+��k"%�+r�0(��s�����L�?�HO>u���Y�5��+0�� U�x�P�v��S����DA
�ʕV8�T	� /f%���O�Z	���AI@h�A�(-�l!���d�m����^�Of���"I%�j:�M��G�1OhFz���]SCp4�PA��ֵ�r�����T���L�9�*��6φpHM�*_T͙S�'���Dy��I�2��q�c+�"�E+������-Gy��O1����8V�T�;�%H?hx�-{��r����zc�,[A�A-G=Q#e��L�>�OQ �����3`-٢3
r��S8u �(p9Q��|r��K��h��䊀�p�`H��wp�6-7?)��¡ma�T�Jk,Fp� �Q�_��!$e��d��<aXw����\�'TsLA��)k����K��b��K%�Ġ�ēO�����i�)�$��~xZ���$Фx/|hJ>���$x.��}��'Wy�`B2cN�\���D7_)�!�'x��I	n����Ox�V"ĹP�(��_�a$*��F�?u��@V2Oj�)�'�ʠ(�BN^#��	(!�F��!?O*@�'n��	M>���B8���i�N���6���M�6��<Ŏu��)��<ɥ�t��4\�Q��d\�S��=�'�P<ZL���ȓ*�Ԙt���uC��J���(nd��JӬA���<$�Y'O�(GK^e�ȓ���S��ٞ
����S�'�B(�ȓ��i҆"~F���C�X��ȓY�LՒ�hJ6^�����nfE���ȓ8iFU#U��1"�2�����U���+01CQ�W�&�`c��C��5�ȓ10P��.L�X,x)a��w� �ȓG�t��Ӌ�JШG@�e ܬ�ȓ1F9q��rdtEKی<8���'4F��d��(F��i&&K�}���i�'�D�1q���wX����}���R�'Hd�jq�ʊi��Q�bG뮹�
�'��q4�AͤdR��O�|&���'�N]k� #r`���%{��h�'���[�J;y��qYs�C5
*l1�'�U�T�D�U����gŐ�Y����'��C"���.EkBC/O��C�'�p�P,��w�x$tX�'؄�	��[d��'��@[��;�'Ұ�G�M�0��S8�^�
�'�XaPa�ǵG���x3�_	Gt
�'�J����^4:f`MIPj؎|g�q��'z�5#^�F3b�i6��%"�a��'2t�E/V!�HII�k��4�R�''�d�g�\�5Tɪ�%����L`�'�����֜f  q�c�$B����'�(!�X�S�Ӈ'g�ʵI��� c�H�������	d���Ҡ"Ol�C��QeR�u*s��vp�hbf"O����F��l�J��m�`�A��"OR�Ců�=�T�0�m��Yt!	"Oj����M']�6)�Dm�c�A�E"OVL�҃�
���ٰ�%^�B�"O$p6o
q�P�2dq�D
�'>�52� F�!H�R��M#<�R}�	�'\d�E�@�_6�������x�'Q���Pꏘ(��	�N�
~!�'B�A�Re��7�^̙4����Pm2�'m.�R`A6�������:}�����'ʬ)�e�^�H������/y��1�'�f�j &R�>�lQA �> N�
�'ͰUx���:�4� JE8w �	Z�'U������0���9wH���'��ղ�L�g% ��2}Z�c�'�0q�����-(�k�-F�I�	�'D�
C.�7 ��]#�o�+Y(4
�'�8���d�X����F�����'����F \�@^
�x'M	�~�@��'z�P
���I^Yr`H<uR��S�'~�H
�bߏ<��I���V����'����ecF*�B�9W��9y�`��')z�X��ڳ���RUnƈ'���Q�'������5�1hK'���'Fr�0K܈Y�k֎Q*Qy��;�'����욳1�¨���P'z���'k�@��ǈ�*.�����BJ�P
�' �$�vN�*n0�+��؊8����	�'����H�|[ҰS$�M�^^���"O.�c1h�1t�ҕB���YcpX
�"O��쁛g	̑��nY�DY����"O�X��L*<��y�/ܘ����p"O6����yz�-�2d��O.-�S"O*ubc�A<X��ÃC+HV���"O��QdY�v�����Z�1ZjpJ "O�Ԑ�l�;e3F�)@G �&���"O�����~��l�"ƍl�t"&"OTl᳌2+�����L�A����"O�9J�	�N��4�6$ܢx8�dh�"O�)����TG2h	�-\�F(�	Є"O��K<4&N-?kHyXP"O>x�a�Q�Ĳ���:^.
H�v"OR��c��A�D��˘VJ�8�6"O��B)�,X5rA{���Fꤰ�A"O�mK��7-��� ׬+��A"Ox�VoƁ�*tC��)ux<0"O�,�#��&<4�hBH�Q���Z"OqK��Y�l��i���0u3�"O�x���Gt��	"��9�B��T"O��gbP�9��9�'MJ���[0"O�M���-c����+F�8
��1"O`�#�L�}4.�2�Y���� "Oؐ���I�N�AfHT7Rh�pz"O��C�.�*�>!� .BL�v�"O�ԛ�T�	L��r�#7�Dm"2"O.���aS:�0Iz�!B;7����"O�xx�D�t�I�Q�j�D��U"O̴�q�	Â�b��2T~��3"O�$�$�\�� x�s�ћkT�� "O�!6��:�\��X�1X��"O���E�
-\��3��#����"O���Bh�'�1���Y jlYcd"O� @ur0��-��Uɓ��)Ejh��"O�y�!�	�{�X�jq��%��K!"O��Cə0�&$ZE��;�68d"O��C0a׷^ N9�w*#�����"ODP��C�5c�fi�0�"x˘��2"OM�Q�H�H�t��I��L��I�"O�}@!�V""$��S�Fu�0�"O���GK̀ft��`断,�n�*"O�m��$3dh8���&�+`|�t"O@˳$�+s�b��d����"O�eڤND� U�)�R�G�%&zHC"O�a0��ËHz"(����<[6c�"O�rř�9I≛���3�|��"O	����oRt	v&�:C���"Ob�`�ITt:�Y�ņ�6��`��"O\�x�NQt�Z�"���$'��Z"O��i�
��c�j���=P��r"O�I��,�P���B ��� {�"O�<���2�� :���S��Pu"O�<��K�!dU�`�fK���"O�}3�隁�p}K�L�-+4u1w"O��Y �U���;��Z�>a�"Ol���E!bt�Xs	C�vv�l�d"O2�ӧ�>oф 
�h��x�fp��"O��P� A�6�#(�mXrz"O�`��X� �ē�h@�A��"O>]�))Y�
`#���,�L9"OR�B���q��p�M)r$��C�"O�X�"�1	>����2�RL��"OZ�8G���l���sԌ��>����"O<��,
�¨��p�B�cEJ�J!�C�Q�Q�!,'?����t�*@	!��b���B�;i���`B_;uY!�D� DCz���%�F���@��J�!��֋7;z82G@�!s� 8�!��C�bjQ���Ė����5�Q�{�!� *�PVN�B��نG<L�!�$]<:+�,�GA�J��c�%_*.�!���/�b�����,���b��Q?^ !�C	�證C
�2:��%�A�!��*E�`<ѥ��M�T�xL��U!�䓰[D�VZ�t��)! !��#�x�q�����D$�:!�$��UgV�;J��`PA�B
��!��SUr`5�θ��qp���9�!�͸�h���"�8X��Li1�F	~�!��k1 Pnސ?��𳠇RP�!��W�8�����G�/e�\#�'Gkm!�ϟ_X(u�6*F2����7QV!���9G�X�Ê�r���FJ�9!��X<.jn}qpN['�h�)�!�d2 m����:t���9�!�dGz�,X��A�p @/Q�7z!�^x/>�˵��Q����A�rq!�DR�D�8�5
�%�̘S��6C�!�dX�*��D"�"��WU�Lq�B�9t�!�$�I�~� �j��d����&sg!�$�B~��ˀ��>i�p���9%�!�d QL�8�ɀ�%Z���E�R<L!��&��&�ů�:Y�`�S��!��KȰ���/G�X$���̒U!�d��'.(b�B�/Bx81f�ǒ�!�dP�@�X�*��ۓw*��/#�!���%�t*��5@�S.H]!�� pl�@�O�?q
�sjU�}�� 8`"O�PWA�xmp�hG�S�!�"O��2k�46Ӛ���,N8���"O��S�	�1|�3$��/�\R0"O�𲀡�5*�>Dra��]�4��"Oҹ�$DQ��E�B٬�2�"O��+�
ցC�p��wD̎rȄ���"OR]o�\�I_#�,�`"O���ʃ�&rB�S�Į}�l��"O�X��w�� C6+
�F�0p"OTM�u�H�D6� ����U"#"O��H��Ǐ%>��@d��-s4Q"O��P����p��u@���Xex�9"O��%�ƴ\X�ׯ;]�""O�T�N��&0l̈�+ <32��"OV�*D��O�\����߂/8L�b"OH�0�@هv',�Ӈ�X�}��1"O��U1^~ܱE�@-0�,q��"O�9����v�8��2O��T�V�;"O�����P�7��#���bE8�1�"Or�3E@ОK�fqcU�'[�� "O�̃�h�?k�<��U��=@e�eH�"O��q��!:���>p肥��"O�<y4�$&,S�+8Kk��"O"	9� q����)��i�� �"OF�!���#��A����d�7"O���"��#]p� ӯϠb�.�Je"O.�	C�,j��Nߨ}����g"O�t��a�)�P�C�A�(���u"O<�i���L�e����0�
E"�"O�X��IN�u-4iCn�[K�D�"OΨ�d�K�>�l�l�R�p"OH�h�)
�	T&�����w���"Ox	5��3Jk2�B�~�D�1$"O�EѣLC67x���'�q�IpS"O |���?�0�ͩg���e"O�̢�S����4D�("p"O6q��lP3LtN�6d�Ÿ�*`"Od��#�>%-%����FTHH�!"O>�*�-��o�x3do�5Q$s�"OPГ��,"��`���M�I@qP�"Ov���@6$~�a`�㗦o����`��<�	'c�,	sS�i�?�ie��2IH�Ї�)D��8�c�����>��� r�
/Kt ���E�L��냉��'=��p�G�#[�	�%Y�~��h%�����8��)����*,��W�B$V�R$�X>���疾`eTh�Q���s+񤆮+�b�'q��N�����L���+�i�3b6(�QR��O���'�(ҵHC1e��+���?�(n��d���i��4�ē3���q�gÕ�P	"$�Գ��P���|����<y����ʋ�dؙ	�<��!1pʴDp��Ħ.�}���5(W�r��EsԀ8Ҭ5*�'�tїBtމ�%��tݎ�Ӆ���S �M�Ba��m�b�핦d6�E=;�D���d�9{���N�L�����.K�*���HS���R�i�h6M�Ov)���O��6�Y�X�1opv�:���E� �z®�08?@��O怚@��xʘرT W�-¦ti��>Iĺi�6�)��� ��> dϩ4��aєjΖ[��*5�X�Dp��z�^��D�O�})�>@�@��g���j�NA�˟	�>�St�Jg�I���P4Y�"Qm�:O岣<�viއf�jͻ0*��y���bv�Գq�Y�4n�,����􉒬F�������_��U�A �	/C��������\�7*��C	
�zĨ�O��l���?�����'b� `��	F�]Yti�09�(��#�+$���W!I�b�Ly�S���@{��*�;��5h�&rӌ˓{�� �i/�i�����&a�N1�����YM"���O�d� 6�Z�$�O��B�U�XHP���#4��#1lJhB���/ŽKTp`��-ّ{�(��Z�.��x§�	�HT�๱+�I�j1�Ɨ������K�%+V��0��A�d 0��U�
ӆ�ۑ�3Ѯ�y��Xy�G�?�!�i�N�	&(��h#7*�(X�޴z��܊�@��F�Q�L�ǉ��o��Qm �����Iy(<��9� �xЋ�]�-�D���g���M)O�|"����m��n�'�M3fb�����c�ذ�\0�k�Z?y���T���ݺnJ<�2�ӕ5�%���UGGFU�Oh:�+S��%\������
Z�xY�I<ѕk_�'�i�u >k	�����A�����򩝯4$�yf�Y2�p	�	ƭ��'`$�����g�B��.��W���#��T3JQ&xjg�ϼ<PqO��d4,O���4%	���妗�y���ǲi�������ZnZd≠I>tDP�AܫY�~YC��i�xybf�i.��'$�`�A>���'�2�'"���|����/97�  �K׃U�,�+��iuD�pcƛq���)dh�8&�$x�O�� :q�J���G`d�"�6�l���֣^��r���%X9�ჳ)�5U}:��ծp��JC^�5���i�9!;ZY�;#��'�Y3m��!Pa�� �1+i���'J �(�S�矨��¦�����9Q��A�u+�.�9�#���0=�{�ğ v*dGL.B�haӧ����I'�M{C�iV�'P�T�O�I�2Sx-2�kA2p,�R#ؠJT\�	U؟�q-   ��     '  �  0   S+  v7  �B  �L  GW  �`  �k  �w  J~  ��  2�  v�  ��  ��  >�  ��  İ  �  H�  ��  ��  �  W�  ��  ��  ��  k�  ��  �	 � � �, �6 > UD �J �N  Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�� |d��"O
`�(�;���8���-0��1%"Oj4��ND^[��"3/9�0|H�"OB���H��*�ʞRy=a"O�味V�!X��!&F�:J�$���"O,��a
���C�Ą�M�"O,$3%o�-���p���+Ն�:1"O��ݢ1����`���y14]2��i�<�6��{_���c�H�`�fX�$Kn�<��A̼VI�xR[�)�Ć�pඤ�ȓA5��('nߡ4�� �)˩%� ���,��r�؊b#`T�eT09���ȓ!�b��g��}�8�F��-? �ȓ
K|m�ș�VṔ���2�%�ȓ"R�X�j�4JN�1�˘X�i����̹	_�jZ��1!g��zܶ��ȓgil,*�J�
j�Ne��i�J%b���f	�(U��:���G��$Y^م�~r�� S�%T"���k\�jx�ȓ|4�1�îJb��@ӵ�ݩn�V��/[`�"�v4�R�!ʎ<��M�ȓ`:��z�ؚh�J�Z��$HY:	��H��p�m�C1��!��B:��0��EnjZA V;9����J[
2���	��4'J�EA�IVW&��~�(aZ��ӹ�>� o�Y�|�ȓ�f�A�
Ο7�H��M�$�����mޠP����/���ANXo*�ȓTv�����{ ��-7�*h��I��sB�8�8���3����ȓNe*M�悡;������X�o��!�ȓ'lj�#F�m�+R&;�|��2)n�C��0S4���T:
b���:�0!��e֊��)��ͷV��,�ȓ0�&�8#���� ع�L�����;�P�AFd���,w�6d��r�EQ�( �gVlɦ�M,H��,DP���|�I	$G#\���ȓ"�)���E�B	yt&B�^�LɅ�4�� ��eëF�ڙ��n��R�p�ȓp`@}bŇ�=�$�AUN��P����L��p���_�a�)�Y�!��-��u�5���o}�`iF�@A�p �O��Fz����ٷ"��#떏*��=����y��Ȃ!'%8����FV��y2K_�Q�m� �,)�����-�HOf�=�OSb��$I�\� WI�"�b�Z�'�6@����:M�f�.d�cL>эb�ӣo�
|��.R5/,��ȓOݡD�C�@<t���b#,1�dK�n5ܒO��=�}JYI0����DE�rc*t���-[T!���%�t�Mb:t�A�ǔ>!���/��T���V.[ft:�e�N�!�U�BX<���yT��cΔ%xqO�Ї�If0H1�T(G:�@����-vb���3�G2�5�D@�3��2��G$�<)3�'�5���ƅ}���!`��/&�I�J<�����4ϐ�^
	8 �I�x��A�'-v���'�F	+Fd��R��&mR�*��B�'$M�L�4AL����.� :��'u�,�e�I��n`0'���.`�'/2I�p��]oZr�CY:'���;
��� ���7"�&���k�
i,r0�T"Ojĉ��fg�X����)]����S�>����*�I5��q�"�q�t�x���2z�C�	,:8�
& ��a^��`th\�@���O0,����Q�n��Q��8.<-�3Nó1�yb�6��0�V؂Qă	}a��" �*B^������4\O��C��>ow�%%�@��'@�	�;"��s�aW*2�
�+�#X�3�������$|Ojh�S��NQ�uCS(ʕE�|��G�ɍ��?� sǏw�|)�O>%ǖ�	��$D�D�1�нc `ە��ix&�U��?!H<	�����dR�v���WI��DII쀤!5a|�|"���m����A�:�1 �S7��' ў���E)��*ntA�'��tp�D�I��HO�S-&���Ђ�/f��q�O��"<��?V��X#ʝS��"�H�����!�	�qb�zp@�s��0Sy����x�Ɋ2)��0�j�%<s3뛸>C�I�L���� � `���`�eժh_�B�ɨ+�,0ؤ��I���A��@j������O̱)���̡Ȕ.ʐ�*�8�"O�m��� �	��Mb��!�ղi��'���I�x?@�Gh���80�,Bs�b� $��b�� xİԲ�M��S4t� �'�B�I�w��ɩ�N�?����Kʭ?q��hO�m~�NVe������Y�x	�r�똟�y£'-̨�:�B��h�5��⎬�OP��A�yҢ`��/����s⡃'i!��	'0i��K�,��}���˘+ !�d�O_��F�V��ZA"g
Q�!�DA�X��t5��!A4��AJ�!�0
A�I0eF
�}%�	���ĜMy��)�i*>Gt��`hY`r|@�S(θb�!�$6�h���)l��Ł�)�!�dR�4�D� �M�{&	�%"B-�Q�DF{*�])�˃�e���"!ILi`]�$D{��/a)d��C���-f�HU�J._@�6��<�'��)�3}�+h�|��dUJ�j�	��Z���x2�6�Nĩ�⃹G�d�b@�8�dz����I	�1R�L��A:򤌼&h$��d���x���9�[��B�Sm�#�\�1� ?9ٴ�䓬��۳e��d�1��]���@��QC��)K2����ˊ8O:���`��Z��B�ɞ~���	�&y]�X1��Q<CF�C��
x(QF�ʩ.��\�#��k��C�	ݦ��&�}�
5	 �ڼrC�/D��`�U�4�����Bڔ��% �gU�듿?	+����&�#8��5p#0�X�3�MIH<�Jȼp�B��z�9��}�'�ў�l�J�z��GD��'<
i��F�0�'�;
 =�V%���b������}�'���?|�8ل&k�9z�'��%� H�K=�(RQ�T��~X�'Ԭu{�����q��:#��'��ِ
D9Sٶ]�M|#�Y��'��Qq�h]!� ���V�u��Jϓ0D�O��R�&�#v�|5	ѨDh��	2"O���Dc
!/��#�.�҈yI��IJ>EQ��v��@�2J�9sh�C�O>B�	O�r��kX�[5X-�W�,�n6M�V?��y2L�~�J>��$fz�h�*Pl�(Uj���\#���J'r�YTϝ�l�,�AFV>.�`�Gx��)���/:L��E�s]�q�nRq�<��$��͚���RP�u�ǥNi�<� ��B2m�Qڲ�G"j��`�p
O@`q�@������$ �(K�"�y�+�+0e#g���x�n�0�b��p<	��,�n��|�Ea���;�,0?bQ�ȓKY:��E�X4I�j�g���>��*��{��I��2P�t�wi�=唵���9(@a{���@�e��j*�s�p��ƈ�3ў@��	"L��}Y7�ƔIgj)��e'�!ډy�_�"~�	4'�l!�C.VB���*sC��<hd��Xg���M͑ ��f�B�I3#u��L֦�� �J�r��B�	o%($��lݜn>����
٬B䉤Ak�9	G�\�b[���D F��B䉸(�9��&Y�J^�)�偁����5�g?�֩E�8G�����/�,`�+O�'Iv#=a)O��	T�Q��� ^(S� �
U"O��r��G��X�Oɚ�P�J���TH<�2	ք$�)�%�%BB�P���'Z�� �2qT�q�ʉ/��Ij�'" d*����zA���^(n���'*��a����~��%��暔|�1�'^�=)�w��	���K�j(	�	�'J�Qqsd�D����Bϗe."U	�'v�����ʜ>�����<:���'��� �/_�7��������'`�a�/ʪD�4�XC� }@�y�'�h�hG���!�@٧�Q��:�K�'UZI�d#Y���J�E�y��I�'-��@\$����c�F�}<�H	�'��备+~&����<mz�!Q�'�`���W�'�(S���R�4��'�(��	܂seP��Bn�P��xC�'�B�h��7TkR�#2�В9��)�'����%Ȓ!�&Ȱ��ڲ5'��Z�'�0X
1�3Li�ጔ7$ڔr�'����Æ�B��ś �R�e�}S�'K��8���P��K�$�3h�x�
�'�X��� �1e���X#�&-N���'���:B�YZ@�#�4c�3�'Y����/��]D��
󄀺]�B1a�'O�2@�#�v�K��1P��\�'�l�t���
YN��!��Er~�H�'m`աB+vm�� ˔@^r�'�����瀷]=\ԓW=����'tiҠDެ@}D])�fܧ/Y�8
�' �I 4cċxf0!�$���|���'�RL�Vl�.D,�dx�)�>�T9�'mCE"�(N˸-zp\���l��'D2p�!�,RB�i�A�;5����'�T�q׍�1b�*��G��.4;z%�
�'KP�C�c
�t +�:>�K	�'�R��ʎx�����Ş1���i�'�t������8Yc��!T0��'�ZT�Dg˖Lw
I��)Gk�65��'P�A�A��!|���{ ��,��S	�'���	��OH|s�H�6,�xs�'�X��W8��l�RbH�(pR��	�'U��B�J��f�ˁ�_%�.��'U`�$(^�cLt���p�X��'ed���,ʻf�E*�)�kR6h��'�J���gϊ1u~��g,0!��'�ڑ�' ŒcD^r��+0�X	A�' h�X&��,R��#�\.p����'�6�u�Z'cђ���Ǣ6ƾ����� ��Hr%[c��qB�K˨nj&�!"O�};���-ƮISrk���jዲ"O��F��� <��p�@1�p���"OL�Y!��W�� ��E��^�.Tʑ"O8HEg�,D'���ߴ^�~�	��'~B�'_��'M��'
�'���'i������WN=��6>�4u���'<��'2�'���'-�'���'	����+ٴY��	5"B�	�ԭr!�'�r�'.��'#b�'��'N��'�H�(���I[�mQS�؃{�����'���'��'�r�',��'���'��}��j� �ǥ"ۢ��W�'���'V��'���'���'�b�'�N��'U�=�!q3��]��a#��'0��'��'!B�'4b�'���'%~���g�[x�t���C��B�S!�'b2�'��'.��'B�'�r�'4�(�F�1>R����*����'��'<��'db�'ob�'�"�'���b(�O�r��t!^10·�'�2�'�"�'""�'7��'��' �%���ǃ�hq�Q-�?��#v�'rb�'%��'-�'���'���'l.ɣ��z��Q9��O(|�@ G�'���'��'��'���'���'��L��c
)_�a�ui\3!N��`�'#�'���'�b�'��'D��'-2�!%Ɩ_w��A KI���U3"�'-��'�2�'���'��`iӌ�d�O��h� �����.�7�R$��`yB�'��)�3?�t�i� %	ef1�:���ɠ���R���D�ͦ��?��<I�i9n-���?j�����B}×�v�2��ЫDV7m;?����#=F59��"���"+`t�%e�g�J{wl^���'�b\��D���t(iЏ�>Y�Hq .�;ƞ7% 1O��?i�����,\#�(m��D�6�
1ŜI��&Od�`�	v}���bB�Xʛ�;O�U��D؞"�W���|]��3O��)7`Ϗù�0r�7��|"�G��DS�.�����I�i���̓���#�$Cڦ�pq�$扖(=8�JF��[�2��燾t0l�?fY��A�4e���:O(�.Mr����ܞ�j$�"�mWq��I]�V"X�̺��$��
^��
ןr�F{r�����*C�lЈ6�DayBZ���)��<��i��:�e��9��̠�@�<ّ�i���+�OJ�o�N��|�G� #}e���KO�n�,�@#S�<�A�i�x7�O�J��bӠ�q�l���cRb�0�3�Ƕ<�4=p��u�2�JgJ[��hO�	�<QO~*��ܧN2u"���E�,v'�x~�ea�t3W�������aD�&� �J�c�z�u1�[s}�v��lZ�<yN|z�'�?q��Q� TX!�f5&*��8���2R��J%�u}�nD]��u��-�뺣��>������C���7�&�PO��lx�l�GA؟�'�	X�	�M[ �<�@A�i����U�P��>=�E��<Q��i�b�|��yb�u��oZ��hB7��v/l�a�	�e#bPq �R���n��<��3@a.�)#����'L��I}���vLٖ$������I7[*t��,q�h�	Ky�Y�"~B��(��p��cH4F��08g*FZ̓K��v�T���$�ЦY&��0��"o��oY�$;�J�<��O��n�M;�����۴�yB�'̨�vg�M��h�Q⋼H���r��>!��	�"$ў�S{y������R��;T�ؠ\mp�K�<!M>��iY����y�R>�!.�6J"%q���+,.d��`??�Q�d��4>5��1O&��I[�s qj���]�����Pl]�A|R��uo�I�?��ׇO#�.���g�JMj�:���x!���p���?X���ΕZ�r�h�������0��b��,I���l	ġ򭆦3g�ɕ�Ïn͢a�U�юeOf�SG��!!z�B#��~(�AgfS0f! ��EJ';��A�'��9A �.Z(�!D����̫���G��a���όj���r���Hh���+P��|�w
܉*�`=����S�Bc�ĚF�8mI�� ���[&�I�	�>���&X-N<ɷ%Q�(���z!nE�d@�%��E��vG*�i"�L�7�����ӎ.������6\@���z2瀘B"<Qe�_����y��x��'x��'N������7$ hh��-��.r�5��EH3����"�G�	�����ɟ��'�܄����k�n�dǒ>t���-Z�Y�m�F_���I�����vy��'��(�;��)�=yH�H@@�i����'���ȟD����<�'L\�S��7��^>��i�JO�S�咁ǾI�Ao�����Iay2�'d�8��O>
g��~�4	Wz��)�4�?Y������#j
\�'>u���?�X�_��1c$�%t�4x��E^y�87m�<i���?�@jḩ�?q�禕�"�b���x������q�@ʓR?���!�i\��?	�'h���?`�Nx1͝%8�(��'��)��6M�O����<��S����ē'���9���eZ1$޶F�Vm�	-��ٴ�?���?�'W8���4��:M5�PCĮ�<�"���.^1l6�نB����?�����<��� ]�%��K��M�J��	�9�c�i���'B#��@�jO��O"���f�F�`�i�����˕!�?}"4��'
��'�
�s�y"�'���'"R`@FHŵ{D��Q!�S� �ǣv��.J���&��S����	DyRH��}��k��J�_�$E��dʤ/ 7��Of������O����O�� �2LpO�|u��IfjMZ9\-��b7t�'���'��_����ǟx�	� v�HA�ϨM�@0v�W������Z��?����?�(O�8"`G��|ʤ��;� �ĆW�E�v���h}B�'���'��I���I�YDh�
P�pVA�;o�DP�(()L�'"��'rR�4�	�(��'=��K�G 7���p�\�%�Qz1�i���'�˟��	�7xc>��c*c]�Z��&;�`�ze�J'�M����?�,O�y��Hq����s�=[�\�S�dt�Eˀgh�W m�"ʓ�?I�'��0G�t��M�'̳j�����V3x�a�女�'�R�a�m�H��O���O��Z�Je�n �Ra!�o�P��n�h�I)Z�2����i���'�* ���Ý��q�a�+^�Uaݴ��Ap��?9��?y����4���ą�B]z�	� �?���,��i�nڨm^��"�?�)�'�?��FR6<�b�r%�:h�҃�\?Z��&�'���'.B\�WZ��Sϟ<�Im?�r����ʕJ���"Ftּ��^P�1Ob���`�c�Sޟ��IE?ARjC�V�B����Q�b�zqf�ݦa�I�c�lq�'���'����Z1>!���G`TnTH�6 y�	�{���X�L=?���?	)O�$2o��Ty0�L�{A��4iM�<����?����'2"��2�L��Z��F-Y�&·}k<<�Џ���$�Ob�d�<��-���S�O��"#n�0j�P0"�O�G[� �ش�?1���?I���'E�m�s����MW�+݂	��6P$�(RC�^}}��'�bT���I!Z�ʘ�O�����gG6�����*�;D���۴�?��b�'n�]�����5U"\xW�-H���z��LLTYm�ҟT�'f"̔--�S]yb�O.HБ��Z"7�Xô\a�'�����N�x��c��'=��D��F�x��L�A �8=n��'�¨H;2�'W�' �dP��ݿ�5r�#w�np��b1`v꓈?D�Ϣh�v��<�~�r�N�R� �1��C
cyZP2�����:e]͟��	ɟ���?�����'ZbE��@K�FA:��D�I��х.{�[rʗ�}.1O>�	-C,�P�m�6��� ��u� ��ݴ�?����?�0a�#��4�����OX���9I�\�Dh�?ƚ	8s� �pʔ�c��Fm�S��L�IG?���>O��f�5\�h����a��5+ ��'v��'����FFR�p���;.,���j��'�����OB���O˓�?A�d۲��a�#�]� W<�s"��,0��(O��$�O�D �	@?Af-D=D\�)�4�Ȭ��!�F�M�ySpg4?���?�/O���ސ���SC�4��'U�q2�T�{��6M�O����O���'29��4Oh���j�GW&|��( ��Z��'2�'/�	ן|+��D�D�'XD	� �?vH���߅*�b���g����-�	ZyC :�ē.D>	����<!3"H�r2�z�r��<��l.\-�,�.��z$dH�
P�e�n���#��F*�OJ˓xh��GxZw�����F�=C�F�Zt��E���r�O��ė:P����O���O��i�<�;��WG�>ʌA�1�L!L�6��'9�	&=g�"<%>�s ��/F�:�� ���"��0�7�x�`IR2H�O����O����&��|���.��5ib`��u_���8<q�PPVR�P ��0�S�'�?�b�N�d`!!����,��6�'�r�'���h�T���П��IV?Q��

��%A��@F��qRς�Z���kK|Z���?��'A���'�?�	0�$"`U��4�?�rH�����Ov���O�\��B��?$�p�WgԠ\���D�>y��2ŵf����џؖ'A�aL�;����VDտg�̲s�/���]�������	s��?1�KB ~[ �S �R�� ���L�z�@�B~��'��S���	���d�'H�^(9�ؿg/f`��'	s�Ym�ɟ��ԟ$�?��8��Ѩ��Mɦ�¥�^:8��=��
Yd���v��>���?y,O�dY
~�R�'�?It��#b@l	8���t�r=(��>s\�V�'w�OH��Yj,�0�x�V��|`���I�B����M���D�O�a)�|:��?)��n-&��dm��>F���s��9�Hv�d�O��+�`L
N�1O�S=�&|�0�*@��u0Wkҧi�*��?!�X:�?Q�������Ӻ����1S�$a�%	37�T��n�~}2�'����OŻ����O���*�Cۚ,��B�	+��iڴ<s�U���?q��?�����4����R�Ov %�VW�&�Df��>�H�l��0&<%�)�)§�?� d͂/�X\TF[�X�𥐿*2���'�B�'ELىGT��㟐�	U?��
�7G�<�E!�	S�1�%a� P1OF��6�D�ɟ<�	X?��ō�n�D��J��JE��*�GC�����T%@M�'��'{2�ę >�RD�)U�2K)@0}��']d�U�bf'?y��?�(O���αe$�`aΟ^m�J�������`�<i��?Y����'�"���N��H'bDb@�/WK��xT?����O&�$�<)�f�΅R�Oh@mE�kdj�`�O/ƭ��4�?1��?a�2�'Q
̂F�ɥ�Ms&��)A�����D7��<�E
h}"�'�S�8�	�t�Ȕ�O�b���Q����׮:y頕P����g��6M�O��L�ɠa��Yx��:�� �Y��ˋ%o6��;�3Y�l��6�i}bY���Ʌ"���O�R�'�����`��th�C�8���`�	CBc���ɀ�1i$N6�~�ֺ'��#� �;6���{v\h}2�',|�'���'Fr�O�i��C1gN��:�����>���"��(�*SZ�S�O�$�p�ۤp�x�W��7ɜ�m��p�������''��^����IF���s�}��@�� \Y�D�&�M{�P?pd���<E�D�'��AIW(�i�D(#W�1J%���Ӓ��O���	]����|���?Y�'X*���`ץd�2�شO;z9�A�pJ-�I�),��1O|Z���?�'�$�KR��w�e*��(�X�;޴�?ypa�2��d�O����O0��"wAۍ �|�V]5@-����û>���5mT��';r�'��	ϟLQ�Qu\a䥟�J�z5iT9�'o2�'$���OD$��`� C��	Y��\[���%�ׯl
��Ӗ�������	}yb�6Ux�S��=�^	i�M�={��-��`�.��$�O.�;��O,��_a�@���KԬxG>@��(�gk�6e�,nZӟ���ןD��zy2`�i��7�O����
v椨�VI�����Z
�0\�$�m�̟��Iޟ\�'2�㋑��d�'���P�����b����v!0#��to��'"�'gҌ�c�7�O���Ob�iF�B���b�%/H���2?6��m����'�� ��D�'�b�F���ܴ_u`Pc�l��9����2jI+I2(mZ̟�	�/�XMrݴ�?���?�������g�d�B��)#y҄pa�,5�Đ��R���$O��'j�i>�Ӻ�1�D9s`����X�=�d�;7n�Ħ���ϝ�Mk���?���z�'�?a��?�P.
�Jގ�����4Wj�Y)A�S-C�fD]�`���''�i>A'?��I0o���D�R�̤��� :"y��4�?���?�%Û's��I^y��'����z��`)J*Mp�e:�K
)/}�6�'y��d���)��?a�z��h�N���p~\x�+U�i_2�L��d���D�OJ��?����xcU&á����.]X�'���k�'���'^��'X�^��iF�蚸&a���8�b�B;Q���OV��?9+OT���O�$X�>���B�/�3A�b���ߊ*l� B69O ��O����Ox��<I�!�[���?<��ZT�L*�"7�75_�6W����}y"�'���'/4���'t*�:S�FE�&d��ү q�j�b�>9���?�����$Y�v�FP�O&B�F<C�%�(�6�V�3�(��6�|7M�O&˓�?a���?a��<Q��~��R|��+p�	: ��W�)�M����?I*O�i� ��i�$�'h��OlJQCV�ޥ1az�X��R�p�� ��>��?1�`׾�Γ�?A(O���P���� w�� 1�H��8}h6-�OB�R�L$n�֟��Iʟ����?i�ɗmyt�b�ăI�(��2�ڠ5"�Y{�O����=����O@�V�k�I0��m�>����D�,�*8p����M���I� :���'�'n���O��')򀏝1��y���f[jU�b쁒55v6�P�d���D�<QF,�|�K~b�'cۆb5��6o�(�`�4ffx��i�b�'�B�µ9�7��O@���O��$�O�N�y4n��F�^k���{��)K��'��ɬ�6�)z��?��y4Ҹ*���)F�eI	,_�42�i��� +�$7��O ���O��$�d���OBx:�펮R�Hz�e��TѡQ�X�"�u����Ο��	П��L�����h������>z�~$��e���vco�����O����ON��O��	៬�I>y6�4�d����Â�ԭ������	�������8�����[�&��M�'oF'��-s�	ƅS
��M�N���'gb�'���'G���Z"`v>IV�A�|�N��b������̮����OR�d�Ot���O��@F��Ħ���쟰�w��I������
:6�� ,�'�M;��?I������O\�"�<��'�l���V�2�<�ȓdӝZ�\*�4�?����?��Y��1�i@�'~��O�`���o�=�A摵\C~8âe�|��<��/[�D�'���|n�S������Q��pHP�E)rQ�7��OZ���t�ii��'&�O����'y��v��<8�8�cˍ0�\,�4�>)��U$����?�.O�i4�t'�:xԦ��e�t�\�IP���M#e�'c�F�'q�'��t�O�B�'�$�C��'q���R��tp7MC�Tp��2�4�p����䗓5�����6U�h�a.�2o�ݟ��	ӟ|XF�^�M����?)��?��Ӻ;D%G�NH�� ��gsr�R LU���Iɟ�K �Q�P�$�)�'�?����3��V�*9*(��ŕ+�ll���i��A�B�6��O����O@��B���O�(��J�N�d�I��8H4!�V��U�#?1��?!��?����?�� Y�A\��V�"~L#�hx��i���'N�'k��'���O���W$ש���6@��^t���ɘ~,�D�<�@ �+�?����?�.2z�"�i�N��I�.Wڡ�W%��4�����d�����Oh�D�O\�Ĳ<���>9(�ͧJ�"4�c'�� �T�ږO�>t�bR������I����I�c^D��ߴ�?1�;v���:o����n�2`"E��i;��'��S���I+&�Sϟ��p���6�e�T��dN��M��n�������l��>o���P�4�?���?9��ni�h�)�f*�}c�'2�����i�2S���	(jJ��M�i>7��B�C6��r���!�#Ov�V�'���ۣ6�p6��O�D�O~���j�dO}G��&OT=L��p���]o�<�'���]'2�'��i>���� �%[�,�;&+LAr�J�+�X�Ƴi.t��e�H�$�O��DꟀ���O����Of$�lC�My$�� �)Qzq�Dɦ�Ȥc���'}�q��O��O��t�N*O�4@�]�h5��Q�P6��O���O��K�ʟæ��ʟ��I�i�Ƀu�ЧVB��ZP��C.�P�w�jӬ�d�<�����<�O���'\�)�"bK�����H�J�0F�V�r�4�?qD��nJ�&�'D��'��L�~��'�L$�c�t4��7ED9����4��q*EW�<���?a�'�?�����<i��pČ����;�cH#H?�Pq�J�IП��	D�	П��ɀm2����	8�(Q6,W�:�Ĭ���h�\�'pb�'�bU����� ���d
����rd'I&��Մ���d�O0��"�D�O2������Mv�pd�!��'~9�;Bh��-�<�'��'�2V��������'�t�K׌ۥR�Dc��&5�iS�i�R�|��'�"h�>�y��>�u敫Z#h	�b�6<�.�a��Ħ��I��'�jAs�5��O ��+U%����(��y��D�cn^��H�'�������kp����(&���|�;�G/_���� �\{��n�oy"ަ6�n���'f�d*?A�E�8�^����9�l� WK�������ڦt�D&�b?-9�eK?jt�H�UaL'?�Z|�6�y�\�k�mVԦ���� ���?-�J<��-[�t��/y�eq2��>��d d�id��x0��S����g(�V�j1��¡2P�TW��Dl�ȟ4�	ҟ��)���?���~��lw\��e��1������I!�M�I>�Ѯ�<�O��'��#�3�ؙ����>Z�1xb[�&�7��Ov�2�@�y�	��h��l�i�ix�D]�4CY�%��uɄ�>��Д�?�-O��d�O����<I���-��Y����7�� 9���,[�@%u�xR�'�2�|B�'��%Ζ;ǼuyrG��8b$��}]rE�c�'s�	ş�	�ȕ'�^@�WKw>�A"�-֤	A(�\a��h�B�>����?�K>���?) '�?���K�ؚ����?!$�3n�!n�	͟�	ԟ�'�*��vI$�	��yy���ϰ h]p��I�hm����%������<!�O��'���W,{����H�,$��4�?I����d+ �<�'>i���?�Xf�rȰ�Q�j��t�@,e~b��'���'�q�Rm��*^���A5��v4���i��.c%�p�۴%P����x����></#�$�)U#�а�f�
IH�IIy��'������u�DYrL$ H��� Y��o^)/�7��Op�D�O:���q�i>q30�V#0i���DW�Y|<���������Oj�$�OV�D�T�'�����ETE�`�iЧa=���!d�����O:�$�c��$�O��'�?��'���rP�R�UK$��Ć�2�&�}"b�Ƙ'y��'����!5\�q@�(��X��G����'62��V��8��,��?��.پ1��-K�
nZ�Kâ]?8R���O6��r���i�������LyR�'8�P���E��A)�H�d	��"ڰ2��	�P�����<�,O��3,M06Hh���
�:��/k�m*�8�I����'^.�4��ɇ ?�J(
�
R�),� z� �y��FW����g�	xybΞ�W��۴\����e�T߲ b���%Sa<�'���'��џ0�:*��!>�� ��J8$&���E�f{�3d�i���|rX����CǓQ-6O#2'Γc��d��%�^h�zнi��'9�I�K萱�K|������(��37�� ��Y�c_vpMozy��'��k:�~�D� U�~;C��Q�=�q"�9���Z�0#� �M\?��	�?�9�Of��J�(F�iʔ��d��i#�i��'��\���T�'����Qh䵈�a؜^�,�Q�gV����U��ʉAD����uǍ� �AX���\��3�O*���I=oO��8�$�H^�aE"O ��i�:#���a�
��\�J2m��z����"+��p�@M��>�n	J&k�07���:����,,
�o��n�V(Rf�R�L��ч�΋0�2ybC�'o��(T�Y�mr��x���*,���b��Y1���Ʌ,�B�"��-{�@�0�B@H�c�Y�,\feЪ^@�ن��O��D�O*��Ǻs���?ќOs�M�� �F��iK���64�V9�vf�'�x���tݐ�b��;�p�쐊L�h�h�'ژĪH�< �D�['�DQ�9�dA��?ٷ�'AP��7�ȥ^]���aR�E��j�'&>��-Ή���!p\�pBޔ �y��#�	(�����O����U� I��)�#-��5q���x���O�����O��df>	����\��pw��?H���ٟ5�b��w��;�$���ַA$�x��� Z�28�'�B�k�đ��+Bʽ�g�
�+�����m�$!��I�+L��d�O��o&TɓE�͝�������#�T@�<�ߓ���M�-� �+c�]H�H��o��@H �%sFBJ'n�~ ãI��y�S�PP'�@�MS���?!+� �j�Of�V�ԏFkЙQU��� �
}�v)�O��_�b�Ɯ��S�����i֟�'��I�a���
�U�F��Q/F����sD��&�	a��@��ar�lQ43a�Ep>p��[�|�Q���1P~]��F<}ҪM��?��y��� ��g]O�C�G1v�$Ũ "Oؽ���ׁo�N���n�Ϡ�Ҁ�'A�#=�P�
n,�l�!��RĪ#j�����'��'4�<�QO���'EB�yW�_�S�ȬA3�B}a"��nH�4�{G��� ���$�#:�X� @�|"�:���qB+O)f��CF���<�� ��L��<�d&^�D�Ɋ�L>��<j�Ei��29����BmQ(�?1�O%Ae���t�	 �h!�%�Zr�y��75'�B�IM]~�[0,�$l8�� d�/,�������'��|�	f�_ {��|*㯚����jBC�Mk��d�O$�d�O�;�?�����O�Oj�`����(�U₁���ڧf"�PȈ"�?�y҂ρ{°�KR*}��@
����P	+ƥ�fɚ���p�r����I�b��)Xpܓb5�5Jb��U?�a���>tʴ)jH�0[�s:ܵ��f�+���J��4^���ȓ*��\�p₶n\�p�`�É,�L�<I��iX�'�dI�t�~b�g/�ɳ����Q�bL�PtN6���?����'�?)������1H���3��D/�H
��i��\��j��u&��􂖩&���t%�h��,i�TJs ������ W{�|��^��$Q%�a<��SHZY�$�=���� �4Y��	�|;M5��b�T"���,_>c���mx� �C�S�0*d�0Dʽ��Hwf3��a�4S��iW�Z-��J��������?�-O��#�J�u��󟔔O��=��'�*���ϐ84� �Kɩl�c�'a���T�r�T>�u[p$S�w<#���4%LƘ�O��S�)��P��q9���'/ä�s��JT
�'Y�Ic��Ԙ��O�h�ڦ�pɱp�*Zʐ�1G�a�<��F�\��T�oƜ����(�[����DF�	��Mլ�)��؃�ߩ2| l����Iޟ؈�猣:H�������ɟ�^�����/xIN������<9�d�@x�Jf��?k[��C�/Rв��%�	�c���$�5"�IbS$?T,��ôe]'��1���Oq��'#��S��+�b ��F[�4��' tIjaB���d����Q�O��Gz��I/G(M��G5aY����!�'�J�"��u��$�Oj���O0I�;�?��������Y�r��!��=�n]�∏b�T�f(�-,n6��k���y̞�~Υ �E_�]�`ܣ���r�,�[�fq!��6k��D��b��0��aR>��=��ʧc�i	�,(����L8��l����?��B�z�D�+�ML:Ԃ��H�M�<ɰ�ҽ}��WL�}ZD F�21O��oZP�	�!�tx{ߴ�?���{�D[agR+S�ք�+�w�������?�@��?!�����_0?��0�w-R�H�nx���)*'����A2%�r&�W'\y��d#�.gJ�@e�T8{��p�LGxT�X�JN�o������l��l����B����֪A'(>�yPM>���A柸XM<a�gFU�� �� �UNn�	�Fm�<�t��jC��K�˛+`pѢ�WP<9��ixP(4E�]����S�S�}Ϫ�Y"�|��Cè6�O��$�|�����?	�P/��lR7�]��������?Q�}� �bMc�0qD5�*�F�'>��Ր�h_���ЉG�E�cF�!�O���P�  �B�;��V�#��I� �Z:���2넫��4!mѡ�
3Q��8ږ�F�1̦��O>]q��'1��O�y�E؄`�<d�1a�"b�3�"O�8�4I���������(�֜��'��"=�i�!u&8-Wl��{�D���E����'���'H��h�KE���'����y稒5u��XK�ƈ$@�������&���r���. B��L}�5)��|���_�L R�͢A�L�7��'2��6Ȑ�6�S��p$�ɓ�)�I� ��w e�b��\��+�7FSx�#'0�D6FW��L>��	�. <xIҬB�mH��;`�X�<	�3r�*0܇M1�E�֫�T~��!�S�O[�*�m�:W�`���9g+`���Q- iL���'���'zRMzݝ�I�p�'d����D��+����A�K\u��&Sf<����	�:�V���3k��IC��PB�X��
�:X�+\?.a��BJ��|a�� ����������[��ϥ&�h� �רu{�B�	>a�`��o6dj��P|��b����}"�h&6��O����E���5���s��2�E�>3���D�O�x�U��OP��s>�����O��O����ַC��	���&A�)i��'�ЕC��m�-�h Q�D߈3H��Ca�N�p<��D�ӟ�J<y&gէ8���q�W�t����C Uz�<� ܹ���8����Y�-"�i$O"Dm�3
!�L�"��
L A/D�t��9'�h�S� �M#���?*�bt�w��O��1��j���C�Ƚd�\�h׌�O8��L*�F�;Uȓf�"��2(�]�� ��O/��b���s.�4^�Z�
�FX�~3��'��+, ���� ��,7MZ�VĂ8����lם�Y� H�"қv�N� ���0F�v�'��̟xhL>��&�9�Фp fL�Q��Q4�K�<Y����!B	�蹻j�A�4ي�DƇ .2��$�v��94��+xxl�䟰�	�4�T��5ZFH��ޟ�I��]2wCx��.B��R����|�����/���C��N���G�r�g��.�<���� 3 ]2 LM�-d�U+R,N8Z*�+`a�?��Ba�ܳ!���OAZ(�ņ�3p�Ϗ��z��y��(��g��'��(��S�g�ɨV��XP���(��y�%�B�	>�(���`���qm΍e���J?���k�ILsp�
�C2�$��G�h�D/�Z�*`��ǟ�����^wR�'�ۦnc�ɱA�G�EL��9gH��\�w����pY�b� GXN��V-��բă�Ly�q����$�6��d;�����x��Bch�&lY0ZS��a�{¬��0C 
��^�>������05�A�a¯��h��m�à
�ߊ�	�m��yB�O)i�� �b�EKQ�����'��6�-�䍎�t�mZٟ��	�^X��ʎ|,8�1�=Pj����ssbC�����|�L�)7Kv��2U�#<���snK�M���1k�"�\��Dd[+8*�GIH%�J�<i0+�;��Gf�|�I�D�Ʒ<�ȥ��Έ7� a���,96زp�'�d�<�QH���hH<䫊;D�H֊�-�ni:�BUx�<���Cm�<�FɈ=�j��pu<Yp�i��=˧�Ů)�����)6����|B�;$8�7m�O^�D�|�.�?�FaO=;a hp�R=o}�9	��+�?��o������򙟄�,�#Mp㋀�<�\
��2}��[�O���1G��"A�' Ź?lt� �>��O�ԟ���4{x���'��r)#������N��U#��
���O���$ʥ���CMH)+���R@ C%ax'ғ%���7�;a�8���Y2}֚�3�i���'��b �����'F�'���wp�Hx�Q�t���au��]�p������1�ԅ��W�e���>j�p��|&����!�"#�9	b������5o@��玳�4��Qgټv��5���#�$��@�5λ[�@3Ѓ� W{T·/$�|
���D\_I�O"��ֵ?��ya@e�2M��`���;-�!򄄥p�|ܻ���0L̙���ۂW��(�HO���O˓fI���7�J�s������	csR	R��>l����?���?�'����$�O(�ӇQ���ZҀ�/	[D�c��oRY�bD�5@�X�e��6��ae�^�'���gO^ ���&l=�]!��H����xeb�]��B$�ֈ2�џ�������l�s��?x�����g�����yO<����?1�b��\��e�V�ֿrI� �'����y2l��l��&��g�5�A�����'/F6��O ˓/Y$y� �i���'�aC�
�:j�s5�T�����'�2*H�QR�'���ǂ�{����j��}�����,Q ����:	�C�' l�H���8#~���G

7�A'L^�{�T|0�/��WjΜ��"�N� �J�c���閑|bʈ�?1��x2$W<5��E��懷6M�9���yS�[�|ɰ�Yj|���d��x��lӂ�w�N?c�+DL��k$�ɱ(��L?K�m�ҟ$�	M�$��K��X�;,U@�ɔS�(��e����'Q�X���->�yA�T9"��T>m�O��%j@f�J���.�:i��`*O�,zA�Q�C�DM藈�0sk�<gE�/0I[ʞu��ID-W�:��`W�4[�I�!�.��m�`�I���S�'q<����	.��1'���$~�T�v��@|��Gŋ,��>OB Dz�똼n�Y�/X�� �bU`�����?���E��% 3!��?����?��Ӽ��b^#6�
|q"��a-<��$�͠M+<5J�)�e�F%p����L>!�/�؀3&���^�;�D�s�D#�,�
 ��A�E!Vz̸gFs��ѐB^J� �w#���ʞKr�5��M�:���k�2Dm�ܟL���Nӟ�>��?ɰjÈ&ʱ���gz`�9S�����xBn�&��H7D�J�z�KM�.���WO�'`���'��	�l���+��X�t�ڠ)d��`��uR�R�p┽��ȟ��I��#\wc��'��)*|�&�POΚ^h�"��-(sv@1�A��
���g��=��p+Q���s�Έ���D3m(a�"Â6�j$i����=�dk�CRxKpȳ�
*�`����C6M���Dɨ�O���D�D�	�a�q���Z\Q��"��'O7��Ox��?��"��K�U0���(1Ɛ$q���'R�}
� ~�cs�;4�
x�C�E `vx��l7�$�Ŧ��ش��d?W�]l�˟���)k�@Ibi�2j�����ʹI��	�	П��������|r���!E�=�@�
"y�`1�۴�X,�k�y�z�bЉ�c@�܅�=#,�K�h�>V$^����,-n�0H�Zx141�3�����F�ߦ�� O��6��T�'D�OZ�%���r�R!�$�K�-�8%��,D��p �O��}��M��C��p�)��ܴt48�a�!n�#��!����I>1� �'��f�',bV>��&��͟�s�A˂_\�aiW��>[&��!P�����	U��|�E%D�+��`R�aF�?�Oi��. �H��d�4�6��w��v���'}��a�o��$̈ɠ&cU{66��D�m��xqҨ��|
 ��&������� B|0��U��H��I���(���ڻ
(��c�K�!H �� ��αd!�v��P�d���"�!@Ӯ��K�ax�j5ғ< n���	��G�]�4LW�3�� ��iV2�'�b�~]Z�[!�'$"�'��wрI���Y� @���7E�,����B���ˍ�d�6�27��&K�1��O��Ye�M�R�@`�{�:h�#gfD@`�06eƀ�m@�w.hd�V�~�ڴ8��u�;a�&ܚǅ��W���[��: �|3�i��ʓ�X��)��O��$�O��Q�n�$W��л�BX��\R��%4���/����]ا��N�� e%?AG�I�?}��iyB�,z�r��Ө��5݊P�u�K�
�|��'Ϻ;��'���'�p֝�p�	�|�sB4P@;�B@�O5�{��D� @��@�p��eJ)7����d�xPz|���Xb�\���[U�W�'1��B��;(u���Z��M��#��kI���=�1Ç�\���w�^�T����0	�ze��	Ο�'���	̟��?���4��#���@�MI�9�B�>��,� ȇq��u8P�²4�>c����4�?!(O��
�h]���I�����W>?۾Ͱ�	�9{�`�!F�U���#A����	ٟ�Χ�f�$+T�R��X E�ر�Mc#NM=3�j|���s>�̐@�e8�h�2ޛuk*y�@��/��!(\Y�D���*�8zȱ3�)����
JO�Z���D��n)�h.��*Qtl�"��G0ԅ�3�_6x!�d�,�F��1D)}��ء �ӘVh!������B�Јp&�TyׄN�1��Ji�&�| 9ش�?���� ���O�4;wm�; )f����_�N�~MJ���O&�d�H 6�uk�?"IR�Z�_��'��)�?��y���@NAh��f�L
95��Z@)��'R�|1�Z�~��!/�k�
A@�h>���K,���*����a(e�$}�U&�?�r�|��H͡5��@����<(���FD��y�k$�9�=2R��e�0<ن��	@!�C؋l��@�hZ�S����ش�?���?	���s��2��?!���?ͻ+爍�T��1� p)�g�7 -Ļ��(v	f�KC�O�B@��b�d/��O. �' m�|
�T)R.�7����ܭ`�>��4f�ͦq�@�$t� �{j�e�$�ă[� �λ�vdjG�N�~ \�@�-M�O9�a*Ǻi�˓lkZ��)��O����Or$�֧D�C#�>�T�QB� 4���#���4�6�J�H�s�0?����?��I`yLÎ0������m� Is��Q��y�M�"�X����E.dD@��Q��y�f73:��d��X#$`�D�A�yb�@���J�*��G�����(�y��K���V�]V�|�*�	�/�y��4b�H����р���!��y"�0 �T�h�Za���&�y��?�Jm��O_� -�J�y��S��FxHT$O�:}�k�2�y�-Td�Щ���ӵ9`R%�w���y��ԩ<�" I��^cZ)wB��y"Č�H����\�Yj�, �C��y2NO�t8"oV�cU���/�?�y���}ňu�rW:��� �^9�yぱ����g� ?Ț��g�߀�yRL�����#�jU%:NP(��K·�yrC'8u�1�����[��0��[,�yBg�/<��Y��}A�L�B�?�yR�wE�S!���T����I�TB�	zc�9�q�B�3�`�aJ� A��B�ɰQ>�[�LV$5�J��5��:"g�C�	�%bF���NXgL���e�;y�dC�	U�෣пv:�|BVGMTC�)� �$X��å2{�!�a��,i��� "O6�������9��ˀ�^PJ��c"O��GU�u�|e 5�Y�<O`)�s"OƩ�%�U���G	,C�n��G"O|����C�u-�1�hԛ���6"O���/<�� *��R�Sd P"O�{�S.Yaδ` �4H
f���"O�@����'@-��O�*L���"O��ѥ���%1��kH��@F���g"O0,�̄�/yHE8��31R:U��"O`�0��8|��Pt�I,A�9C"O&	SWD�K�P!I�K(��h�"O¸�DaN0��,�0K��,�z�"Oba��+7.�a�L|�T�"O�ő�f�)1�T�(��Kdm�pK�"O���NE�d�X�����6>�5�R"OJ����T%i�J#@4.�a�"Op�#�D�=5?2|[��Q�bƶ�3"O[ �	�6Y���7�X�I�"OtPb��V?a��Ē�Z*��y8��'}���C�*Ũ� ��]!���4+&`�q��E=z̲TE�o�<I3j�\?z׊_@{d(Dj�l~��V ��R��&�Fl��#o񟞤���1c�����ۖL/�X��'�2��gI\�g�i�OR�wy��{D��F}R��dEKC~����z���F@�H��&2��Đ|��Rp�t��ʅ�ҴuM��O�H����m$��bI�+=��h�""��dD<-p�B�Ǖ�f��YZ� 	QF�ѶW	$�\Xhbb��5����$��@��F��"TL�ᡂ��LB AL�!Ei
D&��R��e���y�i @.��E�=��T$O�{d�p�n�]����Nš�
b��5:��CtF��J4�3h�"�G^�S����@���@��(&q��c�H$Ѕ��y�
H��;B�QW, A'�6�0>Ad	�r��!q�̼˱�
��]: C�?:eB�ΓC8��a���<��&U)u�ܜ�g���4r��Κ,"�Q���Dte�]� $+~��j�*�u�T��2��xh�E���<�g�S�M4���5C��`�<�eحz�*��ģN�Y;�(�=�U/݌]���XhCn��R���ud� �קzS@�gR��N0���1@q�U�td�8�УW�SL��9O,1A�u����5����^ �S��J�"hR,��&}��>�ХZ$��c��`������']����gɅ� `"Ꮏ'�`9���ω8]�'~���jw^�����X�a�*\F��9	�U���n8N �b�C�x���HL�k+n���B�'�z����	~dQWK%7�Q;���tVb(��.O��y��w���C��$R�s`��D�i�R�R�IX�:�t9	
J�����B���Z�>#<1Q�×x���p.����������T�,�1�W�,_:`�c���Z]�<�����J}l�g:����Z%���:�G�K �xrrIؾ}��ҵ��0zAx�y󄛞VW�ؑc] �(�����sϸ�kq�Oy2��R?9FE^�B��2/�+ �~����.��$#�H�/�R�nڭ�,=�F�� ,ȳdmN�4ܸe���,4�I��  ���kK�'����H[�4�� ��T�~�M4B�J���$B)c`�(B!�6=�0����>�2%Ӷ�f��i�+!ړd�Lqsg���(	���!"&a��������Fn�xÚ'�8���O15KE��f�&" �t�c9�LyDi_?��H�%2�X)0E�2�$������ÜV�~�����la{�KD.i	r����A�#���Aa�@~̓'�����A�����-P,~�jpL���s���.Ас ��t��A�,�����=yո�C$�R%H�T!�fH��n_�ԉ-`�uäI��~r������P������ %0d���J��ߦ��bN�Q��%AD��ѡW�M@��O��֍N �Rp�d��3
��u�Aɏ!]h44!�n.j9��Ye����y��UrcI�e ��a�5e@��N>=k@��Q�_��x�Ԏ$�hO0���C�*p���@�L�O
YcQ
�(������f��O��I�3��	�p)A#o$Z����A���6�O�>�dH�#!D�(�E��T��Y�'3ܡ!Eň<'��BU���w�4e�2�O�r@��2DN�� tn��xH^��	d�N2�~x
g���$���?�I�-i��a�
�D<(�Q� Y	9���as��3^���˄�;$��D*V���:�Iŝ>L��G
i>�cw��s���R��rP×��f]��BY�'T������(=l7MԮO�N	)v��?>��Xᨖ1�D������7#P�Q�%*d�]Q�M�l}1�̀}��Q�D��%p�0xҘO�R�5
,x}@��I�|]q�H�����d�"�VXf�ˌ������
P- ��ɿ5���4��0Q~��"���hC�#�y6�]h�Ȁ2�Z�uap���cͧb�c����Hr+�=��6-�!�Vjo��vd[>s���A�Nr�'h6�J ��)^yh��NA�E����a�Ph�h�	%)�R�)M<� [���;	���i.�%?�9�,u��{0�_�8��逶�Z*!ڪ�ۦ���G�~4�%G�>[������-��7mҟ&�d���~�� (l��I0h���$�P�l�HuZ���ԦI�-�v�8(��
� Q�#��$X�Oژi���C�jD���K!��Pr���Vx�N�O]�7-�6T��=��O)��򨜻Rp� ���m�v� ��'������I�Q�"3���2�=����(1<Ec��R����pI�8]$V��O���qh�I�>O�'�)�T���9>	S'�Ũ��Ir�4A���ٻYi&�*Ga07xĄX�c�U �,"�T�3;�m�Q��. ����lw�4y3#�������k[�d(�M� j�?%��P��)1�4Bކ
�vٳ��p�zy�O��L�b�O���ԃX�Y�$!��B�63ּ����kܔ�!B�36�>�k�k�)>qh�25�\�*4#��R�v���:��d��( �Ѫ$��61@�@���g.̭B�4^�Ԝ��+�W ��tĔ��"���A=���q�,3$�Y�Q��4��#=$N�X���0G���[E�ڲM�����e�y�'�y2l2�)�@%�2Q�� _cX� mA�1" JЪ
Wz-�1�0ړ�8AlݤLkӭ$1�|��ă�,�N�pf��,N ��+߅;A,苂2O����
c.��I�?Y�T�ԯ 2�L��3A����<V�t������t�ۀ �!T�(�Ok
��wϛ*dHQ�%������{����Ŏ7*i>�2�I�8m�7��邾e��Ł�2?w��
E�O�+h�����5:x�	0K����U���
�?p�W�ֿD;d�K��^G}�P>�P��J�� 	���&Dn}�B�I�qp���K���ֳc��㵯0`��9�`�8���'yJDJ4▨S������.}o�8:�U�@+~�zU`�97�����MyR��3c=o�5���A��N�Z��

H��0Z'I�8��õ��I�'��谆
��5�A�!�D���9{KR!G۱3�9�DBŒe���7$�<	��)U˖�IH��O:��  $[^t��t�T�)�0)�����{�e��Ú�v��谭a��ě�XFNy-��՛�m8:��#��'�Nx/��������?��
�Tڐz��]#z��ք��z�Q���O/� ���*)�x��c�%Z�a��
0��S��'��9w̪lN����}4��CD�<9QhBP����20A�����{�'�8�)T��9�s�HI�P�C���W�HH�\�~2�~��C7��)�&``�Λr���s& Z��d�ſs�Сv�'SN�I�iH�N+ek$��oTx0�ݰ�~�P����'�U�
A��
���؟t���F�=<>�K��Q��e�ቃl�t�0凝n�x}H� Ӄ���<�
yʶ�C,y���3"�������~b��/.��q�>�3���2�n�r$_5jv���E�\2Bi*�䖾h��T�b/Y(�P�!+$�?�ɍb�t�a� Ԡc�g��%�T19��2eKL`x�Ě�j��Z<0�A>(l��bOE�)(F�Ol��bGu��I�GF�s���2�Y���� #�r�[��F0z�0��dY�ZA�����%�]�C������k�<�2t�۴�H1�N<v�ɽ�~rQvF���L]�IޞLx�(3k�m(�������g�a{�U5<�p��D��}��)�D%2Ѧ�K��U�rw�dJ���OLU�t.�����F�� (��O���#�����Q�Qa���!�$\��d�!��?q��[giӃ��<m��S�*��G��q����MK.���>O��{`�H���ڰ��ssGIK�'��$y�)�htJq0P�T7M���
C^�gb��B�'CENt�$;}�g�Y*�pE쒗Ee"�����ȸ���
�D.x[P.2�O
����4{�3c�|�4T��@X��$�(O�������rՂ�*_7
�>\B�e�*%:a{B	���MZ�L�8e
������]~v@����jƎ�c�5�ɱ9������vA����-*F����_L�P	�f	�eu&}� ��ۄ��8��a��  B-H�e|�ԛ�-��g� �Ӻ�0ϔ�r�8���)H�#XT1�e �Ns��T�A:æ��CA�ם	MepDy�@�0i'v��n���R��/ė���rjG n6��C&E!yB}�M|����ghV�j������^�@n�r�n�.;)�ɲ����i�͓�D�j��T��8u e����O<�J`�F��̃W�O�5E�T�i^<�q`[�Rت<"q�7;t�}��g=O�R����أ��C6~k��:��?x�0� ���-%�$s�.� 0`���2Z��V�ZgirG��?����2]�#cg���
\������
���6L#_��p[��"���Sⓧ_$v0�p�S:`x�7�?��x�Aj�~��y���ӣ���{�lU�M48zP�C �1�am�>-NV$��
�r��Mz�c>i*�엕������X����b�� Cp�Rj�/�=���ʿjF�0�Ӽ;$g��C<���@d�5H�NIf���C��;�뿟@�q�X;���O�.tU>���,T�w�E�Y0���+���Ra�'��ͨ�����^��K���g�ް̢�	�b�-r!��$N�16���,��p��� jߋbԙ��O�>����N�
EZM���sLщu!+?����?Nf ���>�T�%?�Os�P��n��G��e���6{��6�5Jj)�I��`q�o�=��g�{�t����ka�.��t��nȴ;%t�{��S���:�P�O���q�`OAqj���>I�č?W����V�p=�;u� ��T/�8S8�Y��cɠx��:	�	/TG�@�&�?�1�+P�U��'�R� 6��?	��VL��/�l�b'5O�HJ���"��|C*Of�i���E���R��=OĝB�`؛��,R��'���� H�	4�����O��P���%M�%=L�J��F���	������s^ȓ"�e~R#=}*�X�qуF�F���G`�71����9W�h5�Bk�����=��g�#w��@cF6,(Hƨ@�8$�$�P�*Of'?aP��)\��酤C�� �da�Z����"��|"��D�� *�1� ��@FH��L�Oy֥
ųi��O�I�W����hƘ�H�BVCTr�c���	��C�ɯh��H!�b�}UD����Kf�~C�	V��V�#er(�K1|�HC�I0e`I���r� ���Ƈs(C䉨\O���@/�����ŅɓP�B�	��b $�8����N
<T�B�	=U@yaCL=K�PŸG���,��B�I���YRM�'��Y�&����'�Va#�	Â�a[�c�T6r�'R00Z����l_��Ad-9�����'�,\`Q��5��6L�&-ԑZ�'�|d�Щ=W~�C��/��x
�'�l���Q�~�X��&ׯҒ���'�����05����S!����1P�'R��VF�}h��6��L��'�l�Q�(}S�q�'ҷ5t�
�'.�x��M�{�`�8Q%M*�T	
�'���l,%M���!ZH}{�'��p펪!��rUL��i�A��'���m^]%2�C��Z��p��'�E)5�A�e�:<��oːV��'J�$	�Ͻ1�Ht���K�� ���'҅�f�v�B�0�.�|�bMK	�'�T ��`�g�Z1�A�G�ƠZ�''�N�H��K�h��8�'�����R /K@$�V�Z^H�
�'Gt���DҐ+�N��@U�NCR��
�'N�q���3	]�P��b�A�F�;	�'���mU��8��3� �	�'��ܒU`��<��c���U��A�'G^e$n�5zz�i���GP��'����5F�=5�&�a��D�9��3�'�25[w�	�(� �;�IG(F�nq�
�'B-��N�d�f���@FZ��	�'$���1�K%`��S�-B�lX�'�"!�I�WS�H	��ބqT-#�'e�Đ'  "3����lS�|I���'\�Jq�Q?G.Hx�BF�{4t ��'��awG�3�pcR�	W���'s^�`��o���B�N&!B6�0�'=p$�&��{7�}�@��mjB�'tԉ�K�2!r`���\���'����!��U����
�"�B��'Dؕ͎�Y!�1+Cd��.�F���'���6A���B�*&S���'�^,�'�R��$ �A*� !�'/�1i�l�>^���΢S��4B
�'�$��c ��(��7A�L�v�;
�'%�0xS��	Zn���7���'`��
')�
�R\S��,z؈h�'=�Yg�? �|�'��w��ݸ�'z�4'�$a$&�"�.�8_5�%3�'���"��K�c�>�:V#J��8!�'=r��5O"�I��Y�
���'B�4��+�aP �Q��1X�(��'L�Xyf���(İj����ל��'���c E�Ҧ	�P��1�����'w�	Z�KF�{�,k� �5*����'\.�rP�B9�:<�`š%D=q�'L�)	UmJ�c�KAl߾-V�'h���pMH�h��怄	�(*�'X���CO$6V�lj��R�p
��'ljƩ1/�q���~C��*
��� ��H�A-e$te��� $�0`��"O<�s�*Ҩi�ʔ�� 1y�)�"O:!��$@N�|�@ z��@@"O���&LX�4[$�����X�b"O��R0���q0yR�+�:6����@"O��	6`��|Q���+K8Y�v��t"O�"Єy��A{&֦n�*���"O$A��W04A<��1I�T��(J$"O\����Xtp���Ղ�%[����!"OFip`���_���9��h��E�G"O��,�!\�Ν���y��I`�"O�� ���p̾pzc�Q�g�𠩐"O�i�EΞ!a��\J"��lwZ@�"O����).c�q�&KY�ɫ�"O�i��"@�A��m��ʈ�2��Q"Oz|i���.��m Ul�%R�Jd!��Fr�*���l��-�DՒq��lS!�̚`�,%D3d���z�*�CR!�$;R�x�Ө�^���Ʉ�o;!��	1B����v����q7r�!�$�0�:�PF��4Us�(��U�;�!�M��V�av�D��>x�툕^]!�پH��t�K�d� (@��[(9^!򄘃}� ����n�f09�ÕG!��`�z��f�
�X�$:!��Ҳ'ƠMP�*N�G�����//�!�X8y��brF�
	LAz�+;�!��5<����r&�ɘw�S�Li!�$4>��Ԁ ���vD�A���Z>-f!��P��36ݥY22E��
Dd!�dOHC
�� *ɇ$Cz�u-\�"^�&�)��m
b�M�Y!��I�F�<�|�!O-D�t)`gΚr��P*g'҇W��u�+D�HH�OY~��0����Sz�Ȁ�
7D��9�I�</�j%�]���
teL�~��O���$�/H dR�F��Z�Fa���/��}r����T$Y�|G$�C��!+��r� 2D��uCڊ`E}�S�\#|m�Z�/D���wc�$��	"��1��q��G"D��اoL�p(�(2�7gu�{�� D��R�A��9�h�$��9��O:D��#5����� Q�ۦ0��{��7D��{c���C���Ӹ0Ap!��j��B�	4g�#��|�yg��/U��B�	�S8�r�(
D�	t�˪1v�B䉫v��X�TK�}L��D�%p�HB�I�(V�-8�C�*��kU	�M`6⟘��I�Okڈ;�C�Yp X�!X�C�	�BV� j3��i�r�Ĺ��C�	.���p���_��|��@qшC�ɭdĤ��!�uz�D �I@!�6�	X���� ?�5'��lA��A��.D���g�h�q��ᅦ:ب��K+D��p��I!�XI*J��d�Pq#(ғ)$Q?�n�A���c��-� �8��T�>VPB��ޟ\�qO�p(�)EL�*nQ���~�R)Ez���i�t	��$ܬ���**�ARߓ��'q�⢨;Y���Kb�P��'��p5��/f���D �C\.�
��o%�S��T�5����ꙬwnN1��P�|�!��ьW���bd@*�z|qE��<*��=E��'�Q�@ŕ%a�,�#@T&�@�'�V��t<���8�Bٱ#�r���':p0{1�4���V�� V���d��TD�� �8yA(�PD*��q��%�["�'��O2�}�^4��t�Y�G�z�A%r�@�ȓ
�@`�c��4�\<#A��x��z/r,�B�8P� hA�@N�d�V݄ȓn^��c�T�R5�Њ^�K����*�y۰ȞNʜ����B�&��ȓ*h�{���1T�>��Sa��J��ȓ :�LR��W3��٢�E�=;5���HeP`�d+B(�iRC�=.">̇�m팭�WI�~�����{�$D��;� ��T�S&�Rys`N_� ����m�ΑB��@�U�&ݰ��օ%5�u�ȓ2�r��C �;Zb2t���DM��ȓpҨ���̮+���2��|wdE��	@�I	&�L�a�̈́�NP���� L�z��<��m|�Lc���`�SC��݄�/~��Af��'-܌ Gɋ!��ȓ4���'`-�hXwfU#�ȅȓC��-P'�	Uo&E��D�G���ȓJׄ�9���	q1`�%�-M���ȓ̴��װ5����+t~�ȓNlB!:j��u��	B�%z��F~���v�������`N�T�vdI�Td$C�	�dITǕ2@�@u���ɵCG���/D�4�3�� 0r�J�ɺGXQ�D'*D� K�)J�@<)0��:Ur$@Ъ2���	�U�%�-��E5��W8Z�˓�0?���^?�v\�C�� ��y�f�g�<�tc�+	z����g��X�����d�<�$�G����C)�:b�N�(�j	xy��)ʧC�8���@��fʄK7K�=����i�0���Do����ʋ7��o�O�������yϐ9�4�������'㈛�yr��2a�Й#!,|)
&�܊�~R�'m� A"�-l̨AA�畷T��ay	�'*ZmS��#����D��y��'=���N�kͺ٪#f#?��@Y�'C���.M��Q;��H-|�q�'����@�!"��`R��IGj����S��!�:'|漃k�3|���0q��C�<�3M�Ɛ@ Ů���Yx0�IZ�'?u��jݡu�L]��j���T��-D�hrt�M�j���&��x�ޭ1�-+D��xV�q�#�Ne���t�(LO�㟴��)�9�3D�/Jb�-a$d&D� �e�����%Y��T�R� Q�7-8D�C���4[~�-(�^/mH,
q�7D��0�K�a�B�h���e�Pe7D���C$\U���e��8��� Q�2D�;$(�!4 �	�d͚~���C�=D��!$F��99�a�Qj�#U2�R�;D�H�@�_�X���Ѡ��1S�2�Y׈+D�,��h�+ST��3SD׳W�@X�/+D���b���ڑ���.BLe�3�3D�h�ץB)��q��B�
Hy	g�1D��KG�M�D}
�`"<iH1�0D�`PtO�-V&t �Ŵj �`7�!D�<�1*	�e�(Q9!/�i��2�4D�dq [
ê$��B�7�𔘅�3D�4���A�xj�\H�&(mߺ�J��<D��;�"G�r�SW�@�%��i�*0D�@R`l�x�0c��X�/���8�$��x��;2|���A�!a�ɳe���y���;�	�.��`�r=Rn���y
� HT���3�A9�œ"\k�,8�"O��ٷ�X�grXUsVоB_���"O��1vm�)��C�b�LT��"On5�f�I�Yb!�7ѬI2�	�"O8� �C�&�f�Yq��s��<T"O�AP+ȴ2�b���+�Pּ�F"OD��u�C�q#\�*��M
{�b0W"O�!�uoݕ4��4���fWK���y�	WCޚ�kdÕ~P���b���y!E�5^y��+w��赯ތ�yB	��h)�թ%��m(�<��Ź�yR�4��$�Ӂ]���@u���yB́�d� `��V�}*�H�B�y2���)%�m�0$ޤ͖xy�K���y2�eҦ���ߞN�n�'/��y�c�IÞ�{0��.>LZG@:�yoΘX�����:q�Ç�<�y �2lj�gӶr�j��C��yaܶa�:5�%��r�,m���L��y��Fye���;�(��b̀>�yi��\	�%-���ZA��$�y�$�
6J|�ȴg���%��G�ybCA�6�6����q�%���@�y�#R�K���FUA�4���U��yr��kvL�طJ\'��L[��V��y�$rVNŊwMR�H�����'�yr�X�m�` p@
B��XPQ�7�y��2!=�Ek��Q�@�TQ�$ԃ�y2kT�(�Y�W%K.?L���ʁ�y"c]�4�`4j��3l�0�����yB���4��� ��1��y��ybH�}�X����W�*� �
Q�y҃ùM�p��!M  � �!ߋ�y2 ��~&h�j�N�h���X��yBc�� )�`z�&3��R��Y�y��%5�z��gʇ@y�2���y2�,M�J����|j�߸�y�-3l�Y§���3�Z��.�yrD�#������x�M��h ��yrj�%%8��	��U'wYV�ɕ9�yBė2( H@��oقxkF$�y��]�������"y��1٢�5�yBm(~���XFl��k^���2ϓ=�y��k�N���DhW(L+e�Z��y2*G�4��!�L��NW� �����y�C�3'"$�T�����Hd�ѕ�y��Fh�a�GO�
<Ƞ��4�yү��e��(*Q&��D�)P!���y��P�-�.ے�ȸn@�����y�-�z����C!yT�����y�hɅ<�v���%��rD�ы6jI��yȋ��nx2�$ |aą`B��y��Q�JT��c�mHwB��ug���yR�3X���	W�EѤ�̱�y�
@��9
�gG��ʩ$F�y"��3�4ě�㜋3�hTs���y���0*V�:��mYQh�y�CK_���2���cU$��0���y�L�+p�}0e1W@`���L��y��ͲH"��^n��
��yr�׵���ʢ�U:^el=�7����y�+��tC�l(�#��`�x-���3�yb�њO#��"��C�[��a���C��yrfF�9N�ӧI��M)գ��y
� @]X�g7w��F��9;��[d"OН[��ݭ!"�Ls���eR��g"Of��j��
��:���Kr\��"Oέ*Q�/1��Q��8f��!d"O6	B//���	͒��u�F"O8!T��-eI.�Q�J^
��y"O���r#L�-0|	K��[�F0q�"O�YQ�CS��VLнe�|x@"Oڰ��������b�ˎ�B杰�"O��P�ȱ`N`�Z�
�0��"O�QP��!49�01�;4$$��u"O`���cK�臯F@<8��"O��r �u�����*.��"O� �K#��� ��J�y !R&"O\<!����u���qg�u��"O�ٳ�� ���kfkΩb_* �t"OH-���T�S�Q���˜]��� "O:@$�3 y���'ؼMhIy�"Ox�b����32b�Bg@�b2��"O�ݻ�F�Bb�P��;u��Tr�"O智�l�-z�<�۔o\,�\��5"O���̄�:���0R�Q�L�&�r"O�A�.�1� 	PP�ߠ!�~�ó"OL�p�`�1pݸ	X�C˃���2`"Of5ɶ΂�pаQ�	`�l�C"Od��A	�h�F�81��X�Bx�W"O���4gM���0��D���%s�"O���HҺ�@�B
�9��p�"O�*��E����.Fb���J�"O�PJ�l�(�ҹ8"�g)3g*r�<i�)K �����%�8D�1�Tw�<Q�M�h!�a� �>�V�%IHs�<���� �ҽb��^-H�D�ЄAW�<a��#"h��C�+¿�niQ�.�M�<Y��W�l��y�bD"(x�)�C\b�<���\�gB��t fo0�S,�V�<!�%�/x����!�d ��b��S�<1#.P���4k�
^�4��{"h�<��"B�����TD*Y�Kgc�g�<)��ߢ7q�����;6�(��Cg�<�U�]?���
,=���We�\�!�H�}P �J5��z~����3�!�P�}\�=�0;^��&��=�!�X�:�� �'�ʠS�8P��b��g�!��v
�PqvE��|��`a�1>!�$��h��H �埒`ǈ�"`.!���&�f��&[�F#��Z�/T>!��/q����%c�0 �i�Q�R�!�DV.kޤ���n��N�F�!�Zs��(�X4IO> �'k�!��B�"OԵ��MƇ,O�ts1���!��;�Is ��:�<;`�O&2&!��8Z��6�#8<�(��N�!{!�䐝HO��1ԇS� �h�4)�:g�!���3!~,�yTj[Yl���J���!�$�( ���Y��UH�� �3,��!�dX�&3�X���#7L�m����*�!�� іUBԂC
����ٙP!�DR�K��u�f����Rt��:>!�dM�ll�����2�
�I��)�!��4�{�`�1`��s���>�Pyb(�,z�̴�@�U+`��Yb0#���y�C"���$	�[�8"���yҪā J�4O�Tӆ�2���y
� �!kU�X }�v�XQ���7W�	�f"O��� �М)î��'��3G21��"O�����
���+ �m7�"�"O�в�7)�<�P�I4Oq"O`]����)h�컁��$Y&p��"O�=�u�q���Jg�E�{����v"O�EQ�$z>�$Q%��/wE u��"O��Cq�!i��H�ퟵ:B~pP�"O��k�!V�� �Ц�m\t��"O�������^��4�%��ӧ"ODh�r �,d��	#J�N�N��"O��Q�_5�l��0�Lv5txg"O�]x�P�L��蕨ԁ�PF"O��jV 3�X�x�B�K�2%9`"O����S�-�r�*	�a�j%��"O��a�_�.�N�ꥨ:
�4ɓ�"Oh���!T��j;�LR� �N��F"O�b4ꜝ~�.1"l�_���0%"O��#Ȇr�6m��śD��H!"O6 ��>;	x��i�}�<�"O|��k�9^Ζ�c��&tx�"O~��eg�<0hԅ�!b�(X�4��"O訢f)�V{���G�jIKuŁ��yR��6���BE��s���(5ز�yb�C#��iC��[�܃�y�mٲs�qy4�X�*ZH����R��y�#A9]���MF���:Cgҫ�y�a!�8�7�H���B疊�y柤oL��G�ڥ*�x�bb�Ʒ�y�MK�#�(aBP�%��\(�َ�y��h��bf�	�JW<,(�����y�.S�L�r<�nߜK��(��X��y⮏4f���p���"3Jf,�Ӛ�yҧ�h JR6���p����yr,D>ad�!#��;@��2���y�jH$e�8���HGIk�����y��J5]����	� ?�>r�CU��y����F�X�����P�N��yb���
�:��፟���A����y���.&�"D:UFMnZy���ؘ�y��AUdqA��w� c��y�j��fIr�c�<w��*ƤX4�y�ÒF'�	�V��y�>Y&��y� �	�
�! �wJ��j�ybo�0!`V�;O��n�
�2Akʤ�yҢA,=WX�����t�$����y�b�71x1�V��3lG�\!��]��y���Fm��"gK�]ɕ�^��y�苕2^��R�)�.{T�3dCO��yR�ق'V���,)z�h�(�y�V��#&��1\��'����y�P�
my� �/�P��HO3�yҁ�
�������jP��P��yR��D6���s��%��k��yb�O *�ٓ�J�3 ����]��y���4�<�U��N� ��͗�y��Ҡ����'}ʾܻ�
J��y��C��I��dɡg^�kT���y��F( �^����R���Cʚ3�yT�mIr�H��ݤQQ�ȑ�
F��y�A��
�ج	��İ_�x8�R�T��y'Yò�6�^�X��I�S�Y5�y2J� i��sPxā�b��y�5p�#�G�t`�Ly�N��y
� p��c"�Y�漰�C�KE.h��"O�����@�V�p�ǔ�&��p"O��c��*R��C�;�p`@�"O&`���!$�A��e�(}�����"O�(X`Jˁ�Y�eŊ�
�����yR�^�p@��)�⇵mNش!'-�(�y��MfS$�@��Qi�P<c�	P�yb�$\d�,��إ`z�͒"���y"�60�y�'��^kP�`��y�XA2��Sf�͘S�f�����<�y��cu�E���H�a��<s�/�#�yB$�(.��!'�K�V��1OC�y�
].��y��J�S����o���y�M��(�C���O����AV>�y��G*P�8�Ru��Lt��RV��-�yR��%�� 1p!<jJ����O �y��TԲ�F�4�zAQgΑ�y���ow�x.Q�3n��	�D1�y2� T�)�hH�(�J!S���2�yB&��< ��Y���T2���1�y ��t�w�ţH,H!#��y2#�T�+G���t9@H̫�y"�Hvd�ba�+F{���<�y���&U�������<}z�B��y�A�3����gJ	��	�&	��yB��6B���kF:1t�y0@���y�$Zv2��юT��u+@��
�yb/-4�(�T)@��A `Ֆ�y�#8���ب0��`�FP"�y��
-H���� 8"vYCG��<�y� 
*^@0���#�/*�ܠ �
��yb��1N���h�J��
2KP��ybNVj�Z�󁪂Ct����,�yҤNX��v���nTlMp`�^��y2׉�q��f�)m�� �4͟	�y򍚾.�Ց�C�)TpF��7� (�y�@���
�G�[ �m��)��y�Q<���P�\�Ap�c2+���y2�H ��	���.p@
@��,M��y	/N�*ܛ��4����C��yr � _�f@D��>>H`9q)�y��ϊ8���V0,@Zs�ԛyg�B�	�0���eT����0��D;%�B�I8!����'�9M>���(]��B�	�b����Q�T�g_�X
rC�I�
e�'�͢c���MAy�DC��"���hs�Ш*~�5X⯙���B�	�y��r1j�ct���O��B��4��:�)��)�6���C8$��B�ɨH�.�*���nc4�*"�B��hB��:�bXpt�P�{2�)�̟�-��B�gg��:�K�K´ �BȊi8�B�ɀ<��)�W��c��"��3X�B�I�[�$]@T��4K"M
8�C�6<$0(��K�&�ha!2N��AC䉿N�H��L��p����KV�r��B䉫*�Դs�G�t ��甠O[�B��P��Z?E7l�8!c��z @C�I.|:�T���·!e8H�.�8H4�C�1��]�f�P�J�Z�`�l�l>�B䉐!.���Ϛ�d�Fd�P�2��B�	<+�P|�T&��u�@���[`�B䉗t9"�;���Qԧh��C�I$.4�i
�,Z�T̚�����<?xC�)� �}srj��kV h!��%�T��"OޘᵎH�tJݲ���$���"O̘2�H?q�b�)��������"O쬠��	�w��=K0._'W���`�"O<�ӆ�4|@� �-�q��a@"O�{T��1�$ �g�Z�F�k�"O��1GV6!2�yR�0zd�J�"O���E=o�ʜ��%�&�>I��"O�IلkEA��h�Ӥ	E����"Ovp�V˛{���S�L���a�"OH�	�k_S�:%(�%�s��,�b"Or�sv�ɪ�������bg�0�"OFa�w�	�v�@HS�c�� n` K�"O�9�m�>9��b	�7k���"O��S��ǌ]�2@�bџ ��
�"O��p��$H#��˵�ЋY�rj�"O���G��
I��&'ς}3�"Ov�a�f��\�v����+�괠""O�U�v%N*GgD�"��^����"OV����;z����G�׿Q� ��t"O� 3��]&L�IA�o���l��"Oġ�a"L���K�eK9�(ѡ"O��Ѕ��S ��GE:7p+f"O�iWKE�L�꒣�:0@Hh�"O�<¥�S*fR�q�$˪T' �C�"O6���� �(�¢!���0�"OT�:��L��u
�+�\�2���"O��S�@B��nXz@�J#k`�D�t"O��:���*i�s��MX�m`R"Of���
r] d��^�!�N�*�����J�a�zxqa�#[�!���2X*�cB�B�6�ge2:!�D1id�Acf��+���C�B8Q/!�\f���2Wb�&�t�� �h�!�D*E �y3�J ��-ٰ.��W�!�DӞ^*�,ܭju�B7��"�!���/I��M�MA7 �t�C��X�@F!�LMgR����7_ߺ��2.�Z�!� i!���'�|���݈vV!�6N���S���>q�d+�X?!��y��0"*��{p֌���[!��i�Da1΍H�d;�kP�v�!��	/P�E��-� L>��#tj�9�!�LP{2Q���xD2��0U�!�O�he`��3� `�]�����Y���$D�*q�*� %�բ�y҆�G�`jvE^3�����&٩�y�J$V�� ��a'+!t	y�)�&�yrH��-|�bV蒘!�R��EC���yR ��X���� _��P�k��V�y�:p���ڶ����m(,Y	�':�%�'�u�����)Rl����'����	Q�_/�Uj0"�"\t�e��'D�R�@p.�!�d+B?�B��'�\��t�ض~|�)��Fp�Y�'�<�
4fR�TFdhc�*s��D�'n�c�Q-lw�!�ÂS�o�zT��'8�����3�ر�-ˍn� s�'�̈��ŗ��E;�c�jƞ J�'���xD���.$�Qy"bJ�^�$H��'� q2�쉐1�B�0�n��^h~P�')�D���
1w�F��ÅN�HTrȱ�'���P�J��Kd� qH��!�'t�(+�#��?�iأ�B �֠P
��� �a@��C�B�q�GH373n�!"O½��g6pm&|b��ɢ 5���a"O Ly@� p��@�%	3H3�(W"OLH	��߳[dd���bNqS�"Of��F��!�D�Q�0�Dp�"O�%����jyr��`����Z��p"OF(��Ɩ�
�h��Ul�f����"O�8x��M)sxv䐑kK���H{7"O򭲥)
�:�J5��hy��*�"Ot�1��B�S,�4�ӈN�Tl`A�"O���"��	Tt��	�> K��y�d��s�\�RU'��14��xw`I��y�ƞ'�<0"I��'�"40�O���y"�H(��Ё�(;	�����ɴ�yC��ve�%9U��)T+ M	����y�=
����.\��%p�d�"�y�l,�V�JwJM�x�a3NT)�y�Z��1kV�s���"�Ȏ�y�S�<"족$G�=�^�����y���'Ԟ��-�	�.���L��y�M+[�~���H�$�n�Hr/ܩ�y�f�^;���&�<q�Mȵ�y�fS3ވl��	ֲ�H���嚴�yR'�nv�ԬߝwP �P���y�-�(d���׉@��m�'B_�yb�# {�v�p�0��&�^�y�G��<zV��V˕�c@�H�#
��y�� �`YU�WNI0s�E��y�E�2��RqL�K�T@�B�Ӏ�yr*��D�b���n�Q��k� 
�y��Z�Ip��e�Ϝ�l�%��y��,5�ύf�l����0�y�af��lR") �4Kp��A��yR��|9F�Z�&C��8%�])�yb�? �Tb"��St��(�y2��#�JH�7�:�D�2���y�R�>"*L��ϗ;�~�(�b*�ymΗ
�D��A@�4(&H`b�)�y��E�hꖃ�$+��h;sJ�1�y����j��ä�%*t��3b��yR`��BL�#	*�0��a�9�yr/_+B���&`&��� ���y⢝�&��8��CF��"�{`���yb�T������8y��g���yb�#I���"E�9vLp0���y�i�h+�D��KwPX�79�y≔�+sz��w(��r�8��$�^�y�,^^�4�Tj�[��E���_�y҂�XV���� )��^'�y��K�Zl��&"����5��-�y�\�*��Bf�θ0~4eRFU��y��E����"��!��yQ�yC����:�e�-(<��A �>�y��-[0xS��I�{�jҘ�ybK�[�D��ȀH����2E�y��@%�RA��X=WUN-�s�Q.�yR!�
����g��<�ɹ�%]��y�iL�w.��a�ʥ \r��1!E��y��Sz�4d�#'�DlQq!��y�fÍ$�h:�$�B}y	a�܈�y�U)$M����(J$�\���)ɥ�y2Y6�����3i@�P����y¨�FA<|
�I��A�&���1�yR���A�A�ԇIN0�`���y
� ,P����r�h�{ub�<"���$"O�T�o�{m��t����\y�"O��g�R������[m�	�p"O�����C�v�ih._�I� A;"OVjr��A��E��*Ś=w��k�"O"��cFN ����@I�k`:A�"O|ˁ�?7!8� h�P��!�"O�E���c��F/�=[0))�I5�y"lK}4c��1BP��gE��yΨT=����3YN���y��D���$ĸ%�"�+��ӿ�y2O�'0B��·GO6�� ����yr!S�7K��ET�X�nE"�yb��z� � �n�T�N,�y2]$~� q���3)l�a�k��yҀ��Ex�����Y��h[�!ě�y�鑡Y�@�x4瀺R�,y*����y"Z�#/G1G�z����y��7�(��U��bH(�$�2D����G@�o�Sǉ���:j�-2D��E(���}���0Ca��H�O1D�|*��Q�p�`�CU�!V���Y�,D��(rkU�n3T!��hК
v�e��o6D�0���-��([$f�o`���j0D��벬�
vz�D+�� ;#�Q�c$D�\���$S��=���k���x�=D� "�NN����x�L�<��xCGa&D�x�D�:1B����aT$
!j"D��恝�m��e�����"�B��$D�H1�S޾������?�^d!a�"D��!	w^�i1bZ>��Z��=D��� �M�l4�͖�+��d��1D���@S,�8�HS�G�� �z��+D��*Y<E��)�J�wo���a *D�P�����&�jM��lD�+�I�f�4D��Bm˥]���d�G+F�f ��	'D� Yu��]+RI��Y�c��$��O(D����l�T@�"��&M���S+&D��(�ɂ0J[@-c��	;"�v���7D��y!o/?Ԏг�������)5D���/Ͳ�z�𲅟�i�𼂶?D��!dS�G�(e	����X��Qn=D�z4�	>@���ڧ ����:D�$h��X;v���˵�J��L�s��7D���u铓=�p�ó,�'/.Y��4D�D�#�\	�]���.C2DA'B4D�:3Gֳhox�P���]�pA�h2D��;0��-,x@,Z1f��=0�ec1D��DZ�m2��/��e]�ـ�`1D�t9��*P0e;�c�ZO]cs�.D�P��CG|>�5��\�\I,D�(�3����sd��C��\zA7D�p�3��#+d~���؇&6D�:�+D��A�z�`�*U�^MVp�Vn+D�ȹC؈&�� ��'!E �(D��)3"V��:]�0��}gT�
:D��z��	=I$���4�����2D�P��C��L !U)ټ���ɕJ;D��ҕc�7i�^�R�Č	�0T+s�8D����=2m D��\�"n�'�!D�`�PL�T� W)�/9�)���2D�dr�S#5gN��Z�I�ر�3J=D��9D��;���� J�/�1	�L6D�d��
P�$�Uñ���bD�IR,!D�� �!s�_8�����x&1+�"O���ᄚ�VVNSPć�G>�"�"O��8�S$Cn���� )%Hm�"O��a�fP�w��a�/~���1B"O��I0�ȟ@� ��I�7F�h1#�"O�	�3��-�"D�WhE��"	�"O�u��^�5�d4Q�Gԯ_����T"O~hr&Ǜ��L����*J|@�S�"OHS&!OrX�0�͞ka͸�"Oz�YÅ"��S�.#�4��"O��7f�!��Y V��tʕ��"Ox	%�����+2 �7Q��4��"O��9$��&$n��P���!a�D �"OF9�E��?[�B\��@X������"O�1F�L��QS�:��=��"OH�5�Ǣ\~�K��;$�1�"OP��3G�\��	`��0��5��"O��:Tj&uc��Zd��
!p�%	f"O$5����Kj�]�EF¬S"a�"O4�@��M�exbE0a�Ĩ>�ڒ"O��R$!P��p+�,�(	lQ��"O���mI�,	7�H�i�"OB #V��q���ݒ�l�"O��veԝ1~�0,�\�U"O���,�=��,D���Y֪82!򴴱z%jX�3�� ���H#P��Tc	�'�6���NT��s5��	j���'t(�*���6@XU���K� ��`1�'��0'$�����Ä�Z� 5���'&�����o�\91%m��$"�0�'��P�F+�3d�v��t�>! x���'�4d3v�؇M�Xzt嗵<��'F���t�S��%���ͳJ��y�'�Ji��N����j�@(�^���U�f���K�2hl��d!��@{z8�ȓ��h�^T����E_�fZ��ȓ4��1��U66@��G�%3�����Sb�@8XK��@a�7��ȓ9�DqӉW�}�j�2����D�p܇ȓ1j(�B߀&����dͿ���h^�Ct��|�P����4�u�ȓ�l��@���)L�(��G�-���ȓ��X����q����u+1Q�ȓk���	�6h섉�D��R$(�� ,H�QD(X����U�W���ȓ)M�@:���!#Y|]2A���|r6��ȓd_ʥ�=^f�œ���
�.D����K� �T�ٽ^��|(r� D���lO�}h�=� #֖JL�X�s#?D� "G���9kƸ��&�+C+����:D�T�o��`�-�r�a���W �y��ѱ�B�E~�Ӏc߫�y��8��ܢ��!�h���#�y� �6B0����4�-y�M��y��",�D�$�9<B4	�����y�hx��4b� ˽~Ɣ}�p���y�,7а%�R��*G���'��y�	؞oC�Y9@nO�@��S@�L��y�C�������̺&[��H�*I�y	[��4p
'�ۧ(<�!��DV��y"�,_�p���2�ٷ垢�y�K�0�n�ڲ֗	܈�� U��y"Fř2��R�f�}K~��A�y�HԢ~���ei�xѴؠe���y
� �L&OV�~k��z��+l��� g"Ol�J��]�h�sr�[�PP�"Oz|q�+"���E��S���z�"O��Vf�:L��y"Ӄڕ	V�i �"O����n�� c�}�U#��]LDL�"O\d��"]B�%A��04�Q�"OTm��6\]����!��@�"O�1q�nM�b7��'oׄJ�h�"OX8r�ںsq��PA�6�@�Q"O0}��f��:m�=�����v�3�"O6D��Ŕ8Tz��R��*3R��&"O�㦉�UP<�!l��<p,z4"O�H�����6�P�*Cʚ�j"O�eb�D�Z<���&H8!�����"O|�E�2-���@i�P��%�"O" SD���c�1Ӈ��T��5�"Ox8���^:��sp&G�J�N�"O���E�	*������8����4"Oz�K���lp���G@A)j���"O\ak6�X����AC>x)��"OJ����@���T� %ˣ"OȬ���[����),߶}q�"Olɩ��.Iĥj1��d�"Ik�"O�4�a�?ԙs���Q�j�02"O�5R6iHU4԰j#i� �ԅ�"O"iX���
���8 i߯l�(B�"O�|�&K�V���fG�
���"ORL(��#��-��FO|��!"O�qp�Z?���A���>{�E	�"O��F#c���y��E�Fφ�yu"O$�0�"	HS�rѢ�W�� �"O����/�S�P��֎}�Pau"O�T�"k�$j\
@�ڙ8"Ol�ەL�RJpm��nY�.�[�"O�`H�� "�X�re�D�c$Ե2"O��at��A�ȵj�MN�J��"O�4Ʉ΂�x)�9��e�S����"O(��t��vg2�P��ΓJT��"O��@���'k
���c��XO��"O��s��˥,0P5�"G֐�D)�"O�ax&���	��)k�:I�i2"O�\�� >b��au/�1CZ��"OL4k"$�P�T�sI�>V:P��"OՊU�H"Y帤jB��*w�2��B"O
�X�B5��� 	G%W�h#�"O���Am��'��d��@l�ޡ�f"O� )s�:�֡�dŮS��h2�"O�1��H D�$���bX��NȒ"O@)j%�$*HD �c�(F���"OpMp媉�G�"��a��Il�M�"O ��w��zV>���!H6Y��""O^Q��<�t$"%G�O�
��$"O̠rgRo��<�0˄�@'α��"O�)` 垇,9��C�-u8�كc"O�Xv#޼PȞ��WGX$9a�"O����cg�1QbQ�U�I��"O>fj�I:v��,kp�
'd���!�'5̱
�'�@*�"�9\g!�D�>��|���0fe*L!�lڹnf!�d\3vs�!L>}�Fys6k�;NU!�ڛ�"`� �'�*h�穇yj!�$ēF(�j�@Uw���{''ؿlB!���0ta�++x�Ц�!g2!��A6�����I7ll�Pf��ZB!�� 0��MR�q/�%{� CkԱ�U"O -{gl���u�$dOX����"Op�щ�op,8Ţ��<ٜY�"O^)
C��t�j���ŀr(��0r"O�P��".`+�a�$-�L�"O4���3a�Tp ˭em��ȧ"O�QR�ɸx#�Љ���"jlt�i$"O���[��`�ՉR�
M:�A�"O���h�V�0x	E��+SKA��"O����ܔf���Ӈ��U8\ ��"O#��҂Fa�����2oL4��"O�,I��N�;~�er���<:E���"O��9�E�7	.�Jwo�H%&�y�"O"�p�	?$P\:��2L��"OV�ඡ��9p���&�@�yf@i�"O��+`��	� d��%K�+��H��"O���ҋ�4I�k֤\0V�V��"O���
3]�ȸ�խ�';L�I(�"O��aa�QF��``$n_�E*ej3"Oʽr�m�?,4���%�*�be"O 4�MՍF�K"gZ9}�X�6"O����O�:���Gݒq�1��"O���v+���  b.)d"On9�cLȻM�\�{!j�-w�FU��"OZ��e �
b^i�	�9���yC"O�1��фz�j *��au6%{�"OxŲ򁃢gE9�"$Qh6!2�"OdP�E �n'N\���9CGr4r�"O:d@��*Ew���!���
c����y�@<&�@���V'2�y��'�y�d�)'��2�%?{ԥ8�D�5�y�#d�@Y����kqD	�y��M.P)f-"$h�.8� !�)�y"O_�+X�`�B�-�����ی�yR�+.:�� �c��-8�̨�O��y"
��)*��p��6-�fP(�����yȋ�hY��r�Ǩ28P��J�y��E�D{�#BN�;�~�x���yr�ѲRZ��f�*%(�&B���y�E�:� ɺ�H߆_f�Hb��yRF�?�8�Kh\�lM�9ss�E��y�C\�"b���=^Q�pKD+���yb$@�s�4�����H� 
�.��y�.�����x� UZ��y�E�J�Nu�$�:���
��&�yrϏ�C�pP�V��BL�A�-�y"Α�l��ma�@�8gؑխA�yB'�m3 �@B
R0a�DJQ��y��.����'#F�(4���y2J�K[f��ӧݯ I���)���y��E1���4�\�������yR�vS,	��ѭ<x���I�y��oh^hytH��$��ip#��yª�0&���b�s�����<�yR`Q>K��Hd�ގ���
�&���y��]j�<Ati�?�$h�q�R��y2�^*���KF��w�1� ��:�y"o�>7l��q"	C.�|!@W�9�yr��" �p&�\��&+��yr��-;�`G��`�Va���yB+ևd� � cC�'�
��plC��yb�i�@<6��@�$���ó�y���a�T�����6�\���ǉ��y���Y>蠷'ϴ�^��2#D��y
� �����	T�ʙؓ�K�0�Q�G"O�t��А ��mڄS�*�R-�d"O���������� �E6"�0s"O���|xH�1d�H
2x��"O��*w�M�5�f�Zs�1+d>d�T"O`ᡱ�4�};��Zx� V"OFǒF죥�\i�n��c"O�8�E��P��d!Ǚ+��,�!�#�, ����]����2�!��Wʖl��Nj��9�fÔ�_�!�$?y+,QX��߱,a�0�&#C�3�!�ێF��pC�*�Kꘐ�⋖E�!�D9)�bu�g��R8��ȗi!�D�F����> 7��E�_$P!��'^�\�q�<����A��--!�D�3�^%q�l�XK�`P��:	!�d" �$Ez0�̉.9�$��N�m�!�D�>���\06��C4oB��!�䙎7Z� sG��hX\�7L"7!���m��5H`���F�
�HM8!��Ҏ-d�5&.C�����CW!�DH�@��+T=o=SĄ_ !�LFyb�����u\�m�3"!�d5.��/LxM�L<�`� u"O�@+G�-~h�tK�8+,x�S�"O�A:H�c���k��82�q��"O���V�(���V��'^d�m�f"OV�&߀�n!�EFŎkP�;"O�qӢ�28���2�Ė=O��m8�"O�|����=W6���E�"�  �"O��H	%�(��	
2��|r�"OڈCEAG�%�Q���p���9f"OD9�Ca������+�:�"�"O�eT�6��y�r"��+�@@'"OuJ �G7$��#��Tm><�"O��f��"���� Mw1�s�"O��ɗĄ�m���+!�O�-�(��"O��k�D�}A��ru��v\� ""O:hA��ި. 1i�&8�n��"O���E����ff:}�j�Z�"O�dP�`� {,�%Ѷ�l��"OFj2]&�Rp����+���c�"O��yB�Hy���Af`ҢS��-�b"O��F.@�	x�	���E<#���""O��(VH�Ĭ��#
!�xhH�"O0@�`��]�BZ6)H^$2!x�"O%X�[a6F<���e�\�6"OB@2&�]�C�vс���T�.pH�"O졋�H5��=�2��Y$��J�"O*�h�)ſ:��y�`�.}%�p"O��@n���M����!���)S"O\b0�Y���9�/;���q�"O�\��o¿��h���A
�@d��"O�Y��F�+r�X"��U�قp"Oܐj�F~��� O�l(LS�"Oʙ��ӎv	NA@�۸�2ԩ�"O�Mң�M.��Y����,���I"O�!#��9Z�=�G.O&Mu�<z�"O�\Qu��:j� C,<���T"OP�`�$ܪpJeh`���"���r"O�9pV6�h�u��	�r"O�q�`�݇JF�iѧ�#�>�;"O���"�W	;Jx����<w�xU��"O0 C��T�k�cϙ=��uIS"O� ��C7}��sǮܫ*�A��"OpD�EL��_�"�r �E��Ӥ"O����Q~����sH �i�:�"O��b�N
Pέ���7�(\�"Oԭ��pg&ā���?KD$#"ON��NAB��"F�1�. �c"Oڼ�Ӳ@�8A; �ˑ��P"O���0㏛>��ʇ�0P��P�w"O��1C�֙5	HAaeW�u �'"OB���VLHCᢔ^�����"O^1(�.��DQ�p+�#R"i�"O�p$ɐ�*��H�oV�ec<�Y�"OR�)J?J ���D�0i`x4�#"OB)��k#L�^y�6�!Dz��V"O~�@�dΥDn��3�Nڇ`5�pC"O*�b�.�ā���k����"O�p1�G MH�
3�`���"O��DA�9o�2̻��&�t�A"Or;5���NS���I@�j�(#"OtLC�D<?%Fe���\���E"O]ʶ�ץY'�kwI��V!"OX� �j:�*;��5X�vѱ"O6�I��;�ީGX�GE�x�4"O��c/��d����:SD��3"OȴZ6%�3<\�A�$��&�=)"O����"K)��;�b����"OPp����Yl���Q��+[�ȡzv"O�@�@
�q���l�y}6���"OąX�՚*��Fk��o�lj�"O��˶���u۶�C�i�1Oft�8""Oj́�bRK�t bi�:d��[q"O%X'xӦ���#]|I�B"O�HR�7#��aT
G�`���R"On�Ӧ��	 ����O�\��U`�"O^T1��yר�ёH	� ��P3�"O�K�����x��S�ul)C"O��U3U�^����	R��"O�ݪ��F�z+,�C�O��t����"O���7��,�u�n�t
i�"Oĩ`�g�>$r.m�č�XVVX��"O�=���۱�P�('�6nبd"O&��uMZ�ȓ���n�b�"OU�F�B<�^��!@��s"l%2 "O� 9!��r�*E�>"�-�S"Of�ЊX@�'l\�-��)��"O�I�t� m�~\�2j��:͸�"O0a�u�"O�y��O�jI"@1�"O�l���pY�@r�OH/B��� "OVH.t��z��
��9 ԨW0W:!��E�}q�� �&� ����hR�C$!���Q@��Q�n@�T��e��	�~$!�>6P}� ,�}�А�ޮk!�D 7.�"�	��*�h *��:+!�䜨P���%BTP���w�]?!�d8(!��Zi崕!Q p	!�F�&V�`��o3D\0���I�!򤏌@T���)P�Eٷ��%s�!�W$ ���ZB<;7��+�!���!�i@el��p�Ś�+�<�!�
V����]�*RZQI�k�$9!�ď��֕&aQ�Y^U�5ˀ�K�!� �V�b&�И-s@r��L!�B�j�֝���O���a��,"�!�D�8�,M2 o��8��!���2f�!�� �A���2N�L#�@&`��)P"O8L�#V8>���a�H�(Aƌ0�"O~�A��Ɩ�hp 3�E�LD��"O�i����}���Է/�0��"O�1c#6��\�ӄΟ
��0�V"O�ԠcD�2d���a�<���"O&l9���|ٸ�!ў)���#"O���d�a��6���}Ծ� �"Ol���ϟ+���*Ԣَl��aؠ"O� �G�(�9��˜FŬH�$"O��� vE�,� i<��F"O�3π19������@�f��T"O�)z�N�%քX��Ϝ	$����a"O"]�s����D��nї0��$��"O���� X+F�
���D�jSl�"Ol`�.�
2�i�R���
=rU"O�p�t�8��%Ps抮}	*�"O<X����g�64; �ZG�,�"OF�2�������ץ��*���r�"O`�Z�KN�gHJ4���3}���R"O�Ề�#������/0�V"OȅZfF��C�
}�� �!9�2"Oh8��ʑ�S[0:E�� bDx-��"O*��v(A�;���0O?2+�xc�"O�ě��K	���R���UB2u��"O�X;V�Q7��5�`e��zTx"T"O!���L�5`#��
V��"O��:'��d�L):$G�;i9z%s"O��H�I4� Є4��Kw"O8|0�ɔ�}�Na)�X;h$H(Ñ"O�J7
X�d�S�A� Xh�"O��k�#�:B$��jˣb6�(�"OƑ�� [�\H�E	����͒�"O�\s�j\/V��|����O����"O\�j�
	5p�ˇ���w�0��"O��!#�w��ћ1�4O���a"O.�Fa��E4��3�^�k^Z�@�"O�	�e�'���b�,rm^}��"O��*�F/"!t��#Of�{�"O�]��mF�`d҄���N1�ĳR"OP�FlF�(j��4��]�(�&"O��:s�DK��!�?.���u"O�qRǐ#b�j�`S~߼�Z�"O�t�#� p�x�Q��#�4���"O�9��]p0��p�I9�Iy�"O��vCA%u��mab�ȡ:� �E"OX�LJGaHP󢢚�6��=r"O�5:���C�}�% ��:���(%"O�ق���nR� �q/ߔR!�$W+���"���4K�5a��L�!�d���i�a��/3]���LQ�!�d�6z���
�-@�9��`E���!�DP�`�,X�C˨8��I��	ڧU�!��	X��b��; ���GS�U!�D@�a`|x��A�?q��v !�H
oy��z6$�*~�����"=t!򄂒x�z��D8O����*]?O�!�V��DQ�vd݋Q�~�q��N�Gw!�Y�#�T)�����cx���1��,Df!�D
7m��ɶ�ü�~��%J�#O!��v.u�$���eC���0D-!�N
i��yc�
�9��}0� �G	!��
?����G�&]�Y�i֥]�!�� |���nюg����r�W�&!�� ^�т�
U�$��&* �pr���"OJ<@�M*@̐�Z`
	8�I�"Od|БOM� �����0���	D"O�DzgER�@���CC�TqB�a"O���#�Ha�-Z@E�!5�<�"Ol�� �� 0���#���F( ,*s"O� ��8�bh�AmA�8�-!A"O0}�R��Є��+��1Qɘr"O������Ti�
�"=�i16"OR���B˘\�A���H�N3p"O�Y�#� G2�8���`3"O�͚ ��~T����L*J̨��"O"�qDn� Y�,����Q�@9�"O�[Pm�yJ9B!� f�:��"OXFk] $��r`RY[��)�"O�Z$�ۈE.�3���#H.�[A"OH��f�	��hg�Ɠm�t�E"Oh�3��T9�H�2B���z�،x#"Oh��2 S�Y�H	o�G��P	�"O:��cE�>A�x���T��d��"O.d����h���*	
�t<8�"O6�Qe_-y������A/9�h�x4"O�p�W �2��!�2� �D�͛"OT�:a���i/yN6B��\h�"O�q`/��w(��cNZ����"�"O����C1I<��F�����"OB��vCJ+kC:�qE�BC�2ٺ�"O��ҎMz�";���j�"O���7��'X�L�0(����a"O|I�¬װ:��dc(K� ɺك�"O"=�G� ���'�챙'"O`�h����);��S��Q�|�k�"O��K�GQ�WH��pm�<R�"OX�Ǎ�k\!��<@��"OEc�GH=~}��:�	ͪUG|�Q�"OX�V��#|��8��b��i1�5b�"Oੋ##V�I���֛=���"O�8���;�|���hN5r	>a� "O���w�N:�~��5���/��XF"O"�1+�
[Q0��gȔF�=��"O����(	�i"�9�&���"O�-�`ɀ8;x��P�ΰT�&�@"Od����A�4�AD�.(zPa"O���ա�*BD�Ł6�T�D}�x)�O<u����l���COGX��]rB��_�<9 *ud��ө	q9zPo\�<�`A¬`G��;�\�2d=h�X��x�'Q8L#�C�-���:Q���+�p5�>y���)�e}1#��N�<�17S�4�!���-��Ppb^S���`��!�Q�6��!�M�j�F0a�@�v�!�d�%$����
���l�`OΞM�!�$5^nXa�*��?�X���m4_!��I1'�]�fe�"�*�ۤ��J5!�O�d�2�Х��!� ��5x0���OZ��g���~���Fl�&ZxK& �|�<Q����
�cF�}�l�*"�<لO�g�XM���_l��i��Ϙe�<ADg�*b)[V3O@Хz¢�dyB�)ʧ}��@���E����#+�JxEy��'ŋ��U�!Z��d�ګ;��R�'��ᑔZ5(�`d�)hj`���y�!�W`\E�"L7<4�1�łV�ye �*��Y��U!3�|�.�=�y
�  yP���-)��@�TdW{ i��=�S��y��L�:�1g�6$��g�V��y"�)|��r�
	s���� μ�0=Q� �i��c-ׯlx�P&�2�ybbT?N�ri;��M�`�.������'�"=%>���κh���(iV�R���>D�i��ވ=�h� nИ^��	3s�&���<I�͇�PN���2�htS�
XF�'�qO�!��&�/ѽ&q��daҾT:��-h3�F�!?9	ߓ&�<��K�#2*`��P�UX��'L����Ϗ$��q�Bk��W���""��]M�|"���0�I3"�b�Ç6o��YV�׏c�B�	<������U>$80K�0GV��?	R�=�''T 2Έ ^��s�)�N<�'b��'��h&�G""Z	r'L�3$x�,O�=E�d�.Ie��Q�a��m3�yz�&���y�]�p	�7-��d�����+�yR�܎��M��F�ox�M�����y���l!Py��0g��Es����'���Gy��TOʽTP�DCaN�a5�ǉ��y"I�2w{x	ET�1�θ����(OZ8��:�MY,q�]�#
˱%\�qY�#�>�J>��y��E�T��Ak��WN�(� F"A)�Op��d�cW~�`�#� ����<.�!�RxR ��Î�/פy邉�$.�!�N�v;ؕ�$7m�@�v�Fh�qO����
t� eꐶ=T�-k`盧���1@�T�7"ԇ���y�	B3[c�8��		^��� .S�
��/��i "O�
��Z��(j�i�����r"O�X�� ȝ:n�hҷxo�ёv"O��[�h��I��Ƃ'io�-)"O��3���K�.���K�{��If��؄�	91pl�BC�"Q@2w�͢G����D5�i�D���� ��O���d�'D�,jqަ=&�t�2W�H�t�s M*D�4�@�-����uI88@(-c 6D�$��6n�y3r�5[̲L��O��=E�T�d�h�˵��c�p|`��9C�va��'�'�.e#F��D��#-F��e(1��j�`#<q�I�>Ϭ!u��0GB%��}�<	!��x̸pCI&q��@�J���������>��e 0PŒ\�ǤR1b.�2�%�*��'�xR���W��y�V/{���$CA�U��xXB��M;�$�O���W�+���&(�2:Dh���"O�w럿\,����)0Cv��'9�N,���w�R�1�N%p���t=��i�ў"}�qX�~��X񁟯Ra�|�`OCF�<���']��Iq�Y�aDH���~�<��"��ZL�#t�U,&��h�%KF�'оDyʟ.�p�Sp���⪎�؁�*O9������z��tL�MJ` I�'�0	���35l�YJ���y,�y��'yt<��$�1���{����=6��C�'X0y�`i��(h�s냏9�K
�'�Pa��ֶC�0d�bi�C6���'�^8i��
�<�YkF�d�����<��I��SV:i��W�Te���T�D9}��O���'��0�a@�@JTY$ ��'n��'��iZ���%�l!H���9�'�0QC��R;%�M##�,p�]x�4�?A���'��|ZcjB��	LV9�d��p�ziz�'2�����iա#�A6XА!��On�j���Z?��K��=�X��e��{~BG�/¸π N�Z��/ښcdE�@e�i��H���$��YY��!� �}ٗ�Q�}!�D����PaɆ�"V��+��R�~!�A���\5D�?/P���
��]�����<qF��6K�ـAdJ ��UC�<���%�xA��%��.}J��K�i�<��G¯N��ș&��81���Nh̓��'����}�զL�z󸝢c+K��0`�A���A�A�)��={���6�tL)�A�r*\�S�/D� ���qzmQTn0� �;D���\"��I�7 ["" �1!�:D��k���&_|Ѩ�S�3Ȳi�6`9D� `����o����	�PYc�+D�P���ߥ����ggZ�}�T�:u.ʓ�hO�jEx�Ġ�On�P�N�J��B�	!P+�@�4a�h yI�T)F� C��$]z�	�a��0���� �:�B�	�H�09�Ϟ��|�+сP�t6�:LO�b�HQ�oC�4^i@�i���g�$T�4��_���J񊒶|2:����$V��(O�OL���]�YD0�s�'I����'��$��"�]RpI_�DL*���'�����kCfU[T`��=�=��'���@��tZ�@zt��4
���P�'h�����	r��= ac���T!�';ܼ�5�Y�n�[�d^��'(�Qjр�b���/�(�#�'^��Z�֪>�9�fn�����	�'T�jFdǥQ\
P��ɛ��ع8	�'}�5�9��m���(@3"O\)�׈Ȧ[��Њ� �If(�"Ob�"J%29��S��7O�m�"O��ّB�-qХ��dA�5��e"O�AI�X ��'�E�30�E�'"O�$2qǞ%,BL��@L7����"O���/�1u���Bd�D�{nXc"O|�3��ܬ:e\�Y �L�n�~p�"O����M�,+��ʀ��`=(�"O>�@B�lN����H%\"�Y�0"O����\w7ִڢ��-h����"O8��� Y6���a��Eq�"O�Th���Ol5�tF�*L��x"OR a�k�,Z�$��C/B�����'���O�_� B���&ec�'&�H�B�J�QHN١4�&����
�'T|�d�5�vy�/˨h�P�
�'����Č�qT�ř��Y�\��'��� �c�3E��h�u�]�M��x��'�\i�7��r�t��Ej��y2��'yZA����4k��$�����?²���'��i���~n�����Ӹ6�P�8
�'��}��-�=k����Co��5&� �	�'�y[��ݑof�!�D���<�T�9	�'sjL[a��&�J�j�lǞ~<0%K�'�Fl��( [�
X���"6�a�	�'���10B��)�� ��̇��80�'XƩ´�ш�pT��G�f�"<��'�>a��O�Qkd,��Ζ\��\+�'[� �S�F+�da�W�_�A�	�'�E �z=BDq�J�c�"�	�'Frl���ûb�\� K�\�����'Q�}t�ۊ@�^�((ZuT��'>�X5D޳^�T��cʕ�VV����'O-��[�}B��Y&g_RLU���� ]R���'����I>4�V��"O2yTĔ���C�%z��2"O>�GM��5�Z���"dq���7"O���%j�n���A�ƶ3Eİ�0"O���!�J�o�r
�E2X���"O�I�V�Gx���G�	Rܡ`F"O���eO��p;����.VʐHB"O>X��&JL�0�K�U
��"O�#uL�ш1I ��1n�!�"O�T1�*�������mk�	�"Ohtz�E�H, �,\5SU�86"O`ĳ��A�=Ð9�s�K�yLRu"OJ�wSuc8�C@��=���b"O�G��IϚ�*2�*6"O^ �BM��3�Pρ�4̋@"Ole0�h�0
�[�3�\���"OJd{�dH	�x��>2�ڵ*w"Op�K�#[�X���	�Ei���@"Onp�D��7�(�ˡ�M�G�xs"O��;B͝0B3䐹�f�0Z8��f"ONP��!{�P�;'%ʵiF��F"O�J��[!U���cQe�\�U;�"O���4/�,a��J#�{9�9 "OD�!Nѳ�4��)��^���#�"OZ� Q��_M��S����n��T�"OF�h�k��= �s`f��p�P�Rc"On|J��+e�|AY�$Ρ}hъ�"O؄�S!�8Zq܄�A�ُ5�P8�*O&|� ���, B��v�T���'� �#��)���hÒn�����'�ր��mA=_�|�� ��f�hp��'�v�Zvi�4m8pUM˷P�|x��'L�x�A�6vh �A�G������'���&�5t���3Y!��FQN�<Q5��?�
��+܀_(Zl[�B>T����.-g���΄��}��1D�D	pb����/*LƸ0�
C0���T�*f�0�� �x�����4��L� �j5a`˷�x�dS�lftɀ�3�ά2ǆݶ��'�ܸ�f�	&-#���aۋ	d��%>GE��0;���y]��;.,D����&-X�Yz�B3A��t��C�`y��E]�e?* �A��L�x"}��'�l�%N���C�aTbFM
�'����t�J�hي��T��#G7�-�Q*�be�5o��|�2+Q"ߚ�%�]d�'�����37�Pa�6fB�*�<��Uۤ��e��?�j�S�̋�:,9Z�,�"`z��H�lA*��h!#��ƒO�xcR"�?	����E���7���u�H�<h�F���d|�@Z��Җ��'}�P�OR���[�U�Ph�q ؞5�4�O􈥰�B�D�,��Έ�{.�1B��
*(�X�A*�$��"�"�����N�ĸϿ3�0w���8Y��`P�]	5j�-�������EhJ�1+Ё����E��y'�/v��}y5
�d�
�@�P}�F�BG�^WS�(r�-� ' 1��O��qYe�J"f��'�8ܫ��P۶��L��t
Q�	ý89ia�ڲZ��e#� ч�>ȓ3P��:��[��00���^�Qtn]1�/T*���*7BھdA��;'��N��M�q&��[�x"bTY�Xh�G�ɶy�����Gͨ�BH@� �[E����'�"rμzY�.�A�O��iШ��7�N�]�7�H�դK	|r�L�jj��1���f�ِ�	p�D�h��6�dY� �n�z���u>0�DB��7�%	0��|2'��������.R=ZE�ŘפA;q�4�A�۹Z�,����ݎ|G
�{��������|b�>��T13)G�=˘����L8����6�j��#�:mC�� C�:+���?Ii7y�]a�c��,�)aB�+yo$��U�ؖ3�c��"~��W�[��]@�N���ǅ�����'�:��th��/� ��&��$z���@�+L����MC	h*6i��`��>��$���HK�S�xrQF�B�^t2��=�J��zU`����G�\�S��-R���Ѕ��Ăd�ꀄ���>(�'�� (&u�P6h��}BRM 4��R`�����v}o@��PA@����a�'N�l�����������+�hP0��C�o6�(��l-~���1%�h�A��e�f��@��T3&s�!7b�S6x7(R�D� .C*][#"��d�q���S�s@�!��Dҷ0)h,��F��~:2-
wD�,@.�'3��Ӵ6K�E���`d�%z碑<4*m+���oTD(���t.�[�S>qpaA��}�ڭXTO�<�2@P�[��)����X�LL �O���.�\��1�&iazEjq�=d��n�Y���^itQrQ1O�84�;�έ�����
��s �3�`���ä�
��> �7m_�>����q#B�gA?o�颃�;��Sl��>�f.�h^y�(؁��Zf��7�l%�eUs�/݂��Zf��2�d,�i^y�'Պ��\cY�L��4�X����1Yj�X~�M��7�Y����7Xi�Us�A��1�Q����>Pb�Pw�A��  ��]gj�Yd��,���#"��]do�Qn��'���)(��[bl�^c��.���''v��Ѭl�ƯK ��<�?��1=r��ӭl�ĭM��;�9��64z��ۦ`�ˬM��>�>��1<p���f d��?j��t�1��I�4�ih��4a��|�5��I�0�`g��9m��|�:��G�;�eg�K��A�=�2���:�w;d�L ��I�5�=���;�t?a�I��@�9�7���>�t?a�K�ո����#t$��NoI;��ź����+{-��LlK6��Ƿ����-|*��EdC?��̳����V�b:
qF��h��xY��U�g=xL��`��zX��U�b;
qF��j��tU��]�.pwq		>����3�"O�Q�,puu0����6�*E�[�%x~|7����6�-B�R�/}zZ��4O���{O�P���^�	�4O��
�|G�Z���R��8E���vB�X���[�����Jن�g���
SB}�
���GҌ�o���TD}����@׈�m���UF~����j�}�P�;|�#,�G���b�w�]�6w�+$��N���b�x��W�1q�.#�I���`�t�~�����~�zxo~!�Vy�����z �{xo~!�Vy�����~�zxo~!�Vy����n�����x(Hj*��ᡝ�`�����}-Oj,� �孒�m�����q Ba'
�
�<�B+h|/P�n��lE�4�<�B+h|.R�m��nD�4�<�B+h|/P�i���gN�?�6�J,q�3V�Pl��ˉ߁�wb��pu�2P�Vm����ҏ�yn��yy�9]�[f��͌ڇ�~i��y{�8]'g'�X����I��ZP'g'�X����K��^꧐X.m-�P����C��R覑U#b �����T.�8h'S����(`�����^#�5d(^����!h���^#�5d(^����!h�����~W'"T��"�r9(9dT��y_	/*\��$�z1 0n_�	yQ!%\��*�y4%5mZ��
uw�[Ҿ�C25
�=?V��{�Qڸ�@35
�=?V��{�Qڸ�@35
�=?V��{�Q�b疕�e� d	��:�"�Е5�h쟛�i�!f
��;�!�ܘ6�i잝�k�+n��;�%�Ւ=�b�Ĩ� 99`�)쒽�v�+W-D�Ĩ� 99`�)쒽�v�+W-D�Ĩ� 99`�)쓿�u�.R(A����#=�N��&��PmH^���?�O��'��VjCW���y:�F��-��ZeN[���z8�F���N~��	�E�T���ss�j��N~��	�E�T���rr�i��Jz��
�@�^���~~�`��K}مp���/�MU�?Y݃w���'�E]
	�4Sچt���'�E]
	�4SچtL2�U��ܫs^����<�`^M0�V��ߩq]����0�oSA8�R��ީq]����;�fYE9������)�1\�A�L$|0����妭�(�1\�A�L$|0����妭�(�1\�A�L$|0�����U2�v���P���V۷i2-�X?�{���V���Uڱj?"�P7�q���[���Pڳn:'�U2�E��P�M�+S֦vX1��-E��P�M�+S֦vX1��-E��P�M�+RפtZ0��-E�
�)c�_���yx���b���H�.g�U���vr���b���L�,e�V���rt���j���H�,e�VJ`�&h���T�6#���bJ`�&h���T�6"���aHa�&i���Q�1+���hMe�$|��c�ʰ
()߂�Y�Vy��b�ɰ
-.ۇ�_�S}��b�Ȳ,,م�^�S}���.�ɦ�h����`�H�y�\�+�ʤ�i����g�O�u�S�$�Ϣ�j����`�I�}�[�*�Y=��)t���#bdÛ�C\_:�*v���  ag���@_\8�*v���  ag���@_\9��ئ���⥬����z��O�ԭ���㥬����p��I�ޠ���奭����r��M�ۤ�]��k̠�1&e��V�̲�X�nȣ�1&e��V�̲�X�nʠ�6.m��Q�ȱ�_��Pd��l}�QN^��:�3b�\h��hx �_CU��:�4f�_k��o}�XES��;�2a�\h����jb|� 8�W�9�Ai��jb|�=�_�3�K`��hg{�	
?�_�5�Mc��i4Kh���IGN -�>F�l�1Mn�� �BLE+'�5J�l�5Hh���JDM#/�=B�j�6Jh�ﵷGPRRh�7�+��|�㾽NVWQo�:�%��z�㿿OWTVj�7�)��s�건CrC�!��40�4������y�}L�,��36�3������s�tD�)��36�3������s�vG�.�1)��
�B��n������6+���M��j������=#���M��b������6/ߡF�_�	F��|�_��Λ5�ժJ�U�@��}�_��Λ5�ժJ�W�G��q�R�Ɯ0�ׯM���>��T������aϪR�7���2��P������aͧ[�<���?��U������bϫR�4���5t���I4�:x�!�#����t���I4�8{�&�(����| ���L3�6t�,�(��������ām���=��u?��Ǝo���8�ʃ�u<����e���4�Ŏ�4���;�������6���l�l�`�6�������2��ʟ�f�k�`�6�������5��œ�b�m�f�2���{����X�ܡ�+�+wS�01A�{����V�Ԧ�!�&z^�=<L�q����T�Ԧ�!�&z^�=<L�r��%�-�A҄����V�\��}�. �-�Aԃ����Q�[��p�)&�+�Fщ����Y�R��p�*'�*F1��;
�=K�ˀ�/�ޑL:��1�;zH�ɂ�/�ޑL:��0 �=rA��%�ؔM9��0�3ߏ5o���/�d��=�1ޏ3l���-�f��0�>܊4i���,�k��;�8ԐRDs,�o�_(���6��{z�RDs,�o�],���?��rr�W@q-�j�W!���;��qp�ZCv��j:f���䟖�v&+�q���a8d���ᚕ�v)$�~���l;b���钝�~!,�x���i�Ċ˱Ә��|{.�F���Ìϲј��x}
 �L���̂ùԞ��~
#�J����Ҕl{����6Sd	dx`͑x�ܛl{����6Scbg˖p�ԓds���0W`bg˖p�Ԓfp�(�W���D�	c��c�.�#�Z���O�g��a�,�$�X���@�e��g� �+�V�:�tp�l��b!����74�^�0�~y�f��j&����74�^�0�~x�e��o#��
��64�_�3J]��2{�;3ۭ*dyM�3Aa L_��0x�81ա%mwB�>Ba'L_��=u�61ۭ*dyM�7Ln*G]��H��yi��^>K����$� I��yi��^?I����'�K��xk}�|�[
6B����.�D��s��x��\}�J���r+��;���x��^�J���}#��7���q��]{�M���v.�<���{�Fm7�v�"�\X4�i���Dl6�v� �	Y]1
�`���La:�{�(�
YZ6�m���Bk0���39��OB����$����43��AB����.����;>��IE����.�������D���&��<��������M���+��
>��������@���/��1����������_N	_M�����=�ul����TCRF������8�wl����TCRF������8�wn����\K �Tل$��,E���h��I��(�I@�u��.�}��֏X�(��Pɤ���(�~�>L�d�%!P�4@��B!-�6��D�$RV ��|R��>�r'AMAI)ǥoK��"��- 8u!��5F�����S'���1��U���C��_��Q���4Q���3J�����Q �����P�2噹Aq�L�c#WL�R��E.��<$'N<?fy�4j��Y��嘻Ey�l��#�O�T��UnP�+T����F�z��A����iV�B5��(n�Չ��i��(��mˡP����L�>�F�r�J2��'�̭C�Ñ\>m�B�ŏH#�; k��b6����ѵ+�X������̥[�#�Y7M�r��M& �`k8a���g�*@���*"Jݾ&�$j�y��Rԭ��&����w�I	e�J�̟6/�,]8So�}vNX��˝��Ht�2�6�p�g�l��Q�alE7-�.E83/@�|uVb>�j%���C�!��0*��:�C�l�'�\]�࣑%C��T{���������T��aPl׆t@px��(�,y�e�g��2�h] �D���^�҂���ħO�Z�i��y� �4;]p1���&*
N5��ϔ�n�$דY� H�`�!l�\��F���ˈ�[,a�J�5|���A)�M{�
C	Y����#Ѱ�[��́G�8Щ0eʹ,�$dj�Z86��48t
B^���������l�v1�)���h�RL;!O �x��)�#��w��쐶�D��uGo��sG��h���%12��2�M�?��:⧊�n�"�gf�w_LIX ��( y������tlV�Xǅ4��)"�$��^������}�|k� ȔmĪ)��)�9'�� �g��@�h���[�X���K B	�~q���b�l[�m�:d(�CϐG�%���>�^��}��m��ol�q" �`R�ūU�X8&�08;�i�0SH6��X�"�.�#"(�2p�4+�$�1X���q��3�,F��	Gi�@6Aj�oDh���3&U/o.�a[�D�W͟3�jQq�]�0��WB6y���!�*W7��)_+ �\�"b��2��4��B�Z^�*���&��3��:"�e`+�X�*�'2��b�0:��!0�``�G�v�A� Q U6J9qc� t��qh�A��z���@��%%g�p�J�J��)1�Sg��\ZR�ۀE��l��,:��D��m�v͹�K�=fv� j�o�42�L���.֞^�\�3���!D��Y�j��I�f�'�c>UKTi�<a|�,���6 �)�7j.O��	�l�� 6Ψ & ��;�Y�� ��(��<���z h �@�9`�r�.}��Upa����ZU����(�$}c^,"�˟���H�Τ`Ħ�=u�zm�e�
�"�h̤��O�,� ԆL}Z�['U�4�δ�U�Ao<�Ɍ{���'�R�9P�B��L8��N�}�:��6�՚  �1��O���aLw�g��,L��x��/w�J�{���)�`C�	U*�H����T^��j6GN,p��B�"Ʌm��h��k�xH4�Ɍi�@p��Ą�	����4LO:�ZR�zsЅp�'��#�� #�M�ekG:3.�0S�'��X7$�	�>� �d��/_J욋}��K���F��Nˤ��=���@K*����֧�y"b\TU�b
C�9%u���E�y�]WT�:�Y�;K0�)�O�%�yB�R�5�L[��y���@B�^��y��B�=�4i�T�&e�hQ�$Ŕ�y��Ra������S�R�q�Y�y��ʌh�.�26I��ޙ�Ȏ��yR)������	۴q��1A��y2�H#
�Zug㚀x)�i�����y���@���R� �#�hї��5�y�2<��(���"��] ��y¤S+�h2�%L�w�жH���y X=��pr�ɥ �`%�yr�ÜZM�4z���� ?@�"e��.�y�V	Y!�u���T�v�,ڡ���y���W$-�R��F	ۡ�O��y�A��0�������E;�S��y�AķJ�4�!cʽ?�V%�0ʅ��y��VP\�B�AV�+^]C1���y�)� s���pg��e��U���-�y"�Z�L�^���jT�U?�icBNL�y���{�8����2s�~�`�L��y�M4n�YRF,�w�R%����yb�EEX�M��g�x�F��fȓ��y���=7�+N�Nx`);c(S�JwfC䉺	ԵpE�0�n-J#cP!z�C�		��RC�G�q�A#i��e�B�,\j��U��.�^�Q`�͹U��B�I4]4pYaF"W#,,D���r�-D�0��WO�@aXԧ�6=�Px�"*D��ӕ`Z�B0H{Q��D@��¤�(D���B $Iꜵ
uI[�Xz,C�&D�� B�R'�B�JP�E��� �f)��HW"O� ��dߪ �R �V�ڵ"O,��� �B�$:TO��;�.���"O�dSv��).vLL@�D��P\T�ڧ"O0�n� w��=i�
��NO�"Ode4��h�P��)D$[���X�"O��V���(#*V���"Of9�Cg�j� +�e�̍�d"O&�Y3��F@L��!�٧?��<R"O��[6�V�E{<՚Gȇ�`����"Oh 36*S?ff��3i	�	��"OZ�z��|A<m��G�
��2"O��1��,b�r@��15����G"O�0;� E(��S�ͨD��aa"OP�����t؄�J3dީH�v�@�"Or�J�h�+�����~�8�g"O����*�^��99"bޮ$��+g"O�dM̋IE���	��hA�"O��25�T��� `P 0a��x9S"Oh�������S�@]����B"O�}S��ӧ|H��r�J�t�pR�"OЕ"`�X@,x�oږ_֡y�"O�Ő��KĈ��N�r���"O��1��ڊ.&��	�(տ�5
�"Ob��F��7��Mbq$��AT��U"O��;�@� *��*��B�s��9%"O��
҇@=G�3��HBT"O,8SQ�ŸS��T�4H,�""OnT����'>[е�@���fM�L!p"O��/ո�� 7/A�U�rL8�"OZ,*ԁ��C��DB�$�"/t���g"O\y���`�0���1��Drd"O:���I������=	�=�C"O�0Ҁ.�%/����A�/�XMS�"O��`���7^�����QA"O´!҇޸z���7`B �� c�"O�"H�m:񯗟2�R��$"OT�����?YY�I�M]�Z����4"O���5$��NɊ��4��1z��j"O����YJ��ꅉ����HɅ"Ov�Z��٫&�TQ�գ�$����'�(s�FԻ�Te�e\���`T�J>\�b���Zdb���x_(|�4�h-4����a�l�?��l�\�`)R�5�\db�):�	�Gc���6D��!�0�ē�!򤇖M��$�5H<T.��[�ȮX|x�j�^���k��=wN�����?Y�m�0\9.|�JT\��X7B�L�<�v�6c5^���nO@�ȹ�V�Zm�`#����!�I\�i2�a�fAHv�'��7��!��Q9�oߎ	_|��
ד}W���7c�[~��*�LU��d�)O�3�����(zG�������O�� �O���?1���+����W�K��u��<���c/�<l�|`��2��'��D�d����C�|�֤�7J�[��{.��I��B$�Xg+�6J4�D�SH޴-�.�X�A���u���2���MK�#�h�}���p�Tiz��SSx14�F#�̨@�+�%b
\-y��0D�|�"l�H�'E��ͻJcx��6���GBXj�Ā�A�U�d&ǚl4t�Ja�D�$O
� �,�|��+BHLBJ>�pÜ6�4��"�rQ�¯30�9� �;L	R�N�>Ժ@����d�v6�x�AV���t��(>�d��5E
�0���H
+/4�Dj�["`Q���� z�O@̊"E��G�*�)���F�B!a,ÅU��0P�WSp����U�"@p��>���6��� ^w�vyY �
����cE�)'.���j�Q���;Q�I�4��D�Ë	�ē?jj��@EƔ�@����|*���V����Rg]fad�1��Qd�&i�&!IVE��4J$q�@�I�O2@����bWtA#S���i����QÝ3Ĳ)�Kݱ}����AT�<�Q�l�5��1�g+�JDa���)é�yW��%|o4k n�E@``q�Zq�FA�'�a���yI_w���	P��qP&�Y�����ӥ(0���c֍Wh(��Ќ8�<A�!4t���0/z�3N�$�~��G,5�U�3�F�t�*1A�L,d���Є�D�D�>�HsHa���*[�K�PH$Ӌ6���@�TLՂ
!}�N�i�LH�ab� `皮H0d��U��#2��da�DYq���$S��1��!� �Ӎ��:D�BK�WI�"b�@�<dV�j�0S�n���>{�8&ƕ-�~bk�=A��c��2�`�ن�X(c����qD�A�� �3w%A<-���%� ���b��0w]�"��_�|XYB<$��![���>(���]?)�wO�|z��ƃA�@�*9ZYTCu��%T�d(8�
��f�\����ų��I�*G��Je.֗�@�ɮ`�p��� �<��bz�jݲ��P-��d2R�ӢL!>0���w݅y�£:��|�Ĉ���y��CE�L�Ůٝ=Jn	����G��`Ũ�#^����d(��I�F/�2w�'�@�X84h��G)C&��gfلOK0�Н7������~n�e�d���ʉ,��9�JB) 1AP�u�"�/p������(C�H젃fQ02jll:3`C?؆�2$L8l+��F&2:�ˡ�ɫE�R七��6b~Db�=Җ�J��	c'��#�N?A��듦ܜu�Ή(V2O`�a$M<;d����]	`&��3��F>F����&�t�ʅ�)�EI!�p<f��#cߗ+���GQ���0ף�:4�a�m*z�u)�l�p<b��3�O���hB C�P�Z�E�9͆x0gl5s�80P�*']��K�숆u��X�B�B�V�j�E�;ŒTXg���t� l� T�ʜ�&�M�o!h����͘F�`��ͻn��L��"W�>oڀI���ug�Z$5ش��u�y"@>1%L�Q�#�-��u��U0łu��g2B=�B���[�.�ES,Y*R�#��*��U�S�Q&�����cª���W�+ъe�X�cʬ���Z�qzp�����U��5�L���y�gW*�
�ؑdǨ����r=�i�'�GE�p�gO�g�$��c�yd� Ԡ�z�n�1��@�l4�I���ƊA
�`��֜`�4��ܕ~.�BUI,Df�P�ʟ�.�����bHa?9S(ƻW��]F�F����#7�|�+5/�ayxl{A�����}b	ɸ[�L�+7ִ��s /�'�������v�pQqoM���UI��H;^�^�I�zh�1�_w3�z��v�%��(S�8<X]��^"t6&�p�!�i�"��S�ԴP;�bW�s��6Ȓ�?0BY���sǈHy�K#)dvp�Q�mx�lXHtƴ$����˓ W�	���
"Z͂2)>9)%���}�`� /(�.�3� (\h�W��%B���=;-=�rA�x�B@��tJ��D�9l9"�dA娣>Iwb�P�>}Zw�P� �%H�(ͣ�TxXC�}z�b"d�/H�2�9�"T�m^��a�+$G����B�$&\��Ɓ��xl�*���.J�>�qb�iJ̉�J 6sI>�aƊ��w� Y�QMD���w�$U�a-��S�6I�2�V�zRΐ�o<����Ձo�$0"8S�RQ;v���ȌL�R��!+��SE�T�e��mH �I�)��B�b)ړ"���:�O�*0���� :{��H9�oIn?���W���tKzB~�GaR�d�����>BD� �d��t���z�H�;(�,���ƍmiF�W.��$䊠��ɻR����S���5h1bŉ5/,�ˁeK*9S��؂&^�8#��8X���Q 1��XAbE7(<�93�l̸�#�(QD�Q��gL��B�I�>XL�fƾ(���yBi²4�"���C��h&b����ٙ%�0;sn��X9Tl��b�=-���1©��6�(푵�'� �	����L�x!�a���Q����.�ƣ]���P�+�%6b@�PS��!��I��BQ�tA8e�V�`#g
%��i�FB�<qL"Q��i��4qR�=1�D?XC��Z�&>77�-���E�Ɋ}k`���5)D�����8X��6M�pL*����)���{1��<P��܇U� +5��:H���#�O
��Sb�Ls���Cϙ�@�n�*�A(<(�옔�ʈ=��I�,.t� �����Hy����/مC�f�j�>�
��3�J:2;�ER��Exq6�'�֡�a!Q?��B7;vĢ�+P���.+iu�h �lq��膆y��I�c�5;P��!cקZ�bt��-�6u:Zם�<��A�.�L�D�E�I3�U`�Ϟz�	�H1�Yx��:���e����h�)�F��w �M>~�����@�l�D�F�V����
-��d�i�b�(�!@�V�~�s��	r	9� K}�&�0������L� �� �O�Sk�x`0�;HنX������AEfʄ6������q���6]<48Bc\>)Eh=ض�A�M�$H�Ý� 3��r���m������e:���\�'0����o�=[¹��Qi%�,ڴ��J�0����MbmĚ@�����5��9�\1R�A���`��"���u�s},Q�FS!vA���Pʏ�\b�� �����D`"Č�F�8;�TF�B�⦣�Ue��+�bZ� ����6�(k<����?(�%:��o�\���Ê�Sn��C�"#������<	���+D���"c �*>���O���& �:%@T�3�� ���(E�޾Yc�fg��	vx�o�(
rL�GV�a(l��M��%��Z����?tlQC6�����;�i�	��4`+j�	�M�'�� b��i���S��'��T���uO�i�ڿ:m"iJ��=3�!�$�5����R&���ɞtB�3�=<�H�-61ї�ƛW@�Rm�-7����y�x�I�E".�F�Z�o�o�j�)gBm�<`�M���ʤ*Ŧs�.L��&1���k�.�K�BPZ��Öh�"\b�-������s�.\1�K�.���1/�=-�F���#F��u��� -���PY7`}l�UY�B��F�9��B�]�B샢b�|��CVd�2����ſ).NY�gΟ8dG<U���Z�Y�@�BT��[VDr�Ŝ��Z?p�4B�j�bY�������	.6������R�Uza󳧀�L�R��-��yA׶9v�zF!3+6�Q�� ),������`�@"C�6���AbL��i�,&��A++���dh�-f�F�MX"m��ɂ�ը��cH���%�X���/��T�KR2q� �	���#a@-z�(]�ga�Jp�Z� �.Xf�ڍ*���� p��C�M	8�8&�)`l��<)�(�"�т&��X�N��!	׿.9
9�w>O�D�UN��~�B�P�~�.���FΆX�Rى�ɖ��MS�/��9]���4b�j���סnW.EHr%�:SBlvʆ�;�~O���F��|J�jD�K$
J��i5'�>-��#�pdM�6�P*v)h��b��0>�д��֔kn�"7"W�+��3�M�qbI��Ыu.dŋ�����	AL˃n���iF�
;�ɖ�0)Cj�I���<%�u9@�3��d���b�����n1^yCd"Lb��i�)x�|���CT�F#��$&�a����Wn֫l;HU+���Ij��)Vi�}�lU!Nln\�����(h
�y�P�%��&��5h��p�2f�r�
eJ�!Oh`D���Η*c��h�'%�\�u ë~�PS�/X2cn8d;RI���ğ�g��l���H�@85Îi��Ox5� -	�͊�Aao�mM�A���L4݂�:	���ݓ���h9�x���*Ô譻f��)QF�Z�0�(LKr�19s�m	ܴ!���#1���G�(��]�/q���EM,}���Q��g
Zk���g�0j`���R!�W	z5�uoӼx4�&.-�miu ��]�(��gA���ue�*��S�z*4�f����Dϡ�!8#gHh��K��?�dN����[� �?Q��)d�ý`�(9��?q��s��H�HM��	�);�ؐ�!�p�`����T��������.�LZM�Ze��ɉ�<������'s�n���4� �T�rh��x1�Q!�' c�bٲU"ȵ,��o=(��0(lV�_�^,�FE�O�v����A�`ђ%K��h^ 86�r���s���r��&O a��q��\�8�8y�W�l��8x�� �q���� S�$OTUC���(7��k��R9�m�� 71Aֹ�Q�'�&Q�3 X�NREk�ĝ�2���R�>�a��@ԴUn��`�D�i:���2@P.e��mU�

�V`��,,�F|�L�n�� 
퇆Y;�Y�f�=��)��:u�lH�%c�bd"���۝sf���Z;�I���#�\8o2 x���V@�J���+'f��@��G�'b��@�T�%����a�
_7"��V!G	���rBQ$J��V�W��J�af���.+a/@?exb�ipHĝe���B�ѥK��'W��P�	�΀-�8���&��F��y6�*v�6�!�'m�LY��b>�2͂�4�,��D&��B��AV�*�u����:�k�IV*b��pc&Z+Ă�x���?d�n�2�4`�x��2��x�LүR�\}a@Fw�P�Q��4S�� ���2{T�X�o٘0�(�a�%N
 Μ{3���P�y���0]�ȩ �:0|T�h��Xi�=:��8�0P��@������" ��x�� 1 @���D"(.`��WӅ7������'��%`��">q0�/�{$=zr�܂��8��ӄ4����7��#��O�N��3Dx�����b�7(Vܚ"�	4Rd�Pa��&.�|��U�L���hk�f�0z$y�E[�5�j� WE�x߀�_��4�2�H�f�F��ҤK<oG�O�n�'EI�}Ք<�gӚXw�z�h�.� �g�,�p��+F�j�zp) �|�k
�1clűg�� �D ��$*�N��M�'�"]�i��R��p!߿|05zp���49� j�!��ዧ�  ZKEs�H$����`(1���@� L�����r@�x��4�@"z2UA�#�.���)[&.�K@�I]�h����v}��qnH&a'�m���I�#]�]@T+�xR�k���{��ňO��@�c�K�6�ۇKB�m��Ͳ� �?
�D2��:y�<h�F�-j��� ��V�.��gkÇj����}Rq˅� 6��!B��5gM��C$���Ol��Pd:C�6�}��I���	vI�f��jY;���~\��`V�un�-��V�b*�Hч���OG�����6��&F-L!��W�S75���J�[}�O�x���9����W�@�u�'F��gI�ES��'Z�0����+g�xВ��I� 8я�>�J�-�-Y�5��l���8����zԂ�y�ʌ���ArCNZ8Z`�(�&���B�oݥ5஝�Uf�@���:J~�%��B���2�'|��a&"^3L��l��qm�idG}{�����3:8dX�$O��Q�OB�&�+��6�H!K��D��0�+��S�g�zu��T3-B ��OyyZ�b>1�m�R�����m���z����%OJ�۳�5�.آnZ��DlC�E8 3z	�4�m�0�P#A�%��8!1x�'G24�0�Oa���G"9AK��j� ��&�>I9M<���lEh]�����L *(	P,1�t5�a�$���:VJ_�JX �BrH#���H���O���pb�>;�}�vDMC7���g=!��뱟���M<���ē �� kΝt��H��O��(��?V~A��܇o�Z��M:�z-�F��v��i���� �0>yŮJ�i�L��T�׊rڐ�i��Ls��|����lK�<H@�O�(�2�յaѤAR�A j��*%"O�@��DӍ*849Z�!*|I	P���^P�#����蔴h�h]4�.��o��?�!򤏍?�D�U���o�T�eΚ7Y�!�d}e�Tcv���G��@q�'�!�I s��� �(Ƥic�̢|�!�d�(23v�G��<P@���r����']E��)'��@*��׮>������o��8�.L+�m�e��m�<yvaE�l 2��@��l�yBM̶�X�X�L�"�Bc���y�k]����wH�v�f����y"�	[�X1�&�dI��C��_�y���)J,�9�+B�Y����+�y"�J>,
� AW��t�ԟ�y��۪S��e�� !x.��C��yB��pk�5�	.Aأ�	�yB�W',0I���d��K��y�.-)tX��s/X'=�=��D��y��J�V��a�KȾm	��k���)�yr�ރ'e�I{KD$d'���֌�y2��)p`v��AÑ�@G�0ywo���yB�3�,�Y�FA�4�l!�ǒ��y�K��Q�Ā�Jߘ�fp���.�yB��Z(�Q4D�y"wL��y�NR,[��%`��^4W���{�R��yRđs/P�9ċ\�AJ| �&㜤�y���>������Ć/(0���C��y�d\&t����c�\(3Y��Ô�E��yB��5y�	��'j�C7�y
� �m���>#߆�����+.l�s�"O$d����K�P�چ�v�x��S"O������~[ !0d�<O�pXzc"O�ȓ��=߆)JT$�f.�Y�"Ol���/w�,���D^�BH�xY�"O4����-�� x��2*�>�B�"OB��Bɲ[��M� �Q,lu�X�"O���T��,e{�<��@E�*�|1"O�,*�/��P�H%`#��٢ "Ol����.��+Fo� h�}�C"O��)6�Q�!I'Kb��@��"O�ah�N*lm���0�ːG\��"O`H�-ߤL���R&.�
B:�|s0"O�ٺp��k��U1���ի�"O�tҒ	ނ��|Bt��"v�D!�"Or��a���d6\ R�usޜ��Op(��BJ��ĝp���8���6H���\�{P���̱W��h���̡̓8m�s�
/�\xЊ�6���T*�0[@T���'�J"=E�4��" ,�%r�ǘ��R��"b����S�c�m�݌Pq�ɷI�AT���?%�)�&�1$. ����f|�7A�������>�2��H'i.������k$t 5�<���)�'G��tK��8?��G�;uZ\|�	7�(O�pG��!Ĝ(~HX6��*v��a�&l��Q�9ç}<iQw���]�1���Y�z �>��L6�S��J�`q�m�j��4�Dn�./�OV�a����I>E]JM�"J�j�tH��*� Z���Q�Q�"}J6�ԒXH�c�� d
�4��&����Z��)�iA&��@نLv�h�4�X�B�n�!
2< �/!? cT�e|H�t�O���ӛ'^a�wHL�b?��f�[I��q��5�$�� ��\��>K�n���M��m��eZ6	[:��O؅äLR6����Ot��T� FTr}��i�-p�lY�O5Γ̸�H���	���"'�x2c	XW:�H���i�0�ɧ3��䯟֝U�O&� ;��ׯ#G�����(�$�p2O|�2�';��E�'����1�=�|p,9Jd��*�d˥`r�执�yR�I�<E����d�����_R6�T9%v��7����+|O��Gڣ^)�ʑb�"IM���"OfhA��"3\�ZwB�j����"Oԙ�4�I�S�(�9��&��`ڳ"O M)�g�4g>&D"�!)ߦ�Q�"O�:�%L/Z!����,"E��4��"O��S��,&Q�!�q+�*S�|#�"O�B�О>�'�ǣ-�B�"O���aڱ3�������iV�M��"O�0
%�֥��yr!���Q��G"O�J�A�I`D� �X�~�9"O��R�ʎ�)p���ϜsX0"OZH���ϊ:�D��Q$FC|2"O @���t�) Fi+\�X)b�"O�y5� (G��Q*B�O,,�"OV		u��[V�H���2E�~���"O�Y��F�Q��1����c�QW"OL�y�Ď	Rh�`���BN�P"O,ec��;�(�r�ϙ>Ev�s�"OT���E{�iP�#R7M*�,��"OT!q�4:1b�#P�(w!���"O��
��άN8�0����L��I�"O`\老֬��!y�iը$�b"OL��w`����Mۼ]�<�2"O �	&+��r^��e|^a��ł>�yR@�>i��i���0&�EhFM��y�O ;t�R���O�(JL�����yr�^�a�h]1���(��-�A�L2�y�@��!��	�f�6y��A��h�"�y
� v���Ŕ^�I�F'J���:�"OR��E� �G	@�!Tb��q&"O�#�#Sxܑ�Wg�<L�bXq"O�����=J(U�BOq� 8	"O�K&�L2s�Z�+SeEZؐ�a�"OZD)R�I�p��`��ƏX�Z��"O"��P@�)Ia~%C7��)��ňa"O�D[�i��Qc\�: �_^  "O@����/JR�ؖɄ)#.�3�"O�x�&�� d��`�G�<�ȴ�s"O�9�Nz�0���  �`)��"O�,Q@g�4�E��2��j�"O����h�� p��"���#"O4 +�3%ێqs�)ɞ�y�"OB�zhۤq�إ!Ɓ4i�"��"O؉0�)N�=��ꗥc�(��"O
U��ŧ/�J	����+���� "Ob(1fkؚ\�
xq��/H��"O����i[>#xqa���7O[N<�"O�}��X�f��[1G�,wf�@b"O$mb��ʊe����!s�UY�"OjȊ�� ��Ћ���3k]lL��"O�  wA��R	�PQ�"H�i3=��"O@5��LN5PjZxHYQ�^� "O��X���r~�əԏ�99Ӛ���"ON��/P�E�z̉���>��|Ʉ"O)��d�:�ȡ-2���4"O����Ρ�!��F�5"y慂1"Or�h��G"`�����UN�(#"O�hA��2~q��#�P�yia"Ohaz��	X7v�3�E,�P�)�"O,�����Ш�Qt��<�RA��"O~<�"e�oh<�Ҁ@M�ߺ���"O����8lǲ�d�/V��X�"O٫fI� 4 kfLG;�X�Cs"OLEx��K�VF�t����`QIp"OLE��ُ} qz�D�� �0�*F"O�s����c�Ƭ01Ja�ڍ�"O<���EO�;M��rWHP?(z���"O�P��	��jg�] �"��"O|H4��vm�|�%Z6U���BF"O$%�#�� `���z�đ�d��А#"O0aJV�F�s�F�ɂ�E�V�	�"O�����Q�	���Y1�ő,���k"O��p�MD.b�ĺ�� ��a�"Op�ip���`
Bz���93"O��iFM��D�}�bF5 �v�e"O�
�) r�p�ٟg����g"O�M�a��졐4bӊJ�*)�"O>���X�.�B�PB ʜ'w����"O����-]jC�<SAY�nb9�@"O��cf\ �Ճ�Μ$'��B "O�yB�^�@�Ҩ�@�@�.xL�Yd"ONu��G�#��P	�K�L!�"O܀�'��d���0̝�?��}I�*Oz���E F@Z\���9_
�X�'x�tk�>b[�Ѻ
��B>b�'z�l
� 4Kz���'V�*��T��'d�A)����[Y�u�����Q�	�'"� ���ҊU��|��fX7 ��'3��*�1G�Z��ǝQa���'RP��M�g
���Ry��D��'���������3��.׀��
�'���"Q�߯q����fe4k��
��� ��)�W4�CD-�	^ih�"O�,i�BO/F�,�0l��Zo����"O$ Z�;<(��͆,:Q�qӡ"OԱ�M�yP��m�;,P*�"O���(ɉ%u4�'-@�M*��8�"O��� ݪy��I�B�ܸ�Vu9�"O��֭D�9s2���n�_�6<��"Oț�/��zVՒ`)�\��"O��91����{���Rh"v"Oz����!8��2띎8&��1"O.X{㦖�Y�8�I��ջ�X		�"Om*g+\I	���/��@"On�Ґ���,u�h\�@� �"O��r�K(7x�a#gJ�U�����"OD%0tƌ?V|p�)G<|��	H�"O��y�+&\Qۥi^#^_±�"O���ϸw`Ν����51$��#�"O\H��b��	c��y%�yp�"O"��s"��1>�c0�W2�(9�"OjY��!6bԤ�ȧ�F�Yh+ܽ�yRhYK)� ����+%�dA#O��y��ŀ(����_�rF�2
���yb�5c��ٖh	�9M��r�L���y���+HA���)�z+�����y"ň!{�T���@�?s���։@��y�HD��I D���)iժ���y"lB�N'h�
T�cP9z�KQ��y!*f��$h�.q[ʥ���yr�
)���d�\� gb@r�f@��y�|�l���L�&�аGm���y�
�Z�b�r�T��D`�c��y���&�	�����~O�������yb�4~{���rk�`���'�_�yrCV�:����YD��u[g���yrkߔAb�E*��*O`�\0�F�8�y��T�Z��Y&'F���`�h�6�yb޹Y$θ�Eȧd>�`B"Ͻ�y҄>-"2�jуНdqjt8"+Q��y�d�@h��HR=1�(\�!���y� X��Xg�T�T�Pő�A���y�
�Z~{���� _�|J�a@��yR�I*Rf���^�5PH���9�y�B��,�t�A!Iܕt_b���D��y�S=wnʍ��fbǶ�KF&�yR��R��ClЕ^&�yp���yr�N�(�rQ�A	�a�קB��y��H'IV�H&�(@*"��)Ō�y��ڊ<��+s���=W��H�E�yeK /(0��mí.2��V-�y�
�<��E�%(���m��	ݷ�yB�.4S:L��L�`_��3#b9�yR�ԫz���*�B���}�c���y��'��rT4���I�
�y*ΤF3�9�c�^�gh,�Cn�<����5ޖq8&�'=�^��4�J�<��%[H�0ȇFǢ �2Ċ�&I�<)��ŰJ>�D&O�y_��@��A�<��V�
`4�9�D+:M̉�"�w�<�&�X�ҡ�B�R�sl���6!�t�<A�bD�y*Dx0���9S�ZDjw�NZ�<���;�X��A�]�L���S�<��<�ֹ1n� W��"¬�O�<�eA�:J0D!`X�Q�6�r%��J�<���y��;Om�x�B�[�<� ��k@�9`-6T�p��D�BI�6"O`��%JҖb���g'X�+r�};�"Od����so؁�TM��	��v"O$(�.� e~v�FL�?<��#"O
T1��R�	�eJ���27"Ox����=cȖ���bP)6��0�"O�IR$%��0�4H���l�%Y"O�d�V��Zb��Hp*��!d��S`"O:�2f�_"o\D�"#�7;N ��A"O��(H�� 5S`S7v.&�Y�"O���Ӄ�q;(�2`D�64L��"O��A"c�f \	kf%8@����"Ol��ᇐ ê����7Za��"O�Lh"A��8В��,Q�5K�4"4"O|Ȳ�A�=o`	 ���*.�1"O���5�L Xhh+�@�,�<�b"O�������ctE3 僌[Dli"O<dy�Գ}��8���7sb��"O p��f)(倆�M��6� �yBgX���<9�d�	M{��W#��y2%�5��$8!��X;�)��� ��y2ʊ_��sp���8y��C�8�y���9��nV�>���.�y�D
5\���7\�hRsÙ�y�KFT�9@�
}��u�K��y���T�#0v0\�D��y�gƗX��8( �N?q���B��N��yR��@|�(�wb�o��� ��ջ�y2$Q�`�Ԍ�t��$aO����yb#-Lt��\�]fR(��"�yϋ�Z�@�i�cˁb9��r1G���y�K��B?�h�w"�)������y��'�x͢%���,��a��cV*�y�7(�fxP��G%9����Ԧ�y���ld
��F�&�Е�B�9�ybҕc��e�po?F�,P3DA��y2�U�8�RqGnս2$����#N?�yrAH�}�s�c��%��5�a#W��y¤��^BT���Oт8��� 7�y�l�;��0��o[�z3���c�y�M#/�rM��&�%�@d��9�C�	7-3�ܣ��q!�|!%C�"y�lC䉥x�h   �