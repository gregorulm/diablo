MPQ    OC-    h�  h                                                                                 �1@=�_��LI�VA���3�ƕ�Չd�i�b;T`$�98��Tr>Q��/p�4[D�bK���T�A���e�GL��&�2�d�5y��Y���,a1�!�T���/ӦYK5;:0�f����mؤ��)yDK����jChc����Y��f}I��)���ˍ�\@�1��>fm�3�StU�G�g#j�De���T�3��\Q5q�������o�3s���u��P��ŭ���Ł_I$T[J0d�x�򅢀�ʂ��T�0n�AsM]ux��l�2y)����m��n�?��E���(dx߁o�i��&�)�b�d점+q��{�5�7-Z{��]����^� (��c;�B� '�� �i#+U����/��m�%�-W����L-������5�vڴ�Bbs�hx˅}�q+���������H��h�Дd/?��-S���BE*�u��R,�(�˜��rP@くp��̓�vL{�#��bݳx���3��C�Pz��f�"�i�&X	��I�rB`����PP8V6���G����WsV+w�G�F)O���m�.%E��Ed`|��<hb{q�6�G(VMqk(��ӛ��a��gҺ�ʞ\߃�ބ�|%�-'�¼���1� ����
U�|}�2�5���R�"���57o}�&+�$�(��P�+/�>En� ��zsn@��Yq+�Z�~�G��4�޶��g�en�=2���^�4�Ǫk7�С��찻���
�3`�QZ�/�5��ooUyt2��&x �b~��,������K�↧Y`ZvUt������W3���Mf��"S�lE��j�tB��_��H��Hu��|Al��y٠+`�xD�z�S�-$���Ƶ��fw6V����d����#@w�a�"NX�W��m����f����f���5D
 �B쬼Z����Қ��;�k��ܟxG�Pa��REzS�˗��i��/�z.��Y�I0Ԉ<�����%Wqo�&cf�da�x�2�>D6)q�%�>!��QFT8�2|�t��g2��C���=PP���(��P*|�ݑ�y��� A#�����`~��1֢/����u�q<ϓ2�[g���%Irغe�	��M��î�
���L���?��V8\*j�Z(�B �n���&�T�Q�`��lޞяv_�8��ɫ����
n֐hE&+l�H����!9�=zS̈���;�u�Y	e$P�<�P��}fB!B �1����ڜp ��).Tl8��۶���N��X���C����^��!��-�D�?��'��r$��m�������ԭ4�%D�̡�ˇ�H����а$��t�&e�
�\��� =���j&N�s��[�S� �2��:v�HB��鞃1���j{����|Z-�zC���Wf����e�3�;v��vF���a�i8ԊT��=�$Hّ�C��f�Z���	X����3u�8��^�:����N�v煃��K�ŏ��TO�RӖj������͟9]{�|�ʭ$P� f�`��b<"�rȱ�����np>���*�?�?�ߧgx�6L��tl��̟�rNSy?����Qdp,L�a*k�*Bus��׍�w�Q�S��F��
`�8�h:,� 회�C����C�+C�� �p�ļ��c*?��m� L
������&ǣ#Y�%mu�Qg�C��\ͥ6O`h�+���z3�\8<cxh$�$]ō
�acVp�t����`l�H+���{2����O�$���|Y&)�B��1�N�M�B��]��ڲ�����4˲_'+[ۄR�Of�8�̱��#� ���9�8H�X��)^�n �D��8���gm�,#�]4�T�����
	��?%��.�rU�b�B�]���L������6*����D+�91��+u��� ��]�z6��6>k����Ɩ���V,3KR�R]����EO���!G��e���ע�ɳ��8�0��՘�:��;<1M��-�|����ړv��m����([C�J��/�5n�Ӭ���R���SV����Ւ0�d�K�b�m�z˂���دs�����ڞ�`��p+f�rS�%�ʭ��B^�	�N�u
�+���b�~�1'w��FU�z���X�,Ȳ^�y����	��,7<��:�-�R�;��Y��L�c�0��Y8p]&�H�K�Jsm���$r�`୨:�N&)H���ڀ1��{Z�O�&�x�\e=��C 6&f�i�3ą~�A
ar�*Y`�l8�_-#;�{���H��� =��"��	��rq��6�sW��|�Ζ�z�X�~P�`]5'�,��B��4;|��F]�ұ�A��_]��U�R���If�,�DfZ�7����Pb�P 	
��Ѥ���ꗭMjId�X�g���	�n��$0`2�M�J�?���+	P�d߬���*�_5�vHėP<�)P�N����\��:��~�j���nH+��DK�!��0��c�<)eFw�D�S{BQ�׮�>�P;���Ph<�ʬ�Aƿ�`����7����˲�Fw���������w�c.��q��M�Btg]+��؂N���^6B�ۭS?r-�F��~���)N,��/ɟ���߈t9߉rrO��x�2� .�5���ъ�F�n��u����5���%��জ�^���L�_����+D�C�昴V~�,��9N���On�vá�Y�׹�L��J�[Ob�4u�my��	�sY�F�Nh��]Xu/;Z��I���a�U�6����C.(�w��Q�p_�g�.!bYl�QĒ�3F��*y5CP��O$�u."���:�Y�|�=�o��K�����[XBI]02�@22���_�$�y;��p�9���B�mhQ���e��7>�6��D����S-=��\Q���m3���g��� ���gT!�G3�#��Rr�m�0������
��.��&�Y/!�h�O~���~IFK@3�-��*�����~e���%t9�d�)��Em�i��Ԏ������,��)TW2��dtJ[�^C1�����̎�u=1�;�@Z�/�;��VX:#1��]_�5B�9�m�	H�L��P�gR?2�Lq�Y��(��!�h��|���8ú"3���A����ʺiٟm�p	�#iۢr�שP.o>���!c��-�}@ݎ�Xj�'$?$�^�D����m��3$�޻��H����g�j�ϭGm��`��y���a��u���hUE����p��c��n{a������;	��MV�f�(#�M�����~@�A�7�L�JL�\k��ZpW4r ����.���b��ԛүx��C:�hZܵja�v�"�V�j���F'x޴֛�
Y�F�po%x>��^|{;�ԏ
VDBĉ��!��-K4 �2���JK$��nY�'�T[4�ݪ��yh�c<@G<B�p����G�4�1���Iۅ���x�D��Ggul,T��C����.PR�a=��}pR�y�
�X�"~��d�(�WpQq3����e��@�v�<��y̓Q�i�&x.Q���"t��2P&^��+��Ƀ�W�,�ƭ�y��dy:9̮^Up�+�A"�����2�<�51/��,,�ZL��q
�8����x�PbAv�P�?��Z�hfY�(@";�,st�����B�54x\z��OUcH�-�wT��|Ⱥ_�a����0�D�w�2;��:�x�=��ʰ��}�*���I(�,c�&iR>��� b��s�|v��0=�5T�܂�\4��'��l��
Z\m���!Œ��F����e��z)���{
2����J�X��UTy|��� A�@~�B���"؋%�K��U�� 	v0$��U\�j!��h�������#�l`�<j`[���ă�����ޓwr��0�'�滪x_�<z�H-��.�w �`�V�
�E������#[5�aN3�f�6:���"f���Weȵg3�D%�7Bgy�Z����9�9�T�Ckh��7q�x�CP|�R��#��j�L����*.�[Ƥ,5��lT���W�ѐ&>�d���͘�>?^}q/���3����g2W��t���g���C����F��P�D�(�4�*�t��ly%��������w�y�`9F��L�/,�Pl�<
�H��<����Ì�e�����xB�>=
�>�L���?N#�3�j]��(�V� ΄�H�3�/�QCż`tv:ޙ�vz]�8������|$/�k��Ufl'_k���P!��C=5h�̣w�ʶ��4h�$�(�t ��2B|�� �n��j�+8���)i�\8U�Զ�e�N�q?�[��^�g�K�Z������}�D`�	�"/��bQ��k��Pʢ6�����`oU�gd�˂���C؟C�?߲�.<e����p>Nt����&pN��.�}[���{�}���ă�e�}V�~ݟ�9�p퐀z|u��z��,�2���>Y0� ��6��ќ������o��m�=�0��h��.�-f��h�������3�P	���*^�D`�����~v�ͩ�T�J�Tj�3RN�;j�,�$pʟ�}�{�T�����(`љ�b�����
���']>���օ���[h5�Hg�\6'U�t����:��NN�F�����=,g�W*��BP��L}wJ��S��m�Gc`�w�8&�n:����u�։P��(���/%��pl�/��)�?;�Wj�-LE�n��4{&�r[Y�Ӟu�tpld��p�[�\��O�.+�1z�j�8�g/��V�|��h�a�i'p1�������p�H�3�������	n$��|���=͢1�}�M�]��x��-6��U�4��'�GV�!RݩA!� ��Mꞗh�c�P9�CZHBˇ�$�
^b� hu>�S+��������J�T]�����	�oc%��ȴ�����E:�8[�n��t8�1j�*4���R�6�TOB¦�uf��R3� [�ΞX-6"���k��Bږb��NF�,�i�MO���Ao�c�N�����������N�=�����0����V��o����Mq� ��3�{ϒv�jv�~Ѓ��C�㟪�<n�r��w�G����͹��W�M.@d� +bU�z���/�^�Z��3������R/pFTr�zN%����%�EФ��N�^�憓�������ww�F0c&��t|��hE^}-l��ƭ?˚<�;�:g�Ri��Mݿ�珐c����h��pP�Hˬ�J��h��8\��oڨ�k&$�D�M0���󖦢O����7�\���P%M6!{ki/诅9�1A��*4��ls��_�S�;�����]Hj~� X��"�>����q�[���w����.Xi�x�{jh'�l���4v7(��i�'AV*M];���m���a��D� _7�=�b^�� �uH�쇑�E1<��b�I��zXO`����n�)O0��h�E����Π��T,wdz�����D!5E�@Ĳ	E¤�o�ṧס��� �5:�e��%ΨЉ���})�bn!-�10��O�7��FҶ%�<V{]���)F�+���9N<o�<�����W�ǜ�����H�ĳ������zft�Џ��.k۪�|�]Z������l䆣���ì���SZ�p��0�~�Qk�'5_�3�� X ��`��p��tT=r|j��y��Z[/����0���
��Àۛ]�Ê5�,��`��AX6^����&�`�}+_��a��VY�9�y��t��n�p��A�8��BL��jJt�Sb��	��÷��A�sT�$©̜�{�X��ZU���'�Hܸ�QJ6�1Ξ��2pl�H_	}Y.�&nl���-O�F��y�������$3�"tAh:�ɪ|��}o��K�+��P�X��0Msw2����:�����Q��l�����fhڻۀ$7�ׇ��gD!x��յ|?�Q�7m�W���^u�{ڪ��@T\��G��#�4nr��0���J�
8[��B�Yj�vh|�2�I~��@�wγ�~rqu��Y,�/c�t�"��_%�)FښE(F���{ҋ>g�i�,�J0���L�J��)���2o�t:ϕ���1(��@��x�6lV�L�؎]��r��0�i����D�L�ͩ�K*]�|�j5��t�i��1½�07��&d�3�"u��ವ#���Ժ�'�mc-�	���v�b�ҽ@.�ђ�ɶfc����\��!��b$an��?�������m��|
������ܥ ��HI�
d�;cʸTv�����\��E֬>�j���]nv֠����Ç/;$����Нf��<���d�A�=~;�j��!��wY\�`mZ��r�A�#?ݧ�,Z��ߖ�
�W����huI�j�#Q����^ȏ�F"Nz�l��řEa��o�j�>u�r|�aU�*�;V?�3�T��_�&4.�2��J&�h������{[/$���h���@bjBdb��ӷ�oՁ�(��ּ\�>�.xτ~�'$G�?�P8�T���.KT�a���}����}$
S�="YD4d7{6W��3�o/��j@jn�W�A����^s�iU�x�U+����ufQP������h���2��,*/Ȅn_܏9'q`U+�e�\��~����<ͨ�/\���Y\Z���,���Sby�X��r�AC��Pr�H�U��f�#y(�E�G��W�m�Np��\���zJ��a-�&��	������d�k���!k�r{�2��z���b�Xi��+@�}�N�9C�(#�ͦ!�>��  L�s�ب�O��#ܽ0�4������\�E����h��*,��!*����]��k
������eBX��:�U/���6�� �v�~��OJ��F�FK	��O��v��!�/����T���ݘ�l{��j�k`�t5�ľ�(�~��r���:���7Gxz�hz���-��#�<X�؜h�V�'��{ �x��#v�W��NY%�q&Z�GN�f��|��+�"�&D@r�B�e�Z�{Üt�����k�Ⱥ�b�x�`FP��LR;�_��-�JN�e S.��@��H�������WgT�&�d��ԼhM�>:�mqiv���f�FoJ��22vRt2�gh�LC�㒡)Pm�(��m*����G5y`a�66f����f�`��gv)/fO�+?!<E�Ҕ�2g~0�I(I�eN��������
��sL��d?��.$j��
(_�� �{��l�
E�Q~	`B@ޔ/�v�{R8>����d�s��F�-��uld���p!�;e=��̾�d�1�~��$�t�r(��"B�
H Y���oڒ܍��1)��`8��e���NLF�恃y�����i�J�8�&D�?�����������آ�}e���O����G��}J����Z��ZӉ�j�=e�@��x�ٛ��� &�n�����[z���Ԇ��UľD�<6۞y��є��K7�|�)�z9��H��y�Ǜ�%�1���,�d$���
S�J
.=�\��G��f��Z�Q,��Kb3��u�.m#^�v�L@��evݿ��s���v�T�?�R���j���_-۟<�{�L��c�׈v``�ӛb2��f�d�E\����>�Q����-���cP	�gnV�6-t�x����RNIu*�Z'N��5
,��5*a�~B+Y��M*pw�|JS�<���۝`���8A�|:"[��P�O���?�ï#�S#�w'�p'�F���?�2mE��L����.�_&�a�YI��u��������\\C�rO��+}�z�c�8����|V���CHla�s�p��_����6H�セ�`��7��$&�|���81@�2Mc��ܓ��ڨ��h�v4A��'ODQ�zR8$��V�����|�>��9/o�H�]����^��3 #�%�n���]$�⸦�ӀT��1ּ?�	?@%=k洨ۘ�X�=��7G����8�,�C*�������o���!�)uA�;�� �yB�Sd6lH����k3@�ǽi9�=�Kԉ�J,i�خHag�E�(�2��[�0F�ƋF�T����Ü�b,�G�ܘ���1��ML$��<���)v��#�,�>.>C �؟%�n�OլG��1a���T^��Ld�Պb�>oz�r��jn9��D<�����T� ����pa��rI>k%_��`?��?4�N�g������6�g�w���FAb�4�b)�^xo�k9$����<��:��|RD-O�������Sc�N²�5�pә�H�-Ji�n�yl��ۨp$&�-���'�z���	O�"~Y\ۑ��&�6��i�����p
L�=hMz*T�l��B_c�g;��V�:�H%i� s�i"�� ՜�qTs����'�rg��w��X$J�˖�c'�����gh4���|�ȽA��]�������?}��~eD��7L�D�w�b�~� '��A����ǘTI���X�x���A�nN�0�*Σ��h��q�{͆�(�d�i�{���5 ��������ڼE��u=����~�:@g���\Ф�6��p����)!h�S03Q��2#�F-���\{x��פ�٦���tk�<�3 �7V��&�|���&���@��O  �5�����GG�J�I�1�8��]5U���U�ކ��(qw�Q?�Su2��<�~�43�bs#_9̖���U9D�+��tou�r�ΐ���̕���6@ɛ+j��e�ڨ�p����c���Y5xehћ7l��3�^[h�����+z��!�V4f�X�l�=BnǊ���I�M�~L�8J�z�b}2���-Η?�hsO~~�Q3�6'X�EZ�~b�a��A�j�=n�6����l5��\���_���.��lV2���֞F�[�y��3�w��$1J"��:xY|94�oP�K{q���X��
0h;�2(T��▁�Gj��N��+��
�h�[ۛג74����gD\霉�Fw�QB��m�v�����;�{�T�O�GiK%#���rZZf0BQ�-�_
��ӽp~%Y�o�hm?杻�~���@�TS����l��4�j%�tR,��Zb%)���E�t�s���g���,�K� ���T�J������|���ǻ���	1c�:@�ay�1?/VQ���ݧ1��]������L#r�F�.��%>o��<�)G�fk%����.�.u"�#�mIC����_�:m>kb	)���j���L.%�%���Oc
��s���
 ̝�$��&�:��v�Q�ng{�^͂>����������}�z���lָ�-��f���CE�����J�,�nqkD37�~G�;?@U�Ck�f}�f�����i�~6Q0������\��Zf�r֨��^oG�d
��
N�em����h�־jWT,�R����*3nFD��j!����^|So�t>P��|�V���eV:���l4i��46�H2�c�J0���ۊ]a�[*��<��hk1�@}�;B�s,������1���o1�鶙�Ex��|��`�G��%+$�T'U��S�.Fvua�G�}|iӡ+
·)"4۔dr�W���3�\H��8@%��r�Lo�Z�9��i��xdz��rg���P��� ��$���,e����'Z_�9�S�U����w�E���nB�<<�/�ł���Z��[,�n2��,��̵�A~�ZP��P�Xf\�(��w�b�=�����;��f�\���u�Z�-X�c�$�ǺUyFұ�O�_�P]��m*2��J�s�tʦ�}g�!tK(�Y��=%>V: �0hs�TC�����,���74��q���!鷲1�,_���)��v�����K�$߰���{�
�dȂ�m���e�NБU
��qg� w^&~��{�P1��K$:L�ʡ�v���N
�Ŕ��^6E�S%�l��,j��Q�Oо����N8�m49���D�\�gx���z�V�-�?��wY��7��V�cT��6�3��#�I�fbN�I���2�����f��=�̵�vED[[�B]r�Z�������?k��1��sTx>�lP��:R� h@ᡅp � ��.�u��Z���m�a�srW���&�ۛd��"�>5�q���o�#(�Š26tm rg7�C�:����P(�1(�>�*v�)�"}7y�D������ў��@`���ӂ�H/��^�2!<�є,H/y��I�1�e	�c��.��4�h
xZ�L3U?�?)�j��(4� �>�ѵ��Q�m+`�-~ޏ��v0��8��j�4��2�!�r�Yl]���#�!J�f=�q2�ٯeʬV��ꅊ$�T������B2�� 1<�8��� ��
a)߃y8������N��lK�����g�AYW�D�'�s~�D��,�%;��tU��
��,��e-U�օt�I��x�Y�S�oT�u����+e��y�t	ˎ��&&���?�[)=�q8�o����^�x�t����L;��|��z�x���Դ���6�r�,;�򇩴��ӈ��~����=^�:�B׆�d�Ff�������O3�8J��t�^�|������v�֩ΰl����T��RD.<jsP���
 ��f�{�d�ʾ
̈1�`.�b���A����DQ�]�^>�4��;$��pW�kN�g�>D6�$�tl_�pI�ND#ꁵ���Nm,�'�*��
B����(�w�B�S�����s�`K��8\�:��h�+Y���r�^�˗=���*p���?1�� �sL��n��K|&�pY��BuLȋ���|ڮ���\~��O1x+x�rzD}�8m�I�X����;a��pgi>��A��q�wH\���'X�DT�j��$a6�|*\��3�-1�<�M�2ܮ_v�#��C�4|�'ꋧL,�R��z�<\�)��\��9j��Hx'�˒^�& �6q��m�د�������T�Xַ�	�0+%�f���Nz���M��B���)��'� *�����x9���zu%��� �m�N�E6ǎ9�g�kN�\�8���d���, �C�����ٻ���?���g��2��2��s���_IIT�g��7����M'b7�-���Yv��~������C	w��OOn{L���q}�܆׬�P��É<d˲bKוz\���h�DO?��Z گ��DĲp|�Er�!t%:c����p�کsNΐr�<���7Y�2Uw��F�>.�H���	�^s���Ƭ!��hN<2� ::�R�<��EQ�Oc�'���p�2HϬJ�Z��T�����&�s���5�l�̞�O���Y�\l紆H6ri將���tg�㧃*��2l�f_�Ln;�/���H�sB �I�"'��wHq�cA�D�R�mR8���|X�ߕ˱�&'����g34�*�%��s�A�G]��=���꺸��)4D37�i���b| :���"���;����I��X����ɍ8n���0�a�������S�V���Dd�7t�v�t;�5�[~���.�ڗ�NMЦ��U��`	:����G�п���s�d����!�j0�ʐ�-�3F�/�K�g{�^6�T����䯨�<Q��2���q�)�nT�5Qǚ�#;�z���H���b��
�r*��ۺ�d�P����]�O�8r<¯���1o>���cS�¯��7�~t7k���[�^���ɰ1(��%t��rr�Êe�s��d��к�&���r�w�W�H����T5S���֫��w/�^ʁ�]e��ּ+�`h�W�kVjÔ�W�쪣?n�ĭ��e;�H�L�QmJj:�bX���ؗ���sJ�T�_�ɀ�L�X�DZK�X��>�|R�ت�6����T<l��rm���_�.�(l�ҳ�c~hF���yF��2>�$L�"jb�:S	�|t��o���Kv���sXs[w0�#�2�?���<��*���A̻ ��S[�h�q~۶�!7�$N]��D��y�$��rZQ�rmd������q��V�T��G��#��Yr� s0��\H|/
���KڃY�F�h�+��M�~ZZW@dQ��ӆg������t�U��U�%)���E�5 �-��ҁ���`��,8z%����|}Jl"�����juT��+�1�Ĵ@+a2�,2Vi�HN�܋��F�&��ʬ����L���A��cWB�f���K���lI�sY��3V�M���)�"+���(���� ��$�mɳ	d$����Eu.�XX�?�c%�T��l������0�$��ߦ5N�ѓ��)1M�/_؂��m��af�?��~+	�u�%��¸�����R��RW]E�J��1�}�4�nl ���x�9';Z=��%�fX栤�\G�wVm~1ё�H ��{,�\�ĢZ��r�]`���姷�r��U���ѐt�}h��ojҤ�H�lC����FZ�����;{���@o��U>+��|,��`-�V5���4ͥ��j4Q�2J�J��}�M���[%\i���yh&�@@�&�BZ����Y���>�^s�̊���=xE�>�۹�Gv�0�Tb�.�Q�D.A�VaN�}7S��
IO�"��d�WA~3�i݂v�o@�������S��i��x�����JK�+��PWFG�(^�����t,�_��J��Uo9�U$U�4���Q∯�I�<C�>/����%Z]ݬ�4���"S�1��*A�PdP�p��K1�fj�k(q�[�}���MWz��I��/}\K�]�p��tr\-��?o���Ҍ���3��a�h��2L/t�kăȎ�6�!Ʌ}B���(Y ��ט>�� �5*s��E�E/��� F�3�4T�J��;!����˔�V(� Ἢ�^���x�K�j�䫵
C1P�=ࠛ�Ʌ�U�G{�g� f-~��c �ؼ��K?�s�E��v��v���eb���Z���"�Vql� �jx�.�*�E�4�p��+Y�h�u�A{��x���zy�k-���ɲz���پVǿ#�Vְ�#�/(MH%N�Z���^��}��f��:�hn��H(DvdB؞lZ��:����%��k����H��x��vP͒�R1�C�������.�2Ƶ�X�(��� R�W]�&��dMS����>0�"qeJ�*,�C�8@��2��It�x�g���C����WGP���(��*�����y֧/�l�	��Ȟ�`j�ӝ�P/u�Z��D�<��C��}�t�XI�9JeĘ�����!
S�Ln�-?��$lHjn�:(��# ���c����Q���`E9�ފv��8��}�"��\�����1�l�b_�m�!�.H=f&E�����'&8��Dw$<��������B�Su �p��S�ڈȍ�t�))�8&UP����N��\�����߼�W��4�.RD1^��З�s�fm9��L���X�@��A��8l��s������O󰐣��`�e^��H���ꎊ$�&���_�![D ,��K��J�u�4ǹr-�o�G�J���#|ƥhz/
�é"�����T��'���_!��׈�\�@��=9��}������f�"T����[�3�܆�$�Y^})r��A����v�y��)���{�T�=�R��jN��9�r/{��B���0r`"��b(X�f���L����s>�7{֖��+'���gdGj6�<�tX)�ēN?�"�=�4,�w�*W�B� ��F�w(�S�N̢X,;`c*8w�:xN���(:��0d��s�-�-p�?a�2<^?�����L����d�&��kY���u�?����|G�\���O�B�+s��z���8(6��T������aO�Rp�������=�H�Z������E��$���|�XX�.�1��UM�m��1�ڞi�D�4�s'���G�aR�xwRB��8�2�Y	��	9�%1H�:�� ^smy �� ����S[޾�Ύ�IM�T.Pvֲ�	�@�%������c�N�i��L��� �E���">�*E��1��i��J�u���x ,�ҞIR�6"�p�"E	ki�ǳbܖ��M����,����>�)���;��x����9����|�����`�wP�|V���e��wܚ'�M�Z�hw��Lm v�·�l�д��C63���ZnVi���?���_��
c��~�d �bƏ�z7�Լ����y���`�
 a���
p���r?%i%�b�ֻ��u?1N����lx�N���w�F�\����_ܘ
�^n	ɑ!@��pg�<M^P:���R��ڔ�)���r�c��ǲy��pI��H��J_?^�/4��L�X���Y&0�^����� ��JO��44�\Qf��!��6z�i@�s�j����:^"*��wl$l�_��;�O���T�H��� ���"����R��q�s���5�h]~�-d�X�����Q�'������N4')�����I�Ag�U]l���P��5v��rDR3K7����Rboߊ �xp�=����q�}dIPcX 
�����n��0L�����&�
E��1����dK���q�'�5v=����A��r����s��b}:���V�q�ژ���_���fp!�_t0id�(�F���v{�M$ך&���/���<���-f���4���P�P+T��@c�U��Ű6�k���C��`�����Z7�.V�]�$��s�w��Y����+-��PLS�r��2�~OZ��O��L���Z�J�塮t���r��@����\�l�ě!�K���2���,��v?|5.7��@��K�^Y��������+����*�V�@�����E*�n���R����L�
J��b3�g�Ybחu��sE��º�`���X�oZƳ�y5��ĸs*6���ί+ÐcM���_z}�.�5�l̒���E�F���y����$g*�"�"�:.ٳ|���o�	�Kq]�a<X.LH0�+�2K��˷Ɂe����i�QN���Rh=�%�ѝ�7*{�8�Dһ�����m3<Q���m��Ә���^�1��TG�0#��)r�?0�T�cEG
~���&V�Y>�hM
a��~�K�@n	��:⻊��@��	9t����P<�)WϾEYݏ�H�p��e�;�,s��i4��ĸJ�i�JN�/q���B�����1��b@ƀ��'E�V�C�	h�r$�ש�������LY��<df������ū���7�N,l�ak�覬�$�8"��2����G#�U�m�F�	�H5GeÖù�.�K+��rc@۱�if�h<V�u�$2qЦ0CX�,�5���J�+�45%�i5�V�F�b�pȐ�Lߎ��t���^�����Eg��l���O-ng�`�����&s;u��9 Ff3�9���c�~,q����R�6��\צ9Z\-�r�28��/��R3��������/�3h�P�jMl��ùB�3�`ؕF��� �f�����Vo=">�N|g����z�V0�k�"U����4l�2�PJ����Z�q���[ (Ъ�4�h�~�@��B��$�dژ� J������!��O��x ����27G��[�T��%��P.<�a�j�}��p	Jr
�6E"�h&d�1mW�w�3����o�@���"�e#����i�x�#���Bˎ��mP)��CT�� ��,�'P��|�P��98x�U\����%�xn�$�w<~��/-9�SZ�*�]-��2���2�����A�.�PC�F�9f�,�(,qě��'�ȵƮwN!�\���k���-���ZUg�K���g��(w�41�c�N2���&^�ȩ|@ʜ��}z����(���h>� NZ�s�����n���OP�n��4�6������m�	Hl<�����k��8`������[ջ��w
��\��?v���x�D[U�̅��6 ���~��[%@�w|�KZc��¼v�#:��B �J��@#�a`�ɦcl̈�j�M��f<�o�B�O)r�cv��Kb��j5x�z��:-k+d����mB�V�;�1��o�#�m/�IN����"�]�iMf�7t��>еS:�D���BS�Z`���%G���4�k�����<x�veP�NR�/�.���6��.���^�����;QNW؛&��d��u�9+h>+>�qz���^����W2ì�t��g90C� *��OP���(�u*l����l�y+������w�V`%)�ӸV@/�PB��wq<�*�bӧo�I9bne�1�2eP�*��
.��L�gp?�eR@�j�LC(��6 :C4p ��Q/�j`�d�ޅ�xv��8oU�=����+mlR�l��`���! �	=!�;�h�ʢ7�#T$wCRC�o��F^B�' ���n;��U�f��)U��8������kN]��F��'�7D���q���5D�50�������Ⱔ�D��"����P�L��Ӯ<�n��C�؋P���������e9��ˣ�D����&܏��7[_#G�g�"�%^�o�� ��jͷѥ���|N|��z��R�����*���lص�"	h�=6N������5�����=��ٸł蚅�f��Z�b���|��3��+���^X`X����UP�v�ϩ���6=T��%R:3mj)�M�%���{���t���s1`=B�b�5\���t���A>�Z���������8�g�o\6�t�t��G̦^xN:���kώ���_,��@*ҍ�B�����w�-S�䢳J`�F8�x�:�6@���<q����(�Ʈ���pX�d�M��?'���yL1#?���]&��YZ��u���rcW+\�AOg�@+n�Hz�I8���p��:�Ԕ�a�R�p��c���b�'��HҲ̻8w�1� 1V$� �|`u��)�(1Q{M����#��L���(64��t' {�B�RIS�h��S��ف���9��H��&�7�^�r, Tx4������&��s	����Tɭ�֭�	Pq�%n�X���U��ߑʤ2�2����c��*�fv�>�������u�&I>$e Ǵ�D�N6}{h�ݖ�k�{��. ����:cp,:$��9W�VG��OU5�Ŋ���W� ���ש�^��%����x͇�5ֻ��H�M�e��DR���v��4t��o��CQ}���Jn1�@����p���2�e�_�9eId;[bAhGz�n����z�͋�v}�e]����p���r�HJ%�hh��l���N�BO���q�	?*&)Gwq#F��v�����3+�^i= �|���+��<hT�:	�\RՇ(�9.��S��c�뤲�p'p7�H7q�J�CH�
�%���ըA�x&�����������O~Gs\������6ii��_�%PV�]ټ:*���l_��_4�C;ݯ��K�HV�n �m�"���-]q���z-��c������XUk����'�޸��ǹ4bd|�MJC�?&A�?�]'["���R갏5s�!D�y�7���Z	bʿ �d��XT��1�F�X��I�h�X���ֿ�n_�:0/�����V��0l@�{d��1�lg��]�51?��.9���M�6�~�`
��M:Q+��A����T�if����!�r0��#�F>(��ۉ{�\��ݦ�De�%��<�A¾(��'��C�q�k%��x~7�0�a� 9�b�� �o��M�{���?檩�']Ƽ���xU�ۆ�-�%9��	�S�B����n~*�+��(0
�����f�p�\�wt�F[rh�M�qA�F@�R����v����|}�Gtg���5	Й�L��୆^i�bĸLP�+�b�M�V�э�	�����Bn�������~�L*J`�b����,ʗ��s@�t����guX��PZA��T�ݩ�܎��O6���
;:�H��T9_�[.hz�ls{ę-$F��#y�&j��)�$�gP"`�:	�|ꕴo!\Kl���ydX�\}0�Sc2�vG�R���l�w'��٦	\Lh��Q��W7��D/�D�W�Z��ho:QSe]m�2���g )��TH�G:�	#��5rk��0s�~.�
����YVU�h�v���~]@ڪ:�	e]��Ň�,�t#	 �Kٚ)��E�#�cP}�w��q,�?[>q��,�J"�z�^�Jm�`0��dE�1E@a�̾"x�V���El�.����)�0X�L����7b��-V۬�+#��S�)������_�pN"�|��ĺ��M�С}m��	ڡ�����M.6_����c[17���C���N�C$�\��+��ه�G��$=�e�Ƃ��(�D)vܑ��ϴ�)�k�W��H;�@	.���)�H��EBh<᧓��j�nb�CU��ȯF�;�%����@fZE�tGz����~'1)��^$��a�\�xZ�rrg'@������k��K��v�J��.h�=)jȥ��g��}�x���mF��{J����{To��>�2#|�:Ԗ�V+�ˉ}��Kh�4�z�2wJJ��ӌ���.�
[S�M��h�Ux@�b�BPh��?{%�[̠��1�����Jx�K���Glq~��1T�J��3.7�-a,�}��r$α
?>u"�_Wd#�Ww�23�{�,\�@V�Ñ��u���:iA��x5�H�}Z��P�+'�^��T��P�,;��l�K�>9���U0���;��~`����9<���/�uX�Q^Z�FJ�b��wf�]>5A/-�P��>�A�f �^(�������C4�Ɖł\"e\��C�fc6*��-�!ʼu[��u��B�1W<�!�8�^�I2�m�����m���Y}�i% �(��k�>g&\ 	�Zs���;��|�Jܩ(4��e��e����<��*Ž� ��2=��/]߁8ػ�k�
��ȳ�0��J~��P�U�q��"�� H�c~�)h����2bKu��;hvwsM������q��F �o&�݄�l��jn٭��`�Ī(���F��^G���;1��f�x�izoz-Fљ�(���V���),�d�*#��^Ck/Nz��]��\�f����L:D��hB�WZ;��`���[��k�!���g�xo8P�tR'��ԛ�6��ц�.���k�����Vp�WS��&�q&d�M~��_�>&Hq����q�y��6)�2��t��gԵ�C~�d��PY9�((�*�.�ݳ�yL�N����`K����`����6/k4����<1Ʉ��HXj�I��e: _�M0(��
	��L� G?UF 4 j$��(Kp� U����	�v(QjZ�`{��ހk(vA5p8*��X���Ťֲ"�!�l.���a�![��=���*���%��{"!$����w�jBC� EP�؉���~��A�O)��;8\N��|ŎN�Ρ|QU���߲�\��(��$�MDg-F�	���)P�xl��࢝|���F����n��ib�j�<�Fq]���E�V~e,���E���&70����x[zFj��8�� ^�Ī�+�XߞeD� O��7R|���z%�ʒy�V�e���|�� �,;�Pk*�/��6�q=�K~���>�5�f�ƽ����7�H3�8�K@^3�.�8I���ɲvɳ���5��/T��R��Wj���Kb矨��{�l���i�b�`X��b3�ҟޱ1���.l�>���L�������'gZ�6n�Vt���A5N5�Q�Ɯd��X�,�w�*M!8B��v�9��wQS6S������`|J�8��:>�Չwڄ�/2�#5���p=�h�h?�}�5Ll�5���"&�]�Y��u}���mO���2/�\/��O�(+i>zU��8�_ 
�f��ůCJa�܉p8~�������f<H��B�=t�����8$��|����$�1�J�MO���57ڔ����-�4-�'�"�=�8R�M1ȭ��n���zƝ��j9\�HI�����^)�? I���s
�IP�Nd7����Td+�֨Cz	���%)��hO�D��8�3���{����*����������-su�׭y�_ bC�?�-6�! ���k�$4ǩۯ��Y��u:%,���4�\���
R��1�����U�2�I�@y �D���qZ�x�3U�PU#��M����1��vwv{����(�*��Cl�A��un�3�Np���%(�����6dVj�b�`�z��X�V��/Y��4v���!�u��p��r5�%���L��ЫʔN�˷�M�����AT�w��MFw�������k�^d�����ڭ��*<�jh:�f�R��&�tRr�c�
��/odp� |HRr6JUh~��{ ��'�ܜ�&�l��C�fM5��O��+�с\ǺE�Wm76Ği�ML��/��4XTw�*{�1l���_ϲ;�/`��3KHT; �/�"}�_��/q@� ��$�^�>��SXa@��!'y/J�d'u4�����V�U�A�]�۪��`��++�N�@D���7���;�b%�( kp��s�R��q'�3��I��7XVֺ1�n�0�ŷ�� �-���{Y�d����g��L�+5�`��9�����(�b�3��h���y:�������/��Έ�f�w!Tde0�����_F�Ԍ|�{䋘א+��r���` �<"�(�#������V���?f��۷����;�����h�;�z�6dV��D]�$�]�tE��+��5���u�fc�=�IS�2[�(��~ ��N��ˏ���4������Vgt�!7r����~�́	
��B �������k�b:�l2O5�
ч�R�H�^��6�nL��G+��ȳ�V�5��D���{�Hn�2ա�P�9�YL8�}J�8�b��������s;R��p���"��Xz�Z�h�/�ũ-�m�� 6z�:�ejѐ�bx��Y_pȉ.CߧlBs-�45F��VyW���cσ$���"��:�؟|%�o��}Kg�.���X��0ԛ"2�������U���Ra�d�h�D���7 ���DHޤ�� {c�TQ�@�m�y"�	�V�����T�@~G�Y#��}rƳ0.���7O
t֯�ܭY��lh�'����~k�D@�P�$&؊�ޠ�sVn{t��#�F�)h�Eό��~/������U,��2F�ִJ}X_���e���='�?�1Om[@�����Vz��C�I�7�h&�[���k�rL���2�t�����˕�
���22W���
�Y`"<�P�Y��:=��K�m��	}�|���.����p�]cv��_�p��l̉]�$hhZ�&!!��N�ZN[��"��*x�=��̌��O/��f<{��Ǹ��K�����e2E'T��-���n]���D=�j�_;�\%�/�f�ï���1�Hܩ~"_�Y>ͬ,�\�_ZR��rB<x�Jp������������琥\lh�J2jCV��'u��=Ȗ�F	\g��6��l���s:o�>��g|� ��1v�V&�'������/4�]2���Jm�V��`�Ƀ�[ �+hWL
@�0�B����<b��⠠/>���s�$xv��,��G�M4��T2��"ί.2>#a_`}h�X?rY
�e"�vxd^� W��3zP���h@%+� �[�ͥ�Yi|��x�L��x���<;�P�N��y(L�Z��y��,QZ�|�F�@9�+U�݅��&��h����K<��A/c�O�EZn%��~�ڲ���6�8�AjK:Py�h�<�
f{}�(��!���1���g�d3G�K�\��aǷ���-Dp4�����A_!����p���x�Y&�2]����s��~,ʒ6}���`??(*4�e>�_� ��s+��϶M��W5��c`4%:���*�#���+*�E�T���s�hL*�7���5s����
T��n��,�:f)Uv6+�](� �<�~܄�zO��g�K�n���c�vR㰴:�V6zp��l�����?�tl��j�O��{z��C�����Y8�RL��H�x%�z�p�-!�_�c�IأsbV��:�gdǰ�-#�I���vNUM1�����Np�f�%��y�Ե�}iD�?~BI��Z���UY��Yk�sr�Y��x*��P/R���ԛ�q9��lp&.�)~�ƶ}�Y;��q�JW���&`�td����o�4>!�Dq0���[D���S��X2yƥtYA�gou�CyF[�h�P�V(C�c*b�Wݎ�)y��\�=����֞-	�`����6�/�7��r=�<l�S��� e]�I�7e���h� 4�
�vL��?�F�H�jS4(oH p��*��Q��Q�>z`��{Jv���8�P�sx'�֍��0lɆl�w!��-=���E�{ʘTy�VA�$� y���B�0:  �	ؤI���)E�r�)�ؤ8��$�wNNI7|� I�-�a���|�_��DE������A.l�*�֢�@�����2��	���d8��M���(��Ky��se����u���{��&��萮j[����]�=�������BC�ܞ`���[:R��|Њz�~n�T�xԠ�Ǣ?٣W���B�Mz�&H����@=�5�.4���f��|�3P��A�32�����U^.��s�$�c�vĀ��:��ŬIT�OR0��j�ଆ�\�C��{���*�݈Y`s��b�P��l5�l%����>� 	֧mc�\�Jעyg� �6ID.t	y�����N0��!���n��,	(&*��tBr�I�ta�w�]S���i�`7nt8Ȏ<:�H헍��c�����翮>8�p��W�n*?bo��@L�+�5�&��Y��u8���Vhl�S�\j`�O�vi+dm�z�"b8Y$0%	o���Ŋ�a �p�oi��!��*~HH2��8�8m.@��+$MK|�����1:�M
�Y�hr�I�R�4hT�'V�	8X>R�g��E��!�:ם���9V'�H���#�^�ݲ �9���{d���)�3��o9T�ȡ֣�T	2�%�9�/[Q��l�Z^n�S����2*V}w������E�su����� �{Ϟ:�H63��S�k���$ȋ����԰1�,p���/� �
���n�LP�w(�c�{{>������8��/�����k���-�M��%�?��+vv:v��w����C�q���Ņn�#�n(����8�Z�կ�fdq�#b7y)z������k������K�x��0'kp�f
r���%������8�F�:N�t�e��\�Yw���FRv��4�w�i̯^_#�2�X��#g<��0:�_�R��Ԕ��凉umc�I���apz�Hm��JЬ ��O��jL�wӾ&�"�o��!�8#Ot|�P�\���56�PiQ�8��/H�+3�Q"*V�l�;�_j�y;�Ϩ�ӧH��+ ��"�����2q{d~���/�Y>��>cX�v�Y'����?��4�:���@���Ax
�]�|��l��x)�DfL7S/��<kb�� &�=��z+�'x��xIk�X��rֵ�Vnq0}|�
q�{ي������d��buJ�*n5��*�T d�m��^9��D]��(:N,���?�+eq�_��A��!�L0:�ĻF��n7k�{���^�M(���<��&��}�ݺ�9��y�nY����v�_�<�)��+]������g��i���O�]|L��$�"��g��)�۳���^S�B����~�������f5Җ⍒�S�����t�r^g�ѬO̼�=Sr�޳�,��cz3�} ݂���5�a+�¼���]K^��@��ޓ��c�+劇C��V{����9�~�n���c�½�LS�SJVxMb��6�
!��FK�s6ׅ���%��KhX2!�Z7�
c��h�`�D�b6u1H�������Y"_�d.d�l}���\�F��Ey��Ε��$�A="V$o:��|`��oWa�Kb���r��X_�0��2�-��\�ށ�����妿ܿhn 5�"7�7�>l��D����i�^G�Q	<�mP���$���]q���T���Gp-e#��r!�&0�ɋ�`?
�"����Y���hf���>~��S@P�I�?OS")�{u2��
tY<��As )h��E��Wԙ./�m���̴�,$���G���\J��c{�m���\�Vkp��R1��@��G�>�V�Z�:a�d�m���6���>cL*m�-�,ό��I¬�𪅺���d=��c��G��bn"�����U躺ƞ�m���	P��G����/.��d�+O{c�=������v ���$��!���=ͬ��=���Ղ����p��<��Ū�a���]{4���M�2C:�>U�E�\�����5nX4~�%��;Ƴ-��O�f�M*�����H�~1��=(�g'\(�Z�]Zrqഅ@h�#ZE�����,Ő`��hxj�&�sF����1@�F���1�0�'���o�/>�(|�*��#�V!I��3v^��_$4�`�2�#�JH�i�R#d�b[L���;hc@@�BF����O���)���J��,�`��x1o��G^�GbJ6r��TN9����.- ua��}#	#Z6i
5�"{��d�9W�$/3u�
��K@��G��}�z�̀޵i��hxkh�s�󎗒�PC��Ô�^J8.�TJ�,�@�����A��9I��U��X��%S�t�A���</��/���Z�����R��"��m-f�� A��PǊ�7Umf�UR(]���P��9�$�?��Ҕ�\����\KU��-��B��ǃ��h���ٍ���Wg��Tu�2�(h�W������[^}������(�z�� >�J �sF�a�1팞2��Ό4��`����~�y;��`�s��s�C�'�r��߷Q��Ыg
�.B�)������=UQ�񘨀 ~�z~��\lT7ب��K�K�1�"v-sd�u�|�lG�����%Z��X�l��jdP݂���� 5r� ⍓TIA�|O���x�ze��-�|�ɞ?\�><�V�oz�¿��c�#�59�N0���O��飺f�̈��qw���\D���BĐ�Z���ŏ��;k�娺���x嬉P9��R����s���ڰz.�f��!�߈�K���WI.&;u�d9�˼
)>��q��q�7��"�,$�2Tzt�4g
U�Ct��P�P�
(^�*ݿ��i��y�t���r�|>��fH`V���	W�/a[��Mв<����3��`�MIJ��e�'F�&��~
�O�LZ�?�g�|(j�(��G ��s�<a�,�]Q�B`����vI<v���8��s��Y�����h�� 8ld}v�տ!��=R9y�`l�����1��$(2u����B�d� ���ؿ ��t�1��[?)�!8��F�re�Nnm�Ɨ��eߨ���2J�/D�|����c��D����E�����к�,#��m�6%�_.� ؼX��Ô�L�e��Y4>�{�vh�&����K��[��ȷإ݆�iw� L��)�[�ѶE���|2�z�>�/�J��>"�=#?���NyU��N��A���,U\=���i�3�k�f���s�����;3M���z�^�ī����&�v�mg��.*�g$gT'�0R���j�YA��<��݂{ϼ�ʅ_r���G`�Ёb�5�Y����>�dk�>����P�����gP��6$�UtD��w�6N+i��|�0�)�:,$�t*C��BM
�����w��|S����Mw`��8�I{:2^�r{��� �e���f���zp��G�?�ˍgG,L��>��5U&��uYk�u�H�)p�� ���\�	O8+_�<zܾ8	$@����I�eZa;Q�pn����Z:�8�H�;�S��x汞-$� k|1�	���1bIMŘ��5�Uڊ��򊗦4�4�'��.33 RZ��>���W����`�9��Hm����^�B� �Jȓ���?Ir�z��5f9T���֞+	a�`%�1p�Jn[�:�R�5���֗���g�nU*�8��o�x������uc����q ���5��6����LCk�ցǟԳ�_q��H,���*m �g����=�g$؊�\f��Tl䶝p�z]Y��/|7����W������ZMnۉ�Tl����.vq��EJ�Р>JC�g��An�]��`�����k��v��j��d�t4b��Lz�A��!?�Kd�����v5c��Sp��r+sv%����4M����N�=}�N_�:��w
�ww|�F-��oE��M�^Z�Α��v�\�G<�� :zy�Rf3����$a�cҨ����p5�H���JK���C��8�E�*�&5��q��V��S;�O��8��6\=����Ъ6��~i�V%�VO��B�JL�*1/,l�+_�x;Ώ��\�$H��@ �"sB�վ�eq���K���T�M#X���8F�'o0��G�4������A�M]X=��*���!��`�D>57�]b� � ��4��=�����{�I<]X���ְ�$npy�08S�%Ä��JΝ���bd�I��],��p5b��o�e�s���,+tt
�.�ݪ�:b��B�L�F��ڽ��?!��&0�
��FO�P���{J-׆�ͦ(�h�ֺ<Xo����8�Zt<����������-��������\������Ь_��뮣�8�]WD��_�&Gr���D6!���Ss���~�%�ĈC���H�w��}�t8r��w��������؃ܛ"d�lͨ���&Ԃb��5�Z����~�~�=^�Ԇ�$͛�}�+�G���9VV]V����채\n��f�����_�Ln^�J��Fb�+\�EK[�Ἑs1|��&����XM�%Z��\�\ũ�h�߹P6p���)`�O��)�_f��.�Cl��-�j�"F}��y���z$��_"�d�:�X�|��o��K]���iXOu0
�Y2
��7�p�Qm��H ���d��9h)��=�e7��9D����+�Y��QdWomgQ�?Qc��$W�vT���G!�#�e�r| �0��ϩw
j�潒��Y[5h����~!QC@!'�ZK�����V��R�t���<pm)À�EE��ԴM�����,_��,|���$�J3ǈ6Y+�����Ѹe����1�}$@2?���JV0M���B��k�yӶ�'���L�w��('*���̬1l3� �*º���ZI�T�I��x"��n��_׸p���A�-m`~�	�mC�'�����.GY���-=c��U����D���Q$��Ħ�٘k���䄶DI� ����Ħ�B�υ|�\0���D��q�3�M�ޒ�d2E�T�X���;)nS��f���e\;�*��%�zf����%���~��~1��]Z�""�\Co&ZH~r��x��0��QF���҇K�h�h2Ŝj9�Ng�.?�̢F��dތ4���-ľo�j�>r�@|S���g�V�ԉ�C�|�4؃#2x�J#S�Fc1��2[���^��h͙@-�B�|'����f�ee+��!��͓x�0��bWBG�f�MK�T�`I�X˯.(�"a0T}�U�u�
��"V�d�:eWH��3p��=�@��h��Q-g�[�!i�Ux���nb��	�P��ï|�5@�/�+,ǈ4�Q��<y9�ApUH�o��G������q`<jO�/�E���Z$�oIP�����������A��bP���2.�f1N�(����\��o��o��\RR�W�;��-�m���-��7���2D9D�b��O�2w�>�9ʈ��}���2(`�Z���@>x2� :-Rsa�lϬ���K��ZX�4[���{d�٬�4k(�{�������4쭏J�R�q��{�

����j8�"!��0��U, ���H� l~Қ��N_�c��K�H򧬄2v#h��/�l���@��6ݵ)l8i�j�;W�qy�[���_��Ozj�͞��x7�z��-ׂ��� ��$HV�k��;ް�J#3�����N���<���fۓ��/ڵ?AD�q�B?]9Z�^����,ovk�w;�|�x��PT7XR�����ǡ�ݯ����.��.�|�A��*����gW�eP&'Bdt����a>q��K��I�ʌ���	2/`~t��g�TCo}��P��(y]r*X�7�D�y�wt�s��~:����`��$�/ܞ�(�S<�M��i:[OI�C ek����Q��1t
��4L�D?&����j5ڥ(|�� ��~ ϵ�QgZ`LS��qh�vR��8[�[��Z�����C;#XOl���d!l��=� �{X�ʎl��($cl��a�ZxBT�h v�	���u��~���e�)AC�8-� �m�N����1o�6p*�#�o�f�G���D8����m�:����7�`9�-���	�8ɴ�?�"�ZDy{؆�w��\��Ǌe��o�;�qI�&Hц���[�o�S������[�-y��V���q��h�c|M��z��:�
N������&ݣ%y�ς��pf�\�n����=�٤"l���f},��/�h{�3h�Ϗ�A�^�{R��+����v�z���ڶ�"\�TB�R&�`j�����ك�y"�{ʔO��6'����`���b��cfs��U����>�&�]RӘ�I��ug�Q6���t�	�	|N&�v���&���,?�*���B(m@���w"��S�+���`��8�$�:p��M�c�(�˘ �+��)���pD����%?U�B �L�Q�k��&�j�Y��0u��@D!>^����D\��]O���+Z�Fzf��8��[!�w�5�@�av;p	�O�пφ�H�1��nrYc�~�X@$��|�'���p1�x_M��E�P,��b��e��4�40'��..~R��(�>��wT�v]�;��9�H�G����^:ȹ @{l�+��ﺔ��4}�p|�T5d�֙��	�r�%Z�*�e�m��y��
U��o�L�C�	ʺ*��*A��,���~q�u>��*� 3Ð�0�26�����<k�ߔ�(�:-�&�<,���%_\��L��;^���m��ûe��ߖ��G���;k���d���������VMI��鏹��S��vl*W��v�[��C�������n��Ƭ�+/݆����ўi�%��d�)b-
<z~����f��.��.�������p��r�%\�������|oN�&��^VY�������w�jF�Ȅ��lܟ�>^UM��� 5�A�<�l9:���RAkA�%臿l�c�'r�@*�p��H�5IJƕ��vW�si���e&�a��%�I���n�9Oj�a{�y\x)9�(��6��(i��J	z��f:*��lKfn_�8;�o��q�HBTy 06�"�ՙ��q�Հ�Ko�Ot��WkXAP�SS%'������4N�����W�A.U;]��E�%ꜽl��>Dyґ7�*�͞�b6�V �S��� ����đDIw��X'�p֫�n�(0�I��@���q���xs�,��dR�N�X�]w35��ĊR��|O#ڹ���[4zڔ��L':������=�a�.�U�y����!��0pD��~�F��2�z�{5���#6�����Z<��>��	�/_]��M�d�A�������r�G��;LX��gW�s��@O]2\�����T�{�v����n,�S2�/��L~�����4���؟��ң�HANt,s�rT��h��2%�s�^��0��O&���y��L�ݎ�5us}�8#��h^�	��c�8�X+7�L�9��V1!�����L�jn��9��F�j�L�Z7JLW�bz�q����|N�s,A�oT�SlXh�'Z-h��vݩ�q��z��6k17�v�W�
s�Dݫ_�.���l�3|�=Fx8XyhP4����$�J"L�':u�Z|ւ-o��KX��(O�X��:0%4�2�dq��r���ɐ�]����u�3h�7)�X=%7���*D��ƚ�T�LQ���m�_�Z�%�Sfix��T4�[G�4�#��r׆�0_<��
�t�m��YB�WhTC;�zY-~|�@���u��I��1��t����7�V)=�E ��ό�cҼ�x�,�4:��U��J����+���L&����1 6�@������V�_W������1�2\��{���@L`���#����B�9�Ll^�{��*�)���R���~"M^>��ӓ���H���m;�n	�F9N(G��ݵ.���,�c��ݿ�%����7�:��$9KΦ^��)���N����k/��8W�}��� S��W��.��,���h{�4��E�#<ᓼ���W�nN���!ț�;��֗�$�fz�O�`����?~q��j����L7\^�Z��Mr�:A��@�Yi�������?���hM2�j�'>)'عi/��g%?F�}��疗��9]ox��>M��|��߯Vk%��֧�7י4�ƹ2�P|J��@�����-[x���]h��@:[�B<n���>9�G7X� )D��R���x���}p�GX�(�Tħd���3.#�,apq�}��c��
+�n"1{|d��W�73kW���M�@B��/�}����6�i-lUx����i�p�M��P�v���V|@S��
ĭ,���j(7t�9�sU���4��jB �k�b<��9/4 G�I"Z�P���+c��ct���	�Af%PJ2��-''f�fF(�㌛g��/n���<�H�&\��1�R���&P-uL�᳴����Ү��C�y�~��Js�2n�b��>I�0r��d�}d���i(�g����>�˹ ��ls|9��'�ޞ��ܕ�4��<�v9L�4q�ﺭ��!J� ��YR��D���Ի�ki
e�{ȟE��=S&��fjUE��	 �3r~�UB"i��9.K�eʧ'Ev������}������{6�p�lSq�jZG��L��Ė�+�V�x�Jˏ�c=n�y��xR��z[�-����=�t-�V��N�x�Y�PQ#N��/1UN�_��Iv�kqf�z������ҏD;oB�I�Z��#�L���M	k�)*�jmTx[�kPo�Rve��"�x�=�y.�@A�׫���Ғ��,�W?��&���d��i�@r�>f�qA1F��|�X"��2
ݲt
*�g@tbCj��y�PEp=(��%*��Y��hy8�~�7y��>�`�T��?��/W��Vd<�x�i_�V��I �e&�=������u
u+lL�Ek?��D�j���(7+2 ���i��`QV�X`�S�l�@v��8p��{�w����l�ʒ��e!��=�l̖d��	����]�$���J�I�/uB�-  1����λ�jY����o)|�X8��R�h�4N$��h�j�QR�ߞ�x�A�u��D�K���q2���Ur�{k���U�b@�sD������Uz��_�24�2��BF�e�^�*���lJ�&������X[�H�ΒA�l�XĖN{e�Q���l�4�#m�|hzc�����QWs�sJ��	��Fp�<��wS��"nw=[;:���x�wfx���)�n�#H�3�U}�)^�R�$R��\��v��9�K�C�ݳ�T]8�R��{jp=4�7�5���{Ōe�;.��N�`�$�b
ix>�Z�����>��3ָt똍��(�gF6�k�t���̭C�N!e;�2}��{,Z��*9��B�c�%�[w�)�S�� �z`h�c8 :�ή�(�]�c����h���O�ap�����_?��N�LX��h&�Y�Y!�#ui\�_���e�~]\��On�;+U;�z��8�2�v���7��?*a�Eip�w��D��7DHy�D����mp�g2c$�*S|g����1��M;���k�ڀ76�@�74U�''�)I�Rw��������;ҝ��9I�H�rl��t�^�mM ��t�FT��5 E�������T�a�֔G�	C*%�i���00��P9���e8�F<*g���u�G�d��r~u�!eaT ΖŞ+6D����k	�ǕM�	��a�A,A�� q��w���b��,���k'��BO�,B�װ�����w�V�������	u�M$���&���Gvgұ�x&�DoC��,���nx�`�130�y(�2��so���N����@��c�{��~-��I�)��mQivސ�#�f=\�$G�Ѣ���Y���}atlf�&��;]���{��R��k�*G�<�g���@e�fp��K�ox允��(��a�
-���8"p,Ś����	���S4>��50��O/RZn߱
C��z��Z=NR�E_�!�^5�g.�s�����1�:�,� �Ĉt�lw�7ZmgCDl�}��|Zu�y~�A�s<_O�tX�hjZw	�(�c�����/��AC}�������f����Q�(W0F�S�7��Y&�B����$(�ݕ���Y�FĠ Em���,���Ķ�6F�)(&�M�������T�O�c"N��<��]��5H�����v0P��G�O�h�B�|����3ԣ�ܕD��34~��1p�i�n! �`jPC��j	_��O���N�"nz�HM.��63�D�|!�(ȼ�@*N{����o����8��ݪ�6�}��AH�9g~䐧tJ1|f������'�˅㔬�]z�➨�@��狵�?"=W�GP�r�(˲ME]%{"�<b/��o.���7��l��{�Zp�O��������DB�e���7ƌ�<������n��-�_ �#*D�Q����[���<���5����~� VC�8�	8b��s���t6�j�0���9�M�5�i�i�ހu���-�̤pm�%=w/�����şq/{&����DC���q��'RU�3�R��2 X���T�����g��b�� ���R֓��kdvG����)�|R�/ɽ�&Lo�V�0��sy<��:�߬�!�Qg��>���-�Z�g}�yC���_sK�|��X��S�[�T:.��lC�a]��/�7�w`��-5P�S��_ػ�Q��&UdM�o-5�?n��;`�/ۅ}9��E/QD֍�	��#��-��#�я�2/P����TO������o��d��?�k�d-\5�6�	�\-��Y*�d�ۊl�Ԣ��]��H���Y�n�_����nVFϥu�x�s&�-���2u���V/мw�nA��Sr5�
��!�ȝyIi9
����@z5,�EC#�:�a�ov�ȃ�^���.ZY�Ź��"}�}?8���kZS��g�ufͯ�o��R�E#�"����4�b��=��|3[F��oRf�t����mhF �J�IG
h�|��!@p6����G��@N�7>seIR?���!�v&�k#p�$W�M�TQ7����ɦ�0%�_ѭ�\#�4!��!@u}
4�������>�#C0��U\-�B:�!W��`]�kTf������]��q���Y�׆��XD/���n���8��;0�r.^�Y,��܉E<)!�h��d�tq�r����/�T�	vAvU�	>ܓ�Fl<�3l���O���k������z[�7�>؏e#��P�
�os3����9�(����GM�݄�����e��֦$H����.�(��*�&����S�ţ��$e�r�*�(R79j]6ƅ�?�dg��Z\�#(W��p��G��N�L"G�mN�+?5	�D����DO��<Y�P�7YpLL����=~�R����Ɨ� ����^��n�&�jj���2��3���+*�Ch�q.׍gr �����M���2xUX�E`�8ω����'�l "�(%e�0�e4�}��Zwk�;E7�������˟p�����y��(�EEZ�n���?lу�e���AE��ZJ��W��1�מ8=N��<�B���S2 Y���F�9�%�Hc��o��5��\ƁOSf/�F��[\̧\ʴ�/���| ���?��h[l�	�T�[%a.����cl��75��v�w|h��6�{��AY�K�ª� }5��L�����f�?�ߏj���'F���f��s���șs	R�KF�Ǌ�pxC?�ކ�m�$�������D�29쩑�G]��f����qm�O�2ڡ�?|�>jGG�ZB�x���;�_�K��@T�V(uz�;G�7�L.���S���,\b!��IeT�������懎'��3��~�K7$�!2"�fyŻ���r���������������C
�P߯&��"k��������;i�M�'Wl��s��(��-�XD�2�����b�3VCU%�'��f��k����D��z�0�1
b��{�Ug�tjx�Zg�<�(ݶ�I��6��$i���-z�w��'�?!~�0��+ΣO�Y"�*	�)��Aȡ^�GC���p㐀�������Y^ӫB�a0�`��\���b�h��,Vƈ($�����%cJ����)���ՅH��J\��WAM�V�ɤ_X*�Fҡ<�w�6�$L5��6�[lJ@��z��_���d���|߱�x�c9�8����}l�&_%V<�"A���9��?��'�9�\�~�LH���Q��O(lN�ChG���,����aN�S��)�׌1�\���jp�d�C�d�7�9�XW���[	��ϑ�)��;���e��Td׾Kܜ \)�Z�h�籧׭r�)q�����B�v��BU�P>O��{�fU��?_i��m[Q�>���� �t>KS;#��P�v'o&���9�ы��ZQ����f�Yְe�ǡ����Kr�{!�*Ow���5C�&���P�e���*k��7,5W6��?{���i
#9GZ!G]���������Su���|$d�}��3'���ӕ=��~+R/�}�!�R��6��Ö?BB� ˸�̴[�~gI�cZ�ؐe����[�K7�y�}\��P.ETt�=l�4>��aT�A�3�j��ɮ��2�5�Kb��#�j���w���v]��G�r ��2sS<���D� i��;�%g���\��~���uc�HYq�L��{S1��RDA�����(�Gv��YX��fJ�+����D�32�4[Ƨ����:�E��λU��@3���}u43S�����!�D,k
ӦN.��@.�e<M��$51%TN���{�<�eK��	,ߟ�t�E��x%hx�Κ�=��tNu�pC�K���iJ����
��ͨ$9��x4����F$�����r��d��S"�e*A�N����2�����d���5��ʜq@/N��B3�ړ`MR�_p����yI�P��$� �A �z��>c8uO�� x��P���h�R:�-p�����9�ܹvu�ly:�[�G��P�)S_�g��:K�9�fu�|<��'���WQ���քd�)B(������`�\�zt�X�'kp��<[�r�8�a$��޸�& X�D�%Q l���a���s��O����-��r~{ѲxS:H��2������rg&��~GEƇre��:�k;��8�L:p���KҔb��88���j��t��h.���kah�"W�B�T��9�&z&�*��P��Ӊ�O4!�a׾	���93��>�C��;���<3>�0Ӏ�+ ��j=q<H�����;�g�h�����L�;����V��H�רm�$����9YXY���Z��|Wc����Ja�r ����p4���ې�S	�Z|Slp}�1�T�>���:�d�A�c��v:�%p_���U��;�������m��V��շ���|6�c�����S �� ���'V��M;R�h��
�w�װ�r�Q�#أ�(����dC�<�%}���� ����*mB�ԡoG�
�[\�b,�}�/!B�?O��N`�BW��h�2�
�#�o���U��^L�dq�ȅ�)�W��A\�Bt�_��躨�1S��Bd38�	����_6(��֤������1�!v�f<�h���Q���|Aq��ģ�GZЁli�!��}���(�q�5�]C0H���pf&S�<��=���:�	���r���S#�������Sӷ��������@�8�r����3�;�
ju#��� �~��Z����N����PK̙��"Z���ʤ�q'��^q&>=�x&�h�Mar����"k%
=�8#Ts���t��&
�\RI�8�uW<���ZJ!5��s�T��CP����]7�MII��U�o� 1��3�3pq���ڵw��S�QM䬶q����9�H'��8�JTڍ	?L�#�/�]����4@#U)�E'md.,O�yX#�K/�>` {p4�f�����ꥱZ��!ײ�5�F����qLRhP���3�8��m+�s"�����ݿ�����߉����CJ`��-j`�B�����iJ����z=5��R��B�d#��쵑��z� ��`���G"��gAλvB��y�Ԟ�Tşa��l��-O��D=�vP�K�3�lq ��i{a�*����I!A�D=.����+��̜W��>irs?��>&;t=��a��C��D?���@i��b��'�آP!��-X_C�uȰ�(�%O	T>�D6�^�[�PH�u�����BA)��	������b
����%.�J�x�,�45c�8¼�x�[�f4�]�T*�hHArg�l��;+����.&�d�'y�=���Y	���rH�S9�w�|���M�l��*��-E@7B�r8 ��Id_��#Wd��v��2!���������3|Pa�x��_Z|+J� �q=�^GA�=�>P&�7.�c�����ޣ�Fk{m��N��sgA�t8��&`��h2�8ť2W�2��X�y!K{�s�[���1W�t�*6��uiFLu��������n��M!s$6����/��;���L�{�	�����=*҄��6�ED|�H#+�g�c2�zU1�t���������_�]���������
F@��]��uaNs�iD$)�6�f�8�D[K�7�|��07�f��"K#�ڨz�2u+�K4 �?�A�
>d4q08�U��"��q;!Ӏ�r��k�L���X��/��σӝ�c��KgXY����N�Z��1};7��=�Kfם"[�[ӷ)3exh����-r�#���Ɖ�Ȁv�`U�R�>��v���X��r��~(ȃ�^�P
u��z��(�>�4#5��P5�oE�C�.��9�ϋ�#��ݖ:���aOe'����R��νzT�*.
��Y$���՜�f�?eZ�h*�{7K3�6q�?Z����b$�5*�W��Y>�Y�d�L4�m���?��bD�F��VC$Ў�"��H�	�pL^���*����Xv��I����v�TKB^���8%9j��������O���'�����_� ���8�6�e�1x'(jErSu!���|���� 4 %��������OFZ�'�;�u�͗�����R��w�<�ͧ�a(cy�Z���xlc�@7�ִS��լ���`���x�$��>�8����(�Bě�e�YU�Ff�%��:umo���@�X�S�hS(�>Ҙ��[�#�\���AI�e�� ���?���hm��	�3*[�*������l��5B�vk�h�΍c���0?`Y���¼Vs�7��5Ei����H*�,�,A-�<������\l'�Y�����sy�m�� =)�$j���[�a�������.0O��=�g�����W�^����v`� �Q|�}:.f������:��d����Ģ�Yv,�[�׈ͦ~��T�д�q1k�xH�H���yml��o�w7D�M���"do�ETb����k|*`�H��b�-b���oA��n�Ϥw���oe�*��S��8�<�p*�+e��0����w�c�|U=��`S�*Q�V�15���)Xo����^���#�):7��B�yQn]>~W��rk��g�y����&�dKZ���	�S~�T+}O��j�,�L�A75c�`�V�O=S��ج�c��Ԝd~=�-�+n.�`~}�ĝ%�|�Q5���w�T�~-ք�)���~���+�%������Ҕ�-�6�,8�k,�}C5z���?Z��Y;³�ޡ��ų��4g��L�w�?�-��bn&z��i���\&	�׳�Y�2&_��'j�nR�S���iE:�����.��i���PDO@k+0/���vy镋��������o�Z*�*����"��5���S�Z�.g�-�f~��o��K�6��".����;D4�Ӯ�C|ı��6G3o#��t����~� �cyI�|
��|9�!�q����X�QG7o-0IoRa�[��)�ɚ��y#Aŀ$Hʡ�e��#4���ޜ:��0��V�^S?#R6U��]�u*7F4���� 3�>�0�g�U�t�}�!��v�q�+k���K��α����&��W%xX5-���JV�-�G�;�P7���cH����E�z��)2Z�h�ts��6�r^l��Eo����v|�U��h>�QY�w싱��4��˃8���4������W�>���#	�P�Q�o�d��'�9Czh��9�8�ݕ�"��C�e��R��Z��c$ν��*mﲉx����3�E<�e<O*I/7���6wh?�nA���w�4�W֍l�nģ#�L���m�< ?T3D�1��U�"�m��cڨ L�Z-���#����d�����F�
�%^Pz����j���2�$U���p1�t�W�a>���� �ꡗ�O��wxF nEqO� x�;xP��g ��%d�6���n��Z��!;v``�V旒3������/
�JI&(���Z�6��o�l"��옴ҭ���*��ݮ������8n���pBc��?Y~u+F�K`%���tQ�o�ܺ���A��+xS��C���3[-�\�a�@��Du ?D�?���h���	\2�[��������/�l��5��v
�hrNH��yJ�o�_Yպ�»;���5�{��'��?P0	�lUe��_���O'wMBԷ"RsNb7l=������zpa��E��,{���)�\�m��z �����҄+v_Er�0N��d�X.Ub�s:DqL������vM [�L"��2��I��3��q��÷�oH��ex���a�6�k���С�0���Hb�(��F�*_B�'��!ǨbX�o�9�n4F^w�2����*�XU�o��<������D�a淥t�w"u�|tv��_k���	Q�I(�ƄC��)�Ú�`��`T[޺�?�:%Q:�����#�l� ��+P��,8)��V�	�5;�Ic�y<8�ݡ�4��+�uа��}���<y����fF?/N8A�?]k�)�2G&)�e�rf�s��P�=�ʒPN�G��֨�%����`�E��m��z��2��C�V%��Z��z���䊁�1Cٮp���8��z2��욟8���D~��]_�AF�5L�1C۹ o�y�K�c�
-�e�	�$�F
+V]Xw.Vw�ё�1�AI��02��p�>�J���m�s~�OU�P�*�g�w2��7������G�ۗ��m��Z2=��??��>�jNGp���[�6��3_�
����>PT�4.u�'�Ge��L<x���E��Kx!�W��]TbvB�����
����q��qi��!5Y�f��O�Ğr�K��2���t�`�-�������ڹ��j�9��:Kd�Эr�_���>e�GH`��3����h_��`�0B�W#�T���uu��G=h�L�̼�n�اr$!����T:N���r���ť�D��u���!�mf�q��pr�v �
q��LPE�����싣��݊�����N]�s�2��E~M"+�c(�N�s��-�����q&��wjb���C�G�����/4Χ~�Z���,�)��0B$b�#����@tE�%Z2R�ףnݱ{K�i���2��@��A��TJo��q��a�U�N�1�-�8$Eo�wʴ��2��Ά�
[��)ڭ��c�g�d���Rg��J(��PG�t�p�/{�}�c��D�ҵ���t�Fb=DD�~�)�p��"��v���a=��$�:�� �=ϫ���|V �~ߨ{������m/�+�
�g{���$�8kE^��@+[F�ie��x���i��+�$E�@�ඵ�ƕ��~`�"�R߁��@�6ɶ	�K�B*TS˭���IR~��c/��wOk��K� ��y�O�����P� e�?�����͟��ߡ��N	�Ԋ+j�c�CZ:2��[�DݥX�j���w��1v�}�<Z� ��2�KK���D@��l��ŭz�o�N����ӭ��Y�?u��%�0C1E�G����r�����GK�jY���{�;+K�}���3'�14�Zu�0L����d��jX�@����e�3H�~�Q�I��KD�>7@�NC��@�̆e��X�;71�r��;��{�T�]5�v��T`��V?�mP�h���ӓ�Ikn���K,��e�r|��t��bQ�9�gx	���s���n�������N�H��e��"N�N���,�B���ك��3�s���s�N�J\3`�`��dt�y�?��I_,��� P9S����u�<ж52��ͽMH:�+��z�������u]):�ZMG|�Fk�Ox�����o)�gR���d����\u+}c�O�:�T�M��2���Zm)q���xK�\�1h��f�~�]*+�R�f��B)(l�n0N���:�z?b�j���:V�FI� �aȏa��Y������Z[�ሾ�U�rP����yb?�4�X�5Z���}d�jjw����O��MU\-V�����͐��T����黽�A�*��m�j����ZӨ��e�U�*lna7MbU6Z�w?ܱ=�FJ��7
�W9�����&�/L6m��m?I*TDt�ёX��Є�&Eo��F`L`���l��f⽨u���P�Sͱ��^s%��:�Wj����E����߉��"~�$��!�� ��ȡz���}Xx�`Et�9c������mC 6��%�h�y�>�)�Z�q�;���r��Vm���՞~�����J(%-�Z�HD�Q��l�2D�c@�U	#���%J�:?���L58ѾT�3��B�#�gʮYat�F�&U%W�ow	Ao;�j�³����S*Ү����[p��\^�C���& �?�pbho��	?�d[9�"�gz����lk5ă�v-Y=h�������l�Yxז¾�G�y�M5Ǉ5����,����|��sov���o'��b�z3�s;w_�$=k~��q}�a�Q��Ad��ª������ū��J��uz�vb�ד8��' .(d����:'՛�I���d�vJ�[��v�OM����жf�qs���_HV��{m��C�"��?W��G�$�f���1b\�*�N�*b�+��6�b{p9oC�-nCXw@�6�1�*�NZ��|�<�=�������%~�W?Kwe��|+��b��"#Q��[K0��ư)�&@; ���޽�Z?\W�Q��͖�V}#YR��q.+���,��5�Y�Ø�H��*��8n�G��B+,[ư��}���<�#��ŃFb�8��]N�&�u��)����u�vs
�^rcʵj����r֋�E�A��``�,��U��:c-���C��S�f�s@�Naz�-�1Fbprq���>zU���G�ބ4~G�]�iF�������B;��� ~��:
b�L���p�F _+�^7X:\�w뷊��۷A,���͇\����A�g��Q�m����$�נ�#�v\��.W嫕|��ƄI��6�Z)�	MH�o�g�C����1�6|��.�H�շ�ǔ:/]f��m�������+")ai��Z�^�L� �]�"@Z/��<.�K7����Vo��FѸO'W��lb��r��D9�e�T7��<�!�߇W�6X�K�_ҏ�XD�t��f<�GN���������0��j��V�
�����b:��_���?lԞVk��-33�9�_��z����R�Һ븊@p�>J=c@X�0!�ŋmp�{���o�ɧ��g�yܾR�p3-��H���YtZ��\�mJ��N+����.F��g�ǍW���L�x«�J�v��[B\��S���I���X�-}��TN��C���(Zrqڋ�2d��\�I�J�6��p�R ����_��qYp����	C=�K��K��L�x��M	m�����/��Xr�5����K�\���P����D\t[L%;�f�TtX�[*}�5n�!�I�SԲ��4�¤�%.�{�������S���ca��!���΅8���cp�V��-��+�:���U�Q�/ːj�����\���������g�q}�h�f��Ǭ!��^�2=���<�*8���xΆ�q�hf���K�$xv�l���}�Y�at ���8S�_��<N�<#�����!岦XRk�3�;���rmύ��R`M�_�#^���g?�p�W����T,w����tW�B�(s�gTO�l��͙u�꧞A��I��t)2*[�h�I������/�A��x�_���ϒ��=b����iΤsƳAE������b�(��Vɸ2;� ͠Q{em��,u\��U�6��^(�.]M�j��$�."f���P�c��W�k{�:+���������2�P�듂��<�є�,�3��T�f	��$�f��ndԚ��!Q�`ۿ3���j�n�� ���?��n��mM_�6�����qʩ�&D��Z�{�߲�`����w���6����\H��g0Б�x��1m��,mR�o���l�&t]ϞYn�����{"a"N�K�xv4��k��#A�]���"��6/��.��-7򄽸�v��qO,���y���o�D��e���7��<�'��DFB�;� �p����iD�����&�l�ʵm搞_ڃ�5�a#V�߇��Jb�t �.��\���S*�2(m��T���X���G���A��j�p�#K=Ƚu�5K��0��,;F��9�mT��D��>�&RW��3$�P�Ç��?�6���ؖ��c�sH� ʳ�R'�+���dooZ$Ӭ�����(�δ	����|��-%�'�'b9��~��}ڢ���sQ��V��1�[�m!��~u���b �W�� ��R�M����e��@$���x
C.y�� ��nE��F�/����z�y[�����2�4ǉ�&Ԉ�d-�7 Hd�z�]��Gm9��<-+��J�ju��	+Ǭ���H���pX���q�b��t�I[>y�!f�xE�g.i~�q����-m�SBs,�9� ��{z�y|��.U��W�@~�_
҈���)�S{c� ց�������U����
È7�O�+C��ly[w��8��]U!9O�T'�K�&��q/�y�!/��p��G�5��H����<g�]1�/v��4?�f������r	KU�ʎ[q<�D��1�΃���cݖ�U���	�
N&�T�Kq�Z-o��{S�r:˖��]{�Y�)���ę�����h����~h��U5mc��y�s��z��M6��&w����f M��bJt;�+�E��Y���4�e���}�N�j/ �yJ�$	�H&\�h��kT�&3��i���U����*�(�Utq�2�2�(C-I@�6��T�e�/��_\�qwU9�ha\C۴�©$�K�5L�@����m�n����/�$0X�
��gpK�ިТ��X&\�^%YQ�f`��X�|}Tj��?۪I�|�G2Փ ؃%LS*��m��z�����+af���:�w��q����qcN_%Vo�-����X�|zQX낐�*V���I/@�C�D<��6��!�s���U�ԝq&�[��*tS���7b���:v��9�Uƛ��6�.��M8wm5���qrVj�J\K}��?,ڢ>�n_ப!b�;}|8��jU+����|zR��O���*締9���ʵ	nH5H�*T�y��R�o��q�ei�CV��5�y	.�L3�E��-E�cD��60kN�l���x3��0hj�Oԋ"x�,J��k')�����q4 |�|E:��e�x/�	�!
;
�tbi8�&Ҁ�س}��EM�
��v�0�O��i$�C����=%7�T��6��o,?('M�
��$Q��q�3��e�5�V����B,I��q]��2{�eGW�TZ����ݱU>�J��SJ�9BӇ�_�d�[�N�k,n��Z�.qO�@��?�H�7Xf %���@@��y��ྜ���Or���n7{:�K��ʭʭ8r#�F�n�~!	��gb�x:�}��F�#Lv\�R���h�S���֌W+�٤���%�a� �"r]��+79��&�uzT?���O�r�aHꦂ�+33�f��X�;1�<;��9m��_8�@�*eQ���<�����^�βd��rϝ��-�X��	�cvN�2;ۺ�gZ|{��B䁖C����{����՚�Sek�6���S}�HSh���5\��H�}����� 
�yW�����{�Jc�+�`H����h v��3��̂�������J���\i;��|Ϥ�B��,�E�ޮ/�����(�m7q�D�2x6l��|I�l�6�$z��4�2�_��Kq&����CJ���j�KL��L�V��ڤ1�=�^Vk�/~�{X ��L��K�Pб�^�Gh�\�EA% @f�}LX��}�n��ni�I�kM�6ѓ�k�%�`s�b������ �E�Z�̀��j�f!�@�Ğ9�c�A&ţ�-Iya�����7QG��|���5��BKu�*J��݇�e�I}W�f�m�����+�h���IP8*�-�����^�fN�KPlxCz�����f��a!
'�f�38@Ϥ���if��Y��q���ķ��_�R���(�?z6��bz��-�R�A0_ӡ�^��Hg��4�����p]��,DF�/�{td�ѕՓg��5lі޹Z�w�W�AR`�}��t6.�Rg��孺uΥ6/BhrA����8@�x�Ad2�Uu���1�#�n��ࠢ��"˿(�U��ej�8.��>RYmn�I,����"�6d(b�M����q�� �-Bc��b���꺧�A���Aƹ���-ZVP��)�-���/�Y2�3�Q3�s�s�����*�zԇU�!�,6`�q�Od{j'K��-'%��i�n���ML]6-��,u��&F�^T{�4��*��V���16���/XHn��g�渐��1N0�y�e��թ���J��]�	i�ơ���Q�(�T"����e�#�P�l�P�]�S"� �/�e9.>��7?�/�?+�8��OYۉ��l��$�nD� e>>7$�)<��^����h�����Av'D��A�@�pֹ�O�Z߷�����bk��N	Va�+��bbJ�+��:w���f�H�p�_�}���:��RZ  ��	�
G����`�%u�<@�]]�,/"�4k�d�-7��C�	�?pʺ��<-����,��/���������5�	�c�NR2����ZY֝��.���'?{*w�Ղq���D��;o�+�h���5w���.���)��y���Ҁ64���%��ț�J ;H+�W����ُ�܎���@�̟�Jh�tz�\f����
���6�	��[؜ѡ��`(�"Dq���2�{��Il��6Q����ۜ�_>�rq#�𶔕�C�n���<Kɴ�Lժ3��|��l\S&�/�*X��Y�)ÓK��7���#��g\�!�%�f���X2�}�1��뇕I�Y����LU�%�u�����X�2������؀�� �#@>���ě��czC.��-&Vp����/qQK]��|����ߙ?�L^�pG ��[�}��Pfgf<�6���(/G0	��_�*�$�B�Ѵ{�f/K{m�x@Ci������a�������8]��`�u�Ɛ���ϩ�(�����<)R5�Eg�7v���č�P�Rj��_xd^�Nig	Ei�C�O5$�,A������t��T����gvl��/����t��AOݪ�ts��	��l�����b�g/��gA���i�����9,�D�����ލ��B��yK���0(���B<��;��[Nm+!�,����6"&(A�Mi^ɺ�Q�,d����cj���$�D��7�Ɩ��Ϫ��P�S���G��=�^�V�3��ܰ���Z.ϧ'%Ԥy�!���`e<H�L�%j�5��je���ocnU��MiN�6�A��wد��^�����{�1���@n����r�6B,��h�t�����u4��`�zc{���
�����t�7i=�Mf~�c8p�Yp�N�s}Z�a�~�*u��fw�=Uۯ ��\)�D)x�ի���Q/O�ܐK{�#$�zE$X���Y���ik�>^�N����$���#RJ@�����)pcq3���SlK��S�����LV��� Z�R������Ud����*c�e�����|��NC�煥�7i0�dy]�:�F.��"Q�vn>Nz|��;��g~�yd����BmK*���١�SN�T�ɝ���b����7�<`羥��eS��P�|�Y�s�VdNΝ-V�-n���`�օ����Q�r��z��$5-�P����O����ytb�)��x�t���8��N����k���ż5J��rA�$hY�2��������R�7'R�k���B�jkn���Ϧ:C��&�6��Y8<2�9��<2��8�n"��Ssk��9 ������{�i�Xٻ �/@;(%�U��F��[Yְ��䎿�ȩZ������>"^.�WY����Z��g{| fN�oV8�xB"�＇�LS4���~ZZ|��{�@�o��td!�N�	 �D�Ih�
T�z|�'!��`A7�����!�7?�fI?n�+"*��4��!<#x�$�m�51T�����y�
�T0����.�5#"��i:(u���4�A!�Н>Ӵ0TƽU��n���! �A�kU$��&F��@�Β/��'HX����a9���]��;q���Ӊ)3!c׬���J�B)Agh�5ű�Br.���>L��]�v�>U��[>���G}��T����i{^^��T ��D>�U�#�i�P�̝o�9͘}�J9å�������e3-��tIe�+N�e��3cǽ�&�*="��H>Q�-O�==e�V*�7��K6G=?iq��s�)��W�^)�Y��g�L��_m��X?�&�D�^ �%Y��=R�3���x#TL�	�Y�}��M����V��!	��5�&^ _�i�j�n��r��!妬״�D*H�1��Γ� �3e�g�t1�x��EA���"���ha� ��%���4�>+=ZX��;FA��&��c����R�k�%�,�(R)Z�v�� 0l�^�����l��]��o�!�g�K����8>:9�@�6B3��*�YN��Fu΀%�qD��o�-���Y����jSw/�����[�q\�Wg�ƪ�����4(��Xٚ$q!-��G�	n�+��ZT����+\��}����#��QGk�MN���t�-��|��v�F��ݓ���{���r����.�k�L���5��;M���=tYn"�D|���ڢl5CZչ_�x��l^�mסnY��i�἗Z&\쥳<�)29:ӻ�����-n�iS6��\��Rdy��|i���D@>:�b��	�͕~�T�3=���Z
��NZ�Oֹ�"�3����ᘊZ�g^{^f���o�S��	0$"a�Շ��4�h��\�|w0�I�8o��ytg���z P2I��K
׺�|ь�!���*���[lք��7ɕIb`z��ɾ�%^�ŵ�#���$�@֘}�����/��N0iY��q�w#�ȟ�l>�u]24rR����>V�07�hU �y�t!������kHE�>��!gJϵq]��|���=�XTw�,L���./�:-�;�����av��O���M�@)e�$hp6����r�gw��ԏ�тv��U�?|> Yڟ
�-�w��p>���2M�di�=#l����>YA#��dP�4�o7��`�-9V\�6^����9�J��e�b��>���>��R	*����K���������e��*��7}=�6���?f�v�1�g��Wi��O�VM�Lf�mH�?y�HD�MY��(I� �V�;����L��I�|ޖ�ҽ�"��+�������w^��i�jemj.��6�b���ɦ,���T�-�Q�Y �bn��C���x��E�n��=�.0�뒄 fgB%)�����C�Af9Z�T<;	I��I�㒆gX��~+��)���(U��Z\���;l��)���4��"ȧ���j����-8hU�c��B���%uY�5F%��v�|!oknY���EnSZ]��
�[���\���s�����3 2Kw?܅�h�g}	o�2[i=���GU��`�lKS�5��fv]�Kh%���b?����Y�4���� ��J'5�<��R�\�gCU��#������.�'
k�Ԫ��sk2�K=�/����:�a�ؠq-e�����	nh���n�	R��gFv�����1"�W�.Xi����:W���y׻Ĕ#?vFO[)���� ���A�q��!�*ǈH�	��`��sJC�)���?��T�n��;b�,b�~�*���wo��b��os�enG�wp�j�a^�*����6)<���O�����w��>|G
ɒ7R��Q��C{%ʄ�K:)�'|kG��3	&��U�?�ppQ-����{�#�ע�0+�+,�މ����'`�<G+A
8�� �G";+\�ʰ�}��<�.�d�F�[�8�D�]~@Eʥv�)����>rs:p���;�����B�ֻv��qt�`�_֒����j<�%�,C@�@�0�d;�~x��]�:1v�]p�z��+��z����M_����~<�`]2*�F��ç��>�r�C��E���%^
@���|A����5F=+��sXj�w-����!A\,i��.��k��q̤��m�s��TM͠o��z��2/bđ{|��(2l�*��m�Ѐ2�A�?��>��jG�f��.�k� _Cg�҂�Tc�u��wG�ٜL�q0����bB!������TH��§�}ƐŠj����m�G!(eof/gT�ws�rܶ���X�G*x�`ꨓy���)W�e�]̩��V�MU��K�M}�����i�+�v���-��o�(�3��Hb�ZC�C��,G��
%�Y����%���
�0=��b�>�ǋ{t`Q�S鼲�����0��\y��M��/@��(�6�J��߼L�	a��6N/��-j���w�Q�M����s[�����MTc?1�d�B����y*[(��G w�pd���
nc��Z�ˮ��eNtu��=_N�~)wXprӒ�Þ���_a8$���ë[^F=�=5�1����� ���_-�G�/D���%�;{G�%$r��E�V�۠A�i�g=�34`���<�DZ�$�8�{�3�P�p����~�)ǹu�� �RL��32"������t4����9gqT�l�?a�*ZO��s�A"�MX@t�v�VJ7X[�}3<�uɘ/U�Aqn0���6��ϒ9D��E��NG�>k)�p����1(��G�5Dm�km>��,r/���C[64�(�|{M\t�A&���D�c�A����e�w��ʓUƉ�}��8P�����A�<v�)���DY�r�iT�Z�j�G�;���u��W�<�p�]�/��4\VӁ>H�t$	H�=�+_<��Xሐh� �@���ϖ�R���	�	߽xN�ֈۈ�iZ
[��;䏑���:�{[콨&�A�a7���I(�v�9�a��h���5*���D½���� 
�c�y徨�������J1PE+=������v.D��#��Zl
��.�7�Jy�l����\�M��ٹ�c �ź�7�,8T���q(&q�Ŀ2����eHI��6"�t���4 _o/qt� ��+C�a^K�UnL�eA�����˧���/���XM�6��.KS�Iпr�Gy\/�%V��f���X�HQ}1�r꼪�I����l�}�%I�5�p���3�������]n��oB�4ܻο/����c���-�$w��6��nfQh��%?��J;�P�}�u�!7��A�}�L�fx��g�2�yt��`C��u*s5��
\�l��fN�K�n�x�j\�&�_�4�'a��+��,�8N �qP��2w�+�3�����A��pvR�
�6*�H���-����Rۗl_���^3��g�.!�	gO`�gfX,�;�=�|t2��cSIg�6�l�q~�(���-�A��yt"C�����]�Î�sa=/���A��Z����Zܒ����c��������c��&��0��(�%���3�)1�L�Nm<��,0���p6rZ+(��Mw�����my��6}cNs,�3T溵7���T��G���{1�Pؽ3�����nL��� 3 �2�APf�_�8�x�zԕD�!��\`��r����j5����Áz�1n&�5MZz[6�렗��Ʃ����lH{f|���ݑ�V���	�"6SW���qH��kg�U�SD�1�+]��.�m��wKݔ؎�]&�d���������p"魉�s?5�T���4&]�G" �/`�.�%�7�����0O�+*�,�5�2�eD���e��7r��<��ȉ���������OP�Dc��O�53��k=�"%K��,9]��w{!�vGI�\8oƹ8�����h�+�� �59}��%<��[=�F�l8�{�],Um�!�)���<�s�+! r����D�iYK�߬�`��*��Ԫ������|Cnv��qjm�#��>��y�1d��pP���B�z���;�ᑼ$~��]`/F���r�ƹ�u����׋���
�����#Δ��F+9&+���X�TcwI�C��s�A
G�k�=����_L�¬mRkx��2�����(�w2�`0��H������c
mV�2�t�?�2:>Nc�GQ��\���}�_�{*y @� �TQ��u^Q�GF��L�Z��B|�nz!gV��-�qT���p�d��n��� ���`(�<!��f]�n�e6r��!��2�u.��Nt�'[1�u�"ߓ��K�|���!�|~��8Mk�;j������/�q��-��ݚ��X����b
)C9���z����Gsm�����2�0k�cb���9��t�z��<���ݚ@��ˡ���{�
@A�މ�ÓJ��:��a�� N��-��,���w3���|�/q�[���ږB�c���d<���̴�'�F(���GN�pR����c�������Q|t#c|=���~W�p`��q/� D�af���m�]�	�=X�=c���g���4���!��5�8/��Kܓ^�{u3$`�iEG��Ic�o)�i�}9����Q*��r�c$�v	�)�0�����'~�M�߻_��P΂6r����9B��˶)��r�H~��c�� � Vگx���_�y絢���$P섺�H��{7p�2MM�iP�ؿ���ɧj�'g�l��2A�J����Pj]��wf4�v��EoL ش�2��d��D�k|�W���
M�c���\��EX�Q���E�Yo*T=����G1.�>P����Z4�4ؕG�;YYV)��$�)+�%��R[30ٛ4\�XV6�x~���s��S@����� 3Q�H�z�R�-xDD����N쳑@���eza�"-J1�����{���c,�������?mo�v;3h6��e/��e�nBgK�d��. H��T�X싶9e�PxrO���c<�w@���$���Q�:e�,N0��S���-�GDؓ��\8��j8�/
NN<�:3��`K��龨3rI ���"�
 y�S��>��|��uMhi��Ξ��!�ͦ� :�����C28�P��uu�V:��GE˦FT�O9���<�P�g������l�f\>�}�QO���TB�C�蒆�b��)�v}�!�4\x�������1�͆>ڶ�5��E)�{n�N��bP�z(1�s|��gǶ��ߛ��������Ќӱ��Mdq)���OU4~%;�dtAA	~�\5CM�� qzj[��K��~�-pz������V���B�)Y8Cj�j�)��3�X|	�6�!�Ľ{ �XP8���m�h� 	���H�DG�gR<������i��IV��H5�/�wH�=�������p�c���dݭk<�?l�>S!,���0V�O��vx\�9�k�#��˙��j�|=�<E()���sx���Ou�
�Ei��������+�E;�
�|��7!���HU���>�	7�3���x�As,��M5����$�-�q?(��p��D����.",�~�џ����,8���������=���s�>NJ�q�Jݕ�u�'��$��J�kZ���*m��>��@f�m�6�6�8X�C%�����4��W��U�@�,���Яr�p���:�c�?r����r�-�[}~1����� K:*$џt�Ld�t�S<����뭇�Җ��i��`���a�h"�wq����9�#A&��+0�}V6O�	a^e"�[s��߬%g�� �4�Z)�)��]�}�r,��c4R��F�C;p4w�zVm*5�,ޮ\�ް�6�)�(���M���-)
K#ł�?c�l>���7��T Ƕ������g�P�1��y��=���3.U��/!�������Ö�!��E`Dn��jc����(�<n�ӗM�6͑�V(�B���OZ{Tij�Ih-�ė��7��6Auk�H*�g�]�A?�1V�w�5�����eX����]�������o�εd��"W����� �$ˌ]?��".��/N�.z�7����D�����O��2���Q�`�D��Rez��7��;<ꬮ��pJȤVyQ��}ݡDQ	�|�!�u�%���K��=���O���WV�jG���b�M��$M�-���g��M^�g'����(�x'�zs���Yp��f=�����Ź#C�����i�q���,��g� R���3�cI�LL���2×U��nU\�|)� �jRp��}��d������C�V*��I�Ϥ�����HF0u;�yV�:8e�(�7QA&>ǀ�n��VXgW�ky]T	�=,Kcz�2�0S�rT�(8���;V�D>7�|` %�&�S_C[f`�1�e�b��~_�8�GNe�d3��`����I}����Iɗ��� �f��!]����u��v�g�U�w,6�o�:�L=�ҹ\a��c�u���:+�&G�n�F!mOk��(�ᠭgZ�c��rI\��M}�QO~��TKLC��r�RH)c�(��J\!d�PEz��͏�!�ķ+>�),8nb6���z�t�\90��?��pc����ȁ��� *�y���}��MɈ�M�U]2�nR��k�N��/'�Y5��)�j���K���ݖ+��u�����d��ul�P�8L�j���|j?|r��(���fN3�!x��w��q�v	�H)%��p�R��ĈW�i���V���5�f��`&����oy��d�c[�N�-w�k%��l�D�|RM��0��O��x��T���k��������I|�*�E�����0�xF�����
��ei���	���3E���
0{�����_��/���,�g�7e�L�g鱃��d,Vj�M�����$BMqh���ܪ���,R�O�,`���h鷾�<{��X��vD�>���4P}>׳�U�J����^�L��憯�k���l_>�e!��WtZ�6\��ZX�%$�Q����&�������z�2r����%�:]Se]ǭ!��rZ�tM~��q���<�:S6>��]�L�;o�܉̔��3�J�����t��;�x�a���"J>I��~�9��$&��lOgLajP=����3J8����;��<�:�RN�ӳu_ �R0xHo�y�:��;���� *��B0Lm�,4RV��H�_�m����
�9�c�����E������0���u�����'p�����-��@���w�S_@^��r� ���"��mA���0�ɸpފ���^�|�A���)Mmi8hV�kE��B����j�� �����!i��8��Vf�;4h��j6��)IQ��v���z(
�����̴o�}�+-�t~IC��˿�+��{)�������H^�m}��2.�9?PW9>��G������Y�~Y�_a��؄�pʕT�>%u�s�G�d�L�X��'��؀H!�~�❶$Ts������[Ow�>׮R��${!-f�*i�ժTr��_��?1��a���������������q�������=��l�M�$�����GPg%�Y��-�2�J�?'bz5C�A�����Hv��7�����00�\JbZo�ǩ��t>Ӥs��$-�
گ�E�x�����@�o���J�k��S�a&`N+-��)w�	S�+��Ο��[��k��[c��d���R�I�� u(�Y�G�l@p�*$�߱cnU�=`<�V��t�-�==r~�*�p��K���p a�vx��w]�y�=�V�ӌ�M��Ӵ�t%�Yp�ʥ�/b�L�W�{�$Ю�E�������i
d�Q"[������GP$R��ə��.�j�kV@~J!�+�R����6��HÄ~*B�#��&����[*~UO�c�Ðp����@�9��yWh=�_�P\��B%����������/i@�-�EjI����ur2�W�����yj��rw�8�v(�O� H��2a�"��LkD9���_q��~s�ӻ�b�����\����b fY�2��늌i�1�B���5�))c�t�G$fuYơM��7�+�P�o5g3�	$4�����b����]\����@!s	�+4@3�0r�ꥰ����D��rx�N\@��Oe��CҒ=��i���%! ����|�|\m�Z�"27����lVo^��C�[1p.�"�b-�����Y�Z�+�0�����H��M:��@���3O��Ŭ����J���&�73����I��M�J]6WL$�V=�B_#�h�qQ����w�,<$������lU�*�噑_�M�d�`���cT9���G�l�����[��<���O�ʷ'�9�E(~n_)�s�A���I�S�~��݅���9�[�>�<�� �����������e�+$V��U�j.�y� �/�E|���`�=�gz�� [�SI�H������C�]�!1�ǔ{*HK�z2$�߄Ԍ|+t���47c��z��	HM�E��[��X$2���Jb!:��f��yD��f/�E��6.�Ꮾ&��)�й�sI���7I{�YF|��.�;��@��_��È�1)b�?{��c ��͎�>��c�U�s�(�ۈT؂��?�Zcdy�f�)�L�>U��A̹q'�o&v#�/v���$�rG�]���=@�v̽<��M]�/�c�4<;X��%�T�T	(���-<���h����pw�`aۖ���Ɔ�	�֘N���h��Z�G��pk}�o63��{�{;Im����AL���d�V��A��h�U�5
,������������CFI�kj��
~�7�JQ2+Є��JJ�V����Ҏ:����F��|�JY�<����\��E��x�Cq`Ś�v�A������Qڟ(��q�=2fU֤Ey�I��S6��yP���5_O��qT�A���wC��<�f�IKzQL�J}��R�D�� �/l��X-���;�K3*WП�4����\{�%6ef��X��}�-�3�I�{E��˓]/6%)�'�P4����nRq���q������<����̸:c˦s��-��/��Uy��Q�h~�\���Ú0�+]�αĦ��jE}m�hfX�P�G�u�Y_�9���!*S�ճ�`0�\�ج%����'�wK�a�ü�����j�'n	�Ԏ]�s������=�_� ��a�L���Y��n�D�8��t�Y���2��	evv,g�'U�;�#.�x����#:�^�]\���DFv*[:[|~�c��:4|����qx����H�N��R^��x���CޣX��8�Y�UȎbp�-���b*v��ʴ���yb��oWɸn��GwT����*��(�f�<<�_�ہ&��5���wy�/|���v���sQ�ռ��_��{�).T�O a������ר?�.�Q�}�>c&#m�2�(~GTn��9ʓ!��V�Qő�W�0��M|���N5��
��bW��	q���(��&m�M�D	��OU� u'KX�\��T;���W���uFB{y���@ci�5����"y�9j�PK�l�C�3����r'�.��?�H8�ijYC�ω|�2u���Spn��D��D�>6l	r$�H�S�}��R���u�i1B�V���5kZ�������AֱycHb�PkR�:l�����V�*0l�KOX�=x���/��k+���▽u\9|���E>���<,x3Qߝ���
���i�Z�҄ث�F/EQ}C
}��z:�#^��Ha�ǽ����7r������,C:8M��GHo$զPqէ+��v�Zz���"3,M����������&�X���K:�����>$�s�_�Jg2Ӌ�J����JZk�ꛘg߷�B�D\�����LpX���%��v�ȭ�J��+p�¾�"�r��P��J�:���r<��B�r��K�T�~��1���@�e:��2��ڃLzZ��)~攢i����!��̌���٨Ƚ*��a�Y"�/����V9*)"&�t-��Q�ddOtC�a)M���37����9;5bI<�~�4j��)� 7��}c�H\���ǁ�;�1���ʟ�F_L޽��OV��PH�Q�m��7��9��u��#�R .���AB��K�[t!�&&ptE�k��+m�O��S�"g�q�!��]�0sB�Q6�A�&v��ذ�e�����K�ѡ΁����m6�iV?�~��cɼ Y����fY��N�T�%�V�<�;A4mh��ه����,�Q<&r��d�(�]'�?ٴ|�v}N�+� ӱ�1��jMB!!u���
�uH뢎_}�|BLzO0��N�W��r�
�}:o˗������~�d�xn���EW��.\8���b����1����/ds�J	㝡�����i��گ�#1ҁ�v��ba���;L�ܾV��1������a��UŹ nxQ���u0�]�e�U�m�3[&�5h=7ǉ�zԈ	68r2eSch���냪��������T��&I�@��Mr"�2�s�~�J�#2-�`���\���Ď���4P�h-�0��Z&��
ߘqg�^��=C�j&�i���2�W��M�Ske���x�sѺ�t�q�&J%g�+D8/ďW|��B�!u��s2�-�����^Y܄�Y�M��^���=�`+�s�6D��q,�����q��-�M$W]�� /��yO�'�d���\���k?�B��o�*����4���Ui�'�n�,U��yV���[>i����4!R�[���2�(��츎a���u:KM �F�f��Tk)RU���:8�x�C��E�sbXL�������3�9h�ۃ�T`�-����U俵N�������� uWz}?ْ
B)� #4~<�ѻ�z�����J���N7B�L���T
T�K�(���2��ڮ�����Y�� �%ai�\*�圉X�A��p.$�O>��L&\W�L�i�]>�q;�����cC��D����]ۢ��Zv'K�Pa�,�mZ�CE���d��e)�T~*����^�(POBUu<���&7yAi���#��D�����T1��"������x�>Ȫt���e�
c�[ȘI�R%�6��/���1�I�w���E�Ѩ'���y&q%!��0>��i�u�n�^�h���Fч�M�����	"^�] ��hJ^���CS4p�G�k\���Ypf�v�_0OuU��Eʼ̈�)ux�<w���թ����J@0A�����T��A��|��J~ Wuf�V�	9_�`0���Dp%
wu0G$�e�����l~Mi�.Z�_2dHWm��f��,!9]��ZMl�'$�}��V_�ݜ��s�'σ^9�tZ~wk�� �������Ŀ�w��s#W�D��E�� @dW�&IL� ��e,��$i$�>��.�w� ��E�+����Bf�zc+'[���y߲����l�s�j_��H���z�� *챥�pHǥı����"O�m�L�Q9��&��.��~��L'O,Ca�m��v	3�t��;�B;��u<w�<�wU�xa� ﶻ5i�H����
;����`쨍Ԟ�L�M��-6V�<HzF�m�r����l9Q����w�
�vt w���S�1��8g��`$p,׸��3�K޴�eSdЎ�)?L�'���K�	 �A�'�����)�����X��������m���V�!���L�tg����;Yȁ��ᜤ�^AV���;���h|aD�oeF��9�Q����](����煴4��}��ŤT�Zw��
��?TTe��KF�^�lwP�u�u����mhOA�J����ы+z�6��|j,�t��x����X x���{E��QڼѶ�[oe��9z%9���vg.�X��I�D0�ó��oR[�L������9Ֆ̟Bu�m^�Lp�}?��N��,͢�
��"Ŏ����Ӭ�M^��,C:��p޽�N*��6JYyg�����0v�#��Wf�����$a����u�}�/_(J�k��ְ���I󫋐�Cx�J��tW���V��#_��w�!�~wew\qd$GøÑ Gl9�����_` odoiG�����I�9͑��V(�lO�@Q`���0��g��z��'���9���~�J���7�^\;E��~\ëZI'������ ����
�_Ӈ�D�ze3K�$���m�.�j0 �6iE,d��[��2zj�e[�*�@���aXa��R�ѽ�D�'H��#z���4l��,J+$��;�a��ǹ����ԕX�)ơ��ab�:��.y���fߐ�E2��.��ُ^��I���j,s�����{��|Yz\.�<�-�@��_7{�^��)R{p�� �U��>,�~�YU��`��쀈�ɭ�<
�y����](����yU�'�|z�'[�	&&н/&�M�μ���G}�
�X-�&=N<4�]�ku/�VN4���'���	�ܷʻԻ<N�a���ΐ2�Z�a��vk�	oQENS�����Z�Q� �G��G�5:o������S��$�K��Q�GfԆ�� ��j�#����B�ߵw�����)�{_\�Hu����aHr'"7�4�9ʹ�&mUxnO$a����1�3׌��#�;զ�<_��_!`�`�\ ���1H�59�gRh;~��HCY���GL���y��V~�UHb.:m�Wx��sI99��P|���\V��~U�x�������J�p�ɢ�753�Դ�8,SL+)��$4z���7��^A����z�>�/���l���w��n�ގ�Fm���V��q��H��\�����v�A�����)$k��Ǐ�I�D>���|m	M�K�h%��/�2�E��Է���ۯQ�m��82U4Q?W�=>�dpG�S�sm����_�P�0���j�T��>u��#G}g�L)����_���)J!�e�čTz�<�����"),��!'�ل��|!M��f�8@��}r�3�J�j��VѮE�'����,�V�*�°���%S��Y�6�FMb��۷Վc�L2���-쬦��pB��^bb�C���1X��o����Oɦ�i�i�b0�K�b�2X��Vt�����¼S����F蘴N�r8>@{�[��J��Q����a�,zN���-�߹���w
,T�r$���[�.����ec�f�dS��!�����(: �G���pɞ��Բc5�8��*N�ݭ�t�=�=�#~��opׅ��ȝ�7}�a}���d.���W�=˻��-��������� �d�,@%/ɢ��J"@{@�$�g�E����*����i�����L�	��$Y��ɀS7�����Z~�Őߒֱ� 6	~ËejBj�,��~�̉��~�a�co�_��n%�I�@�By>'��&�+P������R|_��,%� '��6~c���jɃA=28��!�6�\�Aj�?yw�dgv���|�� �%62�Z&���D������Ì���_�)�̈́\��H"D�?>Y&_�Ԡp�p2�1�ݮ��P����+zVG�.Y%��#�+��ĪV��3g�40BE�O��OF1��6 �ߜ@(����3�����-�$��D6��~N�tJ@|�e�YL�Y��1��ʚ{?�{ы�}I�^}qߔOgޖ���hMb��#���>�%Z�KAs����G���Bs��8T9\s�xI�E��B҂�"��.���jK���~e���N'������"ޠu�����b�P{�F��N3��3�=X`&��^��IW6p�Yx� ������S�u�\�uy��E3��d�:+B��a�/���uG��:9��G�O�F��OO����s�8g���;D���X\��B}C��O̹NTYP�߁��9��)��\�R\� �ޛ7��=�͝ю��+?��,)h��np����i�zy���*�!����\�`���ϲ��.��G-�'�²9ܤ����~��rj��B�Tl�S3����c,�0"t׭<n ���j���!,xu��E������
�{Gy� B�%��Q���K�4Z���;e�H�%�������L��
�0��:(���Z﷕��El��ִam�zG��m�����[8]�1�?mCBr��s+Y��pF��U%�-���o�}��έơĚS6��f:_[|�\깺On=�3�� b?8xh{��	˱@[Eb���ǭ�,nl���5��v�,h;�1����$�Y�����6�.5�e��<}�8K���������$�
�'f��Ԇ]�s���a@=��T� ��a��:��H鼈J�<���O�Q�*���O���vn����k�3�.�g����:���U�J���v"eM[tf�[[�2�&��'�q�|����H�q������9h��Eޛ7�0�S�ME�bh��ږ�*n��̝��wb�koO��n���wL�����*�M��^]�<�/��y�f����ㅝwq�y|�D��n����Q���/(�ҡY)&9�G�������9?�ϛQ	DA�6"b#e�l�oPt+���,gum�e�G�$#3��]�E�8z�٣k�+8WM�@��}�)�<h4���F�9G8��Y]�%�ʁ[)!�1��vAs��x~���A���������M!`������q��XC����_�5@���ZA����1R'�p�哹��z���)]	�j_-~s�]��F�"O� �;�N���(���?D
�B�XBY�M�F��+Ek@XF�ww	��,A�P��K$a�M�K�p*;m��v���R������9�2�֑����ۆ��m{|2�c�?��>��`G��QȊ�����_����o�.A�T?��u�?G�J]L@�����ؾU�!�3��[�T����	��YS����r���ɏ! f�]|�S5�r8�
��a7���+�<:Փ��t�������(9��<3���M�M��MY\�黄�E_��F_�F-C!�p���D$b�
�C��������̧5�-�P�V��0�X�b��k���t<�1�s��&��HU�}u�6�ki�@�U���JF�(�(�raC��N��-�:�|��w�v�)<w�]W[s�D�c��dj"F��5���(��G|�*p@W1L@clIu�����y�tш=;Ƀ~�MpNuڕ|!n&a��q�[�����=�7���f=�_�5����#r/����V+{��$Ne_E�kT�a���i�϶���񿯯���$����fԶ,h'�)B�~����i�����6�v��q�B�ew�$D:̠%�~�PcF�}�n�����طy�
�]�vP;A��.�)1}��|��m1ح���k��jG^Yɚ��2/�0��K��j�-$wTpvI���3� <2�^�ȗ�D7�E�rr�}閭v|`�6�s��?-j��%Y��k�ٌ��@1�ZU�����H�"��Gbm�YĐJ�R�+������3�G�4G�m�FL�&~��[i}Ai�@����i3������y��oD�T�v�N�-@}�e(�Ґ�E1~r�rf�{����=���T����/��S�hd-Ě
Qu�`�����K��I�S^�1�y�~�*W9S�x ���j�T����n��PR����ge��N�i��X��9�um��qBq
e��,Ҝ] N*�N3w�"`��DK`Y���[I��՛�ؾ �G���b��*�Cu�?��������T�$:J�z���J&��ju�f�:У�G3DXF��O����2����gij�up���\,Bl}���O��Tp,[�������)h���Ob�\f#(5�$�0��ʹ�������)��nL��P��z�1��:�K��}?j�7��Ȇ9���>�==�bR��È-U"��ӎ^�p�o��l�'5���sNWN�jIAkKY��ݛ)���}��#��)#�R�gjC����s�6xvj��kB�����T�xQ#~���cJАF���~؏gdym���5�[P�������x���o�؅B�C�!j&�r�_2�0��V��z[jc5�w,�v!�f�L �:K2�ޗ�!�D|b�]�'�UD���+	8 Z�K���4-x�IY� QC�}���[1�h���Y��,���_G:�eY�F�*�+����3vh�4ԋ��1��d�36�Ѩ@w��A��3��������D�>~N>N�d�@Uzde "��h�61�i}�J� {��"�����l���,��ŝ��|Qh<q�����8i=����K�a=����vٿ�Q��Ʈ9+�Mx�x{�B���}���F�(�(p:���Ne��N�fj�����n�M�œI]=��^�_]�5f$N��3O�i`��_#�Ϩ��I��ɛha, ������u�t¶�c��Wq�,��:"����[����h�u��:��8GgF��O^���
y~_�gA�i�Ze�r��\�-}r��O��TH�ء�����p)@5a�':�\>����#͌��a�{y�)��n�{`�(6z��o��<��߶U �>��^&)������:0s������U�$�����HԘG��Dz^5�&�K?�&�-j!��K1)E�s����Ư�Vk�^�K�o�8I��j���Ϲ�|O���%ă���nݷ����nY�	��8HI6đ�%!RB8Nĥ�@ia	PV�[5��x=�d����L����2cx�H��G�k�kl�8pƢ@��0��6O�<�x��D_��k[���˕���u�|���En�m�6xc�"��+k
�̖i�=�Ҵ!��1�E��R
����S��w���v�g|7���D_��G�,s˗M���>��$��qQP�F���/���}�,}�x�%ۆ�;f(����k��{9��)>T?^�7P�J�+�ӻ�G��H�LS�k��I|w�����t<N��'�|�X��%���K`.����[����tRk�r�������o+o��KW�E�C��}"�<+9*΄GFq{@8�`{]���$~�)$&��!�sY����N�Į׹�6�Z9�����`�E���z���6��$.Cǽ�B�L�V����伺�1�8�p�#�*�fzddG�h_���D~�£]��F�楧�"k�q����!R��}\
�b���x�P��F|"�+ωXi։w�w:���_A��[�|������3�m���3���d��Z�2������g�:�I9�m���2ojg?��>?��Gb�Sȍ ��_��_b2�
� ���T"��uO�_GWY�LC�I�0L؁H!���޷T�*��a�"��TE���e�3��R�!'�f�P�6�2r{ ��$Vw��wj���䓘�y�nv�D��Щ2����|�P�M��k��X�h`CfʷB��-��f��J� t�b[C�����v���@�� ����C��   �  �    �  b+  �3  �>  �I  �O  <V  �\  �b  +i  oo  �u  �{  6�  z�  ��  ��  <�  ~�  ��  �  [�  �  A�  ��  ��  �  V�  ��  y�  R�  � �
 O  Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�� |d��"O
`�(�;���8���-0��1%"Oj4��ND^[��"3/9�0|H�"OB���H��*�ʞRy=a"O�味V�!X��!&F�:J�$���"O,��a
���C�Ą�M�"O,$3%o�-���p���+Ն�:1"O��ݢ1����`���y14]2��i�<�6��{_���c�H�`�fX�$Kn�<��A̼VI�xR[�)�Ć�pඤ�ȓA5��('nߡ4�� �)˩%� ���,��r�؊b#`T�eT09���ȓ!�b��g��}�8�F��-? �ȓ
K|m�ș�VṔ���2�%�ȓ"R�X�j�4JN�1�˘X�i����̹	_�jZ��1!g��zܶ��ȓgil,*�J�
j�Ne��i�J%b���f	�(U��:���G��$Y^م�~r�� S�%T"���k\�jx�ȓ|4�1�îJb��@ӵ�ݩn�V��/[`�"�v4�R�!ʎ<��M�ȓ`:��z�ؚh�J�Z��$HY:	��H��p�m�C1��!��B:��0��EnjZA V;9����J[
2���	��4'J�EA�IVW&��~�(aZ��ӹ�>� o�Y�|�ȓ�f�A�
Ο7�H��M�$�����mޠP����/���ANXo*�ȓTv�����{ ��-7�*h��I��sB�8�8���3����ȓNe*M�悡;������X�o��!�ȓ'lj�#F�m�+R&;�|��2)n�C��0S4���T:
b���:�0!��e֊��)��ͷV��,�ȓ0�&�8#���� ع�L�����;�P�AFd���,w�6d��r�EQ�( �gVlɦ�M,H��,DP���|�I	$G#\���ȓ"�)���E�B	yt&B�^�LɅ�4�� ��eC�F�ڙ��n��R�p�'�a~r��I`e��Qk�Mq�C1��>�M��j�jG';���@���}�>���*D��R&�! |��&�I4wAzׇ)򓳨�p�x%�	2�@�{ģ��M|.E*F"O�m[�FƩS��A�-�<Zq�m*�O������$Ya��І�P%��i�g%�06.C�	�KҔ�B��*ڱXa�%�C�Ʉ\��1(ɸ��s��&��B��0\�&���+4H�KC���/x�'4a}R
<Q��ip�-X#!��=q�E��p?qu�}��e���0%�4+`.�#>��@�r�%T��3�JR�C~�X[A���2E�$�R"OV��l>_���å�Y/C�Ѫ�"O��ƈ��a���Ǆ5#<���"O(eӐ`��f��3�f�F�L�c"O�Ȗ�F�
;L{>;`̩�!� 4�й��ķ��T��܂9ن�H�*D��S���2_�Q��q�X���'D�@)!� J��Py�*Ç\�0�J�.3�IG���>S,M����tD��q��
2l���re�`*�)7�D�E�Ģp.��}rn�\���&��/�,��L���p?	�O� �}:iI�Y�t����ҕ�H��"O�L�r�O�x��8�u��l���(d�D�>�'�\�O��i�����ҧ�*����$>�!��	F��:&*R�7�^��k_�j"��!���,�~&��s�/��@u�T?4E��Ы5D�[� ?�T�*��� 2��C�-6}�)�O��ږ�:3��JD���)�V�Sp�'�\���M�y��2tnD<�!!�2i��U�ȓ�b�Z`n�<t�����U'���ȓg���riGd�^�F`�V6���Q.�"G��!�@Q(2��d��m���hO�>:AmB�������0�㰧4D�����ŋx0�I�7u{���3D�<s˜�{�f5��!���)0�O��I�6T���@_8)�����߱W>�B�'@����,��UM���GݮPzB�I}�~ș�F�	q�Y����C�^B�	�MT��*r�0p�-h�b�!
x�B�I�z������]�w�dB�	t��)�����r��G�Z(�tC䉹l���#���)!��S�+؀:_�B�ɳsk���c!´>*�Y��B�'�B�	�O����f�A.Ʈ-���_ƬC�?���BΰQW���f��eQ�C䉬B�!�e�ؖ^�xQ��"�C䉣)��s�ϙ7S8aP��"W�l����O
c`E��@^���(9G⌉��3D�����^I[���Ȟ�|��B#�2D��Г
.���a�N�+bƴT�ì+D�4�QEVm��5
O�z��8a��<���S+[�8Y���iu��#/�(��C�I�q�a#�K�&A����J�=[�C��$[^|0Z@�1[L�P��gZ3&�`B��(Lҁ�B���)�v�����JlC�I)Jl�K��6d����1�dC�I��|p�VD��R�i���Q�ZC�IJRi#v�ɉa�I�5D�n�dB�!�&�bbI� ^������DB��=v ^�E	��Bx��H�@��:���g��[
!�OY �8A�ȓ@��t�ȹ_�n�iC���s��i�ȓ������]�dAR���$��q��	�"��IҀ�3��MC	Z����R�h�Ƈ'|���sU��N�І��Y}��!h�BJt�U>�ɓ.%�y�]�b����Ԝ��p�ӆ�3�y�ᘐ��\Z�ǚ��@�z�BO��yҥ1�bPp��I��|	�ȥ�?�M2�S�Ob�h�4�D@\x���pFV)��"O�d�R�Zҵa�M�a2�|��Y�d��I�b��$D��.�ډ{��Ŋ2�'?�x☟��P �48t����-CF@ 遃<D��7V�G�Hx�kG� eJ僶I?D��A*	�b�Z��LR	a]��c �7���(���/[�ܛ���c�칙f�i�ў"~n�=�,�c6��Z *�	@����$�>Ɉ�ɇ.�
\JT�	 	��b��֢8���I���)�.5q����9�	i��??����d�
��-!*��	v%;^��}Ro�<9��s�|P MH
5�By'
U��I��eXQ�˫I	\�As"R�2|�h��IA≡s��Rg�нK�������$xs���;�S�O~X�پ�<�C*Z�n]h����	k>�J�'�
�^%r�T�/�^x�Χ>Y�S�? b����z¸��c4:&dL�pQ��'���?�N?�@Fn�d�xS��l�&��W4�OvO�]�p�< �L�ÆKL_��E	e����RGA�!3ء�-��M�*�i�$S��y���J�jU���ΒQ�N�ط�y҉U{�1�nOD>�0h�AK���'nў��OT@c�A�<5�:���'�
�n��'�q�@@��7�H�s(�[U|�����|�"���.����B�^(��	ҧ3_�d�ȓ1
P�8�@I/�,���j�>��>!�*RQ���'�J�����Z�.Lz3 m�Q�'��y�s �R�Ĥ��b�+8d�������'Sax"�ߑD��ʠ��0q����;��;�S�ON� ����D�'��#�P�	�'�P�!�%qܫe��J�<�	�'����'%։g<�u�TEKޮ�0
�'�\���� .E\��J�8E]��	�'�Hl��ɨyW�x"s��pT��'���D@P�3���אQN�b�'��J��!u�P]�#�Ҫ�
�'��}Э��jȳ��;g���;�'J�B�
zb�RU덝NP1�'Q��HX�>.�$kq��?0l��
�'��i�En<69�Í"O2h�	�'{�a�w� �)\���/L"�x��'I� сF8� aa�J�v�h�!
�'e��ȄA�>T�H��T&vwy�'@.ayd�?��e	�i�J)�'y`���7rRa�D�߾s�"E��'�l!��;O�T T��h��D��'�ؤⓨB�x�+^ӐI�'�ֹQ�u=$�s�G�T㴽�'/ B� V�S�<��f�+^��@�'�@�B�� 6�T�F�Y'^<�(�
�'�(��1*���ZС�eZ�Y�µI�'��yt�)2����&��9[z��'���:T����Tŀ��I�Y�<q��'�n-R�ADZER����;Q�d�	�'*
�
��LQ�PMc"K�:����'��ڒ��?�tK��F�|���'�< ���J8o�`�순g�ma�'����7���R��Y`a@3t��`�'�n�ҵ���c�l%��/�>&e��'Վy�r�7A2�<9��҇B��hS�'lp��dø$^�u�����u���
�'[�5�fI	e���c���O�*y�
�'�z�����[_|��S��W+4��'��P`�@�v���CdmU	Y��8;�'�ya7���g�0�C��~���y�'\��Ī	o��iARG8�ԬJ�'���"�����L�f��'����H�kW��8C�#tDܑ��'�����e��j�P:��#Z����'rL��%�:������X�[\`�9�'J��pr��P=\BbO\�NF �'��+�bR�[����qa\�HFy#�'8@�PsB�S�(�p1(��L�X���K���愝>F) )4ǉU�����ru,�DH� (�;�A?m
�ȓ(Ē��E�'#pQ���?|r���a8�5!E��zR4YDP:*L�܄ȓi(`t`N�8!,�����[�$��ȓrH<۰���%�"	�ύ�'	q�ȓL-��6i9B�C'�^�*
���S�? ����*#��0�o�7A��0��"O�]����>Ü�Ã�K�oq�2"O���ञ(�8�メR�&��X�"O<]���;/C�q� ����M �"O���G	��lҗQ�{Ϊ�;�'���'���'`B�'"�'���'ܮ1��*V�D��$�ض:�����'9��'�R�'UR�'��'���'N���׈��qd �F!��'�B�'ar�'gb�'	��'�2�'����+�z��-kpǇY��-h'�'��'l��'���'���'��'��h���)(�,[/(:�*#�'�'��'�2�'r�',��'���d�^4ز��m%�!���'"�'�"�'B�'��'���'ld�Ї��-��I[���_�V��'��'#B�'X"�'���'�R�'�6Y)��@9��d��̋��з�'���'J2�'L�'�r��Uݴ�?Y$�s�0�xdu'J�xe'�&�?���?���?����?���?)��?��l�O0�Ai������!ؾ�?	��?���?��?����?����?y�@�%>��ܢҨ(Q�Ah�D>�?���?���?)��?��?9��?i��Āj���8a
Ƿc����T���?Q��?���?a���?����?����?!&�)N}})W�A/:*dҖ���?��?)���?1��?���@;���'��|j<+f�F!cV%a��\˓�?Q-O1��I��M�b\��������j��0�2�)0����'`7��OO��O�DP�d�L�"q��q���w��V17��O��r6�#��I'SrF�gȖ'E�'N���&Q�����iFb$�<�����?ڧg�0B��H�����2
l�ƻis�=��y��OB�O�r6=�\- 4�(LXR�xRX����1Õ�n�<+O�O�01�����y��P	,"������e�t�K����y��	�{jƴ��ǵD*ў�۟��Q�	�R��B�^::�H piy���'��'4�6��1OX�7��9e�)�C
  �����OؓO�'���iE�d�> ��=� �BkG�C�V���Rb~�:LhR5đ)˘OG@p�wDQ%K�iBn,|�@�]p���{@�����IiyR�����d��,U��qp%Ջд8�	9V���ʦaz�J:?)սi���|�O���#$�ΉK�2�F��q	��+�'t��i��i�#1u����Ot��E���v0(a�F�=�""ٓ���JǰA/�uxPiļ
QL��b�%�L|�4�BlL?�a-H.}W�.�E3L��J�p�x�R�l�?s�!�Z�s-�9�u�R�]��ْ�/#�]a� ^��B�h�'���� �|���4n� N�^0�	�%7 ½��a	�5���)�;g�ݠ��C>%�n ��o#2�Z���@@���j�о�BB,�-K3�}�E�F41��yA��ar��>
YT�B��f���� }6�	�M�"�V�'���'�Ī ?	� �l�|�`(ͅ7D�c���%�Iٟ�p�Cyʟ��)�O���!<���3����1�D�AڇLR7�o�1l�şD�Iԟ�������|������MZ�@����J�W����ʪ_��	����I�?��?)���ԕY�O�.ܦ��bj��
�&���i���'Y�c�zO�	�O�$�>	@���>
|JŻ�%�e�'�B�'���O���O�$�OBkE-Q+2����Û g�=��o��5�I��X�H<�'�?����Q+S�BuCgbѼ0 ��S�aV���l�\@P�$?����?���?�-���ؖ�X�|K�(і�_1�h���~9X�'��������	\y��'����Q��eBQ9(jq8�
�*6�q��yR�'b�''�0R���{�O���!��P-�� �\iI���Ob���O����<����?��x��KƠ5nU���
e���rMP�����O����O��D�O�5��oX���	ޟ(Z��7�n�(V��%T%�)Hb�<�M��?������O|� 6���'A�ͺ�b��I�x���h�Qxz�4�?���?)�[�̸�B�i�'-��O��m���>�"Iz�C�*���k'u����<���#����'�?���H�����׳V�$(3v�դa3ؔ��`ӂ���O�p�5m�ۦM�I����?�������ӊ$��Hr6��I�)��ң��d�OL���k�O�O�i)��$���H�R&&�,�:�"��
�M#)-ɛ6�'��'����OR��'+� &�T���D�JF�Ѓ�\�V>�7����D�O��$،��I=�����9C�R��H��ť�HI���v��I�	럔�ɀf��|�ݴ�?���?���?��pt B!Q�x$�o&_�M�'��>'����|*���?��\�pP�F	�tZ<)
��H(5I�`�i�RHM.M�P7-�O��$�O��$j���O|I�H�6T,����L+���W�����=���@��Ɵ\�Iן�:W��^-���n
)�x���.2����4�?	���?)�w���OyB�'gL�:i!j	�����<�F���y�P���şL��$�	��q�ڴHc��I�7S�)[J\�%���i�b�'���'?�Q�,�	����SMEA���	x��Q�4�Mb��d��4�?����?I��?�����㡹i`�'[>����:\$�iP�%H�k��yӞ�D�O>�D�<q�H�& �,O���Xs��y�ʛ�0��� խ��{x7M�O���O���	�>�6Em����	�����)K���S�q58c���b�p)�ݴ�?*O>�$�����O��|n:� ���v�G3IE���#eY<|��S�i�2�'Rx��%w����O0���@���O@�a��HU�T2F��k���JRkm}r�'��qT�4��'_����� .(&!*�-J+M�!b�4������i���'�b�O-�b���NC��!D#�0��-��	��M�%��+�?!N>����'n݀�g�	v���
�>���,v�b�d�O��D� jqf�&�|��ȟ���w��iҠ5'� �3c*%�l^��'��)*���?1�?f�aR�éxR���q���4�Lx���iI҈R�y��O����O��Ok��t,���2�����P3��y��ɓW6��Zy��'j�TO]1i��"��}yXA���`v��fd)���O.��*���O,�D�/or��c.�������\xSd0O\ʓ�?���?y)O���!�X�|Z����t;��f�n��E0� Jv}��'Y�|��'X"j��P�D��hl =�"#Ƚcߐip�"U��	ԟ��	ҟ��'I�9��;���+`�B҉���� e��7sҘn�şp'����ş`F-i��O��)��¦� M%!�[\�u���ir�'��	�,z�4CK|��������N�|I��!�s��T�����'�"�'Ȇ���'<ɧ�)NaT\XSԯ	��2���
��6\��{ָ�Mc�Y?-���?m��O6}�cNO�9U���L�%�J�F�iv"�'��˟'��'Zq�.��u�T0GG\�ՋM��n�*�i��ƅh�F���O�����H%�����[(�T�3�x�ID���Z��4Z,ft	����S�O ҁ:&.z� ��U�(!���!\�6��O~�D�O ���\�	ȟ���y?����%h��}��)����G��ۦ�'��]�JO��4�$�O����b4�5q'ĺw�����bb~6��Ox�k��O|�I͟t��[�i�ى�a��є,ӱ�Zv�Ɂ��>��E�<����?����?I���iV��l��7$C�g��J�Gķ�,���	Z�Iɟ���W�	ɟ��I�#���Rǉ���܂��6Q>,C�O�\�'���'�bQ���������Th�5�d�6O�HvvUjA.N����O���0���O���Fab^�D���Ji��':�N	23�W�Rx���'��'��]���`ؓ��'S�uX#j�T�`4Ke%1K�����i
��|��'�$R�b�2�>�d��d%�< 6�'�ڕ�#�YҦ���ݟ��'|��!�i�OT�	�kF�E`�����.����ޱR5X�$�X����8XY���	e�~�P��"C~�5H8J���WU2���'<>uQBcآ&�&��O�aH�d��A���~V�1"O^�!Pkنbi� z�T�tA�dy �T���-���L�]u`5��eO�`U)q	�pO�T;��Q�`i�����S��eZg�C-�b�1!�A2K^�Or�԰��+l$r@��C.�����H 1u�I"�� 	%	L��h��SJ"� hŞyL��d�4P`�ڐ��p$���iJ�;��O��d�O(�$�캋��?���bcb 	��I�~"hӶ��)؛Vꋗ.<�0�"CI�����O3��@raDL��&�1T�حV�|�0S��*D�����i�r�K�=	���Η���TE�0bӠP�<�Rʉ{��A�Խ�y��$�U?��ƟT�	A�'��,|[>X��'R	o�)Ѐ^�; �B䉦-�~���Q��!��eB7'Z�!���?��'s4I�i{�����
?ͅ:�|y
%�	F�����O����O���K�O��de>9sf �F�(��BLb�X�0!�	86��=I'	��>�A�KRx�|0S ČH��M@d�US� lӇ��1����&N$���(%/}���F��/o�TLe���H\��'��Z�2�I��G;�n��,S:R�ўtGҊנ�ȡ�u�2�]�_�\@���\�	Č��Od��ÌS�`��?3��Zy�ō�tf듲?+�J�9�f�.��<�ƃ!0m�(��%Ydc���O��䌦/@Y15�C7�*��� B��ʧZ%��*P�n4���@F�1Ey��nJrR3\U.Y�p���M�>`�|�K�B�"|�h�m��(OHx��'�"��[����͌�{V�;�(�I.�d/�O<�C!oV<WB�s�@M-u��,�a�'��O~��Iq̲,���O�rQ��ȵ;O�(�+���������O��Q� �'���'G`���
?�2a�����se\�{�B`���#2����V
W�O�� k��	^x�飆�f�^����2_SRYAVc��J�����H*�~�d	d`�Y�|������e�M�8��U��:8��I����4V����'J?���:5������(��,�Р#=�d�O�����D��b�'V�Pp�&a*qL1O\���U�'XP�bB�'����	�y�0���6F�("�'�"I)-�@�*��'��'��$l��	Ɵ�kA��,���-J&qaxc�� tb8aU&�`La3�ܛ7���3�To�m�4o��B�Z�� U���XI��&��+��T(D�)B.�L
�!��g�0�$��[��f����%gߚGBu��K��<k��O���+��O��D�<aW��mO#�E�\�����
��Γ9�Z�{�Ԏ3gD��Ϙ'��c�Q4�]��G-;z�r�AR�L�~�D�$��T�'H�S&.�ݴzb���(T�B0�h���L�5K������?a���?9����?����D��*P�����GW�? �`��B�N�r|
$*����BM�A��y��J{�'Tj �q"\̍b�%��5c:Pb h�we���f

Z|Ay0�M�1�Lq�'�O ����'��旵(Fu��C�o3l=ZW�œ��';��'��O��Z�ܢF�	>B~����E����$6ړR����'I.�~Ia!�NyJ<Γ����'i�ɲQ{= ܴ�?1����I��H�i���D��A*4�A#��ؐRd�O
���O8(KN��eRɠW%]y*�&� C$}|,�A)B�2݀%���j�jI�I��~*��O�n�3��\�_ ٣E�W�'W,|	��e�>�h *x��QfiN�V����Ԋ?D���5L� ��	CT@�I���!�=�OD�%�,� A]�ke�aI����{�|�����M��?A,��QI\�?����?�G��wD��$L�b���B�?s���XDDFf&�R���BN`(:�X?��|�]�b�`p n�1�肕Pƅ��������H�n`"���h���٪KE���j�mu�0O^�6o����'���O?��ߌ�|9��A<)Mq�@/m!�^�Vn���fT�3"4�Q5��[�Dy���?=jd�*j/8Y�!bR��� k��H��	 �~�ȃ	��|���@�I6�u���y�nV�s*��{2E�X�Y2���?���Y����:������-'�Z���hOJ��� '����2��)	.18iI':�ZAqrH�-���D^�5��	J�p"�Ԙ#�"���1.�ݺ�%S*&m 1�����-�"�'�ў��'~����ΣDNt��n��$�S
�'U�OV"(����&�>�����S��"=ͧ�?�+O���R.G�Փ�j�	�<$�P刕b��QTi����	ٟ��z�����؟�'KzZe��Ț&�����$"�و��@�7X`!��o�*!]���3,Ox�v�_�y�H��f�^}v��;�F�M��$K�`�Al��L�d�'ON{�'��i���~��V|ݘ�2�'ȅ}(P�x�K��T�j7�9�I��H���F�E&p��/ϩ1�&�Kuj�1H!��@x�l���Y�C��a�v�7o*�^�9�IlyҀ�T�J��?!,�bI(4��!:�B`m�bn��i��1u^���O���͉~�R֠FE +c�E˟�'h�DYD�P�C+��Q���LXP1Dy�Aۘ'���~!��1��ˡ�0�h�B:$��c ŗO��T�r�@�C�$�q�c~Rŀ�?9ѳib6��O�˧s`��iK v������}�(����������DR�����4b8�	c�K�X�a|2�2��ˤ]$<H��+�0�w�C�/����� ��Yx�����.Ml85���)�̑aF`"D��Yk���Hց�����	+D�����> �\��W�\#��r�*D��P)�TYX�B�$/=�8a#D��P4fXFx:���A�G �XQ�>D��h�D�_z�Mv/�L-x��F2D�,�g�Q5c����nU26�����2D�pRA#Z�d�|�÷R�!+�[�b1D�xP�h�3n���PDN;fd�X	��/D������_��Y�Ť��s[(�ٱ�)D� 9��f�h�YVD<))҅�B�3D��:�ڤr�r��D������e1D�������J&4��f�Z�;<���FD3D����b\�W[r�x�/��K����1D�<�ˆ�1HU��C �pYf=D��p��I:-�4������J�႗�(D����]�c8�����d �0)b�$D�DcA��!tM��w�,z��?D���I�5s��D�f$�`�|d�V!=D����ѬS�|Be�+su��[!�:D��x��W�5nԨ�O��}/\y��@8D��0��#�!� /w���6�4D�k�� p�1 ��׉;M��'8D��J֩xK�uccԁgCc�h D�08"G�ўDc.V�m2��p��?D�,	R�@��bB���N�����C D��z�A��\����v��t�}��*D�`���P�JT��F�0<���*D��ȓ!��9�¤OJ�P�j Ad&D��c��A�%� �$/[�CXC��%D�� �d(q�ҍ&���2���+��+Q"O 0���-�ZD�s+Y�C�25ʅ�	&H�L7�۶��Ż���d�Z�O������~�&u������yr�P�8�@�ږ��~�:��3��M��	�[���gF'?�� �S��M�)ѽ{5N)(��&�^����D��L�!��1pb!D��`?�1IE�^�' ��'�4�u�Y
Bt<[�߸C8�F{r�C�bM���'fS�#Pk���O�9:c�e�80�����1��i����߇V�:�)W�ߤ��}�qG�
<��|j��3�O�5x�`�SL�|��N>�r���S��`���7R�誐��\Q�s��&�~��
N#�,�wHԠ!$�x����K�<!����Di�W��((�ސr�*�M��m|�<$�h��F@���#�T��\� � ~������%��B�	%Ss9����(B0���:Ұ��v|�Ј&�kOz͢'[ʦ�q���?O�\�$� y��E�	���*�D4��P��ɍn�|I�Fe�@Q� 5d x��jK�Z�T5���Q#=-�C��<����'�Rl�U㉊�OF��'�ޖ�����h`�@����!�?Q,�*�dèq|D���J,?�)O�q���xelD��C��|���q(=Q�Y�S�V�;�a|"'C�v��TZ��ƕNR�Pm���MѦ��
�\ٺ֑��ˌ�4�&�+�0GyiP�2) v�'�&�)��Aq8��{����l�nx@��ֵ2��$/���U}�/�#|M�d�s���uWE�hbpm�f�ҋu���Yi�y�C($�^����ȴNH�I�@ƃ=�M�b� 8RVA�f��u2��0`+8s��'=O��S#+X:A����7/�V@�b��P��l����!eR�Pc��
�u��=(��
L��|���O�m1�&J��@P�'{t�3�F_��`��$����vJQ)���#x�`t����&(6d�b㘟���=?)A�̆�p�O�~�]�o����$	��q����'TB���Z�z_9h���$�����?H��իUe}�gH8=��d�M?9+�G�k��ѢB��MG.��I�P���ϞjD�����NA�'��M�ʇ�W��U!�'�
�!۴>���CRX�ib��C����:����'���sI�?~꽰֮�?o�U���<Y����0 �?+n��b�ǁ�B}�ɤA`�XsW�i�7��ɸ�O4�i��mZ�?�.��`p����M�6�e����Z ���	7LO�^��&��l̾6H8�˞�zK�� ��⟜͓�M;t>O���WHM~�����h֪y�fQa�(	�R#����3V�10��<u&���Ԋ��W���2G��n��5O�O6���[#aZ��ă_ӆ�j՘>Y�-�N*ܴ3����TN����"TO~b"]	)��ScKu�D��A���ē��imZ�5j�R1�\9imq��	�5�p�X���	U�Ȕ���P1Gٞ�Y 'O�2QȘ%&v"��'"	�c$�}����<af/�?��'�
�X�O�A0c
Q�a����w���<��H�`$s&�~���z\�R����X�
�}KV���2�L�B1L�<AK<�� ��ٳl�UWz]3��o�� 2�Ğ=HV����m8�� ��\$R����ByC.�;uw
�C'�O�}H�����7�?QK<Q���/�¤z��^!=h$��G��'�pYg���S�.p�dY�j��0�O<\��-ؒU ��5v�v�x��H�?A�Tl�83-������!;+��K�&$EV�1׊�O����͜d���D�?�Y��ʜ�5)2�R�F�b7$�D|�/�O\�1�.�<��'W��HC���4 `�Ġ&´�u���p?��=/hj,�t圙~�"�j!!T�/��ɲ
�2"R�V�B��ݦ�֧�)Z�W��xCW+X�(�DѴ��0A!�C�Y@�x�iG�9z��<�'Q��'��s��1@�]���ѝ'�}3�'x��H@���h���E|�˒�j<*A�P�*,�L�!A������
UXa��K�0����
��~R=O�)�Ŧ	����EQ���W	�D�pW!��oQYY�'�TA2P+ ���BQo�4@���BC5 �u�/����dj?���^*�MK卂�< 1����M�n�GM_�^(���w��i;��%I\�S�?�� {��',|P�'�"�oڿ�^���Q����' ����r�E̄*����l��s�?����$D�\�ubǈ�K��3�.�"Hf��p�O�4 1�	�4�&|��.,�Mcw���dr�֝	d^�#<PJ�a�Ik�G�6
q��j���(�Ƶ�A�7���z��i!H��/�lh�B)^����=�I1hP2T�"a�"Pt�AE/� ~�l�I����G:�Ia�h�*TGz�
�'���d���4QX]Г�ԭ$ޠ�y�		�	��H�?��������[�&x行��>������/�0��ad����=���d����'�e�����"��4�dE~D��$���f��K��`�fn��2!���a;,ON`Ð��.o�B�+V�Ӗ^�1����d�tp\�1%�,�'V�'�!�b��#`R�+�m�}ٰIJ�4�� Vm[0	i�}8T te2c�|:�4zh�eX�gU@�l	")�Ѧ��'K�d��b�l��!]8[�T�����:�ɶOi�؀��M�-�`ҵ�NL�6#=� $����	�q6��rt��0RW����8O��c�x!qm��Z	$������&�\
�������&Ƒ;7��k��Ѕ@��@��F����>���.e��@�@/E�*��XYT(J��(�P���˰=)�wcl����׭�����FR0 Pϓ]T����N2� Q0�V) ��봇�1̩�v+L$Q�����{.�H~���&q�̨�r�O2����ߚh(٢umU$�6=S�b�5F�k�(�䉪Ts�0�[��Q�A�ʊ�>l�<�;T7�P��َU
ʼ�VL(l:h�'�V(*��J= ��a ŭ@�Ըs��ѝz�lu+%'�3��C�NØquܫ��F��R��5�K���(O&�PÇ�.%�J8zɄ8TT�y��`�+u���P��'|�u�r�6s��e�Q �M_8�XC�'�ў�>q ��ޔN�NiR�O�5*��*�(T���%9��;LO|R�M�m�Q�E��=z@H�$�T* qHS@��f�̱W�	()ĔH(�!)��T3�˜�yv��I$��%v��i���'�[�Gp�c���#�K���B�!M�!g�p��h(�	�=�U�e��*Kp�x�Äʷp�I�F\�� G�7|̨}��	�M��">9!NזC.̑��'X�h����㓋Sbtl;��9��ԉ��$j�|p�'� 4�"N߆Z�`�;W6)(���R�ob�l�	�Ӽc�_�/2�x��e�flx�/�U�'a���Oe�	qq�\c�D�L;��P�)���pR ÓX4���ɡE2M�����B��Š�%�*��<Qr�Pf>A�C�.,h��@�qӮ���g�	�ϔ7��O���%E6A4je�'z����06ee,*?�ֈCH�<�0�H(�r��H����1�I�����@�x�4�'e���(�	^8k�
����� -%'��F��W#P~Աb��A^A�7'ܙh�|4�W=k���!lOfi�S��e<��;���z:�h�e�6x�aZcfM�e�-I����f���j�\��ߓ.��b��fL�&��$J��Qcs� �#*>@5�_��<����!R�T}"�bԟH��ؚ@�j�
$�B�O�80��H�S��O�e:V��h��T(���*m�<��t�x"ዖ��$��83�T�j�$��zun{(��
%零_c�� �6��)�8��U��*%�$�|c�m���Щ#�\�4�B�� �˓��q��ǐ�{��+�x�#j]^há�>��1��LX؞H3#`^+Դ@`N�%>��r��s�洄�i�Q�T��=$5+u��f6����*�OlY�[5Jʐ��Ƴ/ضl�%O�:=i�9��A�j�'O�aٶI�Ak�����&m+�`���wy�(%ĜSV�IQse�xQ�Pr�OP��B�;a�4u�֑H���O��)@�db�E��;��)cq_�$y��*����F	�;^� $=�M $�c���i[�~��m�ğ�aU(�#r̀`)��_@I��b5ғey889��%��t9���/̎tY����cˎIRf�Iw̓=;\���lN�fe�Ԋ�	ğ 6]۷��MO�iR�'W��Ͻh��!凴:���b��P�,C�D{Zwن���F\������ 'C�ⴣF#�8G���$�$}�88�Z9��;���>[0Č��u�ktZ8v���� &��Ī'OH�#������4
7��� '���n�=VȊ�ʄX���$R�z��#�)]0����_t�"<iV�� /��l�� ر#�����X}�oۜD@��Fm��5)�m���HO��4,̚wt6��2�H0;����oO�C­{CoS�o�a|bI�e�(�&��|������/֐�Z�/�2P����4降b�"��%L���#&�6��)BO��`�
éX?�U�e#�N��� � Mџ��Rɇ� �8�Fg 8� 5�t"Ư9�<\ɣ'2�P�9G�ZY��H�'�
b���
iݡ�w�ؕj2漓6���k��	�鋆g�����^�l���O4=�cn��M����b�̴MU��X��i��5J��Pg[9�b	���L�6!sQ�d�Ē�4a8"�Е�$����S��(O�m��N\�5��MAΕ2?a�l�b�V~�,�OB��i�ex#��:n��S�U[�Y���ي�79|	R��Dt&�ڐ+��(P��$�C7n��K��=���ƋxyT���i�>#�v���gW��z'�*��d�ẳ�O�i��<��GV�S��(3���b�*l��/�-��ON0P��.j��b>9��Ȃ�}���@�?2���>��~}o<?ͧG���u��x)�`�'JJ��q�YWM4,���m�0"�ݘ'$r�H3?�j�i+�x�5A�L�^L�F
`�zuS�&:�$�4Z@ ���'!Р2#�[8�qP��ԓi/��h�O` �$,�G�u���I(t(�y�&��0v���'�/n㨴�$����>)�IK)k�u��H��Š�!a��T9G�=q;>"?�DO�xz�y����E�aPQ^�l��G|�C-]g4���0�=�Ö�H<;�&8r�	C�dB�	_���QDȥ(�����C�,��ɘ�}���B.^��S�O5���c
3Z�|�##�'�%eIc�<A��͹f~D���Sڰ{�g_�I�c�&�b���z8�� d<ea��1�1kK�=�y2G�'�d<c_��i��#�_�����J�p���'W�D��"�5Dl
�oڞy��4�'�����ǜ6�8��nڑvH���'~2p@k0Ѝ�M�i�� c�'Ռ�3��T�Q\�a��
I�5�01J�'u��dmY"P�h�Y3+?1�ls�'F��d���*kjxq�*D��R���'�(��&E3�B�k�b"�%�
�'x*�j�����tH
b�Q�&h��'>�)9qB	ظ����:
�Lj�'*��0.������j�]2���'�tBP��/��m!C뎵����'�6ْN�Rަp�W$�%�F�P�'I�8W�Ą�=q�G��trh��'9�K�&�(3�h!r7����d0	�'w¼����3���/�<
-��'�x���"$�U�� U!%j�'fL���E�&%%�Ӣ�z�.:
�'n<E@p��N��sҤ�ru���	�'\¡0����x�L��Ωm�I�	�'��� ����q�R�kS�<S�'��Q���A�X��)[9h��a�'C4���f
�L��@ဋ,��q�'�ꕳ��L"I�>ŉ"���s�*��'Etu�3DQ�~Shŉ&J�?#��a��'g��a�țL�h0z�ȉ�S����'r�}f�_?EFpk5�2B����'�q��YKg�p�J�=h}�
�'���i4P�H0�q�
)uP�'hT�� 
�r8p!�W��=k2!�'� �E}�� 'C�>e��'#��D�H73=�dy����v�C
�'��p�CLO!h`���ǎ0��HC�'
�@m���� #!h�' ��'nL dm���M+�I~�X��'6�%����w	D���DF!py����'gB�R�l,]�D2b�K�g���'���pb��5#͘ArB.�[��M�'��<�D��<�,��q��O�y��'T�(����;rb|�%ʺ<�H2�'JL� ��a&�jpɒ�3��0��'��-
v�«Ǭ��`�V�*^v��'���P.SFa>eC" x� ��'/��AD*PtΔa��.E�|9
�'R�u��N��D�JpA� ��8
�'C6u���)f��=��NܱNr��a�'y�T1ŭU=o#��`#D"J X9@�'愀I%�._t�#�� HK���'���g���"{�%P�'8���J�'�h9
��D��B ��3�M��'��EK�(ʷ<a.`�0L��$1�'���s��ǀ~��x5���!�dܚ�'�Ԙ�q�&TTH�C�#����'�����+x�*�h�eԗs�*���'e�O�^�<�� 9 ���'�|� ���+�7G�,��'{H����_�8��� D�����'��p+��L�2�V�gc�=,i~(��'"`|��o�+kg���!a�!��'tM��B�l 0�����@
�'N�!h�G]]fY�em�,ZqT+
�'`����Sc���s�\B,� 
�'źqI2�B�� 4�)%AY���� � �PIJ<2<��d�Y�;b"O��(����P�����R]q�"O��a��&L�<)c"���`4@)@"OpRh1��ݲ4[.4��i��"O������q��3�c�60B�"Ov�q�.Vf���%ds�|(�"O�Y��È�6��
F�Z] �s"O2���YhPR�@�VH�-�v"O��c�"ڞ-����%x���c���y�H��n�`�h�*�>�tD{����y�j˥N(eRf��(�00�y�P$}�2� )�;*v�x`"���yR[���i"�=2��`��M�"�yb�+_�ظxF`�>*+�}���yR��#vK8J ����bA��*��y" 6=��jt����e�Z��yҎ�<@LFp7ʐ%u��rp ��y�@�_�@}���Z*tZ����g
�yB�!��uY�� \^>�)��y"���@���]��h��ب�y
^�qф�!���@�1���L�yf!)�UY�o�K��b��P��O�=�O�4�"�/M�s��*ħ[V�Z��	�'��y���A3J����JH�0��'Br���יYb��c��9
4Q�'pzM�0EK�3V]���ξ4I�ĸ�'& �"���{=�����͍`�4���'�Д���Hdif��AdE-X�K	�'v0M� ��9[�*�Q�*ɚ\M�M��'���E�L=Fh�2DDD�@�~9�'C*����V�LҖ]X�Ϝ@��l��'��9�שOxZ���� 1F\)c�'�r`*F&~$R����,�`i��'���;��%J�mu�!Bs�<���+&|�`�6Di+�ǃZ�<���&��D�́;�P7�X�b�!�$ �U&�X��0x�3e��68!�D0#@2������cO�a�!�$ʗVF�)�
`�93���,c�!��1*���Ո��&*�r)\6[!�3�*�um��P�X�seS�u�!��u�� ����P��rԡ���!��N�j,��o��m�:�/ �X�!���|C8I򲬀�R�����)J�k�!��,;4e��d�1{���1t�!��"_��H[�-یpg���J6�!�d����V�G$PK����Ra!�D8Jn���f�0[cu(�K�20W!�K	���x���F]��4��DC!���tSt�F(�XAD�A�l�<@!�^ܹk`��2���|0!�$л��DB��R*m�6b�*�B!�Ċ-WE�3�0��%��!�%vZ}�&�=;Ì�P��N�!�D�"�I��>��$R�B$3�!��c�qY�A:O�N��挞{�!�d�#U�>��У=L�(�#�k��!��R� a�-X�`�5(�(m@��,�!���>��)��j�(��)G�H!!�ϱ>��k �Нz�D-JC��T!�$�9�,�=u�J�+��ˬqH!�dZ�U�y�ED)�~xhR!L�Y�!�vM&�H���=?�&$��� %!�I�'�T�dN�5�n����I�r�!�� �r�lԤw���突"F���{�"OՒ����T� v�4/����Q"Oly�'A'�|��VCK�\� ��"O��)� Ҟ�v�	�[= ���p"OxA�7|w�1Y��Gm�Իg"O \�pN�	�-���:[�q)a"O����B�Jqr���	J�4R�"O\�c�Q����V'��8��T�A"O�����1��=��gA%�Ԁ��"O��
5��:[|X��w �$�"a;G"OVi�a�dHnq�/߿j��`��"O%3�iͧ/�J�
��T�`x�F"O��U���3Xe��	�
զ��"O�X# HY9y��1���f)*(��"O�U��D82[����Ŧw�pu�T"O�A��΅�i��\�S��&+n����"O��;r/��Wc(�)�J��Rirx"r"ORuy�AK�}%x�H��K$GZ<�B�"O�| r*K,2(�ڃF/]�L��"O��%.:�4����lsK1�yHX�?ޤev�<v���5JV���rX���փ�\�\
��9lҌ��u�+,OТ<�H�NZ��豊6���U�<��1k��cW,zq��# �\�<���rN��6�	.v��(�K�[�<��ĕa�L�:t����9G�r�<i@1�X�ӧ��n�����Ax�<����-��a8aΛ'��Z�gsx��ExR�W�n4� �ի �4�����y�cP6"�ґr�$(oS`@X'���M#���sӔ�ywN��G��*q�Fm	���p��#�S�Sp�|�g�G=��I�a�0��B�=H�� !r@ԁ@	��Ç%&RB�7C*�� ��J8� �"��T B�	�X.Z��%��9���ĭ��e���+�5(UP�R�G :�;T�/<��ȓ
��:ƀ�<��zGiT	� �ȓ#"x��T��xF���"1j�� �ȓ]<��$��OE�I����9$n�t�?��4�p<Q7
��ot��K�fW�q��F@f�<a�Dߛ2��5���Z�8��m[rh�Z�<����a�d�n�K��a�'��Y~R�)§R�p��c��wWf����&*�ЄȓZG"�5��{�p�c���=B�)��Gڸ]��hNqV�P2T�0_NQ���fЈ���,%�Zre���n�t��<�ߓ5c2�  $2Sx��f,)|�9�����#tJD�)�8xɑ�ӥ4����q����H�AIŧٟ#@1���F4cWIx�Bdi���4Sb|���k x����pl@-9"&����J�H%�d��i挀2!Z�wxt��T��:�N��E�b¯~�vY��o}�$@�d�d�p�s�ȸ�ȓ3=@��4g�r�9��A28�=���r���fۯUز(	M�V����I���ʤ�]�p��5��d_��rI�ȓg2����H����G�:�P�ȓMΙ� %��o8   �DT&M̔u��c�F�CpGHun͓��:qfh��ȓKg���'gϡ`��D��kD�#A����.��!"��H��H��C��9�ȓG��u�vNU�G)>��&뒄~<�9�ȓYaF�Μ��^�5ʤY���S�? t$����1$�
(c�����p�"O:�H����Q�n�aR��&s��}cG"O����H��\�*�k�%�ޑ��"O�m���'{�� �O�:~�С�"O�0�3���CD.Z�N� ��"O���/�8`��a��:�����"O����L��^��=I��6A�,yW"O�e�u����P:���K����"Oz�Rč�*+� ��i$z�T�"O �5j�h#�4��)Y+h�ٱ1"O�ycm��sʊ�ժ��I�(0D"O.سg����`Y$��K
M�"O6��'&˖j�:�� ��k>L�"O��*�m�+|�J�Qf댘z���G"O`D��d-�����5O&���"O8EIB-L"n��E�S�B�(P6"On�S�����@̐-/'�à"OhbQ�Ő:�p��*�8�@�y�"O���r�G�_ 22sȇ)|r�lY"O���UHK+#]�+䦋�adX�"OjD��#���L�!�J2E�1��"O�� ��n�Ȑ�M;'|sd"O�����;V����҃<!<ȳ"O(y�q-�딜J��� �.)��"O��w�Ğ.`^�[Q�]��ʠ"O����J�w��ɠiď,�:["ObE "��Z^���BY���"Ol��e�+UT����G�RA6�*@"O4,�ыȻC��+ġߴR0@ٰ�"O���1CĂc�*͚瀝�\Y��"O��@ԎZ�$R�� M�|���A"O(�K��'T�(��3n��3�8��r"Oʥ�&�هu���(̓�;����3"O�0�ff� S�M���A�m��f"Ov��_�fZ�33����+&"O���ǩ�9+�����H�kzʸJQ"OL<0gF�C���1G��,p����"OFXj4 Bp8�pv�J�26�Y`�"OriH����P!�b3,Y�n*�A��"O.d�5m�1������2s�F`R7"O��.�H8��Z_Ҁ�X�"O^m	�JўD�~�K�$A?��!��"O.�"ˑ$�\h�㚹/0=ra"O�I�C	�-��bU��w�x���"O����ێ~!���D��%�$�kU"O�4����`�FHX��Q���S�"O�љP��Wj@�p�20�J$�A"O
`Ƌ�+Z�)J`��-��Y�w"O�I�V+H2)P��FLޤSyr(��"O`�X���K(�1��1
�E�F"O�����>�t9���;��=�"O�5��ߟ-��`��� �;�>$�"O�R�C�_�&44A���L���"O�-Jm�3r:�(�oˉH� i��"O�m	運hP�Za��#{�n��R"OlE�b�T?$��m�W�H�c���(#"O�MX��F5M��p��d��k��yCT;P��	���~%B�aM�yR�M#4X�	j� �'L�<�#��!�yB�x(���eB�B�V�8�	���yR툣% �E��ZU�'l��y� �3^x���1�ސkgmT�y2��,2vl�a�؇*�6ԡF����y���NbE�S�Aޖ\+wJ���y
� X �ed��0�M��л{�����"OV�Q���	f�)B��F��{�"O `��M�ht
����ҖѬ�2G"O6� ��C�}uڹ.��o��q{P"OЈ�M�bJ\C"�J����"O���f� 6|d� ��v~J���"O�tJ`͇�T�d�����?�r�@�"O��RT�M+s]�D��͎D��`�"O��Я��#t\�0�����"O`P��Sp�����\�� C"O@��`كW٬�2@���ڥ�G"Ob�hռ���af� �)����"O��cM� M�^�sY�TUQ�aS'�y"Ŗ�]�yxe'�A�1�i�:�yrnդN�ڵ��e��@��à���yb_�N�0��bd��?��������yR� �¼k�$�.`f�+3�U��y"IO�=�*�U쎕A�M�eY(�y"��7"`��h�!�e⠢A��y�'�(Nf\Ia#ˏp��m�����yr�70�[
ʏW��0��1�yr`>V��̪E�M�x`�
����y�-?R�L��Lz��a��y,O�*Hr=ضUv�>��k!�y�$�5��=��� �j�n� ��D1�yr�F4A�����S�Ys��
�y�c�s�|����I�,��H��y��	�j�|)�*�Q�D�`�Q$�y�+û4���y'�ݩQ�1�w�׾�yD� �ա�.���������yR�F�:;�� BT��eD�y��	��q��Y�Dv �������yi�22�����-�3bf��AD)�y2��
T�H��G�t<��z4lE+�y�W�h��(J�S<eV.`"��G,�yR(
-L��A�Q�Ȩc�x����$�y"�^74����4"�c���* ���y�j�9�t��'B�``�(�ǻ�y��� �����@�(�����%�yǦcj��(t*��0<Qo��y2HV�%4<�`4
��� #���y�)�-�XL��9<gε������y�� ;�*�q��-2�ʌ��G��y��^����e�^�-8B�)�	�y���tָ��å$E���CÃ��y���J����1�J=p��I�EL��y�C�0q���;�ŀ�ra��:�l���y2���t�   e덕;H��� ��y��Q�j��AZ
��X���5�y�5Y���P�� +��!@�H��y�0a����gI۠w=,���˯�y"�V���<���8"��0���3�y���Q}H�@��c$�S�B���yB�߼E[h=0+�Z���r��ԗ�yb+��gn�e"b>f�Ʊ��$4�y��A����fR�U�8���ڑ�y�
h	���D�;8��YV#C�y"#�-+Y&��D�~�����:�y���%6�Z]�t�Y�Hpb3�;�y�OW��lآ�N� )�(�bJ��yR��~|x�$<"$
���y!�!dUD�	�fÊ��s��y"�P���s+I�Y���!���/�yiE=4������I�������y
� ]�#��_�&]6�
���$"O4��mW9X��҇H�_��3�"O$�Q�f��t� ���݅��mx�"Om�DKW�<�,�飬�uG���"O�lzSMU�&�txс�&?d��"Oܱ�Â��o�`A5�F�!,*�5"O28 Jڋ|޼�	��t!Zd"OF���(C�e��L%u2)a�"O���a�({���A��eU�q"O�@ɦ�5�u�Ƨ5���"O�X1�EӢ-��ؖ��U���˅"O����G�?�6��B��R�Ą"�"O@��h\��X�1��@D�qu"O@��t��7,�F����J9e���"O.P`c���T���kT�P+e���s"OB��g�� E͠%"�ꁉV܈h"O�A��ҥIn�� S)T�5�2"Ot����ƀC�{�ţ}��Ia�"O8؉���X�H�L�MƤi��"O��`�Rft.Q@�ǕrF ��"OL���C<%`T���]�(P"O�
���?�f��©R�yT�e�b"OVjP9�����N�!R�a@v"O��@�^�XZ���ŕ`��P�1"O|�Ş�Zn���U�n}D��r"O��3ĨBs�d05�_�i��"Oj�q��^64��GoN\r����"O8Y��S��6��5�Fr|����"Of�T	�(x<�� F><x���"O\d�2D�8�$�i4C�<-y:L`W"O��� NU0�B7 ��y'"O�A�� D��X&"ʿv�@��"O�2��>|��6n��@��tp�"OD��Z���O
�d��tB%"O=aV�/Y���B�
Y����D"O�p2 �:?�F]#ScY�k:�u1""OfHpf�8
�,��ȝ *B%{a"O�U�	�=U�%)�g\���;5"O��2e�l�l9CR`��"����"O8�3��HWީ�&��Ƭ��"O�	�'+q̭8R-Z�N�Z Ia"O( Bf*��`¼}SU���>d	�"O�y�L[�h��;�@���]�"Ovc�����̈��֗h�b�"O*j&&�>�E���+H��M¥"O�����K?'����oGG�>���"O���C�	z:��u)~��:"O�Lh�h��l�Z񨌸4�f@��"O�Y`�R�?e0�����Ґl��"O��bGmߢ���D�X4�4���"O^��`��5�8�`��Q��\C�"Od� ��V0�YR�.���S�"O�8M�|�б�ި=�E9 "O�jФQ�@�ܚ���TA��r�"O�ذ �3E�=*0��Y�9�!򄂏 ���3�*���� ��`�yN!�dR�m��<I�#�
���B�E�%B!���������̟.���{$��:1!!���0q�QS��G	<��	C�V-�!�$�H�~}��QH�:�q���]�!�$��~ؘ��L�){*A��!��J�!�A�q :4PV��S� �1��=�!�$E�v)!�0!?��@��]�'�!��Żd6�q0�jB����M&J�!�� ��@E�t��raƸ33L��f"O�9�A+��)�nX�á�(2n�H"O"t�*��:����n���"O�U`'�ֱmOL�&�a��u"O*8EK�9ze��t��I�S"OБR�I�sˢ���)nk�M�"OA�!bG&2���Rh��T��e1�"Orl�,�t�D�3�1p�P���"Oj$1���s̸ԋ�$^�.�P "Oj����0�I�%�M�%�.-��"O��ͯ �+� p����c
i�<�TAY���0��b��k0f`+��a�<ɦe� no���U�ɕy�\u��[�<	�K�J3��X�*�Y����W!򤈵��Qɲ	�<�����A:fI!��?���:V��N�4HR�Fe�!�N����������oٮ)!�$޾T�6q*�I¥C�����+h
!�$��n�zB��(M��1SFA�t�!�R�J���V�4rv��AfQ�3}!�ϙ6|��EΈ�PF�ݓ�q@!򄈇(��Aw� 'C.&}�EE�#5!��ҒF�V� $&\' ^���W0/!�Dʷ_�:Q	1�\�r)�;!�$�
b�r��חq�<�`Th^#i!�D1�\����Hg�`U�CJ��Q!�$N�D�>a1®��b+>!C3���V!�ۮ*��� i��\��À
_!��R�|����#`� a˔Zo!��*<n�Ac�H�n:�I˚S�!�Ȑ40���Lj:\!�J�TT!��dz���(#07�����BQ!��F6�r�n��y� ��G���V;!򤟬D�~�	�h�8"ɠ�*��ڔ !!�A�T_�D�rA�!6�"aSr��F!�d� �p�P�A�2h�<=#�@r�!��\�3F���Fc��U�́å�4Y�!���;�H� ��Τ��� �qR!�_ l�|���d��bl81+�b%!�L�p��$�sH8T� yك�1.!�d8o�AS�'M��X�B�%�!�D́iVt��p皺��5�TG��2Z!�$� F"��!�Z&F�t�c��٬�Py2�i�R}sBKR+�lu[sʁ��y�Î��:;�&�Eq>��B��y�LL6o˒��'G����b*��yRMŽ���V���th��ҳ�yRBՓ_ZN�kr,�)H�~(��҃�yR�T�u�(����*��q��+�y�o8VA����ɡ#��yB(����4#��"� ���yB!�7a��� G�݌F���p 	��yrg4�Ds�Q����ǋ�y�F�	W�H	�m�?j݋҆K��yrN�"�"�(��Ț��qr�!�y���;���� v R 
R��y5B�X��^,cն�ˑ�E��yM��i9��R�\�j���sP��y��ȓ0�Z�) cC�_�,\�WoY��y�ʍ)\.�<�R"[�k�������y���7�R�h�	_�Yz�L����y�F����+���f( y��Ƌ��y��U�W��b�Z<O�5#`m�2�y"�7p���Gc�M�J���,��y
� (]����eIJ�(����"O���Bc�F��XZ��މQ�8�@"O�<�BKX!�l�3'!�9]r�p�"O.y�&C��\�'N��iW�yy�"O�4 ��7V�f�S#K�hTT�0�"O�`م�N�g��Ȩ�M��
��\�A"O6���ݔ�4��	�!-/l)�"O��`L�푓.@':��"Or�K �љm���$(J�"�Q9�"Oً�-��a
p��'�	BzT��"Op)2 �i��Dy���5Zj�Ф"O
8d�޷!��m�V�Q.CLr)�"O�]S�o�g�0�X����y�p"O��u,ZJ�J���ƏS�~LS"Ov@j�)1!��(�c�J�/�6���"O>�2ő��!�6 �;{Hx�E"O&���I^8uw �qeh�zs�:!"O"8��oξo�rd�C�2F�yk5"Of��e���e�5�Az!I"Oic��.0bd��2E�_��؇"O
���$N��)���/x���P"O�i��&�*\��P���*vܱr@"OB%b�L=|7T��V,�HQ�j�"O�HT# :��Uˉ37b!��"O�|�q���*1hM��|�X�"O�<FkX��V���=�	iW"O@�p�?;�9G�Ĳ%\Y0�"O~�����z�H�ǌ@��5�U"O(0����^9
�I��<��"OQ� �I�*�I($F�(+&Mb�"Od<
�-�(�zE�/ `:@P�"OĹ�S�K6nj��a󫖠}L��U"O&s`��
���+�?�,�p`"O��:��"��Հr��3�:�B�"O�!�#��7�((��H<}�	��"O���uL\�#'�H9 g7>I�%xf"O����^;>j���担!0l5H�"O����M�"n���,Ob"�]��"O��ۦ`M��>Q'!
�y�D"O�t�(�5V܈�G)��,h�xr"O ���G�/|�4 ��~�|�S�"O:Ip�@>X�[�	����ˇ"O���e�D�^�*[�B�/>�Z"O� q����N���3��%}:"O��ȕ��aS����ː�E"O��y)�3,E�}�E��
J��P�"Oz������s�����E�h�q"O�,#���9{F�4K��KT"O���	�9{',E���ـ?�`��"O�x�tiN�+t��+a&W,	�`{Q"O��`�X$3F@�4f��R��t3v"O��`��S�Uh��B�)v�R�Z�"O\�3�1Ȑ���.t`mp�"OT|�g��}�~T�Ri�2k`<�3V"OhH���9��J��KeM>�
"OP���ȇ?z����H=y ���"ODtmĪe���z��Ί8�
7K>D�4i l��R�M��L+(��(%';D�T�4���X��=��)Вh_�<�f�3D��y���:e�rQ+u�O5�X�E�,D�\�@H4C�����|^��c�?D�pkf�${���F�'y���UA9D��Q��
g���6͉W�du(b�5D�be�.vJ����R�	�V�цH)D�� �i���z�X@g[���"O^=���*�BX�hj�`6"O��`��H�b����d�'gJ �y�"O��ɢc� ,w�q@�!�>�|	�"O��+�b��J�T;�F'ΰ�t"O��;�
	��9�bK�1>��R"OHX��i;jy�0X�b2{g�1��"O��+�?Dy�����nZ�<8B"O6�h�j 7(lM�щ�gH��u"O�aP��ՙr�|���'&� -;r"O@<���r)��(d��ޠ�Z�"O��S%�Q�);sk� �&iS�"O
D0�J�(IҠ�C%�P���U�u"O�uJؗG�9Ќ�@�@M�9�ȓXe����iҙ2����c8�����X@|hV�\^���0�f^�S�����?V
����JD�:�DE�kg�Їȓ&S�	� gn5+d�O W���)�|Y��D���b�Ðh�$0��X�<�9��5���@�A4"lC�I	e��6#�����b߮B�\B�I(y4t���X��tH$<>B�I�C�������M����>o� B��?��M�A�߾|$��$�̿׬B�	�A� {2�Yڴ�
5�� ��"O� #�E��ՁBJ�e<V$��"O��F�ǉ{��X��Cc1�S�"O�+��mX!H4B
wF�"OμaFKOl�
,��a�69��e"OH��$O_�{�fY�q����l@S"O����"/L�;� ٗ���3"OTA�2��m��	D�0t��"O����Q�@����ж-s���"O`q6j�&Q{z��/Y�+W��Rt"O��VO,:���V�]]�
@��"O,C�ؕ.�x;�-ڛQh���6"O��[&�NK:���I�M7VpQ"O�K�H�#�*�J ���v��"O��ST]�?��Yٓ�Γc9JĈ�"OH�@�⇋,Q�T��F=L/�H�p"O����U��l���G%~�`"O�uCO��Sq�͡��6#$ܰ��"O� �h��ih0����.-,�u"O(!�EQ�DK�%\.I��	r"O���S��q�Ĺ�L�n�.�8t"O�����ȁ:{"���>4z
\K�"Oh1-F�\�F�)W̤SKT��y2�
�+E�1≪Aѐ�`���y���;.<�eOɀ1�4y�![��yb�Ճ[)�E8��M!&]:���(ˮ�y��O��2� K̀@Je�k���y�B�t��ġIB�A9"����yR+߹.ɬY�����D�>(H�*�y�H%9.U@a��C�tX�q�
�y�'��Y�pt����7ؔ(��m=�y�Ɂ�,��P��A�
rp[�0�y#ֲT:��1Q��  ������y�)�)Q$j��~t��z�NU��y�*�p�v f��3q��r`E>�yRd��nxh��2Gs�,�:��O,�y�/E�z�D(H#JؤV����!�S�y"�#X�B8�@2#���Cg?�yR ���L�r�f��<]	�y+�H?p�;�c�>���ۤMɚ�y
� �� (P)��u!$�D8ol$"O�`�Kp;9���P1r�}S�"O�-2d�����S��9Dd�)hA"O��0q�΋�Td���= �4�S"Oht�U�&a���c��)ziܱ�"O ��ᄘ��.�2fJ:z��a�"O� ��'S6+��)s�i��"X�E��"OX��b��[g��cw鈮.�>ɸ�"OI�`�ݥ;�Պe+�0�f0��"O~��iQFuڰzШ>�ޡ�"O�0{����
CdHDG�;�6pZ�"O|�c_;���#1fQ0I�� ��"O���^ A�\�:lĜ~�x�bP"O�� ��� �T�B�K��5��a�"O�{ubV16��b4��$�=�C"O�X{c��r������N�p8���"Ob�����3Ex09C�n��"7"O��Q7OTMp3��\;�Q)�"O�x��(@e]$-3�&~2H�G"O5�#�<V�!�Gݮ7h���"OJ h&b���t��E��06���"ON��¦�c�i�E���dX��"O���cB-!dM6��1ir"OƝJ5Ί�Z��1�i�nHȆ"O�i��I�da`�ʟ�e�̴�2"O81t��M&6A�I
'��e��"O�@۳g�M�����'R����;"Od�7JI�6���,Ɋt.Y1�"O���g�^�Q����&�H%a��{#"O���G	eS�ċ��&t����"O�Y�1��]�dm9��O����Xp"O�8����@���g�g�4MK2"O��1І@��L��e S��0U"O�|Q'� c��q0$Q��8]��"O��c� ��)A�c�>�=��"O��(��ގ=�
�:�'V�o���`"O�x$o����85d�:��<`�"O���%bM���8 ��u��2�"O���T�D�v�@Q$�3x.	S"O��i�#�nX�I�vm��8]�C�"O �0a-�>&�$��`9j��@"O�
��k���È#-Pp�`"OrY����^;B��AOȆM�Z�u"O��@u�Q
<�d���1�~8��"OΡ*��%��$ر)�5o����'"OLhx��/N4�d3k��T��H�"O��ٗ̋ ���p!j�(c�	y�"O�ÆD��,X�UV!cb\��"Oh�bR�ߑL�r=9�`B� ���Z�"O,�R��Oq���2�IO�و�$"O.T�ՠ^|/���S�P��@F"O�EZ�OetnM �Fګn�D��"O=�&A=p߬��w��7E����"O�$Ae�2i�N�i�N�,��`�"O�1�2J�=�~�U��+�p�a"O� ��P��B�%�2R�P"Ob�a��P�V�F�Vk݅
䀈�5"OV�්�"?It�����=^�t�Ht"O��"fK1�}�#�N.5�L���"OJ�"aSr�~p�DJS8FQ,��"O��I��] J��1��j���e"O �왬O�@�) ��1+����"O�Ӵk��gW��Q��B�8�"O2TS@k�;(�BG闲n� ��4"O� �4nٙ9���F	"#@d�@"O���P	�1�u��!l$ِ"Of�I�����'E6tz��1�"O m
���"<DT�ku�D�/cHxa"O���5���l��Y�UPa� "O��h��I�p���1�C�rC��3�"O��QjW9a�,ehŌ]�?�b1"OVDyVA�W��xg���o2��6"O.h����I�􉂬VL0��"O|��f51�R�r�ڪ���"O�<�&��0z:�!�ǩ-N1`&"OV�Ǫ�%UD���$��b��` "O
�s�&���H�� &�8i�Z� �"O��2��-,�8q�%+W1���3"O��CS��aaF���JM'|��L"O���c$��U�ńW����S"O� ��I�=�}� \���7h�0%�ȓ'��� ��7�PYy�+��obm��B��-;w���QiR�ЭpFX�ȓnT= `��Q�]��喕F}�ȓL��(i�AL<T�X�ʑ'�@��(Ąqɑ�8��E[���8m�X�ȓ"$
�0rk/}R��ۈ0���R�"�pՂW�/TAsA`/Cp�ȓKXTaq,ԧC��X�DI�Y`���ȓ{ء���H����F��'t�h��m�ܑ	"ϗ�'�D�B���K4D���oV�j�b�JC�	3)(����.D��Y�H�0lNU��!ѲzZ ���+D�x)��,z(z�*gA�Tei��)D� �(�y�Q���6$ɨQC#D�
�͑0"6��/I�w�̓f�?D�HC�^8�RddFE�2UH�#D�4 SDW�X��Ŵ"4����,D�( GL'>�E��$
�.D���ᯌ>CM�<ɢ�D�}}�ł&�*D��(��R��f%+7n���(D�䚄@�%E�hJ`�+MC�]��(D��+�$6p��P6kЂ)(�&D���c,$)��$v����k
�{*!�D"�:�ZӠJ?qr�ͺ�IѝJ!�[�7z����m�=O4Ґ���D�l�!�ě�X�V����0|&��!�ꄆ8!��K"?�����d�<hZ�Q*�"!�M�<lJ�Q�B  H2�	qC��I!�Q�(��X9��Z�f�~��b��y�!��	7p�xPS�rͲp �o E�!�͝0>b	�Fk���H���I��!�$ƏW����וzx
�����%j!�@����6�Y���8����9�!�dZ<�C@��a�������!�D�	_�2�%�IS��@�$�ʷut!�9eo|�Y/B1'����䈧%!��	:s.��!�Λi��ITdG&=!!��';
nP�D�������� !�	4��b�!� 4v�Q+�ƞ�Z!�P��X0"!ŎXb�ڒ�z!���3y�<�0��N�l�,�b!�d���0Y���Y�i��e�ɕr�!�N<�&�
�"P�8���)_�C�!�I	����E�h��b�(|�!��L�+����oP:ʘ��6�ˡ�!�׈'Fdx0S�[(e
�-!'g���!�d�Pͼ$�A�V��,!9w�T�R�!�� D	�S�\��`�� 6TJ���"O��"�	�`��M:�M�G!q�b"Otٻ'b�.�ļ���G�`�HR"O�e�ŋ��|��Y�t�.W���3�"O`8�Bە Ɲ`�+�%��H�"O.�ӡ�G>I����*K9)UN�11"OB)���oR�SP��P<L)�"O���$�k9�gCԋ7H�#7"O� �P�J+	���`6 J4�ʰ"O���ŭ��ޙ;VΓ##/�D�U"O*�����"t�b�OM|i*@"Oj�@�D
>9d(������o/X�j�"O��;���\�j�C�Ҝ;=��s`"O<��4"�:>�Œ����-����"O~����L�U��8�P됂�����"O���C"S�*���
��"�"O��2�'���=����C��^P��j��x�Nƾ*��+��D ��ȓ3:­�  �=���� H:���+�U4E\�n6R�B��'ոp��.+�
T��'*\BdPR<�0��<vл`I~ϋV���U�!�d�1��Lb&��_lP$tJ��TS!�d�
��d�NO[H)��@�SL!���,/D�w&�r>��� g��^4!�� z��42Ek��rC��	0#K�()!�d�H��% G���L+�!]�m{!� o��̢Sf��95!��q!�D�K���T!��8'��j����q�!��O���yp1d@4�x`Ae�]�@�!�$F�[/.)��Q:F	�� ��/Q�!��B*%gĜ��oʕ>�����G�>�!򤈘x�\%B0(�Kp��fd�U�!�Y�=�XpZV�G(d�l��s�ѹ�!�ۇ{�� �U��2��"ԯL!�$_��uj�*D�>W�D@�'O�x�!�DŤ�|q)�ϔ�P�6FϜ5�!��/FG���%i��)���Ӏ��b�!��4i1���@,D�Jt~8ˁ+ .�!��	#l,8(A��Ȑ�N���IK,C�!��8Du�W�ϟ����$<#!�$��e�n�0�M�R"��/�	���b;��!��#RP�rt(��y�/���k��WZ1�4�]��yr��+ tH��̝�Ns�xѰĊ�yBKbq�ᱰ[�S�
C��W��y��E�J۷�K~2E#��}{<B�	
TV�Qu��3H�t(��n��B�	�<��c'Ş,[���3��CR�B�	�I�:��e��������5B�IIɦ��`-��:��Q����>:
"C�ɎVRN� �L2nЅ2Q�V�.C�%B��͋t��v��e,��f:�B�ɟ<�&�R&��T.Y�%b�X�hC�1p�z`�U�̳Xoh􉙗=TC��/�l� D��YLzP�q��vC�I�u�l���#���1�(!�LC�Ɂ&0�xh�B�3�	2���=�jC�	LD0�0��k)4�iGc�V�TC�I�jԂ�,/yM��AMɧ �C�ə{&���]y������B�B��;�,�B��
65�D���L(�B��~t� 4KW'8R̀:'�R�:��B�t�\�z`���}����/�k�B�)� P�kU�ǅ.�x��b���8��o�.ukƀ�d2@hH�DM,C�2���\��@�����n7́��(o9\l�ȓd4 ���Y"  )�T�J^0��=yib�@�f%��hԗe�\q��;��"�-S�;��RQc-p���ȓ�T��a�&���w'��Qʴ4���@�j3���g`�<��@!l�|Ʌȓ|�~�Q ҈�,�����V��	��)|*�ե��jH���+��>�$�ȓ8�Ԕ@��T�^a�@o�ְ�ȓ1:d�臢n�L4"ǩU&�pm��7 f���Zei��y���9��!��Xd
�" ��8A<�Y� �M�Ԅȓm�b��͋��(k#ǌ�^4�ȓa�d飶� <S�P�Ҡ	`f���ȓ5�������O�X��ƅS<^�U��1Β͚RňZ��܂�)��E�ȓ@V|b��ū?v�5k�g�1Q�L���_H��wjK*6���]z��ćȓ��)����wQ�ʷc��rNF݇ȓ}������h��j��O�}�H��7D����G�
|��c�(t��l�ȓ)s��F�΁Hw"�B�K�.9�T���$?T��%�����쉬v�@t�ȓ^���M���p����>u�ȓM�¹
�bM{*h�@4��C�B��'Ϙ�����$u�@���ȯW��B�I�����K=r ��nD���B䉠XB�=3!��3Br8�Ҥ���B�	)I�`�z�"ȣn���*��X+8erB�	�0W�y#uo˕`|���p��\�dB�	>h0k�K_?rz���g��;�XB�.H��M��&'�:��.�#IB�	�����h�<�,�el۹u��C�I*_�plq�aM=^3��w�hP�C�IqV��'�����C@xNC�I�T��K�ڐI����n.C�I5oڲŉ��t!�V>*m"a{�D0T�LRS��;c9�Đ�(Y,3x��K�"O����_���?�(C��S2�y�gV;WK���`��xX�e�S����yRk�"}������$(�s3�ֶ�yr)G	U�Z��ʤ�Iq�/�y�@�k��)�$�F�s��!3���y��ϯ'��D��i�����Β�y͗7(Y� #a�S�Y A��$٦�y �>�V`�ǐ3i�~5�2�y"���ul�8Z��6BM��y�ɛjX��xUn���y�Š^��y�?��S���6������ybLԉ-�2�Z�F D����!�y",[�p�f|���GrW���˧�y��T�y�(��a&��Г�ɝ�ybO+b��	�!��A��,��yR��;���k^�0�ڥ�y"₤T�A�蓠r~�)�ϭ�y�Ǝ�@�<Ĉw��f���(���y���V�*�
�΢^1x�J��ĝ�y2�E�f��1�������ʕ%���y.J:eC���S��	�:|� ���yrJ�vst�j"��
��Hcp��+�y��,=ʶ���Ù3?�{23�yraB.�t���G�y#�x�!J��y
� ��yq���g�湘/۰qG�E�"OT��f#�Od���l_�@0X��"O|MKV��.P>i�2F�4�es�"O.��1D�!;݈r*+��`"O�̹�B+cJxT��F�itf��"O��6l�^�u�Z3xa��a�"Ojq�S��]���&�WSf�(""Oh�V��iZz�X��A�CN��"O�<�uAΔMKx�*D�w�H���"Odū����c���+U��x�۔"O^Yɔ/��:�2 cLL�� �"O,ـq��'6M�uH6ĕFo�E8�"O�d"�Cζ]���b�/�(��"O��ѥػkS��!���f
""O^X`B��?Z#��i�K��`�"Oč0��/�N� 0�ʝpy1��"O�� �O�2�yc�J"O���BF/'�����
 F�13e"O���%��s��E�&��:D���"O�	@̕�~܀� �)���"O2YBQË�-]�d�v��MA��"O��lM,x,l��b����w"Ob9Ұ`��	�j��`����%�P��y⧊
yh�I1𯇓id�+plY��yB@�`&�5�-Z�ʂy���A��yra .h�.$ys(E�@1f(��ʩ�y�J��P�t�<h�t�{�L��y��9�`���B�Y��h�@ʐO�<��b�~lt@�ؿ90�
_�<�%!yw���3��?J]%JDm�Z�<Y��E3q�Yx�O��E���1bh^�<��܁JΜ�C`,t)�AWD�<)f&T1*�d$�S#R'O=x�sʙ{�<9��4��`��N�*��E�g�O�<� �ܛ/��($�)t9���h�`�<�R#W+G)��u�G%NfZ�p�@�E�<�#��"Rf � �ȟ_:(�AF�<���0C��-��E��d�)��E�<�QA+I ���K�*��d/�}�<Q�O�U��B�$,����Nx�<	�EFS�� MxR
`X(�N�<Y� $鶅Z��'F�	6��F�<�b���G^���Umы`��x��_l�<	�^�fT ��IC�D�����@k�<��b_�SnL@gl��O�����
k�<�G�h�fAC�O>@��)�F��e�<�2�Z= �H�r��O7<FTt��CGd�<���'[ \��@J���زL�]�<�0��Gmt	 �O�mD��n�_�<y3&�%z���sj��Ub�R��Ad�<7E�@�0���[pڸ,j ��b�<E�>4�A�S�ܘCm��C�+�W�<�f)��^$0PEO�!� Ř��T�<�C�>��P�5qL�@���R�<i �\�@d���ԈH�=�9��YM�<IC�ThS$��P�Dّ�JI�<!�W���݋v��|�<с��\�<�D��,��{skG3+|!��Q\�<���R�Fah��H�U��8�OV�<)�e�TO����.�]W�^O�<�&�."�@�Z�(�+`�0��%�@�<���6���c���rr�:f�@�<��/��J���3I-@�>��C�&T�0��D�vb =�p�*Fe� �"D�� 0���f^� �K�葏_���"O�e ��X1LA��g�6K�L� �"Oh$��Q2*�H���f���JlK�"O��Rd�Ľy�,� ���W�$��"O 쩰 ,RҼ��.�	@�$�jd"O�bP"�.�r�k��6{N��"O��G�J��PY"��M":_�hA"O�c�ŧ0dQcd��^(�j1"O��a�֖]r��V�@_f�a�"O�EH�J��I�ru(��0mcȐ�c"Oh%C4��?0jt�Д��K9x�X�"OR@siz\!���ą$��"V"O�1t˭ʴ`���!D*��R"O���KC�[�uJ����5A��"O��x��ڱ5���SN��=P	�'���Å�F�|rJ@a�·�uIxh��'��1�ɓ�M�Pm 6�Vk�)��'l�X`�$e�F a��H�'��1a�%�>	�d�bG�#_lP9�'����R�ʈ8�@ ��'�
SjU�
�'}�Qm<J�h��s���w=ā��'��<Iv��n����D �м��'m^9�����*ǔ=(э�I�F��')��?W��M��#��;]��+�'4μP�mJm(�a ��;0��:�'\�IF)G�0<���ˉ-�p���'\6e�p��1�*�%��7"W�I�
�'GX}2��/�@�I�9k�b�C	�'i�Cé�~_Tɢ�ȗ�W185J�'��,�#��g��4�G>T1z��'K�Ɂ3I�A�*�[�m߽?�6��'���ҡ�̌\�� ��͋�_ző�'�B�c[�_�2pZ%�R��`[�'��0��̐X��Z���K�� 9�'�b�ixZ� ��`�3E�V���'�9��@���}��K����'�p��ꅗ90�[D�ƌ �p%P�'�VA&�KI܁0�L=y�]�
�'�l4���-a88��"���Ш1
�'{��4�\8{�$���Y�Q��'_|5z"l �Qn<���eK8vH�'`��ѧ-O$���C3��-�'ZY�"��,s���1cm�v��9�'ȘH�j=�8���o����'SB�h�^4hBA1�N� Inx�'_ީh4�!d:�6�������'R,�BG�#xLzi�l	#����'":pR5d�(��HC��{����'�R��gƾ��@��߼tɡ�'�Dљӎ�6 L|�Q�_Ɉ�A�'�4�A�E��M��q��;QT\�B�'	�
Ak	- ����3I�:!�'���w���V�>�"C�L(E�"�'��)5��R�ru[�J Si�0�'4�%HsY3^0
��@�J��t��'�N)�@�/`��'���B.Pp�<�D�$��Ir��L�.��lb�J�C�<��a�Q*T�A�`@�x����'F~�<YQl"V���7��-J� |K��Kv�<醉CiR��C",��3y勄��\�<�g�( X �K��D��ہNn�<Q��+~BV�S��VBl�'�t�<9�(8f���V'���:RG�Ys�<�m�2ք��(��g+���c@z�<� �h���+U~��'P.M[^��2*Oܨ���F*�4d�Ǡy���'$����}^5(sfôn�NP
�'��(����v��zSJ`�����'Ŏ��`��E���(2��H��A�'�`T�t+.>��	�۲,;����'L���_���b���'�h#�'|�*�g�.ȑ�g��&12�'Bf��U��-&Yqgԍ]�
хȓ��[�k��i�� j��8��G*q0�fʞk��+���>\�����rZ�c��T��г1��%]NȅȓJ:t���)"�����/�䔅ȓ|;�Ku�G�tx#�*�"cH�A��bV�a��2�8\;��!~Vl@��uIRi�"�<#�<8S�g�}l�8��JS���"���Y;�j�؀t��3ۀ��!,��DטȪ �H/r��u�ȓ"���aG׆pX<�p�1]�)��h�$��gG�E�i+� ��`d}�ȓt��D�Kd�(C��,s���ȓ[�Tp#WAX�[�2�r�,�Y�����t� ���7yȠs�X}���&���
6$�c}�	���ȓ� ]��lN�g��h°hL��<�ȓGH=��ӱ#���	@k����ȓ"=B=�g�ʬBH��S�/�4���YWJX�4��r90e	P�
�ȓ�uz�D�J@0���+G5X��ȓ,첐�0찕��)@&;׆��ȓ�ش'L�UQ��ʒ-N=a3�9�ȓL�!�0�(Sj�mB�n�!2:D�����6��39k��*�U�%�j���0d��k�K� cZ ����jJ>͇ȓ��x�s-�t =g&ɠep&h�ȓM��@�D�-dY �)���:�½��e��A��ćI� X�+ �	[Vi�ȓ�`����:B%����݁'�:\�ȓ|��=#i���HQ�O;g(�ȓi��G膋t*���.�7X	��:90�sS�Xd.!�D@7L����d!�T���  �� �J�0H�6E��($�|�E�\�w�T(x�`.amT��ȓ V:�3!螏V�>Eԅ�,v�"8��Cn��c�ͺ$jT��%�1h*��:1��d�/K�z�sҬA�ݐE��iعr�`�P�n0�Q�J�=��ȓRhZ6 D�@}��(`�
e��{j�h`��*��=R�`&/�(t��O~l�J 'i�\m@�� ~L]�ȓV�����怣k��  �o�v]20�ȓL��3e�{Z((��@PPu�ȓX�="���,:^Sr�܊"fTl��@���w�֬A�@��pG
h@��ȓZ*���e�7�$�B�)G���W������;b��u!�!'^|�ȓm�|Uj5���#Hh���6a*Q��0�έ�6O�2��}�ꁌ_h��ȓR0~��ȕ�y!|	�I�
^�l�ȓq��'�x�b�<����ȓmv�X�4��8Y���@�OX�f�lI�ȓ
�NU%�Ĵ$}��V��?s"̈́�S�� 4�/=k��9P�2]��2���@լA4��������(����S�? ���Z��堠'ӡK^� "OD�{���z���9#%��.����"O�(2WN�?8�-I&��h���H�"O b4��"��E��c.
�v�0C"O�� .��I!l\�Sϒ$�b"O��1A
��Oy>���e�z�h�ɓ"OT4�u�U�d�c�+K�~�JE�$"O�d:���
3?l�j�� �D��P"O��A�3c>�I��7�α*�*O�(6��M�:�ʅ)S�8B�؈�'u��k����804KN�2�rUA
�'@�lx�Ɣ0G�r�FH����"
�'Z ��͒�'��ljvCMdii�'8�����A?n�{aS�X��i�'o��qVX��h �QL�4Q;	�'�VH´���l�hT3w�W�����'nȋCJ�_y^P�F"���*
�'p�æ8�����R4 �Fd��'�bx��(C��r�X� ��h��'��!j��F�#Gf<��	Ԗ���'�  @D�C=(�Z��	?n~ ��'`��E!}��Y��ʏ_�V�	
�'�6�[�
%���p�`��|r	�'�X%��70�`��U�_5T�4��'�pq�'Ŀe��ݳ.��P�*I��'dh�Xr`�%<�VdD�B�
�'q�����cu��[�O@lAq	�'EB��s�_/Qʤ0 �ȉ�
��r	�'���"�lZaQ�t�4%Y �"���'E�U:Eݪ�cDe�%LPXȋ�$.O�q3�ζH�X+׆��f�P!"Or�
AH���y�!��1�6ԓ�"O���F�B��}�k�PI�!�|�)�()��F�ˉf.�]P%C9�C�v���ٶm������ϟ NxB�	*p�������-4��p�ɱ.H�C�I�"��eJ��o��QAÈ�ƂC�3{�&p���9Pֈ��˘quzC�	�s-,�"�E $GX!�aD��`C�mL�1f*��;���焰n&C�ɦN'��;5 ��g���cuE:>�2C�	�KOz�1o &���#���<
(C�"	�@[�� ���ܘq,�eؾC�	�C������EC��8T%üoZfB�I:d̅I��'[�d��4`��\4DB�	�<3�!��b�k�(H�D�� g����0?�v�D�:)��r�d�2�˖A�~�<��(Γ@b��$M׺y��0�'~�<�F��!'�� µ"�adR�B��y�<�"�I'o�萋0�B�d�4ie�@q�<YS�Ќ|S~�aAꌗ%��4���Bk�<�`��=���0�҇>�z�3�Ue�<'�X�L�p$��`�� ;Jt�7Cd���=�C�_<?l�D?f�	,_'�B�	��J+e�	���F >� �'D��%��n������S��1:7h'�IY��L�% *M5ReIwƛ�����2D���B�:]�V�A0,؜A�,��b/D��`�ӭ�
�I�l-	��|ط�+D�h���>L��aa�^< ���tJ!��O��GG.VS��3A��Q��hO�'vΪ}�5\#eLƤ�P��5C�,�ȓ�B�SpW�*�P�RQ��r�X���I]�'AHpԈ]F$=��2V���� ��b%���s�9YH�8+z���"O���M�]�бi�u�y�d"OX0�QC-�V�@!���<\���P"O�D�DH2Km� x��ѱCHh1d"O�	�す;70Z�E�\`���"Oj����J� p�w��rc�	D8�P(�`@�Oa 9Y���+~���*D�<��H|=2�J�O�~Ϯq:ԉ*D�`��f4� 9�k�0+�r���-D��TƓ`kBH���ٱaDl���7D�,qg֬�@}'$�I��u��� D��S�N@�Wx�HQ��y�ac�� D��"ī 5�`��b
ӟk��I�/>D�̸q
Ĕokl��Q��W���Q� *D�T�󢆍n6��zw$[uKJqa�ciӜO�S�3��޿l<Ru���!�`���BJ�Z9!�ĝ�)�^h�f��) �|C5"ک<>�܆牪H�����5�p�b�?<`\�b����O�D��O�l+d@ڀ��5]��F"OR@��k�+�ؙA����DQ����"Ore���'B�nH��=�j8"O 1��<*�*\;S��YXn��%"O�����ҋX)z<{��\�SP�	e"O��B\�4�P��aؖ�h"O�!�JW�<�t�pGA�&���Z�"O�qBe�½J�Pqg�#h�d!�"O>| �@
?8�V5q���*^� �s"O��FC�9&�y�the}q�HI�<q@E�
�L���`P	v��g��E?��(j�!�b]:}�V<�͎�tT�ȓ@4��H}��x0I�% ,~�ȓ+@si��12<7g�)�I��	I�d�Zlf�0F+M<\'p�@�2h!��
I���A���X����N3az2����'k�	�ъ
.O|EȰ���!�� x
�=��E�:ꈍ�¡@h'!�d�t�$�q�&B��� �AQ !��G�`�jUi�7u�Nq��aVz1!�dW�>�����舫)��- !�KG!�M;]��$��?2txj	�_1!�D��W��5�p�0_qFU��*�!�ԣ+=Խ[t�͉Mp��������{��H;���B�߻Q�tbr�L&(�qO����-I�R$b0E�~�RU� X�L�!�&1C��[WEߡg��)���S.�!���b���-`�ӆ�?~!�Q�	�M�c�ƽ!�Li�D�3p!�֦PD��J@*99Z1@VfЭEY�ɝn�|×�&�"}��h�5O ���ӿ�0?A-O�P���A$�� I�`D�w����"O<���\&/6�P��͡�@��R�'�����&[8.ܸ!a�¼E�h=zF,2D�\���9%iᐋ��b�t���:D���A����b�_3] �c��:D��� ׄ���ʝ�9���8LO*�>��BX�R��Q����D������m�<Y�,P�\�<c���!�z� ��X�<�O�O?�ؗ��,���'�J��Dd� ,6D��r�e@�F�$1�fć��:*��<Y��'7�4�1��o����.���\�����	zy�lԣnΊ�4�LS&�a��V��y��ާn1�!y��ӿ<��L{����y���1B��f�2�)B�!Э�y�Se�� �{;
�X�"\��HO�=�π ��1���.&� 4K�<��@�"O�Q� ĂP�������Nh5�K�<��`�� �Z���V�jя�b�<i�ŝ=P�����!���0=�Q@�g�<a�#�.~W��G�,@f4�CLk�<)foU����K6#�fP�ɖ��<�&c7�.��0��dE
��+�V���0=Q��Ƭ#�z���œ���E��E�l�<�4#F#x�,,i���Y�H�j�jSe�<Ico
qВ���&�0>��ӂ�]�<�4�,T�	B��{>�0c�T�<�
+&4 i��Y2^�Q�3�T�<��M�)x���t��Z�J�-�6C�ɨz:���C6Y}��yG�C�	�"8$ۄ%� )mڄ�ㆇ�/��C�ɝ����͆
�8�Q!�8#n�C�ɷc-�t��M�hx�@{1 �(��C�	)Q�X=谊̌V�nD�TD�h��C�?�p`���P�I!��,|�B�O~���� J�
�h��A��C�1s|(P%�KE�`x�DIX�c�C�ɭ\,��b�3tH���\]�B�'g��L҄ �{.!ЩL�>QvB�	i�r��eլw,cօ�uFB��X?�\3��l�<H�"�I�$B�	4;N�IVI�8���
$*ȩ&��B��*ff�xÃ�y��p� ǂpˆB䉐~v���b�0�CB��Q��B�	�g��tb�4�J<�U�V?f�rC��=e>r2�N �Z��fG�
4�@C�d��-�v��z]x��@`��Z�C�ɀg:d�IфP^����RG�?bDB�	
.�L��1�(��p ���$v�C�5&Q���V�jt��c�0�C�I�)�|��g�jC^x�%�e
�X��,�`��֬�8HF����}n�p��O�x=cbŘ�l&�y"u�P�t�>5��3�-��(��"j�ˇ� �T��ȓ\�y 3����7�V�\^�E�ȓ.�8���?-v2�jJ�3u�4��f�F�YW�F,Gƒ�yUf#R�E��GyplKg�M��Qb�����ȓUiPh
�)s�� 'F�~��ȓ��5��"�0Xxm�����tu��b5 A���/^�my�e]�v~rЅ�EC�y�m֌N�p�%%Ѩ-K��ȓy�����/E89��Tࡀ�/u��ȓ}l�u� O�1:Fr��1Ɏ)a5����9mH!	 �{ˌ�HDO�R�J���E�e ��S���Ɨ�7o�X��Fޝ@�l0f/$E�a鐙V% ��ȓ
.�ɻ���*y��-�O@�+la�ȓ�04V�L?v�r�Y�`�:L2��ȓsN���)J�H�a��A ���ȓl�,U� �]m~<	"b �#GH��ȓxOnH���/8�����1!q `��m*4��s�̶y�j ��ۮ�|�ȓf�B��гZ��*C���X���ȓ^H0�Rs���k=�0�th�*hT���ȓ<��pQ�dG4~�81mՍT8R���!|���ˑ�#Qΐ8��Q�"��Շ�E �8gĆo^ҹ��!�"p�T�tIr��\���G�� J�D|Й�dqg�۟�:m��n���y���,,�E�2e�O�Z`L��y
� �pr��@�ZT1����${���"Oq(&��fDd"�^"l�@��"OD}Xa�V�I�����a_�B[�"O"p��Q,w��j@-U�@���'�)ࡂt�H�/�U���'��ݸfLK��-aw�.N�UI�'�D�i�B��4�4��A��;���Y�'���W�&F8 @�(���@�'}�8��۷@����P8���x�'y4j �)J�l�RHߨ̾գ�'�l� �?]���;�Ŷ��x�'m$e���O�x�6yp�����i
�'�# �Cr\Z�˧	 y{P���'�� )$�
>x
�����|\���'����D,V�r�rFk�/l�\Ƞ�'���Ci�h!SD��3=�T;�'}��٢�L瞔R�E�7Ԁ���'|��E�@��h�9�(ƚ!PP�@�'���*��T���MQ�X�����'z�h3�S�b꾸)G��P	�'[�LH�Z?]�Lx�!��P�d`�'Zް�Fa�z��q0sgT�����':d�&�D��b��"�[rP8�'^�Ё%2B4��FPQԐp��',r��qG�H��I!陊~�v,��'�
Lr��C�|�`����j=��
�'k�\�3��)u0��IP<]O�R�'���K-t� %b 5V#�@��'<j%�Vf��P\���܃B>��2�'}�Qc&���D�ڥ�Ɔ9����'db���,'o���D�S6�0�2�'�6b ��!������̳(����'-B�fc�.o����3�ȹ)�(�'�>�Iw�2nhe����d��'{:!��&\�0���҂
[(
�'K@��1���w�d�+刋H�<�u����8)�4Nǅ&:Q+0el�<IJ�͊����b��J��s�<�pHQ7w-Hڱ�E�VQ�
��n�<A�d[�<�ǀK�1Jp�	��n�<yDk���t���OE0;ޘQ��G�<QD�F&`z�$qwd�.`炜���T|�<i�FԸШHH�NڞMX��ⷬ�~�<1�.�'���Ѝ_xh�*1�c�<Q�HD�y���2�J�q�\`�&��V�<���-~���.@�*��D�V�<!�N:��}*�EגUMH��WJ�L�<�RB�0�X��$� ���B��E�<qvCӁT2��d@\���	Z1NOE�<9b�!o������� e�Xik��F�<ɗ�U�4Q���f�>�JтB��A�<��jSҢ�4DB�sM̰��}�<Y���8h����PH8,�rFf�z�<��kZ8��dX�L�_ (�"�K�<ye�"n��0���6���h�n�B=���ݚi64P�$BD~�:� �u�!�s��p��Ɓ�L=�F�\2���W),�\��-H2�r"�dЀ`�`� �!O���ݒ��';)
 i�>$D!��Ê g�
�2�'�8���9GJ�LyS�±P�<�XO���BF�`�qO��1�&�3;O<D� �ޚ� (J "O���Ƨ�V��,g䁿ba����D�05KXe)ÓbH-�cl�+A�vԠ��]�XB�0����@�3��T�sE�z�!R��H*B�)� <��mΝ!i��ZVF�l�ځ���'v��1C�Y̓C�����C��I��6�4(J���,�6X��/,$q��n��ep���O>���*�Sܧn3Z����#Z��B�I�i�< �ȓ#��D�/q�l�7��++z8��y�xH�LS�xؠ��펩zg
���U�l��t��5<2�@Oӈ)��������BjB�,/j�YwoM�a͜X���Z(ЃG�?ll�c�iةYT���~L�@K��Z�;#j�;Ո>Е�ȓ*�� CbC� H�S�İR���ȓJ�H���6�D��$Ҥ�t��9�zq�Q�^Br��`Ɯ	��q�ȓ,�L	�>���!�Ʌ>����Bm^��nX�A�H�+ҏ-�Xх�l�T��b���5(��ܔ�� ^l�#��B΀���P�y����@EI7!��	a��2��7?�؄��]	%����<��V6&nz(��fh쌑3�ۈs���P�/w�(̆�@6� !�ȞP���'�Q �
$�ȓ=�H�I��,Yrk  ������p�#$�	?$d1�7e���u�����U��T.
q�1��W�Vt�ȓ2��Փ���{�Z������u�l�ȓc"��"�(O�9��J;mV�<�"��6�:�xbᑄ��p�WW�'�H�x���&M�I~�4�P�Q�v�8ЅޭLW���f�L�<�@(��v`0���Ш#��@$��<y7f�0h� ����@��)�'�ƽ�4`�U�)hQ�ix��*�vM�V�W��9Q�cL�Zc��2*���M;ĊU?$r��0������	�GAXDCl��(*r4b�(�
d���$�8��Ȋ�>��B�z%���,�M����U2=����@GiX���'�G0
?F)��ۥC|����;�`������6T����@z������x�~|�&�Q�[e@Pҵ'�>�F�VKj�M�E�'k̘PpHƦC��@.�f��B����tD�D��t51�!٫'mĈp0(�G�� NV���w���QJ߫Uk&��I�d-���	�'��Y0�
0_Ś)�v�g�6��q�G� ��,�l\X�)n���N(�r5#�o��������$-R�}�ذ&L(��Őu�'|O��:��܎\,b�p�͓�;ΐ���J)�L����#\x��S��*n��j�*��H��-�E`W
<Æ���؇z�*P����U.@C��Q�xu�O�)ze�ϲ	�Hi�b双@�2h�F�!P��$���7#rDj�ѲT[�H�#.W�i��3��r=S�=�pq���8@�
�z� �;Q<���j٢&ǂ�3�A,��k5�L":���	�E��*q`�T7�4�s���$Î�#�ɀ<�h�B���i���7l즕��'u*��2l���C��J�6*v��G��,� (��Kιum�,x���)ds&��lA����+'F�1%h�z��*�:���
��G�f��ƭ�3>��|:ߓn؆$��I$d�$��%�[�^��X�J����ᐓ��Y�ͫ��M��Dً�ۍ=bV@��.�>Y��\�Jų��ی?fPL�'��(a쇘S��Ҡ��.5�z�����Ў4���S�"�6�h�ST��$[g��/�>(�uC�(� �]�IIL�!3T�.H�r@M2E����$����$c��"ړ�5���,G�\�˗mC5z����� ���k�9{��,H����x``�@�B�o���~�H��-@�ᝄ�Rp�!Iǔs�%���;�U`�Ň��>i�̈́�pj����Ț�X���C�0�Z(i&�;h���e�iVf��aF�
%��H[g�5^�"t�����;��ɞ
2!JB'�"Jr�9��ϲ��=���pE�san�6�͢ �~�ikd�G�w�`��	v0���Et�JWA�'	<�����Ɛx�]�!-q�\�����j�Q��B��m�<��wH�����(>����@���{րER��N�8�&��C+�v"dBR+�+y�Bmh#�8x���,Q>9酣T?s�,�i\p�����W(��#��'b���	zr�%K� ��
?�q0df�������1# � �ZEm�)���J�~y�#�yr���<��r䈆'V``3L
*i� ����$G�`��I7��Lr�+�l�,��C���i�K�F}0�ŉ�7K�L� �DR6H�B�3N��B�b�$�R85�]��hT�c�. ��`�C�D���(ÒIx�� �!���rW�5SB�Z�L>pg�����Q1vmFY2eD�$"��o�6Wu�!j��M�N-���E�{��\+���!a�ȠҴ��^)ɻ��V�t50(`�^)Ns�|�K�hH��ʼQ��С��Ģ~�j�RbNǅü�S5��(xH4��>df9"�L�R�`8pr���W��r������G<opz����f_*}JGnQ�G�zMP�i��cV�0&E$s�! T	և`�v�x�%�	aP0Q7���C�le86��e\��*� n#��Jt!��h�g�#x�d�s��T�8	gB���0=)�Y�)�i�C�M8;�	#��'6����>2���#Ι4	�]"� X)(�a�۴!v~��S�LduŃ�	s@Y��#��9X.�A��o�AS����xс��-����[�*�6Ɂ��"(p�(cF�T��Tibh/W��ʂ�A��Mk�j��)Eу���C_�С&M50�PM�п\���!�eX�N�`2ւX�j��p�Q��2f��DS��t��Dӌ��̀$p*%�L�6Cz��P��0~�P�pN�0T�T�օ��>��+$���)�z%[a%τ��"�f��!z*�p�����'"�����hոK�� K��<;�����\">�H��T��#�.���㌜��-�H�I����Þ:?��ͧ'ڶM2 !� ]	(�iGJJ�EմAR��`���2O�!���
n� ��B�Ȗ�Wm�UHB�)%llA��� zҶ9u�@�"����Q&�遀MCz-I��EkN�QՁ��d��ɟ��tFy2G�jK
,��n���X�Fi�;�n(�V$���I�N8`�]ȶ�:P�Ԍ)�^Qꐕ#�фn��CuM���)5nX�d�
y�6@�;R���z{�B��CP�i�  �*r�ѱg����2�9Հ���	�}��������.�-�DX )�:������^��ؑ������'�ί	��S���
� ⁎��x��� �� ����K`�'��$����=Di�F�֒b�]Ac�0s�E�s�U5n�`5�@fZ�1��<���>Ju���k�Ia3�lݭҕg�^wP�Y�b[7e><0CA��Yp�Y���D*�d��Gb 2�H��O�Y ��1�W! F�"��3zD�؅���D^`�A��A{.@	��T\	��Q�e�|�@E̟R>x=��g�f
x8R�S� �:�d57�O2(y��!Y��1���Jp�l��냓�E(F+��z �Ђ$�l�T�&����c��4 9@B��B@eQ��=B��n��L��"���/Lt�'A��U�N�A�.�a������d""�ʓ]��dATM��Q&�Ԙ`I��!�����C�&�A��M��u��h�B�S'/M���Q�_'�<�D� �>�&��QbHC�EH�g�'�a���91'�R7�;~��T�@�V�p�S�Z�r�ą�g�J��u��U#�а���2p��nZ� qԴ�G��T���G"��u�Z���ʁzf��[E�8��M���+E�?,
�Io]�Z\�<r���UVԡ�/�;�̩�Ȣ6Ia~�I�:7BN����7�(��i�?��'b�U�`O�3��4A����2�� �$�~�K��d�œ%`Ӭ~�B��RN�i�<၈<mNjP��J�]{�E+�)̿��!�"���ř-8��$�?�'�~R%�x�\A�(b#��xF'���y���N� �!�\Ҍ�إH
=Z��T�Ԩҟkhܩ�-�
[����]w�Q�\ ��D�l�@FR
!�,щ��:|O �0�/|W�iH�!�� p���R��d���4�=�`.O�-�~�17ᆥ�5B�<3�<�-���'c�	�Sife�!�K�z`XuHM?u��n� +���C�	x��1Vm<D�xc�品4��D�rJ�"b���hE%�77[6p�M&+�4&����MG��'l����+'�]��.J&m`��
�';��r!N	��Ѷ�R���e�3O&�8

�nL ���Z��z1N2�/X�S�G�.~��d��c�%t�jY"
�u�bM�BU�GP���`�ҋ(N�@6��:d��p�@e��x���M�I$�� ]�V̀�����OX�9�	�#k��y��Ć[K@&-@��ϯQ�R�8��?�y�%��d� |�&cP�y{�@ʰ����~�C7�N�Ӌy���R�?�j�0��)s��7`!^x!��S-�,���V5��0k�C�[6!�í5�j�9�
.�"��Sָ?!�d�>��9¤�� �ē���y��xb�HS�'�h�FI+q"�Q�TE�J�
��'W(��eꇫ/K( T�؅\��lj�'xX�[�'[��j����۬O�4P�'E�9��g��eQƘ�'�ܛ8D��'�(@�� ��a;T�1ʹd"�'b\}�ƃG9��p'.D�$D�
�'v< �R�_�b%3�eL��	�'�$�SU�|��	S�k�y�8�	�'t�z���Sn���ҭB-uB���'(�t��/�9h��}c�I�b�}�'�����78_6"�D
3Z�6�A�'���Bs�ϼ@���g䚏_���'j"��%��-$��ǧ��<��P��'>�ɓ��I�+�D �f��>x�8���'���X��ʉ\�P�����p���'}
E�h���9MѺ|��<j�'��Z�81
�0�e�$�X�'�ȣ���7�t�:�/�,/P*��'���)u�� D�h8�ᝯ3�
���'|r]�#��),���8��Q�9H�}�	��� ��FK!$.rtH1�Ǔr)�4"O�=����Hh�׎�).�d�+�"O�kIKN�9�s-ȭF����e"Oƕ� ��E1F����+d�� ��"Ox�BM޷I��ȚVNų@��{�"O^4d��h���p�N\��P���"O�U���:s:��%m��b�\#T"O�e�g�ҹ�'Lϡb����"O��kW �9MZ�\�+��z|�a"O��x͐S��)���
l⬈�%"O�hA�+֖`��� C�mжū!"O챰�� $4�����U�6����"O@A#0㔣"Шi���ξ&�T�A�"O�]��͜w4���!ț��pLI�"O~�cg�n�q!�AY��P;�!���u������ �ȃ��
�(I!�^��I���3P�1�raɶ6D!��E�>�P�N-T����D��!��ƾ��}�����\~�3��#q!���]��@EH�[FF k�˞�!򄘐��cgχt<x1���7�!��:8�`,1�.߹�k��?�!��\(l��0�J+��ؕ�M�wx!�͋O˖�pU�P�O��Bae
2�!�DB�E�e�C@Ч.bd
��T�%�!���SHՒц
S1�蘱�\��!��j��!L�{��Q�B�!�$W�$��'C�#
,4���q�!�Db��ᲅ��k�d�`�8Y�!��X�k��Ku�MD�6��D�W�!�d��kӨ�# 'A4L\x��aC@b�!�D�s����ܪ I��C�B�/(1!��;?5)a��|;�$���G�[�!�D���qskѐ)���KY�!�
�,6� qpO����6e<iKE"O2t��aP(<důٙz�K"Op$�%��	�,��I�jh��"OZY�p�S�b��l�E��9���c"O��{�R����
D��pD: "O�D�s�S�Zg����" ��E"OB�c��ԫV-�L��R�j�Bs"O�P���-L�X|�
�%q~t�R�"O�XT��N�,�WI��fV4J"O��;�eH���$#iW�gA�}� "O�%��Q�SHe��"�"H��$"O��S�TҌm�2��6Z@A�"Oj���cO�y ��$�g����W"O
YV�̾It 	�W��6����"OJ8c���=nę�$*�~x,\��"O�E��(C 5:,A( "��q��"O�!���	!>��y Vl@�^��p�"O����5KqD��d+�35��d(�"OB��!�B/�J�(����Τ�1"O2PP0��o�P��7��e��H2"OP�Y����I��0:R��$;ĕr�"O���'���؅����n
=@s"O���ӹ���ڱ�� {��H6��Q�<� �A4KZ�����u�ZDH�BJI�<�1�#dP<�j"�é/ �\(ALR�<I�ܕq#�<0�Y�#t
P�e�M�<�%�J��R��3&Ԫnv ���M�<�����n�`͚g% �� m�<I���?A�< ����2lBni�<�fC����Y&`K!pz��Sx�<� ,��$l��z��T0���-�l���"O0Y�!ڱg����%�Y�jO�Q "O����ܙ�$́d�� 3�T��"O�C �-We,<"�`�xh�"O���� ðD�"EZ�!B\�B=;�"O��C@ƻE'���aЁ�R��"Op��C3?(���-G�V,��"O�`��H�� C�4z",�l�hM�"OnPa`mоu�� `bP/���&"O��:gW�̘3F���Q�"O­(��+YmJ ��@�'�
<`"O����k�+?1�x�P��<�lD�`"O4��f�̣J��p��O��ʽ��"O��!�$��X�D�NL\K���"O� 1Ƌ�Qz2�[׬ۅ#�`#A"O�(�R昷~�"G(�B# �(%�!��9e��U8Ԅ�0U%VDZ��U�!�нT/Z� F�N������ۈ�!��>C�b3V@Ԩ�f8h��EZn!��Ӌ]Y��.Qm��KB�O$*\!�dR=�yˀ-�'hty1�矽]]!���
��ˀ�	Ki@�ˣ�D�c1!�䕞Lmؐ�F[�.GI���ǋL5!�d�2Z����0$!T�2� �;!򄟣o���Fh u����.�=!�Č=@�
Yp�,�=U?��脬O,�!��(*s
`f 	L?Fu��L�,Ey!�^#8��l�f3�Xie��>G�!򤙫��i�C&��,CE D��!�d�;�d	ѸPd��!Ol�!�$Kh�T�q�cL���Q���6���ed:!�$��Q`in	I��߲�@���C�R_!�D8u�V�8b�J�a���b��WK�$�	"b�T:�(�)՜9ק��*��q� �:��G`އb����5"O�H����>3A�y	�T5D�&�"�M4j�^6mH3-�����hRSN�g�'�\ȃ �ܼZ:tȥ.܎Im����Ҍ��[�z k l\�y��|;qǂ>=i(���0�ʵ�w,NwX��`όs�|�ԋ	�^Ҳl)L?ʓ3�����͙z�X�D�Ȯ]Ը|13��ȬZ�@�%�%p�C�2�"���*[� U���'�y��oQ�/�5��U-x���a���&J��@�1�J���e�i����+�%+���-���wc�˅	�lM0��W�ض|���y�'�н�fc�X���H���u��Ȑe+��h2���u�L�q�f� ���]��.[�#anC�\�Z3̱��3ﲵxp�O�o0�xSc["3�y��a>|O��B#+�� �EN0tyX�����1'�E�5�_;jY�� f��#⟅]��Y�#V�HO|�l�02���j�*�:�k%��Xw���h���fk"��G��X�QGjۍ��e1V�Ԫ_�=�F.��Bn	�`c�g�^���IЂj�qz ��`x����=�|����|=Y�$.
Z�<�#/�
W���1� RG���`��8�j�P�̛r)y��.Y�̈�ËwT��o�8�^�+Eo���x©ҞƒD��܌w,��S��]�4ى�L�[���`�BJ >��Ԑ�iR�Ē@�u̝q!�4��h�ڿ�j��6*���ŜaoHLR���?��=�F�1����u�K1�reЄ�m<`@��
V�S�����I���F�[�~9s��L�\�lY�tZ�k3~|�uj�2U���۝'�5Y��Xn�Y��ŭI/�i�iŵN�
�B�%���{C�P]�@x��j�= ��QCd�oɎ�egϥ��Ċe���aM����[��I�4�nڷ��hO�)��+��@�$
�U���:ҡ"3����M7kO��#�n̯%�aR�[���|o�s�ڑ�ń�� H`D���1g �����1x �y�rF]&i��Kf��а>y*J)i�P)v�F�#$yP��6����6
�`#`$��i�}�F��T�B�b���GLh�h��#�iP"?B�)c1�J"CzU��o/��=9�!ה������9qΑ��욜}�L �a��	e�U�}ˢ���C� �0��$D{֡��[r�xh$�� h�iz�]�x������4:����-��|�8�����2���O�dj�C)�� M(aI9Z��zTN�8h<�̂h�;�N��"ѭD햡�c������ӏ�V%
�����(O��biA'�%��X�FPt Q�(��\IĂ!hu�i�a��&G���	��E.��v���f�	q E�1_��1�	�N��A�G \�
�ZH��cHP>��d:��ٝmG��	f���C���SJM'q����N>�#�ͦr��ř�dgI��C�jȄB���x"c�X��C�&_�Ұ<��$Ə�47j=�F1�� p�xニ-0���XElW�b�� �K��6<��S�i����6�TAVtŸ!&Ɣ\o��YAj�-m�R�I��׍`bX���7[R^:�$�5�1��.}R,I�#l�9�lʞ\
I���FȊ�jR�ݡ%ɮ�٠e�&����BH�6������I3�V�a���L#��3�-�(k�ˡ������t")ʓ=Q���G�H��(���;fq��38�b��d�H�z�|a0c:^�1��膭K���� N5~Ym�?d���x��<ZA��+jx�*��&-�]���Nc���@��4���&��R2ػՅěY,z@zs�Q<o���9��?^VX��E��3��o>5��i��3�N��� &Is�`�#
j�)'a :!p�Њ�Z;U� �k���=���A����S�ĳn�h!�EJ9A��C�ݓa�R��֦A	G(vjV�s2�X`�.����Ju�8@w�$ł� �c\�n�<p���v�J0��Ų�~��\Аc�" �a!�q��Θ4g�����8D*�6��7�i��N_���Pk@�Gf�P�C̮Tt���\<�p��W�5����e�L[ʣ<��G�'>;��-ͶL6\��dJ�^p�E�C��8&��@+��ÄO�,�%��$80��;r��7F*h�����|"��\�,kD��aI���"�6�։E����fU����d\��@�NƜW�tm��(Bd��*M�5!��I5��'?�ȑ
4f��&���3�Y�U�p���k��3?�P�C'�|��8ɲ###p%�`	�q�'��ı���b���+K\�"baS�eo�n���B�bʷ@� ���¼3���FX� �t#Ԉ  *� �s��(f��*p�5D�4���7���;`�
�kǬ:}����nK=*,9D��O~ ��'ڻ�8!C�FϾ�3w��?w���0� 5$04l�:u�r�*��I)otD�Su�G�s��f������f��>Q�lHa�J�=k@�:��owQ�H��
Y
h��B*¾G`�R'UA��5��+/�"�[T�'*Dx���[j��2
�AD���uGK 2��0�Ge��{9�2�j��A�V$j���~P�l��	�V�)�e� ��a�4g�}ܙk����8JR�J}^��gA�8u���(�!%��Q�䇥|b��������6a	'G 0���32}���cZ�Mܑ�d���J'���0F;{l�QmV'mM�,	�@�ּy等�):4����͋f�h�1@�uڒh��S(8֬pưi1 �YÎ�Qpl:͟b�D�ۿ>��\��K�]�xLZ�լA�����
�9�p�%��&v�P�2�>?��L�CGK%\�|���֑:��D�x�|�dK�����q��)"��d�LB�4��Oʻ��33b����%7Q���A�Z��eC�>H�.LZ�Ѝ*`��^tbV!R�,�j\3@�M+f\�4�d(㳪�3
zh��Х[30[2?�x��D��H�t4 f�яcjMv) :��б��)+tƬ�r��&b�����Z$�Ι�!��8�]8�\Dyb�K��Lz.X*�V�=�ԇ����3���MQ ��(�yr�"Jy���i�'�`Y�D��}gJ8��g �<��%	�jחlFaڏ��'���J@U�l�&�آ�O�cr̹�';|��A!X���0e?S�^�(�C��9dk�G�0��j	����5y�09	�U&'c^�{C�A/����U>���߷I���� �`���C%ź|��Bv�N�؄�	�s?�L�W�X�8A�;`�,�<	�k¿w5�`����4Q�~r��N�~�$���z�t�A"��F�<A"��[D��If�����,�W�$C��5�`�0��ͳ{g���'\��*2W�q`f��U�ňH�>5��'��ZƔ�f5dd��[8:�A��O(9�A�˱F���I����O�����s��	��K�	t䔹��'vℑ�/\	�ج�b�
8�� ���Be@E� .$!�D��>��ٰ��=V��(��D�H"����gÜ=pء��i��:�*�[$�d)�cH6#� ���'xzu�S�ʓLN�ɠ��֎]N\��'U�lb�F����h�>D;�恟.u���uM�
y6���"O�����+���p�'I8-z~�q�"O��
�@�O�҈�U��4T��p"Oؓg�̿P�������,����"O�MZrF��J�4�hC'F��@��"OL��DA�$C�Yrͥ+�6���"O��lY(�<��(,��Qu"O\@�(Z~�,Y�)���v�/D�8���"��]���Y�J^T�+�*D������:�|,`G�	z��k4�+D�|�O�"��J�)
��r&H;D��aedI���3_,�Z���2\,!�dF:,m�D���O8�)����D;!��.d���"aaZ�T,�<���77�!��8�Ԍ
s�_�U/�$���"v�!�D��?�p�3b��V��!%O( �!��~����%%�R��	�9e%!���6ӆ������tj���gJ"9H!�d[2�Z]� �=dN�!�B��� �!�ğ��`cĆʄ6-�L�_��Qt"O� >y��"�1���A��(~�1�"O�0��A	�2���� �,t"O���e�).�p�&�V�&��a�"O�U���ł&#F�k)J���"Od|#&�&�R$$�NM� ��"O��ƈM<LEF@� B���̕hg5O������/���!-��qX��&H��qY��6�\a��yrόN��X�0��<Ẕ?O�����	���۰����4e�Lң��X�h��J�7�h扤=�>�a�%ϖ@���r#�&?�
 LI�Lr�x��J�r�y���~���`��Q�덛|�
 D�4ƙ�40���̥����E�ӓ�M{�Іf~>��� �>_��)�'�Q��L��k!���b��dL�1@_�J����W?�!&ʧ���ܧF����p��O&�EK�n�������:A�@,���	�@��`l�"�0�8��H�I�9[s�L�xA-�L}��	�(k�����O�#�9���ՆS�b��6	�{��P�!��>!����̽'����d���%>
!s1ꜫq3X�#�M�O�T�I���>��'(v��%MM�c�\��d,�#?�j��r@ǩ��?�h�F��W>�*SNڝE�e� �0.�	F� /��0/�V�`ݑG��n&l����+�tL�I�RR��@��8EU��?�O���?ٴ�m���Z��W�z�ɸƠZi}r���e����v�|��)�p�	:!�5k�vࢲ�K� 5@lH'� ��Oa�t�Ⱦ&z���S�P�x��J��D�V��c��:��	Z8�'�~��?�W(�@n���T�4fP���������h#Τ
C��O>���>͆b��N/��=jDF�>a&�P�wx����S�%}���'@Z���t
Ŧ�q0�I�Ӡp �3�)ڧ$9^��c�[�����0��H��E9���I�y*�qO���P�"]L��
�
�Ј�&�&r��#�}��<�@f���0�n`	���3s}��"S�䲑�i-��������?�i>EvF# �R�O�k
`ٓF���kb4*B�m�	�c�$�`�g�)ji�aD�l��Ǖ;R����$ÅxܓQl�}��J~���v1��(�dL�:�-�cf�l�<��)� ~| �kģR��$Q��b�<����	�H$� ��YO8T�f�^�<iUN��jA
�#�)�#4K<��qJf�<��F� 2�Z�8�KE]�,R$%�c�<A���@'JeQ�E2mR$2LGw�<�,݆ o�E�AfWkd��a� Lp�<��f�f������<Q��0�w�<q&
Z-Qr��� G;kG�+bt�<�`�)	gu��� 9:�����Us�<2C��5C�I@��@Ɗ�2��m�<�ק�o�~!R���:1�4MCh
i�<AK5g%&�9#�F�q*�p��Kc�<�@�ŝ0�(a��U0i�����DUe�<Ym�L����qM20�x�He�<����;E����N\�0�
��WFe�<��	4^`������N�+�]�<ѵɄ� � H��=k�|3S�N]�<���	h�zƢ�o 0�2j]V�<��J]�_l��dD�&؋�,�Q�<9�
MG_�1���m&���^f�<�pU9x�ִ��HA�o��8%&�_�<)������DH(�P�`e͗D�<)�E˞xD����W�:�X�v~�<yѢ�o΀0���:)��0��.Bz�<��OÀ}>h�rq��U_�QD�y�<VS�X���"B�� E�2�Y{�<Q��ɫl�H�A!@�|j^ J���x�<)0d�8k��|ʱ*�)L�r�sbL�<����o���@�'[����&L�<��(Й25�`�Ԇ��A0��\�<��#ʭM;��Qrg�n!�#*f�<���1r�"��gb�L�l��'+�_�<��,�S.P��fE	�[�v���s�<��H�}]@�ׂ�5ML0�#�	�E�<� ��s`ƃ�A.������+�)T"O��@D�g5���&a�x�l�"O$u�t�?<�~A�����r��"O(]����"Y�2-�"�67��8�q"O�0q �?w}�$���S-��p�"O�y{g�T�U�}B'��*F(>pkb"O���!��9?>)�&>!�$cV"O��Yt'րoT��6�U�>(��Q�"OL�k�� 5 �E��`�9S&ܐ�"O��0S��G��`���KgF�3�"Oxu��Ď]Xb2DB��R��x�"O��/P� �[�A�D�\��"O��B�ֶ�P�A�)��C&�)4"O~ya�N�7�6[ph%\����"O�y`�'k���T�]:K���3"OJ�:�B�6O�{���!F��@`"O$��l����%�~��e��&�y�A��*Գ��ҵ�N�Hr�
�y���mV��c䂀+d������y���cMr�B2�������y�G�H0�x���9!���bR̆�yR+ۨ)ah
f�I�|Z�����yB�S�O��A�.Ae�y񨘭�y��H	)Ŕ0�" A=F�ea��y� ��x=:ȋɝ�|���d�^4�yF�c\����Ώi���%\0�y��Jb�p	A��ӧM8����O$�y��_�O|Xl�Ʈ�"z|9Su�U�y�.�_M|��P��a+�ԢQ���y�iӞH�h���JҪm���sR`B>�y�n�9#�$A�A7h����e���yB�Z�6hаpt	�N 4�׫�-�y"�ǜ<@�CDoɖ P.h�D���yR��6p�>r
[�i�b�[r$�yb��6��Yk�h��h�>P9A	��yҪ�9V���xǣZet� �^�yb ż@!j�Z�*��Mc��*�dx���E�P�	^��s��4M��}�� D�����-Qs��S�A�T`�M ��+D�T�ǥ�k�D5�FC�@X���Ԋ7D��@Xe#(�IFa�9A���2�J D�DZ �zHLU�!�H�E����'@!D�|q�I�#aġ���?&4�n2D� Z�L�P*� ���Rc�f�%D��Va=n���"���#ټ݊q�8D�� �Z�A��ձvH�
0�}Q�"D��pt�H!�`�Uk�V�ԫ5D��xS,���Am^����l3D�00#I��ST�aT��'($D�����a� ���DY�#�� �qd<D���Q#O	� �PS瘺9���p��8D��6+? �$ș��V�P���sS�2D��a�P5V@P��53i��`@�2D��B��,N?�aH,�Qr�Ґ0D���<m�x��_��V�f!3D����&B,{=Xy�7�E��7�.D����)�c�	p��*��-D�$��/�_e�`�V�V��(ց.D�`��fh��{����T<��`b,D�P�Ģ��73v��nף����F+D�(Rsf��nf��8ĭ_?�B���i<D��2f����(���k�&18�F5D��õ��g��3��m���� D��#CW�&L�:��ߋ�,,�V=D�� Ӄʜu��qE$[l̩ط"O|-Pcg�gWЍS��#d,�H�"Om����IRVp�ucY�QI�y�"Oys@� (eόE3c�U3g<�P�""O2 {���uQ�%�a��@K%Q"O�pb���B��q��0Zժ)	�"O�ը
W*1���J�)�>k���[V"Oi	�م|� $���W�,E;�"OR��W��p��9vC��t�:I�3"O�|���"�$(c�(�)�2�)"O��CA���͈�۳�(v&�0"OJ�j���u�6�sb�њ[��E"O��r1Ǒ�yլ��/W�"H�@��"O^��6*�f�rSD�n�,�"O<\i@��45l�C�
(\@aH�"Ol�!t� �v�CF�e��"O�$�$ើk�a��V���1c"O�m� (wV�r���H�P0�"O
DC�+¿J<
e��A�R6*�i�"O��zf"�! �ZA�`[5$��yA"O��*���*6F�1�`�
k�x"OT�	�#]�PLs5NZ	<�T4k�"O`0g������#� ���	�"O�`#��y����Ԙ`ƺ�8!"O��lO��"����	i�,�i�"O��j�Z�V,�Ťը��l��"O�H�eb�3Ij4���uʔ���"OT���(�5m�R�0�IG��(�s"OTD��Ǎ�eA�UZ�FQ�E{�P�"O���ھ��Aڇ���!��"O>5Z �B6Q���E_+v��v"O̙P� O7c�@h�c[ �"OD��횐T`�8��"�[�p�!"OP�A��	b��QE��. �"A��"O8Y�
\"fx�ԂRV�	����"Ot<ٰ��MLF��#�XQh!�1"OPMzC��7f��t��/Ш����"O 	���˰=���oͶ*��)"OV����$ծ,��/Лnz�+A"OYi�*-��DY�oQ�i0�'"O4tj'�,�"ix���Y�h�4"O�P�c��'�`X��C�*4�1"O~���O50�r��5M#�E��"O0)���'~�
��@�ޙ'`��"O�;�CB:x?4D8V"���!�"O��v�X)��E���̐%�}y5"O¼�A�����Q)tZ(��"O�|�4`�U�h�D�B8Fc��"O�RB�x8�mG,0]T�
E"O�HĢI�f��T2PjW�.�fxJ�"O����Ȋ#U��@�4��{E"Odm�W�Z
��,!#g�4kJ�0W"Oj!�@aB53�*���eG�rQ�%�r"O�=����E����d�-aM��Ђ"O~������}����*�u�"O�!:b���!�M���/s�&�!�"O��Ĭ�-I��HS���,"�0�a"O(�H�1L^��%kQ�"��8�"OJp��*�Q*�d>��d"O����%G�L����J�&��a"OPh�7j�B������	^HI��"Oh�y���p��S�GE$l�Ȓ"OT 1jַJj� �̗�f|�Y�"O�l�g▵kg���SI�h��5��"O�  x ���g���N�0(�P���"O2u1�܉2f,�
��X�v����"Ox��qC��X��[�؉�"O��Y�C%�)YE��9fघ�f"O,ђg��G	��+�&0}tSP"O���a��6�*�k��4�愨W"O�@�/�4@� �'�2(BS"O����x$�!�V��� f)`$"O����JNi#v�J%�N< �"OZYU(����ͳ!d?l�Tm!d"O���M5apի0m�>���c�"O��H��2O^A��
�x� h8$"O.q�D+b���"J_�S ^E9�"O��׫cv8SS�	�3�hz�"O�c#�3�
#d�ө>���D"O�4[���Oʦc�#�3�@9K"O��z�ꔅ4m���	<���pT"O6��͞?V`�hsq�{vp�1"O�-hBW�¦��2I��	��22�!��9"�Ya��	I�ݹRƇr!��P^�n�)d,�j�4��
�\!�DQ�5i.(����+�L��R��jI!��W����)3�JM�r��'	@!��	,+|=��'D�C�*o��"O.�s�)/���͞
�jYs�m.D�8�.ݶ^����	�gy�(�!�>D�X���4R Pa'o���1Պ)D���
��@(�����vs8��,D��(����b!2�a����f�{�k%D�d��S�CE�pu��t�Z���d"D����G�*`x��� 	�v�2SG D��"���92������@�m�0h?D�\�"I�u_F�0��2/��=�d�>D�\YC��k;	BS�̑6 <�s�6D��I.
;d��q ��I��Q��5D��(0   ��     
  (#  �-  �7  �B  �N  SW  c  Vi  �o  y  9�  z�    �  H�  ��  ݥ  �  a�  ��  �  %�  i�  ��  ��  1�  t�  ��  ��  =�  ��  / r
 � % i �% �/ 6 J< �B �H SP �V �\ Le �g  `� u�	����Zv�B�'ln\�0"Hz+��D��g�2TX���#Ĵ!�ڛ�?YV����?��抋<+��:���4.������uO�i1W@M4N��5ۥF	0A��q·�ݴ5뎜����G>2�0��\A�ZM*6�4<��Q�p+�(W64�dB�E1��� BM`Tr��u(�ů�\�Ne+�'w��&#��L��`$$��B�Z!�0�ډ,m򤩐�*"B�D�q,0`3%�%uF*�nڝzR��	̟��	��l��g[���W��x�!E�O�p���ɎOG�`{�eH�M���?9�'@3��J���?��f����T�(��X8`|����?����?���?���#��;EH|��1��c8PP�b[�'�P�ԎW�TDQ�b�@�/��	0��d� �<q7m�(Qɰ�� 9`��@̣MC�1��O�Il�'�d�{������.��҂$1����$Lh��Iԟ��	��I����I؟<�O[��)/��� ���@�cg�#_c��OR7͆��٣۴�?�ҷi���h@�p�Z99��ŹJ�<��Ş�x�ꔫ�`R!4ֱ��AW}b���y��Op����x����� �5�7�?�� M��X��ǁ 'TW���g��f��I�
�Vq£��O��l���M�����D�O��S}���*#��)-����)T�m87MB?1hd�sEȱڌ�Z��P��M�G������3�4/����s� )�m/~�+W ��!���v�r`��� l��Ms�iSxM�e�d� �h �L@&�����	9t�Y�g �n�<�V�Y����0f��5�4醆o�z0o��M��� NACѧ��F;�`�/c�I�@���9B��yg� zx2�a%�Ԧ����<3v���N�X���2,���?���4���8���d6iҴW��?���'��'�6�3������OH4na���ɟ��'��'E�GK�vK&}"A�	i�`7���~��0� jS�d�-E�̔*2K&O���q�Q;(���7 yӶdrs�TgE�����B)��{"nɔ!_��ݞ'C����Ā�pb���C��2����'�B�|�'��U�@��_��p�K�sa�a+�̊B���ǟ����^�>�$�@�s��S��?!%$�6r@��tIeټ�8&o���P�'F��;��x���D;�������yzn�ؖ�Od D�@��\�I�D07O��pW�κ�M�q����OVR�UD�S"�P��� p�:��بQ�#Z�X�v�ٳ�Z����� 1&?i�%l_M��vH�(#/�hx�d6?��ß0��4sk�>��'^'x���<�D�k���(L$���I�p�	By2�)7�ʬ��e�:v1��� ��.ў �I?�M�`�i3	w�8擗d���X� ��PLZ��G,P9T&"|mן��'�y�P�O]��'Mr]�@��bG�{�6�b��]�D~:h�H�7a\����4g)�,b��^a�q�/�N���״*�>q���0
:�JV�V#Qʞ��ܸ�@�8%o\�ƌ�8b�1��0;%�<Yt�!p(��eb���DBw�W�M�\����O
��3&���
/&�е�����IdH:7��q�'�ax��Iی	"�OK4>Jf�J�陼�?Q��M��hӜ�O��8~l 9)H�/V,�:���`�9�Ԋ�+�������I`y"U>�'vaj�@�h<�$�� ��&|u`E�u��v���Y��^$�M��)u8����Am��"��R���u�߷J|x���F@+���a�*�J2�MFMQ��y��${��9Y�7;,t��i�I9���Ҧ�ڋ��<	�O~IA�d�=6�j�2� �A:��A�'@�y����(�.��'��f� ���څ
��c�L�Ц��4���� ��mӟ��	+Q�!����Hp�*���:�nI�	ƟX;�^�$��̟(��Ƀ=Zt(��Od�]%� C&N��z��0��܀%�V��D�)Cz*L2��͉��`��k���!��`�ۑevN����e��JeӾ�o�˟@��'�:��	��R]�R\���DƟd�I�����0�O���'��0O�9h�Bߏ�R�����6	���j��r�"#<�O"�ȗG>��g��p%xT2�&W7��Z��YG�@��M����䧻Z�wt�qj��Ȭ#�`�M/(��6�'b%I�Fv<q�Ò���T�U�K�o>��}j��EQt�`�H�k�H��� �(��$�	o�X5�p�že0A���sc�h�2�\|c���Fp�c��{i��C�Vy�q�吟$��OV�o��ħ�Os��҆  ����Ǐ#.��}�L>)��䓲?����Ě>PI$��ņI�CqjG	��~�.�G~�A�O7-�O�0m䟸�ӬK�v��`�ը���f�Y�*�M���?)��X���D���?����?	��y���*	��2�NIk�c�g�!{t�y�SΌ�+n��$\=hx�%3-��i�p�HE�u�OJ�F�Q8n�̩:D�[�r������ ]��M��0p�5��
<?1�5 
�~�axÂ�rL־%��� b�9 �f�<QD$P���|����\�	�[����	ؓP8h�@���F�"ܕ'\ў�|�Oʢg�����i��{�`^ܟ<���M3'�i��'���O��(v����dԓA�!X�ÇIHTiB�M���?����󉊟!X��:���|v�yB�͇��x2�hǳULR�����>����N�|�lȗ4�F��BϚf��0�d�N
=�"Ty�HM�RBX���p$ �p@jL�'	N���E7sV=ٗ]0���Aa�>�?��?)����)P���U�ު�`BL�?b��d*�	�?���	�Y/@�����M@.�Ovdo�ß8�'�{�{���O:Y{E�J�L�C4-�fπ�=:���O���c�O���O��*�o̯ZX���5i
p��B^� �1�D�(���f݃@�Qr�'V�	u����"�@��X�;�c�g�r�S�w�apf�%0I
4	E�I�{�D�� ���+Oh!
e	FFҀ�o	HM�@)T�|��'5V����4}�� ���:!��(�����>᧼i�����)��<��dA�J�HA\ٳ�z�ʓr�Z���i��Y����y�P�%�4��ǔ7vR��d H�J�"�'n����� MiNT��ܜ��Ѐ��i\""0ܥ��͒t2����Tڈ� ��H�p�
��^�bơG������J
��$�OBP��C���>�����28����Op����'�F7-N]�O���R#Ao�,�b�ȋ{���j��D���}B���2D��������R�2N J�;ړ�?y��i�6�2����-2z��p��C�	�?A����ā�ZaV�$�OP���O>�2�y3�C��Ij�y�%a&(�Q&'�%1[(��`g"�+e����I�qOf%�RG!�j��� _��ʩ���;z����o� Oz���iܿ]�1�pѪ�钢d���.D��ԅ��0޺	1��-�*6m�ry�-���?��'���|�!ˠi�n��K��cZ��5�έz����8��؟x���W���{(��T�,��f*L<]
�d�Od�l��M��rz�T>]��}�tB=[qd�{FAO�l&@��B@��$����R"ar�'"�'|f�]Ɵ(��ٟLvlۆ;��2d� �,��ԫBm��-y�9��M��j"�T��4N0p���	[���m��-��"t�(�%�a�X1 �Z�ۓ��&s%��q�ܩ/Q� �+8���S�H�5<��#��N}�������D�<q�O��ӄ&a���zā.����'@�yr�D�
�t���ѽ.��9�w��+x�"Bl���I��9��4���1Qv�o�㟤�E�<a�e�lР�*BkI�~���Wy��'q��'N>�H3�/x�FP�S�^�%����ɥ.���]�l�����G	a�ax��8�Z�����[��z��}�VX'$Ac8l�	�#_�����'�6���?��O�5A�
��]%���V�M�(G�T���|�'BazRAS�|���C�Ŗ 2����O���?���'\��#'�h>(��0�2�h������4����OX�D�|B`#
��?y�F5	��o@#���I�l��?��)��䛣�ђ�6HHw`5�����Y?��OUV�󢧛����sG�31t�L��O$)x� �w$��"a�|0:t3��5�S��*��qń������F�3yC��F���	ԟ�E��5O�3�#M-N^� �ʁP�p��"O �+�OGQ�� P#�#0N�mA%�ɀ�h��q����}�0� �M��L�:ge{�n��<!��� �������Imy��H�!@���kU2`	p��ƀQ�BR@R'ؚ�؛-����Y>��3��v{x��q�M&�F1��]$2g@	� ��%'LI���c��a�<�Z��Bp�,`ƀT|�!� 2�l�g-�æ��*O��a�'	�đ?�O� @I�# <5��˔.|���2�e_�>`�ʇ	t�HZ���=\�Z�P�Op��@ަ}s�4���|��'��+PH+ѡH����,B�Qf�XԂ��*��D�O����O L���?����?��^>JTdJ�욇.���t��Vע *�FO=�d��
AJ�������{ex ʷ�ޠ<%��e��/H�<��cO.zt�Uʢ�V�nozA#w�	�M8@��A�y�ɸL��3/ͳY�\�l�E/p��3��OXo��" ��?���䓘?��J߀$��݈R�_�?�؅B����y���h��da(?�$�:)��?ɒ�i+"b�fIn�M��MԲ~w�6�OD�DЈln�:�'�"D����'K�ަ���OZ;�O��df>�Cp!	�E�|<����.��m9�z����̨=��@���
b���ɒ��%.��<٠�̱=m~�/�T�P��?DG\���}��jF��:a�9���~��ܘ$.2�>]nb���w�ɯj���[S�3:B@%��N�)��B��;YF�� %tpTi�%�M3����ğس`�'R]�ŘbBՎG���'f5�!:���m��`��p�4B��7�2�:�2�aɒ�'��q��D���'������G����r*���arN�~�ϟ�}K�C�8*fEX�I�	�21��������%.�!#��X��T`A`�w��9c��ia-��O���.Ϲ+�VD�'��y���?Ɏ���OO6�z �Ǐ�+��(`qg%1!�dZ,%#X|��J]c ���dg̅b�џp����õB\�!.6�)���� ��'���'K�9ɒ�)DP�'m��'}�V��:��*8�*؂Յ9o���rC*�6|�@A����7o:�!������R�,����Sm���Qw��S�αZ�ӣ���Q�˦��l4�3�Ɂn����Ⱦ(쮉�2Κ�W��l����䜕q��O��3�DZ3t*�ā2��Xx&��|���"�S�O2�sOų~J��1"��T�J���U���4YěƜ|�O��U���"�Ҏ~�p��V� %ʥ��>.�z�tʀ�x��������?y��ğ���>
�M2�@�*d.���#NH�xe�J�D(|�aC�F:�F��T���&�8���EO�� r(��U
��(SOC�n�,�у�Fj�<�x#�ݖ"�� ���Lh��N�Q�)=j=��T�J<�xP�I�G_\p�5�_���4m;�v�'Y�����I~�I5�~���Ĝ.{�L�I6�x�Y�ȓMM
)!�H�	<�iW)�q8����M�<�lEX��i���"��_w���'~d�"�FW�P�T�æ�X���Y��'��D�9`b�'��&�h�J�p���j�NlF�J�f��6i�7A�v$M;ۆ(�'�~�!q�ݭ3�� ����(I�p�d����.t��櫀�0<	� K�\����$ڋ{֘X�fѩqyX��kѬ3�r�'�R��	r��G.��`�>�3����s����0�;�I{����l�"ah W�O�P!iaIϬ3^�(jŦ%�'v�͈��'z��'��ӰA@Z���+\>	��:�L(@ ���M�fM���� !�Jʘ3
p�̟,ku>1��,U��i>�r�
*}� �ւՇ[ބ�S�K~BH6;�`�#�X�&4lT�1���p���Q� �+(|I����Z�^Ţ����b��O��$?ڧ�y�p�p�R�em�L��k(�yb!K,�Y�C���k|���-��O�LG�$엜5��X�J�%k��d"gkG$"Û��'�b�'C��1�mγ?g��'�2�'Z󮛢1�H�Ѡ�H 	�Ĵ�əZ�6�P��7B�ma���AX1�1O֜kC�O$���@�ܫ:�%�$��"�,����&J8�c>c���&�>7���P1+U�u�����A���M+/O���w�'��t�OH�O>u{�F=�M��N��>a���f�u�<�ȑ-{�:�S�#]�w�(�k�̕Zy�&ғp��F�'���W�t,��Ug:P��..�<�)R��-�DE���,��ޟl�П���|��f����e�tgN�$Hhx��ǅ3o^��/�-W|`8�dO��Y��Ā�^��rhĺ_�v=۲�[;c.��YfƂ3;�,�Ǫ��-Uv���D2����<KÍ��o~~��'I�ڵ 	ݟ`��U�'Q�����f��,��*�?��z��*D� #�`�RQ�ر6�� x�rź�'�d
����	Iy��P+\�6M�O��Ѡm�=��j	78�5���S;����ONM���O�$g>!�Vlؤ9!��"#.a��o�9r�Mk��I��I+�T���(ҠS$��Gy2FG�G�$�*G�WD�(�p�gw�KU���<��9B�W�DѤ�����n�����(QzܓUm���	���m3P�h�@X�5��@��":90U��C|Z�#�X ��11��b��Y��I��?���N��WbJ�9!j����x�I�E_����4�?a����I$^���$F�#8T�$DD)2���S�i>����Of��P�4m���P�92O��D�|/��,�J�+1���Z������3g??��.�"[���A�#��qxT ��e�Ɛ��Ѐw:<�����ڂ��#kr茓u�K�����'��С��6�6k@�i4�S�?�B�a�$}��]	'�I�&˓�?�����|R�y2+\��6		�^�4Rtl�4����O^N���4�?� �i\2'�"K܂Ж��jaF]��ӓ2�	ǟ��	<_�9��n�|�I������?u�%o~gH����	�|\K�(�o���d��mY�MzH�/#��t�|J>)�aF}|X�W�/��B���!;� �ԁ�*J����m**�|rH>��l?H�,�ď�lr�X��f ��8�'��p���?я��_='�j���Y.I����BlC�I�.;8��
i����q�<˓Gˑ���ן��'k�}B�B�1q4�pFWXӊ%�G�:�:����'"�'lrBz����̟ Χ2�2YBŕX�d4�j�:Z[��j�fhM\W�"=h��ShzӾ�;0D��Q�0�".B��j$�Ta�RR��T^f8�����E��X���O�Y�fM/~L\+w�ă?"�	� I_�#'�0*���O��ر�'����䓻=���2�mS�(���u
:Z=!�$T&c�L�RpMZQ+�,�'��6�6�dP�\��Ob
Ѡ�`�ဍ�9{�<ċ�jQ�*_r�'<�%ڷ�'��3��x�CdӾm��D��,?��3r��@�T ϔ p�(i�$�E�$�0=T&��(O�X8��<`���6/	;����W���٨T�J87V��R�.�= gl`��Q�}%D$Z`�4C���"-��ğ�	�,OZi3&��V��)�Se�(>��QB�|��'�^⁣ɉ�J8�ҧT7M�T���2B"�^ ���!&,ĝz48��Q����?�*OL��IE٦9��̟��O�v)�5�'*i���;z��a�ɍ,����'P�fQ�R6Jɣ�0�́�ۦ.j@Y`^��ܨ̟^��j$�h���F]!|�}KG��ī� ;b&H�G��w�T�c#�6/Y0RÂ�[�`K��Y�^IyCb�|�h���ox@��x�	��MC����|���R�#g����JCw��й�LZ�<��ّ_=�P2�c��p��q��Y�'���}��+�2K���r�L'hL�q!�M���?�2��#��?I��?����yW/[:"�ipTĊ.J�bi�q����
�h�p"��o,{*||�P�7{^����'k��Im����dKlE� �Aǃd������t��$@Ƣ0x4����H���-`�� t a�d	�Z|~�� ��c^��0�a'�d� cZ���$ݻ^A���ΰ��$`�̟MK!�$�)]��SRg�):�#s�U b8�"�HO�i'�$8�uIk��]�e���TAP$þ�>��ȟ�Iџ|X]w
��'"�I
8g�``�@��,�
K$���@P�r��	�#ӈ$�d����/fUcd�%ʓd����
SW��#o�a��Y��̭:���a^�1�Q��ޟ����� `w,e��	C~��3?�<��H�i��<�g�Ŝ����*I��?ғ�O��jׂ��J�%�A�O 셊�"O\8I�,O7D�.$AÄ-��A�p�|�,{Ӽ�d(�i>a�	?yz�u� �΄L�W���N��I埀01��֟����|27ʌ #@􈖅P�&Ť�͓OzPpu�A�p��d� i
���I�Io.<�I�/eL��3�q�i#�@�=q��C�H�Ia�H3��"O����	�'f��B����1>r�B�D��:B�	o�����E�wV� 3�.u����d��BcgZ �� �� U?Vq�E�O��u����ųi���'S��	J�x�i��P��hD�\��5�f�V�s��'���M��Z��qI��Ԥ'��u"��	�k��t[>�d��J�Y�4*ؽj�H{�`Vb~B��+N����'FM7t���[�O+����T�ۛZG�t/'"�tt��K(2�;Ӓe�����O�=	�'K(7-Zc�OI�ԫD��IE��j�]C3όN!��Y&v^�\b
��W�NA�g��3џ�*���օ� �2��Y�ђй0/�;|�7M�OV���O��N3d�$�Ob�$�O��i� 1$$C�G̍z��0�TJ�l���gΩ{*�`ܴ0�=�OSv�g̓R���#�(~.h�"�\J�����U&x`\S���.9p��t���h�a�a���|�A��M3�wI��pA�C+F~D�f$J�"������$��4br�'(ў�胧90�I�(��sv�T����W�<�G �+�<��6$ߥK��3eVxy�L$��|���� u��B�̕*/����u��B���bR�L�l�|�d�OT�D�O����O�Dy>�n�4&_x�q�Č.!
��I׺*���g P�`���<i�d�.%�� ��hC�\�@	�6���E�vAФ�����b�]��M{��3D$�ODd�@4@�޵���_�R�ݣc�A�i���'lў�ExB���i�d;�W�!c2Iqd��&�y2����0��O/��t������i=��'�� �
u멟�����@.����kݧB��j3N&����O�ɣ���O���v>����T'M��k�"��)*��7�l�� ��܈/������
1�@�G�aO�DLbh��@9~��U��X�o�-�:!�O�[q|`Jg�Z�L��R��]k����N�O��D5?�էI��<�����E�����@`�IQ����iدe�}r�k����Ja#�IZ���t�O��V�q�VX�&�Q�T k5�'x�%��9������Iz�D�-Pوi?�E��	=5���; �#���'k>l�p��L�Pϔ�i
��@��~�ϟ�a�ק����g�A�2;�TiB������͘uE����ܢ<B��k�ء_���w�+�BN�R���!�ϣoA"�@U�H~2h��?����h�J�	�d�z57�M� �C$9U� C��5)t��Պ��3U���뀦,��=���"����a�O��\<�šX3_y��sS�@����Uy")Û���'W��'��	>S}I"��7�t� )$ b.0�|��ϖ�z�f�H�ŌƜ˧���yB�Սu�����(T�r{���"U��Q�U��4C�ˊ,#U6�*���yR��7��jW K_.Ѐ��_��?��O�P�q�'���ɛ�������!&�0��a�L\�ȓҖs���n�0��X{Z���'/�#=�O8剑z�>��q��&��u/՝ٴ(Z'-�ϟ��I��\��fyʟ��dѮ^���XP&9R�4Hb��tW$I��N�2E,"$#�ƚ�!4�'���@Q�_��� ��\}����c"$cȥ��=:�����p8��9��^i����]L��))��M�w�R�D�O��=ю�D���]�� t{���aZH]�6"O.������U�E[���(K���t�|"�>q(O`���z�ӫ9��0	����rb ����$�����<����?��>���m�?�`T�%�*d�>��Ӌڞ{�L���� �~/b1���W �0<I����SjPHJ)5��Æ��=#r:�[`'�3��a��ŏ*-2)��	�:���D�O0�n��� Ŧ�;&`4L17@ݛj-.|&�T��I!ZrN�i D�K �a�cኞU����ޟ jd+�5S���g��g#>ёvk�OPʓ-@r@�,O��|�4�'0X��"�.H���䎎�\�H�G�'NR�S�{�6�ɔOX)Z���g��5z��ġd�V�3��:S�ٻ#�탒�5?a� ~	K�]'8$�}�g��,WQ>���V�#}ƴ�W��^�,Q�=?Qǯ�埐�Iw�O��� ���`�ˢ��f)̚y��cT"O��3R�o�6�sш����#q���h�ԴB�A�jf�!�	���zcDe�F�s��<9�f	����	z�
!��R��J.��C�88|�� �ҟ�r$�c��g�g̓L0�	�e�+9OT�9���xe:����eR�p۰c�qS���t��c�g̓]�ܪ�G�=JM T�f�ɃB��Cݴ�剶zOV���v�g�ɭ76�q�wD�5ft�x�T1q�rL��c��y�íɬZ��u�3H��M]� �'L�"=�O��ɥu@��[�苂B���ؖ��C��m��\��M��'�B��؛�(��@���BǞZ�p��<0t���7?h���=$�x�!G�[�L�pi�,�P����w��� ׊�� ����!F@Ft��㉪k
�, �Źyq�����Cc�=:3��OJ�o��HO�"<�!6S�h:������ȀK�Z�<����8}���R-*�b)3^�����<)G�Ϋ"��V#������S�a$�qgC�#���I�H^��hO�扉>	#|B�-��v�:�l�}�;���\���u�8,i������0^>!b���	���	v��$T�IqF�B7cF%Z4�:q� ��B�	�,Ǡ9��V��m��G٢I�����X�@��"&���b^?�����1��܆;Ո�mڝ�֢~Ⰾ��Oִ�B-�"�$a$LEZ~R4N,h�B�N�d>�Ia/�D�O3�$�Ԧ��}��J���O���D�HH�]3Ea��A�򩓱c@pYu��o(��v���m<���_�D��Qզ�r��	f>%�����R4��%�@&��rE'D���w�I"I�ȱ��]�e����d0��Y��>]bSMDR����ǛE��9󢍍�u��cy��jn�3ʓ)���kUn�ag�M����b�<�Bx��4j1O�#*��Q'@U�|]^Q�C)'�K1�����q�t�j�9na�V)����O`q�6�'1�1OB`��a��B$$���	� ݮ��#"O���k�#	ӈ��Rn��sm�
$_��؉��S����ؑ>G0M�0��G��oZ�B^���j��v'_Ϧ	PD6�7���U�������������;e(9�7��}��Y�/�Ob�c��O@�$�O���[ H졀�/�O}�����|JE��n
NXa "d��"	LD�'�~8�%�́�@�Ig���M�P��d�H�NwW u��A��nxr���/�4��Yt瞼=y���1i���O�b>����5<к�	�>�$�n�vy��'M�!"�a>����a�C.�@�<���5���Re�� (��
a͉�f�x�G@f���XdD�����	T"۾���Oxd!X/SeD%�a�Ҝk�n�@���O��Ka��,��U�7�J�T8�� B/Vt�t�S�5HT5ca��>f���CZ:;��D�(,�@9뒀&+Px!�so_�)��}zA��~���k�dԒZv4h��k��<�G�����	J~J~��O<*qM��t[4��d
�@�I��"O�cE䕲b��$�$r3�`�7�ȟ���'	e�%�^�1UT�8Ѕ ���$�O�-�� q��	�O��D�Ot�I�O }�vl�9"��D�" ��84qj� �țu%�I��8OF��Jȟ��4�w��#B�0 �mO��
̘Kw"�#T�7Ī��&Ҷ }�'��':�	����F>"���	� ��R�OrH(C�'s��	�<Ѧ&��]��D�c�^�A�)�x�<��"��s�^k'��/�5����N���t�'A�ɮ`�Aʗ��>f�e����r+P%�,�zD��_џ��I������T�I�|���M#K� ��1�	� �<�t�Qh���B���,- ��FI�|�����j�a��F<p���h�����B�����Z7�|!�o3��>h���C�ֈ9���y�2%Z�Oκ\�����U�'P�`��䆑2e`	�$,��Qp5��E7D�4���/5S��7���n_�	@cA�<���iN]�p�b� ٟ��'�柄�'h`�@��Ιg%�QRȒ7�ڀ�	����	џX�	,@tT���T"�`A���2D��' �*y{!1��UX��R�p�F|�V�[��ĸA��-:e^Q�`C g,�t EJPI��a֧~h��3��O ���'%��W�ex����_�#�l�ʋ�m��	C����^��Q�J0k�����:�O�'g��+��g9�@�Ћ��t�fQ.O�@�O���O��';R�����?)#���mJ�-�aԞo��]3�b*�?Y��?-��m��M��@��BT��8U&��w�'� ��d�˗)�i[h�$Hz�̓`�V��Q,U�F��u9����"��1���@��Q��K�:����3B�k�݅�r�'�)��$?� &����%�p�'Q&�0�"O�����V~�����	@]XW�
�ȟ6�!�bM�Ȅ��>~�HK�N�OB���O�U� ���D�O�D�O��i�O�$���׊=��<�`�r�\ã�)9�1�#.�,9̍P�G,,����'��c5$��S�2J���~�0ѢĊ�:a$�0V�^=p���4W���)=�ɩc��ͳ���wwʉ���D���g���	ştG{�=O*��pŞt��`3 ,Չg �t@6"Ob��6`��Z_<%p�kw��L���'�"=�'�?-OZ��Gn��H�B�W�Þ1�&E�Κq��١�(�O���O�����@���O�瓃F���WʙhI�vG�0E���H��ĉ[W�q���Yw��RT��T�'w�� 5��G����Z�w���7ȟ�?2�-9��2*�bE�aځN�џ�з�O�L �kw�t�0K�3b�ة���ON�=	��C/��=��	�Ifys�E�>�!�dU2S`b|I#���)Pr����]?S��I7�M�����uf���O���q>���y��ʆ�I&rՄУ�&�O25�!�O��D�Op���_Qw,pjԅ�G��D:e@y>�8F�ʽ1�fl��$�`p �X��4�=��̸ƀфVVxA,�/LT�';��(�NX�=]�cE�� �D�F|R��?Y����O.hA$EԪ0���JOOJY���'T����+?YWW�cU-q��ǿ}r�bdJVG�Ip����r�:�o��G��4� �=>־X�B�$VO�D�'��'�2�'_�_>I�ɩG��nK�0�.�RH�v�RQ�U�Q+�џl�ش��(a �@��p�6����h���Dx�O^pL|
d��1ЗB�{�̸7뎠k���'�R�r!1Ov�	�'�"�O2O�O�Z�[>~� �7��(�KL�A�ru�ƴi3B���`�r(�O���ޟ�^w�Γ�y�O�u_Lav�P2�������+��(�	џ�!�U�<�Zw5��'a���'󄜌�䡺�ŋt9�w�"^���h��'b�Aגr��:O๢ ۟�^w��Γy|XP�D������8#p<�#��I�nq��ퟴ3rGR>��i�O4�D�����%p���c�gV�I���Z4�Ƈ[���>r}����O@|X���O���	"M�8�s� �K�D�>������H�6����s���o��?�u\ɟ|�	�p�˩���D�O&�i^�R-��mٛ�h�J	�qy^�Z!�u������O�������y�I
���ܴV
����E�F���#��cH=)�H�]��?O ��@d�� oڄ,w
�ϓ�u��O_�D��h%�e��M�J(�"��Q�4��ڞ'A�·iQF7�矨��ß́���?����Y�����[�:i�`���!��˂�M��^��i�'�M�2�O��韾���L,R�)@s��7f4��̗R�<Y�
zjb�	 ��`��ͦ�����	��P�IΟ�	؟��	Ο  ��Q9\��9�U0 �� �ȣ�M����?I��?I��?����?���?q��
$oL�P�M�I,X�`P�+�V�'#��'��'���'���'`"덷wTQ�DI:g�Jq����9�
6�OB��O��$�O�ʓ��	�����$��,�� �p�\9P����`�����O��D�Oj�=Y�!aL�����+�L�DJm�s(������dy��'���'���?�сjD<���ѣq�J���L>J�V�'@��'�r�'�W>��5�CU@c�!F�οZ��ԫG����y��I&}Ɩy��IC;Ymv�+s�ȓ^n
p�"H�250��5S����ȓ��u)V
��]�dԳ%�4|���ȓ9X
y#� E�*�b�SsN�0����ȓ��d�t�2�v�rѢ0K0G~��'���'�r�'|�U�p)]�R��ROU�s������v�4�d�O��D�O��d�O����O0���Ob�#��,X"�T��@�o2Ze���%��ܟ(��������	����Iҟ��hG�  0�V��7s��i��D��Mc���?���?!���?����?I���?��b���D����'n亝f$���&�'���'�b�'b�'���'S�gݺb��仇E�7Ŵ�Q6%�x�D7��O��D�O����O6�D�O����Of��sO�
����qrH����*R��nZ��`��ϟ���П��ɟ�	Ɵ��0Q&l�S�o�1ZTv�D�+M<���4�?���?����?I��?����?�w��9xT)�+ �+�C�;�%�i�r�'""�'M��'���'���'~*EA1��XAf�a�N���;�o�p���O��D�O����O��D�O�$�OD�:V	أz���cOy�=�@��ڦ-�����I��X��������h�����{4ň'jb@�� Är��3Ȑ5�M����?���?i��?����?��?yD�ѫ ���^*E�y��H6L���'���'r�'7B�'�"�'�(�ֽ�t+�
G��q2�I-=�,6�$?1����D=�?L�ٕ�->dl[w�p���4#�(��<9����	��f>��`;�Ǆ�_Y,a��m�"C�4��P�ON6�i�ė��'p�fd޴�~«R�[�T��v�'nx���D`5�?aL�?G�$��ǜ��hO�l������p�8�ғ/Y;k�Bl�o�On���J��"Յ��'�� :8!OP?�B�lP�UC�@�V�'��'�ʓ�?ٴ�y�T�dr@��X���Uꄁ7 ���s�<��n�({�ށ� ��}~�O�F��C�����}�V-;B�Քb� Dr�ĘF��ٕ'R�؟�E��'x���TdN�`XvQ#�ǿ9c��;��^^��5����ۦ��I|�i>��D��3�<�x��������F�<1��M[�pt `�4���
+�`ȳ7&�)�u��Iqq 惀��^��҇W)�hO�D�<a��� �=��4�Ő^L,X.-��֦e�$!��?�$?�`�n�-Q���Q�cɆf��i�n���d�O�7�a��G�d�@�*�����)�&��&`T�C��@�T�����$èt��������&���Iq"?/��#��ь���x��4k��7�����e��.�����6D��� �<Q�����C�0�g�)�I6��EI-���E�b�����wL��b�!�1(AX�p �1�ns(�<�\I#R	�L�m�*!�z�K�+)� 1��ϟ�����/�&.���b��44��y�BgM� ��H9�,MD �Z�/g�p��k����ݬ�F�+�/�'R�,�X1����?��4 �(� ���)��K#�O?V��b�0ب�W�~U��I⟼��ȟ�MyZcX��$���m�l�{��F4Y}��c�$����Ms���ߴ��I�?l�6Ύ9����a[\�1��Ε<�h*Ox��f��U�֍Z���O�ʓ�j����!ug�5r�x|Yq��H���R��?���?i�mK��?i����9O�t�$��%R�k a:��qX̑�M�\y��'�	ҟ��B�4l�	��E�&u��Iңʑd^ְj�fXRU�Ы6G��?�O�ɬ[��D4h���AUk�f��Ɔ��� ��şؕ���'�O @ ��WJBL�2�є5�M�g�Od�$�O���<��F �Ճӡ�7����	�K���BL�O�2Q�1��\LB��~T�b
�.���e��&?6���UR{fdY.�,fe.�����69yS�%ǁe�d��0��
8�l�qn�8{f���&�� ��Ɂ�^�''̗I�԰���vv̩�h�&G�M��ak��5��!Q����݋G'^!��E�2HLQB�4���؄aX:+���9+3�0�𫐑r�d�9�ߐۺl�a�\�;!�([r�>TH�O@���O��D;���O8t��H؄^n� 	���T ̕i��d�O���O���O��'|��=;�Olx�f�G�Rk��;��ݐ<9@A�,OH���O���3���O���5ܟ�1��(���F&�g�@��'.��'Fr�'��S�"�5�O|z�\+�����v�B�8��C�?I��?iO>A�TwX��?i�=���B��3#x�r	9q�H�����?Y��?	��	i����D�'���G�Q~X+Ԯ45�!�rn5N��'4b�'2��BV�'0��'��S�y�t�����~:�|0q蟙'-N�d�O��DW�T��mZb�D�'N�TϬ<Aw��o��ص��>^�k΅�L�I͟�R'O�N���O��@���+�*i��LW'ǚe��'^��B�r�����O �D�XU�>'�> xтcKA�w��dmE��?��Ab������K�1ɾ�ؠ��{��	[�!�=[blZܟ��	��(�������|"��?�Cj�����%n�*?NZ�� ����'Y�XЉyr�'u�'>X%(U�=�DS�(�$O8yB��'����bvO��d�O̒Oʭ bJܜ�XD�P w����h�O��d��g���O���O�d�|z�;H�%���@02�D��k]a��Фό�VZ�'/��'�R�|��'�n�@T���j�0��0ォ#�������'���'��Z��0�o�R�)=yF�As�Ղ1b�����JHyR�'J��' �	ٟ,�	(G<�I�M6�`G��}�xȆ���C����'���'g�I˟ H�G���'$B%�t���Ѯ	��`ȺN�jHc��'�O��d�O!�!�䂾1�F�JP-Ւl��m��G�q!����O˓�?�7&#����OB��e�=��j�(Wd~|XB��
 �BH��>���OR���/���O@�'(q���b�
�%��lcdB�������Hy��Ҩv�6M�|�����pP���P�����F�*c��p2��O���O,d�p��O쒟\�I�|b!>o��p6��Td�2(���?DG��@���'Y��'d��m(�4�J��&Ԗn>����?x��8ʅG�O|�i3�O����O��d��<�g~	s@����Y;�4��£ȑ	f6��O��D�O�yf#L�i>e��������w���B�Ǘ;��4����������	�hKB��y��'�R�'I���káfux�KfD˘%h3�'��c��O�)�OZ�Oz��Q��Sf��pB��W�Xy!�"�<��%��?	L<���<��Ԋ�H��ā@����e���ِ��9qn����5%8
bf��V\���FS/ u��'�R�'h�'����Ĉ
�4���x��<j�P� �'���'o��'Q�']��'g�+ڵI�NY�� kt�eB�	�E��'��'2��'�|�M�41�U��K�)/��qHS��L�*e�b�'��X>��$�	��!Ƒ�?h���d-$����Z����y�������P�	\~�o��W�
5AX�N�Xh��7��D�Oz�$�O8�$4�D�O��P/e2쩗�Aj���J��N�$�O���7�d�~z�'0w��'>H{�[1]|�Pkլ�-G"�"��'EB�|��'"��2F�Ak��O���cܪb������)�,P���%D�� �+rô�~��%D��h�Y����c����%H�t��(C�M��E���E�
7����\-O<H�v	�.G$T	1�ښ�����E��`K��K2�@�&ot}h�W75'����?Դ�B�^�~Nbq_-,?�y�뇪��eY�d�* K��b��L8�J�:!L�L�l��#T�]v0P�0-�B�0E'�6N]�]�v��f��&I�):���������ןp�e��M�� ���х(��Ő�S��ܻ��Hb�!�.K���gU5�HO�s�ݘ\1豛�B�>JF�a0�4����N���`]���-P@A��i�k�,�b���]V�	2ט���O����7M$<�!��	�y�	y�R�,�M��S�S��?��FY�-�A��ӞS�oJm8���M�0���P�k8 U fn<�n��ε��i����M���?!(�h���/�O��Dj�b�g��!��sB�O�G����,V:X�ލ!���&l�r�M�!Ȋ!r���c>��K_����N����E��=|�7��+!����1�W6>�
��Ua�16�f�}��D1�����<BV`��d(�"�o�7?���O���?9D�ܴV�:���J
'V2�;���8m(����?q
�TW@�k�H�$dE��� 5��4Fyr@0��|��4S$���Tk����ly�
�20�6�3��'���@��h��'R�'�"+`ݡ�IǦY�B��) j�]+1A��Hh4-C���<�
1ē�.z@���@&ݴ맗(O�m�v��)zf5�d�ղ1�Ե ��?W�nh�cA[�|��*p,W+���E�'�ؠtN˿^>�(�M��Z�4�ҭO�����'J�7Cn�'��?jY�m���$\I�sdԙ~�\C�	;��՚S�^�ya�-ka�S�?|,����)-O��q�F�f����N?�6��#J1@{��ǯ�O���O��DK�G����O@�ӡwbDw	խM;ډ*�h�/`�t�7g\�77��bS�� �$ice�' `�$i�V��$���{��6�P
l+(�AS&�����
����ӂ툼3H"�;��c��	�xg<�$��	��1"��דEa��٦�Ϭl`ԍ������?�#��ON7��'N:��Y��+4�o:D�|��/O�3 �Xxde�tbl|�T ��`2�4�?9,O�6�	�oW.�?�IDX���"���e�H)��ަ��?���OJ�>�I7aP��"m��r�J�?��:��$���tc�C7�~�*���+DZb+I�H�Ȱ��Z�:�h0���yb�b��T�4c��&�Vj���ȓ}X��,��4�h�3r��8[êȆ�L���y���/� �q&+��K�A��|�d�b���|�a�Ѕ��6��U�ԥ�Pc��7Yf��	Y�1� �� ���qOR,��l�`�&s�tɄ�rL�����T|#a�"1j!�ȓ�4Q����>M�,��m��d��Y�ȓ �l`)�*��(��Ԃ�c��V^�L�ȓ55p�Yt͍:0w�Ur����)�x�ȓ���D
�Lmh��Œ;���ȓIXt�yb��gS:PRB�+-�||�ȓ����bǐi`��2����8��ȓ.�R����� N,�H�"qD�ȓ|�����,�8��&7��e�ȓS*�h�5@�C���0�,gҐ���A`�Cc�Z��qE31�A��`�������DN Au�W29� �ȓU1�!3�8j�`&�+��Y�ȓ+I�N�3Y@ҹ�`���N �݅�w��]��o�%Yk���-�:�ȓVBA�D�B84=SEL�O}@���]��	"q/�\�^L2�E�Q�� ��aۤ�P�ꚤ��=��"�mF*I��eo\DDD��4<$r�m��E_NM�ȓD(ʬ�!��#j����O|�9�ȓY�|=@B�T8� �c-�/Xf!�ȓ(PI���9{�-��L��a�ȓTB`��F`O48F��` /K*~��ȓfG��.Y
�����c�� ��L�H�qe0rR@��%��a���Ez��M��m騒�M�9(q���k'�ձa�`@YT��l��"Or]��/KV��b�JS��i��^����dE�8-�$%�O?�I�^Ȑ��r/P����a�FB�I�9��P�NαYh�}ҳi�L��͐��^ ����F��?�>t�$���Q�� &�*vϝ7<U�욦k�<<�:�:��'�p����^�]A�Q5L^"��X:���Z��*�14L���"��~"'E�1������R�l��˸'y2i���$:.��yvO�KPd��'Sv������8i0,I�K*l���O>�y�j�<���UF�,��]*����N%�C�f����F+w�½p�E@j��� �;h�b ���B�,��ـ�:GZ5�Ɠ A:xP����P����<��rd�&��p+Ī��x �+C>tp�0�B�m�J̇V�~!���ҹ3�)�片W�v1��c�7�	�DY�Cp�E��J�����'�42��XAć =T�e�d�'K\5!ǾY �ՙ�(G�}o�\jI<����(��́Tb�`L<и��?9񈂯����O�|��i(wCZ_��g	���y���. nP)�@٪U�x��QdE1}�P����4��
U�F@T���KG�S�F^�8�w�֐3��H���u�C�\�Dy�Mp�'刼2���5�V1x������@�*n�HK�N��RFv��Qm�:�n��FL��Q�<A�	�')P9B��N�"Q���Ũ8,OV�R�ʝkM��IP�!d"��W�$XjY�ʌ�Y���y�Q zO�h���I����$]-��䩶M[5Z��a�l��	5mۨ���M	8@�D%.�}Y�d��[�e
ܔ�3��6T�h-���~D���e+^���X�&�V���H!S���U���,��17K�{��4Z�E[	\�d���(�v�R�7(�! P���eΗ)-��)��x���F�/��bT��0�>4�"!�-6�a}Re¨ZoV�h����.w�y  ɟ�F��kԞct0��rg^���+T@P�y�\�i��>,q�e`��^�@��W�\y��p{��V�τm���C����(O��p�kE��5Wl =�ٻ�Oйe1�
�]`�8���\�p�>�Dp�Y������(�J�E��1����O ���˚�d�e�N��*ʞы��_����!���J�M��?f6��5kۯh�Mل��)ϖŻ�撊]���Aq�G) T�
� Z:�`I�	�|����871`A A��}^��s��3dޔ3��� ���W�?9���946D���}\�����2g��ݷ?Y����M8�C	?,���$F�!��Z���}�@��� �6t�$"��P��yų@�p���t!��P�(��!K��$��¥Z��"���j?YT'Ǖ=fhc�J��
�,yZ���N��O)ޥ����.l��V�T^(y�$)�������� 7`��[���'R��H*�mq����i�u�09a$��O���l��`z �A2L^
h���R��=[��"��ࡕg �v��@L�3ds�yR��\yL�Q犌V�6��dB�;��¬��0n�iѱ,�K A���'�6 ���J�7&׵���s�h{��,	7bO�}`zu���>6Z�h�0�K�s&���Fַ���C�%�祿yPj�T�6� E)��.!V�{f#|O@��B�վrj.���- �r�0�fE�W}X�5�R���r�,W�fBP:E�T]�*͡q�J/%�|�Ц�&TzV�EH����	SO(,�7g�Dg<��7><����'9��`0�ωO��dP�D�lzt��*��;.��/{��a��B�DB�e�� B�)�:�'[�p�2�ę�8$�D|�,ݨi&l��΂C��9"Sk�7�ڙ��◝+�4h���!1��h���]�j `��Rn�A��-�K5�ʽ�&�Ʋ^)h"�I�@�T r疀�~�`P�0?��N^9%����Ơ��G�u`P�X�~��c�n�P#��P8��X�����+Oh�X+�ě���-�96����À)>A�C�(üY��D��D�Ղu��H�`4I@��]n��  �����Oӑ�e�q���
j���._��a*�@��?��"�� /���G��$0�`	.$6��eIT�kmJf�0�@�*	b n�X@|\�qj�);��,��R!� �R##uS^�`�C%v�j��]0*5�5Z���TX4tBAa+m��rc<�b�0����,\��	L	'8�"�n�-r�$x�A)B]�ȄhҠíb�4�7̂6�.��1!�$� kX�O���A�&������B!���̘X<��ɱB����p
Y$-T�}j��@9��#����I��&dm��/�@���� ��%-R�aJ�;���]?Sg�y���	St�p�bírŊ�����Z��'j�8ZT�$b�$�EJ�M���zI�e�A�N!�Q�WY%E���c�'�}������M�$'���G�I!?�Lp�1�R�'�����d�;�9mڶ�nP��4�N]���2)r����ޒ@�J�ഓ�\����<$�D����'�6�sb�2���#(M��$�O2�􍌘�y���"C�5�|��Y!G�=�#���g�j��!D��G[|1���x2NV��4��4�97(fhhc��+�l�2�/ҍ��*�j�R�L���A�H�m�U��퍩cszE�Č"D� ) �/!L�l �Jl�x���O��ZD��$�B�O�.Ȓ4���=�%#αy��x��׆L���g�D8��{�g�d�z֘d����ph-����	9n�I�k��Q�ŀ>\O�]x����H��Ȟn�rUa鉋!�(4�<y��ˉ%� 0[D�'*�l�`�|7��wNڸ�y�@^h�d�fwx��A��hO�!(�gכ!�Q>���㕣#P���ˍ�1]� į>D�h{��L�᪡dD�<�@D��Mz�x�$�ڮ�ا���	" H �^Y0Ja�9��y�A"O� �e�w焋O�.k�Nۺ�:��$"O�h�2/M W��C��RM�ܩ�"O� ��� �+�F9�˒k_:ds�"O��1A�N?�4e�DK�QA�u`Q"OPU�B�Q�b������E|4i"O���#'ŤLf�0��7L�0#�"O�;w�F�5���q�≆P����1"OD\�&ޝV|L�;�bܤ=՘�3"O艘��ρ�J���S8e̲��"Oʹ�W��i����Af���>�{�"O�3�J�e�����A/Q��1{`"O, �'-:[�B��C�I�C���R"OH(�hαA�!¥��P{V��'f��*N�8l�g�,H��'�F��t��pG��&�
�uP��'�^tD�J�#�a&G�w�Lj�'Z�](T�vD����I��r���'��PE�+8�D����.g��Y	�'�r �� x�ɲ�k�Y�RL��'���G���Ȱ��ˤW����'�,��d24݀R ��A�|
�'u�z��¾yo2:#'�N;�	�'!�����Ϡ* ��5l$qh*5��J�4��4�	:���N�Ĥ�Ac>_� t��	���ұ"Q�1%:%:/��^]^Y�ȓ�U��G�����`�?�P��4:Ub�\~x��ѐD��*#����)ӆ���	ʗF�x��LJ�h��h���F�r󅔀WXp1����=p9����L�ڐK���@�Xu�H,��M��|�fL*�(��f��1�δB�\��=B2\��[�tT��Z0�0F@��Q�
%*�F��[@�0	��_-^d���o쩫��L�!�%N
�6����>��T�f�Q,'A �3@脡e���ȓ(!���S�Z#o�zy�����e�ȓK�Z�*󣗥s�\�dA�Z��p�ȓ<����+�kj�Z��̗ނ�ȓo\�\��i�,u5J�B��_(e�ȓ]�N���	HnM��2'�&'��1�ȓL�B���Y��K$�!����ȓJ�`�Ң�*}��q����wC���ȓ<t��V膁lX�4i��n숄�y�"m��1?��p��_�hz�8��:�� b�"A*3X��d�@�U�i�ȓvgL ����4�r6!��K�r܅�0;�u+"�o���z���%F��Յ�Tf��ɰ���o�h��0c�5}���ȓ+ � D)�yJ� R�LQ�w����j��x6�Z.^�\�P�)b��ȓ1~Xm�g/W�:A�]�('4��%l�# ͕�]q ��Η\�b��� (����l��nK�ht�чȓ	��gbG�zԄco�7Bw��ȓY7��`��\�f�1�U'�żx��(�HC��3%\t�;ӧ+c���ȓr�&0:�JI�PԔݎE� ��5�xR#�͵Mx6��v���#�Ly����\냧Ҁ�ő$(Ӈ=d��ȓ�n�����^�ApA۫+j�=�ȓs9�Tb@T�T�x�ۅ�*C��ȓN�j�#�ޓWP����G�4��ȓ,��vkKP�Y��Ʌ�T�B���(N�1�^K���*\2F�Ĩ��S�? ��bGN��h�<`*���M�6X�"O:��7F����ɲW���S"O��2�慤R�L��D��cZV��7"O�y�ĔBB@��aP�*V �"O
��4���hqRd�V�R�c+Z�C�"O���@��	7T�hC��Q����4"O�Y���o-��7G֯Rp2�3P"O���TH`i��K&���w���Z�"O���oً\QP	��j�g�b��"O��'M�z�lEaE"�/'��:G$(D��   �g� �S3��}۴���)D���d�	�Q��@
#
��vz��0�&D�Ȩ���.<R� ����г &0D�Hz�����H:���`��h
��1D�`;�@��	y�=ʂ�#8�|@,0D���˗�ss�5bU�υI�`T��%D�4�f`M�4H� ���dV�D �"D�4�c �J١�m��B�['^�!��>�4��#c�$4��$�!�
�}|�)Sވx��ԡ!n�!�d�j(�"���0�l����`!�P?	���#��Uѐl���4F]!�q͆���A�j�\Ex�-��!��8PJ�`��$��҄	G�
�!��01��0�B����k����Ay!�D�~9���O�]��"�	��>d!�_3	,����	�6b{�#�h�-}_!�d�Rc: ��
0CZ�K��Q�!��\8!ܠYX�fؒe#ơ�$��?�!�$\eDF*3�+q�n�s�F�/�!�$F�%�0D�5*ǩb �J5�	\A!�[�<l�d9���
b��"�vLQ�X�3f��n4�Q�W9.m 7��O@����K�b���������i�"O����2A�:�!҉v�nU��"O(!J��%\�
9kg��%�R���"O�5�@H�~|=�FD�p�ȓw"Otl��h��{�n�(#el�(M��"O�LB��T�6���.��5�"O8�(���3<�����z��Pb"Of�Zc*�8	P
����a_���"OX���!�<d1 O�o�(��A"O4��VI&Le�$��(y���h"Ot���*�m<�sc��d��"O(����SB� 	�+D,*&0�R"O~�ڐ-�*�q�Hf �\ �"O`ԃe(ΑY�fe��ń+%N�"O��ۀ�U?S�S�e�q(�
f"O�C#+΂wsԄ�5���4�"#"O�PP��	�u#w�Q�߬��u"OL��¦?d2��� I�S�XY#�"O�Wɋ4#���uB˩7� 1��\�<!����;�~ �^�;d�A�U�t�<I7H-*9�P
`@�!/�69S��El�<���,�����T�M냧�g�<�2�<j�"|`b���,���Fc�<�"��<�T����z �qʱ��b�<��N׆`���+�'S"y���5li�<AadW�eH���׍D;qݎ��O�@�<)���.hV��� ڍ5�ph�z�<�� Wi�	��Y	PH���u�<9�j�1<��a�n_�M����r�<i���@22)�i�'K���[ #[W�<q񢞳2���{�>x`�(y!�N�<Dm�P��ty�EE9;@��`�$[G�<� 2�j6�ժ��M��t#��"O�d��3�����%�qsެ0 "O4Y����Q�H���B�b�^M�#"O�t�ևU&��(���A�"��J��xB�ãh��zr�% mJy!q/�[2�IE͋�p?��=\V��C�l�:{ܙ���ۀRv�(��3D�X���T�x�^!�V`Z�a��4�u�2�h��Ԋa�-§L"�L�Í?b���������"sP�9�'Ɇ�@T����-g�9��^��}� �:�)ڧl��݊DO"!��8#�>Q,P�ē(7$�����;��t���Q�X���$_�|�I
'=��	p,�*$�>ʓP�i���UL��һ�ч�|�V2�+[�6d�yB#�����r�S^�����/�Ay�NOmg��4��N!a|��ѐI ͉���
���#m����;.���!DO�<Kl16a�y��O�L��@@���BI'Zِ�%1�!��( ��9d��,�����OL0� t �3!�<�ɴ��?��������נ�4u�S�,w)�Sv��+G���d���:}҄�mjd��&��+��O��y�A��S�X�%FK�o����ቪL��,�2v��#�a��GWJ���$Kش0Ԇ��"�\*�f]43����CF%հI2G�MT� hʋ�d�SV��0>9�O6��4�Ԋȕ܌���JB���k�.�e%_�D�����jL�渧�vF�U����Ռ!�@H��d�<q�i��Y�����(�=#&����g6��CЎ~N���=�O�&������%���������.Ay1�z(<��M�5x�q#��M}D`��(oǊ�'[z�	�Q^�˶nR O�n%Exb��/C٦ 9���'%��/J�p<��@J���J&�H��Y���ȁR����G�T�5hv�!t$��(E�+�z%K�(�Ob%p��N�j$L���ę6'����>���W�s�NU��Q�D�r��P�4�� �Q�~��H�u�Ƕ5k���=D��8�㏌)%��P�Ņ�y�����L���ɘV�J-�\��9O����|ޑ:��Y���	8WM6PcL�d�(����$�t�  ��	:}d`iU�ś���'������EѦ�z�E9� �Y���	,�p�c��4{�4���F�2��x���~R�I�r���ƦI�X���`�trt�)��$u�	�U��ȇ�	�>��E��o#7��x"�KZ�J̾��f��@����_�$%C&�X��AmK'P�Ԭ����mct�{�jU�S!�$UX�	��KG5#dЄ��k�f��'�Ѕ��c
�f$R���h��H?ɧ�t�T��ڽ��n��p�������
��?�p�D�X�`��v�� ��L*�KH9b9�B��:-W�
v�ل��S�Oں��5m�)u����a$t���"5�ɔQ'ԤPV�ɗ*F|��hkL�LIp�:� ��^W�	�q52$�!�b��X04�A�4���0'&~����ǥ<	S'м ��Kf4J��h��S���ΓN&�C ' �s|lA����"Ռ%��t`��;���"[S���Pm˥Jdl4�ɟ#��,�1�T g�pT��O�6U�v���/��5G��Jǿи�J�|*�'��Xwڌ��}.������]o9ٔ��|h�'1����΀�y�v(ٺKS�Dg�/_v��X/[��qŪ-9�$G���.#��m����v4�m�P�۷<�e�?w�=@��ek-`)a��JoKZ�q��#TiX���'��s%��Ι����0R%ԩK-Ov�9c��gCH�R�.�|!�]K��O���Z?��H&e��3�)z_L�
snQ�<v/*��x��H[Q6H� '�*!w"Q�6b��y��	y?���'�	_��EQ�w `�#1#����!f�Y!]P�`z��G�`�!�"�7b��
7�ߓ����&$B��D����c�R�\�J䅈�@����l7�ɥa����	/"TJ��,]?��?�'`�g<�Q+�G� �t��raz"���ū�;[��pk�%�$'���%��긱A�F�LpӓcB0)�׉X L�8LjуE�_I�(�'dp�Ъ�0?���0��t 8O��'ɸ牂[� `S)ʳ�T�H��׵�<u��KI�,�aU�=�X���,$�ɢ]VP4ٗ曥�?�u�R���T>�B�'��n̲]��*f� $,X֑�@%�%;�8�O�[��Z�mW9:-F�C f+�ˎ2�Z����6GZ��@q#�9�O�	��$1vT��ѥ�H�g�U��'D�P�O��c��`�S	_)B�4#LH����-M�:��|:�,� pB���壜*]����'DJ����eu�� 7g�Nݰ)AO� �Ef�:�`Q��X�w�� ���>�i���&�U�4Z^$��5��!Qd.D�� �� 5B���B��B�*֔9Z"n,�t�x$&�1l�*�ʧzլ(q�Ll���7 ؂}R��D B�/���E�(���(��)E�!s���P�?ĉ'��M+d�Y�P���C�%8�:���}b�G?v�򈉳��%d��c�^�p<�'.޲��	�b�L����ρf�ڔ�g���>�4�J�=剁&Z�%X��'jT9�2��i�nI-B`
鈴�U��b��>Q�$ڠ/�����PS�'-�L�B��2$�D�3�M�-��o�Z�"lX�f���.Q�\�2 � C���4�%�)ڧb?�1�Q�R (���aE�-UhՄȓ^Щ�R��0b��F��6~&�$�<�!�LC��X�%*��h!Qb�Un��d�,D��[V̝%���#�`p���%D�X2�K�y�`xgJK�dqd@@��#D�J���,Xvvu �'�6q�\|@wC D���@��Sa�	���f;pt�5�>D���WIHӸ9:�%��
���:D�����ŭ);:]Q��e���ǭ:D�К���	?�p0G�Q�{Ď����9D��"��@��xܓ m�6�x�d7D�$�iҲ8M���O�M\4�&�1D�T9V�J<z1���P���
�3�-.D���N�Tn��)���F��x��!D�������(��8���;��#D�� ���*i��Pg�PsmsN"D�<�򥔧]h�*&
�O��96�4D�$��nH�yi��a���6L�@zd�.D��٥���w�z,v��b��QD1D�X�7m���ҥ�V�ρ=R!"@0D���(�\���MΞ2Ȅ,2D�T�3��z��i*�#�uf:�"4�.D�8� �)ʔ�K �(S����G.D�䀃"ѩ])0l�#�K�z�Ԙ�TJ*D��R� �mR�ԏ�E�x9a�:D�pO� d8�qs��ANV�`H5D�tbG�ґLzt��.� q4R��%2D��R힅%L��҆��g"\���0D�Th��O�q��ؓ��s����DK1D�иrk�(KØ���Q�s����E/D��
Ѡ��z��u�P,;߂Qy��7D� 0Cj��V� �Ӡ�T4r�`u�b1D��@��ކPxRs�R;}$�c�9D�xB��F$3,ȼ�͐�U��/��C�ɪed$�2�-���Hp	4.͝QStC�ɷr;x�`K�/�@<�w�K�^+RC�	
���A�O�Jm���I*�C�	����i��Q�LH#i�B�I�Z�r�o��><��@�D�O�B�$
7��y"1E�����$`�B�ɸiR=�U�=X��C�,��~rxB�	6>dy7�� ����Z�?jB�9M�����6G�����P��C�I>+tz#f-&�ܩ�BO�Ya�C�I*.�y�S��_o��c�G�z1�C�	6D�Kw���X��M���bC��44A���1��g����IF�OC�ɟJ�t�ig��Jp�sʤG9�B��#L�Z-ȕKS 2�l ��B�*}�|�C���`��h�o3��C�	!�#�BN7>��PP�όQK^B�	�e<���l�~��@�D%�ZB䉁jv\�#CE���*��^�4H�C��6J1�@�["�y�ԡ� ҒC�ɂhUV�Ag��3k�Ju�_�h�RC�ɷI��M*���#[V�q��7��B�)� FU�5�V�h@z���`բ���"Oꄣ��@�O��b��r���"O���*L.	Cx��$�ʲ_���w"OJ�ٔL�1S�b��eY���g"O*m���H�=�Iyv$I-���"O,4�f�=�T��B΅q�b�x�"OH$a���l"���I���E"O�����ӵ8ݸ��E�lw^��c"O|$J4�M���5Qf9wW��"O��c(ɱ7ļ���7F|��"Oz�R��P����@���X��"O�DT�-^�މZ��6S�j��"O,�8R��F�ݛ��	�W�J貴"O��9Q�K� Ph�LYu�@:�"OR�i��Ǭ%�z�RSj� F�p}��"O́daT�>�0;�hS��! �-�yb��-6�H<�F�A/>@@Y��7�y� K�|�c`�<א�B��\��y�؁i	�偂d4Iؐ �$ʭ�y�BA]t�-ua�(q���8}-�ȓhѮ��G��6���k��GGV��ȓ�<Y+���=�!�G_�b���ȓ���"��W�B:2ѐA���!j����1(���El��p>�h��*��6O�|�ȓm:�c��F����K����X��a2�[!~����f�	�vu����4�"J	'XH��3�Θxl�ȓX:%��׆A�VԪ(����a�� *���(0|	H�}�ȓ,F�;��O����1ˇ�wg����ޡ�'i�Xg��#�?|��p	�'4Tea��7C�r�n �1��ܚ�'��XH���#��(� �ɾw<���'�.�; H�9��Q3��tl�8
�'֦�!��1��Yb�F������	�'/`$Fܺe��}��L	ȌP
�'H���ht`:��E�(>�d�	�'\h�BĬj("�)�a�k*9	�'�q�sa	�W�)	\�؋�'����U��C�S���}��QY
�'u�<qRc�*'�QѢ��6@<���	�'{b�)�aR&`���Z9����yBlݺx<Æ ��j�YB+��y��Y��БY���*^��E)�V��y���s;8Q�! �N�L����y2+!x��QF�[�B*j	s�V�y��%��A[��D����7bM��y&L�,�9��8��8Hd��y�K��p1h�>(&<�p��y�#��=ڸR�1�V��O	�y�M*IpP�G�C�$��ݻ�M��y	;Wwndz�`� i<с ���yr
à,�6!�fa_���p��bϮ�y����<�q�O
=�i�@�ߞ�yr���] �F}ߜY�h/�y�B�>��!�gb�$
�*����y�$ 3�ɉ��Q�4ܔ9��S��yr�w��p��
�wT�U��ّ�yR
H!w�3E�Y�uu
�jWo���y���d�4E� �]A:����P��yҭءu�I@�X����գ���ybf�蚠��ˮP�| p%!Ҳ�yr��-	v90�Աyx5�գܗ�y��LF@�| V�M�G��e�+�y
� u�C��{�P�;т�N��0;�"O���	�O�m+�"�rn�xa0"OFhR����t'��JR��I��Y�"O�!Q
! � @ǂ��2PU"O2��X晘p���|�D��"O�5��-A9�$�iW�T$n�8ȩu"O(ré�/U�]��(Ld�~�(G"O6�KfB�4,^�@z��� �6*1D�0�Â�8�����9rSl`p0�+D���a�4��$:C�G$v;>H
W�*D�ԃ"̊�M�p�Gb�@6�qu�,D�;B��9&���KDKD0J<Aɠ,>D���Q���~/�A��֋2��[a*D�(���ȹ!��`��ծ�ȅQq�-D��"L=w[�(Y`/'Vё�L)D����[�#�b�P4	C�{똕�UO%D�����YIb�	�A�lI�Iۃ�$D�D���[�"Sh�(�g���֨!O4�=��K�F�b�βs���RF'B~�<�a&��|�b�-�+;��|~��)�'Q�ֽX��9w�P�`c&W�J��HԖ=)#���,�q2������HFr%�4m�<>���5<����c�t@���k��Q�A�*-B}��q������˅eS~�[w��"�x�ʓ�%ȃ��#	^�SslܮH�FC��!j��u��C�h�j$�X*^C�ɝ\���`��L�_���`�?6RC��Q���s�e�^�9��F`�B�IE��3FI��!*^M���'�-�3%��z����g_D��x��'
�ӓS\ņD�4NʇG��'&h0C�I��/':,�����o�4Z�'_��������X�ٛ>���	�'"��Rm��(4�a��
�2-����'_��H` ���KD�%�&u��'���� �oѰd)wN@�Y�\��'�d��&i�m�Xa���X���'���k��Hm���e�
�x�����'�:���Ў�]�`No����'�@��-�.|F�@k\�
�'}�����Z�;�����]��|��'q�E�g2&^2L�4i�WR�2�'(���/��+��@�P	�}bH�
�'L�E�8Z�4h IzA��"�'=�ܐ����Y�̋�m�d���'�"$�0\��3@�hy��')`ų�bNE,}��][�$j
�'x��đ�tp�`��X,Z0R��	�'>���(ǵiMJA�1�X��4	�'Mn ��ݻvxh�a�� F���'�Ԩ8&�M+aS8Ճ��رA�qa�'��xh��8�0lɖ2P���'��cg�A\;��W�Ɲ#���'��4���F�g�4J���X(�',�a��<UUT ȶ�ƵM)���'���Ra*9��IcHJ�U���R�'h��CY�:e���"GB
J�޼��'���A�<R�J���/��RW�!j�'pL8�p�É!{nܐ@슦BN,p
�'�pX����!�b�hE	oF��*
�'$�;���U2�݇>�|�i��!D�P�@��%>� J%$V�z�1�=D�\��ֈO�#&<��iQ$�&-�xC�)� PiS�Пt�B�iЯ�"B˜qr�"O�|C#nI�<����M�(���@"O^���-N���aQ�0^��Se"O, r.B	���M+n~�!�"OLi���S�4�A�Mf���"O�9��"_�Jq 	9E�ԲN����"O�,C�!�`��&�+Dpx2�"O�d�2���oCڔ����5)���#"Oԭk�D�M*��$_�f���3"O:(��j�Hk�:1DͶp��@�"OD��
��T��1�A�}��"O�v��" �xb!J)lƝ�G"O�uZ���,odt����cK"O���m�{��Ȩ�Ƒ��O�*�y��M�8�0S��v3����y��C�P�x�S��#D����dS�y� ��R���[�>y,x۔�/�yB�R�p>��)&��7�ʩ�2aհ�y�R�G�n)����2�@1hL���y2��^���qlՍ
vf!#��ybǐ8R{����'	����y2iM1M����e�l*�1��6�y�_!!�:]�#.ǉ~z��5,���y����~�z��J�jY$�B�Ф�y�l��\�8#Z�dZ�1����y�
?U�XeS�+IM`�t���y��8�6�{t�KTZ�N���yr
�'):�Z	��nUb"JG��yr��<C��G�~�R�8��Ѳ�y" �X{��"�Οu��պ���ym��S�e�p�5�DzrJ��y��w�PY1����h��R�˲�yr�C�Ȝ��o��Ԭ;��\1�y�<㆕�AjSG��;qF���y���d�\4Q�eT�B�x0L�'�y��D#�bp��۲�S@ _��y�DѬJ"D����'=b�X�ӕ�yLA'ROB���`�`l�x�+��y�'�!E:�Lҡ����!fKE �y2�̅[������
�ʩk`$ϫ�yҢ�j���֋�\�zB-��y�ʌ[�����J��ج�y��G���H��Ɇ6�xdR��T;�yb٣A��#��_���%���;�y�Z>t!��3e�yp�eʡ�yBDߧ���(�	�� �F#�+�yb.�J�(QC��	�XtF�1�y"m�4���G�L~7�:ՏU �yB����S%���y�@`�$��y& ���e9JC�?l`��À¸�yb��)���k��#-ք���Z��yBK-	����C1R����l%�y�LH�]�P�҉�F��a������y�J�SejA�6�A@��<[��݂�y�ϑ�4$��E	؄�u! �y�^+,��K!I� �d�#��K�yr��"	�$!��(�q�İ���?�y"(ga�)�)pX&��#���Z���q�'~�c/�2v����ǓM*���'�BUS��\	�,)q2��G#ص��'%Hax&�fgΤ ҆F�X���'^ �sCj�	r�e��A_�`
�'�D�1��ے��03����8�v�1�' Y3��cu4�[k��5]�
��� ����V��c�΄�^�Q�"O��7JO	x��i�%B�V����"O|�TFҎj� ���I3Ov�q�&"O D��� �{�N�b��j�0Jc"O�q��ÙgQT��ÉJ�a���"O����U4��\� �K9֨���"OF��F@4	<��R�Z 
�v1R�"OI�@�ƜsU����'�'Ro.�2"O2P: ���3>�e`�!� gZ�2�"Od�rs*�
nB�9����> �ꈱ�"O���������*w�<A~���"O��r�V�O&�9�EEO}b h�e"O����Ô�M�`��T�ƥ�l��'"ON�3'3��)
F�#��� U"O�1`�CY�V�	�	�1�v� "O:)2B�W*|����=���A�"O�t0A'�86����֦D��B��V"O��"Ģ��u�HY �k��D�jh�'"O>5�ɜ�^i�y�
9F��)8t"O�(��I?ez##G{�Ve���/D�L�q����$p�f ��@�ܙ�V�-D��{���"z�zHy���$B��;�,D�$��[!N�Sw�L*�puR�<D��q�	�2iэN�c씁��"?D���BL].wnR��SjȰx���;��8D������	00UI��	b�Xi�)5D���ʓBH�=�n�;� J�o2D�d�a@۽(S@b��@ZC���� 2D���CK�<;q�]��Lə0MQȒ�.D���3!�1÷C�[-&��N+D��Y2Ϛ+�n���ǕA�Psgm+D��wk��[Sv��!�>��}��"'D�\��ϳk�� #
_�;���h�'&D���֙K �CU�ۏ:�<Xش�"D��� iԀ<P!�.Z� $�s�!D�x��A��N\ڠVƃv!�!��,$D� �/�Inҝ��-Cavt��c�%D�̒$Ȩ�Z,c䮂�=�@I)W�"D�x�(1_A�q�V���L�q�cO"D��!l�� �F���$��Q�VO.D��zP*�a�nl��S �I3�,D�P�@�͹��\6N� aA)d!��[qtMz��) 
*�����)�!��בy3v�#dL�d�BboT9c�!�DV	&8�M�P�	������!�dP�#C��:d*��+�Z=2GJ'\�!�ǔ@2�����"6�<�� }�!��,n�ְ��$X��J`Is��$x�!��I�;>LP6 �h�R�DT�!��0~EH0�t��1fp0�b�X�!��$^|")���O6.�>��5�ک �!�Y�_Z� �V*�%u�𥛷�Q�*b!�q����q�ܿa�Q���3BF!��ڛd�V���*�|���G��!d7!�䃻U��鹗gZ�4��))$!��39m���-�8Z٨�H'
�!��"{��!���+o��t��.W10�!��M�Bi�d�G�0؀<�p���9�!�� �j���R%M	u��4j_�6�!�DI� �@,�a҇^�zT:"'�n�!�3�Q�%iW;q�9�--�!�$Y
{8|��bj�N\���1��<�!���y�ҁA���@.<;�lW�b�!�D ���Q��@ '.>0�D,%|A!�� �t�Z�yw�huAI�|�F8�"O��!�h��9�G@׾�jң"Ov�8�� px�I����.�FhK$"OT=���
**X�r��	;��}� "O��y̢8���RR+�-��D��"Ove�W�K�
*��IζA�I`�"OB�p�j�H�X�"&������"O��a�ߗ������G�"�"O����/��%�2��8m۬�0�"O�$Q���n^%Q�`J�C�Mc"O� �KZ�HF 9`�H�"OR�� ��>0����̈́=I�)C"O2A�e�i�@	�Ĥv�-p"O��S�야`{�1ҡc��Jg@�(A"O~��4L�2w.�c*b]0��"O>����ӭW�b9�p̑}>$д"O���Xi�X�3��!'�f��S"O\$ � ��%�LT�1��(x�H�U"OD�׃ߕ�)�)�
��!�"O.h����-3
�!x&�J{�iD"O���4Փ�B�Up\]�w"O��+$�5} ijK�8b&�b�"ON�K$��.]Y���gP�'=:��"O�y�m�  �B����4s@"O�e�6I��Di��Vg�jZb�"OZ���ʡ,��D̆c��*U"O�a#!�3_�p�YQ��7}킹��"O,���Ã�	�d@Q�h��k��5br�'B!��D>~� bv�УU����Y�!�[<u���'�Їoqd�w�K:|�!�䚙6Ἄ��S�	kt��"ę#�!��bBp�w��|��}��b�'�!�D�
��a$�5֌��W�W�!�D��m�D
�!���9jR�$�!�D����c��j`��;�/9ao!�d�,�Z]���6lMa�U�xe!���:t}�qe��"g��V���YT!�"f><����>c��d�8!�D'pBR�B�!ѡy��d�d$��/!��W]耻'j@�}j�Xs�!�C�c�i��Eɺg�<<�dT�8�!�d25<�����϶@�����-_9z�!�dZG�.�s#�N)&�N���f�@w!�d�s%:����� -( b�d�!�M�h�<{�ڃE!XS�㟺F&!�D�	�d\	ө�'v��9a��n!���%l�܉B��:K�jA�CP3@W!��Dae+����)�ܔ�Ƌ�R!�I}��9���8 |�@.=:!�DUb�&�@�N��ba�ѹ�k!5�!�Ā ���F�g`���K��i!�D�'_d���k��� 3
MSL��d�3I
D2�������TJڦ�y��"Z6��I� �#{� ��^��y�Gۓu�t)�eE� V��y�Ղ�y��*XA2�"v�${�����@��yb����P����rdqpgH�y�nFlA����!h��"ñ�y�K�&/�%Q`	��ZA�8�e��y�˚�qu�0��+ټQ�f��">�y��N��8�N�2�� �ς�y�6�΍���	�=x4S�_��y�D��j�d��V��0���z��3�yB[!
X|�Ȕ� ;�nubf�I�y
� �ڵ��3����`���jf"O�����c����3x��"ORu�Ђ���l�㍋���B�"OpY�'�
��taȃbM�T=�U �"O&��1]�
�����X�*��9�"O$e�I�5�PE�e�?_��<  "ON�Q�!;+^��Q�>ao���a�x��D2ҧ(�̝��Z|W.1:��޼w`���ȓ
�(5���ߋd��K�$��~�u��X�F�w��3 ,�)K��̭g��لȓ%�0ݺ�n��S3�Q�� \�=@p��J���%C��L��P�F�hޤ��z����y�Ft��6V���Hab��M�vN��@5/�d+�܄�Y��yr"$�;ލ�iw">��ȓC5l�Yt"D zɒ��
�6��t�'Yў"|�D��-h�h�b(خ;���J�o�K�<��	*z~��a�
�)5�t��fMD�<�rLà.�iA�HЄ{���!�h�x�<Q�a�
�p��� ���c3��u�<�G�U	A�fyS���"�X�/w�<���0� C!�Ը#8�DH�Gq�<��o�(#��)��;j�!�`ąm�<����2$d�CgE9
��Qk0m�@�<�C�st���A�ش�N����H�<���]�����+~�bxℍ�M�<�E�e���jR�������L�<�B!�2<��-q�g�f|HYcFD�<!��^��z<h�iխUp��&��|�<a�+H�D[r|0�D�&W�fp8v(�|�<R��9�
�8E'�!Pq����w�<16Z�z�x0M}�\�!PJx�<Y��E�(��C��0��z�M_H�<�1���AE�@I��*�`�E�<���Q["q�'��"P�z�Y���k�<��I\�	��L#�H�=�ڭ�A�`�<I$+Y�N�԰X"���f|��i�__�<ɁA^��"�)�@M���@g`�U�<�!��3�9x〒+e��9��LL[�<���]O�Y�1�G(¡�׬�O�<����>�&a1���Q�P	��l�L�<A1XI1f� J �����1b�<Abn¾:m|�+DfV<LV�YTb	V�<A�A҅/��R��դl_B	8$��R�<�q�S�1Î�2HP����QN�<	e�ш&:�X3o� -�Ll���H�<)�Ր[,��1���3B�� #G`�<1b��oT��"6D�@5�E'FD�<��E"A�� ��.	��
��&�g�<�u��Yau�ƪ��7�0D���`�<)��;72��`v钲⪨�t�d�<ɑ�۱,�MpeB��>pk��O_�<� �� x_@�I�)� \T��CH[�<���'6P# C�
b�q�C|�<�eC�+Ix����H����x�eGy�<�5�K�Y�0`�#�@��S�*]w�<9@ۍ����nK3�R�KG]�<I��)�.%�HM+	�L�Ӆ�R�<�d
��|xWc�O$��U��Q�<�T�u�q���	=���k��x�<!V��8k$N�"�cA�j/u��@Is�<�!ǋU�6d�T�G29\|�`�r�<a%��/X�s�ĕ{n�u��H�U�<)����\$݂G��]�å�W�<� Nd�1�ްfG:���B`x2"O 8r�D���6�U�L�(V"OL��bEV��Ԝ��	_Z��!j�"O�����!Z���Y�I��Tv�mY"O���G�E�\��s�"��Ow�H@"O(�9%o�5>�9+��Y�Z�c$"O��I���H�&-8�/=lP��"OP)sR�G�ʽ��M�5J�@��'1�h#S�G�3�.��&12)� ��'Y�Ha�U�f�Ԅ�GC�/w
 ��'#�)�$A'9| ��� ���S�'�&aP�J�Mv � nV������'L���&㉊F}��������p;�'��!2Ѭ��@���SE@C�_��Z�'(P����&�6�JՅR�/0�0)	�'�A�S!]?ul�3���)�t��'�
0��Im�`=8$�Z�(�0Y�'1�T�g�C�=l��i���nf$ix�'����.U�#��u"r� lބ���'�fq�`κ	�h!��L؇w�}
�''��`⑄	PT1�%ŶW�t�X�'���$�U�w�^ȣG끠:�Z���'X��J5W�?��P�A�ͧ9� ��
�'����N�(��L�Ə� -�Zy�	�'Y/}��3`���wl�)hLD�<iЫY��US6�܊9d����EDA�<	��4�d�4,��"��EM�@�<�bL2��!CF˛���Y��f }�<It��@�V�c I��ŒQ��c�Q�<��"E�u(����X6P1X��Q�<���-����
=7�! ���r�<YQ��*U2��Q��:H].10d�<qBB�z�����L�D���&�b�<C����� ė�(�����[�<��L�/a1f=�!�I�|�H�r'DB�<�Bn�~��P��23.*�)�dh�<���U!
�������X��!�Ȗy�<yCB ^�������PAIV&y�<Ys��>L�&�3$'�q߆Q:�`�<�"�Y)t]F
[!N�d�W�<!@���tj()4�ʀ g��ihFL�<�GIo#��[�޵B��1�I�<��K�(:�SÁ�9E�A�<C�I a��E����#̀0-?߰C�� 3�T�@��!z�Yh��VB��C�I�7��	TN_�j����w��&�C�=j�ԸRi�/|F��r&V�e��B�U�X��E�� �9��C�I�#Դ� EE�|�l��C�'zC䉆B�B��f
>s��g V�>�dC䉥wO�y�@V"|ժ`��^2A'C�I*~l�
"/کH�|���)Q;��B�	[Њu�sKN;'J�RhΆ
�ZC�ɾW��*P�@�AZ�$ZA(� 9�8C�I&d2J1r� �f���ȡe�ZC�Irwh�cDAfT����)Z>�B� *��a�i�H���*5�'k�B�I&IE���5�6��x�5j<}ަC�IaS�P;"c=�����iU�FC��.~C4ؓ��E�utLCAɍ�,C�ɶ4�nqS�
^6��@᧙C�@C�	�����3H�LvI�4�b�ZB�5dV�0:�'^�iBn�
v휼+�B��2X1S`O�gr��8�گ)ӆB�)� hM��$��hs�8��闄��);�"O��XW�Y�B�. ���Yƞ��b"O~##�B�:�01�����*�v�`�"O��i���*x.�\��
ئMX���"O6��3Jߛ"D�U�˙m#��e"O�U��cȯW~��ڕ� 5�(��"O`�;*������+}����&"O��c4�,��袗	�^��=�"O�Y!%U�6�&�s�mw[.��"O����㉼!�0ၷ�I$GQ�y�A"OQ��*P��ų�M�{L�a��"O�i�O�.n�e��6=;.t÷"O��;�"�
k�tz�H�	7*|��"O0���ʚ)��q��+ʛA1~DX�"O���#��RA"l�rK� 9��c�"O"��&�L�Tא��S���~�K�"O
�2�팣n&�!� /��#}�A�C"O�%��#Pz���,L�G����"O��80�ޝD�Rr�,EQ%�D"O
����,U�8%����2,y�"O�$	�G���H\���U-(��)"Ox�XRa��7��AG4_���"O�2���}b\ ���C�z�S�"ObI*0�V�~A�u*�+�(J
#Q"OF�(��ڎ�P��l�7|*���T"O��A��}i~�I��C�2+ؘ�"OΡs�o�9
9��A�	�$k��(*O�I�@�/|���oلH����'2��QC��&v��p�3#X;@�&!2�'c��%d��k��R-��0$h8�'�v {e�3�ѻ�j� #�HE�'������̸]
��)�CUz��'>�z�K��D�܉2e��
�`�'���Ld��(�lW�\�s�'��%�KLi��<}��8��'K���&>j?���UnT�n�]�
�'�bT��/��.8�!EbCrx�
�'h^�%�	x������W��
�'��됩�+�>�[Ď�z�����'ɞ���k�=�,����n�^�[�'Ԝkj
Rl�����c�ʼ��'��X2iH
=-V��$�[�*S`I�'��Q�@O���Q�D�'_�dK�'��C슞[��s��W�s�,I��';9s��Q^=�3CRl�@��'7n�te�.c��+��n��DJ�'��4�!M�32�R�cc	�b��'���kr�����,Tǜ��&����&�H�B�d ֮qQu��aj��P�^28L,d`�%S�2�b���q�:��f	�̰��6'Y�E��l����<�炍&]mBM���3a8q��	�M*���xT҅�@��J����A���FF4�̐����I�u�ȓ�2��a��o�1��đW�r���\�8���N��e^���ؔ1EXԆȓIc���cb�D^!�P(�amJ���,.��	�I٭b��q�H؉5�dM��P�B|`Vh��y��=�
R��`�ȓ�iQ��W��15k ue� �ȓ�<I� Z ,���k7��
R�D�ȓt��)� � %{da�";Mj�ńȓ{�~�Ö�FsY0�@O�4���ȓ,��Y�.P!x��%"�3T�ND��S�? B���̌.F�HIDJڈ1�8��"O<���+TJh�5�0��"O���g�ǾV�Z)� f�w߲["OX�hG��m���E�S6;ն��`"O�H�
�$WR���I
��� c"O����ꆃ*V�}q@S#Ј��@"O(;�B&`�|C����rщ	�'�j���gO4r�Zy��b�<DBzY��'T��`�d���k���O�npx�'��$�J��p�@�ő�trj �	�'�����L<����Y�X���Y�'2���Rl�.f:b�Pb
D�;"�(�'��$�'�,FIY2�(ܿe���'��m���؆R2n�pP� c�"��'�`\B��-@�p�B��䢘8�'����W�3n�T�c'������'�T�S� I/s������C���P��'�);��˄,�������N4��'�Ӣ�l����J\���,x�']���c�K#mDR���@K��)�'�(x`,�	,�`�e���z��2
�'�`��2�N�:�F�8��Q�"6B��
�'��h�Eγ�`9���!�|�x
�'.��yw�χ.@���ň��	�'�\)�7���&�
�
�`�>e�	�'�H�xf�P�d��s�T;/�����'�X#ɇ?$� �R#I˔-oh��
�'�����G~	�'�˭W#De�
�'5��U�&͖���4P0��'�����䉀I��Q��JB��(�'��u�*�N�])�W���'%��1w�'Q�,�㠆�V�l���'XV��W�	��q�2�	�f`>��'���Y5$�8�%��L!W�����'7.�;w�Ɇ�*yʱh�� ����'�<�0E�������p욨#>A�
�'kh$*�G����%L�z��:	�'���ņ̀�p�GH�`����'3�|���F�@�YQ�RA8���'��K��N� �����5d� �'���3�dK����Z�CҮW#�1K�'�D�3���`?ڝJ���.Q��|��'	�H�(��(zlkp�;w�~�*�'N���BҚ!`�� 0���|=�'�Je��l�.�9�E��@��p�'
���뀞Tw�L w"͎*c��p�'Ѽe�����G�|=H�IKx	��'�&y:�/�)���g��x�؁�'��M�MA�̩� ��&T8��'<Ԑ�ҁ� ��!2
M�'q��'�TrE7�b-"ď����'z�M�E0v� �����7D��#�'sl�#��1�� B#-����'ǀ4�W���L��^,<��1"�'�ԅ3���$),��`R��>����	�'�� &�M�H���J�a>0���'����I�'JR)R6� ��:�y�DǋTi�)��T76�A��W��y�h �_�z�{���U�ސ�����y���s�0@�ON/0m*1IU?�y%Վf�j�t�D�Ӓx����yR"0�r��a3�V��AǴ�y�2A�*��dN�<} dp��K+�y�f�5-@�(cW�m�� a	��y
� Эr���:*
:#�C��`zU"O&�:r��R�6���H9@ H7"O��T��oӬ��.�u#|݋�"O�a�oR<� �R�>I��"O�U��aU9{[�a�R�G$���"O�Y�%	ƚ`���R%nÌHJl���"OR�%Ɛ�PasG�/P�}`"O�	�ݍ;��$��E֟=��u��"O�#�ɐ�j*e��˙$�Nl��"O�Հ��
|�HČ�_���z�"O�Yȇ�B�Oú�ц�4J��0iR"O���.e�$ث ��5�8�X"O�XJbfT��#�!�9~�0	�"O�$E�>v��SK�.y21˃"Of�J��Mk��rr��hz�A��"O:�zd�7�܁di�fa���"O2�2�!�#�FH��
<oL�9`�"O������o�(Ayd�K92D�9z�"OKϣ?F�3	Y��%q"��yr�D3o>y���\s��£�D��y�T�-��pi2A�$VQDMB�kF��yB�U)�pm2�J	�>(�����y�E K�x@)���9�<��]��y2�Ü�:�{�c��p�!��4�y�ZEC\��B�%���bQ)�y��ï{XE�B*�v��J����y�j.:�༺Pj ~�p[,T�y�j\�C&�Ã�]�P��A��y��r�\�D&~�*���eF�y���D�&��R$�^}p ӭ�y�l�e�� X�X�~���JЁߛ�y2��Z^e1deD�#� Hj'�T��y�NZ�C͞<�QEN�\F�1����yBdڝ��3T+���9#]��y�Ŭ'���`���u2���!��yB@Ȯ-�(:)�u��Hn2�y���m��Ir��]mEB`��C���yR@'��QALP8l��4!&�_��y���&�8��d��wV��e�
?�yN
�[�h]2�Df�0$�@�y2cN��tm-(�&U�6�J�ybm�N��HI�Ź7�Ľ�b�,�y2$Af�<�R���>p&�i����yro@M���'ئ� �0�A��y��Ė ���1��'a*=��<�\��0
�B����MH�OA��]0��q���/J(�BO�ȹ�ȓMhM�رM���b�
��ȓp>X�ʗ�)"8�	���
J�@��S%"�2L�E�蹣W�� W� �� ��dʃT��yD�ܽ�>d��U�fq{�ŀ0 �~���Á0ׂ���]b�T�*V(��c��o$��ȓ60�h́^Dȼ��0k�хȓk_�1��C�5V�Ո͑?H<�ȓpu
�� ��[�tLaW�P�dK���G� h�qD@�`ˆ`�i᪒��y����45��z�*�@�d�Iq���yrAD9��Yb�oI�4� ��bH��yF��h\���V�
	�U����y�B���Y��ɾ9�dQ��,�y��W�� p��:3Z��{3d̶�yreF8%>J�	�Ȁ70�$C�O�y�KR~��e�m҉,k�ًu@�y
� ~� � �x@00�T�V�`щ�"O�ͺ@�Fy� ��Y�<�He"OrEf�3m���%)Vn���"O����ڬhh�1��5W���R"O^A҇i�J�T̀1т/:��2�"O�8�Ï�(FK�[�T𛡎[�yRF��Lq0�%A۠p����-"�y�DS�x�L(�_��UXa#��T��^���`��ʬx��Ѣ2�U:|�^C�I�g:$�H%���;� ��qI\</|B�I�N�tBg&��\���g�4\�C�ɦ���B��~��h��A�F�ZC�Ih�������ywv��S,�pC�I�0�6�"�얰n�2�DBQ�LNJC�	�y�\A2��%9 d���7{>>C�	K'�rF$�P*�W7n�C�$whN81�06������?�C�w&d� B�����)%)�C�13F� Y�";���1�4;bC�I�(�D���hV'TqcV��3�NC�I���c�lİ:HIz�&ˍ�0C�ɍJ5L�a2DC2I�R��aH�cpC�ɤ ���y�Mĳ+�����+YHB�.I#�k�Ǉ�=p���Rl�6(�C�I6Y��u�D#��58��^�%�C�
�&}i��-C�py���&�B�ɹ�̝"����,B�N�+�^C䉚6�PEB�NE(M�Tq�`�[dlB�I0����f儋�X�%��B�����'��%S;�U�cY?
�|B�2|�y��M��e�`�&k:�B�	�iFd��	�T������
�bB�	g@M�v��74&!KU+��T�B�I<h�V�2�$�"F�
Cd��:s�B�	 ���	�m�n�4I��#D�B�ɧO�6��5cٔl��-�S��i�B�ɰ0�|	+S ��$�Z�	�i�83lB�	'�J�O�-[�&]�wC@0q� C�	�h�fY��. c��C���:�B�I�w�X��LU�H���o^$? DC�Iu���L��y�(#sl�mC�IMi4;P�>�
�r�/'!C�Id����N� P[��*���61� C�	�p-�a�D^�ͺPB�z��B䉔{�@! ץ|6V�x��[�H;�B�I�M��P��$9�@�%$i�tB䉴+�@�FA�:HX�e��z�B�I~.>�u��)#?2�+ө��@��B�	"%��ppNF�I�D�36�"|ovB��9���3�
��p��`ŏ��cWjB�I�,�J�8B�R.#�@���>�C�	 f�(Ð�DHz 1��҄Lu�C�7=\.�0%O�4E�j:G*N<3�C�	%h�ꌓe���bDB����m�D"O�B�')K���2���1D� ��c"On�2�JF*}�H�s`ڍ1{R�J�"O�Sb��/��]��O��-n�5��"O�D�r�α2�� ��6�1��"OPe�!Z</��4��Ѳm x��"O�d�Em^�\E�w� X`��"O���Ş=Li8�qǊ�3�0��"O�̩��F�(�4�tI�Q	R"O(,a�>.���Tn����"O كD$йO�h�q3-ɀY����@"O� ���G�U�́�"تK?�pp�"O�U�@A�<:��aX�B�,a�2"O&�DC��K�f�@�۾j�
|�6"OR��&��B��Ba]�4�H�`"Ox)��A���f����]� ��E"O�]�&o[�@K~D����0�
��"O���!��:� � פ��=w^��"Oz��Ќ_�"Y����_��|���"O���Kڰ$���V�c��rt"O2T��� &��iH��ѓN���#q"O�|R��H?/:0�qC Ӭ�B� �"O�P���SSLct�#�h�pq"O�HA%��8w�8$SO�3�謑�"O��
�8�.�2#L�&��r"Oh�│ȔU�	������Y�a"O�ԉb��?�iB��3?�X��w"O�}3sC�^P<
b��b�Hm"O�� �&��`,z�3ĥ� c�z�	""Oz\�D*M�g��1���c��I��"O>;��9?1���F�5a�	q�"Ox̪2K̲C�ћ5��k�P27"O
�"@s*�3��	-RB�PD"O:|���؊ZЪP�����Y<�!C�"O�sr��G�,��ԫ��n.F�s"Ob���jٳX�J��
Y./�^�Yt"O��&�E��}��N-����"Ob�[T�׉pH�@B'5\���"O�HX�B�)fu����>8I���"O��QIإtFJ�YEd	1nH2��S"O��bw�[#C�(��cC.n>�	��"O�����	2\`�2wB�2�!+�"O��*g�ı��B���1{Dh�1"Oh�yF@�(ZgT��V��4,d��b"OR�q`�N�WW��왷n���*�"OѪ�ċS���`�j��	 ��#"O.�`t��>e:��#�H�rK~Z�"O,ai�[�%ќ5c�(��OBP� P"O*��S#�(vQ�1`�F��H�Dd"O�#��.WX|@P'W� n�|�"O����L�N�$)b��רAL�8�W"O���1��8F<P�P��v8�"OPȒ��_5d��Q6�ȗR�j�1�"O���e�(|��E���v	x�"O��1A�֢_~ )s��>↔Z�"Oɪ��/95х!&P:f��q"O�aQ��0�f<�A0"0<��"OT�t�ݖT��M[D��#y@+e"O�H�k�� BJ0to�.^<�2"OP�,]'cM@-�W��><�4X�"O�����HEac�G����"O�p96 
���5�vOA2'ĸ)�4"OtHj�D]�Vts�$��Z��l[�"Oj�(6L�� �t\����	����`"O���Dl_jC^�Q�S ~��"OT��AB�:�2 Y4�
���{G"O�y8�5�lr�L@-*SL�@"O�i���)����g��(d����'"O����M��T
	@B�R	���Pp"O."�|?�T��J��)�H1�"OX���dP����
x��!�"O��X%�ӫe3����	�C�.D��"Oh钔&�(14b����b���5"Oh��_�S����
�S�b��T"O�AX�	:)�%�g� �A�w"O� ��S��שJҾujp�"�҈;�"OB��q�U�!g�yy���;1��8�"Oh�J_�@T�ˠ�D%H2Z��"O�ɀ.J�˂���1
1l��"Ox �E��-�pR� �G}u�`"O|̳�ߍm:<)��$��3�Mڇ"O�1I�`�0j�2H�㒍[T�V"O.���
����s�D�n0v�3"O\�,-����y�VɃ���.J�!�D`)�X��Ϟp�$�e�W%!�J�oϚ��e�@-Ђe� �ƫ/!��|��i���ɓM��P�e�C{&!򄔶k�x)��M�yVX��a]�=!�D��\m�c���"$��X����#!�_�X���Ƚ�,�2!	� !�z/Đ�� ��\�J�˧'I&V�!�$˔k� ��2��?���4G�+~�!�F�$�%C�&�R)���pOS!!�_���׉̅o�bI��G�8�!��Md��a��e�a�"瓭6o!���\�ntad��9lϺ�Dγ^P!�d��~E��l(��b���F7!��7����mH�by�@�J!��NrfF29rDDH��"I.!�D�Zg8��-p�J6��/9!򤀧7�=:������
L1".!�$ʕS#fy�2,�-�:��Ǌ�P!�.0V� &��*����H�1|R!�dª7�`� ��-����b��3!��N&o��m�����e������N�!!�DǴ��0���5VA�V0z!�䑌w8�ɛ�*�e=�xjf��3`!�T'"��m�M�&p5�
1|!�J)��$q�����S��'g!�d�Puƙ�$,I���Lc��]4Lm!�5���S(�?w����s��2@:!�D	�jQ�|��1���+�J�D,!��#u<���A�
I�,�����%!�d߳3�b�(C�Użiȃn��N!�D���R��Jҙ��E��-�X!�D��v!|$����f��H���3�!��J7���x��1#�L9�u�R�aE!�Xg�!��C�6%�H5�K�=!�dZ�nvTr�յ}���(e��"&!��g}B�)5�^���[��)g!�$X6y��y8��}�Q����<*!�M�/ּ��&W�� %��
	3p!��JM��r�I�38�AZ��Z�PyB$_J4H�(�2E�Cb��y��Cԁ��Ί!r�� %�?�y��[)V���)��)r�`(G�#�y�c��5�}��'T�	 ������y�K_�BA�C���T���ܠ�yb��!*�$�%�]G~�&ȓ�y"�Y*J���!�r2T���W�y�"�0X4tR�F=P��A5%��yR"D�gI|:��N+<X#"��y��C���h�b�DDp0i2B�/�yB"E�*,�AkvGQ 6GT��D�U��y"��V�V�2 o��%tNt��cU��y�j�3N�~x`1$J��|X�6�4�y$__�̭;g�P/&Y�e�V��y"�O�q��:�`_	M��je��yr�B�SH�g�B#{�	�1G��y
� ҄��B�QH�Is A�<
`)!"O�(#chM�j
��R0�]�4"O�uZ�Nǂ]���Ǒ�ĭ@!"O���!�G�=��f"5�l&�'D�$A�%M�|Z#A�0G���3�8D��օ�rvh��A8�=5
7D��b䭀���6�S�Q���!5D��*B�R2v�v�[p	ӸYRݫ�1D�<`⃚�#���G�ҞR�v�+#D���`���/����T'�Z]~����?D����7��0X���[@ ySd8D����<r��|�L0B�vf7D��q��:5�����ޘ%� Jqa1D����g��\�4PG�9S��$�Q�0D�ʦ1E�xp��`ٯd�D�A�:D�����%?�Bp���Տfk�˱�2D����������F=��J��=D�hk��Z:�%u���0��e+)D�d��FU=�������zU#I%D����ʓ0�F@H���|b�"D��*���.�(9�KȌ*���!D��&(�O�VQy�E0�����=D��@4
�
a�}jÍ�p,�5�(D�0;B�UD
�arF�d
<P�W�'D�<jD	@�R�n�S� �	�Tt�!�$D�2�,\�x���(�/ϩ	�n\��+$D�����E��1�$��<�6��#"D�01B�#3Aj$�^
T��qpC�=D��f�(=`�"�Ѹ6е���;D�heG�TNz9����<OΉ��'D��� �Wɒw��4G[(�y�N��^!��ZE�� !Q��ǵ&�!�$�0���ba^J�Vx� l�y�!�ڀ#�	���s���Ka+��_z!��_��~ȁ�J����Y��B�^�!�ۣS,�e!7�
�M�.]�aN��!�d��f�PnS#e�>��q���?w!�ҡ�^%���X0;�Z�au!�$q�L�˓
�]&�a[�Y�!�
���U�Cؚ��F�!��&k�,�"���\UP��S,�!�E;%����ǂ+6���� Q�-�!�d�6X�0�p7a>��W�!�R�G�eZG£q����b(޾c�!�θWWP�bU�( �,�0�\�!���<N���b�E,3���څ���!�d	����B](�c�я]:!�$�<��}�Pd�PgN�8��l�!�DH�V�uo�:[Hu��1�!���IR�j���N��'b�)�!�}t$�)��8�A�&L�!�ќ2�D�ҪѰz��Qk�&֌�!�D�3$b���#�Ĕ'�����+I�?!�Ši2<Xoͨg�5y�o �Vr!��b���qK����Za��4�!�$G+���c��"|w�h��K�%�!��T�Aj�L�#�Z���	Ԣ[�!��Ċ<�zHc#�ɒ8Y�pc��Z=:�!��>7�p�UP�MC>�;p��m�!�P	g0ؔM�8@�-�/ �.E�� �2Q0�"5Z��lh$k��qh����8�<��c�#^�^��q���Z�l��`�>�j�➐lc��Zcm^�sl�9�ȓ�����.H��� ��o�z��S�? ���j�X�4[��i�tay�"OpI�1�I�,]�%�B��5+ ꠐ�"Oʕ�C�?4�J�rs@_���0i�"OΡ	���x\@9���7�!:�"OX�Ӊޞ1'zx����Y�a:"O888+ٸJ��+Ў���"l�"Ot@����f��Nњ6��P"O�ܲp#�4#R^L+ƛP���"O"9����i.���cMd�h���"OZY07S�OuN\�&��	���aF"Odx9�ɩC�t�qR���\�X�3�"O�]������Ce	U�v�$q�"O�͓�)��/����S�`��KG"O 1����ma��b#'�9�"O��Z�m�2�8M��@�"�1`G"O�E�1��?t�$��,-=���"O�u�%�C�Х�̍X�%�c"Oƙ+�'g�x́I���˳"On�8�h@�~�ܭ
�a������"Ov=���<
������Y�20Ӑ"Of4𖯚�6ٮ���_���e�g"Od�@#�?��!�f�u����"Ox��o�o����fN�Y>̩��"O�a�6��&�.�a�儢�R���"O�Ye�ȵ`gz� �D	%VÀU��"OBTP���/S���FN%{J����"O�8��]�W��@�$�5L�(b"O��0��öV�X0��X�~u(�"Ov H&hP��Y��J6	��"Ol��š���캓.�*f@�Zf"O�hZWC��晣���&T��i�"OLt�/��|��-�k�,e6���f"O*���L	�/e���)��l�h!��"O�=�f�\�����P2JVRL�"O^��F��+4�B�'V�k��9��"ON�3��n���We�. w�pt"O~� ���aǐ���$A�}t�$r�"Ol�C"�478������0f"���"O&-�5�_�D5���KK��#"OH�{�P��Ɂ��v4ƵQ#"O,�p�ʁd�8�0�ޯ`��cc"O�|i$�8�l���U� �HR"O>���'o0�D2���7v�!�c"O 4k�
b�.���L�xqpeI�"O�P�%iŔ4�V�R*�F�@D�@"O���5�=�u)B�b}J��6"O�9���-e����*ʤ:`
	`�"OP�#�Q;$U|��c^,H����"O*Xh�m�:�;֌�0$ ��"O %��B�"�(�l��Vl5��"O�TZd@	�(d ��3JE�
Eh��"O>1i�o�=�$��HLHS��"O�0b�Ejq�|c��OL�=�"O�d�u,̤"ߦ@[t!D�<z���"O�8�B#�$��,P��Fզ5�@"O.!2�)��(t�� b�,��f"Oj|��E�\/T`ʑHW�m��u��"O���E ��z��ţ���#Y(Np@"O���`@�e���'�6S%V���"O��� 00:�"�%L*tAr(�"O&��ǰ�V� e�> ݰ�:4"O&1�����jw�<V�9�0h�"Oj�·D��B*��x VQ�(��`!�D� h�Ƚx��9\������G!�� =�Fǟ�d��!3퐶r]��	5"O䅱�^��@4"W��&~=����"O~�z��n[����hA>����A"O8+1oː|��!��g�7.�E�t"O4��D�z��p��G='��:�"O84�dÕ)%�4�k��4g��}�"O�<�ŀ��H�Q Y/t�J�3"O�x ���%�>}Y��
�uGB�V"OF�iI--E��@�,�<.����"O$�x�����ӕlR�OP��v"OLa��A-��p���  �~�{�"O8�U$�d��1�ꔖN�8`�f"O��r�)v\!;`����H�"O$����=�F|�Տ�5�9��"OL����ޢ �FY0!m��4��;"OD��$����:N�����"Oĕ�3�F�\OxA3�퓛k ��G"OD��1�(
�n X�̍�]��3�"O����>	� ��*�r46y�C"Oڹ�(�J��� �N=L,8��"O��3s� 0,���ES	3	��Z�"OD!qb��1DR]�W�̂��Y��"O��H����ƌC��W�بѤ"O<����'D��3�%
 6x2"O��PI'@���ã@�,(��"c"O0ˠ�"(�����_����"O�yy4��_�
@�2і�Av"O̽)H��e���@�V�"v"OXa&�%C��� ����d"�"Ou���[�>�*�ȶMD�Zlh`"S"O��HQE.z�Q�&m�zو�"O�P�� ���@��J�<��P��"O"�K�+#�����)��0�#V"O,���٣�ޘ����g��	X"Ox�Ad�;�zU@R�J�l̄��e"O��G�5OZ����/e��DXf"O,�BCD���b��H�,�(�"O(a��*��l$hBgRc�<��#"O\�'FC�cWĀ�0f1�T1S1"O"\ء�_B���0�_�<�c!"O69x�$H�i�� 1kȇLnr�"O ��M�0h�n�˒�խuj,�B�"O��U�O�(0a��'A\��u"O�,�Q�۵c)��B�? 1�"O�@�1�)wd�q�Az+pqK�"O���b�ƑP0f��p��3p�-A�"Or	��G�`������vUX��T"OX��#���f�h�I3L�9T Ԓ�"O������u�2�I'
��/@�s7"O>�����}^T�/� ����"O��顄�,=<3��E>J�xP�"O�X�AF̼+ bp��LRll�1z "O��³.��C4�M����\0�0˖"O�xc�d9���`A�_"�4��"OZ-Kcˇ��}��o��v�$�"�"O8 �v�U%�.�#�g��
���a�"Ojl����� �EsKܦ�R"Ot���
��:ָ����k��A1E"O$Y{���0�Ҵ��&��#�2��A"O�x	��	,�t!�! @&_��I3w"O�:ղ�q�T�^�NQ�(��!��p�`I�K*e�È�4!�D�`��=�I�$&�b��T�m�!�D�{��q!�(Y��!��@��!�� ��QT�Y�d�\A�Bj-iR��R�"O���%� ;:3���:Y"�9��"OaC�Y��
e� �^�{j�jR"O�Y�/�4��T���$Z5T�:�"O��$�$I�qh&.��f�U�T"O�
��Ŕ(��y�O�#,ty�"O<Y2I�C�`y+&�ݕ^?^!p&"O������|�p�I����^$�L��"O �!D��9O�Q�t�NAV�B�"O�D�M�#y�]D#H�"'d�"O�p�fm��1������8"`	��"O�yG�=w5���1F�,M6�!"O������@c2w��9*��%"O����Ï;A�j��ȼGbf��R"O�-�Iݧ3@ԕx�
^�;z�q�"O�������Nn,Zլ�;xGH���"O�<�pmJ1LXX`b��.*�]�2"O`i@���p��5Jp�X���"O�|'*Q_?p�ˁoA��[�"O��)JEP>�X����@��1"O�Z���)V��r°!9�s"O����¨�,Z��̗1�� "OvP�Ad� |�� �g����r"OJt�q/
0r-w�1y]�� 3"O]{$�M��Xtc'M�!YipeP�"O�<�ę�L��BK��),L� "O��Bm��t�����?X���ycT*r��5IR�ЇJ�d�0�	�yR)Pr�-�堑�5�x�sׂ�yrBL)׈��g�����mݩ�y�A<J���ŧ�!�`	X�ߍ�yr(N�s�i�q���5f@�dŒ:�y�`� �b�Iǭ 0\�seA�1�y��@=8�4y���l;�u�d���yh	�m��'�(:f��RÉ	��y!�y����+WX,Ks!��y�.2q�8T�킸x�����E��yb��!����S�`$t�Z#F��y���vs�h��j�
aBX�Z�g��yrǞ�M"\��c�Ľ_W�}k"+��yb�܍*r��ը +3�3����y�aQ�I�[��G�/���f��y2�!PHNjg�].�o˸�y��9*Vas �ͩN��usPD�y��J�N�#�	.T�J슧�ü�y"H�} �%����$GB�A�ņ���y�*�;�Ƒ:�C
5V$dI����y�/ �p�f&#�"i�t�ɥ�y�(˫Gn4�[C靧�4�+�/�y��X(FN����9?���Q%�y2�F�2���P $\�@Q0�����yrf˫N�X@�*�<~A��@��y�\�_x���X,F�8K�m�"�yR*J����@"(�@YC��_��yBe�j!ɇ	ÛK(*�q�G���y�'E�-hT���o�L4� R5�R��y2D�Fl�P�ު�`5A��E��y���
n��%��b����4���y2�T�G���ǉYl���S� �ybF�,��K�藖V%��S�Q�y��
_:�p�Ć ���9�& V�y�GȦz�Y�v��r|M;�kO��yª���Z��8`J�4&���y�悉i�F<����;5����e��y
� >d���Ȝj�HEG��q��c"OZ�IEfV*}�^�BF���u�P�"O� ��0j�.��e��u�"O���̘��j��5��/
�"O$��1��&k����ODS�H�R"O��[�ˎx``)<|�"O"���Rk6r	3 � �|�3%"OjT�`&L\�<����0��aG"O-���ܵ��]Ѷ�A�s�`T�"O�L�oެRl��s�R�Q�$��c"O�� �!^ ����'ОnTѺ�"O�d;� �S�h GΙ:_��y�"O.� f��t̬e贃���y1�"O|�w��,),\z!�J# ��$"O
�q׉�R�����J�BИ�"O�hæފm�8�qH�f���S"OR| Q=(v��Xc�	ڣ"OȔ1��C�@��͚�){��T�"O�ѐ�͞�\���6)_%[�̻#"O�$�%�D����-ݏa��=p�"O�=)g�O)i>,Њ�K^]ot�Q"O�	���R#:�<�����2J6�b"O���PÑ>�9��R�(<���"O������**��$;��?<1@a��"O��t� �K��@	�2*@��!"O�c�eS�$�~��?U,@�S�"OrzW��blt=af�Cm(@�96"O�ł�������<( uP�"Oބ
qS�|�	��O�}kV��q"OԨ+��.?&���BKV�X��"O�TEAܫ8��l1)�"\p���"O��xeB� ��
�2R���"O��9&�њx*�pgjZ
qpN��"O��#��?s耤kwI�"a���a�"OĄ�uAE��t�a�Ŋ�O���W"O�}�K��(4�%F(�"O���dca]���T�
�*�r�"Ol���$�2pze;���L,B��`"O ���]a��SU��2�(��'v�|CƏܑZ��Y�q�rJ��L�<AG�¥s�L+яN	���3�H�<q��Ű(��4��F�����z�τD�<�4d�%��<�a�	(�X"��J�<)�dQ
 f#�I�*D�"���LAE�<�-ͻW�敲S�W*@gr}*HA�<�R��<?jl�:�&��b��j�\|�<a"`� z�"��'�»q3�R��E|�<�3���������E�Nx��M�<�n�7`P5ඡi��}��ȗM�<A��5y*1z��L>K��C��\F�<Y�G�yq�cDM8�08��K�<i��p�X�q���*kyJ�x��Q�<���
����@�JqS�m`w+�P�<a2�O).6f�B4`�;D�(0p@�K�<���ٮ&��u��(�5B�H�<i�
;Y0�(��ǟ�V
v�hVLDl�<�b�� A����q'���s"Hh�<�!L��RC>|�-+֦ԢS��g�<a���(=��
�bG���	��e�L�<�!����јF_������)D��T�R�V�ne��%�0�.�i�J;D��*��ѩ-,��e��{T8����9D��"�!�ݻw�¬+�H5Pdl7D�8����z�!��TgLt���6D�� �$v�ިQrzP �i��'Bp�P1"O&8ۇI@�~9��b�_���"OFE�3D9 �����_� �=(g"O�������ܰ��\M�\��"O�0Q�&#Q>͘e�A�t���s"O��Pk�6�D��Y�y�&"O����gW��L��m.N�@��"O�$�Iu�D-�G�S�4����"O��׌ǐO���z�d�(z�Ȁ8U"O|�yw��0�jvBۣ;&F�"O�$���;c!���f�J�r"ؙ�"O,�;��	�B�����!*."��V"O�UA�%�!J7 ��b�ۚEa"O ��׍EW��I��	�;���D"O$%I�(�	�V0��T�~���w"O�8�e���$8(d�E�SD"�q�"ON�8��R̒��]�Zv�a�A�W��y2던9{�xPC�C|h1	
��y��	'L�B�b�DY�>s��s �Y��y���h}�d�Z�7���Ԡ��y���B}4L)4�=/��� ���	�y�I�� �0	��l��:��g���y�U��Q��*���ï\!�y��-~:�؅�FS�e �&͠�y�#bz4��bJ�GS|��a'�yB)!b!�T�^8J�}�G+A��y2/��V��tD�4>p0��bۅ�y�A�-	&@Q�#;4<b�VY�y���hfր�1$��Z�r�Ke	�3�y�jحZ�64:��NK��Xb$�$�y�A)sR�)��D (J�9�q%I-�y�o���a�g��jt��Yf"Ы�y�y���(�@������:�yeO�`Z�
�hֶ�25H�����y"��A��E�1�2-�%Q'
[��y"狪~�Ν'L߶0X�Pgث�y"�*�r)KOǒ#���[�)<�yRo�8^K�{E-Ϡ�����@��y���K5"�B��Y �QSL_��yr�Z�%��!I`I�8���BD���yB�P�TґB�O� :Rܲb��y"Z�g�\� �� �8��&�y���
 ���Y�Ȋ
A�x@`/̙�yB
���ś��ܧ�J �6�́�y��W�A�& /�=P�Q�����y�-��yn�5��a�<���Be@��y��Z
�����o+w�>��"��y�Ɋ�B�\�Kǂ�k�*�fo]��y���^*��t��,]��8�[��y"��#Z�����@�fè���]��yr'�<�f�Q��ܙ��G&1�y���&/��z��	(#��f
��y�"��G�0)wL��o��a�N��yBH�)lM�FB�x�"�Qa@���ybF����1�b܉td�����yr�Q9|DM���Z�r2��3Ce��yb�ّD6~��!SeX�=r��M��yR��q�,`T��2O�6��`_	�yr(���azEh uf�h�-��y2�L&g��!�g9i-����#�y"��f0��4 ۹[�&�/��yB�~�2�F�$�Ĩ�'����yr(�Q�`��Aj@�S�X�'K�2�y�֣'��K�k��9(�J�y
� *4w.5{L��&o���ɫ�"O�5��#ۭtv�����Q(հ��"OT���#M�Q,�T/]3�����"O�ˇo�)h2�#���J�J���"O�����2n��a�M�w:l�a�"O(����;�m��F�
&�1��"O�+)BH��BIנeg��b�"Ol���߇6�^0�2Cԫct��*�"O2A P��K�nQ���ޒPYpE�"O�E� KE�>N��ɣË!m�p�q"O:�QrF1}�4�� ĩJ�JHJu"Oyx�ǟz��id��$�y�F"Ol�a�� %Rܒ��E蒰6���8"O.�QtE1�٣��E�
t�`"O\#paB�yȼ����%��%�"O,�Z&�?��c�W���"O&�c�ņ��`@�LZ�f���"O���B�,u��8�� ��=��"O.��F�w�P� � �C�h�+�"O��@QHҧHr�AT 1��r�"O����
������O�{6���"O�EGB  wx�-\&|y�"OV� ǅŁW�v����{�TI��"O���g��-��5���]�"�`�"O$�"� �0���8�"oj}p"O��r���
@�5� �!0X�Dq�"O����)�D��+��Y�0�$"Oڐ��#�$��!�
" ݄+�"O�!�tI��J�ʡ�u@���z��"O"eٷ �aa��2�`ٓ�%b��y"�'�h J��݂���d�_��yr�1\|�U�ݡ{�x��K�yR"��Sߘa�v�z�b�(�>�xb�'��c�j]=O��x�"'�zP�'>���'P��zu�J��(��
�'j�����P�Y8�5��	ͬF]��
�'����˕]����7#v�&A�	�'#�q��-������F�R7q�h@�'�^{5��q���3�J>w�V9��'Z���F�2E�|���I�$uu �(�'Q���ԁV�E��YƌZ�Ü<@�'ORl�vAr���@� l����wn6D�p��+I���-Y�咳H���b�&D���	�$I� �s��&% ,�XPŅX�'����9O�4���,����*5Rk�<�'"O<�i����N���f�*q���t:O����ԝdx�K����d,#&���{r�$�)Yj�IsΒ:Q��Z��\#�
O^؛F�g*�QQ��+_�5���'�'pV��rP38>\��<�YC	!D��1aea�@�vW���G�$��C��)P�����ނdS�q���ޚh��C�	�L>fY+S�١A��Eh� �L��B䉀'���Ћ�7O� � TG1*G�B�I%/� <jW�2$=ƀ:Vo�6"�Z�	K��܉�o�,�F�X���5<l��W�"�O�O>!�o��a1Xd� �D�e�V���"O�ȣ��A79ȨE,�"]�&%���H��䓼?���Sm?�f_�QdL�C O@��ly�<�rGĒ��5t�\�?Ȑ�Ey�<��-W�=�B��Q���?�vu0�$�P�<bDJ�*eHP��D��̅��/v�<�bt�xe�"'RL\��k�<���6$�|��̝GH+w�d�<� �RG��v� EM�J�X��7"O��Pg(#'N�B�
fJ�L �"O����8~y�e%ɞ['L��0�� D{��)!{�����[�������r�xB�I)& ��g(�#TJMXT�[7f��C� ��[�)��r\ᡶ%Yg��B�I������O�0�т�n�v�Z�1Є(D�DB�i  O��K��`BX�!M(D�L�T)ݺNF�H +��=u$����2$��J'�&Gz���
zM@���y2��e@d1 Kx}z܋�����y���D�h( ���(�4]����y��N��"&��:^��h���'�ў����]�}��Ԡ��B�jR��"O�I3m�"Ev"d@�/$:^��X��d�<��4��1 �τ"sM���a�QPb}HG"Oz�	dgV*�䩗�_ 8c����>َ����*m����N�jg�aj���a�!�!,P��S��\�yb�]R���a�!��H�B=+�`����њB�a~�P���"nE� ��ɛ�,_�h��{�-#D�T�sgW5g�$��ҫj����d�LD{��	K�� ۥ	G.w���;���!�d-%0��GY
)��lC�d	���ɟ�HO�>y��L�5Z�>Q�/<JpȷJ><O�#<y\��P�k��A���ī^�-�PM'��#�l���+� �%0���O���q���h�INyR�B�KY� x� H�h0TD����w�<Q�#A�G� �sP�>8%"��*u�Iϟ��?��{�/B/7������7^7���L���y��Z���=�q��)f�R�s�Q��3�S�O��4R�m�,-�l$��^+&$�S� i�đ�X�2�"b�&<��aBCէ~�!�$L�O&F�3&T���bÐ	]�џF�.�8}�����MC�pC�Ў�>�yi��{Z �[�b��,�%�B�	�	|8�
WGWC~H1���B�	�fC�eh&�R A�jHQA惘-�B�I�yfj�����d��	H�-A�5�C�T@\;�M�(1������C�	w�"�q���w��eQ�ü#,FC��-�&,�r����;�Èr@C�Iv	(i�#��0ZA�A�o��N�C�I�0lZ '��*@�t�z�g�9O��C���(jd��E�@�y��1��C�	�?j�����F=�jE��M�}�B��.~iH\Ƌ��J����&�  DTC�(:N1�'.��5c�`u��)Z�8C��495����^ǀ� J�5$6C�ɾC��D��J�,�l9�s&ި'*�C�:)��Z�-�@q`�
5`>��B䉼|�:!�A�CR=S��٫U��B�	 5<(���a%�JA�R"F��B� >��j����J����!!)ߚB�9/R���#�k��Tɂ
6�hB�ɔg�y�#�	�O��٣$��fDB�(!6d����^�=x� ݿP�FC�I?|�!��d�!�X�g&�j��C�ɍ/|)SB��B���A2u�fB�Z��CN�%�� ��9��<�ȓS��(�A�i�)ϐ�y�D�ȓ �L�U@�$�8#��C�7����)��t�����A`T�@D��X���`S��;)F���4��*!����S�? p�x�i��|�:p(K�-��г�"O�j+��?~�a�! �3(�V�H"O�Ĩ�hѩi���,���8p"O�=YQnٚ*W��B�z�f��"OH}R郘[I�q�@�+F"^I�"O��Ah�-n^���aϞv�}p�"O΁:M�p����$OP�B��r�"O�I��	m�D$j�.�:D���"O��%�+�"���X�A b�"O�8cK��c�f������1in0z�"O�q�T�Ӄ,\f,۷�0\Y�uPT"O�TD!F������_�!��b'"O������u���lʘ>Hi�"O E��߰l�|1���{�:�8#"O��"kI:r���FKѥp�aR�"Oh Ç	"j�mp&K�O�䁴"Oh��P��v1�Siߺ~����"O�8�G9f4��AH�b0��"O�(��l
@\F��0c]�f(�x�w"O1��N73���8#��ʖ"O���'E��_�(�j6b�-xTZ�"Op}��	"�q�#+C�l{b"O���MA�hM\0X�H����s"Oq1��K)�M2�C��o��q�B)D���0$�'�Te�� M����c�;D�,��h\M��+�iO$Ş� Q�;D�ةr��z� 0���T�l� �&D���CÐ[�C�G��py��8��7D�d[&��;Y�V���<fz���O5D�,��υ&>�y��@_�]�h��3F2D�d�ecM�*�H��#C�C,�dCO.D���`[�D�I����TV���,D�,0�	|`�����1F�v��)D�TJ�θ��i+a�^�	j*�"PO&D�� �B%�(����?w�:�s� &D��2�νs�L�	�G�M^�ɉ�>D�@Bd�Gi���顯T�y�5��:D�P+F��E3�[�ҫ;���:� 8D�\���߻sx�s���6��x	��*D������2vG �ƘA,
����5D��*6��Ar4P"�����!��?D��r#T�3��W�lR�����>D��C��< x1�׮��u	� =D���`mĤQ��m�4�C��[�N?D�p��ܩFǎ���e�A�5���;D�;R��$ �Z��C��U���5D�Tc�N
]o�q37&�,v�^���K4D��C�x�F�(�m�>�L���3D�l�3�{�h�k�I��g\<�!�0D��v�� m"a�>j�,x��2D�����L�nH�����ti\� f1D�� ��c��(w�ĩtX8�`C0D� XA��C�:��G&�TL��G D��r��բD��`	�C�d�8t'+D���`��~n2$	c���9N՚#�(D��)�I�TB(�qc������*D� 	���Nce��j�����(D���#� cj�h��l�G�Qá�3D�z0�-\m:l��ח6*�h�r.&D���VLI������yY�%��#D�9Я��`�t������`!��*5D��RU� ��~]k'��)r�*9;G�3D�k��8B�w�0� ���TC䉱͈\�"�Wy��i�U)�* ^B�)� ��r䕩h���q)}��L��"O��t�Y��j�`�%�R���"O��KCb��f����րT�йj�"On��q�ܤg&9y@�^&��	�@"Oj�CW�M9n~�: R�=���H�"O��C"K�g"ECq�M`D��"O�C%'	@9 ��e0^L� �"O.�I!OG$K ���ɂ}�f�Ѧ"O6���gG8sid9xsCժ@: ��"Ot���mX���A�-a�Pj�"O���ꂡ.f��!�O�	O:@J"O���Gk��l|i��̉b?vuI"OjH �#�6w�dH��o"*�X�Qt"O�]��f���@Y"�C K�f�{�"O� ����y7^]
`��9�^P�"OP����(L4�1@��R�U��I%"O1"原�*w�mңm_�"��PB"O�(`6 ӽ&Td�S-ܣ!�,���"O�y)`��O�`��+ja�#ԛ�yr.��E��ӥQ�P��{��ٹ�y��WX�U;I�H��F�F�yb�;(��{�ҫ?�y6����y��X�m�X���@!h%�1�uN���y�ҡJ����3�4�ܭ�R�P��y����Z�pɪ�OX ̸�:BHͭ�y�Z��ӑ���pH*��p.�'�yr�N;y@b���:rh�0ӨӦ�y򬂽b��ph�䇂xv����醘�y����ZR'M jsH}�����y�@J=Dez��EZ:rUIs��yIU*3�pɒ�d̔\`v�#F�y���2[ľ �g�.T<*�֟�y�D\isM�,M��`���y���C&�j���4t�^������ya��B��q�n���!p��9�y����s Y�aSH�����y�j�dj���	iP��(���yR�H 21��$�	]G
I�����y$Z�5�Mʁ�$�,Mk�ƞS�<��_��>�)���t�8�QQ`�@�<�a%�T�d�1sL�b��Jf�}�<٠��^��2�	D�ڨ%CF)�]�<Q+�	�Bј���?<*�!�׀N[�<�6��Zr>E���4f��R`_Z�<�Ђ�'v�F�"��6>�T��Y�<���_�9�L�c��б�R��Y�D{ĺ�С�`E�2��PKŋ��yr\�]T�i�1ĝ 1"��5b֋�y�A[?c�\���Ȅ9����FJ�y"�ʷh7@	*aNU�������ן�yR,nvXPC�'s����ŕ�0>iO>�Ƿo�غ@/� BV��)$�B�<�
��W���`��Hbr�!��B>� �ȓS"�)�� g���R$U�6��ȓK�X�W��Y�
�TkǍTy�Ą�nͨv�$K���R�]����l-8s`<v�ԫ�D@+P����ȓ*���<����@��	����K��ix�FL�Oa�����(JS�ȓkʬ@@G�&Y���˝+�؇ȓ�M��ߑ_s��Y�HՑ=
���'��a�O�R���'�.�@	�'����"�wa�5�P���u:�� 	�'%�z$.��.�@DK�Mh$M��yr��� ��P	�Zh޹C��\*���B"OV%�tmN�#t��TE�=IyBU��"OJ�@��5����F�D�7Z���"O�iD!����pQkE%�|�kv"O�i�T��5sH�s�	�F�$��Q"O��r�Fbk�2�x�'�:S�P�
O�7���"�̱ȡ�K�,N��Mϧ K��hO��M�3B
�@r�yA焛�v-��"Oj�S�����AdA�zw
��"Ou�QgV�{dv��t��	D�̰�W"O�ib�c.hр*���d"OV=��(#���R��?-a���"O�=p`n�r�X2,�Yjy�'O0=�c�� �L��RE�E���8$%�J�	�Q�"|��'\"g�vE9wE��3|���`�{���<� (^�S/Z�i�큂7&8�h �y�<�t�--��d��JQބ�Q��u����d���E��¼\KP��b`�#X����Bݝt�!��hX\�����$�֨;#+�f����F{��� ��΀:P& *�/Y�8N��g"O.�����$���e��/L���B"OPH�� �q��Qr�+	�m�#"O�i���H�('EC+i���V"O��J��'��9���Ǐ�2�d"O"2�D)O���"@%� �b-Q�"O\�s��W�Ne#���(��	�"O$A���]�Y�d�%=m>�"O��v�@,#����)Y�f��4"O�M;�$�M}�i�bE* .R�x�"O��3��|�B�7��9m�!�"O�A5$�%j�Xc��t��d�V"Oz���P
 �e��߳}8`�3"O�1-_�)z��EF�4����F"O>�����>���@`�W>宵�""O$�E4I}�Э}�B�"O�H�K��M#���g�!G�0,;s"O������#�B�J�ƕ��`) "O��"cV�d�xZd���FNDD�"O>��Di�_X���U�*D:�"O&���G�4>���i�>T"O���EN		K09a�Ǟ?1�p!��"OZh��M
4i�>�;BH���F��"O�x�@F(DNa��m�D��B"OHd� �϶ �.i�g�Z`+D"O|�6�+)5@�3���]zn���"O����*�{�:4�W �] �R"O��)#B�Q�M��Ȓ�($�8A"O�:g�,R���ևCi�P9�"OV�+�k��2�q��.Ҡ��"O(af�Ƃi��Pa���Jr8�f"OT[���M��!j-�Ld�T1�"O^(��!��Iފ`�v-	-l���#"O���P�C=c��M�ąAiʆ���"O�@+�$��5j�%M0��5�>�y��єG��5CFA�?��U��F���y҇�8 ������4�qč
��y��6pT��	�(�{��E���yB,�[���YvG�4p��-P���y�B#P��L[�A�1k�vE�-��y���G��Q���0j��@8����y���P!0X��B�LcBT!fO<�yR��6@�M�h�1A�8I�u
��yb�ǰ]�4�#K��@��!�T爎�yB*�$Nrp	Ue�'�Ar$�M&�y
� ���L��to\e�v@��`Ԅk�"O�)��&��DnË3Z�}��"O���C�0G���#��\��"OI��*��u~��A	�li�L�S"Oҕ���@b�lc��\3Fj�*�"O�۵��#k�YB�-�k"-ؓ"O}���^�vZ����O�fV6��"O$y���V���d띊 7��#!"ONM���ʶ�ީ[S*�<J)�ј "O��b�IM�,��A��7/�<U*T"O pj��Z�98i�R���<�%��"O��(���1���C��@6��X"O������.MraɄ�J0u�"OnɁV 
!fe�*W�ڞ+9���"Of�ѐ�'(�Y�*�LQ����"OR���|er���ݧB�q2�"Of��r&K;\E�-z�*�G�hH(�"O����V�,�@[a�2o2|�"Op�s�D�&T�~�R��Zɔ}Z2"O�L���%����+��!�"O,�I5%Ngzm�B�5��t"O�L��Es��,3Մنl�-�d"O�\�ebP�vE�i�P��Y����"O�\aD,/-󠈊�c��;S����"O̹��/���Qg�ɧ6��I"O��XR��?^@ ƍI�E��xv"O�y��/G$� ��P�E8ST��6"O40�%#S�M0ܒSm80rj衢"Op1�%��_y�0�!���"��Q'"O�ĳq��iz�Ŗ��p��"O�L3e�g�X����K�S���0"Ob��B��Uv�iA��L�$�A�"O�4��L'��H7Б$���"O��@BbK�)������1"O�T5���t��%����2	��!�%"OV�Ss!6.�K G1P���"O�p�SH	/;��6 RJp	z�"O�� $�JC���i�oX�@��x#"O2��$ʞ97
 ���(H|�A"O�ykW�^�l��K `[6���y"O"��d�L���K�$2�����"O��S�X�lp���dV (�V"O*x#��	?R����EA�
"Od�7�,2�� �.�<*��"O4�!���T��K�|S�)Q�"O���Gl*������Sז���"O�!R��Pǖ�uK�31[<�Z"OT��Q�E�|��Ll�tQ#"O����C���m�P�5jQ���0"O�%��k�PI�'E��"�
]J�"O���Ĉ\(_�U�DÌ�fz��b"O�L�֯\ \�d$�փ�)>;�I�"O�9UMv����w�B�
&���"O��1��<b�V�ضHR<(
*�#�"O�����(9M�1 G-�0ܪ|�""OК�X4K�u��,�8W�^��%"O�%1#[l �� Cˏ#,�1"O��v�E!0�
�o%Z��&"Oȉ
fgȟϪ��4�S�be��"O��p7̎,\�|�`��y��)"O�y:�
�@���*��2upW"O���0bQ� ��W�X�6�i�a"O8���S�D'N�C��(�t�)�"O������0��{r!�;8�Hiy@"O� �a�Q�U�Ԇ "C�C�b®Pc�"O4�bN�3�z��t�� �6�Q�"O^y��B:H�Zu�k�2**��A"O��	���'�v�;B)ͨ}�)���'�b����9$�̰��O�5՘��E�a(���0�ܰ��X^M�!�ȓ;�(����Ҁtuθ[��QhZA�ȓ� �e�בB����4*E�ެ�ȓ�Ƭ�P!ӋY�T�[�y%Z���'*�Dʑ)��ADbA�S,~�8ez�'v\)�]��C��L�����{�<��@����Ӓ���p�<i��P����Fn?>��t�*HI�<��D�{쬄�0�G?D9�R^> B�	%�<�%�|}�]B��"�8C�)+�3t�4����WD�	_�C�($��h�(��^�Q���B�ɝpC��Ȑ5�Q5	�;3��C�ɰB��HA�̃w鲱�#�,{��C�, '8U��h566ni���_OxC䉕o���+(�:!њ���O��b��C�	�11�Ј5H��s��"��}�C�ɮ��I��^���Q�Ro*�C��38r�mY�Ch)����-6$�C�	�FF8��J	m8A	��ΈZZJB��`7� 1�&��zZT���k�+��B�I�9�񃃆,7^D�V��r�B�I8Yz�y�K>A.�uQ�d��xs�B�ɫg�F��i�)���b�	��B�ɽxU�@�$nا'��kW�D�O�>B�	 Gve@UL�#b �(T5��C�	�K>�lKB'
"�"�AV���O�B�	�
� ��a�U*	�� �@�<C�I�w�4Z�郌��X��I�RB�IRr��F-�7 ^�h׃�kp�B�7_�$��ʒr��8;�薈e�lB��$a@��'f>x��B! .6T"=��1 �bT�S���Ow����L�wz��@6x?�L[	�'0���6iC
:��2R��'j0�����l�0�����"Lu�󧈟��Q�:-��q�@݇Z%xQ�欌�5!�Ğ #�QP�Rz� �r�,���"��d�,e��O3-�]��ϨO�p��db~�YF�T>aΌ���'���L��!T�!�@���n�*#B�M�elD�1P��?��~�d!)��y��&�t��ܚӆ]!׸'Hj�q�.�*'�iy̒�5\��㴤�\��*�F�6�b'{�12saC��y�C�(ބ���Fݻv|��� 99��Z�M	�=g��+�a�Ĉ	���	�1@q�	l��i�Lw�2T�U ^"!���ď�+hn9X�*���6��&���>� ���&�7���b@
�+o��س��*kf)p���26�!�a
"��/�#bz�y�!�"��#f/E�gw�y����vr`���+*X\5c�N�4^�x�QG�F�H�����Ig@ �+!�	1p�pƦ؅*O���6t�@�It(�a���8������?����3OJ�����J�pMB&�:D�(�fD ,L�U"!ȩg`�P6�jN��r�'��:&��e�j%�v���A�	g�b��Z��M"A�������gB@C�	#a>�1�2��9H��R�٨I�Flʤc�*g�C��.�����I�$O=�%�B�P�'��ł�a�ٛQ�OE]�h�e�R!�WC�,��Rh�!�^A9�L��m�4���3۾mb���7�Z���Ǝ3�p>�V/x ���Í��\���M}b ��lڅh�☡avz@��"N�zѠqƜw(�B�ǆ6z ��`��ӎL�P36,��K1�,
U̓Oh<y�� -	��,g����U.491Rb¼=1֩:Z粉X#CQ!.
��Lڐf������ɼs�/WKܰAtEU�gi�l�'g�IX��/��t���&��I2j8A�O��ʶ��0
6l�(��c����å	��� ��J5zF�ΝŪ���Z�hr��K:L\+p*<e��ak>���eR�J�NH��=a�$���%P�����J�<'lD21�ʊJ������9���K��!�����,�*y,����䎴B�a�"K�1!�0�Um�
[��L3t�P�(��+�ϓ�Y�h��U���D�U��+�%�>���X��TT� XD;g�U�7	�L�Cm��g;�]�sA�q�Za��	=$���V�́
`2\��9mc̣�B�*l��8��FC�H��dA<#����LM�
b*p��8nf杨;�zL3�"�� �p��H
N����Ĕ�G\l�UU�m4���bD<d���G�R7���cB�8a.D�I�\<
�±MO�]�[A���EC�������\��U�v�\�Z&'�^�n��?��+���x5H�DȨ�$��լN$���Z1˗�LHl�"==���i�Z�^�1 �E$-T*���Z�U�`�� EXLڊ�D��<P�r�E-R�^=�
��\�`��B)K�O��(qe��/Z  p�K%z�.=J���6g�/
 s	?K*���Q�Т^�f$��FM85�p���Z����gO[�u�| ���̔`z�	��Ь�U8�, Y��dA'ړG
����ڇp�j���͖et�)Y@������W
(�����vg@-���:|O��A'�� 	a���SF�'7���HƋp;|�K7��y��D�Sl�lA'�F?r�x���M%2���`uK�s<r�sGoׯz���	5�D	̈́V��XeP�����2��nҹz��h=	����)<���)E��	y���*����H��|;�8I�jؑ\��ǈ�:}����MF��E|RޤU�.�I! �<h��ȫ�nP�A��Yj�����ۆɍ�9�8�^�V�"�aq��=j��ܛCNтD��}e�!f1�@Z�-�9d��]Bso��/�^1RF��$�0?�'�GG�UR7�8 �M�Cc��{!ZLHD�%t��{��<?�9���DCO�e"7h;�a�Ã��] �]z�R�kBgN�X)�4Q�����I&*H�(�eO ;�l̓u�܀J/th�í��;^,-�3�F<[-�)�↕9�X$l�Dq.͸�9 �V��B[�t��ɤm�j��q.�A�,����V�x"<���K���q�] "�0A$I �����퐍w��Y�҈U]�L� v"��J�Dp�ܥ/�^�E.�f/"���H�v�Σ>�4�R'&xf�צC
V�X�ӐdZ	M�(eBҧ�yj4�P��H�����''zb�ǆc��z���j#:��	��jٌh����<@z��b��C�N<m�֭�v؟t�����L��iBhJ%�aɣ���?�L�$���y�NX>�:x��¶N��i"���?��c�Q�5��%vݸ��:^����E(=�O5��P;�n�"���i�U��%q��#�Q  .K��R�AO��~b���qZ���Ԛ��4``��p���(&�@��5�� 2`�D|L��mܕ��_Ȧ��@h��#�	ƾ!�m)��c�\���4+��I��F��dN�hW�xr萮U<,��͘p�`�����DA�fiĀ�'�`Ԩj�'A�4 Th�*LB �X�����@��	�]~�=��'���pY$�,�j��N&>�4�2��^9H��aJ>!^9@���~�]�2c8�`&#�_�@9��N�ݜB�I�	.�IU�_���[�DO�p�x���P)h��i(���T��5��gܓu-R�Rt�ٌhnp S�B؇��-ivp A?O��A���}o |B�.D�z���*]��9@�9����&E�Š�-N�T�������@⑞
jb�~�(J��S�Н3�%f�]���M7{�t�`�'Q"DsGb�>=�e�w�@q�`�0����ҍp��S�IRxU夅�n9�%Jd��V6B�	&<�8H:�*�7ξ�Iv�����	$b�J}k�}��iS����[�m�����M8G8!��]�].�6�ۧk���D�_8!�dL"Cd9����#GH��͉!��խhЈ��rI)I��D�r��&h�!��	���6��@��LgK�P*!���tY8��0-�9RILy!�Ǎ`������q��l��iR�!�DX*�za��բ]���R.�<i!򤚢_g��ǈ�hw��V+�&B�!�ܨ0$p{���-r`��q�j�4f!��1���CHVg�a��U� �!�DO�# �-�:nF<ZwH�!yX!��=�lL��CKF&v��5���0!�$	!����菑1&�ٔ-��4 !��3<2������

�a5E��@-!�M9Z3�	�O�H�ID�G�!�Ą�;��9򲆘�[	T���CԏI�!�5.�,,+�M�"��p��ŏ'f�!��Zސ�##yӆ���DW%r!��;xͰ�s͔�jҨ �XKE!�	��tk��ɐm� ���ӂ@�!��[��Dd��#L"� ��M�!�D��7,N�3���gMt�`�)J�!��ÇH�`[�g@�\D8(ӤF�~����	�蘉�T"!�(h{W�0�y
� �pah7��0)4��4{�.�%"O�	"��x�

�(�^}ٗ"O��C4wq@�`��̾Q
�
t"O�����	� +��$��g�:I�6"O
�{e)b���a�R��V"Oı�7O�B�~E	aF�_�^�Ц"O%A�m	�7)�u�O�T���"O�q٧蒇9>t ��K09��E�$"OnI����o��q��g�<&�>�Q"O�C���1Q`ZY�df�5V�r�K�"O<DP�Q�o#�(j�E�&�y��"O� "'��%�~Y�TD�8b���W"O��q'"M�|�rdB#�22���F"OD�eBF�D��B��
$�4��1"O�!;Ć��Z�v�
be��)�"O��%���Tт',�"R\� �"O�j*��7�Hfx(�q�R�{!�"XD���CK�u���)� ۏ|%!�/*���@�Km��ӱ�E�!�D�(	@�+��כU&�=ё)ڑ}�!�$�Rc� A��'$*�eCi�)�!�� *��!B��	"�R)�hp!�䚖 7�:oX��2�8�N$Dv!�D ?>�\A* H���#�V�!�D
|Nr1�d鑢,o^3����!��OZ���(ٞ\M��T���!� ���)A����ɥ��rR!�ă�]���E�B�NJ�j��<3�!�\(F+��b�� �`��b'��L�!�dΛMX,y�@��c�������=#�!��Exy���W�I"6��q�i[�%�!��47ix�£D#?��q����+z!�d�9d��p�M�2�h!H�h9_}!�dH�K�p+S��X�j!�3�̫�!�ӭ<}�|bA��'=�`����:8�!�΂P$���1n�V�I�X�B�!򄟨e8�|�G)^'.���I�� �%�!�$W�C&���Μy�ڠ�E㕍x!��Y;.]~�;bJ�8+z�H��A�F!�$�z��Es�`�-g�
�CR�T�!�L�iǒ�J�a�4m���n�!�$���xb	�mn�K# �.g�!��$`yb7H�)_p0���U7]!��Ol��B���'R��p�� D'!�DY�'F����
2�����A(}!��-�}F툈e�^)X5��=�!�Dݰr\q�al���SJ� �!�D@�.��C�
8VH��w�M�!�$�	�nh#�&��tvȒ�IN��!���q�@������j54�4J�!�dK�d�\P���59^)�7]4�!��6+�y��͘q��+ ���!�ڙXe2w
	���LR�
�c�!�E����:��<x��Щ�K�r�!�$�uؾ����� �<�Ӆ�ٟ<!�D͒Yx�%0!.��!�A��3!�H5��u��X�g�9R!������B#�L�Vƌ) �!��Đ;��e�s�Րt���h�e�$p!�dY%)�e�l�?R̢ �aCZ�.i!�X���<XqB�*�r��ܫx�!�( ��P��_@�1� �!�d
?֤,z"+�X;"q�4ς*6!�� 2��Tn�		�yhRĒ4Q!�� �Q@ʛ|ZT����H=4"Oftx�G�2�t9�@N]�`@����"O�Y�׍�)���y��?C�v�8�"O@�����e���&͈!�lu��"OT��@N�.G��f/H/5��5�"O���̲s^&��h�2<�l��"O
��&GB><x��M )�tA#�"O:i�so�O��Y�@-��;&�Q�"Oz���BR()ؼ
�lؿ"t4��"O�B�T	O%���"�5�\HX"OH���WN4�7�5VĴ�C"O��`l)G+�	 v�U%)m�v"O�h�Ɓ6!��
3��v<J�c�"Om����4fw�D��-؆vZ�{E"O�YY�n�',���$I��Q�(�!"OF娤×F��x�'�!ĺE�W"O�\CO�S'<t�ܛ}�����"O.� 
�,?I���d��5p��R�"O��v�5)43c�X&yk�`��"Ot�h�@!lzT�����".�Z�"O�-��"�6p�X��c������"O6L�aE�,nT���"H &��āe"O�1�W�ǫ7������P?!����"O�mff�в�h?°�T�P��y�I�c_��A��{�mG���yB�H�Z�P#D6���x��S�yR�N"?���#7�̀?��a偎�yBlZ"� Ń`lS�E���8DHˁ�yr'8&.���!�� :�;��%�y��F|� �:�/ۡ7#��� �6�y�H		!����%�M�&��yCĝ%9��5�9ACfI����y��*@���-9ܺų��ҕ�yR	�4���Y )�>�~tY��Ҕ�yr���5	����nˎ3*J�����yR�ϡKN�My�拸8:��`�[��y�X�VE�;0"�>7�@1b͜��y���a� yC��Ո'�4�9�F��y��@7Z�I�&C�/�dX�NZ��y����:��\c d���P⠇�y"�у~Y2����&Eh#���y�aȇg�)��,�/>�F�kpAR��y"��YN�<Q��K�\p
G�*�yF�FJ��m�#zjQ��"O��y©�����5�D%y��д�_&�yr#M�q�m�Ќ�jΖ��� �y���R�<r Ǖ����!֜�y�	�n�*�h%L)����ؒ�y"JB�U��
Ç�p�&ً�.±�y�*�~l�3T�\<�!���y2+�s�����k�޴,�`�N�yR&Z�X���I���i(FTP�Z��y��Xav4uC4J��BCEf¹��'�41��fH`���K�{����
�'�N��� Fa�A/!^�
�'�x�2� @ĸ(��$*  �k�'���{E���vf�Hs�M
Z�&���'x��꒘n��ٛ������8�'���w傥K���,a�}C�'����E!�H�x�c��	����'qb�l��*)�$��"�����'Ҙ���B
*dH(�4c�7	��'�L�5%�3��Zw隅�|��'Ƃ�A`��HXRK����"��� bd`oD��
���Ч;JB�b"O` aFO.Ib�C����F;�M�A"O�-�ħM-|�8R(�jz(-�"O�/�-s~j�ئ-�"^����"OvI*ĭ�kIްZ�I#��ݠ7"O�P���39�>sBW����)"O���DMP�;F4��C��y6e�7"O��z�JG?i���Z@�dkzI�T"OHl����	P�f ���P0�KV"O���G_)M���XWh�!JO���p"O��BwOZ�h�=S�	E�w�$2"O�(�TH���,�eB'pe�+�"O�����;��+������"O��������*BG��%~L��"O$�2��R�V��|��& �3�걺"O�܉���8${b��*�y3�"O��@�OއM<HT�K�R�iS�"OL$�B�3}*d����B�� kP"Ox�
Ae1Y�r�N�"4`ʼ2W"O4 �T)C�r�����cX,Y^�)�"OP�pJ�>3X\1��*0RR�"O:�(Vn���M��L_�d*|8zu"O@�&{��\��kS�sh[2"O���
�aC�C�Gz ��"O:��Э��r\>3����Ga4M�T"Od� �5J��0����G]����"Od�X&�	�F���
���$B�*�"O� '��7�T �S�K�,� "O�8Q��F�JG�X�H0�|�7"O����,�I��*C5\H��"O|��BȑT����_
B$�� 4"O�!�"č=ut�zC�?M, x�"O�4:c儦(oX�9�dB|T�Q��"OƍR�o
8>&�e�2���LW�-�"O�@�醊	���1AJ�yGfM"5"O*m��E��bo�%�w�Nj��"O�M�2(U�E�8b5霅k��L·"O4�`��=:o"D�uh�Xk<���"O�����*弅�է״OW��:6"O�4J�=|ޅ"�(Ne1`Y��"O���¬��dOx�ևE�r5���"O��I��9A��<����r��"O&mBA֘���"�+�u�G"O@�{2��;;��bg!�02v��h�"O�qZ�'�1�`��T���p"O��I��vJ�Nb\���E"O4j0�G��9�!LJ�M��X!"O -�&Fԑ&�����,>A@�9s"O�p���F4$r,�Q7�['HF��x�"O�}Q������$;_2�����tB!�䌽u��Yʒ.ϷO7X��A�5;K!��V��ƭ���T�	�$�ܑQ!��SZJa�b��&y���2&�!���ՠg̝%O�޴Ҧˣv!���}'�Q����d㪅�K�<c!�dZ�%�@�꣪A>ѪTi���!�M>�уg�N�V���k}D!�$T,i�0k�䜰rvd�s��85!���
�d)�H�;GX��'�O� !�Dا �J��B�ɕu���ʞ�`�!�D*+�&�*ˤE���(���L�!�D��b�LW�X29�4MJ���!�$�j̬�I�%�X����N2r�!��
E�P����-]	
�&�L�r~!�� ~�Y�K�0/��V�T(.���%"O���dF76lQ����27Nj���"O�5�QDC������ Z7��Y�"O�eR�Ф�;@H
^�¹�a"O�bf��J=�i��Փq��T�0"O�ā�W�/��{eC�:6c�Qp"Ov�����X<�|S��qBlt�T"O �SO�Q��1��#ыF461pQ"OB�|?`���\8��Zt"O��#�Ǚ�=X�	��ˆw�D�"ON}�g �Z� G68�陱"O��I OW!���Ү�r/�@�!�G�.�t`������qQ�9[!��ڂt��B�&K �� �O��PG!�D�:�s�E��H�:�cM��!�E�.�j�hŧ
�(�<�xD�ڷ`�!�Ĉ�Cf�3�%�7d.t�@�)�!� d*D���9`�y��B?\�!���O�N`��$�++6�Ӭ
r�!�d:+u�e��K�-2d� ��=!��
a�r8�vhŁc-$5�j��4�!��Su)&0cE��&Q�F�b0b��H!��M>*�8��g�K+|��%JA89!��W�x����G����釼�!�DF�'�ށ[t,�7d��'G��&�!��(e"ZP�v��~s�r�A��#z!���8�yӧ�F.3R��җ��c!�DȎanZ������`�$��%r�!�Z�h��!�t�Ċ��Wctw!��\;3�jՑ'a{ǤZ+ӓG`!�d<q%�L�EÞvn\���*�Vd!�]G�,��V��=/#<�(�6�!��?T�0k@�ΫA.n��ꍊh�!��ZTɐ%���!: �
H(�!�N�^��4*m���uN��O!�ڌ>J��˵ ܦs2L��@�U'*!�G�4p`�L$�]�Q�ͣ]!�D_�m-zx�(� ppԏ		!�Q"�L��Kx�H �b�!���a��Nn���n�����"O�����g���p�k׉\�0@��"O�@i$+�6%�ݨQLV��ly:@"O,��g	�3.���A\�Q�za�"Of��oL�R���z�J� p����"O�,zw�_	(`5Y�	��`�u"O��b�n�b��O(���p�"O��S����D�^A����SqV=[�"O�B��҆w� ��%��O�D�1"O�q�s´B��`�c�ۅ#0�0I�"O\��!�U9RFp)�@�#o���Y�"O�ͪR���5������Ys�H�:�"O\��3CD1C�l+���+��&"O�	H�@ӗ��!P�����"O�ո$�M�>��Uх+�g4r���"O�<9B�"�V�zD�R�VL���"O⩱&Ü�(�I��J1t���"O�����G�Y9#��p�@�#"O
P{2��T&Ȃ�����w"Ox���\�*C*Ѩ�EU-:�ܕ��"O� ȑ(��OU�d���9O�v�Y�"Oΰ"�.kA�MJ-y?��"O~�Y4Kȏ(޽;&�M�f����P"O�������TF���g��'��#!"Oah�Ɉ3`� �B�ň�f?r�k`"O� .l�C�C Nz��%�I	x��q"O��e*قS?X� DW.��"O�Ѹ��9F/�91Aȴv�Y��"O�H�5�\�L����� +�l�b"O��[SL�*}Yn}@15�D�"OF�2�FԤW�PP�eɀZ�mpV"O�a�(��$�(�BKٴ��p��"O ���,\C�5��$A�&�:�A&"O�I�JH42L|�⤊�j�j��0"O��C�-@���D�w�9��!�"OEQ��ї1b8�i	N#vd�
�"O�]��@%t���@W鎫K�p����	&�h:W��s������8Ӗ�D
����Ó��2j�|�F�ڑ*,�	�<x��"~�� �M�^T�%`�zX4h��/� {
�$�L�l�������^4�>9���-X�p�y�&˻)��j�n�H��Ԋ��'i����-�!V�4��	Ø1����r �N��8��N�l�2��/Rh�d/�
����O���Z�m\po�ɗ�	^� �3�4WJ��#� ��](�kQ�x�a����#J���^/t���zF���{��9��I �O���JG��챏�~�w�G.M�$��4I�闸�2�`Ē4L3�H��1p����MG�4M� ���`m�S&|����;"� @�ˋFФ�1u�W�^�򄱋�Ě~Z#M�5��}�@�֥F26�2t�5�eP���lYb4CèCf>5���x��ݸ�Ā�^j� A����J����n�KI���O�D�:M�d�1�d��V˝�yl��4 �X��u�Vf�i�ލ��Hb�%��odQ>q�Or�|��L�.�~�@���Kt��3G��k���ڑ�G��Ma�β8ca�DJ�C��D�N���%cd�(_��41��Mà�9d�.�����?7��H��x "ŏ
*�[ƨR�X!�����;?���%����O��.D�p��!N��F���s	�'{$�S!�O0!T �Ыժ:4��q�'A����*��0��0�d�Hq��'��ɨ��"Z��A�P"�:a�<h��'|RR�K� M�0H�[�>L��'�412��#ZK@�kP��(�"�Y�'u���PϜ��pR�E5\>E�'���aF��;Q	��A��
 ����'���B�&sy2"r��FtA�'��Yq�=VxE�Q��#v�%��'��*2ńu��DJd�^�)s���'3���Bq�dz�+-+zL1�,D��BL�31_*u�	_! �XP���+D�@Kp���!qRLBB�,P��$D�X:tÅ?Rjh� ��f(� 3�#D�3���D�,�D���w�T2�!D���"E��r�@�F�
=GJ��C�>D�����;h�Ȁ��T�4Դ�&�>D�@J��,
�R�`�ԇ��}c��=D�����G�B����Q����#�:D� �Z6�����gL�e��c�9D�x��'�9��챠��.j���� 7D���&�@�.�.풴OũF@*�X�J4D��k����4���.'2�˔�0D�Hj�ͳkÆ���)`��0��.D��ಏơ@�%[�f� ���+D�8b��V�>�� �AW�0y�a�VK*D�4 é��cg@Y�Ġ �9�ҷ�)D�(�T�S!-<����b��$,���DG)D�d�0�¯F?�`�$ي�V���%D��P#GN6�$�D��w��J�"D�� `��`鈙��`Ɛx����?D�D��� �piD�n�6:6q�� �y�<����M@��k�'β��m���o�<�f%i��H���ǣ=�j�����<!%�$�z���`�Y���9�oU�<��]9ʜ���D��y+��Y�AM�<i2�n�d"k�0Q�~aAq��L�<� �22�P�n^ޭ�b�;'G�]�1"O�qq�/����ؒ�F�%E��"�"O�Q�r!я.�`I���	*R�� "O���D$:Z�4IvG� I �
�"O�	��cՈ['��+\����"ON		uh92�[BjЍNeB={c"OzXAd�Ă
�D�s��5$B�"O�"�#O�@�@A�&6Ȯ�9�"O�Ps�h�?F�TLC֭�6T�i�"O�8W���<f��Mɩ@T��"O�4QĨZ9a�F��$��� "O�l���1��u�&$A��)sd"O��b��m˔�
 ���J���"O�[
�~�d f�^�U�8:�"O���I�\��t��Y,=��aJ�"O��S�X �� sX���%��"O�B�*��G��9���=����u"O�����$:�H�/{ �`�"O����љsL�&k[�\#8�"O�Y:�@�6m~��t��q���4"O\Ie�Y�bO�xӧܿ�����pE{���_���Ye�}������M!�dE�,��L�(�,A�V9#�.�*}!���S�^��E�y���rm� ,!�d["�̍��C!Ʈ���Ɔ(!�7F���Y��V1H�ј?5�!�D%N �p$�(�ܡ�V���7!�d��[P����Ǉ�tU&��W)Px1!�D��^�Rq��c�bRb%�֧�!���<���qg�ެo���R�d�?�1OB��D�	L����a��)���!5ʕ{!�d�F�h����"�Ā&��,!��^c$�0�gW�x�t��&��;h�!�ğ�'����Sヮe��y�5�!�R�r�$Q�`A�	���:�k	�/\!�dT�bh�%��%p@�ԪA��3L!�d� Ru�a �N��(L�v��vD!�@��~��R
G?b`�󫄺	�!�ߚ#��D�'G0{�*,�hT�Ik!�$�)9t��b�	}��p�h�,p^!�$�1(o(�P��N1|s��eȄ5ez!����x�!�Bi��q�]/#t!�Ć9-INÒg�7+|���& H�2!����k҂θeV����U�!���H�����yT��ʄ	[��!���$ �����[W~��e���pI!�Q }����@%�`\�E�c!�,1�6���a�%ANEI�M�6�!�DQ�;$16�p%�@��/;���ȓza3S�ux���,�s)�}��1o�Q	�J>ww�xyB��|>���c����э�(O�x�@�lj���L�6�J��J�0���0,�����ȓB�V�xG�#�ً��_R�<� &ב�U�e	/���!��L�<�E�9\K�L��
�K%��9�K�<�g U,%hv�f�4�*H�2 �G�<!AM�-���r�Ϥ��8���E�<Ien]1�LT1��P�igBuA�nk�<q�	_/v`��d
E�j�y%bTp�<) !wE�����6V�Z؀a�i�<�fO(l��i��gݪh�r��w c�<	SoZ�c:.�0go�N�*T*NE�<YVI�9c�b���b	�*yL�RじY�<� ��b�/Ȕd��0������"O�upRDT�V�Di�V�ڣg���bs"Or�����=e� 4 �˙n�H��"Oz0����0D��ǦJ7��,�T"O�`�À��u�P��fD�L�2�	"O2h�
��a4��)�X$x��"O4I�V���=�T�ɲN��P&"O�iu(�[`���K[�K&"O�A��ዹu�j] ����eX�t�"O^�+v�	�y� �("j�k��E"Oh8��ٛQ�������)�L}c "O��ac0���,!����E���y��X� �d���ny��9�OZ7�y�1�Ș�`�׸7�����M��yb���6O��z��	�C���y"DR�n_8���#�B����ycV���t�A 	ȵ ��yb.oì�xUCP�'h �p�[
�yr�o��j%��>5�*�n܅�y2��0w�X�4�K�)`��Ɖ�=�y��� �x �3�Y
1U�\�㋋��y".ѣ@F|���J&鞵["̴�yrJ�=�J�D��2�zT9��y�:�J�Ô5y�������yb�^7'J��$[�(�DA�q�G�y�j[WD�����Rtx �0!��y�P)��B`�O�K�Ze
U؛�y̚�z�!�"9�2��I��y�%��j���a�N:+y�a'�y�a�o���2b6z:�uB�$�4�ya�0A,�BaF��x,����G��y��I2�<�V3wbڭ�6��y�o��\��50���9�f��FmE��y$6�@ ���/��8*����yB

&f�x�� 4& Tt���̇�y���e_��x�DY��<�"#�܎�y���k 5��W�B��R(��y�ܬ4:f�6@x���# �"�y�
gO�I8'#բ
s�p��6�y�O��Zh�C�����'����y�oF�=���q��<
��(X���y�3T"�4,&`���g�y&���}UMV� �0h�e�"�y�
�g���"���hu���h��y�$H%)��yQ�j�d,�9PV�y��3=���C�L�l%�����yrlݱxi���F��;H4������"�y¦�;ц\c��R�P̚�P�#�y�BJ����T��$sJ\��yCփrr��C`ǌ��T�C�y"���.V��@�HW2B��y��o��y�e�F"0LP6dJ�:~�H �����y�#܀����ێ/�	Y ���y�F#���%�]($$$Qxf�!�y$[9QfXر�+�j�Nq�B.D�yr�3v���n�O�cW���y�2F��P��!��`��C��yB���"�$���&'�����y�A�c_V�� p:4xuF,�y�!���A��8QT94mǬ�y��N1gLH�P����&��$��8�yB �3r6��x��}�<P�I��y"kǧ��l����g��m�����yB�V&V���2��]�5���NK��y
� 歱rGP�p6VՂ� j�:I��"O8�#�,�#O�H8�"@}��@P�"O8q�!G�(vJY /55|R<�`"Od�	w�ԑD�,CE.ϜD~
Y��"O,��c��g/r��m�1tF� ��"OFPÑb��:�f�
#)IC:��&"OI8�E�<��S(�RU,A0�"O����	,\�v�+�l��l\ř"O%���,�nš0��NB��"O�]x7bP�pd��dǏ(��cq"OZ!Q���`��@���y�x��"O\%���L>n_��q�M�� �q"O� RF�
$����V�H�n�����"O2�B�#��L0N��h�=�����"O¥�F�=��Qd.
8y+j�"OBx�V�ŐZb����� �f"O�}Ra��4&��]Бm�
�mH�"OXMraM�0$؄y����"O؜[EɏV�iC�̏����"O���v��V䘊ekT ��	ڂ"O���f��/D��Ո!��1�1"OڙH�w��%��bZ4F�~��&"O�[��߲u�x����M��p�"O0�A�t�Z�68p�=q�"O��$�r�Ұ#�F3��0�"O��)Z8��&�#Mo~m:7�	=X�!��Rι�T%I�&n�r�F�t�!�CiΊ�
"�.H�9A���=�!�#6��P3�\ A�=�SJRM�!�ά'�.t�5eϼV(���
G?!�O�P'@�{Q�?8�vt��N�%A!�䔈q\��
��5��e�CL�1!�K�!�y�a�0}���	F�_8F�!��9a$	H#uP���'v!���������v��`gf��!򤃂3�R1�� �5)�,�"'儓A !�r@�)J���2b5j���c�I�!�D�f���s�03�����\�!�$ǕK��eR&A�MH2ɑ�δX�!�$A�#6d��WK!(�H��Q�ƖH�!�$кX�	�� �/E�P�25axr�'���qc��Ħ������Y�Ι�Xmΐ�ƞ�~��2d _��?	�2 S��?��X!( ��<^"8g��9�^��5b3f|}�0GZ!W#�
��&jLZ0�U!\\�'W���V)oQ,�C���=]L�xҰDo+,�j�@؊Y-���DD˾<"�ĉU�r�'G. ���1*�6B`��6-�-0��B���I��������K��'l"��?Q�'��ʀ�N'��mҕC�3OQ�ٹ��D8��|�q*"@|��@[�$�qb��E�;���i��ɼ Y�U��ӟ$��A��@�>P��!QbB��� �O����I=P2��Ob!��Ȕ�7�FL��_X'�iA��x�j}��~��Ld�J�"�&�F�P���@�I'!����:)(�rjS�g����/{��
Z.x�abHE~���Q�?q�\L
n�$/@�I�~�H������)k�S!Mt�v�i�*�k���&%�������QGJ��&aqk_�GݰEh���~8�#ش��f�'3�6Mn�<%���ѵmd�Tѥ@ �Aqi��M����?9�3y*5G� �?����?����}{�]9.^
la�m�dv�0����?�E��%͞?�B8�ee�h�r+�Z�)�)|i���'
�s�Ep��S�L?B
��Cf�n�2 J�A��@3��9eq��H��ռ���ٿ�����O5H����̋���7-M@y�D\$�?�}��ԟ�lښ.�d+���ha���9R���i�R�'���0�K�$�(h�"�&R��aI�'[R/c�&Un�~��?A�So}�bڼ.��e6Ö���\�w*X�,�r�S�S>F���O��D�O�E�;�?����?�/X�V�*i�V"�a��s���3� ��*�CM�$y5^#'E�x��&D�b���Eyb��(%{|�� ��_� �[@hĀd2l���i8
Q*���yX�)1Sʊ�e'D)�#<�I�)H�e#ql["X].��sJ����؁��ONn��ē�?����'�(ڇ
3�X-�B,E�M���X��/,O�<3��E�EA
}0�Ú� ŀF�Is���M��i������ߴ�?��t�? h!!1�ѫ+�hr��ާ/<	�u��ٟ����w8�9������?G �S���;#C<�#6&�&�4S��\4d���bf��n!D� F�%�
�&ʓx��hKe��~U����)��0%�b�Ȏ$j�a�mj�0���<�g�|ШR�GY~2b϶�?aF�i�����3Hh�rIJ�T�0����1l���ܟ���b�S�';�fū��]f�B��P�Qd��EyB�*�
��!x!Q�*H�5��ថ�� 7	,%��Q��H���M����?a,�hiQ iӞL�C-Z�n4N�*dG�b�D���П���,d�m�8�|�qСW����*]�.vX���<��/�=�(*5m�wm�S�x��W8+�<��e��p�<� 1�q�d���c�M��	�zt��o�;s��p�!���� D'�����O�lڰ�M����O�~��`EֽL�@�مN��  ��ON˓�?Q��?�-O����O��2n���i���T�&���N���p<�7�ixV6��O��nZ¦90���[l��C��9���eA���?���䓈�O�A���  ��     �  �  %  �'  �1  8  [>  �D  �J  -Q  pW  �]  �c  6j  wp  �v  �|  >�  ��  ��  �  H�  ��  ��  J�  :�  ��  ��  �  S�  ��   �  C�  ��  f�   Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�� |d��"O
`�(�;���8���-0��1%"Oj4��ND^[��"3/9�0|H�"OB���H��*�ʞRy=a"O�味V�!X��!&F�:J�$���"O,��a
���C�Ą�M�"O,$3%o�-���p���+Ն�:1"O��ݢ1����`���y14]2��i�<�6��{_���c�H�`�fX�$Kn�<��A̼VI�xR[�)�Ć�pඤ�ȓA5��('nߡ4�� �)˩%� ���,��r�؊b#`T�eT09���ȓ!�b��g��}�8�F��-? �ȓ
K|m�ș�VṔ���2�%�ȓ"R�X�j�4JN�1�˘X�i����̹	_�jZ��1!g��zܶ��ȓgil,*�J�
j�Ne��i�J%b���f	�(U��:���G��$Y^م�~r�� S�%T"���k\�jx�ȓ|4�1�îJb��@ӵ�ݩn�V��/[`�"�v4�R�!ʎ<��M�ȓ`:��z�ؚh�J�Z��$HY:	��H��p�m�C1��!��B:��0��EnjZA V;9����J[
2���	��4'J�EA�IVW&��~�(aZ��ӹ�>� o�Y�|�ȓ�f�A�
Ο7�H��M�$�����mޠP����/���ANXo*�ȓTv�����{ ��-7�*h��I��sB�8�8���3����ȓNe*M�悡;������X�o��!�ȓ'lj�#F�m�+R&;�|��2)n�C��0S4���T:
b���:�0!��e֊��)��ͷV��,�ȓ0�&�8#���� ع�L�����;�P�AFd���,w�6�F{��'O��V���&�;�+0:��x	�'%��"J�[�]�R�K2r��"
�'Oe#W烹�R}aC��z��
�'��;��7�������L	�'�:<*b&K"4����M����9	�'نx!c̓>�D �,ݻ2zX�R�'��@ �F�9<�m�7I�"+�a�'ր����>��Y�
�%&���'��0��3L�r5��M/� HJ�'U����J08fx����I$p:<���0��j&a��'�L-�I��w$��
��Ig�<A(K74~<X��.>IG�t2QI�~yR�)ʧi�n��EiY����3e��c&�D��f4���W��'^�4�KR"l&I��y���.��~#S�˩y��)\ ; \���EU"�D`A�w+ Q��\ ��/��i���bND��xၜ �.���+D������..r��nE"gp�`*�H)D���C���*����e��b���S$D�0�@%������ٰ �4D���HݦeF����� <����ķ<����,f�Z%F��T�:��4��4z�^C��*RA�C�呅[w  Rcífc����Y.< (��x5\;��*�ڢ>����*���?�Yw�6�MðQp4c�#��5>�K�'4�� M�G(�X��ա-�c
��� r��QIG��L�I����"OZ�����y�S�+�1tYL�p!"O��`qaʜg0�bj��X���"OTQ���[(�qJ2`ʉARb�H%"O"9 MP� ��#3!+L�"O�����@�Jl�2B�� �|J5"O���6f�M�0��jI6�b����'(1O� 
����8�bgJP2I�Ѫ�"O�)@!+��9tL��(� ��X/�y��'�=�����r���#�6�K�'�8L�W�>R\��I�6tP���?O҉#�CĵOH�p%��.^hpf"O�q#��p�4#5�۫ߢ��"O�<�bi�(�¤@�EL8#��R��[�����)�~�FJ%ᖰ'Ƥ��bC��y�m��Kk�Y��� �^�)��T��y"����<�W*:o�̩�l��0?I/O�H��kA�<P#�0C��p�"O���B��A�b�,B�@M����>�S�4g�9j<��UϞ>7�
t�T�_!򤑦nRȅI��Q+Lߴ$��삂z�a|��|� fT�!�n�a�Z3���8�yo�,1H���ǡh�8��D֔�y2�K=h�&�)[��$۵�	�
�챇�%�Ȳ���	�L�3e��K����?�����w�ɟUp��o�5w��Ԇ�In�'�*�y��(��Գ �U�vi
�'��m��C�`����	��Q��-�ד�qOH��c��,X$�� �ιVd>�pR"O>�!��<��;�!��7R�l8�U���'��#=%?u��k-@k�਷"B�n��>D�X0����bp��@6�0�􌼟p$���I'Nn�����T3������>���<�ґ��Puv�����.wBjq�CMY*�y���[�p�Q���!w��QRbQ���=!�{��5;z"�!GanU����ٸ�yb&�.Z����#�ֱ!A�*�(O�,��	!d�t�"Ai�9[�&�xB��FB�I6	:�+�Oʇ)�|P�N �2�D6-3��f,�7$�\#v��S��`&$D�X	dj�1~� ��5k���Ab4D��"���5r���5�#y���c�/D��"C�./����c����ts�1D��B�k��}��I�����P�^pPC ;D�y��_1Bvb\ägU3w�6��7�+D�|�Q��`"��G'u.8ʂ�?D�P��O�2(0�q�i��y�c<D��Qv�I�/( KEb	�rvx� 0D�����G�0�n|�� ��t��h@�0D�d;����#�4|Y��C�*����2�/T��{��.	�Frc��ukVt�7"Oʹi���G����̩ikX�f"O�\@�G���I.
�TRh�z�"O�@`�c4*��آ��\`pV"O|=� #D� �����:LMv��q"O-9&J&T_�ePL7 H��"Ot�b@�J34'��:K��-�A"O1�rJ�!.2$U��i�v�.�@"O�D��&��ݡ�gƥ|�ɰW"O�:�lW�nht`2`��gxN {D"O���W5 ��8�e �+��T"O���� )O7���@�jz|T�"OF,�L�5%�~��F`օ1wx ��"O��a7!��.ծ�fO\�g011"O� $���%%
���iᤋ$?yTв"OLRg�\�+�y �)G�=]*�ӱ"O���L�5I��9��(��<Ph0�"O8yk!���)�J�:Db�+�2x�"O*`��e�lJ<�q���!K�����"Oz�av,�� vN��o��r�"�w"O���W��\�Bq)���1��`�""O��`IZ�Mh�ڦ�ƴiW�|C�"O�%��$�>6Ac#��A%bP�"O�}��Ƚg$:�D�
:	x�@"O��k�kʱ2 A�u�Y:6�N���"O*��T/��p�  �2�K�����"O<pHpċ��u�0ퟆ9M��qQ"O�Q;���"]h
@:b-�mC�t�U"O&t�/ߨ�2��+1@�9�e"O~<�����*d�2�+'W�:�"O"���\�>��uc+,�lZs"O�<s��SD��CE����"O��Y���
A8�i�!� ���"�"O����[h^�Ғ��n�|(�b"O�@jsO��zUd��E�<����f"O��0�P7M�V�	F�(F��"O�&8�!)@$]�&�J��R"O���GΏ�+*�]�g�]�s{����"Or0P�&%�{$�"-4�I�"O�X7Q�4�l���?3 �RR"O� U�Z�kМ1j���j�AF"Of`���L��A�"��2w�����"O�X�A�)y���!�M�� "O&�F�x(qP7�U�R���"O���@��U�� ��0H��7"O�@��ߢ5���B�D�z���"O�yxqڎm��%��cH�� @��"O��� (UJCN�'|�pA�"OZ�eߵE�,$�ʫ
q�}�"OB�ؒ��a2����O�b�X�C"O*���M�)${�{pb�9,:�(F"Ov4{�*L��0�@^$n�s"OX	ch0,..��ϊ�!��)95"O���G���&u�p�6�U��y�Y�7����`ċ�f2)2q�B��y�"��XZ��	Pf�(�n r���y�f�%"�����)U�'��Q����yrh .o@<��!\!����`!��yr!�01�����K�����DѦ�yBH��%���Ť��,����'�3�y�)�
�5ӔR p�(b��"�y�f�Nh~�p�F�0a�ɠHI$�yb�V=+2��@ɚ�q:�$���y��0Y@�A���iـ� vf	)�y��ؿO� �ݺo����%`J��y�U������G*n���r%*O��y�̀/�`�3�U$k:�mb�L�yr�����Æ��z���Iԇ��y2���#���I\wj$�b'��yB��Q�D؊a�E6&7�M�R�Q�y���13�P�i �V	$@�I"�=�yB*vOb�Dk�/S�CB�L��y��0Tf~�h��͵O�����ާ�y��S0{���R�H�1նL�AMP�y��ٰJ�F3"��U�֬��R��yR�G#X"<�'̉�b�6m�%B�=�y�n���0���i<By�4����y�"\�&����gE�93�8�y
� �8��ß�Ti\�Q�΄�
uri�3"O&M�3��>��@���s��*4"O�4+Γc��$�U�	!
e��94"O��T
@�oN���H�=6�1��"O��8��*��S���/e*6x���'�'���'y��'���',��'#��
�*i���"��
M ��Jr�'���'���'e2�'���'(��'�r}Hq�?'�Da�A�#�����'���';R�'|��'��'��'�.e�˔a�Z�W͚��8���'db�'���'��'�2�'�2�'j&l��B�i�8����P9���:t�'��'��'���'���'���'���(P�<]Q���V�J�,�0q�'���'��'���'G2�'��'��� 2�Rx�hX� �ͤqcT�'�R�'7��'���'N��'���'�H�3�͍v�L��L�O�8���'���'���'�b�'���'Er�'͌}8F/C$R��ABX��hr��'��'���'\��'�"�'��'"�bW�0_�@qc�I<j["��'�"�'���'*��'I�'Qr�'�n��B�&U�A���o���w�'��'�R�'0�'c��'��'*�hI�0d`2��h7m�L�"�'���'���'���'vr�'���'�D�@�!�j�|F
Y��Q��'gr�'���'�"�'��!yӰ���OJU�����-���Tֽ1g|�+��EyR�'��)�3?�q�i
n�i�*D�x24�P z������d���N�i>����SѶ]�0��ҥi�H```���Ms����<޴����.c[���Wl�5��6�^;b�,T�c E�Ͳb���	syb�ӠI�B�N ;�xli���68~��ݴ[���<�'��'z��w.��J��{�|���B>Q>�J��Of6�b�P���'��%8�4�yBG�X�>�y�IT)U#���"X��yr�C/D�H��w�: ў�Sݟ��W��GQr���AA�sX���$�l�t�'��'>^7m��91O
p��◭\A�(h� �9�-z6��O|�O�p�'���i��ĳ>a�υ�*���(Q�{(�=��D{~�nQO'\Ѡs����OrP�1��4���7������\� u2�ݖ!�>��'U�֟"~�7�h] B�Կ}�}:�Ҵ+����1t�����������r�i>}�㉸��q)�4?��m����@��ͦ�I���m|~�͏q���H��ȃ'�z1#�o0�(A�k�;O��:GjY.�z�'�$�㳣�g�g�-�i�e�T-r�t�F��z�B�I^�4�r� ��	۔��#`�|��@����)p�\
�,�6�I!��Q�t,b�Ψ�P��b�h���p�E�y���
�+.1�l���0I!��y�G�	��E˓t�xsԣ[�Mi,�q`�=i�̩v�:]	��UD�~�*�p�+́1v�,�b`�k�uY���J�*��`K�)� 6M�O��$�O����D~���:s��$X!��>�H�2 M�����O�H�0!6�I�?�	Ɵ�3���5Q&H����Ͱ8�@(�+���M� !�
���'��'��$,#�4��Z�H\�$[ꉠr(_�E4�I��Eۦ��e	}����'���'��Ò�\>r=`t�J�.��;���:���O��ư4��'���՟�	'r�1�lY�P�\�@�̂_[��{�4�?����?��ފx���ן���ҟp��su��b�W?WMz郳�D�&@��ܴ�?I��,s�'���'ɧ5v�֍?�R���쀖,��AQq���M��
:�����?���?q�����OF5(&gS�hB�S�ji���w�Rl&���������S����i�N����d�JP�B��$ˮb����՟��	Oyb�J1M���%im����a��5��]�@BO��$�D�O��Ĕ�@��	�B���7l�C^�M�f��+~^��?���?Q(O�9���zⓁx�R��q+�?r�HB��=f2,�ܴ�?q�����?q5�M[��9)t�*peka偾�L��2ks�6���O��$�)�f��d�'��d��z�Ʈ#
����(Ȋ=
O���O	�#��O����O�OrQS��1R)�ѳ����	��	۴�?1��D� p�ih���?	�'[��7d� �Bg�s3ȍ9���kH�ꓺ?a@�����'2�L<)�gē]x�+d�׸RՀ���%�զ���,�M+���?)�����x�O ���pOʬdI@��a�q�p�P�dv�D����Oz�$�O������ʧ��)��*�@Q���>"�|��a��04�l���	[��fyʟL�'�Xq�7��b�"D��V���JI<��<?�����'�����|�Kwl�%�a �+�K��F�'5�$�4P�4z���⟰ � �%�6*�F�|,xl��M���'�@9*N>���?I���$�7�` �VD�l�8k�lϣ/��,R��B��ߟ����L�'~"�'���`êL�I��QzC��5"�P슁.�<5��Z���I����	ky2d� �Ӫv�|�H6�WS�\�)�$�%�&듋?I��?�,O,��O�Y3A��O������,�ZA0v%�F��+�Nd�柴��Fy�`�,A��Ri�#�&���a�a�)fM Lӱ�Lަ��ߟ�'g�'0pSQ�'=�Em���e`G6�J��Pi�-��m���\�	iyb�17��R�D�k���C��՚u{]��L^�\�z�CH<�.O��!���O�����3� |��@,ԉ/�0gɠa~�%s��x��Z�� ���)��� ���=�����ە_�0B��(m� ic1�R8�J��a��-4>����Q5���`)V	0�yxb/}�D�C`	���e�2c��1N@rG�րHr�$R�i��������
�"�)g�C?3��lp��X.���@ѫ��d*`D�l�	���`�� �R���	n "���M�0?���
S�V<@��)�'�S�� @E�rI�Iן��Iğ�[w^�'P��1�ަO�x��%ġ&2D����OL����=0��*�O������Z�,I�a�;eK�hs�jCeP����t
~	�2����d>Y@�z��/'��@��0�d������D��%��A9��z��OVUu�'���|R�'��]��1ҥ"*�T�#�=�H���<D�,9���0h�����C�db�"�& -�HO��By� =W�7�B�E-^�s��\<�1� ݧ8�:���O ���O8x�/�Ot�~>�H�&��7��<YU��S>��D��3 8�Ks�E��ЅYv�ĘO �F2�@%$�"�;t`�H��4�ToE�	���޹�r���|�VD�#�	�z�����O4Cd�_���cun{���I��(���O���+�)�����"�����e�); ��+�b�<�c(ڷ,�>9�NI�d�H��0N��<1%�i�_�� �ɘ�����OJ�'=�d��b�0Oc�M)��'� ��r�O;�?q���?�"��4$}~������~Ԝ�FI�>7r,P�A+C��<�Gf�L�sŋV<G�\as��f��S2O$r��f��~Ř5��� >�ģ<�I����c�4hس!\0D!l� �u�B=O����O�fX�1�ǂO�t�9�#b�a|R,2��N}*iɳ#�' ��ͩ�����B�0)�x�'�rR>�s�����	ߟ|�U�M�B�� �3R^�g�ϳ{���е�X�+�V�1�H�H:0<�Oe1�B�Z��$�Ӊ�(_���y�Ç8�*�@�Ȅ	���V�ΎCW�x�Xw+�S�N/8ʶ�
q`�|�]�?~hxX��M/�=]�p�kL%<}h �	��M{fT������<A㈚�~s�ق����6IȰ�_S�<�ԀK/K��ӄN۬H
myw��N�'0#=y�i�҃ G��s�*~�@��S�o2�B�I*Y�Y�I�f��%�Ǉ�=~��B�	)),ijb��}��9"��fB�ɭ���3`A*C���t�O�}�nB�	!20*�k�O���5�SG-Q�B�� FjŠ�G�[���S��ۖ2АB�I�Fi�E�r�<=|N@j�iF�K�,B�Is�&e��c^+d+,��6�I��B��T`� HR�����qa�T��C�ɰD��Ḳ*��N�����z�C�I���<���M�(��YF�
Q�DC�I�&�R3��u�h�P�d�&ks,C�ɉ5�>E��W�,�v3�+ˬ[�4B�		9��4���� � h�,�NC䉅
L �T�`>�y����:�~C�I	m6���!ԡȠճ����eqHC�)X�j���/�K�ʔ���
3AQ�B䉨[8�*��J9�t��IrH�B�ɀ\�+������*^?C��/�lC�k&KG��`��]��C��3m����'�Z�c�d�P��>ְB��3Zw����.A6�jD��a�jTrB��W�Ѩ�#R�k�0QdAK�7�:B�	[ؐP�ω[Z����4f0B�4�����2"Af��DĊni�C��8^���;���W���a+C��C��	o�$ I� :�b��ǈ)�C�>V�����jJ�4��H�@D�b�C�I��,��8�� �E� ,~�RC�	�<"}�HA�����&Y.d�*C�	���x23��:�NE{d��0��B�	 _` ���G�?UN9�s�T�I�"C��/Uu�1���B,|�0�g��~�C�I�_ls%UZ�HiȳT�9~�C�I0ZE (#���0�<�y����4�C��*�s�J3 } �3�	:&��>!Ԣ��H�{��Z��� .�^�#����y
� x�Iģ�,5���굡Y 1�f�=Oz�P�!��������Pu���@x��� �"�`��T"O�u��oU����H%Ό�*���8�E��L��z�E�
��%ɲ���Fi��녯���0?�S��8�
T𢤕3!�j�C�v��u�`�<�5�\.�rM0v���l�@����D��'{Yڀ�1��)I7���#�C�IF�S�4APcb����,h�<dpF���y�j�#�н)Ph[�3,Z|��=.��9�ͻb��:O>��X�� �
x����i��#QHZ.^èL�g
+h�!���)����4$[:�V��g��+>D��Z� Y�K�QZr��%
/�0˒�>ʓ1q�U��hґi���	��� ?T��H���e�"DبX+*���vs����@��)��IG)9!LNXb3Oغ:��|N@��6�7p�Ƥ��ߑ��dP'.`��Ks�c�@���C�����Ċ�i\�]1!#�`D�쩑�Ɗ�y�T�����FA�I�6\�3	 /�H� "�/���=�O6]�7:�y7Ô�]���tc�9s,�)b�uEC��,�v�r�KՉ~Y^mZ)F_p 1��$?ٲJ�l~`b0jE)Nz�8�';ʓn*P�Pb΁�lCf��`͎$w�L@��23�le6C�&+�$� aJu�L�H`Q�z0as6�ٶ+yꈨS�Ϊ�䛥'��|�	[�1B���$�c����e���DY<G�����et4`�7jZ��������=j��"s��X�̡i��G��y��/om,�7��^���e�1z����	���=�O��m��ywk�m=��iS�^�Y�HU���D�xrc�-7��s��&P)0��rAIh*r<��O�aqE隢L�T�z���9��È�DFkbS�t:��1�+rAax"Ȉ�m Xɢ��i�ܐ$/�1\z,�f+�<A����AR�a�`h�ƭע.6�� `8�4�w7�(�b��J��Y�@ -?A�hǵn�	��i�l\�ȕȺ�O�'��xc��[1��C#�Qt�C�ɀ3:a�L�;Q�L��E8	X�	�Q���D�.�T ���Šs��g}���5����R���a�T�/%���!�'��4��
�:�Ɓ��V���ɨ5�ނ9��p��`�n����|~*��c�P�U�B6���C+4ZDJ�%%�������7��7�F0k�{}��w& в�ȨO\t�
s�%דu6p�E�)V�z�ѢH�0����'�L���ßv�S�� V�*�����U)Y��i�m�5��y5���"C�I8�M2ro�Y,���>P"ZO�Y4e�+=�D�
㧇�	��O���	x���P��(��AagL���)D���1T�^�y��rr���B~��#�F������j��)�/�B��ԟZ8�d����:-���028�}�Sc�-5 ���ku��8u@�D_�-6�⡳i���C��]�T�C��ӳ~M��	�C˟0�CD�8<��	#��A�H� �� XE=>�����@�
jh���	,c=�@�u�:���0k��/D�!#��O}|� �g"O�($�M�
0���ҰA������2 2�E���S?��'J��O7>\2�Μ_��]�E�PI�s)۴8�)��H'����DF�N��`w	
+`���h��m��* ��d?�'�d
���3��\��� kd=؉{�K�k���iF�n��0�`)F��Ox\)�L�5�Zt���&�bA�!�i2�=q���'�����،�1�#k�7��{6f�1ji�̆�	Htb)r��ͮA�$��c(ư�t�v4/�=\{A1��z1����~�Ob!�����n�~�YAL	h䁄�*D�T� U"P�J�� �V�H��U���T%2P$ ��D8�~r�O<�韠�Ǖ
|��̻�aBTo.�.9����:2x��ɞH��`�`b�F}H��VU�LT��͏�?d<OnTR!�T_�7��&�u��S���'v&|Qfa��+��41dL�h��KSD\����O�ErDc@'{��))L���t�sq`^�v�3�lL�b@��DGW����Z��y
�a�(Ww&�q�o��i���'.�Mb� �1�ҁaE�F�:M�{���(LK2��dw�T��Oԛ�j���m��1�F��&?��ՃڸL�X��b�3a�j�kq�S�ģ�1��0�w=0��5
�mFx]�Q�ĳR��	�'�0����A!v���rHE=l%�d��L���:XJ�$ቢc09*���Z��t���e% �5ȖZƬ�yѩ��0<�U ��6��0b-ޫ����Vk�+a��X�Z�t�4�����#AP�nެ5���JE)��=��T
L|5�s�'r������Pt~"�DdpE�(1��H�a������@�Ώ���}�D��E��!�>�h���iR ie�,ؔs��F.&�RF|H�L;7��1~Sh�g}r֟� F�BN QtQ����N5�`�$
O��S�NƘe�a�2G�<b��r!k'tld�YR�m��1$nM~��O�a�k	vL��	�(>���1�'\�Ț��/��<hF��3W�� x�j̝�Ɂ�'ø��e�V;7����ú
L!�����vh"}*BK3�����kX	v^&1@��[�<3��,(A�����:sV�S�F^�<1a̍.C��"��C�m��l۔$�X�<����4k��4���A���0�z�<�����M\��ʱnӕg�)#o�q�<�+��ް�:�Ĕ/0�=a��	m�<!E�1{�y���\�U������D^�<�K_�M`���C�Iܮ�+���V�<�',�?R<�����9ό]k���S�<q�/�^%aS��O�b����Vw�<�g�K�0�#�R��%�@L�t�<��Ȗ�FR���4bR�:��a"��x�<iUk�5�h\+�7X:��لiQt�<���	 H��!1��/s����J�z�<����zVii�I�������z�<���b�\� 	�\D��u��o�<y��
�V��dс���Z�)����i�<)��5D��2WO�0MP�i����b�<��j�����Ái����E�'œ]�<yP�!Q� �C�� �$ѓl
W�<)T$�8,���`�hk�!�V�<y���D��S��R�ow>�x�@U�<�����w�]B��B7{0
 B*�x�<q6�+c��X���'lMÐA�n�<�ƪǧUʲ�q�l������n�<�E&%L����U�z�F��m�<V�Ź�2@���E�Da@q�<)���(ۖ�{� ǚ�5i'@�i�<�k�#-E��	t&͘M��-�P�Z�<���NB�@݋��[�L�I"a,�U�<�4�P�j!(�s��(fڜ��GQ�<�d��2>��黃�#�Z���!�P�<9�À,Y�60s.��3��S��CU�<I��C�)�ڵ�vi��Eru���X�<��l&���'Z�s����	n�<A��0*AHi�Ǒ��^�"WA�j�<Q�dYx�tc��z�̽�&�Bg�<�A�d.(Z/ʉ!kF���Z�<�w��N|�����ńM�P���EX�<���� �S��;<�JD����h�<��)T@�p+	�)��q#�e�<�cN�m�0* oC6W�*0���Hd�<�NU�[� ��F�Da��BnX�<Q�g�fMpSÞ%E��2��^�<�&�+ k��@�c�d�du2��Q�<�f�}N���a�P
 ���z���Q�<	�Eڼo�����	B�(����O�<�&��i (�:� 6���c*M�<��eیl�n�p�-N=&�(��p�<���I.V����5&+� ���c�<1A#�g��x�a�B�Ha� e�<����=X�����b��d�`�<���9�>�v�4v�-(UL8�ȓ�DqҤ�rlz���G����m��0�
���o�	x�t�*��$a|��@(Na��(�Q�2�Ȣ�̛{`�D�ȓ��"����|5�l��.[�E�ņȓ;�88�ဒNCЁc�ӧ*|8��ȓf�D;���$Ĩ��Ԟh4�9��S�? Fĺ"�W�:�� ЀQ�NOd���"O
Ij&��=G$�Ii�f�[T|XF"O*x1�]�|g��aҮȄMc(�"OV���H:>@�a��P?���A"O�e�e�=kB�Ѣ+P^'��+�*O<�"0�ݗ�൪��߲�
��'�<�qׄ�91�T��J�0>ꖙ��'1��K���7[N�ICtM��=i�@�'*�pXQo��D�Za@u���X�'�Z��G��U�%�I��T^x�x�'>�����=�p���@�)x&��	�';� U��]36xA�� o>���'�,ܑ� �	(tq�c��i�D(�'E�� � Jm��X�BE�Z�8��'��u�悈2c>��jg�.�z���'�֤[U)��}h` �Jڕ1=h��
�' ��3h� BJ���L2:�� 
�'̖(6�Z�]F���F	�.�D�	�'x����&$��[FhЯ*ܺ�S�'�n ���	�|F~qN�?*h��'�ne�De�W����*m6���'K� �U�ןY ��R߼v&�r�'�>��UM<uW�X�"T0q���Y�'WX�$�/�� Aacŏ3�z��
�'m6  ��	 $9�ʂ�'�T�	�'�B��O��)G�u�M@r����	�'��]���ݎ|�f��VjG�j�� Z	�'�I m���:�#��ُi���'`RDx&���#<�h�G
h�����'8T
�ŝ6�p���J�b�  �'>����H�#,�\@�+��r5��'r�
��M�.`p���F��D��'�����R#ެ16����
�'���q0 �/E�*B��EW�1�'�vTs�����"E�� xk�E�
�'���X���n�.��d�L�h����'m�}��'e۲X8A_ D�8�'�"�lT3{��3�G�(ZZ��G"O��`wJ��f��%��/Q<޽�"Od��2�69u��۵�CBIQ�"O��w��]����煷~� ��"O������"��� Ƈs���ۃ"OPDړE�1�:Y;��A"p���"Ojd ���	
t�q��.P`c�a"O��W��{��y� �M x���"Ob"B��	{Pz���9:���CG"O ���MG'
��a�Q�<�4�P"O�X�A%P���-Ş\��SU"O����$��y\�����]6{��=�"OH�y2�
(Net�XC�� ��A��"O������e�4��5cHIXh�+S"O ��"���|"�G$R��`�"O�Qz���Y�I��O��1)!"O��ె%`r@G�q �� "O��uSk�FUA��V�G��D�R"Ov-RG*P�uvx�����n����V"O� 2&�	it,�ӋS��q��"OJX�����fߐ���ᄂ<v䘈a"OإP����H ����	m��c"O�K�g@�r�`)����4X�=��"O�ʀGG�<Y�ZP�E�mJ4ݒw"O�u�&/ǀ6!���ت|�ر�"O�hBUn/+�t�2��1�8\�"Ox!i�5�0��,I�X�is"O�  ��q/ή{�\���I�d��EC�"O�b�-�F�z�3>�8�H�"O�3b�ҶN�D���Gˊ>�R��"O���C�4NQ�UR�����dɓ"O���!�L�B��)>p$�b3"Od�A�
�{x�̙�2�
첅"O���M��������"O���"��YKVq�D�;S�Q9r"OԈ+֗@[�\�s��<���"Ob�!�HB@V�M;S��3�����'8^Tʴ����y��['o%v8�	�'� �(�
n�>q!�]�7
��'6�e�f�8}N�E�#�D,�":�'p�h9�JXj2�ask�Bq	�'����a��͢D��fY(}��ܻ�'��d�L�ۀLr�BM�{3��1�'Ul�Q�]�2��8I2K����'����lX0����h���`�^�<Q􂂺ox>��b���K&�\y��N]��hO�O��U�b.R���ې��+Gv���'hp)	�hG���������P��'�r	�Beԇز�!��P���
�'(��ۆf�*&��y �aK�\�4�'8��r��R��� �!At��	�'�
��7�H5yw���ꑚ�8�'xD4�K�i�"���mV�Z���'NR%ɱDO�K4t��ܨ9�X�'�Ĭ��� =�$�y�`	�M�
�'�Х*fGZ:3�۳!��14�����'���yN3X(i�6��w6F-k�'��$��䀨�
b�M�/�ȡ�'̌��V�B���"�jB K�'��ͺ#�ϊ#,�!�DU�+b$�'�n=�� �&���A"S�'
�|��'����B����:4mA�j�us�'��!6��)��8Ӥ׵0a���
�'�$Ȃ�Ir��@�ȬS�n}1
�'�B�Aá��.]j��R�ԚM�~ �']�!24�_� 7�=`W�HZ��	�'�d(C�Ƀ�B�����A;�(�`	�'Z(u�K�~K�.>���'���Z��Կ>F��i�Z� ���j�'!�Y�JW�FXd�!V�Nl�P��'��xoJ	W[2�+�M�` ���'���BK�6V��e�?^L�
�'�@�x��-�q�wi�0gX� �
�'���K¼0�F���i��Xj�-
�'����r(� "�N�k�mM0b5x���'�v�c%bì$٬`���C�SI���	�'L6����J���B�X3Wn^l8	�'����&��:|�)�eG%WB���'I���Өة�`�Wޮ�Q�'g��U���`���H�O�����'��	�'��6d*�q�Ȝ0ܖ��	�'��@�u��B��xe�	A	�'v�#1�!k΁r�#��Y�>HR�'r�(&��;�P���-� xVE�
�'	l̓Ԫ����\"�E ��%�	�'���P�#W(~$I������m!	�'�`�[�eO	���B���3)��'(�� /-�Ј�0�r�'UN1��I��m�1�,�LU�'���K�])��Sp%���p)rf����'��{�,�J�(�E��m��#3b)�y
� z�0Ac�tf�X`L�����f"O�@��T�+�B���վg؆�0�"O�P �.N�4 �6D*h���zA"O�@r ϵXN}�IE�>�`u�S"O�\!�,�y�����;N��}S0"O��I �N*a,�m��DM��I��"O�I���h�`�!�j�5��<p@�'Y�$D�0� �V	�W��D�rK�2!���#��2�h�
��3%],x0!��L�'�@) ����{e�����/�!�[>�(@�3�ӵ[]0���+��.�!���Xۘ 8v��!o�<��+ ,Dh!��ƻ=?h�8�#�MaF�pbh�Z�!����r�EfU�옖g�$;�!�<��=����_&�$�v̉{b!�$�7
Jh1õJC�3 �T�`���.5!�� �l�{1&�{,����1�!��;F�č�w�<x�Q�ME�{I!��J4	�f%ꇥ��<X�-�;1!��Ѭ<JL
��P�s��%�
3 !��2�D�R������lY
Oh!�$N�u,92ׂ_S�050�.�O!򄟼c���1�O�ɬ�C#H�D!�H%,��P��1͒�C_��!�DR3 Ȇm'�l�����/_'�Pyr�#-8"�\�R�8��̐�y��E���(2/@a���f"���y"�����d#� �>Gg��f�H(�y�%:Һ�J�ӽ�ǣ)u�1��'�N�����Yaب$*Ϝ �ti2�'��(jƉE�!q2�mϮ�{�B�PK��!���B.��)��� hz�B�M��D��I�1,��bV��$6�|B�I���Xc�̈{҈�9�,B�	�T��(�5LՒKXlc��܄&�B�	O%J��$��58�`��V?~�C䉈��Sb⃛���y�/�/@b�B�I�V�@U q&�#�5�4��_-�C�I5}:B!��/?�X���+#(pC�I.2���� �p5d�� ,C.Z8C�	)6u���s�!'�P�j����C��%s�(Zg�Dwq0�q �3~�C�	���i�{�&����x�C�I�
��4 U���84 AH��8T�C�!Hl1� �\�p��d��I�.��C䉦B 嘰�N6��"�J$(@C�I%z ��E�I��h����k��B�I�[3���2�Sz���Z�dH~z�C�	2.�!v�7D�<rg�J�L��C�	0	��5�%�9�p$���	�-+�C�IMZ4[Ѵ\��I3u�G�U��C��T��jBB_�dŊER�=fC^C����)���t�PY�c�VC�I=���5�.kh�C��K�p7�C�I�n�� ��i\�ق���-)!�$ l��pR�k%�\H���1}]!��

R�(P���>D�`����!�Ĉ%%H`�TQ���p!���1�!���UiL	��
>g+�d���+Bz!���A"�c a�!=6��U&K7\!���=?��dyׁ�v��QT��HE!�D�%I�v�2� <5��`��e�+rR!�DOZ/���I��$�L��B?o9!��,��do�%fOt����=A�!�� Tܩ�	�)�R(����\x�t�"Otm�Tj�$bN�趌�
]z���"O��������
��!V�@�i"O�(W""P< �rE���ѐG"Ob�	#țP�4p@0��"lxp2�"Op���L�����Y����`�"OdSr��8c,ػ��߮I����"Ox[�ψ�8�<�C���+���S"O��Ff�[�(��"Ǜ#�0]�%"O��R�j��4����!Q�4�+�"O�����K�/�!x����Tve� "OR�{�i�^�0�(2GZ�h��1"O��y�.A�+�0����s����"O��@�Q�n��eϛ�8X
�h�"O�WJ��;��`��R�p��{�"ON�`�mN�8��$��,�9���E"O�T��X.e�6������y ��"O��p�čK�<02P�5l�X�"OF��+R�h�FA��O�
dM*�"O�M�d�6#�r�ф��,R� �р"O��h1e\7J8l��� �$�"O|���D��X�1C$Ӧ*�Z=�"OD����
�F���CQl�mw"OJ �g�	(&��q�h #s��p�"O޼A�,�X��lH

5��T
�"O"U۰�B�T2���(�	{�r�c"OP0 ��>U	0����M6�Q9"O@e#"�N:��s!��E�R<1c"O*�3G��mr���↷#3�lH�"OJp�p��P�
�l)��>u���"On8���ѐ(D:�,b�!y5"O"Xq�
C�Ě���*
 ^��%"O��gE_����4)��y&"Ol��L
	�H%�P�:#����"OhA��؞v��`���x2��"OP�*� �_C*�"`�%��"O�1#�� m���kૐ�����"O�-�Ʈ3|"��i�ZlP�"On�Ѥm�#��C�q�����"O�I� ά2	(|J���H���"OP��V+�2U¢@���;�����"Oȍ[���2D`����?��m{�"O�Xi$�N>���6��;<j�"ON�0'���fq�キq �$X�"O�ؠ7Ig�4��UqҞ]˦"Oh��$�Ѵ5��M���&�)y�"OĤ��n\8,�<!7��j�zQD"O���F��Xv\:4��9!V��"O,��P�U0�04G�28��F"Oh���3�Z��Ƃ��,��"O
��4�ڪ0y�$
4��o�ʤ@�"O�a��C��t6H�V�7��� �"O�M�r�M�>�`)3��5�@}��"O@�PtG�`��M0��N� �"\j�"OZ���N�Bgn�:��Mu�8�"O��"��]$�JE���N?r�ԫT"ObC��
4��a�%B ~�T�"O�𛤣̚S֐U��e�2.l�"O�B�L�a�<e��%�b&��"O.股9n�����.�%t�="�"O�)S�)�T��Ǝ�=*LxRu"O�Ah�å^q���mW�

V@ۦ"O�$ɴ#Tk�d�1V��3�.�г"O�h�2�M�\a�5�e+�Q��<8�"O� ���,8Kg`T8gj�;R�R���"O MRԮ
(�ĳDɔ�J���A�"OLqr��Ir��p/M�n��Ph�"O��2PN4V!p%(��O�i�Y�"O�iR�O;A����Ä%�F"O��#�鍡	�Y�G"�J�T�#�"O��YC��i:����"�B����#"O>��b�Q�-B�-[���!~�|�:�"O:|���������L� �+D"O�XG��=p0Ը�a`)<�Dc7"O�˅�Κ5���7i^�ob� "O�ػ�(�;��4#��)p�8h��"O ر�+@%<z���A�;|��
 "Oi���g��-��*[�\_� "O�(
�n
3k�6A���E1�P��"OR�z�K�*O��d��bF�?M�l)�"O�@������:��W���_[�`�"O�(�^�n�2�s���;�l���"OjTb�%��Ѣ�AN�`���"ON�9�ы,��)��lθi+�"Oޔ��gː�숙��N�.�" "O���-��Ie���)uL�2"OH������$i6fO�oH��t"Or��o���qRB�%b'(�	1"O�y)�`�=C�:q���wi��a�"OL�jD�V�@��	(0����2"O�3Ƃ�5�����c��?�U��"Ox��Ȑw�F(�B	�(�9"O"Th5
š%@z�ې��=�@T�P"OR��UT=U���̞/���"OLL��l�;"��9��EA�L��F"OҝpOE78��K<u���d"O4��W�ǀ�:�Y
�"O��#ԃ5���q E�/�VD�"O�0y�^�{��A�A���"�n`�'��*.�搬�J�+B���'�4��,	�K�D�C��!d�<���'ޞ�$DI�r���r�Ѝ`��\:�'Kީ@�I]�j��	��!^ذh�'��xS� G��$s��/ZF*��'�n���愱:�% \'�mS�'��8�#�ע�;T�\>M��'�nũtm�79���� �(\��Q��'��ҵ%۞b�mЃ̛��=��'���#�L��D�#��6�rH�'Y��3�a�~��g q����'���ǃ�<�3�ߣp�zA��'72�BE��x��H
�gK�m-n(��'! ����J�2,�s�_�h4$���'��I��ꍋ([�c醽ao�H�
�':�J��R�?���BT#U*�J�'�1A��,ǔMiF��x�'� ��J�d��g�+(J��
�'ZHp�.L�Z#0�����%�h�X
�'��I��I��wN�AO�6R�š�'�ƌ��@g�����V�R�z���'�Z5SE��& Y�W"V�R�8���']�|Z��2�
 WH�wXt��'d"\/�b�:�O�>"�t�h
�'�*2�O�	�P�R0�=ζ��'� �w�͵VS��bb���|x�'A��U��>~�0)R�7��0i�'lj���Q���1��r���
�'ո$Ӥ�#6��Q�� sZ�@��� lSIġiT��8&Ç�R*�kg"O`q��_b-
(i��E�U����"O����(�?@68��ѴM2԰%"OLu*v������A�oI7DrIb"O����F�=?���Q�ҽ&?����"O�Ͱ��=k^�]iB' �ي�"O ���%�0H���t�J�z$�E�""O�)�B�֦P�Q��K��@0T"O4��c儱OA6\y
�d�$���*O ���$�1�6��j̰-��m��'v<��Q�S>� �M� �6��'�e�VcP���ɒ"��7R���'�H�Ф�V913dpQ2郸
~Z
�'Q
��ݭ.נ��M�	p�ȨZ	�'���2b���AY$��)n-��@	�'+\Uh�FU<w�l�V�=_e��A�'�z��r��'
��cu-@�N��A��'	쐓�^�H��@�㟝?|���
�'�� i�D�f��q�kB
1�HU�
�'�^9�M�O`����8��;�'�@�y��U2#'j�K����byDk�'PX�6�\�1��}�5���V�����'��4�E	M	7�>�Y�!���"�'� e���@x&U��Ĕ-�����'+�'��&	(�����(`���'3`�	�bA�G�Bi:#VS��'������3Hf����C����']0�fm�C�h}#���?�h�k�'w����L0�i��)9۠]��'��a(�M�	k��H���25�tr�' �=���W�^Td�"�oL�J)��'/l�B�B�:V-���y�y��'��I ��ӈ1�<�i��~Z�8��'�ẗ	��) �z�I��d�j�'�N<s��%h}0�!�E��B	p�'d�4�v��hL�c1b�l���'�J\[���/����ؘ$GB�Y�'3�����D�ӓ.��r�`�'+�ER�
	�@/�!�c�J�-~i��'^��z�'E6Y��\)V�V�y��J�'�"�b��1��]ڐ�*h~���'�L�c�?o�&�[0/�8��!"	�']���aU2w�rI{�Jߚ�1"�'�bT�3ㅞ.LDyK'(�P�  ��'�d��$5���g�L6Bn�3�'�����01�([��͋5wF�Z�'Q��B��	fxI�AJ-ni�'r�)z�X2f�ļRĄ�$X�3�'�00aII;cRl�K�.�-�J���'���@"�}Nr��b��u���'�\��&䑒V��"�^���LH
�'a�@IU���h7�Vb�R	�'F��q�� �a���*�ñQ��	0�'m���i��9� Y{v���B��
�'�"�K�+�Sf�d�
�&A����'y� 1��tӪ1��ߥi$(���'[�+�.\�>C��w ��c��Y�'N����/�>�4<��C�*M^���'�ʽ�g���6��` t��*"X��'���PU�
�J�0ٹvBϤ*��%��'�x-ɇK�%�V\06�X&/�`0�'4.@ɓ���%�>����" ��'v����6AT���L��FEY�'��`���V�v춤e�f�,l:��� <EPu��=
�5a��T'�%��"Oj=����F���r�[1
�L�U"O8�7�LG���ՠ� k�&��"O�TZW*?J�h+�H��<-p�"O��T��m����f��f|xr""O(�a��xpT���ϟ� ���%"O�0�6Ξ#@�c��Gg�I�"OzL�p�=g�V�{W`��bK�Ѡ"O�e����'x�*A8�iI�I���0F"O\BT�1�%0�!��J�{"O(Y�MK-�~RP΍%=��D2"O�9�2��7@B���@D�)w]�yJ@"O�$��XY`�ac��KM^���"O���́�t�nu�t!�&5\�p��"OP����-|$D!��D�Vu��"Ov,��R7B�*p@�ǝ	���B"Of !�Qh�@!�i9Z��Y�"O"i��&הAe�p(P�j�%"OF���l��'J�8�!�%L �h "O� ��dI�+�^��b��96 ���"O�	H�T:���0���w!�*O(L��C83�h��amY�E��h)�'5��;@�A>"�Fab�ƕ�N{\i�'�R���X1,��U�@��Fyj��'�
�3�ED	P� y�%МS�]:
�'kl`��e�W�����T�QP����'/v��%��7,0�QH���H��II�''nͫ�᚜Gh�W��P�D9#�'Dq�K=���h�@�/~1H)h�'�����鋀	Fmce�
/J�
|:�'3�q�̖H��i:�nFĲ� �'>�PY��K274�T���!A[`���'J���%���d档RG֢c\�r�'=Fq��/��S���Rd��yֽ��'!��C�@#	W���cE��=�2B�	�'M&�A6ŏ;��{�Gʋ��B�H\	٧A��.�8p �	5K��B��V�N�:��Q#.C�0�%%F�of�B�	�3dP拣h1$Ԃ�N�u �C�I�;RLE�e�9M-�i�1�Z�7p�C�3��`Y @H�i���X=�C�ɘn�T|q�FPQX� 1��Q�RB�I.���Ы�$1���R��ɖI}�C�	.K�x#� ���0/�	%��C�ɦ}�Fy��ƬX0�{@i�x��B�	U3H`y���hX��� �O�jC�I(ȡ����/4LT�q�4iRC�ɯgU��+�j̹z�h���C�C��u\�h�lJ5D��/ibC�I2=��*҇�.gD�3���B�-, �\@�-U��ԥ1��"V��B�ɔe,^��
�-'ض�q�ܸd�B�I�`�E�ElV�J�r�z�Z;H��C�	�W���"�'�-h���?�C�	 Sx�XŅ����s��3ec�C�	/Ѥ@��F�b��q��Kҋ vB�ɵS�.����5�Q
d$��,C䉱,P�eW�4y��c4㐧a��B䉑Q
,}aPN;\!�9Ч�P�0*B��I��Q���ڙP=`eA�D�t\�C�	W��e����|���V�I2c�C�	h���s"�Qz��Щ�aǕ�dC�	 LAZ�OՆ<ʼ�3��Z�^C�I�Ms��z�����1p��ukJC�)� ��K��M�1��'Ң�p�"O��Sb
�$��� ��4li�H�'"O�*�c� M{���Ն%e�EIr"O�1i��
��v�"�χE}�(p�"Ov)��
şYŜݰ礜���"O�1:�I�[�Z����ݲD�H"�"O�e9.0*`���!
'�A¦"O~(�$�ӄ@EN,BD���Ƶ)�"O��[5�[�E��9�0��9U��0*O���A�W2�:i��F�����'h��k�ŉ�U ^	���8���'��qSBϒ�D�z���.F
Da�'��	;�e �]#<�j.6+Fvy�	�'���� �����#��9�,H��'eVA����AFH��Q�O�AH�
�'�<�-��'��q@�!7L4-R�'��1����/#���ŋ�/�!�'���Q�Y�=ΐ1����,�Ή9�'2aA�c׉Ps�ph�m�z�z���'�n��`���yb· �U��'A2��L?"Q.���e��f|	�
�'? D裀ݿ0K�s!�P��9
�'�,5�`�Z�n���"��Zn�-k�'M�쐱lX�,`��Dŀ2K�&��
�'��q�3�l��H��D#H��U�	�'���ڄ5iآa$nՎ?����'�A�a��[1��ӏ��<t>�*�'��@ C�d
�,8S�)��1D��0���!l�� "V��h�!-D���Q�~�<!�ʏ0��4�f8D�8��
o���˥,3�Ʊ)��"D���0F��PY�`�Ǥo�z@�!�?D��kPC�ut�1�R�p�B�
U.!D����g�?~9: Y5j]�?� ���"D�̻���4��Q��+[U��+E%#D�XӲ� ����s�%ٳ�!D����@�rnJ�@$!q
���g#%D�h cTઁ�hC�����i$D�$##IS��4H�f
B2No� ��H$D�Њ��P&��K�(<�tH��=D�x�*C$���6��y��9*)D�PI���8t�ݢa���1F�<�+3D��[�F9[�L�c�۔òxH��$D�d�P����0����% �T��%D�L��#_�O-�,���Jdr�#C,%D�������D�T�'�	4�80�5�8D��@��;#��}�'�H9}�,0�o8D��ՃC$@|�\K"��Q�
���9D�؃�C=?[�.�2�΁Ss�6D� !F��5�������x��� D�X�2\<W-�� �� eJ�)�$+D�İbd[=z�đ�"jmi�9c��6D���L/P1�� ��p��6D�Tr���= �N�0�H:ْ�$3D�X����k�DR�k�Z�`1D����'I�����Jӡ(�$����:D�����$͘��aʍ%x��a K6D��r�`[6c�p#WD̬�vu+�?D� ���I϶l!3�H�uYx؈��;D��*	�) >�(��;7�dlR��7D��� �"8A��gyzP	��'D�ԃs̤��x�����a |, Ɓ D��Y�o,-z�����e|&��9D���!mO��8l���(#
a�� 8D�� ޔ�C-�	eA���H��S�q�!"OHP�B�?#���ђ��-��9p"O���M3� Ȁ%҉&��!�q"O��!���4N�8���U�(p�P"O4\���"�������̌b`"O 0�/�A��)�B*K��ڤ"O��L&l�i�aB�[+�L0�"OFY �Ē1Rb�q� [�%0-�W"O��it�ȠS�L�BB_4Q��p�"O�L �@(;��-� �I�*S���"O
�a�	M�p|.���Ǎ8yCԵ��"O��iV�^��[�U�-�b�"*O��U.�$rJ �R�*:E��
�'�R�!j[��R0�Ƃ�4ԑ�
�'�����(!`v��{�/у/5���	�'m"9�3iP75>�I���5,�H��	�' b��l(o���d ��*���'	\�s%F���4�4<�"�'O�(��N.7��hQg�	���I�"O0e��ܥz0|�P6�1V�r"OB�BtK��p�ՠ���V��"O\�g�2 ����f�ȴ`��-�c"O�ty6�#Zp�QǋF�6%�!"O��"�Gt�r0��X<��H�"O@)���QRoJ|Q6(J�StD��0"OE�D�:_�2���'��%{�ň�"O���7�Ǚ[��m�'�,0�*�{�"O������x����_?�,-+"O2����~��ݙ���7L�8e"O4��A��|I��1v߲w����"O�i�BI�F�
5K4�?*~\�"O�e��y
����x��p�"O��C`�ǋy�r���J6R�*9Y�"Oh�ABJE)s}x�+2��7}x�`�"O6y�4)Ƅ�>\����F��3�"OP�g: Mbh�/�/Vc���U"O��{'Y0Kp�q��Ȓgb� {�"O}��¼dl�@j�,�Yw��t"OС�/
SlR�
㊗@c
{s"O�e�!M�?�9�	�+vG��Q�"OZ�j���3��}귇΋v!R���"Oܬ��lJ�b��UYG,��$$�E"O��k�F�+t	���]g���A"O�3��@�XS�����i��
�"O��C� �rt���H6Jb��ɡ"O$D���8P� �A�6WX2q�"O(��3'N�QQ��D�d:!�E"O��憜4CTʹꧣ��Hf�d��"O2�1�H�dY��f�ŇqR1��"O�!�B�����
Ƙ7k6P"Oj��g$|7>��V
I�=,�*"OL�hR��.�XI��+]�_ɎM
r"OT���+Կ�h��l��"Ol�sqA)�Y��j�&)�2�("OP|i�'O��LiW)W
^{4�!"O��[!��.]���R��wx��t"O��QB��H�IY�J��K���"O�a���ڌ>�
\����*b9�R"On0*� � ���9b!Q�f��!"O��إ�ǵ	n���"z����"O.h�r¾J�����ܪR��@�!*O�`p��@�`�fU��Q7|�4|�'�fhґ���&:�H�Rf�%i�j	�'* �
f�,*�`����d�|9B��� "E{�� s��y3d�D�s�~�3�"O�i��]�v!kGI�'��S�"O��`�$շ<z%h��ҹ?�0Lp"O��@�LS�<��'���8�ʹ
�"ODha���bعE�Pd"O�ɢ��ݺz@
pp��T���;2"Od�����C�^!�d��='܎���"O:`�U!C�*I��ǯ6��h�"OB��D��2�� �D�$E���"Oh|#���<<a6�:�F4�"O�5�"I�i�\8���$���0c"OZ�¥�V�b�R���*A�.n����"O�i��&KZ�15�S�"k40�3"O��Q%��+[�\(�b�<\^��)�"O��ʐ��?B�� ���[uNM�T"O�҆�:6�z5��U�C�,CS"O�@��N1�q�H�'�	�!"O�T!�GUu0��׌� qB�I�"O�����&�&���(�bL�2"O�U���~��G-M�ͮ��"O�heŜ�L�X��NĠ�@�"O�x�k]uĂ�ۗ U-
�:|��"Op)�5��<7M,1����cF"9��"O�tIU�P�QT�p��ᛲ����"O�ĩr"6�	�`�L�J]�"O����~,Hj�o�?�@�Ȣ"O�88�O�|�l=�x�X\2�"Of@s-U/
R`@�JP���"O�`w�Q�����kӪ^��t
�"O��)�f��J*�C��`�e"OZ0KQ�Z`=,�b,4�2`"O��"�O��Xʨ|�P̂�]�2���"O>�䣓?vp�]��
)�M@�"O�P٣��:��U��ʞ�G�Z��"O,h�� ����GOU�]�<�u"OH�3+�-w��[��9��Eh�"O�@:D�Y�Ѓ�P�7��a��"D��р��g݂i�c�·2��!�$D��)��<-�����3l�<)r"�>D�x��i�D�,9���;x`=@I8D����?9��0�l�1qS���7D�T�p'W$|#�-H��[�rH�yt�1D�(:�e72�ݡ�荾b"��뗋0D���I�]#�\�P�)z��}٦)D�����>+�\��� ?;�	ª%D��a6%�R����#|�p��%D��X§G�{�y��k0[Av�36O!D����X�~�V�!��ؽaf=PB*D���Ɔ�s".ف5Ҷ,�J��N-D� ��bՉ�H��(M*~h{D6D��+tf�!y�4X���C JX��f`1D�`
��1Ð�GDE)�&\	�K.D���O�Ac�3�	��V�b A.D�j�$_!3�|��F��c|��x@D-D�Բ�o��X��Ո ��a����*D��A�.ݙ�Y%-�2v|��4O#D��Q@�'�R��7�
4U���4D��u��K�4,a�!ߴ>)R��`>D�
�&ɑ/dD�S@�
�o�@q��G=D��`��1������ڬ@a5D�T�7J	�[�	��7o-��a�@/D��2`(E�^�j�pd��9P��hi��.D���c �q��x
ql��3�N ��:D�L�`�=r���jـ";H�c�4D�� �!A��_���t���=X����"O8H����0:1�$�$J��`���"O$܃RSX0�c2��'=0*�"Ox�SfJE%�+����(U��Q5"O�%(�!� �򑲆�O<9:��8"Oq���5Hc|�a&o�CBD��*O�pw�U#tt��G/����'���ȳ�	1m���cP�[&U��'�̑��RKi:q�E�1p[���'3<X&M#U�j���c��UB�'�8XanS�V�N4I�i��i�d��'��2v�4Y��L"�(��_�^ �
�'~��Q��\���E%i! �@�'��}�1��X��v�ԪO��`Q	�'�x4C�D��7K���� ۞LC"��'*1��c �0����K��q�'�0��p���.=H z%��8�R���'l�+���Lc�!u&]�w@���'y�سQ$�,� �X�dZ?ĭ9�'�&CCcXL}V�X�k(p��
�'�:�HC�6@x`��|2��	�'mD�)�H��5�$����{��(	�'�����9V&P+�._>z$Z�'�����L	���Lb��A
�'�4�r���pF�ܙ���|M(���'�Lu���׵!��c�7 �z|��'װ8�CٵT���A6N�g�\e�'�x̋��o��� �$h�-{�'��(��	<�8��F[�HЪ
�'�`�U��"
Zq�Q�N�e��J�'�5��c��
1�I#�EAu��]
�'�f%�g�E�Y�*�x�>q�bA
�'�*9	%��{x�O@�*$
�'#Ԁ��+�
{����O�1T����'�v�۰�U�|q���f91��MK�'
:�7K��
ަ$��޹�'2��eiJ;^'By�fۚY����'�$�"Ț1�z�ρG1$�q�'�I���[���@��@N����'o�8Jb��h��GA�/4��P*]n�<QW��j; ̸����$�r�yS�P�<aׄ�=v��(�I֬�L4ID#H�<	C� ���k�伜���G�<a���"	p�"c�r��+d�N�<a gV,L��)�bL����Ã��U�<�*nm���L�,���S�[N�<	���z�ei��[�5�h�7F�P�<�5 =;����V+}`�Ͱ� �K�<��JLMÎ���@�%<?�d`6�YH�<ᰯ�6u�Z�K�<�Q�w�SE�<@�бs�0�� g��(�N�C�<a�Ô�XĩvCO'$	��ƌT�<�t��$� �"�ϟ�3���D�O�<��E9gݛ���pq �h7@^S�<�#G�R7�%��(�-�|�r�O�<���υ�Q��	��0���Z0�A�<�k�h�`	Ca]�_�tڦn�s�<�R�2`���s�ُR��M���Io�<�k�WdL�"��!A>��/IF�<!s�g�+�ꋚu|�A �j[B�<�I�XhZ�R��sn��cs�<)�KT�:p��S�k�I�~!�"��f�<0�=��7�PL�椹�BZc�<as�W-d&(�'�Ӌ��%ig�U�<� ����՚+д�btA�6S&q۔"O�A����F@�	6�C�"O��3��$K����aЕC�x1�"O�)� Ͱߔ�HǁV�Dz�"O�!A#GEL��
�!K-����"OH�Ʋ~=��Q�`H 	Z�"O���&�ǚc�^y�FiO�j*Ba��"O2�ȳ�ߴl�h]rr��(f�D�7"ON�q@��)-^���%�:�t�a"O���7g����{p�Ե~��{�"OT��”�8��t��2�N���"O.%2�GC>vH4i�aR�l�`Ԁ$"O`q�H��c��m�/�sj"�c"O�,8%���><�*1n���1B"O��B*y�j�S� %F���+�'��z��5b��R��T�	�'M�� �E�8i �a��@TP)��'@�q�)L6�T�! �*a:�'e�I �gM>}��%��]���]��'8�t�S�L:�\��&��h\n�q�'��t���K1�2�@�T�g����'Ili)��BI�nd2/׺X�r�[�'@̹[�`�%���Z��Z�[���'�Z����,x�Q�+�V�p�S�'ߊh��m�e���P/��C'0���'���w��PW�J�#΀i2�A�'=b8i�h\�:������+N9 �'2�uU�7�!)�
-,�� ��'2�adD�i"^A3 (�t*�'0$�ӆƳn4iz���ت�P�'zZ�PȝF�
�����At���'�T͈��
'A����J��	�\	�'E�!���s�fy�a��<{$��	�'��e[s�;"�Nerp�Ng~����'PT5�����j}����,�_lb,��'L,���I�y�Hy�W��(]��{�'���c��E��{7+��,��u��'<V����Q��}�5G"#X�	��'�j	�v���q�8�D��m!���'�n`��dxhڤ��Y�Z(��'����\�k�D�-`��)b�'B�]������TPe�Ŝo�4A�'u||�$�P�g�|1�A��p�����'�P-��͒CYr�r����o�^� �'A@��gF�D��n�`��@Z�'�H�ծB�i�j�HY^��a	�'��$��mΞc"d���[@���q�'�f�Ԯ1�*)Я �On����'[ s��^�).�MS&�$F*h-��'I$]�5�/	�:�A�D B[�'hP�h'��)}6ݣ��	�2ۼ1��'�$���R/Mm`��!)�)��E�'$�	2Ɣ�>�0T Z<\z��'�`=��kn�f��F��h�����'T�9j^�c^dB֯B�_}ة@�'�n�j�''"��y�f��3$�Y�'i�
�E�-�8�l�4L��"O\�acɘ[��;��ݧ���V"O^� �o�/<pG	I�9�6�y�"O�,��H�w���G&Aq�X�a "O��3S�G!�|�i��Ѩ���"OH�9�	W�F�DD����º�"O^i��KC�qh����Օb�P�"OD\�᧌ d0h-:R�I�=�zY�"O� ���c�Ҭ<�Ҩ��h �EG�p�"O6��g�c���Z$&�3T4~��"O��3p&.M�>tɦ�T%B	�3"O4�@O |�C�
.E�@pV"ON1��d������ҧ��"Oz��,H�P�زI__�@5x1"O􍫡֞(ɴ,R1�ȟrv���"O���'�Ձn�=c#���Zr� "O8I�U�SEE�Mĕl8p`�"O�h%��su��*�Z!iW�IQ"OЙCa��<��r�[Q69��"O �YIv�rW8!��0!�͛�y���
���5�\v��$zpȓ5�yB���h�)���G�sE�4�עF:�y"�>#yn�B0�ϧdr�rwFT5�y��N�B���"ֱ],m`-͚�y�*E�y��vN��_�sF(��yBD�9u}`C�Y@�t��y��+--"�
�N�]�.�[K~C�IX9�c
̳c�
8��	�`�B�	p���B4�K��3Pm3et�B��&�����'Z4혧o�o�|B�	?��Y҃��8@���{�pB�	�X�<y#�_�br8�U��2WŮB�IT��qR���Ah��J[PB�	q� bTG�8h$B�x��:EaB�	 <O�����ZB� 	S�d�B�	5���7G�I��hʐ�Q??r�C䉩8���aG- E�jQ;L��C䉽
7����?�V5V�hC�	66��P�h�>!�F���q�bC�	�nV�%��+F�V�z����>@B�I�X����Am�gʰ�Q��78cJC��(u���JP�>�tl1�%�;a>zB�I�-ބQӐ�P�]�(��e ��o4C�	�`6��xg��=��i��-M�C�I9.��y`]�n0�|9W�R�C�	�Q�x�s�Θ7|���pG�E,o7�B��<�2<@Dɒ�6�5�i��[h�C�ɏB+�eQ��t��i��?A�C�I7Xf����nߺ=�2%g�v��C�^u�$�6d� >�$��j�X/dC��,�&� T���*���`T�_�XC�ɘ8����F	s��TeZ���B��M��0�䪛�u$�t2mD2fV�C�	�#(����,�#.�eP6��0�C�	Xh�����HJǤ���IǢv�\B�I�?8��@�W6)�2�;e��	��C�	��:�K +o!Nyb&��-�JC�I%K����T�[;<)!�ۇCbC�I�f
�y�C*�� �dj(/|#RC�	�>�`���)I�!QO��CGHC䉞��%QG�|٬�8�o��U�FC�Ɋ<vZQX��5ol
�%ǰ&��C䉣.�ؙ+���	3%^�{D-ȵ*�`B�I�F����NH<&��dB�/*xB�ɛ!�d�)Pv
�[�	���pB�	!Q�\�
g��8��׊�$-~�C䉺9W�U��C�i�Ҁ#iU���C�I�"��%h��|1z����"qzC��<54���D��dT#S�S lAPC�I3]%j��ƉE�2��S�ÐZ�>C�	�4�v5��@�"`��1#ĭgg�B䉊i��0�cߢ&����*{OTC�)� �Y�''
���N�*�T�"O�8��ѣ'�4���ω�?��E3"O����nF��X)� �;� �r`"O �B�mB�{��ʚ2��س�*OF8X!D̤t#�%(��K�]���i�'
���	I�(b�`v�.X��Ͱ�'�1�Fݺ:,�j"R5L�h="�'�LL�tE>h�2� EEL'o��@�' $9��E�2h%���d�x�X�'ޔ�[d��7�j�:�*��=(
�'�l���͍�z5�ڐhE���'�X|j&�Mx�\mۧ��/�2l+�'�̩0 HSh�D��p�`�'n2�:"�@�k�LJ֋��,#	�'Id�됏�����P'ç��
	�'*>�iÃ·��)�Q*��\���'�0l�D ����bql@����c�'5�u�Qi&0f� ��"
��'��D���áXAX���)���rę
�',�8Ҏ�?=D�.�#7����	�'L�%�w�պPZ��	��¬����	�'���I@ۚm�.��'�;K�M��'(P󠩆��BI� G�N�<�b�'A� �C�]!|�eq�	E�y3�'R�\�CE%�&,h��&6�6��'v��5C�<�t�{��.��ȓ,_y�3C��?t���@��*C��a��l�<��?*�!�%��$6%��ȓzv�}���>m���f<d4�ȓ&ж$�b�B=(^�A�w�ηcC
8�ȓ0z ���+��vA(��W2x���ȓs�b�#��D<irV�s!�T.��ȓ8� y��k�X(KF�Tb��ȓM�� ��Ȕ7re�B  ����q$e�Diۿ���#���,A���,t*0Nޜn�)5�uΨ�ȓf��pIH9P���W�=����P��uA \Vgxm1�8���ȓ��54
�7��]�t�F�8̇ȓ�-QGL�gd���SB���Y�X ��C�*Ā���d��p�ȓkРX�bĢ���Jκ3Aj��ȓ]��a�d����8��cC8Gb`����4�U�V1X!GH�^�20�ȓ,Q�)cA�_�;q�TP� @y��͇�1,.�+��<�hАR�1@��`��m�~U��HH�R+2Ma�-V,w#ʝ��L��i	*Ċd���f�A�'d�ȓ)"�!*aʁW,@�&O#*�̅ȓI�A1Չ@M��8��@"#7:��=<J�8��V�`��hpq�M�D����>�p{�.�m&�JA���(��O�l�yT�S�>����@�Pąȓk���r-��p���! ���U�B����Pъ�D�y��\�P+J����Y��#
�2_���s�*ȓ��`��h~,�3�.?�t[�jA+?�@I�ȓ	W��0���<5JVS2��'�Pt�ȓo�2����
`�����T%=T���J�Պ��XWh��-�9O�,��M��%�baT�h.�B�!�#�<��ȓ[%jtgX��� �/��H�C�	�x���ɡ
,tB�� ~dPB�I�f���A���#�J(#��pXXB�)� PyXg�S�m���BX;j��	0�"O*]Х�LѮ4����,�T�s"O���H�j`D!�䅯P��yA4"O�I�����"<���	�0��"OMS!�܈Ix`C�!ˆ���"O��TM^���J%��t�5�"O����c�%Ғ*�?k��A��"OV���E�#�4����t\&)zE"O����aӬt2��� DW�Z�"OF��N��=�ΥE�[%d^�y"O�+.�v^d��#K�Q���;�"O6h卖"8��@)�F`��C"O��Rq�½%�F�D�wxxS"ONHx�X!Ou�4zt�J�i�q�F"O64Pa&�|�`(d'
�_��M0R"O��X�#��D�@��4�=׎5�P"O<]��`�7����W�̚`���pa"O�1�_b <3�R2v��q��"O�� �JJ�Q�ڐ�w�
����{U"Oԭ�`I�4M�����:*ird��"O��ӔoBX(J���#?��p��"O�����n�r�K��V9\��"O��X�X�w��i��Ȗ�&訴"OD`� � �����,�R��t"O�Ie#��
��-"k�!���R�"O T��n�
m>�
P��F1�"O<��O�O)�s�)D>b��e�"O��y��GX]AS���-�$8�v"O�Ի#苺_~�����W�z�J,c�"OL�c� ȮR�ĐPc�Z�U�n��"O4Ix��φ�<��fY,_���`�"Ot��`�l�x��A�F�&c�5��"O}��S%����}Q���v"O��#$�J4A�L�R[Uq��"Oj��խZ�Un���`��SV�	�"OJ��Y0m�Vl @��v?x@	w"O��ۤ(��_ht)E�NF�i��"O��ӒBڬp��c�O,q�L��f"O��v*M�:���rWgՉ:��|�%"O*A	��8V{��&КLpz�"O���c��N+ȵcD卽,F~<�"O(�� ��}.܀�vnѲ+�Uّ"O2P�Uo��,J�9�1.0G��`�"O.1�u��D�Dpr�M�� ޠ�"O{d�ӿ%\���Ɖ���p��"O��Q�F6O����A�O�_��q� "Ob�bQǚ�ylT�&J4.尿2�'���K@�O	x��`��I5oT�'��YZ@��[��1�h��^L���
�'_x�ip�W#Hnd0�P�����'� �� �x(���#9�"�"�',H5+ф�F�pZΐ�DXR���'��l+"ω�?�
i�Հ/8��@s�'u2�{p�7P
���n�� �p�<颫����M�C��G($|�'�Qb�<ɠD˾e4�P�dA�g`N 9fHGa�<��虳? ^�K�S�c�$P�x�<Ib��M�t�[�.]�P���c�AI�<Yf�Q&b��XҒn�?+��h��ÞE�<�c
�_�燆!��%+��	V�<��JA.^�h�2oЖ|� ���S�<��"2n `ˆ���Z�j�ÜK�<Y�	�:+F���� 5"�P�jV_�<�` U=m��0Z��
@������X�<� h�ӂ�ķA����� �m"(#�"O☉F��^|p8@ŝbbxrV"O���dB��eLˢ+o��)��"O:��U ��(ږ�Cpe��Y��� "O�bQ"��]I�ꎚ0�8���"O�T��i^�r~8�2���:*b�"OFi�֢̹I�|�5�-A�1"O�����1j��X96 ��/�� �p"O���eY�jQ����o��
�TY�a"O�v&K�|;s̏h�tQ"OغE/F�&��Ȃ�	��	��8C�"O� Q���;:������*�c�"Od�A�Z��]����"0��h�"O�y�qmY�z5`0���=��3V"O��#�@�!�>�� $~��q��"O��BF&8�I@�^923.�3�"O|T{��2�Cg�,"�v5��"O�u�V�Ј�"؂#hW:7t1@"O��yfL?X}6A�Hך~b��"O��p��Ӯ+��	"�#��h�"O��R��� 1q� F�j5n���"O��K"��@!�6�W-q���"Ox���nċ26�i��G/nﲜ8S"Oyh�N�h� !a��/�f�+�"O�+��@ǌ���J+k��I �"O @BTn�H�N�0�̔�V��� e"O1b�O��d��Ɗ�&l��!�q"OV�"hĨ0М���
��@qұr"O<e�#��
W�P���]�lh��p@"O�q�g��wkB��Q�LRL��""OL�zҏT�n�0sCEQ�`J3"O��{�.��f���ᢤ'SmJ�3�"O� ��ַ2��D8S�D8s�h��"O(��\+}�v��&��B�����"O�(Db^�~���@1�lM�v"Ó���ӃOYTU�р�2ky�1+�"Oz�� ̰?,�� �wi�<�W"O�d( 	�W��"#MW�<�Jl��"O��0���"k̞!C�pU0!
""O"t�@e�Z#�`�p��%G!��"O��p`�Q1_&�$o{:�4+ "O�	�U��+T�*C#�6@)v}S"O̬��"��uެL�d��-�I�"O���d�PO�Vi{�e]L���B"O �1$ؒH��J��D�L��"O�V�2�Y��U�x�$��}�!�Ĝ"���o߮X�\�[�C!��6@����EO8$���h�!�;�XM;��7c�h�sԡ�	�!�ě�(��I��6 ��)	� �6�!�$
T��;Ac��s�إKg��~�!���N�P(�'�=�8�e���!�$C�b�x�"�%9�|Q�EADY�!�$�+$�!�3B&Q�����Ԇw�!��
�Yڔ�1 �FB�Y��N�.B�!��1�X�I��}ٖxi�N�z�!�T?;�P���
J�8������!� a{��XC�	C�,�iT&'W!�D�=bT��x�^��;��-o!��W�����hS!R�5rW��8<!�D�B/&\�6�O�"SZ����S��!�$T�\�fM�eL�v@��2a��)�!�d�{�Bj�5~=��jw���!��S?wf�K���, Jx�1$߈�!�� ��k�ES k����0��h��"O���ĕ�t*�z�`ȩ.���"O����
 f���_�_	TP3"O�Qp0oX�c��p��ɐ	Xl�C�"O�1���02�����I�5oWV�Q�"OT�*%O�6{r���B��/����"OڈZ�I0q�eA�bG�'���""O�m0��C�x��݁s�L�$��4X�"On�b�+�#�`UȵL�1�HXs�"Olp�ˊ*zp
$Pq�/_�,�"O��!�O2}�A���ӂQI5"O"� �e��Uv�<H��w�i��"O~�W�L�N����B�ڪ��S"O��kՌč<�^%��#چ5aB���"OU�V��@��_�fU�A"O�\K@i���:��*�.?��e"O�a�槉�(]4I2�JI5+��a"O���1oy�}�5,��W#��r2"O  @BC�O�i��K�
�e�F"O"�rT%�B�����H�0��*�"OB��R(F��D�&aY�A�����"OHJCiW2d�"�9��^}Z�"ONq;�G�-�n����$y��	��"O�0�&�C/� !��ͼm�`�t"O@��E�g�`�����n�� 9�"O���r I�<m���5��b�XV"O�xp�j�AZ��Bad�f��@A"O�|*���G��³��%2�b�"O&0������d����a�"Ob���� z1dp1��B�|H(��P"O�Q�@#�C�Va	�*Ʊ03�pA"O08��ŗn�P�Ï�T.ڠ@a"O�"2(}`��e��v>l��"O�)cVlA�*R�J��3AY�M�F�|��'�l;���2��Q҅J��7&�
�'�Nء�h�.�8��C�:��0	�'���R`�N1���u".o��uq�'�,p` �!�l�c�o��#�'&h{2o�J��nV�~pD�X�"�'j�>�	�P����ߣEh��a_�Q��B�	(p���B,DR�H�nȟ@(�B�ɀ-d�yU˕����J���|I~B�I�_"��1��v7H�JE\�\B�I7h�𰰥[�o�.�d��!�B�I�,�(H�S�D*b��0S� �t��C�:��)I�OC*T��Ă5\��C�	SJ�@�W+��x�A�k�fB�ɡ7�~��bc�&nБp�!�&b�`B� S��AB���g� u@3&�P�C�Ɉ#�6��5�_�5��{�!t��B�	0i�^���@CK\�S�O�2&��?�����3l(�TA��Ul����c!!��
0��|�bK�3#�|Y��βR'!�d��H\,i(��v|B�c�P3h!��ƫ\0�i���}_����1]!�^�<�b���I�}N`�%���!��<����$����Ny�G��(A!�"tGȅ��@<�H}���F�	o���O�� 	�֥�c?������-!��U��1;H�aw�]c�ة��&!�H���Bg$�X��
6u>��"Z���IN�f�Y�Y�UCgF�X�f���{b~es�۪-I!ctc��9AɄ�l��{ ��ʘ�t.�/\!����S�? "}:���P0q�K,��8�S��A��)擓H�f#ײ[O�Yu�^����!�?�y�̏;I�h��'Qw�y$���HO6��Dـ}����䅹k�\��RgJ N�!�D��"mѹ�dԩx�����t�ɩO��kL�D~r.Rp��6BF;.=\<��j���y��!K�:l1B�[Z6+�f�6�~R�'�v)z�@���Z�f��J����'�ޤ3�ǝ�k���z� I�F�0�'��,�@���S��A��*����'��L5��!��DQ�ƞ6\"Y��'{L�PP�nc��AǪ�T5R�'|FꆗgEl�b7ϔ�	'�T��'g(!ᜮ.���-S���'�-��MI�X=^����s��i:�'��9�P��?~+�)5!͢ �l��'u�0�ǼP�Č���H���'��|���l����d� �z��s�'ɦԫ���&^�j4����z�m �'Q�����M��'�{��%��'N�����P�*����!1nvֵx�'��A��7R�����+��K8���'XD���'�? �d/�a�ES�'���sf�M;%VX�CC��X�
�'�FIyR�Qz� 9A��\� b�\�	�'Ǟ����ք>�ֱ���Y | ə	�'v�3֪��X��(�]��))	�'�,E�S$>����Yi�D��'�LQ�c���0,bAhB��S��\��'�D[�MF=Im�!�"�R&@�
�'U*l�sc����U�y$�a"O����f�J`P��ԦNtF@�`"O�$7�و���JP�_Jo��is"O,14�	6U*zu;�� mVv�2""O��� �wY�x��#@ZC���@"Ofъ'�J,�f(��OկG���6"OL�+D�J>'�@��ĕ04\\� "OXa1U� �*���?ʎ)�0"O���	��P�8v�E5/er�P"O���1DT�n�D5���Ų(�Lp��"O�9�gԷ{���2�P�<�p,�"Oz��	��yzhL��O�4"�"OL �$#�>Nn|��=���q�"OZ�1f���0ӈ(�)Wa����"O~2��=4�(u��]��H""O�h�Z�3�G�>ƽk��[9U!�ē5G�8�P��=�����R�	D!�$�v��m���
I ��x�I	2I�!����l���)�mZ1j�7�!�Đ�DR��#%�Ʉ���f"��A!!�$��6ܪ=a�c�%4�s�`�	!�T� X�X�kF%\m���  �]T!�d�-���A�\��Y2q�S�^!��U��0��F� �n�3W�|@!�DȾW�e0 �̠F�\ēE٠E,!�ɰC�`!��A=@���*@�_!��ʡ;��u���XQ�\D(�+��D�!�d)io���g���P�JY�I�!�d�`�*�%fįŅ�8��+ "Ot�V�[l�"7ĝ�",���"O@�C����z�*5DɅ!�ah�"O�5v�G�;��)��:?�t	2"O���fJ7Ŋ�������"O�s�O��w~�]aF��R�@,��"O� B���Ԛ)��ɕd�if��"OpIu�]�wN�`�I�P�ི�"O��AU K�@�"U��뙐��}g"O0�%�N|Ƅۅ+�9 ���А"OA��՞iUص;�_mhb$k�"O^��u�ƙ<:MR�č�;��j"O�K#g�cʝ��F�7�Mc"O������{5�QA �T'5�`"ON��mѠMw$�h�,i>D�"O��)cL�n欲���0l�ܫ�"OP�� >X���b	�]�lD��"O��8��I�h��a�@��H�"O�ɠ Ǘ6�y��""��4�"O���&��	��h�2F�b����"O�y�w-5����eW�2]��"O^��Ed[bJ�5�g�\�"}���"O��y���!N�T�H`G���1�""O$��R�
xk*�"E	���e"O�$KaBǙV Dȹ���&I.�R�"O|mQv�^�L}(PP�h�
~�*�
�"O&��u��5*q�r��V��F�2f"O�8��LZ�v�:���sȈ�(g"O"ܚq�ó��y:C�֐;��)	�"O���aÂ'RAԴh��\�ru�E��"O��ZU�ރ	�Y;a��GB�"O5�V�٠8�|=a�ω�~d]H�"OJy@񪖩F��ر�/ǰ��9�t"O���
�Es����m�.+^R@"OL�Q����}X��*�gҝb(��"Ol��fBݰ6B�y!�DsY*p90"O���+�l��借�&@$ T"O��Q3�I�K��!�OU(Q^��"O$)�fA�8�`��� ��M^���t"O�@���g����!B\+��`�4"OD�S��� �xM�堎�`�Q�1"O�������D(�0ǹws��"O�݃BFB�i��P�@�ʀPp*��Q"O�� �C�$�\|`$dڨW����!"O�H ��Wh&h0�Y�N��9zd"O�8q�Y{�c�l�8F� �"ON�3m\ &�hV��U��A+�"Ob�BwdW�(��ܰ���b(��"O�a,V�A�쵫�f�'@�d��"OA`�L�xV	��g:�F=�"O�!Z�&�>�P �%F�;R�^ݒ"O䌘�/�7Je<@��e�|y��"O�@��|����MMUDl��"O� 
��|��壶�L;6�l�"O"L�%�-(��YrէT�8��͡�"O�5�dK�!e��p�F��E�ȸJ�"O��0A!�/Z$F�.!�$H�1"OZ� �R��*�rEN˥�f��#"Obi`.�%l�	�pL�5MxxȚ�"OФ��e��(�sE
�< 9�7"O΅��
�)ֆ�1��vT�-��"O�5���C ��"��C&]�<h���_d&(x��'�2ãnP�p��
եHiV�*	�'r.�A�+��9&Zk䨎"o�~0�	�'��!�G��>a���⋇o_pS	�'cJh�W#T5a?+EO��9��'5 ׭����D\�r����'���˴.ҒA��j��՟m�d$��'�|�9C���h`K�+0�e��'��:�ǜ67�MK�%�S������  �y��f�$|�����-D^�"Op��K��j��ɐ�5b�"O8p��D�C��T�A��'H�TP�!"O�	A��>7�M�C�IQu���"O�(PbK�z{؁˴�֞S��P�"O=�oF!m�!�5"��a��MkV"ON�R�O�ȩB�O[r¶��`"OjlѠ"Q0J�����.��v���p�"O"}��G�,2�r`��Z�,jN�2"O�I���>%��X�" �i�r-d"Oh��U"L?nf�� Q�7Ѻ�c�"OL)��/թ<�>X��V���2$"O�h	FݬN^����%�!t"OF��ċ�X���J�&=겤��"O~���,�!609:��M.c�|h�"O�l� �Q�����%:(hj�"Ov%k��'6�0�RVL�4��C�"O��WG�	q�Z}h���4�|�k�"O����Ռ<c̈y ##��M��"O�����ǨkF�h����X��`"O�-�j����]b�!$V:`EhC"O�UA�
%����� #�DYW"O�pyŊH�&�h��7���"O��"R�}(���+o+z�yq�O��`�� 7-ZqS��/,O���E'��1�����!�Rl
p�'k�O&d���e�-��T��K!r ��)&��/)E^�z�O�\�A	\�-��	�ň֫>�h��@��/.�3�$r���@����E���C�,EzR\���Γ+y8E��N�lu���Le�pP��6\����OV����x�$	2qp��^�O]��/3��4Xm�)�0�ʳl3]s�B䉩ʂ]�$샏X`�4k���0
�
�LؔN�4�e�o� Rg���F G}"ER�V��q�1i�2.�|1	��<�)V2,�h#Q�ȊU(Y�ھI�5����!��`�Mݥ|��������0?)���+[� �b��O�H�8��t�	�����!b]�jB��A�� T !��ɟ)&��?N�V1#f�W�(2�A�K�2e��C�I(�ub Ԯ%����&���|��� \%2	R�r/�n5����+hܧ�p`�;�,*�g٪�$�S�k�!T�
�*�
O�sB�9�`��CBȮf��`�v�O"!��3��֩=-��"�jN$nO�LB��8�n#=�4CL8Ql>� ��+_.hi���O8�����	q.�\�0嘴46�@�nr��%�R��J��0���r�bS*^Y�T5��kX����"��	���Ƣ�x�<U���!}�ͅ�'��e��t�Hȋ���F�VhkR]�k��ӎ>���X�6ĆY𡋠�B�	�?�0����#�~�I���8c�1�C@ΑN���Qb��A@|�3F�ޱ��EHr�~ޭ�pk�'|�����!�ɀl=�O0$S�"��R4B ��+�y��G
���!R�(��Y���r�4Kr��� O�v�^,z��_�.�M��ym��-GX�P*;;�P�c\��hO�M��W�6�:�.>4+��pw&�7gF�4ѧ� d^� ���
)��#���!u��f�8,��­����<����J�z�14�U�#U���� (�\x��)�A7R52E�D�!�B)ĄM�b�a��� S����!*�V|�� �+�rݚS>n�`u�G,4^����_�j�C�#M��<�M@�j
����G?^	��(K�g�<J��0]�`�8t�T"M�� !�� "lϻm���Q�"^�i�������	�n��� ���K[t�P�F��y lO8Hm�T�����fִ$�����TƉ�o2a�0�:B����;Na�|�'[P5˂���99(hE$}�Л���Oxv��*t><B ��M6����
)cS�(� 댦3:fL�u݀	��P��� ��|��Z�-�/� W��D~�,�FJ�'N��JYI�Ћ_�z�P�$�z��yѡnw���ULV�CAԴ��N��@My�'�V��<aK@E��MQ�/����H�ז���'ئ��cD<��`�!�&��R�m��:OZ��� Gd�/��Eд��;��=$�"��b\c���x`� 5j�f�+��دH�@x)��3lO��E��+�D�1����<TP�cw�-,H���g����<l("�u�!�c^�x�T���
�&8f08�A��+3ꁨm��\��M	q�R �e�)�%�%�6��Mr�Ս�1+�M!��/��t����_�� H���qx��*�&2 �mc��K8be9�g
�&g�k��е�p��CV�' -Kn:�Ya�D�W`J]`Eb�`��Г�|^�RUfT'1sf�̓9 �y!G��Sj\i��1aG>Up�'+K����5A^ ��䒄}d����#n�氛4"�� L��O7>)ʖ͎;H#Lݨ�o�x�Lk�#�k���ۄB���d�ׁ�59�7�� �ͰE�̫2�*���>#D�P��'���Io�����˛�1���B��AU1�y��%��=R�lrS��/C����_�Y��sɧ5���b�lV7�a���ɰ?V��R ���i���x<�Pà�&�O�8p�	��Ot,"��P Jc�)���d�@��� !k(|�u�R�v�hbrIݖbd�XJ��B7Y� ���'H�#��Ii6F�$h.�>3ČPfaY����Dg��0gJ��E��@�ɨ�K@8Kv�0s�č TnmA4A�����G�4iR��T �#l<�i���6OET���fłN,���'(r���/�;�LPSFGܤ�|�"�bW(��|�J�7`~�i�a
G)q.|��WO
�:�H`�g�&�v�:�;~�VU�Hzh)����P b�x#l���ѢW���F�K Qfzͳda�/
���w�1mS�0FW�I���`��������G�B\���_����'y��	0,�;2�����c6sq|�
gg�L��9" ظ��':B��cΨIf�$,0�YC��C��?�Co�Kc�0�S��4v�8<���< bC���|��͖�_N���#�� 4�Ԑ
�J'x�lA�d�N�'x�jE٥�>#���2K�"(�L=HS��P�����͈�,�!�$�V�؁��
�t���L��9xE�I:���P+י)޼e�l]�U�ԙ���_�x�=�A��J.�]� �V2+P�&�6�O�ͣ�G~�8��V'R�*%�E
����L���y��nu$M�҂�$��ov,]��ḑo�:Hص�? T��Y�9o���g��!3Ƿ�����7e
�Âi�]k� ��>� `ߗO,v���ɭ����;>:<��5g�#<YƦM�^ړO���:X��ƛW.6$H��7"����j��!�D-���	�sg0��3J��E��̀��H��m�b�@���
��b�L�zQŸ6�]
�y��S�W� �@B�%$̬��ə?�M���S&F x�<���Lt�>ѷ��ʈ�(��A|�����v�<I��E����PuKſS�䙹��z}��F+X-���ۓWD2$(�통�����2�>���I�3�6�k����P�F,p4d�Ĕ�E�����f�H�� ��:�4�%J�;'����$�XId�D ��s3d��>h�ȓ3,{�$�*\���Lg�.a�ȓr���IY�=�|���M�A@�E��P]JTs��Z�����\� [���ȓhaN���.D-8q`!3�9d�p��m
|�X��.+�9�$�EL+��ȓdK
�Xl����@�F)��	��vfHX`p@?xG����i%MX���ȓ!�I��a�6�t�Cfk�#fĈ�ȓm�
UeB�fLP�ۧ��k�(�ȓ�`ѐ���S��+�e��]�`	���0s��L�6[N=sׇ֬P�dY��C��P�!�$d�܂1D�<.6訇ȓ�I;Q�ɬbK>(ac+T8���':BM	v�X�0!v��4"�/����ȓ��$S��P%=4��g�E�J�z$�ȓc�~�� �4ydĠB��rm�����I�5AQ>�z4�.Հa�Y��F R�.�F�$-�&
R�C䉯O�\� G�Ts�+�]��C�(�J�R��c�a��� rTB�ɗnn���ˆ�V��C&�M�B�O:�YKs�τ��1a�($��54v�H�?E�$�]!f ʴ�#K۴9�e;��P��y���@��l�v�X7��Pf�yr�K!<� �(
� ��*P��0�yrkX:^\m�åӟ���hE�U�yBJ@�PDr�� �M�|�����9�y�h�3)Ԩ�d��9]��)��&�y�Û6J�,��OU.*:z�pC�M��y�	D�K�ڼ�����)tf���%_8�y�FA�����&*G%(��M�����y�̙�.�08��ݾ�c�j�(�y��H�5ɨ) B�7�%�6�؛�y�c��~��H�dJ�~EĘ�� �>�yb��/e2V���m^H8R�D��y
� �p��7W~t:��i�
���"O�l�$[0=���Q�˖.�R�"Ol�r�
�(A�tyv�
�XF���"OF�S�yH��[7#��uN�ys7"OpT�g��5	YZ�r2��SV�!("O�a�D�Q��;o �u�0"O.$���_r�B���LO�o�5�W"O*�i��"] ��!M#.�1�U"O��p� �2"�x��D=R,��3"O�����E2L?��������1��"O�س�CAUP|�3�|s�	�D"OJ5K�֝3n���'5j�H�"O   Q�R�b����ab��}͛$"O|%x��m`(ru!��X���"O�YV!�TZ0yt*#I1�]�"OdU[�<�zxCi��Ѩy��"Ollsr�.@�nL£nAV�4�p`"O����HZȪU/�;&ô��"O���q��7./� �1���<�b�p"O��!��ߣ?b���k6ҭk&"Or���'Z�~��-V:���1�"O<�2'�\�|(��ߏR6���"O��:}� ��
�%D����"O�57#$qf�@T�]�DL:(�"O\�k��1,��Ppp I!$ƌT"O�t3��N�h6��1�D�	���:�"OQ��80�|J7DN�:���"O�:��n�����R�x��Q"O���q�G�Z+&�Q)t��i"Oj�{d�����B�C�20��0�"OR��􎋶�*$�g)M$8e��"O|8u�ĉv����S+E,��i�"Oh�l�5@���"Mޡ�l��s"O���o 6�B]rmS/)#����"O,��J 1b��½�0�E�T�<�E%�����E��5�*0{�C�R�<�vc�2h�c��Ѷ�*���Q�<�%��ۈ�2�N�T�	"&dHy�<��(�;�i�$i�fNH�<񠢟�1r���O* �"�H��I�<��	I�L7*�p��)A�tu��UJ�<�Ɯ�kʪ]���� d���y�<�O;P�C���'-G��+D�Wm�<�3��4� �[Dҡ����b�d�<�g-�Ph�kp�ן$�R��j^f�<�U�Q�n�*�:7jR�j�P!A��X~�<i�(�V��F��̀ӉQf�<Y���4���:�#?p�|��2̏]�<A�*�C�h���lQ�SE�����G�<	P�A���)rl�
n���RW�<��$#5��
cY[\D�t�f�<���E/\�]�č���e��u�<a�jTOBĵ�p왐rv���
�J�<A6&����p1
�+ �.�jD�<�o��XH��B4AC��D�<�v��/.����`��\b�}��ŗE�<��ʰ\�쌒wd��P�(�����_�<�di��K˸(��J�4���q�/�V�<ɦB�2�]+���8�
�BD�_�<�"�0���#�L<J4��A�Z�<��(C�fo���� h����RcP�<	�g�/߀���X=\�h��w�Xt�<�"؄^醩k�����U� u�<a�/����İ�%7v&��$!�l�<� @�hS$*M���뀌Te�r�"Od�H7�?x&ڰ�%H�;d�$���"OR�3�l�-�%BӨS<u��l�"O�X�Fe	�/���gɴe�j��"O��ZG�,,��=J��Ej���Bd"O$���'2��$�b抯6d|���"O��)�Z8B��`+���7����"O��w�KH��P�E�r0��9�"Ox�k�����9 �"Rt�Yv"O�����~d��jݗWf�B"O�]Bw#**,��$�سa*��KR"O�<�c��.�j�R�_r2�U"O(��˒�,0E۷n�!�BĢ"O�U�%��	p85����h��<;r"O<YBF3K���s����VP@"Od���˯\r�h ��6R	��"�"O�5ȣƂ:g�h0��E�xl���4"O�hQ��/|9�	p�B6j��*�"O$�@�$T들��dx���a"Ob�!�n
W���P`L���=Xs"Of����~-R�:a���ً""OVu�bI<%!�$k� F��:�"O��R��B����J���L��T"O�QJB�Z�dĨd�P�0^0� ��"O�P ط	q�l�GÉ"2ft�2"O���+�',�ʴ��i�@��"O�T�&/�3��=r�W�&P晒3"OVY2Sk�pߒ@2B�+,@Be90"O�12���}W.�@E�**ry1�"Oإ�q������b�	U�e;�"O��:�%�!�����!P�	���"O�u ��J7Ix4( �}�LS"Oڽ���B5�P4F<wK�H�f"O&xAMzƈ�Qt�Ğo
 �Y�"OL���6��B�mшhԻ�"O��ZՈ��/4��F�c,9!p"O"�2co�8�@*����{a0�"O�8�"$м(&�,�Ӄ�[��$�0"Oڈ$��!6 �[FA�E���"O@�aEHT=T���룦��KM��K"O���a�ODk�Q��FC�
���"O�����@�s�T�FD�&W,`{�"O ���.x���EJ�`I�0"O�dZEo��iˤ4	���p����"O|Yٕ��'/|��΁0K��)6"O��0A�%s�f���Q Q}�,A�"OB����c�PD����QQ,�"O��i�K�1)�T����B\T�"a"O\������. ŧ؟mG��)�"O�Y!R"�f�Fi5��=4��"O0(���$H�pH��_����"O�]�#�:<��t��,O�h`�"O��`��T�n��Sb�L�B��"O6٤�� S��AE���'=f=0"O&����PX��Z�j�#q��<b�"O���=�i� �S�2j��"OԡOŔK'^@�!f	!B���"Ob}���T>3�� ��Ɋ,�h�c"O����	M/&<�f:t�>T"O�=����ERz��CEM�6��U�"O܀0F���X`�QI<����"O�0#Y98�������#"O$pᇪX�DZ�MI�&�g�bQX�"O�t�J\�o���ㄜ7o����"O�  Ц��3=?�t+��q��j�"O&�b�iǍp��T�1t��ɑ"O���eC�� QB(�dx�"O���!͠~�y0�	A�8�vE��"O��+B�+�LDòN�'���q�"O&�K�	ϩ`���#�/�8�"O.�(b��"|� ���6@��W"O�A���V2��(1蝖C;��Q�"O���C	L�"M3�J�d*�P�"O@��ץ*̸��U��|��	7"ODS����=HzPrRc�d���6"O&��+�~����XX��"O��֦�d㮡
�߲L%*m�!"O��R-W�o	�u�$c�u�~�Q"O����QRA�uZ���遂"O�d��̵qO^$�֤(E����a"O6��PI4'������;M�"�K�"O$�K3NL+~�Ȉ+�,��h�"O���풹]�@�a0A�>N:�3�"O0)�R�F�R�	�j�D",Xj�"O�^ʐ	�(��g�1X�AD��!��8���A�\�Y^Ƅ0q�g�!�d2	k��X�ND�~�`%���!)�!��r����H�/!���U�ķ?�!�d�C�Ze"cK�3|v@��d�̈́8�!�d)9K|YI��R5{䌂#l��!�$G�SVH�C��ivkXBt!���%�q�UT2iG�I1cXO!�d��*�E��M͑9��3�#TA!��\����P�@F?�xS�R	D7!�dM�
vtR2 �	g'0$y��1�!�ҋ>�h0@A�1��%�
! �!�$
.-�m؀h�?CTH�-y!�%n���b���JPT�i��Ӫ]!�DY�^{&�: �J����K�!�X�)|*�`6�T�Y�Ƽ�EԷ.�!�E.[Df�`��r�<����)t`!�$&`̄ZS@�6[u���jчS�!��ă9p�@5`%5��1H��!�L.3��Q�0q��%؄ag!�d�u�Xܩ6`��Ien%cW#�Bm!�DԀQ�����%|~hr�c��f#!�䃪X�(�g�ξ�t���,!򄓆���#�ʝ�@��%z%`�6	!�d )�L�%��7i�	�R�ø=�!�K�5�e�
��)�S�'!����*���2��|���S6u���ȓ3����Cm�\�(�9�DY0b��-�ȓ�f�AB�)H}V1IP��2e/���FIޕ�t��'ay����	3�8��'K�����TW|ɠR K4	$^��ȓ"�V�5gӕO ��F
aa���$� #�26p0`3���xj�(��v��is�f��>�X��;���ȓa�,Tӣ#B,i�A�	�
3�|���NL*HY1`H+%��"���Ն�/B���/Ȱ*¸P!�Ș�)�ꥆ� �h��gbC���e$1!��ȓX�d`�FE�q2�,
E�T Rղ���8tF�26F=�l��3��,��<i�Ub�%֖,�A��ܟ9Р��ȓJ6�cL؟Kc4�D��1�⌆ȓ��4�۶1��)9E�(tFl �ȓq���@�F�E����C�|��S�? �]�c�ˣE�0ق�\�,���"O��*U��M
V�g@�k�e�"O� �s��lP�{� #yi>���"O�s����&\��O�T:��"O¬zT A/\!A�臁TCn���"O�L�D�0�����AN�{7��"O�����LqLm9����Y8Ĭq�"OĴ0���y�-6() F졓�"O��)��$nJk�Y%x2ސɃ"O:�A�ѝR���H10 �xg"OT�m
�F$� ��<4�<�"O�Jp�`d�;1+�6|:�	5"O���F�D�W��y�$ˍ��k�"O�qQD��t����@&|>��"O�X�b�P�N�z�ʑ,��p۱"O]Q"��	ވ8ځg�,M���t"O� �K�LX�Iyg�*s��"O< K�}�`�xS!��b��Ia�"O��y�*J�F�J�A�*�)KA"O�=���7Na��y��p>	�Q"O����Q�%���(� � �y2&K) f��H�a@=mF����ۻ�yr	׽Ka�� �Վb��A2؜�y��7h�LA嬖;Z/,�r��y�,�6��h�䆋V��l�A�O��y�U�KN����ŉ}9���)�y2L%	���y�2�����=�y"�[�ut�ݺb��!q��a�A%N;�y��V�M��5�W�Q-h5$��pO�yC<g�|LQ�-�,;��u	0(N��yҭ߮\T4�H����:u��w
K�y�f�,�p�g�Ĉ�����Py��S�x�̨�6!;ID�+��GV�<qpa�~78� �K7��C'�Q�<����p����� ���s�(R�<I�(�]�N�z1 �}<x=��I�d�<	��?pFR�ZB,�'�=9��NO�<1��@��h!0�RR��x�H�<�0�J�BD�DXl6�`�n�H�<駬K!�@�
�h�?[�:m���]N�<����"wi�L���?*l�[4�m�<���]?�,�ॎ�>R��#�R�<�P�\S����rj�'�<�Is*H`�<����_�Q� �8D�ysLX�<�0J��?�Y�^$c"Ly�s�<!W��`Z`�� ��&�܀��Q�<����HN�]�Gl
K�^�y�d�I�<�R��>
���sp?$C��N�<�d���P�P�+��Zs��Y�Wo�I�<1D�ŤԪ):�A-��l�UE�<��E�1B
�ڐcP"��k��Z�<��B�;sg<��פ�;���@W�<��
�O`Ld�w��>�8��j�<)P�����Uk>m��Z"ȖC�<1U�Y;K �L;�A��A�����W�<�i�6J����p(9��#EX�<!���>����2	�A�lQ�ӥ�T�<���#
ZF�:��������2�^Q�<���M.R�m҃Ꭾr@��r桍Q�<Y��2j��D_ryҊ�N�<15L�I���4���|m^��`�E�<	��\�v�����JK����{0Ɉ|�<�'���Faԝb�$��o�Nhӡ@|�<!u���t�b�N��V���ظUH�����cx������<�  aDmؽg��ܳ�e[�����|�E���Oq�t�yW-�s�Z�31ԍ%��H��FGw���0��ջ2B�P�M�����Q�U�� �t� ֢,��JX�ĸuY��I�IF��q�'����ᓖ���T�^�H���FO�V�m�����N����l��%cE@:���
v��0 �p��^�b������+`����	�WZ�a!��\��a�tA�erZ�3�b�t�jl)��tF7muGP�)��-��i����,G��Q?`h�e@��Fp�p!�C��^���iI<���iF�����~��O�r��q��`I�r���Xǒբ�'�[��<Yr�.6�,�e�jxP)��'`q�5�%o[1Ԍr���	N���[��x c��G�*��$\N>q��Cư����t�2`��/HN\�� DL;z�EAWC�|����i��vv�a��(��.���a
�FIy¾i�l5B��˅75tA���a��o�)p�L���	uh���"H�E�g�$9o��H@�֍)��Q�':���c�Mك"C>Ac� c:8�soȺ6ޖ9l��h���n�OQ>�u'��K"��g��9	��E���dbM?�xr�N��]�%�A�A�v�x���y� � I��=��K�;�H�2��-�yҩ�o���*a�M�g`���p��&�y"cK�W��˗*�6\2�"�� �y�
"3b8*�#_�YR�I�IA��y�g]
�4I����P�N4���
)�y�k�(֑��2Y��ԫg!� �y���1a��ې A�R޺���
�yrFD�ǞQ��.�MX��X�� �yi��;idH[�� KH��6�_)�y�`�24,��+���9;�.�k1E���yr�P�sXy"�
M�9Z(���bK��y"���R8�Ce2ئ�@ *C'�yR#��[�l��0�L�.V����+�y2�'!���P揌4\�|�&cޱ�y"�(��⦇N<,��9fή�yr/ɐmhh�O��*!L<�_��y�'ݑII�P��$�rXJBa��y���(FHzv�"d�S%���y��^Pl�Qp4X�[a`2`1�y� �SVa��J!S�^q����I�<�W�
�*�x��"W�
���N�<�w��nZX�t�E1�p����A�<�C$[@ǒ�9f�&�����^I�<�k��V�xm  �$pT��(HH�<�LŹP�<q3G��L�T�5@DA�<��ȅ8z7�� AQ��0��D�<�v�>��£@�3��$��@�<�A
�:JtF1��I~�$,�A�<���T�4�p{��r��� �^T�<�g*����� ST:=!GI'D�`��#Q��2$֯R"�0��8D�LY���`h4$�3'Q-L���#$b;D�0˕�]&'t:t*����dD�9��,D�\k"O�Q��ak��
#m,�� b.D��0�T2�Lm��^I�l�" 1D��YS�U=*r�y�R$̋.��Z��-D�tQ��­`�2D埦��xK`�1D�̉�C&r�H "f�m�xpC��#D��yR.��3�y�4K� q^
�8�7D�|�D_�etȹ��\t0�]3�$*D��1JA�qJn0@bQX|a�f3D����+ə+g.����:�n�p�k.D�4�S�Nnt�D"T�Z"4a8���!+D� �c�u2�c&D̏�&�
� -D��z�?�4��-Q���C�)D����jUE��x!*^)�ڸa�d'D�XH�B�7q�]c�-"GK�l�'�&D�$���Q8?��T�R0�i�ed'D��$���&��d��O������"D�� ���O��Z!�L���I�t��"O� I�蛶r8ndj��?)���"O@��#�ȊC�m��b	���"Onp)��LE�����A�̰�"O�� "a�,���è��xt�T"O�%�D�
�\����!�R��2"O#�H/{VXz4��]�%��"O؄!S����0A�K~xt��"O�@Ӄ��9��Y��D[�'J4�1�"OTcClX���1�T��)X�"O��Ptb�u��,�7��-w��sq"O�h��NC�,8��蘝-�i"Opաsh��!���cgN�&���!"O�� L�dl�|a�*Fм]c�"O�%I�Ȕ� ~�@�5��j�a�"Ob�Ig��Sk�q�dE�.�	ic"O�]��H�m�uI�A�	��x�V"Or�H$k�cQz9�%���u�B�AR"O�5�TiR�Xq蝻�Iϼm��Ф"O��i�郓*����ӄk	RqK�"O@IH�IS�P#JL�ą�/��"O����H�;j�q �dN�e����"O���#aP����EF! İZC"O�"g 2%�A���@�"O\�
�C�[>��� �І�2e(�"O�Yef�#n�Ѷh��wT���"O�e��S�aufq�M��eR���"O�j� <Lp�)���<'M�xx�"OȔʐ":-,XU�W%YB�$ �"O2�X��\2c��yc�5J8�,9&"O.c��U������Ĵ��P"O�L[��.dk�X"v��0�P�"OD�kX]�n����RX�"Oܔ��ፏ���`ťS*.hڕ��"O�lqf$A�q���%��}�<""OЉ�MC?g�v��GJ�k;��d"O"`i`g��$��z��+} (�I"OV�CcP�a��C�����lx�"O��!n�i�9"��V�v�Ь9�"O�I(s!�z�F�f`W�+�z��"O>1�"�E�_٩��7�� �"OR��a�=X�qx���,2�� b"O�HC#�S�an�H�Q���e����"O0l��n؆+��PQ׫/�9��"O�l�S�V�5Q�r��R2��d��"O@�0v(K�{�j��3AO�;�8�s"O:��%�ZP��{vʈ.@��"O4�R񤅢Z���0�)����Xs"O�0�ҩ^;uRJ���m���""O��׌B��>H�f�]":���� "ONa��7�(� ��#N6A�"Obez"@��l���h��8HH<��u"O�lAQcX�#��tт
׆=tua�"O<l*h�<'`�[�jA!d��Y"O����e�b9 ����A�k�"OL�RL2m�,y���\�
�I�"O��B#]%U���&ҦV�~QR�"O���@`EU0�cpn����"O��p�O�|.͒ @��?�8I0"OFv��L���o 7Qnn��"O�x;�(�s��q��H�9kX��"O� Q�\���!�h��h�@�"O�Ԃb��6K�������`_��"OZ0E�W�aK�ebF� TL��P"O� @��ҬW$�����4�m�"O���k�>#�����-A&�ဦ"O�Ѳ�_�)bB��`J� �.9�f"O�-;2
ݻ(�BP��Q�0�ҨP�"Oʵ�4[�2� ]��NРs��pz�"O��2o�j_���P�����`"O�%ӕ(�
A]d:�gSB�|���"Ot]+�t���$\?uzv��"OST
Ց:#D-ء�V�Htv�u"O����Ѵ2^�"�#DpL4��"O����/3��УE#[?�J�F"OҘ�F��+J0�/� -(
���!�M/ ��1��H�GD�ᇈ��q�!��8b~���8
�����h�!����mD���?XM0mց���!���Z�"DZUo^ g�ޱ1�BVc=!��/Na��U�-�(e����9 !!��Z&~�y �\�0�bRC�X�!!�DԨO��y1��>q[�*�w�!�$�7I���V��28��(c�C�(�!��)4��q�0g�L���� !�$?c���1�܄5=��#c�.v:!��˖T:��DR�R7|���ᘽ �!�� �.MI`�1f���8�!��V��V�Q�	j`Ȅ��n!��S(PTp	��$؍H`HR#���c�!�N9%Jʉ��ꈷ�֩	tV�N!��T3D�,��.ݰlS��͏)L!�]92kliD��/�%r��׋;!�D�!Z�u��8*�� 
�� qơ�dM!�z��5���'ʙ�rNB�y"��$Ȳ����t�Dh"c���y�f�?�A�u/�]c�L�1D��y�dϖ@���'H�&r��M��y����O2�\��/ێ!�r]�oP=�y�)N>p���i����l�����y"��x�X���� ����ʌ�y�ƞ�^�\[u��)��!�p�V��y҄�<Lt�Ac��J�t7� ��؜�yrV����1��d ��j��y"
�h��Di�d�D�z��W�_��y2O�'=3xL�u�J�@K�4r���y򄐀.���{牾$��\H�����y��E5,�v!(򀋐k0N�Y'�L0�yrDHӒ�	�G �H��3c�r ��B��{�kG��ȳ"�p�ȓ5��5�5��k�����ށ��fhz����[=[��3/��*o<��ȓ/l�i���D("a �߲����ȓ5;��m^���Y���YAn��
�'h ��B�L�a����I�x
�'Z�Ԛ���.{z�I��F�G6��
�'�D�Y F���1���V!M�>��
�'Vx����.'���ˡ�ۅ����'����X=%��쪱ٟ� ���'oX%؃�P��Z�W���
�'~���J�h�J@��R+<U
�'�zH�@�X(&�u�� :�̕�	�'¨3@	��p������2A��z	�'�:pBDD[�sN��4��%5}����'�2�ӏܶ8�.[*�ڨI�'��i��c9!�%oK�|���
�'6�()7�[@���5�ز	B^��	�'NF��SA��) ��O�Rk�Ѡ	��� �푶�a���C�
/+�4�"O�1*dmD�j�f�KC�V�4�v�I"O0]�5��/���	��ŃV�ƙ�"O����c�L��Bԋk��Y'"O� ��Ŏ@lܭ0�*Z�8�Pyya"OP�;��J���1a��v�����"O�����)|�ްQ�i�d����"O��!���z�������b���"OT �E��1@XL�u�]�X��XS�"OZ�a�C� 5�p#�iZ p��@�"O�U�[�h@8c�I�?�N}��"O����F6Y��a�H�%�(u�1"O�A��I����s��?P�蕒�"O���'��*F��J� j`�"Oܨz���U'��k������E"Oh�����ڍ�jس�H�XS),D�ܡ�*�<r�x��Ivt�7C<D��9��-vR��4��-p�B''D��ZW�Y��у��w�Z��� D��2Sْ�@p���	� ժ"�)D�4�üb*��
՜M��4�I)D�p�eƁ�Ah֘9�HԡGg�$ʷ�&D�xs`H&�^U�ŏK n���H&D�̻���(�\�q���4uh��Q�%D�8sbď-QT��b.W:R��?D�
����x,��g�qDVjw�:D�8e�j�L1��ўL�2��5�9D��* &�vd�'J�6t�GF7D�L�&M S����
����6D�4��g   �P   �  �  �"  Y-  �7  �A  H  WN  �T  �^  Uj  �r  y  d  ��  �  -�  q�  ��   `� u�	����Zv)C�'ll\�0"Kz+��D:}"a��6���S65O
1S�5O�\q�g�:{`l���H�j�풁F͐5<:�� `E�JNd+T{��kc��Q�V�?�˖/��?�(#�E���!�1k��e���&Ot�/�Ip �tϔ�Kv�c���uG�K�`'���'�d��J�~��؇�	.���*r&��#Bl(�
�O`=�e]�E�U��Ʀ=�G���l�I���	ݟl���0��f�&�2����v6Z��Iԟ��4E���.O��DՍ6�)�Ot��7�4�cnNI����<���O��d�O��d�O�����6��.�ggD�03_��o��z���Z�,���QP�]^?	g_�dCӠʻ<��Oĭ��`ּ)��UYIſ"��h ����9,��yB�dſ&�N�I�G�\��!1���2W$�J=��'�*l�����O���O��D�O��d�O��'�y�DɶTRh�7-I|Ǝ^�?yS�i=66�Jۦ`ܴ�?���i�L���`Ӏ�@�� �:dSGi�ik ���ɕ
��Q�"�Hu�'D������45ii��
d�6���ם�K�~$ʖ��);w��Rӣ]0^�@�*��[���"�Ǖ/\0j o�M;��i"���w>���ԁM��$9���S���
�SQ���Ej�R���j����@�c*�WV�MyشwLm:�O\��M���i9�6-�
�ՈS��>b�X��v��N���h��VVH�������qK�4"*���F%$����C�;�KF"v*�u81�Z'X�	��J��a,Tq�A��3!�uB�ϐ�
�
��ղi��6M�������Q!V�D�c$�2��钧��|��V��hf;�Ú�v�$��wӊU+�ԌʂY+ �)�����O��dS�
�X����p����0�VhZQz逅�I���	��M{�'���E8T0�a�����?Q �B�H��w%�M��(�c)Z�?�,O.���O���н 2ݱQ�V�o �oڭ2��s@X�iXx��"Ǉb���Ics��aPD�#_~X��C���ʰ�T�D���p�KD�Yx�!��H�����\"�/i�I�x�\!x����0z�%��P�2���O���.��O���<��G�6q8ǁûY��2A�C��\�1���?����S<���H>	��<ͧL4���+gJ�CsG-z� x+u��6�?	.O^�q,�ݦ���s�'�yG#3 L���Q�$�,�(�N��?	��g��/��B��<��iIR ��	#���&!
�:]��@b�3?�d��
�bW4����૛3�:(���F�8xe%?A�H�4\h�h��3s�6	�W�2?� ����	ܴa�>=�'8kn��q䕮y"0�i�!��Tp0&���I���	zy���>
,��q�dgr�h��i�ў<�I��M+��ie�Ӷ�Ӕ>I�]rbVTm�OG�S��Hm�����'}�D�7�O��'��V��3S(�!���j��#�@X��I�񈈃ڴah��IU���0����*�T��ڸ^$=k&�L ��-I&#K5H;F1z��^/Zr��Na;買�i��SU��j��v��Uf�Z���(2Z8E�޴L�剫=>^�$�4�g�ɀt��У�F@4����$e*>yD{��'z�����l.2A  ��<������?1��iB�6�/�4��)�<A���3���F�ن|�Q���B�8�[���IΟP�'���|�O��Y~I���0��]�G�TQÖ�a��G]>t���4_����"S.�P$�83^^��PN�<`i�����@8� C	��,t� �����ɑ=a��Gc�:!�0����p]��9�I�O�o�>�HO������+F��a��![�&}z'N՟u���'�1O��B�g�!%ft� �'T 9ބdS�'�6Ml��nڵ�MK)�NA��L�I�	�XAa��>�V`AE�]t\�a��]����	+I;.���ڟP�����$���k\�h1JP%'�k�Gb�H`��W#
�!DFʎ`�ax���i-�% @9&��ǇO?=N1��� !E{�Mս�j-1ĥڟ}�P\ S%���m
�O����'��I}��d+4�E0���=������# K��?)��ᓯ~88��2�I 6��M��#�0���L�q�G�P%#�D��D��3Cv�]�VD���M�(O> +�/�����I���Ok��x7�'��!� ��O�l-�Ŋ;��#�'`�-�`Ěm�R�S�>*!����O��������s����D�,���Q����O`�y����!R�%Ś>�0a 璅3֬7m�z�t+X g�±��gD��k������O*�rӬ\&>�|����~r8���F�S��00�I�	��H$�Ex�m��1�V���<	Δ������O�pm��M�K>��eɦp���@��K7��ڃ�N?YX���'�B�' ( ���K���'��'��.�]�
p��Hj]xB��+!�:��D�L�-��E�:B��s1X>�<i���_
$u(V�I����J��>���ئ�ߞr��h�%K���� �K����i
�[�5�@x�j^�*��` �wqx1#Ӂk�J�;�O�)qg�'y1�b�'C2� �
��0��8ey��Q���fk�'��'� �x�W,`�	��̤q����-O��mZ��Ms��ۛ��'��O���&�%���&o�
]HQ����)2GP��M���?Y����ɏ�DY�d��su6`�u�j�� r�&�cox�9��O�o�@i˓=�:L�u��z�:����T�F�XӁbP�m�ܚ��#	���[g�'����'ǈZà�2˜t9́w��-�?����?i�Bᓫ]�F�i�$Q9x�$˕a�g8�C�I�Y�p2��-%}�\*�
E�O�m�ϟ��'K�18�)m�f���O�� ��^�<(k���V��@�OJ�D�n�&���O���V�j�:��d�� c��rGN��5� ���f�I�Hpf��'��f@�!��'��� ̚�"0�!NF�r3����QP/�y�4�jG�ӵD�\�q�	1`i�DC�u.O����.�`�0�0�!'���ԕ|��'� `2��M!'7���8|�L�����>�#�i� iQƍѰ=~�tK�����#v�qӌʓ+tbI�׶i��]�h��y��֕r�"��p�M�#(}Ӌ��ikb�'�^@��'ފ1Ҕ���@Z�H��q�p��^d�`���M H� /�c��G���1C�S�����@�L9"�-ʕ.3` 1�O���
;��K���'P.��Oz�E�'06�XH�O8���%��X�R��l-����8��}"�����G0L�j�ha�Ւ?b�c�*ړ�?��i�46�5��G��x�� -�"����:r2�D�O:˓>���P���?����?a+O��� ǅuR�wd��w�|���1XA��� MG�1�*ۛO�^�'��=��B� } 5I]�y��ZT�ޘzH�|!���a��u8V�Q�F@���|�u]�|5N)�L���ci!���@U-s��ܸ���'������J˟�'p���r/ٕ"Z�Y�oKS"ٓ�\�0�	��H�	v>���˟�'�L��P���{�$`��O��������޴�?�f�i����?�O��C�@��#z<,Q�ና?z�q�@�Tr��P��'	��'�bai���	��h�I)RI�šco3:� ��M�1�D(��
:���������`k(OL���4		:��Ԇ  5��"�ӛb 3�$0{M��	3V�;1н��H/:)� �E�D8rc~����U�\����|����O��o�7�HO��h���+M�с'a�c[2�y������IޟlE{��me<t��)!)�.Eib���'D7���'��t:`�q�|�D�O�(8����'��c�I�K L!��/�On���
n����O��)�l�5bƏ[f�����՚djNu�BOaٰ�뱨�#�L!��)<OH�j�ДU:�q@5�Ԯ\�xը$)F^~��ζxq���#)��c�ax�+����	A~�b�8 7��I�!�-C쀩i4B����0>�G�]�Kc�l�v�ClҪ��+Cd���a��:2�a��J-j�zL�U�Ȕ,��!�ILy⋂�	M�6-�O��$�|:�ߵ�?�S�^&<���(�m��3j�� ��?���j���r�g��+gй��.S�*�"m�.�p�%t��˶eE�e�|%�0��^�0��'��)�Ӌ�fy+p�U�j(i�ض$k�iɟ�D�G�	_(0��U"y5����L0�'�b���<��TI7Z4�&�zTv�0c�B�<9Qf]'������Oi��z�D�~�'�"f>�Ӧ[�FB?h�0h����v��u�CLm���$�<�$Aǂik�	���	ay�� �։"΀y?Ja�-��-�v CP�3(�����\�{��آ^>��3�	0/̸
"M��{f��#ŘG�&�i�E���6� ��H4?VZ���*�)3ZmH�if�P�e�\xh1��ȶ-SR%������(O�a�B�',�d�?�O��!�Ӣ@�%�b�[��Pi��'���>}�ň=|���r�/E�/
Ԩ�+�O���Ҧ�B�4���|B�'��dM�u�TU���nW�c$ W�s�~i�ߔ�N���O����OXQ�;�?���������bkT��1OH�BL摑7 Z�E�>ݣE��!.�Č���_b|1��	��jx3mN#q�� g��!⸋��H��8���G�vuk��'66��br����D3֞�2��»@B�'ў�ExbƓ�\M\	8�nS�m6�]�U��3�y�&�.\�m�U�>��-ɔ�ۯ��r���'��Y�T���4�?��J����" �$�x7��:CB5���?!7����?���?�3��?DO��4ꖁ/���'M<��h��N�v4n��w"�27א��	ÓV�Bxb�62�t9�墙Y�m
���y��҄�E:��'���9��d
Nr�'�H����?qS]�x�@���:0�\��E�OL���O����r̓N�^D+po׶H��#�ҋ�t�'��IJ���tq�:���a�P�\k�A��H :QlEæE��-�M��I���'���'���C�d'��&�tY�&�/@k:�hO�`Er�'�6u���I�8��?-���'k��Q07,@X�80�%H&o8�%Z�O��A����\��:O�"|³�V�[�8H'`�����LTD~�n��?��i��7-�O<����C2����'b�:b�yi�9� �$�OB���O:�$�O���?����4��$g	�1��LXS���hO����z}"V�,��hC0�8��N6�丸u���ҨY��4�?y*O� ���~���O��d�<�q,�!�D�����1�']`�@�d�~B�6�Z�XU�U���Κ!������۾04�"��g�",Qp���r�p	
��BN����)�;pNZz�9OJ�+�><���U���QȈ���'����,��D�O��$'�I0{��q7ǺB� %{�#Ĥb�����}�:�F��|ov��5H·>�6I��џ�0��4���Ĩ<i���	2��ps�&�m$ܤ��m�p��F��?y���?y��z��?�O�Р��Ē� 7�9���-ja��H0�5`!��q��q1x6�AX�Ĺ��(� ��	��
�D��ˌ�7��$�ɟ`���qo~�*h�`&S�x�Fd�%И��{~BBC0S-�1���~�f�0�*vi��	���?A���9�����T;��J�J�`0Y�ȓ+>P�C�	C�Դ� "Z�@�%�H[ߴ�?+Od������}�Iϟ�Zf�T'��H�6- �H�: ���S؟4��+U������̧0�H(S�-�4z�:��B���M����Vf��@���U���CB�r������V�'H��`��q�DQ�$D@b�R�s��A(�aL�J!��ݓ��8�Kӟ5t�sJکg��I�=k4���w�	�-41�K�A��Y��Ԁ^�C�ɏ��d���׸}�<E��Q�9�N���S+Je����ʐ�0g� ɧH0��O�,ma��a���'P.����-4�R�q�'
�6Q�8j��']�菇c��X��>D�7��m�?qQ���Ɂ3nRx��l��B�\~b���9��L�	ƛV 	�(� )PHM�KK�A"N׹ ���K�����D��<	ҟ�4_���'���XCg<k����f��-�*�'���'��I̟������I>~FT���F��J�Q���=t+���V�2k�Iן��O�������v�a ��ѿ_�|9��Ë7"��v�'�B�'��51$ǝ9�2�'��'^�n��}��Jce9_�Q�oD!3-z듫?�҅np�X��	�r>�4ZVB!��@B�J�1O�#�>v ��T�d�|�<AB�K���%
R^���K%���Msw�i��Ƣ@��O~���'4B�'{"��9 �L���I��&��r�ǁ<b�'��Iߟ|��`�3}B�@d���"�G��h2A���?��W]�	Syr�'O���'��	�'�>T;��u?��!�Ě$0�<��C�Lrd�����,��ǟ;��$F�^F�YB2$^�$�<�# P�3��g�%��AQ�N9v�7mۦ��e剚i߾��&^��#C�6�tQ�æB;AK<m2hP�=��(�4]��}�ްP��ɂ(����vKx�e�� �� ��a*��×��O�@nZ��HO�#<�rƍ�^cB؃�@Z/�ީ�g��O�<i�C(WC����X�^L��(�IT��M3����D�A�`m˟T��;|F�-"_x�����	P�F���l��CT�	�ϧQ��a!L�?���Y`R��Mǭ�1*�	PN�l��Zw/�h��ݱF�B�'&*�)S.� H�R�sT(\Z����5AG�Uȣ�_:`�Mٙ\� �4c��:���VB͍��	-?x��U^�I�<8�lK��D�<��#�X��@C�	�8��I�и@�nO�1i�.�OM�I�%���*�Ȅ�"W�4��RQ�̒O`hȀ Ц����<�?1S$ĄC��y��^�-���ʋ�?���/=4���ѡ���H��J-fT�QaS��%���Y�W�%�\�(KHb��I����1Z���@��}lV�+B����)Gl�/b`��V�/w89#�&%�����ç*D($�w��p��O�}$�"|:���C�l�``� =���N�}�<q���m?~��w��&	y�%8�Y@�']H�}���o�Ψ  LD�46u��W$�M����?���lҨ;F�A�?����?I���y��H6m�S�ìu�|�rR-�~�I w�ޞ��H[�*
��8����yB�7T��� G��#n� ���/��h�FNƄT�����_	�vx�}�<!�f������a�-we<�S��K��P�'����ߟD{"��)\�8��$N�x��ѓ��,yj!��	kW�	i�!A�Oi�<;���h�	8�HO�	�OvʓZ^t�'��(�#a֑<���ro͌5S�Ey��?���?y'���d�O��S-\Ŋ��+�(����QL�X��W$o���(^�a!f6���O��:���'yC4K���D]��s@��*��Y�4�3_�FyIt�ib��b�-x�� !����b�X�(Ѹ��M�n��� �{��I�6a����4]��DTG��U�Dy@���$��@�d��pɇ�IK��xy�!�ޠ
6��'dQ�Y��'�T�'��+[��,�O���\=3�njF������l`���O�-��O��z>YS�)I�<���Z7:QBp얀Tk��j�,��l�f���J�"��dܓj���pT�O> ���e�1��@)���/1G��4#J�=�� �P@�@�-� �I3�~R�'I�I�n�J�����4��V<B�D�O:���Tx���Ɯv�� �,��OH�=ͧY���s�e*T�7	��C�H�?�+Or50
S�5�bs�A�?���y�x#�/�&(�x<y����?	�j�z�Ca�� �^С H� bx�%�&�x������Aֹ[����T�z~PD��8��!F�}��d�ӬXa2{t+�hpN���� ��o)q&.8h�<�U�ϟ>F��jg��Ta���O�5m���H�Z�S�V�r{Cѿl���y'��g�FB��D٢����R~XȚ�&�eΣ?���4�E�3�C8A�R�ëdV�Uo�,�	런��k�\:P�	֟��	ϟϻb:�*�f�^�䰁b�F�A� �E��k�Kf�itpɠ�(˘Ϙ'C�u�#������&�z�zW✳BBxY�Smv����']��c>���ƺg� �)� N]�+'3�0���Q;:^@���v�rȖ'���)���͟�'�4�X��<<�X��:\�"O�V��a����vJՀ"�i�'s�� ��|2���"?�i�O� �L̓��2O�T`�5-H�>����O��D�O:���?����ԭ��2YL8i��\�W����3Ã�� DY�e A�qq6J�=G�h03�M�_0��EyR�}���rp�̥FO�MÓ�U
)Y$Y��ȹ0q�hc��,<���a�M�_�R$FyOE�!�B-h�h7Z~:�����j�y�����.)��O�ٛ�,N<y���!�O#<�$��"O�Y����7o���Ŭ��Q�X�{"�|2Cy���Ī<��˃���SΟ�*�AP ���6c��۟\�	�G �����<�'4.�� �$��/>���	�l����r_���@�]:I�\ʧj�7��Oh�8����g�Ф`�Ҳy�����ʺy�l5kP�8 B0�C����t�?�嬁ԟ���R~�$Rφ�qq眏�h�$P�䓆0>	\�� S���|��3j=L��$�ߟP��#V�!�a���o��`�OP���ؤ�i��'���]� \�	�;�.0;�a1(�
�K�.ՠ$f�I�P��N��T���"���+���5��8��`���ܣA��Mq1�F�J3&P"t�اpO��A����'��"�\㶎��J�uaį�l� �Z��"t�F��f�ô*M����ɵ}V^ո�"-?QՃ�ǟ�Xشt��>��S�Y�:�p���R�>}b5(%L��(��5�:��Ă��/2��21��v~�QD"E-ڧi"M1P+
�8^�v+��F��(q�4�?����?�i�//�p��?9��?���)�ص
po�I������XV��q�80��@"��wӴ@�!�F1CW1�1O̼Z��bҜ�¤�Bb�ţ��#3-��yP!ͱ-~9�TF�'
r$s��ژ1�٨x67Mj�-��&fuz�*
	^.���2N�O.��\`�	ȟ�F{RJ�$��+L�ҌG'	!�$�+q���t۶���Jf��sP����4���<���K�P\�4B�쇳��Ps���I����	 �?��?���J���?�O�(��JC��~� eн�؀;���D��4���>>��s¨",O>mȱ X�i����� [4̈ځkI�m8�혧���0�V�)�r�e�uӴ�A��_�1���T8��k$�١!䰥�@�UP6�Q�Rԟ��Iw�'�����Ǒ��ܤB����E���!��x����4��*]s�)��M?7��'�<6�O�e��Q?a�	( V$  T��:�|�q�e�# >)�	ğ<{�i�ٟ|���|��N�) �&%@�ǐ?7_)B�ϛ�8�b�+0���BD�u���������˧n�6�
i[@��8���H��H���<(���Ac��DI#�I)i��d�O�G�dP
r�S?)��䐡�Ãq��X$����	�bv :�&�z�Z���,�+�\�<D{�O�v��Pr(��x��ӟ!?XqRC풾LS�,c�g���D��ڟ��O��-��'8����*Z�ϸ!`�=.͜��q�'���I�e�3
�9�(4��=(�\�'��	�(!pJ|�����%������z���O�6@ 3Ȗ0!Pȴqu���5���iv�?�I�d�llz ��J�{�m�4�/?y��ܟ���S�Oz�$Ėn�����3�Ly{Պ��?!�8X��P��	Y?P~dl� ��
9ў��ɓ�HO`������V��pԉ�y@���P��O�d�<�����?���?����� 9�B�y�E[0<g�����&Nِb
� WYd��0��W-: �b �|ڞϘ'T�K��W(}�����?�T�jG�-d����4�йk1 ����%�Ϙ'�5[�eP�Z{I�.��\�������8\B�'�ў�2��K�
�4mc�E���̻�MH�<a�#"ym  J`("� �F�^y��>�S��Y�(��D֠k��c�#�J�`�  h�=�	�4�I��H���	�O@8 ��	VR� ��B�+kH�ᗪY�c��!&�-�챱�H��x����0a��ru�Wh�%X�6��)��@��`Q��x��	2:Z���I�H�̉�����pR�Bu	
�{ܐh �C�Oj��3ړ�Old�EņV4r"#B>*9�B"O���3�ܰ���:�-
?�M�`�|B¥>�-O,YKR�K�t�iy6Ε}�@P:VZ.q���Ĺ<����?A�o
@]:�	_䝯�k���;T��7m��+���w<��� -}�@���I�g!� ������Q���/8�����Ͻ��q�ʀ�P~�ɑ�"O���D�'4����%g֤Z��{խDo ڄ�G, �d$�OX�8E�#G!iQ�!��ld t�d�'���Ć�I��L���'ute�@���Q#�\�t��.Byʟ�ʧ�?�6dX�plh��@/A22���S4��?�����j����r��h�BT	t	�Ty��H|%�À�\:��p�g��1{�	- �I�#-�b.4����ɫT|Q>��v�C�-r��)gT�  ?a�&������L�O�� ��jW��� L ��朩gMT��6"O절7�J�x�6ԋ�J�JfT*w�	��h��D)�
�@Z��H��:��W�g�\�Z!-�<1���9���	�m"���1|/��r��l�X�g�\�
4\�bd�>�ʵ���#�3�	.��k����_e��!/��Z#.��c�U�l:L�Z�A	�/��-:6 ?�3�	#C�*1"B����`ek;@S�}nZ���d�+[R�O��3��t���g����;�$�s#�B��*�}��c�S���y��
�
�j�fɑ��'��$\�b�( @��B2v��b�5xiT��akҦ���)1\O�Y�6&�6_�hH�b�/���烏�u�p��HʈfMVi���յ�p<�G��<%��U���rM�0f) e�P�1���m4e�͖W�����nD�EL�;2yNJ$%A�L$�%�g�'L�7�M�'����Fj�2<�g�1rUj1	f�7D���6�� '*��'�2�d�P��"��UM}"T���l	��Mk�Qr��
\������J�� Q�LL�'0���%P�>���&�5�ș3a`���|���!OVp�I	Bٚ�Rq��$�L���-����D��S:RG0����Y��T��*�Q��.�!��ϕ���
7`��&��9���v���O�\�i!ʩ8ǧR� �
��g�|�f�><�6-�/T�Q?q��
�z�(�4D %Р-3�-?y�O��t8��j3�NRMt�h�-�'���	�
�rR���`�7V��y�'�|�أ��4X�6���e&�
�D���@�X1�� �e�u�fѐ�Ы������%i�n�D�43�A��&
�}|<�pЭ�-Vh|�""O��y�Ì?@\x��չPX��x��	��h���� gS�:��� ��0��o���h�<y�FS*���	#8a�c1@ʍ,T�AHS(_�H
"b�\-�:��֗�~u�b��.)��L�c�I+1Ot� �'�̅ˇȷ.`�6IC�A�E�S�|B�C��?����yb�F�zc,1z�E�d��r�ӟ�y��əp�a�Q��	,@�6�ʕ���N���Z� g�).�F�A >`�r���ɜ�v2�R�1O ȣ�ԟ�WFWV�䀾}����a�e(OK��$��Y�s���O��87)�O����OZ �^%Gͺ�V�\/!�T�y��iʉ,�1�2�O�r,{wm/x��@҂U91}�`�!g�U�J��5葌**�1����'<��
�n��KnI؄�
8Xl��~�\j�O^����'����T4x%|xA&�
3�H PЩU=d��	q��\;�H�.Ĩ�K /ֺi���`�6�O�l�'T�뱍��M���5�ҙSS���-O�ui�d�OL�d�O ʧC�ȩ���?�bh�2R����
�:J� �T��.�?��Ȍ�J��-�G��q���Nq��Se�4ԟ5�7f�2p�(�;�� �"���2�'3��J�M�0tJL�"q	/��p$ J.p��;��M�2�<A�O��M�#�U7������	|��qU$�O��.?%?�'�N(��X�b� �$�
�+�'h@�%�$T{�8��؃dw6 ��d�e�O�xD�' -����#�2Hrs�'&R�'�6A����6���'��'�d�'z�tE�&S<Hy�M�R	u�aZ�HV��n��;��SȌ�^n���j>#<��C{f(YjuȜ�
KS$Bj���ae���IS�]2�[6�������O��Iڥ�O�u�H�(�wx�z����TEy&|���O<,���'���	�<�d�h�V\����Y���Ju��{�<aF�R8@@-b���#t� ,2&E�x���4��Ĳ<	Fꁫw�a���%�R�yP�æ6��.	��p��ٟ�Iߟ$�S�����|����f�ʌScJ��E:�ؓ�"��wZ������ν*�E��\�D؊��"Ơ;�F�J��I e�P�v�VU�5e��DW�t����R��-�.[�iS�m�'�	8,�*�dۆ@�(��`��Y`�q9����&R�$���O\Tbʔ�JeT� ��\Q��:A�'c�4R���E7���4 &t��!�<Qq�i�U��b�	�����O^�ӽ �u��Ρ�;aK��>K����b'����OT��)?t}Yu�A��^�2bK��&.��4�2����ցn�lE��'*J">ad �%��e�/��:��<�f�Wi�e"�	W[ydt��	� �*,���>h�1Dxr-���?y���O�4�ز� �������ƶW.r�B.O~��ā5ޔ0R���W!t�
 '���''ў��#���	E�XAs�!P!4� م�֦D��ɗc�F��I֟���n�aF[I��'�|	�B�� n������P#52Z�0��'��A%µ|�µ:1e��������~��Dl��6xZ�j�*�Wg�X�����y�B0R��	@
7ȼ[W(�
ZEk֍��O4�,�c��0b�|Q�⒁Ow�K�'��	��?i�O�O��)� �e�e�ٲ23�Y�ňɯ�l�!�"Ot����\G@��)X"x~]9��$�O�Ez�Omh�YA F�_�PX��E�-������'&�'���9�J�5:n��'�2�'����'��/�Ċ	Z�� 15tYIgF!0���q��\�O�����Rw�Se�Z���Ē�`��J6!�	;T$�Vϑ"I2���l�3if�,Zg��H�<3�'R~r�S�Y��h�,�F ����!��D�8b�r�'Hў8��N����)[n���T�l����[��D�:	2�Ux�.ϟ~�=I��4둞��ğX�'��T���ӒL����@�!{���3�̛E1��T�'$�'PR�O�B�'���|�ȥÑ8���㗟N̔�0��67Z�����]�~�1�Ǉ"��4̈���,��`�!�7��XVj�����cj�a{�L9RdӖ\�<��I�Q�'p&I
��*��8UC߫X��2	��|����hO*#>ac&E(�bm�-\�聚�'px�tExB��6`��[2!J�/�uړ.�?����y��Xy2f�?@��7��O~�|>�[T�VN_*=z�>Z���O�'��O����O*�"��MI?���jF&l|n�N���R�o�p�C`/Y��TQ�@m���9�9�D���4�HQy��M㧅��bT� �-C�!���#���베X�2P3jQ:���A�&��5�4�DPh!N�>w�a���D���3�"O��N<}8	�I�6p���'���>�ⵚ���mvf��D�M��՗'"B�'���ȕO~��G��W
[+\>�H g3=��?a���ߌaJ�Iozi"��#���n�G�I�7?�O�!G��b�$�t���:�H�aF�k�F�DPd��	�;�6���O*���O����1縙���9'*�B��.|I�DJ
Ѧ�� Z*� �I�?aBm�dnz����7O��]v�
�Q�`�B�i��00$h��'R(Te���b��I̟H���H�E���a�> 9�0D��e*��I�I��@0��3�������(W��D�'���A	
���2�'�7J��d�{���'qBe��$�~�Ϧ���?�	�t�åc%B�F�q���I���_2 ���ӟ�4a�쟌���@�@q����g��_��@�_�q��]��ŘjҴ�
ڴc��н�?)��ZAhifQ?��	ڟ��3V:����ȽF����/��5���!�eN�<�NM��l�	�ug�'��d�����i�b�jB�`�9��ڴc��y ����"6�l�\�V�[릕��4P��'��������VO������R�v��E8{6oZ4�J��_:�`��4�f�Of���Ov������@�x���{N�˂��Z�cF#~�<)�悏�q����M˰�O��6���p만J�� Bo�kua!D���3�	�!����jD��9 ��F�,��&�'�2�'���'U��'F��'q¦�-�8EI����J�Q腇cZ7��O�D�O���O���O$���O8���"	�����\��G�@��m����П��	�t�I럤����P�	A��Ԉ�J�r5�9�#�/�:|۴�?���?i��?�(OTʧ�~R��3li�w���lZ!�7)�6�M���?����?q���O�!t�J.\�P�2{u(,�U�Ѧ=�	My��'����'�?��ך+�M@��	�6�Z%EVB�ưi����O����O����|�)�k̑� o4 ��[�,�`���>zI!��=[��)Ӥ��p���2��N/C!�D̰,A8yx������/�!��n�j�hP)T<�� +�M���!�M3X��v�ӶV��y0%,E��!�DJ*�FUK��z�����Z�x�O�%24��8"��*=�
����[���@�A"��E���[�v�P֥hx&Q�̑� ��dh�)�O.����H,:�� �G�[�~<����X�f0��'[�'��\3䃊 )D�K���Fe�U���
 4���֩h4.�3FJ}�Y	@��VSF�*b*�� � ��>H�A�v�ٷTL����̓m/t]0�$�|���#ŤɅb���2Mcy鸧���QT�H�wa�@bSna �20蘊wn�nZͦ����j4U�7 �+x~�a4��&U�'��i�'1O�4&?9Q�J�v(��d�6@���9D�lZ�f �XTh(B�M�B��h�C�I90��i�H۞ KҬ2cl�:��C�I�VԨ �s$�Z�RpӆW�g_rC䉱2������w�2�&�0x DC�I�zȲ�xb��z�%yc���8q�C�I,;}R��S"N�Y�L@x��9��C�I(D�քy։��_^
E�w*��d�|B�I:KES�EP�TZhx3���6�jB�7t�� G�G�~�NU�U'�[�B�	#b2��VbO�dy��:�`B�ɪ��9#�Ìvh�ypA QM�C�)� 
�C#����Ȋ�\��'"O�t��$��i|�GE���1R@"O��gYM8AnM%��PrC"Ou�_�Rl���*
#tؔ�U"O�!���@uD�<2���-fw"O4:�J	>��5Hԁ������`"OܥYsQ\gUB�N�\�"O
d�f;T[�L�_>n9�"O<�R%�:tT�0���L�:�H@5"O��8�G�7�b]�VYO����"O�\bqŜ; ���P��I�IKT��"OL� A���2��҂޴^�Qy�"OJM@Qd�$w}V��F��;��"O��Y3��^�T�2�j��`r"O�k4�J"��J�e��(. s"Or�(�*��H�4((���D�W"O4}���I�-F@�D�D�1�"O�\B+�;>o��Cuo�ْP3�"O�
� V�mj�M§����Вq"O:m�ש��Xt���Z�$ɬ`�"O M14J!�|p�`׺5�:*�"O��8���P���B' ��)�}�$"O0LH�N��GIƘ�2�G��a��"O@;A%^�@��K+�4�id"O��h0�Fz�e�a 6#�4@9V"OF�+�4Y�C�.���u�Ǵ�y��F�'X�)Wl��g����Q7�y� 'D�A@��^�a�����$�y"�0`�Z�"I�W��!�U�<�y�U�L�.��G�t�85)Ő�y�*ؗ,r0���C�L�����y���
�Hh���l0��y��Pb�6�Q6��a�0�D�9�yr���>�����Õ'A��Tʴi�!�y�'
&e�(��F^4��UK����yr�4fʤc��&�H�T�y� B4��E�$ƽ�����C��y���D���B��%�PA�!a��yb!9:{�q�V:țQA�y2`�ml��Q��
yq�R(�yr��
\��0�6�F9Q� fC�y��%7�j�q���9Z0�j��V��yr�Y%������M��h��զ�ybύX3Ԁ�5�A�IVt�r����yba
�1y�d�S�q���C�m���y�,G�K��:s�0d��Pm�*�y��`ؔ��Ҩ�H���:�I�"�y�ȧ�X���X'>��3'X�y��S�Id^�q�a�<�t�W-U(�y2�?/�:5�uNM"f�*�x�-�%�y2焳3?(x����n�J8yŇ��y���B��E��Gh���h�yR�ƍRɹ��̎p�	�@�,�y/�N%8��ݚw�|y"L���y���G�t ���l~:�bB�y�A�����P�3`X�k4=�yr���;yR��N�S0�׈� �y"���N�L�S��[��v�jVbZ��yF��l5�=2k �O|@�۵�y��14��ga՘2���5c�+�yB� k�z����Z?%�Э��)�ybi�ZE*H#w���E��0�F�Z6�y2�S/�) m�E�X]ۥÔ��y"A^+C�� w��tY�IB�y
� ��/�b
̑���x�0�sF"O4��
�a�	̀�	��:�"O��b7#RU�Q��������a"O��a��j>��ߐk8��Qe"O4�Ac-��@GJ�d��5��#F"OhA`�h��l�����&�-��"O^��!ՁK�d�[�bUZb�X�"O|��B`�-[�X�K�A*9_�E+�"O����j�B��Q�mX02�"O�@�`k��QI��C"ɓ:�B��"O`�S�w��թ��@΢-P�"O�U�Af��hܘ� &M��4�C"O~m�)Q�(��<SP�ՙe�h8�"O�`����)"�|pX��9B$T���"O
	��Ʌc���t��@ �a"Ot{B��c��8�ܣ{�!�"OYYw�<v�@AX��;s��2�"O��@��6�2��`�"u�P�Q�"O:��`Ó�/��2@�N��"O"Px��[�V���F�� 7xp��"OHl�c{�Xp�m+��uɖ"O�m!��&~ �5�M͌\"O���e�7'��s�
V�tt��B"O��K��-?w|�2 f�q��"Ol��_x��,Qԍ��^�c"Ot-H��sGh���� L"O�цƸ_AD�T�,yz1�#"O��cʊo�j��
�m�@���"O6\`�.˪K\pU��P�cg<�C�"Oh]�5��CIH�`Ġ�0��r"O- t�I�B��9�ӌeb9�"OMp����>S���V�aRL0"O(�js��A@p��rL3���ۥ"O~�{f*��q%E��Pf����"O���%*	:;j���ՄLaQԩr"O�5�AkF-�2�x�N7+G�$��"O�aۖ�-\���zF,R.tC�"O��P��2��5b'd+X��U�"O�pǨ��G����N<r���:5"Ot�i�����8����=�yC�"Or�[��M7;�H�Q�	a��"O��AL����@_�1�-�#"Ol+����׬Ԧ_Lq��S
�y�ʍ�i]5���r-�ek�=�yRI#(=�c��X
��W�R1�B�I��^$�s�S&{�rX��'2w�C��;8�>�qs���'N�%��)N��C�+�Lm	�/(�<9��rќC�I�ge�I���X�7t~tؖ��,�C�I�K�PJ �ȇP�N�!R���~,�C䉏f�h(��N�\�"G,Z�>C��>o���s�,�w�b4c�S���B��^�& p�I��>Z�� �U-x��B��^b��@�ǿ?!�ڂ��-$�B�i��܂�'�"�J@�lO��tB�I�0
�M�vד4w<0c��)�B�	�c�+emQW,&X�S��<��C�ɽv����`���Z��-#��Ȑ��B�I��D��Ȝ$$�I�����"�`B�ɚ�>)d
Υe�=;f�UD^B䉓`�&Ѐ�(�-�5�E�'RB�	���Y��ȿ<S��0R�FHB�n���hF I=:�h�s�õ!�B�I1&�[#�V
U�X�6�3}��B�)� ��G�Ɛ�����˪o���I%"OpB7 x�a��F�U��xx"O��궡Y�lY��Y�Z���q"O����ޢ R�r��V�ȉk�"O$�y!mR��l��%�:8X��2�"O2Ṁ��|�p1E��3S���"O���O=�q���p"� �"O��)*��f�R��'0��h"O�,(5���
Iy�'ڴ7��ʇ"O@��H�d�fK ���1�"O�Yy��8lUz�*�<h�����"Ot�x��Wa��У".X�<�Ma�"Of 
�F�5�@��5k�l��"Ol�'���X9�ǥ�@��e�@"OJʓd��I��Geϕ��y2"O��1C&Ƣk^"�dZ�a|UQv"O��#r��S �g�ʥYD�x�"O�jr)�@A�A�3#-r��{�"O�48'�-Q�FLˠ�D17�� "Oz�A���6'�ʄ�ga�IL�\s"Op�v�V��D��f��%!f,��"OZ4�@m@�:�J��Q �!]�<(�"OʉB$(Vo�	!��;A����"O�%�EmO q�8̲�C�g����"O��ad��Y��B��G�|��S"OLX��,�K˰���LE�~�9�"O�`Ċي^��� ��3Y����"O�L��jB.�^a��G�=��B�*O��i��v�� �;6��a	�'�J��s(�-VΰC�'r0��'��A�$�Y���\@�� �L`��'L|��d�o�8jP�ߎ��i��'ø�I�W�3y���V ����'��2�OM&by����k=#Ҹ��'���y6���
G钜QWtp�'P�8BH�w��X*%II��'�l;�����.���B�
j,:)��'B�I '"��qsĔ�WŊ�d��*	�'��eѓC$2�;��d�b���''&�[��F���87�.
���'��A�R��
x��/ ����'�Lu��'� ;d�#'�N�Bo�-I�'��M�jPYB�$
S���S�'��5)wG�~�"�E�F*x�R��
�'���H�DC2�ĉ4��wh����'+�\R�B�>���:�7Gq8��ȓw'�ٗ;��"T�]�5�b���2�����8�"�Y���g��Xb�'.�̙�EJ�=�L��$���t����'r�ӂN˻>l�j'�I>�$LX
�'6`� cK/ZK�ѕ�Ȥ�h�r	�'�Ҙyݘ+���Qm
����	�'��(A�r�(�j����
�' 60t�ԏ'������	�l\��'{��(�Û�_x��R�	�1 �'>�ۖ�X]�H�MG�'��	�'�z�����0`��[BiFs4Ii�{2���/�$�ׯ\\,n� A(���Z��L��݅sȤ9$�
"?^���r�6��$:t}Y��M;j���]�̴H� �-h�>i�F��j��D�ȓ;H|U�&�1t�
a��j��`pY����E��*0Hd�W�����Q3�	�çS��f������W&8ńȓ����,��I��xC��Y�~�q��S�? tptN�n�y���,z�x�S�"O^� ���|����Ulӓu���&"O򐻇HO��x��0,�B��5�!"OJ��6�@�G�b#Vh-��T�"O�u��I��V!` �2Y��!�"Ob|��A�3<��e��Ո�z%"O��&�?�$�PN#:k�Q�"O�  ËBT��y��7T���"O� ��ʕ�|�)�`����S@"O�5�$k=�rl���v�\ĉ�"O�dA!�S:yr�-qd ��C���1�"O�s���'[�k���6���%"O\�@��CT���e٢4欰sp"O�SF�/e[�X����x�n$G"O�0KQl���\yU�U���T!��	���"�H���aW-N��S�n)�t`CeŊI�I�ҫL���C�	m6@���c�-K��ʘ ��d�1*H�3�ɒܬ�8ͨ�6�*�M��xӢ�t-^�,�ף=D�Xh��F����9���-c`��2.��F{�8�Ìc�lL�0�*kc��g�':��z�F�i��q�&L<��2�l|(�3��R�gN�SЫ�yT� �C���E=�Y�Ea �OK�Q�(�k�ł�{,K'Ŋ
�hO`R�E�v�U7K*"�P$�����\o�%A�i|��q��$�!�$�P_�5���ٸtZǤ��*��R��`�ɒ�[�5̺���$�U�O_���QlR�k�Fy��C�<2��'"O����& xls��iƺm�a�8QΚl��N �:A�d�ˆ��3����ل	��teЦ-K7��M��I'2�0M3��.����$R�n*�XKA�Q�Hny��䍍~�a}R���U�@a3)==��=��Ǔ�hO8�) /I%n��M�FG�#Ϻ����J����H�%�a4
���'1��%��q5,ҪVZT��1O�L�Z��'��O��i�ME:^s*nZ��#��;���"-��៸NV�xh��W��lʁ�;�Ɍ|r#<%>QKc�W��p �D�.�e���
�tx�Ԫ 7b�t���M	��g�'�0�;�$�w0�#�Y�t��� 3��.S����'9'd����!pKp<9Uȍ[��\��C8
�p ��sX�̛���
��E�!	ߚZ~dJ"���I|�����ɬ���'R.	x���'#@B�T��Vy���n�����b���0=с�Rwl��'uȸKE�V�������d5���t���c�f��>���BF3;5H�~J�E��f5�e�|�|`
�*��'|a�"���,����=�F�A�eM JAXЙpnh��ہk�T�����Ig����Q� q↎�d���+gE��-�t���� 2g��Oh�RsO�a��a]�2���l�>����Y�|�p,(;���"i;5LI�щ�IG��	��ߩi3'ŊO�14	Ҥf$Nxrs
��v�R��  LhB�w' �j]w�>�/O�xs��F�!�b�!���A��J�p��	*���c��BGQ�O�|�'�%W�CSa�.3�$j�Ň1�\p���Q�d��	]�U��ͪ��m�A�4��$Y�Aq�M0T]�9�৫>ɖ��k삠�ř%]�>u��a#cS�9x�J@-,���`���2i܈���j`�';Tn��K�N��ix=E{��S;ϔ���Ƌ��*��	��r[<��'b^��������]8{O�����;N�ش�&T�n�B��h��Pό�� �]�*B@$�
ӓ'F|�#f�v����O+� A攜u��1a�g�^P���n t���[#�$"�a�4`���NZ)L|�4�V!���p��N��H2p�[�'���'�ųV.��K�	?	��=VT��+5�Z�j��"R�v�aA��2�(�c��~��g9m{谢�	W�)��0KQ�Ȁ������5޴�rp�'lJ�i���q���_��`rƮԼ�����Ȟ��S���P�%V�ɂ���iO�T(��dl@�m ��C(�4b�vtKG�bA`dP�-���A �"]vuIC�Ɏ���\�{�jŀVE�6�N�Z5��t��F,(�m���ܾu���D�[��c>u3�"ªN���1��KFt8��T3�"��`�(LO:�KG2�*��Ͼ^�ٹ"�)
=�q3��j����a��Kr�Z�%\�(����
���?�ST�@�x�Ja�ŋ�G;�尅B���Ta��$@	l��y�`�\6P	��
�|�5BFI�V�;�DM�M�\�aΈ�����l�s	T��&��!PYf��;9}�%[�L"U���ps D��~�B5�H�F��(S�2���~B�j=F�`���<��$>�3�$K1YP����N5U����C��)$fl�Њ�k�h$�#���[TN���O-���V�~Bz#?��J��S���S����E[s�G�	+D˓.�
��a�5>%����́$hr�D���
7FRys�_�/�p]���I�t٠qa�'i��] Y����̶'�	ÈV �*���|XHmxb�QL��%��|"��YX�$�Z ��� Z�X"Q(0�� �g(FE��)����(!��8���X��Om�}(nǩ��t�q��+�����ȷ ��+��B�?����d�E��u���=g�!���?�I4s�|D1�`����Y�$hMp�F�'�"���A�zܓ�zY�&lU-(�E0��$Kڎ���(�0f�HY'�i��A����:
�a�Ɛ�52����	�4�N�i!L>/�:i�G�V��c�������Rq9S�� )8<u颭�?����É+�y���L�$@\�:���-�F�*�'?X�H�JB�}(���#w�� #�ݙtj��ہ.�_��sQ� B�X�J�BR�=���'@�.��E9��DC!6j2����	9}!��	�t��ʆ���J!r#I�)���J��ɛ��<��2w�Ś��Ris�.�|��})��-}��� �j)�C�\������)��=y�O�.cv�:�mY�!�����Ӟ|�WJ�M\l�d G�^�l��?/p������r���6.2�z0�;r��5YC�$l`�O��S6�28q�B��,t.H���lA,E��+��'u�1#ܺ0U�eҲ�4@���@Uo0�t�!�{�$�t��w4���[��Rк1B�<!W��vK�,0u
�)�;c$�pQ>qw�̍
�%�' e�B�#�E��!�'��i"P�܍!)ޥj�F� /�P!��d�b�H���U�F*T����u��H��{���*U��:�p�d���qO�ɲLA�0�5��I�%��㐠Y=���hFĊ��ȱ������mqrꌯ&Ĭ):��-�~�b��6�<1��ն�}x�AZsT�H�R�'���c�b�,>��$��jߤ�J�Oj�1S�
3b��p��s5<��C�64����ٮj�~2 �V�Eh^�2�ew��5�Q�ȏ���H� ����%V��>ט']z��9��E!kF1#�E?�lC�5�6@�U�I� Ј	���oJ�hQ7a$՚牸0�l�S�T� ��'��}"�G��x��F-���I�{	<��@f��0@m���Na߬U"5�ѨV��	{Ʉ|�R�'%L����Y0��&تG	L!*�D&)��	LD\3e�	f&�`cbʠ@h�	�ȓp�0���m2Am ���üU��ȓtnr�1���dM"p��*�U��̈́Ɠ��A�a��*d���v��TA�iq����1YP����D.8�v]�_�Ď�N��,�Vf� Eg����ǀ���yRb�e'.���È�_�i�vLW�'�����D$�~��㋵-db�R�a_��A�}|>X�@B_���O��ʰ��J��183$'LM8�Đ|2 7l�8����Lk� � ���~�ȉ�y�C�6��(s��Yo��2�/
�kQI�b��x{u#W�,hE�󣇏X�,��j��w��ɆnAz�z����'oyyq+�<��i2�Ay�0�@a����B,� �=5|�2O\��P*��kp�it�6�̄ �e��dq�>1��6,��� �<<���]s�Ȁ��s@R94mW�$͊e����2
����I��
d����?���;,��!�a�&�;A�����/��D[�J&��P�:N�P��]�U�.�>���B�.dr�`e�����p�|b��sc��tE�J��+f��)"�L��'�z��(K�EnT�s�߻B�u���G�j2Ԇ�ɜd]c�&� 0�j�1�B�&Ϧ�K�mv�	Ǡ�:��lp��D��m�Lͻ���	�V�=B���M8w*�ɄƓi�!@bFH_�88J�(��1���
��R�>!R�@�̜�~>�pr��A"!�r4��'�:��6�9g(�����o��-��G�����"/z�,�t�ө.�9yp��K�`\
�M�)"�1��G�x���օP��U�&�_0��8G}b-:7����eD�[�Z��k\=�~r��c�݋Ѯ�'c��������F�V=�!�!�e+��m��㇁#�p)�6��d
�_����'�����O���e�ȡI>&�y1��9�y�M���q��_N�W�47#��@�瞟?xB�ДDֱh�88Db,a�8Xx�}CHN���aKC2YG�<�T� i�Ɏ6
V8�"e�7}��u�Z�_�
�d�s�� ޔ�s�M�:/z ��0�p?���1|��bP��b��sˊ~����:@���d&�~����C�]q�4,D6q��֧�4E��JI;g�Ҍ9����� �?�$���3&,̚����
��	 3M�N�'#�t{�!F���X�R��4ж��6�'�b�9�B�5O�L�Y��]h�O@ع�b�E��@QA�P'{j�����{��|D}��4U�
t������y'͘g�^=��C�=�~���J�z�P�\��XC��5���?��� z�.�!ݸ'8)hb/�QI:���k�,I>��+Z,���fv�`��Ch}�OJ���$�%3&��)�-�	��,��ɒ��\3g�>Y�v�}B��)s���ɐ���E��'Ѡ�hR�EJ�pI�!^V� A
�f�ZU�@��	�ⴗ��T�=|R&D�њ~2��b��p� ��6�JjT1Yb��S�X]�B]X�.�����ďʈO�q��oS;G*>�) k�m8RE˳��>Q�	^!8Ci��*B�-�駢�O��Y8S��+�������<Ӻ`������ME|b�8z�����oJ7l�w�T�T`H�cN�I�����CV�e�'��s#��`�J�OP�p%�� GJ��G�I�P�V@k���M��AL�,�*�OL��I\�lC*U�b�V1���P����� v�1�!��^6nP�%ǂ�Bk. رh�,s�qO��[�O��-�~��u��y��Xw	�n?�B)T�-4� @�3"�>�3�`�=nB�F�/2��9!��Z}�O���
���o_T�' ѐ@
��ÓB���R%�L�T�rLm"�6yyPL�?*d���BE�i�� G}�I�H�!�  �}�醍� ����:"� !��٠��S�iX��Ƀ�]:�CṔLh.]qB@:+<�8ԭCY�'�0��p�(Ai �λo�qp ۝9J�ɁC�G�,���⠟��Ub\.\j9yc�W�,O8{g�ij�p`���rg�����M	'`��h����z&��R�Ȝ�⧏3w��An�~"��V6��EN��p.�S�F��d0�"����M��Ɍ�Pd搑� �+FD��G���<yW�PU���1�@Q��,��)P�7�
�S���C��(��� ��O�vI��\�=��$o>�K��]:б�֡�Q��\R�����M+G�v_:u�6�N��VQ��[�'Q���rl��3M:y�A��*��d����y�G��O���v�Ox�2׬�|���XU�����Fd��ı$A�.}=���Q��
jjn���H�$oh�M&t����R˛���&>P�a@�GǪJu<�S��Yn≞u՛fGɲ&9��Sd.A�.'�m�&��_9^�q�f���x�C�A�2�c�IK�P<��bS�?d%K*��$�m!�6-�(�R0�¬�����A�%T�_����D�l��Q�@T,�h*�E�o�ay򧈑$��I�R��r_�q���}e|�kq T�S�����%��vX��UƇޟ�:1f�?ےi�� ��Q��B��/��`B/KQep�� �/�V�(�J� �I
��Ё��*P8����B��2� �J��sb�ܺ�Q�Cg*�i�!�k؟�zp��Xu͕
	.90���Gg�h�)���ܩ��4'f��M�\q��R��~��z�6�^�HX��X�B��ɶ�mH<�n̑j�E���*~�ؔ�6U�F�t�X�~�ܖl�6�k�O`����ge�e�(OF��rOEUz�����HJ&5��"OrP�'�nB���o�9�H���d�B��I�	Ǔ$�4�
�>`���iV!}i����R�p�6��/2
�{ԫ�^
���/���x�h�[�LYW� �?$XP����y�-�"s�x����A�3Vis�-�y2��&��|�uG1���S�ʎ�y"�%p�ph���$^T]�C 6�y2�Ɲ9���Kw���\���)�A��y2㘶U�D��4�SND��(R���y���o��C%&ӏ2��T C���y�dk'�e�q���{ܔ� EH��yb�ҍ~�VĘ�b�=3�yx4��y�סF�z���[!=��`eO#�ybN��eA�5���e����⅊�y��c���
��IK�'��y"�W��\�v�+.�xR򁔟�y���&��,:�ƃ�'����1�y��F��9�rc��vA*@H�"�(�ylr�l�4�` ����
��y֡[,�x*UmX �6<�	��y#]�6hx}s�+�-@D���yr�](48�������:R�D��y���%F�LؓdD(劜9M���ybi9N_|J�ޤ?�hFj	�y�)�-BX0�)s�S�d@����A��yRLJ�t�Ц^'m$$BB+�*�yR�X�D[�5�2϶b&��u�\��y��H1$M��'��|,��рۥ�y��Ο�R�������Z"-���y�Z4N�D�p�l��,2�%�UF�y"�A'xWu��K�0���*��y�	�;0H#�^+.~a��n���yr�7x�Z�q�9L��yQ���y�%�1<���L�6�Գ�yBnՏ�س����7V��ʀ��yBl?X��J �F��,9pK�;�y��P' ����Av�8أ����y��[	 �U�H�7扰�F��'��XI!H�\�� !B��`ʮ��K>A�(ڷ`sHсъUg?��@���Z�<�wb��]pa��x�(�h�R�<�����N��pq�$�)��� �*�L�<� ��� �&%"���4�X�Ět��"O���S�X=��ex@��[�h�"O���']/eҤQh�Dg� ��"O�yXwI�$}�����i���$"Oz��o� I���Ã�I�(�p��"O�P6��^�WQ�v��"O���q�@I''"m��v"Ot����!��z��]/f��"OJ����~I��S��Z:(���@�"O��鑭�%t2Z���i�/#Zj�@"O�	i��̴�0d)��P?�e��"Oj�(&!�!a�D|s��w^���"O�Y�X�}�"����@�"OPTy#��E-$q!��J�䀡�"O0����!����H�#H��us�"O�8Ó�89.ԲSB���ȑ�"O�\:���qP6��A�Ta���ɐ"Oӡ�Ir��W�U�S(D�"O �s���)���T��(R�jU"OBN��ul���-Hิ ""On��b�̹*b�	˵�  t�2m��"O�3Sf5-^���y��X�"ORi@-
U�a�!�9���"O:� E��krq�W'y)Q���/�yB�-(�f�#��I�+V�pY��G�y"jÃVe�x#�S)���1k�y���%�ذ�j�%��(�f;�yba$�4��/'���`Ǒ�y�/�q@`H�!���Uf� ���y�g�)d*��p���*J��XQ�ʉ�y2 �t"t�c�I$6�%#�h���y��͆noĨ)PDI�.z��{����y"�܏8��@̈)�L�c�^��y���ƥ��EA�=��R�O�9�ybjՔinh��BnJ��I����!�yR��2Bz�]S�d-�b�2����yR�A�W��t0B�|���7�Ԥ�y��$*��S�/L��x`mT%�yb�Ү�h�-T '���"����y�/P <ᄧ�(�̩iG��*�y�)��k��؃u@�� �H,�.,�y���c[�J��˒	�=�hY=�yB�M�at��j�|��T�2���yrW�~�V!J�@{N�%jr$B��y������H���T:z�t�H �y� x|,\��� <מ�K�ƺ�yR�]�ENU��O�,%��C�@_3�y2�H GF�xЅ�;!i�8� �O�y¬N�L�0��&ҕL	VYaD ��y���gl"$j"�%	���7�I?�y@�=L��0Y�n�6C�j��>�yB-_��� �B&��2�I'�H>�yR�Ie��Q�6��7�4CJ�y����S�@$bv/Ɋ6��;#��1�y�#�En��֌�86A*Ȃܮ�y��� �|Պ��6 �)��� �y�F�gӤ��5S�f��Q�4�y���8b�`�2�.�l�XUĕ�y�N�}�4�a6g��#V��� .�y��Q�:#b�hY�-��:�ȅ��yBeСi.�dy3mF1*V.@Yƌ͍�yr#��7=�0�4� vFX�����yb�O�ލb�	�h������ybe ;a�HUЂɟ�`) ��I��y
� D���E�Hd.�����Q1�7"O��Y�E�7?�[�Òt �p�"Ot�q�+�V�`�E�ܡK��B"O� Ӯ�8�Ȑ�&��-rS<Pp�"ONy���/L��aQ�i��x�4"O8��Q	�)i�햪<���"O�U�!
ǬYN�k�a(m칚�O���
g��C$D[�>�8��Z�)�!�X Y� ��g��84N�b.a�!�dU	*�@�-
F�S�C�c�!��9�|���Ȗb|E�wNR<`�!��_�"<P��AO�(���!�d�.;%>03Rj���l��� !��L21â��4�[0�Dq%�(2!�䄕:�z���Ӳ7�0]��(!��[>n�����⊊R�\Mp�� �h�!����5�'�P�0��u�s��L�!�˛f��Z���-\Vҙ#o1	N!�䝿,ʤ9!�Cr�I#H9!�d�b�ڥ���D��f'N�@ȡ�]�q��b��<!|�:�A�/�yB��~{��ka@�,7�ȁ�e&�y�NFp}���$�#&Ǌ�IwAG=�ybE�b
��Ԩ�"Da��,�<�y�)ģ_l1bA��,���Kµ�y��6h��3"Ƈv���L���ybgV�Kv���Dop@U�4����y�f�~��Q�,@{6��j�D(�y  ��y��T�e�r9؅Ꝫ�y2dA�t_T�z�ś�`�1�D���y�爄,V&�@6�J�^��mY����yb������G�ύ�P�u���yr%P>b(�j�"\{�Q
�H��yb�)0P&E���${���R�)Ȳ�y�IA�I��1@��h��9�jV�y2�ټ*
��d�7UXvI� 	�/�y,&!���($�G�b�1�I���y�m��:��@�d �Db�c3C��yR��7G�	H�a��S�dC� ߷�y�4#��l��o�y�@x�f���yb͍�jv�jJU�	���`�	�y�χ l��(�2�R�{��s�d�9�y���#Z�� �M�;pr�P�@��yRe=1><E�wD�.a��< �Ŭ�y2���c�Ƒ�d�]F}�	�=�y2/�h�.!���?R��1J7�ü�y@?4���#�ϭJm�i�e��y�B�X�d��	G&>mLk��[��y�(~>f�(��Z7��h���8�y2(F�1R�!��ƥ#�}�偈	�y�+�+���a�C�t��b��"�y�K��%¼�
�GG}�4E��N%�y� ݩu�H���n���H��]2�ybo�d#����!`
29���ڱ�y«��7��(�qA\�]�T��J��y�$ڽ=��t.���T�bGaH��y`�1�Ѓ�Ÿ}F&)��i�y��]�3�l�Z#�՞o6ܔ�v&��y���,`��h[�!ϫf��j�f1�y2.�;?y�sl�f��J ���y�n�r]�"�	\ ������ �y�/�I�N�ʀm�=+E�ܒt�D��yR'[>?M�0��Z�M:�xKD��,�yBiW;Y����6BE&JT� �)��y
� j�c����4jp�P'k�J)&"O*��7�	���`.
%�hl��"O��7#�&��`'`����"O.9��I�j�l���4����"O�$�0*O#�J8�
�8O^�+"O8�i�8e{~,�Ah3e�a�"O�:s�މ?���GŰT2�]zS"O��Д.B�k�\�!6)�b "O �i5C� OH�i��萙N8��"O�h3O��_,N�Y'��)#>Y2�"O�s��̋Oi���F�u�m�f"O��IG�:|���Pe�#?�H��"O�qy5�N��V8���_P025Æ"O��i0�F�V�I����&�d�)"O(d��Nr����&?�^y�"OFQ)�\
kx����Dv~\ S"O4<��d��U�1 ߏ*LD��T"O*q�Q�p��+"�
8֠k""O<P��
A&�|��n�#l5��"O~��䮑12���@��1!$���"O�����_�Oa"�2��L�'`xj�"OfIjV`��*�t\�V)_�D�$E"Ol�� �� Pw8���(�.Br����"O
Ua.^�\��Ss�(3Ȏd&"O�ՊhǼ�$	����
E�"OP�bHܨfEZ9ks��=BK�P��"Otx���4y�գ�-��|�R"O����ݱ�URa�?��<�U#�t�<��n�|���ʖ!l��Eb�`TF�<!�Y� ��Y1�R[�J�x�GC�<A��T�F���9E��ęA�<!EH°b�8|D�Ӆ]:p����M{�<V��6!���@��O?訅3�CH@�<!�'��H��y�g�H,��z�<�W�3b��`���Ln��m�Wg^w�<�u�:&^�d�GW�ت��h�<��)�2J��`��KC8[wJ1���|�<C�Z�=���-��l.�3�C�<��Z�[>"M��H�5~� R� @�<AFY0!S���S��1���,B�<��፟K�ށ�`g�(1'f�:���<�s��1uvm�3+_�;`����G�~�<�e�E�9��)c��t��Ab���w�<�c*4x�9�d�170\ɰ��g�<�g�JZ�u���
��ρJ�<�Un�$`5�Ȇ%�M�F]�Ļ�ȓ#Xd-�$��%U��i�
�3�DQ�ȓs�԰�K��bHh�SHZ��32HU�
�U�X��UCDTP�T��Z���C�,�:���
�g�Q�^q��'kXś ��8Ft�3��kla�ȓ"��H� FѠ��Q!��)D.����I�4�a�[�q�dD� ���fr���|��!2KH�j��m��f;ޔ�ȓ+��4���C5R�)�aV�p~Ʉȓ;�21�3���+�a�v�ġ������.q22`��*d��8a��Ը9��,^������p���p�g��;��e�ȓv׶�$J��o^J��b��3\X4��?D���w�0��G���Y��|�ȓz�R � �'�.H&	YH����c�8��F�}t��K)�r��ȓN�q�\zq$��`�LOX��I�����Ɯ[���P5I&��T��S�? �mѓ/تfѮ��H5��Q[�"O��萄M�	��]��W�T�PL{w"OzWF��)�s&<8x%Â"O�Żֆ?�
�)u�4Re։��"O6=9�"?B@�0!���%b�1!�"O°��AJ6y4�aA��~NZ)R4"O쉴NA�sg����5p>>��"O>��e�H�69.�1��f7���"O��u�*C��X�*�4!x�"O�E�LH�+�%1ɴ�yR$~�<	����0��	����!d�q���P�<p)�>�2�X���d�:���(LP�<	��@�M�.���ě@�LA��MJ�<q��� BT��sS�/�`����<䆋"LdIƨG?Dv��y�<9��ɗ��
if���D�u�<YDɄ�j��D
� ���4 �g�<�'��t�ܽ�`�_.� 0y�
K^�<�ׄT�����&[�ELba92B\�<��+�-IAf�+��+
ĸb�jBV�<q��G$?m@@Q��[�+y�T �{�<)3�K���P�	�	)�Ă{�<��k�/~��1��v�����[}�<Ar���9�TMJ�H/� I�Տx�<i&��24"�,��ȇ.G\��7��]�<ib@�B��uB�F�(�8��B Z�<A"H5e/0���.
�r"5�Q.�a�<�������H#J�P�x�_#+K!�ߢ~(a�j�#.��PTi�-!�D�;��I0*���a�Y�*+!�D��}��I�  E��"���!o!�� [� ��@hU�L��S�'�zE!�ė \��C���5� ԣ�'�4�!�T�!#�@�c��H�%F�$p!��,��X��l[I��s��iJ!��Ʋg)n��L�UGRT�!�L1!�$H*_�TU���F
. =��ܳW!�C�<���l_	t�y��ܽ_!�S	'���A��bb����2�!�$)c��g�6 o����Ј�!�	>��Hp���0��]��d��uo!�@�>=���!7BBu� �����'� �������J��aE9*R@)�ȓ��D���ܖK�$�򤑳K"B��6��X�A�E%�8H���Z�S�̩�ȓ��l[�I9^�M�6�^![��ȓ,�b�!r���
~\��o\":�(l�ȓC��Ҳ"Y$3�h��E�ot"���A2��D���:�D�T�xQ�ȓar�!���/E�H��N�*��X�ȓ<�*EX�(�j�m�6.���4�ȓ_H�!�FH�[�j�Z�ҍ=&ȕ��>�x�î�,LʹU��$Y�\�6���K�4�yD�].WdT��`����Ѕ�Ab|b6Aϫ7e�i�@D�?�Dp��>ed|��-�x�:isP�ӫm�Ɇȓ$��p#��Xq��(��5����z��1��5���S������ȓU�����#D�`sa�8T�6<�ȓ)��4�&�q�~=��M�����r��Pt��c�fE���7S��`��b\r��f�4B��[��I�ҝ��C�8K��
Nt���TgH�v�}�ȓ��9�V�`Dl�0�+KU�>x��S�? �9IF@�*&��5��K۸P�$K�"O^8ăH.J+ܜc ʇ41�$"Ot�	�AC�5�4���\4R���+�"O���s�+��{%��H�l	��"O�p���ЫK��kN.b�Fqc�"O^	1�	Pu����������"O4�F�%I	���4$�tuX	� "OĀBE�n�@H#��ǌLA($s"O(T�mV#V�4|�@��X^����"O�$���"���ݢ{���"Od������h����6�L`"O���AF�<���q�MNb|��I�"O�i�agJ�w�� Eʃ�X�(�"OjT���0r����R+�4u����"OXeD�>����ʁ��|��"O��wE�H����`[�;Y8��"O�y� 0V�zR�^9z���`r"Ox�Jnd�����;Uĺ�P�"O�-���HIً�(m�&\0Q"O��蝅9�\LҢ�E�Xx�"O��ʋ�9��䫳�70|�@�A"O����ĝ$�T�d�<4�Ơ3"O6	�l@ �.͛�� [ ��W"O�1;��^�n-*2��a�"OTeiԏ�:�>[D,��l�d��"O&8j"��&��ia*
)QՆ��U"O�����K��̹�GJ�r�����"Oz�q��I��мK%*�*�z�H�"O�l ��ث(����)O##+HKb"O|��S�C`�d��[�18E�"O�-�UG)f�@5�VE,X�"OlSEV�<!NA@��$�T���"O&%�概�+\��K���I�N���"O Tju�X,{EHҳb爬Ie"O|1�0N���c����Mn�"O��
���9C^���&I<^�xɁ�"O���nO���q�Hc����"O@S�a�	bqNC'�$.g���"O���E��I��U[s	��nT���"O̓�
M� X�ĴZhT��e"O���2�+:�Ç� 6��Q�"O.P��Y�cޘ	����V�`�#"ON���.(L�:2t��S��0BS"OTxk@��>-�rtSD@؃��"O��%���!� [v��4�6�c�"O c� ZEg6��1.C ��ejt"O��YC�Vi�������%^�
��"O�m���`݌\��K8yS�3"O�53�").�`+�%�*.�Z�"ON%��Jյ$N���`
J?X؀"O�+5�ʒĆ�#���5��j2"O`�L2;��ac��ՓK�l�4"OVM�p"��^��%���Й�"O^�0h�O�BqK��(py��"O��`+��}���6�\Uz�"O�T$ſvD6���ខ
�t�"ON��g�Z7.���7`�V��"O|��C�) � �B�Pf��Q%"O��;��SC�~Rv�tW���r"O�m� �T�]�̴gD�6u�[�"O*�j�k�����P1_
����"O�ahB� �	r@H	���`"O��z��K��75�%[�"O��h�1��=[bB7m�����"O� ��±�1X�H1�������"O�u��˝F���А���i�"O�yG#
�S�()@怳1  (�U"On�۳M�%?�`��r*���y�t"O:�Q�]�sD�}����j�|4Y�"O�@ӄj]�2 �8a�W
y�6�h�"O^ՁP��:|�Ԍ!����;����"O�86��'������Z�\2jy��"O�� �Q�[�-�3dE%D|Ƞ"OP�;a-D>hH�i6�̈́E�,7"O����.ٽS�z$0�]	*t�"OD�3���ة� {밀�r"O>��&�N�3��� F���E"OZ0Eg�>���[�E�  "O��I�0�D��,�̘h�"O��#Rb��;[����M�ܜ�
P"O��5!:*�N�#U��66���u"O�"K�v$b�j��pਗ"O�Q�ҋھߘ� TiOQ�t1Zf"O�	��/R����
� lھ	R�"O|A��lԱ?�l����N���9@"Oz�B�ꊴi����M�I��"O�P3�	>V(��c��t�B-�V"O���6l�\��TRaI7Pˎ9�s"O4�"�B�5 ��p:��K�r��"O� G/ߴ;7p�Rt�S�S���r "O�|kPƃ,ap���h� ��=��"O�䁡f��@o|I��ǅ�o�.$�v"O�RF�_��� }I�d"O���`Hʥ;�N�*e�7af	�"O��MG+=���t&\�$F�tr"O(!FFQ�yJ�d�c�/;?~0�u"Ǒ	���t|�;�f�Q����"OjěH��u攵�!�JG�&ݒ�"O��z�)��H2�d�t'�T��@�P"O ��w)��3(<3q$�3��l�A"O��U��[P�LX�lE:~���"O e �Ǝ�l4���
�$8@ѪR"O�h��c
2� xyfl�=O�X;$"OF4��J�v��ᒥ��6: ���"O�x�����ٺ�p�� -ġ�"O���Ɓ7SH�8aP�ҍPfL)"O4��&�ލ#��h
��Ĩ'�T���"O8A	ᚎ?��M3cֆ ��y�`"O,� �(^\��z4�̓[fE�"O�(�!o�#:�zp�R�1X�٨�"O�x��З^��帆)C$I��"O�@�����>�nP����/\6d���"OZ|��>�t��֊J�s)J�Bu"O(�#���
!�
�<( +�"O�D�*!���w�ŽQby�"O0)�W�P,y����AM� n�w"O���SD�Ae�b�JU�]s�"ON�u�M�+bt��� .U�Q�`"O��c�D>vn*���S\6���6"O�I'E;���y� �G,��x�"O���T��G����5*�$�uyW"OL<;ס����5N]�a�A2�"O�y����`����q� 7^&a�@"O:E�Ԭ�� 
�A A��FwRI#�"O���@$@�l"$ q�	�0qp.�{1"O04S�F� ".��ֈ�SXH,�4"O"E�I�
Jo��r ('���X�"O.�����$S�����$p�"O� zH��NZ�y��|B�Z){��#�"O��{���,M�P7g]5����c"O|x��A(Ҥ �6�Tj��E�"O������20S��HA�F�Dm$=HW"O��0��C�4��F���2����	ן8K��������'���^?���eԐv�A��4"�*d�C�	��9���?)�4a\)0�O� .�#�-+�JC�u�����W�g�
ْ4�# �0ps W.�(O�U�ƥ[2P�J	�g�(�	��� 7׮���НW
���ug^�t��D�RD�+�`ex��O 8�x�O��ʀ�'g"6-�P�S禵A�-	�8�pu&L$iҨ�;��P��?щ���'�IJQb\�(���Ȳ�&T�N�08��D�i��4�MS$�.OT�q*�8"h<��S�s?ɐʛ�B��V�'�W>;6)	ٟ��IȦA)ڝ�<-�3�-s'�Hjf&�|�pe@s�	�ɛ��,OV�pD=�╠+���	�m2�N16�y��fף��E��`h��dX��"|�4LS� %{T��WI�[(� ���\c�D�
`ȟ(
w,+b��}>,�4\���?�MӡQ�����禁��h�BS:�ƨdWv}��+�O˸��$�ע3	�s��"C"��#I/ʓD���*y���?��{WDT����-.!Ny"6�ĸ{�I���'��慲L��7�'���'y��e�I����{q�}�i!�+S�f���	pe�%C��i�����a%��&6��s��}�v�@[w�'s�s4-���8����P	RT0�#2���u��,�C�~/�����!��ɕ�Cx&8nQ��6v���H�sP��'�!b0I��/]/���I�M�J�~�'"�'E�&��,O�(�#�`_�_d�$�d?0R8��?���?���$Ϯ~�d�����tB21 �N/Z^��2�4H���',�6�O�����ʧ6*�I(U/�=�����)��'�^�����?����?����?����?�GK��y�8�ЯX�9�ur�m�x���J����}#pT��=P����\Z}��!��D�������z��RG�G*{�|с���D��F
B*C��6MU4��T����1_��1�.:?�0�	�xo y�Z�P@�s32�;!�}&��A�x��'���T>��'��F�j��Ў�
�j�f�8}R�'���D��|�x�3�XS�2���'�7�Φ��'̈�&.p�h��OH�'q��bp@>}:mIu�H"P� |�m� �'�iȝ��Am�[��T���#㪥�g�+=�2e�#�\�.��PAg��s��9���>ʓi�p��1���@F��I�.��pP6=�%#
r��1�*cȲ��7"-ʓy"Ҙ��'�M��i��^?��l߮�bj� .5��{ d�>�?����S��?���I$��#a�,���C��u8����4AÛ6�i�]����iu���D��i��@?A�!o08A���?).��0q3$�O��d}��q`�
�@f^�!��L�7�rP��!\�o�p8�g�M.�xBɊ蟔��
"t	���O�°��:d[(=6����D�l}��i�2�
TA�e��j��P6ޔy��/g8��enͨ�Ri˙�5��O �QG�^\v�UH5�M��ȟ�rش9��'y?7-�V���k��R�6=���'r����O�ʓ�hO��0�RUٗl:X�,9�Ǡ̿Lԣ<P�i�l7�?�$l�r�ݭhO�2"�C�<=�BL]% qX��J>1�=�� �  @�?�	uL@h`We����=E`�4   �5A���W�HH}�� )�?I�i��"=��O���0@�/&H`������n�3����������F��/$�A���5)�h�iB�O$�M�4�iuɧ���O��	�b@@��F.�,{a��f���]ҪMB��J���	��D�����h�"�ퟠ�	̟H* HԦu�&��'A����$��us����ѠL���z��7O�(��d�CεGy�ѧ~�f��x�ڨY�(�&,x�xlA�����vj��o���сBu��6:�I�<���
�ȲY���3;p�c�90�}*�,R�E�	Ky�'��'9�	�xn�$\�:�3r.PR�4���H�b�LL�����?��!�<!:N��Z�|�>�@ �� <
��g�Jo�˟ݴg��� A�i�2�'�;p�0�K"��-e�(4�P)Q f��ag��#"	��'�bV+Fz�Av���	�g���y�d��B�~8k��U����,P�3s�=�G/*ʓT�f�j�)[�*�MiG*��M3EIS]�lq�m
	UBl��6'��#��d�a��+��QT#ۣ��D�8�'xl��6�k͍
c�_�E��#".ڢI�x��'E�O>��'iD̡�o�(}���f�J�Lߤ��/:��%�N6MRxRM!`��">�PT��֒�'~@e�n�.�D�OX�'z�����?��4.�)� /�D�<��a�һ]|�s�Ð=���XOM�*n���G�=H`��C̜s���?��1z8H�����6`:b E��k3$�mڽD5V��D��xLHC`눹�0�;DCI�^q�klǧ�~�ICM�:~n���M�g�v�ӏ�?!��i+h6��O0#~nX�֔aG�Θ�K�c���	ß���v؞@��K"h}� �Q�L���
)�T��jӖ�O\��Mdݩu�Y�Q����߬�z�	�f��?i��XF�9�L��?1���?	����n�OX6�^�bZ�mx�
�G ���0K6}�ɜ�>ę���7�敲��h�B�C} ��O� l�KdM�U(�	Pb���-�4.�T��	��Y�+B���n\�tδ$�'tG^�(��9���:�h,"cS�] ��#�Ό�#���j������ҟ�)�4|�4�gy��'���4���"IT�g�����ֹh��؋���O8m�堀C��}���_%B?(㡈��M�v�iX�'x�(��O��')kl26Z �  �  �O�Mb B�x��*2�۲4�5Sw���M�i��'�@�v�O(�'�klњcZ �  ����t�ro/�j�[�����Xڴ��G�0x��'���5d�Z |  �O��'5k���Jd �  ��=t����G�q� � �'��f�	~6���Qיf#D��'7���l9�P�ޑ
�L��'��p9�A֙9 ���v��Y�Z��'�����֏tj�b�+�&<�b�'AT�h��H��B�r6��hp�'�n�hF_�- �Q�H�)^��'ڄ�J֪O�(q�K~w��:�'�"�P�N�$�>�H�
oݴa+�'�d�:��(�YP��5m
���'8�E��(G�F�H�w�ř1�9�'� ��!I\�	��D�w���+�4!��'�.�;b��%Z߀�jg�ڍ$I�p#�'`��r0���Ag&�_tEy
�'����RG ����'�
�̨�	�'Y��7�N�$��ؙ7B��&�k	�'ɢ\i6D^�YG~А�i���Rh��'��e��ʶt"�X�i	4"p�p�'e����+z��)��l%S���
�'#���uÜ2Dv��UC�N*\�B��� �TH+YV���ƨ��I��]I�"OPD����\�3���K�"0#�"OT�I�aA�&�3soԽ.K����"O�	5�U1@/��CO[T7��5"O�A!���<�X܁ �@78�A$"O��;a��Y����TMq�xA��"Oܱ�"[z�V8y���f�"}�"O
�Ӡ"	�f�As�fI��
i�$"Oޅ�e�h늩9P�Ȝ2��XS�"OԠ��&	4���g��+׊���"O�#'��,ͰA���30��(b"O�(���6q�l󢋚�$ʀ��"O�1 �lϳH
���	]4���`"OA؅���9�h�3�'_(�J�;�"O�)���4)�|0��H.2֌:"OR�k%,�: m���+�; v��҅"O@�x��-�����J�#!���F"OLP����N�ƤXw,�(FԖ��"O��!D[�pfԬ�s�1`� 1@�"OԱ�A�R�aFi�,� �����"O�%@/ɸ;��bA�ϴ	h�"O޹I�a٭X��)��%&����"O�er��$ lu��0Z����"O�1�Ņ�4<D骥�J(����"O|���͞�0Yस���\� ��w"OB�Y�2H�9�V)Nn�lK�"O��G�K�*�N,ZbHȳ+c�\"O*�	��ۉ;�
�[G�+�A��'��ţ�2z�$��BC^��)�'w��ˑꞹ?�b�҅�l�6"O�bЎ�}�yIդO�h)�X��PyRk_84Nfy�T���X2@XA�	]�<y�)_�eB�=��-\#p�@��D�<�w���nq��! �̛�jAH�<� ��<04����'T�f,�B�<u��Ά(ŏ �\�Ӄ�|�<I�]ebQ�fBL�F+%��!�$�|�� �,Z�I�~Y ���o�!���_U�əq �!D��E!Z!"��^ dܴ�?�޴I�Ӡ$}���I埜m�La����*:B1h�����-H�S$�
ՠ1�T2�()co�D87͘2U���?!��e(P�����PЀ �V�v��-n��"�� x�Q�C���EG��'٩eK�q�RG�0?���s�a��j]8~]��a2ń�"/�M�4�'�҅��ZB��Ϻ<��s��M+��T������ ��W�[�O�W?q����<�E�O�xA�DG?��H��� e]tԉ��"�MC»i*�'I����	3�,;L�h%��� $Eΐ��4�?��BdZ棆��?a��?��N@�.�O7Mˁ��(q0k�L@~�C���w��P�-G��(��g�G dKv�M��?-᢭ΗL)��O�����V��a@O(��	r���+���g�ٟPq���(���?l�� ���|NE�u�Tb@��
�a� ����*9noӞHEzbU���� �v+�	i��7,�Ѕ2AE6�~[Q?��G��>_ ��aq�F�m�ukcԙ��ig�J�O����j˓~��`��&�&��b ߘH�LDzf�V��M����?���?��'���?Y���?q���M�����(tTJp���P4��i� J+M� ��e�24I	%$G&{r���N+C}���]��T�F�\�d�j+G�kJ�e�«؃q����t�Z�ծHo�j��*Ӯ��	c�e�B-����f<u��Ij��[��M����OF�d�O
ʓ�?�ش_?n�p�I�9Nq-)�J���]��'�a¯�?W ���-m:%c�M���d禵sڴ�?%�i�� ���r�����O���w�:�� Ѩr_��#Y�ȺQb�{�B,��n�O����O��ɚ��9oڨEH|��41U0ɪ"��[V��ɜY�m�U );<��Gy�&%g5��c��k��m�v�i���7��Cx���KY�tr:�A��V<J�*2$K�(�z�)D���U�O��$v��Ҧ�2��C9_����L��o��I#��֭�?���	�>pbG5t��Z�M�0Z��,X�
�a8��ݴRě&�i[�bu�t�L6���h�@�:�'��}��e{�,��O�˧�b����?�ܴNnȹi��Q�`��:�
�.5/p����!=��;�ǵuΠ�+��t`�㜯%a��?��1Fd|�u ܰh��]�A"� w`�ylZ_��2��%p;�D�*���g����\� ^��! �1���%��v��Ͱ �i> ��f��J{�`�D$�禹Br#S82И�acɬCe�u�����4�	Ɵ���I�~7�=�C�K�7�x��	�:	5��<���i�x6m.��A=a��ݼa�0j"G�/|'r�0'�J �6�K���?��k "NrPH���?i��?������i��miA�A,�X��C��DĄܨ�Q˟d�Pj�Epܽ�˅�*��i�	�;ˆ��0�d��f�2IUPo���[�/�h$��':�tY蕀� y���@Yl0� ~��<K g��N�|��w'�!�6샳,�xQ2c�5�d uB�O00����OZil�����<����ą�nu�qyC'��$�z!e��\�D{���'�Z�굄�+$�0� j�7�Rt�&O��I��4���-=�*'�|�1�x�� @�?*|�!��;�.Y��G�+F$\ �H<����i��'&��Οh%�0R2!   �*;6e���<a���Y>"�EQ�Q(�j2u�=>۸�+"�نS�"��Bj�`�2'i� WvJ��$��d}�$q�*lZ�p�O�XbL�R�|I`wʊ:=�Y���O���8���O�Y�gG	>3A�p�0md�<X0�'J�7M��em��,MT{�"!e6�Ia���JN��'�l��&�'�'ԱO,��d�  ��$��aZ?˓�?���M�bO�K����I��SJ�[#��k�<�3by�$GND�jQHPN� >!�7MPӦ�%��� B��?�'�D�1�d� @�?Lk�A�� �  �8��F,S��pǋ� �!�Љ/0fxA1�r�Ҝ��
_�p!�Z���8ao��d�M�V�1:�!��ѶH�ļ��_�� r�XZ9!�Hy*�౶d[�D��0�ǁԊ,!�E�,�.� 3'���3��*O<!��*��'�׫Xi��d�(6!�@�P]0���#s^ls�!򤒍{�)@�gKO�ѳٷ�!���:�~thw+�	33�3�ˁ�!�d�?ha(L
�����6�<�!�Z�w��)q��$]�Ԕ����r�!�ğ�Y�� -�)8H
��@"s�!�X�Z�ųC-!Z��AW�,!�B���2���~��!��+C4!�D�%;���PaK*���em��!�DQ�wS�0�E��>՞���MϜ(�!�����zT�Ĳ��kWlR�F�!�$9!�J��g��|��Ja�6�!�$D�6��<	U!M�<v����!�-�!򤑾j�TdhC�ưW����@�"}!�%-�N- )�+:ԁ��!i!�$ŭ}D �3f��9{ �B�`G�I�!�Ē�Z=���HA0uZpYu��`�!�$�9b8A��o�xT)�b� �!�DLj^������Q�naxց*�!��d	N`��EF�>yR�!u�!��NlS&Hjף[�y��G�!�k��՘�O�"w�<�b�+]w!�dMt��*��:I��A�5�!�D'	��4���	16�Jy���Շy�1OH��$�6SQ����K��B��`��%�.tg!�]�;BL钔暆Xi�|qp��WV!�$�D��i"�G! m�	{`�ԴQC!��07@�����ύC(!��@. ��ԛf#ľSn�Yqu�Q;$ !���5M*��W�I{V��R#!��X&#�P�aK�h�D�w�L�|�!�Ԯ+}�P����@�p�(n�!��Ӕ�z��d��2Z��\[�kߥ�!�ăa�u���Vw6h�M
}�!�$ѫ�^e�YP`�e�� `�!�$�nX�y���\E���+&�!��њ@�:M�?;JJ������!�^�gk  r '�8[7t�&���^�!�d�F��Ȟ�7M��z�"1�!�ē���EJ�%I�ZJ��� b�G�!��3���qˊ�2�~��e��W!�4(�n�"NS�N�J�`��3!�� &���i�-[��Ӵ�H9%> |��"Ou9$�Ă:��M�M2!NP��"OD���G�>��a㩎�a:��"O�Y�g77��,��Ǡ~����"O:��W�ζ*14qҖL��B�ܻA"O}bp �+u���r���Tt�P%*Ov����*Q��Ybd�� 3��
�'r��҂�T>w��h�
��+�h�	�'�vihF�]?5|�i0�ͅ�j�9�'Ip��&J ����Aϩz�
�'��0�D��4�1;�b�7o�-�
�'���g|tN��D�?li�1j	�'��*ǎ�*�)��ȏ7WN�C�'e@�x�_�z/�X�-ě$�4T�'9�j��ڐfj.(��2%4�r�'eR- 񍕔[�j��$��
1r���'�䌱��'o�<!ĉSvR�8��'Z�%�? xq�3��=lȸ�'Kd��bܧ�Aq��dS6=��'��)c-�U]���!DXV��'���w�̸\�,šd��{���	�'�(�Q��W5�̵R�&�( L=�	�'c*q7�@�.}iD�ڄn�P��'������)��
��goT���'B����F�C5<÷-�`�D`�'�l�G�W���pwB�)Z�Q��'EŢpdE�i��Y��H Gj�P��'?� ��h�<@��u��A��
�'N�Ժp��8
�:��EF,;�ĕ�'J���q��(��e9�OC*-��a;�'&��{����h�#' �&r��|H�'� ��Eʵ0�h`Vi��R���'5�9g�'Pи(`��/<�1�'(�p0��߷?%����cͨe��'!0�+��MG�&�ʅϐV����
�'�z�;5�߯!fN��N�[�*��	�'��Ps��^) MX�M�8Md䬀�'B�<`6�<bW]*4� 9|� ��'�踈D,�^,Uc#&�t��(	�'�������@
��
#>�� �	�'t��-Ʈ,��yy���0?&mJ	�'��(�����&�@ѸwĹ�'���"dւ$���%m��J����'�*b�S�xh���,�84ƙ8�'=�K�H�dɎӢF�wo�$��',�e(wd���H`�"F�u����'��E�#&M�gd���B?\�0�'���C�^=$�F�����f���
�'ʼ9�3.�k~�i�I��X�h��
�'B��	���s$H��T�)M��
�'D|�[ᧀ�_���h��J�N�xm�	�'�|A�E�q}�u�nIT����	�'��Hah�F�D숷B��IǞ<�'��P١LYc,��7˃�>�r ��'{���fB9Ƞ����3m8@��'��AR���0}vdA���K)[ީ�
�'�BP
e��6.}���@6�1�	�'��'(ЗQ���5������'ǐ�����L(�9�Evvp�'���L�!gLX�B3O@�@�\��'��H��G:
a�R
X.=H ��''�����8m�!AS:$��Ĉ�'�\�'��*6,X{�O�N��]�
�'18�kCt<=	�%Y<Js���
��� 0PH�e����P�FJ�Uy�Mp�"O��C	�;��E��C�0-�@"O�8���w�T�y����t�E�"O܌�Fi�o�d�bG��envMP"O���+l�ĉB��$6`��"O�����,�%@�U�1b�"O�u�T��*�(�7X4P��0"G"O���!�Y*7�aq�D�!0,yd"O��BA�߱)��p��N��q�Ʊ�"O�z�U�W�L��H�|Z���"O���Ə�x<SR��>?�"��"Oh��A�-)!Hљb`��_�N�hR"O!Rbk҅_�����O�S��1T"O��#����iEnQ2�j��"OH�Q�@&��<M��h�"OL(��cG�5hܰ��k 9O�� G"Ox�䫟�c����+�r�vH�"O\�f(�	 �M��i�lR�g"O��R� �)Κ@iV�(UJ�h��"O �3e�GCM���Ǎ;R)
���"O�G�1E�RȢD�Ǣ4��C "Opز��Q�%{>�Zb-X�Fx�4��"OX���-+V��!P�^l�x"O�1�%t��D��e�2p�`)g"O���DJ�5�\I�
�`�e"OrI��нp[���!S�,�2��"O:��p���h��v������Yq"O|�ZW�I1n�(� a�=9|����"O`h�"� D/aÀƅa@��"O*��˹�ʖ/X�GA\��"O��@iתp�tTP�l�c/V];�"O=��N$��`��	:B����"O¥s����@�+!K-�p���"O�aв� lf�ԙ�Ú-(����5"O���E������z���"O���R�Zy��y�m�$V�d�"OL�AbM�^���9u,W+�V���"OnDHgB�)L��E�?+lN9j"Or@�jj�Ă�jQ�6a�|@�"O��%�P�%��Ѫ�*�Y]$Mʒ"O�vgܔ����.�*>(`f"O����[j��U���-7X�"O>�@���*�4���LEJ��#"O����j�h"H H&m:�)r"O�%��ѪyV���Fh�%l�X�"O���׀����VfY�*�h�"O���%%¤#������4 ���"OZi��D�Ӭ\zW��5��`*O4�0��v�����B��~Lx�'/<cC'ͣ	^xxӭ�z��a+
�'����TL�bd �2`P�\ db
�'���v��D�k��ŕCY���	�'P�@��Y,U�Ȇ�B�J��L�	�'�,<
Ӧ�b�f!q�S@�����'-*0@�뎑�pe�6(:ֈ9��'Ìep�`[�E`�ҍE�1��@�'pi�
#Hg^�S��+:����'0����CB�x�v�Wc�| C�'�b��ևW�F�F��&��i\f[�'
��K2���.�̙�e��8[�ؤ#�'}v�3C)*VK>�ĥE�QEB�B
�'{5=J'����
6DMZ	�	�'�x=0g&�\s�SP@^7H��0i
�'V��)#-S|���J\	,���C
��� 8�s$�  W�0��Ŧ*^Z���"O��2F�Z�)ke,w�F4�W"OJ��ԤʆjLĔ�e�ĤK:��3"O��aA�=>Ԣ}����1v ��8T"O�qʇ��':��2@GV�><���R"OԙCD�V�vZ��a�F�()�ISE"O����˅�E`*hA��]�R��"Oz)�bKTQ��F�,���S"O��)u�V��^<{��X�f���'"O���0$$~�>d�͜L��G"O �rt'�' o�=�m!��]C"O�xa�C$Af�(�lN!��5b"O���E�N%rT��FE��q�V8c�"O�D2�Ƒ�tϒ��IG.� tx�"Of�@��o4�6Ɓ�B�ܙj�"O@XX7�� 9�֐�'&�?ndR��"O���V��"`�Ft��gA.Maj�`�"O�@@Վכ'���W�"l��#�"Om��,������q3�AB�"OB0��n�"�(�j�CF�`�"O�`�&-E%x	��Q��]�J�p�� "O�8�Q&��QlXH���T��\�r"O0��7��-Ɲ��J���t�"O�M��l�4	�����g�xXs"O~��a�W݂�Se^  ��*OJ,ȷN	�l9 @Ac�2�0,j�'�j!�ڹ>p)�//U�����'�ԭ��G�
�ĜbƧ��R�xaY�'"����&̫e��I�mB�J�f��'�qoK�}�t�Y@��E�����'f�*R��*?O�i��V#C��p��'��4{q�>8�M����
�&q��'.4���Q�Mӈ�(5궼��'�J��W��7n$����O�h��'�\(��d���J��T��' �թ�gR�.���q#.^����'ɸ`��M�#&�(B�3W�rX`�'��À&�4z���i^�G�M:�'�TDh��6  ��s �?�4���'���sjU�,�2C�K�*J	
�'�\2��=&˔(#7�����'��xyG�׽x�X`xዎ'��ر	�'�D �vHE�aR)�%I��M΂�(	�'!�y�!G���F8�eKoC\Xr�'_��MF�S�E�<Zݼep�E]��y��!tp��ℍM5�Mʒ+M(��O���	TO8I`�ٶ}����U�P!�d
�~Oĝ!��e�\�h���B�C�A�<��>E���̉D�dDȦ ��+b؈��X��yB/�A*z����tD޵b3�^6��dI9D�n
�QFt-�Nׁu���#'D
�F��-��	�x̌\[vm"<�n�@�߾p
�gA��yR㐶i�&%�UI�J��R�O���O��R5�S'I����djL�e��1��'3��B�6-�Ep��O8���C�J	{zt�-��"}�&ʶP6����ߢ[Bit�<Y�C��R�q���Q�Xq�Ѥ�n����0>��Q6a^��� �|��yYaaVn�<gޓ;�.�9D���B���a�d��d)�-�qK��L}Jݘ�'Y;q�v}��pY�p��C̿-�}@����Y�ʠ�ȓI1d�����������х�lȐ�A!�ϒU� X�O�1�VI��{���A7"�#�l#�t��S�? ��3%��7a��p�bM�"n�^���"O^`QEbƫY	� ��X)R�j	 �"O�=��I��t��AV$O~*��"O t
�Ϝ	C�E"֭c�K6"Oԍ��⑙q��AA�L/sb$�Ȗ"O��z�H�+)� 
K�<�9�"O��T(֨p6���u�ϴ]m���"O�$!��_1Q�����UmиrU"O���G����ɕ�?����"Or@�gC�8�豒%CD�QbD"O��D�>#ôX�bY�z��X��"O�x�F(X�Ѫq���#Z1@�"O���c
ߑ@����d�
J�E"Oh����ީL�&��S��"ܘ��"O������+���cB>o��"OrH0K	S:&����Q!Zc
��2"O� "��q,���c�UcZI{f"O�݉�擿T���*R���p^~�+�"Od��S�V�^��@�>'4��A�"O*�2D%�&�	S�C"q"��(f"Oz���HV�b��m� �>���"O�1� ���"�a@Πn��=
�"O`��s��Ow�<8D"-��S"O�*��K6�X@� 	5\X8�"OE�'K��z��l�� �+lޖ��"O���6)<��q��J��$�"O��6J��^0Ytk'b�l�i�"O��Ї[�\8�zT�&0�`1�"OD�p��<D���1bjP�F��Y��"O�M��Ǐ*QQ��r�IC-.��ܺ�"O�5e��-g ��j��O��8jv"O0�	�C�&���h��$��z�"O0�#B��!%�f�"!�P�rGLtP"Ob�a�iZ<;��҅��cFR��2"O&��Nf�dE)&E�o.�&"OZ$�d+[!�����A;,9�tZC"O%�7m�!�I8s���
c"O��P�/ذ/�3#�*h�Zx�!"O�0��:
��P+�g*y.B�T"O@��LT�q�m#���"O�`�bS�JL�8��(a+�]�"O�-�SJ��S�f��v��
+V=�"O8h��j�nՓ��1�� "O�YQ���K+d`Xǩ�5 :I "O�Tq�k�µ��i:6���4"O�a��aN�Ẍ{��r��+�"O��X Htе�HzT�"O 9�6��.�p�Df��0�JX�"O*���N(23rE�`J�]�̼�"OҤ����>Y��1qoY�Ut���"O�Y�s�:BI���cJ�8e��"O`�K1��uX�K@�{����"O͒Gn�>/Y
��B)I��"O,�t�',!2�����0�*�"Op�����~>��هHFt�f"O�q�f���c
r��� ! b�0�"O
l�WOK2rF�U��L�95]6<hW"O����(��M�w�%Dz�"OڝpqC�.[�h��O�5e5\)h�"O,Q�1A�������~���t"O�%�5��$~R�d�2�7`V1	W"O� ��IZ^��Q���T\t(p"Ob(A�ͤZ	�l޲�d���"O��;�	�*���l��!߾�I""O� &HA�F:���B���5qޝ�D"Op9bBLZ�b�H6��R�C"O�zpW�SJH}	@\1",D�s"O��C���)x|���ŏ�Y�p3"O@q(���?H���c�c�H$"O���EM�$��e������#Q�!��حbsVX�4CQ�.~�i�R#�!�$�8[�R�k�c�6P ��E�"�!��{��0:���	6N8�!	�Uk!��dl]2R)֏`��J! �{�!�Ē2"K
$��Cȯ|�6dЃ�Л!���*�Ɖ�:�, ��1�!��@*.,��:�i�7mvLQ2�
�&�!�� ��l��4�͝��9YGŋ�!�D�<O���"�S�n$Jnߌ�!�DD9Q>@|5i�3G�vu`�k�L�!�$�h��pæ��!'mNDI���A�!��
v}>dr�.�7�ȵ"�f�?�!�Si�<�#��G�HT��DIv!�
D����2r�vѢ�hL1�!�$�'u����՘%H| q&f�(;!�00�!�F�+*��	a�*��!�Zu�Jx���95����G6E�!��Vj枹��ٿ&f��f\�f`!�Č�	�9Y��184����7'O!�$W���9Q���r� 3���$2!�$�E?p���M�r�5�f��0B!�䛼a,��)���sm`p�� �-�!�$�`<"�D�S�uK����!�D�>J��I�	�"=6���6፰ �!�$ԛN����0�$lň��[�Py�]�c�(T�rl�����f���yR�ZC�v��E(	+y3Ќx���)�y�A�$f�jEjG�o�|�å���y��b��Y���0�L{�iT��y"b�@���5�'�����k�>�yR���5�hY�3�="���8�yb��Wz�Z��0`H�ɥE���O��DՔ	<|�zݴ��Ogh4�dJ@���dI�/��OUȠ#q�>m����O���ή#�x����7� d���!:Rr���Z�}:�+E�4�\����FZƈ����;/F�B�-�5隕jVǘ,w?"l��`�=����i��h���Q�AD�.ɪP��"Y���M<�F#�Ο�	ݴ<�O_���bLN�������g�Ȇ�8�c������t��3�戹����m�a �k �������!�ܴ�MsĀS9%�ҵ@(2�L��C)�t?i�/ ^��'�S>���C��	ۦY��E�n(��)��]�p�6F���N����-��q�'��]��*o�ٰ��)����a����	�s�T<�.×�t���-c���I�0������ٖXe������	��\c��g��[��i`	Ơ��=�۴w�D�	ß�),O�t�sӮ8H��ֹu �l!� � f6d)�O0��4�O�X��E�<Si���w�[�Q�2yҡ�d�O�|l���M�O>ͧ�u'�Ǜ|�q1�S�n� ���
5B8���O^�"��d���O����O��;�?Q�4D�����I�{��iz�N�$�p ��얕U���4��.W�^H�#LJD��l�j�'&���C�G"]	.8�Go"@F�b��	4� c��JI� Q�9��	�067�6,�D�����`(�%%f���K�X+������bd�I8L�k��J�,OTa����d�\��@pĎZ^$�lhf�עB��j�8�ʷØ'C�ʓ~ n���Ҝ	��o���M[J>�/���)&���oG�$����F��:dz��!�dW�����?a���?!�!A��?����?���
*w�@��LO(�R�[�-�����(��&r��k�*U�<���Is.�I�Dy��J{�ۼ�\E�se��}��ʣ�ü%K�f�ձR�$a�H�&s���$ �N����1*\j	C%!�+zbq�`��:|�Bs�"�d�<�������)V�}�(��m_P`� ���ZSqO�O�"=��k�2A�eK-�'�S?�`�`}��V�dv���u'�'��^?=��,�%���pV�&����³�����?Q�q�����(4IU��8|�QP"ϳ&��!�A�ǟ}��Pq�[��$8�e�y�'(Eʰ˗En:uB��l��!F�#+Z|D�a��;F<i;ㅛ+R�ܤ
�e��'Z��[�SA�6c�J��~� ��Ben�,\�Y�+�
H:܍C�����?�O�O����ξ0��1㊈$���֕>���4��l��M��4p��,ɂ�M�u�&	�@�_�(kn��UX��I���?�����~h�D�O47M��`?h��Â^��Ȥ[�@B�^�l�$��X�QI��UcdH�&�;RQ�]�0DA��O�kl�.Uu���v�@N�0� `@R�p��/�c�N�y�K]�!j�+d���j��1f]Z��� )�-x.]QG�؅H��P�E�\������O�1o�����O>7�׿9f�Hz�
�Ј��\�WQ�d�O��Gz����R���[�u�%&�����'�"�uӊDm�[�I�?�;R5��!�&L����'(M!E�|2�'i�LS� ��(     �  �  C)  �/  �5  N<  �B  G   Ĵ���	����Z6)���P��@ZT*B��5Q�����0N��?]�P�	W&��t����%��X� ڳnS�q52�ȓR���a�����5`G�8� �c�lH�"�h�!iYd\�c��;\ޮti�`� ��E!��8��FIޞ$���#���|!����$�Uk� �h�rKZ
`8H���P�.X�Q�7��Q������t�a�F-n���b�$�ʇ* �Ƥ�E`� �p��u�]�C�������[R�'���'��֝�� ��酬C�p�%ټ���#�e��
��с$*XIz2+�$t4���Zw�����_��a�'�=�H�X�!�*iD�af�_ lTd�@��S?��	�|�AG�L˞�bř��y���.#vn$���צ@�2���dգ��$�
^�����$���I���9��St� r�	R�8UUj%m�_y�'9�+)����:����Kyeh�Η�3�Io�"�M�Ĺi��'G���O��I2Tt���V�@�W�x<� ��"
V���ŋ/���������,�^w!r�'g���6 g�UBd9I�vm�P/~�f�I��VVl��eL��(�����9�8�Bl��D��M(q���pvL�JB2[X��*�+j�&�و,�������l�"�rd*?1%K̟��/�6K>�X�Lۚ_�Td�����MC��"}��'("�T?Ix��m������7u ��i�<��O�b�dExb̏:YHT\�O��v�6����ї�Mk�b��
u����DЦ=1���%�M���?���c@ʭW�Ÿ���F�*�f�֦��D���\��ʟ��0�a$� �r��(r�j���Cb
`R�a�!�tQ�↦��xqCFٶ#pڣ<�!�!�H�`� λ9��0X��W+�X���&w�I���Y��T�5I���<�A)O�hA����z}��26a�W��uDA!򄈵X���O!��Bݻ6(�'�ў����dZ�����^�V��lba_Nm��/�|��4�?9����)0�N���O���*Fq�P��ǎp��Fᦡz7��%�:����9��`�S�t�	Ն&�YyVGU�$$A`_�;0��P�QT��%>8n(Ѹ���v@��U�؎��;���e�)�;�TJ�!K�so��Ņ��y}��I�rN-���[@�=�"��?��!7+ǈo[ �ȓ�F�j�@S�=�(|�G��QjiGz��$�'��!��/u���,�k���4�iJb�'���1�I�y��'���'�
�]�֘�6���ȓF@`Dȑ�L4U ~Xh��,�ȗ�˟�cWg�|FyBF�YYp�t/�$�h����,-�v^����ܽ}<|�)��aj�/!J��6�\�#��Ӆ0H�jQ�n�>��'���˟8F{��OD,���_q����cT��)��Ob����~�~�{�B(�ق��Ħ���4�|�D�<q�	G�0�t���Y��.3q�A7,	���
�?���?A��o��n�O<�a>9a�m�OT���/E�{�@�f�
 �VX����Ox�D�V���ˆ �/��
V-��+ ���2�O.����'�6 N�-y>�qR��ޑ2��Y[��2D��f��i�2��`L�N�e�$�%D�|Q#�
g�J H��N%gi�Y��Τ>��i��'˜���c{ӌ�d�O���&0R  ��O(:N��	��T�)L.6�Q�3N���O~���e!���4�?��W�S�L�NT:?�*�K��"ړ(� ED���y!D5tA>��}ZT�hO�uje�'E"#|1�F�m�DY��>�4�� ��s�<!C��-ߚ�as�
5=N���bAeX�`q�O�� �-Z6'$�%R�(���-T%8@m۟X��C�Ī�?&mb�'@���m�,d7Z���!I�Z���pӂ��Fj�O:b��g�����L")lT<���
�=���m"<E�"��b~m�¬%g�:���n�%{SRf׆�?�1�|��I�D�m�b��=��Yk1&���xB䉽N6���$ o��@�e��}{<"=!����1�A�D���O����1ٴ�?A��Ggb����>�?����?���{*�.�OkL��u�V}��B� $�����Ȉ0A�H3U��|��y��F'I̔��R>�<!�m�6e��K�nU�eu��0��,�@�	.C���(U%�3XJ���(O��j"��i���֠K�IZfرUR���'r�	H?1�I*a�`8���&V4��B�Z�<�nىT����;{2�Xj�AԦ����4����<a��̯d&\H�1J��MFŊE�xhXr���?���?	��P�n�OD�Ds>�F�� 2� .�$rD֩8eDֱR���
����H�CD�Ԓd'�x��M�U�Z��ә�v��P�
D����lG�(~� �ꊰ.��$���3�~b-d_��P�еDwD�H���6�9ړ�O@��fK�.����c�Ǥz�"O@5+5�!��aT�����eS�\cߴ�?�+O61��*Z{���'��)@f�1R�
�<JHx��,���@f��'b�*���@ S��(��$�="W�$��*ι"l��B@R8n>����j�!Z��պ,�ٳ�^�X �#��Pq&!r" <� �4�����D��T!�ΗW9�0��CI�'�<�����?a��G@�I{�Qp��(4lԝ��$���$�ON���)��T�BK+0�ĹҦA�o��'dў�S����(�x@(����˄��|��	�.��ܴ�?�����ICM�*��O`3���m��戢K�.���������A�9��X0gO�<x��T������(��>ܐ�Ɏ'NQ�<�%�F�0�	�.�<��Ǩh��T�#,���ȟn�SqNMY�$A��O�����YPa�OҜ���'��7�ty�'��Ԩ[�*ގuB�쁕���`� 8g�>����p>��i�3br|:��.^�|�P/I]�'�#=��O���(�kҺT�VA���N�8� ���4�?���m��-9D`U��?����?Y��p��O��+��\�5�TXb�k��5��B�VlymL��p>��0��C4�s-��
gy��ܫ�p>1�F)K�=A�B�A� ���_y��:�?"�'O�Ir�)B�FF�`��
N�Xs�'(� ��ցv����K���D�ߴ���A�I�4��4��&�$�����rI�(	 oZ���	ğ ��֟�^w���'���ȧOȀ�F��%��q%��0cn�yC���3b4�!��Q@؞a����$���w��?d߶UZT얳]�vT��Em)�$J�i0©�I4M$Z�ڀ��@��|Z��;(�]#�'��� b�P (�:�(��Ҕ ��� �'��hcw��P���+H)�$�*�Oxm�{�	�#	f��4�?)���E�k��׀�bfm�����M'��?����?1�釅�?i�y�O������PKֶM��h�M��M!��dеQ?�qqO�/!�ʥ������*ӯ1�E}\��I��d�Ԇ�=rg`;�e�Fh,ɡ�"OfU��b��X@H��ws��k��'�4<�j���.L$� �kYR,�' HM���'�B�'2� R#��IΟ�ef/F
��ţQ?�ܜ��K0�M�� E�+ܤ������t��c���<��̩�J<�]&8p�L�jnp�� �����ED�N��E憫gs�8�1��N@���8Qj���'(��Q��)Ǯ`��	���¸d�0���_�rp�	��D����IBrS��O�xn�S��ub�B��=Et��ʤÌ=l^���O2'�8"=a1�S9���e�
�o���S�� �I��4�?Y�&΢\B �Ͱ�?���?��~��O`ВłN4��#���/>���V �����I#]%xx��	�w����4�]@�ʈ�g��s� ����&tCpI�g�)	KʱX��3ʓB=�������b���E��'Pt�+���?ق�x��'�B�O�	DŖ�o'�5%B,�X{��i�ў�'.ݺ=�'Ĩ �IY�a�Q��*� :O�y��h����'�剿����O6�a������\��@Z��M��,̣��-"$����?q��?9g��d�D�O�ә�Y���[�\�P0'�]7-�p�q� ���DKErz႑�I `�5x�� HɺG���G�<����lU`X�(Iw:�zul:l�}���<w��e�剗|6�d̾-~a�Èy�������tp�ȓ]e�ᩅ"�I��u�F!�!ebb���K�'G�0��VN����#���O��mZL�ɽ`μ5۴�?y����@����)����m�qH���M�7���?i���?Q!��'Ms$q��<bD��6�ޕ"��i�(Mx�A�e�A
j-�&��H�ў�����ɓ�5\�����߄Z��m�wL�Q�Q�%�1R�fX	�b�
��D�2�0�kPF�I���)� )˲~4x����^8y�����"O��g%Y@4�z�cK�
�Vx��i>���O��
���"�2MӤ$�+̂���]�����\�	�<�O�N �q�'�LI!V�l �#C�P��-9��e�6m��w���Y��5j�:�� �M�O����|���m���I@	�*)�F
���?�#�ťz�D(��ۚZŠ����'P��gO@ ��`���|rq�Lf�T�Ҋ\a�2����?��`ȟd�	a~J~�M� �0�h��"�T�?=&�R�	5D��h���v��H	��,���R�i6ғ0L�?e�+׷Y��P0F�#V�Υ��)�M����?Iwط"8رC��?���?	���?16����EI�eT>!"x�D�K�4��0b��r�0k�����A��qݱ�g�'[�D�H°k�r���-7����Ψe���2g�ǚ0r����\�46�ΧC���i@�\6$ �қw����.�(!��I�w@Q�k_ �J*O� �V�'���If?y�C�i� ��@˹>jhOW�<�Gj^h����6�jy�L�e���1Џ�4���$�<�&��}J!����P-:1�>i�љ�HY��?���?���g���Oh�Da>�ЅaվB�p% �b
�8�28��NL 3�!�wDh@l0���m�
9����Ѥ~��p�!��9�E��N�;ȗ�G���c��
d)�fD�|�'�d<2�w�� �Ma�Z�8���J��R!��"O�L!�@�m:�8���.fH��x�"Of�1 �05X �tn]�]��uɤ\�T2�4��P6���t�i��'���'Ul<Q��#�3����sjC�<��fC�L�"�'��:xr0x��)O�U_<��pgنi�	�{)few'�߀M�����ў�z6GR
n���(���.W�$:���$kz0i���V y���3�i�00�R�;�C�a�'�b9���5�>5��̚3ʼ%�t%�^�a	�$.D��5o�*}��X�g�,��I��*��/��|R����PLT�.���B�Ɵ�4���>�@C֤?����'��^>�{"�ğ��I)QY4A1��J�fv�lp�l׏H,̒�4 $J�P�.�H@%�R�Ýo>��*�4b>��6m�%� �0��j�0�������P[�	�=5�����$,D�6��< ����cc2�%P������!�}��Z�_�����Xނ���R,O�O����O�aܪ�+�'�T>*}�GC�f~!�X�X-zm��Q�::�5�W�[�Xj�O���Ie�'���=�d��4fP.S
�4����
_w�6��O��$Utt  2��O
�d�Or��ݺ���G2�I)�ھl]|��,6%���C%������,L��`��;�3ʓ�,X˅��7-�q�F.�,BA��
O�\���#K�����"H����' A@q���ޓt���;2��l:t�O�$��)Y���y�'� 2�?az�N��V��9rC<-�ذX��y�o �B@|��(��2R���M�i>y'� x�m�OwVD���N2#H�WS!�P�р�ğ ��ٟ��	1�u��'b0�
#�M�u���'	2l���U�o�	��@XF�r�(չ 4�-��'S��(O�	�����lq�,+v
Kn��WR��(4ӲK���"�P��M!�J]��(O�UYW�'�ҵ"��Щl-�Iہ&N��x����+D�0��&�A�
�s���$6�qt),Ol�<��g��>����M�=eT�3A�K}�i�ڒO���&[��'�Iɠ#����#oR�B� @�c`I0'"�6� �~|��'�L	v�N|�ԅ��E�2��ǀ̦�(om~��U�e�����D�l��=i�,��.h<Z�*W1H�&�o��In��j3%( m��h���[���B�җU��L�KZ��r:?�� �͟��4H�1���qeF˛~�(�vJ
B��S�[���	v8�����0�u�W�S-A����6�O�x�'&z(Y���:JzΙ�ܤg����O&�`��E��a�IΟ��O��9[��'�b��k�Ƽ���q��x�▙r�H6	 M
�"0�S��lSP,PP�<�R���c>��������+A��/7`��B��ğ|��?%b*)3P N�g�L��%\�0�|UR��	Ӽ0{r�)t1q�
�^�Up��'�����Rɧ��r���5+�0]�C��<G��%���?D�,�o˨N�֐؅&�O�~5�5�<�	�����4��m9���n)��mY^e8�S2N��c� ���ꞢZ�a}��	S� ��I7^ꍸG͝�y���~f�+ff�3\�I�h��yB'�$SBNC�)����&a���y҃�,�*��sa��j�H���K!�y���~0VA�E�V���FD��yr��GHi"���.v!�bdR.�y�]	6h�LC�ф��<R掐�y�I%�4C���(�d�%�ؘ�y��-8X ��7NMX�F,H�y򆌲$��P���40��mɔJ�)�yBN)[�	� ��%��ɠc��yB�F8c���xUjK�	�^��C�O��yb��s������k�J-�R��yr�Ȱw�����w�3#\�v�4t�� �p���&7�X�L(#�f��ȓ�X���� ��Xp�Ѩ}�x���i�$-����V��P���])�`q��_I21P1���Ɏ���&�6"1��B�T�P�nĒ,��������8�ȓB8�=�Q��ʒ�e�'g�\�k3c4D��j�^	�ZPגl8\���4D�P�wN�ND���P
֦�6�p���_�$8�F �-��m[�ig��#|�'��7��Рd#���l��'�=:�ID��x(r# E�"����1�ӳS��D겄�w�Д( 	X8��
�垃L�Tm�VȞ�Z����$ 0LO6|*fKO=y��a`D��n�`��7/�p���S4:������Px
� �E`hR�G�� P9�uH'�$pyTuI% M�A&�x`�Ȑ��O}G�R#y8�)�i�d��6D��s� $3 r�c�Z�G��Y#�Q,w>�@0(G��Dzf	�%��#|�'�^}�AR#UPVlk���x^.��'Қi�Â�e躁@J

"� �^WZD豢i�.�P����h �x�ƻ����)OQ�^��`��	r�E`Rnpa��Zov-1&��;s���F��J�z8��N�2#����/>id +�[�V����L� eI1Oz���H�0E	����N�2��h���BĝL�j|�ʃ�N�z4�DN��yb]�}%� ��\�{dP�	?D�P�S��P��ԹH�K�@�A��lۦ-ёN6�`B��S�
婦��<��9�S�O����L4�Z�Yq���Bڊe8P�Y9/��E����U��+��(O�s�J�z���x$�G�+re��|"�W��'
�=�'y�i �ݸ]:���bW>+������@,813խSOx�01�wM��ŉĚG��9ڰ�	�h�y� �)Z��j��H�{�$�Cܧ#����2lܝz)2���C c���D~�ʹ!c�#|Z���3K>� �*,h�l]� ��%��=�@�-`,�����^AP�D��O�5��lW�Y~鋒L]�-�r�;��O
��CO�$j1O�>�Ѫ�cL�Ց�!�/e��Z�O�,1�
�9�LM=I�r�`T.�5��xb��8i�U�`Hǵaa��J�����+C��)�f�O�p#�O��0؟��[�'�ћ���)j�����,^G8�em��8�I� hKh̪�I��y�r�k�/�8 I�1�NN��M7B;m�6@�R����W���~��Wr�'1^ʙ[��,1�SѧK����<ғe��1���Ob�?�#bZT�ar7FR(s��-ْ�*�����QR@Rg��D���8܌��B�d� o���A��ww ���F�
yF��.-��zK�b>A2��U����c�6=W��:~i�ɗ�B*(��:�kۣQuح��\i��� �'D��/�� �k%�`�R�J��-p"�h�	��r~� U�T�D����?��W�W�|^ұb�IК眅Zf`!|O��u�I�%���S�G�V.x�(�me����Ƕ��k�ǯA"0�R�O��~2��"P�^�%��f��
UL*���(1B�ƂP�K�xxRc��$��
W$��-���g��da9!D�90�Pöf���yruB��p<	��.7H���g̍E�~]�B�W�0y �p��I�<���Z �'dx$��>��cԽ%P�\�D�_��B��Ɲ����D
��:P�"�
d�jC�71虫�e�5�I���_8y7���:�&lR��	�D[`	��/�Sh��O�%�G�O��O=0c���a�Ȩ��i�^&�p=)6��?�A���~u��SEdF�ͩ`" X ��p��,u��E���J��ч	
9*<�QI?��#}�&V�A�{�N�0*$LB�m���'���Z@�s�ݯ`Ď<h#�~"�"^�?�6����#6�Pr5�B'Y�co�	 ���2d/73(up���U8���c����<�"��V?E�� �91���I%��l�\qi�m�"�i��4�\<� ��6��D��$��?ip�-j��1��x���ji�&אx҈6Qz��a��EG���A�I8�M�"B���������#5�0
�	L�t擉i
�=S!��|Qm�l��T��2b�E^�����]cV\�A+�XEX�N/"��	ؒ+�Cy4�p��M�E*��!t&��M�2a:�C�X򓐍�Kn�p@����L�C��%T�?� *�
b�)*�R'��'�\()�ʙ�l��p�N�ʑ"��Z��`��N�onţ7�	�0=ɤHA==q����.N�<E�`0�i�
��/۟n�ӧ��#F�_�\�h��@l����Ea�E�"+ļW���E
N�t�4�6D����_2l���ӭ�6�,Thփ�>!�I���4@ie�J�>��y�#aӺ	�ץ�V�S~B�!U��2V�������#������[���I*�$K�e{�Tz&�ǥv�v�У�C�6�l��j�D��j�^�3�	�em&]���J�}喭`d.�80%���D�E-�-Zt�I�T�x䀧���Π�&i˲e7�I�OX�x@��I�_�f��p���|k��N��?���˝v�TJ�A�s*�����OɊt�c�רh;%qIZ�D3*��
���V��!���e�<p�����H�6�}R�ĉ�kh�bS�OL2U�u"WF/d̉q��589����'��"��f=Z�C���A@�S�
b !�S�i+�|I�U-H�ϸ'�8(�G�\�X��@�	�[O(a�v��(�E"Q;:�,�;��F�r�*�k��T�[d�����ڮS��D)��'�\S�-7L��kW= }�+��DU��\T1W���}���0B�\�?1�×�"�� �уWT��!%,&D����	�?*�����S3j��`$D����958�i��P��H��bl#D���Ѵ5�}е�ʕF>��E�/D�� `͸�E
h�^��D�*d��A� "O��0��݈_d`*V�}� �"O����L�{t�؆C�j��(Ir"Ox���ٯ5*�c<6�r��"O| �"l\6��'aܒA�
�pp"O^yF�;���� Б!(�k�"ON%�f⅜S����Ҳd��"O������vظ�ᒠ�0_en\"O�����^Js����?o���"O��H��2B�@dro�_.u�r"O�m��J�nhڭa���D�����"O	8�
d�]@2�y�l�F"O^9���a�P�4牅R֬� �"O���h�8Z�((㆜>\)�6"Op���O��i�9Y��'���B"O�xb���ɀS��O��Lq"O��R�d��I;2t�9I?`P��"O�a  b]���b�&�pV`Us "O�a���7pe�Ȱ`��]���k�"O��6�Z>sA��I�'��?l(]k�"O��s�b�Hyh�,Ҩ#erP�A"O�e��q����#��h�u��"Oz�Ҫ�U�i�F��	h�T!�"O��ԥY(*}�;Cũg\|��p"O,�膧�1CxLd�C��1n�:��"O��s�*R�w��1`=�A� "O�(*qD����w(O�,;
4С"OTy�MQ�4y
(����I$�tq"O��Q�	=m$�4r������B"O������4pPE�4
�E�W"O�YP�������$��qd��"Ox �"�ϐz�y!��EUֹˀ"O�@�&+&ez��`���L�"O��&�]b@0� ����4"OXl�AWt�6���"���i�"O��L�P��8�D�K���Z�"OK��J�kuA� BF0z7˗/�y��Z#�4X�lF ^ز�c�'��y�h-+��A�&ő�j �`�!e.�y���<`�l��a
�
`��HBa�&�yb�-�����]�.���#@D��y2�M�[��t��˲:l�2��>�y�̏%�H�g/3��:�����yR�S6,�!�J�+���@W8�y��R�K�&�y0l3+u�4h'a���yR��"d�6�r�F2�V1z6���y�	NH�3CB�)S�$@����y�
�>,U����G1L`���$��y����b��`�L�H��z��^��y�D[�����ܽ|�H@��0�y�a׊h���gb{Z��4�!���u�0�i�����cG?7�!���&��p���D-�v1�d� 3 !���5-�0���G��-�l�bY-FH!�$S�x$��b�ع/����D䞕�!�$�`w*�y�gW.S�>���LN��!�J�t2E��y�HP�l�6u�!��Փ,(�
M
�u馕�AFޠn!�DĦ2��mzA�A�',�@ 0!��>u��}&ى]}���ՒO}!�Dܟu��P�4DNIu�ԫBz!�$��j� 1�P,&��"f�B�n!�$U�%���E�	�m��� �Y!�Wb��B$ L�VkXd�ŊPR!�� ���� /,�2ѱb�XTK"Oڹ�p�Ex��q9�)���ek�"O�L����%ʌ�a�&J(F���"O.8ʇeW�b���&#��29>�y�"O����OO�5�xds5䏍g� ���"O@�3�[ ��@$яy�B�	�"O ��F�*u�r��KS�s:�{U"O��0���'i���Sj%Y<|B"O&,I@+,m���;�H/,M^1r"O��5�0ѫMU�FZ	)�"O92D+��>���pF��k_�ၒ"O�DҗΘ�|Tɒ" �9*IN�AC"Ob���e`��B_��*@"OJ���ѩH��PI0�CI�~LH"O"0ʡ`;D�8bḷB��	�t"O&a�C��[;�$�c��s{4� 6"O��j"��7i���H�PiP�#�"O.(p'�6\���D�ua�؂U"O>]PM!RX��S.�>@DX��`"O�3g$���,]#��V�E���s"O��Z���mu6��+ы2�p`�"O\ �MU�h�|e�7�M
��1�w"OX�c J|['I�R��q��"On�;��&�\��#&��x��Q��"OJ� b( �G��<E�<8�`"O �A��_�:+1�'2��b"O�=SqV�8��<�$�Z�z�P�"O>��!��A_�񰕢
,s��̒4"OR,�û�,Wf	SDB,�~���"O���B��3\~��B,B�,�Z%"O|Ȉ��M9�)��K�"��af"O�y��HF��Bl���^����'"O��Ɂ3���b�JR�m��Q"Oȩ 撫J��� $���1�0"O��{�i�"Tj(��po�0SB���w"Oճ�"΀:�#d��>�D��"Obl
��X�(dJ��R-@q�Uk�"Of��e�ǉ0N$@�i��U��[�"O��Zʉ�p�f���o]�_I��`R"O���^i��`��^G�� "O��B�O��=�����K���"O���r�_3W� �07�'O0]�t B�7~5r'�ZX��H���"}���׮�n  ��?D�8�a�6%�@�3�l��B0X�k D�(j��J�.q��8Z����<D�x���_<}��m�W	��) ,�0�;D����&������4,y�MA�%D�(����6X���s�*ʸ{D�9���=D�t��M1#��r���!D�Dr�ˬ;3��҇���k�YH��!D��$�3/�m��%1���[��3D�pB��	/s+6��p��7s���R�1D�L����}�m��Q�D�3(0D�8���M��`k��tef@�$")D���B���e�Pa��<%��b!�%D� Ye`��H�T�B�/w�Lqbq�.D��D���X���̜W� �;ӈ,D� {��׹v0�X�C�'��tA��(D��A��A	�&OX�4���P�'D�����Y�������Hxx�8D��QT��g6r�B`���1�2,ѧ":D��� �7ѲiQ�jЛ9�$L��k8D�����(��}1��N�*<�Ӷ6D����b��`zo���w�5D�� ��`���&,Z�ʙ7�MI�"O��!&� E�\;�IR�K �YR"O�p��
��|<���˝��}��"O$���c��H iT�5|x�"OF�H�+vZ��ĂY�vmLY�"O 8Z�P�`��	#A�	f�l�"O0�%_�{��h���Na�`�"Otɐ�Ց1�4��A/	LS܀�"O�M�QA��M�w��T����"Oj���w����Ar����"O|�ӷ����<�[���^1��"O0��r�J�h�N���
�;J65I�"O�i���0y�`b��W�����"O��� �3�l���dY2x���"O�4P�o6�q�BC�k��#�"OȜ!�B�P��4]h����Ԣ]�!��M1<�S��!'D<h���e�!�ʺs����O׊&�n�#��[��!�d�!e��H1RH�_@�q�+- !�d������%e��\<��!]2!
!��j���c�H�|=�I𕣓�W�!�$
���eN�$���#��\�!��[�)1f�M|#<T�T�-cs!�dO'�����^����8Z\!�$ �/�RPb�O�F��L���C��!�S�r�(��ľ�j8J3#��j!�D�D�B�x���4H��!�N>"�� �dwd��D��!�S�H��$S��ђDN��`Iښz�!�Ę����+�9>��Ч�H!�Ĕe a�&�V"��@����>(!�$ �'���f��(f�3��=�!�DG� hz�I�g�by��ɒ�Y�!�dĽh1��:��E� q8ah΄-!�P�#��Ѣ*3$V�<��,z�!�$����#j6H��H��P�!���Yb��
�EK�v��qҲt�!�D�q"�U�%Ո51r�́8O�!�ۧ8h�|��,N�k0J�2AK�c^!��Y0c�FǘUtx�	�*E�4;!�m4Z0�d]5Th�vKQ/7 !�EEU�qb=L8�����N!򄍒�@��v-HA<�(���8$�!��4�
�����0 �څ��&�!��-j�>8�p�
^�f0��V)T�!��._=�d��l�?�D��b���!�d
�l,ܼF&��pS�Y��`��s�!�D�0.�y����RA�J�O h�!���"^���2�^X02�p��F4�!�$�f��)�%��G:"���ƀB�I_r�AT�YR6t��s��Mt�C�$_^��t�
�)�4���p�<��T>(�,�5N��f`��98.�a�*5D�<bc��4!ְ�H�?@�	�*8�(Oܢ}��+T�Q���3��xc��X�D��o�6(y"����� ��?[W�m�%3m�	��`D�E��W�v�RS��8S��ɲ�<����0B����y���6#�\��C��"D��BuO�nd�����B���a",�� "�4��Ӕsi��%�]�D,�maF۶(ըB��)R�6D#�#�]dr�a�j�xs��d�H���߰{xhȹE��<G%`c��Ώe!�D�+t>���0�:4� �Y�,W.��3�O^�13��4����6�p���'��U&�� ���j�#Y�2�b�-�0����@"O��lErB���̕t�>�kP"O.��P�?w�T�`C��i�"O����L���X6F��yO�8�"O�Y:�ȝ�6H���q%�$�jH"G"O�D�q'�l���tIV�M����"O�h�N�	J(���b(�-spZ9!�DCp�[�)F
w��0RF��:�!�d�T�� Ƣ�%@i��(r�F/�!��$�ř�#�Ea|<�$��!�D�x,��� ��H~$�3ED0�!�dT'U�~U�r�؉_2�K.�o�!��gP��d�/u`q�CB�<;!��B?kE��kGh��`aǦQ�#E!��][�t���QsD ��OB.6!�B�.����t>X>H�fi�2,3!�DA?
T*t�ΒI����O!�D���5۰F3),�9R��$ !�EJ0`9񑁇�t��aU��:K�!�d&m�ʁ*��f��B�K�~�!�$�7[fT�R��U �a1!��5�!�DVx��
`k��w�!/�!�$P�=8�5�c�ūB��� !-�!�Ċ�U� ��g?Rd60�R�޿Q�!�DO<J�������z0�M�$Q!��u��	p�6R�� ����o�!��͞
�$ դ� e� ��7��S�!�$1�n2 k��|�0A��O�#|!��^��K׏y$e1��׬R!����z��L[H�Ġ#R�".!�$@���qa���v�Vi@Ҫߡg�!��C�v�QtdF(m|d"�/(/�!��T-h��;�!G#8o��Z�M��k!��:K��;!�F\.4�:r!�	tt�:�E�K�����l͕i~!��ސo|���� ���'��(RF!��S�fa� ���e��x�$l��	"!�d3-\�L1n��\rD1��A�#g!�ܸ/<�A�T	)&z"��� ��}!�dښ]����� �r���o�*�!�DA����AF\2�$��dW�+�!��#e۰�)���
�����?A�!򄂮X�� ��ESu�	�B�(1�!�Q�-8�2�-Ra F�G�'�!�$I�w� dMbR��"E*E1!�ݍzt������'9�4�3( !��E�Ciʝ�t����dA� �;M�!�2���j��3��l:@��&|!�Uu��q��*I�Ԅ��
�\u!��5y�l8�w��'�d�R䓸QY!����l�;҅N�|�Q����;�!�d�
8�bi8�#߼kh�l�3M!�D��1$�@�g�(R J��.!�U�QV���G^2Z8� p)׃r!�@���a�1B�
U6�}���T:!�31�F���F�%6&=[LY�`�!�`Ǟ1ْ.�<<�e��E��rR!�d�9}�J	�$��}3�$X#J!�X,FaJqA`�4$�1��L�kV!�$ٯ��j��ă
؄�%O	$7!�d�a蘰(@L�,d�����4!�X��`!�v�j�@�˳GI!��(��L��'�*C��c�υ2!<!���	L�F��_C���N�!�� ��G��i�Pp���P�A��8�"OlTB��_}��d�T+"@���"O��3��.�^9��ϯ�L���"O\�+rO�h��a*R��N��k�"O��5� �\1�g"P%x>@�"O�I�;el��ˢ��u`@��"OZ}{5& ��j�	E,6)E�<Pd"O�R@�А!@��ɒ��&m��"O�����
 9�lS�fNm�n��R"OLP��5�t��hĕ^0lP�"O��0&&K�rBߴ)�f���"O���B�
Hܝ���(q��3s"OX�a�q���j� ̑(h�q"O�5��iع� X[����-�"T@"O<`KT�l|��@�-�"2�l�F"O>l�A�]l�^]Q2�z��x��"O�d�㐟-�x��p�5�,�hB"O�� Q�� @����`)�{���"O��3Gj[޶�ҁi�$K�XCw"O0a: ͈$���d�F&"�ЅH"O.`�t�U4��l��(�6M�J��p"Or�։ν]֔5U�\%�0Ez�"O���q�C"+�NX���Z��is�"O>e8&bޕR	��fۛ~�1�&"On�K@i�?�ljS�ư#�h�4"O� I����@^�F��8��"O���#���sH4yR��F�� �"O����O�,�hD"V  c9��@"O�Q[�FA;AҨehs�<^��2"O���q��;��5��C��u�c&"O� �M��}�|l $�Z�[Ȕ�u"O���E	�bt��3%Ê,M~ы�"O��@�#̞v�N$ �B��nR�"O�|B$#����{��8C
�F"OH ��)}�X�#*!A�0x+"O�-�5%@��<�pt+�y<�#g"O�Q��8�r����
��Q"Ol٠u�&YZ�)A ��>!E�A�"O���*�4�I��nߞn:,=��"OҬ�*['��ipe-��I5�)�"O� �(�*s�h�Є�־P%�}�u"O��Q
x�q��.�B�
T"O0�P�܊26����\�2\c"O� ��#�>8��C�BU��i��"OT��,]p����:�\d`�"OL8�!�&L���C�T�Zt"O
y���  ��a�D@�]:\)�'�2q�T��cf(L���Pp��'��y�+T6F�$�3�fN?�ظ��'�t2�҃\&��c��#�D��'����%�*ƶ���)7��I�
�'}��Vǅd�xA�'9/�z\"�'���6'9"%r�i� �\$`Q�
�'�AQ,�j C Zw�MI
�'��!@�����e!#�(Y�jT��'��ʧn$fِ�a�hA�DJ��'h�@$J�Ap�{UE+Ќ��'���-ȂcP<L[f�Ɓz��u�'8�t��L[�&�8�!&�u��t�
�'�&�:����m]ґ"����n`h`��'��ٛ�!ȓ?�j��u�A.a��P��'&�`d�� u�a{Ud�-�&�C�'�\9�K�^�d��[��E�'Ƞ<��� �
מ��T*߾9��0�'d��*�ߠ'�� �"�10���	�'Ƭp0"� ;�Pw)َ��Ԅȓ!Fxcl	D d��aE�4�x܆ȓ!�H'N^�1�xrB��ڐ��ȓ�>\�s��$���q�",���;�lt��	�
���b�:t�x�� �x�Pi�< MR4��_\%��8�.d��Ϋ1b��#���3F��ȓi�>Ij�j�13C���'!�AF�Ňȓ^����`S�����j�^�ȓ.��36a��E��(H0W(;Zz�ȓd�-�
�e��x�g��l�BņȓlDP����X��ep�)�wYn ��D�Z	qPϝ o�f,衦�`sT$�ȓV<1q��Z�g=~�	ƃI�����ȓ�>e�2�"S�tI�B�p����Wqb��G�@,֜!�Ѕ(�R ��ה��UM۴��;��Dq7�X��TU����	�`0��Y�N�^�ȓ)a��Q6�� �
x9���d`��z%ҽ�qٛ��DYdN
Tw
t�ȓ>�pT��b��\�ZƬ�<Q���{]ܚ��ԭӐ|�V��5;��-�ȓ%t��@��1/���_w#Bp�ȓ&".�p�b�B"� :�+�^2��ȓ|θ9�3%;c���l�
,����ȓ&���q�"�	f�C�R
!�쌆ȓ|h,i`�ۙj�"��B���\h@��S�? ���v,׭<s,ű�͊%���5"O<� r*��&�HC􎍫�Y�"O���f+�����.��Q���!�"O���W�]�k��A��CT8�ʁ"ORyp�N�B��5{p��� �A�c"O��Kg�	�~Dr���Z�a�i�d"OR���ț�i}�Dڦ�!K�,� q"O�Yxq�H2B���Q��Çb����$"Ozu�A�J5,>TpB�FD3��%+p"O��Z�G��{`�I�ܬ��"O�Q��K���;��M����"O6�� ĄZZ�I�R�A�F�� "O^� kO�\��@�C]?e���"O�,`��ӕBY�I���J9:�`��"O���D��zwp�U�ŊH���E"Ov��W��`�F�!�D1+��s�"O�Y����DR,����!:�� "Ob�rTLT�g�4����-u�ʡ��"O�pP���.�qȁW�����R�'���;E˒i���b���Z���B�I0D� �� C���^���Tk�B�ɦ^eF0�Q��,���C�QA��B�I5<��As%EM$Gf�⏚{+�B�I�TX���AF_�5?@B�X57�B��31������yxX2@V .�B�I9�:���ܕx�.�H�i:L��B䉊
�-����b5��+�B�	70*V8��j�;�
�KGTB��"�@�i�o<=$��B�ȷtdJB�Ɂ)��}�v�[<j~Uje��/olB�	82��Ti�M Q��%��}6zB�I�Eˬ]�&BAd��!te��L�bB䉁5hR�P��#h	�x�"��x�0B�I�5ޘI�^�	�0#�9$yō+D��a"��1�ހr��K�P��KǪ*D��	�D�3���G�&Y4��ق&,D��	���U�-"��A�ti8�,D�,A�C_�fQeF?�PeI(D��C0��&&�īa/_�y�N i��%D�HXg ݹ@L3��ީ2�X����!D�� �ǟ[H�@g�v�TS�a?D��X3NK�P���3�=h+Գ��?D�(`$���e@�ئ�)����<D�p�BےtQ��>��ͫæ'D�p��IdI2p+�?�� ��"D����%o��A(�W�,s�3��=D��S5Έ'��p���(*|�h�/8D��k�Μ<�r�����=prY�ã3D� !�EU�(@�, `H\� �L2D�)���6H:�DH�J[V�>D���S僾y�D�� �,6B`�C8D���I�dTyWNC9�&})��6D���D)G<;�F|��m_�H�\�76D����fN�?M�����A���M9��?D�p[*_%l��1ơ�(E�#BJ!D��fσ�
∵�a_.U:����1D��9�Å�\d�0�u3c	��A�"D�����&���HT�=r�2��>D���@�ۍ
nV��P�h�y�W)>D�P�c��=��h3�P�0���<D��Zb- <y�š-����5�n�V�=E��4��(�/Y�P:¤�V����@�ȓAM�!��� 9V Q+��@�	�ȓ6�K�\={���Oo�!j�6D�� ��@��]<}l,��A�@�3ΒH1�"O>��#�Q�	־;0�P�6�8�ٵ"O~%���U9c9��᫅�&�X�"O������|�f�x�(G^���p"Oԡ�&�ǞuW����ڴ��S�"O�5�ꓑ8�c�F).~m1R"O�p��Z*3uv�DÁ�,Dt�"O.8�Ȕ,��#�bD�"�P�yp"O��t�,�  s� 3��`�"O���	 �O>U:���fo��h"O��2Qo΁R�
���߯I3�@�V"Ov�˲�Z�B� SOV�q�t��"O$�xq��!5��q�.V� %�%"O�$�H�-,�J,9�'��[��q�"O<lzǡ]%&f.���&�;��n"Oz����H �u�|��2�"On���/	�w�.@�&K�z��ps�"Ot@B�)`����D�*�ȹ�"ON䪷�	Cp��I�
/@���"O�����Y�zx�1E΀FHBS"O\8��D�V�i���@6b��F�<��.M�_��Y%��f`�L]�<)��G"o)pT��A�]���,U}�<��\�Y����$�&:|zD����u�<�ң�(���풫&��Y!"�r�<A���";X�����%R���.MT�<Q1%��y1��@ T����!/�g�<q�f;~d|1˚�J�yCf�<A!�Ly�L�b2��)�%�b�<y�:D��Y #Y�m.�9e(Rd�<AC���22DTzOO�X���cW\�<qv��9z���i���U"ׯ�ҟ@nZ~�� �@��s��!Ӳ��H�BU�9lO�pQBc.}�X u�H"t(�8"l6�(�F��y�G
@�*�ˡ ��X�% ���'�FyJ|B�cX'T���D�T�����K�<р�]�]�\Ts�	�>��i׋V�HOd�}��x�(�u���t��8�WJdnp��/@�ES�0[����Ii��X̓��?qp� b��QIWl\�	2�1�C@�<��	�?l��� @�n$�Ya� Cx�<���$���y��߼OftIy�OE{�<IR`ʨ6@���A�>{��uȝv�<���r��L�a��
���3�Is�<T��|Ij=90�@A
t��ep�<U-P��D��=�9[�MBm�<�E�1[6ҝ����RF�nB�=k�2Eӓ�ËH�Ukj�U��C�I�|C�{���@aZYx�F_8f*B䉍m�����F��<�Ȳ��>jB�	�uL�(ygB՜1�8�S%	�p��B�;8YdU�vO��o���0��*rB�8�"��O�Z
ȼ����P�C��KY��3���]f�Q+7��$z��B�8����sf�Y ��MP�B�ɀhy���B���j��ia�aN�}��B�r�`�[5��Н�BґQ�C�Ɋb��q0Ge�����O|ˮC�ɂg?�ɓE�;`� �&��f�rC�>��2a�[5��Ф��@��B�*�V�B�$��K%����>�pB�I��@���.]7? �� �#'4�C�ɕD�dX�']3q �G�Cl(C�	�O�T#Wh��-�ڹ��G[9�C�)� d��$�/4�����4�|i"O�D:$�O�Rp����AU�V�<��"On�W��J.��f��.��d��"O�9�G�9Fs��s�Å~5t�d"On�p�Dڇl"&Yv���_)a1"O���jC�B�@�h���mА��"O����*_���+ɓMm��"O�=�Se:̼�hB9vg�ȸ�"OXѓ���'IFi��%iJ��Y�"Or�zn��6�c� k�,Q�4"O�uk�[^r�@r�.\rN���"O4X��%<B��ō�=��`"O� ����-�� ÁT!�p"t"O���d-IH�Є+=au��#�"O6���LW"!�ͺQE"76�;�"OJ��sLB��qFÝ.* ��%"O@�їo �'�F�+D�G���]z!"O4 G T�_��zԎ��E�j|g"O���
���Ե3��S�fɫ�"O.�P/�/AҺ�q�1-��@�c"O�EtCO-N-6��E 1\����"O��3QD�0
����!$U����0"O�����0��@A������"O�5/Q�����X�w<�se"O�0f��]�n��"���Edn<�s"ON�Un�tF��ٖ+ޓI)x}��"O�٪s W <^D��`��U�(� "O�$q��+s��D(ϐa���"O*� WC�75:>�HC�PG�h+�"O��`A�ۛ5�y��G�4x,�P�%"O  kuV4#�fyAS�-2@KA"On���81D�4�O�a�@�D"Ot��� l��s&dҴj�����"O�xyD� 'ι��b:eٸ��R"OZ�k�I���D� :l����"O*��U�.�� �1dW �#"O���T(��Q�8`#쇝,[�U��"O:�����T��|Bvˀ�@_�$�#"Ob4�a��q�r���[�V��E��"O��B*T�8��J���X��"O�ճ��'-��zV㐖L.���"O�<�5n(?D�0�4$�>,�Ó"OH�J��� MN41�7���)�b"O�-�#��9Q�a���Y�0�r��"O<�Q��&J{��b�N�.'"& �1"O���8�P��¬Y>Pk�`�"O����#5RH���:W8Y��"O���b��b�6�c�T�>Lfe�p"O�)�6�K�&洽P[)K�q�`"O�t)��[�=�p)�`��%B��`"O0�[B��&p�����a��A��"O,�d�ͭr�x�c��&0��[�"O��9VBǦn \�b�6_�3t"OHݸr/��W�P:5(ϒi���"O@��T���u���6�
�[hJ5Ha"OP9���L�]2^p��?S@)c"O�!̃Ldĩ�"��'�x�"O~0{��X�GL�*�aۦʌ�v"OT,:M�5&����� >�����"O ����L�A J�y2�ʀ)�Ѕ3�"O~��`$Z�xS��hRDY eܹ��"O:�K B�xx�L����.dv��"O��[�FM&���l�B���&W�)D!�$�
�ޝYP$N�>��X��'�*�!�� v����9�E��r��A"OZ\���j�}(�E� 80�J�"O.���oJ=+M~4s�� %.h�y�*O�dxAL�i�������]p�C�ɯp�J���������p	�	/ZB�Ƀe7�@y�E0	�4�bH�BN�B�&Y���5˅ ��l��g�B�	;V��� P5צh�Q���LB䉝KXN��5���tD���@i�:(�B�	aT��@'��;e�TDJ��A)'�FB�	���<�Tb\�z`}ٳo�D2jB�ɸt�D��E݊f(P	ք��:`B�� j�ĸ�@� �d��	�2�( 0zC䉠C��a9Í��Ec�����$q)RC䉌T�
� �BIV�~�H��
14C���Z�t!N�bK�tk��T�9�BB�	�w
�u�D��}�ȸ�i�B�I�sZ�K�]�JI��"G!~�C�I���Yv��*x����D��C�	.Z����4V��4���8PdC��9 k�L�cBE�91���@�]. ��C��7$FI�E	�#R�����*	�C�Ix�`h�5�H.,�~  6$���B��Q�> �  �   "   Ĵ���	��Z�"w��9A�����@}"�ײK*<ac�ʄ��	�$P�h<xbK\�	"��~�"�� �"�ƬQ'%��M�Y�7�@��4,*@*dӬ� iO��3w�E�z뎔�
�D�����P�B�,�M���k�pu���ʣdz��"�R��s�a�%��O�4ڃ͌�:�I������#g`P#�ϖY��5&s�P�@�!��	5C��c��<4��n��� ��4��i��"?����D�^��4'���'C�u&(%>i���G"0�n=��J�;(0����۷tY�c��c����,�P��U��m��K�.h�8w�~��Q!Gͅ��lj�ڍlP�h�S)��`���"�\d���~���J�y���O��
=)���:��P���)Ab˾?���w�;P\�'�LjDX9_?�'R�=�W6~E^9�1��G����0�=0,�q�D�>)�
DGhj��ę>���j�x��OV��Gh8A�T����"O:��b�'�Fq��!����'˞s�MR�j/�����l��ޏ�l �u�ǆ4���p@<!RBݠ��F`���rр�M����+���u�A/&3̕���L8ڰe ����'̺�!�b��L-8�'���(Fm��1�Xʓ%�d��bT�:�b��@Q$ZCB[bi�\V�a&}��U��2Ȫ�&6}��,!� 9��ܣR�&<d�θF�r	UdHs�0����Ҋ�(��1�����V�-Q��nם#���`�c� T��B�T=���r@J�Z��O���K<��C�0rGL��%ap�p �3=Fb�	.��
�Q�����	���(�Ō 8��m��V	so�T���ߎUS�#ɟ�%�F;��Ɋ �(��B���TA'h��W��8[��ǽrP\�Z�Ąky�/��%��K9}"���dG уbc7?��柪_��]Xem��'��9a��
{Ri��ʘU��q����ַ��'�nI���ŏ,��(ь��(Pw[::�!�$�b �  �� @�?�s�I.',Tp�Q��ϧ:��)�!�@�	?r��)9vFU5h���,�`\6� "�O~�'�6�("�ې��,��� ��m��*�ˉ�Zf���)�"�u%�y�"90-*㕟����5�l�v0���	�#@�q��-��F�l���'��!�L^yfT�(O��z���6i
H��	��y�*�V�8�V�1�ФP)w�����L�>0O�O�\jT��	(       	  '  b-  �3  ):  l@  �A   Ĵ���	����Z6)Ú��P��@Zz`�B�4S���y��ƕ	#��?]�P�x�Oֵy��#�ęOfr�k����y��!y|a8&4F�B=+�I��r�,{Bօ{p����ֶ�Lx�7Oȷ1X8�F�Ƚf��kAK��n��̻�(�Qfxz�O�Q�4U�I�D����&ᏺ!�ܡ��Q0$����$.�}>��#J�E�d��K�X��pp��C� =,d+4&�%��	0&��E��,�A���|���Fa9 �Hp�����	ڟ�XwP"/�`��Q'ͥF�\�	�
��x`%J5p\�CJ�$�ȅ:�{݉�3�,�l�g'�/Z������~˞=cA��y�]:P�G+om�dٍL���^=��jCI%W�x�,\��mS��M�5���hq���5����I�MK��x��'-R�Oi2�E��ɗ�T�M���iK�	��H����g�MZ�<�fc 3��!C�]~ZqlZ*�M�c�i��'d���O��	:3Y" q�Md�s́`�@����d`�%Qp�Dܟ��	矠�I!�u��'?��'yU ��X"'��:UB�w�x�`���fq�b۱Ch����yX�����,W�,��(�����Sf�|�RA�e�Ǜt������0(��&��oV>lt�=&b�?ݬ �	��y�,ʈE,�|k���m�z"�4vɞ�'���'��O���$��X�/ �]@PrW!=����$�I@�'�(#b��v����@ >a����ٴ�?�3�iy�7m�O�l��o�6٘�O����Okl��1N`a�$��R��Q�Uؒ�2ڴ']~tb���?��Z��"�ʾV��S�(ӸN�B7ݟZ�sNE+
@���w��c��I!���FUvq���&Bp�8���E�E���y�m��\*&��7j���I_�}����KHx~���>�?���i��c> �)[�"E�%jՙ���(PC�>���p>	�m�-5f��D ta�$��$�O��'� DZ���wFБ�@�xq����O�u�Il}�'���(Jb$�Iğ�[���s�"l�Mӂ{�z H��McC�?z�*ɕ�tx�i�Qā����B̧s��8����
��A��X�h(�Z�,ɃJۏ�(I�c u�:���b�O�X�SNʳ+��,A�1a���?�՟��	a~J~���~�65P5��Q���!E�Ƌ�y�I�g͖H�����O���1�,�Dz�8�M�������YԆ��"�D�qv%rӸ���O��+2A�uˎ���O���OL��;�?1Ӄ��+|21�iY���ed�������9�Dq�e��l v�H�X>�<y'ˑ�STph��/�w)l�I��A���JV�&������4ZY�O
|,Bt/P���I�݅U�*���@OV���L�<� �O��+��~b�@�$�9�Ba�"�{��0@�!� _��e��.�"<�� +$
A"2� %oZ�HO�	�O�C攢�M��6rְ�.VTQj0
��K��`��?1���?YU�����O��|(��Č���-���ȱ�ÙgFń�	Pq��I9Uޝf��h/�	��]&:�8��$]':����(_��JgB����+F�ݛ8�B�Io�.(b�NT"�f�ئ�d��C�IA�.�1�ag��ⒹZ|9�^��#�4��3�T�W�i��'���\.r�d ��-lv����Jڛ���bH"�'4R��j���ԟ �ƅ O��ճi����ɹph��~���C"���MW;RY�){�'릥���s>��D�`/�d�' �)\f��%'D��Bq�~o�}9�ȴ|-1 Ӫ �O���'�����F�w�"M�FȒ>D���OR�A������ΟH�O�0$��'�	�4A?��$[�36r��F!8DT7�E�>H��&�|�>� �
4@�0i�ʩ���y�X�\�%�S�O��<PM-2 ���i��s4��Ys�'��@���ɧ����{$�J,A+\ e	�=)�P�$�0D�X�R7Xʼh�8E�4Xȓ�"�[�?m��hO�^�V����a.���#���M#���?�S�S�G�bQ���?����?������Ƅ<��� &���%��v$�s�śh|\`'ַm]&�0AƐ��3�x fyJ%a�7 vlhA��x�����߿csf<z!@�!$����nUC����8�$  :|c�x�(Ϥq\�I��~��'rў�����4�v�y�(�a*Az3���ȓ>�����*_�I�p
R�
�n��HO���Ol���$S���L��@L�>8+��$M�yZf� ���?���?y ��b�$�O�����t������pPAp�
�O�`�(H��	�	2�4�y��'��٠�M$^���)[�@�)�D�����f̒J��R8�q�'[�YiFI�9L���ks��B��!�z�
�=����q,DyID+Yv��J�d�!����=X��٭.��`8����K��	=�M�����$V$+s��O��۟0�a��9��@�[0"nM��i���+1�'��'*d�Yp��]��٣�֬pΚ;���J�+W璛�ֽ:'�XO$Qj���(O �˧a���=��癿H����#w�� �0�&�ۆm9��1%��>'eC�bI�'(p�����?q����kbd��O�eh|��KL8����On��d�+�����]���ځ�*D'ў����dĥh�Hic�( tA���/l��I==�5	ش�?����;*��Ob���[%}c��`�R�e&�V�L�!�V�%tp�����=9��=�f���2�S���8�U�1+��8� �ț4�@�I�m����a
��;fF�AP)��ȟ��#�癹/��)�i��cY��iF@�O���R�'�6-Ty�����=�%��,;��MB&H����d@�>A��p>�i^�LeV5�$e� ]ֶUAҪ�@�'J�#=)�O���4U1�1h#$]�$�F�Kڴ�?���0X�J�h�	�?I��?�������\T� Xp`K4٢�;W�ߣ
X`<� �aD6-��F�t@z��|x֝�|Fy�fТ�<5bNɫ9"VdKgԛ*
�#��]9����b��]9�`B�]�|�X�80Y`�Ywv�]�6n�{P̟0
{ra������ʓ|�(p��ޟ$G{��O�i�`�:����$�2lOp@��"O���(`.��$�.`�I��i��"=ͧ�?,O��#� *L4��BA<~!���f�96����v��OJ�d�O�$�ߺ;���?Q�O���A��$뀈���o�Hl�n�w9� �;q��6-ZWX��9�h���K$$Ʉ����d&޷&�B�͇�`j(h�)� K
�zRf5�<I� E!��i-�����>[��/��Wa|}x��L2ю�sٴ�hO��>�3�42��=00�ћN�t	��d	I�<���CQte�"B�����K�A}R�|�"�Ī<�'��&��ܟ\�'B����%��%1�|��.�4"� �o�>79n���П��	$W��M
p��x:�����]Z=��O��T(�kY/K�m��`.skP=��D�1|�@['�B�$�٥�Қm�iP!�	1H�*�D A���1s�[:�5�nBh݀@���]|~�+��?���O��p�G�F�y|��#X�6*8X�O���DO�]]����ɓ�l*`�z�a}��??�(� \z6.ۧ1�.���
�a}��O�m�b�'�R^>u��.�៶ٴT�4M��lOX�F���9�8�S�i�>Q��MX���[T�pf�o�|/���ӳ*%��KSvK�m�R2o
 ��I�+��9��W 5���@ޓ*Vn�S"LSEK�@���Xf��S�zm��Ҡ��e�e	%K��^��I�.D���O��S��W��ظ?3�āGh�O�|h[!˖j!��V�gW��܍�UIǍHb�����)��t�Ģ��E�nH�����ie�]m�ӟ�	�;<<���������ӟ��	�?��	�X�ġ2��Ձ"s��Q3'������L\*PV�V�C
:D"�	o8�.u>�<	�IҼ((�㥌W���\�	> �����ӽPͪ�y�jD�:Q�s �~>Y�櫚�4���@#��3f���i!*�y2�|:,��a�cyR�ɰ�?!���hO����]���6�0�l�#�\�p�B��dH����3h����cG4'1�6m�v�����'���5?�D�!A�=M�T�+%P�#V.?�r�Z5I�O����O2��غ���?!�O|"���@��V���F䋚z�� �ΠE< ���DL^*|6��^X��yS�	E�1q�^
N�l��a��ByڼAv%s�b���ND>l�ݺ��� WW`q+ґ~�������ɨ#�������v�:��EA$|�\I��4�hO��>yQ	^��\����+�h� �m�<	#�F.\�H3E-ȤRT��蠈�i}�eӀ���<�
�/S-��ޟ��'�r�fc��nfZ�Keퟜ��qnZ�0Lf��Iϟx��3fq�Qs b#B�Vp!���'
J��O�ec�g�Oԩb�(�7�A���U�\��!�S�D��C�C0��a��)=lvsdR/~-n�x��'�� ���	g�I������g�O��$/�� C;2�{��	�y1��>I ��p?��A� A� !Z��(	i��sX����O�8�UN͖F| �E[��f�S�V�!RN㟨��˟l�O�6U���'R�܅g������D�d�j��DJQ5�6��**�!����4ӊ�㡆� �M�O���|�cc7%D��"[���@4a2�?���;}D�yKS��srf�*`�"W���$[�=��I����|"�d 5��FFN�j1AƩ��?�`#�����_~J~RJ���N�!!(T��wg�7_�U*�'0D�d�ұ6��v�0羅V4�_�?}���ަ%(�	!�9�i�.!�M���?��

�<��p���?����?����?��O3f6zp���Ȳ,���&�>4k�h�ؤ�Í�F���g�w�5�g�'<��q��Fb���" ��V�N}(ӥ�.ϊ4��������>Sp�'J�(q[� e���Y�w��Dk���J)�� ��M�,и,O$���'A�A?Y& N�Lj��� >��I[�<�V��$E
�N!:NtA��֦�i��4� �d�<q4�ڻJ��(*�M�e
`�uJ��+&R�˗�#�?����?9��b,���O��$s>�1f)�6�ޭ��#
/6�Myd�W&'ɎD�Q�PWh����w�Ak��Ċ��� �P�65<q��ϝbBa�dD�O�z�20Ǘ7~���JNu�'p|���}�� �Б'��);�h����2.��u"O��P���R�S���0��"O���Ujʻd�h��M��C�s[��`�4��}�&��Ä��
��W��d���[d�i���H`(|��&�O^p��	�'�$�[�*ir�%z$ U�J�X���'��(����1~%j$��J���0�'�\9�!L\(~�"��LӦ{��|)�'��%P֬�����Oa�j�'��P�q)Dj��4�p܌��'��
/��iO�07���r�"�'�� $�ۛB�j��X�x���
�'	l�ǎ6���y!-�Y䤌��'ixq��1^Ҁ:v!ͮ\j�T��'TI@�Q� 6���A�T&�, 	�'@���0�х����R:�����'omy`ǁV}�)�dd�/8�ΉH�'��$a�] EH��7/P�eB��'��5� ;TT�M�ᬘ�
�'?�`#��#J$�q��E5���
�'\X1�$M�.�|�J,c>:T�
�'�Pa���H'?�bQ	%ր^�YQ�'d�U3�c��A�ts�m�5z��y��'\Vu���D �0"�e�'����'<�X"#�D:O�JP(s�N�~a��'S0xr���j���D"0иӓZ��D �c21X�ܚ�ś�Um���g�SB?p��AG�99F�[ׂ7��k�&�"-����Gm�(-°���#(�8�0���' �V��-ѐ��/\�q�t��m��n���j���=�h�g"O8(�6 ��t��$0��L�/=p�����2HC��J��_2s�J���ߙH�>�^�,�O�\<P7A��z��&2D��0������)�58N�jU�h@��M��ob\��lF�ve�x"!�>,��0��E�y��c�
�0=q��Q�8t�0v�IY� 
phH�#Ԃu��.�%�hQ���`�B�	\,l�Q5�ٶic���<9q�b��� ,1N����8��l�4�	(G�%�e'ǣY�±�K��`!����t�N�S�:� �-��HK"N_h�A:�C ����3?�f��).��`j� G�y 7	|�<�7A�?I��T�Ǫ��{yt��coѷ^S�����E;,j9��OG�zv��Ĝ5=��Xjs*A3>y���i�az��	��p@�⏟f��#��B���B���42E�JCF��DJ̇պ�ȡ�Az։	K�,)�l�<	C�4l��m9T���\�� �o-�ӿ	�����������2AgfBC䉨 �:���nD�p�s�Xe�H���9oF%�5	ׯp��5Q"�$�g~2/FBdȐ �'����Y��y��$P�f�:���.�|����
 /�@ �g��SN`I�v�G�@���ɤ, �LKC�Ҿh2@{A��s����dW$Y ����	љ�&d��\-���q�Ȣxf�M�� .d�-��'��;s��7�١�˿(�ݢ�y�ïA��ܠ��[�s�(�#t�Mܧ[��-� I�)Pwf$�֯���H؆ȓS1�P
co���1��،zc<�8k�pv�!�c+ͨ5�Km�4J
q��Oи�2�בU���GK��=+�L(��'cz+T��iնIe:�sٴ(�Ό��iT�:���K��(��p�ĸiFd9�K
�y0԰Y��*Od��u�ABb�)u� *�����Y�x�\�{H�DN��ܸ�|��;=�'���yB�� �n��g	ˍ)�R��`�
	�ju@�.\O4x�JR� �7˖&1y�X+po �Z�(���><�lh�/��Bw��х�m\~���2O2Y*rk���sޱ��X!��9Q1c،4�:�/��"' �c3"�z�(E��i��P�%R�  W`h ��yRAe�
r���F��y��ݧI7:�ٵ���G-�6f��|�p�ӻ{��K,O����`��Z��F�q���z���*L~\2ЃU�l�lՄ�y�@�҄�8�j`I�"ΟD�d}o� ��E=L�����̉�2���]?aK�*޿��	@���	W�
$ƤDQ`D�
N��z�
�i���@�b-�D��	wm��h�L\s� l�ꘂn���s��º6NĴ2�ض!�(�@�~jaJP��%Z�|�I# ��s�Rb�l��^�qO0q2�T �(�`�\:A�L�O��P��Ȑ5 (�L��k��'���d�8�Y�n�{�Xz���}��(�S�? �1y�oM?�92�˚?�t���y��'C�Sﰭ�I��kE�93�
Ӫ}�4u���`���7<��5C����m���?�Px�Qe�8��Uő)V+�l�䎋=j��RR�C�?���a���&o�8ؠ��YE���Uնxp�]?���!ɽ^R����C�:8�53�	%\O�x�.7M�u@���d��@ !͑/�x0G'8�`���4p�8� ��u����>��O� �%��B�@'���AW�P4�8ĀC!��N��A�&�C圱 ���U :G�����(�>�+�O?0r�D�1 �){��m�$���~�'�<<OL�@�b��>�[OPT[E
#S�+Ԕ�p|"d�<a�'4�~0�����r�]�5� 13��`��)�FT��� c�A�)Nz*E��'�Q���,��X�E��!^)�.���"��9��M4�"�P���Ol�Y�A��4���R�T���c��|+��Bc�ޘ,�a|��:w�e�A!G
B��@��i �a��	*� �B%Ǡo�z�
P�8���������gܓ.h mӀD��(!N[|c�mFzbf�W�4��~���-~�8���J�J)�F����FQ��Ø�Sx�0�����D�{�+Է Mh��A�ž?�<�Ь^�?	֌V���'�	чޛ]?�y#ԥQ�*(��.Q����ɡ��4o��9�gǏ!e!�$�(�F@3wi�#k��*C�,7�ɵy��0d�;��܉ ���h����!Q�)�Y@�F��Mh$"O���!%	�Qx�;��
?�I���C�:��fӀ�T�,I8��qO>�B&gXg�:�X��� h�9@�'$��C$��r��y��,��S0���G�32E*�(E+��Z��i:'#|Oj��׊�+P�I#dU*~<��&�I;B��@�%��uQ(��2o���2����Kv2��$f��-
�YQ�\h�<�G�<l�Рb��'?Ȃ��)_[y��5n�| 
�F�\-lѡ3�'[u�8��[t�x!钅!�Q�ȓ%�8��L�<Pi���rُP\
�X�KO����4n!��C���gܓD>�MJ"�n^98DG�$��(��z�^a�'�֢Rzp4I.bN�q�ȓ%�p�jâ0f�J��d.� ��,�ȓj� 	I�TX�2����&_G��ȓ3I2A��-O�4pҥL x�e��5�ٹ4a�-%�V� �i��E\�u�ȓ�L� *X<M�xyP�7X�j���&pq�J *� p7ϻ0H��2`+�*��1c�u�O��Iϒ؆�D�-0�d-¸-�&ʓ�S��!�ȓ	Xi ���Gڜ� �/N7���ȓ��+�NɘW��%�ĊP>�)�ȓ.��ѥ"G�����0OP��*܅ȓv�虐ȑB`Yc�	��5��xdZ��K�YϪl׍�n�ތ��N_Vsu#ץH���`WI��?�*p�ȓ.��|8�<{O0��m��>�����0�*A	���l8&�޺=����?�t[���;�V�� �1v����F�Rs���-v��`V� &ਅȓ
81Ȇ�_�>WD���.o����--Ȱ:�@�2K$�})F��..�x�ȓ��q�7�X�WG� AՈ̧sˎ��ȓT�%��f
��l9�կ֣I�̜���0��l��
�Z�A�?�@���<�ذ�ȿHR�`S��In�T�ȓwR��3��ؙ/�,�PoU+�v���U�t��~�� b��S�c˾���i�%9�j�/0�(M9g.  i"Y�ȓh��l;�"B)U�t	i�iH0;������F�� �X��ubԀ"���ȓ' M�A�ʍw,�5"�h�/(����O"��L-7�vpSc`)s�`��I�l��*�vȔd;a�,},Q�ȓA_�����u��u�J��D9�ȓ���P�C͜ouQ�4,��Dm���ȓH��8��к	^����A����Bkx����\�B�C��O�EdB���S�? ��E�ǘd�PR&�/!`��1"O�)2��KD��Bb�\�0� �"O���G�źZ�8l�sL��f
�pp"O�|`���y$"1�ʎ���a�"O$U�U�^-q�p� �	6�p���"OTQ04	QJy!R$�#c;�y�c"O
5"�������?!�*�"OvLp�Nr��	�G�42y�1�"Oj) ��ٜdP�A���)^ m��"O*$�t��?^������X��1"O�%�.V:�=
aK2S��"OZ1���R̶lCk]�NQ0�ia"O��vDزgTH�C��'7%Xq�"O �*�����Qg(f1K�"OP	��).8JUhՀ�Rz�P�"O`9tO��u�|@�qI� Z`��B"O(\��f��o؀{G
�:z2��;�"O��0�d��=	2ES0�ȗ 4�A"O�I�1��FPh���c�E���r@"O�̰"��P�� $�Q�|ne�"O�I�f�{�RŠc*Y,q48��"O�����"t���6II={m���"OF����8@@I�	?.�eCT"OabE	�C�X��)j!���a"OX��Ђ�?��#�H�Q�R�xp"O6��� M[�̽C���&=/4h"�"O*hR��Z�_*P�T K�y���r"Oz}!d�C�V�ɀ'	� }��x��"O]�t� 
eC���qeS-�=a"O�L�JǴ'ݲ��KR�P��Lh'"O�1�./��"qɋ�=̜"�"O���fN ZV����>��zv"O~�;3��|*l���@�i@0"O��ӵ��^ZxIs��1�0�"O��H0A�8aY����Ҡ�t�Z�"O�AY %*Ք��-��J���"Od�H�4)��l*1B�Aҥ��"Oh�qE�އc3|����8JR��+U*O����F͇!n����\#�����'!�(��M]t݃�H�I$�i��'ێ{��K�R��L"�eU5�V-��'^m��"��1h.E�!��17����'?�Mh��R����+��6�Ms
�'2d,qq��!,btx(�bLi	��R
�'o�z�Uku�Q��)a@~���'~8}��� ,����¦`��D��'(r��+�3Ӯ���BFa�Έ��'��L8�+U,_��܃`����'&�DRC�+�	���J�b񞰫
�'�X�M+Q�%a2P�	�(�
�'*�`�H�0 ��Y���?��c	�'k:H�a�� ��	�sB�<�jx		�'�ڱb�
�*�xQ2�ގ9�� �'��H�e�8����U�S�3��(��'�H��T�L�fSt)��<X'J$��'��|D��D�`�c ��+m��`�'@���T]�;����ղ)�'�HH��R8j���,M�NB�'��1�3��;#\�X�COG5R���'��43"��>�����rI�H��'�d1���g���8e�N�? �`�<��R?||�����&?hzwh\N�<�w��{h��h��%&��1�b(�S�<i���D��@P�H�zE�����m�<� D�С'�
Q�E��@�I�20�"O.�h�EJ:FE��d�:=0�X�"O��.� T�� SueԣU N���"O�;�L� %/X���4X0�QW"O>`aRD��H�<���^N���xA"O2͂�mW�]r�RFj�l�~m�t"O6,���XZ}�M��0(_��	HɘSlց�akR�^WA��eq�,��PoHi�I�wϚ��+�"O��4��-��U����/
�$��f"O@U7Hۉz�\4��^�x����"O�pѤ�[�R�MH�
�b�Ab"O�ȢqA�624���d�P�SZ5x""O���IP;���{�g�r�]`f"O�̨`G�>~�� pl�m�����"O��(��v��y���U�� "O����ϢV9(x�gD�%'*�x[�"OД1��7#�R�!��=0&J-`�"O�X9��յf��x��*-h�X�"Oک�%L�]��Jv	fLrA�B"O���1�X:
T��3��1(�4�a"O���j��u� ƅX��Z��"O��y6+�$M��ӄ�H�l����"OHYS`�E<�����X
*��"O|�XD��%u�d��d`��^���k�"O����  �.��C 	'
�V�C"O��*�ˑ:��	"O+w��t�1"OvЙ0J�N��m�R�˕} �}�A"O��U�!ht��)�F�2�"O��H��p��&�
�t�đ�"O�(a!P�w���Uǂ<!����"O�¤��"x�1ƌ"�|e�a"O�9��T�*�ڴb�
��б"O�H��]��j� @�U�o�i�"O�prş�HtzC��=IUt<Ba"O>�Г),�@\
�h�I�L�r"O�]� �'}�U�ThZ%L�(�""O���5�F�7��IxD!�'|�j`��"O�Y���|�d�T̀�|%r�y&"O�<���G��)��%�>���p"O���'�A�E�B�(�CAu��i[�"O>���b��dl��뇤�)8��@�"O2��˙�\6��1*�i0Fh+#"OV���hF;R�񰐊IN���4"O�2����l��`J��Sg��P"Ox�iG��
��-����V.iȒ"O2���j���M���/8�*�"O�U���7�e�eMцs��uR�"Om!�פu�8��w���v�v���"O���W*�
T`��*�	�"O8��0��8�hA�섿gr��"O.���h��MSfj��?JZ�R7"O^��ŏL 8�Zi/J��x�$"Of���B��&�t�JT�^<~��]�!"O��b��P��4)rƇ,��)1f"OY�&a�9�z;3F,�����"OB��p�hz �vE�)����"O,�Æ�C4gؐh�dM�^��CU"O��Kģ��{�8����Ԑ #"OnYR6nۥWW��`늎4���"O��a��8D�4��t�>(�q`"Od�3e��LX-h�5��*�"O�Q�5ǒ
qb
Ժ�
�<H\���"O��[Ec[nH6U��IߜsB"��"O�|�Ҏٷ
,m�� �4��@$"O� �I{�E�<�@2�k�0��I�"O|[��9N�釉�3����"O�-���	�}�"ic���%`�pSD"Oء1��'	J ��G�	2^���"ON�#E���PL��P�W[���s"O���/�.@`#El�/A�\D�"O��X�!B�%�'a����"O�eJ�+�QDL�(�L̘��"O��Y�B�j�|Ւ��7@_pQ��"O���r��� /�<@J�R��{"O�ݳ��6u*�q�jķa@�U�E"O@��U�^�|C��;�[%\�W"O(�R�Jǝ����A�3��U�g"O�1Y�![G�)��I�6 ����"O@���$V� ���斆U��@�"O�8�&��k3T�9r�W�s�>Dʖ"O����ϒ�r�X������*5�"Oq��bĢ�( 4�;�^%��"OR��f�γZS�!��e�� ���'+�V�>���أg�h��R!�8<n��ӋLq�<ab�ۀA4��J�(I���7�q�Y� �ZW�n�O�&T��	�f\�t��fP�`��'��D�ȃ]� ���KI�4Y,�B����z�p�O�����Y��y���#f5(5g	�x֗�d!��Ѐb���b��dH���e�T�1�af�V� �\,����猻��r�K޸4�fy���M�;Z �	�^���ye��1)�
B�#m�괩Dسx��E
��D�n1�C䉀(&~��3Qsq6Щ�oC�!>B�ɦG��X�����.%**��L��lC�s��Iqn�&x�+7��W�hC�ɡ��U3`@];�  �5J�#:�BC�	/�I�2`�BҘ����u
C�ɣyJ<$˒�[?{,h)�R.��B���$X	����@�F�ەa]36�B�	�D*X�bL">Z���A].p�\B�	N��7�ȋh�$d�'��k:0B�I&R��dC�;�R��VH3&
B�	�-T�\:�VM"�۳��X��C�p�Ι��Ih����n"�C�I�.Rt���i� 5� ���B䉯A�)q�� �z���⅏�V��B�9> ���e�,W4L00c�$+|B�	�n<�غ�I�&IxDLZņ)lXB��ώm�`�S�Ku ����=\��B��2FP�˕a	g`z�B�h�C��
-�HM4���㭑�>E�C�I
]�U�s��Z���Q;��B�I�,��:�#�c��Ch�	�^C䉑�֨*A.�+�E��R܆B��3v@f��5D *�ܡ�%i��oovB��C \"��\�[��A� �Q�F�0C䉟f?�	��ᗅ�A9!��c*nC�I%��]�PZ&f(�HI@�WD�`C�	�E���
eM�N����åQ>��C�ɞYZ�	��%LZE���¹|�C�	eWdԋCi@(=�$h�3�nB�	�L�b)�f
B�x�W�6sO�B�	}��b�mMG�l��F14�zB�	�(�(Y���@j�Ÿ��(4hB�	;���2ߕy(��Bc�+TD�C��^�R�(ej�If��r�	;�TC�I(a��`��w�����	>�B�I7�r)x�c͖B��Qo�!/|�B�)� ���2��>=H�5�5M��E"Ov):Dh�
d��Ѱ׃0*L���q"O�l���4�MR��T,9��h�"Ot����֩v�T�[��Aծ�1�"OAP�$��qt)��lЪy����"O����A�46�`��@�T.5��Ӆ"O^�۠b�/�zӈȑ-���j�"OR	�BM�f�>�3���2e�q"O8���7�I�Rf�f.y�r"O�yY mYa�8-�#7~��Z�"O�q`Q�G�]C�I�P.g|�I �"O�=@ K�?#�6�Y�J����`��"OJx����;�r!�$�D�c�:�"O\�bf��2z� 1�@1Bq"OTuU[-h[��0g��@`��!$"O]C�oY�S�\��p�ۇMԻ�"O����q�8�K1G׺C�q�"OȌ�AR�F��!���8I��e"O��R�#)B<e(R��Q�<�c"O��ڤK��;�¥r� ݤ�H�7"O�y����i���# �I�"ɤ�Yf"O�I�&U���`����	���"OpxX��Q(_]*�x�n�� ��) �"Ö��'P< �<�,���H��"O�Wh�1x�ڡ+ӥ�z��!"O8�ڂB%3T�h�D�9�H��5"O�
ԯR�<��}�a��J��lR"O��F#)G�J)q.��A�t�"Oź&E�.C� D N�l�W"O���6����
���M�4~d���"OP4(�k�>r��0q	�#��
�"O\���l�[u�V#2fk�!��"O8�p"nV�z<)E���ZG��B"O4�z�k�k ��R����&ab��`"O�qy�
 �O��!f�_!z�X�"OF�Zw(��~�T�j���z�$�"O
=cB`��%����f!�*�в5"Of�d��z+��_��"O���7+�>�if�-�@�J�"O~���&4-/�%��fЦm����"OvH�0 ����`�^�q���#"O�䟁Zx�Ep0f�d�"O�����
� ��,y`��Q�H�G"O���� �`aRQ�c�:\�"Od�8��9�I���Z�W���"O>0����*Q�ܛ�(�G e�U"O~Reǋ*x[�t�ҭ@.���"O�Y��^�" ��#D� �>@2"O���/�93�P(7-;|�m��"O>@k����m��$��f�_���"O�� G�l���Z�DՏJV���"O�|yR*ߊiںEÅiٛ W��r"O�\ ��$1�Z��#��0S�~@3"Ol�x �@(�R`���l����""O����ɞ�N`�)``�pu�k�"O��(�˧_��x���рw*5��"O<]J_3����t�I���@"O��@�:)�Hpb%�8k�h蚴"O�,�[�z�=�E�9�B��"O�5�eZh���#����X��1"O�D�AkD:y]����V)�h�Q"O�pxa�î3`6���ީj���H�"OĴ�s�J*9�b�Y⼕J�2��7"O�B2l��=0�+݈0��eQCB.D�� P-�i)J?~8v��53���h"O<Y�D�0�½e�jl)�"O�����ƫC��#�熏.��C2"O<Y�כz-���@Mt���"O�t5Ov@B�R�ݓZVu�s"O0�+ׄT�A��}@���F5s�"O����� v�� ��ԗ
��"Op�`��Ĺ*�}�F�|�d c"OA���R�G��(�!U�L;b@ce"Ol\S��)^�9
���[$*xhB"OP(����Q�zx���="&p�	�"O�M��
  �   ,   Ĵ���	��Zc��4p�����@}"�ײK*<ac�ʄ��	�$P�h<x�� �	��6Mƍ`� ��d��>!<�H�Z>�X��QJ����CӦ�4��u��F� P��]Q�������?)�����"CG?t�|���O�>_���b0c�<�3�
�W�Np@��>�ծ �d�����FW�D�ɂ
{�2�ʑ{ʖ���%�u�.��Ja��ڇ`�-T.�Fn���d:I��P"��
�n|�ɺ�MՏ��F�W H�ħb���@O�R�"ݛ�nܒ<���s�B�X6��9M�$�W�_�^��K�\�u��96�`���~٠��F�+	lāzBۚ(��I�&/��17.ң��DA1O�m
3�Л~�$��?�a�+/K�,�5aֺ�`]���ƽo���a��|�*_�i޴��x��+�%���d-��A�	*�*#�R3��>8�ч✪�'m:�����U�;���c�C۾�:N_�3�����=N��9��O����`	��g�<����Ti��[$X\���a��6���A�W��$YI�ʓ�PF�.��M]���J8^
|��a�~ep���-=<$�#�'m8��I�k�]a� �!?��I+a��k�d����%���v�G=L��蚠�+Dt���mL��L��
�*>���O����m� &���tD�H�`�T.n�"0��Øl�DL�t u� ��q�$�<̴ "� �Ϧ�� J��&���Ů��XT�q#� �<IqHɷ`u�Pa��j�I�^�HE��9.���gJ�5A��I*���鲚x2)�hL���0j	�@|0�@dF�O�h:��J����ӈ̷;��`��/W��L�!��	�<��`��(��N��d�M��8~��x�1�H�^anm(���]y"��M���<�D�
s�]X�		bmNh��Ґ��z`#�)j��� ЏfꌓOPa0���N�1O��0���4T�}I���Ӣ��DH
8:TC�I0%��  �?����y�$ |�X�{�h�'^�JY8�A��y�-H+
܌#��J�k�A��y�_q��L��!�8u���&ė��y�Ȅ�7�&�ڢ��ԀA� �T��yb̛���� r�걸`��7�y"LU95AV-�DI�oOJ`�S��yr��p
6���b�t�+��.�y�-I\i@OǸ�Mɳi��ybk�5J�
|Q�È���   �  �  �  =   �+  �7  �B  �M  �U  .c  �l  �r  Ky  �  ؅  �  ^�  ��  �  (�  j�  ��  �  3�  u�  ��  ��  ��  ��  ��  ��   � O F* �2 �8 ? cE F  Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�� |d��"O
`�(�;���8���-0��1%"Oj4��ND^[��"3/9�0|H�"OB���H��*�ʞRy=a"O�味V�!X��!&F�:J�$���"O,��a
���C�Ą�M�"O,$3%o�-���p���+Ն�:1"O��ݢ1����`���y14]2��i�<�6��{_���c�H�`�fX�$Kn�<��A̼VI�xR[�)�Ć�pඤ�ȓA5��('nߡ4�� �)˩%� ���,��r�؊b#`T�eT09���ȓ!�b��g��}�8�F��-? �ȓ
K|m�ș�VṔ���2�%�ȓ"R�X�j�4JN�1�˘X�i����̹	_�jZ��1!g��zܶ��ȓgil,*�J�
j�Ne��i�J%b���f	�(U��:���G��$Y^م�~r�� S�%T"���k\�jx�ȓ|4�1�îJb��@ӵ�ݩn�V��/[`�"�v4�R�!ʎ<��M�ȓ`:��z�ؚh�J�Z��$HY:	��H��p�m�C1��!��B:��0��EnjZA V;9����J[
2���	��4'J�EA�IVW&��~�(aZ��ӹ�>� o�Y�|�ȓ�f�A�
Ο7�H��M�$�����mޠP����/���ANXo*�ȓTv�����{ ��-7�*h��I��sB�8�8���3����ȓNe*M�悡;������X�o��!�ȓ'lj�#F�m�+R&;�|��2)n�C��0S4���T:
b���:�0!��e֊��)��ͷV��,�ȓ0�&�8#���� ع�L�����;�P�AFd���,w�6d��r�EQ�( �gVlɦ�M,H��,DP���|�I	$G#\���ȓ"�)���E�B	yt&B�^�LɅ�4�� ��eëF�ڙ��n��R�p�ȓp`@}bŇ�=�$�AUN��P����L��p���_�a�)�Y�!��-��u�5���o}�`iF�@A�p ��F�\�0��[���IF/5���k>bTؖ�;K'DT`�^��@��fnV���Y�b�lI��	����ȓ,nٛ��Ć3���kC��8�m�ȓ'� I ���x<=���޳{��	��6��(� N�����
�y2<��ȓx;6q��I�
=  yG�O�,�!�ȓW�>���.؜ɰB��;�����`9"�ˁl�$@��- G��D�ȓ���zF"� ~\�`%�[�ل�E�1�N�;f��P7�.
�T̈́�4 ��QS�[@��o�|h���h�c�A�,#p�+1�֧jN��O�l��Yl�=�QO����]RB����`���T�	�<��A�]�J�@d/��y�@k�+Ye�<QQ��&X�1�U, 8����L�˦a�>I��T>1b��&8�<I[v�"	!L�1��.D�p���̤A�����[�s��<"!)D��P�O�^	*��D�,�1*B�3D�� PQ�WjF�=�$��F�6t����"O�˳d֨l����6��������HO?�ă�Psf�zҠZ�9��I� �Қ��䒡qx���U)�}�e�O�fR�B���"�aX	JT��
U- ��s�E"LO�㟼!�EٴO���]�+7!��f��5�B(��([����!��(w��A0������h_��Py"�I�5b'��L�˳jݴ�O�=�O>^0�M��Z��3�k� d�ɺ�'&x0QkҊ2d�����K&�D���'!�d� l
���ä� 9Z��!�$�]'�=��shA#�"�-?�!��7{��d愨thd`� �&�a}B�>���5�Rl����%?��Y���~�<av,�.�Q�"�ݦq�81�#z��?�"�'lDUIE�E>�h�E��&%"��'7R��V�W	f�iS��_7V�]x��<��4�2ǇT� -��ŵsJ.��ȓ���
T�& ��p�ӮQ���F{"�Og\�ræY,���`�:c\�q��'����B6QF(S��YÊx�ߴPr֣<E��4�EzVM�V}0 ��F/�8�ȓ
�j�-�v�"����:�����b����.IL6�8�h3oX�� �	�N�p$�L2e��X�vP2��Գb>ṯ4f$�D�b%F���J�X��L�t0a�V5�~�x2�)��WO�����)�:�d�ڴl[q�DS_���O�MR�0���"wL\�>9��'�`b� �I��=�R�4X��Q���#�S�䎆"h9Z(R��C�=�9�.5�yB�@1sَ����D�̋r�^��Ƣ<���Ob��k��j��X
��-�d��3�Id�O����Wc�mw�9�d��M4��'Q�b�^8-^�؉@�yE�B ��~r�)�'Hul0؅/X;q�fc�Rt�Y��z�YWkVfn���'q�n	�ȓ~�x�b&f^�0�J%!�y%����|Oh�K�DӢ��Q��H��Q�ǰ?!�+�]��� ӯfsB@"ccr8�@'�x�eICq�AS��3H��Scn�<)�I��?qI>	/O�'>���:E!O,M��� ۜa�$�Fy��"�S�ԡ��=6�2c/�<�������Ķ�|��ɀ�jMsɅ�[�t[RE� Y;����)v�l�05�b�8�� �V��C���`T����'��I�h�>��TH� J�JmZ�ažC�<�IM؟�[F၏ry.!RB�H���G3LO��$�V��-~�@hf����2�p�L���m�'$�<#��Ԝ#���Te��AZ��$�>��?j�"d�Gߏ�x��#��R̓��=�A�{���'>�Xy�%$�M��r�$F{J|
ŇG�r���P�ʛ0Z|��&a�A�<9�,E�/�D�irL�P^mZ0Gz?!	�;�=+ �S-8pi3c�WO�	��IA~����u˔�>"���Pg��y���62��*�C��P�A�m���yR��&8 n�37H�*��p9&��y��%2�Jĳ��T��i&����'�ў���'�ke�R�`�"T�fl�"O޼��,�8j�J�W��0�E"OT]���ݢ�0�Xv��a1jL
�"O����ޥ��4��h�3E4R��"O�������C*_�y#�D��"O�X"`n�����( ��/���1��0�S��y
� Zh�3O�p�n��A��&w���g"O��
�Ü� Hb�����"��Y{�i�!��A�h�dԋWkL4k(Tt�4�@%��=��y�Ƙ,��(�c�6\���K����y`V�z�.ղv'��X0��	D����I�d�����Do :Ĩ��挊Q��T;������ў�(O��.��g�`�C'�7 �F��b�Ϗ^��GzR�'� `4�āP[�iH'��"��(�N<�κ��E{��n�k�a�.j��a���9>� ӱi��}B(�ԟ(RtDR7���ˊ!7��5ZT�#\Ob�����Z<��t� ��=]�e�I!D����'�8].X�P��E=K��i�t#:�I��hO�O���Y�唭,�"�`�/��g�`4�����&ɨ��5�Ҡ�_�x�`�!�*����o���p�܀#P�h�O�Q�"������F{��)T�/�*��'�
�s��=�e��
�"Oxع�#6� !UJRLt�x�"O4C䢎
y���ㄙw5 9�6"O���%����EX�~��	@"O�rB���b���A�ĕ!jQa�"O���+��D��9W � l��z�"O<\0�g�8eI�k'�H;wm&� A_��s�Z�"A�D"+\׌̂�������I_y��ͭ[纘�Vk�B�(�A˔7�p=9�}2(�%B1�`�RC�'z� A���yB��}�"��X<p&x:e�>�y�	��I�T]9"�N:O�%�$��)�y�#�!���R� �	�RJѬ��yB #C2��2��6"y; g���y�&��l8pM��䬄"e*��y�M�g;�����2�bls����y��ʻt�=�ȍr�6l�`˩�y��+d,,ȊDb�0:&�1�ɫ�y҈צ#wm�%��9t���CA�y��X�kmz���)W3aP����G�7�yRF��k�*�:�aN����R�Z�yr�K�p19��v���
C���y"�A8B��}°c��s!୲s�O�y��J�*TJ5�L�N�c+U��y2���wk5Y�n 
��Iܢ�y���b���x�!���M�B��y�M�E��`�ճen���Aܺ�y��Fy�2�ش��0y����U!�y2��M]hᨦǟu~��3�ģ�y���4�,��$�/m���!TN�.�y���@h��P��X�^�|�ڣf���y�B�N���S�jIG+�fgY��y"��ax���f��?m��3t
�yrb	�U���A4�01�"�0n�(�y"��=R,�تT���$��Җ�W/�y�ܱ�� �F��֕���<�y��N��fFO����:e��3�y��ǋ9� ��|��| Ģ ��yB�¿76�!��Ɗ/tP���cj��y"d�.\�����:߸,!pn8�y*� 5n(H�Ȫ9���Ѥ�L:�y(��Q�����0��T{��'�y��^��(���Ҏ=Z(�2�L��yʃ99�Qإ��_�� ��I,�y�+��*`@w� $_���P矖�y�j���v�W.�V�81R5���y򠍃p6D��E/\�Q.dIu��;�y�eG&.&��3�JL<���y�N	/x�6�K#"A�2�R�G�#�y
� 6�i��J�rW��hQ�):0��"O|����\����� E���h�a"O��eF f||k�R�<� �"OZ�B	å'J�³#�5�4��"O���J�-d�&$0�ٿo��`��'���'�b�'_��'[��'���'�(<itǞ�Uא� 1�g�ֹ�3�'x"�'�'���'���'���'<~|x��A	^��t1��%B �_���蟄�	Ο��I՟�������I��X�"	E"�	�ό<�87i���	ҟ���ʟ,�	ß8�	ϟ����ԩ����A�89�C�$Yo,�㰇������I�0���p�I�@�I����Ϩ
��$Y��p���̟��I����۟,��П��	����˟Ha�ˑo{lM��(DM>���M͟���؟4�Iџ��������ԟH!���aAbC����zL ��e�֟����t��ܟ���֟��	ȟ ��˟t!�N/#�fe�H�)|Ƙ�����Iȟ<�����ן,���������PI��8Z�#���4`�x�養Pǟ����� ��؟h�I��T�I���şȻ���{�2rG��Zg�L��g ��`���t��՟��Iן��	ԟd����XaFL.<x ��q�����m�ǟ���韼�	П`��蟰��؟<�Iş�:�	+8�f�:G��C[Dx0V���L����T��Ɵ���P�I��M���?�M�"�ZQ�B�=\���H�\��ʟ8�����$^̦A���R*��ىz윪&ES�Z-����f�'�ɧ��'��V�@�v��M�P0��/{��E�Q�nӤ��EB�Z6�??I`�p$�"��1�doW�n�hu`ѫ�5%��:7�݋��'$"U��F�4��<H�� �G"ݴ/�Ft	7)�:�,6-ݝq�1O��	;�	Sߦ�]�A pn�0��l	��L	-Ā���Mۘ'c�)�IN=R.6�`�X�u��FPZ�N�f�5���?�y"b6�x`#�/)(ў��՟�R�mns�a�d͉�tV(n��$�<�J>	r�ih.�R�y�k��
:1���!��0��oQ2c���|b�<Y���M��'��ɍ@���y���E�\�s
C��Z�:(*}1�C���|�`[�uw��Of�$Ä>.~��G��|S^�хH�<�-O\��s����|>�� ��!��(s�xߴ����'�L6��Oh�O�+8�i{��	�Eׄ�w��7��d�O
7��O�;�}�d�f|F ���)l�J�p6`	���xc΂�M�f �\u|P�� ���g��>|>�iF�+�F����=f:@S�d�@M�Y��Ș����ㆵ8��Q���K�0t|�l~R��*cI�W�4A�ł(��)g捣,����1�L: ���H�)�H��$��X ��6,O;\c�4�oUF�.�)E��g���cu�K89�U�EkT�L(�Lѷ.J5@[���c ҡIg&-q�gV�1���j� z��;7��	!�����
�>١�߷e?�M�b]�%�FxP h�B�-����d���C.x:f��*0t<��*	��#W�Yئ9����0�I�?��O�ݠ��R��0�i��4�v sV�i�"�'	&�s`�'�"�'#2�Ol��5Fa]�_���dʍB��@�'��nڬa�x��4�?���?y�'{�������zR|�7�_.If�� ��	�.�:7�0y�d��?���'z��'\R��������q��;**�<��t����d�Ol�8fCi�i>���Ɵ�!t���4���ʍ43Q���&A�.����O��$�xu�	���I�@�I���f�
9��Ss�ZF���4�?��@B�	i���t�'�W����	�D��	:��N%��mjdB���M+�|��'���'.��'���z�,�wԿc��X��ǲn��"s!�(�ē�?9���?�/O����O&�Cv�E���<ۃ/L�O���(T�0�1O����O>�$�<���.8Y��£W��o\+�U1�@G'3t�ꓶ?)��?�+O����OD�b�T?�'�Ѯ+�,�����\ePH
w��>9���?����Ƌ�&&>k�h"^��0�ō?T��P�Ր�MK��?�)O���O�K�I�z������$$�L�)҇=/K �nZݟt��iyb�X?C�P�N�D��k,�����u푁y^,p�@��\���R����ğ��r�;§�n��";b��7&ӈy��h��Z1A6M�<q$b�ԛ �~:��"w��@[b���ȉ�(�*pZ1��}ӎ�$�O� �V#�<ͧ�?i�g�	Z	z�Z���!M��� ��5
�7�_0^Ă|l�ß���ß��S*���|�k���\�6NE�%9�,�
''ۛf�;&��П<�I�?c����OU�
F��  �����A�"�v]�ش�?���?!�#����T�'=B.�:!�90�[X�L�{���u:D��?��.&��<���?���V<(q�ר.�1BdB�=2J� ��i&СA`JO�	�O��d�<!qDZ�g��-av�ŋ9�8D�	�ܴ�?��"NA̓�?����?-O&$��B�/i��|���R0����т�M'd�&�T�I۟��IPyB�'l��֮|ZH|�	N-N[ T:�,�8����y2�'�T�h�	�(~���.1}�f'@p�ʜ�3l?��%_��O�d2�I���B��7MԮ+~�y��$_�Y�R<
��	�H�	Ry��';JA��[>u�	�����Q��8Qz�{��s̀�+ܴ�?���'Z^i�WB���mb8TIՃN(2&pE�2�LAo�����'����6����	�?1�RGR�Hd���2��E�J��6*���'�čY��l�y��� �u0da����c�gÊ��@Y�@�ɽkR�4����<�IƟ��gyZw���H"��|���K�D@8`b$��O4��B?x<��������%ۂ�I�&x"�AZH��V+�8c 2�'�"�'a�Q��S� ���)u��A�g_���`��J��MK7���7�
�<E���'���0�䈟��h�,��B���k�����O����):��|B���?i�'�2v�!"0��ܟgRb�#��>�	�NxI�K|��?��'f�2�"�نݳ�
�Gn�X�4�?7�3����Od�$�O��t�Gː�w���	�~����gF�>��"17��	�'���'H��ٟ �4с�����U�l*P� B ��Y�'���'b���O ���M)�Q�F�1h���F��(Lb"i	�������Ж'C��Q�U���� *�"��&�L&z���;�+I�*0���'�R�'��O(���5T=�÷i���[R L�h�x���M�$8�� �On�D�OB��?i����i�O�-�1(Ԝ�J3,�%	�U����¦�IM���?y�)A0i��'�D0T��!z�՚dm%!�:�Z�~ӄ�Ī<���0$�/�����O����8��})�/J�Z���v�ƃ$F���>��Y
��� J�@�S���H�0�� �'��jh�d�7H���$�O �cF�O|���O�����F�Ӻ�, }�l�� ��H,�fge}r�'.��A����Ę��O�&L��DɺRJB�K�,N>g�4�ڴ$������?���?�����4�z��G-L���`�� -^DlXEAA:h��l=`�`!�S*4�)§�?��"Й1rt� gT+N���E�:�&�'2�'#�P��R���՟��O?���P;P���Z�M>=V�����T�1O��tGOt�П|��P?��#h��0�i��'YB���S���Ʌ�&��'���'v�����
�/3� C�'�Av�I%}"�}c�FΟ�	ğ����� �'J*��g �1�P(��b�+{�	ߟ��Iğ�?���I@���/ǧG,�\+ퟍj�b�s�Ҏf���'��'��	韄2Wj�kz�i�1���1�;�8�S4,Sߦ	�Iޟ$�	C��?j	 3���m(D������i���sš7,����?�����O���|��!�d�2�>�y!��zMU�u�[��M+����'�ҩŮ���K<@� ;]LH�7"�L(��b�Ѧ��	Fyr�'��P�EP>�'��T��N�����Y��PR���#�2b�h�	�[
e��%�~"�����x#�+��7�]�g�S^}r�'�����'��^����kyZw1�]�0O�'j�����8popj�O>��L��8|�����
9���v۾0��(񣬆�*���G�T���'w��'Y�TY��ǟ�ȁc��A���jS�I�W2�[��C��M��(�!�t��<E�d�'�]$!�%@�0�0A��RVm���tӤ���O���и
����|*���?Y�'�\}8D�)��� �@Ց��ӷ%*扎p��,(H|���?Y�'��B� �>/`�ٓ#P�F�aߴ�?�S#į��$�Ol�$�O����S-�;o,	*��� }����K�>A�OîA���'�"�'��	��N�0�zث�s��Q*��R�ŗ'q��'i��Op � 
�L�Q4�S�SfM��Hl�}[��������8�'�o�������4�F鋗N؄̒b$�]�Y_��'�b�'��O����?~ט���iG� ��Kŵ_��tJ$�<i2���O����Oʓ�?sO�����O|k�M�61��
5�օq�*	�����b��yn��c�*e%�p*g�Q�$�v�C���m��9�S.a� ��<��?A$��)�����OT��#&��u@fj��3c*���0M�T��>	��#e��� �FV�S�t�B��T(�V�ڠh�x0H2�S��d�O0d�5c�OV��O�����D�Ӻ+$)��dJ�X�i���Z��o}R�'4�|��B�����O��*h�@pÂI�Ycm�4�(�r��?����?Q����4���dQ9`i��X��D�Cb�!B^4"*z%n'�`��'?�)§�?���Kg������� N�Mj�9x��&�'r�'���J^��П��I|?�E��vG(��#m��Rnj!�h�##�1O��r�.	ܺk���?)��?�Ӻ�en�6-�Pn��X����+a�νm۟���[y��'j��'~qO:��@�'!��!!��)6�\��CV�,���&!ж�?�����D�O�|�2�ԥ-�2m�`��_�<=:��G�$�j˓�?����?)���'�A�%b&-n6!B����,�ބ��nY�Gݘ�)�Op���O˓�?��ƞ��)��� ��Ǭ�b�:�&�M���?����'0�G�	y���qڴl��\�F�@�8�rHbbL��,��'+�'1�	؟L��n���'g.�Q��0_�PA�!��&rv0�@|�(��)�Iş�h]`�s�N6��ř$�x3���8&�$�S���pƛ�'5����XR�T�'���OY��2ND9<�V��Ԫ��W:&,�vk+��Ο̐1�ɇnc��'.b�lS?�����8x�'���+W�B�'T��'���^��]�yJdJƦҊ?@`hwH���U���������e�>�)��Z)lݒ�*$nPa�����7��\�hm���T�I������?��蟰�I[h��
 )O�&�l�oѣ.i��޴LN�8 ���?i,O�	$���O�� ܡk����`��8��ې@a�mKc�i���'���>j�J7��O~���O8�$�O���c$�2��͂IMvAHGkW�
��V�'�剘��)R��?��c�8�N��p���S�d�&[̩#'�iOR��yR�6��O$���Oh�DR���O �b�@�;s�Z�QQ$��>��R�i�U��LF/�]�T��� ��Ky�ϐs�	`'�� ���Ӂ%тK% 4A��}���D�O����O���O��Iџ@Y�BA�O�B,
�%Ğb!�,�O˻xJ�(�������#.JU�I��O�$\Pu@~�}z�8aFJB1�8��-Y�`�������������UyB�'s�)��OQ����L�c�$��s$��*f��!�f�4���O��$�OF��O`���J{�>�d�O&�م�Η:JZ�u!^w"`,3 �AƦQ�Iϟ���syR�'
���O���'�@m����1'kĠ�b�­E\a��.9p���'�B�'��{�q�����O��$���=���Ժ
5@�"�@LP`����J\�����Wy��'�d��OW2�'����M3���:�b@�#jڼ!�����f���U�	̟�Ԅ�M���?���b�'�?Y��M�<d�x���5Nf<���G��ß�'���|�'�HaB�O��'3Q� �3�#lQJ5H��Gg{NUo�-z��i�4�?����?���*���?1��1@f|)�^�2�	��O�/X��T���i��Q�B�'��	0+�@�Y�S�?�
b�4�FP�Q&��B�T�k�a� �MS���?i�L��7�i��'g��'�Zw�X5:�H[��\i��$�v�tջ�4��}�
-�S�4�'�B�'�� �2KO�3qn<����BN�� n�v��X�@���l�ӟX��쟐�	��)��bc��/j�`�Ez� u��a�>���<���?a��?�����IQ�.��j�'T+vL*���+)m��X���	؟���؟�í�>��?4g1P�h��wL��A��uX򨀹��E��?��?1���?�/�>�[����:t-�p�8H3��tEV4*��&�M����?)���?�����O Yc>��h��i��Y���� ��������I�� �I͟�	̟�{*$�M���?�!bЮ(�2Y�$ل ~��H�]p��'{�'k�I̟��F�a>���n?�qb��^�"T/ſ%2^�҄���M��ڟ������Ų�Ms��?1����!���a�r�JB�T	w�(ˇ��3-��&�'��	���sgu>��	{y��MK�n�״	�v�Q�Tz��bj�i�����9t��M{��?����'�?!�CP��l�w��4j�bM2$$�#������q�����$���a�IM+Z�p��TW�|�{��]�'8����i}�6-�O����O���X}�V�0`N\]����6y��j$���M��H�<9O>��T�'R|��\����f�n7`��na�����O��dP�  l�ܟ���ݟ��	���ݖ	%d�q�)ǜh`��pRɈE��6�O4˓<7T�S���'P��'$d�CDRi)�*Bێ5TH�c&xӊ��J3TJ�m�'m�	͟��'lZcN�8��'&yP�*ɉ����O
��>OB���On���O���O��D[�
�y��� ��a�E�M�rp� �Oئy�Iߟ��	֟�	��˓�?�FC�fȁUb��px��{SJD@�'��'.��'qb[>�em<�M#a&���J���Ǔ,RZ�� &*����'XR�'�R�' �	��Ib>��kV"4ˌ�q �˪qn\�����3�MC���?a��?qfQ?���h��Ms��?	��J�r�(��ƃ:i}�����	#7�F�'12�'��Iោ���r>��	[?�T�\�d'
{!���W��bGަ������'*0}R��4�i�O���^�f��"B0܌;�i�p7\�%�������
Пl&����je�����
,*�s���h�mZsyB��8�6M�Z���'���!?��7#�" �5��#5�%�B�G��e�	ğ�{f�'�S�'���&�9�UC1gۧp�nڷnٺ��ٴ�?����?Y�'I6�'9��9WG"h:���0P�xw�P�S�B7�N�<���� ��S�����=&TX�S��#P���iB�MK��?i�Fs,q��x��'��O�e��΁�rq,�$���An�ѱ�i��'!�,��c-�	�Or�d�O���v��5~8u��(V,���ǃ����I=s�UM<���?)J>��]nJ�0�N�4K^02��ׇ�h�'$��h�'����(�	Y�Sd����Hk�d�Qd��1$l���!���?������?��n_:P�k-U�@(R�[,q4����ݳ�?Y-O��D�Od�����`�|BC⁨**-j�.1�*�Ya��@}r�'HR�|b�'I�탋�y�@T�j�x�� jO�(8�䃑�J�����?!���?�.OxX��ZR� ^cXd ���x!z���&ʦ4��	�4�?�H>����?ٴ����'��1U�,T�)�ND�+�x�ݴ�?i����Ȕpx�'>��	�?�1gO�k�R����1^m���V����ē�?�h$�3���䓃�T���#pP��C>Y�:p����?�M�*O�]a$�C���ï�������i�'�v5�$)]0������(Se�d��4�?�ooH�������+sM���P��>U��ف�@��`�J6�,|o�� �I����S=�ē�?YRE�Mt}A�lF����iD�֮��	2�|����O~�3"�:��i@�I�#h�@2�M���������	�1W��	H<���?��'�@x"��Z
?ظ1!7�T�%��I��4��lT6e�V����'��'�H��B�S>g�=)T��,<�T%8$�m��d�
/�:q'���̟4&�֘R��aE����0�RI�z���@�`�����$�O`���O.˓%[� �D��AB!���@�U%��� Ǯ�'|�'2R�	��@���2mk�^�3�v���ɥ=)�X�������� �Iҟ���˟��He� n�6Nd��B�~���YwK�ঽ�Iɟ��p�	ɟ��:9&���C�cӖ�pR;|y��
vLjpQ�Y�$��۟���zy"�$���� ��FB4'��� gFR� �0��[����I����?13Q�"�s���-g��\▆�8�o����Iޟ��ɪHZ��	ϟ���۟��S�a$��/u�(I[+s6<%*���z�I��|�	
a��%��+�~���+*��A�#}�D�3w������'�����|�ؘ�O�O��sK�9v��>
|�6��214Ҩm��	�nU$"<�~���_�m�ٱ"R�v8�z����Y1�6M�O�d�O��	�]�Iʟ�J� E�p���a�&�ID@��M�"�^s�����K8J��Ѝ޲ 4���ێ&*�8n�ȟ��I�c�����ē�?��~����V� �oY#A fԢ��'ގ��y��'���'OF�8��],)��!H *G�e�����iӴ�D�"��$�`��� %���2h���a��",�
l�H
f�z��.T�<���?q����] g��l�bP0=�ni��4�Fnv�Ο���b��Ο��ɚm��ڇ�^�'.�x2��·D�1�N(���H�	�З'��h��d>�p����H���U[Md�>Q���?YJ>Y��?10�]r}"䔝&`Du�E�'4�8X0�b����D�O���O����O��ҍ�O.���O�4��D�Jb�YdoӕWl��e���Ih�Ɵ �ɞ/gNU�=���4@� ����P�Ʈ��M����?���?I�,�9�?��?�����M�"�h<#r�+G&Ҭ+gk� q��'�B^��B�&�Ӻ[F��-O�hG,�$I�Q��#���M�'��-12�b� �$�O������Qԧ5���V��ل�E9���m.�'��GҚ>q�G��6���
̍TZ�3T%S��}��#�֟d�	ʟl���?%�',��B���(��|�U'�&q[���O~���)�����@�E @��8 ���VE���PT��M����?��Wp�����?I)���䠟h��.2^�"%I`��1�Hs��D	�O�a'>%�	П0���txZ���&��-v4p�4k�
!�4���4�?�w@OR����d�'���>�df�8j�=�f+E<��4��q}�Z��'�b�'b�'rm�w�~�a��~D�|0��$/�pi'_� �I��`��x�	��d�I�-I�u9F/Y�F,�����9A���(�ě(l��?y��?�*O4U딍��|�%�����P)4��0�� �ƐM}��'}B�|��'|�����Ȝp��BjA�
_�I*!g�<V��Ɵ`�IƟ��'&�}0ӏ+�	�=���Y"-)�21�T*����o�ß $����ß����2��)T|�@l� �fLj�
\T�7m�O��D�<A3�H^��O�B�OD|Q�qC��N5�"J�ul��{
#�d�O����m��'`�Q(�(�36Ū!ÑNO�?M*�o�ty��sԼ7my�$�'��Ģ;?�b 38�B�7l��u�㪗����Iǟ����4�S�'+ ��Q���|dzdñ,ͼ2�xo+v-�uJ޴�?A���?���2ʉ'�m׵:�����9�����큶t7��3i��"|Z�$�Z�!����'�dJeꇢn�� q�i���'��ܨOP��O��ɭy.Pə��Հ,���#;�c����b�T������T�F�&�҂+��<@�ߛ�l��ߴ�?�  ��[�'!b�'�ɧ5�#�/f�@Ēn(UlxK�.�!���q1O���O<��<��L
cJ��(G�#N��ɛ������x�'^�|�'_�fϋP�Xh@(��:4���	V�] ���y��'��'�R�'�*ԡ%�'��	$nUK�
�@�GO� /�H3g���D�O8��'�d�O:�d��^r��	�co�pP�� {Ԩa�Y�;�$���������Dp�4XQ?1�ЇA;����ǣ	-�:�6/D��Pt.�4C,���'M1yI�;bŭ��kQ�Ǽ[n��bޒ-`Rh�7(��aT�[%Ǜ;*�ȝ�ä�+a�ds�&�d=�9B��D�	 �3�C3xʡ*e�>n�4{��߼�Ԅ�C!�XE>��I�=}�}��H%! V�?67\�7�X�YZ��I
1�eG݅Jh��B,�0������}�(�2lլ�z<��ğ,�ɳ�r�)6���K�$l�w�q�}siI�T�ڀ����D�<p�����!��O�`��ӟl�hSOX��Zdg����M�s"��&�V�x�FֵsvQ?����θ�R��9[���p`Z����Ba��O�wӤє��'��.Or,a'�	L�T��WD��0pG"O(�rϓ�*���"Dۙ}{x)�ɐ�HOxUmZş$�D�I�2���v�
n錝;G.�ϟ���3�J�{"K�����I��x���ug�'j� 'T4�ԅ����X�t΃#��ċ(q46p�Ꮖ-m���y��hO���g�0p�D8q0I��6��A���Af�{E�D���*!��(+瓤G��� 3�L�&�@��q4�a�@$D�/���i�	p��`��O�pq��'~�Py��/yw��J��A&OU�)�B���y".��\A@��HH0A�p���-l"=�O��I-��C�t�? Z9Q�)�=H�:BW�<[CF���O���O���!@DX���Op��l,X�z'�Q1���;��	�6�Te)��_�I)H��2��%a��H@�;O��3�d�*��b$I�:w0�	�f��;c�|+G�)�*8R�V+_htz3��;��Hu��OXl�8V^Z�S���W�Ճ ��)�@Lx�4��'^#}�	B<���6T�\��E	���X��IM�'�Xd�s�\�Y�����d�'�J7��O��~V���S?!��l�d�]�`�a����:���I��٨#��YI�'}"�'K<1�1�B�Y���1�H��B�(�,�8�k�/Ld�î��,�B�3�(OЀ����?#������"����ʳ̤���ȗ1LR�a�Fq�ft��l�'xf�h��?i���	��gL�ԆV�f�
u0�h	:�y��'�*U$�?���5B��h5J���n]�'>lH�Iљ5�ic��RR �;�'4�J��6�$�OVʧT�����?��%�b]���	�_��ѥB�( �f��B���?�y*��̉a��b�֦�"S�SA�;iPEx���'�����[��$�ᄤ©.y�=CO��K��h2���O���2l�%jRt+tK�
&���G"O-�V�T�g��Q���&z��јE�I��HO��O�ӇcՅ�lijeƟ���@�O��Z-�Ո���O��d�ON���ݺ��Ӽ�(�&\���wmL���4E����Å� G�ThC�_�wU���g�'���FW#8�Dh�G�v]^����[	E
	ZSD�_ˠp%#ہ���Ν jN�i�<���E�j���Ͱ`z*�s�Z{?�d�ǟT�۴*�f�D�J��Q�M��� ���xq�F��xr�'��x��&��gυ�VX�#�B�'��7��O�˓I�=`U�i�jȣ��&K��LGeFU��e"!�'r�'D�o�0���'��	L�e���{�� n�;!��Rxn%��d
�~!�D�'G�"$ވi� �8a#9�BX!���{�b���& J�U8���p�>��*K��2ٛ��$ΒyxB�|ӊT�qe:z'��h�u���ZE`�O(���O��D�O����Oē������T7�sb��GN����4E�ax�.�J ��4z2J���h�u��I��M����$S�t	��o��|�	o��/ؚbY��a���ҩ�!i~��V�'�'�����P&T���'�@9��X>}��iߌ4��hǀ2rX�4{��8ʓA�VỵLS�$�� i%+b+d�Rթ�s�<�z��9|��3�[zt\H;�F�p�'������v�n�x���|�u��~_\E	���G_A�c)�*�?���9O�THፖ%j'Ɛ�����(Y6��֗��E{�O��O0���{��w�/l\�`R.���yR��Y������'G�Z>٫F؟��	��������� �lЊ��f��-Q[\��c�_QL t�ŋE�?�O&1��Mũ(��]q�a� "*�u!aH���-�w��`�DT�~���O��5�C���Q��!2+�2�瀛[c<��O��S�ٟ �'r��TC4g�z���D	+� �
�'V�)t��,NM��q��{��x*���b���t�'�,�r4Hԓ7���2�J��|�d��$�'�"<~v��g�'�2�'rbj�~R��|�`�٣J�>0�h82Ǯ�$^s䵀4*i��M�4@\�p����֭ä������h� e�0bWN�:�P2��6B�
 Hݴp�`kS��<j��U�?�=���k�2$x���1QE��d��?��
C��?����?�gy��'o剙a<x[�G�8�h��d�S�Bd�C�	�&R��S�D��$�H�"f�0"�~=���Ľ|�-O
l��oӦqqV����#3h��X���	�@�՟�����*QLm�I<�'q�b<CC�A�L��"aXErܙ���mt��o��wb�Y`P��O�y���c*�H�F�H��n�:��&1d�b�ˇ�6 ^�hR�N65�4l:��H7������Ox�l'U�B��!K9���Λ31ƀ@M<����?i�ʟZY��>m?�3!���4��,�'�'�ў*B+$� �bh�HVXI��c��9޴�?	-OL�abc�q��'��$# z-p�"T�b���Ф�T-k ^�"�%�����	П�*4�K0402�A� !R�"��LڴYN�hk3�)J���I1������3��=�<��_2|�tx2��4�F
��	�#S�I��n!ve )	�F-�������' �<I2�P��	_�'6
M:0!ɕ|��I��	��P��?��h�D�sЍ�ypfI���g�B��񉝺ē[����+����vMJ=l�^l�B����X����b�����R�'���R%���,��h	�Ca&!b����$Q��"��9wA߾f��'ØϿ@D<'�(bĬ� T<\Jq�* g�
ህ�q��)�#���/�x{�����Zfx����i>���>[X��V�4*�j�xч�(r������O�IoZ����Ou�ɞw��4��/��#�q��/��B��?�����g}�J��*Zt"<�鉪����"E#
,��")�|�ja�>�?Q��b�2@K\.�?y���?I����O��� �I#�S/nwf5Y�˝2۸���Q-"�8��U�[����PiƬJ{��I+j7����P�r�h	��ؼG���uC�%_ &y�Ϝ�sqʗ
�?-�b�["B�V�Oм�E���6@01��K�wP�e�H?��H� ��4o���dG�+L�2``��ǽ$͎�!bL�xr�'�:�E�����Cw-܏88�a@G,ғE����'�1O��%j�x�@���`h�\hw����y���@\�fm��H��0����y�J�.+���/ρ=Bf�!�G5�y�`=��	S��5D��i����yҌ�6�QX�9B�5b�䒄�y�$��7z�k"�ޣz�i��&A�y�jM�)���р@Q�^"|��-"�y�i�N���/Б	:�m�q���y��2=�\ѳ��1	��h@���4�yrNK�zDH4y��dК��Ž�yBkLM,F����Ã���! 	N:�y��X�ZUޱ���+�p��I0�y"��^��i����i�`��d�C�y��ѯ"N�	���4��1C�A��yB�n�b,+"��?`V�#�/�yr*I�0��j�o�VL� C�M$�yB�blB(��  ��ؓ��ybㅰK:�|�c*@�'��hȵ��y�M�V� �c"��%ڸP�Q��yB��	B�$��rB�7-��Ek���D��s`T٪&��>N�X+Ҿ/�t��/.1��Y�CE^�H�k�(�x��ȓj�B�С�?e
���4���#5�х�JP����DTw��1���hݒq�ȓ�p�!ׄQ.zV:�+ʳ-�T��ȓp��� 4>% g̈�������)�UF,�"��j �"�~��ȓ\���P��B#2��\6+��4��w~T�E�V�B���=S	Lx�ȓ2Z}eJˉA�p���W<n�ȓFF$a1K�vs*mB��'��Q�ȓB;�M�d@��?����@�+�:X�ȓt0�Dco�t��U�T
�8��ȓ����L��,���| ���{�LD��&orT1��"�&zI�ȓ8CA��%/�#`̖V�"X�7L N��9S�jb��mk�'�u��~r�թ}�B��V��g�"�����yb@X^ꢘ�S��5Ol(��fQ9'��T�"�	|E~\�ʙ*v�q^w�Q��i��E�z`�])1/H�9̠����5lOf
1�	��z���`��B�����
f��p��Ȓs�z�$L� ���.o���@�m�[6E4�OLA�;<�1$�9�lMB4d)����"	^�㥪1nD�4!�yb��;��Ѧ �f��e��p6x����P,ʠ�i��J6Q/|� �􉴟|�L�SUB\�V�Q<��V�#D�x�@ǜ%&�lek��P�\�c%�7N4LXA�N�44~V�	��]�0�m�'C2�P�
�Y��
E�D�P= 	�#ah�kf��c�e�����RŮ*�k54��q��Hŵg|��)Q�ʀ�p?q�@��6�����	��cbR=ڐf]�O��Z������/*` f���E� ��rE ��;��3,C�I{��Hj���>m�A�Al�5�$ճ!������@��4XD6X�uH*ҧ�~r`���a���	eȹ�f@��y"����hڴ�҂9l�E[6%X��M�C��)����*E�� ��&�>Ir�Ϋm�p�׍��?x�{���D؞pPT���Tږ�έ7��q�.�f��A�A�=���,OX%��g��HO���ʽQ|$ V���9�F+4�HP��׋,�OTa��*�'"�eZ��+X-d�R&I�|R��a̘PcD#�E|�k�
��(�Q����!L�Qa@+���i��<�,5���c�
�h���*��jB���\tf����O~U^E�J���x�r�7��]��L�Fh��@�!�)@"�>��1Eߤ.Y
��	�!E"6�#�Ӽ��%1�$��f��4>�j���<Yܲm�z����'~����HO� ��9Ԁ_' ����$�6%�,���n�����=����Fp�4˶EXO�h��;Q,�a��O��8�4{��05�5Ŋ�('��+��(��G�e�������f"Wl��U����"�д���d!y�DZ�a&����KP�JC6��Q�Td�\>�b�$͑��M1��	o��i��4Y��yr�Ѻ-��qza�Sm�<}���Y�c�
��f��S^:�g:��!nS���sb�!D�Pr���]j&d:�g G���F,Ŧ�"K̆�~J?7-C�f��b�R"/Yhx�ÈѰB�b2 f�j<����y,i�&6�Ӽ���Jh8�ʰnHi���hG��.��n%[�-	�'�� ������r�� �c�K	�����」j�Z9���#om y�d�Έ�hO"�:d�ʂN���A�J9<س7��<K$ ����/c�n��'@�s�ͱ@
`��L<q'������-g�n��#H�<3�����Y�N�:�fO�
&�H㧀!��ɾ�m��^#������)���O��Bc��P�0m7���WΖ�:�����*wYF!#��N.9m|8�A�= oQ>��ܜ Љ��4Y:@�ĩ�<Yb`k���+D��J���Mz�!-�Xܝԁ��|��Og��a������Q�[��$���HV�p����-���e\�.��.�ў��Yc�����@�������FJ(_��$ÇD^(]�$�yp�-串��>Q��9Z��.��T����;`0(��#�:�三��C�M�A2���hO��ʃ�_}�r���`)ΐ� ���7z�C�;B�jY0��A��7�V�"��`xC�K�Ms��'2�����7H�Y�e��^�k@h8* ��*L��"&Gq���R�&&���Ǣ^XpUR%Eئ�a@D��^��T�٬y� \L\�x�Χ?$���ŋ����@��>x�}�Cʝm������k	�DS�a�y\�,�ק��UDX��H_u�f@�í�r��?�[��_W+�睢Qx��1����T����]�<|��A�(|�����TLl�����5+��=Q0�Ʀ��"�ҚKĄM�P7%�@P����R� (
1e�79�] "dj>yha��T��Yѧ��+�Dr ��r�"ܙ���+��Q�V�I�E��`��H�&(��B�6Ծ0y�ȝ,'��xq�J�H����`��'
�X�v��WǬE���M(9&Ȝ(/��8��K���O��E��Ph2I� �.Q*Y9�O�e��%P:ZݢU�vB��B?hub]f�q:D���I/ �$U�C�X|Y�KU�.���@�BC���"�Ň��(����W�
�ࣉ�R�����V�6�
x:��(E��Y+��Ҫ��
��y>�oZ��Z4�;d�� ����*ѺU$ΦE2X$0D�
+ �@H�E����mX �U"�hO���`��X�"I�z��Tz�m��g�H]o�\R)��P�NO��s��'Ab���-U�}�4�����O~�� ���TFX��W"Q1�ڹ"��X-p�ўp�D �1Vx�
ЄQ�2&��]�;S��
�8��`3�ʛp8l��ɍ`A�!�w�3N���0�����?��^>���H`Fp�vi[2a���C�A2?�$�$B��H��V�.��(�n�&}i�Pj�f� �q�a�
LI��&�N�r�����OTaH�M(�)ҧB���ǚ#��1箒)*��kP�U�`�;�"0�*ȓ��ξ��
��<��'���ͻu.n���ƛ.L���pB��,�$$���匔kx��rG�n8��#�
"��0�G���a ꇁm4"���'��#�m�a/Q�l��������VPZ�B!�	:
�bV�C�Aoay�J�34�25rA���V�����>:K��^+�Y�eNB#V��죷�i��O��������c�K=�Hj�"���e,�	�N���u�4
bC�Y�	jk�+�̗�w9�Dz�
��}r���ӻ�l�8�H�S.���KE�0�ظ@��ըL> ���'�
��	n.Fd���WL���'�\㞨�0Or��HPҊ�,Rn��F��L;��cc�$e-���&�F�*�`��L>�"�f���|�� YG��,�dj%IS���uF��5�(��EQ�4��i��� IY�*��m86GT!V1*C�H����J>)c��?w��Q-�0�D�� �
���c��6�:�iD�׶���s��L���ª��L�B�G�$S��+"ٱ�#ء(���zd(Z2ɛFa�>��C�$��,N�2��s+ɃhY��x������D�ɽ(a����g�fa��&�`SC���b�NN�Fh���@�ٝh��i�&��I(����US�hՉf�̺1^(��q������F�,^ލYg�S^?���+qO<�v'�Ũ��E�8�`���#.~�:��@��\�ʁ+{<&��ȅ�O�:a���U�����N/Z�+��44`�1a�Y�
�����	t2�4�0�Cp�Thd
���� +[�
[*�O���X�M�O� ਐ�
��?���Q�i�ʬ됂�b�r]�s���<Y�)# E6���d�<h0�ˊ$�����,DQF����hFq���J������H���6r�H�P�I���I�P"�Ma����pbt�1q�0YA�ޱ.�D�!'̀�.��O�"GF�!I�z�!"�kH��9�-'J�i���F(shQ��h�>@˾�x"$��ke|���f�A0�ڮc��h���O�hP�=�����C�L���-�' ԁ׍:���;0Ĕ	^^��rf@=8]�O �ϟ� 2b� #qӾ����2^ܨE�( cV13�-� �	��;5�� o2�c��\%}��Q��Nސ�O����i�O`@��\<���v�S0eU�a�r�#<O��r�C%վ`�v�&4(��{2
V�h�	��3t�Q2b�g#�#<�O4܅{Q�	�L��)�>��|��m�1�8	����8��S��	�/�L�2�A��/G:"������Ӑ�H�
W4D"����C��H��4ɮd,p�$�+.�8uKT�4�B�8�	'Cuְ`�+�n��)fN�,[
�	+V8r0���"f$�@�� �����,O��R�	��,������?w�f�ѕgX
e������]���q�Z>r@�vb��!�v�A5J���Y��+�-�ָ��>#x��Ǝe�4l�Ny�OPd�8$"<Y���r��Վо���'pd�HV�	�BA�
FY��� ��L�o�JeK���PȔ%{���q����D������Zw����*
�}��@W!�`��`��OR��"�R�}@̜Ö���~b\D���|�O]М��)W�X��$\�J�Q�O�ŸdH=�)�'0j4��i^!Y��e���n���VI�$�mQ�)����-L�����wR<�;�-��P�Qz�R�-Czu�N�D���M�:ۆ�D~"����`R!�ɪ+�pu� »#ɌZ*O����I[�Ho�%1V`�sT	`��>�O`����ϛ �|q3��,,/�I��X\�'����&�5s���vJ��h��۶��+(�c��q���AIJ��D�8Cn~�a���bi&?�'����Fc��E����.X6PqD@�?���#sܠM�f���;�����4��&j)����LF(�
�nI4A�"��#xu�j��Ҍpk�3>��'ˢ�I�pܧHT��+���w���p����G�F%���H�&� ;��<9�mU�Ԟ�)���7(��ywN<���١oɨ%�� a���Dϲː�!	���O���܈>[f�ť1�H�-�9*'ޭ�3e׫5�@|Z#�AN�dڎ����N�\���'"d|m��+�LD�c𥉔G[�"F�'�>"ɳDL�B׊i;0́
&l|m���e�4PA��Ѻ@�H��3�AyBYk�!�#߄.����ɠ����-?(8��>_Gf|���/?V886��Љ�{Y�$��
�<���ج��%K ��y�F�H7�)���2�RM ��A{y����ɫwB@D����-u�i2�h���|j�#}��p���W�[$0OB��꟞h0�`�r�b޹���͑-vHЖ%]�f�iQ$-?��%[�~M��8�7���P5I
�,Һu��R5"�5N��ɀ�d�2��>�%�'I�d3����I�3br,���3%?��Cf�N/'_4<!��Ē8m�v�] ���0vM�1b�*Ip�:vZ�"�'��Y�_��k��[� ��6o^��Y����@�>r��H)��[�C��r�1���ѳ,��Y�Z���ڥ
<�%ms�(��D�?}*��]F��z 
Ǯ^b���ϗ

�N��aL�<�N�_���#�vt��t�YF��Ȓ���n(T:��7���c "�i�Lp9�O���g?��� ~���Z�MN�s�
��eE0?�����gv:��:�r���������������kR��9]�I�(�?�
h#E$��f%��<���s�=�� �Ư0P�x���`	"'� �>a�.|
 q�ׯK��!���83���� 
�sL��� B��2Ġ�7�*��?����3̀�>9brʕ�"�z�s�E. ���[�)?	%�̫� ��3�N�0SLB��>-�5&R)oc�Т cD>A�:L�`�a���2J�F���>E��ۤ{ Y��B�! � �X#�P�S��L��	�5N�� �4V�D�p�)`�	UKH��N�4�� 3ʌh�H�4�8��n�9OPޢ>!�b�VU�)[6�S:Аġ�e�5�hQM��%#:4��?��λ&b�a��D�)��i�H<h�ƁhF(&�-��M��^?���n���gl�#���� �̸t�MD}�0;F�3f���[:���m]:hïإ�!�Ąq�2�
��3DZ�E1��ǳt�!�,9h�w%	1~�Z�����!�D�S��ez�N59զ��1�ͣX�!���p��$K��� h��1BM��q�!�䜐6���f�
4ID�X�L�!򄊳
�T��rA�?*V0E`��5�!�$G�j&�����Џm>�P�`=H�!�D���i@���)X4�ia�aK�hS!�D� 	����G1��J E:�!�$I�'ݲXY2�ҥ)Z�+�O[�:r!�:��z�m��|�H��)�!�4~F����n��:t �)�MO�`�!���ݒ��R?yg���&4�!�Dވς���o��i��l�12!򄏛~�a�X�d9||���0d'!�$�k���c��)H���$F!򤃸U�X|��Z�}k�	k��W;D!�D!d��h�V��)7>�maӈC~!��-_v4���%:0iC&�]�!�("�ސ��/O�	�U
����x�!�dZ� AEg^�DB���cI�!��2}iH�еgy�RH��.!�D̤�p��T��O�t����3�!��S?j r4؂e�1}"H$��N-�Py����TcJa05�*s��;��̈�y��[�i�E�hYmy��!o�'�y�_V>�$rt��*k.�Jw���y
� p	z����$�X�2��0�"O����+�:5�S2�߈v׀�5"Oi� >pӲQ[�J�!�J���"O��S��_��I��Ȃ�k�TțS"O��c�G>���07G@�<���"O����	πq�0�#� �	�803�"O6�0 �X��Q��A�U��ɂB"O&��q��!1�x�3��#]8b"OQ��d�< ����� @�1!"O~M�V+Z5T���ɷh�!V�N���"O��⪚�C��ɡGܐKƖٙ0"O���P�J+\0�P��'�Au"O�4�5&�ܖ٪%.�2c(�B"O���������X�|!�ek*D�2�Gս2�|�"�A �:��i.D���*](L��a�(�c��x*,D��{��P9L����Q?g���<D������26|�}�%k��(JTl�P9D��I�O��#T"X�@B�!!�v��1D� ���8z������|	2	P&K0D���7��o{hl�r�΅*�H1�Ҍ0D�䣐��'r��hq	�b�i�	-D���5�� ;��:���)+�|�zBK>D�p��GEO���A暨XA,��+<D��ç����I��d�m�Z��4D��q��^�-H��
t�W�Z]R�$4D���b�9d-r]��&��(*�r�(D�|��Nǂ%���;�b�O �]�DM1D�����7M���L�=�$4.D�\[ׁK8al�"��:R��1D$9D��f!ߟA7���@G�"!&�����5D��k�Q#
:|Z��(~����`0D�l22jQ�|Ĥ��i�?j����&0D��bT!˨F��Ik/�'n	Z�zpO.D�4R�OΏ7+,9aO�Y�BhyP�-D���&1��@;�c�l��p" (D�4;ņ� E{���`BI>b�h3+D�p(q*��/���g�ۂH%�<���'D�4��& �#
�y`�d��8Y�`�Ԭ D�@�ң�2g���R�)Y�t��J$(?D� ��a��� �F�\)�0�S"�1D��(Ҡ8"|ɪ�,���LMQq�0D������&z��v-0l�,em�t�<V
U�83�)�`*Q)3&xrT$A[�<A���&`�U0�ě�+�>ዷB�V�<T�z��s�Ǚ*��Cf�R�<Q�A�)�^�U�#0<4�$ǆP��}�d��D�1�X�@Q���J�i3D�@���q��}��NRDk��b�<aġʇL[n�w��xe��Z�^�<A� ;��ܺ2F	�B�h1�g�X�<9��Li�y܍_^6�h�^Q�<��� ed@�ത�3��x�MMN�<�!��s�5��bF(u��a$�\H�<��*��I:�=9�A���8�/�\�<ق���*m�-�%"кf�}���IA�<�M��W�a[P#Uy^�� m�A�<�� �6�����ϙ\�����A�<����0sw�a`��
X*�C u�<�`���(Z�I+Bˏ:9̺(B��x�<��b)I.�� 〝�qW�\S��LK�<a0'�e�İk���4�J��6d`�<��]N]����#��h� ��s�<1Ҡ��.�.����'2 ��	Yx�8Fx
� 9����1�r0�1H�wܲē�"O����f����J�mi~�I�"O&�cR�T�0B�H��@�����"O x�Ce��UZ��;�N�=D�R5�'�6c��ʗ
G�B��}h�!�!�NdX� D��b2��9yLv��W��/q�JD���?D�D����P�P�u"M(�(�5�<D�ؓf�P�5��C�֛=�Hv�'D��K@.ۆi=HU0��`��-
��&�d?�S�'�4<i!O��JQ�GŊ�*)L\��|'½pK��PTA��Έ$B:R�>�a�'���R�)D���m��9�'� � �Ƀ ��0ʲ��9�F���?D�<bbH*O����a�[��As�2D�<;1�O��fQ棌!j��ܲ�b0D��1)�#�z�1�	K/$T�e00�(D�h�CW$@JP
� ʛ
.0���%D��j���6d����Ş@ALC��#D� JH��}9ȀJB�Bi\��6�4D��� �@V�� �9[X����&D��{ �oCx<ia�\�e}����/D��@VI�<�Z�����e&f�Ic).D����A&��qJ���1 �@q#,D����ܦ��%iUO���-D�7D�P#B ��%[��� �ȍY0�3D���p��VV�@��g0sǤɀ��2D����a?"(�K1җ�j�B��5D�8y�A�2k�4LP�*�Y-�)���1D�pX1Gȅm���`2K�f#�Q�F�#D��b���vG�ͫQ���/dJ C�N#D�����5�8ɉ6�	8<`���
"D�0�r,P iRܙQI�S�]2��>D���T-Q�P�X(F?;��U8rn(D���H�W�ɐc,ÙP-l��*3D� ��&"y2u(ǣ@�&[�=D�̣�ã*�Υ�E�A�� ��m<D�(jҨ�&?�Ƥ�ZB0�<ʁ'?D��Sa��Qb>�p6��Tf��	=D��0`� �RDFܮBK�D��(�}��G��(�48�4��!�f�[�#΀_~LD8�"O �ǎ�:-����7���B�T�"O��:f$%-,d EᐔE��:B"ON���h�o���ƃ* N��"O�a(D�S�i�n}C�
�<�����"Of%C �L�dpY��.�,ߨ��S"Oh�J܍f�t�7�Q.{�`���"O�U[e�S�*�E��	��m``�ڠ"O��iC�=:��9Zu�ٖlQ�\��"O,�DJ��*���g�[�<�l�Pq"ON�熑�q3 P[Q�_�:�̑�1�v�����oĉmyl$�@�خ���D���y�H�_�T"�"̞	~�;�c��yB��PO$�f�1��)Peϸװ<����8l�P���MR3�,$GބI�!��4��3�B��� @(�!�$�ug��9v�Jm�`�a/�+}!�dD�f�zH9��PWv�f`�4�!�䚟I:D��6DF�dY��3%+j7!�؆?w��s��_3d�(�#ЛJ!򤎌�I�\��D̛c�O�&�!��cr��:Qh?B��F���V�!��b�ƽ�i|ɒ�yd䍧s�!�H/wvH��fɚ[b�!`�@<s�!�/*r���
�B {Be
�G!�� �JT�A�\2�(H�5g�)�`"O4��Lv퀴Bb�BN^f(�"O��Z�$��X����9L�T�"O��Ջ�nOr�pU��xZ4�R"OZu �o�@׮0��@�cu��i�']\��Q �bJ6�(�@߅/m�i��'���a7k�X hy[���.Ø]z�'"j�#��[�%"����׻-��yk�'����`��"��B��+ں�b�'�����Z�dxȁ��'����'�|�d�@J,���Q�Ȩ���u�<�%�*��e�a��y:TDj�$FX�<A�.D!=^��@A���Ppp��BJ�<$�ʊh�Bx!ࢊ>j�����[G�<!�k�{?� dj�!+|����[�<y���/��\æ�  
?L��E��K�<���ǂ-�xq����E�Q�Fl�<�AiI�q�� �I�D{�����i�<I�D#0EQw��҈�E��L�<��'��6:vy���^KR6:�"<����?�r�N�)Ug�pZaσb��d�6%>D��P��P8������' 8<O0#<Q!	��IC�DA�bX?v����kܓ��=��"	=~���+��ú9�|Ђ�{�<A��ìdO65J���7<� U �El�<���D䪨s�ج$��t�p��g�<��͹#�Z +ѥF ̠Y�T`�<4��:������ϡk���7�Y�<� aߏ`�:�p�^3�` D��i�<��!��|DH��c�(Uhf,�[�<9�o.Ar5�)�)!� ��IY�<��J����
#��i�*3�Nm�<y��G#�|��
$����S�l�<���ğuNܭ"�C�yv�^g�<y���g�x�ã��L���S�"�d�<��K��/Cؑ�����hV�Cf��v�<�"h?3� B�a��J]S �Ts�<q�BCXZ��5���E��\Å��k�<�P��Z~d�5g@���Sg�b�<�TB�/d���F�B
�\�v�C�<���҉Y�z�� HZ�V|��	�v�<���\/53��sp��@&!y�		s�<���ӥy4�	��5u邅��h�<A��T�{Tf���͖a̞�����L�<�P䈦h��	I V�,{B�s��O~�<G�
t���#�f'fy
Aq�<a�
@�-�$�(��_�bs���j�<�3�=B��!
���m��2�	f�<1`)��<� (�c�Պ���kb�<Ivl�#U�\��(MZ��=Y��H�<��#�;i�lP�M������D�<I�D��&�f��1'�	C".�X���|�<�ԏ��l�����=op���@�m�<ْ�۪=�B����^=`%p 1�R�<�T��,7�4k>B�1�i�K�<����\TS�D��U�N�K�<��N�J�KӉ��%�;9|B�I(%��4�v	T2T��=xύ1X^`B��.FՌ�ɴ-Рm�QQ�c�q�C��e2x��.�fK�P�gE7r��C�ɫ�:@H���!�Dt�͹\�|B�	�4�,00�T�~�bS$M�
�rB�ɂ@���b�V�;P|I��bB�I�:7ι0e'Y/�^�`0�C�)� l���(�5T %�B���w�DвV"Od�Ũ��p�*v B�7�عs "O8�c�+3[� 6o�%𨅐!"O�����Z�
�M��8�Tt�v"O��@W�k͐Ȉv��% �m��"O�X�r�ӕh�(AK���"�4�� "O2S��aa�!��A�0!Q`!�D
9�x��K�Cp�ؑM�:S�!��H���}���M
F͊ �f!�dC3g�aa�H>��4!#��m�!��nބ���Ɍ"/����oS!�Py�Ϟw�����*9�d��*٤�y�O�-�1��6z����꟰�ybH�tZ!x�(@>D*�x@�/�y�I����셑E^�TҌT�#��ȓ=4v%+P(H�*��'��c�4��W&H]��	��Z��t�����h��z��8��g��z��&l٣O�Մȓ<�:�{��3)�ر�PmW��Ʉ�Q�F]���6f\&D�f��b����ȓ4����0$6�PI�$��-*RŅ�[*�QɁ��m~��bDΏR��`��eqz��@�ŰrU� �u�%A�z���8v�|B���%	P8��!U:B��Z�܈�`�G.@��841݄ȓ'���E*Do:��q��;�`��ȓg�|��o� �B�J�mN6\晇����+L�qc�9��	ڼ%�Z	�ȓ%���pW圇n>|%J7��7�,�ȓx��}���}O�	t�Z
�V��ȓ�Z�aV�L�\�+�mDpo���ȓa�vhKE�N�+ �=㣈�>�-�ȓ|�Ȥ�v�Y*)��D�BȀ<��ȓ�l����Q.  �� 6̍��|̅�#H�h��D��n��搅�n��rt�D=;�09t`�D��ȓL��QǨR�3��fH�	��Ii��14B�Xj
�i��H��� �ȓ?��q��S�=3г�NE�%����ȓjX��s���/}�b��F#LH72��ȓL���h��� D��ũt,�,�v,�ȓ7���O�1<��P�2F��AN�]�ȓ{��1�EH׸��3�MK#4�l���:��%����:.��!���".�H��������00>��aǢy�r���K�zͩ�g.x��ݙ䣆F�Je��9F5+Q�^B1B�iV��"�@�ȓ2&r�c$�i��#O�FWD��:�`�!k^bxV�Q�J�P% $�ȓ�t([�H�Z�̑�E��B�x��ȓ�̠dE�V��L���B�tp ���F;
\a��,��I��16���ȓ��X��GFZĳQ�Y�by�"O6���ƍ�r��!롡X��x���"Ol��p���r@L�**��B�"O0iؓ�ݷ/Y@�!�`w"O���f��^�u�A�3�����"O�b櫛

HQy��B�h�sT"O���ì7�]	�@�a�L
�"O���c��fz�\s��X]�|���"O��Ӓ�Į��9��Ē!�����"O.�z*K�06!Y�/��� a"O\� �7�8*P�
�#���*�"O�-p���m�L-�M�E���*B"O� ���/�{H��8̈́�=sRQG"Ox�$8-N�#2i\� Z �"OLx�� ͣK46M��H<Q�A"O�t�Bb��@�܄��Ǡ_,�b"Ob}@SJ3u��<eC�HW栲�"O�!ЄԿ!����sdD>/c��"OR��Ј��$�l�+ӅN�3��i"O�=�k�$���K]K�R���"O�[bE�V��=pD Č,�8���"O0ѓ�*T�$����s�$m/"D�`"O`��@��+(�2=h��@>"��C"O��bO�&~��XJu߷�8 �v"Oj$I Aߚ}놵����+C�����"O��k���L!�t�����Lv�Yi4"OP�[�
ծK�6|�GE ^���"O~�tEF}��r��83����"O�	����D�=y�@�b..��c"O�Q鳌Y�+�H���Ұa.2uyW"Oҙ�cE�O%��A܆b��93�"O4�qm�=l�j��� ډ"��ĩ"O@1���L�vy��玎E�B��"O�풆n
+Z! �r�^�3�� ��"Oڙ[��Z�x��TW �4�ҡ"O���4�F�3��8/��cq&��q"Of�!��G�_�,p��I`P�w"O����X���F(QX��)7"O4I��Xye�Y��%׺0�e��"OR p�l�w h��
�`�"Ox�6�  Jݙ��U�]MR"Oܰ����5���ô�[�h�����"OP��&L
yV��ؕ�Δa�*="�"O
�1X�@HƝ�BȐ�p�$�a"O�l�!g!I�X�%�P�+q"O�U�`U�DArL�_�
lZ5"OzxF��e�D�Y�K�9��$1f"O�����r��h��
��tqX<�"O���6D։Z��@�WO��2X���"O�8vÙ,PO:��7MSZ��	"O`,c�L6H�x�(A*9�"OD$�3�Y�U�K5H�I1h9�"O�J�a �#���g�H(T���"O ���� A�saR�0u6��"OPQ�G-ʯ�u��P2L�����"O�,
QB@ $B��`�!�(|fD��"O�Y�=@J��R5��P�V��f"O��q��S�~c*���(C|��QV"OFh�2Y�<脴G!4�B"O�=�éB�=�1��&FP[�"O����N�4	J)j3f�E�7"O2٢�SO�8��a��j�E�"O�Sq�דB܁�J�/J�P��"OL�Ӌ�3Q}b�p	�>!���7"OTI���	?EݎQkç\�+Q84Y�"O���I*9���p��?V���0"O��B&�[�M�,���E���ey�"O�iR�G�k2N5��e�m�:h�"OF�h���'*��U�^�`��!2"O�5hE�ԐH�y�s�>j�^`:�"OB��3�%`��L��,șPx�}�"O��R��`!<����(<�v"Oh�s�Ɂ+!b
qkJ�D���g"OR0楛�nCx��%�D{l�Kg"O�-�U�KL�<JQd�	?Y��Z@"OpCʚ"{\d�Ӣ�1|kb��t"O� ���+M�[�E�ŻQX����"O�k&OW+u�>����?`��|"Oҍ�T �8�T� �I�>�t �"O�����C�a�,�	��0#U"O�s���t��aSeG�Qs�"OԽk�h�4Z��(2�°Z�i#�"O�+�_�$��"�:RYشA�"O$q����W�f��肄dR��3V"OT�p�H�v",U����: P�did"O� ʐ*+H��e�U@W�@��T"Obt鱣�K�< �n���0�"O���Ś�x�T4�׫�m�~�V"ON4��GU�x��1�(T�{�"O�}+�����gG?`����"Otܒ��	=4�t��F�
&Ӟ�W"O*���oˮY���"U'ޅU���qu"O�P%_+M \�flϤc,T�%"OxYVc�p�P�ɗ-4)Z��"OR�*$L&c��AX��Z1��h�"O6��b
2r[茐�K^V��L0F"O�]B7/Z�8�����`�"&�d���"Ob<��M*b�.mӓbS QeM��"O*�1�-�9=����Q�	S���!"O�^H�	xP)�I��`��D4{�!�D�Gf�=K���l��BE�F2!�d
j \�K�o\/���fC��:)!�D�*0P�ۅ�U.���@"� 7!�dn�VJ��Ө~��h���.C"!�$�p#��;��Ȩ[���B��6!򤌪6�h�2�߸.B0��s���l�!�w<� bqǍ�:tY� �Y�!�Ѩ
���X�G�pH*`X�`��e!�$ԉ5S4��mؿuG�(�B���S!�dGѪa��N�?Ͳ�)��7�!�K�|��I��@<^���aj		Ai!��ƆlZX\�ǀ��u* �ebʺkh!�d�G9l��7lY�	h� �=a!�$�3��R�F&]�,�" ި1Y!�dU?�L@�/�-8Yqc�J<-M!�$Ù�Tc�MY�GK~QYgm�d�!��Qʽ
��֏04��WN6x{!�$�p����wgז>/�IC��G,F�!��6<d<86f�����Ap���Py�/r���*�M�������y"��<[��㕧	 PI� ��&��y"�R�i���r#��~�rxBn���y�Z!J�F�	���InI ��y�a�)Y�Deyb)���d=�"_��y���!o)6��8MXx��a@�y��Ƿ7���J1N]y���n��y2,�?#���	�F
S%B�@#��y"LƎ����Å��J�Ya�*��y�ʊ�X�r���-G��� �b΂�yi^�����=#�����yr�'�FA)"�M6b�8����y���jGҹ�V�Q	Kr�3�y���`,�k����h��SeH��y"l�j7���N(C���c
�y�R$n丒&��l�ꥳ@�%�y"Fy���[r��$P�&��&��y� �頥;v�>J��%#r��y�hM7qD~�8G��z�"ݢ*"�y�Jəi������\����"o�:�y�ĆD�F<jC �fȅӗ��>�y
� j���m�ҝ3v�(F�$A"O��p�˰�t-P��Z��4W"O~E���5xG�y:DE+]� �K�"OR���B� 5����N�:��D9@"O<�k�b !".���@@Q�	�"O�XI@NB��������u��"OR#U��P��I�L�B�J��"Ov����G4+&E8Vi�$"�*�:�"O�9�%V�ؠ���A�a��!xs"OqH�$�M=>��E��fg���"O<�Yl��%�&�`{��S�"O0��#E�O�s /�-���� "OR��垁y�"�HĜ5zҸ#e"Oz��
�,tB�K��,R��E�!"O"	2���� V��x�"O�試 X�m	�Ma���3"O���+@r���T�X�J�e"OLQ:�M��@���cj�B�&9v"O�w�V?)���QǇ�3G�`�jP"O��豏<x���&���嘠"Oh���J �!��%(+FH[�"O$�u+U:
h��#L�/%��"O���g��+&I���"�!��B"Or	20�@4RA���>�E@�"O�(��z�l`����z�ऐS�<�dC94<�0OɮV^�@�3�I�<�C�>	hh�@'Y�!��]o�<�򀁕r~�I��A��2rl�T��k�<��i�����9&`�V����7IV^�< P8+WP�醅�"atH �I�Y�<���Z�>��y��ET:�`g��X�<9�O�~�����R�"����NS�<@B=��H�fV.w������[Q�<�!'&[1ӡ�ì��	S/�G�<�c�6s�$M0<TԱ1�CB�<��K�:M1"���
�D|z��G��f�<IĬ�>G�8B�E 
�xa�%��w�<�����#A��t������t�<��<�4`%�B�;�(�zgL�y�<Q���Q�]s�
�7`)��M�u�<Q�,-8�Q�Fƚ�X��%��O�l�<����g��r�$Ѿn-��i���k�<A�`Ƿ6��k�.�Y�;��d�<��ۥuRq{uj�a%�|zwoJ�<ق��V���b���T}��0�l�a�<aATҾ�Y���=��`�v�<�׏Y�M���Q	Cc�
`�*h�<�d =6c5����s����Df�<I���0`rHl��n��)Hj�<y�B�ERx�(���4��}�ëYA�<Y��_� R�Z)Rz��M	d�<!��=��0�`��ޕ�K\�<��O6x!����0����_�<y#gɶ�RL� ���]���^�<�JL�V�ِ����m)��u�ZV�<��� ���Q�?���uJ�O�<� iZ9I@���p蚳g��Y�O_f�<�&�7�$�I�	֮�6:��[e�<�w�'py���d�(p�.����Je�<!F��7e�P���<��,� -l�<�vB*]�<T@͗����aJ�A�<���\2U���Bd��h�0Ic`B�A�<1��B�^��!���:�$@Q@�<����I���	����A�e�^y�<� �T��퓳�Zq4M��&���"O���Bo�gRX�'���	UH�Q�"O�P1�D�k2b�8�n@}V�,I"O"� B��$5.i+C���j?iJ�"O�h�TO>@v��+���@���"�"O�q'l�pI�uP�%Ҧ9��	�"O�m��..H���C�#w1���1"OZ4k1�%7P�@ �"	�)+�pa�"O~��ť�S�F�i�cJ���
@"O���7�	vJ9���cSt]ɖ"O5�HЅU��yk�F�)4���G"OP����	�Ѹ%c�10ȡr1"O$���J(	�0�;s��J%0��"O�iH%�~����"��5	����"O.d��U+z	p��'�" JH"O&�s�ӌk���FcY�@H�EC�"O���K��(�p�h��E�AN�SA"O.�eh(�T+#lH�Unۡ"O4x�T�%ZC�p�"lZ1PB�X��"O�@p��/��;0,C6BE��"OV=�s`�Q�����5O�6�*G"O@`vhˡG�r]"W��.6�BL`2"O���tN�$L����'O�_6�5�@"O�y�B͇�T�j%�EE��ح:1"O���`WC� �ǜ&k�(A"O΅[��@������-2"�'"Od�3%���|C@DF�My��"Oh�c1$ B�%jH��"OF��2!�]bJ�9hE-3/��"OH�	6��%b!��&��t�$J"O^��E��H(V�R�PR���"O(E���#Y�P�ЅJ#	�)c�"O$ ���Sq92.ȟ`��0��"O4�������BMX0#!e��"O��cv!�x���ƫA�m���"Onܐ4�۪8�VLh�IR����"O� G,�QF|q�h�B���Kf"O>��+4:<�p��Y�P��`"O^�r�`Wcl���݀	2蝋`"O*xAO^^!���2!U�Zu����"O��Æ�ۃ��*Q8`dp���"Om#�ye�k�=ءq��OO�<9d^�p$h����Q�N"�L�K�<Y#`��M(� �����%CJ'!�<B��:UT�Y�/P+�Tx��Ƃ � B�2T,�Q��ME+m@L0C��37	.B�	�N/|
6f*�敘D�R�"B�	���08�g	>i.�m�Ї��,4�C�I?K�Z�Y���ol�u�%�]CݖC�I� C�HJuhT�*�X8��Fb�XC�	��6u� ㆥ�2c�)!~�"C��Ċ��]�x�p!ƈ�&�C䉓D�Z ��M��pc�%��+�B�	�Ǟ0��AJ	ԅ��M�O�B�I�x��ՅO�@�TYZAlЧk8C�I�?+*��qL�vZEH��rC�	2yR�(I�:M�����a�o��C�ɢC����l������"ڴ^
�C�ɰ�P#��V�]<�T{�ςW/(B�I�"�:��֊�5{��t��A!�bB�I�H�r}� �۳dp�Dۢj�7I�8B�%z�v�����{P����!,/jC��$$,I���ɪ�&� �VC�8=`���o����Ym�6C�)� xl����]0���$�oM�iS�"O���ģE$�"a�$�#&8:��"OPh�f(��IJ D��I(]�F"O.1,]̵��j*�&�"1�ש�y�L,6B�K7��R+(�2�'��yR�N%��%	�C����(�V(�!�y�g�� 5��-CAr%�jV1�y�웴��ȋ���%(����1g]��y"���H�b�
� �?TXਁA�K5�yB�������A#�!A��uyR�B��y��DW���3���>�>0���'�y�@�-�֬h�,͈>��m8�%��yF� �r|wIE�#�9R!Ŀ�y2�
�G����k�2K��!B	��y�A�A� �g�]�I�<݉���y"���*�� ��J�J�r��yB(�*�6��f�I�~���(��yB�mf�a��МD���`CH��y��Z��`�#	o���(�ϲ�y2��|�*dx6�ұSf8`2�
�y� C�x0�9B�ȎC���	"jU5�yb��B��LpMX�:.tP��N��y��ϏsRaj��G�t�����8�y�]�yg�,8B�D�L1�ᨳ�y���%|DLuɖ��|�ҡsIX�y�ʛ�$��
��o`ta��H�y��OH�� �D�sJ��Q��ٸ�y"n�_��R⠙��12M�8�yB���  M	�y��\!"�Ĥ�y�J1��:�C�0y��̠ ���y"fZ)"}�X�A��4lm�0a&P�y�\8>m� ޭg��D�7���y�ߙ]�~�O��va~�3,ġ�y�oޡ[�2�ŧ�3s�����^$�yR)�  npv�R�qs$���A3�y��	�k�6 8�kn>U�-I�y���4�Hq!��.��� /�yr��t�h��B�B�d# ���yr ���P �I��V�Z홧lA��y�QO3�P�&�P%��5̓�yŔA�P1� J�D��d�L!�y�%)v���p���=%^q���#�yb��u`v$!� ?�x�G.ަ�yR��|�n��I�=(\p�ν�y�eƲEZ�1T,Пz	V@���yrd� ������ܬD�<��0&Զ�yB��^ u�]�$3@�5���(	�'ߎ�ҥ<7�B-�e\�(��5J�'�&�i#h��M$f A�G�����'
��{&�߄Y �<I'MX.t����'Ȇ}y�*Yk(Ĵ(�K�("pv���'܀8�F9vĎ5A ��d`VI�'���gځ>��="�F�(S�<(��'��q���B��I���#Ҫ�#�'n�P�q��-,,�Ԃ�Æ/��a�
�' V�����u3��+��\�~�^4�'�~���[�@ɠ x�Ȃ*k���	�'�,-Cc)�S݊��
C�U��Щ�'����2  �]��RjT�U�2Uc�'F��@m4
]Ju!�� G��k�'r\t�cML�N���牉�qst��'�LI6�L�F��S.̒j�	�'�, �B�q��ܲ��'j�X1��'x�xu���P(,��	Q:c������ �Ԩr��7);���D��I���Z"O�p���ǥD�h� ���ph2"O��𑋌�+v�� ��S��1�"O�q)�@�(+GV�yGoF��1��"O�-;�z��t:U��  �Py�"O 9% ^'�	�ah�&�n�"T"O�q�@o��V��ї&�1w���P�"OTĘj�����3���"�"O�4	"kV�m{���1 �#<jz]�"O��q�>&H����ݟB0l�h"O��s��B��y*����k$�`�"O6<��#鞥S�/�%e��y�"Ot��g-���8<k�ME�4���iE"Oj�S�!����,Q��	�D��7�y��sΞ�T���b܌�$��yr�0fS@��b�g�*�(�f
�y��Z6*A�fd� X6��0DI��yrC��<��"*6Q�)��cU��yRcO�,�� q#H% � �p�ў�yBD�43�^��	�,�H����Y1�y��IN�Y1�܆2�Y������y B���°�	)^����&ʃ��y�Y�d=q�,U@p0s�(@��y�
G
'.2�{�/�4I�^*7/֊�y�`�1Hprs"�^JX�m��@�<� �!�����<O����e�e�<�Nߎq�����O4g���C�U�<1�퐕^�0��E_,<��r *PQ�<I���?��P�g&Y+S���Jb[P�<I��;\ Ւ"��)szt�2���W�<�̋�w��UI�D#-D�
�Z�<Q'ᘑH��%&�$u(�t�WT�<q�	�tW$�fe��2a&�"E�Q�<�&P2a�)�3��=~�j�L�<х��(VsN�i���O�6샡��A�<��#V(c&� i��S-.�C�+Gh�<ǃ.b��h/��Z쉳�+�N�<�A�:~<��e�%��Nv�<�恍�/w@�ȀDQ�ƸV�z�<!���6f�ı!%�2z�@z�m�x�<�����&�|$���E.]�	*C�^r�<����\�<����i�Z4vFo�<�ۈ(���+��n���D��l�<Ɂ�Yc���i@k��q��"S�<)`ɍ�ٰC�L?�f�P���R�<i�J�(tB�	�U��f��t�<�va�3�]�t��*Fp H�#�t�<Y��G:rQ��b��0�� P�h�n�<�Ҥ[	x1�r痒AO��k�N�m�<�!bA	k-D���W3BPs��<�d�*x6�kS�.l3��b�<�BB��b�P��6��lI�%�[�<14�P�C3��S�i�
[�>,��f^T�<��e��`���jڄCO��8�%�G�<auO�)F�f��%����`F��|�<�	���Q��L�bA�k��B�<I��ƏR���XA�*���Db~�<��@�XR8�#�f�v�̔
d!T�z��ڑl����5䟠(�h�F�&D���5�E/�� ���8&Z&M�`�7D�,J��*z�}���XJ�ˣc(D�dg�LIYȩR�#Q�17�&D�D�C�Q�{�ZmYS$�B�
N%D�
���2'�a�Z��l(�%)D�� ԽBa�P"J�fQ�V+þ�L9�"O�}���׃��<H5�%,$v��"O6��Y�P{>p'�!�a�"O$��wG/_y�(�CM��9oY@"Ot�aˋ�)�.�X�N�y���G"OZXktc�x�NC�,C�7��7"O�\�B �+h0ƍ9J�k���!"O�A8v�ĳ!sB�I�
)/�D"O��)K"r�Qo_;�.cQ"O
���]g��J#�ڠ|���"O���X�X� ��	���{�"O�)��`�v� ����
c�Hd�^Y�<A5���qi�	k��^�B\1� �W�<a���D���T�k&q���Q�<�F��"��L�5o�L�.y!!'Q�<Y�F�`��i���M�K7<����w�<A!i�
ek���Ǆ>="�
�E�I�<ѵ�ζ,6P��p�_<��iю�j�<�u!�=
��� 9al��Y�ƅh�<9t'�����*7p��}�֣�H�<9v�V��x�hb�2I�h))'��G�<�A! L|� F� �iS%	D�<����B��k���RH�A �~�<��I�p����DϝEmXH����e�<y�� 'U����aoHDҌ��΃e�<�ŌU9t:v���	�*<�e�@�L�<��KƎ23�L�{�-)��_D�<�R�'N�&E��Z�,A� l�<���ǐ}��LP���(>��h��I\�<�6�_@�h���O�
I�ã�_�<Qb&��*b���X�/��싴�KA�<1�.�DҢ�"�*�.K\}�kAt�<)��-m���UI֭\r��)�jp�<�"��4A���á̛������PW�<�AL�J0�庂�1�z �GCBV�<iQ�k(�bY-g�hP*@�SO�<)4�4 /���s%��n�\�{"h�`�<	ƌ�F�H�K���[4�̓��[�<y�F�&C �I�-�V	��X��Ba�<�D$ƻ;��l��FAK�6����Z�<��DM�X\x��6k��ڠ�Z�<	��R�-Bp�C�)$����`�<�� �KD��)G�1 �ڨi2Đ]�<y�͌�8{�abD�ծ�dq�T��X�<!��6[M�5h�C�'^�j�0 ��]�<)��O�d�p�����t�p}�M�X�<Q$��E����$[f�X$�S�<5M��|�6\i�ϯ`Ƹ`CM�U�<���T46xT
A�̬����A�[�<Ac���}n�%�Bj$��+Ԣn�<9e'ϑAPF`��A���D{PLR^�<y�/;/��T�� F2ق4�Y�<i%ѵjQ,ѳ��_��[���V�<A��%u���2,��ޕz�FV�<!��0Vy@- � O	^��7,�S�<���+mz�X���[�|�w,Cg�<�6��E*@��n�v�=�j�<yS�ѪoV8X4��R����B@�<�F�m�9b�hF�����0�Jx�<��y��ʅb�H���5�@�<i��zm��I�F�u4t��`y�<qe�1o�ڼ:s�H+����mXv�<IUɂP*Ҭ��օ5�J4'/�G�<!�ҙV����Aj��}�Po�<� �U1"�A)g���#IMC��Y�"O��3��ԫY�}��_4c�,��"O�	Zӯ]+�v���Fޮgbr�ۇ"O������)
XH��A�
9YT�'"O�0I�T#s�N#�CA7F��ܸ&"OA��ьa�y�#���@Xy�"O�4��mϳQ�`8�2eL�R���D"OT�5$޴:#`Dh$�� ���R�"O���5b��"�}N�?>~ Y:%"O�m &�H�v�b!�n�a�ͣ�"O|qvHL�|�٘��;ReL�K"O���&�b��7��� r4�ia"O�W�j`tb��2��4["Ol��G�X{��0�цP�QȂa�a"O�]3���<���k
@���J5"O�y;��\�O���Qj$ɨ�Q�"O0U�G��=aZ��<T�����"O�eJuEҽ]�28�g@7���;�"ON����C�1ݺH��߭ ���;"OTpB�E�N�pb�Cʦk�.H{0"O��pFM\�Ux�����W�;��E��"O�t���
y�@U�a�?�X���"O|,�ϓNX0"-'h��p�"OjlX-W72@���֩_&g=@��W"O��P��g����1c^�q62��"O��������뒰?�(��"O�Ai��'m�F<�S�߇&Y	�"O��� @S�EK	<Z����"O�RǛ`�� �,TϚe�t�J�<!�,�8�2�x�4)	�Q��C�<A�%;h���5(1FۦA���<�2�ή$��!CԄU��T�ٱI
D�<i�fCi����o7����vc�k�<��*� 0lh5)G-�.n�ʱ��F�`�<�c��_u�0���K�k08��Lu�<��N츤 a�I>Ȭ��F�<���T}�U���2�J�� ̚j�<a$-A�5z��n@�,�V�r�<���	�� S��HАRuJg�<����&�Di�S$'Q1���s�b�<	�g��g�zjb�R�J��ḱ�V\�<���u�VQ��X�jd�XU�b�<!c�B bRDY�SƄx��90�/@b�<!a%t���N����d�W�<Y!�gb�Uqv�˴D�,9p]B�B�I+3ݢsB@�/��R��V�|B�I�jG��{�R���X#'ɤ+xLB�I�>\���EV�WD��Y�EwRB�ɄW��$��0W�����_�T��C�I�g�B����=��.j��C�	z��9C�ĔlEY���!��C�	>3�����W~����k�t��C�nOi�eR�*�� �D�ń_�*C�ɀ��<B��:XF����#�(D�`C�ɱmr�0�$8�c���JC䉉na�e���WM2X���-ΓTk,C�	k� �0�nC�3�������R�0B��/���n{7B��B��ccZ�KQl��=e�!hT ^��fB�	� ��kJ�x�QgǛ j�lC�I�^�l��C]Ԗ�c`e�(TNC�RK�	�⃮(��ݨ�&����B�ɷ,	���Z�A�EhPH�T�C�ɮ?5���h̯;h�y���~�XC�)� �mɆL��a傭:�b3|]("O"����� ��k�K�%B��0s"O4!��%��V���g� Z.x�#�"OX��m�.T���a�Q�h|�0�"O��1T
  ��X�d֋pX�c"O����#c�l��%�d�q��"OH1�띬~`��"%�O@���R"O@�`��F�hqU��UΌ���"O�%L
�5"�`!�C�D�j��d"O����JU��0b�L���"O:R蝉"�(-0'�Om:2���'��CRŋ�ZY��j���7Q��'����gX��µ[�0,�'�dt󵇑ye �x�	$G%6���'؈S"Ό<�$����Lf���	�'�Nx�����@y4="(�:I�B��	�'`�3e�ґ����ɂ/����'Zȑ�i��R��Zx�I"�'���!�~mY��b�KJN��
�'���;���	bz�"�a z8�Ѱ
�'��g�I�=�l$���nE�k
�'�n�6�DԆ�f��jp"Ob�1q�� .�z���^&3��1˦"O-YV��;����r"8B"O�|1%��>�@�U*�t�x�"O��H���SbY[o�^�&<��"OH�D�[�wG�Y�����2LKS"O�qpǫ��T��a�D$X`"O����/x��ic�Щp�(Y��"O2���	V |�.�E�B,>l ��"OPxa"�G�`��S�%�#lĔ�;"O��A$��S��d���N�n���"O0p�d\�%�:I���BzF	�u"O�q��\UBf� ^��9�5"O���N s�~9kcAK� u���"Ol�u�0m�\�ԁ\�tw����"Ot�����<ф5+��Sh*q��"O�0pMʮ@.䐤��-���%"O���&�\�|�黡�gĸ	!�"O�i�JV=��y����w��-p "O���d_!}�`���
%��4�C"OHu
�I�<)n���)Xz���bG"O�ŐQ����i(@0`��@X�"O�$���J�֠���d� \C�"O@�P�Sv�إ�[�
�~���"O��!ƠLC��`@���6��3�"Oδ�&"7Q�8١C���8mH��"O�x��R�/D�Z$c�U��8h�"O``��#
o38qT�@i<&QR"Ox�P�А/���b
�A4�|�"O���؝E����Ǉ~"�]b"O8��$bӧS��d; F�7d-�S"O����
�8���Cg���KG"O�4-G4(��k�g�t�����"O�i���V�����eZT��)jr"O�����z�DݲA��_���I�"O@yq��SÊ�
��XA��E1�"ORq�󂃊T>���g�"]N�)��"O�1��F� v��E��W�CZ� (�"O���u%�3-�P�V�F<Z�Y�"O���ԎH�@UC�
:��h�"O�M�Aëfj�вb
"s�h�"O޸����Fc�� b�#O��y��"Olta��F�yq:-`�&>*��1t"O� T�{7Ə ~GJ O��H�:�3�"O������v�ڐ��G�=0��P9�"Oh0�i!}�"�R�Ɵ�(�r��V"Oj�c�mK;��1$��L��@�V"Oz���
b���̪d�P0�c"O�ѱ�MޝG�����bD.>��s"O��`��.t��y��<*H��"O�u�T��,yhJ��6jV(U�@M��"O�٠���{����f�Yo�,T�f"OԼ1��p8��;B
[-c]�)7"O���B�/;5�=P%
�)/N����"O�-�bNN5!��eɄ�0UR�'"Ofp��ӽ1�p`��r>����"O�] hE�#;�ђ���"+@�{�"O�@�!�ÍlH��g�:E��"O��K��Y�C��$�@ J#:�H��"OR�ڡO>a�E�Ō `��P��"O(xZA-6dQ� agIߕJ�\IB�"O�h@�휇a`�v�#��H;�"O��ht"��#!�s�O�8z����"O�#��Y�Bb�yth¿z�lLC�"OЬ��G> DN���(uz���"OH=i��G�j��%����=�\E�d"Oth�G��0�v��u�Ȕ9j��"O���!��8�ε%%ޙP��;�"O�T��#�6{p�+pCҰL@���@"Ot����#>]���&��/<0�s"O��IƫO�H>̑�,�8C#lŉ�"Oj�#b�*F��;k��)y�"O���F�ׄ"#��cۉ7�i��"O��(Ƃi�D��_/#���10"Ol��ڬ#��A��H1?�R�P�"Ov|�6�4����o��h�pB"OBL01FYl�@�୉�a����"O^��ؚ�4���M�ϔ�ö"OHy���7
Y@J2Y��� B"O���@@ؐQ:D4k�GõN�%��"O�� �g؁~~.��ǅ�?Y>)�"Ot ��/]&,�=��I%`���{�"O�`�G�%PUF���ǕUBJx
�"ON	`��]�-vHm��	��M`S� D���M+:BM�ׄV������$D�lsgD�x�!�'@<aنe@�`"D�,H�	D��9��X�bƲ��A*O�-j����V��	���"LT�#�"O"��D�'[��P -��>� �B"OȨʐ��1{ z;����Z/�	r"O�\:�cÂ��@@���M-(ذ"O�u���W�
X$g܁�ЬZ""OQz"���S�bU�g��A�@���"O���:����F�t�%��"O~�sN��G=���eポe!�Q"Ob(�&�^	�D�KrE	��@$"OuS��C&� ����֮e[�D"u"O�|G�D���a�E� I(��"Odi�a��0�����i��@/pT��"Oʐ9bAg,�BE�
�1 �TP3"Oѻ�ݳB�ⅲ�H�s4tR�"O�E���V(&i�}�g�1?�钕"O"<�q�
�6��xh�����`u"O�9jc �U[�hY��M*!ĝ; "ODY��n[�1�@�@R���k�B7"ONEa5%A)V��	�6c 6Ф}�"O\T�"��Q�R Da�y��"O� &	А�P�p�� '��0��V"OԀgkS�=�>��O_�_�ȘXE"O�,	���4����h��+�"O  �j�|1�DK)s*�X*�"O~Qِ�L*��9�Dʳ��535"O�y:ƁG&��@� a��Y�r�0�"O>%�!f�
P��8�P�s�p��"O� ��mXJH�TSS�R.s|�w"On=8d�t����+�8z��s"Ot$�2M 'm`ٱ�T���c�"O8�2�H �����������"O�`#%�̽<ͪ�i�ʄt���#"O
���Ch�r�a��8Q�e� "O�k@�³�*
D��5T�y4"O( �FH�<|-ă��6[��e"O
��3Y�9[���a�8Y\�Qe"O�ఴ�D�J�F>; ´�q"OB����d\qfg��?S6HY���
�y2B��:l�9p ��I��d9����y�J�)��-k�$�۲�͆�y��'Z�N���B�&v�,�8�����y�C5Cz�q�ˎ� ��d�.�yrcЧE=2��wi��v	�|Q�,@��y�l�g�P��FR39�a#����y�K�E��%I�5鐤zEAZ�yb�۾��I���	W�����T6�y���>cE�����0w/V���`G��y� Ҥk�N��p��v�"���H0�y­V64ֲ=RwϨn�T�zԬP��yiՓ;�"�:Ĉ�z�Ri�S����y�8_͐@ط��jO��a�E��y���U��̨�#8��0��C��y�$TJ�붎Ѹ����D.��yM�*o�<,
�-��{� |;�_��yB�،:�i D޳uW ��DI��y�BQ�L�𡃛o<
�xIK��yRL�0�d,�� R*<L��T��y2d�*��mIu��%1@x)�N��y�D�c)�� ��m^��B���yR�4U�%�$bf؄e��,���y" �-\rL���+Hp9r���yb%EAv�l���-EKJ��"���yrC�B*��¤K�ȡ3%B�y��
�	r���ӜE�,H��x������#q-TS���0� Gut�����H��eΘ9�V,�Aj�4�D@��e����򎁤@z.���:ق0�ȓ|fN5�R�к*���2�gE��ȓj��H{CN�*Ny
����؅ȓl�� N�P�1� �6�ȓF ���u(Ív��	CȔc �d�ȓ'�j�{��N*F�`�Y� �gt����ȖXс*�2#ۊ�b�BD?�؅ȓ)��n0t�9�����݅ȓM��)��`��
B��"�X���B�2 �)d�� \	]pD�4"Otm��"�9r��i�Q'�CMT�"O��h���	VxB�왟")���"O�4[7#����@nȦ;Ę@��"O�$IBK�R�NH�v�ƿ)��aP"O�]��Ծh��}����*oB�V"O����/�O���@��~�����"Of�Iu�Z�`��ѧNG�x�����"O�r&��n�8�OQ5�x�B"O� �T`'�pĶQ�C��*,,;�"O�$�)	�:Y�0�A�ņ'X���"Op�`�i	D���K4�N�7�v]i�"O�4� 
lj���3�"D��"Od��集.�d%)�J�4p��ۅ"OR �vu\�pᨇ?SY���"O��
�b6�n�a#�M�V��T��"Op�@��@���},%נ�sJ��y�f�R<;&ٿm��{�I��y�
'.�8 ��˰� ,�uN��y��t"�J���aZD�s%J��y��3mV�$�@�}	��K��y�(6�����-T��&���y�ɫtZ��K"��>(g�i6�U��y⨍6�H��O��h b�k�(��yb�Q$٠�)"-^6.֊�+F_��y��Nd��7&˿&���	�#��y�?I�a�2J��iP���y�ƛ$��iQSND�f,Ueވ�y��J�����'|�T�
<u��1��'!�@RWA�dlH�j��;j�8�c�'�N���N	\<Bm�-������'l
��Ӄ5�`L�EG˽z�}r�'9�-a%@��5��m��`�t�0��
�'Dt�w̑?;�n4�5A�h��=!�'�ldP᪁�'tJP�
�`r� P
�'L֡2*ې%����W�f���b	�'��P��=g��9���[�&��'�0��[�\���rh�����'�h�	�n�w�TSeL]8��-0�'��`�g�ٛWs�P�c��V���'�\�%n�!�8ջ"R��Сy�'�(�1u�#f�l<�-�:����'RtTQ�^�qh:�!�lĵ/�ʑ��'�P)�M����ҁ&�`�)
�'��Y��N�
=&8yc�O�!0 �8	�'�9��D�� Sށ���ۗRr�X�'� ��N9l&�˔"�:{��H��'I4�H�@U�x�R��^�['r���'3x����S,��TMJ�X�'GPxۥ��*q�٢ʜ.I�(���'g� �����2���'>v����'F����E@"?0����d�$i����'`���&H�j�r%�5��]� Y�'L�iqq�ui�!i�I�"̨�
�'�$<��Km4TpB�D&'��1�	�'���qQ(�#c���;u���L��=x	�'L�b���?vsNE�� R?�p��'�p�x�̚4f�x��"I���`(�'���q�,@�^  u��߷�(l��'�\\	�I
0�#w�ؕ���q�'8戹C��Ue*B1h�?.Dt9�'+�����%m� Ѣ�V/k�b�'��U��n�.�%B�,;!��{eC�h�<����]څ�e^[R�D[�"Nc�<����yĺXK�i޺0��K�͟i�<�T�[��=��L6�2-�X\�C�,	�I�)�-{����	���C䉜 �URr�iXb�BRCC��C��' Lt��*�n�>1dC��hʬC��<a�h�Q��E"��త-�"O�Tr&ΒDC�P�v��k�"Q��"O:  �G.����ݵR����"O&]㕪��uq��*R��P"O� ��X��ֵ
�	��J�/*�����$�O��b>�G�;� �!�C�ZD6�X�g:D���� V�H�a�#nΕMR�<�E9D����ӻ~R�P�5�ߡ̘3�7lO�'"���XK�S�f�<w��Aq�ؑ�PyB�$�Z��V������i�<QSM��a]b�a�KƇ(�����B{�<)êS~�8YAV!Xi3��hf(�w�<9DI�:\$L��B�LRd9�eYi�<9�$���	�����Ԃ�{�<�d(=4��p� �YIB����Hp�<��ț�J�D���X1�J)8���A�<!��5s�xQ9�oH8A��̣5 �}�<!�e˸bT�1c���3���Q��w�<I�aM5+�^I�2���k>ԳNK��hO?�	=
ݦP�@E�L��म��q��B�IusV�q!�X{��Ы��i�jb�,��)4�x��s����OA�R�PB�	����ԃ~�R\Hg�����z��=�'��'���U�D0ZU��m�9fd8����ډ�ȟ��B�)��4ޖ�'`�_еp �-��MG�,O�B�R�_/�1#�N�'7�,�b"OR�ò�	x̨����s�z)�1�i'�4��Ɇ|���tl��i]H��C7}_����>�`�$W7�#a/PX x�(�~�<�ClN!KHJhfEu�̓⪂}≙�HO��� q�E �=o��hZ�Q��x:�IQ�O���@g�I�|�Z�0e�Q r���"���?<OF��e�K^�8��+�#I6���W�h��)�'|SLDȈ�_�V`!G���)���.kFP�8�j� W��8�2L�>q����$�/w�aԠ�	���h`�H��p?�4�?�1 �Ac��ꐡ�: إ�p'Mc~�'���HU�N�2Ɩ(*���QwT%�'�����C�Ы��<4��<��'��=P�C�X����茮�y"�)��~4��+�+{D�h�G_l|A�ȓ��Ѵ��x������� ��ȓb7DP3��0r�ZpzP"M�X{�h���dy�M�)`$TmR�̩qH�B��<����O������M����L�?^���	A�@l!��Y ��	s��g�̱#��� a!�������&C R�:C�n��yr�� 	4Xb�`��,�X1Bi:;�\���f�:�@SiI8�>0@���&���ȓ���8�F�_�T`:S��z(p1�ȓ%�hQ�%X,3�62B�k�*�l�O(<I�U�]��gZ3LBN@��]�<!7d+�����ګ+��37��[�<si�;`���� �*23����GCZ�'��S#4	��Vj@?(l4-Qd/.R��B��F��U�M�B��:TN�}���D:�|l艳��;e�Q��&�8Nax��)m��D��
Rbk�"ǘvkX��$4�8������j�0�;ã�	yREy�|j2��[�����"I6�($��K�<y�OV�Цd@�j	�*ĨcI�<�5ߐl���,&q�]8UK�C�<y�&Y���%*H��})צ�~�<�3꒤u�P<`�EK'O-��T�p�<)�@�4#h̹��=�HI��G�k�<�Qc̲1{�I!C��! ��GB��,�' ��T�'E���ŀ�$���'���X�����B�兢�b��O��Ҧ!&��g~
� ���įĘ���P�)��G!�(a"Oz"!#О^L��&���5�r	��^��1$�)ʧ�̹sA!�f���ς'�q�ȓ+M�	"ñS��8P� uh\�'|�~R�On7䱩Q���r�q�nS�yҨ��c���'��'���%h� ��'[2���	�9�LФD��q�z�`���/tV�#=��y��i̩	��%��<Y/����ȹ
J�N�Q�a~��,��@�f	�
�zAx3�Y��y��@4�ᑂ�\��pps��,�y2� 3��,s��\�q��\th���y⭋�oZئEZu���|���1�T�E/þ�l�Յ��C�Ɉ&�8��'Ҩ��ҧ[�hј7�-���� b;2a��g�&o�����8�3{�D�Mܧ}�������,���ӡذI��	o�B,p��	*P��1�
�
������&Z�	�$2�)�'_x���(�5`��B��E�Y�ȓ�.1Ju)��l�N�HV*Vcz�Q&�@��ɬ0W<��P �>H��s��Z~0#?!��	�B�`y`˔psv}����1}��X��	t���S!�[.E@p����">��ɞ,O&8!�I�O1�i��g7)!�d'/�����4x��K���o��~����V�i��%h��|�b%�=9�>l���,�O���g]\����h��<�3-��'����{��t{�j������3m�,���*D�8��D�tm<��D�A�9q$5���+D�`(�I�:�.����WL\� ���>A�'e�IJ�3?�' �"����3Jv����b���Dx��'�Щ���סj��	���B�	Z\�Q	�'R��8�eӅ��(C$.gZL��'� \���&�G&9�dQ0FH-�M{H>i�'�q��iމ��E�6t8��(=��Y�b�8�O��'&pr!)Q@�1k��B�L8i�'��E)�%E��v�b2��p�b=q�yR��V��%}J|�# K; l�P'�����b�
�d�<�r�֡��كd�L�^����ڟP��4���G�rq�rf^�0��ȓ-�uڳ�ܜhǚU8�9Jr�G|��S�p�l����[l��m�2��-l��C�I��l��j]���@i�=^/�C�ɐ_J6���IT� {��$��*svc��d�|b[��:�	㦕�Kوi�T P'��@"O>ѐW韲tL��o���Ek�"O���	O�(��\�oX�,���r"O�9��;E�"�i �
�>�j�2�'=�O��� l��lh��j � �:��ht�'R�4�>�@��^Qx�JRzD��������xR�)}�Xz3�'�)� T7��?���>Yە��%3~�����-/�x�%�=D��AGDú5�6�;�'��
p���Щ<D�la�k�
pޑg	�=v`u�:D���e�84),�0�Q0]{����9D����jܻ/��rn9��$���8�D.�SܧLM���)��g:��bS�EFl�'�ў"|:���X[0P(N�;�Ԭ�gH�F�<i�(�9s*@���)�����FZC~��'�J�5�ڲ}M-�5ō�}+�Q	�'����&R�L9���)��n4`�9
�'�ܝp�Ѿ8�����fAT��'&�4���D'F9�R�H.Yg�@�'TH��p�O��zu�ǞNC�x��'b\2SR4)�Є��
�E8���
�'ӀKC�q�l��lG�<��m*	��� �U�u��`#����E	Ϙ��F"O�I����U��-���+% �jw"On��6�� D���	D̽��=²"O8X��NE������^g�*��"O��F¦>B& ���72� Yqc"O����mRd,� �E�i��E�"O�d�"z�:Y���#RX�Q"O���%(�#6��r$��7���y"O���ֺa�֨��b[-S���Ѐ"O4�0���[٘����]�l3�0�"ORyuOɟO!x�J��Q�)���"OP}�T����� h�!($XZ�"Ob�����9Z��q�G�z:`��5"O��s�Β	�0��Q�H�+M�yK�"O>ub7�B�j�.��lҴxE�D�a"OB��"�_J.�z�dK0���"O
�u✭�j�`u�˻5@bp��"O(��p��w#T�bCZ�#Tj���*O:pk�� *�Qadd+d���'�hSb���;9Z���㇢$�j�'��8��׎SPZH#���'H�h}2�'D�t�q�N�s��F:���'N^쉴�#-�"%vA
#u����'Lr :��Ƨ~��S�҃2Ht��'���$�:�0ԣ�/Jx��'���(��\�w����3N�	6�x��'�4��E=s�����.D��'5�	ƃ	7��2��@�Pv���
�'����+]�n��ALѴ4HB�9
�'!Ԭ��E8Y�&u�V�'��h��.ݑ\�t� F�!u��-��'^�$�$m
)fHA�0�g���i�'�m��&[7;�D���B�Z_� r�(EP�
n��-�GdӼH���cV�T�T�ȓL�~�p�%��J}>dS�8U��-�ȓV:�K ��6~�JIK5�W[����ȓ�j8�ݷ^���ӍX�:����?�>U��K�|B�8�# f�ҕ�ȓb�xT`^�-J��A�7�T�ȓzO�!Y�"�3q���ѦBf��ȇ�Q@<�s'th��rN�$�����es:9:ր�Q��ZTo�l��W�����H�`�
�qb��$�Іȓ�\�g<SH�&4�ި��D�8$B�L���"��ʉp�6��ȓT�5��(��]�2�!K�����QO ���.L�vݺ}Іh�?m��ȓK�
�%��9��h�'o�<}W8��ȓKs||AE'�oB��Aa��J!�)��?X})$
]�r������*��ȓN��m���XPP��HE�`��ȓml��05m/r�r�#��C�l ����m9� Ӥ�6sr�Ӂ�рD���|E."7
#+00|+���7x�y��e ���#Ԣrg%���h�jm�O�Z��_
e�T���'X�< �D��37G ZC��=�ti��`�~���4�F%��<�6 V��J���$I�����a0���cӠ��樑�I|-+Ri�`�y��H~)ϓb��f�7zA��M�9�<��dZ(6�h�G��+ޢ�k	��b��cՕ&[6b�m�Mn���O�d*��o��L	� �,Zj����K'@+������O��G�r���B���-�%ʒ����y��>��ˣ��z�aRI� �@��P��>,�щ0��$3��up���i���R�X%�yW��?��X��,���c�W6��?�v�3=*:@��a���x���d�b���������!#PXh�"!�{:��� �Г䙓F�(`�p�W P1���fJq� ��'[PX�̟�A2��G�/L�\B��&2����D~߬�RqĊ'�m*�Gf�U*�aظ&\�I�t�+6�'��%ɂN�.eHU�aF��2�$5����(�q�B��dH0��K,����3wJL��ѫ{�NC䉡u)"Uj�7u��C�I/q�p1"�GУS��Y�A�1���"�*�#p!��N̹���V�S��.\(u�����O�;�0�'#�aBD9S�l)`D�,̸�#B�Z�`��)b0H���� !��[fIء'M*i����)Ķ��?��2��l�3.Y�5���bf
�b�'Mʄ1$wƨ��U�ֲP���S��8X�8`�)�7	���郧Q��Z�!Eʀr�T\��IY_���$��fa2>|�'R��/�(�E��	���Ot��5�ݪ��x���D �V��)[�ޭ�Ǫ�GP�H�'`a��@BΦ$k-Q��_
/WD`��p2)ISH��=�Vt�"#}���4x���O4��A�\&-��(0�o��v��#X~�A�R�ɀ�j)@��2�������+ �5J����ak���c�5:9X����
���9�^���D��Wx"��"G8�Y�L�c����������1J�
"����� -��@+��N?���bhɬ>	���'�������BHn�i�Ɩ�9m���{��c3�X�P�Z��&��M<������ &E�@�#d�d�x��f�I�6l��$0�vMї�Ҍ1|\R�*.ACujc���!��~2h��"�,���<�v�ѣ"B?	ħ�R ��"���2N%�c E[��򤐷^�2�`0o�h�����
g�}��	�@ٮ��Q	�ɘ�8h�Ÿ&�قuA�J�i�<	{pGL6��0K`�I�]o����'v�t��O�� ��֟�pk�mչHv��H��xH��qtˊ5#�L���猑=�R���	E��O�У��4�vQ�Vě.���b$Fm�y�0#�*Zu�J˫ D���&;@�0a�ԅ/��3�ċ*/N 5�'���BV1��_\�}��d�|�� ���4�6���LF���KFC3/Þ^^�u����y��������T��a��I�/S�(�J�
_2��q�k����'�~e�D'�Y��!0&�Գ�j�i�N�A_�Y٤T+8I41:m�b��jE�IJ���$�#r�l�q&,�#EW�e�d���=C>):'�îK2�T9?�~�iW!øL���s�8�ɦXHԑ`�,����呥����7͉�#�[@�">�؄�I�p�lC����V�n�BANb��ZWH��g��H*헾"07�S��&L��O�����<-P�q����9T豹��B;9A����Tqg����e��)h(��c��	>(X�i�&:S�ėsx�C��+8u��NB�?��Y6"��%� qp�P%]�"�nڹ*�J�$V#$v4���':n��q�ؙiW �{r�E�5x�C�)֖���;!ծQ�	�"3z�����ڦ!ZW�۷$�.B��L����� ��iG4 L4�P�.N)s }ذb�5u�IGz�Z%Z�G�<�, ;�Dƨv�>�ʧOZ�{���pa_�tJb��{��A����!ׄ��w�>�ڗ/&|�����Ol��Qmϴ/]�T��$�rƍ�c�?���P}�ÛoR�d�%	�=5��K5��7<�ɱ+�o�L��P�)a$H�c��8�ʬ�������b�B>B@������ J(b!@�s�Q?�󕉌�{�I*��7Mȁo_�^�����_�dgp�30���ཫ5��=x�eJf�G�>Y��ϟ9]�̜�C��0H����+�*1�Ȼ�≻9����O�Y���'G̓��^�D���eH$Gβ50'��6P�$��d�-�h*4�� txY�qeO8L�L�ҁȤFͰ1G�V�]��dO�/�Hj���(up�s`/��^=��e�	<�@h�"���4��-Oj��a����� ���\��۷�ͬ&�6d+#�8BH:�P��ӹ{���"��µ4n8��B�C5&���M�.#�*Hk�&C;CD(�0�O�љ ៚`����d���B�e�_���9�	L� �8���m>��р�d�����
G�Q��ޜ�ls�C�e*���͛�o�Y@b4!5 �Ƃ	�Q۸�ψ�&��'�q��#�A X�v|j]2I���;�(�c_��$p�����N=7��$s&�¦ѐ$n��d�2��W�q�I����l�iBH�0HRTd:U�q�qO0�:`�i�$+/>�r�K:pp��g偃`� #&%O�m�Ha�+}^P� 1d_��(��ex��G���a�0v�i�p��馵�r�	�|��"������-{P�)��K �Hq��D�.2ܩ��tS�$���-c�.U#�$�Kf��!��C�;��b��S7@�}�䦋6�*l����/g����'6^Ҽ�g!K�M���m��ys�bG�� 8�g`T�xyv|���޴'`<���B�McO�ި�vD��]H�/ �"��̨pKI�uf�*L�I���JgY���(9W��/��ֺ
�(����8�
�<�֯��O$�Y�KN�l2��vb��?�T������ ӈm)�ȆO��K4�q���h,���n��D�fED��P��#�Z�%,�褮��jSH���ž<A�aE|r�����{���8,t���'K%�,��ЈZntX���X{����ý7��(`��$z��g�'�"�S#j�W|�{|"�s���k�0�3�@9/�@�Fx�_	_��l�'�ޟ=ޜu�eןD욷'S�'�ԸQT�=!a�v�C�h�(��A��P)�c�P%j�Z�8�"����?$A�։�F�z����2:,B�ԎZ��T�ʢ�A �C��w�Z���߉B��$�Ӻ#���9V1|�'"ѯ.� 
t���vE�$��J��š\�[B(Y���N�!�$a�O��E���P�ba�T�K����"��=��i�-�!l���H7�ߟ�KP.݅V���O�
sn���bW� ��i��#h�xg�ڟ.�r�Y@F�(c��Q����p�0�HV� on�ZƎ�X�,�E{�4��Ň�;��C�I���e ��Lw޹�#�<G��h
�އ��\���\)E3��[�h	'��QxP�vąJ�'I��;ԥ� �T+p����Y��=#�����H
�G�-�f��~J�ĝ?@sl���@*p��5�B��Vt:�������"w��*x i)ŧ�sr�ñ�'��=�GSTq0����g��d��%@j|q�._�4�W�B����IQ�YѼ��W�ǲLqZwW�P"��6j��-��,q�,�]:C��3���r�t�jgEZG�k��Z29JT�3��'W�@T@�:3@��#T>c���A��?c_��P�I3<�8$��Jɟ�+��ʊ��!�㭃Ѧ���ܝ~ǰPi!B�4ar�UR�U=��)����h � �*Ȏ��J�<f����6ԉ��8ړc:�ыRd���x��4H��)p���:Jm� �«� ��X�o߃>ƨ�����*��$HQkO�H��9@�Í�Lb��"�K�?	����F_
U��&ڨ=J���`EE|�'TR�;犑�BWI��FZh?���޹P��� � ���Ђ�(�B��dnh�Nx����S�#���H��Y���G�i;zu�Sd2����T�\"��QNN+Fe����fh��&+����т��Bϲ<��N���0wG���<"v%�s9�|��T�wz@��BK�30���Y��0"��@Bb�)�L(;S�'J>e sBH�&!L��2��2���A��ӆ��	�]&��`I=5*n�@�=4c@��L�)�#Yf'��q��\��v�	0�i't0�`���7gL��%��G��r�Η�����EvDh��"�!v`�Rǋ��u7F�q4�D6+�O��6��A��z�F\��Tŉ(&���R�!��|0�!DHN��bb�)�x�J���CH̸!�Ⱥ��K��M�'�C:a���9�*�F�zBь4�0��*�v�U	cJ1}"C�1�)�6��LqX��7I3�01�0n�Dq�D'@4^R#�u�v$���u�L�@R4N?�y���k�VQ�� խUK\�s�B�~Vt��Dg�'T�r��T:"Z:���喃F�Y�7@�/":�A�BK��v�9wo�^.��Abc�A#��l.6���%��8NbpYR��n�*�߉�H�.���K�$ȉ"$!�@�+����'CHIP	��BJ�H���{@�hb�œ�]j ��WJ�@�G��ur �s3�FP}�+�$�!{fU	�Q;3�|4AE��G�8�����O�����$�R�Y�gQz`\�:�jN��	��&vYෆT.2��ĠaO��!�F�B'Ѕ}l@�*��i2�Q�bA&��,H�¨∖�,޼Q�ZܴTPcju��-"���(�x
���L�|Pi��A�x�2�
%A�>�𔪇v��%*�AI�)�`J4�J�h`��I3sS�8 ��))`�郯˭�0<���#�Pd�K�yW~az�Y��ݩ&�NҼ�tl֕%+��A�j�l�����2�ĂS;R	���)	خ.@L�5Y�h�nW��fxh!�8�@e�O������%zԱ�
�H��:��
g6K�G�*Hb��I�O�=�j|�T)N�~ ��(F@�,��C	�H��л�`Ѝ$�r�)t�2�	�A;��G��#��uU#>���;��y�2Ab�-ܕTm�$�c��?a��5�w뒤'��U9%��;���c�(�~�,EnZ8*�&�A�LY{IjbТ��=�Eh��Vʖc�@x�R�TϜQ���V`�'W0�Y�̯O�XX�F�D̔д`�?�4�j�V��0��J*��'q-*��GdO|j��o��"nJ�7]<!;��:M�(���A-`�(B�S�!����S�Ĩ�M͂�:֎#Hr�yF��*1{J�V¡j��,*F.)tpֈZ#�=h�F�T�E��eSU��Ta���wM�@�F�a��]�T���I�~���6�	- �KA.��	6 J��  H��X�>B��߉>�@t+��̎�$��'}���3�Ac� ���k܏?��s��*Fx �A�kш����#I93Y��"�� �e���"sb��[ը9�`i���2���ac��O�0u��'��)8�^�5Qv0�$KR#�l�;s����挖@,yЂ��9�.�z�,]��Uj���B�(�Bʮb�J��\�GY�I�)���b1+�4w�EA���w���.[�F�Jf��*D`V�ˣ�I�u��| F�E.bk��rtF�:;���JW�L��?Y���@oH���))p��d8��D,fTF4��Q8:������nT��`�]�Wޅ%��X{���՟��W�E��p"/��A��C�Gle�2ŏ$#��a0F�c��ɑ/*]�D2r�[m��yv����H�B��1qd-�3���`lO�xi �$�%V�ι�RO"�z�+5�*h�F��\++�B M��P��6��H�P�3�%�E��hWJVS�j������}��؉v#ȫZ%��7"Ҳ2�b���h	l=������|/8C#j~����'�����LL*[a�R	�z~A���\�h8��/�������t��-;���%@Ker���k�9e���C��}^X�TFǌ'MV��G탗SO�Q�A�@�w�X�y�4t)-O�E[ AI��a�@�U�h�t�Ӄ
G���� A�_��"��T�c�*��֏
x��I��b�@=J�Fɣon�Б�A7_��J�!g�<Za�׍D��↓M � ����v@(���=,h,�@A�V'B���Gs|ZwL08�CU�P}H(��A��\��1�Ҹ0���2&C�/c�(�P��*T�c��)c4��"(�>x$���E�5���Z��K-f�&�p��3+Z��ɇ��ՙ��WQ�������%j\nt���tqy�+�LrL�e������ O֔P������G%mQdh0�+�7Ip C�B�#�&�S���|��`�d��!2*pKC�&P��w	��H|�qN�c��S�i�<�ЁjŐMn�4��f�*9�dhݚ�L�fH�Dz =6HM�ر�q*E�Nl�44� `�,%�d��Cq��o�< ��mϢH�m�����p��&l�i��ʓ~/����JZ�ϲ]�ӈ�����oT�RЖM�o�{̱8�'ޡ1����FY��!AP���@z�5B��1�|X�Oy���H�?DmX�q&�ڌ��'�K����*Wc�a$�y�႐p���K�*t8�UP6"Y�?��/G&���ݏ`��X��G@�ղ�D0F�k��̲=��!�����)�3F 
u!��Iv��4n ��f�8h�8�b�g8[w�(�y n�:��dT/��	�� ?%�0AT��OB��"˟�%��s�i��x*�!�)1Rt�#B��?DwT0y�
�?]�1L%\�.ݹ�nV�m���B�*ۧ�b|�%��~�t囶�_-B��Y�a����d4g�z9B�m��f>8��'�E�48$i�t��D �N ��M�hC�0��u�Q��X0���?qy0Ȓ�]��᠈܀ ��L��Bo=B�¬��\hJ��A*��N#6���Y��O���,J) ���E�*�\M�O�>��p/ɻ2ؼ��)S1~��h�� ٪����!+;�4�g���j����3���C�R�{��X�q���#�E�q���	^j@�!�,���D�����K��,��'��!�:���S�Ff�:��a�iD`,h:Q�ݏa�8��LZv<	y'���t�X)B�i����ŧ�q/�q3���f�,(�V��M���C.Λ֮Îf̠q�B�	�6Ҍq�/�~"��)H���1&�2�~�z���2b�(Y�R��	f�(����$X� ����w�י8b�%c��"k�� 2O�8~on��[^@����1�\�7\������]H��;4X��䚄�h�i�,R+H��c��ոXB�Q8p͗�p�6���Lݱ�?�'�`�QG�)M��1[���:U��t�D��9����n�/J*�X	K3�������6�R�(�l֝iq�F�x���H����0&�+��Y7��uJ���+f�A�bJY�q�^�(KȘ���&_�-��qK�=�6���C
N���V�4�3P�'�jQ)��!~Yd%�O����֩�2Y
J%��K�p��Yz��Rct`�^
b�Z.�(j�R|�D���h�.s���09:}��D�nū�D�)-���)�\ĦO&��+.2��X��EyB�
�Li��~r��[92l�4>�މ��,$-��уÀ�J.����Mݩ���bښX�'�
��ť�F�n�PjM,N�V}b�Q�Y9��rC 3<�i�a����0�"9HcC�(�l�(ŦO�s����+WS���&iSo�*��'1���LM e�l��ނrT�2#?}�IV�� Pp�Ǽy���A3��L�d�C`�J  \�� ���� /u���eg���Vp+�
Op�A��R�TLj@�/M�p�C����pe
���4��'�\q�a�QҘ��d`
HY��Vt�da#�C�!�dK g��Pd�g�����mZ�M��j��� My0��[n�az�#�*#선��CI��aȀ�p=��P3tY R��iR��"aV-F����@H�4��"�+D��B�"	70�|�I��]�qN�@`�f&��>���Ѫ��&��HG�n+w0ZD��k�~|뵪͒�y�O�?*�IJ��U�i��HB�^ D�����NX�u�Z�'��>�I"/<��1o�/
�)�B�F.lJB�ɱi��1�@ �=h�*��>����  ��P�'�r3ԭA�{��UI���־�y��50�zA��=�"�x��ȩ�yB%ʶBW�mc!`.3@���kA��yB�J.>�B�r`��7�B؁�$ڋ�yF���Ȫ�(S�<�X���,R��y"�\�_����I�7"��w���yB�aE���Ǉ�2�> �&^��y�F\6HR��eb6vƔ��,R9�yRnDi�8��C>(1�����yR��jPA h�3(hJ�H���y�#S�Iz�	k�N�Uv�i�i��yr�߬+����H���dYw.S��y�����X��6K�-�zW���yB��~�h��k�:� Y�d��y҂û#�8TsF�� 6�!�eG^��y���&'��M��B�*r�E�e͍��yB�B�{2\�QM��-�1h�HH�y�+W%"U���R�ĥ/"^Q��oY(�y�ʃ
G_"UNZy۰�M�y���(���PB $0��٪�y��ߐ7ɨ�NP��4�K
��y�*�9�	i�d�+3�j �i�>�ybgMw��=I�!R�!9v���I��y���$Tr>�j�&��!�>]s����y�.��P(�8�rꋿ"M��CR����yb�I�&��|Qta%I�L�ys,��yb� S�:���W7tax}�S��8�y���\>�8�ɜb�	�agҟ�yr��=���ՄY�\>��#�H.�y��G,��P�b�ӕ^y�4B�M���y�/2n�`E*`�&ِDS�ܦ�y¥Y�8�R	X�	ג�����y���+l�#�(�� ���yr��:X��K�O�RΥ�
S�y���~���g�1}t"䍂��y��еO�+�&�X�%�(���yҩV*/���E�ޮ]�9)EFn�<	GH)���"�Z"β��7��F�<��%^��<9�U����SG B�<���ߏJY�0%�_x̘�z�i_P�<1Gg�99,��)Sg=toJ�R/F�<����#m�V��1�baZC��D�<r ���Q��9\�qrLTF�<�6͞
�^�s�f�0�A���Qu�<��J�:y@ ��,�3!�<�`��[�<qt��d3��N.|�բ$�L�<�eK�.�؅� �C�#���*�*�L�<m�d���oI�v�~͐�a��<����iC�?a�t�S7z@a�u��r�S�ԵH9RB��-~q�A�@�&4� ��g��7l��'����~�M�b$��8P���{r�/raY�d�N����sj[���<Q�$��O���	�_Tx�QF$�Jm���p�Zy����M�j@iB��ns~m��Ɋ 0� S �>S�С�Q�<J�'��['È�y���XaBĦe�*ѻw6�`����� ���Ra޶>���-8KCP"O��S�I���j�{G�\�<A�!s�Ú�D�6aq�iֺs,�]���_�A?���?������f�p�!n Ib�ח?u��e�Ǔ6�0��$��o*�8�C̤_��Yy���	�x��S%	e1�Hn�*�:l!"�-1t��rG�J�й��҈��b�p�p0'G���da ��O�9�"� 4�<��NRd� j��5�@DGW,j�^l�0���%���� �E~f咦��F���8���HN�!!(�. ����>�P�N�Bd�P�-ɒO�p����&���HD�V�ې���矂|Xs��{C<����KɆ�"f"O�$�X �숱�EH�N���� %y��(���mW��ɤjб*�88��?]�rdO�S��e��w�\yp֏�r��ЫA-Z�M�ZY��
���@,�2�l`Ks	 ��IW���g>�өF52�.z��@qx��"�AB4�zH�"�	�zLP���C�
��-H�`L25�V"?q� � za���0d��YՂ?# �s���!l�݋'}:qj�b2"p&�Xb� �R�xG$|9�K�	\vay KEO�Z}�%�Q����Y)�d�t�Z�?�����.���b
�H����Cȏ�z�B��Ʋx������8$�N)� �½:�d��%�tjY8���I��[��2s�1WA�Uc���A�J�vD��3�`8;���7��H"Ʌ�fG��"C��0UB��'L&Fcr�V�t>���[�T��,���h��i�-&���Ai�<����'{����N~�'_Bl���;�����<}���!�:/=��K;xK���� ������Ѹ�����Ğ��~��]��Ν��%�5'�6:fg�e�
��E���AK����aur�=��IP19����'*(PpŎ����P:c�tKF��^���a@ 0��S�藱fW����a��WH]1E���"�.}E���Ag� S#��,&gH�Y@�1�$˓c���	e��(e�2��d�>��*�	�Sc�zf��~�s�Z8����@&4��-˳��U�@��"5Oh-؄F5bt�x����(B�$�Ia�ys�'Mf�j�P�Є1ŪY"?���z�-��X���35�͙Q��-�ë�)D�*�$>1S�V��a���2w����b�
5��@u�V�Q~|̩�n��) ����URf%RE�������9@>X�rC��$|�� �E�%���鴮I5-4� r��	(N�hRL�M�x��cˀ%fā��č'�����	�.<��˗�0��i����Pm����a8z��-�@���⟘�S|��x��B�s�5��Pkd�S�.C�#��X� �%���`u��=B� ����!
�Q���O�Rmv�#t�B�%��p)� \��Q	��%G@|�cሒ!��<��b���ا%IE&S62�Pȉ,v$A"D�\@J�㒊rO��u'	e��)�nN�P� 7��Rr�L��f[ ��؈��	v+��1�i4�x���<��jaޟ� ����=i��S�L�ٖ��u㌲>$�\�3f?a�̴��I�_7����?l��k޴7;��a+��dy\,���"a*�H�d��2G�$T��0]j�	"�rӔ��0�ɕa���pf�|�>�Bo�iB�aZ��M�F�ٖ ^(���ۥ"�� YA��j�I��o�j�޴Qf��`�m	7�0֝5��L"�%��h���A��+�V��J��$Q�Ɇ�
��HOBՈ0+A~�P�1�A�jyi�C�Q�F�JQ:y*��V�q1ҩհ���b�3E�`aAǃ/Q�@-��P�~%�=���r��`�!^T$� �A�B4��?�qF� �pII�`�G��`VC��|q"�V�&���U�?~ I" ��X��X+ ��X_�1��g$^���uK�7�Չ��<x.U`%΍Y���'^�D���"��f�Z?���ץ�MZ��⎃ks�|�e<yU�`�t�A�z.�$��片X:��ۧe�p�,���K�4,��spOk���K�/B\� �	z>,D��l^x��O.L����zbT{eg�cV��%��:2NPa�k�7R}=I��_�^ᦩ#�`��HkUQcQ�5ѕ.��4ZpY���5Vu�E�Ȕ��J�'Æ�W�Ca4��k�j�8I�bp)O���*3���0c��Q���<r�HIrA��?Z��a�،X�$X���E$)^��Ce�@͚��C7?�FhB8:T��!���Y�6|��OhP	�ȅ+�nUga �@�ÀF�Q�T�R���r�b�*D�>	fpAU���`A0a���Z8�c�ǔT�@A�d�ԃ	̖ #�&s
j'DՖImXؠ��2l&-�� �w@V�'q�\akW���aI��J0�R)?{��Õ6wq�BVD]�L4���gP
X9DM;ǧ@ꦭ�� H�Rq�<�Kfޝ.]i�	�HóQJ��Dޣ49J�:�{2�њ��O$^xBϐ��F=
�S
i+�����Թ ����#ғ`� ����y�V����Y
m3"9�LSh*��؇i8�����c�07M�mQ`��_�+�q8��f���+�l��NѴ<��F��5P��`J�<Ƞ����
���� ���-7�b%�p�E�S���Ѭ�#!�2����F�qU�����8�'��l��L+fh�l�"K 2$���S�-�0%j7�I
GR�$�T�C0|�$�BHR u���l��D�hhv��% Q
IT����,	ԩP`.<�P@�78z���g�/�t@�à
@x�'JpX!C�5Y �	%/���#EC�;h��h�����Y�	!?V<�æ��59��;��^�-��9��E�8n��(c�?��Q����Lܒ4af$E^]��SuOK
 ����͉�e@X����;�r��u	��X����"I�5���q��8?ɰY��d:/���i3kO�ⴳSL�zGڜ�R�4���+��9ưm�gT���� �	US(`�d�ju&T2�>�*C�;�����t�`i�.����?�	��6����o��@�8#Ҍ �TR�Y��oAI�|!�	���IU�������o׳E�sB��VQ��*�C12�"\��3L��Y�E�c�4cjC'%'@%���՟֝<�ƀ���ɈR�$��7������@L%u&8@�(/N7����KG*��X"��õ�bc�f��l�v#0H��D�^�0�"�@�6Vp;d�Ș0��$��)whzá�@䊰a3���\�<���� %0FP{��I2�,��j�-�$���cä6�&�A&�?	�)�B��93&PB�."ړ	i�U�B/CgǶ��RfʽQ6�0�P9g� E�(>/j��+U ��e�k�NR7<��ɻ"�
�Q<�&��b�6M���Z��?YԪJ�V  Pb�M��Dz���W�RB�'�lLr0�T6�Z0�D�ۑv���D���q���-"�3&B�Y4)��Ô;2��țR�K�c#�*a���4R�sS�L��?)ި\>=�CT;3���-{O�$�Ug��;�V�S���1|*Ԛ��ΐYx���jĿg+�����5�Ӥ�B%���~�V�	�o��c��!���H��U�ԅ��E^�-Ib*U��,�xW�݃2� ��3�)� ����D!n�����%3^z�s�E�OL�f̏�W{�P"�EvӾx �	Bێ�)�*��Nm���@�����`EÔ@b k���%u�v���	_ dy�$�1�XF{r	]9k��+�/��&��E��& ����´9`p#�+�~\�=@RB	|&`�� �G�,ѧX�$&�Ġ� ô>	|T{T�'e�]�#��%s��k�Ԕd��3����;ac�}ң�&u��{�'����� *5� �R9%��!p&#��ɚX�B!H8�r��f0�����/8n�'vC*��d5́��Y ,<"b,O 7������5(���� "��R��˸���a�N?!��P�RR�5l��f\:vL�fs�� .]�>�	*��C��F�2苺��Eɓ��O0�#��.����PΝ�=�2�`=���4A�1SD��FgX>&�P��>��B��^7?��1U
� R���yӐ�Ö'�>%�X��� �E�6�w��9s��fY��i��S��g߸Re�{�hY��`-�;�hQ�#���/f��P��0��m�u�o}�I	' �ؠls#	�6\#�a�v��p�<��MK�2��M��]֦��R����.��"��)Z3��
��3V��4�p�	f
UH1�>��,��8�2LaPGцN	��S���4Db!�SC�w}�䠟;�?y���8;fu1�7O��3B%��2Hv��� ~ e�FDB���oy�-8F1�@nL�dM4�b]���k M[dFE�y#d�f�X;|��fWWZt���2gl�7G�mZ��:��-�\�b��L�.�d0�֥�2��Cp��9�+T�X��I�¢&m#^�\�2�z�OC�(]c!B#<Wր��R�R�>D1a�R�%D(�Å_�@+���b�J�X���sg����
a`&�E@@�'�_�'
��w��1���i����jT� <w|ޡ#�iٜ0Nؠ+�58��K�睺4���)1�D��t\��4x�:M�7�q.�58���<Q�҆}&����I�J����.%Q���@Ľx((Sj	=��M
��ءOD��g"@�1����Sn��Q���$�E�{/J�
�8��yr���%˚��B?��U[aI[�(I�Ę	�Ա�@Ԭ�%�V� �P�� �ְ��lֽ@��E@5�L�
d$6��7����稘>����M�G; �!��X.~��ɓO�"�AET�x�d�"7+λ+T�'�Z͢NW�r\�*b�م0���҂��\�p����#��m𥈙�!�p8dJ�QpdÅ˘�X��M���O�E�&a��eƴX���u�D�,Y��",%i�D��b L�1�l_(f�}����l-,B��_�s���
���l�X�&"âA�`���i�7�_D(�4�� ;�m(�-�_�X��1$� M�1OZ��q���O����n0�S D���`�&�s��`���7jD�h4��͟Kg�b��	CfU�@����k��Ԁ��7�t,�w䇅[�j09D�2a��jw-�&G6VX���A��4+��� w����~ʂ,�:r��As�i�h���Kל?2�A�GN�@� %��Dȗ�f��_�M�6h���0�2W.8|lг@�O�i�(
���(�D��ʱ��.�m�,P�q��Ֆ5�~�8.��a�`�+p�N�{�VyqcnG�,����8��ɓ
|7pdJV��{�l֤�!{�.���CF�`�f��W��$eE�<�Gi҉���ҁKτ1��S&�.����1T�e�ʗ��\��o»���1%^�S�l��j̄j�,�?b|�t�W�U�/W.�3�Z��6����H#dR��2�Y;O
%��O��z��zv��������q"�h���TA��|�w�I�F+!$J"K��%�_ J�I�!�3A�<.���KߠJ�u��0O� �ďށ1��)��^5L+���	PJHQ�b��	��Q*����s_�@���C#�p��Nܥ�?��	QI \a��M�
��]
�H�0vV������IR�$\0w�fA���M�0���G�eJ�%;��W'Q�z�t*
u�a�1u�j]RE���?ёb׎ u��k��'8����?`GN>S.Y�3�~u��u�ǋY2���U�L�� �*��Y%~���cE#q�2��䂆5|�q��C�J4Wn�dF6DS�3�͑����r�"�yUzШ�'�ܱ[@͞&[�΁0sꞰj$���*���q�eꝊ6��5Ӷ�i�̅A�m��X�ȑ#jޱl+��
����Qr�	HuTT�S�����8�eC�!�F��$���Č���KU�R����?i�eܪ��F��";��c��h!b����(:i2� �Y<a|0�V"V�-뮁��F
$2��{�fo,v�BN�<>��o.H�IQS�	U�ӛ3Fn<	 FC�{��(e�u�f�L����&@5BEx�(Ig�t��b�s
Rf*%� պC͐7X/�e�QG!d�(|,�8�]�E"�~1��C�$�"ݢ-���l��Mh�t��CH )E(I��)M�|��̇�:�
�R�a�%N��x"e�Ll�l���@(F*A�4���PO����ңl���Q 靠4�$�I��=-�&�&	� ��)rI� f���R.2?AԦR6���7�ݦ �c3�O2j.u���[�������5F�h�58�����9 �S�O3i e�����̘�1A�<����/y�, %s��]��(�h˴�W��<�G_�+��6k���O�q �MX5t�8A����Q6|iQd˒�^Z<\[WR��(#�@�2)��4w�:7m���pĪBHW'`��d�6�ݥS؝X�̺�6��@�e)R�; %�Q�֘��+X_J�ӺkW�ջ3�d`��* ���hUo r/��abf�4E��c�Wa6�C��'l0d3��G:D!�&º0���!��F��:4#�ֺ����4;~��e�!�Hp�����������e\r�Dn��	�	��M�ƬK5G ��BMT�.(51���hʾ�ɖ=���"��+7VQZ�`�		�|��@k]3.	�"�a'0�Ȱ�V���1�'�>0 )�[��Q�5�ޝt�PI櫏�H���8���mZ�(�lѡ�I�u�$�C�<8=����m���A�B;7x��s���a�1a�'�%���d�:f��ѡf�~�T�'���L�0�����fR	Y��S�49ܸ��/�'�4y7`R,NP�1��ƨj���A��v(墄%�1I�d��Fo��.�� �,O\�	�TL�*i����J9A�X�4��=����m
Ŧ�уd�Ij�������Ӝ!c�i��Td�U�F��f[V��E̠P�`P��zo���TD.kT���'���G��?NcN��6�rH1�ɟ�m2C�w�R��v��ZI�A	B OgX\BB�Obt@��J�NQ�B�3+JXi��R�����Ѥ1(&7=�\���ջEl�2�ќ;C��*씬|�T�����))��H,�\���,zy���� �P4Kջ�1�j�YB�� 8n�:�����h��'!
� ��+AY�4��QbB@ɂ{2z�r$%�.��3��-!�p�Q���$g��ԥC8<��:�O�\~r鋇r}>l�]w9�,�}g-��! H��cJ�U7>���*�s�*���,9�@h�c���a�mӫ%h���U9$ũ@
ҼS���Q!���%�2aCQ�ȟty0� �sH�KB�>�~:r�N䨘k�Ԙ4��P��ur�=`2B���T����/�|MiW��%%^�+!�T�6���OL�p���N�!Ql� F�j�B2��2w� )�O^�ȥ$@��~B���*Z�J/'n�π �y��"ad��3��k���g�d.�r���:��4���\x�Q���	,���2 Kٌ�3󆕥'۞�X�`�`��5�*5�.O�.��!j�h�^|�e�|rVxi O> �%)	�W�P�'�p?�r�Mp�
�+��6A�ř`�*�l�$<��a�<+Z8�a�n�zg���(�29��w��\�&F#��4c	>b�<�	�'U,���ƈ"Y�ƌˣZ3��1���d��L�:?o��9���֘����b�g~�*�D�@J$腡tڈ8�E��y"��V����)ڐ�GC�p���=Q~�١�0=vE�W����
S�

���w���ҤEŭ�Lq��l^%���͚���1��]wY��"O�`�5��7�����	X )S>�j'�dJN���֥rޢ|�T�w��鉕��`E��)��Q~�<1D���874)X��<b���d���e���$�N�XG��'��!�J�Xp��✠#/�P��'r�d��h�0h�qzG��'u\�M��'��QS��{������/
TU�Ӥ�Dev�ؕ!D�l,��9��#�!^�d�B蘳;�!��͉V�6�ۃ�%l>�t�1�!�Du�(02����6<0P􊎪y!�D��'���y�ქ3�(3���xR!���0D�9lN=`rh��*Y(P1!�d	���M��Þ.F��жJʔ?$!�A��H ��w?	�@ۖ�!��DXN���HH�d9�Qhb�$$�!�$�-j�ިq���d��(ElC�E�!�PRT�s��B3��a1���5�!�,_D�j�/}�V�놆�:�!��2 £��D��WdѺ.�!�] �:�ï���!���]�!򄇴/�*����5mM}���"O}��؝R�2������u"OJ���O�N�ʠ
gн: ��G"Ob����;��`� č��"OV���E�|;G#��O���"O�l�`AҮ?�(��A�o�Q��"O,�لbQ�,�8h%?�N��!"O@��Z��trao�g��9��"OZq�&��*�"�yС� %�pс"Ou���0��`K��P&9�Be��"ORAs��#;L���AX2P���J"O�x`�s�"�OÐ}��g�'��KAD�,bH��Kկ�~� kŬJ/�u��ą1N�Ɣ�3��*_>q�L�M͈T�o�9d��]�3Mn[��s�p��GFZ>�0���G�3�W�Oβ��@'?�w�O.x��a+�	�N>U!���J8�|D"șP'BA8d�f������A%��e4?�~:D���܊�a�&�	Xl�ٶ"�;@��=a0�D�q���Ӯ}���y��ƙ8�0�9��Q 4rV�O2��<q��3M��i`���k��I0�gL=��1��:O�,�<���[c���0� c��XQ�F�"&:�Ӻ#EAZ���c>��#!�\h�ah� �j���*A
@9�ɕ�?�$ ����\ib�p!X� �Q�!i���M>	�4�0|�p�N+���B�%�`�>�Pĉq�I-`�<�XԩXq���OԺu�@&,i,}���Hb`$��-O���?)�'g�]�>)�e�$XF�8�OҔ~'X\�pIFYdI�u��OD$`�Fg�_~2��1G��8�T�0Ud"�I�5N���?CM p��E�3bR�5�4'��^�1O�1�$�d�S�'}Wb�Id.޳qg�q���Iu����'���낣%�)§r�z��BˁQ2XLi�^5	� �.�5�%�)�'dVͲ�E�)�\�q��2]%d�o�*Y֠� $� K2L���uw�O��9P�
:\����H�T�%-�����Hy"j:�&|�t@�-�������%�I�r�i����R�� �O�?�;�燡5���`C��R�4(`��S=s{�I����g>�C �x����6�V-M�
�G�>Q���0�"��ȟ �iԝ KZ<����f�����j��D	Rr9{�" ٟx��g�? �����*#� y��nX.:��,���Iέ:�(p��	�UR����O>@���֑P3��:F�G	>��'�D��Qj�?t�`��$��)=� ���'�j�RP�ڜYN�a��ޯ.ŉ�'�J�@�/�d��to~��'}2h�'М+@�m�aǄ�|�́�'�"h�����Mzʘ���{2��a�'���I���RB�� �\nE���'{28qP�V��HY@�J��*!+�' 6Ձ��ֺU�����10��
�'b"\�p��.�҆&ۛ�v|2	�'0�k���{j�pӊ 8	Ӑ-!	�'�z��e
3zBL���{5��Z�'��Ag@�K�@�+�  h����'����2�Ɩ0pPX ��0�4���'��P��*E;#�R�h��8#���'�48�R��z:���l��b��T
	�'͔����ܑ�b� ��
��Y�'�2E�`ս8\��D��*h 
�'����ɉ�]+.��``z��%D��b�"�%7��@lE.S�@���%D�DS���^��l@��C�E���{�)/D��k��!f��AL����%��i.D�HӲ���^4]��342����*D�L9��^�1���r�F2^���5D���D���^�J1#gi��x��`Rb	5D�䢁���%��p�B�s5��Q��3D�`�pe�S��Uaj�E�h�a��2D����  }������&�`K�b0D����-ɂ �����o�"�9D�@�(��Z��iZƤ��d����4D����)]jv�㐏ِO�p���5D�Di�c([��`kT�hy�렡.D�ȲA돾">X�%��&�na�e?D�@"�K$Y�(��GF�&�p�8�a=D�D0�=�p�x����u�1�;D�<�t#�"gK�e�l�n�&q��&8D�T2�H�'�꼨$�D�{a�H�G0D����f��`UFκ�0JA-0D�d�4�.T}��b�L:qϊٱb)D��I�g�*n7$���ɶ�@�TM+D�qS���Il!҆���6� 6D�0+�F�4h��pz&����RF&3D�\�e&6�cψ�1�Ԃ��5D�p2�ʷ	�*)b�ɓ�Jp�`�'2T��pvW��,��N	5��0u"Oę��d`��+�K�"k8� �"O�m@�eH~��A�jc ��8�"Oyr�o]�VmAwC�e�T�a"O��R��^�[X�a�"�*���"O��Ch��g�(�(#!���%����y/�\S��+�|x�S@H �y�Ƌ�4Z��e�()'`�a�=�y��T�DQk��W���RU��yr�.h� ܂L���BP��y��)���`��B/��ڕÀ�y�L �F!��d ���A(d�`��w�L1�-D	v��0$>�x�ȓL1�ըc�ڜ{i��kC�`���ȓ'Dt5��=��=*0/\2O\��D��d�Ђ����� O��uN�t�ȓy͎(A��ŋ�����H$����(���F�m����ۻ�<<�ȓg�b���*Ӎ"Pb�C���v�����S�? |u�q�U�q���	��̀�$"O�2cX��P1,��Ҹ��"O&��cP��hMu+��i%(kG"O���h�q@��(��T"O� N��l�A��wK�( �"O4P*vGG�r ��, f�L��b"Onu@!&��-�ra٤�V>d�V�ٴ"O�u�͈R��!���G¨���"O%H6�W�5MJpp&�� �dr"OJ%���� $j�8�I��&���"O�8����-er�h���P��X"O��hq�*~�ۢ��[��)[P"O��3lô�9[AIߐ��Q"O�Dc�k�7`�R��5H��(րxx�"OVdpTޢV��:A�&d�2"O�P!�N#B��*��?�]��"Ov�k�����<}'�:5"O*�X��$Y�:�ÏhXk�"O�IBW�52�%��'Z���"O~<�u�W� �2�kҶ�$���"O
�z��,1~�lP��Rd�0W"OT��7��"�i[�\CT"O��h��SM�vH1��:���2c"Or�㡆F��I���	^<!�G"OH�{v��&.� �@\���r "O6�	��	&�NmZGS�*�ŀq"O���E ��]SqD�0_4�m�1"O�,0��Q�;���ren<����"O�$Y�MG�4���m&W�lc"O�5�En� �+-S=�ah�"Ov��UJ� �O���p3#E?/!�Άu6��%S<:,�ba�Y�!�E<���s�hG�~*N�x��!��ɏz�̽��l��F|�+��;v!��ʟb��[�g�0��)��	X�d�!��/=Y��Rw�i#��"�\'�Py��'f�����A�#$��ShP�y"� &M�욇�x�lIq�\��y���<e�HmS�On*�0"�@;�y`^k����[�Z6a��H֬�y2�@<9��K�}gb�A�!@"�y"JC 7 h�Q6�J�b1 ���4�y���p_���ƋH@�D��@"�yr������=H�t:,Ҏ�y�B�>@Y�G�:�@SuD��yBH*%~�#��N�2��M���(�y�$؉8��ۖ���ܱ��.���ybꅤy����ʺ|�I����y���2�x�#���_�4sU��yb��q�@X9�F�*PZ�Dr"�Z*�y2��/6�(ᒅ��L��*���u�<ᢡ�(~.
�U�#�z�(u�L�<�'얇f]���Є޶=G8EH��p�<�$�I�wjp0��:Y�Є�gWT�<I�dQ�C�ɣ���-W�����L�<W�״�V�* �G�+����I�<���Q�{_¹1tFE�[�
09��D�<Q�!Y�([� 1�F�hW�p���
I�<�3Ǆ�q��i�ua�@�P颴��D�<�)^n���u↖V�"�E�F�<Ѷ�D�-�i�@	�:||�!`�K�<��H
��F�9a�T �6=��n�n�<!��?K��ъ)�*|�d��P�<9�̀9L�pu� (�<R}�0	BL\d�<� 0ܒ�jJ!	8�yI?��9�G"O�X ��Z.g9��y!��-t��  �"ONܘ�鎩~�\�8�/a����"O~:�"��j�&YIǌxN�T��"O�|P.كdv��f꒰8I�j�"Oz�"��<���0��	�FP2���"Oj�8M��M�ല��Yz��k�"O`���^�h�P��"����s"O�Y)���Q~��	�].���qe"Of����&|�~d�Qi�?m���"O�Q'�M�7x��;ph@= Ʈ��W"O:0+���N�4�Ӳf�9!���"O�P��� 8�U"reGT�+�"OfP����֍�i�ka���"O��s�*~`��n[.b>�I�"O��6a̶P��T@�lO�},%�5"Oj=8P�Z

֠ �5�1H �3"O����x�-�!����B�"OXhW)�
����#	���Y�"O��2�)Ƚ⦄����H�L���"O��v*ɖq���b�Q�9�<l0"OƸ���p�����-.��a�"O
 ��	���D��#eZ�Q���[�"OT�2���/g���A�Ǎ�<�R�"O�QkEd�!p���b!�L�<��"O�:�CFw�(`G!Wrݨ$"O���&,ֲp���=id���"O�����Gn�,��d��{���"O���Wž�`)D�L���52"OB���@Q>HlĊ)͢)ǌ(��"OT�2�$i0�Q�+M7eϊ�K�"O����A�;����)��(Ȥ@k�"O&D���Մ4>^)��O2W�M��"O�pb΄�6Y��c���C�qS"OZ��jc�����ϝFgX���"O�]Cu�
�#I8�Y�`I�w��D"O0�@��@$E��pt)-8�h���"O�i��ES�<L�mՠk�H�a�"O��aC��7�NpAҢ=5֬� E"O�m��f��uJ7���6���z�"O�`��א'vP�B"�$�h�Ѳ"O�0�s`~���C�K{�P�"O�P�³G��R�ѓ��<'&!�շ!Z�����̙Y� ��=!�D.
g�"`ӡC�d�����x�!�$N�+!��(�هzp�]��M9�!򤓙 �<�������>=x&+��!��O�h���!7�Վ'2ࢩR�x�!��B�lr\��D܈V)�)V璳h�!�D�uKY��〨4��a8�.W�!���|�K!�	�Ŭ�7�*[{!�$��b�����3t�@U��'��D!��@f��[7HW%%�f���F��!򄍅Yl��D@�M��XS�	/�!�֠�2"�֖hd�³��c�!�DR�J��YHƊ�5H�|�cA�W�!����B�` �X��rx��oP�4�!��_$1�H��G����n)K�!�DY�:#lm��Ǝ:n��hydM��!�Dۏjr�*S����ˈ�?!�D$z�͒4ϐ14<�8��i��`!��	�5N�hwC�#u.ǈ%�!�DT G��ّp*˿B"�@	�M«l�!�υ0-���홨b~t�Xp�8Z�!��  Cb�߮dXHt`�力#�H`1�"O��ɝ?.��z�/ܽbf�Ж"O^�pW�_5M��)���%h��`r�"Of�:A�DG��@t-���a�a"Ox�Y��['F���*g���x�"O���g�ǂ}&|���+e{,�D"O�x�   �   �   Ĵ���	��Z�Zw)Ė;"�����@}"�ײK*<ac�ʄ��	�$5�Z,x2�L	q�6͞�:~�x!kWu����A0�󡌌�.`E'צ	p����u'&F�Z��]�Y�.�i��?I5��cm�����y*Ȓ�oY��]ve�<�B��8O	V�G�>aLZ:g�&͚�;��������<���@�v���'!��3�� �L9QΟ���!���S6�
b�ǓQP��`�O��`!cV�Y:!��0%��;��0|خ�%>�{���j7��CX�~�� �ߒ_��es 
�A��6s����	�x��^���a��s�px��{�K'���(���(
'i�3�:-�H��r�
�";��O�xɷ+��T3JG�&3ژ����3m��I>�`���d�0�$�(zģ�l�i �ػi"��p�Ώ�eT��Kc����'}P���LWy�O��A*A��V�,�� b #e� K���C��âJs&�J>A��UHc`$�P����LR�+�3He.PR�ᘊ}p!�/O���	��vmA�E4���7B-C��ilL��9��BGA)aX����Y�2l4�1H>��,��:L�T9�O��EMZ�EZp�W����h'��4e���4$$��_P�����|b�@ �ƌХI��J��%$�~���B����	Y2���EƘ��'~�@�����
1:��

�2%蒥-���B����D�0���	!*5�	�2މ'�|@�p��#? �����6��XZ�' Fx�\�If?-̐��UD�{���P�]�$ �)
aL��ZDY�wɐ(yN$ز�"ԔєO�:(@���{�B��F���L����5*�L``��$fk�(�⬲�.���2T��z��x2	,_6>�(�T�T��8���5� ������G�� ���H̓5�Z$��.ȷW�eP����Sx$;!˞�y2��0 d  �� �  ���h�E)�g�<!a� 2  �@�?�  �U d  �-��!ӂv!�$O'��=`g�o���G�^(i!�dY;*�� ��,�U�r���'��!�dE;�r�!��tzܒ¦Y�]r!�d�+>��ex�g��{��4��DڍCw!�D�NV6�x��X�B�d���2U�!�d�!Fpj8�i�(l�>}�`,2�!��
L��� o��N��hx���" $!�DO=@���n�b�bӴ��!�ċ�2�hxtk�&�(   �  �  X   �+  �3  ):  �@  �F  �F   Ĵ���	����Z6)��,p��@UT��C�ֹS��ԡ@#L%~�@�$�.?���D.C�'ll\�02�hY�`C�a34����U�=7JY�d"OH��-nq~�Y��-H�x*Q� 6%\p���L1��"�����"0���U4]aՠ'\�R�jЮ89d敋D�ńN��q4 �Uo0���Q�vж�Iw�0w��MEJ��GK�+f��@���	�kp1�u�)z�v�҆N�xR|�E_G�t�SCW''�h��∑p(
�d#�)K��A"���?i��?�S���Đ�?�P��\R"��3kG�OrR�"�N�����ɚ7Ҟ��v�� �b�]�?#=�CD	�1�l�m�_�(��bJ�%pCL;A�\����O�q@�2����	4U4��A2Gt�Q��a�=	D�0)��F-{nA���<����(��4&8�'b�'p�䂢 �F�ȣ]@A� �*(��P����ƟtAI|�>������I2��5����RЦ[�40��v�|��O���[�t�ql����P�F�
6����&��`�:x�eI�ϟ@�������>�u'�'�8�"i��h�1	RƈQBkԳ2d�@�=HՀ�ҷc�CX�@���'�)����kx4��W���f��r�Wݰ>����`9)Zy֦1� �� x�p�k],F�nZ��ē�?I�����	��B��!aY�  S�D���u�"O�zQ�_�c�ѫQ�!0�V��W�8�4�?)O�|�!τѦ���՟��'c��0���*���)�)�X�lڈX�� �	���I�?�&=�dL80`$#�+^>7*���)����k�01�������JB(�D{�GƷPhl<30NF�XV��� ��~L�`��f�'Qd�kp���T��ψ�]z�pSB[�`����O4����'I�6�E ��S��ꀘ�(;V��|X E�(d�tt
�4�?������4}��Q!�M������+o4\'��G~B�ӠHn� 7x�`ď�Mټ\@���`�!�4,��f#�"3E�Iϟ��I�?�)C��ß@�	L〬�#�Ѿg�$sր]��H�޴}*��)A�S�Z�i@�i�47]>!�O��IY'<��UE�tY�����6����Y0c<�AfcQ	hB)`���`S�qV�ty2�Б ���Ӂ9	a�d�Zkȅ���ìn�~�dѦL���']�)�)-}��4|ܹ �j������y�`D�}x8Pr���a5�D�g�T��HO�hE��b��3�����2;��hSw��30�7��O:��^�,�����&�OL�$�O��$����[� K'i��a�
�HJ:P�B����8R�J�KCS<D�x${6.� ��3�C�]��!�#��TB�$˥/�S7��}Rt�R(��Y��ۑFNg��� ����I�J1�V�6�*�ᷩ!C���ԧ�<�p�O`��=ړ�~�ȍjVXic���g ���u���x��Q4��CV!9t)�
ݒ¶i��#=�'�?�*O��y䋆T<��3�݊s��J@�[��a(���O����O`��[ݺ����?9�O�}��ᘉx�(kA$R%Q��M�A�&N4q��F�!&*�Ut*vџx����F0i�@�(��8ʲ�Ȣe�Qy�ț6E&4�3�ͳfR�[��BD"<9�CH���hVe@/$�|���^
c�� �'N��MK���1�Ld � @ہ^�<J�D���T��	w�'A�@k�#��4X;�#�gn����O6�o����'h�p)U��~����DG\ 2őfc�%(���97Eܶ�M+Q%%�?9���?Y�c�%&:N�r@˂s>�+a*�#R�铈W��ǚH���-0lў��g��KJ�]�w�����}:���6^�`K�n�Da���N"B�Kp#�>;�>#<�W��@�IQܧst5����͈�� G��D7|��'��~R�K�5<|\����6��l0�A����hO�\^~���d�D|3�	&0�H�J��V6��y,�d�O��d�|�� J��?������(Ѝ)5:�d3b�
F�"��r�i��6�ʃ|(`ԉ�n<Z}L$(��~:���-ֱ1�@���^	$H4�ģ�E���	��48�B�.pR�aX%h�*�@4�C.Е��O��@1�ޭW�Z��=�qg�'���B���?�O�O�$�1&��wK�}�@8p��6D��r�ś�@��y�a<D�,(:��.���S��4��xS�a �`]B��B��N��	8eόæ��	㟌Kd�)b����������Xwg�L�DB��=�鐆�W��$H��L�q���C%y���𲭠|Fy2�A�e�:rF+
t�%M�:KZ�0�`�,�C��l�y�/�Q��1�&�$9���ˋ�4[�)�Qơ<���O���>ړ�~2�A�/���f� 1R����F��yMC;pBDj�/W�,R$�D$���M���i>A�Ipy�@U�'��!��4Xdx�г(�/N�Dܳ��j���'�R�'���]�t�	�|��IP���=�g�w���b`I�־ ���*Q
ux��L�hT����(�t�(%'!tX 	�۲N'��R�#@	|f6�r��Pmz���&�dJ@V�p�@�)��,ھe�l�n�'�Q�\K����QL�5��I��E?D�d���>i�F̈́�&p��cš>���i�R��d $����O��2V�8١��{c��yŚ�n3�7M�6����O`�dĬUD�H�b��<�� L.R��0Bv��Igz�R�Q�xXA��ʗ�X3����*O{�3ܦ,�����]�aG^U��fs�? <$�BX Fđ��ꓼ>�"y�%NMH�'�҄���?���oY�k(Qr��H�xc����$�O����~����g"{}��|̉'ў�ӧ���ψI��=���U�4xD�BB����������4�?a����H)�r�$�O��A����0�Fv\I�G�Q����W� B  �Ѣ�+�M#hV��)�|j���k�%�NMh	��Z�Y:���d��OZ��g"�Y��ƥ�!}���僁N>�� ��)M
?�X�Y�ʲ{p!�R�H�lh��՞u�R�'��6��O��O ���O�
i�`�@ ���*Ր�J8 �S�d�	C�'}�zT��aB��H�y���`�a(������۴(�6�'�
7ͼ|V�\w����,s�j}H�'ߪA���'��.��X2%�'!2�'�r�o�%�Ɋ;!���]w�{�ی?�>5A)O�`X�'~�i!C��$��M@����KHy���p>	"e�6����  �)�Dy2l��?At�'�����	*cf��N�O$��'g�AP�H�q�p� ��Ҡ��شw����S@�I"N;PX I S�l3�E�w9�sA�  5c�,�	˟��I����_w�'B�σ90�ppƚ%^� ݓ�����@J�"��E�Xҷ��&i%��y�4��pp�Ҧ_��S�[�/4��k oQ�/,����S�3���aDE�?�m��$E�'8�$p�$�"kſ�������p0� _��0�D�O �D)�i>5!�䄾P�|!!�P!%4�i�a���HO�˓�(OZy�ݒ1 �(����.sI�R��i��f��al��0Cٴ%�la9��?����?��^�Ur�`�-i��́��J�
tlZ:|������I�&�� ��l;h�@Y��ͩ� �y�O�ʰ�wB�]p�!���)i h��d���>%QF�Wipx{ d>5"���/G�����+a��X�J� �%�G��?e�f�d�O��>ᡕ�2{�2��s&P�(�n��Ⱥ>	��I>��`'؂ �t�<�8Uq��m���N:?y�)BKEp����M�=�'�D}ǋ�q�2�'�S>Q[������I�>�����팋4�4`B(�k�8�ߴv�jM8b`��6*H��+N���7]>	�O��W�Y\S"�<���U��>^����*��y�`����i��'V7-���!o�%�ZQ�VO%hh�ɕ*0��Lt�	6Ӏ�Ӆ��**؈�D�@��':�)��!}"��F^���,�fC�f�C��y��2
vf$`�#�[E�ixf����HO E���¨#)p�
f@N*842D�-��pLR7�OR�d��R�i����Oz���O�����[�����R,Ά{��=��&$3&�y)��i^R/� B�|2��d��1ő����c�8>�lP�.X�2<�18�D0�n4�(�Q�L:/�C@tTS�) �-C��
�l�<�qM��I����?���~Bb�<P�E�՞�:��h	�M3���?�A<?IBE-7���C!��,�<�V����>�*O��O)�V�ܙ�T��}���ל_f �+G�N�J�ˆ���|�	ӟT��2�u��'O�2��i�&j��}�� ���1FV�*�7 �ց6�0%cFM7z�?��"H�oi���W鞁<KF�T�
�F�v�C�M�T�t���bĹm�v����<���Gx���?�r�����͓"�U�I�n�
dj�����G�'��8�����y�=a'�\�$�(���(ON�	抜-J=ZÍ�l"��!�R���4�?	.OX'j�x�T�'*�i�^,
�a�� V�:���B�L=��)H�9���'���/B�\��2�/'݊���M�����$��<�1Y&b��H�,3F�=�C�9a80�d�ߑog��K3�!9v4�Ü�!�ܸ��O�8W	�M���^V�)��l��!���'���k��?����iʐU��Q*E%�#2AÂٗ��D2�O�H�tÊ��Zَ%��J��r�a}�*?��L��+��0��0A�mZ Xt}¨ܿ0��7�O��d�|"G^��?��)��@����SLٰ��8E���ih��Ì�;(����ΐn����Y�t_>}ϧJL�ҥ��1��;��l|d�	�2T�데p8n����Ŧ%�d��-Wf%6-��&x�OZ�ywk֡p�
�t�ܬd�0IA�'�`���j��h�<%?E�K?y�Y;'���ӅBǾGH`�3���i�<�r��V��1�V1����i����P���O�	��L�e���G����� �ɒ�IN$Yt*OX���M���ypQ��|f���â+D�d�1͆�zV���C�	eJ��o7D��J�EH	V^Pt�'+��[�J;D���s"�3r�x��͘� �}X��&D�4�4kP�V@�Q�̽M,��Jr�%D����+��Q�<j�%�q�J���&8D� q�A�	�8�8G�qU�� &D���2�Y\��+�B?�
�1��#D�� 歋� 	�bz��!�D���"O�]��Ă� �z�3��\%�60�"OX���&}´�(��R�b,P�"O� @"!�^�P;�菸3P΍��"Ozш�C�A��j�M���څ"O����Q9(��8QQ,�%Dʘ��"O��!����8dY�b��k�� A"OD��aϜ���p����@]'"O����M�d�ǂ/H	0"O�P�#lA"�!b5��:V	�x1�"O2�xd��<Y�E��`�.\�48�0"O�H��&	R�x��@���d��"OZ��&��i���)T�T�z$��"OB�YV��qR9۔b�#��5�f(L�Eȁ#��mi�}0P+P�K�>�d�ZQe��3?@ ��(N�ЄȓvxT钀k+�!EM%xv�j�C�>)��ap�
�1���X�c/O�����$��c.ܳD=2�'���0��$"��D6ͨ	���y��D��n�4O�K׈�P(<)p�1,3����F°�#v��x�f�0�"t���Bg��6��(��>�5��w
�tS4&�����Aq�$D�|���а o*XYF剣rq��3��)�	����%Ԟ9(Þ���"|�'��I�D�)wXLU�a[%'�~q+
�'��h���TE���*��A�kF�V��KW��^)ޡ��'d8�D"Ac�/�.IsB'^�R갪3LO�8���m�tZ�!)Z[�,i���")���9%�,-*wI۲�Px�א}�zm{5b�;`	��Z1Qژ'I:�[3Yz^p�Ӣǖ�ƽ�}��]F@�bT��4�ԍ�t�<�&P/���P����.���aiƜK� ����.U���AI&Qf�D��OL��bֺ}���ҐEN-\g.#�X�(PV�)ʧJ�(��ƚ ��8󀪜�k���k�۠Rj�c�O(�ػr&.O.-��ǽ1h� �5R� �|�ظ'Hڑ�'il�sa���*�Q6�ގxI0����3^�,p�v��{x�p�w�jm���2��B�o^�cx�t0�y�kF�#��u2���&Ox� 4aA�'_Cp��FQ�%�,a�m�YӰ�D~�+� t
j"|��k��=���Z�)�*=wRLY���)
;�I�wcˌ%B��w/͔UܜD��Of���^� �W���U�!�Oh�AL�
�1O�>�Ӏ�J�wJlݠ��ڲ���)���)-*%{���-��,	e���R��xĖe
H���ٌD�W[5k�'Of�"������mK*�Dуye�	Ӻ�yc@�D��� �fܚb�(;��$���4�@؃1,Y�%�4|��!$H�n�A#�	�d+�9Y޴O:�� �`�PHi�-ɪ(Ζ4��'Ј��|���1���n�53F�=�rGљ�HO���V�ƣ�?	��� �nI�%�O�2(��fF²��A�\�ȣ.�	)�6�ӑD���qK��I7�|�%��"5�`%��l
@�t�ߧ�.)P��>�|Ji�$V���'&��2j97��R.ԙ�(!�Gd��o#Ɛq�H�meB����:O����+ղ!��ЧM4#�(�q �'<R,ƈϑH��E1���;G��ۈ��O|૶ @
)kf���) �q�$�^��X�%k�!\0H��*���s�!� T��JÔ!lx���G��@qᑏ`0M�ɖ7��S��u��1�J h�`hd��5	&�	�AhvL�u �<j�D�a���X�4!���80)��k#�8mV��J!r�܍�f��b���b� � � ���P�V�h%�	X≏��j���8W谅�0$G'z��%(��&~\�q�K�?q��2�k���(w(0��6(_'A�����R�6�p׮�Xh�� � II(�a�,7mZx�1��HB\��zI���m_�-�,�t�)^\���\\�T�4��*7���	Ë����՘�a��Y�6�c��a�  XgnG���<a��<!] Zcfw�i�@!�S��M(C�v���0�$^Tr�:��ŴR��Xb���lc.A�_w�N�q3��c���,�.@�C)o�e�G�'9jl�!R�E���t`9�I�b�NH8�$�/}rx=�Ukx�iQ6?:d��%��E1�� ��;�ޕ�q��|��Zgՠ,�H�G�M�Y'���#��%�V��1�I	ri(�J`$��TQ�h!Ӣ
����"���DƲ�H��6�?�t����Kb ��4�8i"ծ�-�0����?|�×��?梉Pf/[9��)�ǧ<I�I�g&�(%v����K?]k�<�a�U4}T���vЛ�c]�'�����B�Q����§�V4̧(z���/6P��ѵ�,dC�I#΅c�4�����&1_�{2D�|�m��$��$B�˨|3�9��ɚ>R:���UA8��1�x^,� �/��%@��~�f�O@�̻���P��ΐ\lh��wDQ.jʁ�?�aK]P�t٥NO���'0e���/��8�0��>4F�PGƏlĆD�r�ȇ��}@g�<��9�O�(3	Vw
����Ns��h�(�r`$s���
��韦�K�J35r � �e�|��䬻ɀ �i��O�)�A���F>
Q,8�S"O�<4J²V2tQt�P�$���`�X�������{�Z$�#��'�#mi�e��VA�ӡ+�� ��HU$z�\�q��R�*a����B�j���	��(Cd*Л�~|��*e���'��$f�����7_@��WJ ��/�ɌWD�|㗆A 0h!�F26����$Ɯw:8�C͜gGr-P.Y�&�>���H�S�T�zp(�2%!j��#LO�xG
�V @�)Q��l�ش"��	9tF�'�\1g�2�aՆZ�ސP5�Y�7������U�!Hpa�!@MG�<�WH�=�5�F�7YX��pP��IyҌ�+�`�0�Y�S�`Q�OW$&>�B���m�f�9b*]|*��VF$D�Ă�A�!zAҝ���2^�x����Wۤ�(ř|�^ �3��O����qO��K�/�-���LP�Y��'�h��g[�C:|��fUX���\�6��7��'(�6��WI���p=�$/��m�P�
#f�c���Cp&D�'6-A&���X�٩8Фȭ���@x�D�z�Z(v�R8_0�ȓF)v�:Q�gt��RA��8��Y�O�C��L1����� ��*"}b��G|x�Y�υ��H<s�L_�<idC�\���Z�F�(+��1wa	��6�����Lyb�̥e��&DX�]�YZ��XQ$�\�*e��+<�q9���,R���$���T��X����C�~� ��(�0>�1�5XN��2`�|<�m��H�K��Z�/5l<�'�,�0�Q�6~�r��	�'���Ql�UT�,XB�S�;f̋�k׬91a��([�SCpP�A��_*�=������y���3ߊM a�@)t$d1�"�y'�A�
�)pNrQK5LX�y2 ��m�*v��Dɪ�buoϫ�y�-�� V���0u�r��)���O<�pT�:6���
Z���e�3O��i�I�4JE
us�o�{Z��g�C��TH�V�X'G����e�'��hC��z΄@���d�Ƽ��'T�	�5�Dt�\�H�cԛz�i)OP(p�'I���d�7R��Xz��+��}S��۰v�!�$%���5��b���V*ަr
��StlW�|���և21��R�����yR�!A�l|*k[	�y�-�N�� B�1>ڭ�u( 9�0?9���hZ��v�yF�LI��y��Η�Up�Pch_�'ě&��)O���в�C�����P���'JJh�f)>W,��F�.K�zxQ��DAM��e��뒕{�T��c�J?��e�ȸ��j�
�IelZC��9b��@,&QŦ��t�az�$�GC��%��\#	#�yr�Y $1�Q$��R�1��(�.'G�A��!e�]!l͒�pv�ޡX��bbR�"i�l+à���yr&��c�&,�UY-6KԸ�j13�2I8 a�:U��a�@��h�f2q.��#R&-�WQ=V�T��f�yg�W�t����6DB��EF���0?!!��*�CelP�4����0�ۥz>F�&M�t���K���-S:]��oԭ!R4�Cc`H�TI��6��U̓zOP)z�k�8d�`�����EG|R�%/�� �2l�P=���ۈ5�P�+���zՏ�U����C0c>��EH�}8L2U�9�0=�Յ�+���
M�X���<�n.�Ӣ��(က�Ӊ�(o���**X��
 (��k��Z�/h<��Sh� a�i�A�_X�x����F�u1m�� �1}�y�9��R��*�0��Y�7���"ə;5�l���]A�z�	r��ͻڦ��AIPl�7�X�	��-�O��� g���y�H˔Bs�O����d��	��`�3�CD��pCK�9_�x��A&��$A&��i��͚j�Ta�5�[2$��sE��ʯ�$��@nL�<���pG�`����@B*Md�U�s���O��0
��|M���FbT�\GJ��rC�@�.����ɷC��pH�ś�v�4laA�E�Kb�}9�G�t߼�h�@�6VTџ�ϻ'.�I�C ��l������{�|y�*��_DP�ʔI��<���اn2�>��c�{�a�[�M�H1R��2
fmв/.�dX�l�C���L�P2w`��=�o�Rњ-3RCɲW�>���K*3H] ��C�-xs�[(Az�I�&K��R��ݝ/!���2����{R�
�^�Ġ�b���~��F�wp��b�(�U�n�KA��y��(�YroU2�,���	�!���B��޶j�v�2d&?���ߍ-U���mجe��9�6LN88H���<9g�!L�h���A�{7��cA�3|� ��F}��>K���2�i���OV���ذ5����,9iAIʴK�0p˄	K�Y>��%Ɂ�V�$">�r!�À��S���fE*e�ܰ�&ϝ?_^�3�IJ V�SdY�Lz�ü|Rȟ���p��ñM�w^(�CO�9��dF|�D� ��Ȁ����H1$o���y҃�t��Q8���,J �k&_��?Is'	�C��¤����V"*G�8��A0m��	��?*�r.C>!º�
�i��]�Ƭ�Q�t��&�� ֩��f�]UJ�Ι��4�F��S�\�����/B�
�nX#W�r@��C�ɀ&n�rC�5g0���'Rز�fHO1O�U:F�%}1&�a���P�V\s �M�#tP�[�Yu��W��zN<��V�If�Ș0�F��N
�]��m��$6��{�	+�\}��ɵ<]�� (h�T�
�ewH���� j<ڌ�����
�(�Yp�~θ���9O��<)�d6!�1�pNԨ)����S<��O��w�	�3"FL[�O��J��i��<� 2s� Q�Œ(�F��ݴ'`eCb�E! b
�Y�yb�U�?Ym�_2b��1�@v,�xey�D��xX�'1 �!t ۣd���
�˒+FqX!9�S��(N>V�0��H!D����5_��0����(�Z�<����Ȧ�0!���p�⣁7��'�ְ�&o�2�.a�.N7:��Re�*rV<#G�����BO�*"�`UIֺ��ԟ��S��* 9�آR�}8�i�A��%����,(�&�������vhPo�:h�$�/:�a)�oْ]��؂��O��ϓ2z�,ۡ%H���g?��>3��رÅ��$��Ч�#\�Fp���.W�
�̓&pDũ�:�č��e@�Ba��t����< \x�Y �I O�V0�K<��i�<PY�`_]�(<�;S�"=@͇$�����d�MĬF|b"F���'`�4��Lܦ��JF�x�e�)ibup�6?��!bӤT�������ɒ�m�>EZc�|R��6{�ՒD�� l�Q򑄇��hO��b�Aݮu$�q�)�*T�%�'#A6ZTI��/8A��#��"�A.��t�����Xr�ɓ%�}x�lJtS�j~�;G�W�(4h��O�ũ�����Y�JS�v�PlIrC��:C����ڄfC�+d�{F�7h�db�$��gD@"�"O�K�I�Q<9�7@PP� I�@��d�L�4g���O>�&w?��4p��ΐ8�D�tc�!�� c����}��}����]ތ)�w��`�h=���N�!���P�		q�'[�"�'b �9d	�'0<�H0�dV$��p���G}�bYi�O��ў���I����JϚZ�R"l��$+H�x">�R1��-b2���`�M��?�#�U��� "+;lO����#��G����,͔n����'Ӻ0bV.K�<�ŋ�+1��@6#�
;�D��@c�<aF�
[q�W_1r t��j�'�T0!�����!�����3�	'<��B��70L�Rp�� 1���X7O�$B�jC�I2fR��Rg��n�6 {��ID�B�I�[���N�q�lYѵF�	v��B�3�v��Gψ�0o&	r�Ǜ�{��B�	h	�L� n�@�!	�f�i8tB�	>(�!����gkF6�C�I5t�x��L.tP�AL�h�B�*}�7�ǋBd�T
��%��B�	P��b�!>$(�N�#��B��8zx<((P��b�4+�בNMC�I6Y	��/�:eȼ�U�Rn�C��ll\�,M�ty(G�Brd#�"O����Ĥ^��a*ŧmJ���"O�T�f�5$��`8ł�3�"$��"O�0 ��n�P� مD- ��a"Oؕ;����@�`@��u�"O*�Sei�8
܂�'K��yf"O*1S�d@�z��qZ���^n̸W"O,���@��0�'B�#[z6�z"O�[��S���ur�댄-J(I�"O@e������2���m�M�7"O�AQ��RiP#5+H���<I�"O�"ᢟ(~�ձ檞 S>��G"ONe���	W�vpC�i� W�,$�E"O��D(�nu��;��H-,�<�f"O�\q�S-WP!�@�)e3�)��"O�d���ڄr��y�!�׌YQ���"Od�! D'g<q���S�P���Pf"O����	�sH���k���y��"Oxd�1��tpb���c~Ȩ��"OЕc��׮r��� O�j��aZ0"O܃�ҳoI0�����3$T�A�"Oh��B(!$�t�&��B"O-#��&�|{��*LZe�"O�)�d�\DL,�ņ�"讴s���K ���G��BX���Rjߕi��4�D�Ϛł��;D�TJ��E�i���	�� �-i�C9D�����O`���I2Got�[��8D�aƎ�+JZ0�B�	ǣ+�RI�d�:D�� ��Cm��q�!R"���I�s"O��;���9��(1�oȳ=Ȟu�T"O��c������p�ݡ{Qn%�@"O��g�
�l?�Q�F^	
g$���"O~tdh�TP0��EK���*Op�$�ȃ7�����J�����'��`�����r����\h��'�ҍ�ģۓm�� O�ǬY��'�ޅ+a�7���(��qw�0��'��X���P�lS��k���w��ĩ�'����"��3⼛R�U.8$�(�'��%XbOX�����!!��fJh��'\d�	��9>)�A���XTI�
�'�j��9��JH�:V�(�
�'�h�AQLtZ�4�KXp�J
�'@��bq�٭J;F1"&��m���X	�'4\��ET�of�!�HV�j���	�'��zvGƗE��HE�d<B)`
�'�� �Opx1��JDW�.	�	�'|*�bU�u;z�A�O�8`c�h��']Z�1��X�؎�2�F��)��q�'��a�`�..�̌S`&^�`��'�~�k���n	�E��2��'��8*L�'`���0P4��	�'�`����� lrD�Sܡ�ƌ��'Q�=[�����u)2�!tȣ�'�N���J�~�
\����8��]�	�'�8�tk�m��E���%��y#�'s�AÂ�P	 ��c��E�F��'�nȸ��7d���	�?+(D�p2����Y:�R'� Uc�@;D�����El 8$^�!�4���4D�� `ՊRZj���'ǍHX�3D���V1�&9x�A�
^�vd���,D���ː����M�7�:����'D��� d�;I�Tt��E^E� n%D��h�"�)<��)�*�4@� [V� D�Lb%�=o�T���!V�N,U�>D���1C��HT��FU�,�쉺W�<D����צ	ƴE�wƓ�@��A�k;D���3b�r�8bW�N�)����:D���eO�m��S!.DA�ub�:D��X��']�v�x\ܬh
s�4D��CQ�I�_UdŃGE��D��]H7)2D� B��X�7�,��,����f0D�4�B��b`�\#�퇞U<�E�b1D���rC�6�����Ǎ!��	i �4D���'�ԛi��P�'��$_eN8[��3D���U�%Ii�e*
�ub�	a,3D��r`�pH�x����,e0�qv�+D�@�Q̚�7�D|:Ӂ�9L�� >D��p�U)F�Bv������z�<1����SO�� ��_|p:�v�<	q��i?�����@� �����y�<� B���Z\S�A����$w�<��Eō�5K�d�)5����F�[�<�udV���
��?Fhp롄Ca�<с@P0��)sg���D��j�W]�<9T`]!-���:���[��E
䧜C�<���t<��H!F	���Z�<Q��˯|%P ��S=���&M@�<�U*J.NC
H�J$A&�] ���~�<9W�98��Sn;I.ޥsM�A�<) ,��S��Q����T]�"a~�<� zA$MɝAo������#a@ ������HO?�D�SlY1)X���ů�j�!�K�l�� ׫��K��		0���Ln�����	])WLHKs��<���A�0LO@�DL����=7T~i����J6R��K*-C��Cm��S�*Q)Q�$�����)nE�➠G{J~ʧ䏀Ajպ d�r���4GT�<���ҸS��x���5M��Ń$�UQ�'2axb��J��1��$��c4J��'�yI� ���f�[�X�`�$��M��{�a~��Д�Qb��F S���i��8��=�ia���e|�ߐr�@�BЮޑy�C�I�����q/��;������D&�=a�']����v\��U��WWJ��ȓ0�%b�Ȍ�s�"���I�5!:�EzR�'��`*'�E#5)�ᚢ�R�^�V��
�'��xqac]�Q�b�"��Pb��X	�'�����-W�j�w�K)c>������V; 4�V)EA�|3ԡ����]��P�����Ttlp+��+�N]�ȓ!.0@�biK3P����A�s������X��}�k3�$\]���!8�h���+M�X$���Dj1��!�V�Z��Y�xV�l)�� Tf�ȓ�f�������8d�L�2-���ȓ[mzur0f��k�D�4�H�� �ȓ.�0� �o:;Ș#�̝}$&��ȓ`����w'�`�8���I^�p�p8�ȓ9�F�@�$\��VÆDO�[���ȓ&6�	1m��h^U�g��$H6i��-U��Ѻ�8� ��G$2E꽇�;�`U�d�St�����<-Ph�ȓB��!��e�-�V���J����:�8���J�4�h�:�EM;c|��]�& �1]��1����:|���	~��5M��+E�x�񯇴o����ȓ|P��h7��
_��1�'V&Ld�ȓek��g �j�F���� U�,t��U��em͋\h<�$V'k���a>&*�)����D�8����ȓ!��#6�[�rU��ɢo]�InD��q��K3ē�;�Tz���9쩅�N�I� �tuF�37MZ"=ߨ���L������8u�V<S�
��]6B����Z8v�}T�4���ܞ �Zчȓ�:��sdP% y��D��
z9�ȓy5����iN�?��APa�B�.i��pz�͈��� �B�@Ǔbedq�ȓ wl:`Ƽ{`�M��_�m�2A�ȓ+��W4n�p�j�6����i������D��$x��T0{¼�ȓQK�%�/͏z��t#�EC�"𦁆ȓ��ʦ���g)���P�xj����X�FE�yc�+ÊO,=v���`ƌ+P�úZVԝi�	��U.���ȓ;@�1s��qM�0!��� `�bE���D)��D0hl�P��'�_zDЄȓ]����
�_�}���@�tƂI�ȓe����GƟ r�:dP�*$����.��Qw�M�=h�����'��0��xTTPG!�V}4��ǫ��Z�^�ȓ5 XYٕd�vC^��P�N8Ye���n1�$�ʏh�hTkŭ&��Q�ȓs\��hF��CA�q��c�i�l���S�? h�z��Ivn��;#N;� @��"O�Hj�
U�?Y��x��"d{�X�"O��ysi�$O�hq<=��V"O���AZ��vC�n92�rQ"Of�Q�I;YZ^�A������M��"O�� �O�T�Oϸ�NU��"Oh�+Taׂ_����܃'�ܹ��"O�4�v�^���d���.yl�A�"O�Y��@�^-���K,H]0e0"O��AfAM�dxµ� �̼z�"Oh��/D�
4�i��R�P�*A"OD�y"G&5����,�aq��@@"O� 0�cЖ�Pm�g��*0f.m�"OPaK�V4��-[ֈ�
 � 
�"O�|��Ɔ�w0�����
�D!��"Ol]����H8Ɔ	5��C�'+&,{�]�O�8D�ׇ��L�J1�
�'�\�(�%��~�Na
¬K�=�H�S�'���Ԟ� �Rr�,�B��
�'�����<ղ���)"zp|(
�'4
��G�5���Q�e�&'�E��'XV(!HA�Itٖ܎:���'�����AMp���.1�	Z�'�&���.H; aA%;�nH*�'d@Y����pۈӥ$�5�Ψ"	�'{ ��UM�+P���A2g�.	�A��'�ĄRR�O�$ަ��q�Q�*����'���q�ڤ4�V�p&�W HIZ�'���SD�A���)�:6��b�'ZdqjA�!2@Լ��)��(�	�'y�� C	Bzdl��e��$��$Q	�'�Z���E�8�3���M3�'������3�(���-�{��E8�',�p��le�u���@��س��>D�h��F���tS󤆞SJ:�CS$>D��s��٢]~���'���ZF�SM<D��3t�"��x�k�0�2͊� ��yR�*
��crǜ�yBl���ԧ�y�NP�]:~��4U@����7���y�&��kQ����,�R�Dن,	��yr�ΨP�H���D��tl�u����yR-\2������pd�i*ФW'�y����z �q ]��n�#PKR�y�
 l������'����F��y2�24L��a����� ��M��y򩘱�؉"�#	<�� ���y�NЪ|h��G��h̉ÅHF��yr&S�r4Г3,�.�`��B�D��yb�W)"�~�I�u:�զ�y�5.�.�*CkĆ?֐��e�:�y��f\�TquG��{O�5����yb��	�t�ˏ$A2����V��y �/~.�2�L�2jH�#b��y��9y� q�6hշ,X|Ⓢ�+�y�P�˧eJ�u[Μ� �yr�ѝ=c\��i��C���%kI�y��ԯ���J4=��a�q�y�%�� 8��EKd�1�f��<�y� Y� �ā�*Ǿ1v" �w���yBo_2FzE�F�1`n��Ëĝ�y�/F�Ol��֍W�<Bh`2��ؔ�y��6qc	56@��)W��݇ȓv����� �(3�x���U����ȓ/t�@�Y+"�Ъ&C#n���S�?���� 
     �   Ĵ���	��Z��wID:F�����@}"�ײK*<ac�ʄ��	�$1�Z(x��	��6��"������ �<.���s���(�I���kl����u#Z�u7mƷ?���y���?�G��:��EBJ�S֨�C�MP8s�@����<�t��G�����>at Ҭt�̜#�<iV88�A�^���3�U7�	�'E��OSTغ1���Uq┨Ze�1�-O����Iߺ'SVة�#ӿx�XH�&l�!�l��� %��7x����$!�iP�Y�R%{ӏ�s�D����/�<���NT0|�^�'���CϜ>+���'6\�"���~�aǡh����ԡݙ*���E�5�~�+��ऀTI5}r��8j$��I>y!Et�'G\
���J@�Z�Q|P��V����,���(!E]�I?4-. �� Ɛ=�e���*F�2�AG�NOF���ˆ
��'B����ā��d� ��1���*S�\|�ѯIs�&^2+�0��M>��l7��&�,�SG��Y:Ș���ϑ�t��S�]���P5�|RhW��͘M>Q���w抩lZ-=X�P1`� e����`�����j'*�}�I6+��1���}~��E�\<�����X�l��B ?i�A���,Us�'� �D�����E鐩 �ǝ�?W�%���|�l� bg�4a�-&��A��)q��'>u*��<[J��ߴV���yb���n�:�k���(@rm�'>�p�OB'o!�OHK<3�
�A����J9@�<��fT?��.)�> �<I/�%�,�����U&��JSc\8▉aR�ª^ɴ�iB��[�Sn�[�͏+`*�)1��ޟ�UB�;�qe�I�c�$YP�d�<�1�<Q�'��1BC4H�OP��e��.�f p!�F:r���S���~�&�:!�|��D'\���y���N�ؼ;� Ȩ��0��pX�D�A"ODh�W�  �'~��K @ ��� ����d  ��jHx!H��d\b0"�(G�Y�f��'��Q�!���x�L�q���(�zXqs �2ָ'}�6�7��|�aa�>+���s�D�D�:tk�&?���V�i��'w���U
���U�Iן$���?	�����i*+;�v�
ޮK�4���D���?���0�>]�������Y���W�C�b��ѷ]��U -����Y��b?
U�"b�V�$�f�Ă��)����;��)S(   �  k  1   k+  U4  �:  A  RG  �G   Ĵ���	����Z6)��,p��@UT��C�ֹS�ԡ@#L%~�@�$�.?���D.C�'ll\�02�cm���r�ږ��?H	� f"O������B�,��7�X4J��ي���_��	P�/v�蛪6��[�ΘS�f!��]>^��y���C���8�Eȗ7K����ل)��]s�.ǐm.l��p�)��3�;4����@J�9c*�'��3c�Avj�*Ι'o�L���&��(�r11U��E�n�K�j��b��qk��Z�?����?���$���Oda�j��2����%gS�d�vcӔ:�T0�`@π@]r�s_�jԺaMfݩ�3ғN��5'�@A�)�S�O�3LX��B֜\ z����8��D
��		��TX�N+J�+ `R�th�g�p*��J�6n\ʓҞ��	��M�4�xB�'�"�Oh�`�m�(|+��58�@�տi��ڟ��	���g�,4��G	sZ�K�%?/ݾ�oZ �M�5�i��'����O��L���#bJO�֑+�)X��h���=.����	����I�@�^w5��'�B��u��ٳP��.1� �GX��]SC�Zx�����@LL���!����� É+.Lax�E�H)F}r٪&m�({s�܆�u��e��0`N[ц��B��Q��0?!�������#dU?���mٻg�bPq����M{d6}2�'UR�T?�;�O�[�F9+��؉#�l�ȫ<Q�O,b��Fx���t�V�R ��wⶭ���(�MK��w�Ffu�P�DԦi�P��*�Mk���?���S�Z�p��ȥ����
�*ҦţХ�ן������p�eD'"��M�eF���IJ�,E�x�n��T�D$"�EK�'��:��ӢK�t}��-�
z�F�%D�� ktE�:2^$pT�\xy�]�9u>6P�|�����?!��iK.����k�<iI�i\�/X9�4��* RZ6M�O��Oz�d6���t�ӸHR�����FN���)^X���ݴ6{�i�+nn&!�T��A��I�N�ON�6��թ�i�wyR�'�"�O��5 ��'b��-�)z�(6?�傰(C,4t�6mߦr��ٰE!��L]�݁��Ό�M�O>�S�|Z���p���HcDWgV��R�I��?�EP(4�Ae'0����>@��( BW]>2��o��|
�@�}?@4*�*�<f+�!ӉC��?������W~J~ZK�P0�dg��3������!�'D��G���Il�1�t�0S՚Pr()�?��?����(f"AJ5mR�Nʬ�H���9�M+��?��#	�8�֨����?���?)������G'<�ř��4F D$���MBF����~���&�v���E��s����@�S�IH *D8tk',Ԫ|�R	��I"u��@�����s��c�^>)kQ��
9��'(�xQk ����+��]H�y�.O4<���?y����d2p�0w`�QsAd/Q5&$�С8$�D��@�c1�т��`�2ԪP˳�Mۆ�i>��	Wy����*��r�*֣FXT{d*��~ì�ڵ[�q���'�2�'�j�]�����|20�)mʜ�BT +_<i��A�{+�!�L�Iށ��Ó�9n�� ��D�)���y��˲7��@d��	��F�̬�b���_KR�@��-�&�Gx���?�?!��ϿR�aAJ�=?�$D��/-\����G�'ʙ����g�;\ ��J���<���Պ8!��&g�3��Z1T ��R�x�ܴ�?a-O��*e���'���R�X1�u��d��-h����#��V�K+HR�'�r%��f��FŦOT�T�����8f��yu m��f��$G�h�%�t2�=I���w�| (���	�nI�áʆ5t,ա���t�T�9�*I�(�6�ː��9 J��Fxr �7�?9��˸O��u1�EϺu�j�(�ؐ)ϖ���=�O0q:l�+?XĽ�a����첆�xr�i>�;�O:|넢ҭ>�ܳ���9�$m��]���ޟ��	�ԖOR�t3�'���q���d�C�}7HUBt"S0="D7MY�.����-��ZŌ��G�8�J-�O61��8���%�Nx�5��5�
Q���O0���	�I�I81l])o���D� ���f�	I)���9w���i��|���Q�!zB�'��)�	5}b)9i\dhB�_%v����#���yR�![��B�Z�	��@C�%��')�f&��|*dK��,I*h۴mX�u��L��$��Sě��'���e%�s�'P��'�iݙ�	�$�j\Za�¯OY�Q;�
�"Y(H�F�� ���R��4mD)'v�g�'�uc�	���]�@Q�1I���f���R ����xdT�)�f3���I��(���\"	|����n�6/�0�q����O>�=��'W^����.�`���o��
�'����?*o����*�dK(Y�4dÑ������'`l�V��:�0Џʁ8�LȨ�Gڐ)@m*�'���'jB�h��	� �'A,N�YQ��lRY�Bڪ���u��4���h���8G䙓2�-O�L��E��g��`9���!\{�p:���I@bg� o¬�d�<�p<q0�O��.�Ow%;�`����c#E֦AD{r�	5�`�ÍD�]�|qz���Z�~B�ɥXѲDp��E�ռ졀C� �0�ћF�'h���d����D�?��fg�Th�G��ZKT �A�b�T4�Q*�O��d�O(9��H�)��H#��@���U��r���H!�ьz~�p $]-`l�#�X#�Q�8)�ܗL^�qA��0'@�t�`�T#��Q� ��!�K5x|ڦ@O'cG҉��p�'�����?���4/@�f�I��x\&`P!����d�O����v�%��������]ǉ'2ў�S
��䀋<�	[Q��0�r�PqHܫV��	�R��с޴�?A����	�d!L���O��`4C3>�q!u�K�UDex���%�$�$��`�l���M3
�!��|z��)Aa�X����!�"d���O�9��� 21$�[sL�.6���2fX��S��P����m�?^�SDk�$�x�č )��'rX7��O:�O���OlZ�cC�!A �̠Q��nj9[VR�l�IK�'���I���IƢ�^~�ЀD�Q�b�>A����nӨ���ʦ�O�԰h�D�~8�`��M�TM�J�t���D�O���t��?d���d�O����O�,���?ɦD�*^p�!h�;T� �H�bx�I1�̈́�7j�ԅ�"V�=���[+8�˓{�.��I�=F -� �4/ڰ3�.��T��"0d�O�-���+A%�)#~��9J��� ��C�I#@�A�	R�I�h���ۈ3|f6�Wi���ę|B�V4'U���MR�N�tq F��T)ɴJLg�R�'���'O�������	��`���H �7Ϟ�Ѩ)H�S�.��QK� Zs�`�ҋ�4���D�Tz$I�vJB:lB�X8�O:ot��z���v� B%f �s�:h��Բ�U��ተ�H�d� ��Q�c@�G*����֩)�l�l4�ē�?������4L��M�<ҧ��E끫��V�T"=�/O��<����oAV��T���o~���cͦ-�I��M��i�R�dӐ�$��O �$�OD���1��	9�(A�Q���%� � V�i4hEK1�' ��'Ъ���eۯ���d/i*����n>�Q�![v&���F�@>zmi��)�	|�q"�R�:���%�~)��a�U�*rLh� NM���a'X�V��r��_�'DP����?Y���e���4��1�ܩ	�͂QI���7�Os!�%
�4P'ژLIUH�x��i>���O����
�InB���oT�&. ���^�h����0�	����O�"I#��'�B�\x�0s��ƌT��!����k��7������%�@h��S�+C��.���'��d����S�B��\�w"w9��s`qP�'�Y,�]J��	�R�Ve���V�rb|EF�5(�@ �'[���q� �u��5���4�ؑ���4���ߟ��'��I!7�R=��fQ>�� �J�;1�C��0[��|a��� [����AcՑS�F#=y��S�6�@���B��x&�!�䦝�	ן��Q$	��f\����L�I̟PZw����f��T�f�6�X������I��6-�O�D� <�OB �B�	`ID��#��l����.��?T�Q֡Y<{���ŏ�6��3ʓG��0� ��%���9UM��Ԉ�'�4�+���?��x��'���O����.zR�c�n�3C�I��i�ў�)X��'�2x9�K�
4���L^"
A4t��e���'����i�O��3Dj����ǢD5GgK�+�6Q�a"I4}����?����?a�����O��9J����\F<8�����[�m�m�)H.xa�ϣP{:](��TZ�'����CX	� �B��� �zU[cG��w��I6dL��jh��.�{�H��O%�'�!C1FF�fm��r&ɝ:���3��dӮ�=�����>P|���XW��0�d\�˓�(Of�smK!�*M��K�%��%#�W��:�4�?�*Ov��R��I�d�'���Ւ$d� �MZ����j+ u��&�Fl��'����xi%��<z��S�m�����V%i2FN�e��ҦiƴQ~�=y�-�s���P�P�䴡2�Q	/ļ� �N�$|KD�	��-� �zQ)��D�b4☩%��0�'9����?��T�s����Z������D'�ORp:썽G����B�.��v�'���$���$X�L�p�B����'�&��'̼1�Cw�8���ON�'6������?q���@]z���V(	��R:ݴH�}��D��jO��Ŗ.��x��0j�|hi'��Fܭ`��3
يEm�B>�����t�� (OT�@Ё���#������Oƈ�4�' �6msy�'������Bi��9�fNm�ajc[����H8�P�G���*i\͂�Ċ<86��.�?�����S1N_�q!!
*=^0��׃Y7uO��ܴ�?	�bU��K��G!�?���?���f��N�O>������{~LL�N֙�Y���
v�7M��^se;"��4h�M�[w��):�$j�Q�@�_?$���,�>.ٴH�&k�D� mD�q�X�I��٧
'�Lͧ;Р�{��U�^5V��w�\ݱ�KKs�x�`4�SӘ�a*O�u�1�'/r7-�Ԧ��?I�Ӻ�/F�-�U`��E�a��|ړ��Y�<�,U�WZ�E#��b�L;�|XEz\���'qp��(]�K�d	8@`_E���HDي�'�*���^� M�A�ДJ�z�'�ԕ��ױXhi9w*݌M��}*
��� nTV�\P�A�W�Z� �F�� "O�H�J�6�DH�K��x��"O�m*0�Ȩ!1�e�&���"Ond�S���,$����\�n��dy"O`�[��ܰh�p��֍Y�F�B�!�חO�(ɀq-1L��y���!L6!�Xg����J�Aq.%l�%<B�ɩ
Q�X⣞�r�bPM	"4B�I�>٢��1�A�$U�Q+YrC䉢@K���D��(f4�r@�ʘ�hC�d��j����-n�#m
}g�B��0�<����3%:0�R��*"��C�I�;�|���E�a�Ҡ�ሗ`}~B�	�1���6L�W��#�J�}�
B䉅c�D�Q�V�V��� �1�B�I-X.4���,�!�P��� >\`C�I���3�M�Z ܵ���@�=]�B�ZՒ(�#G]Q���EoZ;;�dC�I�O�rl2��*���!�E�#�2C�)k�$m2EA�� �xqf��}yH���Mچ�$�r
J�7'vؕ�'Uv�06�(K�T�R#�*I˔��ӓmG*@�o��%J�Ũ��!uBzT� �Q�]�����4��eR%�/���2�Aq��%�<$g|]r1�<��,'�]s3��i���>8q�D4ٳ�پ���P�M�	��]Yr"O� y ��Z���Q�)��(�Hh*m�'���AJ8e���`���R�>�sO����/� a.z	j�d�9�ȇȓy+�k5�_$���	��V��؛���v|@F�ɹ`�j���.&O��t$����	�5��\E�'�F��\ȭ(��2�
�X��R7}FFX�F@�;k6%&k
Z�u���ո@�\�G�f�Y#Y(���<Y'Q88?L�H�'K�K�δx d>�� ^-�\�t���kޞ@	��.{�C�ɦS.���=H���X���::�"l;����݁��X�E	H���-*�g~�n�'k!��Z�ҽ��q�S��ynϾ(U��	 DN�����.�v�P�@��E��A�io����*]�X̻�L>4Nԥ@W�O�p�OԤB�}���?Հ���\+t0a�I�C qkP�����r�A:�AV���;@A ����=&R�1C�+gր�<3O�'�ցR�o� �a�(%�S/f^Y�@����zF�� ti�"?���J&�(�ص�BÚ$mp��2fG�o��I:ՀM�k��H��[#�p���H���>�z4:ٹ�i.���AC�C�4�'��qC�>�)�'�l���ꀧ?���;��O N)P���^�++y��ݜc]��
=OF��V��>ѢSLE�@sҭ��>! ���d�%�D "��?��f)����whQ�`�]jDg<�*��ۘܰ>�Q&�q9��6��Q�((dcȲ9{�4�SJ_�@��,��#U�y%���2귟����!B
K�;V̗�EӂQ��C��hO�l����yE��zg�[���
�=c�IS�a[�7���I���%J��/��˧A��A�o�x����	-��0n�)3%��BPn�
gś6�U���L�I_���Q�9������~��ti�|�4�*�K��H^LD
��O�lvH�F��8�؋��L��p<ٶʞ�
��09 �$j�`��M��<�D'���L��F X�)ڲ�|:ܟ��H︘�c��x�p�HW��!�<���#LO@��߰1�Ez���nȶMXe���#�(|鴧���P�dˤ��8Ƅҷ��9I��1���w��8顢ȟwG8mQ�nӞzd�A�R�(c�s�KU�o>q\���;��'L���8cM8 `N>�#��Dጞ���x�l^|�	{�p�`�04�t(��F	fZ*0�s)'N�PAC�B?�V�O�p��N
8�����U��Y�x�L�s�ٶz��j�ڃS[�Ԋ��$��l�c�L�f	�<��I�k��pb��<Y���_�@�~�R�@�fQ
�Ë�~�
��O�K�n��}J���
����]B���9�.)̎��ƪ�[x��;�&	UL���²Ʀ�Y��A�T�dAB��@'~�����%]�%I#Bt�
u�aE��1� ���G	R����xYS%c��u�1<�||8�F-wƕ1aDI	\Rd�=1��i�2���ә,�j��O?e�!��P�݋Gќ{ff�Ydm��	+b|�Dխx0�͸eb��eV����*�p�T܈Kɬ��ZJ>��ї\˦�[�a �,P3T-
?|˱d����F�'c@��Ӈ|�&�X�m�L��5
\=�w�G%ަ�1�ɑ�0vԺ j�1�|U�e�=ShgOPM�� ��E�h���`2h�>�,]�RH X�PE�⥕>FC6a�1��5E� ��Md(�
� �;QK�8PQ��D4�UY!�^(e�(ل퉜j���	�$["�s� �`#�`M�8�����MoFř��"�V��a,?X��`�Y���`!�h]�����O�Ě������aD�	M� ���!��C�{v�d�2O�=�˘�Sh��.<�ϐ%d�D��y��#3D�A��8RD�F�XZ���r�@��R�"���4���* �)��3W��8ahQ`���ʍ�`�j1q�ǽ<A�'W�a���W��YR
���$���8>��k�bʋDo6}1t��*��	�i����WX����H�\�V�EL�dP<O4�R��!L IS��O88f���-�upE+�d͏:�n��è�u����װ>���i.���Ғg a`��B
\^3�]�F]�,z�
6&������!\diҙ����f���6I���P�;oX�É�W�IL|���4���B�x�@��z����q��7PS��(B���=�t��1 �|��x�鉦g4�)P��{*��ڂǈ�>�?��D]��gCݬ9�pgN�7-Oh�y6Oߨ@1h\X�� v͠��@�<�d�����F�:���*��;I#��'jl"��̻,��seH��2:���Ӡ)�f7&D�:$z�H�,]�x�*C䉿bغp���Qw�)�!� N,��(��`��8q�C�R\��2��3�I�a�BQ�*�
~��q�XZ���Y�]�H�'�ͨ|v��'*I._+v�����X���k߿b���'(�BA��I�J��@H�c�����(�H��"w��7J:P���ED@�22�N%YiR��$D�谒͖� ��)ʴ��;�ppRG�<��,˦�n����Q-Y�,e��"8�'g���ԃ�;�n�3L�'>�]�ȓSը�h �Z)+��I�`�\*��;Q���F"���V�'��t�fĝQ�g�I���ɱ$
 (�e�bőf4�B�6D��!�#Z�@T�"U��J?��bG��;B���LJ�`��B�-Mb4 �E�8ܔ� w�1<Ob5�M�x\��s�a�Xi��I� ~�8EC#O�t  �E?D�@s��X�����b���:��0�I �Vpg �C�O/�����ϩH r�q���=��}��'�r)�OCH�j�у�$h$� G���'9�>��#r_���T�*�jx"�i�wTB�:K���a�-{*��Ø�R�C�	�H�j0@�Jc�(9h���/��B䉑X�`a�K�0d�(��� �Ov�C�ɜ2]�G
�� 1� a�8��	�k1$p8
�/Rfш1�،�">G�G�ZFB�2ׂ!2-�Kƍ�~�<ႬQ�NFh�#`�ޫv2������N�e�f�iy�_�W8 �'D�z�JN~����w�Ę�"藀~���ƅ��Z��1��k��A�'��I��#��(�0a��T�4��<�r�1Rn��>@�EJ�Cܣi���%��'��a�<���sd$���P+; �{�k�'  �u���ico����=�����F~�rb�#S
���Q�ݡ1h�`i@�Ǟag&83���$�e�!�ajBO�A�֨̓~6@C��F4���`�:b7&$��T;`hFG�;I֩"r�i�|��ߥ#��EJ�]
6Fq��'+m�-+R^���!��v�~a����6[B0�$�<��i���X�l�%ް��%��,�`��w*�@G��(��*�%bЌ
	�+(ƅ�V��{=ք�`�B�d>���W���gE�.��H��S(Ha~4)ށ�V��f�Z�Ͼ��<A �]�$:%�0�m_*	KOu�'H �Ȗ�W�Dަ�, >U��>
� ���G�?1Kz�����?>1�2È[��t�����L���A�0=��i���3��$nx��AR���<q���
3pI��-De���e�3wi�1��.���CV�ɫO�=��� �^��P�PwzX�S�]�<q�G?A�KFG��-��,�2��򋄁4a�4��jײ=��-r�W��IJ_#y*v,�� �¼����a�T2������uF�d�i���?�'|�NɒG�7xj�R�䔏�8d��¼y��8u��Y#�јcV����&ܻG���Q�茿u2�;�y2
_o��D"T'[��a~B
�̓2�"��'0���#�йq8ry(�*
�Z��o^���#��|� ,�'kEQ��m��e��R��1ʃ Ҳ82V%��˶Z�9F�0�5YR&^�~�v�ᐤ��f�(I�@�e�b���n�.	*�i`��$_;�5XP"V���
����;2�D̉׬�4TŠt� Ō�ȌG2/N�^RP��!�q��!7�\ Q�\�	&˙�t�z����t���(��Ū r�I�����A��O���DG�%}��r�e�=�b�X�w@��xtL�1u�H��k+��R�O��1� P�'͆YY��*`�V=8�����ҚNo�����Hڴ��B��i���Z�P���WBS�\Ȏ�тCA�ZPA-��>e1O���R���VI���WrY��)H�h�x�be��y�(��(]��T��'���O��E��_p$Лs��Jy��p6���юE�O�y7�آ��H,'�*F|R*ʑ�yG��.��2$�ͱ�NqB��ͻ����#;c�\��O�d���|:�>qt���EF��Fdʰ�t1���o10�����BlڐA!t0�īAa@q��PA՗E��X��C��  "��U��OT|[���=�T�(*}�`k����X�:*p7��j�? ����=ۆL �
Y�d��,[�7O��ӷe�$P)�dKbfݒ����\�擩���XϏ�-lL�*� 98��jg BsX�X�'��eY���rf��������"�W���'H��7��+RQ|t*�d�/\�*��		0��� )O�q�C�G�@�$��OQ��s�ғ}�TqB�Y�AAZ]*�z7(<��G�`4���$X���
Z��9��y@� �T�ުS����!ń#a�hOv�}�	)�~x`f�.yPb=�茤e^�,ʊ�䗠G��-ƣ+ �IX�܂l]r�ڶ���{�F�y�*Ƀ�W;�?�tC�7���I�\ȉ'�T�q!k]� 9��h��H�-~]��j
q3,�a�/��('�� �S���e�<i�D;�g(]?��h1�r���]s���w^	�q�����@M�IFo^+���&�KBg�O�����	�]���L8��(�J�����^�F�[�Ȑ �P�`ġ�()iz`���%�8&�ʉ�������BD����[�(�:�
���i �iR��P�;��R�-�O����o�)�RC�
q��t*��~���"���I���-���ɢ���c?�i����FK;:pNuhV���XfF�x�Ѓw�S�r���z��s��pi���n< ���'e�jh�yjHb���}Q���&��$���M��zD���g�S���a���@� Z%K̻r�����|≸7euϓ9��Q��,�4�'0��X�&#�+f�r(�4���6c�}�D<r�y-���O:PqH�K��I�\�<̡&��8��(�r!��*60l�ȕ���e�Rp� �@�`O<�U>$ ����^92Up�`B:.���@`Ⱦ}��(f<�i2������h�ma A�f�C�f#�y�*�?B�� �㒗� �AG �?!L�8p��x�T�[�� #�&����wy�T�0~l��e��T���+�*�q�Bk�fh<�񣋿>r驱F�P�ؐ�!W�Y�:���/��z�T��a�]?����&_9t�Y�H���Д�g��y4M�d��X�O���1�#�O���3��S����gCW�3W&��� k0}b�T��~"c �n�6�r1�S%qOI��eE�r��q�Γ�kh�,��퉊a�}X�0t����
�K�6�O�rl�bEYtr�y�i\�*��� ڴ۬)��FP�4��דX'ʱB���U>�ge�l�z��	;t�L�[7�� <�V0ˢ��xgJ7]?�-=@�8]c����uK
3O�6��� 
��	�'*�a���M�F��fm�]$r,���ɒ[}T�@�ӡ�H��fj��1;�	1@F5�B�	%�$�JD�.n����&4z7-� �@�"~n6s�"��6?V$�3�C/o��C䉥V��H%(�/uB���nB9|�B䉔U�\`Qe�9D�����}Q�C�I�Q+v!��
�J����N6.B�I�u6���
�rӺ ���M4uVB�'AXxC �U I��ȡ�'J�'�ZC��>�v�SW��1��-˴�V�h;,C�I[;��� "kl���ҫ�8cdVC�9!��;��7q趵��^_��B䉘�2E��\3�Q�7޼g�(B�	�B<�g�²����q��C�I�J��T ��3��	"�*`B��4��l#��\�1o���RGK!zbB䉖V�!�f��#���C%�@�XB�IDʔ��������ڴ�W�w8B䉃'����&V������Ј\�$B��8I���@�.H��ѐ4j(1HB�F�5�Ϗ�k���G�5!)�B�ɑ&l��R���t�v�A���B�	lBB|�c������ϊt��B�	5E���h͏Q�)ㄯ�8��C�&60��n�d�\���@W�Z(�B��j�F��!�]�g�pe!�iR�0�LC�ɊQCn4Q�	�/40`!�d�˕t���䐖 �0:3�Q�>��c�i�!�D�<AP(t��Ȍj��H�	��C�!����x�R�B�v뜝:VH��!�dm�L[��kI�Q錈]�!�dۢ[��raӋ_L�\� 6|�!�D��V���@0iЮ:J���� V�Z�!��ێ9Ӯ��Gk�A������Py�0��%y�J,bV�%�t���yb�
�e�.L� B����环�y�+���,sjP�钬 ���y
� ��f� -7��C��_�K��T���'����R�s������C�p�{ro�=Or�C䉵����F�/zt���)��` B��')6H��j��$Re�m��B�ɣ~�iU�^�'D�j�(�1;�xB�I�S��yR#J\5[���1&J�HB�B�	�+�h�R)L�0iy  �-#�!�d��f�	H�5y����N�$5u!��lc�O�t��k"́�~t!�� �"�Ū{VB�zSA�>U!��6 ��t�B�Ll�C`΁�!򄕵1^�]�A�7wӬ�)�΅2p1!�$��U�j����-!��i�.̌d*!�D7VOZ�Z&ڷA�<�CF�N%k�!�d�dd<cą�<p���;��Jv!���I�h�e�'��UID�ڢ.\!��%r2�h`aY�-�
!�i� +!��06y�aƂ;�XQpǗ6!��[Q�J�`�炜C�(,[��1 �!���>a��ctFQ<I�1c�Z'i�!�$�(]�P��%m�$�ħ��5=!�$qe����ˬh�UbDR�v*!��N	��D����J�VXz��ժ�!�$�d�t��I�9C6�)C�v!��4�>Q�d	d@BୄY.d0�ȓ!:�������4u��HW7��цȓqNm�S�]?�L1rd��1r->0�ȓ+��j��� '��i��.0V�ć�`���5�5�c�Oq�^��ȓyj$ꦪ��D?�ܲFg%q��y�ȓAB rU��5��Hg JE0��ȓW�Ru0��
T	���ef[�<�Ňȓ=�VyZsR9dp�ͩB��9��ć�?ٺ�Ka� G�����ӫ�����"AHp�Æ�+Źw�?�zчȓ@c�!�#I� �Y �ăԾE��to.�SA�Hv���T �8��r.��A!��S�P�Uȍ�^:���ȓ���KCb�2�r�ed�����,D�T�����a�\�Z�AE�}5�Pc0�-D���PΌi��� VO��M.��7D�̚p 4C\U���2��)r!D��K��jf��Ã\�lO�A�>D����1&
��h[�8,,	�#�<D��Y��a4h�Q1 L,V���Q6(:D�+&S�~T��{G�1>�Ȩ1�a7D���eo��s�صP��ݿc����5g*D�y�n�.f[��o��?��8۱�(D�`˔gǆ{�V����vO�|��'D� {Q{x�<�p��jЊ'D�da��c4 LJ �ɏn%hH�)D�$Rb �B�~�#��D��r�'%D�P� նy\�`�却o\�87D��;�@�M���5��*cdPh1�H6D���� �b�vxF�n�F�#�!D�X -�3���Z�����2lXCO D���$$`��VS-X�& �m?D�yB�!c~��nL�� B2�2D� C��b� 8���O�L�
��R -D� �Qi�5	���qĂ�ap0x�7�?D� Qb��	�u! +ۏA?��<Q�fD�C�~MI#lK��z�Q(�e�<���]�L8
1�1K�zw�ψF�<��#\�ul���SnP�`������i�<� �)�$z�6,� �_�>Ճ"O�U�M�j-n̪����p��,��"O����G��%��	߮�2�ء"O����e��@z踔�N:i`("O4�FaQl�AN�5"e�y�"OJ9�q�W�J���@h�����"O&����E�GYxa�({�Fm��OnX����ed�,KԻ�9n>�	��L��p>B�>iBƟ-�%���~�#BNA\�<��bpi�@�������Z��MSD��t�Ş;����Q��\��q����_�����>��q�п{JD����,4���D{��'�n2ǂD)F���a
ߑ����
�'+� ΏSy M���S8�<���x�4"+���qN�[��t�k���=�fK�U����T��Cv��9D&��tA�@B�	,�č�Ӭ��?tf�xCS�Q�^⟀�ݴ�0|r@���4�l�&!�u���'�p�<���(�F`�Ć��x� �Qt�ğ�F{���7� �CD�nx>M*CP��NB� ci���șd��0g

#5t�7- ���3Ț�"��尲�M�S9j<@�
=D�H��g˜m��a�żGBL��Cn9D���&�Ղ���UMv!0t"S`$��hO�Ӣ�l��O�\�Թ¢B���C䉮

xZcBה���i'啼��C�	zS���⤏�K���XA�|�"O��@�ǅ�^y��'�6�R�"OTaSb�Ы�Q���c���"O�5���@�A�A ����ƴ��"Od�[�(��C�NUP�
Uq��b"O��2e��
H�P�j�O�v��$"OD9���X+�(�Ύ!<v*p��"O�d�� ΢<�
�0�-M���"O(�qUh��v����L �8��!�$"O�4��A�T`���|���b�"O�$�섌_��{�j�-nĴ�!"OluCOH]ǰ	�©ϕC�؁�1"O>��u���3����Ũ��Y����d"Od�ڧZ�3�^P�4�ͫ]���E"O���C�9j�n�+� s:|��"O:h
��\"�%{6.�$jz��K�<��Kʏ1���x��E�3#t$K�Gp�<�2��Y�!�P�s�\���k�<A�\$bU.��N˧eε�&��~�<�w�K�iZ�̇�1G��@U�Pq�<�EiM�-)VQ ���<����!Yo�<)��Q�| 1"e�A��mh5��r�<��$K>o��`v�92�N�Q���k�<i��""1��r+��*��]Q��j�<A �8N�<�I� ��'`�M��h�<W�O�C:�)���6a�U�TK�<�VA�)�2���7i񦜂%�QG�<��E�/Z�mရ�@�.�r��i�<�eNI:&���C:U�j�ȗ_�<�ǁ�T"b���;�&�Q�@�]�<��:.)vȱ�$\2]1*,�sX�<1E_@`��CUa�+y%�Q�d�Q�<�Γ*9�L4��.F��!q��N�<YJ�#n
� +��N9��AŬ�d�<��Ř�'����T��y���F�<QRl��X���E�Q��;��UZ�<іj�?s�q��jV�;�ժ���Y�<A�	�3|����dЎd�\��c�T�<� b�����kg��#�/4��)�"O��х�FJ���f"1�C�"O2!8���8a�=����)O-���U"O�0a���}c�p ���.~P��Q"O�e�Mزj<������<�H�"O��P��2R�v�" �/T��C�"OBt� �"8L���`�K����"O�<Q�W�!��X�`��C��P0�"O��hbQ���U˰n�*_7P)��"O��chW3o{�U�M��)>���"O�%��Cj���{�았v�P�	�"OXX9� �5զ!���j��̃'"Oh%k��U�G|>��wgZ�!�@��"Oʐ22	�TN�}q�ůlĦ�'"O4H�T�ZT(�Z���+w�tdq�"O��ZîϮhl�[�U�bT�P�7"O���+č	�5���Z_�X""O4���qXaq�e[���`"Of��aN!��ɠa�J-|1fY,�y��O���&�R�x���a�@$�y"U�9����dS==��1���y2���$�%l�4a9�Ł��y��;����cxPɷ��y�cWFш݉� ��RJ9Ѧ���yR����7	�1b���ѡ�#�y�ŗ��Ji�%[U�dDȗ`�,�yB	��|���UW�`����yr"\�D #4��-�#E��y��4i��Ҳ��-2ȻC�9�ybd�:eDPP�� 1�r(��yb++�tS�� 
��ę��y�@[�~�x�I�N^ ��`G��y�k�=*[�� �EK���RGӃ�y�Q�l�tA��+·6�K�� �y�mW�1�̴����$�l�� 	���ybj���p8��/Y����	��y�_v�������d9*���y�"�fİ���@	�d5@qW���ybo�Wb�Q$/J>+&-�Q�S��yb睒f����	��Q���	t��W�<	�e�,��%B��٢`Ɗ�U$^i�<Ĥ�
�@HÅ�,��-�g�<��ہ�Vu�����ܤ�y�GE��r�� o�+lX��G�J�y�)5i:q��cxZ��z牞(�y���:;��yu%�u<L00"���y����̮d���Q�6}&t��Z�yR�֖,ƒ� @�2��5{���y2Ȑ~����]9VH)�!���y"(Z�Y6Z	rT�RF�K����yr*U�WFʡ� ��!C������y�g��KV�ʞ5~��Q��y�J]6�9���S4��U��N�'�y+��Aab�8ӌ�'7�D�`PC�yb��2v��A�J��9�aҶ�>�yb��KHb�0���P�cߺ�yjI!���wC@�	[2�!E�1�Py2����a�̜?@�i8V�K�<�N�m[n�c�͞���f�TF�<1��C5Z���f�F���#�Om�<QE�84���+�P4& x����D�<i ���1M�Vڄ��P+��y2NE�l�E�U�^��� e9�y"�Z�	��hf?X�ŰC'�"�y
�  ��&� 4`�B�ȬX�Da��"O|�p3�M@��K�:`�4"O��x��27e�̀&/��dL)+W"O�e�,B�RH�w�J�Tn�p�"O>���cW�$k��%��$l( �q"O�u�S�  �      Ĵ���	��Z�"wi��:G�����@}"�ײK*<ac�ʄ��	ڤ<�Z(x�*�	
�6͞~��#t��iR8] �H��_�P��G�9C�A�6E�ߦ]�1B��uW��#X�"Mo$-�D���ԟL� D5�q�ʘ�F�V�SFAf���P�@�`�Z�3Ѩ�N�\+�>��\���A����\�=�H�ۓ��8oj�	(u�ђQ
�.���G����O�}����'�𽢴�A�f����K�O}��KS@;lgСd�xRB�b��\bw���JIy��� ��8��R¤C-\:ެ��	����.�a��8�K�(�*��@&�y�c��v6h��6��M��C��~�3S��{�*}RGS��c�B;}b�PR4��FH�4��펾! �%E"��@a�#~z�� ��u��2O���`	Z�n�PG=Q)�$P�4���M�ؠ�^a?d��K��O� �L̪�'(5R�*��iNe�U�gD�����	Vܑ��� XT�/���Y֊��@��L�"Lie��ntfX�EU�[�IV�^�l���Z��y: 8 e�.��IJ�h���뒍��� #�ת�xED��#K���'A\�6����D+zAJ7I�����S'5��Mɔ
B�#N�9�F��<q�e�O�D��O�D�����|��C�l��mb��F
B^$E-��`��ڦ����ēd�dA umT���'X�\R�ʙ.~��6/Y�
���Ahh��
DE��OblE�oY���'?��$�4	B@D�v�pB��Ԅl����e��HG�$	Q�؊�'(\��kC".�%u$T*Btp��5@	94':�`���MWh��W?�������
�:�J� >�̤����@�������T�>5;%U�$�2�.N`��L�pA�	T����O�`2��6~`�x�HM(�Z����hl�,+���G�Ě�c:hl���U�	�s@���wʨ�F�B���q�Xc4!�,J� �  �QȂ��4H��8������%"Ol�zG�0*9ȓ�HK�"}��C"O�Ĳv��]m�	� ]"Ox�Sdmt,�m��؍&��"OlH�����$сJ�O��˳"OPcˇ�&tH�����DY��"OrX�A�^<86еc�ʋ3jF`#6"O����� ejԩ���:4@���"OJdn?���S�!]'��"��)D�Ѓ�S�4�[v��;���$   �    u   �,  �3   :  h@  �E   Ĵ���	����Z6)Ò�,p��@UT��CnѶS�ԡ@#L%~�@�$�.?���D.C�'ll\�02�Z���E��_���QVI�	rh0t"O�1*���>�nu4��4B�#�!'dꠒC�ԳI�� ѡK$:*�I҂$!/�$�;�
�)Ҕb �/;\
�)?
��<X�cU%���a'Oo�Z!�(��3/~�PI�\���W,ѯ*�@H�BQ)�����ɋt�����X�9]X���o�K�6�$"6�x}#"�Sh iY���?���?���G���O����6
�$��e��OF��'� ���j�o��?�H��@�LR�4�;�Fz���<mw�MI���80,|�oŹ�(�W'�-xr�G�~b�Ʈ��(�CQ���GOZQ�N)h���Sf�)wE ���ۡ<�O����%�I<a���?��'��0�GO�)��B X<a����4��D�O��D�E�3�I,%���Qp��+.����#�U�t!�7M����ܴ���2����dXndJ�㲆�37���'�3w�S��f2���O��$�O@I���?�����d���e�f4���ēX��$�SdňN"�Yc5�>�����D��M{��)��@).e�b=[���ꐢŖ !�����6V^ "6/�='ZDmZ*V1 |�GT�61��I����؎�b	L�{*��Qi�]�2���&�:.��7MNŦe�?QS�sӘ͛�
28�2������Q�^��y�� @�(�����q;�0h�‿����<+O��:��I}�'���%mNj�k�ː<��� ��X���o�z\��'s�Z<p����&c��_]��:&�Hݦ�S*�)��^�L���N�HAD�=�c��:s�4����N1��}�sa\�!ۆ*7e��"&8à#� x�b��'e�55v���$Ϲ7U
��''l����?�����ï�J� 3�_�h���RG*����'�Oxm���H�5�I� ��	 �J��'���%�t�#&?��l�"��>��' �'���'W�{%^5���h�D#��i��B��x0b��'K:�M�4�d'$Q`	'���J�i��SY��>��Q0�㙟\_��#U�H�:`�鉴��O>EhfC�#BzD���׆HiJQ���e_B"UF@NU��7��IS�LS�*�`q`�*JL����)�O�]�?��������>I�eM�&ȸ��pɏ0�.��O^�<C�мo pp�ԡT�'V��:�X]�':#24��
*M"���a��x��w�_��v�'�Ҁï[�����']��'��h���I�&r��F�щ���􍙗?���QT'��_�ڝ(���~����pm ���4n|���<~�ƙ������iA2�J�x@&�kW_� �&̰��|2�	Q=FHfئO�y(�Lβ�,�Qs�)p�p��Z�t��'���Ij?�m��H�4qq��E�aF��jH<)�"�a���� I/E�D��5�:|��c ��|�������6"X�I�|��* �5j'(ϤQ.����O��$�O���;�?�����M�=�xpu�?q_fI&_�c����n�	 �C��P �C���.f2���'�ݕk�eX��C"���,�T��e$��&:�Q��2A�VC�Hc4"<R��ʟ��c��u���# �Y�B�����M���D:��6�A�蜣b}.,��;^�i��Ix�'~����?����G�Hn���(�O�o��P�'������~�����$�S0̒)���
 ~�H���M+7���?���?A��:F����%:-n>��H��)�X2��2!&J�Yͺ%[k�Aўx�[���CK�(^���K���hab�a������`�J��t��Q�8'�@#<9ׄ��4��YܧW+�ޣQ��pQ�Δ�k���[��>���)���b�iD%E��l��Oڝdٜ�'�`E{�O-�|� ��,N�[@Pɀ�䄗^]���'�֐R`�'&�'(��/������)�N�}^R�*ua�~�2��֚�M;�*F7k��쫢�Eq���Z��#4���N�'}0�)��յNB�Ѳ��!3́�2t����'�KƘC@��aBf�0��ٵt`��|�n��j��@Q���Xl�lȂ)��?�6�ݟp�IJ~J~�H����h��$+�fT�*�T�a6D��A7'��z��[���S96U�
0��ϟX���4��$x�	-T��mA�&��	�����	ޟ��2�R�Wp ��I����	̟TB[w���iT�별G9F��S <!�H��e	'K�1��%MI#�|Fy"G�X^`��	�~�29�!b�)c$E�f�	�V�,��(W�*JLS-�Q� �bf�$��)$
�B��b�<�3�OT�� ��~bL�,yH�����6bwV�jʕ%�y���CvR��v�Ia �bCF;�M���i>��IEy��C�E="�&G� N:0��	a���v'ӿDyr�'�2�'#��ڟ����|�h���H�H[.�݋��ѤT�|��t똋�(��&��.hU�����YG�8�e��Y��yʴ��XH8)aF�Z��笖�\����Ǔ�K�N� �BQ �!<�u�N�sט�mZ@�'Q�(����E������5Kf����.D��C�b�8;襰���\��5���>	��i��X�@��E�9��I�O��S6U���4�*/�����ǅ-��6-�E�^���O>��=̬1+XD
��Y�Y�2/��(Ҡ��A@�@S���!zL�+���6(�a��ɍG\�2�A8.�	Z�P-f* `���m�? �|h�C�;�K2��]8��]�'�V�a��?Y��M���D��?rt|ks+B�����O���܂}�n@z�+֕ٮ�q T���'ў�S���D��>|*@f�˃5���j��4;��I<{j>�!�4�?������,T�B���O:�9��M�S�y��̖�!�`��C���1��(5W0���M�5mٶ���|����F���!���s�_�`�@v$�O�P�״wڀ���
�S!r���!bZE�0�6�&e�eE�C�ThˀD!>�l�$�[;B�'.>6-�OR�O�2��O��i��MWh^�����"J�$���Q�$�	B�'���Kn���K	�l4��ɻX���>Q�{���EdӨ�ĎĦ	�O�x�hs*��t��-㴢
0$dx]�� u����O@,xb�Z2|����O���O�����?��n�"o8��A�
�?�$)� �َ:剻;�6������曙A0��Ag�%hyr/O�}�!�'n��K��_$�1�� 2[G��.O��S��'@J��d"6�܂LW� 3���E�!��F����%�N4�
��h�%���/.��|�M>�`͒��IP��Z4Q�̺��X�Zd��,��?y��?�+U��O�d�Ob]3�FGoQ��WKX�`5�q��Y�t(BSq�n�iU�T@��x�(B�t=}��Cˠ')!#�N/]�|9����6qv�{�&���x��3��ڌ���T�bg��i�^�d��8���@�EY�,�47-TF�I֟��Im��|�����`� M�g%��EC�+�����'�Q��ʠOΘg�<��qc��L�B� g�����¦��ܴ�?1��i�h���'{��'�ZcΠ\q�@Z��;D��w��i�ݴ9c@M����?��E�B����٬��D�\�*�<�28P��K4%ER�����v��XE{b���`b�+1"��|�b�S�$2�Q�Ǖ-��j�DQIi.��M�7`;�����6bX��'�q�,`��G�FT�Dr!eD��̪VR�,��Iy�"���c�a	ʌ� Qs5 O�=ͧyw�	=fGn%0�mK2W�@��#�>I� �	�������?	����i��0�Z���ON�2Չ�IP$�q�� �w�����Cަ��ӏľ ����X(4U|����ɠ|��O.�³*L&�X$C�:n��U�T�'���#JH�"���5�Pwc�l�:��$�#~��џO�-څ�R*0�d�2!�J��)S�'�.�:��?1�O�O���4�1�X�E6X�`&CK�!��ȇȓo8�X5�͞2B��I��.�Gz�N �$�KM�L��e���^U
5i�i��'��p�(= ]�'���'����'��&BG
����K�_F"u[��W	k�ȓ�+'T`����^?#9��'�O�<C�� h���S�'Q�{u�ٛ���3t�����b$��7��.Y���'@�X8W3}R� ���u�۱Nd�!`���!n��'TўH��<�z�jtN]"'����ھ}���ē�Ȕ���֋$��*�0�!B�ʟ�M[!�i>!�	Ty"Gם^�<�zӭP/�N(" $B=��a����51���'	�'��ם��T�	ڟ���Ð�U���A�}�r��sa�	n�y�����>�$��5|d���
��������do6��U�Q
(���D�GU"F�p:BɻG��(�p� ԃ��@�6MUæe�	��<��ן��	꟔�O��A����b�N0,x��.�v�6��Oޣ=����G'��0*6�H5i]Lis�Je-���'$�6m�O���0���@%I�l�BEm��m��6�,<��I\�	Q`�[f�Q$:C�	�  ���r	��A�&��Z5e�C䉁$�����#�77^�I�k)A��C�I��܅���>Aq�)b�( �_��C�	�>,�i�V��$@�=3��M�C�	Dm\���ѮB��)�G%ՄvK�C�I�1[N�A�Q&�ʹ�a-H�6*B�I�V$����ޔva��w��`�B��f`�P*���^�Z�Y�MՄ_��B�I�K֐S�b� O�p�b��-^(C�	�<.�y3ňl�&LSF3C�	;bI��a�퓻y.��ra� ɨC�� <�r�[V�	rv^<��l��x�XB�	�/v6�o֍"+(("GDɉh<B��t�(!Ӕ�θ9wT�7��
B�I=V\2�`�G&�·Z$4�B䉩G�`@���X��p;%*ƅ?NVC�ɜ0��xk�@	�֜:P���
?�C�Ɂ-��Lڐ!�"Ӽ�A�ŇG��C�Ɂ=>(:�Ǥ&�ܤSƇ�<�<B�)� j��̹F7�t��1�9Q"O�����H2V� ���A�\��5�'��� �߰���0H�74����'� ����*����H(<�Ŏ�zz���s�	2%0iCb�`�e�iB`�0lx<��c��'��>e���I���iB%:r�a��>D���L :	��P𧒇c&:d��N٘apN��H�/E?�y9d�C\�#|�'�N����P�%�1*�h����'����w#�#�e�h��{Pf��^w�8��N6
6�a^q8��%c˲b�40��[�Ei��b�3LO��x��ٲ+a3�!Y�
qr�	3^�ީXF�2"`����  �Pxb$���H���
+S�-s���?Ƙ'F-r���/f�����4�~��}�慚�;d���I���`Ʌ|�<�g��j
�SV��_p�qh2Ł']�ڝ��(�%�������|�'m���Ү5ɖD�	V>LP��'�
�{ՆK�����r��ȭw-8Th���AN0is�'�K8���������Qmؙy�$�­>LOl��2�Č���R�ܾfļ�lL��fd�e�1R%l�S@��0?)\�M���\I@���#�	$P�WY\�<�$Q�S	I<�̄�@	D?(���>Q���7T$L(b	X	7� �e�*�g^@QG��
^5�� ���NLMP�፰,�TA�G2}���R���$eY^	���آ�CG%.��|��u�<��`�>������H��@Pm��zy��C�C��@U�\�E��L�4�2���p<�&�G�U*�8BC�Bj�h���w�ɥPTT�ҏy���U��/�~��#�)M��*b��%;����g�1;�B��d�2�5�wV�5q�
�� ,ͨd@�f�Y'�̩fD�&r�XycMM3'*@ٸ����YJ�Ip�原��jk�#.%Q�蘡L�$7���?�K��ٟP��\H����?�(E[�Z�Z���D����G)Ҳ�ӥT*J8�3?��D׽EyN(R��A�h{�|:�oC���Y��eŉJ<�|�p�Ϧ0ݞ7- �ov�Y*�+��sh���]͂��d/��">}8�N��1|���Eb�A���AKr��	uCQ��m�'��Y��m]ȟ��"f�q\ D�^wVd}��[
"��'��S0-ݍ2��H7�O�w� ]	P�a�����U�D@A��X�����Nƺ��$�f.�	���;���`��h��Hb�9}��0��w\ȉ03�Q�ll:����^aKF-��"dو%3��en�Y>1���ޕ) �Y� 4"#^UX���z��OF������|�6xKa�B�x2�Z_H���a%D"
�P�@� c���,�[�B%�,O��(BG�+����f��uP�D�nd��cZ���k��N'%�0�B.Op�T��Ƀ>��P�Z2"\T	�Pn����7�W=�*\H@��a�J��U.��g��tҍ�T*��G�k��D�@�/�v��&$	�-�y��	�6���",�mgkA'2T��4���N���G�=��4p G</Î���+.H����CӺS�àf:`���2<�v���̙��Ů��*h.l9�m�e�X|2ghܓ �>����6��TCwiہ���}��2P�Ŕ:`��ʫ5]����c�L��N?l�.�[ѥݮ@��02R�ݤZ������қU݉'���K�O38t��QSo��R|v�T�H�k�5�G��<uu�d��J�
G#4j�RUc��2���V�O^� [Ώ8A��I穖+w�������U`��Pa��1j�p��'l����R�@�@,9f�ߝih�Ɔ�0ZH.�ܢCfxݘ��N�
�x���)O���/֏Q��l�5�.��i��r��y��� *Ú���d��&	�瞁C�.$hu,�y ��n���e����8�ͬЈ�Q]waˊ�Z�t(�Y����b����b_�a���qD;
б���EM�4,�|aU+F�=1�`��7�N�t;�$�!' >:/��ˢ
��pl�PX�:2���¬�q�e�Ɵ$�'+Z� �Ȥ��@�I]p�*DcK:����\k5������ӥ[�D�S||���K��6�=��B�����8@���F"U�wd��5�
$>N����).�RDyߓ�Ĉ�%Yv�r����|��5�I�ڒtbQDX;��ɱ�F�z�ŉO~ʳ�N�|Jp��L����e	}�z�	b���T��X$��犄F9�J�N^�v�؝{��ɘ	��Hk�O��(d�h��ŉw���b�d��So�85��AÝiu�ɋ$�ف6� x�"�|�'�����ƚT�'X`踲�]�Y�H!���	^�P=���E C�\����>O`���œ:�^0�E�9�"=y��ҏ!T��-@.8i������F-A��?($ �/B�T��q��3/�Y�դ^.p?̍"�L_�/6j�Ye��y��� ���RK���D�3rp��U�T�PZp��`�$&��Ir�i�s��S�3ɔ,�x�"�-�6\�� 2��?m*劏%ɦDK5-I9��s
4D� i���h\>�QժC"�vA����V�����S?-�%��f^n k獱|�K�}�x�3�w4��K'X�]�ȣ�`Tn�z��Ot,�Ja/D��a�Ӣ�{dL�b 	t��T�r)���O�$i���Cc#\5hb`���	�6ۢ1Ȱ%j��;�@�$H*��?��Y�M��խG���E�>d8�m�bj�0�0���� 8���b֗j&V0g�h���)� $9��D6~�h��@c��	�U��P����c��@�+X&)N`!�Œ?e��i;��e�'0�.H+��D�t�\�qJ��g�݅�P��Ep��B�uwd)��{N�s�F4w\��XsO�2a+�l����;w�D�OJ��¶�Ʒso�.��<����u���V��z&�K�8ɡ�DV>2�Q�L��j��L{!b��"����-O�4�7啨I�9���7T(Q��I�*�4��[�1O\SD�m<��K�q�\WL�0F�<u�)9	L��81DC�#8�1I砀 -�Ԑ���I�S�4�;� ��%^� ���'��� �W��U	����U��<�OAΌò��>n�`w�]�Z���'�(���\�2��(e��]K���	�"Z��	�2�9۱<O>1Y�5�\i���e\�9��۲9�P��S"O��B���x�ar䚘z,����
L~(r����K7���Q�9��ƫF=�y�ejJrӈI ��*D�\���0b}aW�V�/5����o��	Q�q�"h��ոɺ��֍:v���&�5x� ^7z׈����2��0�ȓUK�5+$CK�N��@�J_v�h[��V�br4E|ҍ	H���
��ywl�&l�P;��H(A��-В�T&�0?Ig.�C۶a����'2�j��"�)%�\� �ȗk�Jx#�T�(�.�)�]IR�)�ND��<��
�mRSG6XV�]�b	2F�#>YCD��m*J���ҀK���C���<&����Q�5I��nA�s�
@��m2���iA��T��x��K�"df�@.�|IQ��e�(Cd�I�/�r r&ď$u��y��O�O�D&0G|HS�̕��M3�B�cǆ�@u���H�*E!�E�<ad�=q\���էU��a1�.&�ܠk��|Y�-
6��c`�:1�����o�D@�n�3�yW�C�������0aO��I��P��0?�`�ת_B\��!ʕGT������.p@�
�(Y"\x�E]\J܈SR��!G����-ҥ'�Դ¡̅h�$�m2��S���.�4���D|� ٱ-�vu	��=7Z�`
w����P �c�Ș)(�bT%��:Q���6	�8���=�0=���ܡiy�,*�a�v� ��<���Ғ�j0pbO?�ͺ��đ	��-(�3!gv�Ѽ����!��"Lʑ3%�6A�pH� �Y�<1�E-9LV�#��X�W����O$3��Б�h�	"K%y�ꈾ\�A3�My�V�"��@�7-����C Լ+W/F�L}�`$-�O�)!�C�e���ҧ�J�����*=,�q0NU���Rgˡz0������!`�S�#k����	]�lp6	6扟[{�0�b�G�	�L�	ǉ"_bc�p ƍطx>����)~E�q0�*7|���ξh&xI�".ƦkH,�Õ�?^f�d���ibbm��̒���	����I��^Iv�BqNՎ�J��A���_@��h�94���ig�\�|���H�	�>�v�S+�Z��:�@�P�`Oք� ��s��=
3�I8��<[���0���x� �P��A& r$���ŇZ�$|�!eƽ8�e�-_2o�^}��N�<�܊��Q@�r%���ͷ:n�}�'iލX��N�>Z��a����)X<)B�O�b7�Ɏ*��a� �a`��R��6h��O��(pO�d���Y�W1M���Pg��.Z_�X��O
i�(�*�v���R��%c��AO�m̓\�ܭ�����48�x��)A�bXȡ�͚/)��I��'Ϊ��#��|�\�����>qR�0q�ɖ�Nl�	�&ƺ��4��.ş�l���Ί�X�b��$�\#�Q����wƨ)���^��!��<j�zg��2X�~���a�N}R��C�b?��w� �7��	U�|A���6+��()E�	�"r�98��h�<��b4e%�I�����C��8"-��##n�<$��6ƓS���A�[$�,�O�c1�@;F6H�X4})2�)&>��U�6?���H��(��	�5�`����DHA�f!	f�>��|"!��$$u�6�� wI�Kv	�&2���b���	���*h�F8�&Y0I.`�B���o�r��� 	gEf�3.V�q����#�`K�ɘq�PC���@h1�i�?�"B�A&x�Ą��MȘ@xsׄPbe��D\�{X���s,�/n�̻/���p���:i�PD!4%�:k(L���_;�̬�H<���iڧ>�ڝ��)O)#��Sp�9(���an#��4�+�i�6�<11r��lΓ�ΰK��K�6 rW� �0T�=�	�d���h���'ҵ�r��B�X���A$#�����%	VLA)@��_�D�K�L����fZ!d��"M"$�l�ɖ��>�'q�� �a�W�l�H�: ��Z贩�bA�� ^�t�P�x"ɒ4A<��&����} S�5�1O�AAq,��	����a�	Ȧ��d	
4TG"ș��@�<��d��
V A@s(����~:�I�3G
rT$%��Y�\��e>�Ms�@Q�
�%r7���O�� �Ɔ�z.��zѻ��D"J�5mu��x"�<vt�и��O�i�ϟzЕ��$S��X�% �<��k��{џtig�
 -�����A"n�E�D�0��42�EF�*!�f�Uy��
��\#��/6Uy��&'�Dv�fUC��λ\r֬!�w�XXb�G�r(}��Gɽ)�<iH�P��ퟲ;��y� +L�);DV>MP�M�Ll�0��IT�Iͬ�󃃓6�5�l�?I��<ܛ^#M���`F&4��>.ZH�O�%qv��5��e� i����'ל=�U+@�<	�Nh%pt��#�?��m�?���H2'�lte�?ɦ��Qn��Eep���V7 Л�)i�j��#`A9��<�lڔX�F}����3E�,�"���ɟL��o�j�b
b;Z��`´=F|�gy�)Ȕ� m�$�`���Q!K����!4�JAڎE�\ �Ř�F�t�PGπ4�$�[���5r�h�^�D��k�禑�d@V6�z��?�Jeo��
�R�bR�L�C�^��gg"�O޽�ecJ��t1��"����������L-(촟�􋔵 v���I	 '��x�Jϻ?HX	f�$G2	�|��U�	)9�Qe�לXўɓHJ>�xT8CJZ�6�T�1#~��Th���t�����k(�A�����Ms7ȏ.q[ �vU�p=1�$+gs�pb�O�D}��՟�s4�U���HЯ��K;@Q0� y���>�f�YV�؝(�F[�-����0a�0��'Fh9���r�l�1�b�H�m�`���|��}l�f� �Oh8���R��I�6qλ�-�g.'\��!���n#ʩ��bql��`	L?."�ۗ,��&�t�"�F�K�%�=E��"�����͌e'�q{0ρ�7[����n��.�/�T��BI�V���'� |۠�'�j�"�'X*BF�]1�$�C����'0:�Bf(��A}^��d��P
Ͱ�'��l���ðGX�R�W<4GrAy�'�-c�jԔ>��Y���տ)�P
�'F�T���K�@n�M��N._���'�\a�p��0�رz�^�]V��'@��K�k.��{�H��&�2@b�'&�T�� ߕ�&\�� �Hx �'q|�
�j4 D10N�_�R���'�`��r%)S�P��P"�%�ub�'!�#�Ę"�"��S�σ^(P�c�'����Q!�_��X(��ӧV�E�
�'ʦyC�ʦ ~Nti��+G���'��Q������yqAH3��x��'�,9W�2���@�',&��'��D;�C�]0N��h��J�U�;D�H���˿�H�:C$ǬM9z�Y3�,D�"sl�)-�.=��d �[�p�4�*D���2DO�@����Mr�!�O>D��!��"Nyv �!Fϩ`Ӥ�:�@1D�� t�z��,䲙f�DS�@B�o-���/�1_��mB�� �KV$B�	�y(��[��8CB��Kq�Q,F�B�ɚq����$̑.@2�)�`�,_�~C�I%|G�H[ B�bKn R�o �B�Ʉ@�m�I��]����M-9�B�Ʉ0;�a�A��(~_�1	Я
_jC�	C
�\� �P.lǰm����=#fHC�d�t�s��3*�l5�P�*d�B�=��z�	��Dm:7���:0�B��1i�9rՇ��v�%�E���B�Aw��;Ռ�$`��Ԃ���C��e���x�%�;ಔP�ϸq��C�I?30^8��jZS�#� ��_4�C�I8Ht�JU;_d�3#a�"?A��]*(�Z�k"��	Y��*e�	̦):T�Z�-< Q�3�,��d�%D��5	H�XJ�"o̊��&k$D��q$��KGnh��M�UD�(3��!D�(�&(S,0�2����N��p�!"D�xx�-«1�AS*�C�U1d*D�DY��R6T�"3/@�@�<�H�/*D�T���Oo1;� �S���r�$)D�`�� 	� �Ҙ��`��A���Rg
&D�x��VTD��C�0ʃ�0D�@�Q�� S�%r'�ER��p`��!D��@���t�p_6Ϫ��%�>D�0��� �V�Rd��W|H)�!D�������x[�݋���v�i�Qa>D��R���<8l1��F�l��x��/D��(��R{�	��d�L�-D�8c�-�%'d>��\�&�l�0�@.D�� ع���?k�(#ح`z<!�s"O��R^]��!4�7/y(���"O�e��+�F5��Vj�-��"O��1��w6�٥R�v>�cC"O��;6�4Z-�����!d!l]�"OP�P�*6qǮȋ����P[`"O�=�pg�~�����6��]H�"O��[e@GSD�-�$�Y�� h�c"O�A�$X�M.�Hs&G�7�=�G"Oji��Mq�9;�[�;����"O|J��	:!G<l�e8�X�R�"O%�a���9�
tX��Ք3�ZݒF"O�u��i�Tl|����%�nlJR*Op���ǋ�B�hC���,;���'+��9�a�)&�@�掎�py��x�'AP�cb��T�2��Ң�,|�ơ�'��h� �P8N!�BjFx8A!
�'>�pY�	#_vh�B��p��0s�'�jU���Q#|� �c�c�~��'5���7��]Ԑ�c��M7GbM��'�&}�����{���� ��'�6�"5�ˏI^�˷f]-lJ�	�'�&AWbY';����H�9�j	�'L��▵B�����Bq�����'є�ӖT�5K"�Ka�-g���'�8��/�_`ͫ`������yr�������3}�^Y�t�.�yRmSk�|m{�(�5n�f���oڛ�yҧ\1qP]2��;7�l,�"oW��yr�^-z9�0�2��4�����y�ʖ��2-�7â/�Z\�l�!�yB�1_�q�F� L� ���՝�y��a�!�D��c�^L�3�/�y��7���R�ϲa}�5�ש�"�y�/�
jp�!#�-\vdqC��G?�yr�G"]�Q`�e�Wќ�H�ɇ��y�'��,H ꓟL{�DKӥ܂�yRf�=f(�� �	L�XT9��'�y�	�$Q���>E��	2sg��yR�H ,���1�B58�Đ�2J&�y��\��18 Ȗ6����+ݴ�yB�G"kV�ѥ�Z�1��A{��1�yR��wa�����/�HU�T��y.֏!h�`���/�F1��-�y2-�93}�P��@�O�������yBԣyԼ�qI@�D�49����y£��u��rRK����m!#�_��yr��^�ry���ɨ7��u�R!���yr�	�d�PP9 ��1R��0�G
��y"��sӦ��U�\�/ֆl�V��y�B��>zX�%F��")��萇��y��Ñ R"���*�B��v�W-�y2։B,@CC�"q���f)׾�p>�T�>�uDɒt�R�y�dʫd�̰P@�l�<qsA&;c �h�|�N�8�I�f�'�#=�O�i�n�>h,�J�hZ �V�#�'fh���jT�B�^��R�{���Y�����dD&����:A%(�S@)dm!��J?�j�X��v$�e"���E�!�D�F�p�,��7�vL�5�6��{��+�dG{�`q����ll)b�^�.W!�J�^~��kD�Ҭ|���`X;\J�O�-Z�v���@�-�$�iqO��`���a&j֒s�!��E�y�N�+��A�}H�?����n�0��D�지 ����ȉ>~�4�:� ��"O0J�
͠	|(`.�~���s�Q�D��ɍJ��� �gǉ״���ȪHt,B�5o%Ո0+JsFP;���<E�B�I6].�G�>8Ё#E�+vB䉞f%�%��'�c]�C�韊

NB��\�Ĺ��L�Wa�i��e^�o�6�D{��9O\���K$�aQ���P�u�C"O��ʾFK�X�l �&|��7"OL�0��JO|�(el̄|`Le��"O�t8�L�v.AyB���b9)�"ON�pc��|��� *׷h��l`!"O4�
@.����j�h�q�ĔP�"O�4r��[�T
"n�;*�(���"O�px�E]X�U��*=���J1"O�2�늚_�����ϸL�����"O�L����V$�H`jsw�B"O��2'��}KF���Y��"OZy!��ҥ7�0��G��dĨ�"O��F�=�V=[��'dV �"O:ղ�C�4!t��6a7[ah�[0"O�tb�R�Yw.P��/N�,(�"O2m��� �����cX����"O���3c�_!�= `�	�A��d�"O`M�#����f��5.T^��Ac"O�A�K�6.��Kl�f��1"O�DQ᎛�������!�"Opgl�;
m��	+nxf"O�1�!,��*:�ŋ ��.�"�y�"ONy�˴]���"3NM"��"OX�P��M�l�D������Y�"O0P NSm�L!I��
n���7D��:7���>�VmJ��K�eѶe2�I4D�`��ʼY��*�()���Kg�>D��#��YufHAX/R���!D�dy�@���V�@��P&Fv�t	�C)D�XYrjR�='�ܹ�\�qŔ8z�,D�ly�Fپ1���@��{�n ��,D�(�×�U�v�4�5ds�鈱�(D��B��ۧS��x���/_!�Q���)D��!
��I�� D�߰, V�Z��'D�x�#!�$�~�� �&�(�d$&D��A''��mph��$�L',��D���#D��&�]�83��h���Y��Q���-D�D�d�c�:Q�dǑ�H	S&D�$����O	����ƪB���I%�$D���SG��)�Dłb*�k\$�;n-D��x��D�y3"��&�`@X��8D��#Ԭ2*$�p�%g�0N�iW�6D��YrH΀O3`|�dϞ*�<J��/D�Sa#�8�m��
�>��y��.D���������A�GZ�jA��9%�+D�,;����IQF��*u�$� *O��8`m�;4oB��ՂR�=Rm3�"O���F�M�:}������� ����"O��r��#LmFmq�a�$���Q�"O؝��A�%L�x���D�2�IW"O0J�d�.j�{bj��Z|`D��"OL1t�S�F���	��H|�Р"OI�!V�m��AriF'^�§"O� ��)�?>�$���D��w"O��s�)VQX,+��U,x~RJ�"O  ��F���$H�/a8��D"O(!C�T:Qw�@'g\?S�DQ�"O� H�2aCT"q������ίJ��P�"O@m�֧J�$�FZ��vpHU"O(E�H8��#e�%P�b�1�"O,����%"7�=q�<b-�չ2"O�9v�F�GFx6�I,�MP�"O��.��Q�n�t@ߵ6�|z2"O���X+8FY�<8h �"Oh\��F T�-�g�(y��8�"O��jŁI7JS�}�Х_�\�B"O`(��b�C
*�9�$2$S��K�"O�]j�FG�x�B�;�ܐ&PN���"O 0J��ߤDb�(��"�F��JE"OԤ
�5|d ���4C �$bP"Otj���<7/b5q��x�qxg"O��S3�Wp�9Fȟ�~5��"O^�rT��0-�T�U��V���qp"Ol��'C�� ��`zeJ��(ŎT��"OxU����h���Q�bJ�BT�y�"Of����¨+a����T�L��!"O,٥-�,c�y�� �/M���"O���'S�(�b⁉�g�b��"O�U��D��<���S0��4�l�ڤ"Od	����_���!��ibi��"O����e7JΌ
�f�!L�,l��"O&1�5JH�5�8������<E"O�E ��Wz�a��E�	�&�F"O$���ir^ݐ�C[/��J�"O����n4`"�t��l����1"O��Q��(p��ytI����x'"O�)Q1L�o���ʆ�9Q�l�	5"O�̡�,���KaF\� �&�"OF�b���B�:U#�&��c��2W"O�+g�߬%�P�@爑�PrP�C"O���LT2{�t��G�;kd`a�"O��Y�C_�Z�4L�&
�QB�C"O�5B@Y�sgf����7`S~�"O6��� �-7��R�J�E�r�"O�=�"��%6|���l/��#�"O&�s�Iy��:�1k�e�1"O��7)��˖<k ��]ג]�&"Ox1Jr�J�E[�={���2ȸ���"OB}z� R 6��M�d�-S����"O���OR�m�
h�0�ޕA:q��"O��y�����SۻVD�ՠ�"O8�ju�NPe���28�f� �"O�����
�2�j�a�ED?8����"OȰ�RZ���d�'F]'p�D��"O����P�ۺ(1�F��:�	7"O(�3�tJ�8�c��?ef�Q�"OUj ��Aզ �Q� �p��"O�]Bra6@��͡�OZa�%"O ���Mb&���3a�88��A"O�A�	�
  �   $   Ĵ���	��Z�JtI�:F�����@}"�ײK*<ac�ʄ��	ڤ�Z�xm1	��6��o7$H�p�O
�2l�V�J~�n��VCI�ڱ�`��I	A��,�u��`��PlږP�N���˟г�A5I����������p%ЈRW�tʑ���pH��A��J��:�)� ؗ��#��I�x~Z��Ɯ� �<�A�ڛl%|�HW�����kV~e�'�L�dKˏ a�\�dhΡ(Q*�0E7n����"�x�oS��+�c+��L�	��+�o��A"JP,ōt�uB�9�@�'�����Ǫir��'���2��[��~�T�Zъ����#�����+�~b([\�X�o/}�J� |i�P1�[~�C:�
����4G��k���":�"��[M)xl���Oh09K�r�@O�Ĥ�>3�q��ކ\��GO�a�8��������v!��-Q3'�%��O���A� C�a�w{ �U&Ht�$�`E×s?��u�8ۤn�>�$`�O��󮜠���G�Ku�ۑ
�����ƪG���K�bq �Y)��|����f:��P�|�ӓ@~���ڴQxH+�lX�]V*� �ШQ��p�'^�C����nx@���[1��D�4	Ԑ3�m�-�V*co;G)�����9[�ĒOv �c➽W��'݄�!M��ő�AD�8���IV��4@� �I<AG��a��	J|���	$�*E@�i��t�ѭ��hr�B��i��B/O�P�$��%{/��l���xB���q@T8�$�L����ei؞�~R�	X�'���&��p4A�O"��UN^P%��>$�ڕ:�� w���Q�Yad��s,]�G�,:�o��<�u&%3���:$�!s��U[��*��ǽo�Q;�Y���%Q�QN�ī��1-�OHDCvF�� *4����;�tN�Hq�|�@�!b7R���y�D%G9F��r�_:S����	��!����"O�%zr�  ���?�	ퟌM|�>�fK�+�����#k9
ͺW�̦5[�43S���|�O��_��#`ҎHh�3ꋷv������=i�`P�'����韘�	�u��'�b<����"�|�0����;0�0�h^3+&v�$dX��C��X=X���aQ�^�:Dؗ�X�/� :7!�(�>YTn�ϟ�ᔥ��n�Z��
��4&�B�)z�4]̉'�r�'��O�S�G �aq    �	  !  �  %%  i+  �1  �2   Ĵ���	����Z6����0S�@UT��CnѶS�ԡ@#L%~�@�$�.?���D.C�'ll\�02�8���w�� {�ۑsr8xP`"O�4yR�ž2�Hx�a%(m@(t��"iD�S���^~^ "���L�L�R�A6#��@$d/<E�h���>Q���Q����bpC>����%S &�����60#ܱ�㝲}tHݬP`�!�c]�ېQp h[<3�.|���*(��x�A]�e��\[��?R�xZ3K	(�������y�Z��b̐���6IN	8�!�$�;/�,����L�%jP�"	�_!��� �Z�υ<*sH �"n��aq!�Dy���S$_�_IH���T�`W!��ʵ��0|}�&�V1�,��"O���S',�
�[ )�
Mb��"O|�"�رp
�;Q��./j���""O,eB�LTtR� p��V�}��}Z�"O�#��H�<TJ�j�M��T��e"O� ���.��Ma+�v�vAs�"O�y���[�Ό	����Z��գ�"Oά�#����u��o��A�"O��:D)��~8�eH3�xc"O��¨dt���O��(x����"O�}��oY�21r�c�iW,aav�p"Of��R��jw$ͫ5IۑjUfI�"O������q�Z	0 	 ?\��IX�"O� ��i��e4�1����v�r�"OT�ۇ��R&���S"@��"O��s`)_ v���'�9�I{""O�]xg���z��C,�w����"Op����\�1�����SO�u�2_��=�7%3;*98��R�c>���	��	Q�4�JՎZ��*��ȓD�F5�ee�xrvLB�� UOPmI�l\�y���#o�a��S� =O& ��fO2gb4����>Uj�@c�'�@t�ŋM�
5D�37	��$(t��|�勦��*&�'K�(�7S*lҖ�V go�h{A셮�H��<yC荾:���{7��-	jp�b%|�T�G��?]�H	G*�(VgC��8|6�]AAm@5zA�JFAN�3�l��e�5TTU��X�DT��;a�>�g~� �
f�rR響_���5�yriH�*;D���싋U�(u�\/j�Ԩ�G�	N���U�GN���Ɇ6b�	؆BHf6Yh�5;�@��$ 4[,�ϊ�1 6�秋�be���3 ��� xs�X�Y��	+�'�h�"��G���r��G�R�|HA�y��O�r��H@����k
�r�cXI�'_�����D�|Ϭ��֥A�I��L��%N��"�\<|k���E4M�buP�(@iR�����Y�q�PE��!FW����1Z���dm�*K{�lk!�*%f剕a+Q��|2V/W��,�1'�3ZX�!4�C5rDhD�B�P�r=�!�:� ��$�<nŐQ�cN�?3Թ�a�9C��'�Ը��{�E��|2b����p)2'�%s� ��u�]�4�v#��J�Y�����ywW��B��塍�NT�����%��'��p�pdX4!T����}:C��wˆ��ve^
,;ި��&�Z�'мY2$$�'L����(��U��z�DŁE�DN��\�ŀ)�L��OL|���dڢv����G*�%
�ᨣ��<���U9.�R4��&ؘ�S���R
�M�A�R��P`���E[��(�Δ[D.�I3�'ú�Ң�6n��,��BY%CN�\�H��[+��
��dHڔ�d\�%q�i�5�yr�(qmv Q�ʯR�(�0���#�'��VŽ;���qT��l%��h)�%WL������M���T�]M 6��_����Q1�~�Zx̧+�d�够�-@`��h�*�D ���U�2�p���O] � ��%=�Ż)�N4�A8�-J��I��8С�?y��O��8w"$�M�XrR$�:�����	�� �CU��g��1�ܰ9_�S�'��@���|�ҀW)*��Y%�A�F�ꭂe�
�JMx���Q���jP��
V(��D�+ae�B��E*�@hEυ�|�RQ?aD �[�*�t\��A�����D�+]�ly��2t`,W���K���s�%���P�17PqX�d�6+D6�𷅈�2*�À�Eˆi�Fl/?ۈ	�$����S�	a�3S�	3�r��`�C�z�@�n+�	�^�Ш�V�\�[�̱ȵ������*w������Lc�̆�����U�ph������LlxECX�i\���<q<Me��f≌Dۚ�b�b+ͮ�ٶ��K��J��	
V�������?��L��c�f;,.�ڰ��_���-RO�\�6C��:����nL*� �L؅,��ؤ	�����
�S�? �)��Z�&�h�Bv�h���a`ر"��i�^�� ����9z�(��2�-CC���o��58�II.~.�P� R�R���DY\�.�R�(B��5��˴ܭ�b*��P��+�e�L����:Nf�uB%~b|�Ub`�1r������N?�b}�QjД�56�T+Zԁ�Q�čD��1!V+��'"�����I%Z���L�z��'Sʵ��:�f`�l^1[\R��ԡV�e��m�&�f��)՘�j�Z�!Z\�c�`F��'�L!7KI <�l8q0�R-0��0����423��gŖ3G�,�$�|"5OA0\�9r6�JPb0���O ^�*�\�ni��"iQ�:��Bq�DJ�醦j�� �
ӓ|�i��O�O�B� 𯁗YZ0}n@T���eP85D~5�0O�/9�!�8���P�O�0|�3�G�X�bb��tX�c�U�z����\���\?~X���P�|@�`0B�	05��Ar��'ȈD�(6C�P��4G �x��@����4ma �(r^���?��b��ܑq�ja1�Ę�N�O�Q�)���{�`!��6	�<��i�i����1ċ�1.���&�ǡo�V����{�<���H�/Rz��e�)	[8#<IU��@`y�Dd,yCL��4$���̽ ��Ħҧz2/YM�#c��?Z�R��O�zQ���L�
հ�8K�� ��%�`��`�'y���%�.�h ,�$7�FX��O�As�d]3@Ѥ��3Β�\8F��Q>E��n�h�k�&;�PY@�QI�.�ɢ�[)��>ɦ�K	�ybǽ�r@q�O�]�Х����.{���x�%$WQ���cE*l*��j7����XT�c3�$�ցE-�I���їWA�!:u�'W�$����2x%�[to�7Ѻy�D�#a��-�U�e7�hs�ӱΔ8"��吰X��$�!F�İp@��-t���e�ݱrџ���	)�4�b�ϏJ�d�ST���0h��d2�D��,�=uLPS��Ӏ]�>���'c��M4=�u�B#�~�t��*OP�	���4�xѣ+�(f>x�]�0]��Jq�� ����i��P;� ��I�#᜝j�B�	�/��ҧ(4!Yd*.k���T�	�L�Z`�6I�e��o�o�'m���I����y��3f$x�q��(4� q1ƚ���?ٔ�����7�W��d�J�4J�4�*!� *\S�e��Y�H`H��EC�Rb
��1�O��OڤpFO�:|����HD6(��Z��	-=*p�!�q Q��fъV��Й�$+f@�J��1��E��e\�)�b��eĉq�0��	����H%+#L�d�W�@�g�f�'Ƙ��?��{�g�H��J!#t�?a���i)�<�bM�;��0��4D����C�.U��q�r�M-9L^4�n՞m���P�b
�i��Ր�\��>�j�m�ʼ{�ƛ�8A �9�HYBG���b��mh<��͆�j�P��Y6V�<X��aD������tM���ɊO�Bt�bKX�C5��0 ��B�"^6��ԭ^4Z���z�h4\O0t���p2^��+K+f� ��X�k`.`�FL,2SԬ�U�?#������^�ZY!���P�����W�!�x��(6,O~�	�'%/>q��N��V��h���J1��!/�z��%"O�� dP��LH�HS�[��au�$č	D�㟒�lm��@��LRN��3(�,s&<�!�"O��q�j�9rT����s} ��"ON���D �~���F����i���ɹx�!ҋ[�h����)W��ɟi{�e�搳�@�&�X;M�����W&*�9�#��M���$ޜO!�Ҍ�lHt��+g���U�X<�L�|� �p/֌oa�	;R]���c?��_>m<tm����-t�h 
�i�<A1J/*d��7��;�|�!� T����@n?I�gI?��?Ot��M2#H)�:�4���� e� x�HPZ����'4�٥-^rlkY-� h���%�@1�Q����4D�ɒ�9O��4��$�6����<��ÐS�.u���� np|��N�~�'ZBtp�۵N�T����2�F���V㒢g���؅X���%B>.�.(x�B����d��QY��H�B*�R�s�,��w��c�d�<e���5/�|�zJ�
Z:v��P��|�
a��p�1�ؘt�hD�6"ל;0vC�ɹe����ӫk�
��M)O7`�YB	�
h0���|�T��]�U� /�Hx�;�<q`�	�"^���DD�m�~�"e�'�Α1㩘#s|��)���
ԏ�թF��=l�'��ժB��,���W�ٝC��~I>!f�E�8�D���O+x�8E��g	�'����������c��HX�-�C���q��	�Y>��e�N6�	s� �0'���[��SM��i�� :����) ia�)� �O9>���̓[�����OB���wG�+@�����%`�'�l�����*�\����Q�ft�8
�`ը�*�{	3�0:5�K�X��|��� +L�2�À3�����d� qB��`-̟A��N%N���� �j܂S�W!/��f��%��t�(��!B�S�E<U̓E�`b�l�UZ:A�e��<y���<�a��9�[��VOf[��T̓s7��e虗%�<�z�F�cyf-9sˉ��x[6�S�W�t,2�oƢS���'����Y�E�P�H)�2W����1��U�Xe����	� q$�{�'��.��%^�;5��(fߴ�qǥ��`vbyZ�šs�
��'������ $Ͱu�\�>Y\9�% ��dsT���f���6�ڙn� ��/��rf7 ��f�v��b$Y�
� ��I.!���k�J�q�d�OL���b��#׌%�R���I;� �0�4����x0��堟x���A$UŰ�r�7l��Q�Oh��'>L>`:&�2|�)�ֈ ��z�:!�A&)�.�9�O���wN
��.\w&�ER�p*O/?�1O|�p���[��,=. ڀ) �>z9z�����&�p�����#8��0������9kywl��]t�z� Ѳu4"$��7G6I�A/Ί'��-F|��V��5vL Z�M�J�L� ��)���$`�FL�F�l�ʓ# h�Od�sӀh!%�����ů�~�� @f���O�`t��9:�4��g��C���;ON9�R���R�"P�˚) 7TP�'�<Y(#Z0U{��p��x�V^� *�Y1�΢
�*�p����4�2x{��dx�H�厙�U�.牗W�XC����n�([�悉ty2��|b�`ݪk�Ң�4s.��������ĉd�ȍ���:3�,����[�Z5�b��3�\�2����2?�c��Y.[w>)���;�P+�+HV:�I \�sE�ğ��S�	��B ��iF'jXlӅE��AP����'�f5r���}Q�H =��ځE�l��c�%�ei�6��]��aɰ�A �����9O��<��G��_�B�!�mU*�k�ڜ��O|����] i�V!NoP��'�i��
GMZx֘�gJ��- ٴah�kE�*3[bL��yBgs�!Z������e��8� �¤Vj�� ��^�Ļ�4f5�Q�!ɷ6	��0��O�S?�>�J�Þ�]-<��" D�1���4�i�bL�<0��Ś����v���6��2��'jfУ��@�d��9%�	
H�p��n
�%IҀ�æ=�G	Y9nT̡Eͅ�D	�ԟ8��Wg�}��-q2�pʐ��N��sq.ȷ,^�1#+�Li:����q��+�]�f��j�&Ī���	-�ȹ$�K�dR�J>q���3��O��J��]�%YQF��.1���RbVJ8���lU�<�F�[���7M>y�9{A��1iV4�S��%K���C��w���j]���'���bD�5�jUk�K��3M�i����T��3��p�'�ț'�xRh�0fMlZ�!>���V�ϥ	�Z=b�W1r��kSp7M�%E�d�c��"��we���'�.e�EÃ�C�PR���g��dp��đ�k�����%װ~d�w�Oٜ����V;!���s`GsM�͸")�&O��&��vU3�̬k"m��	>b@䘣$��m���YPP:0�L�
���#��EU ��fw�@���-|���&K��JY1n�v�P���v�ĨKE�ܑ9p!�DW���g+ԓ'�RkG+��t42�d���M{�@V���Qa���64�(E5�"�y7C�2Ag,�+��"B*4�q�'j��s-J�7����e�O�Yf��c�� Qʉy�Z��Ѓ�'�~�Fş<��K0�Ġ^lqO|���'9d^�a4)Tƽ��I,?��$��M��LH���Q�6�OFn�II�S3�Y"���,����$�;1�2����M?OE�`@O}�,,�1aЉ0��|��֤���̓�2�r#$�q�~}C��� '�ч�'X�!W�z;:�ۗ�� z�lmGzbc�S,Q?!x`�C�r�9S ��vǢ|2�i$D����όP��pQO��8tR@�4D�вQC�`~n|����9�P A�3D�$�co	� M�� "_��$�D�0D��C�"R�R�6Pôd�/K�|���=D�Й�J� '*<{��Mh���@:D�P)���T�QI��CO���g�8D�h0�mSJ��J�j_1q�9�"D��qk�=_�x���C[������4D� �wW� ν�F^�i+p�bq�2D��k�`� z!���O�-��1D�<����d3�� .G�`��Y���>D��P㚇XY�II�ǂ4����G�/D�I�a�19��c�˰C�!��!!D���ȡ'��`%�JS��뷈4D��iW�
�@Yɦ�����ًp�4D�`3�����uCcj�$k��%�rO=D�4���	�rO<��Lb��qn@�!�dH?�Fq`�"o �B�R�h?!�2�l�g��<���@�A�'�' 9~��2���#I�qJ�'������"HS%�Ce��'��,wO
��D�����p�'w8T�EJ����5*��'�^�XEj)\����ֽ}0�C�'�|�Jd�=@=�!s�i�J  :�'�9�G�@(&L���J������� ~�Y��	�L���F��Er��"Ol�� �p�����ˣ;�`�&"O���t���v����NZ ��pX"Ol�x2�]2v���"vNJ>M'�\��"O�q�-e�,1:��ڝk-�i7"O֘�'�&j8dACc" F#�"O�*]�6Ei�!�1m`Ie"OL(��%�1\N<�2&��v�R"O��B�����sG��-+*h�jS:d�N�˳mDnX�x*�1ZZ���R?A�6���.D�(����%�����fQa�4TЗ�+D�|[���:B?��P3�ME����)D�x+� \�]��݀C�J>y��,D��'��ԒYH��	�n�Ӳ�+D�hK�韕w�SD�Ի4��u ��.D� q��S�n�kūҸ���a�-D���$��gy�ʥ&�y.!��8D�D@6�B�q��Q�`�4�ȣ�4D�����ɏp*@��/`lj&"&D��8�$�4TY@���'>�JP�d%D�p����XW�4���ѡ3rH���=D�H�Tіm�$�T�T	(��]�R�9D��5��qx�۳�V _`�c�6D�hA�.dn���(�UUv9� 3D�����?{U�T  �D�0�
��>D��J̈́[$�[�e�*WY��r6�;D���3�\H��� ��6}���D$D�4�DHD����%G�)���7�"D�Lڃ��}Pr��E+e���Z#o!D��I'�8TR� Hv��U�xz�>D��K��	G-̨��.��Y��\��i<D��B�Jݴh,X��F]yϔuPe/D���&�H�P��.9�JQ�+D���#���B�Đ�,+
�L0�M4D���K߶$� ��+�,����2D�������A�@�����F��"�1D�;����bi�A�LʥK��	qǆ.D���F�>}N�XR���;[�zhp�!0D��	$�EQ�Y�t��|�:���-D��h�E�l�����D�U�*<c��6D��ʲ`�6Q��4��A�j��MҎ2D��(E.�	�М�d�}��`�;D�T�1H���|,ˆH]1i���7D���4�	�V*��%�Ͷb��P �)D�D1W��D�"Q��`��
�XJ3�$D� �Bg\Xe-��ej���=)q&B��K�:���Ԋ=�$	���2TC�&O<Zdj� R/���#�DA�HC䉤i6j(�#d�Z���eP�Iu�B䉾���C�S�Q?�h�mQ�{Q�B䉢��U�B���#(ܠ+�B�	?E�J!g(1\�	�0�2�B�	:���
d�@
��]jEHV�L<B�� /���2 $�']��X@O�
B�	�,܌�Q U�B�"I���^��C�I��M�f�7p�A���P�C�I�M�d@��-8S�Eid
� ��B�('��p��F�C
f�����mNbB�	 8��iT�����[5ɕ"h@B�/A|���ӭ\0W����%�3;�
B�ɀw���&��*{R ���׋M�B�I�i�~ �TĂ?�00q��CYw�B��y	���t��(�i3��N�lB�	?c*�A�v%U�f��� ���CbB�)� \�*�OЗXj�Ȉ���@�rUʥ"O�)�g�%{̲A��(�qW��"O��������i`�"&����"O�,��� ќt3 ��fn%Bd"O�͸�`M�\7]
��ȻQ���#�"O�с�/#b���@p��n鄤ѥ"OV��p�H�f#�t�B�j�^mi�"Or,)t�͇;�ޤZ�O�wo����"OD��[w�$��thE�[|�s�"O�{b��?4�\: N~Szh*B"OF5��	)_B�#�˟-5����"O��`3L'r3
I�u������J�"OP�;�/L�C��p.
 �bգ�"O�0�1
^��ٔ� H�6t�"O��Y$�d��A�I�=�"OZ�`�K( B4���"��I)�-�"O��3 +��/�"8�dbW3��"O�e3�ҙw�优� ²X<��c"Oh�F�U7#�;�.R#0_X�"Or ���
�*Q���$2��pS"O��AT�N�m����v���y�FP��"OlQ
���1Y���WF#�6UH�"O��UJ�F� .غb�P�;D"O�!p4�g���&�e�F-��"O� @��B,�^8S�EY2�Ԩ��"O��Y��R�Dń�yХ�3a���A"O �J�ƱqX�����^g�'"Olq��!/H���ibCI#oKDš�"O�ؚ��X��uc�aF�]i���"O�t�GF�rd�i��
C"NQ�<I��+wP�:�. �LqR@�R�<aԇI�3Uh��`-B$^RPڑ�Ye�<��Y�7_v���Q�Q}����b�<�u��5eJ�t�ac��-�e�<Yf��)��hh���w)�a�`�<Y�$�r� �r�&тI���I�Q�<�vi�/CAdLSF��iz��iM�<i1)�
>�J� 1�<X���:��s�<��$�ܭb�ȵ`�"`�֢GJ�<)4�K���]�䉯P� �R�%H�<��X)�r��tK(!Ѳ�x0�@�<��ŔD�eR���/E����$��<!hĵT.���!%>�N�)���_�<��S�<Ȑ���c�>2��a�<yue[4�"�_d:�)�/�h�<aDF+ ��<�NC��NL)3D�m�<Q�l��g��s,)�L�86�P�<��ꁂ@�����Z1`���G�O�<a���!d�0�$J�T�tpf�I�<���ŅŒ�� �`��e���G~�<���@>i�(I���	)�8 �bU�<��Qh���3�ٺm�C��y�<)�6.��|�q��8&��ݩrhFz�<��O�k�xd�B��514�25/@u�<��N�#���e��0K�&���Om�<��@�MR�bԄƬW�N��IXD�<Y'��V4�E��=@�`�sJ�<�B��!��IAAh@0 /�I��cB~�<Q%Ĉ�|X.]"��פQ���q�%b�<!%O�<w&J+�+I�$B�A�^d�<���f�z�x��`�ԭK0Qd�<I�����h��A�+J�Z�[Dk{�<1$`�*|B�����Ǽt��	�{�<�Ve��w�L���
8�c��z�<� �`�C�M�}�8!qA�ɠMא��"O���l �<	�����Нs�]A"O��K���	b��QNϷW�V"O
�����-����AL�p$��h "O�ų'ذV�t��� �<��C�"O����쉝J�)�AJC)c����s"OX�KPĖb �*IX�d����T"OVI��Ա?i�L�chW/g�ؠ�"ONh��(*�bi2�f�5ሴ"O(`쀛L������ކ�DUj4"O��в���>�2��%�2T0�8"Or �b��8_�41�DҸ(R݋r"O����!޲&,�1�td_�zsf�Cg"Od�#��
i1����MUP�PU"O<m�%��#�p�ZŠ2k0�)x"O�8�N�4��	{�ů?'�Tc�"O�ph�o�d���P��(*Z-2�"O0L8��ʬv�&�+��n���%"OJ-[t��y�paғ �M�� hV"O���W��3M������?2� lK"O��aadt^&Uk�V]��Upq"ON�cfR8��x��.�4j�uS"O�I��?�>��:`_���F"OL�@�L�'U����lM�)Wly&"O��&_4;���.R';Al���"O̵�r��Y�J���MZ{?рE"O��3��G#��%[��D�b0�I�"O%9���3������
�;�����"Od��EF
:2��"��4Hn
u��"OB0��1~��dH���Fn�t�"O��A��6P���p���Q��!��"O4��$�>O�(��J.�m��"O ]����& ���Y|�@ɱ�"O0t�wDK�b��. n��"O�q�$+D�|�� ��5u���g"O����%zE��;����l`�"O*�m�^�|5#G螒4�� �"O�4�Dg��k�-���'f��x�"O� ���R�D��1�ђ����"O�`��j�' �ȸ҂K�hUxq�""O, �f���v�Z�b`��X8
8��"O��9n�'7�L��r5B(J��U"O�m;V�CVa��R��"Od�[�E�V���
F�E-ل�C"OVL 7@_�s���!���9p"<�7"O�m����^WR}�'�ܲ�||��"O������[O�����s�<�0�"O~5�CC��)�hQfɅ�a�6�QV"O j ����Pq��P�x�� �P"OX�)q��JQ�z���Va��"O|Y����L%T�c) Gւ���"O�=R0_ϐ�G�gm||yF"Ov��6F��RU�����Zr(�w"O��"��ɨ`-�A��-^�c"Ohȓ��D-ZZx��B.�Œ5"O^���ŇF�><�K�&@1)�"O�5@%χ�R�Z����01
���"O|!���M���8ȰN�%�$"O�d��
O�Td�ieMǂa�n�4"O��I�h�$|���s�Fm��"Oh0��J�r�f��I��2%"OR���AȚP	�鑻F���ze"O�T۰�V)�A��h����k�"Oz�h���*��]�3ə�:<�"O� `�q��W.,D|y��*T���Z�"Ob�X�^� �bJ��^"f�X�ʔ"O*\Ag�̶�\u ��3u� �J�"Ov��a-��
� C�-L!��PM;D���]%DLpс��?3��6�#D���`d��%y���
��)��C�	���0f�\�����g�1 �C��<PF�[���5E����"�7C��n~��J7-�f���aQ�� ZC����q{��ؘy�ne[���(h�C�	�!~i@�h\gob[6Ϗm��B�	�8����̗��Ny1pN&�B�	`��X�W���"�JU{���x8�B䉵L� P   �      Ĵ���	�����t苑?�����@}"�ײK*<ac�ʄ��	ڤ�Z�x�͉0	��6��1:����K�E�a�dj�0(� �p�Ã�I�(0�@���yq�eP��u��ߦC\lv�V$��̟,`voК<��ya�K�	?�8���+� �"X�X����$t���L��V�(Cr"0�7�ͯ2��y�����xY��������	*)⚠9�f�D8�`�İ�s'|���'ܘ�Cn�"p b1������X�f���H�5�x"�H17l�S���t$Ԋ�D0����(2$*�B��,D\Ăs���8�*�ޅ���N�m2��\�R͇I?!�%
%rap��7�Z(�Q��e?QR�1���"��>ab�AF-���%�3?���Y�Q�& b��G�@��7�ݚoJ �¥��#=�8��'gPh:ì�q��'},��%�[�\txMZ�/�(o�`��D����O���	�&{��	��]�^?R��'�jayC�����;=È�K�iS=mm�X�L�[Ez���/F:*�V�@0��' (y���eyb��OB��K�]B��v��y
 ��ᜏ5_�d �4}ROF�s-pHJ>I�H�Q<$ m��1�Ry��`̵K"T�S�<�j�4�����E�I(��K�DE~l�O�Dl+a�ͯR��j7$�:��s��2��'�F��%����qA^2��M�O� aEe��J(2��$h�
�� %�l�̋
\r�%>�PD��*�۴at5��m (��S���$��P�'I ��Z,K�O(T�O<�r�\�������^�1��6
QA?���)�e O�����'��M �H�aŲ���/��m��r��Xzk�L���^�����8?��;�4O���'�O"��4m�ͫ�iO-Kʦ-Sv((SZ0��'���XWL�'k_�'�R���mٴ��u>JɐƄ�h��z�LW"�� �2��gBj�$���&��`[Xb� Q�G�w�"(FL� A�9��` ��4����  @�?��J���'��3zQ�B�1�|9!�/�(e��U���G�Z➄F{J~�l�
VQB<2S8R*l}a�IG�<1�aG�C1�H e´��HQ�J�p�'�ax"V\@�#� ;��`�҉��y��"1jF�-[nPQ���P��M�0�^$}�a~r�� �2�"�,Ob9����?��=1��iV�ɦh�d����^~n^���E�Y�C�	�.>��i��	4aXra�C�\0��=a�'E��P�kC? �bY'#=b�2���7��TɰŖz��a�ŋ78s�Ez"�'�8){r�E	}'�Ȼ�+X�n<X<��'�~	#��$�&�Qi�j.���'ݘI������@_&]W��	���=l[y2,T!S$dp�#�D����ȓY��1C��H�U���&�O���Q�ȓ#��r5�N?�d�3̅�o�d���I��,!wn�
�N���H=m����I���Rd)�	���Q�	�����ȓ,\q`��2}�5X��@��ȓ�v�j"/ͅx�n	 ���~� u�ȓ�"���j���N�C�>M������
�җF�<@�=�KE�lS��ȓ?l��k䗍7O.傶�Z6[C�@��j5  ��Ą�R4�1!��6l^��ȓ-�`�o/�(�'.#�\�ȓV�Di�2
8\���7�#PT�ȓ�TdcpFݲ+��m0��@�(��4�ȓ\L"`i�2x�;��7N��ȓQZnܑtᔍk�H0K��Q�r=N}��6��d�,(���b���X�����8�����G�rLB���J2OX���g�R$�0F�R�.m��@ V���ȓ+]�H%��Z�J��3�2(�$�ȓWŖX�Q��-�8̱�e�o��!��`H"�ƙ{�"��DA*dt ]��č1��:>x����.P� Ć�*?X���JD:E�q���Q.���B;�%Y$C�X�a@"Ž]I����@6DI���\.<J��xH��fM�$�� �~Y	�85r��9��U5mz���ȓL	ި��lۨR�D�@��gۚ4��;bh��Æ V"L��H�+����nR��D,7$ݳ ���_\q�ȓp"�I$@@��,�A��+=Dq��]L��1�S�)I:u5��!i�i�ȓ=����a#C8}�0���GMi�̄�	����]��:ID,H�o��a�ȓ"� h�rf��0�|��]!���ȓN���"��`M�h�'Ɠ$�pm�������
T$I��A oT]�x-�ȓ )�`�$It�dq9`LϵQ�(E�ȓ,k�M�E'�5'lq��O�	L`i�ȓAI@��!�O-)��a4�\�P��ȓD���
E��;�(�a��� L�i�ȓf\,���\���P�W0���Vl6��Ëӯ�`%���U�K��������I�$Zo�5�����<���ȓ1Ѩ(�3���p�|��40<����e);��3;ˊe����,⸁��S�? �0k�m�FH~����O�a`R<�"O�� ć�Jd�d���UL���"O���f�_HCh�K��9��i�"O�8d�!1�FE�@
�e�N���"O$��G�$x�в̙�.�h	�""O�Dآm��dQ�@(ѹ��|;�"O�t���.j�l}&�_�}"�]S�"OpQB�� �T=bg��u4�1F"O�-���d
(`����m4��"O*uar� 0~	F��/;n��ܛ�"O>�k��H�N�Q��M�:n j,�`"O(urR��9<� �T�Ĵ ı�"O��c*�5D�|�����Xq"O��ꟅzqR��c�w�ތR""O�j�H%yĨ^�f��j"O>�9���(�v,���%}���"O���(�/4�R��F�:���j�"O�i���T ����¤@?y�h�S�"O�H2��6����	�u��"O�*��F� ��u��hӟ��(C�"O�;Fi�7W��Ƨ�>ouFو�"O�}p�3���Њ`�Ԃ�"O*�����Pr�hy %�a��H"O�Y4��y%�P�Dڐf`b���"O��
�@�<	��� ��P�>��"OY�� �?]�` ����N�T���"O�@���4� xU�3�|�pa"O�����V��2�̑~>�"O����@36x�P��ټ p�Mu"Ovy��"+���k�ɞ.3V�4�"O�"��<|^$�w(�*JS�ɛ "O�������(&*�x#Z��e"O����D�|j���5"Z�;'"OP����Yt�5���ЦFf*��"O����ބ\6j�3A��{We�2"Ojذ���=� %0R�ʣ'Pj�"O]*T�ӷ6� ��ao�|��J�"O ����&/��\��(�b���"O��ɘ���d�>���"O�Ɉ'�P���R�Ť�Ru
�"O��c5��g�
D�U�=
Ɉ�˱"O�d`oͼZED�K�&Ǳ7�d��"O:DQsd�R�,�	�b ��@�c�"OT�� k͚S�*�����N�x"Ont���߮)E�C�Đ,Ob�Q�"O�uJqK�,P6�e���I�[���t"Ozzwb��%ɚ�d"�DX��"O�S�mY<��Y�'��/YJ��*�"O��b�Eη~5]��h4��a�"O��b ��BY��`���?�9�"O�`i���)�>�0�@�ND@���"O$=�gP�u��}X��@ lA� 2"O�y�v��9Tf�=�h�A���P"O6����5282!y��[�H^�iF"O޹Ӏ)Q:c`<M)e���(4Mp2"Op���cԇI%��C���`s"OJM�w��_0�]�臗����"O�����Z�n|���3T�J�YD"O�4!�ٟZ�4��$��8��4"O��#W#��D�|�#��n�|A��"O�͛6�D�*3�hJ���8�LѴ"O�`�Ó7�@��c��"i�1"O���wF6!�~���i�dc
�yr
� *�%�G˦dg�|��E���y
�	}� 
     �   Ĵ���	��Z��w�D:G�����@}"�ײK*<ac�ʄ��	�$(�Z,x2n�	A�6�^�2��hxG�W.:�0و5%J�5Hcn�vq���3��ڦQ	4f���u��A�9���]�Bϖ����?� �F:"0�dYp��"hPi�p����r� �<a��P�8EБ�>Q�E��j����#�6�Y�㓑"v�͓g+ѕQ����'K,�I����DR�Ӯ��Ax�"V�F��)O:��c�ܴ<"<�\��=�F�@h�>�P�
�=�'�
��Pd�<x�Oީ��
�3��haVKQ$]���8a�a)p�>qԋџrΊ��b�>��9�q@�'�:��o̠F�8@��%Y"t����'��a��X�b�t�D��<	CJ�wc��Sr�H���
G�
�t��.0R��-�d�,E>tEa�|2����CfЍK�m��@
Y�F�ġYO<r&9�6�'���C��7��|� ܩ��J�I���D��4 �i��9b��0�-=�D]*��p�t�|b��D�0��r!E8�[�Nϲbz@�S�. m�	�a(��D#�S�'Xh�Ծi�P�E��5s�(�����@ia�O�M�lC-'�'$��ȓoŶ&��_p���ޠWz�]��.��9w(��O��i&�lp���G��O��.��$B$=!4<~��!�!	����2�xr��w-�����̈́��B���jӆ� dK�'y�f�A�<�V��U�(�P��b��H�?IWL(�d��[���92�X2B��튷@)U*����O �$�N�䱠�ʵ7�㇅��]f舻��B�s�hC�	.��%�O�$��OD\]��	��5޴>!��:�={R8��
�5x�⥕'�2T�1�����
XD�1��j�Ɏ%JHIÌ����R���JDl���+��<�ړO���1�0�1Ol��� !��3`�'*�	7��,1�C�	>fE��  � � � ���O^���S�Y�V��$~>,H$��/L��ebHH��y��0p�(�«��G������y��rWd��`�D0G.J\2��Q3�0=�K<��'�p� ��=Z�V�{3�6bDv�K�'��Q��δcuj�#�>E=(�J�'�0DQs�m�٣��#��h��'���c��Q= �>�S��=����'T:p'#]؜�7e]s{��k�'p�8)�:�<а���S���
*&!��4_r��?sh�2&,Q�z�������"G�:�N ��jݭ8!�$��·�%T��a�'\�A�!�MJ��0悒]�He�3E�$�!�$�8R}��1���)3�L8�u�
�=!��S�]��B��O��]�����\�!�˽3ݔ݀���I�Ld�p䘡�!�M�# ���s���/��M���H�OR!���>i�� E�n��C��^>_E!�ȑ4CJɨ����9��d��A�>�!�� (phU�V�G��2r�V�G�=�F"O�i�D�'4�rY���ƿ|�}I�Z�4F{��)$ 6①�h̢E�Z�!�M��i�!�&Z�m{�W�:_�\��ǔA-�'{����+o��i�UqX�X���so!�D�O�͘��/xP��$͈}�X���"O0)���]��x��AJ2e�����'�ў�k/OsD�n΅ �`�g��i�<A��-V @���]:�@���FSl�<yQDF'Uv�)۱'�>Q$4��(�B�<iU���N*8��H;u�`��~�<i�烦I�:1
��X��Yە�Vy�<�#��&8�IBG �e���rGy�<q�b&��� ��.�m@��p�<��Z�v�4YG+��YO�A�ri�D�<��фl�^U"�*N�)r���%��C�	}���O�<0ڰ�؃��p�+��W���'�=�H�\��@i�#�\h:��'�0@��;U���)���G��mK�'��ZK�
Ai�)A�-����憪�y�� g�2@�Ba��]WHmk��� �yRd�!�x����
vb���S�yr
���,, �OY�T������D�+�(O>�e��3Y5������D������(D�xxB�K6T�~b�a�'2F�!96�*D���ԫܙ CJ��Sd�- �Us�i(D�@�2	�{��A�E���rQ� D��k�BZ�!���N��n�ks)=D�XU&�]�"��Ë���[8D�`��P��z�q�M�p��gJ"D��:����??ʬ���MV��k� D���Dj����B��T�℁R.?D���aO���~u��(V�y�Ac?D��c䉉@q,����0���0�!D�t9��V7޵zr�On� �q�>D��*�K��gN��#)L�R%R)1*O�\*���v �=�R�!|�g"O��`�Հ276U���O�{=HY��"O�)[E �%>z��B-ʟ-<4��s"Ox�C�a��L�M�ǉ�\ZX]�7"O��1�o�
+�i�\> ���"O����-�p�bI�V�O�?*2���"O�4(��@|��x��W�0@�R"O&� '�]�RL2�����F	�"O,��u��m�H�PJ҃K��e9�"OHY��΍��];�.FK~0�yQ"O����/�>D.4y1��iP.Ͳ�"O0	�BK�$�q*�m@�<M�5"ODD�a��E�����L¨D��"OL-��^l:�sL�[8h�k�"O�sA������8�K�Bʈd "Od���H�2��� fk,zJl�""O418W�
�7�EP�O�<8a�C"O2���ϛ�H	 �y���x#�`�<pON�[�+�N�S�4�Kǧ��|!��y��bR&3]�=J fM{>!�d�7TR��(���'<g����c.!�䎐'�	a`�"UO��A���	|!�DX!�gےYH�!����!�!�$@��x%����2��C.�]�!�F s,9
�dƓ�� �-3}�!�$(���a���J\�e�ֲ?�!�\.�LL����&V<�æ9Z�!򄈉n���4ޖ9��B!ŧy�!�� �x�q"�6|H�u"�.k93"O�=is��|xD�+4��92��"O
�#�G���t��c_9y�����"O ��i��5�N�W���!"Ox9N����(��]�_�"D!�"O(M:",O�}"�u�#L�O�V�ca"O�a����x8�<p$	�Yo�س"O&��"��J�@���� �{`���A"O�A�V��8��d�"�� �v��"O�	�VGz���sv�R&H�\H��"O���G�X�XY�@У
&�:�"O����l�Ƀ�Ol��p"O6�j���xr����3��G"O(���W�D�P�B^'�h�Zu"Oj,h`��!��a�lT5M�(�z�"OHjf�s� A;g,@V�P=�R"O����Ir/������N�n��"O��PQeY �zi��뙺fv�B"O�)6"�c}~�Ô툦.���4"O~��Ǜ:��i�k����KA"O�l�GƙوfHPd�삠"O�d+��  ��t��1>�$u��"O��s䇀 u�p�`��
�N��"O�8��M�Q��Y�c�#�n)�D"O�Ӥ�r�PP9S���0�"��B"OX��`�XBD��3�&x��`��"Oތ�֯S�<a�B���l���	�"O�Ղ�
�(?�^���NST�R�2�"O�d��	:,���эߒ(��|3r"ON���A�8
Q2d�h8��5"O"�"C׼[� s��Y�S_|��p"O�����]��t% w��hn�H�"O���G�  � �� �S�{0"O~%���U�'s�9���]�UJ�� "O4S���5M����C��ּD"O��H�,R�k L<A"�����"O�u�_�(,�T�̥z��"O�P^�Y�ٺw҅l�M�f"O$�(�`�60�ɐ�b�F��1b�"Oڼ�@O
�p�$pA�M�$�v�b"OB���e���L������	j6C�ɠ��D2țiv�(���o"C䉅��8wGR8b�4])b�H�>�LB䉠y"ּ���Ќ� ��ȱP�HB�I+>'���uAP�����Aȱ�>B���dx��\:4�,(���4�8B�I�;�>�bV� �"�Kt.\�Q.B�ɏI��pB�g¸[����JY�m�,B�I�K-��2�/�/g�a���?a��C�	�W#��Ǘ�\�� �ʑ���B�I2br�$�q���D
\T��7��C�I,g̰Yv�G�c���Q��	I��C䉗s@r]2g��JTVd���6B�p8���v[*9�a�d� ��<C�I�(�N����O0�5�K��C�	�2;���#e:�D��(K;T�C�ɯ�\,�7�ś'G����3^EB�ɝF���˒�P�7����tHUs��C䉩L8x�cEI'/#ZM6�5"�C�?�t��RG�
Ti���Q9##�C�I.~k�ܢ��TY,"�b7'O/`�B�	�D� *��
�`�����8j�LB�	 td]Cb�G$��=�6DJ �B䉴)�������+l~�Ĉ7�PC�)� <�WaH
���K�Ql�)�V"O�m���A�w}	`
1K��|�2"O8)zC�J�,�n��h��,����"O�ږf�3y���''[.3�̄�"O|�JtىU�Ƞ{�`��+��'"O��:�͖Sc�pr��7$����"Orl���6$��h va(t��x,!��˞	����0e��8 ,̃J]{�!�D�)9�N���N"P����![�O�!�D�(� F���xU�Å�(�!�ě��2��#���q�V0��%Y?�!򤙸��#�]� &�sϙ�i�!���
+�|����0����LݲG~!�d	�0� B�[�m$�i�wɛ�-a!�DJ�e�����ӺNo�i;T�O+!򤆉G[Py�nޛYA���'޻u!�$%�ڄl�:�*�K��!�$�"2���P}�.<R�䓮g9!��N?O��{�ƕ0'�X {ׂ��f�!�$y�l��� y�J��Hʐ^5!򄂭7t��`Q+X!*��l�#�C�"!�d�7�`Y��&Β5���(���!�$)j�є ]�(|ؤr�N�i�!��L(c"Dj�F� o��q�Ҏ�!�ʊS���VCN�ua\tہ-�%F�!��*��_Sq��: ̇�Er!�DV���S-e,����'b!�K�yl�y�FEC�F5Z=��$عZ�!��	F��X��o.8$v��F�5Nr!��[�W���C�C}L1ʝ2V!��,]
� �fF�� ��A�2K!�$�(w����Ǝ�\��T�U	�!�$§x�Ѷ��Bf���ŤN!���?x̬��˛0>n9���ٵ�!���g�ּ[!�Kc��@�#kͼ�!��Ǒ�Dp�#�ɜZ�K��̸+�!�d�e:>i�kP<��p��^�[�!�$�IЬ����8��̸�&���!��5��<1隘L� }�#�,S�!�Ā`G�!YtF�����k�k�!�$x�@m��=t��`�d�@\!�.n�XU8����q�8��gnH!�D�C�<���l��gu�I�m��12!�.Dъ�
FDK/,���bI�r�!��1&�j�BQH?� !��'װ_!�����KcGT=r�VU�C.!�$�0p��Q�lA� �d��AխWp!�$��Dn�0ũ��2�l��DE�!�d̲/N�g'�~�H�SԚ2�!�)"j8��g��S#�9��D&`h!�նv#�	K�N�\���� 
gg!�Ē2
cJ]��L�Lz=��b�))D��{�-^9;���yF �1��-:�E&D���GD	�Zp���L=��=
�A7D��kpI�	B�P�U
�et��b!7D����Y'Vu�2�!����4D�`I� L��Z(`&���G�!8�)5D��C�&Y�Lh�M�c�u׀��6�4D�H@CG"p\���W�wjl	{��/D��hӀ�Z�P��&�X8;Q����)D������m���iW\��q':D��i�HA8`6�1�aW>�ΑQ�&7D�̊��Q����{u��r@�q9ҥ7D����-'wҘSW��'qb�e�$�6D�� �+T��=���t�����LCt"O�M�6gO�Jc.|°ȓbdJa�S"O�ĳ�E_�",~)� -QR>��P"OH=Z�`Y�p)�M;��Z <��h�a"O��`�dT$�VI&�{��	""O�K�%�4��n��Z��yǫ8D�+��� 5ߌ�*�)Z�Z�I�1
#D�h�H�I�Ω
A��6M���k�5D����ȩ+.�T;q���1��uc�!D��� 	^B�r􌔁t.j-S �9D��K�M���5A򥓄�2���H8D���g���0�NA���X���hV�*D��k� C�!cs���B���&5D���G�ݽ*�D��"ܺ1���؅�2D����I!SE���ƛE'�I���/D�p���v
���7�τ6u��(D�\s�D[��ȳ �"[ T:�g$D�l .���PTj� 7�.ݘ��!T�(�WIɶ%md��]6`:1"OT���`ҡd��[��C�"-��V"O����c7oX�ɺ�Lǋd9����"O48`�ҕ>��4�s��1kTX	�"O~�h�G� lfҜ�V��G�|ٵ"O��3�o�g
@	�7B�M��d"OD��#�(?zH j� ]�NAx��"Op�*��G�[���?��ȑ�"O:���W�(A��J�$��Z�` "OYdŏ#Y��@ ��
5��|�"O���."�8�ɑ��+q�Z��P"O���c�!V��&�8r��R�"O&�8�M]��<��B	k���V"O��D��i�ҁ��Y	��Y�"OB����M	 Al�X`!Ұ���SF"OԭH�$A�� 2�_�"q`"Od��� %jT�U��gж(!�"Ou�5��f�|1%I+A�����"O������E�,\��b~���"O���#�- 0�.`�IP�"ObɣQ�z��$8����W]��`3"O�5��Ds8��$-EqgT�z�"O�Qg�U'cs6�uA�w[PK�"O�0�',Qf<�q!Z�XZ=��"ON�����,#���΄�V>�J�"O4� ��զW���;Tm
:;&ɪs"O����Y�h�0ub���� ��|"P"O<l���ߗ�ȡ[ՠR0{Wpm��"O�ܐ�FQ�_�v��J$O���"O�����c�]��I��LEk"O�]�J�*"��iصi�}FZ�a�"O�9z�B�I�D�G�,D0��"Ox�3�Mn�h�U;SR�X�"O��Ȧ �v|��kF��
	�d��"O�9r!�&)2ԭ��F�Y&�<y�"O֝�A F���"�!����"O�X�c��W�����;h�D	t"O.��5� 6H�bY�6���d��"Of�qUi1D�J	��G�-K�(�#"O�!W�S
o�2$����Tr6̲V"O�	��?#d�Y⠫T2hh+�"Oj���(�=
�(ґv-���"O4�#I�)<�`z��1u�yz�"O<�C��	
�\5Ae�E�����"O�ZWg�+�ℚS��7B���D"O6@H���nA�����9:u�q"O� �Pre�LA@�,	�H��o��j�"O. +��2t�)a�I�/���"Od����S.9�V��/�xP"OP0��^"���t��3J���"O������G�����^�f�RD"O�d
��ֱ�y�C�ļs�"d�"O��B	�R,�Y+t$�g�&�ۆ"O�1�t)��w0c�!�d �<�g"OtDz!MZ�-���sa�$2j]�p"O�`�JV�| )[
�7���)"O�IJ��˸3+�4�@i����h g"O��p��Չ �T���HW�i�B@"O\%�Rɓ��h zpGѯ�,�
"O
mx5��t��aB�e�r��d��"O�1����C<r�:P�͒&�xl��"O,xЭ�
M͒)�
E�
���!Q"O�b��"a��LR$&�=�x:%"Ov8�S�>D�D�1F���a���G
O��"�H�Ԩ�@4��iXR�D��yRo�<HM�;�oL#�q��)�/�yrȂDp���l͗?�2"����y�EҦ,P:�k�
O�Pq��a�ƕ�y�-(�5i�ZS+ óL��yRݟ q��i$�T@��+�i԰�y�@�n��w�+w�(���/��y��Z2Vyv���T�1�֌R慑��yr�*�,��Η<��@��`�>�y�
!4r��gh@�<��-@���2�y���cZR�\�6� 񪖎���y2 $P��x���.�h�����y�Lĭk}�	�G._�q��m0-�?�yR�H/��L5 �s-��l�5�y"�IE$p��I��b�E����y�kG����z�_!�	Z4����y����YT�ق$#VCx��� ��y�ڹ#E�h<6��[Ujן�yªķ6��`6,ҲD͜\�t%�(�y�KH!qGޤX󁏻G���FI��yr(ǪX��1H��(3��9�(���y'@(�� Q�ǅ/H���l���y���Y�� l9z���� K��y"B0d� YU�B��(�g��#�	S�H�5И����DI��`I�dh[�k��I�Oѓj�!�d�d :�d�<i�~�0���n�b&��AK؋�7|O�y�C��+�:I��ǂ�R��5�'�H�6
�T��-1�4?�0���b�iΠ	�IP	h�8����#e��D��a ��%���=�S�WXІ�`��j?Q>I(' �j�T*��Q;O.9��n0D��s��0u�p�		�a q���N;#��%���A	e���I7��"|�'�{�b�,�����4Tڮi��'L���[Y�dAk�-P�J�6���D�Ic�9ȵ,��b�i��c|ʍ����U|�Ӱ�C�J�p���I$.���3��8aJ7kE0=�C���5>�̘wV�\|�Q��#D��X��F�.9Z�b"(fH�%H�<y��b����֣**��acK���� 1o�
u�b��QE�|%Hؕ"OjU�#!�|���a�k�祌Y�<���+�<CS�(���L2#tبM|r��dN$F@hQO��p�RAH�:��~2�N�:�Z!v�wj)v��iش� NL�a p�9�Qf���V �k��l��@�W���XtaD	'�,���7�m��s*T=�<�`Q�Z�1���fI��.�=�N�tr�X��	/+��ԇ�'� ���
�Q�ΕK1�2?s��ϓN��PQ���;X���� ����NT�Od�8A �f_��qweA�[��\��'��yW��O���f'�^5HDY%��p�`��T
	�hļ��#��I� �1O68� ���U���j^��a��'��q(�HB��� ��iQ t9�P��玫_�PL��B�/�98g�M�hu����'e�}j���w���Q��+h�+��䘉0�0�*�!<g����7E��soӫ�B�C�1�D]!wM�0r���ȓ$0Xi5M�o�~�"2*3 [lXoڃ*����A�,WKXY��J�lFz�������56����
�EI��{6/��yR��4}S(0�A�(=�ҁ�%�ڋA��p��%�e���S�\�\}��`���PlU\�5x���)�i��p	D�Үey 8����_��d(�AǬZ�l��6�A����"�3Tܲ��n(k��xT��<(~(SӓvKYі�Ȩ}4KW�̥z��pFz��:&��\���=���ᆓ�CA(�sB芸1E�I-^�4�A�Q��h�!"O(��Ż?����Ҏ�P9ָi���@g�ds�l����.�xЪ��u|�c?�؛,,�hg�3P)�y1fڹx>B䉴H5��k�&��98��xRm�6]�U�$C:hH��#�Z
"ސ8s�~z#j��'�!��b�(�&�Hv�d������H)��ӡ@1�=�oJ�uQ��a���&<��:�L���|kw叞$�d�퉫s��9h��׳;ĀW��@��,����V�q��%P�n28Ì!i��,;�j����A8�ip䘐/�f��0�E�~C䉉b簱�@�����$)Ivn��й��.��EꝂD��c�#~�R��r���E�x�+���i�<nأ���cv���$t��Ɵ����#YȦ�E��3�	�}���2/N!���9}�����s������!9�<�q䎙&�	���mR��<���"��\/�⍑�MľG
H�ȓa��IY"e��b�4 C�P(�̴�ȓz�3�$A�]��x��&Z��u��=,EcUG��}i�љFGV<OҢ��L'81�D��=t�,���(G>H��\��+sT�ʛ7BvP��<B>���Td
Y�@[	L���qOS%y*:��8b�ʑ�S�R�q��"(|�ȓG*1�D��l�T��#�u6�؄ȓA�]�0�H�vŦ�� "ٗx������M����EZxqs��0�1��vf��(����FEܙ��ꘙL�й�ȓ[_&t�B]�Xs��KT�.,j �ȓu�%��'�0���)J��-z*Ņ�	N��ir���Vޛ[����"O��$��2n:mv&���x���"O����.ٸ| �Mr���cܰ�yP"O����<Gʶ�xT�vϮ�3�"O�s��Q=9q�֋\CF�ce"O�Q����Qs��P�̑)��1�"Ol��#끩	��rd	��V�༛�"Ov�H�*8��j�iٮhj���"O�(Kc�.$���B�\"����"O �@��oNL�B!�
'=��S�"O�(�P%�U���z#��= �%+!"O�Pp��ЈP��92Ҏ͙}.h�A�"O�|j!kS0v᰽9�"H���R�"OҬ*��N�2ppbg��l� 2"OnW�I�b [��W����d"�{�<q�NV�x)�œ�
ۧZ�Px{%a�u�<���υ��A�Q��bM*����n�<�+��|ꁣ�l�?����"��B�<)W��"a9VPk����ep�ѤIy�<��u��X!J��T��tC�'�v�<�7�0Sx潩��W�-`Di0��p�<�5hB ���RRL�2y9���c�e�<�጗9pl:���$90�{e�b�<)ff�oDD9�*�a�hXDl\�<����
f�k". �ltt`�LU�<	���!��ؔ��>Č���VE�<C�X�Cm�}�s�>Tc>�s0�j��<��E�#� ��0,ҰW�r��FGۍZ��3���hh<� |(Q�jſNb\���MQ��8Y�鉂/<�$b���'0��c?��V ��j%"���X�&z�h�f&D�|[v�ʗT �1��f�3o^����7eu�piE��Jj�(�Ƶ�"~���$:T9���P(���q�~B�	q Q1��ރ\EJ�{p@��E�IR��)�5dD�B
�c�T�'xV���5w�]�0�Ύ}����ߓ!���	�8Xܙ�H�jֵ��ʍV� �2�W2<ˈT��'�(A���$J��m@�I�Z\��T
)��-(ܽM������[R��5Z�A��F�V礽[f*ݡ1��C�2jgp-0'ϩݼ�e����$��׀y��A��Y��]��J+�g}�`����%M�Y'^�P�˝�y��^�F̌��ŝvr�#�� �Us�lH�m�L���GV�fH�  Zw�Q�80$^�?Y��s$ũm�F1�&-lO���Ѫ'�̔q� ɾQ
���?�n��a�� C�*�P� �sn,����bp�
�/��i���4�ȡV��O,H��^sZ��a��<TN�Y�C�2��l��z�I�iX
|6H��-ք�y��W��v�rp��!��!����NYp�F. X�,�
��.������������exĐ�L��d��@��.D�lH�	�`�~(S�ݡn>h8���%:�P:V��7i�)���W��N�'�dL	r�V/O;Pa@ХF5�f1jۓ���&�\�C>���P�37	���:��YP@ ,�9#���p?�A!\���ׇ_3�0���m�g���0k��6X��랞|�b\&>�(��W�M0�Å��#�b�!�'(D�$��U��T�������d�B��cXR��amԋ���p��-�"}�'�9q��@v��{QI�2T��e��'�<0�%eH$*�X���p�����YP�T���Q�H��W;�F}r�#|�r�k"���P�|�9 `M:�0>!ԣ΀m�JQ�q/��8�\#K�yr�m�=$�40�b^	��?V�l�(� 	S�e�@�s��[�'sjxas,ZݼE(r!�&��O@Pq@�C*p��'T ^Y	�'��p�7*]�E�<�S�ػh<�Q�L�~��z;g��ק��"�/x XéC<�<�ф�0�y�ʚ=5��A�oU!]�����$��T�pc @�̰<�U�)���Ʉ�{$������V����%�p�䂒�8��������.|�g"O��@U��N"*��������"O ���:@9L�0�'�U�R�r�"O�e���%��ؒ��""�:Pj�"O����֬`��x
�Rr�+�"O�U!T��$�.8���͉$%4a0g"O�����X�P!���`)�e"O��;t'�&K��x��� $����"O��c�#n,0�(@9S�$Eӕ"O��kd��m|j�i�R%0bpau"OnQ���ʒp>H�F%4d �`"O�5�Fh��[$蕂��YPty�"O6����Z�.�n�Z��_�h> � "O��A�͛BR��s��?���t"O�  f�KNB���#J�<����"Old��7Up��cr���gl��"O���s�΄!��ਲo�&T�n�P"O��bRbڥ�>�`��#sF�a%"O��( �L�)�\(p&B��P*�*O��PB�@QžP��J/DQ~��'D㓡�XA��r��̻����
�'Y� 0L�(���shڳ��
�'��p��S���tJ�@iB`y�'z�5�m;'�ܵ��&�u��a�'-���d�װ���z�n���C�'�}q���({�*�)Ŧ� 5;���'��a�ȹ"��!�X8zt�)�'b���FR'p�nA�C�����
�'�qA#L�Z�t(q Q$-�
�'K�t&�WF�s�gT7������� �j��#s~����S�$&�C�"O��Pb,I�|f��Ȏ�~-F��`"O�|ʳG��X�b͂�G��" ��PV"O�Q*0�Y'R��m�� 9Xf�Br"O����W�3`t�jt��&E���!"O&@)�kc��А.�8#4ى�"O�����a.DY�w"\�L���G"O��q��2'(��a�g���Q7"OPl�k��?8�]Jc�г����"O�h�rH��jdբ�G2���B�"O�p�UkҶ@��8��ЦGtСZ0"O�s�̓T��2�F�(S\1�a"O�8�p(�2_'J�{���K%���"Ot��N�m���w��h X�Q"O@��(���Z��'��(VJ�SG"O,8hC��P�`�8�)86�m�p"O��1���`��d��� �;�<h2"O��fBR.o�m����e^
H�g"O��8Ã	4I�����NFN�)g"O��B��K�P��܄|UR��"O�����Q�c�a`\P�@�x�"O�Tr�mE�I����FR2-��y!b"O\)b��̣s��ɸ%n�!?�V�cs"O����)󂁣vg_=�u�Q"ObI�S�8��mx���nb�T�u"O�dz�n� ������c1�a"O�`��/ ��p���,V*���U"O$UQ�/O�;���R�(�)x�-P�"O�ģ��<x��8��G��Dj^�b"OРô@R�5$���2P�8�"O���B�
�h��P3"' Z���I�"Od��钋p��c@@�&E��Q	"O�h���V.��$pq.��iJ`"O:�z���_��@�7�՛&m
e"O@P�u�[8�QI�Cќ��@U"O�}�&Y�"�ش��"aٸ���"O�x ��϶DL�k��Q0a�����"O�,��i��/��<[���"�n�q�"OT�i�jդx#��:��L�mtnHP�"OZI��3)��4�EVG|�(a�"O|؃B!L,r�
�.Y� ��"O^qB%K�$0V#Q�z�|l`�"O�a�$��3 �ըEo͍a9�4�"O�!Г�J��,��m3|wp���"O ��F�P8E��&f�<o��$"O���Q��+�^���^2!Ult�b����L�z���s�����Y-t� 6��3j�*hiGi7D�|�K�,pɰ���$�`�P����O0�׌ۺ}L%��ɒ~���arn^2P���s�_�I4����W{��ց�'$��ƏQ�޴EC&
��tA���fd�	�y����yDd`�����hT�`����'�ܕ3@� 
�2�C#�'r���b�	E�a�'��6g�^܅ȓ{X�h��E &Kj�S�J�$m�9���z'JP��V�<ن�R�����^0�[�JN�m��y�aҪ`2!�d�X�l����O���Q	%�

d���ǟy7��`�\Paz�h�(!�0쀥n����<�š�7�0<��!�,t�`�hf��Q�}PT�{;JA{"A�B��脌�)P�JD�ȓ6l�x��-ՙw���[pG�+l��'e��"g��Z��ţcNL�.jxkU�c���XQo�T�g�GL��C�ID��z�6l�$�{&g�q��1�oM#!��p�vj=etZx*7(=�iTd�XR��h�+1�$�RC��U�L(��	��lU�G&ȹ|G���B��pnZ�a�I}����dػ,�`ESwF�4�azd�'�����A��$����_�шO��"�ğ�v����[�J����H+2M��{�C��`�Rw&�bi"O� �1�P���y��d�j�l�S�:O��1��	FP}�F�׸#��i�П�>��E
�0 d4X2�ө0���4D�0��/�t�a&))��]�cMV�����lV?d����Ș�;�~�'}$���<yfA&=����*[1���ϙ}x����Y<c~]�m٦7��0{6��
c>*��B[>ވQ#N�0`^J��#Rp���(�F LR�`���*48�i��I=ғN�f��Ѥ/l�Ł�ԙϪy�4ưj4
8��ĺA�I)e��O��qc"O�I�D�ԟx���2T�`�.�:S�i����?Z������WhT�2�˨<�Jc?��CִYad��4}Fi�dR�[�
C��'"��@Z'$ZA�mS%+�Ra�@Z���'sK�tHѵS���P�&�~Rm@�A�1OF�U̅�=�r8�fm�9ۖ$�'�'�5q�/������É\��0"'�@��d�)k�*��E)@e*��A��/LO��鐦X4���@$-�h؃��4w� q�������\��@Sd?�i�H��M	6��CKF���e�^0+6*���'!Jp��4]�}y��,`"�ڴ 
����")�`�z %YP�X� ˬi���k��6�n�=r|a�˓/R!���=j��	ad�ۚ$l~�X����o��yE��f�Z"�,3�(V�Ԩ�66AqOj�+D,�P%N�xwe��]l֘a6�'�޼��U��1j���12g2�p2�E-trL�B ��y�.<��$�V@�rg'lO�qE\/l�����2��ۂ퉾 �N@)�+�o��� c凍/���'���ID�U�>����&
AE���I��K�.�24�
أ�MG_\�̓u�9s3k <)�~$xЅ�K��G��Q1
QX��	J�ikL��G�S��y����[,@�ᐦ
6k��0W�A�ɕm�QAD.����g��i� C��7�j��#Ҕ��	������&y�N��'�9\;��:Ê��1�\i��'C ݃&̈́8X�����;*F��
�' @mX�Cʭ@�č��jY9.r����'H�%��S%]���A��y�@@�'9j�hc�7��]3��6|���'��R�h(u�F�P��V=�(�'��]��c�
F��JU�H	C�|A��'&�E�\/	�llX`��C����
�'�BL��X1'bm'�K�(|�i�	�'��t*s���1*0�7�X!!���	�'�n��Ə��H���S� ���'��uZ� �:j�JarF���9ϰ��	�'�0Y��C�i����:�D��'j�]�@fX�l��DlE(��I�'8��6��/bPX���ߞ-�@��'M�e*��Ğ���f@�=�<��'-b�� ��:Sc.ߗ.�>-��'Xޥj���Q��U9�՞[����'_J�Q�^'nMc���1t=%y�'��
� $!��D� ����yr��y�� O�E?��1���y���t� ��e��E�<9�'�y�c�x���a��>],��P���y�9e �U��&�~�(�I/�y�X*.l�"� 'S�p��[�y�B�3����'��	�%�Fc��y2�]2J]���]?W2�s�
ˡ�yBU�c	�< #�J�V�M�V�<�yb���"��P��5^�x�2��<�y��%5bp�2�_���Ԑ5���y��*�4���,G�N�@����y�*б2d���i��.�jt��c�4�y�B-&�F4@FO����q��#�y��=:��	��j:��׊�yBh� 7���Z4�I��x*p.�yR�ږ;a��q����<`{@����yb�%4��Cu*ٌ��y�GD�yB���m"�*D.?O�T���7�yB�k� Ie͞*�lIX�L�y
� �Qq"�����s�+[?�>�d"O�� d�IiqjMv�޴"ONģ�E6�\�k��#��ș�"O@��do�%���E�|����r"OL�(�eV�VpȈԊ��]�h�d"OV�aO���j�|����R"O
�X��Y�QV�9j��yV �"O���o�_P�97�B%tV�k"Oz5�s��J��|0���Alfdap"O�\�W��P=�Dc��[����#"OeѨD�9���Z��[u��-Z�"O���Q����ji)�ڡ�b�[�"Oδ���N.C�by�R��j�ƈ�`"OԨk���
4~컆�L�f�E��"Oxu�ΘZ��y�3�ߝ!?�A�C"O:�Y��Ј\�"a��g��,""Ofujf�/1:�!�`\/^R��"O$`���5��O�Zg����"O��r`AAd~�	cp/SS���B"O�S��S0���x$�t��l��"D��@��&W��Ps�O:`�PIRc D���#���PtP�̸\:��IT�*D�\qW�?s�>ȨPl߶
~n��VE(D�X��i��b8��I����:5M=D��95c��r\ =���703��2F�.D� ԇ�<8��q�@�C8��;�M D��P#ŘZ�,`6��IRh��� D�(�!�?Ql湃�	]�+�P%��o8D��JTMG�TP��?�f�@�5D��#RAί=9��4D�q(T�v�2D�����{�	"A�O�$!�W`/D��ɟ��WDҿp��<���/D�Pz� X�h��I�̀d؈��p*D��uń�(���A�1.qg(D�l��l��$d�8c�$o��q��-D���%*S�ijH(��.6g����*D���̍0v���ɷM�d��4�g�(D�p R+��-����J�An�[%�"D�\�M},<�@2�^�JdG:D��K@cBL�V�� �6�K��%D�p0�L1r�0��J&59Rٻ�"<D�pyf	 ,=��mF��|�X!"<D�4*\�Zy��(�oI�<Ƒ�`�/D�|
D��'$�AQa�H�lQڣn,D�4q�h�h��Ӭ��*y�1I.D������~��@ٶ��.m�����,D�У���C��$����5*��*��+D��{���<i�*�Y�e*�ĚC�&D�,��.ނ^IN`���־Q�,���%D�H VYqUB(����o��c�-=D��q��3]�6���-�"�� �:D��q%#�.�F�S��_4"E��/;D�hsvo'�lA)�j�,!��7D����ኡ�L@�%S?a8�0��(D�H�f��6��LPp'ӄf,�)��$D�,k��U�f��d�6�P�R�H�(%D���d�:t�·}_BĨT� D�0�C��0Uh�����QD�Ӳm<D�,�����`0B��.�\0�d)D�+��ގC^�)T�q�X�L'D�PD��D떌`>~��U�%D�(�4'�2M�`�Rǃ�i��XP�#D���L:^n!Pe�1�H�Y�E-D�XֶR�j65�(��`��
�y
� �$�2��'�����Mn���""O�p�R-�9��#�иcj��"Ob-�Y��b !��If�"E"O|e@��Ҕd�l�%�� K7d�2"O8�#7焤2S��[F��1p=^Dˀ"OZ��W��\;]Ƭ�9.z���"O��P�&�+E�l�P�@��@��"O�18t�M�Y�j�*�'U�{�X��"O�=�1'�5rK��2'�_cb�5�"OL�A��>A3B���ȍ�	5^�06"OT�/x@~��f\	Xف"Oyòe�Xr\������"OJ@���eڰ�wFڜUth{f"O�@�p��.<�ے�	�Cx�Q6"O�����G� 
�F�^ҽx"O�0�Ȗ:V����E	�i�2�X�"Oƙ�D�����2��%���"O�h��M�,��I�#��u���y"O*��N��Ld�s��Ȭjy��AU"O����#kW6%��n$GZ�"O^���ǂ�$����K� �̈�"O�er���x�1�Gn�`�A"O�!��!҄߄H���:�"Or���ϟN���9�DE�E�F@� "O���!��,:��# \t��t
"O��a��F-��\ږM�Ny 8y6
O�����h���N%0�� ��ѦD��d��u�O0��0���O��*�d��D��)�"Xf��g%("Md�R��
D�)ڧ���F��W�EӲC��AP"�ߚ!n8�aet~�d�?5Ba�D._	s
���>=�4�����OZm�[� �?7m�2�½�%d�q�,�!�66���2�(Q4)���S�O}�,�'$��̨�R��)~ox�S��zC0%�P��
,�(ӧ��^�|l��J��.d�H�ɐ1n�� ��F:��Z�O�6��_6{���9Qd*
��I��=4(���I�O*P��c��$6���Z�n����
��Mg���?i�)��@�C3!�d١a��lI�b
%?j�fHƣ�?1$��U��ӉLo��ر�ǔ!�X�q���1>UX����xH���>��:�P�'=�O/&��!$�� DhI0M(j4S�B�.C`H9�� ��)�)f�a���-U��\Ä��6�(��s��R�\�Zu��Ŧu��&S�3pl��E�Oz\� �°

 ������-c��ͦEFa� �R|�b�P1e�����O�)Ҽr�,�����/T�X�pN�0/H"�#��RYL��'�}A
çH:$h��G:x������0����c�Q@��?a���O�S�tjX�PؿpC�4�*��:sXPB������0|r$�i���MDrtِ�H�\4 ��J|r `I�t�ٚ���?6^�:��@�ɗ?7\#<�}�3��8KP|sֈX>tZ��g�ay���b��OQ>��eʍ�&�Āxe��0��؃��O��a"j,�i>#<y	M��P�̆Ft����)T�R4Ex��S�|ҧL�#Z�\i�!�9�����$�L�<�E�e�`�T�B�G�<) L�V��̹�[h"�1A��_�<�O�xS��BR��-��Ŏd�<�slڃM#������
|��ܘ�c�<iR&J�o��,Y�!�LX�e�x�<)��9@�L�A�Dr�̘T�O�<� 	�#lM���wo4S!�` f�E�<A! Jgp�V��2w�T�GW~�<�A��( $��a.�	5< G~�<��g��;���Y�#?N�c��`�<��ЂU������U�ܤ�&��`�<	���B ,���
 4^�����\�<)��?�,4��#:@l[�B�W�<	uH�J8��*ը�O�1s�HVL�<�a�܄#\A�C��/T��EL�<� �0�E3A����$�/��L��"OH��T�Ԇ>z2�*
�4h�a"Oz��&@.��aiGh�:%�| "O:��4m�_� e��$��.ّb"OL)�ՋTv�����U6A��\c�"ORY����4|g^i��LƊO~l��p"Oha�E����4ՋFK3b�m(�"O��TM/4�v�S��#V��IЀ"O���%��$���x"� ����#"O����*֪+&�Xr(�1x�t� D"OLD�
�#}n�a[���0���)�"O6��"C�7k�b�Ct�jA��3�"O��4g��e�t���O�@$�`7"OX��� �{���1T$\�a�vp��"O��5H��>�H�`�U4xBj��q"O����O
�J���Ue�
0^��E"O�P��-*s|�z��[:K�����"O����b `ahm��aO��P�"O�Q�e���@"���i��3�"O X��g��~P:�@ҺD�FP��"Of��w�Ӵ/�\s�h �g@dUR$"O��Ad�J�P�G	X�
Q�rR"O ]h0\��p��(��K9B�Ҳ"O@��a׊Pl Z�ô$ִ(�"O�������&%�����. ��B�"O�L�G.V�1P��tf�}��E"O){�l�'=r�����](8�B@��"OTE`����)�	�d�$�n��D"O*�s㩟"=RNL*s��"qy,HkD"O����	+����\�T`Z�(�"O�1 �H�K�T����p�Z�"O̅�c
�(;�� u�;_t� ��"OR�x���/�Ju��w5 ��"OFX��МG�xm�1�
<W�v�R"O��Z����q�/.BmP\�`"O0��Ĥ^�v�x��
>e0k�"O��rgo�|(93¡޳ jzxf"O�كJ˿;[ш��L#"e��Zf"O0��#Y1hj��3�#]u���t"O���)�I�(DƇK^�AB�"O�(ˢ��!^aȅ�<U����"O8�{�	�?h@`�x�F==Inq"O:��!�[9X�cfn@�����"O��8q��'�h2�"��K؂��"Oea�GYŬD��#�%;�b8�"O �P�GTt��e�-��{�"On����� d^bՠ���&����1"OxHK2lQy��I�@��}0�aW"O,є$6�JH�" ��^`J�"OFq��)�(�9�5.�f��"OT���L;\2�j��;] ��"OBB^�ˣ��\�P�R"OĘ'�����dC��QT���"O�q�� 
:+<H:�[�+=V �$"Od�A�M��R  R�ش~�Hb1"O$�k���:�tT��J�C��P3�"O�AڷR�s9��WȤW�0�#�"O��ص@ŘF`�S�bY��"O��@5ĉ�c���S�tq�"O��bmG_0��(R�[P��;"OeCB�V�
��Ȁ��Z?G���C@"ON��Ӄ۳3�V�Rw,׾)�؍BB"Oޠ���{�Ā��k�O��ц"O�q��)���Պ������"O� �����TY�ՙ7	8j����"O��&�@�1���h�A]�����"O�(s�i2j����t��2A�R"Oxm!�k\�!��(�=m���"Oj�;u�3(	��攚h��B�"O��r�D�;o���qďS���j�"O<�ل�H�I���JW��#� -�@"OLa�fM
')�qY�H]���at"O�ѺħԢ|||QW�8s��E��"O�d"gɆ�p�D�"�EL���q��"O ɉ %��%�xȺ��  ���2"O��Ao��4�RF��)��\A�"O2���(�x&��â�4Rr�В"O�Lq���&VJ�3f"��a�)H�"O�E��M��	<A�s���W=�y�S"O4�IvkZ�uj U鳍�5*=@ux�"O�ԙt�D=w��ċ&#%�H��"O������)1KI?c�l"O��Q��	 d.����R {�)�B"O��	�J;-�Qqg�ǕY~�,�a"OHx�pQ�BϚ�R�h��9f�\23"O�J�a�t�$�;��s�(�!"O�9rbB����b3�B2�n<�2"O8�y��[�J�,iF�� ��@�"O��q�
9Q��JamX#69��"O�I��eX)YS���e�^�C�� ��"O@�2b�@9����"^��@"O� ��MZ���(�ro�JW����"O�(�e�� q[���92���"O��+'�!RZ��Bn�V ���b"O��I&ӳG�5�w���pw��H0"O�E�E��.w���Hή:�`��"O�tA�'R_8%{�G���z�"O<�ӱ�� Y���e�,����U"O*-ScA�a�D�)�d��0�B"O�a��$��dp�d�߭[�J�p�"O� o�7}�Tae.�L�"O�����3�ZdH��hA�,Pf"OƱ�5Ő.t�4Y �Ɇ}?�hT"O2T���f�J�[*K!�l�"OdŢ��2.)�Ct�;?�l"OZ��ҁ�e�$eaB+C���"O�P��E9V̞}����<>�\��v"O�H��"M�f��#ŦK1<�kW"OJ��W䓪�I�R 6���kE"O��QE��Q�x� "ݽH���ig"O��E�M�`5���c^��֬�"O�]��-O
eh���G��j�(��"O��x� cBН���J&</\�j�"O�H���	j�4,��OƓY&j�*�"O�����:/k2dӖ����Ub�"O��z��ڼT�D�gmB�08�V"O�)[�N�;e"tJV���S����"OfT���<���Q��1z "O��qt`Z)G�
5�f+&%��s*O6��� �J��-`U��E�J��'�[�	�6��P�,[0&[���'_^�-��f�h�2�W�t,`-	�'[ `��TǴ�"���i��[�'wl1Q���N��P�H!))&�
�'ю۔.���,�@G��i�H��'_�X��"���A�$�u�RD�	�'��@��0���˷K�:oGTx�
�'4,=��#�N�Y��ţ���	��� ��Gîs ܐ�ەK5����"O��H��lrZ�QBY/b�(t*"OB��K=fb!��Ҍ[�h�"Or$�VU	3L!`XAu8���"OH��a?4�"�J��U:���1`"O��8�iԁ% �f��.fS*��4"O� K0���u�f0)��:D�9 "OV��ef��_fze#�[� ̠�f"O�5�h3a�Y��mߤt
��k�"O�Ƞ/�e���D�=>���"O�	��9S�:���,sג�s"ON�rD�%@��%���>Sf��"Oč���Fx:��m�.4��"O,8Y�J0��"'�DB��	��"O�$&��-{ ������'^�`�ۄ"OJ��[���A�hSdI�"O��1q�IMB~��5!X�;�t��c"O�K�ƛ�I8�XS��P9���e"Oxó$�/H����ˤh!B���"OhQ"�	SP��ɂ7蒸 �.Z"O��B�2/4|
!�Ґf�`�"O�(ȥ䝻�,�"�d�4=��"O��-�I��d#TI/b�ȸV"O�t�`N@�q�\h�`���Q"O�X��蘦S��rՎ����XBp"O���ؕp�
гBC�DvxAR"O��C$bkp���+��6J`ܢ#"O��Seʹ{S�x���ճ� �!"O�� ��0]\����H_�::��"O�yAO���I�3H�
J*��;4"O�Pra	�U2�Kԇ������T"O����D�r�ـ�fުqB�%�$"O��w#Ѣz7*�����c$�`a"O�Y����v]rt&�%,D"O��"�׺�ِ��\+ꜹF"O�@��K�O�8l�5�	
Uy�Y%"O�Q��	_�?�p��ue]��=9�"O��tk�'����dħ;���@u"O��v���<���1�#�2Qʨa
�"O9��L�P�N9PpD���0}�"O�i��f1
"���b�Տ81���t"O@�ʗI�=!!���V�V�`=��xc"O�D��,R6$��lQW�R��$<D�`�D��v��h�C21E鷄<D������D�p�B��A����/D� 3��¢�4���C���p"� D����JY83��K��k�<�w�*D�@S��O�� h���:w�@���3D����BO�N\qud�����u�-D����",y���G��\�� 2�
+D��ao
��s�Ǆ�5PP�`�H(D�<`���8B)�bb��V�|Ԉ�i$D�xXRA�2p2�%�m�m �24�?D�$��Ė7o�	� �,��5���?D��Ò/�	$��hI�nD�]��P�>D�x�C�jƂp���H��4��gI��8���$��&�'n��nD�4PDyыT	{�X�򐌛>#���y#GK���I��,�19�du2�N����O�m�"�E�Z�8	�r����7)j�{���#��(6�� 4�� ���)���z����w@�A�*9�@��e��a��I
�zqB�'8H6M�O6��?1)O<7���^�h�)S�K���`Y|�Q0�'T`EQ��<{ޭJFC%Q�$�@�Ԧ��<I޴��/Op���	Bp?�3����SV�X15��DR7�9=&��'e∋'v�b�'�B�)�rxb�M1S�� "M��I<�%�4�F�w����ˠ�ډ:W�i�'dp5��AK<}�eI��6+�|���,Ǒ@l��'% �@�����_����'G;�b����OV���� F��%�V�Am� 2[h�@d���p�'������їt���t��5i�Xu�w�I��y���7/�](�e��R�L�'��YZ�oZ�x�'Ǝ�r1�~�8�$=�	r�%)C"֤)�N0�m�~�y��-'}2�'Z̊�jU��7�ޒrrM�G'Bm�$�*J��Q
�u�a�¢���'P�#M[�ĕcU�A&�cEպ3qg��sf|ę��bʄ�*�c�)x���}2c
��?1��7y��'�O�n��A��p3@b�5"��!�%����'��']H��SE��V����P�
��T�����@b�P�9m�J�ˊ�P]
��uf!С�9��(H��kӰ��O�4�UIs��O
���O�6�K�)<��&F<-���'�J�0^|;�;rL�PڱiBBcRԟ��'�B5be�,��曬I]bu�'� *ș$�C�>KiӇ�[�l�� �s��~��,��&�5p4�����;5��p����/����`�ڡQ��'�r��<a�Fs��~���Ll�t�
�Dn�r7/�W�A+���&���I�F
��-{���聍S}����4�?)�cћF_>��	Ц�	ƅV����Y�o��`�ժ͞�?��B]7^���p���?	��?��Y?5�	�!G���@c��)�~p01?EH���s����y��lJ$�� w"$�:`N���x��kpN����P�� �Q&H�um��?�T@��iB��k�4xD#%�3�ɻ`p�X�sCp���bFj�(F��KG�%�?Q�E����'���ٟ��	f}�A�)	} ��q�B03gl���S��p=��}�����܀�*��2F���dAq�҅nZݟ�!�4�?�pE�?�O)B\���k��7-=��0�Ǜ�K"p�JU1��%�I֟8�	Q�XQ�I֟���/*�6#]V���ϸ���B2$æ
����qG�	�(Z����,�"?9ע�	�Fȑ&�\mn}�4jذ,4*iQ�މZ�:lJ�E�z�V����; Q���$EHB�'�]��m��<���0I�Z��,���Q�$�Oj��8�)��_/]&L� K� �4�[��m*�A��я���P��SDC�L���N-/^Ԁ��s��dl��� �	ן4�I؟�'���
 �  ��   �  e  �    �%  �.  �5  �;  B  ]H  �N  �T  ![  da  �g  �m  .t  rz  ��  ��  7�  y�  ��  ��  ?�  ��  G�  .�  1�  �  `�  ��  1�  u�  �   Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�� |d��"O
`�(�;���8���-0��1%"Oj4��ND^[��"3/9�0|H�"OB���H��*�ʞRy=a"O�味V�!X��!&F�:J�$���"O,��a
���C�Ą�M�"O,$3%o�-���p���+Ն�:1"O��ݢ1����`���y14]2��i�<�6��{_���c�H�`�fX�$Kn�<��A̼VI�xR[�)�Ć�pඤ�ȓA5��('nߡ4�� �)˩%� ���,��r�؊b#`T�eT09���ȓ!�b��g��}�8�F��-? �ȓ
K|m�ș�VṔ���2�%�ȓ"R�X�j�4JN�1�˘X�i����̹	_�jZ��1!g��zܶ��ȓgil,*�J�
j�Ne��i�J%b���f	�(U��:���G��$Y^م�~r�� S�%T"���k\�jx�ȓ|4�1�îJb��@ӵ�ݩn�V��/[`�"�v4�R�!ʎ<��M�ȓ`:��z�ؚh�J�Z��$HY:	��H��p�m�C1��!��B:��0��EnjZA V;9����J[
2���	��4'J�EA�IVW&��~�(aZ��ӹ�>� o�Y�|�ȓ�f�A�
Ο7�H��M�$�����mޠP����/���ANXo*�ȓTv�����{ ��-7�*h��I��sB�8�8���3����ȓNe*M�悡;������X�o��!�ȓ'lj�#F�m�+R&;�|��2)n�C��0S4���T:
b���:�0!��e֊��)��ͷV��,�ȓ0�&�8#���� ع�L�����;�P�AFd���,w�6d��r�EQ�( �gVlɦ�M,H��,DP���|�I	$G#\���ȓ"�)���E�B	yt&B�^�LɅ��N~��\	?Cv@ӎҿF��(8`����y�DG�|�mYDG1E�>-��'��y"	�*]�MYԤG,Czr��v���y�M��ۗU�~L�S�Q���(�'j6�!�j�Sy���(�GD�A�'�l�`���!AnU1�V�GH���'8 81����u���Q�J�5o|��'�QIE
�8��Ё�۵4jxq��'��aj֕yn~,�0�]*� ���'�Hc���e����%0����'���	��g��ۣ%�� �`��']T�BEL IPZ���!R�����	�'��eX�_�\Y�;0 �[�0�H���	}^Щ��*�
�Q#AZ�oL:B�'ȒmIA����{�̾&�fB�ɪD����I#dIh$���/WN�B�I�5�R���
,a6j H����6��B�ɑ�>�� ą-��9�I�d&~B�4x�����S�
��gK:l�lB䉫:\F(���i������W2:B䉁OJx T <\�8�����C	xC�	s=h�s�ߑc�
�3��\1tC�;]$6ih�+�B��q�g��=�c�dE{��� Ԝ��GA��mAPˋ:r"���"O����C�I�BP�W��"H��z���-LO����(��Ml:��mDڬ�1"O�阱-�`��"A�k�|�2tM(4��u-��Ju���@Ўe�4 ;LO0��Q�� Q�2��0DA��Rݡ�d7D��ke	�|,ĺflA�|�j ���3D�P(Ri�B5E^�^���'<D�����Ձ'-��o�*fZF����:�U����dN78@\���KM�m"D !�h��!�!�䞠hHD� !�)��"$G��@�!�$��7����Si�x�P&Ƈ�~�!���T�ȼ�zMp��V�!���%���#�ϋ ]��cá��d�!�D�;��rs�۴��!$ ��!��T�JT�J5n�q��`2�N�.1�!�A�Z5�����*k`����ӣ}�!�H�U��Z^�Z ����K;h���I�*��p�[�7�� ���5c�݄����s I��qPt�Z�d������4OmX��;�NM�t����B����^4StoB�*�ʄ+�IYHq�1p��%D���D�_�-��w�!c�XD	J7D���g��i���7�$��V�6D�a�EL�~����P5h�}a�)4D�PK���	>)�����B]��r�4D���׎��l�^�1.Z 9b���2j1D�|�GB��Nk�2�̗'�¡x��)D��B����Mx@ӥ״��H��#D��(�G�H �����N@ �K��m�:�=E�ܴn�6q�0CP��8� ���s>���ȓ1o
�P!"R+<��e-'-IR���iODЇ��.
��%q�O�9 a^��0��f����O�y�-O����҈����EXjs�"ON`
T#X�f�����7@À	A�j,�2?E��'��Q0v���l��ms�=/Ӹe��'��E�#�z:���S���x��(��'#��Y"ߤ�"u��M؍|7J`Bߓ�ē%K⩀e�A
�l�qG���@JP"O܍�v�݉�\��F�� ����"OP�D�D��̒Q�[>��"O`����R0 ��UM�'gI�"O�9p��I�7��	d��5~4@�"O~��"�7T�n�`��^�0�9�Q�'���d��T�f=Bp͈:N�>��Ńga||r�ֈd�~���n��Xp8D��F=�y����7#� Dt�Y�#폲�ybDt�X1���S�@�Bh�����y�dJ��B4s�oJ�h���Ɋ-�y2D-�L��ۜQ��pi�Ā��y���LV�
Ê�J���J -W��y�i+D j��жH��́�y�+��rJ\X1	��BB�P롫���y�j�u\��"�j�iRjL�
��y2�>L$���A�[81Y#���y�
U#��=8�W,bӜhQ�f[��IW���O$��BO�~0*�"%��\~l��'���c���)�� 2`�r�� �}�&4LO�a`���\�I�(��+�O�Z0���;�J��D�)G0�c�6D�Q�/Q�:0����Λ*@N��Q�!<OB#<yT��IמD{&��E��)Wjd�<�S�)$�a0$��LB#X�<��
�9O�D��C�-� k )@U�<� z��G�T��pC�V�P��4"O@�SrL�+i?`ґ�
���aT"O���D  q@]�s!Ta��K�"O� 3��C4<->x	� M{�j�q"O��3e.R���*�I\�j��hJf"O�A��I6=��)s�>��Z0��/�S��5��"AU��:-�KY�4��B䉪B��IG]J�
�(�/�pD�B�	�6L8���f	��X� � !�C�	.p�^@�t���!G�hB��ȓ3J*i�D��$�X�ǜ	�ɇ�$��X�w˚B�@�.�)8�1����(0�e�b��g�9 Xi&� ��)��x�����Pd�~AQUC0��C�ɭox��g0w�J��	X�<e�C�I�o�$��v���+6�#�2�C�ɏa˚�Q��82�p�����C�I�f?�p�pD�3$8 �kŊP>�*C�ɐ�(����J�8S�o�#v3�B�I3$�R�� �0>OY�B�,)7�B��l/��(s��/Av����@ӆ���=�Ѓ�!
�T����;DVy���n���ˬ<e.�1��!<����} c�yyz��"�t3�]�ȓ}��!AB�'(f0is�B*Sd8���p���a�$e�z��v��?n \���;�Lp��]�Y� ɦ�H�|�������C��h��� ��n���ȓC�@q�v'Y�U���0a�R�iq<U��I`j��e�}[�`,��P9��E�<���!p��+�De��ɒJ�<�A΋��p%��i���"�J�<i3�͟E�\۠��+�2a��h�K�<���5j$��gєZ����b�<i��K�(�B�j!�RX4ڈ��E�<��LWe�XRh�ք1R��\v�<�FNʗ���uM�P��e
�CD[�<�Ë�_bVq�c��"����nOW�<i3H	�[��B�܅aI��G��U�<�2�ܛEP�����U]8��j�l�<Q��]JXRB틶CS�U;@QC�<�ec��m�L�g�*ќX�qH�<1F��
VƎY�W��R>AAP�XE�<�"�ў'���g=0�8�	�E�<�s���{�b�p��L�ss*���Qj�<��
=vČZ�\�!]�P�%��p�<�T��2�,�ǅ����ʁ�h�<�Z�����%�IX�0�|�<�䂒�F��j"T�5R�5BRit�<Y@(�Y��Y�	�1>�2����r�<��	�]��i��0�����]m�<����=6u�$��j\��(�㴮R�<����>� ��e��;
�lS��J�<�k��=�<�!��,����NLo�<y-^u��0:��ϓ�hx��nEu�<QsMT�4*0�ѫæ3fh{R��r�<�����a6Bź.���� �Fm�<���V
Ƹ鱵-8{Gne�O�l�<��ޜa�Ľ�B鉰=�F��j�<��h92�,�#B+8�� Rh�<���M.XKp���[2,3�F��f�<� ,S�!�$�Zd�J�PҦ�傖\�<Q�a�(2VF͡GA��TP�T�DU�<A���>q�QH @ ^eqƟE�<� z)�� &'Ȥ@���(U2a��"On��'ɑH��5��$0�d\p"O7B[
 �z�b6.��MN��`w�6D�h�0K��u������8�tM�Ħ'D��s��n#$�@i�[�Xq���O���?Q���?I���?����?A��wٌ)\<p�૓�,6�P\@���?Q��?1���?���?!��?1��>+FDY��Ɍ)�L�k�n̶<�5{���?A���?����?����?���?��/��
F�S�:���w�R>h�2EC��?A��?����?����?���?�h�����Cִ4$k���[1�����?���?���?���?����?���5ЈE�#�K<MT0i�tJ��Y������?9���?���?��?a���?��4XҘ����uL ���T;Q�L�[���?���?9��?Q���?���?	�� ��09U�/*g>����ҋg-�3��?I���?Q���?���?q���?a�[��U�۴	�B�E�JEL����?q��?����?���?���?���%�� ���>L��8����?���?����?����?)��?Q��zUV�G���5K�US�!J������?����?���?����?����?Y�i��5jv�H9]�J���'V�P��?9���?9���?���?!��?�n�n�U%^�|�@J���6��q���?!��?y���?���?���i���'~���h�V�#
P�N�	���<Q����󙟄۴)�$��)Z(t�哹L�*E#��H~"(i�0��s���	�)�P�A��!~?4mj�$6Vd������r7m(?��O�|�)+�$�۠>�X`Vg�O�03A�,��'�RQ��D��B"\o��wB`:��@!���6�l�1O��?�����SI5z�� �&#�3hØ!��Û�?����y\�b>]���ަ��?ނd�.�-��i+[�"ɶ���yR/�O��#��4���Đ�
����F�L�A� N$j}�D�<1O>!��iJ�ӈy#]�m���s�/�}q�h!�i�*0�OZm�'���'d�$�>B�_��P)D��|���C�t~��'ߠ5AŅB���Oߢ1�	�!A",�G�;p�d@T|ң�1��]y��������!k��!.��r�Ju����Z���ɦ�2�(5?q�i��O�)L�d.8r@�)���� �ˎtC���Ot���O����h� ������M�Q�T �"	࣎�i?B@f&IO�<��+��f�9��Ɣ)s|iKG�d�<�K�� ����9	��s�HI�ub��uT�$�rΙ��ɛd��?;Gz�0��M�4Әl	A���Sb�LӲ&U�_��AB���Fq0d
���u=���9~�(ׁA����R�k�!�����j)`�J��avE�w�S
7m��6gD��T��b��f�:p���G]���"�J�=���V,����]\?�M��/�B�<�NL&CY�	������D��]d��\J���X����L�S��U��lȮR}��*ԃ��ܢ䚔�Zxخ�"ƌQ�uc�I��Y2��f,*\��p��], ��)8�B�7e�
�bE�Z1���K��M����/$@��E�jZ6\���ir���P΄9 �f�7[�T�J �Ό �p� �?!���?	�Q��S�� �<@�p�3&d��-��o	�";~R�K��� W+�ٲ� ET�����(O�AJ�	 �IF�aʷL�a�!�	W�S� ���e<����d��t��Ƀ<��A���x�$��MD��%[�-;�Ti�b�j�D?iP����O"�ԟ�	��'���i��"q&�Gp0�y��'�M��Ў%���ǔ3�(���F.���<�H���e9wu0PxfHY3���R(�"R��'�R�'QJ8��'R;�jX1�T">Ɛ3��˯1l>�*��ˢ�p�� zLS  /<O�����!{�Lr�C�t�w���taP˅}R�xW�+<OveP3�'F�Þ �6���*Q�.�>��"��b?��'��I��?�O�Iq�+D�pY�Ő�	D�<�<���'A�9��b�K���˱6��ڙ'И7m�OʓA�2��ּi�b�'�Ӓe�� b7��3l�����7)�0<'����ԟ<�0�ήC@��cmFm~*���`+ֱI?�$���2Z� �r�	�^}IعhPD�?�����((�u;���u;z8y�=ʓ1�1�� �Md�i�T>��d�%%�j�h��V��������?E��'�vLم��&=j4P�gY�$��A4�'�ҵ�`LN�u�p�A�M�/p�|��O���'��y�(�iސ�TOÝ�xqK1"��y�B^�>Z꥙������� HD��y�J�-�����NȰ������!�yb���W6��D�J���AB��yR�^�*��
ꀮ|�vaQ��R%�yR�Ơ
�N���`ҼQ��;�
M5�y"��	'���p-��1�9s��+�y���/V(հ���"dd|b�Θ�y
� �dz��Q�XY8Q�����tF��"O�3��A`�@�Q�TK�B���"O:�P�E�HQ�)y��8��a"O��;�Ȝ.S�vp1A��%��ȅ"O(b&d<N+1Kˆ�[� �"Oh<�qNW�,��с�j؞K��(�"Oz��%%�n,&u*�I�}&�k�"O����W�"���Ks��;dƙ[�"O�00g$� q� �c7�$MQY�"O��OA�:2b�:!KB�rC��:D"O��c�d�e�����)�3t^�B�"Oܥ�ŕ� ;�����9�`:�"O ,	��ؼj�V�cՆA�nR��"O>|�`ˎJ��D��R��5��"O2<����a�\�" �N���j&"OL�@�\wԤ��R�K�,�*�"O��ĮG;
-�	iק�=ɀ�
�"O���
X�=o(��0�>Y%�X�C"OvTQ2��Q�R\Rh�/v��"Ope��ݦI/=�S�H�n��]��"O��L�0�f�HfM�[phi�d"O&x؂��=S p�4���`~���'�Q�@:5Bu��EP��Fe�A���.D��1jT�Rp.�H�t�n��',�<�`@\bI�OQ>Ś�e��6.re(GdF }Oh�%f'D�l��ǁfH�Ba&O�cs:E��*8��\�HG�u�$�'�p�n�N2td�D*�r����{�~���W�?�@Z%(!3R1��W3�V��gT����	C�Z�Ƙ�T�L�B�1RL&#>ae�A�A"����Ӿi�\�8BR?A��02fYR�ʕP��@��=D��Q�k��|h���ȮTu��Bn�0�#ėJ{��HQK���S��S�?�"t���d���Θ�|@tB�	�Cd��@&�[�d����F�ĉ7�Xq9@n�/$"�$J��X8+�N�z��%Fx2��:20�D�a��z��ȄM���>ɀE�>Ic8�!G�aK��R�����27.���u�LȲ!7`�&4�O�D;�D�Nf���qi��/���@���	`�ZsC�к�MʪWq�7=����V��1wY8x �v*�m*�"O�%Y�����H��
��j#�i�p�Zd�F;_	�yG	ӵ��`I�t��5�!ګ#DJ1��#ظ3d��lN��yb.D�b���R��G�o��t0��ʿ4fB�+R�%-|���E\'L��I/�Q�Px1�߀R�"E�tD6�,��7H8�O�� �ҫY���T�L1nFRA�� � i�8j2�����b,dX� ���Z��1 q�
ؑP*� �:��E�GF��Q�&�!{��� ����DȅV�v���!ڒB�I�} �z�IK�Oh0k�l�#Z���	�7������fMv=���J��ȟ"�0#zհ��w��~0bIn�<V�&]$B�B �1#?�iES	 %�`�A�i�@�1b엣�i(͟� �]�E��k�4�` .C�[�r��$�9 �x�A��tjI�R�]�81p��7�;Ĵ9K�oE���	�E���IA�=SZB0��˂6��#>��ɿw��9�cB[(&��|[,�����JQ�&�p'��><<2e��"O"���J62��<S�iD�U-|�#��'`�e!��F�Y�Z�"~7)�]"��1�L��PIW&�yr��0p3���C'�r�l7�� ��DF?z	ح��o�����}�Q�#�<����^�~Wa}�ĝ$}�U�ܴ�RUS�ULz|(fM�#��P������@�4V��zQFD�!� �Dzi��MxdF��d�h���AMت|!s���yB��\���TGM�x�Į�M��#�������Vͅ�d�4���R	:���M���y"��/s�*3��me�����&��d��\��i��/#�0h���Jd�8э�o������{^޼1�;�؅cCC�
�Jq��Y%x��$�ȓ�tيwa<x4p�ꉢz�MFz�`�(/:lĹ��� ~Yx ���jh я�� 8@"O�}��鎖@�T����#W�c6�i�:�����55ɧ���F��.t_t@�7-�C=i��G��y�q7�+���]�h,�0��'��Hv�v���d2LO�-h�/U?ni#w�JN����4�'��-�I�d@fQ3�e�֑ARD���̹8����SZ�<���Ԓz��:���Q[B!�S~rb�["���ꈑ��&���1T k�	�>I��a�R}y�jަe��sI[3`�'s6�*� ľZ����O�3扪?����h�6A .�(r�I E�C���H���z�Ɔ!+R X� ӀAu��{�f�����A�)��	9o�&�7(^�j�Z-3Bf�jR���DP�q�U�'U�!�eȤcz���I�!BQ�%�A|X��Ӣ/P�C��`�G�5Q�d����6?��� +"�	� -  ��i�F<�����+f�(Zw�U"=�!��ï0r����� �H��@Ɓ�\��I�g���B�ҟ�P���N��'
���[�>WE� A�F$[�P=��JY����O�HGY�aޥ|��u�A���O�\ȓ�I禡A�;�>1#�H�`���O>i��cE�D�&��$�J�b%b��O&�a&m�G�2�d�Y�Py�`�� R���I"w����vO���.&MPN�&m���^�$p�ŀ�n~�7	0h�v:�d�+�)��I�R�K��eh�"O�X�6m�DZ���#��=^�CR)�%+S0H�!��Y��?�O�����?��� ?xt�-���R�"�X�6oa���A�&��q�R�":��Ja��(�ް�$~�N\�������;V��qǻ�B�u� _PRX�AŽ6@�(Ѣܢ��"?���
�H��oZ�R��,X�ǚ �M��C	�<��t�-Ctt.�[R	@�h��ɗ\�Z2���	�{ިa�,9Zel�q���R�:� a��(g��O���Ӊ�/T0��'n0|��|��͘S�����F 	��)S�j�n�<�ǢӘ������3a�0eJU+8�:���n~2��y��J0Ri�|λYa������	Kgh%$���*q��I3µ��̂;x����% 
"Qb��DU���v?O�B�'h�h�7��-a��2@Yf��5t��POq��#?ɔ	���dX�:rx��O��5:�g7d��d��fJ�xFT��M�����'*��ؖ+�6�N(����v��us�O<��sJ�<)���U���O^r@���:<M0�P�MS�zw��b�' .�A�V4I��`3�	:��R8$�j�	# p���ϐ ��ɧ��%�b<���6b���_E؟��![QA<ő��V%���*&�Z�pI0���C<)���=�ɍ
����1
����SQ,ҕX�Q�Uh&��<�Z�Č�"��H3��O���K�E&��3`��2�>�������7�a|����hM8������1L�*���Бl \�����1 �T�Y��������8�Ԑ�LWJ�ȡ��yr���hYR����#E\L��.#��kņf�9V�Ք@��0N|�>��!��`U|Ԉ�j͢:��1�Dw��t��4_/¹��)��Z��24H�(�}b�*�+\��a@!�O�̓���%E�"�I�A��J/°ZG�'�0�2S�U8k���,h�"I�e:V�a�B�+d�!�D�)i���{��ƗF���%�ܑm��Od�9�E�&RN"~2Q*C,���9��Y�6�F�1q�O0	x�	<����!�4y#�i3 ��G����G�|�h�U�5~K�j�D_�G�f���E+D�d�0��s�T�e��*>�f��e!j�&�#u��J5�x��ɲ{������. �Q`g�	�},���Jll4�����<��� 4E��q9e܇tP�)y���v�<��)g�^�0GCŋQ"� á�u�U�8��@�����DR��d&(�@P+@p �"O�ˀ��M����O�S%ZX:��i�pX��!#�)��ɫ�IR/2��id��^<��� #D�L�f����ӂ�#k�x�n�>餄G�vTa|���|P�$E�!�4�����>Q�#dx��
�<��Y�b	�h`��+�'�!�䑱$/�l�F�މ'�~i{6��.֑�0���@�����Cf���[��Q���A�*]��"O� |Q��E��
��ya�s x�P�i����V
N�S��M+����*���Q0[�]��*\K�<Aw"((��8�D���^��a��D}��J�|�9
�r� �S*߂%�| #!я�����I�_��A�gӬ��<T�ehk��4f`��"O�����R1[����o�2�*d�2�ɴY�M�u�ӀG�H(��Ս��i�#�c��B��'zk��˥m1���$�$!�6m*y4��>E��4܈���(I>m��ɴ��
5�ȓM�r� %̫�x&I�;ŒM�'��,��� �Ot�j���)<����`�Z�����'�4@U�y��ڇ
�K `0�j_���ȘD�?D�,x)Օ^�x0k,?��@�8�, �=����j�F��CaO�SM���6�X*�~C�ɂ8$����)�/	�zu9��U�UJ7�T5���>E��4~Q��O˱8���*E(֮lJ����N6�3�	=)���G\+HP̗'t$�qd�;�E>p�fYZ��[�t�]�ȓc�!�M)9�Z�
�#�0xvɇȓpVn�����*Ҙ��7��:���	4D�3"�Vz�ԥ�C�64��ȓd8J�f��%J(D8�L�1z�N<��~+$���.�nH�ti0n֩��9��[- �qͥtW��B�פ ��ȓ2��M��� &����Wĺb����~~2a���Ec���Q��v��ȓ-�8%ag��j�<s��,F�H�ȓ^�h[Ԡ�7e�"��AL�	��J�NLp�H�=�f����M��,�ȓN2L�8C����$z�lm ���D�F�1�,	� "��M�Z�p�ȓR5�L��^JK1��95ۂĄȓ�p���74�)�u�J2|#U�ȓv����B�1���K-q��u��u��" cA�X��� @���a�ȓ�]�!O�Q��	�b���/n-���(yb�b qt~�����F3��ȓ=�
��K�k*f�s Ψ
����ȓ)>� @�=���A��NFH��Q¶�ɢ�Kvzr�ЦG���ȓ7�d��$	գy_��B��;5pn�ȓZ�dH��T�?�y4
Ւ����+���pnءl@,��A>kj���Nw6�˗�\R��S)��zu(��U���` �}���2ơ]�e0�y�ȓ|Ӽ��%�����yo� �NZ�<��MO�MrF��2���Xca��M�<y��Q77<8�jĬ�^)�V�]G�<ф}��LX㢉�F�$xyA��@�<1f� �T���R�i�p�=D��ᓀ��S�z�;��4P�<��C/D���A�q|�Y��8� �S/D�`��aV4@��ѰX'{$L�b)D��q�a£@Zl�%��P�&D��y e�B�B�㲩��>!��"D�k�\mD���Eҫs>��)!D��)bÈ�"��A���M�>��Ӣn:D�,�ql��W}�U�a���m��Y�T�8D�lHPL*N�\hRI�Xd��ю:D�X�D�^<.�8���H76�����):D�$`4��ih�Zp�E.\#��;D�$�ah�L ��('�$-)�!�%8D��2�H%V9�Ajb�ܒ�Rq9�h!D����K��p� ���$?�L��?D�� i"�	�M�!n�j�4�A"O�MH�/{�����N�ACb��U"O`U��B��H`F�]L;ԑQ�"O���f��w=��8A$��:f���"O�i$e��(f�`���d�̺�"O�Mp��{Z�%���5%"�ږ"O�u��윐f�>q+5���w�`��"O0�g!
��~|�Ģ80�=Q�"OD���&`�>	O�n=NM �"O�2��Q�UE�d�1���r����"O��A�s�99f&ZS�T�B"Od�X��4!֔!�q"2Lw�T@�"Oȴ��䞓`�B��o��#b"O`�@�rq鑡M�!^�qr�"OVILΩ�T�j"��.q[p�)U"O�I����T��90 �U�+B\1�"OL��B�ޒl����GnVGK�<T"O�p��@�M�|p(�-ِL."}�"O޴bN����e�W'ډ�g"O$(�F��C:�S��.:��@"OjE�쌫+�B4�Q9�v��"O��y��V�]��Q�B��2�\�"OԈ�2��^��F�Vׂً�"O:���MJ�`E�0f:*�����"O��Zb%�.;����r�1c��|a@"O$�{���� �ţ�!'w��0��"O�"eÁ"ؕآ���K��P�"OΙQB+�*#��%j��O@D���"O�Q;����$4��AE�V���""O�U��fX+6LhYc�!�������"O���b"S/"E�M��Ώ����)�"O~�PD�L�F�4Pi׎�R�b��"O"��DMқO�|���Wr�^1x�"Oθ���	�Q���v�!�"O�$pV�(#A��c�b�S!�|��)��`��q�«ˉ��C�*� B�I`ߢm ��� �� ��N�0p�C�U����u�4-����b�-?�B�	�CV-q� �j��T9#��25,�B��0Y!��!�J�f�Q�!��u"LB��*o�I��^�&|��A�f�FB䉛8�di��!n����d�C�oHB��~Z�!Mɕ~v� ��E�C�I$Qʈi��	|��"�۳m��C�I.$�%��#�:� 5	3���S*��F���0���݀D�!�WF�n���j�VHj|��Nq�!��3���iu��6D��тlڢy�!����pf��|C�:5l�d!��{��8��e'T�A���2^-!���~5ҐAJ9��#a�ʹP!�d_�l'z9�%ڪO��9��1"t!���.�4q#B��A@@r����n�!��չ"�|uxb�I��rU��FW�S�!�K�O�t�@�\�t�9b�םwY!�d�64�⽻6��wK��-�*M!�D��q�� �q�KaA\-;�,��<S!���U/���I�k*�e!Ŭ�O8!��Ș(Lr	��HU�S�����Z7!�d�+W�Ч�ʀ!�� �'��+F!���^2Xm���y�~����!�މs��:!�� ?�>�r(:5�!�ʃ/�vԒ�F��*���9��U)i!�dR�՘ͺ&U�Q�����$,�!�� z��Ԋ��q��2�hξ]N�T"Ot$��Q�MG�`+Vh�5=K���"Ot4�A)I�6���ƥ$��X��"Oތhs��0���J���"ON���Q�f���X�Άg]��"O�8��	�fw�ؚV�Ƚfg��ْ"O�GK�	f��Y�5��	b�-�"O�Yk3(�x�IQ�ԅZ�8� "O��3s*��X���R�ρWD�=4"OL�q�-��Y���S��T'���"Oj����KLP�c�n�:0�쀲"O�t
T�� !�Z�cd<�2�"O��%�,Y�2����m�2��"O��H��ڣh�D��"���
��m	&"Oz}�3K�A�ա��$�a�"O� CP�ĥP!�����\�I�"�"O�4�6C�7-J�E���RI�4i��"O8 ��ƌ�H��=:�T3_�ܘ:�"O��j�a�!�v�W�)r�v�"OtZӬ�3	�Dŀ��"K�̈�v"O�1Ƣ[;E�0�+R�A�`�\�Q"O����i��-�e�Ζ �j��"On�9���7x��t  ��5Z唄Q�"Oj(*Sg�=~�� �I�)�x�#!"O�����7�9�Cʏ�.�L�1"O
�j��L��M�5��D���1�*O*�G��}�zɖ�"�@�M>1���	��kh�\�0�]�f��@�$�_�!�ȶ<!���D&ut-�5B͙EN!�G��wU�Zh,y�G�Pc!�$P�Eo���,��� ��oX!��Ie�T�s�e���K�!���J�� K
UD��C�@�)�!�䚵x���U%	�G/�i�P�4�!�DՐP�RT;���>*�%`�..�!�䖖3G�@�i�M����ݐ�!�؛Q��D��J�g�HUљ�!��P�7�i�M�,�]�2���ct!��Q<c����dO>v�V
�Q!�_;P�P�
� �y�PT(�e�!�H�m�u�$���)�yi2�$U�!��3:}�Q)ڣL��4pQ� �
�!�d	w< {unJ�xoR�q3�L(
I!������ɚ=HŐ��@j݁�!�V�������`���#o�;Qe!�DU�l����Bc�1������ L[!��{ 6���n��l�|AGh�*OO!�$�;H�c�'̓�M�40B!򄖕e|����V�ed�U���(!�$���6!��g�'{%�ԛ&�9*�!�R�_���+�(ҒhpLj���G�!���j��9�а*���PRbR	SD!�$��g 2iD��w랁	"��/!�D��P�$���@˴!�%i�
A�o+!�քY[��Tc�(>�n��&�ƕ���)�-���sC셳��ȰAݙL�i��'N��#���;�x0>���'���Ht���c�0�K�3r��k�'����^'9�8���b�4Dh̉�'Ҵ��^��� rf^�-&2A)�'���{Р�;nF�Q��|���'*�YR�ȉ�J�|8��A�{Ĵ��'��Zbꇚ*�RjΨ}�9�'� �
#	؊]����,�I���
��� >�RF�S�]�����ڰ}���ZR"O����$V���!ᆘ0p�ɪ�"On�zTL�)o���)ǲMcD�R�"O|i�m� M�<�����Q�2)��"O�1q��;_��`b���7V	HEC"Ox�X����>�h3�@��!�$�4p��M0tȑ'.hLe!�Ą+e!���;v��������=�>dt�C�I�!�d�_Oࠐ�ώIndQ+u分:�!���h8�� �S!rB$y�p�W�2!�o�����"Ɖ(Yl��DZ8�!�_�g�򹊤�݂c�^,�b�D�@]!�dȳ,p&ؒ�h�#,��M��㚌CG!���-1�!�E���G�ν`!�$�;ys��S- ?�E�r�A'
c!�$��3��U(QE��x����FC!�$�3�L��Si�ؽ3�j�.O�!��,uQ��ª�79�4���"82!�DEвq�P��T��=	�惊�!�D�  ������(����R��C�!�$������;n��=��N21�!��j,&|�����D"�L��-�!��#��T��	 Zr��#�UKr!��@�A�����	 '�F@H��S:6!��V�-�T�1��I�W��̡ `�&E!�J:Z�X��Q�F	� ��!��8r�W��-,h�a���<\!�\�u:1!�폺BImPхg��"O��I���Q��]�!�ԑBGx��"Of��`Oɋ`��E2��
�,*
��"O���w��d��5��o�>5�jȐ"O�X�����qb�]D��"O����bS�	D>�U'�;3Ҍ��R"Of��B[�P`�Ч�$uμ���"OV�@%+�V��IX�Uʺ�s�"OXc�ϓ3m��as+��zh�F"O`
f��� $�����RK�y)�"O��rFb
��*���m܉u���P"O��p�C
~W�8Mg4BT�"Ox٨���0M����Z��<q"O<T�R�f�*tR��Sp�h��"O�!p0��%�B��R�Y�	�1"O�1"��A��d���ĥQ�"O�����ZK��t���F���pV"O� yf��W�Xq���#��R�^�!�Z�]l���PcH/e���`I��u!�$Ij������9�DP�h�	b_!�T�i$�ve�2���h_jM!��@���q5�a�H�!��^L!򄄔?�����C�]6nT<1!�DO�
�p��w��H0��:�l
L=!��-*\k�e���b��\f0!�D��|�� ��?����"#,!�D˭b,t!�O�K�8�`Ë!1!�D�.Q��0���X��Y�s��g$!򤕧Ff���i�:�v��r��`!��[�2�Dб'"a���B��Ռj�!�$@;=@�J���[��!T����!��	��Z�!
Q�"t��J9I�!�����]�FCHxh�j�L�!��\.\�(���@iz9Qʇ�!�dM�`�z`[%��:Ailp��)��(�!��^,G�t#̹'E�u�bOI$;�!�	�=CzHyAE� ]H��� �<^!�� ڠ���ݍo�nU�����r�Y�"O��HЈS�Wb�{�Cӹ:����"O�� ��� ��+e#�䶹r"O�x�T.�&C�2���+#�@�j "O���vA��pq�u��$p0"O� ���ΕE��I5@�Q@xt�V"O.z�I�J�r�شNZ [3�ab"O�(�a�P�xYjl$ZCBى�"Od ���4[D���
�w/��s"O���K�	;{�*�1�@�"OVM��/)b�E:G)ǯi���6"Op����K�t1��	[)�c"Oz�8�dRF�|��`@�5JҰPF"O(��1D�aI捂b�?t�D)q"O֤� �~*���W
���A"O8���B
Y��e�I� [|��"O��C�j]>%^)jU�}��%�T"OF�D��R�`H����6�yBZ��P��$���E��Xd[��yB-���GE�=cT5r��~�<ɃJM�J2F�s�.@����WfWE�<Q��fn�ꡪ�H��-J���{�<�Ф�� ��a��R˼�	��w�<���E�r�x; ��a���`�M�<Y�����{�$�F�<DC��I�<���ɸ@�m���jx0s�H
H�<qfIñ}��]�� e%� ����_�<�3½OG��r�^�W�Ԙ(�d�<�����DP`��k���K��a�<q���	B/�(��I^�0�	MF�<AP�]�H?L��3�PN�<��T��\�<�0HB"U�lM
�^���Q#�Q�<YP�R8aSV)[�@��#H}��-�f�<Ѵ��'����#@�K�B]X3IIw�<YըʇE��a�el�/'d��� N�<U�^ �u���͑��*�DEJ�<A5�]B�<s�oWa�0�#���}<�x�� "��@�J�̇ȓ��1���RYs�9�)V�VI:��ȓiD�$RЊٞ-�vT{�% H��i�ȓ s��u�T��(�砗`1Fm���T٠��P��l��������a6�X��ש_$�PKb�Ƒ?H��ȓ!~T�k�W[���c���0���By�PH*Z7������w����ȓ9�^��J�+�D�0ՎO�;�0��=, Л���s�8h��P����d �L�<��U�կǄy���ȓU`�p"ƬX�k������ ���9��Uh�i���5����b��j�=�ȓwg~���#9��!�DNJ�_����'�0WM�*���
T$L9)qŇȓ]Tv�a�㉒Y��ab��"D��"OPx	JO!�����ߓFaB��Q"O���j�2H��U��	͏
m�䢳"OάH�+� ��ܪe��c^@-qE"O�ᧂ8bE��5fG�U�V"O���f��(=���a�%.&�"O"1zT��fuv�Y4�Ȓ'?�r�"O�I��F��[��i[���4")9�"OJ�ڤ�
VG�A�b�[f���"O�@�!a�gK���CM�"��"O�DHaC��b$�m����[��A0"O�eHR�O+}��m�Qႝ8*:I)�"O� ��iZ�vz���f�2_&��ږ"O� W痾=���]�:��(�"O�����)uj�@���;~��"�"O 9�D�0]�eߡ;��{�"O���ҭX���*�A��0�\x�"OlRd�ӥP�J �I�7H��2"O�x��Ι�pj�3O@%a�*<ڳ"O��p�ꇎExX)a�M� 1�����"O
��d׷	ڦ]��ؕ4�&��r"Oha��.S)u�0w�#">�)`"O��7���e���KP�<�mZ�"O��c�.Ϛ=�<���\6k�P��"OF�J�L�[�.t�T(5 �}*'"O��V&L�
N1�H�s���s"O�9��-�9-OB�h7�U? � ��"O��Y�Aߖ�`����"Ae(8��"O�a1����1��mi��U@T�	"O��J���&�l�:�B�lLhp�"O�tP�T<. ��r�y�Q�"O�c#�$Dx�u�� Ի:�Fl"Ot�%�45����4b�6ђ�"Op���Ң`<h�Q�֬P�"h`E"O 8��P�LK��GeĒ)�L�@"O�)D�"�UJsj
,�uY�"O��A�*^�4��5,��~�P�"O18g�#ϔ91�R�y����"OtSd�Q�ܕ��!���eA�"O�SUg�jv���ǁ
݊��V"OƘ¤��AaD�M?/��@�"O�����ӾM��R�Aمj�¥"OL��D�xN���f��I�`I�c"O�X!'�P9#1���/ڙu<;�"O����0V�|m	�L��[�"O�� �	�j�U��N©}�$$��"O4��f���fe��!���9q��&D�������Y�d+%̚)HrMpW�%D��8�k��p��T�;T�q�3%)D��9�� ?��Y��GI�fl~i�Q�%D��K�	JI�Is�)F�Zz]c��&D�غ� ,��p�B�<�<��v�)D�<1�$'��+�4iO�y��(D���!m��l��uD�r#�P��-+D���/�*�=�s�$D���G5D�ti��I�}_�D���s�<�vK2D�Jׅ��D�\0�烔�MɔH��<D����+Ug���Z֫�.Q�B�R5%;D�����3f?)bȒ�WTpT��G5D��V�9�Xdfѧ�|@Q�F7D�<�`EQ��B�-*@���wsx\�ȓC堨�	_���@@�	@���h��R��Z��ϑA��"��'P$��ȓP,�����05��e5)��Du�8��'X�� -B5��U'�1�ȓ_���wލ-�n����:�d�ȓp0�t��!�/7|DE)���7��Me\� @��5�%a��4gp��ȓRj����ʅ�<)u���0l��X*�eH3爑R[�����o�HȆ�o����p�_���5"��fb ݆ʓ�FA󦌾.�LDK"��Y
4C�4�t!�ɀ�z�fPx�-�t$�B�	tL@᦮�D�z� #�${�B�ɶ@J���d�]' Ղ�IS0�BC�x��1�`�8�N��0����C�)� `��E�؀"�"%�' �1
1�U f"O@��~���c�*.4A"OP-�!�-N��Q3�I!:*� �"O�kuEJ���ѫX T@�@��"O���D�$ͤA
F(��(�"O�h	� �.+��C��8���"O�0:��Ճ3'�Q�g%��a�*�2"ObmI�b�e}($2�#�� ����w"O��҄扃\���Q#ٯ"N��D"O�uip/�1u�0Բ�dY*S/���"OrQ��i\�cŃ�(��"ODY(�C�	.l��-<���6"O�Y�&�Vb�!��>%C@���"O~}����$H��� �Z!T2�`�"O`;��Y����BS� ?�y)�"OZ����B��a���NLTE[�"O�Xaq�J�e<�)���Rv���yR���>�t���۬qv.1�����y���8d�����NN�U�p��Gj��y��6J�p�A���#`���I�ɍ��y���0)�Աis�k,�2��[��y�O4����0Z��v�-�y(Ϫ6.�����ڭUʜ��y���NP����[���Q霂�y2n��{:j�EG[�<=xf���y�J�tir��1@�t�"��"���y2$�6.��(krIQ	n\&�C����yH��i!h�x�# f�1c��yBl>k��p�D5 ֑���0�yb�!:�@��U��
+�v5bM��y�*U6\P��x�-M?"��['�ɾ�yb(�),0��(����u���y�M6!�r��r闐��`Hډ�y��/r�|KT���
����&��y��&d�����5�����#^(�yr�E�1�"��%�Ԟ1Z8�J�D��y[�~�F0(�}���:� 	�Py¯�5,q��ₛ>N�@���c�<����m#���QF�K�
�k�s�<b?y�STB��2�p��0p�<Y$�� kt��JC�%}2!9���P�<qt�H�V������U�AAH���Wd�<�anB<C��IX�mN�F�!�FNQX�<Y�g��%06��S
!=p����W�<Y�_**~@fȆ��0�
�Z�<yS@V:c(H᪑���~�R�C}�<���ܮE_\L:��] �� *�n�<�񠒠*�Tx"f�X�zL���F��C�<9Wg�%1�� ���l�l	׊�x�<Q"G��3u8 ��ݫ9KT%��#�Z�<1W��Gf���HS�7e��9$��U�<���fT��'��/y����G[�<�PΛ�^(.pS,V�pC*�jR[�<�2�3�����	����R�n�<��㟏<��Qs�e��F�@��sΕ@�<i�͒%ov�8ȱ匰]������
V�<�TBŗ�°l�!J�c�S�<ك.ߝd��9G�Y*�Q�dM�<�G�C4©B6AX�j:0}iҊNP�<iu�O<D�-a��3V�!���AO�<!��<�ڀ�f�0{��8�'H�<����Z�^iI�
�> s	�y�<��팏l��y!l�"x]�0��s�<QU픆jC�q�-!8�����u�<� �)3�� A�}3�@�+;4��"O�A#�S6N�Z�{W���O�p=#�"O�(p��#�*�H��$��%"O��v�L
6SD rG'��]��"O,L���I�#`�A�FΆ ��"O*5���u�2P�T*��̥qT"O�1�a�D/)�x���h��de��"Od"��1b󨕛D�Ǝ=�V8��"O��Q��+��ě4��8͎�`"O��FGW7	j�U#G�:c�x�5"O�d����(�$rUܢL���R"O�um�u+R�c��ܝ""Oh�A�N�a��Yamˊ#�x5"OZ��u#E2����5�!��A�"O$iBjע�X��#��8m�f��"O�h����=��b���X��"O�-QW�7dV,�����R�"O��K���4H�l�3�ݱW��$!�"O�����5�
U��NN�5bt"O������J
x�A-՗r|��"O�8�6ME�J��t���Z]���3U"O �HЏRX��t�E�g�8��"O�stJқZ#�A	��S
;�L�	�"O�q�	�X�p���]c7"On�x��_7 ǆ8�Ba�O0֗��y���c� �F��-+ "�����d���[��)9�yk����مȓ#?�ysc��MgF��6��?-=l�ȓ�2̻�.��( ����J�CJ���7,���W��/P�@ͻ3�@6y����<�6aQC�\%BT�ۧꐲqz�Ņ���y��+�z�iX��PQN!��A��D-�	q<�]�R��SY���V���l�|�<X��؍uR�ȓ- ��@$��z���$@H�z2���84 �� ]	���mX8��p�ȓy�Ԥ;7# }�H�Y�T
>V)��?�B�Jp�ȜV	�1ʖ�sHn���k�@A��jQ�g��#OB&�4��&P��PD��R�NG�E��%��gp�y�"��+	�����.�,y��ȓ6���ƕ'id���3c¯=��u�ȓz��Q+��ՐY��}p���
����($�L��ˡ$� ���D�,��ȓZ�)��=|f��P�;�Hԇȓ(���0@A�t���aߤF�}�ȓz6��Q��P�r(�L�����ȓ��@��'6���s�H
TsҔ��/���Y ���X@��d�P��+��E����&y�X遨��;��A�ȓa\�}y�i��=ffl�1aA��m�ȓq���7&�)6 �P�̒8yW�-�ȓLiH�ˀ��^\�5�LK��b���mI$���˖�f��
N	>����8�As�E6$	�X0���6ل�ȓ`<ıXF(^�z2��!1b��,��ȓ:��$j�n0:T�q�@ĩ@&Q�ȓz��y:_h��T�>R�1Bw�K@�<� ��AJ��C��2 �} �O@�<qs�įa���@�G2(��ux�ʂ~�<YD��bxr}	C�׉	;$ �_�<��H��P�"�� %���q��X�<ѳ%2w�e�Ҋޥ�eC�R�<���O%,�� �!3戙N�<� ������/}x�Y�"��b�l���"O\��׉U��)1F� ���J#"OR��Ҿ$��e�3��Q�^�"O���g�5rS�h�(�0�#"O�-�)�K��h[�lŏ}�`��"O��[��G��"��Q+�9Kw`�bF"Ott��A
S����l�(�h��@"O	��Y�4g*8��뛑
fH �"O4�B2�� F��J�
̝��P�"Or5k�n�!-��̛�IQ�[���	C"O�([�f��G�i��h?��B�"O�0���F�Bu���޸kJ�)�A"O�ࡗ��$�L���W�Y<�,1�"O�)���[�рJ+m$���"O���7���Y���ge�H-p'"O�@�f���������q��s!"O&<:!��7[L1#�J��h��"O�@�+�)rː��ꋼC�"*�"Ov�F�,/]�p�T���
Z���D"O�PaU�5�4h��
PJ�"O��� �~�r���5�"O����ӪBH�z��Ї_	�-['"O�`*�DJ>yÂ�܎5�v�8�"O�qJB��f�6�� ��X��5��"O��eB]�gg���c�(5cN ��"O��beJD 6i�0k�D�D�"O!Ԅ͍d ���
I2A��"O�йcGFp!d���֏^��B"O�� ����0����YvX�S"Oޭ��U3����ƊU���c"O����
��,_�xAjS!��\��"O���1c�>1`���կX=T�{"OB��\+rS��dΒ7]"���"OPQ3!ԼF�l��U�?��]2 "Oި���E-v�
�F�Md,���"Or冈$�6�Kӌ�M����"O���kq-�St�^�G�9Ѡ"O��Ȱ'��h\D��$ ��M��"O�I�E��6%��-�ю�#8���$"O~��G���$f\yq�l��#"O*��o r���4�&kzd��"O�P�T�EH�͡cʅ�wm��l2D��0���?q�0��쓬?wXj�!D�кG*��h5���Ԋש>��-j3h?D�T���F)��0)��_�T�ȥ�'&=D�|2d�B��h��@$.�N�1�:D�$��$>9}.��dǱ6(PݹD�4D��`"�Z��iLS�I�0I��0D�l�0%�<5�t�B�h��Ȧ�)D�4t�ã6|2��ԉk���A�&D�@;�jE�E�ܭ��!� e��A!�"D�YO�&w�:�"֑�օ�WM D�ѭ��5���0����ɋ��"D��2"�̚��7���)S
A�<1�n�=7���)Z�vIp�G��Q�<��@�S������T&�b��s�<�JU3-���+1�G�mذ)E�z�<	�!�aٖ�`�i�"(�z�<	d@�v���!�<'�j�ih�u�<� T1bG�T��oڶj��	u�Su�<�A�ȑu>��AK�Ff$D	7�n�<ys	�{+��Ç�U;"H�xJդTm�<1���,&�b�%7p+��7�Po�<�c�s BsSaIOt��Lh�<�  I�F��_��`��6B�����"O�����M{ZnBB%�0p&Ψ�`"OL�'L� )���$BB\�"O�<B�K1ж����	%p!�U"ON	v��<(b1q�BW���"O��26��Oܾ$�\#k����`"Oƅ���23�U�$Ճl�P�ʧ"O��ôD/IL� �Ë��DT�w"OD��&G�)ܲ�S�c̶`���y2"Oz�{1d�-<4�Z�b�]�&�K!"O��;�'�X��1���~�04�"O��EݮZ�)P�ǉ4�:pY�"Or}C��W-?����G��1o�>|��"O�}�����Km����dU�Po ��"O�U��.ٚzD�h�#c��a<rv"ODD���,o;�̃���x����F"OF1`ӫQ�N�8$� 2��z7"O�e7t9��R+N��mu��F�!�d� R�Az�H�u(��a#��D�!�	h��,�Dg�^*b����Z�t�!�K��J��ĉ	�T�C܃	!�dϞ
:�5�ÁL�3��JR�X�!��K�-���B �w�� mπu�!�Ўe�nۢ�A�1�x�	��!�$C'j��E�%էa�F�Y��6�!�$(H֘��ĀQaɇ�!����'v�qӧ�ǩp�Ŋ�&�z�`�'Y�\B\p����(�@r���'��L1��� �`Ԁ�1�^4+�'6> ��c�`�����
$��=�'� [�M�Hefi��RJ��'g0$��S��0a�(�*h@��'�^a� K��:@ex̏
�>�+�'�v ��]3d�ɠ!�M�5�p���'8��[BO�;=|��A1�I]q\���'wL��r�K ��h:A+ΓT�JP�	�'�8�z�i�!��K��R�f�@�<���S��p�C�6u��ӣD�<�( %("�T�Q�������WF�V�<��S�?�\�R͂�(�$9Ǥ@^�<�'�6D#"�H���\�B���V�<����7�P���a��:��ұ��R�<Ip�U�S���P,&�	���O�<�dᄐ /�����ż2��D�֯Q�<����P�0E�#oL�]���0+Dh�<Y�푒nPF��f
ͷ#o�gh�<$&Y�0�V���H�6L�`�<	���v�\q�E�2A�!�r��^�<����X�2}��H1t�`Z5��v�<�s)L�h)VU;QdG-i/l�Y'��u�<��cC�i�,9�QAH'Q�ܑ1��v�<���	��@՘#!&��1х�h�<!��S�p�����hW�J
��xӈ�g�<)3��"���r�_L>��& _g�<ᧉ�����%���T�$x!�`�<�ꂍqh��[ҭ�0-X�l�!e�<��INP���eƬa\A9��G�<�TER$\�5�f@�'d.4P����k�<Q�hJ�a28P���`B�����Mj�<��l��R4а�r��U3�`�c�<9�C��&��D��ĸ?���I�k�]�<��iS�3�4|��Q*h3n}A �s�<i�kȈ}�6�0��V�J��hIGCX[�<1-E�L����EC�QD��g��Y�<� xi	�b��IQDAB�Ez9��"Ov�!kD��0��$�Ыa�b2b"O@�{RdR�n�"���M]�zx�Q"O��I��[$��s%�E�Gj�t"O"����7\]��#1U���E"O���aBiހ�Q�e�'Cb%��"O.�W��"���rY�.4qX�"Oze�I�[FB���.d��"O��ɀYڮ��G�Y�Bԡ#�"O� �-z�^�`�}�*p"O�e#�� cP�q�*�S_���"O�@���2�LPZ��U:{�j	�"O,��8?`ؠ��=sڔxre"O̽s��o�J9!m�р�R�"O��F�Znx���k�Ԉ�"O�a��$oǪ͘1 �2p8<�9�"O21���
h���o�2X��"OP]@b��
��l�G!�-W�M��"O���SaC
a��I2�҅U6t��"OΜ�5NՆ�ڝq�L�V'�Y�"O���E�F���:� P!.�����"O>�#㫝�+����	�b�0	��"O�L�#,u�E@&�D5T��@A&"O���u&�px�t2W���y�f"OP1��A^s^)�ө�tJ88a�"O��R6�۩!%v�ʣ�I#ybإ�"O�����/T� �J�:
]rU�Q"O�� cf����)��G,��"O�a ,&q2&)ȠiyGj���"O8�D�� j����u�F�`S"O�*׍يH"L����d��M�u"O��e�����Q�JS��L�1"O������8��UQ���Z�ڼ:�"Or����I2)X4�Q�R(��"O���/ 
"9�衣ϣ\��`�"O,z'}l݊�m��"��-:4"OJU�ǯĪ`%@���+}�9"O��1���yUj��Ujq[� �w"OJP���f2| Z��4#0ր!�"O�u���L�&"��Ã�@�(:ԻP"O��%��4����E.�*�2��p"O�����ԌYݶE�欁	{�M�p"O�:�GJ�K�>|1��5J��tQE"O�	���T�;l� �+�|2�Q'"O6i�W
6EeĕZJA01���"O^XkP�:���Kj�=���""O��)Sc��+݂�i��c�� �R"O��5.Uy���(�G�MP�"O%P�Ƴ����|,6� "O �z�V��J�
%��,�Q"O�mů� ?ц�Q���3�5�4"O��Ag�9��(چ)�2j�Հ�"O����VY�)+����@i�a"O�EiEJ�1s�x�oa�f��0"O4YG��L��z A�Wj��2V"O&��L�k�ve�J FD��2"O�i��-TRN��i��,�x�HP"Ol����?H�|�z�gې9��Q�"Ol�:"iK��̽;�Ƅ�}$��2'"O�X��[9M��EҠ��4p�"O�tpBߙR���3D	�鼐��"O�P�s�Ğ�<�&�O�z�� �"O�0�p���G��Y��E�gm �"O\�!���,�J0��TN��@�"O� 2�J�@��B|�ї)D�\`�"O��9�$�;LH�kQ� >��H� "O �T,��CL�d6
+�$�+�"OXDS�e��s[>(zҎ��
�Z��S"O$���+�&*ǂ�#��+~Gf劔"O��D�B?{�	�fK�c.>�Zt"O����/�^���c�K�o�V��"Oh��U*͎}�
T��C�-���8"Ox����9��������)���1�"O���Mr�69��������*A"O>L��I2h�����+�QHB"O�|��-�P�L	�B��A<��v"O6�K�"Nl����'�O�x,|i�"O�A:��I<���S:v����"O�q3�]��C�H[5$�̱�"O��q�#��.���g�P��|:�"O
��V�"I��: ,�&dC��"O�Kp��X����+G�,���"O��:���i{�u�F��P��x�"OLM���I�2R@�h`V
R�DaC"O�-8�{ܨ�1���U�L��2"OX��#)]��p)�CC��s�"Or��M^�xZ��"��i�ڐ*@"O�t+#cQ=���N<Tp2D"O�*qj�9/��+� Ѳ/4-b�"O���P��RC�m�Q�m�̉y"O k Dޕ�Zy�`�H��\x"OvD��,J�1l�x1�G� v0ܱ�"O�Y�s5
�*t����� "Oѩ�!9��Tn�;:��ڑ
;D�|1�i�4u����9[�|X���8D�̠C���R���Q%�&0h�Y��5D�$��cG"K���z�G���J$ 5D��³�4
���[��D�0�qʖO3D�(����#�,�����#A�A�3�+D�T�S�\�Q��^�L1�u���<D��ag̈́�PEr��0!��!s���u�9D��R+�)�`���M@�Q�C�2D��:%Eg�!��?C�V��<D�P��=�.M�'Ý^��[��9D�D(n�	T�d��1(޴x�U�7�7D�`P��Cc����]"2Nv���c6D�dFM���(d�������3D�dxt�A?dֈ#V(V�~��L%D�<(�CطE�L� ���p�k�'D��Aq.�k:lu�T�N�J�h�A*D���s�YD��t�M(�,��!.D�X0V�רKjX�AlJ�)�$���,D���pCB#S@0����6~V1���*D���ŉ F
d�$;�*Y�m)D��s�@�e��p6�M"/0��`�3D�<�cL�>�N��&��L�e'3D�� ��_�L1���#Hr���j%D���C`J�I�`��fڨ6�9��!D��2�J�nD|�be��{�l�A`?D�\��GT�Y�����&��g�R���<D��CFiR01$��Ӯ>X�<��J9D�T��ĝs`�Y�o�8"i�|!-D�,���"6JXy"�E�11�l��o+D�"�i�%���%�l��@1%�.D��B�%��@ �'�<L�r�@�8D�T�CcM�F�L��1	<���'+D�������1RL]IE�ì}�ֹ�'D���1��<d�Zt9�L��w0��9� D�� F�p�O�#�Lx�T�V�b�m�"OlP�,�j�<���J9e��ա "OZ���LG6:���ѩ�++�� ��"O�9B��R��{�P?)��a��"O<|�1�\�}j����-����=3�"O��M>T˄]p-V! ��] ""O
!���уY=|/��҇�f�!���J�I� ��f����G�	!��W�E����0�·^U�lq��(�!�Dߨc�,x���
SDE"����P!��OL�yP�bN�tEb`�� 9�!��JE��0x\× ǣ8����� Z�}���;sj>p�v��#nY|��ȓe��3Eo�n��J;J,��n�s�<!�˖�es&AKd�X�+�x%r lX[�<Yç}F�xsre�O�n��%U�<ٰO�KJ��P�C�XA���l�<�t_6j��L�2����2r�Tf�<��`�R�1�|'������J�<	�!�`��)��(N�]5 ��bSC�<i�	k0�IP�R$f!�l�ok�<��aL�A�U��RuE�T�[�<і��~�� "B@�iт�pe	W�<1��"n�d�AT'�Zi���}�<y���;���J���RC�R�<!aiɍe�8�2��zZ����W�<)&˕#;��)Pː+J���2�SO�<C�>O�,  
̣X#"��T��J�<�P�C�c}8!�Y	u"�Q�)M�<y���Ü�"_�Z�\̲f$D�<�c�G(9|��#�R=�I(�|�<3g�u�����		�d���Uu�<aC�~�*,!�c\b{���b%s�<aak�.j�$*�Iφ1�~�kUNz�<��څ|MT��3�9O|�8ra��Q�<Y  H3:(��ô�4^h���-�N�<�O\�L�\���N6P�����IH�<Y�l�t�����f"���A^�<��V)����b�,"�ป���b�<a����i��f��Pv�A��Z�<Ʌ�3
��(��#A�7\pD2�KW�<�'�+�H�?�Zt��� +W!��+�t��"�+��i#u�]�!�dR>6g�"qG_� �*x�� �	i!�ρN�P�u���3y�V�P$!�d��x:|����@ =�L�8�!��[�K�f�s�Mc'�����Y4�!�Ă9ˠ�vO�2k�6�QOR@�!�]7,ޢ +6!��0L�r'�)�!�dEb�@qV��(B���:��J&y�!�!n��ř	SJ��fK�w�!�$Kl����7��c���冗Q9!�Đi�&ɂ��J��������!��ׇp�H�)�f�(��Oз,!��/,�D� D�)�]#Ӎ�;0!���)��$���R�='v�W��V{!�D�4}�V��7�Q�t8�������V!����e�6B*�D�"P!�	9*��"�M~P8�I�!�D�+1��e��▜p/�͐���4!� +jW����� �t����kY1!�d�+�l�r��؟5�H0�W�^(S�!�dJz�4d�� xBl�	
Y!�;,X�B��Ű}��鑳M�ka!�� �53�lO[v����-\�F�4Ƀ�"O��0���dC`����Ը����S"O�9� #�P�z}�!�����̸�"O~�2���?j�x�i=yQjA8�"O��yv� 	p�G�qK1"Or��0�B�$����}��1�"O��eN�sˆJ`��/v�Zl�G"O&Ai�i�d80�U,�S�Q�"O���)Y�=��U#�,M�~<��P"O�;#�Zh��ak.V���a"O���Z�˲ă\w�A�"O^��	+g�]r�#ݲ{�`])W"OX���φ���������҆"O�A�󂖾OF�!P���cT��sP"O�p�A�?:�q���� .e����"O\h��Ņ�Cn@�{� 2\TLa"O�T �aȄѦ)��Q��m��"O��cA�N#M~Z�(�-ϊ\4���"O�$��"�����M�N<AQ""O��ӡf�-3X\�#�J�q�͡W"Ox���οL��i�#�;eߤ@�@"O���eo�Ğ�o�*`��$	"OT�Ӄ�u�ȱcg؎f�By"O�$·=�E��,�&Q���k*O�P�`H�>(�����5fEH\{�'�4�fW ]�䀁��K2[B2aR�'�P�ق!T$�TZr玳]b��r�'�L ���Ǝ?x�81�0%��0
�'9�2��#7 QK�%L��8��'��H
�m��	�xIի�	�nM��'��H5/�+�P���(X� ��S	�'���b+=��<��)C�K	�4��'#4L�#���eC�`(u ֧1��@��'����dG	�Zg3�f[�'(�e��'����td�cۦ�;�nM,�@E#	�'�Z�EoQI!vQy��_�G[���'H�sF��vĚ�*�6J��	y�'� qL\0�Ι�֍ǽ@,!p	�'�l���',�$sF.��8�l��'F�=krD��|��@	
4�����'�te��P�g�E�,�}	�'���іK�(�ܬ��c�Mm"��'�5�э���f= S�S�	�ũ�'��GO�l|���[	g Ћ�'8 M � l����r�@�~���'f�U9!��P�Ԩ�C&|R:)q�'.p,�κ�Z��@
�wW���'�t,�Qf�Lvlc�ǥ8�A3�'{ν`�Dֵ�4��,^�f�j!�'��{�q>���L��c���
�'BnM��A�,�̴��,q����'�<�AP��$�XI�m�%^z@i�'����K	6�6lPTƙ�U�a
�'�b�C�̯��@��K�I'���'M �ec� xh<w�^I��Q�'�V�P ��6Nה���dU5C��k�'����m�
87PлT	[	.%�L��'�xe�TقצA	��͢nPV��'�V�9��JH4s�е4^
�;�'ؒ݁��.
�j8Ӳk
�1�&�!�'�:3�kG7:v�����Y�F���'P�z�σ�OOt��a�^�|�m�
�'�R�p��_�)�dqрv� ��
�'>��R�,&M�i �*�n��4���� 0���Ϛ8�h���R�����"O4��CDɈW�����E�fئ��b"Or�C"��.��"��]f�$h��"O&��$a��o�TdX5ᓴia����"O��Z���#�6�: �M�T��"OL���f]--��k#���U::I��"O^0R��@�_?������2P"�p"Ov� ��߯T�ڀS�1O�z�"Oj�+�J�X1���7��ճu"O�(J���,|b$�r�ʚ�u�ŋ�"O�P!S�
6r�x,\*8*14"O2$�+]8g����:IA�y�"O*h�C��(XȤM�`�'R\�'"O�ع��F�a�(ưJXb%�j�<Q�j:/"�����%����i�<6�=9=��4c�	#�Ȋ�f�<yAȜJ�q���-����T��f�<�1%�3\u��/nB��"˅a�<� ��%D���ᆭ�+���DW�<Q��A�,�e!����(`�	^�<��&rp-�FT��(0�F�U�<A�o��K��t�	 ���	���(D��r� �1F*�C�JF��5#�&D��Q5�� N-<�CH�&7r)�f D��Z��SO�I���3&t��A:D��+�:o�P�ac�.n.>4rC�9D��s���';^D���B hH�1�;D��3���.i�$���L�"�"]��8D�dH�mMg��� z6Ub��"D��a��h�<�p�M�xT
�r D�0�e��}.�ˣD�)U�����>D����@2Ȅ���zV��#g�=D� ��#YZ�2A(�/�92l�$r'/:D�d�&&K���2V*����@"D��G���s:$+�'lG��Qp+"D����2\:�pا�L��H���!D�`�5���F�X�O/$�4� D�H�,N�L7Ҥ���OO��x�p>D�\�aχ(d�z�@�9c��`�(D�����
��B�j�-��i%'%D�|�JB��7CƜ"ܒ�J�MX3�y��\�ZHh�V$!��wJC:�yB���T�d��a�-���� (�y��"9�L��BP�r�J��ٗ�y2+�(y����E�^t��E���yB��h��5�@�I�ʄ ���E��yr�C;hY Sa�>&�"I��y�T�c��Ss���
�c���y��ػ-\�,3II�z��*�F���y��=|h��Bg�Y9~�����ʺ�yreX��ed��r]�������yr�E�������q���ˁ����y/�}��Ćz�|)����y��F6k�3#�rGP�I�	G�y���H�ň�����K�V���'n�Veǡ�@YFO؊�����'�d�"L�|�ȡ��f�+�Q��'��	��* (dB���Ҡ*����'�hc�WY��;3h�/�����'���� �J<@�I"��	�'�X�+�%�M�dE(�(т�.��'��;u�RGrؠ�
�'{����'y�A�b`��U�Pk���5`� !�'b^�!/K7Af� ��B�n���� f��BbNA����A�2�
��"O�	��S�b: Xt��Xp"O�Y���O�_�B���E7!z��A"Of�Z�0=YF �R�I5.j�6"O���Z�[�,� �_"<D��"OzA:� m���S���Q���"Oڅ��A��W�&�X%Ms[^�3�"O܈yB�؁ _�0tЏJ��pv"O�\J"a�0��\	7�UX0��S"O��a��&���Y���v@��"Ox��tBBV�����zIHB�"O-���A�R�� �u�ܳ/:h��"O���3nY7�"��G%��Cf"O�-Bd�H�5d89�F[�����"O(�� m�)}�8b�%�f�-a"O`X�I�J��5���|Fm`#"O��3bdզ5�D��Qc�|��"O�^%�����V�N�\tp!�MD�<��
N�q�>�C�i��3�Nyku��z�<�%�?����M9f]�`�`�<���XG����Լ4)N��Ua�[�<	��٭���9� �X���"�cX�<�l�M���
%�s�J�b��}�<�s�̯4�@Mq�G_�R�8tz�� |�<��H�5�$��
3�HtԌ�t�<I�@�#=�	 �/��(`��s�<dkL�t9�y�V�ʷR�x�t��m�<����3.0@ᢥJ�m��ILQl�<a`��&�.����b (���,�i�<!��kDR��!Z}t�ثcϑA�<i��Ɖk�к���	4ޠ�PE�A�<��*Q!�Mӧ�F�@�j���~�<i���s��Q�H��2"$�P�<	��P)\� �G�'x���P�<��nlj,@��"T�2@M�w�<����t�X�� 
uh�\���[�<���(}"���1�K��Tȧ'ES�<�Ճ�%�Z� ��z����2L�<I��:�$����\�N�F�Q��F�<��A@�C7�M�&Y�uR�U�$�K}�<���"N�4a`����pc�{�<�sMC.y1z���,E	?8�A��DN�<F��
���bO�#Ŷh�@�V�<�4唹dh�k@j�&(��ah�QO�<1":
�A�"�dL�C�M�<�By`8X�6)8]2�*@��o�<�U�#rd8�n�7P:��y��o�<�`�.>�Y�dM�@
��Id`@�<IG,� v,�*�-�\�=U_p�<���F�C}��0�- �c��(iBa�`�<�����h�17�L�G'�o�)bi!�$��&��*�C�?vf�[�bE��!�E4
d�t�`��,n~����\R�!��8��:UQ/Bs����+��8!�D��WV8�xKQNS����<m�!��F�P48E�G�-%Ox)� �Ey!��	�dgR!kw�*?��-q�@RrL!�A+�"��ә.r��z͋8!�$��I��2�.��dY2�P�e�{R��D��Qz�qz��#f,�����y�".{�tE#F 	��q�����yrCS>oe�%N��D3ț�y���s�Xb)0f�r�9�	д�y�4dR`��$ŠS^�H5!̆�y
� �Ț�m�8mj��'@F�6���q"O�����(�>t���^	(�t��"O��;0���1YEď#��"Ol<j�kU�C��K����U�<I"ʘ�Bi��[��S|��!���[�<���\b��#k�?����B��l�<I�V>����K�@�^��f�<����X+�̲@`�D�:aed�<Y2��7P.̨1O��c*T��	Wk�<�&"�kߨ�!+ي{�zh�f�<��&�*V�����k���CըFf�<Q��������] �4��6m�<	���g���8*��	5� 3qI�T�<1��Z� 5���@:u���2��v�<�w�5,�Q��\�i���Zp�<���\\:����⦭��i�<��%�(ڝ�%,lL`S���n�<D�	2!�~�㷆��d�@&�]b�<�S���#88���) n'��gU`�<I6�V?���a��D�WS��r/K^�<Y�B4E�$�qC�S��y�RM�Z�<	#n�y˘ �D��0"��1HK l�<Y埃`������/v�`�C��d�<�7玂M� �e,B�r�,�^�<��	F d�5pУ��&��D�d��Z�<It�V�g�Ţ$�$|�#�<`�!�D�5:��%�����6���e{!��o��0G'ƷHfj�h��_�j�!�$�#&
�|3ANN]BNY�护n{!�$�"gS I[R��`��AST��<�!�$�u�|�iT�=4}��K�L��qL!�]#�SҪ�"�XDz��^�!�D��\6�q��	2��B7��F�!��ʗ4p�x5��;x�-I��J�P�!�d���Z(��"m��Ѣ"��]�!�D��@���`���.b��@⠔�sV!�U�ebP��&�z^��p�
ݹ<C!�ď+��T:ĭK���K#,�!�����ً���M���%���b�!򄞰4�@����C�� pW��i}!��ƫS_49����0yf���ϗFS!���^�`�@`,��cҡQ%�d�!�؎m3���G�Eb`@ ��!�d]�21����f�C[��ĂF3e!�Ğ�hn��� 
Dr���da�\8!�DI+��,��ސGW�\��@Q�+!�_ |er���%GX<0KR`�&!�$şE�fI`�$W>?'��k�?D�!�dO[K�h �(B�6o@)��]?S�!�D��fS��`HĽQ��B���#!�$�E(N]2C
���0�9N6A!�dJ�vI�A��*�
[��5��'T�7]!�5{�V��'c_u�d�l�0|f�B�	-a�
��ƒI�����S�KNB�i���� ,����-�q��X�\B�;�H003&؛�����׀]�2B�	:$����fnɥ2Druh�R�d�B��$����+�s��T*�R��C�I(�H�t��w������qs�B�IS�XY�eb�.|�`�� ��<�vB�I_������Ƌ$�B���o��BBB�	�&��$�m>��΄�3�B�I- �!�E.ȣf���
�Īt��B䉢'����R�� ar�2�C�=�HC�)� ��At/#t� jW�h#t�b@"O��c�֭r�2Hba�
�|����"O��0��L/������|��с"O��(���7�0-���dh�V"O�1I�m�*$�Zco͡	�m��"O�Q��%(K�(9�u�_�1���"O�l3���
s��c��$ )�"O��6iV�B�H��,Z�	a"O��j#�E��])"C��Z'Kg"O��dIG~�Sc��r��"G"O�}R�A�,���a�9�RD²"OjQ�C�,<��#��ݸF�Z��s"O�W���L,{6�ё@W����h�<���.��L�`��ek��A�d�b�<i��biА'�-EP9����X�<IתɳUn��+�:B�6���U�<���\���x䀋�4fdJbT�<Y&L��O$�P�DX�8�����NL{�<9#B\91C` �dWG\���vmWO�<y�A۳)�8H���&wڍ�A��L�<��oĺ`�>��IIh����o�<av��6��+C/�i��rg/�c�<A�,[�JM��k6�5:!X0���Ju�<�夂=MxPce"�F4I%Gp�<�T���e��K�H�;m=
3�Qn�<1QaP�!��t�v�!#}���ʄi�<i�n�~��6@�: z�`�h�<1s[�����b�:�f���}�<iQ�x��6�)&Ֆ�����d�<s(KH&�$B���"�Ap�ib�<i�)�1�,hQ��(>@T��`�<���U z��%��7������OU�<����x� �J~���+K\�<��@�)��PB�oL�DR� 6�XC�<�6RAA�%��0>��ѐ��{�<!��'o0��äH��(�R0�y�<�5.ޕ=bn͙��/b 80MA�<9E�Q��p4�� �s���Dɘw�<�r��.=����qg�'w.�̑�M�s�<�W����@��%{ �Q�#T���DR=T��Q�a�S� �0��g.8D� `R ��T4�W	&�L�Z�:D��) ��S{�]�M�6,�6�+D�p�l�8�F5r'`B�	 ���7D�4곆	��v���/��)�2D�̉2�{/4�ڔ^=X���(��#D����,҂'{�A�C��;_p��!�4D�tK����DB�s���n�r�;#1D�؂�c�7W�}�MH�hɂ�a�3D�0�
�Ӏ}�L-޾��2�5D������'�`i��_�V{��
`,7D����)Vo��!b^?6��3��6D�����H��]��윭R,�S�3D��Z�cߚK�豢w�ڐf.�i�C%D��Æ��z�05��6N�|j��=D�d��%U��y�"�F#V�L<I��!D�d�ઋ IުH1�	1t,�	F�<D�<�׌��;N��+�!�$8ze
;D��#2�4��2�
=KMb��e�4D��A��ϴ|�����E.Duy��/D��b!ņ(�v񊱍Y��bQ�.D�rU�1�R���)��-���e�.D��`���K�r�� #"I�G/D��AT.��a����1�����-D�� �,)��3:���4M����`t"O�@q�j�3b6I(��E6��D��"O��s	V�)���C7鎯	���P"O� ��a���d5:�P�J����4"O��I�M�9*bR �F��@{��0�"O�(ȆJ.��AG�Dy9+d"OL	A(��ζ`C`�S`�*�@�"O�,�ᮃ�_�e:1
W��$��"O �11h�  �x��&�D|����"O�mą�_O���iIܦ���"O%���a�.���ߋ�&q "O2M!�D�2`��ɰG+&`58�"Ot4��fOx����1g�7C�T"O��Ə�/ˬ,xFE�*7nF�"O!c%W,��9��d>Z"Mp�"ORQQ#��o��R�B����v"O�Š����:���F�U�A�丢"O�X�!��`8�8) !L�M&Y�"O:%0R�]���Zr` �^	;�"O��@�h�5Q�%b �B<��(ɑ"O��gI�b�4��5�Ŏ3�\�b"OԸ!V�K5_���g��1e�0���"OX����ɽweX�&��5���"O���0o�@݃Uט �t�[&"Ol�˔�H�|H�P�m�	q�"O��y��/� ����źC�z=z#"O2��*�o��-k@o�I�"O ��@��Q�߼r�8��v"O\t����/af��BԜ�
G"OF���l�vBb��u��n��sC"O�q�2�3:�艈�΄�O1��"O"� �d�%�6%���S$K~��"O�0�f��T�hpˡ�v�%1D��l�<ir'�IN��(�!B�Y:SeGm�<QF�ȾJy"P
� ��qu@�M�<�1�Z�,�jh��)C/���'�B�<9D�םE�:LQR�ĉXpd���A}�<�0/Z5h4Z�i+��5O��H�d�Q�<A3G� ��*^=%椔��T�<�GsRy	U�D<&��đq`�L�<aFc�?���GQ�'@b���!�H�<�C�+[��y����a���j��H�<)��,VCbl�Ҡ�r�h8���C�<����i�0�
1�Y�>(���@B�<i��~�,�V ��7ުpb����<���9$Ǻ�`����(z"��Az�<��N��@���beꖷ5n��Y�Gw�<��j�0A�c�γ׭ �D"~�<Aǟ!(�B��3��
@�,�1��y�<a #F68�$A����G��u��#Uq�<�E"��Zi�x��\q��b#T�TAa	��d�MEJ����i4D��iã^%"ʨ9�n�)=����,D�Ԛ�)�2O9 $sG���`�2q )D��؄]�^��Y(�<-�xc�k%D�\�%m�)���1D�)����U��yR(Y7_��1��_��-!�ѐ�y�d@�
���`jN�Vsz�V�I	�y���2S\��S2�ڱ=E�����yb���Zd��k&+K�0jȴ  #���y��H	~����n">�j��)�y2�F3<�YRA <�,��
��y"��0�'��4�B��oT�y�
)xPW���+$8�Pw�T��y
� 4�Y�	�<7z0��RY3Ҝ4:V"O����w��ЃD�1�Ψ&"O����22�D5�b���@�"O`�U+�5* ��ԭ	�_��4�"O$�ɳ�^����0O~w��"O",1��+q����̎�crj��s"O��P��C�.T����_T�|8�"O^���
�sú	��c�=Ɛic"OP�f��ǶE�%�ĲZO��w"O�@ bA
w�
\��ۼ޾�+$"O��拉G�(�Pa[:p]�"O���j�z6E�� '& �P"O �J�LԜ����cE�<��"OH�8p��?����*D����"O�̣A��T�V��$a $i��"Ofщ�\��h��̇u�Z�"O�X
���Ts��2�o	5E�,��"O� %�2B��a�([��mc"O)���&b��))e�7t��Bf"O^�IY���u�QD3U�:"0O�9��뚄J+eIR2&@0�G�I�e�~��W�,^:�j�J+��C�	�Wd���G�@�ZQ�"�/F�a�C�I�.w �;�瞊-5�CAC�q$�B�q,��s�X	Y�,��ǃ="m�B�ɣgR�-r�	 o{`{­��B�ɭH̐]1��ǣE(I��H�lĴB䉰@�ب*��T�x���"��FS�B�I[�!��bF
W\��҆j��B�IzL���!/[e���
�8�B�ɮZO�x��hI�X��Pu��/D�C䉸E&=@7	�>h���6�Y�"�C�	-5PqP�]�p�Ĉ��O�0C�	f����/2�ĉu#�d?0C�I'h]9#��R1�PZ"�lc6C�	>K���k�`��
pt(d����C�
(�m�b�
0ml>�K�ݒw�B�ɧ~��U�&A�~�E*�	�'8ވB��q��y�4.�d>��"/�h��C�ɞ1��K�$zúhҀk�?��C��WO����̕HFj����;�'�&(``e^S�����W�,�0)��'���d��c��LR�"�$��!�'���Ӂ�M�>�8�A�׹l <���>� 0�a��y�$ҐG�B�b
�(JK��)���ew!�Dr�8)KA<\�E����N�'� ��͍�-2����5���h�l~�����eF�5#!�?����Íl^��ڵEG�p}Ftѳ.?Ʌ�ˏM���>�O�XJS?����-�
�`��O�Tj3���?c��U���h���QKB֔�C*R!� ��I����W�
ɜYQ!�;�?Q�\�8 ;�d��+�|��`��-A+5�\=���
��Q�ȓBz��� n]*���눩L��(�'L�t��N,&�$u{�P����l)�Q��)%"v�eW�3����"Od	A�Bs����s�3"<�`V�W� � �!�-މ90x	��`��3�O�R��s��<Jm��;"��Z�L(��ɽ�J�p���+4����D¿��A���0��(�p@Y�
C2�3� Z8�p���˪.�\C�l*H�P�)>�~��e��*K�-�p+w�S�M�HЗٟP�˦dO�e㐤`���N6Ip�"O
qKdb��w�2�)æ9��S��зF �EAW��1e̤!H�:a[��9�`P��B*6w�c�E)~i2�a"OԹ+��U�<�n-�SޕgS��"�\9f�TE�� ;��y1�e
�/-�ĈU��(OUYPe@5a��k#�H%_"6�2��'s�@ʥ"�F%y�E�%.��Z�H�m\$0���l�Bi��	#Q����%D��fI�	j�b|a��jd���?� M�<A� Z�m��.�����	��d�g�? <	pe�TLi<��C7[�XUH&"OI��m�g��"���`�D(j!�9��T6 ��uS��p�E vY����"n�rn!!����nܝu��X &	*D����ܓm�n��Q*�4�ܔ�Tψ�+��=�f�	��P9�,��L����H\n����0#�T0q�`���a{|��'B$BA/�Z6p�3"M�L��L7%���|P1�*,K��py�ʬi|���>�N�td���A�
qO
\�� �����
�/���[����>�\�'l mI��̩$!Y �a�b�|�<I�O�L� u�D���#/�	��(&w��Ų�L�8P"Bڳm�Xdz�:�Ӣ��ë;ʂԣ���d��h�C.�!�$�Of.�+�SZȢ�z�`���$�t���$��u��)�t�@-��M` �s������I�3̒�N�j�1��S1��z%/}ZX��l�5�@(��7 �\�hر}��"����Z0�UK�@H������4�%�KB����*���qOn�K��؅W��=���Y�2[<%%�9Tژ�3���`���!�0Z�� �
���H��(�T7�Z�I��9����Dn�F^Q�GH��=<�����veC�w�
�q1&����r���I�*�:
�'��j�˂�;�ܪP�@2��Y��� ,&� 4�s�	,	" ,3���u7�)�TF|P�M�M�r1�1"яcS�H��'�Ve%WCp���@�wDJI�Ƅ�Y9��lU!YI
�iW�4�O�m#�`���i�I7).��)e�I�:�$�� a����� �Ԉ�'B�?6�� �(=�BB��
��Z(�ؠ�sJ�������萱`��=���x���'�t(�l�-*�=���J�b�'e>�A��C�n�kwsZt���'4��3��ܠ!'*98� [�n>��'��Q��G#s�|pHL1iK�'4�X�']�u�|��싏/⺴��'޼�"J�=��놺hu�s�',z�[���g�T�y��~���
�'�n}3P
�V�tH�a
��ؔ�	�'+�-�ԏy�� yd�]1�h2	�'�!頄�x���S���L��'g|I�(֋7������x�C
�'h�	�ŋ��:)�	s���yQ��
�'>E�&d�0%���b	�r�¹s
�'�AӋ^p	��1�T�g�~,��'��	x ��*X����]On4A#�'�%y3��%0�� �����
�' �0�AA	+I x��ӥU_��8�'��0&Í+\z}�֊_E:�9�	�'�"�qw!��<�0�[8A�9)
�'��X�.Z#	&�Zs��D��, �'a�U�*1���af�]�C�����'��5h%'F=(r�[�E��}�
�'�:]��\�	�H��#ntJ�
�'�(E��Jɛ��6�]�Y[lI�	�'� \:G��wW��
vIҀ'=�L	�'�D�؅�N�e��d�UĒ�A��c	�'I0E ��>H�l��Ϫ8��83�'
v�A�T�Hj��M�2�60��'�����W�u"z�H� [�P��X��'�z$�`fܵ	��06���K����'~�!�s�ߤ}k���
��:d.���'�p��S"����E �O�1~"�@�'p��7��Z5
iѡ&"��AP�'/�9�3�IF���E�S�$/�P�'l h���Ę+Q�u���&��%C�'Q�j��Bv��A[u�,��u�'��ܰ� @�>&΅q"(Qa5��	
�'�����!��}\u[�TwhB�	�w�-L���*A�AP(w�B�ɷ3\�=HuI+X���ـ�bzB��;�d�4k[9K��A�N	!IB�)� �ZĩV5�HD3���}w�u��"O����劒y�4S@�Q��d{�"O����� �faӳ�ؙO�^ؘ�"Of���a9���������JP"O����I�"E��8��S�5� 8�"O�0��R�����D(nͦ�A�"OƽH���N����,�U
�"O���k�&}��TfS:e�4���"O�P�S.5y�@���T
G0ti"O\����\��l�1s��5:2��P"O��i���6^|��D�|��*�"Ob�;�Fߤ�p��b��!n��Q"O<�����//n��u#�F�6m��"Obh��J���9��l�!Y��aU"O�`�r�Ō�;� ;�ұ�"Od�y�e�%"z���5	����"O��H#͗�ZOD���=9��Zt"OU)�,m��=p�'��`��"O�8c�D��cg
C��q�`s"O>�˖!K�q$�ϸ`� ����d_$s��x���iA�J�"|Jbaض>�l ��Թ�Py��E/R�ld!�/<�uxG��:�Z�:��Ɩ���'gwQ>˓jN~u`���$�J��EM�3ZkR�����-�B�Cbyȣ��Ye����:�(�d&Q�=����� C�,�s�'k�x	�a�/�ay�.�lK���B���
[<9tH�9j��r& 5b�L���@�wk�B�Ih�b���̷y�,� MP	9|O�Xy���|�:c�_�v��|��ğ�S����+��'����Q�<�@�"yԴA%OQ�fl�Z��$Q�i�V�!i�&L�Wk��}&�lJ���'h(�ࣕ�0R"x! F%�,J�C	�?����ǉ\�n�PuL�s�h�
��4[n��I��T�azb���$Wz� �L��8�H�@'��0<��E�eT�i�?��!��Œ?�Ty�F�^Ad�A�C���
��_h<9d��7�^�i��ɔN�HY;�SN~�.�+�j���F���Ё��Ѫ<��ؔ��d������T�Y�@J!D�B��4��͂�b\���ىD# �2 �|+���z+�E !�[�L>b>A$�lIΚ%�pӔ�+�����!�hQA�N	>T0j�g�D���c�A[,~?����e�1u*A���$����I�^4\�j�&V�Q6�1C�*X�P6���$�;4�Ԭ�1XQ�ک�!�.���+$S�����C*W� ��n<4���gG�(s��a��"�0k��,?��(OMM�	9h^�t��h(5.]���O�x�CJ�Y��b����h#
�' n�S'�͈MCBXrRBۇ8Q���p�ά,O$*1)���	����|"I>��L�'e�@�3���]I�����j(<a�fӴA2T���jDe�DL
$�L(z��X+TCT+^�R�6���B!���� ,.�m�qF�vb���ҠtX�x�is�֕�VCML��u	0Ë �V���@�qT���"
D�����xa�����l���P#K*�D	�{�� � |�hA��0�'�VM��$S�=�T�'7C�i��of��I�O�k�r�1Be &���6��6������Ozb��`�g�ɼ2I�x��ΌѾ���l* q�B�	V��р��tob�c�b[�49v�i��l@aj�FF�+a{�ƆfL�ȂB�W�v_�T�AS��p=�5�7րy�4@g��'����d��%�V��Qc�)D�\Q0��5l���䩈�
���qa;�	�5,h����x��L��Z8!@� ��ɘ5kI�C�I�zv�˖bH��v�	g�ֽ��C�85� (�� B�.�w*��B�ɟv�i��U�I}X�d��F2�B�I�mN�$����o�"A�ï�'�TC�I*@����)ɲhK4��1+'>�JC��5@W��b��3u�X9V�L+��C䉢K�R��Ԣ�
X��I�SֲjqbC�I$��u腯D�K��i�@���QP�B�)� x�5������;�,c�N��"O���`$�yG���ʘ����є"O���tH9<4:��d�N��x�"O<E��E^X`�e{���(t��d"O��v,�$I��br��.�%J�"O�\��ܴ(����7mH��*�"O�);��ޡ7��`�%�G%b���s"O�qJp��CK��� �x��tP$"OV�0��3BP���O��e��X�"O�)t៩D�Zlӄ�@2���Q""O��GKN�<�I�-�y����"O� K����.�HLC)H-x�)"�'[���p��*SB����BI�+iʥ 
�'OB���1cH>=0Tf'vh	�'y���L��m�b���.��#�'���)��3y� � t�鈐!�'y�9:B$��ǈ	B�i�c�����@�F(��悤D�Fb�o�c�0T�ȓ2R������2����KY�$Qz�ȓ_�0���J=\N��1�W3�z�����$iu�P�?<�q�b<�f��ȓK�|UJ¢�5XB|��U \�\�p��z��j� B3MZJ��$.��s8��ȓ"p�a
�@��w�
<��)ńL�4��0}`���@ Th�X�>D<�ȓwͬţ�Ji�ضN׾	������ ��"W�h�4hğ!M]�ȓG�}+���L	 ���G������ȓ5����i����'�R�P&p��$f�݉7���� ��C�;FńȓO\�ձ����	�~}�%�*�����$�rl�`�V&p$j�a���u�ԍ�ȓM��:��R��b��w$V)�Zx�ȓFմ�H��*K��iG�E q�:T��j�i�%��V6��	�!jz�	�ȓk�@ ��&�n��)�
L�ȓ{F�F!'|U���<(�☆��1��@���d��ƅZ���ȓ{�.�B��}��i�=C	�$��/y��W*�Y�������,����$Z���P��P�_3��ȓp֔`���5s1ڂ�4P�����|����A�������V1�mʑ��� ;�g��w�)�ȓh�&�����x"��˫/,&��ȓ/�$4��c>��M��+B-8 �`�ȓ/��!z��ˇ/9Bx9��P�����/;Fp)��!}rnĄ������9��iU��y��0c-.���D� i3�DS��ē�vQ�&�I&k[a������Q�A� �遇��y"j�*|�Ԅy�1#��e�V P���ڧ��mʐYL�>�O��SO�7x�Hذ�'�(e�D���O��3�,զ�+$�ޠXm�}�v
�%l�j �Z�A6���I	X?��;0� 0(H��:��2K<У?�o@Ȳ���"C�*���4�&�9e�@2qT��*#/��f�܇ȓC>VD�$f��>X��H�0<% 0�'�h0���O�8��@�HP���pA�G��z�f\�hP.Z�T"Oh�ƒ�N�����((c(����
Bh Y�d��,k�J�
�Y#(��3ʓ� Փ�a�z�[P�x�^��c"��*����C���"����[\��kr�B�s���ޮ3"%�E���p>���	�i���J�}�P4
��M�'�Ȱ��O�M�u�8{�B(:Q�?	�EN� N�F50�ꛎF��e"D�p�ӄK�+'��" jV�	f�$��7<I���ɯ�t9��t`h���s��a%GV�x��!�'�(da�� 'D�� RT�BG��&�8yWĞ�Llv9Џ�'(r޹J���sL���T���T'���(O�h"�ܤ2e%o|X)�t�'P E�F�T I��DzC#D�
#�|J�&'� �FP�T0���%0N,\y
�t\��&�@�K��Y@�Tdve�?y��/�� ���"��P�V*%�:���p%�����
'p��
qh�ȓHf�X3�Q*�$�0��i"�M8�0~ �jѮ�l~��bڅLb�?i��w�+�$
�b�0T�g#0}0��'[*=rQ�ߝ��G��8)���A`�S�E��aѪJv���BL��[(1R1�_�'�� �e+��Z!:6�6�
�V���B�MF:d�2s���j��8´�	W���"U����4��-ΠI�`�P��'�0�ɰ�I�+�h1b�g.>��{b���}�UI�
CDa�ǠJ���$C�!�?��a�^�hŉb�ǩEv�@p#D����,8.��0��S�LA�-��=�"��^��TtYei�U�@����	Զ�y�d�;vс�rH����4�y������ĺ��"=��%��>Q
�q�K�.��: ���Yi���������Fy"�� mlL��Þ�L���5cA��p=�' �p2b�0@��A(1l�.��9�l� ��w K�4��oR �|2ް?R�m�b&͠LW�	i�%����'���Ғ��l���ɢl�0ny��H*/�S$QrA�W�V ��4� �/E��B䉒Op<srI�d�����aӉg�0��!��#��56��:�X�'	R�O��(�;S�$��C/��,���I��I	L�j���P^@#�٨+�!RPE�!Q��"1�E4 Z�����ѣR�y0R��k1�I.�xLk"��j��8� ˓T#����N�!
�$yU�܊,�~P�u͒�FuZ��u�M�:�b`��m��]�(�bD�'�q!qφ������Ea�@����ݨR�>��b^�=>QH���!1>Xi��N� �P�`n4D�T�w�T��� ��N2$C�aR5xfNj�`ߠ	�����✃O�F�Y��	:�ŭX�,' ��t����k�*M���1!��*s�T�ȓ"���1�C�(6���y�!��}�E��o
�S0�лT>�M��
" B���1ZU��4����ѶC�T���^$y�W�
����K쟰jB��ȓ��0�d��Qg�I;�!Qo"�|��$�Z��D�Ήd@� `��ji�D�ȓ�^��QBK<���ե\r�І�o8v��poQ:���؃i��S.���~��\Z�́>�4�*7#�$rx̆��.�C�f�-�01�^� ��ȓ��8�׀��A�Ph�ȇ�e�4d!v��9C�Vq��8CK�=��g��m��gC�t�P�&Z�r���ȓR���JB/� �N1(d#E#f��=��Ufka��6b�x�[�N�h���ȓj
5Q�����z��Є�5�H���n��0G�5�l�:#)��+���ȓz@�V扖I�0��Ė�.���h�V��@���D"��Ja�T��	@�DÐ�N/e�����`�D�D��h`�4�GH{�FɃ�
ŉ*r.u�ȓ+E*u*gc��G�\\R�o�@(��!��bQ��$�a����4d��ȓ+�T��aMY ? dq ���`���ȓe������,^0T�T�;FL�̅ȓRX��(]b�Z�$�7*t��ȓF�Vm�6�:��Mʁ��fxJԆȓe�r��խW�m:��5a�7��!��o�.�*�k�&8�u���,=Q�)���~IK��ޕ!��8X�5yͅȓ��a)rE�_;����a�5�V؅�t|�`�U�N�����n ���Wތ�7�S���RP�z	�ե+D�ģ@̝��Q���:y�AY �(D����G�>6��l����1
+�9�@'D�� �@�ǁ�:a�a�b"��M��"Of����I. �@a�T��%�G"Oz%�'���[Z, ���)Vj2\;Q"O 1�G�_n��"��LG�\��"OzD���
:5�1B�@uh�"O�౰�$.�f��c�6.���"OF�Z���o��D�"(F�2-8Hhr"OL,��(
���(7kz�B�"O.5��U_�!0��]�	�"OE��	�YZ]���Ɛb�d�X�"OD�S�/âC�rP󶍋�k�z$²"O�[�+!�]:�閲��*�"O(�w��n8Tn@ ����"O��ã�4#�a�dM��T��=��"O�a1�nU�^�vi�ek�tl��"OH%��f�m���+ԫK&[u�T�"Oh��gF�x�d����"aw ��ȓoj�Xf�Q�@�"�K��NA�ȓ>܀R�9r���ꤤ'[�����l @e�*�R�-�9>꜇�bu��Vf
�D�7��N�D(�ȓ���"�$H����ꋮ 2���@�8�/Y0M�w�L[2��rA/D�`�F	@;�f�LA�G�<���)D�,#B+���*,H�	R:�*i�[HB�	�K	��z���[��(!�ڞB䉻`�|DZ�47���#�΁C��C�2I�k$�ޯI��F��)��I%D��;���[^<����x״����<D���3��-K���J1g��zZ���k8D�Ժ�Cր
��0D�,s���i��,D���W,�a��q�U
D>Wh�%K&D� 3��܄*���iE�1tvӥ'D�@��!��Ghhњ��2I�~E��9D��3�{ ��D��G'ru� 9D��@uH��%hxQV&�/;9�\�(D����"N�`Pz$�M=>�8��:D�h�C�;- �`�6�Ě!��`A�9D��PCȀ1]�
A�5"�8b�6D�����,9CF����[����e�(D��i3�E�f�ިJ�\(�} ��)D�hv�$4b\Ԩ7��y`����$D���d�E9 =�6+K��q0t D� ����5/�u�g��p�"�>D�,���/��2V��=G�^� g$<D��j¦W�x����ɗ8�b�`�9D����m�;0�d�Q�kF�R�Qї�5D�����G�3�4T��`C,�x��4G1D���V� �~L9���*8Z0�#ԫ,D�� �;����jH�;6���L&D�d���/�,�y���0��$D����e�����O�n��7o0D�@�`�l�RP�dA'io^�2�m.D�|hhRu�͒�+q�>lA!�!D�T���ج4Є��֢|>x�R�"D�`�3(� t�@�p撔L	&0+��/D�̓f���^j��Q4(�tc�Y#Ek*D�܊�eC�VBٱwO�$D���˓�=D���*D�Δ5s���rc�}�2�$D���u`�4S�urQ�͋-t�	�r�!D��2v,�4�8�(��X3�!D�(y�e?��eh���\��Mr�H<D����k�+1��� �&P)֍p�8D����o�^"��a�#�l9D�� ��6T��§֯]��<��"O@��COV�Q���D�����"O)T�ۢc�6�%�l*�Ɋ�"O��C�`���x�G<ML�"O\e���ȾkM�}�wX����"O�<@��B*,�
�`ae�3^���@"O��	s��O8��*U�SI���i�"O(� &��9��h��?�� �v"O�*c��w�$����G�V��q"O��	�*C�IcX]��,3����"O@I��/��h��D4wD��"O$!��-@^p��! �"���Z�<��	L/P�v\s��)BPy֊�X�<9��� D�V��+�&)�nYAD%�m�<ɣ	
>a��4��C6a`+c�<a��D�=a��FO�-gR�d�[�<�BCǫaR� p/�-7z��U#�U�<i5���n�h��ܫj��E��E�U�<�1o[=	¥J�nX��>�qBgTQ�<YCLQ�N�&DQ�!G�uW�q�<���0t��L1$�Z��f�KB�T�<��L�1H������`�,��o^k�<�jڒ���{3b�O0�b�<��
4mٔ&��"�,��aZ�<�T�{����&� �.Uf�k���b�<1��I�u�Xa���2u.�|�v�V�<a��B)��ҳ�3-` XY� �n�<Q$�T0�LQb����(�@j�,Y�<y#*զ1����BN�'aČ�*�*�Q~�ܖ��dB$j������2�n�@5�'���+Ȩ��#�H�)��V� Z�o��iJ�]�i�DX�vӜ�Z��M�⼣'��"��ա[�h4I�Ϗ3aܔ�" @�@�Z���$���0|b���\6>)��W������& ���M<Yw����0|�"ڿ7��Db؂E�.�Ъ����0��Y�3���0|*G�8���͝�9�ؔy��X}��Ԉn��a�y�ϸ'��(ز
�M���b ۳87��:ڴZTeFx��i�Cw�����wm��AG��*6��8L<q�(�On��.�'@dH��1bjM!�IY�U�O�ВR�'3:��ç6���JbYh��P��t��^�l�	;o�(hէ#�&U˱�����1O��Zcc5*7�S�^<:�� ՟HΧ[(�O���'���@�6�>xa��Q��}z�
!>f�h�×�M���Pr>)�"�[lK G��DQ2rMܲ(C�lh��6�Mہ��"JG��������@d&Ӎ84�,B�VL�4����'g0�lZEi��B���f}���7�+ᢀ5IAH!8c!V��(�lZ1b$^�6	Hiy
�'ka�������)'���Q�Vo�)��OرO���Ʉ�B��\�5و?�D�s�"�*�Nl�>E��O�ԠM�>S_��bO�E���k-�v|a�d��7�>��␒!�I[U(:��'�TB��4����?:0$quΆ U5�Qr�QI�2Oh̫�6�)���d���Vc���ZV ��D���Fx��	
J:�=q�J�&������B;mk�C�S����t$�b��J��1�E����L0D��Q2G�� ���4Ԗ,8v�@��y2	�x�Q�*J=f��	��햊�y�Ö�0�E����ko���f�$�y�t!�� D�8-�4���@���ykҀ)�Hɉ�D�N��	ɷ�y�/�/����%�d6�%��4�yB���VG�y��P:3�r��e�P1�y���{P�(y���6o�?����h>�p�7$�}�������}���@�p�BӉ_"�8	B��(_�
}�ȓ�
p2'�I�a���$�f68��r��% �z����X>H���I)� ׄA�'�`��Ä׼&���S�? Ll��!�8�>8�����qE�c�"O��A(Y�
U9��ٌ.�<g"O�PJ��	�0�q/V3�x�"Oh|����jdr��%ND?/���&"O࠶�#Tgth��TDL1�V"OZ�)cn̩l��i3Uf��xL���"O�� �Ʌ6'�-�C$�f<b�p�"OtsT�v ��٣rD�8�"O�A ��'a]� Y%C�4"<йf"O ��'oE�/��	�#rB`��"O�-Q&L.N����!�_:M��"OF `�L�#y���3�՜I�h4P""OAfK�� �⮊.P��!� "Oʍ�!�ϙ-cb��p���vȋS"O�:�F�$'�(CL1A��s�"O�`�(^�`0n�k`b�{+����"OZ�B.� ���͔Q|��"O�EgEي"�t���O�7n��,�'"Op1�$
1#�2(�CeX�X��5�r"O��Ӗ�ݶ,]�Qy��̯b�~�q�"OVT`p�F�t��RRd����
"O�����hZbP#�b��KW"O��Ҵ��`fL�E�D��ػ�"Oj���勻Q�9����"��LKU"O�)U&W����4f�}��"OR���`�$�e��F��OΘ��"O�qVNؐy�z��0��S^�Y`"O��A)SM~@����
Lt({s"OB]w���w���g&V8�3B"O�8�J&��x�%�`��I�"OL%��!@���$Q&��)�nTр"Oj�y >u����я��*vjLp"OFᰐa�:sl^�f]p(�"O�Az���B���F���U�@A�"O�T��G�B��1��[��d�'"O"��4ꚨj}Pu��Ԭ>���H�"O�m"5jJ$E�XLK�K�2G[���"O��F�t&z�aب'���p� D�����ajꅠ�"�9I�9yCa:D���D)��F�L��ȝ ��a�]�C�ɡ
 ���Z<e�m�#*ˤK�"B��	V��DZ��=�v}��J��yrÓG���;cϖ&3tQ ME�yR�͓d�ly���/� TQ��]�yb���=u����_ ����U�y�肌]}�I2@�W� ��ǌ��y"��йQ�`V�^m�fC�-Z|FP"���4jVM�䊥3�B�I�7頼�	�4Fi0�+�LɰL:C�I7G���r�;<nTq��9�ZC�ɉR���B�K
%m�TĢ��$&�C��w�t��N< (C��,	d���"O������7���ȣ!�TP�R"O0�36l+ �$� q ^3-AJ��2"O��Ԁ�9M���s���
Y���"O�@�"c YfrpΗ/-P��S�"O�ɶ �/dw�}3�AI �E"O4����L	� ��i�?	^\U!�"O�%�7�2l�$�k\%qbN�k�"OTYg��NО�SԠ&C��R�"O�	�Ɂ<\.m�`ЛQ�P9�3"O.<���7���/�e�q�!"O`�+���-�:=9��e°�ۀ"O�8t`��m�ʕ���Ѹ'��5T"O� FtY�ϯxW���o4-îe@F"O���J�����N$���B"O���% ���g�]�Ltv�1�"O�=��(��%Q� �u�ƺ��$�4"O�P �,n׾�q"_�jB�"O5��4j�V��P�0B�`E�s"O<�ⲮX'N��� 9�@���"On(з(]�~�p��
��Ě "O��qňLǸ�Iԁ�<[�ڀC�"O�9�R�V�<��,S@�	��p��"O�����>P!"0�ŀӜP��1"O\��爥sh�5+��G���`8f"Or��D��=b���"� F��H�a"O���`S���%�ՠ�>c�U�a"O�=�tn��jD%�2B�0Z�(��"ODD�e��:l�����W���d"O�0�V�V�)�����Ⱦn��"Oب��I�6b���$5&��"O��	pȞ� �10��11v"O �e� �����ℜ%��q�"O(��倏&O@Ċ�[�L�x�2"OL��p玈G��1�c,�^0a#�"O���rg�!zn^�bu��~BL)"q"O��C���5�vA�B�	RS(v"O�tµ�RPZ�`��)�8C<F=I�"O��iR�ݍm؜��ӊЁ 
$u�"OЌ�D��\���i�3G��(X�"Ox����-zK�Y��K�r��"O�a�σn�|��ڨn�>�xP"OV%��(�.H��\	��!"O8�i�#K ���5Fޅt�L�b"O|�q7�]!|z��a�f	�v�H$��"O�AB%�S�xr@#�㜨K���V"O�l�fi޵L썁����p�!H"O^�6a�wg�u���*l��@�"O���Hβ8T �Kp�^x{�"O��BtΝeJDݨ�(J�U,�H��"O@AJ�U)Y�0� F�4��:�"OlL��膻R���9��]!s�|xy�"O���)H ��HR�*ҁw��I�""O��*�ŕ#�����+N� �H5��"O�8��d#-q��,� ��q�!"OX��+[,l�H�ѥJ"���9�"O�l�Ո�g�ƈZW$���v�c3"O:]�3�L:�~��n#7`�p�E"O�u�E�wqD��oHE�ڲ"O���n�Ԗ���N5�'"OD�V+B�@}��KK&tu28�"Orl��G�p{©RDKk�|���"O2L*5J�WGAy��:Hs����"O������#��%�Ԇa��aT"O:0W�#Hږ���LfXt���"OΘ"S��.^
m�CհKA�,A"Or�j�l��&h q@�D=3�9V"Oʰyȣf� 1���_$'�����"O���hQ�	o2m
�(�%u��lk@"O��Ң�	�h$~�9A���_֠�1�"O���p.�/<|)�qe��NĨP+3"Oz�h
03:}"D4.�@%�"O��d�ڎ��E�78�Mj�"O��j4F?r���&�'Y���"Ob�����S�(�J��؜m{ 5!�"O �A�ᆏ$����$D�\]��*�"O�5b#�V6v�d����>m$��&"O� `d�@н4D���-�h���"Ol���LC�X� I�٬��e�G"O$��w�ۉO鈑aR�{t,�q"O�|��A�{{�txB��Ej�p�"O`a�C>&�ЙBS�hK���"O��¬��*9�R�E_��J�"OTl9b��2Qk�j� j�δ��"O��P��^�౉��U�����"O�ђ��*�FL�h' Nj)��"Oz0ST�ð]{z�M	�=���"O,59�O֣n!*�ɏ
~2��"O�H����l�� BD�,t��;�"O��!jԋ"F D�%��y~��5"OUcs�+,R��eE�&q�4"G"O:��@�C��@0�-�7eR �"OuQu�Y�t� v
�	vءz�"Of���L�:^�*A#��,C|l:u"O1ː�F �~�"v,��+2�ʑ"O��P�욥nen!�֡O+� �"O
]�Т%!'a:gAj)�@���y�+��"�h�@�,����wIF��y҈�$����AY:|��V�$�yB�W�x/8P����w1�J ��8�y��8
�y�GH<U:�*����y�쁪KMd%��$��i�81XDC��y�O/U��4��@1`��4;���yr�]h5���o�P�̌z3���yR�Fn��ٳmI�N�E8`�[��y���5\��=�&	C/�Q8� M)�y�"�;t�$y�U4:O�IQVD�.�y"f�#����j��%IF��yb]�Τi�� ��rTB��e;�yR銣s�^!�� �!�biR%�Ӑ�yb��O
�,�nN5P[̭�t���y"fܵP��������f��eKL��1F�{�nf)���ۡV�qE!D�p��hB��̄#��n��Z�b?D�0��a
�3f� z&/��I�d젂�?D��ʐ�.#�ahRC��.0	ef9D�0)��ݡ-k�Ƞ�m((� �"D�@�VC�j�xU��@�7��!� D�����v���P��V�7����;D��3�	�h/|H`TO��\��x�'�=D�����Z!�h�2����B��"�:D��(�g

⶝C�A�	G�9B�:D�����N!D8�
��8C��XP�%D�$�PM7>�& �]e�k�"D��r�3o�� WNK�'�� �ń#D��"`��.B&�,����&V����`?D���7j�"��i� ń'���@�<D�h�#��	r�F�s*L��&D������d¹b��6q�"49p-?T�T���5!z�!���f� HA"O� �ЛnD��˜� �-*!"O��+���K����' �8X���c"Ox13��(ta���;�.�It"O���(΃Q����#��O��4!�"OR�z�   ��   :    �  �   ,  �7  5C  N  X  �`  l  �x  �  	�  ��  ˒  �  O�  ��  ӫ  �  X�  ��  ��  !�  d�  ��  ��  |�  T�  ��  Y�  
 a � �+ �6 �> �D 	K �N  Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�� |d��"O
`�(�;���8���-0��1%"Oj4��ND^[��"3/9�0|H�"OB���H��*�ʞRy=a"O�味V�!X��!&F�:J�$���"O,��a
���C�Ą�M�"O,$3%o�-���p���+Ն�:1"O��ݢ1����`���y14]2��i�<�6��{_���c�H�`�fX�$Kn�<��A̼VI�xR[�)�Ć�pඤ�ȓA5��('nߡ4�� �)˩%� ���,��r�؊b#`T�eT09���ȓ!�b��g��}�8�F��-? �ȓ
K|m�ș�VṔ���2�%�ȓ"R�X�j�4JN�1�˘X�i����̹	_�jZ��1!g��zܶ��ȓgil,*�J�
j�Ne��i�J%b���f	�(U��:���G��$Y^م�~r�� S�%T"���k\�jx�ȓ|4�1�îJb��@ӵ�ݩn�V��/[`�"�v4�R�!ʎ<��M�ȓ`:��z�ؚh�J�Z��$HY:	��H��p�m�C1��!��B:��0��EnjZA V;9����J[
2���	��4'J�EA�IVW&��~�(aZ��ӹ�>� o�Y�|�ȓ�f�A�
Ο7�H��M�$�����mޠP����/���ANXo*�ȓTv�����{ ��-7�*h��I��sB�8�8���3����ȓNe*M�悡;������X�o��!�ȓ'lj�#F�m�+R&;�|��2)n�C��0S4���T:
b���:�0!��e֊��)��ͷV��,�ȓ0�&�8#���� ع�L�����;�P�AFd���,w�6dΓ\y��"~�ӡ��x� \��EB"�Mj�j�^�<Yk�!( Ӱ��9xrr�ay2�/�Oΐ�%爉e^��Pӥ~R���$"OE!�c�hV�Jc���� i"O�PAiI;i�Z���U'c��2"O�!�≘�r��h����h�X��"Oz�J%�%�`�(r�Ѕ^e��A"O�����)��#�$�i���"O�|�ǣ��{�h�����aZ� %�	ɦ�G��.�!�ā["�R����&I
�p>qJ<)1'\8|�����-c�$�.Qw�<��ϭ:����oY�630�' w����(�f]�S���`d��F\K'�`#�"O(| aA�3��8�`Lޱh���&�S��yr��E�D;媅,pJ$�
G7�y�&��\����"\0jG�M����M���Pqy�l�q���R1�B�_^6A҄'j!܀�D5|O�a�"�<��,]�`�H��͊���}�F�I=�? f-�S�O!������{B�p��c��V�`2�I4&'a�ԈE�N͠	8afF��xԨ��U����HDX���!P?ȉ����%L���ڰf��]ԛ�}r��R�mX�o@��D-yڱ��*D��x���.m�v�	ş7�� ��+�<�p�'6�؛�Q�i���'�:�21i
�'�<��R��.r>ވ��IA�t�Ҽ���d),O�M����hE� �S��}�h\��"O� �� �aC-?zȘ�s�7l��U�"O�="�E�l����nՋC�F1��"O ]�بA�V�ö�Z�/ebx�P&7D���")�)cX�J��֩(�4�As�6D���&��R��6�I $8s��4D� ��	]O.�e�D�XrnP�i��`�'V(ҧ�3��O�2��&�P:W��0�Ȱ.!�$M�M�n� ��/�|E���L�e@�'}�|�H�\�D�j���P|Sd��8�p=�)O��(�`�Q%�����pBĉ�F`��sX��@�
�H�D�ȢH��H��h�<���)�S"�
E!3��0|%*L�sA��$�C��)x�|��喃tĢR�H�6x^B��;Y2��J��F�
�֝ڄ�r�B���<��o���������pe�� X!�Ā3d�Kc�̭�����)$�!�dܩ�H�A"%��L "�!#Y��p��e�̀=�rN�	V��p�R�	]8�t��j�>O�^�!3C�G)tq#d�4D����G�+��i���9�r���fqӸB�	@��D3�!F+d{(A(�U�tG�b��Dy��i�1e>�U�.�R�cJ�bA!�d��PQ3�Cof*�X�Fw��O����	,�<��j�	����`�ρ<s��ā�Z�vuH���^yV���a��C�IK��X�A�Q�%�,�KS�������1�,q��@�"�1N��1lˁJC�� �"���N�3m�֨���b��HD{J?qe�S��B���@��+D�`��Oؒq�`X�,�3S�t �4�}�$K<-O1��I�f����Q5����G�/'�C�)�\��,ٌ`gt�����X�f˓5��}�,��1="4Q E�l!� �Bیհ<y� �B?�O4H�䂦RM��0ŋ�(^�v�K"O�$�M��q� ����^��=����W>��b����
��:]Ƹ���K+D��;T���T�$� Cn�||x��d�O|5�'ʛ��Ld?��1O"X�����t Q"�� ��"O�K����	��!��D�4�C�>�)OX�FzJ?���%�.%�ԃ2��2��h`k$D��K�+��$�KE-���h�Hs�'f�>���'i�-��G�.�Qd��G�
"=ɋ�T?��qj�.�6����	Rh��������	$
�jl�f��Pq���uiQ�K[�B�	;��j���tN:�Z����x7�B�I<��8 O,��@��N
 z�!�'	R�C�CX )�ݰ��0F�h�	ߓژ'頰y2,�=#�K��۞j0d���'�P��RK�[c�4��F�_���
�'ǚ����E1Vp� �Ӌ����#
�'���I�=Y���wm^�F�B�	J>љ'm�y�Jƨq�d�qQ�� =�2��6/ֈ�yF���zdB��1펰� ���y�b��N�ԛ��M�0�4��@`ŉ��=�yfO;,�HL�p䀂,�䰠���yr�2Vf�ѠfUq�@�RG�Ŏ���hOq����d�ð
�$m��@��a�P"O �#JK Ѻl�f� �t1"OH\�5$��&]��st�\�{�nQ�"O�|0�đ�}6JdB��?Ў���"O�y��'Fc$�I�u)F(R؄�"O��cP��[�|POԺ'�(�p�I'a�t!D�i�z��։#�\����N��'�ўb>Պ�cbҞ�b�I$)��9TlN4�HO?�)� ��A�K*#M�Y	�H�Ej.%3�"O�y%��I&�$hb=8�~ઓZ�D��I88RAxtǬw,�J���(���M��;�:O��L<�O]�I�|����M6DB��� 3V[XB�	�Ԇ�bv�	�E��Y�4)�;}�R��<�v�'�O�O֝��ٺv�F�it!��y.�	[�'�a`V��?���A\1�ܑ�r+:ʓ��<9�㖃 :���J�)G���ˋ{���"�x���;'b��%h�zxRf$Y"�y�%�7X���c+��V~)��ި�'Z��=%?�sa�9Y�a��є��a���7���������e ����`�e&�-oC��n��-���D�.��@!�j�"��㞜E{J~
[�F�� ㄇcyR����q�<��XB}�ĹE�&e����A�^m��0=���O�k,�M$�T)1�0�Fm�<#��,��[��.T��T����l�	�fב�b>%�2i�c)�*e�R�haD��B�7<OZ�1"����O����)1�>e��B	�` d�"O��F��aF���ۘI�r��$�ɔ�M3S��y�O�\i�3�L�F�R���ѵ^��ԩM<� 5|Oܑ��m_�(v�1v`�0�ti�ĝ���'���9O\牍j�(�5�$ �=R�n�,~��B�'<�҅X���,w PRR�ӥ!Y�B�	�0pF����XB���Ⴅ������x�|`��i��d�.�T	���[�9�W!�L���u�'��O���H1y���t+�/ ��������<���
�~�%�T.(���"�U)&��m�b�<�Qg��P�qs��<LZ�8� o�^x��m�C?a檓&�&=��m�!	6xLQ�,�r�<�W���X��b��NlZ����B~I0�$pӪ�}:%���U�����<8*8��}�<qt1<D��Sc�?�>̋�n�<1 DW*H�t�e��/T@�v�N�<!U�Ҟ& `낋_(n`D�c`�D�<��C��De��e�(��FG�e�<	�n�`=�ak�ãr5R5�5�W[�<Q�3Y�@����!l�L�SE/UX�<'(��<.
��q�ޠH�������Z�<A���x�&�+dm�>��EM't�!�!Μ�0&	�
��9
Rҧ!�$�?5�j�ْ�O�Dfڤ�`�H!���"`���b��9.c�u#� E�;$!�Dȕ)�X@C@�R�C�ۢ}�!��W��\W	 �����!�$S?$�[�I�r�:l��2>�!�D֔7�����[�5��T��g 0q�!���.'�hB2�
$�:���S����$R�v��1�֧dq�|K����y��O-�AЅ@U�o���RPh��yB��5B(%��h���0���y���2���:SM�/��x0�:�yb'�(i�������&�t�7aS��ybe�J� �`2��.�]����*�y����7�jQh�e�#�xd�g-
�yB�^.e�P0ip��7G�$��*�6�y���o���f-Ю�� �Gԅ�y�I�jK�L�u���D��,d��1�yB/F�!Hd�2RdϾj��q*���y��۸*Ȕ�V��w�c�L���y� �B?��0E�V�Ct�Ջ�����yB"U�"j����bT6�r$�r�Ϩ�y�n�,!�r%����z��4��Ο��yr��EJ�8��<(:��O��y
� .��enǙ>�ܩ�@���[V
�y�"O���Ä�=Z|i�&��H�0� �"O�`�b�X*'��*��8���{�"O�pX�Y�W_��;��
;S�Q8"O*��Z�wT4�&�X� %J��'���'zb�'�2�'���'��'""K�����d8�e�,��1`�'�R�'���'���'c��'V��'��0I`��Sq��2�mJ�JP�g�'���'�"�'�R�'B�'%��'�"�,]n�P�L̓w�	��+��?���?���?����?y��?Q���?I���d��+0�N�n']6�?A��?����?���?I���?����?��ƒS_-xAA׷*]Z�06�Y �?Y���?1��?Y��?����?���?�)���R�f�����6�?i��?I��?Q��?A��?����?!�C.�;ƌ��M �ԩ�?9��?���?A���?y���?���?�7!��]h�:ԍ�}����Fo���?	���?1��?a���?��?9��?A$W�)n��r
mf��A��1�?a��?a��?Y��?q��?����?�E�1;�82�����<i��
�?���?����?���?����?���?�֎]=-��i�R�L�>~:䁡�P��?���?���?��?a��?!���?�B
±	P%���(�*���@��?��?����?a���?���o����'J"dܬ�����LՒ���Q����^��˓�?a.O1���*�M{ph�	����A��;��L �f��'�(|F�|��~b�i��y�Ea�j��������{����C�{����3d�6� ?�0�4QSt=Q�#�4$Y�����\.�
��7i����'�"Y�DG��-�*y����L����_�%�,6͘�1O���>�	K������ A3�����'�~ ����MK�'��)���$h_�7�y�8(��ϖD�a�1˕
<��{�h� I�-_������Xz�����'Dfm�_ �Rg�Ʉ�\!�'���E�I&�M���z̓;V�L�A���@}[VH[�upN1�����>�Iğ�n��<��O�	�pdǴ�Za*ûaN���$��`
�/�	y�,
j$�6<�����_���u�[N�� 2�m	���Uy�������k,�Q�PG+h��I�y��Ħ`�/?1Ӷi�"�|�Op(CW��/l�f0��,{f�[�',"�i�b�[�)훖���:!&ޔ��|���wl��U+S�/�ޑil4}ї�i>ŕ'R�O�� 8��p��,pE�@�g���Or�l=�c���Sq�c�꼱��� u`��U�]�v@Z-O��Dv� �Ij��?9�I ���s��Ҕk�N$��i�����J��K�`/N�3�����	��$Xu�Ra�%kK�>A`!� ��82р��<�-O��O�=nZ/q���W@��;c�I�v؀[�����M���~�'����'Qm �Zo�|��CD���<�4 Єd��2O ���/��H-�$��?	��R�5�ن#�t�ЄΆ��}z�g_&�yB�'L�	^y��)Շ �� ��C)B(��j1O�4l�'���t���|����T�S��D��8�bI�V��<��4J���'G4*#�i��$��?�`��s`�<�0h��B����G�}��� W��"��O6��|�+O��Ċ$|� cJ��0�&�Q��D-���æ���/�Ic�t#"��y��,`�Ey��7���tyB�'���9O�����3=��{Tƀ���he@��"�4U��C��6O���?)
4E�!RLn�`uMNn���u!�%1t����\��<CW�-����B�P�zEb��$k�6~Ab1�h�/%0$�ɔ���p��ԣ�~M3���7`N:h�d��}��6�1P����''De��i��>c>�}��
=ugL�`f�[��cV��4Z�Д�G'���t���P�9e�A�!h\�8��J� =T�;Q�S#K	�ibD��ti�[�)a��SWG�;\4|�0�� �����S�����]8 �0�C	G4"�Q4j{Dh9:E�b1�c��1����� ��u���	�q���9�a��%x���#'Vc�v�ѡ�͘7�'���'m�T���ޟ�@�{x��g �0�p�1u�(,P������	֟X��џ��O�~<:Fkj�k�!�u*��(+�h��W�L�UG�I�\�	����'�b�'�,ʨ�8�H�M�uL�/]��ā�i~2�'P��'Ѽ�'\R5R$���;��9�V/O�(,,aG���|ƺ7��O����<9���?YwȊI̧jÖ|���B^dX��6N�Ľ0F����4�?Q���?��d�?��O����5�3EF� ֘9�񠲫��M�)O����Od�����O\��i����AðB�f5Q��I�#6Ve޴�?�i�bxIF�i��'�?1��G�I	M���

��>Mh�h����#�26��O@���C����|���&�"���:_�m��,"˦س��cӪ��JJ㦁���d�I�?�rL<�'0e��S@_�Sv�谠�ȭ&;�a
U�iQ�x`Z�0�	���3��⟬(����p�����7zޔq,�Ms���?���H��E�ԙx�O���'/"ȸ��{���Af^�V,� �T�>)��?��k@k��?Q���?�S��$�\=�hzF�y�K�t����'�"�C�-/�4�*�D�O��$�b��M��"w�AqbI��y� LR��i��Ҵ��'���'"_��0&�	m
�y��@J�A��\��1H2=�N<����?i�����O0��D�? ����AA&on�E������S%EU̓�?����d�Ox��b�?U�T(уyJ���l �4+��4�g��D�O\�d'���PDja��6-�2= �)��Ƈ��Lq����	ޟ,��~y��'Өx@R>��I v�-�"U0A%�H�Y1Ў�Rav���$:��ڟ��Q�I�`��OJu�l�(;7bu���)t�����i�bU�������O��'V��
X�8��`��n\��x�ôg�)�
c���I~C�8�uf9�~���T�>����!�R��ä��]}��'m��'m��'���O�iݑkrO]�0Ԗ��Á���U��>���(xJ�CG�S�6�)E�:1�����cD�7����	�F�N���OT���O��ɦ<ͧ�?9e ���c��O�[�P��,t=��JW�z�$ҍy����OXT�I�1h2��*��N������˦��㟈�	�S�~�����'MR�OJ�q�� /���&�<'��D�AG�c̓s�JD(�����'���O�E9D����������"e�vQ(��i�r'G77 �	����ş@�=�kW3�T��#�l[���5�i}�c���� �O.�D�Od˓�y��J
}�lU�C!�#3���"$@�T���X/O��$�O��d?�I� �c�5dZbE���\3N����f�&����Q�)?���?(O��D_,�2��%����IA	_�v��׫Ţ ��7-�O2��OZ㟄��8.�h���~�4R����\��p���5@�t��dS�\�Iܟ��'RfV�S�@�eлIe��ٿF���u���Ms����'���T�` �qM<	��V�~���FF�h3�c��G��y��[yR0O���c[>�������өP�2L��"O!' �����%rvҝ�}b�'�>a�f�4Ø��I�P9*�bp��:���B����Iß@ �˟��	�(�	�?���uwo��V�Ԩ���7N]*Q 1G����d�O����m�6F]1O����i��~U�q&Z�Q�@�ӹi�@)�0�'��'{"�OB�i>���>(�%O�0#�Π��J�*�ٻ�4t�&Q⑫	f�S�O��֒M�Yô'SC��xC���\}�7-�O����Ox� ���<ͧ�?���~R[")�(@g.��B�jpH��7�Nb���0*S��ħ�?!���~�O�� >L���kH�;��A��䞎�M�n4M�/Of���Oz��<��/&�H���+5� %���		\��Bb|��Ɩc~��'��U����(~m3�AӪce� rc�3L�2��ECuyr�'���'��O���[-Ҙ8�h��e�~�J�@�[�"iV,"~�I����|y��'^�:�ן��r��9N_\�a gֈl�)���ig��'m����Orrs)MKI�f��u�p qB*�  �	{Rő�����O��D�<��f�,�,�����:CYw�T�
ק�2<�q��4�?�r�'L���ǃ �ēf���B�7"���XΒ�>��n�ß �'��BǿXH���L�I�?e9E���r�Xy�i��&V���ָ��'��b�i4���y�O���[CK��$`#�ӕ�� 0�~ӊ�H=������?a��?a�����^E� ��EϢpYs�-�6�^�,��WA��ZA?�)��l�Z�"u"؅,HP�� Z�V��C$Z��'��'���Q����k5�NV(f��ņ����u�Y4�M�.�m^L%�<E���'OXU �M��nj�\C+2L[Xl���y�0�d�Ox�䀣[�8��|���?a�'N8	;Fo�#:�e�E��*C��k,��B�5I|����?)�' (�0�Rj@<���'I�4e�ش�?	`�����d�O���OR��9s��r\t�;�
�x���2���>Ai�')w�8�')"�'�	��&G��~1���a�
m\H��\�^���'wr�'�2���O.�H�����y�$^4{p(K��&4[��1��X�Iԟh�'�B M1ON���:�(�{Pf�<��7,� 0���'��'��OX�dó#2�=���i>�4:1�O*k(��X�͝��0��O�d�ON��?�D�@9���O��e	�>Jj��E�\3"���¦��	U��?I���0�2u'�8Y��k���c܈=�Ƽ!��i�RX���u��(�Or2�'���Q$6��
Ae@���+��Y(Gߔb���ɾ	d�9��;�~b���#rIHዕ>Z�q3K�w}�;O�pP�'���'��O��i�!�J wI�酯��QC�ЊW�>A���=�Eh�C�S�m[
A���+��@�0
��n��m�lcݴ�?���?����'A2�%9��E���ʘe]����;�6�L� �����Ob��Oh�I�OX���OH���b֦�h�A��&�v-�Fdπ�V�m�ޟd�	�����ٔ�M���?���?�Ӻ{�I$����Ï�/��(�C�Q٦%%�̰Acp��'�?���?a��)j�0�׬�� ^"�"��5����'�8�P��kӊ���O��$�ORu�Oa���	\K�4"�CU��N@Q IT����kqz�ß��I����ş<��꟰��ɝ�`aj�=E���Ud�@��<r�4�?���?���O��y2�'�"L��N�]Z�4���g?f1)��L�����O���O��d�O8�d;�m�;9v`��r�ǥZ����2^*Xʦ���4�?���?���?�-O.�gw���F�TJ"�,�Cʪ;�|��i���)�'���'�8��5�i
r�'�(D:�M_�R;"�! @��I�S	l�p�d�O��<��a���ͧ��)� �p���˸]Cn�c�ݵ[rdŐp�i��'���_�`�ٴ�?����?Y�'p86\��c�=ix��Rf�iɨ�W�i5�R�Hϓ���Sʟ �nZ6P֥��J�v@ȴkB�")X6��O���ͫk���nzoZş�I�?���ϟ�[�h�7����H�#=�q� �������O8˕��O��Ļ<ͧ���$At�I2���^��@JCÜ�P7�M.Y*YlZ���	��`�S�?!���4�I]�~u�F�ZR��S��A��C�4M؈)���?1+O�i#�	�O@#��>�8�De��`�
���Oئ��	ܟ,�I���)�4�?1��?���?�;����t`##O����J(�ؐoS�I���)b���?���%,��H-��:[�L��d�.dXҼJ#�i� ���6-�O>��O���S��O|M�#�D2W~)�q��+mC8���]��G#r�|�'IB�'��'�reڷ �n�B�U�$qR�V��U�ʑ�B�fӖ���O��d�O���O{��|@V�P�
=� �4霎l�����l(������	��H��ǟ�IΟ��g��M�RA�;�-�ą�e�����a�9M!���'��'"��'���ꟸ�U�x>��Yh��f�
�0���,_
��ࢫO��d�O��$�O|���h���m����k�.@��KQ*$<�94���/j���ٴ�?����?)+O��ĝ6'��	�O��	�
���p
�!�HC%iJBS�6��O����O&��$%�o�����(��b�\	j�%O��(�qd�N�J�b۴�?�/O���(���ӡVe�H���˃S3���αI�*޴��Mf�@n������p���?=�I����������B��!��Od�D,,�"�$1�4�$�OG^$Ib,�=��l"m�8�̜s�42��% ��i��'��O��d�'�b�'q�§�G6KJi����f���۔�q��]#�B�O�O�I)�	�O����Gˈ�N8I��Á)�4�7�ئ���˟X��$�fp۴�?����?y��?��L�Ɯx]Z�Yp捗9X{��oZٟ��'T<�b�����O����OĜȀ��.���a�C�;b�I�#˖ߦu�I+���3�4�?���?a��z��o?i�+�zZ��*V%��6�}g�J����()����P�	�?�I��|�O-�UCd�>9��xkG&X�|� �ī�;LNh7��O$���O���m��V�p��;y:���h�5m�P���J{��`�u�r�D�I՟`����l�	t�T��::0t7m7�*\��.؃k�.4`"�7Ajҡn��� ��ݟ��	��p�'wؚ�����,<"h�i�`�#��ո�L�*c8j7�Oh��O��$�OB�$4V��oZ���I
Z,Mˆ�O�=� ��%&p��4�?)���?�-Of��!t�I�O���	H(n�B��E�@v�SC��i�-xs��O�D�O��$�*Ǿ�n�˟��	�T��	]��\�BF�y���6���HFh1�4�?�,OF�䌞]}��3�4��fK�"є��Ed�V\�GB?�M3*O0��C�ߦu������d��'�F�A�H�����v�')��ii�4�?��A�0�������i�� cqԇ_,�<{��65��;��oӌm��Ԧ9��(���?���}2�2B���C�1M�4Q�e*/��6M@N�|�d6��8�S㟤Sd&�W�Z�8����Dgp]1&���M���?q��A=�[��x��'���O�u����%;���Ҧ34�4�	��i��'�V ������O���O,�i���-Ǹ)@U���b��B�ܦ	�	�x�J K<9���?�(O��Ǝ,;DcI�M�� 1�� ��$`�X�@Q�lf���'���'*�R��x��ލH�L����J^$ D�)u�=�L<a���?�N>i��?q�(Ե^/�h�RU�p�{�FF����Γ��D�O��D�O�ʓM�<d�6>�<��*ɠ!���e�A˚2�\���	֟L&���I֟��m�>�t� 5�ek�È�;L� �b�Xz}��'t��'��^��N|"����J�C�j�n;d원 �%=���'��ğ��	ԟ���ch�P�O���!	F)}����b�ogb�ʓ�i��'x�ɐh�FT�L|����j!Im�Ah�(�3�P�~R��D}�'q��'�4-Ù'2�'2��̷i����B'	�.$��q�	|,�&]���Ύ��M�R?q���?��O~`���Q
G�<�i��� ;1V�xԲi���'�u@s�'�ɧ�O\ ������&���������ش.O��b�iF��'@�OԚb���g�u	h�0�Dj�Y�lɑ�M�����?!K>�(��ʓ�?�.�y��%2�M�Af�����;`R���'GR�'eP���#*�D�O�����ՉH؅z�mK,G
�C�g�<�On��5O�S�������pbU�E�ᰰ-",x0�l*�M�Vb�Ect���O:˓�?�1*�Fɢ4�_�F,�g�69�b1�'a�HKr�'a�I��|��쟀�'W���N��F�<JC��%��p��*ڦ3�Ov��O�Ot�$�O4`�0(������Bo�(b�b4sGQ�T��$�<���?yK~*�C�1��
|���ta�j�����"ё3��'��|B�'�Bk1f�Ӎs�E���KT(�C�٢@! ��?a��?)OZP3b��E�ӹd~�F�U�VwTҐ�Wc�*��4�hO�d�eAN���O��	p�Yb��4�����%/��6�O��<A1� L��O�B��5Ƥ$��s���.̅������'��ŅuN"�'F�~�goF;(�PW�L����C�V��ɔ'�M�%dm�FE�OJ�O�����y*�B)3��m�b��Q���'��I����'�Q?� �U'	>�T5{wO,��:A�ii� A�NwӚ�$�OJ����&��5I'�$�sd�'JO�U�G�J18�R���4
������S�OUR�i@�G�S:\Q���=g*0o����럌s`N����|M�4
CcL ^Q  ��+u��)��$i�2�Ī<���é=I�O���'IRcLC��	��#k��GIɛ`��6-�O #e�^�i>Gy���-�(bI�+;��k��Ҕ���հ:p�d�O����Of���O��'A��8:�K#;6�����s@X|ҵK���?���?���?)N>��?u�ˡw��p#�\>��iÐb��rt��g�H~r�';��'%�	1A~0�OD�u�l��6	𔏑�{��X�O<�D�O��$&�ɵ9�8�'Kun���k)1�<�9���(O�)�'���'D�'6�k~����(7�B�6���QB��V��Ƀ��7�M����%�x�Iǟ$���I
~�Ox�H!�¼S�X���05Wn9��i��'=��04TL|J����!��6{0��)7���]�����$K5I�'���'�
���T?5���\$�J�8(����`��ʓ�����i%�'�?i��L�I8Th�E��#�Q���e��7�\6��O����)�S�$֎���	�䢥MZ�7MJ!L!1m��l�I�������ē�?�t�@3X*���	K̋���hy�v��O>A��
, qP��"t�)�oȮ�ȍ��4�?y���?��g�M_�'���'��$B2A�l���<<5f�4#�	:w�ON�I%��Op�$�OCb�P�hp��eF$|<=�'�����	$O!�,�K<����?�N>�1�FP��S����)���'=�5�'l
)��y2�'N"�'���9k���겆�-�8�ϐ��t������?�����?���1Z� w	�4�TXY��T1��@@��P��?a��?�/Oȹ�1��|����
w�)X����HG*��1�AB}��'�R�|��'�r��.���99c̰h���Z����,B�[��I��	ȟؖ'I�8@-+�)Θy��Q1�S�@��-i��0�f�o�˟0&����˟�kD�7��=f?���!��)��]�1+��7��O�D�<у��k�O���O/���[�>�X�A���p��Tj7���O$������'R¸Xq*F�����/#���mXyB�ר'^z7�[_�T�'��d�7?��T)	=���筞2S9�T*7�榝�I؟rD�-�S�M����ޤDھ%��o�@nZj��ܴ�?y���?i��`��'�� B�S�׫,���K6ƀ�,��6-Cp�"|��l	 �I�=�S'ĄW Z��A�i�'��흁Y"��^���'2��=1�D�*_k��0���*���>a���?���?��F�"��� �T?	/zQa5l�1�f�'�UjP�����"��H3.��%�3�ڽVa�%钥˯a���%���%�4?��?���dN�f�h�z��ƚ
�y�t��`����k}��'���'�B���+\��ロ��`� i�&�l���l�|�IƟx����p�I���y�nUП��-5PJPɣ���QڜY�H��M����?������?�*O
�8v�i�����G�Zp�T"��,�ѭO����Oh�d�O��LH=<�D�O��$�8��lۅ
0�N�IP�V+ %oZß@%�D�	Cy���=�ē>~�����	�@a"��+�vMx0n۟�	dy���7�R���d쟰���.�<P]��9 �S�'UzP!��A�?q�%�b��M��?Τ�E(6t ��ئ���ٟ���Cǟ(�	������?=��56��C�9��A>KH؁h$�D��M����?q%ǉ�orzh�<�~چDN|@P�gԝ`殮x&����;
��M���?����A�x��'3
��bĕaZ�± N&MU\@� ~�ZyI��)§�?q0b	�7�d�Qe�G(L_�`��(�;���'���'w�%��( �$�O,�ĳ��J7H�G�Xݺ¦H�xՒر�B+��-[<Rb�������� I�ĽS�(�[��� �֒EcӦ���8,c�4�I<q���?�N>��-��0h�b��"S�����ժ��'��;�yb�'���'�� '�Q���w8!� �K<���o;���?i��䓽?a�m���9�D�jj� ��ۙn��@���V̓�?����?�)O2H+ �|⇀��J��3�Gu��R[`)�'���'��'���'�z�*�O��a��O�
�6�K�Sd>��Z�D������I\y�HP�)��^`kB	�+t,X�Ŧ�.��<Y��ܦE�	ş�'��'� �k��$�α<�\���#�j��	�H��6M�O��d�<���] X�O=b��5�]�q���Bp�A�|iz��A��Е'���'9��@��	��mQ�״�
��"Ri��Q���ꢬ��D*�AE�ڳwW*�$>�ˀ׬V�H��;x# 9���*Zеp�D|�ЇȓU�p�G����M
�e�" e�Wj�iap挋�f� 'Z�2���[�H�`O�q�R���<��j���@�((����r�b#�i@�<P��a�
P�(���'�D4�\��2J�i�f�h�%i�����F�E� D�\*#-��(�猶9����(�i�4]�ɔ�\���?����?�������OV��Uu����C�-�$�$Ĭ0I��[UbT&W(ࠡ'I�R/�h�g��� 0�`�e˰`�CT�v�6��"͞&9~թ�-� #cPjf�ߣ��	��_1�͈М|��M=�ҡ����4|�J�#%g�V}�n�'�?����hO�� I���X%w&ـ�� D��	�O�D�plI�%���;�m�a��f<�|Ez�O�BW���OK-�Mk�,�''�0hX ��3c�0p�e��?���?��)��`���?��O��ڑGP1��]T$�$�$B4������*b�p�#Ѫĝ��<�K��U�0(ҨM9C� ��fw���#�g\��j��ĮB(i��Y�"D�8��s���'�4��Od�D���樠��}��	��׮{�F�=��$�$rD�dc�B$�"�bZ�O�!�Dɂ"2��R�l�?1� �I�I$���W}�P�,s�����O�˧-u:$"���>m��`h�G�i����C��?Q���?�$�4oU8��ӎެW� ����	.���r�L�8{������7�Q�0Js.��^st�� M�\]&>m����WXB�ɴj[�C`6衣�0ʓ9���I˟t�j��%v�:�*T�3Z��b�)��<y��_�$ـ�Fѽj6L[Ҩ_�SnVu��	-��^�֬��#:hM�(���#DV0̓g:L��\���g��C@�c���'�"�Ƣ}�� ���i��4;��3/�ʐ{tG;dp���D(G��0S1-�"�5���B���-�9S����IC�5���p�ݢy(5J�.Ԃ{��`S���t4�{�'�g���>����2�[��+��bp֝��|�XH�D�O��S�S|�o-nhil�"��;��&))C�I#$�T�ૅ�.aȽ�N�+q�"<���)��A�ii<}S��i�a
T��?���a]*�iL�2�?1���?���l���O��$݈��x	����,1|�@�g*T!��Y�Mğ*������f>k6՟"=u��� D�Sh��v͘��v��@�n�2����Ii(� S?K�?�FzB�Q\p��[)l�L��'���~����?�B�iN�O ��O�ʓ:mp�q�QӰ�T]~���Q%;3N�\K��[�`)`d����?��Iay���(�6�;y�@� �o�g�V�k�di��?i��?��D��?��������kZ�x�j�.D8�ѣ*�+�Є6�Gz$H�j��E
�:-��I4)">X2�"[����3��MB��Z
k,������x�fM�`�=F�He��$$�/����	��MC�ND�wI�܀��Z�n������l���{��~���
6���hن5��,�UmA}�HD{"�X�mu��j7�۔:����U �y��>)+O�)n}��'��I�*(�tK�Nf�4�2h���L�h�d�O���5_�� ��K}��`��t�2����H!_vN�y&c�:��&�VV���	���Q��A%�U	}�=���c�jdx�jZP\ڝ��H�:!��*o�"v�	�c����AҦEc��ԁ�T�ѰwbB�V��4����:�y��'2�}2�٭ P�A����>Hj�ȹ�\��0>�ԛx�㞹N\�B��@ �k�4�y2c4eW7M�O��$�|P���?���?iS��0\\H
��F�E6�|R&��>��y C��w�.� ��>�O�1�b�XdR��ӪĽiC8��1
L�<�L����.\��B�t}���'�����Kɮ6N�$�ea]�*H�\���l����䧁b-O�)�����$8s)�3R��u0"O����h�nQ�4y��[-Vy�s�	��HOV�n�֟��$nP*~(^��g�>sm0p�@(���	�6'xU$���d�I�@�I��u��'���Ҷ��0JS �~
,���D���~bb�:�T�3oP�ayRfO	 |@�C��r՞���5�~2�R!(Ȯ1
�J8jaay��&�0���%Į?�� s�h��*�BHӭ��,jӨEl�?��?�/OLac��*Ax���ǌeU�H��"O@|ۦ�@�@64�1���]<�!Q�H�'9������K\x�;V~� �j �#���$ՌS�>����?���?pN�?A�����X2�d@�ff���uS0�Y�"�4���N�E�dQx�E�*�|Pq�	�s��Wg�c�.-�'C�)0:M�!`�uK�i ��Vw2��E^�g�����4�r@���M+D�K4�P4�A�1R��ȤIE�6'���'i����|�?�O��pcQ�9W6�КfB>=`Ó�hOj5z� ue@Y���+�A��=O�m�V&�O$˓%�h���Y?��	y�db:7$x'^�0��`��kz�ȳ�'|"�'��+U! �,Uޤ`G�0B�9��L�3_֝�[zT�
�K�l�e�2��<��i@�mQ;���{���xg���00�^w���� �1��+j�tm���8��B�N0�~�mKw�DAR$��9@h�#Q��<����>�0ѥ%�d�� ]4'��� |~��i>��N<�֥_0K D|�H�6>:i��
Q�<I�<,����'�R^>)��ܟ����E �0q�`=z��Y8%��ի֌vg�r4R�4�5ZAi�lςI���c>��ԚBS���۔<���+da��ML�05|Pb�Ȃ� {~�Ƅ2��>�� PE;S)R #�蒆�,T�!���52� �D��ɉ-O�O���]�0`rᛁg���'NB����!b)$D�1��gnސ�oێ)	�0�GL4 ��0S�4�?q��
ֲ���	ϊ��E���/�?��t���	f7�?���?�����N�O����8ؐ�1(̟d�a�͟=h@شCX�%���ȇpI��tF{���-%ʼ	���8!VMԤz��<oZ�V׊�Z�B��ro�?�=Au �:Im�ie�Qjh8��']y?ac��ʟx۴Gr�'9b�'��9COf=@ԯ��\��� ӌf�C�ɿ}�D! #��&� J։]�5� ���|�(O�qc+���=�6F�Cl ����[kΡ�7Vџ����h�	3�z%�I���'�1#��	YC��T?����Z�>	��2T�-ϛ�4,Oj����@�z�CG(�y�	� �Sɸ]�"�ӸA�@%���YD�裖V<-"�-2W�	yz�	�yZ����O����� ���+G�x���׊-���O��D.�)����/i��}{E�T�ґ���C�ɬq�z��G�O31�-�s�'Z���Mc�����C�-%�l�P��I����`9�T(@I�X�<� fйh���`V�'�r�'r�-��� �@U`�%��'A���e�,5�iJ3�A�wݖ�Fy��0#$�� �8�'i���A��Ũj���Rd҇.���Fy�J\��?���i-���KTj��U�o!���x��B��O��"~Γ#1��􀝽CD`
hM?V�
���7�ē7w(c��3�|��#�D�1�ֹ̓n�6}j!�i{2�'8哾�Z��I˟<�	'M�j=���$_�~�J��S6N"B0rL��?+���f��8����S���'R<�a��7�x9�GZ)FQ��@ E�&�H| P,��C-J)�W3O?��J�s����	G�B ��3a�͋9U��0w��O`�lڼ�M+������ND*)`�r�'Fq( LK�
��yB�'7�}2�׭a����3_�9���O�Ez�[>�+�ܯ4�b�1"ǏgܪE�a��	�
׆���
�֟|������I�uw�'�R�T�c��Hڤc=�=y�ʗ�~2�&�a}���� .�
���R�x�LJ��~�,�= a}2��r�xj�.�3ej� ��aC��~��S+�?�����?I����d�4'6� ��D�Y��7�/N!�#o�HŊ	"-��b���&P���Ezʟ��2p�z�i_N�@�� �l��%)�҃q��<�U�'R�'��d\YR�'��ɚ�G'֡�FCi��S��m�0DB�)�����'�L�:�%SB��bX� =�,�FO'S�R���mܶ�p>i������l+���t$_�.�\�Xd�3��q%����͟��?�O�Hu D@O��I!�C/I���'a�y��U�XZ1� �M uy^�K�'C����۩��Dm�ԟ|��J�To�Db��CPi�OH��y�ƓI��"��'���'z����'h1O��u��#bGJ}
Q+��>��<�NS�O�$|z�+(/��c���S�dۏ��A�}���Ӻ;�|d���p���㥎E�u C�	Mb�8��h�Hyl���g������Y�	5\@H��K]Z�����ӣ�T�	�q�]�ݴ�?A����|���D�Oh�%~E�t�Ư�37�X���I?=�X�D�Φq�<��OB�K���/�
<��m�(�00-Z!b���6�)��X���Q�	�hX�a#��mF(e��C�5/u����MS��iZ���Ob��b
�f���6A�(��=O���)�OA�5�πL�5�2K�/Ou��3�	��HO����'�X�Q�Ǚ�8�7,��+n�͐F�'����:C����2�'�R�'��wݽ�	�d�$/ӽ!'�h�ªJ�a�0H`��۝�?�@$@��H+5ʝV5j�3�<����Dڑwp��dG�:|��5���'b�@��
�zd�ꄭiF{���m�ȼ��LB�6Av=�DB���~2��,�?����?ًbQ>e2�MǢ  pM9�(˻>�āJ�3D��q���y��Eav �gp5�����HO��Ayd�f`�7-Y� ��u[�14�� �h���D�O���O�y%+�O���}>��C�ԭa� �3�_�SO�{AH�#\%��ٗ	H�k�0��$�v(0Ѣ���� P|�G'O*V
\�[<w��])S�'�����7�)��i��L	$'P������H��1�\O���Oj��'d5��`_�:*��c-\Bl��]a�#ƕN�K��ǧB%|�̓a��	Cy���6����?q.�H1�^	�9jb/��s��5�b+�����O��ğ�HRh �1���ʥ+!�֗D���'M�\t1i��,o���kȹ&B��Dy!�z���Iao�9Xz2�`����P�S� �{2����S��(O2�j��'N2�� �)EI��	e�ÐJ䖭z>O~�D.�O�Ա��ب	찤�6��>9}(��'s
OȽ"��G�\q�%5W5T�ð6O6�H��T�i��🴖O
�ŪB�'�B�'��#P*W��t0���g����1-��5�
��GOA�B�S�T��'S�}	�a�LP�����R����4�gl�y�Ÿ���S��?9dk\�&'�P��0��L�u�
�C�ĵA����k�n��1��y����7n;|v�`a�l�X�	Mx����Q�+��p��/B>��U�/�_��H5�O(��(Q&<�QD�6d�ji(��O��D�3qZ��5��O�$�O$�$������?A���-=���J@�Z���0(T��B?��K�$�v��d )��|�f�-P=v@c�J;)�����B��{
��Lq�R��h�pP��?G.������	ğP$����ş�'�x@��S<H�^�I��J̭��'B�`�F?I:��㎞+�:ͫ�k.�S��W�`ұ`\��M�ₐ�pp����IN�v����0�	��?����?���]�F$���?�O�JJ&h��\H����̖U��ȫ�i��<iVX��kBx
�{�cH��f(���HH��Lr@��%5��M[��Ic��g�'	�t�����K{�8s��Num*(�QE��f7��O�ʓ�?َʟ4`����i���Rh�Z�%��"O�Iv�(nP�UK4
܃?TBQ�?Ob|��'p��C� |�p�$�|⡎��YF1�g╾MȬU���U\[�=:���?���5��陶gT:����$X�}�b7]>)P��C��i�^�*=R]q��>�F'4�Q�G�g~>e mR�T���e���u ��@Q�\�����g"	�d�ʾ�(O���u�'��6M�i�W憜(��ʖNRP�*�N@�p��Γ�?��#��iˢ�<ha��F+5>�E��ɫ��F�\QG/H	n��a�F��B�� �1��Y�\��L�(�j���'x"㉥&�ri��ұjSV��`�	%"8�����@����4���>*]�qT>1�|�I"+��t��
ŒG�ƙ+�o�;j�p$*�,��<��HwL�%5�$j5i	{��?!#+R�*�y�4�3@�!�	2�$���&��%�<%?U��vy⯜�i���Å��Z�9�K��y"��
GR�0�7H��N��|��ѐ��'�2.�N��I�[�������z1Z��PB����I�4r��Հ-\��	���I�R_w<��'8���d] F��0�(ɩ,�h)�4OT����8k��E�8џdK��I�]�4�Ze�� �<Ty!S��H�i�!o�^-�!T:��;���mQ�E c�I+�y���� �`AwHɿ;�D��cŕ��~rf:�?��i�Z7M)������үlI�t3��^�,o�����@�%[!���O.���B�8,wԥis�^/X��A�A��ɥ���0������O[�5@��ڠa�"O�qI� G�nD��8#�W��qbf"O�á�O�3OhP���X<���"Oz�#@��(\�p{G�S� ���T"O��� [�x�p%@�[y�Āu"ORU[2��>���Ӵd�(0]N��"O|,ۆ��V�d���.DƩ#T"ONQ�PIӆ8y�)4(E2%X�"OX�J��I�3Vv03@�3	bD"O�th�B��%|����� �!�lM��"O����	���E��.��,3�"O ����0dXi
ƕ������"O@��(E���麒�ܥ&ޤ��S"O~�+�)UA��D��J�VюyQ�"O�5A@��L����
�m��Q�w"O �S�.Je�<H�����"O�m���p�.��i��"�K�"O��{��O�-9'Y%��E"O���!ݤ;���+#��!�X�
�"O� �b��(),~��@$�y��}�U"OD��D��A����A̓�ew�(v"O.< ��]���嬆,s\�t8�"OX1&l�	}K��*�,�%����"O�rSΞ��F���
5e�X�8�"O�d�,�>K E�S̸n4H�p"O���j� R7P��G�Ĉ��@��"O6�9w`�3�s1�D�L�@AY�"O� �01�ᄘn`��H��31m~��"O��	ui�&s� h�'�>[썉%"OF-�W*ˠ@*>��ԥ�M��9Xs"O@�(PjZ'@E~aB!$&s�a
�"O����R�Un����5c���"O��c�뀍`�.�`2ȃ���x��"O���uD���J���e��Jf"O��aE�JJT�H2lʁ�@(�"O^t��Z��b���M�FI�G�U�^O�3�MHY`�ِe$��~��t�q`uM@��m��-��8~M���0D�|��C+��u�(�+��h$j>)`51�Ӱ�Z@���C� Q>�O�1�F�M%&�8�r�B
�9�E�'�R8b%
�&C�� =�H6��hQ��'�>a���+͡$�����
�P��'��h�doF0'lM;IA"G�H��yAQ-bǴI��C��vfw�ƔӘ'��xؕ�B �f=���?����O�u���֦��1�	�Et���J�I��e��_���Y�8O�t�
��YV��'��$�H�FD����oО���o	��)��eTo�|���'���k&�چv�� ց_�38`��'J�M(g�2e�t8����'��S�2M�L��h�r�uHvÈ/`�d8�b�'A:%�����D�o����0���#�����Y�@�����и'B|��'c���Q�gC7'��OH�\� �f�츉�hоp#��S�y�`��0����ܧM�0�j�Þ��y2J�u��]�$I]�D`��
�$;�6mq�" �s�ԔE� 	� I�Wf�67��8#Q>��?y���1��l��=U��	 �D��~�S7�ޔX���Q�e�<y���;q�mɍ��-ȹV%�pal�!�0A��L��V��)�J["SF���'����	�8@���DÓ֘���'3��� ;C$=�e��,��OGf��#Lm�b��10͠P �J��v��%���'�({!NZ
S}��b
4c���JX�v�)� ��Q��,s`h�;�y�m� �j�[�����$$])QЃ͈���'L��Q�ޤ>x�A"�.V	�1O�@ �&G9MGȱ����_��L�?Ob����M��y�abښR#����A:D~�3Θ�Y���+1*��P����2zk�ʧ��'<������(U l��+D�^�PEzC�M;�j���Ӧ,>B��'�������h��6Er�֑k��P96�S5�8@�dnB�e�~<�2 �#c>����+0�T��eL�}J6!�wX�F[�DD.R�Ě'd�87��h��)�or�H�p�p�Q1.�`I�&Y�T!���$�>U�H�.I���d
�G:WL5�t�0{����3��qSrU�'��Q���&��l��O�b��3���'z�L�Y�
�sC&Qy�	�-�g3��2H��X ކq�+�ܙa������l	�f-��f�^��H�!�G��'�v��3N�L��Y�'3qx�_/Se��C����M�����0Q.�y�4x�Aτ^P�I���S"@��?���s EE��N\�ǝ�L�|����C�D%���ԅ�p=��o^AIh@�DM��{}.i� h�"��S�6
Tt���K ����7YJ���$�b?�s�GLaj��"�Q����d�'B"Ղ�M�)^*��I���Gwh��SD�>	b�)��Jȑ7�03׮�O����(��<i��w���$qj�aK!�X�[ט�iӬ�b�j�poB�>��k�f�  �E�x�#�0NE``B �F�U��L`F`ħ9b7�	H p�Ʌ9�8�b��͋�.
�&�*AH|�㊲���p�A
r��tK���<^����5��x�y֏��y:6
`bB%�XS���!}8h��kӀ@&67�Eo��c�l�'*Q���·O�&I��M��H
��5J�}��b��}��zZc����c�[��L���]�L�t���4uxtC�y�	?5�
<�p�W�;��� �ns4<�F�'�:T�E��Pf
izօ^���)�0��&k��!�
�H7(iɲ�O��>�҂���(h˶	�"OӬ�It�0CX�V��w�&�K�#���Ao�L���W"w��%8��l�K����'�$�f��t5���LiF�1�@[�~���8�8dH7꜁��wn-��'�:Y��+[	g����\Y0�ꃦ�'^0��2�C@�-�(��4Yu�t�D��RNb���|�'�f�r^�d �0�m���]�g�
W���ZE/��=�1'~�ё�W1��<{a�D(j�o�=2�Ԋ�FY�c'�
A�S v�:��'+X�X��;r�|���3P�h�(����Pg�;ð<i��M+R�$��5�ߌ32�)�0:<��$n�Z�y�m�0q"���/+j�@�B���\6��$�8�6�BH��J��ܙ���n��'$@��#*UxĀ��̈́��SAr�f����x����e��QeD#[%�ْ�"��xb�V���c�7:a�U�r�8���\�xs��&���`g�,Z����g��ۼ;-z�4����T��*��'*�~H<�G�Ån�}��CV�F%h���	0>:]Zen�5� !%kU@?�]w+�M����b$d����S���\�v2X�b���v��c �(ay"� )U��	��Q8J�@���FVn*���`����bA[�u�����+�f�i�	6���Z�c?���t䵫2��R��Jb���b��O�3��-QMz��F���2�&���J�?�*R�6N�䨚dg=8i8Ar F�TY�n��	�Ё��G��|
� ���sꉄp�Mc5�4+$A�B+�<z/�i*���S�M�BH�j<���w♤F��L��?U��'�pH��aޗ.Z�3�i��N �	�'�bxI�b�A���`�C�3wi�a%M��$�v�X0��,2��1�N�:�t֝�]�M"7�>��O��M3A��'���+s�P�j���˓�~h+��݃h��]͜)��CF�b��<���R)RI�Pz�A4�T�"rܳ/�.�'��>7-�?k���X�ի8�!���X�b��'�J8@&琓vMĳ�eŝV�x�i��n��Y��n�b�0K%�_��I&730�ďI
��y��:�n�C�#�SBZ2�H���� ��p�#��q��db��)�E,Р"p��q��\���Æv�I�h�3�PxR��L�0y�2�"�0�f��$�`q����kK�mc�B/%�x�I�fݵ�d��2 [���4JZ�X綜�Q$�=z�$�눰ʰ<9a�X�;��=K)�1!FH����'�j�c��ȝ?�~�Zc�C(��E�65��B�޿:?��h����ͨ1G|��RID4rm�-K�m��ē(d�Y���J��1�/?�*������T�$U¡�7-���e����.��h� ��<�b�E�|��RƎ�C���F�kFZ��ŏX5��y:p	`�$����)�$i٠n�A b�N
<�Vœ@A��x2�,��ͫ�o��i,�#��L:>�� !Μ:}�x��*�<)K?�$e�����O⤕Q��;	a@��'��6j���˓7���G #���)�E��r
 �a�˘�����%��5)���'9��9D�b.�dѿo� �c���O�-P�M��}}�Ԁ��D<~�L�%�xˉ�8��u��CƛEj�(Ұ�_�Z�q��5N�&d�q���t>00z��P.c�l@"��Z� �C�3<O�,cfgگ+���0�	��f;bm�w �&�����g�(s Hk�+Ɩ>���yJ?�am��F8,<�#O�)(>-�#<VQ�i��2�Ok��>	�l9e*Pc�f|��A�GS<�DĆSܓ�"dϱ�h���'���$� aF���~`[4�o�V���C���²`�r^�� 	M5�l�M�.����u��i��=�	�KQ���O>H
U�icl˧a>p\��MJ�:L�؂T%��'-�0�lS4�ZZ�'�`-ۢ`��F4� Y��T�vc���Y>�2������J�u&��jޘ{p:d(!�f��\뵦�4X��w^�l��؃��`�VDH��/7�ĨH�j�sK�<`U�4	�pgG���Vq8��z��I B4��Q'*D����pA�Q�lA`�:7$Z����O�b����#`6��pE�'�p�f�a�V����Z2Je�Չ�D7���'Ծ��f^�L@�PQ$b�E�Ɣ�G�S"j%vՈ�ܟ:p{tG�j�R4P�O�`{(Q0Q�'TB�j��A�Q�d�H'.񨁵X���+��,X���v)��
y�ѣ��������L�Ⱞ�F�b��"�H3AkfˇXlf=h�_hp�eIʸ <�s7��%ˉ'�x�fH1Yʖ|��-.?,HX>牍B�\1�bZ=,ؘ��JW&8�� !�ˌW#����X8��E��"V{L9s3jKhP���$FNT��U�E�^88��I�.z��1��Q�`1Z�Z0㕣Z����;�*OH9V���k��!�$Q�2��ycgX)~>(!P���?�&�ȪS�����"bU�I��(͠!2��?Y�g�
R�<�Cu�_2 Q��IM^���'�p���$f�N�5R���
�$�� ɮ��y�
P]�9VN�gᶤ�1� �ll���ɑ2$9	�-U�)��d�2��L�梖y��@�eV/Y�\�bCoφj&�Y�E�`���7Ϝ|�+�v��1Är|�M�3�̂�vt�B*$J1���|�'��unQ��:�	�
�R%��{�'��P4��:`��\���^�N� ���Xa;ȈCvMη>�|5���O����$W�}�W�G�*8�X`��U���RI�e ����Si��o#|0*5RS"�LDt�Ru"]�?0��I!1-���D)Q/��1X��E�����4Ђ�ku�ثM����A.��iH%ؚ���ؐ�X|8�Lbq�u��Ś)B���dOE�xM`u�e�'J���OD�|m ��D�{S�iѢ䄬�ħM�~����^4:����H#.�ۀ�'|O�5���ӟI�n��6�R�rԘ	qs�[���c �[ڦq
ӎ�,�jX�nd��H[L?5"u#]BH�����B�]�B�iL�.�\�X�M�1K�f`Gz2�Mq ���D5+�J��"�����mi<MX�%IJI��w���17����ҦQׂ�@�x-[��
�)�,�$X!� ��K��#V.��XF���5CA�R�2�mv���R�Y{5v�@��A
�̨C��@���äM�5ST�y Hֻ��-Ҁ���%����M�Gd�)�M8؈Z��+O*E�=m��H�o;6|r�B$x@0��<1��C&|H ��S��ͦ� �ÄN �w��q���ܺ!��[T�T�L��s��'�N��`��s�� y0�ʷ���у�ď2wj
aMo�6t�#U=9r ��Ѷi�Rx��Фj_�	��_���@�ʋ<�?�5�	�l�҈��J�
W�X���z�'�Șw�U�5�Tq0G-^�kR-b�OV�$K����nJ�M��űlT�I���d�[�Ed��� �O>oIF4��C.�b���ET����GaN�*�F�l��sW �J�ó~8�kU��XD�b��+խ�
\L�8z(N�0kXt�D�\;D�Hp�1�IF	�J��U���}��R99U�8�f����.��OK|;.��?ioƇ6��M3��撚�P�>i����)����@c�,nN��H
#oR���$,^�mC7m�7��! �#��>�0]{4��P%;�j V4�ثwҷC{�F��`oJ�AD�W�?a��`�y�����'�,����вeT�\��F8w�v`Q���*~|HA`�jڮ��D+�<�Y���+�L��iF\^4X�3�M��r92%ɕ�Yv��aM��|k�5�t#'ړ|�r0�.��.��a�gB��%@�oZ�B&�$��m�LsL�1�X\y�O�~ �q%��0dy����1� ����FZ�V;*myvNZJ�3%��*h�tk��"�OtA��`�ci��(c�� Z��+uI��򤍛N�H�ׯ�'�"���Y�9&��OuJ\̻5B��p%��RcC��2$��Ć��d^��X'[*_LtL����Pxh���y�'�0łN>a�k����K�5H^tɁ���ϟ���=k���I5�� �<���N2�O�H���A�2D�s1gF`Q�a�Χu�~@��[��81��,�>���� �"�G{r��u��o_B�(�� � ��O��ɚ�=�8��J�"� �C�!�):}J4��hO9,��4{a� "R���ׯTX���dF/[�4�ZVd��X���ʰ�:r�!�dԆ,��	c����$y��#5�!�D��NM�ㅆ�7F|��s��?fv!�2f�@r�P3K' X�,S�J!�䆧-��īG)N54��l�B�!�W3��d�g�����1AU�r{!�$ �dm��Òeȹ5��5���υx!�dѮ���+�����@�J�]�!�̖0]���40+���[S%��^�!�DR�T��ʋ>kl�x�[*!�$L�*dH���E�]�� �'Ą<x!�$��႐���
��|� bK^'!��ԕ��-�@�8I�V�Ae.��!�$�6R��"4OM�B��,�.�!�D7�q8r)�53;|4�JG4.4!��ة{�vQ� ���L�h�p'��H!��^�bwGO|���b�ܨ�!���!e�ʣH�EH,`��G��!�D�/R}����ڲG0�ceL�!��KZ��<Z �
�EM\�)%��Et!�Č,hІO@�{ELE��*� 3�!��� y,��Ӓ�Ԧ$(�գQ��&�!򤂁R���EoH�C"\��	_)<!�$�V�tq1"&G�c��ZG���=J!��$#B�i��t�Tu�G�>G!�DS�^6�zw'�/,� ����;G!�ώSђ�c���� �QҀ(V�!�܏<S��BC��%^��I��[2!��1� �{�iC�K�0JҤ�v!�8N��Y8�K��pE���b�B"&b!�d:�FɁWN&UO����/�9>!�d	P�8��Q���ʔZ���4L!�Xm���F�O"��Aw� �#G!��O<�e�����A<!��O!)/\<סb���Yg{,!�d9o��P	���$��=(C���&!�I�J�P���re �R��m!�DUqJ�2����!������ԵR!�AVZ.0q�-ߘN����4�	!�
?F�K���\^���b��/!�DL�U���Y5EG�~G@�XG���C�!���J ��c�Z�X0N���	�?�!�D[%b�L����=h'�U�V �
�!�ò[u,x� iV)K�j9���56!�d��-~|sFJ�/���@3��g0!�Č�4g�1����( �8�� �!�$�E������C�Ut|t��⋶2!�D@3\}����fj���_�<!�$·%�*D1�l�
+�)3��.!�d�%c[�����G�^��SA.
�!��R�Sn1I��kfH�u��a�!���Q� %:vEǷ9�x�e�:�!��/��a@�/�+V��D�P*�C�!�$�����	�1m},,$�X�!�$�)����׈�=��	*df��p�!��-R��K���'g�f�k����!�� ���"�]6:���C�8*@0�R"O�]���߫�x�S2Ձ`.\�sV"O M�b�µO8@��U�D)��
�"O>4�V�!��k���&twh#�"O���j(p&P-�SC�'X�<��"O8��2n(��bU`[=`�؝C�"O���Fb�n����y����1"O���CM�"M1p4��ωh��W"OZ���J�([`\�R!�(y�|y�"O:���O� L��X�i�u��-i�"O^�y&d�)
��k$*34.ll�Q"O���v(^�W{�y�V	yp��""O�h�x@D���E"���{"OH��g�S�fSPYp��x�"�`�"O��@C���p��bJ2�|S"OD�{����C@�H7C	y�XL�c"O�h��&
?7��'%����M�p"O��y��FU�5��)�4z��2�"O|�f��83:HcUh�?�X	p�"O�����Z�l@H�π�(V"O���+�_�H �$F)����`"Oh��CƸ$���������â"O�� �M��}��5��#&!�""O�<S��d�X�K��;b���
q*O��2��3�Jyu�BB�p�'���C㋞=b8pE��:?��9��1�S��?ah�0� i�΍H���j�v�<�C�A'
��-�B��గG�W�<�mUKp�1&�Ş8!�\���U�<�o s���h J�R����lx���'W�DXE���R���p�9�=)w"O��3�
�
��E�H�tp�M���'���0v$���K@=z�Ɓ�b�K�bB��)�@ur��&a7���p�C�j��c�@D{��t���H�i@�(�1[% �����y�#ׂ�X4xW�Z�N�(��߸'�a{"$�`ո@�9QIı�6%�%��=��yR#�n�f]��B�A��I���Í�y�c��̨#�Q�>cd�%N��ybIVu$X���F�/�Z�ȇd
 �y�f;�(�dkέ/x�q����y�����Kw
M�~T�U@��H��y�I�"H��uZM�<��#�?�y��NA<P��p�]&��(��eس�yR��o��������b=r`g��y’iL��$#�lx}3 �y���E�p+Ĭ�/u���E��y�MĪK�,��2�N\�$�B��Q,�yr TkS��H�cR#MI*8j�N��y2+�$%,�QF��7�B���o���OzO@�O��̐���T��`�b��=Y`��
�'V$@D�ܰ5Q�!X��`��\��'���8b�a4L��4/ֲVR��'��V���d�0�
�.�HArD����y/F0�:ѫVb�KTvX�dm��yr�
'4C� B��,A���� ���y�g'MzF Y�&L#>$VE-�y�
h-p�C!�P�/��q�O��y�l�^%��ae]8PL�a���۶�y�lNA:�&ْFW Q�-�y�D!=J��р9nz����ů�y�"��A��8^bQy�鄺v/����:�8���@ɐr��hW&�*d0��ȓ\Sr���,����@�!;�t��S�? � �&T�&=l��)Y)5%0��"O�Cm\27�eJtg�"���1"O��D�C�(JUY̛�t�f�aR"Oެ�wj
FG�� �S�qL�k6"O$A����`�Ԁ�JQ��=��"O 85JN�T.�@��)��m�8��"O��K�B� $F1��N��`�#"Od�ӃS��:C�,�*�:2!�$I�Y|���EM
��,�cӲ-�!��(�4\q��;�r X��ގ�!�R�vG��q�K�$t�@PӒa�'?�!�Č5=� UQ%�@A�����*F1OV�=�|z�ƒ��~H�^ s�� Zį�K�<�W����T�;��<n�*SHDp~R%�>��!�f�K]!t����vH�1q�-��>�4�*rAN�d�l���P��*W{�<Q���y�I���'`�!Auh�z�<�p�Dm�N�#��&W��A�Fw�<��	�
���qT�F\C��l�<�d�O;�H��s.�$�P!E^�<9@�̷i���� ��|7�|�pD�u�<�!�3e"�J�ȉU� ��[]8�|'��q��5��8p2��?b��r1n-D�h+@�W�l��(e�	-9:$�%D�\x��S�L����M�< �(q��(D��A+lN>؃��'ES��‧4D��q� �i��yf2V�$���0D� ɗIҍS^��$J��H�R�Q/.D�xx�aU*XC<xk7���B �5 7D���ϖ**Ӿd8�_�G�.4s�6D����OZ�(���2��)fz:l���5D� C��I�"�c���O�ԕh7�5D�4r��y��,3WJ\�4��2�+4D�ph� ��%�B`xM��#��a�f2D� ���U��LL�E풽)�:`�C�3D�$�lF�Px��&m�5/(x��3D����eث������^�N�ڷ�3D����HM�k�U	W"0�pp��2D��Bv(_+'�j5�a�� x9%3D����
�2Ky�x��K��B���/ON�=�`.��m�^����=|��@�CI�F�'�yҮʪJ�x@�#���(svY��
��y��i�"~��)�6
"��g-%L���PfD�<��ی<��Q��[O^ 9І��<Ѱ�����X��՘X�Zm�3�z��<�'8��c�O�h�!�g�[P����'����+C!ex��@G�Qq���' �Ъs� �?��I˕NB e�T*�'
�PC���;G2��DNE�Y�h2�'�Й��&o>1q��(y2�t�V�*D��)�YZ��� ]��h��#L'D�Hp`��U�t1�-&8\��G#D������~����#Q?� �#7D���r�%a���YR�+L��5���6��hO�SY���e[K
�m��E��
@C�I%J�I GH�WB�� &t�nC�I$�޽�'�HE��:&��[BdC�4PG|t�@&
�4]��! �-)jBC�ɹ�z��BhN8=�2dX�,�����q�$�$ ���(n�T�7�K�M�TUiS"4D�|�ԁY�i����d�4�
V��OF�=E���"'7�=t�O. ��  ��b!�A:w;l��F?:z`kӮ�.�=E��'�0lI��Oq���bcE�|��aR�'�� �-z2R	m&�us����'���d"64�|I� ��w���+VB�?Q�!�$=�و���q/1( 2�S�sT�I�"O��ٴƘ.W�l[u	�����'�O��0Gڴ0��i�A;
p��8�"O Bu�-- �aD�;n�M�e"O(ݪ��@�*��dρ)��x("O��t͘<4�z��زy���U"O���sb��u(�J��5o���y�l��Y����,�*:��i�d(�$�yB�B'W��E�!� :`����lW�y���>s!�u�$	˷JT��Ȑ	�y�nW�,���J�vpdqf�$�y�kL$S����u@���z1q�6�y��	�:��|�=�dK�%O�y�$V!��J���H���@C�&�yn]�D���E�L$ �g�̳�y�mL�g֢��L�?�Li��-N5�y�XB��)����
<%�郇��y���|�����@Uh^T����.�y"H��b"(@�ϝ�,��Y��gů�y�;U�ea`*�.@��#�E�$�yRK�
VB
̻�b�P!��XTc[��y����9��D~f@9��"Ư�y���6|#��σu�M���*�yR���$�R!�*E�jXUMA�y"� %�݂��C��l%nï�y��D�K�H	xCoC�B�X�qET �yr�Y��,8�bNL�n4Ybe��y� ��w����˓�l\j�`��0�y�)�(@�x��Hy�Iȓ����y�. #����1�Y+E��s�X��y��ͪ2��+ģ@	j�zб2�Ƶ�y�e���\ n��`
bɋb��yCI8 �����L( r�ά�ybJ��rh\0@d��j����y"�'$(��`ŷ9ց+Ō��y+ܡl�d�Ƣ��^)Б�# ^�y�AiE�5��(.P|����̽�y�"� r�x�c�+A�n)p"A�4�yBB��<͂}:T���#�He��!ɑ�y�邂h]�8@#��TP��`�y��N/b!����)��jd��yrJH�^#�Qس�����)�y2��D�fkFaD��͒!�3�!�d�*�q�2�F-nB��S /r!�Y�5 ğW��I7o�0K�!�$MW��Ѻ��TY�d�P!(�d@!�DJp�T�X��Ȇ���c3��
+�!�ŹF<�0�I�0���27�!��3�R��� ^������!�d��U�x����2��}(Q,��	9!��R2X�d�1�J�>�@�9�+�3�!��	.b�f�A�KM�)u�Y�����3�!�dC%��Qp�`d�y�#��I{!�Dӗ��=8� !;�V�:�쌚-C!��G��:߳�J�@�	Z+!���}|@ı�L޿�Txr��&!��rn��d��~]���wƇ(e�!��?2|��ZRm����f�!���z\@�
�;)�b�:C��#2r!�։3Ҥ��lӳ+ǰ%1VO^� <!�$�0:|)��зqU������x�!��,Y�JG���b	!b�!�� &�����LΝ�`쐂w-����"O�h)EIP%q�rE�vk��V%�0H�"O`�)J�S
 ��p��[6�d�"O���ED�^����"�;H��"Or8���B_���q�O�i���R"Op�S�l��&+H�r̒�*��t��"O\���$+��]� aߡz�$�"O8���`�#h��h)C�ډOk��K�"O�� ���i|�1����9m�8r�"O��Hʣ-���ITiB4n3xPÃ"O�cgH�9zR��J�g�b���"O��QC�6A�"m�S�-V��r"O����o%3���F�T�R�	�"O�}Y���1�-R�� t����c"O:�`�Kȝݺ4�p��4tP��g"O���O�(X�XI�@��E��"O��x�Z}f��pA�ɔ7�F"O`���������D���W�"D���"�1D_�}" ٿs�ܘp!O%D� HP��$W!�50�J�,���($9D�8�̉�|��(T�/SV��%!D����z�\�)�덾�, �d D��+���p3zT������@r�<y0��8�� C�%W�	B7�I�<���7�>H�c�X�FL,�sE-T�<#���+�Z4�hF9�q�8D��(�F�����c�GO��2d7D�����f_�d�2�&C?��r6h)D��ң�$U*.ቤ�W������&D�Xj���^�B��ZR�
�9D��H7h��
�H7��;b��u#*D���b�
aQ��� [č:t(5D�� �LŢa�Nd(�eЬ}\����6D��g��Dyvĉ�����t@;�O6D��pV�Xf�t�Ӡ�L&*�����>D�܈�	2!����f�8^8���0D�jb$މ���1�
�R[�E�$�-D��#���cXƁ�C�̱	�VqSN)D���#�+E.d��BJ�`�2�ء�<D�Li��@�}>Z8�D���<3�?D���E�
p�(�Ӯ�?h\&�W�/D�|*��qM���ޯ2��-D��*���.!��*���'s� P8ƌ%D���� /B�m:"^�"Y���0D��9�A�/?v�����5�Ա��a)D���v��`p�ن��J���L)D���	T��	[�+@6���)D���QːB��=��iݹjx�)�V )D�dy0M�N$�H����r�P��%%D���0 /*!�pX��ˣ��0R#�"D���E�KԮ�(]��XW(!D�\yv���N�zl;u��=��tAf=D�l(ň�	8 ר@����v&?D���dW��bp�d^bT&���?D��� O9!Q�YE��l<D��f�� # � prb-t֑��:D���KB2s��{1�15�k0�$D����(8 J��\��m*W!"D�D��oQ,�Z}����o,��Jө?D�h���W�G����B�f��ZT9D�4ѤɊH��
�� S4\�J��8D�ȸ�킞8��я_�X}��[t*O>�x�E��b$> �W�Ȓ�
���"O�����5N�L��J/�1��"O� �Q�//)��h�ˉ5�m�A"O	��JJ)��8C��:&fx��"O�&����R�fݜS!�Pb"O�$8`b[#���H�E��K��e�"O����͔�lx��(��Ș�ՙ"Ox��r���F=�D�C��m�"O�Ȓ���x��P��"2���SP"O�L�a)S�o0Xi�w��sv�)��"O��[�k_�"�
U-@d���"O�-� �)��q��3?�]p�"O���7�\V|M�L�����"O�hӁ�N�uq B�'n��m!�"O|��0�o���� Q5��L3�"Oĩ��*E�S�乸��R��mc"O��C�>2��X��>�x��"OQ�hä� 8Z�lR�3�vŋ5"Oʠc"�J8"�Bq��ʍ2�8�"O�}zu��?"�^���)F���x�"O8�����
i(ۤZ��ͲT"OX0��ψo#��Z��X"�>�i�"O���C��R��Dif�V/B�FШ�"O����	�*��M�|��U"O�8��/M�3��mJď :D���"O:%�!ا[�9@Ԡ��2���U"O�L
�,̟N�:�a�3�H�)w"O0�ʔ��HS��!�*`@�"O��#PIJ��׀�7 �R"O(�x��Ց�` ���X�=���A�"OF`�6� ح����:ݫ�"OX=p��
�t*B�L�d"OBXS�$I�]0b��œ�d����"O�@�Q@��"%&b
��"O�M��ڑY���c�"��B�"OܐAq����H�0#��(����"O���GOG=N�u��!ذ�-Sb"O�4i���1':E�nچU�|��"OZ�"q+W�~��+��K�JyP"O\,B�	�,p~��ۖA_��+�"Ox`���+��@YK�k~b``"O�œ�!˥6{��A���zw�X��"O& 8��ߧAf%`�K�PsJ X�"Oԁ��c��v��Y�j���1"O�Y���!$��� p�	T��Y3"Ol�8�O��&�^u+%��00 X�U"ObiS�B�X�hШ�͇���xp"O꽢Я�$S��i[�뇣!����"Oe�����QJe�W-ɰ����"OBD�5�H�c�\�"/��,�LX@"O��*ƃZ60����#���*b��"O`�q�-�J�|Ö��'�Mk"O���扄>Y���`2#��x���"O��ÊA�.��mx��=.�5�0"OR��D]�h2���0�^'�@���"O�D��'�73J|IP���0�ld�`"O�-JT��!s8@�J�E�<p(�"O��X�,\5A`d
��H'u�zI�S"O�\�d�Ȏ@���d��&m��"O����D[�#d�@�+H��hV"O$0%�ARD��!W2q�&aڇ"O��ɒC�%P��p(�B\�iZ�uh�"O��W�� "�Pr�09�-�"O�[v�ЭSզ�0� +c.��T"O��r!��#� �y4�ʹ}���6"O:i�/��400`Ȍ;m��urs"O� 8��� �
h�e���K64�^Mt"O"����/{� l���J6�ʐ"O��@uɅ�>�V��&�ɉ9�r�"ON��RG'dN�k�(`�h���.*D����W���Äf577 �!&�=D��H0oT3%:�ȷ)E���TCq�(D����#�"l�8yP��/�]��)D��Rv��].�TZ�LA&���*�"&D���#d�=$�\S�߭cp�$��C(D�(���<10A@�o�#N�XP��8D���6eS� D���["=RH�)D�(�wiD*�h96料 %�E�&*&D���P��V�*Њr!�%P�2A�¬)D��QD"�'t>�9��G�J,�a&D����E�B��S��p ��i%D�@1�-�g�2�[�)ε=�U9�g"D�X���4w�؀"�� s��i�n#D���s&A�e�X)�T���'�����#D��
R��S�@����S�iW�1���-D��a��{/�l�Ј��`�VI�R�/D�,{c�T}���e�U�:��� �-D�[�BR9(2%R�@��X{�K?D� ��Ϛ�6Hȸy��9#�@�a !�/'�T�W�AUv�Ш&d˾�!�׶<�L��IWC9� �C���!򄚌{d���7$BQ��Z}!�΄��)��R
"V��r M_!�ĉB�l)��i �$�O�!���<l�EPr�D%qG�0��mY�c!�dA6x'HXr䄱X1�D!g�ؖ=R!�D��Cbd�" P�r�M�9!�$��]L�f/��O����?�!�dJ���I��V
`�i��*
!򄅣:�[�ȗ�KA
�+ԃ�+!�dI�0k�\��GZ>S#V�+X�=��'�8Hc�!}p-�7�ЬJb|��'9B�� Eѳ-.R��(�Rh^\��'8�$��Y�^:�����G`h 9�'����W�_"�0*�b�=��}:
�'�,�Sǭw*� ̓���Ĩ�'�TMY����C'�A&��ْ�'�>UR@���o���яK�\��'t4x�$MT�Z��,�Q��ٞ<��'����<1��rbΟ{F�i�'������y�%2bF��m��d��'����b��)��x�`��>QKB�y�'@���fU!f
j��F��y�'�t!�!���#-n��@ �=8<��I�'�iS���X���C�ߣ-|$�
�'��'Eʇ#����'�(Q�Q�
�'%d�⣇�N�:��iP*���'\TAWCQe���󪑧i}Ɣ��'�<��S����6���Y6a81�'��j�R�|����`��EMn���'�fLC����n͸�g��3T����'��$X�B:��UCbޫc�����'�J�#Z*�`b#Ԓb�n���'$�-�@�)oG�9BK�_�L���'t\���MnЕSa��S,&,��'�׬ޒe"�ԉ�QK��C�'$t�h��I�(
�Q�CJ�����'�,S �A4I�����$�/=�����'��٢�J%2R&��a��0l�J!��'ǀ�B�ㆇMF4,1&MB:^�Ȥ���� ��s�ȝc��b2j�
'���v"O�y���_k<��TnP��b�h�"O�d�2/'%)�6���N=b"O<y
���t� �&-�H�� "O�LdN4�@��Ѭ �N�4�"O�] `�D�4�$L	��@�L��8�"O�!����7Y�^�GLQ5J��|�2"On�y�l�0nzT�E�Q(G����"O��xf���U脌M=>�lӵ"O�����y�-�'l�$rK�Kv"O�x`N-�XYd�M��е9�"O��q'�N�<Y)W�E<1��ە"O���7"\�7pH-`6KX�=�����"O��i�5}�������rv�Xc"OZѻ��Y�/�"�1!��"?�~��7"OL�A�L�Rũ2� n�	A"Oֈ��#�b�J�;B�x0F\9"O��2�]|�e6�_�Q��;1"O�+��]�Z�er�)	�1%��B�"O�Y���Y ��mCTH��$fx�"O�8��WʂɃV��:�!�5"O ��!��~l�����ê~Q�5z�"O:���F��	[ -5f&`Ę"O���&��|J����&R8k���"O�K��A_��{  �g<UC"O$��O^�0� ��/[mF<i3"O�ZvCA�4�����L
EGDL�6"O8Y�����*0�Q��D/7@,��0"O�ыd-�������;�$�"OT4 Q�H:M<�2�	؈�>Tyw"O����$=~8ʶ�l�u#0"OKCVf�
t��	f�P�r#D�y�$d@�1O�^���"ԑ�y�\� ���8�`�\L@�P*���y")q0�M`��@7�
��V���yBI.:v�H�+tT�F	ǰ�yr�^�b�@��D�z��*�y�'�_8z=sb�|`:@�GX�y��JV+�%��N��{��թG�L�y�^�_�^��A� z���KYs�<��!�[���_q�e��٣m�!򄁫�
�R(Q�`�m��n�!�dU���;����&9ö��9�!�D���� B�B2���ӊ@�]�!��54-(#% _ ��j@�%-!�D�G�$݊�FJU�d$��,!�ݕLЌ�Ch�!��i4�!�d�}�����Z��  �)�S�!�ğ�-ٞ��'K�Z�RmHg��N�!�dX��FaZ�J[�UqDղ���x�!��;aR&E���M&in(9b@2K�!�D�h,�U%�:+ 9rN�;p!�	f( ���eJv �eǇ�#!��)�PXac�l, x)���@&!�D�H�BJJ �M�'$n!��)9�P0�գ���vB
�4�!��_f�=XbCֻ/�X�Z�A@�E!���F[,\zU�/O�XNS�Y�!���b4��W�sh|m�@/ڇ^�!�$@-,��*!`N�}uj��V �%!�$�<�l(HQdM0X�Ƭ���>$!�#9�H3��>g�&H��hƨ�!���1��$�`���/�|(�A!ďA�!�D�5W�z$)ŁU�-@l� ��!�� �P��nר�>L0"ԔM"��"OpiRSB�\˚T��K�2��F"Oj������$!H���/�3=ŌD��"O�4K��SB�̣F-˸g���'"O��hp��?xV�=���V�e�6�[�"O�Sp�]�]��.ɶ9L��"O��9v�Y�j�B�M��.���;&"O���@8�,)��L�5�2�J�"O�(F�R��z=��lJ�x��"O���	�U��	�2� �"O�)*7&ǚ~ߊ���-�T���ؔ"Ot(��T�r$P�'X�/NN�s�"O� �B��>vP�5�̸t@H]�"O��Hp��^{f�I���^,���"O8`�g� C	6�bH���1 �"O� Vk��z�ǌ�U���!1"O��r��[�-�B�*tIJ>
�����"O�諴/�9�*�k���(,�X��"O@%��$�X��M׶C��9v"O�yA�Β��,��eBl��{C"O�Ժ��+����؛ICd�8�"O";�(TaBT����.ruQ�"O�){�IY�o*�A��l��W)u�G"O�XR0]�h���
�8��1"O�M�$�W�C���+E=y��YS"Oa�@�#W����%#0��Ң"O�<˔�E�I�> �ac�<.���a�"O}�#��9>�thc[13�r�pR"O�FjX2��À�d��-#�"O\�(��߈pk
D�Qv`���"O"8�M[� ��I�-�h��"O������(�t��I�^�P��"O8I{dh�xv�)i��Q����"O��q�Ϡ0cZl{E��_h5!�"OrlvFʹe�Z/�|��!C�Oz���]�dq�b��?o�j�@��yR
�8M� ��jӚg �1�O
��y"�M��<p�J����ۓdا�y���1
(/��`��g��ݛ
�'_Ш�Uf[�
����S�FTp
�'���H3K(X6d����@.4� �')��q��7{'��h���"n,Ř�'rި �b^�-�f��`^h���
�'�+��|�K�	�_���:��$D�hQ��[�AU:0Z��lڄ=�R&!D�(��� 9�J2)�w�d�R��4D��R�DZ2�~�#���25�3D�����X-�T�a���	Lf:	ؒo2D��Pa�˥U�����cI�%r```��/D�x�V�]�^��eF�G2_4���+D�|)T+��Du�p�sE¸j	�t��+D���u�]��pD�D���N��Q��c5D��c��P�!"T�*L%om<A�4D�4K@��<=L8Y�(�B��좆.2D��R`�C+5�>�hpB~��@���*D�8�Q��-φ����_���)��(D�tb�
A.P)`f�		�Ѣ�,D��;�Ŕ� �NB��˦U��X0da,D�d"��׋2̼h%lU#_5�����>D����C�_�XYIeiUE^+��<D�H�v�..�� 1�ő""Z��6�-D���v�խD�@�)�J��f�0��ԃ+D��a5l$$+`��LN�����i+D��e���c��7�7j_��Ҧ$%D�� �`0ѡ�/p��!��±54Li f"O��C����i�HC��	\�\�js"O�5�Qi׽�+��/c�5Y�"O�`����
 Q)�∽'�F�	u"O`5*4�R�$�Li�OͤxaE�"O��n��@pDlI����n]�|iw"O��pL�>��H7c��I�hbF"Ox�I��%6��d�:'̀���"OXqX��-$�����;�q�"O�,b��]�Ι�+�6��xQA"ORA��ڝ"khpb�-������"O�u��0U�X�������P��"O`���c�!*G��I�m 
ᰌq�"O
u�g�79(N�
Q����h	*e"OLQX�M��4bf%��z4"O�,��JM/<ޘх��4�x"O��8&'�(�2Hx�4:&d�"O�)�ҩT�U�	��_�z��"O�yj��7��@3�S.b�]!"O^m���έF�F=��I�4����"O����&++
hȓ&�K�,@�D�5"Od(��H��k'��+Hx	BiqA"O�L�'�Rc�X���б{�h�C"O��� n8<G� K%CR�J�E�R"Ob9�P쒌^�8%�h���C�)9D�|���`��tsQ�M�"+4Dy5$7D��s��	\��Y�tK9��G6D��أ��)&�`��{O��5�2D�x	�R0S
�5�f��<x���J�k&D��*�����(�!nS���&D��$$��P�VgŬJ�Y��?D��(4�.Ca�tY0��ܙ�a?D�X�v�)v���0GF�r��� � D�49#�25+������9;����>D�t����7.@� �bM	#U:ȓQ�<D����iP�t}Ji!W�Ռ�>��'-D� ����:R������0;,��*D����KT��|��P<i4(�WN*D����T9�v�#7P+ay��A�)D��	@͔H|n(0#�X�#% YԆ=D�{b'Q�.XI�U�,x"my6':D�,`fG�\����T�h"����+5D��I'@�d�2eR�N�#S��d���0D�py�I$��}���D ����3D�d������r�C�c�ڱZ�$2D����/29��uE=��%�62D�ȫVL�A���I��
GȂ��CB,D��s'��#P� �`6d+7��52�(D�h�vI��6�Cǯ�W�B�9� (D�$�p��B6\�J�hmBx�)D�ha�
Q�T��c�v�^�pb�$D��;��˂s�����hR �D��$D��K`��.�i��{�X%�ר$D��:Q-�g�P�pU�A�>�h�Q�&D��ru!576�LU�2�BL9 �!D�|��"YX��0+Z,h趉>D�ܲgT]v�h��Lh	G)*D�̐s��6d���9a�D�,�S�(D���5K��48Rq+&iE�Q\��
$d(D�Z���H�Nm;�aE9H��d�%D�\	��3l�Pb�A";�5�"D��Z��D�����#L1
F�$D��p��ϻSҍ�%���Wi"D[T#"D�8�T��/|2���f��:��1��4D�� ���we&S��cԣC�L"��"O|�Ia�?�$��e��d2�B"O��g��4pԶ����OF"(��"O�����M�P�(T/	�*
z)��"OP��%��cc�E�ևJ)'2���"OD�+����8��r �̠S�tL+T"O�y&G�*U[V�bc���z�t�9U"O��ȖA��/S�=�""�8e�Zx�"O�=��Gσ� ��$!P�qҮlBg"Ox�!J�7���Ӄ!N�'U��!"O����#:�ؑ@״`:�Qb"O"QZtc�.*#x����V>/���%"O�t;wh�P��P� ���� �d"O|@�7AN��8��F�"O&h#�V!81���@�i�~��"O��zeĊu?0�����֌cD"O�҆a�}� 8 ���r�"O65�#�&xTpұ����"O�"0~�,!�Wk���Acd"O:�X+��!�	Zf�\�l�5�f"O��T� +/�"9rD� =R��|"O"P�g�$6���"����jA�S"O�3��&-V�i�����`��"O�m��H�{�Y�(ēal�Q"O����e�*gsp�tlȗY��!�"O���Q@ԎЬAcW���3��k�"Ohl
q�	+~�
���V_j�L8%"Oj�XJ�Od���<h��9�"O�ĘT ש~ b%p�oJ6�$�Q"O��� ��(Q���X�L�3�"OF8D�^.|��9V�	�eըDp3"O��{��#q
�p0$J�1��e��"O���ă@���Tㄦ����"O��"SE��F_@�����&CK"�"O�Z3��-c��m#6DdAXs"Ot�bb�\@y�)��O8Zn;t"O��Bc�$[�]ʄ�ޖl��4��"O-*�
�L�j�`�){�|A'"O�����_?l������A�^�0�r"OhP2�Fʹ�l�h�#=�x԰"ON�SУڼ;*�R���m%���B"O��P�#� "�T��d#�iR�r�"O�c'��}��%��h�1M��@!"OԂ($�$�ȉ�]��8�!"O��ʴ�)N�)S$Μ5�V��"O� ��D��r�q$�V�V���٠"O
�K�M�c�|��f��o-����"O��@ǀ�O����
֍ "=0"Oj���f�j0���h#o��@"O
�Z�ۇP��e��$��>��"OJ !�d�{ )��m��b)1�"O:�j���&K8^M�D.��z��(d"Orp�H
%��1�r�U�L�x8�"O()�uǛ�"ayD��?�k"O���BD{�Z�+U��\�T!�"O&���!W����F�`���C"O�8�.I6w�t�cMh�����"O`�ᗅR	���f T������"O$�i��$�{�ÑEf8����3�yRޘ1�x�JrT�@� ̉��:�yRIS�WNh�`2�Յ%D����ɘ�y�Y	>�6)�஄�z ��I�5�y�.�)rbl(uj��Df��q֌�y����U�k�~�>����)(��B�)� j�'��YZhP�-6��'"Oԙ���D�#�v�)C%L%H�� �%"O�b5KX�^1ޤ�gC�.8��ݰ�"O^����V�"��{��Kj4��c"O����Q�=��JY`Ld1G"O���q��7KX&��1
15�S"OLX�$À1�4�{�(��4�eQU"O	i'�H�fG6���<�X��"O����͐�@�)Q�O���J@7"OF-QC��@v��fIT�\I�"O�@���iN�q��*��$��p�"O=��y:�bI��	�4ţ"Oę��k�n^�t��(�m��T"�"O�a�CdD?&�*<�A�B�W۰-�"O��bv#�0u�����H��k� p�"Ov !��%^�Б�E� �#�`�� "O�	ˡ��<.6@��h���t��"Oq!�6^�> ���Η9� �cG"O����nl�T���\*��q"Op-a�,6�|����'\"�2"O�`8�!֦ j�T`")\�~�\�kr"O(x�T�ܕh4�rW͋ *�"O�}��E��%�`�R�Ǉr���@P"O�e��)�pd(5̀$1��1H�"OIcQ��T�PՂR쟈L�fL��"O0}�5����aa��L�xq�|� "O�� �� wX�Tk��Ή:�pi2�"O|��A(��<�u���PE B�!��X�&�����U�v�L@��ȼB�!�Vv��1���+\̸ 2��0j�!�dU�	60E���ihyh&��:�!��?u"��k�nV�pv��p#��gr!�$ײ)�l�T��o&���%Ӂn!�ޑI�0��R 
�T������5b!��5Q��!���ܔST�YV�!�������\0u�mӀ�]�!�4m��D�Y��B�ѝ�!���$�|JA�Z>yᶙi�����'q ��E�&_���VAB�f"Փ�'p�h�$jæ#rܬ��B�
����'��a����Q�s%�.�*�;�'����m�&h������n �'�f��@G	�cuf��򏖞�- �'�\0V��'6Y��I1�5���Z�'�N�[���[�i�5 X�'j�I
�'�|�1󆙽w�p��h��78��	�'���(R,	�pH@��K[d�`5�	�'|`�A�`ϧC�Np�Ј\��U�
�'{��0�F��6@rHJ7 �`�1�'Q��	�6=��*5뎻%�i�
�'��L ��Y^�m�*�:����'����#C]��E��,A�~j�� �'��I��d�q�p���K�Kf��'o�@�7A�VP\|:��KCV�!�'ӊ]+ug9,( c��G��I�'|���!���D�e��m�*L�*`�'�i	��Ĉ��1
�hӭ?�̬��'����@��"]�S���'�(d�� �8�x��� :(�i�	�'< ��5'
�.s� �����l�",��'���w)�)|��Q�X�k�|���'6VH&e��+$���j�XPS�'T�ቂ�Ĳ9�p�2���zc~5Z
�'��`3LF���'-�)֨��y
� ؅y� S4$�pQ$�O.:���8"O�ӧG�Ak�|�2N�YB$�4"O�1M�W�i����2@z��"OrÔH�Fbe���l,��c%"Oy���(�\p�i�Kt~�4"O�2֦ðc�:� ���~\��9�"Ox��*�8uf.���aB=y2RS�"O��r��!d7���bA�%@�r���"O���Fb���"�@Q*H7� ��"O���kܣ`�t���G��A8�ԋ�"OLU��
��#�����
�,��+�"O�{@����a(v卷[�8)�"O�|(��$��xbuN�+1�L ��"O�c0�ө"�܁I2N̜9ŒHpf"Odi�
ɑE��ĲX2"�V ���y��ǥ2A�����2+P�,�����y��A�����I0a�+�yR��{K8-Jsd�����M�:�y"�R�Z&����Omb�ɢ�y�!�n�&p9&��{Z��5�N�y2C�L�`D��&���NQ�y+��3��;��ȽG�`2�e[��y�'�2.�0�T�5<r���gh)�y��P�H�j��C܆:���DF�+�y���"h�H%��M�,6ϔl�6e���y�Eҽ��� d��'�b���ϱ�y�@Ԋ���%�-(f�Y4�	�y"Η�eatP�w٨{�*�m����t��;R%a�LB�P�0ͅȓOIi)6#���z���ۼ!��K*tL�P��74���3�!�;AV���j���{��L�$���莺Ke�Ćȓ/�j��O*bߔ RY�
d�ȓ9{~����\�'��偀aԳ;fN �ȓ6�X��ц�>Z�Hb'�ò3~P�ȓc0m� }�)r�Юp����P���04^���ɨ
F���;#�AӃ�?Q�\%P��Z����ȓ{3�T�AN�/� �Cqa�'V�b��ȓY r$�a��>��ya+	�Fo�|��[�������PT����R�/�vD�ȓ%5zQi&'V!95n�x�m� |��ɇ�U���q�����i@4�Ǳo����#)�u�sB��Nl�a�EA	p�d ��CՎz�!Y�06�(	��ǅ3�HІȓ:]��P �dͬL0�jԁ44l5�ȓ ت9�g ���Q�D?�h���C�ތ(Ī���T�%�	KH�����G@U&�$:�O13<5�ȓ���qC@���l��͐����{L(�P$�$�����D���t��z�e� bQ=�\)@�	J�Նȓ?�X�k�g�zaz#B�5t4!��;���W�U08gZ�^�A}��������<.Z0*�oʼ+ڬ��.
�9*�"U���s�]����ȓ&<���c1Y����6ʱ)���ȓ>O�|���M!%��;'%@'=�tՇȓ{W�eJ�.�8^�ǁX'Fm�t�ȓ38�QقK�>� q�� hB]�ȓWvx|��"��Dcg#�_�"1���6�(rC�v�ZhF͆q�d���V���bX�zz�]9�/��+�>h�ȓm�6����L3&]B!I�!�>��Q��S�? �1Qpf]:T���u�^�>���"O|�)��R����PBR�;�j���"OЩ����O��P�U�Am�腺�"O��R*J*
�6`ш
4���Y"O�C��K�(*ȝ��,�:�^��R"O��FL�|@.��!K�A�41�"O�����aBV�����A�U3"O�E!������3��P#	A Yj�"Ox��C�Z x�jt	�G�OM,�yg"OR�s�"��4�:���,94����"OD	فC��FZ�a�I	�;'¨��"O�̓��G�0�����=3P�x�"O %��aU
g~hi �A.�ͳ""O����	M�x����dՎ$̢x�F"O���b�+2��(ڴ�;���"O�JC%L�"�(	d�X�"OD���nQ�0f��X�ȊP��mB "O��8$��a#��1B-C�\�@"Oq�q�J٤�
`�D�
��7"O�tB�O�~�$b�"�.�Q�"O��d^�
�.xAB�\	+a*���"Op(X7
V =�ޠ����!xv<���"O��§���YՌP���܈.7�<*�"O	�!e��ݲ��@6i	6MBt"O ]�'��7��xS�` 3-$1!�"O���D�G�P؁sȍ��m�f"O��r�/e��0�C�!.��`�"O�����+�5S6�3t>�"O�ł�O(L��G*?p����"O.���*^���v�7?�t�"O�	SV)�#�T]���((��]B�"O� @�"�Y���B��Q00Z���"O��[Re��|u�K��O�.��dA�"O� ���]�}�x�iEE�S��T��"O��ף� �m!��
�lM�U"O�up�ζ{�c��4���yg"O�4%lJ�QDΉJf�ѻ��4�$"O����[�����C	�v���"Oz�A�'T<�v�pb�Ǭ[��ф"O��5i�:j��$[D�� q�m:�"Ohu�d,?}���#Ϯ@m|]C�"O�U���@�J�}���$%frP!u"O���&/EC$ ��D\�(T�Ey"On�/önl>u���ǼfJ�!B"O&D&	^�8��C@7]9�AG"O�g�Q+�B=��A��0+� H6"O,1Iϊ�MN�p��!	Hxa�"OpM@��1d>=A$��r9�"Ot"�+��	fMr��X�X�,�"OL��A�|�R%��LDn��"O )`f]�1;B�@l �9
�"O2p0� g�p=k!ő�A��x��"O����_y�Xa8��L (2D���"O�t��l	�h�x=��6,�m�C*O�ɳGg�xp�1Q��p���'���A��9a��D�aS�R،a�'���#z���Ɉ�bHX�
�'ꜹ�pKA7�V�j��U�F�*
�'�����	�P��,�>��$	�'¼MZ�(� d�XJ��4)�'�: S'��K�"Ȱ�%V8>�v!i�'M6@CC��Z�����![$n���+�'����UC�/{I�v�Ӎ84y1�'L�)���A�D�j�K`^g/ ���� �a���b̥�"�[�B�̉�5"Op�%�-��p�3Ŕ�{���"O���`��0c�|YU	�]��U"O��0$�1#H� *Ȧ �$4 �"O�8�"��f���`�Ɗ�1X��k!"O
9�G��,v`5�eFɞW]D���"OHhq`	/d(��h�M�SbĨa"O���DkZ�8s@��A��U*��"OV|r�d���$���� Dr5�"O��(�Ś�v p��4GAn%�!"Of�d(Y̪ݒ��R�	��[1"O6���MB�R��Q��?��A�"Of����c�֠�VDZ�q���Ar"O��`#K����hD�iy֙�A"OlA�Q�E({6ᙖ��y^��!�"O��;��8kB��eh!S�V1l_!�N(, \�q�Z9wD��h1�Ρ9�!�T�jE�t"� ѥ)*��Ph�� �!�D\8l�f�;0�ˌp0v1���,&�!��ܸ��h�QnG}�*��3�ϵw�!��0r*`N1>~��ϙ p!��D�*�����	6.�F}뢥�5D!�DG�T�4p�
@��!t�!򄃁hF�XU�-~b�� ޭ3�!�Ssvq��7q�s �J-�!�Ĉ7��{3��%Z8�h�NL��!�R�^lu�L�Q��%Y�m��w!��)��1��6׬�#d�Iq!�-Hot]8��@�.~$�i��Z]!��]�fv���ё[8;Tǟ 3!��H�5�d]�5h|]���˟!�DЪT���BE��/:i�ͩ П*�!��ąXw���܁gb�<�be�@�!��P���ق�.ݧsUD����N�!�$-�r�i�@P=+8��y�D]�m�!��6N����ĩĿ[:Px�bćF�!��V�6XIB킢*�4/U�!��I)&u�4�Ȉ�y f<a��Am!�$ע�(E!Wΐ�}��ԍۇ l!�8X��
�F�5~�a!�.��!���S&�=��;C�
�%LK2{�!�X�b4�y��G�^�$mzъE-�!�d�ET��@FA�;�@X��Q!�䙭|� Y�+V�@��Yd�YV!�
�Z�h0V�G)��x3c��'f�!��Ҷ%+�e��t݄�Æ��L!�D�p��h��`���I��	>!��#Q߸��c)"��k5ʕv!�Y.�h��j�a
I`A�h�!�Ę P�zL	v
�MXHY��F�( �!�8lTTU��o�0O^�g��JC!�DXfT �CPN�k�oԧ&B!�$�O����,Ũ����2��J#!��;Ɣ$C��P��!�ܪB/!��8�f#��72�lq��ŁI!�ъ������(8�ȕ!���dT�,CD��<T�h-�g�-!��Y)Bʄ�Ȕ�L��\Թ'ݶbx!�� �!��p㏒�i�HP�d��}�!�� 25I�(R�ЍDo� ��X1�!��D1V��z爟�sl`�Ȣ�%�!�D�d��c�D�8a��R#��$�!�ė*'��x� O>e؁GO�&5!�W,0��
���5WL�I�hU[N!�� إ�D8G�h���cR>_@�U"O�h�.���#�̾k�x��"O�,�Y3 Y��֝F�fĀ�"Ol`[1��N�4{S� %C�P�Hg"O>ha�Gŗi�� 4��< ��6"O*�r��K�{	p���M��~��p��'XXX$��S�M�TɏC����'I,`Y�`P�f��AŅB�$�':�H��cF&�b4�C,>6V�\�	�'p����ء2������ߞSL��'u��p 'J��<QBk�/y
N�
�'�D�Ć��*��A�]�G��-Z�'���E0Q�P�+�	�:�Z�q�'��!p�	!�"{�iI�6�@T��'�J���˖ j?��0�.�����	�'�B)��GY�x����mԶ[$��	�'!H!��a�<�R����ȃ�~@��'�f�����g�b�J� ރ}@,H�'�"�c��V�
\���.s[T�'�����L�Nؘ㙛r�Bt��'+vY˧�ߍj���BĨ[8o�(P��'�؜������A���)y�z%�'��)��߮��	�#�n��A��'�buӐ�I["L�bG��Z���' ���%�#S�p�'���:"��'����KB�q��!�Gʅ�;�y��'Cn��1����"�(GG�~
&<A
�'�^qK�m��F!tj�
,k�<j�'͐����W�T���� �0�2�'~z��
#g�)8�@�8z��'oj�)q(e����(Q�B9!�'�"���N�Q�a��& ����' �7(�)�9�4L�b���'Y�\; j���PbʱA�:��'r���0�� A2]���f�x!�'�H��.�
��t#���O+�uH�'���(�؉n r]¬��D�X|��'>ش�ɜ�ΐ��ĥ��	����'�a2bn�?f� A1�-/� q)�'��,2�P�ev��cA�!�
�'9Q�� Je���C�{T��k�'�@4����37��؀g��qL�Ѣ�'��1�� ȃ���NF3�p))�')x�0��ڔd`��&fT0/�m��'f�h�d�0j⾀�" ,*0L(��'1tmhUfX >\���NYg��
�'��hv� k4T�� َS�V���'`�|�vD�O0�l��N[:8Yȩ��'J���͞�&F�L�����CL�$�	�'���)% ��J�`����>߀���'�0�s�A�'zU�P�%��/�DM��'��T
���4+���.J(��'K�LA2��DgD��S���+����'�ɐ5�Dt���C�V��D��'~����+�$q1�L�"�� z�'�x1T�  :*�E��$:	�'
�I�T�L>�0	P����6�Y �'�(�3+��J>�\7�M�s��ʓo�%x%E֝6g�;UK�-lN���)��`��N�$w0x+��Ƨj�R�ȓ䢑C"�#.�l9�n@<"ԆȓKP��u��>J��B���P
�k�<�`
 �9"4AU�,eƜ$A�D�d�<)&�+`I"Q ^�Df0��S�UY�<� 4!!ϖy/� zOK� )�1"O�҇q��P�4!�9P�!y�"O�I�e��=h��a��D&3,tr�"OV�!7*JW��@�@O�7J.��Ӆ"O^y�ѦR�z�@Z!�WM\���"Ox�4c�w>y
"��TK�Ā�"O�ay�L�#g���p��/DF��"O̴qc�9<��q���7l���D"O��[$NĐP����$�$2���g"Of���>��ƢĚId��"O^�0=
�B�� ٸ*@U`�"O`����R��x�CW��2R�A� "OR����sL����N%?��}�"O���� ���n��E��A@"O褉FĜ�W�Z�p�\!�0P�"O�p���q?���5��V�:eI�"O*I�AF�0'����M�(����"O� �7.H8{����@MC��:-��"O�uȓóg��ۡ���6顳"OiS�H	4]�cDo�\��D� "O���LZ�2֊��t�H�^�ĉ2�"O!���=�dq����-.����"O�%��
�Z�~�S�B��ܨK"O���d�W�|�Sg]�jC~=B"Oкuk�)�p;�lٹ_��<��"OT�	�ȉ�i�d��	�qt��Ks"O���*�n�d�S���tz��A"O��HG���m�>��u�R�h�h�rF"O�gMS2��d2!��4�f��C"O�E80��.R�e� ���Q"O�� bD!!ֈ�r�Mڅ�819�"O:\���I�L��CG5v�f��'"O*$�U/N'���g��f���S�9O�c�,���OF����(��w_)D_J�R�'�@ku)	U3�2DA� =��`2�'��M��m�`!�C�Q*1��L�'���Ҧږ��@��k�t\R����y2��?�Q2��u�P5��C����'�ў�'�~b�<q%����T�k��e�P�y'ŕ|Xx�A�\�i��(+PJ���y�C�'d���\9�*|p3'�2N��C�	0y����wEJ6s��`�L� "���3}�˓��<��ޞ ���BŠc�@�2"l _<y�����J���4£��65�b���#b��O�ӧ��:䀃)ǩ.�H1�v�݀0e1G�I�[Q?eP�e��`��1�a��Xv:rEH>D�l�FV�n1�p�Ň��u?�y˳�<?����{a��K�~ D����H�eq�B�	�t)�y"D�A���i�5�HW�����'$��x��	*p���J���x���oFTB����8�%Nq�̑$)46+"H3�!#D�t�c�)'��y���"�/E�	������S�:Z��@!�
=%�.�a�e�=g �#<�ϓ PPBgNA#(r�@�E����Q�'.�Ex"���U��zҎ�;]6
Y�c	��n�"��T�9D��ʔ)ud�ae�m7<9Id#D�����#(��u��!ѝ����.�O��I7�`�����Eh �B��g^�B�	5Q���*G�Le�DЂC�2
9�B�	�9����·�,:$�� ��Z�B�	2%����cOD��RlK !O�`��%}2(��SC��r��ԉ9�jx3���ybbK:C�ؠc1̾/���L��y�H�t{��3r��&L.���aŁ4�y
� �1��	K|��6��2 ~K�"O��G�U�89k�%�,J�be�0"O0 {�%ּ1�bԢR��1(f��Zq"O�1c�
@� @��CY�OOHT���xb�c����O�xa�V�(_��L@�r��ٴ�?����4($����z�K����$��oZ@�OrY8O<��`�=XI��
�AG��uPqH~�<)� �2�p��̍S�$aXN��r|�v�|��)�c��
ec�M�2HK� ��� ��x�<)3dI#��Ѥ��44J-�'Pe}��d8O�l�@�:}�p����I�j�r�d��a��$��2��4e��c,��i�p��>D�Hh��	�
+�Q8���yT�L���v/ܐS�'���?�S�s�h��/Wg|�1�@[`^n��P-$�LʅKڏ.�.�z�L�_߀�9�蘜�y�kv��E�L�jWZ<I��ؔ�y��D�gX$��┵���r���yb@3?>��a���(���,����'y��l�O)P����C���5��.''�,�'���8��02+&a[�BKά���'�Z���Exh��bŬ��`�j�'��`�#�ـ/.�`�F�M�9HJ`���MIyB�'�4�zf_>�l�!Q����	�'��|V�M��`� �b@�N$��'�. �ݝQa`�K��Ȩ�'��n���4A���A�fy�g���yb@�+`[>�.��H!��۔B��a��'���:�j�k4F��q�N�Az��r�'�6dy$E^B��D�#O�<}����'S�� ��� !0�3#T�3���'�P�k ,�^ �I2���';J��{��'j5[W@���kr��/1��a��'J�Z#�ɒK�܂�n�$NQ�'���H ����4��!��&v�LB�'����S J.I�dѨ�Ԣ"����$ڡTF��rwKD�'�n��r#ǹR�!�D��}�l���Ά�.9#$� %}!�U���Q��ܾm�$�����(?!��$m
���뉾EZ
��F@@%A	a{^��K��'h���6f@'a�x٫�*�+.�X��'LMi��6TꌂB�N:)5P���'�r@Z���	KG|�`.Z*�\(�}t�˓T'jT*qkW�>���ˁ@�%��	������?n��!3� ��|mEx��O�7�<�'-�����Z6HE��э�6ct�!�ȓ%~�{�� a
�
�O�t�H`��������G?i᧍?$'�z�=gU\�s"����لȓ2�̳Bo�;�b���$�*	�4�ȓL�Z���jK23TC�,�s<ԅȓ]Mf	����(=�Rl��A߸�6%�ȓ �z4���< ��3`	>�M�<�����N�k�\�*����q�`��!!��&.$���*d���:��!hd�O���$$Q�B�(Ӣ�~��(��M��<[!��V��h�ƯF�Fz*u�#M�!]!���-�� ;�������#�!�L40�a��/Z��-�OH�����'��|Rh�:��G�K�Z ���ǌ4�y��	�*-��!dȁ$��y��Z-[4�����z����1O[2�y�΂EO�hq�Ԝ"�8��������Ov��D�(�E`î=<&�<����^�!��	u�:|RD�Ex�0IB��!�Ĕ32��5��B �A$�a�3���aΛ&W��O����Ӽ� ���c�U���V@���J�"O��QM_1M7^��"��a��iQE"O��r��i'� �H�/!m��ۣ"O�)��h-RB�������$y��d��	`?L=�`�5
e`�	F46�X��DJ���6�>�[S�£ ϖqȑ-EKVC�	d�Q�W-�3D^񩡪ջA�R#<5�?�S���?9 �xэ[+Pܰ�D��$��Op����	��]>D���ؚ]�t�;��;'�!�R�8a�� ��'��m� ��������oQy���i�̠S��1���]�S�ԙ��'��j��<�Z�B�E'��K�{��'�U�ܐ����3ŉ@m&���'�FHR�A�<���S뛨2�Z�ɓ�O�c��H��ɋ?�t���brܐr`X�>w�xR�	24E6�����W��⧀܀[g�C�I�Xs"���A2� K��̥8l�O.�=�}��b��b3dȁ��Q�
���g�<Y��M�+j�ib 	��nEZTb+�k�<yEšs̲���E��k/����Hr�<�I�c��t@U��A�m�'$l?Q���M�'A��f��ĎĲS����ȓ'n�0�aaӾ/ʞ��S��/�B�I�!�f0H�A��m*�Y�9��B�I�Z�&H�TG]>q-�ҍU�C��+G:�j�HP�$���E/��o��B��<u(�ah�:C'���(�0J�B�Ɋ4g �Q��b��ٕ�u��C�8k��p�F��m�������B�
 �9��F�Rʮ��E���.�rB�'[m0y��B0z��12�� �lB�	X}X�3�Ϙ&(����7휃YU,B�ɗ2�2�`�L>l�TL��<c�C�F�bd6�=PP l��?F�C�I�M�q!R����%�gD�D�~B�I�8
$�'A�%m���ID��SJB�Iz��}��bղ;ҚIs�G�	4�C�I�ARxIy�JT�7QN��V���B�	>g�d2�'�F�.�۴��&�PB�	�I�LD�U%e�tHbѝE.�B�ɐ"J� ��A&*�����9[U�C��9U�`����]%O"Y��� S��C䉬�T���\0q�VHAeC3�jC�	,|���8�Ɍ:=b��p�_%�B�ɰ-�l�uSY%8�����6� B�	�]�0����.�4<�����o�:C�I�1u�̑���[ �!#$.bC��.vT�����%��i2�Eоk�B�I$](���#ڲ|����8ӤC�	��z�9�`��g&x���c�-@�C�	 j4�Sp�
�d����dB�	�t ���a��+m�6�3'�ۓ�NB�.&��sL�72�I��._�/�tC�ɝv<�0����2p.`9$菍7��C�	-F|	aJ�\�����J�H�vC䉥D� �Sv��U��p�2BJ&Q2C�!z�J�����&EE���&ӯ`��B�4uo���Qj@8Rp@(��mE.1 C�H����FV9��ჿD��B�ɞy�Ҡ�V�:;"�c��E�B�IE��1�O(��9- �=Ҩ(D����SeR����˺=��5�Ђ;D�t��Ϧ9�4�g�2j'��h�O$D�����*Q¶y��a�7 o���Ť4D�� ��y�
Y�-�
�s��L?#��iP�'�9�4-�R(d�fʴAn�M��e�;K����'Řl3��^�Hb��2�C5��k�'C�P���P<N�
��`-^$%�����'zM�êש�Z9HJ�=���'�N���%�=0s8Õ�QC��h
�'�����Hۢf�lE�Z�W  0�'p����E��#T���\���'*��h^2_XX3*1\���'g4�u��ʜ�*���J���'i�x{��J�x�qHƩ>���'I��z��Zj��C.��>-���'ji�f 5U Je�p|��#D�e�<!��ك-� �1������,�b�<�W�"[�Pm��O'S����D(Y�<��-Rsx0!��G/E�-�Ń�m�<	D�)�z�ck���d!�̛Q�<IdeB�_[��>�J��R�<q4i�O����"��x�� �S�<!��+b��S@��y�i��]s�<9J�gD�p�F�w`�9��j�<�-�=�B�z1"	���H��k�<)S��������d�S��t�lŃ2���)1��Oy�E���PF��;&�fxB���>[>�(3��T�x*���Q�j#B�b������S�b�� E*6"�8(�.n�2&��?�z"QK�'MеAЏy���䈋�c4��ۓ3�a���}���c5BU�����p(� |&��J�ܳ+�V���虘���G,|O����'\_(�$�H�!���[S��T^�Ƶ��̟�a>��� ٤sBD�ul����ݽ<y�e:�H=e�ƝXU��'�C�I�_~9�����U����n4��eǐ1O����a�]�2n����R=\x5�L~�&�s��R�A�% ����F*�z�R�3D�t� bB=R�����o�v-��aN%,8,ѳ�Č#h��6-ף:�p�`9F��!��T���+6E���ĉ`az�kۣy} "$��4��GEV#0��x*4�Ɖ�
��bӳ3QhJ��$Gy~�����[���cd#�$䄌��'O6&xL�Y�,�ɶ'}B�	$�ͽ@=�)y.�	[q�HRg�@���{D#�=՜ɒ�A�oFl��GLύ!��B�G��pJ��
�2\�ī�1��� 4��$bg����@B���`sI�B��dR��~��Ӽ���u�T�Q ��J�<	r!Z
H�5�]#�mm�$��� �*���ABОJ��B��L���o<��?4u �`Z[��R��9]@��L�q�[Ug]�+)>��qH���=yC�K�!���s��E� �1���1o� [2�޽�p=A�iP!7Sn�:��I�+­��g�D�)ʵ�r'	A�5JceF�!(��ab](-u�\`�IP!2f�)3G�t�Xq�\�����t~�t˰
#s*��BP�˶&�΀'�K�
�4-��Q�p+bM�;py�dӐZ>Q���	�1��(uŶ1c Āf�p���]�d�!�d�{s��`��_�nts@��f��]�7'����ԪEH�7�M��,�)�����A��~R�ڥd��A�Gg�wD  �.�'��ǀy�zbJ  9Z�Q`��sYn�y� @!f� ��� �Lq�t��V����0�C��~BK��ݰ`�G1^qO�i���9T���gA\�Y�Q��D�/~��x� N!|ĸ��>
�Lx�R�����ʓ�8�n��֫��7�s1�N0:�>��SO�?o�1�0�	��0=�ŊG���YU�Ď,Y�Վ�&Z�vX���X�TT��@-w�:�j-������ˀ��Y�DՏ	s�L����i��ف� ���'��y���΢+@F��pFB,�^�@۴>��q$��	4�@(�e�)b��`�_EP���,�)�K%(��?�~]�dCA�;(�{��W�L4ܨ�2O(i��I�NW�xce腂O;��H�ӄ������T�\���>�n�th�5���$ja�X�b]ꩆ��N��fiF�Qhe���L�7��Q�LԪm�p s5�ׄo,�		ϓ%D�I�����l6��pH�q$H��ɶ��Eh���
>��,Z�Wrؗ%FP%��0���H��o� ���@�'��ԩ��¢R)�$)�cMg2�y��o&$��O��o&82�bɒs>�x�@f ����6a����­'��I0+N7��x�m�
\�\�s4��R`l;�ba0��U�ĺCh|�u`��2��fC_�\�c$�6ja���~���N: �4m[�(�Z�AD'~���h� hؔHQ�*����D�8L���Q�H7F@%h5eL�p�:��$��c8�x9���TQ�8(�i8Nŀ����W�S�? ��Cb�/Q�\��##ݿ@�2���Y��c����v�����&|���']zn�ӷ($60��'�D ��@��(�H0�qF�=UQ�q�Ⴂm	��
ĳ��OVMT��
���(.�� X�5�ՏyLBS�I̍0���iٴK�B�������Ŭ
�r����}:��6Ip��iUL�l�X]��Ꙩy��#>�i71��P�M�+�~"n�7Jw��Sb_�E.�tEe@��'��7*�m24�&RV�� q��.y~�
S�&@'�l2u%�B��R�/4-�Y2��7h� �[0�̓4�\UC���O�p����9��$a��յ�?9��϶k�2���M�1�LIk�����#�33�Ւe-��4���%�M'G
�c�nQ�^�jhh3i� Zg�T" ��0�����FܓS� �3`&q��G	��h�� :�V�ÆSXy�����U��.�0a$M���(�j	*Yw��Й��Df�>d�dĈ=S��d�t�ȜmvV6h�NA��#����?4\0}{�'��I��?c`4�F(�nj:{�.�2��� ��k����ƆC1�	I�o;gx�ȟ�mm0$;����&;�|��BC/[i�uDz��Ëq��x3�JF��r�a׬6�4�h��ɇ~@}�$�* � ����=o�e(ٴM9�08E�؁gV���'�<!�����QG�PE�/y�(���bN������͚J�6�sK�Pj$enZ�T�N�	㉓%|%t���
�H=.�UK�V2�W(��\Ҕcr���V�z
����/j
�RqeT�Bh�r!���_Y�9�搬PV���W*u�����9<(��|�TjL�l�*���"�?6&��0O�.�Č��R({+*����Bk�D&�6H�@�+��\�d�B���\�а��H�kTܨY��'(lh�5��y��">�G-J1!�I��eU��RD1~�b�8��T�90MP,@+j	���A����4=��U��,a����h[#���`'o��dSu��n�����Z$"=)� 6DF���ŧ��]��, M{$��>$(��W�rsՂ�k��J�20��3`�B��,H�T8�Ԯ� 64�`�V�vtŚ���"I� �A��Ej�X�p��KW��3� 零͕)�Ԋ©�t~r�C�!���`�RAO,+��0@��'­�h�X TB_�)�Q*�,v��N�B!���A]���R�aހ��H0$B^ �)b�:��YQ��'&$��!a\h�3@/8uC���M��=q�&�9��aq��5 8�Hْ&n^\l^�,��wK��p�LT���װ(H��� H���xB��?]�.�b�
����Pĝ��ı	�&%B��J	*P�����]pZ<�`kS 0���r�J�\	G�E��<*C�ˋ/]�1�@������Ҷ��8w�a�C��4G���`��V���n�#nt&h#����%�.����b�@b��� ��"�h�9>�\�k��M�oT�BGuzWZ	$�l	��N�;��ĉ<L\�*��9x��pM�a�DP'Q:b�1�CD�?s�D�$��U���0�����c-�i�ϓ|���y�MZ,8�Q0l�
��ɞf؎�����e'-�����O~]iE镭S�5��n�`��`�u2O\�"���i�ddP��[,fq9��,Q�=����c��L����P�$�eJb9x�c^�i��t��D�Re���d΂1K��Q��A�=D�i��5y%�P�_�!�D�ش>+�0��Ğ h��dЁix�����3h�F�� ��XK�`�{�^��i��Z����%!���(�b�_�9�V�}F| 2���,�Yzх�n��9�$�q(d� �'W���o�Et4�'��V�� ``i �(������r��3+�D��� �(�l�+v�)N�`5�wb����DhC�^a`�����z/v�R�AM��Վ��ңW�r�qɆ+a�V�p�үs6�'���'���]�fHR�
�{$ �0�,�r u���ǧC��m2�I�]Xx١%�l?uiգN'��C�I�<�80"!�+,,Yb��йa����C��3!������'C��[�O�9�,KR���-
.�'�y�jN��h`C폵F��̉��y��M<(�QWI
4/��x��[;3���"!^�u��l�M�+ڨ�k�O����e��Gl,U�.O�E������Psf�jWF���'VB��G%�%(�t��jߙp��U�E�L<,Y�,[CDK�N��I�
�_I���e��7G�@E~�njs��G�v-ΘA�-˪��v,ʐQ�֪ �n����H�u�KQ8o؀�V���p��p��G�;���4�G�9������y���#�'YNY����<G���9�D�.D;���J@�U�litOY�QK��
#ˬL��KC���aE�@3���j�|Z6єJ(�H	A�ЈX0H$��҇+��$�b��+$B:!KFI��R
d~�I�(��L�RaE	R|�aV!�Q�xȃ���Q�x�XEG�4ez�A�F>N�BEI���Ww����yo�@�FnC�en��Prl/���D�i�<b�f��'�@���'k"L3�A�6Gl )"׏k���c�-XU���Fg�<�(Ѻ��ɫ2�\������hy�	�#,S.=�j�nE/ݨO ãe�hB��ؗ�R�
��)�ë�r?	B,E�m��aЧ͑^���򫍷&�@ԣ&	�y�թ�؝+1��t�֜4u�ԍ�|ޅ�cQOrj�Y�'��O�4����"�VP�wh��]?px%�Ǝ_�F�2�[���gq��K�gV�i��u9�K¾B�h(F�=yr=Ѧ._�D�:�s�-G;;�YG��B`o�f4�E"5�,�g������%�V�ק���?	p&��I@���G�.�{2F�O�8�a�EZ�D|�oҼ%a�X�4lR� S�}(0�� ��	�5p�M*f)+�4 8����V!��P'L�+*0Ȑ����M�犄����e�V�h�s�4�R�d2���3��z��ȹ�T�u5~@{��I�`�L��cR�b��H1G�7A'�pñ&I|62hvN�q2nd+��i�b�� W��
n �٘ԪřY��d��E��s���-@��X� #k���p��.��@�1i�1�@�� �K��X��B�H_�Dy����b뚨	�#��*��4��N��,�^���	Z�'L�ˑ���YC�hS���L}4�)�\�cl�6�v)�$�&wt��(25̾]+P�V�Iu"�aR��\�;#���fic�BJ�[4m �EPC9��@�k�v�'�pySab�W"EhD��B8��n�/n$Hx���c�%9u�
�	��Yi7��?�����&�Q��0���p�����ڼm�Q�jK��EAw�پ�����^�f��ixTk��]�DȒ�^Ǧ�ۖl�9	�~�a'K^�[�d�o��zܔ�SA.7�b�S�+[|���M�j�Hb�n�
?�yF�3kΔ� 'b䀸p�Оa��%Q�ͫk�Dz�I�8�O�05��..�K�
h��RօQR�8y�BA�*V�b��V�Q-bP
�P��*"�"ekGm��J��P�V�� �� ��4�%�ժ���ຂ��d G1Z����	)?�N�xR�kJ�`�0tK K�p��A��,OwZ`�%ɹ��][�n ��$�DJS��s`kY6u��9!�P�Iz\p��	��[�M��R̃�e�<J��UGg��@�a�'�H���^�,��]:eZ�8^ qXFʁXY��r��1�^EUָ6\b`a%�/cy(qs��Q�z�s%�0^��b'R3�NeH��V�4^d�]s�9kC��Д�C��ڨ�����*�,����ު�L��N/;̖���K��kM�z�O�5c*	�E.�qB�a���j[7dWs���14%`��G�qKf�yϟ> 0�S���4"?n���'1ڥӗ�6b"�ar�W�5,�m*@ݻy3I�&�� :d�2�✧�u�n�G�~��T��X������K�go&Ѓa��|Ϭ�*� M�.�$)F��?�)���*?A���ˆ=�V��'�F�J�04��*�Ҡ�#n/u�}1���FYH��Pm��?�Z�J �[@�T�X�U��Ԩ���.3��5�f��%[b�EF͔��E�Y8��4�L7˾��t+RnkJ;����;c)2q��4�����4u�����P2mH��)�H ����=o!e�6�ޔ*��1G25�(�=a��iYq�x�'x��ɻbB�W��,J&ȁ$`p	觌�,)�i��|�z]z�+#���QqJ�R��}��薧�x!r��[�������|�	�BU0a�iA�<����$��Pl��B�� p����ώN;��hU�.�ħ4�n�ۡ�w����7L�36f����>N��5I~�F;��A�tR��$�'��q-5(���	�^���bA��S�����A��_!���uO	.>ldS�*�(|>���(X���Z1c�4P���ڷ���<�<8�".Ӯo��r"�"�ayB%�^���;%J�<A>,�i�֨�]X�!2f�H�9z楒�\1�<�@A	6&�#q�)�i8a�O`�$?��5��=k��!
�hT9M��XGF:�Q�p�T���|����7�W�@K�z�T ��X�7���,J����@"b	�3b��_� ��*�t' ��0���k��L�xh�f�5R�B�J�vy1զ��bf|%�1���o�W`�](�����S�.�֨��E��(A��+Q�P�n�B���Jo�� �~�JU�o�8���	I�d��)V1���g���M?F��p��\��hHe#HŠ|�t#�)J�p��ɏT0�ذ�LKK>B���DM�d�xР���*s���拤� ����+M7�yQ��R�����Y���#��S$���P� 6[���A�k�D>qB�:�@�hX����[�'���r�(DJ='���H��p����c����A���)�kġR��5��ƨ�´S�͎��M�; &u;t�.���Y����O����Qo�Bp��|>�3ݸu�1�?@T�YjG�B��E9��۷�R%��V�d�q����7մa�!�	j�]��b�<"�V��ĆC>V:� ��M�%-,`�2�ŜLh>�k��,LO���^�m�EV%u�y��ޭE�J�3Z`Q�I�&[�������.�83N�����	ߟ���g�9x0�A�.�,H#jx�J%$��AȒ0-�聋У| �e��'1� �AS�J��-�'�'yc(\�S���^�n�N<�D�֢92f��n����<qr�,Guj�@Q(ݽ_2����R�&�`�o��kd��s0�� 7!�ړ�B� &`���0Ӱg�h:�'��<��Ǐ�j?�1���ӟ@�ND��		Nz�8�%kL�C�C�I��t��'�Ƽ���1Z�*y��-׎I�c��YF��O��򔅇�?X�9�#�޻
U��a2"O05��C����PB&Z�f!j��i0p�#]Qx���g(M�Z�֠���C):�JI��f/D���I��8��e��iM'G����,D�<�"	�n�n5�r�T�g0��)D�|��#x T��OS�~�މa��%D�8��N�9�ճ�S;�%1`�5D���t�%P}�q��M�
�`9���,D��3��H�%�P
槈EUxA��g?D�h�$#�z� �#W��li$-�� D����.^�u�X	d+�G�ś�;D�,  F(�����@�r��aA��;D���D�"G�1gJU�e�����6D�|�� � ������^��Sr2D�|�A��7@HԚs! .�xX�U�1D���K96��\��)�e|>��Ӊ/D�@�%31;d�˫t^��TK/D��K7G��a�~Лbo"I��ǣ-D�<q�dǦ;� ��B�ǹ.,��#҈'D�$[3+m\iU��L���H>D�l�4�s<�]3gc�,4D( c8D�<��`�:�Vu�K�������7D�����6^z<Y)4 0l�R�m3D��D�hJ栈e�&	l\�r�3D����
׊-|�!�a�_��prN1D�����%��L"�* 1%\��C.D���烟�-��ckØ?�2h*��"D�� ���C��=c��XV� �,�8P"O*8�tJA�L�Zy��\�T��"O�r���fƠ�$Q�K�Y@�"O�yd�9n���D������"OR�1��6l�|�������$8z'"O2 �M�hx�)�Cͼ[���1d"OХ��	�$,�u��HJ�>��p"O���wckb�,0m@s��Qu"Ot�)2�0йa�]%W�d���"Oj�q��&��sUXy��"O�]Z᥆�_�%�� M1E��Z�"O�Ex�hV�@?�h�/�:;����"O��#�;h@`Ж�X3ku�4��"O�4���,�r&G
%�d$["O��p4N 9"���%�S��3)�`���� Cn�Oz���/�h(�$���̱H0�F*F��W�7^��l�ȓeNx�@b.�7M� �&��Z���ȓAC�e�7eB�R�RD!��RvhZ��y� ӐE��qr��Yq���.�*]�ȓ>
� YD�ڲ;0TqYT#�^�h�ȓGt(��#����|9�,��F�j��\��r`�ο�`iC-�:��]��6�����dba@�k��m��ȓ_��ɠ�>2%
l�fCD�n�����?��`��4A����(����ȓkk��vEǲXq�HF>��M�����kUv(�'�b�S͚Z�ϿAF��\ݺ��=1���Ǫ�s�<A��K�K���u�>`d��r,Q�M�̳��K�]$��#�'���J�� Fx�ȹp��Ƀe.�U��)��=���!H��T�Bsᰡ�2�_2K>�S��_�Yx���&�)��Q�D�D-���3)?�����_�:&0
�dAtqO�b�,�9_�Q�1�ŷ'�űPa�)$�R���y��0�iޕ�^m%�\�'�|`��,D�Pr���v�p&�
+��DX���T2m� ��5b���BHI� 0�qJ�c��$8���(^,�󐩄���X��nɈ!Z�C�!�:���6[��q���]�p92�M] �Y��޶��q�!�0Ԑu4^�qO�࠷�(rT@�W�d��q�'�'�F�0v�.�[t�G<t����3�N�[2%�E-K'w�\u��I�=y��cQYѴp��I�s0�
�IYl@x��a+��R.�b���1˚�W%� �G�)3��������uye�q0qj���"���mS�V)T"/D��ʲ�� ��bo��DW�0�d	�)7TE�!N��/�0r���dF��2Ԇ��'Œ0ͻub���K-Z�L�Ջ�5P~t��J�e�f�+q�H�wE̶�`�4kФmF�R��ō|P�`�P@�$K�y�ƄQ�w�^���!��a+����&?<��`���&LOTMJ�^zk(d���
R� C�O�/,*��â%:k(�,�1@��\�r�;=*�\�ד� � 7�A�� ��h�yY���<��菋}S��j-�s�lq�	�+���e
��"�0��D�v�H\��� ����6��h�<�T��W�R��s��>������N����hT=êY����H����$��X�O��ѤM]޼[� �e�R��U�
]N�Y�<���)s[
Ls@�����u���M_���R'��Y���N|�����Q�(� ��p�\������\�+��!h��"�\S��c����ŉ�*�L�P��si�5Y����)Ej�3
P0�\��ْvNBdF?:��	d˞�[b� 0���=A��]�y�t�/ăi��iH�� v�a�8���@������|#@�.��]���1�zIk��y1eZ�dA��\��ϗ5$���wcQ'$H��V.��a{Q�֛+`j���i/f+l����۷�h���L*~1c�|jC�̌;� ��e,��_r��ĪS�66n��,�IH�a&/,D��j'ER����ӄ�L&l�V�S�nӦ@j�bT�|���ɤm��|b��uN&U)N]����'"��Q���Lk��s&�0��=��I=f0d����<���V+3���!��Wt<�	�O.�~�R�݃=(�s�"�lD��O�42 !ލ���1`N�*@}$�Y"Oށ�CE@&��3���.>[��� ��<SL���fG��ʃ%=<O鉐��v&|�&�.o����'�E���4z�\�\Z(hzC�b�*���Ǖ)x���22�Y��MR,�^������=�qY��]�M� �+�+�8rV1O$��+_�w[��#��'_���ti<3��3w5�� (#EƜ�=��x�צ;�r�B�OJ�х#�s#�3�2'A0��wD.X3��K�M3w�b,{2dC	yA4���;r!��O��|�K�0wFp�FTi�2���\�.�|B�7��D�����i�-`U���r��&N��R�E��wa2����jS�K�������2h���EŔ1�:Q���h�R��1�����5z2�ƾd_PԔ'�j�ۗh	���mi�T���	?DH,��
��%g��P��6b�i2v�íl�A�`H
R�@=����Ń�fٸI�(����9r��b�"�\W�����3��6mN�[�^,��*?i���,���(���d�&]@�G��VLӲ���8�Bp�@OΓ҈O���3�k_e
1糟41L����	��!u��(So�7j4T�g�_g(JWl	 2�i0#FBz��y6���vƒ8��7h2D�K��dќi0�N�M �N�,w��A��s�����B�.�ސ�Rg�O�a��N?G40��L�(p��Q����r��6q��qic�+x�1�i��S��m��[�4B(5��[�h���R�4u��QQ����S��d�VΗ'Mo� ��	@&�(%˶l�vI�$�)�Xa�� Qðd�V.קM`�(��)Ր@'���0L{��z�Iܴ++V��ǃ �P��G����y�bDx?<�=�$H�<(��j�2o_܄��.(}_��p�
ج�N<�e�J�B�����v����Ĳh\ܜ���){P��H��-�^ۦ�΍���HJA�ǝ�jӑ�P�'Ǝז]�� �'��l�N�4j}~�0¸S�"D�I9,�(*ӠOuU$6͂�Q�r$���@o�鱎�s�0�Q切p[ �Ad���|p�*I�r�e�ǁ�vV  S���v�0�,��n�a��h�b��0�8���B؟t(N�(	�-![wxh�&�D]�>ѩa+��/�(�Gg �k�D4�u�R�D��.�+t}H��J��[�*��=��β0Q�,�d�ܔuJ�4a)Q���F03W���b\uH�0a���<3U?�S��ɺH����p'�*��H��!ʇdp��Ȳ1�,e����\pf�	���OqF�'	]iq�G�怜ps���joƩ�)ׇw|$��N	�6C>�FƜ�r�p7폁��=y�fH�"�ʤ�N���8 �74Ϣ��a�'M�R&�؎�HOt����Z�bZ~��t���H+'lF>����-A2/�!e���{��
��C����Z�V���1�g�-p�<PK -@0'�B�Z���*�hC4�K�'R,Yt�Q��f���D4�aJ��A�e+8N]�dC��:X�q�&O�]��˔Ō�4���gn�T�����dj\�WBB�1��R�AY�Ƽ���G�}-*�#�+Ψ7�܁�
|lz|я�
�G��(�f@� W\��Q�A�m�kƭY�eU(Q��� ˒B��0�v`ݘU@������ 9��U�p� 9Re%Q�CF�4	R5g.#TrT��Ie�0x��\8<�8p�J7RXEUAZ�q��٣î�s��ICU��T�	Yw�<�7��S^mY��w���c�Ȃ1�Z�Rק݂b����c�^�N=E|"���S��s �ؿtq��"Z($k��J��ѱc,r���BH�q����A%[�Bװo�$X3�d{Ӿpr�@� f�J�JF�_n��t����<�P��T| ��J|��, &A�?���9$W���F�O�}0��C�",���ea4���^!z6�K7�?Zv���*N�6{�"�O��5��*��P�+�2)��G��k�8i�V:!:���T�l��'�4IR ��%3���Ā)VsHq��J�'h���J�OވRG�n��L�ߩ���M�X�ɑդ��X�!�'a�Y�a�+f��Ӄ��G���f���p��n�!�M��q>��)�ǜg�d�!t�P�v 	��{���&S&8d�J��$ �����*�O�څ�S�Gy��:ȩ[Gbɐ�4\<�er���$���U�(�V]땃'E|���ɫ_OlѰ��uy�C��P��]�⋢`a�q�����0<�G��\	+�M�%l	��`)\L]1���.w�5��J!)���e 0@���'�1o�f0��]0��OJ�qDn���t�b�W\DL�:Ǚx䖯=���h%.6��ar�O�QH|���k��P�(�ch"xk�:%�#.&)�򍆗�:9��&1��j�`E:.Uޘ!�ɖ_��aN�WP��b��� �|m�U�P=��:e 8*RԈ9��|��wlA��IU�\���
H���,��'��4�g\6
�n�鷉�p�ڥ�T+O�t�Q�p�����X��\���$��^����hG:��DZ�O�X����"�PU���7J��}ҍ�7H����dJ[fԠ�G�Jy��x�#�"���	�m[}κ@�w,_�=>�B(\�'�.�*�'�ZF�,1G����K>9Wğ����k)qr���
uI�I��A��8�:�j�!H� ��7��i.��0P
W
Z��) !|Or��%��2%)����>UXe��Td��z�j�CO��Q�҇`[��"����b�,I��.IpF%�l����d�HP��ʕW�\A��S5LT#>1�,�he�H��
���Ӫ�i�͢=D-�DU:
IZ3���$гMtTuɓ��'D�a���"<A��gT�?y���2Q����;�T|b�Ќ@>��I{��5�c�&u ���O(�K�oI)8�c`!�X�E)C�*���0�� ���,[!�j,�¡���2�0��"*��A�N��/Q��b���5gL�}|� �ő�$����8df�SDA+��$@��;d�	���=<M ��2��^2���]�2?<�
��9bbXQ��D��~
�yÃ���ʔG~��
�'L���R�e���r^U� PiF�
 &�	C��ذ'�����a�4a�Ò1;�+9~�tA&!��$�c�L�1%ʀ�# I��TP��=������$�g��5Y0�K&Uf� T��ODppf������ΜPa��N"6��cq��f�4:!L�T���̾�A)�`�!Ɍp!e��$=��#�Y`	��8F���*6�\���pľi�.[����_���;�␃����ğp�뙾wJH ����.2�y� .��[v������d�\46���`Tʵ̮G��6�ġeP���Ά$_|��Z$�@x�y�X�C��!��s E�'Oe�`ۧGn�j���6s	�ô��k���鄧G�;N2\[��J1M��ܹf/O�RР�� Kx�{vI_0!�d˅X���@2�;d�hL���$�$-��H�5�G/�L�����=@��H�d�>�<|{���X@���^
TC�ѹ#�´�L�d�>G��	؞=�4p�!��
Z��Ư�s������F=���D�J��v/q�0�&1����	N�� �)s�X���Xh��$h���1�P�6~��p@錇\x�6��8��#����l@`�&l���q4{��Z��׉p�����~�. ��i*p�a¡2΅�����&
ů\/�M$ƃ9r�㰠�1g�F�Z��Qh�P\��Q�@.�����.�	�F�7(U�BQj��r��уi�VP�2��5��K�}ɒHA�'������/G�赢DP,�RB��|�z�I�N�Q�H@�$�μ[!�@�C�歪�'	�Փ&k�#��+! ɗD��@�<m�^�񁝼�p����&phhЮr�}Aת�H�$| �ܱV@\(0��[�p��PДl��)�5;�䄀p�qY��χH�"Hi0"0UAZ�]�jX0���o�s�HB -�&`Cr܃���M�n�s�G�=�T�橘���y��nמAYFu[��̝f�8��п��0�ޜEQVik�̟b�(Ԁ���"	��1�%�4%z���ɍ	��¨�DUZ+:|�b%��r�.�@r�OZ���#իpt���i�H� 9�U'U9Z�*�*?y&넚�$��E˭4��iБ��"+�Z��`�>[~��b���O�%����Z�g~�ĝƼ��V�F�/��D��	�3�\���,�hdHɂ��;�&�)Cl�	ô��F�j3�'Jp�松	,�i%��4,#|$9E�� ��탐BQR8�y���F�P�����	
Do>�h�#Z����G��y.'F�
 1��	ѭ.v�0� ���tk4�(Rc�_���L�z.
���#������k�u�Ad��0$k�'}��:Tm�L*�hP,\#G3�X����+x�7�ȓN�� �'XPzI����x��0��!D�pQE%-���'l�6�H+�Ad��X B�6y.6P'�������h�FX�6-Յ�~��(� T��v�EF�P�;w�ic�R1}��{VJ�<
l<�#׎Q�4Z,�I�f�����O
,��A]M�!r�ҙu�P�QA/��+�-��A1'�2�1�-��  �����Z>"���Ê6���:e�L�
��薦Ih�i*�M)(�ZuPc能Hlde�˓SS	�m� �
�h��{��p��h݊{�I��u�r�(H&���X0� (b�h�3x��h0Rh�mؤ$�̐NYּA�ǉ�F�ܜ��'���I��j�6�qs�B'��	`��Z�[����B�&T&e�4h�S�]��
%�mj�g�4H�(X���]��$f�ӤEi����f[l�u���t�DO����9���4�͑<�tA�p,
/F�����Α�H���sof�$��>J����AI92�ΝP'Ɨ2J����4�'����>�@'�V�Fu�k��Kh8A�QDE|R�+�T�p��E��6MN ���D?W��'i5��P��|&�8�Ƶ^�P�n�+j�T�PQ�܀�tp�Q��a�,���)����b�1�DD����=dU�i`��K#H- C�D5h��k&�+��ᔂ2�F@� �]�cX�	�"Y�N����v̘�aV&�`uJ�1R %�ӓ+`�ubX���I��·�h���)HgR�5�m٥~(9��ȓv���!�E�\ОE����!���$%�~�k:�I��´X' �q��e�.sqO��"DfW9>A:PP��O����^�Fm`������!A��I�}��͘ p�@KgI�j��Nڶhݎ�	:J!�"|�'��y��Ãdi���G
�|vJ�9i'q�<��[�y����'f��a*��#��S%�7��)�u�U�3qBy�ō�U�x]P��ރYRR�+�'�YR�`Q����9%d��S��V��!6��O�s����ħ���)�D�Pk��ڇI�2��EX?�b0s��D�Qk!�$��(c�,I�v�tm@�
[?!L0��b�3Â�RG��?� ���|/��'P�$0���59󺰃5DW�b=>a���kq�aQw�H�q�rp��'��i���ٱa�`��3�H�l���8�'Q*X�6[�r\�Z낳m�. I>Q#��2o�$Q�%눟�]Д��-�hm����f��Q#�"O�T�B��TЀ�F��vb&��5-'��9I��:�,6�g~��(�JgI4lxl1�W�y�H˓�i:��O�]G�L�Ф )�Msb!A5L������/�TЊ��N��3ơ�H�!�$M��Bl�e��tUtE�bN�
�!���a��|��P��&��� �!�$̐Nr�0pq)W�
~Q�D��
�!�F�I0� �I\3¤�dAJ�Lc!�d�.w	ԥr#�׶T��c����o�!�d�>E|�B*^p�ʂ��(q!�$£,3ٰ����yY���;g!�ثTc>��T!��)� �3g[�O�!�D��|�<�R��8�4|�F,H'�!�DX{��s,Έx܈0�Vf;R�!�$��3�@�bdK�	l�1%:-�!�D$�f̑�cY�F�f YƄ�9�!�D��\x��{f\�{�C2`�!�$��D�`���I�<��=���/�!�F#Rjf�Ժ��+�K]�!��գa�h ����p�NpWf()�!��6*V*B�R�e��,��h׈\�!�[5Anx����:4���AV�u!��T�XBH�&o�w�PZ4��z�!�dH�-�U��OW:���K`-��)�!�� @a#�ǒ�l���%�(�rLY�"O`��!Yh\8J�a��l�b��"O"����D�DD��r���B�TX"O�yRF"G�|~B�Qn��5�L�z2"Obq�ӯ�S(�24H�2˦""Ovly��Lo��I�B?/E�"O�5Z��ڪ_m��xɈ����"Od���-��aN�
�c��W�L��"O��p&i��n���x�]~�T<2p�'% %@��E�NB��ZQ,��554����)I�4y�2	R&Ά�����qjhl�!f9�)WD0!4��^@���B�pAI ��BR�6�ˁH�6=�Q�9�Ȉw����j�C0�A��a9Ų̆q6xc�4��1T�$���	S>.�6���AQ�1��>YD� ��0|z��3C4f���ܼ#�\J��\]�<#�^B�}*���	�4�xY@g��S_���A�O���	kLy� �)ʧ0�0U��#�(hȹڷW1���	h9 �����ӴvM�un�:qz{EH֮:Hc�D���'a��K�/#��B0F�
nN��@S�3���D��	�Y>�%�ټ`C���`&Ñc�(ٖ*��c�,ў'��&�[�gq��	��n�#�^�I�@�'Q�t��"؀:�d�3R�T
xΓ/*��Q��O�$�ח�ʥJwEAnή�s@��ZS|}q0�*tVʓQ+h�z@oK�6|��WƸ:W��˸'b^�#������ݤN�0@���-�#6O�?���_�@���'a��%�Ԉ����>�$XCEg��~�f�l��foµTuĒO�R 2�>/)��@@'h��5Z��O�7�(/p&��}Rv��
Đ���n�5��3NTe&�V�X2=Y�c�S�t��M���.�^$1a5�z$XV"�ΦezÅ3�S�OE$ԫ!�ǩ/�Tp�J�, H�HDd"����Q<�>����Hjֽ�Ԁ&]�@��)��'\�D��9�};�lG�O� Y�<"=�4���x�,P4yEx�a�y��TK�6�28���68�\�����Q?���W�2ҦF�O�, �ܖ"�"�R�6}�Ӥ�"Q�i!��<aPl3��q�"Q�%N*���#N�d)��E[�l ��'�:i�� �W���	T����)jÎ(':ִAəe�&�Y���6�j�z�C���>Q��<GFp#q�d�i !�[�<q��	$3��uYn�<�V��U�<�0�ق\<�hI��_�\���hSKH�<� 	IMB����]Ͼ��ЉGY�<A�%�	dV���DI?�Y@Q�y�<�SdSO��{��R�9$)�~�<���-�z\��
$\\T�g�b�<!�$7cg��`�����C��[�<��� ž�2�E͋KWb�'}�<q���#*��0���	%�����(v�<��aڤT�v��C�O9B�9ⳋ�[�<��B�2
дy6�Ͻ<c8��)�b�<i�a�
�� *�A�}�.5��O�y�<Y�kU1<�d1hTF��]\����}�<��-T4��l[�K����DAR�<Ia��d�F,IĮΦfMle�q��C�<	@���:ϺY� -��ntj�b�,�@�<q�JU�C_<�mБI �|�U��@�<��e�7=�U�j#UHF�5�W�<��/)S��" eٖ١�!WP�<-�� $e��?�(�i���k��Ԅ�."�ס�:o9�4��IԂoz��ȓ[���з
�Q߰�!3JQ�h��5��-����E���KĨu��}��#D��`�A�� W`��AO�
 ,d\�ȓj=<z�J�d@�[c��-��ȓ,^���o�q�|�CvJ�n�©�ȓ��ĹcM[^��	!,�N�D��3B�}rc�ȃ*ꉉoE3/��y�ȓYl��B��Q#p澝�T��2 �H���S�? x�R��W���� 
�y��4�"OD�Ոы	���S�A?�̵3%"O�Eh�g ~����ՁG� Ժ�"OtQ� ��#�������%z�x�g"O���U(�R�-�1-ŸM�t��"O����8����R�ݩ?Z��J�"O��!I�8}�L�)V�	*v�L�0"O�Ļ�ߌk�h��F8�� �"O� �欘`��@���9 *V�HC"O$@��G��4�L�۵h�9zM��"O�x�E��Y�\�6\tg"O���1cњ¸eR����3�"O�L�g&����E �Һ�XL�"O���ȱ+J
�cqB5W�> hA"O�ሰj�7� �F�ڙm.�c"O�[�	�n��\2�"�(F(v��"O=�#aL9oC���bT�F���"O����&^9Q0h�����k�"O(��'*B	X�@��!�jΖ��P"O�����-K뚱 �E��|\H��"O.a�W��*�>�����'5N�@CR"O8�@l�!p��1�����"Oܕ�S�IL�-�jڿi�e&"O�Q�+B�C��H��G�H���k%"OjT�V"�# �,����|�䴠�"Of�kC ��dP��@�8���"O�
%�S(+�H*���I���q"O^���OH�B���۰�V,\�t�"O&��p�֪�(�2�G�y�mb"O���t��>�٢%�A�)���"ORiQ^&x�B�S3	��U��"O,��jV82m��g^+6���B"O��`+Q	u6��h�>e���"Ohaq�(/'�@Ɇ&V�q2@�s#"O~�pW��2G���"S�x$�¶"O�x7D��s�h���`�1a^�"Ox�D�в&@d��
�~��[�"O�-��Ǌ�XE�Y��nҪUd>�p"O��5g��������
7"O
�j���qj(��a�֔�� "O�٤�
><����e`�;��! "O�¦�B+#T�҂iW�u��8�"Op�0׉�s��Sb)͙5�
���"O�M`"nS9V��]3P�P���j0"O��!��� H � ��X�<*�3"O�E��D�y�d�8dO�0P��"O,�z�H���9��K(���"O��'�:0��"t���O9��0"O"���h:=AteuHDa�yH�"O�T1ҭ�A"y�e���Mۚ���"O�)r2MI(iሄ��"��J���3"OVYId���� �@h�$��u�r"O�;!�H�sx%��Z�T� Ay�"O|����(t@��wԧFW�g"O�!R,r�Х{�G�c͊C"O�[����JS���� �!쁛�"O�A��� ڐH� �9U�z5"Of��!FP#)�n��!���#Q֑"OF�k�f�o*QCe� ?��"O���&,��ʘ��}΄��d�e�<Yĩ��-Ͱ "6�Z�iJ(��d�l�<9.��BF�	*�(�(���g�<��܋�7$�i�D��Iظ�y����V�4���ɓ�W���6����y
� ��(�c�.,��H�\�w�r�yD"O�u"ց��1@-��L�T���2"OP!P��F;^*�"X�����0"O,Rwj�%gf��у@��9�1�"O�46S��;%J�>K�,Pb"O�(� ҫy:��󁆊��xb"O�M����7(^@UH�F�0���B�"O��c�w�����O��h	�"O��!P��8V�����5Pr��"O0��,B��t��2�1I@	�"O*�ӑ�U�"��!!��xX$��6"OL���K	o�R-y T�rn��`R"Od���S����,[�I�-�"O@�2�MXO���8%�g�H�"O���]��y'�(!�pc"O�pǉֵ�,�V�3�Z4��"O,���C�Sp>r��B%`�"U�@"O��  .��'��hKi;qt$��@"O��i��P�3X�8��ر����"O�
���E1B�����j$~�y "OtxQ#,C8A@�dj֤'��t�"Oj��KD#M�$�X�U�p	�"O��5#���j�	�(ѕkf\�1�"O����D�Pi���[�~��=�$"O��I�G�i$��t���J7�)�R"O�l(F�L�{�Э����4�~��"O��
�D#7
�{�D�B(P6"O��JT�P��p�x$f��:�t Q"Oh���+Q�kQ��sORk� �R�"O`x�&�C0=�h��.��!��:�"O�`���
� D���"�/q�E�R"O��s�e �#�F��b�#<�|DB�"O��U�$��h� Ş��"OZ�P͟�H�s��#�rS"O$�b$Y�~R\�� lK�c�l�b�"Of%K򇁉S�e����p���k�"O0��-ا�\`�l�Lc͡�"O���B.:�P PP���;[baKs"O��� �o�V������^�����"O~(H"`Վ-�6����^���R�"O6�X���L;Z�A˚
�*��"ODicN�2)L�+�*٪6��uj�"O�t��Б':�ݲ��O4p <���"O�����& 2�
dGR�	�"O�BȒ�:r��F]�D���Mf!�ٿ�B�����dE܀���F �!��B�{��� � �sBܡ�NX�\!�d�@H����g`������!�dU�o�Hi���B!��џ)!�B�[�X,b�[00���7g�
)!��0c����ڮs����'L�M!��ʎ|m�={0lD4�<�H��ÏT
!�_�g���S�g�hn1$�$K!��܂5��rᢈo�〘�S!��^��=	���/��Sg`��!���R/6ـ��� ���"N4!�$� �t��ָ.�8:���	S�!�d�	;�qvK�Xl�!��۸6}!�D�pg"�r#ӆ�J�@I�.W!�$�0��1Є���V���E!�d<�6,���6=�ԁ���	�7C!�D �0*����*�<lɆ�S�:!�Č�Ԩt��l�6+���c #!��l�rq��!6 ����얂.!�� ���§�,T(4��-��m���D"ODA{�� x_�%���ކq{ "O^%�C�
��ya$�B!�d���"Ob�*Q��IL� �g�k��`"O.=AF���)G�,�R��0'4�§"O�M�QjV�{j���P��"D+t`��"O�)���E�F���ɃL�8�t�3D����+	%n��0�W��!� 䋥�5D�,�2.ѿ_$����4$�ĝy�B)D�����_�`젨��(��L�=J��<D�Y6�g:�Bg8Y�p8�`-D��
�j�3\����>0E��,D�,9�
�a�ڵ����W}�=��&D�K'�˂g�~ {6�*?�d�b(&D��EL	+&�L� 0kM/a�\1 #D�Y��0i�
8���W��ҀQ!�3D��1��@9|]�!@�*��v�n�g+2D�l�#��N}�QƩ�F�� dD/D�l�6��`.#`c�b�&� �.D���C��b�"h@����h�-D���	ђVٚNIf�[��'D�`+��������:�Bf*'D�T���D#6���(��K� �x0@$D������+ �\��o��c�B\�0D���vn�:J1���eJ�-_p���1D��K�/H9s0�d�ągxPx��:D��9%`M,��t���=��b7D�l
g�F�^��� �ׁ!����5D���wcŗY$
p��O	t\�ԫ2D���f"0c@��!Ȉ)�<ٚ�F>D�|�2握�.�2㈌N���Cb;D�Lb@O�~H���h�>1����U6D�4ss���4UЏ	E��|2D/D����cɄL��ɉJ9`(�P���)D������$��JG��=���*D�4���^�0�0}IrbO�-Mj �'-'D�8�3EʵK�6�3AL�G�^d���1D��
��ڭGĖe�R	's�(� �.D�@�0�   �����ȓN&z���+����C�+M�2��!�ȓ O" ��" ���EdH�u֤��K�HK���B���e�ͫA֦d��X}�l��$�!et��Z"��'.>���D����A�&B�
F��"t�p����f�ٗJ	h��͹��<�	x�'ۢi��C�L���!@�+mB�'�P��S�S�T��T.E' c�!�
�'Sڔ��A�
�,I�C	�R��Q�
�'�4{��_�W.Y�S��L�l��'1z��a!�/\ Y��\q��U��'���"� ��\���a�AplMj�'��u��X&,��+��GR�U�'"����@�9��c���5���'7|� �9f����Ąڎ+�Z���'��l�C�#L&|��%X<b�'H,�Q�L�eB࣢�ߌ%�`yZ�{��'����&	��`���G�${���?�S�)�x��1��؋o�B����֞vD�'���j���-������������jx�@+�L�pÑ��>Y�C��Z��dRH>E�tD��2E)@2^)����� �M+�(PP�*@N>��zc>Ձ�+��r0�b�Sy���#��X�@)�a	GC�d�u>M��!�*uC8\��E�>
��F˗49�Z'��*\���j�~��O>m{ O܂O��Q�I\vx�)����(@�d˟5���h�'ޢ;�l��we�i�t9�MɁć�"���H`9�T�H��I~��O�r�(7n��a^�i��%��Ke�P��Wr�l���i\B&H��0|
#��B�O�[x�,"�&�&@1 ��a���?��Ǎ�rn@i���,v�$���B�'�~��6i�0�0�j�mR۟yb��l�P-��<��b3�'�U�BI=��@takz2��t_���5�D"b:\ۃ�>E�d��Q��	��"`��sPI���M+DJ04���J� ,}��	�{��K�ՎRet��&�)������:$Z��'S��)1>����`JˎG~\4[6��/
	��/�x~�L�_���ηvDA��i��l��*4��x�'�0<:l�i���iM�dZ��k�ちT����A C�E'�	+��G�ō��S�O8��R�!P�yu��`�k�0
TH@ �4W8 B'����~)�ȟ� �ipA�/4�6�s�˛mgJ}�ن���J#JSz~�-��d��C�W*٪R2,9k�%&�Be�'�f\z�+�3�V�gB��# �K3��4�"Mt!�$�q�������-pv�@����Et!�DE�|I޴@j�2\��*�iR]!��E˼�@&Z���9'ɑ5�!�)��
D�A�-T�����We~!򤘜kd����[�=��&�s>!�d�s�����i�:q�.4�VÛj+!��D	;b�AĞd�D-��C�$3!�d�S7�1I�Î�+�<`�a���w-!���xPL1�5�Ԋe�� �c�j!��ώ�0)*j��X��\@�U�e�!�$L!���A���'V�,�ꕭ�4�!���;]z|iy�ܔU��-��A��-!�S?gdu�� �*�����Py�"o�q�G�L�DE����yBaC�$x5a���"H��]����	�y�,ʌW}���H��6.�X&�G��y���[AD�Q$������F��y"�L�]��a���'�e*vű�y���Q`Q��%~,JU����y�,Nܜ����w��2���=�yr�?U�Z(1�O�j� �D͙��y�bʚ%�p�욱fR^�IP
�y�G��+>t4҇�_�V�t�{�-��yRf�'pK�D�BOȜ2Y*�#���y��Ƒ*`� ���wȊ�x��I0�yr(
;�\d�3 Ri���A�3�y2o�<�Ҝ�p"�2^?�����y"#��a�>��2�D0"�/�=℆ȓA5T)V/>�I!��u�V�ȓ:*�i��"`�!a6(��@��iÄ�6c��2/����I@�`pl��Q���'�G�&�0`!�8\�ȓ6�vJ�$jC��c4e�!I�P��ȓ��ɰ��J����ϛjð4�ȓ[:���L
J���Y��[[0
�ȓ6d��pi�i`��gO�qӎ�ȓu�\肂C�U�����J�oQz��ɼA�b㇥4�3v�	]�4���0�,wD|DI���T����#�.$�,�H�^�/"�ȓ\>�l��c<t��QcO�"�`���B0Sك$P���$K�h$ܜ�ȓ;�Z�;ta�~�&,���1J�]��n{��(�C�')p�&�)
Ԛ �ȓh��p���YѸ]	bݪar\��2�P�"U&5q$�� �Fx�Ʉ�A��Bm�b���,��@�.��Vv��D�:q��ts���VL�5��0�y�c��t:ՠb��(-��ȓV25z���,z씘E�D!y�$%�ȓC�r��q$O�"N��Dd�bS�)�ȓiY 8Ղ�q��!C�~P�͆�#1���"W$8������6j�ȓD�>A1��ؽJ���V,(-������8�!��ߣy��C�(נRު ��P���H#��
w���0bg��_��%�ȓ@Ԟ��e.���8ҺЉa��<�U�7	i(FjąK�B%{��Zx�<� �U�T�����)E,�[�C�r�<q��'W#� 3�:o�`��It�<�vMEd^��  �] ��j��Z�<� yP2]��x5n�
��ht"O�Qqbl�!�NY)�#м]P�d��"O8��dGؙ*`�#�Y89FB$�"OP�Ղ��8�FDȲ���|�"OP�Ăߴ��2�jԱui�<2s"O�eԃN/y^��Ш�OVq�"OD}�S��WUN�.��('���y�#����c���</�>P��I]'�y2,ԉm�� �怺7β�Y,��y��Q�l���B�ވgo����'�y�^V��tA5�DY{��pO��y��R�*�+ݷW#��eޥ�y2���e��`AHIxs���y&N�wºȒ!;G�ʄ����ykͺ&0<�֯�1�B�G�4�yR��3>(�҆;	�6�şY}!�$ķSJ]	b 6NӜ���gգ3{!�d��J��%E�k�����)n!���ކ��g�M�0�N��/^e�!�$)�(I� ��-|�X �uh�,�!�䞾!��@T+x�!9�&U�&�!���]�N�;��_�7v�1朽kt!�ě?�B����1����Ď]!򤐯��葆�@��P�7cC�!�D��v�b�	�I�2Qb�����!�DĊ��aU��[s��r$����!���.�>�I�l��7`�%����!�$�&[ȘH����{F�P{�
��!�d����s��b@���A�H�v�!�DL7"�B��A�� $M��Y�/Q}!�d�d\$�%�Q�AXth��D:[p!�$�:$�h���("$MA��� !�䛜PLIA�R�+��Y;�䉼\�!���8���B�b� Oh5�1�Q�r!�d�0z[�a��Q�BP�7��o�!�C7e{��z,�+�eEP{!���$wR&���yWtXG��J!���=l2�0�,a1��)��/M!���,a�0�aEG�2ϒ��c�>w5!�D�sf
-[5�ŷY����0�7,!��ir lk凁�	�l�!,�m�!�$��I~�0G铖A�Xً#E�#�!��Э:E(@�K%j�{��қG�!�X"��pR�&Гk"ʼ��Bѡ+�!�zt��*��;����aR75w!���}
�����86����@�:4Y!��~�l�&��z�X�/�1�!������`�?J���g��0�!�DܟPA\ͺ� S�-U��� ���!��Ʈ�F{dߺW9(���H�!�dV�&�P
q�I'���K@�rd!�D@(!{�y[%��\Pа�L�y4!�$�%O��RqH�J�1iV�]5%!�D�O���aL6���
0�Ӌk!��SOJȐ4LW<А�g!�>t�!�$�\�8���\�l���¯+�!�$�e>���Ɛ�|��.]/�!�&�20Id+�2JC��#�S1�!�E�L|�YPK'3ֽ��U�rء��9\����I�_�|!fA���y��XG9z�ѷ�:������y��ŭ_��8b����3���y�˜,�~$�S��
�m��c]��y2#���VJ	��3���y
� ��c�̛]2T����F(��"Of�憖PD��V�F�tz|U��"O��s�M8i��L:�4(_����"OL�cn� <$yf�D[Lv��"O��dѧA�a�G��Tڊ0��"O<͚􄏄NvU��OB9}��`��"O`�*g癰D�l��.���N�Y�"O�D�bIǯD F�$o�%+`mt"O�jU�F�B+O�|N=y!\3f!�D v�9�W��%u|\s��ݓT!�D��LLq03�9\�h��cٚ	7!�$�b���zP�)$Vư@c�ͣ�!�D�+sKf�G�>$�}�SAX,:!�$�s�ʐ$]'Y��+'�͌x�!�dȢD�>�A�!�:u���#�k��l�!�D�#!�\��E��
'� ���	-�!���s�F�qe�L/x,�x��C�$�!�$�&@����
R�$#��2`!�d];�(�wɞ����u�52Z!�$�$�l�b$��%��D�NQ!�͌N�@	��&̘[-�x�*B�4!�@;k��ܐ���=��炁'!�dJ�}���0g��u$ZaA��-{!!�dϵf_H		H/t�P��L0W!���v�:csꐭ,��4$X#O!�DĞZ�VA���y:@$.� !H!�Ą0U���C�Vt�X#����6F!��M�Q�d�#Bl����GlƦfQ!��Q��EK�+�#�`�8��7V4!�E�:+������P����U�>!�������A�sh,y'J��}i!�D٣%!����`���,� �W�mL!�d�oD��y�V*k@�h��F�!���)�d�vi�
kx�!+�	�)F�!��0��R1L;7p ��P�!��?g2H@���Io�ܑ6n�D!���hz&=2!���,UR�s�/X`�!�Ē�J�A�(��Lصplի?�!�d<Vn�	'BV��ɐm�7�!���&#ؤ���P���I�.x�!��,'�&Y`���n�x9qS�!�D����E�6xpv�9P� -!�$ڍ;�(���
k=t����	�!�D��e�p�t"ǘ='΁2��
b!�$���-����*��x�$�!�d˄gW�����1:	��'��!�d !���J���7�ə� �4!�ߙid�Z'-�D� ��
!�d��E���Q�l�1�|�P�*6�!�ę
Den��-�}1�@si��_L!�{	t]��B��7'j�;p�\7<!�dA�D5v���I{*ԉ�f�� ��C�	�"��ݛ1H´����!��zC�I5D�$T	SˆA���ए�8EPC�	p��d�cD��*��aF�)|�:C䉩e�p��+�[۪8���(f\C��#��UʕgbP����#*OB�I�̘3�g�9q"+���6W�B��&q6��c�^9L�⳪\�8 dB�	<��@����tJ�sV��?)�B�	%A�n(��ӗl'~!@�MH��B�I�MݰiȰC�M��ҥ��-ibB�	$ef��k$�/kz �E���C��O�T��9&������Q2�B�)� Je��ޅ5�Ƥ�q�ǚOyZ�#'"O�]��hU�( �Q6j�|�� "OFIBNG[3�p*�BSa���"O,JD��0%��2��1^��5"O�=@'��u-(��*F!%���"O��S���:�d�������"O��k��U����3�M�jݜ��g"O��ar   �"O��P�.��=�
�����\�P�"O�X0���b�5z -#�,ɩs"O.10@��:Tt*��$7j�Q��"On�³�N�����U��'����"OƴI!"�S����7�݄X�(!9V"O�D{k�� @��y�Fě"O��)`f��_��1��E"�.�I�'
�}��E�;� i3G�7:�(���'��{AhP�ti �����<K�}`�'{IkFoE��VP����-^��B�'�t��Ff�<`�`!��q���	�'�푷ĝ�'�bH`A�؍�j��'
���%e��W�]��Дhg�tb�'��Eh�E�|����
ظl}��	�'�%���)K�Ҙ�僂�h�aS�'��ȩuʞl����[!i�]��'a^0Q��jdaĀ n�y�'�u��o�m~�s���+P�xX0
�'"Rq���-�\�K��ڑc��(�
�',��-Jx��
 &�;Y��i�	�'�0H�u�F�f�Z�##)U4Z��a	�'d��J	H
^]��i�P|���	�'��h�@I�9�@�2���O�|�<��*��0H*�*�?I"�X�CV�<����(�8�)�Bn�$��3ςV�<��m?x��Y� �O�NHA`�P�<)�%��]��,I��BBz$y�Oz�<�Q�ɰ+��S���TDp��6Éu�<!d�> _�r�k�Z�ڀ�c��q�<YU���i�ڝ`"d۲0��J�`Hf�<)䆞;=pd11�*	:��
�D�a�<���\d� 'j s�j�Q��Y�<�͎����S�EČ;���T�<qb<>��Z'��X��aY�<9�� f�����S�=��f��<���? ø�;B�;c�dq� ��<	��"V���D��|T�DbU@�R8�����o��{��,_t�=OP���B�3t�P��M�R6|��P"O��!�v�����S�:'Jy�t�xBÍ�qvN���	°5��R�^��)AZ>-3`�ʣ�N�X��'v:H$�>�OFȃ�l�)�MBn[�Q~r�� ��E�(P%�m�@e���d��C�>�����lb���/Y�C��YG|b"��tf�1�P�|�'.���`�JM�M&TL��+Y�o��N�iw�E
^s��'ڞx��mڝ=?P̨��ӂ?K�S�'ޮřSCD�m0%�O�Sl,�s�<`Ў`��/��Nn�͒b1=��ɺ��9Y���dZ��ڽHs/�2,S�x��@&'���g_����� K@L}[u�T�n�%�.�pb�OW �+E�����u�x��^�����	�;b #�`� a�  '%	}ɰc!�2~�a�FJ�~��3��I7gZ�9 ��
78�Qd���^pz">����<�Hx�Vg<��XS��kW��z�}2�"W�R�66MJ�w�!XR�N�Il^�	�gLL;5���43":d�ϓR�L�p�(I1`U�ӧ��*��a3 1"��c�'�Lc�H'a�P�&4iEh<Yv.��2, 1�	O.1���33ln~rjS�_eR��'f]��9J!F�!��ɘ`z���;
�20��������w  �H
�~�k�h�"@�FS&ml��MM+o�<l�ül�0aƋ0�m�&�"~�$o� �x{f��9�	
���O����[�K�ȡ��o0�4�2zq:���(2f�ؑ�����2e (�z	דia-��$ �e�BG
L0�x'�`���N4�|���)���@]5|�r� ��kjC�	�ASڐ"%\�>g�D����w�zM(d�My�䉸o����~&�� �����"{̐�4��l:�O��p&��c@�t��*ފOޜ���c�8dHa�K���>��2P&�1�"+�	�܃�L�oX��K�W'(�']��
�`((ܤ��G�M1y%�����9D��3֪�?e���5��Rqj81 5�$P�7����� +��FXC HP��x
%,ZVx"O�t���W�He��¦D90��14'Ʌi|�'pj���/�3�d@��@Q�4���&�տ	g!�DE&
�~����8u�b�M�"�����Db�	��E�f5�'�i`�A�̍B��F|�P�g����emÍ?OД�AX>eY����.`	R��(�*܊�4D��!w#T�3��Qa�
�$1�����O@mC�_t���kB�b�\�
5�	3R�f�ӈ ��Yc�A�"�y�̜�L��)�����R�R(_�ȍ�ɐo�E��N��,�*�⭟��: ���4�O���!��f���F+P�yIZ�+7�'�x�.��\:�r(�h���R��ʙU�&���� u�P�O$��G�a�g���v��P��`Z6�:ܰ�h�QR������ �|Y<�k���=55&����"��Xc�xƂy3��9k7)"
�<�yIˉۀ�#��
Z�o�-n�QA�!�x���|�2��4%�\ɃBƶ<a2�ՉO8����g��PmV<#Yz�<��)5"S��oz�t� G	H}�ј�Q�#��<MJ�O�1�����i�"��P�D��"y��q���W+a}�Λ(B�B��#$қRK	w�i�񈑊�`��ăU�WL�OL��	ƨ���ē3d���+_�x�5@�,-0v�Fz�딍5t�����o�'�! "�W5,Ǹ�x�m�%j�VtI�(� $�`}�"�;�O$T��C�;�MV,����*b�';@�k ��`�ɧR��d�vYi0@�<A�jbq�Hsp"ͫ+�~5p�j[V�<9�5"��1�e�#�T����XQ~rlG%2��w%ɰ#F�8�@|B��|���/����M <6a���R���*�D
�"������E�c*�6o�:�Jy�M��|~�'�Ni8��N�g��Ԍf��#�O�ؔ�Ŭ�����L�u�r����)�13;�m+���4�x ��ƥ 4�#�c\6�p?i�FZ�f���3!,h��`��<�u���X#��6}��IC�B��w-�	y�bU��f܁,*!�$�`�.?.~`#*B�p��OX�
`�^����i�8E�$�Њc�^�:��1��͆�	J�ry�iӳ6X����)m��|��-�e�f C�
O��B��Pw�VZ�%SL�d���I�Z� j!��A)q��H�T(��*~�BD�3t��Q�P"OP�@Gq1⹛G���M��j9OА!�c�|���L�"~�&m
�v^���,�A��=[�L�k�<!��~*��r�ٜ준����M~���:�U1��]8�x��Q�[)	&N�2)�x�X#6�OԀ����E�F��eH	.,t�#�K���,��K4$���B��x���;�!�	w-���@�9�R���s�d?�S���QP��zr Y��ϫ@;&B�,_�J1;�e�	�|��J$��B�+w}b�8c�8�4�c��Vl�C�IF���c�D��氢�i��do�C䉲N�^h1� F��1��'7lvC�#���CH[�zG��� �Σ?�BC�o��t�B/tȩ�c�
&�TC�	z9���ʂuI�q��`��LC�ɽ9R|�R��ϩ�;��s,C��k!���ţ`����W�[2:C�ɯuJy�w��1 ',iZ��_=Tw��J���g�;z�>�[.L���.[���´�H�C@��ȓ;V,�	QeЈu{d�#wI3$��D�s��P�H��'s")6$�;�(�3
�T�����uK��!u���~LJ�I�2�2`d�>6Ȳ8С&_�?:�C�)m�\	i�ᐍh����Q$�c�ش�T.���F�S�F���R$�6X��&�[NH�B䉅l�DɓtlϢ!F�Q7G��{ejh�&U�K�� ���D��Of�1"��� i2�OŅ��U"�"O� *����u�XK�ؽ+X�p���-��m8��ɴ�p>�@B�K2���ሐ�2y��2�Lo���X4\�:�U�c�O֥��D��i�A@�14�a�u"O�	�F(�2]����Ϙ�V�)��󄘽U��uƞ�D����;hܢ�b�+��l丗"O~�w���]hjIYg
��?.^���s�0��M���/7�g~�iNFΰ͐4mR�K�2�(K>�yB+�C��Hq�ʴMp�p�@��� $.Ќ5�����=k�k�����M��G*a{��Q�(����'�� "a�L$dYR�{D��*�
��'���a��3 G|IP�e�0�+�'�`�)'.����I�wC3\|��	�'Òـ�$�,7D@�J�#�%J;���'�nU���.I,b���e�JT�
�'tub�*����ã L�0*	�'� �V/ī������Fw<���'o��9�@Ā<�Y��R�/�����'7ڰ ҆I:L@���n�)$�9��'l}#r�_|ƈ�@B�%6#\��	�'�@C�� Xup%�6;�`���'5���)I暱ʇIS�M�pu�'J�lI@o>^5(�J )�,�ɛ�'��!J�	�	�DZe��:&�Z�[�'�б*1H=Y֜���iږK�L��'���dZ�8���d�Oۜ=+
�'���a�͞ �`ೠȊ�E����	�'8�a�0I-+�xЀB���1��
�':^��2�G�70 ���/�R��	�'�V��QC�&�:��Q�D Z ���'=FM� �I#FL��Z���%#�'����B��"Fp�jd��,e`����'.B��"E�z%�8��N�MX���'����Z�֤��m�0)�F�{�'W-�a�� q��iS��2 F�9
�'+� ��fߊ{�ЉE#�u梐r
�'�,����D��Y�n�c���	�'<��pv��KhԈ�%��)�b]
�'��X4U#�q�Ŧ>p�A���3 ��(�˛R-�I�%f�=�ɛx�pAt�OMB,���G�p�6�_����a�iȅ��)�~l޵Ca�$H�d!p���X^
�����tL�L�r��?yH�-VE��-ʰD^\lj@����4�`1Y�'��bC#ڮ_�a�Āͷ5Z���D�w;�xJ�ʙ�m��ɾ'�ӑ��T϶i��ӌ1���E�*2T������rw��d?Y�L�*Se�/\N� ������Ih� �3L��ii3a��,��Œ�L�aH"5�T��V?��.v�ӧ���5����`tz�����	��pIZ�<�O,�=�4]��AHN�?`нC��T+t�����2}�
Ei���O���o���c�	P`8�B,OJ�=E����8Ed�G �@��D���_;�?Y�{�]�-̑?�b�nZ�>(�ܣ6��uA.mpw�-�: �Q�����: @
%5���Z"�(��U������ӉPh�(�jM�4�*�E��4W���H����Z�zW��\��E���^����h���Q���O�x���j�+r�x4�ۊXl �O DyR�>]��)��p�Fܺ�K"#���P�(OQ?�p���#� بăL+<�:5����'>��'ya{ba�B��I��=�0zcdL>�y�N׬u�]����*0�J���*��p?w琺]�L�2険w4("Io���Ytŏz̓o���Qd�/��$��)�&[l���Үn4�"��>$��%]�jT9TF-�gy���Yސ��ŗ�k1 ��~�Ȯ.)���y��IM4�:��1̈#%�I0��3R�@뀋S)6�������$Y��0�o�h�tQ �ۭ&\2L���Φ�]�0��Oy� 瓗*��=�B%\ψ5#����y�'c*�rV�YY��J&hNf�$�8J k�7V>LH1�S+E�^M�%�*D�� YY )Źu��Բ�.��=�$���"O6����&$��L޶|�j��"O����W��  H+y����"O�-�цHh��z���m&`���"Ot�۴�F�_Kt�����$~�&li�"O�|ڄ/�|�`|�kH����""O<Q(��.*�}�(�H% @��"O���q��z�s�-\�w��ə4"On0p �&6x0��l�Cʪ�ц"O�Y0��P�6�8d�'h\,["O��3 h�l��c'*ܒ4 6���"O�	+�-.lVZ%*�;u��d*V"O.��j�4�XH1b�*v�Hݐ�"O���D�%]�h���A*;���E"O���g�!3�ga[�I�4�C"O0�GM��
r��� �^��"O`:�bb6pX�U�R�\Au"O�yR��Q�P�R횤��c�����"O����.�lϼ���� ��0�"O04�����	�\�p�߬8���Q"O^�З�I5S^N��D�Y���3U"OJ�� B�6=�� �� f޸�"Ob p�Y�4Ң�� 5N��"O^�x��4��RP�כ}�ԍ�f"O� ���B����/�t�1�"O2y�@G�u5dU�p�@?J����&"O��u��h��=Z��G�e~� 2q"O�0�F�]o]:�z�ԩkRe�"O�������a���K�a'Z ��"OD]
��P�=�ĸ�J��N�Ma�"O$Qó���W��ERr*R�W����"O��K��v�`E��*�c����"O�@䔋v-h�*5�H5��'"O�@k�#
�]u"�8�g!q��<��"OnU#w��y����a&V��Z�"Oh�s����P��U�!�Z}��"O ���<H����B�FW�r8i�"O(�� � c���9G���,��#V"OlM� b�C��d)��._�^��u"O��е
@� a���͸m��3"O��1N>P�64�@^$*T��3�"O�U� G<3��T���|���k���y*5�vL3u���z�6Y
�����y�!׹:Ӭ�E�
m�����?�y"��=�<H
U�����;dOH�y2NI-hh5�"�6FDpY[$�\�y��̀[X�  OL7	┙t%�3�yL�,H.B�!�9T:T��y��ƾ�`6	�(���!�a[$�yr��_@��0!�� �!��yr*��Nf���MW%O���b/�>�y�+8b�Y�E�"�D0��KX,�y2@޾u�:Ր6�
��u�1�F��y�72t�"@�����@b����y-T!p� b&F�&2dI�#��y�.�u�@�C�T%dbr���*�y�L�\�2�Ռ��[ �R�mͣ�y�""dS��_5B����C���y⡎�댅 eP(8b��y"�?\t��Y ��3d\��a��(�y��O��t ���̵��x�'H�yr�G�	Zl��E4�d`�%A��y"�R5�PA�R@B����pl��y]�bv��
�)G+v�>@X!�Ƀ�y
� �hql��s^��-A�+�!Ca"Ol؄ɟ�l�Hx��.i&^tE"O�q�d2%�^$h4�7P&���"O�]ٗC��,'�����7��L��"O��x�]�uێH� �ÃXX�"O2���Ƶr7ڱb��&p��8�F"O��G�+"@��%hSj�&�h"O�qB'"�,��e&�΢�҆"O2�!W�(J0x� #&`��"O&��'�N�:2��qȓ3I�|��"O��Fl�n��aQ����(#"O�1`��ƏhD�!�D�^  ��"O"�DKR0�@A҂�	(�"O���OK�x&~E0�(+����"Oh���)�I(�ı3+��b`e��"O�DX�, 
K�R�cG)	k� P"O �y7�o�r񋔧HPT>�s "O�sF�G�bp�ԫV,�9e��12"OF��U�@\�B���*�� ���"O�Q	��|�b�A�
�/B��a�"O,�J���	h�B����"���
E"O
\��Bm��M�P�r���"OđB�I�"q��SM�#`mZf"O*S�$w!�y ���O�@R"O���GD��M�r g�AF����"O�P��'ߴN�]�`��a��""O��b�IֲC}���S8��5j2D��b-�?n���B��l�I�t�"D��:��µx��X(���>��-�U�5D������ei�HL�Qe��n4D��0� ���͚BJ����zg�1D��c�I��6���çG2o�����$D��#��S�d��3�ē4;:�Y�&&D��%�U�m������N�H��ԃ'D�,{�"�9���A�:,"�XUg&D����D>X�� b#H�Xʹ�8g-%D��`������1��J��:mrL>D�(x!�ر1��d8�	��8���K;D����ӵ�)j�oC�6� �Ae�7D�$8��#s=P����0��
8D�`ɖ�R	#}J�22˝Y�r� �5D���R�%傥�	�Z�B�qT�6D�� םu}����#��=R^��5D�x��Ðþ��f�u>M��"4D�01��T~x�QUef�x�<D�`��N�J:�š���-��1�G=D�d��A�4=�y���^ǎ� �;D�DiSj�mS���m�������;D����6�Z��k�c �0�V�9D���w,� $�Ԛ� �`�~��f6D��p�� ;��#NO�*

4��E3D��@�l�Y���ߺ4��*� &D����S�[�=KEk(wD1p �.D�	��D&N����~o�-���7D�<i ��l�t�JP'I �f��E8D�z�Z����ʊ� H9��+D�(ؕ���ӄ���Ά=hT����'D��Ռ�19���Th	W�@�0D�0鱧['���+F �=wl|�J4D�,��3uv�pE��'xoV�y�=D�$0��g�����#�r   �k&D�h(r��Ta<sPC��
=�ɠ�.D�H)TK¼��9r���L**HR�A+D��KCL�e~�"֦Ƭs�����<D�� �XPD�=H����$
,d|���"O�����ӆ�f�CRS^y��"O�\��_�9 �E��a�\8b�2%"O��c��"J�2� `�!FH�6"O��b �����%�KL���"O���'C�b�d�ɒbȒf�I��"OFPQG
X�n��٘�&��7d�P�2"O�%�Dg�1
�Ѕ��E���ء"O(�)��� %��q��;O��鰢"O�U�LܵaB(�b�(dӨ!��"O��A�݈Sq�H��`�5N����b"O�a�P�+�<���D�$(�f"OhQ�ƯU#6��EW���=�-{!"O�1�&&�#k��a���`���	�"O�h�����h뒠_1B��Th�"O�\1$�X(W��e���"^����"O�]��,�4:�N�aҁ��5q�\x2"O���D��l#����Lh��k"Oȱ�3KG�\�,f��/G�=` "O z�+ܦ>O��1�B<H*bUs�"O��!e��0��!��?�T�h$"O����2{��a���C6m1C"O��ĭK� ��p�a�
�I�n!��"O����7C���q�2(�Dx��"O:U�t���{͈���\�?l��"O�@W�D*@s�ىW�$=/&��"O~�9�կ[8�L襏.+0H+S"O����@�?o@-��c�5����"Ov騴 5���f�sp@Ȁ"O&}@�C֘y�&��E�b�T��"O�% �E�:�fd�s>i�0䳴"OB�(e�ڦp� �b͇b����"O^l0%��2"�np+�&:s� �"O6��']M�2�޶MY:�"O�ty�)�1o�8������-P��3"O�H�c�X��81���}4T):�"O�����	BsfE"`[d*�e��"OZ+��U?��T�dK��Ћ4"O�Y
�a߰���D�{����"O�Ŭ�z����@��_�&�9�"O ����6����F&Z�֬=�C"OA�diU�[��\R7�I���|�""O��s��%к�Y��#q<�;P"O��9t��9����NПr��Bp"O~��1��R�psĊ�Jo���&"O�`��F�He֙�p���yjD%�"O�E��!6��i7BR�uc�5��"O��*��� ~�B���]��,��y��L�5��˂%B;{8m��F���y��Ō#�^�S��̓`����+��yrE�t���d"�l�(c�K��y��)��rvșe�n�HЯ�2�y�Rm����D��Uar0s4���y�`��
 L�8�lPRJ��Cb@��y�d�/�luxE��-?����-�:�y�CX�TT�	�a��4u�̸���y�%Z�~��g�.�Bm�4ʞ�yR�L�-����G��r�@0�y�%50Y�D%vx�`B��y�6�"���������d�3�yROS.o^}��oF�W48hr��=�y2G��&�R�fM"
u��VH"�y"�ǕE�Bx9s��1��A�ԫ��y�C�<�e[t�V�t��-�����y
� �Iy$�J�)t`�R�z4��"O�(�#���b�����npsP"OF��(l�f-q�� )��	��Iɟ��'O*,f�V�'E�Իia^����)�<E:���PŢ��O������O��$�O\���G@���Gh��*�Z}�V��!UЬ���/Q���I����p����T���Y1Q��F��6k�0hH҃��`�: ����YE���5^*�d��%� h�!QdѣmF�}���? �i�F�OPP@�C��{�j���4E[8x�K����	1zW2�Z����ʮ��Bb��t!��dG����� ����z��wE6���'P�R�j�z���O��'8��=K���M+��ӓoh`B6�;x�*��2���8]S�5�C�Ҷr`��N��U��Cv�� <y���C�-]��Qu��3i� ���K~}�B2�v�ʄ�B�:��3Z�+����e��'g=p���Ei�䠲6�Zd>P�'-pH���m���h�p�8zI?��+h��!A��Ǫ<z��e�<}��'1R�'��D��*�"��E+I^\	����`ݴ�?g�i�Ҵ�PQ���/<�R�8Y2L�u��D�O��dI[���R��O����O���x��û}�vh��#!}��Q��$y��k��>!U�-J�0������Ⱬ\�4�8�'�P�q $�)3F
�a`/^Z&�����>@��B�������B[�ħ{2�@)I*k��S�x��$0WL%~Q��إ� �z5>��޴�?��J�?Aa�&�Y�P�IЦE2��O�\���D�F;aL��h�K���F{��I#pg�,���?S4�ȖgT?$����æ�B�4����i�<9�aB�y�V���|��r�O9���Y�я�?����?��s���O����O����0,�����z�L�dv�������<t����M�o4�l*Ղi�Q�$�u�=�d�����/C�=C��O�X��#�L֙��21�ֻ=U(B��?��90�}�oE+�M�C#լ,����Wh�9��H9��<lV7ME����by�'�O�D`�t�n0!(��� �Bo 0�C�I:z��A:�22����"FM6^p��'��ӥ�m�l�z�H�s�����O�7�кsVJ�y�MޠA��-��E��'���	-n}�I��������[:���E�<u���⒂Ƥ��	B��<H�@q$��_���oŰӌʷ�9�]�N����w���ό(:�����F5��}�w�]����L�2�n����K4�O |��'$T7͙n����v`8�!�"�Vl$�P�lϠ'�
���ϟ��?E���i�R�x4�T:8j@0�MT8W x����6ţb�U����?b����=-�d�*�\�������M+��?�*�x��r��O:7m�.N.iHE��F�@�X��[�v��m�ɂe#�Io"�t7�[�_���c)�~9�)��ם b5�$]�s�l�K�� 3�j�p��U�gIқw���$��<�F�^w��aä����Y�=���j�%;�ebTG��D�P�2`s���l��xG�)[��,H��*K�S��t�S����ޟH�?Y�}R ��O� TC�u�6M��X#��O��m�)�MkJ>�Xw#v|��Ԁu�܁�wc�.4�X,�2B�O��O<���,J7 H  ��   >    �  �  �+  e7  �A  L  U  0a  �j  �p  Jw  �}  ܃  �  b�  ��  �  (�  g�  ��   �  D�  ��  ��  !�  ��  l�  C�  ��  K�  ��  ` � � �   ^& �&  Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�� |d��"O
`�(�;���8���-0��1%"Oj4��ND^[��"3/9�0|H�"OB���H��*�ʞRy=a"O�味V�!X��!&F�:J�$���"O,��a
���C�Ą�M�"O,$3%o�-���p���+Ն�:1"O��ݢ1����`���y14]2��i�<�6��{_���c�H�`�fX�$Kn�<��A̼VI�xR[�)�Ć�pඤ�ȓA5��('nߡ4�� �)˩%� ���,��r�؊b#`T�eT09���ȓ!�b��g��}�8�F��-? �ȓ
K|m�ș�VṔ���2�%�ȓ"R�X�j�4JN�1�˘X�i����̹	_�jZ��1!g��zܶ��ȓgil,*�J�
j�Ne��i�J%b���f	�(U��:���G��$Y^م�~r�� S�%T"���k\�jx�ȓ|4�1�îJb��@ӵ�ݩn�V��/[`�"�v4�R�!ʎ<��M�ȓ`:��z�ؚh�J�Z��$HY:	��H��p�m�C1��!��B:��0��EnjZA V;9����J[
2���	��4'J�EA�IVW&��~�(aZ��ӹ�>� o�Y�|�ȓ�f�A�
Ο7�H��M�$�����mޠP����/���ANXo*�ȓTv�����{ ��-7�*h��I��sB�8�8���3������X?4`�v�)���ɑ��]zR�d?��FJ���g䙇f��1��]$F{��d�P�Ӥh,�����$f�Z����&��F��LG�$(��A�B�I�JO"���)e�D��|�A!��\�$e�33��"@��1OeD�Jǣ߂�y�@)>t��@e�3V8L������?�g�|�I��"~�SF��>^56�S,Sۨ�j��џ�p?A�O��0R��)q�B�J ���6p��"O8�S�g�c�<5hd�ԡf@~!A�I;z��O6ʧvԎ1X�R�J�"X2�C]�[�݅�(�0À��
a�a(F�k� qE{�IC!����	� h�$=��(�w�*G켜�"OI3�l�iGv(����Kt�8V�'��v�|d��`����:\�����y�`�G�xA����
���\��'9E�����B�c�f��#i�vP��CC�/Z!��C���R1/^�9逘��H�S�Q�0 ��' �Q�L�%�P��fُ3��|�'�0	`�M	�虡V*������'���B"�6A�f}��B_���@��'�vaJB�@#?@��ZB�J(X(i#�'��p1Y-B��0P�,��M����'��x�!�S����H�J��Й�'��Jw��2t[�iC<��Y{�ON�� �4�������jg�����'�qO�@�1b�,B�h��!��eRJ�
Ik�<1�Bǟ��E��B�c��9�QA̓ N�<�|�ߒj�����΄={W�A���D�<)�焨X�a`t�ߤjn�����Zd�<�Q�ǓRüQ����"(�.Kb�SZ�<Av�G2m�а��c
�Ki��rec�U�<)4���p᠁g��t�쌂r��L�<� ��"��7����R�Ls2"Or0��*
���e�r
tڥ�	^���i�j��@����b�^�2%o�~�!�$�/_r��b�]�F��!��-��nw!�D��T%x���Ǚ���9�f],W[!�B�m��8�m�&(��P����.CG!�D��z��!��5 �R�	��|,�{b��5����Pc�97"&D+!�T�:�\Y���|A��#1���G�'��Ih���)ޭ-y���ʐ�'�tD �I��!�$��f���W��q̦�sBhE�i!�d[=A��1vh�3��B�J�!�d�^�ԀC ��N��C�%:B����>if�=�ЧǕ�t�t�
�σXX��Ot=4m�?zcH�`G�ט��H;%"Op8�Ё�;0�D�ce����Q��$��|6D���S�5�z���㓾i���Ջͣ}uB�	�p�&E2���$8���/˖�ģ=9����a��M�1lua�O>{����`٬�B1��q���1w+ �whh���ʰ?��S�E�m�'��09�E�g�b��4��ж���h5)��O3IЅ�a�*���.��Y��Pu�ب2e��Gz"�� G��⌄ &�iT�PB��5,��x��'A
l���H$As��2$��SR��k
�'���K��O%�mI�C�Qj8Ѻ	�'j��(��xV��3�.D�C
nx��'�R��k��pI>�� ��nF��'茘�嘷;���J��YWЁ	�'>@�є�@:�|5K�Wb�-�'�6�#LIS��4W)Cϊ��
�''h ��GY5E�5��!!G�� s��䪟�F����Wju��-W
8���:Tkʚ��=Q�{R�
�*��`]�<�}K�J<��l��m�Z�H�'
n����,H#X��#��"�y�#VO���O���a�+9_�Ѩ�`�,Ltt1�'Wđ(!��<6IX���(���bI<����O���剞r�Q���K;�qY�II�l��D��d[��#��PQl�
��&#D�L&��V��t{g�K:���*?|O6b��@����d��a�4n����J7D��96d:�,%�'��>�4y2Q��'�)�������kj4��#��E:D�<p�^�T1P��t������#D�8v�V9F�f�Yf��#�.����;D���d��R�.�ri�3"��>�t!�<�I���ɴ_R�`1������5�c��B�	-K�Zhj��Y�r㘭�1�ތ81�6m�C~��'T4)���R�kڢ����&n�ek�'�~92Cf^)9�pPJ�FQ�iN����'�qO�F��O�t�V�5�ja�U�N�J����yӄ��ç&�@D� "ľZZ0
piU64�4Γ�?���'���1^�x:���j�5f��4[��1,O��� N�3�1F��b����d>�S�i/��, ���� �KB �J����?�(Т4� 1�5&ڧ�ҭ�g&D��ط&NC]\4ۤ�ҁ��ȃ��%D��)�IНKeFI��mQ.n��̚�-"D���T�#w�^=8 kYQ��"D� ����FI"aH�hF� R �U#3D�� ��^-"5���c�x�P���$<O#<!�"�5�py�Эח~�N����Ll�<B��9GR���IB�&�PX�0j]_~��'�S�O}��h�G�#!�TA٘�8
��� �Y�c�
�#�P҇��4 ��h���?�D,�3�x��!��}�5w�/���':�U��O�3N��p�7|:a�v�Hp�<yqkU�:vD�vMJ�o	飆E�i8��o�m��V(`� ��pB�I�/$|�ȓ�Y�"�L�Nߊ,zB�ҫT�ѦO2�=�:5)��H��Ao�'1{�T��(Mf�<��O����"ΟD��q��S!ıO��~b��D��`#�܈��y�<�ڔ+o!�$C�Q�<]�׋ɜJ���A�k�Dj��D{��D�%yD4��V�ݶ%"����6�y��Ǖ�
]	u�����$cc�T#�y"KF��!9��S�!֞�����cH<�ٴV�ebe�#�x��B���o��{�'z^�t�ŞUO"�p0�A�9��i�˓L�Z�l �W�
R|����>��G!#D�ha ��*�t�y��(jS�\�f�;�	!�HO1�$�$HėTe�R�=s!ᒠ�'��'!
 �TD��[�H
�Ɏ���4�ɹ�p<�bH�
2Ўhr�#�e0�h:%�k�<f���X�鉱$�\���.�d�<�F�����X����S���	�f�'y��w�']�Ap�inRt�R�ͬ/D��'�T����֋>���pB�Gy"�j�4�M��'�h��'��)��i�������$����	��eR�'U�ԛ��ƈ*t	s$N:~9:���'H$�;�Aњl����"I}�
���}�+�Sⓞ	�ؘ[�b��m9�0����B�I�y�p��SÏr1�xZ�kWee�B䉦:c��;���W�v��(� ��B�	�a�%��"�n��
�N�HB��&�Y{6����jAd���TB�0vP�!�ǜ�]�h-�
ܨ�0D���Wa�|0D	�a�<�ؕCC/D���(݁v9���W����� �/#D��Æ��A�R�z%A� ��ҋ<D�x��+�U�����O��kT\�S�:D��*�,�f�<lr��>��æ�7D��,���H�A"R�?Q�� ��*D��H0��g��lh#BQ�i�~��&D��*bN<!ene	7l�dSl��V�$D�4������!�?�Vy�	=D���͑yI"dQ0(��[L�;e.D��`d7A"�S��M�h�(��� D���!��!&�~̀#� 9��ٳ�L>D��b�'*U�؀�RދN�D �J>D�|87%H�K2T8T
<A�ڲ�<D�8�ԇP�	��%�텻D���7�;D�̀`�2�RoB:$�zL��O;D���Ǘ�]x�Y��M�X\v�y5B;D�t���4j��:�F;�nl��.D�, �/�/���C�K��`�.D�p�����	�:�����F9;�l,D�@ʰ�Y�:7Ph⮛�S#��1.*D�`���*U)��S�l�=b)�(H�''D�Ȩ��Ǘz6H�
#+Qג�Z��$D�D��B��=ê*{�@���!D���"@�.�d����>)rJd��`?D�x;pn0�㇛`��ydn)D�\
4LI�/�.�� �F#t���C):D�D(@n� ��J6%��{6�"D�pz� �z<<���63Yl��i;D��!�@�7�A۷�~�<��3T�<P�l�T�\J��Q�v�����"O� �}�ӂGf���"�!�4g�Px�3"OEq�Ш�zPR3��;�v�˵"O�\IW�6A�eF�@4z""O�!�e�\�q�\uPPFH�]t��g"OV8Qs�����[����}m>$b��'U��'d�'���'Cr�'���'�ĲWo�0u��Ǹ|�V�'P��'o�'���'�r�'Sr�'f��:��C�K�	�Iڟ-R����'��'B�'�2�'\��'�b�'r����;���zA  >�>%:�',��'qb�'��'���'�R�'b�ia*֨"�D(Q�#��R9ґ�'�2�'1��'���'j��'���'6&���Jʴ��������r�'�'?"�'�2�'��'��'vrԙő8X�b�XA!cyDݣ�'F�'e"�'���'���'���'<�] ��SuQ����18ov5�T�'���'b�'���'ir�'�2�'֔0�{#�\�1���\�SKX�����������	ȟ�����`��՟H�BnSb��t��+\ (�����J������� �	ן0��ן �	֟<�I柘� �Z<��q�6Ɂ�?�ޅ��&ɟ��I؟��	ɟ����	Ο���˟��g/<��	'ctkF#՟��	ڟL�	��L��ɟ���ǟ\��ן��@蚨q>}ƭ_n�Ltʅ��ğt��؟(�	�T�	�������M����?��.���9��ǐQ����a*ݙb��IƟ������TӦ�c4��� ����W�Z�����0FM�
����4��D�O�@�CG�G�@���c��H�On�ė�u��6M9?ٙOS�I!���n��)�K� .ePa"K���'!rR��F��7����Bi��xh�,3�쀰hX6m�6?V1O@�?�h����BҨ@ۘ�hm�8h��u��l���lZ��ϓ���S�&F6�i��*���"7�y�o��=�B��Տ{���G�+_�����'��Q��T���5 P$H<X�'~�p���M+a��n̓T��X��j�0L��p��mW&@�N�@�RƸ>���?9�'��	�AU�}3�!˳
/
�ёJW)����?��)
*T��|ѫ�OV����,�e��A��RPtUu�\�W*��*OH��?E��'y<l�t��!lx�P�$_���'�7-�h�	'�M��Os�lk�ۡ\8��� g�rlT��'*��'e�&V���F���ͧT���3)�7�ī1k<C�,Xwv4'����Ϙ'�p�2" ���.3�f@�0���#�Ov�nږe�\�	��8��|�'GӔ��rl��'�E��fT�?z��Z�_��3�4Kj��'/��i?_`����HXf�hl�$��
���/C��q*�X��a��R7U�2��p��wy��YH�ZQ`�H�u���@�@���'���'��&��7��	�M�gA�!�2�f��D�6�F&�T(�I�?)�iY�'�"H�>����y��i����acf��M	.��ͩ�G�S�v9Ȓ<O��ٜWm�-R��)`�������Hd��c
����a��y͓�?���?��?�)O��ȟLC�-U40�9�
	 =���#G�%����؟0�ڴy�J�(���?9Q�iI�'}�\�ըݫ���A�$��j@x���'*�ئ5��4������B����?��ͯ~Y�ر�&�P�l�"\\�`����O6)IO>�/O��$�O��D�O�]s��)-H��A�%^�;ȸH�fNx�a)uk�<i!�i\.�	���y��'l��w˼�Af�L4I ��♒# ���'�"A�>�i����,�4� �I��c	��E+:���6!�l:�,闠Ϳ+���ӡ��<q��2���������Y�W��B���H��ӽk�d����?y.O:�4�,h@�m�K�@�(���$�Isʝ��Í��lu��C��'�B��t�'>�v�p�O~�Đm}b
t�X�DΝ� �y(���`Ό@p�!ϦE{ݴtL,Ȗ ��<a�v�r ������9s(O�(4�ux�g����e)EƉn�<qߓvr����h� n0�!7��D� �ihM�2�'�R�'���oz�Ec���P��ՈXxj ��4�_��Mc��i�hO1��٘�땦9T�$(j�JRN��,��ܩP��0G��d԰$�V|��e��OR��?1��!������b0Y��aX�}v�C���?!3�L��?�-Op�n�:� E����	(�Z��7�G-!���E��hh��	^y��'�h���Vo�OnO�Cg���4 ��#\�AH"���3O��
<$R^d�£>�~��
�E�O�P��I͢$�3%�( � laT�Y�����	�ȳ���~�j1�^m8�`��oB��LW'&��'��7�;�i�}㲬˼6��p��(t���E������Ǧ��ڴN
���e}~�F
=�n���.�� '�$.�e��ն:2͢d�|"Q���Ο��	֟��Iß��F/սpv (��A�vpt��Cky2lsӒ����bu^���O��P�D�V���O�؊�����!��6όI�+m} o�he��D�i>i�S�?!s6�<t:~t! �� ;���@7D���\�J�REy]5�Xp��K\�'���W�:�,gi��P�	�*7(��$˦A��)ڟ�;�ǟ_ �p���$!�xP������ܴ��'|�8C��oq����)2}B��1�(cvB�y@�
o���Cܼ��I ���O4f'?��=� Zq����v�����(u�T<�5O����O����O���O䒟���'H�/4�*��YW���2	�DP� �,�O���֦�`@�����M������4�MȑK�sV��2pᜩj�^�&� ��4E���O�����׹�yr�'-pM�Ў��
7
9!7����x�Ӧ���&�. �	rJ�'���ҟ<�Iԟ���#$��L�b�9%l=)�T����^�3�M�'��6-���9O
�d�������6.��f,��*���OT �'0�6�_̟�'����?h@��Fъ���fbj���V�ޘe@V�	�u2�'?�4��3�S@ׅ X�3eL"P���7���w�D3��?doP���H�c�`���ʑ&���6�+n��DH��Eဝ ��(J4���
b�2���˰W�tԋb�-F��8����+.�X��1ϊ�0�a��&U���&��b�Vm����:M1��`#*b]�Y�'���"�sTB�X-��$��N��p"�� yY<]!�%4^%��@
P7�A�w-9xv����ͮ_0�0�4�?hT�2��E3�ZE��|m61
�G��	�t�$�4kZ�CVEO1\����cĹLQX�V@�-NQ���?A���?�K>I��?��Ƣ��1��mH�q���W�v�#���?��?Y��?�-�8I!����d&��^LtUie
 -��'����M�-O�$$���O �d�_��Ix:�XP���6:�@ ��*VM���?��ӆ7��<	��_���	�O~�!�@�F�����2=��j�CW����	\���I�X ���S���&��M��+G0K���"�����'�rY����)��i�OJ����<j�FS�����&/��4膤��	��ɏWZPx�?��O����
�]
� E �?ST��޴��d� (5Z�n矬�I˟<�S9�����s��~X��0��!�~�x"�i���'�@�u��,�3�h�3F�Ѡº�K�;Xf7�фY����Oz���O��I�<���?AG��*"�� � HF;?ejMyU��;Ǜ�J��l�O>	��z�x��a�3�~��Ӣn)l�:ݴ�?Y���?���������O����Oz�	�![�mC�g\�̣WΊ�#"X6-0��oRT�$>��I��D�	�i3��w���T��G�+3���4�?��i������O��$�OV�OkL^?Q���2I�<=Ҍxԅ�'��I�b�H��؟���cyb�E#n<���D����5ndC`��>�(Oh��0���Oj���wQpuj�
�������4.9�a��7���O��$�O��-w�(�1�Ѕ�D(��	�nU�6�A� ��� E�i���ן�$�H��ן�i$`�8 DE��|B�c7���
��t�%���d�O�d�O�ʓKK�EReQ?��ɱ|����)�L_�̨�J�-%���޴�?aJ>��?�`
Q���'�b�"kT1s��F�D�J�4�?�����d�c��	�Ou�'�T!��:$U���&]�^��%cE1ߺO��d�O���t�#�	w��fֿ8=ji���0�\�����ɖ'+f�8�G`�x���Oh����dԧ5���@�������b���M��?�Bm���'pq�j�ر�rʱ��@_�<>-s�ioxQ#@�'���'��OG�	ޟ<�����X�_�g��4s �'F�x���4)Il�Gx����OT��R@�<jOl�	�i�K �Bč�ߦq��͟<�	�9ϰ��K<ͧ�?���.�{�`_ԩ�$�ԲdK(=�1�i���'��o��@꧝��O`��:�>�z�K�}y"��Ѱ�Ëp��d����S���Z�A�>�*��4O�t��K�cϲ=�^��¥�� ���?����?1.OB�!P���a����!�;=��"@e߬!1��'����'���'�����?-&=1�'�F�j��c�P-_e�|��'K��ߟ����q��kľLj��ڰV�%r��Ȱb����	ԟ��?���?�'�|TmZ�j(N]��E�U! ,�2���h!�O����<I�D��)�v��)T��cs�L3!�np���	�5��Po�@��?����C6��D�I�8̱Ձ�eL��:���'�.7�O^���<9���w�O�2��5�|�.� �JP�(GL
�oZBy�'��-K*X&��t��5fBP��9´�)X�.���A�����O�d�7��Ob�D�O>�����Ӻ��06�RP#��K)ǜ9�iPϦ��	ʟ�r��X�x\�b�b?�p-��/����d�ҬH��d�d]+�Ҧ���$���?�XJ<��CB*i`H%���NI����hAǦm¥"C�p��ٟ(���?��Of�S54\�� ��g�Ќ2.����۴�?���?�Rؾ��?u�O����5w�����}�4`[��~̓`������O���>�T���N#)�az�m�9	m��/��Y�/O����'�TM��H�*�F��F+�x��c� �>�ر%��=�'��'Q��c���_���D�8.f�\���@��Љ�M<����?	M>�,O,!�L�$x#,�K���
��9P0��}�8�d'���O���?�q��1����`�<!��ωNwY'lK7�M����?1���'g���("��Rش&��SP��/��$��b�9A�q�'�B�'��_����#�ħG�T�"�C:c� �����;�t �a�i�B�'p�̟��"��t�IW��ҟZ�N�8�T�m%��˔;�v�'t�]�$ImO�ħ�?i��Sa���� ���-$�b��Fڦٕ'2�'=T��'G�S���S��*��N��0�ܚ@�-&�ػڴ��d�>�����O����O����<�{�? ������lJ���).K��৵i��'o!7��瘧�O@"�	$c�ς���a��OX�޴��\:�i��'F��O���I�F 
QA`�����6���>��)o��+��������	۟�:�RT��23�ˋh4IyG͕K��E�E�i[��'��A̧*M.7M�O^���O����O�B�7��!#A�>@������Wޛf�'&2�'㐄���)�O��D�O�<�"Ƃ{����E�%��ٸfM����I0��@�Ot��?,Ov�����bAɅNTR�{���=:�50Y�p��"w����ٟ��	�����]y��џE��aFͰp��E X.!���(��>a/O��ĵ<i���?)��V�Vk�((61q��*7	v$1�l��<����?���?�����D$;M�(�';g�݋��� <�D6H�#:�}ouyb�'��I��d��������~2'�2"P*���#NT�AĜئ}�	�8��؟��'y�u����~z�/�|�V��'�6a���8X��r�i�2R����֟����xb��zqB��J��5+L�F�!�B�j���$�Od˓��xV?��	�t��1����A>m� ��M� EMH���O��D�O��C.>"��?��?�9"� M�+��+^�8c�`�2�M�-O�=��&�ۦ1���$���?%b�O�.S++4h�bCK�sP��3�Ɋa��v�'X��Be?9����<�S_�n��G�	�4b#�P-@�7͍���m����������� ��D�<t+V�x�>h8��@ҥ��z"N8E�i�q��O����O�r
:S�n�G쐸+I�Pb�Q����'���'Z,�(�c�>!.Ov�ĥ�����Q�V�H���,4L��%j�
�O���=O������ڟ pq+_}"����<P�P���M����LS0Z� �'M�Q��i�з�
cˠ9a��
$�Y9'�>'�J�<9)O�d�O��Ĥ<�r�Y>�pg�3(Ƚ��O@�e�FP�`�'�R\�d�	ݟ��ɸ;r4�#P!�>��a��Fңf��%i4br����֟��	ޟH�INy�]3j�瓩*TJ�Ac�!� 1�d$o$D6�<I������Oj��O���c=O���$I;r�
���ēa��\���Ǧ%�	ϟ���џ��'��yJb'�~:��{u����vnU�s�
���¦q�IgyR�'���'�RX��O��	�P�������>Ty!䓀g(6�O��$�<�ըR)*�S�����?�"XI:��Y�O�
'��1f�R	=H��?q���?��(�}��<��O2Q넁�<C�Ĕ�g�ɻs��ݴ����]J8�oZڟt�������������1�J8<, x�o�5ӌPh��?9��[C�͓��9O��>y����d�2%߷�-he�~Ӓ���L¦��	���I�?iX�O��R���i��2)=X5Z!.�#a��
��i��MK�'(�'N�0�D
��Z6e	'
��(B�@�b<��l���I֟$�.��d�<A���~���%R4����d�)�0&�Mk��?��K �S�T�'���'E�Ԑ��,���d��� ��%eӜ���?�`A'�$�	ퟀ&�֘�uF�z�� �kG�`�>��_�ܩ��y��'CR�'tr\����eܧ��. �K�Ɣ�K��܀g���ē�?�����?���[����4���\�T1��N*ab\��E�<�-O:���O��ķ<���$i�)Y5L~^l�A�_tV eq���J��'��|B�'�B}���L~�ȁ��&$������A�1]��J�^�4���l�	RyB�\�\��(0�V	���F=�$	�'d�ԩG+U�����l�	꟠�I�\�z��S�X���l�@E������Z�&����'��X���Ũ�9�ħ�?A����8��Òǌ���9/N�Ոp�x"�'_�Ď0�y�|���$�u���{,N%�N�
6�`��i��ɭb<R�ٴ_����������)��-��j@&h���q��ߞ|m�6�'��oǭ�y�|�IɁ7Lv�1TN͋C��L���ɛ�P7R�7��On���O�IUy�˟�a@�.���Yג�r@�M+ck+�?�J>E���'8 8f�-7����և
�Y#��r�
���O��$
L��]&� �	ܟ ��{p5���ʤ���t�P(n�n�I�Ĝ�)���?!��\M��BP�-_����/��a�0�i�b&o�O�d�O��Ok,T4G�V9 D$B���*�@�3k���$]�$�$�����	iy"��#�L'[3*g���$� 4e�r��$��Oz��/���Ox���	����a�>�(!�l�9Gv��,OoR_���I۟��	}yrM09�f�SsBDHǁBn�A���>k� 듍?a�����?i��I���J��!Լs��@2=�)ӣW�&�	�W� �	ʟ �	py���B�6��?y�&YT

������{�P1�-��;{���'���ȟ��	���EKd���	]?a���(6Sv�@q�U�\�Uk0��ئ��	ş��'s�d{��~2���?��'R��l  'C��˅�7��TI7U��	�ɼC�����D�?���܆^�JQ�V�v�ج�Gg��x/n�3�ik�'���O���Ӻ#�#͘A�� �PC��!lh�y�"Ǧ���۟�sd�d��᨟�$/�  �*�A% \ ��*s|�����Ӑ� �J���u��ݟ��	�?)�O�ʓV&��R)����c(�H��u��i�H��'aY�t�jRɍ��XXp�EmQҍc�O4@�Z$[�넂�t$H5#3�*����'�N��jKZ��� :��&�)VT���#���!�LE�D�'� �t�4[�u���V%ֱ�Ǉ�!
ش��\2eu�q	��a@@�B��� c��3��J��F��+��aq�W�K���F�ff��Z�FZ� �$�*��A>)PW��S@܁둮� s�xAE�zN�tD_�!���# S�*�哆]����a����x���?I��?���$�?I����4<('����mU+`�"(��G���h*�6g�qz��:u�T���<e��,���/������h"�[� ^�4��!B�Ɂ0+`�U�f�'.�\S��?yC	]5;x\��a��WU�d#�KT$�?i�r�s��)��:Cv�z�G�%l��8��<D����)
c����� .�}Xԣ{�|˩O��6-���[�p��M�� h285�U�V:nL��B\�s@�i�6�'��'�`y����~M����Z�ZB(�T>ݐ@� �s#��@��Y;9�^���@/ʓUbx飃ċ@HIIF�Ԡ��'�yZ�j�D�T(S#�^"r\t�Ey�%G�?�����OG<��A��NG6�ەd 5�F@ʝ'7��� p����;��T�#��	�0>A�x�&��fw��%�w;Thcc�W��yoO�&X"7M�OR�D�|��8�?���?QCXv�D�ţ�,eZŸ��Zv�>���f*g[*�c>�d�>^Oz��2�ɨ<Mp���@�6�F�����$�D�R�K�I��X�)��|�����xMRD�Fܗ)�n�1������������'����1�K�k��It�S�@�ȓpV�a��!]!��QQ߀ x�����P����'�`�ǚ�A:$X;bc��r�C�'g�$��%YֱsA�'���'ZRci��I� ;M��Lؐ�
s+L�i���̅+�?Iv�0قx��$�9_���3�z }(!�u�j��a�/�}�D�'A��dl[')�8Ћ��MF{bIT�0��y�HM�E���K��~ �;�?��hO�F�b�`D�4�8U�"��"i���ȓ�XhcgH���I���9d���G�i>���Dyr'����JT�H��|���F?9_8��ꁴ|��'��'0Xq���'���'^���1�ռH��q�g�(d��e����4ΌI�Wm$]j�9{ד@ 0�:�I�^]�7�Fg����Ï�},�ы�KھJ������mt��'�RY�6L�3�b����I�W��c�5�d�O�?��+�iV�V_]H�g�Ip�ԋXH�!�DS�U�0��0:�IBWHXt���̦��4��d%!l��nϟ��	b��+^<��P���г}�"q*s��2�h��!�'P�'7����Ƣ:��O��=F�v�óŎ3"9�\��ײmp�<����$F��z��iȕ{V�e���Qr�:+a뎭u�Q��z���O��}� ?���[BɅ�@ D��"�s�<C�.�y����+W�Ns�H<�Kա
��Rrƀ&~�J����<��M!&���'��X>���Rß�����"��!z�h�����!�	��"������[�S���	@Ўɲ���B怆�b��ܘw�F#<E��!Ӓ���1y�DxӆO����B����?	�y���'��;���<S�l���nTE�	�'�H���Ӊq�y�����A�����H���t�'� Is�͂*�,��B�(�E�v�'l2Ђt\�9��'�r�'c�bm݉�i��c�F�^i�@��]8Ը�ee�$\lL�����/D����g 7o4���>�(O8���
 ̼�%O�(Ls���<i��	@JW�H��	�� ����K�'c����)X�X8a�s��$*5��'ƒ������=af�)2�� Q�7{�N�2�a�p�<���0G ��шY�.%�IZTA�㑞�SX�I��JY�ܴw��8�%���D���&�{�q��?���?Y&`���?q������Wj�Y��
:9� �O�Yx��RW�K/E��PE �q�0X!ց7O\`�Ey���E|Y�B�̖1���r�J�B���iF�)e�inC22��'�0S��Fy"ˡ�?���5W昪ebJ����Vl�2.U��ȓ"C��ZV�K�m��ȑ�P-g����k�|����!It`a��(Q�&�ϓV��|�&� "�.�'�?A/�m��NK/eSR��u��`����������O��$�X��]�dgР,X�" .K�'Bm�iV%�>y��I��:��Q�Io�'͒8���[�1�~]����)U�h9q�6Z��URG�Ȼd0&�	oӺ �\;+�c�'�T<Z���?)���kA�dit`�U�R�o�h�B���y��'A�}R���k�r����n�<�3'dΜ�0>��x��e|r�$�jg I�g��.�y�B%TO&7��O ���|�s�K6�?���?�2��	�F��! Ͳ!BLTZ�
S0&�-�������	R�	+����C>$bp�$�f���×i�������M6QZA�Wz��T�7P� �y��'1O?�� ęa�+Df�h��9��=�"O��ɓME�Z�Y9�$���'�ɋ�HO���O�HJv(��m���P#l������O��䆓0m4x����O��$�ON��ú��Ӽcr�"o�H-#���-���r(f?�GM�m�~|	� #LO2 0W��]J �8&��<1p���0�Ov,�n�(!5>]��^@���pG�n<�HQ)R�A�lt���v�����?�S�'�bW���f����������"p~��`4D�tXEÀ;'ڮ4�A��;"ǘ�^������|Z*Oƭ8Eh�ʦ���s��Ck��$��(�$����P��ڟ8��.X�����,�'�~H�b�]�s��	���T�{� }a�A
"Ugļ��.�n
�U�E��J��C�`	E{��R��'l|��ʗr<�(�d%��ke ���B2@��Y$+Mb�'㬕�
�G�P⑏@<u"���'��P��A���X)Q��o��M�
��hO�i�H��p;T�8����5OrI�>1�׭_S���'��Y>	&��2�6X��
��z����q���!�	矨�	�>��i0`l�	Ǻ���(H�X�ڟ4\���<^iε�%nЌ(#�<ʀ�	2;��\�O%N/$�&l�OR���OG���D�=/Y� ��}�P���4zC���=���D�JY^�q�7&7w�C��C�L��ƥ\:$�� S6΍�w�����FM� �ft���*��E������y"k�B�"��?)�X��֌�O����O�\JUn�=1�H� , +Bی���1e��mrpII"��S���-&��O%1�wa�g8\�$@0U�H�i֢�
%�d�u�͎/.΄��jI T�}�A�(����)$C�8'��v
A�S��Ys�m�A1�����M�EZ����ɻ<A�,U�h.�8ۥ��46�����T�<�Á��dțr獖>W�Gf�P�'6#=WT�L�.Ф_T�h7bD3j�޸���ʟ|�ɫa�~<��*�؟�������ɲ�u��'7�΃�7�=��Cǐr1��(���l�#6.�Xy�C;xF�Fԟў��Dk�d#-�]�\��*_�M0�Vh07|��Í�T0�E�g�'��dB�	x�H-�q�\�$N^���'�N�c�����u�\��r��@�G�ѫq�,!�k_�{��S"O��E�7�^��1
��w,�Q�dID�'��듸��̸@��oQ��X�P/�>U/h}x�!�0R@:��	���ß����۟4���x8�捤;hnq��iD�m��B?%�,���H�QJ�}��B��Oay�n�Ԁ�AJ�9V�p��L��~�u���Y�^P���L��z�򤃳f��yӜ�PA��x{L<���Dcxj0�����'#���0�'.�FP���j�q����!xEȻ�"O�+S<~n��c,��?��2=O9��g�=�'���B��aݙ������O� �a&�y��U v� Y>z���C�jr�'W��O}W\�1��ލ_�&�&CW8cG�(�'���p%�Kr@f��)v Fy2��3�$qE�G�{e�h����B~��S&]���A�ޜ���S�N�4<£<I�#�ǟ��I[��ӟ<�3��&&�xd@_%K����ҟ,�?E��'0P1(ㅋ"v�U�wʟ5�^)�,�'��q��˗\d���眱[���'����%F�����O��'|XV@����?��P@�� F���J�	��M�yVU�%a�Y��m1'��"yN��T���2��O�غfg��6�L-�Q�BN]r��b�9[�X�)Y�.��|��"
 >k`�e��|���ar�#Ьh疭 ��ͳl������69���˟(�����'QJe�� � z"���͆� բ�'	��'c�	be� �| r���0t;>-����X����]>h�J�2dǽV,x���B{��$�O�@���R�F���O��$�O |�O�r���T-ȁ����<&�ǆ�~b�ɟM���p���9Q���d�?Oy��W��g��+�)H�{�D�'���;R�P!j �p��	�n�B�k�#[�}vR�rU���'�X��V�'�^7��ʦ��<�����<	���Ҡӂ"����dZ4;�!�D��#�� F��/p��1���o��Dz�B_V?Q/O�q�u�����Ag
�NDQaa[�N����Q��?����?���$߀���?ٞON�I`��?I�мm]QC�C5�f��j�p8� ���<���:Y1P9�E	/l��"Ni8��Q��O��d�a7pݰ@�>AR��@��[��OV���O
��'I��37%$_Nv����;n,�ȓe�)�DIA�&C��@�
�}*��5k��oyB�T"qo�6��OZ�D�|V��8]�Zظ�튭X�6a�`� 27��;�?����?���@3� f��t�dH���=���^�?ɠ������U|@̐�g��2Q��B�R��N�ё�G,g ��a�|�ϕ%f/X��5 ��t�0�!���Q�';����?	��?+���" nL�O�:����?rX�|���O��"~�S�? 6�A��Z�8� 貄���Z�b����'�JOJ�H�,D�gtJ��
/E���╟�0t�O���DE�mW��ipH��SJ�i�\�!�]�[-lI��@�h�� �!��7S&m��hV�1t���F�.-�!�Ďwܦ�Z�E�%)�����,�!�<M2�8Y@ �`�*�nD%j�!��:�zA�`H.�<}
�.F4�!��@�-̢����ص?�pU2+K�!�d�	F⸸9�腺,�fJ���r�!��C��� ʗ�ڱA����bH�L�!��R�\��h0-�!�(,���ܴ#�!�D�?EʨMX�-FF�:i
�oU=S�!�d� /b�'�^9������x�!�DS�Po�t�Z�;��G��G}!�0f�`R� �$0�M;�㕕Dh!�D+`>=�!�G�5$��W�,�!�S�r% =Ht홷��	�f���R�!�$�o|��`ƪ��,>�)r6�Jjq!�d @�*t�%DZ�hUɱ�G�8p!�dL�L��4[@�Ȇgi��CI�*@Q!�$��MJ�A%p �H'�F+6B!��I&G<E+�.�"�αZ�H �!��3NN$@2&���ƴj2DW�,!�D�=|�h(��H��	ہH�/(!��)@P�AF��m+��&��n}!�dJ�d]�taN��o��-�W&�+Z!�D�7 �.@�� �0h�ʝQ�D;v�!�$£oj�����X�'d&%��͚�J{!�DK"W@��ȸYc�����т=�џ\uBD�ccf�c����IЖ�ӵ#7����R6b�p��"D:3z��ϓn
,d�8�B�1��ٛc���-�F����'����e	�Mz��*Ę�<�H�O�m��MG�`F����iT2;��M��InP2�&l�#5��e�	��Q7t��-S B�=PW�N~ M��	,P"�����}r�yk_-�r� !��.?���3�2Zv ��/SJ4hw���	vf� ����h� ؿ&`ʈ��j" o��Y'�_�b��z� �;,������ ���fE�0G� e8.�=K���E͂O�'"�8�!ӱ0)�X�� �*�|i��4W�t�2mT>���AN�;�&�=�$/̽���4�۶)#��Sn�H�Kl���ʍ�b���ӡJ69%
���� ��Nղ�+UH�v��Ez(�0A�l�p!���4�8a����  ���,W��K��3V��yr�@p��­�(�=��6L�
��� a\����	2}%X1��.Q�5p�DM�:��!��	2=�Xzf@E��9Ӈ�85�zP��O�SP�иs������O��xT�W�g��z���Plz=��k�aA���3OP�`�㑶�ēWYz�K�$����%�*[��s��"��� bm����l1j����H+lO�P
�S2h�����;���q���B7�CJ��I,��'`��s���p�*�ң�{���.�-�5���R	}�x�Cȉ�)a�Z��J�p<���ݱ1OhP���F�~\l�@��\~"!E���d�tl��{F�2xܚ��A,�4u�FH�@#&nFֵ�å)�O�ȋ9`Z\{��^�4�)q�@�#;��ՕW:�D�E�	�,��<����`��a���a���!��~ՙ��C{��
H�7OQ�V[p2a.\������)L0�C�a�W�2�4��f� 8��	%G=Әa�O=����� s ��c<MzG��2�P$5��R::�'�<LxC��_@��5��0zF�ip��N�.<��C�?3�c��&�����p<�5��,g2����H"xR2\0g"�I��ͱ���T�Q�d8��'�M�<6�4����2p�A`i��	R�g��5&���:��@K������*��Hs���N4�h��޼�����"����4���&�³��5Z��l����7y	L������ШH>91I��XT�	��,�,�@P��
�qOX!*Pd��<�¦�^�mha�b�|��э#��Icģ��tc0a�%���
���4�J>i�^�0�4�:nc�F Y�xsw"��"6%ʕ�,���a��7���(fk@���<-ٛEa ]� E�
Bh<z�Jq�U�Z0P��[JұO���e��&��{�Aۢ!��Q�+Μ=戩���0\���p��������\��A�Og�|�������?}����:��	��M�� ���r�ռA�����������'s��r��ڹF������V�d���#� R �%�'풼��̒h}�t9��!�S�^�:m�u�\���.[+!����D��ᩓ����%�	�'�B�e��K�B�7��A'Nښ.�.�S��[%$>xtj�����D.���ӭ��Ј�����Kf����~*+�dmJ�F�Z�ԩ�e%�S!b���CƆd�أ	�g&B�aCo�){t �g&W&����N����M�����d��+1�H���c��(O����;"<b����$Y*��q�ֵ	ӌ�!��d����Q�2i��$QA�����lH�yP��\uM��:FBԨr��A˂��'���әVj���q���e���;d,0�!�e��V�a3��Vy�I��=�?yskM�qi��Dl���)�����HC�
ý+lܣ�&�,U�Н[1)ţ����'�d����̪	�,"��ũU���`/O��On��7�����cS�J*]R��N9Z�@��b�N���ɢ��5%Nn��3����%_6EU�(�Q��`h�?u�0�Z�'Ŧv�1��.Kv�Q�R�X��dC۟��i�DR����J�`��y��% #�<�a@�a8*u
��I�R2&��0 ��O�iP�e��]	�샳p�F��(��MpkI��'nb��B(FW�*�V�-`����:��%�ƞ(Zې�pC�M����R�M"<�술��O[��rG�
53���V3� L���,�db�O��WG���Q�d�s �[|�{���,@�̀H~:�؄L�&̓��9& ,���2e�Q��F	���P�8�ؔ+�ʦO�J!x�3@����D"����7'��%aƪS�k�P rL�O�qr`R B䪴�@ A���Gv "@�O�Q��	9�܁�$m̧#.����	%y�В���0=��,+b�HiV�ّP�D�S���=x����E
F�%���ԋ��piFzKR7�H��J�I�슄ǂ�0n�3�5���<nR4
q�-y�/+FB�ʙ'�L���~Q~�����t$��W�� ��p��B�,��uKV�R�N�)�w9��v�
Hb-k�bU�,��ؑ�8�?� .آFmV���F�=���J~��J��y�G��R͊`� r��Vb�7���<H�xW��0/�I懭|2��<}��e�v8k���)6�`���g�hX*O��B�7L���.'��1����PV��@	�̓"X�Q�F*��3�c�'� ^�'o,"�'��{T^r>�Ơ1�k��M���;Wi��hCX�` e:<���ɘ3vȋ2�E*F�Ƣ>qAC<S��ԪӨ?�QK)R�O��%�PI!B�E�C_�z�)�$�-�r}B���0Ů1���&]�@���ɓ!��\a0�:���P��%�r�cw�Aڶ��'c*�{r��-[}0���'h�uA���
T���э3?X`I���`H�+O7m�B!���Y]1OR�0e�F�̌��c� �$����$�e�F�2���C����Z��p�P"  d�a�L�ƞ,�#7K�B2&�NH4X��	�i�0�"��Μd70��c.�U�@0�"�B���KrS�|fR9S��'#jX�ōR���)ч(I`>T���'ʄ�X�j��25�إ��Q��M� %Bn#>Y�b��25�ȅV(�P��E��߭��DG=LqJ��U�p��4H���	�~�lA�p!�!�t�i���?B6����ZG�0A"�t}�� X-��8��)RA�4HP��HO�5�c�p���^G������ą�Q2�b�VF8�$!�h�1��p0B�'�ZU�U���n�,��A.G��|`��''ʩ;�.��-�~��6	T d�h�p���#k8�f�G
(@TD.?�m��nK%EX}�R���B )	�2�qO�� o�%�?�&����~�$�]ֆ���+0�nl�ӊð~��=I�H��!���Ն[���4��L��kQ:�v�
t��[�����l1�`׊ ��I0V&��|����۟��&`t��bJ.lm�BM1vJ��4���rec�6*r��QFz��3�	�CC�,PT�c�X���۫):f�80L�<a�f ./����E
�� u!�S8�ԩA���%w4�P��1W1&�1E@�:t���D*%��c�\Pt�?M��pW���+ ^\D=j6l������)\=B��Mă&�F��0������9�����m^�qt�ȓ�'Z�_�B��.s���M��}Q:��B�O�=��/ם0�D|�W.Z�vL<��tI�&r��C�W�S�S&J�6��Ok�pԈj�Fe�K��D1�.��?����?��!*�Ѽ��W,, 8�N۵`~�tZ%�O}��0Z���J�T?���G������.3���F(˂-a��`d���p��'��	�j;�Ip$��l���9����_���I�T'b`��_) �\�ېKT5<��4Jq*��?v�řM9DT�O��)I?���'�ƑBHV�>�(�3f�
I,�H��d���#��!�����x9Ɛ�=�O���#酘N��c��t��z�� ;x�I�u��@�&�9��y��ƙL�t���d)KK.(���E!8n�� F�y�S���"�]Rm����Ǉ�B�IBO��~�m8�nQ�|�G|B�A~��ɉ4�8�̻
m�!�G�SGz�i�G�b|pq̓;�>�t��F���+��J��>�D
U.� ?������B/mP|�,O�U)�ÿ<�Ш@pa����zh�꫟ȉ�oI�\bm�5���_���ѥ┼H}��k�-֖c���A�8�Nʓ��>I���'��	zu�U\���crvb���^D�1��*�V�H��6�|��
u��yȂ�_�
TI��0,~,�R+O~�)T-U:B�`�;"���F�?N�\�R���4�Y!��˘�$��'?����dO�Q������ ~�ҥ���D��٢�X/c�>P��1O��I@�;�S���'js0��C��|Q<ܱ��	*�!`�I�^^F��=K����J
"V�9��m��<�<#>��催S��͋���)H)�cL��/T>�z�O��JEJ�g�d]�vI�	
\��	G�O$�s��Or��7ȉ�1�(T ��ܵ�(�"�88��G�'�k΂3
��SAS�>l	�J�&(�͹��Qy�$�x�Ѷ@-�l�v�ͼK��O�S�ZnL��	,�zTEB�ٍ�d�D�ث�->9Q�o�;St��
��F�W6�p"EX� �7�#� �j�{ak�!gRPe��«0�>��ɤ���!f�ԙP\��0��g���BD2�#2T�):��O�扫[�����D��	�dcPC�|� ��[��UD^,@��X�>��x��R ,�@���j`Gq�I�;�P蔪�/|\��ȕ
�1Jz�"<q�I��Z�vA��!E#x��h��i�6Tl9*I�KH�c��)v�cG��S ��*���ܨO�H�fi&p֊	�eW�'Oʩ#u �b@��0Vp4y�����zR� hȈ9�@睷x  ��M�:��>������x��y�b�XSԇ��x���k�j��&��{�@ߟf/f�h&�(B�Ri�Q�>GU�;�m��A;PxG��TK�J�D�j]��вIπ]�<���BӮZV0���"ځaBV�)�hQ�������B 
Qp���H5�-bJ��C�|��I����<K�&�c9�f��(�w$\�T��:�Ȁ��q�c7�IO�XM�f��=Ԃ�����]�(�ɤ-Ɯ��G%X�Y����R3IX"<)f!	)1���b�/ ��h�a��?�N��kȫp��� ���&?����;y�47�9�A�X�p�.��#X�1say��ȋ�Y�w��s��L*f0Ks�HQ����v�X O��b)�����s�	d�
a�:���D�~� �E�ۀP���`!��	��布h�?V�a	��(��">�3	��\������x�,��M��<�$U/��1���Q�	³�L����'�vEc" ߪs]$HAOū!����{¦F�_j�M��I�hθqDJ�k�je��NȄXt���1$�`��ɏ/P(TO�>ٶP��GT������
šu���e5_��zrAw�Nٙrl��,֠@ ���<.W�>qsᄽiG�iȎy��;D��E�!�,z��8�B��߰=�A�C9'ڈ����S�7��#�Kl�b�]8�"Bm52%�ɂX��Ĩ">�D�\)?ě�N0J�ޥ���0{� ��m����'w�l�#{A(�x�n�#WC�H<a$�\�(0@8@4�ZT�g�'L�eQf���]�f�=��@�YQ� ��T��$�F�A�o�$0�	0@��aI�`Z2(�Q���;[�9!w$�;�paY�Z��D�2�"�7�eZ����\Aӈ=������s�(r��dG}2��a>Ь#��;~"R��T�[�*�6})�-؄	�{"b÷2\�L:��>��=��f\��<��G&p興�X�x�-\Ș�G|BOT�l�Ti7M�g�2q��+QPd�SHB���O�9a��۽�����(ۿ�ę"�i�xC�f΄X!H����Ea!:����K#/��͛#	�'��R��"_d��c�-V���-O�}��b��76X�#F��6��U���>IC\?A��M�/+ĵ��ćc�E�B���|[%�M�e����Ɂ]��иa$͒dh�v��UJB䉡aX	��#Ma�RD�ܹ$tC�		&��A��P�D�Mq"�_[DC�9=�l�Q��d����ǃ�6�B�I=']�y���P�)��X+I�VB�	�1��L$A�6_z�A�խ�|��B�	�L��@v�>z��K���H0B�	�*�}�$ � kCXy�6!E�C�	@�i[E.��pIva�se�'7a�C䉚Z�>�
�H��+<D���ęh0,C䉾h�^\�DT8N����1�K^B�I�~+Ti
�Ӽ#x�u����j�&B�	*"fƸssA��=�e!f(�2b�C�	46Z1`�n�^����l\�T7�C�	����u��V3rl�Y~�C�IP�"�K̪x���B1��C�7S���Q�OԀw=���"�*r�B��8{�H�G��T�`S��B�${6ιx�ǂU��x�蔺L0JC�	�1�ʅ�+��REr�x��Q�"�C䉽L��aq+@�DЂ�D̔Tp�B�ɓD�(����d�pX�C�˰J�LB��5OD*4�JF��B@�v��0U	�B䉔Q����i�\6$�k�
I+� C�)� �@Kk��R��y5N�:7^j��"O�XgP�`+��K��Z�A5��#�"Ox��e㑸�� kg�K�4�u"O����O>JjLB������"OT�Ak�/G#��ɣh�u�Ҁi!"O�����A�[5��y�^�B`"OF�)1b�MaեR.�L�;U"O�A�Ć�,%�.7)�`�x�"O����@!n�i��sђ��"O�\��l�6W�-i�F�=� E��"OHI��NO 9/h��N��:��a "O�Mq�O�e�ޅ�čԦj�F���"O��`1`�f�q�0��_�����"O� R� W2!�K�cs\���"O�Ds7-��(���<ke�@��"O��2�eҧ7t�ɔ��&:.��*�"OR�����2l���U"F�|1��"O����3(~n�p��֖Q���q"O<(ӂ�A�Z ����r��q��"O4!�@�ԧ3�6(ц��W&B��"O�I��'�d|	�<z�pH4"O�A1n��A)��:R� �Y�"OZ�۷GA)a�&��fL8g&�d`"O, ����,FZ8�2�'$�`Y�"O�A�E���]G@�#��G�E�4��s"O �xwi\3%�1���>䆠�"OTZ�-�~>�� �D7� S"OΰR�IV�?5��P/��0����"Ol��4�[���{d.
���{�"O�]���L�Z���It��8e���@"O$��dƛB�X(�" 5�~9��"O�%�2��,�<+�/�����cg"O��R6iT�?�4�u��$$��i�"O�p�a�F�5� ��@���q�"Ojh��*�^���C<"���C"Ob���#�6DY�#dƝZL����'��� {��2`��2��)���%D�\AmߐW�С�V�԰Ni���1M#�-�S�n�Ҳ.� =����:(��Ʉȓs&ͪ��]�V �)�`8D�ȓh���A�HJa;R���D�� ��ȓ+�N8B���b��TB�|#͇�H�������FT����ŽU�|��>Ͷ�7�T���h�( 0	�0��d��-�"���r��/^d����,C} $�@Pç����Ɠ<28�r��ӗAbxd�l^%��+�'>��·!�.�ָ`�/V�"e�H��'�>�9 ��X�	�E�T�0�'.��A��0��5�)�غ��
�'-B�� ��;BJ2�zɶ}�*T�
�'h�x�eT�e��pЀ�*�ZA�'f�H3%G�G�� uJ�5T[����'>@8�SHS�l��
dCMUvލ��';��4�6d�lI5Μ�x�'kr�J��9����rgF�Z�ȵF;�S��?�A*k#�[éB�Aƽ`�om�<5��'By.�4�׷'�L� $ �q�<!6F���v5h�W(`�X��W��i��`�'����2�@#p4nI�l�:ʐ��'�
D��J�=e"`�-s��=�
�'�0�rWjτ[�bb`h�}r�'\ �yt*�		�vL�$*Ҷe�tm(�'��&�&���F���DPF����y
� ht�Q�B���Cm��@�"O�@4nW�G�pi���X�9�0�b�"Or%-�T^<d3E^,k�&�{2"Obt�viR&(�
4�ע�.z�d���"O@�9��جBC�ț��ʟ��̀"OԌ�0`
$#�P��aG�H���C"OH���(�䈉�,W����)0"OB9چ!�"k9*�a��Ge�$(�"OZ�IF@'��Y�$�a619F"Of�J��@:s��8s�A�0/u� �"O<x��dG�K�Z\t���s�3�"O� ��%O�Az*C'�Z�~�*��t�'��4�*͑i	�%��%B�� ?=�8d��)6��;�c	[��ɇ&�H<����e]�B�NV�`ZF�X��$/���H�@��2 ѵ|�̸S�
�ht�G{�'�� �a�@':Yb��0lώrba��'G���G�EfL���" a�@���'�Hx�D�$P�J�藨Q�@�	�'��D`T�*Mk�J$,?tJ�R	�'&ڐ��-����5�,�>���
�'[���b|���&H�8d���'(Ѕ��`R��#L�m \h�'��Ͱ�����L�� 
n��%��''00Rg�����wfKSJ�� �'#����hI" wT˃SP���'��Y�ΐ/~6(٢�"@-��b�'
l1���-9�p!E)M�0A6�+���)�T�G�6nꄪ�坷5�,�Hu���y⁗77e�L���	� � �A��ybM�F�\q�%��~��	8���?�y"���\ܺe�Ոn{��)�c6�y�
�?lG��H�γ�8�C��[��y��%�m��d�g� *��I2�y�,M*R�MҤ�){Rd��"�0�yR �"���H�D|/�܊Ǆ+�yMǜo���v�SnA��;�y���f_謠�K)IЁ�#C�y���1����+���3d����y�M�!�<��v����R�(A/�yBH»iB�����V�O��3�Η�y"�̖E �h����A;n��Hɠ��Oh�~�C6����O��kJ�-˶��^�<��	���#AAU�m�h�d�</�$8ش�M�L���F�<ɡkB���b�^�I�v�c���C�<���%l�>Q��Fйa�R�+@�<��.̕2�>� ���6�"I!���y�<��d��	�h��j��n}����Us�<1���0]Yz˖@ۆ<"���S��p�<�$�ױg��hx`���0j�I����n�<AS�&I'�<P%B%� x@D#�j�<1�A̦@�4%ف-��q���B��HL�<����+{�l���SO�D����F�<с-׼?�0�7�K�P]��"�MQ�ē���s�P`��ߐ\�Z��êH3�Ph��4D���cD��
�]��k�,��3D� ���ؖ �(H�JP�)y�Ł��2D��@��ɡ����
Ԅr6���g4D�8#��E3kz��Ӡ�Q4=��m�@m1D��z�+P�Ǥ�Q�E;r�i�`�1D���!D R �bvB���R�,D�D�3�ŐER0�cg���a;�"��(D�t���5(W�0��H�iJ���` &D�� ��t�<]�j��ł?3"0�"O0$r'��ξu�5D��l�*m�v"Oh��se�P'�Ԍ6��Z�y�<�p E�8� ��5 R���	Zx�<1��}�!ٓkP�J��!c���!�!�d\�t���,ɔ"=�P�6���!�� �`Ȱ�Pl�![P�tj�7w�!��?~壦I����(���gݡ��(��)s�
�1n�n�ª\z��TK���/��~��ν� ���+B�UnfQ⥊��0=�f3�I�Q�J���*шf�� T�Y|��5���6.t�9��R�sL}$�ÛR�!�$E1k��3� &_.�y�(F!J�!�K��R��󮖡!�p4"4%��!�D�&	hhɱ(Ӱ]��Ѥ��T�!�T���}�%&X�%հ����/rq!���� *-ƀO��5��D4T!�A�x/��2i�k�*�C�#F�GK!��*h���)�-M���� B�+d6���m��5��F[n}��B��y2/R�}#t�!��Y+P��Q �G?�y�eD8%�"�"7J�4Jς�x�e��y�!��=�|��0��H������	�y��.�"5P��>N9"C�$�y�O��
��R�/�5��@�2H��y�ς�o���b�Y*3n�q�!�$�y�NP�9:�
V���z��
! ��y��_�F�!!�F�+���.���Ē ��I��BYb�jO�ja~�P�L��Hŀ]Ej���#E�J(�{q�)D��xqKW�#��"$/}+._�y� ͱYv0Z������2=�����'��i1Co ����̓bK�p�''��w��Cn,�'�p̜yB�'�r���KTd�c��n�P�'9H5뗢E6&6s�3B����'����o�޴�W��_�Ƙ��'l=)�gJ$w?��G���V��E��'�4��!��ݳsgW�V��mi
�'20}�0� !3��S7}�$��'�v�qAҳ^�P�c���y`��	�'��!�e�]*�]y�Еj�p�k	�'�LpY��Ɍ��A���[�sb�%	�'kNeᑃ^�*5�����غkC���F6l��L��6�$�z��	n�ƙ�ȓI��	�-&m�9��ÁCCr���>�� �UȰ	cn�����>.JC�I�m�DhgB�I�j̹��.=RB�I�E�������$*�>�����mdC�9J��]�7�����Mԕ�.C��9d1P�	�DB30��q(%�Q0.S�B�	�0P�D��̇���5[�ۜb�C�	�����4$�(D�: J˚-8ZC�ɮ45�!	���:���Ş�B�I�6ޒ`% O`Ҥ����V
B�	�>.5��@ *����	ͦ~�B䉩1LY����60�6��`��d�C�I<"Ǧ�	�Z��<�Ĭ�*��C䉺"����G���JRgk�"n���'���j�oB���&���'����R��yW

0n����']D��]?vllB4hV�+Mf��'��T#,qW6q[�%i�0�
�'�(�q�� i����R���+BT��
��� ReH���d��4J���Y�"O�����NȾ��֨"<zHp��"O&$ő'P�e��8� ���"Or)���+N� D��W�Ъ�(Q"Onu�)g���	)f&�bS"O��J��;��{a�f5Ku"O�9����XKJ�b��:8���"O�ي�̊	{�5����P�ږ"O�\��������´C�
́�"OyJ�lW7�}�q+�s����`"O�`��ĂqNt̩��F|���"O�1�G�ʂ+~��;0HS�6]xa[�"O웗h�0UIZ!��l���y�"O��9ҡ���B�kI8v�hÅ"O����^�5�Ĩ�IA�n��,�""O��*l�+b�@�zk���QI�"OP�y#�ݦ	!輑���
l{��3�"OV ��L�bsN���h^fc��"O��O��b�X  ��7zLtp"O�L�'�_�3ȢaC�$m\��)"Or�@&섢H�����C�LK �4"O����C���.�D�C�9a��ZC"O��b	�<I��%m'��:"OQؤ�L�j�5�㬙(&��s0"OnЕE����,Ⱕ!��mD"O�����Wd@��%��K� �b�"O\�Z5b� `�l��82<��"O�}iE��A�6�kd%7R،��"Oܘh�L����[��H�xaQC"O�3dʉ� LR$�̘G�2h��"O�m!T�-nΦݚ�n�*c��q6"O��q��*�N䡵n 95V|�1"Ovġ�lV=b��c�-�3!H��I�"O�qzD"�&[�H[Y�n�~,�"O����"�����J
?y�p��'"O:٩`K�|EX���'N�g���"O��($/9�"]kd!�7Dɚ�#"Ojh�eB-g?P�s��Ih��"Ol��䄛>b��u�Wć�n�ʩR�"OH�j4d	-p+^	�T��f�� ��"O� �� 53  q�ș+xt�j "O0��P%"8p$�CH��xo\���"O��#"(��f���`$D	(F,XP"O2 ��)/d�	�Ì%md�l�"OP�eD��J���Y�}[N��"O̕��N�1f��B��9OS��{Q"Oh��D(�+���3I94���"O�Ty�	Y���Q)g݉�J���"Oν��Ȟ"}ܕP$�7^�ԥ��"O�T��A��\0��0B@0�""Or�P q�t��aT����07"OR�33ϲj~\Asb>)b @
"O�3u��Y���A�Q���"O�$臏p�`���b�9Z� �f"O�Eb��+]����Pk!��R~!��gJf�X�B�v�81��U�q!��CZ�V�3��	�1��e�V���jT!�$�#�0��1�h�4"��#7E!��^�z+\���ޢ~IB�i���!/B!�_:Z��Y �/A�.f�[dҸ5>!�d�.p������2o'�43�L�UU!�d�"6��g�W����g,� H!�\%
����Y���I&i/!�d���`Y�ِ���
v��uI&"O� H���o�&-���Q����y"O� �V�^��bI�ɗ�Q��4��"O�e��M,]8���w��`��D��"O֭��*_���(��Ap�e��"O�Œ��	�tH� w�ƛ_���ˢ"O�pq�I:�8x�����h��"O�� ��#0*��2nȁ`�T(@2"O�1��ٷJ�����ܝ&��T��"O�����<$����j��Y�DAʴ"O^���+�2=����'�T�G"O�����dG�,x$��`kح��"OB튷�Ɖ>�!�4ԜEc��95"Oxt��)>h��læ˟��&"O�A�G�-dX�RG��;rלTQ�"O������I)����į2�xZ�"O�3��(*��S��Y�]84@[�"O��+���� ֔�J�j�8+ֶIs"O��@���(`("g��.�Bd ""O�PG�F��L*`��l��+%"OPӢ�K�(�BͲ��K�O�~d�"O�̫�!V
>p�&�Ք�5"O�	)&��<t�D����F�,�"O���C_;��qe�ՔOp�qT"O�l� ^sw
Ă��_-5B`D��"OP@6��(�<�$E���{aÐ�y�l��,,���ElY�@��)�5@&�yBC�G��!�b��5�*�� ��yr�Ļ 7��qe�-	nѺ�Fή�yrg�`�Rps��T&,3� ��G͏�y�#�>�.��'K�&���o4�y����k���,�9v�5#Ң��y򇚍qXXdj��9b,-��"*�yR�� U| ����52V���
�8�y"̟9utl鲄m�1���Qg����yBcO��ƍ�Ƭ��'�b�x#%���ybGA�}w���NѯMV,����Z8�y�S�/�XP�>�ɂi�)�y�)�<7ш4��މ3ݐ�@�`��yr�Q+\9�Q�2;�Zv ���y�&˟u5�m�`k�<��<ڄm��y��>��+&l]�l�b���[��y�E
!���y��Z�8OT�dl�y"K_)r@|���C"fܤ��jW-�y�N3F�����T�]�(���-]��y�E5���Zr��Su��sF��y(T���MRgƏ�W ����`�+�y����	X�x���"#[����,�y��F<0�vD�(�l��I7e��y���-v
�tr�ORL1���<�y҄E=6A�h�7^��u�p���y"$K$:����B�r(�g��-�y�)�%%3�(2I˴�� ��Ȑ��yB�I���b�3. ��\��ybe� �[D�H$�vl`a����yr�!kZ�࣌ٗ��m�F�y2̋)VQ����6�8�c���y���*,�id��}>�a+����y�0Tv4H����r�@�9Q	��y���1n&!�#*eV�h@�\��y���< ���C� 4��(����y�#�9{����H�*�n��t-Ʈ�y�'R�0�$9KǏ�'�m�#-�)�y2�4YuT��t�V::���e�[�yr�T�8�<a���Y���DM��y
� ����9*K��
F��!p�&b�"O<tѶM�qV�x{"��$�L�B"OP�����C�ؠu ڷO=����"OzL"`H�.� X�4�<v�a�"Oh��VA�)\� ��fd���"O����ٯOc�	�B/ު>֠���"O�	
V�Zu�L�cm�BДas�"O����X�V�9�K�N�P��"O�e���4_� R ���E:X1;�"O�-qaC��|b4���	�RK�Ԙ�"O��S�уu�^�b�03���qE"OİX�۶��i�a�[�۩�"O2!a"ŉ�g���a�6k�QG"O"�2��K4���b@�n�|���"O�d�#+ؒ$�~��0 QoʨQ�"O�E�V����Y�𡖽|��'"O����)!z���̸֡M���X%"O2�	��d�Hz�._wZԁ�"Od�2�̄Q��eI�⋓IA�A{�"O�\Jd�i�����|̴!9c"O�8�Ƿ+�B��Vd\77W�ٸc"O�t0�!�:&Rڽxd�D8���E"O���c��?F\�Kub�J�hq`�"O���-45�A���"Of�	�-�E��ɓ��:Yipl��"Oڜ���ϔ��H��e�HS �hg"O(���N��I|<¡��V�컄"OD��YT�A�O�:
�LB�"O�D�/	X�.��5Q�
�b��"O��)��N4����E0V��`�B"O�E�"ДH�r�3B�&���"O|���FJ�t� x�Y4"Oʉ;�̎�5�L�#��4Ǻx��"O)���Ѣ*�&��b�8��t#"O���Q�Q�]ބ��bߤ[Y�U"O��x�JW't޾B�!A�@hūU"O���df	2-f6}r���/����"O*|0�Ki}*t���հO�p0@"O0}�P�W7e��m�1�E ���IF"O.�� �Q���!�ǃ|n����"O2�Qm
c��ɦ.�MV|��"OXH��� 5�̛䌎 !?~��"O~� 
��>}=�w�߶:Ʀ��"OJd�g19��R�B�����"Ox���PZJ��6��o����"O
�{��:d�0��J�h�S"O�UzsJ�G8��P��c�W"O�H� �1��=c X%�@"Ol��P�L�x�yaC :�H"O��[0d6	V�X��o^�9��"O��Ba�������ښY��p""O�h:Sʃ�E$� 3K���"OxT����v��%+K�i��\ɐ"O�}�t��2�,Q+ސN�28�u"O 8��O�/D����h�0Y�"O�t�� �,38�d����?��y�"O����:":Ȋ��D}B4��"O��x1e��J(p�a�Խ?��E�"OscFˉJ�Y;���%n����"OPK�ē#'V5�`	:6�Nka"OR�Rh<�<��3e�0}�R�A�"O�8"�^�A�-���� s<�5�G"O���B��=�ؘ!��ގ{6���"O�p�)¬b�; 䇇�H8�c"O� J����>F#���a��<��}��*O~T��&U�!����`+��)���"�'� �r�-o�x�Qw��K��p�'(*���q֎`1'��ʎ��'�ޠ�ȋ)`, ���	����'�}���_�\X�&A�6.X
�'���$��,+#�tIV-�|S�`�	�'�F��Ba�5f��R&��z�9Q
�'N�d�#Y��ىu^��~\:
�'4^��#�=Yņ���I^�x�|�`�'�ʀy��\�}��A��l�>u�(	�''�D�Q�@-{�~�l׵o�ԕ��'~�١�+�+@|�s񫞯hE�@�'V�e!�E�T��k�eH��	�';|��')հh���gFO%_`xa
�'�v��w���6�v��6"ڔQ�(iH
�'��J�E���R�Ȳ~�Dx[�'��r�M�
bBu��hrt���'*��R�Nk��0��[�X���'��@(�NG*]E���aD
<�@Y��'a�öI�i��!!��W�J�Y��'<�B�
@�m�f�������'��{3�2a�6���J
�=ֆ��'�$�C cԟN��d���F8�A	�'��	��$v;B�C�Ȳgp؈�'�>y��+";e�`�S�`]��'�Z$� ȝ�i)�X��M�O��<��'��i+w͑0r�0��a:=	�D��'��49Y�52 �qJ��0}��0
�'&�,�rjU-X�$5�q�-�M(
�'�h"��ьe��mj4� �%�v�	�'D�m+��A8>xp7��QG Y�"O���ϟ.6	�4�f��G/^E@�"O�}��h��o�6����ɔ0�\��V"O��ś����Vh�5R��ZP"O&5y�`)*(X��ٗoYZt�R"O�Q�E<x7��y4��z[<ݫu"OҐ1i@��+b��"�Z)a���^�<)��D�wP� hb���`�d�]�<��	:0r��3(A �pQ@Z�<A��H�I/�Z2`�#B&�䢞S�<I��-nO��X���� -�d�I�<���-+VD9i�oS�Z�����AB�<!6�мG�y1e���a�&�ǁG�<)V��6!r�Ƀ,��.����J�<�S�6�4�x�	ݸ+`(A�$)Sp�<��i�;��4�$O�@q>�
�o�h�<�3��*U�����,��pڶ��\�<���E=t��( �ǔ*P��Js�<i ��(E�G�.'�"����Fl�<1�GV�_�]����=��'�d�<9��B�t�U��#r�Q����k�<�@��_H��@L��=��%��[d�<�@��8E��M˕-��E�)PF�<)Ш�7_h� �+㮽�MWH�<�q(�':�8x����	(�i�i�E�<�D/���>�Ч��+h�2���Q\�<�� �?��p��<�<I ��Z�<�cŝ$W	ε�q�Glv�� �@�<�m$B�P�A�
Iøm����<��iY&u�j4���0���R�<�'�& <� Kľ@��q�hN�<���K�2�t�؅a��V�D@��e�I�<��ʐtP�gj��hq �VhPB�<� ƕBRh��:D�a#EАh���yv"O�d['"̮o���f�G>Q�tX�"O��P5,�`}$Lp�,I�8�QR"O�Tja�>�T�y��ܗ�q1�"O.����`��A�ǚ�9����A"O&���	�^ގ�y6	L�0�\]��"O�̑��M��n�8ǷmKfE��y�G*#������B�)��c�˘(�y��T�f��,�t8Lغ��S�	8!�D[�� 0+��Ϣ z� �ˊ�%!��� <N�Y��(^h�࢓k�lf!�d�)w�\ 1mGTLe��pe!���;�4����0J���)�`�2>!�DNO��a0Ș�0�6p�m��?!�D�$wQؑSV�<��5����#Z!�dZ%�0hɂZq��x�����!�[>7������e�X=�&M��!���V���d����K�V(<C䉳	߼�C�)K|��y#�/�(C䉇>ӌ�	)L9-p}*S ���C䉘5�pPDd߿}�85h�%��sC�I�18>(��(2�a�T5&�0B�7k�z��ł�2?�Z�a��T>m�
B�ɴ#
@���K��h}(��sgӔ2G�C��!J�^1��`2bBL�G���j�zB䉼XP��H�� .<0n�R����]�B�	?^�z�Cr`=k�\
(ױ7ZB�+8���z�(I�8&�У���>�"B�9{��ӳg�%@`���P�B�ɰ���@�ѨNMrdz�뀖��B�	�����#GT8_!<�p̓_�B䉿vd-Ӱe�x����~B�I�pT}P�A�/2N���	O�#�4C��`d�A$�B�����lJ�#gLC�I&'Y��Ƀ� ���Y���f�:C�0C�&�tN�ut�[�`���B�	�c���cg�=�Ρd��.�RC�	
'6�X a҃��u��R!��C��?P{@0���!�ћ��ۂ6'xC�ɈZ�P�8�cA�,l一�f��C�	jy��i� 5��f#ջ^C��f!�D#6C�*pmlԋ3�Q�3XC�ɁG�8!s7+��\�Pd�̌Y��C�	:Jgހ!&,H�|S"�1�MF!3�^C�$P-R���H�u�TX�c'��}XC��),��t���yVE`��;~y�B䉓|\051�JP0_P)���9�$C�I��^� �l� ngn�"ፗ�!�C�	V�Ƞx� M ˣ0G�,���[�<��K �1a�$� Gۆ@#<���R`�<Q��ϱz�T����:Vݩ��[b�<A�E�8 ������+d`�e釯I_�<!�i�D��}Au����x}	Lp�<a1ƒ%G9x`�gֶ<��|�%�D�<�0��k6re3����[�8�e-}�<��*K�|��Х����2(�z�<��蛐"[P��$�n��d2�$�^�<��JX+��tb0I�'Fp�`�j\a�<����k���[�-A1)�p(d��\�<�1���2b��06�[�E�X�<�E�:wx&	��GA�=�1�"M[�<!��t:5�^�����YP�<�B����q�-0������a�<�E	�]�v�bT� \+�ɹC�DT�<� �Xt�B\��!Iq���"Ojm+��i(��8�@T�+P9C"O��{7�J���̀�2��4;�"OTh�bA���&TXul��IQ����"O<�� ��P
H���b��"O iτ���*�3њ��V"O�+�&�aĽ�fH���˰"O4��w�'�������-�*�B1"O�5;�d�3.,���D�#��`�u"O������I���X��\���щ#"OR�
�+^��"��nt�,�D"O�3��ߤA1p!���,S�q	�"O�81� �
�Y葦E�=�0��"O\eH�� (��CQ��p3�9�#"OB(Z�N?�ɚV���n��Xu"O�y1�Z0"��w�R�I�d�2"O�@!�̞\��7DDf�
��"O4�	k��"�H���H�p��iD"Ov̒�m�6t���tH�:a�-��"O�5�$-�d~�"����uG�}�d"O��3A t.j�+r�^�y,��;W"Ot��e�;4�2��&��B�M��"O��o�c���`nW:/~��G"O,pY����]_���kޤ[�	Y�"O���g�;["4�u"
�&�bA"O�|s�H�0�J19���)�z���"Oġ�뒂
����-Ύ��	`"Oz�cv�q��QgR� ���"OhL�6��n F@ɑ�Ȇ0�jd��"OHH( ۿ��1I�"ێ�2���"O(X�i�lQi�h߹v)f�c"OB�c��l�]�bξ;/�:�"O=�V�4�P2aD�y谓�"Op�#燗��(�&�)G.q!3"O�V
�z�<���P?"��3&_�<��ĝZ����U�3*)sT��c�<)���N씰A`�&^�����o�w�<i��ʈ3m��j�#7b�O�<2Δ�F�I�e%�2AauIV�<�0�Ćr�¨���n���ȅ�F{�<QЍ�!ʶT2�	��*DD}�Yx�<���G�1�ҸQv�[5,*�YxL
]�<���̨W碍7,J;�6�E�U�<�
�S���A*��K�|p�RG�j�<I�	ύH�(4I74�P�M�c�<1uC�o8�l(e��3X�0иE�E]�<AFMˉo?���@����i��Q[�<	q�cÈmh AA9	L�9��C�S�<	���HN:��$,�AFXI�5��S�<Q��^�#���.�;���ct�Q�<�UkK�&y�e9%&�]D�y�@(�q�<9��F*g:�Qb���M{`Ho�<��gW	/���2��Hv����'j�<���S2�~���C|�)��_h�<)s��(��H[�̐�Z�Ȝ���`�<	�n��(��P*�\*��$����e�<�4�O/j����0ɟ�x�X:��Ax�<�O��G~z���/ 8Z� %J3C�v�<i��=OR��0���s�����Rr�<�gM �J�����I�e����@i�<)"b˥�|����"��Ac��b�<!q
�%Q�KT��7mnⰲl�^�<��� 8���0�>����W�<	��Y	 i>D*��_�v�1{UH|�<� ��\A����G��iMp���"O*]!WIT��<�S��p���"O�aY��=j�R6� 7����"O��Ө5z����1�αX)8�RW"O��gA�Ks��D��%��� "O�)��R�*�b�@��"�P�HR"O24e��X��نnW*�
���"OZ��B���a�А���kzy��"O�-Y�F_.m�^A�^78:dr"O$	� �"O�l�d�٬X* ���"O�L�f�C�axq�i\��q��'������#����M����'�KÂI��(��C�8e`��p�m�<��%%ٶ�p��-mR,���S�<� I��e�@\�� �'O:`�
t�Y�<I "[�Y�%N��6�|��K�Q�<9�I�ZAn@�	h����tL�<�m��z�qr�5�\�P�O�F�<��!@�\�n���D,d���?D�\��#m�͘,L�^�)G�=D������@�Q2@˕B�L,[�g.D����GсI�����C�T�W� D��fH�-^>"���k�ڌ*&�+D��CVeJ�`�,�jr��)�t&�*D�8aӭ	�P�j�)^TL"0�*D�d3���<�����m�52B.D��iq���xJ4*�	�#I, 3�E-D���%��ek���Q�N�9k�F�*D�����Y2f4�0�L Y*�9t�*D��� �>�2�(��v�ءS�=D���f҅iP �H�冫t\h`�';D�<SM�j��b`�-9�D܃�F6D�ȱ��J�>"�Q��.IA�F��&0D��	�GI:Y,&�[$OTq�*�G,D��8������15a=B��a'�.D�,�e\�H2P� r�Y=X���BDL+D��7� �5v�0�:�t�Bb*D��2��S�S�@� ����ԣ��(D��+hr���2��ɾ�����a1D� �5��$B�`���Ŝ�m_ҁI�n0D��S�N져���/<��e�T�"D��H�K��0 O�� 겱�B.=D� C7jEc��~^��I�C�ﲕZ�h�)D���%�Y��|C�ɉR���4�Q)\�t��E��)6�XC��46��i��jJ�S1VTB����]A�B�0o:�y�E�F�$ܱ`ۃ=�B�ɀK�E9��C n��=
�M�Ҋ�	�'��4���4RZ��h��� Tʜ��
�'C������k� ��eϙ^Y Qx
�'z��jr��+V���i��$XG�,�	�'R ����=WTJ�0G�J���	�'%���ZR8@���I�37��	�'7~�կOE��r�� Z����'���[���8GA���"T��
�'f�0aG���\��#KT#M�Ơ8	�'?���rh�Y�tU
sCU�v�rl��'#\���&�����֒��Ђ�'�����	�h�Qr$O-]���k�''ܰ+�l�!!�fq��1M��b�'����V#x�49X�e�@�4L	
�'q)�d��[�J�7�U�#�0,�	�'zq8R/Q9wf�M�Ph����'�p ����$\ Hd���Eڀ��� �X����u<�q�fPb�c�"O�As�D��Zt0��@�P<�#"O��y�I02�<}�d%�=)2���s"O���`�*k+�A���Ɛ}|�8��"OFQ�Um��)��DZ�&'o^�)�a"Ou3��?� ���13RER�"O%8���nA�lh���N4}C�"OxD3"$@�Fn	
 �0R]��"O���d�<�45�S<X<p}2E"O̔�E��0;Ц@p@���E2,s�"O>p��oK5t��l1灓�&�<��"OH�qq�"z�J�oVb<K�"O�e)�+��~���ûV2ʌ��"O��jp�4�&���S�~ ބKd"O��P��T𜅠$G��8�xg"O�p���ύ��W��H�L}�"OJ�CL�K��8�n�7w%���"O���1a�:f|�tL%\�� �"O�$��C)t��'%RJ��٣"O2��� 7�6Ő�(�}Fz�	W"O� �%��J�X�'��j,|y�V"O0䁱%X�Փc�ݦ1���"O4i:��RHoD8�TD� ��#"O�j�l.8��̪��H(�$�Ip"Ox�zF�]�(�vL��.��QX�"O6�)Q�SZ���0�kB ����"O���/c+j� q�>�g"O^ٺ�T�w_��ꀡ�Wraa�"Or�S��ϥ>`�7AՀ7�4}��"O����%��bi2ri�/r�`$"O��Ȣ.ً}��y�
�`}�Pz�"OZ�a��"8HD�ó�:x�"OFYb��Ʋ*NЂ·pw)�0"O��;���/�@X�/C�!s@5��"O�,�.L�������=VZ���"O�����]�Ep1bT+�a]��h"O��c�2��-�	�3�6���*O��#+K�e#���~����'>*9cFˮ8���J���3�'�M�Q"�.gT�I@��I	�L��'q��QƪO�@�.���MH����'�����m}������80���	�'�����/T��ZP��ªDIf��	�'}ePn�	h<���a�(l��C	�'���6'�h��1�4F�7X��	�'d;����jp��P�̇ .QZ	�'MvI�� ��8Y �ɉ%NT���'��Y:�Ꝛ��8E,˿i��K�'>H9X�iO ��ュ��w7
���'�n�`�oʌE-�9	���j�8��'�
`ak[ �d|uʕ\�֙�ʓ=���`�F�2I�@GT�W |͆ȓ��L1���vG�̩�N2z�ȓp�8a�Ve�H%y4E,S�65��S�ڱ,׌U�N1�A *iJ��ȓEB�YXuF*@W� �b�Ĩ b�M��h����&Kr���ƕ"7�td�ȓ"�`��a$Et��9�ڮD�!�b,e�6d�r�E	!C�3a�!�-N!�1��$>� (�O-�!�$S'2��iPcE'=��҇�ǅx�!��-r�rѣ��/����9M�!��Nq ��	J�MbrA�e@M��!�'l���K����@�2}Y��ϝ�!�� �<���v�"EQ$�R8WK��ʣ"OUj��I� Y�-s����-Z��"O^y���@p*a�f�x ��2"O�$@�@1nsQ�G¡P���R"O�9�P��w���G��#��`X"O:��t�QZʎ�xï
;�UA�"O��u�<����	}R��a"O�ϵ0�����u{"O�]���ш�d��T��
����"O�� ��<�Br�h^!a����w"OإsSbO�=����!A�zJ�9v"O�Ż��Lcڄ-K��v�^�k�"Ol��B�ρ�Q��'T({b�'��	�����蟗N��q"��:o����y�	\���s�I�8�,���`��2�(qA (D�<�R&�h��Ѓbo�����%D������2x�Zwk�|���-&D���S!�kN�ҕ��>��q��)$D�XAC�;&�!�aI� ��"D�[��MI'�P��D�uj	�F<D����Q6\ߞMQ��R9���v��O*��0>1���
Urpa <N���1W�Pu�<q��B��W��'���!�-�L�<b��k]�d��qg6�9�G�L�<YD$4�|ɁVӑG̕q��c�<�2�ܚS���S2�@��p	t�WI�<�'�ִ~�PȩSB�j
�h�B�Hh<yrƔ%A��*�$}dm�ŏ8�?���@U�*�a����,]*�ф�u���U��n� (0��i������QZ�Ƙ����2�	=$����ȓK��۵�1+qK�� �4�.Ѕȓ_��C�ЎbR��vg�W^�ȓYQ��Z��P~�"-֑j�����؅�!₍,iL�.8�k�D�F�<�'i�;Oy.�����RvF�k�<!C.F&@��dڶ�����sc/Sn�<�vQ�[[����˗w=f��lC�<�dhF�$�J�����"=�g��w�<�"��u�t����X�'�w�<a��ƭn�,���D"95��B��n�<!fdP#��be�hll��*�k�<���ŇNq��ĭ\U x���<Y�*�3a5$�"@�-?��K�)�z�<Q��8N��C �K"�W��o�<13hԉ%�4\IR劋$��(�N�i�<�U�J�j�T���!��_2�k0a�n�<�ň@�pzH"í6p�
1D�Wd�<�A����V��4�t�]�<�0��}U������|@�)�Z�<�a�C�]-� !�
(#��a�c�_�<�h�#B�l�(���4��pj�E�<a�d�<b><p@��~������D�<��Ñ� ��(��I�|m�}�&i�C�<����&A��H���B_�A���C�<�'Q`�`p`@��?.��2׏�J�<��JN�#�P@Eh�RH�tmH�<�w,�3I�ԁ ���� �굆�{�<y�!�(%��
Sƍ�!�f�rp��k�<1F'�$U��l1.�IF��b�)Md�<)��INwx=�C "nz�B�.�`�<	T���;Ǩ"�#Ӕ&]N�*a�_�<�d��$ ��[v`
�?�4"O]�<a1/�"cY����J�n@��ր�q�<� �`3�/�5?%2�胨 �V��C"O�t���3=��R'�4D�f�d"O�q��،_�zq�#[� �"O��ZD��4�&��3���<��	�"O�upG�O0"\�� ���;B�h�"O��
�O���)Y���H@vi3g"O�IƑ2Vf��S�G�5�6T�"O@4�aәE��@[;4U�R"O�@АKH_��ٸ!�S(���c"O���#P1�r����܏� ���"O2p��/V��ĩ�L��DHx�"OZ,��ջ� tRa�ԇf�9"O�	���_7�M��*@g�6eZu"OU
�Ȉ�h��}�b�5��3�"On5��A.)�f$S���#� 5x�"Oz=���zE>A:���%r�! @"O,}Q'���v�($�c+@�}�ܡ�"O��y��V�3��|�f$�%gq�i�"Oح&�&<0���"_~]�ȡ"O��`#�6�-1��SP2�Y�"O�0C���V1��O�a��yQ�"O$��Œa��ea�}�<�Q�"O�-pg�a
F,aǣFh\���d"O��9�⇾K��a*�3�����"O��!�!X����J�$�V����g"O��@s&^�4$8Z���@Ӱ"O�=xcϔ�i��h�b��Q�4IQ"OT��\@8�qd&4Pc0��F"O����4 nrpc�]&rZ�r"O�'f��<�}��=V6�g"Oh��&A	�_���aU�AG�麆"O�I	�d�$V��]���"/34�)"O̝jA�#��$c��k�0�p"O���a�C7G�ʡ���1~X@�0"O&A���ԍKb2�j��Ǣ�pP�"O$�˰r�Ę�0�p�@"O�ز����.����V	-��2U"O\t��`&�CpȜ06�E;"OB)!<LwJ�S$���I'�kV"O,0S
 +eCp|���C.]$z��"O����&C��M��$L�S��� �"Ol\�EE�
EP�TD���~�:%"O�e�a���f��iQ���4b��:�"O\��Ə�@��x2q�̵lD�Q33"O���m/m��H�%`U��@+�"O(�Sc��<i���t�A�k!���G"O������RAT����.;|��"O,�p���V�p�T@�00�ly�"O�!C	�/8�vT1��!)�hB"O0l�t+\��TL@�Q � �"O%�����"�d���c�.;*T��"O襫��,����ƾwxTr�"Ox�#�I�2�n�Rg��k�y��"OX-3����>8xW�ޘ M���"O�-+�e�'�>I *\6+�nH "O���g��mTHi÷�X�H���Ґ"O`�നՉYp���ˆG�^@�"O@�ĉ�p0�qz�֐<��JU"O���G�d�b)�6`^J��� "O�tB��O�u�� b=`Ej�J�"O\T Cm��GK�蒷���R-��f"Ov\ZV	M7-x�cӈB�Y�1"O�ݣa�KZ�dAW-�V����"O����V e�z`��ߐ|	�-x�"O� <�aW��'vR�[�l־��aJ"O��9�N�_��q�gE�
��\jS"OJ��S"6v������m��"O��2!�v""�c�%�%#�Za��"O(P��,�(��aC�`���"O�4UnL����VdM�H^�a	'"O*��cF\�>(�%C���D0��"O����冫{^d%����k�"O���q$�#6�eaQ���m�Q�`"On���UU�`q��_�#�.���"OVYq�)�9Gz�1���	��-��"O�]�!]���WO.!а%�Q"O��8R��g��ތD��q�2"O�����,���d/>�bm�"O��`L�mT �&#J�4$�w"O�=8ek 902����z8!5"OE ��C��ʼ!�J�*w�S�"OZ���Q�_�l�j�h���֑�"O�*�8d8���e��Op�"O��Y$_96k����!�np��"O�����:\�\y`!�<Tݛ1"O6��^�$�5�ӼH��"O:�hQLV�_��h8����J�$(J�"O��a�2S�d�����5ڴm2&"O�{f�ɟ6!�8!(�	$5T��"Oj��4FK��|���Y-��&"O�4�� jdHA挲G:�҅"OzX���u\"�2��F�kQJ�xV"O^-��_�]�h�Ē2NU$�"Oܹ"W�s���Xad�IBpd�4"O|q���b�ՠ��@4F8|��"O�r�%L�	���������̓T"O�蒐�P/�� �������'"Ox�	����8T(N�k�8��q"O�Ђ��1^%v�s���1�pP�"Oʤ@��"U/����=����"O�)�Ș�pn�3��K�k����"O�����M}(��b�ʪ%U�e9�"O,�H��d �Ҧa8ve;�"O���'� O�\�D�ځC	�$Sq"O��AG��8 �r���<�`"OH�U,�:�٣'T  z"O�<���2)Ul���GKAPHPv"O<�R��TN�+c�@<�@r�"Otq�A߷s�]8�X�v�Xw"O��� U����1.�~��ͳ"O
Uz��4.���yG�D� 7&�bw"O"5[ƈG)*�Mq4m¸�J�"O��s��Tvة��B.s����"OK<8D$P��$�H��P�b\�P"O:,��%U���Ʉ�QY�"�1"O�y�v���M�vl�ڰp�"O��a0����.�x�
��^�r�	�"O�����S f�
l���Y<�a�"O�9��B�2�.�*���!~���g"OF%{To�;0�̈�A�ox����"O0őv�2\�ԑYCA��z@��A"O6�����0��M�g��S��"O���������u���֡'����"O��D���<�r���U�U"O֙#�ő�:�8r�ѳ�>u��"O�5+B�צ\��i���7Ӏ�02"O>�;F���u���bI�B��ac�"O�X�g۾,Qڝ9b ܂[�"<�!"O� |Щ�n�`��9�դ/�.ɣS"O>��쀓_%�5;$&`nD�"O�b�k��x�F�#�dZ�@�f��4"OP�x %H�)F-֊���34"O��1����)��ڕ	
6,Ȕ(�&"O��Ub�8e��Y�'k�N��"O���a�1?�ȡ@t�	�@̲��F"Oj��'m��?�x�P�!�&n)d���"O�|���P]!�s��1��s"O"��d*ӹ!�U�W�C�ix�Q"O88@�$B�ɬ�c�Q�h,8m9q"O<��LR�~�]��3&��ۧ"O�X#q��q����3�OS��ȧ"O�A���[�z�[d*�4tMS�"O�XQjH����*M�Z�qd"O�rGƍi�lu�FU#5J�L�%"O��2�˨Q����v�G�s�^1��"O*��A D%l����̓�~j���"Of��a�9��pqo��/;�� �"ONU ���b��	5%��+Τ�q�"O�$"V��!a9!n�rͰQ�"Oʜ7�� /�y1�� p��qK�"Oh]{b�VΚQ���,�lL��"Oʔ��\TZ�<�5A R��u��"O@l�wo�/��	>f
m��lA,�!�ȣ�vyjF.M��L�;�؇�!�dV�Q�"���I�>^��[դ�f�!�$�;J���Hԇ�.^��h�F�W"�!��K�/��觮��uٴ�ׂIi�!�d�#Mʬ��"��-Nd���!̮:l!��!,�vȠ��Hl�Fd���#IS!�\�Yk�T���ְg���@EKH!�DL13�1�&H�*s3�(�/L)e�!�S(��)J���8�"�r�n�30�!�]�?��(�*�$B=ࠀ��!�䞜X@gّX`����r!�Ē�˄ y�^���3�1!�dO�>�@�i$�^x��%�A�^�!�d�S�$�"&Pb$<A����2=!��s<^}��+AHK�����-!򄄂M��4�P�p���`��w!�ʽ=�~���+����" C��!��}{��e�^!t���BBֵ4!�D�(4[<5��-L*��84!�d!��5���R�[;_�0e���^�5U!��a�Nx�f��!v��(��΃�Yp!�Q��^pi�,E~��JA��$4!��T?�B)hAH	�	���2%���!�d>Wxx�t�Ҵy��Hwc_. !��
�j�����L7ri6���o��}E!�Dɿ:{^���Iʔ8W,D8N�R+!�Dʇ �a��'ʮ�@Oլ5!�ݯ�"p�U!���I
�
w!���3R1��csa(f��Tr'6%�!��Y*����I�-.�\��+��*�!���1I�P��BۗJ�Ь��KJ'.�!�Q�m�X
��S�J�:AB�@� �!���y�hI���LҸ��#I��!��*`�̤+&(IT��W�+�!��-8;�%.@�\mL��m�!�:k.�%�[�V�c�Ǳ ~�x��'�䔚%�?]h��HM� U��0�'Wj9aA׬1�Ni#l��#�q�'����Q���BJ*&��=a
��� @�pVЮ��y�1E�}9��)E"O"Yڡ��$@E"	��c�ph 4"O&x�2 �R��"�"�\0s"O��Iš\�%t�L��ᄣsy0I�"OH��6Ł<D��e- >X���"Ox���	�B�~�[�I�k'�a9�"Or���艑f�N����Ԓ;�p��"O�� 윗��񀅋ę���R3"O�H�W�Ϋ7A�܀���0<�\%�g"O����H>Z��]�v�t�;"O���j�7<�R�t�)@���"O��Ǥ͵#-.��3$]�KoLՠA"OJ�ٖaM�9ܼL:��3o�|��"Oƴ��i[�U(Q'� <v�q�"O���Á?���Xî�4JJ�"OX�!R<�¸`R T�4�*h#"O��p�A�0�4�iaNȋp��"Oi�kh����)(�|X��"O������!�f����ײ,�0���"O6�3!L��/�@��}����"Op=a�%�&�C�l�6uz�B�"O���́�a�`b��C�~�T�W"O<�f�Kh��%A�,�B�"O��[�6���1n�/ܱ��"Ol���e��c`~@YCιJ̩ p"O~uyp��ytX�@�Yz��Q"Oɀ��C�k#�aB"���s� ���"O>aIƁG�����쏩=�x-�F"O�U@j�7���R��];�Tڢ"O�=��H�5�-�J�[��	�"OZ]��B0A4Č{`�(˪B�"O�ݱ#�{i�!ZC�^$L��"O�E���:>̘��(Ҫ%T� �"O*�x��V"N���9岹�'"O���mX�.5��� �ہ��y�"O����m�b�4�t$�t��"O�ڃ�ŀo����m��E;�"OXll8Q��G�G�)�5�"O&���=-���0�.[�!E"O���%Q�p�Ի��]�x[�"O��B/�To�q��n�N���"O���c*ܯk�l٣��X� T"O��:`%˃%���+��7�Jh �"O�Eٕ��J㈴��1���"O���7���@��舯
4�H "O�]�t@,N ~,R�a@^"R�"OVU%"�76bd��!�j�I��"O" �3�R�`�0����|H
`"O\�z2&A%~m�� 
ѭ0��"Oν��k<�rEh�/R��-�"O�RlI0$��� �N���8�"O��R��3���:2o	9\��X�f"O�� 6�� ��1b4�4e,�A!"Oi��,S� ����ɋ	2����"O0ċ�e�,5bT�� J�-^���"O��$�Z*#y�30@ ����'o���'1����ƥÌq"��VM��!�Ĝ(Ca�J�M�s<V0p��0,�!��H�w4���GP4d�h#�� (�!�d��<���CÍ%G����#g�Nn�I���=��ϸ'�Z��D��PA���ݖ I�D�
���y�@ṳy�s�O.	x��b�N�䓲0>1p�˺d��+G�!�̜ �!�w�<���Цmx�:4���"�r����L���=� $ �1.����r dR�]�D��R
O|7P�Z��ge�FjH˲� 9!��!.��p�$�,;D��ƝV�!�L�;���gc2�00D[�p�!��-�b��6��� J)��c\�7�!���
��<)���h�*!�d$u��l��i
/w�УuW>�!�dυ�+��C�&�����l!��;a�ȫ�䎌$��䍶c�!�D_�2�t1f4?$�C��D,&�Q��G{*�P��5Q�Wyi֧� HdJ�"O��@�!pz�`!�^�Ф"O佐��gmb���v^`L��"Olps��C	fT�"@�JoB@T��"O~��$�]�$x��!ZX&�� ��>�S�gL�$�2�E�@���S�J�nw>C䉓t���zQ�ɱ\��dy'^z!C�	Y�$��B.��r}� ��иn�C�I�_J��U	̜+��y�g7!�B�I�\pLՃB�&&�A���E�R��B�	�"�f��������1*Ġ)��B�<[���5#�
z�Pа��4I�B�	�D��  ��G�1ت|��7ݤB�I�?� �갃�6H�(pR)\�`3�B�	*�5h3�=U�j$y�d�-U^�B�ɾ5�4X�7�D�M��W3c��B�Ɂmax$�gg��2��i�[�g(�C�I�!&Ҹs@�͌otl�[�a�#��C�I�/oZ7`��RL|UC�j�nxC��&�f��O� &��P��)f�C�8Jzf�`�ML<���;gE�7{�C�I';v��j��H0�����zzC�	M0�1{��U�N�!bA��B�?8*�ݹF�R�<���rp���$6ʓf�:��㗷TZ�(�SJ	0��������h��D6pl�)���&�E{��d$�&L�
|J�K�E(T��kM�yR�D"6T�'K�? P�۱Θ��y_�(xX\!�#U�>.�������Px�i}t)�@BЧK���s��8/��(��d?�c�8bfU A���H�/�l݅ȓc��t"�hl⌹�,ٺN]��ȓ4��#`'�41J�S�	�J�x��?�yr��R�K�v�KG-ڱj2:��}��'Z�}ۀ&�=��5�E*԰m~T=K��h�<�&��%BҥʡGC�l�ҙ���a�<��iں N���$4�@a@a��b�<Y���g��@�%N\&�܉R@�j̓�hO1�R��E���[�R2��`j\�"O�Z'��y^ ,���x;`��"O$�k��]����㩒�`8������*LO�˔,c$����Ǘ>#8���"O6�`f��	7n��g��oA8(�"O���ٽ6�&]�ÈF�Xh�)��>�,q*����կv$��ࢃ�Iπi��ɲ���װ$���&`AvT�b�m�!�ā�Ӝ%���_�`E�����C�,��Iqܓ��Z��gԜ)�d6(��Wz␪֎1D�,�!N��&lZ��!�E}
�S��-D�(�h�n[ ������49"&D�l�@�D�Qa䪃>uD�Y��gd�آ=��q�'j"������o�Z-3��#g���)��hO� Z2o��Ce �.��92"O
����c�hw���1����Op#<�I?�'?�  }[r���T��Y	���"zj勦"O$r4�
y0Py�Ӫ0��W�DɃ��>aK���O��J�n��dI�I�8�V� ���$]?�E�"|���pkU�4�f�BAOX�<���ʢFaX��� E��b�Z�'K�?ٳ��̨M
���I���ݱ���O�C���Aۄ���(_:h��e9F�% Ġ��d5扈ub*A�k�eDt�hF!�3���Ox�/LOF�t͎�E�R��щ�P]�E�"�'��*h�bB��w��a1T�N�{�!�$&o��p��1rޙ�Pd�̱O�����/���a�܀_�����ԍD!�D�2&~ջv/�
.Uh��4�W1~�!�dշ&�,�SÂ��@������!�$A�}��A����a2N��5 *]�	e��p2P2CRQ3��ؒp�Ҩf�5D�8���&�&�RG̓��z�)��4D���暉[g���uGB{�4��F=�����!����	&�hW��7B<,��w"OR��S'ņM�����,�8ؤB�_�G{��K�����M�H$RPS�ؔ'!�ۙ�䰛+Q�C��@z�ɢL�$�P�S�g�	\p�B�Z'x��PЎ��0$�B�.d�-�DX�=<��凋"m�t��S"O�e	TM�tж��dǣA�@��e�	`≁��OT����.T�R�q�	-q|D�
�'�Xp�ӣ�?ZC~|Qs*�e����'>���&� Gc T���#r��D;��$��sD�'��Ov4���5-vi���V�����'����eG[�(AL Vv�i2�'ў0D{nȫV�����l��tC��+٥��=эy��C�>D���� �nȞ�x�a�&�y��3�6|�'�H�d)dL1�����'�ў�O��b"ύ~(ф�=��h�'��i��6-;�p	��~����b�)��<���ʰsq �ŌQ�|t�cUiYU�<�#�
P@�ȡ�ן""�-���j��D�'Ê����S{(�Z'Fe���3�'@���#D?T���J#��Yz,���'���sgML)���,Y?FA Ժ�'Z��j�-̶u�QP�H�l�h��	�'�v`ѱo�7�;�/	fv�T	�'�|�alF�@�T��jGa���S�'{@����&�H�ZҬ�S̬�8�Oh�H�������%.Þ�6ea���W�"��Q"O�$���j犡�&�)��kg�\���	>@����	\;���x�%�k�!��R�؉�R�K>dHa�q@!�$�*���m�#4-X)�W��i���8�a�G�A>��� ��h�#�"O<(�B����0o��&@��:D�t� .,����B**� ��=D�x:E����ɻ檊:��i�O:D�r�nYH��a�?�в�6D�(x���(�l��7��/S4̡�E'D�Di���MAHH�����L���:�O�˓B��	C���)ds��C�B\�U�2-�ȓ$S�}�Հڏ.�4Q�jF�CMDy�� ���DR	A�:���g'-\�����"O�A��K�%�f�aӏD��l��i%��dݿw�D��1��;JX�P�Ϛ�!�;���Y&�� :�
gH�
�!�D\e��s��p����R��H�!�Y)+�v�à ��#�X��Fm\�9�!�� ����Fr�����,4�V0� "O� 2���3r"�e���-N!z1"O�0�e]�lN��ɇ|����"O~���V7p�(8��A$�x��q"Oȼ��I�, �5� �./}�ܹ5"O2�JGH����1���z
��s"O*Qh�F�
K^a[C�19w����"OJ(��aQ�F:��m��¬�&"O��JW�.m*mN�5��X�R"O8D��B˻jEFqkG��UYd� "Op�X��C�a��'/��J�"O�}`@,��j^����N��~�s�"O�E�E�F'UF�ҕ��qJ���"O�%�7��ok��Xo�]1F	��"Oa{0I[�I8��RW��#T��	`"O&�&�rH�$k�K�
1��I��"OA�+H�b��i���+;lP@�T"Ob��ׯ]�G����th�/U���7"O`5���Td��GǓ!Tܡ�"O�[1Nԗ{�d34菔"7fU;�"O0�S@��N(c���Np��!"OFp�!*~�R�jbe� �:|��"O�tJWo:N�-q��
�B �q�"O|��P�"��y�����4��ݱq"O�e���Ǫe��q��Mٰ4��	1"O��H6dM�D3�����L�@� "O�e�r��`�ɗΝ;?�!�"O��cHt,4[CM��r�\р"O�t��"%?��y����J z��"O���O�/F©m�-l���rI{�tJ%��2s���2��*��z�>��swڠ?x�h���a���ȓZ��環+ļ1�R������JzqRf�+b�I�R�TPψ��ȓd���^�x��eI
רM��^�Xq��=1��1q�L��ȓirl�HV�Z�=;P�� �F�.8��'!2��C��I2ȁE�! k��ȓ"��(�p��0 �!'#>��}�ȓ+)��am�
l4p\Hd�H2/,8���8�hq���� 2@9�5� )�8���%t�!���W�"�É0'R�	��V!�D��f�jy��lC�^x� ��Z���7�+,�9�a �+m��݇�k�м�u˕�_9:�Z �A��,x�����agL#Q�ꠋ��e���w�4�'�hP
���>Y�+�$�N�{���Z�:%����Q(<хC��R��Y#G�X,�����D�܌�9�jX�s����2kM���=�'��c��A���2-~U��@�����*l�րI�+B	e�G��;�����^���sЭ��B�	D��aT�LD�P�E�^H�C��&� F@�f\�s4�Nc��C�	�/����ŕ�uu|�VcJ�$˶B�I:��ZCa�XT�&������>y�̠�Z��D	��\w�Uh�N�<7.Ñ.�T`���1�h��F�'��#� ���$0U0Q%<*({d���9��K_V!"Q� k3�w�ֲiI�����v�9Ꞥ�����@�R3![v�v���ɻ8P�
I+Z�(|
��L&Z!�� �t�h7��������(\6�e�'E ���T���=�J����\=Ӹ�D,N�BE��&���TW����
�+�>aP����mi4e@1;����'������c�S�O���Id�^�9DH0eF�J-�1�ܴ?�!��؍���㏋p�20�E�эl��'�
I"k�b�s�1O� ^���ȋ�Fq����I������'{V�xcm� $�
%h�%
,G��h!NU�_!4 �=	��)�IT3!D��5ł>U'xe�
ހYS�� �P�F/+�$���hU�Q�j�
��W�x�u�ɭ�0<Y�[{���S�ޒX�@l��Zy�.�yI�OQ>U�1�v�:�0��۱|�����fmӀ����$k`L�&��^�vh!�Ι�*�f�E|�(��V̧i�ig��(J:F�fd3/B"p�ȓ�0u�2r�|�%d�f=�	�Q�5{7O�I����D̠� X�% �䆃`K^(:�K2D��;B�ލ6޸c7�~� ��7$�<a��.A}��	��0<� �ۥ���q���6���PO�hx��:��f�6C�D�օ�����#!"���޾�MK�OEP����aQ1R��}V�p�E�0O���|�7,�*C6ʼ��N�	"y���W
YK�<�J8M�>]Aǯ� J�-2������v���??E�N�^�L-��͗�,�j`�D�6"O�@c0��2%r!�A-�$WX�M˦���Z��B���� ��3?xUk )e(�
TL'D�Tq��o�� @!G�7�hTh�c1D��s�/	/�Jɋ�@�KZ��l.D�����N�u��ؙ�M�8o�Ո�e.D�HPP+�!�
��
I�f���1�.D��Ð	��^�)�p7TR��.D���l� _��1��~W��ٴ(#D�8�1��2e�&$����)`d"�2$��9P
� bvHyc4��_��@QV�<��(v�'�q/R/>3 =���GC��Y	Óx�~��1��'v= ҧ�!�d��Y��K���*��i�<i�A�,<V��!�5��,bF��s}�M8L����ѳ3�1F���WX%hf�E�.�bŏ��y"O�*q✲�L�,`����(̕\'��2�O���*��C��H�M?�0J��	�G������#���9#�8�O�D���"%�.�y�OM�@}�����ʢH�� ��d�ޤ(��;�O��1W�Q�Z� a��L�tހ�@�I�9�b):"�"�2��� 1,i�[w��-�!�	�{��A!!��0)�YR�'S(�a�OZ�B4����>�����'��E $C�_��5�c�[�KW"�I�E�O�E�d�#��5N�+��r�'ߦQ���ܧ�Q��%�T�X��2�Y�r�aځ���Y�=i���/������?U���]�Wۉ'?��3E��<F�"MÖa���A	Ó*��%
F�6�Mk�j\7��kU�-d4�`��q��9���BaG8�4�QfI��U��ɵ7��鑶AA\�VH+�dD=pB�˓Wz�bQM��	�Fmͨjr�A0��V�ٞ!񏝓k�Є��,�]: �����2���E�I�hI��'�J�	g�9_Dt��D��Z�ʧ�r����$��G�`0�i��x�bO�v��4Ȓ#	� ��:�?�<I��Ț� ���a��0(H���'K6U�%�I#y�D #W�p
���O[�!��\ ���v<`%@��?���rR)H&~�L CWr��P����RCC
�>x�sj5O�1�
.�4�oB?��E����l����#�M�2���Fr�m�+�3)���TH҃)���;��[���Rn0O����h+;�f����&�v�ygW���1C�t����ݝ,3> "C�8?&)c@	�^o�ŉ�Â  �)H˾d�t���
̴B&&�Q@@�[<�!��*�Ek�+�.Ȉ9��ޚ0�V#�3jkz[1���f��C��F!?@ �V�W3Y�1#����y���zx� �G�->,!�����?��G@�y��yX��|������O�䍑�ɑ'���B`kG�y�,�$H���Q2,x�����	9.��J���F�r��s���"�L��	%4v*���O��<�P�B�D#��S�) ����8W�I`ΐbǥ�F������s��t�WF(w]�x��(�E#�F�@�[�'����
?��;�����E��!jAԼH���9c��qэ�$P0�:񃉍b0�����W�V�V�QoH<q�	�$=�ޘb1ȗwR:��n�!U��]�c��)��lYg%SY�z��IἯ�7�$h&���4+�p��_�)&!򤝞'�4�Z2+� ��Q�d�2Q���a��+&��p@��TJ�$��ݞ��O�����2�B�&}K����'F��C#^3��Hnچ>�$� e^Y��t�G0&Y�jR1Q��ɿ,��iz�`YAȰ���!�Ǹ'�Fa�P
� *J�mE�$D��I)����Č�V)�գ�˛��y
� bEI!gS(�Ai�~'2�C�iW�T�Y�>Y�h3�gy�6{i�1�M1t���q1��5�yR�X�����͙�m@hX����5ŊQ/ZZђ}��>��m��͓N��9��'�:? a��(w� �YA�OJZ󄛾8�2į��@¸�v ϴ4�!�$M�S�ً֤�6@9�a����0r��	�C��X�I9���{C�|�O��
�.j�Zx��97�L԰�'������r΄���ޥ+��*\�Z��I�I���I������g�
�~�!��s�h�g�Q�b�E��ɽA�&|��f�c#�9tn�.97 ����,(��9���B��OR�SL��HO�X��Ь�|�1�O�q�I���ʑ H�A1�`�"�*V�[�v%�b;v��'�i%X�B%Kٯr�|ʘT�p,�V�x��a��<�~��I	s�*Րc��K�4�bm���ޟ\��˞'��		RB��9AT(��"�����x�'�z����J�S +C;yj`!J���� �#|���ێ0R�
B�̑��h>���9���*�@ل1��%$�O(d1��(w��`���B?h	�֢��[~v��s�L>���8L��@S���zq�剁z�������l�x��#�վH�,�>�Gيz渱���'�����!��޷	0^l��Ѡs �!a
d��U�P�%�O>�)�/A#d�F�# +�
�@��Q�O)V
ހZ�\��N��S� �f��MU;g�䓱CS���P'�(����#��,�!�dH�iL�(�CB�
W�(0�A�>!��'�$AX��xI�-9u�)}�@G0����������N�ȡµ�0����Y�����	��/�-��\P�� ����j�� Ң�0}B_34�2E�}�'��i�}���#�O�!/Lũ�����d͟��^��	r,�4���ۀ�ں9,Tqm�8E�Q����U8�h+U�
5�tmGꞯm���<ٕ��(x��!h&`"}�O�xec���8q�ő�*G�=
f�_�>�6t��"D�h�֊Z�C~\`�s���{��C�K����q��	h'$A�3�I�s�#�����Q��_�Z����y�l�Х�7)�4��ܜR~>0)Jå	W�l�
��oQ��
� �'e$]�ڈu��=k��d�kp I�	��ħk�F�����>6^�B�H��B�`��ȓ?�
��/��
@��
��T*?�P�'  �ëEV��<�OQ>]��S�Si����<C$l��A�)D�0􄁾m\��܈(Ύ�beK"��ɹW�5#e�e�3��7{�bЁ��ؿco�YE�]�j����P�y�lLA6m��b0c��V?��UjC��g���	�x!G�B�$!�`(V��2wpx���I9s�1!!Dq� S0l�Nͅ'&֬IB`-��B�	�VB���!�3����� �RJ�'�>�١��A�S�'kR�uia�D41(��� �P���
 \���\�T�ҵ91��'!�ȓ�������-\(�1c�aOԄȓ5�Z�Ғ�޵Y��0��NN��ȓr��}�sG4e�~�tGT�PD�ن�-=fU��ըg<xY�kC51��ه�j�E����{غ�x4�G0H�<��$����s懫pj,p"g&V��U�ȓ�携��ҴK�r�)�
	�9 ���FU��0"(̓OQ���D�o��Zw�D����!�Fa��E P�B��o�2 �*;�O�t��,� \�|	�L� 4P�e��' ����C]Z���ؖ59�ɟb��!�1�L�y��s4��s5d�Y�,٣q����'5J ��6(�l�E�4	Ǯ6��N�[ِprF5�y"�\��j�p'�ǹ7��#�>rF��!�Wt6z�'��>�ɝ0��6�S� ?L '�2�C��#�K4��[��5��_";����1GI�م���=�G䇙�"t��!Z*��K�n����B�?F�p��g�i�ք��;=_"�p��߷s�^4K�'��J��y+`l�B��h+*!#�2ͅ$a�2L�a�R�Oi��Q�	��54P�6K�]�"���'$�����&	���f�E+W���H���:��I�p(!}��� �<�!�P�7VF����̈́e�J$!�"O�|�Dя0���c�MH
mx�����'A�8#�X9e؀���ɽ~����& ��,�"�Y\���D�|���r��O�}�u'�$\tt$�6^hNtI�"Oz�ؒI�a����qĄ��� ��I�~�Ȃ��en"�2[�Mr���Na�z1"O
���Ϣt���2��W�)v0B�"O�q�"�8N�<�E��jT���"O�܋u�D=A_F!Q$$	�!�LB�"OD��h�2��9��$�7E* P��"O�D���ܻ-� 仠cS>(f�Ӷ"O�5M���[�w#�|���"OZY�Ѯ�% �\}�>J��e��"OL]�"���gO��%�ıHʞ��"O���N�q�"��g �(w�J�ف"ON ����#�t���($����"O�Ar�ƊQ��m��i5� :�"O�� �͡@<����G^�Ȩ�"Ov��7�0s��I��U�R��D"Oz�`�B�;OG���A���ȩ�"OH�0�n] �@���]�f�:�2e"O4�����M�ܡ���+i ���"OV��rC�$T�&�QPL�4oH�Y�"OZ0�V�2arY�G*M	u r�1�"O��"���5���թX>�R��"Opp�c(L�$���KG��*��=�"O�i[r�'q����`���S���"O�5�P�7a
�B�/$���"O��P�������fݽ	;6}rR"O�]���+6���B�&T�t�w"Op���-J?@�P]j�"��n����q"O=h"h��a������R~Z��p"O�h��"��S&��Q�R�j��"O �%��P�Rd���>����$"O�9Q�/0nV���͏��j�"O�L��ɝ�7;p���T#R�	b"O�@�V'�%6�K2�O�$J�d"O84q2��	B\KFȏ�,�ؑ�3"O��y�Bި|��jT%a���c"O̤!S�	g����<:��p�"O2Q!�OT�{���)��Rg���u"O���2�3� r3H_� ��}""Onh K\VFtXs���$�t�:"O�z"��"5IL`�rb��f�J�"O��1 Y�9k�8"�k��2�Lҕ"O*���$ȡ@�X�����9q�Ա�"O��K��j��EhX"�-�e"O��H!.�)v[بwh��j&02Q"OJ�r'�D
@j�q����6 ���"O>��2��9D�dJe�0[B<`�"O�I�� 
8�Q�3n���Jyi�"O����������5ɀ5"O`�ר��]��آL�y����"O�1�R�[��0Ak�[���s"Op�2#-W�T�@D�%g���²"O�%9Ѝ4�9`1b8$,� RT"O$�I��,v�iZ�bD�:c>�"O�i[ 
&2b�g1BƘ��"O��ZD�ۢ^d`a� A,}�1�"O�u��E�n�"1{�/87����"O�PH�(�W,n�CM_.��S�"O*�����B�:U��!�T��"Oԁ��W�$&�9�5K�C�  �"ORe���y�
E*&��1�"O� 8M;A�ɵ)>&8��ɗ�$f-� "OZlbt�M�:��Au�[!
�Q�U"O��ɣ�\-V����?��q�"O�q��D�:>�8r3�E�m�eҒ"O�Ed��x�D��׹0 �L�G"OЩ�BKmhN����9$��l�w"O�Di7eU$7������8�z"O(�z�E�8|���C�={�4�"O�ĳ�jӰT��E� ,��V�:�"OjiSW���@z�H�"kO)��"O�l��W�Z2�<@F�a��U"O��ir�۪j�|i�#(ɶv:��� "OB�WH�S٘��FB(Ͳ!��"O�@Y���g@�Ct�H<o��M��"Oz�s���X�&�R�Ǝ�WFU�4"Oĭ���˟3�X���(J�8���s"O��Zb�ΩC�l���	B�Z���Bp"O~E��K�'1>����I2��%�W"O�p���7)z�cA	�al�"Obu����U2����B� A���"O�T�0��n�A�`�F�+�u2"O��@�����ִ{T�L�Dd.�+�"O�q�+6��5�ۏ7�l���"O~�Pgꆰ UHkB��6��q "Oz��R]�|s��;��͸%��58�"O �����+����5�ȣN ��V"O2��
�"YFN���e�x1�"O��A�,\&T��Q��ǃ] �`�G"Oڤ��S�.1*-��.`iA�"O�x/��P�@	'h	@�Ҵ@"O
��4�O��v�*2�؎x��cr"O����*�jE��  ^�b�"O���&(V-w~�����4^6@H�"O�Q:`޼3�� 1���L%F�R2"O13`�	l��I���<.6��"O}���ct����ӓn���"Or�K���5u�؋���,`��|��"O|�:Td��px�y�sJN��~���"OE �^&}�����|k�}n0�OԼ�d�!�M�ƌ��Sܸ����X�$ea��}�<��S'�vYq-�&��@���Ft�'5�iq�	�I�Q>-��ݐbP���Q"˚��$���>������4�]�U��*,;:�P�X�;��@���Y▹Ғ�PyM�n��?�'.A'I�~��GnU�`�U)!)y�L���οp�� '�H1�+��
���mZ#4�|qGe��h�7�.k�
A��e��p<�7aO�+��L�w	2xz��C�_y"��$��U��bL�T?A��bWs�Q�c���4A�8�3�AD�����A��9�dYOz�񶦋�@8�}i'l��t 8�(^��9l� X��;��\�H�,��I�7��n��DX��-	�:���aɢr����ǰ��B�Y���V/�f�ؕ���w��ɚ�- �l�
A
�j��~���k��#���������N|��s� ���OB�:RJʸ%4�AJ|��lU,OLh�
��@0�?B>M�'�J%
�B�"��)�)*O��S����R��F &�RYB���ٖ��|*ōH���~BE͈�3�x#g� -r�p�1Ð�v<h0��N���G�(�D�@NF�n�"�ΈR�f_5��I
G0L�A�̿j��飁ɒfʭ�'g��])\~<:��
{�\��p�����ɩ	Zp��OؘR����"���Х��R���15��!i��0걮�<9�4ʧc��UA�`ϫUbJ\�`ʚ�s|�5�	ÓyV &]8M>��
hz��5��M���c�E�Iq�����F8����* =��(��kF9`8.=@��!}ҭW�s�tXj�"3�Q>=0��0��� ���[��IG�&}��A`O�@��K�n�()��ə� Ӥ�0խOl?�,�N>9��>�@Q�/=��P��۝sO�qK�i�q�<!�"V5��i��G_�u�R�wg.B-fac�^lx��)� Nm�U�Sz��9@$�/Q�X��'�IP��0.��VƦ4x�O��;�b]�@��=r^�)�ȓQR^=!E�ȹkp��0D�1at@y�=	�2<������)�'a���qd�GlǢY���K&()�ȓ��(�*̘f�����s���q�،7�Ȅ�O d��Y���'Ry��P8a��TfPjU�$D���w��=���WUJreJ�%���乸3�#y�T���Z�fe���a�*	"@�)K�z�N�\-Ч�J�<Q��%W����q]�6��p�<a��.�%b�ӂ0Ŷԫ�Ky�,�O	��oޅ+)T<���� t�PK�@Wc�	`��VB�I�4�Jq�R�F���k���H�֕b�,T�L�:+��/=��$#"�@��!	�gW��&�_�:��~�펱�6�p�
Ѻ���Ė��l�@.F ���A	�� (^)R��2ғ���LϨ[.���wgN�Zi�G}�!����b	Ņ|��T�[0+x�L����m���`e#&%Bo8���d v*��0$Uu|�YЅg���{�M�'����S�>ͧ
AXMi��_z��I�7��a�nC$Jd(1@0�"lC䉌q����Aoãz�8��o�<<x�'�8mJ3I_x9f��Q�Q]�$���f��O�p��E<��ܫ(D'Xͤ�Z�(��B �K�	t)bVzYʬQ�ɛRf���g�e���'�ƀYF!�c�gy⅓�O��$�V�+F�C1�Y.��O<���H�l=r)���$bǋ'=��v�$q�����B-="r�@r�Ͻg��T�,��9�4�JA���2_�l�H�AT����^��ҧ��ω�$赙6� �<^e��H4��+�:B4&X=@!�St�:�W���w���L�1�'��Nb��A#��v��0�Ȑ�#֟L��uTḙ���҇K�b���'H��U��,V�4��@��S�H2�I)`��J��,m�R��=��=�<Ww䙂�mD�:i 8 -x��s`oT�o'��%���)�7��tI��<q� ���i�2��v S�,���dZ�C%�Yp���c,DQ��+,�	�7o��(5�TVe��|j��(�����H������4V����Xi!�DW�U�
ĩׄ�;C��+�����|��O���l�v���qO0I"ajC�8Mz�k�f�,��b�'T:Ur�
�5o�
Y�g�X�@���.[�Hl�Ve؟��hV��ȁ���8$���0��DaV��Ӈ��\��������d�f��JQ�AD>��W"O�9sGT�v��'��e��	�^�h�3(�V�*�I�>E��D�Q9 MI!˄��rY"��yB�[�.�j�4
�K�4U%P7`���'��9(��ˢj��ϸ'd�@q�A�,�<�Pa�G4J	��A	��f�XIf�T#y�z����&׺����A�&!B-��'�OX9ؠ�Py'A:i�}��0M<ax"eź��Y�W�|��
/G�nq9S���r����҅U��y���k�z���W.Ԕ��P���ɯ]0�9��)'EE@%8��8$/F�`ŦZ<!�D�'Fh�a ��7���H Q�m	!�d�h8��3,Gm�xc&�^ �!�$��ZHI+3N�3�6H)�ΰ#r!�d�.)�r�kq�2���9�d�(;�!��T�+�L4@��ϭ|���j��_%g�!�$-�.�4�H�h�C�kb!���$@~]ۣ+��b@l�+� O!��9R�<�z��	@�f�a��CM!�dJ:���"�M\�=K.4C�a
�J�!��Wˊ��B�۸1%@��o�="��E�!	�x��q��)T�hqA�'�XɆ�	�
f�)��
V� "K��&1��O�d�ީ�cg7D�\"�.�|Q%K�����E�]r����N+H�ұ���S�Ūc�ߊ���	SoP�-B�I?Y�����.��.ﰐ�`D����5k]�=�^Y�J��G��'�8��P�˰'���Zb��#V@��'ʄ]c��R�\��#Pk_�'��l���&��@����������Q�ʊP��x�(,{��{�J��b�<������ f��ACѲB;
����͏,�\4�"O^�I�8Z_.dQ��C��@�$�r���3.�H�(�	�&�7g��	S"�՟L<���"OF��7B߮2��ȱ�JG����h��D�x)��jc,\��1�g?Ѡ!%���5��$3w���g�\�<����D�@�����m�Q�b�ԟQ��T.~@��V�'_�!���.�Rщ��Tz>e��]�H�����=�?Qbl��idXE�4�����u*hFV�<��I��8��!� �6:	��w��Q�'&|��	�T�O��2��LMw�H����?�~�	�'|�8�J�p��S�����t��'oʈxЭ��P�4�3g	�{�(4��'��!i��ښu�r�c�F̐qF�)�	�'{�u1��*9)Xt���Ǯ`��=C	�'�d%:Um�y���j��*gT@k	�'���� a�eѼ�X�
ə"�^�8�'cte�+�4�.e�C��67"���'H2U{4/Qj[�؈�)�)	��'��|i�A�+)���Q�.����`�'^R�j%�
�Qo"!��@ `,���'<�]k˔1)x�Zr(JcDi
�'��ّo��dq��ȑ�z	t��'��5��
�0��Ȇ~�q�'O��J� ɦ>_$����B6Fk�(
�'�R刵��X��`���G�>R�(p	�'�a8ŪS��b�#8\���'Ռ�DB�w\I{�Z�+P�m[�'�F�资Ƭx�T�i�Z),w��	�'��a�Q钨-��Ĉ�R� � 5�	�'p�������C
X�d]�U��	�'�X�$Z6o��pb�z�>�'��a��'�$�����A�t>���'�F��Ӎ)�h@S�&�&o�B�k�'�ڸ�6����M
7�
o�09*�'����B̉�R�c�y���ʥiZ�<� lW+w���(A
X��dd�0�H}�<!���)n� =x�5L��C�z�<y���s��p�EKь���(��<AGʌ�Z��8�!�.&�~�#@N��8]M�@fP � t���!M%�"T�Z�f��-�H�3T��5j�riS��O��	���c�>`j�ѩo&H�r�'D^��!�Ly'��N�	`�h1#�a�>
#H�3�֚���j1�V�B�� ��>1��$K>Y��8#����ȋ'@5x\K�%zOڅ;J�Z?���XKa�d�E�33xM�eđ.��|;p�S, �^ 2#�O�p��Ǜk�`�~n:���,7��6�R�7�����Ô�~�e�4���hO�)�t�pk�:i�BI��!�!�$�f�h�q7��}�0 ��� ��t�牰]�<�XvkN7T� ��Tm#{2VB�	�0x�/�5��Q�Է1P�ɗ1�`��?E��E^�5spS��21Q�m
&���]�Gy
ç_� ����E�ih���ǈ��>���)�� ;���*5�*߼�B0�3t�'T�#=�~'`�@�iG�׊�ur��:�HO���ޞ;^*43D���)1�E�%Jشc�hYq�)�� ���ABκkL^��� ��}�'֚�Dy����f�tݨW��8#��`Pa�G�_��b�'�x��5��4,%|xc선Cp=��'�24Q!KP�8��%�*L�]���ÓY� ���g�g�e,fJ�q1 �`��z� �L���<��S$�Ф�T�ȩ����@��d.�I�.�M$��X�g�S�T����2F%�:$�d�jv�R���'�f�bf��0|�2䅂OVԺ�)��M�;��n��[��MP��H�y�ç���9���^#Z��0�ܮ`�XY�C�܄�%������\����Ο�<cˌ:G��Ro���$\����1�ά{��<�k�%<`ax��aT\��W���t����,E��y
� ,db��֝y�X��"�ޜ3��h�"O�pf�'l�h��X�r�l�"O�{eL>ks 9z�m�e~�Y��"O�)�Ƌ5M-����o��aA6q��"O�[r�[,'��i��	�Jy+p"OޅB)�6R�&�	�/M�c�^Uۃ"O�x)�K�%g
t����';���xD"O�59�C�(x��+��	l%"O|�3�F��k,�2g�C#�^� �"Oz��$�q5Du��꒙㒍�A"O^���ņ���D����o٤���"O(I[��1�j����-W�Z���"O��b�ETh7$q)�%�pX�c"O>ḁ�c��s��] �m�"O9I��}w.����eI
gk��y2��Q��2�(�qhe���[	�yBh�!a�1ڕcC�$z�,��O�y"jϧ�t�	0��@���F��9�yr� �
B�S�� ��%*&��yrh��p]��	�cU4�8yDa�y"`�/P�2��X9:_� �d���y�Ɖ�j��M�UE�.�$�`č�6�ybE��<�u&Z����4��
	�'4����/Ò{G:�q)��0�X�*�'t�e�œ;�n����
T<�ʓp���p@��w��x�\�:�����NƜ���!k*�4�4I����ȓV���P�T�5�p�.W;��ه���]�RC�jj\0��,��|��}��3���:�j!���G�1l%��w,��qi�:`N9:�)Ϟ`Zr��ȓ�f�$�l��	�pbL1p愡���,tKQ����	q������1�0$�� ��$�PX���P�uH�ȓ)�JI��E�I(�)����6=��P�ȓVcQ`��B�vz����Ol%B��ȓ@�X0 u���b�I�N�)O��ȓh��]���
�|�H���ja��7.����e�	  �<p��t���ȓZ�EQ4"�)?����+Z���ȓd�Rq�rD�	}�n��p�ڳ�⍄�/z�AJ�l��{��,/�X����'�!c2Q��'F�V���ȓx�b1��n��x��d���ȓ(���IT��6���{��� �VY��|5����+]����{��Ѕȓ�!�b'jm:���mG	E����5���2"
T��2����$JT�ȓe���{u!�~V�$,�('|̆ȓ@+�Y�� �<�d��G��>s�0��ȓ"nty�F�L 8q�U-;(���ȓy�X�RAI/M/�4����5v^��p��C"����0���Ͳ�ń�j��wC	�}�ZLb%�1�M�ȓ0�D�`FэVt��[���7U����_�bi{��B'H�@���ۆ	��F{D"�A$z����.G��ԇȓ' �<:f��8%Θa3w���p6�مȓl�&����A�:���j��G�kU��ȓ jn���CD1k"�dp��, ��L��h!���'�tp)�RD���@���M<s߆0���_֢��B :�+��K�TV})6i����ȓ]�.��)I� B�Y�$'�D��S�? ���"/Y O8��ce�Mp!D"O>iS�GِC��\a��1c��q*f"O&�2L� �j�ecǼ<N^��"OxE�S
� f�� ��K�[��H'"O UإIj����t#X�D�THT"O�<�	�.���M��r��"O�=ȗF��"��HP�}ɪ5�"O�0`ue!)�I6FX(�d $"OB���S'x2¨i�d����%[F"On��0F�O[J�17��-9�Lic"O�S#�2rq�e�e�l�tA�"O�([�N�� b��R�Yp"OFEꗌ�#��	���@�z6�K�"O����H��T�nȠ�
�"���"O��i/Ճ!�������@P�"O�a3tJ&��y�j��>8hW"O�2槇�f���#(�5=>��*r"Oq3EEP%��,@�O�/b�u"O����F*8�m�p�:K�;�y�N ;��<b�;`�la �Ā�y�m1!��� �i��u��i��yR�͑)q�q��B9[QN�	���y�ʑ�wS,iQ� V5)Ci(D��y���P�Ҕ�2$Yx$P83sa��y���+�,x*B�ۇB�ά3o]��yR�.E�޹�W�� E��!�NA�yR�2?��Ly�\���p��$�y����XS����M�zM��ѠQ�y���*|� ��pL�
r�ɥ�B��y�+�xz0�P%�7s-�8(E /�y��#}Lv����'9R$�K+���y��(�Q�64R�z�M[&�y�^<Ly�P'L (F$�2� "�y�i�)ĴLs*\:M�.1a�-�y!�
M(Y�fH.A�D���m���y�ʀx�*�z&��<@����y/Q��lD��ݘ4������y��Ӿ�(���	�%0���3u�G��y"���:���Acm��,�l��agB��y�d9 �es�Ȇ�-��	a�ʯ�yrb[�e�oT'xφ�)� �<�y�*��<�p,��D�r�:m�E�ܧ�y�b�Y�f���(P�|x�` ���y2	����S�V�{�Hp�rM�>�yRF�}�t��0��zan�bR��y���?�F�	g�K�I����G^��y���^�DK>�>�#���y�MBJ,�!:-vL��0LX�y�[� �
,r��ъZ]�E����y�h� y<�f䂡WJ���Z�y���u���A'U�Q������y��3�hhP��ёutFU{�� ��y�`����E{'�&v�:a(�Ý+�y�N�P>���:`�\ja	)�y����U��z�֮IL1
�AT��y�錮;��`�׎�<���)�cF��y���:CZ*q3��1��%C��W��y��!p`�`Ԏ�?at}��	!�y2/��$�F<ӎ�0�z�a�/�y��͇jp�1��>b8�*���y!�(K+�iQG��`j��,Ÿ�y�V:D�U�!צo�~q�@�H��y��؅vш)
�mH�s]�� ���yBIڮǖ���;Z�� ɗ���y
� \T��"�4h��#���d����"O�9ɦ�^)o�Uk��]�Rq3D"O���q��"
*�\H��C�艡�"O�԰��֚fD<5*�+ׅ����"O�e��
�iԼ��g�E3e�JQ��"O�)��#��1&]j�ɱqg���E"O�<�R�>-�h� �E�3 y{�"O41�S&s�(X���|n!��"O�@E��p���@�ɸGI0��c"O`h��ŔQ>|��4c�&89͈G"ODI"a�M�1%R�b�?P�F"O>-ׇ�����Ѷm�b�s"O�T�uC]<�����@R�(~�U��"O��XT¬4*B]��*�8B���R"OjP�G-ھq�~�h4
�PNMK�"O@eɓ�-R2��BN�1D�)"O-�k�o��	�%-��)-�Y�"OR�[���/$���٣�( &E(�"O~샤AǑWX�J��3# ͊�"O�`9�`H2RрY��T��]{�"OPk� �d��AbҊ��U�6�0�"Or��Q(�%C��񩒦R�2�[`"O����6�̄�PU+x`"O�){��϶e_��[%��&�88�A"Oti��.\!|� ���/	'vj(U�'"O�2�H53��U& C9Z�t)G"ON�9R�T�Z���2���*9f��0�"O�E�Rb�0!�6��t�848�#�"O����FT"�����C(�b�"Ot�yRCM%4O� 3r�L<]�֬�#"OɃ!�֔/����u�C�x}b��"O��YsMް�F��R��b^>�C"OT�֍�N"�sp��cṔ��"Oj ��Y�xlC���R:��7"O�dұ�`2l�����T)2�g"Oc �J�Ri
��N�)�\�"Oj,i�aU=@\L}ڤ�ִ*��kt"O䑀���5='����P
`�8�"OX���� y�\+�K̑p�Ha��"OЅ��A��j�� �ՠ�/ty1�V"On�tfC7~-R�1UE׆x��S�"O ���NC!θi�w$� l�]�"OT��FF[n�)�B�LR><��"O��9�0�&ѓ�W$?hL� "O^ �%C�%&�4��U�`]2�f"Od��D(�+chrE���r����"O��*�C� �r�y�o���!��"OjL�و3P~�Z��ӽ<�^�!"Ol�˴"w��`PP�@>��J!"O��2U�əu�`�Ȇ��L��)"c"O�UYa��`��	�����Ԓ"Oʤ��	[b �a��!L)4
D�"O�����b��]"��Q1d(H� '"O��g�C�`��# ��,Ȁe"OR�х�>M �(�8Kzƴ��"OT��ѧi���� Ot�l�%"ONm��B�V�"g���sd���"O�@27h�0;�B���rZ^]cV"OZܘ��*,"� �0(Z �9�"O�U�t��'����6 �4iZc"O�쑢bڶ+f�J�ۚrD9�"O����c5` ��.�.��-×"O���`O�,��}y҂��0��Р�"O`�hD�~����U��#.�0ěR"O� ��R].^��r��=o���"OPq�5�pp2a�@��O"��"O��P=#Xjm��M;pFza�V"OҴ3�	   ��     �  �    6'  `1  �7  �=  /D  sJ  �P  �V  ;]  c  �i  p  Hv  �|  ͂  �  S�  ��  ٛ  H�  ��  �  ��  $�  h�  ��  ��  ��  ��  ��  *�  v�   Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�� |d��"O
`�(�;���8���-0��1%"Oj4��ND^[��"3/9�0|H�"OB���H��*�ʞRy=a"O�味V�!X��!&F�:J�$���"O,��a
���C�Ą�M�"O,$3%o�-���p���+Ն�:1"O��ݢ1����`���y14]2��i�<�6��{_���c�H�`�fX�$Kn�<��A̼VI�xR[�)�Ć�pඤ�ȓA5��('nߡ4�� �)˩%� ���,��r�؊b#`T�eT09���ȓ!�b��g��}�8�F��-? �ȓ
K|m�ș�VṔ���2�%�ȓ"R�X�j�4JN�1�˘X�i����̹	_�jZ��1!g��zܶ��ȓgil,*�J�
j�Ne��i�J%b���f	�(U��:���G��$Y^م�~r�� S�%T"���k\�jx�ȓ|4�1�îJb��@ӵ�ݩn�V��/[`�"�v4�R�!ʎ<��M�ȓ`:��z�ؚh�J�Z��$HY:	��H��p�m�C1��!��B:��0��EnjZA V;9����J[
2���	��4'J�EA�IVW&��~�(aZ��ӹ�>� o�Y�|�ȓ�f�A�
Ο7�H��M�$�����mޠP����/���ANXo*�ȓTv�����{ ��-7�*h��I��sB�8�8���3����ȓNe*M�悡;������X�o��!�ȓ'lj�#F�m�+R&;�|��2)n�C��0S4���T:
b���:�0!��e֊��)��ͷV��,�ȓ0�&�8#���� ع�L�����;�P�AFd���,w�6�F{��'O��V���&�;�+0:��x	�'%��"J�[�]�R�K2r��"
�'Oe#W烹�R}aC��z��
�'��;��7�������L	�'�:<*b&K"4����M����9	�'نx!c̓>�D �,ݻ2zX�R�'��@ �F�9<�m�7I�"+�a�'ր����>��Y�
�%&���'��0��3L�r5��M/� HJ�'U����J08fx����I$p:<����Ojb�X��tO��S��Y��X��%~!*C�I*(��(�g��j�:����ݩ
��B�9�p��v�Yz�<h�$��f��C�	6�@	�6G�v9&�PF��S��˓,:^�<я�d>##
) ��V5� �R�m��%�!�d�#o���V#7���Y,*�<i�����5-�(ء�͉�F�6M�ȓI5ļ��-��wX��q���!�Y��.�*Q�%K�BǮL	�-�5
�M�ȓQ�6�N�~�H�@MX�$�����a�,�u�H<8�@bf'Sh�4�'�bloڢ�����{��6���8�`ƮS0V��$B���x2�'��1I��.���TD�I�.���yb�'���"M�1��y��χ�Q���!���6�IO���$a��v��I�<��EJԧ�y�l�PA��!�܄F��t�����y
�  4i�Ώ�B�iW��g@��"O�ɨ�f�;e$M�g�(FPhv"O>�+3���!�>i�!�Y h��k&"O�;JU��ʴ�S��b?:���"Od��#[?c�a��DV�X/8a"OvuC�`[ &��%+�#�,=8@�#4�X!-�cN�\2��O�;mV�C�$4D����g�fA��"r�p  krg2D����W�(H1��˕�ԀCq�<D���JӋ{j��h�M�u���[&�9D��ӷB_�\�@��]aA���-��0<�0�S��h+���5`�`�+f�p���'��vtH�!�~UCR-,M��d��"O��]e�=c���4$�2��CT@�<��K}aU�DCT�r�H�`���ȓ^ю���ħ�p8�%�G[Е�'C�'>ўʧv��Q�gdM�zW��۱kѾ���|y�D�.%�Jy1��>}X��
��y�N���҆��3y;���dZ?�y��,q|�j�BvH\�p�B	 �y��	z�0�V�S�I�m�P��4�y2��1���� �%}�L,���yR�Z��!XEg#v������D(�?��y��)�Fl�4N�앸�d@	�h@!ϛS�<yb��7قr�
�x%���R�<	0oѰ	�D��7m\� (�BLK�<��K]��B�Xb̝�n`�z��^�<I+�|f�D7%��zc�_x�4Dx��R��mH�b�8`�44��dHD�<qC{)L�K�
����we�f?	V<O�㞤(��雥kU�D�4.�gR�xI��"�!���g�k&��)�4��OWsr�	U?�g%#<O��#E�ژ0��%b���5BQ�Lb �	\�����P� �����i�v��PZ�a�!��~ߨ�z3k�[���J���/Z�a{B��b�ެy��ԋil�Y�V�!��]��X���UWL,j!o���F�<q��>�"n\F>�qE |#�<�"^�<�pb��
������Y.��!���ܦ�f�'�d�#�)D;�>�z`DI�r<�P8�'�b�R��,sιy '��|��܁
�'G����ݬ=�t`���u�P�
�'��E�`�-(�ݐ4�Y�knhPj	�'VD����	�cGf�k����'�h�nZ�����v��f/��c�'�l1�QkV�e�@m�f�'l�X��'X�m��B�%�l����U�R�&���'zT`u�j�H�7�` p	�'S�U�F�U1Q�A�5"E�E2	�'��y��F+W�X9{H�����'=xم&ǁYi���qJ�"�3'�!��"������p�r���^�!��c�L)�a�Z�����.E�!�ė�d���%r^�Z?M�Ԭ���/D�(!��M�fdQ�u�U�*7�8�N9D� ����8�}B0S���0*P�7D�dӥ�����[���Y��J�N4D�x����+YN���!J0���	1D���g̒7n�\�C��P�o��h��-D��1Ð:�
Zp̈́6�Τ�wl?D���"AK&�ܑ��@U�fN�yrG D�R$#��n�>���S)�p��h!D�HQ�L�J¼\�����hP~���.>D��j D�G�^(��6-���7D�� ��j�DE�����*���z���"O<P� ��|���%4�b2�"O|�p&&�"�����EE��b�RA"OX�Kg%F�;(^ RR��� ��A"OI����d����!.��.īf"O
d�C�e�}{�R>"�}�"OF��g�L�6�BT)�Xe#���s"O��0���Yhj�����!
�"OL��ov����_���	�"O�m��OYn���E�(RX %F"O���'!�-D��4���>gQb-Q"O���'Ń�d���[���q����"O��q�A��:��p$<D����"O���T ��sJ^h�I	#!^���"O�h���ז�hI�燐%V��"O  �7F��1l��;��X�[�$Y[�"O$p�1d�]�S�F�%L�����"O&�!*œY�z��� .D��\�#"O��xפ�	t�A�S%OمT�bo!�dļ���	�/j�]�5�N�.b!�$@Z::��B@3�lYʲ�ܤGY!�d�j2�ϊP[d��D\6@!�]
��J�hV�o`����]�!�D��NL|�K�-�-�(�)����!�DF�r*���4���
�.���!�n�8���C,�Dx�F�L!a�!�䔻5?@\˲	/p�d���,N7�!�$J0T�  ��̵}3r�"�;�!��X�)2���--��+�+�)_q!��?�l�`�I	�?3��ӅK� �!�Җ U>Q��`��iK���*�>�!�d��hQOX9`�4�;ŧ�>�!�$O�dn��h�,kk �,��N�!򄀾M�p�ֲ8�0��v��6�!�ׂBl�s���4Y9��5��4n!��J�����V�K���S���`3!�D�&��[���!zǞ��� A77!�D7R�-$Dv�����/]�:�!�J�1���	RZ���� �!��:{l�`�v�&&�*�x���h�!�A&j��D2!�N�y�:�ⷩ�%�!򄋩^�����FF�b��@�'��O!�D�;k&0P2iV+6$�y���j�!��F�/4��y�� �t����:A�!�D�P@�0ZDn�������".�!�$�5j��hF���!�������r!��<���{q�� ���8t�C6X!�D5<� <�fDT:Mf���"�!{8!�D�M�9)�ό'"�t���W�!�� %�E�b�ڢߎmZf"Ĉ5!����PX����oe�h)2�|���'`�1�r���yxك����l+�'�x3%� 3�(g
���� �'8v��@�4?����l��8�Ű���B�U�y�!��#���M?D�$�3�G�\�*	q�bSg��:�l>D�ԣ��H� �왑��M����TI<D�LA6+N�x��da�eK("K<��Ql8D�(�0�ߎ{��q����|��2$2D�4A��4�P�
w���l��d�U!4D�|�'�^�h��w�+"͊Q�F8D��#V�1CS�h�G�-4��y�a6D�\���,F̈́�����1l�����,0D����ɄT�B���37;��C$e8D�� ��J�N	A��T�E� ;�ԙ��"O�(*wOִ�����^�:��t��"O�	ڔ �9&�^ܑѯ�9>��U@"O�m��/P�O�T�b�m�'W�\P�v"OŁԌ��F@lu�Um�5~xq��'��I�h�	ꟼ�	ٟ��	ן��	8����D�,3��_~���	��|��ڟP���L���������I5ߨp��G�eȥaã�>l\���ş��Iٟ��I̟��ϟ��I��0�	�-L��G��4���˂F�8Q�����ݟ��	����IΟ�������	����	b��Agė�!���P��U.�e������I�H��矨�	ݟp�IןL�I�T� �Q��Y�;��9���9�����ٟ��I埈��ߟ�����`�I���I�[��ը��N%-���3Q�"������I��4��џ<���@����,�	k����/_{p��I4n'\J�����`�	ߟd��ߟ���ğ������	.p�fi �M��ئ�k����w2r5�I��|��ş���⟀�	�l�	ڟ�ɺ	Y�Q�'N����� ��$�I��ҟ\�����I�8�	ǟ��	ߟ`�Ie2}9Q
@>9x$	��K�x�	؟�I�I֟�������؟P���:_X�m��xQ0PX)����?���?)���?���?���?���8���R���R��%蕅��h%��3���?���?����?����?��ir�'WJ�j�GɄd���iV0��6��<������rܴ1��b�oǰY�|, g$F�njq�r �h~��lӸ��s�L�ɷ3�Ƅ���BH(���Z�j��}�	ퟰ�wD�,l���T!�Z�O�L�rmF�Z{Z�iP�GD�x�yB�'�u�O���0�\0P���	O&����u�F�sU�=���M�;k� L��hɏC�.tcD�� �������?��'��)�>�4 'gr��q��x	���_蕺R�}�8�}�i�����'Grt�%̈́7)(�/�7j^0�'Y�I~򉞤M� ^Y�F���	�N���('gŴg��i�rH�>����?��'8�	&EĈ�Q�J��(�HP��g@�
��?94��8��|:$��O:����}�ys�#��v���d#�,z��<q)O�˓�?E��'#����aT��@�a Ó)@�0��'?7-(*�ɚ�M��O֠���]g�h�c���4�b���'���'��Q\0����O��"�/3 ���J�L۴7�P���$1A���Q2L��$�+|�ˏ�L>�A-�\=���͑(m�p���|�<�����ΐ�V��c��EH6K��H��Ȕ`G�͚� R�R(�4tJ�/�֜�7٣w7Xe��M8W�ܨ��*��z� hHK4 � ��%&4պ�	����R�h����<"Mj1�,��VƐ��@>�p��'((��Y��ʇ�!���o�7-�x]"�`�hC��������'����'IR�'o�t�2?)�#��co�`�iʯ#"�1�y}b�'��9i��D��D�O 9J��7/*�X��.��%ps����J�D���M+���?1���rA�x�O
�-#�#>^����YGpF��nt���y�'�	�?c�����t4��\"�895�¦r�́�4�?I���?�ܣE����d�'��mT:a~�<+&��U{�J�_I�6��O�$�O�k���]��'bB�'1��Jc�`���
�<R(�!�D.'�6m�O-XDG�e����n�i�)1b��9\�R��CL>*s�)5�{Ӹ��K;X��D�O��d�O��d�|��-
p�)I݁�8x��f�~�P!��˙N��'���'���|��'2I��툿Nc��vGA(�|@��Y��'���'�"V��2������ 8W���C���v�ިI �N9���?QJ>����?����D}��ڵd[DlP��
m=Ҝ�������O��$�OZʓK��da���d-e��8�-�>h��rGNA�K�2�?A����?�#�U��i!G�
-�V0I�оW�)� ls����O�ʓr�z�k��$�'��T�[?#Sz�h M�� .䋥j]�/� O�d�O4 ���O����OB�OnZ������RCK�>���;ܴ�?��;��=x��i�막?���|�ɏLډΒ�p��,gf�HASX����[:� �?��g�I��Bݚ�f�!��DR�d�]6�6MK/h^Dn�4��̟x������|��Ґ$F�PW&F.+��µJ;~y��"4���'���'��^>�OH��voܜ�̀��6kD�qӾ���O��DN�@���S�4�>�v�U�ȴ�!2*���L�A�Rc��ן [a\d��?��'�2����C�"L�	��ZGD�J�4�?��I����Wb����܌[.$�;�"ۚ:4�a�'-�qn� P�H�f��l����'�)�4-ǯm��P���9lVY��U�L;tO����Or���<I��?I���.k��U@5�ӖY��0k`
�e��������O����O��D���:���B�����츖�3~}R�Z����埔��ryB�'�r��_�R.��:���օ�Z�ͳO$���?Q���?q-O��x�+`�#w���vJ��+��EI���,^=rQ�4�?����OJ�I&����3��UXi�&�ДE�Tt����M���?�*O0��N�M�S��p�s��&��`��w�:��b��rӆ��?i�b��Tb������q�? ��p��#���BJt��@À�x"�J��=��	!G�bpp�	҃/���(Q�I�lo�B䉙b[�4
_�_r�iT"CAގ�Ife��8A�)[��E�H9
T��lJ�rz�*RǛ�w"$)� F]��T��f�+ٮ=�E)I/a�찻�H�HL*`�jԞj�JD��L�%��x!�% ��]	�,B9u��sJ�TtZ��Pi�-���E�B}p��|`�@ Q��`$�i�r�S�)�	ʟx���^w�R�'���.`
lM��mK�c.4��M(6�0H{�G�,�R)����D�ɖTS4����D�����2x#��p6��KR,��~� (#�GéC#L�SI�'���˖&���&	1�_��,��A�'aL���'c�7�Ħ��<�����$�9>�❫���h��y�mB4!�d��4�p�����s�Dd�pL�/&��Dz���G�_�`��؅�u�\��\�ˠL:@BRQ�`)F	V���'�"�'��D��'�"?���X�m�A��qr�+$V<R���;����
��4C��M��p<I���4!F8$#Ѯ }������ę'B|��Ʉ`P�5�t/�8���'m��'����ǜ=���PB [&>4���Ib�'��
Cl�b�,=෤��(%4Q�'H��� -[�:q*F���
FHY�'�6��O�˓g�z<j��?����	O�(�Җ��e�X�����E	�O����Or<8CM.�r�s��S�)��	�|�ƣ,_/j�S�O$xoP� &Dj�'/�(��A�5O[�PR���Ao���1����Ն�k�`Y:1d� 2(E�V#R\�'4 �)��}��6ai�����|W�Đ^�H��^j�*����?����9O��V�f�h��撳E��P�'h�7Mɦ�IDx�*�ʙ0i�d��r��2#��?�����<I��id���L��\��!�{�<	�-GyC����H�	z84���v�<9��T�5ꫠ�9,\>D�g���!�D�"�yy`� 	J����%
�!��#QYb�q���h?vp��#:!�D�7Nz�����K0P7�ف3� �oQ!��P�]����G	�K9����'\q�!�R�-�t` .]F�<5�DfU-�!�$V�f�J�s��A�ltAjTc�!RO!��'?̬��G�7M!��O�R:!�dC�5��#��9�V��qo�69!��)H` �� �z�H�� D�!��A�Zlȃ��J
}�䣓�w�!��6]��z�(e%�"�[�����ȓθuSQ�M�U\N��fN�b��ȓ,��`�M>�V)�DI �M�؍�ȓ��Y�cЮ"�2\Y��э�%�5D�@�N K#`ʥ+�{�L��8D�\�&�W U|���<��#�7D�z
��Q ��}��yԆ Y��B�I	F�e����2"�蔠�N�sB��lh�wΙ�/jH�v*Ɋv��C�I�d.HhR�ơ�!�U��� B䉗@�d�x��P$���A�NG*�>C�	M��DE��ZVr�0�f)0� C�m�p�G땴a�%��Q4A�B�Im0.�P�
g�f���Os��B�&lb�Xñ�ܼ /���@AAòB��c^�R%�:��٘�(�LpvB�	-i�{w�XC�I�V"a�B�	�Q�9�Y����s��A��B�	�5☠�DըH�j�����Hi�B�	Z<�Bf̙	�~$)$�S`�B䉟n��m	�/ɘW݈�`銈A��B�I�Y��2�(�1e��.E'f\P���	7Taf6͙5��1cNS �-Rc@�'W!�+j��)!�Ӯ/p�z��Q#`���rAOe�Q>)��M620��%� p��H�N1D��1aK]%]���R�[+��!�Pam�T��g��qO?A�  �ip��q�^�ZUc�F'D�d��kڪ`^��˶�ӽ$�0Q#�c*?��e�;�h����(Tr�B��s$��uB��(�xr)\�X���)"�33Bu�? �)!$�U�<�@�`�$H!PТ�2�nQR�ǃlX�x��쓁x2xa�!G��b;T�P�F$?��K� Ev�z��(oؒ|1GO�?a%J,�-�5J^"͂��� !D�<P3��)8j��q���r�aCa�#u�����*�,g^��O�'{���ǎ����čP�=�I˃�C�=�u��Hz<���@�hp���5�Ҋ)lT�5�^�'�X�)  <림 ^<<fUDy��Ɠ0��i��+ϴ{�n� k��0<�3F���ܡs�8CP��t�Q��
�X��5&R� �d��+�~�y� �e��Pa&M8�O�ĢW ��0J�#Չ[	,�Z� ֕���C��R��Z�˧84�!�s�4��� ��P�~:�0��� > �I�"OlPiuC	��P(�
�
%����7�v�����	+J+
$��8���l�-�<1� B�'F���O���8C9d���­-h��`�!<H�I�;���{�	�*��c �,�Q��� N�� ��nQ@���5OBiz��m\�q�*�lm��{'�)�`�R̔�o�`8���S$}�����I�hEL��
�Q���3�IL9yM����R�qX���'r���!$��Nc�ɻ#��(����=�'|HN���^6J|>�znչ ժ�ȓ&ʂ��u�NC��P�C@�-FYj�$:�n%2��7�)�KP�D�FX�;�F�� e�`)�;�
T%X",��Z}F�۵��,�x��WoؚUMx�Y��Ih~B�ƀUk��߳;�1Z��O�'�4�����U�z��$H��5鴠�Ó7��� У�$���B�j,5�T
����Y �SCD�+Ԉ�� i[%���E�8$��	�?;��rFABi�Xq#gή#���H��a�.O`��ǉ���I޼�x�ӑ0Y�5$��O6��䌁9��C�	02������8 iJ�¬�8� ��}�F KS�0&������Z��gy���`�-.���O)b����%�'?����[s#��x� Ưj�@�9%�<hּE37Jɫw�b��B�|���i ���`�\@A��37�M���N�E[h�"�����n�@d�ˢG*b ���V���� [�<P!\O�%���$AK� & ͭZ,#@]�X6/A�qO��)G���2&Q�mՖ��㨀�+\= �B���`�'�4�91�Һ@g>$r򅚬T�����S�,�	p�s��Ha�.!&4���?%p��j���	-��帴��P[QL@?Jl��������Y`���� �ȒD%A�W@���Q(���UN�j���4���{�d3�	 (�ع�Ć�%g�~���J��+\6#?��vl.8��i(��m �MKנ�cx�(�6�CD�4��7�����+�f���ӤlO&-��M���I��ce�>��d�'G5I���+#��hP�/�v?��',�dO�$�|͂�E��h*=C1�ډ5o(B�I3 �z���D�S�h��m�, �
5���;I�@�9�'�����	�`���E��sb�B���ۄ���M% ��|؟X��̊�S�=0���W'd
����T��'��$�6�^��V�ڴ2�����ũFqO<��ы�)\ތ�b��8�L5�0�I��L��bL+0u�Ca���)�D7��
��u�.��\L����
a��`�d�L7m`"������p=If�M�%A�&W�@� ��c}� �(R`6�� J@&p<$1�b���~��O����Tѳq�˽[
NT2��#Gt���9Έ�s3�4L��H��
�S�h�o?�Fᒂ! �<�s�'��?I��i�4�b�w%YS�%Ȧ&\���[9Zp�0�'�XQ"e�/93�q�Vg�0~�:С���_���d�>b:ѣ� �����)��O&�HԤ�b�|,�fݩ	
�` E�'ͬ��k�vkNLRt	:�Z%h6��V{�!;m�"A��q��b�o��Z���B�'.�CH��Vet�s_W��hSc>?)���&���ծ�W�x�# �UK��?�xU �^�
�!M]-ft� �P;D��$dҘc�Z�SK@Ov���G�	�&�;r��y5�ʧh읙�I�Ƽke���� �� �5�*���J^<ia��/nd0��w�[��	��=nDa�Or��:\,�����]z.}Bd�Ė�m)�M��ķA�6ii��I�z\ax�e´W����A[�n�:��fCܖT\�1H��
�\��ŪBcC�%(���-�X�����H�j��{��<EڀMQ)�����V�R�'����!J�M?�Z�"l¢P>و�iF�`X��h�#�bå^7M�t�b�R��y�XQ�$�އU%$D�hŸ�y�� %��|n��(���.�7v0�g}�O�v+��>-@��KE�]�b+�	a�'Nh|�a��>V�� hаr���x�O��uI���p=�ĭW�q���@��x3EBb���҆�צ!넯� ���7Nڨ�¡�A�.D�� %�BZ�"�a�f�s"O6%�F��0~��0MV�H-�m�"O�l�ԡ����3"2@dq�"O8��3"�;$\�1Њ�r4�S"OpYhc�׆eA���e��6`����"O  !�i���Wj�4~tNq�"O483H`�؁�Щ�[��)�"O�����E�k���%\0EU��Q�"OV�!u��,��dS�ҐBDb䠔"O���U�E��T��O�C��=�P"O�P ����<�҇u�.m��"O<	�p�ȶ�@t`c'� ���d"O��z��
#�: rL9��{2"O2�@P�"f�З�ñro�hZQ"OT 9%�E�I��i�.�Ni֥sA"O�A���B$�$��\��"OrQ�D4VV� !O�`M�"O��Q� f�H$�%Â���̉�"OJ}�Da�w��5J���-<<��8�"O���H��
��]8=�*}�"O��Ye靓>��]($ ����"OMDЖ1�ݚ�"X>eٌd��"ODl@捌1(� u��&�;�����"O ��Rf�J �qc^5k�H�"O�$ç$L7<e1��W�|Y0"O ��N
���q�!Tp�$�у"OJة �N �
��CZ'_���� "O�L�`��)��
a�CC�Nm3"ONs7���0:�A��)<��b"O�Tc�$H_۠���
�/&퀳"O��r�
y��ъu�ˢ<�UIw"O��)� K;N�\���ӞH��P"O�@�ˤd<n��P��D���u"O>uP�g� GWHy۶ W6�Z�+�"O�D�4ޡb��85���T��i"G"OU�EG���.!3�%}��["O�"�`'D��YG��P����"O�E/M�+Xa`M[?fY��g"O<�H�ŧ*|M�W�U:E�\;R"O��Bb�֡DIg���"O�MP�a��K �'JjQ`�"O����mU�_�l�ꃥ�[-��Q"O��wo(qxN�R�ƽnq(<�"O�����(���CM<<	~�x"O6�S�?9��j���3`�^��"O�p��]���Z�x�t�����yb�Ш�Uȇ˙.n&,�DM�y�G ���h�eբYM�Q�E/�y2 9(q�m�ס�Q�)Xg�Ѧ�ybaFjk��#gK�&�pYC�%�y��υ8J����irv�9f�L3�y�Ĥ$gU���N���̮�yBOH�wv
� 4O���VX Ǜ�y�n�\��!m�>4�YH�KJ/�ybÙ��t�DG:��y�u#M,�y �$(?��"7C�=`��Q6�	��yr-�< ���F�A=m�� �1�y2-)���Ѐ���Y�P]�T�͹�y� ��QTA`!O2�J���y2H�.�����_�A�L\{�$
��y2@�.�8�{2"L�<@H�[Ff���yBg^	-܌��>3��2�
C��yb�P�]vM�@��7�V�rr����y���pk���DZ-*�^)���)�y
� �8')K�r}9�#�0~��w"O
\��dѶǢXp�Cؒ2ϔ�Cd"O��2�AX@�"�q���P5"O������:FA͹�Kji����"O^E�pO��qÀ��<�H,b�"OD� E��"���*؞|K�!�"O��C.R�D����zӴ�{�"O�)Fnп+9�\*�M*E�ܸ21"O�Hj2�J��@M�,Fb|2���"OĤ�1ℽU`�-(q�@E���T"O��H�(�Yk8���`a֠�t"OΕ���Z[c�ܩ@��Bi���"O�QR��H����m�)#�ؘ��"O����eCD�\}V��4"ON ��M� 	���D&�/a�+7"O�|bb���S�p��d'�,��C"O:ܪa��$�\}x�M�<3���cs"OB�3t-�EuD�ꆭA2�:���"O�e���H�2�ӋT('��,�"O	s7��L!��a�Q�<aK0"O��FO_�*ILxT��Ez~�U"O��/ϙA��2b�9�|��"O(��W��bh�ܑ�J�?N���z@"O~�@,�����2�h�ʕ"O�� �2z�^鲣&R(^<Ȕ�q"O"��'<:H���_s����"O��!�NZtm�J6M?e�ܐ�"O���� 64��e��'�(��"O��q��
�b6�X�l��h�"O� ��M�2),�s�)�$��1"Oe��j�-��aÖ:B���k�"O@���ھ)� �RE�*}����"O𼨆��3� �@�~y�))0"O0@�th��uuЉ�p"��s�x��"O���gG�u\�]2c�o �(�"O���Al�)-9 h���6�@q��"O����Э0���hl�0�tQ��"O�i���%{��誓)B^!�-�"O
)J��C�f=��RB�@�(R0+p"O�L�si��*~l��e�H�PV(��!"O4�j�'�;��L��'��Mqj�0�"O|�`���Z>n�Ǉݡ-f&i�5"O�YA�Bө*��d�$gFR^1 4"O�B�]�W@
[9��-�m!��H�'���/M&M�|*�j��A!�$�L�HՀ��щY�T�B�	�*/$!�$.V�qpa�	9�6��g��0)!��و=���U�F�/���ǉ1[�!�9d{����m��x	çE-Bm!�$�'\�μ����!���ƘU�!�D��kwޭ{��E>$|�)�$	�i�!�ԯJ�@�0��B{�=	R���?�!�>� �Bȍ�d�r�Ń}�!����
:<P�A�-?���P�\!�$U}L���(�D���H�!�$�dZ.�KdK^:��d�R@N)�!�
	Dx�p�a�3����"�H��!�N�kv�Za@ڔu׾�����.�!��H� DSqC�.�>qʶ�%%V!�Ď�Z�J� 瀅T�-��ӟC^!�K"�V��A�D0QTB�Vd݇S&!�$�=\���È�S�r#C�T�!�P�<h`��Tm�y��|!�07|0�1�к�����R:%�!�� J9��%��<Έ�C&�Ϯ l��b"O=򰩁?8�𢖨� ���Jp"O�Av��(2��І$#�ȠZ�"O���A\e,|#��Y
�ȐX%"O�`��Ը����t�G"�\��g"O�#5l�����J2�?b��*O�D1�ꃐ_9D�i��sQDA��')؈�����,�lG�kX�B�'�.��w�O���!W#y��╧�y��V"(BraH�}��$R�ɂ �y(^�z��5��B^v潹gK���y��[	_!�"�s鄥s�y�#y�n0��iF?_���o�y��ݴP�,�
Fl6JO�� ��@��y���#ݣC��݈�'X�y���W]�P�"�É/T�5Xvk:�y���-S��Q�}u��Ս��y��;i	�A@ -��t��)��̘�y�@[��:����g�e�tB�4�yrІ:k���F��V�[ǎ�yҨ�P��aC	@}x�(4NR��y�N������y���H����yr$ܛa7�yأ,��u����Ch��y���'�N�-сt\>%A$f��y2kS�Q� ۠c�[��!�s�V��yRZ;g�$(��Z樥��Ԯ�y�fO�|��j�!��X�beZ d]B�ɾ}�I���0��ջA+�4�B�Ir�v�(�ABbL���l	"dk�B�ɇZ�`�R�h���CƟR�8B�	�#���AIN8%������$I$pB�ɜ�\�8sH�r�y�DN�xB�t��q#�+�iR��X�\ZZB�ə<�8���i��aB��/;��C�	�,����@�$�J�����C�I4�~����.H���@�R(M0�C�ɨLRbEZb�N.�*���cd�B�I X��E��k��{sl��q�nB�?�L57(�|1OP6_�(C�	092�=Pʋ�^H�d�R!�)�B��#W�5��)Q5,4��_�N�B�I�T�~��D�d�B��s�Vp�"O�r��0^���au���Z��<3��'�����F�X�)Y��
r���6��";D��S�ϓ9�,`C#�EG��#�.D����F!L l-�r@�=v(�V� D����֩Sv
B�Ôy� A��=D��X �6v�+7�A&u+��� /D�d�B�S	�0��#C"���!�1D��r��[M7FA�B�B�p��"D�PsP+#����"�T�t���J4D�4Zơ�^��9���Ѥt�*�j�0D�l3s�@P��JW�O=1�D�S�<D� �ȉ�)�Fb!-�>�!@ �_h<�P�ݳ	�B�bfL�H,!�6��V�<QtCZ*MUD@��O%5m�@ǩi�<AH�}3@Yy�@�i�0,��O�e�<Y�kڧa�jxI�f�L���H�n�a�<��"�2L�\|�B��kQB�X��^�<!T�Ƀ|��y���ߖ~1�ē�@LW<��,��tc��f���fY��L�ȓ]-։k�&�Ir��9�+�.Qd�Ԅ��@����
��̱t�	�(�r���J��m�N�����/��̇�S�? ����& � +�&�R�}�e"O>�Ƌ
�Ey�0�Q���X:$��""O�P3��5zB���-MDc"O�I��ɛ�>�� ��F�v�ړ"O�l�VaõX�2!�n�tM�Q"O�ŧ�`&!b6*|r@l8�"O��k�4���!c�_*�A�r�)D���R���@��zf/��c؀M��!D�`pQQ3���sFY'� �8P�4D�)��Y?�X!8�U�����'D��J��L�����B%  ��$�(D��+�J�)B��R0�"Z���r�B"D�tHQ坞5�$i����M�|���?D�T`�טA()	�ND7*��: i9D�D����;�6�s���""fi�l9D�(���/V���O��{�0M�f9D�pb�$Ԙo���
U�_�(��.3D�$Qg����ȑ��}� ���2D��'�L�'N���P�˸��̘T)=D�H��U�IF@a�g�EDta��9D����K�-L�2kஏ9F}�-=D������>ߜ��7i�?������5D��! Q�0�x8HQ`O3�j 60D�t:2�ҺrL0�bO��~���*D����-4���jB�^c�)JA.)D�4�$@�:9B`(*��D�PH��M%D�̈c� 	z"��� 	���7D�@�iГc}��A���uqv,1D�hIc��s{�m_.Ia�Q#An.D�HZ�/P	0�,���	��u�2k+D�43�g�>)!x���(��DXb���g*D�܊х�4@��ӁF��Wl0u�*-D�0�ViL���1��m��eSGN=D�x�MA� �,4	$�T�<��m���;D��P��Q�LGf�4E�ѲI��.D�8�� ��9���D�;�5��m+D��æ�]�@4�S郧)1�t��E*D�X������JU$�( ���{��%D��G��Q��O���)�I#D�<�mf���@�L!p���6D�,��c�>=�2�Jad���4*0+'D�x���_��#�`Q0W>��"�c%D� �B�(q�!iR �g����B#D��c��,#���@���x0�e� D��A��S;i����Qɗ�(蜰�!�!D��a� �G�r')�9m�|̋��3D�PBS�93�%�d�1t���>D�0 ��Q���Q�DV�`;jp���)D��cw����]��K�^�X�z3�'D��#�'�H��`iҁ̢z�@�(e$D�D3�#�'��D*MżT��TrU�&D��{U�]�����:;����l D����&}�$9�ee��d�4-��,"D���A������!V98�0�f� D���l����U� /!ɮT�`g D�@0t����&�i0�E
rS2h<D��+�`�"J{�Y� ��L�r�vo7D�����&����^:LP��F�6D��#�
z]�9;�I�3�R�hՍ"D����9v�5R��՘[^6e�B?D�����ҔZ��q R$�a��N<D����ڀ[F��%�@U��x O;D��ٓ㍾e�M������q��9D���i�i9�i( ��*hvrE��,$D�� �,{�f�"@���SU�.m�N�"O>���.o�i��'��]����"O�,���34ɶg:��Q�"O�0��+��!��@�J����"O�l�ܜasE֮r��Ib""O����;U*�y����	�@��"O8����)���8I"*t�a"O~Q�v�%cK`�r]���"��e!�B'�* h�oJ�� Q�$�!�'��	�T�ؾ`�-C��	�!��, ��MV�n�|�)AR�\�!���p΄��»1�rᡇ�=f!�؁�^]�1��	������IP!�B�a?4��ٶEm�!�p�ͩEL!��!Ol5[6U�w�GNT!�d�b�ҨP����SӎHh��R.(>!��\��=��֥9� ����R(!�$��ay�ds��nC�d# S�"O�(��mθTD�T"�NyhT�W"O�و���	p L+kLTȧ"O����g	3�h�3�JjX� {�"Ohѱw��0Ezt�'-E�x!Y�"O4�(6�� �Ti6�їD�~��"Oƥ�a萢q>N�g�S8���"OdZ��߇E���פ�o���q0"O��c �^�}�.��҄U-a�� � "O���@��B�X�3���7}�*�"O�l�Ê�%�l���9�\�&"O�����I��-����"��{�"O��K �Y�KfX���JڃC���ӧ"O�C&<�\m���@�xa�h�g"O�Tac�C&E�F��#�J\O�b�"ON�(��� D�⼫%j�*9� ��3"O���ǈž~ b�����ot�Y�`"O�9��T�g �)��
�:��!��"O�ਰ�F�{��$,��{�"OH�s��ȩάeh�O6ۆ��w"ON�Ɇ,�1~F���+X ��"O�W���rнZ��2m^�д"OH���H�]�j����ap�h�"O�)5��!�vp˥鎆i��C"O�T ��4�P��%IW�[rY��"O��Y2)�J� ��e&(gH<��"O(��$�=2 1X �J�mRi�r"O$�����A����W��P�:må"O­F��<X�����	���Ó"O�l�v��!(�"���?8��PC"O�d:�.îa�Ѝ��kӜ6݆!P�"O�� V,���6ez�x��"O� �$��k�M��9n�8�xv"OD#է�-;5|�SŬU�/$X�"O(��dC>S,��x��2X� G"On-ANZ�5�� 2�d<$F\ �"O��(��";��x���ɔ,�D$��"O�`�
n�vP�g$^�Z�����"Ob�j�ǖ4Jq�\��$��D�"O�9�a�4Ӿ!äf;�P�"O
I8�A$���FH�,)�u"O�A��~��y4K���X͹!"OTɨ�⛚v%n@b(�\���F"O�	JQ"o3���fF�"Z�SG"O���I��r;L�����OGv�V"OJY+p��i|j�1 ��&c�����"O~���џiy�[�'3C�!"O� (-���B0L(4L0f�L?
��q �"O�5���ǺT�Z�ZEf�9�*P�"OHA�D\�L�<�i�D��i�~ S�"O���7Z�pD&��ꓳx�)�2"O!R�c�)b��0�r��)�Nlj�"O��q.Ѡ?�~١&-
�>q�9@"O����,Z$�R$�j�<^Z�S�"OPd�m[E�@���ƽuQ�SU"O�e`̛����ⒿI���"O� 2&o�&1k>���q@n˶"O0a��	�6����bO�� U"OHh����g����B�~��1"O��� "�h�4�MͼKa+�J�<�s���Je�u:��תN�&��
�C�<qSED$��� Q R#q�9��TB�<���Q4z����#�G�|2��lV(�y�ʱb�����;FA�P D%�yR��yl�ѐ�m˺?���bP�<�yҦZ0z�
ņ�4jLlP!�Ń�y򣙨}��蒃��*����W��#�y�ϒl)bE��a�.��`H��T��yA�BP9�k��-=��:����y�1T�FYR�K1s55�pP��y�E��{#�yL 9SWj��*���yB#[�E ����b�6,ed��ybឋ*Fl��O��Lmp͠E.�3�y2�L�SDe�������񅢞 �y�����V��gc��Bl�� d�Tx�'cT�ɂ�W�kI�i�å �bW����'�N�Kc$N�5̒���̴[hJ���'?��#�#�  _��V;}jJ��'5 �kǫ^s>��AŧA��+
�'=XU)R�HH  ��k@�
r�
�'(F���@� �Q۠��2ztti2
�'�B(�,�>9D�z��P5j� �	�'����)�f	A���P�,���'3��HԮ�}_@�+�#N��݁�'E��z� ߇Bdh�� YW�%��'(��WI��1�\z�$��UQ�'�N��%��Tz�[(E���A,�y2�*G�ad���^����a��y2'�<�2�{P#��!� �ϝ��y"fW��E���ǫP�hp[$�ynD9ndL8���[����EF���y2����Q�(܃YE��S���yr�U .�(-�N�SQz�!$���y2�2)3������7��Hk#�H��yr����KD���U��բ
��y�ȏ�*c~isi	,}��fB��y�S$-5
�*&�HK�d���$�y�H�(`��(z�U�I�HM��e���y�@SI�u 6/)�%S���y��t������!�UiB����y�+@<*�,)wJ��
����l���y2kX�<\�cC
-�Ԩ�'!Т�y���
�r$�E��x��r0
�yR��)�pѹ�n�:�+�Μ��yr�>��i��OlFe�gC���y��Ҡ3$�42���s�Pp�
��y��$o�v�bRÛkN��_�}VC�>_
�RD��� M�5��0�$C�I  [H�!0��\�J�N� wM�B��`���r���+(�8��Ca 1ڔB�	85
J��L�;Jm)p�@�sBC�)� ��ɰ���r/����#�<����u"O�u��F�\E����bE-�4�3"O���*V:w���Рb(���"Ob�* ,9���À�+x��B"O�5�ݐ[F��`�N�g�8LS!"O8ث/���H�e��_�>��"O ���Iףx8�9���.�T�K"OF(���P�-�l��a��BԚ�"O�C���r4$��#��M�PkD"O"�2��A=��1��_�<�\���"O��c��S�B��7ĉa�^}�f"O�(��/J"TW�x�J�I��r�"Oz��!����9x����h��إ"OV���.��m�P@�te�	���6"O����Ӓ+�P`i��̖U��=:�"O������g�H�@�jlVL�F"O& ��[9]�
�e��9J�B��"O�	��=0X�I��A�T��eqp"O�� -S�{��J���C�<�J�"OB�S�d��8lrES�.V È�{T"O�cۍC�h�P�E��RQ�"O���E�J�X�@l��-���"O�@��-�73m�[cM*>���"O�4KCl����m�DL�Q�v2"Orh�7�W�T����`�M�zf�0��"O�h�$�.d����[�>:��I"O�`��ڻA[2�x���d9�#q"O�-�EEK�8Dʤ�ׂ?��Q5"Oe`rM�c�(Xӣ�٧yT���"O��NݪUƤ%���̠<�(6"OY��ڰ8���P;5���"O|��w	4vuC�C�U�}C�"O~���m��ykP �_��q"O��i����"6!��L��]V���R"O�i��%T�u��E:�K36!v"On��tL��$���E*���"OL��T�_9v�xb��7֩�""ORh:3n�:0�����D	6�.�ӥ"O�pQw-���a
�'���"Oĉ�e��.;�܍���ƀ�!�"OL�â.Ph�Dpn�>.Q�e�P"OP㕏�%R�$�RE(?�`��"O8��)G:]�<�q�,%<M��"ODi��Y6P���i��	h�h�"O����!�0f�P���[�3�@�`'"O���3�J�u7�����m���J�"O�]���2S��`�s��g�f���"O�aAG/.i��l�s���}l]Pd"O&H��E�[B(A!P�P���5�A"O����\�3�����(ωN��'"O�1q&a838\�*�JM�0u!�"O*��q#S� ^&��C��0��)�"O^�`�iz������� �P�{�"OL�p7M��b�~����Ĭtꚙ�"O�}�%S
=9�y���Ǟ\�S"OԴ�7B�O`�,؄�ۚ-���D"O���@b��V��yR��lF���"O H�Q$�3W����,�j"Od ��h�B���`��/�^�i�"O��6�6bfhXt.S�E�*��"OdIbH�9qJ4�Ƭ�$~�} �"O�������(��k�QΥR�"O����j�B
��x�[B��E}!�dZX`P���?:���sea�]!�� �-�3��C�1��>d*��q"Ol��b�̾:-Z�gŵ3���h%"O������>%�,�V$��!�$ �p"OX-(B-��E0q���Dh����yR�� �VT	�L��_e"|(3�=�y2�W�--��XwK�*cn�q����y��J��jT�0Î�*�xa�cȸ�yRӷbN��� E��U���	"��y����.01'�M�<p����y�L�:N�b�"I53q˳���y��ۑ7��yu*˂&���hR�߹�y�B��6|b�8GIҭg��!���$�y"ɑ�@�L��`�?��l��O	��yRN�{9�e
Hv :VK��y�l�����ᎏ_Jlk�kU��y����hE,��A ��^'��&N��y�m\�Bj� �D�"��{����y�D�:��<�Q��6"А ��[��yʊ>Zp�q��ذ�jD�2�y��Ý5�p�;���^�Hq���y"G�#`rV�p�^�1�BJP%�y��ێP��RWH�}{l���ȁ+�yR�XP�qb�R��"��%�J �y��bt@���*q��hش�J��y� U;l8�q��Үc����E�6�y���B�M��-�`n�S%���y��Y�l�r5X�QW�\!'��y��."�:�(��ȘG!z���ʕ��yb%6=�`����	����pM�0�y��[  �L�;��,wf`� �y�@��`o�)���3(<������3�y���
Q,e�Э/&��J����ybFմV)6\	���2��݄�y�	�,�]jġ/D�Q'C��y� .��%�T���%z���E� �y"fOyȤP+%�ڟ!�6��&JƇ�yb@E%)����G�3�Ɉv+��yrAF<.�j,:bC��R_�H2�`��y��D�E0�h�-Imʔ/ٲ�y�O�h2�2�O��1�l��è�y£�$ͪͳ�hG9"�<
��@��y����K;,�q�
�P'�YÁE�y��0*��%�Bw:q��l���y"&��<Z,���N$c�P8:1�.�y��lb��:��L�_I��@ E���y�O7�3�!�l[8���C"�y"��iT؉��)eeF���`Ӷ�y҂B����޾iG 9����y2aC�/n\:AhLKP<�	�y��$F�R��ą�>K�K�j���yb�8<.zE�f셏4��Y���T��y�@�xz�
��+�
5���y����! @"˓ ��Ab�l���y�d-3���A�H��Ω�v��y	��v�MH���7Ӫ��5)B�yR�H�Vf< )��?|��E@e�͊�ybF�W�Zp���; �F��y�*�>�:�����xN���mǽ�y-,d±� ۔x�Jq���F��y�+�"1z���f&(#bm����y�G�
�R�D��%��#��)�y��:5BH6��$�l���#L�yɄ�s:8qa�O��I{5ET�y�*�
l��!g�~S�@��9�y
� ꔪ4�W�B��,qLX d6���"O��u��"�2�&H�>>���C�"OH�qR�mm��ǟ9�88�"OPH��O�=r��23�W�+��`ht"O�u��g$�����Q�0�G"O,�
 ��� ;����a�a�z���"O��w��S$��Vi�1 �"O�(
s��&�v9x�,L�T��"OBD�d������K�� Pć�L���;O�0e�2H�����̄ȓM��I"f]%R����˹S`B�ȓe"�e{�-6B����!%Gґ�ȓ(����y�*�s� ?�JM�ȓ [�E�g��$ǀp0�$���G�D} !g�"�+�I�!+LH�ȓO_dX!%o��4~ p��j7Ͼ��ȓ^��pǖ�z�^�[��]N3
-�ȓp�e���Y�x-S�'��	��1��ja��[m�9a�ːT�q��d��mj��n A2M�i�>u��u�����׸~��Pt�I		 f`�ȓ<s,`(��h���2F��,Oȓk�t�����J��B�)��,�ȓ.5n��t,�mܬyR��1z����P���I����SD��J�$;̍��
��� 7a 	wP��D�:�4m�ȓ&�<�3c��R ����rx^u��$��ht�ρ`���+rD�\��,��z�tc��bI�ɓU�54��ȓnx�x�T�%�ԢR͗)A����9~ɰ3M
;)�`dT&X�䡆�L��[���9z���5� *��\�ȓ)�:1c#���[�4y f�K�1� ȅȓ�"��0ș�@�� S�š(��ȓ?�x� WIօ's��f^�o�d��������N(I;T(05����ȓX��| P��$�`$�&�]�h�ā��F�fh����!o��u��#)T*���}d�s�^�8�\�[瀈5i�y�������Xu�i{��E�WXRЄ�5R��̀nn
�UDQ�M!�5��?��(RӷX"�P�hW��́�ȓ��dɦO��B��\��@�hz�1��G�|%�V Y�<|	bf�0�2}��p��1"R\�+k��y���
r����oSj��"�c}
��7�5k>r ��O�@��(H�E.L�����0p� �ȓ/�r�p��=�R�@R,lS����sT�8�'A�W(c�O�(�>A��J<���'7 X��
@2�9�ȓ9����ު<n�YA@�}t��ȓa�m�S/G�+y��h��хN7"I�ȓe�^�"��@�vl�"`��xd�e�ȓKp�%z���"9�L�h�@�	� �ȓvy6��U�E&R|���n��kv��ȓ0L&�
�j��VxR����u��X���@�c�>�Hd�Al9G��ȓ�"�X�E�V`9���~���P�D���*@��hp�R0Mh���z�.�`aɆU�&�0F�+=�ȓG覈"#�
 +�]��G�"��a�ȓ(X.p��皍#+n9(P#S�Q�Ta�ȓ`�t�#"�.�X���\$�ȓ'X�(�dZ,#�ָ�P&��h��S�? :�3�m�30�q!���Ug��"�"Oʭ34D��RT	��EI	\���i�"O�Գ`��� ,����5N�ڜ�"O����DJ�Jk>	Xc@�`�!6"OFX�d;w����G�7x� ���"O�E8�̄7��S���'=�^!HE"O<`�c9!�Xe�$.`�6X�"O虹�m���BF�آ,���d"O�|�P�A;BP�:���h�n5��"O.�*��߀+(��3���U�H q"O�ܓlE�&�pcr�]�J�8�(�"O�@
��4�NyɓO��=-���p"O��z�5C�p�y&�
�����a"O|)�F��h&y�����*�����"O&��#%��E� �픖� 
%"O������75����f����M!�O%UX>L����84�0��@��-�!���X��"C�2� XYga�K�!�䒀g-��NG�T֨@�
��X!�^�T�u�D/��o6p�$ �hH!�D.H��P��&m~�C����5!��л576�P�UU�̙�ҍ��tG!�D��)@����]�.�yP4&Ƅ>!�$� ��͋�k��F��Ő�!��	
�uQ���y�:xУ.�!�X]��\��H�';N"����?b!���U��#GN0E�$9ū͂Y!�$�>8��(�/�;q+:L�Ɖ݇*�!����(^>���k0���N�r�!�Ǉ+
��l�l�rz���m!�d��͐|�����@���-Xt!��â"��D(�I�5?�}���Ѥt�!�䐓9��u�5*	��鷧��J�!��A��U10\�'��Q�D��Z�!򄇾5n�ö���	4��}p!�d0	Q��U�=�����Gi!�԰B�~�2�
)sqБ��bN�W!�dN x��x�n�
[px5!0IG!�R�'�蠠�$�2qpq���A&�!����h   �E�|��R">!�O	��ivVr*&h��ʙ1!��Bo(A{Ǩ��:�z�I�H�!�$�q�"�W`j�d�D*�-�!��A4l��ީ/�Z�b���!��5$�"��*
�l�Ӓi��r�!�D�!.��5����x�pF�Ya�!�DD�{�� '��s��C���!��I�L�]s6k��2T�5����!��#\�vqC�Ǘ55VD�w�	�v�!�����k�a�:.ƍ���-z�!�>Lsd�a�ޛ\{�0�p�ĕY�!��[��@��#�;|޽��"��&�!�D��������;m@�i���a1!���Z�<�Y+�:Xh�����ī#!��L�L�,�ΚL��S�+C!��O�+b=r��?4J8x ���R!��6r�,���^0#2l%��+YSg!�ˡ5�h���jQ�j�6��&� �Xb���<|8|zD(�7{�	0��
�y+M:&���0J�z5
y��:�y�ʖ)8��%��D߄x�N{qD�yR�Ⱥf�^h�U"S m�T�Jө�yRf8L!�lX��d�n�C$*U6�y�	�o-� ;E���a����V���y
� �y��AkFk�*ŀ�b�"O h��I�	�T��Q��,4�"OF�;a�ޖD�ԥ�5L��V��A�"O,����g4h�p�O�[��rf"O�P_1AtU���C�6���o�o�<A ���uj��W�?4
ܹ�l@i�<I�A�49X��������}yÍ
A�<ᢢ�f��śf�߄e���b�(G~�<�� �c^����J���"�q3�Dx�<A�U%JzTB&�Nz�l�����N�<�g�Qo��1 ' ����L�<q�j=f"}�#�W}8* � " D�<Y�\�_�QG�qMȬ���e�<AUA�u���+��|xЪS&d�<Q��/_���Xv���doμ�W�Lt�<!�aۄ�Z%PT��(Ԓd�0��I�<�w(�g,A#CX#r���ҠC�<��L��|4�Yh����I��a鱭U�<�DN�>ID�
����"f�5YG�q�<1��4a#&P��쑅X�>EȆ��v�<!b�M�W%�m��
LAV���ׂ�u�<���X�TD��{�z@�$�e�<Q�
�]>�J�(N�a:��ՅNK�<����W�a���`<L���_�<��(^S�<�AD/G�Hi��e�^�<�!=ɲ-�A�(t��}�aD�\�<��*Y�挃cb�(:�l����[@�<!�[f'�[)��pnXِ��@�<	���WM@��!�E#Q9N�@��S�<Qe`�)P5�Ya�� 2���su�<qWI�Ұ�0P�Q�o7�����Z�<AG���2ږ<��e˕@o.�X*�\�<���E�$V
��ԉ̑~�,�BG@�<kҤ\��@u�J����g�D�<9���irZu�r�UB}����
�J�<�uE�t�1�u�-����QH�<���Rti��#�� [=^�r#��B�<��Q���UF�?K0����LC�<9e�"���[�e��l{֨^~�<�$�\�5�<�H���$3�����{�<I�d��3�zE��'8�`<C���w�<V�O7+%��s S�-0�Ԃ�Ɯt�<AP�ڰvt�1À 9,�2q��J�<���W� AzMhc��K.���#�<I�e>%ơ���[ BT�X��p�<I#&�.��J���@��̘!OWW�<�«��iҵ{C�A,R�] r&�P�<!1Q0:��sԢ�=�����`�<i ��ܭ��P�z4~av.�w�<4"��b�����M��)�&��t�<yd_�iF�Qo� P���rc��p�<IQ�0��ŒE���9��2�MVm�<��&y��1�� |��}�fi�<Y��=j�9C�	�/m��)Ԯh�<���h���A���^ѬQ�E�a�<�~a%���c�ĩztN�:SV>���x5\Tz�ă;z%�@��6$��Շȓ��uڔ�Ry�P���6CoF��ȓ$�2�)��c>����W�1���z�����z&�W<:|4�ȓ�"H� &�)_d85���68>��v(�X¨B3���r�ǰ#Z !�ȓF4>9x�-M$O -�3%E�VM���ȓf��<r�dM.O`>T(Yo����S�? l�Y3N^�l�Af�ې-O��I�"O��r�	�˦x��M݋N0���D"O,��n�xC��Qo�"0v~xZ�"O�y�����>t���TN�NQV�5"O�E:��D;+�L��F��N�84"O��j�b^"g�Ȅb�KW' ����u"O\5�dC�0z���A��(^���v"O�p1u�ϨXqx�Kd�H�N��;�"O�x���ZG_���B�ZU��@'"OX08â۰�c�і<�:T)�"O|	�G�b�����͛># ��S�"O��	���
`q��4]F��xp"On;.�"�%DHՎ�k�"O2�c�-���S���4��ٳU"O*�ʃN��1C2(��X��:��"Obq��*��?�a��jC�)E�%J�"O6���O�_�����	�!9�V%�"Ox�A"o�;�Ճ"J[#�J�j�"ODL��O7l
̭kg�ק7�"P F"O\�"#�E�0>Xp�̂ ����"O�q(���@��ȉ$�N�/S"�[a"OHlA��#hϺ �B@W",���"OX8"E*ߞ_�&�c'������@"O��kQ7P�Fa����U�	��"OJYA'a�5W�L(��	��Hr�"ON1aw�Qv�˳
��wϐ0[&"O0L��@�xO:9��B	05�|���"O>aR4"ʟU�����CF�Ԙ�`"O\PH�2zB|X��
!/�nU e"O ��B�F�鎍+6J����"ON�WK���y!Ó6r�0�$"O~A�GY��BdO��|�^9��"Or��ר�	�b����<D���0"O|`�1���[�ȵx쟜C��+�"Od)b��O��� �r�2��"O. `�M=����5D�0�"O*hJ�D�M����f��-�Ҹ[�"O�9ca��7\�|{3��a��8�T"OA�!�ҹJ4�A�!��$1t2 ��"O}����F�f��֡JjԠ��"O^�cq
�VZH�j#�8=6"���"O�	�.�	x�Ľ��'�"Y��$�E"O��D%�*@с�>{�0!&"Op�1�iB�.��i�$�:⨸c�"O�9����b�f�Cd$�c��|;0"Or4���+rd�у�)��*��	R&"ON		g'V���ZΓ�W��1p�"OJ��uKPij�9�$x�.p��"O|�jGIęv�:؂pC�	R����"OP${�Ȅ4|�p�!��sv.L�!�$A6awа�B���|�\�'hԔAl!�*#@mP����\p(a��F
}�!�dƏv��t[įD����U����!�ėn�R��eY*!��!���*^�!�D�63ҽ�נ� ��0	f��+�!�(h>:y��@�J��e¤���!�DE'�ؕ8M�GZ��D*ɗq�!򤍘|���{Qn�HH���j�*�!�d#pܴ� .ֽ~�a�&�J�M�!�D�l$� �v�����MD�!��~�Iz��_�b���*'�T�Py���)xD��V�t�x���4�y��%�1�N�?|�� ��Ů�yR`�g>�}1����l�YXDk��y
� T�C���:
��i($�����R�"O��P�!k�*h�$�v�"O.kl�1���&���_�
���"O��� X1O�%Qn7B�b �"O2�h��\���l[�N�W��X
"O�"复,f�Qy��C�`�^H�E"O�(xdhOI�dœ(V9c���c�"O��<K����^���Aa"O�ܠ'g�ovnp���;;�^��"On��uɁ�y 0�L?
5!"O�I��iK�i�(��m�a	���f"OJ����ŏoP6�GjQ�"�P�"OL���մ4���i����;�"O@A�%g}�qR��1׼i "OƄY"�Ñ{��Pӱ�@1;&<�p"O5�S���<T����#$�hP*O��� .,8$<J %��8���'n-���?|�Eiԋ�3>vb���'C��jA��g&� -�m��0�'��(2nJNt��X7Ҳ}��'��5QV��;+�4A����	��'\xe�e�ËNrάP`E�逑��'�6��w@P�V����g_3"�s�'�Pd�c:D,��!ӊM߈�a�'@ eWʇ�'޼���>G�D�S�'[�ɂD=t:��&ʾ=IP�x�'3`h��8_��e@��l��'�\��R0Vz�4�5�>r���	�'��1�B
	�z��T�i+��a	�'��ܒ�'��?KxX���T�
* �q�'�4͐��]�|���хƀA�`�'[��J�+ٱc�ȱ���F�5�:�i�'����i�� p:��LO�.��B�'�`��d9;��`�����!
�'���"�CCd�M`�,��y�^�Z�'�$��lT�d�*�J�;fp����'���׮ު�<
WQW��0"�'4U)����`�/�
x���'p�ia����*�`��4~"��;�'��:ԌW�X��6�%w��j�'7X�Df�1g�TX�+�uN��(�'��l3B@�l-0�AE�gʵ��''��BCi��'��i�L0��'��l����
QP���oXR�|���'�٫W����|@!l�?���'���!��P��x�"!OW�	�	�'��]���ŕoՊ�3׬�
0mQ	�'���LJq���� 2i[X8��'�Y�_L���`�]��'�����ɤw��Y�m˔T��a
�'�u�eH=}@�@f��SY�9��'�J` F�ӊ�`�
�9�f��B?D�D2�i��<i@a�qnɋp�����<D�` Gđs��9�Vab���>D�ā5W;9���H�WyF|{�!D�,��T8Sְ �4 r� D�Pk /_h��HT��.Iq`۷#3D�4��擥?8�T�A��Bx��$1D�t"�g�10aZ�#r I�@�Ε��-D����IӥY6�|Q��ڦ%Mt|{G�+D��鶄L��6�S0'���7�T�<��A�G'thP���	����g��{�<�4�4 *�6�S�]=��	�u�<A��P(SF� ��~u6����Gp�<� � ���N+�ii'.% :0"Ovqb2Kߟjk�-���,*T�"O�; i��g�8b���B"ORl�A�_�Rmx�"�
� _���*�"OX�hˌ]Il��fIPZ��@�"O~y�G�	c�lBNϣ8�~��"O���͒�z�Z,�,�&*l�I84"O8=8�۲L#��������*�1�"Ox��ٌ$%���B0㐍"OKI�v['�	
�ƌ�jH��y��Ť4؀����z"�Th�(�y��P�p$�:Rb�n���c�F
�y"G������V	c %2��X��y2(�)%�5� ���R&��y은L�֔� ��*i���ϝ�y���#W�{Ħ�#hp!�;�y�mԈ�q�%�%*��8�s�	�yR�4$��dD�[�(X�イ���y�Ms�ƝCg���V/ɣ���+�y��C?@�����O�K� E��,�,�y�Mޚ	U(���D�"Fe 	�B���y�K\�6?Q���+���"��yB�D R����bf�#���1GY��y�Ӂ`��q��H�H	h�cS�y"��WɮE#RBM)}�0@f���yb�S��~5�̘\T�@e�Q��yҋ�����N& ZL���L,�y��M$r�Y�R,�*t���j� �y"�S�8��Q�7c
pym��͛�y�$�)cF�(�r)��j�&0���X/�y
�7���B�Ͷ��P�����yBJ%U�9�G�E��r�
��y��&_qD"�	H�}�`�`���yB�P� Ҵk%�i
U"�G�y�X~�4c��'iպ�p���yB�NM =2�ᒴPP`=`�G��y��_�	��@b�4{�H�6K���yr�p	�1r��Ou)T	6H�4�y���+?`���E\�c;��A����y�iC8�©L�X�.�cѠ�y���$&)@u��&Xu0!5/��y��A8!�r�e�G�T�|��+�-�yr'O:v�Tpp� T�XzĂG�y
ЎR�D`�ǂ��hP�DhEL�<	w$�:c�����Ƚm�l"��w�<��H9���G�<hy�4J�{�<��m
^n�"�7M.���t�<���*:@l��_�sr�p@d�s�<ɂ��d�Ҁj�D�?�:���#]z�<y��$Sx^���b(c�D`�Ms�<���?�y"�N���r�iCE�<9b蘼	VP�E*G�#d=����B�<A"�>djIK D��I|�� U�<�T� +n*�J��	�4��#PT�<����!'Ψ�d�Ǐ9Y��#2 XN�<!�0Ja6���"Uu^����G�<��/7!኱��e�7L!vόD�<y0J��\h,�� �K:\���p�+Mi�<�$ˋ�..�1�f�� e�`��T �c�<��gZt��H1�^�EX�z��LD�<q���"���yp&�<jn�dMy�<�R�Z��\4i���7dyҁ^�<��B%<L��a��z)�
T�<�M�g��0F,U���V��W�<� |���^�i�z E!�@3�"O*	 �ˍF ��ȏ� �Eh�"Of}z���a���JTh\'(Q�"O�Ā1A�W�$��'7�,	�7"O&4�r�µa�dpFk�5:�
��"O2q%�ЎC�i��B�4�.h�"O�<�*LO�"�3�h~�`M��"OƝ9g�4M���IU��V���ڲ"O�����< �Lʒ�׈!��V"Oz����E<XTp܂�A��{hQA�"ON=!aN�0)4�%Rǀ�@_>��"Oz�q�K�_�
���N[N@E)U"O�Xa�a�*7��`��nM"6:��9f"O0�Y�C�!|.��D�R5�4��"O����"M%8���Q�j�`�s5"OЈ"&�Ũ:&ta��f�=/rK��yr���>��5PČٛ~02|{����y�D�r4�0��E܋o��	Y����y"H�/sX@hKM�_ꔜ���	�yr�B�Prb�bOM�.MZ��RJ���y�)��H����B�Wo�2���H���y�ƅ���ZG�g��"�͂��y�bV�oLJ���Q3af�1�G+S�y��ǏSU4��g��� E��y"fW@"�$�"�Ҟ]���6�I&�y�0�)���*ZX
$��e���y��_dzCh>e�X�fҧ�y��3oqJ�!1�]?+��]d��y��ݧU2Aذ�E7"j@ˁ����y�(�<\��x�"���ƱJ6���y�@�!;��M�S�b� ��V�y��Y5�ܩa N;H�|I��M�y2����`飍E�{@��@��yҊ��������wRDi	1/�y��9!�lL!7@Ƃv�
Yۡ`\��y���@r����çf@�U*-�y���R�*�гŁ9f��*�����y/(��J�*^�`O"���(�y��_ $欉Ģ�3o8�\P��ƪ�y������Ӝa3��F �y�H�>"����\�4������y�N�Wa"�W���S�*%8ND�y�49�f�׷P(څ��y�兤x, aN*M����/E��yr�U<]�8�e�܊�ƴ�d�
�yB�2j�q��ɟv���Ƴ�yr�/=��1s�0ѰJ���y�/B+K�ΐ1ώ#,�M�I��y�.M 7zt �G��; Dp�U��y'�$$� �㒈�<�Qe��yҩ�6:�� �X� F�{1,L��yBÌ߸P�$'ͳY��� C�5�y"l�C+�����BPn�
�y�m x�P��6�*����B��y��$�!�����l�'�:�yB(�'-Ԩ�29����EÒ�o^�}�ȓ ���DH9���[��x�^I��@�8Q�U��`d�#��Q�8��ȓ-�v-rᬏ�w���* ^�F��Є�x��H&��JGV	+hQ�ȓ"!���q�N�s���0MG0,�r��ȓgl���u�R?"�r��V�ȃ\��ȓx,Dq��՛E�rl�$.D�M�؄�ȓ@`�����;_|R)���`��S�? 2L�r�9X�z9�4nοO��:�"OT��ZO�ԎM�o^���E"O��"���S�d��䌈9xU��Q�"Of`{)�6����L؞+b�!�"O6��ٗB,"U���\Љ!"Ohȱ$��
�~A�wP�L��"O�0� K��\_rܸrÚ$lK���"O��;�*N*�Xp�r���NE��"O�)9s��ksli`4�,1����4"O�Mࠪ�6E�.��AK/�(��"O����A� ��34L(��|@2"O��D�	6e\�e�X@`"Oz�h	c��,
'�ǣ3fͰ�"O����܎N�f!`��ʿg��\�""O�0M�$`,��4d���vy&"O��a4��'"�$��	�+gm�DS$"O�i��Eհ
AJ8��n�3>X �
�"OR8�M.M���ԍ��U�@��"O��cva��CI&q�Њ�)D ���"O&�k�A�c� �A�ˎ��aa"O���]2EjR@X��
3=���"O$�U��&�0܉@Oߩ{���c�"O�� �ѥ1�t9å3m���"OXl�vG�f <��d��5xP����"O\���ݹC�
�8B�O(,HB�"O�y��~#�u��g�2:zAJ�"Ol�SH������AR� 8Tu(�"O��U�rR$�4C�'�A�"OűDW<V��sU@�%��"v"O(a�e��� ��,q�jpK�"O@@���5ۚM�P@Q�"O����-O,(��K�!�H5"OH�ea�cU8Ey#+�q�,!"O`aٳh��&m4q�2���7.q�"O����?��	p��(���P�"O���@��$J@�隗�R�ߦ �"O yIR��
ȸ4��!"����"O`�bT� ��ܣ3�#U���a&"O�( �/">2��ցW;l%�"O,�괃��U��� �-"^@$��"O���;�t��o��C�"D�D"O8$�	�}����ؔt�Ac�"OU1���F��|@`-�����R�"O��Y5G�
+.0�æ���4��"O�\R��-`�
��ȅ70�<��"Od����J�Q�"�K���;5����"Oby��ϩ+��8AAڀ2%�4hS"O��S��X�py,��El|��q"O^���.��D,��0ra_���k�"O4�9+G�d��/�=m�j\��"O���h��<�TLS��N?�Ha��"O�HI� ��D��H��Ƭ�b@�""O�T��}QB�N��Z����T"O�� �۠	������nxl�"O�%��
�
���h��%\`cG"O�q��	1i��Ȇ�xH¨�!"O��&#A0n�!D�K�[ fI""O��`��rZY۷,Åo�@@"O���^3P� 1CRn^�/�6���"O����t���/I��8,�B"O���r.V"s� � ��[��6T�"O�Q�G'Y`�J!-�|�D���"O>p��W r8�p1��C�{��ԙ�"O� ��O-b����%%�?�6-�C"O� (0����'= �[�3mr~�
�"O� s�m�~}���M#�ɫF"O4qR�O�;d�y U��E"O������5ȥ�� `��QU"O�x����YކP�#�<W��R"OP�[�"�����Д�]	$؎x��"OP��0��2@����ց?��,��"O$����\����"F-=N<AS�"O̥A��I�zFX`���gH�=R"OTؚ�]��h� �م0�l��U"OrL��oR@��� �_%i�� U"O��"�¿T7L�&J�	V�A"O�C�&,E��s���>D�xG"OX�)T��6@��<�X5��)V"Ov(�t��=o��}H�� :a,���"O�d00#
�Q`� 倈�>T���"O�$Q�i�e�0)2t�ݔ\bT���"OxH�/��6��<SUM�1pj�8"O\$"W���;�@*A���p6��"O� ��A?H�l�F�K#/����"O�H�--[ �ᶣ�!6�qz"OP���AQ�n8���u`�&?2��c"O� ����G�@㉝ z����"O�$�D���;B�u�S��]=(�'"O.e6���Gs�<p����)LP!�ƻ<S��A�hV�+�ڥ�s�R@N!�d��s�vh�W�ƌ+��C� ]�7b!�d�t8�Q��
�y&�=32 ���!��\N�\3��Q )������̇j�!�dڴ H᳓i�&�\�x$�V(�!����`H�#L��ts���k!��T-$1�$��A��!�\�~�!�0�&�S�lO�1�Z����Z�~�!��ͣ|m]�"��Z��.{U!�LC�hh����$HP���-lF!�$R4a��M"&��gp:��Յ��rB!�?�dh�B��U_�����ՆA[!�D
2'e�{�K��M^�|Quk�!�Dĺ, �!��G�wCܙjaي.�!�$"j�!!�@��?��a��)�!�H�
�b`�FA�k~v�b3&J"9�!�5?�<y��U�M�W+�{�!�3V�D9�u�9.ob�� �ر+�!���)/P���խ� Fi^U���Ϗ7�!�,(J��5��d�D��@'<�!�dA�&T�P�fT�S�1X`aͶ�!�ϥ��SZZ��C��/$ P��"O�"J�1 �d�g�m3,p�s"O�+`�A	chq2���)��Kt"O�|��M�$8E���ș	�P��"O0k�g��%�R��D���T*�"O��35nH�m�89Ӌ�>����C"O$�iS�BҐ9P���7��`�6"O�$i'ǖ�E���r�#C��>�(�"OޡITG��ad(!�v"L�mI~�
�"O���d�E�;>�Js�ԠD9���'�����2�{ЈO���l��'Ӵ8k&�.=��IsgW�St��
�'-�����_5D��2�C>M���
�'�`�q.:f(�����>�x�'i��#&-��X$�S	�Ki�
�'�tɋ#憱�P�r��A�@B�	�'�
�sfA��GF8��� �?:�
�'FZt���X�ll��]�;��Ÿ
��� ����J�L>�pt���8l.4��"O H��F�}�40�Jʰd} �{"O ��&�&��%�3�)Y�H݋�"O:��C*�*x�BMM���s!"OL��ި,%k��Y�v�9"O>l��9Z��Q� ;H�"ODuc�"�����[�)$~�1�"O,���=��,�cU�c��Yq"O�)KEƝ�h��{�AU|>�[@"Ox�t�[ L����^�NS"O���	R&VJ�"�,5u���'"O���)r�H��m4g�Ea�"O���"��p:��sw-�W�P�"O���2i	��KClX)(.�2$"O*�!UIח$���is)�mr�As"O֤�5�ޓ�
���(��G\" ��"O����lt��� sI���"Ol�����,��Ⰾ�1e����"O y���?�F�02�85Xd(a`"O�!��L�o�FM)����K/*�t"Oj��m�=.����4>��"O~��g��n1������ј4p@"O"M�1�D	)��=Pr�D�M�.��"O$��c%�hU$P9J t�*��"O�!8��ҫP�:ՁR^�J���'"O�M�3��'e��f:n}L���"O���kBFn��Q�l��t"O�L��M��#x���dX�c$���W�PE{��U^v��a5<�j��{!���=،��Gڏh��-��j�!��s6z1�s�@U�t��%�K!�!�D�c��4��w�v�󵋉 0�!��	F�FȢQ�ɷ6]�Lr�j?`y�O\㟈�|"WǇ{Gh��CQfaD�bQ,P[�<��]/UWV���FG�F�pԓ�y���+=;f� Ƌ������"��y��S�b��8�K�
 �D˃EV�y2g��pd�b,�.|�n��2j���y��	a���b#�ՂP���b�	��y�0���2@P��L�À'I��Pyk��fن�E�U<Ț�D�i�<��E)7x�y���̸X*���6&�e�<���7c�X]�D*"��\�c��e�<��e8b��Ep���qI�����De�<Y�o�=��%��@�"/,��+G�X��x̓)��4Td.hp(����5J�tɄ�h��8�gZ<J%P��7=��ȓ/hP�h�ጭa|F���!K5r�&��0z݈e�E� �����D0	�6Ѕ�_���U��O�b��5(Z5i�DІȓp���%�;dUZ�1��rb���oZd����c�,,���X�����	i�'�Ey0�po�]��֝��D��yB�'9\�aBwn@�`F��9��r�'cȌ�P�M�L���%�B��p�'H�u٣��O��L��J[4��)
�'�L=�s�Ӕ.��᫐N�;0px�+	�',Q9���B�� ��jԳ*r<���'&���&W�H�0�:�'֬!�j������H��-��k��q�`�(-E�
`�|�/Lq؞�C���)�@\P��I�I94 ��(�	Q��ħHl�aȤ��3Csb\�i�G�,�ȓb�b���oɩ>��@
�m��OO�0�BK��'60G��O��^��̚S�48�)�"O� ���ҦL!H���$����3n�b����R �& �ZȻ�O�>,��]0�k�&�y"G�<EQ%r�|��D�.�yr2?Ȥ�Of�4`�yc�%���?Ze�o�y"��i�tc2��!�1���yb�Y�m�݂�.���؂�D��y�_c
�0��m�3.p3�-	�y�OY�]4Ĉ���wlP�4�6�y�a��pY��ǎ�_x��a�
���y��N?^5B�d+9�����؞�y"� 8�p� 7�,|��	��#�8�y�n��_jeɷ(B�ՠ��r����yrN_�KI��0�Ů1�PH�H�y2�� ��)�Jӡa<e�Ci[-�y��ˎB�2�HC��T(C��Z��H��M��a��g\�t�p�ɀ[�<��+L���֥�4
�h��!��3t���0P��p&ʀG�f�Z�g����.������r�}��Pt���|�
�B"�ԉ	�<�A��M�ԩ��O�ȌP��Vk�)��Ж~R��ȓG�X�[&��P%d@a��� ��8�ȓ����)�qWB19���
Ϯ��ȓ'�
Pz�>r�R�Ȃɞ�/@�a�ȓwȾ�{�+R�d�N�!�W�W:&=�ʓr��-��V2tbF��0�+mBC��?{�s�jD=3&�ɵ!	�C��B��Yhz\ZUj�:jhƵ��R\&B�	4
z kTk��*ݠm���D� B�JU����lӴB�bI�ah�"&B�I�XK�i�T*F�9�L;��ܟn
B�'�n���GC?h����\�X��B�	�.�8Z�J�M+\�T���f��B�I�pW��c"�:p)I�`U\�B�������;��KF��G�:B�	�@d�Ԙ��Z(G�����*D����ki���DKʜS0����=�!�
�,X�0�<M&&��-P|�!�d^#>_,a�ĕ�G#*3�MR�]�!��%������87`���0?!�M%lĔ,ᢟ�az$1�� �7F
!�y?������>�Z�yeNO�d!�$ߗd��$�>uf�*��,c�!��!�v�����,N;0)'�;�!�$�Cٸ1��5u��0d�	�"!�d��f��Ŭ�#
P��{�/��8q!�$��}n5P��/9�BXjtϥi!�D�����+͕$؈tq4�Սl!�W`�� ��[}��0�ͳ)�!���#{���cC�S�t��Y��BJ?�!�V�}ٶ0 �f��*�4ə� �e�!��ϩ{�� �A�@e�(D�ק�!��]r�򁌢6�&X����Y�!�$�<�����Z%w���X5%N�t�!���K��9�B<nirT£�#�!�F�*U@�C��;R����ރ�!�dE�Cl�l2�� �� b_�g�!�D��;�ؐx����b�{����!��'���`*R�L���K�F
��!򤔔CŶ�K�̟�.��&&T�}j!�$_�qTH\ L�
�؄rs#V7"!�ߧ:�&�G
�9v|�r%�� c!�$�YD6Y��Z.&]@C2'*q!�� ȉ1��ЀNE1�e�"S���"2"O�%���� yJ٫S��8Y�.ݹ�"O>�R� եƄ�PR�_<�!��"O
��#V�#K� Ywo��<���e"O �9PO_?>���%/݁*���;�"O���,���@Rc�_<�@Q( "OTx�F��	;^�`����,��L�"O`����)S�z ;�D�K�h8sd"O����!3t\� ��ͳ{�6�0"Ov8���5#���F�U�#��"O�QPJJ8*��l�&���0"O*���4v|����] ��	� "O
ä"��T��� iT�<�tiH"OJI���H�h��p�p�.'��pW"O i"�\�5f� ��D"-�y�"O��D�C}�D+�U�1)4�Cr"OޱŊXsH\����(%���"OdA��ri&�1`��U{�}P"O�{�G�+{Ӝ���S�ubdab"O||ٖ��
k�f�`L��(L�� "O��0"#	6+-f�˱��5"�H=�v"O�d��V@�QL�'n�=��"ORD`� H+tVH��喙gk����"O0�0�ؙ~�Xa2T�6FE�P�d"Om0G�$ev��#O�h<� �"O��J�"HR��BY(Z!�Ѕ*Otm �64����ql�4Q�'�@t+�N�L�����ȡe�����']�6%�ZT�c���VeD��'=A9d�G�D�`[�Ă�Nk����'~�9���0%��q	��F��T�'��"Q�#[|�B�[76J)��'���s�+��nj��j�}u��Q�'%��v�N�fC�q���K>^>�}@
�'��ɳI�2�UI`@A�U��i3
�'��h��1e�\��Dl
��x��	�'�b�ri86$^l;���[�Xx	�'cz�(t�KZDT`�a[�LO���'�^E� @P�N��$c�ċ�L��L��'�tHj1��)]HV��FG̈́U;B���'�pQZ��B�.�I���G�j��'x��q�ٕ�fؓv���v��-9�'�%�Dc?�4����W!9;y�'I��+Rdݨ(���8��ʷ]O��[�'�\L
��V�D�
e�UCN�W��hq
�'��u�Z.,�x�E��T7�	�'ATHI��!��Pō'K}�0z�'�<�ѭ��VM��<b�k�'��HpQe�e�R���2ζ�R�'��"��H
f��廔e�*�D��'���ƌ�=LVH�XQM��0Z����T�b��; ��>r!�䚑zF��IRσ1t���� k!�D�&k�t]!��B���-9&�Ѝ�!�dM)*:���6{�`�1�C��U�!�¥��x��t�xG�
p\!�$�@٬q{V�<~��`�L�	@!���I%�y�@�C���q�d]
zJ!�^���Dh5��^����ף�PK!��s�M���k���W ޺l'!�$�7`>� �Ō2w;P�U�0!���B�@!�ō9?�>eІy�!�D��Y�z���J����� �!��߄q!@���Z�,X3��"8�!�d�"wA�q�b)�8HO����ձ�!�� ��[�f�\���sDؖX�} �"O�I��l@0���:q�F��T��"O���L��E��	�)՟��}؇"O�BeE^��T�Sw���Z���d"O��R��lu�pc/�	K3��"O��B���Iem�<Q����p"O�\��ҲJ��u{���� ���"O�X�P��/H��D�"�ܥK�:��"O��[q�Z���q��Pp"O"a�ċ�%-��z���V�\$ӷ"Oh��&$ب�&��.�@ǐ)��"O<�:A�QC��H� �e�,ɀS"O��ʀƄ'Y��aA�H^��x�"O]Z�Mތy�N�0�+L,�|�A"OB[�BE�dlҹ1��Mf�x@b""O�E��}�e�6dߴY�"O�w�²BMt	��ԌB�F�¡"O�Y���z�<����^�Iߦ�@�� ����W�C:<�A������_�EU&	v��R��P�R��y����2�TI�@�Ϙ�0��pċ��?!S�w����n��E�܀���(Ȥ�'��}��	�p����ɷ1<M*#��2q4��IPl��n��AP.�$� �MR��R��f�'��:0�~�0�ȋ}��S�{�>��9xg�� s��� ��=A_�O�]���J�#���W��w"�U#�'S@�X%�D�?rl�6C�15�p=�u�TW@��C�?h6�K3���j�'.:y���0N; xC��� 5d� �'��X��۰
� a5�Ҷg�S�O�E���P��U�$u��_:��@��ɋk�P�e�0h@ =a��Cw���K�`ӈPR�(��5��,@�֠lݬ�Bd%T<B�j��` �:	\���m�/FUF�+�[�txi�\�J�h�#�iS�
�R�$�Ԣw��'lR���K�+�f�S"���y@<a�FQ>)�CKI.	��@&S5���$�"D�@�oԴc �85)΃�2ED���h�Vis���W��H��ӵ@�rH�N~r�h��B�v�$��Ǉ�~�>�"AEϛcm&B�IY4���AL����Hנm���ueîn�BdPTd��`%��8]Q<��viF�'�Iz���,m�8�3�TA�6<
�^������V@��@L��D��yf�P5�<!�+�]W��:#� C-д�:)�mL~��w�$w��1D�\�n�ܥO��CP(83+Μ��,��P�D����+��~2��	(��II3 �F0�i�7AG�<�� �7�����Y�1�q�L�h&Q��X�8���C�� ��Ba�� �������+>1�Y�׼s���!?��ɥ�޵ ��DPx����$ÐV���B�&Ɔ�+u΂�ߌ�P�嚓x�,h3�LY8U�6H�0M	 V�%��i��"ϒ�K��҉'Ǻ�#_!R��f!PZ�q��\H�'�ʍ ��8AzZ�9Æ� TS�]�"M��dPܽ��)F)�J��ŅE;��SgF�X�r��p�\_P��- ?wd���IϞiE-�6��ͫ�n�/-D&�����RѸyIS̝�I��ٚ�C���Qi�MZ�2��ћ�/A,�)�L� H��%蘨K�aQ�-�
{*l�0��j��|��ֈg�p�1�W���YXc#�5$�z� V!��f�]�554h;�,V�e�p�l�2��Mh�c�Uiq'�pyx9� דuʜ� �!|Op5A�lٌq t)��B���U8V�B]<q�U�1t��7-���Y��+A%�ԑbNY�'
E����H����)g��i	�eK��F�F��ҢN�l�����U�z�����J��(��N�A�N��A�8�x�Hc�M5CZ��"
��j}|}� �[�1�LkadU�/���F���������x��캕k�

�	�eC��%�=hd���t�
��¡$V��蛧&V/XSFL8���-8Ire,�>x?����� t���ұ�(� i�t�;l�����	VlX�)��T�F,�V�D�3�@�XU�ԟ4&,�X��ģn8T�RS˅SfF�aC��U�T����7�L�X�W�P��+G�h�F���
S_�	�RVu�c�@�g-,`��-�,r�~�
��ޗW�����*8(�"�o,U��iY��9H�&���b��q�r�2��ߕS�����B+�~2���v�68+���7$��}�b����'^b�0��@'Vƙ� �Ŝ'ؚ�R���	9��E��vN$��'�'h&Zd㤌@��1@���8B�Tڦb�5I�l� �uKQ� �r@�3Fɰ��-�.O2|����+ �;T��X��Ĳ���&]�=��2Eϼ����̯M"T�!��/Ҵ���L�$=3�A�b#tȓ��ڙ-]�H �'�Ե�3��+/�	p�� ����ݪ>L ��"�#`�EHB1Y���ڳ�P�*/�=8%���]c�����%V�.Ĉ��R� < m���!lOH4	Ч��	���1�
��p=�G��O��)�CE�	��CQW�Eu^����1>VpL���|)ħT+H��=�Ň���ɋ1�Ti�W��+mIB�RfK�,P��d�Х�<kx��f��	Tܘ��EL	S��[q&V�7�*�/�(s���˳hۍq
~�o��A��q*NP�|sI�A���|l"?� ,bҧ�.��q����Q*���-"$x&e�r*�%��;��J <�0J��R�/��y� �S/��Sm� "z\�fH�+{�pa�h�n� �i�U�b�й��ɈQ������9B�����{�Z�%I�y��$� �R��H��R���ѧ�9C��#�4��λd��=�U�A17]BఆT7/K.%��I�4��iq"��P��R��b����	�6 �ұ���%�(��@�m��y0n]۟�J�O�C��<���.����㙾ˎy벦P�'jX	�'N�*������~̧4�"P
b�T�rrQ&L�6F%p���n���c�3c��=:�K(O�p����j�l���Ǡ|���@T�'�^T�� �Z=x�O1�h=�Ȉ�o�i2Ɉ9'&���0�Hᅬ��xBI�%xnN��	����!ȂmC��I�#��S��O�\���D)�?��-]��i�O�*��4�\��*�k�.�!�$�/�Lm���[��1��7[��7LT������bE�~&�\I�Ü9rX���,,���	�L$$���f݈iopr5䟃S�L�(�	�c���Ʀ��TD�1��ɹ1� 4!BTiKp�/_Z��򤀝mM����1[���I0�<u1�`F��\e	�9@ �B��Q%� !@�ڞ~�f!R��6ʠO���اo'�}�Q*$�8+��$A�%/�	�i�Q; 5��4eZX��L±G�z�����%++l<Z#�D'|�"�G�������x2�W�c������3�!I��:��xRl��DYD49a�Z��8]Rb�[(0��R�Q��h�-8Z�+�	��Kf���) W<��I&�Zy�'���E��3���:S|p�$NP,�yb���%D��W-�d˚�P���y�N�&_��+��@�dtLRJ��yҬ��=���C�k�\T̜��ʉ*�Mۈ��s�$���!˿*�x�r��T0Ҙ�""O d��$;��X�V�!Vkf�h�[�܅��0@o0<��Ē��yw���O� C�4ʹ}JG��*k��|c�*�	n�<C��(8�H� ��4ᚤ+��ȏ'�C�I0r�����	V�P�{���(F`"C�ɺsJ�iq��4$��C�+�C�I�\l\�p%4?�P��'E3��B�I���i ��
?�(�o0@�B�	�=��H󄃗S�l�`b]7:GDC�Ie{��i��<����T�&��C�	l+jTcŽK���s���<��˓�,��6���.�nqaA�)f.�}a�ȁ��C䉆�"=�@��PM0�'�0:��C�I%�bH��$�����r�ݿ��C䉓X� �J�o��4	ޭ�V㆙MPC�Ɋ:��eB��H�rU��IWꇗ7��C�	` ���@S�]�X�C��

��C�Im�$���m��r&i�s��@��C�I)(02#�? #
=	 �R��a�<1�ʏW�T1`iH�t�&Hc6��Z�<1�W7&̈�����Ӗ�2��"Oԅ{ԢD)f�1��ɧc�*}x�"O�Ly&�
q�\$#�����m�"O�=p���8"Pظ6�H��x�"O�r��ҵ�d���n�4[@��"O�%��ДT�,$���>����"O0��fN�]DN�Ä�գP���"O�A���Q(b'�8��J�<-�r�
7"O��y���L���yQ瘞hF~�"O�� �kV�^���Ԧ�/���'�,���Ӽ&Y^�AGb�3�|�Q�''��H�������ȋ+punu!�'�v逃�_-(
�m����rT2�'aZQ !mV=of�ٲDድ{xyj�',��h�!�q�@q�D��]Ϩ�b�',��bÀ�+Ɯ5�m]�Ta�X@
�'v�QR��=?�b�#wFO�H]��y��� "��kT�x"�@�p. :#��b0"O�=*�K K�0���Mƣ3, ���"O�y��dɘ��0��/T�,}��"ON�#`A�8�8=��@�v���'"O�@��"D��Q�P�Bm�
���"OE�������г.��<��"O0Ys��.�4�*t��;�h��"O謂��ۦz����H#_�H�pw"OF
�%ڒl5b��mؙ;R(|Q�"O���0�8gu(E���F�)@���"OX@�F-:J���#��>,�9	�"O5)/*F��7��H���"Ot�$�D/؀��#I�7K���"O$`A��ʥN{Ty4*Q�c��Ҵ"O��A�64��j3�����$S"O�����V�f���+��X�az"OjT��DH-w$x0�ˊI�Qj�"O����a�*w��y	F
\�5@�iI�"O�Q��ȳ-bD�glψ!a��"O��{V�S�HQ��16eQ��E��"O ��@-$�0�Dـ�I+#"Od�4 ��4�$5��%W0�Ĭ��"Oh	���ܬ3���Z����^��0h�"O�8�d�¤p4D]!7�ԏN�~@�A"ODQiE�	������1�y�T"O�,��K�:e�����)U�B��"O&Q��-G�_mR�p�o�?�DkE"O�e�'��
/�фdR�51�d8&"O^d�#Q	�� S`�!9�q��"O2L�%N��)�<Cu⟙M*y�"O��8a6=��8�!!��[�"O�9`�b��Lu�ASo��R�l�K0"OD8����0���B-B7$,���"OU�f�D?O�EKȯG�x�"O�$k�Ժw� z'�LTɼ��"O�Ћ��5}d@ �j
�~m@�JA"O@܉�,X�I��$��
_�>�Q�"O�!�l�.}xHp	E"@��t"OM�vK�Z��T��A/(��0�"OJ���G!O����� ,�R�"O�U��g�R���+�
��02e"OVL�Ƨ�7.�A'�U&��� D"O�xS��J5��x����qp];c"O�qЈ�"_dl�!q�B5y8��p"O>Q0Z5�y i^�P�"�Ir#�^�<A�Gɪp�����灭%!��QQ Z�<)q���.j�Ě"�����}�ǫn�<�c��h���WKC=a��"$Nk�<�r)�X��t+���?����a�b�<9b�ĝ9��1�ҁU�XdZ�*�%�V�<95i��m�
,SF���]�l�rS��W�<�� ؤN�a�Ε�KߊPB��k�<��o��<{�t�B3f�l�R��o�<�����m~��1�b�*~4�,�3��j�<�R*�JK^U�S��j\q#�$�o�<��@H�&��Т"��_���DnFi�<Y�J)rޘs�+ר!*h���a�<�c��AEX1e�P�D��+Gu�<`��9�q"���v���tğq�<��ىakDH�tH��Ymպ��h�<a�H�,Ȁck_�h9�r�Af�<����{պ�R�A�W��\�E^_�<��`U�:� I!D�;
mb���Y�<�Ն�S��5�Ɓ=\��a�P�<�  tj$�G����j�nX�#�ꕂ0"O��;"C�h���2�%d�L�"O�زG������G�էr6�1��"O�=9��T�.N�KC�;��u�"ODa�A�'*)+�HG1� �`"O� IWZP41�,�� �FM�R"O$��CcܟA}���5b�x�V�p�"O��2C	O	9�䡉��$��"O�D�5��]q4"���  �0�i "O��rD.��]��5��g��w�jurg"O��iu��d���d��W��5��"OFX��*;P˒0) dƨH�t$��"O���T���IH��E�]��H���"OT�A�'�������f� �W"OLUP�U��P��ƞb�ؠh6"Oh��s��<"L�EO/��uQ"O�!w��a�4��P�e.�a"Of�	%�ّi*��ƚ�/���"O֡��D>��d����F��"O:�[�D�DUz)Х�C�c	�� 0"O~;��@�	*�����/q��p{v"OH��� �(�S J)'�N|��"O�5�Ԍm�̒獦}��"O�8���	�
��A愧Kb6�
"O^��"��TluR�E]+V�HsC"OF	�,�>"t�T�f:�H�"O|4A�F��8�`���a"O��C�+&��	`A
Ɖ��"O�2'jY�=����b�;�� #�'8� ;U�G8OkF��bi�*��'��k�fS�6��e;�J&^�bP)�'GؐP�d����2�ĸTk�8�'�y�EƜ�%���a�рTsx`��'�ij5 ��]A'�^#�� 	�'��y!�D�D��%�gC�^-r�z�')���e]�x|��E�!E�|�K�'�Z�iP�T�F�
%��"(r1�'X�: ���� �A�NF <j��'?�p�E!�F��x֤�=�&�r�'��̡����o�N���H�7L�*�'p|Йv.�w�pr�.,���I�'���H2OF�;��ub�`��$�����'s�\���#edaP!ǽ%�T)	�' �'��T�R >����'p}�EH�;XZ��&Ú$��X�
�'N�����R}���@����'���1U	�2]��̱T�	����q�'o�0珐�9l2��G�H�����'D\ݘ��G	hr������<B�|��'6	 S��7�hcai��9��Ur�'���@��[|�H�@ E��*�'��k�\�z���y�@�8n;:���'����TE��V�ڧc��F�X�''�A A�5ut �W�ʂ���p�' ��Q,�5TBx��� �.�����'��|˧'ҹ_���
����.VF�(�'"DmHB�X��p����K�:L]��'��-���Ѯ��V�ǠG4�
�'w �)s-\((�����̨(���9
�'�������UȘ��N�%�J��'��`���ϊL�	FFM@���'l.x�p�
�KI���5��J��A��'f8�Cg�5k~�A�DBԗCS�=��'; b��Ua �v"�EE>����� U���	�e9P,��r�F���"O�RE�D�4�0i�j��~��e"Ob���U�u�]+�ؼ@�nQk`"O��Z�'Ьf����HM�Q�Fx#�"O�����Ī{f�X�ǢS�L4(}
q"O�	���.�
��ᓿa�-�"O��R��ϖU&`��.�w���;�"O65@ୁ�����Mƻ[�z�A"OZ�2SN�&�S���b��<�t"O����Ď0N��=�V��ߐL"O���e�,$S��p�BR�U���"O�}`'a�VerB&T�`(Z��"ON���zgU� �\��M�e)6D��R��%��*��#U/TC�7D�h��mˆ/��ёE��:����3�3D���%��n2��Q�� @LK0D2D��y�O �-��݁p�0��3*3D� ����,N��!����V�,S��1D����ו��}�sDŻq�$��b�8D� Y%�џ(���B�
V�=ci�o7D��iEe��Yg�}��cT
B
�y�6H4D��(��$EF��B�ҳ8<$���4D��%��-�pXy�喨B
&��Ua)D���i֪&-�0��W�Y�0�ꇅ%D���o]�k��E���$5�2�/D�h��ZS��i�mM14^����)D�82����u)����:~�j��=D��	��AX�XC$�B.Pː�&D����#�9GԸ�GLB���m&D�`�F�E0sƚ�:T��Sʚ���.8D����A�Lč�ŋ8n-�}Sa4D�<s7ā�D���W�(!�L��g&2D�TyvN�}Y�ugD��\���a4D�`��J��r��LI�~�{u`4D�$�q�}�z��K1}�:y,2D��nփ(�d�ƀӅh9P�\�<aB���]����A]�H�k#E_�<9Wo٦��x�ehS�P�[�d(T����T�0���C��[
my��c�-D��Rp�ī(g(l� Le@�&�6D�0��=)ZT	�fؑO;q�L4D��I3�J�r�.�C�x�ܬ�gn9D���Ɏ&|�qA��{���l4D��[�� �0����8�n(RPB>D�H
�b�U�ؙ�Ǯ�3Gu�1�9D��r-_��&�J��\��@��(4D�����(i�`�S���y�<:1�4D��𩂰 ʥ1�k�<rc~���1D�8Z�#�	l�B��^�D�D�* J!D�����;	,I5�\"4���ai(D��� ��vZtc���3�~p�$3D������1]^��"A��S�Z<�-/D�����&����߬ �઒�6D��U�ý(\�H��F0�Mz�	5D�D��:w���ڕ�$H��m�a+3D�LA�J�qifl���Ԡwb�����,D�4k��VB��8�2\� ��6�)�y2.�t�R�!���
Q|�49f����yBě�2<�d2��$��+���y��A+8�|3��Q�@�(��e�.�y"��X/�����=��ZR�y�#[��0��B�_��X� 'B"�yҋRHp8Ń5怟Nh �
`I��y"��!�(\8����k�>��W�Z��y
� �@��,Z�C�a�!Տ��"OBuʲ�(	G�$zW@��Aڨ�Y�"O�قG�W=C�V��n�>�&Mr�"Orh����/�L$��J/V�&b`"O�	��/eN,�bi��!A"O8��W�0k��a@�A��	��"O*)�J��~�*��ة=�D%3�"OzH�����ּ���Ֆ���9�"O^�ٻz�D-��Ò�y7��s"O�m�W��r����"�7�l�&"O��*wK>w�4�2��4e��s"O�	�EV�&\��S >f���""Oh)��@�J8�H�� T�k�@J>D�l��Ox��1�!G� �p`>D��*��͚`Y�IQ�E�+� J'<D�L��)�D���Z1�7@��Y %�=D���g�#LdT�-�:��19D�E"ǐ�>�#$/0?�fm �/(D�X������|*p�G�D��*#D�̉2	Zc�NL�&�U)�4��;D��C'��lJ���d��5���� 8D���c�P����$��$�<����"D�p���r�~�G�ܦ�0��@� D�����з
��H�D.�Y2Nł�<D�t �	 @&=c��!n`��;D��Ѥ��
��� ���}+����8D��Z�I	�>=|��w�Ɩ ��P���*D�d
t
�_L�uXrB9^jTsA'+D�Ȓ�f�O{��aPG�2 �����&D���'����;�GƀemR`�`�'úi�@��@�mC1�C�qU�Ш
�'�.	x�*�^��p�H�;��1��'����(oȬ��2�z8X�'�^�Ye�	pvLB�}cL���'�ȥ qo�0kF|�����	r�ʸq�'��Qg�ϑ$5����#�0l�l�	�'}�m0�ݸC��5I꜡[�`��'��qX�,\7RNa�3-��Rs�(��'�>Ta��-D�μ���A/� �'��adjF����	9F�ڥ*�'��("A�+.�Z�!�ؕ4�P���'T0��ub�n=R���.�A��'��X��KL8Wh)#q���/j��9	�'0�Y6cڂ�j-+�`��Mu`���'�$q:���-�uQ��.k���S�'; ��>9Rr�+�74@&�	�':t�J���Oq�L 4��\�T��
�'0ЭS�C�w"�iZ�Y�F(\X�'��[r#��^��h���4�@�S
�'N�
ՌNmB8���E E���	�'h�ڢ/Ze�탕�>c�\�	�'G��z��_��A�D��6�@8�	�'�ZH	Q�]7v�y�pm�$lV�
�'�W"�+M���0�֣%S��I
�'��Z���r�N$SA��;`0	�'`y���_	���8�ݑd�J(��'BU��L�&/P8��#�� $�0��'�Tu��� �n(; Ä#$rTE��'gd�yG1?R:ҧ�7,�JIj���ɭm��P3��?Z��bS���F��?�jI�?E�D��-xHKg����`�w�֨)�Ψ٢��4t�P+�Ol��
ç/3:��T䑠Sbڠk1�E����"�ӯND25�'"ZP��[l>=3b�	�0y6e���[� ��m��#����~��� 2N
hф��iʚuI �P�Z!����F9g�����0	D�*��Q=NAh�{��O�- A�Ե�Q:�'		66�C�N���HY�p�X%sy���pCc�ڣ|�<�� �����-�ZH.܂,JEr�j��8���w�P��@FR�XF�cO(<��̬//�����4��*O�82�닪,��@C{b����2ض��VI�k�����ŀH���!�M�m�vE�f̟�Z^���O�-r֧�&L�s�Ьtӂ5�D២g|�yh��λ'.
�B'��0|�ub�$�p�z��"�s��7]&L��*.G(<"�a�1F7�ӺȖ�����Y/���8J~��Lə|.X$����Zh�Vi�O>��B�Nb4/�[?�(`���@�|}(D��F�fˇ�-r���#}��^9�8��	1?7�y�*�o��_T�D�L���EL#iz5���(�����,6D���u�^�R!B�����6��b�c2D���¨�D��X�L�n�	�0D�Xr��Y��2B�&��a���-D�h��I�%���|4���b,D��b֨�40�ف���k{�uP`,D���.��o��l�5��>2X�e���*D�8KeMJ#	��)P�/M�,�0�� 
(D�Ѓ�kP p�
��C�ё��%D�8)��Z�W��̨�d���uj�h"D��`�̾k�BDH̙"9�$��>D���CE�,� ϋ��0��G>D�,)����B��p�r%��_5�]C%�:D��؀H,iTt����w�X��%D�((G��$D.<�yG2���3��=D� ����$2��%
�*<NGZ���:D��RE�Q-;`�2F)�&Y�i��$9D�ha2�Fp��Q�S�,�]� 6D�l�u$�	;_��ʅ�V�3[H���4D�|�a��Bv��Y3էn�%!�=D�d!�ې!�T=�@�)���e.D��
�-�)n^�����"7z�D9D�� D�
��m�Rϑ�Y�)*�L8D����'�r�p�.W�z	���5D��Z"#m��q�ꊺN���c�#5D�\i4��X����!���0F.D����D�@Q�4jn�����y��n2�	Bb��`�Ԡ�OB��y���!LZ�k���&��i��y�ˡb9��զ@,*�H5�լ���y"�^�d��I!$œ�m��dz�C͇�y�M�3r��@p#V�P~�	�O_!�y��ɖ����T\<Cl����B ��y�홠$�(��ެmh�����
�yrc84��/I�<.�yB����h*� ��~f��7,Ʊ�y�"<FH�m#V�Դx'^�PsgX�y��6|��t-�>��ҏ�0�y2��dpI��7E����,V,�yBh�8��y�L�(`���)�y�Ě	N�hh�s$���FaÃeǇ�y��� p�R�o�k��i��T<�yIT+P�a��m�6XiC;�yr�%z�ݪ$NO<eIY���yR�&w�P(c5�
�����(�y"�Z�P��9�7��A)Ue��y��]��e�$
?]��h;�ϓ��y�J�+j�L���M�� .�3�y�9��y�s���M_�s��2�y�ژ�8�a��syJ@�bЧ�y�Ν;ed�c��)y'��kӢ�0�y�f����� �\���I��yRޮT��H���/S"�0H��̈�y�(O�L�h�Y�.�v�������y�X"-�
ِ�(�h���5�N �y�DE >W*񡀉3aKP�c��y
� �`�k',Tz��B ¶OY���"O♡�
�F�T��lzX*�"O q$A[�m�<�x�KVW�I��"OQ��AѪbv#��۬M�`���"O�� �I�u���x����J�9�"O|h'�">�Y� �?P�6mV"O:�+�F�F8x}� ��<4����c"O����mI�VD�#@ϑV��$"O�Dp􋎁o�vPp&ņ�f�b���"O^]i�
 g*R��6J[
7�Vyy "O��(&�F,>k*T�q��t��`"O���vEHT	��!��b��"O��[����;�X�O�)�*�Y!"Onu2"矆"4�[D ��1E"O�T���c�.`��.�/�Z[�"Ob��1�3S��`i�휀j���q "O�p��JNsn,I3�+A� �}�'"O�m��*�-L?R���J��`4��r"Oz����'��K�iͷc$\�#"O,���Ď-h�Zi(L2,]�"OeH�<q�h`	Ї{��q�"O��b��فd���f�ki�Js"O��p�ɑ,r8���EWZ��y�"O^$B6�4��7�{�TpA�n��y�	��2 �G��}��$8��8�y�N�Jmzi%�R!q�Z!��K��yҌ@y�0��?}T89)W�?�y��?�Ш%畐&�@��Fͷ�y���2C��(�M��+�l�a��O��y��փ�F���V�[�Y���7�y��ѝS�h� ��Sr~9�ˑ��y��|l��O©Rf @+W���y�oU���X�!��|���K1,P�y��N=)���!ؙt����+���y�&�,dSQK%���d�J=�cd��y��Z��RTׂéc)�`;D��y�<7�Š@�o;� P��ٰ�y"��'R{ �"O\*h`Tm�0���yb'��1���D�[�
?6=�-�y"�ɳP&��'��r��[t���y2l� p��D��	;.(����A��y B.=�)s�؃��k���;�y�)&	�ڡ���|�x���y��'4��wH�/D^����� �y���*[T���ʝ'��0�*���yҩ��� B�A߼(�,eKg�y�D�-W��Š�vT¤��Dۨ�y¤�up!ZDNY%n%�������y2Ѝ'f�Z���Q�T��׀ʜ�y���d�Dظ�N��Z���p�"H��y���5(�洱G�Z�}����)�yb&�7M���x����M*z�S��J��y���]������R�tm"tY3��*�yr��fn4�*��Zj��Qʍ�yr�O�~<�R�R�iuz���P�y��4k2f5�Z/ZZ¥9�Q��y�j� 3�f\��ҫS�FHEI7�y�/14)����"Ҭ�y�X �y�)	�j��P&H�+'�d)"O� �ybN�S,��mǕ5I
���N��y�`N�o��RC:�V��P!Q��yB,P2�-���.�̺G.E�y�B��yG���I���"�,Y��y��C�T�R����tiǭΊ�y
�  �PRE 0V��=�A�O%��� �"O2!Y��jE`D`]�1� a�"O4ٻ T�s~�ŨP$UR%�&"O��z�g�-T��R'�,,��	0�"Ot�	!�L���ڲ�*o����e"OJ}{w���1v2�cŌ�z�#�"O���� C��MBS+E�]�p���"OT�Y`�S'Ini(AK$j����"Od�w鉤,�l�x�\.�=cE"O����~X��bK4`j�%"O���0�����e,�S����s"Or�)�!�"�<`��K�(�)��"O���k'�R�#��3?'�x22"O����-�;�F[3!40��T)�"O,����֭M��ܳ1�8N�e�F"O�u�f�Gw�*�W*`G�8�"O�P8TDQq�hx�&p؄E:"O����)���
B�Xy/"M��"O9	�-��P�Bdό�Z���`"O�-P���q��]W��"J>�ٻ7"O���"�
R������ħH���"OJ�B�^�q�^�b��B�a��"O�H8׮ޓ�zK$+͒F�j���"O�mp��G�(Ҍ�0�*� ƈ��"O�0K�֞@�0aS���'��R�"O��
�C��k�^$30 �-O2��"ON�!��..V�y1�т4���"O�t����0iZ�q��ȃ���:r"Oni&�ɺ6r��l�>#|����"Oz��Ӯx�`t%�:Eh�4��"O:�+W��R2�TA���"в�"O��[�FS�<�hA���5�2�0"O����E�.W�&p�Fokd|�`"Ol���Ș�sv��:Eejإ��"O�t���]*cAbX�0�X� �R,ڥ"Om�ԎM�ޡ�B�\.;���W"O�qWM�^M��#DJ�
�̓�"Oڌ�c�_�+`��g��
(�a�D"O�d3VAL�6�޸`���x\�"O���`�I�p��C���-k6D��"O�P�%�3(�n�yT�+�̴23"O0�A�^/];�e
�iǌ�T(y�"O���ŅA�e�z�5)H�x����"OZ h���>%*|x�e�|K�"O�Q�3A�4!���Yt�D�@�0"O���Q#��0�*�j�!�D���Q"Oİ��@9$��0�@�N�Sb"O q� �j"�8���;�
95"O�8xST��\���gJ*;H�y�"O��0��O5zmzuhT3��h"O�Aӂ�q������JL|rb"O�5FOӝh��XkT�*+=��3"O��1�,�j���Q��9I�dYr"O��� ��y'x9X1�!a��	�"OF	2S�._��a��8����"O>P)B"�TrV���O�.h�B"O���u�A�=�Ц⍷|��Hg"O��Ӧl&>�쑘�o�v|5�"O:�˕�_�M�L�Z�LK ^l�r�"OV"���'u>Y�c9}@.I@�"O�DAg5zϦ!*�ĝ]=�[c"O�| �m� ceqH�L��-��X`P"O��nďORTa!C-��Ta�H/D��Sg�ʹd�6�ZB�0� �",D�� ����% &��W�C�:TN��"O�1ȣ�
=5�(�� ��Kd�X�"O��CԭL��  �bL�d;�)��"O8����ޓ9���f5$"� "O�Q�fK�y��M�2�q��T"OT�K�4 t<ʴA }RV�˗"O�A�$�D�,�D�
1��'>c��F"O���픨3]p@Y!�]�(@""O�B� c�=[�I��e�����"O\���j�-F~�5��Ω<�eie"O��ɣh�H��PA�(p�5i"O���vO�4�N,� n[�&�6E2�"Ot9: ��,�cL'u��1*"On��GC�#�@�bKV�glh�:�"O�䊡�VEx$���n\�2r"O�X�A� �r�1�锢xO�`C�"O��TH��[a�9��_�9�J�"OP�	@«R�$D W%��p 2�*�"OZT���PI��Ӗ2� I�"ODs��2/ � r¬*,\��K�"O8<��K:K��+"%E�Hka"O�yj"��mTA���W�0��[�"On`8"/S-^����v �'h�B�"O��3�   ��   3  �  �  �   A,  �6  3B  \L  �V  �`  �h  o  _u  �{  �  4�  w�  ��  �  E�  ��  ʭ  �  R�  ��  ��  <�  �  ��  ��  ��  ��  ��  '�  j R	 � � A  Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�� |d��"O
`�(�;���8���-0��1%"Oj4��ND^[��"3/9�0|H�"OB���H��*�ʞRy=a"O�味V�!X��!&F�:J�$���"O,��a
���C�Ą�M�"O,$3%o�-���p���+Ն�:1"O��ݢ1����`���y14]2��i�<�6��{_���c�H�`�fX�$Kn�<��A̼VI�xR[�)�Ć�pඤ�ȓA5��('nߡ4�� �)˩%� ���,��r�؊b#`T�eT09���ȓ!�b��g��}�8�F��-? �ȓ
K|m�ș�VṔ���2�%�ȓ"R�X�j�4JN�1�˘X�i����̹	_�jZ��1!g��zܶ��ȓgil,*�J�
j�Ne��i�J%b���f	�(U��:���G��$Y^م�~r�� S�%T"���k\�jx�ȓ|4�1�îJb��@ӵ�ݩn�V��/[`�"�v4�R�!ʎ<��M�ȓ`:��z�ؚh�J�Z��$HY:	��H��p�m�C1��!��B:��0��EnjZA V;9����J[
2���	��4'J�EA�IVW&��~�(aZ��ӹ�>� o�Y�|�ȓ�f�A�
Ο7�H��M�$�����mޠP����/���ANXo*�ȓTv�����{ ��-7�*h��I��sB�8�8���3����ȓNe*M�悡;������X�o��!�ȓ'lj�#F�m�+R&;�|��2)n�C��0S4���T:
b���:�0!��e֊��)��ͷV��,�ȓ0�&�8#���� ع�L�����;�P�AFd���,w�6d����?�ЂY��)"��Q0�]2�K�]�<!�aؽJ��ab�I`x��c/[�'~�f?Ojb?)��"Ln{��ǺjP�՘�,<O�"<AvF�:-�D%Q���8m&��� Y~��)�'S  Yiϊ"`NQ3BY�
G����i��L�ѳF��Y:Ԋ�KA����l���׃XQr�[���;����<A�U�Tq�@�
|.�N�9c�9�ȓ��Aq�G\�e��T��o�-H�<l�_���hO��/w\AsB%
@<iR���!\�C�0mT`�!S;24�񰕫J�{��C�	����c�~o�%�pfӖOUpC�I���y࠮л'�T�5 T"8�t�IW��hjR.��O�z���&�� �Re�3�I����@D�;E¨Y�bc =��cB1D�`��̞5
n�Aң!�Lo$�*J϶��<��O̍�d F�4���Y�gO[e�n�Ey�|��EZ!X:���tg�:^Rq�ĉ[�'�DE�����_�R��q��g$�6���'���F�Ou��kOP�l"�����a�
��'ў�}҂-��E/v���� �J}�!n�V�'�ax�lZ)	��$	,!�A@�)��>��O�=�f_�o:Q���T�*`�'�'��%�O8�R�6	X,��e�m��jD"O<	1GL &�����D:	��Bq"O�y�O�\>訃%D�"|4R�9O #<	� /�g�? ���5��������@�l���JJPH<����UJ�J'�f��RM[�<i��"Rx@=je�`����2ˋ`�<9p�GI�yZ2��:1�Ȉ�dK_���hO�C���@-3v����	�BĈI��PT�JdbQ�e��	0�պR�d��-V	�tB�!��,I�HՀr��(���G�'���q�P�_I��P��	2t�����'�zH�Tf�ⶅ
��y)�Dj�O��=E�B��\���ڧ7�*d!�i�-�y2m�l�b���E׃=NR��Q�	�y�!��43��"�$_H�BQ�H�y�鞿e�脙�KݩSZ�$� B3�y�,�3����G4�L��pc���y��B�9s��s�iӜ��� %��yB�0s��.V��+������<!��@�/<B����2�Am�&3~铘�>���Օi��l�b�6}�00Sb�E��hO&O^@k��l�-��L�� �L�"OJX6�8U����aZ1��,Z��	Z8�x�3���phZ4��?m��s3E&D����ua�mD�c �  a��K!��T�e2�op����
 �D��J� m�P�I���ٖ$�>/�����IJ@v�13!K1!�$Б�K(D���Ǎ�(ЬY����"�%D�����<C�H�`���JI�娢�"D�4h��K�#�`�g*i��Xjc�2D�4��*_�7l�x�!�d�ȣ&�p!�[� A>H�$�; ,��H D:mK���.$2�I���9�Ȅȗfм�y��nIFA
F�D��\���'��"=%?m)��
�?�irQ�]o���;�C>$�`�����~�L��@��g�x�CD���yB���0����Ra�������y�Bԯ!��ĳFhNZ�`� ����y���,jB�����CS�<x�%K���	9�Q�t�~�#��ON<t����?*��q%]t�<uN�^:p�QRGJ�Rqlqa�`L���=I���5��-���?Yq�%4ɅJ�<�% [;*��Ҥ'�!��\8���_�'$0���MJ{�$��J�>��0!B"!�P�L�X(@6�Ƚ1
�	�f���!�Д]peI�T��m؀膝3��p��H�xa��ߊ�$#�KM�k�!R"O~q�b�G�&4t�P�
,��H�>I�x�V܂v]
��0�t�_06���A4Bҋ��lfpy ��D����*�
-C�c�+|��%9���p����j�'/(TYfdUJ�,0��X�3=��Pٴ�Px�j�X��qa�=�8�WM�p=��}����c�8BGB�,�׋���� �OD��&?2a���M�@�xl�"O:,��.9�Ta��fq���"O�ĸ�*�Y�"� �#(S����n��D{�O^�9��"l��Bc���(��"	��hO��H�`٦f�������0�P�a�"O ��� �q�T��>��h�"O�ᑣ�ݞ^��5��@��E�4� �"O>�R�	��4�I�FJ�'�v1��|��)�����	�ӏY���Q�!��"YVB䉕EQ��	!!H����+3!���DB�I70���D�*��Xr�I�ls$B�ɜF�bX9�?c�Bp+p���Ai B�)� $�B���9TNqr���<;��;�	b��<��z�Mϟ#( ���.��ȓM�b5�c�҄[�r�s0
O�	Y��%��F{����$`J��Y�Ǝ���P��2�y�c/bۢ�kEa͐o�>�CQ��3�y�Z/N�Pa�T�͊\^��������ܑ��>	�r�Y�[>p ��*G�4�2g2D�3#��<Y	���c��2� l� /.��X����Mc�`]:t���9$oX�z�z���M[��?��5,���Q
L�vᑠ�	M�<�RL�x�D���-�h|	� �H�']R�S$ʅ�f� ���EK�|AT=���>I��hO���EPĂ�4i����q�x�i6�x2�7�S2��Ëi3V�;ã��,}y�Q��y$�& MF0+3%V�LQ�ܸ��Ѣ��3���IBܓ�~��4�r��[`o�e�$��+D��a�"Or���Ѱ;�	H�I�[������L&���ቆq���� ��-�Cʏ[�����&ғ#�и�
�8]`:�v*��y>��>��HSX`xD�	�$K|��	�#P��UE|"���!^b�kA	���׀0f�xB�	�mJ~�xa��.�8!dNX�gHZ"<y�O:7�p���'/�i�*���b��H!*f�i8A�
�R!�D�3E����g"z~v0���w���hO��(�ǮP.|}XDbS��)rú��'ۛ�i7:'�8Q��>C�����$��RX){�6O$6��d�S�Op2��!d3�6)JA��$S���1�"O��Q��*�P�ig����4"O�4��;buVIW	�}�p���l�c̓�~*�.����_��xm�+ѭK��|qRIU.~�:C�ɽA�v�Y�A+u;Lp������>y��$�3�� I��̀Z#�8���yR�Z�xG��9�c�4������yB|��M��"2��%�U��yR���8�l�J2o�xz�!�%ͅ��y2!�95�0�B�䕮u�)�����yB���~d�c�Z�,��:B�yB�.m� 3���Z��(2o��yb��,>Gp�ѐg��A�i��
�y"��h��}�qǞ3N%؅����y��a�|d	"���.$h#����y"Q�|҇�^��(+�	O �y�(әl�����픯?V$A��y�Ǔ-8�h�Z��+�P�y�v&�0* ��=��`ٲ��	�y�*+H��S��,	��݉�@��y"NC���̊�2�]�V���y�\��t\�q	С'����r'W-�y�	H��[�o���^̊����yB��,y��B3Ecu���y��L�[��XQ�K�`��j5�֫�yC�>�̲��*!^u��Ր�yR�e�i�"�G����ᲅ��y"��[�"�0A�R�h se��yBΔ,������E�0�P�K�& ��yb'�Z�[ W��W0��4�y��WG��{QI� &vR��3���y�Oz��o�kA��wF&(!���K�~�׮χHXpȃ��6�!�I�uBU:�C�$S�!Ib�^'Y3!�(Z��I����,1��"G!�ĀWô� T�[�~���`VED�O0!��)Z��U떬�8���D6#!�j�����2H�f�I'��n!�� �� �'	 �����فz<�+�"Ob� �"	�W5X��u�� "�����"O������Bq���v<��"O�`HwE�0�zT��oݝ7K [�"O��+��1ExH��� �QFD��V�'���'���';�'p�'p2�'�$�u��"�B���Zo��M���'���'���'
2�'�"�'�2�'��h%m��m)h��C��[Jy#�'�b�'r�'B�'r��'p��'��;���V2��c�&(��2��'��'�"�'Z2�' ��'��'fL�V/T�m��)�2���Kmb��'��'�b�'�"�'���'42�'�ذp"�S���C�jE�p_��'�2�'���'���'���'0R�'��8+H��L�h"���z"�U�G�'�r�'���'���'�B�'P"�'�"�/H9i��� GW�I�@��e�'���'�R�'�b�'��'�2�'�Nm��-�|x0�e@��r�\0�'%�'�r�'��'��'x��'+�	�ϑ[B2�b3��;yN����'���'���'�B�'TR�'sr�'��(qff 7z�V�*V�XGD�Y���'Y"�'>�'���'�2�'Nr�'W:�2D\~�y����ą�b�'.�'5R�'���'J��'�����^r2B�J�吷L�X��E��iy��''B�'���'HB�'`Z6��Op���.	��4 &oX�L�䦵�'r_�b>�!F�f�]G���P䒑:�h���؏-�ء`�OtEmޟ�&�泟�oZ;#`
��OL�`_�d�C�>`�;�4�?iEē�c~�'aĽ(çX��ܤ��H��������ksk�N�̑��D�O�ʓ�h�^�S��Qu�y�`��*��lI)�����pi#��?=&?������gc�#��t�h�S�^��v)�x72�i���<%?��!�T�J�|�	szI�%��j��s����f�I�[R~-��,;U�ʕE{�Or�S'~��*��P8L�����p?�.Or�O�o�:Dc�Dr�%�YΦ�25�� Xdp����x$� �,Of��t�,�Id}KH[��Xa��Z0Ѯ�%$�����Bg��9�̗m#1�6�	FI�t#`���4 Ԃ��"��c�&�r�琸6ʓ����O?�	~�d��J^�x?��QE�M
z��M�O�r~�$s���$2�4�ΰ�����-,IeKM�{ Hе�O^�dz���dܤn����ᔟ�Iu�����A���<�LQ
��V/0yaƪ� /�(&�|�����'�'$2�'e����)��ԉdi��R�qDT�h��4Cj̀���?������<��I����ڀK�*QP��b��B�ɶ�M���iN��� ��㟒�IK�"�@��'B� ��YR�&J��8�'� �?��d�%vj�D�Cc�L;�h���%��뤡�	Y@ak����N�(��A@�9�|m����=eJ��W�(\Y1CHԁ2���݃My��I�E�
����C��#Y2�mx��:@���5i��vG6U��r3��@���L��OZ�˱H��v�#dn��m̾ds�Ĺ�l�Q 蕰E4:I*B��@h��åq��;�!��(�k���|���{�a��il��kA�O�,����t�̻-	nz'\,O͢Y2�e�A���l��Z*�IV�b��<�E�Ӂ0rRy:&�P���u�D�g�������j�A�ٴI����`�� �f��������	��i���'RR�'�bQ�L�IZO|�S#�\|c⧓���$:p/���*!��4�?���?�����ċ�H~�l�ß���5&� �Rs�Q�P����tDѕ�M{���?�������Oth�*�<��'�ĚC�^�=�D=����G���`ٴ�?Q��?��O}*a��i�R�'z"�O��,F���l,>��ѦI�k���a@)bӊ�d�<A��!�r��'�?a+O�i�:ܣ���"i2��U \&X]��4�?���P*����i(��'���O����'h���G�=@~zxRoS��<͐�>���&_�dy.O���|�'����Q���2�)�E��ه.d�zxP�������	��I�?������I���j�AD�c L���F��عhF�˅�M�GL��?���4�ڒ�\�D`��8@ՃO��昳@�k��hp�4�?���?�DQq����'#r�'�"��ug"
�%n�� F�6�����M�I>�7��<�O{��'4��d�҄"-�oj��:E��m��'��QXt"m�L���O��$�On��O����^��	�cmԑq±�ԃ���	>�J��?1��?����	Ʋ)��c'n�n"�qQW�D�H�&�� G��i�������ܟ�h���˓�?y宒�n�*���MN@-�d�ȗ�������OR���O����O"�Z�q�D#^N� Q�ؚj��X(� ��M3���?Q��?�����d�OB�4����##I����EO�V���EMp}"�'���'k��'\X�'df����O�t2g���bV���D�
O����q��Ο���]y��'l�U��Op�A��0�/�l��YБ�wI��l���(����I=�*Hh�4�?9��?��'���޽ �V(s �J?:N�H����M������O6�P�>�`���<��Ł'm^�H[>\`��N%Gt��R�}Ӧ�D�O�aSdW�9����H���?��󟴘��	<��aK�i_0.���3�����$�Or�� �O�Ĩ<ͧ����m�4���4aU��V���>�Z7�@	mHo�ߟt�������?���ʟX�� �Ԋa�߸mj��3�b��>���bڴ���/O���|��4�'�b�a�_6W�):��H�y�T��bh�
���On���Xޤm��L��������o���qSÑW�x��"Ѡ&�,6�<�1,����|�S���OS��'���  P�T!��-Xڌ�Fd
a7L	��i�r+v'�6m�O����O����Q���O�z����=)`��!H�S'U���Ѫf��	��X��ȟȔO��B�H\�!u�@�6�X`8�+�g�	 �uӌ�d�Ol���O@��O��������
D���H)�N�Nb�������Ty��'�Q>���,t喀2�4lP�操9b�a`W�D-n�Y�E�i\��'���'�2Z�0�	�Pr:�ө7_��� U�]��I槉�hi�y�O ��O����O����a)o���<��:{U~��G�$ŀj[�b���4�?���?�*O��$��'�I�O��I�qh:��-�
PzBACD�D6-�O��d�O���Tn� yl����Iߟ��� S3!F�V,4���)0�K^Ȧ��Uyr�'�j�КOUb\��sӰ}�rnލAM&�B3�N�kYB̲׺i\"�'� E��GkӚ���O�$����OD���d�.�.5��J%t����mNR}b�'T����'{�'i�5��O��^d�5���\�W%�0��ES�&Yl�Q�lش�?����?�������?���o�ܰ2J�~�~L@ᅉW�<إ�im�`Y��'�ɧ�ԟ�$�'@FAP�@̍3�v��#=�t,d�ӄ���O�D@
w�|�o�П��	�����]>Nh-�b��mBCiBpF�6-)�þ/��?a��ß(��Zx432�� ���{��ۼjHμ�ܴ�?Y4��?�&�'��'��~2�'�E`uEZ.>�1��Y;\k����4wSP��@Ň�<)/OP�)�O����O���ү�i�5�-^dEi�jJ'cb�q��OƦe�	џh�	ڟ�ɨ�v˓�?���3�^Ȉ���)2>��	L-ZY��?����?i���	�O��H��˦�	%B73O�ѳ#\��40���D�MK��?��?���$�Ox�"7�����D��u�T�P�n�s2������I��p�I��|��ɟ|a�O	�M���?aQ��,�����0Q�`(؂Ò*$͛��'�2�'��	Ο ��,r>���R?�n@�=j$��M��'X����f��i�	ٟ����X*tH�:�M����?9�����/h9�X@bM�D~*|�Qb�R���'��̟�rT,s>��Iby��M���ɤF޸bd��[-�]���G�9��۟�R"M��Mc���?)������?�5)G�d}R3 ��0�vP`d��G���ڟT��I� ��Cy�O���O8�n[�mZ�zJ� @,T AǼi���2�`�x��O����$���O��$�O����N�4��P8Te̡>HH����%�ݟ���Iy�Ot�O.ҢGZ��CXB���z�F��ALf7��Oj���O�ƈ�Q����I����i�y��b�+D(���.j�!"dap�T�$�<���^�<�O���'D�b%� Ʃ����8��� J�7m�O��HAaA��a������IƟl(����ɯ~	�PE@1M�a����21��W�~͓�?���?!����9Oz��[���`΋05e�� �EކA �$���ܟ�$��'U<`����6���՞qE@�Yq���'b��'�R_�ċF�ć����E>Z���!"���d)n�#���3����O���9�į<Y���}��%R�(v� �0M c	Ʋ��$�O��d�O�˓I4�QӐ�t��I����������H�B�7-�O֒O��K�@P�>!�LF��)���n�B�R��5��ڟ`�'�1&l/��Of�I�qa��k���/���EAS�)��$���'������T?U�KZ&#�,()%�=8��	j�`˓q� ����iW���?��'<J�ɮ
��ѨO]Px��#��>6�<䋘T���Oj<+�.�e�u�qƫI6E�ٴ/4����i5��'P��OX�c��+F�N�E��
��(������MKs o����D��C�N�[��5A^�����r�XoZ⟄��˟()����'�B�OlmŭC?��=��ϊ���-���F���$�O��d�O����OBq��*�(z���;UC@0S�LЕ.^�����t(�}��'�ɧ5�ć�L\�x
�Y��t�Ī����D͙61O$�$�O,���<q�O�D����بt}���g�11Ӭ<	��x"�'��|2Y��*��Z�<�&�� �;��LR���'NH�c���	���{yrb�/Mw>�.`�Q��ݻ`z��P�JT�'� ��?���䓾�X�?5�Ƀ_$&��3OJ6!���)��j׮��?Q���?�.O���դQ�S�I,����³}�J�MS.in����4�?yO>q/O*�����4N�"a탥R�<�����&�'lBZ� ��N��ħ�?���$N��˖!Ҝ �
���/��)����x�W���5��|���3k�a�6�H&[���1��lR�v�'�b�
[��7-�O,�'��2��رdV	���F�\�(����vndӎ�bbnDx��D�������2^)L%�B��(�M��/s�F�'�b�' �D.�D�O 5HfÆR)�b�ҧt�p�2K��Q��"�S�O/�G�7o���h4�D5}`����s�6-�O$���O�%��n
B�	ş��\?Yŏ�@�`�F�+_J��c�|�L���<����?��<
0zU8N+00�@�C�y�`U1�i��J�!�nO\��O��Ok�6%�� �e�_M8�C��P�E@�ɿ0c����럤�IBy�oH�5�ra�$N�C<h� �z��#�C7���O$�$#�Ĳ<)����@{�cУ�?eJ�Ѐ�*0e(�<���?9����L3T���g�? ���NW;Ul6 y��j����Дx��'��'�剷O=��m�(ըb	�ly��[�NT���'��'��^�ܹu��8�ħJ5��rDԂ�-u��ELU�is��i���|�X�pɇ�?�	�:�ܝ;2NVqf�,5��:n��6��Of��<�׉�2�O�b�O�܍�7͒�s2��i��P�f6(�	b&�ĵ<�6�Te���	T�b)�x�'�E:g�q��B�s�F\�88%i/�Ms1W?����?�	�O�I�@��r��B�DJ�f��u`�i�	�dl&1�?ͧ�?������crD�S͋8��������q"6�O'�M{��?�����x��'�Ѐ�!²o�50���*}4 +A�}�6p��O!�i>%$�����nD%)D��En8��Ŵi=<,�4�?���?�1!K�!�'Or�'cr�!G¨1�䀤"���ke�߶F�c�X)P!8�I�I����l/#���sת^δ�4���M���	.��5�x��'��'�i�ai��G�e�.�V+�]����'��>	��Ph̓�?���?�.O����ŋZx�yB$%6t�hC$T�U,�$���Iȟ�&���O�����"p���g�J�h���D�O$���O�ʓx/ˈ����,Ϻ1�vi Ӧ��If&%hg�����O�$%�$#ʓW?�-�D �`�08BC�+_P��'7B�'U�R�0�D����'xh)A�/�+?Ʀ�0w蝞AK*� ��i��|R�'	���S�5)��HɠiQ+�^�!�4�?I�����6�$�%>��	�?i��ב6���I�"[<T�:'�����p>ag�B2���y��ނ/*X��I�U�'���(�f|Ӓ��O��O���]����H�le���1���u��nZ[(<�sAU�u�p9�e��2פ�Bu���������M����?A��B�x��'�2���)��:�aJ�F��~/���E1�O��P�b�ԣ7d��L*��#CĲk���mڟh�I�[0�����?1��~�* �s0��!��X��灅$ʰ=q��?���,�p8;Í�(�*=����'n� �X��icB+C< O����Oj�Ok�S�>�z�+���?�t�S���t�Iɟ���Xy��N8����e|"%��=+��U�c�-��O���*��8}®ٮY���#4㏟:����cn����'�r�'�"^��C%����d+�'@��\�獗	�pY�B��3���?�M>�.O衱s_��E`�*���hA�������>��?����P�)"X�$>X��ѷ>z)QE�&P����K��M����䓛�<2�O��fÝ�a���S�Z'D6�ᤸi�R�'q�I>+��̨I|�����gc�+<FڠiV��05�`l36�0^��'k�	��X#<�υ9ZmViP&'Ʋ'٬z���M+/OZMꕭۦ�x��0�$�*��'(�`�2���4��i��)CM,!;޴�򤘭}G�b?�$Α(�\9��&����Cs�^���B����ߟ����?ysM<���5q���M\�sÆd�� =���Ҹi<L�����S؟<���׍ �ّ�IV�zG^0Q��ٹ�M����?y�D6�{�x��'��O@�h�A�fqP��'��و��$
�D(1O��D�O��Y�8Ĕ�#��?%a6��
M_�
Qm؟���͔�ē�?A������$�7��P(�iܑ-�����&�G}��T�٘'���'�W��#!�Z��A�fB�")�43��Q�8�M<q��?qM>y.O���%�X�����rݪ-v��WcʢNH1O����O����<�ą��]��)�&�ɨs)h��I��h��2s��ݟ@�Il�]y҆F�����_�BE�2��)|�xeGN�{d�	ߟ��I��ؗ'�ڱ�/�W�s�e� ��S�yY�j��5Q�EmZҟ�&���'F8�}��N:��`g�'5Daˢm�9�Mc��?Q*O !C�E�A�������xL��D�#Rd�x��Y�ܘRO<�)O���V�~��͕8�@��煛�R���(�/Uᦹ�'����kg��O#��Orp�'J��(�M�}�ԉ�j�{�p�m�Xy�>�O���@���1x6u���O�;.�찐�iy��pjoӆ���O*������%�\�I�of���ǻOf�������4�R�Ex���O�6m�s'a�riLo��S��W��M����?��4-���xR�'	��'V������A}��SE�N����b�"�I�;b�X�	͟��	'8: �E,E�DPq"�W�)��bݴ�?ɆLOVM�'I��'��U���V���R*N�p �p8
Z/�j�e����<����?	�����"n��+����cR�|��d�'�����}��?!L>/O����� 5�DƯ��J_j͊e+�)t�1O����O���<Iu�Z.���g��D�d�c��(Tf	�����d�O��D"�D�<��j��~��ױI���U�N��V]�P� ���$�O��D�O��`߂쉠��4lҮv��q���g�`8Y6�͇Sp�7��O�O����O Ā@��];v�
кE�c"�l�K1qƛ��'�r\�,"�H��'�?9�'~�� F�Ȳ�W�^<A�']5���3�x��'�H'�y��|��F�#�lS�~a,1su�	$f���0�i�剡
)>�a�4��S��(�������Z�
�ْ�O3l�0��)AқV�'Z"�C"��|�]>���q��I�"�O�
H d[(D�,�m�&�B4��4�?���?���Z{�'�b�L�M?Ҡ��LRP�m�ǌ�xC�7���W��<��џHӌ�"g�~i�0⎞W�¸s'�2�M����?��Q &8�1�x��'�2R�X٥�h5��0!,�z����c�i��'�ܭi��:�i�O6�d�Ot)H�4-���jЫ\V��S��A�ɾkidu9H<���?aJ>��%��A���LZ�32*�B&h�'_�P���';�	���I���'�2�dMYd��P����N�, k��9O.�Or��O|�Op�$�O�!@�JU:�XuJ�2b_�m���ŅVl�<Q���?YI~��N4b�K� ��\�R��운a�PdQ����ȟ�$����ȟh�"�c� Y EcJeJ�A�:Y��cѢʤ����O|���O$˓2?����$DQ�6�6\�M҄$�(��@^(��7M�O��O�d�O��Pd�O�'��0DUd���a=k�����4�?����
�ET�$>��I�?�0�l��"���p�ˀ�hd kF���ē�?1�K�f���S�����>[��Q�X*&�Õ'�M[(O*s�����0����$�|��'�(����CEa��J��UQH�d8ٴ�?A��i�<�����D-ʧ�h܉6�s+0e��J^Yl�� ��J�4�?9���?���<j�'�2㎗k�P����7B����lvB6�G�9�6�"|"��g��4E�r)��9gAӼE� ��ѵi�R�'�r��̼O����O��ɹ/0�i��T"�d��%�;S�b���e�(�	��������p���>7����"�P�e8B%��M��H���04�xR�'�b�|Zcni��2y�<�B�^g>���Ob顱��O4�$�O0ʓ/�<SF�ٔv�Nd�Vm��0@q��0w�'c��'"�'b��'k��1��en��x�'��.����b�L�a�'�B�'^�V�����'��TÒ3Q@ISr
ʑN!(�ZA%�����OL��7���ON��O4R���
3,��B���������a(�X�'f�ԁ�a� Dz�;R��1f�D��	Ot4�JT�N�,���yLԎh�Rԁe�?P�������~r���B����/ú5z&KŰJ=������.a�j �.^�q�<ܓ�+�5?٨��Ն�+`}N} ��Z'�*SS��i l�`�.(@��1,�+�X	8V��1T��AB�Q��h�"d�j�j��&��RX�Y�I$V�{�-�W�t�����np	�B�/_��H��Gٚ�?����?�Q�/j���!�_R�����F��]�a��^{r5�6#�{#�@ ����N:���Tl8.k7�H�Wiġghr�FR���uA �n֖�3e Ӳ{��I���˺kb���@��Ͽd�HZV�h�~�P���@q(����!\�&��<%?���^y����[p��Z�̽�ЉZC/M��y��V�;� Q��	+V�:���,��O`Gz�L�>�*>Bн{w�1`�x��@ç�?�)�\�r��?���?� a�N�O,��ѴB��+G�+I�h�5��%V���
a"[,F�T1
�gǟk':��؟ўt�� :is���t��x��C�k>J�psC3Olc�`�t���S��r��Li�eh���pdZ�L1��/ٌ�I�"�d�d�����I<���?!(O�ݓ�S)�4�$�јē6O���B4u���a�^88���b�&vlйDzR�O}�[��(�K��M1
X�.�5�f�E�E�ڵ����?Q���?��o�����?�O�e�%mU&'��Yc�� Y�lu�`"ʇk��P�@�����'_�A��*M�0�ҍ"!Ã4��!��jc�2]�� S��10�ip���jV.6���{BK	�?���J��;`NF,d��:3� ;v���s���%��s_\��蜛'�}��
2�̇��]�'��� n�0�%Apx�`����y�dӦ��<��ɇ����̖۟O�~��6���9m*�P�Î O�����nR��'\ۡG�����C���8##�O�����K�.6��-@�KS�9E�<��ј6ø,�I���,�y�+]
	7)p��O2���IpS*V�qu�T^��u���?x�=�'�.�����?��$+L�L<���/�=ľ9j4!���y��' ��#�B	е)����7�Ĵ;�h��'�*�XV��<p��e����Q�'=T�D�qӾ���Od�'�fE���?Y���.YG �+?���'ݘU ~�qύBm ��L��fp
1$�����/��O:u�2�U��%�X�{�I��0���6�P�vz,���'��P-�����'y�q�\�T�zu�.�&1�tA��^�I���wӎ�lZ���E���>��;����fC��{U�	 M0�̓�?)�IQ<pGd��L W�.ii��$�^�'4�$�'�2(�t/r ~��Ř�7����'�⃆+AN�'Xr�'.R�x�u�I՟�j�H�1EX�%k�E�����ͷ 曖m�(S�b�@����)�g�'��q�󈅸Q5��x ��4�t��qO���	MK
&/ZI����cX���Dی<SKM$�X��!�C8:�	[j ���ߦ�3ܴ��'��g�? j8sT6�v����N)�9�f"O&�p����\|\-�����)PaR��r�'�V���$+z��l��I0�e  沌�6�ߚPŨ-��̟���̟�	R+�џ����|"����@#��t���Z0"�Z*��ÇkI��z8t��19S�<��ɪm9�E�ԉM�s_@�)4bUfNZ�j�cF���q	 sB���9O~<��' 6핗^���K!N�-���xE�·
��dm�r��?Y�>�I0o��D#���%>Ѩ��ơ�C䉕?�Dгk��<Z��τ����;�M�������ep�nZ͟���W��LVDteZ��Z�}J��xE�9Cde���'���'���BV�	&����hԦmz<<�V��~�׍A��Z�a�aԸo���z@jb�'�L���L!����ٰG�48s�\?5��HU�`8�v �D	�s�*ʓ>��|�Iʟ8%?-�I�-h�);���7��@RAI�5v阐�	u�S��yR��L�m�3Dكw��e�u�����/��|���x��,d5f�s�A�8�4(�W�M��y"�ڹz�6�O��$�|����?9���?�ʈ-�B��Pn[�	ZU�'8�R����0:��A�m��}����0��
ۜ9ڈ��;u��I�1�V�P�)ՠ~!��S�L-%��8ipj��5�j��A�E��j�ϋA���}Z��D�u��3+F�	ʔXa�'VN��Iݟ������,AS6�ؚ:H�癑O����0)PA�x[�]ɱ�P�^��<��/	����ß�iEC
n6R���5&��=K���֟����@TqWl���Iҟ�I��u��'rBB��~�x��/G ��4{dd�M!���ӽ6���!Cj*w2V�H�O$�LY�JDƸbA&R�h^����X�K�N١��2g��K7`�gb���'c0,(C�^�Nk�,�ՠv��g"�7d����d��x)�sA`��,��o�O��oZ���?����\[�
�WO�59ƀ�Qfkq�!�d��4�r�z��@�eZX�D$X�h��Fz��O��S����ש�M���J�"h@t��	%-|�����?Y���?���~)�����?)�O`�p���Ŗ8{��6)��/�xO���1��]�Yz��џ)@�6Bk�	�'��N�����1�:����4qWe��HB'T�FR��3�?9��iB4ɋ�C?<����1hPw�ࠁb,s�x�ĸ<������)p|����;��4$�5OX!�d��������4�V��PI�@¦��vy��q��'�?�.�L�3��K�����)H���!d̼n�d�O��䝝+6p��DL[�|QbQ �)<%�"�&9 �E�e�@8uT��Q^�d�d�I�}�\��f�(=��bq�˽Q*N��gi.jx�j�z-@ȣ��E�\�R��	 �P�D�O$�?�
� ��+�敱b�')��2@s�����V�h���ᔆ-�X�����B��hO�)�z≸D�� #��)08��ZAɧoK8�	�kix�
�O����|a	�?Q��?!�#]�?��"&�o��d�"�Zz
��J�BV|@�E-���FU?	�|�� � !c$cط-ᴨ{�o� y�*��)�t2l��3�F�W�*���L�9���eX��rx2G��?�.g���G��AD�����Ӊb�y���O~�lZ��M�������jS.W�T�W"��Ύ�1����y��';�}BdP;!�����mW�d���@�<�O�DGz�ʅ;Ee�o�@pyҭ^�@0�0%� v"�'���ӥnF�Uz��'���'.�םݟ���'E�� ��BF|��9��H	��	� S�P
j���U�'/�IBТ#U3b4�îbWڝ�?H���S�Lx����I3g|xsMє���sE,�����j�z�d�OԓOt���O���E!�a�I��ꐻS�*dcd ;D����,xSTx���-E։��
��HOD�)�O,ʓ}Rܼ+��ix݀�L�Sn��p�c��ݑT�'�2�'+"ḾOy��'C�	ݜ&���u�܅iz��g,ΐj�k��jeH�󗆋#M�z��UN$"��=���d����*[<>����Z���;�Ś9w�e�ǀ�k�n՛�G+�hOq�v�'w>6ܠj`�S��1.���Hv��+�0n�o���>�	 !S5E2���F`^���e�C"O�UQ�*��O��u���B>4-�A�7;O\Xo�����<���i�	s� 푁nW��jMX+"�!�3JA�e"1'��5�`�a�,N2�!��Z� nv���G*[&�P�r��}�!���/9��	Tl_>��P��'��A�!��\��� ��B�Ki�F4j�'c�I�t��`*�	�ߖV:��'�Rq���:;�^�����V"���'�ba�hI8u�
�k���J�Z���'L���7�8�6�z&[�A� y(�'�܁��@�%')⠈6C�/I��(��� ���g��m(�����GyM�@R""O�����Ҥ� �xVJ���m˕"O�Y�d�|Ή��m���՘"O.�ӵǄ�<�J�# ��5>2\��"O��1�WMJΝP�[�P2¤D"O���u���5|�]��h?�aأ"O����а'�2)PDk	*<�В"Oj$22�N��@U�t�M�Jب��"Oޔ�D�ŋ�Ay���>�Pxi�"O����%L� A9;g�p��"O@I@􄆚4j�̘��@�gG¼�F"O8��2�Q�(T���9h@r1"O|D�2i�&Dȥ���W�Q�L��"O������J� ��d��r�n@ʆ"Ox�P��3QX ) �h�6~�td��"O�2d�K*H���'F��⽊�"O�%�W�,��-����$��2"O�t3u�L�?,� 5��0~�d�0"O���f��c,ق��պW�BѢ�"O� !���0OYZ�B�S0,�`�"O�HRV�����l�ĸU� "OPM�
�d���g�ۋLE�8�����<g<<��&4��);�ǈ�W�4�TU��`��%a��Y��:P!Be���AtBiA��NTD����9ږ�Gx�.U�IxZDq��
�'p��C��1
jR���U4G��y/IT����2O�Y�<s��TĹ�*�'���w0y�FU�{*"A�u�] :�����x~��HR�s2�Uh��=�������$8#�Me?�� <�禁���UD���+��� X�ڼ�6-X3�a{#C�Q�i�)��Bz0����	����E?��ɴ��;�ܚ��n�mP�띿��dڋB� �ٟ��avk0)t�ҷY#uW�E�7��q~|��>9n�?_��ы#B�:$T\��Ǭ3�F��K�Ih�k��|�ᄥF
"����@πdyR��Z���)�oݺk�c�(E$|� ��N�jG�\J
���P���?n$h�rL܅ 0��$5zЊ!��B�vn�(P	�Q������"��VFT�p�7N����o�i�8]caL�*A����o���&�	\lĆQ KA0�.z-Ҝ���ΐ ���@�!���?�'P�%��@>�����,P�h�>�+�K"�HO�.�v������I�Q$|8Sʗ$��)x���d�Q#t%]�"��L�#͐�G�0iTi%bR�(d�D����O�e> �'L��d��=he�:w3~9��>���Qkи��Ù� ����ML�=-������}wY� �!"Bk�3�(+6����4%i��I��1��9IҔ�DEV�(�	y��z�ǘ>��*����r{$����H�7����'��������\���4��O�l ��#J�k Q�r�
�b�4 T"c�I �� (V�B��<����g-m�@9U�p1]*�g�%3�Ӣ�s�~7-V�k�t�cK?���{B�
':�~(�����8��1bE�q��q�w��~)�����xV�3fU�1�q�q���4��W��?zF��mӈ%GȈ;��[}���e��y�'f�p�0j�1rb���G�s��Y�Ɩh*!#�"�>�c'�G���BW	VA�	Ы`�l�Z�ަ~��  �.���M�Ȝ�~�X��M��1Բ�X���N�'�tE`Fc�2g�-*�Q�Fj�<�o7���Ӕ�E�Ju>����/z�pѥ ��?�V㋬}~���c�y��i�3J=pbn��f%�T����V�F�� ,¬�ФԲ*� Q���Z��rZc�Y� $�2�$��q"L�E䓥)B� �:O 6mK�i����' ��''�0NJ-1+A�.�t8�*X�0�Q��)�G�J,3#Q�nt9��'
pѐ�KO�Xu�\A↕�Uy�T � �t��W���X)Z��:��|�DDz�2�h�+Z4k�>��ʏZ��Y�S���0��2k�j �b�����j�(����'?"L9�pyX�Zq� =bS�4�'���`��.Ѵ`(Q��ՎU�
��'���Á�3X��h�ܛ4-�Ŏ.{��=��(��FQ�6͊�%4���?�S�	gƐ�K����][D�U�7<N�sf��4���۵MD1e<qE~���t�I�v���� f��0��h�����hO1�K<q�]���g� ����j�"g�pFzZw:2@�QǄ!@�� "^���vL��B�9�FˤH����+ �O|.����Ŵp�w#��,�~ ��#¬U��'!�d��H>^�f\�6�O�',t�/�;N��	
��8c�Sn�'�:ŉ�Ȟ�t�R�A����!���+Ob���Cm�K(y�tE "��?��HM������}i��"��D}B�ǌ4p�I��l'$�Fy����؈��Y�$���h�I�%�P�z�,?}�f�h�'",�&�LcF-6p44	ҫW�6D)��&�ЀFy�'m�p506E+����$��)�9��#��5!u.��#�:�I�K��#<�'qT��b�81y�1�'eW+X�������i;Z��󤔰x��ɲ�i��|}��� <فu`�\�t�!�R�|��R�Ã}�'Jx��C[�Т�	_��W_���P#�$��Y����L� ��O�b�KBPz��h���ㅛ�F�9�Ձg]��'�i�q5�X'3:�c��y�<Ey���5vϓ5Agl���<H>ehb(ǹ��ɽ9���<��G≖x�j��G#׭m$>��Q�LV7Nh�#�F}���C+Ǎ-�>��U�\/�Ni�����uP���R\|�@����;w�b��!��>��|��OJ�#a��AgH�h*���g��U�0^�D�HC�.@$=����1
�Ѣ���O��(�4�J8P�������G8��u�d�<$�(�D�Z.t�E�'Ը�1�ůON��1 H���,�B�K?3��2�ɻ7u��ڥ�Y�䖑 ����d�O"��&Dٌ����O�޼���N^*��Ri��t�(]0�k�R�<y��Q�?v2��'˅V�(h↬��G�D����O�2��/ۥ!(i�*O���կ�!4�$U��I* �Yp�'�.L���"b*����'V�����F�-G�ʓ2Xx���K:=6�X�{�r���瘤Q�,��t2z�8�F��#Fx����\H���Z�$��O��f��9+���O��c�p�e��9џ�;+���5�W�V�Z��L1D�,Yg�H�Z#D�j�#P9��
-޲5f���	��y��Q�_$����S�D�x���� �y���cڀX�3♜4y&�P[��Oh�̒���'*�x���F�b����⮓|-t�
���tP���<��怽e��"b.��>A�"�KP}� 13����I�z��(C,�C��vEU�z�c�\S�Ⓘ.�џTP��V��T���;&����:D�(�$� ��-ڳ*���ӧP9WJ<���'e\��u���GM��7��Uҁ)�I�<B�ɯJ��*�����z���l�=�$"?Is�D�-Ť⟐J�@P6g���aJ/$촹p��5lOL�������$U�������J�>���nG�F��	�'�R��d�'RY*v�З\���Z�k�lR�}��J�hTiF��D ?g�Yq�Gb������ ��?���T [�zS��+F�`J	��Z�1	�'�!�eh�s�!Q5�ӚILص�d)2�HO���$c~�QA�b҇u��0W���lɧLR8�5�tS����	�>�-Ɓ��cktё�*O�n(�yՈ�?�������uA5`ߋL������9'Ƞ"`�	 y`��c�W'���8�D!S� �� �?K<�	�Ү,��!U)-kJ��BӵM��A�$��B���б� �XhGC/N(}P�˵>i�R;x��ysFᓊ.\�<���]G$�P���z=2=J%@�0<��))��>y�B0���O��	� �4�� �����.p�ʱ.�����<��X?������E�p�ȵ&�O�Y�Wn��8�s4����>����dS�Of��<fM��)�D@�(AP8H��M�|q"�h��� ���Q�|�b�ɗ�W]L�P&(C���$O�H����FP�+���y����<J�@�3b�a�'�Fם��*��%t7p�S�]������$j�d��G*͚v�,��.�+/xXM�bC�J}�aq���L����F�!,0���y�p�!n|�"ъ7�%F�z�s%G .~�����O3"���w�B�2-�VXV���.�Y��(��Dy�'�ē)��Շ
y�I[�ء8n�����(O�ԏ =��hY�ȁx���Pe�!P3�?Rn`���K_�@�>�S�PP���dR�r{Uj��RNjq��=�.�P�b�>qV���pX�����:W*��t[�@q�o�E?��x���a���<�tHؓ��j�fx���dvݩ�����.���%i_6��I�@�4��2&�g�\�Xq�[��t0@�[�����*���9,Y>yN���N�>���߁ I���t�U�6��<�S� ,��)U�M�$n�+�c�:@�X@�f"O8�p�+����9A��	.��9�w��)w>�<���_n�8C��[M��?��b7$Z�uX�x�cF�1� ��	�@�~��qV�H���c2O�I�Eo�2��$®	H=�#��]J��opӆb���R�#���p3��9p���PI��*t�>�޴�uwL�S�F�@3�^�*�9�vM�G*&��h+�YM&�L��jǔq�p�`�4-���?����'�e��c˳q����$��/���ChY���=�[^�2����	>Kk��-5�rX8R�%!	Ra�gǲ����Dy�'�ēS����T�
����{��9@PZ��u+Ɖ~����-0w��w�'L���+q��p&�M$v3�� �}��,�O��I&\�(��Y�.��Ƅ�\�p��/�}ra v�����̦8�[��L�'�N�x�m�Ok�9;b�ݫ,#�8����='J��2͚�uc����E���� �qb�&�-w�,=;�_�cQ�Q�tkv�R�p��"ⓧ�'R�U��됿r3���p���6(^%H޴j�t�Sf�^����ՋDI��<��SуIl����6��DB���3��F���'��O��8Ѯ4XE���f���s&P#�ثSmZ�<�Š��b���B�&Q!��O�d�� �j�
�Mď�%M	)�'��.ؔ��R,K.8�H����n
�L" X
2���2�OuQm1FER��g��!��|���Ʊsk���qC֑{�l�:���Z����F�șu�B��%��6~X�R�lR�֖D6�hDΕ>q�L��/�UllK`o�'�O�@�2�݀:J,ô�\DF��U�i�&�TO�%v5���؈w;
QGy�'�5Vf��P-�4�U��, 9�q�K��'
�O�b�y���-p�	�r�{\���L�w���Dy�'0i�v�/;�\���\П�ԃH9*:�Ԃ`JY�#������;�	==�"<ͧ'_� �El�<Lު��Eǔ +�ib��
ia�6]ӂ���i��C���� ��*A�c��	Ӆ b�륤E}z��p
��r�0\�>� ��к&�Z��Zcԯ(L'���,
�3��(
���l"Π����s(���d�M�mL&�#.O����<<%����W��W���@������C*�n=r��.|OP%�Q��p@�Z �f~��ӐEby�c�$X�O1���T&�<$�[`!N"J���"�8�=��AT	2^Z�c�\�[�����$U�n�`}C���N�(q��N"�ʓp]����^u�=��eyVɓ;�j,��M�'x�0�@����!ʓ�I=d���a��6�"�ɏ4�l�!�E�
�UI�fCLy���6IT:)bS-���#���;t8l�ęw��?������mC��J�9N!��kб1hxA���ԟ�O0}�⏇"X~VS��]s-L�1
�n~x)��o�����$���$5ps��J%���S
�g�IY�'8�T(��~�S��ߵ���ϸY" mB�e�=����a�<9ć� 7�$Ct��R���Z� Z�<�dB�p�T 2ע8�@�ͅ}�<��dØ�N� &j"g︼Re�{�<i��I.�v��`���Q �@3E�r�<Q��U�&**��I�
`�Ν0c��c�<a��-;�Q@��	m"Z Ȇ��b�<	$�28�n���g]�)�$���D�<�Ge�mL:�0B��.,m���\�<!��D.�n`�4J��To&��֋�V�<�de�-s�
ɐW�\✘
�-�U�<��\�- jx;�f�0+Ұ����Z�<Yt핉h�ЙI��5t��ۑQX�<)t
�I�T��ɱV�<٣�*VP�<a��Ց�K�(�H�!���C�<)s.K� h##M+� x�c�Ei�<��43�f���js�	���b�<�1dS?p1vT��A�9+^D�T�b�<95��r��q��Ś!Bx����I�<����#k�~y
#��0
����m�<a'�JI�PR_YO�xB�H0�!��=t-*=a�  P����o�D]!��D�6�����
�.b���O]uX!��Tt݀!��\�@� �ܺ4q!�ę�kb�yA�NIPF�he!�$�701��vO�4O*da�weU4	?!�d�#dFz�+�Ï�5�F��A��j$!��N�cK���h �C��$�҃�!�}��p�刄-j�6Р���2a�!�$m�b��Ԅٍm�Bħ�G�!�$�	O�l��$п_��Pk�67w!�d�y�P`��46���(�ʜeq!��=y�T��ʋ��:V/��?!�$Y�)�D��������&:G!�dx^ܵ�P�B  {�Pt�I.!�dT�n��)su�P<��^r�$��'m��`a�_M%���a�B J<Mc�'h�<겋Z2'�j1�"�"@
 � �'�����!l*���&�#"�T��5�>�Rp�ȉJ.@d�����Ն�S�? Z��7�Q�vG ��a*"tJ1�"OԼbdC�nj�a���?j>��07"Or���!�5��\���8�eYF"O�Րa"��<�@��K(t7���"O������ ]H�C�--
*(j`"O���pQ8%�+�&�|z#"O�m��I�%���K`*��Y�@�3`"O��I�N0U/TuqRc &�ZDH�"O�DZ_��QҮE%C�L�pnD�a�!��׭R8l9*��O�3���f���!�$��^{�e�u��>S���Ó��$5�!�$�)���sa��q�`ء��3&!���mХb�4#�4U�e���#!��^?o� ��7Z"�(��"!�Ҡ59�x"�Bū@�0�FFԄ�!�D��s*-A!�R�*�������!��	;93���6Ĉ3K�N��f��p!�$̬Pi�sߊ6l� �"��9Tn!�$�11RV�be��m	it(M�6!�D[�'z\q��ǆm!"i�2�W=W!򤆎r�q�ٽxw�<���d�!��:����o�qg&혤�C6�!�D�j��c��\�@�����P�!�$\�C�j�0�E�S������%!�$�:2���@O�>�B���	+k�!�@�kM��W�V�B��a���!���'0�tm�����H�Z���͓2#!�D\�&nF�j$ȉ#�.�AEᕖR!򄃫	w���I��b�
�b�j$N�!���$�&�1smY�{�$��Jt�B�ɦZҌ�iW��2%� qp�D���0C�ɩ}F��ѱ�[$URP��P�ܫQ�B�	@A�XѦ��/}R���+��B�I+g���9l�#5غ���śR�rB䉍<s�� �\<tR����+��|�B�� W-��x�ȗ5@$d�Z���	T
B䉀*)��"&W;(��T�=�(C��%]��E�VȞe�$h��g����a�\�K�QF�8��
�'tE�G�+D�s�)���^��	L�KZ��I�5D�� 5G�)� Ȗ��>v}`0��'�J%��k�>��x��)��m!�'2��9ej�0���w��/�"��'O��:�,�2I�i���� >�(+O����\cBp!˖K��b:$a�g`�|�!���.2�I$D֦m"I��芪��pF��N͵Oyp)ؤ �)jb@����yRHE(}����J&FEXș�U�y�O�S:j$�Ė*q~ʜ�@�Q*���hOq�` ��)X�Tz*��E-���ݪ0"O�����H ^��Ɍ���H��"ONap�L�0/�0k0	\K(�8"O��S���-VP��$h	��"O�, pE {�N�J�5���
�"OXP����v���R܊{%"O,@����&�Jt�@�>�M����@�<���V<,��hκG�Lc�}�<cI�<��H���?o�v��0��v�<f!-ʩ�D̹|A���qIo�<�0d'R�$�!�:u��@
�fEf�<yw���4��I��׵V��<z�Țc�<Q�
9ur2��3M�(��I�]�<Q�g�$,޼*$X2�$t�׏ZZ�<�E
��>�3�V-\�P,IW�<� �,��'!~��]S+��%8͙c"O������8���p�#X%S"O
��T� PR�e�4��I��"OJU��e֫X�r �P��3j��D��"O�II��A*t߂d#�nH@�"OV,���*r�d��#�C�9�ݐ"O�PQ��D
�(��p띖(�`�"OXA��T��H���Y3\�Fղ#"O�C�퀆Il�6�ݺ\2HXhs"O���c�H7PI R��	�Bi�s�'���"(�$�0t�cN6w��=�N?D����DR8�4�8#�˖4Dz��((D����a�
�0�B�
D>�
Q9D�|�o���$ƌF�䚓+��4�!�������cA�78���9�!�2%%�e����,)� u�đ,�!�S9#1ڭ�G�&j^��G�-�!��@���-\1N@�H�ʍ
�!�T�-p�����q�$|� g�'�!��2�R�+4)L97� /	 Oe!�d��[��]"1��/" e��]!�)x*�:t��|`�h�5�Ȓ2�!�[�@?6�����c�������!��#?d�s �K_�l�ӂl��=�!���83&�@K���&���#a&��nG!�D,t<�C���L��u�־/\�	8��>iF�ՠd�H�+�Gн"������T�<��W��P���5+�d�D�\�<��@�$t��X� �<�%7��D{���i��h�#k�.>����W�ѱ�����'�8�4,Q�-��9$j�2lڈ�q�'�t�8��+�.L��nٚX�>��'I�\��R81Ox�!s�\�X��iI�'LH�X��@3��̉�OB�q��'0m�tm��CߴUYR暣w���'�ZS�(��T�R".ݦq�V�y�'���� ^1&������gI~�0�'� K���?�zpJ�BR=-�m��'HH퐣�W )mr	!S�?U�
4#�'"�B���0��\8�Hfz�Z
�'�Pp�/�"��l�L�L�E�	�'h�lR6h��+7���Q�� (A����'��!UH�!(�e��J�wd��Y���#O��"q�H��@̒0��'J�rɘb"O<M��m�0)D.*��ω<���J�"O~��r �.o��(I#"� 7�`��"OȽ{���}�
u�d�P� b"ONE��K׶\��� I�\���q���D���IHxz,�A2�������S��r!!򄙠Q���Ib�K~�������!�Y/3�D����5���y� �!�����	�Q�ӄJ�XT�C�F2{�!�dT�|g�QBG����%0��(y�!�X�:�J)�QE�}���:C�+�!򄌠
����#�&{��
T�I=?g!�E�W%@`֊<��h҆@H�EO!�d4Q����L��3�ʑ
�nZ�/;!�$��i]���FF�3�L�(P�5!��0�j�ڗ�Ȃ���a��ւ"O�	(ḯu0�����07`�4"O�]8���.k.0��j�U��K�"OR T��2.V�Uhӏ�"S�(%@a"O�=��HpP�d��(�p%�Q"O4|�B+B� ��z��z�8H��"O� ����M�3n\6d�� 	�:I%"O�ɒ��U�4	(���Q:l����@�Oȣ=E��͎5z!�@���@L�0	�͛�y2���\���Ǆ�?*��C�N��yR�ǐ*����ff��8�4e�"N�y�&��[�=�K�;dB\����y��e;�q�(;9V�Æ�yb�Ҷ	�"���AP kR��\�<�#��0�$Q����~>jS�+D�l�A�4�zanD g�`x��QW��x�'��a�v�$qD��vj�;2�4K
�'	��˖$/DTdM�G�9w�4uۉ{�)�)�=y\`H�EΡp�堤�l!��qu�p$�24��a!�H�'8�IN���8a�1Cx���1!Ѕxg���N D�4ÐIE� f�d��J��Q0̌�Ek+D�D���_�(TRL��%M���c��&D�XpQ��(7{�t1���:�`����'D�4S$D�m�@T�@[2"^8�b�!D�d�3�7f���1A��0*�;�a5D��3���J��z�샵X(1���2D��@˗A���ʤ�e�J�x&-1D��ȣ.��Y#��GoE���!�+�1�O���s�H��[D��j:<��"O�Y٥�ݰ�Š�$L+pށ�%"O^�3v�0i0i �b�����"O�̓�`��,���0%!�%|O�ѓ"OL���E��9(�`�y�|��6"OR][�!A��<���n�=]���d"O��P�aջ}��!�O��a~��!�"Ot͂笖
>:���#t|p�4"O~����92�A;Q�{d�I1q"O*�����G L+�ŞN��H�"O�Ey��Ίc���A}aҏT/WC!�$�9<�kDG�.P DKn	�2a!�d��iN�I�b��8�D`3��O�!��C/s���b���l�������5NA!�dR"$���HfE�E��M���(a!��G��P���I+m�D	���, !��k\%[��C9n�Dڀ�V�JO!��W9	�6h�a�9t�����BO!�����ўzrjpR�b��ȓ u�)��)��_��9T�30G)��K��|{���Z��0�/',�фȓb�������(��W`Q%$i�4��LRpp(���v�ȩuL�}<y����؀!A�Ę��[�C����ȓZ����kQ=2���X3�Qu�X��ȓEsx�Z�. 8;���J$�ըqe,��ȓm� kU�M�~W�D P�&��Y��Y���'Ζ��P�I�:9F9��H%� �F��\�)HEj�8H9�ȓ9R�Y�f�,<���t_�x�dԆȓx�pqr#�)H
��%�B+\1��ȓ62�ݓ�k�70r�uaƂ�,q_r��ȓm�-�$&d�Fa	����C�I�(�yH䯂4z���!�Gɇq��C�	[����aBҴSZV΁&吝��'�\X��\�v%����Q�:$K�'
P�qiE�o qp��*y_�ٹ	�'�R�d�-Z��E˒G�P�	�'�~���A�6=�UUH��'(J0A	�'S���(ߤ!��h��*B	K�0:	�'̎9���)vޜɩc`P/G�|8�	��� ��×⛕PU�����T�B���"O�Y�ŕ)4��TIQDƵ�z���"Oj�
��,Hڔ񨷈��Ł�"O*�b���J��(�ӨE��m�2"O���M�&: � Tij��kR"O&�i��)Q}:�s�[2+�u+%"O����\?h�(Av�Yts�5{�"ÒC�K�.�^���A�Ps �XD"O�ٱVJ�b�naq@g@"tS��b"OJ�:'�"Lv
�P�ȢcfԈ1�"O���B�r��\���)� 8�P"O
 ��M�c=`�"�aդO����a"O"� �d��2��)g��4�FM��"Ob�K�DH�o�|��`��r�"O�]��P#8���2Y��"O��y��pA�-����p�Z��q"O�E��FN�r�V$q����1"O�(�"�N�:`ѷ⅌q��(�"OtI�U����3ThE&3��lr�"O@��"jQ'p�4�f�ܚ	�D �b"OD%�J��<[b0ת
��dek�"OP�Q�,�vFR�@Ĥ���h�T"O�����!: �-mTjW"O�e("��84/�,R'Iā*��e"Ov���R� �U��J]��"O�U:v��>ϸ.�ȴpc�WR�!�/M%D`�4��:L�r@� eN��!��2Wa]1��g�\0q��ҬG�!��]�o�r��'*ИK���OU5}p!�$��"�� �]EnXxӮM-e^!��P"8L`�@�!�!/N�b��lv!��D ���@- )蠀TI]0+I!�d��B~����^#o1�}��.�n*!�݀h���um��a���S�a"!�D� y���-� �|�pŬV�R!�Ă��Vl��+��+@�Cv%d!�ǹw�����?=��$J�Q�!�Ć�]�0T֯7��a���n�!��V�9�:)�7�×V��=�,��3R!���b�
q�e�²R��|�7�#[I!��
�D#�\��@���<���ט45!򤂤{.D5��(��l˔ȻD�I�K!�U&����U�|�$��DD-<�!��Fy��q�j�9����AM��!��C-D�2�IA_{ؼ��ʓ6G�!�D�	(ph�A�$^��2J^�!�$R�J����W����`o!^d!�0A�d؊w�^/ؠ�YQ���C�I�}Z��#rEۍb\J<hC����8C�ɟU����S�g�T��-º0�B�I
@��Ģeӧ@�аѧ���
�B䉫h�p�5��=@�k�O�yK�C�	s�sANQ$rH�Q�A�s!�C�	/!�B�;+C7�n��
¿�C�	�Vܚ0��oۃ?wD<*�D�6�zC�I�h{�@����K�t=h�O2~>�C�ɰp�|�a��H11��Q��&�	b�`C�Il�T�d�J-5劣Xq��1V�LC�I#ZN}#���4]�RI�2"^sxC��Q��Ht���i*��U+�%qw�B�	9H��teߚ	�̅K���)~�B�@�@:�"@�r��aX#D�B䉜c���k�:�<�7�V�E|B�	�b�$#��\\�p%���LbB�)� �I��҂.�n����
�4��8�"O�U�oD2:M�	� �Ľ�u"Or�:nI�	[Ef�?UT��r"O��1�!�fL�B����S���7"O|9GD-c<�(�'�w(%X�"Ox� B(�3
�|)RE? �r�"OZP��*L�$i`e`�胓$�|ɧ"O4 �K0)��ɇA *�r� E"O�|�FR�GK�:$��癧�y�!R���0f�88��lğ�yBē���8Z��&����)�*�yBm�9@��@������˱���y��
0
l�l�2��u���B�̔0�y�aB�T�����ΰ��0b�'L��y��>��鋴c��
�Vt��N��y�D�I�'�s���@L��y��F"DF�b�\*���E��y����D��uk� DZE"0OQ��y"����e��	�o:�)��.S��y� W��ܣ�JŪ^�-�����y�+��%D��B�כc���iVa+�y2'�C�6��i ��HH�%��y&�(F�8PV��;��{U�Z�y�	o���[�b�B���Iܚ�y�dZx��ł��0!����y�_�SD� �g�xӖ-zB��)�yf�p�~Ĩ&��Ȗ�X�،�ȓ1 >�bo=y�P���eō:@���?����"I�9�,�K��T�1��ԄȓO⾨�r��	����h�u@V̄ȓ:e��� �Kz&Q����v���ȓV�(���
:Ɍ�� �
�M�ȓwZ�PZ����b���Q�A?f9 ݇�$v���D��)��tQM $�@��ȓT=��Ʉ(s�\��ED�7uV�ȓ[�<��䌶��ݺ7k_� �8�ȓ"����%�(#~��dD�J��ȓ6Q��%�� ��!��_�I����e�G�0�z�0"bC�q��Ą��~E���17l�dȓ�S�@��ȓ�8�3��܄v�أ�cP.6����ȓjP!�Cm��S�r$��eЭVZvI�ȓ�4�i�F�%�^�rW����P�ȓj56@����9�3�׿'�Ň�sM2�:�����������G�d��oM�8#΄�F]9�ʇ7$6�I�ȓWbB��Dᔛsy ��d�ּ.�nX�ȓ8���4�)����!�u+.��$,a*���MfT���۝�B%��CRz\����]%Z�h�&��R@�ȓ&L�l25	�����H6�Q��Ȅ�Rh:�"J3K��mΊb٠U�ȓJ�L	9@�
���`ݑ9S*	�ȓ?.���`�D���Ƌ[�؇ȓ&�&�ॉ��-��|�Q`F	w� ���L��6)�����b#�&�N��ȓ3�R�[�Z�S
���0�ڍn��S���K��"�lݨ���"���ȓ���#���2h�38�Ё��>��:@�-y�b���f��nd�Շ�e:2�:�i�J�t,Q�I�I=ڼ��i��I��H�)b6nU�Po��"Z���0	V%#B�HI�<�#DC�u^�<�ȓ0͑S�M�(�Ԝ#6��V�����S�? D�Ʉ�vY�8c�lz>�(��"O���
Ҩ����>j��x�"O>̨��?)�!ޙ\ �g"OvQXW��/|O*��!C��� h#�"OA��%ߺ�p��	F=B^���"Oaq����##h��M*�5��"OF�FG��B�NX��lO�!�iQ"OQ��[���;�)�}
�As�"O,�P�+�;uZ��K�H�B��bB"Ofe���?x���!�է �(Mk�"O��f�5@�����m���B�"O���a`Sy�I��L�^���"OJ��f�t�\z����XB4"O�ѓ"�|ɰ!��0k��y�"Obm�RŅ�|4��y���$�D�kG"O*���ާ`�T�q�F&�~hط"Ov�;�n-<@A �]�g���"O,����QH"U���\<ĨIw"O�,��C�E�d���kΒ<#bmy�"Oё0j�==f��٣!�>B.�{�"O� �f͗�xb1o P��-U"Oj��*� {�x�"�ͨ�h=T"O<Mc���x�Hᣗ��p~""�"OL]Qw��{��Y궄�:ZKN@�A"O�����KX>�#��=/�p"O,�B���%O �x��ʠa{��!"O�z�n�x����g�� �"O�	�&(�5���@�-�|��"O�0q��7\� �� QX�=!b"O8�&T�rϔ�AtMQ�__>H3�"O6<�mE�~�p�P�Il��`�"O���D�J��hQB�O��n�P"OxM�Ff�3��#X
R�� "O����#�'i��Ƭ�=MtE�"OZ���/�gQDY��ryk�	P�<���۫L�6!�mS�K6T����N�<�4��7tX
}{QhI�OB��KJ��<9�+P���I���K�:t��E�y�<��F�/.�s&/����|�o�}�<ɓ��4 x��J�m�'�ᩄj�A�<�.� H~��bS�E�	�d}q���~�<Y�hm��h�����͒a	�Q�<)���B���Bh�lC0:���f�<�$��y�e��&SpԵy�Af�<�ؽ0��H�5'U�v60�A(A`�<Q�'!>Iy��V�1�.qI� �[�<���ޒ��D���a���B䉸6�Uyg�#!� �Y4ĈDv\C�I���h:�k�j����A��.|�B�	z�*�d�D�(������	 w�B�	Y6 �Κ�a�l��g��t�C䉧hp�����%xp9W�7P��B�ɗNVr��g�r��⦞)�B�ɻ�NE��#�f����d�Q�gVB䉗B�"T�	A�r[����B�	�M����Uh�0`��(0C�G$~BB�ɢb�j��h5+V��:U`E=Q��B�	5��e`3+D:^;�p2W��5c�C�	$}���P�lʃ �l��!A��C�I2tT���E��B��2&�bB�	(A�����'r*�8�m��"lC��($���{P�M4�d����\�xXC�I�+�F4�p-W�v0� ��ծ-�6B�ɴl^��kw,��`�$�˒0WdB�)� x���e>[�����dA�#gށp "O���dfӔC��!��B�v^���"Of�Ge��KY�6kB$Pp
E	"Oa	��,y
A2��SS�$*R"O�4��	8[�\Y��iГG�Y�@"O�)[3�\)&Ej��Q�>���"O�YuΊ�^- 䡃�
`�8�q"O�]�A�� L��,9����/R|�1�"O���-[�'urL���ɂq�y�T"O(��V�ɒ0��5R�\�V9��e"OΑ�!� �Ѝ�+t�nEQ�"O��2(P%_�D�Iq.J�#��t8�"OTa&H�B��0����x���V"OBD���JN�`����e�N���"O:eY�CY�Z�t���Ut =�5"O�])pG]
Gs�z�F�#UU2�(�"O��!�	(m]|�(e�K%T7�š0"O��s�$��%h��Z�.�g�A��"O=���͔m�Zq�
4�h�BP"O^M�R�
2��`f圛�:M�"O� ��\<4��#���I�L�C"O�L���ڋ~l%�2��.s8 aZ�"O�$r�����^�*c�ɬP��1b"OV=�D낂c2(t�B��V7���v"O���6Ɣ�Wc^�� g�xͪ���"O�H�ƚZ�0���5��A9t"O��q��J�-� �%i�,��"O<h�c$ٞ�$Jb�C�hces "Ot�䎙K̔Y
A�Z',.n�E"O��'�vp��R��3y8���a"O�)�BМr"���_�^�DD��"O&xIG��2U�O��4#H�a"O�E��	%oӐ���/��^�X3�"O�5��n�@ἩCSDAJ��Qx�"OX�[�U��� �8��ݒ�"Oxl��[�;�̤Z��A�N��a�"O��`����Y��>*ͨ��R"Ox�CPÅ/@7$a�DCҬ]_����"O��;�ؽfJ`Dp��K�QO�k�"O�!�ef��W� i�t$Ǡh?�l0d"O޼[R�1,���#A��JU)"O�mH��&��:����<v���E"O��E�m�j��l�.ph�"Ot�{�
�*9X��E-\P��a�"O
�2� W��Ps�#�<5@&3t"O�la�I�8�ʭ�3#��P�"O�)�3NĦqA�\sԦ�j�8P�"O�q34�HC1�u� &�,zx��`"O ��F���@�R�ԏw�����IZ>M���*�E �I�R�F,h��+D���l*:+���2�^�&sD<��(D� �a-�n��!�F�	�+RP��%D���'[���	ug�5vA6x���%D�(�b�9��҄X�
�(lɄ-$D��[�N�&�p��@�b�(`׮&D���Gf�*N=���a ��Zi2��&D�tY�N ��0A� 	BkPS�%#D�؉FƔ�s��pn��4?�b�"D��1`kE�}N0�ᆅ��=<�qHU�?D�x��苮{���fz""�>D����.¬9�����D,V&@�h5�)D��\h0�<bC�/[g q��g+D���A�˅mXv=��߱^J`I��-D�P����7^��eY�.^*4�Z�j!@-D�� ����ə�.ƴI�5Ⱥ
:��a"O$0h�L�>���c��=n �Y�'"O��p �1ri�\Z1�O�*t,��"O�k�JJ�?�<�h!H�+��kg"OJ�;AB	��Ѕi�8q�:� �"O����4rb2H����	;� w"O���ec��Z�+$�/�*�"O �O�/�ԁV��ޮ�%"OdB�k��hH�a�ѥ�M��X�E"O��h�17]Bm�ׅA0q�X�p�"OJ�+���/��)d$����A�q"O�$ ���\t\ 3��/��HS�"O*����[
�,��㍉f�����"O�l�ǐ1%��{6e�&0��"OAOр#�b0P�)
�q��"O�B5��{�Ȥ��*��^��d
Q"O(ͩ硍L���d�������"OVqZ����8�(��&��Y���!"O��Ӗ��{�̹�gkˠV���"O�� b�θ7kn�����;��h&"O������E�Dի`�̈́.�0y��"O�e�U��'p�0��+BҐ�g"OJI�͕�/���ru_�S�(�p"O4�1r�� ��Z�#�4W�""O�q�c@6X��8i��$��@ɷ"O�e)ѭ|1R9h��\���Ȅ"OZH2���Z*��� � �a"Oxܫ�mN�v&��xbOR;>�<p�"OZ)PW��
�P$B�,.l�Q�"OHXAn�?���!ҋJ��%"O��s�R�.��M�*��>y�3"O:��m7�P��g)�I�v��"O��/�
&(��"��(c�m8'"O<z4�9cWx��&'٥7����r"O�	��M�2̘	�,>�2��"O$AM�+� ��A�]}X0�"ON���杤[Z�w� �gz6�u"O�a�`��>m�<@��rQ:�I"O��PUdG�;��5��س@��م"OD�0��1SEbj�	q�2	K�"On��A\�UlN�����g4,�"O�(�4�@�T���%��!rA0�"OV��hI�|�b4Ӄ;�옛�"O�����6< �����/�@��"O(��t� /���b��!+�X��"O2t��+x�%:Z` \��"O"8c�$n��ara]�#\	y"OK��b
����hJ æ��Rbď�ybE��m�\!�3"@7�ހ끨"�y�+�1̢PCc�,g���p%�y���\Ov�B"�ߊ�壤ƕ�y��K`�L��T����W�Ť�yB�W��L����}���p�m��y��J`V}R�B�tת�i� ν�yR'E	{���Y�	$[�N�8�y�L��[���Z�z.�u	��yRK�f{�Y�P�ä(ZJ88��y%Ә+T� 3*�J�2r���y���-{�$e�fψ��R���J��y��fe\ �T���h����y��=D$aT���<�M32�>�y¦R�Z�� ��R4�0�a�Σ�yB�e:؂�t ��;@����y�Hp���$�+�>1�H�6�y
� �tz�i�y(T��@آS�fT
$"O~=Y�#���b���4�����"O2Q+�G}ve�� n��H �Rz�<9�P*4n�l#�'?Dw8�"j�l�<��A��s�.3�'k�"�	@�<)�
�>*Ƽ]�1Ɛ�5�6�x�<�qEΰ6"��3��Y3$�"-T�z��$s��A'"�d4 W/��C�ɽPr�ܳBb�L ��SB
W��C�I!e)�e���d (��!AB�ɵ`*���ES=Ӹ�t�[&i��C�	3Րd*��~q�����7�C��<T%�81ЃU�����`�=��B��)}�Ecgiƅ*�RI��!*-��B�	�+]���D N�x5|��냽(��B�ɏ��[F)γ���aC�/%#B䉋;�I(��Vu�р�G=7S�C��'J|8�"Ͼ4;���� �B��B�Ʉ@g�=�E�� P:Fir�͝y C�	�=����Df$-)3�]^h�B��Y�|�j�H'g,���j�C�ɐ.�6\B������z'ES9n�B�ɫ(���tC��$���Z�a��B��9c�2���	\�o��yPg�1d�B�ɽF���
�p��9�.͕tdB��o��HS��X������hY^B䉽qjV�b� @� �1�6�L,3�PB��u�z�ʁ�bk�(�J�(XBB�ɛwWt4��"+S�D9�MU�zdDC�	�d'�,����s�T��l�0C�	t�V<��JFg��[s�{ۦC�IW�f��G
�y���R18�TC�I�C�<����\섡{�h�S{HC��
C_\����5�,��4!�6H�RB�I7lBr<�aŜ��6������4�B�
������ب-�@���]�DC䉍FHr�#�ݼz�@�"���N$rC䉽Z~%S0�D�1
0ȡB���8B�IL�Ht�r ��R_�i�bH͏y}�C�I�~�p�XUnÖT�H� O�n��C��p�i�9$GL	�S��70��B��	zn�H{4d��>�8�����$��C��9+(�y�%��KL2��3�L�BX�C�	+CW
�┯R�z%�*�(�+֤C�I��QCƓ1m�2��^�ِC䉔p�p�h��1u�0��lN��B�ɿ�Je9���+A��fG�S,C�I�R���0���&��P���(�$C�	
2LMps�Ȏj�0"�/��9��B�I�4��5!4!O zj@��ܸp�B�	?$a��;��	d?f0�	 ��B�	�n8t����˟Y_�R�(��B�I�<\T���J�I��$QF�ՑV,�B�	�6l"��ē	���8�IG+]"�B�		� ��h�{LHz���PC�MM�h�5��+q����:z�B�	�caZ��J�h��)��
�Di�B�I??n�!�<E�9G�&!��C�I�H	���抛����k��[�)�B�	:��xUG��>v�h�KY	܌B�	�M^�P@G$p��@h�	ZxB�I�(9�Y1a���fM�<�����~�NB�	<
���V�!3/$L3��Ko�VB�	x�2|q�H�Cs�Q����^�VB�)� |,Ȇ[|�t��-+i��Q	%"Oh��"��<x:1m[�8��I��"Oа����5qzy�ݛA�hU��"O�))�Ζ3V<�Aj2~XL �"O����i��S��L�Q�ޭ]����"Ol�P͆�E�Zh[*ϹX2<0�"O,��2Ꮃ���h�#�7+�� S"Oj��&)�:}R���s�N�Z_�!�(_+h����'I$�
�!Q�!�D ]tԒ! �f��l�G��0�!�dJ2DtLxc�g�%�~[��X�'fj�����rp��W�Z'% �I �'P��c���� NyS�n	���	�'����B�$*�.�sEɇ%~�b	�'2�`�Qݴ}t\ɧ���M�����'Y�%r���z]�ƌѧ.�5H�'�"����YĮ-`��3GƬ���'��B΄9{�l�gD�A~���'��	g
�8�b����'L��a�'F�y�7FU,>�\�慍1-��'#�Uj���*4�.耔�B�m4�(�'/��d�E)b��͐�g��`f�D��'`V�Ǉ˞l��MPS��p�~�A�'	(����4��3$/��%�SZ�<)S��)9P�:d*
^�D!`�[o�<q�E����5�( �`3n�r�<a�"Ɋr����Y<,5�a�Qp�<���.�鸀�E:`) K[B�<q%�W�A?�l�VcL3�D]��J�S�<���<��$�'�ٰY���"Y�<����<T案2��X�ڽsd �Q�<��T*7�q ���y�pk3&�c�<�▴:�^9��@��|�@ ��B^�<��ʋ!�Ub�oI��h��t�<Y�8bC��!5��E/rD���o�<��]3'�����K_�F]��5�
k�<11jI�x,��곇ڄ����GLe�<A7��R@�c���	j�*}��%�c�<a"�,�,9*7O�h�N����j�<Y4$�,h*��׀�	:��ahD�j�<QB�ITr�D�?���Q��b�<��(7?���ЋT�]��A�K�_�<�F�˶E����f�'Rl��$ q�<��'Z�	<�����
YT^@y��W�<����
�l��\N�0�BTV�<9�_�o��xh3��J����N�Q�<��(�;(���@h�?p)��㭐O�<��ZN.@dArfG9EBL�I#��d�<! O�B�8(�oI�$� ���k�V�<���̧j��D2��� ,�d	��DR�<!BEL�D-��R�
��B@���&F�<�-�6�ѧ�C"���#�PL�<aq	N{y���@�N��r���<���6w�,��Eٶ���7G�~�<I�I���H�/A��ÐHF�<�1
��$g�$���o@��cpB�A�<A���.��Т�9?�vՐsc�@�<�RLL^�B1Ǐ�U;�t�n|�<Im�e�( ��&�0'h1�F�n�<9�R6A[*E�g��`rc�q�<�6�����0�#c�
w��=*�a�j�<����6>���!)tE�	bU��i�<��c)?S�D���͆!�(=���g�<� l�8T�ĘbA��+?D�Kc��l�<� ��*7/ +�T�O(*�(	�"O@k��7B�����h3��"OR�Q!��X�3�%ˀXwd�k�"O4MB�O�j���q��!%Xꀁ"O8ce.�4�X¦ł;'T(��"O\��  ��D|y�_(V5��"O��,�sA�Q(�D'�dI��"O~�q�y�������z�2��"O��h߀C,��B,D��P"O ��`��6�1� ߱k&vpÄ"O���qg�h��R��-e�)t"O�D���R�_%�`��K3V�PL8s"O0���0X*B���f�w����"O��J�4'�^9eD�-��-�"O8�I��/E]>�ٕC��0��D"�"O���K9n-|=�%C��:��\��"O`H��Ƈ3��p���X1��h "O��ӆ��2�.Թ��G0�xy�"O8�+���g����P���f'�95"O�e�T�͸i�Je��*K�B\�2"OzR�ˎh_ Pz'�9����e"O^Qb��?��t�bꙴ�l5k!"O@d$
�&%j|h�h�7F�xxz�"O�I �Ŗ9�p9�Hۢ%���A�"O��B�/�1
�!��r��I1�"O�QǖB�x!���/��5�5"O���%��fʡ�6&�k����@"On�RDR�V��	F�^vB�d"O�J�c�4&lX#���6zp��
�"O~���̩Q��591�
ivp��"O��!&ۖ(��E �!�Y���"O�咒�]}B8�������P"O����V*V:B�Q'݊"߀�S�"O����)m��"w� m�08��"OZ�УÚ}�,$;�J	 �dq"ONY(��7l�e�Q��D�d�c"O�,�6��E�l	T H<j���s"O��1�@G�h��o�zeR(�P"O<�Qԍ�`��T�.�1[��"O�," �$O���tƙ3ߢ��"O:|Y��A^ڤh�ݻMvJ-`�"O�k�OŅ��	�u��*͢��F"O���NB�$L��������"OB�Lh�W'`���w~%��'�(�(qFU������Þ�
T0��'���
>�
e!�J��)�'��|��ʕ�+<���Ͻo�5��'.Kb��?+<�y2���~�t��
�'�Lԅ!Q|� a��ihh(
�'�R耐Hӌ�=����(��5��'��ģ�^�D��4+�4��+	�'���K����8S�M \Yc�'��A������rbͫ	�ƭ"	�'S6%#�L<e�|]05���&�	�'��yuk�c�J`j���{W��'�X��tԈ2�l���hF<D�|e��'`���V���&xTP`�V�C��I	�'��!B�rE�SV��B��p��' �z�$�$�e���3sl���'�&�*&'�*&v"m���ڏ��Р�'��i�wGT!R�9�Vd�8w����'v 1!�?�b���U�\}��'���Bf�W���5��ʙ, �8�'H�(ѲB	�s��z6nT�v������� rx��ń� ���[b���9��e�U"O�a*���2��p*۰˰TB�"O�X!�c�{�:�i!
O'2�F�#w"O�����"2��B��;F� 9�E"O� �+(.i�|�#� �"O��4�ѹ9�ek�Ã�#�>�*�"O��h��G�&�ғCFh8� A"O(ţ�a�?(<2��&b^'N�HIr"O����&ԯ��7OdS~A4�(D���7.�.��*V��& tB�"D�hAWʟ,,�:�������q� �$D�x�J[8%x0K7N������i$D���(ħA�{��$U�����5D�����(��Ф�p��ee>D��J@�D�?>d���OI4�6�H�!;D�(�g*��xkR*�_r�,�V�-D��(0�\��l� �U�i��[֣6D�L �CQ��cU�N6���pA5D��ђĈ�o���XE�!r�Ib(.D�Ē�<�al
j�D|3�*D��*@䊠m����e��72t
 "*D��b��G���x���9eT8e�)D��	��&ކ�2�LV�26�!��h&D�S�ƌ?E��ђ�-T.E���v'*D���d�D�=�.�bӭ�N�Z���,,D�����$���˴	�"6i�%*D��`#�Ŋ&���S�%Z����<D�TB�,�:Z�@\!��
�s/���S�$D�,����c�Ω�T��4U^pU�!�"D��p�(C1^�aBfO݄U��$k$D��tJ���Th���A6pB�'D������t� ��l�浘�`#D��2��=L���#B)AU��]꓈?D�������� �Æ� Q��ՋW�'D���ĥ����IӒ��sC^]�d'D����8j[L�J 7l��X�A$D���%aԽY�$�k��̐tn4|(U�#D��*�!U\�Y��
^�n'��H"D������.x[�9���ܡg��ѥ	!D��y�,��!Á^�d=��+�>D�H��O9x 8���3-[�ȔL;D���Cb� ��a�"R6�	I��&D���U�8x�F��G�F&�d�!r�?D�ܣ��Mp�ED.�Z *��2D�l��-C�T�z#���P@�=���0D�j�E�\5N�Y�����`��.D�`h���'V�5҆B��D�1�.D�8�d�"^b0J�''̄�Ģ,D�; �̧m��&ԭ<�� ��)D�����
=M\�%��a�k���k�.'D�(���(J�Hś�Aσt���Y�h%D��9N�/�x��� l̴�f`%D�a���>���]���� #D�� ;gE�h�Q�>kf�y2�6D���p$�oR���b�<�j��M)D��p5l�3k�{tF�$9r�@QI:D���ز'�r��e+P=z���J9D��E�!7�,U9��n'����5D���$��%#�@q)R��m�R1�3D�0�j�q��0� G]�G;��6�2D�PIf�ćH��}�B��3��hR�1D�(����:��Dw��{,���b/D�8���hV&L+�/$)�Zq+;D��B̌9���:"�h����7�3D�� 8y�@lCF=�ݡ�NB��T�S"O Y��K��"6س8�098�"O.!	�BG�(��J�8�r�Р"ON{ŢN�����oc�18�"OL�k7�ƱTj`D�W�F���c4"O���D���"{0ё�&��l?�X��"O\Ő#G��;�R�����8�I`�"O
8��`D1{�tzY7R0S"O, ��ϒ�\>���V�5��C�"O�<���E�u�(��!�/m�Y@�"O�L�D��5�4(+��O���"OF�p "Y.qX<s`F�R�L`��"Or1�R�R�KмX��J	E�LPI�"OB�KУ��M�h���cN�AVfiX�"OR]�������t��G�"Od<�A�B�:�f�hacL��lxQ"O��Y�U"~ޙ�A�~�tZ�"O�d��I\�'d|m�Ǧƕ? J���"Ov1�7͇c��k��Z��&��"Op�z�P:H���I��G�{谔BE"O�����٭#�LIïX�v�VT��"O�܁�%�}����%9�Bʲ"O��ae)Ğq����3�L:4���cc"O�I*g��&f����e��oG�x"O�xZ��وPJ�``⊉w-t�R�"O��[`G���b�=J� "O��:�K�2
P0"���I�@"O���Οkc���`Ƅ�i�$�Q1"O�I	��`B}���[�D݀aT"O�l�IJ_e�dzGj8̊�3 "O�@d$�<Q���T)�r�����"O�la@��%V��bΎ>&�^d:�"O�)���S�j���c�ĵ\�x�г"O��f��
V%���(I��՚E"OʈJ��u�(����
W�j��C"O���.H�7>8��Ao�i�����"O�)Sd�sX�C(�*bt�̓T"O\�Ԃ�8Q����6��PǬ�1'"O~M���9qA�� &A�k��́�"O.���`U�Z�8��&i�8�  ��"O
�"�i®l���"�qq3"O�{7c�=B�)�g4j�$F"O��i�"��+�H(3g�N���§"Olh3t�]X/Z������t߶5��"OTe�-�:{?B�P#
�h����"O�8���J�X�J�X�k꘴hB"O赩A�J �L$�
��Fd"O���c�íE�>I��Y8�By0@"O�ᢗ$	��q�u�U�.�ʷ"O�ĀB&V�N8�a/+v�P"O2Q���H$�q����}>�J�"O�Ec7�B�."$pj� ɍvVl�"O2�C&��k��a;�o��l��v"O�$"��9�0e��-�[��a��"Ox]����X)�@o��R��	�"O��	��ҏ)�r�`SGL�X�	W"O��Q��E�����X�y�,��"O�x�����r���4�J:/J`!�"Oڌ� ��(�B�abx��f"O���(�?��A��ʐ�=Б#�"O|�Cs��-���21'O�b@5��"OxR&�՞��దWI�b�X�"O��B'�䨂�Aԗc�*�J��C��y��x�m�rl�,\�<����y
� <I�&�K�m\� �0���"G�p��"O.��!	3k|����cN""БAS"O&Y8..������v3�"O@��$ѧNo�p�sG��O$�:&"O��H�ès���p1���_���"O�ݳ�_75I�0 ���	|z�ڇ"O����WtDyQ�� ���"O�P+b'��D��a��@�ABC"OV]�1�\7��P��ʣ9npd0�"Ò�3H�	�&u"� SĜ
�"O@����FV��f�ܘIp�`�W"O����O g�����qh��G"O�,���(w�4]����=yUT[B"O:��Th�q�:4�5�>%��ф"O8c���- 4�x�+��&��E(�"OغuNL)Z�^d�q�!2O��+c"O|`��ol�S�*��d<�"O�� 7���@s6�����h+"O4JS!�8�Be	���[v����"Oi)Ci���j,P���1��!a1"OfU��.�`.P���`�.�i�"O ;vB�.rܵ�P��l��ո�"ORp��D�Q�������*!� L��"On%���x)�z��kp|��W"Or����-e�ny���d�"O�q!PMֹ���f��8N�r�C�"O�@�0��i�&="��7s��!�"O�M2�M�0@:�r�⎄�JX�!"O����$�>r���YŢ3C�eX�"O�C�׹"�B�C��$(�|J�"OX��U���VL�Ч��b"Ov *��h�^��' �8V�e"OD�b�䓡-%�M`v�AX\%�#"O����ͭk�P�km�'�$ţ"O�$x�*ԕƒ%:�b�=�z�C�"O>m;�� ^NN�բ��E��"O"���O�.E�B"��~%�Lr"Or��⋛�X��	�7��:21!r"OQ υ�P㜔���ۧ+�vI�"Oک�#�y�P�KG�~��1"O&�h�Ȍ,�����.�ܔ@�"OQ�0�@:����$j�u���S"O�-�4E $ZT��ꌔuh���3"O���Þ�*��|3���;5e�-�"O0��(�8���ϼP��\��"OV���L0tGF8KPnK ���x#"O�)����1l�X���U�$�� �g"O� ��,�|�����͕O�l�'.���i��i�R� ���5 e���'�A˓��7N�L��GU�Fgֱx�'N� S�
YqN]0oN�O^b��'��1%E%q���3��D�RPi�'>ft���u a3�,h����qj�u�'/�a���JA�ȓ1^W��#�ry�p�а!K ���"Or�"�eJ�
x*����_�E6r�"O����ޢTF����$"F13�"OT�钀g.���F�N�@54)@�"O��!lϦw|��v"�`$u`"O���6�P�0�C��m��"O�}S�]9�~�{��N�Yc�,��"O��gĬ	ώE��ޑW��A&"O~��0IZk��k���v�D��&"O��0s \-���-U0��G"O� �9�+A-�h�Pt��@��"O����B�n�2��tg8 ZPt�"O�I ����a�X�yc�F%h0��"O�d2��m���)���N`��"OVu#u �6Q�X��FS�`��X�"ODi���U�\�����2D�S�"O�A椘:1�:y�U⃘l0��u"O�A(��A.TBE⊿r��"OؠB�Ҵ8��`�ҫ 0q����"O�J���4XI��1߆yE"ODU�c�V&��h�#�pѮq�"O^�#H	̈u��ְt4��t"O>��p�!-L��3#��0.��q"O� 1�-�-Zn�lit�e�z��5"Oyې�ԤIΖ�	9h�b��Ќ�yR�ʞ`|Y��Y	�]��Ԃ�y���Z����dW�W`��(s�P�yr��>L ڔ�7J��V���q��y� � P��ƄG�\�p�����y�j.dz�@B�F4�xp��B)�y�OI�w�^y����7�2���yr�I�!�A��%/$͢�L��yb�[�k&H%k$�ܻ*'> A���y"��=~��k�J^�+eT͂q#B�y"�����A�R� \�����yj��lE��8�d�1�\8���
�yb�[2�H8�W'ؼy�Zm��&F��yR� ]��JfO@$h�裃��y��B2In��IE���总Sa��y��"I�>T����*��<��� �y��%�<����+�ڀa�f �yr��r��
vᖂ&�����ȱ�y�&�u8 	pA@�9�PkA���y�N�{5���B
�mH@9��ˡ�y"���&!�F�R=ؽ`ը�0�yr�ݳDB��Wȇ�K�F�SU�ͼ�y���0W��}"e�×A�"}��Ԩ�y2
 2��	 �i�
A<V8�`%�y"G�=_�m��۳blb�M�$�y��[0T��I���X#�m	�h@
�y�K6��Ef�-EH��g��y���a<����0oE��&��yrF$+�2Qcb,<�b1*��X��yB�pm4F̚�6U��Z�K�+�y�ѥ>�&ňE�}q�����;�yR��9$x����% l�,�D�=�y���Sþ��*b����T�F��y�琱X; d��L5\�0���iK
�y�
�"1���SQ� H����y�#)r�A)�K�pMx���)�y���8��t��D4I�Ġӌ�7�y2��;^TMѣO�SH5���W��yʜ"�lu8#N��N�H�r"G�1�y�/�_a&��ƯtU#%�>�y2��)j�+�Ҳ[#�I�5�Ӷ`k�B�)n���*�X�#�C�@�~B�I(�9dhT.�L�b`@�>�bB�ɾu
Ȃ���=U��9e됢tB�	?0��d{P�ŒF�n�P ė)�C�	�Zd����+Z�6����
Ô1�vC�I\p�J��A�"�ty�qO��A�B�I$�܂�"���ٸ���h&�B�I ��P�En���r��Ӎx$C�M��Ma��ĝ5�1`�&{�C�)� H�����!�]9`�ÒFk�I�"O�8Yd.B[�pܚ��ɡH�� �"O���a��A�Tq�Ѯ\愠�"O�q�� c6BEx�hԳ{[��"O~��7C��_��z�Y�]G^9`A"O$ r��I΄�#�̆I��iٷ"O�9@�4o�(qB�&���!�"O&ݺ�e�n
��� �+Z�\d�"O�1�A���tI�N� ?��ȱ�"O@@�f\�{�Y�MبS��h�"Oּ�D���&0RH���:����"O�D���$#L|c���#]��w"O��!7�38�����i�ZY�"O���C�~e�ݓk�ڡӓ"O����A���"ؠ"�aq�"O���V@�e�b��"Ou���V4ѐ�{"jS�{8� �7"O��j@o�:x�T�Ǉ��cHUx"O��*�	�h.b�!aH�5	Q�Y��"O���[H\P��Q(�o�R�za"Ox���	B�[m�yɂ�	�
��=��"O�5ˣk��>?�u[�$7a�N��"O�����6Ҭl2�"O�����}<"�S�b�d����d"O���@ �r�:�H�"Ȩd���"O�D�^(s ��� ݢ���"O�9���щ;����lQ�\ʲ!q�"O��jC��:P�j=zW˖ s�j�2"O⽸�Ej��9W��yp���y��~kJ������,j���y���=}�Tr#�+e1*�(��/�yb�L*�z�,F��uF�r6�]��'�TauN	L �(��Q(z�p|�'k1�tOK(WhAcS.V6t�D5�'���w���E9�IXfB�{�Ɖ�
�'�����.ڡ7��B󂅥rBQ;
�'V<{%eȾ"���.�[�t(�'��끮��!@D�@�؅Y��Iz�'�<��e���	*�㐗UeR�p�'�!��*��c�0(��!��h��'7$���o�6 B��� ��
>�y�'=��!���X�Z�頪 :
8d���'�	�A� b�� IבK�6��
�'I@`{��ĀY\峀�H�;���	�'�J�A���<���Ӈ��1��
�'y4u�t��*��&���{<t��
�'���	^k:�U�v��/�,���d0O8�Apb�D0�l�5#��q$�C�HO?�$W1�AP��F��Q!�ƌ~!�$<$�L��h��r�x��ԗc�Ipx��O��&��i1���9����6"O�|B�g�;K�*�36�^>A��rd"OL8��M�P�h7F�;�R��	L~"��t$[9XV��r�%�Y�Ʃ�a���'��{��$ 쭂�	�:r"�R@l��y�l��P��+O4.?u�D��$�y��_�WA�e���*����#$X<�y2�SyV�huO���X
(�=W�<ل�@��<�M�%&`K��ƹ̄���?3d�aQ/��l��Ձt��/C[Rm��	M�'6���ڰs�R�i�JѣB�N=��}"�)�	��&������&�ڴ�/e�!��f�HaY0k[9E�i���H�!�ĕ"Lw&,#I�|����{�!�� �9ӡ�NFp��i�O[`�x�d"OZ)3�/�VWN�;p�3{֕33"O����l-;�h0s�C-~`\t��
O�6��"_�R���
U�0�,���Q!W!��G:����� �n�x��ƕN~��=��'�O��?�'�$V��0Wb̡e�i���PU���=�'�{�lܨ5��&~��I��&�O�'ta��A��=R�Պ?暥�q�O��yI�5�bT�3��+3~(�t���?b@�S ��Dz��Y�M��q��3�� �Fj���y�� {��\����&#��h��!�yƗ�b���hՃ�g;ġ�p�E-�y�ʌ=���0�)���@%`��y"IIx��hc���L��*�+���yR"�h���3'�Q�4�@��WA	��y�'�?D{��Z�i��܍�⭒��ē�hO���;!@ڢX�h\�D�P��hf,#���$-�'in J��	.`N�2w�ɆQ��y�ȓyڔ� �#QJ��)�n�Іȓ+8�Q2
V�S�ne�v��(lf�?yӓ Cp�#һ~8<L��K��z�l�?q�O��}��ÿy�2u��W�j �|s�GS�<�#��(���e��D����E�П,�	d���O"d0WW�km��C�U Uh�higR�dH��!�S�O�2X�Y�L�| cfW�`��=K�'��	W���O��r�/D. p, Rzt
I>�s�e�~�=�O��h�R,�nQ��TA�'�(�ca���l��$$M4^t���D&�����íJ?
uC�&ҜB�\xeI�y��R�dw�iR:����E�R��y,34�8�b�B$8���+D����<A��dp@L娠f�Mm0�X"[�7	!��~�xZ��H6d\d)��3B��|"�xr.APS�iJ�۵/@pə�≢�y����+����@$B�}���W���>y�OB0b2$�{����Qd��[J��ò"O�Y���9^�tMp��^>6�@�"O��5	@�*����.r�|<�"O�D+gfB���Ď1^6���"O���E�R[�p���uTЀ� "O�yc�� �:>>�+ *;Qʙ�"O���3�F�|��p07�UZM���"Oj����=P<��厄RD&UZU"O0U�"O�,O�^a��.�,K�"Onl���c�M�@(�,B��H���'�1O�!�a����pr�'Ċqyl�P�x��'�����K�#W��ӓ�1��l������l �`��v<i1�O/0�!�DQ;�*����U\��s�Rr>ў��'��|��̜|�P���B�ӥ�W�<	�Ǡpȝ��NS�Zd-�O?ً��o�����ש-Ђ�9"a��y�xB�gk�A�A��(qx����H���'=a}2%�9V�2�&������y 	�D�̸��{?�i(ąA�y��5k�ҥY#��w��9h�A�|�<� ��Ę�Ƃ7'�x����J�<U�?PX���G/ٍ0�j��C�<�j��'��05�ƣ�V����f�<�O�E�f����_Z�d�cb��hO�2C�1�cd��.�,P�6���L��?щ��~b�6D�dA��(?]�< �PR�IR?A?On�����hSr�a.��X�V�$2LO޵I�JP;0���7K��tY���e�'���T� ��3��O�"�(=Y�$Z�A;8ep�/�O���G�'u��Q)Øi/�MCɄ �!�ă-H��)��� �L
f	!�$[S��Xb�Â'*_
A
&��!�!�D�@2� I�$Q��;�	��I�!�dEz�`(%��jĘ�C�=
�!�$ؓz���:�$��ff�@�TAO|x!�X"L	p��`�rZ��Hu��Qn!�D�c��0���S{�o�jP���G{��j!郄��
��bEQ�2�}*ӕ|��)�3D����B�6��ʍg/D#>Q��	��.5�x�K�9�JQ���ۄ1�!��·c�epQ��CㇾX��O��������d׏I&��7Eœf��l����El!�T�k�B<��G�M��l��߽_�!��>p:Tٖ�Ďv }� ,!�dԈrPx"��%Y�(Ys��Y�!�d�3�=�� ��2�"�rĊ�L�!򤟫s�H|*��T�%�JD�'� �ġ񤖻]����L���+egӊ%��<�?ٍ�b2��)�jG2B�m��9�p<!d�ɐ+�b���]�fL6ĩshY0#�~��&ғ�2�{����,Ɣ��e �vl5'��x������P5)��Uܰ��$�X-���>y� #GzT�P�/�^m�Bg�'�ў�'U�����0H���REB�'�j����?A��_�`��K+%<�1+���{?1���08��d-Z}0� �W(~�C�I�}qpM�s��f?��z��ԝ���d�V�_�0�4���:����UjE�,�ȓ+��\�#-\J�j��+����<Q�	�S���O!k�,�5|��!�͠�8�(��D<�S���ʱ#��T�d��D%t �iD�'s�x�/b��K��(��U���0�HOУ=�O@�M�A/wK�
E)^nR`�k�'�D�a�-�w= �:G-ԇl��A�O^�=E�D��*� )#�I��ָr� C��y2�0�	��郇#����>�y"�)�'hT��

p��m "(
�6цȓw\�8�JZz�R�+�,Q843�8��'�\�n��8�:�nմ)+ �ȓr��1��X�0�3�֭(��� ��Ћ6�H�^n���Jը7�"<�O���$��X�0pi )Q�1;��ą�X!�DN<b冔3Ҧ�<C��Q�h��+!��<	l.��6���I@�P�g��!�,1p��tJ�g��|0�c��a!�䙷a�*�[Cc�V���� c_�L�!�D]ܪ\0�mM��"��ا4�!��քh�H�:�+ʴ]R<18ҀOm�!�D�4R4��DV,nL Ct-ّe�!�S�B032�	EFգ��
�!�IM͐�JcĒ/:D@8�щ�� �!�$�=�Jr�/
��%)H�!�$�!F���h$���Z�,y�7��ek!��A�0��ˡ���b��%�'*ݑ �!���}�V�j�,2�@�#��1]�!�䊕Y����+�&��# �(<!�D�.HB���E�lb6(�R�֮}	!�d^��zT�Іc@,`#ǌ,�!�䑄B�Di�E��H�R��#g�!�$���L� Q��+T�>��'�OU�!��8��6o^�M�z����Z�!�	4��]k�/Mw�U0�H�f�!�� �!%`g4t�fG�b��\S�"O:T0`a�*5�T� &߀c�ٴ"O쫣��1?~P3%%�5k��u��"O|I��&��t�P��	�(�l}9�"O��zQm�X{J��4�R�F�܁��"Opta5K��]�8}cE$K�2�XlJ�"O����̉[���cQ��0a��"O0�A��(w��XВ�\�A\��"O̠���\��j���w,m��"O�TH�lN}ZDX2R"�G�
)"O�-1@��%X����aQ(AVt"OlQy$�ϔh҈�� )`�Rt"O~��$�M����R)�&T��'"Od1q��?(���S�f�,W��]��"O��z��P�%F��D�D�\�R�"O
�h��0V�E��D7t��@k"Oz���^�����܂X�.���"OX%�O.sz�"Ac�&ʐQ���(�\ȱ�N��Z+v�1�ر$���I*L�iҨB�dN�,�f�W� ��C�	8�rTC$�֜	�h4�Sm�2T6B䉎6 �eZ�k�,Y�(�`��N�C䉽TYr�;�� ��αs�M(hd�C�	:?h���N5@j����.ކB�	3	Մ(�3cW4[��eE�PRB��/a�H%�·�D��!RA�B2"�C�5���Hw���Kcde�MM;v��C�ɻH`�Z��� �t����2͒C䉤h5j@X��x*h�A!^B�.iW�LY�Û�1L�:�:T��C�I�G���ǒ�Y���F�3��B�I�J�*��
_�jD.Xpt�ͳn�nB��0��l�6�G7��[��8�DB䉶N�|���fB�E��a ��ILB�)��@�B�Kؾ�(�`Ѐt$`C�I.��܂�@��_S��h1ꅌ/FC�'X��8�mȶZ-d1��j]�LC�	.p�v�s���	aD��4-�pavB�ɤ*���ЄKי�4]k�J$h�B�ɽvk�q���:{z4���M;P�C�	�?y�O��@�^�S�iJ�f|�B�	���t20�9>0��g��\�BB�	�Cx�A��Z1��l�T,I�h� B�I=f��A: �]=$�$�+�Ʉ[{LB��y8�U��@��ݚQ@��)s6B�IDD� "���m�gM<B�IG�f9��l	�L���q��B�x<A�B�v��	Ar�ʧ	1�B�ɼ_��X kJ�
��R���y@
B�I�-���fύ�����C��t��B�	���cl�4/�H�+/+�B�I�_r�!dI�D�p��j��r�LB�	'4�<#�O4>|$�	�c�t㟄+C�Ni�?�K�"�Z'65*Is��'�7D�`:# V/dżt�PhK5~v�}z&�&2d�Rv�+}��f����0=F*��4�X�Q`�Y�m\��!�ƀ
Q�P�NJA^�L����h�j�P�O�,�T	�%,|O���+ΦkxA
%�_�	��LK�'
|M*ub�
��Xk%�������R{ IK`��	^Y.��G�2D��Ȇ��F~�e����p�8�9w*3��F�r�6�y�*�
o�fy����o����� ���A�Dl�!�ď4@D@زmX�1\��@�%L2��`S� .ގ���d_�`���xB)G�,8ґxT.�������(H��xBOˤ��$�wFU�@� @�3��7%��X�GHːxkB@��B8��z��(K9F� `�]2�Ñg����<�q� �6�P8WCNqB*�e� H�	6�W�Z�����
0F���1s"O���'�r�^��f���$Њ�a��x�^�NA�%Y3�H�>�J�b�>%�8YǍ�_��YW�^��B�ɦb���(�LB�!nJ����ݠY��AB�L	�g�*���'����=�3��X���BG���.b���-W�rM!�V'~��L�a���L�A�@�
N)�'��&���!������D�7U/�Q2�O�pI��g�*ayr@N�r�f�3S2X��g���ː��P�R��KA=a�B�ɠVnzT���m�}��m�X��O
q����	\��-R�&���H��\��-��|	6F��*x�"OBi���$ ���
�.�k��϶4�����l1xo�	}����O��P�'bqD��a�Y%$��T"O�t;a��Y�H�:�@йM�$3�"�7b�|��/�+b��$S42�j-Q/H�hl�@C��zBdڅ�\�p%��<����,{��S���n���:��{�<��Y���u�܂(2�웣Fw�}r�`��a-�pv�p��S�-[nU!"�>F��ȓ�T�&#;�h�P����m ���s���W��=:��q��M+|�T}�F+<D�hI��C>��-��
�U�x�do����ɤnnt�,<IQX�:V&˗S�B�ɴH��بP�1@&>	�2�I=M�fB��o�T<[�&C$��۔Ǿ$�C䉞.f����0��m�EML�nC�	�*� ��ΟJ��9��iL>VC�1=x�p2����n���XR~B�I(@�.��u�:5p�{E�q( B�I(���J��K���P`��v��C䉵��(sK�!}d�r��d�C䉳<*��2�ϝBtࣲg؆7��#<ш��?m���"OttZ�F�%:��`qխ$D��Ӣ�nY�|;@�;0I�TA��D}�����䋹l��9֡�^Nl`83�/]!�dV�@���CK��u#�-�"��V��-�O4Y	�o!'�*]05!ЎI�6`C��'��|�ޅ&��a@B���ڌ,25E�y�EP�s.��;���&pf�t ) ��'g��-��%3rCH�,�Fܲǜ�J�!�#yM�X����%�2͐ǧ	��=E��'o����rL$,�`��5)�@B	�'8�ʰE��Iaq�*.����'Z1O���97��3�AS�#�RL���S�!�Ĉ;.���" "�a���A��k쌼��<O���uG�����E�]&.$P�����0D�MIIϊ0����ߊd�$��o��"Ee�v��tEs�B͆ȓF��<)�^	!ht�X�	ڽ4\Rȅ�=��
�=n���`��Gr�:�"O ��W��((�N��Ar����I k�z!���S<8 a�t�r!;����~ 
C�ɶ`4QAJҞ0j �����K-�B�	�-5Z�qVmV����H���B�I1A��J-��p���W��B�I��je#RK�X���ӣXx�!�ߗ5bj���ƧX�L��b�Om�!�䖘A��5�cάo\����;�a}R	�w��	�,Y�L�եڍ0ҙK���%�Ɠ��I�GE�"��Tb��*I|T��IQ��g!�Eb�O�o�)�u�V)I|)��)�J��qɰ�&��I2N5Y�?D�t`�	ŉ|� X������@�<D����EB>ptxA#��3���8D���X&n^�P##�b�X����0D��z�d�W
|A�M�!P��)Q@3D�� |q���)>�<5{$F�#�$p���Ʉ�<�5��5p��,ʄ�Ę/\�5:���K�<qek�
�(��G
�.ET)���M�<�G�	��|��m�6�T1�gA�<9�NȠ2h��g$2e�(��#�Fk}R�����>i7N�}@,�G�zA�)��BFX�<)'�D�kǏ�(t��,�@�C�<y��� ���(S�$\mj��s̓��=�@kG�v�鈰H�$:�nE�ת�a����B�������A��� �3��������m:҂�IA�
M�EEH4ڧ�����Ջ�t���oۄz��(EB�F�U->E����}ctBO/3hI�$D�Hb�Qa���Q7M��~�\�fϢ>��O;jH�"}Z�2(�	rL�'�,�!�HB�<�!a]p�q1@�K� Q���o�C�IG�LK%�'+�-���� l-!�AJ�����@4��1 ��H�b�xql����5��C�	�c�%��U S��0a
��q��#?�`o@=x��?�P��.{{�apu���3�rp�%�+D�lI�N+Pɖ�-�Vt��%	�>Y�D�'k�4�"}z�LE�$��I�P7Oc,�8�HIz�<AW��1hh��,���,�kO}�0��$��I&[�]�7a��]8�!�@)M� �B�ɄV��A_�
Ԛ���l�DB��[Ă�e�Dz��.�~ �"O"iʡCԂ:l���+7)��X�"O�AKB���|z�0
�
2U@@�"O.�s�)�b&�8
��>A���"O��3�瓢)�]`�N��4"O<��TI��'��y�e]���ct��l���Kz���@V�M�X@4!�"OE?g�H8�.�OL,!��N�MCČ�撜���9G�a��@N[�<�c ��h�+������qm^S�'N�0�aj�Ot�0T�������أ2�~5c�':t)j���I���'�"��A���t[Z!ɤ
=�)�v���c��=D���)^*
*
�q
�'<�����X���"R�hϢx�*O$h(�l�
ɰ=1�dͲX�6ex!�E+:�Ӭex�� �LդAO��cݼ] ]`-D�/!���yb�S�+�4<� 3�|pt$ؠ�O�y�D%?ڧp��ⅧOz��u0��6D� 8��#���`6��|�X1#�)3�La�ȓC���A�aR�R7P����� ZM�����8��c���f��f�܇ȓ|�^ �r@	_�1�'��d�����B���w'�rZ�R�M��T��3�>$[�K\6�y2B"�00�ȓY�b�3��E8���Յي��L�ȓ#ʀ�G	�*aI����ˣK�T��ȓz��e!So�fs�+S��
,х�z|�!�;�0$q��؄'j���#f��T�H�o8�x�B�=@b�̓��?`�%�|Ę�j������$�g��$��0���2��@�U~���q��/D� ���V� ��&\5����E* D��Ȗ��azrb�iF� ��I D�����BT>��ń-����B�3D���s��s,b=�k?�jI�c3D�<!혀n��	�ab%��!��'�)s�NҬZ��,��H��mf!�DƏK7�%[e �5'���3R�;5k!�A�~a��xU!4p�f�����?9P!��(_ �(���|��|��}!C"O� �!�>�>���M�Z�b�$�p=p ��61V8�w�0h``cm�b�<��L�<%vȢANǠ��@��^�<���	�ܰ�A���8���S���\�<cJ˙ᚠ���k�衃�eI^�<��$[��e��I�?�QK�U�<)���&�N�I�^�O���p���[�<)����f�@h1%��f�2P���	k�<1P�� G�B4��I"�'�e�<��I�VO� �γF�����MUu�<ɓ�Ұi�� �Q�Kt�:�q`X�<10N�*r�S�N�;B�2D�Hp�<����	O��Q9��Q����`�g�<1�`2 V�߿{$�c2��c�<	�F�{e�#��Q4Mܦ�kE��v�<yHT�8
�Aȷh����3`u�<���B�v���B�OSx����o�<���V�4�*�T'�,�L�SN�_�<�P�F�"��Q;J��-+��W}�<�u��8{�b- ��E�:v$$�d��r�<��ҏXR
�r�I�z5�����T�<y�j�0?�YA�#ӭR�6�i�g�U�<	��"E ��+�
(�V�B���K�<��CY/C�̙��'�(XZB�E�<�M�$N~���Ə
���E�H�<Y��
#bEP�������P(6fWJ�<���]�]���ۣb��A��Ö�L�<YF(�5]��i��q�B��C�<QeD�^�L�B@�S� �Tie�L�<qafC$�zvD �8�"a�<s�$@�ŋP �f�<�#ji�<a�O�>w8�Sᨂ�4��Q�$�f�<)����!*�C�4)�:Q��-�`�<��ш����l28DHh�c�<����v�X��/e�h!�g]�<�����~REQ��Ɛ/fUa�+Q�<)�
���*=c�+��gu��P�IJ�<�HE�p����ĪS�az�2��K�<��W���Cp��5���u�Oz�<�0P�.^	��&T^��A�}�<����G|�93w�؞	�҅apb_S�<a��Q%��J�SX���O\H�<�$-D+.m1u@ϗ�����!M�<�#��*�H,
Rf��+�� S�<y'͉.L����mԗm�DH�7"BJ�<���5��I�A�����z�y�<q�O_�|#<I��	"}��Ą�t�<!��\��H����"j�^\٥ w�<��&M-'��Y��d�%5�@��ТSq�<ٕ��"��X��B�|R2(��>T�(r��/
���8���1M�����0D��Ӌ��>��s�E�|X��ql,D���ûr��3U��'!�\��*D�qS��+X�5ydKM�A���x��5D��$n�Q -��A�ob:�B�O3D���4i�Q�RE ��٢yG�(زI3D���AF>Wm�����	nӤ��e�?D�� &�J,2�v�2�' u^�vI<D�\��EP4d^`!Y�@�n�Trsc&D�l���@�#f�q FH�w��0�!�(D��#! I/���VM
#�h8��$D���bE��g�.%#�eɵF�n�#"D��zvm��s[�t�4D&Hp��Q!�$Ƣy,�Q�EX�7q�<��)ʫSh!�� �|IH�:�F�2�G70�Nds�"O��� ̄Av�X�gVv�%!"O�����1s�V�Ie� �,�@R@"O��S�P3�ʀزkWK��Y�"O����A,*&�x�'����8A�"O65@6�ž>� IA�n�6�l�"O�%�"���������=���Yp"O8ݺ� S�|���E��<�D	�"Oz�h#oO��>ݳ����rś�"O\��勗 ������Ye"O
�
k2-�@(���׹-���"Od	��0@�fD���C �~09p"O�1FfO.T�|�����&�:�"O
-������ G�7.�08�"O���ț�W�j�&�u(�bc"O�ɒ�ɛ�D���X0h2�xr�"O*���e�%~�$�1Dֈ~��r"OFp��.E�%e>E��M� |8�R�"O�%��NX�:̜��f��Q� ,��"O:�SEDl����!�0H�h;"O>`i5�F�~2��Fo�2_���Ґ"O��1�����őCߴ0}:�3�"Od���aV�=}��00�5w��#A"O�0jq��>܂�C�${�<r"O�S��F3?�"�R��>��`Jw"O���Dߐ�$PK��`���"O>А��G/9�h�gj�L|d|*�"O���.�@l�|��� ����"O(��Alɫ`�D��#t��!�"O(0P��$���rAO�¢�8`"O��)B�N:h\Zy���ܞ=k��c"Oz�*�+�3MI���m@t��4"O���c%]�ȲFM�mf\�"O������ 5��RA͝�=_^8"OluЋҖ �y+��XY�❑$"O���oƚ�M�i��Z����"O~�����������.t@u�@"O��䧏,u5���B��c�Ik6"O��r1��!�z����3ƈ���"O\,;!�I�-��{�%��d�p-S�"O�����Ն[D��$d�"O|�!��qS��b�%N.�4Ѣ"O�h��K�QR���;�9�"O��F�-1�@8���
�`	��"O�e�7�@	��y`���f�A"O�s�hE��v�� �[��ހ��"O0��e��=���ߗG�+7"Oܽ	&�8���M_?I�\@"O��hqf
�o^Ȁ��oS"���"O� Ъݥ*��j �Y�5�D�B�"ONusf�O��m;�˙1
6$ T"O����m�L��X0�j�6U��0� "OTQqui[={,=���%q�ԭ�"OŃ�H��"%ر���^���"OR���mqj4@%G�hb�"OЈ���,H�bm�⠗���K"O�����p�:���`՛��yb�@QUh�C���2K��	����y	�"ZO�1�F����iŋ���y�d��<�|�cť_^4�A,÷�y��X�6?���Ñ/q���Ң��yRHV  �*�����~+�X���$�y��ɹ!CR���i��'ӈ�9aLN��y2�R�K^D��̮i��i��'�y
� 
���jQ}<*�z�LO9|�Be�t"O<��LZ�Y�>	�4DW #Զ{�"O��e�XYb5��#�m�0ұ"O��ᄊ;=Ch���+tu�"O|�#J�W�D�g�I;���p"O����H9���`��a����4"OV��Nȩs<(����f�J!s�"OVD��̳&�������)�n��t"O���3��G�YUh�C�έ��"OʐH�N[�8��Z��Z�h� �)"O��b�B��zh�Cn�(v�@ ""O��re��z����+nR� *�"O�U���M�uNJ�
�Qs�A�"O֠K�
738f8J�솣}ζ���"OT�x��U(o�����'�H4��"O���B�,0X�bN> �&���"O��c���H����P҂aH⍹P"Ō��$t��&���˶C�!�D�g�Dk���\�R��CV��!��	��[����hr�d�.�!�DZ�-|�p���͔�"��Gޣf)!�D�#�F��5d�$����A
z�!�9v�����5��e2�#�!��S��C��C�v��nǶ2s!�$�Of�_)]��sg̴*7 Y�ȓX0rX�"+�6��Q!����/����1���ӐZ�0��(��,.\��ȓ%6��/��%���`a�b�z]��pfN��D�]��^����AN��|��R�b?T>�z���C��%�ȓ �2 Q( 2����e�]7$��a�ȓMF>Es�L��'WX�R!�-<�F��?����2c���v��O%�|	��hP<�BD¶[�2-�&J)d�ȓ$���A�l��6:)ʃO6����ȓO�޵��*^%�,���5�Z���OȮ��'B#`�\�i"�J�y�J-��W�|]8d��Y���I������4��P +ٗ`�d$�Ӕ>�ꑄȓW}��df��w���kGD��@ZhI��l���bw��8�fa�`iH� ��ՄȓEٶx�e�5$2�jƃ��`~�9��t!�΄ '�)���ď4x�ȓVb�h�D'8F<~�(�������p���`D%��n���H�Kx#ẗ́ȓ2����T[�bp���4!���ȓK�����!['i&@0��@̆ȓv6D��cC�sH  Q�_�SS�y��%0V[S��cW��̔�4ql��d�Ax�ƄJ!����X3QK�X�ȓNʠcg2R�T-���Os�̈́�g�*��Fi�$�=i�U�J��H�ȓD�1 _6�p=��'r�"���CX��zAƣmĴ8�$.�j��ȓeY��#3�D&��Yx6��Z��P�ȓV̬��9�1�r	[ q%�5��*W���6Jг��˔nD+UXp���=m���C\=��4�U�Y?�i��6V���E,�,�l�Ҡ+�G����ȓI5⭪��FI�4�@�����ȓ8�`*�d̚~��+���	u֑�ȓ@�8�r��0��M���f��ՄȓM2p	 
މ`�N� �� Z�@]��a��ra��^�Xݢ�о�ʘ��S�? V���mҞ6��]���A�N�P�"O,qi2���r(�X�e����A�E"OJd�S�4.�u���Z���KG"Oz �ܒlf��[�o~��{�"O�h8�F� /�B}��N	Jl���"O&�b��޶g���k�lT�EZ�䁰"O�q��[0�f%�KٺAH��R"O��k�"Eo�R<�	����Q�"O���i�*wx��NԂS�tR"O�ۂ!^�0�����@�a�`�a"Oz�X�Ħ*2���ZWҜ�1"O��v��%4�H�ia	�PL�	�E"O��`ŗ,S'h�P*Y�~��"O>�x��14м��j[�`��S"O��C���%�nL
��73�i�"O�I�q�ƨt�D@2��6�n�"O�D*��)fU�ӄf���@"O�aC��B`-#�$�*O|���"O�U�Ώ�Cζ�H�iI;LA4"O�P�R+ �&O�l���� 5��S�"O��&�YT ��h�!Gy���"O�0��$Q������DRSN`��"O@]rOY�}�lцjL6{b�jr"Od
v��Q"�F&��&!�<��"O|�q�愛kLstG��F�´�"O����<YN���
�$��� u��<�~��v�J*E��l�t��p��C�G�s��z4�R;��h�Z)=bO&�(�5R9x�$��>��7B�>�z�.E?hy�!��h�<�,{��(�إ��b�t��1G�F���sV�����9& �xe��]�ډ�UV�`��$0�S�O�x���_�Ht*�
M�l���d*������Zc'��4A�:1��2T"O��+�,L�j,}ɷ�׿��9f"O�a�d�e����.$�d�ȶ"Oə��Վ!�~�H�i�J��=�"O(%����v����-B��Y���'3�O�(��?z-���qa�&yy�\hW\�ԇ�vĖ,���C����e�mb�d�2'�*R�$�*[���9JQ�
çM���;�gS7"_ �g��c�|�ӄ�9�~r �8R��?��'��#}>]�rd�_�)c�Y�L���'�Y��(�9���핤�l	0aCsJ&������e"�#]�4��g#Վzܡ�ȓt���X`��(����Ї�2]@�ń�6uJ�* r�&�K�/�/|C��ȓx6�ZF͌��uC"��v�IDR�S�P��p��������5'îW;�=Yçi���PeĈr	�tI!͊�{&@�?و��~z�!ъ&F�! �9(�y�
Vc��hO1��� �X-���`AM�Wؼ)K���hA�"�d�1[Q>=��n��&�x�e[<U��u�u��j�v�`«Wq�I�|����ҙ*�p۶��=�qcD)��i�!��E>
$(D�I΅&k�!�d�E3�=���3s�ڤ�Rl��;9!�d�M��E���!"Р��_$!�$�1`�T,�qL�8(3�L���M� !�D��XS�a�.I:��Uq"���U�!�䂒{u��PqO�Kx�C!�� �h�8���
=�&������!��CJ��ݯҴ%���P��!�dƥT%L	[2�/W޸�����X�!�D��!��D:"3�X���]=R-!򄁩!!@`�'�^�1;�uz /G)l*!����c@O/�����+!�Ԇ+Լ��F��K
�i���g!�� �,X҄��ծ,��`��ɳ"O`�jc
Q�a�Q�c�C;_�@�[�"O��y�$.f�3��"�@��"O��q#΍�js�m"���� �"Ob��T`�g�>d:���]���"g"O�@�&��.(��c��ڵ��5ڀ"O��ڶ�3�R���*
���"Ot�te��w���A�L�9>�ZH�s"Oz�4�X� �f�YKCb�y�"O ��`��4�2ɫ�i֊!�d�v"OL(0���P<z,q@JB�h�A�"OT�c��,3�q�T)K)1a�T�'��h���1![�����%�,`��'{f���量s��l�&ʣ���	�'�ژÔaħ4-&D�Q菊?��`��'����(�(F�-��,�+?D�xx�A˜���S�CZ�0}|�J��2D�(q�M�,oeP�rV+�/�8}�6�/D����jK�#��19�� ��4}2�n-D�3��Hc���"��/�@�"�M1D��	�8�$�i��޶d6��.D��R���F���ق�]7(��dۇl.D���B��=e^��"��}��آ3+D�,��ܬ���p�Y*7\�s��$D��Wo� e( ���S�R�$x�S�0D��Bl]�[e�	3b�ДU����;D���b"�H��dED��N����� :D��"!��@����p�>�z1���3D�`z�g�jr.+�"�3�����$,D� �5��0Nh�MTdAу(D���-_J�z�c)^�Y��9�ѩ)D���śjk��S��H1?Ծ��&D�@����$}�jT�H�e��K�#D�HP�.S��!p�mۀI౎+D���pJa��(�2,��A�R�f�'D���犋)<bA�diQ3@�H5D%D�xY�ǀ-9|��Ȑ
�n��81�"D�dq�n�5:<Bݚ׆��u�(��k+D� ����<�QDG�WRPP��+D� 3k�K�R��
ǜH��a+��&D��jp���0"�aB��+~���*T�7D��!�ޒA-��4L�16���i11D���é�(��3`aN�=�~I	�"D��#�O2# �X�2d�Y.�	�>D�8Q �ʏ��kIzi"p���;D�lc�� y.1�d^�V��'D�T	/�(*3���$ ��\ٚ¬&D�D��N�
V�t�����3��D#D��)��F�t�(��J���bej"D�����r�5�P�N ��$���#D�|�%
.C�^J�o��^t1g D�l�f���u���+����F0�#?D���H��qb�P 0�(0� �`Po=D��S�U�G(0�@���Hh���P%;D�X��+�+����1L����-D�x�@b�]�4�+r�E#)�,�K��,D��zB"��$f	��F>t� I�f+D�X��0j��P���H�_�L�X3+D�dçA��O��҅ǻ8�~<��'D�dӠ�/XH���HP�1� `k��&D���D���2!��)�B��TL�b� D�<9p(�R�X�I6N'��;�f*D�LA��'�|��C���jqhv�+D��б�Ҏ_�d��6s�Jq��G.D�� np+�앒>�j���/T�b��"O<�%�K�tY!iD�М|s�-�&"O��S+�>e�pK�J�+U"O���cNpkz���J�����A"Ol�c.G�Ĵ�6
ȵ!ʆ�q�"O� 슢\pԢ��� 3�(��"O2�%L�<�(P�r"6#�T�
W"Ol@`Tf2�������
rٴ�""O�q+�Aܵ28r�h�.8���W"OB�r4�w
  ȟ!f~Q�"O��i�_�V�� $@�����"OV��Тd�&y��W����b"Oԝ��e�ih���p��83"O�d���Шs��傤�C}ʬM{2"O����G��6��O�F�q�"O^| A�O/|�j���ǭ:�b�I�"O����Q�3wZ��e�ͱd��Y��"OJ��O����m�eI��6��P�"O )j2%��p�"}�(Y|r=��"O�1)@��?2،���|c"d w"O\�1��׃E���WeSA_�U��"O�Id�+xR֬҄���IV�գ�"O�ᠶX!]����Z6D�Ę�"O�)p���g��\@�V,|Ȕ��r"O䪀�
=��q��%��w�|�	�"O�I�-�4Yd u��	�-��"O�����+I/��эPV��(��"O�@���S�v6��R��d�ҵ��"O����`Md��&� <2"O�<*$�N?""6�¥�B�w����"Oԍ{���T`�|�^8���y� @�I�"�����o���#�Ȉ�y�Y"U�v��fHP)c�R䩆"���y2&H��B|��*��C�fV Y�f�ȓ¤$��
_D����X!1��ȓk�����_��az�L�{+�x�ȓ%�ȃ��W�V��R��]�!��o�����N�A�����y!䠅���ږ�(���KQ�����&�21-N�Q�Pɐ��A
yj��ȓN�-9/�S��Ũ7&�<�μ�ȓE䂵��B�?S��H�)�19�p��ȓC[|��d��5���gE�d�6ɇȓL��ˢM�S
���Z{/V%��x3 x*�F��CV�̕H�4d�ȓ�Z�Y�aJ�#��a{A�ύ5��م�C �3�X+{yS��?~����gS\����� =����oվ6���ȓ-�<-Z�j�u�x2�7C�v��	�H*��W*8iR�	G�O�Ƽ�ȓ
��8۵�V�Z
�����*�ڽ�ȓ��u['@]�Y��u�7�<°���=8���&S�.�;���ިŅ�^��i[��ߝ;*~�3�QkM����)�R�k��A�WlJ=8��Ïg���ȓz�)����d�P@E��Lf؜�ȓxdQYP�˶o�j�W� +҈��ȓf�<���MbH��g�8k�2фȓ5�� b��8%��id"6L*��ȓ�F|�elW�J���H�y��6�K��m�ʽ�qP
&��ąȓa���1�I�IM`y�F\��浅�1�P�z�Q3��r��BS�!�ȓ0��ɹ������	πv��݇�S�? $�+�6~�@t�4�טO���T"O���2�3Z��s��u�0���"OH���]4@�v����ܺt�����"O��h7��?�8�H$ç7��]��"O����<l:D K�~ȼ�s"O¬���ŉl�&�����}de��"OJ��T�ձ�Z���H�-7����"O�`6�̗��Ly0G8-�r�(�'~�@��-~��`&Gʚd]>LS�'+6�yc£7�t�r�����(q�'�����/ˆ<u�XVM#�n��	�'yvT"����^�tAz@n� :��a��'ڢ�B����H/ iq��Q�)y��!�'���!)��{$�%�VA� ��% �'#�|1`�+x*�9��`����'�zb,I&X)�(���~=֝�'���n-�iP��G���o��i��'�p(4J_
��H� 	K�;�8�'R�Tx0�-*w��Ip, 7�����'�pԂP,"	]4=��'&'A�]�
�'�Dp�D#W�t�P���(����'x�!�fL;v�4H��O��!򲭒�'����͊G�~ ���N1�	�'�rH9�h
�@��	c��7d���'�A��O�G�XXQG�+y��'�<41`�1Hq�ņ�QR���'�h��M&9����b� �&���'�,���
��s��EC!��'u�H@�	�'�¡J�.#}HL�PJشm�$��'^I���%3�axp�d���'�F��ueO>��5S%�\V�`#
�'i��#J�*?@H�� A�%��I�<���R�d$��� �1	�G�<���A\(����ɰ�C"�h�<!��ʐ[����c&�[$hI�D�g�<��!�%<�����BAMZ�JW�<��mȜaG^0pI�x�&���n]�<�D���F��ڶ��uxΡ1��Y�<y�&��E��D��şl��X��K�<!��@��0�%^�c��h�NPw�<�A�<h,��PN�\d��1��\�<�V�qMx��p͎�D��%�}�<�����$�S�VG`z��s
�v�<yAE���a�ː�vޤ�v�<9壔'^0����HH,0�.�[ n�<A����4%�#����q�mi�<�3�́w��G�i�Lʰ"�h�<��2�����p㦐��F�]�<��/@�1� D���ɿ5B����s�<a�^������� y��/�k�<���$"B���
�48]�vM�g�<��H� 0����L�h�s&��e�<q�@�k�0��r��c�������\�<���f��Q:!�[�x-�i���Y[�<iW�P���1 q��q��r�IXT�<	��C��@�?���G�#]z���_)7АC�	�,ʹ�Č
w���p�oN|C�I�9e��o���¡���8bdC�ɶ*�����aV�>Z$X�eҢp�C�ɓG�l��������Ηe��B�	2S�T�`ω �v)A��G�bB䉓UD�MP)�(8Hw�L�DB䉔qz��v�"�&8u ̄�B�I�:ȸ�q D�T�d�i��ȫdͦC�	�{�t��$��%�(�B�'Y�xC�)^Щ�ѫ@Y(8�a�����"O�q�ǔ�f�d@r� �/t<����"O�c�F�n�9PD���R.~�X�"O,X����7S��J"��>��ـ�"O� 01�A�Xi��xp!�oEڼ1�"O^;B�\�"���A![��2��']1O�غB��d:���&n;'~�A�"O��7@X-D�a�(W
~����"Oh%��JA
��֦ ��cp"O�a�۳0L��6��:�<��%"O(� ���PW
p:WK� �Ƞ��"O���dF��En+Q%�yf�Ӆ"O�bT��h�0!��*F,M��"O�]��`�۠0A��_ C5�a"O������D:ȌS�D�A� 3�"OD�*� �
,n�h�3!����g"O�����S0jn��ہ�ԾV�x���"OT�(�ć����q�[U���(�"O0@[	�B�^�2�x#���"O���K�m.� ���=|y��"O4X��H�vbވځ�L��R�r�"O@b�Z@c�Z��Ӄ{84��S"O���D�$_�UN�d�*��w"O�T�B���� H��デp��41"O,-c�j��QL��ZS�1�\�!�"O���ZO�^�B�*�9O�
�)"OX	 a`؁w�$P4���J�"O��YWbοT��;�"߻-�֤"7"O ���\��|p"��}26"O.3"��_d$e����W@ָc"O�C�K��X̱��P�!7�`�"O�`�g�X�n)�Y�G�"&��"O^���t]�mI�)���"O��J��=�*`��d�i��"O����34�9�beJ�ox��"O�uSwLӕ_(T��v�D?	��"O����JO�ao���FCM-Op��"On%[�T�D��\��0T����"O�sa��Ss	Z���-�v-h�"OY�t�)�p��$/�	R�p���"O��+�H��z ����hdR];!"O��z���=ae��Ȋ2�E�U"O����ݞ�̀��턖���"O`���7?b0J�L�)}�p�"O�|���Pbv:��kN���6"Ohթ�I� _^��J�9}�0��"O*Q����4D����ygĸk�"O�=K�G�g.�
�Gޏ;��{c"O�<�Ǡ�%vj0Ц'Ա�,"�"O�4�U�[�W`�A�&
�L�t@�U"Of�k"��Xz"��cL@�<��k$"Otq�1�qܔ���+�5m��ia"O�Ydb�a ҥ鳫�	����"O����A5�V���i�;Sx�X�"O=2�䙛<�Y�(RGT\��"O�5�plR ��}���x�D��"O��R]$�`F��
$9�S"OR "ԫ)V�����ҥ"O�1W&Hz���� S�
��I�"O�YT,�<�ȹ��e�> *╱�"O|�c�MW>eL�4�o@$��t��"OT�Q�JF�����D�v����"O<�ʶ��9&T��a����a�"OԈ��٠i��$�WW%u�����"OT�0���u��v)�$>���"O0 QP �fPƵ��H��tq��"O|$0��L<O��e�f�(&�J�5"O�T� �X9
耗�@k�ڬb"O� �qI§B�4p�!���*���"O�łq�^6L��퀱.��i�@�PD"O(������22��2-N��Ż�"O���g��."gr�`a�DQ�]��"O��DCE�	���� �e�Qv"O��t� 3��A�LN� ��Z�"Oh��k�8�I�#�A�8 ���D"O�k��|e�]S̏�Y�M@�"O�LSWEѹ!V�1  kBD	b�)r"O��0� �QBU���u*��6"O]�(���q  *�-N����"O���H����k�5j4"O�j�鈚�V='l�YKL� "Ox4JQ�
��h"	��	��|Hs"O�Tq�&ԈҴ�����"0zX��"OX����>Y�� ���E/6�(�"O�h���߸����H�d���"O�1�!�ڔzyP�ۑ����i�"OŻ�b;��Ti㦓�1��1�C"O���u��3��I�f�2%�VQ�"O���j�n<b�����0\�"O�Q�B�S��q��
1�n}��"O�)���ܶw�hpxU&�+?��X"O"����*+UdA�tI�U����"O�������(XuĚ+O~����"O,���X$UĆ����H&zvBqQ�"O �T�E�eN0��e��4�ڹ��"O �"�wA,L��2���"OL��aO�?���ad�V�V�"O&\6ꏚy&��D-`��8��"O��+b쓛:�v-��d=��`�g"O�d+��:q��,�bܚi�~���"Of}А��$%�0��ܜ<к��!"O���QK	 2����+a�X̠�"Ot���W#n$�C���a���x"O���0K��-�raքm(��X"Oj�*V�UXߠ9����9�52"O�4@r�82jD�0M�=yp��"O�\��+��~�u�l>5K��Å"O���ٻ(as`�P;��a"OVy8ǋۺ� DRB�ؒ61
�"O��3���zE�y��ZS*ԉ�6"OT|Ud��ob��0��:���*"O�	;kF��l982�E ڠeٔ"O���.
�R ً�O	�4���3b"Oĸ����+��SmI�%!`��"Ox�H!/�#D��bL3b�x��"OH���!��n�J��6T�=|��@r"O�A�P� �6�!c�ȶ9o&�
a"O�i�C
��}ў0C���5U���"O��х�
�-��RF�ƬH�,Y�U"O��H'�%�1�r�܊]"�"O�!8����m*2%�*��e�Q{B"O`���G�)֌	���5Ѯ,B�*OJ}y�iL���1�O6g���'�(Z�LD<j�R� ��N�Z;h���'D��� n�3W�^Qqpeړd��-��'-f�֨��J2<��ʆ=e�F�yr
̣u��`���SV��U�yOZt� �&��N��9*�	8�y"͊<p�T�bb8�ꡪ��y"/_)eh���O\=\Y
6G'�y2��+�D��M[X�@u�=�yBo�U�~E��՞L��k��y
� �D���8�0$��!{&:��C"OT��Ak��+[�%��)M:0tx��"O
,�2��b��cPj�'&`�h�"O:�a��Zex��8_Qz�)�"O�I:#��~w.5R	
�n�f��"O�9�Q�ܛs*l$�PH�B�ʩ�"O�|:W�M���t��F\�)'*!9�"O�,�0J,G��Us�Dţg�D+�"O����#��5ȺO��U�"Oh��p�T&+�8�2�J�Vh�І"Oz���(�rT9p�S�|��ؠ"O�ĚqAU�~��K!Ykn��"O�!��9p�L�#RMQ�{�"O������d����V�D(�}U"O�#$��)m��R6�	Z.�|(�"O"��"�F+\���ae��5p�>|��"O̒t�M V��0��=���:�"O&�kv��6$��*�!���a"O��9qc[��=����
Qa�I�"O����Ë2A�Ƥ�R�
"O����كG}Zc�C�N<D�ʳ"O:P`�hE,qq�wa��!��|`�"O�(�pɪ%Jx�Aw�lXd��"O$E��d�%	/�	�<c�j� ""O�!*s�ǣ#ì �k�;�.Y1"O�"��)~�	cJ�\�6yRt"O�(����By��#c��!l��p�"O��s��8ED�Mz���$hR��"OD��&�h��@ ?0܄d"O��īZ<wXX5����Y����"O�|�*֍[>��$�Q�cv"O���B]?�*ȳ��j�6ht"O@�z�b��3pnY�u%��QR�� "O��@��g��X�w�4K@@�"O��R��T?UĴ�Jq̤l�'"O���M <sT r�� z�� "O"H���6�I�c��b\p���"O�m����HrP���tI81�"OԠC"*��0��"D�|Mȓ"Od�2B�\�i��P�M�42)��"O�z6�8�	 ֏G�KE,az""O���fԏi��I�U�	=r=���"O���n����Y��
V'����"OFi���<v�Fp�$G[�b�`cR"O��@"��g�����9��g"Oh��@bQY�l�@��,Y�A"O��33��4q�^���9�,��"O�as3`ڮ����]9�"O�|aO�p������Щf^H"�"O����do H5бEQ{J(��T"O�؊Јԡe�(�dӽ,6,�e"O����Ѣ���#d�*l$�Dq"OИy�̟�<�"Ă�3�)��"OU�3"�>�^Y�,�_~!B�"O�IK)��Et%�Fk��7W��"O��r�Y�mA�IѠ#T1n�n(�2"O2���
�dT�"p�Ҷ+2	1"O��q�GK1b��"O͖ 4�z�"O��xR�b��40�����d"O�i�B�*��$��#�J��E"O�-!Õ�]g\U�&"�[��#�"O��z�*�$sl58g�?p��CW"O�չV�� ������z `�QT"O"a��&Ƕ��qX`JT~I���"O� �%jB"�4	av����;o�"���"Oڬ�5��>�xa��	:��zF"O�5�Q#�"2��J\�*�
Tc�"O�@��̿/
��4�߂CZ҅p"O�:�d�[�Ȃ�gXE��b�"O�EQ��^�s����.��"O�L����P�ma���"PXӕ"O���51W9j9j`r��cT"O8�!��;_�$��������"O��k�G��qA@R MΜ�j�"OĜ�g`�+6݋%�So���{�"Od���A\,��1��� �i��"O�����G̸#�-Ep S&"O����)�	�J����K�y=
��"O��qc\9Q�&I�ܜz��E"O���!��"�=å �����v"Ox����,�
p.�23
9Y�"O`��b+�I����b�Ќ��"O��KBF�7�b�
�ر�"O>�X�i��h��\��\�5Қ�)�"O�y����Y�>�놟h!����"O�I�.��+3 E��@( �2=y@"OP�pgl��2�x�����m��"ON@��,�/|��(6"ۭ>i�Q"OJ i��%Vf��a�؇_����"O.�kͲH�pQeN�t��C$"Oz�I� ��_���'ˇ�~>@yC"O�]�"�I�\*�ИS'JA�R"O�����W6/�u�ʪ@|�A�"O8XyR�A �����F:5`l�"O���+�B�T�rY/:�.��"OIh�O�N�"E!�Z����"O��Ď� �<B+�g#�( �"O�(��O)&μ��1���"O�IQ��$Y
�L���ڬ0
`,��"OrE��Jѡi�ڌ���P
Lb%"O(Y���Q�(~��V� r�v�"O�X��gC,J�����N6er蠡S"O��j@�S7V�l5RćQ7]W�p��"Oz	���N�6�^���g\'Kq�b"O\�aM0~|ZĦ��2HX�h�"O��T��5F6]S�&�?O�|;"OH�c�	1Rc��u燰:/ta�"O�����H�v@l���Y�X�p"O�9'J�.,\�y�eWO��@�"O���@�1Q�n�zW�ɊRK2m��"O:��K�bXL��4Ɂ�:2�q'"O��k$  @A�0�ߝ��P�"O:)�`��}�ƹYehݭc�a�F"O���W�T:,�I�L�u�̱D"O8u˅-|�:MS���c�	R"OT��V��+<l����R��A� "Of�	f��0
j��c����b��� �"O,�����m���Z���?���"O6�� °���� -=�b(A"O��ц�!���5�Y� �`I`"O|9��cmn�Ȧ�,fl�"O��a�.n�h�`DC&xC΍#s"O|��Pf¢x�xE���h9���"O�h�d����³DY�b(N��@"O" ����	`+��ͥ,'���'\�*�f͏,Ԗ)��G�
�
�'�cۼk�a#t�E2"� 7"Oh<��/�'t��9d1\L�"O� �X:��@�-J�z �i!6T�"O��@$@�</����o�+��"Olm #I^�*�T]�����je�\"OЈYflE�>���펒O�x("O&���(57:!�T�8,;$#�"O�H3hɚ)I>��3JG��@��"OT �rhO2 ��9'ϥ[c`q�"O:�*#	.uuw�ɤh�03"O�y��Ô3�4)D�<��z�"OཡCHͼY��(�.��+f�YK"O�HP�	^�W&�񘔪�Oz@�Ȁ"O�M��ӭ`f�LC`j��cZ�C"O�7��f�=�%U<oL�Q@"O��q���R�u1tL�jQ�E��"O�(���08���BlZ�F"O�<�ᡕ�U����,�(^]ȻQ"O �P5iU5�8]{�)�+cYbE��"Oj�ᤏ�{{
�:V�ݮ!��1P�"O�Mc��Ǟ?��@���	�R���"OL�F��02�F�B�YFjl!I3"O(}��@I ��c�"�gs���C"O�G!�L�Iv�O-gܠ�"O�ݸuhT�4�Ր0k]!"7`H��"O0�Շ�j�V��e��.eJ��D"OH�'Cܛv�J�(C�&�`H(q"O����'/m�@�aǆ0���"O�jH��PvՓ ��N7�|j�"O80�fB������#A�9-���u"O�5��d��1�V��],R&na�%"OE���Y�=�J�J�eSBbt�"OTͫ��/����%�/j,f��"O�(�5GR�?�@�ˣ�@�Tx& �"Ob���/i���3�HJ�Bq��B"Od`�����Eh�P�	/�4` "O�#�C��T�����zo6���"O���
R�h������V����"Oll0���O ,�J!�Ek���d"O���?+~�b�ދQ�@)�"Od�JڋA�`���P+3��""OD��@ �9B����T�r�5�"O�	"��A8�:5�P���SW"O�y��⌣P�pt{���*�(�"Ol�Y6�(P$<�A�<ې$H�"O�q2��
:y���!AI]�8��4"O ب�W�`	�`�f��#"O��FE;�mAC�_����"O<ٓ��*�	Z���>����"O��Cd^�f���w×�-F��P"O��ѩV�mn* ��G��k'��8%"Ob��:K�,HC_�ax�� "O�Q�'oW���t�Ia[NUq�"O#��N��I&aݕXx�""O�V�jT�Ö � =�Q�"O������JV �4-���`"O֌��L1(�)���١Lv(�"O�8 %�,)��0%�Dl4�8B�"O�]RC �<YY4ɐ��}�T"O���p�"*�� fضW�8��"O.`#���%l�!���"<���"O�0�&@\V�U���׬c$.��"O"��Џ�96��q���-[�m�g"O��з��<U� (��
��a��"O�W�]c-(,��a7"�8�Ps"O�ls��Ԯiݤ�
E'p�X"O� �D:���%�-B���"O=�t��L���դH�EFa�"O�᪗�[�}�R9idb��~�v"O,uc�� %�fi��x�&��"O�uB�D�A�b�� ��VP�\�p"O����ޣQ�L0�@f�""O�Y��?!wx,#Ӎ��|�a"Op �#W'��1��s��I�"Oj�j֤|��Y1��b����"Oa; �Ω}���ᐣ`���w"O��C42� 4@w.-L�`9�"OT ����!i��d�c�?�D�;Q"OT)"'�71؍�⍄���t""OL��A��>C����P�Ң�.X�"O��Y�@�j>�AA�ʿH|��y7"O�� �\+\�μ��O�@S,�{1"O,�0�i� �@Iah[Rڼf"O��G�ʪ}Id��g��,
Ip"OX��ʈ"R�V�K4d�w'&�4"O��h�a� u29�"d*,!S3"Om۠/��"����Q<�tP["O���0#�J�r��v���0�ؐ��"Oh�jǉ���0�ja �O�lp�"Oȍ�"��()������"�""O�%�Q홵J�f��%�`�FU�S"O�'��&6�ew��59�1j�"O2����(^��kse�w�Qa�"OhP�X�c�[2GG�jޢ���"OxI�F��?-v��(�Ƙ�8"O&�R��K!��D�qB@��L`"O�� b�2.1�5� n��=Y�"O������s��q���}���B"O�`��~�ti�ƞ�8��8��"O<���0j��t���3�"O2R�
M�� a#��OJ��#"O���@��w�h��7�S\���"O���ffǽ16�QJ��C�C��02"OH1�,G�(2ܸ�`��5D����`"O"1ض�9ٌ��сD�!�\@
"OZthD�A2�2%����7є y%"O:I #J�2�:�f�#�X]S�"Oh(qTH�N��(� 0}T�s�"O\Dk���A��;���_EA�"O<���$@�~&�aw��}S�`��"On���*�+Rڴ�,��7bPye"O�	jbk��i�p5bq���\����"O��2���i��x��ݱ{����v"OT�a�G	;U(����5˰z�"O� ����X&��Í 9[�Y�C"O؜�Ѯ�zQ�M�-d�Iv"O
ͱf�U�z�xb֌�
�e��"O�d��a־vfA���W�1U��"Od|B��Ƶ�,R&���O�F|��"O~IqV,Q)8�C��T%|���[�"O�IE�n�D��IN1����f"O�D���~Z�i��F�0CS��	3"OL������r�5ݏr���c"O�l3����l{�M�f��`��"O��C�V'�,c�b�*r�z��4"O�a��'����qk4A��ǔ\s�"O����J�@�*�����HĶ� "Oz)�tĢ`s�8R1a�6���R"O��n��K�����Z D0U"Ov���h�&��U���O�2a��"O� `��AY�;R�u1A�<��@Z�"O�� ��;;�Z�����2��q"OR�b��ƧND��A��)y����"O<M!&�A!�@����%:xy
3"O
�����)5�Yp ��j��"O�`���Ѧ_R��R*K2X؛"O>	�t
�:}�t��G��G��<�4"O2	qvJӨf:�[a	ѸM��!��"O�\��M%_X�0� gl�z"O�1��ȟ�%�y ���0|L ���"O\q�&)Y�d��qK*�> T��@"O*�j�3��ܒV��,z�,-��"O(f�y|(��U�4n��Z'"O@�:!N�|����L�`Z���"O��4揼�H��C�V�At�-	�"OT��b�g�jDh��!^�&
v"OR�G�Ҿa��`37�W�^O|u@�"OԸq�OS:D�v����(c�x�6"O�TS����w*����RB��j�"ObiKv�E�HXzTP�G<b�x�"O��Cg���
�I!���p#����"ORT����$�@�8b��o�}�!"Ob�YT ��ab�1;FL��OkD��"Ot�cu���~���KI�����"Or5ɱ����!�%�	�ɡ�"O�c$�T�x���*D�H�ID"O�9r�%	P�8�զP&q��!""Ox  M�N>��b�@=Mǖ|��"O�B3��[jUㄚ�l�����"O�T�6�l��MR�B�4��(�A"O�)H��:d�"��Ԁ�6,�\�F"O�M�'Ѻ�&���ܯ���"OJ�)#
M4:���s��և�D�Q"O��P�����T`��& H"O6d�G��p��%��L�ZD"O�Q��C�l�L��D��	2���"O�g��@<˒a	*���Q"O����ɓ{����W�y�a�g"Ox<If��
1,}HM˼S�܅��"O�YH�oŃ<|�ږiP��"Oj��ȝ�s&��
�m�xcv"O�T�%�M	�BPr �ɑi�N�t"O�1x�E���f�k-D���"O��21֟sb���aoĻPΨ�q"O�P�2D� y�0�@�g�/�x��"O��!O['m�hkA7��$"O���q vV��+�k�$ ��؛F"O�%�� �$'��x�k��z]7"O�ݹ���%-�%�W	�.cL�B"O�� �oCw:�1(�AփO4$�x�"O
��3nP���Z��y"O��YE���y�X��@�%,Ve��"O���aC�<�V9jUI f<�Q#"Oڠ;�ˇ8�$�ʋF=�5��"O����ԓo0�� ��@�H\)q"O�R1k���D���@bFq�"OBxo4"h�p ��F)k���4�+D��C脫����� �o�lN4D�x�n�J���ȑ)b/(Y���.D�����߫u�>-: f�:(������*D�T���4L�MI�IR�|��T�S3D�(	@J�TVepU�J>��a��4D� ��I���u�G�sf�s�2D��ڠ�	�=�������)��\�1<D�� �t:g��t3L�0"���'U��"O���&��Ai
���@�,@�@�v"ONp��fVV� T !4!)>�2e"O0��C�IQJ Rb�T�uC ���"O0�$��F],�@G%B�:5��"O�����Vs��7�J�"Z	�'��Q�d��.�U3qV��'���W).���
[���'�	i�GB�p[R�e�� hY�A��'e��R�gޫ'y��/�i?�x��'��y�FA/$EY��ٺh}����'�,���`�/���R ȹf���'�hQ�&��#U�`eСj�(Z�@eH�'Z�P9�%�&�h�	�A�<W�����'�nh`�T�Ჱ�@�Ƞ�0���'�p3  ���}�Ϝ}�J��'��!�N�$I.ljT�ؿF9����'�2�j%�T�e���JG�	E�4���',d�3a�v�P��6/f�� �'�x��>*����@�eC
�'�5����<Ut0Ш�-7it���'����mP6@�FFW�du�	��'����w�F�=�@�M�n#��
�'���@��M�\H�cD63g~��
�'�zA`�j�&:~�`z6F�>+�nq�
�'!�Y�SZ�H�R�ɛ,~��)�'�|t�`���s8����MV��S�'����F��.�1�xS����'�b�3�ꂺf�� k7<<��'e`	����q�`9�#ʁ1H�:@p�'dv�Qf�ъS�I�UӺD�0�	�'�6�j���3�n @�m��<�.л�'���c�x:�Ƞb
�G66��	�'�����Ƃ	t`aJ׍
^B���'P���G]#;��t���8�ڑ��O�����FN�ȣ�X8# �A��y�!�$+Uv���"��T�|��nM7;�!�T�9�4��7�z ���nO�i�Q�pE{*�&�"�H]2:�$��6�R2[�z���'�qO��P�  ?E�TDJd�!(�ri��	b�8��i�y˄\)�J=#��q��!Ⓨ蟮�f��%�����$Ŋȸ�"O��BfK6<q J���>������$#�S⓲q���ەٗpN�dK@��2W8�C�ɏyk�ͻ���O��t� �M���8��	,iUTݱ�ސx{h��Я�m�,�<Y�����,�ic��
�����Y�K!*"<!	�6Z�v��e��Ɔ	f5��L\Ti���v���` X:��%���I�L��!	ӧ���J�v�
�/�����&��%$��HF�Q����\9Q�j��/����/��Bm�&�����X9%��c��D|��x�iس(���d�&/8X�u��y�� P�5��B�P�vf��y�C�7��9	օ��n��U����'�ў����ӊ<y��ꆡ���ȨXB"O�q
`���%]�=��/��xH.xzV"OȱѲ�'v�xa����/HT��"OⱹuO
�jc�Ũѭ��}Ӛh&"O�ā%LF�.ԛ��/m��$��"O���ם~Ot�R&�	Kd�35"O��L��7+��"ǅ�6�� c"O����ѥv{�PB���q��* "OA�qG�(&����3�ʘr�ѩ�"O� n�Y
�b�ʬ �b	;;���p"O,���: s�)���A!8&jp��"Ot0!��7�� C�*�X��"OB5�c
ȨS8� 2���D[c"O����Cň?j(�2�, ,� 1"O� U+N{�3�Dr�DB"On9��*�x^�:�䃜b����T��W�DI}���3�7�&���$6O�YK�ڻ�"C�>'����-�����A�Y��#=)��T?�s�Z8�CB�4I���-�$o�W�:yY3"1#>����`o���=���[�d$ʓ$�@X ��38)�ң�I����\ �XX�F�P����2�H�V��h�)7D�����5r<x�ą8[��#8���>=�qE
$�FC��s�Z��y"� N_6a�Ï �/�|�����y� C�	KN9[��3	��}3�b��yb��#�"rBI*	|�Ƞ����y"��|�
I��/�4T���oN;�yB*�=��Xbl�w�p[��C�yBnKt�9�h�b��p�$

�0=9�̠o���$�]�*��3�J�yҩ��fr�5�q�$RZ�䁃/��y�i�g���ga�#���eɼ�y.H�< � ¬��p��������yc��`)���T0�� eGR=�y���){f=뢌��&�	E��y�h�+B�b�У��wH�%��#�>�0=9��I��}a� S`�ԵkЊQ�C΋�y�.F��8j�!I�l<l膄G��y��(��x5EцctfܢG�V��yB��%I�̙��ϓ$$O%�U�N0�Z㞈��	0:����IG
2�0(	���p��C��/�D̹dC�	;������V6<3�C�	�6ɾ=��e�#]���E��;5�B�	�x zlj$���,��`�ۃu�C�	}��	�sL(0
�р��.�VC�:8�Ȱj���� ���uzC�	&c;| ���%X0Ȩ�`��1<Z�'�ў�?��&��P���T�H�3�|y��1����ħV�J`SA�O�6i�� ��.BC�E�ȓӢEy��^qrz�(Fnʣr� ��b�0�ضE�&t��)�S�	�xVQ������dJk�n(�uD옆ȓ'M�iJ���_<
T�6�H��Z	���Uy�恍'��ȉ��\
+�`���k[��yb���a��HGٛ���KA��0<��Ė*|��X�&��.��Rvn�u!�$�S]�|���Kq&��G��=+!�D �)"�hXQ\�2)BP�T�^'!�$����I��T�<�E�RE\�!���y� ���e[�%�X6�_F�!�ą�2?��C��
WdD8T�;x�O��$-����/��y�#K�d!�d�.$
jDM����k�E!�F/~�ޅ�Ѡ]!6����Y�"3O`d
��)z�x��AmH�V(yE"O^8�(�Harh"ͩC�4��#"O�5���Ֆ\W���JB;����"O�$��B��E�M�e��:-�8 "O�AH��d�X���:z�F��$"O�E�r�3~�LBB��MȔ4��"O��I��IQR�$�@*�1TP>Isv�>Y�x��P	�@Ew���R�^5z� U��S�? `��w���7��q롉PG
��>9�<�O  ����������)7UJ�'*F�O��  ����i�$KU�9��ĭl%!�$�"G���m�06�����b�'L� '�ډ��!C��y��ʹ{\��g�w�!��5��P�p�׍O%<t��ɒ�qO��=ͧ��d�Rrh�d^?++��b�(" %�OʙƧ�<BI���إYr�m�"O�D���i,�,�P��@��=��"O2,ٖeÁ����5
MD|����|����E{�O��!9�熠�ih&�LQ��
�'᫅�L�[�Fm/���#/M�yR�_�h$���M�6��������y�.̙+u���k��X��A�(N<�p?1�O�t��˙�
K*����U�B�3��'|O� 	6��UG�Y��%Q�L�P��'�Q�(�A��z��M�4j_~�bl#�C=�8�S����"�ֻ`P��P陓#ꞹ�ȓ`z�����V�oO i����6�F}�ȓ����Y,=i���c��1�
���즩�OX�a���ѫ'�H� � ��8����>���$r��Qg���}���!�.WX��Fy�,��n:��h&�^�J�C���yr�@+R	�5����W�"�P���y2oE�D��ua�,C�M������yrk��X�x�8���w�t��h�y�(�2�*d(�E^"uِ ��1�y2��A��+�AӢub|�%���y���>M@�X��	�E�R�@Dd	��yK:Fb��y�_�T��q�����yIܙ/�Ѝ�sLRO����F�� �y⇍ ��!iBh):*�x�v��y¡�*7h�@D�+��XAv���y��Pq��D���"���ϥ�y�m�?I���A�(kn��ۡ� �yl >M� �!r$�5h���1Ě��yrJ�J&\��ݣ���@�˜�y���-���i���z�2�j��R��y��"8f�:Bƛ:}����?�yB�.f(p�{��z9Љv�
7�yRKR�vǚ�0�&�w�P:Ae���yҡ��@~�5a�� h�RXUI��y�ԅz&��	]�c2z���@���yR�V3Xy��r�<Y���E��ybF�~Qv-�e�����b���y��a��8Q�� &�p�CV��y�(ܕ;�x�񣀌���C#I��yr�æ
/⑈��0[����"	�y��	P[�pi�PN�k�����y��D*���`/O�Z�D�ц��yb�=���a
I2)vV�Q��y�n�?+�ȭ�V���Ӕk��y��Z�G��0i�A�E�mi�GO�y"aAi�F�`�SO������yr��0��C���f��#�h[�y�	 J�0@ ���&fzNl8���%�y(�~��!sD�Z��0�7n��yrJ�U޵
T`�V�lU�R�M�y�KJ/V�{#��
ODtd*Q����y�o�-%)�1�F�]<*�[`�ۥ�y"�>%��%�Ę�1��t�az�%�jq�|��+R�$h�&��FDC2	���w��9�y�O�x�ҩI��Hx�ek�m���y��H���i��o�x��9�y
� p钳J�)(
�R�l�?)B,���"O����!�(!↠�Ы<D�hq@l�N�z�za��txh4��@?D���r�."�!h����.����:D���C��(R��i�j�#c�. �Ǭ:D���`�H�M冰�!H�	fPr���H8D����M�a��;�F� I��8D��ز-�*4x( �/���rl(D�TI5�[��f`af�"_m��R�4D��r�B])�� .� � ��#�9D�����7PV��� �^��0`aD#D��rS*�BK�4*���+Dv�)a�>D��x��ةo:&�W=;���;��+D�<��F�H'P���c���*��%D���p�IWhF����U$�[��!D� �SΊ9vl$٤&\�D�0hچf*D�x�h��{�l��o��WN*0)0I?D��H��¹t;3K[f�����=D��zA�û*���e�"܌�N9D�l+��I�SsV���N@y�؛�;D�x��#d����C�M(0`R��q�7D��ʁM�9144��B\JٚT,8D� �Wg�t`Ԑ���%'�,�-6D���$�mm* �v呒�,�q�m!D�kℬSQ�9��N�J�\����>D��t�  `�HIuǙ��H�+��;D�X���8�D4I�E�>���r�$D����(� �Y��R93�hҤ&#D�4�3��>^x�hCU�:�He[3�!D��0��5oz�t���s(V�F!�$[�6L���)ux�(�Ķ%�!��#<��)#��-Z��� %�!�$�K�(��E_�Z(J4!(�=c�!��*�1NG_��!S����tJ!�D�,-���T�q����f�$�!��A�X4
��Â�?��r��	f!�$ˏ ʝ+�"��A@iu�]3b�!�d�t����V��}窵���צG�!�䕴e{b��� >4��Rӧ�e�!�$�P�lĈf@�"T���� �7�!���a�t%+�N�r��H�`Ȉ>�!�$Y':�N���o�}�~��B�A!gj!�$C, =|��R��E��Ă�I�!S!�� K+�MC��L��a���_12l!�Y�Cq�#%ۛk˶��ViB�)G!�D�$'��R䈟�6	���*�%=J!�d=��k�C@�*
8D��F?uW!��>+�*e�D�Z,�!�+N�s>!����;��a2�B�JSR�ՋO%{2!�F�R	���@xƉ��A�!��9�A�_KjQ)Bʊ�!��H!��=�@��	"(T�җ���X�!�DR�\�F�I#�ձ1����(N��!��Kb�(`b&�X����0Ȇ��!�D 'd�ۥ
��R%�A��C�!�DC$YrPB��q��Yh��.�!�D�~T*SCN@�!y� CvDD��!���=E"�2I�Ur��0B'9�!��=r���a�
"n���CF*1�!�d� ��]!�f��h�x���(w!��*F�69�H](�68�T�B�}a!�$D4^�$	�%eM�W�Tdq�d9H[!�d��Cd��@ФӴ.Q��F�5!�
���$��(x���b,rK!�� XD2�
��+��Iqp}���"O��v-X�3����n	.T]t�a�"O�%9v�Z4n���@爻�\���"O�Zv)	,�8 	���=2�4]�6"O�EM˰-�M���� $Ly"Od�I���/���j�匑M�-�R"O��C�oK"eA�(yq��v�(���"O���B-�<b$�I4n�=�&��%"O��ze��.tVQŧ�(��"O6Q#� �w�� +��=O�*d!�D�?(ѐ ��@����Q�!�dFG:�Qoˣ$/>Ղ��͍D!��@?�u��L�!�6��g5!�$M�,)��2�g_�'�0C̞��!��S�r]���߭#���kL;6��'�	����)ɥRF�jQĈ.x�۱�Bb�!�dR�0���QvD�IU���sf� uZ"��äP������>dY�RE��-)��
|VU��^���'z����գ\_�,`i�4�>���	8K�yj��6G�]�ӣC�ay��Գj�$�'�D�Q�^Gؑ����%�4(�g�<D���A�O�)،I �o��e�G$�$.4՘�ӊ{����,���D��P.��37,�
�y"۱*2��a�A�2VB�@qOp�c�F�g�I�^qx%��`�Ne��!r��C B㉯d��h�b�i4���
�5LP0Pv�v<#'I�
��PH�~B��j#)Ae�I~C��b3�'N A�֍�"��ȠQ�Z�SU�Ԑ
�77�4�4��?�Y{5������_�!�<��:��#d��^8�s�!�r}Y�'&�F�&���J���Sh!��٨7��u��ʀ��=A��L�'6!�8K��l��H�6]���1 +�v)�Lڊ�K� �!`%��isF�)>U���A�'q��#GN%D��x��"-����h�2tllRp
 b]�|��4{�&V!�8�g�'%���h���@�L�-� ���A�Ъ��_�yth�&�J�AT@F�	�0�P"��(bT�4�1d%�OiQ�FČu�`�Y^<BA��$PhqiVfE�p�-X��Y�_>�S�G` -xP1X|XI2k��(E�B䉽W�.I�A�T1�Pdl�%_�H��j�$
7��z� ߈	X�@"��
��h��nY�qX11p��[�}Ɂ�#F0!�$S�����X�e���Ý�N>!� iY�J�����ȝ0����0���=q'�K�6�H���m�D��B��Q�l�f�~M��{'%�]��M:aG/|���$�G""��5�%r�����I�Eb�<��Gh�Âh�"�	�L^�Ū0['!�X�P�����Ov}c0�ۃ'���c�	8d-���	�'\�"�j�F?ձ�a���`ѥѫ �&�84�ў- �j�)7]�>睼%��2�n���E��=v�B�I2X��\�J'��ti���
=�e�ʕ0��l�ш�� �֝!�q>YE{RɌ9"�,$��dǆ�>���D�0>IՉ�7[!��Ԧ�0J�R�i�����Q��
�Q#��)��1��#�h�3���v�L��lыw�UEyR�\!�f�Q��~�T��QK�ԄXs��Ui7e	?*<tq�J��yRaV8>O*0��GV�R�T��Z2d����ut�i�ʤZ+��)���'}<0Y��dJ�T+�_̼"�'"�����[1q9����"ܕgЦt�c�[ȟ׃��/�AAf�
���IP��T�Q�zᤥ�4�3]G��DT�f�� �S��D�&�0Ə2j%�AҒ���5ߴ\i���a���dCVH,q����P�
%���!cў�Ѱ��I�|�`RD�;B��OdBe�d�=:��Ä�(,F��B�'�����0"�a����5�����'E��	�l���⬥O�>#c������)Z���AG��$�y2W�&uS,��b���Ư ��b���֏:,O��KW�N�7l�y��K�-\B��s"O,9�CJ�.���g)r3H�Q�"O� &�Q&���}���#�%�T"O�A&D��%���\~zlq)�"O���#���Ek�,I�/�8)U��:�"O�p+�!N26�� h��׭fJ��%"OPQ�@
Ҕ?��H�!ჱ63��J�"O�С��OK�>� W!Xn@$Av"Oh۱��4~�f�x7 M�k��L"O BW�qͨ1a1�
�v��""O��H�jT�����D�V	�G"O6x�A�51p�L�b.Z�f��'"O�ls�	�=j���"��U��`��"O�qAwh��,�(��mO�;p^P2�"O���6h�%�CE��9m� �"Oޝ1W��"����РS�Y]p���"O�dS���A>�|Yd���T;<#5"O��0c��<��-�|T�1"O���$D�f@dF�L��v��A"O��F�(�^=��eEv�LK�"Oؑ�G��M�Z�(u�Ͽ%5�ى��',�OX�C�.ӀV1lu(B�V�?�AkA"ONxc�f�)��d*��+y)1����#�ŞnBr���V=�`�P!��(�ȓW5
x��*ݫ����su�Exr�'m�5���ܓk���p�KG�o����'�HԨ��Y0RYJ��F._�Z=�WO�sdcɨlN��G�C] c��`��t�?�"�>Q:�rT��2�8�p��]�<1Wk??�H��HM2���B��Z̓�hO1�j�`�m��y�ԙ �e�����"O*<C��rY�)�Cj���D"O���ʺtp��k�HA�KG��"O^�+3E�/�����"E3\5�]Bu"O�a�7d0Ѯ\A���@v�sQ�@G{��)��xŠ��a��2i`J%�T'u!��R:|��B��=^v��S̈�v�'wa|bjŨD<@�7��(t��Uʭ��?џ'I���J�)�D����R/�(��'z m�%�:tҚ�AS囲JMN(q�')�9�0I͟p���ʍ"2���
�'F��Q@���S�µ����'-�qxCe,i���ڔ��
lȝ3�'�2Q#@�\" b@���ѕJ��y"��DUh��)�	Ή���B��y��[r��tIP*Oy���&M&�y�BѢn֒�	��`^�۲!��MS���6 ֥��!�+pZ4����"n4���ǆ7e���DFV�%� ��T����x�I �V%N@���a>X�&�y2Y�I�z��v��.� �[�AE.�y��ҡ����K��� ��6!#�yR]�7[$\+e�Fb*|�&���y"Ǉ5H��2&��)��y�����y#��UY\���I�S� �F���y2��vJ��I��]���D�� �y��ݒ@���b�	2M#��0�yb�@=g����׌�$yJ�a��yR����=��٨	�t�u���y"�\�R�v�Pw�G��du��a��yB鏫F����5�!�g�yr$�'�@sFΨ%wD@1"	��y��̷l��ٶV�����.��y�T�\]C��S>�*ٔ���y2FK5+t\T[f�	�x�d��sD�y�h޿)]��20ိB����OF��yb瀄b��@�U VK��q��S��y
� �X4�9	�mq G݋K@���"O8���C�^�]�7�N&���E"O̜�J�h���ICP�y��P"O�{���4_�H�{��ÜUl`�R"OTy�/[�z��p+^- Z�5X�"O4ʃVj�ԙ��V�(D�͛�"Oh(�æ
5  �)�J@+�����"O2IY�Bįt���Y�o�j�:�"O����ou�H`�e�^�Bg��) "OD�����<M1��E�D?z=�"O6D���S ��l�'&WB~�I��"O0������
64i9�f�=Qa�L+"O�@����s�!ghxG"O��Ё��*>�Y��#3���"O�XrQ�ؒEJ����L �D#g"O���s�,]��18@��m�"O|��0��!|`�R |���"O@U!6M��h�d`���\#"O� �ȃB�xr�&z�
��"O�=�Ua�D7 #�A�:�s5"Ozt���ȯY��I���2쨵"O����	Lz�AD��8+���0W"O��¤�� �l����|�"O��*P�ʕB�c��)z��@�"O�)�B,^�	fr���,��h��e�t"O���'�;q����Q*[�u��1C7"O,����*d<~98R(�u�\ "O�Y��Gb�����g���"O豪Bɓ���2Eh׷=h�|!�"O&��0�͠-,����L6lRd�"OT▍V�h��X ��[� z�"O�T���"�$��c�KBL����"O<��-ȉ3��1�a߳�0�["O5�2  )��1�ъ[�Ĉ@V"On`��h�.f������s���j"O��,^�L�n58�� ����d"O�9p�lШ4u� @է�[�Ԑ�d"O�}  ��
F��=+r�4j%�8qR"O�h8ԏA2R�P$ q�ޢoJ���"Ob�D�m��D�@#�.1��"Of0�0�Ä��))����!�&$��"O<���a�c�����Q�6A��"OTI����pD�h�eNG*�(l�3"OhY��ۧw��臉p��D�d"O���'�;�F�ȱ�O�77T14"O���!�� aT����'Ĕs�"OR@K�雁s�h�8��b�H+�"Oȩ�ɁcP½@Vh]���a�"O�B+��@�Ku%��]�F���"O`�c�B۬P���㊵(�@�r�"O�P@�G0aL�iP�ˉN�ܸ��"O�\�#�6W�d{1�ks��[A"O�쨔dı(�U!k���H%"O�YB&IH�^�@�@��"b��K"O6�т╧h���h�闂mpP)3"O���u�<,
ukv�ʝ!K6��"Of�2@G/09L�rͭ
lyi�"O\U�W�c���Q�"dTԫ�"O���C�ػ,#�y�C�G+9���"OX�X4�MD�$�p��� ���T"O��p���u�6����Ş p�d��"O�pa��7%!Ƒ�c���hrx�A�"O�eA�+�
\ �B�垅C:e	e"O��:7�:�D�@I\�<TRݙ�"O� �l���ͲQ�`��ӿUT�	P�"O�d�W#��(Y���u���[6�*""OИ�B�4�D��c��n*D�<���ӘF�Ƚِ��>B/| 8��9D���C�!v8�٥c�-Rb��'F#D�����M�]cx
�7V� b�>D��� Lƅy|d��#��j����A)+D�l�@�g��D�w�qx4�(@h�<�t�U;bx%���ц~��$��/�g�<iX4�tcܲi��8��%�6XΘ�ȓ��q��
Y�[���H֘��^¤@�'���sjC��Nup>���>��9 	_
%�Ʃ�3n��ȓZU̙�Q)� -)�]����"݈��pn�����X#tو�1��@:D�`����h�S�,Y�MТmc��8[����(�@�fm'�Hk��O5N��ȓ��ĸC,��~x�;��ϟ1�U��3Ô���kC=Q��cN�g��ȓ?fD��N�K� da�⇵�t�ȓ&���9�̓�E�����*��i6D��ȓ3,-r��IV��Ԙ	}���ȓ[ l]�qnՒ
�biCR(�2bԂ���_� 13KZ�Y����7{�0ԆȓgrFy��j٧k��MA�+�+V��D�ȓ$?���/�.^��t9�.Šw慅�	��E��:Zf�`�*#|ty��h��Z�A͂'�>-�T�S�lԌ�ȓ��q����|���(ռLGl���AwB��S�òK+^U�"ڬJ�T<��υ%)f� �,�%ev>��1.T�<�$+�'טxY��!Kx�0n�W�<���Nfv���B�q4d C�]Q�<quύ	J��K�$�b�m��(_O�<y���:4�vX�0ؕ~�T�9O�<�MT<�@]�1ŋ���Q��I�<�g.�$1k�e�Oi��ـ�.T��A�.׵ m܍J6%#[b�8��;D����B�H�6`	CPp�"�8D�D���A�'0 0h�F>
ψ���8D��褌�ne��xfK�r��1���6D���@�W�r=x)вT�J���'5D����70>tm�$E���#��3D�00��5=�T;�NMP�i(2�"D�`��Ch��h&���N�Np��2T���,p be��{<uy�"OfE�s/�D^j��D�!ho\9IW"Op5�  M&<� �� ��V��$"O6|���Ě}� }"�#G�	y���5"O��c�4v���Y�߆��"O�]�g�	?��P�Հ�-��<�"OB1��E�!m�@0�D,�"O����Вgb�˅�;fҤR�"O���@��Ru���^�x�"O��h�<m>���Q֙}FP=(A"Oج'���/��3�e@�J�H��"O�T�����A��@�F�@��9��"O���b�*k�&�2�3\t��"O�� H�so8�A�K��|*\q3r"O��	F���[7i@�O����"OU�ψ�<"��),Y&A�"O�e��W�ƭHAȔ�J�؃a"Oj�2ʁ+�ޅJP�F>�V�q0"Of�juG�	(e^aۗ�Q�rؼ��"O� ��z���o�0PH�F�wނ��"O���`&N�:X�5��(�^���"O�A{��(4}�؁CЭ@�|� �"OhXB���0�4̐�G�. �"O`8��HB�r����*¹G��1��"O��ӬȮN��ô/K� �R���"O�5�r"(���;q�5z�����"O�8ZA�'Va("��:4
����"O,`��t���i���+��8&"O�h�r��N�(ݘ$
S$J����"O������/��i�÷B�p�a"O��'m�h���D���}��"O�,8gHG=j�B������P���	�"O��s��	9'X���H(f���3"O䄲�i�&p!�u҆˔�G6�q��"Oޕ�"HϛM�&�Qj�;eq�Dx#"O��{3i�.4l�$NGh�"O��v
6RL6� ��� S�V"O�����P��͘���+t��}�u"O@*S�7|��H]��J�qv"O���ר�A4a*�M�3t#4C�"O\Ź� %��X�1��0u'"O��1W�W�!��D3$��*范r"O�5`��Om���Zs�'x��"OH�3���?�@H���Դ	��Y�"O��z�o��4
�O�(md�AQ�"O�@q&hªh箃�%��ax�"O��h��69ܴIҪ\H���#"O�DXE�̤}{(-;��	$���y���.@�a;���27���0e،�y�1tQА���87C�x���̥�y�#E�e���I@W!v���@W��yr
]� �"��B�  t)�u�C��y��F�
V��:!$��n� 4����yR�ЙowrܹE��d���شk���y���)�6� ��Ѩo1X�n���y¯Q�t�S��B�dTR�Ӡ���y�+��e
xY��MU�n6�W(�6�y�ME�@�V�
2��J��#���+�yrG�J)��R�
ا&i���y�hI80)�(Qc�A�!���؅���y�{&�@�r��txRZ��y��׻}��#p�Ć���krbҿ�y����+�rA	���;p�:�{�	��y2�D�NY To�vP��#�d��ybJ9d̼KbOS�q߲e@�	�yB�����ԻT�%����׭ʫ�yb�ňc�T<���|�� 7(ɷ�yB�S���x��7s���G��y�I�v�^�����>g�l1���G��y�CF��,��G�J�b�������y�%KXa�4�\Vv�4(Ԋ��y�)��Pza;�*�{�P}jc(P��y)���"�̋7Qꡛ�AX)�yR�OҮ�@-�-{>��ҲN]�<��˜M��y	@�%$&i��@�<��=���sȂ�c3$�H\X�<����`i�ɺ ��Z(���o�<��b�Z�Rh�B�nt�[��k�<y MG�|��A0%>�,�5�F_�<�'��8�f�(B�
)��xg͚U�<�+!xa�<�� Bn���x��OQ�<��-%8�8��OЃxƹ�1�Oe�<9�W�}����"[�9��BL�K�<� Ta�靴p��U����A���(V"O�りR�
V�D+Sʙ��F�)!"Of\H��Z�U��mKc	�8�Q�'9&u(�l�@��k�(7b��z�'i���G_X�lr�m^�$;�x*���M�,L�%:�E݌gg��ԫG~�(�3�ǒ \yf�i���9���w&��I��)�"u���R!���w���0|*�����Xd��ԄJqK3	�m�R�Т<%>�:��:?�J�/Ū:߄X�� �d_
�(O���d#��.xSjt �5t�p�1�^�ěB�韸c����
\�*I��N�dɢq�E*|�|I��)�'�u��Y� �lZ)klr�	��F�t٘��>��%�������E-i�������NsRlJ��J,��:��Єj	2Y�O����C@ �;JPVY!�)_��l�]�DQu)�c�~m&��|�A*^�R�h���Hi�Hc�۟�"�F����%��~B��A�k��q�M�
p`(���-��&�]W�Is>ՙv)o��%:L��@�\L�-i�b�&���2�[X���"��O|JT`�D��W���x�ā�ڠ��'S6�*���$6�x�&�O�)�Ӈ"Q�E�`G(-in����ǘ|}Rʓ���������S�Ok�����߰}�4��P���FT��*��	�7h��S�OŀA!�̄ʒ��A���!d0I�F,X��H I>��'w*N���	��x�\��(M'�ȵz�����N!8�k�O��>mJPD[����VbGGj>Հ3�5}r��*��|������5ɡǐ2a+�h[�(�27�e�VlEx���o̯.<B!ZG�ɝvߘ=:�)���~*Ѻ�(O�>�ä#V:�T�
߳2��z��c�v�"���S�PQ��{���p5�5x�LM3a] Fy��!�3�k1"3j��u8��.V�O̠	����̅91,p̺r �=��Dib�P��{t�ExZw��O�zpѤ���-���X� Ò/��%8ՊG�Mkz��DU+/.X�e�A=|θ��A�=�yra�]3�da� G+\�H��@��y��Ϙ�:��d@�*f	������yBkʅ�r�j�D�'e^�7���yBh�s�$��	C���xFmP��Py�'ٰ�&ɲb�	.eA�+�m�<u`�?e8�+�jB�n��8�g�o�<�T$��Ml�cԎ�Cr>����m�<�*Ҹ&3�<!��	�A�f\�A��m�<�ۙ?�t'	�(��jq&^�<Q�,�h��e��/��w#�[�<)���/,dAxe���d%c�Ɇp�<yQg�8hht(���	4��*�bCf�<A�o�!==�6�	t�<J-�k�<d��<@3 �����W�Eg�<�vJO�A��U�fk�(WC�w�<1��_��x��I�$Lfy(R��s�<A�W2��bg
؅i��婣��E�<qv�[�\�N��aG��hI�,�H�<����?n<��!!JBT��� %�W|�<1g��	L0@���F�@<ЄH��q�<y����td���ڸ
�r�xW�l�<A ���x��ݫNKxU��@�<B���ք��Kv� uJ�q�<�E4�f8P�Fĺ<��@��v�<	�1D}4d��#S6����fs�<1$�B�����/G��{c/�o�<���\N� ����pp�*Tk�<ɗ�K.?�~�z-'9)d�0p �{�<�q��{�4H ��炨GغC�;dVJ�x .�-sJ4iAA�,@��C��|'��#��Nc��8��
!wi�C�I&4C�ɉ�(_	X�J�9jN�txB�	4�p�D�zF��V`_ �8B�)� `�QaNgM
��_�P�H��"O �Gʅ		��ؒ�ȧE`�]�t"On=D�>r]0T�bn�-=�p�"O\l��.]�P*L�D�_27�}�V"OX�S�dE&�=�W�B&�ؒ"O<!!�eQ\���샹-�l��B"O¬ʄ�҆<�h5���
�f��Pg"Ot�cb@܋��u[1�/�ޘ)�"O2$Q-�f�"l�D��4YÃ"Oj�C%��[Ǆ��s�̚T�
�;"O���EπC�	�_�x���*�"O^Y��f�w[tK��8.���"O�paC�h�R��rɗ(��BE"O��p�.ܴ}A��ڇ��d��"O|�֌� Y�@��U6%�rqE"O��� "�=z඄�Ҡ�+\tę�"O$��$�2�@ W(�Ұ+]�!�ą��\:��`����Ç)r�P�ȓuJ���Q�n�4t��Ɍ��6$�ȓ=��qBB��
��T�Y (�I��
g�9�(8Y������I X��ȓnG�)����v�D+�C�\T�����KV�A<�`�!���H��ȓBsZE��ʛA�vi�Β?z��ȓ_�X1QQH�0��Pa�3Fq4��ȓ_�bL�WFب&��q��p����ȓ!�b�)�M3q'�<�gΙ|I^%��r�T̙��Pd�^yҢ��^M������"�[�'�V���j�e8�t��+�8���S]�d�{��I�
D�ȓô4��ڑOIB���O)0͆ȓwx<�6jۘ!���	���nG��[I���g . ;X�9��m?\݇ȓf*�l��A�H=�A"l��n8�ȓzPzJ�OO}W�Y���O'
���P��b��4l0�����P��@��u,h�a�#Y�"F��H��w �uY�����q�W����ȓ��}�a.^�R��Y�b�k,0�ȓ�B\y�$C5�u�#�g>=�ȓZ����lH�
�v�����n�TH�ȓ9Y�$:�'
�Nm�0g�?kA¤��~��6'=��tk2+�<rF�����(a�E�@t	YU,�,aNB�	.�*�0�c�
m�\`'��-w>�C䉨&fd#�ĕ@~���6�RcC䉩zUl�����0RL�pȄ�1�B��n0�H��L�;���2��j�fB�ɑ]���:��F�X�rC$�+cIC�	
{h$yh��L=	IN�2�� �B�	%q*>�����8d�@R(P���B�I�y��E:Ѯ:dr�A�\�B��Z�<y��ٍ&O�I��NU*V�I,�z�<���ѢX+�D�w|�\8���Q|�<1@�ޮR/�X1�
˅E6ѓ�Dy�<��m�Het�k&DOQ��s�Ri�<�-G���y��/ٚ*���"��a�<!�@Q:Q"����+ �^�P!VZ�<�g���n�<��3 �$F
�3$��W�<�`fɮ�Z�����h����,�R�<�!�×6�&a�5d��sh��D�LZ�<!�-��5�Խ��I�(g�V�)�`R\�<9 ˊV��KU�xo�MIp�r�<�N(�N��f޹R���sm�o�<� �pҏ7C1),ڜ(ۂ��"O��X��(u`<�7�0I���b�"O�%�3.L/t� ]t);H۸��1"O�i1���_^|�St)[�c���w"O��C�3t5N4�E*A�ƙ�d"O>X
!A�,��9rB�H�BsB�"O@��6 3X��2���Fc����"O��!V�ЗP���f���a�"O� yϴ.<`e�V��e�̐�"O��Rq%�y0l!QB�({��i"O8L��j̑a��ȣ׋>�d8�"O��p �~�|���I�*���R"O�����߰;��������;y��%"Ob@�R ��d���
,lBT�"Od��gW�}������.&
�b�"O���T,$b���!��Y
|}��"O��8�!S�O�j�"V	�X�@�"O�Qh�haic��ݭ��	k��Ӛ�y�!@"t�^�xfƽOm�6`��y��(T'�)��h
�=�h(!��y�'\�V!�V�03Pz}@�"��y�\�n���؁*���զߝ�yҧ�#������B��B튻�y��D�|�PSf!J4���X�Ց�y�Ш.� ��$�0[��Z����y�MV�#���Q�"�����/�yZ���6��L��m�v�,�р	�'��h��iضwR8�FAԼ'.p	�'��x��Ë�f�x�g4]XB��7\n�Lp0�)܎4sE���o'&B�	w5��a"�/��|Q�6�B�	�{�R͢�-�a���p�_"=�B�>?Ė�2�R�x,���B�3GNB�ɑ1�Ts��Ԉ9t���|�^B�ɪo�4a���W��Ks,�.x�nC�ɇ�Pˡ�X�u�p9����lC�I;N�L���a	6mDr8�@(A�bC�ɟ{�~��r�ŗ.�d� �I3~dC��*_M0Q�NW�)B��E�L�+H.B�	Ĉ�6*�,(^�P�P�0n�
B�I'(�V��@�)H�xɑe�ݺB�oxD�C�æ7l�x��!��>v<B�	7	P��1$
D �jp
g�y�\C�I�x��Ɂ��=$�P�!en�2_��B��! Fj�E	I�?�N01��	+[�C�I~r�Zk(*�	��9IxC�	 ��eBa��8�Т�0;��B�I[Τa�6L��@J �B䉪�f)Z�Eɛe��0�bL�]�rB�#Y�Zx��	�+<L���l��BLhB�I%��� � ]�JdS�&B�\FHB�ɪ��Y�2N��5� CC�j4B䉙(>�k j�a��IX0�Z+^�B�I���\@6�V3"��ScGK� 5�B�I�Qp0'�S,,�Q�A�+XۂB�I8X�V��1a1V;�5��N�6:�C䉌x<pAãп%��I�R'�&q+hC�Ik�����e�)$�����+]ؤC�	_�:��W❤xR ']�?��C��+#p�2�Q�n<5��`�C��!E��}I�ǖ�ENT)��/ؑ8�����!;�5�a��6�ġ9�Jؿp�!���,]]�M�b傤Y���٠g_R!�Dת>�|c��R�S�
�a�F�)VF!�� ���wh�pg,x�&��rN���E"O���O� =ZdxG%�zH(%Z"OR-B��SaZ� �.^hԠ�"O��F��v.($·:���{7"O����n�7 �.�k��K�P}��"OBp1��N/R�����r*���"O<hY��Pp��$r$�UU����"O�u� �RX�1�Wiθ"BAFx�<"���f�vq# Glt��"�r�<��bG2�\|C�(ކ>,a�b@E�<�I�nJ*��fN�h���"S/�D�<	�Ɨ/p��fY�P�!�BLD�<Q�N�9\t2����@���I�<��H��mO�C�f�j�<YԮ��p1f���g�V8�ڠ��j�<��#� ^Di���K�i.�	�	�i�<�W�*�L|qlS"4<�c�|�<q�K��aJd��r�`��D
{�<��ڨ!N<0���%M&N �ed�k�<��gE(h�Pu�r/R�xft9w�g�<&AK)#��y8S�Y�r+n���`�<�'&0P�שC�Id<P+G^�<A��õ,�XQ���>A�H���W�<�rhYg$� ���6 ����s�S�<Q��,r��if)�;E�䚥�d�<a��[	j�2x�7�M�M�R�Zgɐ[�<�4��%��Å��1}f�����S�<ɢ�'1"�P�� �ހ�b5ePT�<!��"J����"�*4]BL7�GU�<��m��wH!�
R��Fa{m\T�<Y##)�p�(�G��XF����JF�<9wd��NXE�Q!OB���gAK}�<i�dY�!���s&	�0��Y�Wv�<� �	&]��z�茷@|"A�e��m�<���� 0  ��     �  z  \   -+  e6  	?  0J  7V  {\  �b  *i  jo  �u  �{  0�  t�  ��  ��  <�  �  ��  �  C�  ��  ��  ��  *�  l�  ��  ��  A�  ��  ��  H�  � �	 �  Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�� |d��"O
`�(�;���8���-0��1%"Oj4��ND^[��"3/9�0|H�"OB���H��*�ʞRy=a"O�味V�!X��!&F�:J�$���"O,��a
���C�Ą�M�"O,$3%o�-���p���+Ն�:1"O��ݢ1����`���y14]2��i�<�6��{_���c�H�`�fX�$Kn�<��A̼VI�xR[�)�Ć�pඤ�ȓA5��('nߡ4�� �)˩%� ���,��r�؊b#`T�eT09���ȓ!�b��g��}�8�F��-? �ȓ
K|m�ș�VṔ���2�%�ȓ"R�X�j�4JN�1�˘X�i����̹	_�jZ��1!g��zܶ��ȓgil,*�J�
j�Ne��i�J%b���f	�(U��:���G��$Y^م�~r�� S�%T"���k\�jx�ȓ|4�1�îJb��@ӵ�ݩn�V��/[`�"�v4�R�!ʎ<��M�ȓ`:��z�ؚh�J�Z��$HY:	��H��p�m�C1��!��B:��0��EnjZA V;9����J[
2���	��4'J�EA�IVW&��~�(aZ��ӹ�>� o�Y�|�ȓ�f�A�
Ο7�H��M�$�����mޠP����/���ANXo*�ȓTv�����{ ��-7�*h��I��sB�8�8���3����ȓNe*M�悡;������X�o��!�ȓ'lj�#F�m�+R&;�|��2)n�C��0S4���T:
b���:�0!��e֊��)��ͷV��,�ȓ0�&�8#���� ع�L���mL�����&m,B	Ġ�C��
�l���$�/�y�ƕ,v�FAj=	ݶ�2g���~�'Irqˠ��lh�Ӱ�Z7	S�'
h�)֠�	z�	G�;lta�'#@��a��~��p�FB�66�N>a	�X�L�(���^H���vNU:2�h5��uK�x�1K��{#�d�b � ^�
�B���s��� ��*zz�!e O!kY�áD5D�Ъ�╭U��9��AQ2{���(�On�6���Z/Y���MK�����GԽ�!'����u!H���T��Id�'�$*ס!���-^	vsl1��O�ץl�$c�"}�UG�R"ȼ�2%��s�$APR��hO�O9H(bM�]�A��@�O�ujI<q��'Faz�H߲���*�Ցp ��1��?!�'��a��;�
��7�2�R�!�'���s�N3x�܀J�(��;^h){�'N�d�M�5a\��KvK��ae�9��(O���f��
�y�-�\�B1"Oj�"��CF�cU�}k6�Y "Ov��t̞,\���SW�N�~�����"Oz�3��X V ��q��U�t^���'⑞�yqNڲ|�ع���C��51f�6D��;���`�T����#'�eH��3D����l�.>�ec1�S��3D��{JJ�%�\hÂ @�0a�,?D�����&�R��D�K7����bE8D�� ��C�.@�C�a��$�&Q�*�g"O��ऊ�%�vh Đ&t¬HcS"O� aA�77�(]�"��	��)�%"O���PAM�8wpـ$�]�5��m�a"O-)���U��;vdq
�L�%r�!��;w�R	��>l�v���o|!�Z�Cq
��%��9�>�l�9Le�b<O�ěU�_:R���D��V��z�$5|O>�y���%'�Q`#JJ�a���E{���>
�<��JI�P*6�3��8�!�$��mcҴ��@3.(P���O�;m�!�DO)T�zg�Y�jb�rg���.�!� 7Ā�b��3�6���L���!��2p^��rk zB�$�S0�az��������W �����*�5N�!�8�\yre�'<��8�R*֋X�qO����<���١^+��Qt�@?�ܹ�� |!�DE%)�0m�#�܀mDP��4)EGbTX�'a���s��"}�'�z���@3	���)GA	�y���	6Lٓ��E�xf0�נ�<9��6�Y�J�Z���}�g�'fƜZ� �2hFa')�$�y����dO�e��I{ �I�o�D�わ��L����b� ��$" ?xt�@ɀ��J�Exr�x�  o��c����F�}:���nZ5Hx�P���.D���6��7:��w�>$l��a!��!�HO�O�D`��'<�f���*�`F=�
�'LB�Y����8zΩS���Z�	�'�R���C�uY�'З�R�:�'0|,XF�6=r��V�B�1����4�PxB�.;�Yb4��eP�]���C�y���(.�<((B�Z�Z<Xq��y2G$�-�B�A��|k7���'oў�OgFTa�T�9�[�c�y��'H M"S@S�� �#DD�����$6O�y	b�	�8������axHۅ"O���D��D2z��%rG  "O\C��q��X!�S�Fn���'e�Oj���bo�v!eʵ:x5�q"O�Eˤ��.U;��_.P3�1��d�H���'F/ڸ�T����� �/Q�>����oy��ғ8b�%I��D$��8�G�]��y��1�F �"$�|Ya�����xR��>>kh�K{a��
$�\Ÿe`(D��J2e�g�$����>S�xpF�$��=�Idz�__yC�-�� �D�U4��a�	8�y2h��EQ�h�D��r`����u�B"=	��4�J a��5}L��r��</�eq�O�a�6*�9��p�s� h<�B�'�����D�S�O���g��2�L��ۋ�`��O��=E��eҒ2��)�Ɂ=�4�J	��'��{b�� ,�DE�<��������?1,O��O?���J�K�@zӈ [�����"HY�<�g�	YOR��'_�?8��m�T�<� !�MPVq��D;eY48(EhJRX��O�]#2cǊ���.K,X�h��"O�$�f`[!��H�&�E 'DT��"O�x[�+^-:�ĵ2�āC���d"O�%	#��W1Z=is�Y�M�Œ�"Od��	[�G�(���n��$��"O>Q��	�+i|���&�*�t)ڧ�e~�i�ў�����G)P0k�z�Z�0a���D�'Tb�`[��I�V�h�D	�!Ix��WO&D�d�RI[�ϖ8��?d*9�De#��\W��ħ�Mc&&5w"T������S�d�~�<� >�� N@��0�T�_�b{�}��$V�Ø'=P�i��L�1!���`�Vء�'�Lɀ����?��d ��:��eQb�$4��x�/ߨUN ���ܧTE���4�O�5�̤X���d�*�B�E�`T~}�?I��0< �k��ش�G�K/�}c�f���"�'}���G�I00h����6E|�a���s�ܐq���EC2�T
 �4��q�-,Ol�<S�fx1��B��l����ӟpx��|��l��.ϵk��*�!�)�I��'"b}����=�`ؖoW�7�p���(OHC0Q�-�0���5d^f}�c���b���o�J�Mգ^��9����Z�r��ȓ�6���Œ~��٠ǝ�*���EzR�'I(1�1	;�r���@&�i�+Ot�=E��^�D�f����"�tb�y2d9G��lRc�[o��$ ���y��15v�3�ިt���fB��y"#�j����ߢ]M
0Q�C�yB��w��M3C�$��x��K]?�yB��1E�r�����U  a�y�JGcҁ�L� �2a9�Q�y�

T����b���\ɢg�6�y�Xwp�0ɀ�n��R�y��L��A�a��LyP!U?ШO��@#�S�"����R-R�v��5`���<4C䉎�25IeK���a;����|��ʓm��<E�䌁#	^��Xs���_� ������y��[�G��P%A�C�y2�:�y�M��!�l����\7��Д�yҋ[?�]y�iW:)�ʥ���7�y�톶'b=��\�@� �@�@��y��V�s��4���\�k����yr�̀wp|�J��S78-j�*����y��@��l/,�3��7lDxy�'6`��ff�/:�ⅺ�/Ʋ]�
�'�aE�an6��Eg.|��
�'׸\�����~�+����]݈�h	�'U�A���]!I� &IT�U��z�']d�`&��,,�E�� G�X`�'haj���'?��1��B�c����'����Z��ad���^C���'�����t�����,Ԑ}B�'�Vd��N�>
$P+em��(���q�'�4���Ì��F���H+"�
�'�f�B�ۄ஄������!��'�3ЌA3��2%���m�'%̰��UGY~x����yD\<�'i�y��C��O1T��N�HG�tz�'�$Q�łX�4�����
�'��qH���r�.�+�D��z�#�'X>��6A� Z�� Q
|�
�'Z�X��\�JD����y�A�	�'!�@6�IU����$�wb9�'�|�U�I�x��W��
E� ��
�'t�$"�"۫`�|+7D��@e��y
�'$������QA�j��Ϥ-w�I�	�'��r �ޭz�؍��-]p� ;�'l�ɂN.����Y�*���
�'���swh�PَH�b��	4��5�
�'
r�B4�4'2��Q�`f��
�'|^X�ueF�tZ4�N�/c>ԁ
�'�HY���C��R`�2ě.F���)�'��a C"M�싂�9��0��� �娡 >F5	$X&L�T��"On���Y�}�@��E	*%~h�"O������n� �k分��M�1"O�@j�A�s۬ea6�
c.���"O�sA�P���ʱ�X�)��	���'b��'B�'�b�'���'���'�0Ȑ� sϜA:A��4�N�+��'6��'R�'��'���'�2�'jvZ!�c�P�B"عL��A`��'B�'b��'1B�'jr�'���'K���A9�Ȃ�E��q�F͐4�'�b�'W��'���'h�'���'�������"%|4��r�5��h	��'��'���'$��'_"�'���'��,��N�a�q��њ@�v�96�'�r�'��'�'�r�'���'�bs�d �3�����~����'A��'ab�'j�'���'�2�'�$��:�ޙ���[�_�r��E�'=��'��'S��'���'���'3�S��+�P�TMW�N�09���'W2�'.B�'�"�'h2�'�R�'Yd����U�bd�� C� ��[�'���'+��'WB�'rb�'���'��[�!�p�@B�n��$F�'nb�'��'c��'="�'���'`� �cP���i��O>I�J5�u�' ��'b����T�'���'���'.�+T��%��eBS�H�{��c��'j��'.�'���'*��h�j���OPe��`�%i���DZ�V���gJfy��'�)�3?�ոi6�(Z�C�<[r��%ȇz��a������ԦE�?��<1��1jF%PI+4�Puz�G9G�ļ���?�o��`}x�'3�[�?���0$y'gKb�-+&��/X�����O���h��5�@�A�`I�5�p�p~����̦�h��)��v��j���w�����$
�H���8���U�'�0O:�S�'9�&�Q�W�<��c	�6(p�H�k��}����<q�'�&����hO��O�r1k��D�:��a���
�24��2O����n�֪���'ݜ��#�=�^�85��T0���I}��'�B2OH�C��\���܌~(M�%�$�i�'�"��]��	�$�Bß�q�'�������S�P8n�
X ��P� �'!��9OHͻQ.٦ehP7LF3a�
L/�yb�t�fh�v�� �ܴ������O.2!�|I�G�N	�)�ϖ$�y�'��'�����O.��b>՚�'\d,�S�l��K��!#a���!U�(`/̠� p2�͐�$ꎨ������\Z��,e�dI��m��5}@8h�-ˮ���r) 5H�.� ̨u�(P�aѓߌH��� La|"�F�X��������M0B,���z��Պ���MCa��-ؚ�j�(��H��a��	�9
���p�.���
8)T�H�x�TP��Hɀ.}��:#�̃_�p�l�:��x�$�8S{�陰�����a����-u�x��D���"(�ͨ\�t����f�P[1�2�:T{�nX�v*�Q�@@�w ���'�R�'��t�Om�ݚ����ƑT����3���M@��?� ��?�(O�$�e5����O����4z��eCF�@0r�V'��-�Hvioҟ���|���?%�	������i�V�a��4G_��U4z�ɘ�4��t���?�.O�i:�i�O�0��"��kL1x��
b3z`�b�ZѦ9��런�I�y%V�0ڴ�?����?����?��
�>LfN��v���8v��lZƟĕ'A������I�O����O<L�L�*�uj`	[�:_��L�Ȧ���({y6�Pٴ�?����?�*��@?Y�#Y����cÔx:�����K}�F��y��'m�'G��'���'�� �n��T�T����K�|�b$����v`6��O���O��D L�D_����f�*�*)�Z���E%
Ę@��p���I�I��(�Iɟ��I�?����4C%(L�W��52Rv4���Q���jC�i��'�"�'l_���	�M��瓼Z�n5kđ~3ZHp�'ũx��ɰ�4�?����?A��V��KG@�k�4�?����bM`Q��@ nI��iĄG�`��iM�'UW�0��`~4P�'m�$R�TL�@�b�1y8h2r���*���'f��'G$H9�6-�OJ���O��)�t��B�/�&\T���M�8I�]l�����'sR�؍����'m�i>7���A>Z�ڠ+�*Ev1(���&��&�'�ų �~7m�O�D�O������%�L����U^���@������'�BC��.,"�|�O,�'a�|0Xf��i]͛�エk 6]nڒ3�6�C�4�?����?9������?������aM�f��$��c��Z׷i���Y��'�ɧ����$�'�> ����a
�@=b��iz�MlӾ�d�Or�/w�H�m�ן��	쟄�	͟�ݢ&h<Ia��A�A�G�].`6-�O��Ǟ7���W>O���?��ǟ��ԍV����Z!ů@\ a�Ǒ
�MK��H�ʐ�ݦ�	����	��\��F�	>� ��pK��&����ve X�*6mƛ�n�34O��$�O��I�O���|�o9��#pǜ��U� =� ��!�"�Mk��?I���?�[?��'��p�R�ĆX5"u)H`�LEB�x�O����O����O����OT��S��ȦEJ�c��q��I��@Z�ؓ�kM�M��?���?������Oءr�7����L�Z�H$J����I���צ��Iǟ������ٟ�׫S��Mc��?q����= |ҁ	�iW��3e��=Y���'*"�'Y��Ɵ��(e>}�	K?�`��(ff�(p��C$���0WA�̦q��ݟ|�'���Ya4�	�O����(Uy�� ��)��� �f́X� '���'�~U#��T?� |�ӳ� V�j�Z�l�V�`aC��i{�m&Di�4;���럸�S&��D	�Y�<�K�ҫ�r�6���~��&[�d+�;�S�NV������*HX�p2�	�1���n�eZ��Cݴ�?����?!�'��'�B�F�<�`���8Nh��Jm�67M��"|���}�5���&	�!9a��DМHrp�i>2�'%B��O��OL���O��ɢo�Ա��+#H(��g� ��b�k��'�I������N� �0��; f;�i�(�M�����	#D�x��'�B�|Zc^p���Z;:;�͋�g��$-6塬O���#�$�O����O��H��H���_��B�'�!��b@\�@>�'A��'��'@�ɧR� 27j�pE��2�<���5o5�����I�ԕ'>����$w>%qҀ��UK9�\�7%6���?)M>�.O�䀂_��1�&^=Fi�\�"*E.x����H�>i���?����ԧX_��$>���="�ȸ�*Y�(���«�M���������O(���KW8baj�?3�.т³i�R�'-�	-`�Q�I|���c�\Y�L�o�Dj\��
��H��'.�	�2#<�O!(��d*C�:$J���R�aܴ��dL��,�n���i�O^��[i~Ba�,J'Da1�'�	Z�i�S�O6�M�-O애V�)���>*�H��C�(��q ���QC�6�Z+d<pl��	П`������?�PIK&6�Ƚ�ѥĶkٚ�*V 	�(O��(@��O>1�IaŰ��	B�4�����N�bL��4�?���?����m<�O �d��lhƝ6I޽+cB[� IZ=1"i%�I� �6b����џ8�	w�ސ CUJ905퓌���ݴ�?ဧ� c��O8��<�����DĻ9�P�b������`�Y�ع�"�ß��I�|�	̟��	C���S	\W:uz�O�7	�TC�գu	���3�I���&��'��p����#L%�wi^�%�1�J̙��'8B�'��T�d�a����E�9��U���9qp� 3����ē�?	I>�*O|q�qU�L`F熕���90��"ؔ zB;>����?	����D��
��'>ٹ1lm���Iխڈs�b�Ёƈ*�M���?)OV�&�����䀧v�r!��n��]ݞ�(Vڳ*|�V�'��[��rfR�ħ�?Y��f���1���_b$ Q�Ζ�v�,��#�i���By�������sӼ���,A82�6��� [hQ�آa�i�4m��@��4;v�؟�����d�09:���e�t-s�#O�Ce�6W������s��|&�h���n�qȃM_2��` �k���{������̟L���?��N<���O.b�N�4r$�+��)@"P}���i�(���4�1O�� �^<�Ҕ�һW,4�HC�߈Y�mn��X�IƟ�G���ē�?��~��5M�^L�L�Ѱ�8#�]%��'���=��?)���MC&̐�?U��c*��E*��#{ӂ�$*sq��%��I�8%���m������C)>=�ړ!�l>v�]و�<���?�����)��d���R�``#`�Ӎ9T�a��K�v�I���b�	fyB��zuJ��K~�� �D�j~b=@�y��'=B�'?�{��Y��OhԬzT�� ˲�D�Q&�E�O�D�Or�OʓHϢ��'Y,��d�T9��Z�Á1`R�Q:�O����O����<��OΒ h�Om8e�$�@(x� �!l���na�S�`�$�;���<ɲ �e�<�n��e��.%8��mҭH��o�����IGyr �d_��$�d��.�/PДS���O����ꐅt��'���'�VUэ�T?q R�ܭ3�Æ@��*(QUjv�ʓ:��xc�i�f맍?I��S�I�>�ȕr4_�v��a��Y>l7�<��J���O8ir�ʶ�y!A [�_��Y�4�"hQA�iB�'ab�O�.O���L�Ne��&o�z�EX�FEM�ƅn�e8�#<E��'�p�զ]��y$	�B�a�"�pӆ���O �A[T&�L�	�(��
E� ���BIGx��wK��yM&4�>�W��?����?���?i�! p�"�,�LKp'�g/L|��iTB�d��O����OOk�ڲK�"�̒"4̔h3&b�$�I�Q��c���Iӟ���qy��� P)��{����n�eǃ�OJ�iN9��O��$8���<�p)B�^h��
�U�N��򑁀0\�L��<���?1���D�?1Ϡ��'a@h��1o�Be<�+U�|��'��'-�'�I�h�)%0, Ŏ�T*�횆�ݶt%�Y�'5��'�b]�X���ħn��G��h���c]�7dm�D�i��'Z�I�L�����g}2� �Bt��' ����@3�fF��M��?Y+O��
� �a���x��Bb��#�EР@䰤)�W�F���ش���O����0��3?��]@���>r���0�e���<`(d%e�|�4�p� ѱiKR�'�?��'l��%c��Y(���w-�'�6m�OV�/XӬ��3��-u��	�KN>;1���o�>�րQ�5�z7-�Ol���O2�i�o�<u���ŏ�)�}�dH�?u�<{��iZ�т��4�1OX�$�? �
�ܩf!����A�u��}Y�i��'��*)�DO*���O���O�UlR�bE`�#T�v��@N"5f��>qe�B̓�?����?AE˜;f8x��G	 H�`(:d"z���'�$�h�5�����%��X];�y �*j��5�@��U���P����<����?������^�^�B�/�'5�%��π9H���FɎ`����X��Y���\�	�oȶU��V�M��� ��"8�eSV�r���'���'!V����Z�����(���`q�&
��h�ꓛ?�����?��S��\j�PF�YbR(��<�2�܂3��k#U�|��ٟ,�	[ybma���ԅ��[(�90�G7i�F@e�Φ���D�����	3f��IH�	 |��s�ҳK�� DA�u$���'NbY��8"��ħ�?q�'t�� gv�ʗl� d? l �@���?���,�1(���䓂�dʘ/Zzd�;ǃ �c1�-�n@�M�-Oj��b̅�������$�E�'+D��D���B�݁Y�@Zܴ�?���L�Ia�)�S�>�)���M֠�A���)V7�"6lz�m�����˟l�S���?ѱn
�'_���p�谉����p�֭���y"�|���O�|�ay� e����Y�<ݑ �ߦ1�I��p����`�K<����?A�'l.�JGK+�<�b�,�<<�%�۴��"#2�Cp��t�'�'��	)6�4=v9��=k�Hh�`�m�d�$��*Hx�>������uc�"&��|xE*� +xQ�2F�T}݇�y�[�����(��ny�O^3l6�@&J6ҭ�4.����YC	#�����'"�'���Ȁ#��Y[��ϐɞ)���(�F}�'��	ݟ����d�'�D�t>�����:.^4�`����R�n�>����?YO>���?Y��@*�?��k�5�؁t�#>̴��b�FD���������4�'��	D�9�i�)����d�I��Zu���&|oϟH�'�R�'=��[�V�Z�֝�_>���5�_9�q8�(�9ˤ7�O6�$�<�u�,kh�O���O.ֈ#E��8L��jW��ql�-��9��O���I���d)���?�����dۈ<���k�,Q2)��R�I� |T)c�FH���g�]���jOk)Pt��E�)�'/>u�#
�68�4�٤�W�g��Ab�;�p(����G�@���@��0~����?+��I�%�R�s9�Y��a�'�W�� d
���#�zI\̻���K�f��� Ra)
�AWEǹq}������6<Z5�W!�na,,C	V�� s�bQ.Fd�1gF�%�D욕��9c���CV=B-�A!2�'��'-gp���	�L*�f�/kp�|� '# ��r�F?8��gq~�3���DH��S�	�����;-Wf��!Ԍ�#�����cƭI:��	�� �.��q"ݟ��ۂ���O�lJt,ѣZ ��Q�Ո6r��C�O�"�':2�'x�O�ʧ��	��ᇉz��	�d�N�|��|�T81&ӋH�9�o$s���9`�i>��IryBa#��6���i�.\����;:��g��$K����O���O�t#��O`��t>��$%�,E�4��GL�{��He� H�|�����X��E�$a�Tx���S��o�@ݘ��9~�a�7�Q�k�Z��%����r!�?y�^��i�&j���?�t�韬�ɂ<��!J�6[¼�3#P	T���D{��� �`7�	�	��C���' �C�.PTIx���5Ǣ`�[	|72�I;�M������ы���m�� �IE�Ԩ�$E.�xŷZĈ˖�9u)P�#d�'��'��%"���u`.-��,$T
�T>A�)kv���J�#_���&6ʓJ}�����4ku��2lL��ħ&��	��(&B@y��[9J���Dy2�܏�?����?q����>uh��'��2^4��#s�ʸk���2�)��<1��]�H8��)(
��تPm�U�,KK<!w,��7aFR�F�8~�ڠ&X�<t��"��E/�?Y�����.���D�O�d4#�6X3a���<��Ʀ9N&q:���,����/N�XL� �Co�D��wd�=��b��U/�1�V�^�|�8B&��I\XPwe��0�����,�r�}�]0|��!
�c�L�H ���Vk���(������4S0�6�'�?�Y�sL������xd3��_��d�OH����D��|��D��5�* �.�����㟺�$�	dzx�偂s�(��0ꁭn�T�$�O8�����	7��d�O����O��;�?��N�l͸���Yz���UN!B.6d�E��|iT�u�M����g��jڠJ�5�b�تDa��8I ��lġ0�H��c"�%jf����$�R�BүؔC�����eYu�TK�ɭ~��ّ�CQ��9��m��	�5��d[ɦ��N<1��?y,O�  �n̏���3bb��C@ΰR"O�=˒lɁ9�Z�҅��;;=v({G%L�'����'��Iu
 s��
�T�I*���r]��8�$٫�?)��?���4t����?�O%���Z�8��0#&S�n�b���}��T$�� 걘�'�������g��1Ś,�:(�eH�!O�Rt�SIޔ10tݰ��'�Tt����?qF�s�Z�c�L�U޶	Y"����?!���s��q�"j{n�3.�.4�S�'D�� <� ��=O(D3�ʹs�*q�d3O�%lZş �'��q�a�&���O\˧L�x(���$�l *��A����@��?!���?�d��/d�!䙨���j���}�����{.�`)ނ��(Q��u9�<iń��
3䥫c閟9Һ,BD_�B^��	�7�ly�t�˳q_�1�7O���Q��x���O��� �	�Oj�! ��D��BF�!�-�g��O��"~Γ3�lUb�2U��m�����c�)��I��ēe��0����"��Ժ�	C(B��ϓ+��S�iV��'��uvm���I79���r@�T	}�=r�?~[�5�N51�-��ש2p�%�P)�2UKC,I���Y�d��7��Q�GH7;��<ː䜕ge�BKfZԺ0���*  �@���%�,�yN~��3���0��\�X��+�q�m	��ȟ��ݴJ��)����ʓgx���3Թ��FBu���P�(-2AP��FtqB��u�ƬFxB�-ғu���'ELz�nR�
����ǑrA<��'�R@��-���X��'-��'�g��	ȟ�C`�:�!���m�(��b)����b�,�|hb���IX�X ��ތXǜ�H��:/Bay�p�0�$��0$��хٍN��S?Q���C�ŖU�Z�B�ڑC.���Q����B�J�O�n��ē�?����\�P�\�ȁo^7�"�p�R�c!��'��3�N��!��z��݆-���Ezʟ˓S�(��iޘ�a���nz�y$eJ�pN)"�'Tb�'BBM>E���'6�	@ :�laC�G ���Bk�7����܅7\ �fI��ÆBd=��Z����=o��H���֡�@,$GP�E�0�r���Zy����M
��OiÐ�'�l7�#Y 8�C+*z�()��f̡oS<5n�ğ8�'{2��?�x7헣[�F�C!�?|j�����%D��(��j�����i�p8ԣb�T[��џ��'�R<QMe�	��ş�Ox.Az�cV$G|6��b���F�H�`@m��1�'�M?�l��E=q6EP1gʠ|��8a JG�'�L����>Wp@�[�A� =��dڎ��T��u�&�'a@L���ܯ�g��IS�O)]���r��-	5ҰS6�+ʓea���I۟�'?���%��#�g�04���T��#L͒��Ip�S��y�o�a�8(���pd�Q!T��0>٤�x�ϴݰ�`�G�g9B!��������Op��,<OR�zV��X�PH뢬�3)�f8�a"O���#�ɽ���՜Gs�[&"O�+�C��.8Ѕ�ӴT�p|��"O��ǅ��%&�(�s)KGD��"O0���
�b�����9KN��`�"O����9a �u��'U�>t���"O����	^5!F`[�E�7�Ha��"O�̓2��sT�Q�!#&�`�J0"Oj5�Ӊ�$>����8*hD2W"Op�kB�[(�N��!��0�	��"O�;!S/�}J��b�M��"O|����J���k�&CX����"O��� �K�:���O�%�0��"O��"I��ykx�qdNآKBH�"O��Jg�9#DI��Ңj#sv"O����ɿ[4e�#E�����"O�	e���D=�P �D�n�C1"Ox�zŢ�"��� !F--bj�"O� YThI6Xe2a�BL%@lԥb"O�$��'U�s�v�+��|�"O`푠׹F*QU��	y�͐@"OVh�q���I;����@�op|�b"O��p-�$<|q�'��
Z�Ȱ"OB��N��O�S!n '��xb"O`4�t�[�|���+�ڽK�"O*�����7eT����iC\�*���"OYhu Q8?�l�Є�ȝ!���p"O��"hJ;vs���Fe�_�pZ�"O�H퓽�$j�M(2�䱺�"O.TK�!OI����ݘ���(�"O�ӣ,Y�c��	궧S9e�|���"O�D�U凋.�z$�\�B��j�E�Q헫nFz%�,�T>㞈��#Wrg2pH`R�/��)R���y�rT#s.�D� ��f���OD�Nנ?�4D9f��o�� eK�|�g_(������ �0A`��C�	��F�Gb<�4�!ӨO��8�#� (��9r �S0�G�̜@�p�q,ޕm���	��?pxqO�a��/�����y�����"_\ԉ��g�h����*?���+KN,�B�ω�b�4#R�k��?���!V�6��(U	obEk��>��'1�4Xd��"�3����7���'�=}2�hh6��v�ӕ�*e��Jc�n�.�8\��{���'.�ᆇX1V�`#�����J�>.���gp���E��~ԧyW�:��L���W)N��JFʦ��ɏpҜ5�?����3o�pt��/V�Ӕ�)N�#?����(h(|�����4L��I������5,)���c㚜A� ��uE�@̓T����H�^�	�&ٴY� 蛃C�b�ʩS����4E��Q��#}�g.���"o�2թ^��Hx�Ox� �&b�M;�cry����7zDaÄ�|�"�A� �&O�5>7��q�퍥T�����!rt\�w�ԟ�O<�R�k�(x�$���7lD�T��S%:���sC��N��y�B�_U�y�c�M`�:Z�:�S&�4he�O�u��D.�)��&�b$s%�5_2��
����s��=cv�I2q�b\�!�ډP��8����b�	�S�ck�,bU��v
�͠�(�	E}f��=��ݟ���g�pH����F9�hQ� =
fP�'rAӦ�,:�͢��.	<\���{�'I��Q��
E�K/C*��.�3O�qO�HY��i�5k'�J6^!�q��gXE�dCAW������1Kh\IS)H2e�65p-/�����ԟ�O�Td�4j0�h��P�3��-�6!^ �L���M= �8�����O�n�R�B��j�[F�!�hǳ��@����G���B�4�`��R��:�Q�
ɳT�*�J��ď�R4�R�A��Ȟ�@��)��UR�]6Ҝ9�!��LN��{�OH�1O���O���`Ra��R�.m ��طL���@ĉ��J��O`D��Q���T"ɅMD���|�'pxF"���>���+�
	{$���|�;�ݬ��d뷎_�%eʒO�ٳ��G)8*ҵ2��ˊV{�8�+��|���*MC&���!��&7(��c�;zzD����^%f��Pr��Q�����OT�Y�T`���56�NBrp�pɐ�h����
��}�8�J1�|�Y>�'�XsȃX%�E�S(��b���'0J���P+E�S�C����p�Ӯ0��8�􉂩q!^�������6ǀ�O�L�	�B��<9�'�<|l�?) �oө;�{�nU>���'��LU�p�􄕫]G��Y��GRx���C�n���
yV�ɱj�[E�(���)�6����'+�Ql��z�>�dCȺ[�/7�;�x���ɭ@�xXqU!SQ�`l/[�01��'���(`"�4H�R�ԟxY��h�0��ˆ�w��\Q�jí?x��˂
�9�27mȹkjRl�	�I��8R�i�U�Ь)�bї(v2ə �A�ݺ(|�4�(�0E���B�{��]�!jv<0���y��
R���'����1���ٴ]-J�yT��&pS���1�О�VH��'�$��2�i��;�`�OJ�{P��4ۆ��5ݟ$�i�7�lx�J���u�7B��z�)GzbE�;+�6�C��߬6R:��HT"�?�SM�
R#��X��pBp���{.|���`�R��a@D�(����w�53S�	0�j���*���y �[�]��קV/"�I�B�G��d�AV��3��9���tGļ'wRP����������X��D�yv/5�O�P9,U�^2���CN�p1>Y�bcuyR�x��O1��҅�3L����N�!&��b�GGѰ=�4̔>���&��w�m��)P�v�01zv+�Ym��4�'��l���ɍ`�f��Oø$�hm���D�{e�D+P�N�}NY+�o�\�V��!�RR��P�z�8'��e��a�:��Re� 7E��dn;}��ڴA�%[3�̖b8�P2dF��'�0�`%�W?R�ƀ����gQlXh�*b|�!�b-�z�6,O�}r��U�-d@���uO�qxD��W�^��F.����ʅ^h$���Q�FKr�C�9Gɪ]��Ʌ�z�ƭ���Ё�"��S30���'lOV�pub�Qu���K�&��K����5���DkC����T\������d�+Ƙ��L�ic��^�f��P���@�1��3��'�L ���=^$z ���R42"�I<a$��S�
�c��t�t���#�M��8Xi���W�[$�AuM�<��OXL.��,@���_����̜�&���"T~����>���X-?��pb ֔3D���O�����F0`L;�H$|O*5Qe���$0�\��BЫ^�����Bsyr�+/�O1������%}i�I�d�0Ua!����;��=Q� �o������=��3&G��(d��#�Z����{��7���,\})���So�7��#Fhx�Dk�p��UbĮ�J�a��'���V�Ԩ�;q,Z��	:z�|����$l��#ߦ6��6m�/�|Y����Cx��ϓ|��A���Yd�R-2�o�d_��&��X`��MH�9둧E���'��:��	��L�[%h0Peh�
\�*��']���Ui��,����Ǟ9J���:������;<*�S�$�i�E��
�ܠd��PN���aQ8$�d�� �p�����!���	\X�ØG�Z@����8�Z�_F�9 �
B�����Ӓ|"�C<:h���ɍD����7`Ȱ<9��+WH��j�c�>HP�D9�������*N�p���^|�F��:x�=@WMЩWn���Iz�l�Eև�����-wf���Ѧ�`|ڴ́^:�qa�W1�m��MND��������T ���FL4kJ"p{��~�N$2лX��E�
�]���u&+VB,ѭفt�����)�x'b0�`-ԒQI��@?��O��I�,�lqP���&c<n�� �F-&p\u�'�d����K!���F��v�6�G�+�����֤�x-��l�K#�����/@J��'F�riM� �ݙP�E��i�%J9�����Bܝ��#�t�7�|�
6�I�������32��)2���@d�ïD4e��-	�y�$Ml���v�9�A�$tXN�k��\:����?���D2p���B��(4��;��K�{�N%�\�A�L �W�,T���\@�A��t���9�[?�A��
:%(���ߛ+R�s��@ Z����W���Q�����	�t4���1h7���;����,(~ ���8�v�p1	�o}�IZ��MKG�ٶ�\� ���>�����N�_-4���C�p{��K񣕦��s��)�xQ4�І��݈��"�@�Р
�aÎm���Н��D$KB��MG�{1��R��(Q,α҆.�5�6�_�q9�!��}iL� ��:�B�L`V�2D��V��$�l4t�#�^p��� �ECb�V��զIg~B���pDr����]��D���	���'	��!�*Ev�(7���ya�l�(��o�"|�Vl�3Jɚ*�qɒ��-�7J�v�*3���9���e�x�ꖋ�#,2���biT)��[��G�.9�=�&��/��=!�+	�|�Q�A`���Ͱ3��-2zP��#59���څE�3�#����]��JF��hg�!���%��=�.�qQ�{R�ϣo"������PD�#dLX���
��T�t	2G�*t=CĀ�.]ﰈH�D�@}��	F�t�x�ݟ�����Z!c��(K��b�8�!�[����GzRǎ�ǔ���FY�*�L�ᄡN3/5l�Ӑ-�¡@]���5�BO~��\��T�	
��0m#��gݵ�V�	�e����vE�z�-��gO�V��7�=X^��aݴ,K���U�� �ߟ�eYЋ߾
-V`A��B�|��t"m�;G���K\�B�獞< ���V� v�s��
PF���ؚ9���
tmW;, m�k�
���F�`�v�q���?��ɪYz��N$hy�b��B���Y��śha}�
W�wQa���xPj��v�� �2�Q�2��6:bM8���*6TF1hP�'�p�!Ҍ8-��4���s��i�~Ti׀֦!����>J��Gz�%�8����ɰ%����i/�?��*��y'��'o�t�2��ͅCT)���i`��e�F�d��?���L�d�z��e�1S3 ���?z��4Kҡ+V�m�@��|������N�6M�aZ8Hq�A{E�Ą{4�ɀl�4z�������NM����Ď<,���ʑ�B9���"�e���?r%sO>	(��k��c5��}QZPQ�����
�6��DkEMU;�j�9���n��T�RE��C�pZQ�D�CMXt{֔|R�D��Xu%�pXU��?=i��¶j�tA��l��I�D�#k�2N<Y�(�����a��hÜ�̓a�韒hRp�ІM�M��'�`���"�F��1P`����� �iØ.��KO>��.�L�J��� �=,�t�Jҁ��>n� �p��Y�p���y���'�"�!�'	hx�H���O�j��" B<2h�p���G�$�p��p�&�Ӽ��l�'$ڜP+��伔�c��j�$F*!����?-���R�}T�ax
�14v2�;Q�2>�Q���C�� `Ag/��Su�H[��#�����A�mrϕ׸'(�L��=y�ߟ���aU�pѪ�hN�hsnQ	 �Q"1����'Q�ݠ��`��̋�{�'������|]Q�b�i�ճ����BH��]�5�����сkj^��O4�a�֤RFn��;t:�#MS>Fq� ��i]
%dqO���,O���p����`|lBc�<W���pC�)G�̙���t���4��U:4m*_s���G�I�Zl����>IQ������O)�� ��D?�t��_�^��Lm�'�!����K,$����ߑ�Iӝ}�9����=q�0Itg�oܓx��%��yb�j����F͸2�ۃ��8��V=�i�ѐx"*%t-zy�OB�y�T�h��h�O����	G	Xc�F�
7)Q�i@2-OT�#D�>q��E���O�m�$�V;O?2U{Q��mMH8�r͖
�j���+C�WEXb��3��Wqe����
���P��C6L�9s�A�o|q��bK(5J:e���4�R�QR�V~��]�-
��S��>��)J>����O6��G'@r����`"�D��b+�~�'��#`\�L�2�H0(O�c/�\fm��_�?��ؐ�g] �'�lIٷ��A
 �N&t�� 	� Ϥ%�D��o"K�~��T���j'��j���<`困l �韒Y���tK~�	���:t#9ö)�eܓQ�`�Xw�U��f�|a��[��>R�]���#��>C�Nł"�#ae~@�A&ܞp�J��=�g�"!x��,�:�LP鴯ߤXZ�I)�ם.A⽢���{�L��m*�Ӽ��F�0�4� ZJ3��`#�Xq��Q�^f��?�$V%�Fi�`떀P
.�jՠF� ���8B1BC'7�PtaE�F�kL.WH�W� yB"I�W�T�Y��T�=�`"�-��'$ʧ
ܮ�� ԴȤk���t��s��;#�=�"O (�ҍʲ':�(��,W6�@"O~��G� ���c��>DP*�"OFaPd&��5/�0!�ā	i�i�"O�q�'@X�R#�� c�Y�5"O��B�G�$�Nx����[\|��"Or�"��H�}��$B�Vo��;�"O�P �T�e�G��Om�(��"O���aF�$7����Ɖ	�l�PF"O�����,~{��ĩ��S����"O�u���R�"�"�T���L{Q"O~9��.J!*G҈� W�`�1�"Oj��Da	;8�~�Ⓞ� i� �Rs"O��ښ:� �cf�ϞI�(A�"O&��B�v��#�ɂ=�ä"OΘ�T�ض���֘:+�!r"OT�����b`@=e`��`"O����熙x�}1��A"OD4��'F�ʶQ��M˸H��K�"O��&c�7p������8&(�d"O��/�FB`���-W�.��"O:xh5FM(+R�d`�)T����"O��ϓh ��d��`��AQ"OЅ��N��UӅ$�L��bf"O"	K�eD�*jԥ��^�p��-�e"O|࠵�ʂ6��1J/Q����"O��S"�	<Q�.  ��Ґ*��R"O�P)�C9Q��"P�v���"O��@te��wB�B&ʓzÜ�٣"OXyJ��^�f�Ű%8Q�T��"OH<����� kZ%�c�(P�Dh�"O���Wo�*��E#q�X"O^M�%"QWp����z����"OrР,�t2֨��G�s��0k%"O�ѫ̳w��X#f�õ����%"O�M���A�_e°��Q t�}��"O� �"iɍfw�1#���7V����"OD����#v�I��c�re
!"O�$`"���Lpl�૒Rmj�	�"OX�X�ߦ ���b�͑$eV\ �"Oh�fY)U(y�f�=5T6��"O�� CR�T���ႉP�Z]�A"O�p�)}�%�ӡ�>Z�8q�"On�J�I��g~�H�D�QF�(v"O�< G�RB�\��M-���"O"�9��*�qa��Q�o��A�"O�RL�ޞ0��.X�:X#�"O�Q�h���$���+J&pd]�"O��⊗* ���B�3�d��"O.A��Jg�H�	��ٜ/"i��"OZuZc�&S��%kg��9Iv�Ĺ"O7��H���S�@�� L~�@��:D��e㋪�r�BǠSoJ`M��H:D� �E-���th*�*̨S2��A�$D�r��[y���0�I\W1B�.D�X�a�o��G郯`U�U"c2D��
[]�}�S,�	l�t�B�*D�``V	�-�����@x��2�'D�ĲE(I�܈Ӥ�H *�^��*D�Ӳ˕)&����ǆX�"��#
(D�P�A�ΨX��,��ķ$u	�;D��0��a[,�G�C	S�)j�,;D��Y@_�Չ�[��P"�&9D� �c_�Y�$�~ȸ�B�8D�� �h�!˟Yt`	P�F^�k@�x��"O��1�s�ν��%3����"O&8�dЉP��d��&#��"O��j�3�\)���̤Q�U�7"O�Ep&ӌz0R�e�<4�]�"O��+�(^$^��ё�Y�N��ѱ�"O�t��ĦL��aJq�@�+�֬x�"O�9����K谴j�叙a��4"OnhK� Ӎw��u�2�!u:`��"O(�`q#��!3��G�p(Ԡ�"O+bA2!:��i�a���18ԧ�P�<����D$��l�	x&� M�<�gΝJB�Z�U�j�c�b�<�'H�U�*����{��l;B��S�<���F�FE`�KZ�F�x���D�<� *\�TT�t�Da ���H�<�!�Ú}T��У�T��$�kA�I@�<!$� %D��[T�M<����@P~�<Q@$�
F�:ts���
x9��d�o�<1�+��d���J .�C�t��7�F�<	5JM�y�Q�T�Q{��ӬB�<��� 1+�=*�"��[A��D�f�<ɷ�y��
ǎ�]&<|Rp'�w�<��o�1RYz�1�M��x��TZ��]�<᧢�:t�Bb�
��!��Y�<!���>(�4i�g	�2S�-᧧�V�<qw�kJ�H��gM\��*W)IR�<���K-*2��*Wn�;��9���Q�<����u F(	��U-���O�<�C�W�Z"pM���&Xx	TJWN�<��AL�Ƙ�2��).l9B��F�<��k?2B^�hǡ�34yÄN�Z�<%JS���$�۰-�<�Dd@N�<ɴ,��Y ��;���>�$e;rd�G�<!U_+ct9	�H�*�B����z�<i#Jϒ VҘ�&��(T���"Gy�<�Ң��pY�D���l�yeM{�<��$C�Ql1����Q[p �v�<i5�S%A���:'@Ѝ.�@��`�Zo�'nў�'ޠ��s-�8k�aBIY�"9@���I>vUIpcR�25~�r�C@55$�ɇȓF�L[p�L����XMh��(�ȓ�@��f!�~�48%��3 ꄆȓ̬�82)�"~�L�S�9DSh��ȓS=�����0}� }���6+�Z�ȓ�1`�%ѽ8*"T{���20Z��ȓK�x+�� 45���́��$ф�E���2��~�T��#��g&�=����s����#�"����m[�{��z�=D�䛖 ؔ �8 JφL�v���:D�(��Q:D�rɅK�'D���$D�$b4D,��i�#A�"2��R��!D�(�ʁ�dD�-�@C�?4���0!D� Z�#E�}��QA���ys���0�"D�<�'
?#S�Y��bM�M��A� ��"�Sܧ/@�ܻ�Hw��}iT���*���^�n�	Bק?���6@B�&>�U�����l�6Au�b%�H`���ȓ*�����1��Q� N�+�:1��.��Pd����6RIE}r��= ��	:�72M(C�Z��2C�ɹ�\ݪ�f	�8U�M�dL��c��x�n 5_~xa����r�
v�?�y2��,7�����_�cY��&&P;�y
� @�p��4e�hE#!0i��0�Q"O��
���|@tҋ����"O ��t(��~@�g��d��%"O������RgN����l��9"O�$��� 5�>� ��#K� x�7"O ��cR4*��Pѐ�,~(u��"O�8ra���ŉ�
Η�t���>Q�%ߤ�R�I�?X�~����
xm�=�����D$��nZ̰���@�Q�ؤS�����y�`V�j�6�"돇DC�l��P���'	��.��|j� Ǡ`�,�t��E�.(5(�`�<��níH�Ṿ戔�9�Q�! [�<Q��-@�l��� &�^��RNI{�<�Q�ڪy�n钶LSzo|�!�x�<YGmAi�H��	��#�ࠢ�~�<ywA]=s�4�Tė!k��cS�<aB(`�]�G&�3�CΗN�<�����ˀ�G�
��A�<ٗBڭKs|�j_NE)�Տ�T�<!% "'�F��É�	F�0�We�I�<I2l�
t;���š	�o8�Q��K�<�g��C;�K`�UV�beE
�r�<1uEAcޙ[$�{���8�r�<�pc���r��B`V�Lk�s�Eq�<�#鞁�6����ɨTȢ�* E�v�<�oA�5 x��v)§v��I�fu�<��i��1��⅍JZ���B��w�<$M�J,�Ԡ@��a�r���r�<���D�<BT%F�+Q*(��`�I�<��.4f�ڜr� �oPh�w&�E�<�$m;�T�떯����7�~�<���HSNF�Z���@ȸ�F{����'d�ݒA��9����éɉ
�x���'%�yA㧁�U�%��D���l��'��\e*�Ti>	+��P  �� �'�h����K�1Tl��G�u��5��'<B���Bөa����� t� ���'�H��PΈ/OjX  ��`�=r��$5,O|�!�D�vre�����7���C"OĬ���P�LI�@�C�W=���dM�WH<a���w�	!���TTʐ"`�k�<a��/���2�Q3>�'�q�<����C�\(V`&�p��A�x�<9&�_X=���،9��
�l�<�S�Ɍe#�@���!>�Z�C�Cj�<R6?/��`3n��JH�ۖ��J�<�ukI8"d<ب��
:���Q�E`�<����K�B��h Rd���%�R�<�4���}����K�xp���L�D�<y�������S8���ñ�@B�<���0NmJ�k�)K0��B}�<��hC:(~� `(��=��w�<	�!��CPY���m�\����u�<�Fn4�,5�bKA�`�N-�q�<)���;Z6ƥK��"7zi�`�A�<�Ė�	2�,�犋o�}aը�z�<�v�^x��q��
1��x�!�	]�<�É�:w! �2n��%��2���M�<ٕ��t��H"/�>�|��M�F�<���,H��)��O@HZNM*M�<Ѵ����d�!� ':8��F\H�<�w�
�@�
X%m���!���[�<��O=T<�8c攟t����o�W�<��&
��@pF�M3@$������w�<� V���¹�JQR.���"O�0��!�p�H�׭N�_1�"OD�˵�O�H	 s��ąT󆘱"OȀ0����i����u��Tj�*O� s��Єhcūۏh���'�>�x���Qab�����dĊK�'�B���.w���9bE�&}�!��'��i�A�b�fA�Y`v$��0D�����Q
'p�Q��0Szl��r�+D�,�*X�1Zt��׸u�N��G)4D�+�H��9s�"J*$F����2D��P��H�
�NX�TL��4I�.<D��A�+Zl�ȸT�ߣ�$�C8D���GށXv��� �@�=���()D�T��i��Q��]���S��� ��(D��QdM
gv>��OT�!2�q0�#D����³$�t��BT c�%�R�,D��x�;�����ϝX���rF�0D����.�J��i6$�30V%��H-D�����
xj�EK�`X�N�p!�!�8D��� ��7H�=��'�8$4���H9D���B/�2mjTy����,]�C�)D�X���=t=��K�@�~��hCn'D�R��8vꢶ'�Љ����&D�|�`C��B��0��N$<頀�d�$D�X�4����͐��9>Jx@�"D�88�d��[d
���
�t�i�g$D�$$R�:^��D�A�` %96�%D��iP�	")�6m2�E1˸L�6�"D�P�'�נs}F��s�$r���p��?D�����T�$B�,A�"�b�5�?D����<L�@�r	�pH,BP+2D�����\a	�L��A�TZ8���.D����ƣC�i�a�@	pi^!@G,D�d8F���z���Ta�6+z&��p**D���e'�}�8)�k��� �1f(D��C�'��9�g�W�h�=C�%D�dC��L&�嘃��'~eQ�� D��#�kK�ܩ�E�vx�,{��>D��
d���[�P��Q/ؖ7�0�1D���ďՓj]�W��j<
d�5}Y!��N�|�0�E]�4�X�Z����KD!�Ýd9v��ѬՐ}��A3JZ"2!��G#t�S��H�/���q�8D%!�+U��L!���D �-�!�,!�Ě آ�S���I]( �Z
!�DF('�L�Ӥ$�锍�}�!�Ɠ�\9P�cڙ=̜h��	~!�Dۯ1�� ɇ(Z�vh�,hǋٖ&!�d־NGj!���I�Hcj%!P���r�!�D�C�`�3��f�6S�C
n7!�D���L(Z�`��^N�����xJ!�d/	d��K�x�Q���o=!�LsQ�`��j�B���yb#Y|3!�D5�%�a���u�VU�R��H!�$�d�N�o�n�a @L��S�!�ݡ0K�\�u�� g�6�ӡ��	~!���!�Δ�.�;��z$��>j!�dk�j���@?���S��!򄚁9�&i����)^��7�Z�0�!򄐇=©{�d�"v_���T�p!7"Ok�G�=������#ۄ<�D"O8��t =��`'.<&0 B"O�X tGԓfV�y%��"z���"O� ����7v�X�%� �捛E"O�Ի��O�2
h�a��f�$�q"Ob͊�gņt]����d��P��"O
�:�A_�T�P�v�a�^���"Of��뗂��X��o�Mg>�U"O�ĺD�o���� �~�f�I�"O⽈�T�l|���ò'>���"ObK�'�*2(�����_~%rE"O؀��O��b�JH#k;V��� "O(�M�|���"+��kJ�=��"O�(1B�'RB=�Y�n1t�Hv"O�����	8��%��P9̰�9 "OZ�F�\&Kﲄx�H�	o���(�"O`�Z$(ٸ@ pҳJ�5���J'"O�Hp7g[�	�	�
�,;����`"O %y�J�#{�\�PHїlj&�У"O���p 2�`J�g˩(�^(r�"O5�q*�ޑj�ݷ{�"OD4��*�(7�j���g�J�@�1�"OtiaG#��k
�� �E��0�"O�|0�	�:,a:)+ՏC�d�$��"O�l)��=d	�� `^>�����"O"D�B̒^��أ��Y��:�"OpU9�EO!/� @K �Ͽ-���kb"O���F�Y�2漀��Ӓ-�$y�"OHDΖe��=2T�7��t8q"O�!Q�`���"H�.�Qj܏z!�$�<O>D�"sBl�`*s�Ƙ[i!�dȎEZL�!��Ǹ?��u�ʇ�B[!��N5lha���G2�yBg
�uW!�ă��b���<<֍8'�"�!�
�w �x�N8/#��@�G�?�!�#B�}؀�D�[�°��y]!��"�B�)ۮdD�R��C�!�ø �8�X���sR�p@3�̢[�!�	�`D�k4��7v��2�AM�!��W����(R�A�#���0BO]z!�D� MҜS��2qf�ku@
��!�d�6���9��_�` �m��x}!��O�rHx'�����YS�H�}!�� 7����$!0�"vKuz!�$�73��B�c˖"Ϫ�P��k�!�ğ�K����!����Jw���<�!��Z?9	���B��n��x���9B!��	��XHtm�P��V� ,F
!��M)a/d�X��n$�9�ϙ$2�!�\�-�H����N>5�pC!�d�rgj��Ǽ2*�u��v!�\ I/>��t�߀21�X	�Y21�����2���p�@d{(���)�"�y��D%z"��Ls�X(b�4�y��$C�48�Hy5d�8�Օ�y2`�?*��{t�8o����A�
��y��Ì ����%߃g.> ��d��yZ��a2te�b\{T�Ѳ��H�ȓ0&�H��ռ!ϊ�"�A�1'�,���a�= �J
o�V��6�N�ek,-�ȓdB��"$�a�PP"���.b9l�ȓm��\�NHQNzȱ��8Ψu�ȓ15��6Ɍ ��ٸ�o����y �%�9B>��E	pȬ ��U<�""�Z�"4�h	�m	�6�䍄�8~<ktBX�R�������z)��ȓU�x�F��	N� ��̌28���S�? ��çk��L�2')6ƥ`F"O����ܤ0�J� ����Z�"O���h��(cg�3l����"O���敭0���e$�&-wpm� "O�� ��>ij�q$Rv�[t"O�:`��^h�cU�9�� �"1D��c��5.���l.4����0D�0�!�ŧ`�CQPugv��d3D���Jd>�i�
<��I���/D��� ��3���H�`Ҽ+����F2D���p�_�C��z�ᏙT���`3D���Q�T*XIX�)��&V����0D����6P����G��=�U�:D�ຢ匼?�R�{�b�./�P+d+>D��*��H~x��5C�I�s�/D��Ι�68��5 .j!�l��$'D��A��u��#�wL�� �/D��P�j���a�-O-t�Ą��m/D��C��A�;&u�s%�f3�!�*0D��ɖhJ*"�iK�ʘ4�^�#��,D����&�.i�MT�X���iSq�<!F�M3S���(�ր ��T�B�k�<��˵G��]`���U%�,S��Kh�<q���8Q��LhF�Bf�� �f\�<�gk=�X9�um�N����`�<��W	.�Ip��Q�����A�<���;:��XB�H�
�d!���b�<�$�-Nԑ�@瓯v�^,:�&�_�<)�Ʉo>��f�#5i��� �c�<�D�E�T��Ȓ�a(��0��T�<y�. 5�>�0���G=�8q�@k�<yR�ľr�����F̤D\�!�Uf�<!WcԸ}�Z)p�Aơ;���c�<��ټ"��1������itet�<�$�X/`��̚nP��:�3#u�<�4
��.�h��J�k��1
Ct�<�ƃ	suܔ����
~�) �@e�<�G�ʆ:+���d*щZ�X�QuV[�<A�hWB�&\a�jMY� 3ѡ�^�<i�-H�&�vA�  ɂys�(��/0T�,J�Z4&��m�$c���yb�T�
P�=hG$��.�#gf*�yB��B6dq��1*� ��1$E4�y�*ܲ:�@��'E�-���G��yR��"�>�Z'c��136`:b���y�G��G*D!%�U*T+��u��(�yb.W�-�<�Qk��E�8@3����y�H�	��%B�7�ܩR��0�y��ऻa�en|A� @��y"��J�Vaa����VG����n(D����*Ӥ5�<Ka�ޝR�b`�7�0D�@�'�U��I��;��9xJ/D��BE��3?���A��2}d#�+/D��a��#PԽ����C�Nݓ��9D� ���>�`u���e�pU�B<D�� �Ӫ4�^����\3n�.��FB:D�j�J��3z$j�ֳ{��-3D��P1��1�m�D�l�蹃0�3D���0 E*B�1��gލD��-�L4D�d����V�	y�ݴx�u�W
=D�h���H�V�{e+]3/�z�wi;D���A�W�:>@�#��(E�V�(��7D�P�ѯ�9+ZZ��7k����T "D��0� �&�$�1�FV�O���i� D�� �I�7�&1�XC��L�^$�"ON�Z`&�/2�����X-c�p��g"O�9T���D�^!;!Cݻ<U�,��"Oz'bߋM�Yx�"Ƶ>��v"O&�1CEB����+p��
=���`"O����T7<�E�)6&D�C"O�m�����i�JF#���"O��Qf �#L�f��C΍nf�"S"O�ڠHT�&��5爎O���"O�4�T
H�sYX`#�Vh8����"O*8H�I��/�|<�'�ֈY �(!T"OЬQ�&P ���P
XP@i�"O�XY�n��ǎ�3��|ڼ��"O|�!C.@#����Ս�`Z�,j�"Of]� jA�=Bh|["����8�[e"O�,Ie���q���x<2�"O���Uu�t	�ƤQb���"O8T��.Z�R	$FƱ,NT`3"O�]�Ek��r�l(2��,8;PIb�"O����	�U�� ��a(N(A6"O4X
T��{� @Bӯ�v*x��"OjT��پs�>�k���af,��"Ol%��KA�j��E��k�>`�8*�"O���HX��[B�ģ7N|hK�"O�Hbr�?f`�Xڄ)�=x*�A�b"Ox�`�-�>8��t�pE0x��\��"O�H�b!Y5�4%�G�G�"O�캲�ٵ-m*< ��K�,���"O�q���'(!�ITn˰zy�LP�"Od9A䠄�p0�U/C�D �y��"O��P-O'gL��"����۷"O=��+�e�j����A��Ȁ�"O�u0��3�>�� ��}�<�32"O�L+ÄU�_V&��U[�;�f��f"O��Q2Oǖo -j"À"W�@	��"O�s�D�$q��Ӈ	�]�xX7"On���N@�.�Q��Za�h� V"O����@�xV�U82Y
H�rع�"OV�i��>U>B��CJ��*���"O,��/׉�HKPh��S��آ�"O� �jZ�hE9'\�  B"O:ES�[鬄�t��x��d�E"O��@!��~��0�
y@@"O��U��6��I�cx��B"O��k�Eє`�Ⴤ��1Al��"O��*�Y��D�Y�&�` 
,:2"Oڨ
�!�/'�Ss�VJ$�z�"ObUK�/0��1ှq2Ɂ"Oڤ���T|����G�b�z�"O8�kgM�\��5kf�ؽl��) �"O	c����]����d@� e$�xp"O�$q����w(}Hp� T�����"O-�F✻I����U��4y�
��"O�@� .�$�*h�g��;��y�"O�ې��2���R�DCi�x��"OF��W˖Z�V����� %�"O��x%ψҬY ���^���c�"O4�U�IRވq#�X�ֈ��"O�)I�F՚D84)R�W�;P��V"O�i�4oL)�U�� 
�B��e�P"Oz@��Ø�����\0[n(C"O� j����(��$�K+H[L�2"O~u@�OY�0:N��7m�/h�j�`"ON�F��G�4pHf��7�^��"O� ��a����u�*����Nh:,HK�"O��2 ��U�̐,[ʂ	v"O!���� ���:�eV�I�1a�"OL]������ȩ�鎞,���5"O���w�4d�����jᎹ�$"Oʌ 3g�7�B�'�T��"O��5(�-�t��w��m��8q"O�i*N��б���-��C�"O~e�r+�;7�nm9$��5u�V1QQ"OV�)� �%g��1D�'/�\�$"O����
�? T]i �@�,��@"O�YhI]�<�4�ha ňD5z��%"O�y���K��)1��'GĨµ"O��U�T�l�#+E0m��{#"O
�0B�P!{�(Ze��܅ "O<����K!(G^i9+,(Ԍ�i$"O��Y#l�-o�8iLT[/x�
�"O쨓MUm")�q�@�0{��/T!��FvZ�)�g ���ز����!�Ώg)���Ү�Q��"�;f�!��Y���vƘ��&W��(G�!�Z�]@RiJ�<�h=�s�� �!�M�Hu-�i[����a]|!��L�m���D���܊T�>DA!�$8��hS�DD'�"�c�/NTT!��Y��y�W�"����t�Z�97!�d�TrY E&G�g��3��ߘ;!��'^걈��Z=�,�p��S;!�d��dE ��f]��` ��rM!��V�)�F$T�mz
8@�y1!�$�{5>5�4Y0! �4H�M�)!��=�Fx	dB^�<��qbRm� At!���^�݂秐*�� ��
JE!�X�Y�D���JM
�x�7K3!�d��0@�Y"�fƾ�e�ҟb*!�d��FJ��k�=*��HB�4!���6y�n���̶7�t}2�ud!�4D�� P��9�8��
�)!�U9 ���6)�n���zj�+!�1JOZ�	�@�H��4�	Ò�!�D�M��!�٧ǂ�X�*�X!򄕆��1���ߚh��!f��!�$�p��$�\���%C�پ !���~�L����<�����L�h�!���"u��R���0�p�C�$I��!��0�`�;�,���Ĩ'�H1 �!�D# FH��A��,q��M
(�!�䀆/�Hmc��{�6q���F C!�D,(V��5B�^�r�ѥ��S!�$� /�\i0��W�]������D�!�O+;l��!�,~b�Eh[�t�!��5 ����6g�:�n���M�b�!���0�I�T��I��m��H��LF!��j: �	�n����h�WgAD!�$�>¹�Ն�7X�M����$8!���!��d��$ՋL}N���V�H�!��27�f9XP-�Xt�X%+��"�!��<4�Ʃ��MJ$Y7||�u�Û�!��?;�P��h-��E�CZ!�d�� ���Z'MWDՠaFʾc@!��3r���p����\�X��Ő�&-!�$gW2(@���&! �(���ţ^6!�dJ74Ӭt��MŤ<�4�n�!��PA�a#�X1N�Vu��+e�!�� ���c��D�(�kC��6ɔ�S�"OIZ�τ�.`�9�B��qh"O$u�%�C-+%@@4�ȘE�F,�"O ��dT�">^ݡ��1A�L@�""O���H�%WڑJ�f�c��h�E"O\�����Y`��P��4�Ie"Or�C��Z�4EЁ�Q#ƒd�p���"Oz�KD�(>�����#T-w��C�"O\)"�m�5�%�V9k�z���G��yB$�6W\�#�ҟeM��-M-�y�[�$=he��n`)*����yrO֐���-[#W���Gi�1�y��Q.SO�l���VE#.(s���y�"�*�C�@C8l̺a����y��J\˒�ܕ.�������
�BC�	�Wn�p�r�L=&���ĉ�6@�PB�I�7|�+faV��ò� ?�B�I\3|�@�i%0~@�s���-��B�$z�#��ףw����Fmu�B�ɵ7�p��t䆼W�~0s �:7XB�=&
�	�`T�\OB�ҧŜ0B�I�ΐQ�P&����q3g�+x�<C�ɮl�b\HF���[�`Ǻh
VB�	�_O��:�(&ɴh�a�Y63 $B�ɚrF�NS=Ƚy7����C��:<\�Ѡ�N�'=	N�2�*�c�C��1_�"��ɦ�dء'ē 1��B䉭%I6m22jL�D5&��G���B�	3F-������J�ZzVB��+è�Z@Ć�.Ff��Wr\B�	nH������S���q#$��9�:B�	2Wh���E�Z�f�X���#�C�I���E�j,Ś���lmlB��-C�J���G���Q�0�bB䉻�P��雳Kʊ��1b	.B�I?(���#�Y�t���&J�=1}<C䉿�~��cR$ִ�K�LD/:C�	�+���A핾UD����Tu~�C�	?�H���M�gn�� ��އ8�PC�I�H�]	Z�1�Q�V���5a&D������2��%*�ԓP��̸�$D��x#���?b��2���v S�"%D��*� �)@P�%�qiA�5Ln��(D�lqE
M�@�0��%^$l����8D��r�K�~jd��!�]�&K��6�"D���͚�Yv�����'=^8l#��?D�t���Isߤ{1��?���3� D�b����Z�T�R��o��Y�"D��0��NKLq`i��M .Q{Ƣ?D�H�1N̿U��@��A��0rq�#D�,p�C r��9����nJvXbU& D���D c�X#U��I�B4�QE0D�D���@�R���'S:�BVe.D�\`���a�R�����&8t��0D�x3a*$O`��r�U�;��!��*D��c�F��^ճ# m�q��<D����R/M��T�(�5��6�!򤁧@������ˢx~�@��зC�!��<`",����\?C� �eA�)�!�ӧ�ȝ�a�:@���媍c�!�D�,s���`!j�,�Ĵ8w*F�<!�É*w
Q��g]!T��1��>%�!�DK�_Ƭ���9cL��k��P�H�!��Nڍs��!�%z���)��B�)� @ĈbnPIz*�S�(��J�"O���`n\L��;�g�.
�,�P"O�
ۮZ�v@��%�а`�"O�� �e���4u1�b�.�K��y�J���
�r+P0�U�U2�yr�Mc �b"@#
"�i��Z��y򨊿��Q��"Ў }���ᮗ��yR��G�2�����+.��E����y�ˑ�
g�(A���vJ�b`����y�GQu����ɸj�p\��"�y�f�,�|��(
�b ����Ɏ�yŃ%&�XPh�k��p�
	��ܕ�y�GQ�'z� ��
k=��)ç�>�y�N��e��s_H���K!�y Q���,)����Y��͂1�Q-�y¢	�v�
h�7�T"K]��ʑ а�y���K��t����A���
0ŋ
�y¢�/�(U�!
F�7��)ׇ1�y���_� ����}�F4A�-��y����H`��m���mܜ�y�*(���i���i3��W,M��y"� ;h���Ŕ3gp��Վ���y҄#���z��S�KJ���$�݄�y�V�]O�P6W"2�<C����y�40��QJB囶d�]�3*��y�NM�UR�y�eݦ�\UBg���y��ưVi�4�2��P3Mc5�Y��y�*�2Td��{0�.L������R��y-��! !͆�0�p��+�yү��X��]�Sbޟ\!��#�ږ�yb�7kNQkSMZQ��:�kA�y��^U~��^
Q;ȵ�`����y�̄�
G���?�*)� !��y��G w&��i�� �<�9p���y� �����7��d,�8WO���y�M�&l���)��#	I�)RuF\��y�N�O�vss���Ԕc��M=�y$��j��*	қ�����I�7�y2	[�2����D�'\�ͰS/T��y���0F� BJT�D�6x�K��y���K�z����T�(5�E&��ybg	_�q�#�DV0X
�"�y�kD:%��ٺG�
m�u�d͑�yRcL�yn�� A���j�l��y�@p�bİ0K�ǌ�[��%�y2�RV�%R�9�x��N���yr醑g�:e3��A21�(9q�ϗ?�yN� L���÷�0>�e3��(�ybq�L�Tl�Xs�ջ/� �B	�'�P8q �?Q�С�CE����Q�'�&1 ��-��X��&�+=68 �'�y�qLHnެ��)��q4��'{��[.R�Lta3� >��
�'����
jPf⚰v����'i��t�E�"�r�"�C�)r�.��'K���Эӡ;���##��=6;�$��'����2�ϔ$39���3/�,���'q���D z^H�Y��/'����'@���
����*�ߐN2p���'��D�P'ϥ4��t�aC�;8�>���'�0�IW�Z�xA�.W�ع
�'�X�"O�FG�8�ᖆ<7���
�'�,��%+����I��+�O�y2�L����C`���|��.��y
� t�{��Q��t;4&�*�d"O�`1J�
j��U��e�0K��(��"Op�T��;��q���co���5"O��r�EQ?Onz�@rBH�so �C�"Oh]Qg�U�I��m�SB��Yz���"O���*��j�z\Vk���Tp"Ol]�~un�
#-C9wd���"OJ)K�� 4�ʳ�ׅdm��"O���Q#</B Ja(ͅi��@bU"O.�d!�A��%B��͟B�����"Oz��A6cڢ��	��p��D"O�]{��>���9xκ��"OX�:w��2fW*`�k[��9�r"O`�QG�)�B�(F܎pSP%�"O.|
��ߑdqT�Xˆ���у"O�L:�[[,VE�R���@�r"O0T�'��[Ҡ����� �t9�C"O:��d�ҩg�@	�!<wt�=��"O�e��d	�qXm��sb����"O.�P��P?��u �e��p��"O2=�6�L��X�� @�rUPp"O��R��1�襃���M�fi9�"OV�+$B�aFLqg�*[�$�C"Oh�d���-ɔ@�g�4}"O�p�Q�ʓD�\���6���"O���%7���@m�5�y�"O�y�QD��@��IQ��X�"O.M�*�/wtp�@ba�5C^9��"O��9b�O���@Q"�f���6"O�PA�\�;���c�#�5a��\`"O��`AٰX�����
���"Oځ!��ƮUpI�F+��'"O
���aU�$笌X�E���k"O�X��A\�1N^�QTCP#���HF"O�\���V ����H��x�<�#�"OP��q� *1nt+@H�!9��y"Op�*�N _dBܢbE��v����"O�Ĺ%kY�
[�Y:��4-�t���"O�yq'�5K���b�<F$T�;p"O�dj�ďuB�$��A��}ĉ`�"O:`��9а×D�
��D�"Oz�{#�Zd��:�OצSOyB"O|=�gO-/ϲ�S�#`I�e�W"O���W�JȒ��u�ԭ���1!"O�����W1���� �U�&u#F"OH�(��P 	��a�
`���1"O3W�2��Y�*�4I���""OΘw�_0H���
��b�ԍ�"OP�{����xaT�2p�2)�"O�uhጚ�fVui3��2�*mq"O����D\���h�MI�p�Y"O��9��P��;�ƒd���G"O층�J.b]�#�$ʝ��i7"O���4s.�a�F"� �`kc"O>�Ył]�	��أ֣�<�Nl4"O�i	S�"��Y�핕\ }P�"O�x��6q��{��<N��"0"OT	�3��?F\�+JQ�t4XR"O��̋)�ܠ���U��=2�"O�tʦ�5���h�BV���"�"O^H�ӣ]�$+���!�5�*e`7"O�4�mؠvS���`��l7L�q�"O�t��O�$-LDЗ��N��"O2����Wj�qև�	��8`"O� ��N�'��8#�ě�F�,8��"OF�jED�2u"��!��$��QD"O�a��kQ!q�<�u눕H�&)��"O��PI��B�l�!�+&2`e"O ��&�^����R�=��Xw"O`�q��ɂg�37�&q�(���"Of�J�'ܖ��PP%Jy�$A�"O���V��o���+�rU�"O��6B�jb\д B�pd�Yhc"O���˞�I�e
WE:o��Y�"Oz��G��P/b�9A ��I"O����G�+�*H����h� I4"O|I;gaN- �HC�A��?�؀�"O>ģ'��z�҄��jŒ{�N$1�"OrX���=N�@��gh��"O�`��hƽQ������\�)df�"O�AGDY�P�0��p+�d+ ��"O𱡱�I�%�ri2a��F�0�"O��� 	`�eۑ�2*$xK�"OZM����H�L�c �
:��i�"OH����7L_�]�� �P���U"O��T�K#g�<`Ӕ�^*�:�q"O@��!�:+��(�1NY�}l��y�"OX�(ǚ�HTL�run��u���S"O�$�W�HHd03&M�c���"OX-
"ā~
piD��%MK���"On��cb�~G�h��DW�.�Ɲ�"O><yb��
�����N�1�D}c�"O�� Cʫ�*t�p��*#�bhr"O6	B�m^�q�Xt�1�d�("O��Q�� ;�*�B����&�.j�"Or��Eg�rR``�C�J<� �"Op	y��T2v$R���$];��
�"O8HEH��xLR"i�s�>��D"O�y�U"C�	L�0YF.�$>���"OʬJ����V�2M�p,$�Ɣ�"Ox�jV�R!q�b� U�U,.�=QP"Of��0���~� s&��q���"OT�1��37Ը�*�"��h�Tm�"O����įW�*	��L$ͪh""O¤��M�yP�e��Z�P0"O��u��#=�(]ȓ�(��1"O���"K��D�*���)J|) "O�N��t�:�R��8����Æ$D�d��\�c��3�/D�p�Rhs�
-D������
&��¢�B�O� ��+D��+2O ���X�iu���7�C;�y�i/�D|@�L�P$y�U�\�y�Cȸń�;�희9�Vɹ���yb�E����K5�i������y�i�:���B��YO� ��פ�y2�7q��u��l��Q��@�'���yb�,&<���	HS�xA�-޲�y�/ۀ6��`,��^:"�f%���yr�PG?F�q�	QŪe�$�y�
�m��+ŝQ���Q�҅�y-����)��ƱM�l!j��:�y�n>d�J��ˊw���7hS��y�,_�i�"M���!뎍!R�B=�yb%��`|�g�*rE�IbI���y¬%W����ȰdYL�[�b �yr��+'���F/Z��)�F��y�E��:���"�l��Lu��Q/�y"�Ǉ^&�<�DH�G�~� @E�'�y
� lh�Qo�,!�1�#
�y�´�"Op:G�RI�ܝ��O_�L��H�"O�1��(�e6�D"B�$��4@�"O���B�&�y�ū&_��s4"O���l���尃H4^���"O�l���_�FtjAC�&�"~�YJ"O&���86_��4#��.r�Mz"O��(`(��@疜h��	'h:x���"Ob�I1��%��Y�@f�>7/*	�G"O����%�A��d�(Z���"O���w��:��̠�T.	����"O��ic��bm� �#i�(W�x$0V"O�#e#B���D:7�H�]��<�*O����m�Œ`.fP�03���a�<F�Xe�mq�ː.c�ق�JD�<�d큧*��H�5�	++����"#w�<)��դS�����GO֑�BE@y�<Q�e�MR��Y�Ȏ�tc�yJ��E{�<GK��S����BD��"0��u�<ّL�TuL�;�W�k�Dt2 �p�<	�a�!e��@�'O � ��Xk�<���M�G����惕� E	�Gk�<��n]'�x�!m5�T��(��<Q 䛱hg0Q���g��Pk��|�<��iD�Zx���iJ�Bf�*t��v�<��� D\Lb7�Rcۺ���p�<)�V?0Y�5S,U9 v���p�<y��дzXIڗ�YA�u�.k�<�#)�?G�LU�A�I�܀�C�c�<�2�%�8�K���/_��Vc�<�f���g �i
R"�X"�DBCd�`�<��%�=kN��F��8:R��_�<y �S3*v�u�ӭH�$�tj#*BC�<�G*��,��y�s	�qj� � �k�<��Ǭv�x��]�]G���s�M�<1Giޟw�83�h@�Z�>��\%!�O�gg�=Q#�\����5��;�!��$��ȡ�'.jo�q���'���Ą�Yܠ��qj��"X١o���y�peؠ���g����۬�y�d��@�\�g>4 ���D.�	�y"�C�Z���I&�^"WL�� �˗�y�
P�=���ѷQ�Rq��Ϳ�y���7I?����C3�
]P1���y�� <4����K��f��qKG8�yBGm�$q��bG���!�Dͪ�yB�ȿ�<��R��!V}��ᄸ�y��к֬(˕I���I�	\��y�t�U��!((H�����y",�;-˨@$��R����f��y�KՋD"�]�e#D�(A������y��u�$d�r�8kbܸ4!T�y�mD�T�=�W���2�6ł���;�y���8�R��W,J$7���O�'I�B�I+���$�S�*3Ą2B����B�[��1��q��2琽P��B�	�pxpڠ��4hd��JΔW��B�I(�b�
pb
z?2%!u�0SfB�� M���(\�/�1��E��2�6B�I&U��"2��j�aZ�TB�ɤyڜm�@�N�(�jɛ��٘GM�B��*3U�\Q�$ �%>T�i���]�B䉧]�Z���Ŕ�m�ޙ�#(�npB��%���FW�?ju{ ����� D�� �t)�@܆�`� �) j����"O0����@r�J��Ȑ�4���P"O��⦪Q��n��e�̶n�i�q"O����	�6D888�  Ix�`rq"O�ฅ����RxZZi�B|�1�XX�<��#S%9��@�C^�(��#��y�<���8;;ȁ`����1�D��0�[[�<y�)�,i �εd�Fh#P�WV�<I� J�48�lR2��.Y�`=#��U�<�񅑚N�BYJ�ڦ3:�G��M�<Q��)6Z��2�"]�zM!4�OU�<y�b�,z�|k�%G�C�i2��f�<Yf�:5�6�i���{�p4���H�<a��߽ym���? �Fȁ��G�<!萀JҬ���ٲ��,b@��X�<�6H
�`�����@[�lx�yҊ�Q�<I �&�^�@֩�	��y⍚N�<��!G
�d�����R���.HD�<yS候B�x��H�1LP	�B�<�!�H�s�|�c��`S�e�����<ї �9�|��"�*I�`b�Me�<�� �6cJ��� MP�Y�vr�-�K�<�pJ�(xeʝ�q�%R����g�q�<��.3�ܐ0���Y%8X��Rc�<Ag��(������3e�q0��Ay�<q��U��$�KPMЅdlɂ�	R@�<!�D�A�Ɓ��cJg�B=����s�<�
��i����%��T��ATnh�<��U�Bp�����ɭ^Sb��L�<�ʊ�E`��w$M!]TLA����F�<!1�H#"�Āh�d�a�5K5A�<�@I��r�`[d\.=y��}�<�@��Z�����}Lّ́d�<1vL~*@,;���0$��bwe�v�<�&��x��K�,�x:P�]p�<)��E�f�$�*@YF-ʐ@�m�<ij�jyv��"/Ȑ�a�e�<�@�4���XG�@`�F=[��e�<1v��Jd�(�&��g ��ꕢw�<�A���ic��t��%���J���v�<Q��D�t�XE�KD�^��c*Cq�<��$�[�ĩ��*t�=*&(p�<��/B�5$�A�ٮd�8�9�h�<iRW!d4 ���a4l�13�K`�<9�#�+ ̀�C�+-ZcHLcw��f�<���^�. ��\*<�^�js��^�<�b�G�	�p2�$ԧe���}x�"O��F�ܲ,) %����={V��6"OV�
 	�vi@wHz�v��"OP �1��3{��``�' 1!��}�Q"O� A��]�U�*��dW,G�>�h�"OP��IB�M�@p��Y�ȂD�A"O�AR��R/=�]Q�����hC"O����LZ�XKܐٗ�R����"OV�"�%N	(�B��4��0h7���"O����B@aP�q�3�U��"O�9��b�"Cd\k�E�6e2��"Or�R��d)H�K���Z\�e"Oz��g

�$�LB�l�7z�>4*t"O(�!B(XNd]�u��<D�jHB"OL� �)>2t���$dݺ��%"O6M��'s�*�jqhV8� �)�"O0��k�JE@u�R�G�l�.0xs"ON=�@�%p�0 qoߵ} �M(�"O� �ER�L6_)�0e#o�Ĩ"O�� �J9y�	2���U;�uz�"Of��wcF��@�`��۴6����"O~����,/P�(�7�/H4��"O@�Q��X��\넡Ěa��v"O���ǎ�4@R�"�)Ȅhif1Q"O�y���H�41	 T��gUZ�P�"O��Sd��<Ji��N���� d"O�y'� ���H���2�TH	�"OJs��CnF�y5#I�1��$�R"OT;2��"x�2��(!F8U�"OF�rK?n���؝RD�a�"O�$��)͏ qR�ƅ:e�e�"O��2m��ء21�D�L����B"O������+�� {#�Q<.�z�j�"OrhJ�IŊpw��r��c֬
�"Oθ1��}&��.]8J�eT"O��ш�rG���޽1<p ##"O�HfG&̔�!Ð�U:NUcg"O�D*S,^=n�昳�˕s+z�x�"O��S��'B�X�K�>C�4�2"O֑��]:g����J�]�pi'"O�A��X�nb��;!HW�c|�[�"Ob�Y�D�[�@��1�^�Oi��r"Oz�2����!��t;7GD�Ku�д"O���d�M��; ��5_�q)"Od`�e���U�EȐ枠1=.q	!"O�� K��:���d�c'�ћ�"O�p)��k�h}1靤O�ȥ"O�m��♄XT|�q�Ϊzy��"O �qϯo#� R	ôY�N�h�"Oʍb��R���dF��@�WD�<��۠,��yR��Y�:s�ia�S�<A"����L�sV��oo~ 9a%y�<)�@d�̝���	%(����k�<�g��5p-���̄bb��C��m�<�B���������B�l��OA�<���x) �AuZ�Kg�S�׊C䉪,4��@ǫ�;
���%�n�LC䉀-Wʀ��,� ��Q�ÐQ�XC�	�W��T�t��+S�6�U��*�2C�$'O�p�6�޵|ལ�%��`�lB�	#����$�K4�n�S�R�}-C�	8��a�����"�n��>C��5�I�(@-z]X=#U+lm$C�.9�n� `�#@��螑5fC��p�������h�0���[�*lC�	&;�`!9Bd�9����G�g C�	�+��m���X�"L�g 8ww�B�	`�v�+B��{�V@Ӱ@�5��B�	�l�B���FY%4td����H�z�\B�<Mf\Q��b�+�*�(u� B�I��4��h�:��D����3N�LB�	)��5��4M\�g*Ӭ6>B�ɿ��!j�/z0��Qm�/w"B�~Vx��.Y�VLQA阐4`�C��2�lT�I�Rw��E->?��C��2m�̙��o[�p��L�.m�B�I�pm�I"���4��%+��+��C�	'$��2mM�/��j�b�E!�Dɧ/mR��/�1_�R�Ͳ	'!�[�Eފ�12&J�LY�(SR
!�Ͱ�BsI�xԤP�BDצ�!���
��%Dޡ\��l����j�!�� �+�ł9T��7K��`,��"O��c5��
_�XkKĶ+T.���"OV���:��gOX;y���P"O��[���D� �s��P|��:�"O���g-�Y�Lq��[�~J=��"OI٢ː�RD6�A$E�!_L��"Of���C�ڭ�%S�W<��'"O`,J���?C��EX7oЩ}�8�"O�� � 㪍�٘��p"O^�k�j�&l#xy7M�'_�V\+D"O0�J�&(�����>:��Eð"O�P��O�t����ʼ#w  Q�"O��8���Y���c��W�h�&	ٳ"O
�����?It`Ƀ��*Y#�5��"O���C�� lvA�� K�����Q"O1�cgïTR���υ� .L��"O�m0E�ض�Ό��-	!x�^ec "O~h��k,��0��l����X��"OPQR@'E#��(���c���z"O�A2���<b ��F+�k�"O6�c�Y�M9��cC3W��}�`"O���w58��ZB�ؿh�Zy�"Ojq�����7�˽{��}�5"O�,��%9|
h
6C�%���C�"Od���E��z�.�Q�B�~��(�"O@@ "ǯ-jyq�C�&O���:!"O����
Z�@���W)�5Rք��"O��H�.�ҵ��ы9Ȁ�Ѧ"O�� 
�1Y�Lt�f w�P�[!"O��f̍|�D�pT\ A]���"O��z�BϜYV�@dC�� \���5"O�+����L��t����du���"O������	DL[�Q�f8"O�ұ�S�c�$mk+�Jr"OR�{��C�S��-���N)���"OXŸ�
�2�	C�
Cp����"O�8C�&C�:!�҉"{�@SU"O4��F�t���@ޤa �a�"OR�SbG��Y���ҠNR�aG*�"O����`M�t����N_8:/`�"O����!�p���i����<���W"O�H��/Ϥ�YVd��� �R"O"qJDIʖ/UX��%��]���"O�I���*�Aƈ9��9"OX�1ui�-�u��a3޼�"O4yC�Cu3N���훟;D�Q�"O�-�#A^oU����L׿DQ���"O,�(ԵR��$AA�(s��Ȁ�"Ot�s,�Iˆ (W�Ŷ>��[""O��*ܳhv��&��I����G"O�$S�i_=��( %ϔ��5H�"O��ywm݄o��T)U���N���a "Ohm����H�֜��c:,����"O� ��.Œb�j]SȈ77�1�"OvF�Ӫ}Q����M(�ȉз"O��8v�
�^���ك$��X��"O�9���X� 33B�/X_`iA"O�A�wi�5��C���]qz��"O��;G�.a��,)& X/;SZH��"O�t��aY8!C ��MW�P&�4@�"O�$1�B�]Qz�;��S5#�x��"OlL��!ZA"�Q�4#"��"OQ�����.�t(��`�"��`d"O;M��M�����N	���җ"O� z} ��q�t�p�N�>����"OV}r��Րg*���◀H.��'�a�fH3v��ӯ<H8��	�'x�zTጥB�Ŭ�o�J (�'��bvK��f�&�BE!�#q��)	�'�VhPp��>)���3�����'�vU�e]"=c��"�Т)h�|��'������ɖ0�R�sc��<5@�'y�|Q�hɐ.%�
2!<%D����'��W������Ra*�k��c�'�J����P�|&��;�iȸi+4���'b�<�CKG�<x���	_�@	��'\<��3���i�
��+�10����'b���NO�pRԇ��vqnA��'J\Sd�   ��U�b�O�hw %B�'AĠB�b�td�0����[�����'��L�`<qi�N�L͚�'��C��FQ�b��фĆ>"�
�'�j�YD��H�p��V''Rl��'k����M�%Yz���%Z�/��-�'�Ƅ�3�ڿC�0���iL&<�*�0�'f���0	P>~��C'b!7զB�'���#��ތ$0ԛ�k��D�0�
�'��u����kB�}����/��E�	�'�(�X��L0J<�1��fC"p��1�
�'	�yD	Poܼ;c�@�er.���'Ϣ X�那D��5��GJ=Y>ള�'t=���4D�R!��*U3~���'6�H;"IJ�W�p��b��[� x
�'����Z���+��]��ȡ�'�Hy��X�C�n��vI�+V�4ѣ
˓�(OL� � AD�>M�$�	n�H��"O�M+��ʧ��5�bq	S���y���0�`1���E&�d���R��yb�O("��2C �|]z2����'da{�@�,�4KM�q�b����'��D/�Sܧ�y-�(!0^!I����d;^��bnP��y��Z�Y�zE@�/^|| ���ڋ�O���ڈG�-`v���Z|[���d6!�!G�y��D�9'��H�a��0��'+�|�Î�:�( �W�I�<�*��`�Z��p>)J<abkQʾ9� �R�,�(�w�<�6�	 _eJ�ʐ �[e
ZO�5l�=��_�(p���S�\M󐀈5xUɓ%D�4I���dP�	�#Ǳv���S�$lO��`sRFA;dٓ�ƙ^� �"D���t��h��4�PƉ�.D��{`�t��Gz��ӛvJ�1�v�J��-"�QA:^���:���Cz��g�2R#��8�i�'���hO�\y�����rK@�Qa�D\6yF"O�I1�ůA���ܻf\< 4"O���!.ަGo���e���m�����x�'(^�H�bR�
���cw��7�xy	�'nLE��	�Q^8DX'O�*��\��'�>�#O�:���f�� +|����'K.���]"G8���_&Lh�ab�'�n%c��/8�tC���=SRi��'Iڐ�#O�6���85�U�6�BtI�'�D�@��_�}m`I]+���
�'��7#�P�Gʒk�b�8�'�0��S��61� h�Q��/jNa{�'���SL��6�pe�tDM�C8i��'�\%"0��,F0��(�l�I�2=@�'SL��+Q'W
�bsJ�7<�x�	��� 8����d�VH��nf�)p"O�DҴEƹo��@QeN� Z<�pX#"O$ t�^G(�	M�b��*��'���n?"L�$�	��@�bwV8H��Lğ Kr�'�{R.Z3#�Όug�!0����'Bf��D�į{Q�h@U�F�&�j�B�}��'���F��?rȐx7䖭������6}b��d�O��Y2r`��c�,c� �F#�4�Px���Ub@ �:��)@n��(O��)�'���P�� �Dcȝ1�E�	z����P�2��U-_�W�Ϣz$1ҋ�$?�g?A���bd�h[���/+Xj��"̈y�<	��G;Tu
t��(6|PuP��|�<�ϸ�U9# ��~s&ESu�<�5��|��+��@ GVQ�.�n�<1i�T��i�&O%pT��.Cm�<���\�C���C ��r�D�S�<1�MY<+Q����`�s����MJ�<����<򨹉ԮH.R��H��� (
~C�I�R��)�ϔ7?�$�I��B䉶?"T��ᝪU��A��<��C�I�/���:�	�%ܲ|���C��C�Tmj��y�r�8�ȅ�7tC䉀�
�����R@ʍHx0[�"O`��u�_i>M�r���n	6�� <O"�=E�ć�q��{a��&ZZyqT�S��y�/E�r#X��lI�a:�Q7eҦ�y�J@&�bd���M�z`�`!�ިO��x�O�,�P�o�9�v�)����'�l��'Vy0卆�>3��+Ư�k�(x�'R��2M	F].2�� h�p��'l�����-��M�Ԧ+`����'5�=���L���AĎŇX��Ek
�'\��!�ԦY��QvEB&H�0��'�ļ��/[:[L��R��"l�D{�'�Pp�Q7+K�(��ęQ��'�a"		Qa@i�'l^��A����ē�p>2�S�'�(�Z&��
��q���_�<	��ɰ9Ѵ� cD�h)��\�<ɁNζv`��R	� h�)�r�c�<q��*2.� �͏;?ݚ�{¬t�<AfH���P�&��8k�j@X6�n��hO1���:�A�9,b!i�lU:e�QQE"O�a�(R.VH��ʀ�A�����8�S��yB�,>�>��6�K9!W���CKò�y���;�pp�uM�e�\89�ʐ�y"�+a(q�%X�`���dG��y�
΋c�H��%�v���&�yr�Zb,�"���lD�uCΆ��O&O�b>�rQ)Y;�ع3�v�i�d5D�x�7�O�V��aඌ]]&���1D�s��jO��ŏN��*��*D�H�S��_�P��SjF#])��-�I[���� �^��oX�u��y���'�B䉢Y^ih��S�%cF(��B䉾zk<��b�PƎ��!$�4W�B�	x*��U��<#��1ĨP=zn�B��-jp�D��t���*թ�1?�C���p�c U+f�\�4 �+�����.�	� ���"sP�8��fM	c�B�	�K�j] T������a��e^���Ĉ/��'D��Ad�N�Pt�hb�\ށ�
�'�~�t'��'��U s�]1	���ə' �O��S�O��� ���d0\XZ"
�X�ܰZ��� ����ȓ#@�Q�A�R�}�V�g�s?�S�=�T>�<Qe&�{��*��A��
�QT�R^�<Q�&3��UawK�_,|PY&a�\�D�O��'��S�%D�H Rq�5l��P�S#�z?�B䉐3�&����K��Xð�E=HʔB�	:z�@�ZՂ��Hb�bn�?[G���+�ɳ5F�#Ôh��B1z�d"<)�1р�H&'�����r��(a,V��+�r����T��l�#�W�Sĺ=�ȓ�*��`�ZQ��}��`�3Sb0�ȓu�̝�I�n0�뚣e�9�=1��D2�	�Z�Έb�c]�����%K�[�!�׿?x0�A�K	&rV��vdX�P�v�)���F�'S��p���'�dP�E��>A�`Kčp2팝c{��R���ȅ�w�FK�)E�U��8HL?H����
`؁2 ��J'&\����a�~�'ɛ&�$��O�4�ɢ-E;_����1�_�o2�A�'(���fY $��J�(N3��\�4�hO?7��8o�Y�Ѕˋ ���)`�Fq!�$fj��p��P�L�p�Re�i!��#G���IÁK����a��8B!�@>q��ڄ�u�JDz�ݹ@!�d�_�4Y���^�eyt�j 散X�!�$ըb������97_��胅�	O�!��,�~ �RM�uEhݑ�N�8!�䝹eJ� �b� �v/�AQ�Q$t.!�D��^:��:�d�(�L�����!��ֽ$"��5LTX�.Z�-Rp�!�$Z�d,������rB$�5�P�u!�_�:��t�5m�����m֪(�!�$ӗ2֌�d���A�nسq�ٌ.�!򄀆V��1f-S$`ʰ���Ȕ.!��<7>� �J�q�6)����?-!�DU�~��*4ʀ�z�D
K!�DQ*(-��	RS#DȈ�r�䌼h�!�J�\�� s&ŉ?�D}��W`!�䊺x�<�Y�o	}����q�@�d�!�$���r���-��q�M�*a�!���+Z����&f�2f�|�`m��"�!�$�$[�.��f��!�ep��5n�!�D���p�$�0$ݦ���Nƪ$�!�d�([Ɏ��f�/6��h��H�h{!�D�>F����D��Єy���!��T�N��Q�o�>x���2��>`�!�ƺ_2)�S�g3�l��c��u�!��T+��c����:zQل�#d[!�d�('Ҍ�7c�-{�=�U�[5%G!�X9�Ȍ�"(�*y�r���A��\P!򤁢8����#�\���A0�R�2l!��j&�� ef�[:���B�|!��^F�@��-1��"�,Y�{�!��A�B#�طe� �4f�!��EK���ABE/v��!'�G�R!�4i��m�Î�Y��&RX	1�'��`@ED�0(��ߠ#)�Xi"O��qggѼGSj�+��� Tq�(ZW"Oh8rIY�T�f����7]
��?O�)0列9:!�L #E��v-@��Z�!�TI̹_=4T;Pk��n�zC�	{�@����W� ���ā2�C䉃Vc�\��/ݕ���1)�$vC�	�c�JL��"ԕk���Q��/)��C䉟(�Ɛ�6�H�,S8U� wifC�x�#���&�P�g�*:��B�)� ��[�B�6)�Q ��^�mʜ9��"O�\3!�'_n"Tڃ�Ĵ+|tٶ"O	��h��=8��slÌ<�y�D"O\t(�@�O�z!q+�I�|��"O���⅒ �XH�׊'��)R"O�9��p�ʰ��mU����"O��R�Sk�V�V�FO�AB2"O��B�B�O���h7�D0u=�9+�"O����C��䒗�D8��#�"O~��7	�$&���>w�,�#"O��[���8P�H�1�%B���:�"Oh1�F��D�x(��>]G�<�U"O ��FI�7R'�T[q�(���{�"O���r�^�J�n0[a�ȟ5x΄�u"O�(!#�4��̀fj��*x*�"O8"�*�(=D�%k�CC���2�"O���I�!�8��[�Z\�% �"O2�':��}���*_x1v"O�x���
,)�B͛�j�h:�
�"OtdŰ8�����W"F����"Oޝ���5V�`���+�,�'"O�sф�d��+M�C��b�"O�h
d�-w�"��#�~�X$"OnI�Q㘪M�z���]�k�"O�a�GBH�Lyu�ڭ>�P8��"O��!w"�=!@�Ay���zӘ�0�"O��8�F�	/`\���F/M���	�"O���F��.Zu\��"��~���B"O��a1 ����$lV�E�:�85"O&���� 2h��Pn�G��]�"O:��5���<N̽c�-�"J�I"O��L����`�R&�_���[E�&D���KX=_0�\������E1�$D�\�e]�5̵ GiX�-���5m%D��yS �+�L	�A[�.@�90"D�<��� 
o�U@��L�%GTț4� D��J��;G��K��M�&���y��-D����e�5� XSd�9g��yH �-D�������EǨ���T �d��*+D����ó2}*0��l�%�L))bK,D�4���l��"�M]&~|��)D��;b��K���S��q d�;D���ԏ�6+��l�A��o���[��6D���e���7~݈�d�#�i c�3D�0h
L�Y=΁S����}$��e�.D�[�ME�`�hك!!�<Q܌;�*O��	� a��X��C�&�"L)s"O�ũhry��@�0`�"Ё�"O��U�M'G�%.ħ7$�7"OұA�]�8�e���X�D����"O�M�VOEG:���1�1w�0H"OV�S1�F5y�ٗe�9�6H��"OT%� ��4z�Ȅ��$I&!�0��"O��W�,Z�xJBS�X<ziZ5"Ot�D+Ú/iB�ɠ��bͰa"O^�ic�we�R�e@�E��q��"O0l%���`qjS�ۗu�"O���v��x��`@�<,�nm�"O\ܺO�-0b�Ca�7nQ�D"O��ڇ��k^�����%dd���"O�������9!jү�z���"O|=�0^{�}q�	���"��Q"OФ��`F70�f�T��#��ԋ"O�!ɲ��^%�&D�.�P��"O� �2�i���±�`�Ǥ/�hpS�"O��I�m���� ��	bʦ���"O� ��

p�>-�g�ޘtt�j""O�EK�'<�Z 
��=SRF"O��1�%@�oV�%Sq�fB�D��"Oi���G<{|<� rɒ�RC ���"Oڝ�d�+� �۲�ͱfU��kc"OXtY`��!r&�t��M�)P���"O�K@_�B���r��	�`�1"O(�S�.fMf-����
��'"OL�c�G�56����ՊC L�"O0���ܸv��h ��04^%�R�[�) P�,�.�12ȝ8�E�� � ����/�O�U gY��?�qG��	D|䱰O����ҢJG�<� @��jL@���L����aBj�'�^UX�'�u�O$�z ɏ-+@�@h�셅v���j
�'<xy��Z�sF`����w�,u��4M�d��#�)��}J�m^#{�N��v��^ߨ��%D�,�AV�j�6��7�U������O�>i��־�l���4.�
���5&!xW�"�a}���G��Ie��
L4 T��h�M�C�	�Ȍ�ӂ�ר?�F��C�V�jiB�=1��2∟�8��ȴv�V�{�
�.�޸#��'��t���{}�cל2�:�a&��#AM||�(��ybbS�uO����	IP`Ѱ�`�1��'�l�@��X����G����'�*�P�'�G�P����y�,S�����&��)7�4����:�1L,nCL�ɮ>����O�����<aج�R��Pa��H��O�(+���G��h���4~P��C�+,:T��'��T]�E�'�/\O�H��a�${6�"̀>E�����'�j ��~�`}QU$I�(0T�d��:V�L]���ܻ0Wp�)�3D�\�A�E�_�ڸʵ�]�J�PA�RF3}�+�f���v���o3$����[�O�
N*||S�/Z&M-,X(�'\0{�g����
�*�@�&��U%��"s�k �A�A�f�(d��(ڸ����J��T����b��y�pT����"D�ǰ?_fP��($4 ᑆ�@3Ach(�CǧN�R\r#`����<U�&/"y�K��R]|Xɡ�On��`Qi�\{P��"C�@tb��l)8�Bx��E��<I$�R�fN�����0�����jA �_:��?��U��l�h̓���{��ˉ�t�ΐ6�"Tz2*N�`�
�ɓ����yRkٟ �8m�R�ړ5i��HJL���y��R�.�-A��@ M��,�����|�KΥXg�Y��#;xu�Y=�C���8�hB��+�LH�V�T����B�  �ȉJ�N�!z�ai�Jx�qq,N�����oյO����P�-OX� g��x��MZǧ�d��&�>�~��P·�>�����)��h�.C���	�1�
0|B>-qpC�:�f�`��hj���-~0�h35"= Q	����'ouUF��T��"��/�y�F]\�T8���\�O��L �b�.	f���UHD8�y�p+��҈�L>�&
�(0���j*��q+eR|(<%��L��d0��1^���k�6�(��tLO�ێQ�qC��x�d��d�Τ���Ω����ט}	ay"�ϜQ(��G*ծ2��`p���R-�U�� K�%�T�+PFܦy��B�	'S
�� ��,]� ,�Ҧ��j�pOI@�%�I�2���!1"�|r���j�5i�)��v�,��pF�<��!�'wS����Q$  ��I3H��-�lR���d�@9��?�'�@��G�߷b;��+��(�uH�'������O�g_z1��G�	_Tj��6��yY�b��#�0>� N�B��y�,���:d�Pv�����\/C��	���,���N�z)r$�����"Ot�'l�9Q��$Ӗ��"�U�t"Otp:KT�&���%FD�"O�Q�ff��+��X���g���b�"OM��-ިkB	��쑏	�Љ"O
�q�����t��0+�0)�4�t"O� ��2�ߡk��UӰ�U(}���X"O�M�^.~�f�`��ĺ6"O8IQr��;d.8= ŪR��i�"O�b��i�`%O� ?	2�T"O��ñ@ܤ-�R0�c�,\#�"O\��c�'J�=�Pㄵl\�|��"ONh����w��R���?w�(���"OZJV�A�����Kſ<�B���"O����a�o?�'#�[��0�"O�y���*d����3�B��h�"OXh[�M'�p�#.Z"|�0Q�"O.����c�L�WMJDRv��"O0����Z=<tI�.��6��Ī�"OB](�Ń=LvlX�1,�-uT�"O����̇$�x�3�_$ې���"O�!5�@�^�P��D�p� ]�"O����/�xg���K�h�s "OH 1C�D�<0���N-��Pk�"O�dXuCR4^�#sAE*�BM��"OR��P�� Rv��f���r�8�"O�Y��o��y���p�
d���z�"O���S�N�}��p;���M����"O����CP8Z�Tc�L7z��W"OԀ�4��00�h���qZ~U�"O�lJ*5_�0���E%`@��S"OB�{b�S&�t᳑���	0@5��"OT,��X3l�I�fe�Ȳ���"OZQ�׈%�(pjb�G����Zp"O��sbN[���Z\��'"O�� �N�&�iV��=d���	��'�!�D�<X1ν��aֵ6�4�:��^;Y��{��ƕ?�tѺ$#�:R
r�Cr�Q;�!�D��c85��P�<����B�C��OX�=���E��!l"؊mZ�tv��b"O�pŠ�/n�H�U�Ӛ���"O����ΧB�&���CX1�,�x7"O����\�)5��Qd�H5m�`= �"O�I���T4��C�Z�c����'"Oz8��*]:ݒ�9f,���m�S"O �����9�t�CD)�l���+�"O|ݒ��Ib���Ў*�;rO��k�gO5��9�dh��R���V,F�P����I�d"El���g�S:Q��?VZ�(�HF���*�R�<QT�L�I=~��An�$3�BR�b�<���4m!�3�־U��	A�v�<qv#��}�4A&�5Tld1��Ir�<�-�v���Hր߬b�R,c�eQ�<��[�ym��d<%����M�<Y�L�g����s%L�-l��F��E�<Y���Lu+�G]m��sec	C�<��l7Df��q���% �@p�A�D�<��#�za�H2� VȒQ�V�|�<	�&O�[�i��׌_�H�"0'Ft�<��D�b�0��c#��Y�t�X�<�� lD좲�N	H��PrĊT�<���[-B��@
�O������z�<񴏂�\F���͸^l��!x�<Y&��/E������7�.=��+�L�<�띛�@x�Qk�8}��X#q)SS�<�s�#���r�'�;/�r�w	�M�<a�H {��X+���0��@����K�<I��G����oW70hF�9c��C�<�&L�O��8�	�f����q~�<���eL�<�p+�-?0�ۓiAP�<� �B%�wD�,Bt�"�.DH�"O%xf�ϓz�D�C�I�g���s"O������Zxj���KwԈ
�"O|�ˇ�]4t���E�4��e��"O��
�@Z=�,����?R��"O��vF�0n��3��W��ucc"O �@D��#) ��A�A�p�8M�!"O�h��;v<4$�	}��lk4"OBA�4f��ULxD���&�j���"O�1����L����_4l
�R�"O��0OrI�p#@ַn�����"OBт��/���qOC,qk����"O�F��)4�+�.9oR(��"O^y�A�]O4��IW�M`I ��A"Ol�*�)� O/f�� n$���"O�HZ�)[�L��=	dN�6j�����"O(5z0��n����N���]`5"OxѥgZ$n�hu�X�i"�Ö"OZ�3UB
T�����R(KM��0�"O���V��2d/�͘`�_�P�ޑ�"O�5h�D�R�tĈ �=q��0�v"OJ	��/%���CȆ�nLiR"O�ੱi��-����6&C��й:	�'R�� ��ܨ k���.?ъ���'��4D��5еJ��U*�ܤ��'ɰݫІ��*����`��Y�'�|�a��ta�@�:��)�f�E��y�Ԓ{��P�p!�4mv,kG��yݖer�S�*T\�5���y�Lٳz��-[3ԍ4��}�7�A��y�Kgh���Ș�k8��2����y�-��NNc�FܒMy�q�gK��ybKʶ.?��FS�A�|�щ�'�y���	�L���E���`�a���yb��6S� �B�,Z�weH��y�Dߦ`b��D`ӆprf��#U��y�gH�(r
�!�E(c�p�M���y��Vj:u�r⑚k�Z��7A[��yR&�<W�lX���(e@ƅ��Z��yRGܽv��왥Oאo�j�V��y��~��A���Y*�X�ֈ��y�׮Ae�aE	I�`+�E�Uϝ&�y2�Λ\����c�P<o��35��y���f��z� c�ػ�F ��y���\9Q�BįJ��)jt����y��!
'DQh�D�;9��������y�aT;L����F '&�����y�]$j��A�C���#���yb�õ>&�� �'Z�6� ���yr�Y�Y~+�@ڸU�"𫷭�(�y"�4p~�8Aj�7e��@S2�y���,�H�l@6z/��`�l�)�y�N +��u�$�R�h�PD	A���y��&�,ʔ	 S�L�`�܅�y���$����4lGM����[�yR�� �ްJ4��g<��Gc��y' �Q
"!�£��Z�y����y�d�F����
���U��(�!�y"L�
=��!�`/؋r�����yRf��D�| *�O�/u�칲�MN��yR	!&��R����f���@P��y��}�l���~ؤ��E5�yR�X*8��Y��!?�H�$�!�y��X�L�p��#萀!�����y
� ��Aׯ�"S�y�����fU["O��B��G�W6X��r�>���C��h�<ِ�@�tӜMRT� W�
����b�<�	,��t�$���5x�"�t�<�$�]1Z�R���'�e�v :p�<�����8�!h�Cf�,�@�Vp�<��K�7�T�P6*2�qa��[�<�A��,<�i1�S;���@Y�<�"%�x�ܨ�IƒFej�,[�<I���Z -���N.�ݫP��R�<y�(H0������qp�p���A{�<)0�9	
P	cV��%c��E�n�{�<�g�ɔw-,��!Lҥd���Y@kFr�<�ѧ�>UVt)��T��i1�QP�<��UG����UI���M�<�UL��3@��$3z����J�<)V'U�O
�!�όm��J�<q�M�C��7��A�8J��n�<qՂK	OX~��'��Q�M9���V�<e#�z3p�E_509q�$U{�<�W)H2게�#Y� q
]9'��c�<х�O�CȰ��bI�:K�mYs#�F�<��%56�|x��DjX�h����F�<ѓ-�>�r���Y��ȀB��j�<�@o�%P���#��l>f����a�<�F$�	&+H�4M��k��{!�B�I< &RѪ���1���A�M4c�B�	��q&P^��Z�l�:��B�	qѤqi��c�
���ƆQ��B�qN������G�����Į ��B�	WlJh��L�P��#��.#�BB�	�D`4��kR�g4�D�m� �vB�ɶ"��"��q���B��#aB�I�V���BfJ�=l�BS�:��B�	55����E�v.�ԫ�*�vB�ɵ^w�˶ň:�X ͈/�nB�	�i�P��&�
�d	HvF�C䉎��Z�������	1F/;ZC��?s!����.I�O��u	0.I�FY�C��
c ȁ c׊O�Dĳ���wC�I	C9��"I�4y�^ԓ��
�9��C�I��Lq����E�
*w�Hd��C�	���0E�<���R���$�Y��'A�q��5D�Z]b@�l}[�'�`$���(_H�]��K�@tj�'�]:��ޞ!qr80���KVJ�9�'�Јy�+�'�T�5��E1�y�'x\@FO�8C����N��I��'�P�"�Ĝp;�V*Ө=�x�
�'-8=[@C�$nT��*6-�-�	�'�ٙVˎ�e�E+ Z7(4}�'���G�D�V>�؃�.T�$�����'�.��s��&.�)Ї*�:i��'>f���HL-m��S��>�,�
�'<,p�V�9W�U���[��� 1
�'��8����/ƀ1��/8��i
�'N�����M��T��ϙ&4�l��
�'l.�D��_�\�S��V�W���'D4A%�(0��@��y����'L�1��ϱN�@S��uH5��'a��*SMǀn=Lx�)�b��P�'�pi)5h�?x%z�@c�ĴY��U0
�'hZš���]`|y;"��Z��,Y
�')��a,� %����1���Q�@i��� �uX0E�?x��HpQ[����@"O\z!�ς3�p��zsJ�2�"O��r��D�z4�B o֎e����"O���+����'o5R���"O:d�o�*�����E�J�tҕ"O�h0��t�tH�Ō�i�"O�@swO� Ee
��d�-k�"OX@Q�gΡZH�X��N�Q�!!�"O�Ȳ2jF%bz�����r$(5"O�|QCc"s�Z�q�f^�a\r�س"Oh#rkJ�?���Y��	�;��L�T"O�U
���/Y�$+Վ]8qzQ��"O8�봢Y>(�V�Ӗ���"O�۔C�!+���2`�'/r�2�"O�)�#M�]���ǁ iD1S�"O8�����QjOl6a��"O�=���F�V�dX���։�NAf"O,0�lܾsr�J&
׮t`(��"O0CES.f��7iچ4HB��t"O�AFBCZ��JdIEN2*M�g"O��y�b��H�Ԑ��6I�1��"O�e��ǃ)���H��2:0��"O��qV E+�)vY"4D�D�T"O�Ȃ��] M�B���π76��A"O�A1riؽS=fL+�`�9u���"O!X`�YA3p%b�Nf|�bF"OFb���`���V	����#"O�P����=�ؓ��<-�-j�"O�h�V��C$��&F��V�8B"O�Ms&�V��Jeąe��H2"O�I@���Q�R��([;R���f"O Y:p�\�eY��bG��-C��D"O�d�F艔!�E+5CQ1%>�L#4"Ox1c�ͤ��l��Z�B"O���֫QF �I5�қ>�ѫ�"O�a�I���,�`��T��S#"O��3#�>gs�5±c�,�z"O�\�gԷQ<�p����V����"OL���/��L��;l��91"OD�a֋�:Kݢ�[��8�ڠ��"Or��4���b^�"t��Ie�(Ce"OB��A�"/��pă\�4�����"O�%i���Xfy��e߮^��嘔"O���3E�sw�	��V&9�m��"OxΚ{�mG��=;,ꍂ!"O\� ����$�UcYZ�B�"O޹B�e�^�V�r5lˇj�`B�"OH\�5��
�TkP��$���"O��H!�ŬG���1��Q�y�""OP�����V5�a���52��"O�p�g��Lq��&$�&1��i
"O�)����sv
��sÎ1U��Tʄ"O���1ۀ2$��;��B�p�,�1�"O�\Q��P�8�8ѿKblIX"O�h����Z��B�E�*0q�X�""OL�*��@�J�{S��ptj`8"O�]j4D �r�����DA 	dD�yE"O�x�GbS�HQ\��^e]r�!b"O�����F��ayf�M]�<��"O@�c��� l�Ԁ[�®d�Ƚ�"O4���EǶr� ă��6oժS�"Ox�����ʔ!�y(F�`"O2	B*�o�6�#�"_�m:$@�"Ol|��̕�`ڝ1��;�4]�"O� zIӰ��U �]:u�\L��"O�%����?p�L����6L̢�`�5O��s�H�8e�U�$�[	!P��59��M��I�Q/����hj��ҒA��(O���R-���³l����U�M'hw,b��j��)񉗖qД�L�l?�t�$0AZ�'�~�Ey����%)����ժP!o���Q)����\.�(O�>=1DH�)F�����2�d%|�
)0��)�'d�lr!��D@x�fI�"��TK�D��uw��?�$�p.\p�0�B�q���K>� q��O�e.����H��4�R89e�p�dIɊ.�	$I���)������S"��T�	r�^\zsbF>*~R��F�?)W΅%7&d�J>E�h[![iV�$ [�Z�*����X����F����0|��+J�?��+�کL�.=*#�I����'�8"3�	�|���9��(��
�5����Z�gO �`2�"�BX��O�(9{IF��d��.B���y�I]�@��� ��L�B�|�у�(��F�ud���L�?�|b��D�0���D�ՠc�) 5������ݎJ�\	&��~j�Қ�N��a	:���K��46�.��Pϔp�t>9Z���qȭXU$�;$��+�#%��O ��|>�~�O}���C�#�Eä(J5Oy�e��'+}�ij����P�~�]>�M�DйQ�8"h�1BpIàj��d�'EҴc��2�)§91����[����	��[�e� �����Dx���H'��Q�@���J��L>E:��d�z��ȟ��SJM�?\B�IU8fH�L0�k.ʓ#�a�D��(~���3%��H��N����'B��GyJ|z�%��.�4�Ӗ��H��(��J��;.Q�b?y��AًQkl:�"O��t.�>Q�4�O�	�D� s��O8,32oB4c�*) 4N� �
��[f�<)2��f�jiB��ɋ\�t
 G�<���PNU\�bŢW!-�@�"��F�<������jPk�*���sYX�<A��پO�R�*�
Ln�*T��g�R�<�����x�x�ҍ�(�s��K�<ig�J�Q<2�CRg�3GA����C�M�<��f$cb�$����0g)�iS��t�<��Ą�^������/�*l��a�G�<�g��x`Lh�'�������J�<��(�����
<� �AÌq�<��$��?A���6�S�X�R��ѯ�a�<���Oh�&��$�׳i����!F�\�<	eO[�vKT��%C.@�Ή��g�A�<��G��W@�j��(a�~�J�b�r�<	�M�!��&=�6�FjXe�<���L�RH���D%u�H��0aQi�<��m\�3����fe �fje��O�h�<Q�K�N �1��`��b�HD��*�c�<� n
�3�l���A�8Z�6����U�<Y�$0�x��!1��J��NF�<�ch��4Z&�F�T(����A�<Q�K�M���BiC�C���c�Dt�<Y��T/+��������H�M!!Kt�<YF"Ξ1D�y�F-
+4���`A�o�<��¾;o�U��&�P�|�2��l�<�$]^�m[@�)K�n�v/If�<����`��*w���Ԣ9�,T���V3$����A|M��(D����U����I Ӡ��D&D�  �gǦ[`�8��O1���B1D�<@��ϓP����I<5zrz�j/D�C7��/0,2M��.04��,6�-D��6@T!k�rI�#Ӭٚ@W�*D����͆d>P�@WBP��8|3sO6D�4��ܮF��L8�f���Җ��!���W�Ҥb���T¨���dP	"�!�d��D��ٙM�&�j�,T"�!�� ����98q$�2@B:�t!p"O�4���[�b��tf��ghPؑ�"OzH���e^H����5J��Ȃ"O(����(6Y)�"��Rd�@�P"OR�{�nI�_q�@ :.Y��
g"O�51I��R���v [4s@0hq"OL�g ��[�񖌇�k`�!Ё"Of�)�ʚQ>�@���W=rp<ڵ"O�x�2�X�9�H��D� Vp|tr�"O��3��G�	R�D�D� �
�E��"O��3�� �Ny��������"O���ԧ�<�<�� ���8���"On�g���^���*��UQ"O�׌H$%2ykAG�.����"Ol���ӇL�E����d�P�.�yri�{p��zvk
�3�\XP�8�y!�1���D�N�+��U �����y�� �_BqJ�Gµm]��q���y�BB.C`M��K��f\ڭm�:�y���#a,i(U���tc���yY�[L�3G�(\�L}��J4�y�%�����Q'OUĈ�b���y�e۽DT� ���!L�#�*L��y�Q��<H7.Sh��������yRB̰\�8�`�E&d�x5(�鞁�y��ߘ-j��Jsn/�������yc"5/����*�3&�� ����y�m�t'.���˜%XNu�@-S��y2�ΐ|��XƇ #
��+@fC��y�猶d=�x���Ԙ�$yrgY��y�o�2<�<AJW9H�t��	�%�y�j'_)�D0�iV"	?Z$����yë���㒽?�}ڐl�&�y�I�0]:1��%H�
�z�̈�yr�S�Ey����mL�	@g̕�y2lR1B�Y�F�
]=�q
Ј�y�H�'4	�5�Q�[pPA�%ڐ�y����kA� ��OP N���h�B���yK�oqX��/�XcL�����0�y��ғB���X�e�((8����y�ꈦQ�(�:W��9n |�
���y�jHT�d���X:�+����y�
![Є�f�YfVQ8�JϜ�y�'E sv�G&�"&������H��y�����89�ӎ�r4(�����y�fƍk���� R�|;����F��yb��+pI��ۤ(L�(܀��{J�M�ȓ-%r5��-��dDm{�fIZu������A�J�N�9P
��>��P�ȓz�2! I��zS��|t\��ȓF-�a�DA�u�V��FLJ�$�ȓ���(�(�= �Aa`�>�,q�ȓ�b!Rŵ7RI�Տ'&�p������؍{��p`ӉA~z����t��/�xi6���a��ư�ȓWQ��{��S)���"���A-
��}d<"TɃ5��к��"h���3/L-�Q�7Y�2��G�(����K�Ҩra�<Y����r�1g䀆ȓ7Ą|�+J�L쨚�,�x|����1�� ��HL�l k�ϟ�z�
����?/��C��.^�����z�<�p"�'>(��b�ք� m�)�y�<��U�gL�����:�� }�<� \LZևS�~��@�T����4"O���S�Kd�(�.ߢw��	��"OD����<F�л�B�W�08K�"O$�9C��G|P�� �C�x�Ĺɢ"O�衤��[����U,P6�97"OB��p�N
X\B�c��R�"Od4
�,<z�akQ�% iq�"OVT�q�߹X,@!��
Rl��R"O6ЉgE�rI�i�F'=4�hQ"O���S�S�F�!NL6%Ⱃ#"O��iơږuR�1Îƽje6��c"O91�^�2���y��ɥl6�`�"O�}�$��X;�Ђ��R��{u"O�c�6�|����Ӏ/+Ρr@"O�����/z��U�ܟmL+2"O�A@G��tNz����#�$0"OF��J[S�.�!D쌊�ļ[�"O��[f�%I�,�pu+�!3��!�"O��R̄�I���3�S�z�21qc"O�r���0~�� nܨK�,��"O��"�
�M9`%���
�.K�1(1"O,�ӡN��"��G��+��t�@"O��hR/�|�*���(|Y�"O�9����uIȠ�����K_�Q�"O���a�9T��`�%�ȃXQ6�:�"O~���i�hHY�SGJ4y�4��"Oԅj�.�s|�����w��P�C"O,��p���\p��ꚰU��C"O0��V�K�:r��A���
9�!��$R�Q ��6�.Xi1m��!�D��"j$�q�Q�QZ
lY"*9�!�䔺gø	z@/O)SQ� �ƫ��!��62HP4
'�&Gޘh�Jʘ�!�S}TX�3�K>zT�5�4XQ!��K�\M�����K�:9(Ш
	5!�Ě�F+�t* ��Z��%
�I<K!�D�!3R�mX��߂i0���!`J!�OD������lb��h �@�X�!��P�eM�HB�gЛK�F�qNД�!�ĘH	p����7�������mn!�dN( J�����U�ȁ
�{�!�dF=s�ZI�ʖ:�@ɰ��˯.h!�$�L�CѠ��y�(գ�&��xf!���Ed��,G���ѷ�F:1X!�D�7���2�`�.~��9�խ߻D!��Ƈ]�,8*�d�<�����+F!��ԡ{�hH(%h^&m�}!�U�a�!��P�M(���@ͅ;L_��Y4N̞&U!���1x���W�ЩeUε�n��mL!�� �, �_���h{��3-!��$t�H��'fL�skʹ�!�B�/�&�k���v!
����!!�:FR�`S�C E6r�Y�*N!� V=z�@4)�2? ��+�.K�!��9h�`�㔼3��0f��5o�!�D�1:��Є��"�Bq�\&Rv!�_*egxH 1`x��Y�!�$�DX��+ޜbBVu�K��E�!�d� ?�9Gf?8!b�/v�!�d��@[��AA��>z$訁�k�k!�dˠ<�X��f�J�����IJ�R�!�D*VK�E�w��:0���@�S	!򤘔4��؄�L ��ȵ��D��Y{�!p���r��U��I�(�y
� �Ys�$V�*`p! nՆttX	G"O�H@�mB�]c������5��5"O�hȠ+I�l�x�M4Wؠ��"O�M��C
�n���M5*� �2"Or�Q���6 6��r	6-�p�q�"OmRL��v�zI�h��.�CR"Or�`��T?L��P�&�4���P""Ot�#��	p��Yo�/ B���"O�ؑ�b��`��2�H͠���"O�I"�
@�5�T��M̡^ȋH�"On��"^�Y���Ӷ��Z�v�ش"O@��a�H���"��;_�N%[�"O�q�����,&Ľ[e`��qC�"O� �5��`L���E�W�F��a� "O��(�ΪD	L�0C���X�"O�� %Ũ4��L2�I#i:	�"O����6(�nA���#j��ڧ"O�9���R>��*�I��-a��h�"O�(��e٪��qrg(͐]WX�R"O��ʫD�P��p,>T
��C"OZ����-�VX��*_�R���z�"O����O'͆�˶�ʠ�l��%"O�x��ɞ ��I����X���1�"O��z����6��@e�(�a"O&���K�#�"=
s Ѯ`�X�pa"O��c`-C/)�T�jS	��bך���"O ��D�R�8��9�ȁ)F^�l�P"O���!� V��X����}�N��"O�I!�Ʒ ������_6l�f"Ox��t��)NlVH9�kO+��a"O��C�A�]~��e��!}��D"O��	�   ��   �  �  �  ,   n+  7  B  LJ  +W  �c  �i  p  }v  �|   �  A�  ��  ƕ  
�  L�  ��  Ү  �  U�  ��  ��  i�  N�  ��  ��  ��  � g g �' �. @5 �; �>  Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�� |d��"O
`�(�;���8���-0��1%"Oj4��ND^[��"3/9�0|H�"OB���H��*�ʞRy=a"O�味V�!X��!&F�:J�$���"O,��a
���C�Ą�M�"O,$3%o�-���p���+Ն�:1"O��ݢ1����`���y14]2��i�<�6��{_���c�H�`�fX�$Kn�<��A̼VI�xR[�)�Ć�pඤ�ȓA5��('nߡ4�� �)˩%� ���,��r�؊b#`T�eT09���ȓ!�b��g��}�8�F��-? �ȓ
K|m�ș�VṔ���2�%�ȓ"R�X�j�4JN�1�˘X�i����̹	_�jZ��1!g��zܶ��ȓgil,*�J�
j�Ne��i�J%b���f	�(U��:���G��$Y^م�~r�� S�%T"���k\�jx�ȓ|4�1�îJb��@ӵ�ݩn�V��/[`�"�v4�R�!ʎ<��M�ȓ`:��z�ؚh�J�Z��$HY:	��H��p�m�C1��!��B:��0��EnjZA V;9����J[
2���	��4'J�EA�IVW&��~�(aZ��ӹ�>� o�Y�|�ȓ�f�A�
Ο7�H��M�$�����mޠP����/���ANXo*�ȓTv�����{ ��-7�*h��I��sB�8�8���3����ȓNe*M�悡;������X�o��!�ȓ'lj�#F�m�+R&;�|��2)n�C��0S4���T:
b���:�0!��e֊��)��ͷV��,�ȓ0�&�8#���� ع�L�����;�P�AFd���,w�6d��r�EQ�( �gVlɦ�M,H��,DP���|�I	$G#\���ȓ"�)���E�B	yt&B�^�LɅ�4�� ��eëF�ڙ��n��R�p�ȓp`@}bŇ�=�$�AUN��P����L��p���_�a�)�Y�!��-��u�5���o}�`iF�@A�p ��F�\�0��[���IF/5���k>bTؖ�;K'DT@%^��@�<a�>\OЭS��g 4�0C@�;nG"aq5O��D��S��Ѫ׮�J�fT�� ٗ&Ԅ,�ē������(#�|Cu�Cn��4��ɝ�HO��'R.
hh���^7���"OX��g��N�`��<=6$\["OR7+��	p<fl�/@V60
v�:D�t1���`)<���"��.��.4D�$0Ί/8�j��
Y�bd�v�%D��"�o�=W��X�J�;Q��	�&%ғ�hO�����G� t�Rc��%fC�I� ����x�.T�Pc�/z�C�ɵ��s�)���`��C�I8�V1I�l��9 �*���<�0B�	�bY
D?y��C�A/@3�"?���'��-��E�$��,��ɀ5fa�B�	J܈4��ɆS�~0��݂;���hO�>��@��;K2�9	��r��	�3�,D�� `�z����P��B�4V�- Ŕx��'�
���n˓|��x��E��n�FL���y���)Wp��WD��Ĝ��y�%�`���#BEV^)	�!�����hO��Q�&,j)�ԩ�7�6�!�j�N,��:O�H2f��,�j]y��׫8t���"ObX@w�ƺ*�rj&	O}�=�!"O�Xzp�
}d>yc���sk���"OJL2��5KԌ�bul�%��%i7"ODE���(!]�����[�M�����"O�R%��^lh����3E���#�	矤�'�j�>qQ'��=G�nE*`͕n��m�B D����Y$M2���K�)��!B�>��OleP� ?E��c�dߺ���X!f�{�*7�y�Z�e���J󉆫Vj���e.�����}�)��B*ԛ8&XX���B�H��i��N��y����9������v7�$Z��ã�y�bC�Pjq�e���q��r���*��=E��T@������{68#�mTS�l�ȓ@����@�R%���S�[�^��ȓ�(Mh��DT�Tc����R���G|r<��g^%��%� ΁�X:J0�ȓ:��!�O��xc�D�0��!��	>��'0�)���@]���x����'�l	F�&>4��&���5�I<a���a��uw��d`�yd�1
�R�)��@���=�yRA�{t�U&�#�0%R�	�!�D��(	��n�,�.�ٶ�؁Q��xr�I"���:�&�_�a'h��I��9�Ɠj@�XPQ�Թ4��t�3�������Z~�P�xy�i�4�ȲHX%��m����[X��)�	ܒ&B�8��T�V٘��3���l&���O����x!�b�����Ǔ�N^C���B��K�*h8�,Q�F�"=	Ǔv(����Њ|4��횕'�`L��m�������.����.ܚ2������z�Yb���U�Q�>��P�[3��d�&$�4it��;��(E��m+`%H�e���yr��]]�M��%+2��[$�����&�S�O��A냂L�-z�����1�0�'��U)J3o,B��@�Z%d�G8�S��?�OH��$��B ܊���V�<	a����E��9tP��'&L��M �@�r8n�;󇙥*��D�'�vPDy��	��(\�0J�K	��ӗ�e�}�<��^9 �¨���B*?�ى ,\A���=��Ƅ�U��8�j��~Jdq���s�<����.9��%
r��UbN�D�p�<y�i�j:t��B P�J[��vI�H�<I�_�O�����l��J��KC�<��㜉1��H�o�E)z�R�E�g�<�&)^< 0��撀n��׆Kd�<y2�!	Xv|��E־C>��!!e�<A�)�0ww�͡�/�n���`nAa�<��X:?������Wp� b��\f�<�DהY�I��`+q���S���L�<1�nې.*�4�#)J�<; �r�R�<���ʹ�0�B������F��h�[��)��l3��",������A�p���	>D�hI�M�5).��H��	Y��Q��O�?����Ȑ�HdrկW@�S3@Ak�!�D�D�mKr
X/�`�⑮�w�!��77xph��U阥�&��Z��TD{ʟ$��b��1?�U3�N��4O6��)� @E	VSn49i M��<f�}˷�0�8OtU�pC��� r�+B�,e(`�0�x��'��H�C&��c4J����I�H���!���Ĵ}a��O��U@$��WA*t�d�
�:;���
���K#�$|��+�=n��	v!Q�"|�q�Rx+6X��(�llV$��Cm�'���(�
�s�� �\E��ے`��t�`9OF��S<?x�
 �^&4MܬCW�D�zq��)Z�y��ʤŨ�`�F+a�!Rs�N,�yG<7U4�YWEW�Nȃg."�~��>����~�#d�>�~�u�9��8)��b�<��E3
vYs���o�^A1ot�'vaxrF ;���֠F$R�i�Kמ�HO�6�.�=�����!l�T� .@h�ȓ���c�2~P����9m�|��'^.�'��eS��)V=��D2��\�E) ���&����PyR�X
1��c�^5c �A!�F���%6�(�<y��d���P���W�y�ƍ)�C��bLa|B��`�$װ==\�� G�1�T�6��g=�'ў�>m�`��5tݚP�U�ޢ=i.�K@�'�I�{�Q��O#Π�����/a�́dd�!��%�	�'j�p�ALc�Z���/�	~�IJ޴�y��s���2�I3y�`��ǽoԘ��"O��h��#<>@�f��J��Դin����=�r�Ѽ8��mh�#T�/��훢�K����<�g�_	pp��e�aQ����ZF��hO�O.j��� �Vm�LZq)��~bRtӎ�<�S��̑�gL�%�_b��2$��y%K=T�R�Pԯ�o= (�V�S��y"&�
k���֎̝fR�q�F�́�yҨ�B�XM!W��/�0��5�A��y���/� xp���
�
���e���y�A�$�~�X�ҏ��FD6�y�트ew��"%#��}�J�c�ȟ,�y��ǭ� 41��y��}�����y�'xM�}�	�jYz���DL!�y�J�%��Q#
���I��E[��y,�S\tBD�܂l�:iC*���y�W�Qu�`�b	Zb��d�`��2�y�����dC<=@)c@�Ҽ�yRbĻ
xe1���u�oT��y��Ĉ9��[���vjH
"-Z��y�N7@��EjH�~J굑a%��y�(�/��(4E�8,M����ܵ�y"e�=X�d�U �u(�hE��yb$�X��p�m���Q����yRL� Ɯ��sLRu64���y�I^�ʑYc�G��Vh�v�ж�y�O �D`��+ަ7p�XR�����yRf֍8 �	r�L�~�ڨ�$�� �y�H6�,8��u�X�@����y 9�@���/k�v-:���y��,X�~�p%�_&a�t���y���%`���
�-A3R������y�c�<n��-Р胥\L�u2�o��yblɿgR��'�\Kb�����y"N�*X�fɋj.�E���@@B�I�,�-;qɒWJR��ҋS$h�B䉲l��Q0��}�00`cL3e	�B䉡i%�a1��W�<��@��l���lB䉖 #Pm���f���a���h2�B�	9R����C�4���!x�\B�9���1��F�p�@ eL$g:0B��7j��!p��~�*SE���^B�)� �8x�Η]���{&��$kvY��"O�)q��$�ژ@���12��h�"Or�2ĕ�d+�4�oCq����"O��u�:Q\�:AOO�v���"O�x37�μ|;�`�v�N(Yj����'�2�'8��'���'�'*��'�i�����,�� c4�R	�@�'���'*b�'���'���'J��'���vl=���
-j]���'���'��'@"�'���'��'����T'�j�\X�$��
?z��*0�'=b�'���'���'���'��'e�S��ՒfV�mB�;,�dI��'R�'�b�'�r�'��'
�'o�0����F�	�Q�Ć�,���'
R�'�R�'�2�'�'�b�'@��3�[;`ظ����j����'4��'���'���'���'�'RtAX犃y��R�K6��6�'�"�'��'��'L��'��'����3�F�;�`@�C �hQ�A�'��'�r�'���'pr�'xb�' �7K� �kV�}4Y��'���'���'���'r�'w�'�x)����$߸T�w!l1�L��?��?a���?����?I���?���?q�M�9� y�!ʓm@�����?����?���?���?Q���?����?�`,Pw��\2��I,n�x�kBK��?����?9��?���?���1����'�2E��f����N�oX���pf�9�F��?*O1��	��M�o�	J��UX��ԉ"-��M��)����'��6��O��O��O�7�M0LP��`�W	j	(-X�≐v�� o�џ��'!B���.��JBH��O�tS�K�#�h�)������E��y��'���n�O
:��A(J�Jh��� ��(��g�P���d�2��,�lzީs�ܹ��`���?} C��*�?q�4�y�W����x�֌�b����6�������`�b��{U�Ȼ7ƒ1I��ƨO�2�=�'�?ɵ�M-<R�:����a�@���m�<�+O��O��m�=�Tc�@��� P�z��uo 1I�Jm��	Jԟ&�4�-OB��vӢ�In}�AU�{��A�p�5~b��������M#������2�1��×j�+�>�䈌u������*�P����0l��ʓ���O?�	:*I��ի��R�{D��g�@�	��M+� ZK~��c�r�� �4����P&C�dA���&.����O0�$z����d�� �e�����HصS$��1҈Y�B_��9��H�-�D,���ZB�F{�Oa�b�S�O��в�KH5KF@�
W�4�g���(�+ޘ'�� ��G�9(Q$�R��	JhX�ɐmy��'�3Oh���	�O�d`�M�A�p�R&��Q�`��"��L�eS� �Ψ	��� �����x��-�򋔯r5(j�+T�	j����By"X��$�`bߴj����� �d}蘛�OLp(�͓K���4����O
6-�OV-���Z���[�k��c�%�eý5���u4O\M(0f_@W�=�Ջ������O�D��*y�	Qf�P+{2R�ȃMr6��2d`{���	Jy�[�"~��m���3�ሣt?��˰�K�y��b���զ�'�|�� F!~��h�Q�om��Pb���<�)O�7�Ҧ�	�=z�x�n��H��X�l�p��{�S1n
-=2���
}r��
A��'��i>Ֆ'sn��6X�@y�K��di*��O&�y��|"�kӢ(��$�������
��ϺW4j ���9��;��$�O�6b��&>��
:\�0��#ǐ�#J?������ BO&?���:����×in����߽z��y��F)l���ظ$8i�3��yt�1�EǍ��=��0d!8�F4�li�Ӯ!L�ɡ���E�40�{8b���9�BQf̑�\��E$�-��P����7{��Xr͛+<��R3�&=��3��T"�2i�*_;
O��r� N45������������,!e:��P�_��ɺ�,R!67X}�r&��Bw�P���`,z¦��([*(�5D���AG�)pb8)�$��n.X\�3"�[�`I�2��(D�d<��6��K��2Pf���qSN<���?�����O6��N1,����G��+#*T*�Q;Q�`p��*�O����OH���O����|�T�$l_�^cX��� /�zmFI���֡%�8��O��d�O
�Ŀ<i��?�$�	u���8On��r�g!H��4���)�M��?����?9�T?�� ����'r�2�¦"��J�����n�B4Iǹi���'�	��`�	F�b?�(0��,�f���0j�� j�g�B�d�O��O����`�o����B�daa1�K0�91�R*n�&!o�ly��'��`F$��"��i,1ȕM�&A�����c�#�Tqݴ�?��L���R�is\���)�A~"dôo���"��ɁP:�y(`AN>�M���?�UJ����4�x�����'�\�TG̋�6L!�Y*y���{�4P�0���io��'���OZO�W�S�Z���΀4"o�!baN�q�̜mZ R$��'rr�'/��y��'^P�#�H5c��&LP���uӄ��O����Y��&���� ��"U�Hق"����	h�(KP�M�O.�d�O�����$�O��d�O�l�댍h��E���%%G4|�2�	䦍�	�D=�ݨL<ͧ�?�����ČG�Ũ� %�!j'GC{k��m����0u+�I˟��	�l�'��a�ę�Y�ܭ;v�9	�qtH� Q��O|���OJ��<����?aB�  ����_�Q����E�{u�3g�Za̓�?A���?-OԵH�A�|� QǠ�( ۙ�\�p/JO}B�'���'P�I՟`�I�F^v�	12ٷ�3Dװ�����L����'U��'��]���T&,�ħA���5��"
��[v�Wߐ%��i�r�|�U�����8�S,��9��<sr�dbڌ�,6��O@�d�<	䄗2ȉO"���56)�!]�t�7�S���j���M�,O����O �i��S�?7-�'\�4�ɣG�0A(4�zu ��@��	ޟ�t��T�I���I�?m��uWO؄W#�Չĉ϶=V�P������O�ɑ��[=(q1O��l��1��6jȎe�Q�Z� ��8#�iI6�v�',��'b��O��i>��	�Yp6��$LD,�)��#�@��0�4$��uj�A�S�O 2�R,Px���B��Xov��Ɖ_�7-�OJ��O��k��<�'�?����~rc<Y��`a�_���Q=�(c�hkg����ħ�?I��~BI�',�XA���>_@b��@��M��R,R/O����O��D?�I�fUF����*ېК�፩D���P6^�!qk	c~��'��S���I�r���	�"Z,��̈́�Ek�b�E�Uyr�'���'G�O���!�,ႀ"ݴA*8ݱN�l��bD.͑w��	ן���\y��'��Р�П"���h刷��4H��ZR�ix��'��$�O��Sǉ�>w;��,H�a_�HÁ.?F���+-��d�O����<��(�R �-�z�$ʰab�!���ASqF��W�ǈt$�o��|�?y�no���fɀr≬u%��(&�E�EE���b�m��7-�O�˓�?i�K9���OP�$��j�32;(��U�їov�� 䃀n��?ɇ��o�]�<�O�h�aL�w�����=
M�A�O�����^a���O��d�O�	�<�;aǪ�ѳ.JJ�8D̛�a�5�'Pr␛E!���y����з���baJ��|�A�Ǖ�M�W.�?�?���?����/O���O���}yL���ɘ?&c$X��F�ݦ���M6H��b�"|r��|�!����>=���5%Y'S�d�2�iQ2W�H�6��Sy�O�2�'_���`cH�]�>(
5T�	�F���<ɷT19b�OR��'V�$_&fͪ rH>X��֣t�V�'�R<��V���I�l�I_�Ҷti�Ə'��mK��&l���L���H"��}~��'��V�x���N���C�drW���j̱Q��dy�'�"�'��O&�dS�0�T�CS�� M��pk����iq�ڇK��Iȟp�Iyr�'Z��ݟ֑2#�Vv�,H�lO�A.n���i���'�2�$�On[�C	
[�6Aʫ^\RU Ƭv�XQ'U���D�O�$�<q�� lB�(*����U�`�2��d�(\��耲c�0_�`mޟ��?���bC�u�T�q�	�`����RDT0�4X0��UQ�>7-�O�ʓ�?�v��3��	�<1��^C���A��T��p�u�����- @�D�O�I3���-�1O�)����0�g��}[6U�S$��0��mZFy�kڥ%*��'��'���S��]	�Ȣ���4{�����I���?�D�
�sy*��<�~"KE�}Zųc�Z
T@��yd�UҦEig�����I]yR�O��i>��	�"}�����_�F��<8aO�!�`��ٴjָ�%��e�S�O]�dӈtz�1+�>7V\�!Q��h�26��Ot�D�O�����<ͧ�?��~	��R���Z0�A�w�ld�u��Hn~c�����-�ħ�?Y���~"hN��xb��k4�4�%I���M��yj�L(O����O&�$"�	��N�f�¯zx\��Ǚ+��L���;p~�'��Z��	�+��k��D9��Պ�
�(�J2��zy��'8R�'��O���r�!x�C�.^q3�Y?1���(k�=h!�I�����Ry��'��<
�֟n�c ��8�Pd�T�B����%�i�'�r���O�	���H3$���D�f)�v�؅@k �Bd��*����Ov���<��ox!�(�D��S"����@-V�%-Ju*�lS�<�hnZퟄ�?��n����"FL�IX(�H�T�C��8�{t��9��7��ON��?1$������Od�D��p(�iE�J�Lh��'o֎h���u��?QD�1j���<�O�X��%6fh!��ā�M|��O��DMS >���Od�D�O�ɡ<��*ll+�R�hQ1
Q"� ]��A�'�R�ͣ$��y�y��䎉&�x���U��I�!��M�匬�?���?���,O��On�PЋ�-	i>0���D�Kє�0(�Φ�[&`�y b�"|������Rf�(M���c��((��8q�im2�'��#�" �i>��Iן���Ot��p�MJ��a;#�"�FQ���ԹQ\V�����O���$E 0�c��������÷�i@�lW:��I���	��=�`��|�μ���"ey|�'A�n}�ȅ�>���0�O����O�˓�?��O8ޖ�k�!vƸ�[��C�$�K(O��D�O��$#��ٟX+FK�KDC��_��XU;�E�X��K�+?����?�.OX�$[�[l\�S8V���]�e�́t��*qh6-�O��d�O�(��j��8Z�aj���0�9:hy��t�n�RQ�d����P�'b�6�����p��X!<BΘ��"= ������<�M#���'��O~�M<� �A��!��Y����	�4&o	p��ib�'g�	��L��ퟸ��ӟ ���fč��W=Tʬ��3I³6�Ly��}��'H�0ǡ�����iM�
.!� ��R{��g%����IğtX�	ǟ\�I�?���uG�[���6\:�z�F[
����O�(�	�I%1O��~=;�ڼ|��ՄP��a��i�L����'���'���O?�i>��	*p�ઃ��!�B�P��Q�^�Hߴ0 ���s.�W�S�O���>�ҰÏ�3� (@�A
 0��7m�Od��O�Pj㦲<�'�?����~/�5��3B�YbT�	�D.Ɓ�c���3&>�ħ�?I��~��^V��u%AP��\zr	F��M��&�t�+O�$�OZ�,�I�!/ܪf��!a����D�ƯRv�). !�A�AZ~"�'2W�p��E`|��3HI�>��B#j< ���Z�VHy��'���'1�O����?+'�-R7�l�؅q!(�"
��e�7��
�Iɟ,��Vy��'���۵ߟ )��FT�Jø��ND�Bz h�p�i�'�R�D�O�e����7���`�}�
	a�hN�\���ã�6����O����<��d��a(����>^t��@�,۞T*��׀0��n��$�?	��p�l%PÄ�G��Id��!ݔ~(	A�ԗI*<7��O��į<�b�P��O9"�OYdɃd�Wf�V���5�s�\]��'�B�'�$���'�b�'a��O�~	3�d��nz��gk�V�X��n�t�d�O�p!$C�M�������?IY�O�=PWCK�HRH{ �aŸ<�&�i��'J��'���'��p���&��"�/s
J��j @��#��{�B6��O��$�O(�I�H}T����)#�AsǪ���&�rԨ�)�M�U��i~[�����~"����@�Y�s7��lةr��զe�����J�r��4�?i���?���?��=G����,��W� ����8t��<mZџ��'� ���)�Oj���O��S"+�C� P����p���AO̦��I�u�J0	ٴ�?a��?��.!��\?�d�	� �	#�_��1P-�G}2j��yr�'Xr�'�r�'�哴c�!	�#G�-2rl� %^j*U�À,�M����?I��?%T?I�'�r�J�>��5�楖�dvV���e��1?���'X�Iٟ��I�d��ݟ,Ї�͵�M3$�	��<@����',��c6-
s���'u��'���'3�	Ο4##c>��t��8��B��V ���Դ�M��?Q��?�vV?�[�l���MK��?Y���,[�*���,�@T:c��_�v�'���'�����Cǉ`>m�IE?	A˟���h�Amī0Cvl�įզ-�	ן���Ο,��L���MC���?����r����h�:�J�'/�V�C�G=�f�'���X�6�q>�&��s��X
\�%:v𩠨
'Be�вij��'`��3��d�T�D�O����`�i�O(�:���AT�Q5l�-\~M�cI�Q}��'p0UH��'��U��o�I;_��ܢ��Č:V�1&@�+X��¡\�z6m�O���O��)Ꞔ��OR���<)a��" +�]�t���X=x�Am��J��A�'��i>��|��*��ect��5�D�!%O�)�u���i���'�����	ȐOJ�D�O��ɮI���!c.;��)��!T��`61�$l�?A�Iџ ��"~.��(ɖ>�����$Kd��,ٴ�?���݉'0b�'ɧ5��&r��4z1NN%Q�I���ţ����^�Ĳ<���?1������r����D��D"x Ekĭ#���H��@K�	ɟ���E�Iɟ��	/�1+��?adDK�AW4(�����y�_�P��͟x�	yҍ@F���S��0)�.�m�p0	PKK����?������?��!��I�G��3�αn�~�i�gE:>�x
u^�`�	��	hy�ߔ6����0�W�*X�؁(�+��$0�]�b�B����I�Iş��ɇ����	|�$��'��d�qa6m"��M�^����'�V�Њ׋����'�?���/�N�ҢNս.'�1��V�Z&�x�'*bHQ�J[��|��h��.Y�x���̖I���$�i剎
���شF"���X�����$).�ȵ��qZP[��1,�6��O��D-r��%��ɔou|%��-^(4�	� ��9�v-��#�\6��O���Ov�	JK�ܟh����
����C.�4�BЅS&�M+�h��<�M>E���'.�j��a��#��Vd�\�5��6���Ot�A�]���'���Iڟ���'��cI�(Dw,��V�kzDo�`��y���)����?Y��CkDmi���q��P����o5N��v�i�� MF~OX���O��Ok�E�&S����$߹M45������%@De��_y��'���'�I�,@KbFTv��+��̀�
�ē�?	����?���M0F�!�ѫG�FJ�hA��Oy��?a��?�)O�aD��|�N�'���sb؄`(Ł�m}��'��|��'��ĕ+�y�7���J%��j[�5�u��ySJ��?Y��?�*O��A�m�z��!;��0�׉_����"(~��$�4�?�I>A���?���[�?1M���	� g�R���3`�����z��$�O|�Vp�A�3��4�'��\cȶ��sŞ'ՠ�A�똠2�P3�}2�'.�`��'�Q>�9p��i����5���o��D�f��>!�f^�D����?a���?�����^�z���qo��	� L%F�a��i"�'~��Q+׆Ә��π 4(ċ4h:���`�y\:yr�i4��V!gӒ�d�O������$���I6 K������ ���m�
a�q�4r��Ex��)�O<a[v�ߋ� �f	�u~Hi�֎�������4�	 @2Ʊ!H<Q���?��'�%���l�����V�4�%@�}R푮˘'�2�'M�l��w��Z��Ɣjf�Iel����7��O�I�@L쓡?�������R�g�+ys����_��&S��);�	ݟD�����'��H�WE�cޔq��,��J0�¯|��O�d�Oz�D�<),O҉�0���ƒ�3�K�3p~ē`�['.91OB�D�O���<�w�����:�0B�d���0��0g��'�b�'��Ibyb	Ť��)U3RlX�W�Z3��0(mN!b�I����Iɟ�'����5�$LA3��>&U*�"��ְc��m�����	Ey�'�r%���O}����B3���4J;X/4;�4�?����7HSD%>��	�?��>Upmx�o�4d�M�j��ĜO˓p��PD�tܟ)'f㎼��[2`�\�ɵ�i#�ɘ5��ܴy����������DV��C���t��8��� 3����'��ΐ��)Z�g�	�l������Y�$sG76t�6�b�����O��$�O��ɾ<ͧ�?���];<��`GQ=.��(Bn�]��߬`<�Q�y���OR���I�������Y���!f���y���� �Ɍgi������'R"�O�	/��T+X<�`
�f.��G�e̓a�`�S����'���O`U��^.?Bah۟<���K�i�"a3d3�	П���ܟ��=1RK	�>,��Y"I`zD��b�`}2o:l7���O��D�O��?�Aj��v�Ep�o�9 ��-I5m���/O��$�O��=��sA�L#A��][�!(²����[J��c !?Y��?Q*O�$ɟh��S,��z5#Ƭk(P��W�@	T�
7m�Ov�$�O*� ��2OBI��d|Ӏi��"&d�<�N��BHG�Mj��؟���fy��'��
$^>I�	�|����)i0����	�m~�c�4�?��r�'�|yxA	ę�ēss��FV&-��3�(49"hѤ�P�RL��c��$���$�g?A�BWA��̡��G�2sb`��In�<�/N.Z�zP$�:}��h��fX'J��l�b�D,I(��G��Q	�%�͑#`��PG�l���Tc]-^ݸ���-�$�e��͛��J���i>H�
���,^�6�T�J�)Y�)�.�#t+�����#Ȑ�2���8ck4\�Za�ARl�%{aD�&{�8��u'��(� L��A�/7<����)�>Z^T���?9���?i�*�K�+p��+^��(1���;s�ll�%Y�>H1�[T�B�,+�3��V�"���c��y���8���x���+�O�f��GN�}(�@X�/:��DM����8��`�f;��d/-=.��&�O��]Yz��i>UG{"2�x�����6 ��� ���y"�I.zVRyc�;���׫C�y�'��"=�'�?!-O�x��d 0P�D"`���l�k@�]�;Xz�H�O��D�O��� к��?јO�0�pB�Y(d.8��G�0�R�;���+B:��G;.��'{�իR���D�F��oS0?���@/L�)�i3�i�0`�*���i ���L�6s��wI_0���Y:m�T �2�x��F����B�'7���g����%�0�۩3ϴ���? ��!�ȓE�����oZ�o��-���P1�t�<[�H�'��!w�>y��R�8���N�-��\9�l��,�0�����?��D��?I����ԫ&���j�9����)��J��î/��� &�[�uPY�㉾8�l ��a1��If�Ҩ���4�F�`�<�3��o�mH���e ҟ(�	qyRE�3F(�52C̊XI(p�����'O�{BbQ���}#E�]"��E�V��x��nӪu������I
����i���Ѱ2O��ChL��i���'��cW^`�	8*t|p� ��=xzՉ�ώ4���	ߟ��U���(�.tA���q鰇}���K�DJQB�����\-I!&�2����I*m��̈�#�m��7͜��$�J�m�>�|�[UD���ÌV��ӀL��s���OV�K��'7@7�Ԧ���h���^9�,މj�m���O̜��<�����<�U��\TY����&�t�Z��(�hO��z�'a�������%����S���A|:]�$L�"�'rB� pJ��@�'R�'��l���G)�m�L$ʲ!Ύ(
�Y�òM��8ٕ��9*��r$�u����|&�x	��Ԥ{�r聄��.�@��@�
7��M��
�{8f��P���O,b�>�O6Ӱ-H�}	�#t*^d6��"�.�f6���|�G�;�n�����d5��͏�yF����p�țAN�]��E�yB�'Hp#=ͧ��y6=R!��Y�D㭔<c@0Xj���:��a����?����?1��b��O<�=�6=���t�`�җ*V�6��Eu�ߛ�@��d�t��`{���Q[�{�k۝)�t��um�&pKa~d8�����R����C���)Rl����?����?�*O:��/��>���/@< �@ZV%ǎ\BC�)� �P`E�/ܐ!�Q�%��t�D���~b^�Ī�О�u�'HR��
�Q��<Ϩ�C�Ȅ�2�'�jY�3�'�"7���27�V ���:T_�t����Mi ���2�bX�G�'O�!8w S>���^����\5+��Pf��0]` �B�#O^�`��'��T���5��8����JK�P��Íb�\�	ϟ��?E����r�`�b�Q�!�6E��&ƞ�xbHx�~X���>SP�CO#x�<��<O�˓#��T�X����l����-e2B�1�\HFȄ2b���r�τaY�'��"�@�?�2�Pt#��f����;~=�a\> p�Z{0�� ����k�j2}2D�"4\4�Ѵ�4f
�:�i��J~d��%SK��
�U(��n�&눑"Aޏ��	�;M��$	���ӏ�I��4�(���=<(  �����>�QTg"4���J]98{(83B�R�A���N*O4<Fz�kM����a��A;Mp�`�L���6��O,���O�)�dķc^�d�OZ���O~�;e
dx�����G�6� �c��SqHDY��nʛ��_�$�<xoM�c>��6eZ� #�D�7mvzi����6�L4;r��o�yB�A���ߑv"����\ܧ@"�����c���ԧ��!�`�B�-íR�0�! �M�!T������Oq�R�'��٧Mz�����?��QBV( á�����Z"MB�A��u��(l��I;�HO��By��-T��c#����}�C��&]�T��S�O�4���'R�'Y��]�@���|2���%#i�"�ږRl�ʑN�\���s� ���tѸ�1i�-��C�%�O��4HI���/l^�ܚ�fP*��=�����r�p�"BB�q�bL�����	��M3U�x�'R��G�"H�qh�m����A���j!�D�3]��e��M.X��e`֢ C1O|��'�剈Y���8ߴ�?i��]������a�
������=ܺ����?�"h��?����ĮG?��t���	�f��Q<��,0�`Ք v�QM\�#���Ie!B�h��-HM�DAc �4cJ�Ƥ4ds���.��9A	P)�F{"*��?�T�i�6��O�,�LU�m8��)�
�	�bM�u��<�������v9K�Lߋ���H%��m�e���	p���D$fӆ���bI�d}Np	��ه}O -nK�O��OP��3?�7�Χ7r0j��
�|��D\o�<A�d%��=�c�k��8Q�`�<��Z�TXu��j@�|`�NY�<�B
@�����^)<��gHa�<a4��r�8źuKkm��a�c�<��%D+B��b!��jk��gW�<�rȟ�,�R���$ ����g��T�<QK��
�t8D`���0��S�<���@�<p3D`��&��-2@XN�<i!�ŷd��� �6ڝ��&N�<IuN'`�%�tC��]*y�G��<���� �pm���ތ�Ԙ�wG�R�<���j�Q1+ʡ*#*�iD�?9!�Ċ	*0	s�[�_P���d���!�V�dT�m"�,Q�8^����[<?�!��� ���B�IR-z���1E!�D�Z!�r�S��A����(l,!��=s"�97����-Sj35�!����4Ь�	pa��>M��B�OB� �!� ��#&��
i�8ؒt:�PyK�P��uxFL��aXMbfT(�y�)��D�  ���ȭ/u, j�'�y�+A�e��t(�#�u ��E�<�yRN�2z�P�Pl�9�"��$�y�+��j�ڐ3pk��q2�"�;�yr�Y�v�@�o�e��+�/��y�h(@��o�h���F삸�y�$�'�l *��2`���B�yR ɦr���
'C� �*���&�.�y����|̐%�%m��z�)�P�y��]<JHxZ�J��§����y�J�#��$�#DFh�l֏�!G$C�	%4x��όW�tQ	��ƅa�B�I�|��|�QE�-(��$aP�����S�? 
�Xw ?N
��p�v�[w�'��C�fͱ��so5e~��dO>|>d����/pwvQQ��(�����K��8�����}kz!�E�.
����B�V"<R��*Yz��F ����;Ã�g~�όW�Xea �5%�f��AgW���z��'��Q �Ɂ.�IY�b��h1��5@�����UϨ�"b�6����9�Y�'Fċu�p���A�==�@�`"O1���Y &ܐ�f�sl� ���x�qOf�O�� 4閤t���a�X�T���F�>z~�]�od��r�-�OB}!g����*E�`����c�^�_��� G�̠뮹؆�a���I���_lX��h���O�0��L�H)T|��M�*Gܲ����I3�>c���_R��VO���6��g��Q!�Qgx՘�/��L)�%W(U��3�A6�#� �?��%Z.,:R4�`�O2�P�A�AM�ua���'MS˦�I�&(�~*��n	,��,Ȇ��!qU�]X	�!�6���S�ΥU���U�~�?c�"2�� ��L�0���p����qv�( 3�  )Ŕ9�΃Ox��'rs!��D�1pk<��O�$���O�*u0<$XMF�{�v,�qE�*y�P�Sb�'�u��e�2_פ���bȐ��2#�M��^qsM�2Ml����s��U��3sWt,���~� �	'f�����v���,�T�Hl��dȋ*ݚ�B�I�B�����I�Oh��"�ٰWպ4+ƍ�u��� ��;n@���mKf	c���/N�ظ��O Z�q�@i�F�<���[�OI\AI�ƭ�`ȑDôdG�1Z���$�l�(5�|��MIr�5�\`��׏V��aʕ\>�Qu��@�!/�J��I����Q���I��`��;��8Fx2�Z�T����HPn�,ؐ�AK ���I�/����e�Ȋ9]4��Oz2�˅DI4
�ٓ�E�~�/��>*��0/H#�~�yl:ғFB?U������?�2��A��]�����ʩN�@����%�So��zL����D�m��aY�NuqD���Pݺ���%A�"�ji�9)�(Ag��\�'h,ё��ȑ/JD1��O�)Cc���q\����2(����`�<�Ɯ��I�.H(�-�I�?�6!ɷg�	����hQҢ|����m��tK'��7RW��h�,9����V�B�x �'cd��ËĖ9���P��k��9�&$�1�2^���y����w���kR2^� �K�G,�xu�+Q>�3��<�"�!S�.��R�� OՖpn�'��`f�5T
x����� )�������B���cs��T�t��
�AD#04�qRfb�#+�N�I��P�D5 ����8�D�\�T��	�Ƣ�D����F��O��4Z�/��?Ip��/+hL��B\�e{r6�U'��d��	�����9"�	��+��pb�D�T6�DC�k(��rB�'�� �'��EA5c�F@��B�b��a�'�,,v�\X$/�1�4�I0����fo�ey���O�Ob bc&�8{!�bC�A(V�$jV�R���XVt�$� q� �sF��P�B���(�?��m�8��͈�a��-yƁ���Q�'��ٲ�8G�^��˟���`�=#����\;F�(gq��cͤE�@�j�̋E`,�����a�'Z0��'FA�;s�!��L��H�0Ax`F��uό��5�	2�0=1'�֊F�șYc�$�)�IN�{�(� H�cX�(�G����ӆѡ����'E4��~λ`Ԧ�h�H�5+ l���耎+����!]�;�ʴ]\��Z�K9I�x��&L�`[�dx/O$��jN�py�l{.O��%?ez�mȌ�d�3L��2w�ώLɴ8���ĉ=2
��,f�n�9�o7�4��K�Lmb���)��1�gfE�k�������¨��U5���5-Ll`���YD��n�5v���N��71`%+Õ:G;~��T�*���ɘ'��n��}N�$��c��/f}�D�����lX�8���Fi&|OTHY��%�#�Ȟ,8F4!�F��uBPR����VeDi'�W�$cQɜ(0V���v��ai�m��H0*F��H�p�'���B��¬(���h��W�J轰�ő2o2@7�2e�ܪ�H�S��bE�]Y���ۏ���,3�� "I��A�L���ɴ X� 9��S4��O��
&n��<Ϧ�F����ú^*Ia����`B>'�,��%"��P��YX�#y�6�1��z�
d,���'���Pp���Y��ܘԦZ�GӚ%��Ot��"�քvUj<��$���s�$[��C�+Ay(xxq��F8� ��aP�p�>�A���S��) �2o��H�˧{h�p�p�ڋy/����g޹gN�K���ce��~s��gm���wɨ���9b$߲`��m�ӫ9�jx�'��Su���vf^6D)�I�V�	S��(��_'��;g�ܜ,��O`l�vG]�}*ũ���n>�;�i����6O�<��Q3@�Fzo����*{T!�W�G\|�s��-P�����x�l��%[�iDvy[u�J�lm ͈3eжٲ$�Bl��G��=����'
8Y��낔D�t��	�P!����>i��HQ��.���U�8x�����(j����O8 �v�M+]8��+�¦�pv	b�	�|�'�^�)%� f�h�s	��E'<���B����[0�K3��ʒ2:o(uG{ҥыt���\&|��͓�@�,����-l괈/O$��OJ�c�	*i�$$��΂LL!��Oވ��go�Q�Q{A�eP�};PcD[�'�j�j���$U��a��
�hK�q�s����$��~�����U%Vμ%�Hw�W�^�=TNu"e�Z�:)�����?����EN�$�
-����(K�q[�`IU� )X��I�-L�����M!c��Ջ�������[�"���'h�i��X��ͪW#�%�ݢgO��>�9�E�߮~=BhC�J�>~�8��f��l����+4�	$n������5	� ��-�-ΚA���
�M�A@�����'�%��X1T|�ȑ�F6�=��%	�ʶI�Uś�UH+�+Α}Ԓ�+�����-�dT�"k!CR� ֵC�1z �ݟN�>p2�Z� r�[�ppqj\9 �0=�Ȑ���ݩ���?�A�	�=����ˎ� �q���������3D�֤�1��=a�@������$�-��P��R�N��8 ���oY"���8ժ$	��� �%��?Q��B��9"���/�"�R����?DZDˆ%��f���z�	E�R����G�U�,�r�h��όP�+���h��e>��u���DȈ���/43`C�A�X
��pN��p�� ��@����q��OgT��?��+Ƹ:�~d�q	Ӎ�A@v �:;b���W�d�O��)����4��$�kM3g�X�`d�׍7`�r�L*P�1⃄-�h��ua�'�]#��.Ō�"Ub�6s�hl ��/h������G���D>�D���^͊��&��<Pd[�)|���U��h1��$r*n�� k��"��Q����O2�@��	dTݠ�	� �r`��g}b�X� � x��B�q�Ta�![F��K� ��5�>tȐ�^7R��0��I�@ x��R�H����㿣�܋	��4�� #�`�u�j`̼��b\�_ 1 �?��`��O�Y����=�|��@�l�Z�R�R`������8$8Ċ"�T�k]<�C������.��'��x(R.Q�'p�"�f*(��� ��be�xf	נm"��c���<��TACL'Ux��Ԍ�*�l����,7< (�⊼�XP�n����v�3\O��
7$��-C�����I��r��0���I�g�NMp�8���[�NŔ%���;���&C�\��c	K��uN�;��f`M#q���5
Y#�<���к��53�c�X��3d�*F���Wd�|�Fy��kį8<X� @'^�~M���e�5�V��C�|��Sl���)/ֿ����="���SaZ.'@�a�Q�a�ɔ΀Ɂ��A��]�C�F�5��IY��S�K�(M�"ƒ�w}�E�PD�(!�,�����&)j<;SOH�M�ĬP��c�Q�0A�:F�O��	��\�8/X�@�R�r+�}� ���d�����.$J (������.�R�݈z��S�Z�ص�եکa�j��C)d�8���L�պ�X��O���#7�D*z>������ر/�` I5�T(~.̂���?q�6M,`!v��O�.0���92p!K1�T>��W��8�ؐ���H0h��L��(4,O��#ecR�$X��mA��?i��r?@Q�G�K�^n���QOpks}��$�aN��^}>h(q�2?@P�C»|�$9�V]S�GX �c�đ�U��-���x�J�'#~���Ċ�q��V�`�L�?e��ၵ*R(��4L�RD�fNY�;x� T�FS�a����uq#��6=�RmQ���'$��U7];6Bf�M�mB6��>8>�a�c����.�%���O��jW'E���)Ϳg��T[1	ٛ\5�0��ʞ_���9R&_�Q���Q�8\O��[�GG�q6Tt�W�]�+��i`�ڷ�duY�CT�8���1O�\uW?��d.�I�$Ae���놎Ϸ\�����ő8��tKƍ��<��M�g�`�Cᆬ[�����㇂L�H"�C�b&�a���+��i�<lb	����p$ \:Ab��6��}b�◢@�dkg��B%=@(���S'��:��Q�⒅
|A�`c��J֨���4�O�zt��8A�ݚC���2k���W@V"D5�iLΏ}��Hi_w=�4ґ Am�b���T]�(2��Q��1Zh����
5�T�&�߯PU(��.z�s�px��~�7�>(ٚx�¬{����ٞ=K������o4(��דo�4���a������Rr��Fӡ��`��.
�*�!���u7+M;,3Ғ���',�lY�͑P�F���l��"h&���I�c!�� �e�$��M,_l{1�AXmT� �HݮZ�����dԟt��NU+b��Q�_���)��6h��8��ċ�%Z@x�� I9T�t���c�'�ē2(J�p�#��y��L(%+��dd�8{�"=ZwmϳQ����-�ʓ}OEG�t78��;"<Xs�D�*;
�YaC T,$�\鱦�\��'ȋ5v�B�@���>k��$�������A�
{��YsBJ_<������3�x\�ˊg$��× �9m~z���Ǝx��+��;�0c`F�^�$pp��79"ٻW�p�f%�'}�>��'@������>�a!2';Cl܇��'P���Fl^*B��ٺ������8���KD��!A�xF���w��c�Y�`iQ����O?�`ᅑ%��p��&?&���p9��ʹ�L%Ç��]�"�2�T5<���>%rAIֹH�ޜV���6(A&D<?9!�t��lR�D8O`�äm�znTX�5m
3(��@�Z6���N�S�1����(dѱ��a�Og x�bN��`��\��PT�0%�u�g��x�Ɖ�n��l:&-�9%�4S�O�P���Rކ#R��QVFCEy��n:�<��9c�H$Ar�Y�zF�qf��8v!j����8u�� Đ1lB�:c�)k��`�Ó�;)��2r
X�~urx��ᡟ�K�l��@�����>E�4& �.^H�#d�2_����o��ē%>�8Y7$Ϩcp��V��+i�[����P1$�K�i�%_�����7��O`X��	T�1�1O=�dL��=Ғ�!��c�v)W��3Fd8�'%I:"9@�;f`װ2ձ���i>�2`lٳW5I�2���<}@�n�	CF�<yQާ56�.�.$i��j,m�B��S@��&�R�FQ �ۥ�y����S�3}����&�*���Z�*d�� �*��<YQ�	 5�Tʶ������iH	V}�p��s��b�b�(���b�'פ�Q���T�E�O>QK��
�>�1���Ua^T��0����^U�� ��L�rE�;��OUB)ђ��_ �GD3J<XQ-$�DTC�<Y��L>A��Mv��A������!E�YN�<����+����T�ȑ�lP��VG�<���ޡG���r4�ۢ|Z� ׁz�<� Dɲ�ɖ�hlD-�aJ�&!.Nݛ "O�ɡ�ʟ�t�����'�Z�"Of9�F�4WJ&Ti!	��""O�$Q���o�4kv'��^�hA�"On��t�åvΖ� �%�'Xڢ�r"O�<��^!9��� �B��3��Uq�"O���Р��
"�L	�,��u�a"Or�+���*	�-� ��4O���2�"O�8&�-���Chն;��#r"OMie-�3x<� �� B��Ҥ"O�l!U�S)e.����W��4Ra"OŻr�H�2�`���j����"O�ܙ3e�-Mn�<c�ȈĶ5Y"O���ĉe�j����H�3�1�"O�԰����� ��A;M�>��"O�D����}�LωN�|�6"O %CEh

L�xq ��<:�tmآ"O��sS�,r��hfK�!(��R"OJ��@
�n?�� �ɗ;r��J�"O�J�- &Ȥ3g\�j���"O��s�/%L�D)	ΩG[��B�"O(�b����I(H�Ԩ�fN �"O��r�K�S�~ �1�%S�ݺ"O6\�#O�,�R��pES��C�"O\��6��8x���񕄌�%"�1[f"ON��b�?!F����_\��w"Op(�"��~���K����=�t�@"OHD�Aj-	��)g��2�8� �"OD��qd��j�L�y���[�"O���#Ȧ�Dt�0�Q
#2qsW"O4P#P&L6`�����T-t��"OJ�[�A`H;ʅ9M���$"Ol���E.nhQ�K�٤A��"On�q�ק"��� fH�^�DH��"O��*Ů}K�5���q��-�$"O�cJڮ](��W��%s�&``"OJ���. y�8�C�e�Mx�"OJ��*̌e���cb�
-ܠŪ�"O�� �e�%9hjH��֢�JlÂ"O\UpJU3?�z�ҥ�J�O�(ۅ"O6���̝8m����U�_ JY"O�!��M�I��i�ݥF߆v^@���j8�qJ�Œ�JX�K^�P�D��ȓ���+	� �lT��	�@��T��]��`�F��<h0����*ʎX��r����4Ć
<�!��9/c^@��D	�=�Uđ�l�Ј4�K8o��U�ȓ\/������j-�"�3iFq��bz�&�O�KoJ}��h�0p)h1��m�ri�B��
뾕�F_�Y^U��u��\��^��Q�&B>k����`�΁�4�P%O�t�"h�<𐥄�$/\1�Æ1fghJwE� (Xޥ�ȓ$��"◸��d���R�4P�ȓJ�bA;�@�mxvX�bk�	p��� 7.��s�O�9d�{�ܑAд���
P�Y��	��%d\n�x�ؓ�;D���@(�3T0��kY""�qC�8D�ТŤ��:����/�p\ *$l5D�d9�F10v��%�C�@��EhĂ0D��"`%:��rէ�'��� l.D�t��d
;�:`��,q\~�1&.D���/Q9"����ӣ��"��X�e�+D������gV���N/~����(D�� �I0u���@�QI�g^�3�D�z"O �K��q�n�٣k�/ռ6�<D�
�E
!�2���� �v��u�:D����J�2LP@� �#���#�9D���$�U�"�<�8`��)ҲY8�*O:�Rҁ� :o�,�Ӣ��l����"O���LR"G���tA�u$X"O8���϶�D1�`K�k��b"OΝ�el�%}g����4c3�T	�"O�y�D��9j��;�GQ�$\L@P"O�B�傿=~e�&��:�B�"Oh���(+O�.�k��=�g"Od���-M0-{�*��B�X�;�"O�{��ީ
�2�V�T�1��8��"O�P8�̩F@(��r�մ�����"O�@
;38�D�I�򘨧�'Q����A�{����f'A�	��5�4D�ĩ�fֈ�4�X�������L D��sp%�2,t��CND3A�N0�i<D���;5\`�Ҁ�.8���`'%D��"�ˀ#W4��D�>�%��!D�Sm�� i�($��-C�4��=D�yÄ�u 1�чƱbg���Ԫ?D���u��#�D9ۦ+D74�"���"D��24�.,} 9ڕ+�5H�@��� D�x� �W<� �S���9WI>�cG>D�����Q�f��[�a^0=o
8�0�;D�h���E�5�L����?�M��:D���7J��rG��ȁ��5Dyܡb�J7D�4�w'�*K�M#�����K4D��Y�$�_/<\ѷ��bA�0��0D�,d�#f�49[�I� ��Xv�(D�43Tᒣ5��%`G�ͥ�p�sTc(D�`��@�#&���>�%&P,s(!�$�Y�ʼ��+�&P�t㓫	6�!�䛯0�u��ǒ�I)�tۗI7!�!�d֙������<i�&��P�!���,Px�pyU���:�6l
�e	��'E�$�B��_��	���W\6C�'��!�hʋ\*�DQ�|5�'w�#ä�o���+�ϕ,L���'�j���U�`q�B��0���'64m:��T�S%�;{6Nţ�'�\�R�k�%S�&�pg"��Cx&���'���4*Ӏ�����/�*S0��'���hs*Äj}>y%OX! RE�'�� p&�Q�]����?~Q��'@����.��Cf��Vh�����y"M�J���N�\E�|+��z�<v�NUN�!u+�%~Gh�ғ��^�<I��!C}\ ���(/�BU���Z�<��IŅ.�Hi��O��L���"��T�<�p���U�ŹR�z�0,����R�<��F�p�,M�wnX�AL+�Q�<)����3�`|���ٗ����#�	q�<y�A�s� �ʧ��<w�)�O@k�<�u�?b�.`3q�7���!,j�<1��C�0��q2B˯/4쳄�Vp�<���ʓ1���8�F�I�&�SA�D�<	@�Z,�zɑ��R�.�3҆�<���V�KH���P�K7n�b�<���V��9����� dC$��^�<�T�.�z}�P�����B��X�<Y�Ș�/�4�*�M�v���E.�z�<� b�	Ξ�g6��a`���:��	��"O4� 5���R�8UcG�eG��t"O>}�`��,�l#�l�
�)�O���e�ǏL.�U�Zi��[���U�$,�O(
�bR�4E$�R�W�z	��"O� ��J�J�D��&Ü�,�-:P"OXu8c'D9~��+����h�]:��}x�T�㪖�so�qU �; N��׍;D���V��I�x|�W�ݛl�{��8D�`���h?�1�,�|v�`9�:꓎ȟ6@��U8v6��@��l]��R5"O��)��:����n_<}2t8`"O�m�����]]ȁb�N�3d�|Ȣ"O6��+�%1j�J Ӱ ��Ұ"OTL��CÏmp��j�
:��h���|����Ѿbx����K�UĤ�+�#�!�$d��� A�<(Q��T�*��U"O �+�l��eg�m�s�����b"Ohe��ϟɴ��_�OU�i(5�>�	�y���2ǊM�����Ɇ���,�ȓ{�f��5��g���K�GR�nj�m��E
v�0��T,5���#'cÜr%nЇ�7)��������4�L<:pB䉔sW���d��-?�P��*�M#dB��;6h�Ӳ�41��rS���!�<B�4N�,t�eDӇ
��)Sl��C�I�'E�(�s�	[��0�ϻ7��C�IC �|1�l���$-���� ;�d+�Sܧ YּA#��`����ѥx~��ȓ%J���	�.�	'�D�j�X\�ȓw�Ĵ
�掕>�$"�T ?���ȓ��\`�B:jbn����<, �H��x�ܼ����W��-	��^7l%ܹ��-îx�g�%j���䉉wĄ�ȓ;�yh�@ʃL� ��� ��хȓQk������?J�r�`^,4����(��u���zԑ���&��Ʉȓ7����4� �`Z��q A08v
�ȓ,�!�JY2m`�t����mN���KÅ�BLae�͛a}
#G1D��&��#9��q��qx�m�Pg4D����((_��0GO	�p-�c0D���bC�IRH�r��NF�@�1D� 1Q,�kΎu��Q!m��͉`'1D����e�]����̄���5��0D�pPc�~E�`%EA8=��҂�/D���D������C�T��1�i3D��e��3v�~,b�`��� ЀT
3D��J3JJ&㚘*�C��r_�4��1D�D�3�A0eP�Vǚ�)������/D�h*���$%x��!bG�)'�e�e -D��膤_�ga�a�˽f�W�*D��S#��#��Hq֭�(VX�S�&D�P�O��g������zjF� r(D�H�蘜K�ZԨg@�O�N�sh$D��ZW@��5�0L��q2]8�#(D�`8�f�06 �[�C(h��+D�̲�	ɑg�����3��|��k+D��9u\5&�0hW_Cd�`R��$��p<Q��,A���p�N"zSxlY!�@A�<a��ڃa�r����6�ܐ�o������Vi`\��_!](��R�@�Tjهȓ<��g��y�c�6��=D����M�9��x�5��;.��bg�;D�� �y�6²k[<U��S�\����4"O��3*	�	#¹g�ɧau���R"O��b��G����[ *ent�4"O>��o�/y����oԨ.=����"O��"ch)bco�o�l��I]��y�gS�E1 `ʷ�A4�L�ړf��y�Q+��b0_4��0��@�y�bR9Il�Q��
��Vb��S���y��ڃ9�n ��Q�8��Uk��y��Ԙ>�̩�����:�ݑ��M-�y�j�lb��{eF��H�t������y2��5��m�g�ۋW�p���Ȕ�yR�8m?.!
AP!nX�S��y�M�1P5>���T�r�`�FZ��y�nZY��z#�R*e2���y��N�m�
HQFQ99^��tG���y��;�p�h"�i�&�� I��y�Ȃ�t�1��<]4��C�"F2�y��ױ*gF����U�
����J��yB/  J~�9������
��yR*��tV���@2w�P��Ƶ�y"n�2d�|���:e@ʥ�!e��y��["I`��b��Q�܌Yth��yb�Q1���)VJ	F��Pb���y�ɘ+P;��U�;:F��p��y����Qf�L����5���{DO��y2+�C�vݡ�ə0[fy j�9�y�
4u��|Ц)	"%�ȍ�����y��W�;%&Ź����\�'���y�UrڼU����:"wf��e���y���\9ޝ�&�Һ-�:�@�g���y�$Q=�2��eɑ�}|^�ią��y2�J`\a��ֱv<X�y3Ĉ'�y�hM�&�@��A�x�TJ�H;�y@C��VE�4�~������y�f-u�r!�K�ue���sÃ��y�N�wT�Z�IXm�d��@��yr�I:t�tC�#�(V��谢�X��yr�G�O�@:�hZ�M�\I�O��y���;#�^$`�MJ���0��X��y�/@'gf� UiS�;��� �.V�y��
4D�! �9,�b\�t�·�y2lڞ@m҈�F�9&�Ҙc�i��y�DߗWݾ���Ǚ�&��zѤ�yrl��Sa���w�&�0��bN-�y�ܳ=H$��"�	5�Yg$Q��y���8*ر'-�.x�������ybDO �U
*K�s�!x	]��y���7'b����#nҮE�����y�/$s�� ��	`޸<�q�ׂ�y�@�m��m��'�9lb2!B����y�S�mp,1)�Hc��%�F
�y�D;I�:�;@��1e]� .�;�y�A C��h9�b�`h�i�Vc��y"�E�V�(���;bt�3Ƥ՚�y���e�����"�,AQ6<�y^=p�V�1�ɞ�!P.Y�RM�	�yI��s�n�"�Oȶ)i4<��`�=�y��?~pX�7m�����E<�y�T�A�1账��}�L�!�ه�y2��7!X ��t�@u��g�y����Y�WB��!�����V7�y�G2^�]�u鏄H%ʈ��&<�y"M^�0�A����o������(�y
� L�����$eÄ�v+�P�d"O��Æ�f���ʖ�� "
(Q�"O��2�0'VкAF.B�(���"O��;�A�d�L���A兀0p"Ov8���le�t�@c�{�Ȥ�"O�-���w|�c����J183"OHb� �1tN
�[��\����"O����ʓV��u���"01�9Xr"O�0B$�+����cL�3����"O�pF@�R� �sYY�p���U�<9���*�`%�s���Jk�'�R�<�W
Fx�$)�$mՖy
(�jv�i�<�6G]��Z,(%�
�cJ�mR5Dc�<�K��H ���ω�:I���3� c�<��*Ҹ[���JD�ɔ)c��؂��S�<i1�%/|!����A��q��k�<�1-N6)@�0�o��;5�,�o�L�<�Q�:��8r��6:�2�c�m�<�p!�z��cᕮs���`�h�<�&�T�]�ଣA�.1k�Ũ�f�< ��-y�8۵G�-nRE	�`�<�t-Έ&yj��e�ƣ"0Q��Z�<	���\�(��񠒝l_��hp�X�<IӍ'v��9�7n/UJA��	Q�<�Ā[�p\�qc��/|�J��	T�<i����\I�A��+�nؚ�I�U�<�w啛k�A+�&L�8�4���P�<����)`��`a8��5jt�<�si��'S�ء���1{!x`{��D�<����0��0�҄Ho�`YC��^g�<1�,Bt�n!a��X�hHz���c�<9E�/��I$iۛ\�"}��bGc�<����H|�a�B�@��tB�lPF�<�ℝ�R����ɐ{��{��F@�<�t��#�V�IE*[�J=��I�<�q�P�	�t�j��
,Ǧ�����B�I�auQ��D<m<|���Pa`C�	�:��s6Y!�2���Y�?'"C䉓6����dKg!�񙇈�g�B�>t�H�$w�ԩ2�&��C�I�K�b�z���!�Z#�t1�C��8{b���#�bx8��\�?\C�I�>�BAx�A_�:J�b�MEs�!���h�Z�A��&+xm�D҄X�!�$F:a�*U�SfJ>!"��r���A�!��D�ڢ�P��Y��V�T�q�!�C����Y$���j��r��+�!�V�f9�]S��3�
p�Q���!�АO[��ڑ�>Bn��A��s�!�����RG"{�fq��S�!�_�G���C�T6ɾ9�2�� L�!�M��h�!���=~ʚ�b�ƮP�!�$E1�$]r�gV|�-J�鉻1�!�d��2ۑ�O`q~8�wH�*`�!�$U�2<D�H���(m���B��$o!�dB�@"�X�ؒS�dI�D�ra���'?����î�~�#čP��y��_��^LH��	�H���P�oƇ�yBj:M�9 e�E.C�|Șq���y��"Zt�s'C@rը%Rr�Y��yrb̓*ed�VL��R1�`!�mÍ�y��Ҷi1�P����3�Py�鈉rT2���������g�<A�l�#b�"�y4��
 �<�cp�W�<� "I�T�Ж�Ș���eQ"] "O�}*�H�;s��	6�Ē-Th�"O���ȹ@=���e �*ͩ�"O��ze�T-+���JU���H1�lx�"O�	b�E�W\��1百)z%ۆ"O�t�OY�g�R�P�ܖ����"O
ՙB���	��eӳ��P���"O��c�b��lw�%�2o
�N�!�'"O��dbR/&k6Rf��jBM�"O^��vLN�i�zm̜-1m��"O�������+l\,+��KM:@��"O����.z�@!P���bhUc"O�k��ĲB�>P���Q�  �Z"O|RtԖ�>;&�ݿW�B1�"O����L̢bK\��6l�5[s�X2#"Oz%�uǃ�x�ڴ*�*��Hn>L��"O�D�e�S��eK���bL\{E"O��꓃V�M4yEd3@M��Q�"O�RB�W[� �c�� �UM��#R"O���OD��q�@2l�%"O�@����9�m�!ˇ/r|��"O|X1�%�G����%1v~�Bt"O�1I�oF!p�Cf$��hn��R�"O���I=Y摲�-��.O*T�"O�Y�#Õ� VЩR5���j�q��"O6�KH��pE6��ʖ5���:�*O|d��DW_��u0퐰^�\��'��<�D��m��G��7�й �'��eh�C�h{.��#�g��5�ȓbD�2d<D����]�?�%�ȓA��F�Y�+͘��ZeI�"O�p��aR5	��P��L�$��d(p"O�s�b��P-h��H"]u"O �QG�^�V�������"O�BbJ�|w
�E慐 �4Qt"O��0aS$F�ҝx���Rm	&"O��:fH�'���ZQ�T�N���"O�)���E4IJ���@�AK��T"O92@O	2W�qѶ�@^/���u"OJ]!*�3��-��@���t+ "O�q���y�ȕ2`GRtp�Y�"O\z�h[k�R�
��C�D�����"O�p��g�{�(�э�)9�b}9d"O�d��'ɶx�đ�g-+CS�Q��"O��c�N�%-L� ��O�dˢ"O��+��� �|�:�k�~G�(g"O�ht��6��<�"�Ӆm�岣"Or�BFf�:Y�Zdz��R����"OJeBN#b`��b���Y)"AR"O���A�JL�
�a���xy��"O�q#e#�]ub��J�Y�"O���GNԴ|�D�@�	�K�
܃�"OiP���4(=Z�b��N�Jwla�"OnP� ¨Y=,�ǡʬt��[�"O���
`�\�D!����3"O���2�Z�(�`;�Z�s͌�S"O��B�
2E����6%D"�X�x"O ��`M���5�D��s���A�"O����Z�6�z���L��p&"OP�q�(��V=q���"OoD]�"Ol��MV�<�T��F	4�dU�b"O��:�R%�l��g�D	h� 1aU"O�p�`
�+i�(� F٬#~��y`"O6aa�)�%PJN= r�ЍN�U�"O� lq���ŉZ@�A��U���!3�"O�e�Ăأ'j2I�Ҋ$(��$"O�e"D���B�t[���%�2}�@"OX�S%K�:��p �� ��@1�"O�U��$�1f��u�� �(H* ��"OV�2�D�.K�&�)Q@�
=NI�"O0��bm�E!��k�E@�jTp�"O�1��3%���0���iH(!�"O"����	x-���f/[>�dEXC"O��Q$+Lq�c����1 "O:�	M�@LP�:D"�s�|�Pa"O`hKRc	�:2�DK������w"O��Sa�^�G�Ĝ�T)�0Xb�|�F"OX�2��%Vi`UR=p�10'"O��і�ЩwqJm{�b�6�ł#"O$���@\�'Fp䣷'X�$�+3"OJ ��`�zMh�ʳᐝ:@D`��"O���7Y�z�9�bܖn��%�F"O�`;��LK4�!��!B�n���3�"O��'��?	����GO1%���`"O��+��W6Pv)R� R�0�Eõ"O���oI=>�N5��Aոߖ��w"O�k� ��~U���%�R6F�8�iv"OB!�OO�p������1����"O*�Y�g1��pp'
�G�T��"O�Y�c��5,y��)�R74��ID"OV�t&߈8���@I8	n�Y�"O��A��1��H�?gl����"Ov�q�hʌZq�	�r�-0pFP�"O�K��7<�u* <]<5:c"O$�2�Rp! �3F
� X89ҷ"O�b��-O��"�'��g�j� v"O�-�q��\e��PG���< [�"O
� �@)�P��ՠTL�2h��"O���$]�(d�� s�G�*���"OX�!`�.��ځQ$��)�"O�T�1,L,KF���Gg
;����C"O.���BˮA�$��L;��K�"O�Ygh��F���Ef^V�lt�r"O|)��,ϯBt�ٙ�dы!�lIi2"O<��W+�,[�hY���R��z�"O�͚�`��p�L�;�ܠ���X�"O��s���5NN6����,3����5"O�}q�)ިN�Q�sA1"����D"O8���h�%�4�  �-�*�r�"OJk%.�)�`X�s(�Z��yx0"O:����=}�,)�G˷yJ��"O2	
#��7w������pD�lc�"OT��C�U97��9��!S t3t "O���$n0��mL�`����&�@�<��Yr�%�bnݧ!#�J�x�<tӿ8��TG�$Ud+�w�<3�%11�*Ǥ��4�ҍw�C�	�t����C�2l�I�!�xC�ɰx.M"���<}qd<i0	�"[FC�I�mtђ��4T �ʎ�y��B�I#;��� [��I�f�r�B�	�N�lH�Q"z��L�ڳ�͟�y�ص9����2�Ф_�&�+�ʅ<�ybh�n�R�k%.�T[9����yr���ko��� �)J��Tk#���y"I�-& ɠ��A����C��`C!�D�H�>I��D�7	Zhb�7I�!�dNB� �H`�[����w"�p�!�� �eI�BԢW��i�q��fE!Q�"O��R�g�`HI��7?@�"Ox����%4D��W�־s����W"OF<�$�ЄRq��a�A�C�b���"O�5+C+�py�à��+kVՋt"O�����^<v��`M� ��]�"O��E=��@�d"�tAY"O��p�*�%�xQ��(<vx��q"O>��F�1FC���f$%&X��"O\��VCL�C���D��To� ��"Ohtq�b�5;��u�ei؎`���rf"O�5����#E���!�#庭��"O� s%��?}5�$��f��>��$��"O����#��
#D�V�� �tJS"Od�QCk�� ��h�.s|X@zb"O��抔	p�3� G�T�"Ob 7�ڹJ9�9y��Q	 0�"O���S��L��E��"Y1Z�Z�"O��h���y8�a5�K�L��	�"O�U�p:j3�)��f֦O�v܂�"O�L�ץ�j�p�sQ�]ZD�p�"O����=	\�u�����g6��"O��x!�ۿn��}#B��>,L���D"O�Q�@�!	P���_e@F9�V"O��TᏚr��SG�E{�� (�"O$컔��b��Pґ��W�u�"Oj�aן<�$���ʴ:F�X0"O�1Bm�	 *���@E�Zh�"O譣� �>r
q8�xa~	j"OL�s/��{��h�b��@3^�(�"O0�k��F"����'!r(6ܣ�"Oʑ˴���|��򶇐�lƅ��"O�Yu*�0�4��p&ݲk��"OP�x6䜈h,��sE M��2�"Oθ�ҫ�@����ڛI�̠�"O��sD��.��8�1�у&W��Q�"O�Q@�	y�%��	�
0`��AR"ON(#5�A#Z�ܰ�GhS"/a~� "O$�Q�L��6�@%6�VL�ejp"O��j�ʩԶ����\@�4Z�"O�` F��Q�q��t|M#�"O.8��H�q*Ӝz��0P���yRGC/,m@)�V�\@E���w��>�ybG�K�$� �Нo=.%A�@\��y�eB�^���2�@��V]�X)!O�>�y�,J�~U f.۫S���8����y��1y¸qc��(N�g˾�y�h��	�ՀB�߀b(��gC�y2R'�d`䐢3p BH��y�cÔ�6L3�j��z^�Is���y넶]�j��Dټvb�򏝨�yR����S�����8T�ҢD��y�KD�u�2��&�HԮPJ2e�'�y��	.���g�M$u	�9���Е�y���7s��B� 2jǚ娡�ů�y�"�!m[���nS.!lL�@�F&�y2���[�(���`!lH��W�y�G	)�ڈ[ �KK�@���ؒ�yR�@�=�(@Ұi��9�������yb*��KąѤc�����yB	�	{1s��ǇY�����Y��yRY|� u�P"O���{���yB�Y�ps\̺��³2qa�Y��y�)ر}����0
;�����/�y
� |��`���B��[��	�NV�+�"Od����L�T=��B`�2 $2���"O�9T�29{Z�i��?V܀*t"OR��F��~�F��W��%r�BTs�"O~�c���
0�RP���@�#�"O��,��,�xm�D��
iȐi�"O�Y�Ą�<��c6c�lI<U��"O,�bQm��-�
��ѦCHрr"Ob���N��k#,�F8I�"O`�+���^�Ir�S�L7`9�"O�e��!ѣ���h	B"O��H��g�-���E|���"O~p����x�������.%�s"OX��LK#Kr�<��	7_����"O`I��`�0�J0bbO�FP�DI�"O�	����*��d��,L��"OZ���!YK����_!�4B�"O����s��&BZ�*<06"Oֵ#4��
�̴��e	����R"O��q"��\��9a3eT�A��a�U"O6�:�E�+pA�-xG�N ��1�"OxRr����v)�P������"O$���dVڍ����~��Y�B"Oxa��B()#R�� ���4�(7"O"m���*DK���'^�_���@"O��B�NO�`\�(J$�P`� hP3"O2��4kX�p�����7�6q�P"O��ZCeH��m���Cknt
�"O�!�0��2�pI8#�s~8!e"OJ1�j&^�<����h��T"O�D;DN[�6�V�gFn�p�B"O$��r�K�&�� #Շ�Iuj�#p"O�D�dj��7MZ�Q&HĢ7u�ٵ"O��P�N�gu<�3r��:����"O����+�0�P�*5d�=��"O��˂B�F�z��2�_>t��)٦"O��!	مh��p�G�KZ���c"O*�&�X'^B��!�g�;��ڀ"O�e ����a�p ҳ4l���"O^���mҶJ�QS  .
2�`
�"O\P�����&��%�p�q�"O����#�63�����I$m����"O�0��h\й�R�Y�WX�1"O�XB��Z���qͭ�����"O�����8�z	z5��,�6"OJ�]t�6ш'�%e'����"O�!�RqG��~���6"O�Q��c�;]i�V�U�+7�=S�"O
����?4Ԯ�)ШU�N��SP"O
�a���5s�l@H�N�;���"Oh8r(�}�2��Ȼ:�T<�"OrەLI �t��C0�*�0v"O G#� ���X�gן$����"O^(�Bz���H��J�y|ؙ�f"O2	�ÊL<f2X��6��?q.�z�"O���lN�z�p��7A��_2��h�"OF$�T��U*�ݤ- L��"O�5:1�P�����#	ƪ�#�"O,9��&N�2��ŬU���`"O��~(*��P�V�p�@"O�]�&�e-��3�W3 J�� "O�����4'�^��t�G�Q��D�"O�Qb�({Z�ECd�55�1��"O(��P�ˊ2�QR�̓uF:� E"O� B�S#���7��헊.����"Oʥ����s���S[����"O�z�O"\�aR���gn�Q�g"O2}�q�Ҥ�ZMi%��f����t"O��a�!�o��E�4�ٶnvQ"Ox\���I�.�0�C!d�3��p�"OR�q��"gN4�b"K5+�N�g"O���
��[������ vD��	�"O��;�$87��9e	�>-�pa�C"OL�j��P�(�$����<!�B�e"O�Uh����&��h��3ˀ���"Ob䁄@�B�u� �8y���"O����o�5�n)�0[�Q�le��"O�X�QjԟE4*��NĴ�Ѓa"OK�=`��(���2s��x�F���y2�Q�9�� �.�!d��1��[�yr��A�\���!����d��)
�'L��a��O��N]h��H�^D�	�'���	oX�DSjh(RF�5;\|l��'�dEZ�c�H�Ν5DF�4DN�p�'��@�G��dn���ؽ0tբ
�'J��r!	�cT,T3с�9r�I0
�'~:��*��b��e)�A��_a�	�'��m�r,ǑP�>4	0�$T�@�Q�'�:����8��8���3� !�'X�d�	�s踨c~r#�'~Q��k�,+�h$��#�%�)�'�Z����2[�Y� A1�X٫
�'w����HKK�:�X'��2l��'8�X�K1X���&�R���n�<9�����cD&R3�z�g��j�<�"��0x#����@���p��Xq�<�1�t�@e�ÅJ=�̬:A��j�<����2���q��D6y�"u��k�l�<9��әW) �H�8v��IbCfKN�<	���X��9�C�ʶ@b�y���FK�<ɠh���ͺ���4}콠�F`�<�U�ɗ%2i���W/0�`�Q�_�<	`��:���� KZ�mʢ��Q�<u,��Y�J�r�d�p�MP�<�4�A\�x��k��P��#I�<�0�0>K�AB��O!b��p8� H{�<�wm�i&� @��}|��G��Q�<��,�j�*�%"x��KS��P�<��n]�5�4�����	)jܩ�K�S�<��̗<�)��,WFC4ݚ7�RP�<Ii�'=�DiKC��CH4��/	K�<�RP�+6�i�d��Y`�!�1A�m�<aP�4�^U��@֓	����H�h�<1	�m�
��CL�7���f�c�<)׼%�iYVe<(���fK���y�m�8X#�tH�Ջ�R!�v�@��yrb �C%�W�<��d�2�Z�y�%\=�a�q�ą'������0�y�Bƙ�x@c�AHx��Ĩ���y�*]�g\����@X��	(�F��yB��;Sp]��;R�2� A�y��N3a�b��P+��Y�A5�yB�ju�Բ`�EbYIAG0�y�* �c��ɻ'�^0> �( �	�yr�����dC\�"Q�b�W�yB�M$#���:�"�o�~��T	�:�yre	-�����"R5o.�P��W��y�UJc�K7%J`Az�+� ��y
� �d
g��!$�׉� W׈)��"O�e�Ǌ�Vq@�S��D�h�@���"O�� ��A�i�Vف�
�e�� D"Of,�`N�Q̜`g�L�qXE��"O�Iц�J)'M�i�@��2�&�a*O�")�mޠ E�C�^Ѥ�1
�'�e[`fP�8��@U.0\:Yy	�':��`�Y�)���5�Q~����	�'CȔ{C-�zx�Y�ԧ֟)u�E{	�'�$��Q�E&<�:L�� #R��	�'Վ3���'%ʌ$�� +)Ȉk�'B	j��/i�D@����'r�H�'����"�n�Cq-^7�h���'�4i���J��W�%W����^`�<ɠ膣K��"�(h�t���[X�<!'�!6�¹kƆ�#>wNY`��i�<�Z&JI����6��yRփ�{�<�ӏ��NY���q A�2���@�f�L�<���:
hP�Y��S�yE����nI�<S���~s�A߸4ǆ���o�\�<1G�� Wa�p -�y'�\ �	X�<�W��'c�D ��n	���#V�<�k�6=˞ȱ��ǃ
Y�,�"��L�<n�4СԠJ�D�8�ÉVK�<AC�>�NѐP��/\;r��l�<��G"Pt���4jQ4ā���e�<��ɝ�%�� ¡�4���� ʋe�<1��#M�� ��P.%�T|���f�<�eF��g����^��P0�*Ga�<Qf&^;$(*3
MS�L�H�l�E�<���PV��)H�x�g�~�<I"N�u������<nZ�q��v�<a�J�)t�j1�С�c78u�ч�s�<���M�>_ DZ�'�"��r�i�g�<�i�<o���j��"�Ej2�Lb�<)G�ǈ'�h+gJ������W[�<�p�:������ (�e;T-�V�<��^�t�d��E�1Ue�@�hQ�<�b+T#>�q�(T�=���:�RJ�<�(�&:�&�j�Eϫq�2L1��E�<����:'��*1�
-Fi��. �<yd�� �-�T�ٌ"��P�Ôd�<YN_apRU�pH�0���HPc�<)�ڈD���S$�)/2Չ�%e�<q��ݿ`�jS�F�,�@��%'�J�<A�ؙb'�ӎ-!�A���I�<�s/�
�΅����/n�
R)�\�<	��0B�,EϜ�U�"W'�T�<	&n$?Ϣ�xר�J���rb�S�<�(R�\�j��1��9nE`�+���Q�<�ˆ��8а-Q� ����A�Q�<1��9V�� &�1�2��DL�<����4�ʠ�DƯ	�� ���r�<Au̛q�z���^�?T�'�l�<!ce6ji�y��å�����g�<��S�?BCe�̻5?���d!D}�<�2(��6(���5 9���r�<��Е'#�9JIZ�m>R<b��\o�<1`f̟}���Re���kr���W�m�<A�!]�=>l���^�:��Xa�BE�<���"+X-�r�Jk��Y�Ф��<��T�5�DX�W����Z 	{�<����q6�����5o@��P�a�<��	>����q��-$KĴ���F]�<� ^�A��1NQ��hG��<���"O�0�fKUH��Pro��?9�$�R"O��4'��bbL@�R�[�x���"Oi��m�ll(+��C�M���"O���uO>ZE�iQ��.F��d�2"OHy�l�_�漒�Uw�p��"O��R�A?/(�� �ǜ��s'"O�jA��:��58�4i�]�S"O�X#1���/�0���_�u�6�ұ"O@a�lÐs��@A�T%u|�)H�"O�AڱK�\���y��2c`��"O\9� 2%�rX��˹PD 9�"O��S�%O@��[)��D���"O�{�G�*T ��xEe�=����"O�ͱf���S�za�$J��]�G"OPɸ "ײ,O��S�$�C���"O`�2!/�%P{f�y&\6q0�"�"OQ@�<z�̸ACN&*P ���"O<�T%ǋ�Ȑے��5/N
��7"ON��J!lr�
�	R3r��W"O�M��!�kD�E�t�$�.-�V"O�5�KZ��$�P��Ӕ'v�d�"O����A,K�X�3	Ƅr\���"O&����Y(v��EgDC���"Oґ��*oF 0k#H��`�<��G"O����*=����g�{t�M��"O�T��J�y@��$@�#l�QR�"O�Q�����)ж :2�"Oj �Q��($���:"(N@(f�V"ORirD1r��鐔�ލnwx�"O��Ì��^�L�D g�q�W"O.����K�6����8[\��"OlK�bƸKoR�A�+>���"O�5S�J�;��M00~�LU�b"OD����q-nȈ���T��!�s"O@�s��Ҡt�Ju��Z�����"Od�ǃ���
ȺL�+J����"O�ܚ��,,��}GL�>���b�"O"p2s��x��@�py��:�"O�*5.�>�*c�i�����!D��كJɬ��x@�)�1*��p�Eo$D�0�D%0,�&�ȡm"(���G� D���h��	h$�[&���|֌��p* D�d	��ԍvL�O�?�<�c 2D��R$&ץ=i����
Z�X)�s�"D�D��뜊J��1��̙o�&CƏ.D����B�&J����h�٢ra8D���� o�>�[a���J]�`:@G5D���CG� ��QY�ڇ��MY�&D��P���%-+����{����
$D�ؓQ�u�`=�*O�\f����<D�,����-#�����L.H�bQ(��<D�L�F�ph�ဆn��Bd�ѳ�6D�8.=���A5C�;K���@�E�!��U�D|ㆊ֡HW !�@lê�!���%1g<�@ב|9.MHR����!��M���.�L&0L��*��h�!�$GD�$�ň��{E�� )V!��t�py[�b�-FkH]RCh��\j!��;��,�wD��Pf8�[�M�5K!���.��pN$c�����%�!�dƥ:OХ�F��;fV�1�IJ}�!�$��{6|{6d��:��u����i�!�DH�q��=6nU�L�
��xU!�� r�3��J�
�`����Kn,��"O��˲	ݰ!�Vd6�P$u*pp�"O6Xb���w��QW���!<��	�"Oz�r���h�j��$�&.8�@"Oڝ����D�D���"J^T*�"O^��ŏ�����"�xؖ��f�<�e���:xrTMJ"\�K�g�b�<�Uf�:����T]-$q#H�[�<��F2TF�L��+��K>��g�@�<1d��%)� �J�1r�ap��U{�<y�+�H>�d�g�^�\fx<���y�<a�/F�<�	����y������_n�<�U�P>�B;0�Y��0 �o�<�Ę=5��iCb�Z|k� Yi�<)�!�5��%�����Z���Ŋb�<���#7���5B��\mV͓��Bd�<)�,��d�+`�Ե*�Xp��^�<Q���<� 	��iö��0C�CX�<����G\)k2d�5r�f��v.�R�<�w�}�D��R��2t A�AD�<)@A�(|�Ԅ���ߧe�(&�}�<yc�.2+Փ� ��>}�P�u�<����b���{��-_�ܴP�Xm�<q��]�.T� rfN��`S�S�r�<ч��c�2Y�7�'9�6i�Αp�<�C�:p� e��X�� ��UA�<Y�$]�b�$�x#��Z����*T���1�ϥF�9q�bH p�����M=D���!Ǔ�G�$!��-�=Fv��gB;D�9���,�`S��-�x��%�;D�\r�F��	�V��dj	+Q�-�e�6D��HF�P%Gȹ�W ͝T��p��4D�HG�'HԬt����>rܢ�)�b.D���� .A�P�8�-Id����+D���!A����.�#DL6�� �+D� ���U����H�e�3 p<�D!&D��KAH�b��<��'�!�80)&D�d�TJ��''8Q��b �h�޵R�*.D�$Y��&`m�ACv����8D�����W�=��ym �'���d*8D�8`fT�pzް2�$��Pi�� ��8D�����bu�[)���� 7D�D��P�o�T�2�3pF��3e"D�lxV
2!W(�����c(�YB�� D���҂ך$�h�:#@�l��3��"D� b���\=0h�F��#Jr\	"D�����$�Bq��%-*l`���!"D�`�cN�q��<��E��uB`s�<D�|+� 	/r��E�]�T�{6�-D������I����(��&�<��2#6D�H�K�\3Bis�t�bikU5D�dA P�0���� �6U˳!3D�İ7DB�ImCL���B�C/D�Pa��I!����uJ$���cUe'D�\J��ud��#H� ?/xۣ�2D��4B �����$�5Q�.hSFH5D��!ր�lR ���NƗ?8·�.D���-�3-pι��(��O�@)*4 ?D���R�ʖpJdp�nY�"P�>D�@31�V�h��)�g�D�1�e�"D���7��^az���iͷF�UZR�!D�Lc� �*%dR�{�� �ZEB��!D��{2ğ3�(�BVN�T!�&#D�au�ՙK�|9;�Iӯ���@��=D�� "�!ä�TXq)B�	nP�X� "O�d�
�D��@rF��dQ�R"O�Tӄ�F�$�M�#&��X��9�"Oz!:�j�<��R0��!�"O��t��*�08���I�%�d��"O�u���Ҧ����H�*��-��"OH��R9o�x��aɂ�w،` w"O�0ө��j��Wk���=�S"Oʙh�1k�H ����H9"O�|�p�J�+�nٓ�� �
e�f"OT���	?2L�XU��;4���"O��x�"�.�p�����""O8yڔ�V�=NX�`�Y�{�"Oՙ�b�^X����k�@�h8f"O��������t�B�h��Z
�"O�X��r�طi�'		����"O��1���R�Mr���*H��P�'"O(門�&a�{�( 8ow4�"O��Ca���2�����	�de*q�C"O(U��aQ�]��,k
�	�y��"O�D@�M����"E�"@yS0"OL��d�B1��d(��>N���"OĖ�=S��Q�nd��a�!�yG�a(�d�&�9z��w� �yBѓ,��"��Bo���al�y���$Nl!�����2���Q���yR ��O6�a!G 1`�1�!�Ӣ�y�F�)t�t�8^��9��D��J�>e��u���9Si3Z�1��-��}�ȓ$��iY��n�  
�?'+��ȓ�.|c�g%]n�Z�F�#x����s��{!ܾ\�[&�A�r���ȓ)*��#l��T�^�v/kȄU��v}<�{c$�-eS�p2�OYm�.��bْUK��ŭQ|&5*6LK5*����;޸�!	�zQ|tSq�_-5l�����͸ч�.��@3#��8�>��ȓ�|A:%#'!@u����,��ȓe�P��d؍u��1"�豄ȓ`�DeA��mh��ʁa�0kZ���|N�i(
��ڄ���V�܇�r@��
كt����W�uGR���-ܫT**�p��,	�:�4���1�vu�'L3CWx10�S���#�l`�G%��B 8¤�$���k�l``��U)$��ii��Q�A
�'h�NO�A���p]P�s��y��X�rFi�c��k��8�C���yR��n3��$�� �"����޾�y���#�ʵ����x�+��7�y����ȔC&�J�`�K���y��\i��AO�++4�ʤb]��y�C^3 ;�-�WKW�cDe�W?�yBb[8|�U!�F5U�q���]��yb��!ȡ����J�K���yR�[�QԬh�W�D&] 2ib�N٣�y�
�\:���E�_:U�ȅ@�@��yB&��'��!����9=�:x�S��#�y�g/F�;��\��핮/LH��'~lB�ʐ4#�TJՍ�3.��
�'�Zܫ���5�4)��[�6f�P	�'Z��qb|��L�&y|U��'C�� ��ܞn��Y��o�_p�y��'��H��M>o��Hx#D[d
R
��� �X�)�+tr���>t$HH�"O����@ux�ZV ��}��G"O��[�$�\=)!�[�c�8 #"OT�#�,pA@l(�x����S"O8��ȴъ�s��:n~ջa"OM��K'Z�
8 k�QV�	B"O�(�bf��1�Xpo-:����"O����K�:$<\�2���8*t���"O�9�ç��@eڑR�߉U�`��"O����k .nX�Zp�� �=�""O���!@�d��`�B�e���*u"O<��MPQ���c�!φ!R"OH�2\�8il�0���q�\mrT"O��uAͫ�,C��ͤ"� %3f"O(,���]�q�F�m�,�p� �F'D�xC�'�2�*L
Ԃ�u��&�'D�s���9Ů"�Ɂ6T��ɛ+$D���1�м?��� ���5�$�#D�d���e�^>g�=�����I/D�XJC� �8|�@�t��pavF(D�8JCH�<�2�0��r��,�f&D��:�&��G������S(�4s�+7D�DЗ,ђ:g�d+�L�C��h��5D�l&N��@�8�"N�+�8�;��2D�C���X�!%k�� ��+D���׋ 6Y��u���rc�I�*D�I�gUB,��p�U��5�!d&D�P��L�mqV|x� r�px�u%D��X��&3�$SlǵJ'��i"� D��Վ�k2��J�����P�9D���NM+{E��i��b�|(!"D���Q�ɈN����
=<�L-"�,D��z��C(R�37l�:NB�H��+T�Hr7�҄'3�P�Q ���j�"O2��s�O#���� ��x��&"Ot��P"�9j��q�O��T~�=s�"OpI1u�ݾa��j��	�mm0�"OX�
".d�c�G#[p���"O����� +�)�aĎ4Xzh�p"O����fP�#=`��Q'�F���"O�5+���� ��aI??R�٥"O�����ǹAO�8Kg��?����"O�;�`I�A��(#��K�񆬈5"O@M�E����aK��Z�2��"O<�zVF�w[���Pa�ʌ��"OL�h#,�0�X�ō�h�w"O\��� ��ɂ���LX�:$�S�"OZ��X:Tta��0}����F"O�9�A�^��*L3�f��c���!d"O��"I�z�i E՗��1��"O��A��jsD�A&�w1�<�q"O*I�l�4� ��$Ț(���!"O�D@�K�9An42�E�Y��#f"O�q�vb�R3���wĪb��, �"O���%
�cg�S�d�yU"O�02G��j|�`�vK�Bi��Ô"O�FDP]�r0�����OP��ar"O�@���E���ӗɕ�
�\�3"O���M��=
���$t�����}�!΍<�`��[�h�bԄȓ(1���u*ОJ*�x[2@ ����ȓA:��ⴤ݉ �$�Qo� �6\�ȓI~�HS��f|��F�]ca�ȓB)ƈ(�M���%0����.���S�? �ɳ���&�,|jf��99#<dˢ"O����(6�5��g�*>���"O���W���X@��e�3��B"O8���JԼ���X��'2���P	�'�z�J���BU�� �^�]�pЫ�'1\��aH�?�}rq��4W��Q��'����DgҰ
���l5Ya����'������fzlh���YR�S�'�p����ܙ�8��ᄎUX����'` �;h����)z�RIeY	�'��Z*C:�N��"fS�Hi����'�2��!¡��`���i�����'l��5C�
m�ȹ��*[r���'��	�QÒ�34�#�"U3X�Ԥ��')���D��M�R���$�Ҩ��'|,�S����h�3���1R\���'�T�[b���U��H[$JX��'�:ĻӪF�h	`���$��
�'���Q*?9����%�$���
�'���3UI.e	�K��g���''p���%֙M�޽��kV�2�q�
�'��]0��Jv��y���M�h6�p�
�'�����r�t�K���\��]I	�'
�j�c�E."�y4�,?�����'���x�kN7$�<�j�
-��@:�'�м!����H�{*٦�	f"O�xf��*nI��Tnʐ&�J�bE"O�Ty�k�4Xb]fm�2@�#C"O��!�	Yfx�����l�2ES"O���K�8�������m�D�Q�"OnT�r���'�ݎow�U�
�'��d�2B��~GD��S�0C����ڢ0���6$n��C_Elh!��J��� ��}��C��˛��rh�Râ�N�Q(�Y|��ȓ[�,q�w�	������\$_�F���7\��!G� %^��@����6���#���� �AsV��%X��n�ȓ|���̎Y��-r�AsV @�ȓ] ���L�5t�9RD7��\��Ga��u�ݥ>8�\�iEp�X�ȓ1T����I��	5z��#J<��ȓ^�$�����K�~�D敠\r��3��a��� �c�e@�ѷ"�dy�ȓPDq�I�)M�F=��N��:�Rd�ȓ���w�'J:��D�j����&�HD�Ҁyz�cC˼'��ȓ[�Ɉ2D�#}�Q� �2�X�ȓt ��rtǋ%����n�����O���;��Am��!P�Y-x��ȓ# e�c�%��Ʉ#'e2чȓ�#!иqGbL�h�%TQ�<a�@
5�D��R�QŪ[N�<f(קf���[$Xx���+�^�<9!����@����Eޜ+��LA�<��-�T�(��w�z�c���R�<����i�t���/� 9R@k�"Fj�<1Ƃ��,���mŜp��k"�d�<����7Th�i��Fy*�RtN�l�<yG�͋r�М�Lɳ80�yqN�e�<��n���e��.;�l@A��z�<Ɂ��05����2�yKeA�x�<Q"�֙t�����P��sIt�<�,TO�ȃcѩCh�X��h�<� 8](F�1B��1��ٿ[>Z]1p"O�+v"���ͣ�#�W&�� "Or�x��P�U�p���׸Y�i��"O�)ԫ�E@~0�a�oN$�"O`�qGX�X�����!��1���"O6�;DB�9���"�	xy@�i�"Ofaᣅ�;m>0[ ��6	l�� �"O�I��M���Y�҂�,wx�ص"Oh�����J�q���Hf�i�"O��� F�m{.䨖�*Z4��9e"O8��!�qv��1�L,23|鐡"Oā�G�;Y���)H�sP"O���.η'���#`L�4�rDs@"O��ش̗z4���CI�iP���E"O4���oG�&���R�@X4Bf"OP��sf��~ꔬkUg�
{�C�"ODh�R�^�r�4=�B�O����"OP0�
@�}At\IGÆ��$s@"O�;F���J��P�\�M�`�� "O@P9�b��Tj^}��J�$�@"O�ű�ƙ)�ĺp ͙u�D�"O�����<0m&A�J�V�D�CD"O
�jg"ώC�L��0i�0D���t"O�4rC A��#���:��X�"Ol�8⩇�Xѡ�W�c�����"Ob(���Zv�M�F4v��+ 8O@�؅�I�ͮ��
T�̘ѠI�.��B������BĎ�Ç 	�=��=�Ō+D���P�Ȳq�$�2&E�.���`ꨟ|G{��i�*5���	r%�A&�0
�[Z�!��)$�����)<ص�g�ʥ+�iF{���'��ʔ-Y�3�M�&�K��	����a�\�gS/��y9rhX5D��Es��,��0<����q�@�Wh�N
N|�`�C(<A�4X��1�c��>{	�B៰�(x��F�X��쁝Y�Ԑ��H�&9����i�<��)gVХ �>etX�Am��D{���i[<P`Pa�Zl�8G��f�`H��F{����<qQf�1�Z8�>�Yv�O��M��'b@�BO��!�
�C,˞H"2� 
�'D4���"���p�ƂxX�Ī	�'(�v`�m�(艓��v*�����є�y�,�'��qpG� 9�TC#�O��y�@��NE�𯈷}d��1�aS��yo�#v��2�mT*+�z)��y�l�.=f,m�3�F�&->�jr@���yr�'��X0G1aLi12&Á���*�'��*qW"M��dΔ�H݀��'rz��[ꌐWn��}���s �W�<�Ul�@N���C�:�Ek7h�ē���~�N|���k�N@�+Ϡ����]%S�$�'<�}��.Mw��
A�;;�e�f&�y�G'bY �'+-�l��6+S'�ybIϛQ,>�6�o��,�E-ޏ� �=��V�%�֝�?J����:��q��_�oO
B�	�dsz�1��$�,E�f�I <F�B�	Qن��@K���b�cH2vxB��x����0cD� �� ����8w���>က�F�ypB D������\�<1f�ޮ$$�$㠯�3��I���W�<�f	G;s���9dDUx҆�Y�'���`�Om ��g
˟	q�)a�i�6~���'�(I�(ί+m0�p���<z��(�'�<�p�&Vo0Ђ�LY�r��0���� L��q��.1*,���5g)<`�iU��O%�S�O]��q3K�8D�Pă�����ա
�'&�p�C��uK>l�D��R:`��N<��'b�m+�J�w��u�Ch`)s�yB��C
�y�N��qC�= 3�!��E�E��y"�ݔh�(D�!A����!R��y2)b}���L�$#C�y�@˽�<]�v�N�]�������M��'�ў�|z­F.rɪ�V��B@�]��D�e�<�ЍŦQLZ� �@����g��j؟���'-�]Z�	#e��g`R����	�y��'��y��.Ւ�+uE�Pd�H��yR�ՙx�r�P���zĪ�8s�1�y�*ߞv�p<����ly��1���}�ў���O��c*\�=�������@ d���<����Dń��7�Zru�a���'��:c��,5��*�&	y�P�T(9D���7 g\��TĆ0R����lz����7Olc��qde1�*�
D (ٸf"4D��SR��|9�����8AV�t 7 ����	4<c�Ԣ�LX�m�X���B�)D��1�?��Ş��9OX�ֆT'N2)�'�S.p���{w=O&��yr�'#����${�\ *����2嶡ڍҥf�����c�h�c�4\!d�C�!�D��
�ӳ�{��(�&-���O7�������' ~x����EK�,ҕ�� h���C���j���� D)I�`�S�*���烜[�<)ׁ�5;J���L��P9(��B�`x��DxRB�013ș�����G����ύ��y�K�
8p4̠�`�CN@{�ǈ���'a{�	 `P�C$�48�8��7����0>�M>鄦 
f�,!�\�n�r��l}�P�4$��9��C�O]�����
nJ�U@�E�6/F�,E��H�5�<) ��6T�Z12���y �S��� b�#@�\�sd�)�yr��<m�
9��
�=<�j�����y��
M�:�CK	�=�l@a�E��y�K�
g`���T���� �Аx�G�){P$�b�	8����%�T.Z��qy"�|Zw�Q�X�V�փP^4�y�ˆ��<Zd�2D�X��)T��@K�.T
N0�2 �+D�@���1�����G,/j�H��'D��a@h��8�ap��2z+j� 0 �<A����$L���U*����%W�6�B�I����f�ȯ.�F��P�y��C�ɕ"Nl5�&�ђs�F�d�zPU��E|��	��;�LN�G���AF��aȪB�16��b�E^�0`3iU�vj�B�
\8i(�'��}�Fٙg�N�@#>ɋ{B�~�g�+]3���%O��8��{�IBWy��)�'�:$�Ț�Z���9F���FO�͇�g����&��[���ق���UƼŇ�e�D	�΅��,�B)ZQs:��'�~�� [�-�3�ʜ�J�%� �yʙ%?�V���|�&H�5e8�y���)&�c7�΀{\P8;TΚ��O��=�O��͐�(�El�
�I�A�.�Y�}b�ix�T��D�2�μ�e�E����)�F-D�@�	����� �D?;�(�!D)D�����Zyp �{u�	�򔢄O:D�t#6�s&�
i�)�$�B$c9D�DY���7F��;�A�9L���X��1D����F�$�)2���{�̐��/.D���W�Ց9�de��#��Zf1Z�a9D�� �5`%��8_D%i�G��!tr�"O��I�#� _�d�����&�Nm�Q����� o���'˚Y~E!��n*�#?ɋ���"� �yr��.Y�@� "T�!��V�
��a��Ȏt,T�xV�H G!��O/j>��6�D&HFQyG׮I0!�d:<��b�E>��sDĜv�!��_�[��bf��4%�����T�2�!�$	�9��=�'@Տ^F�a�G5]!�dB�����vɞ6n�&P g
Q�l�>�J>���]..�M�C��.$:T8p����<a�䑄`�fezm��+rZ��f��z�<	��*]��q��د ��ě6nK�<���M�$�!�m�g�����K�<iE��L�$,�� X�zm�i�F�a�<!E*L C캜�Bʁ<P��@����x��!b�6��˅h��,1w
��y򊘟jT��pB]1q���I��#�yR�Q�>`�Y4�ؗX�����,� �y���B�q���S��QEOO4�y�����3��V-G�����F��yrH7T��8S#O�A<v��C�y��0Y�d��	�Eoڝ� #�y"F�K
�YP ��4>���P�����yFߛ.��*��W�	�Y���ʊ�y2�]�}�:J�OЖ�갤õ�ybD�>h����%�N0H! �A;�yBlԿ_f�A'BP5h|�Gh͢�y"E]�L��\[n�u�c�N��y"M�?�Լa1MS�Z P�K2���y"��'��i��͋�V?��W6�y���N�Ĥ�iߦFn$܊2�г�y�O�1VZ;@k�(C����1�6�yR���	�TE�fE%T��̪�yf��}���[� @.q����0�ҍ�y�Hf ��9���p5Ju���-�yr˚'�l�b�J�
pʚy�C�	�P��][�$�D��e�/\RB�I��⡺��LK�a8���'�FB�&X��Y.�88��tb�O�]�:B�	�w��؛qn�=*���M�Gq�B�I�<ͼܨ"�بJ�vl0a� 	@��B�	�}���$K=\p�c���O�BC�	.�y��ƃW	��*C�ݤ<[>C�I�G�D��Y=?��$�U�ܒu�"C䉙-M&��'�'[���9��T�]C��@������T1�ץ�T�|lh@"Ol���O���y�%�A d��3"Ojd'ӪG�L�BЌfX^��"O��)B �p'T�C^J�4"O��`�dG(,��`��Ĉ�c4����"O�(A�(A�(#�W4K&�8�"OΘR�C��X^��ɆL^/,��"c"O���[�f��j])pv�EQ�"O��z �;n��h I�?j*8�Q"O�����W��l%� 'SfPTXC�"O�rV���\@0�q�+�l.���"O�Q��ŉ,0�b�HpJ�u�!����r��f�ކNV��z���1O��rQAX�KH�:&ܳ�"O49W�ʓ^��t�ƌ�9h�ڱ"Ov�RWg=t�
�a��_�xH��"OH4A'ԕj�iᗂ�4w����"O�� -�?�VX���ݤ+d�eZ�"O>��蟰64��EeX �;�"O� H؉�"R-s�vsrG6oW�U��"O����[�]���9q��U��"Oޭ���J.ֆM2sAI56��R"O�h93�sid�{6��4tf��"O��3P�Ff��2`n�7Ah�i!t"OzL�w%�F!�q)���F^~�"O�Z�,h��,WL�!"}�v"O�d�aՠM����a'�
�"O^����^�q4�-��Ǵ909��"O�@�3�7	�x6�ʥ7�L��"O�\a��I,�-	Ҍ�h�XTA"O:�ÕD�	ӄ�S��!s�lq�"O�@��nf�(K70y�v�Q�GJ�<qE'�>x��5���3Oi� B.EG�<q���"]j�g�>}��/YH�<9p\�7N蝐q(��Vl;vh�	�hä�Iy��X�$�F~�NPm�5�eU�n��Ť���<�%�� �h����O��E�i��Ԃ���s:6h�v��v��݈�	̭�0?	ծ-��=�5��?6�T��� q�ɱ~o2�X7�A	`��1��Ø��ӗ&S
vw�ӗ�4	ؤ�d��@�흨	�C�	�F������\�pM\;���Q��̀^��)�!	O$�̽s�ə���¥[��y�j�n"1�y�ђe��\Ȃ�B�i_�l�1���xw��B7��hƬ��:h��a���ƈP���b�Vi��� f�QiM	F?��Dz�I0\�[5Cظx\HK5�Ё��x^LS��9-�6MA�p�h(S�ϊ�g��0gc�`��Ɖ�TE�I��ӌ	��:�-G�m���s��p>��g��1,��4��2]��qM�[|�P0��I��aC�^#ؚl���A
7<���m7T��͈ԼS�B�LR,�z�A�=$�`j�+1�(�4��5��ѣ dSr�B��=F��f�3~�$���?(2�Q����e�<�wK�
u
�Cܔ<G�)�fM�{�>��P'B�}�ʥa����I��$�"0ɇ͜�w~���;����O�DI,�p5�	�o�H�:�'^57c�%�צŕ3A��`��ft�m#��yhT|i�	�@�\�R�_62j�=���4H����'�LI
(�!4��,7��\I6 p�O8�yR��u��DH`�(KC���R ��4K7+����Ҵ�±&�j�`���?	�}��H�lr:(��2\2샀���8�Vg�3"�x�����O�E
�HX>Nw���!B�V�X.�&����d�#b!$J�*E�4�Q*ѨX�J}�r&�"E�N��w��uA�742�ˀ�A�d#]��`�`���d Y�g?�7�	 �0ц���C��j�+]5 ��� "Lh��uA��R��u3b	�/��V��G��z���6(���"�|u&��D�#��@2P�W=o�1���tC`�yRHM%�~�'�Ժs�L���g����\�a��3 4�B�ǟ>S���F��O�z�;��B�6~��u�N
d�$�(�7$�b��߽T���&aN K�d�{S*Gk��2��"U�.������$ǅV�s Mzv�߇V��D�'䘀F�jARG �&a��I5h��h󤨛(��#�S�l���I4J����A��:v��Yըד}��H����1��(��!�5W`�8�G,6��Aq�O��xCe֌2| �b�.[�X�<�0��3Z~�P�ӯ1��	�5�V��Q�V/F����K:Hq�u� �D��H!����:X�&I�0��SV-B��K������O@)�c�2,7,Ypӊ�<�X`P� ;(z��Ó�3�İ�P���M0�ŭg]dH��֟�\p@$U�j�4��gn߱K+\����I�� A��8��N#R���x��<e�V�(��R��p�Z�^���AaW�=�<`ആY& !:I�%�ʘr�ˣ,�Hg�Az�b�����fݍ��,�Ml���O�zm��TW��R�S-D? QYЫ^;]z�Z�xP��@�<u����bj\�h��h�$+
z�K�KN�+����Z�]P��`��N#GE�ܡH	2�q���N�E=�$Z$d��?����0C�7XY��,Ow����40.���L��y��Pȡᗐ7�d�IG���.�Ti�l���떒3�p�Yg �*�@]�����'T�.��٫5`��e���+�&�?��	����] 4��X>ӥl�}��$�@/^��O�ip�R:5_.�Z���'NN�ZѤ�&i�.�C�/ �� "D(@0Q��i`�p�% @�F��x���2M�V��(F�|	�⁤r!��+l�,`��	c)T�L�#=�OP,�D�B�7Lb41%�݆*����,��Hޢ| �^�"$2�0�&C�8����
�a<�!bbC
l(��3��8I߾p�_&.$�(Xw��Z���J�����[i@��4��}����'І� )Ϥ'�uq�H33ܠA#�mI<��l�ݺ+�I�7�H����Z��,����:��/9]V�]�ݴD*��a��9��hgk�:n��qt��Ϻ���N6y#��Z��I>m{��`��;D�mppB�2R��̋f��cqt�;@� (�'=�H(��\  �,<(�h�fN�i��+�,^�Ip�zĲ81�	��m� ��% {���
�V�va����.[qO��M�0�Zxȵ��V�rk�<���I��Y���8��T1.�&�͝6�FD�5���R�ZwF�lr�G�)F����	fN�%d� h²��4 ,�X�1�	��j�p�I�v�>�R� T��IU�@?RM�d�J?q輒�/�V�Ke��L��H�C��I��Ae���T	}��o�;z��$���Q��6aH�LtʀF �X���.?ᴁM�:���ԟU�6,)�b�K�� �ς
\�5�P�� ��!��2�@`"֫�t�@�q��Ӧ=�T暋K�fQ�Bnы7��Bg�No���t�W�*��@sjѝ!�ZT��HܷC\�j�j	�)L�����D�h��a�A��r��P��D]��R@���6EL�:G��.C���ٴI��<���͊a�lH��	��P�槍ZB��hvlGR�R���͗nu��E��g�r0(M<1��(��I���e}�Qдc%n��,����%=jiI�G��M4�e�6�)�7��.*��\�)F6O��m)�C�	3�0R6"�:dXD���Κ@=0hѐ#��a+ܸ�p慔+��L��a�a��+R��i3�ǆ,x��,c��h��h�=�7I�DU!n�m��h�?�3J�CP%k��e��h�=�9E�IX,c��>�#vu�.
�|╰=4Ci��<�#vu�.
�|┲>7@j��?� uv�-	����91Da��6�*|`��L#�+Ŏ��?6�/�/�a��@)� ͇��26�"�'�o��L"�)È��:1�%�"�j��X���D�LX[��S�[�[e�Z���A�I]_��Q�Z�Za�P���H�FSP��[�^�_f�]����Mdr��X���Ƹ4
K#���Doy��\���˰<C%���@k��T���ʹ?C%���@k~)������,�"���F�����)������$�(���I�����)������#�(���H�����!���@B�[&U����߫@���GG�X"P�����׬E���GG�X"Q�����ѫM���O@�C}�1Pݩ+��=r�=VH�֠Fx�2T٤'��8t�;SL�ԠIu�:]ݧ%��1z�8PO�УKt�y����nZ���/5ؙS�����nZ�����)2ߞT�v����i^���*2ГX�r�ԟ�q&��p�gL_����'\�-���r+��r�bK[����/T�'���w!���bI^����-W� ���z,	����k�P t�Yh?�,������`�Z)|�\i;�(������`�\+~�Ql8�+������a�[�5���*=/�a!yç��i�]�0���%0-�g'z��·l�W�=���/8*�d%z��¶n��OT��"R�"��y���DX��%T�%��v���G_��"R�"��y� ��D^�
c��7�Ɵ mѧE�Þ�b��0�̔-`ڭM�Ɲ�b��5�ĝ&lѧG�˒�h͊g<�����
C�.hv���`=���
E�/jw���g<���K�,it���n7���쩄�[k��Z�a�ϕ��宅�Yh���P�l�ğ��⥏�^h��Y�f�Ę���c�dַ�^�8����Z�>�+b�eַ�_�8��
��S�0�&c�hٹ�X�<��
��R�4�!k�b�];�aVT���6H�Xz+���R6�k\_���?@�_z/���U2�jZ_���0M�_}-��� ^?�f�=���� %����؛�O(�6���.)����ڛ�O(�5���&!����؛�O(�6��x��Z<@Z�� �v��\�q��R9BY��/�t��Y�r��V2OU��-�p��]�p��WR�h����#���	��h�R�h����% �����i�R�h����,
�����a�Z�n�b��9�~�h\���0�g��:�}�oW���<�`��9�}�nT���=�e���׭�EՎ�as����	�G!��֭�EՎ�cp�����J,��Ѫ�CЊ�cr�����C$��ߧ��PR��c'�������}�XZ��k"�������Y[��h ������~�ZX��+�O�#�e���A��@b�'�G�&�f���F��Mm�-�F�/�i���@��Mo�(�~O���f؁C������5�J{J���cف@������5�J{J���bۃB������5�JyI��Wh�4�"qs��H��%V@�)_b�;	� s��F��)]J�.Za�8�-s��M��'TA�)_b�9�$��d���M(�J�}R��$��d���M(�J�}R��$��a���G#�A�uU��&���f`~A��y.������(� ���ae}C��x/Ά����"�	���f`~A��|)Ɏ����%����f�]c�"z@�;��X P��b�y��]c�"z@�:Ó]X��h�p��Uk�$~C�8ÕY P��a�~��Vnό��'j
Ȁ������g�u����(bυ|������m�����,`υ|������m�����l�pC<~9���)���^�)91_`�zI6t0���,���X� 0;Vo�wK6r4���%��S�$3:Wi�xJ�¨�GK_�u��Se�����_�ɤ�LCU�r��Se�����_�ɤ�MBW�p��Se�����_�ʡ�UÀ.lb~������ȕd�%`_ȋ!bjr�	�����Řk�&fYˉ dh}������Ǖg�#c]ɋ#�t�>y�B���t{��V���t�>y�@���wy��V���t�<z�H���xu��[���|�B�M�#x*�\�-���L�}B�M�#z,�R�(���K�rO �I�!x)�Z�$���C�pO�J�L��qO�����NAHLWm�M��qO�����DJEAZ`�@��{E������L@INSj�D��[�A��tB����*����OZ�A��rD����)����
FT�N��wC����)����	BQ�I�pNPň`*��ܫ-^|E䒨[ςk!��ܦ'WrM뙢X̀h.��آ%VuH疥�ϣ��s����/�kSA2��Ǯ ���x����-�kSA2��è���p����/�kSA2��ǭ�l;�A�w�5&3�������*�g1�H�x�8+>�������.�f0�O�t�4&3�򸛹��-�d2��F��?]���֌��m(?=�3�F��=Y���߆��e/:9�2�F��=[���؎��l%03�8�KΩ.Wj����Բ���X!Uj����׾���Z &Po����
ѵ���W .X���;���L��Yb���{
���;���M��\d���s���0���F��\d���}��ے�^����������ƌo�*���^����������j�*���W���􇹎���i�-���Z��Sj��M6A����x	�?�Vl��E?K����|�2�[b��N4B����r�<�Qi���3�+1۷z�U/T�\%��1�$9պvs�R	,V�\%��6�.5ص{�U/T�\%��6áh�G��P�x@@赭k�-��b�N��\�z@C⸢i�/� �b�A��W�~FD㿥`�%�
�j�D� ��/vc�n�~�9J���%}n�c�t�<I���%|o�a�w�8O�
��׺��7��0=��`~m���ݷ��:��;4��azj���Ѽ��<��:6��kra���شo�F���}횵��}�� ڮ�i�E���}횵��}�� ۯ�k�A���zꜰ��u��-ץ�a�@�'������;ۿ�ɤN�3 �������3ܺ�˦M�;	+��
�����0޺�ˤN�3 ���N���#�g@j�,�EMA�M�N��� �bEo�)�@EK�@�B���&�bGb� �JAK�J�L�����`'� u%�<�AK�9���j+�-
-�9�AK�;����`'� u%�<�AK�;�����M�(p�@d��L/��My�w�F�%}�Hc��H$��Cq�t�E�-s�@f��O,��N|��M�(	�"�y�o:���ۖ,�(	� �~�e1��t�ӑ)�(	� �~�e1��t�ӑ)�)�"��H�xĒ<����ݰ(�,�z��A�zƟ5���۵+�*�s��M�pΙ0���޳#� ���D��O����j�<�U�,T��o�J����j�<�U�,T��o�J����h�9�]�&^��g�O��|h�Zg�8��)����tb�So�=��+����~j�Vk�<��(����t=��u`��>�B�����6�d=��u`��>�B�����1�l5��sc��:�E�����1�`>��A��%���Z����N:�~G��"���R����L9�{A��%���Z����L9�{A��%gU8����l��f�K��^m�UcP?����h��g�H��Xk�QaP;����l��f�K��^l�VgU:�2h�˚�jDd}B�X��;毒6n�Ò�wbCczE�]��9篒6n�Ò�wbCczE�]��9篒6n�:ɹ��r��!� �Ԕc�+��?;��t��$��֕b�)��:Ȼ��v��!��ܟh�!��?̸ $��Ҧ�p�q��OsK
U��A��8೦C�je�d ԛ�b�����6��K���S90AbaHV�XK�!�A��<�*�`%��&�t���Ě4���|�w��
��i�A?�Ĭp��O��m�=�U�F-f�(i��A!0)�1�OYVIh�U�%b��6bH�]�D�&�� dD3BFߟõ������$���b��
WE�a)��H�y�t��'�R�
͋gG�œ��EŖd@�ѳ��{�����Tn�t��1\�la*v�Ez�XE���J�OIP���<�w�ԝnm�H��$><
xqG%Ko��	D?�a@[0:y:3��55N$tQ��������7�PC��,���R�5V�戋���"8�x����4�H}��'��(( ʂM��@"���n!� ��cMtB9p�Y 5�i�&"H�4���U�N��(b#��o ��p�V�@2k�L�AB&��{���pI<�䍑���I1mp�����!n��wN�L�����L�����2(| ig���=f�{�Ε-mMI ��G�u^�P����y�K�H�h�r�'�8)�@�0�˜�~b׺<1�e���!^�� ㅛ�4"#[���K�%`@(�Oڻ2��z�"B7q��R�`G$���k�,P*/�y���A*��"���#M�^L�W�0x�n�zT
�(���%{��8��N��B-��2�B"I�@l�,�z�~�:Ĳik����BX�'^b�Z���n(�˓OL���O � �fH9*��(�f�ר&���!�ɾ[��@j�1j�h�Bb/	�A����eπ�����'��b?�iGoXjB\C����"y:��<�v��-��`7"D��*��R'��	Ⱦz��͓6 Y�@]���I�9����'�]�k ��D˛��4���D��Q�:a�d><�ʳh1����d��@��]s�xr���H�F08�I��A�����V'����30�Z�S�ϋ�}x�,HU����p=q�'�,
���܏}lDA@�ę4~�Ĳ�'�x�S�  f-��S0xN�PG�^ sѶihd9s���bߌɘ��B2Y^�@�w�?�OL�k����Im.KA��*Ÿ���>	HU���0Ь�/Լ8�D�=DA��F��]o:�Ӿ��A��PZ�u��EC<���?AbgѲ|~J}��֖}��']'�t�Ї��(��)�P���l�
e�%�L�
�Mn���� ���ēo���kw�-}�yb3�/��9�'����H�	\�ou�S��ӿo ��񀃀#����4��?{x��&@��;0R@�]ܦ���	���Ї]�e8�`[d�V>"�L%���䀭}F:����堣-q�� �R#�#e��Yr!��~12"O����{�$�ŪÖ%��Eڷ�'�Q���pF�8xH������UUrMu*,D�h������H�)PZV1 V&D��Pu��'�Z(���_	K=�H��%D���R�\�'ln�E�3/B0
��%D��Yp	t)rM:$Lz����ƒ�I��'s�՚�T&8���C� #r��I!�r��M�QԎ�h0M�pR���QG|	���p�z�53��|bq���"�$)Fy�mҢ�r�nZ�jg6���'��<�(�j!e�bf�S���*,|���ӭ"�IV��~��6E�B�	� b&�J��yB��<a��uC7]�H�����^
�yR��|�=[a'�6��� ���y�k��]������J���0 �E9�yB	��}"u"͆ָ!��y��>A�$��"Ĵ�����
��yrO�&*d��pG�#�z���T��y2�G�t4��A���}M@l�����y��ԽN�5���rn�l�k�=�yRQ�
�eI��?dr��ǯ�y"
RW�m �'�Qȵ5	L��yr��� yv|*1�ٽ|�.-��I܆�y�+DAވmY�
9}~T��4bS��yR L�DQ��ӷ'�Y����y�I�l�4lagcɲjH��oP��yb��1'ߒ�	&(�R&@QP�y�Ȉ6p:u���~���'L��y��-%���X�#�O��J�ݒ�yZj�t��+Y�֭����q�"O h�A��� �@�J�%�H�"Ob��#hN����ɗ�ά�'"O��K��/gu�uIcE�.�
D*�"OB0b�㝁Ӣ@��\�z����@"O��PAEJ6v��ԓu��_�Z��f"O���Q��9y?p@�%�TP���x�"O� �L�!A� ,6@&��z���y�"OZ��@̆qx4Y���F�u��e� "O<3��!�0�r��5>8�h�"O���f�C$��ǅMp��P�a"O��ɡ�ҿ(J~`ɑߗ8��bv"O������3:�H��M y ��d"O
,cA�M>�ڴ���
0t��7"O|�B�DN5A�İ�s��2:XR#"O�\�b��1G
\��
��f8��"O����.d�5��+T�S�
�ِ"O��Їf�:u���3	��>|��"O\P��b�k=,9�D�
�h��RC"OFA��--U�l�H��?P��k�"OFh��G<6��1藍�p4 �"O~� DFժHb���A�JI
P"O`���E���J1�C�A9���"O���9	>r0��iA=>��H�"O�� �h�ur���if��	U"OL�%��"V�T,��H�'X{�"Of��ց���I�K�CM"��N�old��[�0�N��Ye����QCIS
�I��")�<����;<O�Y��C�(�8����7��h�(:�t�@*^e]��I��\=`�����i'�O0�s��ɧ49�`�%OHGZa�a�x^����TC�}��9餦�n����0�k����_T�qr��-#i��A�߀�y�iz��'M��	��}�B���9j�1�D�G�y�p��Pj�6.��Ɉ���L��O��ո���{��U�E*|���EԬ'[�` C�p��x�I�-�$���:��GO^�0��ϙ� �5���{��5�q��Q�������]�4љ�O?�),Dh(�*·+V�bҁB�Dެ�'��r�� Eݪ܃ҲidV�� e��QF.tH�h��{VR���F\�9F.E�RE� Q��=Pj�`�����%(Q@���I
���F]w� ���U+6H��$��(k��hg��.�|!E��L��"f܎r�6��H�V/<�)/P\dJƄ����
��+��Rܓ�h���EJ����
�"��
�`�n�9r�5�!
�/w.4 �Pn�4+��;��!���2��À�d�"�8v���j�G[�����=�H�P�5J�y��O)Z*��C��t�v��ge��>.���`�O�,{D���h��<.U6��W^�1�
��0�Q�c����D�uq����@:"q+VK�Z@�y'gK�,��*��=�f��ƥ�-zX��BO2?y��S�8奟&�R-#��s��
� V�(5%^$�J�D�H!2M���o��b8h�eĦOi� zs����)�ÇVHp���ɢ6F�d)�Sv�ڔ[�\-효���/7N9�L�6���ʀnɈ�R�bS�Tu�Ҍc+ݯႀ��NE�jk�w\���q�ƺQ8vP���JDE[,�d�;�#�� p�E�c�g?��Wp��9$�M��@`����p�����F����E�M!�P7���w��)Q��̈�Jl��B��s��8B���Z�v=�DM���P�"(��B�݉Ŋ�N� ����M,���'�����.W�A҈6:�\�R�;AB$4f�E�"�B���jC�^(��䃑c�P0�U��. �1�9EJ41V�!%�F���� V6�SԦX�{+�Z��ĞU�t���6��D�	?�b��EP�i&��E/�@������W�:Y��F��3[��� �h�p����\i�j�I�4²��V�!K(ra�5�_#g��S���?�����Zc�a�q�ſ�ՠV���V���F��X�{p`�jF��b��TYi�Q��J�< 
��ض*��N�$�Va��"�\j�E���Gy�\�2���Y(��ӵ�i2�쐣O�?e��b�<���QMƹ(��݈J����A�Ƿ ����3ʅ
WP̭�4Jޝlb@{�J��<�J�@ݴ�H���L�o@���
VQ΍��A���0a��g.�i ċ��*X
x�a��
9iƒx£�+,(2R��3�~=� u �H�K)U�s
�S̚u#��O������bї=��A5l����eݽȡb��8��.�3g�����J�=!p�'��Fh&��i!O����\�A�A��A���D�`g��#��>�����=qV� a��/
�z8+dIȔPt�r#���
t�����3A��\!5gϩ2�J�0� ��t,Di�?���J����h�,UU��@��Hc�-�D���^�q�,&Z0p��ڣH���@�̕Q��O�?O�
��5j
��.�ǇY*RO�У�(Q\��̋��!x��
��?N����j��ē~��g��;;k�@!�oĀ-Whi{B�[y\���C�@��%�5!ʢ�m�+s}¸�"H�� T�ܮ�c���ۀ*܅��t��IA7`j& O�-�E@�/�6o�l+����m�<-�ƌ�&$
���E�#"������	W�|X1��s(`��Pb\���X@�K���	*�*�W�~L��%ÈM��[1��N��C�ށD�Ac׌��u��x�T<4?�Ѹ�OX9��+}ed��х��k�}Yen��������OV�����Շ2�F�J�n��_
,�Y��8Z<DI0s�D.d���@�>!�pXgˇ+o���5lܔD�P�[w��ڡ
Ce��9:@!B�OM����D�'T�؈�,h�t�
~F�@:E�O�����%S���'R)rx�(7Α.�pD��%L�*uxIKG��&"i����4�5CX���7ɉ�f����a�����yW蛹42�����W	�e���M3L���3��J``�E��HO�(�t���0<��4&V�P�}�;4�4�V�M�v�]��)�bI	F���i�p��y@�ڱ���>&R��ˋ2'�lTC�:�`���Fs\����T�h�B�*���?X�v�G��h�BI�f˅�n��(�vD��	U7m�F�jq`G�^�V0�����!VR�r��:��h�����QD�?u|P!��A�ds>8���I �3wglҠxV�Áp�<�MH�G��q�u�_&hE�$7*aӬ�Ԉ�>j��ܣ�MI��T��[�I����&k��Oׄ�A�?2:����+8% ��a�/:2����
-?-(��k
�}+Ȃ1>����.>-)��o�p ̅1>�����C�����"�9�,�ݢۍ���L�����.�2�&�ש׆���J�����/�2�&�ש׆���I�6ߠ{�qBP��	�7.�2ܢx�tAR���8#	�5ܢ
v�xL^���?'�;����r��<Q�ŸS��o����z��8R�ƻQ��o����z��;W�þT��m����)��o���=��X+�`�$��j���=��[/�e�!��b���=��W '�m�)��Ml�1��]n,F��m���BLl�1��]n,G��n���@Oo�2��^m.D��i���HFe�5t�O��k�����Ej[�>4s�E��c�����HgS�7:x�N��m�����OaV�3?~*K�$&��IF��p�<(��
(I� #��LC��r�<)��"B�/*��BJ��x�9,��/L�.�����7a9������������4c:������������<k2����������zp3@9��O�J� �T~�{��zq5D2��G�@�+�[w�}��zp2@?��@�@�-�Zw�p��rx9K�쩱�l7�&T���R��&��魲�h2�/^���U��$��魲�h3�+[���R��,�������`ah�����F�e!p�������cel�����@�c$t�������klh�����N�`'w������׉}{���Ȥ$���\t7�ь~z���ȥ&���Zs	0�؆tp���̦%���Ys<�܁uw�5��5����ʂ��x�"CΦ2��5����΄��r�*I˧3��9���˃��p�/Ní8��S$p+�!����x�3����[,x"�*����~�2����[-z �*����q�7���V#x!W�Z0p|�p��x��΄{X�_6vy�x��u��͆z[�W<zt�u��}���͆zZ�R�y��R����C�{M�M�.��t��P����D�{L�O�(��p��S����C�{M�M�/��q���3���1���hiαa<`�ô�1���;���ebĹf9c�ô�1��	�3���iiγj4l�Ͼ�6�^�z�x�/y���>DQ�6��_�x�|�"u���8DP�6��^�z�|�'s���6NS�5��U�I����I8H�룢�
A_x�W�O����I8H�覥� JRu�\�D����C0O�衢�	DXp�\�B����c|`�e�UZ��\�&:���l}`�f�U[��[�-4���mpn�o�QY��[�/0���dz��'|��3�[D8B� ��,p��;�\D?K�+��,v��6�\C=K�/��.�{�$����d��MO���$�w�+����`��MO���&�s�,����d��MO���$�v���fLר�"��pc�03��
��nFҪ�!��rm�21ǡ	��jC٧�-��}l�65å
��k����x[5KV��% ����{_0LQ ��'!����~Y8FZ��/)����i8-2g��A�:S��u10Sb=)1g��F�1_��x<<Xk:-2e��G�2[��~==^o?.l"{W�l�����H��:GF��n#{W�l�����O��1JK��f$|P�i�����H��8DB��f*q]��������byh)�ċ�ؗ������`xh(�ƈ�ږ������`xh(�ƈ�۔���ؤ�,�g����K-�h{��ը�$�b�zę�H.�oq��ݢ�%�l�t˖�C'�ir��ڧ�����Nt����� xKpOl����Ku����� xKpOl����Jw����� xKpOl�����}Y#�S�&�y�N+Q�����	sQ/�Q�.�w�A'Zʘ���
rW,�]�$�|�H)S��������a�7mMi�'��/�1���a�7mMi�'��/�1���`�1eDc�+��'�4���G)�~���ő-���$��J!�}���ʓ)���.�E)�~���͛!���)��F)SN&z��M���Q����%��SN&z��M���U�����/��[F.}��N���S����� ��YE+w��^ƺ�ڽ�
+8'�U/����Vɲ�߾�/= �\%����SͰ�߾�/= �\%����S!��8�r�8~���A&�*��2�u�=y���H,�$��4��4t���K-�'��fO�����X��6��
mE� ����X��6��
mG�����X��6��j,ܒ��3+��4�X�g|}'Қ��5,��8�U�j{% Ԙ��4	,��9�X�az~'��dD�s�ϴ]�e�5�\��dD�r�ͷ^�f�7�\��dF�w�ŽR�i	�:���V��l	ۜ"t��͚i����-�X�Nۜ"t��˘g����,�X�Aߘ&w��Οo����"�W�Cٞ%���U7|�s������7�O7���U7|�s������:�B:���_>v�y������6�K0���_�\��m!�JL0��D5A)���_��n'�I	M2��C=K#���S��l"�M
O3��C=K"���U��
z�op���Ћ���;]�;�q�b}���ۇ�
��;P�0�y�iw���،���?T�0�|�f�ֆ�u�l}�f�s�%/O��ގ�x�ls�`�w�'/O��݊��d{�g�s�%/O��ߎܔ{�]�Fb�����F|9�
�p�T�Om�̿��Nt0��q�S�Ka�����L	s1��s���3�P$�-��/Ǚ��6�Y.�'
��*Û��5�^&�/�� ɒ��>����T�ձ�b��7����W�ټ�o��1����Q�ұ�n��9�
�ď�� ]P�V���������� ]R�RŅ����Ʉ�t�VX�SŅ�����Ȳ�[^��I"�ͷUu�G��ʹ�]Z��N$�εVqx�E�����SU��F#�̵Vqz�@��˱�^8+6����-SKF�g%m�?��=-1����'XGM�n,i�<��0#1����.WMA�o,g�<��:(2u�X�}TZ=a�9�i��� �s�Z�r
ZW1m�1�l ��� �p�]�xWX<a�9�i��� �p�]��A}h���{"N}F��{��
Oqe���q/CF§t��Gzo���p(FvOȭ~���Z��w�;}t
q�8-�tiF�Z��t�<u|�3'�sjD�Z��t�<u~~�1$�plC�R��Vr�@��w�/�\#ն[D��-�Zx�B��z�'�T*ѱZ@��$�Qt�H��|�$�T(ֵPH��(�[}�=�|��2���wA__1��8�}��2���wA__1�� ;�x��5���pIUT<��	
?�~!��t'Q=:`�@���+e�|�$��~,\07k�G���)f�{�.��s!W:?l�E���+e�|�$��~GW�4j�`fZ�D;����9��GW�4k�cb_�A>Ń��1��HZ�>b�ee_�L1̊��5��BT�4�0x��ZB�r��4���/�wݪ5��VO���3���/�wߩ0x��ZB�r��4���/�wߩ0x��Pn)S�p1lSѥ���;G��Ze$^�z9jTס���5O��Zf	,P�p1mQҦ���8B��PnP�3+2a��'.��=>_T��P�3	(7f��,#��66XQ��P�3	(7f��,#��66XQ��Q�1��v�@dB���B�i�T$K�����BfO��K�o�W!M����s�HnI��I�j�_(G����z�f�ׯJunU�EI�] ��c�֯JunU�EI�] ��c�֯JuoW�BA�W
��f�Կ�n���Z�i�#��(4Wu��i���P�a�&��*0Rr��c���X�e�'��)4Wu��i��bзR�
��5b����֟U�bзR�
��5b����ї]�jױV�	��2j����љQ�b� @�z�OP�f��3B��_�@��U͔+�
�a!oG�?%<���K�\�������t`J n���*e�*^O��s��(N ���j�Sń�ҕ�<����d�����ߙZR\���-D&d����k�`D�!	dNā|wRDz����^mV����L���ifOvB�����7o�RL�$	��d��D�A�8[�,i�;�4YRf��==Yl�Q���H��E%s&v*���(�t\9�#�6��� w�'V�ᐖm�&/̕�5�� Gȹ��䊖c�Թز�A�y:B�\�ZN�`!F��)�
H���B�%BĹ�Ť
�b�1����")�"6�D��@�A��u�R�	-���2iQ"4�N �C��@��q�O��%H�]��d��(���C�A,W9���LL��d�"ʋ>����1��u��U	M%DB��q���'�Nd
q��L@������X�O��y��$��2��X��
��ї�S�(N��H���];�]���1\O̕�V�#|x������rG�4 ܘo�\�	�-X��{2hѤ���h�2x�D�RǝD�61g&[�}�h8��O�?��arn#P�����%-@�5�q ͮI{�9#!�٫�d�Q�3z4���$�^�V����kA$o.��#�Ht�)a�k�'U
����K�ZxR�0��VtD}B��9J��L�EG�K̈�\?���(��R״�H!셋-U��+��Ez�Xh�[��^��E�:v�Jb>c�� c.�k0�0`��~I)��P��Ɇ� z�FK�[}z�E��c�8?�8��!�0�ڷ(CZ-�C��"�B@��S�����ɦ��ȾM��8c����wǄL�����t͍1�e����Ԩ�$}H�Q�f���C�Ds�*d*��8(�r���/�7I�^q�r�'��Ȓ�Y�_6�� A�Z���e�}�쒵�߯�I��@��[0ɘ �H,]<��Z��[��.��iG�'0V�:cC�0|�t�#�ɺ�zd2�T/F:$;��	g�č̎\��hZ)^�O��݉A �<8��Ā��'�BꝜ��ۋ��y�̋FѼ�A�h�G��I���ٺ�~�%+G\N�?@�܍Q��S2.j�'g
k�B��1�L�q�L�@M�t{҈��.U�΀��"#E��	������U�Z�H��4��_?Q�L/�BeuԟFm##D� `�h��v���yҨ]�rO���7�1S'�1'���ϰ?���Q:n��a�kH���YPɒ��\��Wʌ�E����A�ݜ�$�(�.Ży��I��O���4	�8YJW�V9f�*�{W�	�;�,H�4� X�=�O�zyh�Z���:����Kbj!
׆d���'C*E�%�3�$и.*T��b�<�4u�dM����dE�x9�e�����)���Q�F�\�;fn`0�ޣq*J�9�A�%h'�M�s�'��B��J�#^X:���;w��c��ݻt󂄥�\\*��w��0�b�@LH�	�)	�9�6@��W�J͹�Љ~k�1&AV�i�	��R'd�����+q(�K��<|�fy�ȓ3o��ڦ-D-q�d��eV��لȓ6�� ��<k���C��%��q�ȓYgXa!��Y0)��Eb�ΦWn̆�v��"'A ��}"�%�?1��d�ȓ~�a)d��'��%��˺W�>܇ȓ�P]�h�K��QKC�_p�9�ȓw��
pPR��(]�--���8D��a�&�9�p4h5��-�9!�<D�@��L&;�3�3A2�����:D��+e�h%���L֡
Ŧ����_!�y2��H���� 3&��e��yb*FQ� �&Fۼ[�x�QD�#�yr,%Q�4('"@!K/���kƆ�y�͝7���r.^:$6���"Ƌ�y�2�>�Ç�>ӆ��fI��y2��0q(R���yl^��R�y���9R�ҐeR�-��XR�`æ�yҁ�mx��Z�B: �����B7�y��$��UqU�۠аa3�Z��y2䉘3�����ց�0��o)�y�GA>*$��3�ՙG{X�[�ψ��y�fY+n��A�.h�t��e�7�y�fX�؁���b��b �ֿ�y"JI�x>PP��Y�NTg�A��y�-
��f�r�@��&��VY��y����{��С�G���Ś	�y��ܰY]�x�R���r�%���V�yR&֡%��9����Śpŀ5�y�R(.#�!1���w�ZA�F8�y
� �h�"�v��c�L�n�ZT"O�����	�����(�'Ld�UZ2���Kk�i"���D�h��L�1O"���._��64��UJ��;��+���4f�9�jI�vF���/IN�xb�;R<�X4-e����ܴO���8cgʇ��a�6��M���Q3@�
����?e���h�1L>�O_ZXiP�"����H��"c5I��U����=b��O	��r��BГ���KܒU�L<�7O�`��!�J>�~�w��^�% ��ӄ\1vHZ�U}��F�$����i��)ҧ�fA!G�^�G�,t1���B��l��(�Ѓ�H�Ŧ����O�YQF�����4�T A�UJ��Ei�o��"}R9ONH;PH �I�O�x��U@����,C�E6ܻ��ȷh�^1�O�h�)�'{�4手sV��sEH~<���B�A�O>�Fz����F$(w�9���x(��S�?�t�'��"=E�D��.&x�M^R.���ś��?i��)�'^�]jգ�t"��z�Kd�T��"�t9j��{#fx1
�/�<�����_�����B��� M��K�E����LH��'�F-�c��p�ɧ�O8�\�ס3g<���&�L�z�'��1��i�8�O�>�b3�T	&�����͎6YI���%�Q�6�J�h�4�qOQ?�B�-��pl Y3�кKq��P��M���0ҧ�~2�V�gz��R5/��Gϊ�;���<<�hc���S>Ż���	!e���уēoj�`A ,񄧟dI�y��4#��� ��$���K�����<�M���O�Odu!�%B]J�A�*C��S�1?L���e$?9�D�����e?�&�;U	�>	Wo�<ig��"}Z���#lM�x���d8��0#m�B?a��U����I%~NA�1��Ez��f��6$!��#m��
� �=tc�����'!�$�(-��%X���Sڕ ĩ�"I\!�$G��v��҈��L@�=`b(Z`W!��0W�ɴ/.tA��m\�Q>!���~!�]���84�8ҎI2!򄁲P^P(5�;Y҉ڔ�,8�!�d
x����hٟ5 rQ6.��0�!��4~P�e&��V�ش ���7~�!�dG	;�`Ն� ��h0W��2"�!�d\�b�P�CFf�8n�`ի]�q!�D��xq9�O�bE��8fk�hB!�$	�_UM�����G'�$�bJ��`3!���>A5���DU4dxzTrr�PF/���(��e#��/1K���� �ybO�AGDesd���(S"'8�yrf��wƀ��A._#( ��m�(�y�����a1�2,q�؉S#��y��3$	r�ǁw[��ВK
��y�A�*��aZ�K�q
d��7O��y"���cGd��$IG3��љV�G��yR� zϘ�����('�|�BADˉ�yU�"�(�Q@ Pj�B'����y�/]C��dے���H�I�i �yb�������20�P�1d����y���c�.E�V�.s���S&�2�y���/�Vh�6��1���ʈ��y��څ=��q�@�\��+g���y��*g��%HqǟT#��X����y"N,�p-�ԅ���X�{% S��yBIU!�z��祔2e7���H?�y�'S�EH	���	X@,��E��y2.�!3=f�wM��U�(蚣��5�yr�ǭ������cM��a]�yB�F�+Q��9��M�U�)�ϗ�y��<Y��!��Y�Q%���"��y�!��}����U%�;;�0��ؐ�y"�Ķ8}�+�B�+�!�V�$�y
� <lX�鞕q�&b��`�"O��f�72����5r�`���"O4����0�Z\���^1H�8�V"O��wڄ8��"'�$Q��k�"O��
 	�F�����v� I��"Oܹ��	��&�ەE(���P�"O��"��%�8qw�Z���ԂU"O��kt-gE����H��JFKp�<�6"�.o�f�ʳ�$�j��֮UD�<�E��'6� C7�T< �<Ȃ��G�<i��+��0�搱N*��PV)�h�<9p���.V�
�d0)�4!��C�c�<	p�Y�?4��KW劗x(��u��a�<��i��C��x:n�6�r�{�BMT�<�U/ń&�&@�#��.:)F��N�<��[J(L�e�ֆh�^���B�<Y �9}?l��ĀY�G�9�F�H}�<��
�*�m���ݩ%�R�[�T|�<�4	.,e�8P�L��OA΁�G�L�<i�c��yfM�mQ$�YU*�K�<QQ���ĤieF�/N[Դ�C!�c�<���5*��:�g�&0���`�a�<a�g�Y0dȵ`���]�ǈ\�<1�ph��a�D��-�y�\T�<���JAB�*e2�h�2bO�<)&�R�_�`uv���/f��Wb�F�<��k�`�a�ɲ/�0;��|�<a/��v�^}A��,it��RCk�n�<	Q,�B"��#(�b�(�;K�k�<�b�W"���q��ݰ*HęS��Qo�<q,̔B���Ñ*�~��giYo�<)�nR>��,p�Z���8��k�<q3ɍ�L�t9���X|�:�"��He�<���;��!��ib�@L���`�<QQhE=;��l��aA�P9�EjB,D[�<�Ԅ^�h+�rK��n z���EZ�<qg�I$"�k���	;�d��M�<��cʀ#��4B�"ub�9A*�G�<A1���#V89�@��3T0���a�E�<A���$?���$0ua|�ǯ�B�<YWd����B-9���ᢟ|�<a1`�-4���i��F� 0��m�x�<�#��q���;b, F5���Eq�<�@�L�:M�U`��uw<U	&K�j�<�s��(l$h�#�M� ��G�q�<�ŃJ6���-U<x�� gN&Y�H����d�ϖ,W~����R�J� ��CR�������=��÷`Y^��D�ȓiϤ�����+�:�" FG1A���ȓ2�$)rN�	
_�!�gM�"�J!�ȓ:�*Z�A q�~!���"Y�|@��u8�U[d������W�F��M2���,�8`P��(��l��^� �t)��Kx6h(RܾTrE��=B�"c]�2�l��&���P�8D�����S7|)R +g���)(9�N<D�|A$�h���Y�
OJ���u�;D�D�0��	*�D-�x�tB�a:D�L�Hb��L�C��o[=��d9D�,3���0Np�/�'Q�$0p�7D�tQ���*���cզZ�*��ڢ�3D�<�� �T����c�ԱA�U7D��҄a��^��6Q~ܽ�V�5D�����u�~��$�
i�]a$5D�� PL$�ʨd?rѡc 
�@!d"O�Hs6J݂��7kO�وS"OD�P�LG�7m��qG�_
s]��"O����!Ө�2�b ��Z���"O�ÃB�ey��m��(=�2�"Oj�{����H8��=Z�5�W"O�PҮ$���:�����	�"O&9cb��@����%��2�Hm "O ���e� ���Aրyl��"O��r���p\�ux����t��ً�"O���O��B�N:�@�?*4�"O��P��9G϶���!�?�Tt �"O�*�%D�^�rt��aĤ/�z� "O���2���`�����ޕ�H��1"O�`�OS�zո�h"G6]���Z"O|�jq.�!�9p�\�*��P�f"O���BL�8Wh�9�@��#�J-�6"O��+�;#)$HϜ#/��!*"O��r�E[�2]���dQ'��l�%"O����N
�:j8y2'�1wxܲQ"Oތ(Q��w�x��A�_e���"O@$��޸Wk4	bB!C�1K�8�"Opax%��qL��
��#5.4�;w"O"����ɭW^��V���:)�e��"O��؃���"}�U��둹F����"O�аV����Lq�#B�j|B�"O|lx#��\�D�A�� �q�a"O���%�mX�+q��\b���u"ON�JAJ�=�^��S
P/�.��"O2`)�Ix����ƈoV�Ce"O�a׭�|rh1T�1;`tY�G"OZ�s�	-@Ϭ0Є�(T]|HrG"O�r�#�CO��#��4����"O=s��D&_���҃�0`���%"O���C�
)�P��6CӷT���"O��:�#	�N�x��aI:�Y{�"O>�SB(R�xH�cP$Z+@M��"O�ap�<nK��(���/%<���"O*��E��p[J��F��g�G"Oz�'g�*��X�m��U��0"O�IHE�ϼJ*:��2��<9d�"OD4�SW;4+>eS$�<a�r�U"O�}+�/NISv�JVJW�[傀�v"Or�T�&r�d�!�.�6z	R"O,�+��89Τ�b,ǎ�J�"OB�q�I\gM���U��&I�xq�6"O�h�6V��P���ߥz��!�%"O�4�ࠜ1�΅�T�ۛO���"O`<A0C �3_�̸g��
+M���"Of��f,��M0�y*"&E�9�"Ox���J�@v8qS'�Ķo'HŒ�"O���ԭ���z��^�W&�m"O�1s�(�5Y��Y���]��B�"O�`$�~�����㛝A�-!Q"O +��hW��;u����´x�"O�1B�-ȳ4�,$�`畭>�
W"Ol����^b�h� J$*X4(�"O��{���R���B��-G�a�"Ox�a���]�h���J[-�%��"OX�3R��n�c��]�>B�Z0"Ox���{#�$[�D�?,V9[4"Oh����P5D��'̞q�iD"O6th�I�t~H@fӮ2��q"OX��B �&�̑��+��hÅ"O� ��I��MtH�LX62��Ɉ4"O�q �dUR�8� p΅��r|�0"O!����I��h��~r:�c"O~`ks�(Nx|�GI�*	����"O���� ݨ5�-��f[�b�ą��"O�j�,{ݼ�cp�Ͼ{F��*�"Of�2v�S�?{>��gO�i)�QY5"O�aА.H,u��je�C�^-���U"O�<����A���~1�;2"O��2�mA�KF�ɲ3� ���"O�`��Â�t?� f��w�`���"O�8��S<�`!p�N��|��"OD%��O z�^�Af��Q��,;P"O����- =\t|����:c&h�"O�ea��	g ���$V�	��A	�"O�RU��?��AQd�/���a�"O��b$
,��HaY1C����"OP�Q��D�����O�K��""OP�#����L� oV>o0��"O½��&�Ve��Z�Ƌa�T P�"O ygB�!���D0��d"OR��(ѷ�|�"��ƌˊ��"Ol0�j�,*>�{!�h�Z�re"O�
���gr�s ,Cb� �g"O4��Z:X �*g�C$rf�X@"OJً7���P��IE#%n�ag"O8�
�cN3 5���	�u����"O�]���Đt�`��n�&�$|@�"On=pA%�<yY��;PM-|�T]�f"O���右8ێX�Vfߎe�ڜ3�"O����F�Wĸ��ӧ#>�ũ""O��(�   ��   �  �  $#  �-  r7  SB  ]N  �Y  fe  Ap  �{  4�  ޓ  &�  ��  �  ��  �  O�  ��  ��  -�  ��  ��  �  S�  ��  �  Y � � #$ g* �0 �6 c= D �J \Q PX �^ �g �w �� � � >� �� � 5� �� ��  `� u�	����Zv)B�'lh\�0"Ez+��D��g�2T����	#ĴYT�?YV����y�抋<+,e�A��[�R�(UN��[�
IQ���.%8*�������"5�ֶSz�N�h�4��T<h���	&��<8A�K�V�|��eÑq<�B��4&F�r�GE���6cƦk��p��,����'r�v�֪d|Fa�$�H%`�����W�p,b%hJ.1I`�$�6Ε���)}L�n�5?���	�,�	�� ��}�2,� Ŵ�FQЕ@��:�%+ ��0���;ش/����'=���O�Pr��O~R�'��b��9��jv��2J�ڵ�P�'���'Pr�'�r�'b�	�Yw�8eK�n��@礈��/ȓE,�0H5��E=��!��z��8͓Va�I�Nu��Gy�IQ�Ol�O P�����̐<��1�X��Γ�(O�]ctn�6�`�'��=#V�߈	..����]�t!hQ����?���?����?y��?�/����4;lbp�LI�%+���MZ�:9��æ)��4mz��iCGa�`����٦i��/��pDNX���%�N�{��G��,�ge�����־�*-[�f�On�ʕ%��l&l����7M�?�Vǧ��)!ꚳu��1
#gȁ+xp}
���1��8k���Ovl�M#�'��T�O��Μ�"k��G/�+:������V,H^�7mY�*����F�l}j�*$ɚ9G���A��Mv>AmZ+�M�A�i��ڇ*٦x���ك"�B+�t�Є@6z�����:P 7m�֦U)�4����g$\�>ڴ�@�~��s%�{��<�1G=WȮ��g nVL�xŪ�3Hs�ѳ��i��6��զ�a� 9��YBjL�8���M�=�fD 3/\<�I�!-т�hشX`�"��֢L	(Qa�e3;������'��Y"�z=x9�E,g#�@/�����O0�d�OĭlI�$h�5��X��ܧYv�8r����?�)O|���O����PXΰB��S	��l��sf��ˍ�*P��*��;k
�k��q�Ty�b�<�� �SЦ���M��b^Ѐ`bb�4[���a�1�I��	��0���(}�VhJ"D915��A`B&O.��$�Od��-���O
�$�<Q��$��C	̗T$���#&H�1��?���]31����I>i��<ͧ,��ȟ�N��0��䄿&[h�u�
 �?�,O,�i1(�����	g�'�yG"��}3����Z6#�
��"����?���B�|�
1J]�;�0M���i�E�iS�rS`Dxn�.5aR c�I=9"�{" ����M�9U�:��Ɓ����'�>h�J�\�L��*#���'�x��� E��3ҧ���+�L�D`��s(J�����?1��?�,O�c>eA�eQ7���C%��1W�Dh[0�=ړ�?d�i=�7��OPn��|Z��Q�DZ@����	{6�Q�'�M�����D��Ix���O����O&�h��CD�'���!�_�@Y�:h �(�vS�; T�`.b���?��Bƀ�szl��)��`p��# I��\�4��-�����*d�b>B��Evy"�؆�±�E���a�f�+a�v+�<�C�͟��M�L>i�Ѱ(В�s���T�6�.I��hO���Y�4� 9"ꋑ"���C��
r�"�']�6m�ҦM$���?1�'�@�1��.0nb�S ͆ 4�)m^W�x��?y����d�|r�O�pl�P-��9분WU��c 	a��5�c	�*\'�v!�p<��)���1�'J� Ұ-3��Y�qy!k�(P�uz �#�V+C?z�{TA\�1�ȣ<)�.���@�L�r�Q���;3�l��%�M"�	Vyҟ���*^�z�h���L�:H�e��O���,�I3Re��!������C�k�1���$�ئe̓�M��i��31v%�޴�?	�d�>a����B�^��¨g��t���?A5�˛�?���?���	m��� �n��a�����<>>�2!�{��&+�D��I&���0<��
��k*8�����Q<�f��zG܍���3x�8�tkėII���4���0�FxR���?���L��&�'J�z�o�f�<4b�*R�t�剡k�4�?���Q�<i��I�Zp*���~J,M�P�v�	%�M���4��]lZ���(�S)Y*�f�@�%]yz�.!e"�$�Ҧ���F��M��͌���$�|�'�X�j���-_�uP�!� ~%S��?Q� ��7j�Y�F[)��i*F��1�>5bé��2�N-�2L�4k_�!���/8���%OZ�^��H /�0Sp��^����E�]�ҥ,�c��۷����)� V\~�/�;�?� �i��&b>��ш�5�����`.�ڴ�,���O��O���O��k,�cթԚ���'��i�5��)�?��4�?�ױi����j�x�@�:�޴�b��3;6M�O��d�O�%�0Ś8:��d�O��d�O4�<t���WCߣ.>��`N�Q�d"L<�搹.�X��|�<Q2AJ�$���� &UV�0'-���'r(#2H���Ϙ'�¬GV�,�2dҖb!��Hf�i
�i�$�IL�矔�Iޟ����6TD,� *R7Z��Q k�o�<!��½_������H: E@����r�'V���'�剶?:J����ne�}�mNA1L��&�M{��?�����	P����rO��xʰ�9Q�28�S�H��� �6���$�D�˓MRJi@�d\�(�F Y���*�xqi�7HWbM�1LW'De���
,��p#'b�]�'�B�A�/�Ѣ�[.]����OL�?����?�����!B^((��,�(I �A�n[H��D2�*q�Z�
�#��Q��b�ȓO�n����'V�:��'��ӶNc&�9�%ΘL����&0iǞ�D�<q��?q�O)�ذ0��� U��,c�ȍ�� d1�P�T�G�,H���\D���'�Pt`Ŏ@(`JC��,l��}�`N.'B$�Q��U�&��D�T ��usb���Of�0�'B7�wy�B�<vV<�Q ���\�t�C/;����<���~Bތ���	�kZtu;$A������?1.O�=�'[[���.���� �2gd ��a
�6ǔ7M�O�|mZU�1�ڴ�?�-O���<�u�U�* ʆ	S>'����"^��?Y�d��11�^/mO�z#`�Q�� J���,�6�H͹�f��̚rIn���� R�$Z
i?n�Ԫ�W$	�po�-QD�0B>��m˹ �U�Tl�+Fdi���D~��� �?Q��i�"}J�O#@́BN2W�6�����s\y�����]*;�8 ��`܋ma� x�L�	�ў�����MӦ�ib�'�\�r�ဝn�&5s�^��ț�e�*�D�<yr�������?	���$�e^r$�4M҄t7�<��˦*�ByYw��}��Ձt�M�~�~l
�˹|��g�QU6i�q��+���A�H/#�R-`&c��,��C,���<��(�A�';�b<�o��<q�Q�,y4Ӕ�������ȩ�MóT���ԇ�O��	;&�s����� ���|�Z8�aKe��hO�'
Q.�Z%c����U���[0`����	�|��4^|�6�|�OT��U�h���:_��I����]٨���[5�����Or���O�˓���t>��Gb�-�����iݲ��+�GE�$D��xao�'<��ʢMF)ް<���q�V��@�ʨh��웡	Vhw2��GKž+�B<��̊�*�`�)U�ߨC��#@°��D��O̺�k�
݊�9�!�\��4'.��PExB�?*��=)�
]����F���I������B�=`�5�a�ں?a����Z�HU�'@^7mG��'�8�bA�u�t��k��@�m��h�|"�EkK�4I�D�O�˓�?���?QM��PlQrǞ (���0%j� ��'mחTDha3�ֶ;7�  �'�xl[���V����B��f$6��F,Ȍ��Mӡ|��:c��?Sax2���?�����$�#'I�H�m��Y����E�UM�'L��'ӔC���P����◔<Pz�X�J,��@$}ph�$�
�",k@�  �?�(O����O����Oh˧����ӟ`I�<�nXW�X��ͻ���D�	�]�8����Z��M; �$L��.���'H*V|s`�q���q�U�q�l��O�ݸ���\�����o|ʠ�a	�
86V �0��?�����>}�r �L+3�L�t-��uL�I�Wf|���O��}R�'w�|���1"ZĂ�o��h�]*	�'K���ʡyd�4Ϛ&_�(�؋���u�O�B�p���~Sd�H3a�	-IDY����?)/OjC�'�z��\1ALU �B���nTR[�D�5�>�$��A&&��|��x��N�w�ĳ�ꗔ8X&���[�[���Pt*ϡ)����pFR]�`Î���?��)X��I��
(fX�|:�Ƀ,>���0�t
�O��$0ړI_� b�"��4�,8*\M8.�C
�'���1�ϹRȂ��y��|3*O��Dz�O�2Z���	-a5ԩa�m�7����6lIvd�����ݸ08��/X�\Y��NFvQ�Cc��3�y���B^PӉ�dL�	��4�e8��aQwh�0(���8A1�1!+RN�:�"Rg�K�'9�	���1a��ڑ̀>�ʒd�+�?����hO�"<�m�f0��S�T���:�G�t�<!Gh:���!+��caz��&r�I�M������A>I�:�nZ��@�	�}�nq�,,�"�ۄdF0�R��	�X��������	�|"䋚��xA�&��iX�=l��@%g=lx-a�`A�.C��� `O�`Z�<1$'$>��X� �66a�3�	#ʠѺ2* �r<�|3C��\	.�JA
0�ޢ<Ɂ�MzK>���ОF��8ǎP�o����A
j�<apS> ��̺�8$�-��^f���hO������Iq�1;�!��K�@�N�!2�,�䇵L�n�mٟ��I}�4biRj]��U��L=�jߕaR�'P�\C��}�z�xC`ލm�U+U>��O٬X�C�>X����S<Z��ћ�O4�9@�K��2d#_�[��B���4���?�qE�0�nh����#/�P���3?�P[�`K�4vz�>��;H3��3�f�'(m��+g��7�Z���0�F��0��-"���� @�G{b�'�#=1g+�f���d�M��t���¤Z�I���>Z1je�m�����؟��I�?5�%�����&@�<I�.�h��n��M�R��^{�&,�8"BB4�-��3�I�]sذ{b%L�>{��
&C���䣁 V&8�`&.f�-q�-E�i�l��`>�sQ�	t�杕]@�dH�/P4ڞ�(r,]�38&��)?)a���I^�'\��'JX�jo�a����)a�Ti*#"O�����ԙ��h��J�P���eR����4�\�$�<Ad0�4�i�_�½����`[fP��i]3�?���?�����?ɝO�����7F4Ɂ� L�(�>0P�N�W,� B׏Xd 6͞YX�H��-� tE��e�+�Z]+��<B��5�)W����S�V�DU�̻��П����!�����*7��H��B�B}ұ8��ל�:��Ã�H:�d�O�=q���U*nH	�`O;3u~�8��9j�!���E}�U�7K�W�x|d�5��'5�7-�O�˓V���!�iC��':n q���4jg�M{T�ӉE�ř�'�2�/AIB�'��陮]��qvb݉|qA���F�#BA�~ :Ur�m�'c���W�Vi��z��V][z�P�Y&i�������= �R�*L�H��������f���@4&���gLI.�4�iMP���˟Hj�4�?!�m�?/hu�#/X�hR�I���9��D�O�㟢|Z��R�9h��b��-�v��� 	@�'ў�۴Z��|`#�HN�e!rZ�)�P�B�i��	�W��y�ش�?������ٴ�D��361�����bzx���J>x���O� b5F�]�쨂C'�ѦJ7�S�d�?�b������1c�'{ĩ�AH%?	���$0j�a�Hn�9���YP��>�[SҤ@�4᠊Œ'J�Yr�$?A�Aȟ4��4F��>��'x��C��7�2���(J�Z<"���w�	By��)س�z<2"��-����·,�
�=�'����dӶ��G��̓/�v�ԯDP�T
��hlB0�Od�d�O, q��"g6��d�ON���O�]�%�v��Rn�$7u�a�W���-{���O�!H��IB=��B�U��T �h�,g����T"B�`�K� �ms&mɍIW XW�����	|_d��"�M�Vy�*Z�u�$elZ�M��PD�j�f������F�:�߳Py
��,R�n[�ٸ��*D��SJ�q6�(%!�&_Exh��O��@Ħ�8ܴ��s)vI �'��$	�r�+B`�
�6�:�J7,^d8����	����O����OR��;�?�����Y1!��Dq���W����J5�D���*�,�e	AҨԄ�I:+X���D0e\�9��̝p�hQ�)�</�2��JZlw+�	n�ΌE{BFϋN��A��6�.�3��F $;�J�͛�w��㟠���*Q� ��0��|<��a􊉌��=�yJ�f�`y�RB� ��1R'4��X���'+��ԟ�sٴ�?��BS�@�!�V�}��ꄬc@�ȱ��?�Ǘ$�?Q���?QF%��y<M��m�5_@8ȱV�~���G,�"}3�@8E��$���a�7O�):BcΡ*�.� f�N�4�:���E���q���ՑW�<�@��O�G����
��8��P�)�b����\qN�������*O�AH�x*ha��ȔwF�i�0�|�Ie�C��h����O�XPՆ̑-����I,@���'D�S�'Cy�Et����о2�f��&�@�?/O��&&�ܦ�������	�?�;Cڟ�34��qV&`�����~�@}�pMܟ��I"V��$ڤ�.�&]pw�F1& �O��S�~�$v-A6�m��?���<����&DSҸ"��B�`�)! �!��' ��]����<f7н"WK��#��'�l�K�3@���'������'�x%�A��(�����K)K�:���'���'�B��!v�����l�{t.K-Ǹt*TlG�'��I���d�>��ɏ9�9P��ÔNc�:P&6�H0۴�?����?��D��r���?1��?�p�wd��5�_�ς鹑��j������m��ʔj�%��HJ��gܓ:z9���>b<R���޼f�V�:�e�zBlhCT�	h#��k�o�y�'RM4QR/O*<�B`L~~8넊ٿa)�dH�Cb�
�d�OD9�7��O��i�O��D�Oz��ORth�ϑ�R�k�ԳPq0
?����D��`��Kk�ԓP�@�N� �r# Ȕ���J}��/��DB�q��~�����(����3*���p6D҃#�
�8;r�'
B�'6,��͟���ڟ�V�@-Kl=�N�|���B��}q����$����,�����I�D�`�P�K�8 ��\r�;.n:���i8O����:�!��Ƹ ��m��� ;�R�'�NOv�D�O⟔:p酋o��q��덣<���@� m�	ay��~b�i�1���;��O3L� (�ɞ /� бT�`����MS�����'JN� l��<��3����ѯĵ1��hab7+WP���˟���EΟX���|�#)Ƀ92�XYb�L.6�	�<�ޝ�!�M�mT�QR�X;`d��w
b��Q$��=�6��'M�$Yb��2*�����ʚi3@�iÓ@P�A�I8����C�^���0��4R���ȓa�Ji��A��zH��Y��}��	�?qu��k��]�G����K�p�wl4��4�?I�����=u~��d�#6:��BA�ZhP̆����wzx���ȋ2����M�Bh�O[��-Fy� ���R�V�|,q0b�3.��]�jM�������v�^�s�ꕏhF��`ɹ`�*h0���*�Fm���Mx�^���Ck~�'G�?A��i��6��O�#|ڶ�zu D�˙�	���X�i�g��H$�<Dxb-:+e���s嘂BEV�ɤD<��O�hn3�M;L>y2I�0~�z�K��²D��[�%�Y�4	����?���!d嚱�?q���?�\��_6�( ��k��p�G��4�}�B,�8i���(%��6M��00j4�3�	�5�छR�
;R���5Z�h) ��"�h�1�%���������xn��|�դ<kۜQ�{�? �
'㑻��5�g���ȍ��+�D����d��"�L����`���aUn�!�dٴO�"`B���`СÕ��2~�I��HO�),��[k�0�(�������[�6���H�ÉU�Z���O�d�O$����?	���?QCF984a��1lP<�"�W(w����B��f��)3� ɸ����D@1���
7h߿M�p���fB�y���S���J���s	��u�h9D���XH7m.O�`]K0g"?E�R� ���ԭ���A�(�����O��k�ӟ��	w�	�|�CD]/��D-\�:pة�KS��D�DK�bZ�:X�:e��F��S��O�oZܟ���4��P>P�O8�MK���?�I*A�hЋ�ᅙϜE����<�?����B�����?!��AѺh��ِN��q�T�l��ͮ1|���TF�7-��Td�F-���ɱt����`-F�k��>�,�9Eatt Q�1Ѳ�q�X�,bFC&�H���'?q�.�ş0�ݴuJ�ɞ�����(D�0���l� ���O:��hO���<�x�Ū	En%��E�d�JC�����[b�8A�S��؛00t@eˣ�M���Sc�6j�/��'���'k�	�.��N?�dȴ$�!f\��uJ��w~"�'[���U#A�����Q'�Ԁm�|2-�f��͐>���6G	���=�4�.?����m(eJa�o�ԍ^"�,�i@	�2����g�J�O����r�ͭ�\��>-�(�ɀK7?1�ǉƟ��	b�O��D��p\��rK�130B�з@��>�!��A�8��|�H�����\�џ8���iC��zl����c ��0��]/xfR�'���'�h�C&n�5}���'`��'n���G*.�!�K؆;��ݲ&%Ð2 ��$�R�H�m�/l�v�iQ��|ڝϘ'�8t"� �6�xĪ!�D.�J���2e�P�@��� �r�A��6���#�����$oI��	a�w�.�2�
�����i�7Z�������;!��'`ў�QTCW2iy���A�݋on,�8��Z�<q7.L/8�B��OR�.��ą|y�5��|������}�v8b���))���K���	i��#!��$�O\��Of���O���y>I�IK�c�#�e�2
v@i��W4Xpؙ3ē("����4tayb�Í{ 41��E�C7���F��j*l��0B�+O��9�B�#*0��H�O豺�C��sYz���O��c�
�x�\i�)ŷ�*1�c�X2r�'�ў�FxBn�2�b1R��Ҭ{���X��
�y�%���ai�77%��(2���HڛF�'��	+%��u�N~*��!^ҜeI�|��5��������'���'��CB�Κ��1�ӮS�j�xe��9Ҁ�4�M�m��l@f�\ ��'X��{S�VPeJ$�7`����O0���I�_x���!ĝ�0<Q���?a����S#��5�� U�,�!��B�J�'�a| ]�o���R*�4Z% h�e�6��?���'��##'��,u,c�� ��͟��'�83�R��'���Oʤ B� ���2�����e�%�O��Dٿt���9"-�/.P	b�>Ô�?�#��ř&KV����rSx��"�f~2�Q�/�zp2DC��}
��p���s�O��rQ��f�ʹ�EB��kg�"�O��s��'�b��<�'DS�;4LJtCߕu�L��5s�<�ǣ�9�H�q�V(�dN�r�'��}Z��P�5���oG�Z-�lP�h�Jy�[�����ɟ$�	��	Zy�Iɚ ����hV87�nD�1�E�{`X,�$�l�5R�&:���P>%�g�Wo�)�*מT�8� ��ʱA����%�rI`F(�Ke�yh��@�g̓
&�B΅�J����G�*��|�IG~�����?i���hO^���6[x4��eK�! ��c3�>D���#)]z��ZDn��{���(���<q��)�*O�����60�d����~����N�Y��D�OJ�$�O��S��'v�i1�P�zrX�Q�s{���t�X�%K��P�K	3q�A9'�ք�p<��"�f�������6@��		1�IP<Ie)�+���r'��
"_���T�|d<�� f�:�0 �#TGI��B��'P��w�'�&�R��ϊ�*5I1��/1S���'�HaR���f!>
�N���K>�R���'�d�$+$���fめQǩ�?�P���
d"_���I����H<Փ��6g�p�����@R�{��P��ٶˁ^b=�F�U�P���
x�ls����|����#Kt`�ը�,��`�T�5T���S�FBR�'�����s�I�w �,
�
<N$�O���$ك=Bp��a�c3J��f�D��B��O����R..�"��2e@�j����p�'�ɾR{�ɗ��I�|��� �t����Sl���Ѩ[�(U�����?A�K��)�fu�1��;[��ų�H^��O��=afL��d�5C�H��9�����LK�0Nx��+�^=ar�S.�t�1f/��n�*��)3`�~޶��IßF�d;O� �@�҈�8F}�a$חc�<� "O\sF'��[�]6J�wrD���"�h���HA!�$�M`�ӍC��ۃG`��y�t+�<�2�����	�r�1ڥC�p�B�#��զn2�+��g_���)T*$��{�.�3扪$��+Jj`<�p��/20�`�{�F����!`Y�#-�3�
<�F��P�oy��,����l�
��$��f�"�O��3�d&N1��yb��y\���O'�hC�	5=|R�""H��6�����
ww˓b����Ԫ1��y��K���(8e, ���ㄈ�צ��"�<\Ol�G���^��۔��*�� w��"_��ꔬ �o�|�fĖ�p<��^�(o�<�t�4u�,�K�q�x-��!��RՒ$iލJ�B��䇇 Z4����!6K���a吊-L�	f�'@�7�YV�'���Q���*HyP,�숮r*BP���1D� "�^�w��
 ����P��:��A}2X�,x�cד�MC�B�C�v��
Ln%H.K"
�4�a�BJ�'(�Dʈmm>�sp
��v��d2+� 4��<B��?O�	���)Ύ8'Dގ5�b؉ K #-����8!���,�䓖EB.�g��m�4��O�
�!�
b�QI3$�u4��8��٠>��f�O(y�r&�(S��0=<5�����|R�ک :7mҚ0�Q?{�U�D��@�E�v�L��*?�𭁙�t%��M�];�yC��:�'B�:<�&ƌ�XW��҄;����'�v@6O�A~�@���~�,|D���+y��@�	ȸS������dӐq��cf�l0G�$;�Y��o�� $�Z����<�1W"O`a�SK��c~�`��)P���Q8�����h����D7���	RNޒ3�n)��q�(i�i�<1e�R���	r|A��>9l�EYQ��P�yb��?�0=���?T�8��E�۵k'����b�u�HHT ���12�pô�����ڦJ�c@P'������OPc>c�l�c��Q�
�#�U�$ܞ��1D��u�Q��B��c+R8fŐd�E��<�r�)§Nj�P�rk�?$�J��ϐ��DH故P����,n�
�rf'j�\���¤"���'����w�B|#D�H�����Gj�;�40;��'�R ���'���'�����̈�t\�U�^h}�Oh �a��5H8X!F�E�����~[������&>	�b���Z>�٦�ÅV���M3�bY��I럼�|*g!X;
jh-�3+R�Cn$j�}y��'5ܴ#Q�Cz�ĺ�G��s�&e����bh.$�%'N�(�h�@����*ʓ��<��w��)����	��I�O�8I1畕7*���0�zm�7��O~ �œ�;,�1p�[-L�:���t��W>u�'o�H z�M]�Be�tكIç��ϓo�<�S�@�������GˢV���s�*S�t��y ��/Dwl|Χ�|���d�-��nD�	�y�Ҭ��Iޟ�������	jP$[w�1Hn`1W��*�!򤏂N4��EJ�{�~)���
0�ў������EPʩ���5`��Z�nJ,X�⤣�<��h��<q�g�'/����˿3�֡�q�E!f�xWS�r~,r�O�*H��j����Ia��V����ݪo���r��	�>����};2	���j��t.5�Ο��>�p/_8}F�rDB?;�:�Hj~�L��?���hO�牿b� ���N�:[�,x���*��B�>E��Q�Į��X"�&�oHn�D�Z�����'�I`�E^�����&Oͨ\. %�C��)Q|b ��p=��Z�N˾�Q��T?O�Bd�� �7}���`a&��a�G�
�;oh�0�I�<�r��W�^91x��>�.�ybdУQ�v��2��-,�������O�J��'��Kb@w�l�n�pd����'lў�E|B)D,9�0 �7����0���y��Ɇh0�UH���,b�V$17b����Jɦ��my�%3�y��5��S��(��,�;������=92�">)C�T?J��9�u%��H�� �4��-U�N�P��T�`I!D�M�>�h�!$̑JAkѦ������J��uW��R�*�hCh�+�������OD�!�'��1vp,��X�MU"e1�O�	��K�� ڱ�<^�J��P@I
{�u �6�Oy��ϿQ֨�UGH-N$�7��?������$�O��?�'�T�IA�Ov5Ld&�T�j҆4�'� �(�IVT́���><��U �("ҧ�13�mJ�-3��(���mR���{�N��ѥ��!��M�u���8t�J6��N�rC��/���*�
�x�I�6�����O��S��J~
� H4�"��%����eI�9���"OA��JߝX�Z����:��-K��I8�ȟZ�D�O��4J!cI4*�D�h�K�OX��r�?\O��(gɎ^�jD�d��u�.�Q��iJhI&Ls_�APF(�,��S��'� �`!
Yj����Է�������$�R��숢%����-�����TJ�Y�d����̚ ��LS5<�(�'>(1���?��Df���`�W���ՠ�PUxIR��(D�P�c�7T�C�NbQcf��Ox�Ez�O�bT��@#��D0��҂�@!������[%v؅��	/5����NۨGet|�4�ֳj�@�R�F2�{u�K�u�����M���O2�3�KU�4虖fHt ���"SD�����W��!@%≭��c��9�Ed(�	�P������w��hh��Ӟ�t���e�'�� ��/�)*^�C��ë6��	E�2D�ء�3@�l<J%ǴV�\�%�<I�i9�P�h0$��M���?a�O�z��"� ��(�8�8�d�µ�?1g�J3�?����?Y�O�2AFt������k6蒤�¬��t�A�
��8*���?^���rti>��O��)�tT��mүf����N{TmR��΁D��T�7j ��-��!;�o���	4��OԐ*ī��[@0�%M[���Y(	�'�ؐ��)�h����ԇ��&�8M>���4����'��i�G�a��<�T��z�b��-O���O�˓�?A.���
�ȉ����Vv�ѝ�>����(O�HlZ_�O	P8'�	 7B���1�T�k�r�i�'Ҋp'>m%�#f��X��U)b��8���4�M;����8�'\�8{��?y���?a�'�����L[0Y�0���R�5pQ�Ў�Os���'�T���'��dO6a����u���<��w��P�΍�?W�����:$���@ˉϟ���������u�'*��O��3O&L�e+	l�zd�D�L�8S�Y���'�RF��@�5O��F֟�^w��H�$�L� Dʒ]fL�r�/�>�V��RG���I��S��=����O�����d�G�T���C���P;ҥ�[�vE�I�u8����O(���OP��	�>�s�tE24`|�Pӭ,�b=f��:GnZ��?х��Ɵ��	�B�rm������OJ��K�@�Έ�0�ݽ,O���
�i
-Q�l����OZ���Һ���y�+���ܴ2�t�r���17:����D�*0�����(D���6Oz�4@j�(�m�#O`½��u�O��tJS�d�a��\� VN9�`J�@�6M��3�\�	(`1l���M[�'�?��'dr�1�p�l��j��ڄiX>t#�8)�i�+3�'��	��޴j���Y����C���@���:82�ʜ� ��j�^�{Ӭ]4C��U(������nZ�X�����������������(��?�f�f�A8>���1���Py�Y�4�?����?����?!���?i���?)�U�X�t�J#k��1(��ǐ}�t-`S�i���'��'+R�'�B�'���'h�a���'_2Lâ�ЮD��Lu�4�d�O����O��ı<�*�����fD�!��Տ���q��P�,#D듵?���?���$M:i���r
�l�:q"gy�	n����' �I�l%���	- �OԤD�v�җ'��R޴�?q��?�+O�ɷ|�H�8�@�'
���hN� [��X�7D��χ������*X�p��3D�h�n�;p��;���N�d�0
3D�d��O��Х�'Ժp\DP�Ճ1D��򡨗�/1<H����i�x|�dI.D�Hh��K/w`���j��PFh� ,��?���?����?��������V�>����`ʸy3���'���'���'�r�'�R�'�"�� j���֣'�����퉉3nH6-�O����O�$�O��d�O8�D�O���	� ��0���ڢ>Đ�	1�����l�̟l���$�	ܟ��I�p�Iܟ0��f��`2��S��*Y �c�d��A��4�?a��?����?����?����?��a�|o5��My��"\�FD+�i���'�B�'\�'qR�'�r�'���8�hR�(����
�Xa
��'�"�'���'�B�',Zf���'�"m�g��I�7IٻQ�l��cR+9#l6-�O���O����O����O���O���Y?HP�$�d���, �P��NӞqMo�ڟ��I՟��	�� �	�p��ݟ����dw.�`A��9�ش�s�1.j(��4�?��?	���?����?���?��,9Q������47�$m��K���M���?���?i��?q��?)��?ّ��tXl�T/X�VY�;��ߞY���'���'���'<B�'���'����5_�6�Y#�ͯW�8l�b �vϮ6��O.�D�O���O���O��Ob���&X�0�.ܳ;� ����Jo�m�i~��'�IS�O�vy�A�dZ�)�t� ����i�4H��'��'
��\>�(�Ms�w��%:!<)�]IT	��~|j�a��'��6O.�S�S�*C���Sk���b��Q�G�8y�#%L5�ѱ!�O*���+�d�AZU�8��|B�'��q��X������F�X;|j����&�d���-�G�/�[�? v��҄׾Jx���"YZH|���'L�'��ʓ�?��4�y�V�H�穛��� �Cߠw+l�Z%B�<����#R��g
SR~�O�HsNԪ$s�dݔ"���pfד2���%�J2cc�Yy2�'b�>��YǠD�˳M�@h��IT$G���C殮y��>?��i��|�O��I�
�'�Ƚh����F�p(�2O���|�2�D�{.�P�#��peDQ,L*����&%R"m�Ri"��PO�
&ͮq@e��şL�'�1���B^�;NQ��E���DP��YܴD0�!�<��'��'}�Zm-A�x���M��R@������O6�w��G��a�Ty蔋OF�BI��h�?T��� �P����4���с� ��'���'h�ث�o�tJd�%�V�S�$��'l�&W��>���L�6��1�y"k� ��))���d�j�����B��1�ଡ଼�\V���X�L� |`��TU]60�OF�Qʠ�i�� (�f���^U����f�U�x���!q�[i%���uIK�e�p%(�o�'"�B�Igi��7��x�/ď��)��	GG��p#���p��4���� l|�������qS���Ol�;��l�� fC"*��k+�>�n��ֆV�w��a�C
�O����OL�4�����+� $@�gIХnr��[��½��'�7FB��Ҧa�O��Iv�N���l�/��i��W����w�.�a��;~��d��@�)&����j@ BhC��MC0\I�c��
k����c�4^pa�ԯP~��Ը�O�0��2��{�ҥ@��H�U�<]���"5�V�[j��t�TM�>��r��+nJ����͎/I4��+�!W�H��A&�?n�X�eC�b��H��"H
-㠥Ȅ;a^��g)�/K�6TX���&G�- �-�TqSw&�-H�������\9�0{s��"����m*����M�-����#T4�=w�HR9L˃픿}��QK/|\�Vd��U}�+�i�r�'���O=�ʓ6�b�*���'/����%���D��P�I�x�ɡ]�h��Iʟ���柴��ȟ��;kz�1"�  >ִ�@�Kޜ[��Ʌw*B���ȟ��	����̟���\��S�G�t��1"$���&�-�2�ܫh�D��y����'�R&6��� ˏ^�R�K�d���'��'�H��'�P>��I�<��EI��l
TBȋd��9��W�jc�h��Cf���'x��'��J��ĝ9��;hp�AO�2}���'�m0��'�RY>���C�6Aр��8/�����e]�/r��'JU�&a@(�y��'��'�'��	BC�(݉#C�`4����6��$�'�B�'���'��'���'B�=A�̓����#��$7%Z�M۹m&¥��O����Ob���Op�$�)p����ă1�5r��C�rD@�	�Z������O>�$�O��O<��O��Bk<{��	ȇώ��(EC��!b(�C$�<��?a���?��,�)���?!��:�t8SpF�vݎI
ñ%=7`4h���?�O>a��?I7��*O�bԧO�K���!CRvA@RyƐs��'�"�'�I,LٲI�I|����y�(8kn��ȉ,j���0㏛�?�+O����OH�9��３�G�.*��0�AGY���H$œ����'�Ne�wOq�T�'�?�����+����)�[���Ґ��-J��d�O �$T�&I*��|����O�YY���2,�A�F�db[��'�ZT�#�~�v�$�O������'��Ӆ���( �T	t
��l�ƍ�I7C؅�'S�'&��y��':�!`��e��d��,F>��cl{Ӝ�d�O�����Kb\`'��矰��3Q������,T���ԫN#I���'���'|VD�y"�'\"�'��*�@�'���Z�$����"��'	b�ɥ�O���OH�$�<Y�JH��yY�A�Dݶ������?9�ke���<y��?i���$��i^�8�ɗ3���� ◃'���@�	�,��Ο$�'���'������!UP�"U�� V���e����'|"�'BU�L����-�O�>u���Bk�h���TPy��'��'@���	��N������0���Yp����H��;$rʓ�?i��?�)O���O⓿p�6�q��m���
g��\��T��ϟ��	myB�'>̚���OR��S���;68P|х�ďo��� ��?-�M�-O�9�NTg�S���λ@ʀ� i	 �\�@�U�.xy'�X�'���(��{>Q�����-MܰYP�0&�1��D�O��{%��8�i��S۟���+��$�-r���pA�o����I�h���'b����)j�g�D�,=�Z�Y)K(%a�g\+"i��}��7��O����O��Ir�i>]"�ڶD>� ����o�d�1aG�џX�IMRy��'D��Ϙ'l2�ؘ&�D��T%�Eb~AP���9��7��O��$�O0�)2F�q�i>e�	П���6	4h�4��I"5"0�	Byb�'@���=��'hb�'D�-�O��(e���0�X="��<$�r�'¶T�C�5�4����O�˓
YX1��AN�_xq���$m�-��?��Y̓�?����?�.O"�{��@� ,"KQ�0a`$!�>$0(�$�l�	��X�IDy��'��ܛ-� |�'���\�0��2I�-2����y��'��'�I�{��T��'th�P�6�Ϳ ��ys�a��EN���'���'tbZ�����P"���?e9 �@��φ �H�+'e8Y���H��Qy��'	���[>}���%�
bK��v l`uhL84��]������?1���E 7g�Đ0~*h8�Ƅ��OR��&��\C��'X�	ڟ@W��J���'a��O:2�:�
&::�s��O�*����O�� Oʵ3�1O�� �8��n��M؃o�Lf���\���G(�������I�����Hy�Θ��h c�㐾R�v��6BO���IΟDC���B��c��>}���� Rv��I�1>�.���/�O���@�O,���O��D�&��|���uW,x�aL�
y�X�3�D1|�V ���u��QghWj�S�O�2�2w�dH�,�QwR�	�k�2�'�R�'��0�Z��ݟ��I�<y��ư��s����	��[V (��c��C���i�ݟ����<Q��3'��c@�{�>�/����O`�!��<��?�����'�乣��f~Ԑ'�#6�-O  )��A(s:���O����O^���<��N�}1xݣ��2f�T���</���R/O����O~�D?��ϟk�я�݊�J� BT�*� M1:o�C��.?i���?/O��y��S3XSn����s��P4CL�p.���O����O�⟸�	7*�f���*�4aď^�_���ؗF��}�'�"�'}�I����D�~�d1O��@LԎt�ބ#���'I>53��'�����OP���,V��lQ��/�TI�H�ьu�|���埰�'2ҋ���Sß��I�?��tYw1�d�f�R=bnR A��J@���?�C�I4S���<�'�Z�z0�[��eZt��x��ї'���j6��'���'��tR����SBؠU����^{�
�o�oyB�'������ ꘧�O���d(H6�R�p�_;�vu"�b�����?����?��'��4�J�$VԢ,�C"�61qiB"�����!tql��������A�)H)+��I�ѢW�N��!@���$�	؟�	%�엧���'�>O�C�N�3Si���	Y�-G~���AN���':���e��t�'�<O�I8�L�(�`݈�����(�[���!�fy�'���'�1O�T��/B�IÖt*A	ߡA��@hZ���Q`Ϛx���?�����$�O��a��\�4E��̺z�v%[Qf]�%<r˓�?���?I���'p~�Sv+���b����>�> �c��SH|%��Oj���O���?1��ě����_���Q�1�W�,@Ʃ�䎉��?Q��?�����'9Be@� �≑0�m��eD5�<(��^�9"�'vb�'��\���3͟0�I🬪rK�����)6��۴�+�K���I\��?q��ܺW H��O8%3ve�8`C�mص#�Ԫ�y�'RW�T���|�Y�O2b�'�tW;�(A�7c?�<���A��O��D
K��yS�ԟ�9���`�9���DL���T����4}0���ܟ�������SJy�IYZ
����2�\�!2ʮv_�Iǟl����WD$b��>��E��6�Ԩb(a��}����O&�Q�n�O���O�����T��|��WD΀�֫���ר�a�RЬ�Mh�"~eRl�<E���'����t��4Ut��4��1y�=���'Y��'�R
�sL�i>��	�p�.��q(��(�����hλB�r�U�!扁F��(�����	ן �IܼA��2Tܩpꟴ 0FTYc�şL��*8���'R�'�2�d�K��Ŋ&!�C~hr1� �3f��&|{x+����	���'gjH�s����#F!	N��:ÂT4e1�)�']���ʟ@��p���?��%42O �ȃ��(�Ԡ�%)��~m��p~��'b�]�@�	����̧M�͹wK�a�� �%�M�(9��ޟ��	П�?	��!��y�!OV=��Hw`[� H�T[Z�qh�퀁����O��$�<A��:��S*���$ܪ;Xa�Ŏ���)sa����O�⟄�I*��a��	=}��n^9S�`T0p�F`ZǏ�?Y���D�O������|J��?�����5S����9
�1�kM:�.��R�'�\�Tᔢ�����ϋ��4��R�R�
��d���d�O�=�b�O��D�O��d��T˓��`���&6�v��#�X8\��.O��䆣Jd�����IIh����ā�j0�m�G�M�6�B��G��'�B�'��dQ��������&+���b�`TBgC��X��}@�b�"|��q��y蒸9���X���?���?�6hA4��4�����O8�I&e�$=i�g�	]��xF��' ˮ��a�$V9�P����$�O��	q�6�@���e�z�B&�3XV��}j�c)O��D�O6��'�/{BR�jj̋H�N���k!
�`O���U��?!���?���?�(O����б)w�,c��q��P�R)V�-�(˓�?���?!��'�n����]�n���)��� U��ۗ/�}#�Ob���O�ʓ�?QO��?�`'��O)�۴o�/wxF9jw���?����?y����'�B�W/g��a	̼RȨ�	B��suʄ�$���v-�I��`�I����I� 
��^'�M��?	惞�*eT�c:�hq�b�\)�?���?������O�Q�5�T��d�Dr�E�9�Tp�*[�.A�c��O ��O����O��I���զ9�Iٟx�I�?�8.�Y��0��c2�4⣦H����ly��'���O�ɧ���L�!�H��E@ծ\�r���k��7�"�'ҏ3'xP6-�O���O��	�����_��(�nZ��$e�GOоP����?WH{�?1���?i�Y�|L?�R1���"D�s�˦cv��%�'�`Ũb-`Ӭ���O��D��\���O�d�Ov�͗�g4P�dF9ϼ��Ѩ�Or�9`�On�O�i#���O� .����0@}�t��/��pCtM
p�bӌ���O���O�]����O���O<���O����-ЕP�N%�@��+�O�D�<��ϊ����?A�Ӽ{D�R���������|`{a,�*�?a�A�H��i.��'�2�'�맲ybO�;wDȢ��K�c,��M���N;K��O����O��$�Oh�D�O�ԡa$�,{��T۳M�"j�>�����	V"�n�ٟp�����I ��i�<��=aNLh�����1�1��D�}�1��<a���?q��8�?Q���?���T���iL
x:1�D6kﰌ2�I�	O����'eb�'���';�Y���	�q
��$Z����7@��H��� �!� ��Iڟ�s�%�����	K�i��P6��OH��	pz���A|¥{'��-v2���O��Orʓ�?�Pn��|��O�]{O�!CW����^8����'��'���'��O�6��Of�$�O0�)��%^����
�$��p�j �f=���OR��?y��|���?��O��|*��[�<�Xr���;��(�H֑�?����?��ȉ����'sB�'-���O�b��Y���#S'A';?tБ/Z��	ݟ�KAH��@$��~���۳9E�-bEϋ<����'.���?� j٦?����'���'*�t�O>��'��dU<�*is�K0�X��.ZW�B��vR�'��i>�%?I�	�T���W��7B*p"&F!rp!Q�4�?���?���
*�����?���?�IB�ʄO�b�����H�LZ����?).O�9ړ�'�	�O��dc>yW�˞O��c �I�|�*�J�O��D1rj)n�|�	ןl�I)��	d���P�P���aө?�&Y���<9�@�x~��'���'�"Y�n���z��&up�)I��mR�Q����<A����$�O�$�O4hÃD�Q��Pj#KA�=��� i�lp�<A���?�����D��F������FV�$�0ݫ��H��<�����$�Of��O�٩4Oe�T�[�J���S�!ڼj���03O�O��$�O��D�O&��<�_?m�I7v_
�Z2ȅ9TT��"W�^r������ԗ'Y�'�biO��y�U>y�!�KD๷�rC`�����	ԟ<�I�t�V���M����?�������<8��â`)|�jQ�E	���?������O���t0�B�$�<ͧ<*�m����,�m�%��6X�"u9���?���k'-�ia��'P2�O���'ϊ���`Ɩ[�
E��1x���R���]����I˟,���Ğ?�K�'�'6��J��;�ERE@�Ox�JcBC��I����	�?���l��쟤�5�G��)#��/:�=���\�$���d�Isy�O��O�b�ˆAZ�lD�\Qf���I_�4��6��O���OT}p�����D�O2�d�O<�ď�d�k%�Z�~�>��s�/���$&���V�̓�4���O��d�{��8�iMv��i��ӆ.X��O.(R��Z�����	l�!R�rՠ�A��j}>�J��N����'�ԁIv�'g�Iܟ���')�<�&O�)m���z�뀍�2�
�Xg
2OX�$�O4�OZ��O�s�FE�6z<�����i?�]cTh<ugV��<����?�����U����)w�p��7'T�r��)�d�B�D����?����?��^wN3��]�v�sbn�z����A�
� ��L+O��$�O��$�<A��șig�OM�E�Giٱ(EN})V#� ~B��v�'�R�|b�'��� k4�t��A\�D���2��- �j����OH���OJ��1P���4�'Z�$��S2�p2A}d�=3�)��c��'e��'$�ڙ'ɧ����(A7���҅�!"H��i�1�?,O��B!d��}�O_r�O;8�t�A�6�R�p�,@1���u�p�I��p��4#6�	v�IŢ@i4$�D߼ <|2�HŭA�p�	$fԭڴ�?���?a��iA�'��(�)�ĉ
V��A��kvK\4����y��|���Ot��Lzg�LAA,��e�j���-�����؟@�I2ؘ��}��'��Ā�O
��a;��D���Q�$���|�Ԑ4��O�"�'��i(Q��<���Ԅ"��Ks�����' Ԉ��<�D�O��D9�d�<\a�%�U@�C�6h�#ٱ`��@�Γ����O��d�O��:<�ؠT��%�IR@k?t�JUJ0��	6�'���'|�'���'��`JwEµ >�8�b��/ո=K�&R��y�S�L�Iӟ��INy�gN�L�$���[�Yc�݀T�p�@��d�'�R�|�'���_#e����Ld�ӥ=O��
�2��D�O����O�ʓlR��;e��Ό#�TC�a�>#��|����@Bb�'�'Cr�'zu��'���2�d��Y�.{��3�JP�i���d�O��d�O�$��`�$�O����O��ID�s�2A	VÈ/*��t�3��O(�$�O�U����+�1O�	�6<�$42���3e�d���?z�BX����R�M�,���d��*��'r������5.��ZT��-P�5�K>ѡ�����L�	Y+xh0����5v���P��O����'�OR���O��$��f���	�O�XQ�\;�P�2iTKn�D��W^2K��������v_�{EZ%qÏ�K��]I���M���?��}:�ⵝx"�'��:O�̂�S����AC7}���J$�dK��1O����OP�M�g���e元tt�(J�<�d���O	��@�G�	՟���t�Ik\�8��"\2>�FU�4�N*|�'^Ԣ�y��'E��'i�@�? �-Cd�ېq'ƨXE)%{�I1r�A;LN�O����O��O����O��S	'(�����Nb����K�+1Oj���O�d�<�E��[��4��5Y�ș�w��u��ř�
D���O�d,���O�$����&.J\�x���0_�����3Nt�	ޟ���ܟԕ'�V�s5O:�)������LN��4���J����d�OĒO��D�OBU	�����k`�����:�6)c5�T���'��X��I�iƠ��'�?)��=;���!��V^�a���%���L>���?IP�]���D���u �=�4�C�P���?Q/O\yp@����їO�"�O������M�p�i���RkR�E�	�����)-B�#<�}r6'b�`��5mˬB���;���C�>�Ms���?���0�x��'!�8AX�<�Fo\�s��@减!�"��O>��ɤs���$͂}tZa�0*&<=�1!�4�?Q���?�Ak�8Z�'�R�'���b�DQ !��K�f{S�Y ��O~d���O��O,Q�q�>tYp��R៭"~`Ac��O����=�&���I��\$���B��"#�ā��޻(�@�@Dy¡ܨĘ'�b�'�2S��%��H�F,K4z��P��yr<�I<���?�N>��?1�����g�+[(���'�f�*�<����?�����ҬWTJ��S1#��ᨵkڛG�TAq��9�R˓�?Y����?Q�O���RPƨ`��x��MIE��%
.�'.��'��[���1)�.�ħ$ ��&�0�aFr�̋��?�I>����?A��q�]x�㑍��!;�e�GQ�ot\U�����	fy�Ŏ~�������a^n�A�-�J��j&1��O��(��Ӿ!7����e���hBu�
\���<d��5e+�&R>a�	�?�@)O~�m@v��Hr�ɣ&(<jC�'�"�'su���)�M�Y�����A^�c� �7���`h�6��O�$�O��	R_����0X�bB?b� =����5@�P�)�(N���f�6�S�O�lS5��(įV=��`��!$07��O����O� e��f���	�<7I�6dPx�9cM�2-޴�玐m��o� ��<Y��?���m�!��K&��`�%�?l��� ���?A��
j\�'���'��'�~���JG��SB���8�$X�X�(s&+ �I��l�I�x��⟀��ŜS_�\x�ڜa�R���yp��'w��'S�|��'R��.!� (7�ÒB����!=�M�?���O����O�˓-LFL���O�n}��dHF�X�� �+ϴ%
)O�D�O��$���}�Z��8��e���9Q��&�H��>ʓ�?����?����?�Ǯ@��i�O��^v�����25��a�a�O��d%�D�O�ʓe�4)�OT� �^vYZ���Gޯm�Z����'a"�'~��sh�O|r�����)Y�2h��	;M�,[T��䓻?Q�V��Fx�O���֎�*Sm���AĆ
ݖ������":yo�C�T�'����<���\�RP��3T?c���b�A؟@�����s@�5�S�'A�L+CNݩZ`T���<(P�I�T��qPٴ�?����?)�'r)�'UBȈ�Ttd�h1� �!�#i�S����O>E�I�V�F�`��E���s�*��I͟<�����k�NyRT>���<9D�_K��	G@�g�!B��H��j҄�<���?��>;�@#T� FX������\P!���?�u���?���i�O��O
�z&Ɠ���`8���G �YH/��]4q��I蟄����D�'*ơ�U��u��xPo��*
���bȣR=�O���OZ�D5��)g~% �S�8��+��R<T�TU:4�0�	�`�	������EJ��|Q�́&
��1�Ʊ�������	ݟ���|�Iݟ��'P�i�4�^?qtɺ��"4�pI� �%*��Iן��IΟ`�'�6�£e'�I���ْ����xQF� $Qm<���O�O>���ON�P�Ę!`�:}�vk��	N��bS�)���'��T��Q 
���'�?��'eĐ�#�J"����N�,�hH>���?YסIF���Ԯ!�=�'��(.��s�@1�?�)O*���+���O���O9�?����D��L�li���
X�^4�	ޟ���0@�f#<�}��@6#���26�T;L=��ǣ�ܟPQ��؅�M����?���zg�x"�'�z)G\���m�M��h���E�'T� ���ɟ���,(����Ʌ��{1Ȝ��M���?��4�Jٓ�x��'	"4O����,֟gB�!@CO�	Vm�5���:,�1O��$�Op��ْx�bq��ˑa�H<IA'� �����O�(Q���O����|�����Xd`��4U�����ĜX�~�`+O�T����O����O`���O�E��l�\��ik�ABl56�@Æ�}����?����?�K>���y���G��E�ōS�`����?�ӡ�[~2�'2�'��	�7C �Z��J��Ȣ��	[6(�B�+��n�"є'$�'JR��R�k���0f��}�@Q�.�DL3�cѹ?�ӟ�	ޟl���$�Ia���'�� b����&0-`l�'G�l�΀�$�'�ғ|2�'��� c�L�'�&�XlRIt9�Ȗ�v5�X�۴+�E2��	�$�G�L`�2�Z!	栀�������w#�,�! �'@."u�极7�0�R��'.b�'�䃜'���'2�V>牀{���.����@1�G�6!���'[´i��7-������ԟ4�Sv�dAwp<��3�����-�?)�.=��3�_�[]�[�ώ�y����'RgB$�uM�"����`9Jô�B�'�l袣��;XE�c@b�;Kc�y9�O�:NX��}J�N�B9T��Ua_�)��U�nޢ>���@U�S4��[GW�M�v$K�d��=,��������ޢ'�:�"aH1� x�ia��}�*��!�Tq���<$�L	peȄ9q1����iA%uJ(	��]�d��6�����c���e1��I#G\D�I��O����I��a��B�\�b`�X��R�	�16�Qc��`�U�6�M-"����)��b>7��>��1ȥe`�tD����қ�B_�2�hL`��8���REڿ	αbX\�%�|�1A�.���o�B�E��oυv�bMn�1���$�O��S��~≖Jk��� *�S�P��@&��C�I��֌3��E�`�!���L�I��HO�)gӼqH����*r)�^��u�[˟<�I#H�0��ΟT�	�t�	��u��'���x�����P�@��c�S�F��	J��y�,��Nt��Q����T+ n _Y�H��H_:wE�i.�5��ѱ��C$O��%u�D����O	~���R�@#N�@�vޙ�" �.O喡� �U�|����ɨ>��Ο,�IS�'N���<����P]�<=)0�Y(A�<C��:XF|�AQ˅�D(M��nW�a6̬{��)�,OLX�����F G���*Ʋ�AsjFNS>�f(�O����OF�dO'X�J���O��w64��4,X�FLmX���P��`�3M �KCа�c�P�.$���j�'�ʙH�዗q5��r��c���.5	���5�H�f9Bt���C�Eɗ �f�شDx����?��B�=�R��g \h�إ"�˟(��E[ךx��'Mr�T>)c�;?R�x�Κ�<��D�!<O�"=���
�R!��]�:e��E��N?b�i+U�ԒF���M��?᪟Vu��d� Z(QՋ�q[h�+�eU�1:=��ӟ���=+-�])�!:Je܁X�鋀E>�I�O�c7�Q�+���:�cل{��H��$�D)N1c�.��u(�j3J�$T�S:�E���.fA� ���"=iu%FƟ��ڴ�?������b!\x{�!L=o���h7G�6jf<d�	�����͟|�i>%Gz����
��Ԉg�˺Vl(� ��O�p>Yc�>1!�I7w��ܡ�I�$->L�7K�$�!�)m������}�$�Ƹ+��'���B/bfx�*BH"�*��?��;E!�!�^y �!O7;��d��|��ܴy�f@��%���L!`�׿w��m�y�j����ҏ9T�xcd]��ȟ�fXK��Pí�	+��:���M[3k��t�Ih~J~�����
4Q��sg�8!,�y���\!򄑯;|��l¨$�Mqs��(Q�{��DGR?3 ׀5|�  RC��'FR�«�;0]�'�����-���'B�'VP�]mZ'�����۪N4b�J�g�T���q�'�|e���&C��iF��~FzB�$���G��%Ñ�O;�R��I�p}�"l�+�60����H���4^������y�x�Wˤ>I��� �I����?a���!b4�&eT4c�#M�y�I��"O2�a_�a!Ё� �&�v���'��HO��]y��n�E���@�����*@���c�BmD��'�R��e��5�?)����$�ԃ*�3�ByȆ�KD��<��i�&�Z���є
�s����]��ڊ��Y��(R��e� �C�œ28{&�X`I�<XR��$)L�p4�7Mßjč���	�Oަ�Dk�x�rr��Gv:y���3^�>@�Џ�ߟ��?Q���'Ԉ�Kҡ3~������jk.�0�'n-���9L�(��nX�+]l%;�'�<����.�nџ���k�4��<�ڡ*g��>����A`�"�D�3�-�O���Ot`c"� 3�!J�����B`�~�pl{i��N�r��KF�H�= #=�#�(~����sa� H��C��Η$�����1I����2�Z�w�d0��#V����l(T,�OZtm۟$��h�ĤD�f�����e�2*�x�� �
Ll���O����O�4��#=��?d��u�!/P<v����m?�@q�P	�O�\X��04̓/i���ڦ㉣	�j	(�8O"�ѐ���9��ܟ��O���1�',�ibUR��= 윜�#ȍ�Rـ%擱4��`b�D�*��A&Q�h��ݶ0�^z��ܴd���B
�/zf�Yf�^�u"V�m�p*�1�F�O5"�Q�H ?�*�]eG�q�}n�1��I9`�V�9sZ\Q'��S��7T>)�/n��@���'�B�O�QէGZ.Ě�b
-ur ��W"OX!�����V` `oڍ(nj�[r�d�O*�Fz��jӒ7�A�Nxa���N!6բA�S;p�	ʟ0"��p; e�����	�઩��7MǯI����aA��yR��@�5B�L��/��Vw�,���Q�.��[RQ?#=���͹@y�̈�3t��-�j��)����A�o�X-��U�2��t�O?�x����.��NY��k�$GVIV�{� ��	6`���'Jp�a��'q����,O��Ī>� N  �?n�rPq���l�sD
O6��XR��@]��C�W� +��k��$�n��<�PJ��3�lqQCK(gx�m�m�.QP,m��ን�?����?��rbNly��?��O�[�`ɞ S�(�b�B�d�d`��Ni�X9Ѣ���7�p:�'���a.�*Q�(@����k���q!�.��!��@�6X�6���"��e)�;��hՈ�����w��i`~�{f��}:q���@<�l�F�O���E��5�}���47Z��3��Ӗu2�ȓ�N(А^�n�Lk�&�a.�=�s���'�ɏئ�sش�?A�����?"��"���4�H!�u#�/d�> ( ���H�	ꟸZ��M��&��o͝��5S�E�+��$"�R�B��s�.<����#O=�HOl���aβi�IXR,Z[`�Q�'�?�k� Az���)��+Q��c�h9ғD��m�	�,&?1l�&`���)�!��@�hQ�>)�Zi2����������;Z�J��!`ثU8<,��.�p>	G�>��ќ9�n���LT�K��m��^?�
��`����'��]>�9&M�����I����ΚU��g�>
9�@�ä�'�r��bc�6�y���i?�O1���'� (`��4͘[�>��AI��Ms���J�dp���߯=W��)���c�gHMp,1Sh�-IX8v+`��p�'�7MOǦ��a��M�Dϔ R��9�\ht��TM�E?����>ɗe�X��aS&��c2ZŲ��K�'��"=`b���	2L��ܠ�
�������M��?��hR�@��՛�?���?�y���O�7-]RqVtɠ�K�2Oܑ�F�X6*�I�_0� ���=C�\��D�Zw6X �I�7gZ�ŋ􍚬��	vV�BaMP�N�����İ@Mp���$9J5F�� ��_�L���L�	�I��M��~�'��W� `��I�LU�-����j�� �=D�����
�9�`�h�@E���"(]@����aB�O�|l��x��
{~(��V3X���S�,ƳS�be����?���?���?a��?Y�)�8����`Eh��E	�EW� �0%дH�2I���U�i�~XKǓm�Tq)a�w�aɥK(0��-����{,
�"�~9@nT�.7�$�ZS@��L>4�\����L�X�l���ď<;P�xb�2R4��4�?�/O���1��|Bǥ �N+����ő}.��+ŉQ�'��IK�'X�1;��Iu�Ai��Q�it>�%�Oz��V'�֦y��3�MC��Q�	l�n�O��$�O��1(F�1�0��¯��@D:s�gO��?y���?��@��tYr��U���'��P��)����)VS�Ը��J1�P���S�{
���*����0��55(q щ��4��D+O-�4�!�����d��O��HO� ���'��6��ĦQ��\���P o$p�D��D�ڣ@Ԓ�4�$�)�� ��+)pU�ɫФ\1X�0
��?}2�i>=�O����X�]�&a�����yc'%���nZ&$�P�����4����(���Q.%3�X�l��Â9�' ўb?	��F�)��쨠�׽2���#ˣ�p����Z�����^���>����̥�j5Qva�<dj�U�ȓ|����MD/	���%�a{r���
a�Yu�����%��&{�,��Qh��3I��Lpr	*3C�$8�T����pQ����i$�u�E),L��~@A�%��&>�Ĉ��f�����c�ڶaəY��e�� �Ʉȓ�r��ĩ �g�\�)U����܄ȓ�Ll�tJ�pG�@���c)�0�ȓE���a��!'L(�
���/ �<��ȓ|�x���P��:�l���~��ȓW \���㙇F�`�
ң|�Du�ȓu"q��A�~@:(͟+���$��x�d�645|�a�	E8j`�ȓ,c���
K�h�!ڑ_"ll��\�`���L�$!��ЈNY����h2�����M:r�h�C��V����ȓ��P��O�/c^�VK �#|��ȓ-n��J�Æ�=|�(��
:w<�d�ȓ	6��{ U��dcL�4OMn���Z�Xa��	����ֈ��Q:��ȓe���$ήiA�=+`�y|HS��jK��D��#�������O䭈�ďe�޸���5Mo"���'�r����BVX�C!�	3�b=���z����7A	�)sKV-�����DPr�cE�K��1ۆK��i>��=�,ǵ���c"�
.�H��-ٷ]�pD�!H}>� �IaV��w�
,bǪ�2 \�"Oh�������dGG�(��1�� F�I���ypH��Lqz������+
n��$�8�	��)	�.�i.H�tH�X]�����4E!���i��ҕY����0K�,���q� Y$.E4}��i^�	�d̀r��
�I�r3����Z�Rm�0m��$c���i����D^0o��+eB7m���9��İe�j��k�8
����S
Z�$��Ǚ3�ޙ�۴��=���E��7JB +(��"����++��b������?u{<(��ɩPÊ�]�?a
Rb`�pA�*�;@��0G%,D��(���?x8p��s�A�i�[�z �g�>3R�A�$T�4KH��F�y�T�+ d��ڧ-|�E)�۫i�`25d�9n ~��'=�O��xgE��o�F<H��K=G'ʨBŧ�/|S����B���"(Rq�ɺ�e�>v�H($�=��v�L �S�i�Й���W�0�ӃA���O�u���W�?�p�p���`x`8cG^%<�:I��ܭz���BjÙpu��X$ җX4���	,F�4�'�l��%OS�ژ�M[u-
Ecvp�WjG��ॉ����<ID&�5}�hx
��^|������@o`@�
�'�챑�Y?�v�RNr�qE*���삄efӬD�q�	�8�F� �Ñ\�ay�O���Ġ��W�E�&�9����HqO�$br4j!�����A�~z��!U��8�$�OrZ��E-D����&,�28�#cOTxY���;�&܊��K���}24%7dKP�@�kʂb�X�`*\'F[BP�$����`� $��Q�D4aM@� akK�d�h������[O��S�^.b���.>�|����_gLmآ+�����Q`�(6?x��M��
Xs�Ǐs��C�9b����A�E�~�(�[33f�sVP���G��D��~u����_�4�RaǂLZ�� /��ss�U7p/�����|p���^�2�JQC�"̏ZP��g����5�XR�h
+2r�٧���sЁSǍ&3���s��|��"?��K%:�ȡ�Ueqɨ8����8h�D���܊ZT�HI��*a����A��;�α�M��Mp̕u� @��OE�w�"�i�� ) �����&w�X�[gj��0?)Ǣگ���� d�H��N0w#���W-�	<r�Xf�I���0cGB�|���S`�d�T;�N��cuf43H%:.�8��x��+�s؞`� �T�nvv�J�
#ed��!U�\��@B[�mi`�Q�F��Vqȵ*��)�9ц�Gbl�Ӂm�_� �0���nnp�	 �f� ����^�UWF���AU�*�z4��]�|)�T���k���B�֤l����MPt�V�Y8 \�<{��|��)����}*��C 厰1�L��'!��T���'��:Q�"=��]:<��14��5M;������޹[���F)x�ģM ��86��q����j[�08��99�dQ�%�"N�8�qW�Ƣiih�����!P,9�ԩ3�OrMXr�8+= �j��$c���W&tZ���c@�G,0[2�8Dda@�'�):
�B��B3%o����d�'q�hɃ%��m�
�1��������<aw��	"ނ͘�C�nF�Й��k��rëNkި�1��T\�|����1��H`��b�,15�ȕh�Z��χ fĜ���ɐPV�T��MX:s�����ã|�΄������|�ĜZ1�M�ѐ�S�J�9Lv  �'��(m� p�9uX=A2��l]
p��b	�@|�Y��#��e�&~"��i$a�sR!��_�'�j��;:N�}Rg��5e��^>h}�G�ܟ�e$p����l��2�7��~�؅y7�)�r��1��sA֚{�(D�B�3>
ț��nr��w.���(O L�b��l�<y1���9�����Q2wc����CL�g��P@c�+~8%{7�ʋ
7�`a� ��6���#�3���b7^�!`'#A�P��f� :d�i	�f6�0�'���2��m�iЧC�
>ڪ0s'L>)��8�6���x2䉰��O�s~�ՊC�\�%�ƈ*c�r���ߴ[|С��D~���z"�\�=����N8q9��K����#���Ck��-r�����9t?����M�#��=�b� ;��k��	=:� A�Z�({�-��8w;�ɳc�"��	����)7Aip��Ylj��%���Yehu�R�r���E��Y���ՆW*3UA�}B�
�C ��XF���E����Q��Er�ݹ�`�c9\@�jY�7�H\���@�e4`H���f�)ќuz49x�#؏~Ƀ��ъztX�J�Ï1I��иǡ�j}���}b�ZE.��!+�<�*=s�����n����8A�B(uǮ(�"�W/�>	�Q
6*�JWL��*?~�r�����(�ètƢ0�rW�+�*!U��)(�	$Ŗ�x6�E� �<iP��b����6<	|aŧ��,!�!dE֒{1�Y�C�W�Sv8����]1_����¼}Υ�sʗ�R��x�Eʞ: �#Ag�<�`����4T���p�C=~Ľ����M��	b��!�Ҕh��=3î��i�:T� g��2a��j�2��&k�&
{R�Ȓk��k�.�3i�"6͏#��TK"n%a�D�� �9S�^�P,�6"��p*�n�옼Su�T���d+�{rJbl>x�@i��5�(����6�K2�5�:h# 	 z��L!Ac޸ o0d�)�2�$���^؀�n	�*H��CX�X�Pbpi�'%6��(��0����K��qO��B�%S��`H�H-r,jr�C�a�.�kJ�]d$ ���LX.�$j���ܙ��!yڰ�� ],��+�Yj:8�G�M�[)�8R`�Ӟ
�D��[L6�B�a�Z
�\�#V�8�`��$Drx���P�˗���	��mJ|Rw	+u�4�¯����c䂜)C���B��R�-�>l1Ы��@,ʩzt�*q� ��r�B����Sd�]+E��6��\*za���ùd���pQg��fk���%�V�	�"�v韍~f 0vV>5�0�Y�9D����!pz����h,P�O�*-�D	�ː>kh����5�>��P�E�1�3FFn 1O9�s�r�`�!�ֈx���0e��Kli�L��E���N�V���)�#:��#����B�ӜO��@b#H�e2��ЦߕXKR	"7�� �6٫�:g�}����'e�m����v�PxK�<9ȼ��f^�:6D�s�M�,�Z �1)
�*=戹#�?3�И�",E!����"cO;0F�3�L�(�J�qIʚ+>ST
("�0�Д_�����Nq���� ����v�Y�j}2�[`��`(�
/m��Ӄ1+P��PLܼ<��Ts� ʱ.�����F�&����C�O����
I�*�l`Rl\<=��@[��0/�����OƦ �"(�y
���Ά�'�y���>s��ո�`�~�~�i�/�v�c7h[�x	����$�Q���<w�k��fg���Il�@�����_#�}J�M�:�̀��D=.�dD�e��&em���*���3b� ΄�!�4�h̛�.W�Z�J�Pi^��S�̆�o�nA��l�0	�д�a<7�n���'[�P-� �_����C7�i���(�HPX�8|�}�g���.��VE7e LT��� Gvt���gSV�M0����3r�!�QL|<9h�Q�b�������d璁U�M8�hK�4|�a�ѝ�"e�9u��6��=���*� `?����}u�m�5��3�����<r@]����\\JS�+���{���.u�b�!rǋ*i1��:���
�*�!s�@lڥ,C�� S���g��ŔLҠ� �*Ƞ\7N�ٰ�˩`Ll�TK
t��<��#����BA�H۴�pw*I�_6F�� �J*d\H�-�kZ����	]������l�ąb0�D�?`���(���<�E{"G�s�����P]���z��B?A�t����_���%�.�,��C��4m[R@�e��X���"qK�<G�h�VD6Z��1TL��D��L�T��F��łu�S�B�����hU�m���(T�[��P����y�x5���ؼ�2%��A|�o!I߄�[���h1: ���9 �n��ٽ�&�F��Dv��c�M�K��y�R@g׾�*��J�4$�\�OB0��e�(nSܽ	�dʖO�Ty�'�1hZT��fE�A�H��nʔ^3�j��*l:���a�-��a�3���Sp��0�a)�i�[+��< $t��x��^ 5��x)V��G ��15����	p���f풀[$bޞP�����߂0��Lq�.ɻD ��Y�ݝ�MK ��~4�� �Y'i���
�o<}�נC)�Q"�IB��Dz"�@7����Jy2s�L�|�P����qp�qiԧ1��`�穄���&�6(8��Ԇ��6���#��[��l[��O�t0 �ɻB*�yc�Q)Z�T���h'�D88p�\#����蔭g�Pix�#�F�j13q@\�x��!�A�Kؽ@����
֭xQ'H�R��J�$�B�|s�\	~��qE� �Lҩp�Bj4��$j$�@�ͽAe�@��OD���EJ��Ðd�V.z��k'�H�OCu�0�âB+x���,�x�
�J.�`�m�P4@���]*�}�u ���	��EpQ����bޖY%�'׺��iO� ���H�D�2b�D�� ��p+� �\8H��I&4Բ�2≏#��� ��2d�T2�-�'k.�S�
�u��a"G+,>h�Ibf�;���h7�$vl`���F\�'\rȰ�� zȠc'��(���R�lA�A�!(�4�I�Q* .�&]�f�&�ȸ(S����28�B/5nF�eh�
0y��9�$쪴r�-�ma��dH��r��O��#��>E�a	E������'vE��@OX�4 ;pkT�-Sh�!�$@����Ah±�\���EןrO���oY��6(#@��.[x�ͻV�`mq�i*&|p3�j�2o�6(�I�&��2�bF�e�B�f�(�4,yu�sʼ�m�)6F���9L��X� M�ڼ�ZaD/_���S��	w
ޔHmZ+3R�ʥ�	A~B��v��L��j�.}A�� ��Y��j�pg��4^�����dXtf�!��'v��T/2�l��l95Ɉ�xģ�9C����֯-!Ià0BQ��x��Q�+d݊�BP�
�!D�N��d��T�q��U�hpc�c�b�F��ƞAy^A`���59j���.ed��yD���bl;Cטe�R�:�f^EsHuq̆�1�vp ��ϛ.[x(���P�9�*������OX��@�I�3U����#u�YB�O�R ��	�#��� ��K�6ʐӲ���
������
U��tC�ͻ.�F�pI�!���8�K��2Ҥ��w�v]��-��޴J�^m��ȟ'ߖ$!.�*��p��~U���c�1_P����ϬQ!�ŋ��	纼�p�/FR��
�)�ֱ���J�04�Bte�/T+����]�	���:�y�%/tK�Ps���҅a�ҞDX��B�D�5E�����A\��g�?��	�-��|lxT@��$Hx�C�
� 9� i�l� -�e�U�ƽ'���(�c�B�v)�b�6�hO~�!	(:�щ2'F�� ��Si�4+��T�c�Q.yri�iC�8��`�Ҭ':�ɉRǆ�(��s	��)��H�kQ3lt!7ݽ=P˴��5�ܑ+�f7�e㬽�� d�����&R;���*֮'K,���]���s6�ыm�r�*DS+E�2!��oμ`� �����/%N&�$�� _���#�,��y�e�6��LS��|�u%K���d
�0B\��"��)'�y���?����G�3�=IV�A;W� �Ǎ�Pd��Q�`� �5n��H�#&I�5��h �Q��OR��W釬�����$"|�&��fH�+~�r�� �'Od4�wM�+m�R��	���ീ4G!z�.��fhD�~��5CtKߙ\ά$���0X��W��`D�O� ��E���0<�3�Y�Y���Æ��_�Z	����b�Z *��<i�n��)���¹y���"7���ˆ���u7��L2ǰi	�#��"�� ��O*eMџ���8��P���-=��9)����qBT� 5��sk��G�|@� Ѻ-R�R�Ë.3��!��V�q�'Y`d�QcH??!FOW�:��1$-z������Zy��_���rv��5mb���͎��ħn���'�[6nw����Cdx�"��ŒL��G����օ��Z�F��q8�x�j!(�d��"BK�
UPa����46�0��. ��� ��?r@�*�� ��Ê
(-,֝�;zPd3�
qx�h��
ٍPyh�Ab�v"h��Ʉ������M�x�ԡ�6�P�ʌz�P�LS�0�'/�n�1��l %u}�DŌ�|�Ɓ���Έ�O�V�8&˰���m��0���;���X�.�Vē"�� %����]5W$����=)v��`��)z��uA�^��ͻ���?
�@���)^����b�����$�晫��6mvBE;d'�<�G.�UӦ�Y���b:�H�w�����O6�h�W�-혝8،Vi,�A�ɟ�/��:��Y	"��p��Z����b�Q,$���z�n��z�,1��M�*+ �"o.�2��	�2=�4�}jz�@���=N��ᙶ��O�H!R�EiJ���c? ��O��PEAԊ�tpp�e[�+��}1&a\)%�N�� ƅW���2baz�@Ty�
���Q9sp�ᣃ�D�p<!T�Z�F���Y7ϔd=8�d^�7"���ł^�?�0�&LM,�B�ɸQPɡ���3t�,�B�̫X^O�I�%�S��J��«;�0=F�t�Ư1����,7�p�jA���y2gо__���F! X�i&	 09tͻuŞ|�l�H��E��OZۇ�p����B��7��ZD"O"E�#n��}�\�@H3�Jq�e
Ҥ<�la�gk@B�<k�S�? ����#���E�h�#-�V`9��'�� :��K8]F��v�iqrӧ�H+(��6��8`cR9�
�'�����#��AC%�@�:�ۉ}���O�p|��J�R�O���!F-�k�2�*�Ǖ�Npl
	�'܂���M��wL 0��*�@����ȫ�&��=E��'�~�Ԩ6y�|@5	G�H�Li��'���t^yt��t ���'ɮ��aA/g�ж�C_�H%�'tp��U�Q)E�(qS���)Q{b=��'��&^5b�Q���^�Q��(8�'8�h�EG
;��1�%_q̔��'i�Z�h�XlxF,K��,��'n8��	��*{�0Uo\�_�0��'-^Ec��Q��/Z�_�E�'�f�#�DޠT�Th����IM��(�'�,���]�!�ld�'O�?]S8$��'n��֤I�/P�	��3VH�)�'��� g�W�8t �@M�KJXi�'�NՊ��Y���積�{g��'d�Th��%L�P҆@]�eǬ���'7�Q�p���!"�+g�V���'��E��Q��rc�M̏LeHiS�'����Q�E)^��e�e�]�_�ptb�'g�#Ǫ��I1B���G�#l�`��'�v�w�
X�dI��֨%Xbiq�'��Þ�j�|�Eؖ*�4-2�'dA��e��BE���c�hب�y�΄qg���۸A�P� ��"O�m�HM?9"��`�ֱ�(`He"O �C��y�4Q��](�%٢"O�P��"k�p¢pgB��"O�<@�.D�kP���B	�JV P�"O�<�
��n0]�F�x]~�j�"O�x��Ӡ2�9�B.
AL�E""Ob)C��"G"�Ӗm�*L:TL	c"O��0�A��[9x�Z�셳iq��Z�"OH���"�5�FR�Kumꄀ�"O"d#&գD�,�����$%D���"O򉹔�V!����1V�]&�e�$"O`�( .ӨH1Z��I�	VG�� "OF��w.��pR�t{��.�d8�"O�h���x,x r�\L���D"Oj�2�(�13_�V�U�z�r�[�O���2(�7�\�;g#w:Z�9d��2�ջ�ǘ�E���AaEH��B�	�h��<K��N�X�C��98B�	�.��d
2G�+![�� ���6m��C�ɓqB1��Hٽu�MؗG�U�xC䉖��H�'�γ4r�s���_ZC�	B���Z��Q"W�:�I� �X�DB�ɂd
�(@E6(�H)��N��QP�C�I�-ND�Q�މR8ڀ�3��C䉎NA����qS0�#E�Tp�@B�I$p��iޫ}E�YAѭ�:�B䉁;P܊D�!ZE��`�(.$C�I�}P�<�E�ަe]0�c��<��C䉴u����-�`�Ax�C䉤l����F�D5\]��Z�J��C�ɢ9�N9�`�e+*��R��*|RC�	�:�v��ӫ�1"$�ؖ�֏X�B��+
ۗ"�(D9���㥏�^U�B�ɂCFA���ԷIͤ���%�IzB�	�zݘ��� Ƞ��"�]�6!B�	�bA����H$�ԏ���C䉆��man�i�,Xc�Z<�C�)� �|�VǓf߂�A�Y�
ba��"O2p��(�D���ݷ9Z��:c"O�XQuώ�%��,�U�T!ao�Ps�"O�`��F��0BHՀU,�O�D�F"Oj��!C�$�#�� �S|Ph�"O�@�����2�F�2?*l�zC"O$DK2]���1Q��=�:���"O�����J�F:H7X�v`$"O��5i��}T �)}�����"OPy2T�P�(˧iM�L��\s�"Oj��0<!�a1��	$%,�3"O��� ��ju윀u`R I%���A"OHh�oe���+  !(��"O%�M
�p���)�n�.eYb�'�lHB��|� �(�L��y��A�F�hSX㞠S�ITܓ1��dGy@`��4?���Z�2�Ѩ0c�H�'��@��+;�+w�	�J��b�a�"4��
0���C��00���ODj�-T�"]���H��đ�e|�P�,����Y� �&{��d�*%�d�q�Z�E�6ر�@�~�ўHʣeZ�'4�0"�I�V�mk����?yFK2o�5k��ʖv�����?8Kx��B�_48]:UG 9|����G�nD��>�A�#��ұzo�$8O�V��M��1C.���'���;rLi����Y��@��`o�b���
)��'%x9sy}�OX ���d�Є�Vr�����G�7AȮ�����Ol4"#˟)��y���I���'� ��0��7cjB��$C��Ă�H��[��$�?!�'��t�F�q)xMХ��i~�"��SPR��
�� h�X�d%��~��Š�Bg̚kA�)SJ�	�yAK"pμi�d�0�?�Zoz4�(���:~[=�fϜ ��a�ɩr���3��!+v�pt�'�zdᐞv���H��ʢe��	U�W�Q��k33O��K�TjE[��Ob%˞��d�w�ȅ��\&F�& 1��z��s��,�O� z�w��1' ��b[,�+qM��f���H��w
 hj6�O�5q�E��ԟ���I0W��g�	�"H8#@)łL��#��Q�pc4$��sB 5�V$ؔ+��8�%��O��١N�8[h�8�V#�0t�NM�b�؝��)rb�O��#D�p�`�j��ȉ{�JtX� S�I�
��ز?���ӺELXR�M0gD������$��!�$3�d�=��`��S��!͈&e���rK�4���D�	?�­*�N�(o7�L��|(���#<�а�	>eNy��*�`��8��'s�����8��@�'�Vi�g}bC�-*u���n Kj}�Rg
xktؠV�'p��26��w�K�_h���̜�f�s�#�/zo��$f�<pC�>��X~��$�l%�T'��ԨA�΅|������(<��öC{`@���V�,\�z��܏\9�ly4f}��O~��Ƀy�0|��#N4jP��`����7������2�¬u�F/��p1$`�[�?�ɝz���ړnT�/�b�I�� ���r���0!���٩Z��	�IW��Bd"(H�����'����JÇ%�@�ٓX+SR8L��;/4}ZF3O��p��҆N~���wڟ�����	i�&T�3%��m�R iw��Q�.M�$�]+G��-�R���$2شt�	�oZ"M��a��G�I,<k@�A�Ѷ}6�� ��xC2�	\ڟxA6(�,F�<yq I�+B(
E Z�e��e��D� ع{���W�9R��lK�a(΁�A�W :?9����R�$��n%�s#���?!��'�ޠ�ų	�e ����U',\.V�a �.�x�YD��>�,],V�c$�'nMx�[@�'�x�H��ܘ�`-��o�7��q���Ǿt}N�
�"Y}�y�U�w8��s�X������%� �vi�G*D1{�џ4K�/��,�ۧy?Yb�� uAX�Ə�2�	k�:�r'p��B���eָp����'�85CW�\}&��h��Ug�	�.���� �n �4E�t�c�دf�Xt���&ez�BA\�/HXh��Z�w�&��?�����?J2���&��"ߐ��0H�gl��'�����.��ީi��[������.�����|Ӷ�ar���C�	Mt�J�Q��d��,�0��$�l�BP�"Ӑ+U���S?0��Y�r �o�0��e��hW�O��0��ð",�T�ԩH��jMs�]�-�(ĮS�*]
5���ϖu'���dE�l���A��� 9��a��f@4xaV������|~Zw,а�"LƧS�d��	W�q1�v�L0k���G��-���Sv�
��=�ƃ%� ��r�|�,xH�$
�I��K��$K4f�cT�L�C.��Y�3o� V�
����x��k���)I2}4y)�h�)Y�vd�Ď��z��?!��K/zi�V��OL��D����"�'�H�K�aΉ	|j��p��-S�~���ܯdZv��F��OG*�0���H�I�i>�d��P� �3PZT��������SC�5I`.1�ME��?I�E�u����D����������w��-+�Ͽ}�&m�F��)Lm���Kǂb|���`�Ԍ����Q�/>axrEm-iz2i[j���F =eN]S�>O�E��H�a���Q��ix6aSJ��DEA��]2URc�ڛjs�5��/�|�Yaz�@��[<��Y:����:b]�uP�LȦk�.-*%��H�!ҍH'N�m���۰r҈	���(fU�U̧o}>h���"^�H�=� 0	8�܍[���D�A�g��9R��ǝr�*a,O I��(��<�Aѫ;����Y�p�� ��T�?�ȴ��:\!��J#�>�H��A,�������
)������eǀ�b������ �H���)��x-O�i!�J��<q�┺8�8�""�?����K�@� �@�($b�ˠ(C9�����,����*�H"�!UL_���'W�#�b1ョ�rgb �3.	��$1:�zQ+s.:C0�)G�cL����y� �e�`iȗ��'��{�B_;I6�<�$�2��s�'z�H�5�	�eI��+��'̼{�f�(U;��a*M�f˪D���̛��P�+��¤mZ�l]
�9wJ� ����E�tE�T�R�����w��0k��ɊP��T�%8��K���$:��+=	�r�'5 �Sr0R"��]���ԃ	�X��ę��0$��a��(	�����\�I�. ����O�I�-Ȁ�c���_�FEz�)ƈBL�ۆ�v�������OV����S�Q�����D7��;C���(���
eӣW98�Jp���s�9�F$�p�6<x���M�'��HkR' �U���#��V
,�D8h��[Q�P'�Y�@(V�O��-1�Fk�MU�e�@����E>��`4�5��@EC�<{��\�M��舍�����ھ	�I��G�+Y���j�C]�OI��O�O�!�f���2��~7
 �W��1��D:aB�>���O�E8iS�z~��s���?�7O&u�g'�x��iֶ (
��
�A��ȋ#��>AU�U�p�`�RGN<9,���0cKp��>?�\8U�-��̟'e�ti�]�m4���W��N��y�t�ƃL<�~�ǃҺ��.���y��y�ѱ�?U����O�2��!��$ =kP��QA�	�j����<=ḏx��U./?`�P��.;�R��G���Nİ�Ƭ@�a{�BA�4H��`�;)]HI��N�8��<��h�m�Xh�WF��7�Ou�����õS��Lc��@�F�!�dUnjP�`w/�xn(�(&�K$O�'�(�*��Z�F��m�O�Pe:�2R��cc�9#�~�b�'��"���{,�"G�:^���[��	���S����P��@�'yB��Ӡ,�\���r��c�Ꝍ(0@�!��ڐxHW�lҜ�Pc �*v����C�ɷ�tˢ�-q���`��Y8��}��Oڌ�� �j?���3�*�c~E�Hi�����'�~D��@0-����YC.HmR�A��>�dT"�̑��i���O��s �b��@���#�AQgyʟ�I+B4P���K��W&n��p����'�n�����X]�� @�+9��z�Sⓚ&�lc�I]LYh�c;Y�d���V�62�5�08r`������Y�t6th���6+� ��u2��IcK��>a��!�?Q#���ĥ<��j�8F�dj�I��ۆ+�>�q
��&�}��iQ�|��v��'�N�p��$^Rܙ qܒ_���JD��Q�o�S��O���b�J���1 ��q�J�6u�*iwuzQV��|�'[�p�`��ݲ��^�y�풉��D[�BƈXk�!h��W��?y!II��qOL�)ʊ�?Y'Q>?�|�r��)�n��c��9����b�B�`X�&���f�R� �� ��F�~vؘ1��O�,OJ���]��0�����|9��Q��ǅصD��<L%��x� �;܈\Iph[���$�Px��2㕟0��uH�fV�?]�	���.l�^�GL�4���[b�s��ݩ�'m�=�d�����Hs`C�k��C�Nσ*�I�5���t�6��r�[�0<����.���"‽�r�9ԯ�8,��p���ɬO�Adh�I��?9�e�ƻn�j`�%��k*��ghί,vn��
ϓ+���c0O�m� Y�~����H�)�:�Y����?�u����O�'(ȭ[ԇ�-s�XN�
؋"�Eh]�I�%CS�)Рej��O,�MF�jP�Q�'�2��⏯QrdyD��)P{���f�D��$F�C܈��	./�N�韏P�bE;������T�)��J3s�vQZ�i�0fl��I� �2z�d��a�.�<����U���Hǀ�Ij��y7Θ�Uaܠ4�8!��.O;���s�y�����B*D��`�%'Zehh["&nL剼(ݔ`�����GAV���AM��`��d1<O� �EE�8�~�@�2_�����7*0���]�a|R�I D'���K��=�4���M�4Zl̢��L?4�6�����wB����fkW��˓AU��	e�L4� �k�O�)�,1�`�&�LT��ڹl�L x���&Ӿ�1����+PnI��DO쪈W� ?���X*��y`S]��`a	���'��+DM\�-��h���d%�H��"N�TĄ�F☖ k\�JRJ�$�0<ɡހO���L�6w�}�؝\Z��y��ݻ�M�; ��4�CE�6��]�	4B֜}���BvMR �ɇay�A!`�'�vLP$�u}���(ܾ�*#�@�BM��]�J� ����ۊr"���&�O�䩈�ܴi�˧KQr�z��=$��{ӫ��9�~��?�3��/|�#�7�Ώ}�u��+�46Ա��mHVyҁK�S�ERÖ|��	��J��M	�)ԇS���:����e*�@�/���H��	.k�TA
���v"^��-E�c���=m��x����FA����_Kظ��E	yјh[�d4J�n��d��~xŀ�G�d�8e3� I�/��z�*�Y9J�U�p����Vb0���S$ F���a-D�P�V�E�<=�h�Ԏ�d��:��)�I8wF���T�π �  !��k@
��'�$U�"O�ٓ�HO�g�����V��`�Ĩ�I��&�`���<����HM^�'��6�(tz��~�<Ʌ�14fb�z��Yv�NY2�FC�\�>Ag.��w�a}R���z�BA��i��:�6D9u@��p='�^�M�N�O0���0�F�����~�" �"O���ԧhi�و�}�~�'����đs,8�'G䥻 O�~�R�C�I�O.����$����8p1���/v����4Gҩ��'��#}�'҄Ȱ�k��U�rm�w�G,H7hQ��'l�%���Q��!Plڣ=�D��	�'b�`UL�J���<%Z�y��'(�iz��Z����P IIE��')��čWI��
���K�F=�
�'��&�[%`�DЎʠD�m:�'5`!Sse_�dE���W$C� ��'*�a+�
�y=��9/�R	�%"�'�𹠤��5:�8���� J�J�	�'$��O�D:��g�8G��R
�'�V�3�Ξ5M���SdfN�u҂8
�'�9H�'M�hp�!l/��'�.�k2�R#W=>1�p��$ P{	�'X,�1�*p<(��0)��u��'O\��[�{�^`	�`�3+a�1�'K�8�7�]�Zx  ��GW.��u��'� Ԁ�ɬR��S�l��)� ���'���� �#C���q�e�l�r@��'j��*�"�~P�pC��Юc�b���'�R!ӡ�#B�:�"�W+�Y�'; �� clPC2��/<��	�'(�)(�S7)�N(#�/[�"`4�	�'I9�w����t���މ¬�)
�'~ڰXr�F�=���iF�iZ=p�'��`{�ڢM�tؓ0A�: @Ą�'/8��"�mN�٢0�v
�Y�'̢��K�M� ��C+��p�@݂�'�PR#���M�dpS#b�o>����'����CƄ)�}�q��dO�͓�'�|`am[6x �h�	J�T���'fyXA�N�<`0������'b@U���<m�����aGr4C�'�w��W>�`���
Y��hP�'}��	�NB6�Գ�O<�����'���X�G yp:�㥫ȫI�bl��'xb5���z�>)�QJ�:D�%�'�"�q����D�r���
+*L�
�'f���N��	�<Ԛ�HR57i~��	�'��]� N�v��t��3�
Qk	�'�z�iՠQ���@4b�w] ��'! ɢ�P! cD�Wm��0
�'�b�`��܆M=ȸ1��Ϡ[X:�
�'�f�HDE3`�4�9��݇[�pt�
�'�"��O,�<3�m�"+p���'��	 ��A�Z:eĎ�'��P8�'�Z,�Ԧ˰R�z3�"����0�'�<q�!�8��c��
��P�'����4��#�XP��"ȱ6�`�'�l���`��p��ߞ,a4-	�'h�|:��a̜�7	G9.����'�dq��:oھ`cwi�!d9��'�
5�`M�3��Yb"�& y�D��':-
���)lD-��i�	�.��'��,���A��H`Q)D���<j�'�a���-RA��0��ѩY�0���� �����]!t�2�h�b������"O� ��Lj�eP�B ����A"Op1ʴmW
~p7�W�`��q�"O@� ��>ީH#��R��x!�"O���և#�%U������+�!�dG�*8�Q!៖�<\��LO�E�!�$G�z��H"�^�8t�"�ڥ�!�Ė1UsJЛ2.[j�(�%B	�!�Ȯ�>��m��������>w!���Dt�!�j�v� )� �Z�!�d��Ag$�
�Ɵi���G(I�$�!�H\y�`��*SL�thC�ǿ?�!��	-����jY�*T�#冝j!��A(�6$8��[4���k� Q!�D�n�H��pJ�O�K&`	|:!�DZ	 ED����Y���ᗄ
-�!�"/p2}��Y��M��B��!��,-�d��N%%��ѧ�U�R�!���M�i�����(�n�(#�Яcn!�$�-t-��q��Ƕ��@�҅�!�$ŧU-���₯K��)�n��!�$B�}�"|c% [i�d�7΅>E�!�P7�t�AM�'j����j�;*�!�d́=��8#$n��ib`@�����!�N5H����dE�l������!��<�@����#�� �
/�!���'
����q�@�1��IK!�D�#��X4�S��t���.�h6!��&��� (د=��QN^,!�ʛ7���"��W9��lA��@�!��m�(\#��	��cћ�!�����[��4�`r� "M�!�H�@���
Yaޝ��+�;���8�'�zm�1��345���'	b�s�'K�eQQ�:)�ʨZ�"J�|=�Q0�'2n�1II#ibR��Q���u��y�'�j�sE��iٌա�Ǌd1(��'L$1 4��N�21i!,R+X는0�'j` C &_;#y�̆�g�x�ȓ_^u#B�N?6��u"�4^�ܼ�ȓ0�M!�nPd�c�a���B��ȓSؙZ��׺H}~-i��
^��ȓ#�����`2q��/� 	��ȓS����Y+N8�[glN=97�5�ȓj�������90nuS1m@��U�ȓH��B��*>�QK�J�A���� �pY�IЦ]��y�ƱݸX�ȓ�.������U2���,=�X���#�TXb,��ʱ��C_2u�����$���3�`@�O� p�I˯!��+���;�#�KW�=
�D�wD���ȓX!(����W���%��B�	���.��A��%��(�<�rԤ�/I<Ņȓ�ԡ�"4Y\�B"�9 �а��7"V�b��;<�ڕ��y?$x�ȓ!��1�SE��<�ع�e�'����� �",��oQ3Md��	`I,K�d�ȓ,2	��&��z}�����#8J���KA�I��D�X��ѱ�#�[V��ȓ|Ⱥ��D�ȜÄ,"�Z(p�-��s����G�\�|���{A�<܀=Fxb�;�S����L�С�1dMg���i�6�y"�ɡzj����e	�^!jyB���y�e�0��IvkN�R{(dje��y
� ��zĖ��6���H�%�,��"O�;pCH#8�]��͟�3�|�Pb"O,3Pb��@�d�(sBފ�£"O��˕���Ogt�p�A�+�$��C"O���
�#~J}s���=�d �"OH9�c�R@rabG_����q"O � �p�#��!e�l�+"OpL*@���4��K�݇;��"O���P���_�Yȣl܂  *`�"O��{!D��>Ay�낐���W"O��ڐ�P�+E��J�� 'd2��s"Oΰ����)'D@E�mF3Gh4��"O�<@���}�0�T��!$AV�Y�"O���7ǋ9a�z��L�m� U	"OބIw� 8g�]H��Q�Mip@�"O�����E�2�5	�ŏ�L�ѹ6"Oj��gIU�u?��j% �(=^�%"O��Um$���c��xd�'"O��*���.v&d�/1k�)rrƞ�y2%F+{��tJ �T!gЉ� ��y�HͯJ�U*խ	�f��SCٕ�y�I�4;`�b�.
(ɜ�C�=�y��(�*U�	��veÖ�y�lE���!����U�M��-'�y��ھp�Ve�֫Q�}xhbgAϾ�y2�X�Q�\ܐ��ˎ���[�f���y2/�>',h�C���GФ�dQ�ybNڦp����=|*X�Yv'��yrOW�v��ثBC�B��	SI��yrf�D@.�;�:5+q�-�yr��[xb�;"���#��<4iR��yBE��my�}iK��tD3�y�W�}⬈+$�t��yB��JF�Q��ӶUz�2⋍�y2�ҡ���G�zKb�J`��y"��bE`�Ǣ��!:hq���y�eݻ[����rU�������y"�!q	� 1o�g���G̎�yD�0ö�[ �S�H�H���"Y�y�l��j��d@��2xl��W��y�	V/1$)�kףC�Z�Y�E1�y�+[X�X�q0��38�E�%�M��y"͞/%N����-��E�[�yRԹH�b�H� ݞB��؍�y���L+��⠩TS mz��[7�y��'��1 ��$�B��^��yb+¸$$�Õ�a�D+�I�5�y�����եS���X�*Ģ�yB��
�!�N�(R��	Xm�&�y"`�9� IW+��I�M� ��yB�Q�`X����X�������y��Ɍ��Q",��ڜ�\8�yҠK}�Z�$Δ�U���raO��y��X2L���Aϓ�a��JR��=�y�(G�H��sH��|���A@�&�yB�I(OC�#䆉z f�mI��y���|є��TM	a�V���	��y�/ԇ[8���gbږe��i`g���y�&�d2
�ҥ��]z�uk�č��y�˗:!�$�Q�`�'��7���y��3&�=0f�˘LJpcq�E/�yK:z1�Q�!��j��mi��y��JO4$Q�6�D�a�dxsP�^��yr�\3[e�0�Ղ��`o�9�2���y
� �o���X��ʏ$:!�\�0"On�RCL˶E���X���?&X��"OhTr'.T�i��A)S�ֺu��9X2"O8ã�P13}����W�w��3"O��Y! �Fo�)X���R�0�R"O���3��>S���B�
}@�l�#"O���c��1R �;Ё�)�r�a'"O��c����Z6�xr��0�(Qc"O^D�EC5l<r�z $D6�����"O�R�?�Ԙ	�a<NP�	�"O��� �3 ΐYչqFtT��f(D��*f�̷!���:T��S�p@8W)%D��Id�	+��ze�Q�f�f\�p	"D���$�B|l2�j�DF挈��G?D��Б%�tHdy`���wXb��u@*D�DQ�N�+,<0�'��:g�d%"�&D� �U�Ԓt�dq����_�"�Q�� D�0�
�2ަ�d�K�Z7H|��g+D�����0tZ�4���n2��)f�>D�xp�D�>C�Z̈ �6Xx�Zч;D��9эQ>Ue�1��f 3�^��4D�h���<7�� ��i�Tw$���3D��sd��q�h�Y$���!��/D��C��6k&��a�#��u  �	/D�Xb!S�3��4T#�W��2��-D��x�J�9;)nt��	3Uc��u-,D���'��+�H� !&�;v˒q���7D������2Y�t���ŗ�4x��7D�Ċ�OD��؁�m ��s1D������U�*U:gfX�U��p���0D������]��׻<V����9D��GmM� `��x É/�Zu�n6D�dQ���.�(�+���rB���4D��j�&��<��Bީ-@m+�(?D��{��B�8��*^_�Y`	 D�2���'�L�A���Ot�t�+D������P�ۖm��w>M��7D��0&$:_�x1���)��x@�1D��wNG2u���2#.ؐR��X��#4D��3 G�+l¢]RvF��d�TG3D�jP��o��q�̙L����G�;D�T��)�	6/��bvc� i��!�E�&D��I��U$51tbؖ*���Be9D��k�Kج[�r����<8�p��J8D�8�)�2����GS3K\�31�5D�|�F�,�Ī2�F�xHT�F�(D�x;����a�	y�tХ�;D���fU�s3,�b�0�q9D� J����N�L�� B�*�V��Q�8D�(j��+�́ѐeC/@:8b` 9D�LN�2���eΝ}p�0�8D�PX�lB�ubƽ�C�L��Uya� D��$��vͪPX#�Z�@���$�?D�8ŇY�QU|��cD��LSV���� D�0q��+�J����<s4`�1"=D��s#2 c�p�f��L�f�1�K:D��e,�J�NTx�S*pDR�Q�:D���/�4C)�X�R%O'W+$$�U(-D������-�� 	U��0)��E�*D����,�<!�̑�GB�tð��A	%D�p!����� 䊴�D�@׬��4&/D�h�V�j)f-�^��`�FE0x!�$��:K��RUnοF��1רMx!�d�-3/|X�0����)ʕh�8Z!�� ��YҨ���Dj�3L����"O�}�q�Y d� ���O�F����"O�c�
�TP¬�i��^�|�!�"O0|�%��@~���
-x}``c�"O���R��u��)�#�ߑ"Sj�5"O,�i��>}���Pf� P2��7"O� �1�ل1آ�2���%�| ""O�I3ჹa��8��,�E4<��"O�Q�1��$�x�hb)55�yA"O������]�rX#`iȔe��£"O��#r�5lQ��F�S�r�C"O��Xd�o�ղ�oW�PD( �"OJ5�ᩈ�Z�!��~@6e1�"O^ ᧪�!\����'��V�tѣ"Oʹ����*Q,}��^�)+���"Ox����Vy�4E��L'" ���"O2Y�DOà]���@$@�Gv� 2�"O6Eq��	(z�i҅R>�(�	�"OB�RF��.550m�����q�p"OPD��F�X�`���� �&��"O��)cBG~������:|�"O��@�I���}�oV�@���"O�ܰR_�Wľq��M׬&7|Ɂ"OB�ђ��+>�e��nW�3��pBs�'��OaH A�?��\�㓘-|��`�"O��:E��c=�6Aͱd��a"O2� ���Ba]Q��"7#*a!�B����u��-"����AZ�dz!�d�U���wf��,a����[9P_!�D3\AT�����M�٣�ԡ�!�d	�:���$�� `�Dc3^{!��ܔ�P�CI�-F�J�����7ebO�#d�����X���s,�0"O�Y3��U�q�|��'��bSX�r�"O��.L�0"0�7N�P���2�g>�pa��(cG&$����# J�\Xw�/D�����"��	g�(5t���V�)D�,��b�A� $�� ���N)D� Q��|`��H@��UA��<9
�5���#�#A$��/i�٩�2D���`��Aq��KEM۝F��.~�!�X(��ɹ"�ɹ�v@�&&D� �!�D]1v��i���4�V�	�c��q�!�$Ɗ,:x�id'J�W����ȋ,B!򤒫.`���	W��@���>�!��K%l�Ȑ��Z�}|��ɰ�S�~�!�D\X���D�
S[Z��ڦo@!�d�%%D6��#�I#/`֐;��;#!�ɘ��p�M)GU�X��)�/1�!�DK�n�T��`��'_㐐��Òb:!���!��qk${̀�1mX�7!�Dy�����@	[��)�L�!�[:x��+�}���cR��!�R$�fY!�`�� ���l�)g�!�Z-H=�#�=ގ�bA)�OA!���o=^%����X[�ɣ�!�Ć3)dVM{sFC. 0���u&!�2}0�Q-�%o���:!OOxk��,��7E�P�R	a�= ` �*���4ʓ\Ș�V�J�X�,�3)ٵ%$★ȓ!��9�T��{M�c��3/�����R�9�P7h�X1�f�P-Di�l��`���k�Y7pX�b�X�8���Ey��'��[��2X@%Je㚇CѾi��� 쬰�L?+��fVk�J`a�"O�`�`�<��|b+Y*2�>�R@"O��XդK��,�kB�]���3V"OZ��Ug��;�TH�S	�	𒝂�"O��a�@.F�![iY��~xP�"O��]�PXt����:τ���"Orp�D�Lf-P�(���B�<��"O��CR���+;t���	՞@d,-���'B�O@�Z�@QR{��z4�@A��""OЭ;D��9Ȅ���Ŕ�U4ݱ��O�6�&�S�O�H����01�gET9�r���.D�d�V��6}�0h��Q�A�`t��H,D��I�Z�\u�c��Yw2h�$D���t�ہW�, �2H� 8��>D���W�*g���	�
�w���jt"<ғ�p<�3�RІ�vg̮+��Pٕ
�t�<��l:R���R%�����C�ʜk�<�lO�<4�0�& �/�YC�gj�<���o����`�pN��0���\�<QT D�&�L�d�1�I���\\�<.F�|H,c��fG�,�b*FW�<wOC]�1t@�=�R�7C�Q�<�c����q�۷-	�5j��t�<�ƭΥ|x���@��Z483hn�<I�튻9��xAB��3��1	���i�<��%D-k'2��'0<�,��U�h�<���ͻc�+�G�+���"@�h�<��ElD�B��!$�y�n�c���>	'`�,H��9Y`-�4f Ԓ�N�^�<�eB��6�"�M�0wZjA��`�X�<� �	e�|Зe_�_ܠ��0-�P�<AG
r�X�bCE�Nw����)�P�<a�g"]Q�H-�v���ŇV�<9���wh�<Y�A0COO\X�B䉕 <\`�%)��JC°B�	\�B�ɢ;U���DM  ��a�GҚG�C�	9^�DA�	H� T��AKĒcG�C䉴x���kqf�Z�	ՄÄ[�ZC��:�* unZ2l�T��׋@;� C�	a׊4�vI�h8љ�)�n
C��	� �p'?%�iɲ@Z<B�I�R��`b��-J��z����dC�	-IƝ����?a|%��Hݵ] B��E�عq�͵[�n��	�0Q��C�,V���cMҚ� �҈Mc�C䉪g�!C���u3��d�JB䉿v�Pc(�<9i`�� -�8�<��p?���
;�\���$]}�� �G�K�<� ϛ����0�hJY�됤BE�<��>~e%��Q�Y�x��O��qD{���i(M�b�2THjXȰᆙ5���@�'�n�W��.G���gϑv�N���'�vh#â$߄l�����f��! 
�'����j	%{��`h3�f,)	�'����d�w^��KR��-[+$Qr�'2>X�"i��y�zj���xE��'��e!b��,!����':Ma�O���ĝ9n��$:a�-w�������~bP�p0��w���D�_�7b�@�;D�xBPj�:xప��ݒe���A�?D�x+��V�[<b�(Y�&��!�>D�`�)��
Ԫ�c�d�Hж�4��[�4q�
O�+�\��bH�5%b`��fȬ�P��`�4ي"�'2	^���S�? �� � �*RN�U*��w��$�3"OP��UJ�8B}�IH��Y'#�	$"O����J�
��ْe�#|�1b"OXqc��<{� �^q��u���F�<WG�JRW�.QSL�1���x!�D^(��"��^�*d|m#BC�B�!�ӎ^��x�#Y(%�P zըAK�!�Dȓ���C��
=������J1!��
�4ja�BĸyQ&ТV5!�d��:��t���ȡ+�r�+R��"%!�X	c\���ē� ՒD��9!򄚷3�Ҙ�7�в�>ṅ��%1!��5t��ÂO����=b&�(B,!��v�L] �&�<G~h�QH��<7!��%wf���a��z����:!�W����2��6xJ�����>p!��G�.�M��(��}:�)q�ޘ"
!�;fud�F�����6��t!���t��d	��vd�PX�+�!�$ΰV\L����٠v98�t��	�!�Ă �2�iR���#4y�ԇ�4&!�d�%=��A��I�= HŬA�K�!�$_�u��B��$=�)RB�n�!򤌈m��k��ĄR1 �Z�`�!�DS�TE	7ř8�@�J@%�!�DB�8�zd���6&0	����!��i;@�P�W��Ta���P�E~!򤎸i�l�2�˅t������+B_!�d���0e.��%�,��S�+�!�D�r��l���(���r��(>F!���D�P��䊅�liea�ˊ�]!�p�~�� $č3V��h�J�!�P�Fʎ�G�E mBԝ��Hɳ!�\�Y���Pj�*R(�H�V���!�$��5�<5C7���.x�E����!򤃁9��L �BҰ%��<[`�B�=�!�$�f�����gt��@��l�!�D�b�q��.L�sv�C�;�!�D�-o�DZ�X-4����K�*�!��آ��@3��&[�pԣ"��7a!!�7�9�%�=qT���j�]!��+#��l1D�Y��K�j�!h!�D�.Of����4<c`a�7'��R�!�DF�V�*�XU!ɀ~Y��B���S�!��(WnP)�
F�K�`��"�O�!��IjT�e���*'T��s�D�h�!��w0ƥ[� \�cF�<R�!��� \{A딏�(e�𒯂�1�!�$�$Dj@Lbu�
*y-��vO��!�L�F�~����!'�H���2�!�^�|>�S�[lEb��h�o�!��'tF��0M�N�'垙l�!��0��]�f▬0�b݊�"æ�!�"x�GɎ�bH{Ћ�v��u��?���D�/ c�|:����k�\ŇȓxY�lB�I�:hx�����?�
�ȓ,�dz��:V�~�sŋ�U�H�ȓq(n�)��C�M_�{ӣ�l,�y��B��u���Q;'�P8��	;>I6���T̤2A��m�Zؚ��H�/�؅�`����VGX |#Z��f�R$K^���ȓT'�e�h�	����" �]"R!�ȓ���I�y��ԫ��R2�d���eg��Hf$F�Mؐ ����.76���S�? F���#=�(�ҊߔD^���"O�i�PEއ �6��U�@�K�j\�"O4))d�?P��i��#��S� \�E"O�|��ʋ/T�$�S6�Z�S�l�P6"O´�q�B�Gx0����Q��)j"O�ke������X��"�h@s"O%AM�Q��)s�kߤv0 %��"O��B�$�����S�i�6�n�;"O`�P�Dʷy~l|�6o�AFuz"O",���W^�m�A�-$���"OX���˜:��X�&T�h���!"O,E8�N#Dx����Hj&"OZPqG�i,ՠ�A\3Q�M!�"O`�9�TA�@�/S3-#�@�Q"O��A��S��[R�P�t�E"O�DK"��2T��#ć�Q�ލ��"O�q�T.U/ "x�['��"�C�"ON���I
�)P�8IG�ӫv*e;"O6QCd��:��9�p�=�3#"O�M���κg�,q�"+��0�""O�X�e�N�|�^\�3��4
�x�6"OR�3����r.���
�=ސ8�%"O&��p�E6D3L4�Ϟ�!*���"OB5[$�T)Ê�%^�	z$Q"OZ��C�:��g�ݽ-�1�D"O�`�F�
 f�D��i�<R�>�*�"O~�#G�@��r<vi�@�"O~`U��5����g���L�B��s"O��(�W6\P.��C� )��3A"O�Yj���H:t�7��^���!"O,y����v>�U˲ņ)E�h @�"O�� b@ήk� CC&�?{n<��"Oj�o�0n8D�kC� ft~!�"Ot��r@ӎ;>����w��!A4"O��ca×�'o�}�E-G�i�����"Od 3DO��Xag��v��A"O<ݛ���4L���{R�B����т"O�`�L�9V��K�kэu��	"O&m�� � ��0K�Ĵ">H�*"Ox�E� 2y��]�6dUb��9"O��F��IC�@�D]�v\
4"O�X9��'�(e��6HG��a�"O 20b]�74��a�eP�f��aSC"O88R '�!^��h󂀞�tT!s"O@���/�3. JѪ�"ř~$I�"OB�S�D)�2-���]7s%C@"O(����ׁ���䈅�OP�]�c"O��Ȁ|n��Ѧ�K;��"OD�Pd*cgF�Ps�ܴY7�t�"O�m��hA�ՈBf�
0�i�"O�X镰}e���^6H)<��s"O�\�U��ju ,l0�� "O��Aa	�� "r�pVc�G�H�"O���AA$���C≰Q�:U8�"O֌y�`�*HE���Q��>'>,Ujs"OJ� ��	"��9�JT8,�@�"O$-���Z��Y�U��x���"ON��ܢ@l��I7Ts�E��"O�1�(��mQ�	����`,�ٴ"OxU !G�(�`���	4<[�("O|�Y�Ӝ6
��K���6-H��u"OHIQ��$���B���.4t칐�"Op�R��D�R.����dHMiU"O����ߊV��رġY�9<��"O� �$ЇOņ��|� *�i�V"O\ţ�9��x��B8C/��q"O�����$ܼ�!�I�%]'��6"O����C
�j̑	Ɖ��'���"O6a�`�1O��#�S?W�8#"O,d����2���i2��*P3.(k%"O<��dƽ2�0�3� _+t�5"O��b�O�[ھx��A�n�d���"O�@⡋I���)�� �U$d��"ODdg+W:Sh�� �fS6�s�"OH��e�B+a��x��d�!E�,��"O	9�e�-@,-H�\�$�\�"O�\k�.����SN�;l @��"On\9W
��B�B卟XY� yU"O�=J�(��*v�(�L�v�F.�!���(a��*��%�N,yR�^�c3!��E 3�J��'N8lV���'5!�] YO1��L��	v�B�e��X!��_��\pK����W8К�M0%�!�@=��R�K�kA@A���?�!���WIh$�2�[,q)�d
�c^g�!�d��w�dmP�W��`�C�(P{!�Ĕ
$$Ne��O��^��h��G)Z`!��I,.��4����ը�Ӷ�!򄋞@<zu���¡ ��"�&�c�!�D�]���P�\�F}z�kf�W4~!򤉊i�@���%Ӑ8�'l�x!�dT.8&�-�"�o	5)ڿn!�͒V�0��B�^H|�C�\]�!�;F�$���±U��X�c� �!��[*u>�a1eCF��� C�!�ӗD��A�����$�R+O",�!�d6��t�ΕX����$���4j!��CH1^�ɶ*�,<��<r ��y2!�G5O���B7�Î4v^�P�ⓗN!�dr��q�q��[\��4��f�!��bV,���̥z7�
4�Ʌ�!��S�m�zuRѥ�N�P��@�[�!�d��Hr����L�v��)T!���&+� ���/f  ���QG!�P&#{��	��6t��Y8`F��g�!�D���Sug8Wƒ�J�ʍ�!���=��t8Ǣ�T*E+"`�z!�D�%�����z;�H�N:U!��Y/\qZ�#A+�'Q8ҍ��^:�!�K�d�NW��q&�L37�!�Ҙ$��p�3eń�ܨہ��kl!���?@��EigZ��m�1�F M!�z���Y�&6�Р3�	�'H!�˟QM6'/V�-����c��Q�<)4ǝ3Lm�\$I4�)���J�<	V�0i�z@	q�+(.^9��&k�<���i:��#n�*1DX[1�i�<Y���<4$�BUoޣ#Jb��c�Dh�<�FA,G���H���2�|�7�@e�<IT��4JHtu$�7(LY�v��z�<��ʄ08E�S!k�2�րBcl`�<���F�z?8X�3Dӣ5��`�H]�<�%�47]~\{ơ��P|pIs��d�<P��j��^V:eȣ)_k�<a�g�I*� �O>����F��j�<���_�-�·�كY��:f�RN�<����/4�dУ��Sppd�vbv�<��F��/�IT�Ǌ.5"d�[n�<� �9`U�*�}r��Vu\Xv"O>uv���8�I�&�������"O�I�f�#FDj��j��2a"O"8H��#Y��Y��W�8��)2"O����"C�d��(J9D٪	J�"O���dm�R
�Q�Pg�k�`��"O�p��KF��"4��;��D@C"OxU@�nî8r��EK!||ܭl<D�� $��-y<�R���4o��-k�)D�l���HDT�Р�S9^����P�*D��S@�i��̑1��BO�4�@5D�0 ��љ �.��ҋ2!5(C�IR��� ��.�0�n¨T.B�I.|M���#��a��Ȱ�n�9U�*B�'}{�L���7��Dk�Ǆa�B�I�oD~�S�K� LP�lyn�:��B�a��T #���OdR쁐�W�m�|B�;8��A)wkU4}zJ*��փ�FB��"\�R�2�ퟩRX|ppkY�YTC�	���(R j\�hKHl)bC2�8C�	_\ �j���X��a!Ԩ�2C�	�b b8��2�0!φ�'�(C�	��C���i��(Y��GC�I�f�pabR&X����˭�B�I �~�b��h�$��IJ"H�B�T����G�"���CFʹ+ѼB�ɲ����bf ,s|��[��G��C�Ies�����bŪ� ����fB�	�#���$@�9$&bH�)��d�B�	�7{�1���
=�>09A�(hU�C�If�A)7�-h( �R��&Q2�C�,�
�J1�]	t�>Ydk48G2B�ɼz�9��]�(
�L�C��hR.�6�]�QI��80��"��C�I4{�����ϥe0�y��	�F�C�!��ԉclW��,��j�>9h�B��<od��ӁJ"�ȕI�ݟ1�<B�I%W:����f%��s��Z�h��C�>��h)wG�k�ޡ��䙧D�C�ɗcy�ˡO��u���9B�V�4�B��=	�ْ��Ǣ7֥�6�U3|��C�	���I�A��d$ԡ�ć�n!�C�u@F�:S	��Ny����ĕ���C䉨]
!QkK!'���sf%��:�xC�7�t�a6�2i2̱�T)S�b�DC�I-D�RY��MJ�Y��"A�C�ɤ"��p1͗�Y|�ؕ,�e(�B�	3y`)����":JX���Ã'+�B�I�N!���"N�/
�<���e�C䉕J��,�G�"��89�)@cX&C��+-��2RdΑ�z$	fH6(S<B�I5HĤX"V���}�L@(��[9��C�ɴx=*�ʷ���'Rt!�0#a'�C�	�B�>\:��æn�~��@iϥxF�C��7`�et��=,�l�Y`���p��B�&>_�r���?7�\��
�	��B�ɸ(���p �;G�R�w�җ5��B�I6 ���@��V��T8T�V�U��B�&#8�����5I�$�b%!o��B�I6'� ,j⌀!B׆0�-����B�hT}hP�jE�[a�P��`_��y�I)��J�A����m�� N!�D��N{�i֌�|��B��&�!��M;���#Uj�Q�ӣ.�.N�!�� Vڔ)ʈ��Up�L�����S"O� �w нa�lY�i�����"O��7(��>�>u
Ձ�T�����"O�80�	�Vz� ��|�Z�R"O�`g+�>q:��#5�9
�bL�"O�(�-�mB�0�	��:,ؠ"Oi��,K�Y˧���/*Lq��"O��p���v�@�BC�Q9,i�"Ox�-y�D)��b�0�b�$	@��y��'+�-#�S�j����N=�y�&�']��)i�GG+bvR��R�Z%�yB�כn�$ �i�i�T���,�y�ʉ�sst��2�F�,K*�ʡ���y����Y{8Y��1�@@1���yBB��Ge��	�
U�6zĢ�g?�yħ�<k��N�	=��R�l��yr�M#+�`-ZvQ�|���1Do���yR �,��W��5n)BDZ��[?�yR� ���J׌�V�dr0���yb�Ǻ{�lD`��L�D���o�y�ׂD��t��L�v�� 2W�I��y����Y��\�-�&G�pAs�4�y"@�+[H�[�O�&Q2a���
�y�G
<m��g	Q!$�b5r����y�Ɖ�b��t)�k�/��S���y"��S��ma�D
-ؘ�v���y�jL�ƄX��(ɞ�@h'��y�O,xR|�ФR�I֜i ���y2��8q����M,�B������y"���/�Fh�F	ʊ�4��e��y��&/�!��b�U��=�yr���^��84�	�9d�`e��?�yr��76t��cFʨL���+���y�iV�F�yq�'W�p��+�k̿�y�g\%h��e�	�p����Y��yrM�4I�e��ŜU��xв���y"OԇW��	�a�6N��4��C��yB�K
C1���Q�B���`�ʥ�y��� ��dZ	�.&0�bd�y���<�(�3�Ĕ��b@z&���y��J�|�p�5�Άy P��T�Ѣ�yr쐏O�v�x�I�n;
a��ޮ�y"J	0ِyi�-R$N���G��yBF?���B_�N d��B��y��[���ĉ�D�Ȩ�7���y�#f{ba����4�f%�-*�y�a�4#����8	���x�%F2�y�+�\:Ġ�69(��%���y§ �����Ʌ`<d��Ta��yD�.]��0��*E=�)Z�J��yBIѲhs�+v�\+	���U<�yrm��L��o��3���5W��y�K$hst@ ��U+��m�s	@�yA!�z!j5�M���y�(�>�y2
� �N��e
K.D��9�%EE)�y�c�T��ۤ�صC��Q���!�y�+ɌKo@	�cA�
0nh��հ�yRI
�p�NL{k,e����y��'e�AK�@�}��!#4'	�y�c�9����� �L����_��yB�� "�,����s`Jt�H��yR�b�p����e�ƱzQe��y� 
�s�:2r畛\���s����y�"j0�tp��Nː`�VjV�y
� �0���\�@�'	�0/�}��"OFQXb��(�J pӊ�)��!b"O �ҡ��:�r2��	�F#c"O�(���L���i�m�ȝ��"O�	[�gT�<0��Ċ��8� p2s"OH)�w��u�]`ֆ�Ɩ��"O� �f�^/"�1eE�,�p�z�"O d��ǦR)��b%e��j�:8�T"O��g��hXX��I�P��J�"Oz�G[�{�=���U�)����'�T�9QJ�Le��#V� �{
�'���b�+���������9
�'m�����`8��Y�ŋ^��	�'�6H����K��Y�#�V#eT@}��'BL��C�oa�����K�O���' ��s��A�r��yd����p:�'ĦD)�/?p(�/���i�'��x�!�-;^D$Y�g�*
%|�`�'v�;��^�G/�h�KZ� \(U��')P��`l�0J��k � ����'z��B��1����!w>*!�'��Yzb�Ƴ3��,�/�gӸɳ�'��-��M�	���B�V�`��Ś�'bM����/W\P�֯H3Dx�Y��'�7MG	�YꂌE?@��b�'�T�kDN�wx8"n�;�p-�	�'����
�#+�"�_!`�.Y 	�'��-(t�0s��DG��_R��R�'x,�'� >1H�iV��Z;r]��'5�PX��ȫp6
ۖ��!&k��X�'�2`*-��}��A�����m*	�'RH;V��!����L�mvM��'��#�F
����C� �	k�Mx�'t�� ��d���(U/t�2�'j`=��i�L��@e"��y!0%x��n�q�
=H�!��y"�I8Yh
��N�j-��׉�=�y2��&[��kɄ%R�21�Šʱ�yB�� S� ��E�V|i%���yB�ś*�A��((�Q��.X��ybf �\b�n�Q�������y��p��@��΄47�Jĭ���y��)zuZ9��oV ,�cv*X?�y��@�@�"�SE�B�z¯ ��y�*�%]���Z�ArJٷ-:��ȓeW��0	�7Vv$ {c���*jX�ȓn4�eg�u��`XL�J����NR�<aGCچb�U����^U!��N�<1�K�K�t)�ˎ1�!B�KM�<�p��	qݜ�ҁ�
3�4��砌K�<��n�g�t��Ĉe�X���`��<��"���
��U
	���'f>D�0��f2qW�L�A%�t�J�Ƞ"*D����N�"<�o�M�(���'D�����7]R�!t�Q���dQv�(D���j̍�JL�̓�>�d8���#D�x��i��<` �'-� Q�F,�+?D�����,�R�����I�.dPl0D�@��NK�k$� ��<4��� ��+D���D��8{i�lQ!'�j������4D�Թ�"��I�3��}3x	�G.D��+�dFS%�ʖ��7)(�i�#*D� )'��&���j�Ծc�����l5D���g`@�7��X�Pѻ��"���y
� x(UhrQ�)�����?<� �r"O���(זT-b�vb�{ lx1"Ot��S�.�,��'�]�7�p�"Ovy���B��qC�L�#	�H""O`���FÅCU<Y�@�)fD��"O���Û�[��Q�sm[���h�"O֍3�Ȍ�m ��X��I)���c4"O����씃ӈ�Z\@�"O�Y�C��!GoF��B��Ym���"Ob�"7$C.��\�v"�rc����"Oz��B��3i�h�RdJ�I���h�"Ol#pN�mRDZ�c/��ۢ"O*͂�!��i���!	���V"O��I H�1h�	�D	,Q�zF"O�a���H�B(�:���o���"OfY"�G�"]\�sVHާ#��"O*�:R��(S�$QR��Y���"O\ƌ�.�z���Ě4g���	�"O��c�Bt���:G�WJ�έq�"O,=���8Mr�q�B�=HB0z""OR�z�A6~O�8�ab5w����R"O���Ŧ±\�r��ơ�>�H�`6D��� J��J5A姜(bŴ��d-)D��i�ӺN=~52U+v&v����(D���T43��P��Ԫ\
 Yr�$D�@� 7egx�{aO9"��� �$&D�đ�얚��jc$�$"�(��h#D��jU�00�@̚2ެH�%,ߑP�B�Ix�zX �e
y�� ��h��E��C�	� aF�ȱ��!r�D蒎X��C��) �R`:��'rs����ث=AnC�(6�V 0`6;E�<sSI���C�	8KA��Ӄ+�����&��C�ɚY;��:G�ۢPhI�o��1��C䉫&���#<�3G�HW7D�pz!O +Iz*}K�(�s{��k4 :D��2��VM�q+���m��tG#D����� ��x��)�bu��!� D��� I���E�W�(��u;fC4D���$vW6�X��Tn~a��m3D������r'Ơe�djR&0D������������٘WK4m6B-D��P�'8��TӄW.<�0���,D�K�-�3t!����0>i&�)D��K��-r\d�"䁛���k_�!�$0_��Q
��Gn�u	��o4!�$B�`;IRv&V��@m�f�Ǣ|,!�d�8P�\��A�"�l��B� m*!�� -b��pi��)Z�<B�b��+!��@Tg�9T$��\L�m� A�+ �!�䓏R�j���&y�L�0��w�!�d�5EY*�R���T�@`0 �]q�!�ΊG�ji��Łj�Cө�!��u6L�I�|Dmb+3�!���p�쨑�F�s,>!���u�!�D£8���"2(y0�kE3O�!�U&
�����[Yw�e� �-8{!�;y���
�A�}���za�8M<!��5�B\v�Z7�V�hP���3!�Ė�.r4��+��@�9R��
7�!�D�8D��A��t�f%xG%,�!��\�r�E�q~��:�&	�H�!�2*�!��+�R}NT3C@K6c!�D�/� ����5HŔ�I铹d!�� �q! P<t�LUb�*SU�6�I$"O�B�-"Op�i�Z����"O�r3e�>U�,�wH��%ߺ��"O�䩒�4sB>�2�B�9�rP*�"O�dXA��4�ыBe�4�j�0�"Oj=��c\/ș35/��d��t�!"O��㑣�j�V�B ��7��Ia"O�I���"'��H3a�T�G��1W"O@�k�B��@E�����H)v�x�G"O(y1qJĄS����$�^r�԰"O<�� �N p��ՠQDXq�i!"OƤ�$��5��碛��N�Q"O���Λq]�{u�čl�l�д"O8H�@�@�OK�q[s��j00��*On�3�E�(ON*�@�S�1�l�Z�'S�`����2IP�U�PMٝ%����'3�$�2�R�K�P�Z7ƵrV))
�'�ڐQ��-��i֏\)a�:�z	�'�ne� &�1m�� "7��.T�����'�"��&S)RrНBÏY�D[��	�'��IkBD�')n����k����'M�T3���:#
��2�͇�����'3�M9�"�h��Ex�)W!3@Ԑ�'��qd���^"��qd}��q�' 6��q�20hb� a��
�'�<�ቬ\L��hk��n�0�	�'�.�{f�ϝi���PQ@�/:]��	�'��@W#H	lE���7�V5�'�H���⌽P�$�fc>cb���'�����7:�q)J�V�z��
�'{r)���	!���3O��C��͐�'12��g�=Y�1�*��:�›	�'t�h�C�	q�0sb�����|�	�'� q8��_�O�ry㋽t�p��'��$�Ս�27��gL�2pq�<��'�aCF��dTt����@x����'�b%YD�D�BQ(�d8ld��'C��3�������$�`���j�'ڢ� ���Hd��RU��8T�5p�'�
�A"ǂ)��d�׈[TF�J�'�D�HA�Ȏ!ՒA���'�&Q���T���t�?6�.Ѹ�'�z���̛�0��tBP>5�"i�	�'���C�81` @S,F��-��'�����^�F <(���ٿ$�|���'�9�g�q�l�c!�:]��'��c"��A�U:Bl�"tE{�'A0ds��%pN�cPV��.i�'v��Xgg�+�����׾��!	�'^�y@ƒ�;*P �w͏>��$��'g>)k�gF�-�@#�jQA�As�'z$a�g^M=6 `�5t�'�fK��'	�9�P�'�8B
�'6�sD��/����(�-0���	�'
�q*caFS|�ْ���|h�	�'G�5&�S�^�Xv�D9!y ���'d���Q��c5lE;V��dm0m��'��ض��FE�|Ȇ	����'QJ�@�傦N1�#�Dܕx����'ZB��sK�6o��j �Y�X@�'zl0�Ui�qC��#MV9��1�'�H�R�Ň/�~�cϊ��X3�'�jʑ΄	W��9�˅���<��';ܠ���s�L�e�G8�&����� p�{�,M#�d1�HQ$TbҤ¶"OL\1a6f��2��:P�ݠ"Ox�1�ӕ+���F��I'.�8�"OZ<0ƇY�t~�sL֎=?d"O`u��7��r ���U&`m+"O0-��
F�4�\zp�%r�0J�"O��ׅ�(8�V�I��A �¸�5"O���s�G�+�~y��L����YR"OZ�i�+�<�V�����b�$�(�"O�	 e�B��6J�h���"O�X˶��M|�)��曅0b(�iP"OP��E� �d184��yظ�"O�I���ɰ�^�	��bV�"OzqiS�Ǽ]�iiR)�iB���`"O�Ȃ�ǣk8R(�Jh;Bq0�"O�u�C
$Q����iӑ\9$`�0"O��WH�<[���e�_T�b"O$��L�&b����PhM�=g�Xc!"O��gBARAS��߮hu�qru"O��;�K!D�2�#U��)c�$�B"O��[�@Zz��0����!9XD�%"O�8y�)J2�D-!C w��1+�y�;+X�7AX �`Hz��D��yB扁n�����H��X	�a���y�k��k��܀֤M���lC���1�y�.24ZDY�r��4;�5�g���y@�1��cj�)y\�&Lڴ�y"�0y�HI�Kp$��ʦ�y�,M{{������x��D�`I_.�y��2���b1��r����(���yR�L<>j9��U�h��dC����y����0�C�YdY��	��y	��E�����Kg���q�ձ�y�ɪk�b���c�A��$0�@Ū�y�o�/S� c%��3�*u#���!�yRȟ$�����$.4�����y"��%0p�ʻ!��37L���yR鎀$�I�TGI!>�e9f��y�N�Z���M0���kd�V�yrI_l���K��O��5�Ħ��y�)ǆ"���1����&��q�S��y2E�9�lu�a��
���RϨ�yBl_�7
�L�en�<J4<�����y2���g@��r�_&& �����;�yb=6p%Ytg� R����޷�y�)ܰ�t���ϰ[������yr�*R`C�m���.QC�L �y+�-f
m��$ψn 8��N�y�cI�}�^	2�+��k��Y����y��S�u�VQ�d^�W^�b��]�yb2.Z�"�$*C�n���/�y�MGE ^PH�Ե@\���t�·�y�n��i���"q�ݢ
���"��yRFZ�$�$���01����3R��y�G��%�R�Y�*o� 3bT��y���iu���Ŏ�$(�d����y�m�%8�	0���3���yRe�_��`�/%���6$�)�y�d�4$>��1��E9#��ш��yR	���=j�I�4:A���H��y�E��H�"mCċ��(��� &��y�a9.N�50Ldh�%`�!�y��"�tAT��]�\��&�yAC�s?|��%�/[Q�9��N��y
� $��Pe˥[��T�$ 1DRش!�"O4�ĤE!"#��Y���u9.�� "O@*AfN�M�t��қ�&`�@"O�Pc�I0i'T�s���a�]��"O�l�u�A*E	���̓!e���ʖ"O`I`����X����P�D*J�Tk6"O�%ZÓ=a�@��)��Z�~�#0"O�(:�����}�f*�i��]�v"OԐ년M���b�ֻ�bmj�"O�-qՀ}F�:rG��Z���"OQ��L���m�sE[3b}���$"O�e#��o�qSOi�NY�"O�} dn�m���qd-��q��"O>M��eJ(4��"u��*���"OD�`�;p��BO�Y�x�c"O���`����W�\�Wu2�"T"O�9���1�B��aA4Y�yڢ"Oj
Pƞ�y�-�&�h����"O����ޣv�fHbb��  ����"O����(�;|~�"� �{�6�a!"Ox�XcK&��q�� �/�v�a"ON�@f@'a�$�;�.��=��A�"OЌz�.�"I��8/�����g3D�|[7FJ7W���A�!��9"B 2D��+��C��!f���[M(S2D�x:&���Ko�XCLV�w���i/D����F��`��XQbiS5ּ!�:D�$P%��� �Z�k��ϕ ɜ)�2e9D��r�k@�;\�Qz4Ȏ?PPlM��#6D�����O��lwKl�a H�t�!�Ď&#"������[�� �̖)iS!�ʺ�HX3�ٹ@�>咂��^�!��'z|q!k�e�4�@���
n�!��D�}A�i8�懑l�ԍ��
�r�!���w9�5Z����ڰ1qG/�!���+&�-�hY�u�����xh!�$�ǎ�	v
���N-@��Kf!�D�lo�9�S�	&UH &h_${x!�ĈY{�-��J�EVh�;�&�)wC!�䒴aò�P�閏AN�m���,TX!��7[
���-L-+G�*��>u�!��C�n<ȵKu �`=n�
+��7�!��8|���ȉi���(I�b*!��_(����bO>#����g�.!�D[�bEr2Iֽ]��T'߃<�!��P���+ Α�[ݦ�`�5u�!�Ӄ3A�P1c���|�DFN�O7!��)
�j�&�>U��X(�
��!��O[��(SEI�ň��UJ�1�!�D��}�*%��̋?����CƉH!�VR��V��� �#.!�ԕFv
�� ��,u<]�`�z!�Dْ7#|@�3 �9�D!��l��~ !��I1�~���_�QKt���#�!��(�h�8�L�LB�@A)Ӱ:�!�$]��*��K��*Ln�@�\(L�!�D�B�Y���E�@7�urU�%E!��Գ/¢�)��I�$d$�&�g1!�M��t�F�G�Y�E)g%!��!X�z}�c�/"��# B_%!��c��Yb��3H�t�R0g�Y!�ċK��t�p.�Wu�Ęd�(�!��ƅ�L��,R=Y���G�O��!�	!A�^ Q��Y�<f1��fO�.a!��  �@��X|jA�!mYx��"O�H�-Pj�\��a�Yn�hI#"Or��g0dU���4GN^=��"O�4cP.F��`t���� C+�m#�"O�(�(�AS
�a�%͇t�$ *�"O�i9��9J�HU�p��l���&"O0�� ϒ�K@p��F��QQ�%�Q"Oq�� �<�T���]!�u��"O�@�n�2F=�Xa���98t�a�"OxQ�t��'V�~���� K0Z�D"O\a�+�&�4$��>FX��"O6��!��:W�9���7qa:1i�"O,QJ��#J�ꔋ�`ވo*2M�"O�0r���!0Sv��FEŏ6�Z�"O���B�_\�NZ`��%��r�"OF� �I�ar6� ��K0��	Y"O^tsa�Q����X5�ѭq���Q"O�H�#��x_���v��;�����"O>	�BU�[i���Bd��)�t"O @`����j�R]�f�2iƚ̐5"O��z�*��^��ј��9�l�F"OpT�G��tW��u%�?�
�%"O��[��&ʚ����V�\���"O�4�M9C� ��Ô�X�"O��e��d�J��ɒ>��E;�"Op%���ʐ-	d�(�,#�V��"O��B�΍A�(ڧ%ߓ	��p�"OP!�e�f)�'g�.Q�ڰ;5"O��ZU���B0ܙ��l�ho��p�"O��r�jE^'8J͗NW�I�"Oz�q�n�,)~��EY�QC��"OL� �`��^$Й��-�H!��4"O� R��njʐ�c���j(��"O|��a�2Dwx@�3$�#jE8�!�"Oz5Y�@�!H�$uHC��n"T0��"O؉zsl�(U�=:`
��$�2"OLm��$F�_Jd��S‎���t"O�=#TCΎiNvk�@S*4�xi`@"O�=SE���/dL;w��?� Å"O쌲�*K,�JY�`��T�6��f"O�$�5�I�O�z��t�Q�_v�Y	b"OP+�d;�8p3.�P����"O���	l�jM���٪����3"O�����A�q�r]��b��8s��[�"O,�[P)i8Z���
\Ur0"OU)^q��@z`L,!?v(�"O	���̸5%$�{�N�?V���w"O����'A(j.(���T;(`�U�G"O�E8C�'u��@�s�F�>��i��"O�L���mz(��e�)6����W"O����D�:#���S�)�%�!"OjY�r�����F$�
�6�c�"O
T2ѡ�>tq�2�ږvD:Y@%"O���5B�!a�^�`t��,P���`"Oj��G��s;z@ۆ/L�7�	�"OnQ�ǐ���mC,H]���b�"O�Y�f�q�t@��R�FNx��"Ov��3ȑ<<�h��`;V00q�"O8�vˣ��IȞ\�haH$"O�At�סY��3�MαFQD�1q"O����_%���el���uv"O"Ͱ'�<Hf���
2x�8a"O>�S�Ƅ�uGd%'̉NdH���"OXV�;W �BǄ���];F"O� d݉���A���&ۦ@r-��"Ofu��(P[�p���^6�p"�"O��	��]�W6qc��ۏp*� "O
��C��)vS2Lz��) �0�"O�X�U�>b�4#�!��"�n�1�"O�,[$��6	X��a�6�����"O��`�$Hg���ʩ)����E*O4 "V�t������Z�
5�0@�'\�Ii��˨=�H��-�1|�Hd��'j�B�#��r��J�_�<W10�'�4�! ř��8�+��.;��'��pF7%(n�ÀMP+;�y+�'������ �j�ǏH�-��'N �J��F��5 �JQ9i4�h�'_Py*���1���б3QV<:�'�%���S�*E�@k������'d��	bł8]�fiC��I0�H�	�'p��p�(g� �פ��$$s�'���f@\�b������G6��8�'�(��+
x�Zr�_+O�$Q8�'%����� �Ef�����¤Dg>a��'d���-MG>1�b-�:N
-y�'�2)k �R��Q�aa	� z�@�'���AP@�PC�Hs4�s���a	�':�+!�?on����ɚr��D�'���2gb/R�ꂤ�n1��
�'��В�"�=�p�W�¬2D��
�'l�ib��5ot�����]4��q�'OFmI�� �}�V�ِe�,R�p��'��eœF�D�" ꃏ ���"�'r��`f����R�I�P���Q
�'b����L��W-H�s��NJHT�
�'�&��K�:�Ґ��Sd�9
�'�����)ΔJ� C�6M����	�'���Kb	�w�ؑ;�/�o�v4��'k������ 'H�#Mx��Q�'���"�]?����b�Ɍ"�� �'�R�TM�9&Ӝ, 2�ϖ�6 �'|�@��՘c#��Y�`T$셙
�'x�-�i�Hl,�[5��
��8i�'ʠ�S�#�?63H]Ǝ��T6"O�}���)yb����(�H�6"O�Q��. ��+$J�Z���E"O�I�Ō��j/HA9�B�!%�,8�""O�PR#kI�k�Vc��)i"Ojd�åH1̾4Z��ԕN�(i;c"OdI���C?��:��L�u)�"O9q������|�F�I%4�^9�W"O�ੀ�ƻjG�d�pkQfӲ�"Oh0�񢊕rD@R(��e(�y��"O�$�Y$I�嚦G�3,9��"O�LH�k;m��QJ�c��|00X�"OD����������A0�n@�V"O��c�^'gPL�!R-�vH:�"O`	
��a�|�h��C��:�;F"Onȁ�P��� pD溵1�"Or<r���!�XX���ڙ{��J�"O�\:uJ�-c�28)��B{���"O�lҁ'UI*lT�I�P�伲�"O�8�S7yz(��g�"�*�T"Of`� �
(��(x�g!5�<;�"O����@%�$�����j�@�a5"O8�JQ�O��:D��M�v؂}S'"O$h�WdŐ_P����D���9[�"O� ��k��rf�)+1kB'M�Z���"Op9�����]��dK�ƔYQ"Olz���x��Pe��uyΔ;�"O (A0�Ӻh�@q�D��iq�
`"O>-	��֮@�\D#�I�\H�"O� �#f�?$tV�K�^9�,1 3"O"�dIG7r��U��ebE�#��Y�<�"�ļBpl���KA�JXR��Hp�<�qaâq�� D���,�8s�UR�<y��L�{�`hc7��0Hq�;���S�<��A��2���"�X��z&�L�<�F�f)��"��=�$���R�`C�ɻWP(0QvOwr��sO[c��C�ɆHd2%"S.MN���c�*��C��E$@��D�%b��1Al�ظC�	(W�^ȱ��_�#F��C0�¦�C�	;M{�Љsm�2Q�b�a���C��)�*��a(G�=�ܵ��O�8Js�B�I�;f�XA�JR�����0H\�D2�B�I��Ɲ�p$� y�i%ß�&��C䉋As�%㰋Z�d�t�è�Yb�C�Ƀ��Z�g�1!T� ��rfC�ɽOS�9�J[Qzh�AE�LC�+jȦ\	�l��*�Td@�e�.C�	Wndk"��ooZ8B�r��B�I�	yR!��)
g�>��f�� n�C�ɐ3�̣5E�A��x���
EϬB�I8i��1),?]�$t�� ���B�ɼ )�eТ�)h��)��߳/�JC�ob0@C@G�;����r�Ľh!��(.�8����S�Ճbm��#�!�ă�-���H�	X�R�A�`MN�,r!�dU�l턅�"BK�C������]]!�D�bt�e�b�_�-�4�	C�S	Q!�$ݠ2jRX�B �w�q9�˙a�!���"ă�Ñ�]v4�J&
�0X�!���-��ٓ�U*U]4�KU��79}!�d:�(����4^D�c�F�>P!�D�?5��[U�U\L��)�FǧR!�d��2 �0k4�O�P-�̓ƦQ�g!�"-��h�
�<p��$
d!�
x@�,S�,N,$�ˀ��(c!��[|��m}��U��beI!�$��*$��R�\ > ��g3!��S�2m���
�D!����m�!������Z{4��Cgdd�!�DI�~0"��T�֠@�Y��$�!�DβdL6���Î$jh�##ύ�!�[���"��������!��,s2��f�Y���m\�!�$�%j^�Ѵ�F
Lh�Q�,ގ)=!���|-x��
Rg��Ku�G�!�dC�HM�x! l�?jU�pjG��G�!���Pd|(٧���~Af}��2K�!�D	0�F��w���O'&mQ��>�!���k��L t"2��	p��.-�!�$t"]��c)�,���ɵL�!��{������^�R2�u�\��'5�0Bv����B� !�n�+�'�D	��#�l��0�T�߅�X�'xf���n�n|��6�Y�;�^�+�'���	!�=cݸ8AD��0w�=��'�`��	CJ%��!埐쪹*
�'��HPU
�)R�t%`7B�@D�1:��� �%�ϮK�����^%Pp�"O��"+�Q�e���:9J�(�"O����Fp	R��������2"Oh}jccT�Ktp	@0�@��R�"Oԑ�&J
)�>��V�
�X}���0"O2E��fD:J�������1ؘ�"O(8Q�/�!7<1��;�dHB"O�����B���ԔOcJePQ"O��{��&ά��B��\+����"O@15�� [�F��V9��"O�E5BY�z(je(��%��q:�"ORi��ǩH�(%��`+P�t��"O���ɀ?%�����^ �rY��"O��Ab�Ԃc�	8u�C��Y�A"O�<�Q	��1Ux�H��"l}:�"O.Y��B�PCh���L'=y�q8"O�����Pb*��R��un���d"Oޡ�s˛�QF���lWg&�R""O⅊#�M�~<��ܮ"f�xv"O��Z�
��%BNA3&)܅8B0��"O�<�!L�E�f��e'�8)՚`7"OvP��!�����f@�V޶	B�"O�����J�IX`Ido�!Z���	�"OD�FN�
ls3�Ά!|¸�"O>��Eg��o�����MØT�^�PS"Ot�ѧa�&�I�r���,Ȁ�J�"O��z+yf�ˉ�-���u"Ov�!坡u�ze�#
�k�"���"O�����6@̉W��1)����6"O��HT�
�N#D����*Nf�8�"O`���$J�_�&Ap7RB��"O��q�/M�{�ތh���M$.�y"OX��'��=��\"fkS��q�"Ox�ògH�Z��Y�
�-B@�A`�"O�T���\2@��c׎r(Z��"O,=�&mK��\�q �݂b"Z��"Of�{�n��e��E�R�K�� q�"Ohx��K�T�z�g�
�~�*}�1"O6�[􅒏=A@�a��ے���rv"O�+��x�Ƥ:��S�V����"O���7�6n��S�aZ�@x8��"O�H�F�H���:Gʏu���X�"O�Q�S����	 mk��R��Lg�<Q�I%e�U BNE�|̸��Zg�<����*EÆ�jG	ʵf�.a����b��L���� ��= r�|��XEa2�O�M��� )vg�|�Ő S�p_�Y��p�&�`�ͪ�bM`eg��C��H��IQ�'���ef��'BLQp��'o�	
�'M>hBdb̾_%�Ui���/i
����'��dđR.Z$���5`�R-A�'�P��'�ۉ�н0)�T�`�	�'-��'m�sV����	M/ag�q0�{��)���T�������"��yئ��
!�Dޱ��,1PJߣ)df�s�#T�!�$�S�����E�Y`���ׄ_ $�!�=8̀3�90~��g�R%���'D���i$��O������2(pP�gY-�i�"Or{S��b��"G���F5��D�
�(O�x��ژ��d���D}�d���h����xr$!r9�uh��Ο[F�%I��8PPb�4����<�E�Ȭ����k^�>��F��M�����i�,|*����tE;��-i�f��
�'lh��R��/-�� 8см\��!{����Ba�>� ���35�D��
^�9��M��"On c"oZPW�����i���q�9?a�)�'n�� ���ײ6����w��@�t�ȓf��E�VC�٪U�q�Q�~��=�ۓ�V��V!ȝ&��	���������0����S����W'K�FTpP�ں�y�`�7�Fh�oR�9�RL�$D���O�"b�LU,`Q�r.F�9ܮ���AC�<�AI@E�]DP�5�~��ca�u?N��O���I,d��Q��@�P�r�cg�6W�B��8,y�`i�*_�rT���D�9�V D���׊-2���r��1m���Um=�	ɦ9ɚ'ћ����#.���1��@��TP�jc
O"�	0�L�m�Ȓ#E� F�hs�m�"��Ě���2�~�'�d�I0՘4�֩��KE&5$���U�c�Ы���$�^���:���a �=��x�yu�����YgB���`Ƹ'�ў���ep���`����d*��!P"O^ͨ �7���%oQawf)1�"O6ի���jL<�u�M,c����0"O.0��Úf{\�6���-�b"O�܁sa��$~`�RbK��Z�s'"OF1��Dy?p	�!7D�T@r"O�ܲE�B�!M��j��ڣz=�Ԁ�"O�|qrB�*+Ī��N�����"Ob5[���4^�4}�7Ƕ=�8�st��;�S���L�#��K�-vd��jXa�C䉏d�l@Å�0@��A�4N$HB䉝^�P����*U# 82�ס'*B�!��0��,S6~o�&m�\@&�'ў�?-i�AK�]���E�:��l�� "D�p@ �Ge�,��%�	{~)�+*�I<L\az��y��`� �M6p��X�B*7��'�j#=%?�P��Ը([�끄֋I�HpQB�*D�$ٵ���R�d�ɂ	�x`pmB�(��<��mۓ>�N�3�h؏�U�@M�<䡈(��Pra�6��q&��c�<�C��'�"����Qp��AA]�<Ѳ��=���5Ҋ?�����E�X�<���Y�pҌ)B �.R�	8A��k�<�a�:�c�/E C��k��e�<�wK������T4R���vNS^�<I��W<h���m�6�4���\�<�	̜7�����	Դ1Պi�f/
[�<q���!C0�@�5�*Ъ��T�< H$��Rc�
)5�� �JK�<�;lӰ%���* �6]�W ^D�<�d��d���*���wG�g���̓V�j��.[�H�I����p-@4���f�K�.��S��SD2!.lE{���O�}
�Q""���'A´P��|rmM}�<I���eḾsf�
z�ٙ7����"�P�S��MÀ�K�/��@�Z0n�"�����<���C-w"�T�W�\�0��T�y�Մ!C޼c���)+"TsjL>�yR�j�Qˀ�W��ta�"jS��y�H)��QA`��4x��tj�kD5��On�~Jd�R�l�"��D�:����DA�z�<9�a�7�$�C��Z���.�by��)ʧa`$��Fʗ�u!ք2ab6=��ȓ{9H8�v�J�xe��Ł:X �Fxb�)��O�/Щ��B�*���iX�D�O8��4����2��/�P���"O,1��H�X��,��Y7w�
0kw"O�  9+�H׷e�&�Ip&��f�Sv"O�8+����$ٖe��-4I�Ix��O[��H��扜O% ����D'����j��L�B�I�%���R�B��╱��O�4zF��~̓�M{��E���>��:1�jX5%"�vXKR�+*jC���`�a���n ���ٜtM�6�f��G{���Y�4��k5�T/=>�����Q
 Ka{�O7扢Uf�B$Ī���bd YݜB�ɴ���"���~͢B�������Ӣ�a�S��6Oa�����Kry���[�5��"O����ꍽ$���S^ڢ�!,�M�ܴ��S��y"fO�CR=�mL�@	KfcJ��y�h	6st�����/z~��JA)�yr�'��)O����|�>1�C�KјͲ!n��0������?)�'�*zea>��Ġ��;�̥9H�HG{��d�"p@v��!gBS��:�&�y��n���R�
83����H���'H~���@�5�^Q�a�Q�7�I�3�!�dQ0���k�j�	A:�2�G�*xX!�\:mI�H#�&>�]�#a��!�d���4�`�9��&@�+`�!�$��H�l����*,��.a�!�dğ+_��4��T�xfKS=�FpG{���'�)#dOқz����h�S�b���'Y���Ȓ+��t��X�DD��'�a�E�~��P&іGSm��/״�p>QI<��E�Dr�����*��Z�*�[�<a5�O��1@b�_�©���V�<	�I�C�ڥ�@_ZD�+��H�<I5��3$w��#�GZ��
��\�<���ֆ4Yh�G)�-t%���p�<ak�-��X=	D���Gj�<y�ϑ0BC�=E�ڝ��ж�p�<����jEFp�@엘n-ڜ�L_U�<Y���#�20�f��E-ZS��N�<A ��v��PA��\��9�+�s�<Y�M�J�(xq���mlP=�R��r�<Qa�y?�AqGbO44>�A���p�<��FC�1��<���5
���#f�WP�<���zx��I�F3_�H�(x�<�Q�MU��r�D�t��!W[�<QK�kI9���,Z Y �$�Z�<a�Q�,�����U�4U01XVɀP�<��`�&z�嚃�ըz����b^L�<�Qg�?~�֙�sn�:<=�&��!��R�k���I��z�l��,v!�Ȫm�"�:A,M0��p�H�J`!��E2T�> �:l,����\+Q!��"��]�B \^� #�K�/_!���M9|�JD�>H�]�!��K.!�):m�@A�,��lN�?!��ё5�̸R��K:=��-��L�_!��I�G@%��*1(D0�%��7!�d�5fm򤻕�k����A�P�ΰ��')|ţ���v��$
�F�6P��k�'��ijgf��"��U/x9}��'Sl���	�pF��c��N	iZc�'��f	�?$6}UH�dl:\@�'��Yq)�	,��5m�!Z�\
�'�
E	q�A-�0+��@��	�'��X�#Jڏ�Ms4IP�\j] ��U��*^�PP�u��ճ5�+D�p��ԦPT:�揉_��p�r?D��wj�:8�Ęwˏ9;�t�U�>D�� ʼ�A`��2���H1ǌA�{�"O�m	ѥ�)z�:l"DE�~�A�""O�D�EX�x���DC��J(�W"O\����z�И�F�L�*��%"O�1�1G�;��		U�Y\�!�f"OSȕ�D2ZŸ��	'����"O��S@�S��
v�^h�\(��"O��jI�-I.�(�Ni�գ�"O�`��X1Qc��.۷F���"O����E�?� 8-�#+H���"O��
G�.x�r�@��mJ���&"O�!��Y�� ���_�F%X�"O�0r�I|�\Y�H�7���d"O���'�G)b��H���!�b� a"O�pR�HK��6�8TBǠ)�fLh�"OL}��n�mF�P���ub!�b"O\m8U��'��$�B�r����"O��$+]���UO�7Rd[�"O��z��D5.
��	��M�yb���E"OT�ee�&p�)��C̃1\��'"O��S3D/s��뒉^�OR�,�v"O0��f��Q����$/P xM�4sc"Ope��o[�V��EP�H2l�V�	�"OJ��S�IB��'ٌ�d�q�"O��(�C٠=h� Mo�P��7"O�`�#�U:$%1���+E���"OB���\��5�B��w0	"Ox5 ��$�PI��O�,F�J�t"O�%��#n�6|I�I�9}�m�D"O6��*ƯB�NX1� LTt�)"O(�zs$ڒ��h���	`b敱�"O<�y�Câ}ڔ �6��9`H���T"O�a�-ҏin]&��->��XB"Oh0�fE��܉�*�b$0�5"O���GC�u}(�P�I�2�}��"O<����:��y���42��P��"O�ٙu	F8N��!��-�p�2�"OJ��aУ}�����ʍ#��[u"O��H���ZU0(���0n�M��"O�t2v"�)�| jAf4uYj�rb"O�z��8���Պ�DI�s2"OeR�e�U�H�"àܨPA|�aw"O��P�/��7cz\ `�T* V"Oz)�o�
۸cp@��nB^�$"O��E��^��B��G%4X�4"O�m;U#˭fvN�i��U�BƁK1"OX�AFA�,;U�PHS�^�.z�wX���r]$#	˓\:�qH_.%�-EK�:)�d�ȓY6� CTʀ�{�~�ش�B<'\�	��v�<����A����Z_	���'�&�l_�S�O��ma�`�(Iz��0ʒ=?�(�R�'aN��/Be dH	�OpQpJ>�gh	�0=�`M!66���P�h"������V����ɂ{>�p뗃B8~�����ip�p�ȓ-���m��3��� ���-9�T`��z�'0�pK!�M=mG���Z���Bݴz*�	��*�S�OAJC����܁e�D��q��/�x7w��BkM'&@�͓���2�B2D� �v�V2'T����%|�Li�ñ>�H���O����D��3p�x�*C�}*����	�N!��W�7t��p�K��P'�|�Ꮬ�ִi\i�>E��4+2����_�'�hhWĝ�*��Ig}B˗CE.u�D� zF�g���?ɜ'�ў"|R1m�1�8�+4�icJ���/�z�,����)%��� ����G�ipg�6^|[��OV��$_uh6����ZC����I�"��O�7�o���~�4��	22�U��$ ��B�p�2D�H GiؔAS��P�b&��y��q�$͓Y(�c�pmO�OmpL���)4ն����Gt&jI��'�����D�8�nԻn�$k�)J�#;p���� Y�ѫC�B�|�����1Oc�x�|�J�ʴ��6`0dYI�J��6��W��`8��CU�է�$!"tē>
��xp�6��ަ��	d�OZ=q�/Ð��,pdB�'Q����'�
�������I8N���(O����(I?F顴Ł!	K<�I��MJ�az����FK�|K�"WJܴ !���!�*�����',�|3�N� 1O���E�$�=Sx^��'��
�%f��A�هȓoE� (�#T'e��,:f��s��'�:�AV�i1O�O~��-K{V􁖀P=AR��C@���PxR�i�QӒ��b�h�o�!a��LYg�'Q����i�Z���x�b��-�u9pg-D�hr񫕬}2���膸W^�c �%D�h� +J�`PHp��`�T�ht /D�tIg�Ǆ/���(еB�90RA1D��Z���z���i#.[=p��2�<ړ�0|�".�>�q��b�nsR���(Wl����'�o���.D1�N�4644�X��_��p=1�}"���,x	{���14�%��d	��y��Ʀ,8\k��˙2E��ږ���y���"h�R!¶l�7~��8�%�����=��y�m�ؓ$`p(�8��y�E��*�H6k�]0��4o�qZ��Gz���':�{� �p7��Ŏ��G�Q�	�'hf�w(NS7Z�H��@Vnic�'6z��DN1	��Y抐>;��|��fJp�!�.k�Z�f�Z�X�p	��)�sg` ���$�S��y"a�?|$bD��	9��ay�#!�y"�_�PP�HⅩ� \���#0��?��DR�E��7m.LO�)�2���lG�J�h�� ;@�B"O^lH�N̛
���bT� .�#��'��x�	�"Q3b��.'Wz�c�AQ���O��0ڧ&�Ci��M�Z1)�	J=纠�ȓZ�T�za�N<9xq�$�9B꼐�ȓok�A���p����q@8�'t�	W?!���S�(��� �5�\[b���U���2v�%p�5�1^�\9{w:D�X����
^�v�2�؞uV� ��8D���f�'qv��b�L`r�7D���P���X��� �KS5lV�P �*9��(O�֝�m�rĹ�sS���&�0	N�	`��h��賆���(�X̃⇉�$��|��iK��HO?�d�5i0I�`i݃f<��Q؜D�!�Y�>���sJ��A��H�ꕩ���A_��0A�G��+Q^�
��C B��Ve>D���E�(�% t/ݛ8��0zWn<D��J#��3$Z;�"��o/�|d�7D�\�핰~-r*���m�N�HT�4D���D�
23Ķ���'�>��)��LD{��d�O���K�Lu�A	�J�lv����-D�0!ꕾR��beG�]V�H��-D� �0��	.ŒR����ڤ�Gn-<O�#<P# Qj��˞1?:�c�Y�<���Z�a���3Re����BI~�<A�E_H�(a���/�z����_e�<1#��|#&��sӽ3be�A/^X�<�R�c�I��֐9�^�h偗R�	D�� te��BZ(��yTf ^xvI	��/zQ?�#Ѓ��U�f�C�H6}���"� &D�hQ@�B��ڡ%���(dHT�#}��O�d U�)�s�� �!i �C9&��)qF�R�Ȅ�G�q�f�&|N�X�q��x�PȄ��@xQ�ǂ�8m�t���P��كA�)�镻���v�����	��/�X����Ik���B"O���G��<QA�uµ�
9j	��I=�HO��0ChܣU��,�r���eG�|,,���>�I�y�:�23`��Y�4�Aw�0��'�b6O�7m6��~ڂ�\"uX^��S"�*S����6� e�<瀣.L쩳#�T�RP�Y
JH�<1UL�Tt0�����������H���'� 1�{��#
�5Enu�6FÊ4�T���C�����ț�`h,��b�ǅ�U�ȓK��SEA^=?��%�3B�%[*�ȓg����׾�sÇ<@7�p�=��'��9OZE�ԬѻM2l�`��-K��!��G=D�0���˿G�p1�®��M��mYP�;D�L���Yfr�fpY�(_1j�=���nPa��OPhȆhM-d�ɇ�x��pIʵs' ���n�fQ0��ȓY��!/�t�p��@+~�����R�<���2��A wD�G�@p��UN�<E�D�;�t�y���$It4�f�u�<�����(�PПM��	���Cn�<��H�k�xXTHO�X$���B��8z�8Gy���'���am�a�sI�;���'����mNs!�6%L-+��'�" q�n5�D@W�J42V���
�'*末Q��X���4�b�R�����y"ǜ7�ȣ��J**������yrf�3f��i��a[5&h !N��y�b�+�����+݅*g&4�ժ
��y̌$�"Eq��%���$$�yb��1(�D���_.Tr��:�@	��yR��,��ѩWD�GT�i�"�y��N�� Bp�P�G�α�r%��y"�-&�9�@ : &�� �L��y�څr���H�%�f��9㰠J��yR��e�)w,6a2��P bX��yҬ�5_IBBN�c_AC�)ǭ�y����0��$`�$NjRCǊ2�y�+�5c֐�F���<�6(i�oŝ�y��M8?"0�;qL���� +�yҊ�F���׭�"{�;�O[��Py�	��U�����^���=X���R�<I.��,���!O�?�����O�<A���d�sǍ�V���#�Ls�<�b��a7��a�/"vc&A�@]t�<�&��	<�&Q��ǩN��yUe�s�<��Z'� 5��Ȑ&@��ճ"�@m�<���/�V�����2���cQ�k�<��l�$d� o�3T�q�4C�f�<� a� )�j�,�)��{�<�a�ݎ�3��,%W�i�d.T��ф�DL�k�ꕛ�z�aAC,D��'ۗP�
 ���S�%Te��,D��s�fb!B��Q#Kr��O)D�l���ejF@�6
*
��0#��+D�d�g+�/>r��a@g�1b2���u�*D�4���$�8�æiה;s�dY�&5D�2�.D,O�$����:cL��֩4D�(ô��R�գ�. �RIY'e1D�� 2]��m�=C*���W��T�"O�5�N��v(��äܼ��%�4"O���iA� ���5��"^xq"O���N
_``�� �5?h�R"O|�to�:1���u␘>إ�Q"O��;4��mJd���m��"OȜ�2J�wi�(�Α�Ha"���"O�g#��P�ېN�$][����"O�%+ȳW���@.��`Ufix "O��4ɐ����*&��MqD<�"O��(��I�x���������"OL|ap,]�(�:<Ju鑮6�,���"Od����݌e�<�Hg�+<��@	�"OZD�UM˺bSJ=��&"d�q�q"O��(v,S�8��\qdo�3U�{��O|���K�|D���2�p�b(Cf�I}��(E���VS�1����*�jC�I��Y�A�F��uQ�?i�vC�	�ɬ�2�B�N*M�$D�r�FC�I9,�(�2%	�,oF$}�e�C?�0C�I;ttA�O�f�V��'�.3�B�	1=��0&��}J�@q�b�* �B��h��L��C�a�|�&H�D��B�*��M����6lV ,���R�B��*!���qeף<�f(#�AT�U��C䉭7��ƌ�&�P�
�CP�G�vB�	He[��2�d!��c[8(B�I#G!1����QY����}B�I�^��;2΋4#�HY���6�B�I5`"��`c�+�2�򡬀�.B�i�Z�{���R��H� aC��^C�I7MO��k��!��� ����P�6C�I8T��8Q��2EQ�l���=`�FC��]����ք��c����.�3=�&C�<GvDCՍ��8G�xq�\�TB�Ɍw9�x�aAU*ּ�v�A�w�B�	8���UG�6B��h� 
\$R �C�	�P���2Q6���ז��E���-1�h#
�	�~e��
d�'��AdY5�d��!�Wnx��l<(�`�
.�<�I7�G"�����	y.�M�������CуU���P�$�OJ�[�+W����tg�=Z�>R��䞭C�=Q�ܛ\|*�B���'9��2�������ЅolqK� �;F�U�����y��Μ��󣍋a�n*F���Ё a�:<ݶ�)�Ơa�TH��N�
�O�DP�w��h$-����v�/R;�ݱ�'�����9 � ��Έ>R�p�H��Z: �h�ȣ�΃N��c�Ɖ ��#���=�O�@��'7��j`�_�D��,���'��B��A���F@�6
� `1-��U`��y-�s�mY�Ϗ �¥qE�ݦ��I3DOD	��R�s�	[��	i��O�swÌl��dU�L�8�y��ڲq7֐�^w���-��]�i�K a�l�c����y2"��1y�u{Ҭ�MIу��Y+)�]pC��5"�p%��P?l���zb9"���"x�X%S�2�\x��L�Y��dRvӵ4Ѵ�z��'��4�
Wo��K�M� `H�C�e�~Y	%FZ=0�.��B�>kj�8vI֖Th��3�Q�Uj�����\�3�2���<n�{SI�'���[��$��A"g��|��Ir�i�:��z�$S4$4�k,��v��@bq�*cG(�A#��'��TĆD���f�禅cS&�4���Z�D�xH��ʄ.b�@y���)PFR��D��I�:�3�f	2���:%�|N��¬���9�J9L��At��+�rh�t�i�`]9�)�1:��}eԎ�<�4�?W� ��h�?8�<:���I���#��}���ۀ#�"ע�\?�+$M��W��6�A�d|���g)�y�����ƞ�o;����L�(��>ѷ�X�T�:���L(<����UI��^�Pq$�W�.{Ԁ�#�Ψ]�Z��U�N�@�n�ٲ�ͪ9��������Z�p!�HV�(w��s�	�J%J��0b�9)J�3��n�'a��IīuH w�I�q�|��Uޒ��Ĺ��Ĳ �l��Gh�l�0hON=N8S0G�r�zh�VM� ����tcE0�h�i��ɏ"rV0Pb�6��x�)�"$F�牃'1@�I� ���9j2���!v\$x2�0��p��#%G��8��=�ŀߏ���4�$��t�A*БY��P�"I�piB����OZ�æ�--�`=��-)����ᕻmND��k�3Lܤ`�2m�_R�Ӗ�D�,�j)�4jӠ%��K©sК��b�W7���ᙢ9z���.�	*�vaU�!�O� `u��ߟU����J��4P����o��=y��aNڎL�"+�e�*�rU��G_P����J²7W���?�r�I�G���ɰ@��22����'�Ia&>�����l� ?�����̼sj4QX�G��-:�Kp�ۘ
���SW�R�qf<���¸:���P,�qo8M`��F�),�#شNDfsf̮�T���h��n	�=i�a�f�`Bњ7kf�0�jŧE*�xKA%&�9j����ĭ��
�@�z!@��A A^��a�]����Q)� �
$*4`E�HOn�x��@(,�r%NB��l��M�	tL����"R�4�A�N���8'��*)�!"�� �D�1��
qF�ȓ3/�+9�b%���U��jO><�����CX��p>I4#�,2+f̘�%R�(�Ӥi�>D1L�*�BFx�>Q2%��:L����C�4/lаWS�R�.���ؿE0JѲq��&9r��F�5~�m���xx�ĻM�4z�E��]�Zp@�͗5��Dqa-��4\�r`��fi;���L��	�4 hcm״��PI�mE.2 F�"�C��rM��ćڄ4pj�//ôm"�[�.ƸMC��n^LpP�I ���,�7#j����ńA����ƇH!h��j�Fٵ6�<E)d
�)ow�4����)"c�m�(�D���.,��<��L��"�)�A�ӡGX]@6�
X���Cr \��$1*D`dt(��UL>$���S DVMp&GB	Y��� ��?T��$�B��#vPh%Hec���%폓)�̢<�b�L#wQj7�z��%��
�
=��c� 3lh�K�bX�*\ι�0/Тj9v2�8C"�٪��:�)����3mb�+$�,(_ȵ��ș}W�!�+��)�.�C�?�ē{Q�Q��J@3N�!��
�E�d���e~��Wd[�6�"�#�ĞU�C��J���AC<!'�V"�0L�ro)Ri�l� 	u{DS&��d&r�j�����Q�ٱU6X�c)�u]�@a$����CE��4:��I���I>L��|��0��H}��� Ɗ".��T�٧<h"� #&�DJ����ł6-:A£�1g��p$�]�[�H S��?l(��}���H�:I���3�̃��\^�4��Nҷ%yH É�X��M�U��<�&I��P2�.��~��@g�;K���%�L�D�!��B�Z�����/zR�Y�T/Ě��'�>�;��͘��QX%�;���تیp�q��ZI�kS�O��PMI��ȵD�87��$��o�*ה\�@�[F�sCϠ���J�ImV���a̴'���XW(�#[��1і�cCܣ�VL�G�P#�EXCM��w<�	r����?"�AŦ�.*(�����L�h|��Ǉ	�,eTԪb��+]¤�'@�xr���&/.!���b��lz���gI�)o@6�ӵM��󑲪6��/�.hVKڥn� 8{GCD�X���*V�,��d��i1r<V���aY-x�~Q�B��9��?��X�F�#~D]P�B��GѠՉ��Z�a�p�jR��p%�1��9qO����D�s�j��da��	���$�b ����=S�B��Μ4��E�@��3�N�%��ea���;�<8ұ��<R"�xS [�4�h���8y� ��2�i`#�6��:�A�+fR��{t����|��]#���Y���}ބ��TM��b�p�I��ٟA���M�K��p�hWQ����j`���l�&i�;$�)[�6�{"a��=b�h	�\Z�}�.O*��aH�  �h]�V����|�C��)&>9����(��:�'݇y�Fa��e���B� �Ex�q��OU�\>|��Oʪ ��b܅z�Ny�@�6���E"7�-����7_����,��C����i8�-rq��Ѩh�!�m���1��J�ꨈ"�j<�Qr����@�䡐�p���&cY���e3���L�P	�o7�a�<Y'iؓm0�E)�%˷i,��[�%�W
�lK��gU�X۶b�:QW�%E���b7�AA6�J5l.���'V�`K��ܗc\NIbᑔbEpԲ5e3C�=��$UDm�%M9�D/_[�� 2i�JA �a;xL�tjK	AKζK������u���"�*E��@�<j���� �ڧWSZH�7J����	�<b��;3aS�(����868�'��`�4�̚X���a�)3�쁡�iN�I�ތ�OD�y'�̉/�5A�Y�_7��6�N+.TH�� b�u����e㊠kf���E�	-�%i�]3����-^P��I!]x��g��@�������0���Xy��C��G��
Q�!\z��%
>A���I$/ ����?�(*a�9u:
�ّ(��1�VYs�"�3�њ�423�7�& J�{�j�j	 �%�=�ڰ�U�Wv�ʢ!�*Rhٚ���_(�� F�/ΩZ0�vqY�f�����C�^1�b�����RcK�����biV��	�)4��Obpj
L/;F�c�ʡT*��G�`Nv����* ;>=�3��x �t�W :ZΨ�c��9����� P?FMn!��EL* :2!�S/{�d�O ����z��c)H�jʍ�'��XVc�ML�@ ӎ���#� �b:X���7���A��ѿ&��ԂP�ԏH����J�]����ˮn\ݰ���Mc��;J U�%��L����;E����K�B���ƉQ9mh��.�'��HPDH�l���f&�9@���(�kF���V�P�il�)��Ң[�,鈅
��>Q���0<��-Ӎ^��0ӡi��hO�%Za�̀Kf(@��} 5�R&E��L!�� R��]���P/aXP��t5�[�"���tiP!�RG��r�N��8���r���q#`iA�:�\M�Q�Q�^Fz��Sn�)&�|�u�E��]�u�:08$�#��<
eX�$Y����B0<����`�A��u�u� ?;"�Ϛ� ix���P@�a�j��{G͎���I?�pA��E:is4%x%d�-*��3/W�[�����SH(�2�YI��M�a�X�	��Ys��^��a�dIݦ˔e����6���ѕ���K��Y�L���O>���A jdȹ�f ʷ3�F��j\��Ɔݩm�x�Ȕ��0̉� �loܝ.|�p+S���6)B4�,��ML��֨��b@1��2�ed -�QS���M�'�j�Q@
,�9�� ��Yg��,2�Ldʰ�^Xt-:p@�s"7���IB���.D����B�^k���$AD�F� \����9�,	RGN+3|�1f�u�'��p�q��cG���#ca��xv��9<s�l�!��'�%D��Dc흝?g0����'-~}��,��7����f��*�@���V<#�/[�M�l�a�L�nT�8v�ޟP˄j�B5+�Q8��Ѳ�P>m�0��u�Q�|B�cX�/r͋�m�W �Mrf�P���Bc�D�֪�I�*5�q�òtMra ���J�D��"0 [ǔ>q�iA�+��	RLB9L�T���k[7D�0�AK �*��T/D���]k���(��9R,:K�V����[6B�X&��VtNq��K� ��L0T��c>�<YG�&	�D�AЯIA�#<�h\�9�j@�	�	��:1ߑ_<���ҕ=�v5� `�/��	ѕ��,v<u����
��B�m^�[;��"��S�8�d�P�߿z3J�3�)
�~Nl{��DP�����h
?}�r����Rw1��֐?���J�"�, ��47�\3���=�Pѐ� t0h;#!��% ����+�0��B�6�@sb�x�� �epf�G�"	���fOF�iI6�'�~��Lm�^�0D��e��|B&�Z�e�^|��z**��L�cc���UOĄ}/l���BR�j̾�x�&^
Y�NX�w��~ >)�FKfi�I&Tn��t�>?L�P���0% |j%�V�O�\��3�	 ��<X��l����8D�P��̀3 (H"ՠעa��F��>`pc'�n�#�����Ō���`���'��pF6 �TA���:7F�	��E�2�

0��t�c��#sHS�cѫ%]�@ys�>8T�9�3:�b¥�5��Ab�E:Mo�����ؕ%Z%)�$\������p��\SwK��2"�����M�U��M�c�S��rc�J�<1�i�7<@�@e�X�9$��$S��i�AU�R|��2��R)�y�Tlv���Fώ�M��=��J�yr�J
j��4���\;�6��T#ԃ��Oi0� � �e!����׆1����.K� ��l(�B��?ӯN�%�,Kp�`,��Ӷ�V�4���-L��	ӂXXuӕ]�SA��<X�����V�6Yy��`�A ��� {�nH�W�>}1ؘ:z44��G˂;�1Ѱ��N����(4�~�:���!`��� (&�S�V�pj��E{�&��Z� ���$�,b~Apg�3���Z�(C��rfg�vM��P�O:UF��ے�,ayu'd���1W*�4yW� y�E[;K%�%@�C�#�l�AU4F_�#>yW	�����/�L�c��|�ci�-��P�@U84�1�Tm@:�����@�;��O���3ɏ���\�@a97���ܼS5�M�h�0ƥ�."���Yy��Xq2�P��ՎnZr��I��1����j�"Ed p��
�
5���6��i�� ِ��p��hy�Aʏ�'OLx�mY/��'g\�CSǃ7*�KPh�o�Zl��;0s6t���|��&�-gX�k#�5'�0#�Ȗm�Pt����;0�ތPc�2(3M��T�Z�(�Xc.͉4�"�Q~LJ���Jᆘ%;]^i�B�j��D�3���D:�}�s�.p��.';x�X#��8\^Ѳ��>ks,�(~�����Y�"�a��$�x���a�G¼a�j�H��/���]\��LS`dP0l%4�)���b�L��i
6M!�BWAJ�Jf�%����'6����';� /� /�>xk��,{A���(O��Ӑ�Ў"��1q��~��3��DDV���G�^�i؄��u!pP%���~��1��M�Z�4B�U#X�2���U(�t���k�pP�EѢ6N�Q�H5B�Ȕ�fmGRQ ��R�@��P44n�y�q��=B�D��W+�(SF��$�ʰt͂l�,$x�-)�O�)y�,0�^�+�l��ز��v��5o�)k�K�;�8 Q�o��Ey��X3�H�S l м��V�;��č�4��A�]�ؙ� h�'6hP�@G�0b�:�������;aC�N��Ya�]�P(Ex�S�h;Q����������4�������U�I���3�@
T��Ջ'JY&1,�-Z�K�o*`�ބ�.�+Bx�D�|zu.R�K��p�7��˱ �Ri�0���	��|[.��	���])7y�% bJ�#�BI8&e�u�̥c�Z���Bd�"�B�������)$�,AX3��k�HFiЂ�܉1NFlr���{�y���J@y���D	vk�ݺ�@C�*P�u�̙�B�0ƛ.m�	�˂E����'�B-{-���b7�9P�(O#�B�&2��(���'������	�Z2^-�"� �@�ĘIr����yblЉ>��Pr���C��"̒�ēA���E�'8��)z��8K>E*&�+��<��B�;n�!��?D���׼5�&����@s���D!�d$`����8��$�>�t\�gnR$uHƸ�W�'��t�ȓ�!�@B� ������k�(<a("��8�ʙq�>���>;Vnܘ�O~2��j�jG�z��_-�0���$5���J�_����Id�\ġ:�y�N�*_n����e`8<���Ԗ��'N�,0�ED�p5�xE��.O�,oJ|qE�@%2�� ��>�yR˞2v(���¨[=i�X��W���!s�"y�S��y��7�i�c�6]���P6"�'�yrP,_�$��Ǯ��@A4�@��yR���[�8l���ܰJ��ԥ�'�y2f� �����!
�o��e3%��yb�Ăg�� �7��bDڠ���T�yb'U������?4�:tz���y�?�B��o�8�v�ಏ%�yB �%,�f:ŧ��=����2GR	�yd��J�t�2"l�*7vP����ybI_�sjz�9%%�/�H�fe�y2��1q.ă4'��qc�Q��	E��yB�VS�޴���'|Y���#@�y�c��3�"�cA���y�����*�y��˪d����'�����'�yG�> !��F<&ݸ�����y�$F�z���$T��*8�c�ه�y��8��t*a�}���3��y2
�qڼ���ʡA7��ʓ���y¢KU2�����h�L��	ڼ�y
� �`��cL�)d�K�+�l �"O��Q��6<��'�1[8p�"O̼��I����CÞ�X��{�"O@����P��Q�� ɭw\�(�"O u�4�J
a���%O��mԔ�[�"OИ Ө�4>��\!gxF"Ot��R%��k��Y�dm "OF��*ŵ^�ٳ�7dF`��'SN�@&� GN���up�L
	�'~��G��<@Y
���B.R, ��'H�`�Aˈr�\p0��-@���@�'N^ԙFN�~
�M*�&�A�~��'l� �,$��H�� �Rs����'������̱M�i��%_<�P�1�'�x�@�
Vu��㇭��c��5��'��:���4w��!9�j��H"����'���q�m
�ck��+%ș�I,��	�'���MO>{�����j�:�l���'�.�2�	A�	`�L�q'� |�L!�'{�"ԩşQ��͒ �$ V-��'u�8(2�]^����D�k�>T��'�K3S�[)�aJ�Ù
	�	�'���u�ݯt����ϳ�����'�peP3�mM`x��铛�.��'E �b�D�kz�H�%U2|^�!��'�:T�T鍣u���̐�@��(��'�R]��*��>�&�QT�^�F;�}�'�8��GAB������ȵ@kj�<Q�A��`��:Ya�%1w By�<A"A���,�gM2�veÈ�p�<����q�bd �Ζ�ƼHd��h�<I����>����@E*U�r�b�Pg�<���UF�[��\$���ţ�g�<q��R�n�U##-�x���w+a�<I�II�j�����)\X��f�<��O$qM��b �:H3
�����]�<�l_�Of�xВ,���;V��]�<1���2W�����
gc�B��+T����ҖX�ʩ�e\�b�	#�)D�(#
��!�\�ipe��")�Hj'D�taMF�$��"O�ҺaE	� A�.ڠ,�8x훦P֒tF��Ymf���nI�q1f�h���=An���MRa�3%��ȴ�ԩPRC�R�Y&�X_h�R�G��t�i�H�N-*f'�-^>���d"��.�Ubbs�X1SI�(G��p�U��G����P�2,Ұ)��`�t��㙀�y��? ~ݨD	��P�&���^r�2�;� ��I��$2u��bM���		=;���N�_�
]��M����WLI=!��ī=���B$�,"��H��FWD��Өɂ*L��RN��u�zT0u��?���=��O�r^�0#`Ǐ�8��h  �LAx�43 gO�<��@p��}� �`q+3w�D4Y�O-&_N|д\1��3W�D�4Qa}"��?��h�E-U�y!��5��U �aa��7aI��c��O�hS��� � aj�'*�
���A�2}�y��L�jǐ�����=�`%��xز��C��J��	��eZ�Y����|��T��?��GX����R0�4�� ��s��Q �M3@l�Y��'o��+�����@� ��=ʱ��d�����(M7���`��9B��(��\>��h��m^~�	>��`#��b� 4s�ѐ���'FX��q��.�����N_��v���D��!0��J�ՋF��D�������J����Y�i��?ҁ
�!�r���i�퐑~f�=�.�1��	��nd��ǆ z�Dh"��=�^�9a�Q�xm���nD�5�����P�Q�f��]!��+"��GBdӨ1��,_�($�E@5���]�ay�E�9F���K��P\V|rO/FV�#��N�\���#�e����)V#-��S�s�ZQ鈼?�QA��I�m�A�ܞ!c.c3I���0���}:.]Xa��8�\��'Ε��r��va-;Ĥ�C�/{�L�:`�ǜh>�Z c�(8�L��g�U+�~ș�a/7ܔ҃L�$'��(������)[R!��p5F|�D�O��K��]=gN&XC��T�EN@P�qĘ6���{� R� w���U�JJ��9�X;B<�0"����Vq��DY0���C�@r>�]�� �hB鏅�^D���h�d��7O�L  
5Z^nę��F�Ju�|8I��Jt�U��m�n��'� ��	h�/��j�n��A��&wm,ÕDXu��i��G8�Y"��3^J�D~װ2�D��K������r&�:-~3�.T� �F�1�-.n��W�0��T2���MpR,�Z&� �%�ez�ƞ,HH��PMX�.��"ݦma~���=E�lYU�	�&�D,A&�� �	�c$HV2��i��őc?�q` ��0>C�D	���'�F4yV��y�&]&(����)�3����V�=qf��5_�D͢.�;O"� 36�	^c�4�ߕo���k2g-^��e摸G�e�f�[~��f��\a�+T l�1���L���b�����i^�r�-	� �	8����S�^[T�(�嗜L�n|�ɩ>�-�����ꅝE,����Fh��$�p`i�B�q��y�z��F�΀	�͡JD^�'M�I�FP�OZ8��v�p(!h��Qi
��łh_2D!��Q¦5����P0#M˄,�Fb�H�3$\��D�,r�"(җ���z�d��,Jf�W���p>���׶4s�s+_�r��UF���raC3�@1=C��]�h��d¤^��� �ϐF�~�ҕN��
K4l�խːsɰi�E�W$�p���fo�y�U#�T�E�N�cd�8Q'�K�p�a�3��V&�m��3a5���gY�8�DY�'�0�c�#u�i�co�S-�Y�C�1e<�4�Qg�)��5Q3��"�q�g��>p�'$�A G1;|���B)��3�8�R�@B�}����\�/�Z�Ed�*��"5OT�l�J��mվ_K<��hM Q�V��).V�NŻ�d��(O�=�0G�)zp%��/v��P��� 0�Jƿ��wd�}�*��b���
R�w��rA*(�g�B_%b��c�˧+��m�p
]DgDѪ���:l�`���=ʓ)��e�`*}�̌�uKE�:�HĂ�nP`��t	��XjԠvHD�>��(�p���`��:a�J����c��l�A�f¼;F(�-<"r@�$��6y=:h�$� �M���x�aX%��V��] vL��6x>0tHDȣ+�T���b�&L��eysu�",+F��/.�X�����M�bn�d�N6틸�Bu��ë́
Z�	�0�����[1�T6\�8�g,!q�H$���E(R��U�PA�2�2g.3T�Eh�
F��,#u�X8��A�Q��Y�pᔱy�9H�lƠZ�ĉ�	A�7�~��'F $�h��+�S��#���sr$x�F���'�(��I_�LЍ� ���,Fmr�$��� ��9�i��]Ȫ��I_�D��L����LK�@nz�D�K�(���D.���q/�0����r�0H�c��2G�ēm�L(b�F<��\�Zc��8Y���4�\pG ��Ķ�i�J	��z	1�L�v~$(�K�4��9�+W6�` g@ǃ¾�Qcj���h���M$nx�v��`� )O6�����+oH8�c�6^�.)(�@�Z���V��0<@|���S�0	H4�W���F��FP"!((h#��E {��y¡�D�g:��2X��_�V�)�&�" )��4T�t,˗Hڥd�^��b��1"Q�iưx��q*���	.5X�q��S�V�| ۷Z%e�P����T�3 Axe)G2i�p���`��!I/^Ց#�F)m�|��ኂ;(<�Db��<�|���ϸ'��	��n.d=HI!��դ{J�Y��[�\�v�26C�6 Le�@g��c��9��֯g8\qi�t��XlP�#����lǖkCfr��S�(�$h��E�0a�X��G"O0Y��{�C� $��|�@�@R&҆L�kBdX�5l_�C�d3��˴vr�#��\���ht� 7!K�Lc� <3��t���G�XCRDJ�ru�3S�Y���q�D <�J��
��=��	��c�<9�.�)L� ���ߌ)ry���6��Đ�4�� ���ʑ��@����Z)"��P�/�1#�i��:亍��Ҿ#�9��1�L�����,(�o��*;��!1	}�B�ښ$Iq@��27�� J3�,���"��|2b�E�`��F��O ��`�R*~ ���Ł���-ɢcS�J]2��Gb\�p ���)1.i�D%ҫ}'�c�l�t��*~�.9;�I�}���D�Ľ(�F�sd��f�tӡG]�H�\��2��?B�,[���7~�����ea"I��3p�Ά����I�L���tc�$��H�*X�!1O�D8��X�)�d���@�L0i"P�NK"���2DR��15
�q�B����� #��'�(;C %M!��a,: dj�o@�4�a�d�<!I,������t��E�����|�8�d�(�2�`U�&�����HL8�0u�,�@��=U��P�6�ߐnM�"\KT�;uJ��i��	pAV5�,�U��=T��D�fm��jI!�#YGJ��^I������ex6���O
��u!���9H��,�g+Y�B��p��J����OI�d>��uOĚ���ؒ?��4��I��4�增�Z���� .��	`���^-�ݣ�E<=���=��^juMP $����Ҷ���*[�e�}8�d�	E�2 )����M��Y0�L��H��C���j�i�m�$ڍ{�j���N�6���S1�Z7y��Ѡ��� J��O�m�E�S)=$�ڳO�h��E"�㟴_��8`GƚG������\˔��� wd�i�ظ)�^��u��,?��-`�F�G�����Lի_Μ����O	\rw��F��P8d4N?�Y��'b!r�&ֺ]�/J� 8��צС@n"�Mڧ��Hp��9䪽�KCE��	(EC֣~񌔚��[�}� �i�^��Mk�^�V�Ecg��L��0��PM��P�D��p�<�0w���.ͶL���pG@�!* ��� H��p�$�t �ʠ���s�q`���.,ݐ!��Og�X�ӇT.LĢ�3G���$
5�hO�MȤ����,듅1�-H��~�̣"���8W&!�Q��'�`E�W�=*��3�0�`�o��|{��뒍��8a�L����8p8t�	�4/��`�"�*�H|�e!���*=,y��%	Q�x�d�X�Gg0��T�Q�4��:��޼0��p�C*NeᱡC*v����c��Co&��T&џ?��R��>5��PD&��D (A��ƤU����4,�		��8 VM�oph�IaE�� (�����b�.|�&�\��80&�i̍�ҭ\�[4H�r�Л a e�v�ݚ.�ԥ�%D�tg�1�&�4kę��M��X1DO���7E���+�c�p���)�zw<MD�O;��	�
��釧R�C���+�+͐b�j��G�i�����N� ����v��,�p�`$�����K Jڽh:L����Ǳ�HO�U(RiU�w�����/r��1�i\�`&��zA� /(��z�O^w���lZ�P%x9��EZ�����8�RlQe�W�ZU�-0&E(>���Jè�x�4�R,��HO�+���WwJ�Y4�<n9)F��82-��E�Aj�~`�G[�^�P�)E��Un
`�FoF�1y��U�DT���C����i�pxCSړ[�@�J?Qd�}�f儦
���P!�6s�H���'WJx2�@�)	6�(C'��9>�u�V�D& ��Χ7p�P�scݕn^�|h�JB
9u|��&E�/����i�BuH�ZKƀ@2�Y��0 ɐ.U�x�̐���%R�i&�e6��f�{��D.C��Р6�a�u8��V?#�X�j�*��h"�}(FMQ `���D.@�����b�E�? j�J¥�	L�h�9�",�|��W�!Tt��k��G�x �bK��Oh��#�,SN�s)�eU �YP	9@۾��SᏲ"�`�a&��
�3��<�CrI�b[��	ѸBް���0&�lԉ�IT2#x9�oT<�|Q�O�:�F� ��ӪaJ�a�*1}��O���@��p���'!� �d�p��[,�[Gi_�v p���W���� »t���A��t�0�w]���խ 0TV���#k�r�VI��_� ��M�<� �h��U�M\Q>M�����]a̡�cb[�)\KsL�&pҌa��F]9;&�A�B ��5ʺHB��+iމ��BZ�,	t�K$���J(��G�	�{=�M ���6Sg�pa�b�(}u�4�W�\�74zE{��O)��ק�}9�M(�#V�Qc�T!��Xծ�YE�_c8h0�VC�2pn��5m
Vl�uXv#�j=z9����/e��$��+��=y�U�Q>��w͉?B#!��:R��{��P�|چ�{��!?~�K�
<����G.ʳ�^�|dmAКXa�4� K�N���a�6�>����1���)6������u�0q0e��(�6�ߎD��9��UJ؅x��� k��� $I�p�(]`�����$�F�^�B����[$Z��1n[�vbbDS���9ό��/�[W�F�q����p,H�Y&Xc?9#�GֈR�r=Z��t9������(r�=[�����$�|�h�� #'vܓ%Ȑ�^n�� *�DM����� 򭇝tT������[f$�3a��#�|�IW�6���&C���H6~�}ƂGIl�ք~ A����	����C��!�j��bnG�'~0��ޏ=�=����-/�pLD{"�	 K>XD��=k�v�bq�ܱ_,ɺ0��D�����,,�5{Q�.�
Y4A�=h�p�
1�\$݊@hѦG��	Iӊ\��&/]�A�,��A��`BabK�'���C�� �F0Χ��i4M������:��q1��D��XQ�<K1m��@���};d������㐗?���;Kg�)�a�,i�J�Ƣ�&x����'������	D��ٲ�"�E}q�~}9�� :z��@t��ms�8JŁ�?f�!xT�[�@����I P|H��X�Ew����A�h~�e�|2"�	c  a�&��U{X�SBO6:(֍�P��?Q�'<!��M�3b\�d0(%��8SrB�s�7:)҉��ș�7� mw�	&3،�AP"��ia��'f�h"��Q�Y��˚o�PI ��O|:�ɦf�:x��KW�������lSc�.T�&��R����;��O�ݒC+�� �qN�4�2��dҜ�(�3�;8q<\����u�������pk�>r�A�b���|+@!�	���Cgٖ >��H?	�ׂ�,���۶  ��2�|��l*o��ʓv�fp�S�1���2�&��/�$>}+���iR������{�nd����f�����U�����~C�AHFO��p<)MY�f�j� ̒XB�re�^&$� ��E��d�$�uĉ"R:�Y�;sl)�e���4Aj�;V2�yr�Ü16��1NZe���h��˪d��
��Zbf P�iBK#Lܑ�aT?��%����/�0���\���m#8��R�ÞN+R�� AU���-�ɟΨ�����(qʅ�o�zh �U����a�"�=|J�m�!�W�0�*�i !ҕ�p}���qO�]�2(Ը*I!��2�	�D��(�H�'?�<���ʪc�F�B3�02��� A�SyrJ͹f�ظ����A �2
�,P�1�85����
Gb�*����+S�z��/Nx�@dƯc90�� �p=�0�=�&�*�
<���J�E�6ߪ�K�.�,1�F��M�-wP�H�O�t�A%*ƞh�l��e�ğ��/�&QF���c� �5�F���g'���D�p����G�!6����N�&���9���={��,H�c_����䃵�Jy�B[� ��JAk�2��x�
o�����J.D��y�0��=:y(�R4���j��<�Pm��z4R�ȓE�r1�ǃ���2"fԤ^���&�(EČ)J�(���S�%�p8[���){��B�N���i��&���!�!|��J�F�8���j��O6 ��0�Wl+'�`(��'|�����m�(�L��h�:2�\��6D�8�2��/d��H)�OۘOQ�YA٣,���rVhJ�a�����'�P���%��̌zq��0�X@�ד3�X�A����x�JٴNa*@r�H����S/ ���[������ha#1$��
���>AB�B�.�j��vO,ڧ*�x!���<r�\+����Uf~ �� y��(�"�����I��!
�'� @��"~Γ�	��}���""ƅ,�B��6 s։`�f�625�2�"B�	�1n��e�$8���V`�C�IY;��h�"TO��!����#Ei�B��->@�-��D˗{���l*i�dB�I���E�� m�9�7i�o<,C�I�_��@�P�s9�9���\ cK�B�	'���
�m��Q����"K:�B�f'�E�&G��j���G\C�I<�5z6�@7@%`��ƈ�._C�	G�x�s�
q.r93uoRo��B�"5��A�v*YS�J��G]���B�ɺj���ѵ%��6�:qac[-s�nB䉜#����d�6Y.�82�d��C�	.H�����CձkN�kE�݊ )B�)� �#M�*U`�"�ြ(є�HS"O�-�vcK�p�=���هsȞ��"O�qY��i�&݋([�&lLU��"O���� (���0��|o`��"O���ŭ��^㒥�UM?CZ0mu"O@��1��1b'
qy'%
�f<�Cu"O�ds�fS�8�`����N<��"OXѸC�0\�vtZ�� o�k1"O�#�D0x��-�۠-	H�yU"O��B���r���m���8
�"O��р��@4ިHG*0� �˶"Of�i�oS�zB�`�S��2I|2��d"O�xG�������,aNY��"O8��ײ@@-`�NV4�X!2"O<�c �	����ț�ET\�%"O��	�L(#���pf
�.i�M3�"OD�Sr%��	zF ���ۜs�R��"O$���Is4���h�b��"O�pe'ъ�t�	���;Q�R=��"O*��7�J��f��BK�1���u"O�0C�-_O&"���)�>m��"O��	Ĝg����U�NaC"OB�q� N)?������$Rp��v�OT�	���y��rK�4\.ڄ2��Ij6��#���9B�3��I' �V��v�N�8�OT���'ؽ��"[�A�@����O�XdsB�|�#�O�a�t��rRb�r�ꖣqb��I!N�!��qc��A1nס�0|Br��Cނ BPOL�F��00��@y�(�1lҐ|�򩚭&�F�a#1vM^��D��l��OԞ0�c��~�
�4d�N�!�IW�|�ք��^�HK�}��O;p���;������Z$ I���V�HG���ih�)օB�z ��p��!*��L�p��i�S�'p0���,��,�v<���&"�4$�'C����,6�)ʧ�D�*^D�x�0a���O �J�D1OQ?ɩ�KUq��PqJ!H��K�J�TA7�d �>�U��g�L�[eƕ�N��ʷ��ј'��·�O|h����9e6���cÏU���iN>��C��U����<�}�R)�7h���Dd�emz���..�`yk��yӊ��'!rӧ��[w,�4�\<���^��0�7'u�p6��Ky�	|}"�'�L�L+���x��9��m
�$�m����&R[�#<�ç{l3��۪Qe�Q�tdH-RB8|�?�UjHG������O,]�	<a=�U.��ǆ�4�|B�Ƅc��>�� �����S�a[�eM�mĀ�<�n]m0��!?E�$@Z�t+ (�Ǉ�5�h�
��
�?A�"R ���5?�s������	����RȤ4c��Ī�;���1)$�H�	�M�hŲ��O�HP��D.��� ��v�,8ѩD,��c���i"Q��R�-���Z��	9��$�>�RbNi>�:q�|/h��"�Z����2��?D�3�I��;j\�T��N��a�7�=D����B�Sl)�w�	H�]R��7D�����P9�Y�t@�Z�-�A1D���������ҝUx��dc9D��� �Cd>��5GOB��Z�f8D��+V�z:��u���#�v�;`E"D��۲I	(y����w�Y^ ���,D�;PCV@h˰-C>D����*D���gڑq�z��ዱHP�a)D���F�"��t`���$ I(D�`!�%�_QTYi�d)Cx\�9 &D�(�3j}%� Q-���.��#U��y2Z�X�xġeÚ
�5� �0�y"CQ\,���d�:m�5"�ɒ��yR
��b���h�/�"%��.�5�y2OR��!3��-:�������y@�|l>	�0nK��,Q�'���y
� N(R�*K_zt@bX�<��0�"O\Z�X\aԛ��.uȆE	a"O��Q�LKX𵸑���I*��"O���e�W�� y��O��e"O��JuI˭o�v�c�d��;�1D�4��=?Lt8��H���I -3D�l��6}z�[�d���:ro/D��F�.$m^��'i�f>�{0�-D��9%�S������ <; 
�,D�l���F�U!P�k���֕9Ƨ&D��`d�Ơo7�D�˪D�ne�@�&D�c�	ÝMG*�fH4oaf�"D���᠛n&�Q1����R��x���%D�(��m�:�	��-R���@1n#D�l��b�P�	R<{婢�c`<D����n048Ȃb �5�ޤ�E&%D�D"7ŇJ�@�*-���da$D��(�_!C��r�^:���P��"D��؅nBG.L����<
��:Wd?D�pH��H���s �غEF��c�1D�H*w<!n |iPJ�3��)�3�0D��h7FR%9������PÞ5��"/D���E����Ad '*�C�?D��C oM�Z��))�]) �V��k>D��R�FO!`U3(�!� �r
;D�j�`E&#�tб��K�,�y��$D�,��[�;��x
��+"���R�8D��!�	 c�P���ID�&�@���!D�ĩ$�؄+TN�TgL�y���fg!D�XG���g	�p[ሏ͢Ղ�)D�!�
�&�Q�� �����"(D�4C���+��}����!Tn�*1�9D���� Ӛ:40y	�*�z�<5�u�;D���Dz:�fdT��"}�í-D�Щ�^)�5��$�� ���)D�ܲ���M��7L��t���3bo;D����L<u	֝��b�-K�ٙ�G8D�@����qhP�2$M����a0D�ԫ�H�~�(@A���-uԨ�c�	.D�̠`�A�N���� �OYNp�+D��B���;������#("��'D��f$
�m�����i¶8b����l'D�p�7ˆ�T?�9�i߉$��i	&D�ثd�73��QClޖ@P�aB
/D�H��ȗ'���Jȥ#`�Mc��?D�C���n�$�Q��'nd����?D���@�^<.|Z���!t�X���=D��旕aô�'�<����;D�Hk�*�%	���K4D-D����I��)�4�#�`K����`6j+D�$2�g1I��i0�.�7dJ�$�'D��Y����O0*)X��(U�Z)`b!D�|��i�q�za���uF2���$D�(���Q��=��#^	#G��:e�0D���,]%	3`E��/[��șr�I0D���s�|�N�C&�Y( �ޭ�	1D�yЪрW�U�Qc�3\Ͳ��)D�\�5C�C^��Gl�I��qiS�#D����C�'s�k�̖�g!Ƚ��5D���ţ
�
�8���@++����!/D���'L��IpǑ2/�-4L-D�8��Չq��c�JO+n�rA"3*ʓ�hO�ӈ@��Y�$L��d�G�rB�	�+$��"F�@1��lіf$B�)� r�QqHĿ\JJ}����;�� �"Ony��ٰY&,�e��2�g"O������(%�hc����4�c�"O�q�$׮"PHV85wn%YE�5�y��/>FNպ�釃0��tn(�y�(^�kz��k�Ç�%3R\I4DȻ�y�ԟv�T=��Z,s+����D�y�gM���
e M��ȉA2���y⨀"28�����DA"R&�y",���5��1��qsaGű�yb��(?5,�ҥ��T.s�ˊ��y�H�U��0C���ƌ��6�y��V�]�QHw��9GL�uX��Д�yõh�ڀg��3;�V�S!)�yB#,$� ��׌�-1<ܐ����y�O�x�z���2�8I2l�
[B������[��x�V��0Q�
B�I�<��}�	0D�����Kܵg��C�ɸU=T�U6��1J�����C�I%=m��9q*ı�P�/=4C�IR����ܯo%��Y��.+�hC�	&�.!1�g^y+�1���"�B�ɚ8��I��.O�}��/*��C�I�W�8w������w,J?*x�C��= ҉�ɖ��4�1k�9��C�ɀ��HI�S	�% ��F�vC�	c�x,&mNV����aj�W�$B䉧c�]�3�� j���P7� ��`B�	�a',xv�>|��4�#)�7&B�v�>-"��s��8A����5��C�əo���dĶ_P�u��'�7t�TB�	 H}�!�J 2n��� �E_�}�jC�	?B���#��>|��xP�ߥE�\C�I-���s`�7@Ġ#� �'�<C䉬w�`��f�3iTE�Ӣهo�2C䉫@��ht�B7&����[�&C�ɱ,U�!e��7c�PgŸn�C�'WK�qR�ѝ'&�و���)�|C�	:.���'�Ǣc
�����@�c�RC�	4����'f̤0˲��g�iRC��5t�%*'�ǁ�6=c4�ݻ6��C��:`�#�C]+1$Y ���-�nC�	�=1�I:����b�����[ �
C�	)������>mCaP�)�[f�B�+�:��e&�o�8��$epB�	��,�@h�*j��1��@5'B䉏M�F��vM�6.ڶ��0��?EB䉱 �f�ئO�^k|�T	^�<B��-@��`:1�%u8n!�Q�[:w+�B�	@F��A�H��(���$�C�I�"8Z�tI!�ʕ���U9M��B�I�wqX�����vm��Pb�ӈ��C�	�靖)��V�F��%:2��4k�nC䉦r��T�񋋟%�.��N�/>C�	,�V�
��OWHQ9�(�,vCdC��5]}�@��
!�Z���B�I�x�@����;z�)���1�B�=9���`��01*����	�n��B�9~�.����^u����B��>*VY���ԬG�ڭ@QiF�aN>B�I���A3bOǜ>d�Թ��H)��B�	/�HY#�KC(�v�eg�5X�C��'G�z��rc��z]f5ᴢP4e̔C�ɯ[K�q���\�r���$�1��C�)� d@�����JU��c��a�W"O��C"�[�<R�!�3�5`v"O(�`ٗ3��jR!@�/���"Oba�ք��Wt�3�aK���q"O�`Q�� PF�c�O]0I�-$"O�\�`H��NvD���n�(9�D"O�Y�(���P�GX����p�"O�����3I5�� �>G��У'"O$��Q�!��	e-N�֘(kC"O��B�6t�ش+����CW"O��hVa�J�R��k�;W��h�0"O��çh�X"5I�D�9�ڬ��"O���NBeb-CW��e��-�$"OB��T��(H�P5�$�[��ܐ"O�ʗ�$;� ���f��!"Or��a�Qd�)���<��yh�"Od!RR�Y#"^��eGʀ��ly"Ox�1R�׉Z�v�i�"�©:�"O�AH�����Jݡ�F��J���+�"O��#�ϗ.i"�-���Ɋ_BDpZ"O�����A��KTJ�D�P"4"O�A���R�m
�s��2-O�Q�5"OX����G�r����3�ލa�$�h�"O�H3���aV����U��@K�"O�]Qfn;R��� r��0"C"OP�Cś�vC�;���C��pt"O��#Q�K({�"��#��{ւm:�"O�����8�FѢIߺ��"Of����#W�\�Y���1m�r�"O<�G/�7�=� �V06k�Q��"O�Eh�iQ%1�꧄Y

L4���"O�)0�"�4��1�#��o�z0"O<Y�@��*>T(@ԫ�I:0��"O�չCg�Dd��C��.���"O���C������`��H.j�`P"OZ=�0eN�n��x;#�^��:H�a"O�e��L�e�rT�gI�PR��"O�-[Շ	�{K�52&ہ��"OD| �d+V8ɑ�%�=6�JA"O�k��I1��]@��j���� "O0�ˤ�V<^����2]�)�y�"Oz�KѫK5:��Y
�eڰ�@QR"O��XVJ�Ȭ�Ad�Z�*��"O��s�Ö�m��a�BN�c��B&"OH�ig��4�Ę��"�X��"Ob4��"o2�}K��Ж	�~p�"O|�cԪ3�D3�/K1ؘ� A"Ot}P�
\6>���54�B"Or1:T�߼��;S,�)u����"O�X�씎v���6l�-| ��z�"O�|�TR(�p��e'�BEba"OD�	�B�j�hQ���/<]�u�����D�F$k�i�f@f�n�ިI	�fܡ:�⇉r@Y`0��ٟ��I�gM�,!e��2HU�G�H4ECg�%��'4y֨�G��� ���?U$`%�V�G��E�S'�`B���2��$�HV#u��h���0�P�$_�6':�	���;����xR����?���p�OS�On��ِ�аw����s��)vB.1��{��'�ў$�'���Q���XEI4L
�vi*Ǔ7��h�O�ٳ�ۿo�X�&�_S�l�A!X=�M���?I�W�윛Cć��?���?����5�7P���4۟J�^����ޟP��*B� (p�xE��H5;{<Y Ǵ|��'�0�ψ��+�;f��\��B>����
V8)�"j�K�%��$0g��/�1���1w��K�Y<ⱋ�虘ND�ad��4q�7�Ky#�?�}����TmZ)|��QKr�ю�S��I�1�Ε�L>ɍ������(l� ��A,Ńg`�t�m���~b�'!�7��Ǧ�$��O~�I�O��(�!�<>9a�Eԁ4��%�Q��M�<����?I���?�E��^�'�?�a�0� Z�B��QV��o�=�N����I-2��d)�c�q��I�2nڅ/W�k�	!� ��u��[h�D�Ǯ�l�V�ä\8��0���&x�H�X��I�L��r%W�Q�����x�ʇ/ d!���ޗF2,K�$�+-{�}�����./��On��:��%T]Rc��R��d�<"����^؟�طF�A�&�(p��=�4�SMZ��S͛�/{�v�B��P�T�i�2�i-.�s���*{�f�#����xpr�b�O<���z�L���OT��:B����
��Ē�۲ř�g�L$�%b��2F�)Q�l{p���G퉩l"^�Q��	
<Gj�P3�ArH�4KE�l�@ɱjC�]��`��<r�!C`,̏+�ް�3�	:93L���O&9�'R�����=�X�5��9�
���?Q�����OqR�� �1�|��7cL�p�I���;��|��Dۍ>ɬ��c��Q�!S"`�;I��� ��iO�I>o� 9�ܴ�?i����A"?2P6-C�
C�H1K��yaE��/�r�����P�V��l�z�ّnv��zP"�|��ɠ~:Q(�x�읣���Nhlݙ�g�k�ɗ5��d�0��&eB;ݤA�y��)������f�s��J�#��m�A ��z?U�q�xr� ��?�@�i��7��O
�O?�I
qG��`+��:�d(P�ы26qO���,,O*��R�"*�H��g��1k��Z�B{���t�m��0o�V≺]�.d1 �eeά�al�O��l��i�'
���uϨ��b�'Yb�'���ƒ �M�^��B��!X�E8� �.h���Ů�մ����� 5N$�O+�d��[v�hI�?�d {��Μ%�T]b'b�$����2H)VP
h !MU�DA�8P����O!��Q�jj޽�r��S��$��S�C~��U(�E �6�}�0�$�_����Y��mZ!%�pɤa��F�A�)H�
�����hO�>=*�o&���͏�V�>IyU���d�	��MKU�i��'���'���L-�8�H����dZ�)ä:�$"�OL��  ��   +  �  i  2   �+  �7  �B  �M  }W  *b  6n  �t  ={  ��  ڇ  �  b�  ��  �  )�  k�  ��  �  1�  r�  ��  ��  ��  ��  �  c�    �
 8 �" 
. m5 �; �A �F  Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�� |d��"O
`�(�;���8���-0��1%"Oj4��ND^[��"3/9�0|H�"OB���H��*�ʞRy=a"O�味V�!X��!&F�:J�$���"O,��a
���C�Ą�M�"O,$3%o�-���p���+Ն�:1"O��ݢ1����`���y14]2��i�<�6��{_���c�H�`�fX�$Kn�<��A̼VI�xR[�)�Ć�pඤ�ȓA5��('nߡ4�� �)˩%� ���,��r�؊b#`T�eT09���ȓ!�b��g��}�8�F��-? �ȓ
K|m�ș�VṔ���2�%�ȓ"R�X�j�4JN�1�˘X�i����̹	_�jZ��1!g��zܶ��ȓgil,*�J�
j�Ne��i�J%b���f	�(U��:���G��$Y^م�~r�� S�%T"���k\�jx�ȓ|4�1�îJb��@ӵ�ݩn�V��/[`�"�v4�R�!ʎ<��M�ȓ`:��z�ؚh�J�Z��$HY:	��H��p�m�C1��!��B:��0��EnjZA V;9����J[
2���	��4'J�EA�IVW&��~�(aZ��ӹ�>� o�Y�|�ȓ�f�A�
Ο7�H��M�$�����mޠP����/���ANXo*�ȓTv�����{ ��-7�*h��I��sB�8�8���3����ȓNe*M�悡;������X�o��!�ȓ'lj�#F�m�+R&;�|��2)n�C��0S4���T:
b���:�0!��e֊��)��ͷV��,�ȓ0�&�8#���� ع�L�����;�P�AFd���,w�6d��u�H�,�fo�5�%���9#n�23�+D�t3��-�(�K�
�f]�f�)�	�iwQ����,K��4QhQ
QF	+-��A�!"O,��r-ӋQ
HzP�B$;6n�b�A"�S��y"�L�"�4�! ��;'ľ�0���6�y2�M%���1M�(�� �֣�yN��{'��
W��j��h�ٹ�y���_�2�c�T�@�x�g@;�y㇙M|H�-�ب'KG,���/�O��q&g���F8���	�t�)�"OR���%��<b�!�e�D���YPP"Oh!��̴w#H���H�r�Q3ROf�$Y�j9З&��Hp�f��G�P�����ԣ<ɉ�d�3�T9�S�&��R�ĦJr�|��x�{��Q��X�6x�D#�	���Jx���`ڲ)�:):Q� ����G�,ʓ�'�rg�|�ҊȽ7�2�Iu��=??����)Q�<QK��t cA�U�u�¸8�$�c�2.F�<%>1�7�8/��U
���N�SO-D����=!������	Bl���m�'��E�,O��{��yM�݋�c]�_g�M�"OB�Ϟ�V�H@�&aS=N�e��'�d��D܈PnNU�A����q�e1*a|B�|��[5�������k����#�y�AN/u�̵��A�0e���YQ�N��'O"#=���a
S�Ar�\��@3a�^�2"O� �<a��� ʖL7EҁsM$���Qx�@sW�C4,D���
n�r����?�O:�'�21�Q��F��QH�>���1gO���B�08��(PC�> q�!�5�IL����ҁ(r��Q����K��0V&x��{¿iE��[��i�RԔJ��7U&�FxҰi�ax"��:>�-�ê�<;�^]�p���O���|��E�v%ؙS��1�����ݟ�kg�'�z�� �[&=weZ�R0�۴2Bc��9���i��k�
z�0�F�Z��u�
�'#�p��EӁtd�YcϕD�FX�O����A�mz�E��,��e��`��8!�^�:����(��ͽm��b'��L�<�Sa�";����Š���1k�N�<�r`�)9H�\r3`׵u�������<)fjߴ`�b��ɜ+(5���	Q�<�u��e*|�v؞<M�%�惁J�<Q�a��9�<]��I@�`Q�)EG�<��
4,�����9��q@1KF�<!#'ɒ*ڴ���"�5�8G���1�O���JH�pd��A�
�l-C�"O�����--�|�`C�'`��x�"OVк��3=�LepE%��VD�A"Oh��]�[��X�N+�4+6=O��dޞ $��� �-��+¬Q1a|� �|�Dܘ~��k��<4�`�Q��O-!��8n�x}S�ӣU�$��b�0_����>�Bj�(	x�Q�&�7%f�885@�zx�(�'Q�-	�ٱQ��9��"@)U�5��'���2��N�[�����zvfģ
�'�0`���ڳ\~I��mZl�a�'�D%�-�e�zxru�el�t�'$䀲��}�4��]�J`�m��'��!  O�EI�1A 5s�͒�'@�UIG,�\����_�]����'� �gڟ���3�*Q%$��	�'�x]�'��^ȄY�F�8H�2���'�u�4���6��������'J���#Ri�
���ŲtV��*�'0����T�#�H�h��i;����'w��r�����!����c���s�'v8�
b�H*$D�&՚i�z�Ɉ}��)�	܈v�n�{����Rk��H!D!��D~��ٔ�" ���1rg�;K]�ODM�Iv��i�OV�1*������=&V�D+5�$�g�5v>���O1!^��%*�2�8ȅēt1*VM]'<nu���,!ԡ��JqX�zU��~(�A�#��2�A��	S���T���l��)#�S�T�����h��!��z<�݆r�m�ȓ2�n��d��[��Hjg��PY\uEy��'0��T��8��{c�	�&�a��'p6\�'%�A
��;�eƇ0"�Lbߴ�Px���N' X�O 2M�L�3��5�y
ͽ�mY�_�o�x0��K����0>��̕2-���eߘK���+$�{��+�S�'i�l<�t�W�0_�c��Ƹ\-���(�� �U��:�j]�u_�Z���ȓt��xxrF�NJ�؛�\�}ոe���?��n�^ r��灃%N����s��r쓾hO�O���"��<~Ԉ�ia疨h�@�Ó��'C���s�\��g�)�⑮�c��'���q�D#|�'w���L������Q�s�P1��D9�'{o0��"̅�~&r��C5F�Z1nO(<� �M9P�ۙj|"�3�.H}X�`�d�O�EEz���Zvf�H5�>G�:͒'&���!�dٲ!B��9V��ֵ �����Ir)�!iA�)��R}$,a�2�S�@y���!	���Ȧp4Q�����@"� n`�C٦����,���f,-`t {C��R��G�?On��*OD�Ӥ�1*��Be��A{Re	#E���1��	�0<�'��*R�vS5� .��`s�E[��hO�O�D�#ܕ=��� �%^��ȡ�'��r-��(�0�D%�a(�( �+�
�0>a՟xBA#��	vk�I6�q۵C��yR��/:Lh�ؚ֤HQ@�6���y"�K9�p5��!�ݢY�5��6�y��T��p��P"KpR4�e���y��
)=�z����<�(�x�e
��y��ȅDQx��_2l�Ht��	�x��'��e�P�\1	���7f���'|X�h"�Q���@A" X��Ó�hOF�X�d˧" �k�c������"O�`j��V=\���SQ�
`��}�`��8G{��IFmƄȠ�(4�x����Tub!�$ݿ#D9�V�R.B�Rn�#_X!�D���q�#5T;�5��.�-G!�$D8�&���(Ӝ";��h��E�u3!򄇳_=d�2d��e.&�[Ҁ-
�!���1�R����X&*mpE`��!�Q���Iu�k �hb�@�*�!�)v���ۖ�<��Zs��!�!�B�,]����s��D@���Py�*�t�	Ä��|v��7j�/�y�*E�-D><ᱧ]�l����'�y"�I92m�U�'�v��7d@�y2d�y�� �gn@8F��!�yl�9M�pȸ�"^�Y�n��򩓉�yr*�,`Z���¬f� �ƍ�y�&5��u�4<]����PJJ)�y�����b�ڃ
Ɯӥ!ߕ��B�-+O�W-J$͐5F��`�2=�'�Pa�"�޻?��T���@�i�0��'�`���ַ������"Z�&���'a�� ���T�'E��K��}
�'J�4#Չٙ}-����܈J�U��'�d03��[Z���)�=�^|��'����0Y�pʕ�0ZM��'�\��1X����KU"sẴ�
�'F&a��P�|�A���֪h>4r�'`��;��)�4��w);\)0�'�hz�#Z�U�p�C��źi�����'Vr9@7�Zu1�)�5� �`��(0	�'N&����BO��1E�^iGl�	�'�������a��E�TI%Z�&��'yj�&�1Liv4�P�O�=,��z�'r�)����=���ЍAH®u��'��Q!�eVg�pL	�S278t���'�d�G� .�p�RV�4z��U��'_j�*U	
XH)��Pr;���	�'h�a��e/nb�%�YU��	�'Z���CH,����C�P����'oր�)^"e� �	���\tJ�Z�'E�Q����n��0��Z�>���'��Qy��g��1iǮ�A�V@Z�'�r�`����lL2$�D�3����'�)��J5F_�E�sꀘS�V��'�4�0g�5z�cTō�C#��s��� :(� �DN����'�U��P�"OL=����3x�T�e����]�7"O6�q���!F ! �$v�t�0"OfX��@�wJ�TC.�4m �BU"OP���!�~sn�Q"�u��<��'�'���'��'O2�'���'chD��T7-XBe�n��`�����'Or�'I��'���'��'d��'�U���c��X9v@I.6��Qt�'t��'\��'���'���'�b�'3������:iΠ�U%��ۂ-���'���'mr�'���'["�'���'� �����႒�W#��Yp�'���'��'���'�b�'�R�'�"!���<sxa���L onl��'$�'B�'���'F�'_��'�D,����gĜ<&x�Ӕ�'%
"�'{��'���'��'=b�'^"⓯J��2��* K��5+�HR�'v��'���'�B�'��'$B��/����n�"�-���n���'�"�'��'(�'�R�']2b�Dn8ź��\��̓�b¶`b�'1��',R�'t��'�2�'h�'�[���9Èź<�<�d�I�z"�'���'��'���'���'p��+{ʁ�g�� �$h�#�H	mB�'g��'���'a��'���'�&Ɵp�\��W�T�N�YCOP�M�R�'��'���'���'tL6��O���)fą�Ĝ�Aʮ$:D�& ��''�X�b>1�'�b6-�3DX�
�)%L�3�ʓ�w�9C����A�4�?�N>��_�<oZ�sP�t�S �C��px��"9�>E3�4�?�E�&N���'��T��FЬ�����<����*+�����B�+�n�����Olʓ�h���C#��<beA�!��e+���b��?��?�&?�������Өd# ��Ɓ�&A��ZS���}�"�i���<%?�B���	�sz��v�N��Ĥq�H�8�`�	8j���Q�Fe�$lE{�Or��t��x�HM�
���`@��ybP��'�P9޴_j��<QEݔN�2%	�C^��&�A$נ�?�L>q�P�`�IϦ���䊎��\��ٓ9+�P;��S%��ɵ'�X x��2H�b>uI���3J8�X�I�Pq��*	�vBD$+1d�2ʜ0�'m�I��"~��\ٲ��\*gY�	!k߃O�@͓r0��/K�����撚���i>ՠ AR�gFI�t]�5��W?q���M�����0SBC~2��H��iY�I�:�)v�M�:�@s`
�9�0I��l]�XD>9S%@/1��̳������E(�f�%aj$��3�`�poZ�DFP�Ri�%��!��,4�ju��C*��0��l��Ƒ��-U�u.���l	�	����p�& �:��&@$B�SJ��n�0̣7��%��D�8g��@HfA�pWd �b�ۊkT��g��~�xT���12�}؇G�6{M�e�c\3��͒ނ�?�@+cVkO.�P`�7c�^�#�	�x%N��7fW�H�ӧ���+&���gQw��qiW/H%�0���ܢﰕ����J�vX����x��Q�4�?Y���?���_)��@��Y$Mʂ	Č B���J7m�O���M'hF�D�O���O����Oj���HD$�.��Ӿ^ԑU�i�<��'�"�'�B�O,�'�S5*J��
C��6�0trR��O�΍��4Z�r5!�/�y�S�'�?��Aa^���J�kF��:���#K���sV�iu"]���O�����uy��'��$��<޺�ON�N:p�9GKC��%�<ɧg��<V���(������	o=��q�`�'�������h����4�?WĔ��?	��������'��qTO�*�:|����r�D �4l���d�5(pm0�=O>���O����O����O��K�.�A�NE��C�] 6NPW����O8ʓ�?�H>A��?Y�2)�ʴ���1���;���ya��j�F�T~�'���'�r�'���'�ڴA&
&9�.��A��|���1�m�L˓�?�L>���?�%�_�$�l5z�5`"L�y�`:E ����?I��?����?q�͸�?����~b�T�u��{���:6���i�M���䓌?����}�0��a≏,�@���[�@{�dذI7h�t6M�O�D�<��"C��O����5&�#=�����0ݸx���M�*O*���O��"�S�?7m��ֆ����ӔV�pd��	]�z>��U���!�?�M��S?����?]��O&��q቎/1���j�]��Dz�i;��'�Ґ�[��ן��3�D�X�2���� H����%-�#r;���/_��6M�Ot���O���R�i>ij�N�?`̘I+R��X͙2a�͟[��ty"�'4��Ϙ'X�+P��@EC�`Vb ���96wT6�O��D�OT��SJ�i>��I��@Ս�@ĉG
�:�2T�d����O���\c�1O����O
��K�f���2F㚨#�OH!L� n�ݟ�j^����|���?*O��k$Ɍ($<4�!ĎD�Ggh�� $ۦ���1ڌc�0�I����Imy"�$� y ��2;�N��EO�;��r�d0���OB�d�O���?�8�Vx1�֛1�����,�H��d&�O̓�?)��?A(O�9@#N�|ZEΑ�(ՌdkV+�3oq�)����_}"�'��'���Пd�ɕr52�]H|�!hO�+5%��.]2a�'sr�'/�Y�tK��R��ħb��Qm�<��$+m
�y[D���i|��'D����I�Tc?�ӄƐH�9��غ#I�$)D�q�D�d�O�ʓm��)T����'�\c�`����K���E�@�.T��L<)O�1�j� 2�� �ܤ4��,RT�!�A▹i�		@@,qz�4J���ڟ�����_C�ڧ9� �#ȉ<D����'a�h�6y�)��g��+��9��ʐ$֐`ҧ�+{�6-��te(\m�۟��	ßt�?���|�6F�X	x�z g�MO��BV(գ]���@�^�I�����?c�D�I��� ��H'	��$B��ȁ4�.�Bܴ�?���?�g�! ����$�'B�؝K�،Z�*�7FYcF��>���?���Rؔ��<����?��@lxt�)A<M�3狛1����W�i�b�A�a��O���O0�D�<��&� |�� �2�	1vf��x�W�f%���'�B��y"�'��'.�	cݤ���+�La�HQr*]=)��:�O�!���?���?i/O&�$|�$�⠗�?�}!Á�[�bt9Ɔ�7^A1O0��O��$�<��6����Ϩ8;lX�#L�u������؟��ݟ��'br�'�~���:�BU�P�b~‚�%�?��:�]���Iן��'��g�Xr�˟�*�� �$��T�K��*�u��II��M+����'$�o��a�Tq8I<Q�O�}�f$��OS�IƖ��CJ��%��Iy��'q���W>M�I��S�8���$,�y��}I�D*�ȋ}B�'Ǝ�h`�M������f�ġ���X	9Yq���Hh�	Ɵ��"J��I�@�I�?���uGAM���1p&�>%|�Ĵ����O���L��H�1O��>�P��Ƽ�4���.g�ةX&�i9�L'�'br�'�R�O�i>)�	!M���n�A��pI�3q��ٴS��8�Ç�g�S�Oh��ϕh>PuZ'��0�!z��6kpN6�O�ʓv��+O��O�$��d�dIܿh嶵[%�`���慞���'�ja�j!���O2�$���)�c����I['wcT�)��r�r��W�z� ʓ�?����?��{rg��P0�U5�˨G=Xk��I���$[������O ��O����O��%"�d�aGu�c����J(f�(N����O(���O�⟔�I�x�ժ�N�g� �� �x^�Z�̓e:��?�����O��!�+�?MI!�(~�-07Hñ��}��Ek�����O��d5����(�MʨR��7m��4�D]��	ɐo���T��_F��ݟ�Imy��'�`���]>��Ix4 tH�d�* ���2[x���4�?���'�v��棅���O�� �2�C�z��c��k��l�֟�'
��K.Et�AyR�OeL�,W�g�f����ۢt�A����'uRgP�>�h��y��:����C5�)Q��+�X�XP��	<d�p�����㟰��DyZw%�����J�AY\���遜p�x�OX����N*� ��<�~"�g·6�@��F��4.��s�������Ο�Iߟt�I�?������'\K�d� ѻ�E�U��;$6�Ȁcf�ف���Pz`�3s{ʀ�-��8���ҥ�-�M���?�����(-O�i�O���������  �(�%G���D玐��'�`�g1���O�����4��� X7��j�≃O�6���mn�B�d�N�x��?I��?a�{"N�R�0�s��RȮQ�C�����W�
m����L�	៤�'#��{��ۢ�_�L�X��@��m�u:Z���Iɟ0�Il���?A�S�ho~I��㇜QuFeļ0�l�p	H[~��'y�Q�����Ɓ��r⼬��J�13�i��܍.&Hn�՟������?q��J�P��FCǦ%���/K\�8H��.T*�2F�cӘ��OZ��OJ�PvR�y��?a��eWf4��3&�\�Th\�;�	�d�i���d�O�P�E�Ɖ'�(uy�!�9C�T:3��$���۴�?�.On�$��i���'�?����j�N� R���֩�=r�ԩ�B�$c�O���Т\���Y��T?婆�11��(@�˔$������>���z�d���?	���?I�����q�� �h����d���OLBL�TZ�@�I�|�恙�5�)�� ]�^(�166����C͔#� 6͙V����On��
+O���O��`��_�` �B�J�����HYԦu���׳[��c�"|*�NP0(
QE�7B�Aq�#>Ȧ�%�ib�'����i>=�I����B13�b�G:Z�0�M�+������d'�&=���?��?)��?�;rK\LS��@*v���$Jx`�o�ʟ��fJ�Jy��'/��':qO���*R�(=^�*R��17���T��C�L�y8�I���~y2�'�P�`�P!��I�
ű6�ܩЊ./�I���	���?i�>KS�4��+��P��˝3vdi�d�??���?�(O���M�>�S�]ql�fkՕNpX8h /Ɓ/1�6�Oj�$�O��@�ə7�8��hӆ|ږ���+����!!Y �b�V���I��ؗ'�2"�7>�S�t˔�� �X�Bⓛ~�b�<�M����'V��^�R�\AL<�p�F��F�XT*A�4@�B��צ���yy�'l���@S>�I���S�jj�� T�[�,\Y�#��P�,Q�}2�' ҅�쏂Ϙ��i�H[��;��ژv�61��H.�����C͟h�I����?���u���T@��P��<�s�ޔ���O*tq � 
1O��ڍcuC�-4���'��H<��5�i�h5:5�'���'�"�Ob�i>��ɠntJ��^�����C�-+��jٴH$�Y�4C�S�O�R*1� �����;K~�q�J�D���A�i���'2"��$�i>=��П���
:n5���-r5�f�/>��SW�CT.)$>Y�	ןt��G?� ���V�Lt� ��~U��o�ٟ�! �KFy��'o��'	qO�IX�o�]���p��Y#�5:�]�d0�J^9L ������������ly�-��y�)¥IB ��eA*��ڀV�,��؟x�	^���?YQ`]�n�� �H�<Z��]�e�T�Ș���Gr~�'%W��������������#HD��Ra	'�.y��
�4�?Y���?Q���'4�(��Þ�M3��L6P:�e�-sB�����I}B�'��'�r�'Y�P���vӈ���O�d�6E��!u|=Kb�Q9Cq����m���$�I_y��'�Vli�Ozb�O8!Ԅ�qO�1�B�0j( �!�i���'_�'[����i�����O����(5�r N?bOJ]kb )�xւ/m��'Z�Iϟ���Oj>m%��s��)Z�#�R�R���f�)IZ~�kG�i�R�'���u%kӸ�D�OZ�$��^���O(�ФAмO�\��e'ҔK�V)���Z}��'��"��'~�'PI�O*�|��@��̶M��))a)�"?�ވm��f�~��޴�?I���?Q�'�2���?q��u(���͇�}��9�W�ܕpt�D �i��£�'�ɧ������'���*��.8(:Ĭ��[��y� i�2��O���5��-mƟ��I������֝$��Ԩ�.�8X��U��f�6��O�˓$^h8�S�t�'}B�'������dQv�"��$$�XBtO}�r����1��	nZɟ�	̟��1��ɿ���a�m�zT�!�ӇK6>��1�>��K�<����?	���?����?��&��b�ƕ.��db���sx�1�)Jm���'2�'XB��~*/O���ߛ7eUa��	
0k@@��aܸ�!�3Op�D�O�U�1B�O^�$�O6�$�3h�mZ�*RXjQ�D�C��Ի��Ո�6���4�?!��?����?�,O*�я=c���!c!N3gb򭁒)�>4�zǵie���Jg��'��2xB¥�i}b�'l,LZP��<0ƨ�� ._�H�j�ehӨ��O��<���_�&�'���|DI�  um�\��� ��6��Ot���O��$Z�>&�lZߟ��	ٟ���:�ǀ:G4<�(��"��4�?�(O4�䛇~r���O���\2;��i�>�7�PY� ���QҼ�yڴ�?�syR��i ��'+��Or��'���be�B�Z�@��4JE`�>���U#h]q�����|rH?���`O1+�VD��,XPٕb��xg$ʦ]�	ԟ�i��]�?Y��� �ɍ=^�+�(���l���>Hn�޴iŶ����?�/O�i;���O��*����j��g.1o��u�@����������0<;h��ݴ�?���?��?��A�.��柤\� $@ũY\�`m�ş��'t�8����i�O���?Q��ßs��aM��H�Eaj�����g%\$lZğ��I۟|�����ɣ����D��<�����iK"h�pp�>bi�X~��'p��'��^�tx��Ȑ9P��{fg�1�K�
�D��Te\}P��	jy�'n"�'�
�3�LՓ2x4����wJx�Tg�y�P���IןT�IByXG� ��=s�T��㛱RT4��5c׀f�.7m�<����D�O|���O(�k�8O�tqW�I9T��`��Y7Qq���u������柸�'�0Ё0��~2�Jv�Y!�L"r>P��7=0���iJrU����ş,�	�P�`�Z�ܴH����@��8��gε��mZП��Iǟ��	*N�8"ܴ�?���?��';��i�����Ѕ�a�V�[��!#�i�B\���I `"���Ԕ��ܴHq���Ǯ�*,h,)G#M�=0,�mZ����IW�H�2�4�?���?i�������6�;�hǋ
�4M�](I��	&l�	ş,sքC�,�Iyy�O��')�0�i �EwJ��@&�{zImZN*��uӮ��Oj�$�0���O,���O@�B��s����Bh�*���dG�Ӧ�
P%��$�	Py�O��O;rO]("{��h(ØKYH�҆�G�F�6��O�$�OhթCЦy��ߟ`�I۟4�i�mkl�	(8�g�-U�졙��dӆ�O�8�D<O��� ����"E�h�t��dޱ^���j �M[�h܌�a�x��'��|Zc�PR�M�]�����DX�Q�܌Z�OH�%h�O���?���?�+O0`S!,�[�ꅈ�l�1t�Cw�� ��%�,�	���'�(�I�����J
e����ͅe�2\9�|����IZy"�'>�'h�>���۟O�,�z�.�)�8�J��Ns��ʫO����O��O����O�Su��Od=p^&(��	�*\�ʽ2րZ}��'���'���mAM|�W�'f�a�gV�
8b˃�Ec�6�'|�'�"�'�����'F�<�l���"Q���5�)&�vn�����Sy"×f^������L��uF2����q�$Mʕc�Q���L�	Q�
�G�~���O8Px8�@"�54�� ,~r6�<��ĉ�-��& �~j�����xa�)L�n\���3��A�� D�c�0���O���y�|"��ߔ(�B�rdD+�l�clC()�����K��6�O����Oh�i�Q��ԟT�F.�I��E���8s<�}�Ţװ�MU`��<9O>���d�'�&aR��*"�����G�ؑ�R`|Ӻ�$�O`���!F���>���~R a��ց�H.p5��ͽ�MH>a��{͉O��'����U�1nʠ�%[��|����'��-:����i���|Zc�*w��]A�FbQ�x�O<y17;Od��?����?�)O(� �-��H�i{>�rb��^ݖH&�F��'���'��'���'X��@`�C�|�`�̓�|�>}R3MP4�y^���I����	xy�F.=;�.XXH@ LN�)t	�D�\~�O��=�d�O��d ����vY�J�	;	�,q"�3���'K��'P�U� �A���ħ?�F,��#�&]�P}jA�:��衽i���|��'���#�y"�>�,�$^��� ��9o5
,K���ۦ�������	���"S#����I�����?eB�˴n�p ive	�='p�����ē�?��4�T�`!"�q�S��+�2~�~q�(@����2�BY��M[.OԽ:nL�1ɫ�<���6�'N����h� `p�Y�!J�Y�m0K<�FA�����L<�g�(�T�vᚬ1^�juGQ֦IY��՟8��Jy��OD�Ky�	��܉	�'[�X�lt"3f &��6M��vj�����S���sGL��;C��3Ir��!d"�M;���?i�� ���ӕx��' �O�â	�>O�*�H"#��)�e���=	r1O���O�$��	��uA��
[��Xp6����oZ���I���ē�?�����kC�.p�b|�`�X1�(1ۡ�l}�ٞ��'���'�RY�H����,:e@x�茀j�d����\�M�,,�K<���?�J>����?i�oU3���w�ŗB���d���X��<���?������ x��ΧQ��"p�$[:6�jG!�;D��m�'���'a�'���'[T�b�O�ZFJ�5Oc�-��O[?�q7Y�x�I꟨��{y"�պM|����b�m��,���J�8PЙ#��)��a�I��,�Iz�b� �ㅁ1c�`C�L�=} A"��b�<���O�˓�\�������'��䄁tafu�HCH,�	eJ´#�(OZ���ODh�R�~�҂ăX�6�%!G(��`�R�K����'�"�Q�lsӄ��O���O50�)\v�#c�X�j:tA11��%p�o����^."<�~�1Eʇ�D�k�/s��U�����y�����M����?���B �x�'>(�$�,μ DE��m(VmyӮ1���)§�?�����OҒ�8t�ڴBmV���˗ ���'�b�'��`2��4��O�������X*�$ �,����a(@�4�	�a'b�8����h�	b@J!�f��q���[#�ɕ���۴�?A��X�h�'���'ɧ5�� y<dI�@�(&�4�j�������I�1O����Oz�$�<qB,�/�8�
�c�(O��w�T�r�0:5�xR�'�r�|B�'��$�<�>���B_��$1v��>k b}ىyr�'B2�'��ɾ݌���OZ�Ւ�
��H�t풬�F����O��d?�$�O���!���!i�~�G��|'h��#�7MyH��?���?�+Op�P���m�S�_5�h���3�bP:T�G/�L�ܴ�?�N>���?%��]�Xo����k�!4�FHS�'Ş��oZ�����Hyr���?'��T�d埾�3��n8	NƯg7�V�!l��'3��'�8���T?�򷏋�4�^���
�B^MR��z��˓��$�ĺiY��'�?��'7����A����⋛�(�J��VTr7�O~�$K�b?{ '#z��PB�O=��h�&�u���PE�F�����D�	�?=�O<������F�G֊�a�V�rY�`�i���ۍ��˟�ysȀv�zͳ卝�U�~��#L��M���?��"�,�	��x��'%�O��	.��u��ś��I²����1O,���O���G�Fmz�l?R�r�ၬ�j[�m�<�!h^0���?q������4��-F渁���TK��уZ}��X���'_��'�"�'�"���,�h-+!�Cd�y����%2��KX���'��|��'����v��Wh����Sq�}���i(PI��O2��Ob�ĵ<���-l�٨&~�����b�h) 䏢S��	����Iş��?	C�k���-"8�L���P4(BfJ���D�O��d�O����O�@C��|��ZD�;!jC!@ٳFV�u5�����iFb�|r�'G�	!JM�Ori��睍^X����^�z��[�iNb�'��V����K|����j�ǃ�A�����`�>q�I�OO�MJ�'}��'L�����T?���D;db� ��-��Q��sӔ�ct ��A�i�>�'�?Q�'d����f�"LJF.�2�^51a��y(7M�O��D�75T�b?���C��{Ʈ� c��B�|�
{�b�u�զ��I�I�?�J<Y�>
��{�B�]�P�8$��QX"�iS������ɟhr�܁"��� 퀸8�@`#r����M����?Q�ݾq�*OBʧ�?y�'9�DX���'zFrUJ3�M!1Ũe�?��KRr��?���?����(M�j(���ݔ
ID)��K=<���'p�%r�'�⇧~�����M�2XS6F�	l�~����J�� �x.����O(�$�O.�?���$&ʐ4\R�{S�<sq��; �U�1a�'�r�'s��10k�;chU�=�Qp�*ؗ��']�'���'�������D��
��1�n�0��ϑd���X�L��u�	��H�'6�h�ڴ �ḍ@�E�}+�F�t�]�'�r�'bX�p�ժ�ħ�� �#��(6�2T�%���N�r'�i�|��'�R�߈��'�`[�L��v�u�;E��3�4�?����$��c V�$>��I�?M[QM k�d�"�]�؅cs����?�s���Dx���� �j���������-�,X���i��I�0�Ne��43���˟d�S����ݜ;��U����}��H)�=��f�'Xr��O����Aþc!p�b-�-���q�i�P�XFd���D�Op�D�0�$����r>�4�؀��%*&b̲Td �4P� Gx��)�O(	2`�94F��8��;��4���X���������I�`����N<���?q�'��=���IE�*��T&Xh��}2I[���'���'M�d �V�Tرd
���<|h��X� 7�O�����Or��d�4�'��'�T�(�P.���H@�TXh1��>�2�@k̓�?!��?���?��c��P� ����XQu��7Hz���.OJʓ�?!N>Y��~� ������vm̤�υ�M���A~b�'F�'f�I�0�|���O褨8����-IP���T���I����	h��6>��O�'��2 Y�F��s�T2�O���O����OH����(˧�?9.K�4.�ʧ�H,f��y��5Y+���'��'��P��ȱ $��X'j��)���%���Z���Rx�K�/�,���̖1�yb�BЂ�:�xy�&
�1-���M+D�(a��]#�����Z�ئ&\"��P��Bi���D��P~�u���S>�����݋
\I�$$Y(���saYH�v��!��3��q�í�� c~u`���"v����l�7�r���gT |��J���%4�^�B���K,�����+��)ys�^,���'�Yj��.Q	k01 �T���؟��	ԟP�	��u�<2���;��
�T넜�3
�6n�@K!jP�C�f�h�N�������|h�� 'j�8`�C��D��r$%{�
�b`dە���0�ꐯ".<"E�I3.�賞w� xPO�>��]!�/U��0��'���+6�4��=AƄ��J�:58� :<E��1R[o�<!v�M�K̂�RreD�^��$�<���Z�����'�|��B�)H���",��䙫h��HϺ �d�'���'�2Bb������<Χ]�ʡ��!	}'v$�2H��#~�EeI�irҜ�t`+�f�	ϓA:����]�F��4�"3p ��������KT�F��
 ���<�C���uю���̓y~���e|\��aV*�ΐx�^^<>�X���?)���,�I8m�:�{2"A%R5�"DfZ�D"O���nF|a���Y��
�����x}B]�l���O��M���?�v���g��D:W�X-O`QB�T?�?����R!���?�O�n��)#�Q`c�"p&,�8"�3U����e]�Nk�{��*��Pȼ�X��L��M�aE�'�a`3��3(2aHĖY�R-"�M�6�( ���?��x�	,�MˡX�1@�L�Y��m�4_�5�Q��#{�<����?E�Ĥݜt�ACpKT!Ggz%��ω�O4�=ͧY�����e���@V���#^�_�"]�Љ��M���?*�J�k'��O�0��z�:i���<wr��`���O���х\��Qr�A��P����E�H���'��)ע4K�ᨰ����V���}�qb5�G�1e8\S�C�(p�e��� ƻ4[��*2bK�����e�FW�$��fLGv�$�d�O�����'4LJ((�.�.�zA�|դ-Y��?!���?	�FGt̰�E��n���ΈC��؄�I��HO�x���T;Z1��dɠ9�p3�
�����	Ɵx�		i���ȣ�����ʟ��	��u�O)L���Ѵ-#��%)���x04B��E�y���D��Kc�����|��T�L@���30bYi� ҵJ���a���(��D\�?c���L>�a+\�_d�A�L�pD��o��?��O 툠���$�'��Ofid!߶X�����9E��J�"O %�vW�I~x�D!�}��=�矟���D�A}�X�(E㈞p� �"V�6��l���ɞ#��������ٟ����uw�'tb0�(�ʣ�2�Xq�R1{�A��= U��b��=4��5XP�-<O ��;7��J�DO�K��IP" 0��	r�FD�/64��-<O�r�$��]�|kW��)!��1�O�K��'�2��2��qWiÝ5�)��ڽ_�hB�	5������4 �j�2oTV�c�xɪO&�E���q�U���	y����g�X�;tP�`���Q���˟4J@��˟����|BU���2h
 Q��O7"%��4p2��sl=P�	�@T�n�a���XhFy��	�8<�xq�FP�Z���z��i���4N�~���C3�[�91��q�f<����I���'��	9ZZ 蹱�D�=��P��U�\��c���Xx��XЯަ1,P�k0�&`���h��3���4hDv��s����,X6j��%��<�(OdT��g���i��ҟ�O��	��'�:�9,R<D��}ऩ  -=B(Ӣ�'���՚~�ƀ��%����H��%D��O�Dٱa褍	���?>������ ��	�F�}�qg qXD�CU
�'f�T��g��h����
�Y.��+&�=�'�^Б����'�������� \dz����`[�%��g{�����O��D�O��$>��6g`sFM,L�M�t�"�yg��j�P��O.�q���Ԫ!D��
,c�����3�.�M���?��G�6PJ�E��?���?���Z!��5�9���)5y̂�iӳ��[R	\	%ٺ�[� �I� )��7�s����r��RgB��5,LPc�[�l	���12@M��:s�Y���M�J����4��i�ZUj�8O��z�-(�\DR��O�� �)���-O�tB4���t�O!�O�Qcs��6De"i렦��[x�ʥ"O.�S�͝7�
QZ��/W'���8O��D�Z�'�7��O�ʓu�P�{O�RrHUB%��>�>%�bM:%JIA���?i���?_?Q�I�|�3��2�e���V���8�nU8�0���M�j-�8J��(���d�Z����D�Q(h<x�4eT:ZfX=4�>Q�m���G"?��#6 �A�>|:6�OǴa36�/+^�
T�U�o����G�O��d�OZ��<�����'�F�C��1j�4�á�$en0"���;&� ; (M�>j~tA/�
$�`)�<)�iIBP��qdMʑ����O@�e�?;�`��gKO8d�e!$�O���]5E�����O"�ӫ
��2�	�!tHJၲ�_禡�H-5������%2�U�c�+OX��	/��h�#C1��,
C�O6a�������^��ԃ��8��eOE'K� S
y[�IO�z���O&˓N��9k�	�#2�(s��U� ��<�����<Y���Ba\$���J�u��
֩ZI<�q�i��=B�"_<_�)��U���]���'O�	(�e���u��ؕOM8��`�'�s�e�#&V�-��
��42�hJG�'<bd��W��y0���Bqx��عF(맙�iM�-�����&]��x���#w��m۞�����m�@9P$�,I��ԣ��d�ÊXb) ʘ��0������I1����Ox�����z��H��v�2��ąӦ5VqXw�D�ON��h&�9�e��Q������[�ax2#>ғp�\,���c2B��2
^9g��cw�i��'BQ�WE&1&�'�2�'��w�6T����}��c�kA�	>"�1��M�k��Lc�'G���Ʃ՘��?A�a���"A"gMW_9T9XP�6����M�.dˀ�-�3���F��	�ֳ���7 ���&c�ΨmZ�0��+П�>��?�U&���tR��Y�$iU��$��xbA���ڼ��M�A��t���DDq�'�t@�����0ob��h�R�j�#G�$�툄�OQ�4���O��d�O��;�?�����4��� 
��D�2 �  UK�My�%����x4��	��dŐB��?:�x	�F����|h%�L��5��jZM�Ը5Hݫ&�b)����w���$&�
����¦�(�4�?a*O��"�	�R;x�#�I̸/��zSG��C�.C�I*WON�h��PUF��R �J�D1 c�T��ODʓ[D�T�B������O(��*ZXr0�O&��I*p��O\�$Ѽ0����O����>3m�
��:��oډW�5��B
�Slz��P�C� ���:O�%�� N=+�����W4Q��`9��'	ܚ�1�$��Ct��h��ū�W������-�D�.RmӜ�l��8�rf�v�آ�A�EC�����qy"�'��O>��Ǉ�:.�!�u��V1���4?�,O�=��UǛ���O��\�n^�90(	��D�Jc6m�Ot�o�w`�H#��R؟X�	ߟL�� �0����R����Q#X�	���A�e�4�'S�
ղ��!HC�S�{��-�0K�R��P�T�_;�}����,^0��Ǝ��I 6r�p�+� ;�*�T�ۺ[�t�` �)�0Fc|,�k	�[wD\���i�'��T�	8�MK�i?�)Z�/ق$#��P��"��DFR.1*1O�4<O����� ��l[�=V���+��|���	�|���eg�*%(��90�$=Hʷ�����ɱifBŰ�(�Y�(��fщtuB�ɤupRD�˄�f���OS�E�C�ɸ*�~U���h!��@nQ#@�C�I*2�ֱu��%�豓4�N jLB�	
�9�VΖX�ʕ�5��JB�ɭ5�JBǉ�'0��("īF�k�pB�IQ�`p�_�D�bH��Ч
jB�	�-nRLӶ펷�lp�!O�-MC�I�c����r�3�F���Ѩ#2�B䉩�tc�d
;.Je������B�	 g2ɒ��yA A�*c֮B�ɆEh�ݠ��2~]$99�
ò-ȤB�Q�hp��gg����A�Ve�nB��1
���;F�,3���BT�
�C���xx��MN	N�@HӨ��y�B�)� ��+�I�yE$0j5��.*�`1۵"O>�����'�ޝ�4cQ-F�K�"OP-�%�Vpa��J�]t�<*v"O0�ن��,j��D�tB
{��,r"O�=��Ɗ 8�T�3�Y�j�XY�p"O�� I�'�l��];��]R�"O�����lw$�a&U;$Θ��s"O�8y��Zo���D�U�\x�"O���Մ�	g6���$<�
���"O��Ж��/j�!Qg���(��H�"ODlӖ鑖 W2U�f	�P��"Oi����b~��Qi!�DW��y⌓���r�6V�"! ��E�y��\�=�d��I�#Q�~yH��Q4�y�`Z�g����1�ى~9�A�M��y23s`,\:Ј˙g��� �5�ybB<(�z��e�b9��mĲ�y�k͍w�|-a�/K�!P��yb�FH�ĥ��D 'Q�����I��yrO6a�V5(��)A٬ +���#�p=�`B@kH
y����9X���DA���aZw��@��!o{�{��F�J��d�=:�P˗�-.(6�\ H�ڦi�B���D0\T1O���@��B��^�-�Y#P�x5�#A�& n�𳎞,Z�$�?����:2Di#���M�<@�0(") ��I=>h���JK�A�*1�*�""������l�'+�U�)����f ǵ�ȣ��O&Le�b[)(�p]��>�O��Y⢂)2�
, Ae��:��}A���e��OHq�IIiv���& �JNd��*C�`����I#e�2�k��I�n�IH�kʻ����v���p �"'�(Jj�F�=����O8��I�?��d>#��˶���iozEpD��K{��Y���qGL��!�o�1�L��%
����o��E���[���0�L�UD�	[`F�y��XM���NmZ5�?�3�'k�hs�h�f"�UQ��l�'��p�w�܀BT��OҀ_À���;��*@�J0Yp$��'!�Q���͢ܸ$��'@��'H8��Ǩ�%4�8V�ЩND�� k	�5��RF+>�O�Pî	c-�d�Fϐ�k�2���3O��qV�Ko���f�O(�c���ԟt	�	�U��ud�+��Z��W!YWb������𣀌k1`��cĉ��IX�  ^��|3`̊��D�*4�Z�O&8����?A��ƂkW�$Z7j�g�V��Y�<����6O[4���#�B@�U����'�R�0����'�/s�D͓xj:%Js	H�'ھD��O9 �B\a�I��lӮd�I:�?A���MX�;&�Z���<Y��#HHn����#%�ȩ���5O�8����oJ�<�U*��<s��~��&��A?�Їz>%i�k܉afTL�f!��
���7�Y�B4ּZbNՔ,��|���n�!q���f�J�2�L��y��W(�(��U-�~�K��|֧�tn�O����� ct\�2&?C�-A'�'8���ǀ!+���f��: N*E�� 9#��u�f�Eb�Fx�8Au��>ɑ�'v���;U�8�CI��\��9���<Z��b�� @B
���%a|R� mm���O@���O��e����v	A�|�d�;�4~W���O. ���.=��sm��(O�*��G�-��h�LI@���q�|�\=	��Y�&'l՘�G_�R�����[�y�$M�e���@�J4���)%��@��UZB�..T!��	��y���;_��1s�?0N��� ��y2	�u�� ���=	���������0w�"�N����?m�%�fiQ�6��dN�'��O�4I���r]��{۴f$y��-k�����;Y�AI�C�$�~����O��ʆK�t��v�F6�?���'x��Hc)J�-�he�ӈ��sn%��f?�5;�H�9��	�O 1�%��9�̰¢�X�y7�x�ӞxE���~� 瑶]ꈰ��e��t�F�A�A3|z�I���x��f(�T1��j��Fyb�O �΁��&�Uhz,i#-��_�Ҥ�([����ȯ`�$�� �I��I`��<SJ��BR�N𰸒��d��t	�w�(x�,L�G�Bc�(N�q�f�8ÓE!"=���g1��	0�ׁB����"O�
} �8S���oA~�ӣ��z�'�U��չ�l}	���>���[�4.��C*�j@��Њ�t
�-�'�*xB�OP)i��ye�����
�G$0�`����~bE�U�Qc�͏����!�ׂ���
3.��%�1M� ?}���ϊJV��bO=�əd������ �0#|�䥓).��H���o�
7Ο� ���dJӹ$)Q�� gC)J�z���HP0��3�l�+A�6��@�ן��@���?9��N��m��9�@�C��n�6�_�$��2Є��m�ń�	C�x�r����j�Ƌ�"h Q�u��"�~���p������pI�ӽf$,�j ��p
�T�ޠ � ��v�i<.�!���9E���R����M3��
":{ށbWlH<�A����-c�L����+����IdZ�Iڰ�Ƕp*��	,E�<�C����m��M����8kM�6�M�J3�H@���<�V����ɀ@□�3왗Z�K�Y٤,H�nh}���� �� #I.y|��K�ܐ\�T��'�=P��ǏL��J��@e���\�'�!-N	V�xI�Ԁ=�}@�'Q��e�~�,�3����#՟�%�ҟ�[&�ԡ)|d����4,����1k�X��y��_)�I��'�{��#���b0��6X������N�RjD��(�,Fm��"X9{��5(!Fu>�c6��&x�����F�RbT0�5 �s'd��0��;lw�xk��	�"�?�1�nn��+�'�Y����)RI�DGxO.�1��9i��X�(��pDd6���qc/Ԥqː�P���~x�]Hgb3��,;F
H�J6d��9&,��K�<c�$�ac���4i�<a�@	I�dҦ�d��c����C2)������V�A�\���M �d!�v���B�FL��%Eb�t�H_>�B�(a[x���סh
牮`t���'�l=�2��6�>���m<�T�SԦI�p�·hI&�1��џNZ����%G�;�]�l�8w���'u\�d��/����"��]-NX�fn  l��	uj�[�2��ꔅ.f*���MC�+T%�J��T=�R���9�p���/��}��82��e �ME{2m^�����c��q�D	(�~Z(�Q���En������V\�l�t7-�[��ũ�#-A.�:d����G���(,hL��Õ�|�8�8���~�6Y�ܴIRp����P��q����O:��'��ɣ����6t�ݧ���*��Q�6�r��g�Ӄj?�]hT�܎bz�k#-:�(�r˯~ҏ���:T�����m��U� V�K�n��	i��I��1!��D[r��J<���]\�BSC�'��H"�*���ȅt�d�?Q3(��2��.�0^�̩1���9\Kq�F���D�1ݸ�Ʌ�J�k�z�O�O+��A�P:G��)�����h��Kڐ	��LrD ��g~�:r�)#�"ex��:6b����&�*
��}��*í+�f�O�|��"Ӎ��4h��,N���~bq�½�N�W)�&���EJ�N��v�̉Tj:�#���71H(�	��y"�B:�L�	�7(��Ug�n�X��'����r�[%s7\�r��ƨup��y��̽l��T0s[?�Ey��R�^�P�
%�D�Hf��`�@�}��e����Z�~R�^Ϻ#B\�`�Y�M���a �.�h�����]����i'X�� �D\���d��	�N<I�C�B�,L��Əd՘� ��Գ�����<\YS���2t
�{"��.ڑ�t�r+j���Q�J9z��O�ܙ�M�Zh�p�c�\�0�\P�'��T�"��.b�μZ�k�*~	�Yشjפ�������~P�'��"~nڬ,���	�3Pe�E��Y.B�	���=q����>j�xt�=�Ұ�-՜���ԁ?���B��O{���'1�N��T�쓑�.�h˖�,Y�Q���pX���ۡ%��@���-'m����Nx���kZ=%cwĆ�v��Qc#$�3Z9��q�i@�~��i͵+d�Rs���UF����$a������ʨQ:r�{@AȊO#��j�nb��ɛ�j��b$����!��1���B塟�jAQoyʟ�D�#�,�ZZ��&A^�y"�<�Ҷ��A�oӴ�tE��\{T-{�]�$����E����^6T; �qă�PJ�|��+X
Z��	/��	�9t����C�'a�B
!Bv����)�d�i�O�h$���
�D�<�?�@��|r��${ȸp�PJh\�X���с`G97�.D�"�/48@��mt��^&5�ڀj"-E$O��AULKh��j&%�O�٢)ѿ7�Z�X�嘇 ���O0d�Z"=����;)�@��v�S/P�P��/ҟ��"6��!�_�n�8Q����qO��hR�݅�?�)�/I
7'�3U�r��	�:���_R���]����ҷ�rӔ!B�C�tb���zV\8`��>ȗ�z�pΫrO� pF�lY�1�'g�(�"'����dɆ%YSz����Q�0��("0�2���g��>4
W��MC3J6�	����Љy�S53��\P�A^�W1�u��!ʰF<T1��%����ɐ��3w�'�`�[M�.:=�4*���KWlr�Of���@{��?QkP�'����ȕ(��2Q>*\c�*v���A�T��yR�XC�U��b�����!�B������yq��rV�d_q����I�'��e�F�j���#�HzC��Ha�������/������l}BlL/�y�I�=�f�2�Ę"���?�	g�0h�%�?����I�2BX&d�����?�� Q��-!�mRi I�-�_�'Q�=�ҢQ-B���@_j�}�%ͣk���%̯<��%Nt�',ҁ�A�c�$Th��."�D���*8O�)3@Rex����w�rPXi�`d^,�R�B�)�%������Q�DٯdC�;��j؆p�r�+�gJ~$FG��`Ɖ�o7�ƺc��hS#`A�b<�1�Q�B/�џ���E��E���ÌV�J=dm��戋�~1Z����|O$4h��ՀHX}�'�L�y&�Qc?a�mד��'�Z��X��3�f����s���/�̼9�<�Ǎ8��0���'ṯ�u	U@�'-�p� ��0E��H@�W��D��4PN���
Fy,
�V�@�=�;d�x{�H��L�^4�ǋ$	��D.��w	���p�5<O��;m���NBG�����C�j�����Ξ�-�$�s�B̡x~>����j?q���
�� �2c�\�)�f.�$a0�ܸ�I�YC���$T���v�B�k�����+?�\:喆z�:y1�̲N������'�nh�C��7S>�-����p��Ga���
Q�H*��B�#B]��EPզ'�)�'G䐹��0Ve#��P;z8z�p�I��J�Oz�F��O� ���n\�-b�3����Je
�ᔒ>�c,Wa���՛
�T*�LO+�0��%��~��EՀrN���>}d�xWi����cJ7Q� �O�i�V�ƓL�X4�c�.2��
���=?�,F|���F�L��A��ŗ~�z�ɇ H��H0�p!����.U��c�-_m�����2yH��B5Y�f��Ѯ:��S<Q� 92�GV�n��t'�.�^B�/F��]i#��U�L؊����z<��$+Z���[9��<i��*���#��v��0bk�P���1cX� ~~!!���)_:ex��ûk.�y�3�rh<�A�J,B0�FщK��-�q!D�'�� 1G�U(f0�|�#s)II5��[�@��v9@ "O�(�$5
	*v�@mn�9z�?O�A�T���"g�O?1kBI ���W�'??�5jR1D�p�	�l�આ��V딼�B�0}ZO_`�X��'���9Mէo��0�T�[�X��`��'4����*f��gW�HjTc	�'��lu���(��NA�	�
�'����+
�q�xx�sfH��^�R	�'Hx��"������#�
uV���'4蠘7��(�"����$zgj���'>F!È�m@JY��K?&�4!j�'���j���87'Տa�J�#d�d�<�Q&,�U����8`-��/�[�<�eJ�1d�1��A;�V� ��V�<�
���S4���nO�<�Ŷ~�Qf#y�4A	W��M�<����'7�Y��kFf���P&*HI�<�$ _j@%�eS�c��T��z�<�^*� �a�?1��S�X�d��C䉪{�l�s[������V�,�C䉜@���U��~������*HrC�ɉ
�l����x~�!���h;�B�� �8EPS��kd�0��xU�B�p�*�a �7D�V�sÏ�cԨB䉯X�¥�a�6-� �cf#�֐B�!+ǘ��Sg	%� �QfB�I�Eb�\��H����c�lB�ɡ|nT�������9@(��l�B��	0	ƨ��K��K`��:f��M�*C䉰~�`�@�ٟ����R��%h�B�	�B�Y�5n*{��ŀQ����C�	 8��,	�D~���G/�`C�	U5��3wCձh��m*����8C�6o�8a��>����c�5SV^B��&Mf�q-�n���-_�g�BB�u���0��[3@[�1pW�@&=�B䉝X	��B c�c{rm�^�a@B䉺q�n0�*�3<�@�ْ-V)��C�IP��9ٷ�^�A?���͏}��C�ɏży[ǭN2��U;�Y�a�C�	s\�Y����-Q�v�0Q�,�DB��9'B�QX��]+7�L�(c�X�D�dC�	M��+� ��� ��-�BC�	.V��e�%
ѯIBPѤ�z��C�I�u�����˭�Йq�P$p��C�	�b��1y�U(l��MfHß$h�C�	�,���$KR�-�qY��7&9�B䉕��36&��	Ud��q�ڙP��B�I�=�u�L�)h\, �L+~-nB䉣F��9�����\��� �G�(B�	
RCj!Q¦X�\C,h#�+@/��C�I'uv8��hӘ5V� q�!� fG�B�	O(D�'Jڰ{*j���G��B�)� �!!�ϒN|"�`p���y���3&"O��� �
`X�C�jE[�h�+�"O�lqW�Q�j �-p��6�X)Zr"O�Q��9E�"}��Ҥ+���%"O�&��%�"�J���"���"O.��e�[�{*6m��;FVx��"O2t�����)ȧmF
"l��"O6LZC��N�:	��C�A���Q"O��;F!ۭ ���Ak�	+��"Onl0U�Ω7p"f)Oi8�j3"O�M�c��T���%�;~ �XX"O��A7�ūI�A��AC�@-@�"O��q�g�l�$1!@��&-�42C"O"h#�IC-��J�%�(\i`"O\��1og��T��#O�B�e�f"OT$�׊O�¤Q���F�\l2�"O�J�.�%l�x�1A�`S�� �"O.y�G �E��)�ݏ4K��"O���Ǥ1�����͘�<����"O&��Pǆ�b�f���%�U���bV"O��{����]�NYZ�#]�-fR���"Oڐ�%�+U46�ri�*+r�݂�"O��f���>� �SG-_f<(W"O��q@"�'v��	# 4.� �"O�0!e�=���� UL�1��3D�T�G��M�<�c �:2�јE�2��0|B����|sdAA�0$��d�	d�<w+\�t��!`eN)AS lx3�b�<aR��
Ma�Q!�:A�h�`�<�6�A)H�Kc�˴ ��6�F`�<�B�ձO�(9��e3/���r�iBZ�<Q��  ����$N�h�:!GAa�<��bJJ���a�D#�����ƓB؟��6�<��\T'��CO(w��\��	$����킴W�Ru�C��9�m��Vb��A�+Waȱ�2�
�y;��ȓ=i�L��呍 70L��.	��$��E{��4���A�i�# �K���;7-�y� *�@IbD�P�J��5a���y¯8Q��P��I������
��x�IT�t�pU8H˘.R�1���ݎS�C�ɰZt� ��&�O:���l�S0.C�Ɇ.Xe�����`�)��0
,<C��6#�h�A�8I�� 0㕓S��C�I#(���9�,�U(�੗A���C�	,Tq6�
ß�P^��� �;��B䉦w�A����s �Å�F>VPC�	4oEr`��ぉ.���C��*C�ɨ���`��ր[#4��aW$4�C�	1fl|T(/�*��1�  �C�ɞ#����RK�>:��1��^A�PB�(��9�#�.b�h�&ǁ;"�0B�	�z�t�xgE�?��H�d�Lw�C�9n^�Z��,���@�^��B䉥����2E� ��i)����BB��4���3 ��'4Р	+���&THB�I-7�n9��O^�rl���j�.B�It =&�V��� �!-��B�Vk~�2�@۸0�fD�D�̘q��C�I��<a�#O��"磉\���'_a}�㍂	Ep�a��P5| Ir���(O4�=�Or��� ��an���U�l��	�'pI��ʸyN.��� 7r�X�'����$�+Ȧ�*%O�{�
� ��� l@
�.����
Ǩ�� �>1j$��(��ɹblQ��J$�c`�l�`C䉯�y�p��#5���D�2�hB�7�H]��S�IQ�ɪ��ЙJ!!�����ibK�=,���SWh~!��.b���c	U?a��dR6�ĺaY!�r������2��kG��I��1��7U>dKK^&(�*�S0��GN�l��.��Z��'�h3�ֻBx�U�� ��� 㜊.�����lڠ50 F{�O������9�����M�,o+����'�ҽAR%ҹp2NP)�)܉e�`1"��Dx�$��$��f��BnL�>hJ�Ђ��*z�!�$J�f�%z� "Y��*�ba!���,8�B��կ<�ҁ�0ᚣ\O!�$�9h!X��V��YSō�o=!�H5�b��,9D���K�䗱(G�̰>aT��6�� ��k�*[����N�<a%F�}�&�Rg�2H輌@w��G�<���Z������`�v9 ��E�<�k5	��;�T� @����f�<�0C�{��)KA'���5�Cm�c�<!GO��+P���.�DF������C�<�ƍ�?����,�[
����FJ�<�"�+䙡4/�u�&����F�<ɵ�Y~�A��`�7-)
�I���B�<�w��K����Ͷb��ء@�HG�<�#�փ8��t�]Lz%��F�m�<�� ��(��P
��b��Br��i�<9#M�tRn��Aʍ<h�B�v��p�'f�?��D@�GLqxB \L��@���#D����ޣ!�4R����LUPd�T�=D��i J@�j���	��� Y`sl;D��	����G{���6Ń#
�*(��j8D�Ps�?E��D3!�Ad�@H$�W�<�*N �|�Bǉ�$S��RBO�R�<�C[�=�(�ڢ�ԡ}����PP�<���T���)�6��Q��	rC�g�<Y'oċ}��86�M�"<��1�[g�<1pi�5_��@Hb�ՙ8ʡH�*\�<A"�U<Rέ0�ܗ/�� ��U�<QU�DM7tݫU�OV�� ��M�<�5�D�!E\Xj���?f�qȀ�F�<y�Ii>ơ�5M	61B\(�N\�<��K��@t���Z3�rg��T�<"�U�i[�m�Mټ��5!�O�< Kf T�� ��6<��:��JM�<A�G9�ơ���	��2��T(<a޴ (�Ҵ$�uPZ1��ؖB,���ȓ#�XT`��ˍ}���[�*̒_W�����Ԙ#FTcP ���ǅR�$�������F��PQ�5�R>9?��=ۓ1F����O7lX���ö{�(�ȓ���h�aB�wN�q�wn�6g*|���3����$B���D�p�B5��}��$��r�Y�m�x�Y��ʊ3��9��G�t��6��V��Y��u�N1��L�l�r��ْ-,�E)�G<;SɆ�o��#ņ$fp��ä[�� ��'���	F�Y�1�.L�#%�^P<�2ӓ��'�x�;e�hg�E�S�G�@���	�'/�AS�([�R �t�>o&�0	�'n�U��� s.�QDJ�~�.Mc�'�	�ΗO�p���P�}�EK
��� 乚��W!j��h��oV93F��s"O2(����P��,ج�r%��"O\iZV���<����eݘ��"O��y���6 <�R̋�����"Oh9Ia	�Z�L�Ytĝ6P$���"O*,��ڴt�N��t�(gHZ$��"O�H�d^�I���2B�DB"O�Ihu @�p�
�j�8R+de��"O�㍮k��ˇ�V������"OJt���)8�
x�-M���y�"OAB#��2&�Q�䪓fe�A�"O����Y�pf@l�P*�5pd]�`"O��s��;D�H�F�Y�K�̘�#"O�5�uN��%+2b="���"O�5��E�?#��P���"r�:�"O	zpG�8�L*�\�TMҧ"Od1w��W�e@D�@�[�n=; "O �c"+��@�ljԍ�)'*|i�"OХ�&_ܰ!��k�#@�*`"O��׊�(PL�M�I\�����"O��*5 �0-d����A�4b� T��"O� �u��%��xa5F��X��"O�@�᐀=X�H����	���"OfA2��޸,� @��oU�i]�X�E"Ov�ؗ�V�=�P���V+�}H*8�ȓ|�t�����8AB<���N]�L�ȓw��Лm�?5�H�8�.�Bp��;H	ѥ�E�{��M���m~`A�ȓ@_.�AC�A�;���%kQ�g�T�ȓ&��H� V�ͤ)��G���FTr}����m�ѩ�D�	k��L��7�P[���0���۫AP8���t�`7�8������ApR�ȓ�� y����2@b8G�G�1�u��)�\�p��?=��'.@�x袝�ȓh�5�2 o��AS���	�����F�2�x"BU*�z��p�A��y��Z9���"�N$$|��0��QJ�2t��{�г�n��
*�i!��ߏd�`��ȓ��4��㎞�v����.�ڔ�ȓI(�a`�؉(�L����Ƅi�Pe��C�����D;GKD�X��_ ����ȓq�j�8��,{	v�i� �=Y�v-��y�u�����Z|9���o�Ѕȓ1�(�A$�2*X��@ьcR�e��r��²"�5:�����r7`���yiV�Z;��A�M�m�؝�ȓ{�,qPɏ+w�{�G��~v4B剀-,�1��2qp`U�5o�c��B䉃無��8v��hc��}=�B�I�F��� *���8Q���/ʖB�	7��x����~��qS#,Y*
RB�I�tn����Z/*S�q���p�zC� ��Г��M�y�mb#`A�@xC�1+�X���ōH��\3dHC�	�D=�$H��@b�}b��Z9e��B��'�l�"�M������3!FB�ɣi�~���)|dI*Q�X�"�B�I�+��y�G�W�v� D)>�C䉏g.����N�7h@�`�@A�C�	z�8�S�L�y0�ٯa�$B��:�����$L�
�跌�"s��C�	8\����5�],Ji63C�T��C��{Ƒ	���e8�jp(ؐ{(�C�)� �ٹ�K�/T(��Z�韖t�diX@"O�k1��-x}BM{$>�X ��"OX���	�z��}���L6U���"O.tCaK�0 ���ḝ"O�d[�m�)%���"ʩsz�#�"O|q����)���Ú���"O4�`FO�������F4H��&"O�u2��3-� 	�%��$�4�sW"O�	�[�^:�9R�HH�ʍ�W"OV���E�𘙡�D�m�4=!�"O�� ʟ_�D�Bk�:P�L��"O��Z/e7X�RQ��!�\���"OĸC�-U�Q����蔋r�4�d"O�ͻgކ[�iC��G��T-S�"OLAR� N�z��	.g0�D�a"O`a2R퐠}d����/hN�0g"O> ���00�X�s��.p�pb�"OĝpF��S�b|[b��,U���W"O^	��㒑�\@���4v|��9�"O p���;M��xWGܾ\_�<Kc"O*mӁ�X#Q>�� �` �;;Q�4"Obt����S"��Iƅ7�h ��"OX��<K=�h��IE(^�D�`"O�U�E��;<��y��S%l��7"O�� �ƞ,J
�-��� �Aΰ#�"O��3���a�đg�\'E�Z<��"O���&�"��}�TG�n�H4xW"O�����Ґ!>V�j��*z꙳V"O�D��ȵ�v���ӫ,c���"O�-��畦� ��V�ղ� M*G"O��;%K�0s�� ;�9���A�"O,�p�+8����gW1iy^%�4"O���4O����E@�V��Ks"O \�%�2%�E�w�5aW�ؖ"OH��0�"o��%Y�h�4.%�i�t"OP�Ʊ�*�XW	%v��ɦ"O� e�F+U��Y Xe���b
`�<iDC�h�����J�j��Y�N�X�<�1EP,OX��H�J�<����m�<aBmT�F0�u�V
M�[��Q&�R�<	2�I@d�4���%+' L"E)�z�<���њy��y�q��6��}hD�Nq�<YUŀL���Q@�*�\�"�f�s�<���@,6���'� @���B�Xm�<!Ǘ�48B�Z�
PR�L)G��j�<m�M��������}�E�@g�<q�)[?1����4`�~��'/^�<94IG�\��!dǞT�37)c�<�V�NnH
��Z�\��T�<1҃��3���p5Ҿ7�:�#���J�<!��<�p���ȏsXh$�F�<Q�5�����M�~�Ji��A�<I1�ýY3j	�f
��H|��G{�<Q�J�Q��Y�.1V�\����s�<���^�q�M��K�Wq�i��V�< ��8%�ҭs�dI>!cN)��AE{�<!�N�GYh�#��D=���9�)�^�<9��Y'q]r@������͓`�<��LB�NmZ����17K�e�<i%	#_�4��#�	w���Blc�<AC�ӱڜ����ïv,�E�s�<�(£4ǜ���
&���ځ�Uh�<�b�́4��Q����Ĳ��b�<i���M^H	CFÃ[ٴuRF'[�<� �E�� � Ϩ�� ����R"O�Z��ڂꚵ"�L��b|˲"O0��bLD=���y�g�`�Ȉ��"O�"ԩP����!���Y���"O��;3n[
i��ek�f�cY��	6"O ����S�8��H����`SN�{�"O|�b�*��ub�mQ&6J��Q�"O�}�&�٭�hT�DKRD���R"O�ѷD�f�P�xs��53,P��"O����n�A7�ij` \�C%�]xp"O���`�Ӳp�pe�n\-!�0d"O�x��ݧ*�<,dm��`t"O��BGm�8']�}�eB�sh���"O���sb����P!a˗ �rtK�"O�eS�C;:h��/B�W���5"O�-�/_)a�ԐH���~�\�i2"OJݛ(��.�����#P��e��"Or�:g�S�#4>�8�M؈SH|e)�"Ob�#l%1x4�X�+�#3��X�"O��Z�B�,N�a��P�hC
�b@"Oة�E��t�J=��A�EQr%"OI��(��V#N9/IPŹ$"O&`� I8l,����eZ8E��"O� ��B&FB�b�%\uFa�'"O����v�b��Dd�WyR�k4"O@�aD#w'��#��	��0��"O��-5��q�%��	-��ĉ���y��X�m^9��H) 3.`1��R��y��r�� �4Ǌ�zB8
4�¼�ybǂ ]�&q �ϱmbֽs����yr䃻(C*=	6���/�pY�r�֠�yR��b�@�#�̎�<��a+&�y��;���䀄�X� d��#�y�-5	�L�5!'z��� _=�y���b(�H��a��o\�	#f�*�y��1��<#+��f����J��y��±"z<��B�q,����@�yk̫� �yD�.6���\�y2煦l��d��,Y1M`�=a��P��yr��&�.8�
p�B�hl��yRO�s�r峖�I�W��Dz`c���y��,J��1�+KJ���bL�y�M�-�������u��Ph'Bс�y��;\����eNָi�0<�w'ʚ�y�ͅ�hX]��IN�g��T�ƬB�y"�=(��ǧI"ZM~4�BB��y�`)���թĳ Bp��KE�y��ҿ,�A�7-
eD�����yN�oM4�Y�$�j�̄@0 �&�y"�/
�́4	�<i&��;��̅�y�AR�'�����T7�� `׃�ybaH>���o�6S��1�l\�y"����x��Qkp�whα�yrBA��ɒЧ_t�d��hC(�y�hO�(et�'h����G�ŵ�yb���n -�Ui-dm`cW,C.�y�μuJH��^�J�0W��#�yR$��|�|�Æ WQ��jGA���y�aK��T@fEߣQ ��j��L��yb�D<(�0�I�mާ1��c'���y��F�zy��#�M��
��y2k�{�X�x��-G��(�a���y���=٘ؐd&E��Y ���y҆�#;RЄ�Q�u�c���y
� ����A%t�(3�l f�J0 �"OH�s�DĂc;`�C K]P7�0I�"Ob\�q�� *D"Ѩ�Bv��"O��Z�O�/�v�Y0��;r"��"Ox<AL�i�T���&^�{�q�"O�5�J�+6���׊�;ks��8�"OZA��� �y<���t�Q,Dvt"O��@Bزy�Y���ōG�z\K�"OD��ϗu<x�6�ѵ[��E��"O�\cI��8ru�!z�xHR�"OX4�P6J�����,�
S�Pò"O^� "(���|(�+�^ў$��"O������[�
0�Fh�X�N!�3"O\IG��{(�t #�IA�d��"O\\���	�+�(���f́Cƾ�'"O�\���N�z)�dU)	�b�"O��3ŀ �^,�X�96���e"O�AH�^�U�@��#��H\�i`"O��˂ugȍ�2c6I8�d=��CMұ�fP�9
F٣�O
f�ń�3��+c��g٤�c��@�R٘��ȓ@G����']!�p�! ��V]&��ȓi�(�@�
�R-xF�F*F�^���*W�`��A��4�J��bJ�B�0�ȓY��ħ@"S�D�G�f0�I�ȓ:�@�!�D�Y��R�"�b�4��7�p9j�/Y46�6H�j�j,�x��=�N"%�L�������y\���ȓ4�,���F	�T����$�F8�ȓy7�Py�jA�*���Z׆!����lg�8H�EM$@G�A26�H�6�$��ȓ`$�<����0���GNݬJ0����
�r� ǇQ�DQTX $C�'.6�ȓ��=��PKi���S�gP�ȓ\!��B2(�"
V���-U�~��c���ˋ�,��]����0iQ���)�n�y�]�0�t0�wʎ�ą�q�������;��2�X(n�Ԅȓ�*�J0�
--�Fa�s�ޗtb�܅���E��<3{�-[�5uK���'k֌�3kQ�k2h�G�f�F��'j<�wI5"� ��	Υ	G:���'V�|���|%��sю�8{����'���E�3��!�pH��x��k�'�^m"��)"2��i��} x��
�'��%Ѡ/	����a�s�d�b�'*Ha{#I�-J�h�6L i ���'$�U,l��2»*����̍��yR�G�_OP%�"��"')��3��_��yrm��<1�]�Nne�\q�e�7�yBj�e�
1{%���`�Gϐ�y�b�0,�H����ӾY	�)ח�y�ꝭ[X29�cc�g����`Y8�yϔ�?�u��Ě�_wZx�BK��y"����q0�	�P@|�g-؈�yR�ٰ.�x��I�r�Vi�d��y��n��ju�34�!1�� �y�B�a	���.�.%� �w	���y�Å:,�%�ǠI�$����lÁ�yb�� Ǣ��/�

m˖-Ȫ�y��29�V\���v%���g�>�y�e�g6��U��o�,U�����y���='G�]���\��$q���y���<RӇ]&<�X���y
� :��%D|�:���J ?�����"O~k@A�"��(�a��k��02"O@�@��5=�A��[7"p;&"O�E�dݑv���H��ֱW>���"O��-Y �l�c�	yP�1�"O@���BŒI���"KX�K瘵��"O&좕MY�F5�#/'tt Ǌ=D�t����sl��Ps"��>^Ttb�=D�LKe���)�� �w/�>{?00�U�>D� :���b]���G<xf�1�<D� �D\'C:���d��]��Ѷ�:D��4nݨ+�L�W���!˾	`��"D� �%��E�4ljqd� B���o D�L��,^S�6�����7�p��?D��i�j�t�	s�^,<�Ђ�<D��(��5f���!�[������%D��"�N�/g��y�LX|zA �o>D��3gR������"��a��=D��)Hi[5�$�_KV�)�:D����~6��3��]^B-��l8D��0c��	V�	�Ro�s��eA�@*D�lHd���-{4�{��^�k��h�D5D���A ��4��@�ݖ<��c�>D�H�E�	3� ����?�|!;c�=D�p)u��-ι���؝^����+;D��H���A�x�X#䖄3r@ � 	,D���b+�$B�6Ȉ_�-z��(� C䉝g[��Q�J�S���9G  T�:C�I�/[��8� ��wx��6�]��:C�����A�As�YS�ښX�(C䉶,l���@ 8Y���s2KU�49C䉶_�e�,� {zI��ݮ�B��
N3�1TD|�F��!c��B�	��>�c��`"� Ε9oɮB�z�rm�g�&sU i�LU�$1XC�I�t@5j %.�8�&U�U*�B��.Yx-���2]�dl���*N�*B��>k����rg�pD�i6Qn�B䉷B� �M�H�R9{� �(�C��,*�``�QN��tU��f�
C�	�{m2qA���v(P��ۙ�C�I�s�����>,�(�RM��B�I�A�����D�V�,A�.:S�C�	N(�|��W?e���i�+y8C�Ɂܟ٠F�ʵg���1'*�a�<��A�e�3Esf9+0'U\�<���	U R����&W~���PW�<!�nW2��x�5l�"z��X�P�<�1�ź�`�0G���%�@B�*�I�<i��\��
0`0�Θ���kI{�<y���� y*�j��KGbE���R�<Q6#��_<"��q�ST(2��w��P�<��JY.p3CZ d��A�<��`�#/�&���6w��L{�u�<)sI��HY�Q����|�.����j�<��FB�X ����E�@yC�A_�<	eKE�$.��r��H�n�(�NPY�<遅��8�Ո�!�71��=�⯝X�<	�B^ROz�F���v,�0�l�<��	@2ޖ(P�ˇK��!A�nKN�<�C�&1Դ� ���/报�1�K�<2@��e)�
�eب�2+�`�<)�Z���qi"⃂��)�V�b�<�vK·Rꞕ�"l*E!h��(�_�<� l	`�e>W��9K#pBR�"ON�3�\�$�bd�G�/|ֱ�"O$-:P����UI���tg(�;2"O&틵)�	R7�ɘ���I&�B"O��c*�fל���#J��
�'��6�&޺9�M�;k
��'��P�S��8PN�q�i��je��{�'L4�҇
p)@K�R���'r��$��G��:D��Q�X�)	�'*���7b��Q,,�����N��I:�'��8��ڒ:zr�j�=u�h�'b,�
�I�z舔����=�j�y	�'i��Aڲ����J95�Z�'ޜ%hT�Т,��L�"�1���0�'v�� f)���;�8��'�}t�80 Р�(Q���
�'��p�ƎR�Z��&-]1{��i8
�'�58')[�p��
��vlJ�`�'N��q.C%+��Q0�W -ި��'�����)3E8E �n��j�����'+�$ ���@q��0�6�P��y�
�J�J���ƚ<�|z����y�oV?6�Xջ�j�&p��OO��yRb_&`4H�k��8F�H�����yb��<|d
�a��� [> نM^�yB���h���s䋬<X�����&�y�M(Zt��`��b�&4��'�y�O�9J��ض��`�bm�oԨ�y�J��D�|B�D̜k��{B܌�y���}���C&�[*[D�1($H��y"G6�j�r��)˘8��	���y�$��v!f0�Oλ����W�ybʙ!nҜY�N��=������y⎘rHژ4�L���b���)�yrfF�T�Ѡ3Δ.H�J�) ���yB�Z(	#�}�7��B,�d
���yB�N'�7�Ԅ5�z����
��y�d�~�QFߠ97��������ybli��a�Ռ5�Ti	#����y2��9^�ՠ�Æ(��1r�]�y�f��V����Ǒ�W��i�D��y����8���K�U�^E�P���y�$C)~;�F59Ml�畩�y2$H�b���	uj�7���2C;�y¡�[���1��<&�l0 ��B�y򊉫7$��&�
(vib��&�yr烄g���òi�D��@�"S,�y����~��Dk�z�x��d�!�yR���|��$92��} �&�y���fR��g���˸�1�����y�Y,XY<�h��I�{ю�p&���y2��'y0�e�vCH)J�G��y��éU��*��>�l���+�y��]2\�*�K0 T8�lBVˇ��y�.�j��슁3K8�h5J\��y���'�|��g�_V���dfO��y�\,tr朡��^I`�i�cǥ�y'Y0oeɳ��4A�Hh��7�y�J?q�B����̩=���Q@ȓ5�y�B&��iQF�ƴ+i�8+p�E��y��ĪP�$�(N��~�Cg�.�y�C��9���b�jֽ Rl1��A�9�yRaD�K��d�t`H�cI(�N�=�y�V�W���`�K8U?�v����y
� �͡eO�$A��d8RJ�7z��F"O�9 �'�y�|J4鉩�r�˴"O�l����P�0����+c�� �R"O,��caR��PŨ!hF�puhL�'"O \ P���l������V�Y����"O��;��L�W�P8�Ff�6Ep ""O��PQ�ǿPuh5���L.&�J�"OjU�UG ��rS1t+H��1"OF �G�!7K��6�s�����y�m��ڑ����y��䩔h 8�yrJ0��� ǧC0�\��p�'oY�n��cW���W?McB���'7��@ŝZ�ZY�#�Ä78���'QDU� i�5Ql �Vd��/�:��'�z��X�V`½{��#�ub
�'�b)�ǣW����l_iӢ��
�'Aj�тC�Uޭ�"L
�*��T��'c�p�E΍;I7�� �H�#�V��	�'IX�́'��4)ֲ"��=��'�L�ӡ�6�^\"�c�j�:l��'|�Xxl�7'R��)�>[�D���'�02+^+8���)�.�U���'�R=�`�	��·'�X
�ȣ�'�^mb�����RP
�!W

�'�>I
���w%"���ᛸe �B�'���P �ہW�2	�m�2�"��'Szd1TdL�R60�t��t�ju��'��j��ϟi�3�k��i����'���qsN�cú�bCDZ]�v�@�'e6�CŢ&����bV7c����'E,5� �H9]f�|��U�ao ���'� Г��EcDD�����N�ޜP�'��4s���7ذ���PMgb�'��)��W�X
��r�A�x�(�'(Ȥ�b�J�t�J�x0�J&i20��	�'���P���2o� +� Y���	�'���C�/y�:���F�V�ds	�'�pD���m����%iT�Q����'���0ݱu�� �p���R]"���'�Q��0���kW�NW�I@�'������nŢ��aO\�I��3�'
��:�f��;���1ጥ,yP��	�'�x��dY�$2�tP��-B��'�����K]?O�Rٛ��,J���'��B�/^���A ׏9@hR	�'��x 0%ޞM@���w��.7��)�'x:��-�/��H#4�T�Fu�)r�'l��
��D�@n4�㉉�t���'�b���)9zD���k���'m^�;��:0^|��>cd>|0�'��e�b��H��-`�&�ZW��#��U��κkH5
5���tA�BI'D�d	�M�4\6$�!�:_%H=��J&D��ǝ��Ldҧ U�C��3�i>D�D�A`.~Gt�����
�pD�@$:D��Q�C������%�Z
p{bD�w�6D�ze���� 3�X�.�(����'D�hZe�2"�Fȃ��4t�qp�%D���"Ŵg�ac Q�/�ʑQ�#D�H�1-�P������`�p#D���� 4n�y������.D��z5��h���p4��f*�'�+D���"_7X_>(36�ӣ���Ӗ�<D��a��-Z^�Lj���'d��]zv+:D�� E����&al�5B(�Z��Y�"OUHcoC������e�3�Hш*Ot�+5,N�h�]R�aD"j�� b�'7��Ɂ闖0� �3�	d�̲�'y��M*z�.5"��P:hjX]`�'�q06��:OT09�V�h��t��'��y�`��x�0(pd��g�Ī�'�v�K.@�')��V%��q���j�'6 pXъ�:�ԭ	��Gg�@���'�Z���Ǉ�Y+�\����m�<,:�'��A N�uG(��'疭t��R�'W�)��g��{���r�σ5�t��
�'��us�ʘ�V�
c��52f�h	�'@hR���-Ip��b�ӳ9��x#�'%�11`@�T,�p�I٬7.JI�'S)"d�R��@iې j���'I�����A>2��0��ȅ$�m�
�'q&��M��ʴ4p��<T���@
�'�8���X*X]H��v���D� ��	�')~|�Ɯl��S��� -ڝc	�'t�2��Jk���`����c�X��'�ꍩ���C���8%�R�� ���'B���+, �8 ��ɶ+��'ټ��Q�P�'��EBT�Ûuc�}�'l��d-����۞$^��|��'�Vh�K�*t��H8�!9P����'w����A�i�J�է�KĠIX
�'wdْ��ےd0>����̔;Sxu�'Zj�r� �{bx�e��0�����'��a0�h��5	�嘧11���'r�����W�E*�e�z����'M>�q6-�?0޸�a��#=D ���'�f�S�&��<qI!JC�8�8s�'�Y�ƌ7٢�c� Ȭ,�vu��'�H�
B����Jt���Q,$��]s�'�� ��ǻHjRI�X���0p���{���/�H!z������V:�ه��D|"�.R�=7�pa	�E�����`�$��'�M���c� V�"�b͆�!�4�*y(J {S͒D���.���㇅�"���3���<	��v�������5�0,����1i� �ȓp>,"7�׆	�F�A��W�1�h�ȓm�뱍�,b���bi�)����-1b�$�]󐈩�ǋ9��ȓu_�񉡤Y�*���ɞ�U���ȓN�����i�'V��QcFܪ
/lH�ȓ]d��k���0iI�8��`ZD�$�ȓs@��坷yl��c0&��}u>ń�IY�eyÃ�{hr�� BF`/���f~����Eр|�8|���K;<WX���W�rEѣ�G6+˜���m�<A�����Og��ea_�e��\���:`Lⴆ�]Ht�AB*Vs��P0$�ȓc��@Q��˲��c5�֖:h ��f��ē g�",=����� >bq�ȓ@�~+'KS�W�aC:'��ȅ�^�t�bB�(�Τ(�!�7C��ȓ%�Hu�4�N�00 0�@��4���2�_7$�{�
/i�H݇ȓ-�*�s�G�b!�%䊧^����ȓp�`d��H�;?�p4k!�^̈́�h�r���ߟ<�l�˰�ّb�"=�ȓ[)������EV��m�����S�?  �����'W�����`�GI�d��"O`!����m:��s X�->��r"O��#E,/7~x<��oI�7-rX�"O)�/xur/\�k3>Z�"O��c��z0���ƌK,��f"O,D��_�|H����1 �P囗"O�C%�[kJ6i��ڒ|�\"O�hz`�Ĺ���ʁ��"ڠ�K"O����H]�01:��C:J�
�۔"O6��W͍Ҽ�: n��MZ�@w"O�49���Adu����?��i� "O.e#�K�p�4I!�l@:o�
81�"Oj�����<R.F�kw�\&t���D"O:Cg�PBs��׺�*� �"O6\�f��,~�b@!��rp��3�"O8����8:�mj
�mYt�1"O����)ܞ��Ph�n��桀d"Or�H��[�Τ[�F�S���y�"O�u�*ڽy/�P��:C��"O���nD�$����� q1�;�"O0�sPiʼb��U!g�Fd|3"O�mxa ��O�`��%@(L�q�"O�qZ���5��mj���, ��� G"O�@	 oآ���M�="C��k�"O�=���!Kc���b8<�"O��@wm���^�[�k�+WW�m��"ON��e�D<F%�Bʛ04&4j"OF��q爫y�j�X�H�~��*`"O���g���*� U�cb��,�̰�f"OҐR!U>%f�G6 ��Ic�"O<1�T�Ο~�H�صFݕ�NL��"O�������Y�7�D�["�ف�"O>�`�N��I�p�>��K�"O 	�V���d8�C6���mJdJ�"O~�3��HG�:S����4 �"O��ǅ{f
V�D��C���y�%��phֹ:!M�}Q�!#���yr��H���2�̼mL걡�c�1�y�m
^���T ��k��Ism�5�y2�Z�J��֡�l͜��w �;�y��.�^���� i�������y�'��`A���1S ��&OG=�y�Ċu���e�Jɉ%eԡ�yҮ��!�0�Ba��6��{u�7�y�&>M��Q�o\>"� hB��.�y¡�r�~L��k�?o���!�P��y�E߇9��0e�ղl��d��I���y��U�D�
!�_���4�!�y���4}mШ+�nZb
�dg��yl#7�@�傴@X��!�mė�yE��N����؍�M���(j!�dU����ACH�0{R�]��'R�K!�DS�yxʴ ��ID��拪k!�䂵L�8XK�'Z�@�VŻ��	O!�dڑr�\0q�G�e�!,��/�!�DQ���<��R9������Q'�!�]�����;A$�Y�� #�!�d@Z��x���.�	��Y.�!�7h_Xu�%kW<"�a��T�T�!�dK��$<p��R�mx��`Y�P�!�D��^sj0���ʯU`�t��*WN!��'�t�)��#Sƀ�����2!��^�cn6�%�F�N����8Z�!�ć	0�ND�&	���-��*��K�!�� D)��(ظa]
�K��)z��8�"O�qA�h�:?��Љ��D/_����a"OJ)r"GR� ���{�j\�C���Y�"O���v,W�:Ͷ%ɥ�D�K��m	�"OF�[FN��"��ő�뀰-�����"O��pϕ�|��
�Û�� �"O81�Ɔ�C�-�Ӣ�6kk���"O��炆���}��a��?����"O4���.чr�4}B��َ)�<`"O���$��Vd��Eɾ<aq�"Oh��e��}Q�����>=��%�C"Ov�zr��+GĭÖ���c�$��"O~��w�n�s�`>X7\!��"O��_i��	w��2"O쑪�Mt՜cm�,%28"O�V��n�x@��b��J���Qj�O�<I�.۱,���
�b�;� �� �N�<1P*�>���q�Tb�P�U�<ɒƃ2JSF�˓�Ԕ(��2s��T�<�㮚�T:�`�%�H�5\�A9f�E�<i F�!�� ���G��<����[�<!�`W��~}�U]�vA��D^�<���=zE��
u
U�cD�@�<��*a�h��
2�Vi�d-��<�S'ͅ:F����@_�@�(�w-�F�<q K�^񡣦�0|"�8Po |�<i�ګe#�����*3$r�H1�u�<��7SCn��6�̫u{@�0���n�<���!^�*i2��qn�d��c�<�W�	5Y���c��{�"d(Sb�\�<��ʃ�h� AU��>�&x�S�a�<9�I�q����"'�>:��ۅ�\�<)e	B%d�E�T	A�. \U�ea�L�<���CH�$�xDI-|��qcI�~�<)��Ǐ
S� vM ��<�y��f�<9�űl.��{�Hڋj=����z�<�tm�?sR��3%�YڐaC�MQ�<�Ԃ߇H�:,ۂ@U�KF�=���GK�<��HK���˜�D'Lňԏ�n�<ٶ�ŀn�rHIC��C��6J�g�<Ѣ曇(��V)K�fol���w�<��(�Eu<����@�'Kv�Q��Jr�<YAF�[��r���<V�F��[u�<Y�Dֺd9:(K�� m��A���r�<9��F4k"tI��(��;N0�s��Y�<b�*����,�)]�I��S�<��A�@�����ˋ1C���BC�O�<�''�?% dX�"&'��l�b�a�<��#*L$��(���m��S ^�<�r/�[��e�#���j���Z�<�Ņ�=�
E�U_�N���
�Y�<�W��(���G؂q)��RƑ[�<���	>E�=��@<@�&;��X�<�懒��ȼk�c��@�J [��T�<QP.� t�^�5�h5�b�S�<a7�рV7�Z`[�"�y4�U�<1��,�=p�͗
%��Y$L[Z�<�[�>vvp �N�"%@�Z�
�m�<I�C��քC�i���M0��B�<1҈���@�Y ��"�A�<��Z_������-s�0S7��}�<�+�'6	�!_�T`z�ڑ"O�$�ԋ:�V	y`uS@Ы�"O��:�+[�Wc<���U���ۆ"O� ^8��n�e�<1�](r
X�r�"O��qF�y2�)��k�){���z�"O΍;s�K�\��Ĕ�6�	hG"O� `����GT ��m�4 K"O�t��u������A��p"O�A"�[&:7ZM�f�30$��*Of�����x���3�S�����'��l@�	C�d|3��jD�e��'M*92��**��SQ����'	XH��!9}�h�Ñ�I�wA����'w̝�p��{�ɳ�G�i��[
�'v M�Y0;
|a�/��]��X@�'�\[@�U�qԬ�+4�C�W�&�
�'��T��k�lF�J��]+�h	�'�V�9S,X�4�yxS.�$Y�걣�'���7 ���0�ҨJ6\{�'��-�̬�Θ�C��G~f�x�'�1ۄ�@ ��PSK�F�h(��'��h�E�8T�$����>��t��'��-�S��<ײ؂���8Ȣ�Z�'#z�Ѯ��|XY5��3�ح��'����d���W�`�e	6 �@���'�Z��Q�]0�M�C� '�Dib�'Xd���/B��r3l���Ts�'θ���Ȭ,���"�bK!�*�'�@��@�%v�8Q��ъX7����'ؼ�!B�ޑ�F�A��@9K� ���'u�Äa�n��}��+ʹC���'ir�Q5���V���0&v�Px��6D�P"�����eٱAJ�H���5D�t(+1����K�'���S�4D��0�FG6�� !F��:��CŎ1D�|���Ø>�>ͻfI���pr��#D�p@CH�Y�4��bȦFKz|sp�4D�ӗ&TW*a8V�H"ɊtpG*1D���ǉ����is�E�+K`�Q�J*D��R�
?R,�h	�IW�6�"�fB&D�P�q�N+f;j��3
J�Y���`%D�8Q���65�(sw��6iİ�jf�0D�$��G�)�������8i��!��.D��1Ci���L��n9����
:�B��3�X*FO�,� x�$ddbB�,a�x���8W�Ι�Go�: C�.,�Щ
�薬OM��{��@�>��B�I�r⽊G�,{���{���*7U!���A�4�b�$>�2�1N�
m�!�d��T��a3�
K���D��O�!򄝙8��d!��,e)�̱�AɲR�!�dF9J۶oX	$m�enA��!�d�(yG����A����Do�E�!�$�2U�DJ�KX�4�FU)@Ř<!�dS5r=X�@1�?648)JfC��%!򤝑,
�;R��)9Vh� ��*!�$�h���1�$��y4�$0�"!�$E�a~���i����0k��x�!�$�?S�hQ�6,��DD{�G�Jg!�
%Y���rb�h~�]���DU!��M|�K��^o�����\�Us!�͍~�D�d>U�hh�k��4�!��(s��`�GV�D�=`�%�#t�!���fxt��.�&5�����$d!���9/��S�h��M9�ه��!���P8Z(�剄3*1�5f4t!�DJ�K��0ׂ�C�NM���l�!�� �=���yJ: �w��SF1v"O�P U��
X=��+��"SiF���"Ot��]о���^5=�J!Bs"Od�p��U�x<��]P��$υe�<Q�	��`���8ńJ�A��r&��H�<��`�*\E��eך\l�	�dR_�<��J���m�}�!�h�Y�<��nY�q�F�`�=ch����M�<)��\N`&�� ,�;�8H��/�I�<1�e�./������^?Hbm��$k�<�"-Oè�s�¼5��E��i�<Qq�t��%� �^|��2M^�,�!�
5,΂�p�c�sn��ެ�!�D��t��%�gA�kD5t���4!򄘦b�P���=�JMxa� E%!���_��FΚ,�dd�C ^�{!�$�Pɬ� �E�!��1B2Ϙ�B!�˺�8uY��[�H�n	=I�!�d� sX$�P�*�?���6���t'!��ԛl̠�i�k֌W_����F$!�#Q��+�)ǩw��@�D��!�E�)-@P�!|XlQ�@:�!��M+D���D�tx*uZ��n�!��̤T_d4�����HYД"5fުd\!�DM4?]04�$�,�Li@D�+�!�d�)_l֨#sl��5�X�r�eɬ
�!�Dcg��%I������P�P�!�?C�Dt�@�8�`��Q�!�ǿEO�i`�)���Y1��ݯZ�!�U	*�8�(���$z>��wk�U{!򄄍cr1����3TL�e�P��rz!�$Ť(ߞ���H��u5n��j��JD!�d�%$��PG��t-x�JTυ�W:!��+b���Ŕ`'p��2I3!�ѓ_8Z̸��Ba��%�#�)L#!�D�
GD�Dƙ������b��j�!��I@��qd�[�R��_9K�!�dR*�i�`�4`>��1�K�G!���;h"m�ք �^��(��A<l�!򤏳RqZ)SDC1zTL���J�q�!�dX>�Yq��6UT�Ր�+�,0�!��1BDa�6i�\y�4*�:'Q!�d�h��GD�kwR}�&�X�cK!��T��A��P�T^���pǒ�n+!��([J4��r�!U\4H�%�!�A�G�!��K#���Fe�]q��d\�W���87/�M��U��"���yr�% *E�)�2}�>��Ӫ ��y�Cf���s!��s��h�t(ۮ�yR��PM�R�'A�NDmQ�,�y�oċU΄1��I���t{Qc�<�y"K���RE�@�~; ������yR%^
	Hp���t�"�x� �*�y�_nm\�(��B�o��]Z��3�y��W�?X�UiM�]K�凰�yr(�4@u���ˌ@�.}�'�Ė�y��K15��)��Ã<P�H��-ގ�yrI^�ph��eHG?;�KV���y2mL�5�.Ĉ�6�����V9�y��/'����"H�3؊m��\��ybH� �!	�Hמ/���t�G �y�k��P��J	&�R1hg����y�ɫ)��J�î�⹑1E��y�H_#)HVH�j�.�&��B���y
� h- �Iʰ�6�8��
�/\L][�"O�)+c�Ѩw��a�/��eJ(P"O�����U��J��O�O��� "ORa�5���8"bH^@/��3v"ORC�̒� �4)J�g%['dء"O~=�v˗35B��r���~$�1�"O~�&Pg���q�������"O`�9b��1d�(�	}�x�(�"O@���+H�`p6�fI��d򅱢"Oz����ǮVŒq��'�
T28� "O�1�1�����%�< ��B"O�U�թP�)�����XF�h@"O.�Z��Z����E �����w"OƉ"�Գ�<	С㔭q"OZKǭ�� p�'�^�8����"O��k�
mւ�bV׌F�H��"O�K�`��+�9Y$�5e��2"O\�֊S)�h1��1��	�U"O*)�'-�0�Q������Q+g"Od Za�:G��ځ/Ҽfݶݠ2"O��r���G(`$(So$�\U�"O^	�eL�i�H)�0��;t�¢"O@H��%�,sB�}a��feR�"Od-�����l�L�$m����Yy�"O4��S ˮIF���¥'4Ԟ�J�"O���ǡW)���4K�'?m&��"OBE� (Wd����bo�
 ��y�0"OFz��5}o�%��Qk���
"O����[?H,��S��7��aiR"O� �)\�FtHp�F�Q�z�(�"O8�`G�C6����R���!�ykT"OD ��բe���1�,�����P�"Ol	x��S#gO�|{	�8��Lg"O�q
��SҀ�R%���0Z�D"O�tSC&�'/��h�ć����"$"O��X�J�9!^�d��f�W�B�r�"OVHQEX7ɞ]���84�y��"OP9��m	CĒ��8��x(�"O���@�b�d|@��&Ep5��"O���K֗&�0`*�KT��2aX�"O��7��p�����LZ�O1�,�y��A#�B@�Q�N�`'4�y1���yb�?��D�Ae�!Pj�=b���,�yrGG�>� X��I@4@�$�P��y�E� Rp�Gd�2j��ЇC��yRN�/Q<�(@BL�}���##琾�y�	œ?@p�i��
u�d�uÝ�y��mC�d`��U)r��U$�;�y"�.�{2&G�s��BcO���ymZ�T�:;F��*��p��)�%�yB_�}���ҁG�]�b�hC���y�G(~�=`��T1�,���!�yc@58�@33kK�^*��a�O6�y�,^�4-
�i��]���i��5�y2�֤.��1�  �VE��0�oד�ybe-W\�
�f���߶�yR瀮�P@y� F��8��	�y�N7t~T\H5���,�Yp�_%�y�d vI:؁��|F 4�feF��y��J�i9������2<P$��E�:�yR�֖r�*ܩ�o�/7YJtrU�ۢ�ybN�I.�
��A�2�I!@�?�yR��|ybM���+ ��*����y��@�E�L�rA ��Zb�0��l�y
� ��:B#Ѧ@\HH��E�(�vD�T"OX}8P(��_|�Y�l�Fh��"OR1�6Dؿ1�`��?	�:���"O䨛W��
�@��Y#�H+W"O �+V�R>S+tL�r!K�_�H�"O�Y��9i(>X)� ��)�ܸad"O�M�(T+9��͑qEӠJ��x��"O�,і��9H������P�'�m@"O���n�2pw� ���	�p	�"O�(��ַh�͒$I�'d��$��"O����ǘ-�h�X�J�'�^�+�"OH��!#A=<9��U��-?!��D�v���V�S�>�:��䃐�Q`!�;�N �卆�84�pE-!�G(l3N�j7`��7�8��f��}'!��=\J~��v��P"uH�͒�c!!��/S��+`��	#۬`k"O���� Н50��#!*Na�2!�Q"O�ĠR�D�[)� ��k��f��8"O�u��䙮?�&͑6 ه%�Ƽ��"O������iV�d!�
o��i�"O.�C��2�\	Sđ�~"OR��'�2���p�)�x�QR"Oh3��=���椔�o��mk"O��K��G�H8@dD��v�v��"OH|JSc�� �S�0MȊ�a�"OP�Ƃ�6����bK�S��"OY�3�>V@����R$j��1R"OnPk�C��y��I�R�PDS"O:�3��/ANjXs��؞D�(��!"Od�5�R�`p[� �Fp�8b"OdY���,2!H§ 0��g"O�:�iG�?:@CE/Kb��a�"Ot���JŔUT$����W��Z�"O�i2�ɚwyH!��,�TГ"Op��r&�jeh��҂G�S�D�t"O\���H�0|��t�g"��!iX�J4"O�t�&O|������ ��P�t"OH�J.�?_� 9q�X>$�v|� "OܩY�ޯ^0��I�ђ ����"O(}�g��vJ�
�ňUi���"O�d�4�ܺ?H�5D��k)d}�"O6���gǃ@�� �����P�ҡ;�"Oԑ��c�` �#gP#4n�9�O�7+Y.�3Ą�/��,B�C��yr��+C+�}��M�7JY��B�,
HLb�#	��yb̍65i�)@cB�7s��ِ����y�FQ�D�I@�U;o4�<{�=o�7-.�IX��~",��m��( -L>c8���K��y��ɒ�p�PujS�
�h�haHK*�M�����p?��f��[V��0gn�Yuh�� v؞��s��׫#�jɻr#�Ei��2��g�!�J�lc$9�@##�f�y�@ŭ(��dD{��S��y \�u��J0�5Q���bU��8�(O��'G�;դ���d�	�PW�%�ǓM"6�<S��YA��G��պ$G�r�B�\j�B����Z�l`00)��ʓ��X�4��b�0yaN�H���rōEA��@�D�&D��Vl:m�ܩ���W�_3 l��%�I����'Ez�%ꃛx��dyơU�w\`����V?��ȐZ,A2�D 3j0T���#�D�'ax�#�w��\xw.�+��HR��D��y�(�Z{�t�I�Um��5F��:�:�f \��B�I�6107*d���l�G���M��'��'��)�� �a�����`�0*��H�y��"O�@��DD?��0���	bX��飭��'M��A;���|Γm��\�����(t� i�D���I�2%�F���s�Έ�����_����c^,!�H�_U��8�-�9��LDx���4��4?J x���3r�-�WV�ְ>�@M�R�c�e�Mu��Ǆx}�iH��+nA��.Ԑ���F0w��ѣd�%$��Ȳ��rX�l���~��D�&��y�$V$_ÌL��χD�zD8v�	�hO�����P\���Ei�B���Šs�!�D��:���u+�Th
	�3��hR����"~��-Ć�8A V X+{�x�����yrl��m�@�`�z������
4 S���<���<�f�3}�4�r��8|6n[D��c� nZ~~2�P6 pZ4i��K�f�ȂjɥbQ��G{*�Z�Z�	�2�
A5�W�	y��"O�����֣Nx��+v�H�Kt��XW"O�����8F>�Cf$����q��"O��K�#:��uM¯4�ڡ�1"O�,���R�La~�{��H�H��8Ca�x"�)��MHl؇!���ةk��W�|h#?��Odc>9�iڮ0#�,rbؤZӜ�M4��蟠��3��B��跋�&��v"O ���%�8A(4;�'��;�\�	"O�q���&F2�ӡ��%>�c��D�Od `I$th�a��	m�0��'��#�S8j �Jg�N�swXyA�y�'lO��ȱ̛i��m���Q�B����OJ�mp���� �w;��`��NU�B�Ʌ!�����*%ʈ�Ԯ�.E����3���>4�ہꕉ?�,lS��@<�'�4@��	%@tݲU(�Y���$U6NB�	�T�*yx��E��f�k�,����tHE��Ŧi��	�:vJ �wAѽi�r���ȗ~�B���H��'�;CpD���l[�N��#>����h�0hʄ�&R���YЊTn���|��'�Oq��0Yv��.4L��G��{���F"Op�uhF�CH�p�w�J�$�<�S"O�!Z�O,������N�I��i�G]�������1��ȋ6g�'V#�逗���?���0�ɒ�y�hѴJ�l�a�lP;0��#����y�.��S�V�96.ݰ,jB��؟�yb�L�t��2���b}�ᑆ�y�IO$��� �M~k�)hAA���'!Q��$?=x���<Ho�Y�Mۋ������ ���<i�A4<Z`ܐNN��l�X̓e�a{�픜:MJ��Ѐ� :��p�s ���xBt�
Y��B��	���$	 cI�"O��I�FY:�T�3��#?n�s�"OX}bA,!:~��
FP�+�$�yb$K�a�v� a�,��lڴC�-�y�.A*�N��Tˬ+[RYp�B��yB� � 3FQ�T�
|K׍��OP�Oj��b�d]�8�60;*G;'m�%��@H!�d=%T@�I��'L��x2j�$82!��[(G�Jq�.���D�5c�1����D{���t+w.
:��k`,F-l��"OL�`�0j:�{D�u2T��@"O�ҶFA,�����ӆ�v��"OڱHţ�+c��#��"�x��t"O�a����CDر�P�Ľ@�[�i���Dȓ,�T"� � yd*0y�B��H�'`,8Ey��0r8���Ċ1�(�Qa!��y
� �!`O�&�`�J�әB��Y�@ᵟ��a�N�T?7&��B�=8��Ң�0%S%r�B�	6sZ�@�&��K��Ѐ�N{�B�I�^�
=�T���TF��b� �4Z��b��O�r.O(��da�ެ.�m��K�*R:F3�"O�a�ǎ�*+w�y�Y@��1AX��h����Z�t�Q�%[LՀs�Z�"?I��iO�G�"i���<6�mzf
�y����'��Du�~�O�>�!�kb�����̻&��jd6D��x��ӇwT�#�F�}�@3@ D�@y��~�8 QÔ3:	�)	�=���d��O���H7�]��+U��1:x��	�'Qh��4n�zZ��q��H'3Eq�'U��7Xƺ�0F�B�"�����'��Y��E�=���!����Z]��'b�D�Ox�'�S��'Jq���ŉE�'`Ż���)x�~B�I�#S�-{��%o����	�D�lB�2��A�R/�'y�k�d� �Of���&A\��뙄x���ㅇ2�!�d�7C�$;V*Wus֩��F:N$!�d���dz��݈l`Z%����:H�!�d�T��9gI)?O�����%3!�d N����FJvʅ�Q!�$״W�¡P�@�EG�U���2Ac!�d���ز��C�"VQ���j1O�Q��gP��i��hPŔ�$ĬT�ȓ_9V���̴l�H���:#됨��R��C4��h<���f��`V����&�	���Hn64�&�V7'��9�ȓr;*-��$X�G�v�� ,$;�]��+:�23&R�c�ԩu�  b�贄ȓODaq	������K�+����sH�z2ƚ#o�P (�'J��V���f��H	�W��8�����q
�U��Pn���d�V�n�\���J1�\̄ȓE�8 ���%_��$�³/�ҡ��hd�sE^�lXIp 3.0Ʉȓ>�D�&D5=tsf�+^����T^4�����h��M�Y�@H�I�ȓ��|��dK�*(�S�O�y�Ԇ�&t���� C���r�(� f�� �ȓpTxɺ+��|���&�|8��i0���!��
�MJ��	26$2@��|�0�s��yd���%J���P�ȓ``��G�A:e�`8�jT�(bm�ȓv�z�8��j�
�*�%�5� ���$��A�u�V�B�!��ONp��ȓ=�6�#��I���@2��!�&�ȓsr�4z��3�X�Rů��'�܄ȓij�D��c�^A�����\5v<�ȓD9�{wo^~�`�#fL�K��ن�<U>ij�C*QC"� G�T;m��'	`A��=cT���B^P��'��\b2B��#?�	O\|��A�'�:�r�ǫw;�a�J�y�����'�.Q�A�sӄ�����!��T��'�F,Hpe�Q>�yGeAP�d`��'Y��� ����H�JR�E2d�{�'�Z�5-4ۊ���*�4`#�'��RBŉ!#f2��PC^<.^ly1�'w�D�)�"(qEHD�\��c	�'f�4PAM�^q�]�J�!� Y
�'3h�S�g��R:��P��zP�t�	�'��ѣ�Z�-=P�q���m��0��� �4�=ءi3��8K�f�81"O����N�<�jUB��;}���"O:Qi��̿$e
�� ��Q^@��"O��S�۔-�uy�锃0%V��"O�0���S�jJ�h0#�]�s
�y��"O�$��&�u���Z� W>|�"O�M" ,!�:5a�-�./��,��"OL�"�G�wخ�ð̂�k�(���"O�pd�\,�L�%��yW���"O�(�JP!)ށ ��>gA���Q"O�x)��qr��jI+f̺Mh�"On$:���#4�nC"3k���"O�k�>񚥳����,��ԁ2q_�ݐ�O��L&��0�'��%�Q'_Ǟ�����x�5��'�̘�Ӏ�r�x�9)V3�'aH8ȴ*�,D(�rbڠv����'�µi������q[�-��h�l(��'������3�
x���E	n���k�'�N}H��%����F
E�Z�$���'�9��+�:C���ask�%��	�'s��u�0]E�Wˮ.�^�X�'c�3��^0b푃��#\��Y�'=�@c���D�A�cHєg*,��'t|��'�P�p�9��hS
�X���'6�2F���Z�K�0-'A�' �#��<�زA��'X���'�H�c��; ��m9oΧ.�>LS�'���#��?yny3�@_3t�Z:
�'�BB�,JLQ���2���'�t�s�)��@���zFV@xnY��'��)��=B=�i;�|���'u"����[�5%�,z�++O����'`� !F�1�v�QW��;v_�9�'N����O��s�5pw�)PE4�3��O���BS�R���d�ͪ:���4!�&p 6!;�l_�L�ڨ�	�NC��	�
5(��D����T���F}"���\�«��K���YN],OA��Y���%jRQFi����7bT)��xb�ђ A$m�C��4�e������y&9���7m�0�!4L��B"e�c�H�'C�Ƙ��W� ��!iANZ/v��ȓ$ĺ�1"�K��v��͓$t`x�q2L˝ ��Yq��	�6QrWF�[���ŸD x�T��<;ԍ�<�|P�􅆜���'/+�O ��G�˱G�ȁ�tbA�[H\"��C=��,:� �H/�1��'f�2�s�"2d��ēW,4i�L�%y"i6�
�̐�i@*�	6�Ð9� !K��|���@�A������i��1�29�B�i%�6O���co�<���,I'2��ҷid�`��ۊa@$Ǖ'X��Q�,ۘ}�����s��m�$����g��U���M�<��e��4��i��E�Bј�Y� ]�-W��:�
�Z_�da�-H ġ���*5��e�E���|+0���
����(غh%����Ʌg~@lSd�5�F�3qi@�Y�ƙ���	�A���va��Pd+Qd������ӈyz�|򨜂ьq�O2C��W�&yᷧ�-]FJ�N>��G�XL\<��*6/t��*S�xv�캵��i欕*jN�2���� �߃����W���#K�0y��4Fc>�O��۰��|jH�҄�KJ��@N=1�7ƕ(K� �čP�c�ċ ��~iJ�k��)����${Aa�t�� �3�⑓bA�3zݰ��',�Q���FYA��E$a^�@U�A�g^(�A�ՖTWJlBF��PN�1v�Â�\e)���$gP�7�	�1Ũ��Ƅ?s"��J�3�j���%<O*���*	�6�|���-Ųktp,aF�]*�Z'a�v���Őeͤ��eA�,q�R�+&H֢�TQ��Y>�:�n��d�|��qR�k��l�1$lP3�X	��*!��2�L�Pj��4����)֟A�)[�ϔ��@���#����0b�}K������"-ڵa��#"��פ[�b`i������
��G%xd�Q���m�uI�� �v@ұǖ�o�����Q�E��-jAF&n�Y�F�l�yI$�ܣ�l��C<J�;@�� ��aQ��h3챐��[��H��	�G�H��f8hn襱��\uԴC��
kH�۶F�[_���%�M:B�Z6m� t����kK��a���	v�ڸئ�^R��Y���`��Iw�Ҭ�dЫ��*РG.P�2��ïMzA����"`�:u,�+9����7�+���@��W�<�҃�xD�ba�XG�=�3g�ԝ���_Q���by�@���L��,����M/� T���-Tn�v������D���T�+�^)�vϖ���E�PJ�,-�\��͔m�f��0l<��(L����jA�l/��P7���O��D	P���b�qk���tI�N���0����h'�G��I�6���*R.:g���k�~�`�)��^��䋏�:i��
`�^�{¨�ϓ*�*@�*
�1��^�~����B���7�Q����A�w�Y�.�<-(ÍP/��PMߕx������N�d�/X�8>@H@�`�\m���'2��B�e�+��$��g߼_,�@��~y�d�2i{����E
���@��cI�0����S:�p! |]@F�0lr��z7%�b6�9��'��6X�)�鉨.Jx�ۂN�3�ĂC�)����D�:*��j3Ö&/^�H1�/��ny��0��p��e
�d�R���GZ&���cW$*V�la&o%�Z��h��1�:����@&7"�V�_�U��&�Y��)�$�����p��onI��ZOfT``�k߈Mm0�z4�֐*id���C�
��T&�,BOr9�B�*f�5!˓
J 0*i��m�i���/����pd�����V�@+�hȒ�ɝM,,q� m�y��Ǧ!��AȅD��(��\=-j`�YF@J5�F����(�=��8��|��ĺ����k�����*`�����~q6�cp%nA��B�iR}����>P��!��V�m$x��U�x} �K@Eۙ~e@q&��l���@E�'�
	���te�e�6V�aR�@�Q2�5�Q/�6\�đ�c!�4A�C�zq#��̜1�2 'B`�2WB��ӮO�q�����X�D���o]Uy��Y� φܲ%�D���CY�C'�O�޲� sA��"�h �E9v蠑ڍ7buKb)�"@]�{wa�ܨ�h�!��#�d<"��i�h�E�)]. ����v�j\-C<�q�b���@�`����'0%8��(z將)ۗ�Ą���O8��bb~�ya/̸)d5����) �b� ������PX-�ǳ�d��^	7lޕ $�@JGp<�T"ۥZ���>�F)V�x,̐9��) 8=�q���o��	�c�%��eƣk �2%ւ%v��)&+�#jYjʓ[��!��/E��m��Hځ8ːd�%`Htt��jt,G�1#J8�vE��j��QDj#j�xxZ���j^�d�V �@���&�G'3%D$��6k��I�]�o�dTB��IBf���_}3���.S��l��D�<O���w�$�T�i������>K���g�|��� f�>�!��!���c�B�O�,):�c�+dF�Y_�!�D$f��E��Ei�8���^	��I�n��G%�,M���y���RȂf� =z_4���O��$*��=���zlxE"�6܄�R�Q���h��DY�|����7���)��P�B�ѓ�
��O����6�,�D���DC����n!��O���'��iQgL�#��E&�[�n(��Й~� @�K8Z*2��$���i�:v`�(9�"�˘'=���ebBI�����B�g
�\���5��!5�t�9&LT�7���x�H[�A�9#��e�Pe8(�!���At!X!��'Lq;�H�3Eaޜ)ǎ�S�J9����*�dX3w�Cz�pj��UMְ�rG7uʸitgN$S�N)8�$-�d�%���Pa�>?�(JvW�`�09��	��$0�C�Ƞ`bM[�R�&���@Qh�;1�ևV�f�(m�j��pv��\�P0���O�&�� ��c<ɘ)���P�<�5I0��t*0!�
g��,�>AN8�F����`�eGDǒ���Ġn�Zph�O^gX~� �'?CP��{�x�2�D�aI(�֎Ė8���u��;;�	@V�2�	�:� ֯�"o�Xp��o�Uψ���@X ���TBf�����[>R�� ��s�B�&Z*-�N��3O(bGU�A`����mœY8\�;Ơ� �y�$����P6Z���B&�=`��e"q�L�n*
u�u�	�g$f���^d��-@K|%��x�ū��@.vE���*(�z�a��j�
��2�Kp���2+�0C�u��@�/tE�Tg(.�1O( ;e!˺&v��X�h�cG��*0�òR��+�G� ��� &��-).%AJ8"~��h�`D��
p"�3W�M3���:6j���Qg�:g�,�{�`5���K��߭q`�{�{;������5V��(! Z�%A�S��Dۂ(�=�r�b�Tx u4-�&��!���U��Tˢ?���R���<�n-�b�,,~��qJѼt��b��!�Ѿq���;A��0-@�R���c׊˼�h�KV��<�2�f�ɍsc�Zq�H<f�0x�C�e���p�fO 5��s&H�6?�8�F�)�iІAGh��'�.L�jT ��˘G�� Y��8|?����IF%s�����BBn��c�/O�zt@�
�E��4�;���`&{��i�
��o~�q������4�� 0HC�γ���	�]T޵B���`	�@61�ba��%�(bW2�Q ˕'�d#sϖ�^U֑V%�= �D)R���4�he���5��8�1
��gk`�0D^�m�BQ�	K���G{b�ٛ�(�w,��T��d�BD�u����w�˱�|��A��IBtL{�~ҰCa��!{Ѝش�F4v�����-�3�v�WaLNbd3���4�u���|�l,[t����'4�=
3�
!�P�q�m~���Cؠ0q��@R��L����S(1c6�kR	ߧY������,j>��F��!��A���
	Iʄ%����*5d<�s��&[�����Jlj\�P����)eK��g'ν��f4� d��_3U� a*��݊HhnX�`o��k���c!�������H`HA��"�9�������)I�)�P&\"��A�����F{��5�^lI���:�P	cc�'!TH�+&y��3(T35<<Mk�4�ZX!2g]Ҧ�r�&%o@B��V�L�/�8%*ybH��c��-Z� ��.�Q�F"=b��3"��	K��,k�\iG�b�H"E)K�G��p���Q���Qf�i� M)V��h��#
�0:�,��jc�|��f  9=�)�3l�0�8�
&l [��&��'n kb��"��� aC�r�B�H��@�'ؕ�;E�*D�K�xg���`N�t�δ�sDM��ĊGƙ�
�,0Y���89\8��k��}m���0p�ژ��C�?iTe��_�%�P�C�Fڸ���I�%B_�3g:|z���N�tb�O�5� �B�BҪ���	 �B_ ��УI�C<��3E��7��Îٺ
5� rc��V�(\H��,4䈱� ��"F1�AD�Y�:3��
?�p5�fܜc� ����� ���ɗ2]n��F�P ^�8���9�l�U]�M�˄:O�,���H9%��/4�́�˅8K�<���(�y�'�q
'�zF��<�t�G��p^�t3��<��!L���)�eͦ2tn��7o+hz�1��iHuV�`:CW�z�(��f�� O���]p6�LRǕ��8�Ĩ4:��O��Y��ny�	)��GkB�"|ڲ['/9�!��EϨ&A~����E+�I���/R�b2�Ǻ?�Z�
�/ۧ.:�9�rEΪ"Il��s�ĩ��y�2o��Y9P�#DKN�&��uʴ�@����%CD�A��aڴO��� �~���ɰu�$�[pA��q�rA�OL2svT��"C�]�"}��gJ_��{�g �K/8��5ht�h���0v|�O��� 00S�DZ&t���Y�AF�}�z|b���21F�I"Ǯ�1n��)G&"C.s�D&t��yca�y�h`R�C35L�y��fL=-�l��ڕaU���L�b����k�(��'Sr�0�'J�.ɾ(���3>�ؒ6��zƩ�A͋H���((T,j�k�w!d`�b�&=:�!Bŋ�)/�4�I�F�)q4y�#�\ Q���X��e!6�W�(����F��N�X�O�������J�H�{0�P�aur9I���g�
1>�2�G3>�B鲒-�Du<������f(��
��(����B�40�ba���8�V��R��5�"�*L(6 �k���lH�)H�w����bB�^���J!�χ5����7/��n")��O�P�DD�5�B{ƈP���B�x ��YQ4����!w����C
Ԡѕ��}˞�<1�h�5M�0�&̐� P=[�eƚ� L{�H�k�ŉ�bT34_t�ip��B�4�6��B��03_n�!�� �/�(�䊬6
�D�Ŏʰ@'�ݸb:F��r��I�<h��ZaT����݁B
걘��`R �P�Ԩb�L%ʆ�߉|J� P!D��^�B/�!k⭀'ď�b\<�0�)c�J5�����y�v`)���h�yb��]\� 8�}�c��l}�qE-¬�c���KA ��q�ƈK�zG� ���h��Y��p�𔯉"p��ⱀ��C��@�)�N��<*�J��	���V�ݠ��;_���A���G�fI0!��lU��5���?ad�?5x�k�1#�sr�V>���fT�#�[<�&-�t'ؓkeX�)A�fإ��@�:II8�Ƅ�WrH">a`��٪�!VEA�F���Q�%��Q��[�?μ0S�P8g��h7`�&�E�l�6�Q��f���dY�o�~���+��C�@�à�RN�����'O��T
����8�6=����5g�**!0�S%k�\�|�����^~���bB�S��x�U��=±�v��5�O�??DiCw�N#�,�P�G|�����$�.D��EA�'?���d#���'R��`�X�e���I'z�n<q�CɹV��h��%��]4�P�w�a1��+���'
Z �<Y��I�0�XxJ�*�?�0D	f��w	��P�(�$�"��󍃔a�z��O(Pu
�GZ�-�8�`����-d�ED�?f�		r���<~���s��\C��C9�OVh���\�.��@� �Fj0 6���5o��i�1d�� g]FH���y�� *��z��@�X��;$�Z�j�h&��攖F�\x��I #]ּ�b�Ј)C^��e�Y7&�V����Ax㒁��m{�qsb�տy�Y!�`��,���瘶$�R�'>,�y�Mϻ���r
��2��	���;��'C�aJD���8�@D��JK�(~���6�~�C̄]��d���a�2��b�F�:��D��h�����/,d4����OV�f�ܓa��<����N����ŝc~�I����l]>@� O�{��OQ,`�T�O{�R�V'P�\�>�jeٮ-_�E('���c����m؟P�F�M/+*�kT�I�d��AEj@h����A�B݊�!�!X�Q�X�V���)-�;č���bE�wm(�v���K�Ӕ:�� �DU��H���ZQIy��(�L�P�v�v!��j=X⩛�@�����d�3C�X1[���!Ĝ������r� �d�N�:vh��K<�!1�~��W3,n&���Z�WN ����H�<q#N2�.��.>$ɾ=��7��c
�%�&��BS�yD���&�D��R�_�&�>� ��E��|�ȓ):<�R��)]i�᫷M�z��q���OH�j�_�iʰ���(�Q��9�KD1~���Ծ�R,{$%[xx�(k�9;`z�0�`%<���U��7r�j|y�"E; ~\�S�'�Ȑ��ψ�*��dR���%������D��s�EYM(���L���.�%ZH��a\78����"O�,*���"W���V�b�0�D�Oj� �6�M��}
�H.@~~Q�sKƫ_�(%c7'j�<1Ť"G`Y��cT�B�iB� a�	
B�aJ��'
2���;C3\LC��*;g ���'Aޤ��l�	3�����X!��(��'�v��&r�ܽ�
Y�`Y����'W�A��J��G����)�Ժ	�'���B�j��/��`R�ှ���'��&�Ύ��0�D���z�`�'f`�X/�^���3�I_�>��'Z���d"��v��ӂ3WJ��J�'��pꎤ7�@s�G�M
�P�'���В�׊W�t���G+~�p�'C&%�.C3-.L]Y|�٨�h9D��b`��8FU�(y���2�p%�/3D�D��,�%W�eJ!�,w��W�4D�� ��S�q�(�`���Jij���5D���f�A6j&��CFX"Ҁ ���6D� U� �I��P��	"`8Dx�R�7D��d&��V�DE�5KJ@���2D� @� X#yNqhf���d�<�Ȗ�-D��
�&�kj�d��O1u,��W�*D��A�eY56811aFlS�};'�LJ�<Q%�](Yj�%i!H�0.�!C�`�@�<� 6�a!����*�)�����"OP� ���H6-������I��"O>��u/���e�w-P�B�n��"O�<���T�Wn��r��0�"O�	��UJ��haU1̐���"O$���SV��bh������u"O�Y��J׸Lق�yGl=^���"O$�cd�Ԟ7�.�r��Px�s"O��{2��_���'*~V�݁7"OfY�� ,���[B�\2Z���@"OD���c� b����^.O��5f"O��!��>ȼU �FA1�`=��"O�H�ż7�9�\+j/�pY�"O. ȆLR�*>,�"A��8��b"Od��׫?o:�!�$��"OBM�Ӧ�0LL0h��J�;���`�"O���(�
O����΁(o���"OL��\�p� p�Q]dp�J�"O�H�lU,8�qbUZ]��c2"OhA;1d��j萜H���4D�a�"OL��CjA��(�� Q�3t��D"O��5�4z �A��U�p��"O"-��!ʣo�1	�.��j�p-�e"O�PZs��+I��`q�m�%8E�i�"O~0�@/��eQ�k3����"O$�{��د%0b��T��^=�\��"O�i���S"2��I�{;̼��"O���Vb��N@0�b����d�A"OM���D�O�V�Ɂ*��h���v"O:�X��I�"���3HL(s�A�"Ojl�DbG$���WA��%�����"O��R���;Zеjǡ���ܱ7"O\���N��7A�$I�NY;t�L-��"O-�7/��2�x�{�/X�3����"O�A��`�5���10�җ��p:�"O���Un
�f�H<�OV*�����"Op�*���!�	�$��7jJ"O0-b����8�V�K/"UԤɂ�'2%r����P,��ӵ"ÀL(�3���6xL��<\)6���'X���"qa�M�K��(B���ʽ/qf]	Waц��|��+H"uZ��ݎ5;�e����"��)�!�GüC�I!�DcH�=��&*�#P�z�	4�<X؀���n�(*u�#�Hs�$F�(]�&��2��u���T�B䉆)�`�rq��6uc��ѢM��]��t��ꆩQ�uSW�]�.�ZP��H�|2�-ݙ��'�D�R �V����	��-{���5C�I�)@�P�T	��q���R�Q�����K��	X�a	-#��T��2�	J�(�8�E���Dzbe +`�X=�$IF�h�d4���AS^�����2��|x\"�+�\����L�� U�[ �4"5*�!2thmZ�A�PC�AC�T��$��(���I�j@6q�k�ٌ{Ŵ��ѩ	td̙�㎃}�!�$�]0ݨGC
�T���*���H�����~=�`#U,,D���)!,�\6Ͱw�ʷP�ƒO(f��2�\@����B��(S�',*Tqv���ft����	�]� ��#��Z�\��K��\v(��/�2h��o�/�t�e��~�I�.�
|�EW>B&)Ҕ.UXgf��>D��(�$S'�(l�P爡g�6a10���pm,U��N't�,zvIҧ=h�,E������ݸ\�j�"��5�q���P�]g�g�	�=^NL��c�B��vh_�g���S��Y0d��	d��yra8T\l���M��O�������o�,'φ^���*bܾ��HA3s ����P?V����M�c�4�!% �N ��[0�;��pR�ȒW�y��@�Z��0�'d�0�1��Ǧ�� !6����!	��ޑ���^�F�`��	-����b�;E�
|#�L�,1�n�;�HҷR����"Bh�Qs��;�>Ac�H�:'&b�d4�~�{HS�T���ȳ�C#���4"� ����X��:vJT�R�d%���*�Q�L���X?�Yp� \-`�J�I���$�.�����#G��,,���/ݚ\Ĵ5P@�0p!D� !
�ʑ��O�Gx2-y;��&Mǽ+��b�h߷+�<���C��c�~ȓ�]�5��}��7��0m��*��R�h4,�"��Jb)4��&�Ɩ?��)��MP�,qAV��hWf`�C��� b�B���2>�ڗ�,7���:S	�+e�x�YsC@�oj��	,0�h�*��ihjX5/L�]j�ɱ�RT����C�/G�!�������pw*�O����Z�d�������-+���%[r:��A�hH
�@ �b"IyS��@wc�e�����K�.,���Ge�p?��i����^�EqK�6~$��t�.�>���4��X���]���iWH\�9����4�Q�2f��=���� ' 1#!X+k���W��!Y��( � @7�q���I^�	� Y���!E�,� �:�`99�N�I� Z ᒬ. ���s��"Z����/�0�z2�;<�TlcR�C�1��6#��ba��+��`�AQ�&S�I��+�N���ɽrB�q�v�ߕp��<�$�y�{���&o��Q�4'ӈpJς��ċd���.�h�b�&�*<�'�� ��A��Vː�"�aU l���'��pwl� cX�(cw@�����wi����`�2vQ��k�}��y�� �<kg�P����GI�������"�0s�1�U�A)j,���BZ�4����1�I�0Ē�jP� 0x�	񍈘S�Z� #��.�"��e,o�,P+��͓L���3��ڟ���Ȃ64��$��
8�6�����.j�<t{q�,�dNw<>�S�ɚ�h1�@8�:J���&~B,qK�MG+:�)�	��~t���7�x`�B�w�4�anG�\L��1�M&Z���&ǵV\$��E�K*/�p�!ď;kxP{�TG�Q;�����Sm�8(�d��ww�P��`�2
&�` ��LP@�Mw'�4��`"�Ǧ�A �ɳh����rhG6Dk$9J2J��u��mA�:ʓ���bHg��Lb�$�$l��M�"��x[􄃷)Y"1�,���_�b~��QA8x��j#� "Nh�a8�\�������"7� 0�Ć�`x��@��n��䊓� ���#؛a4�8��0+�:��0 �z=��I1&C2x� ��j�����Wc��k �x�G�1)�2��paݘKpz��d��\��("�:ҁ����lmz�R��@�+b��0NM'=7�����z≕wxp�Խd�.����+�L0�� eZP�;�+���z �� sr XV��e�4%� !K��P9@'�/a}�I"�Է:���K�I�.��RF^&�^Y��������>��A�$��(h��z�|�c��BB��@IҎ9R�1w��!?�08��
4�>��qÔr�v�-A�BA��XC�:��\)����Iƽ
((�6��'0�F4z�kJ����"%�$���o�'���+�X�d�B̆Eh��&dH6�U�.
�*�n i$ hF�lp�oQ�=�l���F�E d��Vd	3�q�s�J(�f����+O�6%P� ��k�R��lU�-μ��4) !,��j�*)�\���lZ�L�8=x�@R/j�T��Ԛ*ź��PE�5Iɖ��OP*qu��xp��+Pne�4,�*k� �g�_�H��Ѕ״Hʒ���g�I���ԩځR���)e
�9a��hzP��@��!XekOT����%����(�hH�ʓ��@�-C��?8�"���)73�6X�s�G�>���!,S?��]k�	�>_v���ċ-<��	�,�d���h�id�q1q)�QD"	Å O�3�xXP�晗�:�a�D�1_	�l��
��B���3��dbf�@o,�0�ƆK�6aQ�G��eI8'�	�qO �;�f;(h�	�:v>�@#ûr"Jh F#C% ���K��I
����G
B�?4�m ��9^��� �z�4��C#^'���%I���튗�:>�q����U�'���(e��*�-,�lp�霔xX��S1��48�f�Zs��A���t���"��R/K�$aD0S��yh��c�f�̜Q"&7�������b5^�A+� iH$C���{m��&�,��e�	Z�Z!9~����|P@��u�+���{a@�<���
\�B�ϟ�w�qA�z^\$�AJ�����fF[�Z��eC����8S�+�il�e��lv�in�u��l_4!Z��aj�s��]cN@�NCv��o��[��pwJ�6����D�)�u��%��C���NE~�� /�R��X7J�g��|3��ԳYy&���yH��<	 !�qX�1vhɵ .B!�g�����ןHTp#'�^ܖ�u-T�\F(�r��6wp��ȨU�@��U�B/!Xt0S灔_ߒ�:%�?_A$�R�1�$=�hE�B��95m^99����ұ<�Bb���S��;��N/h"5������\�u��%eu�СT	��D�ǝ�|�$�`@��q/˪L�d�i�HV�B�x!!��ԉ���^̓P*miCI[K͢J"�U23���@�Җ0����dl�!vP1�o�	Q	$}1�iZ�LĲ0
B'�23���`E��K��9+a��Gv9pt��bf01�tn�2�p\Y4���Fe2�$���A��U�l�$�5欙�O�8��HC>g?6I�ƕ�a��,�*�1N�8�C�Ӕo`X:��
2����B=a:>Y�6�!b��0�T��ip�Q�A��x0�ɐ�D7 b�p(�)��A;:p���6 !@�M&�1aD#ir�Ҵ�T�jY�����M
^� ��6,ªO|@��veN^�Ȍ�e�.l�&���G�i_􌹵�-�Ϩ<��Dqr�Ǡ*(\ȣeI��?a����J
�!
n$��"�>_�M��&�+?��LqR�ǡ)/L���IQ�=f��;[G"�������c$*:A��T�5D���U!�}�^(��Q��鉧	����EL-u��6N�-aN���A�?q��5NTD����D�L��#w�ʚ]�Nuq��
�fE���߾��9���;B�~!A2j��	��p����Yz8�+����]M��RG*�.$�,d��d��f�,�A���� �z���;6o����t�ŇD6�ʜ!$
>Hkq�A�5ZyD0qs��@���+«�M*h4�Ҁ׺
<N��KV�$L���	JZ�tz!�����y��BE	]����̇.��B�G�H�e;�KBX^I�"�ѳ,W|l����5w�:БU�+�)���F4K�i���ZV]���t����:=9FE���-�䃝+�Y���`\fq�@�QK?کrP[�	�Q�喆�1�'IY��G���)B�T?D�p�� Kv8�
@ڂB�C����C(�=iA!Қ)�N�;��=�����$B5*���	�?`.�����=zK$\#��(�T�SV"n�-�/�m$8dsLX�4��	�(G1![�W`'-ʞ9c�^����p�#ؑ.~���	Sd͚����,Q��@EGB�^��u�ڒ9#��j�4����Hިp�(YSb4Y���q�O����RG�7 P\�ՠD	v�Hh��i��&�9�����.��"D�@G��X��a��r

��!��	��G�A����Â5ޖM�`�|	j��S{�T(F!�nȰY���N� 4%z��Mf����.�����)
ϦqbN�3
���ы�_!��PL˃"�1�@�,�6�ٵ�p>1���7�ẁ˃^.�� �I�_���R�F��K
��׀Z��%*��`2��ԀX�t�a��Z���FxRK��S�]4(Q�['q�n�h�x#~q�僓�}��i*�-�
ZH1���Y1 A�hڤw�x�@ش�����'ۄR{��!NH�E�Ĵ��|s�Q��x�'���)w]p�ҥ9E�Ӟ=��2��	~V��Q�"�sj�P�N�a;���E�#�%���G�1��bfI�|Q��!bZ�
ud�`��p�� ���#Y����l�?(L%�#�x"���7wD�"���3*x0��ᓎz��ـg�9/�j�a�<@`�'���|���֡4<��#��y��՘Q� 8+�z9��C:KD��/X��l���Z-H�  �N.Y 죐a�-��ɪ�J@¦ɱ�����Ӫ 
�Ѫ�
�,p���B���zS�J8�B�	Z�19���3J"��a@2+½�p���G���*��U�y�������fE�y@���,݊��w� �,��1"��.��R��+����l dA�]8�C/ۂ�������TD��g���Y9���2x�p@�D7Nw��P�Ď�3@��ꎂy=j숱 �=pJ-� 1������8%�c�U�d��I�������#��8v@!;� ��4�ڰࡩ�98)�����T!j�􈤂`a��7k��'(,S��5o������ i���~2�e*�Z���Ͼd���
#�H�4V��!��NW��{v�ح3���ߪ�J��厽�e�W_K��X�U#l��w��3W��K���a�ņ�1��s!�Y�w�@��a��8�"�*�D��:Iƪ�)�<�ȃa�"!�BPL�:^��q���TX*�� ) �ޥÕ-Q"�A��e�� ,�<Q��<��X�0j 57��5���Eh��k���|#SJ�#+�r	4H���\� j��5����Dl��`OҝY���:��L��xؑ�.O�4�ٵ*R8ў�8cK )|r��C# =Ix� �'i!u��Hq�
$eA7��x�B8��6�����7v<�0�)�!w��T3*�&fM;g#ʒ|�z��`ۂ[{FX�"�eT,
��$���H��`�k~�1QE+f�>���;+�v��anD'Y1��(FR�	Pn����֋�ZPꅣ�g�25�P���.�d���E�\;���	�d�
��$(��k��Q�C��T~�p��Q�N�H5��^�>��g+"@͚=.t~��A�N��!
d�T N^,�s�J�B���y �L�G�^)�D�C�4;��#*[���`���b�';�u��٦E�ƙX׀��.�X-��4.��-�$h:�
8�e^)�h܃r�Y�O�ؕ3��Ag\��JP�O�P�Z')L	�<�ʶn�k��$,Ůt����	�t_J�#d�'d f����ΝM�dH� c kj8�%d� ����d�G�8�-�v�@]H����.�d2��SG��&lt���d*� ����gY>b��86(Y����=a	���'��Ԃ
0/��MX�F
b�.ڕ���*$� �BOpc"�h��S"X%�0���J1,��eDyB�/[���R�蜕 E2\R�%7�2��em�#��y12�ä^0xh˟��BDHO �L�Pf��Z������O�~�|5p���b��lz�X�}!�`��CX�HKD�{3�l�f��K��4ӡ�H�E֚ň���5lɤl�TM�0�h�M�ͺ��Z�*0UcS���5^w�8
�ş�  �B��@+>��2
ۓRK��¥�?^KT5 ���632�A2��1N�j�勝~0X;Y� I�����5Y����ô07�I:H|��/b�ԻŁ*�@ay!�
�h�Z,0�%��'@	Y� ���*)&TM�$�3�+M�RP���9JA�5�I�E��D��E�h�䌃$��	R&�Pz\wQ��J�D��w���"!���Ys��-FHd(��+ep@ٴf��� A0��Y�f��Z�$���Tp0W�
LX���ԾP�����?!S�ō{��4�U�Ȥ¸%�(D�0^Ԡ�i��Y��dz�l!�P�3s�z�� ���	f?1����j<�O�5}�L���d��E��d�Ư<|O�p@�(˷n��r&�Y�Spyx�K�AT`1K'a��;c�i���V��~K�PiHW�Kp@�JFE���O� �0�4�0� �E*%�ꌪM?ə4e�O/���Bn&� V�<D�����uj�L:gV͠4	�ک�F�Ю6��EpuÒ<쨟b��(%�N-Q�l��F]bA�G�)�yB"L�m����L>,��Ը7�'���/td�}��ǿ]��T��(O����N,�lP��A�1k����d�'����4�ЋM�,8��K"wq�� �)(�a�²-��%��ɕ�8�U�$0!.�"8�j#>�`��������8����#ù&P��S�<ք���A��h�F�)c����go@>GR �0�J���?z�ӧh��53�	�1�Z���"\�<yH�"O������ ���	 �?ux�it�|2&?tz��剆 ������T�F�ig���P)�C�	-i��u��+ tI���i֢C�ɺ������Q��ԧƇNR�C�	�dU�	Sp�W<����Ǫh��C�I�=�欒�&�8C������B� �����*�Gr�����Gh�C�ɾU�Ƙ��䅹"wʡWi�.*�6C�;bd5�悜7���3C��.DC�I>9�ȴ�@%Ȩh��8���%�B�I�NwZ�p+O�W��� �n�lwnB�ə<J���
@:h�R���)K�B��F���c��S>V�KbBSl3�C�	���!�ϩx�����N�'V�C�I80�&�0vE� �$%xga��f��C�ɀ?��h1W��2qݙR*�`��C�	(R��ܣ׭2.9��69��C�(�0����|�0@% R|C�)�  �3�H���hH�L	��y�"Ou�&�o�.�z��@�}�5�"Obm��$өe?y��hX�;��@�""O�yI��rN�!�f�/��4s�"Od�㑬ֿ;�<Yѐ���|JI��"O�Kq-��� ���V�P�^�3�"O,8�� y�*�J�/p�2E�F"Oh}�F��m��pj՚!�t8�"OB,��)Q/7i4i��)[U����"Oty�3J�F_�<���4#�:$�%"OZ��׆��`�]چ��<<j�|:a"O���qdB�J�����\$B<P��"O.��S�)|�s���P&��q"O�9z�Y� ����a.�?O>d���"O���H9&���쒡fz���"O(�Kw�؏`�(ǫ���di�"O����C�����+�7�P��"O�xũK�qR(lj�h�rZ"=��"Op�zj��l�Y�] L�ԉ#�"Ov5�码��Qy���i,T�J�"Oj���d��)��$���EǮ{�D=06�Y1	C�,���'��@��M���!����a�����xR
�C�S1�|��4H։Rh���f�� �hp�v���d��S�:!U�3���l���1��m�x��U��oK�7m��=5�
�m8���,F�t�(���'�Q�r��M���j�i�2I�'����I��>t�L��� j�>T�Sj��X}�O�R�
_>e*4�/i��]CDd? IPq� 񤈠
$�>�~"�jH�*]�p+���s�:�ѩ�@}��_��b�"}*-S�0��yX��V�uP���E2�0��)�G�S��M���~���;����#D��*�����WI� 9�?��,�$]�t���M�?E�r��AA��1Op��aAM�Oh�S�Y�$!����`A�T��Ӟ**�O�P�p�W&=T1O����ie�Fs���d�6 �z�K�_�0��.�'�c�"}�$�ȹ!�V�!b�LU ��)3wEm�A��6��Ӈ �2����Z:f����M��E��y *O���O�O
JT�N?ز��<�%�%�+pn�Hu̵��1^�(�55�SⓉL .=
��!#T�E5��$O��� �)���|��0IF�_��Q�0�5��Z�@Dx�O��c��Y�!�p���H��L'��eV�x�2�NP�S�O8d��	%"��в���%�r��� f?A�Op��ᓺMP�maFlA8bF���G�Z+X)T�Is~R�릭X�)*�jI�-�E���8lBUӶBZ�OH�P��Z��܀��O�yJB�"���a��'l� ��
�#������|-J#��c��>��תL�]�鑆i�IH�e��<�gZ&i�OQ>]Q�����L#*�'�<��	(D�4�L�T�������p-���A�&D���C#��>����c�\���R�n$D������$�4�a�\�bE$���.8D����H�P^�0�`Y�>��k�I7D��H���V��QDð%�01S�H5D��I�!N.X�E�|���I6D�h��#�+j>F0c���x��lрE6D��C &Ӳ|'A��M�V�j "4D�PK��q��E����0�0�c%D�HH���CH����o�-NU�mR��.D����M&F͎�ـD���Q!g�(D�(�3,��\b�b�jZ�<��X��,D�ԭC�e���#C��"nV5S!�'D�<�2Rd{0�*� �!\肶�$D�Ti���Y[̠��� Q�d�Q� D�4�F�Q�(�x�zV�I	+��9�vG>D�������b�	�jL k6���2�<D���)�%���r&&�gL��Gl;D� Cu��&@�-�G���|�n.D��  �{u���U�p(��MS- ��"O܌��b�TbSGY�p�"O�Y	�jh�2�Pf�i�(��"O}2��+O-<�0��@(4����"O��`e�+�b���,	-rhΔb�"OzT��l��1�t�k���xr|�AU"O�5�ᑿ@�A�b�bMb�"O���-�0����h/B���"O`����O�Q^��#q�2tD1�"O.�s��!|�za�O>+��H�"O��ꁎ֡ �L�ir!\�5 ��&"Ot|(�DI�{rZ�C	�j��s"OܳA�W�:��!�ݹ����"O�ؓ����8F��`��Ց� ��"O�����%�rh��B�e�V�"O��qsh
7vX0d���L�K��k0"ON裇�
�AI�y�d6OFڔJs"O�U*&i�0l]�k�d>m*aр"O�@1AM��� 1Dןfj��ag"O��3��[�����b�F,�,�0"O�D�rM�J�I7�w����"O<�x1�E�<Ä@��:�A)F"O
��h��:h�43�%�7�K(�y�u�>Q�4.�Y3hi�r���y�Ő�L]$�k��@�R@��
w�W9�yb�4*�BV"�C$��BV'��y��I�D>����MށFJF��!,�yBF��/���Z�+U�F�B��eoM,�y����=�h���Q���0����y��I�M�x�`�X����,ǀ�y��'d�ď?](Í��y��Y�z�\����,6(�I7���y��\�?����V�~G��x��y�k��5��A�t�3kXr@�'����yҩ�>�HՋ@�16�MxWO �y"A�_���`�T#.�Vf��yb�\8�<PHS�J�kzT0X�ę�y�#��A��d`�c1����̒��yQ�+�l�kPM�r���t`�1�y"j�����g�4hr8D���y���6A�l�X3`ޔnhR��
�9�y�[�0Zxc�c�,jB�|��n���y��I��L�	eL1dN��pb�H��y#	
jozt�#ȵo�
hJrヤ�y��  L���fǏ�`S5I�̆��ybn\�]qp��� B'Zz�yc���y�עK��)��M�R�h a��C�y�)T08�TP��1Q)��b# �%�y�.��r��-\���!��y��N����Ѷ���HQ� �yr�R=|���k1*Ns�:���b�4�y��W���k�$<yj�p�E�y��ǝ'2����� /?���d��y�F\- ��	R3NN�:�*��w	й�y"�-?�a��c�b6��6�H;�y�%��+�0�3*�/>8��%�Q��y��T�+���/ۘ�l驵,�
�y�@

b��5C�DL��XZ2ɿ�y2�/8j�ѤG��Ϙ=�q,ӆ�y҉�G��H���{��9)AK�>�y�*P�n���r��2G�\b��L �y����gO  ���l�(�1�K�3�y�� ͐���@�VULrփ�2�y��<)�HJ` K�7���
�%�y
� ��"�S1 ,U�w�#Q�"88"O���#
4L�k��Rz��0�"OB�[�Ɩ"*�@����#r��8G"O�T� �7��}��@c�X�"O<�IU��-��Kr���a=�Q�r"O�� ���JNvL��)��+̌�"O$��V�ʯ�P�؅�'~vL��"O�9�E�����ڪV�t	1"O�(PR��C~�xI +o����"Ov��ۢr'X��V�qȚ��R"O��ƭ���&��F(���i�"O֑#�J*Tz��� ЫC/���"O4q�d�I5���msށ�"O��۵�8~R9�▚=hx��"O2��`��6s�,)cW($N�2�"OR�#'�˸S����1��(DBX!x�"O��u'ŀE�4y�Ь�;}$m��"O"q #�O�P��H@�kĐ$�[ "O�����4n*�	0��zu�"OҌ�e�n�ʁ�!IF�V�Թ��"O|���9�X�ȓ�UW��ؑF"O.�)d���F��䊀	2ܦ4re"O�8Wd��4���PG	-�`��"OԘ�J�0T3Б����/-ʀP �"O�!���HB�>��Ӈ�KR4a�"O�Xk��]� ��@�T<�!
'"ONm�ӧR[�2ȏ?X?�Q��"O4��'(��0����a�<���"O��j�!ٰK�2E�t��w����t"O�u�lE�H��S*N�Z�""O`+�ջ:��7 6����"Od��@��y M��n�Ml�H0�"O�Q៟E�c�l�,F���r"O��"�(U�v��(� ��Xޜ�pg"OT���(d�h��$%U�E�\�v"O��waT5T�@`��ȯo�F�u"O4鐖E����j��^�M�����"O1��ϗ�bV* � F�Yvؼ:"O���*Z+L�CRO?yZ~�7"OZ-0!$M[��1v.�
a��K�"O�1B(�;KN�R�A67�Ρ��"OBl{�o�[�@X��j�:iR��8�"O��鵭_�J RЃdg�#5I;�"O֜{�!JoF\�7��
F�Ajr"O���BO"$2Qx4&�.��*�"O$ b�ʡ^����*ķYq ��"O���6�H����p#�@\�$R"O̙����av�yQW��I��b&"O��@���~�UHË?м*�"O�%����&��`�Q͂�q*�ѠV"O<��ʡ�D���-�&%���(�"O�i��NSR�
�q�)I���	�"O�Aq��y�2FK�M⦬k�"O���Ɍ�U|�P�H42����"O8�#���w4ثŊ�j�j�	"O���OЏ�Ҭ31$\	!t��	0"O��Y�������d�*NjR�ZQ"O=��
ǭB��չ�X}Mj� �"Oj��s�H�sB �#�8Q��q[�"O��['�% �ac��Y� c�"O��a�HD u��`4��->����@"O�� nƊ`ϼ�����5 ���"O�ؘfD�.c�xA�c�� �`�x�"Of0{W���`�����@ B�4,f"O� ĳM�|z��yT��/,��p�"O6Q��'��p�,J�m	�ea�2"O��{��Z�T�U��|	nmH�"Or�ZBT�[qɡ�:���"OzD�D��p�2�rkA�5����&"O ��w�_'('
p�4�ס?�F0�"OJ!�%�^�=�FQ�E/�l��yId"O:R��C<o���Wn�P�H�ґ"ON���hGw1.y��nչe�ʄY�"O����� l��L�f\6|�1�P"Of����t��U���8Sop�A�"O���� 5u0�q!�,^d�w"O������*=�"�b`�xZdس�"O��p`B�oެ�� �&$E2��U"O�qjC�Ux�#�A>eU~�P&"OxE���./�p��A�\���Jv"Oz1ɱ��	zn���c�'r��"O|��GF�#����M=SN+�"O��aP��Z�駍�5%ٺ�@�"O���,h ������Td	 "O\�S����	!.MZ1#�49�"O M8G�iw2�p�Q2<�Ԅz"O`h��hM�#f,q��V�SO�ؖ"O�\Y�n�|��%J�&��W���"O�K��ǅZH\��dG'OAbY"O*L('B�L��l��	��5Y7"O�L���~�|�0�����6"O�)�dn�w�DȐ�M�;��1"Oh@��f��	RUa�ؖ`0�"O(���l�4"�"��f��5����"O0����Qz �CoM�0�j�"O�̀�%ȓy�h�&�O&����T"O�[�lň!�$;"��]%�m�"O�e4�Z�2�\PC�'��|r���"OƉ��E�[ђ$��R�Cs<��C"O4-Y�L��al.c�/2Mp�%��"Ori�2ETI��IV�I�bz���"O���d@Nh�� A.rH�jV"O0\���8͔� $`)��Kf"O���J�:�z��m�.C(x�G"O�aq�IS�IhB�BGCP/���%"Oe��&�V?fT
���@N��i�"O2�+�C�̈	S��&�Õ"O�m�d�U\t�e�r�	�"OVD�w�'6�I1P��}mF0�"OV��DFz���h��� �� #�y��ѫw�L�������cϥ�yB�N7�܈b�y�U
rˈ��y�Ƈ./��Bp˃ ��Ͱ1R��y"X!.�N���G1��@a�.�y�nH0u    ��   �  /  r    `+  �7  �C  �O  S[  Bd  Ck  �q  �w  #~  n�  ��  ��  6�  z�  �  G�  ��  ��  U�  ��  (�  i�  ��  �  ��  �  ��  6 �	 � N  E) �/ 6 J< �?  Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�� |d��"O
`�(�;���8���-0��1%"Oj4��ND^[��"3/9�0|H�"OB���H��*�ʞRy=a"O�味V�!X��!&F�:J�$���"O,��a
���C�Ą�M�"O,$3%o�-���p���+Ն�:1"O��ݢ1����`���y14]2��i�<�6��{_���c�H�`�fX�$Kn�<��A̼VI�xR[�)�Ć�pඤ�ȓA5��('nߡ4�� �)˩%� ���,��r�؊b#`T�eT09���ȓ!�b��g��}�8�F��-? �ȓ
K|m�ș�VṔ���2�%�ȓ"R�X�j�4JN�1�˘X�i����̹	_�jZ��1!g��zܶ��ȓgil,*�J�
j�Ne��i�J%b���f	�(U��:���G��$Y^م�~r�� S�%T"���k\�jx�ȓ|4�1�îJb��@ӵ�ݩn�V��/[`�"�v4�R�!ʎ<��M�ȓ`:��z�ؚh�J�Z��$HY:	��H��p�m�C1��!��B:��0��EnjZA V;9����J[
2���	��4'J�EA�IVW&��~�(aZ��ӹ�>� o�Y�|�ȓ�f�A�
Ο7�H��M�$�����mޠP����/���ANXo*�ȓTv�����{ ��-7�*h��I��sB�8�8���3����ȓNe*M�悡;������X�o��!�ȓ'lj�#F�m�+R&;�|��2)n�C��0S4���T:
b���:�0!��e֊��)��ͷV��,�ȓ0�&�8#���� ع�L�����;�P�AFd���,w�6d��r�EQ�( �gVlɦ�M,H��,DP���|�I	$G#\���ȓ"�)���E�B	yt&B�^�LɅ�4�� ��eëF�ڙ��n��R�p�ȓp`@}bŇ�=�$�AUN��P����L��p���_�a�)�Y�!��-��u�5���o}�`iF�@A�p ��F�\�0��[���IF/5���k>bTؖ�;K'DT`�^��@��fnV���Y�b�lI��	����ȓ,nٛ��Ć3���kC��8�m�ȓ'� I ���x<=���޳{��	��6��(� N�����
�y2<��ȓx;6q��I�
=  yG�O�,�!�ȓW�>���.؜ɰB��;�����`9"�ˁl�$@��- G��D�ȓ���zF"� ~\�`%�[�ل�E�1�N�;f��P7�.
�T̈́�4 ��QS�[@��o�|h���h�c�A�,@�X*1�֧jN���"�q��� ��Hp%����ȓ]�9+���.E��T�qA:!Θ�ȓ<d���jF�,�*x�d(�9w�Ňȓg�\x�b��/k��<8�ɔ�(��U��Q^��ç�	)��c���d�6�ȓ��-	q �Gp�p�ԭPpGx��S�? ��KG��"����(���sa"OTEq������ �+�+?�2�R�"O��.ܮHְL؃h�2��""Ob�iU�Dt�Z�p��Ը�<Ej"OF�qSƏ��EXQ��'��Y��"O�|c����B�d�c�8X	c"OP��&�\ �za�H�A�P��%"O.��%kְڲ,�+v����"O:  dZ�@β��R=��IrT"O�- �Z\tu�[�輑�"O�×@ RJ���#qRaF"Oz�8�䞐%�L�FnM�blt�i�"O�q�t��|M�j�,�/S&0�"O$�& r�<�J�%kX@x1"O�88Ga��\H&�+�j. ��m�"O�U[�N��`��'��x�t���"Ol�Bp�^*���������Q��"O��E"ěI�d]�@�8n��Zs"O�%�R�U1pС�6�D,�Bzr"O���6�ۖ%�vP0���m���R "O�	�3	�07�Ơ�`"�p����"O�Y����e�@-B�%���q4"O�pZ�=E� �:���?���C"O �g�-d ��IR�Ҁ]�$}��"O�Ѓ�DQT~�Ċ`��"�m��"Oj��&��!U��p�ʽB:Jr"On����&�jE�C' 	v�BE"O�,I�	�(�  H�O^%b^e" "O|h
ĄG�I�&�: ު(�&"O��	DB��g�R%Ң�¹b�̅!e"O8�H��I*Hă�%�it"L�B"O�邵LF�T�"}��ł�e8C�"O���q�˴K;�����\�fz>� "Oy㕋ͻ5�i8��ݮ$`4%#6"Ox�[cG��0��(��&xz�D �"O��;2�"$"�Z�Ub�с"O�t'$ǔk�����O�؉�"O�U��v=z��cB�1�C"O�8����N��ч��؉!"O��6���w�@zU(�?}ʴAS�"O~Ab�ޑYp�yQG٣A�Bbf"O�Ya��=!l���Ɔ�b�V��!"O�!)��Y�fx���eE\z0	J�"O>��pg�0Z�2=�C�A�Hy�"Ob\B��;h�`��Ɇ*���S"O�h�T�ÕZ(jܫ� ��+�Ƚa""O�A���I�{"��qReM.v�\�J"O�I��cR�G�Fm+De����(�"Ov�M�{�Ҵ�U���F�T��"O� ��M�g��l�a��8{�Y*7"O�Z��іh��8`�tm�`�"O&ESS��M�,ɠ��b��b$"O,y0GD�!�<�Y#dYF��c"OV�Wc�6�:�3�	�C��:�"O�`y!�������3-�<�"O��!S��3C����ǇZ��\�C"O�V��vA����EE�@�J�yT"OtXa�Ǫ|�t�2&�ۥF<��BC"O�i�w��&dUj��+,1�4�"O���I�tͰ5���߷O�y9p"O��&�(w�̕Z���
P�C�"O1@ŏΞ
f�}KT��}�P�&"O@%����-Zw*�`C�#���"O01#�m�{�0Rda�#�"O� �	�e���Z� TX�؉B'"Ot�[��*Y�~����4[�h�1P"O��@�K�4Xպs-َbF�ģ"O�-��H�l붼�t,�0F(���!"O�����G>�`R+�0Zy�6"O�eXu럋>���i��wf�%�Q"O����d"�9c*��h>�`;�"O.T���T�`~fM����q)X�h�"O,�YD�#H��k\��t��"O�ɢ%b��/�P5P!m��hb5�%"O���0�φO�Z��k͡1���k�"O�``I�4g$�1шىK�yR�"O6|�D(
46�jf��\��A8�"O�ukg��<Pz�Aa`�#�h��"O@PQ%ƃ^R��p� �p���"O�xjd�j���a�ݾ
L�t�V"O�(Z�[�3p�����CE���r"O.��E�	Sn���
W)^?n��D"O����)�e=!쎷E+���"O����!,\�| �-Z�6xtb�"O ��.X������.��K
�!	�"O���*� �|�S��N ��irU"Ofl0��h=��@�D 5K��� �"O�<kqO�D�
�AۣFj�@2�"O�2���w��"��QL�.a��"ORp�2H��X��a�Ԇ	���A"O�u3o�A�dr�R3�Vy�!"Oؔ�sO]�:��@��z���U"O4�k�a].����E�j	�p"O�1`�	
 ��x1�F�C���XP"O�𪰇O�<�D�8��$m�p��"O����Ȃ0z�L	���K�(��	ˆ"O0���<�*��4bڥ�V<(�"O�m��OE SX�7$�f�31"O�x��R�8�k�]8�U��"O���/�4Q����TdN�lЌ�Qc"Ov���j�3����cč�Dm��"O��ۗ@^�?1�H��ի:�晀0"O8��M�T#Z�h����B0p�r�"OR|q5��*?��ATn�(Ta+�"O��zc��n��w-ݏ���v"O|��u�&�j���?$��q"O~4���7,��)q�V3h���s"OJ�r3M�i�[��V�ZY�u��"Oҍ�dD 0��ER�<hbv�A%"Ohx�  >,jȁ��"){�M{�"O�(�b�Aq�tQR����]���
�')\5fŋQk���M�r���b�'�~-2�+��'4���Ůe9����'��1gOJ)'}.��a��^�F�'W�1�( a��IJ�s�ź�'"D8"�J�,�^P�"�ب@	�'�ʀ�F�9Q�  �����X��'�p�Z�-3�����5{?���'���-c9@yq�U�i���s�'�5��A�g*f�)A��$u���*�'В}�%�G(}b`�e!Эe���Q�'�Xi���2���@�T�^x�a
�'�^dk�D��h�J�Q��B�d�H��	�'o���� ̗Q�l��@R�]� ���'ƶ�3�ʑ�����F`[�J���'��� !L�,Dl�F��6}� ���'�8#R�F!*(@��5CA	z�����'Ϙ�q� ]�h�P�g�fMT���� �ኃ)4�J&ךF�0�x�"O�\��]-|�9���G��0��"OTE�2cQ~B(�b��)��"OD)@p�1�uKЧ{�a� "O؈+q��6#\���<4�d5h��'�B�'���'	�'/�'�B�'�����,�a�Ԍ�fnA�Z��AD�'���'�B�'3R�'��'���'�d �\���Aa2�E�*�D�@e�'O��'��'��'�R�'���'A���Qg;Lۈ�7���@���s�'jb�'�R�' ��'�R�'J��'d�i�a`P|L!�� �
���'y�'��'v��':��'���'w6��0�Q;�蕧S� 耒�'���'��'~��'��'�2�'�R�!$F�2o�H���+'�q5�']"�'r"�'d��'Y��'-��'S@�2�B�;�.��fZ>"V d3��'4��'s2�'��'���'\2�':���B)0��ہ�C��J���'���'���'W��'���'���'��a���.u�6h�4h�.d�,�C��'��'���'\b�'�R�'��'�y�QF�	�pP���4 �HQ1�'ZB�'Cr�'��'?��'���'Tv��"�
>"Y�us����:���'�B�'@��'-��'O��'��'��x*4`�2U�f{%k؅�H C��'|B�'�R�'H��'�@x� ���O|-ۅhϯ#���F$߄zh�a��L�ry��'�)�3?i7�iVf��t"��6j���V���b��x�tf�	����O&��,�� ?��42ˆ���,I7~P�\E&^�+�d#��iD���}����O�4ˤ-%�N�N?ɖ�	�\I܁�!�#lk,�Ҵ�8�����'Y�>j��-��z�I��5�U��)ة�M#R��w���K~2�Ӽ��f¨��o��P��uRD�(92�i��<%?	���7+(�ɟ�v;����i�BJѐz��牶�2��0��)�	E{�O~���)w2�p���k�Bw-S6�ybW�d$�@�ٴm־Q�<y�cʻW Еȁ�Q2���jf�.�?qM>��OB�$��	E}�DP"zx���W�HZ��Dʢ���~�
E�pl\�1��]� ��E����@/3�����%��j�x�m 0q����D�O?�I�:!�4�REGp���BN,U�v牪�M� �U~��'��|�O��	���F�~<˲��!I�� p�'7°inr�ǝ	��	��O��R)[$U���48���̑$A�A�a獥Q^�O���|2��?���?��b�&ijE눷������N��99/Or�n�
uښ|��������?��O���,1Pu 4A,����aJc�ɔ�Mk'�i��)��z���7xM��r7Nԫu6�T�d#G, ���//@KT�	%B(��m��T�p�[2�>�!�<���Ǧz��Q�A3���8���)�?Y���?����?�'����B�L�֟T�Rh������H�D��DFCşd�	L������a�4�?a���!7�Q�9'��Ai�8�@9�P��<���_��"�kK�#3`Q����I���k��i��@ ć�n�l�YE����D�O���O���O*��2���y`�MSQ�K+~����E,�.������	��M#�B�|���?K>�A	��[2 J4%�6O�y�C�!��P�x)ٴ���Oz� �5-J��y2���C(I��ά��piggr[?|��ԁ��4��<���v�'f\˓�?	���?���F�`�u��=E������?)9�t��?.O�Dl�f��������V��N
� �Ul�0t�`p�Ge=��Ģ<�p�i��6m�ܟ0'>m�S
�����զ<}ɶ'$<���� �Z-a�"0�r"Iy��O���lO�TD�'���)��*y�B����ţ$%��"��'!"�'��O/剾�M��F��d��I�"�1u+���A�]m,�X���?�����'�剎�Mu��)�1:����3�J�P����ߛ&�'9�q��X	�y"�'o���G�c�-�!T� ���K��i����(�P(�f�ĕ'���'��'�2�'���ID�yp0�ˮq�Ry���N2X��4�h����?1����'�?��Ӽ;C#�d���
	�@b0��p�c���r�H��X}�O)��'ۀA(f�$�y�HE�C6��R�m��D����FX��y"��s>H�F��l-�'q�	˟d���ml=�f�7,IdM��`�s����矀����8�'��7�� ���O��d�XF�	���	D� ���,3X�@㟈�'��7��¦!̓��Ą?u'����n�S�؝ᴫ��<�d�ODX��h�2�.���ʥ<1��Jw���D+���?����CAd̸t�Z�&�d��Aaߦ�?i���?9���?��I�O�ѹe�ھ hX���S}t�z���O�Mo3k��}�Iß��I|�Ӽ3A�[ 0Q&I�&�et�uI����<�i��6��ݦ�+&AN#�R�����3A�� C(@'!�B��B�)_��qAq'V�p���'�x�'���'��'�"�'<�i�$�y_�ts��O;M�0��P����4y}���?a���䧆?�R�j�J-@3�3O�y��ݐ��YΦ�H�4�yB���O����!"�~����['1<��d�]��(�)�	��+����^u�4$�ȗ'}��Y0Ϥ2$Fu�lR(u�h`��'B�'�B��TR����4NW�����rK�A!E�R�m��峳�\!_DX ���?���Z�X"�4/+���'U��E��"�3�	��-(�(�];g�T�(�'�B�"�|��-�F�œ���O(�8w�x�� Ҥ`'O�ՖT���Ȳa<|�i�7O��$�O����O��d�O��?uCq�L� �x���&6�!#c������˟�"�4Nd��'�?�����v�$�{��I:3:���e�%i ���'�	��M��i�Bn�ppԓ�'2�0Z�l�w�p�˶%_*X��; ��;t��h���7F_��őx��<���?I��?���;�^�釧�Z6�c0����?����D�ʦ�q�ȏ͟H�	�8�O(���%+��DS�@�uė�nCV0��O ˓q���j�T��_���?�(`e˛��&N`L)# ��x)�c��Œ09�k�<	vb�޺�BiG:HFT�љx�e��M��M���"����c���x�d�OH���O6��I�<)g�ipN��'j�lI95��S�\���N#��'X��'(�'��	�M�g�n֐��"����A����Ki���a��:���"d���O�5HFdόn�L��D'�<	�oT2G�B���fp�Ȱ�b�_�<y,O��$�O����O6�d�O,ʧ4c� �È
}����AL<A�Px��i�r,C��'���'k��4�(�Af��+Y)�b�Ҽ22���^Ԧ��ܴN�_����?�S�K���Wj�4��ϛ 1P�w��5-*�2@{�� 0	A;s;~i�#�I�	{yR�'H�?��ț�H��)�H�F��s��?1��?q/O�=m�9O�l�����	�
��U��M�cI�Tjp!9H�1�?9.O�lڍ�M+��'q���6)SF"mk"qr!�U�7���I�0cD�Ӗ,Vf��|Hr+�J?���u�4~�&�i�M�OP�[2�_9�g(X�l�j1��.�Od�D�O���OȢ}Z��\ �%�'^z�)�A�����M�v�,4&B�'���'�ɧy����U ��` � )�Xԙ�E��yJj�T�n���M[��54%��C�
H����4xM��0��*{�6��a\�0TոbAJ�JE�L>�*O.�d�O��$�OX�d�O"�k�LGQ��Jd�Z�u �sr��<a�i�<� �'(b�'��O)ү�uU��aU8���(@�J�L.�	��o�<�O|����?9���H
`I�'*�q���k7+Ȓ,IVoz���{�fM�B�K�O���s�>�bž<�f��8D�3wE]�`ش�8�/�?����?���?ͧ����ACgW���M�	G�:�It�B�*>D�agП��I^����$�ߦE��4�?)�@�37�"%EZ?K>;�z�;0�̃IR�	����S��.��q"kyR�Og��P)����&�F��m8�M&p1���ٟ0��ȟ�	����K�'Z����$�B)���b�������?���HX��a�)����'�r�|�_�K��(*�=�2�	�!�4E�$�>I�i�n6m�OD��d�0{���Ot�{�h�5J B`��E��uhAc��7z��U��\�O���?A���?A�&@ ��b�=;�8�i�&.����?�)O�lڒD
��	̟��IR���Z=�� ��|O���Tb�#��$�<)��iX�7�d��%>���
`p�JG��
7��Y��уe�p� ����/&DASH�_yb�O�(���:qv�'v��` Gy$�ł�5K�5���'H��'2���O7�	�MsVm�u�z@�C�^'9��H�L����K��?i���'~剗�M3�-z�X�����)��x酏�-0��'�X=2���yb�'����c%��RW,��R[�(���J�	�x�[��	�`]d�Q�b�,�'��'�B�'�"�'@�S�zL}p�M�Rvz��@�?|4-�޴O�������?9����'�?��ӼS�-Z?hZ�l��)ֈJ�v��d�K5��n��In}�O����'���:t�ʗ�y��18oJ�x�-�R����`�*�M{gI	괲o=w3�'$$ܕ'�'1���g_*_Ӑ�rh�%3���1�'��'�2Q� �޴(Ț-���?��o�0�{���F��8ꡪ��o 6����P���۴V؛V2O
�A���0&@��"|Uh"�ܼt?���x�Ipa�4�|0��T�~Zw
,آP���l�z(K0�'�Y���D�$CE.Z�]R�"��'iR�'��'>�>睉q��L�%IsBI��HH�}����I��M"�)�?���?�����Ӽ���ܘFD*�yuOK�
��(����<i#�i�7��O�$�G*s����OR���B�����B4fY�ŢIZ�J͚=�H�ab����OL˓�?���?���?��m���rL��q�$�.�l0!T� ~yR�q�^��4��O����O��ɾ|��;�p���ϛTH��I�GxT�+-Ob�l���M��'�O�4�'�0l�W��1H�F��奁�����F�!���1^�ˣ��=��8r�z�IPy��D��L:`�g4�`c(_r�'32�'�O��I��M� �؏�?�RȎ� �E���S�<%X�T��"�?�����'M�I6�M�!�i@R$X�H���'�Fٺ=�n%B0����Կ�y�ۀ��8ʤ�Z�9�@E�"7O�D�� ^c����љBbD��U+� B�'���'&��'H��'B�pl0�@�?'B�B�&ѹ|�0���e�OB�$�OX=oZ���ȟ����`�'*�U�ß�^��8���!X�����O��Gٛ�$l����Sh�>%��6O���A�Cb�eM�J�~%�B�8.a��Ov�	qv�;�ĳ<���?���?aB�ޘ���i��� z]|���9�?�����W�����'����	��t�O�pI#�B�3�jr��T"�V��O����p�<\��m�S�?�A�Өz��"���p3E�Tp%&e�\z2͔';�t�%t:��4�|L�@�F��� � z�I{pe��"�''��'��$R��S�4 ���%�M�Ji��j��-|�����?���?шr]�`��4)��%��K=H���� c�T�u�i�7-E5[���C9O���²e�]9#V1i8@�S�? �
�n�%�$�Sj��L&�}�D2O��?y���?i���?i����
c��9���t����+X%��Plگ5
f�����$�IT�'�?�;Q\Z��ԌR2zd�7��)F2E�iy�7��ٟ@ק�D�O���f��[�
dʙ'in� 6j �K��� �θ3���؞'�8:P�X�^|��:�|B^���ҟT����$[a&*�$K�Y�Ɯ�s��؟������	Uyr�sӜ�0�%�O��d�O&�� c�(Hl9�킹9V���l#��Gy2pӬ�mz��IM}��]�CTte��c�46VtTW`�y�AW�]Z��a���8?j9��O�oݵ��훷9�(�J�o.�Y���Nu��:��7�������?���?I���h���$.O��K&��%�&%	�_������5�"*� ����?�;\�ֵc��&n���3��5=
��Vk�v�p��HmZZ��<뵮h���I)V����M�ڽ�&�V �-��K#&4�h�B*�C�Icy��'2�'�"�'H�BS�.���S�M�p�AAȁ4^q�ɨ�M�୛��?���?�'���O��94+��yBV�z,J�1��P�� �<Y��i1`6��ş�%>��S�?�A��~͔�3��wX�e�ׂD� �`�vI�Ry�K�#o.p�G�_3q+�'n�	+��)� � (�x%�&J������՟`�	�8�i>5�'��7���^�$ǂ�Ac.����b&+���v���O��x�'���i+6-܌Ki���.s�p��c���y���HH�$�O�=@��	�U��Y�<���q0k��M߸$!³ky�%R��֫d��OL���O�d�O���&��2|���E/�"P����g���B�F��ɟ�I��M3P��|:���?�H>�m�(x���艘��Ȑ���y�P��nZ��M[��Ic����<���S�r����d��cr/N
�舦,o�׺�䓭��OH��O���'&�I�a�qp���g�R/29l�D�O�˓X��f�����'fbY>��V�=��0�׹k�|�1"?�)O~Ql���MC�'�O��U������<�
�B������b���%Ɋ�3�my��Ož��`O�V��'�Խr"MN�:�1������N����'���'t����OT�$�M0#ʣT0�i��M0S5���׉\2jV�O����O&㟰�'Y<6-�_���#'_�;o�p�Q�H4 �mZޟ(2��O5��I����� [t�����Sy�N.L�hT9qoE�2��S��y�^���	ן`����|�I��4�O>U�w�ȷSQ2q�w ��]Fx�B�!uӾ�%j�O
�D�Op�����O�n=+��1�0��]��6��
c��mo��M+�'��i>A�͟0S3H���0�If�%aK
�.��f F�X�I���� @�nhb %��'A��'D�`I��%M`���!
Y���	��'���'��X�@�4.������?!�R݆�a��-u� Z@�� ��a9�_�0�4eΛ61O��E)�AY���Q�|�!�SNH�ϓ�?9��ԙB�jT1���d��P<� @�AD��ԗ<�nd($b9sh�7٢*,v���OX���O���1ڧ�?qjCP�,43���[���� ��6�yQ �K�L�����?�;]��p�f��b}`��IW�h�GEr�i(��K�Bs�'��
,�a����+�h���[�Ot!��*F<d���|�Z�`�	�t�I㟼�	[�䚯Yz����6 )^�C#gpy�a�� h�B�O��D�O��I�|��s�|T��F*̨��	�R2p\�)O��lZ�M�'ʉO��$�'b5aG�4G�8��!KcjU�X�y���2Q���țj]LQ"�DF�	\y��&(U��X2Ì�/h�Ѻ���K_��'r�'�OK�I��M�c��$�?qNC+�l���쁹�@��5���?I����'Z�I�M�ֵi�Rm\9=���*bO�m����ū�{�ҽY�����yb�'��Y��^���Q+�T����5�5����<����i *g���ϛ�y��'�b�'���'���	J=�]�$',1Aʸ���#���O:�d�ᦽs�E|>���%�la�b�B�6��'�D�^!� �"���<!�Oln���M��Z��J3O��<A��?�n����YYQT	
��!o.��C�ׅ8��a�U�� ����$�O����O��DP3>#���&MO�}ԭ�s���J���O�ʓ=ʛ֯Y����'��U>��S�A�G�U�2��K0|]qՏ<?1�O�djӪ��IV��?��iY &w"б�"�.%�F�"��ۄ3����>8p�l�'4�TE���H��|"�Ѥ�yR�[ X�N9�W�V(l2�'���'c���Z��!ݴ,�1���Hw�U.AK�%ۅMC� �̔�����	r���$�ʦ���OĽK�d���l^O�8pG�B)�ME�i���B�Ǔ�y��'�(���(�)I4T��V���E��!��(�w��~��Єd|��'���'O��'�R�' 哚R0�Y�0��'
ZrU�ģ� 0�1i�4�x����?1����'�?��Ӽ�+�N�P�83���WV����9.��֣r��@�IU}�O��T�O��"@�y����vn�-Z���BBc��-�y��^�U���*1��'f��'�������ɤ2�,5I�N��}\Lz�J��@��	؟l��� �'FB6mþhz˓�?q'*Z�r��H1! �>\�8D@ ߓ��'��I�M3�i����>qv�؅2��m��B̶]�r$5��<i��:*��+g�,���x-O��i��HH�����O̰Ӷ�Ń:R-i�s���[t��O�$�O0�d�O��}�]?���O�L�ꨩ��� C��t���:Л�>4�B�'i�4��ei1'ՊU�\��ܲix�m�g9ORdl���M[��iDdI�fK��y��'א���0��ܙ� �x
R��,S�$B�����g!�d�<I���?����?I���?I�V)Y)�� �\^��z�C ��d[ʦ��B�cy��'���[>��	�\@���0J^.C�4�3b��%Nm�|�'�J7�[٦����'�z����!� �Mx� �r)>r��A�H�*H�/O��c�A>j�8Iz"m3�d�<A�DP������7E2������?1���?9��?�'��$ͦ!X�ҟ���c�.u5����-A�a�GL
ȟ��I}����ߦa��4��v
ɪ\ch�� ir{F��=�U;��F��y��'�jQ��ʥo ��0S������5f��!4�ŨĔWz}��I��y��'"�'���'���I� Q�x���@�QI��t�\�S��O��$T��#�"c>��I䟤&�h�/�%#]�80�j+b�������?	�O��o��M��''`6)!D���<)��>�ă2��%��M5��~p@��o�~��9bnׄ�����Oz���O~���6k=Ȕ��ӊS�4� �.�������OX˓��FG�,&��'�P>m�Ѣ٥0\̐&R�7@�� �4?/Ov�n��M{�'7�O��4�Ŕ*��+V��mWp�Xv���J'^$A2�mZ�I��U����\y!�k�U�ɾ��)u�V!r���Ѐ$ڌOF���ן�I֟p�)�S\y�me�*�B�m_&5SD�r�.�x�V\@D��-&���d�Ol�D%�Iyy�nsӖE���ނ���&�
�� �C������I�n��`��al�,�I�1<����Xq�!�'�R�����.0h
�8���7Y���Py"�'��'�'rb]>q��%V�f��$C�>��U'ć�M�
�-�?)���?Ɉ�d�y׏��cb\Ic�oF,����3}�6M�榉���4���)�O�#P��g�󤟓MI>��@�J� �
�·튕]��dG(��%i(�(Kۼ�O�˓�?��� �kF�Np����Ͳ DC���?a��?)OR1n9\�P��ɟ�Iv�Xp6n�-Xs��-�JwJ<��E��syr�~�n n��<��O����I�Qд�1� �1t�;W5O���G.�`������<��'p����%�\��?A�R�LtD�#��57p������?���?�����tY�C�<�X\ MTSd0Q��F՟���4 ������?q���?�I>ͻ.�> �"�9w�uB@�Q�;�����M˶�i[�7M%��	� 2O����5��I:r&
�"�  ��b_������r�:�,���<	���?1��?y���?)f@��C��lse��%G1y�bؐ�����9���������㟘&?��I#H4�=��LP�U�V=��W�S�&y�'��i�H��2����陇C�����յ�x��aj��ZcpR�0���n�.��><t�{M>	-O୫��7 �Y�h!>_�0�t��O��D�O����O�I�<�ƺi�u(3�'��,S�݄綉��`H?.k���'�2�'
�'7削�M[R�i��6P0wl��0��Gw��b��$d�B%�ľ����O�iZG�7�tu+2Ʈ<���@�kl� K�6y��֜t?(uckH-P?�D�O��O����OJ�$?��"(aNYc�I�	�T,��#Gj$������	��M�B��|���?iK>�ԫNs�j�����H���aC��D��[�@Y�4`�v�O �S`
U��y��'�z]�"��3r�\�K�/� �~�3$c�q���#"M�d��'������ޟ0�I0+�<��1�C�^@�4R�kJM� �	۟Ė'Vx7��ʓ�?�+����w��):��9b܌d[
��5����'���i5n��.����QJ��͈FH�x�fAV+�в���E����A�6��BJ��u���K>����y�!�'��ic"EwC���O����O���i�<���ilL�sT�C8����M/3�1Z�>���'����<�E�iU��s���)�	<en1!�mӴPmچsR���uz�T�	*�L�� � N}��']\����-��A�d`W'r8�'�����D�Iݟ|�	��(�	M��N�0X6j��R�ssd(0����7��p�����O��$<���O`�4�xp��	ʘ0 -Y;��Q��ʦR�4�y�Q���?��I�,��i8��g�D�N�f�@`[7 ��>�-1F�r��kV���/�)� ��P��]y2�'JI�}��AȄGC���ޛU�R�'A��'��<�M���?1��?A׏��@�
�H�Dd�t(5m���㟀�'�7-�٦����Ė�DBDq'��~(p4�!�Hx�D�Oh����Ύ>����<��'l'����� ��?�)��;t�����!�1XR����?y���?���?���I�O8tȥa�8�)p�oK�P�u"R��O� o���a�I��<�IU�Ӽ�r�  =�֥k�C�#K:�x��W�<Ѧ�i��6ҦٓևQ�bP�I��A�+(+�*h�Ёg7
e3�V<Q�h�;��	�h�%�ȗ'fR�'���'��'s�L@R�2(R=1��U�_�HER�8ܴ`���Z/O�$���O�q���F�^�h7g�
]T���<y��i�6M�џ�%>����?��T"��_�r�rp�ډO7�83� �vq�L�"�'�L�!^=�zy�T�|�Q�0#��N�2�9kU�JJ,0�so�d���(�	֟�SBywӐ�d��O^Պ��<Q�Ā�Սm�ꝸ��O ��.��py��`�jQl�ퟌx��9i��"�iC90�a��I:?*6���~�l�	/|j�0�լ��;���'��Bu��㡢	xϔ�˷� �r2�Y{��e���	�$�����	ٟ���@�<`rJ�+�=rf����X�?���?���i�����O�b�'<�' `hq��6s����@��y�,��0O\�$�&�l�r���w�zdQ�4Of�$ 0� MRaF8I�@HOǥ@ζ<��/�!3\��*�d�<����?i��?�!�_'W���V@�9/���r���?y���]���	S{y"�'��Sq?0��rϏ�C���BMWz~���$��U�޴�yb��T�O������ �`hK[*-^�����t�����֛r���?��I	Y��&�8�@DD�W�Uc2�Z|d��{�E�ß��	埴�I�b>ٔ'hh6�S^ѐɻ��O2/�R���-�.x�|��FM�O����O�⟔�'6M�1*&�4慒�x�*X6
�q3.�oH���Y"
���i�mȎg��E��jry/ �G_�Iz�f#C��x�HՑ�y�U�p����۟���˟P�O#�0�iD?l�r�낥��>(#P�t����m�<����䧬?Y�Ӽ��KV�C�ĉ�N_L�����M?}��v e���IS}�O��$�'�>`�A����yF�:'��Y��\1�`����P�y2`;��R�Fd�'��Iٟ��� �FE�2�G�k�`Q�(A�b�bP���8��ڟt�'��6͎54F��d�O����1J*PSn�C���@�c4��ė'Ur7m�ʦϓ����5�� ��M-jF<�2H<��$�O�Բq'ÔS�ݳc��<��'ZG"�6���?�0�\�V"����J�5I%R�'��'����ğ��e�AMr
�an+�",JA �Ο��ݴ0��?)�����y�,Dx��I�V�ۡ�rP��!R��~R�i3�7��O�lB�ʈX��O.�p���2n���o
Z�;rH9���.,=54�O�˓�?���?Q���?Y�j1���흺��6	�<�Q,On�lZI����I�x�	D��0��l)(�d�c�2M�!���Wy�Av��l�<�J|b���?�&Ռ�$�c=�nȒb��64Cb�HġA��Ď!Ɗ]鄧�1!>�O��� 9���܁:\��� B#=6<�����?��?i��|�+O��lZ=����	:�"���I3Q�������v�d�	ϟ0�?y/O�m���M�<��_�/�^�ȡ�M�S�RX��:!O����?!FlƂO)J�;��R�����d��1_�d:g.�+�&�HV�+�2(��?A���?A��?����O#�R7�ĢQc��P�m��!`���'���'��6דR��	�O`��?���;g!>P���׷�t��
U�X�IU}R�~�8	l����H��͇n��	�@rG�4Z�h�1�iN1���G�	\�e+\���%���'u�'D��'3��9�˃�%i��s��+����'�"R�4��4U����?�����7��$a	@� ���C�B�	fy" t�(�o�<�I|J����i�!X7d�PE��l]WV<p򮊙��az��X���D�$AB��h�����-
qa��'2�Q*b���� EB#�^��� �8��;����/�\BZ&�!�(%���'�X��F���8�6L��:�TTQO8��=����1y���2�Ʌ>i�T�1qesI"�)èp��Չ��܎)z��Xs�)X�Z<j6-]�r>�xb���Z���� �r���!��FSvH��d·�Dh�Ԧ�K�x��r��uz�͊bƃ�SYr�ո��3f�f��j"G�,M5�I��/�l�A�!W5�0���z�D9.>�����ĵx��1�dD�ē�?i�����?a�[Ӡl`F��� ܮd;q8T6�[���?i���?����?����U�R���2I`�AA�F;A�&(�
VnPo�@�����%�D����������l7-� �@lBu.�%0Z���Û&�'���'"�'��&Cb�����DF��f�h4���;�d�6�	'�M������?���aFDL��NS�	�J�FI�f`�!4`±�Q����'?�'	B�ԇB��SIy�O�F��$�,A�@�u���� �w"8���Ol�d�Y��c��T?Q�ȑ�^j!�o�>O�(- ��t��$�OFM��H�O�i���'��]��X u�i�!�	)j��d��@@J7��O"�U�#�r�������:~���s�k[A*�A! �C���J�9sL��'��'���U��O�d��p㇑VL�Fb_�lq�u9�E{�2к U"+1O>5�ɝ���&�?�A"'.�W��x޴�?����?�tL���|����~(�
(Yz�f�3}z��$B�>~|c���ցA����Iϟ��� ӝJ���r1�]�r�D3�l]�M���A1���a�x�O���|Zw���B��l*�9؆�W�])�|��O��[q���O:�d�O �d�Zu(E`#-l���&}��=�A�Q�&�'���'N�'��	�S��`��ʱr �j���Q��l�f�5�	�T��ޟ�'�x��3z>U�F
��D��T�XtTTT��>!���?�J>)/O��R���F�N�>�֡ꡨ[�
�(tY�)�>9���?������D-�x'>���(Q3r�@�ɶoG�h���V��Mk���䓈�ǃzs���� 	�(���S�k 8J��iG��'��IP�r��L|r�����.r�h�dS2F�r5�b/�>nr�(&���'�!����?�����o�(�9�,Q�&�Y�:ᛶX�T�u�Ћ�M^?��I�?�O��ʐ�6�D����f�A�׽i�=>5�S�ě�ܴn�@�k���t�R���L8q�loZq�R�ش�?q���?��'��Yy�����Y��f�#"T4�2D��aA�6mE�f��D*�;�ޟXr�@KV��9G�ϝp�Y0�Hߥ�M3���?��1��{V���'��O��rK�?L�Ǿ�"�%ۻFf���'%�I�/�Z�)"��?���,����	��|����jD�p4
Y8��iA�h�S�\����Of��?�q�? l)�W�ݹ;/b�C��M'� �2T����i{�d��՟0��ߟ��	fynH,l�I����U^`��0�D��>�*O���<����?q�g�^�k�f�: '�):��)���	R�<9(O`���O��Ġ<�p#���IΖ\�>髢n�&�����_�[����dy�'T��'(�e#���Q�WI�Ld{�O�UhR��C]����͟���\ybHW�d��맽?Q�"w$-�S�_
���:��?�������O��D�Ox�Б3O ����pk�G��}zW��Pk`Iêw����OH�M����[?���ڟ��S�Y��8f�J3z�l�	�������k�O��d�O��d��wZ�$�|����h˸VF&�蠡�1=� �l��M/O�a�qA������������?i �O���
�>�b�� )�*H �.�j�v�'��ڇ�yB�|�	�&���@� �,�[��}T����)�6M�O�d�O���@}�P�PP�g��8ڸ���E(��
�=�M�!�<�����%�S�P��((O4��y��b�hѩ�Mk 7-�O����O�=�h�`}RW�@�	`?�1&v�\�"���q��mKoZަ��	Ky�M� �yʟ�$�O���f��$��D��o�^ԣ�g��q�&7��OtP+�l	K}Z�l�	Vy��5ƃ�FqR��#���´����)����ޟ��I����	���'��:1oG�c�y��/$ #��A�k�p����O0��?���?�V̛�	���e��cchKb&?%�6��'�2�'2�'��I&�؉O����I�E�Fpp�j_�$ڄ�ܴ���Ol��?A��?�@D��<�篓�Q����T�EfA8%�Щ�P���'���';Z�Z!"	��	�O@����J�'��E��B�������zy��''r�'��y�'��:fB��&�M11p:���K�x,nZ���	Gy��;I��'�?��������u�F���Αj;���R�&w���T�	֟Щ��a�Ė�y��O�M�#�Ul��1�F�N��es�ml���O.yx�B���Ib���O��Ӻ�6Ȥ���:���dB�YV���'Zr��<�yR˪~���Ouz5����,��F��z�|�*ڴ=���ق�i���'�r�O�V����4$�2�"�^%E�j����B�`w�hl�?J��	�\�'���ą1p�ta�$E�2�P�k���PQ�i�"�'�2*�,���D�O��	�66R2�d3j����.�T7-�O��{��	�S��'���'7RA2��N1l#z<�4-ڜJ�XtP��r����@�VH�'S�͟��'RZc=v�
�%R
3�L P�D	Z�Rp*�O���5ON���O���O��Ĥ<Y��4}�~$0�Q+�ZHs��]�� \��'TQ�����T�ɝGV�ݪ���l�vC��ʊp����F~�|�'��'��Q���׋�!����IM��p %��	Z>�0W����MK)O���<A���?9��`���Γ�P��"��4��I腏A�6��B�iZ�'��'i�I�h�Tٯ���d��Xŀxh�&8B�"�$D>
+օmZȟ0�' ��' ��y2�'���L�IMt8ye��j��ڤ΄�+P�&�'�R]��q�������O4���51RBŁ|����bX�\�l#�N�d}�'�2�'� ��'R\����]��H$��C��kv�޽9v�n�vy�e��s-�7��O����O\���}}Zw���2��"n�T�f�Y�xd�I�4�?y�Q�@]Γ��˸O�2Sc��>QN$����5"dȜ��4ut��1�i���'&��O�`�����NܙS�Q%K���eEVk8(n�}��Iџ@�'$���'�2�'%�掭(ت&g%SZ��3GD��
7m�O��D�O�дa�a}"W���	@?�5@�H���{eÆ�������[}�]���1f%?ͧ�?	��?	Рm�HE�e�ǦP��d�c�f
���'�X���>!.OF�D�<)��c$�8�d-����s��pF�֦��0-L�{���I��<�I�?�����`�'P���A�K1\���X%�3R�0���&F�L������O�ʓ�?����?q�ÈZ�M��oS�J����!��2JT��'�2�'���'?� ��O'J�1���	[r��rj
#����4��d�O>˓�?���?aW��<�cB�^2�{��09�< 򦇄n���'��)�'�'BP�P)"�ħ_���v�ѿU�F�J�@aHJ�i���|��'��ȋ��y�>	�NW�%�#C,�e�4��Aզ��I �	ҟ�{���MK����I�T�蒢È*��D/A�1���O�	؟�	�z#p�I�	K§�݊�(� ��E�a�`2�Ǧ��'�n��ms�}�O���O)0�(����q�1@~��#í��Al�֟$�	7=�`�I|�Oܧ�N][�_O�䒒lC�]RRl��f``�۴�?����?��oa�'(2�ڑ3V	�2�M	a�p��L�Y�7��_�1�d �Ɵ Y�-Z�]��=�G!�H;� "!�۝�M3��?Y�>8{Ĝx��'e��OF�Jb!	��z\�`F�K�t�����\(&�K~����?��$"T�ǎ��s�T���J�/&8�q�i�2*� �b��IDy��5B����)ѫĥu%\ŀ�IP���D9/a,�d�<���?i����JL8�� �R�+/p��g&U$:(���b�K�	럘��n�I럜�I�	�yň@�!�"t{�R<���z�x�'��'3�Y�$��o����@^XG$x!�ĘA�2\ C���d�On�� �D�Ol�ؑ6l�l�? �� �ǀ�p�m	2Fy^��3U���	֟��I_y���%���
��	��>WJ|�"��fi��WѦe�	M�IП`�	�W���=��R�pp�2)R�&�ɈeÙѦ���ڟ@�'T�%X��6�)�OP��P-��K7��=L��0iI��j�ND%����������$$���S4��퐜f�fI)5B�V�d�k�^���Or�C@����K�T�O�V�;*L|{�,�����I��WZ��o�ɟ$�	S>���V�I�?���Y��]z�m�
�O-�(��i}\�@�'o�J���OH�$��
��>���5Qt��+9��U�uǞ� ��v���y|2�' ���'��C?PqR� �GѸu�$$��y�I�6R��5h��2J���X.��p?Q�C�&g�Dř��~��]�!R�\�����ER�3Q���ގZ-J(,Z�3kLeYR�b�ĽH#W�HՊUXp@Y�A�5�uL="���th�iD�8T�FR���⠙Q�>x��S�Y! �@�O!���j �}=5�� �<�P��OS<-�‬�/q���*x�6m�O����Oȸ����O��w>ɚ&�A Z정�v-�{�j	X䞲t�8�e�z@���me֑��I�z$�����[����Dj�**��P�5LG��)�˓3z�����&ܗ2��jWC$S�j�	럴ڂ% �w_f��!�F�	��Rf�'�џسdnQ�T��0�!��nYX�G2O�=a��A	&�gl�m-���<�հi�2\�� ��ǯ��i�O�˧w�8��k�<�<�[g�J׌HPo��?A���?)t(�	5�:�Y�m����p*���C${8�$��e�A�G.ȋ�HO� �A�&��R�J�)M�����BɃr���4u��Ks-�j`��j�`I���zt�����	6|���O�?���	��C�%O:���C�c�0��	��*(IU����j�.�
�t����d�	� �̀��ұb�pu����?<�	l=�-+�O��$�|�*U��?��?�&��0�Ȉ�O(Hͪu8��M�g"��ʳK� h���7�V�TM*�~c>�DO%)�YYҫ��*I!P*T(E��t)�eR��4�� ��2���)�����6o��0�bʑ]+`��B|���ߟp��'��_��(�r��d�h��E#B�vI$e�ȓP�0�pr���"S[diFx��4�S�4��Js�9d��,״yc5@���'�R�92�Q�Pr�'R�'���'�?�5oǷ�I�&tl���o��֤Z�0@"`�c1R�PۛO,r@��'O�}��M;��%���Ȉ	����"����KSH��|I�@����0���Cs�&���y@C�Y�V�Ҳ�W�6ܜ�+�E�56K)-�"�y�.�o�?��?)-O*�	��׃d��M��.�?6�<���'�ў�	ň��
�v� 0K�@��� FdK!�M3�i$�'R�V�i���p-
�4�B��rlؗT���A� 4D�@���:b�i���zcVĘf�3D�l�C��Rx1a�5	� ���N2D��R�oԴa%Z-��N[*|_��C�C2D��Hm\�C'^-���K�~�x��&0D���@i�SԫJ��љ�G.D����n�3�x� ���/z��+F�-D��Abn�"B1�%���#��ȫv)D�ض�����!�$˧5$���2a&D�,�ǌ\7	�> ��%H�x�X�*(D��ċ�ec��/��EՒ0 �+D�Гƌ҈$0zm{�"РXhX�F�)D�$r�&�4�X��N��qֈ@�F�#D���OQ�s���j���:PEz&6D��#��9Z�\ q��W��� �	4D����@�HT�Ix��j��|�%->D��5-ΘAu��2�������#�:D���Cω-�r�"1$׳S�Za	F�8D����,�%K]PH� �6[0��8Q�7D�\ G�9jR��N&|9 ��)D���α���XB��(p��pó	(D�TB]�K(�!P ",��Y�  D��y��Ç"�x��Í�/� �U�"D�����s@��.׋!6�c�O"D�,p @yn�X�GU1��P�e D�����E7R���e]�SZ��i��0D�<z�A��!��:�):�E:D��Z���(;���@ꓚ}d��P�-D�D�7/�3�0�"Ӭ%���A�7D�� F�
� �L�4!�F�W�Kx�M%"Oڡ�u�?�DqZv��C��Ї"O�	��U�}�H��%J�O' D�0"O�����a�*\����>'�8V"O�)��
[�C#�)����o!�%�f"O�H���Y�`Ȥ�0O@-z�m3%"OXM;�,��Q�r�x��8.�ҽh "O
-ss��:mI��^
i�>�"O�q�j	���)��j�GH�:"O��G�A��4���#���	r"O�QV�,a,f0�c�����"O��U���l���"	d��"O�xs�g����ȅO]��lC�"O*KwH&1��1�UoS�KںL��"Od\�q��d�3,�n�T2�"O�eJeD�9}8��{0�լ3@�� ቑ�PG���޷���$�ӍN� ��p�B��y�)��TkfY��Y>AB�9S�@���h	5��s� � ��?*�H�%+��1R����'D��r�D�(3���@�0>X�A�d��r�@�Zx��Z��?9� U��@\�l>,|aq�"�ObE���<��U�)�j�9���# �4�A C�<�d�*[�� �b���!��'�J�'\���6
�mI4�C�_�N�z ���tC�Izx2
�o (���8R�2B�ɧ7�X�
�#�B�Ic�� r��C�	r�X���S�oa�  ��(a�B��>���P�nU-����Eٞ+�tB����+b'�lޘ�9e���m�fB�Il��I�6@�?��� jU�.�BB䉟[�8s�j�/�XISf�хK�rC�ɨ� ��!֙b�X��!OP�\C�ɖ �}���,\���� Z�PC�I�-�ؙj���5-Z���c�]�RB�	,R��
#f<@�$��%B�5ohʓQ��J����J<Z��u똼F�N�s�aQ�!�dØ%NRe3���2�@q��բ>J�'�`2�-<O0���'M�Y`���B�=+�f�5�'���c+4;D��@O $p�0�B�&��A��'k,H���E���TX�΂�&�H�b��D
�;�
����j�'K�D|�͒�G���A� �8tSa�ȓJ�����]�A���h�?�$��'o2-9r�>$�O�>U����g��Hs�*R�Z�n��g<D�òo����B���\{�$ ��L;�I�>�쪕�"��g�R���!6C�C���"��Z����Ie�dʕ��f`
����4e��3d�L+l�zPj ��[�����BN-i�|U���+9�@�*�����v�jH��(��O@�1���O�c�R-R"�%`����'P~�zCn�wՔPAa�@2#>0�I�'�湨�4t��%0䟟�}:���0^��AP�Z�\����c�<��C�e��3��J�x?��H������܆J��6\�>`�g�'�|���J d3(�f)��e�E�����,���P��u�h� �V�M�T%8� ��K96��J��Z?:�H1��<<O��I�}rL@g@���-]%��@ʓ>�y����#��Aч��c_��ɔ�ݘ'�ўb>��*˱M;��A�qmܡ(�*D��Xa^�X�����h��@>D��	G�D�*O�$2�`S�\{93F�>D�|#��D:g4m����/=�F9rK=D�W�i.�h�@'&�=��@:D���B\16��d[w�ݡs���t�8D�L��#ʟU|} ��YE�~i*�g6D���tj��No֍��WDJd*3D�� ��5#_�/����@I��=��$�A"O���2�k������r�0A"O"��Af 𘜻��N-&y�W"O�\3�j����T�A����F"O:L�$�Y�~\�q̜�xl$܃�"O���B�=��Ya���}]b�@�"O@�bb�� v@�TA���!2��q`R"O�i��M^j�%[p�D�tu�	$"O֨ �E2Dl8���T�c
Z0"O�8����'`x\ӄ&����(`"Ov�����_�`�@�0A�nI��"O��'eW�7��UG�����#�'��}�$�	|Rm��Ԗu~:!��'qހ��W��� a�^�$=p�*
�'eX��@�7>���[3�W�e4�	�'�j̈�d
Q�'h��l����	�'��I��3R)��#��^�b�d@�
�'��sD&�>	�rC��C3�̳	�'��Ě��|L�RO�<����'������:�6�r���93���'N\`��]>�]K׋W4�̸�'���b���K!ѫ���|��p��'�؅���JQ�����%Aw�:#�'|�����33�X����^�t!�'��iQU�ܐcƄ�+����X�����'5�aQ�� Y�X��>@�԰�'�4,����[�(1��f�%+Ef���'@�2���]R��S̑y(�}��'�{�!�H+�uj�J�$�"S�'����D�#K�Ĺ�Ķr���'���9�ȕ�0A���N�3����'4��Z�!ׇ+�x�@��cdP��	�'�b�i�P;�d�2��	*%`�#�'�uZ��U�;��U���,s|��J�'�,1�	�I2:(aHɂ8�Yb�'��m)���g$*���-}�0}��'�x��E��@92�̘&B��� 	�'1b�S �F*�����Y�j�T)�'�x�����S�]I��9�8g��2p�	T�"B�	���M���sL�2�H�6���4��I��m���F 5�XJUφ�+�|�����k6�����QRk�o!J�����y�&�$L��E�-Ck�x{Tf���Oʄ���6gaj-y��
 XTH�0��f�|B�	�[�Π�ER�V�2���ΰ+nPB�ə���Uc�\ib�(��H�0�C�	9l��Q�c�*x�b��܂�<D��թH�[2ļCL�� �qR�%-D���b&K8|�bl�V���[h��2�,D��Б�_�0��)�IԩOI�)	f*D��J��S&�pu�W�|�р+D���bԕBۚ�DDʯw��4&E)D�� !P�^���!P$���)��-D����o9�Qi�	�q���T�>D����6���a��ǀ��)J6!<D��
�L��(���R�\(b�8D�d�ǥ�3�`-åI�<~�\�Y�+D��[CHӰ�ذA�%<*^��� 5D����|m��c�0J)C��4D��Ӵ�ї#ݖ4���M/]K"�e�2D���k�~!\��� �SJm�#d4D�R�jF/}��������U �.D��
ӥZ�1 L����Ǹ|CڬHE�'D�,* ��Ă�e��Rz��S� %D�� ����D2Pk �cCJؔ�&�bP"O�00��!$d:���O9^����"O����l���Z1#c"k��1A"O^���ꈫv�j�Y`��3 ���G"O��@���@��j���:��A�"OV%�L��dڠ=:F�Π(���1�"O�(��+�4eB�k9S��X�q"O��S2�B���ʄ��}���qw"O<̘@-874�p���$ކ��v"O���I�\SRM�ŉi�f���"OԽ���ۆ ��[��55R8�9"OU�sJ�7$hQ�0��u��p�"O��`�F�c�=���7j%��z$"OƸe ��Ota�S'�#z�r"O&Djk�!:� ��(C<��"O�cjցh�}���ǬG|�$�u"O ]A@��@P��K�n�X��"O����%Z��1,D�;j��"O�1���5xr4y��.^*`AX%"Ot�3�X�d��K�o�Wq~�Y�*O&T��I.72h�'��/�ֱ�'��)��$X��i�'4$r�9
�'C�+D�B����V-���V�j
�'^�ٵ�ݥKG<Q�,�M:H
�'�:�a���S׮��%��:���	�'�n0�JY�O��8;��&xA	�'m.���fQ�	� ً׈�%~*Nl��'���&�=Z�����Ӆo���'_�ܻ�f���h�Qj��m& H�'�B��«�!Q9�Qi��^�P"��h�'��,Z'B9:=�Pi&C�)=E�ݛ
�'�ԩ�����6)s%��9��|*
�'�`	5��N�*)����
g�Ʃ��'�l�ȔY�6��e`�aQr�'MԨ0%La��Ae/[-���
�'�`���A�OHA*P�Y�"�U)�'0%��(=� a��AC����'���#�W� ��M�6�mfx��'w���6�����bw��^*4��'+��hf$��&��5Y��ug��`�'��<���f����F�6*	Y�'�e�q��/~�h1�v�ݖ��D��'�(�%��&�l�������y�'.�MbP ��s2fʽ�A"OL���	Ŗ"��8� ��==E�XS"Ov�j�@��r׬dJ�B#n(��"O0��`2x��u���9�&|)E"O�A3���3S���P�x��a��"O�0C�ۑSJx\���J�d��a�R"O:�@6A$[�`I�U+n�\�;W"O��X��S/�R� ��Q�/}��"O$���bںS���8#IM|�P�"Op`ۣ� 6�hՃ���,"ش�5"O�H���u��l�s�)�|�v"O�q�`N�;rb���`韍v%T�
�"ORT�t�_;���aȈ0d�5{�"O�\X�îa[��i�!�1�0A�4"OR�cq�޿e儬�� W-	��{�"O�-����(?�4 6O�[�R�yA"Oz�KcY>&i��֘u�>�)"O��z�H�$4'F�P���S���t"O&I��L$�
4K�.[Z6��"O���dN�v��qH�yV2Y�W"O�<�G�(}��I��]�`A�9z"O� R�!  ��~m�$��EɈ.9�ܢ`"O4��ç63��Y0P,G-�R"Om�t+X-Ҫizg�D�����"O��`�ʷ
Aj���&@�D<�1"O�ѫ�FV�0dl�(��@�}dؘ"OjtA����N�̓7�L0Gh�[#*O����E�jR�J�	{T���'{Ā��m^AF64(F-Q�P̭��'Ɗq�f�8/}�LZ�(��X�'�6 +�ć�5��"�F��g��y�'��Y���[�:n�t+P�RA�x�j�'�]���k�H�`w�ĝL)^`��'X:��Ð!<�|�і]�0;J ��'�l�hp�Єk�pF��#��0��'I0��P�ݏp��aYVO���rd��'6��"�T<PHl{�k��]��'�N��'���VGJiP4I]*)K\T�<ᡪ�,��C�bQ80��4(���S�<)S!�WDb��T�4&�P9��i�<)�aI7%��Ҍ/��9��T�ȓ|B�b��E���&̵&�NE�ȓ�$�J���NZ�d��L��fv���)R�eI�H��w�PR��չE��P����i%m@�}>DR��DH�ȓ}��H
�.�Uy��f�^ȇ�S�Ԋ%թs�)YQҢ~ʀ���ck<L���)B���`���7u�Їȓ/]l���ӈ/�J�G�:�6�ȓ2T�Eׄ.h\��6Dú ��Ux�Y� k�HH����ۜt�
��ȓ$�l95FH'J����o��j(����h�h�i��=Ovpu��kדiyh��ȓEhb�@�a:z.Ƭ���~\蘅�X�V�Ф(Q��roV���م�Ib�I.P�H�ଡ଼
^����H�({�B䉏4ۀ� �j�1iN	��J�&��C䉄;��h��A�,�*ъ��ʫjL�C��k�80q0�ŧ�,�5E
�T͂C�	�"��E�D%�*f�x��F4R2�C䉌7��k#KOd��8�1���<�C�IR��)ŊbG�DB�F*l�\C�ɶR��&(̘ISR\*3 Y'�C䉾,*`�7fK6(�����4"�ZC�	�{����I��Q�Jt�7���LK�B�ɟEf��Վ��96�jKj�*B�	� �@rb�)�����J�0`C�I7I�����"�&@l�h�%eʡm�B�ɓ;ҍ�t�G��5k����B�I?L5>u��fNg����  .�zB�ɑ�x��V ߥ	>0�Gŏ/.�DB�	�]��*�b�0v,  ��Z( ��B��Ad�"��Ed̤s�斀)�B��$s()q4@�1z�p�b��.[lB��6��(���f~ X�$3oAbB�	7MZF���hؙ*q�Ӥa�i�@B�	�B�P�7�̻(y
�i�G5a��B�I4<�:᱒V�3ΒԊ�@J�,"�B�	<{$�y�P�^k4� C拜ewfB�I22�\m�u�̅:�I����epB�ɫJ��5&G�9���@߷ibZB�dL�@bw�J�S����:ni�C�I'���A	�|Az��3'��NC�	�@d��-g7�A+FꙤ/[8C��bu���F�gdz=	ťX#L�.C�)� (��[%�HѣK
L����"O��
2&ē@���)g�L(1�B�z'"O6ѡ�݂D<�$�H��mL�T"OTe�.F��%a#ǐ�B|x�`"O���(Zn�±%� tnU��"O�q����-
����ǣYo8��"O���ԯ�w
rDJ� �c�.�R�"O:]�H9%	r�Y��c��a�"O2Y��nf/R�N����h�>��k�]-iS(�4ʛ3�L%��g"D���G�<8Z�4	M�2��:p/!D��J��.%����d]�B$�l�F�;D��C�l�&����C-�xGT}Y��,D��2c���kÊ9��ܡ|�.����>����	;K�ie�ʿ{�
�qCBP�B䉪>Gֹ�S����s����B�	&Т�ˀ/
�I*������,��B�	(qe�tR瀗#L�<��' �7ʪC�I)G������H�-�P�	wyrC�IB�$l�u�=�����MU cdLC��.uFf�g�����#GN7H�.C䉶`�x=�(�:���g_�fB�I�D���sOM�z�V����ٕ9�C�I?B�`�'�~�
�x�kX�kn C�	��8�rfΏ=��!g��w�B��3_�BL2p�M�	pRP.�VM\B䉢�$萵�_1D�(a#J�#y`B�	$0�v�K�bݠ�FU��ïi��C�	�s)��*���<C4E1�m7
��C�ɂn��8b�h^<�(�f၄DÞC�	�g|"����u`��2v�N�rC䉱;rL���e�@I�եX�AdC䉄j�&t�����#�v�Q $I JC�I<۴i�$"X�(�:8�"E�
bbC�I]�
��'���2��)�>�^C��
DO���'Q4&Ʋق /�LCC�	+bO�E)GiF(D��&����B�8�1���D�a�����O�Vt!�dZ��TJ4/B�f��;�@��,!�1�����Ï>B����P&#!�Dټ�4Hs�G�/��t��!��}!�$�5�艛b&Xr�8㳁�\`!�$M��V�Zc�Ii_4|b���J!�d5(:0����GDp��R�̕/!�ĊF�Ը��L���a#H�E!�d�OU2�ˍ7e�� �⨌�U�Yb0"O4Y#e�-?���(��S=I�8 ��"O��)�&\�c��[��T��X�!"O���WM�^8P!R�"�8[�05��"O4	˅I�Q�(����0�*���"O�9����XB�+��?�(��"O��VF޸Sش�;�̎>Ō�� "O��@��'k��@�ӌ o�權"O.�Ǫ�:�<(j��ͥk��|xe"O�y0M��r�,�I�B�6j3@A��"OތP��܆s�ĥ�vÎ[�xU��"O�����B�M��!�>�ҽY�"Oʘ����$T���`��i���D"O�� 1��3:t����1�BE��"O�l� N�����pc��4���K�"O�I���"qP���T�O?g����"O���M5>2F�i��M�/VLD1"OӗAL�U���%b��JF��"Ob��ʋ32��t��&OI:�D"O� 0��摀%�ԝ�����F��Q1�"O�芀bC�tVϛ�i4�]�@"OT�+C$W_�MH�n0~"��s�"O�ܢ��5�F���4x"��"O�9B���$: |\3�Kٵwz���"O�u)�떨 hhb����Pl�p"O��I��7?Hi��c&sV�I�"O��k���H�*�K��R�{�"O*��u̓�Ng�I��5}N	�A"O�Qi��`�HP�D)Zm��P#"O0C%A��kiP-Iصf����"O���������g�M�.���"O>0j��":m��w��1Ǧ�)@"O�����O��Q&�=���g"O "�b6f�`�ɑ��	�2��"OBi2�֙gd�Ԣ/Q3�`
�"O�PBЉ�&G�������>G���6"O�4	 v�j�؃/["hk�\Ö"O���&��:G�@�g�V)Si
��"O2�𵂄�_�HP�HPb�T��"On�3���/Tb����ED�M��"O\ �4(��C	y���vL���"O�#�m!��Y�
�<JZ�"O��zD��]8��Ґ/�*t�y%"O3��̠����9e�ѸS"O��A�@N*~���C��4�(	`"O*�r�B�em���a¿X� ��P"O��8�&X),�H�òN7u5h��"O6I��$��i�^0�\2���F"O����ֶRz|�0ei	<"	*�"O�p`�Y�7@�3��K�,F)�y��K� Ĕ5�,���y ɐ	�y�
�E�hR�o�&�H�CD�y�W�{�(��rV�Y�Hو�y��ք\vL���+ѧbo�Lae��y��5�� �/� U�t�ʱ�޶�y�
�1ohy�W�M������yBnZ�Ke0T�d���@
 ��` G:�y�$۱x-z�:�H\�3��;����yb+��Jݣ�JT-"1�����)�y���0,!�+A�nD��@�ߏ�y"�?g���0`H�}��4q�l��yR�4oU����8a�>|
�!�8�y
���Za~�jBMsh��o���z^պ��=. *م�Du�iK�G�	fD�ʷ��6�&��ȓM��<�Bn\)C\p���H2M���ȓN(�a�G�$_j��oRV�m�ȓ72rq��ZlJ�wѓP�� �ȓOZ|��Ck�@BBt(��طhBNI��b�Y��a@�^��A�S�<��^\&��E��1�֨����N v<�ȓrмY�P��Hs�<;�o�Ն�G5�Qb��(q\#�ܺpO���'B���D׬l3���N3STL���L�($L��e2P��)2�a�ȓG0���GM"R�p�0��&V .���[[�q��'�$uO��A�*`�p��/�&1��,��;�8�;Ѩ� '����=8$�!�J��s# �:�0���~�>��wZ���ū%���z$(`��l���cd�mcP��$��.�H��.��$��n�G�N�B�[�'����� �ܑG�O�n�� ��0��Ї�S�? %v��lv5���U�,�@�"Ox\�`nP9(b�Xc�ʊPB�"OjH{eV+x墼3w-]<DC�r`"OB��W��V�^I����{����#"O�t2��Y�^e �G/&����&"O��!� �t:�*�SQ1ԕ؅"O�as��U{�V@	E�;.��q�"O����ŝa[l�2 
���l�b"Oh��!��3c��+������b"OAQp-��1X��!�E�;a�3�"OJ��"�R# ���U��-<�U�"O�$5aO�[BB�� �|賗"OZh����%-޼�D�FO��J�"O��X��X�Y�n�$��h�:UQ"O���͛���| C4u�-I�"O�$��A�2vZ�I'���T�\�K"O�p�A%´|�s�/�d�h%`"O��ñ��']v�5Rr�0%����"O5���ʕESd��a[�Zvh�1"OMY7"��g6j���il<{r"O��r` �aK���+WȔA�"O�J��6h7��%��3(�"O�}���ܛd�|� ��E�u�3"O<��kԇ~��%��D��2�0E"OJQR��=Pj4Ѣc�V�,�А"OT] ��?\Ή���#X���	�"OL\,	��49�� :�`օ�y�"2�B]C���3�J<kI
�y�Ї;���B�)�+���dH�y�Ś/Z��i���#C0�9w,���y��;N$�Q�'��%�����GT��y�Y� $���A�� h �c��O��yrU�G�h(��|�tW��y���e{�@�vA�,%��Ȳ�o��y"	��n��)qv�S�$��<�tc��y5���%J $/,^�����y"@Ёe'Dd�R��'.09S��3�y��ks\\1�E
#9�$�H��y㇁'Є]U�Y�+�"a8����y"�K'a"���Q-Wsp��T��y�!�2q��tC�"�����X�yB�ß[�r� w�؅e��yq���yr/���b�ADnI0]�,ӰJ�,�y���fE#��@�N?��0!��y�F�:T���a9r$���ɟ��y�E�+1�������n�����%6�y2gCAK�x �$�kª �$�
*�y��˳*�b�В`�`�PE�dc�,�y���8Rː,�`�Nk�h��Kҥ�yrfK�t
bɫ�$���xT�A��y��ԪH����7"y���æ���y�,Y�g�qQ�שA�a��\��y�Xn�~0��W�=�@3⌡�y���q$vM+��.>��Pr�T+�yb$�|�0c�*�wB�T*r���yLX=b���r �O�r�fpZ1���y"j�8����Iԕ7U��� �yR킧������=,�����yҩ>(�(����خz�X��Z��y�KU�f�R�L�|�\$(U����yB�ӂUp��ьgk|�@d�N"�y"A�	 ���{sk�f�nD`3���y2���"mP��Z]�JcK���y��\�S��9yW��P��= oN��y
� *��fDB`���K�r�l��"OX0!wV�$R�\��.V�q��16"OjE�A� 	�nĪ�З�!�2"O@$�A�[�g#~�X5�ʙ)΢UѶ"O ����]ld�Rl>N��4��"O�5C2��"����� �<1�"O̽r�hL�L>����ؽN�IR�"O���э�6�\�5a����s"OV`1��Ż =��ZԀN�E٨d0�"O8i�a�XCOR�;ԭT4~�	�"Op`�΁������f��d�7"O ="w�]-L�*L1U��K��mH�"OZ�����3�
��	�
�ؘ�"O(��`�ѡ��izɡ2%3�"O"����?�B0S�ї7� ��"O(���l�#T���J�@Y�Oq�a�"On��K�,-Ԗ���h�]huX�"O@�B�抏
� G�o��i"O�y@p'ڜ%m����	JJ�tp"Od�8�O�#�9s3���;̰q"O���p��)p�&�C�@-O�zeQ5"O4e���Íh#w�!D�R	Ʉ"O�08u�
�'k��yV�_8l�t��"O�$��@�E(n8��F8}*g"O~�h�-Z4�L݈�@�-I*�A"O�*�Mѡw�^���` �e҄��5"O8DQ�� <��Q�n˚B��EI�"OZ8��EڰB%�Ao��T����"O��1C�U=L�~�U)�N�+D"O��,��$c���a��]�r�%ZD!�/C�]��]�E� Qb�D$#�!�Z�2} ��e�L-���q%� K"!�$ՎL;x:��U��X��x���E˲��1�ۯjYD�!g B�u�(]�ȓY7t����.�L�`��A��ȓ+̈́ʆ��[�Xy �攅�%�>D�����z1H����k(���.9D�l锥�����Q�_:j���!%D�T�F�@�M���j��P +X�3p1D�ȉ����-��NڴY��e,D��qJ@�%}�����f�J5D�����53�ĳ.�:�P�?D����]rf+�&#�"c�8D��Rs�=���򣁎X���q�7D����(-�V���Xs���S�6D�رR���4ȳ��/��D��n6D� a�II82`h�" 
[pl���>D�T�P"���A�CK�=��@{�`=D��(q��� r���n�VӪ`)>D���V
. jF8���0X�lE���;D��$ջF�(���D�S����+9D��p`�+W���J!�0,�0D�5�:D����l��F(��Q����@�j���9D���3�ڽ6`��PbE(#bIs�
<D�,"�]{�R 8� E�"쩠<D���V/d��̋��­j�i1n;D�,Z�,Z�Z�`�5��A�~�萭7D��XEAĸyޘR�m+I���a9D��ZQHS8}��"����y�R躔�6D���i@"b H��iU2=��	���3D�h����w{�9�c�a^�J��&D�H����/x���I�����"D�� �U�i�M rU�6L�Y��
"D�<!�m�nBѲ�CAZd�%�*D�� 8I�v�K�4}�M� 	n�ss"O�H���G6?X��,�9/��p�"O�\0rA�:[�f\C�K#�v��!"O � b�?�HbR�!��=g"O�P۔G��qc��HE�M�j0�"O�cE//8��Es��rq"O�*�@�8Ȧ��Օ{�"O�Aի��?��hD$�F�y;�"O��aFϲX�x���BB�S"O(��N�!�E���^b\��"Oz}���?.�*�6I�L	��c�"Oꁊ�'�&t���[�)�t��"O�����@���D�͆}鬅xD"O\��S���Xq��f�`䲠"O��*�I�����!��0z�d��T"O,�
P���C��Y�6�O�ΠP�"O6��i	^� S�EA�"O�ZT�H:D�D	S0��^Նm��"O�]b��#���:`��]�D=� "OrTHQ.R�j�x��VB׃a~��{�"O�pz#c�9N(Az0����4��"O܉c�D#)� �ń �iovYI�"O (+���	{@��:Cc��b�ZIkR"O�����:1�9B��	�xy���"Oh����C�Pt�lJAlY�W_�j4"O�MBr*��2K���D�̤<���"O��J��Lb  ��L�´Bp"Oj�HE��m�XSЬ~�
�"O��"MI����i�,X:_�� Q�"O<�G���S���4���h��"O����@Ч\��ЉFc֟S��;�"O���ȅ>+��%���ĐM�h� �"O$ѓjN������)1E"O���'X��h�"R�d`ƙ��"O<�VX��p�� uꜹ "O&P�'��?��,+���0�N9ɓ"Od�BE�0�2��� �J�"O�M���)l�;b]	L����"Ox���@|r!�B½o� QSs"O*���G�>rja�3f�m�%"O�聁���X�4��"��ٷ"OR܉%�B"yl��RF�P�l��"O�Q#�QT@SCI�;o���"O9��oE3�xB�k^`c�"O�X��3�\���`^�!O�(K�"O�1�#� �$���:M�h"O�5��҇i\,�$��V?
��1"O����(O�dla�#��*8���"O�![.ݥ`o:a`#�6#6j�*�"O�=2���:Wi���.d@X`v"Ot!�4�ˬW�=c ��H��$"O�M�fPsa�4S�i�
a� "Oz�C22�!�g�����E"O�`�%ǉpż� ��I�*��7"O.��PNY66j�Q�Đ��h`s�"O�t�S肠P��x�����ш�"O4[�.�x2�q"��	x�<��"O IK@$//�����..�p�{t"OH]ɳk�'ck< �РM#˞��a"O 9$fա�ŀ������U��"O֘	C��(�f�r���u����C"O�(Y�g(	����nW[�.eIB"O�a�f`�G�`t`6-���H8b"O܁k��(
�%q��)zp\Q"O� ����ۥ^k��Wb��e�4�p"O6Uz �%�,yiǁ��sh8�4"O��D�0�T}D`н bp���"O���@��x���� ��.f��B"Oܐ���$h)`�(� S�t><�1c"O>yP�*���z\�S��%&ʲ�A"O^�h@��M���q�
�'� xJ�"O�#d�ϫo��(��V;JХ	�"OB��'��(04�p��B�Aç"O�q�2
G?P��`��'iA���S"Of$#�j�#Z�Lu�܎t0��
�"O�����7cH��SW?w�Q�"O|<�G"�LJJ���6%}��p"O��!��8n�AI�Z�80	�"O¡h�$�a�r�a�M�il�#"O�$��,ƙ|�ʓ�G�*��h�5"O�Ps��t��*s��t�@
d"Oj�@��僐�ǹ�rъ�"O��(��\�e�n�����j�
="O�yA�ś@vd�$�7p�vpK2"O�9qƯ@�D����u�;�����"O�0���@		'���ނ5�(��"O��X��	^�FiYS�H���/D���(�eT����ֻ!��S���OC�� 9�5�7� 4�m#E��y�B�$�����oU�BO0}z�̎�u��B�I�W��0��F���C���i� B��	t�L��g�"|j�D�f�)&�C䉨)3L|�Ȍ;ˤ�R�A���C�I� ���[ӨH�8�J��Cy2���D~�4F)L/3��Q
��U�p�+�@�O�B�	>BN� �
�N�"*@C�J-�B��&0�U2��M�e��a��j��`�FB�I9m���j�	Y�E�p�w�#2�~B�	6s��$ ~*�t
ݰ/�hB�ɹS� ��#ݱ:�(�G�_��C�	�a��;h�uzʍ��߱Dθ���<?yC��\��Tr A6/� ɧe�p�<	�h�V����"K�{;a��-k�<!����A�L}Rc��'b̔�֮Ig�<�FhP�0�r1h�ʎ&\>x� �f�<��˝���uBG%E����^�<��J@&d�j�YEC���I��"�W�<i����}�*Xe �(w;l��7�{�<I㥏i�d�CO_��<tj%�Sz�<q���X� t�����H��kA�<!�L�B����$lўim)Z�Ȗ~�<���ϖ0�bY0� �0Zz@@�MLF�<�Eɒbx��g���{�E��<9�b@F������)"��90��Z��8E{��)M$h[�|Xn�f�"���b�hM�C�5	8��	C�H� u�VmGd�C�	}|��[�Q����J�ͰB�ɀg�p�R3��
Q���H��#P�B䉦/�,=
��"E�3�Ū'i�B��Cd�q����F����m�*fߘ���8�I< ,�d$כf��b�]�Vw�ʓ��'�?X�( ca�M�"j��@#D�PX��UJ��!K�1KJPKS�-D� z��>�h����ʜe6vPc7D�*���%8�����I�8���c�6D���tʃ6g܌1 ��Ƴ�R(0�"D�ȃ�'�������#�=7Q�ᡒ/><O��d"��:O��)�&M1�$��/[����hOQ>� H���EW����/����Y"O�M��B�!8�A�1�V9��T"O���o��IQ0|h*���!�u"O i���܏)���c�(.�� ʔ"Ov��b�B�l��x��]�x���7"OtXiΎ]���bϕt�4�*!�'��'��č|(qC�Ü	mt1A���N��'Gў�>�b�&!�Ĝ�����W��E�g�4<O@"<1�玓9ǔ�R��F6�0�n@�<��l�G�4@�M�5�r9Y$�GR�<��,'.�2p/�o��;��T�<���?}���"�
�T>PQ�iR����:�B�ᅰv�Ɯ���U�A�ȓ[�r�I�K�d�\Ur��O�H��T���D�Y �?.fM"S�ɋk�����i�@6k�7�`�hS���N��ĆȓBv2�"�ǫn�؄G<ˆ���S��) �҉-����Q��^>$��}���oFD����� �	�ȓc�&R<2�Pbτ@� �ȓu�FTZsD\<y �ػ����̅�7��Y�p/ֻ=���[�1;��ȓ����RB62�� �Ԡ�*c�����:�n�A��[�J��e�s[�C�	:�
`��aY`�Ak!��C�I�ǜ� ��3X�8�[CK�m����*?�Ц�4OM��Ɂ�~���h�v�<�C!ֶ'Z�T&\�Z`�؀C}�<)g�ߣ$�Y	����p��fOx�<IE-ޝ?;
�TeE9;�t�"�X�<�eM)9��Xx�Ο21�2ps��S�<s��VKX}��
%F����N�<AR�*��`���\�8�bl��Lx���'�@���IG�옆@��z4v���'ܾ�c1n��B�f�Ze@�'�R�H
�'uV�`���Pz�p	�L�2S̘H�	�';�h�b(ȼ�����+U�R�(	�'�����JNU��0�/"��-��'g�EC��\)2���"kH�B�'�)$	N@�N�f��09G�t)�'� ,SB�Z;xF��RlK�,^<�'�d1� %�-��Q��!��s�'|��2%ES!
R>1��b�_t	�'K�9V��~T����є�.���'�Bx
dj�>28�e�	%̭��'�܄P��_�{ =3f�ҋR��(Q�'��+��Op{����FͿu
|D��'��\���(HY	:"\.k%��Z�'���PJ��%���bk��L/
�:���y��U(y��*�ˊ����6�?�'�<͙SꔞD�TA`��;�L\i�'I��pR���-�j�����%)�1�'�Ui���lI����E�& �9��'�`N��O��U����	 �^dX�'}00#�&�TZ�q�c��4�
�'�a� h�nf�E�W�H���
�'.��C7l2:z,]�6 �/iv����'�!�]-�*J�? ��XcC�{�!�C?_�����*J�%��y�AA�	�!�DQ(`����8�"lb��
�"�!�d��>�d��22�T��X ~�!��o۪(�jV���p�Dӳ:!�$�;#	�	���5�����^�7���'v�pU���F��!P�	Ex���'N!�� �0ieJ W��b"�۠6B���"O�d8�jN�P���'�M�X�Q"O��Xv�I�Y)�e�`֕04"Op�j�G�.�L�/�O���:"O�t��Ǟ�I�Сz�`Af"OFl*5Ö�THy���_lV�	R"�'a1O�<0@�΅L$��q�(�49bܸ�"O����%fn ��	P�J��%"Ov���Z�e�(e�W��� �.�&"O��"��Nh�+D�:�\�C�"O$LQ4@�QO�1��$|H�@r*Oi2eb�T���f҇.�hp�
�':��E&��`����R�]z��(
�'� ��',ϸ�y�a w,AI>��?l������_����c2'{�5��On��cIO�K_Xɣ�b�6\��60LT��)�!�܉�u�Wtyr@��}y 홑 F�,��`?Ml็�[�@U�acʄ21%*�隽S��ȓo�"��-N<|L�F�^?H�h��ȓg��!�҆2?�$��:W�����n��@CqCZ�j[�PRQBU��*���xF��x��� �zyi��H>��ȓ���0r��(V%�G�Z�;!����&�H��\=^�v9���7@�Nd��I|~��D,B������7\@�� �y��ͮ}~|�� � :
����
�y�	
�o����b<]�I���מ�y₌,�� ��A4}�,�aW&ϑ�y�d��W�X$�T��=yĶ]�V�_>�y"��R���h"����jk��y��NJL�b
	����2�y�l���@e��B�q�����y�k�l5h̐��*?� ���jJ��y��S�t��|%��0�"�C�y�IC1A⸀qg�-*6������y��
��٧t�\1�քX,�y�[�� rFbV�f_^a�a�D��y�dC�`��萔h\�-����q�ǁ�yBoT^�<)2��ڑ\nz��4���<�O��0D�L�KsD�@D��"*X�[�"OTA�7�C7/���)6�ۜ4Th��%�'�1O��y��R������!J;$��S"O�$1r(݌Fp�h�W
�qH�"O*�Z����H0N��gY.j�ęR"O�l�p��&u�XI&!�ue�\�p�I��|D�"]�$�^��S��.���r�;�yҀ�
>��h�#�ߞ_,�QE�A��yBa�6�������	$�1d \'�y⭅A��1�����0ɳ)���y�$[�~T�9�S1 吕K�	�y�A���qc$Ѩg��`���y�h'.:�p�:\�5�'���'$b�'I?��)�*[X�#T��x5+w!8D���b_�r	�c�B�hꦸ��g4D�0�.��,+�ab7k�^&:xq�/<O�#<ѠN·TV(1�g��g�6����V�<�O�'��{WAK2�^8�ǏU�<��GS
T��4+-�0Ѐ��h�<���#R�d� nY�W���T^�<�ҠK�_� ��M�/B�D0S
�q�<�t�}P���"C74����I�D�<�#�8p��0 �BG�O*����C�<��ʯ� ��DB��Θ��gA�<� ��#���.�q͇�')�i�%"O<�uꆥ4Rb1Ku�ʤC!����"O%!-S�|Q1�	�En2D�@"O�2 �WJ�(��%ܕVz�q6"O�t�qah"E��È�IܶB7"O�@����ZE�F��.	�U��'��@��,�Y`сQ���An=�%&D�\�M�*aά�7jT�#��d*!D�\P��+����#���+0� D�8�!B�Ğ}g�u��"��^�v���'鐩su��?�C�	��S2Дk�'��ac\Z(Eb����R��1	�'FB��t Y�]Ơ�� '��QHI��D4�'<6&	j&+ܯ�n��a�ˤqb`ńȓ	����q�K�xJ�`u�C^(bU��~� �6�@�xP���5�t���ȓ?�H�ʔ�2�Y��  J�f��ȓY �5I!�W������#$)|�ȓW�0����Ҽ��A �ʟ�|��M�ȓ(f��
��D�t�Z �a� �%O���zNH͒rɇ�$H�����$P�}��<=Z�ȡNW4*�`ځ�dN\��S��<S�!�y��T醄^Pwؙ�ȓ;�ڡ��c�?;���KP%M>��ȓ~��AA&&Q�C	�tPa

T(��?�LPьF�Ҹe�����{,�I��/픑 E��x����7�E�!�	��	�<��1^�����I�-`q.Z�<�r(U�/o�|����1sw���w�<�s%K����B*��9&�BB�r�<��gʝ+V�2B-{�jc GH�<����a7<epbʓ�OVt0C6�F�<9vn�%9j��e	��Z�*w��~�<�1�İr�L�YI|����y����	�A���Ӎ֙i-���UO�!jY$���Z�)y3�L�(~�b􍞠 �����U�q�0�}$�F�U &�ɆȓM�d]��/U�d)@��	V���(��Q36b�6f|�[�f��݇ȓ{��1xg���+�ܢ֣A�>d��ȓ��4�&�R�E���3`�H�Rô�ȓL=0����e�t	 ���|�Ȅ�X\�K��'H<����I���ȓy^�1��#�o�Tl�p��4�8}����(Ak�&��;��ɌV�Ɇ�+��,�F2J�*f�܇N��ȓ/Xм14㐑&�(����d������k @��y��h�&ܽ&���� ������ڨ(�*4�Q�B���؄�ey�<C�U��y���N?~��S¦a���T�,���tKJ 4��Ňȓ.��0�"FA'FF�����؇ȓ;~�C�B��\q������|��jbtB��U�\�^u8P�De�ن�7씲�.�q���M�x��(�ȓ�D��.\ A�6i0)Uh���ȓ;=���a�͕k��x06�Ԛq�*��`�f�S�F>�T\P%#Oc�Ї�{3@P�n�"�>��It2^���\Vi�%�ΒrE9�1(Ar-b�ȓR��yg+�
|נ��D#TUB蜆�p`�$��/L=1:�L����l
�˳ ׿=��)Äg7>��ȓ}�J �uچ�v,y�j��V�6���S�? ޤˣE�j0r�@R	њK��})3"O�P��
�^�b��_� |��"O����&ƭl=�ͫ��"'��"O\��䛱S�����'�(��0��"O�;��,o-��ef�^�j"O��e�R�m� ��>�4X��"O�T�p�	�,������h���HB"O�M����*����jH?I�l�s0"Oҙ!���;
X�5@Ëx���b"O�E0�NK7#�����J.��P��"O¸���#jU����K��cJ�D"O�=�7�>1� �p*��H.��"Oj�8��P^2���E�Ҿ+�e�R"Oxl����/f��U*�ˏl�](�"O�XKǅ?\���f	`�͉�"O �g�,EB �A�ӅLWZ�B�"O�	A��Z�5Rp����@��0"O<�@�?5Ҡ@s �!#.��U"OH�d��tnX�!6�pL��`"OZ���'K�V�����SR�TÓ"O%�uᐽ:Æ]�&�Z
RO��[�"O��{���F�$�H�n\�L�ƐJ�"O������dy��˴MY�l�XC�"O���Ю]�#�|�t�O�� "O��4�Cʚ��� &l����"O�D�q��P&H̪��μ[�$�!�"O�)2�"2n1�ha�_�Qv�:b"O�AS�W8��t�1g��+�{ "O�Tt�
�|A�t˱�K*"��ܙU"O����+��h�B�qW��<W
�pA"O(�Җ  $(���ҀED�0@p"OE�a�%Bwd2R�<�a�"O���0�ɪv���Rfްn��\S "O�=�W�_2z"~9�F_���̳t"O(�����m�pD���h{�"O�$R%�Z�R>1��A+�-$�E"OHH�iӠM�|�북�_m�r�"O΅��d��z��ψ$_�Y:&"Opqr��=H��M $��5R����"O����")L�D�F*��=<��R�"O�lJ��-V�(QSB'��"'�+a"OT����~���x�Q�u�1
0"O��������Cd�=j��a"O�]��{~�=Ra�LRT��"O�M�A�˂,,P`��a,8���)@�|��)�S� Db�&�?k0�B��t�B�IX�U���hQ�����]�]8D��ȓe	T9 ���`�0	�q��D���ȓO5�e�*���n�)���7D�4�2���Nl"�DΥc[���P�"D��IQf��.�FPk"e4vt%���4D�H�#ݫr|���+*Nn!H�)�O��ģ<�-O?��ɳ)�Z9ñ怅4z�݈�D�bx�$�'|���#ƭ;��YB ��8�ms�'���q�a�1C2J,IFAԜ�R��'�Ġ���D�% ��N�T`6��'�)d"M�G�tU���N;�X��'�%�w����qj냴@��t8�'��$��� oR��J3��G`a��hO?���k�k���{��
Nf�u�ҠJjx�p�'A�L�ì�	^J��  r��Y�'�̘H�㈫J����Ñf�v�X�' �Bed��#�d}+TDT�l$���
�'�­��E=��;��[>g�PD
��� `؈sHMT��|���H��xk�"O��SDH!Wu2yr�#K)����"O��	�1j������Y
P� �7Q�|F{�OR�¥��W[P����	,X��G� �� �S�'<]XD�V�H�R�@GF=�*���BD��VBѶ)y>��ĦR&'�j��ȓDR�,��a���ׁG�7Q�ԅȓ^��4��!�P`%Z�I4���ȓX����h{��5x�.-=N¤�ȓj�U�E.���`%�"cr`L��>��̺3aN4JJ�3�� +�dp��x�	d����D�>eZ�-��H����6Q/�C�	1P�R���Pi�TAe��H��C�	*=.�q)P��0~���@&�35ȰC�ɇs�\�	w��}<d�D�[�.�vC�'l0pALT�QV������:C䉵s� �a���q�PQr���*��4�	|t���g�p%#A)����@�IY�	a�'r�$� ��`.��J0*�.W ��� (F�5��W=|(���W,W�L���H�ܓ��?	�B4� eT�j�����U���BW)Y��a`�ĝMWp�ȓo$�&��4i���aW�3[8:��72����L0l�IP	-y�f�ȓ"�*ݪ���l�����#�F�H���q�P҅h�:g���8`f�;oɾT�ȓo��-�"f�1�`��Ed䠄ȓHS�0�& +?&l
*]�[bX��6V��7O[}>Q�toR�I��4��G�4Q����?(P�a��D�~�@���}���Xq	�+v,�u�!��
o5���ȓ-q&H��<@��H�o2�
�*D�`a���]��Z�����V�ys�B�ə,qV�X6&�!g�x����_^h�B�I���f�Z#���c� m�fB�	�g,���Ȏ!��q�
�1du��G{J?������n�H7 ��1<n�?D�P�Q���Q'T��͜��|�"8D�8	�E͑c ����a���D��F#D��p�*��B��x�e�S�hx��.D����-e�UqTꞄ�P�E�-D��CR�ц[�<b� C�t�Sj8D�T{&���O�\UI[S�X�Z�4D��	nʞl���j�!Wa�.h�%%D��BmK�r�����z������>D��+l?F���
M��`S�	��D<D��"��V8��\�s
��f�#
<D��#��G%�z�r�?ybh�K�9D���!�LY�U�&d߱eH]H�9D� ��k·Lr�9* mދ`O��I0�5D��Rł+O�Ȇ� �Q��]���4D�D���%�h��n�Sx��Qt�%D�<��d��{Rp�郧]�\��(8D��G�&'K �����c��h�g7D���$�{�d�Oսaq��Q��4D���F�,�5��+��	���Qd�/D��:��I5�͐T�G�?x����f,D�p`bJ��H|�DH��*N4r�01?D�<��.�'�6E�S��(
�Q,)<��7O��A�
&nW�ܪ�U>��`D"OV*�޽4������^�=����"OlM`Ra�I�歚r.D�!����"Ob��!�x��&�T?)��,@"Ov)As�F��� 
wӓ88zh��"O� pyi',Ⱥ`� �LT!..� Z�"O�P��Ƅ4q�h ����QI2%�QO̸���BJhi�����W�,���"D��
�� �}}���@��7{2qs�*!D�08����hza@�e�<Z�>D��Yuk�|�Q���;.����8D�t���P�+� ��"eӝyo�y@�5��ሟ��@�ˉ~:�jS�W�oiL�Q"O)�7��Ř-H�"YƬ2�O6��cG��Z���E��P�Sԅ<D�تGBw� �z&O@�d��:D�(��I�t��D�r3�x��;D�q3�@ '$�I��^�>r��a�;D�Ԣ�M(6�9��<B4P f	$D��*�ɟ+D�b�k�eM�a�v�>�O��N�|P2G���F�r���/ԿvY0���w<!�e7
�!�'�B+��4��	X�����أ��ŕ7�H��Y�/�h�/D� ��B��n�~UbEB��e T��-D�8i�H�}���aK��}�8�R1$*D��Z@��������[���4�%��0|
�G�	[1�u�F���L����~������Elz�����r�*�C��Vė']a~�kQvvȊToهeTZ)������?�I>������ɮ#�v��	�~p`����	 |B�	�jx�-kwFͫ"�8�ɴ�VڦC�ɫ��=��k]#� "cN�?0�C�ɘ#���{�B�K���H�� �*Y£=ç,:��*0�Њ3@D�q��дm��ȓh(N����	H�ܠ�G/Q�Z� �Ɠp���q�.$	l��R<U ��
�'�jQ��G�`!�I����@p�'2=��`���}cզF=�đ��'��5���[�Mp؃���9�>Q!�'7���Ď*"P̽3`�Q:6W, ��'�Y�BJ#W!��ɷ�R����S�'_����N�;��L!g��x�<�[�'~��Rb\c�pi#GX���Hi�'Q��(�IҸ�b�����/��c�'���h�#��Ac�Y�L�;pGv��'6��9��&vQv@[p��iF���'�� e��4u`�P��*1bѢ�'rQ�g&PԘ�ס�)sv��	�'ܺ=��CӪ8B��0nPɠ�'!����G�� �8�a
�m�¬`�'������}ߢ��P��
m��Т
�'���Ď�$a~j�ذbU�:�
�'2�8�F��$�@8y���-+@���'��hs�[/%%�z�ŉ�2�K�'�Z�	��z1��"�~ �'��1���9;��qB;s��]�'�f�YC��'�v����ٟ:��ѳ
�'<�(��Xڤ���Iϰ�ԥA
�'��䒡%T�o�8 aqm�~i�':�Бm�8p$4��uhۖjO~���'�@%jb���dE��)6)H(S�'B��mնf�`�3�>N�lH�'�ڜ֦�yX0
կ{y���'VHX+�&�P��,�Dn�o�d�)�'��Y�P�AVn�(�a�� dܖ���'K���X�.e"}@���kR�;�'c.��HPS�pS+� ]����'��(��K5�)䖾N2DQ�'����NΝo�����G%�T��� B1��A[l8 �*�+qֈ�3"O��y�E�;:���WJ׎d���"O\t{�MΒU
�"�X�T���"O�MQG�w<��C�7gӢ�`�"O���&��>4��ܛQ�<�yf"O�q��;��aah�7!�Lj�"O>Ԙ(�T�f�2ޠ\�}b�� D�pC�#�'7���!�}t*�3��?D�\9 R�Nx�}�eB�;`�s�/?D����[5y�(�k/C1'
J��"D��U�;6�N�Չ�%%����n3D�܋#�֣+Ҡ
5睃��q(��4D��@v$ɍr�d 7BvA��(.D����e�-��Y�%�D�m2M���'D�$2�T!'}0)0�޶9�f=QL+D����^�!S!h���W ���PM+D�б�h������B/�:�T��P�'D�T�1�P!M� dj��
6���)�8D�0R�B3?�la��僷u���db7D�S��=nѾm�⁠��"�rC�ɣ!�`<�7D��}��.��4:�B�	E�	�C.�bb�9��ɈN~C�	5A�fa;�솛fV}���D�w3�B�	�8�f�s5-ϕD���aĞ>lC�I�6�B���'� ��8�BO�rb�B�I�>��X�K��l���BDM�-�C�1 ��5z��.a< 3�*I�QZxC�	 7�b���HXk�HJ� H�7؎B�	_�Qe(Y/���S�[�f{~B�>�>�3�c� !���:с�P�B�ɵJB��25�.o���&תnބB�	�&z�@p��$2�r�GT�5PLB�	&��Z�"��)��@�:43BB�ɉ�v,�Qk	`�Q��
;.qBB�	
;�,JgۈM��`Z�}B䉼B������7�|�{v�8Td�B�	�YCl�Iw��6fc�ѹhJ�B�ɡ	��x�6���\��*�ę]δB�ɧD~� ֫:�am�:2��C�II�QP�/V��,y�AҸi��C�M���箎�)@`5+��
�	�'O�(��R2,�4�C��gK���'�  ���f(��У,Ih@�	�'���h����Ѐ��]kV}��'�� ��o�P��lO&g�>��
�'�6E�&!��|�:de(%gN�z�'��0pqg_�0�"()�Z^4��S
�'���ka��'&kX�Q�lE�[�t��	�'�����ڜ7�u��W�+ �<9
�'t��@&`�,&��� �Up�p
�'f,|C�.ʃv�Q��훬�$չ�'˺�Q���<�ĨuAF	l�
�'Ԁ�r��J�xD�����
�I��'
!BI@�"��CRϐ�~�`�9�'�DA1�ͧAY\l	�̊�F��r
�'uTtH1�=3u´u'�<��u�	�'>�� ֧Pr���#�爩2m4�	�'�՛��= ���3D�)3B����'�AEc >FR�[3 X�w|��8�'��j$��1��h�5	��F
h��'i��p�o۫YY�,
��B�>���'af������zudPc�H��e��'Z[�pIM�b�Ap���b�'ne	���S�ش:p��uNe���� <�w�����0��EP�v ��"O4�x�b�?J"�*���#��Lz"O~T$�؃e���ɑ�
�s���"O�P�b#�I܀�K^�����"O�1��.p��ا�G�!��M
"Ot��ȃ���	s�ªob���"OܔX�H��Dm�Lc��+ae.}!'"O�x���:y1vȪ(L%8]b�SU"OJ��σ�O*}'��TB���"O�`!E�g��F�WHI6�[""O�IS&��,Hq�<x"$�F�ᱴ"Of艒*��[|�U�BC/1:�V"OrQ(Sƌ�8�r��0�p��x�"O�"5 �4<P0����@$I"O�	pF@�\�~PBf$�<}G�Q"O\�hPk��.�Z,rcR�_�Bq"O�(*�&�
��IB��������"OX�p�*Cc�<i !Ť�<��"O��*��ҏZ�L�O�Mon\��"O ���	D�s��%�үÕ�"�i6"Or�S �f��YE(��}}�pS "O�)�tM<2v���Gȫ:b)r�"Or���H�y�&4
6�ջc���A�"O��A�ĝ$2��4���,�N�ZF"O�e�!O	��xR/�?(h�
�"O��8�ڷ:���N����a"Ox�J��E:H!�P��f��j��5�d"OZ� uh�1�� �P���i"O�A��m�ތ�4AݭBW��r`"O3����$��[V	�w)D��"O�1���ڤr��L���Y&Raq�"O^�Ӱb�%�r�Y�쎎8X��"O��"ޭA��;0I�=^� h"OJ�ǳp퐨`�*ōE`p�"Oh�`R5/`%�ԧ��\����"O�mJ���Q�\F��J�X"O��S"r�9x!G�9M��Ջ�"OּC��ں+�"1�̀	�dx��"O^��fOU�&9j�½&:j�jU"O*�Pe�C4Uh���Ƣ��A� "O���5c�$N{���@�*�"'"O�����t�tP���&^-�M�"Omm���dbG?3�<�f�&D�XkS�Ak��x�Jĭ >f��R 2D�l`uo��a��Ѻ%�×B�lik�(/D���4O�}�`ACw�B�9�M�fG.D��7c ��.�P�H];c��3�9D��!��n]  �pIjF�TT�!���>�8��)rb�@���w�!�dG�x	�A��"7�h�d�� |!�ZW���A@P�Ȍ�"�c�:,o!��J� ���+M��0��dg!��rP�J�e�����)B�!�P)�i�e���c@"�J����6�!�$�j���5'��z���y�.�(u!�dZ��*��AF77�Jd�r�=^!�²kQT�`%+�)P8PQ񷃀��!��O�V����C9U#N��W#]�:E!�T�Ud�lrW)�%\�6Th�Lʈ9!�d��k;��qB��6�,T9��ܐk!�dE ���J�fD�Rx �u��Q�!�4u6�%�#��3f��$�ƫ��my!�[���@ю�7.@Z��G�>_!򄆏)�<�ᩑ&�EGO�wN�|��S�? �}BW掍05�ȃ�(\���"ORaBA^<A_��3dG��7|��C�"O� ���:r�+4F�>�N��"O*4$�ê��R'A�L���nT\�<!`�^�&I����� `�0��l�<q�dZ�2����A3fB�e�P@�<��
�&-`-x��
Dpب
sMc�<�!�+jU�$�-c�,���j�<1�KS�]�d��Bc�]���w��e�<Yae�={���"l���K7"m�<i3cL�G|�������P��w�Kq�<�V.�_L�e���d����c�Yu�<1h�([�4�*�!�L6x�5iHh�<Y��G0I�Z�
��Umn��R�N]�<�b��8�VP�e�~
6Dȴ��\�<�GŒ<@��9A"I��M8�D(q�	W�<�E�wm���莠.�(�DaVO�<a��ϩ~5�(A�Ѡ̼��AŊK�<�Eȇ�W�r�Z�:��� b�<I�(.Z��c`����B�<ɰ
� /����hV��}���<����lP�t"wB��'�F��f@�T�<)��k��򌎥CR�"���Q�<�2/�0�l�t�õWdI���C�<I�&�Zz����F��Wgf�)���B�<Y��đZ?
@0#Gϡ�y��RS�<�rN������@Z�_*�
fO�<ᅃGJ�n@��"F ��
��P�<��,��vRA��O�21���N�<��˄Y}����N�� i8��L�<�hs�9i�����Y�Lb�<)pK],�HW��	e�A�`��Y�<��gό~�>|9��$�#-�P�<q�*%2T	�	U'��P��
L�<�nO}%<ܪ�#�(ch[wd��<�f�
�* �+��#��R��C�<a���F�; G��v�vPb���d�<bI�@�2���#8��(CR]�<)��&5v��7���=<�	z4~�<�U��&6����5��3�"���EQA�<����-Z�\SHB$?��Ղ���y�<I�o�58�
hAw��V�1�Y|�<�΀d�L����J�
����s�<��ID$Kj�81�#����m�<ɓ`����$bU)ezꩳsk~�<�C/O��p�lE�4k���W�Q�=��C�ɔ/E�t�3Z���#�JO�z����P���4.7�	�P�M�7ń�z��D��L�9r
�C�	��\t�Ԫ�% ���\Y��;�O�u����%1��b3��	�U���ƀΠB䉇k>�#V�T��A��-�B�ɼ*��,�e�� e�]bc� .s�#=A��T?���
8~�Tz!�D�8'�����4D�H���,I�.�@	�)6g��d*3D�p�,��;�E�(ý=j���X!�d�.ZSR��
�b�&�2Nm!�dۥ�h8�SjL<z��h�q�
�f:!��ћE�>l��lɑC�X�c��`+!�D��D�=��f�#e�>���N��!�䊥9j���&�,2���x�7!��_��Y���w�nq���͸X!�ڿW|Ha@������B䭙�mX!򄅶+_0�P�E8��A5b%R�!�� 씥����-F{�Ic�Js���=O� Rx�2)M�(�|�:t�7ըICR"O��KTB��<QܼɅ� J�0�j"O)���4\�H��u��҄C0"O�$h��He ֈ�r	� #a��p"O��*�7�ތ�@�P�e^��I�"O��sa�2�D�1v�G�?�2"O� U8=8��R-a�p�"O�՛b��񦰒fC۵P�e:4�ID��S4��U�|�OE
�����*D��øi{�Q4"�p2�$�)�h�<��,�K�Hj��A�"�	�d�0'�,pAR�f��ǐ	@�؈�d,D���CA�̬����*(�V�8�,+�s���OU��ǆ�>V;�YP�Y�F���

�'Ҙ�A�cV�'G�IR����z��2^vX�Ѓ§0'����r͑5��u"8D�܂-��<����,��9��th<�bF�$�x#�@�*5����c�� I�{��?[���5�ǉ`�UXj�-�y��6/�8	A���RcP���Ѷ�yb�L�)p|Kv�G�Qff��e
/�yb!�#f!h;4�O; v-Дǋ)�y����g�P���*�� 2'�P��y2o�U��#��!4�a1a���yb��6$�R@!��%!P9��·��y��[:�D��Ѣ�#��`C�y¥#t�A��\�!�n}�b��(O^�=�O�F�j��L?��(��,NxE��!�'�`8*#��&�rD�ǋϧ��A�7+�����d� c`��ؤ��u��'I!�H8.f�+���݈TX��|�!�ċ�)Q��25�̛%��	�AjR��Q� ���z����U�t8��@P�Y�l�!��Г�y2�ߞjx1[!c��$�S�S9g�����s���U��:�r�#i��If�<a��7�Ol�'*
�)Bk�� �t��z �Q�'�B�'���)���9��	A7�P�iG8z�'�n�X`�J�#�`�#)t���r�'�f��JR�r�r`BA�j����˓�~|R�F[��h7��.V8��%��y�Թu��@�B2=-t��H�5�yrh�1�� �bC߄3i��i��A��y�D��2��(c�=&1x��P`7���p>�� �8�� ��Ǒ^�8Yx��|h<	���9Z(���)ҏq�,�C@��y���'^s�l�d�  ��TZ'�� �>O��R�]�CI:eõ΂&V= �pg�?D�\� m[�Ya �k�H���} �<D����"��!5&����@������,4D�<�K�q�\��I��3!��B&�5D�8j'�D `�V�8O]��H�`3D�liĈ.@tԼK�
���͢!2D�a�`O���b!�����-�D+�O�=E��c]�U��f&9C����ڵ:n!�d�cMH�(PE��!*��ʑ�K�O!��)!��9q�=zp���K D!�d�O$X�k�
V�� 0���D��"OD�x��.D|�b�6# ��p��I��h�����@K�"(D��-�-r��pa��̇��Q��k���J���(��O�g��]���|r�
�.!��a�u�T�p
*�	S��t�<爑Z2|=	���J&�+S�n��0=��*�*������"������@f�<yQO *0���9���	:%��0�K}�<� 	���WM|�*L�b����
O�6m �$:>qb�����.���@�&6C!�d^,�����U+�@P�lȄp�!���'����K�?ۂ�r�LE��!�$�)c1peHcC�1ud5:�́�>I!�$
&�Y��jZAe��C6��E�����\u(E1A��������V{�\��� Pd�!W�L:������W�O��,"���	o�j��C�ȱ4�`�ȓ��4�tMѹw+@d{�+a˜�=)bM8�S��5`�l�E�P� �xY)f�&��C�ɤIe��!J-a%X�gO�O� L���D����2��;M��5�rjU�&7����wV(�z�E��3q�̻ᄓ\��1������a��)Su��u�L��9���Stb��N�-�5�ft^��ȓc��ܱ��� 0��)�U7��:�O
)r��A<�TI�[�X;8q2T"Oҵ��,�7<�D�bǂ�U?��iS"O������W�my�o� $\)���/�S�S	<0�5�w*�uz��0e��^:�B�I-L��a��s��U�c5H�NB�ɫU�R�IE��*���I�/:��C�7�X�K@+�@�,��T�egdC�I�t�d�A��>DY} ��O?m��B�I*H���r�I<	&i�#�	0GXB�I�ZL"��&����x!B�k�(B�8G��G煿������&�LB�	=*��Fa�"tj��ӅކL�B��7�2�8.2�H�Y��B�	><H�4�ʝzD�id��
a|�B�I$|W��H���B��1 b��:X�C�#=�,y�#�Tj{��T�U�n��C�	�y�ƍDO�P���CԪƴBHC�	pE���'`�t�  7�'v�C�!
��Z�R�kA:k�BB��<���$خz^D����!wB�I���*�䁆B��L9E�_�l<>B�ɝ�`|��H��U�4#� \�?2B�Ih����ݎH���z�&X�n# B䉤?7*Ђ�Kϲ�f�A�׸��C�I;k�L,˗͞t�2�pP�Ӫp�B��
kSu��m/�B��D|64C�	8>�8Չ�Dƴ8��8@��!\�B���Z����6�:��ǃ����"O��b�h�)�y*��
�G��	�"O���WbO�m�0
!�R�n��%a�"O&\�4 ̮C\�&@X2X ����"O���Ǆ׼*FD��e�^*��"O �@P#���@Q��B3v���f"OlHp����Gb�2���1Wp �)�"O�U�
׍��e�AQ.bu�a��"O�PeiX$0��첣 �$]ú	�D"Ov��W ��](�coL	"��l90"O<%� H�'
$D�`�0d�Q	Q"O"�R�C�}&�aC��	\�T��"O��:3�vZ�Yd�'g=r�zr"O~Qx�H31
`Qa,R�Z��"O8�
�ɒ2�c�
�.��!��"O���3≶2��A��CV&���C"O~�y��mq�y[�`]�y���"O }�� �VgV CQʏ�R���"O��t*`���^@� ���'�F8(�%&�"����30X��!�T�LB��	��� z,���73�BM*��_�Cy�y�"O����P�IZ����U*h�E�"OH�#�`9|=t	!"�36��X�G"O�@�)�6���a2Gwy�"O�|�Ů��-ب��d ئDd�*�"OD�(v�!w�"!v���b"O�4 @Id?��a�HE|�)z�"Of�xcB��k1�A+��ʬ�j)@ "O.���B�n�H#'&_�n� �"O&}�ۈ>8|�r��)�>�1"O���F�I<�����,�61cV"O�U�&��x���cj�p"��"O" c#U�= Z�J�R8���"O��e^IE<`ԉX�I\� �"O�9k��72t{Gh��OK���!"OP�C��JU�2�)"�=�1"O�4)Q%ޙL,��M��?��5"O5�D����m���Ɉ�r)+�"O�Z�#�19�P�r��1t�`��R"OLرA*�	oКir���+�,�"O8t��/�b�X"�T��(u��"O�P��:�0��-�(U���x�"OAw`͢��Ak#d��Qa�'�h�J�H����d׾L=LD���O�7�4]�w��,!�DؤK�@�	�$$¾�m��7
1O��U혞5	�EF�d醲#�`�uV^xx0p���yB��xĴY2P��+FXaP�� %|B�ѣ,e~��рH���m�t�k�ٰbpD PK�,�bȇ�\�>�xp	G	5�p]��`߂C�����h
�~�h�ה*a|B��� ��F	O	4��h���$X%='�8�X��:0� |�$�iq��B�!���y�ŀ4�P܀WN�Q<hT3�"O���"`VF�6��,0v�I��6Ob�yD��8;��0#�g�6^e���@�?����9آ�z�O����"�fm����nb
�������J=y\2p�s8� ����T�+~V��G%8�\���Ȁ
�F��R焼{X4x�;U��O��jԍ�,q���V�%"u`۰�I^����U�\!x�½�d� o�`����2���"�j�5�*I��x�jY�5�څ����j��D��"�3b�v�ScbJ���:���O�4v���1/����/k�\�ʱf�d�3��ʟM����f�����D`�5��2q�=w����F3D���e!�$=Y>��J�g� H ��]P�3�ҲL��J����B���A��L�+E���ېA�<�y'@Ãpiv�I�"�����3�p<�1$H& ��Z7�J"t��$� �ݎow�jb�
���à̇j����6��-'D<���j[9�H�6��j~�J"D�K�fN�`�B�A�Ԩ��V�m�'�|�qS��4& ��ɖH[�����֘6כ�&��gV��r�ݹ�HMQPj�
n�ժe��9Mơ��/��D@��f=|O<�C�[�m��cN���� e�@"<ҰM�aA�82�8K!��
P'��-���Q͓��5B���&#�M/X[@`���6e�#�'���	�m���\�Ku���n�<`�dT�gq~��B��;SR��ʂ$Jp@k�iTj�b�*��X�Be���O+e���:�EV*t�H:qh�
f���S��Q�q$�ɣi��ԫ�K�*�$,Ő��

Dy�����(�,,�ӡ_-$ڌk�g��w�ڝ�0J��?�a���:ct��C�/��O��U�T�P���.Kj�ib��
���:�%�'��i��#M�����M�'W~�(B�ۆ+Cd�!�
����rR�ӑ�X�٤ I�(��)
{l*9���TN���	�"�!����3N��lAI1Zr̨C��P�,���4I��T�����;'��bI�1K��PiI0_yސ#�;����q�V�s�ֽ���ڥ@2��9��M:P�S�������8(,�yU_G�F���J���i�Τ��+H�UĠ�(��։w^F4�JM�����lK�g`�`W �,{(�� �(c�|��a/P���'�p��k����Q��W��ً�F>G�T%(�ϊ�;"�=������+1酗t``�3�'
v��	�3�JT)��A</����GX��(�r8�4�l7T�;U
�������"I�r-��#<U�*����=/�l��.֐k8N�s%�������JF�8�Ty��@Ȳ$ؾ$���!7?.�Ӄ�T<� �-K3��=��j�6��"6@T)>��!�b��;[��1��g	T�ڳ(�-�h��5�2��=�O�� ��U�3AD a���e�08�@�=,��k
�2oj���
W�A�"H�N3>����F���c!Y6iV|���
/<`���)��:����z@:q%Ə*1��g�1k߶ȘAI���~%���X/�̑2�dE$:�y"Dפf@.q��h�U�-Hhu"��#�d���G�av��8�Ν`�䅊b}X�@�Nдd�
��S
��PC@�P&gT�A�
Uk��DۙA�����x�y(����!��2(��G��Wy��ЪF�9�2 N�� EP�g�<A�a�b��`�F�\R.������S��Xf�τo���0�S�? �"�,Qe�h�i��@Ybd,1�-�'��FV$���&f��ݕ'���ɬ27�(���f�0L��	�9Т;5eA.x5 A�iR�����>����W�)�z ����R�ֈRЏ@�,�ve��+G9��fj]P	���4\ݮ؂a�!I8R�3[��%�D�-k^b�r�2x����ָ<�м�Ĩ���'�֬��HU�j�d�KS�Z3nrv��C�8M�L%��hf��L�V)�
o@@�@�>k�!�Ml���0�����C�A�e��x���
�`� ;�`�d2R�s@H�0���c�3���D�>�`k���6]Tca@Z1`9H,⃠�67���y۴c( P3��K�F\�D�AϏ�>��[#���`tK���D 	ߓ6���,_�H���\��l]R���{�j��%n�")ʭ�a�V�t�L���42�ȍd�Ÿ9���$�ߪ7���X��L�Q:H$[�j@0ZG "5A�y��$@u��� �ʐb�!+i��R�%g@�`�X�
��i�2!�.��d��VEp�۔``yAw�G4/d�0�AĪm�`�Vu'&AS��$ ~�\B�+�(d�ZXkA�d(f�P6��&m ����D�M�h�`u��n$�P��X#j�@�4�[I<��aF�V�(�kE�J��e$��i�(�Ѕ��m�^(����:"�y�i�'mi�U��C��i�Sߵ}��Q�&��(7tJT��>%�]�ǉ�jf�˓z���`�$aډ8�☎f��Pb�T:�`rr&]���>�Ĕ;
��[�"Ԑ0Q���8hEP�3Q`�8"�j5��I��� 4wH��:dC["�L�i�MI)u��`C���8n�>lZ�.ك%��(ӓb2�z�,A�t�X0#�&Z�SP ���42n���t�΁��|��X]<7�͔Q��i@�Q)��h���mm�hQ%��� ���}��L��",��GI1n�81�=ك�6r����5��d�&8��aF�:G�U;�)	?[����S�ï�r�a*B��ꂆ�*?�,�B�LƳ�6���[*-n����D�*}2��مn��'���,�Ҽ�wC�^�xtB�BM+���!n+~6��N�$.д������ڴ�GÈ0(��7�J�c*� "#��kƀ�!��2�O8�2+�	R�fD@��>x#��i2B٭,���(�/�D@(�oZ>>GV��0��7������b���*VO�?#)�9�2ë́/�8�FfS ٰ<afʛP�I�m'C��U��d�3t^�`s�l�*���Ai��wE�4Bǜ�����*p � ��sQ�T$Lɸ){���I���	�{)�(p�O?6m.5H�E*}r��|j�@* j�~
$e���!��&'��X� �s�r|X�K͈.�Z"��"QR�h�ǆ7�ܜa`�.$0a{�c ]�NEԆ�H�
�XCn�
n6\�����Ef>1�do1즅�V��_�LA��RI��xΛ�j=�D�gI�]Zg��7�H"�	��?��ċ6d�&�@��Ŗ!�Hi,1p�Ը��7Ux(rQ�B�.,�ԇNE+�!F�"�81�bQ��x�� @N ,R.��OZH	���

=P�3O�v�H�g����Ԓ��\���G4T�	@aHH�o��e��@�l}R, �BFtuGz�! h*�B�mi���������i�?x1*�xq瀋�T����'q�ӇÃ�?i栝�w��)���R���lڔ�a��k���fٸ����k�^��s�Ўh�:� [ �$ɆI+=���iA�u �E�Kh�Z�Sk�,R0�"^��=�P$`ba]<V�B�!��~�#H�U� ����/�<�夕�]�x ��H�(	v(�R#^ELAQ��2\�4���ƀ(�"9�'V�Tx3��0-`  �����nƿ/�D\#���/ώ�>Y���3RppГҭ��Tb� �b�Y�1���B��\ F��Ik#I�?o``�b�(U��r�OY�5�R��(ax�
%��B��#<�P��::�6��cǄ�ɠ��Yd?��)��F|��@Z�l%�q��̸>�8��q��Ր����|Jb ��I��`ɴ�[;0Qr ��"Ѧ$�T�$��K�����	��$,F�]�p^�]IA�$�
�:Z��tR�Y1��ئ�1c^?��ro�
L�,���8�t%��'ΓBw6��g�-ig�9	�'LJ���לy<��q�\E�5�BB	S��H!!�;*�I84i�(-��9��I�q(���R���ԫ%V@؉�.�;8����P3.4ƈ0��;k{Q�����
�t�	���M�$3���F�R�<��Dy���	�*�6�Q�~(�v��g�ř`�"}��*�P��	�4i�0�&ԫ9N|�de�(d<��	�˦�Ȍ4��paul�ef�8aЮ��Tw��>!4 D����Av`c�����>D��`��0�L��<1��%�cl����$Q�c��%$��{C��8�<�O@�zk,�'�0u� /��aH�.�^I��W�t�R���v°$b�"�50�"|�����Nf$9����1#�a{SɃ�_6VA8��'3(�Sd��{w2�+�d�@z����R=Gp���Ҽ4DL�sT� �>>�kd���G�: j�+U�(5Lu�C ��Т!������4�ъ4���{f`��'�P�H��O�#J��[��E�^�Jp�v�ō�q�:i�V����F8V�A�^_��e"O�EHՌ̇�r ���	9$� ��hS��@Pq�ƀ<^�X��B�j��Op� �R�>	�._�Ab%Ą*�X�+Ճ�\����q�ܵ3�H	��� !�u�-*s�镃M�P=j���6�(	�`0�p<�@&N�T[����]*C�����H�>)#���)t�-9"�T"v��Q]px�ǉ�z��eztCI�o"��CKإp�FQ��
O���R�{@����` `�O��Kp�=�>8���B3Ol�1#�ɚ?&���}bwD%尕�"a�-�t)0��a�<�S.�2[`�#�J����#a�Sg�X�7o�!;�M�F�M�a�(��,ʛ��'��4���o���Fl�R����U}2,+4�ө7��)R4A�3zn���O7!��C�_�B� Kq�G[��5i��� �=��+#9�0�����J��I�m���S��9?"�  	UH`����1&_4u1D(P0�H�PWi�S��k
�'��X��C�s�\��%ҡC ���'�4��t��/�!z ��Er�H�Q��L,�d��0�t�ɣtep=���X}F���
��y���8&���'$��H�2��->FT��\�xEڱ�*��.*��K?�CסT+'Y\�7O��C� ��i"|��ïC�B2���@�'q>D�#O� Аu�S�'6� r�@�d�L�i��X:��A���#d�x6��%ۆY���dG�_�j�듁ͼx��`����)|Q�0�Uo�:���W�N�ir]Ҳ��\��P��䋀v��5f�SZBiK�̔J�X�N�CX�L��*#$�����ːY��H:3�>%�>_������f��Q:��PT�tԃ��.~F,��Oc�e;Q�SRX��K���	����'-�P�}�e�)�X�Z#⎨��m�`��Ă��X��bk���=�"E6���Ѫ�V$��'�+8�����'��!A�!)I�����',9`�q��H�Y�� ��^�|��L�B�G��� �ŏϢ.F�ۏ��#g�d�u��5A���4��`�џ �!�G�89V�/4�e(X!�E���%���8�˭0rbɊ�����L��K(�O���A�^�=�`�Y���1��(��Z�أ��Q *�ؔ:S�¨.dd���ξ_`�rKM+7�4�S�Pg�L9��ˍ0#*�M��m�B�	9��5x�a�cЅ�ue����k�� A<�����\_Z9���8����r�������;�֭j�qY�56�( ��}���dD�/��`�B8$N�Y�&��%a�8��P��'��R�Z�m|qJ,��
���1�*ʓl�H�-	?������#	���G�ǜ5'����^0%�6����Vq��K�9L�颵��Oo`"e�9A����$]��p>y��F�e�D���8����l�yy�eS ���
�O�1P�1���k^ 5��	ϩv��=S�O�e�� �
�F����F��ݒ�'�����W��u�)���sf`n��1 F*E޶����my�c��~�������;�w�BP��'��@w� ���J�mBZx*�'�D@��ᆁ9��:gȦG�j����Rj8��
-p0�|Z�)�+���F >ў�Iԣ��d-^�3����(� 2n'O��Xa�E�6�4bH�e���� 4f��s�3$���d׭PCF��=�0?	�Iҁ*e�T��ʈ�2�!��R�	�.f tcV*ώ$b:�	%;��p9S ;��-[m
r�������$ EIʏ�y���!!�v�`���±WR����D�!��'��(f��>����v�"Q���ӡq���F�<��Ӽyh�\[��P�I�0�̇C�<a��=)F���n��)w�m�oF{�<Y6hB. �j��6Kݻ]08��Fp�<1�B�($����#	z�1��G�J�<�e�=~(K̶I���!��inB�!#�T`���.@��$m\-JC�I�A����D�rzi	� �8K%8C䉦Ѥ4�δU��.��B�ɩ-�-�W
�*&|@ 4	�3e�B�ɷD�D��A
a{FlKC�B��B�ɔ7�<����S��5*���OS�B�	w�2���m7�ȩk�$�9j,�B䉗z��d�BD�gE�C��c�C�	n�РBa*NA�&(ҧhSK��B䉧Q8H壛�:}.D�_�d.�B�	S��!����,p�<��	�%ŤB�	 ��]�r��:���wd�l�HB�ɖ�0C���/_��"�C$w�C�I'F���5$�.i�|��e��o"B�	�,tP=�u��3>��0h���C�I��a؅	@~	��@���,��C�I?x�{0��Α�'E�'J�C�I�����C� �v�/�Z�"O���&ơY+ -p���o.��"O�Z���9#���%:-f�Jr"O*M:c'�������dvI�'�'�y�`
X����������`Y�#ɐ�y� $]�P1$��Z"�A�A$�y�W��ñ�6�J��R˙�H�~B�I/KXzph��9,���
A9ZB�)� ��QҫO&]ȼ����1���1"O�$)�!єFH=r����E��UR�'�;5	�Z%ft�q�C�F��	J�'��YRӏ�>S�\��q��-8��M��'}©�����(#��.+�"LX�'xRm�&�Q+S@�p��>p�p���'�ލ�+ֲv�&x�g'	�#�fMj�'�~|��l�#�Ɲ�&�Ű%+�M:	�'/>壒�3Y�F}EfG�7P��'_�R��W�]�҄�t�Q�PU,��ʓDv�3�����tr�ǂ�%����d���z`�N�~l�=Z�C�!0؇�oq@��U�V�)�ĠY�#� V`n�ȓGT����&�70�*�ҮX�U�vĄȓLt ��Ӈ��&����"MZ/X�D��ȓh�庡fB_�.źKǀQ�P]��G@���84��A���_o�l��{��a�@�15�6��gfW����ȓb���*il�x'��n8�t�ȓ{G��*Q� 0y��]�c�ő@ �U��_<@ht�R�S�(��t$՚���f/*TJ����Y Q��{T؄��*OJ%!r Vf�zɓ���&D���I�@e!5/��8���.��C䉣>����dH:,���{V��9J�C�I8����;�ޑ�6�M�M�LB䉸�$�kݟoՔ	�-ʺbA^���5d �L��^�X#Ƅ�$c�\c�Ƙ=ϐ��0o?D�xȦ�¡d
�mp��\�6p`
<�)]�>P j\��ȟ�(�GHWx���bI�He�y!""O�{fޡ��H��'��-b00��M�dS�Z�O�l@d*/�3}�e��2�)`"\�,�9�B� ��x� ěoڔ�;F�_;�q�I�_�t��֭	:`���(�O���A�Q���	�C��/D���U��
wf�t���S�$��ʗ91	b�;e��2]Ӻ$�ӈip�u���D��.D���J"�B�ɫB(&��D��/[�C��گ���I4풥m�1B��Z���)A- ��'o�1�0m�YV�i��8��}�g%	s�rdӴoQF�~�"�OH�#t�Ǵ_��iǈU�F�j�[�Ċ�Ghl�%�]v�R�Yj��B��$��u�=�	�Ll)��	sH0B��&�">�sC.~�P�΂D���!��=32��-��S�D�FFнI���{�i	?ۤ|A%�E�dc͋�6Zlq�O�9F����cA3Qn�H���f�8�#4��=9,3�&�1JH9oһC��͓�À�Ui�X��;`,���B�,��4�Y�;�д���p�@M(�T�P.<C���9 oǠB��"�ġ�*�4	��|\w�^�k���;�q�w7��Ly3��"� jv�ܿo�X�C��'��D�"�Yr��aC��͕=_�8��
���!n�tZZ�*���M��9��ܟ���+�n��1�%R�8HnOI��y"`٢�жJ��yR�N�E����'�X+�$Ɯl�@kq�ĭ_�l=��!73I���Q+g$������+�:#*
5m^x�ѯH�5���
��2t��\a��%|O
83RFɅe�D��3�Ǻez"���k 2 c�D`V)�9;N`�;�'��K�k��b�Z�ϓbv>ţ�����ׄ*�)f�C�sy(���'��=35�ŋ'� ��$f�zh��fO?XaڹhB�Mn� 8l���o��N�z�!��hW-�x�ШC�dڡF"�����y�L��Eo��G}2B���J�ا�U�eS��a�I>C/��#�͔&�!C�ϑ�
��Ua�!M�8�pa��аA����럗C�ӓ��%�GxR��&,l˂�d�,�#���~r�w �k��E

b	s��݋�Y)7 �0G�D�����1e�ҹ�AF�N0ْ�@�)t��p��,m��D�S,:R���$G��`���r+�\���ӠGlp�R�3C��}��AU�m�2j䀆�-�� ���	H!�j���`�&�E#P����l0q�&�'^���)
��؂E뎷�LU�_{��n�^T�d�i�؄S!�$f��S2��]�vቆ.L�Pd���	; vM�E!X�,�X��D˨WI䨂������O�%���MF��e�O������� +��p ��N7j��4�B%!���P�Oǟ���ǘL8xB�iX���DX��W9J<�O��R���ٰ`b֠X� ����T?!RF���r��YyB���U�@�%�rdH�.R�M��K�[4����,2ೣ᏷�@5sC戱F����@B�8�p��	�
 LI�F�E$P��\�f�R��bU7i@pb���7#m��!a�/R}��a$}R��	��s��|c�����<@l�-�Ū�S������' e+ kA^7�,(��	3`�2�IҶ���EcM�c��l�,_�8A���� �v�1��\�i���R&hr� 2]an�z��*���5:_��Z����q�8��$��f��rO����xŅb�,�s�IrP�Q�݉SXxƈ�C��ѧA�
ġ@�eĄd�6�T��X��@H�w����剔��-Cp�Ȉ9�x�S�ǻ}y1�� Ξ��+O���G,��e'^�������,1�옜|�%0��/��$�Y������ 
r� ��1j��(���2��8�����L<����<��0O|q����� W�vQ� �[YJ]"���c<�5��!C1��k����M)�gi��&p6�q�cؿ=���I $�*e �4L`�PF���-��qtD�&�����&�f���kի��?01(�Ē�!B(dx4�	/{���T�I�N/�4� �5�L�:��K�<yg-A�y���X�J��c�`���ғp��7h�b���PF@��	�"1�bҸr�d�St-;+��U �AI���d5V뼰��a��#@lؤ���]�a35.K*~H(ڴ�ة�$�D8����/]�z�j�OmP�a�#o��9��� ,��'��&�a�gc����;��!yr �Pb.�%{?fx{��N���ώ�B�=�$OkD�w� �� &�<vf��0 �&a�p)���,���8Q�dqCT�RW(*0rᯖ�N+��S���a
|�Q�]+_��B�	I������$�ڵ"��C��r��&�E� 4��$Ʌa�'�v��a�ړ� <�D�R���� hD0�"�p�� Z��g����Q�E0g"msGi�!%z� ��ݝZGz�o|;�Er����r�wh	���U/iTJ��""��CW΅}�F���eayR�]8=��ȡ��	�"T8Q�#^�,�5�P�p��p�'����S*mg�[`&�Ij�(%.^�;�ā�Ƒ:m�\�Ė���M�t�,ْ)����C>�`a�D<}Ip� �F��")�(@7�Za���`\R�3��΁I�&���O|�޴q(n�1���$8�ebՌP̮�R���yX�O]�-�L8Z�����Nr�����dεx�� ��[3I�b��:��|���M�ov�����=	���&���p���	�l��PIݮd�m���6S�v�Љ��$s.I��Jk�|I2нr@�P�`B�&Zh)�$f�#��S���%p
"	r%W!Nb�X�/�?wK�X� ΢R��@a�@1WocdM�@�8
��9�O6d࡮Q4��SԀ՝�E�U�҅�u�!�1EZٱ�`\7]�>}��Α4����8���K&>�%�ߡJ��E�À�'6���D�UX����2Lk�ūuh�)8��s��/��|"b8AO�MaЫЪ"g�����O%U->�#�$����[���Lz���9CL�Y�O���d�Zg�q�Ei��|I�>��̊!�聱�[�^q�q̐��܌@�_,oV�EI�**���`d�?'�M�e 	�_v��2 (B��Sbh�߰=��bΣ[&�=r�L�9Y�-�Y�$](����3�㍞+ք�(G&�u�:1��g0�����	tk6q��YW�a�3���]9��zbe��n���D[Q��4�
�<,�u��:#h�*&0Ow������ZJ��K�"*$o�<�����&�?�B�ɃkF� 1�|�#bm�W�' �!U��q8n�Y�lI6rP���T
Z�
h�FΜxb��낒M�V��%/�5m��ŰW`�>���.{
�#=���F�<�RG�� c����py��˜F����F�d�dy9�AP�@��)��	�l���	F����Ų�lS-`��#֯Y�Fx�kA�it�q�uL��{��|�	4U`2@Ƞ�χ!�T��)]Ά|+ՆB
��@h�I��(���l�5Wb��#�`��➫�y7$F�C��-
a��&6�Q[�ʉ��p?yR�C!�H-M��y��-�帩���L��Ȓ�	�4�t,ː���/��!�4���J��M��b�ڀI��|�G̤`V����K��d�a�4�9�p~�PJƥ9�*"�@�K�YJGgM�!�1fΟ�I��xi4�ՍoN$�	�M�2a��U����<ٖ$%�K��>�Mc8t���[)`M��Хb�h�A�$����3	�0!�d��%4(�A4j,�(� �0�k>��A�X$\4����~X���bE�O�A�5�� <�����0餪-k�΍�Ԩ��8#0Y�K����f��O��}"���V�}�@xR�oR��y7��y����E OdZ��3j�p?	 �vO������"��4NҸ<1
�XD�p��"�J�>��C@Q#q|�U�7��DN�F��U�Ń)_�HX�a�-Jb�#)P�FePp��Ċ�&��JPė==�	����ձ���2=���a
�z���E�D�81ӣ�)���O�}B懳Q;H�<� ۺV�nQS�� c�����h�g?16�Ho$���̞B� �p`��g���	a���;L$�I�"ۤ`��5�"*F�Jz!��p�*\ w��
�H�5J��f>��x�N�u�����Y�� 6�~R����u:��4�O�]˪ Gɧvٰ]��	�m�F��P&G�f\Bmh��xYp�1&eR�Hd�3�!�6|�g�V�gU*e�Ǔ$�d�r֠�7 R��k ��V�|D}�+�/d
�]K��< }�墑�"�v�zdMCu�%3d��48��4#_�D��B�I�>68urf�y.DX�`�'��2���KQ�êp(��D@����)qC��=��O�:�t��Be�Ч�ϙ_����'(Ը$'%*x�H���O��z��3"�L}�m�R�I�{������ָ��'�|�1O��Ĉ3%��ݑ;x���h,�O�(:s��'���8$�7 ΐhf鋖^np�
!��E���	� �
a��Lх��j8��a��f�-Vk"������O��s��86/:�Eƃ�V!��� �Ѝ9B��-L���\�!B�M��(股q(<�uNӻ\c����)��|y*GȗW?	���Ij��p+��E���BW	-4T���4�� �)��ċ7�Y��M�bTؓ�"O�tӤ���	�'�G0,�k�%��J%���w��2Cz�Hb�9QP�'`��� ��>)����3vT�u�S+5l D̜S���D��N�R�L?4����K� �^l��,A�"��;��[��$@M��p<q7���:��H�u�ˮN�`�
\f�'�P����ʗXX�В4��5w��I:�m�
{(q��G�̢,[!+"4�,���2��"�V;wg���D��C�:x�3����3씦�V �&!�Fjt �«\�0�FE2�Ʉ���	5Z!y�j;�R�.@�)l�B�	'J��t
tݛx L"0�@ N=�D��L$E.���` � �4�-�4��J0,`	��<�e!��&��|	C�!m
������H����ab��x>��J�6����*�Bn�bqNRg�64�))���� �)�(�P*#�	t���	�by��B�Hr	G}�@�[H�dx&���>��dV�
h��˖�;2�3bl�s�
��WlJ�|�bU���"�a}�͎D$����5>�l�s��=����2�����
p��jwF ��XC��[�o>�!�৾?�`�gƘM|6�37m�7s8���#,D�LRL�"���QՈ��K� �cF��R��Mx"�ϝP��4�4JP�eîXJ�?Y1	U"}��A�;{����
��r�j	a��JJ�����	y�����Ӊ<�
�s��7sZ8gF _<���	ѹA,�m��uk�5��
;��<y%I�0 �dA����=I2X���'�e�'����
 |�:���@uj׬�#c���х۴�Ҕڣh��� J�nP�Z�]�	�K��YX�M�'i����j�1�x͕'��R�l(y�D���&�D��["!�:���&���"��By�D92�_�^�����y����� M-65��Ғb��t�����,�5�DR+<,5i�-�D��)E'%Ybt"�<�B(K��^ ��i�N��Iq��'�J0ss"	86On�2�(јSs�; ��"E���Ss�W�4��a�A>�:�JH�1@p�Z�򄎒]��9���	.e� ��nK�<cџ�;��K^+��Rd_9)���3DV<.��.�F��6/�S&��#+�򈚶fE�l�`�����V��EK���ie��b�M��rU剂!�����ܵI�}�A�/{��0��B�j��i���?ѳ�L]A�x9G��g��Qs�D,D�la��!�t��%��P4Ĕ	���~!���6X�iUC��'�`	I?A�TJF�6H��;k���K䌔�	�`lǈ!~���j���â�·`����c�	;y&\-I���,H�l V�<"���'B���@��$�hO���
3H�l���D��[��'�v0��!��Jq�R/hk����Yh(��S�C+��@��
:ɘ5��BN^��X�bEZ%���ѠxRa���:�d�#@����oO�*P�đ�os���~���E�VC�(Xh�?�>�ӄ��T�<i�Ȍ�>�<�(�L?��A���R�����K<�&�K�����ɔl7�(B!��1����`X���"Ox�(0F���f��Ə�V'���"O�y���K�^�슱`Ҽ	8t��"O���%�1W��hK�"�26Y��"O�d u���t���(p�
Np	�"Of����.K�2��t�֗r��p�"O��xw�@6{�&���	&v��A "O M3Se�${��S�I����۳"O&��f��wVh�J#�<���C�"O�Q�q���P�#�
wv)�w"O>�1��+����@�pTp�Q"O$܉�eO��i��ϻ[A\�1
�'�����n[�#y�T�R���q�L�"
�'Ą �h
>��A��=0���
�'��S��\
WN�#�HM?)�
�'����s��,fXd�'���}M�XY
�'��Pk���t�����wBt��	�'���H�cOlJH�&%?'�K	�'j!i�EŔ*�B�x&��5�6"O�8�A�R0�N���ꅿ ]�!#�"O��3���N�6�UH�J��=��"OT����P/]���\����"O�0��G�$�͈c�?I�P��e"O�ph�cF�D#c�K	p��"O4�q�N�m��Da!%��+�DZ"O�(��ӺU��Ic�d�|Ҁ�C0"O���'	�'z��[ǝF�>�B"O� xX���W���'��Y�F�3"O@���H��Ѳ�B�V�\��"O�%날ˀ,���V@��+�
���"O �Zq�DH�}�����3p"O�(C�ՔgCR��pc�yĢ���"ON@�g5J
BH��(�J�P,"Q"Oȴ�1hF�n�ԅ0�A�!?�����'ِX��FFt��Q�	���ƋFRq�'�ܬ����D'�5`��J�P�
�'E�L���X#6��<�� B ��d�	�'��m�e \�.% �;`kr�^l�'SZ��ǈĚ}Wj��'fKo%���'x*�
`����t�jW�6'�t��'(Pr��� f6L��a��,������=�Q?l03v���`�f�2��d� O`�`:��G '�a��A��s�����S�O&�������	'l�N0���~�O�<��n͉�4K+hj�9>OԘX�lSp�S�O'�03�!���2��Q��.5|.p�'���W'2D�;�
�����'��y��O1H4#�f�	D1hp��`�*�y�ک)��}ӆ��b�G�N�y� Z< Vq�dL,ZN�9��Ə�y2�G� � ���[�V����c���y"����9�4-פA��ѣX	�y,��!��xT�� bu����mR�y�I���G�&������	�y�
�!k8���@�]�d
�P6�y��Z�48+�C@}���cG ӳ�y�/9c>��b"�t���[��C��y2+Ɲi����0�W�=.I2)���yBL+"T x�奅!*���֏O��y��o��Z��݀Ed$�7-�#�yBȟ�Y���{�k�c�H'NP(�y 2}2���n�ȇ���y2J�-��-HD��k�N��w���yR���s�t@�gETkr�XPH� �y���(�r�V��_���qW���y�́R_�TZ�#��R]PS��G>�y��� X<��3".�A��u/d�PQ
�'��<zG
�6��s`R/;-8�q�'Mx!Cu��5f�s�5̨a��'���
��_>r$�Ӯӻ1*�|�'�^D`w��j����*�TM��'�������_��ӌ ]�-��'+�t��M�=_&�cv��/qؠ�'i���5�ɉiR-Z��A�Z-�h��'}���p"D�r-�E��J%A0	��'i�py�B��Q�L���G�N��٢	�'n��Cc
ى6ef����?f�E��'�&��uaW6U��q��^6 �`	�';��+b��1�ꨪ@�y.�@��'͐T8��M�
=�W�w�T��
�'�|ȂK�7Z����g�+~1�б
�'�5��#��^�$�A�m�1��'Z-q&�U��z#��V�2I�' ��C�p�&�؅Qad�I�'��r�O;F�P	U����)S�'s8���q��i�aί+�(a�',xX���,z�f<�R-0,�J��'�D�qd��R-;�(@)5}��{�'h�\�"�6v�����C�,�Z+�'k 9ٓgJ<������84�8A�'���Ћ
3pkl]�5#��&[��j�'�x}@��Z(u�<:���&��u���� �a{�A��4�B�y�*B?L�,�7"O,	��*�	�	��G ~j���"O|�&�%�~��2\zҘ(v"O�(�
v����(w���"O��I�U�,�&n��<u� �"ON��s��8N��[Ŭ��Vq�"ON�#ӂE��V9�T�R3^�2əE"O�� 2�F�$�ޥQ ,>J�����"O�1@Tϑ�BU;p`K��lH�"OL�����8S�}����?0���s"OFXq1��.=-z��'m	@�@�)�"O�8r��(ZZuAT�G�<�6Ţ�"O��r�	4��81����l:�"O� xQ��_�XD���ܰ5����"O~�I@!@)��%�CG�b� �!C"O*�p�������aďU/ۜ�PR"O�u���( ���e� �*]K�"O�]*�&��N9��CeȾUb��ѕ"O:�'�䐁@�Q4T̐!1"O�UB�Aݝ~ˢ�;Ռ*g��2�"O��(R��/{�@��eʰ:�(�4"OB��V�H07����(5�N���"O�E25��8d ���Gl|�"O/Q�8�c&�)褈b#W�[�!���r�4#�!X��x<�r��4&�!�D�&ja��JH"��X��n�b�!�DI�4}[��6'�~�YU����!��dTIR���!l�*�rF-�aw!�ę-Hۆ��ШN	<occJ`@!�ĬU�`��P��5[�4�C��0!���0&
ڬc�OQi¶����U�!��m�V4W
�2�����S!�V�6��
�e������Qm�g"!�D�u	�K4�x���j͎� �!�#�(9ǠF�'Y�%P�Ό�!�dƼMk���RHy?4l��)z!�D��i(� �2�8��D�!�DX�Vl<1����/Z�#GPh!򄄨\����qfМN�4¶��'ўb?�ֈK�L���A��Ž/4�(˄c2D�4[q�ԑA�����!D6�ph)�$D�4t.��m8��0C�6)�,̱#m$D�(9FW;uA8��&{��p���'D� GB	{��+���.L_j8'D!D�X "J�S��` ����T����)D����,�:NU"�ZQD��`�����3D�lp5J�>#�����nq\C2D�Zb�ϔHg�H��*Թ4D�p3/0D��q,{2�"q�V�c��eT�#D����J��a��9�5���'wEQu�6D��!р�$O��"�*�?|���$"D�xb��۷t�9iF�A���2vA D�ȣ�� & �&��"�T%��!b�<D�P��逜"|@��S��H����G%<D�Xz/��\3!Ba���,D�T���nM���P��Z���#i%D�Px�N�7PP|����aT�1r.%D�����٩Y^5��`ʠH(Љ�c�.D���W�8`�r][TS�Ya�5c&)D�P;�IX�PX\�Z A�B:���)"D�$9�* �6u|���F��u�qR�/ D���c*�C��D�q��=���j��<D�Xjc�.�$��s�� [�t�2c>D�����ú6��ء�Ѧq����">D�� Jp9�F�]3r���C!=G�E�"O�����W�R�$u(�L�`�iq"O�%S���� �x`�ڄ��e1�"O���u �L�x�1�O�q��"O��:��� CW"��e��cд�"OLx�G�ՂSg^ydȞ�1�>5��"O����$$Nž-���||4��"O�Y��ϲ+u�)`6�j���w"O�)!�&�f�*��
.{�T-��"Oȍ��Ia����'E[��@�6"Oĸ���T�A���H]R������y�	��m��H7�F�)/�Mr���%�yb蓬u�N�Kbb,����yr N6����$�׌1��Y$cT��yr�R��M�LF�w�ty�C��y� ʄ'�:���kc-sM�0�yB���b�"X�%�V-�y��˛�y��P�pnF�+S�2fG� J!	�2�ybN�ow\����f
�Պ�爇�y"lֲ;���f�U��90LP��y��:?��Q��J�J�F��	�yb*��`d��g��N
]�#���y�U�2�F�:e�]	wf ��C�.�yb�ڔX��X��B�o���{q�[�ybL˫b��BC��&c:� Ѐ7�yr�3I<by(rj�V��{BO�y	�]��C�_J�8����_��y2�A
ePua�Ǝ=���'H��y2hJ���b�H�bK^��p�T��yb�
� z9��(ȱs��S�)Ҍ�y�	�R6XL� ����RX	�K�*�yB*�wN-q��֫�zd�J֣�y"��h�X���*֣���q���y�Fد��8k�IV.��D��"�y2�ݖ3��ZՈ�$xM�ઊ/�y2-	xl�b�G�rc�����y�䝰87m7h+FS�.˦q6!�dҼL���w��vD�� �&C!�٩cH��[�I+y�>l��n�?!�DK�f��L�ã]�D�<�)U�Y 2!��[-PRhR�B��VvM��J�T�!��ӽ(�-���W�!E&dr�$��!�ºuW ���I-r��&ڿEk!�R�F3 �� �8 ��SLСj!�M�i�r]�P�Kj̴0uK�[�!�dP+A���C�_&K>Y`4)ʩ�!�;]g�q*��[$6B��pÈX�!�X+�^�*WcI�IV�A�b⏔?�!�$�M (�쏚@@J�ga�?�!򄛷k��괆��l+
�h��}x!�D�2�d�eB�p��5�bn�9Qq!��CW�|`V�ah�#�+]z]!�k4Щ�ϐ�U��b�<2K!�Ė�Ax�d
�T�&Lp��ܩb!��K�4�#��4�y)��<1!�P�51~�9@չL���I#�!���ek���ċ�N�d�X5��2�!��?G�6!�-ы`����D��-b!�䋱N�����/�>�p����ɧeP!��$'UpX9�i�E�D�Z!&F�O!�N͞�1��.:�Z�R`eſJ�!�Ē�J ���0C�6иA+�i�7�!�V>�H1��ܖZۀ������?�!�4��,:���:vŮiDh�[�!�� T���N�N����3^91"O�@a���Ztb�G�K=~FY!�"O��b��A�7���@$Ö�3�V|C�"O�i����	KD��raB*� \��"O�ВD�&غPɥ	
*}�5�"O���@H̳*|��j�<X�`�"Ob(��,��l̹�ȉ��$!�r"OBDہE�5SĴ�P��f��tj�"O��DK�n~֌��+���R䋦"O|k����<�1e������v"O@��bX�g��U*��
QҒb&"O�tXE�@�qй镤��K"J���"O��q�fI15���0wD�N�V��P"OÇ�B��a���~���s"OX0+C�WF�JCش^���E"OTHDi�,OXY2�ƒ&i��	�"O��%���ll� �\�U��J�"O���ӊݯC/z��e��c���K&"O��Yg��7<;J$�a߸I��D��"Or�{��Y�`�ND� �Z��pw"O��xA�C@גD��>q�l�PT"O�\3d�V�'���V#�qq�x�T"O�d�M�#(�Э���G�g�~���"O�p�«�1bnܬ"Ҩs�8�Z@"ODLH7�U�5@b �ë�*,t"OPX�`�̥~��y@� ,��"O�ȱ�K
&���Eiu�q�"O��"��ہYWD�"i�!V���"OZP�2�&9�A�\:1�\q"O��R��/���3		�a�f!��"O�t�BD�o�B4!GȞ�#�6|R�"O�z���V+�؆l��|��"O4�����5t�l�]2�LP�#ۀ�y2�ÏYF�ZGEL.L�4��*���y��^37�H��b��F�26�A�w�!�	Dt�SԈ��A�����څ1!�d��� �  ��   �  �  +  �  ,  �6   ?  fJ  RS  �Y  �_  7f  {l  �r  �x  A  ��  ŋ  �  J�  ��  Ҥ  �  Z�  ��  �  ��  ��  ��  >�  ��  ��  _ � � 	 M �  Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�� |d��"O
`�(�;���8���-0��1%"Oj4��ND^[��"3/9�0|H�"OB���H��*�ʞRy=a"O�味V�!X��!&F�:J�$���"O,��a
���C�Ą�M�"O,$3%o�-���p���+Ն�:1"O��ݢ1����`���y14]2��i�<�6��{_���c�H�`�fX�$Kn�<��A̼VI�xR[�)�Ć�pඤ�ȓA5��('nߡ4�� �)˩%� ���,��r�؊b#`T�eT09���ȓ!�b��g��}�8�F��-? �ȓ
K|m�ș�VṔ���2�%�ȓ"R�X�j�4JN�1�˘X�i����̹	_�jZ��1!g��zܶ��ȓgil,*�J�
j�Ne��i�J%b���f	�(U��:���G��$Y^م�~r�� S�%T"���k\�jx�ȓ|4�1�îJb��@ӵ�ݩn�V��/[`�"�v4�R�!ʎ<��M�ȓ`:��z�ؚh�J�Z��$HY:	��H��p�m�C1��!��B:��0��EnjZA V;9����J[
2���	��4'J�EA�IVW&��~�(aZ��ӹ�>� o�Y�|�ȓ�f�A�
Ο7�H��M�$�����mޠP����/���ANXo*�ȓTv�����{ ��-7�*h��I��sB�8�8���3����ȓNe*M�悡;������X�o��!�ȓ'lj�#F�m�+R&;�|��2)n�C��0S4���T:
b���:�0!��e֊��)��ͷV��,�ȓ0�&�8#���� ع�L�����;�P�AFd���,w�6d��r�EQ�( �gVlɦ�M,H��,DP���|�I	$G#\���ȓ"�)���E�B	yt&B�^�LɅ�4�� ��eëF�ڙ��n��R�p�ȓp`@}bŇ�=�$�AUN��P����L��p���_�a�)�Y�!��-��u�5���o}�`iF�@A�p ��F�\�0��[���IF/5���k>bTؖ�;K'DT`�^��@��fnV���Y�b�lI��	����ȓ,nٛ��Ć3���kC��8�m�ȓ'� I ���x<=���޳{��	��6��(� N�����
�y2<��ȓx;6q��I�
=  yG�O�,�!���Mӥ��B�X��E�P�+� �q��O�<A�n�u;��a�ወT�ި�.�M�<ѣ��"�By�D���Y��LR�<Y`哨YFeٵ�ؕ6����t%Uy�	M���O���:4%]�q�L�R�)��@�L9��'cNX�� �6$oxA(��ژ,�P��{R�'ŀ0���@��9B�M\�sp:-��'Ox���Hؑ� �HԂ���V�[�@4D�8y�2I�~�A�(�}�j�)Qc'ғ�p<�S�/� �;�,�G"��*!�]M�<9��B�-�C
�ST�m��MЦՇx�
p����1"8!�6�G��)��S�?  9�רW w�DU	'� 9�
�"O�e(��h����Tψl�V(��"Op1�aB�ʠ$��I(H�J��p"Ov � c��r��'�A�^����'ў"~��A�6>���Y�  �Q����y¨'�4��ڴ/���p&\"�yRd�I�b����,Y>����2�yb|��
����%�E��J �y�U5�z1���������A]�E�X�l�w�S��y��g�TԨ���*b�L����yB��i?fݻ4U�w�DD�T3�y��ձg�PQ⇪V��|��.�'�0=Y��Z�I�@j2BؠUbx�c��y�D�6��5։�O�tPN�p<ي����R�0�
�s�z0I!�͚�!���l��` 0�N;k��%�&��+��x�Q��$��Cal!D��]���K�~2�)D��q��M�j�)P� �+!d��w��<i٤���"}��R�O-aak�K���X#�z�������I/ ���b��/=j%*/O�O��'܂E���k�.B*n���y"`&�S�'_��A��[a�q���3FQ@%����u}VPC��cؠ��U�W;N��B��9g�`���dU:m�rxy����x�B�I�"�1#�`3��C��1i}
��'sD�JN�k�`Y�l
*L��'C�a��G�{�0M�G�ҋ|L���'��p1���5i�
�}�r��'��k� '1\q"g�*B:z��'	:��/������.<3�8��'��d����iVy���;"|8p�'��l���9���K�#_|KcC�2�y2�y��� �׷�RPB��&�p<Q��DM4 �t�j!a��v�5Q�h\B��'U�#=�}�#��
�ƹ�RD����@���h�<ᄌ!<�9eК\t�Ӑf�k�<�r'M�C����w�+ 7
�#wd^�<�H��W�Jd�f�T�pO�D���0��x���Tm�Ր���˔Y8 �)�y"��TzꭒFҹf�"��D�^�yP�7ϊ���Ǝ�p5��B���y���ƥ�S�&7��S-�'�yB�Al���R��&_��)��],�y,˫�1[`��0 %�}�GJ��x���2�4O��wT p2s�.7�!�$�;�~�9"E-#�i�5�E �az��dDXS=Sǯ�3t�ɖǔ�!�=~�H��%����Ҡ�V�!�F�3"��)��WS��`�T���`�!��No_������19C��`�!򄍋�z�'	35�@�v�νf�!��###r�Ѐ�ֱV{t���@J=<�!���*��(qŎ�(q�:P�C�x!��R�7�Hy�P�Q"gǪ�``��|@!�G�\<r@�U����P��KT'!�H�Y�\!1�a�4D�ty:t���!����(�x�A"N�
�4�"B�X!^�!��r0	@B	;��q�2d@�d!��@�$�6�q"���QI�&$�83P!�$ѱ��`�����x+����azB��U��5��=D�+��B�!�$2��V��0%bN�b�N��'ў�>�bF88���䩞� 2�[�4lOx�Tk`k�r`$0R�A�Kg��h���=� ȹ�&���J��Ӕu�T�A�'��$	jni)a��e���#Y,1!�	F�a�̍�����L�=f�F�H`�'��>��{����A�*j�"��t)K�a}�xң#?��᪃�BA��0�l�"�~r�i{�}&I�@0�/S�>�vdqSGF<������]^�	"GbT܋�%V�����̝}�xB�I8Jn�����o^���˱X� #=aǓa��0����l�ŀ��to����I�<	�ɓi�>D�F �d!�-y@`��<�O���'/ɧħ4�����R��Ap4m	L�*q��N_����!�}��(�%�N��
i��hO�>YH��B(�>XRR@+F2 `'�3��XܴC�@�jV�Ӣc�ٻ��`���f����Iɑ7���Ĕ�*�DdG�'�?�KF�޻D0 � l[�$��	x��6D����ș�Y����eցvG�qі�9��j����rp�b�B��1��h�ʙ�V�`C��~�<����M�ScJ�!g��d"̱�g"Ou끊�+`����ą@�("�TP��O�=E�4F��'~8 ���W��"I��y \�\O9P7(3c��$�ɚ��ē�HO�c?�� )L>5z��W��E�WD.�h��A�a���G�o
�(fg�C3�#<�ϓg=	4�yo���ր/ke���fn��;��Cb��E&��R��q��'����CTX� S�EK�M����'�ў�}b�B̞Dp�uiK�Ӻ�	6��~?1��'��x��'�VS���IZx���'�n-�Ĥ� i޹	�T{w,)��'�֘X�h�$7�\�cD$y��=��'K�,��e�8OŨ�1�M�k��Y2	�'��n�m_��卟]��Qi�'S0�E-��I�0`�I´Z.8)	�'� �$�R�T�:h�$�?VY�aY�'o��S�E�0�������/B����'O
�qfFK��4��'pҐ��'�q2��I���	$GHc��)�
�'`��xI��.8J#�̉	�1��'��a"u
pe
�U�'ТH	5d	�U���s�����\X�'V؀�s S
Y� �bM[*yѨ��
�'0�1
	n` 9�1 ���@H
�'W�)P�8���X��3h�	�	�'�^����O��z0��	&f�E��'s�a��\�>��qplF��0 i�' n����=�nYs�1��p��'��h�1Ɂ�q��qr���*,�1�'ߤ͐do$qs�"g˓;3�r�'ؽs�1: a��I��=�	�'\4%c"À�4�`s�H�x�k	�'�$"Q�*,ΦQ��֫�@�s�'r��P��)'D�A�������''H����7�<���J�F����'�˳��y$p���N�/7��\��'D�`���$W��4���\���
�'��3��?=zL��6
�J�fE��'�� W�Jm�F �&�@R�	�'Wʩ�
�"u�� 6��&is��r�'��
WkO22�!���7G���'w�8�'゙�`1�fҪm���'%�H��R�4L��xPE���AS�'Bţ�C� �(1�f�� ir|��'ˤ�)���-t��6��}'�� ��� �]3�Gm"�ī���[�du��"ONy`��M�W�H�J�bۨ[�`"�"O�|KĤ�df���R ���Uh!"O�!���BHF����.H	�"Oޥ��k�oBd�TO�f(:����'�R�'�"�'�R�'"�'2�'�����!+�Ԝ��	Ħ�����'+2�'���'�b�'�b�'f��'*ě椊.Zzj���!�C�X�{ �'@��'R�'���'	��'���'F����(}�p�a��=�����'�R�'0�'�b�'P��'��'�t�K��ăb�����ٗ	�N	W�'�r�'d��'���'��'���'�ȹ�̊��P���� `w��a��'���',"�'~��'��'}2�'������|�n-"��F�G���v�'0��'�"�'pR�'���'M��'>` 0��<a5���`�J�/x��Y�'���'��'g�'#�'r��'�Z�SnV���uᒂ�/�fա&�'2�'���'u��'8��'���'�8��m�;��"��F����K�'�b�'��'��'���'���'��$q���+}��Q"���r��b�'d��'I��'��'�B�'���'jȨ��E�xm�%[1�D$�'���'���'E��'�B�'���'�`�R�زOG��MW���x��'$��'�R�'�'�BfwӠ�$�O����I2*��'��BN����Ay��'�)�3?ɑ�i�D�paֆ<
|V�T1Z��8�I������䦡��g�i>��Ȧ)�G�PM���
�c[��჋��M��~���a޴���&)[�2T��0��S�N�I��c�(T���#�L�tV�b����Xy2��D�>��"�*���PC#B�B!�ɒ�4.=�L�<i����~���w02�Ӏ)R�1�HS̄���)��O 7�d�����'s�v�#�4�y�D��%�Y85=�$G ׈�y�c�1P�|�Kr �qў�ҟ�3A)G��G�Ź-ZL�4�m���'��'�*7��4,1OԵ��fՙ_�D��J.j���n�OT�O�'fb�iA�>��0ۤ@6"M?\��91��c~�mD.}gX�Bdӓ�O2T� ���y�I4C<h��^k�	�;[X��'5���"~�-h�Y��D?(� ��jY& �%W��^?��D\צ-�	X�i>�RX2i�zh��`慨m��L�	��U��<j�llZk~�,ztbY�7�	`��x��@�-k���$( ���D�|�T��Sҟ��	ß�	��4�A�PP�q#q�WA�p�b�'�uy"�g��	��#�O����O����dx�r���%��O�ܡ��<����'9J7֦a��ħ�"��B�p���"sG���J�QY��m��s/O|(ї�\���L0�)R�HpcF!
�K%���M�m�Fd�$�E.
�P�H��wol̊��A�X�v�J�o^XQp�ص�L8 ����'�y�'idx脫G	�Ơ�
]���-��U?s���P)�	ҵ9�@�>?!p�������#R �U`�x"մ
 1�R��54�i�����94z0�8!R����	%=�	9�%ڪ6w��ѣ�/ y���胸u��tӆ�R�x�1��៱^�����O0c��
�D��=p~ %2d`W/x�.(�B��Msni����-�������:f�I���A�	� ��� ����	���;�=)P0d��M�\�ڴ�?9���?����k6�$�Ob��U��lz�kD���t��%�6m�O^�O��D�Ov�sl�}c�'
��0g��2���L��ٴ�?���?	��[q���?,���9i]�0Sf��h�A�Ȋ7A��$����՟�C����<�O6-�v*E�~&4ؑt�+X&�K�4�?y���b���?y(���I�O����"�9���@�he�E�&�R�r�i��'*>$�3�������O�"���-t��٥f�WRB֎}Ӳ(�U%�O��$�O���埶�d�O
�'&$]"� ���|��,7o���z"�iT�H'�'И��0���m�f�:gf�.Y<��FJ�q�1o��I矘XR��$��@�t�'���T�~/�t��~��@�B �M.�x�<��P�2щO�b�'^��$��i��g�m�ZA�&��E��7��O�iT��O����z���'��'��E{�H��{��;B��A����>)�X��~�'�R�'2T��B�-�V�LEs��V >���"&�}P\�{M<i���?�����O�䍦ے}AT�\�z iⵉ�&@�����Ov���O��q8��p4�d��Q�2=�� c ��\����s]���Iӟ��	]y��'L�"����	+K��!�o�{�5"@f�$v���ß��Iџ��'i���C/�ʒ77D�ӣ0q�B��O���Um�؟��	Hy2�'bB���O�cw��8A4�[$�ߞh�t=��4�?I����E&
�V�'>��	�?�دv ��B``( ��Tb���2*�6-�<����?��-Vi�O��ܴp%�M��+�<���1����{�"�oZ{yrh�X0�6��z���'����+?��l�-\����M y�$��G[��)�	ߟ�@�.@Uyʟ���x"ݵ_�vMq3�O��(��D��M�ա�Pm�f�'d�'����-�4�8��bW�#hɲ�DԄm%��X������+B�Jmy��'���Ϙ'�B/+ds�c�k�:fs��fM�8&�6��Oh�d�Oh����[Ц��П��I��8�i�k GЏ�ؙ�W�[!�jT�f��O��q�?O�矜�IΟ�� ��� ^-"zX�P�̛5����P�i=	G���7m�O����O��DTr��ODX��Q���H૗�[�h��dP�|T�l���I矜������l��*]!!$���X�d�Z���GͦoK*�k�-r�x���O��D�O�E�O���ʟ4
Q��;b� ��,C�O 9�­Ŭ~�D��ҟ0��͟��I��(�O�,D������יH�(��8@c�ac��Ԧ!��ן��	��x��my��'��MQ�O�δ��.�*7B��uΏh�\��5�>q���?Y��?A��Ac^�z4�i���'���22��/ k��YJk�"4�grӤ�d�O@��<��a��̧��M1d�җu�r �d ��T�7��OR�d�O�ď�>J%n�ٟ���ß��SE����̻N�p ���["��1�۴�?�(Op��K2���O���|nZ�k�X���j��	k��1��%6��OX���9)��lן��������?u��,P�U�?v�<Ღ�%Uș:�O��$ҭ3,�d�O���|�L?������輑H�&s��R��aӘ���ݦA�Iğ�	�?��S�������#��[-=y���L�(��91�V�M�qc�?�K>�'��'�?y�D�<� ��C��_7�U�p ��#ꛦ�'r�'��T*�+}�V�$�O|�$�O^���t@�
�	F�:���*l�E���i+�X�\~���?q���?I�ꏕ �0y�a'G"�h�x4�Gɛ��'\�2$Lz��d�O ���O�I�O��$��w�z��dϙ�"�����H��^��I������������	]���'[@-y���&��j��#k�=a�+�1P�6��O��D�O��$�@��Z�`�I��<�6C��8���2_Z��-v���	ӟ���ß��	�4�	~����۴`����j�P�V�B­H-�N��i���e�i*"�'��	ʟ��"�e>7��+�P���ҡ)]ڥ�t*Y5��F�'��'�r�'UB�M D��6��O8��K0B���U� Xy�Y�RF D��oZȟ@������' �������'��d�p��v_
J��� �@�"��v�'�R�'�L�'.<6M�O:���O8�	^A۪��,��*و���uT~�o��8�'I�D���Ę|��Mc0ꜷZ�x�����"]������Ϧ��I�$��L��M���?��������?��m� >���#��v02#�42M�I�X�A����I_y�O�R�O�M0q�70N,�󇦏�d% p���i����iӠ�D�O0���r�)�On�D�O:\��jU�!���/7��Z�F��A�ED�៼�	Vy�O��O
�)���&��_@�t"�O�`67M�O�D�O2u�������ߟ@�	����i��b#�ن{<���cAUb�T�o�.�ħ<1����<�O/"�'l2�Y�uUpTJIE<!ѥe�.��6��O� �V�P�m�I����	ğ\꬟���/邉
AKI)��uJs�®
��U��h��?���?���?���?�2HQ�@%Dpha���2��P��#SPh�c�i,2�'�r�'iL�'����Ohե�(n���4Gs(!R�L�b$���O ���O����O��$�O@(;L�ڦ1��m�.�{ �V�a/�4hT�M���?a���?a�����O��09�h�$�QE�v '�Up)Zū� �~}"�'���'���'���ib�j�X��O
%(b�	���<
=ڨ�P����ğ���dy�'�B���O�r�OP��b�  8�݃f��5�z4��i`��'���'�x�0��nӂ�$�O��d埀�Y� L���@�m����� �����	iy�'�0��O�S��s����!�R;�E�#k|�+���M����?���f���'1�'$��O=rL�7nU�ۑ�|R8Xw�I�
��?	�A�;�?����4�L�O.��*�M�B�N�HtOמ����ߴΜif�i(2�'���O5���'���'���[ƃ%�t%�UL�Z��Y���r2��O��O��:�	�O$�tś#M
,j�#�(��0q�R����Iß ��%2�P���O
ʓ�?��'� c�Z��`Y�Od�T�޴�?Y.O��c��Ob��O���O��$3L��Xť�[k���`L�-�`%o�ޟd�̤�M��?���?�S?���d����>hO,�����:��p�'�`���O����O�d�O��$�Or��w�T�O��M�ɇ�lxؕ�+��;8�hm��� �I�� �����<I��@�����NV�:�F1���9J?D�!��<����?��K��?A����� h��xoZwU��  @א%l,�2���D�.`@޴�?Q���?q���?�)O�����i��u��%ӳq�2`��F�>́�4�?����?A�9��ӞPj,���4�?���Jv��Ӥ��~����1E�,a"�	��i���'9�S���I'�N�S͟��I�
���	c�+�x���CC�,���E&�ן��	my��8_���L����ڄAE�N3$��`�#D"R���`��g���4��0 �	T�i>�i�W#g������L�>|�]� 
�M���?�DB�0\_���'}��?��OR�&�(������."qB�!A�iR��'� ��T�'!�'6q�0��Db��|���L\O��]ғ�i���W�o�����O������%���I&0Z�"�쓩<��b����� 	�4&R�:���S�OM҉��}�r�:��K�]L�Z�!&~�t7��O�d�O���0Jn�	ןd�	P?)�Ihz�2���t~r4�%d�Ħ]&���!h��'�?q��?�DO{�tJ�'�$=��� �2j���'�J��$H2���O��D2��ƺ�����<Ym�i�t��m�F�!�_�p� �t�'���'��]�p��!zzM@nU-k�նa�|P:I<)��?!L>!���?�b�V� �|�:T��#6�i5��,ਔ �����OL�d�O˓ڶ�7>�� Z����N�����w��{]�d�	ޟ�'�`�IޟT;��}�Ta�!����"g��D���Y9��d�O����O�˓z"%Ӝ�oȩ(G�)z���6L���	QK�7��Ot�OV���O�9���O6�'�� X�6�j��Æɏo�9�۴�?����);���'>��	�?� ���"6�����E��2 x���E��ē�?��<�z�S�������9t8�3E E�je���i��	�v(}AܴEO�S �ө���׷*T��"ϣ0����`�8#7�F�'6"(� I82�|�O?b��56H1�m��R"�hs�^>�M{v�Q#>���'?��'k��'��O��"(p xyS
�Q?���k_ݦ�ٶ�AğX$���D�����"`�a�z��,^a������@4�Mk��?��k�-H����Op���C��h�v�>z�����C�6<��_=G�?�B@�F���pdӢlrVDF�v��t�!�!t��z�"O��av�ܗ\`��.���8,x2�'C���ù�$��'X><<J��6��D�t�㢅���� �'s_�y�����+�[A-�+ 	ҷ��P�Ĝ�a���/�JM�&��3� �h�-�LB� $Mq��[b��^!:���).P����˥.+\`pj'33!'��fZ\�#%��`��@�)2KƫwP� A��؟��ɗ1f���Iȟ̧Ie(�0`�@0CuP �R�50d�!��7��Ⱥ���<�P��&Oxl��M��2s�4��K�-0�l)t�
�
��H��2�L`ړ�H��p<!�#����qٴBO�	."���YnNpe��
�?Q����P�Iy�S�O�0a�e�H=g��|�2W�l4C�4��8۴ �8g ��Y�`1� #�?}!� ����S2媅nz>��	a�T+ЏFQB����u�#�#�`h7 U*0�r�'H�����fm�%B� ,)�T�T>	�OXJg͋+	�DH�ƹ�e���j�DN�Q��ȷ�qj���+�+3��� 5o��l��s�b�B\4acq@��6e[��B�\H����pҶ��O�!ڧ�?��KL<0��Aŭ�@��|�<��Ζ66���į��8}H�c��a�L��$^)Q�6�P6/P��2@
���8�ґn䟠��Ο0��jQ30��E�����	���%t6��v@��ĈG B�Ŵ�jA�J�Zf�83��F[k��ɱJOv�g�	�D���ԡ�L��
��r[Hm�CFA�~|�D�'��)|xъ�^d�'��*W�p�I T�ɓJ���S�H�Zz����Y���Y~���)�3�ظ���,C�0Q�)�(%�!��ǚ���@�g��9���g�(����O(�Gz�Ol�'!�f#ì2qr� �eZ�
��tS���_�pYC�'s��'X�c����؟��'ϖ��q�Y
�b РP?v"Ţs���-9���-O�1a�MZd>OX���(W��K��Y�Y!B%Q�k�P0s�ܶ 9^E���X��ΥE~�♣E�D4k_�(�`h�JG,��D��?����hO\�ĸEF�}I&�#��X#| [�@1D�(��֋pP�D(-֜Tk��a+1�	#�M���Η?�(]m��D��Oz�L:��!�콘 F_;37��������kɟ����|r���|�p#��$[�i�G���=��$�sJһd^&d�4A�	+"���2�����˚yr��²���ҭW�-���ΐ23��!EO#-����B�I60U���]��7K�敂r㓡~Y
�P�o	laC�3 [z��CkJ�u�α��Ԫ;=�"<i��4�b�o;e<2��q��9A�I�%!R�'�ƴ'���F^&��d�Oʧy��	�d�R�+�Q<�����ꏢcX�*���?AÎҢ#پd���Ku�T>�O׬���H�!w�,<Q�%�"2��E�M�9Q�E�U7XM��O�~سU*E�`$1@�E::x$1�K�Lj���O ���ON��,�S&O��ӄfPPm�`����Lc�P��Yx�t�A����4�MT�T�2�M+O��Ezb�Y	$6��F)��Y}b��n�!�7M�OT���O��SFƋ*E.�d�O:���Oh��H�|��58��]�)�z81�%��tP<ɦKК:Z2��Nʜ*��*��(�SG�� �L(	F\e @����ʠD<�s��S&5'��f�H�+��7��h�.��D{�%^�`�ziH��/�h�ڴD�剛i6�4����*�	^ߊ�ۡe[}Rq��.�9w�B�FilH�7�̘E����.�e�n�Nt�����4�?�+ONt:�D��4��A��A���ɰ@mP4�`P(�O����O&����k��?�O-:�iG�J����'�I
a`����)��L�H����A2DBZYE!%,O�E��)P�	g�PK���, _�M�GDѿZ�Ƚ�A��%s�LIcaÐZX��sE�ز!���H�	` �(X�m�-U�F��ΦM*�4�?�/OJ�d7�I�?$1;Ճ��ElO�6����"O>|q�N謠��`Z�R~���	R|���<I�)�'��OZ���<�ʙ�w��8.�]�%E�v�����O���0"�OF��s>�����O�O�0)��\?Y�<���77*Xi R�'z"�`�ҫ�<!��Zw)��1�Í�p<�Rk��h@L<� P�2唉?.pjW��xl��SP"O�������H9v�1�#ˡf���9VOtoځ^#*\	��[!q;�(��$�pC�IH7�%���K=$�b�CbcQ�!�XC�ɓP��H3P��:oX�+�A<*C�ɥ]D�K3�;*�z}�G+ˀ-��B�I�Y=V9��g͎{�$m���B�	C�Lٓ�˕J�9� �߂[�B�	'-VX����ކ���QA��a#B�ɋB�Z'O_�3����F|�B�Ɋl�6H:�m�7���7	<9��B�	�l�@���I9izI��G<Y�xC�	�:�$Q��+̅HsT��iI:x�B�ɸantu���Z�R^$	��.�,D��B���Z�(��T��  �$�T�LC䉘t���1�)̜�p�A:
�B��s~	hc�Ųw�����K�0��B�ɧD���� ֗/v9���Զ6s�B�	� �����6�>Հ��%"8B�I�M�j=�`���M�5��l+\��C�IUq�@�Vf��X�P�R�t��C�	�nt��0�E]�Fb�GӐgBC����q�g�^;|�s�!:��B��G�\x��ˆSc4���!ݙj7�B�	+k�)�7c�O�1�0"�-�B�	�x�Ȱc` ��#*�U	[�@��B�	,jt��g�X�i|�iK�E<T��B�c�L1)���{l1�sEn��C�I�@F�����Z�C��f$Ym�C�ia�苩	�Ɓ㋦���lZQ�<�"B�{'Lu	�Ü���lK�K�M�<ef�>T=T�K^V0��ZL�<�VA��N���jK�z�j�is �M�<��N�@�R4�b�G#E�p�8R�	T�<�W�K�QŒ�{V�&j� I,T4܄ȓD�f��SꞤaZ��h9@=�p�ȓb�&���Z�U� �-���@�{�m���nђ�#��Z�<���G�`�:��_2;��%q����,�=IU��<Q�	O~Q>}S�O #�hJԍ�9�Щ��)D����K�2�y���֔K����M+u�P�yO\�Γ2�bTE��Oj\��Ӿ` ܈�K�g@�"O����c(�CM��-�-�� ��M2�{T$�U�'X����z�lA�BЎ\�y��56 P"`�-nY�d�f�U� ������Z�L9�c�,�%��c�LjS�����(�d�3E/$�2f��v �	�b��8P�NR��d<������S���Ȳ��J�b�Z�"O���6�ǽo�Ѐђ.\>lH����I��H��5+t>���E:p��b��q ��2�L.K4|v.�Y!a/<O��$[<�.�[%i�����snL<&f� �L�%X�*��^'F�0gnF*@I�S��5LO�b
�Fwyۡ�P5	4<$HB�x�K��j�hyJ��D��M�B�ȯ ��1RA�<*�[Ҵ�2�� ��x�c�Ɲt�!򄖘S�� U%�,Kg��{I�1	%h��4��-U2���bĬ7�t��O�E�a�ܺ9�"�1"�t�����H�"��9^0T�74�O��QLR�^��Pb�F*U&�3u��;\M��ⲋQ��Ӈ3p
� �i?B�,��E�ڄ>&>|&��x��U�Ҧ�	����ਢ'1��^4i$e� ���D�j��z�4|y܁��Ov���##P�=5�yÑ���n��`o��4�Wk)O��X�C˅&�d� '��5@����O.5�#�y4���e/\L-إ�R;rȁ�E�|2J%bֆU�6�Y�6�t��!�n#�Q 
�'5$�˄�NFU.�b�g��)D��	RKB���ucP�B�M�2� �i���'i�~��:C��2h��/r��j
)�~����X@���u�|��h�,f]h@�-�	���{e	�#���
O�%̲�=?� 
G�2��f��./9�#CM��n�[�xu{�hع\�jm�+�S�������n�R���&^�|2�	ܫK�.HR��E�� h��9O� ��*�����E
s(X�G\�L
�-h�̠d�.=�<{$�/�4|J�(Fd�P���s�˃*%��Bǯ4��J6��Up�(P`�1L!ZlC�$�P��O]�B���1�a�+�l�*rMF���h&H��k˘E��I�>7��Y�2�F�  ��l3�穌45z�b���A�'�R0;D�7KXf$�C9)�,���O�Xc�1j&NpPu�P!848��$�BO��"�#TL���
[ Bqjt$�O,	[F�ի:=�%3`�\WL	��e��%D\��׫NC�δr�́�yض�� '�P4�E�6O���i�/�z 0U�d@�b�lJ����B� gi���.�.:m�F�B�0���/Uҵ�Or�!�G�A����_������K�_�l4z�� �|}*� ��&���`�R4M��ѩP�=b�!J�D�n�ayR�R���A����Y\�\���ͼ�X�#
���a"���7�㞐����;;
�D��
<0,���#�DU�u���x���+wD�)R��
�'n�W�E����[�PTqY��'����W�.帨uI=2���i�n,~D�V���$�!�t���@���7wvMҰ��=��B�.[^q{wo��&�ӈ�����5�$�
@�E`�jB>��xBM�!o�8�"�A"g�h(���s0�DxrVu����9w���0�9����tlM;69 xp�n�8咈����ذ<��J�:��$u+�H1��kÎ��:O��
C��,�R��3A�,&�����h�o�6�L��b��-+�ɶhn��CX/��d���J3	T�'�ڬ�r�õ&����ݡv�v	�3�U]���īVX̽��<A�(�S����8PH�h��� �0ͅ�	9,#H�6	P1N���5E�5EW���6�ԉ! ���H�$��|ģ��V��I?�N	"��aZcU�m�d�;8H�{�OW�6���6�%�ɢ}�rM>�Q��~�^Z^�a&��S by°�
�}��, ON ���k�b�#g@��y�!R 9צ�ӗ�L�d��`1�	;�"�w�|2�)��4��D��$�Hk~�,�;`h����Q�0�rTrDn����prUp@f�ĦqK|�']�6=:�*'@X�HN Ce�]�״�ҧ��2��t����T�uE;Oh���UG��}R�(�.@�4A���F![�' ������A	�h: �')��A3+pxa�%�.��2�� p�t[A�d�k�̟vk
x�q�Z�o���U*G,PTO�4������ͺB�j,�6�D*��u�P-�i'�1��d�	��ec*5c:Q��l��Si����lI蒃 X���I�sW�b�tB��<I���K�X��N<A�B4B��C�$W�ol��r��ݦA��I60�����"�NU��b+�����Ub��CqY�tɊ�Z�� 9D�i̸�$�.X�Wc#OH������m/��{���VD��ԯ)���m�0:���DƪH���}�ly͟����D��I�z���AM-B�$��c[4za|�/	�y�ʩ#���Ys�K}��̫@D_>q��8f��O���SCߜJ����Ϻ|�)�%m���s���9,�7� ">����S�.���A ��O�Ԉ���SB�}�Ǝ�BL� &P�8�-8!,�>�d�f��q��+�O�A���n��<����,� pF�'�����xML1�6!�>7MO[��D�1 �JQ!iB5b�8��Y�]� �e�1U&U!b� h`ax�[3����%������/��I�4��R�x�t �!~bx{]wM4H��IS�� c� Q0%xRҗ@7he2lOJA��⼻T�eI��9P$W x��J�L� yS�lμC�r��Ϛ�dN�@�����/뢹h��� Eie��2�HO�I��5Q\�Xa	�b̧{� ·B
��aK���,�cI <�4��䑟4ZJ|B�%�G�X��'�j�Sa/�.}�>�C7CŇAb�rش0��$ѡ'�'6hf��,O>�pԢv�����J'Z&�t��I�Y_8�U�u�X\�@Ô���=k0� 9ʴ���I�2�
Qjd��4'�`��ʜ���#�8��<O�)z��(4�}��|����� �g>��6ˑ�V�Ȼf��^����$��}r��ϻ*�8�SG��g��L�ՅÛ�.��F��uTH@x�ބ�8�i>��Sz�iŅ��T�׻G>���c�Q�'u��͎,�hO�U���/3p��pc�i��e����͌8(-N�ArF�K�,�Γ Z̉�'��]�`��L^��V��!;M<��N��@?Rl"G�� ���ɜ�<	�+�2t:aY(Ύ�������'^n$�y� �OI�Tb�.
7X���*V�g�
1��,[Vh�q���?!b���
Q�{��/@�VApA�!x����{r� �uW)� Z���ǐf}�-�3�Y	�G��|k��'�x�h�7�Pe�'^�}�C�Z�_Q����w����ɕ/��P���Ob��^)I8)�S5��YC��H
ԍф勎y#>i��+(x�Dɑ�q�}o�'�y�E�<jmа�L4.�BT2U-ө��D�<1Q%É8ؔ@�īf�m+�[�P�Ic��a���4�Pu�Pؐ=�u�I8V�KE�I�ۗGA�	c�O��O�7�	�I�t���,T�H�B�kO# 0�!�@@�9-��@q�
T>�5 �c�A��0q�� �D�1}	B�5�
��Z ����2d�O�>� pPCslґ@��7�W�J0$ĢDtGa{R�����{ފ��jC=#820�u@U�SMb�0�����!�N4{����"l�lF+K�ZIࣂ�)y�.���d vֶ ��-�+1-$�S�Ǆ:�Zw@��T��Z@H���ȬQ\�i6�I�9�f	(�J`�zՉPl�n���D.$1��r�8ݳ��Fo��m�&b��cG�
�;�t����]p	\���O�y�U�L�>N��'�K��(�q&㙵Υ��딌<B�(���='��XE~2�%���:�Z"e��I��F�S�X u�m�UI��I�n��c�l����	v�0ѭ��$<�Z�j�&9ڙBӓO�Z�j�3逸j��ͣ/��`�&�R��][��$����UJC�+k�QI�插b���BlD�}����B#68�#=�uD�q`�`#2*���P ����}����bpU��_�$~0��!�	�p�4��5$�}D�-������A�'�a�����yy�JM#��=0�4L2~���I�o�T��d���G��mz��'F�	�<����	�8ZyS����<����kϬ^�����5/*��Ǩ*O|�z�I��j
��@H�/�8��G�W���Ҩ�[���6��WIչIqHbr��E8T�ѧ!O�=a|�M�Rט
n��9SB���}�jB�L��y��<�=YJ<QF���=j@�L��9�=�2��|���8�$��K��I�0���+ғU�>U�j�ځڡAZ�d���'���!`��%m#X(����5Ct��q)O��b��R;[W�[��1�bd�	")*�q!I�.TR7K@:Dv7�P%}�$h��-�� jfJ���ґ����)s�}�m�  İ�*u���:���`5/ɗ�>���iт�gG<{�@C	 �Pm��A�=A����y7�C+��iS��D+4���"�kۘڰ>�A�ǖq5u*d�ǔ3+DA�W����Fͮr'�vn5_ӛ&"�(B?�����F�v�v�9�'V\ɒ�i��M�l�؄i��V����/k.d�ʰL�;�`m�0J+-�`��'0��D���=Cp*�����v`J�	ߦ�1 ��8��k��p3�E����	�)�ak���/Zɫ�� d��6�,m���aS9��Ӻ���O�?ϰ�݉XDfT"��kHh!��Z�AlVa� ��
���� 
�dèԂBcL�\�ƴ�'p�%�'9Rȏ�U�@�=}�T?ŐU��m�t�QU퇱#��� <�O���$�X2
����$K�(%v��&��Z0(�O�f��DA8��yJ|�cрH��n�*�*���*�~�l=�r�s����Y0�5�R|Q��F�r�$a�¦&6ꃏ�L�$�'�l7�ޟX�ԪB�ў�:c��N�`�H�'h�x�qӬ ����8l�ȣ�"~nZĺ�� pf0��
��6mӣa2�F�@}���WdE ���������$#R��اuO>�&�W�~����2�Z�<�x��Z�<	4iD%z��P窓�|��T�EF�U�<)Aj	=��ɰC	n�\�Q��R�<�M%\�QSM�O,�T �P�<�s�Ͼi/�@(Fפ)�8(�u��M�<���`�@'T8A��A�/�O�<���Ԭ)ԥ�.T�>�T�Sa�At�<i�b�%3��`C�Z�܌���Y�<q���I4�#�ۮG��Q� �|�<�pM�X����E�I*K�,����{�<�Eɖ�}�n]���#ml�	�Waz�<����9����R�<Y@0E�`�<�#�ՙx!�hq�ԛ gfeR���W�<!��?MB�ڡx� %rtG{�<���Q�n�|��i؂	��@��Δt�<a3��@QȬ��#z����n�<ygM��Fوd9E�E�o��yY�kIn�<���S�B�9�����~��31��~�<�E��s(ҙ��;}�#a��d�<����O����E+7�@];��	d�<qU��
�X]z��1��i!�w�<I��Z
d:�ó`�{Q�AYC�]�<)�k�Q� /D��aW�<y��:
�8"ƍЬr�(�.<T�T�â��r��$)H�k��8R�'D�t����#2x¸��N�=��8�a#D�(�B�V��h$h��h!�ce!D��@�]�)Jȸbdg��N�8$� D�[�f�hn�!�
��z �ȶ�!D��  �𶊖�C,tX{��Q��r�"OH��u�L�Og(H���^�O�@���"O�ء�I�mw�ġ�/�{��1�"O�%X%�K��#���6���B"O���ʛ=^�xa�M�
��hZ�"O�|�g%�4Ayd\ڠ.@�*����f"Or��gHص`%�XR�M�:��x"O�X��CK6VL0A�e'�7ĸ�5"O(Hz�͖�J��1M��+���&"OnZ�e֎>���ţ���t"O4:�
�(\`Ȃ��� U��"O�m����A�Eq�����@d"O�	�j��2F<�3�D1!����"O��Ё��g�����Sk�)(�"O���+A�:� ��p��7{0�!�"O��+�&֎<�h�"�Yk�{�"O8xRF/_+�4 xvEֆwt���"O\�!c�?��-2WF��Tc̠�B"O��6*�A��R�Ň�Qt�d��"O��{s�K'�r��Bj;l�r�"O�pY�%�|0�1�D�8;
j4"O��2#^:7.�$��H�`A�$�"O�0�%��wM����%�X��(��"O�LZs�ϔn�H�,���A C�\�<aR��&R�<Ff���p� D�<�vA��!�� ��ꔫw�4q���R{�<��K�-;pM��)&5�&�RЪSz�<i���w(ȸH����e���z�<i��#E3<	�*g>y�u�b�<����n�~M`S���>Ę��S��u�<1 �_+F�X�a#&ԗ ���E�j�<I3��9q���
���j�a�f�<1�F!jA�(+�HƘ	�*����NJ�<��}*A8e�G�:�����J�<�3���m1
]�F���t1RԦVF�<�A�� G�pQK7D��5ΰ��mD�<�dB��\�F)x0i�	B6�ؑ���C�<q�ɏ��>�*�mI+nzظ���	|�<i#���XX�r/B�z�4�,��C�	%e��A�'ã���C�Z��B�I�tU�腂�%���	�
��B�	�"��X��Ă���X��^�ԺB��i��I���(x����ui�B�ɶx�����2/���,��m��B�I�[Ⱥ6��*�r��MѻF*�B�ɏ|����v�ʭO�L��c)�0�~C�p�R��g%�������g[�AvC�I:�����)Q��h� ؾ=�fC�I�b��Ep��UD|���׵Z�vB�ɺ��S'�_�8�@��D(H�%V>B�ɮ8+R� ���	�jP�!�B�B�4VA���d�~�G��>�FB��4B, �UȚ**u�X�b�[3~�tB��2;��@Ĩ��B�:ɩ�慴HB�	cᐘB�+�.1i�|�C�	� 8¥�3jM�vV��%���C�	�K]&(����\�@�nC�%c �j�)�O�����_2چC�	J\@�3#vȞ�(��:B�IKBX��IU D�M��o�:'�B�	��b��N$E��	S	�HY�B�I��]�# �&t��ty�	�N�C�	&|�v����/"�ĳTc��H�C�+�Fij��U`P(,�c
�9!��C�)� lh����:dl��}.H�"O )9gn�)hrZ��`��3Q�D�	�"O^�)�C�v^�
Ӭ
4bȤ ��'qONH�S�R?E���T�ٌ"R��R"O�a�	�H��B��؊+�~��D%�S�[U�}i�
)��K�(WY�B�	�Zٰx!s��#���p�CX���B��  /.��h�B��ͨB�нtlC��.;�D� $H�A�����R&B B�;�|����=f`��PTI�hB�I)�D�aK��h�q#��vfB�I#wf�2IK3 l\t"� �;��C�A�(���"m���i��_�HK�C�	�k��d�c�ՑW$�$�b��� ��C�Ӥi1�B+$A�b]�p<BB�I~yD�#3n͸K��-�V�Մ��B�	�bK �)���k���SU�KوC��5z.�@��T!�X�����C�I7Yk�-I ��P�X�ΔC��h �8�o��^��衋J�n�:B�I P����ퟍOT�I������C�I3R^�i)��L��PF��U��C�ɜZ�ڗ�l�<�Sd��$�"]{�"Ojlx��Q�d8�HŸhՖ��f"O�� �BX)\�`=�u�:$�6X��"O��M�$YZ�r�mޭe��\�d"O���B�٫|�漩�@�"����"O�3k��wu�%�E�A	[�I#V�'�ўH�"���e���+�R����Y�2D�(a�H�9��<2�gΜ2�: �0D��tE�<S\� ��"6�5`O.D����Η�@ �ib  ̰>�,�`-D�pH�G�VF��c&o���[�j*D��ٷ�
�`5��Ų-5��.D��y1@�����a^bQ#�/7D�D҅E�&w�Pz��*P9���f5D���G�dJ�ͩ��4���t3D���~��q@X�7� ��'�2D�H"��E,%�T�E�Q�`���S��4���<a$a�G�E����{� �w�f���>���T���&��hv�
�O�h�<	!j�B�H�ҍL2���ې�i�<���O�,uȷ�	P�ls��!T����-��!�P)�5�ڐ���2D��Y���&?��z��9-X�����/D��kc��
9�����$�c���q�/D��8R�ЕT
mbG�������.3D���@��%Oh�ds�	Y�~=)d1D�`8'�ڰVl �gK� z���4�2D��A�L-{h�Pr�監�;�O0D�8@��R���`���*z�a8�d D��IҏB
}H�T�`JE�[�$�:D�$(gJ)*,�awk�^�u�
7D����m^Y\(�F�!bF�"�`5D�LS�+�1*�Xq�t��<�t�شO8D�`�vI���	�e�݋hS\�8&�7D��q� S�9���g�)I.���3D���aگpI��ѕ��f	��Y�"?D���0+d�1����t�؝P��=D�h)q��y�M�a�
��8�(D��B�ڈR �{��`���%D��ɠB؜�v��t�V!,���d$D���Rd�e{�f�ӠtRdj *6D�@cTf!(f�q�u�Qa��C>D�� ��cم-^��x��Y�$��4�C"OD���][��e˕ʍ%#��ų�"Ol�i�� �����j�>�8P�"O
u�`�L^��������"O��%(�EG�����k�QC"OX�`��0}(V@) !�`�p�#Q"O"ls�(J���Rm�$.rI�"O,���&�,>u����ϖx̤�e���F{��ɘ��������#2c��D�!�ė$� �Ysb	&T*r� ����!��K5-�5h j�]'�(8�ʙLU!�D͓�$��'��c� ���N�!�Ą 7|�٢^�8l�0K�4�!��d�8,�)9z��CM�2Mo�}��'_��S�	]�5p� "%O��؅��'F��s��7|R��2b�Z�,9(	�'T����C�k���!�W�o�r��']�-j!��4	B|;֋��e�:���'�L����$~�|�@(g3�,��'s�I��D3n^f4� 
F�+��'�֑C� �,��a�	W�y�ƝI�'���Q��_='�B|X ��t��N<9�i�
�G�(:h�˱�=���ȓ�� �B�ʄW��A�-�0$^���;>�p �� {�T�e�U,N�xՄȓ-���Ê�*PD��&ة�>h�����dOëGUP�.�Nq���E�<�3�����Q���Uc~���B�@�<�3��.�;�)�%DOtA1��Qh�<���M���$bS7I�z11%Bi�<ICH% �)�D	�L����^^�<9�n�d�*=��`C�su����]X��'�(x0#-t�Ĭ���������T"O��!�&}��
b��9�`��v"O<�4k�1+��)�!���=i�K���s�O�u2�@��tC81�V���)�h�+�'s����8���P��̹%+&���'
�i���TK�,��	϶�((��'٦��r�D���A+Bo^�����'�u&�� 5��s�'x�45r�'Z�����! ҊL��l�}ӎ�0�'��H@��t���
6	��ap�A1�'��<ো��i�`�{!ǝ���'0��7���焍
� ߮?|���'��I9�(� L3��K��-rPj�H�'����2��Q���)e�,�Z
�'����gSU*�j)6`����	�'(΍0A��C#��p$�)!i��9�'��Qڲr�>��`�P��8� �'FN��PCE7g�:u�w�X�����'�>��DO��A�u��?���'����`��tׄ���Z�F��"�'�tIA�G�D�]H�CA3����'&��)΃L���w�˱$��!:�'':����U�4tZ��͑n� e��'-,����Λ�Vؒ�,ʑk�����'ZX�1Cċ�xe�֍��!�'BnD��KR+o�vA���J��J}��'�"-YTj��;5N��j��y;�'_ (Q�*�g��d��cFs��m��'�0��1KJk�L$�C���a<���' t8�b܃'~�=�W-H�z���'oTɢ����>ɢ�%�K'b�j
�'M�A�'
J�& �E�3r�k��� �!3�F�n�n��H�O��r�"Od<�҈��i�x@qG�A>��!"O�}!�g��1҅
��B:d���"O��+$�P6|�PbD��b�lp"O�Y!�уW�d�aā0U���¡"OD4��NR!]ZX
�i�.6�nL� "Oƽ�'��>�qy�H�%j,v|�f"O\q����^�JS�u`Yp�"OL���x�)8��3 �8�
"ON�8G`�
ڴ�9��M.	�2��q"ODi4�@�<Z]t�Y4��P�D"Oꨊ�a�0P��R�ʛ%n��%�b"OL�S�GC��!0�iIL���"Ox����/JD��<���c"Oj���*�	|(̙�E�C���tK�"Ot8X'��" ��k����k�,C"O^�	QIRWjXŰw�
&6�"4"�"OVER� ��~����#�0C��CD"Ox��'�B�x��5�g"KqOF]�B"O�9� )��a����IV@I6"O�`p1�^�I��S�W�Y.�$�V"O�����k�`�'�Ko����P"O�����wftsq�O�q>��"O̵�q��8gY����M��
H�s�"O��I�〟&����܂��ɳ"OQ���S\i�'
l���"O�9Xw�,�r�c��],]�xE0�"O0��')��U �a
�E��J@���"OF�����3P|0�����`;�4X�"O���	��>噀���US�k�"O��㇢T6]j�M��R�sH�hw"Ol(�slڒ2p�mjѤ�8Wg(8��"O��1���;?^Ș�J�;g@5�"O�����V=%9�ա�IL+j�!x5"O��{qaݿs����iS�E�PM��"O�����E�f���iP�hw��K#"O��R'�<��4�����Y�"OUjt���z�։ �i.�>5��"O�� �͜vT5��U�4���"t"O� ���Y������Xs|��"O��JS`��Z���2QcO)p\��5"O����)U�Y8�(U�� [uZ9C"Ot��CTÈ%��W+nw�P��"O���0�3G* Xq�̈́_d� pe"OT��vEϷF$D 5Dh+�%�"Of��a�%|r��QT�O4΄��"O�Ui���`�ːn*��b�"O*`�e�F�����4+�?�}�"O�h��=q���@ڔ[����"O�Y�&+0(%s`�.R�d=J�"O2T��ɟh��x�ʱM����"O�8��b���81w`WJ*��`"O �ks�Զ#�ڠ;�ĭ��Sq"O��� ��)���T/8؄�1e"Ov����6B	�%a�R�.��ix�"O`�W<���cC��p�����"O6"0*��S�e$rU��"OP�����WRڑ�G!��.Hɛ�"O���K�.�8����� �Mb�"O,�k�kج7���<���"Oܼk�E�%:6����d�Z`Jr"O��q��܆��#�6�t�Cb"O� y�Lշx�l�BRmK����A�"O��6��.~Z$i6��,����"O� �y�	P&�6�`�.��B��UX"O��;�'ǔS�������e}T0�"O�dH�X��X��c�V���"O�3�C��g����W��L��"O`ǅ�'7r���B/ X���"O:@����y�(lʆa�~�tH�"O:�PA�1Նh�q�V'��R'"O~�R1).h��$� j$����"O��ː�E}$`�p0o#la p"O��A��ۄ�pI17M�fp�#"O�]�N�3�,Hê�x���B"O��cU�Ci���9s�!$)3"O"i{ĉ'zl,�A�b�H�"OP-۠#Mt^�C��7J�|I`#"ON����Pf��.ΗHs�	�r"Or|;�K�s�4���,5>^t��"O`(��(@p���럇RP��q�"O���ӌ3@^=*��I
���b"O̵��*�03�Ђ� %u�� 	�'�Z��T��8m���pC��L�`��'�|TےF�D�J�@$�J�8��'���j`lh<���WN��,m��'n��	s��-lq�Ɂ�^��-�'�tec"��9������:IZzT:�'
�1�J�z�*� GS����'Z����b����eP$��>�D��'Hb��K<�l}����0�JP��'}()	���WN|���XQ��(�'h�,�XTm���ł��K}$̓�'��t� ��6�h8��'9gn݊�'�d�i��m��R��1d��)�'Th5+�cNT�W�����'�V�xC�7~&�QӵzW�h�'g��{�n�t��
�G�wx����'):9B׊S�cthĂ '��v&�T��'갨�G��g�<m:`A�q�����'�D4��`��z�X�O�b��y�'\�	 V��r ���[�x%��'�&h���F3e L8�ᑮ��u8�'�p�4H\v,$����5��ԃ�'l�}��.��̓�R�-l��'r��B�P+5��`v��x����'kƈ�A�"x�b���!5�) �'*��1��ļT�xA�b�/@eB�'F�`�7LژD��d;$+H ��ѫ�'tl����?0�$(�m�,o�$�H�'}F�aw�
Bg��E8h�T)�'����5"x�2F�5^�=�
�'<# �-X�N��B��' �
�'���#cX�\6�wk۔fi����'�@(Z�gψ�u����R��L �'�D�i"S�%^�9	�6~İ���'��Yrh�&EL������#��13�'�d�yr��@�2���G����J�'����f��ov�x�� $��z�'���ːA�'l4R�S���I��a��'zIv��]hx�*�)C,(A�'��qS$�͵)�����-I�T��'S�y["��+�xQ.83�'�����w8*��p+7.���`�'EZX���K/1� ���$$���*�'��z�˖�ư��%�C���x�"O�YH�aX�qaĮ��j��F"O�e�$F^�l���M�?>�H���"O� H��G��Ϝ}BG�܏?x4�"O������|Ԯ\ѵJԭOĂ�"O�0Sм��%)@�7�ށx�"O2���aϼB��&G��)���6"OB����S�r�����Ѝm�h[�"O�mr�JҔ���PmS�gn�ܱg"O��r��A>b����V�T2��� "Ox9��Q���ȶ��x0�i��"O�H����`~�@X�@۝���'"On�YP��Sj�00��f��p�"O>4HvG�=gZ&��0o�4�����"OQ3�K�_qpU����(@�"O���r

 6ݲHj��ɝH�8�r "O������8#��p���kӴ�*�"O�U���E#���q��|B蠱"O���Я�#�i���ip�� "OꍚSg�<F>��#�8�zh�"O� ��[+~�FŘ�
ڳu�"���"O��7�X#
��r�>�|��`"O^P)$���(�	�hÝ�LL:�"O�9A�� L6���TG�⨍�T"O>�qb��Nl�Z�EӅZ�Z���"O>8�SG�N�d@2�$X
k�4d`'"O �0��-b�d\` D�$\�0"O�T1P�D0WHP��A-�%�Y��"O(���lj|-#�5�ܩ !"ODu#��D,	,�b��+rn m3A"O�j׈�6Qp��KU!Qe�	*�"O��W���y����{�,yr�"O�Y0L��gy��xg��{��="O�X��ӧ-4�"3!K���H�"O�W˟�
���c�o���ha"O@Ic����Kݽ&��٠�Ox�<YdEʷ
��3�R<:� Y��|�<�u��?v�n ���_/6�a҂��n�<�TFQ[�I�c�ި0�y�"��i�<�6�iq�F[&�~ @Ce�<9a�3#�VUҲ�GZ���6f�]�<!1b͈V#��cZ#��آ3�e�<q�"lB�9�*��qb�$�LY]�<��5ҒXT��H�`iI��r�<9aǇ�-�B@Z��6���T�<9�* �n"(�)Be�O�P�$�L�<��I	�s:`@	�8���c�K�<���\9&��b�4.�gGUP�<a�&�gVґ�̇5#����)�B�<!"��f jP�֫M�(��a��y2�߳0���{�-�-`Y�8
��I��yb(��,��9��=�(��d)ʢ�y����[��Sb�6F2��D.R/�y�FTd4���;jU����y��:�`4�莶Fw`���,��y2�V	d�%(�h(F�3�C���yr���|I�B�E�v�*Ze�S��yb
��s\Q�P�0y# ]����yrV� ��ҢE�m%�Q+��ם�y�o��pU�)�Ĝ�on��&d���y�'�=i���b��*D����͏�y2O]�wZ�hs��?)�y��IY6�yr�R�0fN� �t6�����y�I h~�ȓ�S�+H�qG�@�y2P=�`j�":3&}jf&]�y�[r8R��䂃9�ƍѕ�V8�y�l����d���7@l:�!]��y
� �����3N�M�%�_.��}("OEj�ϊb/�@(d
Q�6�~�1�"OD��&m?��!&	��SxE
�"O@ �q�;&B��D͈��R��"O\`���4U��5��"NnS�u�"OL�Ök�(`���[2��%~�Z�X�"O���Ẅ́���l�G��,�p�"O���1-��|ܚp��B������"O�%B/F�i#�H��"�"���"O�|�6�G(���3�["��l2�"O(h�Sa�.v�r��¯�"r�ȓ=���e��`Tn�{����l���"�\uyE�՝xQ\�����3&H�ȓ�~*r�x�4��-R7r�d��X䄹3A
]VZ� �����i�ȓFv>�L=8x���.��H�F��ȓ&V�]�󫂏n|��1ġ�����ȓ7�4Ҕ�QX�4T�U9�܆�~��mASP��|Z�B�
O��ȓh��Ubb	�P/8�{���8"�D1��hp���Z�z�ѻ�k��	/����'��ɳ�Ϳ#H蛧 �)4r�ȓ% �)�A��074�,��n�p�� �ȓE׌�A���0c�@$b㟟x�~��~YX�����$��<!�Î$x&ɆȓIAĜ��;~4,UIq��p����1 �++��<��������z:ڭ ��A�tƼ(�T�L�p��ȓ,'y��@'f�`h�����KjfA��c�]Y���3�퓴�f����1D���%�?��Q�E먹Ks�0D�\hdQ�	E�r+�,$0�pm/D�����l������A�t�d)CP�.D����`�0��a��-Aw1[ �*D��!'�F'K�`�xC�D`�B*��(D�h;��=<J��@�,�̵�t�<D� �@�G�_Z��cM9PZ~-�r�:D�Tt�͵h��AK#K<u�2*8D�ys)A#��;O�-�d4�U�6D����A��:��bń{������4D�D�vN"V5b�+�do0�#v�/D�����Y�Z+�It�=:)bQO-D� 6��yݸ\�ᇌ�x&2��s	(D��#�F�v����L>A| Yz3" D�#	-'6�JL=,�޽A��<D��PEV&¬�h#�16�� ��#/D���Q��{�6�&NR�`����1D�Tʠ	C�Q���v(� +D�0D�0Qĥ�3!�ő�!*?nN�Y5`3D�t���,$���e�:l�0�P�h0D�l;##�$Nƹ�cM��*}�+D�����UH�j�[d�8� ��R�;D�عV�̭�4Y���F�CTJqKa
;D���K\>D	�	����!�J&�:D� �rjV?p7м6n��"��q	8D��
R���h��]��ꓯ6zv�Z֥5D���I�$�@QY>JL�]{��4D�"��Ț5g��W��^���.D�tJ�I.� U��F�kZJ�q&,D�Ҥ�OYtH��(%�(P��)D�X��♵}��tkA��c��xi5�#D�P���Z-*� �9����( WG-D� ��CE:�h��m:V (�W�*D���d�Ӹ��N6M7*���M)D�� .���[�j�>����O���3"O`��A!8Im��R���4���9Q"O>\s��[V��Q��ё|��)��"OЈ ͼ[A��Ӵ(_��U� "OD�����(X��	8��Μg��y0"O P�˂]9D	hU�+�BQ�1"O��A��	a�!R�!�|�@@"Od����e��"�j���"O pI�-B��@`LȘW\�1�"O���ݷTP��	�f>��3g"O�Pq1@\r���q��b7���T"O<A�2�b�>�P��>4��2�"O ��{(&�JWoݪF��h�c"O��i�y<�� �?,��}��"O�����۹~�ND9��J0��(D"O�!�T_�����=��b�"O��8�ªli����JE��� "O��H�������-t�6aC"O���MB+H=�����jD8�%"O�DȶGŒYtD�2XV3b"O����OU�9��q�Ȁ�"O�8Is�U�yUYR�Tb��ݚ"Oh�*mޕgޠT�B���+Y��["O왨��u�|q�d�KK���f"O	ɣ�ح��m�W�:c2����"Op0�a@�6!d���	K�����"O��҃n��A>v����Y6Il��"O�e�q��[��q!Jy_\�""O�9.N�iVv{��Y^nq��"O zCGќq�乻P(ͷ���� "O��C`	C�:�(c"�ք��Lp"O�8�孆�[0�(RT���m�"O�	4��(��Qga
 ͤ��"O:���'�>D������Nu� (�R"Oȋ�.�w����n�;�`|A�"O<q@�+�)q��q wJ�Y7�e�"O�D)�O�ak"�q���5)Z�"O��R���`�.�qa*	��Xr�"Or}�Uh6�>�3��Y5Z|���"O� �g���Փ��l�"O��L	�b��g�0I��5aa"O�Ţ���7�t|�O�U�49[C"O�$A�hܝz�)5�W�.>��[B"O�=�իH���V��=���"O�p��J
���2�d�&��(�"O�( BD�1D�t�c�S"��; "Of :��L �TAs�� !.�)S"O���4�S�唰�E#�=z�L�SC"OPx!���;��Οj��t�"O���׀>	&�ȶ#D��L��"O�C����b8�`���T�[���J�"O\�J���ꑝ#�^5�b�@)C�I�T�p���"[=]D�2�� %o��C��7m� � Q/L�GƂ� i�B�C��
);,ሥ��f*0"&d�7+��C�I&d�� IAa &Dj6뜚j�C�I�1��t#�[1 ��y���8
�^C�I%��s��	��]y�i�'�P� �Jvz�DҦdӖx��%��'%��a@�T" bp̂�l�d�@�@�'3h�!�e�1z|N�*L/|)��'4d�:bk�͂A�FڐEj�'ޒh1�- .g�j�
�S3(.�'���c�s�ě�Ύ^\�@
��� �c�CJ{�`����U[�� �"O %��� (=e�q��F�R ��0@"O~u�5�A�mh���&N �H1i"Oa�����ف�ŁU�|��6"OV��5�A1�^\�'ѶWYH\�F"O.Tцk˨//0��ҏT�8 *Or�!�׎�v����D�5|�Xi�'�	Id.چl6p�bT-Ȑ'�����'/���Ót�B��Pϝ!��$��'N}
�o��1H�ےA�@�pq�'\��	e��T��x[2 �f��@z�'
(:v��.�Dݙ�d�a�>�'z��r!�)n�bz�P6X�����'�xpۧE��x���4ᔣ<��t3�'���A�+C�@���33:� ��	�'uR��cǜt!� ұJZ�+��mR�'�N�1w�A�DF�Q��0�'��e�e&B�H���G�Ӆ�z��	�'��:b��ug��B(\$�m��'Ab�atE�`�ɫ��U6�h�
�'K�]���)b�}JB5RI> �
�'~^�r��&���&XQ���	�'�,�!O&�HqkM:}}&m��'�R؋���4+���b�	��d�'��9��!ƺF[�8d!B;S�R��'&8�(��Ʈ�ȑh�C�X���K�'P�A�3��oFE�����
�'���t�ơ1���$@�KG�i�'`��Ť��V�xz ȓ�d8Z�'�l���藾im@dI�*�-w����'c�D��.�5�RazP�ݺYp:u��'�2�""o(��GӹMR�x��'gX��)�hg^�&�I9E#��	�'�X�GG�]�5s�+�:cD�2�'���9၏�Yq6M�T��>�n�A
�'�P��Ά4Fk��2��� 4�9B�'���bGj�-eE`G�Dj�C�'�I��͹�L���O�B���s�'�,���U5z��$��##< �'���p�N�H�1��	��!��c�'�JU�C-J��������y�tI��'3�yAS��345��J�'�sk�ݢ�'�պ�eO�@h��㰈�o����'�Ε�s��Dm��bpJ�&T�r�Z�'�j��b��6MG�1Y�H�{�@�"�'Ț}ac��E�~�5.�i/��	�'>�īb‾8z���G���\_��	�'�j�I��yV�xHVɘ,[��Ib
�'��M��.�,	�$٨�C��OS�Y�'�@j��<|e�-����f45��'G�S�K l�fဣ"X�7�@ْ�'��łG��4
�䐅文(���)�'��,Q�]7I�~4:��Em�8��'�bغ���2_2�0�!Wk�:��'E�-A ՁN����@�]✔�
�'9x�i��U�',��1�B�H� �
�'�")`�F��P�L�q2��T;�ܢ�'ߔ�� �FY�^ ���ݕ~8B�'� ��4+h(�q(6�I�{z�@�'�܁"g���@�&4F����'^�R�j�!~�  �$�hc����'SXu���5-ND�Š±b�A�'�*�C獊+�!�FͮL�\ц�h�ᇢcX*i��	�5>�����S�? ���@Bճ
�H3D��R��t�"OF�� #O4w���H����u����"OB8wc԰q;�h�ᝬy�Ѕ"O�%`���z.��J��(ao�YB"O�`i�� �S�|Ez �6�8h�4"OR)��h��Mۮ��!-۔�����"O�}JK�IɖIY2��#=�
�z�"O�� ��a��i���%Y\jR"O܌� a��tD���#��FMP3�"O���è�
Rf\�(���"ܮ���"O��;��m�Դ���Ly��
0"O��5ʑ4w{n�������;6"O�)Yr.���a �۔
�Dy�"O�I(@L��:, �C�G�XU�U"O:x�2�_h�|�zR#":���"O�����/�iPb[�g҂麵"O���cĞ�{��BS�Y 6aJ�z�"O`�!ȜJ�N� ��ɮ_A��"O� �l��k�ّOŴG1�̳�"O,(��<k�B�!�.;H���"O^;���r�����D�Rl�&"O^����I�k��@�͔�*� �"OVȠ6�� ��h���m��8W"O.("Ǩ԰U��C�擯h�X�"O����Cc� ���$=ۈ!� "OP�w��"j���ꥄ��{�h��"O]۶�~8-��M�=e��"O��Z�$��^6	IЍ�	|Q�!�g"ON��ւ���ņ��LV����"O����A�NctpJ�&4/_$���"O����/�N�C��K�fAbP�d"O��P$�/\�֋��شp"O��b���?��ԁ��i�ļȠ"Oj��狔��lYPΈ8	���c�"O�l�7��X��X0G����"O:5x�Z!*^<BR@ Zh�"O��%A� C<��o�3dG����"O�9p��/�"u�RL_�[6���b"Ox�I�cH��;%�B15�:�u"O��f��x��K #}T��"O�H�p
Q6E��a��ȇ0e��
B"Oh�cׯ��z��a�矉ZS��R�*OĘ!���<G�����/jƑ��'�~�����s󰬸J��& ���
�'=�X�r��Z�0S�*�3���'��]�P�N�:J�EJ!B�$����'���8�܆Vp�P�[���H�'����s��q2�Y�� #\�X�`�'$����ɟ!r�-��*�?X���
�'c�4Kt��)����q����z\2
�'N���aR�E�*9��	G���	�'��e�D��[^Le2 �Nt��9�	�'#��%��j�@G��{0 �B	�'��4�U�M�{!�I���x���8�'�-����&7jt�y�-_w¶��ȓ/�ec��� �ִ�5��1����ȓe�hN?cL>����0��h��x��Lp�@�6Uyp���Hk�$��qx��C-�<$�<%!��n���3]�IE'U�A8ZA�aN��N��ȓ|4�A�b�J�"+.� ��\8*�l��'�nH(0ŝ��X䪃�Ɵ6�e��2^Ȼ"�8�r(��$�Tr9�ȓ�l��AHF���*�F�
j���S�? ��gbOR�|t!��	I#�T8�"O�i�mlV�����C	l��!"Ohi��GW�i���󬒄	ۀ\��"O�)�IG<(̎��"�2\�~0K7"OHQ۱�ľkƔ���6{ɠAP�"O�=��Ҭ9�=(G��W۬���"O|]HGڽ<whQr�bS�U�� "O.d�%#�t�d��@�V+�=��"OX��+T�6����!��-Ql�y��"O��� �0x��$�-TR�u�"O�;�l^6���Ӂ�MD4ԲS"Oz��0���o�MyE�	c'�1�"OT9�ao�5ld�b��.-��q`�"OFŻÀs�����(byBAq�"O�e�2f�
�L<i�d�(y�`z#"O������]��\�R�P=hbd��"Oв�!N!f��\��"J(='�R�"O�D�**P�uR��ϯ"%�u"#"O�%A��O3kc��b'ЀY�§"O6�Ң�"SJ�Eb�ƅ-q���d"O����Y2	�V�:�Dα?���+1"O򭓇� �fy�M�q��'I��H�"O��P�Ӎ;kf��dE�%Sn浪"Oؤ�U��z�v`�$�a_b4�Q"Oęp�o5'��I)�$fU��J"O�Pj��{��ț��n@e�c"Or���1��ОD����"O��P�OVJ���£+���Q0"O����Q�D���d�41j��q"O������x`�g$B[&8�x�"O���4�ʦ|�L!��>d5�"O���-�?����
�R���	�'� L3���Ož�ѶN��z���
�'��X�&G]36�Z�aw���n���'�v���kS%|E���H_�u��E��'�����"����ǐr ؠ�'&$�W(8�l�Hp�p����'�꼺 oH=5o�����_�n��q
�'����ŝj�, �E�=g�v!
	�'�f)�g'�:if�a��4�E�'�ޥBA��Y?: ���|��l��'�� #V)C`Mx�B�I�t��8+�'�VD�%N�_,�����eJ���'�Ĝ � >�d*#L��-s����'�8�6�V>w�1�G�q����'0������H�������U�mb�'ABl�gnR<D;�HRL̂>�n0��'ڞ����1<$41�`99i��P�'(�j�HκRJh0���$m���'�~��N/���@��ͺs<��
�'�@yҒBU�g��� �K�P<�	�'cH ���0�ڙ��S�70����'FrA5��&@�f��g؎%l��2�'��I�<��`��\�L��L�
�'�PI��e�m�����-Y�̡*�'���J�#��BsH�R�h7Q��'fUY��H2l9�M��	+	�'�2����:-������\��'c~�P��Y
l����w	�w�}Z�'��vFĹ�a` 'Y�m?fE��'Gj�F�ۚE�
�T�"����'�vY��&(���H����'t���Mȏ�H��gδ� ؀	�'����`�y)8�B�	U9/G.M���� �@� �%
��l��B�ar��s"OL��G�&E�}�ī�Z�1��"O0l��AJp��Т�@�VQ��"OP�)�}�X�臷�Pi�&"O~XC���%j�+f舝H�N\P5"O�K�K�1���3�L�(}N�9�"OJ`#ר��FH��1�ȃ�U||��"O�(�B�D21���3�-��O� �rR"O�$(AcZ?kQ�[���B��Ӄ"OœV�	V+e�B�ƧM,�1u"OBQKwJ0A	H��/ØZU3 "O0�������rO�=��ȥ"O��k���o���#TE@�T�^8��"Oa��)��:|�������@�"O��DE��i}�I ��Ҫt�|0R"O Գ"�I�[(h�٦�]���[�"O���7oW1i���q�h��%�"Ot|��)�y�8��HЀ�X��"Op:��Y+�s��	���k!"O��ç�H
*u��*?s��@�"O�K,76����L�� Z��Y�"O��1P/
T��l��K��~r�yk�"O|�H�y�t�@=���W吗[!򄀲Lz",qdͧrJ�$�!'đD�!�ĕ1�(9�F&�#6����W��w�!�$�#)��dKßV�\���V�"�!��#`�-�#lB,���"o�:c!��_
eZ���2� @c w!�ќSP�|0(>�V�ŦD)!�-F��ݨ�J��o0.��CL�=k�!�ĝx�cAmj��6l'R�!�$P6���`��M���bJ2�!��JFT �.P	h:I� i�u�!��U�}S���c�\�-f\�a�c}!���^A�jAg1ޅH�J�L	!�dk�q�ƈ�}!�2�VsU!�D�>:�0���/�R��G�E!�IY��!q'7��M
�Z�a�!�dF�\N�9�@�m��I:/ң+{!�dn_Ѐ33�)V�du��b !�䜯>8�A!$� F��5YSϒ�o�!��C|T��ѥK�4v���D��y�!���i;~��G\�Gdb}�3Cɮr:!�0	�8���Y]~��b��LS!�$�|kJQ���cU��P��O#!�D�c~�L2�
Tb �]��ܠ�!��D�[1��Ie�(1b�8a-w!3"O�T��l7L��\�CO�R�r�YW"O��I�h�:x�`� �K�'�X�J�"O��&�E<#�6H��ȉ��)P�"OrL㖆�`4�Q"�	,�y�"O�]��c��?��)E�]>*)�p�"Oz�2��?��4+yat�!��N�b�����<]�:)� a��6�!��U����
����T��ȸ6*>!�!�$��xo�XY`�W�NY��#I@�!��82Ju����2an���ձ2�!��:͢���O�z1��U"ɑ2.!�$�!zO�=
���,;��K��
.N!�$�<W� ��닒�r����D\$!��߿'�ޔqvۏH��h��@G!��.G�a҅�I�T�,(�#j�1E!�d���u�늞#�N鸗�3!�ػN4ā�3f /T�)������ $$q��$C��1t햮J8��"O�E)�#��z�=jw.�)��|�"Oj=�� $+��XaJk�rd��"O�(�"�D:��a��]�2�0!"O��SK��p��(��C�R�x87"O��+d��13���PJM�?��X��"O��ٕN�K��S*�p�2���"O0dc�$�q�@�pN�'@�$8i�"O�ӆ�5 ����l�ɦ"O��JuK���ّs�Q"�v�2�"O�"G�2a�u�A@e�"�P1"O��2ӯ�H(.��qoٔ2�@�p"O��ya�V<a@бD.�8�(�u"Od]�L�9F}����JQ+:��ݣ�"ON��⍆D^���l+J�"Ox�"wϕ0(��P�mJ�X>X̉�"OH���KZ��(Rj�=D� �g"O� �e�A����V�'`Jd"OR�����4�z�ʕ̀'o��0"O4Ed��r|�KG<cvջ"OX��0�M�R��ҧ�A0���J"O���Vd�-K�əF��F�Z|r�"O�@:��I���c�@FP���!"O*�3q�c&�}"��L2Y�z���"O��X��2VϤSׄ� �2R�"O�ݪg���q d|�� A����B"Or�ab:�|���	Ϋ6�F���"O�q�G�!j0}��	
��qY�"Oj(C�#U
��xѤ._"��g"O<�Hn��]�,�ce'Ń#o���"O�����ߘճGŋhcp���"O8I���ѼmI:  *�	IG|��"O��`*��,3>l�a��!:��V"O��˗F=L�����/68�<�h�<i���u|�Yz5/�	+�v1�ǋ}�<٣��oB�@�LP����[E�<�I@�:t[��Be�$,Gf�<���?$x�ᭂ�__�� \��B�I�
�ޔ��b�,`���uh�B��(o�T�:EM�E�Z��n��0��B�	!baĥ�������B�ɦ	l���P��ajq�L; �B�qC�(G/t���'�_	}F~B�ɥ#4�<��C�U�ҵ�P��='� C�ɾ"g��+��9+#��V��B�I�VT*<���ŏ!j��Ơ�xu�B�I�"c�I�S.��;{b��a\3��B�ɆH~���;2Q̛�%�&"B��%�hࡠ�J���f���B�ɝH��&	������(�g2�B�ɆJNm��n���
8g�,H%D��@!+�9��}j�n�2Q�8��e!D�H����e$Xɗ�U:|^�h��h<D��+���G:JTP��Ӷ�,��w;D����g�!?�
1�d'G>Zq�IH�N:D���`ˁErĴ�dJ��tܠ�B@7D�x+(ÈI6�iJ猓~*d%#F +D�$8DA1��K%�o��h@�)D�����۠:�|L�FF�\_��`6�(D�D;j1S�r$85��K�踷G1D�@� @��$?�uiG�L�vLsV�#D�,�eҧ"B\���<(G�E8�,ړ�0|RI�,��a���j����N�<�&e?H�h�7��0[#�K�<� ʬ(sI׊Xhh�%��L�Aڶ"O䐃�`@�b��,3W"M��JAR"O���Bj�3) ��ތ���q�"OR#vEЮe&s4��3�@���"O��K+����*s͒(�V��v"OVȸE/ĵ%θ���+��&�䅰 "O�Y�4��g�<y�����u�q"O �x�
݉Y��h"��8�0�1�"OfH�T���	r�h�Ji$�S"O�7n�,�
�Z���d9^�Q"Oε�'�^�C�,�êɳH�TY�"OX}&*]7R�i�J�7g��)j"O�Hb��Y�G�"C�I�N����"OB��Fg֚[����� 8 �$1d"O��4GV�?�����J�Q���3"O�i���,�
�G�$��"OZXHA��>Ғ����jR�P*�"O�@�2�,?n$�¦�X:G&��'"OZ%�'h(1^�Գc,U�98~�إ"Ot�4o�/ �:a�7��;o�^�'"O�tB�cљC��*�KJ�:�6���"OZUi2�ѭ^�"��5�����q�"OX�%g�-P��4�Pቍ��4�`"O��R
<Q�Ʃ�6K	o���Z�"OPpy�G�Y�@���i�^��qv"Oڌ�@M�o�"}����S�"O��Q�ݢ��[�������"O��xЊ���w�@-w�:ċp"O�-r&�:e��bР�+7���b"Ob �R���a0u1�^=`�"Om�%J��2t������bH;�"Om�&xkt���HM�`p��"O��
D ��YU��C����cQ"O�L�슖t'!���O�)�>Ɂ"O�$��)G�r
@�
Xd��#�"O�p��O�-0Ln�z���.V�S�"O�%C�ŏ(z���0���1D�sd"O�U� ��P}�����)�<��"O\��#/Z�Pp�����>��7"O�<�tbӯ"��\�f��	&�.mPW"O�؁���( �h1��S��x+�"O�A3L��F������ �(��ii"O��z�61��\
����l�Q"O�EF�ʨ*U�L@`��M�����"O��P��'Qp�	3Aӏ=���"O���g�U�*�ڠ����6蒒"O�B���h\PXS[�+̮�1s"O2ѣ&�ٹh�D���*�3+��F"O��Y��51[:(¢�I�@V�E�"O8|��ó|�6�@�"���r"O\�Z�/�ʮJ'���*B$��"O��Am�$�8�2�k�0,P 9�"O$�y��SnC�5�#k�:-�]3'"O�1��GSXJ�y�
R.�,
2"O��#%�fab��t(TA+��"O2 0s�Ǫ�a0i�(I���*�"O�9�sC@�o~�,[�%��|iy�"Ot�R���^uX@G[�r�&\�"O&���a��d�B���)6dx�"On�Z������Փ!!�"OY��3֖��E�1h��G"O�1B`(�� ���!�� ��Q"O0�a�a�t-;F�[���2 "O\1AM��(K�g�bK([0"O� ��9�AU�N�<���%���U�B"O,������!T��%�(�-�t"O�� E��n�F�h&.^0&�,�`�"O�
Q�'S`����lX�s���A�"OL�S��.C�8��M�%���d"O<ɨ��M"�ȈmC4k�R�8�"O�\�/�N��U��M���<�"O��1���+>�<SJO*pPm2�"O�;�hA�Ȕc�挩��;s"O���$���d����ڮ�IV"OD�P��ܷwj�|@�%�L�Pp��"OL���� %�}S��>_©�"O4iPQa�!�����|f�(;D"O��Q��N3aT�r�B��dx �a"O
��`�H
`y@�[phJ�A���ʔ"O%Q�-y)ԝ1���@娈h""Od�Y�͔4&[�t�!��{+�Qf"O�t���5�0�R�Q�`���"O]��;w�����@ҳM�!�DJ23�<��
��!&	}g!�$��A�$c�`$	��0T��8E!�$H � äf		�p���R�D+!�Ոy�>��6�L�SV�PsB]�t�!��&����$�J Uנ�!�䊥}T�<��NAL�*Kao��$�!�B�C��G֧)/"��7��:f!�F�df>�R�#,ơ`�(R,8!��X�d=���V�qd��xҡ�l�!���^O����Z�]J��B�O�{�!����$dA���>-� P�.��z�!�d
����ŀ�%�)���!��hZpQ�/��[r��ƒ=�!�&���`wL�!>Yhm
��!�D�.�bѻ��Ljj�B��+�!�d
�w��Sᑱ,m}`$hŀ~�!�//�H�#���pL���p�X�xp!��&jb��J"��"g(]j`��Bq!���w`qr���i�ea�eF>,l!�	�Q2��eF�T$�P d� >`!�dՉ>�!���
�WG�H����2Gy!�=�yx&�Ǽz<���d&w!�DQ>g�|-�F��9�-:��=Z!�d�צ$�֯� �p2b	�lF!�䍼+��{���:�Y ��T!�$����DTC˅_p���|�!�D�%R�5���ħySԡ ��g)!�~a����=��s�C�*!�d޹%H�=YDC�L��<k�@:!�,@<�"g�S0U���R�Ȏ�!�D�^��t����A�J�D�� !���OW�Q@�#S���Y���.'_!�$ɏw�J�ƨ�#���p�D�=�!�D�3�4�ǂ*k|��5�&�!���	{�9��K?�����k��3T!��N�B��v+y�< ���([;!�$Q�RpZY
�F�*�Ĺ�"Mʚw$!��J{3����O��`I��!�dC-Ҥ��HY��X{��!�d�$���CI�+j��*���C!��/��i�84|6�{� �d�!�Ϳ}qPL����"�&���͞�!�d���6��/\�7b�th�lԎ4�!�_�C*trq��r5�<s��=(`!�$+ms���־#������	B!�� Vyr�([-?�@�#aN.(ݞ���"O|	(�'�F.�d)��W{fLAu"O	!r���o�d PD�ad���"O���'�F9z�
�y���[8�蠳"O

�'�9�:��`IZ	S(t�"OMI�"ZX��IP���5���c2"O0ݫECS`8�U�=���ɤ"O�*cO_�A[���!�"��2�"O���C����
C��,���bq"O,�a��S%b���y� ��d��y[`"O�Ī��J+VY��S y1r�{"O�MD�8z�xXd�.�ε93"O��BLM,B�Ԅh�� })�"Om�A] zw5P! �_ż��"OZ� �X)J΄A��/XX��=y0"O���OD,�D)aL��?F^���"O�qf�/&�vp;w�>f7u�U"O,�r͛$W�V�!��~2A��"O^0�C�\�2ǐp�쇤7�ش�"O�D� ��3	�	��K27����"Ob@�TD��i"�ʀg����"OtY�V��>
�� K�HT�G�,��"Oj5y�΍�R���C&hH/}@�ٓF"O�,�����Nز�(�K$>E�u"OęS��\�n��Z3�	V��܉P"O���"�<�`��f+�F�"Oވ���7)�Y�V�!p��*�"O��"+@�z^��C�6U�0Q�"O2u:��� 0���&㗻+�	�"ON�����nAJ,hp�V�t��"O�Q���˴K��á��$�:�`"O>���^ftI�[%U1n��#"O��fb�	>�d:��]5�	�"ORL��	G��J���ME�t
")"Odⷆ�`\�DmP�d �ex�"O`k��=v�U�@R�9)�"O�qj��6T��ۖ��8p���P"O@��t��n�Bm��$ˊwO�|�%"O�b��8l�Se,p4��"Op��@G?+|X�K��D�/ȁ
�"OL�zd�O�1�ȍ��ˁ6�P	S"Oh�D��,��L)1 ��lgR� "OڭYӮ�H��@إ�X��F�`u"OعZ@�S�/���I1�ȸ�$���"O,���������{��k�"O� ��Y#t�y陲b�=�"O���"s+q�z����$�neCG"O�%����	��`;��;�"O4�a�(�*jz̫�AC$r8�x"Oi�2�޲(��(��9K�$�"O>	Z�AV�B%�3��8G��V"O�<B �ҧ#
�U[Х�={~ވn,D��R 	QF<��Ɖ3�ڌ�5� D��C��Bk/�U�ďK�7d�#e@=D�l0gB�h��`'ȫi�H	#c�9D�X��ٮ.h��cG�	M��%D����F�rx�'�ĪV� �ʃ#%D�� av\J\�7�4&W�<Ӣ�!D�4�P�ܪc�qCC��v��a@��#D��;�@EEl�D���
�(T�q��"D����K߯8�`�D�[�2����>D�\����*�X��F3n��a%<D�XQe��o�5
5�E�zB�����5D��:VF��nf�E���>*φ���3D�� �ȋ%��:ݠ��ƫ�U-,IBB"O�@˱OL�)��a�щQ�:�4�!E"O��bӦ��X`>�@�J�n�2lY�"O������w4]��,��v�܌	C"O�1!P�T�s�[�퍆?˶�iF"O1���C/<�耲�lМ��MX�"O��3F���9��4�N8�"O8�d)o�Ӧ1�`�"O�8��EҞZ�Z� �\&��"O0A����-���/ZlZ�q3"OLx��C,Mrn��`�7x�*�	�"Ob�5�Iv$���_1�ɲ�"O�,��HBv���ޤp�����Ʉ���d�p��J�D��4����3�1��"O��ɲ��=�:�Z󍆮W�t�h��w��z��퓺"�@U	0�ĹA��-�e��[����d�w�c���p��l8AÅ#$��ǀ�K���vIti��&r����X� �aŘ��"�EI�sfl�ȓ5S�5r�ç\[��ѥR"XR��>q�vAԭnO��T2D�2F���B��ȓ^���x��D�5�dH��$ߗ%�P���>j�X;��$\��,6�Q>xq�)��<c�Չ�Mϯ2��\���!0�x��
�=	Ё'sV��w,Fd���V�m�"�ͻ2Ұ�a�M���I�ȓ9��(z��ߦc��)�k�M��ȓx&T�Ѵ���Cv�11�X)�p`�ȓ��HJ����G�P�!s F5RXņȓ1LƍHP�]�fd�5�W/9~���9|�P���4'O��EN_Zm.8��^" �r��0�E	�[�*��T�?ш��~�3��M\�1�Чo����	9�y�-ƽGC��h�
D�3�(SB��yR�W�WP����� 0~��3��y����rk|d���{���A셛�yB+�L�TÔ��!6�{O��y��F�M��a;7�DI��h��#ذ�yR�4_��٥��Bb���G����?A�'w:�AF���/l�s m�>�`��'�P=�rEI�5;��Җ.5�	��'"$�9���b�q�6� ��	�'��q[�"ח=���zFk@�*���O�=E�ą\��jIH���cI�E��B*�yB���&{� �k�P(��%���:�O���ï��8�ܑ+0�
X�<1�@�'�<��'"��q�gE�V��!	��ϭe����'DɺD%V�`�>�JФO7N$5��d$�'q�*�ӄ�
%v�l`��u�nl�ȓ5�҅�����`�˭9�R���Bё��}����	��	B�=B���K�<'�U�r`9�!�8)���p`cID�<Aձ*<U�)�Q�֥�'`�:�!���W	�t��l]����@��N�0/!�$�}��e3�B�o��Yj���=+!��	Y�vY1�HQ ��$񶥔��!��6.R��a��$�܈�ã�!��/R����ԟ|�Thd��H !��M0�{DC��q���)����qO>��䉔,���j���x��1K�)�P�!��ǈ�\K�kRE�2�Ӂa�W�Z�Rw"OV���B&=�����<Mc�"Oܩa�LϦ3P؅��O�Yۂ�a�"O8��7���v�l�f��(C���i��7C���%�� r�[��� JWMBE	v�ʱ�DO��S��I.�:@��e��_Bʵ��,�jB�ɼV�qy� c @`B���N�O�➌�	^�'�]����cC$p`��OL�ܤ��T��,�u�Բ%ﾥ��ƍ�#$$���Иr�)zR%�*�5V%��s�'4�=s�� 3Q���G��e��ay޴�~b��s�ZI#r�^?K�m�&oS��t�E"O^�"	Ёt��V��E�B�#e"O져��ج��6�*E��pw�'�qOZ�p��Y��bk�,���BU"O���� �
C�DaZrD�q���	��I_>1�a�% N��``�9	�( �,-D�(	�@Ķ���QЈ�� Ӥ����%�D?�S�)�8�Y��ڏ7i�La��֓�@Їȓ:rЂa��U��1q��
�A�ȓx��B@��IF��aF�K*���J�8@j�����=S��X�ȓ>�I��Ç.�``�j͡uЎ�ȓ�Jy��l'�|�q)�"-��-��%Z�ð�^�lN)A��G8��'`$ HE˭p�Hl�#�
^�؄�
�'D-[�iݙl��a�˟P�б�
�'a�ɄI7@(�I�Gʆ��M����<�S�t��2\^Հd(��t�X��P)��ybEE�^P�cȗ�fmH�`��7��L�O��O@L;��C�|��tAs+Ӕv���"O�1��_`M�H�r��5�v����'�8�����i�d*A/Ĳ[����c�)/�}����!&, `�CM�"I��2�L!D��qꆃ�b�˅��]U耒d
"D�L�d�߬ߨ�j�g���}1�"D�ԙ�޳ \AA�*�	k4Y�k+ʓ�hO�W@���рj���hAoQ�U��B��+J�����h��aӂl�!`z�B��;��\!	Y�h���c�˽_v�B�I;4�(0��"R {||��BF�1|$NB�I58������[9!],1cG�\�&"=��4Ñ�����#+�� G��C{������a	!�d�3mT1�QiW�'^����k�8X��IV��H��� ��T��Sq�Y�<�8�S"O�=���
"�ȹA�e����Ɨ>!1�O�ݫצS�z�|���d�8#�hA���'y���i�b-9����8;B�â��/<�rԂ�'�.�a�IF�M�RE��F�J�~	��'KD9$oQ\�Yrۤ���s�':��s�b!�üct�+�b��yd�Yƀ�[�%�1-��
7��*��Oz#���\4@���\�rx���b�C�<aq� 7x(�сB%9\dc�e�<�u�S����xQ�X�=	�1��_�<��} �R�V�L�j�����@�	q8��i4JZ>��p��*%��ٲ��(D�pK��
NҰ�т���\_��G(D�x����G�|P���ڃo����%D�8� kǖ*N��;"��zєR��0D��jE�	=c�
3U�-vr���,D��KJ�����U�ѓp�V\��,D�X*A(Y�K��J�ώ�p.�	q@=D���Ė�e�ݒ�l�.5� A<D�x(䂘?Ts�Y��Ln��9�6�'D���'��	Yz���E�ĉ��d:D�XyTa�!td�$$D�d�R؈�6D���o�#z��Ӏ �<}� HRJ3D�� faҐ���T�(���T�����"O(�A���1�Q4́��d;T"Ol}[��,��萇���iѠ"O�
�cٮ:���S�Iw�4� �"O��#�:5,����S� 5��"O`�#�,�C&>�0��S��=��"O�d"u�[�Yₘ#���l!"O^t	�(�5�@�ec�����$"O�=9��\c
�,!dbP�?��4��"Oܱ"�_�anDJ��)�T �"Oj�1m8_�.�c��.����"O��(v��*pr@�$�2 ^�U"O�|��Ѣ.lt�$�M ���"OFI����1��XT��?%"����"Oh��V��S2U�e�P�P�*O����S�W�TY�"��zV���'�\`�Ѫ�-��eQ�O	wς�8�'��u����+D�I@ߊW^f-�'F�Մې>�hi`�%]8�'��T�q���@
�e[�%Ќ�.��'
��FcFT���a�)(�\��'b���n�[	zDi1g2p3�р�'�Zth�,8�D�a�N�hHR���'�j(F�Y���h�Y���:	�'�k�-o������V��͸�'J.`���ܱe���a"�:�,h�	�'�}��ڞb�J�!�#,��̲�'�$�S�і*Q�\k�m�*qxHR�'�"�"(II�}���S#;n���'#$�*��	/�$�
��`�(�	�'_�(��H#l�L�Z�\98�1�yH��
7�ceNn^��f-�-��'����Q��6դ�B'����'X($fEZ� D�px�OD tq\(	�'T�)b�%wM��,E�Q��	�'���QdO�zD2���AC\�,���'��`(��g��љ��K^4��'�
�e ����J�L޹E�9�'�� ��@A�	�p5l��>T����'��X�e��6��`JD�2�Dq��'4�M�gʴ1/�!cn��[P`8i�'z~�{�&ԧB<����IE�(�
�'�����ƞ*)�ehWk�!Mhl
�'y��Q��*��ŦR�A|�!�';%�0@�T��=)���?J�t��'���ʅG�5N�I� H!��P��'&=���3��)1�	�
R
���'���I��%����!�c���'�dE��Sx��8�@��f0.l0�'K�tB�T�-��\*A�'Кx�4�G�]��F�+@:<]q�'���GD<^ ��`��;��(�	�'�-)��0n��uP�a��>2e�	�'�NM�#�	S�,�w=�4Q8�'�^�X���H#���O4�&��'D�uJD��(#*݀�`�/#,U�'�DA�F����h�X�c\�h,�4���_="��D"O�����_)K�^�¥ѯo ��ґ��xK�]�>L*˓6<<KEJ\\�Ba&�L�,�>����(-�4�[��2[�,]X�CƐb"hS�@�1���%�2��s �֜]�i�BӺ-�D����8�/��!���-Ղ�H��)ϡ*��l�g�;eZ�h��9X�!�ވmn(H �Ek����n��Ѐƃq
�a4FM�"x,t�F�Oll X7@^$��Y�̂�.�!%�LE��>Q9�$5lO���g� e㘬ΓE�N���ɛ�j)c��B���BT�;��q�Q�3@vxhd����O� :`ё�=Kی�	�
߃]f�`$��. �p("���]m�Q�V$�W�����!'�ؐu�
�� �d*(M��� p��"���'�9�J\?�9�c(D��(��\2i���ӑ!\8�N�@�������!�C�O�.�!�w�<@r7��;Y����ğv�^���'��@� !�ц���Z�2�� I
m0�A�hu�𳥭�95����@��%�$���>X�>˓U0�]��.8�\A��o�3N�4��I�9�Ra�f_�K�(hu�z�ځ���]A���W��/i8�=�g���be�N"���S �$���l>��'��B�c
B�8�c(cp�z�!�.;��04a��q8h�Z�֮!��cF�!P7�G�nn���,`W�Q�6Jt�,�EL''�2uJe���?!f��LhԤH�3�l��u�Љg�VL�L	R�<� -��Z��X��'fʘ �O3�d��H�˼s����RE� p� ������E��t��LOS��E@�%@�%��� .�?,L;Bk͕n�Z,����d�"��|�&΄�&���A���9' hk�����"�N,�d�!d� 5�̭J��ODKҧ9���R4��MH��5�8I�� ɯW�܈[c-v�`�H�I.�*��;29��
�/���٨�bK ��O��5�Ǔu�^a#��5VG:��Z�U�l��T�v��}+���?z��Q�m�r�FQK�^�PL,���'�U�L*aoP/3'��Q��J� ��~�i�0�0��D��:��+w�z��&aAdJ�p���RW��!'� �P�P�I��rG�٩r��-*B+�!c�53L�,����
E!2�~l��` ���T!��&��7ˀ��t�
�L�ʘ 2 =+��@��E��M�� �Dh"h�ۢM�?P`��J�I�Ԥh��?.��l�+O�DえԜ�nq�!��kL�:�P�����'l�)A��ف,�fZŇ�8\l$q0&� ����͆�D��9�$��9����J�� �(Y�\L
�����Xu�)�t����Otܨ�胘h9���?�@�@��_� �!p�P07=����]j��EȂ�a o�et\�����9�,T�S& P����>Ex&Ɂ]�J���'P��ja��@9NX3p`��j3PHz�hѫp~�[4c4$�v�e�D��l ��ǉO�
 m����Ż�D<@�n���:Ac@��lKA6�S`M�9+���B�/���ꎹ��X'�y��ϕ�u�}P���Y�Ll�bWy�ܾS�T
���a�%p�c^��'���A�N�r��Q�"�S+1@Y`c�@8���;���f4*BۻP38��U&�,������ %���s�c�Xj��:Q,ށ��OzI3 AM�;J��Q��SD��!� � �(�3dݟcg"�8�I@�$`}[�� =G��)Vf��B� �m��n2���ě�eꞱ�Q�ǻn�\��bO�8H�ч��X��(⤎&�8�Ã�P��b�����'D�Lz`O�y��w��S�����Sd��.߿��^�>��|�D�>B��;�%�%�0>boޘ/w"�*�O��x���V�gм����NL̓!3�=R���d ��-`Z����_+@ �@�'�@��$�,XB�#*^;7�D�b���R_
�"��9^��p�U?pc0��5 �+&�N ��.[9�p���o֕=��$�2OŃM笩;Q��(M�|i�SO�#)�P�?��a[bLq�DϾxmM���P�nʼ��U�^L���g&�w!�6�͙\mRM��i��4��c�E�*��m�c��uI̸�C\jԾ��F�'���Q�(�
vY��'Rt�B<
�#�&��ᗤx&7MU�$�LY�c��%}*�ʔ�'#�J�0��wK
�ȥ�T�B�8u�f��{�jh��'D��ẇW���U�Å_|�!���l��L��;"�8L�E�3���F-&O-V�[bk[{�[ 
�k��V�K~�%T�p�(���>HM�mcg�C���'�d�d*
+G ��)���x����.	I���nڞX~`�� ��<=�&e�阅e����	�@��
�t��Ipq�'�� ����Ff6h��K[��%�3�����B�Y��p���I�]���Y��ē-�<I��Wg?�E��$��v�d�ȒO��p\���DH<AA�W�*��%�
9|�dD�׈��79�"��S+����"$t��0��$K�r=ɲ�*��w�6="��}r�[3�%~
Rh ��'!(D�7@ąGa(.L�I�H�im�)P!�'WHn���e�(�vFO�xM
uG�NP�	��l`��Q�󄈯	�f��ͩQq��6�O������Y�p���W�0xRlZ�<�v ��.%�A�A�xd��ZA�Y1+�r�:RjP�2$�7
)�zBi�r�J@�� 	%���	���lbW-E�=�� ��8z�P��	�%w�\l�`Ȋ �Ӡ	���֘�;g��`�!V�P�bt0ԅ�a�\��dW�`s�({��\�6�����J��U�JD�B�э��q #)�+�Xaj5+��/��h����5����0�T$R�Ph�2(ь��U�D$����� ���B�Pe�e*J�') �D2Be,ؚ�i�Wf�rw��Va��5j��Y܆�R�Ǐ,0�3�I�M�u+�R���u��Rd( 	 ��^��#<���.��@��_�d��37�Φ�µ����\�S�,ܷ|��ݐa�N.Z%�ʕ�4��u�������e�	��ӡC�3#�hh"��2	�v�H)�>8�=��I�\�����P�]�&�P@��>���x"���s-I��N Iz�3&_
@r��#@�{�0�w:�[�._�+���ʃ�Q����Qԕ�E�ƺ���C��ުɨ�a�M\�q� տ?��yp���)�� 3^����ռ��1��JF�9+O��j횆@7�Y�Āͺ\{0����Dφ4�M�E7�t4��)@s��T��C�[ഉsi�+V���'�3˶�°-ٺD�����	P:�kS)W%�A��I�M�-(5 �"&� ���ݷ��H���فW=Br�T#�I�O��:ШQ&Ԓ���5i�RtHt��=�m�ēK�ʑѣ+� }��h2�dN>~��I]�8�R���'QG�ȋ��"K�΍ɳ+T#{��\Z����?��Y�? �1/KJ�xT����'������8M�3���0B�i�N× F��1�@I�x��a�$�;� `9d��`�w�P�<���&K��Y (?�F͒>l�Dĩ��z6��H��@ܓDx<�u)��l��][���5�����d� [�L��	%�x ��
Pi�b��t!Ůz@@qJ`�G�<��nKL��wd4OEebX�`SҔ�$��!�A�GQ�T-��sƅ
O6pX� ApaR�B?d[܌��b>�a$G��Ӄ�{�,1��:�*U��⅞:�����K������~Nx�)H�f�b��4�]Xc��G��W��M	�W�K�����fOHh�A��XT?Y��N;o)�0��$�&Ԉ`�$ȯ�����	4!�-aD�3⢙�Ӄ������$�d�+v���41�4y�*�'�HB���aL�A��O�� �k@%�h��O��05���J�e
qc��g�ҥ���òX��\ S'E*�iJ��'*����6~D�k�Z�1�GHP��90$E� ���hI\Q ؆���
g���U���H���RESRT����F��^j�E�DN_2+Z.HU%�e���E�?z *ʸ6��ªĥ&�Tlb�*�48H�TSdC�!���$K�y�Ve"'�/lŮx��&R�M#� �I�v�̺�K$}e<,�,�g���(O���hbO
xCv�E j��F�'ܘIa��|ʸ%P���!�9�ph�y@d,�B��A�<���] �T��G&�O hW�ӛn�8�dڀ1�V}hT�D �O�.rw`�9L����&�3!����j�c��ǃz0I�3��Tq8�EAOB�<q��^<5�u���#s�2��P&����,P�������iB�>��B�󎐏oT�9)DĂ_r�`���t-!��J��a�e"e�Zf03%�T�6\!�P�&�#bY^�yó�,	s�M7ʓ9lT���KC�I����e�Ɯ��	�"ܶa�,xP��B7Ԙ�3��3���˒�W�g6(# �<�豇�I�F�����҅]�@���iɄz�X������<t�,�XrM��0��]�vUbR!�xb$��p* �夕�d�jt�i�|�<��bT�oJ~P��=p�*�3&� i"RI�vƆ&΄�{�K��e�*��"4��8���$6�t))�!�!�v���\��!�o�.P�GlNY&�h�C��@��͙6�B�x���镂M5W0*er�m� t����Z3 NF%��#C�b�^qC"Y�c��z2*X#TMʤ0& Y,l�Q�G'����FKɦ:�L DnP�"v���h�(n������:��}P�F�4�d�b�x�qOH!Ӈl�>o����B�2�b�!���}�����?:��9�ꂺ4L�h``[T�~Y���k�'�)6c��X3��(���B�v 8�Ld<h5��C5��q$-ƀ�	�~�A d��0D�9q
,5SQ���-������%}��)�S�<���T��V�"�.��0���޺Hܰ�����E�5�qLB�=�衛�M�qO�Y	 NU�pUtL��I(�ƀ!F��(�I�,-�4�b�M�d�mq�n11zt��M>`�����U��<[#�נ)���㑁��;�az⥇&�`�i���#��ո'���ՇH�*6R�@�I������[s����[04�e-��o��K�����*E��'�����b���G/��W�xl���E�zQ8/��^�05�~��Y�M����e_>�)7��T3N�|m��#�3#WRy�"O~ԈA'ɫz� ɓ��\	':���R�~����J�=Aޭ R�:-�nƝ&�����Ǒu(��'�䙸blT�6ZpI{R��#�ڤ�ߓ&%*���o����rߘ��9PqB#�d�@ǧ79z�AP[�,"h�W�wyLu��!&H����Ĕ1�X<
B�Y�l���8���׵FA�88�a�
/n��$I0�jMSt$���
pB��E�u8r�©���ʱ� ��uꆔ �:�{���!\�P�ףٯ[�|da J9@�"�a2��}2���
��4�[ě?=�;rZ�9�@�!�4�BiN�/C���O8|a@�'|��AO�v� �/IVgܘ�� ����0Y�Y ����&L:����r�!xψY�D�<O}�-��Q�ڜ� 4T�{R)M��V9���Ip*�xd�;,1h���rv�P��A��{`S qv0�i���p<��`��m���s���%Z��9!�MZ��<#h��g �t�J%#W��N�.���G2x
�w�PU��C�,IӢ�tQ�Ȅ�DF��q6���V�D5�Î	�j�^�c�ߘ���(i��)W��r��	j/L����6�?�ϻ`��1�g��'J2�I��Զ ���ȓk�����*C�`�c�W/W� �hQ�*S&�*t��9n]�e��?��E�(F�v8���6}"��&V'��Y'NB����1`����=����� N^h��Ƈ$R�d-���]�"�D���-#��C��V�+Н��}���r�=,O���KQ�h�X�A~��}���6Q��a�gW#5�ܩ,��7�[�2tǍ�_�� sΓc��2@�ʏU�,��O��pi��G.-H��>
,�xc	�v�lPJ�"Q���T�҈f3��PW�F$F,q�w*��%��u���͞�6�p�I��y�FճV`��bP�y[�%ا�_	�?a�P�/G
����^|Y����t)B�4�I�hg��h�˝&��5z�o�'7�~��D�'6�zݙV�;� ���݊;�l`�7A�r-N��7�:4�x(R���0����ݝN0���K2D���4BĮ=��y��b�jx�`��	�>���#�S�O_�����E-c��
u@¢/�Y	�'5�Q��G!A\�·�ޮn� }�	�'�p1��.(����@���gKX���'6ʖbC��\J�e�X~���'�Z��v`�2=<Ġ��Q�q���D��a�ԉ�TH�T�5��}���w-���y��J�D����xҌ�eIՌ�y��K�\Mvij��F��eC�L��yrbǉAꨡ�g�(#<@���H��y� ͢�(��Ț���*T���y2� n�<�ɳg����`���=��>i�����B�1.�\��F
 hr��ԧL��yR���3<��ئCU��:�84O�7�y*��~3@���1|Y�p���\(�yb��'�`Z��O�H��@��y���.�"��v*��G��LR��Q4�y��Xkp�Q�Ê�8w0q��l���y�!��,��8���:�4�����y"�)
�����&�
Ye���'��yB�X d:x@rd�\�:6ZQ�R�yb��S>q��O&I��l�S"D�y2��)""�P�C@<@��]����y�L�90�� ��*\�-w�Bǔ��y"IK��R0h�̍lft�H�����y�h����T�/���1
��y���|�VF88͢X[7���y�EWx����68"�8��yb�P� �V邓'E6��̓R&��y+�0���:�L/�J��nQ2�y��,cz�P�&P&%���1�=�y�NB4<���h��W-M���d���y��Ӻ+y,�� �7�؊E��y�'R�_L�����R�\|�.��y"�T�z�C
/F���x�Aܹ�y"�&'2H�[��];+��Q�Ҍ��y"D�����Cmǰ"Ȥq����yR���{8���F�09�Oً�y2�]�v�AI��/gt��+.^��y�B�|��Dz'Jމ\A�I�rc\�y"i�7e��!����ZgJ)1����y$�$3.��ӄ��D�\��q�\��y.�9���Q�L�j*C�j��y���3^LEx��kU�e[�d�y���y;�=2s�ǍY���s��,�y����x�`+Q��p�7/Ũ�y2
M�JD�Q����T�E	B�5�y2o2fi���O�N�̀B�D��y�hX%2�hq��h�P��%�RBI��y�e�@�r�+�'W2L͈8��e֍�y��c�$`+�̀4o�Qyue>�y��7,4YtS�v]z�U��yB�9"Y@��l�*FT荀�Ɖ3�yRDɋ1�x� Bi�VO48��-�7�yb�P@�J�5��1v���y�?itf�B�/$V>YS��Q$�y�&�Z�*�@S!� n��� ���~BA��C �x�y����38��h17�P�`��+!O#il!���:F!���ʛs�D��4OҼGK�	���X	^���<�1è]C0�A�'F�14�h  GZFx�``�ڇU�� �w�p"s#A:/����Wf�>k�B�+L
Y�pł�#�εheA�7#=�A��%��a��S�1�� �aA�E�C}|D�,�s�|��"O�p0��7�����Q�|�&I
��Ў�h�iJY���O�$`*�$�I7���٭��ɀ({��_=;��`�d�#QH��D�m��-�PD��<�$�'.^̌�c�V�H)S�iܹOQF�2-bJ��ȩU��	�d��g�'�����Đ�u�8�)��:d�p�0�{�h3X�| �mդ�MK���qm�{�+�E����� +>�&a��5�)Aچ &Լ3�bj��ȑ!M��jB�,�R��-��� �D���$�F��,�Z�ዟRmT�ɑ�M mO��2IE�?��Fd�u�B�N�uk�UX����>ȮI���?4��1#��X�c!�N�t}cեM6&<,P� E2�����7TZ�@+R�C�	J�Y�� L�rmS-O�)yg�ݜ|B��k
����Ha�'C �)+����^v#��J�E)��B�D��Uְ��� ��1F� ���sCz0�-Zl��?�%��S\��zD	���6�:�AÐ^X q(�e߬F�� :q��(.8�%Q�PX��B�i�#�,�RA�YVU��$�B�qЭM{k�� ���YI��K	�zڂ�N��x�S`��|^T��w͙�-�����4.{P�'�(����]�z $��'������wΰ�9��Ô��J��$m�n�Jߓ5OhY��.��Gȼ�	�`�D���c,�$��Kǯ�> �@K d{�X ��v�x%���7O����L['��sG_�t��ku����C�)H��T�/!���;���s�.~K��b�o�e�:ۃiI=�$��7�܊���3n�b���� �s�ށ��I_=�HvZ���1)��	8h�vh���Y[.�b3/*����I�^0���u�ڣ2��� `�H�m�ft�壘]#�%�O�"�����G�-�Xt+����q�V�~~��J��7�x�KK4Oڸ0sf\~�H�C�(D��t�훀3d�%��!��;ܕJ4K�6IԸ9P��]�h�@#*A��H۔)�r.X����ʍ�t�"窂/�p=�Z8m���(��Pb�$��b�߃T��="
�i��	�b��s K-OZ�+���@��Y�NG�9�`�b�D�!�'��X��T�Uj�i��m $g�5ى{��0�����.�a���*#�jAc�~�ȓ�N$g��B���$��`2���9�x��K-Q�ڐ��"�������M�=�WC�=LU](��8�݂$��z:�Ụ�t��#�Q,˵���t��戃;����h�%�P��c��m<L��A�/P#������<���FW"d�5�W�� N��e�%�P8Vcj	
��x��$�DLݦ[p�CU�>AT��9J��n�\���7��i"�!焐�pڐ<��i&\O�5	�.�!��A�qB
,��''TT�s%�<�l�������9~=
��Ѣ�F����tJC	Z{��ӗ�<��TC��p�"�F�j�9�ӥUCܓ5���R�@�k�(0*eҗg9�8,�(�����BL�s���Tp�
 �i����D����� 8�V9&���&ʚL�'���*@�	}$�PЪ�<K_���.Q
�xa�S��0��$�K�g���B����q>�( J��MP�6-V1Y�8��V��9K�}����Fט�$E*��?a�J�@iv�ɢ�҅�������zl`$&�(c>E�(OF�Γ����B�E�r�T�w��4�ך4 �I�I�1����'��gH�i�T=b�)�~0$)u+	*O�(z�[<�y"r���tJ� Q���d�H�y=>i��ȩH�
1U��#n�,Cw
P�s�P�O0PP�.7�	������\��(��<� �B��l��ӎ��8�`Yi�n�L��䢕��L2l���W1��}���\�^%�DCF�'f�,��+P`{C��3-V�QH�=� ����50I�hc�k��#�ҌN6m��iD�:�b�`v
�!�6{%3DK�Z|CġQ�a���d�/�\��2�G�?6�h���3��ՠBOD-$v��#�˦����R腈�e�0p|8
!��n��._*9������$�|�C$3i�����G1;C�����?��,a�JR��c���/�h�E]4����A޽D�,��b+�-^�9cK��Y��.�9(�v��6��t�P'SBB����vhQ�?U*��n;�QZ�	�"I���`$ �W����C{Ө$�Å�+l�a��Β�]����2k�!9SF}�2�Z�L�>y�嫚��p<�3�'	�~���P�k��QO��85@]��	�[~	�F�)�5��U���	68�X��HQ�4�YChۖ ��!ʄ�R���$B�O���xbg��b��Q�#�Z	|*��Т$ dq�Q��8��ɒL���2�Y�xW��¦�^	,5�Q���!�%
H��؄g�A�R�Z��7|O��!$�.sg`��n�Y�Z�r5�G�g�ޝ�ee�Z���U-īVl"M��]Y����\�T�:�!� `��c�X�4Lؐd@�0 �bؗuv�)�I8��3G8:-�d��3&ƚ4)��E1,�� ;4��3�?�H�y:���4��,�L0����Wpzy꣫HH��	��ɝumB����@0X��OB�A��i�z�½x��D#[�*�I� 	pfTјG�܊E;N0���C��I_c��T��T�@h 5�Ѵ�P"
�KGj��"/��82���ΟX4�8�a�;JV��。����%">���dՌ8>��a�_;���A̠8NZ٨s�B�,�D(A�����S�!]R;ў訰Kˁ-F���� !w�Hǲ26آ�`�06.�6��1*�d�RaB� 4��s۴�,�6�\R-B 􆓸bjL�w�"�P�j��H�fKx���Փi���m�@n�	��Ɏy�ҼBB-�>��i�Ę��KM�$�P��c� B�rl��!/l��-Z��лM.�x��G'4��FJ�b8��%FK�a���P-
�j5�}ib'�[k��a���	ߺ�٦��#|X�e�K�b���p��o<�Y!�eޙ�$d��k�$�P-D�#=z�`G�.�OVɱ�ƺy}�LJ��}-�i���T�\}Xi�JB� n��GB�o�\	�'ԕ)�4�8���/x&�E�f�0[rFU�2j�<��	 y�8�E��B(@��U������D��nEj�ʧ;'б8Ph�<,�LY� P����M�^k^1�c���X� �z#Ğ\����D�1%�֍�5���u	꽀���%@�k-�]�|� g@�o�"�[�"�ȱ녋W�v��!ф%�V��5{?@٣�b�!m=���c�ƮC�I�J#�``gJ�f��Ћ��?)?TH�ĂȄrx�p��M�����d݅p���.	�Q����'��dĒRFu�%j�Wՠ��
�}�,���?�N��o^�$���B78`@x�cB�'0����A�[ۊE���9!�d2CJYmt(��=OZL���Τ6��с�O2�"A�9b��Ń�_O��Q ���%���'!ԊE��VSi�T�@�H�2�I8��>jx���-D��wjF��������<Y.�~�x�:�+(O iL�e�H�(��Q0.���:Ӣ �S�R�(F+U)�2��6!!�lՏa�F���q>�3��к3vI��*�JQ���$y(LuGҾd�ک��V��-R��L�s��uʠ&�H�\t+�"���hW�Y%	c���T�5V���N��r��Y�p��O?����_:(ݠRf��~~�H��i������䟞2U6A2QĆ�<3`��d��qwlX�%^�Y��47���C[>dI��GO\���e+3s:��'<<P�r�]�^s���'�$5�$&7d��IH-\����{$�/N@�9��I�6���@A�KIx��Ԥ�!z��@��+J/�`d�'��H�z�R �#i��	�Ja,Q�e���
�ax��ɍ;���"�޵(�ء���ě0���Ѓmя,��a�mܙW\��I�:�ɸ2�?�HC�ߓt`Q���N -�r�håR�.$�P�����Px�AX����(�f��s�E4��1 ��'�����=9�Dx��X���Fyr��>@8�`��Vq���͗�p=Q�=QW&A#Ea����T=� �,ɾq�,� ��v7Va�#���C��|2扆	 �� ��ˋ#�Z��Sd_��'�l�2oC 4D"xx &�
Q@ ye�W�!�&�S#�h�b�^�2h�q@� �$w%�B��-FZ��H>����G��D��D�|�[1��vo�$+4�H/D��)�w��	0�&�cl���5��2r��Z	�'|�z7ES��He��H�c0f���ƬuQ0�0�Մ^��QI�����u���N~Q�����<T��+�(��H���%lO���+x����%ř��0�!��̼)(�yg��%.nհ`��D��Ы�"�O����͛HT����Z�8c��u���3M�r4��3Hb�xjPJ�(�$�!��hbW�@�b����%U�~���!0B�@�<9O#M^���C
�Md��3�; H��4��>��\����99ڸBD/��2�����)���0d5�G$,v!�d�Fd�"A$�;���$��xL�TF �H�I�@#��Jm�1�qgUDb�z��ĝ�K�nYc���0d���D�)m�z"���Z�x iW���p�0y*�G٪�����땃ofR�෇V(s��z��(�Z����Ō�{��̕<���A�4s�qO@�Pd[;T TP��ch�Љ� �2G���'S'�}×$�N��	�/�8b�:��ȓ	dl�d��5<��X�Z�+^�p�`'�J��`(3#�s����B��|fb?q�1� 	A���=7atR$A�L]�7"O�d����!7��1��rrE#u[�p��n	�3��j'� Xn
EʶK�8*���+��' bIq��K���#�\"R�s
דf��Ts'��"�4��DH���<I�@a	�#A:�����,trѳo
����;c8h��ኘ�����
�
7�qO��S�L�B3���@W$MВ��<���r�"V䀡7h��>�K4H;
�p�sH���x�A��t�ؽ�-˹~�"Tt*J0�x���8ڨ���N�B��t�J$w�֥�#m�|���l��K0�
3b2���C%q�!��(D�\(lL��9�c��Ԝ�VL��T�!���2�1��i�&ם0\`,�2gEbfȧO�,�F��ԇ�7r��I�R�W.��=1whX�/^d�*�@$'�T�����	xXh���5��q�+�(X�X��1�Dl�YiC�Y8��h�d9��|��f/_��,s�,�ɒg�N��b�u)"���ˌ�X��16�E&�#cϐ�v�P�Q��-��M�R�B?1�C�5=0Np��J^d7�L���	<�I�s��%	��	8�H'��+�\�:?PD� ��f5���������?<eI�,B��DCԁX{�<��B&m����%]�� �e�	%*T�f�[t�E ����J�b�4yK��Ů?�,x�>��/
M�mSdk؏Wr�1�h|���XE�Z�����0�K�X�t��-�&Ip�.�(Fft��e�	�]�8��Q�S�堐R$'O�0��BN�&�!v
��;�V�5�$ҫB��Q	��D15�a��Հ@|0�z��۔c�\��D�EPT���!�2@��`.J	N����P;�!bŀ��+ؖu�`�;DJ m�c��P,�2M5đ�>�	"� @��	i�ٲ0̕�1H��e��mo�A�Ad-D�hg�H�H��e����~�����E�u����d��p�`����۩Z]����J��MA'�V{��9ըdB�m�@H:A&Y1������$`�	�J*=ܺ4�#n�>0Q�݁E-ĝ����cW�<�j�3sE]�[�L�q k��q>ayR�I�w�Z�h�ǧ-��uȴ��)�O���H�Y螩����M_�����˾P��$�Ŏ�!n��xc�eQ�J/ ��V�
$'��C�)� DM�!j��Cq* �6�յEy\Di�FT����tg�kPQK��ŔkB]�a�Y;Bsq����/MQ<��e�������yb`S=D�B�8U���H��!e��?ITmS���j��)QR��d���7��#q��!�Ϝ���1c7�#f�N���D#g�J5 2��"���{#��T�������N)�Ɠ5�.�b�B��13��FpP�ȓoRL@w�2��قuAB+:�X�ȓ,8,M`�1I^|����+0�P�ȓl�mڀĒ�*N��C74`ȅȓulm�к�� �ɚ�"�Z�i(D�h�Ф��[^��ɵ� �Rf���H(D������r��۔�� �
�҆M&D������]\ �;C��$��ݓ�'D�Lxs�ɤbp�I��N[?1����""D����/�~(��eBj�l�e� D���w�'l�jdHA� �.49҄<D�(��d�)U8�!hJ�>� @�:D�xCQ���&�B�٧M�)K���t�$D�x��*RԅC?1��З�!D��s�I!,�q�'.��Ʀ�a�@<D�p �/�#F1��yÉ  &�,P1�;D�q@+@+xpAP,��pÄ)d-"D���I��A<5ڰ�@gpfȣf�#D�(�Ϝy�D�4��6{�(3��-D�������A�r%�	f#�!G�1D�x�S�]?�x���kZ�����)D�0� Ld�ƌ�qJY4~��-RRF%D�X�C@�bų�&�egz�"s-D�@��k Z?� 3*�`gR��/-D���e4o�Zq�]G.�&*D����KMޔ�fg�I�0���C)D��6�Ѭz��pȕŘ0[�E)�� D��ɠ�
=\���3 �u!�j>D���V�LyVm���A>V�8s5�?D����֬>81���¥#	�s4�:D�$�T�&<��(4��
9�G%D���l^�y��|�`e�<C�\;e'#D���.��	?q#&P�_#b��,!D���@��LZ�*�L->T&} )<�ɮ9[8Az��݋�6ṄA�,u�c�x��fϹ ���H�@�`��.�dE3@�h�����*��vn׀x~�%��J�}\�9]��ч(Z?�SŚ"]�Q>A�6č�HoFE�6B�0|y��9�I$kB���F�k"�6O�;&�<%?������K^��=��*ƌ2b���ܰ�@�Ȟ^�`� 3&��1>�	ɟZ�?�����'C_��-K���z�@P�m�%�Pݰ �ɞ,���g�O��Z@���[QM -�2y��4C

]
"t-��6�ցP���E��O�.��;�BЭ/�Q�e�$�`ܰsAШ���'	"��)E�������A�f����*yP�q�k�y��G(
E�����(:,<��DB5*���)C�L�ZA���'Ԫh2�L52�h�
ç%��%��(��t�4�� -&�q��D0���	��j5�/O��?§�����̓�:d�X�b]0yC<��f������)v��(�jW�h�}���;U��YW�i^�=Oc��g}�V��{�O&]2p�A�b\Q1��e	�8�����#���DD��"��x3r�S�R
��	�t��	J��O�q��� ���(�� 1Pb��o�ڑ�b�iAܙqŖ� H������)�m�O���I�B�!�x�g�E�.f0+f	�T,v:�q��R|�L<���
��7��b�=��A���5�!��bE�<�1�Ob?%���BQz`QW��6&��Z ����'�J)U�O�\��t�]�<�i����U���rO>��%� U����>�"'��Uj�`͗�;
n��Qc�>�B�Eh�f��<E�4�� 5��&�Up�  �Shy~	Z�
ܨo�Xq	/O����'y:I��K3�5q�F�#3�P4�7��$Q>���y��)��١�L� NF(�9'D�#�����ݦm%�B4ں����O�uru?+����� ���(t0S.J�W���G�U���)�k�|5Mt�7?!�� Ή���͙#4X9� !�-��D��"O�H2���$�C�GUH*��&"O��	��U�R����7�B"$>�1�"O�1jǮ�*4�(l���"O�������� �ԬM���"O>pJ�AQ$Er��*�&���Bt�"O*��A��K�s�
�b-�IQ%"O���5�
6�� �K��c�P�"O�y+�LŲ$���@3�[:M��$3T"O֤ۇ�S1�-�v��5��Y�F"Ov�!�Ɗ
m���Yw'�D�%��"O�Y�&D��oO���ѐ272��"O�� �I�v�͊�)�	���p"O���
�F`�g�ӆ$��1i%"O�t�M�'K���)۵vj*P��"O���.��p{
철�҈	��"O��{0)ݘ DVH�'C��&���"O�E{T߳:��U% T�|�4$�"O� �(E3Yϸ���/\? ����"O� �E�l��`�R�|�l�p�"O�|2���S�N�$,�P�>h9�"Ol}ejU�/��i��M�=�8E�C"OZ�(@fM�9/T0 � M1���"�"O쉱�ܰ
��A{����%u葃d"OHX*�g�#w��q,�<$�F@3�"O�(�2E�4%騀�����Ji��"O �A��V V_�x��؟8vaz0"O�;B,L�~��瀐0i�Xp�"O6X"�	V����ƀF�`-l�ZT"O@丆�D�	�(�����$�""Oܽcu��'C#: ���E7
�x��R"OP��(�Z�ڱ�¶^@�"O�l����2b���l� ��Lk'"O�$�QbT�o�$�2�l	%����"Ol���7�>�Z��
�81��"O����?c����S{���G"O�!RK�6<Zx��JŰX�$��`"O���h�6J�L�%"�h��!�Q"OȨE��T�D]�$��hDSg"O"��K�7A��`3�l�(�t	�"O����� �ةP%ڨ)��rv"O�4 �#�7^ir�ʖ�1L9�"Ox�x�M	���$Q$�)� �R"O�0��8;���Z����dkg"O�@�EIW�I`��n֧:�f!��"O��q��9�"h��\�J7x���"OBu�'Q�v� aPKQ;a$���"Ot��ֆ��p�~-�5�K�4
�ȂW"O��BǥE+�l 2��ת;_�Hy"OF9�d@1�:d�
�~�Ph�#"O4�9���Z&�\*�*��m6pQ:�"O��	Z6������7 �rT�"OlU�'/05�8P@��� �� )�"Ol���aH#cެRm%8h:�J5"O�U�A��7ULh�bb��9����F"Ob(�&` r��fꝮsH��B�"O�<K���L.�a�I�U0N� �"ONѠ��9+*P��v�߀?*l�7"O�����(O�yE�� D�ąW"OV���J��g�4��DT	D���(C"O~yp���=l���&�k�h��"O��ض�}�@1���l��"O��"C�����ң�Y2��JD"O|��B�=~_~}*e�� E��"O� j)�ea�4"�Б�%-ޯj(����"O�����L
zN&8��lH .�FEI�"O�m�'�*y�r=���Q㮸*a"O�0����n��@���WL;�Q�q"O�ő@,��k+^t*�K8���"O&���!��Nj}��)�/2U�9�"ON�)�T)W|N��c=K��,Q�"O:�y7nt�G�j�,�"O�}���X�j���!�I>R��{�"O �݉P$����e�F�t�3�"O��Z��ö �b��T�-?\�H�"OƩStF�/H��Ups��(v�Q�V"O񰱉�`z��ӃBćW�P<k�"O��)!J�Ix�u[�g�c^f�B"O���FB�	Sf��&�Z2UJ80�"ONე(��O�4����
`J�Dq"O�5��oFXIy��BF!TD��"OĒ��)���Y�/ȬW)8P�"OT�8Ɖ[�F|"Ȃ��"gA�"O�U��<&�P�`�->:T�W"O"����cE�hR'��[����"OT��� T#=�\B"m�'e�(H�"O��kM&1�	C�l@9m�-2"OZ-{j Z�T@k�+L�,��"O4��G1bx ��)�"O(l��A&���C�iBM�BY��"Oj���-fq�d�$�B�r�A9�"Ojib4hܟ
�B�K1 9S�`Z�"O$�o'/�.�B��7t�B�"O���qɕ�bQ���#nը0���"O�m�4e�l?��jr&S�V���@�"O�lP^�((�`B9�}j5�B�*!��-qt8�����@W?;�!��!	(,xj`��g��z�C��g!�3i��1၌vD��C�
+H!�DĖA�L3UN��IA�uZÁD�o.!�$�u��5B�b_�d)�hi�nٳR$!��Ċ1`��Op
�a��y
!��*�=P�a�KI��+�	{�!�䖋9�N��
��H4��XC*U�94!�d^�u��C�	�f������v!��472����F[�#�.3x�!�$5������n���4�$6!��4�͡���
7$ s�� \�!�$*@	�	���D�m���32p!�䉾 �>�ؤ��6r�����m!��-%�橢��E�~�$A,�$L�!�dA/:�$�����@�,\��!��Z<0PH�	�,�"�)P�jWY�!�D�.6
\��ɂ9]��%a�8!�(A�f*��&�i��%��Jk!�$A	v��頦|�n0�5%8+k!���y���Jqg�qk�i�D4{\!�D��25�g��QRF�#B�cT!�D	&}Z5 ��$F�$�Bbñ/!�$�D�9ڑ%I�`Ș� �T�%!�䟈
��t ̟�viӷ�� �!�$�r�&%J�`u�S7]&,0d"O.�G�R2�l�v�T�NY���b"O��{�珡g"�t
��ƒj$���"O"���.�D�$�a4E�L�a�g"OR����8}K$�1!*@�s�"Ol̂�dʩz���C���3G����"OZLؑ-��tH1m��`�P�[d"O� �`��d��;�4�E)��J�vpcA"O�x@��'q�ҍ�¥L:'��=��"OެSӎ�bfqI�D 7J'���"Od��׌t�qj#�Z�+P��T"O�{��F�v�˔Y�n'$�(�"O���6��A6	���N�D4��a"O�EXK�,��aᷭT�
�m��"O�)��K��J�fL��������2"O�xs�,K3-�|��wF͘(L>�!"O0Y���L&l��a�&X"2m�r"O�Y�B�U�
09R���7=pr"O��� M?}o��K�!����P�"OB����%{����H6f�i�"O��2fYR�t�t!׷ Vd��"Oh�� '0��Ƞ�j]�$�길E"Ox�5��m��(�G,��z��\��"OfiZ��3)��@��-�|l���#"O��i�aQ�D°*ؠ`����"O�`��k�L�}�'E�+�Sg"O�jB��S��!��o�)N
�k"O6 9�j�
��f� Q$�a�"O�h ��I��8�r�5�´�u"Oz0��O[�4W�|C�eO62 2!��"O���L/iy�®Ӎ�RU�@"O���rIQQ&���P�(��i"O�l�<|^�M'��:V��"O�Ip [�X& x��E�w�&"OX�l�,vM�%	���$\Jq�#"O����1X"�eOS�vq g"O
�q�?�����/;�����"O���J0]H	E��:y,0�@"Od-�0A�i�p�>T�"Oj�(R�̺{B	�`lޝ`,���"O��8�eH9v���d�)Rm �"O�퉧͐*ɌI��lM�g�J��"Oxy��ꐧ8P�������x�6�S"O:]{�ڼ3@���kҏ0� T��"O:��N@�=V*�� ��{�;�"Ozu�P�܆{v��)�H�~�h"OWʛF
�8��@�4��0�WG�M�<A�T6����a�1���J4��H�<1A�Ȅm��m��jْz+�`���m�<�r�&+��aX`���n=��F]^�<y��R�d���X��N ��#5JTV�<��(�q�؀�,ĩ*�(��NJ|�<��� �:�d����>F, ��2��u�<C���A�@aW�g�.��v��W�<��L�,bg�Ya�m��-�8�gNi�<���!zC����Q�*� �S�g�<� ��#)�$�����k�n��&�\�<��ڞ�[�SY~\	6
�Z�<�&" ?�\��lۛbq�@�u$�_�<��!V)@�B�J5�V�{�J���i�]�<�7.L�9F���*
�7�����_�<���O�
���'�� ��^�<!�=p�"�H%�S���$�]�<y�FY���ƃC�]R6�O�<�P�/:��de�S����t�K_�<a�d��a�0�zb��|Ti��ZW�<�Ul�cʔP( ��<A�#�z�<��Q�L!�=*�KM0�2q��j�t�<yS����a8 ��gA���t�Zo�<Y�Qa��#s��Wz��dd�<!��t�<9*U��?#DAl�<� 0��1 ��6���e�1�"O<Q���	PB�x;��®鎌c�"O�  �(.6#���D+�Z�n��s"O�\ȶ�ϖRӒ�`��1U=(��G"ON���   ���G�K��B�I�=� %�Ũ����:b$R b�B�	3���B3,�3zҦy�@MS�]|LB��(H�-����JJl5�%�+g�B�	���q�)�M���(H�h�$B�	2
���@m�b6T�E���0B䉽ݫM�=r-	B`������'�6�� fΓl�,�q����4�'�i�'����xؐ#�2�x��'��m!�D�7���q kG%���!	�'=�d`�e	8��Q��)Mu�'&
�K@,��e5jL��z���A�'�v�
�.ٗ�\ �2�۹F,"Ѻ�'�-pQ��v:l	Y�L���X�'����`��5o���hN9{�LX�'�n���KۃLF�dpC�J*	��#�'�X��
�W�RM"�>��|(	�'n�X�I�-ْXK���3w��<�	�'I���BjK�<�*�r�k%�`�C(D������rC��#���QCb��!&D����AM�.cxDY����b�"���"$D���֋h�n�ҷ/�0�����o D� ���$,\0�fK�;���cv�2D�P��ɓ.K��XRU������� �0D�8K�%�	8"~�K��_65�n����0D��Af��<Q�P["o��Q�\��%%0D�N}I�`s�fA#-�tqH3�*D��8��"��}H5���XI���)D�Ȋ'E^�V!����/h�N1P�`-D���T+Z>#}�qk؀U�.=
��+D�d ���		� �gY�Uz��;p7D��PF�O�[e��9�؈ �q���(D�$����:��cԬvM,�b�i"D�Hc ��bxS�d�?~z�� �� D���e_=g�H3#"Θc��lK�=D��+��@,-v��Jҭ$���`so;D�T�ǧ��X��	�v��j=D�\�rb�/8^��t�7��`Z7?D�D��D$T	�JL�"U��q�2(/D�� ��S��- !�J_�.ݖ�#�"OL��*E�)ƾ�x�k�3���C"O��*ϙ�����Jj2��"O��B��Z�浫��]�oDL�"O��_�h��'��~���FK�D!�Թx�T���i
#Q��L�n2!�$���ʍ��O�M~�3�͢h&!򄗙�4 ��Z65~�:��օT!��. *z��q��8J�!a��%!�dQDr��cn��d�0H�sH/�!�$�5 �L��ׂ@�	Ȓɜ��!�ć�q \��iO���)H�ȟ�!�wQ"})DjӠ*�X��!ኮD�!�$�,OP���A9p���&�ȇO!�ɪ=�n�������5�� ׁ!�!��˟�2���*�;W���pq�Q2m�!������p���f]��PAT�!�J
��Q9�-�!��� ��I�!�D�-S<�)EO��Q1��Fl!�4Y 0�w�'�����QL!�D�+� �;�o8����.ԒC!�Đ������Ա���r��=�!򤛓_��aprl:V�@�yE��1�!�$��,O��R�ɛK�xD�U�CN�!�T
WdV�[�Ƀ�_�z���Y�!�ċ�[�z����9f�B}A���+w!�D Xdse+_��hK%�3zp!�Acꨪ���6����$qOD|j�4�ا�^mH<�ea\�5s�\ G��x����,���fR�(��I����Bm��mg��fa�k%j�1��:(��ن��M�Vl3MV�HДm[�X5��0˝g�<����p�ղv�� D�Ub؟���s��1��J5;���RbÌ=s^\���I~���ҁM�)]���$$Ԥ*ڽ��Nk�i0�%H����ˊ,�J���3�f���N��V�d��\w"<�ȓ^���O�j����beY�"�j<�ēb�\�  �9w|tZ����c�Τ2��IX�O�`z��8ʂĬ?�T:��%OLGy�+P<YsR��E	�:G��)�̓(�y�&� V��m��@�#����yr�%i�\)�B)p�$}h����y�i��S$u���	kϚ���M���'��z��Z�j�����qk&� �G�y�I�S.�ȉR4xUL]�t�;�y�Ŏ!н��DR>r����yRkđYJA	�m���ЩcI��y2Lٽ���5c�_+ �Z�lҎ�yBB G�|�A�B)�t�o���y�F�8�ڠ #���=�����g��ē�p>)&MI�L���G�/)�(�#Yu؟(��C�~P�GV(�T��ǇuU�5��ẐTJ��%`�ZJ&�	�,u���|Y���@-[�%���	[y�.�"G"Op(����`�v����J:T��"O,�k�˚g_~������+AF���"O�1h��xIywJ�G*J}+@"O���&H�"��=�T	_�	Ft�X�"OV*��J�LJ9(dHV�~���7"O!���Ȭq��\I���}5(Х"O�y�d�	�"�00�B�/+<��"OR�����~\\�a��	xl�"O
0��k�CJ�9J��Z�thx���>|O� Ј���Î@��p��g?�d��
O 7���:����Ja���W8:�!�٘J� t	��VJ��C�ԬS}!�䆩`�0����K-L	 �
Uo!�D��c���光Cάpg�!d!��M�$�ȹ��7B9X�`H)q!�dޏ[ڴ�(��R"'�֫_!�D�5'��(WӁK&E*Gm� ;!�&B�� �6��7Ha3��
�l.!�#g~tPV��5
�A����R*!��-&�2������0�p��T�!���.`��5Eč|J����T�Y!�D�8`��dsF��	:LɈ��*\!�$���� �B>H�����D1N�!�DR�=*�j��]�O�h���m�  ��D~Ӹ�����}Z̵[��B� ��@�"O�UP�-C�\zh�'��S]L���'zў���̊cc>��@�%P<��74�;� �O��eH �q��%��s?a���?\��j��H�f<qqo^���B䉖4<ԙ�P��unlS��Ǡn&���0?Y'�� ��IG
(tJ�N��隣<�ɟ�IQpEE�vˌdh�%"7���"O�HY��=	_R5SAcZB1��� I���'_�&�	@��Ԑ�jD�F�^\��J��Aƌ���
d�'���1�ɕl-���U%%v�Ds�4�Pxr��W;B�:wPN;�8a�/���hOq�������$V ^e�r�	%@X�q�"OH��
�+y�DcЏUv��S����'b���,?y��S6W0� ��=Z��c6�f�<��ΠK1��h�߸3x��0&
a�'3ў�'un�� ��H�)���'d�B�$(p�d�7F	>k%�2� 9���'����D^+>����W:���@����a~r�'��7�%!
�I������ةZ!�$��6��g ھɺ��C!��m�az"��
>]�]x�o�u�v�pgAO;=�!�$�5'
s�f0��
9��1�x�E2�O��4e�&2pa��	-"�����\���	cQ���&�9,|���,@�}G!�Db��4$��s8V��Vk:7�џ�Gz�KL�p	P��`�Ѿ�����&	,PC�	k�4`�qEծ~W����P;���'�ў|�>�sJ�q��8�����i�,����`�<A@S)Y�!K��+*�=��I�r̓��=i���d;�H��BVCr�3m�c�'�ў�~�P��u�$7�\蕄M	#q�Gzb(/OD�ᇉ�����%) �-�Q"OD��mS'^��H4Oǎ8�`�"OBq�v���hӦ�S��D/iX=��"O��<x�ȩ@4��=Hv�"O��Yơ�ٍ�T@P[d��0E�8D�Hj�O��r`C�B�\8��;D�Њׄ�<~��0sÕ49�fHHw�&D���cX�@P��R�K�8P%��S�$D��(�
�3i�ֹ�f�:7��8�w�"D�쳇,��-�Y{'�Ƣp@���#=T���W�@�*�F5�W	E�dUG"O�h3��F.Uˎ�&�,G����""O�$����H�< "E�¾t��	;�"OH�zt��,f��Ѥc� ��"Op��B慞g���c^&����"O��P��
�΄sЁ�t��� "OP��&,�!y�P��Ϙ�0�S"O� |؀��.U ��F�tt���"O|���K��s�Z,°/yP��A"O�,��FW-^�I ��7HJ�	�"OT1JS�אL&�0���.w�X�X�"O"�B�((2,S����=�"ORiAa�
M\j!k��ć*=ʌ �"O�@X� ׮Ix� �Mͧ'd	r�*Ol�D/^j�x�2�a����'|�;u��\MJ�۳lԭ��1�'�L� ��vizJ2�>���
�'0��)vN�%@��"��u�y
�'1��ڣ@��g�4ى�ǉ
B�:AJ�'^�@�f��cCp�*d΍�'i��H�'�
�`�DA�ȓ@?/�]�
�' lbAg�%9Dn�`A��!�`�0
�'?*آ��L�s4z���/L}$�s
�'�@$Y#��p���Bc�%oQDx�	�'>j���!�w�)2���d����'yn�r��O�>����Kۻ]�y��'l�,c�M��I&��@��\�FC&<��'��͎q��(�%gV�8Kr���'�-�U��b���NC7;8"�	�')�ՠ��@z��.,���'($����|�T��O�(�-��'����.��	I0!��őUʨ��'��H�bIV�
��$� �ػ}����'����bT��ՙ�j��)B$��'��Q3'/_*2�&����ZX�<�	��u���i����1��I�<A%@�
�j�{3���[1+�F�<�>p��8!�
:ao��@l�g�<��$�>n�l�Pg���*�:�:Ll�<9�j߀0s�4��N�h5��0���l�<�"�=9��=ҰNG>�x)a�e�<Y�(K$)�Thrs��:(tHx�S��e�<���5p��D M 6Ȥ}��͐b�<ёi�3 �(I�1eZK�4J%�^�<����!f���pOȥ1.�|#��X�<aE��-weX�Q�ō)A�D�1�T�<	�Ł�q00�e&�-d)\T�ɑM�<�d�	&U��F�){"�y�X~�<�F�U2|���@�S"0‌�Po�<A��e�Fp�P�>l:@�Da�j�<�ף 
4 �1��5x�`�&�j�<y"�%:l��D�3[[L9�E�g�<��
�v^apF7g�(��`�<y�)L�����/{Bځw�Z\�<��b/J�85YW�.\�L%HvJS�<a�+�S�<izSݧ|��8���U�<!� Q�+��x�a%wm�pW�^X�<y�΁2�$x��K��\�(U`0��W�<�e`��[MACQ��m4,�����T�<	tŋlD]h��T\Ђ,�6�LR�<!%a� p�+� >�IiP��2A?!򤘱)�,%@�3RISAm?!�D�?�����ȗ_Č�eB�!���;R�%a�/�O���dA`#!��1ĮQyG�X;_#�BK+5x!� c'I���ݖC	.��'�#}�!��xb��6�ԕ}�`q��,Ì�!�dڃ^s"��S�0"��9��	ƎS�!�	��p�/5N��u���Y�a�!򤑏}�n��3��0��ژ{�!�<I��a�������Y� *�\�!�� l�'*G�;.T"���
Y���"O�����ѥ+�4�v �"W���"O�`�%ʑ*_n@�q�`�)H�E�'"O�T�s�Ȩ?P�u�ч�%���y"LF�5��QS�W�w:�y���yB�["N����cd7F�L�[ ��y�M˷2Sxeb��]�
�u�B ��y2`��Nq8��I�Ӝ�aKD��yB�Y�Yd�Ex��H/^-�f �yA���hЋ�C�(!�*���MSc�)��QڡM8b��J��8��!g4O4#=�F��yVI��N�8�Ԙ[��_e}�o1�O��`��Ű���#cO�H�H���>ɕ�)��F:(�	G�
z>i��M
�u�C�ɇ�갓i��|�\M	�l̈́��B�I1B$�A%OZ<pi�Sc�=\h!��e��y���,�&<jԤ�?}c�|[ō-D�0C�[3�<q�%8"\S��*D�t����jz��a��O
m����*D�T0�+�C�N���#�����7�*D�
!=)��X5��}U҅���(D�D��ˌgn>�a��	'Ѱ�h��%D�TXpa��y��ٙ!
�2cLܑ3�"D�0�/�"f�-��oZ�p���!D���,O2�ޱ����r��,�¢1D��0��S�Y~��� R>i��H	��.D��e��} |��b���<���1D���q%B�bQ$��@�
��Za�/D�$��J¾7�����
.k+����+��<Y�,�8J蹰c�8�@�b�	�V�<9�C�Jw��'�e�P��M�<I�&;1���C���dɠ��L�<����?UM�=+1mI*���8��}�<�E�4 �n�a`��>����v�<q��	� ���)E�S�P�L4���Sw�<)��!b��Mi$�P#A xq`�q�'W�?���`��i�B�;����8D��z�Ğ'h4�kN��L�t��,1D��� ��4��sa�ɱz�vq���;D��X��CM�=��͇]Aq+�%9}��'�t��4CK�T̄�!iҩh�V8��ē(9���p�ӝ ��y�&n�%X�C�I�/�dɑ���Y��1+�f"<e�1�S�4D@*ni��)���pC���c U�y�AE�2~��"�:<��3�nO��=E���$�PQB���=�J�#���@py�ȓ\Y�������8	Xp��AP�)�'&.���Ąc�"u�v�ُ�X+�8*k!�W*����KJ>��H� �A�(�!���(��a��a�:�"4�Q?!�D�>0��H"n�`�l������h6!��ÉC�\A��4l��y0.�)c1!�d�3]�"�𓢞�7��'�K�8!�D)e�h�Pq��06$
rLY(K?!���J�����i�+L� Qɢ�^�:�ab�O�Ѻ�/�=�����-�(1z�#"O�s��դ3˦=����y�z��	��?=�D��-7��땠�t���8�6D���ઑ�lHh�@��w��"#9D��+�h�9WlѺ��,��%j$,�Oz�Y��D����[� G� ��g6��H�=!ۓ"�0�hJ!!NP�as5JZ*E}�	Q��>�ȱ��p#�TY� ��۰�I	'D�h�ϧ �h�ĸ���@�d����ɅGtqO�3�)� <͈f @6B��`�q�#(_$�h4"O65����#v��b�A¨m0T�i�"Or��c�ӿ5j.�r�Ï1��ݓb"O��Iw`�7Y�	�m�*l��'�$!�O�Ѣ!��()�腣�L��u��"O�i��W/<XA�򎒓:��ȳ"O���w�O;�4��$(S+[��)���|b�)�Ӡ�n�*"�O3v���b�۶u��C�I����r%���Ԁ��X�^*qE{��9O ]���$ovh�y���)����W"OF�ĪE��(��Gb�����|2�'�N�"W�F�a�,-�A��=Q�B5��'��ɡ��a�bKH��H�����'��C �	lt<�O3y����'�d���EٸA)��!��3n���'\���0@��j��Ђ��.�5k�'
�y�/V�L��é��	`��Ó�hORi��CA�?2�y� A�(
��-S$"O�аA���0 �7拘"�J�Z�"O��ԥ	�ؠ���7l�ls"O�t`���2#��Q蒭�9� 5�p�dX�<)��R�)SJUҐ�cЪ}:V�%D��[�JM$���'n ��%���4�S��8"��RZ�)��z�H��I��'ۀ�"*�"CS�ȃ%�$�n�S	�'E@(���
�59��` "�H�+���'�S��1R�.�a�F�RlYb�RF�<��Jɥ~Ś%�/�����͖}�<�E1�޴��I$I4����G_�<A�e��xtX�s0K�S���D'�Z�'D�x�G�{B��F�Ô?-�}�� �=�y�ۄB7>�����p��Y/�y�G��v`H�υ~H�(�Wř��y�.M�1a��j��z_�}� �N:��xRÇ�G��4�bVA@���4���<�S��M;����R��D�g+&<H.�� T�<Y���b�)�fl�,V�e��n�Vyr�'�����¬w`�!�E�O�Vp3
�:��˓���'I͠bl��4k�c.�ȓC�����31PuԍӍr@�D{��i1Q?mbGdG?4Qx��vMD�c�2� # D��T�^"o����Û)�:E�T�1D���򄑾w�"�[Q#B	
*Q��.D�A��2>�Y���^#E�&9J�J0D�؉w#˙-��RW$[�K� �[�q��=E��4Z�^a�P�	~�Ak�͐e���[l@��G�ްu�G��Q�4��ȓhSf��nO�ZJd�קԋjQ�����V~b��/$�`�BP�
���\�C�!�y���ؠr�cD�\�6-��DG��ym�/H�]��M�}�B�����ybB�K�L�q$�4n�ѫݰf�!�d�>lvT`6h��׊H�!k�;rQ!��`}�F�Y#I*T�AN!���=D8��5Mͮ�<#&N724!�$ΛO�`\�1�U���M�-U[�!�$B6f���-J.E-ڜBF*Z�;T!�
V�؂��>���#w�G!�D�*(�py�X�+�@�[�m� K,!�C�>
Q���clYc[!�䇹S��P�3��I�t�X2�N�,!�R#!TƩJ���.VݠP:C�ŞS�!��r��P�4JF+ {�D	�Ý:i�!��I�<ؙ��<�V$؂�!nZ!�� �xx��܉a�v�P��7J���"O��1T�Ԇx��c񊛩^
�Y��"O��d��Z��I	�����hQ"O����ߣ~B�쐴��Zںa"�"Ob�ʥl�
����$U�|��y�"OP�A�p��2tf�~���A�"O<��(N�������,@�v"O�<��7`��E�t�&'��C"O������bTy�cj�����"O2}� �_0[���
ȕg��l�"Or�a�MH�E�2��c����"O�a@L� e�1�����>� �"O�B�(ҰL�T�����b�`���"O@�;�Ǩ=f�1C�_�k�I�3"O�5;���(fR4�1��)#�P�"O�t��Hӧr�(�L�'c�[2"Od�)"K�Cg�,K�H���"O���EN�E#�!�	�' ێ�E"O,��N�0�"(saÈ#p�@<ht"O�,���Vv��l�!٭O�8���"O:�!s%
�b�
/yެ�"�"O��d�3U���7�k��"v"O�t���Q;�=�r	�D�b"O�Mh�$^8%7�	���&<��Y�"O��x�Av�8�m	KՔ�0�"O��@f�\��1�Q��7��<[$"OF5��F���<�f��C�9�A"O�<r6�P�V��� �7J����f
�`�d�y5��+n<���\
5ԩB�%�Pv��eG�3!�D�-Ϡi� H*e�%B�2G!�d�)A*Hl "���l#(\�`�ϝU�!�D��uq�	�[%�iCe��!��ٯ.s�����^*M8�)17�
=�!�D�l�l��E�Q;(
��%�=w�!�S(7���Ѓ6jsıC����!�DCl�S���oy�!c��T'_�!�DF�{�r��+�	g�eR�&.&P!�E'�Ҹ��fɪAE� H$�N�!�V�*��B���#z�8!��r�!�ˬb��	�dO�@���EaG�3�!�$��H�8։z�=�JH�q!��
�&qf!b�E�^8\����X;Hg!�Ď�d��a��_*d�lPZ�AS!�DŹV��0�0G		*��CՄ���!�d�3*���&�:������O8F�!�G-V�T���O?dݎih�ȨC�!��� �\�@�J HZЭ3�-�!�D�\��P��$YH�}�"OS�Zp!�dA.V���FFְ><��I����Hg!�Đ� C@�:���Y�ĸ�A�!�ċ�C��%��ϓ[��� V9w�!�$��0/8�b`J��X&�E"���Qf�W� lO�9�A�E�k�@���y ��Z��'��ئꙿl�ba���C(hA#�B�XY���z�<a��M�l�����\�Uy��@d��'���ɧ@]�_�R1��	�7��f)Y@��(�G�͡Y�!�$Ți#�:S�*S��x����\����F��*0�t��>1���O�xfb��wl"m����1ɜ����'�4�@�!����ىCx�IJ�K*�J��+:C��W�?����4�̣@����#�'�����E6o�ԁ�lZ %�K>��Z'�c:O��y��H:Ȩ% Ba�=��݋C��1oθ� �2P&xUD��G�XC�	�}�>E1�!�6d(��RWH>&����i��Mö�EY���dQ�0M��Nc-(ϧC��%d6�t��T���sb��K1�S�
O>��&#р
�6��`�($`�z��M$<=ȰoB=9t�br��-��X�A�	�8�� c(%cO� ޡ@׃��69�Ճֹ,��� �'���@/���[�g���\��1�!\ J�yЎ�h{u� ����=�����v���:��򄀝��`JM*b�2��.-����Z�:�
N�YP���" �;`�)�.S��ĺU�ۃ?.kfl������0n������xbg�\[��`ץ��JǌeiR�
j{�(����uY��왔#Q�t�����ZR��@���Kń}Q¥��5W�.���bЧUFx51��P=	x���ўBI� �O]����ڒSXp� 4f^�k��(�!�J�%���Bo�I�vm�7<��P��TWj�HD�^�i��O؈3!g_  ���$M='KP�j��=%N\�Zu@9t�q�J�Nݪ�+"�E�T֨{���`tDUJu%ȑ~Y�0�a_�P�@}s���&SX�(�'��\�剨h㬈�v���J5��!*%2Е�F.J�j@�$�J�L(���\�k梨��d� �P�t��)�MSe���.i�[�`�	h��P���J�1&���'Ǿ�IΚ5y�\�@^��hdxchS�p��u��Ւ'�-�!	Ƈ4�2E9�*۶�@)iR 0�z@0�H�v��A�)���"�$�f�4`���X���x�4I �h��#aҪ9�芥�O����`��0a!Dc��1�p��� (���@��@?��cC�F;��$�r��	� }ԓ|��Т\�,۲�ɪF�N��g����~�%YM^%�B�=ɦq����uQ�]PĔ n*\�k�,���*U`�����[��N�[�X�;W��U
��A�.�?a��P�ENE:r�ayb��'��l���å9@�d*f�\[�R|J�t2AS�'p"={TP�F�0���j�$`��$Υe�b�����|�9$�W3K��:��<� a��a��|⌣��d��]vr�C�(�A��܃Y���W/5�l#*�ހs��!;��恀_h�Ҫ�:� ,��,\\\	)!�Ãa�Kw��) {ayr��HPFN�UM��ukJ���C������-Q%�ʄAH�$��ǚ!G��Q3@��y��xD�#[{�'�xU�1`J�F ���C�F�(�sJ<�! ��d��}�W�-O2pq ����Ip(^xG���dÏ.��mIB$��*��(G��k<��ڱ��"K�uҲo�QvQ�剃|R�$DJ9��S�H��$3J�2%ɒ�)D��rRIH��e!� ӓ.��R������ �*	��T��VH�X��)ܨNt�� cAn(<9�-��zo���p`�<A� �Q��А��WF����/���>�l��1��؋�A���9(�C5�c#C����w�!AE�az�h9���aáb� �gN�8c�}y�+�.g�$��%a�@�͓6����¦1]�mj��ՙ?l�AC��)h�O@�z��&I��8���5���[��Z�Lw����� q(u�7d��"������/|7-�7K��P�$W�F�<�YF�R�T2�A�DɖfAlYԩRf�"-��	�ɨX0@�\+,�J8��5]8��lʇi҉��ŀ{��e����ƶdH��iW��@oֵ�M�� �3)AT��w�̌2�iB��B(Y4Υ0W5$�k@c̽4ht$�!��4o �z4iϳ=��s�ǃ ��f!]�.�a6`�}i���Ź8d�,�E�a`��! d�"�ЂF �8�6�6�*\O��9�-�<��a٢^q���h��,0bF<��"�;Dn
��E���.$Y(�#ܡ0
��r�!X�~�i��>�O���'��)��@(�/�VTV0X��d�USD8 ���}�֕���&������ ������'a8l���4�"(�Ř�5˞Djv� �ܶ�#��JS���D
�Da�i��n���X�Œ�a�\#�FX%M�X,�jՀ=[2�Sơ�4��$�U�����^3
T�)�$
�Q��ң�STH2��gAE�y��9@��ciɩR\�j�L[�[�&u�c�z}�&�c��G���&�ʉ�D��)`I֍�t�$��7��(x�D�D�٘(��q�W��|�����e`�@vG
�/TA.�� H��΄6l����//9thj�@N� ��d #��(X��ŚB�ƥ@�0b*0a��&���7O'{�|A:m��=�v�%�:o������{�\��F2�������$�KR0jΟ����$��@� Dġ3���@q�/OO��O3Jo��r��uF��#R!���$��,N)��Tz:>1��N��Ѳi���SG�E4��QiMzb|�K�f���$�
�νx	�fޕk��x�j3�Ӂ� ѩb�CT$�!֨7�0x0��*�:pP��a�.��T�r}��哆�fc�.T~�H�E�D�`!���PF|���k���#�h�o0h�"�_�ͅT�j�� T�̈�\TĪU�&I�Т%(��F&�0�G�NI#��,Y��8Ԃ�
�NpIT�t�Ii�4��� �'Y�8aY6��	c��+��h	�e�5L��f�p�hF��n�.����&[�6}aF�`� �,C��E���m<�}�S���V*�Q+�
�%Jp���$>nXS���uX���A��nM�m�.�$2V �)��,j�5��j
#��qTd{� =L�F`��F�!g�.����,�T�eh�{ 9��ɄD �Dlɿ
���'F$à����}�d�ӪK�m_zp���[�+V~D���;�����Ƥæ=�EG�{�v����-l[r`�ѧF5y>�XY�fE�G�
mp�Ν!��'�0�q�.P�:?��a��2 L���B�s����C=Jf:�BW(˨A.�Y�CN�yL���4�/p���J�R�U8�����Hd8�RwhK�@*�I��x28;���� :��erÑ4V�`��(�/G��5ʃ�Q= m+��ֻ=��*��~��Ț�S���+_�L�g�Ǚ1�J`R�h��b�k[(g���xC�S�M��y��i5>����	Oh�#�5U`�(�&C��No���A$=m$��6}�]�a�qѢ�bƐ����m�=Ƭm�#%L9\D��v�[
Pt�H#��Vx����Ux�|KPS;]�\�`bT�[!b�1sfM:����)\���"G7mȈqi?K�t��"��],~�I���O���O��DP��ڥR�Ha�U=����!��5���1î��&}<���M��/_��)S
_6�)r�CvtA���u���U��a2���Exl�h�ߜ]�z4P�'r�w����=�W/��}?�U�B�Y�_�`�3&�z��գc��-��Y�%L�=7nʽ��O^�x7�A�R:�d�{�&܋y���� &lB�D�@�J!����S�j���� uJ�'F�z���2i���a pQ�b��<�@�&�g^�Q��&(�x��U1m����Pc�m`�)j�PJ��*'ʑP�H�5&%��@����jPrgB�1�)A��hM�E��?U������'Epd��֧�&_T��3�	:k�ar4��蚒_�L��`��|���H�
��'�2e��@�.��O(�y���@Z�D��b�C*S*B��D�اVp�%��);p 9�Z�n�Z�qAGO(0J�]�]�x�uj�9pT�i��'d��u��5oN����:A�0Qp�@�YX�\#FU9���{�����.*��A�0i 6A�\� \��k���b�(���Cf�p�
O*��=(3.��q#�W���PiN�X! ���Cé9|�ꊂ��Ȫ5�@?/86��>�e���\��FaN�d���˝+by��˓{�`�ك�W�P��(�+W�Ҵ�;���Ux�M��)�"�!ª�;&� �y��'�TŊ%�"s�~���N�H�Z�L<yu R������S)_~�8 �.�S
2�I5�?�A�N#F��@`w	�2�� b�.D��ZD����*�)�NG�p�Ό�'+@>]��KU�j�`�Mo}bb?�"c[��y�+ԊZ��y�k�f���ϋ��x�B¹ Ѱ	�`bV�^�K+�\t�"Mڂ	/p���9c��BpeƸ#֠#>ac蝀G���*&�Y(7�60Ri|x��2f��4�$1h��ѿ1��5���!L ><1D
�?%#
5@��ܕ*��<�dbCS���x���"=����$���!�a�&��ګ}����G�T��m�*Ki���!?.A������!w,	��OP@>PB�
N�G�X�N�|�����4%ڍxPA3���(�;>�ASB�<��2Bט (�'XDĉ���*`D���ӳ>�ֈq�'p�XJvAX�y
�x*Va�(v�$�a
%d���w J$e��
�G����Mr�9�!|��t�ڻZ�$���n�@����ɵu��m��I��&��U�äC,�@c��	y�)zt��L�B!�0!pA��s�LQ��%<�$�a$&��A��%�@����6�FQ��n/t�T�X�=�Ȕ!˟xT@���ANX�(G`P�bdΌ)�"O
}Z�
�QR��mF?cVft#$O�<a����p�s�E�'5豟�I��)M�<9Vc�:o� ���Am<(�0�\p}�)§8�����h�p<zУ��?p�2�,@	~�&����  2���0c�)w���W�ɀfjsD��@42Ƅ�\�xO��1������M�H�0�b`�.�%beÍt̡ͪv�  ����P`�3#U2�X���\X�P�
��,
�b�A�#I�5\�$�4�B�Ґn
�:�� f�i��@2*v,9�ƁA��T����U3�A˷KR��y2,�^Fn	Re�IK�����&�
ȴ�ՄףRY������[l@��P�\Ej�'�Ԙ��1�h)��¥T*m��Iݤ�L�uOe
 I[��<�C��R��D��CɆ=��)X�KR��2��,U<�b�+@�[�*�Ph3��/^hq�T��)x4����1��DT�+~:=�!H��<��5��7y�B�k�c�
T�P��
	/}�Y��
;r3ԍ����9����dν*���#��+Pe8���Ν"1O<���$���K��?	�Z�撳~P��y��<+��EI��W�wDn\3��:^W\x�6"O��� M%D�\8Rj�9n��SB!�<�zm:\�hP��k��]e�a�VK����[8&�E+�
�����;W����Ŏ'f!�d 7K�M�V�҃$���Wi�to\-:3�Yl�8�J�(x�8�0&!4L�a��i #��oS'��dJ9��9��H/)���Qa�1Y�azb$�I����@#Y/c\�M�p��&+L�X�L[�X��0�5�Ře��Q�2$I�v��i���0=��EW��ȼ�'��&q�@vs�p�L	Cƥ�0iQj1�!*�{�TXzg��2gZӆ���H j �N��Y�`�6��(�ȓc��M�P�.�D��uHԞk���p�.�Z&�
�*�Z�R���e��i�0�n�T7�yw��^ƹ�S�S��Bq� ���y�˄
�&����T@��D�W��P��7n��}�^}h��[�N�jq��K�|�0�L��'�����/�m�T)����R0jQ�ӓh��p'���>ͪF�߮�ԉ(E����\!����&	]�%��]	Q��P��)=�h���iJl*4��/Ҋm�0�N�Rخc�h�p��VѼ��6�G"A5v��BmX'����-ڌhHl�IDh��TS�u�Ѭ�+Jr��be�%D��0����a�f/�AЀ�E�ÍPB�Q��7k�jA�Q��[a8� EAD���'Yg4�F@�*�"Y�X�0A�K��B䉷k��%��Cۺ/�0����զ{�.u��O\2?���"ȓ;L�Xe���r��3�Ln��O sH�8l���'�	n����'r���V١%s��DxCc6frR�q+�1��d�06�ik6�';�AC��!a�֤s��P$Z�J��W�rУ��C�O��)E,��uH �r)&8N(��'�a�䗵D@�S�%�,X�U`�'�,��aJ����i� :ް`,Oh4��S�? Hh㕈�!^����Û=���"O��pD,�
|������V�7�E��"O:�K`�ޅ�|*'��0v"OB��3��0�N�!�A�*P@��"Oȱ`�e��3G�M2�$�z�Xҡ<J8�|�'�)b�$�92�ʽ &'�;k�(K�'D�AN�`��zw��F�	�'t +��Z���g�>
�ܫ�'�4Aw+��!D�*�6,2���'pH���Պ(3N����/�ָ`�'RX��l�4��сd�L�D�����ۙܦ�F��Bŝ�%/����5�f'�.�(L��`.��Qb�Q�DJ`/
Z�"��	d��YS+'�&YҒ[�!sP݆ȓ�vA���0w,�c	��6�$��C�<h C�A�ftB�ȕP* �ȓ{�&Y¢���u�`&¼:�ȓ/w�}��K�?�,s�]�Y�L��~"�ӵƊ�F�2AɆ��0G	���+�*126"��f�����F;Gw� ��3�z@R�ɑ������[�8U��`:h�2�L�dݩWNB �z���4��X�iS�By�z E��M8��|�s�f�B��u���V���ȓR�b3�ɞ T��B/��Ȅȓ}f������N �S�G�4�ȓCU|�8�Z �F�{0�4
w5�����z1��hT31KL?+�t4��G�U��٩wU���5G*j	��2���+v����	�0Y�V���K���C� �5(y�A�-u�I�ȓ�� ���/N���n���ȓL�@ـ�N�,e�QæU&X0A��'ż鳗F��v/\���˝H��e�ȓ����K
IPmH��Ԇ�w�l�
Ԃ@6x��#�K�����ȓ'��1�uDJ�shT�D̫0��	�ȓ&�� T盨4����� ����h\�6�ܷhZڵk>N�]�ȓ�@Ix$a�?H�>`seaP B�h�ȓ�q�!���#�ə=HD~L��Z�b�#�f�$)�ܕ��D"S�M�ȓ<r�� ����5�O�b�nX�ȓ\�W��]��zWc˚
_�݅�6��!q3��>�D�JG�M�F9�P�ȓVbt8���]|.�ڒmh��q��{��L�Ä�L5���ǉ�i��ȓKX�#P!�?��1:t�
<X^hX�ȓpHй�셒`<@�I�.�<m����uQ.�)���=d��2���0��|��0h e��MLH|�1�D� �4��H��[@����B�]g�ٸ��P XnT��ȓ	�(�d�W:I2&�`�f�	= ��ȓf��e��#@�ݠw�<&�l<���B5�E�v�� *���<��ȓU�p4����dlp���7��5�'��(s�#�7��=5j<R�P��s��+��<���O8����L�z:F�� O��L�% �-n5�"J�!5!򤋍^ N ��<]&�}K����B*��k���� p�/�'G���h��E�<�D�"t��Ģɇ�o�z,�aɘq'��*"�� ��%��o��E)�̯��d9�g?ɱ���S��p1De�/74�#3�Ti��������^�� �#̖&x���qϘt�t(Wf�2>�dq� L���p�-�@X�h���S�ň�坅0L���(��]	4D�+���<)��_�
Z�A���;e�@���=� l�F�T5#�xAg�ǅc������vH<) F;#Y�h�	(�a�4��dN�+��iCd���E�.��Lh���pM�(�Vdf>���Ɋ�y!U�;��&��T�rG9�Px�J��[%�����($�]��CKD{��ʅB�)~ L���ٴk=�hx�盫X"��� *'�U���xmۧo0��E'�Z�  	� ��0<�! O�9���� �������5{�x�	M�'?^����+=Dh����d�LI���<l���c��'�.RՏE9ޘEw�]�v�����O�=�R�]9M��=;����C��hg��1-�ؑ�$.�2Q��y�ʐ#F���B�%.��C4���<1��r)<����q4���gH�>[��KW������s1����də<]��[g¿z�
�)Gc�?zB���e��� O��=�6��5 JSu&]��8'u�z2���K�H}!fNIc���n	��i$��^�H��bIN[���И@M���u��;/���U�ъ��QDd�]��'[Thk�i k�
)(㮗dD�<��y�Η�fB�$�ׅ������5�`56��y\DL3 '�$w]�4�%�=/$�h��k�M�u
'�� \�D���"H������4	���h��ы!?�,���A1t�`]�P�uM� �C	�f0+�����0&2��@@���F�P#%�����9(
,<#ҀI2A��8
�'$��yS�.Z�SV*19f"x�S H2��!aT=d�� ���:��� �N��
O�=o0\����4��@`�
2̪���O�"oޙ��$,O�Y���@ȐkAŋC�ӡ�UW���p��ЧW�)�Hȉ8P@��X��
m".Y�x����#��P��� Q(&��g�<�P��X�R2�p��C
z�>�%�lȁ���IZ#�$�$�g#�
H(�O�0ƬMB E�[�bxF��j@D�%/L�yNX���e}(� !��5Z�����B�5*A�%z�	����T5Y��� �h!b��w���a�ՒA�`�4,F.ؘ�N��5$ �R2�@�V��|���8d�ĵ��O��Xb�'��0sb�	(u :f�?B�9p�M1#����灣a�����"= �9FD���8�,�x1� ��@AeI�9�ƫ@�r���ƪ`����� [bX�<���P�
��c	@5B�f)�A�<%|�:��O�� ��`,�'"�+��
,)�tzsGE�X*���A�q�ɞ8��d�&O��0�F�K1#�#�8O��(�b�B?>]����*��H�F�w&x!ԣS9z��Ia�T�3���z7-r�@O�*�RuZ��+pܬ�h�'�f�ayb䏱�"d���F~��IB� ]O�<��k�$oEr`�g���"/x)�ՄN3
�4P�fd��x��m�/���	�]�y�n���M!k��,Hu�76M�}��dĸ���:��lI V����q��
�z�*�Ï��5f����ۦ]�S�\$'t�)�B�/v.�E��8�Y�(�2i����Vhܵ{r�R�'��QT.Z�:��xQ 	!A\,Kwdͼ#��-�3B�9/�f��ǅ��<)�Oސ=(*����8|S6 3��?$�����"��l�H���*��pX'� FNqO<���萢$�vQ{�B�@�J�8�g?�
��wӜ�$�^�s?d�K��`�b#��h�b�t0X��+�c����ɇnr�Ҧ��7s���ʅ#A8d�V�@�h'����Y<�F���i}�V�i`�4���T��M�@�Z���b�W7δ)�ON�#R��+=$�4�vBO" ��̛'h�5FZ@���n.�:��H�{���HA
j�RP��B@ 5ɗ��l�
��6��F�F�y牋m�FtH��ZXdZd�R��Y�����.7&$Xq%�IW�4�WI��|dAw%T#T�J'ˢ{�� ���%u^T�@ҡ�*#~���)�sz}j�ŕ��ē}�nQ@cm��Z/�0JSb�A�H�<Y�G�E�|�7I׆3�@͑�"�!2*h�h$@H7z�pm��"͌l?~a�~�B�P�MT�{%��V�D�x��Ǭ���<iq3{ȵ��!��/hj8�Qc�1���Ag�x4���G!>�9��>��)�28����؊YӜ���`֚j��if'_�a^]@�L;D� �(��_x��Qaܜ#�z-Xq��*�ɏ��4�Ջ�j`� ��������\�������@����i|���8(�az�B�=�hE7�ݗX��DX�ɰ;jp��׬�~�j�Hf�Y�GP����}�ԕ��M�b{����2>gn��'=��hH~5z�M� -R7��d|c�$rW!Vaq%�vD�!J�H��h��rr- �O�Ƞ�,N��@3��%)��I�AI��v���6�X���ޤWO�ea�� ~�*Ub ���qz�a%���A-~,��k��iF�C��P	Ĳi�jq�D�L
w����%{7�R��Y�Vcf͇j������@�*ѫ�GW��c��׳��m�'�Eh���Э�kيK�4�AƋ$;��B�l[����DNR>#n�x�#*�s�T�*�萃KV* �	ʉ�d�:DĔ�U쀋.<���E�,G�h�tI�X�T�֣_$I����4�tl��τ�d4�a�$	�%�x�G�[�D�[��if�l�`)�!jH�v��Tz�V���� Qqb�n�(�)UgP�nk�H� ��&dT�O�W}�fǭHu�9�P��Z�DM��/Ѭl�xĪg�"	6����[�z�J�@0"�-W�^u�WϚ�ʮ)�w)�� +��rE�Ux���A�ۑy�@�PB-U�Ta�7/Z��� 1)C�R�vY�Р�:<�a{bjүi�GхDk@ ������e#�%�)s�P��nO#~R*�b�ə�6Q�ba	4N��$�g%�)��YKS�Q�t�C��;GAԦP}, r !	8��i�=� ��^�dH�������
d��O-qW4(�ӯ�|\�e���t̜h�!�rJBH�ץܶ�X��`�L�wp���I�E�j�C�"	��`�-�rOV)d��%�$��a���PgD�0B�p���	 ��i��%��(M��(i«�"y�XlY�'ިR�!��­<�V��%��D�d�s���h{0�C�U_T�@4-�`g���F��-<�N����J�B�z��'h�Y�	�"WT�5�Āe�X6�E	iraz�.Df�N4Sŷ>�~
� �:�� =D�ޤ�4�b��(�� .4����L�M܆yr?1�`ߡ^`Ly�y G<G)��;q-��j��+�ߨ��k��un�+\l�d��=ڸ���8T��ڥ �=D���8V�ޜ
j7Ѫ@K
|��j�āЦ}x�"��'Sn]PVk�<Ps�\R C E�)����b�8�{���R����}Ƙ�C�_ꕂ#5�|8���).�:4;d
�0a�(����2�I�@J%�Px حM���ӱC�s��JU��3E2��DN??��`'��#R^��M�I���G98֑Kרt��X#�S�y'
�;���M�&q Æ�|��}�
�L��Q��L����pEEp����A�3��-�W�L5tR����L#�X�+� |��L3pg��p@�@�ޅ�<y`�'J"u�P����coO(\HrK<)��~�eB�Na�x�&AϴZ1hG�^�V0����I%o�X��Q�Mz�=��Ā*�ɸBT�`��l*�h��'�88{�+�$��*�i�6J��qhB0`�,�1��O)T����dN2�0([�K�\��f�e7mH�,V4���k �B�̊����/b+fC�:�� ����o��#��G&,dA��#��t h�f޹e�b�2��?��HW��`��'>x��n�"����"�\.8Č
���J2ay��8_y*�a�Z�+�z0 ��U-C٠[��E9y�h��C�#���Z$-�F;Z���N;
f�R5�XZ2��>(�'���HW�bpJ��![�،��k
�A�f�'.��E�3�O���/8��Z3d�K�<!��V�@C,�Q��[@��B��R�WPx�`�$��ʆ}��DM-u)2��~
ë݋N��$ԄTG𝰆EM4*�<� ��H�!�1~ P�0$�"��{��8#��
�g�J�U��
8T�1��(3x.pE|"D�A�� {acN,^�� �aږ��<iQ�έ]�$ؠ�MJ@hDK� }J��b㏁h|��U��J��%��DI��0?���P8�`p��FT��$Z�#o�U��8wC�-���C�ǔLg�ux���b���-oN}h$���S"�f+���y"�O�c�^%�')F�T����'�N;�P�J1z�|(3��j|rl���4�۞�*牁w��u
�,��D�p��Y&= lB≤rz[�������hLsz�� �W�!����a˛9m��hH��t5��d��f�8�qAN0Ⱦ���_ayc#i�MA���  �pڲ! `�!h��0�D��c��i�r$����Z����C�����F݌9�'3@ٱ���9>lL;��\;ݦAȦ�՝[f��'<�œs H�a�pr�۹0B^���m��aS����&���0�Ż�@ȟ12M�A�P�di�(��~�'?���?O.�I�_ɰ�8�GF�2���O�3eb̳<ʔ�ϝo�6�
�FS%�s1C��6��Ո�-EI~�Bq�'��(�t@Ֆ���)P�]�DD�
˓,D��ǃ�#Q����%[� �6�ʳ_p7�%���#���7#/?}��W#�20�a|"N��vT�%A�Ӑ9�jt�懗�ē w�ɠ�ƌ�) ��� �lY�%S�;�bd1�fG���f��
�� G�26��dܹ�y���-��a��ehB ;��ٶ�(��K;7�����3��U+�)�,���d$~)�62�F���A��y{l��'��6 �T�&Opu�0nˀ<�.�s�垏0�"��#��s��S���/��w���a��r\�	š^�*�qOL�QhX~�̠X@B�'+X���#�'�ʰh0b%-U����-��d<qP�F��xH�"�M����"m��L��)D�̅(n���'u�����7���b�k��oS(��y��1lZ>���gQs�d!ӎ\��p$��哎r�Ё,Յf��$��B���J�f��y4o$��醆 1�$i6�C��D8�Ӎn�t\`��`L��`č΅0h(�Ο��S8ﾁ d��5A&t��T�V��t}Z�"O씲��ڃ+�&I����g���n��?��%��jӖ?�\�+I�F�脂��-�8u�s���;|��18Yڽ����r�az��/��40-��`����)9m�#���9/��P���E��]�#&й%�rtуb�0=ٱ��g�Nek���m�FH)���`�l�JTaEc#t2IK5 �䈹��EU2*)��GR�x��8j��+�Hq�H�z��l��0ݢ�+!��5�x�h�AI2��Ic�<m����	c�xhS��6Ѵ�A�_�d���y���z,�������'|tm�W���y���:�G'�3�T���Q�$���3`�8y~��I o��KY����ӗ��0��'��I"Ɵ�v�6��o˻6;���	�q�h����BL��E��y|��a��O�h����+m�Ԩ����.���G	?�)��	�ag�С�@��±��D�b����$؏@��S�F�)(( ���L��p	 ;`e�,c�����	���&\lBك	=D�@Y���#(�p�'�
?$��r��vM&!�b�ˆ~��c��ؠ$U�Xi�#��'&S���D!�i�Q�d�h,�����~k�B�I6A�f�Hj�C�F��㦂�_n�h���:�P�s��� ���uG
�F����?�q˛�3�`8s���b��p��{"�E?bi �+-n�]����o�h�q�fӺ��J�7ONU���ka|
� L�Y��6bR��dB'/��4qv�I&̪����9�H���[ B�B	@8��-� (#�"Of1A���>6|ԸRd�����c"Ox<B%� �_n A�U�# ��Q�"O�q���N��\3��_.b���"O�hs�KY'
n0�'��{m��RF"O�\����+����F	*mXi�P"O��ĩQS�l0��� aP:�Y�"O$����Z�:0��($Qź�"O(�3�hM9F�I3����37"O�!(�U�.H��� �>�i��"ON���1�����`�`(�3��*D�<�2$�4Yg�$ҧL;����C)D�<ˠ)C�=u��t�Q J4��'D�hsw��N�<2��[U�&dy��"D�0�4	>r�ة]�{;B���,'D�|�n��Vw���1��&���v�8D�,�!A�Hh��(q�������6D��(�*�$R�6��	�[��5�.D���EzN@�o��p؆���-D�j��;Ԡ�y�Aej����-D��Xq�ۆrZJTy悜O>�J��,D�ؙ6J�d����݄P�H�b�'D��Q���"�TEB!�!#����1D$D�P�o�1|�$P�ϙ:4��i"bh%D�p��7�ݠ��&M���`�>D�T20�I�=R2���(Ԙ�&��J?D��*�L�a{��`L�}�"\;��!D���IN�s[��VA	�g1؋2�#D���@�e�ܵ�V.�+�ʩ�ǥ,D��@rC�!�n��w#P�Bv�y���,D�,���;iU�6�"x���[¤+D��hV�5Q %�3E�B.���B�I�	n��w*�,_���B����n/(C�:�ʠ��T+������\{�C�+��gdY
F^A�GC���t���"vI�����w���ɏf]�I���=zdʸ�w!.D�H��(��)N	ZĨ�i_�X�b)D��;Ią^X`𙳌�]�6t9�.)D���7ؔ�(SEW�U�l��i%D�L�Blܓ1��ڒb�m%��SH.D��⤞��y�Wٓ���F.:�k���	s���D^�8c����Zn�O� Γ2�ܢ}z�fӜ�a@IU�y�Nl0b�Y�Ph-��W�0���R�J~2��y��  �,�A좤AT��ۦ��'���Ԟ����Ӻ�h�';7|Ey���4<4�E�X}�*�S��dW��~K��H� r&����V�=������OD�>�'���+�
�� ��'�'L۴��O`�I6����'>�p�Rj��(Rɏ�J#b�@F�O*ᨦ��?�$���~B�k*>*"A���CFq��J�T�d�4�곲ivRy +O�˧���.���D�}0,���)i���?x�L6-CEQT���'�����AE�T�4��Hp�U�Zf1!J)��@3Ș�<��EVӦE�	����П����W��( *ڕ���T�	�Z������'+�'a���-w̨l��<4�FM��~�.��=��/D>A �	Ƙ�F���3&Va�
<�I�&Ti����]�G���ÎɑEG��k�=��I�&F9�&(?�e�^�O,BuB�M_|	��?�6�k��$��A���QyҎ9��H��ӄo�,DQ�߯o�J�i�j�+:I��Z�xϓ���4��I/]f��WϚ�@�`� �Tq��Fz�O�Zb��Yg���L��i�A�3]��.D�3S蟐NIj�R7��Dq.)ZC#,D��B2�z��d�n\���*��&D�d��΀=Y� SoY>&��p�f%D�04B�X�^�1�aE�Ta��$D�� 4TXc��[�,��u�M�" ��"O���!O=]R�iQ��s0��"OH�vf�C�� ��I �93�y�"O�8#�.�yXHM�sO%�L�u"O�A� m$��V
Ǉh.�}a�"O��1uaŠ\�096�R0p)>��"O�I�/����}�'�.'�x�"O�m����R2	a*Tr7���d"O�e�DO�2<��L�F��/����"O���	�,��I$Ȟ�P�@��B"O1���	O�p�����:{��" "OV�c��%3� ���j��u�t-y�"O����P�K���Q	2z�
u��"OR=�u���,��r����`؁"OM����u��u�� G�fqx"O�	�\�8�f�l�(9��>w�!�L>V�n��s'��ZZ`9�T$D��!�C�F=[�EĿX���p�œ�!�d[a>���!�&<�~D`�#��!���@A���\ P�Yx!�Dԣ}�<i�����a�t-��a�r!��%	����C��o����� U�l]!�Ć�;p��{e�3lV�Җ��z�!�dP���C�`�?;,��c#U$r�!�$�7`�@�yE��=!���e��uk!�d̂)и�+�8����ć��_�!���=C^1����x�KF�t>!�+	�d[NI��Z�+v�4X!�d0,Y[�d���x#ײ>�!��O�Q�U䃲rr����l���!�$�:�RHAc��&*_ � �
ɕ-�!��I2���)�p?(�"f�Ӟn!�DO*_β8xG��G9��	E��fP!�$��u@4�v��8(5�P�W�B:!�טb0�0�'J���5�ՃD!��G)� "3`�&f��컱��=X!�_�s� �b%ِV��p`6M�:0�!�$ӵ6S�����#����lӊz�!�dٸVT{�$���.�'���!�d�B�l8���.���N�Y�!�׉CΠH��͋�'�$���ϗ0t!�I�r �ɉF�R�'2l0�&����!��^��еۓ#	�xMv���BLy!��y�|XT)�b��������O�!�d��>18#�4^����AEʰ1�!���4Xj��r�]�]�>� eC�.H�!��U;S�J�C�K b���ԋ�"/�!�䗮>��]I�Ó��n Yt��|-!�J"Y�0Q�	��` c�*��i!��ƶ/z^����?�4P��	.(!�D��
�(��F��2��wi �!�$_�k��񴢅4W�V܈A�ё�!�I�{:���&�,x�
�M;�!�$� ����Z��p�R�9w�!� ^CN�[��N�*����#�!��.l�\��R&P�i� ��c$�b�!�D^�S�j\�DߚP�`=y�"O�+�!�\�EM����-��$\  �!��!��WSd	r2�]94��|;U���d�!�P�QJ��r�9�bQ����dy!����x��V�u�@	�ƛ*pw!�d�^߄=�c fX5P@�܌u�!��<:Y���W��[�|��#��
�'�����/B�
�8�k���*��#
��� T`6��)}�4tQ�'? ���"O��z'BIT.(
��K O��7"Ol��g��~�"yrO����H"Of�[����9n��t^�,��J���y�I�9�a3-ϒvH���˛��y��\�h#r� � ��t��  �A5�y�L�@��0AE�YN�j�J׍�y2����qQ�ݶ}���"R�͗�y�j	lE�=���*} rE���,�y�#\�#I���!��}VV�2��Ԯ�yR%K���7���a#h�S`��y��D�d����S�(D���K�y҆L�!"�������5�����y"Y�&��q ťqa�5���4�yr��"�L��j[��a� �� �yr�� A����lW�Xh`���<�y�o:r����H
T���vh��yB��87��(�!$�Q��u8�y"d����02��r�� �`���yr�єeѸ�����6Ȑ@`N����wX�����PюQ��ɳ:*Q��8D��)uȘz�r����,��a�8D��H�ˡm�*���I�=����5D��&�TGLȡ%��^���I�-5D��Y`%1%z�@��	�@�x�"��2D�Ĳ�#1v(}�P��>q����#D��@q �n����)*����*OP¥��������MV�`;�"O4)5jT�����ը�-t4$bc"O�j%�Զ1pp���+����"O���ʋTz~�)���m�"O��K��[�lh��f�;o�*p��"O��Ss��Ȑ̚�׀R��W"O�t�W�R�_��=���-D�a�<Ც��I�q�g�N�f���U�JD�<�����Zu�x8��д"H�\�FōC�<�q�L�&;1��pn��;�CYx�<!�jS�"��Ă�g�]�y{�cr�<Ie�S��:��P�$��N@g�<!��]�yR���F �^���:U�Pf�<�V��ԜBq�Z$;�4ᒢe�Y�<ـN���y7Dݦ%�@!�Ca'D�|���0HH�K�"��"�8��e�/D����`��Q��S�KӅH$=��:D��#s���k���m��l+�� #"D��ېGT�;t�r�/�����r��3D�4ktc�6tD�œ�J�d��[��.D�tJ���lRr�h@K�X��C?D�8�b���V����G�=��xJ��;D�di��Ϗ!f�r�ƀo,�9��/$D�@��"�~�kTo�5�4	r�?D�h�$��_2V�K�a��3����*D����J5X|�AD��N�Z�/)D��V� ,����
��?�@�1�e%D���ƀ � ����I�,��&#D�0�3��g��i��ثFl��z�6D�d{6+B&,�|��
�4I��z�b4D��a4�ė6�f�3�x����'.D�x��m[�j�I:"qa�i0D���ů�ܥ��L4s��bA.D����g�'��	�&�G��,BF� D�h1�n�w<�e&��]��=D� q��6|�C���o$�;��;D���`e�&~'ba�!o� ��PA��=D�� H����8��v×�$M((�"O�HVD+<���Ѓ��A3�S�"O�IC�n+?d��Q�	Xx�NY�&"O����i�%z��ͣN  霤�"O���d���KÈ�cV�4DG�HY�"O�x	��ǁ%ΜȺ��06=܄��"O<�"��1�ܘ۱Aނ.7L�R"Op#�h��mq�k�@IB"O�y�Ą�6r�=��L�p,��r"O��vj��l)�� +b���1�"O���qk
�]���R� E�i��"O.I�":�H�q����9څ"O���n�e�
�ʦ L&��yu"O�� 6�ѝ�R�*J"}�r�" "OH9�!K�L@�g�#$*꽉�"O4�$A\V��p�$�'
P�`�"O~��4��bx�D��#6F$Z���"O�,���J�2��-Cu�I�g����"O�Hh�@�,j4�`)�*��)A⼲!"O�ejǠ�}ܶ)����P^��{6"O��E@�`���p�?E �t"O ـ#P#	+&�0�E�G6ʠB�"O�Q&ğ9#�HȺըF���"O�Mjg����X� ��v���"Oz��da�H���cJ|�`��"ONs6������eb�G��MZe"O�U餠�2w�G�K�i�b�"O8��҄9Qؔ�T��$u:���"O��S�A�8�q�ٛz�RE3�"O,!�`L71gPP��	��B!��"O����8Ԑ��� Ykl�P�"O:(H���*��Ǡ�=aP1�G"Oذ���B�<��tω^���w"O���&D�I�Z�p��<�H��"O�X�fo:�"�Z��A�wZ��"OX��.�U(���9dir� "O�ș`C�5T����d�m	bՠ
�y��О<@,���	t��s�J��yR�0�4��堕5q��d@sf��y"��l݂D;`ɓn#�Y���ߢ�y�!Ҝp�Xz��?k�$P��� �y��)�<��� ?q����,���yb��|����d0�@6�-�y����(��� �+Nhnͫ2�	��y%B�$��k�kDzȍ�Aۣ�y��ϛ%�D �N�,��C!����y�$��ځ!�'_�|	�f���y��H1읹��,+�����	W��ybc�3(5�q�MX�N�Y #Q�y-Ͻ&�
�b@�e��PɂeW��y�/�� L����G��[���	�'&�y�(�?~z�����0� �H��y��	�1ѵ�E�ģ +>�y#�+(��)��1���U��yB�M�d�1A�ʕ2i�$�%�Z��y�ME�@,��B����t��yb)B�	Hx;�d�:e��B��ybO�hR�I�r��j�v��CL��y��w��Y��*k��Y�̯�yB�G�ad8��M��~X�B�V�yr�C g�	W���x�
9�yү�uN���X_2p�B/�y�'��P� 5��*7�,b�	��y�KވP�qУ�Y����`+�y
� h1�rf@����Q� >�yb�a�t�8ٴ��$�O�)@&aC����O���s��b��Q#9�� ��`:�#e A�΄�;S���{�'� L��+(<
��u���]�'��ɰ�B]�N�"�˰	 7w�
�a�+^
]��iܣ����t����Jq��$Q4z���'_d��(|>�ѓ+Ƨ*aP�q�ݢrF�D�	!�M��Q��#6���ā w �Г�у)M��� FB@���@�'������R�`%�F��>,��R�"��)�M��i��'{��O��&��1Ur��A��_М0!���0�G�+g&�y�-�O^���OP��ǺC���?)ݴ]��1UE�-,d�B���=n�nez'[�d�^�0�Z M},RU-�]l-H&�H���'-2��Wk	��>l�@�G�q��q��%rڐLB�.�>5�����u�O�6�N�?�g탵f�8��b�9X^�������m���O��CJ�Iҟh��y�ɑ#�t� �ʆ7nlhӁ ɿ�����>��D�S�$��m�R��)�&O�I&D6�3��צ��Sky�'���6�oӢH� f\7�"���DU�w~�`�+Jҟp��ݟ��Oϟ�Iϟ�����4��I�k@�;^z��� ��KVdS�7�����*��0��lyc�	��� ('ѓg��Yd.�x ����K�GP���	O�N��9�"U?Z�r�oQ�'�0Y�^��Fi%UQ�D���J�	���z��DTJ0$R��'W�(]P�?�����Ѽ<�,����s1�$,"Q��G��N��h��̛��\�M`� �0�Ql�M�)OjX
�-Ǧ}���h�Oa���B�'��T׮�38t��!�	O�w<B�'�R�S�t�.�2���rT��ra(�.��@=�n��JOl݈uӐ"�.�j���>qձO]��Q�iP�ᰅE�v&ʸ�S���~����'h� i;v!}���ϔt�.��I#�I?KD�����="�4�?qO|��+���� V?G�`{�`_8|��OJ���O��7��+1̝�����7�tL���OR�=�'ϛ6 iӠ�^�����Ӊg��P�ať-�4M땊W�Be,=x��'�����e�a�r�'��i����$�m ���g�R�Z����ʒ�g(�9��䄋C@�m�f�T5o�
=�w�|��'f�`�]�-4�P��X��Ωz@��$V��9۳�=E�J)�c�Q�0t��{VI4Z���}�:��I�!�X:D�Й�햱B�8�R(^ٟ�x�4`��v�'"�F��O�e��%�d���(�Man.D�Yɟ���N���O�ƕ��;w��-��:(��lRK�����MK��i��'���'�M{sl�'�l�v���p̐&�ͺ7���W�~t��'�r�'��n�A�	�o�wu�-����	�!x�@]<I�V��$Ey�#�O�W|�=0X�`��� ���?�O��1�fX�oD�h�ǂ�����1uD՛���]6��	���1��΂Q�t�Ɉ�U�l�Z�ʠ�ۆO��r ^��M�˟���4#�'4��'\�'��XQ�V�;n�x�R�3E8���'��{�Y�0i���)�� j�����GP���|,iӘ�))�d�O�o�L t  �a��p�N5�/͇B#�uHP˝���'v�Ȅ��@�[�muiP�&E~�')�����3��v�p�I7��-k���
$�ҫW�2��Ϊ6g��'|b��-���;�6Ÿ]<��Ps�
�]��<��D��V�o���O�֝6~��,�G��<�t�s�G vjth�����<A��   ��=*�aߕx}`� �'�'Oay�Ȭm $  �)Ԍ��\��������60I�MG�t��I䟂!��.8YT�I(�������s�X ����1s6![�n��(�2�J�jF
K���?�����J-O�i
�C�m&�����p�9D�����B�[R�y��O���O�7�QK2��R1�o̕�S��z�qO����ūhtnt8'	H�@�\�	� P�^���8�M��i��'5�D�O��'2��)G�n�n%�C���k.r��%#6$�8
a�   ���hO�� M�4�(��吳�;�/�:R�H2��%�'�R���Gc��	���OE�`��S�6��ZaKӉD�.	����8���'��n[]�zP�0��8����2���~��ƍ��.�y〜�f��_�:1[3�33�ORp
��H�@ �lջ7]~m��J �_���x�'[G0t�A)X�A��Ibrn�NI D�>����ϟ\��4���'�Ocj�h�XN��z�J)3��p{5&!�	ԟ�t�'����A�\�wY�A�\��	i�`Fc?	��4�^l��MC�O�RT*���hh��G_�;��9\�F��ŠL�d4����OP�4�.�1�C�Ox��On7퓃Uݮx��\�wkN�s)
O{������#[� Qyw����h}�uƟa�r|�O����[¼��E�S9��k$JO�Ub�Ǧ1=��A���!r�(��C��#8�È��Oh��O�����'��XP@N�a���9�Rt��M�<�]w�>���nV��R����S�9'�����'5�O�"?Y�MV+
-�=���>�f����R�D�O�nڴ�M�N>q�'���46��T�e��0s�,�O_���O���$��F� (  �QZ%-�'0�8� 6/�$�ey҄��\�Q��;6�� W NMw�F�VDAr��_���'1�8ʓ�&����N�G���)$���#Q5~����
s/��$�O����OV���Or���O$˧�yg넑!�>���&ҷ
� ��� ���?�f�i=f6����}��4�?!�i��(�� y�P�2�n�
�;'�Ƃ	Z6�C��%v|�  A{}BF�O��J��'�ڙ�FC��-e6X��O��6џ. i��ÝFL|x�
�Y��;��1 z<�D�.�����'�,6M�Ǧ��g
�'�u�%� V����iЬ]_ I��E�F]��`�XF8E�5�)h��e�T�K@t��e�ӭXۼ6-�����4
nJ8`��B��:�`L�+x�	n�� 4Z��b����7�Wަ1x�4n��ȫ"��>��0�� Ro� %)xG�L,oН��C[8Q����*#J&l��ݧ�MK0�i�$7����xIs%�r�B�ʤIZ�Q8���#.�GE�o�`�կWŦ�yd-�1}�HRe!?�գ���۟��?у$��S��(10�a�0���"A#�?9���'G�'٦7;Ra�XHL&U���̵3�DY�cD���0�'�r�'f��X
}��M��ƿc�>6��M�8�9!��dd!�Ɨw;z���'O��)�%�"ml��jӮ$XV'̵y�*X2t�T%1x��@�h��p��D�#���&��dˤx���wȻ,�+V�O�1��'Q��|b�'hRP�p�	�3{`J�<9�8�A�,�69[F�����h$f�80�t'��s��S�?	��344[�/QD�f��� �'�"uفNx���9�¼��ʙ?f;,�"C@�S��dk�'@՟|�	�[�H;�A>o	���ߴ{���I����6�MAсF7W��끯I�s:�	^�ڼ��&�Ǫ��!ө9@�TY�L�k�S-LT���K��l6�����H�3�8\����M���S�|�s:Z{���3cV`&���f�P���	ӟ��''1�����E2`���$���b�0�hO$��ͦu��4�?��i��S%b�ԙ02ʇH���ŏM�87�Ov���R���?����?9(O��;V�C(+�>Z7Ur��Da�V�Y��4o�r�.���hV�(cnQ�O��{̽�������G�н�f�	S#RLT�;��Q���lB�0���/P�[v�W������ Jn�8q��U�-�\Tl����dI�b�O��3� 5��t3D�kZ�<1G.�sY�=�ÓN�.���<@.p1�&K�&���ȟ0��46���|�OM�Z��!@��RD�m� 
��T�II�{׼��RP�T��՟��'l���|�4ЍwU P�pE����*!:Q�fGQ ��k�/d��:&�'ِ�&��
,q�eژKW��D #Ib�S
Ήe)�1�w�]�
,ܔ�rBA�'!�h��e����x��*
�������M����Qyb�����$ڵ;���Pf(KlH�H���O����-�I�-š�ʆ�8��P	��pT��ަ�̓�Mk�i6�S/Ev9�4�?���Nn�@�3/�?C����2� V4$����?Q���?	��?�*$l��!�^�PX�fm:v�5��뙧��� �DQ�[�e�w�'��C.����ڹty<E��ж+����'� HD����6� ����b��Gxrl��?q�KS��'����Bш`6Q*aU#M�J�P���ĩ�G�Ӻo�A̓hF�	Ё
~� ��Ѩ�<YH�'�̃ٴ�hO��������-2rx���Q�f�|����ؽ�M��[ ��K�O`n6-�v�˓��i����ص�Ԋ*<LmH��2{]�hrj�O�����`���˾Ÿ���P��q��DY��|����@�z��ό�\��	<+�zei�)�� �ص
��D�<2|\�j�t��)c-��?�r!NF�ZG��
�e��S�+?��ݟ`�ݴo�O�1���i1Ƒ�u�f��v�9 p&U
Q�|R�'B�'��'g��8Qo��0�̆61(�HC�B�b�hS���GƟ�o���4�޴�?Y NI�*&� ��'g
kq.ٸ�6�'�'  q0��1T'b�'��'2��7n� 	�K����;�'!'���%���d9Rxc>c����L
PB���A�i� K��$��r h�J�C�g�%����@ߛI|"�K���?�4%H�4,�剢U�j�$>��O2���O������is��Si��z& �V�=D�p�4��
9|%���ڏg A �UG}�.�������d�K�  Z�S�!�PJ�x.L �M@¦u������Dy��$ �(Vm�jwM�4�`M{W���d�� C�f���	�Z�M�D-���Q���4�U�U�V�!u)ל+	LiC������
��A��"��{j�mHǿ"<q�o 0�v5��Ė�Im�!��A�F�,�I�L�	Y�������䀶q���+ ,�T�R7�'�1O^�`##͢HQ�C�o�f��8�p�|r�{���ĵ<p��#�?Yϟ�-�B��Y�2�)�ɉ�O�,M�'e�I埘�I�|�S��L��C!Ě�y��%�$�J]�? ��q ��V��=�"H��>��x�@�'�V<���]�u�"uaT�ǜF"���@"9��H1m���:%`Geа^谓Cfc�D�*�O�o����&#�Аz�$��Gq��2E�ϲ��'h�yB�'�LUȃ�P�[�Z�[󄃶p��Д�'�X�G{�O�~7m��pi��{���0�wd֓#U�%n�򟼑ش��0�i��U� ��y�e�%m;4492 �+X���W�-���'�D�G�l"�呠�P>W2��82�i� �:�b�./��\2$��L���|,XUw��_��C���B|y���q� �O7�� #ؼa�d��Q��1��O��� �'�7m@�OM�I$y;��Q��K}�����I2U�}R��\`�I`�Ld�"&>JX�(ã*ړ�?4�i�`6m/�DQ�I�H#J�r����@����oZ���'�����O��'�X�$���G6��4����Tp�CG����Z�kA)9HEa��Ȟ; $ܖO���{��3v�\Z�R=l�*0o�2a�}Q0!�%a��c���9⬹@����9�Fqi�'�T�(��G�Cn�$bv�ص+D\W�iܐ�	Įm�	�?����2��E��-�j�0�X���)��(Z�n{��8*ۨIĖ@2��"�?��_���y�H�O�I�|˓X/��:����DJ�2�,C7!�"�rGMR08��������yBX>ͧJ�hq`0CU�\)��BN"L 0��R�4GTy�� G������'-j,�'W+z�.�R���]$f�ȧgaֱ�UK5c,��&���d�{V��7�O&t��B�A���`�*���HM�LϺT�Bdo��Ez�����ܑ�ň�]p- �IC�dŢ�c����o̓|ddc��<�����g̥�x$�Jߴ��X����� �M����yR�ΎX*��z�Z�DT�cP����?-O���O��V� ���e��9�Ҁѡ�ѐ�M{Smʍ�`��f�OIV�%8�k�t�X%ĉ,5\Dг����h�v%`ݴ���� �
r��@g�J��m��	A���O��}s�\���3d�'�S?L���%�@�	~����4�� �,�Ȇ<�D)$�&�O����#��Bwnt`�a���A���ġ<�6��?����?�)�6L`��O���N�i�����Dу�	�O4��Mm���CB�$x��$ش��O��8Z�\p� �ɰMR�O=��c$�Qqg_���t��ip\�aP�Ϡ1ؤ�ϟA���_2xe0K��i+���p��|8��O+�i5�>̓�&mjCF�#����㩗�N���ȓF�P��B K)u��Z�Y �G{��'�N#=a3�+T�5��*R�Aꩬ���n�͟��	ϟ���k�c?F�������ޟ0ϻ+ÌEv�e-
h�GI�8]b�(��`���0�"�\���� �m�g̓y �ū�^"m���J6@5�Y "�)
r�]X����?��=�GZG�'�T�V�<�q�H(N6��Y��Imx@)pe����JixX�	^�g�P̲��V�i��86�nX�l��z_>a.J�b��Fb�goFq���O<��YA�����|"�D�!i�)�b`�;hFN���;gL�=@�>(r�'���'d�������4yd�ŀN��l���8�H%pD/��,PJ����W]vu��40�0���6KC�����}��膙p�b����`)�p��՟��(h�0tQ�����p��+��ˤ�$���������C���ێ��<�O��ж`��$��֥-0b�"E�'�y��D�����0R�(X&SP�i��lӂ�ᦱ��4��I�s$�nZȟp�	�52�|�B�� f��Q)AJGv� ��ӟ�Q��֟��I��x� u�<����W�D�+P���<ǡE� 7E���7ur��"�'a���/N Qv�{�
i5����W��TSu���O��1'�X�h&Dv�(/�L���Y*,O�y�D�$.�Y#	�sԀ�h��|��'}�Ղ��^�HxX��ь6�������>Q!�i+<q[G�G<4��&��&P�����S�0s�B�֟��	����O������'� z�C3{K�هB G��X��'^�eڃGA�sU�sz̤oZ=f���'��)��^lޠccb��/��"���D��ɜB+��1F��&�$}Y�4�H��IǪ;ݬ��OW�-��#
7w�,#�g_,H���O�Y6�',�S�<�qME8D^d�:�~wN�P�nl�<�ŁZT���1(�t��b�,�P�'E��*ғ B�U�S� �µx��)t��6�is��'�ba`Ũ1���'T��'�8�aQ���1��	2�ǖ?O��a��F��-�sz�1��J�Fu1�1O��B7�ֲy��hHB�rUp�c5)�%W氝�F�D�A�C�&�1��(�Ú;F���)6"�1S�9<@f5	SC+-�1Oh!	��'����� ~-�mkɗ=|J9�	�'FD󤂃<!V=�������%8��?9��i>e�IKy2c��*
���2��,fYb�"��e��b��4-���'Y��'�֝��I�|1�˘\�p�1 ��%bA�`PD��-�x}�
0rb���"U�17-�����05g� B�s�Z0� ����U�%A���#gof��q�ܵ*OR���(<�e����%��i�p� vBяin��l����������?я��C%]�}��hG+���CU�8~f!�d#_�Tq;`����0�95��Bd�'�6M�Orʓs��H`V?1�ɲhƈ+B�PĹ���_ �|�����a�����p���|�d�R�E���
fe`*�f� S�&8��IN�j\޹�$���@ ��SfH�.�8�<��N^.��'썎yEp\��Nζ"�!H�@C;G��ȢJ��<�X#}�<I�G���Rڴe�I- ��a�G@f B`g92�Or��$M�;�-k�c��A�����D�O0�=�'s�".�)(����Q��|��-���Ԋ�?(O��cV��ۦ���ޟ\�O�6$3��'ZJ	�W��:-@��oܖ#�:�I4�'�e�O�����l��`v����JߺP��r���:) g/		:�����5��$�	$qJP�+O9�ȲC��(�R���Jؑ!/6d����]Փ�p�	�O�Q&�"|ʇh�7"�x�B��7Ӣe�W��V�<���4��`s����͢��P�'-��}�Ġ��n�`���;vz&����͟L�I����! ��X�6���	�\��μ�g�4"">�A����Ĩ�yV)ZN�*�R1�i�r��6f���œ���y�Ffg�0�7�ގf��鶠5%�ei��`ӈ�Ò��?� x3�i��Ȭ�W2O������"B����W��C��iz�'��	��X�d�O~�=�eˇ#����ԉ]�P�l2�EȬ�y�h�L�Bt��J9Bh�0�$^��?��G���S�l�'���	�ǜ/�|�B��P�`:���'��*��p�r�'sB�'n�"gݭ��ߟ��=�tlq�l8�Mt�RL舑 ��+��ei�D��PU�)�'�"O( ����(Gڢe��o�rm�&��?Z�s�
��7�NЉ5*ZRB��PC5�T�\-�S�G�5AV��&��l��PCC�Hş�K�4p��V�'�����4�?�G' ���U(�{%���`i�����0>�&��e�� 3n�a��2�I�h�ɫm��%��4��T�Txm�;�?1�<ِv�.Y4�b� ܬbBj�A��?�e�ޭ�?����t`�ly6]��&�?Z,�6m#)�&i����rN�H�Փf�+�'�fE:�&J����9��t��i���[0��[W V}�@ᖄ�Y�P��3�ԡL`��"���On�d/?eM�,�p�q���d0����Jo�^�,*6���);��F��@N`��� �IH������OT��UO�@R޽�D7B/�����'��	�TQ��hڴ�?!���iQ�"_���7Y���c�-6�dH��'XX�d�O�����t��s�aX�	��u��X>	j	��)N�TذKFT~"�iKd~�%ؑͼLP	qʵr!DI�O��t0f�ȧH�"�+��H	0��x�O�Ab�'8�7����e�O8^	�p���Zq��ȋ<�t�N>q���'P1O���`[�3�D1���3�x3�C}B�dӦ�nZK�	�X�1x��K�IV=�v��D$�4�U�[ß���П��Ì:Z�u�	�٦����?1��˒sp�{&Aلi��`թ'I�*���!Z&�?ϑa����|�<����e�LE���b�`�2�#|?�R��/�?�ԍ�T�܍�|�<Y�A�=$����J;]y�]�t�Y����'��X����?1���:5�9r��W��<�GJ'#�B�ɟe��D
��ܨ��u!��߫E�ʓ\�������'E����s��id��+VY�ʙ>(P8Y�'���'���a������<�	8

���d�S:tr��$_]��0U�������ɜ-��xlۍ[H��㣃��(O*UqPa�6n�h��@ʘ<�$��M�!2D� �tM
lcbXXp*�� �.�+ ��+�(OP��/�5d�,� ���9�l H�nێ'Bmh�`IDz��I.R9��{a�
�f�@=��H�>���OLc��ه�%[CP����'[��d��5�M�E�ܴ��]�E�� n�����	�>*��(��D.��L!��A,s����Iȟ��O֟��I�|eFI=�H��7c�d���"Fzm��Ct.V��s 
����3\L���1�4ZBh���6(��,_����Z7�����H��%3��-�gb��I-��e�0m#4�(�ԸRcZ�L�H��ȓ8F&��N�B|tĎY�2��?Y��4��9��-��	` M�0�;�,H%O��OՉ
�)�IܟܗO��EB�'[���LY�����/
��x�y��'�bAC#�J��I�qȲ��M�-�f��T	��urB"�f>���ω���Č>좜p� S�P�"�S�D��}n��`3�)�	
���`Z(�#�P,3����, ��9F����ݦ)�۴�?9��i��W�2Q�«״d���1sb�^��'��P��F{��&rp4��pCX�M���c�N@#i�џ<ش_ћ��|�
X	�"��4����t��/5ݪ��5�'��'�f=��.Ǉ^��'�b�'Ϩ֝j���c�[�$�����/H㮅�uh�^�fN��Mv(̂�/�ş{v��龟`З*����S�<mf��0�͎m��I"RL�-E�d��&X0�2b>ղ���
��� \Q�&��FV�0�瓾u����w��ї'��{���˟�'r�4r �R:J8l�dF�sj(��"OB�zD"�	Q-h@����cn��' "m9��|���������i�������	�xv���
?~�`��O`�d�O0����?����4LH�8{.�1��1j���h
���HaQႩ(����`�Չk�zԄ�ɕ2�p��J^���H�Q�1�R<qQ&Ś$��-�ୂ?.���`0)�. R|���3�9���6�6p�p��T�Z��D�<�p��	�Us��^A���t$���{r�$��Y�ԥ��.��o� ��Z��'�>7-�O�˓k
�� �iKr�'����V%%���I��ۭ&Br��u�'E�����'����>{.̱S�^
���,Z&�~Uy���yݎѨ�+O�6��0Xe#�z�В�
Jmb,8t �2-�!R��7^��R%�-�tA��^�[I���D�+9��D"�d��Hc��@b��'��] �H�!��C�Z<��7�ΡE����N�>�,�O>=���N���s�.ڤ 0 �u�|RbE�8b�'��Y>�Ї�ʟ��lZ%7�(Mk`�����N�MB�'ú�c�jV,�"���A�i�<o�|�-���g+C�Y!�H�S�A�)�L9���%?�!Ro=�%C'�ޓ�l��3K
�y,1�V��!}:�90�H��
�4��%�x�%�#LV��'L�� ���?1��Iv���Ѐ�40�%�č�,Cj� wb3D��r�/�6�C��۳T���(T�;���>�!�&�
 ����X#F��@�O���O����x1��Q���O����O��D{�!86��.U�0�@G�ք+T�D��A��s�XU[�/���M��	?[x��O���	-�Php )�S��4���$IV\P
����4���N
X�a����4ܾ�c?�f�fa�?Y9���*m$t6�,�R��#�򕟸���O^�d-ړ6�L�����V��#�V�n���s	�'���ubZ3p�:\���K=`��+O>�Dz�Or�]��CM���蹙�lG]��U
��#�vxj� �؟T�I������?��	֟��'��칅A��!�c�W��l���lv�D(`�כfD;,Oep�GӁ5���['ύC��5z�/ȷp,2=XR��1��XwiV#.�@��Ģ^�%�"A3႕C���<5K����C��Q)n��'��FD\�&�O��d0ړ�O�@ᑣ
,�vh��	�|�%"O.Q��%V�B������!��څ�|BK|���$�<��_\��Ou4�F��0�i�Xt�������O����O�Q!c;]�]*�<�|@��IX	<Ƞ9BJ�-������X�|��
h˰���H�)�&�v3d�T�0,��AOF@J���8��$��'VZB��?)�O��v"F3Shu�e�&�D�#�|�'OtB7-�Zq�銥�M<B���?��')��	-kS���T��"<�,b����$ؔ/��S�DY>q�ɏc���%��|�ٶ�y��I֟,A%g�Z%�p�d�H�T����
�R�',Q��c�5p�<�u`	=Ktz�O����M	juZh@��6��<���iCZ��c�Ja�V<'&��/�I?�@��OD�}��'��a�r�T�M��L�s�%J�M8�'�ݺ���n]��3S��9s��ˎ�Ax�O���[���-T��![�[o��(Ob�3������?����?�+O�hp�/�-h�@���1�"�Yt�'�PA�a��R�.�c�_�rgf˧���yB�i ���f��|�pq� d�s0T�处 J	N����*>/
}H���y"���-��7b���� ���?��O>���'k��I� �D��!�ة�0����\U�����'Z���N=aP�����F*�Ԗ'z"=�OF�ɀXѾ$����(t��l[�tV�-xe/A����	ǟ4��FyʟX�D��L}؄���Y�zI�I���.9IrE늳�BݪF�x�d���'���CO̡Cb�A������M���S"�t�B�p�-x8�`zp��s3����#_?P�f$�T�MZ�:�$�O��=Y��D�u�hI�+��e5� �S��m�!�=�lع�Ȑ�RћEN��'!�����S�@ ZX%?��en��Y\ !G���3׭�O���?���?ѣ��<,�Hi�D��u�r� =��<
�#	� $�ف �8��eZ	Ó7&�X���;Dp�*�Jօ�/\�*������+]����I��Ha��O:��>?�g�W�ݚĉ���.���E�	p�HQ��*W��҆ WkCx=Z"�"�Oֵ����VU�� �:q2�'C9��D�<����?q�OM��F	F���1I��$UI��ث\��'��T���ߎt�@=��cF��0�2�ə! h��;��H� �S�K ���D.҉cE�S=s��@��F+��|�ƊӋG��s��EL��c�S~��!�?	���h���)� |��7f�=V4<����Y�!��"O�	����o�ިځ��4� D;a�	�h�>%�١$b8��	S�B�i$�{����cK�<��������ɣ4�y@Ԯ� 6�	�� J�|�� G�~���qfC�v��$1�,*�3�ɻfJ mQ�[�!�y��i[J�%j�ܘ*`\�����&��T!�&6�3�I�i��M�VM@}$�b�\��lXnZ��D�]���O��3����B��FĀ�*������JC��T�YY<�]��V�DL���-O�Gzʟ��"�%��j�`g^A�F�#?��"�e�8H����p=�pG�m���UL!fLu�bFr ��)m圄�#a�+t_����<2�CT�֛d��8`��!tG�i��
N!T��=iT��1��ȋǓ;�P��c�L���<k�@Қ;��������ش%���Ex���O:R�P�(L&=m��@�͍�yB���}ɚ�Ȳa�Mi�������2���Ay2�Ӕk(7��9���,S���6�Y;M8m��n��#^ў|͓OjE��I"C)�pS b��`۾D��D��0<qC�[�'T�g�ʤ'9:�s6�Y(5���Ó(R&%��9���������g�~���+��k:��ȓK>m�� P3�|�!����wzh��I)�?!'Ŋ�  �$-Ӗ7H<�ХSi�i����MӲ�Uj�Oj��iW�;ڮܹb�Y�T��O>�����I�h��OB� ��=�����;�t�c螮lٔ���K�I~��,k�B�X�+�7�68ٔ��Q>1�Uĕ�d�`y���W.X�hu�m(?ɂ����p޴eߑ>=ͧ&��e��)�#�JUJWF«u�Z��3S`"�)N=�ҭ˴פ �n�Frf;�'E���;�J2\�P]S&��-ULZ�Z�4 �l��,O-�&b�|Fy��!?��)@���\�n�����ؘ'���
ӓO�U��i��x:��7JHE��!�<���EM��P*�!��rC�Xr�B�P�O�a�I@�\�D3�3�I�|���5�#Z�j�Ӡ��^\$C�I��LhK��]�I�R�������`�j��"|���׼������Y�H����R�z��g��]���U
_�]�����<p�����O����T��b�N�s��2K�?���5H�1���:�f���OT�$'Dp�⩋�/�P)x��X(�2�Ӕd�\U�A��B�-�Wj]=LQ�0E옞'<�$)����J�
Iן�Ɉ�N=>��4C�d��I��>�d�O$c>YS�@�w��ԋ�l-PW`,�'N�<!�*^��PE�ϐO?�3�OT���5���7��D�As@ճ�+��%�c�4i7�	�(��L�	�l/Z�˦��O2n��s�O?2�Ҹ8r��cʥr��pk��-r!M�Yx�+6� ?@@�lڼq.�'�O(�z�.�:���A\�u����'q�jN5jz���uӞ�!����&]v�9��)��-@��r��71���g⇑B��D�)�R�'�)�	$?yd�n^���4n� ��A�}�<�����,6��'��9md�(+Q�Z@��?��i>�y�d˗r�q�WCŁ��-�<h�H��	��qPH��Hq��՟���ٟ��Sß��U�� �xr�G�
��p[��H���$p,A�'X�YM(@ȟ��
�L9a�p��ゕ���P���0�M$C��<�P�iB[�/�&9�O25�
*����Kଁ�	�QC�4
����>&��?2���d�O$�=��'_�y[�b6'"�����H��'�jP;#S l��z�9 uF�h��'��"=�'�?�*O̘��o� 2�����%��4��k��t��5Y ȍ��4��O�����D�O@�C���Q�*B/V���$�J{,��`��+XNlc��E��M�W�#Oh�`ᄖ�DC��	�ᙇU��2`�N��y�w�xB�m��@e$���oS�U��#<Q�JQ��()�!U�QO�H���A="A�(J6h���E{���lu!�#�Va��Vė V2���<{��!�̟o�Txc`��)��)�'�@6��OʓC�4i�}��1�����E�kA��C�,#(blشJ��?�����?����?�-H)a�A��*P�F�6���|�N�0hB��@o��%�P��{h��з��z�L��3I#�M�C�� ����H�4#�u�a���w�ؐ`!��;��A�����|��L��)0R�!g�S&;���C$�ky��'bYX��G�AC1AO��*�L>q��4����'�>�P��Z<0 9E�"S�`,O�I�C�O��3uN�O�˧5
��'�?Q�HN���X��LE�6#l�X�e��?��*��DP�e5$6���*�[̧]�Y�Oώ�2ь©Rb��i���\4 �[f�iL�Xw�C�Dt�ڎ�i״/�zܹ�]9 �ܕ�4(޽�yb���?��������� �1�U�Q89�c�%H�&v(�jA"O&Ё��եA&x3⅖�Ҙm:����O�Gz�O|8�a��Ԇz8	�!X-�Pʤ�'�B�'��hH���>J�b�'t��' ���'�ڤ� ��	�`���J�AO��dk �BtG8WoH�0
KҮ�g�''P�(bĐ'c�>�*��A���9�$y�B�'� S�D]X� 6f�S?x��Y�'-?�v-��A� `ʥ�$a��0�[~�+��?1��hO�扟`����jD�^����C�bdC�	"6�I���0,�B�j	�l��I+�HO�)�Ot˓OP�ԓ��M��
���2F��ٰΙ��0?�J�wX ���B
!,V����L��^ʶ-Pe*�5o ��1"��/��F���d�~��l��9d`C�>xS�,�<�Iᣖyp�����N,��O.��A�'���7��;Z��& �`ID` �'�ў�F|���jU x��c�t����@cԆ�y�m��&��!���I�j���𧈬����Q�	Ry҆��j7��O@�$w>%2&���U�@� ʨ��6+�Oh��cK�OZ���O�9K����FM�c��8��=�v-{>��daZ7��H���Ͳ�6�Q�m;�~�����f�*�(Xg�޽�X����D(&P�ˋ W��])���;Ѣ����\�'��ء������Rbm�4�AVE�M���p"O|b�dRQ+Va9�c�	n��ǜ|��i>U�+O <�G�G��Bu�,��P�Z����ğ$�'��Z>��O�`C��9q���a@:z��A��'�Q�,�ٴ��}A#��'G&��c�L�@3���|�rO,�I|�!l�;,�ԫҏ�/u#f,�.�$H���'S�U��>O�a���'$���y��Oeb�H  ۨ�#P�=��}ɒ/�Ǩ6��O؀���O���	��H�s��K��yR5����ѿ8���1�ωY�$@*A�?�� ��,��'��.�O�$�l�Di� a N]�$�Ω�"�V9\��[5���*�D�O:�땀�O��Ɉ'�0�s����y0	y� ��h���~��6.+wU����?Q�h�\�jWU?	��ן�����@����c���rE�`�L$��*Z��?	���,�	�_�@����?��%Khn�FN�ȕ3%vaP��?Y&���Կ�Mc��'	�����?�c�=gK�����	�?![2�@�:Y:"œ�\10P�������$�%Y<U�I�|XYwOB9Ot��Pٟ��$����0�a�#~!F�
�G�3$nA�`�k�:�I�_�V�mZ��M��eE �y"��P�	�ru�`�%V�T�v�
m`�sm��u�$��<a�� �M�i����'�Z�dk����gL�)h6�H�5��O��7�(�nZ�d�U�I~y��7mJ�?9��b��-3��hHP��*sh^��0���m�!�d�/Z=�QCD-��� u�ؠDx���'��'���'���'n�'�B�ǌ��1�b�CZ>r�B����n{�6-�O���O����O�D�O��D�Oz�$�>b�~��T�����iǒt:�m������꟰��֟�����I����I�2��sF�<,Xn9�,�V(�4�?����?���?(O�˧�~��_Ť!(F
08�h,XB
�9�M���?��?�����O��Z��VP<���ؿ2?.���.FܦWb���?���?�N>���@@H˥H��a�����	A#�i��'"S��S\�ԕ>�7��?D��V{JL���L�<)�W�̚X�ы	�4�$0����B�<	0e	?�����C�p�
D�y�<i��Z�?1<A:Ҏȍ"k@�u&^w�<�F<t��h�n�1F����t�<��ÐT����e� �09n�*�k�m�'�"�'��'�rJ�Q�ڱBBb�
`�45 �%Vr*v7-�O��d�O����O2���O��D�O��dS;z6 �6C�!b��ܒ%��	%�]m�ݟ���ş��	����I���	�p�� ��d��ҏ<ĸ�a��v����4�?��?a��?���?A���?���L� t�%�ۦ85�l7�M�`�T�t�i�"�'���'�b�'A�'���'�$�:un�A�MjƪM#}�}ʧ�yӼ�$�O$��O �D�O@���O����Ov��%k��4�� 	�l����CƦ��	ߟ��ܟ��I��Iޟ$�	ȟ(s�E�5��� �$%~(��"H9�M����?����?����?���?����?1fb\-Qnbu�"յ+>(uAP1$����'_�'M2�'T�'�b�'�2��LŖ���U�j�Z�!+
X6��O���O4��O��D�O��$�O*���2>-����'D�8��GN�'mH�oߟ�������ǟ��Ɵ��	ӟh���>90l�t�P�3��v�ڍz`�ě�4�?���?���?i���?����?y���m;�"�$'�\L�B�_�T��e�i��'_��'Z�'4"�'���'v\�x%��z"���Y�HH�4Cw�*��?))O�#~�R�'L+�{Q
�Jؼ�p�M���Mc�iUa̓��L~��iP�NP��9g��tƮxڤ�L�x)�Dp�f�IUyJ~zh�4XerM��DM� ),t^���%R;`r�(�ɖbLeq��Ưc"�G{�O�䎣��Q
�&Թ(�l�Q ��
R��\��&�Lc�4-��L�<A� �YԋҽF�fH�P B<Ҽq�e�'��'"�˓�?��4�y"^�|*���!�HU�S"��x�d���<�U�]善8�e�w~�O��5�3b�o��D����h�^1zߴl�dNH4���vyr�'��>��99��z��~�c�&
W˰�DXᦕ��"?A��i�B�|�O��9 �(HV��\�1j��7Dp�j5O���n�l�d�Du8�s ����M^��PA׳��$�Ѯۭ~�:�JH�&�p��	Ο��'�1��]H��ۊF�%�TG�)5x1��R�D�ߴ"RA�<Q�'��'�ArD�ׅb���G':%!�S��Iݦ�̓�H�pu�6lX�4r�2����G��C�j�pz�����Ћ�ϕ"����V�޼m��-�rN�O����I�di�n�0�qy@fX"�LY��@0$7!�+`
��:r��0w�x�ѭ�z�1O|��-�y��R`��$X>��C�Ϣʊq	�,o��
g>0*qI癊�R2�ݬ
en@�"�^eF�ө�<Y�$=K�a	
Xڑ�����0���s��ж>l�	�@;+�l��G��z�7Ô�e(�+Aɾ�H�#�ȠNW���r)��o���&!��M�����sS�;\�Ԭ��B�cAp�1�BC�3�.�U�5r4���?q���?�'���.��N"{��;a�jS���?�	%�Ms���<mr�x��'H���i��e`��C
x��F&�(f��X׈ԛlt�e���'���6�I�{�`�ifX�mV0A�3̖"r?�\�Toz��S�f��n�9��(j�lx �D1D�Ċ&(�|�M25�]�@x�w�O.l��]�Gߠ[����f�lӊ';��vkP5e:�@`��+*�����G۶`�Bđ���l愙��J"GL����Jc&`a���L�#��T�$A֬T��P'��@5�$�#�O(S><}*DK'#�~�+5���Kp��iLXPZ��q̈!o�b��$l�r��'1��'��� �<!�*��O��T�Ɨ1-C�u����,�	ş���DGy�OB�O�7�
�����M�@D�T �}��R��'���QDfd�>���O������$��S=P�BG�L�2$�u��Q�,��	� �^�'S�'���O��D�O8��FL4k�����Bđ<��`��"��5�������uxrDO<ͧ�?��F��T�8]�Dn��r���,O��$�O��D������4�	�`B ��r�&	ے�M�S$��1��ޟ����t��d�H<�'�?�L>I��G%i��cB�Z�P��{!>���+`F��ٟ`���p��K�dɉ3���١��K��8�p_�!����B,���O���%��<�T�]�*����V%@z2�,��Y!���<a���?Q���DĞXn���������oK^�*���D.8�D��?���?-O����O(�Eܟ��cP�Z�̩��3<M9wX�d�I��x��ayb��0!(Z��t�D���$�͒�g�DX$r���O���O�˓�?)�%���}r�Ý{ ���ͅ7ft@WHQ�p�Iݟ|�'�x r�I$�i�O�睲�)*f��bc��j�T5�D�$�<i���?��C^�O���<Vj�p�E p���C̓�Q������M�,���D�0y�'�=�����j1`�JSl)��?��J�4٩,O�	�O��>ae��l�r�,<P 42RgF՟���ć�M��?�����x�O��(�'�ͩ#溈� 
ڟ{�0��'�q^������ �3�I��Y��vg�l�C�G'fZ��k�N��Ms��?�����i[��x�O���'o�\�@�X ��0�C<3�z��Q������Z�b3�	�D�	џ���=g4���tBS�߲��s�ğ��ɿ��H<�'�?Y�����^G�4��*e�4p&��6_��D�O�0�D�O��D�O���ON�*�Ӿ�,�b�K�(�D�OLQp��o�ş���֟�����<����Y���d��+���*C�<!��?y���?A���?	�Y��U�պi�t5r`�A7��i�6D����'��'1B�'@�^����27��S�2�4D�"Z&�Fu�tɊ�y��'D2�'��'��)��Y�(7m�Ob���"��m�S�
�tIV���H'8�d�O����O���?�Fխ��'!���p囄5���Y���\����?q��?���t܎��G�ij"�'��OVx�&�J3p�P��kˑ8n�����'sU���I�r?���d�<�'9qn�1N��H�����p%�x1��?A��"��!Ja�i���' �O��T�'�H����t��t��cF �$_�|�I�X���}�i>�O��I#���N�
m�pHU�vK�(i�Z&�y�i!R�'��O���'��'Q�ɳƋ�\f�I�3��*��|�V�'�&@�w�'pɧ�t����'���s�@�yl�B�f9Q=��������O��$W�/"���O����O��$�O���B�N��h��n�^�h�w��O*���<Q6̋3�䧀?���?���U7���p'��Tጔ�u�N�?)�1��"�i�2�'o2�'A��'�yRC�q!�,�A�w�؄�7��D�3LY�D�O��$�O��D�|Z���H�"��u�>qPC��A6u�Q�*K���'���'_�b�~"(O���"N�~l2Gm˃%#���m�+
C�19O����O����O��|�D��H�惘dltB R�`m�E]�DZ��'-��'A��'����x��i>A��[�������W�z�(ETy��')��'P��'鞍�A�u�n�d�OΔ���N�ȴ� ���Tfj@+���O.���O��D�<��j�8yΧ��D�#kZ&�{m�n��!#Te���y��'�b�'T��^*c� 7�O����O��IɁL@�� Q�^3#�D����O��$�<�]=���'�?1�n�^�ͧ� p-v�T?l^��3k�uPl���'��'n�p��Haӆ���O �D����I�O��	`��/�v�b	CY��:���<��iVZd����?�.O�+�K �:c�T���	�Th�d���ş8s�D�2�MK��?�����'�?9��?Q�w~��k�U�o����g���?	���?�?�N>�'���?ɖC�"�8-�6�	Ѿ�g(
�8:�&�'�R�'oz����OSB�'?��'�"���݀"N�1O�t]��d��"���'�剁L��'?���ɟ��I/iT���ǀQ�#����n��1��͟�°�^��M����?���?IY?͓����"��\I�IY��N��i�'����'���ӟ���Ɵ��'�z�k�̃�A\��y��o^�L�5ض3:6��Op���O$�dDG�tT�L��� 9~<�ڐ�`�P�	�;	D0R#�c��	ϟ�����Iџ��ɬE.d�I�4�P�ã^� �=i�OA;��-��?A��?1��?�+OZ�$26�	�5�V��)G�C9"�EoG�rm��$�Ox�$�O$���<ifT�|�O/*́��7wSL5*��u���3�'�2�|"�'�b�}R���9%̍Nn>��煀�?_���OB���O
�d� ID����'\�'q�4!���@�C�2��rM�'�'�b�'� y��'��)�텺Jv,��`K�7^�,r�T��?�,O>5��)����O��Oqb˓4��9�hPJ��jvA�q�^�����ɼ[8 ���n�)�S0�"�0M�xg*�˷j4(�\�ò`l�ϟd��ş��S��ē�?��,S*]��*��T?R�pr'��?y���$�?�I>E���'+� �í�[��S�BK�@¦�R��l�����OR��
�N%����͟�ϓ ���U��0zk�p@1(��6�t��	�ɓ{~~�&?e�I՟��'d`T���l~�1OR)����՟�������?	����*�0����5<������ "�<�,O��A�>O���?����?1*O@���g��,`aA�XxzB�� �>`$�����<$����ៈ*R�K6/�����،h#Y�D;P��zyR�'H��'��ɩ�R�''aXd(�((tUpBR������'���'�'���'r����'����2K!��`�ٯ�lu��'�r�'"�'*�S�>c�r�4�?Y��v�\)�D�44Զ��d�on�`��?�K>i���?a�l��?��Oh��U���bFǴ��'7R�',�2U}� [M|
�� _�<�*� �i��[��0�Eo�����?���>�d0�Ov���:kLZ��t���F�M����z��oF�T�'��˿<�UkQ�BgD������f%�a$�ğ��	���1���T$��>�X��M� �a�ğLi�=�.�O�E1��������I�?1#N<�4�y ��.\0�B-��n�y�!��IΓ��S�O��b�% �:A�"mC�`b�}3���?.р6�O����OxE��$�P��؟t�I�<y$JSh����l DU�e�䟨%��k3A��d�I����	��<�	�4�إ�l��f� �c��Omv���˟�B`А���?�����B��C���q�2-ken�X�*��*O� 
�;Ob˓�?�����'&o�=�$"�=�<� �JܑJI��[�
�6!�'���'|�'���'��X
3,N�T `�R�~鬼sס�w�Ҕx򮃖�@�0�Dɗ�I�F��q� I�oW�^���h� x���۴�q��9en��>v���O��$�O֒O��'rc�)�ǝ�x��+�-]�� Ծib���O��D�OʓO���, �giW|X�F���f�����<�� aN	�W�:��Ŋ2�O$�`�Ԋ$�Nd�ЅD���9��'B��+2ĕ'Q�U��)yi9K�+ 8�%�@�0Pyr(���.Z��L���^X$�cԦ�'eAF�B�I�!`2E��&|�*s�G�,(���FA�"����إ8�&��áރSl���Ɩd ����@�7�y�qDD�1�݁OS2��(&RL������EBZ�9Vl��?A���?1�@��?����mĘbX�5j��C��Bt�L�0ź�[� �y�\�B�L^4s��t��	#'6Qr��+i�S C"A�H	{򌙿[lL�@�q[H��ڭ��)�a8F�<��	��Xn��)� p#�'W�0@x��g�'C9��<)�	�Yh�C�%N���,BcJ�F}��8<�nq��IE7*>�jf◍M���;D�i��T�d�Ǆ#��	�O�˧5����|Đ��GD�*8�1��H�?I���?!���7T����F�H=�7��i~�pի��\���C�&7*��y4(���]	�qqq"ض^������m�<�� �%���׉� M�O(lK�E� ��:A���>?)2��ɟ��	q�O��|���G�B��d馮��GY��0
($��)�f�)h���a5t��`2l-\Oҁ�=aP��$7dR�c��i|�5�F�
jTs2bf�f���O��4�Iw@�O����O�6�D�z1{�)]"
U�аS�b:�tj�����v��BF�Th��D#2h�5�|T5�,{a��}�F]�3��Iy쌢�ī���)��	&-�A�2n!��2�J!�Ӭ�y�ċ<�Z�%M�P���Y�!?���`򉛣H��ɤ:a^ R�%E�Z�������@?�B䉥b��G�Z}.qS��Ȳ]���'4R	8��|ҭOx�ԫ�)`utaxEI׽k(^4#`/ ܟ4pA"���n��	����Iǟ8qYw������ ��n	�7$�H�,��f ��C�N�`������d�H��" ���Mcժ�
K	��?)Ҡ\+�&��_�2x��$˯8��H�rk	&\�q���>Xx�;3b�q�:��]��RS�P�"K��A�.{͵�&��g���OѦm�4�?I��?����?���M��.�*�8t�e�ь����͞.*�r�'$ɧ��R�W=��uz�ŏ���+��"Zu�Po�}��$��ɬ<mY�.t���i��t�NH��\��F̷tؤ���O��O�m ��O��$�O�@Ó���Ydʆ.C� ����(�/DJ�a�G^-/f�������-��x҃L�K�t��-V�#On��5���N��G�,F ��[��P�n���a%M�FYGy�(�5�?�7�iuZ-��"OW&�!t��!E�-)�Z���O���#�i>��'��!���U&o*�:���2)ۏ�=�'P�@aFӷxx��y�$J&U����fӰEnLy���%Ch6-�O��d�|:W��7x�D F�J L��E��,��M����?��PG��!/�'O� 5X�ʧ�u�O��H���daؚi�:�����'��8���߬w�u���ܜq)x�&?� �CG�;nX`(T��%��d	�E6�I�?Y&��_̦-2K|ү���0ä^7]��H'�Ή h���to�C���?E�,O$1Z�)�=tP�H[��T�`��'-�➠��8eu&��6e�~[�����;x���G�i��'z�O��#�'�2�'q�V� F?�  �e	-G/"�q�	X�6$�aԤ�r\Tg��'��}�OM1���q�>1��&�-HS<��É�A#W(X��Qa�_=�d��Ή�2�>�&�r�+� ��0l���T1ހ�`��'�06-����� 0�>�6H�i&�Ӝ"�.�q?'��h#�'Fa2嘺(���:��U(~Q2p�f(��'�F"=9�'�?yڴqO���E�@k��X�d�Q�n�2���'D�Y8�N.O�"�'/��'����矴���j(8��^d�mj��-N��-���i�h��#� }��8�6o���xnO$(}>�QU��,�x!�&��_��R��^vX��m�m���]w�pp�A:ڔКv�� ��$�5n��E��-F,<���B0u���F���?�"�i�,O ��O�O+�W���P%�]yz��Vq�<�gjE�d�$ �W�U�X-Qb�r�'' 7��O��<:�4x�i��&%؃>G�$
�n�Q���ڣF��cR��D�O��ď�g��d�O�� k�*�rS��s~��@���!�V1أJ�O�H�P4Y �P�	�-����Uh��[�Ҡ�G�BL���R��7�^p�-H/U����'o�x���?�4 k����M��f�1V��-vn9�O�d�O⟒����\]r�ը��B��n�c"Ox��aM�7���j�c�	��}ʇ���M������3�
1�O��Q>1�e��>`c ������>�8�ȲHF��@���ʟ,�I�8�B@&SC�)A��&	��p�����]�FMx4+t��Y��	�����b�� ����	mĭ��I<G�Mr�E������C,y�"aj�A��OTp�q�'8���AK��pÖ�4�#�B�Et:�����?���ĖWS���-��ޤ��#A���0�{'STl���46V���̤qք*��Ʀy����i>YzM��������$n��b�L��ćSu������'U�m���C����*��h)U*��3�>	g�R�!gb��S|Y�)�Ţ��F.--0ݸ��Z9k��3��<����yw
[�'`@��t`�>1��Y"�U#�����j�"�H��ɡ
E,�Ì�]��QkZ�RB�I�w#��ؒ�H-e:r(���p(➼���4���(�hx0 ��H��``k�$E$�d���'=�=ȣ'�� ���'���'^�֝����)(vK�,�z$1�g۠y��hcQ�i��]�#R����R[,8���͌L�a�G�
�ow�3�O�O�8�qe�{��P���Y���nz�m)���&R���6���]���Q�ݍh��ԉ^�=��M�Cco�촻��'77m�g�ݟp��`�I�}t�����"D�TY�^��B�	�#Y ȫ�遥^{�����C�w�Ƣ<�RV�ĕ'�:�갉����Ɛ�m2�٥E40��3'O��?1���?�qɂ3�?a���� ��)���#q!K�A�A��g�?+�jN��-֜����g�(�r�ϸl��ADy�͖c��P`���gH�m_t�z�$�:��9��3b��5C�� *�!Fy��"�?y��M���0R��\{����dXdEy�l�,z�O���<���N6*e�]�CK�k�hpѦ��r�'<�?�����w<�@ �U�`Y�h#�@�pe���'�I���#�4�?�����l���cb��+E"��Z���7~������Ot�d�O��  �2�@\1OS�rUFe/��պے"O
2��5Y&䕲#�R5��k�~�r�vqەKG�E�$���d�1�|�� ��a^n����L���0�d����j�4o�˟H%>A��ـQ4p��J�j�	r���'���Y���%�����Н�@���3\OT}�=�TmL �ɲc���`����%M�b�ў,0r�'P�O�Q��'O��'ś�jۙa�)+�Q7ָ��[~�~�i���r���yش$X�&b�?��|֧� dиw&5hO<�%�2<k���{	���ƈi�X��ͭU���� =R'ܼY� ��|R?�"Pa�W{0�K��M���.B��PxM>�R�>	��]�%}�q��(�"�f����Vr�<��J;|���d�� �dq�eIqܓ����SW}�D_�`��i��0!�rG��~b�i��&�>�i>c�T�B`݈�E��.|�̜�$f4� �O$ (� �]�T�'úx��E�դ�%���[�=vr�Bpɞ/F<\j0M	�
	!��J+�w�&g�c4kP�[_!�D�O�~����{��|x��J#M!��	%'H|�9�D�	^�*�� ��42!��*�NI�# S<W�D"��/],!�d�|��mzŏ�:(R�<���ű[!��|&���4\VB�	��Ӑ*��D�n�I��/C}�<q�A�0�yREІN[ఉ�ϻb�N%��oL��y��?j�f]Q"e �dn��dF�7�yr�ZUؙ���U�^�8�C��yҧ���L�aB��23���J$�yr�U?S\Ȉĩ�!ZH10��O/�yB�E$ʹ�	�Ҙ!�0,�A�&�yr
_���� K�!;��1�b��y�晝P�|8J� $����e-��y��p��U)�F�=W6L*.�9�y�VR(FY��b��K������y&ц4�����Gڃ��h�N��y҃����dy��շ��!��ߗ�yB�� rH2$�S��oT"e#!�D[>'�t�P�a�'
!� ,B	Y$!��5t�HsA��4�Ʌ�K�Ds!�H`L}w+G�t��TI��Mq�!�O z���O2I��,)�#�/�!�SR{.5�'P�?o�� e�̿8q!�d�f��bjS�V�B�����?�!��Ǒ�u(�� <0F�t*۷�!�ĉ.�x��p,�-J ���Ƕw�!�d�29�z�Q7���:Fl��4b�j�!�D�72���'���c�Y+�!��r���1��%�* ���_VZ!��$���1�9q�����va}�)�l� hᢄ�2�x�0�c�[�0���M��8�$�P�w�x�+Ck��|Z����9G���D�-���+n��<�f,�8E��"���/�� �*l�6�S"n��M����H�Գ�ͺ;Z���'�1����(V�T�MO7;Gh$�u��:��R��c��`�C�F�[�)��4S�
�&>�3�Ҥ��>q�^$2%͝?nC�	���q��1
����
� 	!��.�� ^��<�`���}��BZ�	���e�>�`o��/�,Hk0"�:����E�J؞ H��T݊��*���^���^;Tԣ4	��@m����DD�݀�@�N������T�m<<��7q=�H��'?��[�O�=	�O��@΀9���@�I�%�pXFl�<�l��.�G��06��UX�+��u�$�gK�1|f�RdE��6�`�m�!x���FI�nCX��`��@�<��sZP��Ā�$&�Q�vAF�n�K�0�dϻ$gt�j��
X��CP�10�8E��*����n��~��Q�6�-�6m�-�=$��I����i����aMԺCï�:y�Z��?(�~T��'	� `3��:,U򥛄fÍR��A�ۓu��p��j_�/��y0�հV�&�	H�tg�](�gٚ>J)UO�5��@!�fކWr����`�3P�0�Y���sh�ipM����cM�Q�;U�8Ql��
=����w��2�X9H��.=�R�9p�ߨs5j� �c�;D�fyW�ǚ=N%��k�b1�D˖�r�v��caT3x�@�:�f���*Gh�-݆ `L�}%� Q�)*t�8]�"�ɁA�ސ���I�`�ްR��S%+ѐXd�̻~#�Q��L)\���Z�E�	��ЃXI�4ɗ.a����)hg�p��)%�x@Ĭʐ6ʡ����(�B�Fʺ,����jd�r��O� �L84L;kL�4�x�rG/��s?�sPD�;�8���	�cd�x���eͲ��Z�f�)ɐ���� I&Ʉ����!�Y��py꒦d�Ppx�k��`jH�>uz�iEG?ɰN�n�n�!"��Z0��y�����]��5�E'GG!t5���<�(����ѨS��В�d\"3���t�֢X�
�j%�ɯLA�	b�kP+Hz�u�+֨O� ��LT$N�~��gi��B��.H�b�Je��K֌y�X4�@�E�V��8B&,��H�`ň��œ
�X�He�	"gĬ|:�b�O����b�H:!����QM%W*�`��S��˳,Q7j�� ��A)7�I���38�
M�F
��sN�p��T-)~
����./��A��Қ<�
��TII�a|r �%Ivxj�*�B+��(��6R�����KDWT蘬O��"�g��e_ ��'�V(��ګts�0F�!,%j�I�nQ���燽R���zDI�:kl�"<I'MMָ(�B�|�d��%�s9��']��zqh��=[������$��B��-���cP�;e�c��
/����I5閜
���b6��J��_�$
\���+pаX��.3d�	"��4옼Za��g=��c�iF
$ж���[��e�k�t1ӕ��eD���倁�}\�����_Np�{�9D������@�d��u����c�!R�9�XCn�#���9A��8b%![G�󎆯b�z�Hc��}�pe��E.�x��oe�i���H�j���KY�>�sb���M�i�� �Y�CH0%�B���![�y�.��� 1�8+�ʕ
N�yʗR(��#>�2��$�ıF�-q�ғ-}����r�h-JM��c�$�*�C�L�*@�R���䋟:��d��CȘv��H�p_9�8��ƊK&08��Q�͏7Z��񃪒i��|"��(�8��0%��JGP8��&�5}�|�	�A�
Xh4Є�ĀNb�}�W�G<�� ���HCX,�t�X6z�`�Apa��<yԵkp��>*�ًq��)����ǝ��0>)�f�=����!AΛ6�����Ѵ��|�Rゎ�Y#*@9o�qk!JM�*1$����7���(�7��H�cC�H�#�$g¨5Y�N�SH��&>�=��PJ��[�1����`T�nI�e���@�Z�p4h�L��� eY���a4/Ԏ@��1�T��R�#�=���a���e��<�$ۨ2I��za�|��Z׍Q�<!�D�*4Ԙ�g��*v����(�*6@��2�AM�x���B�]?A��g�}��i@�-S_���1�m�����1N�}b��\:ayb�@<y_X��ǃP7:$� �f�F�W� г�eU-~: }���N3l]p*E^>�8�΋8ζy�qHT�����r���!���Q��.��	ab'�O�<��&)H���U�=RqA�Λ�d�0}"1��)vJ���PW갡z&�&GV��b��m≧L"��@�7t㸜�h �Vf@K1� <r">��ܖw69�jNl.��:0 Gl��a)�d���H�3B1��˜AI���@펩O�&<�'^�Zr��ku����dD
�ӓ	��&�� {��A�zO��п?���2"+H32�؃�D�eF�óI�'��'>e�AC^�<���WF��N��1A�G�7�:�㏈~a<��T�Sx�\iD��+<�d�3��/��-��'E�^��	�9F�p����!oq0�'p��� e�@��x�Zw�J� /B ތ�$%P=:���TLX��f�]����ib�� )��k�0�0$�`�X�#�J��ۦ�S�gB�P(P�K6�S�Zr(u�uZ�z���b��Ɣ�>�Җ[��'�ؙ#B�';iZ�a�$H�5�L@#eI��B|h����r@���5Q����A$�t�'$�����``��� !�I��Yo�~��<��ǭ�S��t���S�z4�U�7͎7iVar�
�_�<�
��x��T���Фr��}�����P�axңW#W�ٹ$�8vb��%��?M>~1�'��ԩ��׍�<�S�`r"Հ�Oef�`qo�X�N8�� �N�5!L57��)f`��0���D�1�@�%�A�
~<ȨA�K3:80"bȴ_1l�ش6b`)�ႅIZ0��G J�\�1FW�'�nP�&�&���P��D��؄�IH�� ҆�D��E�Xh�@Ά%  �bu�$R1�� dlD�	�rlZ��)W��eB��I�(U��IQ�� �Fy�D\*(�6B��W�
�"�D�t���.����L�t��/"L�0��Ɵ{����H����̮����KQ�e��Y�3ɑ�f�ax�m	]�dS�.�N��3��X��pTBQ)� �Z\�ֈj�M�3p|0�������
A3isx�稇��'�����;ˊ� ���j �jup�|���F��k��E�AYxp�,�A�<�d
}T����)�QeI��(G����Ը|��ղ���Q�n4�|�bA[~������ŪS	����N���x2�
�R@��H$}�S��G0{��7N7F��x����f(���ޚ�0<q�H�/_y�j���?V� \s��y���C�W�ym�z�[(@����V�.1�Q��~���`V�Bj��˗�2�t�*�=W�`����k�3	&?ɰg&<�B��	�J1�'
��~�q�|ڱ�[A�� ��K���X�Q#�K�<�%�D	u9�܈��ϴ}{H�;��U _=V�(G�-��l�ǇT�@nJ)�}�s
??9FFK�b_�,"5�P�t�,e�w�V~H<�R�ͩU8p��f�%u�͈F�	�Ҁ��B>dm
'@��l�\р`�'�̀�F��vh\��]�XBP��˓.������9u����1-Y�s�ͳc����m�D׈8Ō�F
<�PxbnJ�Y�>�`%o�'�2���ũ��Mf} �	W��iiA�W&���~�6�>$��Lx�_�
t�)*���t�<�S�N<L�8��"4^Q��9���0<�������=/TM��49|(+��L��z1Q��L!-�+i��㢢*D��y�L���Y�A�{Ѐ���V�>`��k]����'-LO�i�b��$Ц�f`���n��$�'���'�ǯ$&E��S�? ,t��E�0v��"�˓d��x"OR�J��+Tb��!%؜h�ZIz��W�ZZ%
{�Ox�����#�,x�%Ȍ%TxX	�'f�yR��1�6,�(SW�J ��'�r��V�	R��lk���(��'B��`6D�|a:���`ysBU��' 8���f�f���ul�l��1�'��q���$O�L4�*J�i�4Ը�'1�=3�H¹}b9+B>b{���	�'����e�L�[�q4MJ�vx~���'� mhu`4q��TJ�<$	+�'�.�Á� 9w�lL�'M��nH
�'SF(�1-�y� 1D+R/+��و�'��ȑ��4��y3�ɳ״�)�'����Dl]�S������ġYl��'�u��ƙ�x�T���"�3ɠ�:�'_n)�a���p6V���7!01�'B�T &"�R4F�J���8xG�)Q	�'~�X�r*W�%7����PN�-��']�M:c�$JǨ��S�
@��Y��'�4��� F�I�0�
R~�ģ�'��x۵+ި-��9! cG�NJ��@	�'TR�`�LR#-�(�P��<:c6���'�=����0QрRǭL�7�l�	�'�9�٘�.U2��"h�+�'��tSנٚ8���b��0J
|A�'ݰ�Ѷ슡[/ZI5�" �nd#�'h��x���b�ч��Vܨ�X�'��X*'B���Y{�lR�M�2���'<4x3�-�5���c`��D��h�'.VA���R0�u��
��Ew8Ah�'��v�@(6�HS`.ڂUղ�p�'��0ے,��yM�P�&�JO��'���P�T�g{8P��i�F���I
�'7�y�Ea)Er�;#���i
�'�F�HŢ�>B��u8���=|�\�	�'8>��/S"Y��X��O�<}lr�j	�'�P�g��[F$pAa˕\lN;�'+�Y0��	�@��*SH��%q�'S�-���B����m��B�H�'Hbe�	1��x����	\��'���A&�u<���̎�-0	��'\ v��'�:��p�Q�����'�68x��r�
Pń�LVry�'
�9i(M�a|����c�B7�m�
�'%yk�d
b��asŒ�.��'�bUP���,"��-�a��%�R���'��A��/l)�i1�M���^!�'Dظ˶+S`'����dF�B���
�'��I��C�9��m�gL��(����'�N�#p�c�2 ��J'<1�r�'�P	�R+�hQW	�6���'a�,"�)V,������rm��',����y��:��~�b�	�'���"BݎA�pu��ǒyr@��'�\Pp'măZ�^��&G���9
�'7���vƂ8GѪU��#\Lur
�'-�xQ���$��	5A\]�D�#�'�j��r,�%�@ͫ�l��Z)�'��QHC�9C6�jJ߮<J�'%��I���n"H��!C�`�y�'� ��萓O dŘ���n"9I�'��M�FN�W�T�ԦK�|��`+�' ����+m5�$#��q0�x���� h݈Ԁ��(��3ub�`�S�"O*T9c�r��⒄Y�u��@�"O�ب�E�63"đ�%�=u#�!�"OJ�� ��z��8P��ؚ|��p��"O�0��L1N�#qE�T�D���"Oh�`j�:0�r1�ƨK�
\�"O*�8s�͜]�F�"�;~8eۗ"O��B��%��a�� � ��ybᛄjJa`6 �:Iq�Uٱ���y��]Ȱ��c 	�Iy~`V�H�y���(V��s�OD�R�Z��J$W@�}��'^��Aa�*@G���@@�$��p
�'������	ny��e����@�
�'�\�ʠ��^Pd!� �RZ|`z
�'
�����=���b膱M7D��	�'�arU:tnɤ�Ӳ@�%z�' ƜP����J�d*DoǺ�	�'
.D�CI�68L�Uy A�8��	�'��9��%�ډ2�,J;RZ�`B�'Y�r�.�&l��Qo�C<p-p�'+R(;��հ?X@�Ӥ�ދrHhq�'G�L�����b檀3�Rn�J�#�'J���HG,_���S�
jޞ��'�&���"Rb9����Z�vP�'T�D�3i(]��X��CP�=�x���'h����C>?~�Xe�, Y��'�ȣ�?^�q(х�� Gdٲ	�'fȵ�ힵI��X�9"W̙�	�'� ��z�Аd	�\��!	�'p�T�G@X�K�2D�楕&U,��'{l����ܕ`�ڴ=e�U� D�d	�h�Q�
 �㙑%%�  �h?D��ˤ���\0�!k�,(`���7D�D�`F�|k�t	i�^���c%
3D�h�O�Q�DH�7J�++${� 2D��!jXN�x�beDF�X�ik0D����^8�����~<X!�H0D��ᴃ��d��Bq�ӏ4Q$ճ��/D�x�S�ܕ9s�E"���6�2��$H1q�����b?�`i�/L�$�U�H�!܎��uaLa�<i�K(7���[�aVe��yb���&���8!SAU�Ol�N^&j���8�R056^ł�h[�f!�
�4^LШ�OH�C��ur�$P)f� �m���)�w�n�(��`���UǏ��MC�1O�ʓ+�e��⅍19Ԝ{ҧP|B�㉪W���Rw�Y����w����U�+�8�!6@�6Б��OR}3B��Ab(�ⴹiJ�����`�t|c��V�P�\e�ԈչB�(!��Ȁ��3��5`���/l���H�i�'~�i��Q
B���s���o���l���IZ#:@�����YQ��'�=�f�1�N��y�-Ky�'��6mf�I�6`��<�+��<-�rq��A7�h4a[�Z K�bĄXִI�tBXnџ��$��Q�bX�"!�)!ٸlڒ��?H�L(6+� 4���+V?�B���Ɍxнxċ�} 	��S���"F��Z�����*^�<�|��Z�0�תۋ8��U!�i$8����&�/�B���]�h�!��Z��E�O����K�%5उ�MI�z� y���˦t[�%� �%AP�Ӥ����mH�MO�L`�X����'�V���L��1pG�DL��KBc�*��e�u��1C�p���$����I\.�As4@%?��I`T�?�O
�k����[dg�n���B�D)�O�(�RI2ed����nܬ�� �#��a���0=�g��	�1SsK��|@Duٳ)�0y��C��>�&� �,�Q}� /?�,��}r��i( ��ďǄ���<5��m�%@�x�f�z�8�qOz<滠���:,o6��
O��'��	���C�tIs2AH�WJ�أ�F޸@hn�8�'��Ux�,��0<�5
����O�����.��AEi���k�kOR��6��d�Ӻ�'F*���|��G��� ��ˁ1c�^�s��k�"t�@/�-D�-��Ir����$R7Kt�c���3�d	^�I͓�� ��j�� ;pd�2M�HPW�'��)������ �q��X��� ���ݴ]>z �L<Ch�~2��;A+�]�l�<�N�@L�����P\�Ժrd�~�'��+�*�i3T10���׎mٛ'T[��ծ,)dg���hAcAU�uO0�cU�ڒ�����4m�,�?q�`N�a�H�f�  N頒��@?)A�P�v��tB�t��Q4/�P�'�`��gídT `�[��<we`��
�'Z�P�a�е<e��T�L֎y���_�
\ɏ����Q*aЇ��/�󮚄Z��0��� �^|�@��U}�}�HЋ��H��eR4@��p6��.&���{�M5J�qO�<�׮
�2��䗓y�v0�C�|�` j���EG��9b|������hO�5��J&,�fГfl�8�n88��O6x� �̰E[*=���;�L��d��I�Y��!o�=���9<OnQ7�� �Z��b�ٓ`}l�c�3O����+l�<����nS3�5UV�R�d�>�H��*I:<ZXQ	�'�V1RuN�%�@�"ggG�Or��85�gYP�O�#<ٕꃼ!�NL �w(&���	86"�8C��Y8	Plb�$`��I�0�����3К$��$B�/"��B�`ؼ{q���d�NӶ4K�Y�r�D́�Bѐ9�E�:|�g�7zD8�q'�ŏ�A�O�q��Fһ�����@�/x�q�B7O����O�����8 D�����I2��U��+N�~�DL?+�,ý�p<����a�\�{ �^*HS�`���8J@
�r���G�꤀�n:���|2�x��H9?�ԭR�� 	��p�Ҫͼ�C�I"0���� �8]<�����d�$(�$K����&�HRtA|�oZ7O���yA/I�<��"�*y�:�˯O� ��$ǿ%,��$�?_�@k7�Q�?�JYR!�K'�H�0�&@���i��,&K�	2T��*Ac���y-R���lY���F�'���aÉM	a�65X�'%��L>Y�3G�p��Bg�>vؕReC�5��02�
�
|R� CL*� �i�Hm2�!��Z�* ���܅���W�l/`%���]������E�_�x���
F�
���:b/ ��U���4�j�o�AB�P�<]PA�����"����!+$���A�၄M�N���g�a>�������mS�qB|U;�/�WS�=��!�	4��'�*�i��Ԕ:����o\�E*�N�'����4N_8�t��df��D��T�� ��c)"t�H[V���{65��*R�_	��#�؞'��Y�u ����O�+��Ȯ�lH��&O:>/J��_���Ϩ\)x�+�n�c�
�9���[�`�˗�߫R�F�9T�i5�2u�
�uS�Q(�.@$T���*Tk�S�!Y�4JE����u?1��D��%-*��
(7�4�Gl%we�XԮZ!)� ���Z�[�6PsUB��e�*�=Ie��".��x`��Fa:\8���G���6�3Ola{'��RBB�"�lDN�`TD��'Yt��-���D�'] u	wK��y�^�)f�Q8u����)�E,8!E§�"�`��@bʗh��lN��D0vf�mp1ٰ������	L��[�J�&�6� ��/`�!�6Y~)���S<s=�Ł!��RU�O��Ome*-1�.�e��p�c�W�x����T��B?����)<2�0��\29�ux?�aЧ9\�y�Ɂ�+8��J�t�'۾�ReW�^)
���)�LI���	fpd��/��`ڸ�͜k[�7�<}>�G��FKp�A��S�Q�(�8�Llb��xX��	~�D�90/ ���XY��M����eH���'��i>��O�<�B��1	��%H�iDP��ŀw�^��Ǔ`I&dG�ӶW��<y�NR"8�d�{��vd�	y��Bʺ@Т�-}�*A��~���'-^�cC΋�|���$��iy�@.|� �HQ/�
a��O������Y&Q��F/}��<!�m��3
�iZ�O�3.z��R+^̦��wN�����w�U�j6�\V�'��q��a͡X����Zp��!	7�p��i݁���&[�p�Y�HO�T ٤	�HAA�D��tP%��p��L�`�tX���$:�n�".(2p�# +��7�F@��0I���D��1
�7V���<6��)�F8{��<x-2O��⣯�:`�(������<�0�Ut�2xB]8r�(�#��	����� �����)պ#S)��^�ҡ�0��(􆒰gb,�P�
_!�jm�O�Y�D�~�T��f�5X�Q�ֽ�d����1?՞-X3IԀ����h�O�W�ɢuD��'��d���I�wn�M��N��e" *U�I!GX^�z�Τyl$xX"*�R����ɧ�'){���r��V�;Ɨ2~�
A��Oȹm��}�;3�tT�bL����RjǱwSD�17BW�lFT�#o��"����~��Y(WE�(P�Γ�IG,�zF�NX��S�B�E�Y��\�>!	J^����#�	:�R !�ֳg ���C�R���'O�O�@�
DJƍ�~⤔�	����k�-t~(H�4���ēh�Q��aMҜ��6I0���~��S, �Ԃũ0���֎�v�D�$@/�bu"����+��
>�D}�)��3bM��A�n�~���"T��4+�$;����旘0��!@���)�)��+�fQ����+�yӥ�2\�y�fa�:��{��o�}�6b��W�0yX�
� �� 
bN#ʓ��O���� f4}�2j	<�U� ͜��,�RA+�|�¢>��IJ�NR��8�ǂU4"�˓'�� ����Z�~�(<p�*Ә�(<	v�?ғ{}`}�P%X:�9`�a�//����*I�`�~v=��ƧZ�d���@#P�����~�>�X"��$DG{�� ƈ�#,�<��C�ͽ�?qd�X�{B���b�T���)��@�'5��q@7��LH�����R�<X�D�s�"8�S��-4?ɶ�J!pQi �"��P�BA�,����'����A؈� ���.G���2�V,��˓:L���>�4 +��ڐ1D���"P,0���B4@�-Z���)
�D������h�.E0&��u�.��dA�*i�B!�5ڶ��ŨC�(0�QAM��~��UΟD�%h�**����:�?aЩ�~�'0�7%	�hPr� ��4T�X0�'�0D���Uv�(�vϒ	X�虎�O3�yI�LXQaa�L19��)2�ͰG4`� 8O���曾b3џh0%(�((Kr�_�U��5Y4m�A�†U��R�����>Y0e�����`�^uHD�g&�of$��g.[�V!��Ɏ~ck�iCp��.Jֵ�Uh�J�)�J��mZ���D�<��'LAX��i+��0CV��N�L�6jV�A���ڊA�d�z4�TP@dh��n�<$��6�S�Y��`�(�0}b.T[0�R$�剃�?��O��h�'��#�B�Ec(D ���ODI�bIԄ"π�ZNʟlBh����O&{dŚ0��eF��"$H� �>�����κ����̴Bɴ}K�#�-� ���H��[]Al�!-'�~�D{�ܨ���abQ�'�8	O˸f���� �P�qOF�>a�	țE�vp��_�&��@r-YV��[ f��0=���v�qh���c,x����`y�Q@�0�O�8�� �����29�!EC< n�����4\�ț�,�h�� st�כ��Z�Јȗ��0�\ܓ����$/��r4���'ݗy����#�N���_���8ia�V
U΄����X�+��I+S5R�p"�W/OF\3��H�М#=a�CE�rx�/���Ȥ�g�FX?����8A�$�c�±ɥ*b�'a�%j��ëg�9B1��3dR�Q�NN��<�xF��S�	5��kQɃ�f9<�� #�R�����勭<)i��
O��y�훍�y��/f����@�F+�"��Ox0id�(�$�~7M�nM �)syΥ� ���XQ���Ҍa�3��L:IbZɈaI�O�9b�%=[d��`o�i�X��W�l��O�払`'BͲ��i�0��iJ1V"�ϓ9B���SJ�u'�\���&^�6M����9�욶6��a�<a�f�G{����3p�lA'aP:ڪ�pу<J�v^�mh$hݴj1 �B�(��r�Q��Z�Ʀ}���óꚲ�ܡ㇅݋U�`m�s���p=a[�M�����nmb��7��\���;����!�O�K�%V���8�b@�-4������Ob���%��]"���6ZZ@q�c�L�o�\L��G�"u������<+�I� �'�^�I���$�H;��Qb|!e��%��}��'�4�X�	e,@b6��J�Q���F�E���#��
u�P������3��z�J��p�y�'F���
ػ'w�L3���&���cǋPhh<)gvK����ꌑd@���[�YP:8j�^��D��ɍ�!���h�m,��ۥ�yr��P�B�R46�`�b�"�y��A6w�PU�$$U
�l	E�H�yU/f��8F���K���#M�yrΝ�L�t�=H�#3�B1�y��ޘ$�
��c��,a��သ�y�	�""XP�%��:��
3'��y��E8T<�$y�R���:�B��y�#�����-Ե�j�"��1�y�틯r�R�˄� ���RJŝ�y���0o~y�sΊ�E�T�X����y2Hņ}'t�f-�p?�<p�㕫�yb��: �Pi��1`LH�"���y��H��*H�'٥-�P�ZƤ	 �y��"5T�!d�X ��pb�(�	�y�O^���gJ�	��x�G�[7�y�E�M]��aA8la��%���y�lU�?���@Sn_�-qzP��G*�ybl��_���P���2r�I��6�yb�2r�!���t�䲀l��y"��7l���Ӽj���/��yrl�[�P��u͆dD���y�cJ!��$�w�O�"�����y�I�G$	�vjY.=�v\[����y®��5���S#@�3�4q����%�y
�  ��'�@�y� ��W=#?���1"O^�e�6�h	�r�Y�"O2Ix��3n����HX"O^��nH%o~E��#���%�%"O�,J���xVzM��e��,�$��"O>��,*\-ք�p��)�~��"OtAs�{�����@[�v��ٹ`"O�Eq�J��@}�$��Ds4 �1"O���;'���ȴO��>dN�S"O�D��@�-fJM�4��S=��!"Ox�bR�J���2�ɺw5<�� "O��zQ�NA�����NT,��zW"O\rt�]H�L���=vnB�"O���SI(��P��"�0��"O<L[t�Ԡ2�1����^��x�""O�xd(QG`x(�-�4O����d"O���m(k��Q���?�&�"&"O�Yz��P�6��4iW�|�.eSf"OT0؄��)M�>+��ſk��Q�r"OP0Q%�Q�4�V�`�G>ly+4"O�� �G�3ʸ2��[�~Z@x�"O�)IGEK�j%��Y��>Xo��ص"O6���k<�zx�Q�^�~E��S�"O�qA�`�=���0d �!k�j�i�"Of�"v��s��z$`�\p�ؚ"Oƈ�%#��en BO[<_���E"O��AOI$D�0 �F@��Qtm�"O8Wb�3"J*TSC�VQ�؊B"Oly'$ġ?����R�$B�y�V"O�股+NAG��� I5#a�\�"OZգ��G��y�v�(oB�}��"Of���o�U�HR�Ɲz"�}+�"Oze��m y:4�1e�%I"O���&�и|�<1�%ژ;�4 9W"O�h�VOC���+�
D��,�$"O���S��.K�� �6��b�ms"OF���'��P�&1�h9�"O�`C6
ˤ�<l��@	���9:�"O*t�SO�b!Խ�e��h��!j�"O~� @,�9��Rd�s�)��"O�pSc�#<]8����%f�*ё"O���'a����B
�x�q��"O�T8��N�Y,~��D����(�"O�Q�ad
2U�u*b��IM���"O�-�g�!|Ҕ��]�%�du�!�$
.^�!���O�Z���"�,�D�!�$\�@�x���иu�J�9 �J�y�!��\wL��_�z��H���,D{!�	.0Y�@�		-��As5��.|!��>s#@q	p)[�o5\��#�Б!��2]+#�-��1TH��,�!��P��S"��E�ĴYV�ЃMt!�$߷(:L���@���c���!��'��C�CY�ag�EC#�J�No!��	�~��QK�`��k�p Eg
?pe!�D*W?<L����(2�u_!�$Ĩe�<mks�^0\� �� f�!�D�@hT ��뛶^(�5"�� �!�d��ax��k���3"ܵ�I��2/!�DR0�đ�Um:g�� 3Sȍ#!!�d�"������ kR$A��]!6!��ɭ�N�f��c�p��S�!�խ|	�#�P�Og��$OX�!�dG���LaT� $l�j!�� �aBר�$�8�5�Q�A���U"O��(`%�"f`��E���f����"O�|C�`�~e0Eh�I<`e��s""O��`v��2G����BW�@2�'���8ĉӫ[*H��+i����'߰��t�h�bq3c�?��!��'v����
������'�Ȑh�'-����i��̡3��u�@h	�'f��%&آj��}C$��ip��x�'�2�FٍRC&˓�"^���
�'-��K"�U%��QS�E��x��'ސH`d��(%Z��KD��.�Y�'��ᐳ%0 ���3���Մ�Q��xS`I̗ �8iZS��j���~�ZX!(�i�h%����&�9�ȓ5LP=�Wa��X�|JUnѩ �����+,���pO�
�Zx9V��"V����g�$�b���tF����,.�"Q��|~=p���
6ۊ�N �y�ȓ4g����� -����سS�=��dK��r!�ݔ��`���a�хȓ
FiY�ǀ&%F<ز̂I3ʱ��lz����H/lFXun��+Ҍ��ȓ	e"I�I�7,Ҵ�;`�V�^�>x�ȓ4���hdŔ��^�����HPԑ��6��q�DL�e�z4����Y�8܆ȓ^������s9���Aב#��ȓT�\M��U9t�~@C��MEt���7V޽{ ���B�� V�ٍETA��, ���v�Ha��c	y)�لȓ]�Y���U�7�u�AI��	��w� ��S��"���u'
.H�ȓn�4�dG�:0pb�e.jvq���+��'(t[EoƭD��\� &F��ޔ��'��5(',I}`m!��y��S�'SBP0 Ge���Ɍ�i�^���'�|1��Ʌ�f9�ܹ�+L�sA��'�tP�L[z�0��#&�?n��'����5�� *o<H�5��3(b���'�Ԉ mC7=|9�ߗ@*8���'"eb��d�6%J��<��9��'.&uy� #|�T$�PK�1��e��'�̛�/���t5r��ϙ|X��0�'���ĩ��m���#b�Īp����'�W�溑�Q�� a��*�'�<�r# ��I���Ċy��M1�'�L�т�G����HT7s�8��'�X�Y6���8G�`���7PX�
�''Xi��!�R�r]��NF�y���'x����d�s����b1f� eH�'�Ti�Wd�F�h͓dI�?d����'�<M�g��5{��A�\ b6���'�h�T��jҌ�;Cl_0V���c�' t���P�xj<k��ok=�� �'V2A;��J
�0;��X����'*���kRoT����	�-eP�
	�'w�=�'��X�9��g�j����'4"�d
!����߼p{Z 	�'����a�ڸ?~�a���։y��h��'��H�bi�I>��)];z6$  �'a5q!$I�F���ߐd�A��"OP튢*�?jMZj����ڄ[1"O�7�͕laH]e�;I�$�"O@��7f��M"���B�5(��b"O� �{ei�.�Ⴃ�
��Q�"O�0�\&u�����-b��"Ot�д�
0�lP�򏃓�\�"�"O������/p��������"O�x"��݌��!e��4^��<�"O��JUO��>Kn��"�(�8la�"O(P��'ʺ"�4eٱ+���-�@"OΘ�Fjػpv@|�*}�$mp�"O�uJ�>T�Hِ�H��P�����"OT!��Ʒ_��3HE���E"OM2�i�$|�Ĳ��٣�@=+"O2�9u�>�Dd�lIe��Hh"O$�ㄒ�W�4�e�'��]�d"O�Ă��87�d�K�gV�V�
�"O@d��O՗[�\�G�	��2�"O�Tb�hT�������>�^�9s"O��4j���#ٿL�䜩�"O��D���i��WL���Ղ"O�q $�=���K[/KD�X��"O~��!��@�\A�kF�J'�E��"OB�p�	�>+,�I��4l@�A"O|�1��U�
�ѵ(�G���"O�ԧQ�]�`�p��jψa�u"O2DH�,~��"���!(�� "Oڡ	��\5f�����7#4m�A"ON�adT�G���;�U6��p"OVxpF�x3�e���'Qƥ0"O�|p����ȋPDւB�{�"O�8�`߄2 TI�C�~�V��"O�E���feשJ�e�4!�2R�!�G6�, ȕJ�o�<Br& ;0�!�.q�ds6,��p�"HP�b���!�Ǯi�x�Q�;k t�����V�!�䏂{�j����:^	������?X�!�$��oK�y�Ub%r��$f�#!�$U�(�\\�">Hɺ"'��`!�4y$�8ҫA�S��stmF !�D͘vL8��$J�<�\�I���*U
!��E+��`f�˹j|@H0�Į9!�dŒ-�\�����.xf8A��V+!���"'�6 x2�V=Ⱥ5��Ļ�!�	o���+2��2'�TA��Rq!�ć�^s����oD2����Eǖ�=S!�$X�w|d<arˎ���AU��GH!�$M�/(���g:j��y0�Q��!�$�A�Y���	3�y�cاyk!�Ğ�c{t���I.q����DY�1��D�;~ң�"Q26T�a�H�y�b�4"�R� �R94x�� (���y"��"]^��,�<� ����V��y­V!*y��.}�U���Ů�y�-F�&$�e��̎t� ɲ%�\��y"�I:�BqC�KH�X�^da��
�y���$*:(�q�e'!"�QeNI��y�,Q2r�#���p���ٵ0�y2�B�U����&L@�f�bf꜏�y��Y�$��E���MW�j����Ň�y��	���ɑbi�:gz$��	� �y���+s(iF��0'�ZԋR��yr��%sb�K�l��)�H�N���yo�(	���K0`&�ε1�$��y��U��i��m�+��c�#N��y�C������`�`�aw����y2!^m��Rc, 8-��C�gɚ�y
� ��!G	��]�m�e��W"O�D�$��"+�8)V��SP�]8�"OI�-�tϘ���Y�'=vux5"O E��`�Ux"��ǲ<#�t�B"O�I"�ĉo�Š O_�{��"O&|�'��<7���e�ԧO(�A�"O<�(t�ӔIZ99wL[�r����T"O�1c��l��,B⛺$�ȁ�"O ��'@�f��q�E��/N��\��"O�r��7ٜ%3pMR7<��考"O|��e�� K�Uc�e��#-�\��"O�q� ˍ�Qh̀���s�ɫ�"O��XDM*Qe��+U6f���K "OV��׋�lt�uا��jq�P�W"O���m&_�d�{�,��/fr�$"O�]CƏ2M��L��lU7J(�0�"Oʴ *�V�p��TF&i���!"O�yr�c�6�ּ�GV�Ry�ա@"O�E8�J�^��zW�G%o]�$��"O�\�o��	f����N;O\h�`�"Oj��f�7G,&����3f*FŪ"O6t9�/D 4�m ��[�s$��1�"O�I؃#
�l����ृ�U\���"O8�p@�S���I�t�O>�34"O&5ل-���x�R��?2���	4"O��� �:k瀍@R�C� �&�i�"O��`�-��h����Hò-A�"Oڬ�f�6��g	�� "O�i��&r���a��� �P0�"OVT�� �2�S�H�`P�9:`"O����Ȓ�c��*�{"OZ�t%)V�Z�=3pd#c"O��'L��y`}"�σ�O3��!�"OD��ba,�����
�g�0Y�v"O���ױ W��	T��vYlYD"O��JrEN>#�(Su��/IT^�9�"O\(��I:�6��$�+rQ�x�E"O� ���U+&2�!���F�'I$��#"O$M9�k��T�Ԝ`��E6]*��I�"O�UA��	0hKD�ː�o?�x(�"Oz�)Af��f��V�"�Ԅ�Q��y��ϊ�ʑpIދq�����8�y2H�%[6�����*q�pY0���yZizt|@w�N�L�u���]�"�RB�ɨ6��
��Z�.����o]�+hfB�ɔ&~>�B���)JǬ��P�QdRB�	�!�|؉P�A*{�PU;w��z�B��8Vo����������"�""O�lYw,L�7� ���M*8nHv"O��(�*B?o.\a� &9#Ը��"O�p�Qݭ}`u��nK���"Ov����M�L�b�-�~�LИa"O�5��	ȕ4QZ�`M�G�ڨ"O&��@�Q
v����GKð`�Ap�"Oj:�HT>2��&�Efl93"O��pf�[��}��0#b���"O��1�)t�p���N$,U�k�"O	�P�I�#դ�w�E�X"4�X5"O!�BA[��9#"N�4�@�"O�̋�),���8D�>��p�"O`�R-��n���
���b+,�h�"Oak��Z�y2�[!U�/̐;t"O�L�m�."X��N�e�)� "O�X��J"%Q�� K�;)�<e�p"O� $ Ch6��� �V�eL%�"O�Lq@"HBft� �g��a� ���"Of�8�*n9< pw�'�`@)�"Oz��蓍N<���	jRpm���	O�OT2�`��&	�h�ꁝ���
�'ux�	RJUv�����
�X�q	�'� �ƃ�<^d 2+�M�أ	�'��Tc����bj�i�AAF��r	�'D�Xn�7EUL4��Fަ|d��	�'�:��BL�&���`n�
��3�':�i$��F���4y��
�'�T����N�V�ZA.�n�pp��'��U�NǷW�P�piT�����'-��I�%ba��C3s���'����(1�H�K��Z���'#6�K#��7UӺ=�1�@=�0���'V�����(Pɨݒ�V+�<�C�'�(,�@m��F�!�CЁ(�V��'� ���.1S�ș �F�).����'8H��$	ݽ<���CiX"S�9[�'h��
+Ҹ<���P�D|(]��a9$�l�C�gV���#	U1�P�`2D�t31��2 �U�3��8_�(��:D�@�6oV	���5�$��b7D��
�=����J]7&�!0��(D�P{GaϾ8rAI,H�E��F(D��*���p�`�Â@�J(�A�	%�	T���'c�d��"ؽ<��тpdO�S2l��A���fú-0L���
�Z/�	�O����	T)v̙2e8̥r��]�!�DO�~��s���)�$"����!��̀R;�a5,=6�\�:�� !�_:J����=�,�����|�!�$�=x�v}��J�x*xs�CN/:&!�d��p��AF=Qf��p�"V�N%!�d�"R�p�(��9-���\-,��(�S�O�6�" ��Z��'S��	�'-�����4^��K��9�V���'����f�9��Ѥ�hݤi��'�؊W"L<N.x�p�]�01�']d���ҫQ����m�)\�p<��'ZN��	�]B00�%ON'>���' hqy��Z�?�b=��-PN���y�,]�6�tQS4!�4cA"!{j���yeM�,*����&r�ʁ�tL�ybN�}
h0�4nT��]{�	#�yb
��2U���R1u����d���yү� Y�X�!�(�e/���f�3�yr�U�T���p!�К.j�Q4Ė��y�*�*2��Y:e͝�
��2ŕ�y2����D2AS�s(Ӳ��<���ƴ�i�SA�	AT�qp�B�9�!�d� WFb��ōU~�r�ÁӉx�!�d��?��@A���#��+�!�:)�!�D��p.�T�M�X�~�Ӥ�ȹ5�!�اbjZew��/p��҆� ^f!�$Ş\2�0��(6�8��GA�Q!���F�������7Q� �N�!��ĘO�r�P��#���B�@�t�!��!#�x�P̓}�T��O�$!��W6�Zf˞��_�~�!�5o�� g�>Q"go�Hf�	B��H���9��R� �	�.�����"O�}�A�5x"��toX
1n�`"�"O� \�zG�уTu4P8�tS�Z%"O  �a� <&�b��ǝW���"Ol1@`��=R 0���HJ�P"O~�0dڂg(�����n����>Y�?�b1)_Q풩�pJ:<�h�"O�y	��A=9S���'�`Z�4�"O<�A�R��~aq�ؤ+E�Qۃ"O���*�;V��h�G��!ޜ� "O��� �\{�I����i���"ONx�	�+p~��rVK�8�ZI�s"O<-@�D�)�� �c�O�\0�bu"O�Mۃ��Z2j$�G�:1�
�"��L8���V��~�J�'Z$J&�-D���7MKQ$Fq���
�>�H�+D�`q���'!��%s&�ʩ#��*�`=D�л��RU�=2�
 ?I���2#;D�ܙ��Q�<:pY�v.�;EF��;D�l����P�I��$XO�v R�,7D���P@B�������`���f�6D� �/
��`��#'�t%p2 0D���6	����Y��ѩ`\`9pR�>��	m�'� %�V�1we}ŇI�%q(�r�'�i"TF	 l�M��dU��=@�'�DЁ�H9C?Uk��`@��'Z֜��,Q7OaV	���%g�X(�'�F%Ig&�$+�3�˟Z�\x��'���U�X�ZFn�k��F=�$�
�'�n]k��9J� �#�;}6��
�'��x"�� 4�!�H[�@&��	�'6 ���;'Җ(�&�N�I���I@���L>�!d�/d��b�L�����
[�'ma���ՍV�����)3DR��bk��y�O�4��U�!��3�_�y�gZ�.qR8���_� 2�Af�<�y�.�5��%���|�J5�ѡ� �y2OW�+�1:B�C1N��NO��y"1�� r&��g��\��+R�y2�EH\�CP�[S"��B��yr��.-�����Dz�@h����y��S�C�-	�M�s�F�x�D�2�hO���i]�>l.��V��A�a��(m!��i� ��r�)++|��W!V�kd!�D ��	`��9�ݡto�KK!򄐃e�ڵ�E��X�@��A�'d!�ĉ;Mm� (�t�^��!dZ�H:!�D�6(��}!!(׭^�h�d�2\}!�H	[~E�iԬɞ,Ic܉"f!�$�,A`P��b�K�"��5!�d��}��eÈ�r�b�q!�K�!�Οu�8	B-��dX ��� p	!��"݌��s�G:7�����]�=�!�Ӂ+Ԩ���<g����4� �y�!򄍒n�-����$<��P�w��h�!�d�!R���#���=����q�!�d�'`&L��U_�0�S��q)!򤊸{�S�����q�P�^o.!�B�/%��c��
�&HIF-!���}�p"u�S�'�Jm�6Eǉi!���P ��ŨI8hTȐB ��,�!���1`l4PkӗbbXU�"ƅJ�!����l�[��ݵmFlqo�Q�!�B^�������.����5+`!�d�!��8j@���LmK���M�!�ǆ7Hۗ�W!d�4g73�!�� �鳥 \�2b�IT��QA.�	"O,L	�%2a��Т�OHL��B�"OP�õ!\�'t����طv�Ja�!"O���Ҹ6��ТG�@��](�"O ��`��q�ђb���@��8S�"O����8ݘp(U{g԰q3"O@Pr�D�a*��"��0e���B'"Ol�`@�K�Kg�8�� /j��"O�����_�DEC�ㅿ6O0�Z�"O�IB��1`-"d�B#<� ��"O�Qc�	с$�LYReY���̂�"O
��~����4
fP�P$"O~�U�A� �bl�(	AL��h"OB�S�ݬMeH�*��V6���Rd"O^��H��R3%�-b��B�#µ�y����J��\s�'S�\6�a�F�]��y��yGT ���
T�jj`�2�y�l�3w���vN?FN�i2�fͫ�y�i�^𞰺��J:8��R�/��yR�C���	WCƑ/CH��$���y�B9Y�P��.ܘ�aE��:�y��J%7��I��悘PȔ=�1���y�a I�z�ؚF�4yѠo�3�y2%E>i<P��H��BE���	�'� �	Pǂ�".�) ���= q����'�L�! CB�A�d�A̊q��x�'n��Y�� ��������rTa�'O��*rJK�#���Gm�$v�j١�'�0���4��iÂ͌�fo��B�'�j�K���@�S"���gbX���'gP���ΙGf|�s!����q��'�6 ��o�'}� `��	��*X��'X$��.�=iR]�ah�*}kP ��'�p1��j�nh�	��M�vJh���'���w�P ���
�?��-;�'Ef��f���#HӢAt���'".-a#�:tUn�N�	
DEP�'��Az%�\�a�R�Q�b48�&��	�'꼱¢Ynä勰�?>kz����*���,5�Tf�T�$r��/!��`���*/z�XC���;� u��Jۺ�0ǐwMX�3��َ��s�h�
VIH0;8l{/ьaBɄȓ#�1"���s��}�ajý6�4���$�iٴCG8��eCaDȄZ���ȓ7S��3�(YQ�Lv�p�$I�ȓ37(-E��5f�j�:C�� ��\�ȓ���t8DF,yz��X�x�ȓb�:��TD �>�p���uT���ȓi' ����%m���x׉�4)���ȓ�xL�獇6� pr��2�T���C�t͡bK	K<�$(T�1NUhĆ�B �;B�.4�hpR�-�5%�HU�ȓ^�&�ZFX�C�.Z��%��l��Q���z��es���(�hU��E�2��Td�:A�Ό[V �'cb�܄�->�[@�UE~j�q��i���ȓ,����pf_��=�i��C�<�gɮ0��}J��I']b� ��&�~�<�f��5$����υ!	p�Q�G�`�<9$�\;b���	6���v��,�q�<�c�#QNM���ʗmh�����q�<�&��2;�!���bM��Dk�<q7a7,j�|!����kE $�С�d�<� l�8DNښPI�4�����
��"O��b�ߒ���	�'���!�"O0�3�Q͜�jЫ�7U5�h�T"OT�ߎ�	�y����\b�K�"Oe�$jWf�Ux���4,1� ��"O��Xa*xz�x��܁s��e"OZ�
��ߩ[��)�0!V�ӗ"O@ؓ�bY(X�zٱG%�$��z�"O `�������pD��0����"O�%��n��&�,]���{�8K"O�q8P����A���9'�"<S�"O��d�8'E!�r O==&@p��"O�@��O�5v�ڄbG��*v�0"OJ
��������L��$��"OB�Qf����X��EH�<uR�Sf"O� 	��Z0Q�����F5S�Q��"O�,��8N,Dp#D��V�]�"OB���U�!��C�e�&�V��"O"E: ��0q�P��D��[����"OH]�v��B6�kTd�~�H�G"O�S5k[2k� ��3�.S�tY"O���KҼXy�jpBHe����"O���M#��*�9�z$a�"O�����b���ȢH��"OL��kʰ.~�R�c���"O�D���R(���hP��F`\娷"O���a�@/~q)���Q&%�"O:|�"��3}~a��e�Dt-I�"On1��^�`d���v/�)-�H"O��X���$��i �
wB��"O�t��eߥZe���`�ǫk6(�"O����$�!|�@�׊d�(�r"O\��!	ҿY�N��g�ׄiMf��"O�d�3`'$
���&�:�"O����"u5�<��L��@�4L��"O2�{�W'5Ēp��-a��:�"O�a��F=}C�e�d��N�`�"OҠ�)A#{�D�#��>'Ŷ���"O��Ht`�b0{�A��i�Pw"O�����7o~��9�E�����"O~(CL$?ll2��х#���1�"O��[ab�o��+�<	}��c�"O�(��(�,�Vq�DL�.Z��,a"O��J��F��:Q�ǫ�?J�b�"O�L)GE��h�@���遍$d*� "O���d�G�6rN��sH��sxd���"O��X$�͈tx�K�&�bn�q"OF��rA�F<� �cfR�M��"O��G�R�q��i�ע��L �С"O�ѡ҅��{�2�1��*�\|�d"O 0��7[@�
��G�z�]k%"O��Ö�2x��xP��,t?�YW"OF�A�c �H� ����e"O>�� %<�F�C�L�6i:T�"O�X�#�oZ�E��P�EM+^S!�䝷f��0IaJ
O�kU"ֿKb!��"^Z�\���M�@�~�4"DCO!�%/� �E�31:��!�<!�+K��h�tBJ7�N�;s�M"!��tv�y1�(��
�@(���%!�+H�Za"Å�;|��y�.�%!���B85k
)�
d�`�2�!�D2T�̅���I�pأ�׻K;!���\�=�G�1�h���k!!�� �A
 �pX"E��h��|��<�"O!�D�٫P%<q��'��Hy.��F"O��a�%P�mN�Pu�0D���q"Oh)a�}9�`���!<>�`e"OT\�A��%R����j�;3*�Pr"O����F�1i�����F;�Z���"O�Qu)E�M�%��Ä��4"O����=0��E��%b��)@"OX)�������d�%yOrxz�"O���󢍃j���w�KK�KE"Oj Be����I��bX2\��V"O�HR��Z�K	���A��fb2"O�eá��=}|@cA�C"�n)HV"O>m�%݄cUn�I�N M3H�E"O����%;F� peZ����""O�	㲪Ǿn�4D1�
���)Q7"O��#�IW�V�"Dq�bF�)ܸ4�p"O���2#\�C�-3��I?&8B,��"O��"�G��V!�t`�	�B>Ȕib"OzP�4���Y�iR�ʉc8�z�"O�઀��(���#�-W�1]ؼ�T"O������W-��0�K�,���kd"O䍢���'�����)�p�b��C"O�H栕�����C\)m�D-�"O@��wnZu�BA����&~����"Of� �G�*b�p�R3�G3&�X���"O�A�f�خ �2u��ܩ(�	�5"OZ����*���:�O�'>jT!A�"O�hYg�2[NYД)�{T���"O�J��[xan$C5h�7]���"OH(h�W�;���G!I i���{C"O�<ib�Nxl���A֨��"O؀a¦���0���k٪t�!y"O�=��搽!c�� �P2b��Y�0"Ota�w�����/њ��L�<	�%<?�m1�]�l��JB,��<�wj,�*Q���>`F̱� �|B�ɡE�J��U ����:f�R2#wRC�I�\* ��HO�����E�Ё76@C�ɜ;���G���x�P��~�B�	�CG��(Q��#A-�x��J�A�B�ɻ'��=�E�"G�xg�].dB�&}d���Dɓ�7~������B�I�i��3 焮0�h���0;��C�		y�,Pˀ!<�q ��?2���d["~*�X6�+��`�$�!��:Q���b�������Z�nH�@�!�(�VH+#��C�<8��CO W�!�5]lɺ!��be���(ͤ%j!�$ő-��t����
`p3���2aQ!�$�a&�i��Ð)I���I�
C!�Ր^��Z���3$/��#��B*!�Q���{��U3y�B��#�!�䌌������$W,�(p"��[�!�$TP�U�r��6tJ���,ٗ)�!�D�=f�z�����P-6\�JOX�!�$(d:	T�%��󨊘;�!�d�c��K��T.I�ݺv�ڑFi!�ܔ=S|���\8�
L8���m!�d�|�����c��X���TF�,R!�CL�b��w�!4�B�c��O�!�D�m��Ɇ��!�\9a����!�C�y�lp�FM����5Ҥ�ƱR�!��N�u�p���X{lMZ``	�"�!�� �t*���!��(N�ށ��"O`,���	��ē�+U*o�N	��"O�p�S@̙Rz>	�f�͊cƌ]��"O �;��\��>i��/^4>�$h�"O�*��ůG:�Y3�퐦!҆�R�"O���D�+��`xp"N=S|�w"O�i1뒧-z��'�����"Ov�У��!h���S��;��p�"O�Y���TXb�mBt�
Ak���q"O�(����f���s��=[1�5"O$9��,���!�mL�6pҵ��"O<1K�fZ>d��QJ��͋z\�t"Od��b�*�X�h���:5C���"O��#�Ȯ|�Tm�dG�t��!�"O<�brM����]��^���!�"O�<���#[{�+'�\l|b�"O:|��g�B�*<�T$ï`k�lQ�"O�y�D�T�?�ʠ��I+Ck��4"O�Br��?�U�q���?Lb�(�"O���2eȋ5����Ӆ^!>�څ�3"O�t���z2��Ҏw��T"O `�nś1��D�l� -~�|R�"O��{�*�L��XP��Of�s"O�����15�Y��B�R�|X6"OH�S���	�$HFk��:��Є"O�H�GbY�d�"	�3�Ծb�ȸc"O���'M�J.�3Q�Ƚs�.�Z"O>�s�&�*Uv�P����7� �9""O���E-H)W��Q�/X2 u8dڑ"O�LX��s�|��+X�t����s"O����X,Aq�ڵ�r"OF��2�Ƶl[��(aHˢtZv�q�"O�`4L�5:|�zԨA 'C��qq"O�@�E�IlY�F��_10�1$"O�y��S^^ �$fI�Ur�m"O t�S�\�Kʼk��}f@�`�"O��錻Z�t	%.�nQ8�"O:�Z4�@�%�>��q��+�>�8�"Ofah��:uV"�ֆԉ]��(`"O"��D�ge �rFY:8����"O����G����䇐3�И�!"O��Ai]:g� ,�d��74� A�1"O� �a@�*j�Qi�S-=KJ%�s"O2Y���-��8E�M4%Fhi�"OF�1U�G����D���9 �[�y��U,V������R��Xg#C�y"�� ��	Ǧ�P���6!ͧ�yRc�/8C$5[�ӵG�l(z�8�y�m�>W�=��;� �q�i§�y���1^	p����-�v�)P���y�nO>q�<������)�7�%�y���2��t�Cj߾1���W$�y�$��l�DD1��3x�$঍ş�ybMNn>B��!�"[=��B��[�y�ߚfI\<��H��U,0p��M��yr��F�h��!Fz�Z�1�� !�y�K�딕�ui��s�0) �A(�y�"JU� �aw��=Z"u�@L;�yb��Y�gƋ��ع篝��yR�K�%_��9�o�h�T p��>�yB/�8uߺdQd�ħf Z�r%&��y�	P�t��,�$�	+�y�����y2�ſa�L�:�M�jib�h��y�a�x�(⤦ض[��1��-�0�y
� ��	��jQt�k!�J<q�m!�"OR��W:hu�x��޼#�Z82&"O���� r�Μ"a�D>$T��w"OX� 0Iվi;ΰ���I�}H�"OT$��%#n� AM�69�<"O���� .�<L��¼f�VU"O���B���@� �AJB	biCa"O�	Б�7���p	��*E2Ñ"OT��fh		�N �v��0HxJ!"O0i�2���W��"&�<%��"Oi)2��#H���5B[�B�9u"O̝�V�
�X?��2�Jڵx�~��"O`c��I�b+��1�BH��B�"O� �gK^��}*B
�Pج��"O���I�,T�pĪ�&N18�*�P""O(�0�"G�9�X�Yq�޺4��, "O��S�\=ĵ��jڀ9S��:S"OJ)�����;rj��yV���"OXA�$��7\���2�OI9K�P14"O�`��eڕ%4�0�rY
5� uچ"OR�V�H��\��`
ә6�\�Sg"ORm��| �
��P�K�F01#"O� �4��N��U�A�FV0ec0"O��IT��>u^`C�m��JI+E"O�;vH�!���A4M&�Y�T"Od� N+ �a�!,�n���W"O���0,M��0���k@}��#T"O�U�1AF�g�~eȱ+Z1l�v4��"O���#)?�ޕ�A�K�v�P	s�"O^P�#G'n��RD��w�t��"O<��g�F�}".�k#�|��a�"Ojtaį6J"�t#0AZ�*���2�"Oh�pB �2_�8�A�1p�l���"O��	��"(�"=b&`�!�45� "O$� r�W:�8��0����"O9���0VD��k�nG�"99�"Ot(�T�0]��)�ƍ��#���!�F�@Up�
��5�DMAB͝�w�!��ֈ6�&��
�'*�)V&�=q�!�^2w�¨����$3
�p��xݴL�ȓ'�2��G�I-�9�7f�x(D��]��p�UH�fn��ȆLǼO��Y��dipa��OZ" �����M>ؐ��x7��*fN�+2ھ���i^�% -��@F6���,D7[�i���S�Whx��ȓ��D0��&�B���w�U�ȓ2�e�` ٬J��0bKK1d���ȓ#A6({S�CY�j�c�E<v���ȓz���c��q�� �6ː7B򢐅ȓW�v���ĬMo��js��:�Ҍ��%����@b�NV����]����	(.}!s!��?�ư�b��"�̇ȓk��e/$6����Ɉm��}ɲO�z�<I����*�9P���.zb��P(OQ�<!���?y$� �'�(OO�㔃PH�<i�	�f�f�Jq��,`��� �AI�<QQB�� �V�kp��+D#8"#�J�<q� �Q���EA�[�8mG�<��o\�-��9��i�P1&�1��]E�<񀨈U�0�%��J\b�qJ@�<�fƨs�ZP2�e�2D&!) �OP�<��b��A+TGX�{��԰`�S�<eB2@��+ԭ��F?��3E�N�<�� 5qr�#���57�����DO�<� f�Jm;-���Z�&�wJ}�"O�@�t�L.[��a���G{�d!k"O�Y�u��"h� ���K�W��uJ"O�UR�E�j�b��2H]	�`@��"O�ЃcR������v�J�r�*O����׮,�>����WF8��
�'�ՠ�L5!�^��c&���E�	�'@Fܡdʌ.u��;�"�;��ղ	�' "y��̧4��icaF���"��'Q�c��]�J}�#�0_�PE��'�6���ުqz����@�Ysz�P�'*u�C���K���+g�йR�'@�W���`U<Q�h�d'Ȁc�'=��	�gƺd
ɐ���K�~es�'��d�Bۗ@BTË�>Đ���'������69���� O��dż;�'�d8�v�П*~.0U�&:����'U<P%%�D;�,��HF�6����'�� �  7���B�����1�'��-�'��"A�h���Ջ
�bu��'F+�	B�I�:\'��8u�r��	�'��` ��s�*��*�!8�x	�'\�E�P��,4.RPvE�1�rx3	�'/�K��A�]�R��)�z!��p�'�t�k[��r��d�mq
�'1lXr4K.�$�sR"����Z
�'�V%�u��?�1´ 9eฉ�	�'�ƅ����D�C�_m���	�'J.���ƄD��`�3O�&����	�'f�3RMZ� ���X3��݂����y��]7J�$�ŬO(+'x��VG��y�	
W��1��K��p�;�-�y�X�{����G�Z,�ѧ��=�y�%�=̢��#�R�!�pǧ��y�H��51�U��	 D*gK���y򩕱u��݂��:M���pCT�yr�-o��4����9K"�K�/�y�cD%o�؄�/�4Hp�ʦ�y��Ўf��X�垒 9���d���ynѓ�dع���K���凷�yB(��`���v�@��Kϙ�0B�I�|��j)q�mh�.͆_B�I��P�z�0���ٝG��A��?D��a�D��V7X��*�"D˺=�<D�h��X�|=\�{����&���$�8D��C��= ��4	���ހ��!D��b�/�)�FcԢ�'x��A�>D�x�GG���<��C�U�l��N0D��@��$;L��*��x����0D� �@�Ҡe�0���?����9D�� �M=
�x��定���YU�6D��"����=��0�S�F+B~nM	��5D�(�G���TThdcP�U��C32D�ta�*'b��iϗMcܨP�!1D�x� ��-u��y��%X�,����5�.D�`a��ĲIf(D��V�EX��C�/D����b�$r��A��^)J�c�.2D�pHB�P�W�������p�|\�q@3D�lQ��ȦR��B̛*PeD���/D�����U�F���i�D��1D�/D��
5挄.��9a/�$`/�2��,D�j��AE�T�j84��VB,D�tQ���ڍ�R��&0!\qR��(D���d�ǅx\UF��L�n)��j3D�� <P(���=g�`��W*$�ԣ "OB��SįX��iX©G�q��x	2"O�I�U�5�b@��̅]~�؂7"OlP
@E"�ذ�0��<d�] "O8:&/B*v,��4-�4H�E��"Oj�p�� ,��$�%� 3�"O�	"'�+Ps.�0J�<%��t"Ot#q`H֌p{��������N]�<I��)a��Q鴆�>��Q� ��Q�<Y��1"F
��M���ȶmXu�<���4YR5� ������(L�<���߽r���3��A��q���F�<)��!��pF��� ���օ�Y�<�V��"0���p`wH����kp�<)0� *w?��{ Ɍ�q�p�,�@�<y`-�?�������&u���
'�p�<y��V�w��°��h|<Y��G�k�<!���	$<�1�PCP�q2�I���j�<Q�e˦0y�=��Ҫa�TA����o�<�C��-���#�U�:teBqB�k�<q3t��B�ߣ�����\n�<�@"����ٳ�ѝ��ŀ���j�<)ce
�(c�I�2O
"�D�Hg�g�<��o�'n����G�s��p�FBd�<90�Y&J+B��lG �^��f�E�<��/M�.��a*��T221RF�OE�<�rHS�}or|j�Zek8 *�l�<����'��tOO�f�2�����<�Q�����8��˘�j�������~�<�B��26�ҷ/��}�1s�z�<��T�_�h�
ą�	k@��b�<q��^E�AʀÊH������`�<a&��rc���e։_��A�w�<q�ӡ(D�!�	�0�(�1�t�<Ac�I��]��S�&Il�(u��n�<���@�`�{ G��w���g�@o�<!��W�_׆Q(QI�k��E��R�<!�욊u�b5��/]���"1�BM�<����;&�nȉB�"Wƴ��&�Os�<)��@�Ru�m���`��m�R��z�<	A�|��@	���f>�����x�<�3�L�2|�sBnH�r5�����o�<� �P�~���F;`��e"�A�o�<��*9j�8������i��i�"�i�<1po��;����hC29�p����g�<)`�ص_`iS��� �d� *�J�<Q&����<j�0�:�P��o�<�C ;kc��#J ,{�4Ђɜk�<�'�7{�PJ��VA�H-xPJ�P�<�D�RQ�@J7`��9�`�IYL�<IPk_�נ%��^9�1�*Nr�<�j@LIpsf�lľ驓��n�<�Bm�c��@kpB�
c�JQY�fj�<A� �v6��X!e�)�鰂���<y��Ճ^�0$�D�0 a��ĎU�<i�/,)���u�r͋�%�F�<��j�$Y��ďJ$y�f�a����<q�._0/���`Å4�ࠉ@��~�<�ル2����I�>k�<�;���o�<yƃ��NՈ �7�ПɆ����m�<AB͆M�� f�f� `�0ɓE�<G(� �Ѐ��M�\F|q��U�<�1��5��̂BFĆ �乓2WY�<�v	߲lf��bb�9�8-�e@n�<� n!ЫX8�<�a���(�|�r"O�л����h���a�b���r2"O�a�C�^����91��[�"OP�2�l�*62�`Fa�=T���V"ODaxa�N�f�iSĮ�0g4!:@"O����_�[��!��ԓZ@���"OxTõ�B5Z�ba���ت��"O8�"!��YG�Y��@�}{N�sG"OI oPx�J1 yvL� "O�t���ʻ"�zXr.�co��Iq"O���CHM;C-��kDmNW�`�"O�q�� �.8�N)YT,�_W֜x�"OVL
'D�
;��`c,)$|�d"O�E�6��>q��}�k]	]�qXs"O�	( �>P��
7+�<+*L�2"O�`���Z�<�
��lG E�b��"OTan�]��͹�Ƣq���"O�����M�K�Ĩ�$ՔE�����"O�0[��o$�=��c�%}�� �"On����4L��3D�Z9i�(.�yR��$^?֠!⤌�Z�*6*G��y� �����	�";����P��y2�ʬ��y���'0B�)�O.�y�Y>XY���M�6[\�`Qj��y"떢L��0*He�4�1q���y��Y ��艵"��-i��"у���y'�9��0��h���`�UeP��y�,״z̄Q���ْ�*�+%���y��� �t�
Fɋ��~9����y���)�Ԋa�[�x.1!�"�9�y2�hX��m��`�4�E��y��X��Cɒ���ݰD�F��yRF&s�©��.�%�`=���Ӂ�y�犍#Uޘ��B k8���X/�y�
N� �uA�MTXx�Z`
�y���DZ~��� �V]ą��bP/�y����1@4U�1���E�,�CG�y2*�-S;�����ܳ9�
2���y"I��_`4�,&�@���y2�T�
b� �ᐯ!aAQ�O�#�y�ɝ�K�ZՋq�N&"��@�iL�yBb��ղMp#���5�`���yR!U#]_�T� ��@(��P��yR��e�^$��E#�6X	VK	��y2�P�Oҹ#���S�`Y��l�%�y�bA�:�Tܢ匘>O�� U(��y�_�G�u�#X�9�V˛��y��57��v��*�pI@�&�y�5hҀ�:�X�x\��7�y2�ϥ6h��O *x\�s��ҧ�y�m�$KJ��s�X�g�б�� ���y�&O3�j��֧Q�V������y�.$�PhaDX�O�Ұs�Jm/D��ZL�R�V��U%P�m�zF�.D�p�dA�����%/͸ej��s��+D�x�Ѫرr_Pm0�e L���R�+D�@q���JC��?g,�0�<D� [��H�U��;��	�26��١�8D��s�Fڥ9�֐j�Ê)B�I��6D������E��17�o5D�x��ْ3�x�T�T�9E��X��&D�D�A
�2ASءj��T��̘Bw&8D�$����w6�����*�`�D*D��1�*H�\hz>�)O$D�� 6�x��j?�Ev��	�(ʗ"O�4� DR�K��$Q%ˁ�F���c"Oh 6X�Z�hy�	J�'B���"O�\K�(��e-q���1q9:�"O�l Ü}{��zsW.Z�C2"O�uk��5��ԁN�uJ���"O� ��b=#�U��ԍR�"O��K�Ł+X���#�K`���C"O�г�  ���v�����G"O���ȅ�Sb7�&p�"OB ��UP�3T�ۚ�����"O~���b߸�:�`��%q��0��"O�ѡ��Z��Q�V̴1PX�G"O̐y��6MX����N9128Q�"O�� ��+�Pd����7�l��"O@x�b�w��jFخb�Puٔ"O�:���0q$�h���[2➤"a"O��EV�
��c��6;,L8�p"O��%�E9Rl�8@��ŻC�}��"O���A�v������Y�d�)!G"O�٘6��_[�A��,c�"�# "O*�P�!�6���)F/Ɛ��Q��"O��"U#�0 Q��΂6�4JA"O8I��D��������k��m[�"O�� �c�7^�D���ا8FdQ2`"O���K����3�(.Hs�"O�$�0��1l|��s�%�"���"O�P�2/�~�RlC�A�:^84]�3"O��S*�?� 8q̚,�(�B"O$i��N8[\�H�C)]`0��C"Ot<�f+>6�<SӋ>\��1�"Ov�ye��.IZ�Iܖ�¥�"OTY�q�E9r���j�K�-�\��`"O�p#@nW��� Sk�ƴѰ"O��r�D��b����&d��3��8�"O.�`��W�_�&�	Rd�@����'"OZ��Ӭ �x�IBl��"O����Q�)td���	�H>���"O0��H	&%�D��/��b�H���"O�P@�ʖFl���e����w"O̐0� �1F8钀T�PL�1"O�T�4&�I
�]�D��)��̳2"Od��c�f85ïԩb�v�("OB|T�Ɔ<;�a��
�b����"O���S�M+H�t��;o�x��"OvxN͋pa�@�0��S��	�"O��9��0n^��AN2T}@�"O�8�$O8*��C�'nL!�"O�9�6��'���b�쌷 ��t�t"O�ʤ�@�,StDz����c��݁�"O^�k���~(��Jfˀ�Z v�3"O(LJ �ץM�T[$���0����g"Ov��d
~Y�(He���y?�!�a"O<T�&�����)������1"O�h"��j�@c@��*t�h`sw"O�=:*��Ym���� R��0""O�QK��	
'h�@����Ū�"O� J�� �d����M!O�9�A"OLE�7aƉ_YB�����m�.�)�"O����R�&����.iDe2�"O���"̡{�H�q��*S�@ �"OZt�ݒ}f��e��17����"O��j�摦V�8�)�f�%n��"O����P��0��7��M��"O� J9!�6u�@����B�c�$���"OFi��۴zn i�`G�%(tb(9�"OX�u���.ň}���ҵPD4�Y�"OHu����c�b��nӍ0���"Ol��Ad�Q�F8��-��n��4�"O����S���A� �&[�`�P"O|�&���6�ik��8}Θ���"O�AH��(�����EG�'ƾM�T"O��S3j��X����/BƦ�B"OH�z��ްY��
�P�MG�� "O��p�ˉ�ArN�3�B�'@�d0�"On9�3
P���Չ�A8%�"O i�p�0;',��y����s"O�0B��!5�jQ��2O�"O8 �iK�¬�W	J���3"O4�a���y� �"h�j�r�"O�1aqś�"��T�B�܋> :��R"O|��e&#�vi�t/�k�Lr�"O����g�h� !P�kZc���h2"Op�*2�= �\��c$��� "Ot� �:$�4бB�����"O�`�g�ӻE?8����#�npc�"O�u��M�c�S�Пm�ԈE"O$r�@�/d�H���!���7"O����P�H����%R����!"O�Y �-0,�&�Z�Q)��D[e"O��%�3�2��ąvK��ipU"O������d�N|�T�}m4Xa�"O���d!A�\�A	�K"DN�$�4"OPq���D���`�@0�i0"O8�(R"�b��5�
��w&p�g"O��C�lݽqq^�B⊌ (`	� "OB���*������Q�Q��0�"O>Xx����D�L�g.M�K*#"O��Y
�,0�Y���^7$��"OL}�"��R����тE�U9��Pd"O(�0�Oء}8�L�p��Q'd�RE"O���,ȜiF��ڒgN{��h��"Oс���y����o�9����u"O��>ZQ�a���UL�rS�"O�<�ծ�DR�
$�Zʐ�ht"OZ�����)mL�ȧ�;2U�$��"Op���\vpx�� N�H4`9�@"O��CӉW##$t)��K�j+����"O$J��\<\�04`!�G LIK�"O�u0��>0&�ѣ�F2�[�"O�"�"F&yq��q\�U�F"O2m���C!4��I�C\�V���a�"Ol0QcN3$~�di�%���h�I�"Ozd���̡ P~�X�D��,�Zg"O��U��/A^�=S��ʮ�|��"O�rO��[J���#�B���"O�P�����`��'��0\�a��"O(���LƨM!�X�a�Dm�@"O�	�@��f(��j'�<3� ��"OP�v(��BP�Hcv �U�pJ�"Or�+%j�^j,u٠ �4r\�M#�"O��a-Ģ!��`X��l�Y"�"O,T��nZ4�|��R��5Ym�%"O@���l	�j~�I��!\6��2"O��"�����ƈ� ��#"O2�����
L\ �Xk�2R�c'"OFa���1�fH��Ժ&�lrr"O&I�6NL)X�!,N�@�n��`"O� �*5�P��h�H��|���ȅ"Ot0����άs���C��ՙ�"O�lKsh��5��!�c�\*X ��"O�U� �[+G��-��h�5]^��"O��c�Кoy������P4"O*l03&�dy��K�:��h�E"O���8.���r@,S�"���	"O-�6�K�MS�y�Лp�"7"Oh@���A/ޡB��V�]�P���"O0y����̸�� �&M���"O
!�q��6�&���Ꮟ<!0�A!"Op݋�a�o���`�O}��iT"Od��&)n��%�	A���!�"O��r�	�Z�zY
�1դ���y�˄!aVۑ1�\�xč�+�#�y�كt`���f^`�����y��Ky��T�vJW��yЦ��y��7���N$��-x�n'^�rB�I�{m��cO]�g��}��B��sfB��>�JxKp��9��Zb�T�T�<B�	��t��o��i�5*�H�v��B�	y9$i[��#d^TU��$O�Ab�B�	&d���v��F�0�XV"��}^�B�I��]��	�)X���&�E|�B�I���� �
��yY6�d�h�"O`�t���QF8	$�d2���"O��CW.		:��sD�=x�G"O|�x��V0&Kt0�Q=*q�E"O���V.%�L48�A�x�0F"O$�h��e�ia�Oȸ��"O��5 �?X`�Y偙�a�U�"O��g� ~ލ��\�T�𠃥"O ]�1�T���Yz��%*}"O�q�aD��&�Ρ�! H=O�$�"ON��b뇠+d�Uro�<v�!�0"O���P ��]O��b7U�8�9�"OP�E �?+��!Q&D�q6�\�"ON�	�jxQGOȏE���"Oڙ(�U�^�J�[Q'M$E1\4a'"Ob-a�G�lp"����W�
�`�"O���%��68�iG&�jp�r�"Ox��$	�#J02i�%�(d��<�A"O������
mu�9¤�y&�a�"O��B ZM�����˙v�A��"O�Lȁ��:V+l���ڬZ�F"O6�V�ߙre��0�E��4���"O\)Ac$� y�<�h�	̃P�y�"O ɖ�Z-"n̺�)�a4@H�%"O�"b[&��&�:mc�!�E�!�D�)2��a�̦Z�8���ޢY�!�dD, �L�/���0%�H�!�$�.X�(���E�&��S�e��b�!�d �Q"�A*p���@���X!�$
@�(8����[��x�"�X��!�$[H��<��9i�ɚb�؎�!��?|�����%bm
7(�7�!�B�ᘔ�� %!�b�sC��<;�!�د(�:��SDQ�K����@���!��*��rE��)�-A���k!��R`�T������ �)/2T!�dܷ+���o�Mqd*�.W�!���aH�̙%(�I5��`�M A�!�DI��k�%�C�9K���6�!�dG�m@pH�i�Zx�`vK�><�!�� d�3Rg�"F:��-L�	�68��"O5C���2����&��R����"O�H'�L+2�"ԫ�唯	Fx��"O�j��J-����Ú)	*9rC"O�X)t.��uerܱ���9� %�"O*	�5�1*�Q����!WsR�"O��R�'��8ؚh���ޚ,�e��"O�t�d��xc�!*����p"O�,r�S,D�(�hѷoH"�"O������8���xC(�HnRp�Q"O(��w���}��Hړ��"Ej�Y��"O����l%a�"M���[UZ(��"O�p����N�ʩ�s ޜ8�Q�"O�A��듹Nw�`��
�в�"O��i�ʘ.9�)b�ϓ
�>t��"O�)2��3bSL���âC�T	�"O*(��-ܷtH��z�˒s�B(�"O@�� Pr�TT(fj�!-��1��"O�����Ã=Զd��(ʐF�:�R"O$ܣ�$\�[�዇�
C +�"O`K�%[�Mݪ�r�ǋ.j%V���"Od@�$@� 
PPb��<3�]ɲ"O��*�
/b�4��2���&i��"O�ECk �g)f�ٲe�&h#�"O.Ykt�� =����f(��<���"O:�K��1��bF���5��b�"O��b�I�l�y`��ۭu���F"O �c�[�y��<zw�\0�8�P�"O;@bL4fR�MH��d�"f"Ob�HP�N7bO`!f�{�h�"ONhH5��^U�ݹ�E����]x�"O�YI��Fhc'ߔ@l��3"Ony���"��:�ș8�|��2"O^�zq�;���:'ME��.��"O�ܓ�H�Uh�"l���!�2"O���7,�Ob.Xg���鹖"O��ʤ倞i$(�lZ��6i��"Ox+��ŐW8����I�4���"O(�	�l��#~܉�0
�px��zV"O6�(1�[;P*
��$ɏR�(��"O*�	�H�"�N�94��<��"O���4�U
b�C�(e�L���"O*�0W�V!"Z��O�JӨ�k'"O�E��W�)w��%�̘03fp�w"Ojxb�aE�!(dt°�_����"O<�B0K�*���{�j^�{5�[P"O@X�5���b~�Z���t"���"Ox30O�n	`�[�,�mS�"O�]Y�P$�1��/��P�3"OD�be��6<�=˄N�2���"O6�T�۹m������~ꪸ��"OT!i�W+c*|�@���&�r�S�"O��:0��"��(S��T����"OM��k��������]ݐq`"O^�!��\�(�ؖ�����AR"O���%N�r�Q�n�&V}Ju��"O���U7q��ٗ�+_JR��t"O
�ڥoS�,�vD�Dl;�ų�"O^�pd�?{\%S�G�L	�q�a"ON[v�*Q�����H�����"O����>�1��#c=��Sb�Ai�<IbBW	?�%��C\���|�P/g�<���:21ЂB=��xˣ-�`�<I�!۱ƾ,�Fc߼V2��vO�Z�<� X쪧��as~tȔ�M� 
l��"OP���U)���4fJ켩"OTP��� /Q� A%F�2��K�"O�a raәE��T9q'�:.�X�"O,ݨ��h4��b�FӢ0��re"O�-�Ǯˈ����be�5�0\��"Ol�S��%��|xT��Q�*��"O|�Q��&�������+=x\P"O{c����ǉ����Ц"O��x��*o˂��'&i�mYF"O
H3L�x<4RF^�{Q�ehq"O��t�1!�퀗dI�34���"O�H��i�R^.Y�5�3&Vh��"O^�Q�D�?��#a�y�4�'"O�����Q�\��@s��[�}�81"O�X��EE�&��E��d�0�1"Oh��f � ���C3jI�G+�u"O�ꀇ�&n��չ��'�^�� "O�42��N7k}F��ѥ'�:d��"O��E˓cYl��UJV)�X(��"O^���ֳXxn���
K`'�!�a"O��:� (Q���	�)�+���E"OZ-x���kOΐA��J,��tR2"Ox�Xa/Ε����Ɗ�#:����4"O �Q�#*�vT�j�iX��"O|���
Yw���1U�Z�fx�Y�"O*MSqM�Uxdj!L�oL:��d"O��	�ȃ�s����� ��O>�H�"O �ط,�r���:'	�($긋 "O����¹;�����v��r "O�:����t:�0!�٘!41��"Oܨy�KI�2�$�Cg"��+ X��"OT��b�C�{�� ��v�c�"O�!�̤�*�K�/By6�q"Oh�a ���j�ޠI�͢&y޸�6"O*��E���6��T�"N�`�V#�"OY�`	1� ���[y<��"O��+�f�H���C,ŗ���"O��H��݂��%�7��CҌ�� "O����yg��;�΀!T�"�ڳ"O��&dR!RR����Ć4���{"OT0g+�b`n���M�~4��"O ����KZ��ҍV,|�:	;�"O��J"��0O�L�Fk +ܢT��"O���D,��RT��~���hf"O�E���"�.����9|��q[�"OD�֌8Z����M���,�;5"ON�;�	�$;����B�4{2�:6"O^�r���1R~�AB��d�vQa"O���D�#R�u�FD"k��a�5"O��B���x(�sF�[>??2D*�"O�Җ�Ŷ<H��"gʯl�h�2"O��[�b��V59uH�0���0�"O�-H��n�,E��@���q�"Ozx�q��h�����Bf�"Q�#"O��a�ͅ.�\&�T.��4�0"ON �p.ì����M�z֞9�2"O��H����$�b�ĥy-l P "O�Ģ�)�pQk�I��f"OD�c��?Dj�:BZ֪�@"OмJ4�6D��@KSӲ%��
�"O�ԣ@�O�	�9��N¬ORn��P"O���/7
� ���7g0��Kr"O�C,ُ@�Tm�@�X�`:�;C"O� &u�kt(���FIx��C"O8�alI�:�l��5~���s�"O �Ӂ�R�x��P��a&FD�i8`"OZ��"��2Q`�bKN$z,��"O�d �J��)8@y�o͇>?�p�"O�M �n�4K`ـ��.S+4Q[�"O��;f�3>"�ū���-�Y�"O�%�D�׸����`�C.`�hX"O��X���)/Ь[���1�˰"O,$$eW�_r�DKr W�E�Ta�"O�(3&�m.V9��#
���"O� ��/^9��b�M�z�A�"Oh�@�ā;�U���
�xͺ��"O\�Y�/B���Rg�!*���"O0��'��(s�ք�#���R�"O�0:@��>��a��� P�b�"O�dR�&�2M˦�X�A
�u�X����'��Il�I�u(�J�u�bYrGP.JB�Iw^���O�t}��H�O��,(��ē�O͉O�(U`�'��t��1B�8j_��'�hp�b6���H���]�ic�'������8o!�@,�Y!�a�'�>%%A,�����@B'��"�'z&���@��[e�E�7����"}�D<��P#/��l�UÏ��|;��صJ�!򄑝5�.A�s�AO��1���4��"�S�O� @��H�\T�@	_7+H��'Ժ�sĴa��ZT+�Q�{R�'#\Q���[=U��l1C�ߠS�
=	�'fP��떥H甕ɢ.^Q5�	��'���#���H�:�i �N␥��',��
�`�=*��C�A�8.�)�'�d�t���f��i��oׁ`������F$>XhհSmD�?���aa�7�y�O���x4��l�%M�Fl��kH$�y�M��Y��pJ��J�B�\�d"z���=����[|)���:b�����޶�y�E��f��� ,�@�Q�C%�yRl�3u>�l�
�� � ��y�O��	{3�b&R����y��� ��gg̴^z����O��yҁX
rV0ȁ,S�4^�Qx�啙���0>	�d�L�`�p×�?!h�H�V�<����4�bf�ݙ��\gCQ�<ѧ+�.W�&�F-�+@Z�J!�AK�<q�	9��\)U*�	|K�D��L�D�<�6k���y��1-�P�b�e?���퓄g>(�C)�/�b�ˣ�b�C䉝.,�z0&[�fa�p1�׭5�*�O�Pڴ�M�Ó�.�b��ʼT�,zb��-K�x���(M��� #>�t��Β�j��u��r�VX��!DC,$B);F�l�ȓf�@X��_��@�����P0��X��5�J�'3t����z���Fz��~�VČb�<��Ʌb�̅K�MGj�<&��#���{�h*F \�� Ob?����<rkD����.r��L[wC��$7s,l��.V@$��G��;#�C� i'��Y�d�6
� ��'����+���V�^@�@$\.�t�'$e�C�I�s�d@� �#zĤ@�� I�B䉡%��\�����c��J�<��B��vf�=h���˾��ɠp�F"<		�I�Ʃ�W�SM�m�a�@[����S�? ��T�
%����éC�T��"O8��Ԛ<� �s��H��%C5"O���D5sӜ$��OU<^ոE��"O����o[�(?���NJ�-��\�D"O��S� E�,yaP��4>����S"O$�����Y��+5�vh2"O�=��P%l�+2��6��b"O����ҨHeD�꒤]�-���"Or�a&[��\܊d�R*!�&���"O����R�{��
S�I�t ����^H<I�����	��&L�Fp�Ѣ\d���'���Igz��cq�
[��PC��0#{!�$
k��y`R��Z�{�"�
W��hO�K�ӽ&���k��=R*th�P"O���S�ĤOR`T"����x
X�F"O�0��%���I�5`ŕe��{�"OʑP�.ٟ_y�}YG.�yG�*�+,R:�������Aͦ=q��K��Y�az��	V(*̹V��"�B'@ i�!��0gS%@��t�H��ᅋ�h�'�"=I�{�OH�~_����cK�%<�s/V��y�	аH�������{�@X�rA	eў"~�>.���'��)�4�sd��n� 0�ȓS�~��ҽ1v��{wM�u,��!�������+j�x�ch[n���w�ҫ@�ay�O̒OB��RƐL`a���ط#�($K"Oܔ ��ˌ���ٔI��.#.��U�'��I6��Ih~�I'�K�Ba��)�9��I ����Ml�B�Iͦ�qf�\�8�x̃c���;+TX��-'D�8j�Aτ#�����V�V��,$��*�;��iK�S�o�,�WOϾ$�!PR�/�>➠��ɡ�p1+�
�(8K�A�#l�������?���囑$�! �΄R�𜊵Q�<�u!��\Y�8���&�r�*�oRW�<	 �64����陧_����e�V�<9�F�E�<#4' � ��8"��V�<�ǘ$;�mP�NT�f`1���P����	�W���C'��^�H�iRŞ=� B�I�'�e w��E�O�7xR.�>��� �|9�� %JX�Nz����_�	Y��ē��!QD۲iHr$��ڔc�FEEx2�)�2Q;"�� �NK�l@�eKT��$�8�A�Y�[�J� �čZjȢ�c"�d2�S� mj1ۓK��O�`��%���m��5�� 8����y�)%5��D{��'7��Iq��0�����G_�=�ϓ�O�����/��PK�OK�?_JuB�"O�����'~[0���.G�cU���:6���ا�b �GO"uN&�)ĉ �,�G"OI���1wd�P{�ӊ�̣��${�܅�I�����eGMY��P��[��:��D*�gG|,bAAޞNB8u�gD5D�:!�'�����7<���G"Y�h��Vj��Z]Q���� @�D���oQ�h+���C��)��B�	���-��m�y�~��Э¡h�@C�	�jǰAXp� bu���W�;-[$C�ɿy��9�̓��n<��&�8L��B�ɚ]!�BA��H|����%f���~�L�� �r���Õ�=I|�(R��/|��D3���5Ć-,YT}C��W�.���#8Ov"=�d�D�w�V�bT��&\����T�<���7�>���ˬK��{��P�<!JԀg��(	�*�-m�Pst�I�<����Mur�ys w���ע�G�<� �ŊpIH������+ F4=�7"O `bŠY=X2t3�CF!/�-i2"OR)�bD�K�\��v!�>tI�"O�DYTbP3����&#b�2�"Oj�bG#V�l`�@2�
�Lc�"O:!;�Jح0Dy"eh#(aӴ"On�4(��D�ġ�M�8P�A3"O�xp��
�.J��QB�ޚ<#��%"O��g�Z�a*dQ��(V7���"O�d����@���
a&�]�F"O$%)F�P^�^�;L��Q%4�a�"O�4r/��(Aۭq�"O�+t�p+��[��5@�,��&"O~=����(���Țx�v}��"O��5�W�%�(�E�ȓQv�Q
R"O���%�3"��-�W�2��M�b"OZ�Jud�s.����݈0|�D�V"Ox��7��x4��<lR�"O��ah̼�V���1tf���%"O*M�p��g���j$YQ��S�"O �+WhG!$�$)5��4Jت#D"O,H��FL<�rt�@�c�L�"OP]��#]_G~8;�� �1�"O��J$o$~��}Z��ϭA�*�+�"O�%:s�^F�D�EG�O�~���"Ox�m�� P�@f��.|`��E"Opu���l,DC�螴e�L���"O6�*��ϗp�� ȁy��=�P"O��y�ˍ}�Rl�@_�H־�"O� ��#Z�Z�����B�:��b"O2�I��6+����Rm˷��H�"Op�1m��F�<c,��l�b)A�"Ohq��V9P�8�k��}��,�1"O�MR��"z�8H�6Jܱq��H��"O��xQ�_3�R�ȴ��;���B�"O��n��{��Ef�>5����%"Oj���HS�XQ+G΄�����"Oj�ퟘ�e�Dc�w<tЋ�"Oʝ�'�<Y��2���&x���"O2�q�Ñ|�F���Jk����"O�X�Q/дB	�(vm�.z�2�x�"O�c��V�b�r��ÊJ����v"O�Aɲ䝁���'ͦ*�>��U"O�}��
y"�!�i҅_����w"OdP����<��ȕ.Ͷ�"O���Q�$	�X��`��P�"U��"O>1a"Ӓ7� �`�9�4���"OX�x�Mày�(%�)ƫ@w�<9�"O��Y@g,Y� �0Æ۩at�K�"Oz����s�h��k �VTr�"OM���Dqj����OK��6"O �≛� j:#*	�-(����"O���OWzp|��eN	+
f��"O� �o�rx�T���+���7"O�rI	�`z>!�ĥ�l@�ap"O���d��kʂ)b�F5%jB5�"O�y	tI�=n8�g�B#|2��"O��۬r�]
�ɇP�hD��"O�����N��@�h֐6�l�e"O� *�Dt�Hš�)#�D���'A\�r'�/3��PS�G�R�8�
�'�����= �m�	(C�<��
�'����LJ/1�pӧ	�:UV��	�'���A��}�P����;c]��Y	��� �d�6��W��"��>nЌI�T"O�YS�CL�d9���C�[ J�"O`��e�>d*�	ጔ@ ��"O�H�!DP��x:�M؅U�n1�"OR�aN^�i�dXc�ށ����"Of���e�YX(��Ƴg���{p"Ob��s,J0>�����U)uz�y $"O�i$X�\����mN�`�]xd"O�!Q �;���b#�F/,T�eq"OD�Ѐ��'Lؔ���{..Y{"O�(�G�2j�`�p��W�����"OY� �I`���1+׬y��5"ODI�G�1;��ʑ� a�"}@�"O���c#]�Nj0��(&n�jd�U"O���7{"�`@I�3vL��0�"O6�K�3�JlZ�H�8E5,0R"OpQ ���3$�0�֌#�$�kB"Oz�bB[�Hj*����n�d"O|}S&�W�A�6��eP~ZT�5�'a�'9����
Ն�sVFK�Gp`��y2�'�����2�x�YhL&I90i��'iJͷV��MY��7Y!��	4j�y�LǖZ��%�u��b��A������Odt�O��a�7����΍� �Ԋ�"OZ��sÒq��Z�J *M��SwP� F{Zwp�O���DٱcH<9���H�)��T��"O�9�&�;��0�gץ]�`�i"O��؁ D�tœ3 O�O��"O\)	�ӳ%��@��o,{}�|Y@"OL�31iǻy����7��@��L��Ii>���b��w&:`C��#i0����;D��2���%����&),9��$�:D�����nm1a�͙t�����-D�����1m@ȫ�� VY��g	!D�8��Aߝ**1ٗHK.:��I�E�*D�D���R	������J�\j@�ڠ`*D��su-͔ I!��FF?\T{��&D��kg@�Rŀ��E"E-�L;$/ D���4��  �@Lx�f�6��ŀ� >D��b��ސ-G�ȇiĆ2/P�0D�hR��2�� UmT�l��U��n-D��ԇ�=u��0R���p���A1D�$P��F�s��t��Ű}��f.D�I�l�C(�����߱�1d�+D���3J��gJf��u[:=N��q�/D�ز�jD�1�&�1O��WTD)�&�+D�����2ndD��&1w>�3�I+D�(	c�P>QP��J�)T0E b0�F�'D��G��^=�2�O�YrkՅ;D�D�U���`!r1T���8pa�L4D�| ��{����񭋤wN�s�A&O(#=с�Ġ6�PM�c�[8e�p�#C�a�<QO@�
Q�i	41����+^�<y�H��QU�c�G$ \L�3Q�\�<Y(
9�
�	���e��"�TX�<��͙�Zh�h��'Q�!�`�_�'"ў� 0�Dl�=8�b\��/�̼����4�S�Wt�(A��� i����oK���������.(#_���]"`r��Q�;82��"U�+����Qf<D�'G�9UҲ��m��T�((���M+F�F�8�v���C�{^ �E[M�<iT�͖d�jM��!��b��̓EH�<!�MB0o�0���O��F�ZY�%�D�<� ^Y{��	wN��t%�
,%��K��IK�O�����b�Tw��3T�$Y�
�'�(#�lD���$A�k�=Ob�l�	�'�:M�. C�<B4��5C?���'��KژsL ���9JJU+�'�dpGӈ&�ʽ �"��-���'�Lh"&�g�0Y�f#��qδ�ʓ\.y�#H����	�'V�d^%�ȓwϊ�	�gE;
"�r�Wg:��ȓm׬�z�v��P�j������VX�'�x�I$CO�^vD��"O\�����X\X��@��jo�I�#"O���bk�?�@
�i�8X��*��4ʓ̸O�,���?p����NP�SL\��'��X\�g�l-����	�
��Oe��#&	�ىs�%�Q�e"O�0؅��<�r�!���r�4�����H���O6����P�||�w@
-^
H���'��`҂I��:�講� �k[��p�O�˓��S��O�M�2h���BP�'���=*hC�"O6��d#�H��0-�Z�Js"O��{��W�e@@UQ��8]� �T�IV�<�e���'�l�K�� �T��;2�(D���#*ז:����B�!x�`q�i"D�����]� �h޲=&ɣ6�3�O��	9E��3FLKAˎ�"0�4_NC���ĄڢMԇ8�t�#��&�4#=1��T?���Z�)��C��|Y�ܲ"C>?��8�A"D.[Q�@�
@̣a���M:�`��LǢ|:����ɘ.=���ȓt��B���
y>Ty�"�J�H�O� zV�ˢ./�]'J�-pV�D�'��f�x��( �,����U�wG:���l3�yB��?�}�$D�(�k5LP���'ߑ�D��2l�d��|E0���� U��xCA"O�9H$�5"� �PH�-&���v+1�S��yB!�NgR-�N� Lj@�E����y��ɓ3�l�2���x����u�	��y�f޵>+$��%�/m.�)$O��yb!�C�Z�{b����md M��yҏ�]��w��4G�R�IS��0=��Y$>��I�Ь�!?�TT���B��yr�ѣ&j@�Sr\�_���tꑼ�?I������x�X<f�i+ӂ�.���&��&�~C�	�g�֐��G�$��X�J�����$[a~�`S%>���b[gc��Ie��y�o�'R�J�a�$ϒp
��奋&�y�`�]��HK�eM&1I���SÈ��yrA%�L=0LC�$�z�Ȇ�y�9O�0�ԣ"_ersH1�y����@��P��RƬhh��̟�~r�'���`ԍVK��bq!T-:I.�X	�'r�E�Ǟ�!���jP�׈}���
��O���N�+���dқW�غF"O�bh�=>\�]ɳ�܅O{2�#��'�1O z4kN/JA2$�'(Ʉ6w̱I�"OTՋ��7Q��(i Ff���a"O�E!��^�dG�W��}��n�I؟���	l<EA� O<dw��c#��~��C��We���d��!�z�9�~�B�I0k��Ɠr\Q�oN�)L(b�,�� E�j9���Y�ZX) �dB�%�a��Oܴ�RI��I��iC.C/�vh=O>����5w��(G�u�4�S�蝧�!�� �Ti��:��1�KE�pz�q�"ODL3� �IO@-�R%T�=GʴB�K(�S��ybdѯ\B�ks�&�Y�MK�ybg�|���q�ڲ������5�yr�5��E��W��K��Y*r@��-j�`��K��0J�HȚy|�ȓ;�H���N��șu��l�(�ȓD��(*�a��u�(�N��M%�ćȓi>p��5c
�`91���
����]��Z����� 9�ָs�x�� ��W�@��֏L��p9����i*�K��n��h N�9J�!�ȓ�8q@V�u�&Xf�ô8�������@�9J�@�_�:��$��D5��C0C��,H�Hc��˷�
��ȓZG��Bf��C�d��l�2-edم�a�����V�s>���O,s� )�ȓ>�)æ
�,+�ԡi�A#�B�� �ʵ�"�;||���Ā*v�Є�ȓ,�T3�Y(�~hPV#Ƥv�!�ȓi��+rAޜZd�y2�]Q�丄ȓ^\�t���9�N]	�Α5�b)��;���,��u�U1f�P�؉��di�(	�I�)�ƝzBC�i�
�'7FL���D�q3��ȧl�R,��'�.��7JGmU�<sƃO�]ӈ���'�x��(ҿIZۋ�b�%]��Is�'d��P�Ud�*���<NK��
�'"P�VB$e@�Ǆ�X���'����4S��d�В!�A
�'["9����98��XEE�J��X�'�F��F7\^��À���n]��'Ub;R_H��![p@5e�&8��'V�=�Q�2*�*����X1Y�@��
�'�fMS��@�����)�� ��h��'0���E��"$\H�B}R�*�'���?C����w.w����'����#��5Yy����u*.�'�$U�#߭"$A��(������
�'&0�P%�ab�����2�8�
�'��hmVZ>ZD�Q�X� ��Z�"O�0�'c־��1zƈ�!v��aJ�"O�8� ���R9��&
�PF$1Ұ"O�RG+��̍���(n�@�"O`�&��V�F!��&�".��'"O��U`��D����0 ����"O^q0wbS�M(��{��]rԄt(���D�8[��U��)0v�"�e�!�d֧G��8@��S�!��y�S�	�!���4���QCA3\T*E"���8k!���#�ԉ��%(1���z�¬!��o�&�rF
�.���h��)-n!�JS�dY[S�A�P	���;N!�P(oV�$p�ʘ�"H8���b��w.!�$ܵ:2"�rR+S�b���!�U!�Ċ�w� $�
���t����2%!�d�k�����N��}� �Qw��a!�D�uN�頕Â�hPR��>[ !�Z�
�׎O��>0i�mE!�L�.������h�&�����#!�1>�X���7@����D�!�$�28���2+	9-<a��_/f�!�ܟc�t�R1��	!�q���� �!��#r�@�ݒ^�q���]�!�� ~��B0�ACv 4��30"O��q�A�Js ��Z1:���"O�h�aGոY��8X��ݒ�bf"O>$��	C�,YL| `L)б�Q"O|]�Y�MQ���\U�tCsˏ�?@!��c;Z<%K9
m�E��kP�uS!���+~��ϛL�2�鍌LU!�$Jo_�U[�Mώ��M��x]!�$��G%�t�%���A�+2�ӥ�!��\�{":u)Q㒓3����YZC��	KE2Ĉ���dv@�	`�!yD�C�I�D�ҝ@��Ʊa��(�6f�X�B�ɸ6h�Z�DW<!w0��#iȫ|�C�	�La��q�lS����S	8�C䉪
a�����Ewڥ�#�Ѹbm�C䉉0B����$��9˼�# J�ZN��$�q��"1�>t�-Q ʃ> 1��݃T��S7��Ҧ}��� g�6�sӓ5����)
��0ǈ�L�|�Gy���7���Ui-���H�N�t�o�<[6lp�#	\޹����F���@@On!C[�ZX����mP�����p4����%��&�	�F��bw�i��0�I|λ:�~UX6&ě"��ĉ���9� ���a�F�����_Pz4��,��剗1J���D9O��pF��r0t���B�ZẢC��fF�U+bM���Y"-��(�����E��	�r��r!R8L�D��b��/s|U9�o�u��h���M/��
�Ǒ�g�����%�֜�ÓF%9h]x*�Q(x2���FYE�>`����@L�"��	A1���p�ט`��@��Ҕb� ���bC�*��C@M�i����E�H5#U��`�B�±��-\m�d[�%�w,�@DL�̘��f	6%^��!W�C��ԭm�qᐠB.Q��SဎI2����=D�D��� �ٚ��݃W����2`�,�|I���~�8�(X�-
���8R����Gp @=:B?w�34ؽ��_;	����e�R^؞�KG��W��m��ѥw��9k��ɪ|��U����GW�H�"��ӊ��wL&hr3�E�)���(y��i�G�q�$E
?X:誁��/XƎ J��V'K�OV-���&�\�PKǕ�~-c�H�]�b1A�ΔOUԁ '��A�ղ%D�\��A���q��8佲d1#�-max��ɧr@.ٺ���� ��2i]���Xr�S.|f4����-�̙``j$uO4��G&��,��R����d׭$}w�$� %�|WZq����7z�KO���?����tg��I�?@��2m��mu����ZE�N�� �ϐ/�����G�9tg����E=M�7:�k�82�v4���B"l�aA�qFn��Ƀv$"�
��	�8iL�F�@'A�̍�#��_�ܲb��&,l2�	�8Re�����/�D�� ��G�ұ�� �X��ʒid?k��C�&Aq�Y.PA�T;ōh�/�Fi[�j.}�����`�^9��MU�p����W�A!|ԼL�p�5�FD��eـ�,���
���s	�OR�%�p+ ���OFL������sEA=un�;rĕ	&�`��i}�})��\��C�Ń�6�yJoL���}����^0�p��޹++\ܣ�g��x���2��6q����%�O�YrM
����b£��)�^�r��#۶���H�/%8�p�*O�p�gC"?���xr�K:���λ)?@��lĲ/���b�N�5n�����uܠU��-��"H��R�\�RDU6Ǻ��bD�>Q�bב&��YVE��%��\iT��S%l!�
ZeR�YI�'V\a�#o�&�d�-��ˌ�d�`���J2��AѪq��(��4SB��$�(�U�r��bEE��D4��b�� �Jq��'��Q[Z%3��.%�r������n=x�kK���fC�,v����!��}�A�i9��:GI@ 	�~ B݆@����4^�$)@��9P������w��p���C8;���S�m|�~Rb��Sv�����R����G�T�7(N�s5g�_!,�x�] z�@�j��T:Uy�ؠ�����%�h�-�y7ć�6'��œ*4����+�p<YB�N7^��D�X�&��0��E�~�|y��![�T���T�>��0�w����(�5AO�.�J���
N�y�fU��K�Y�L��
�����i���14,�3�F��I��剰!q�xe��'@�Bp�wƛ0wq1s�'4TL�h"d��}i�-c#�Ӡ,`	;��1�Z��Mě4e2�B��3|6,+a�i�H�QC��"'�<�2c��7F�2d�&6p�P�H�����mP!
�:4s��D�2������#�0$C���B����0j�L,d`�2����B�QЃ��<��`���'����['!����ѧ!l�b�×+;nS�|q��O�{����G�{�P��f%�&����\!j�|��G�E�h^�L)(�,��ͳFˈ��b(�!F�(Z�E}�,�=h��(k�)G3fn �ś�����*##" ���,,(����ʑL��Z��#��ڲiӴU�锲CLT\Zķ|�'��8���)|Y�����v�8�'M�����؝]U�!'H����U�ȫxP���u�t��n��]��˅�{�,�ʰ�I�eļl�;J�x��oV^=�f�,,O$�;c�F�Yƴꅬ���t`AB�>1"b����_��Q� �. ʧm�p1��C06D���	����I�#{NzF��]��I/�� �m��5�gm��Q�y�N. �.Q�y� I�q�A�d�H�
���1��O<�b��b8�-� zu!� $4r�Q��Q� ֽ01��//�`�$!�-2&�F$:"��l����QK�X�}`4�@3K���끯ɀ� y��`�>1f�}O��M~�'p��ܒ9�A�2k�pVVM��'��9��@ߦ/�ltQ煕%)r��\�8�I�"K'�O�R8��hgJ��=L��ȷN�78��1�#��t��	��L}�p��D�u�(�"FE JΨ��A���p �0y���O����ۨ��Y��?eT���R5����ۺç�����`�-q����I��������Qႅ%I�=��F	!9�1ɍ� Lp�̑"ll�6�"%8(�If�B�M��%j�M͓3@q�Z@!�l�j�ޜ9�Ä=�l����Ϻ����̛w9@��C�?H���^�����Ȉc#���	�`�M�e�	�
C��&�0H�0c?���Opݚг�T�@U��T���Q��h?тB+8�޸�f��?F�~�!�/c��2"��N��XkQ��r�@�
V� �((�T���J7_�|�*4O̽��ʧl,~]Q�
��<�u�\��Dĝ*H�Q�����|�©�
\�V��R�^�>�t�Y7B�@��A#�3<`�#�Q: �0Y0t�Ax�\ T��J��ib��T�"�KFn��;�b���H&gʛ�
u��ኣ���������jUx��l��@cgFg��c���p<)�i�c�ܰVm��B�X�V�T�j��-�Rd��lڨ�P�hĞf�X��&)� ,I�c>��fi>?����|��M��NWr����r<��`ئBƐiӅ�E��t�� ��Y�-cԬX�Z�0�!T
�� �`_r���/P�$���BG�>`h Br�2O4�4-�<e�h;A��W�y�FH���M�j(/-��1��3N$(���'���qr%ջ[Rd-����^+`�a�O��jpMԓ#�H��3H3A��"�
��1�
�R`蓠C�Ar0���D�@�Ҡ"O�1!5�O�&��Ē�鉕oO�I4�ِU�H����P��_F|1��HɆ�� h�GIb��l� �-`���D�,�H��Io� ��P�?��}HQ�TB �6�͊�)��(��,Qe$O��Q %I�SSmD'o�$�;S�'�<q��]o.$E+��]���q&ĵJ��0���X� �c4��)`NL��'O�i�gO�p�t���*�4.i`�O�:�U�LbF8�X� C�+t�x�����" g�^����\�Vᰁq�JW��y�,�!��fәEJ ���9'��]�B ݰf ����3��+���`�Y~B�DezXe+&�ɤi�6�Rd����xr�٬�������a�%� AʲqϚ�2��Ymlҍz�A��4;ǌ)O@ܲ�͒�
�2|��JQSr�P&�'Jq��T����L�	X�E�ӃGA�
�'�>��!�Z�9?���ġ%u�$1��Nܹ�`�5-*�'���C��G*oSF�p4D��$.|Q����TE:>a�`�؝?��񃐠�y�2d	� �	�.�a�Ȋ�k<{� �SU����i#Ia��>a�MI�R�~�S���yЀє�P{�<Q�ۯCڦ4)֢Yf�6��Q�4T��
ĭʒa+��x6O�n�����*��g/�}S��G	g�f��8\O��B٭[���(�'�%8&�xt^}A�,3%����'u��C�CC��Hx��#��7�0���}���.mn��v/)�'J$����.u �ȱ�y�-�ȓU���qփ9b ڠ�[&�$i�ȓ>�����ىVvbX��d��xC ��0��Y��@)9s6t{g́oh\�ȓ/�)"�a]��zae��SIz����|Ԓ�B�~������.�i�ȓt86����!�Z#�.�)���ȓ�X�Z�i�?��1�F
�Rͅȓj��4�'	BqC��r$J��i$t�ȓHo؉��eK�5���
2�@C�޵�ȓH1Gg��'�(U2�j�N�䐄ȓ7�u�L��ZP�C�Ǎ?�~܅�K)BhDKהNQD����,;����;�p!b�)L̓ÅA,:_q��V��ab�L��zt;�%��}��P���!�_�@h��Z�2H8Y��K����# k[�`��YT<�ȓ/��� 偙l�*	BT�[��ɇ�;+�T`��,Y�����4�R���4�tq0$"'lx�I�#�*�Y�ȓ �"\��� q"��9�G�yY�ȓ��xh�H e���5�]�5(��S�? JM��텁T��3pl�<4��p�"O��e�6N�x	�`��86;>��"Oj��g�-$����sh�,57(u �"O���PќV���h�'I�5,�U��"O\��q��!h����J���v"O�l�cD���dX5��g���+�"Ojqbb��
s�(
�ė7�� �"O����ݺ|�~�y�#�<Ә a"OP�{���nb��g�)/Q`K�"O�H3pkL,q���ラ��M��'"O�$���Y*k��	zC��SO~��E"O.��7
�q2~yR�/^��4"OAZE�-[0ps��ݱd��QR"OL�"�%�U����,$���"O�q�m�8o���៩1bF���"O��C��Kt-F�� H0f(Ł�"O����E����:l�-r�E�!��ѨD!�n�/S���D�� L�!�Bt�#BnM�GkT,�7V;k2!�$LS)|�3��	}J����+Ѻ. !��ԫ��l#Ưb'`�P�^�}!�$�=z�\��'�ғ1�}�c���!�0�f�����+��I��� �!򄖾IO��B�.�H�E��t�!� �I�zE�%+��U��p�"B�K�!�ԟ\��u1���cݺ�B�ᛷA�!�$="]�=��dԼy����#`H�n�!�dC"°H*�C�C������!�I&gg�p�C7j���c�%a!��y`�u▭C�O|��6���QP!�Ĉ�(�<9c���q��ZҠ��g[!���+���a$B����;���=~�!�Z ga����M�T9Pw���7�!��MI�����M���8��O?d�!�$��P�d5k�K�x�LG�¦>�!�d�":VD=y�J�M�^!p���v�!�dN<"n�(�˟5�zmPc�
�!�*U��=Ȅ�ȯg�x Z�(A�W�!���_ތ E������Ї���T�!�^:mS@(��@G4A�LqX��R%`�!���#��!��i��}���X�J]5:Y!��;+��ٳ��;��d�a�Ϲl9!�Ĕ�0��f��sA4��o��)!!� v#�ls4O��z t$���!�$�1��u���Ӣ}ɜ`"p��m!�u;�	��eB~@p1ȝ3�!���^�rD�U��V�z`��MҖ'�!�D��JmUB�l�4yB��L .!���v��aӇ�f��FI_�Y{!�EL�z��W��%#*����ze!�dF�H���idd�6JF7^!���y� B��T:2�	��h !򄝶^Qĩ��W"!�hA�W��*�!��H<k�F8;����(u��
o\!��A?>.:d�𩂂K��!R�ǉBY!��EO>@8�D�l�b�c���"6!��|$\��Ӎ&��ɡUE�3F!!��2J?"m���M���b`㛎!�dOqn"\�7jȘ?����O�Ub!�Ĝ�!�TpQ�FU�L���)��ն;�!���(�V�bL��r@)i�!�84��Q	C��֤�h��@&4�!�$Y�	<,����Z�X��)�8�!�_�/;� ��f����SBI�!�� �qzu�ɿ/���!�܉2�^1Y�"OؙA��WU>ä���N{� z�"O^p{$[�|*�U��U%;h����"O������	��b�Oȍm=�`�#"O�)QV�b?x%��	�h�1"O��$�>e㪑&bL�;�ꁊf"O�͠P�m�83u�D������"O�=����>u�.\V/O�B�	"O��X���&~��q��i��w$�p�"O<\+�n�/Mp�EY��,?f$�0""O�	�IU�:�����PB(1(a"O�M ��ʻ͞dÎ�pIH��"OF��7�U?P����"�*J��"O�<��ȷt�dd�& �0�s�"O�M�giA�ag�s��I�}.���a"O�L`�ܤ�l5��K����"Ol��wKG�8�*��a*�N�d�i�"O,��t䃽�lq6"��HC��ʦ"O��X��uz���u�
>�NA �"Ov]r�g �8�za�Pk�4��Tٖ�'h5��mY�J���bl�P�,
d�Y��8(��V/w�T7mڥB�H<{�!SG������5o�1�qd:&J$�(�3ʓ3C:�1��4m�!�A�:'I"�CDsӔ|�d �[����4S�F1�1��x��۹���ɃH�Q>��׋�4l踍Q��?Ό�+ S({��]��.[��M��g�P�s�5Öဍg,@m�V-��*m*Q��;D���E�G�~I��׍Ul>����%C�F��$�Wi01zr�����Q�	W%�~�`��>1O�3r~d{6�C�z%��8�cJ@؞t�o.lhA�ߺcm�$�Q��.-�<�;A��� x(@&K��d����<��H��B�0<A����ȡ@�RRH9�ǋPd�R���b�i�2F��2CF `FUaE(߭G���� E=��)�'�i�6��)��w�6]x䃎]���5��&(z�\p�{QD��O�S��X�rg��q=��Чeřc���k�/�%.q�@@W�����n����@eV�J�݌bt$�F�>T��c�� }�|9V>0^����ι3j ��,A�a3p������|s����	3 ��_�f� �k��$�A蕮B+P ��)�Z08��-lOv���� 誅1$c� �T-���\�'*U�q̚	I�Z	AT���-�6˸��ԨT'�N�ɝ2!4i���;}�oP!K	p骧��\��Y������'(\����<F�2�UK_4Sh�R�a�-}`�s䨓;	#$@��H7c�^�[�o�F�B�ːB�F��d��U�g�n�y�l$O4�Fʐ��ܤY�$�,�\ȓfk�"n�e��.�bC�ZQIĿn� Ҷ*��ƔV�A-�PЫvk��i�f@k��L�y̞l�Q���d���� �F�$)����B\��	V�P~o, xT]>.�68�e�c�
��׆��Es�ţ")��^� �y��њ{f0 �眽)�kLW�R}���OU=;�����U�=�퉃>T� @
^#B���A��K�a���j N�/�jh�A��%	�,9F+X(��(�RH��/�u  �g����� (�tT�g?�gbȷWn��c�@�N\&�h��x�	-�A���%�D����N>.$M�0 q��pퟴZ�l���Rq$�]" b�j��q�E�(y�>I@��+���7ߨO�<#�`JC8�R ��3S�Y�u��2(p�$R��K�\�\Ȏ{0 ÇLL&�:� ��U�i����쑐&c�6�6X�/�oH=�`Iߋm5�y3��2t�+5�Y���K'7��3r/��<ؤ��*�I˶xb�P�x�6�̫GS$=�r��h�೜w��՚@j�a�� ��e�n4��}�$43�#�&M�pq F�×V�vL���O�����jIb}ң
6vpl�Տ�SF-[2�(X0�Tw�%Z�vQE�Ot1�n�B̃�eHG�T(J��	
G��4���ɡE�N����
:��h�'*�0��O�<!L<��]�~��%��1/��`��"�vQ�ɓ��Z1�d����)s��BăQ�9��u�6]�1� ��Rg]�A1)�#K��h��	r�)Q*v��t�#<��Y��il4=
ӅO8H���g%/ܹ�G�.��Uؤj�����DQ�i�~%�&_�޲���'�0����L�i#�El_^����x��qCȶ���&���8����w��t�E�ֈ9X����j^�Ey�=tH�"��Cs$�:0��&2Wv��璱W�(�Nȿ �~a3��~>%���0s��C�J֥7\b��Q���T�&+�^���E��B���[D�6Gs��҂�&Q^�͠S�J��p�QGh�i��;�eݍ<[�pJ���8��Yt�A).����B6�"���C*�����J�$4y��I#Y !���A��D�!ד~~���R�|� h�𩕛eOj��!G�"[$-��oA��J�q�d{h�p��R%}|UK���7�R��2���q�H���u��<s�� _�4A��ԅ�E���#d�u�� ^a ޖ�;���^�6q���qy0k`�e�Į׵*��)ؑ�Հ>U�9[0�O����X�%�$a:g��T1�v,S�1�b������J�`a!p��o�:�:�Hֺ�M�g���/��"�M�&��Y���!)�*{�"�����4��"73�R�y�%c�Q�>a
�#�3n�)0U^?� �M���M88p�k:SN��Y��i���� ��-�~�cW�	5��<�#���8�&��*�����M3:��!�*@�iU��JQIʉ_�L=�K|J�"R���Bv'B�9*Tcb�: ��*4�%>'���
�'�raH4nZ
_ε���C�dI���׆�M[Qa��Us`8QC-�0�ҰH�t�IZ.��;�@�G�J���4R��=I����V�H�ј�N2���7�_ �*򗋑�E9�8�G�}c����>���>s��K~�'����!n؈Oj���ੁ0$��*���Ҳz<��	M?r>1$>�k�`��K����d)3]�X(��ڼ'
0��daNJ���Ex���9wٜ��A��\��(c.6LO���!��/ Wd�w�,"�x�#�b0`�X���AHv��t�}H<R�޾ �T��sJɅ{�z��')Zv�Iz�v��Wɚ�#R��3�(=���>Q�E�Z#�B����*h.��DI;D����"Q1EϾ��PL	�h� ���{% 1d��	͚��H �b��c?=�Od��&�$�<Ex3��`&���
O6�Cc�G"\w�퐰� FX�i��vPr��'�P6!��D�B9DiÓ.�<��	X�nw䀐V�T)���I�O�>i��g�7kސ"}��� L�t�ha��f<D���ib��y�B�	�aZ�T��*�*�12Ɲ�^�=V�I(�M�//&��g��(��3��E�'W�x��M�9n�h�n41٪��.N��^DZB��Aπ0��	�Xv�)9tE�(���A�X̧� �'�TaC�@�	���r��+y����'�\y{�	�c�h����ϰ9��<���܁���@�mǿO5�0�K!]��(�vT��%�۠a��:"OG%En��/;�)s�(�~54ڀ�޸,�d ��+۬d�*�Ca!թ>>-a��K��C�	�av~�a�3�bP���.�%b:�it ��0R8P{�,�=�j�{��X̧�Z<bBMA/���E#G�2����EԶUxa�m�<(V'Ɠ�X�+���9n�F��`wf(�1-�}̧cqn �'��hA��4�U���i��c�'��py�ʙ8X�U��CQ����q/�W����S%��X�"xh��K��npjÓT�+4'��R����P<$�^0��	!8<ʥ� 
�p��ab�����8DϢB�(TSp(�7(���ɳ�N�@p�B�	"�Z�X��#r2�K'�Y�i|��lD�|nC1 ��9��(G�����f�'�:=0�,�yi� g,4�݆�V̜���nY�A�B��J\)r;��
5,�;J�yCTi��s�ā�IiܧT�B�0��RC凞|��-*%#[%z\���ē�6��C��P�hHC�a�[$�����	:ܗ�M9����-ݯyP��	ÓF;�p(��l�Lq�g��?j��e��I��z����7z���������iR�u�X�I���5;}��JW,_(<q4��6,�E�D �Y;�p��Kw�	��zh��֦j�4���E�
�b?�h���2$�:�B!ߑb����y2.M
�<�"g��io�8��dU=d��ؙ�.S(q�`�ֶi������>16�;��%�u�ƶZ�*�Kg�<�G��KE�o�`8�T�W��ػ����<�����2�B��䒀tX�	�S�\�|�
؇����z2D� �qJ�AD��?��N�Q���D�F,ܹCG�\�<�$i�"$2nуS��6v�|��a�_}�4x@�$=�?=�tH�9��Q��MҔ!�D��/D�D���C�5�����jэu���a�6D����Ţq%Txb�0�jqʴ�;D����E�B!�<��C�R�$U�E�7D��i���=�`����[��sRD(D����"VKA@��2g�M�Œ!�&D����\_"Lc#��kf�%�@/'D����ݺ`G�Yq ��w��1���1D�,�� F�2@�"Vi^�*ļ��d+D���a�G͌%°O�2E%��'�&D��FΚ"�Y�!I�+��YI>D���K�|�Z�P�D'P1���֌*D�`X`�� �r�;3E^��� b+D�L�"�.xS�� L���7D�Pӂ�.e�{Fb�^���g�2D� q�kƽ*�.�Ec�$H���0D��*���6�*Ǫ�^V�*��1D���.�XLV��NT�5Ќ.D�� � �f%�:J{b���c��`�-s�"O��X'
����B��`Z��e"O�q��o�\� ��aG9lM�U[T"O<�f��P�59%�1D�̰�"O���׋���9�dKVK�-P"O� J�x�֘����`)���"O�P����K; ��=�LQ�"O��@��N�^k�r�!�Q�q�"O���5,�*��o��m���"Oj�cIO-K̐��(t�l�3�"O����	��H�Je��"OJ@U��#� ��	? �,�"O���6m�;M�UҕJ���0H	�'8�$*r�J���YF�0rvȩ�'=F��p&L*^�$=�Q�҂�I�'"��H2ዸX��X�������'����f��GJ�3AE7�j0��'�-C���xV I�cD	y����'jX+a��#�pب!B�-X���'|L0A����0���"D>�ف�'�d���� �"r�H�F��X��'� `���Ѹ�b�&8 .ma�'��\pw�˺W錙�	W�:�Q��'�����\�8���9�@]�l�n���'K �ui�6 �VpJ&H�;c����'6$Y$/B>�~M�F�f%�2�'� �#��Q������Z�:�
�'8��1$��.��Y��]�S�N�q�'� Q���Ұ�Y%~��t��'��4
V�L�>i�`�T�;k��l��'�%��+�+�����X��m��'L޴(���6}e�0��H̹U*xj�'-`���ܳ(q�����@P���'|��� *�"H�JA�	9�&-"�'���u�ʐ�r�J1�$��=�	�'�����Ξx����ǧ�?&Bp<b	�'� �{���Df���3�!Ae��'�6�y1�FN)V���s����'cF�'E���㲅��jz����'PZ�"���8s� �Ig��q�'������f.��aK!6%jY��'z"��`����q�ԫ.s�a1
�'� ��'��HfpI�
$#e��'��]P�bƗZ�~h+���A��8�'t�5���4G5~��ك9Xx�!�'6�XR��J5q^A����(F|(�'���*�E��u�F$����'�� 3$j��%K���X+�FQ��'m�X9��t+�\���H+{�ڄb�'���@ᄊ�"4���e��o��P��'��is՝Fb(��U_�J�:�'O� 0W�V"?�V��Eă����'h�ᡂ�Z!������x	:�'{n �BhC�+ �e2'H�N��'�����;K��x��6<P�� �LA� ����g N�iC�C�;����n>�v��S':�[d��I�� Q��n&j7��u��[%��=%P�O>Az��^5��TDU�O���a�>���8 �hx�T���"�"�d�?R�xA�EЩb�BM;0 Y?��K�,�L#J����)���QrOI�^�=�1�6����K�%���⅁��Pbojc&���T�� �`K�P�`]��o�<B��,HŬ�� 
� �-��<)ċ*�`M�Á�|>A���̋M�.���!��<����O�q�I�%2_:��b>�x%g���}�Rj/��Y˅�"?����8_H��+�E>�s*S�YT��d.G?\�p��`���U%�M�p ��ᕉw{�3�I���A &^D�!��'~����љBJ j�e�#j}*�'�I��!���O
7��� Z�Bb�D$,|@��72�L�􌕯$�HPHҒ|��O��|{À�>E��*�b@1�ƌ�)�7��1�Ĉ	ç;���"U�$��T�%��u'jd$����kZ-%�L����i�|����`D��a�� ��D}"�D�
4|׌(��$Q���2�S��� ��G�)�*<@�(b�$}�f��=%���?E��+G�n��D��3�
H��� �r���a+打���p֝�Y`�q��'*
,�2ĩ	Y����y҉I�Y������?N>i�&�H2�@%��l�|���_?A6C]($Z��S�'l��-s��SO�?��!����b.b��z����4.�W�S�OG��w���AD�R��a��q�2�qgM<�)�S�V���C\� ���B��ٮiY�m3�Hժo?qO���陨m1 	`��R#�v�)��˛Ҏy�ˋ���e?!ɟ` 9��:�dɑ'�Ac��ģ��]�?��i�F=�p,�x�P���Y�i>7���d36(���獽k\8�񦂙�(�!�V�&hؕp(�X�3�BJ,:!�ē�.��6��EEܡ����K0!�D��<�֡𬟔��ܓQ��!��^	A#�	13
��Ǌ�be]1G�!�$�I��$0qG� �jD9�ܨr�!�D��L�(E3$��M���0/�=u�!��m�.p*W�Z�a��u�UGI?fu!�$�!Eü��o�a�Iw%۷[^!�$J&)���3�+�9F�f���O!�$�*O�P�d�5��=x�ʱ�!�$	�zJ�٢N�<�NO>�!�d� r9��8R�|��w�Y	u�!�$�&&��Zuy�A���B	��P�ȓa���Hp��6��t ��cz���o6�3� �������B�ɇȓx���@��O6`҇+ȥh�y��j$��N�zL�EE�"�!�ȓ-�ptہ�T���"��OP�0��L�8y���&D�hC"(�!����ȓQ�VAӴ���^�T��r��'l����S挬Kp�Ů%+R0"&��2Trهȓ�RE�aj�;}��i��!�\܇ȓ��-*�$T�G[�|ɢ�1� ���H����Cmԕt��wD��:ل�e.�0"ƚV���4�<{8���ȓ�r��q`7y���9@@��ȓ;H�Tj&�R ���PcB�,9b��S��g�uu8@F�)HO8D���¢c�S�RX*Ǔ�"�d�����59'�H7a�t�0Á�a5F�ȓt{D�5F̘>��b ��-�rB����mxP"V.i�J5��"Z��B�I�R�2�X�n��4. RH/7��C䉊/������>	
�@�"d�C�	�@��أ�L��$8�$�lxC�I'Kw�QX�Ii�x�9v@��� B�	]�h�k� ]�j[T�3�m+XB�	9U��!��R�2s$A�Ҁ��P��C��3ma�I�P�b��݂=�rB��5[/@�S��N�W��#�C(R�B�3
Y���gR�!UV�ȃ$ԣ��C�I�0\�MI��ӼNQZ�#C�N�6��C�	�f`.����J�H�:���M�;s��C䉠Eנ�3wƕ.B*�#3�ѐA~C�k�ux���%(��n�~�$C䉘K�fm�'/G8�q��24��B�ɕp{&0�@��[�0�"S(�B䉤�68��ݧ"�v(�v�ԆmĘB�	�~m�岱뛝zb>��t�~bB�ɟa复�u �Q@H*�ϓ=Ne@B�)� �m����ݒc�\e\A��"OJ��@
�p����T=UH��8�"O�ՈV�Y4S)��ȱ��l`��"OmA˟=a�~�X�+PR��k"O4�`�:o{����*C8�u��"O��#DM<@N�g' s2D���"O�e��,�9r�P��0�.�1p�"Ox�ujB-d����"tV� �&"O (��M_=:���*��\%77@<e"O&x���7P�Z�A���5jx��"O��딥S���q�&n��S�"OE0��*��4RGa��*�b���"O�I�T�G8�\���(�н� "O�bb�\1��ej���s����"O �p��E��`%�򁔈	YF(#�"O�e�ڳM�n�Q�&D�b(0��"O��scJ�N��
qc��$Ȃ"O�u�M�2ᾉI6���I�����"O���Ԇ��"څ� ͝��y�B"OB-3�<��g
�0f�,y&"O��9��Ƙf`�rk֣CL�;W"Oq���T�١臫%d�CIL�<1�@�zH�s�ϻ�li;�h�E�<��� ���)*��q�:`��Z[�<�w�s���Q%h&P�@4�c�B�<�c��#LFr !2vx�ao�{�<aq�4��X������i�v�<17�LD�4!��!��X�v��k�y�<yB
�Z���#��{H^\(����<��i����y�#X�|��0�B�<�cI�5�|����+l��[�D�G�<�H
?6d����Ǧ�:f�A�<�-�!s���a��v��Lk���h�<!�i1P�,c$�'h.T���Ed��4�?IQF������_��� W-�9B#!�dWL|nqx0U8M��y),�[�!�䕌��80%E�%�zxQ���O�!�d_4"�I��̓d�h���E�!�DՒf��v)$^�|X�$I1$�!���Zm��'_0hu�p#��!��-؎AA�dҠ* �G(d�!�J3a�Hy���Z3na�Dt!�=!�D]�p�
hZ��CX��ĨaAF�9!�$G#���͉�i4�$Â�k!�dɤX����FFR�J�c*Ʒ9�	��mӎ�ʧ.ύujd�)ggٰ'�\P�ȓ��I�i�*�Ey )G-�L�ȓ@�����!]҆x����//��ȓQI��cGg�	v�U�s�ʷB<|��ȓ�мJ���*yѾܠ�A�'���>��]cW����Az��%]( x��u~�)���ɞ@n!
���4��L��X��Ti̪)\�	��g��؆�=�(y@�؈<�9���Tay�=�ȓqg,Ż�IF5s�80�"M8Y^H�ȓM6�� �%|.vx���?ڈ�ȓS��D	��J
+�++X�bPU��Lx^�s�	x@�DJҡ<T��ȓ �p
f)
5|i�c�F�rJX�ʓ5��H[M�H4�����'��C�	5M|\9�BI>}[|��6�N,}�B�I���9vI	�=j`ܚA�9S�0C�1W�|]�Ԇɘbt~Q�1울18C�	�M���DA:ŜU�G̘~TFC�)� ��*�&6>��0R@��b�"���"O�QcF �%8P�hcK��`yt-�d"OZ-��ÕD��E�q�Z(KL�7"O��e!R�^��$���[2�i�"Oj�k�ғ�rL@�â2M�հ�"O�E 6"\��Ԋ�5�-�%"O6Ԣ4�� ��ر�	..:�x�$"O*�@��S5Q,ҘZ��	�W
�|[�"O���BI�H���sV��#Z��"Od��ՀS(+¼q:``͘~�z4"O�)8�c�&Z����g
�Թ�"OB�c ��5�ND�gO;�6���"ON�9��A��y�u��^�
i�"O�	 RO9)�p����/�" i�"Oj͘��ŊcA�	���/%���
�"O��z�OL�Q�؈ %���
L 	Ҵ"O^��U��-2����&/<�;W"O���F?� LP�P0�"O΄:�A\�4�³+�9,�J�"O"��h�U_VQi��Ӑ;�0��"OTX����3~^m@p��t�]�1"O��Vb̖W�=�D�.@�r5"O|�XR�&p�Y!��r�ڥ"O�4X@cԸM)~	�b�96؈p"O��Z�c-M���C��]?n)���"O(0�W�D���E�͠G�ʸ 4"Ot9ч�&m}h)�#��J��A��"O.artk�73V�xs��R(���"O�����|�"�+�Wܑ�R"O�21���>�$h�.�X���"Old��֔V�LI��́R�Hٕ"O��i���tm1^��ؚ�"O�����'Mn̩�눰u�<�R�"O,��g�E���˔j��&��)Є"O�����=(�x����?]��)�"Oʅ��	�����֩C����&"O<�Y4j� X�]x����,eh�A "O"�� �Z�8���)҃� ��4�"O���g��;�!;3"��s��
�"O��0���i� �g���0��"ON@0S��+$�@ I�6�T]�"OF���ń��I��G_�;��qa"O|t)q�H��b�4'�T����"O�x� A�@F��ϊf�:�hd"O��� ɪ8��)a&A*E�TU�p"O��	@ꏠT:y��F�8F~���"O"�����8����f�8H�$�("O� Sd�T}3�s�`�;W���(#"O�q����b3�0�`�Ep���W"O�U�� �Poj��(*\�	 �"O��(ۘb z��&#Z#mV��"Od,[1D�s��؛�!��x({"O���$K�+��]�PJ g� �:b"O�����WJ�N)�ȃ#==d�"O��qP���/����F �#���7"O� �����:�6t�eS�I�( "O������p�,|qto� ��|�U"ODtc�02� ��Q�ǨQ�9k"O*�:�g^�L�t��n��<þ��"O*��'$�Nd|���B����0"OPh��<n~z�a�$��^�&�g"Oʑ���-I#T�r3��)�8;R"O�  qF�Sa��Y ������Ke"Ol��@FO�GͺĂ%���0�8m�"O� ^�[�,R�y#"<��:j�P1��"OJ�� C���<��@
�v�m "O�\�2�SP�~$IVI���ga�n�<�c)
V��P�F���W��n�<���@(42\�r�Z�RA�"��j�<9�míKP�A�Cߍk]A����f�<�u�ҽ>�܀��f�9�\�Q�a�_�<�1�5mk�A�B�O�S]�`�Q��X�<�Sk]�,�c�C&y�d����{�<1�W�>~ޤ�e#��Ӛ@�"L�S�<ٖ�e�92��3٠�8̉{�<1U��,]���.J�*Q��˜��!�d�2^
eФ�)���"	_q�!���4
�"R�˷x5���%�?i!��,/ ����޳k�n�E���8!��I/Y�
�)�y�t�W��+?M!��U@��!T� X�Qdb��:L!�dC�s4�@���Q��,p:��1l!�d 7v,L��R��D�vOβA�!�DI:&䂕1V�t�`��VG�5z֔��'��J�s;�)���O����O���?�y�MH(V"a2���f��R��V�N�ʖ���s�Xx�-�R+�e�O��T$��n��)+*ONAkHI�6��ī�h�'9ф����,t�f��@-��P��M�����^?a{'j�_�(!�w����l�	G%�i�!�Z��I�Cy���?�Q
8��'�2�'j���םM}���V�Գ�X���(O��$7���h��Tf/Ja�Q��^���֦e޴�䓉��'��{�>��V��s�t�؀M
;?���4
�3PX�D�O���O��;�?���?���y͢I#�J��X�`N�L�xy�ġ����3,�23�68�M�'uuԁEybӃ8�� +�	�h>��2&;@ �!S�.K������r`J��2�l�Fy"��)�M���
8|�e� �b�x�Ѫ�{���/��O��d8��T����Y5Gц�Js�ʪm�d���'��OXi�b�}�uC����Lu �>Ѵi7V6��<�F�&E�F�'r�iW<��
�6�2�I��f2]8ve�O��w��O���O Y@��a��$H����\D�15B�qv0RA�:�t��cc��v�X�����@]I��l��)�A1@�̻8H���Ϝ[��ЁJ�L0q ���&6-8rn9�	��Mӱi2��Y����$:0,��C�2�a!�O�%�� �i��D�4jY&W6es�GRw`���׸' ў���M[d��,�Ԍ0�R1Rq�q�� ��$Z͑.O��@�n��i��ܟؖOˎ�8��'@���÷d��%hQ�t����a
C�UX����!k�����E����X����Q�ā�6�(Cٸʧ�u��!	��=G���2�+�K%����#��%y����02̍���n�9�Ai����/����B
i���hv`�S).y�'`RH���/)�Kw�0�%�'>�`t��Q.�L�򃏀U��O�D"��K�Hn~Y��	@�Y�.�HTFX�.ٶ�Fy��'g�6��ɦ9'�����
-^�H�H�t46 3bJx�����џ$�ɫ���nKɟ<�I����I|��.۪E��y�aQM�=���@��lq[D'��Pz�u�am��ٟ����5?����sV�H³���1�V8��B�4n�ڰ�R�
dj�+�	\�21!��5���t��O4���Z�	KB,:��]k����֝@򬵨�4�?��K͙�?9eH>�Y�l�I�uSD'�o�B��F�K6�c��]7�hO?��A2D�gש6/:)a�%P=%� 9����MշiM�'�x�����D�	.�nZ%��┩Iq�""78�cV�1bߊ��O ���OR,�;�?A���?�t�w���M͛i�L���N2^A��K�
"p�H���N��k�lʶ�C#�l�K�K)ʓl�V,і,��6�аz�n��Jf�eEL�-d��ai(@���i��`�-j�	��3�Q�<oZ�\â��,��9"� S,?�dH��ipJO<�$�O@�`m��:b�
BE$t��E &`�к���=��7a~[��R
�~��T�Bo�ҧ%�i4n7m8�$�Oj�D�>�gg� 2  ��      �  5  �  �+  �6  ~?  �J  �T  �Z  #a  ~g  �m  t  Hz  ��  ˆ  �  S�  ��  ڟ  �  ]�  ��  �  V�  ��  P�   �  4�  w�  m�  [�  � �	 �  �  Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�� |d��"O
`�(�;���8���-0��1%"Oj4��ND^[��"3/9�0|H�"OB���H��*�ʞRy=a"O�味V�!X��!&F�:J�$���"O,��a
���C�Ą�M�"O,$3%o�-���p���+Ն�:1"O��ݢ1����`���y14]2��i�<�6��{_���c�H�`�fX�$Kn�<��A̼VI�xR[�)�Ć�pඤ�ȓA5��('nߡ4�� �)˩%� ���,��r�؊b#`T�eT09���ȓ!�b��g��}�8�F��-? �ȓ
K|m�ș�VṔ���2�%�ȓ"R�X�j�4JN�1�˘X�i����̹	_�jZ��1!g��zܶ��ȓgil,*�J�
j�Ne��i�J%b���f	�(U��:���G��$Y^م�~r�� S�%T"���k\�jx�ȓ|4�1�îJb��@ӵ�ݩn�V��/[`�"�v4�R�!ʎ<��M�ȓ`:��z�ؚh�J�Z��$HY:	��H��p�m�C1��!��B:��0��EnjZA V;9����J[
2���	��4'J�EA�IVW&��~�(aZ��ӹ�>� o�Y�|�ȓ�f�A�
Ο7�H��M�$�����mޠP����/���ANXo*�ȓTv�����{ ��-7�*h��I��sB�8�8���3����ȓNe*M�悡;������X�o��!�ȓ'lj�#F�m�+R&;�|��2)n�C��0S4���T:
b���:�0!��e֊��)��ͷV��,�ȓ0�&�8#���� ع�L�����;�P�AFd���,w�6d��r�EQ�( �gVlɦ�M,H��,DP���|�I	$G#\���ȓ"�)���E�B	yt&B�^�LɅ�4�� ��eëF�ڙ��n��R�p�ȓp`@}bŇ�=�$�AUN��P���G{�Q�\D��cշ F�s�o9L�������y"/�SU*U!�J!9i�1pj��?!J<1�O�	+��)A<u8C��#X1L��V=^ar��ȓ�:��O��S�0�ZƩ;Z�q�ȓKB��'`�	���`w*�7t�Ġ�ȓt�~���̊�TW<l���^�pV�!��B�c��L�E���J�!.N�Dxr�>!�S����0n�M�T���Z��B�ɊF��9���ĎB��$��]3�Z�=q	ÓA1�������F��iPn�)V`���>)�p��`TK�X�yP&�X]$�'u�}��R9<5;� �$�(�����)�y�If� �H��b\kwj��yR���4@C�F�?!�lH�f�?�y��K�'ζ�9V ��]Pu�r��y�`�#�D[DF�$���b��3�y���;��Tj�!�
O1��;q�+�y!�;,�RV�-r��`��y�(L+TnbP�e��u�a	���>�������ɰU���Pgh�=KPƍ&D�x(�m��M�νA��cH�S$D�� �]���J�|hE+�Y�2�"Ob<�1偓`���k4�H�,`m��"OR��%�������i7Y��3"OVq��U9p���脴g�PʵQ�Ć���+��r�eJ�z���s�F�a5�C�	/<�&}R@��{�`͐��t�C�:�zpr�O��f�x�!$l�FC�B�I"BuN�	7A.Y܌(���>DrB�	�dhn��T���_x�!:G�Ƹ@4D�G{��9O4��@A��[���'K\�, �`"O2�b��]^�{R��e�n��Z�����i���'��톶�2�"'�I�@�\D��')���W�=,� ��VFC4kݜPI�'|��J(ŒE]��fe�+�t�A�'��h�%$ $e�5
L )�>�	�'f��� �:#4p�J�|���{b�)��"Br* cfZ�@�j碚�!�ɰH�<�vJ��Il��ġ�/-␣=E��'Q�mbG�� ��q�N�~5����'��ȋglQh�`�iC"�4~�0Ĉ�'Lr�[E�U�wT�@�2�
8�����$%��\�h֩TAƀ�pc� (%�ȓ6��j� Մi�zU�
�8y>0\��߸�)t쒡Y�T���k.����6, �;�$A-R�z8�G�Ō_�%����I�u�p� @>b��5g�0�bB�`�� �d�=�8%Js��*2�C�ɸZ��0J���4X��Aɋ'V?C�	�"����6%I"��ʷf�'Ot�B�I�l�(t���ռU7F$X���8�hB�"B l�'#�\2�(s%`E#cNB�k%��A��!'���(�I
&B�ɺC�,�2pBȇR�~p�NV/�B�ɫ�
ȫG��)SdXai�&W�C�ɴF�����E�	��H�Aӥ_u�B�	���C�#}q8d�S�$Icp {��5D�L+��77�hN/9�\��>O:�O�ʓ_Ѫ��r.Å4Ey&�U-����q*0���(���(�)ә�����hO?}Y�a�#��$95�)��YQ��0D��fAG�&�����"D*k~�@u�0D���F�RP��RB���+�q)t1�O�	�}ܲL���G�-`�,�*[c��`��'fވ��@�sB�i2��-`�j�����&�'1m�P)ɿ\��l�&J��ȓKl�H��[��`1�!D8w;nX�E����Gz��N��tZ��&f�a���0�y�O�
�����nS����`�e���'(az�EАU6��`S�	;]u ]�  ����x�lۻj�p|Q@m�0<��)K� <{K�-�ē:�p�
R��,F�P�鑡��L�z,E}��O`"|����-O�<�A��b�R��֤tH<!pK�QVb���\8���aܱ\\���X��,?!��Jx�RDJ�
�H�Emգ%J����<)�GNT#�B�A�r0�|���a�<iGm��E��t �'��t�h��.J^}�|2_������|*��]�{���r�N�S�ȬYb\~��'UBx᭘�[h��#T�r)k®����鴟���8T|ܵ�e�'���SWC6D��ra��%�e)'��?=r��Ǌ3D��3SF��v��)񎉳^bX�%i6D�3׭λ�Ve�$fɭ7L�)4D���e��0�R��FꅻE�jG�<�#�h#����l�$�C
-F a���Wv�<� ��A��D.��чGġeZ*Qp��}���t�'{��B#��6���OL�H������3D�8b���[C�=HwCʉP��qJC�'��*�S�'�,Yf�	|M�B�F����'��0��E�<U5�}z��^�-�����B�� D{����%0�	k��Y�A�\�r���R�!�D��NL���h�n ��@oB+��O8��� e(*@����21|4Hb�؎T���8E�TH�0�5�aa�&1�}"��yRɎ�m�r`���X k�đ��i�2�?�"�I��O?m[f̛J-�/��b3��'�Їȓ}�<Y��B["k���#�� 	.걗'��d?|O��3$a�!<kV�:Q�1�X�Y��	t�OT��F�C :L4�eK9
��L"۴$�!�$5޴R�C
O>�(���ˢc1O���d�A�Q+���4l�	��(OW!�Εc.<ݹ��
.I���(a`!��V�o�4��#@�X}A�
�
r!��W�H<jsʓ�n{R�3㘫*]!�T/!`Hz�hD \
�;�Ǐ��{��iD�I809(�#$4�H0��#��t� �@�'
�ys�<1 ��a�^�o]R(���$-�'*�=��N�F
� 	��9v���w&�X�/i���gL9'0��ȓo?Fؚ���X+�ɰgK@,Z��]�ȓ@.4
d�����B�h��q��e�ȓo�h �o����`�F�td��yB�t۷'�;y��a�D�V��p��5���cJJ'2 ��Ĥ�:���UX�b�H̭�@<x�D�xb!��M�MЦAL'FT�v���&-�ȓJ�:(��Lŗ��LJ��EX���ȓH�H���kX�FU*��C	�!i�`ɄȓXP��A�GE�l��I�EѤE��I����t�0��(B=R���(�ȓe��<��ܱc�E��(I7`2����n݂e L(@����8
��t����D�W�ܖes.�I�I�7{��U�ȓ��&�e��I&/WA�I��v}�����%�l�d��jq�M��P7�ЈFL�[L��T�Z��P�ȓk��ZC�W�vn�1�'ˈ?�̆�\%� �M8�t�hsE�?\���W��8�� �?/w~�
�I�U
t�ȓ@ �2P��`F<E��5�l1�ȓ67�D ��K��@��BR�4d�ȓ#zHT&!�h��������B"O�L��T$'RpQ� r�.��v"O��#��e����
<v�]�T"O��ѫ�<j�� ä������"O���);|�X3K�U���#���y�ɐ�Fjm���ԆL��=����y� [_��Ł5�J�;�t�����y�I@/SF�NX�59 a`Bc��y򁙜���uO6j3v8�9D��X4��1@up��S�
�2���+D��"��7^(�#�$��4n6�xĩ7D�\�!-�z�ލS���u�%J�4D�����A�Vy�a)U� v!2M$D�Pb �̮y�.�CG`��abd���#D�d��O�~R씩���J�6�[d7D����&ڣc8�X'��t,�@��8D��)��M���PG+�^�&]�e�8D�(;���"������T?�=X4�8D�� �	;����H��5��Lx�t`A"O�aA.$t�B�(M�W8��'"O<�����V���Ûw�j4F"OD�1��9��D���G�%-��i'"O ��0*��@�j��i'��qT�'�"�'�r�'%R�'b�'(B�'�,%��ŨB�.�HvB�%K4E`�'gB�'YB�'���'�2�'�'bd�ii�"O��y�ē�<>E+��'��'�'���'�r�'2��'�LY �"G�FL�R�\�w*�dٟ'a"�'\��'�R�'�"�'M��'N��Cʞ�8�!���}�px�u�'���'U��'���'CB�'�b�'�dM�`�!�h$)� �2]t�E!�'���'�'QR�'�r�'&��'���򬑷~��賵�N�zij��'�r�'`��'�R�'���'B�'�~9�B�F.d�{�i��h)��'�2�'���'���'8��'���'����^�F~�r6*
it�9��'�2�'X��'l"�'�R�'c�'�j���,	?<�F,Z�oV�лP�'���'�2�'r�'���'\��'�d1#f���l�L�b��Jv���'9�'�2�'F��'���'|��'7��A	P�Jy����E�8�'���'@��'���'��'��'�>M;�NP�vA���tC��Tc�����'���'Lb�'kr�'��hg�F���O���c�W�@C�ŏ�=�2u�u�Jy��'��)�3?�Q�i*ʠ�e �k�qxe�
5J�i�����$�ڦe��F�i>�	٦ŀ�EA�L_����R k�� �aE��Mc�n�tSBmY~r%ӣ `�e	V@z�ɕ2i���o�(�RŰ��bTb����Qyb퓠�<�P�DE�U~���`I�t��h�ش����<�'��'֛�wT]`��r���� �۝� IS�a�O�6�p�x���'r��q%H��<q2E�%�(��F�!㔽`&�O�<��!�f`8r.ߋ�hO���OTk7B@�	�f����8Bb!X�2Oʓ���6�^>��'�$�#��E�w��!B7 ��D7���'k�'(�˓�?��4�yB^��
�11� "����}�d4AB4?�D$�n��� T��ļD���Ĭ�?)���d��!�6-_6 K�bۡJ�����D�O?��6�����sj��Eσ�-�d�	��MktNR~�'g�J��1�4�V�i#���=��X��ؔh�X��O���fӢ���	kʘi3��(� �� ڼ �E��h#b [gQ/E�D1���4��:e�Ȭ,�I#�
�i�8Ӑ�M�YB�|���9h��pw��>>���5Sc� ���O�Os�E Ƌ�a0�C�I�W�-�W�~�*�dc�T��q)���1z�:$pi��G"�(��k�X�R��f(Em�޹��a�@����4�W����*��lH�鴣ה8H~�$
Ó;��h�E�_�D/B=iCeU�K�h�ْ/��@���5�Ҟ,`%إ	D2;�ٳ�c�)A� h2/�p%��ذG��\���<]�(oϟ���џ,�Ӭ��d�y��PrS%A4i7�q���ɛ6�'o�G5z{�i>��	�?���xZ��ԖDh�B�ŗ^�Y�ꦩJ��ʥ�M#��?����#�x�O�@���Z�ʂ��4v�0 #����M�����$�O��$������I k�2Y�g%7*�B,���T5;A� Iڴ�?���?�F,�PJ����'���>_q�l�ϒ/{��}iGaܼqDH��?� P�'���'<R�'p�"�HS��YS�ܨB!Pt�%K}Ӽ��*{ڙ'���ş�'�֝*~�26,V9��T�� Y�/J��'Z��'AB�'t����L:rj����%�FMP��ē�?������d2����"�pDږfӰ]��@c�$�O����O�˓oq&E�4=���#G�i@0h���� Y&[��������ry��'���'���R�<n ]z��%��$������Iџ��	��'Jz�� �0�q�j8[�FͥC�Π�DIM%z�@Pnݟ���Yy�'uBO.��Oa���Њɵ<�H4��AK6"���4�?����D�$K�E$>����?�X�W؉��-� (nT*���3f�6m�<���?���Iq�Od�ܴDW�(3�
.ڬI���w�xoZWy��ˆ6m�w�4�'��4(?��P�A�4e�rD:��(*ç������*�$Ty�O�"��ē$�ʵ �/+s�	5�ִ.���n���6t�ݴ�?����?q��:�������;Y\�ǣ�*#��@
@�)U�^7M �r�zʓ�?9����<i�7�Z�ɔ�dh�[��^$b!(V�i���'���+-LO���O^��Y�QHripW��,.��#a��)n�h�'���'�xu1�y�'���'�4�j�a��yJ�Q�N]6DYsQ�o�<���2'��'���ß ��My�a�k^U�h��nrS��>|�6M�O�)��D�O����O��d�OI���Ӑof*\��MT, _ q4n�8�� mşP����I��i�<�����+4�GɅԪL����ݍaR\��?����?a��?���?�'�ىlb�Fh�)����1eދFC,Z�cW'�6M�O��D�OZ���O�˓�?�]�LΧk�p��R"�$J� �AA��9� ��vW����͟x�I��X�	'� ;ش�?��/%�y!f^(3����`O,i�6y�2�iNb�'�R�<�ɟY��Q�=�B��E���U.�M��,{D�����˟`�Iܟěs��M[��?����b��	��ԣ�/� ;6�$92��Q��&�'��џ�r�a>��	]y��M� ��9g��!`�
Hk�a0Pf��*��i��'��Q���l�N���O���� ���O0X�"�سo����OG>6��@�S}b�'���4�'�ɧ�4�~Jt��= $	�h�:l�P<�7]Ԧ�j��4�M��?��R�'�?����?���>9FJiyc%+D��pf��./F�6'��n��|�On�Og�Ĉ�(�چ+Z*��b���!0��6m�O`�$�OPAGNЦI��џ`�I�	�O��r@��/L1�q��?�(�l��'<̌❧���O ���O��!�O�u�!���X�gL�RŦ�I�y��Pݴ�?����?A����Z?���_52���#��H=�x�r%Z}}r�9�y��'�r�'�BQ>I�Iw�z�KH�.?��e���S�|�x'���M���?����?Y�T?M�'Tr�6:P�{Q��?Y�Ne�0CS,�����'0r�'	r�'5S>}	�M{��&(��*@�.F��H�'��⛖�'���'���'�	���{��j>@Q$�>\�4m�.�^��`��{w��ݟ��	����������I��M���?��+��|X��B�L�,~R��MA�[���'���'��I��b�l>-�O�=�5K����t��)ܘ����i���'���'Č�$v�"��Ob��T͢O�#j\@� KMb���h�HȦ��ItyB�'�64;�O���'��I���M��. u(�h�2k>0Z� H¦���x6dO��M���?9������?�e��s��4���H7:��1q(�6��	՟���ɟ��Iyy�O'�z����k����i�,nچJt�|��4�?����?����j���?��{�H�01�7h(�c�l ��d��`�i�NX���'	ɧ�����'Fxh���������)��i@��c�4�D�O(���5�"}l������T�I��֝����$`V !�"=ȵ�M�6� 6�O�XB��S���'���'��x��9l�ҷ���"tb#�{Ӫ��V�D�&�o����ןP�ɀ��	��|b����I��x�\	6	0�j�>I�"
��?�/O��d�O$�d�<�V�`݂�aa�f8�Ӧ(=F�.E��i-��'���')�����O��pD�6��y��܉<ĉ�!��Pg�$�O����OF��O����O�1�� ]�aC#X4NF�V���xX�2]�M;���?	��?!����Ou	R9��qZ���6'����-�}P��̦��	����I�|�'Zec��%�	4>��-!�fV�+��e��.�� ��%nZ柌&���	�X!���T�O>�3�X:aHI�$��'#H�ᙦ�i4��'��ɘ|8&q�K|*���"3�K5(Z�Q���$d����� �'��'�\�8�'q�)�ݙ,��b$@B#u�˂=;�� �4��d�*�:�m�����O���^~�&�����q�㌹@M�h8B��M{���?y�O��?�N>�~*#��O�`��)�z����%���=��@��MK��?Q���J��x��'��L ��$�n�zO	2�vd�G�y��Ѓ�O��O>E�	�GoP�Lŕ��{Fc��Z��۴�?���?gB�	b�'�2�'���+��X�D*ۚuT`2n�&WX�v�|�(ϮO�������O��>b���9��?t8@+d�I	Ŧ6-�O��a��G����0�	g�i���)��r�L	b�W%M�NP#vf�>����<)/O>��O����<q�������A�DYAq寑���V�x��'{|��'z&˝Bnf�;�cӆZ=���@e�(G����':�ԟ|��˟�'�F�dp>�9uE_*U�pʀ���i��֠�>���?�K>��?� �O�<���C�J��S�K�"=4�Jb��<�F�'��'⍧~rT��&I���'�2i���R�Z��B��2%iɿ,�X6�OP�Od�$�O��vg�O"�'��X��g���R�I���(#���kٴ�?a���M!\A�M%>��	�?�˘�~�Yʰ ȹ8-�y�1�ͯ���?���r��ڍ���YÉ`NfP�#\�l�8�9��ib��?e�"q@ܴ_���l�����I�ǎqqE[��|�C�7��f�'Or撕L���|������.B}[&�ƪCA���A#Y
�M�U�F�3țf�'p��'\��i9��Ozt����*�����P�|`pԀԃ��E6@r�&�"|���<�j��Tn$l����5i� =��i���'7b�©O�fO`���O��ɦA)]J��F>@�`(� �K�(7M%���K˚�$�O����O����OP(R6�C%3��a�(	��21���i�IV+0�:I<���?	M>��-���!L�8+�zl�aNa��	�'iv�;�'r�I�����[�@�Xh����H(��_3"�dH{������?�����?���&�X���;u���(Ð,;�)!�Ŭ�?��O����#�n�������p�c>e�b+v����dK�eC
���C6D�0V�İmXJ\B�C��,N:\��'4�	�'�@�s��3F-�]��&��5ٲ 2�2hÔ���@�[�k��V؄��|�r��q�F�{�.����J�)��qht���#{�dTm̴j�t�9�
�Hۢ��׀�%'�6aCP��t�&GW���gɂ;G�^$���G�Gm���"ե@��`�w��/Rt�`��a]�y���c4�'�T!p�	�~�ӆ'D�A�	��'�r�&W�,��әT���h�M?��@��K�]].���eK�_IlH#*���]�@d�1��3>��M�0m�T�8�-���˧M$苵gP��f�2�/�>&� ��O��0e�'~��柬��ʦ7��t�@jS:6���D�>D��ȡ.�' �|�t�R',���c�
AK����?�S�? ��P�f�2�r��1�ԛeM�12P�I�I�I�� �I-tҥS@����I��i���6��0\���d�A�C}h�iV��\�� Cƥ�?�&�Q����|&�d�$��^�*��S�A��8r0 ��{�L��Ǝߪ=KԵ�U���(�kњe��Χi�.��m޹8c��(���I@�����p� ǟD�'<�e��|���Q  ���D�&���s'�#e !�.("�@S7����5�b�7�����HO�tybhS�n�*�
Aq~�)���'{�^���̢V�2�'g��'�(���$���|BwȖ+��11O�v96Xzde�D�	��G �Х:Ĥͼp7�8'�+Ȣ<��A_��ċ@�d�e�ծ���$�&
�';T���h��U��/O_��<ɕ�A�{�D�R�ҽ<��c�X�i���ɦ��?A��Q�d����W���l�J��W�|'��A4�A�µ�0���}TU�F*�I�M�L>1�Oȅ����'ZRBZ�p� 32�̅*�* ��O�.k��'O����'A��'؆�:���j(BA6jx7��a��*�L۟c����.��q�mV�:E�Q��:w�W�sMLd��(_�LQt�u鍼K���F�"a��UM��)flSbA�Q�,���Oj�l�/�MK��D=@uMC�!?bٻ!ޘn�:�����?a���?����'��~5`|[�N[�~����Q�ޱx���?y�rʛ&/����+2�C�l~��`s�Ϳx@7��<q��[�BP���'��S>������KUJ��<�4ɱ��J���x����h�	?d"�跌ϛcPqjVJ�>Rt�O<�^��-�ICvvh��Ʉ
�f�'��H���>s�E�PM"1]��!�n��]���OA��A͐�	��Ij��3s�(�M�$��B�O$lZ���'��'(�v���M�>�����/�d��<���hO�ʓR�9�Љ���a(��������4��!nڧ�MI>�6A�`��qs#�ۨ?&�CI���'R�'6�p�`B����'��'�7��7�hզ�>7Zri�c���Ys��2AG�<Q���:(��I�|&���)_�J?��$+ω.|`hr)�"?��9�dk��p���(�>�O�MQnJ�!2�e2��J?�9���Ʀ�J*OFX�!��?I��?�%_�NV�
�+�� 0�IC3����x�� >3.�*# ��	HJ��E������o�'!���'��	�=K�т$*�(rD��Ca���xmh�d���H���������\w���'c�iKUOƍ@���AM�Ճ�`W5=��Y�g��-�2�[��U�Le�U�ǓdOv$箂�{��q0#�Q�V.�(2S��F�Ψ���W�N�]S�B#O�;�'�/��]�g �h��	(���n��E��l���'Sb�� &J��LYĆ��E�e�*	k!�$����Q�U"�D�t�RWm��H_1O�m�����'���k7�hӶ���OLy��ߛH�.�+V�#[�X���O��d9U�����O���|��(RT-W[b�1�
Q���˷�Z���I#N��l�T`>O���j��
WR�����i� �.X鐍\qR$�[iU�ѫ�L�����D&\>U�f5��OlA#s�'H�7�JT}�� �(�$���:�\�1��y��'�����0�"���[+5.;dd��TmC���M�0E�'r��B��U"o��c�]�?�.OrH�
��I������Ob�y��'�����ˀaSP�۶��u�3�'m2D�%\p���C'�wFESF �ަ�'���
N&:Ջ�Q�csr�!bo[�+��C� H9�жSw�ih"O
�I�Q>U*7��Q�M���� �ġB9}�W#�?�����'��'C"*5:�/D��y��-�ht�<I����<���L8.lAy�a_Ri<G	A�������K��-BBE�Q)�􅌅C��m�����͟��^	�=�	䟨�	��]0tj	�HIE��L�$�F�u���0@%\�;���(G��R!��:$�T�'�ē^�L92�պ@��u�p�[�7�2ܓ&�@��-�F�R�8Hx� ���u�'��d�
�8��	$d|�6�+V� �����W�OR�$�9x:�p�F1�n��e@�;!�$�'*�X*D���g@����1a����HO��O�ʓF�P��4e��]t�`䭉]e������&������?����?I$��b�$�O��5~I�tmH�i����UIAd�pc��^�D�:5)�%~n��'���;cͬSl&u�dI�m[��VBL�V���p�����Q��ɍ��2�e��!58Ш�
��jE������O����B`I�ф��( !S���@�TB�	44��Y'��'fcꄡ�e�SJb�xZݴ��YW��@��i���'�ؙ����	e��QsE�y��A�C�'*R߅3[��'��	��W�8ݸacˏK�T�耋�'i�ꨫb��(<�U���$:���Z� j@�U�3S�"hZ1�@⦙𱁐 ׺lh���`>�� �J�%z�ų�kǆ6��4��G��W�
��k����'������3�ܭ���G�+�2�a�'2�'��O>�*v,�V�H�cK<rP<��!-�,��4r��� ���� `ASB��͓��$A�0<��'�U>���Lğ� �P���G:"�J�ӥ��($)��8T��O�����l�&<#����SB�ö��!Ũҵ	��G�ʧ5�xT���`"��G���}�Of�i¢�1]�U[B���:�(0��A--<x�˟* ����'{2hA�Um.���>�������Iw�O �%����ѬD�V�J�K�XP��
�'���2�KF���Z�o�w� �)b�i>i��ć�.��R֤U�*�z�AEnI=�T<lZԟ�	ڟ�&#��52.|���t�Iԟ�6q��Ⱥ�>>�#��2�\���끤J?��s�i-��k�ٳ��� ض3��F�=V.S.P� 4���)s��	�u�Rٻv,�����$r�RƢ��0�y���]�lE�i"^6�Od-Ʌ��Oq��	՟8+���Kl�`�F>Tz@h<YRec�������������c~2b:�a,��	|y�GE�0�b� ��^�\���s�L�.�1���Ȓ���'x��'�`������	�|�5*!�"��ǃ�g�Z2���e}��s�-;;Y��
U�i ���$�.v��wF�O�D3 ���ةX%��<i(�Y����75d�ݸR�l�T�����i�@�2 ����$�	2g�^ yqM�-���F�ʙK̔��HR؟��� 2���a�^$2�ȥhbN7D��)�a�Z�&�7��Jt�-Ď5��0�MS���?}�Bƥ+�*�+ v讅#�*5D���꒴��@��*��:��3D����?�1� �0e젅���$D���wk��>8��p�k[�f����$D�d3�N$�0h��܏W~E�I.D�l(@+Cj��b��^�`�I;�!-D��i�J^�fE��ڀz��Tلg-D��3��b�Bg���Tjц7D�Ыߌ	��!R2�|�s��U�<I�eX�`s 8��� G�H���R�<�
�?wJ�]��G[>e84�P�<A�I�>BS�)"f�\�"
�L�U�t�<	��љNA��h�n�3PZ�Q�� r�<aF#�%#*���4㉺J�x���m�<�kA�~�T��n��Kv�iUf�<�����UUҥb�@��6Yd��I�<�M
�K�Ճ���04"fG�<�B̕aDd�K��Hh&��g�<	�隵?$��Qg�_�x����d�Z�<�����(q������N�<,�@%Q�<a��6xP�$$t6��� EN�<A1�K%��9�`�D� SGU�<qt���.x��	(�tHh�|�<�V�[
�&I����;L��(x�}�<�fK�;$�Y���_9L5<�Wm�B�<1� V�)i�����.fFr	�U�Cs�<�O6Pe�5ǃ��>!*��W�<Q����}�sD�;%�9�$y�<����8Yܪ ���X%>�H�Z�'�L�t�R���Zw!��'HMJ�[bi5yv$*�)�J�̇ē�U��S�U�H��J:|F��Bg��<��O�,�G?��`�t��Z�I����L/�|8F�	�M�FENr�}p��i��P��m����E4���B�	%�`i���YK�Z7�@�<�ӓ|�~)�&\�`�<�7��&e(�^�´"��=�(mP�R�<~(mz��c遜����#
p���G��G�>�ɴ�L6K��C�ɭb���e��`�X|)Uς7B�$�("(M�|�I�~�1�<)��[�:��P#9�йI4�5Sd*��P��6^-
U�Q�'*�*��]�9����Qkӆ M�̉�d�R����}�dӌ�s��G�6jfn^�e;��Ž>�E��"K�RA�ED ^��b��c�'9h�X`�M
Hᰉ
�c� �a�'���GՔD�!�g�����3�4?bȠ���Q$p���T
�� �8�G~�Ú��D��M�g��qg���yCT�MQ4ys����bSȖ<]V�&���'��%�`f�w��[EO>rB%���KI������x�\	ː��	l���RDf��]��Å�L9ayB���2!Ӵt��1�޹B�2'!�D��H
 ɔ(S�A�@������tF�)�"m��'r�d8'	�4<6�J�
'rH�@ℛP��0�C�69�|���2g\��p�M��^
P����Cd��ƭكBj@�2؂/�y*' U=��'��x(#EK\�<�%�4k��,��y
� ݈s�N=!��y�� 
�D%3�X��
��	v(���P�❳W�4��r V04�Xj@m� ��1��� G�`mZ3����-\OʅHP�Ƹm�٣P	��xm��	��L�D�h����J� S��T�����}�vN����k%b�L(<ae�Oq�5O�֜�K`�V���>'�%�D�'+��$�4v�x�gG��c�q:%�-��	�lY;uZa{Ҩ��s��,i�F��W����0K߄o����U@}�h���ē\ �Q��5Of���V_��<�ԎP�����U�)���*	^��t�T$���`�B(�ţ�J�PХO{�hHwޔ���;k�@<J����π�X�	ӓ`�`���@45��0��.9��Db��EQ�b!sz���`8��~?��'��`	�T;8���	�/�On�y��'4ݩ&�.�=�0�&4����Hý��O�7�&�,�p��81��ݝrV�B�E�,`��3�퀐����$�sY	��#ɽ2�V��g��tXc/>"���3+�<�e��x���g��h((����f�'��Q{�c��Hn��PdT�pS� @�}R#̴y���qC��N"��C�R���dP�����\�������Y,XB��
!�N�ˁf�j�ؙ�j�N��=���z*�P�@��i/ ��C�] �1��/��O�̠[����+�tf@bȚ4\!�$΄j�X�CU.ןkL ��0��w��M���D�29�]a�ݤA�D�q��2{�81db�q(T"V�G�7������s}B���b��.X��M3����Q���s��:L�;�%��ē5���3r[�w>��1b��!��|�>a�\
l+x�V w��3F�<������7��I���&�O�X�sF?�\�qI(���� z��=�v.N�N�u���0{[�	����.ga{RK�>l�y�m�f�Bu9��ݴL5���wɖ��hO�kL�$E�Bq�S���zC�I�a��-a~Rǆ'BJ$(("�ʆ�:(���)�H��Ņ��'b1O:)����	HbH����'yr�m�G��R�j��0F�1B��:�\�ǨOD+A���L�!f��C��T{ �'o��I�����-�1<0<8��'���N�up�$9�?O��9'*�$�(OP����/t7N!�4K�9<F�v�O~��uф"��s4"@�+(N@ R�	050�ņaN@�aM�9��q�P��~B`5+ H�A�AR%��@M.;��Q�
��_4�$] -���O�ɞ�`iH{�.����6�6A��ԛ����.o�3i�B؟Yda�,=6)���g���o�Jh�Rc� ���]�=;��zTJ��^I	�	U�s�O@���4?3�'i�+}�]P�ɝ1	J@�5�Ι1ƹ�3ɅA�@���]�4���4
.*��ŧҩ .�T	�c�+@q����*���ܚ
B 9 �V-7�xL��L6�eiM%�=�d��� ��ux"㲴��0@�I�Q�\Z�*��U�KBi6z$A+��ȷ�@�xv�ّ�xD�.m�<��C�=X��兕�A��Ђ��85��r��,~�x��7?�([X���ECb�(��"I�`G�7;|O4�х��
0v0@�b*�MJRE����.�"@��*@��p<I=O�����@	>��@Tlp9xEo��lﴽ�c�j쑞p#'Vx���1NA�7Zލ���6:��`Wm�>""�bP#G/)�9i�JL��OZ����.e�DE"��V�J�R�q֜�tS�D�yJ�]�@[�>�r��Hy��+�A.��!X?9\����"���Q�ڝ@Z�'�J1#�J�\�ܨ�%MMNd[A�p�eȡĝ*1�P\���T�U�|��D�1vfY�6�N�ܝ��%^$+Tago�5/3����S�>�>��O�H�*6^�e��@�?" �q���Q,�|����İ����8Ɛe�ŗ%9̼JЂ�Ɵ �Or�<��+���Z��DE	 �L9�I	�2A� C�Fdۈ�Dݴ`u�T&�ĺ0@`T�M��)����M
B_��)��?�ݴa���!8rq��!�n�i�|#H<� A�9O����C�:D���э�<�0�Q��!El�]�ъ$A�Y?���|�'���5V.��Ƚ1^�8�і�p]a��®����-���y"��;1|���5��"�5��@��Q"�m���I#6�D�i������!T#[�O颜��C��a��LB~x�`��DR5�S��"[.�,���(���q�+��HO���t�-?��]wYz�YP��!<=.܃�A��0p�8�)1�{��:��ץ;>)r޼C6$�����B�.:��bv�;K�̓z���77��9�)K��u�D7]EN0�M<��)K
<���:�̐�&\�X	$���<�'�^�CI�jƍ�� ��l��![j~Z��&��x� �؃�5���<y��b��7K0�<�EFI�Ml�͑S�'���fX_��ó�N<?L�XK��џ���O��Gzʟp,��Ǩ� 5*�.��@4ěF�rX�h�3�`�A����sd�@{��_#*Xu �ė�b(
�OtΓ����԰�f>��	�I$()�-�7eT6��P"У&S4�F|"�E�D����&�Jx�l�~�(ћ@�t�"�+��C�����n�0S���S*\R����Vrpt�|B+E�P���uj��1ux͐��א�~"ĕ�{4���c��^>�-���Z� \�H���> �K�Ɣ:)�P�*�Å�4���1�4�L���MX�d�N-_kd%H�K
 oz�q��Ra����i�pH�E_N4���Pe�bFX8^�)2�.J�n�BBEvX��؁�n�u3g�R8�h�0Kǃu�bE#6#��vf*ħOfĈBdV {m랟<ZK~�'˃j�fM@p	�Z��K&"F��(Ob5�!Ó:*.fLBt�X�I"�'��aZ�F���x�'@6��у!̉����?�K�3�4M)Ӏ���M����ē9�4	r7�8Riz&�2T���F� 7���+��w��(A�h]ПF{"�ʍ_\�#��1(��$'�����١q�< ���A�p@��	�4q� ��
��Ԋ��ژ�hpI�<����Y�5����&���%�զ�Rq��I�ņD5k,ԓa���� ]? ��&��C��Ȕ'������u��-�M�q�=YCZ qC.Z*|(��K7*g�p)��AH�'�B���))m�>����sԸB/Oz�:w�\��U���'2�l�2��<酆J��`x Fі�?9s�Lz�L>	�G�	T��y�l�[n��-�`���B��߱WM�ɲa�F�=P"�>%>y�� �����h�^�t=�Ѝ��_����Ϙa���qE'LO�!"��
�t��Mi .�~��hU�Bk�O��Suy�P���I�7VC�d���� i�ȴ���H(a|�V�M��E@%��a��1n�",g2�ֶ}�j�(�'cv(�v.�>)SkUI�ܴ!ax�ز7O"�K��"��YAF�)b`��@�� 8�|��즉�o9-'����
V?�tH�Y�؁�E"xj�0�N�T��@���x�@oZ��M��%Ep�b�7qP�᯻L��r���$,��m���鑼ar$� ㄏB�I���ہ�"OR(��'��4��(��E.'�=2���|a"Q��+�2`�\EnZ�fԜ��'\j�~����Z�L�����ʭ[�% ,'ShQ��>Y��'αO�OD�R��wY�p2�G>U��0�Bkaz�+�
8��
�wmAA#!	��T�-P�c�U���!lO��rDM�J��=����$��eAV��3U��$��o�����I	P�zɆ��+��A$?	�G�<x0�����l5(�g�'����.9p`maA#�o��h�O!�LX�ĩ��܃��q� �nA���G��|@�<Z� �;��?�uk�13/�Le��52�1����!7f1�j�&�]!H�;��ɠu6-�3ނ)C����ā0A0XcK�R��,s��>� �R�������xt֭�G�NO2*t��	zk�ġP/{�1��9!�H��� K��0�.�>�I<1�&���X�����'ΰ\�/?Q� ��O��h��m��
=���M^��  ����C��,QF�'�.y8���g�mK%�Ӂ-oʱ��ꂧ,Oޕa寧cu�˖r:��O�q�*�c��z�&�>"��R�K0.�@�3�؍w�b�!�Ùa����2�NᲵe�>kIL<��f��I*��ۛf%��'�tA2�$Z8�La�)�`�`��L�B�o�4�=%?%�O4š �L7;�Q�g,>�㳇�7JP�{"�C~�Xy�1s]��+��*rV))�+Y�YZ�,Sc�:3��DF��)+�#I���-�ɟR�1f��x
՛�AK$ �n� �����7�@����F/r��oZ!:׬�I��Z8<�`e�*��7�5rI"�#R��`���R�H˘���$Y���, �I�B��*2Q���<! 9O^��'+�T��dӢ�ⅵi(�
P�'��y*f�g) �F�D�ᐢC/c<���'5u�2��B�����تR�B1��OA�1OC�%�dA�舟 t�aF(+j��F�&0o.M�u"O`���&�4�J��7x�xX�4Z���'_���e�h�g��w	xi�T���G����*K�b�<C�	�?ƪu��g�d����s�["^ZB�	�v_�r��f�ƌ�f�N3yBB�	�>,�d
�#�6ޢ&��3DB�ɂ3lN}A�@^�T � 0цާ-@�B�	/t�-)]�xׁ�.ĪC䉡_)֍�Wʛ�O�HD��Q�B䉥'~p4��.��|d�!��6��B�t��13�B,�QfM X��B�	4_̄�z�C�31�˃l��/��B��'�rB��p�U� ��B�I�9����4@��Z;�)�F�U�b�B�I%u��xQ3�K5H����+��tպC���@̼oG~�#e���&�C�ɔ"p�5PqU,?���UH�6cdC�	�B�C�@_*M���c�9>C�	�l"�5	�Y�{{��1!�X9C��
�R��R&��!�&�t��.D�� ���w)C�F�`��@H���!"O�d ���O�X�jP�0^���� "O�����FJ��)���G���:D"O�	 c�14����2^�EA"O���!O�T���ɡ/S><	�0�"O�!qQI�
�0x˅]��ݻd"O~��$��P�U�5�^��t�b�"O�u����#Ϙ�����x�B�`�"O����GQ�7;n	�A�@
U�B��"O�	����l�ӯπE���q"O��؂c��z�H*� ��H6��C1"O�
eO�F��PQ ��n�k�"O�i�H�
~T�V*Ƀ	y��"O�$*C�ۨ��ٛb)�@^āK"O�p
�R�.��!�p��i{�Es�"OnH��k��@�L:is�2�"O�eAs��_cjz�m�?~C
���"O��SÆ.*����!�]�=�J]Q$"Oԙ�0iؠU���ZQ��c�!�"Oh�U�ɕ2r���W#�1��$�"Oȸ�#&��He�L�b��@H0��"O�	Z��^=aք�� &_f��"O��;CiUaFAj7 �!��lR�"O�8@��5x�ո��?�*���"O�%�Q�Un�-��ܼt�٨w"OH��:���x�gߠ"��YQg"O�i�₞$;9*�x�&_�$�b"O& �'�e�x%K�E��^!	�"O�8�%-8O�*���؇-
"��"O��1!�-f�ΈH�A\�N8��"O��H��ƨk�ӄᏏ:�jF"O��"g-��:s�D4��}��"Oְ�vI�E>~|�b啄H�f�j�"O�,Bc�86 }Bt��8����"Oh�6m^3�,{���G_����"OLP���|(b���o_��jYS�"OrU�@m�,�b�K֫�
�T�3"O:\ZD�QB���������[�"O��JT!C4JS�l�4X�9 ~ٛ1"Ot���B��;.�49���Z���V"O,	
b%�Uz��$a/;��"O�	*��R�)�y������T�'"O�A;�!3q�,[�$��E����2"O�����[�����Sc*F�J��!"O�P� |^�p��^��B"O�y�t��3��X�4�T�;����f"O���P��r�ԩ���$���R0"O��[r䚮nlpCP���\���"OQX0F��m8�@��dT	S���3"O.��#�5b0�P�嬐"Oj�E��3���2�Q��Z���"OZQ��D�u��sa�+Q*��"O�A�`���!��Ib���YN(�d"O0��qKJ�N����.F�u2���"O�E˱�M]�V�A�k�h ;�"O,����� �4m�4(��z{��r�"O& 酀�2[��P$g�&���T"Ov=���Δ5X�S���U�Ƀ"O�����ͷQ�tL{����⩒"O�豐�Օ+BF<10�^��}ز"O���q�h�t�Ùt�#K(D���c��A,,��@A,I 7m3D�pW�F4��8֮�*9A���0D��@r�D�T`l+t�]+?+�p�0c/D��  �$�L�{y�7��uQ��l.D�d
C��4:����2ў�j�',D�����O4ʩ�T�xƈt���(D���GjJX������f�|Х*4D���UA\�mX��
��DT$3D���a�W�ҪA��PUfظS�2D���DN�>���ـ��I�N�����`�����D˗/)�A��`�rY�� �hM�!��j �ʅƆ�U"�����S�-�!���'*AHqX5��(`2�i�J[(,�!�D��6�~TQ�	���9QDǠ4~!�
#K,pƊx�\!qV@ `!�:JB4Ҕ�.^6H@� Ԅ.3!�D�D�$ݚ�lþw�X`�.��!�D�r��qQrɌUd��Ϩk!�D�`].ͪR�� b��k�-!�$3h�������Ϩ��l+]�!�D�wF(څ���"���XE
A�!���7�P\a��͔B���0��&lm!��Ӗ�X�`$�����.={h!��M�Nu 1��>�\=@�LL�W�!�$J��R�X��	`�����>�!��I�	<���Hk���Xœ!�ax��		u�Rd�懚:,�S�-�rC�I����0��/|�b���Ɔ �B��H�x�J�[N��T�I"=C�}�E!ӠhrxDy�ņ51�B��$%��)�� �4]e�Y�lC�3٬B�7��rB���Q��C)BfH�B�	(�f�(��]�5d��B�ҁQ�j���%4��4@��6a�Seψ(�J��D0�$��=bE�u��*R�S��E3>%!��F+n�|��#Ú}]TR�lQm!�я��B�H/4uJ�:����ob!�҄#�qyड़9;S�yņ��!�� ��\P��'VAhZ0c��+�!�K't�"�����]Y0���CR�!�d�.n���tG��8P$��'��9Q�!�$;�Ue�r,0oX	:;R����?��E��f�K��[IN�cg��r�<��׹r�x�s���m�k���j�<a��ܻ]�T�p �D/7dTT˒�_~�<� ڣSJ��!N�fR��`#!Nb�<��'U'Jc�ѡ�ǧm�1G�Bg�<��'�m�X�Μ9��0�&��a�<Q'��#���W�C2.��ӥ��H�<�D�V��F��u���v9%�UH�<q2�$\F��p�>��Z4$TD�<	Ei�%r�S�h
^w~��O�B�<���^|v��fEDM���d�|�<I�U
i'�J'F�j�
�k� �y�<��Jԡhr��33`�$<3:�t	Vv�<1F�JTҤ�Ԋ�"SDȹ9�L�s�<�D�U���e� q�ܠ9"��j}�)�'
%�)��֧_jf��E� y5J5����\B���(l4��/R�6���}�HH KG�T4����'U&a�ȓ/m.e7"T��z1XD�U�SUĴ��d󸩊S,�� �1눁`��y�ȓQ����e�@[��� ;�0��Z�|t� n+KB���Y9C:� ��U�>|����WD�7�_�q����ȓ7jYIFJ�k����J��O��L��ZT�X�uϷd��z�T(�B�)� nA`�I�0�˵u�bL���O���dG���pa�u�\QՄO.@.!�D^(ܚ���OF�&!N2 !��L�_����`A?R�����M�'Y!�=&�b�`�JO21R��Q,�x:!�Z�d���G�X�5pR%X:a|��|�Ř�!~�B�?�޷�#�y�BB?\Q�AƉҙ����G=�y�/׹n��{G���u�
��y���t!,����ˋ[� q��J��yR�2F���A�ڏ)|�ISB�פ�y�+�|0 V�F,$육�hu�!�$P���ĴBH��%�AN�!��X$`��?=�ɂ%FJ�jq���iӲ� t܇�T�ࡂD�lX�ؚg"O��G�S�Wdb��>e(LՒ�"O6�a�ϛT��)�FlĽ�:�"O�+��2)4�CWH��<�P4j�"O�����͌�8�����Y�p"Oʼ�"P(�=��$Y!`&4<�d"O�p��/ 6x��u�قF�`�H�"O�y�AA[�)2r��D�1��Qv"O�!���
G�Bܩ�(���JE�'!qODy9�k�"{ap!+��N+TQ��Q�O����FCm2E��RW�L@��K�K�!��B������� ��8%Ñ�E�!��M"���
O6o�(E��!�d�5fX�3�Ѳmr���uBN�_f!��:�n���Oϓ`W���ُ}P!��Y���8��0/(h�E �!��L�o|&�Q���;-~�+�K�1!�D���1�D�4�ISvf��W'a~2\��9�A�X;���J@$oנ��bb�bB�I�hO>:��>@��er%�:��#=��	A�M��˙ ���#Q$gE���b�>��� =��t�e�������b�h��eC�E�U��N����Kx��G�?DF$ඏR�,n�܄�d�T�Р\�:�� @5V`��� ���ܟ��Z��N?,��ȓj�����Ў��H:�i�X���-�,16ԂFν��#A�|�4���5I�]�����CH �b�է)�XDzb�'�����Kt�IKQ,DJ!3�'w<��U㕜M�b�I��i�J�3�'��5yE��Ym,M��@�_M�UP�'��8s"I�z��AK4(��Y�����'4h��eY-u���)���M3�ay�'-��A���hP5�7F�.�-Q�'��ș��*u4U8@LQ�z���'��U�&��3{P�b��
D�`�'S��Za�VA5���H�A&���'�\d#s�
�DJ�)�vn	<)����'���-��Zh��⓪M���'�0����V�
\���>l����'I�Aڷꄒx�P�R�ާ4��#�'6f1�dp�Z��>1(�DZ�'�`q[G��<�D``�kѳ`G����'�4[roФ��`A2^��X�'�h�SH>g���	W�I��Ex�'�Dx�F���\��K'���ȉ��'OV!
/\:
��SŨK)Rt�\	�'�*���ğ+�}��Z�BЪ��'b|sU��+H��C� Q/;4:1k
��� N��DŞ8df��fK�cg���a"O��:�JŇV��� 
�QHU��"Oؤq�)��(
 ���&P�~)�IR"O>�z�� 0 /$iP��W����"Oh��ѯ��w���D��؈��"O�����˷3���+鞁9�Ԉ��"O�(i�36,J�FI��t�6��"O>�A!�F#:;�|�&�?��U0"O*s�KK���U�Mm��<r�"O�ka�"{"���QlԐ+y�L8R"O��P�I'Sp��7,�
r,U
�"Ovi��(	��UP3������""O4Q��� ���K��H�4�Ѐ"O~T:��ݟ"ۀ�
���[�:̓b"OyW�Y�q[>�ҡY�s��:�"O��:'
�}/������&U���"O�}��B֣R�rI��T�`1d"O �A���rH�!n��C�"O�m���>(,��ChVX4Ò"Oz���d��(�p�@'.�@;�"O��;DM�7M� ����,p��"O�A�1M�!�R���4�غ�"O ����Sl�q'�H~�� "Oh�h$�?@�4 Wn�>���"O�|h��4�����̊X�l̋�"O���OF9@�L�1��s����"O�4C���X����;�����"Oe��o�$Ze��j��/<���q2"ORUa�ߟ|�����r�]	'"O|QCЎ�(�I�� K&a@%�"OƄQ��H=g���7�����i�"OD�Q7���z�<I���S$���"O\ �h�XE 0;$D����"O^���#��n�ll�gCW�L���"a"O�!��@�=b7��
0i��L-���"O"��u��48\0A�z�@�"Of8k4��(�4�+s��:cy�s"OP�R�(�=(,D��GĈU���P"O���2@I��d(��EV�q���a"OVcT�5�L�{�FX/�2Y�"O,%X��rk�њ��ƅ�T��"O��[��<6|�@	5E���20�"O� J���h�а��������"OAzSœJf����ͅ`�|E"OB("��V�(@X@�9�6�k�"O(�3M�4M�D����_��ɳ�"O�����M*J-� B,�HsE"Ov�!w��1Q��҂�; ar�# "Ol�)�nG�}�P�a�+X�G�Y1g"O<��O��� �@�[�m-:с�"O*�+���5�zP��*�,�x�P"O|�),�G��Ò�P�qU��C1"O��r�c��R��x&h�WJ��[s"O�qʥ��V���*�F��]I���"O}Z3�G/p,|(��77��*U"Oh��Q͆'&���e	� ;��d"OHe�`�����Ƥ����c"OZ5�t�Gf|:��#�܎���"OԸ��ŎY��!+�늎��	�"O,$ d˄�O+���� �4�����"O> ��"[�1�̈�r�_��8hc"Oʸ�$,�:`�lx���`�@0��"O���I*'�����b׵)��X[�"OYpЬ`�h��G:T�x�e"O� ����Nʃc_
􋵩F�xD��3"Oz��q
LKb�0�hˢA��:"O���F��`�Xk�l��\<��q$"O�$K���;a�V���F�%ͪ�2�"OH#��(�Nժ%�I�̤��&"O8(�S�Mǖ��Ɓ�,f�r��7"ONhQ�/.�)2���6��hU"Opis�/�={��=Ӧ��A*`{C"O����B�9<��tJs�֙M�n��"O2���UҪ������=��(��"O�U��LA4���lH�T"O�ȺL��F���:E�p����6"OP���]�p��ٓ�*]!Q&Iqs"O\H��	U#�`��@���"Od�k@/�+���(}��=�"O4Șem
2X�{��Ow�`�`"OJ��qȄTzt���Sª�A�"O��QX�"��p�E��
�`ݚ "O��O�A����&-'W8�,�D"Op-��C#`/�e�̛'|y�Y�"O8���"�u�h��$InX�G"O�Ai���F��0��UX
m��"O���	O���5��k�fQ��i%"OL�pt	�us@k��5����"O@=zA��;���I�N�^��7"OC���:�ڡ��N�a���B"OV��� �,�C�~��` �"O�D�q��'�٦���Z�r��Q"O|qq���aS��g���:�J�g"O=�%�[	II�}ʔe�/7{\	��"O"\KQ�Š^��1�D1�z "O�t���[�	�.�)�S����"O�<��Lġ#����1s��e��"O��YD��4-�XY"E~�����"O��ؓ.�3l�^�+šۖ	��P�"O~t�v��	Q���ҭ�&N#P�aq"O t��O�!�f,2&�2�|8�"O��:��4zVƜ��E3�`h�s"O�@�0ň���,��Jo���P"OlaZd��L�2��t�F��D� "Oް����=*]a�ds���;�"OT��NF��q�S 4����"O�x��E)pj�������"O8exQ��W�,��*��J��"Oj	��3E� ̹6��Vz qV"O�Xô$3;��<r1�͗xP���"Oa���>�� �5C�,@pw"O���C�ًT�\��Bɡ~��2"Od���Z��(Äd	}��"s"O�!���U{�PZs�^�HY�	;�"OPDr�X����&�		F���6"O"X(�OZD�*�ƒA�u��"O��3V�_�nB(H��c��G�բ"OP����T��KuBD�S��!"O�5���M;G`� S(�)(X�9�"Oι[f���Ì�T��
�4�k�"OЁ ��@"J��1�B^�sު��6"O|)�N�v��G[�t-���"O�H�E�-�\�1�f��bD(�"O@h��L�dY9QēwЬ�e"OӃJۗe��E) �]98*���"O���gFW���1Q!����"Oj����*IwHɤm��!Q��y�X�^X�:�lL=7���b��y
� �y��O��~ذ��B�2{P��p6*O֍��k�tNJ����/z�Y�'�����hR/q������: J^1�'$ P�G�3	Q�<"dƭ�� ��'̄�����" �� ٓ�T���'��!��p�Rt�T���Db���'�t	���;;؄�z��X�8uj�"�'�Z���!�?�i�C��5���y�'����%*R�(j0�����(��Q�'
�p5�Q`�P�`s�����' ��q$Ϋ@TX�1$cP�r��)�')N�����+�~��+N�r ��',��˦�ܨ|4���Kӫfb�l��'9�K!�<�RU�&�a���'������ϯ`�� +��T�b�h�'��ˇ.Tt��H��KX����'�\�bE�� x^�Y��=P��uS�'d�P��aP:<�\����]�~J�Y��'w��If�Zg羨	@@H�#�Lb�'��L��L��Q�����=#)�1��'F���/�/�
*��H���'�V@�6l��r^XMس�G�����'�p ��oX�(>Ĉ
R�U�Ҁ��'�|�'�L#��e�"�[�\�~M�'�t4��M]dh=A/ȂYT�`�
�'4�=�թ]�~gb����['T���Q
�'�����H�=t�1L\�Dy� k�'���I&�C�
0�p���BEx�'t�b疼 �:��WU�P��i�'��l��J��-Ŝᙗg� �hY��'����#�<2"�;�mV���)1�'L�*v�ЇOm⁈�ä=[���ʓ�R-C�gJ�Yu~��NZ�v��!�hg��A�)U�B"�ȓ'�X�j��"��­�5T�z�ȓ}�����&^{$�y�@CS�	Wz$��,-�AD�u��C#
�`�@ԇ�9E��p�P+���pׄ�R�Z��ȓg׾�%�l�"��'�ǧ^0 ��a����Λ^g ه/��8z���ȓS D�H1g�2P��H��Z3<�X��ȓhج��D�A�j	�	�0s��ȓG�@��1=5�$бR�Ʊ$�q��;���Tc�?uS���r�)g�r؆ȓV�!����H�D��W��[u�y�ȓ����_90�7%�$Q�ʘ�ȓMZ��`�Q	z��1��6R�lu��O�@X:�	_�n� s�So�y�ȓ�%o'�:2�댘b6��P
:D�pYA'ތ)��Ap��a��c��9D�$�eKA��7��Nz&�!W#<D��"�DȖ��y���K���L$D��R�ϛw֌BQ���M�����?D��QB)D��D�B*�,<���%>D��� !��B��V��vl'D���SIȫHUnpRT��/E�)��m D�l�5 3� � ��&v���-2D�x�1�@$|�����'�<�A1�)1D�xb����2�*�E���X�f�3D���"��b�b��AͼNP	3�<D����� TF��X���0�����:D�x��냚0�^U�e,H�X��}U�8D��y�*S�YlT��� �N���k&�7D� ��()�Ɖɂ	N�-���aO7D�� x�����r�C��;ܴa)�"O���h��<�W��j�@��!"O-�a���a�IG�{� �k�"O(��%!8��q����6#��]"�"O��ĆB��85	K4�����"O�b,X�eߨ�#��] � G"OV�V-�8*-��G�я�v8;q"O",����)$t<��"� ��"O8�*���S���r��h�B�"O2x����B'�8o�$�R ���<D� �a&5���WMJ�fx�R�/D�D����
Q�BL-[Y:|�g! D�L��#ʁ=��X3 ��Q��!*D�Ę5��3O��s��=i���;D�p��q�`�;�DQ#J\����#:D��"�!aR�ţT�Z�@�h\���+D�Bać�� ��j&~�� Iq�>D�@�RKK?0�`����^����N<D�8�M,n�A
7	7d/�e@L%D�\	��[j@:L�g�G9]Ƶ��')D��aQ֒'U>l�CH�x@����'D�,p�/J?�uJh�ٴ�u�)D��`�N���������`Z��&:D�D;���-H����Q�(X�:tf-D�|*Ǘ�O ���͢
�p[�">D����*JL �Jȉ6�,i�U#1D�$���ۣUc�iD�d�f���+D����-�-EU�!Ȁk]�4Wf`3��+D��c�C�.f6 ,����t�����.D������r��X�/�rP�-XUK)D�H�(��@q<��m�F���(��&D� �g5D����Ȩ5��iw�#D���A`�;%�G�zi��C'm!D�H���_�6��lE.%�����)D��(���0a����G��9@�P�j�a4D�(��nJ�u����H�-U<���D'D����B�M�؀;D�T��<{Da&D�����d�Dlp6%?��T�.D�lx��,�y�FmM�*�$	x .D��9�?A�Lr�$�}�P�X��-D�(�p��"�;�<�a�!O�pB�	 H@4�.�]:uXA��4N.HB�I�N�Z�y��ܼc��pb�O�M�B�{�R�K��ܮ6I�q0s,ڦe��B�	Lۜ�2�Ó@%�QH�(#3�nC�I-��i�(�ν�Ȥj��B�	pwV�t)�&�YdېB�I�Fhʱ�G�,}��Q�UKUm��ѐw0����zò��0@�!�$�%�D�������+�jO!1�!�L�3\�qc��!}P�y#+��!�$�8R��z��M %�X˖�l�!�ñ2���$��?n�p�B`,�5)
!��B+�Ƀ,8'��;3Lԁ�!�$Y6��)
d�ܔ70��i���JD!�$��w���#0�[��*9��-V!�d�<��dr�&��h�0��Kb�!��L����W3qd�gI�_�!��9b�l��g�*b��1�T��2�!�$��yh� YT�+.�\�����!y!�d�&$���:+��C[�p� �X�Fa!�Ď�ٞ@��,˄>z����դ	�!�!3� ��M�0L����B"O�ݲ���^k�m��D�>}s♹C"O� �t1�
�D���+ �>Nk詣�"O�%r�H\��bȫC;�}K�"O�$�u¿v4��s��)_!�Đ�"O�hlOK�`h��٢U;Ig%��"Obi�������#c��%`8� �"O�ec@��V���p��	\�{3"O~,��� &i�t8��W���p"O<�QS�Lh���%�˟JF�x8G"O��i�ler���ĘR>@ؚq"O8�(��H���RV�4>7���1"O
1�D\)~�����E�{DZ�sV"O����ߐKZn4Y��)(Xh�"O\a@t΋�<jP���
���a �"OʥK'H�no�}[�
�$�ڹ1"OFI3F��7�<$3�ˆ77I�D�"O~���l�x��ִ9���9T"O�D�`@��q�����	R�j�#"O��AW����([�-Z�R�0qe"OލC��'MG��c!O�66X��"O�Q����WY@�h�2!L�"O4Q3�j�!@<�cBO�:b1� 3"Ol�(�#>k��1c��T�s:��q"OnezS��iZ�i�E/��^֩Q�"O�k$�'��pp�ާEqVHs"O���"@U(��Q�Iɽct2"OVU����P-�:զT�1�.D�`�����@���~�8%�?D�L�K��Ԩ���}9�M�&!D����
őW���P)�5U����E�=D��(�-B;�ѓ��W&��`1G;D�X!�oH�J*a�G�vՒ���9D�p��m�_4�S�jN�,a��-D�4 �"~�|붮�o��5��,D�(B��Ќ~����Ǹ�!U�(D��7hˑ�j�*!aù`~P�U�9D�*u���5W:��e�,g
�����2D��
�"��/�Zi)���+1�T��e>D��A�-��� Y�!@�I�x)�	"D�xA򊞳y�\;��"{T�s7�#D�h�j�/oΘyG���h{%`Q,D���I��%��=0Ud�1f%�ia*D���`�U�U���}u�y��-D��v���F��R�ĎV��|�p�*D��u�W�Q�x�(-ހl��ădB.D���6ˊ^��ea*�?Z�@	��'D�,�A�Y��@��h�|��&D� q�
(�V i�d�	׍a�I�<I&a�.w�d
�/"�Ub��H�<�׮�=1ihx ��%P�[��C�<a2��s�ӲbH�i>�1���U�<!EH�
V��#��T�2L9��FT�<ѣ�Ѫ#�����//!R�����R�<�ł
*��Ɲ�k�d��wcW�<���ȐO�)*�M5<?X �4��Y�<�&��R��h�	8��x�U&��<�s*V�l����G9�@�r��C�<�7�U�h��]`�� 5;���дaUv�<�������\��T���lIs�<�cJ>Q�:�`�!�(�(�BQm�<y�� #~���N �������l�<��!F�`�~Xc��&���0��M�<QM�>*9�i%O�Lg}���M�<����V��Ŋ�ʵ�  H�<��,ɜ�0�*�ds.x�ӣ�Z�<� ���7�E`ޤ�r.��I�ԵW"O�͢�h�����5�
o��zv"Oz���	"���j�)G?u��)"O8���E�Z�fU�U'�0����A"O6�ˢO��]}>hk�Ɲ���}"O@䉳��*��m����h�p$"O~܈��Ѳ'���e1*<B "O��p��`M�q2�T"�t1�"O�أ)V�M���G�
/0� ���"O���(�-��P��A_xFh�&"Odd
�l٩�<�"�#N�L8T"O,����=b���j7�ѿ%��k!"Oƙ"U-U.�|���^�$�z�r"O� 󳆁���%��#߷B����6"O����_:3SRP�� 6��Qؐ"O����U0AL"��@B�/p�Q;�"OXa���J;M�9:O�7uj���g"O m�&@�\��y��N^/,g�8��"OB��nӏu������@�A_b�X�"O����i�I���B�J�J�W"O��ul�?h4p��}+�9r�"O����͒y��D8'NS��H�"O�`�ӆ�>�c��^��p)v"O�C��� T���6���N\��"O.j1�H�>�Y��)2؂��e"O�Ak��
vv6EÃd�/&��[�"O��Y1,�T¡#�s̈�$"O$���� "w�C�(�|�D"Ob��C�wB*i�&"Z({�F�c"O~�c#�ۧ����R�<�x2""Ort+��Wt��{Gn��<Р��0"O"��gD�a�P����2� ��"OF�xeNH"R!RЅ�&��MQ�"O�гw@@�3��k�]:�T��"O����Q�CI�]
V��1p��u�"O(����dt���1���"OD�{�E��bL��a�()HhA�"O���$O�L��*1��SD�i��"Oج��k-g�J�i]u��Ё"Oܩ�����ˇ�r6�����H�<���z`�jd�X���+�G�<��"O�4���S�ePh�@n�<q���(s��G%��1�"Bl�<I2!�@\v��u/A�'�� 	��_f�<A��:vn�$��9�d�ū�V�<��H"<n4�`+.v��L��A�V�<12� l4|�p �#A
����m�<Q`��t�(��jZ8>�)��-f�<qB�J�Fr��N+7\p4c��W�<I��ÞHFå�܎4\R���T�<QPH9k�!"2DHu��f�z�<I�fN�|��ZЭ�q�&	��z�<�ʄ�q`��z嫇�2m��]w�<Q!� n>fa��^5Y�]��Eu�<�Ț8��rf��P����¡_n�<���4g��ղ���X:2�W��N�<�&dCtx���d���l�ޔ�Fh�B�<���*Sњ@�@˦7��Y����}�<���K�v4`��f 2\��;���y�<i��E2�
p*�%ڡ\�R�(���j�<�����Ԣx�D9l�d]3ìLp�<q��N����ēD�p�)R��`�<ya��V脥p ��K�>�9�� F�<1W�[T.�	����\���)�{�<� �}b�6B��\(�&y�h���"O�X;��ݚE~ �
�+��La ȚV"O������h?���R,,,���"O\+��ҽHO�퐆�Q�x�"O�}aR�A3z�xö�^�_�5�"O:a	�MB�^�����.8T��"O@%��p��i���\B�u�"O@qR��+P`��K��P�,�4"O�%[!�7
=z�FK��Czj��F"OL���K�$�[U��9[�@`1"O���r��04�q���{?�d"OP9:k�Q*%A���>-��S"OAh�"T ]"���ޠ&-���"O*$�����4�4�7�6+t��F"O��y�%\xZ��b+B@
�U"O�XH_UB��[�դ6��`��W�<�E��;?�"��S���:Y(Q('��|�<�r�1y ���J(��t�)d�<!@�? ZF���!��<aP4�s�`�<Ys"C:͖�ö��!kJ�&�^�<	�$u��4��d�t��ɱgePA�<b�nn�(�HA���9uA�r�<�aiב�h0(>��8�F��l�<�)X���ڄ�غA�i���	j�<���X-���@Ĵs)�0��k�a�<�r 0� c�%ޤ��,KD�<�tCƤF�X�i��	�=Wحcvlz�<�1��;�F�:�!̄o2�yk��q�<�� �� yR�� �b��k�<�r" %�2�cu�>>����o�<�2�+���Q���	�>9"g�Q�<A�G!�`�D�"5(y� +�O�<y×�d��p�!*Y�D��A%JK�<1 f_�c-��qH�Z��8�A�Q�<ѥB�}	��b�J��;	�����G�<�&�0',R�1U��	9{�	�F��D�<1�HQ�+n�X �>�\����E�<1r�V4p��	&��.j@��Pr�w�<��ۑ2B.�Id0(1x��-t�<��#�H��%A��	�&� �Dl�<Q��A [��a��&B�d�jQa	g�<9��pE�@�m:��j��_�<� ���3��e�m�d�2u�e�<y�DK'e<�7KM����"TN�F�<�a�J�L`F	���G�����̅w�<�4��Y�ع�/�1z��tLv�<��H�4�,��"�k|�
ԅ]n�<q��U�n]d8i4��t����a�<��HG��Π��ǔA;�T���Y�<	�咀ِ-�Qɟ���J��@I�<a�H��Zi�KE����rF��E�<�v��ep"�3C(�+IU�@��A�<)Wn��0�8@��M:K��p���RA�<9����7Ö7)���#�A�<YBI��^��a�g	/z��ț��|�<!6�َj(U9wi,-*��.|�<Y�h�9jRp�ش/�1F̑�R`^^�<�R�׺o�FM@��_�
���$�]�<�"�W��`��Co�K���Ů�~�<��)ԓT ��c=T���Jw�<9��N,6O^Y��g�'cPLh� w�<)�j���(#�	;5lD�s5,q�<�C��q�~��7�B�\�E��Yi�<HӧLN� �.TqB�0�(�e�<� | 6J����r�i�H��"O�p�g���i��Q?S�Њ%"Or���C�Q���'G߁
��`w"O��P,я-�4�9vf�+~��Y�"O��0�g�u��(��_4i�b"O�,�@��.�6%���e��Pz�"O`�9tk��5K,m���՚J�Z%#�"O�L� Ñ�6JD=[U��%�H�{v"Ox���n�_�PU8a�έL����"O����kE�ZUL)�"�J� ��:"OP��W	���Q0aIO��@*`"Obܡ"oF-�nYbba�)F�M��"O���,U�c���U�O�(�n�c6"O��A#;=��ي�$
Z��ۥ"O��˵�&��d�$��o�
T�e"OtIA��Q�+��4�Eŷ�-q3"O6���4t�������ؐ�"O�I��2I��[����� �0�"O@	����+fU��S'O����"OU8%%[>��T�`$Z�~uh]s@"O`T��ʀ��L�e�Hk�,�ڵ"O:A�d֍/C:����B�$o�٫R"O
J��yb-���
�#�>D��"O��!�� ^_�Ђw�H;~�S"O��+Z�c+LT EK�v,�b�"OThj%��M��Iq�����Ԩ�"O��ag�>[�B�rSG¨h� ]�e"OND �����(-�Y휴P�"O���C鄓��x��Z}?\yZr"O����W)���g�ʧ If��F"O�-�A'��6�jh&c�
2���R"O�`�%mv�p�Y7�|�&̘w�!��;`��[�A�K��Qq�h��q�!�DԶ3Yl
C联(�z8#A�?b!���61�t�9 ��/S��%!���<T!��ԡjR���R�<�%���S6H!�7q�4������#!@Fs!�d�oۜMi��-6qd �K�w�!��="����F�v;&��%�6�!���[�xa�RO��g;�Y�3�!�DW�gh�TIp�ꬹ5��~�!�DY�R<6*�`��x���(~C�ɭyBt=��k�6e֊MY�G��k��B�I�d$ ؃&mΣ<�f�� �8<d|C�� [Y�}
 ��4rN]�f�ݘ`{jC�	�,�P���+��Dh�˝�*jBC�	G �6.Ͽy��t���0mWJC�I,��p
��6wդ8�"a���B�I��H�"�/�lZ�2%���gwlC�Iw���׎�j��A�b�$%&B��|E.��(Ɇ&�����B�;�B�ɱ?�P�2�Ɇ@��̫�,�\��C�	�vsP�{ԏ��5u޹�k�-2��C䉫.�.�����(v�yh��(<�C�(<5$�2j@�9:�*�	�C��
@�T��M�P���p�f [��C䉸'G�!;Fɕ�n%����8#�ZC�ɜK6<<xE���U��9 � C�-:�6���p5j���(�>r,C䉶ea�-y��U�ܒ��@���E�B�I�2�h�����{5X�"$��W�rB�Ie~��gM�("�6�1'�	SC�B�	�/dJ�� ͓�2}Ty�`AԪ9zB�<8f�5�KM�0��^�q�B�)� Q��g8B��y )��>E��{"O���j҅P�������<��cU"O��<�x	�E��imp<hg"OT!SA��&HYq&��� ����"Oడ�h�"9���0�ן��[p"OD�����9sZ0����b�L�"O��aZ/����4dH9Ȫ�s�"O�HC�/�)�e�X(6�� �"ObhIdɑ�#�@�QS�P�c�L��w"O��B(���
#���t����T"O�5�&FF�]$�!Q!ޕY}D�"O28@����M���S gW�%BH{t"O��[W�</��10��� @5� "O.�!�%߂����"��,�S&"O�h�R��`��bV�J2\��H� "O����B�i
Ri`Pn[>:���c�"O��IcbU�j�y9��͵~�(�#�"Ozܸ������A� �ϥ��y�R"OHiҡ�� ]��������v�kb"O�L�D��[(��b��Q����g"Od�( )�-y7��>�Rq��"O�PK�(A'$�F	�xH��"O<��A=v����	��y���>D�[ C�p�>��!�h�Ԩ�ca;D�P���=-�ę�a$�6x��81$8D��1�W�X���i���^�V	3��4D�������(�f\!%����6L2D�P0����P���4���}^X���1D���7�G5{��V�#������-D��e��m�����hM�V-D�D�R�T�Hf֘���·XVL�(v'-D��5��=k�R��n?�Z���)D�`�@�՘��P/�>~	�萔n$D�l�"o�5&V:��	rd\Ё!$D��q��Q�Gx�`!݊RlMS2�/D�$���Xa� :'C��@1��.D�X��c+� )0v�ֶrQ���� 9D� +�����M�W��_y�{�F2D�X2� ��P��Ԫ�T*��K�k=D��@@�m�B����#��qg�5D�dP�j�>x��en�/��3�G5D���G���L�Q�&ʔ[�hm��`4D�I�N
�6��I���G���k �3D�p��-J�m]�5yw(|�z�'c2D��J�H�y��Mp�'�C�\��$D��q�g0\K���!m_/�<]�3�&D�(�� [�lS���1��*�}(g�%D�0�����G�&˴I�#vx�5B,7D�|���cZ�p�V�^�Z@A2j/D��Qg$��a��H�2���;�,\�`c.D�  �ɞ�XX�9Yv(ֿ^���%e.D���c��k�`0)���
{0��r�� D�xB��	�t�fi�L֓1
�`�+D��{B�Z����S�"q#P �7D��h��ߑ}�1�������òB7D���AJ� *�:%i�c'G*Ɓs"�4D�`1pB�0p�Ҕ@��i���'D�,QP*G�?�^ypg�?*�%���&D�,��H�=��<���/7����v+%D�\� �|W4\K�ÅPx�y��)"D��	Ə�x-XJ�d���NT�!�-D���%�>ny��ڧʜ�`�V���i.D�$S��ޱL<sg�=+˒!�e�/D�x����\��X7ᙆi�K�)D�� ��!��T;}�V�����j2�4@q"Oz)9r��t�P��	����"O�T�ؤ�2�Z�MǱ'Fd��"O�eQ�gɥu� 3��M�d&��"O�t8��M��:��Vϕn,a9�"O`��d���ue�0��W&L�y�"O�A�&g_�Ic��Z?A0���"O��x�(��p�����A��[`��"O����>�ZP�]�"��#�"O�u��C�2"$Gm��y�T9��"O<��������BRp�H3�	u�<�ed4�0���	���?mh!�DR?CƼ�#O>���7j5!��܈	����/�e�R�Z)!��Q? 	�P�q�{��lb��u�!�d��,��x�TK�.��!a��0n�!��D!F�2T#A��I� �V�	w!��/>z�����1€��'ä2�!�T�y~8pC�(_��虐�v�!�$D�k��J�iY��e�U��!���[ �ق�ȅ�@dFʚ@�!��F�VpCcP�Y& ��"&_
Vi!�^�N�Υ���C���0%�&S!��w,BU[��0|����c<z?!�$Ƅ=�nT৯�b�
�@i�]Z!�$W?UR�1QB�Y>9�2]�b�H1H!�ęzX<����j?2���&=W	!�ě�$���̄BTB\y���R�!�^QMEM
�;Ҍ��\.�!��pY^ub�HB){:Ή��	�0�!�dK!����j�4n1R��+@8�!��Q.�~K�\(|�ðg�u@!��\sy�S�tC��J��c'!��9O%0 B�/�C�%:���$�!򄊸&d�`�Җ.��С�� $�!�DS71��pa@�D�/�vY�f �`�!�DB1Y��i��ֺ=�L��O��!�DR�x81I��ّ$=��cb�\;�!���l(�8G�3GԔmsoG�
�!���.��h�c/�)h�PXh���Q�!򄘲d�	�Q��8fBP+C�@4l�!�dC�x��( F�2O�{�Ɉ� =!�$�q��9DE��~�8#�ƕ!�dL�M���7�^�P�bT˥�}8!�DB�
iʭ��@1=����"��|!�d�$x!���i�]j, 87*��-,!��ǘ#�Ј��k��G����	��!��!XDĘ��P*Q�ma"�^�!�
R'(tK��Y!GI>��b�	�&�!��NS4��Sh�d�xZ��T5NF!��\<�i�!ӳa +��V�W/!��G4���r��/#��,S��¨@!�.E� p4��;x�0�xa+�>	!��wA�gdA369�8�֪e!�d�?c���Q#�_�t2��
։E�!�đw��-Z`��.,-���˞9�!�$��:=��v#M1�	�i�,#!�.��ys��9S�9�V�H>_!��Dw���5h�1@����!�%o�x4���v�lH�R�o�!�CA�J�`�R$܊��
�7!��D�(�dX?Sp��{�`�O1!�$�-Q�,Q1t$=6S��`
��!�dѐ4^� �
J��%��.g�d!	��� R�Zr�K��J1���W����"O(��L_&� �5	��ĉ�"O�5ac��)̞Y��g�?}��z�"O�eh����1��Q � z	��"Oj�Zp�EW�.$
��X�&��!�>D�$��gO����X��:���U�1D�PY�l��ks`H�� X(8��壖h2D����	�:j��a�� )Z`���k1D����?�~Y��iB�G��uE-D��҈ɣ?��kPꞄ=U�:�B?D�@[�ǆ�KĢl�B�&@���>D�`�S+��%��ū��V�M���;D��+aG�%��T��	t��Tk�5D�D�L��'-�{4CZ,Z�A��2D����g�7j>�Z�J�u<L@��0D���)F:¨� F���K�&��E�1D����m	�-0�e�Q��5h(�I�:D����cV�n[�	AE�(�H�h��6D�H��i��Oh�7�߶q�&��ơ�h�<y��B��^�B" ��E�x�3Kc�<a��^�,��I���Z`�ʒ��D�<Q��V 	Gd��m؊So2����K�<a���A��i1��P~]���O S�<	F�C��{�
D�`
̰��j�P�<9 &�% j\b�b#��lI��T�<QV�_)bT�0�#��*��m��g�<��P|<�z$�¹SXEp��
^�<��/	�JY��Iu�4���A~�<Fɓ5o(�<&	���%e^d�<��ď?Z��TX���
���H��E�<I�U�6U�4�Q�3�^���D�<I`N��}.�ӢH�7P�M0p
DB�<��T/]R �6���jvh�cMz�<�dK��_�,]!�.t�dEs���^�<YЃ\�L,�#'09{�P*�Af�<a��	���i�VaI�!X�X�b�d�<��%�3�Y*�#ϧBCzEh��Z�<Y��?�R�A����E
�t�B��`�<!GI�0i�<iRn�<$�4����G�<�*�Wr�i���_ʀ(gC�D�<�V@��5a< �pOP�
f��B�<A�ռG�Јɯ�	�,~�<)S�.Q~V����ݨ]Ҥx�k�a�<Q@�D�W��r�\!-�����\�<�Q���:������uGdT3�AT�<1�!]&2��a%�R[4�MKgKP�<IqmL�`(�}Je����@�Mg�<ٶ���f�	�a��IL����f�<q���ܔ � ��������l�<A&bً[�p��'#`jIJm�<�Q ]~ ��A?5:t�e�<q�MR%��%�׺3��� ��QG�<y�d��,�"���n�8Ҡ���!��<q�IƐh�P�" 
�B�ب�gTf�<�����
ތ�V/�0Nj��	^�<��	��q��L�k)
@�(�W�Td�<9"��~�. KĆ�;"�4�Mc�<� F�,H� 7BɨBm���#�y"���~�&�*�I	8S��5U��y���M�XQƋڐ� Pichβ�y�*�:F4�)�GV�_C���%�y��= �^�!�^1+�v��4��y"�0��g_"� A:sH]�n����'E�<���	�r�R��m7�1���� ��Ѷꂆwz6�`��cƆ%�!"Ob��%M�C��&C8wJ���"OPA�%S�r����Ґx�Vh�C"On�2��P>yB��i��̠��"O� �(E�m��d[�)0�ְ"OH�i㇟�(�آ�(5�x�:4"OԘ�G�ŎH�:+��$Z�� �"Oʽ����h�9�$��n��D{6"OX��p/��Fel� �e˾c��af"O �!H`^Ll�X>T� ��"O���a�Z4W�g�I�sC�0�7"O�]�S�P�I$�a���,<2 "OxDq��Q�",�E*�F}*���"O45���^1+&*�S�
O@��d"O��;ac |�\{��� RM� ��"O.�8# �:l?��AdFի0��i��"O<|	Ƃݲu5�`�� �Nm�a"O>�맣H�{p�� bX+����"OB���̛R��	we�@�"OBԺ!BKw��=!!\�2[0l�"O�(�"��oI���Â֒FEx�P0"O�H�bj�:x�B��rh�%HBb=�"Oj����żi��Ʉ��w7 	"O|p�BS8*T$��
�
'L��E"O�,�@L��8���8ѫ��B�j�"O-��fˉ?�`M � F�r_��"O~m��@5j�A%F<Zu���"Oժ$��0>-��$��h`��"O4�k���%)3X"�ǩ:��J"O��cE	�f��͚�׸�3�"Ol1J nZA�m�4.Q5R�V,�3"O�a�S�J!*Ƹus��i�^ds "O�5LX�[!��G�ӸA��6j.D���p�F�P���Z�K�8�ze��+D�X��˘OQ�`C�,J�	T�(D�d�րD����ʅc��tK�)+D�P��F�W�n�ao�|����f*D�`��_�B༐��oCX��<"�
(D������'*��ǌԏ��{U�1D���Ď>��3�N�P�����.D������z��Y�ŋM�V��n*D��:V��
T����`rЌ:"�&D�����ω?�f����I�t�Ѐ�`,&D�HCe��B[����F�1��P�tB&D���%/��a|䑊6f1`��H)D�`z1�T�[�R�p� �_��$yW
(D�,�TݣQpTE�˙	Ov�pq)'D���vM�D�8`�5�W[V�)cK&D����ĤFdI���%� X��(D���0�+P|� F��� D�!D��"Mϻ���-@,r\�=P�>D��x�.X��4�������[�<D���vJ�=�X�P�Aj�����4D�h��B�zT��I�i��X����P�%D�XY��؁p$��""��(��"D���#ן~�������i�5�c&"D��� �ԦR'Z�#�lۚ,�X�vH5D�(A�N������`�lU���'D��[���$XL����4WB�UqǇ&D� �A.G=r�(2#�!L�1�C&D�0P#fR.ŮQ
��}��D#D���"�q&�$�G�C��}ǫ!D��S�CJ��1�#�����³� D�8
�J��~$�5x!fO9�xEi'>D�� r�(UJ �����4$�`��"O�!#�H�����F�!|�=��"O�sS��zS�$P��Y�" ��"O��7,�����ccȺx�Mڀ"O:�8��J
t�I�않�"O�t���W��r�E��N�bIk"O|)��gR�V1B��e���
�:%"O�K�N_�P ��e#LD}~I�s"Ory��l%�H�Я�J$"O�T���"!64�go�0M�����"Ov\�B煀�x����̧B���"O���Q&�$-荪��O�LӦ%��"O�u�"�*��Vij�.�G"O^غq�ƑSrDd�@k\�&��` "O���郼|�5
��2RVI�F"O`\�rl�7�<P@�I�_�,a�"OJ�	�@֮P!R��D&�/|D0��u"OR���J�<"4�W%� Tʨ�@�"OdzQC��~.�Q��D�Yȴ;�"O聺C�4��[��"w���"O�Y�b.@�a9� X�G�.*ˮ�T"O.e��2<����l9��"O�Ze��.-0l�����`4�w"O�ŉLK+C�I�7�Y�Lun�v"O(�3�n��"(��
G�}@<�"O�q�Uoɐ��@���M�H���"O�W�� e1�U�88��J�"O P��ہ=�v��$�w�r�E"O` C5���F�̵ ��rrl���"O�����W5?l�Ar��F,���"O��S�@:P�h\铣�	��w"O�BR�?�f�s�'���S�"Ox�����c�te��8A�A�W"O����������닞P��h�"OF��`�4�Z�S�j
4d�Ց�"O,�Ce/��i��B��,I�4��"Ot�Qrΐ,Sj���$+�z��"O��Sե�4�|���U
�C�"O&��Q)z�5���C�� "O��eX�	5��z��Q9>�����"OP�$\!^0�\#!��	iIj�H'"O��@F_�#>����K>ZHF"O0�!��4m$;"e�p�2YH�"O
���jNK#!~���"O��C��m��(Cb�* �>L�7"O�p���Z�u���͛l���"O�´&J��j\@" ^�`p�"O�;BFP�:�\�9�%ߧ7WF|�b"O��"BjR�sE��Rċ�aP��h3"O�9�f��-tV���#�)"f83"O�����-:�d�p��rT4�+�"O��&D�2a����$�+m�6�#�"O0�i�jE!H�>C��)*�E�T"O�Z iR'�᱒����1P�"O�Azg,�R�< �qO�8Zi@"Oiq0��S�ԝ�A�U�!1�5�"O��:�I��Jk����,Tp �1sr"ON�@ �C�
�f]�a�Ԗ*\&��"O�Q��T�V H4�@�	4�I;�"O(��v�_��|Ы�	�<|k��I"O�l
CI4_��*��,jkReS�"OV�pI� &�"�A��ӮKzڈ9p"Oԓ��^�]��,�W.��/� �{�"Of�HaE���bs�� 2�L��A"O� R�k�K�b%Y�Ӝ���A"O.0��Gͷ��f�V�Z̳"Obq�&�&<�v4k��E���`1"O�1�eѹ%����F �Bz��F"O� J-jqRmC�`��cv"O��ielE�_���b���=4����"O�����*C�ڜ����6�ģ�"O�1�D>_#MQ6@Z�s�����"OJ��IO30WNغ4,5��5"q"OF]�פf�b�c���P-�$"O.<��̝.<�T���R	b��a"Ol4b��?���CA/G��ЋP"O����-��/L|�A#,���-�"O��ySA6�̘Y�D-#�4��"O�Iل��9R�,"���(|�"O�ik��N-;�,5
B�:kxT�3"OX:�f	�FJ<Z#n!a
,�$"O��A�,H6�����\�;&ҽˢ�|��i>�'����&ȑ�8B�oL�9 	�'��P��gB=mD����|�����(���q%��<y'�EZ��-o0|YI�"O��g�wNHRTGV�q��` �N1���l~���'��D�b.5;�dq�RJ[#zbt�'>D�T�HHo��Y�K��"E��'/r�G{���Rf,\;�@� 	/N`�EK*%!�D/&m@0ƍ�]P!��DT�(!�D�"�<�Q���m�T�pSD�w�!���3}p�r����9����P:�!���^ńx��%��5�~���L)&B��d���?M ��&g .~OX��d��2'�B�hg� 0�]<2X\���;D5�B�ɪpP����ږl� ���M6	�~B��1�RM�/ҟ0� ͋@eͨ�|B�I�(�� TI9�r�f�dELB�I~ZT��Q���\�k�`6B�Ƀr}���HF�2�dL�Tit�
B�	8�r|J��~500*D-�*��B�	\��j� ڍ:8����[:�B�9XX^���e��CP�:�OHB4B�	�DI�P!�_��
t'�&u�B䉎;���0�e��	�@K�(�C�	-��	8��.h�~���ʁ�J��C䉊|�͑�!ߐ)�TH1񋞷��C�>�,94��ld^	1)ȫ fC�	,Z��D�GTy�P勐j�A�ZC��[m" ��F�	g\�#��޷\�"C�IVi���2@M�R��M+"���/�C�ɌQ ���b��,��(�d �E� C�I�;.lAbӇL]�L�w �=��C�I�_Q�� 1΀�]&���r.ި����V����(�֋�
��ذ�a��+�� K�"Oz��ѯR�2y*e뜕b$h3r"O�5�d�Y8��5˒cόZ���"O���Ԣъs��a��E-�ڼ��"O��9!P1�fi�tOX"!>�c�$(LO^tHF6�|R�E/qL�`J�"OB��%�Z5s����?U<x�0c"O>����uzL�PM_	��P�2"OP��M���[!�ёw��C�"O6��r��,z�r9�3J�u�l�%�Iy�O)�S�% �n�����=9]���'�B�"'ۏh��E9s'Ǐe���'t�eh�Nڥ;��±b*�8�'�$�yՊ��xO�y�"IQ�\U��!�4�hO?7� �qp��j ��(���9j@ꉙ�"O�4�'��:Ko^5x��ͷ \�h�"O���E�Ld���,'�Tʇ"Of�i4���Y�R���D�g'��а"O`�r�� M� �O
B #"O>� ��v$C���|˴Ik"OB��s��0�0t*�`��3bΐ��"Ox�iˎ�>�8A�T C7}�X
"OlX1Pd�&���/H�iI�X�"ORX���)j� �ۖ�6��"O�݊Q�8��0�/
\�}C"O�	0��8&� �jw ��'̎�F�>��+ʓ��'G�%j��ϯ	�t B�/\��8�''ZAq�HSgz��a�'�������O��=E��A%e�\*w`<yg�yAb�y�ʀ:Pj��j	N�l�t!��?#�{��g�����ܠ�Д�����?I�'َ�"OA�2/��	`D�)=�N�H-O���}���Hg��-G�.` ��-�!�$�]A�4�lS �1���2q�!��XzR���e�ʕA�8t��ȓT�¼PR�;"�EZ�輇�~�d�E)��R�)R��1j:����=P�])�J�L1��� �+-N-Gz��~B C	>Y^����F
�*d�c�Sz�<!��(�,�C ��x��Ì�[�'�qO*b�<p��-V��X�&��Đ�.D��ɕ�=D�1H5ń�pC�1y�*D� F��0�8�&��2��&O��=�v��8XM��!�%�U���0�PM�<��i�3�])�H�s��XU�A�D�.#<����U!_g�Y:g��~�Hh0�%�z�<Ʌ�D���|Z��P�� -Xt����@%�����yX!��]v7F0�:4�d�B`ѽ'���$�"����B��Y�<���Dw�k%�E���8��T�<����8s�����+�?:��5o\U�<��#̿Ghd��R?c5��N�S�<&HO�'H�����>C4J�P�<i6�	.di��g����$�Hy2�)ʧe�<9���W�Y�JdG��ȓ"E.��t��.3�A�W�Z#`l�\�$)��<ڧc��BV,[r#`8��@L�|z�뉑��'�l5�����`�P��L�~ج�r�'3L�X�ņvT$�z��,,d����'t�c3h9B��Z�0)b�� �'=r%����g莝�a&�l��Z�'��%8���&U����a���\{Լ��'���┦~��U۰�Z5}>6�����'�r�S)�r�d�8`�6%�(�'�5�e���# pG�R)ߨ���'�m`G�??�yVm��z�C�OD�=E���,g��p���B͂1��2
�'���B㇕dł͒ ���4�ZJ<)���i�A��Y�*&'����眄z�!�Џ%�V��s��R�<�A��N��ax��	8�P��a"١WmS�'A�>(�=ç���k�� �65d���:\�J\�ȓix���MՁt3��(F���bT>͆��m~�,V?n���'�4&3���FǙ��y��A �d���J�
@j���(O��'#>�k�֥1�r R�R@j��%�>D�,�Κ�Z�֥Su�X:AP=�0>D���q�C��"��s��Q�&E>4��� �9d��$-�2�X�B�>"q{�"Oz���M[/�
�%!	57 0c�"O�Y3��
C�%s'AF�|6�%"O��J�O�AZ����b�${
^lk�"O��82��4R|�|h6b��zD�a "O��jD(wq\\zR�W_|��"O�)�AE�(�4TQ#ޑ)�֕!�"O`QmG24����-�o��,�3"OX,����(	d���ӻ��T�>D�|��N�9rI℥U�>Ҹ�K��:D�`�ԀJ-Z�h�g"�Vb��9D�0��_�Y �-�%!ΒR-(��
;D�p��'�.G�\�%��i� C�l#D�4�*� Onr&0���!D��C�
6H���p�u�����@#D�8�u��e��Q��p[���j5D�|c$h �'}�4�W͍*S���y5�%D�P�g�B�{�!)pC"D�� %�6D��ؕ��Sf$BF�#�M�v�4D�(�HC�2������\v��b>D���Q)0�p��n�1>��|	<D�t
�	�&�H�j�K�����g:D��s M̓p,y"�GN�e㰉pq�7D��p�G�q,���.�5Ib��B+D�x頍��m'n0��o���" �֮-D� )5��	;�ڇ٬=I@I��>D�`�EN�|3L1vH%	!X$E/D�����H:'d�q���K�l�@�*D������.3J⩋5�т�ܹ��&D�l�V� ���;'��+*�E3#D��R�h�>��\.a�5�b�"D����	F�3�0Gk�0��)���"D���'픔}C�Ġ6oZ�<��c� D�LA�U{ޔ ��cK�6t�3�� D�`񶆈�E�6���C	�Z޲�� D� ��i�H����R�ǂU��2� D�Ld�N-bB���" �t�nh��/1D�̫�*ίq/�|2A�M.sm0����.D��K ��:Z�b��K�-�\�dn'D�L�%9ʜ2�A&a�"�#D��:��X{���	w� Su���2� D��hW��~�4`3�ϛ�{Ƽ�1 H>D�L�7cϹM|����Y�x��@z�@0D��j�x~N9�@�؞]�T �Um9D� � +ʐK��i���t�P,�w�+LO����j�9y'��"噄_^$�3S����tA%�D��9�'"O �W�M�5�p�S/U�$�0C�"O
m�$�lԋ��o���p"OR(�3���9FژX�^JV"O�a+q͕70����F��]u�1�R"O��o�"�uI��ǃ=l�{�"Op�rG�&EGf] Ѐ�8��y#w"O�P���׾hb�I7� �s����S"O�=r����~���t%K:)�>-��"OJ��BXv��*�E�ez�%��"O�r���@��D�]�HV|��"O)�V�<��MqfCY4wN�ա�"O�5���m�e(U"��D�*Q��"O�=�Bb�=D�h��V�#��k�"O�h)�	 �oѠ�@��ԛL����"Oε�6��3�H�*6O�2��"O~�۴gH5{`-iD�Xh��"O�L�'�Eo �ppT�(F;��u"O����o�==�T�G)ՔALTH��"O� L�t�ȝ� ��N�1�P*�"O�@�D�5��4ʴUY�"O���3č�czٲ�m�";Ί�;�"O�ݒ�=hEH��u�z��̙p"Op��g��J��\ ���!@��ap"O�}+��wҮ����J�F��u�v"O� ;��JG۱�9�"O�IIWBI:/�$U1挘�v�Iä"O�UzA
�,U"9���=C&`�"O��ȳȚ�1پXI��/�ʽڲ"O���U�J�E���#�d�,0)ڌ��"O��i�c�2���S�@��B"O�Dsp�&1Z:}��#��T�6�Bc"O�P`w�Խ}�{���
@u��"O�$X�MX�H�p=�A ��S`���䆩2�L�ddAo�xAn���(ݴ!P�	N" ��G�2q����dF�V�!�DH7%�~h��YfkȜ�"Ĕ8��ds2l�'	��y��	.�LP��4oI�c>��"gs�@&��5}���(�n4�UHpd'4��H��@3��������a�����
6�W�~T�1� ޲m�<����Հ5`p����d��Q��Q@6T&}��,;P.ayBÀo#�P��%��u�R0i3���mT:�3�Ë�SL�h�$�b�s��[�)��%(%B2a��	,�2)�+�is������_��'����'=4�x����A�p�Pmϒ^uP6��(�j��D�U:s��� ��I�
��y�-�8�
y�Ӭ?P蠀�I�"�$�҃�Q�?�ޱ�s�Oo���n�$Zv,�dןꬨ�I�.�yǃ,pHRp�O�?�%�F���Px���Ɉņ�6Z�`�	������A��Xj E�.����#��[���&��\�z�iH>��M�Dg��if��HxwK�[8���bF�}M��2��B`��3��.�|5�֤�46Z�E���
nP`���,��kBP`+��%lX���	�r1��r�e2f�^�Y��D�[��'Ό�0#^
S4�t���ǲ\㮠
V,�7�� Cʖ
�lC���(θ�D
t�q��Q�3w�!��۬@�D��`�'2����jR�2L�27́�)�&���X	k�89C�#�v���B��,n?���f*S2 7D�w�A�(�<���l_��:B�E�l]�z��	0�~l��'Dj�#�^8�6�"SE��Y:	��:��-�#/ë3QX��5� eGn��H�=�.�Z��D+^58a&Dƀ=��q�эTu� ;&DYN���'�Kv8�ܱcؒ`m"����_�(�B� �Ì"2}9	R�U3US"� v��bSǐ�$MN�h���'|Z�,M�5rq���<�O�y�fj�={�]��) ��@�V�>�֯4W
�����h�R�[:�a��[���|¦�\�k�h`#D�@'�Ѐs�C
9�Zp�3�G�FMD0�,L�3�̡C�EWX�8�$����Ss���U��L��D�1JY���o��2")�n�OLl��Eȑ��(àBP��xȤ�JU����@���0��C2@�]���x� Úk�xk���\6�yx��W�q0��	�{LX�E#�v�x�9���n�nk0��Z9�E g.�v&���i&��Hd-�^I�}�HC�I2��dV�\N�U���F,]:Ё^�,��#е0nI�a��"Il(�B�
7
]K��W6��4f"*�,؀7 ?pu�I<I����^!z�D�)|���ˑG�]�	)~���Q�26����!!Eұ��'t��1�i�P�j�����3�B�;:@Y2�.Ad�m��@�e 28���#,O�xQ�%���y������Lx��ʔrO~�)�)�p� tbQ	n�H9פך#���m��L*$��P��+��&��:/��Z fO�: ������Pxb)�4Ml,�v���Ie� WhÆrV�I��F�k�����e��C��6c��p��f�ԌI�N�4��� �*��e��-D�X���������.C�<0s���0��'�L�vg?� ��f!�":�!Q��	�k}�������n�:P#ؑ"�T���;���N<)�j�$
�DP�f�Aj
᰷��o��h��gJI,%��pڰ�ŧ�%�B4�|�c%$��VL4��椃"C�Ir���/Q*�A�kA$J�.Y�B�(�B��Px���B�HiZ�@tj �k 0�%�)+�Q�dF��C�$��� �Y�Ԡ�"�ZKnH� ��A#g��Ȍ�, �]q�HY���0G�� 7���0>�b��8���Y� $��'�<b��z���6|�x*�߉wD��ƛ�U_d�w�I% $��X ��m��E倴�t:2�_�\`
�3�V�"��������X�<0���+s���w���(C6Q{�Aր$6T�BG��Q�yr��w��uS*�9!ږ�.&M�(� ��:t���)�)��i�VݳB$HӺ��n�~�ce��7Do��kRBK�s�*�]�{F. ���K1' �k׎��fn�=ȇ$�k��c�OW3�N�*E��P��ʣB��J N�>)�j�n̤|j�$
�@���=�7���sV88�ݼ>�5���;�1R�� �D����[�<�Dd:{��A�B������]�LG����r=�(YêN�$@��a�H�n�r��뉐dw,R��ڳ���؂�<.��x��+�P�7܎%�����(�4��ܘ�1z@��`�L|~�Ӌa�����d|>��f�G���Hv�N�v�8 c�	;�	�w�2<#4I�+h_j耱់eT�PX7K�3E����G��#�A�*[:�z�/ʤO��]i��~�	I�F��/�3}� � �F���9�����n ��A��n<؀�a/CP�����
0�và~��ڤ� ���D�h>��RE�X;aȀIб��#ѻ�p>т�"HL#5픘0�:��lJ�,��<"P��U�\�A�C��M�e��F���J*6mzq(�M�yb�d�T�0��.�&��FD��0=�2�Z�x��	R,S��_�P�2=���ͅr3T���B����	�i"����D�\ 8C���h�O��tF.L/V]��	����y��ʈ�������d���
��)�/L�2�8����xт�-���D�C�P�$���
6*��
 ���}��F�Q���H2Ό�,t(�K����x�B%(X ���R�'+,����i���(�j�<ܘ�Q�=tN���c�M�5�c��;Lx�{��Y��p=�vH�]5�(j�nƲڙ��f̏mu����#��tS! ��?�f���۳����B$��58��)���%��"�
!+���@ΧS��zb(�l3��s�>'�@�E��`����\�
���������X��F8O�U� ��*Q�ȋ�,U�&�'�}Z��Xk^PakӐ����{�)w��ic@,��*6��F��^	,X�l8B�ƍ0�P�!�<c����RŊ� qjȸ�ċy��K.��܉��N"b
r�3F�G�p�' @0K��4
��׺a��)p,O.1�P��b
%;p�?Ш9��n(v�@���,*��̈�m[�z␤Z7�D]���ئm�s�ڸY�OZ�u���� �O�i+��M���~�%E�nâ��F�z�(��樍�^V|æl��BW�(�L?H��xBg��*B�|r���xX��rA@<��-�v�AJ&$KbX$�I#/�\E3��'cM�x��f��tJR �m5§G:X퉃���c�3A�Q?,�$�z
�'���kҲx��ŉ��9��	��x�0	�'/�X����Sk���i�n`qO�$I�B�YUfՠ���WzII��'UrQq�_���5��#Z�l��R���h[Бp���Z�� ��lG�*���דl�������N��h�#	��6	"�D{���)8�"4�IR;7�tz
� L<�����X�aX�4(e�>[R����Л;!�ֈ0�e��iI� ���b"���'���P�H��))�1 
7�u��	FA�S����J�� :AG�C�ɔQ��ys��)���8����T�yq�i��4�$����pC���|�4�hܓ<����cǥmOh�W�ȵO����I'`�l�iwgA@:`��Ď�
��i � BI	f�yT��
d@�d� +ۇ�z��۲D}N]�Iè4tF���תިO�={��7M�.�"�U��h������Dε�T��S�x�r�	º4rو�'y�X�t��cvE����xܶU�'�F! 3k�jr��S)?\�P"��%9�nXHe���wm�����6 C䉗m���CC�>�Lx*�G:A/�\��Y�6�&��K&Qn�[db.�����;�D��E��dyQ�ף��?i�Ƒ�t!����썭kG�](�B	{����ț-��Ċ6�S-a|�f�9K���B��� ��˒�I���O(�Kr��'\E�j�O�6&�����B���&Y~d S���q�!�Լ4��8%�ՋzQN�0F���Y���+���(!J�8����II<^`x)P�MG D��DY�!���5x���s� �"l�����֋"]JX�O<�����G��>�O����I�/u���!2X�2�`��"O��I��BO�b9 ��YD"Ol`�.�+=�4���+�(
(e"O*��G�Ɣf0��m�D� �k�"O*u�WDH�&Ek��ǁ�����"Onh
T�޸b��`��#}w$i��"O�mJ�噑:I����x��:�"OHe˂h��/6z��&�7�D)T"O)��*UV4}p�M{h�ِ�"O�k��b����`��;\[�us�"O|\���U�Ơ�f�,D�0`"O�iô)W&Z�$+�Ԑj�z([�"O��ڰ�ɍC@�!��y�Ľ�1"O�9��>^�,\#�O��H8�"O��!1<i��߶.ÄըF"O  �$ęj�B���&0h�Y�"O�x�Fa��?�@����#G���C"Ol�ɔ�ͻ&���	G�p8�L�G"Of�:�J��<>�q궧OXɪi8�"Ot��+*���kI� �䛕"O���!�B<��ȉv��WP�@"O���H�'�����CI��й"OB1Y�m�7J�p������
�"O� \���"�i�tK!�ؠ��"O��S��#3m3%ʊ��� ��"O"��hW��.��W�����y¡���S�'z���2DS�y�\�}�T��T�������W��y��� �,��g��%���u�غ�yR�f��`�\kƩ����yrL�a>��V۠"��,j��Ɨ�yB�[S�KG�� ���Ff��yBO�]}P��0��>k�iv�4�y�!,P��'d��X|f�k����yR��Us�a��Y˴u�gDV�<��?l���{C�P>P��vcIH�<�/�b!T��ކ8�A`�-@�<�1` �]�!��*�x\�P,��<��k�'S�r ��hӀ��`�_x�<�w�v�Dɠ�JL8+���H�{�<��w����<Kh�1Ջv�<���^�o7J: ]�@�jD$q�<�%��D:��d��yF���o�p�<)``Ԙ=<�y-M�p^ q��'[K�<�TE�&S��@i&�֖���\N�<����)H8����U�*MR�<QU�y`z�;�-�Xg�Dk3od�<#�X�F_�9s�GʳaXL�	Dg�<�/-l�<�H�&��koc�<l�'��z� �'}��[�Hc�<Q���#8�vɸ�Gҫ?w��S5I�_�<ip��!"�&̲�
�P�M���Y�<i�F�-xGa�aB[�' ^����q�<��O�/�T���2q	0P[�JUz�<��I.�F�C���;N�,�Q�{�<)4,��@մ�@�]xpDx�,�]�<�@@��`<q���l|x�f�T�<Y�ь�9�HY�}�.���R�<	cB�e��ܸ��1PQ�#�MM�<����0T���z�e���c�Df�<��.�&�8�A<^�0 :6ITf�<�����zYW�O �Z��b�<)F��)>`˰J��U��y�._�<�W�3.NS�@+Fɰad�\�<	����4�dR�n��,I�@C�<���Q0�Lh���&^sf��0!G�<�w�E��DcTiӏS�J��7"��<�aN�L��Bd�tfd%h�h�u�<�Ʀ��, ���E/�D_�]�5& p�<����_�N�I���U+�k�$Nm�<��(W���,�rE?�f�Rg�	P�<�E��	�8��H>z�z`j�K�<1)�&d����R�z��B�<�Gh]�4��HaLB -�0 ��a�<Q������ٲ���?e�l���A�<yA��	V�WoJe��]��p�<�Q�=b �J�n�l�y!)�V�<qq�Q�9�4I��Ġ|6����V�<�'^3z�AX�HX�b�X���u�<Qg��Yl�58���3)��0����~�<W�ݝK�"��c,� e� �B��x�<�ӈӠz�):$�#Y@���v�<1���7VF�IP��B6s�H�F�T�<�w�F���# �E4"�(Ѐ�\K�<iG�؏\����4Y�N��/D�<I#A��y�k��.�zb�[�<yv.��,��Ef�'jJ����n�P�<� ��dH�O�h��T$:|�qU"O45 �� �V鼅p� \�tlf�"O� �uQ�:�R5#��YQ�Ĺ&"O(��K�{H�첰�ƨL�6�a�"O�=���aG�Q�&�˥�Vxy�"O0�H&B�6Y�Ų`�W/6�X�P"Ol�R�H��@]�p� Vt֍Ya"O��3�U���ퟏ"zZ �"O.�s�ü8Y�p��ɽkƸty�"OfD�G�#Z�i�P�\2Q��8"ORy�ɐ(w@`�v
ٕ-;�ա�"O2�s�O��l��؂eNV�N��Sv"Oz����=L��h��*%(�"O@d�5�N�381b���E��"OIق�\�����W�J�aT"OR�2��($ͦ�� �
03!"O,�+�:֤D�FD0�
-�"O�L���:W�|i۔LT�p^$r�"O>e�IB(�M��+�3-�1q��ٖ>Ɯ0��i�MxDm�$:��0�ڴ&O�)\�	"��KS�ȯ�*y����!���q�z5�L)+!�P"B��(�L0�,W2y�L��2BΥ#`p���4
�c>��Ӄe�uz���3k��zGjD8���T	&4�<��(�&�F%?U5��Â�Υx�6T(&D���
Fp[��t��N"J�zb���F�T�G��0ը��S� �ayB�6g�M	/�&9Fa��H��|f�y���'wr-�d��{���*���D�b H�2�=IE�A�a�Q�4)�>��� �n�D�z�j!!�X�Z �2i�(e9P�!P�Չ�,��^�9]n����OK��#"OD$�U�&�bo�-1� ��%�_��	��<,��Z��0�M��Z�'���ӭ0�!�p5�5a$�C"5�T ����2=<��a
O� "g�B+^j x�)��X`���[�| ���e��B��aeטz������)Sp4p��+T�'�:v�)r����$/�	w�H����e��R?C(�EЍ�/ʔmz`�H(o���1'Ng��a����$m���&n�z�IƏ��<�aB�m}$�R��7�2���hn��<9h�I �+�[;R��e��=K8���1�
����E]f�) 6�7c;�q��h¬5�Z�*&�cQ�y#�Ü>�$��$�0cn<!Ε|<k��BF��py� �B�YpG�1Aq>|A4��5hxXQn�x
8S���A��@3ϱUǊ���ҰkdVʇ�A]��ث`�t8��JV]v�1T��Q�Ա揇 H��p���G�:tA�I�n�jH �K�PRh�I�i�W���oF����f
�L���,�N8Ђ:O� ��3A��TR� ��m͑4��V�!��.n$ ��%�t{j�(���6��ł�bQ	zW̼p�G�Q�1YS	Y�i)�'�$}�E^�3�}��g�B���N��f!� ��D�Y'(Q��#��"h�z�I5}Ӕe�r��5�zx�)�<N �X�����x|�0����� ӈV���I�'�29b�E��8M��g�{?�0��R�QR���#�ޛ{زA�C !�,:e%O?=F⭑��}<�8R�Ӡ@� �r���*S�I�ė/���'�0�� 0���*����|xR ����uӠ팮s�l٧g�P�1h7��0���BGoW{wL)Xe�Z p ���ѽG�c��Ԇ`=6Y�4+:<O�K��Ue6.m���?G�e��Ǔ�_]¸PGT�^���3�D�Z~0ɵ��w�R9���N3?�RP�U��[TД8���ē(�&���*�2Y���0ƆV���%��P&ƐS����B���}�<�e/	#d�M/��֯V�*�p��0_l��V��?5�t9�b�O$8�~=�@�m���򤙒d�8)��ݫG������'[]�1�iR�V ��^
j�8�b�"x%`���k!MK�����1�Lh2֧LB��9𢈖�kRt��'$�9i5�U�w����aNN��zA�r�\�V"^}Y�H����<l�/*[~�;r*�+.�)�#]8T��B�8$�T�{GiR8��4cֆ�P@��b&<O�$S��ڐ�N|� ��9p�<Q�`��,�(�H@�&��%�z��KC���	����l�t`��
�"��Y��n�n��5�9dE��hA���2&,&��H!b�7+2 ��^�м��
' A"�m�`عR���;epŁ�N�A����0$7.Ȧ������}�)X�o?��<��$˶3 �m�p�^8$T��g�^B�PC��%h����U>x��M���K�0&�I��&�)L��(�XI�`'�bb��H �W;]NR��rI���x�E���l�T��:�DQ�M�x3����͎�J���l@������^���H���0=�x9qm]{7����Mժ�b xCb�!G̾�b�^*3t�yb�E�DŨ,��L�5yN��Q쀕�Vj�*�[�dp�"�v�`A�˅�5�X��%,�.�|(��A��R�]*T�j������v�B��n�&�x�`Q5�DD�$�h�8�bT,HDXM0�hE�|�@��O�0-	�捴=�U"��$�����㈻Kn�T�#@���Yr�;lO���ջIL�P"?.1����+�JxJ� �Ŋ!Z���2#K�:�����&#H0��F��\L����'ƛ�Gؐg�Z�rg��N߂�0�"O�  $J��ןV8�܋ K)$�
�ZJ��fYv�Q�#<
�̝Z��P*F�" �'j���٠V�D瓜>�X���	�"��1�@��P���ŁJgl�0�3Wt� KF�&(�l�#��,Ey�}���đI'b�`��x��]�"�J�"�3}%� aa	vb̫G��)sw���'��QA�Z��YpD���'X��RQ��#�}F������+7�42OY`��|RH[�y��`��F�^��5CF��*s����Ό�ho����Z��ϧwg6]Kc�.T��1�RU�<Aw�Ԛy`kB�(2�����h�r�<�rk�3>'R` MB�m��˓�]8��ڵH�R�E�f~�>i� Gɔ9���{ M�[,L�`A%D�lk�'�d�`Cf�)3&5#'�7E~�xF��6eD��Ӂ��qV��O�-񲣊�P�.��W���$�4 -�p?Q2��6&Vd̑�D�
�kb�u?�Ũ ��m�R(a�Ѽ"Q�xI��'2h����	�P�JsƠ�A����O�L�!�!�?Am�Ү��0�$h�Di\�
�N$����pGZаU� s!�$�9V�d �E�|8�P�qkX�SR)�Y�8�G�M&����R�h�����礤�f�roL\y7��4^�C�	�,B*%�Ě�|B2$�Gľfx�M��D[C���w$� z{^�vG�|��_QܓRV�LG��#sx�I�EV�N�.���ɃL� �s�%��o�)6�8�!�-R:S6�	�6�[�g\��y��!�&����WD$MY�@
O5�	�.�1�ў$U�L^��J`"��Emܜ#��1@�ZA�R�Q��8�Ǔ5=���H҃�j�<
 2-��z��,b(�|B�NY�(�R	�#B!�Zv�	��j�*a�T�2e��EP�#r\	��i��9&B��ȓq/t��aK˟;���iRʂ# �d@a��,��詣jJ#�2z���W��g����'�Ԩqd
A�	F��EU�k�܌r
�j�А:��L�@o�S X����ͻX�KQ�2��� YN�Ҵ�뉂z$t�7 ��q舠�L�%t�&�=��`ބ��9`��]�=-6��i�!
�Y�p�ߦE�N�Q$م;lh#s��
�y�Ꜩ_ֽp�mZ&�L��%D��?���
S�Mɕ��,Q\�p��*Y޵D���آ~�v�Xb!Z�c�f�2���Q!�d�1I�A-/	��C�Þ�s��sC�����J�2�%@�Q>U���"�	�G��0hڍ9T�<��#��Wk����7d�z0�,"�" H���x���UaUQ �Z"��q1����G��p=����4����'�I/�!HP�'���sS	Yx�0�DP�z�م�;�7j���&鑁_��X�m�Q�<Y�Ü<3�.��S!�j!<T� &R?aDAΞ+ |SQ��4Q����^��H�r�k���^�xA���*Z@&"Op�����/�:A�SH�s��%)�-L�dڲ�S�>�Ȥq�+ U��g�%* PGm Ge�lyà�&1hD���	�rN*H8p�L�Q����Ɇ�"�䅑	^��H!e2Ζ`�	�<��Js���h$j0��������OJ�����5��C��R8 ���6�v�C�I
8	ڙ�agٮU�!��j���{��S���*e6)����)����ʃmQ����	l��!�Hy�Y)B3s�!�ːU��)��h��o��E )BؼQM<�d� S���>�O��Yb��A�ƨ���� װ}�W"O���
q^�ió,V1wȠ=a�"O"-�v%�a�P	���9� �y�"O�����1I���y��
o�|؂"Ore��IW�YG�F*H�HI�R"Oxdp5��Om|Ah��E�x�fEW"O�p�MR�Ƅ	YD�03lȕk�"O @�C�9\��m���A�'Hn}��"Or�#@�o�&E*���4����"O�@kӯ�" >޴H�'[#XYr�@3"O��B(^�`�G^�L�&}Q�"O����L�<z��!� �$Ff�R�'�Ȉ�B�>zXD
 �\1c�"��'ܴ�%�̺q���C���o�h�'5<��U�4[�щ䋔�X��U��'^�Q�7fA�{�����Ṕ1�'{v��� Ƕ.F�����S�~�H��'{REr`�ܷ��]�&���h�6Ɂ�'u.غce^ �*6A��o7nѳ��� ��S�W9x��!��I��0��@�"O�A��G�b�j&��9"OD��g��&{6t�J+ �@:D"O�ay�C�|`�T���G�%�"O���P2)~���T*[ܩ �"Ob���sr��3���}9.t�"O��Y{���;dڍ`x�m�"O^; � 8�,l"DJ�+W@�3�"OfĀh�
2�����Z�"O�Y�SJˉ�p9뷡�I���3"O�ц#�@䀕�"lJ긒a"ON,���֨N$K��(;l8��"O|$R�c� ��x��N�I�dR�"O�H�?l���폰|����"O����`��Wc�rbBLv�S"O�s�N<��)�ٶ/�nxh�"O>�*���20Xq��)��%�ލAq"OT1���1dk�}2�с\a�i"O�M���ś{|�(�����yҁ�$'k�0����=�9�agP��yB���H�n���(��sq�=�y��l����V�-+f����Z��yEM�C
|�� �I����l��yR�Z8DU��Z�ǃ(��E;����yb�G�Ks�U�Bf@�{n���F�y"�-� ��i|$�Y3P
��<��aʷ3���q��>���##ϕ~�<a�(�#%L�y��LL����Ņ�y�<1%,��R���j���1��M�f�\_�<9� C�'�ĘՌ�
	&$���CT�<)�eQ,De�1���e �b�U�<y$-�!$��:�ā�W�%�ːW�<���)J�)bE�5[���PE�M�<i�-;��)�OG�+����FUK�<aV#\+M�h̰g�#w,=1�L^D�<��K�P4jCG�L�r�@�i�<4�0t!(,���4/F*�����a�<��@P�H�l��R��X)�"I�Y�<Q@iΦ��]�L�s��+Be c�<Q�&��M��Uu��%f��<���_X�<��)�<}g��JpĊ�B�<��g�c���.�<���o�x�<�'ػ6��e86�F>kȌ�3�gN�<y#�
1N�����@[�~wΌ3���b�<	E�Vl��ro�#��0��PZ�<�ElۈwQ���TK���Q�v�Q�<)E$P�|�`5M�[Z���H�<��H�gj)��	I
d���F@F�<�5j۪
�DY�D�T :Y��(�JG�<ɱ��6i�N1�kZ�g�ʱx��A�<!�i�q@��Bd�+�A�x�<!��Ҕ,�hhK������ce�v�<i��H<Ne�p��ɘQ@���{���+�M+	<9��+ܐI��Q� ��`�L̠^�MჀ�1aQ
���������>	��к�����	-����[>t���3��8h�%lZ4@��|×Ο�wdP��OG-�Q�"X��A�+[ +��'���W N2^� ]aХ�`~��d�'@�h�7�ڀN�:	3'Θ=)��Qx�'��	��Ӱs�ݛb)�>E���%z�(�Ad+��p��>1���X�̒ O�H����'���	�|�E��Qc"- tdE0��cᓾIP�%��@FT �0<��~
w�?Y�%��k���q!
I�	�d��&Õ[��v�r�$�&!լS\�`�g}��Tɘ'�L v	�*S�n�	�ż��$���N�1���)��<IQJF5_�9C��$6�кU�Lɦ͠��� f*���ƕ Z�H�)�'2$P��� �|�	
1�$��� ?{%�����C�<1�t�O��x"E,���VH&}0�I�Pm��Qi>�*f=�D�T>� <)zp�V�?M,�+�'�
�a���"��
	�i����|���V�g��M��%oF��L#=�,�j�r�)�S�7d�W�˗ey�m:c�Ѵ[����8j_�(��O��C��S�O��xA��
*$ؙp'Z�@��y�ORT)��4��1O�|IA�*ch>e�#wZ�L��V>���:�����?�Y�)ȥm��)���]����b�B]����	r�"�g?��d̚B���7E��sh�����0hLu{@d���~2F���?Yq�NF:<�8���Δ3&<��ƽ>����Gv��"}Qn#P L� �U�g�d��\ӦIk�"JiqO�?���O�=Q`�;Te	G��aؤ��Z����=YB�Oΰy��b[����`�Ne(���,����;P����c�}���Ol�|�s/ͷ2��C�`4R�*�3��C+OX\���i:b�b?��%��)JV�SqOߖ���K:DB��8+�&�yDJ���%k�P�}��C�	�?�� SW/G�-V���䏋_7�C�I�2��k�~�r��ΫtَC�(e4�3b��?-��3�+ ��C��\x�V��(Ͳ�����%:x B�I�~F�����ے9Nf�i(W%4WB�	�S>E3#���MN�YwnB���C��84�\7�&;��pS��>96�C�	;	�(@��1[�I=u��q"O�i
קÊq�*鹥�	�v��"O�`��,Ji��bF
?&��b"O����."�l���L
<�����"O½K#��4��Z ���Š�"O�s�A?]l*�c�DK�:�"O����/e�(���#ӦoG�{�"O�L�҇V�$N�(q�;�x��&"O����g�>D�C�1S�#�"O��R-ՓeEd�׬�`h�0 F"O��BG.8(|Ä�%E����"O�A0r�؟P��1��*		�zl�"Oq�d��wN \����7��DQ�"ON����ZŒ�
ժͮyɆ���"O��!S'�<�xq������2"O�)	Wh\4v!�l1�F�v�4h�"O�u(�-�>�D8"��#L��a��"O�Mb0@�k��Yg��? ̥��"O�
��7�a�򅊟i$�Pp"O ��.�	%����RE�x�k�"O�X�ə]�����#��
�	1"O�	��Ĳo��Yӑ�Ϝ�Py�r"Oؕ�E`M�g���
çR�t��"O�HZm"w"���)��r��G"OΩ�
D'Z���NO=<J�A1"O�Es@KӍ4P�IA�\"9?T���"O8�s"�['��a�w�ĺ	ѸeY�"O�Ě�\�l<�@	�4i�"=�$"Ox=�τ�l���S�<pz��@t"O���	��(QW�U'h�a�"O~�A!A7"����&��7���ʕ"O"���>�J��KҐ�ʭH�"O�U��ɏG2��1��P b��:"OH��t'�J�2�P�$��;�"O`a`2�g������~�b	ɤ"O�E�q ��:ݶ�O�i��9�"O2qxE�L�O��pyr��@�*)�C"O��QS,Ɩk)jq+@,�	=�p��"O4l�$�I��F)0T�o� ��"O��k$���[�|���È#�����"Ov���Γ�� �z� Y�f@p(�"Ov�F�GC����f��,\`^��0"Or\r��	1��a��O�^�i�p"O� \�8��� @�����*DQ�АF"O�	;�L�aYl8(֎����k�"O�!��i�x�V];"MŔV �0�"OL��b��1�.�a��Db R�"O��d�</X!5؅�"�b�"O4�r@(�F�~8aD@ռ<78U��"Of�Xq��i���@Ɍ��к�"O��4*[�ĜJ�e�"�
���"O��r�MP�f�L�f�֍P��Q�"O�t;Ǧ� 8�s��9F�<�"O4Y�a �m|hjD�Nq�`3�"OR�ZvۘjR
�p���ƪ<��"O4�W#ȂPPL��4��LŰ���"O������D�l�Q��1S�
�S"O :�8���{���?��8R�"OX��Q?*��xR���J�>-�Q"OR�!rɖno�H���,�h��"O�퓐�ͧ4^��y�h�m�M#�"O<m�n��@mXz��	N|�e�e"O�����=J�[/oz��Y�"O Y�ȡ(���
���"O!���\7q�ZhK�/�6!隀c�"O�酇u��iE.=U����'"O�z��[���Vg��*���QW"Op���jQ3q����cW'M��1�R"O�H;%�Fq�H���]�r�b�Q�"On�(Ш8<>|��,\��Y�q"OepQe�#�Y#yΖ��"Oj���9c�r��U�G�� |�"O�,9S�@?!��p�-�(��ѓV"O�裃T+��
gK�5f�6`�"ON0[g�S��\j�HF>#�(h�p"O��k��\�w���۹r�
0��"O��I�AIB��I�,]�\�]x�"OR�&ٍV/�Pl��&.P"f"OL�1�!lCl�DJV�z��`��"O���dj�%g�,r��̮}ݎ͚a"O��P�(I�q���)��9�^m�B"O$��R"ȳ*^a��'�8z�A�"OL�3DIZ�C��r���]�4q��"O���b!R�|t\�#�I3ȩP0"OйB�S�6�l�;��-"�� 4"Oh�� �U� ��f)A�lJ��"O<��eK,F6����E�eb��0V"O�"�DC��h��dɗ��`��1"O$��mG5/����hF<�1��"O^���HP��~x��	wE�a"O$��ALkH���a�'7�p��"O��I'Oʘ0���uAրOO]QV"O���%�K�ـ%��hI�Q��"O���JjG�e�N�D�0@��"O
Љ�CÞE�P���EQ*���a�"O�����5�e��G�d4"O,�i��Lj�8)�+�	 �$!��"O��`�
+,��V �-e�~�"OV�fb���̑86�'J�"O,�QϕJ��8�q$	JŪ#"O����	T� c�b���A
�'�eȶŋ�i�f��0/�-k�=c�'��jfGԝ�H; ��h|b���'���ʥ/jTx��Z�\ 1�'<��{��5>��ZǤS\�|�J
�'Lz�� N�?'��T��/�6P��eA�'� ����n$�3��U�;Q*�
��� ɂv!��/�2}r0@T_�|��"O0ܙ�j�9�8�6�GU~��"OPd���(k2D��gCoXL�R�"O�qg�HS~��F�#�B�7"O�(���?蘍;��Ѭ���"O���Uㆇ$8TE��˿Ex��V"OR�;w�JK����#$4��%"O^M�S!��|⃁�`ⴭ�`"O|��u�F�x�j�:�DU�b��B"O>�#5�L�Iv>93$�Z�_�Lث�"O(��ѦJ)^eǏĚH��p�"O���9A���$AD"C��Pht"O"I��卲i�~�����X~(�"O���i�/x��lbgI�4!R�\{�"O�ac1���6�ڵiR2\℁�"O�`��nʭ(���5�a���"O���zH8�'�ba��;�"O"�ɵ�"~ʵ������ks"O�a�.N�%4͑U�Ͻ?��3"O�LAS^�9���q �������"OX��0���W3z��n�*7�ҕX�"Oz�;�M�>:��H �׉�(�9 "On`���ڰcذ���!�&x�؅�R"O��g��7t����Ҡ1oe`�"O��.�a��F��VVt�"Oʑ���F9���O�o@f�Be"OƁ�RF�p�U9��6�H��"O6蚥)̩Qo� �#a�/u^J�"�"O�iV��y�V�ؐ��a�V��"O��B���$2��EJ�F�V���"O^Td�Y�MPp�n�(��]Pq"O8{C\{1�L��D�p�4��"OH��G�	;�8���BZ/#X$�["O���E�ۀmk1!��\E��H�"O&����ӭ"�X `�����"O޽�uM¤P�>�!1��Y����"O��+HV*����3���P�"O��Q��	�}��q0礊�P�  C"O�����-p:<`���:7���`"OK�c��p\�Y�v����yB�;�<���&gn�h��.V��y��1��%ȷ�O�[Qh�h��y�1&;l� �̥T����Tg��y��ΤX�1��oֱQ���3g��y��N�����*��J*�,�#	�=�y�FE<x�&��G��ȡh��y���^���@R�ѱE2������yҪ�y�a9c�N �T�îU��y�ѳgG|�����v��<[���y�,�12\-"���0rfr�y.Z��yB�3\%�TJd��m�*5�"�O��y�%Y&t�$T��<i �����yBV#F����˃�`}� ����y҃@5�(!xb�E�S{f�bV:�y.P�Wp!�@��X�!�p$���y��ܾ(xR���:a��i	 l�=�y�KF!TPB��pR44��f�:�yrF��y[(�[K�P���r�f!�y��H��L�� N� *�.�y¡ ^mر9V�ӽ�5ڳ�� �yb��%1?μ��
��b	z,2�H�y�Ϣ\<�c SZՌ�#�Bش�y��~����`\�&
�%�E@���y��Yz�(+�P��!��P�y
� ��%�M+m��Ʈ�?��U "Ox(Ȕ+�@ܕ����0M�9�0"O��E�,6�̽�G�#hJL9�0"Oڜ+��	 r�j�pGS|�= �"O� �Տݖ~Pd�V�-O[4L�"OF��g\��!�s+�,- h*4"O�Q0F� |���
ѺZ8��"O|��2��t��Ε�'���"O H(k�*L����G�#���a"O�}JaC	�J~�x�P�E�1��Lj'"Oԝ"FۈGY���qP�N;��s"O`�+��N���D��K-T���"OR�pql].i��%�6L;bJB�b"O�$hu���O�|5��!Na�"O�� ��0��2�ݙm�>u� "O�eCN)I+�U�@�F�vhz�"O΅���	&T�Lq W#Ԭ��d"Ox���ٌm3b���1j&<�7"Oj�CE   ��   +  S       _+  �3  �>  �I  P  LV  �\  �b  #i  fo  �u  �{  ,�  p�  ��  ��  D�  ��  ˧  �  U�  ��  ��  *�  ��  m�  ��  ��  s�  y�  ��  �  J   Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�� |d��"O
`�(�;���8���-0��1%"Oj4��ND^[��"3/9�0|H�"OB���H��*�ʞRy=a"O�味V�!X��!&F�:J�$���"O,��a
���C�Ą�M�"O,$3%o�-���p���+Ն�:1"O��ݢ1����`���y14]2��i�<�6��{_���c�H�`�fX�$Kn�<��A̼VI�xR[�)�Ć�pඤ�ȓA5��('nߡ4�� �)˩%� ���,��r�؊b#`T�eT09���ȓ!�b��g��}�8�F��-? �ȓ
K|m�ș�VṔ���2�%�ȓ"R�X�j�4JN�1�˘X�i����̹	_�jZ��1!g��zܶ��ȓgil,*�J�
j�Ne��i�J%b���f	�(U��:���G��$Y^م�~r�� S�%T"���k\�jx�ȓ|4�1�îJb��@ӵ�ݩn�V��/[`�"�v4�R�!ʎ<��M�ȓ`:��z�ؚh�J�Z��$HY:	��H��p�m�C1��!��B:��0��EnjZA V;9����J[
2���	��4'J�EA�IVW&��~�(aZ��ӹ�>� o�Y�|�ȓ�f�A�
Ο7�H��M�$�����mޠP����/���ANXo*�ȓTv�����{ ��-7�*h��I��sB�8�8���3����ȓNe*M�悡;������X�o��!�ȓ'lj�#F�m�+R&;�|��2)n�C��0S4���T:
b���:�0!��e֊��)��ͷV��,�ȓ0�&�8#���� ع�L�����;�P�AFd���,w�6dnZf�����h�%��p_�E�T
C�8!�$�x�h��(�d" �Q��2��&�	a��~r�){2`�T-܌$N�YUl�%��xr�G�J�6����S;:�����L�E��B�I8ei� 1��0^�+0�]�����`������������	�+��?�~E�ȓ[������Ov�1���H}��Dz��'�����[=V���kCN�6.���'��8��䙢�4�	#Z('���C�O��O4���DBqrg�goVYK�M l!��(+ɬiwb98H؄����z"=y�}|0�,ǵ\��)��oY-|���>I�yR���OpRW
���`+P	�a�|��Qj�Q?0I(Ri�B{�s>�z��H���@�
��o��� t�ڂy����&"O.���$r3��
. ��D"OZ���D� Gr�81∴U3^�a3"O�5��/ �n���c��g�Ji�1^����	-���1̔�*�x���Y@b�pG{���m >`v�mj�)~�Z*4�~�<irE�09P4�i΅M��l�g�s�<�V�ޱ�f�äJ�(4M��o�<ه`�%z�B|Y�� �~�1�[�<����(g@,�V$[tM�5�#hO<6�nB�	џ������P ¿L^�H����y���O�X�6D� �P4��6�+�Q�|$����3� �4C�b�"2$eJw�p��9�v�OR��I�q4��6���0��`��4�2����b?�Ex��吃c���
ɟ7SZ<�ȓz�fd	$��	�~C����T��E��V���%�H8��$c��H���F�ma,6|OT�$9?��a�/��]�aʏw)|��g�?~��IO?�����B
��J��U��@�/�2��f���y�.mP9�S#��(���@��'Ma{���L1^]Yv�^,Ve��f5�?ً��	b�n7�m�\m�r��<1`� �`C=�� /�Py�+�B��@ɤV�aD��s�D]y"��%�<�)BL�\p�.7��r��̴p^!�d�O�]lՙ\f�h[&�U\�.����S�lR@�D�j	�T���nI��Ul',O
�<Y�nF�h[t1rw&5�z!Z#Is�<)TAV�-*6X��Q�U4����m�'�ў�1Fd����ޛ8;�"'"T�]�͓��?a�]U��P��K'B��$"M?ي��S&m%�����ı���kە<�B�I�t;� �6�TwL�M��G]*o{�ER��ʚmp�d6}�.'��`B�'��|�^��W
��u16<��刟x����#X\��"j��KԺ�����4��I�&LҤ���ѩ�,E!��]*Cɉ'���b�S�'<���!�L2a!\ʐ���葅�=�Q�g�	<!��o56���ȓ�"��rL#"���%�C�S�r@�ȓ!�R0���K=��Xy�L�/�d���?v�~�e��&�\����NP��RrF����=�y�o��C8�"Ud��Dܛ��S��Py"�N0h?��c��-(� ��E+`�`���'�� q�EP��B�;f�;�qy�'+����JҊ}Y��$�N(��'�h�1%�0��%;��Ov;���'��*��Q�A�\��3���A�6x�'������"BZ��ǫ�#J?��Ӯ����|xB�C;Di���D,!G����¸�y���zb��"r!�A�N\P�d���(O ����P�Vmh���+�� h�O
�P4C䉉-\��Ҁ��#\H��Ŋ�B ���,�S�OEƠ�"�	t��PŅȚ17P*�"OZx"��(O	Dd0p��*�V��7R����� ���1�:+:0�B�V.� ��ĩ<	��[�s��Y1 D�Y��*	�w�<i�̳�j��kV�5�ՠS�r쓴���O���IߙA�.xS��Ti��p���6��~[����斺X����`�)x�\�0�	�O(7m�ttqO?����}��H��OT��%�H�'�1O$�O�-;�ĕH7h0��.y`<�ش�y�e��Fx���*=�{�D���Y���#��>��O�)�O��/X����D_�"�Jh(c�|��'+�!C����8j����C
Gq�,ʍ�D�ȟ��J��!���Y���mD"O���$�+dTf���_�����9O��=E���R�>a��P�a��W1b��m�/��O��D�d�^�aC���ЩE�H�Ԩ0N��yb�	�<>v��+�D�X�r��]���>i৹>i�(�6d¾�� Y���g�T�<6���w��(̓����b�h�<i�bX��D!�+9?��T!��eH<	�����is�FU�W�����˽g1O�b��Dz�%�(v����9,
Th��x�exӞ�c�l��3?n��g� 'ˈe�"�>���)��(K��EԳ+��Z�G�s`�O.�O�"~*'@ q8Q!�Ϙ0M���k�,�E}B�'$�|
� �I�m� �(���숲^�r�g?O��Ik�S�OeS�g�m�xH��S�k�t���'��+�c��W�Xd�c��(#�{�8OP�Ot�S���\�Lۑ�Ηe��i�Gf@��0?1�'���*`K�g�B�Y�$��j&������B�<��
D:gݦ�[��M)�Aӵk�d�'L@�E��GP�sԄ8 �� �*Ȩ�˜+��d �OԤg�Аd�8��i��6�:ҡ�'�ў�OT<�O���	���(U���H�<�`'"O �j�o���D��5ǃ7�)���'}� �OzPc�]02mx��iN�$��h��'��Ov��d�5nրu�to�u	�l�6Ox���0>9�����Ii�f��%�,Te�o�<�!�'~��xc�.:���*wnIk�<���̸i��8��O�, ��0ч�p�<A�NX�-��܈��c�����l�<!�ϕ ")�!"�h�)�H\H���M}"�)ҧ3�<�3C)�>��T`�=�͸	�'�Wd�D�]@�d�JDڀs�a��~�R}2�1����P�8F1�@�R�xs�W���>i�:6�Ɖn%�|Bcl�Z�����Х4�j���M��O�(��^|��K��9L����$�N�93�c�ī�&�	|�3Q�"�R�ܱo��]�Ҧ�'q�C�ɴ|/D�2�X��=�"��B����7��?�<��P
�K^4JfT�d�I�o����Ms��:��q�!b�'��8 �@}}r�'�0����ބ`��]r���TaF��
�':�3��0����Jޙ�D2�'L��q�M�w<:0񀍻#ұ�'�,�a�Ea��q�s�N �a��'���i��W�|
Z�&��\��%i�'夌#�K������@�I@�-��'u�;"!X28�<y!��7�l�(�'���Ss�C�"r����͒�4��'�0�U�"QD��	��v�p�x	�'����3aZ�:��g��0 C@a[	�'3�u�)SU�\��JQ��F��'W��i����Hu �� ��w���'k&yz�m#!+�Dɲ�(m,a��'Et�$������Q����Ȅv�<�6��g��I ���|Ԇ��ӏ\o�<9c��K���A�U�g�H��
�i�<Y��4R�E�b�F1B�%K�<�\�ll:ȀJ) �����D�<�V���L܄)J�FG�S�(�#&@~�<�� =�8k��6mp<�n�}�<���ٔSf��+@�"�uC�w�<��Ҡbp�敞U$`2��9D���ϒ#n�U�A�;g��]ɶ3D��r�GD<*���cp���@r�1D�d��&5$������&z+���.D�� ��Y�d?(��5�Զ4hx�a��1D������MP ��S$;:�q2�"D�T����a$:��r��6_���v& D�tzP)+̅[�-M)U�Ƥ �$ D��z'�	XL⵰��L<;�̚!m"D�X[��ԭ9�Z���?�(�A/,D��xS!� ���bd��9'zD�v+)D���կC�A6���d�y�,0��(D� h��6f6x#�_�|)�)Ǝ(D�<�1b(i\ ����®(�XP�%D���$�_6J�l�@r(K�F�+��s�!���a���M�+5�j��1D{!�Śjv�i���H�֤���\,!�� L���ř�� ��U�
���%"Od!�'�J�V��)�fB�/16�ZF"O�� ��L�L�[V�� �r �"O��F�.>81ڕ�	�\��j�"O@����7M��y�i��8�͉��'T�T�`�IϟD��ß��	ɟ����/���T�Vw,�4Z4%ͅ��1������`�Iϟ���ȟ���џ��	�=����Sb�Hd%V*q�8��쟌�	ϟ���Ο��	۟�������4#2$2c�U�{IM+tm� ���	�,�	�����,�Iퟸ�������f�0a�Gwx5s���/O�l�	����	��	ߟ��	ן�I����I-M���c\�&&=�IE�C6�Q������	ן$����<�I������0~���I:=x��o�q>p��ҟ���ǟ���韐����\��ҟ���=u��@�� ���y��3P�����ş��	Ꟙ�I�(�	�h��ӟ��	`.�@V�^��b�U�t�	����ԟ��Iݟ|�Iß<�I����	�lx�l��}���ńHs�x��	����I؟���͟���៨������?D��0��S\V��B����68�����Iҟ���ǟt�	ޟ��	�����,sP\��шF��hz��@�]ȥ��џ��	ӟ���˟��I����	��,�I�>R&��n�]ILY��$]�qG�����<�I۟���؟��	㟤�ٴ�?)��>�¤f&Z�iD�$�a��Lo�	:�X���uy���Ob�lZ.C��4�%e�"��*%��,m��!2��+?�b�i���|��~r�i7��+Gۗ|}Y �@;/��#w�j���DL-1RX6/?�����x!�;���]�n�{b+E,p��X��JA��'��Z�4D���1*�th l>���Hi
7-D�
�1Oz�	"�iO����e{�<Af�O�+�T��P��)>��qP���M�'�)���4Pe�6-s�����I6kL�%�����P4(v�����hl�Q)�mAU�����'�:�甁:�)�Հ�l��Hk�'y�	C�ɐ�MS��Fm�}�p����  ��D�&�T^�x�����-���ǟ�oZ�<��O4b
@�18;���	r��E��ppvgÐ$�*�3��=擅'򀁯;w�Lԩp>J�#��ρڨj��ֳs��	{y�����󄝕?����CQ
4>j@�c��5m�d�Φ�JQ�'?�P�i2��|�O�����O��(!&����~|��'$R�i�b���V0�&���"��Zm�	לJ�r-
�	h�J�=&��E{�O��h�S�5Gh����\�@5"%��K�g�b�qÛ��1И'�����4d���Hh�
��U��YA/�4�˓�?yܴ�y�����O�"����aN�xd��I\�` �mRxю��'r� �C�n�8Я;<����I� ��� �i�ࠂ.�"� �IMy�S�$$���4]�5̓߶��S��(c��:��>tN���Gf�v�4��$�O�6M�O�8�1m�;>�ک��g��\�F$9�M ��7s���kW�$���P��ЁuO���$$1�m����\*`���s�IK� ��4fB�<	�����<E���ZdW�y�oH��@���¹��'��6-M-�� �M�N>1���z�>M� ��7�63�
���y�Y��n��M��lW�1ߴ�yb�����U9��H�%Lɞqd�ʯ ]��;q��L�R\�L<��O��<1�&),|:��F-}jL�e랠(�����5���'ŚΘ'P��V�$���b�0��K]��]���n�<QM|*��^.�� �S$!�*P`rK�����ٵም^{��u˄S~�O��c�� %�(���-h�l�qCơ[r�0`D����՟��П��?�lsyO{� l�d��s_����7C+S'��4�d�O�eo� ���Dû>��iCZ ���3\|(㈐X�0���Ʀi�ߴ�5�5V�<�?���c�6@v-p(O �r��8�r0Z���<��<{'���O���h�by�ÂA�F��tre䀕n�����l���O<�	l�'@��w�<%£)�2�̀��@'�a���O�6�c�4���l.�#���<	Wi��O������dW���DO�<!�J��f�и`6e�!�hO�	�O��k3f1i�(	cG��p�C�?O$ʓ����FJX$��'i �"U�lJ�43��3A���K���M^y��'P��4O�����,��e�(�ҡ�O�d�@��'�nsu`ٽ�MB��\Q�԰;
����ק�)~��v�+�^Ejb��̟X�I؟(�I���D���')�)9����V��Y"�FzNfm���'-�6�ÿ<���6�M��w��ypӄJ�R�X�{F�$N���'%F6��7zr7m��5ʎ��@��\�5�ֿLZ�ͻg�M:Ő8R�ǔe9�H���[6Ae��D{2�'���T�S�Y��"��=D��$(a��jZ��fʛ���ޘ'��2�kR�z�)/L��Z�CIyB�'��64OL"}�R�B"G��]h�@(p�j�H�,&�Rr%�_S~bϑ,Z�����R�&�ў��6����X���Laa>)��*Y��x�'|�	~��M�u���<��aİ!t��h	%�����̎�<�&�i�O��OV��y���H-h�5���/iv,��B�%i��A��B:��IKRM�E��Gq��ܮq�? ���eF�0��U:��D�p�0u�!;Od���O���O�D�Ox��$��T::�����܄PĖaH��.��Iʟ|�	>�M�ׅ��<!�D����|�M����Ё��#�V(IA�/F���$�>�ѱi�7��h84��t�D�O����Uz�������%�U;6�O&tz����&8��=9���D�O~���Ĝ�F#�4P�+Y|���<OΓO�l�u��b�����?�s�h!� �V�"~��8dd6?�U[��	ܦi͓��'�J�D�a�~l��J��b�-:�"Ūy��sd��d��0�'�����p��q�	J�p�B@�2�l��k��V��E�'��]�b>�5֛�E46Bȁ���/H^���)R�D0Z�r�Ov1l���$�泟�l��z��ܩ씈*6`�!� �ش�?�rl��M��'#�n�s���`*����X�f��6��6?V�ʢiշ_A1OT�D�<I��IH�~���
"�� '����"4$��oQ<@b��S_��MϻN�4��C��z�,���� 4D����'��>O2��?Q�����W妹͓mвd(�A	 ��E$�մ/=:��4M��L�B�>M��4���D�8�"��V &T��x�EN[g��<aK>Q�i�0U[�yrlȘE{��Э2j��s���#���|���<i��M��'?�	�r���P2�T~�v�Q)s!��	ɟ���W8X��y'�1?a�'Z����Zw�B�d�m'���`J%.����7*�$ʓ����O?�e�y u���/a���e� �I	�Ms���c~�,m�H��;!�`�+�	Q3\9� j�
,h��I����4�?!�,"wBd��?�A?\��P"GZ�h�2�dv�4�q��m�-���4�ʓ��P?�	!������(��e�X�'%�6m�#b�1O<�?)*7�W Z�H,�w�P ��3��K���OB7�|�%>��S�@��'��V��L�+C` {L�YB:?�W����3��	҂�=!6�X�S���S6��
Q�
 �3�ޢ�?1-OF���L��vd¢�y����C�!)C�#G49a����ynoӪ�泟l���9��
fB2�����С��$|V�`1�Ȗ�)���֟��g��`���"?	�':k�vt� zG�\4BX��OƛD���O�˓���Q�}�6�$}8px�ӊg!� 9�I	�MCE��r~2&k�H�$�<Ѱ�W�9��H�(W�H�Ů��y�^�$mZ��Mk�:Ɏ(�(��<�� k�Xh��5J�Hjm˝9"p4j�n�$<2��S�d,�	W���Q�?'�
����M�R��,D�(�^0R��$jJQ)a �"S��p#(Uj�t�VDR��|q +j����J,{iL�B�({�y�HIdQdm
A���¢ҋA��� ףO	{�N��@4��D	|!���k
m�h� ׁU���`�ԐL\D�F�D�3,@�Ð&��>L����AT2�P�p�&3�����z�~�d�O�����X#��,eq�q���*(Cҩ"���e�	ɟ���J����	���	~��V��4�Jt��怸��S�H6m�O��� X$|n�	��h��:��D	�R��s�.��-X��B����'�����2�'
��	��NX���O_�S�0�R��ޒ3��l3a����4�?���?a�'d��'w�� *e-����Bd|`���x�6M�\�����O����A짾?A��#���d����Hss[�aK
��Mk��?a��UjL� �x��'�B�O&��
Lb��ĈơC�G[�Л�i�R�'�r�%OK���?i%�����˓o�{��I�[�q��)k2���ȓW�a���T��.Dh���Bk�ą�I7�diIИ%{HIHf���qC������h�D�!cϋ*@��v'��s(i*��R���򀖿ek��p��D��ey�fđs�)��A  $�"����u�"���b�=0J\���6���Ć) �E�1��}�� �	���!�Х (�@ˀ/U.����3�j�q�W-����Oxi�.�O`��r>5��c���8PL�yIK]|bĉ5�qВ��?O�M�b!�W@ ѦO�Ř%�X(R�lN#�� d�'bR`A����6%e���d����T(ҨD��r�7Ib��?����^JʞZ�`H�Yp9��"�
<*!��覝�f�
6��y��/���Hd���'a��lZ6K"D���O��'�̽P�
9DA��E�fp�B՞�����?��K�JM��򌄚�?	�H���I�|�D ��'��<ѧc�tNu�`bDB�$�=!V0r�牑2�@�����������0s��;-P�xU���-�F��dE�>���'Z����?�J~rM~jm�{J�s��A
0Od�����OT��6\5���%�U82$��D۶�f�=�'\V��D�(��FP�f\�U&~|��,���M����?��-u��3J1�?����?Q�Ŀ{U�C�{t|�����2�Ҥi5��,ט'�,@�\�qkgg�<4܍鑭�f��A�=Y��jx����!��d�I��Xb6�ß��'�4���S��|��ҟ��B 	@�	 D�2|&~��1�NYh<a��R����r	Z{\��� \~B
-�S��P���K��"���U�ĳ(_HՓ��� D~ �"ҭ������L�	�u'�'��;��Y�� Z�RG�!|���!�n
�Z��Ã�X1ey���$/� ��`��C�0L2��[��@Qs�΂"')�(��g�>N.��1�T�.��s�M��n�$�O�e��AҎwb���)�q!�޴lg�n��&���I���?��]��d�ELژqHD� R��o��'��[�$�v cp�
�$��u�D������uy��G���7�OZ�dSM�B yWfP3ni�G��!Fj�$�O~�H0��O~��z> �`K�3C���&I�fa��Α�R�@D��.F�t��v�
�i)��Yf�
.,�Q����J�;"�Y��_	Ti5hJ�R9[JId�5��9UЧ��)bϔ$ �H�gR��P��9�	���=�f��	�)��GU�5�ȓ��97k-H�~�
�	Y6�=��n���/�>n֨`�0 ��cq��U�E�@��'��R��e�����O�ʧ<X�0���c�F}����! � ccD��pN^Ij���?�r)FL�j��T>��O�`li��Y��f�C�!^.J�&4@L���D�O<k�<�)Ӯ��5�T�O��ۼm`��3����E�.5h`�!����'m�����1ɧ�OZ����хܑ!��TN,�P�'g�cm�t����D$
�DX����<���ie��3��yBE?O 1�eJ�Mk���?��T�j���χ	�?���?��ӼKW@�O!��PB�(r�@��_,dG\��W�u�7��6�A���|�D�:@q�i����-H��[p!�n�z硗�Qk�o��Bg�$�a��|�)={S�(÷J,�n��BFɤj���O`�������&��A���a{r�D��]��	�R���Cκl0a�C����'xb"=E��Eգ3/mA��պP�:H�����y��;=TS`-W5C����蓼�y�Ç�@,�� ?۾�[2M[��y�É����&͚9�I1�DƁ�y��9�4�I4�2�J�kb'
��yb�ޕ"+,e�T.�()�@���+�y�"�T`&O6P��SKG�y����\l�v(�	Ѵz�EŃ�yb!��s b}�Cg�yBv��b�
8�y2l�/�����Qp�'��yRJG|�̜
��(oD>�S��2�y���0�#ZG�=Ȃް�y��DN�i�5�\>J���"���y¬�O<0 ;�o�6F�v�x1a�$�y�KCsU ��a�8?m}�cMۀ�y2�ۄs�m��i'�a�P��;�y"�@�f�T"f0Ј�� �yP�w�����C۾W<0Y�j�4�y��/�xk�a�V#j�!R�>�yb-�$JȌm�!+�S�~lz����yr/��6���"S�H�BaJ$�݈�yb�H ���;f�
(e(���2�y���":��, s�H������T��y��� z��[����|�~�C�֟�y�D[&��s��J���쌱�yB����r��E�鷩]��yD+z��A:vĊ0���`d��8�y��*N�i���S��`�a�&���y��'���S�c�y�@4j'i�,�yb�8&�a�V�T�t��"ބ�y2�+�����K�-{$�h�`̦�y��r��0��ȇ^�X|q�%�y�+�N�����S2�i@@����y"!Q�Dl�`���^��W��yb�Ǜ#����	��"黆a��yROŲl�X�Г��5�֌�*�?�r�E.}I(�2TK�*M� PG�R�'r���ȍ�=F^Y;2A��hu��'���g셕c����ՉF�?�r�����/.S��b+��a5�����7C�@��6��{؟�Y����J�2ˉ�2P���I@�E��p�D��@8�B*��y���zѮ�C'-D44)A�
!�p?�F��KH����7�j@:�n��m���i1o<ғ9c�Yp�ϻ� J�DĖpȵ�'��L9���'5&�i!+�\�ꝡ���ܴ3*yPgjA�V2R1���9z]
� z��eR�@C�� �r �z�iۺM�`��R@X"G�$O����Ĕ;�d���Q�I��[�G�vV���O�L�T�΂:(��f!2ў�Qć�"M@�Ҡ����d��GN<��-Ј�D��?�"�0�)�?�y��� ��@&%
%1F��`O��MX���B"�'e�9�)�5v��u�<�CЈ
M����)��'�"=�';$��h�I�I���! �|z��rg(L ��#=�f�� _���}BF�1.k}r�L�
��p{��
�ÁG׋�(Ot��\�JX�qy��*V����O׫;W�j�h�R���Ux�0�Ã��M3�K
Z"|Pa��;&C|y����Z�'����ĉ��R���j���>���i�Ox8)с��/�i����/�����I�^�!+r	Ϧ�>Mȥe�[�U*�	���O2��=��CѬZ=>Ys�C��l�̢� �#~�̨���p<q6�^"h�Ί�B���y�)��+��P3��� �qO��=ͧi��XsS��$_X�@n 9��ܨ֬����"=a���o,v!
3����nUiRL�j}b�џ߸q��oK�V܆����Q*�?)��'.}�5k�e�O����I�/���c�'l���?1QZ���2.onyAc�ϦQ3�/�
�\9[���o�hm��n<�o�
YQS ۻ�!���5-�<��'��6�ӲaD=�ڴb��@+`M=�@T<kf灂t��I��P�Q<�cLՓ&�џ�������x<h8��e�^�� ��Q_�6�-Gu���	t
���O1ڨh�,P͔�P �p�4 �{�O��'��&$cb�SՊ�b|�GL\&U�|D��C�=쑞�cC�@,q���!"&��/��x{�)�>�3k*�i���A�eb�i0Q����O����Ofl!DmQ-��9�D\M�
8���'
	��BJ�?�ꨳ�BW�Tj��4a�TIk�K=5vR�(��P�a�D~򌇭%̠ٖ�9�B�"ff �B�x���mi�-�'"��(����e�ўl+Sl\0�{7����A�&NږrE�D������<9�O0(��]1kB���C�Z�K-�,��"hY��"�/O.�"���.
klZq�9�@�T�@uS3�_4�qO��I�����|���i�X��qJL���m�b' �!���âH�'%@�:!�^�F6i���0%��c�O�lAɪ���"�-� M{.�p��'����%�O�D�O6��n/�t	0HþK*��0�� ���NS�	?���vDٺ,c"=n�0q�h�1�W4VT�)Y�m\��#?yfO�2PhZ��"Cǣ	F��y#뗷gv���o�t=�d,J�w�~xybO��hO\�C���0иSȚ�}h��Q�ED�n�F���3�U�G㗥5�摃u��Z �1�d@%>�~���?�i ����3a��-h�ɣ�*����D>�Iy���w~LY���:V��LRg6j�$i��V�'����o��&(�7 �?���H�O09I�d��^(5x�
��t���������DΆ��щB�g(�7�\>�`���G�!��B[V�t����ݫF-�7��XiI�"��{�X�yѠK�џ�HtK�<n�z� �څQB-B����M��%G/>�X�t*z�tB\w7$�=���5��HR���%�*���H>x��Sw�I"�ըP�F�by�N�+d� �(�B�F�����i��MC&�Ad8������m��טz�Qt�K�k��!��b�7D���D1|��02B����5�н'���s�n�	�HONq!��/X��G�γ���h3Q�Hiq�ޔ8:ni����l�Zt�N%�V��L��떰�J	˒�U	aTI��C\�� wO��>�@A�g�R�,��6��<Xd���(zL]�-=q��H��-
�9���L�t�VZ�ͱ��s��. �<�!���*/$�� �+N���Ћ��ż8���Ҹ(I$ ���[�ΰ?��_N��p"��9xƈ���;l��t���I-�<��y��Nd�����_����.�6�0?y�g��@e�q(3[@�(}��,�%��(P&�[x�|��$�A�)R"���?�l��K���
�ص4�L�3��: H�<Z[w�^]�nF�?E��'���bZL-"0����z��=Sէ*�D/mt ly��_�q�LA	���O�,Y9�J�
# ��N�v�P���4k�XxGi��H�צ!<O���MB���#��X�s״42����z^� "p����%��MF�OR��Q&)&,�|��
_�(�<є"%4���+�=H��a�A�ɏ3O�M(u�>}����L�T�x�Y���L��z����V'0;��R���J�$�Z��Pt�<���*W�q�
�oL ������5`U횃r@���'��m:Fg��y	�e�w�4P�b��M>�s�*b��q�φ��$3��O(^���Ak� jp��&,�[�� �b���FGh���eYpo�4��`��L��F���Д�J�Ew�H!��ԟ�a��x��\62.���Qi�AY�]�b���$9
�p�sq.�m�5POOf�8�7�r(J�A��crT�����!�����^�c����r��������<a����2�����<�y�̅/�ܔ��ߚ\�t#�΋I\��o��ɫ�ug��w��y�.GW�5m\"�)�� gHG�@Yz��$�R���u��45����-܉')�k&G+8E� �Qb�*WC�L+P�ߐ	P�k�>O��p1,ڔB����Vi�U�]�$1��D2q9kJ]�	�ڨ�QF�ēTS:�P���&|�B���nFx� Q�4��3~m����-�>"kf��s5
3�x"NΗ{��]O���C)�m5�0���K�"3>���dѿ�2��T� Cy��ج�<0Z��y�҉���P��r�͞��HO���W�
i��Uh�"h��bW���J�i�T�;�%�����Ʈ�O4ȑTLM�C2�;S(Y��?	�B�<	E��8�)��s�����{w�Ŏ{Р9h	',0�*a�`���u
G- `������@���;lk�9�ővC�( �� A�	����4{�Ȱ2`�ަu$�E!���bG	"Y��WH:ړ'�6P����b�@P1w��3`j�yfd�I��ɥGl@�+���6*�41�R�X�'�8t�TFП{�6�C���fO��S%�S�����.ʘ<�27��т%O��!�s�^�"����eB=x���Q32�I?�(�P�1��9��HӌZ� ;jԖ=:DX*���B�%V��aV���	1b�>]��	���|�VJ��y���
&.��^T6m��O��)p3�@/z�D��˛*2��X�P��"�?�@D�"��b�܀���(�������*qv�lZ�[�ցr�B�~�]yF-ޮTE��|p���R�}�
,�tσ"DZ�)n��R����6��x��(@�E�raf�*�F�OZ��C���Z�=	�	4i���J��l�`"'��@�@�Ҙ>y�@F(g���� ��=�ZH"K?�n�3A�,��m�gXصc ®c6<@�B�.X6����H;�λGZ��3�c׉@@$�b��mT��y�A)~��	�L����5o�h�F�Ј1�"�:�'��ȱ��,
y瑞�9C`�8 v�D�4d��{�
�>��]�$ PG��n��U��<�A 5t`)2��y�M4)%VK�b���S���?�R�U4VXhpq�R
2������Ȅ�+M�N]HE�F�<�1�>��N�0\�<�3��l�ȤXa�>3���H�78��R�'���%�ל�� �5�"2�R�����No�e��㊅O��Y�/Z�z���œ���'Ajծ+YqOԫ_w0`�!�2?U��0�@�"�`r +�
��)�W�']���q�IrGH 3X�2}��Ú5;I�h�O1�C.�G�ğ0�I~J�`�7l���2U��=Q��I(1����`� �#�6��`��"s��q��-~N]�'��i�G����5�=<�|a���69��M� �>�����Ɨ0v��=��q�E�ҭ-�$��B��M���n>�Y���չdR0˼��=�	S��y/�?w�L�I�ㅌt�y�]��~b�^�]�d�yD�C-Xh��Ï��hO�a��P)�����G�]It����T�=�e
����T�UO��	Gʄ�m�"}�ǘ��\T��&O�0$�x��>#^^��{�~T�![8�~t�
�/8���F?��b?��E���D�S�Z'I���r�
�?������	�t�ͫW��^|�[�% ���@���iF,H�P��,�VNB�I�l���ӖsC����p�B�#ׄH�^)�����'�� y,.��1hTRb����4d/b@���յ|���EB2Q�x��=a��*�y�HO<+�M;��F;�ْԮR8��ű��ɔ3�l��'m*t���Onў0��䁍.�����+��~�4q �#_����$����ﮖ�{�e��gXc���,��a��ۮ}a2}�Ǔyc���04���"�� �jl{��.]�]��'�t[�K��v��5s����s̄*���_	��Fz�mF�?_�8�G�Ψy�B�ɄEǏ���-=����k/Y2d�$���Q��Ї��,A=���/S6
�J9se��O��J�☑\DN]r���/D2:d��i)T1��؉N����@V�,crY��$T
~h��!̀Iu�q;BcY3>U�DӜN�M�7��1ZK��"�'�ў�	'.��#�Mj�䌸`�<�3@ǻ0b�:�h�\j���p�%�� 2�6A1�.߅v=���gȭ� =�v��6�C+-M�����Q.v�.j��'d�UN˨ڬ�sI�;b�Z��Pc�3�
�EzR�^�N�V� �-�t�5��9��d�f�X��uH^8T��)w*<�Q��cb����qE팿2'�1�a�O��s�	�Q�t�Ƭ�,H�y(T�i�n1�6�<@����OJ0X���'5�8T+n�%��A�4��|!��J)0��);AR����	uŃ:�ўP;�+��J���PUTy9��@��#:Ȩ��";�0�Wj�:^Vq(Cϐ`;R�*�+�?%6�a˓aAv���w����b��~�q�o'�P
�BȨ�g\5g��[�)��T�c�6Ĝ̆ȓ@x���ch<C�^e�O�?%��ȓy��I�������<1��3F"O�XJb)H65hM�����8Lʐ8!"O�eb���H?�L�c���d���"O2��I�!"ƀir�x~<�D"OX�#����ps�Ż/]�p�"O�	[Ҁ܀t�(��#OM�T��p"OL��'�C*�.0c��S u��"OHa�P��,6\����K.\J)u"O��2�E�lH�P�g�!����a"O� d���W�m�"��tD�*@Vd�v"O�]�-^GY�IcaCT%	.���"O�|r%	Ț�,�����'4��*�"O
����K05����w�M�0ꎔx"O��CB&�rK'��9q˜IE"O�w�J2cdۥ*�- �8}�g"O�}:u��ҍ�шMv���I�"O�5�DC6d*�ᵦC>����C"O�=���7����E��J�D��"Ob��� .K����N�i��%"OLĉ�)��$��S������@"O� �� @�#'� ����;h� ��"O��!�-���5�w��)J\�3V"O�P#b�P�Mh�"֤pC>i�7"O
�J�$FQ����?@P�b"OX��ᩇ(!K$I��h�NQ��ʶ"O�h[�@τ|`���F'��"Oh��F��>x�F@�-���b"ObH(��M1N$pQ9B�Q�Sf�m"O�U���'�d�C��08c2< C"OP���㏂9*��QV���S\�a"O�x�KF0nQ�#d��m���`%"O�U�2�B�S� r���]��tY0*O�a;�C,25"� �R/K�P��'�t8q �1r��E���<�k�'��Ѻ4B�?C*��׮ה!ަe��'@(��GS�@H  -w���'/P���nX<s��y��I��+̲ ��'�� @�l�,Z-�A�,�%r �I��'��+����\��ƃʿx�<��'�R���3��36(�?=~����'A���śS�V�����;��M�'6f�Aj�m������\�<��
�'��$rt��Y���z��UY/�
�'5�y�t)Gd8���,��J��1
�'�$U���@�W0�!X�G1O-h���''����JR�a��?���'�x��1�ܘ8HU����1'�J�'/Δ�W
�> �� �&!6���'O���3Ȕ�-��\Y�p�a1�'�L����i���!�ԪqG����'�q�i�J��Y��)��khv�K�'_6q�D`��@����Z�a�&	��'��5g�Kl׼�լA�X�:k�'�0�JC��5?][��^�T�ntS�'�X�� 1�d�`]}� 8�'��I��a��M��!����B�����'Lݲ��5\H@���x�	�'��q#�*�	.SLQ	�ʚ�̔��'���I&ϋ�+�R�Z2��#�����y�!�)@����ǳ'�f��B�y�L?]Y�}q��9W5�u �B��y��p*5����*b�]��D*�y򮀇7�Ա�v��[H�PD�W/�y��,]�̳I�#*����僶�yb���$��oIU3nE��-	)�yDG7h�p�bALI�����7�ت�yB��%<��ِb�Dj4x{���y�*��E>X�J�ˎ�vo���% W��y��� ��ecU�v�3�.��y��S'l�Ա�R��o`%Z����y�*E9^�JL����5x6$pjĬJ��y��!�,Y��^؜(�f@F��y�HY�[����E�?� �
KZ�y
� pE���5UH�)IE��:��દ"O`up���M�	ʒ(Č8�t�X�"OZPB$��.��0���L�9���)�"O��	���, �y��#&���@"O��Q�^�,�nE��NQ�~��A�"O�HSU��/L�Pt�4gܶ5��=h�"O��2��u��Y�4��p[�"O�ń�o�N9!��� g��\Z2"O��FL	�}��%�5�rϔ���"O���À١^ټ����U�Rq"O�Xpe��\�! A��X�6��"Os���%X�vQH���zo��s�"O�H�q.�䪅F�cA����"O�m�!A�%97KQ:+4f�B����yrȒ�$m��o�ʆ��VC��"�!��bS��;��	��~�iUc_�g,!�� �q��f@IIX���AF�2?!�DW�7�h����'WʄY��L�b�!�$��Yͦ=�r-IV�ع���65�!��O�%{��W���-7����b�!�䌢Q㲭� �W�, ��fHG�~ !��(AhM�u�.T���� � lM!�D2\[��
D�!�W&Ǡ%�!��&�@	���V20IP�*+!�$��s� )��%��M t���!�䊲����!�S�y.A��X��'}2�A��@ >����dk��~O�0	�'�;Ձ�:L�^�
���'R>] t��=�dh��/{��!��'ݐ����n!v�,�<قi��'~�P�r�0)�h�e쏞 �@��'֌{wkW�ĥ�̇q���'/��N��PؽB��-X��
�'9
� �h�ݦ���JB+fg�0��'xF(�aۥ&��M{r�ǩ^"�ի�����[�Z��Q�R:d��:��b�!�D��rWH���:��
@:3�!�Ѵ!�xu3�E�'0\�!#F��5�!��� �rx�`
�)<<�ppF�R��!�$���A�0�0-P��b�OU!��ĴgR��(� J�d.l��W���!�D�&����ܣ�P�2c�A�!��V�l����"�]��(�V$�.o�!�D�;�)�W#<�F�d��!�X�(8H8[3o�y���,м{!�$V*��c�$�!a��fl�=6\!�C�y�$��aV�RE��#���*!�$�-SI��F�'���ɐ`H�U�!�d�/'\h|���V�e��L�����,�!���[����l�!��5ߜt�!�$��(�8���"� f�T]�˓�.l!�^/���$�cq|MӰ��!�$?2�~�˗�mC��$�ف!�!�/|f���i��HFx����ӽ,!���q���P�W�\+�`zT�MN�!��ΐ3_А�rGN=��e��I��=E��']�ٹ�#��7� a蓬��,z�'��2O�y�E2��A�|���
�'�rЈ HG�T���!ɜ�
%��1
�'{><��-� ����z��\�	�'�8R!ǘ�/X��I���A���a	�',��:��

5�qC���u���'y����S#V��Wa�%wf����'����j@�\\{F�_�l������� 聑�O�C���*��"��L!"OD��"?h�j�Yj��~�`�˂"O��	��I�#KJ�6��QQ�)�D"O��Vd̅MWA�W�=^P '�'#�I4!�&T(.M��H{�m��?��B�ɛI�\���%���x@Fl;]*B�	`tX���F8+���I��J#�C�I3Fg�2G������`-[�%<�C�	$XH`�Y���z��\r�l�OB䉯������Se�"����Vf|B�	�k�ް�0� :(�`Ã��!�\B�*_V�ݲ���5u���#��W3.B䉉.O,�w�C),_2��T'�-Q��C䉥�XQV�EҰ"&�ЮoT&B�I�p� )Q����tV �`0B�ɺ^D�)8�a��a���AFcO/��B��/xSb�[(]?�j�����)ÞB�I� _(1�Eϲ^��`�H�"[d�B�I�r�d�Z�-E����R�]p�B�	�G����Q�â_S�y�n�9PxvB�I=K�3{Zps"e^7�ġhF"O
)��A�3]�� ��)U�#n�)�V"O$1B��&9���V��?��ɩ�"O��( m�3銘�cI�/<~�M:F"O�T�� XP���'�8i�0i"OTmJV+Q�]0@+�F��\P�P�"Ov""�P&H�mi�E�>8>�@�4�'���� u܆��RNֻt_~DQQd�n^!�Dt�f�"*NA�y�HȤl\Q��G{*��DXp��'�0�c�b@�Wh>A�"O�X��&p����b�*Z����"O�<zS�Hp�ERb��){�0��"O���p�H�F��tfS:��U$"O4�2'�I�V��(QeA �D��R"O��#Ro��V��$�Y�L��yR�N�
렅��GF�BMV��Heb���S��?!�ՈD�����"��9Z�xҐ@l�<�R!Xb6 	���>	���K���@�<�/�.Y���X�� �J$<�����~�<���p���K^
c�P�� �]F�<Q��؁̈���Åˬ\�q)�v�<��M�s)�%ʡ�7��Q��Ny�<YA �09ֲqJ`&�+���2se�t�<)��XB�T��@#H�j����n�<�4�-��P �IM
��4DZh�<��P�j���#���t|�B�c�<y0J�!Xk"��S�ʚ�HztH�_�<���L$\����Ôi(��o R�<��N�"J��, ���`:�Eb�<��NΪ=�J-�!��]6�l��]�<��HA�t~m�G�H��BօY�<��M�ӂ�1P���pbp$�@��Q�<���+P2|���@�ja:�
J�<Y��5$��HI\��B���E�<�w�Y�l0*@�٭`P�A����Z�<qU�ذD^��i\0Iiꈛ�C	W�<Y���N���35�,0�=�/V�<�-݇B��X@��#�&�BDJ�<��K�ni�{��Y=SO��Q
m�<q!+W-d�85���;n5:��Q�<)�?�����eD��!�h�<a�D�<4K����Hzp=zqi�~�<���<��� ��=N�����K|�<A�.�<S1��H����u�q�o�<� ű��Ű���g/T�Y��J1"O���a�6c��Ԯ�/X �ȃ"O����(OZ� ��C 
˱"O2�apɓ�2�p1X.��l���pf"OB1!�6���b��ߕ�@}��"O�cE�A7���`��ѳL����"O�ѣ@@'GK���,��V~H�
�"Oƹs�<e�@0p�ߠg�uz%"O����j�p�R��N�n�Z�+ "O�̘��3lk�	��ǣ1ml=0u"O�}K���	�.8�F�yW҉p�"O���P�A0��8��ȏ���Q�"O���1��IL��+��4��$:�"O�m������%3�'Q���S�"Ofd9w%�4h�\bq�_�c����y菙m}l�#C@.4�����5�y��J7?��\P��<)M�ðJ�y2�P(,�@ȓJS�-�tʆ-��y�M�&��F�B�8�ԣW�P�y�b̀,+��a�;6�(b�@L'�yri����|����<_*�DÐ�	�y�%�c����\�P����`�L��y�-	�$c��)E�l�CP떴�y��J�y?�t�4�M�?}t�kXq��B�	a޲=���صb���K��R`�B�'�U�4d@���ЀNX�

���q1��4hS<%y�i'[D���'��وFR�s�F�����K(���'k���pB����)� �O\2��ȓxve��%� h>�����;m�~�ȓc�F�(�M����҅
�ird�ȓ7�HH2O�2h�2ς;%L !�ȓ9!rI�RB�?3n����	��z5@̆ȓ�j�C ��_  %S¨
.p�����o���Q��FRR��t@*L9Շ�/��	��P�q�^�$K�'�TQ�ȓk|��2��y�'Ŗ&-�jنȓ,�h����|(c��E�p�r5��E�Tx�d�jHj,`s/��rI>��gU���W��fWH̓R�׺L�(a���p!1�̏GU�eCP��W��\��~��H  �I�4m�d�X�T� ,�ȓ}���`b��&	IB8a� �.?���ȓ_�ޤZǍ��U�t�Ȯ2�X�ȓN,e:U��f��@���ݫ����ȓ0H�-jE�\/L��D3w%E+v�v��ȓr����Q]N�M"f"R(���ȓ~pĸ�2iё/@�Y҈�'d.��ȓ9�ix4�	N��Yh&Aܹ��ȓ1O(��ǿ�6]UL����p��u�fI�<��4�Ꮇ:1�4�ȓ�X������W�V��j�!5�<�ȓd���q�ٱZ�ܣ��G�f�ޅ��r+.�8�� mRH�S�̌<,��l�ȓ�qa���\�ˀ2@�.���}��&��/��]ǗO��P�ȓIIY��Kl=e�4�G�����ȓ9VLYa�,�	&�vi��M�8���?�T<ID���[J��Y�7/����ȓE�\(%�U�\��S`@G����l�p	����K�X���"��{D���. t 7X%	����ም��(�ȓ'l�$��˟d~"�A������>:uZ厔 sF�y�W/�$���S�? �����.;�	��T%�pٔ"O���`D� R@T�D,Z��>�� "OH���*���h��Uʗ>2e�혂"O��YEN��&�aҰɍ�:Fb�p"O��i�%u��4��BD� ��2�"O��:�cK"0F #DoR @��(�"Ox��%)՘)�쑒0.�q�֠�"Otҷ&S2n���Ox*�y0"ON��k�6Z|��1�#� a 0``�"O���̛V6�m3��G��t�2"O��䎔�+���ghˋ'0&Q�"O�5Ώ�[�D=c%��&oN�Q $"O��{6O�,0|�I��� � �a��"Oجjd�M�9!^=�%D�#8d�Kr"OB*�)�A��%P�i��"O�)y6�V�4��!��&?=6��"O(��i|t�����B� n!��"O�4q����L� E2��Q���"Ob9��BC�J1�ܱ���:1Nt="�"Op� `=ig�M?���u"O)�U���}j�p�Ϙ�l��1�"O��HBu���G�
o���I�"ORU���V�=F8�1r���]��h"O�+�4g߸qk��ҨW�R\��"O�AB��"kt�aؗ1��T��"O��S�13+��)VbA�f�V�1v"O���%EY��銃g
�o�(h�"O\����N��Y�h�I�^ػ�"O&( &Iė>��)�1M�z[
%��"O��m\�úՑ�Eǧ\�t�C"OfT�bh	�(2�K��a��C"Oh��k![H�D����!I�F�ɵ"O�a��U�"�F��V��)NNP��"Oi�0��$T�vp9��:~��"O@�"� 	m�e1M� (�p�8Q"O�pHE��P�j��6k��2���"�"O���bfӖ`1 A%O�{�	�Q"O���""��|u��EE�P
VYB�"O���.iڽ�u!�
mRl���"O�e�F[LR�Y�a�-[4V�KW"O�|��Ѣ7�8����j:��"OFm�e��;�Y��n����"O�R���f$`�M��,��m�u"OjȈRj�(�J��
� ?�� X"O$R!��:0�@I�5��}���d"O�=(@(�ö�؂�L3D���P�"O
��A �p0�AD�Tl�Q"O�ġ���gӄ��4o��� "O\�C�͉yo��3�\.ef#"O���Ҥd�(`Sr	�m*v���"O`�V�ި:��c�ܶ$*n�+�"O.ru���F<L�3��5^"����"O����G	�~5�mf��,e�"Ovy
X3z�XAd��<%5|@p"O@�f ^�G�<h�@eQ�:�I��"O�q�DhD?qV��P�Μ�9��u"O�t��]ZL1�w�U����"O>�0A���oD�R�ϖ5�85�"O�!9C��?�(��R/8Ѐ�8�"O^d�D�Վy�Bt!��NQY�܀"Oj�R7��# �(��e�B�gC�8"�"O:��Q�ډQIwk�>zQ	S"O���4.U.2J�����ɘ�P�"O�Q2�����;�k�*W �A�"O� ��*"CڦX�����#E0ȡ�"OlT�Q�Œ9� �Q
rN~��F"O,��`CH2r�lpR`��f�2�"OFX3B�Կ1��ɦ�����[7"On!PT�Z{^-H��,pVR,S2"O�`p3霪\�D�I0�Q7_5��"O�D��)SS�����/-40JF"O,�R���3����B�Q�H��ᛓ"O�t!&�ϳ�a`��r��Ys�"OV�Z��@�,�q��aE�p^ @�4"O�	��޹�NԠw+��-�Y
�"O�8���7�@���H_$BQ�"O���e
 �-%o㤡jr�(�!�هk޹��"Z&cx��q�u�!�D��
 ��M�:~��bv�߄l"!�$���@�2!S5~ݾ3��0�!�V��`���m�%k5k	=>!��7k��܂@*��-��uIG�V*!�و!�!iBf��`�Eʞ�!�$Y15H1bR�R�9�i5CQ�!�$F�@J�p�6�ĕa������+r�!��3��T�7@�7ik�|Z�猹3�!���Uq�0nK*HN��X6I�C�!�d,mP2�aH+ y�A� A�!���{xJ�����2�i��*\/!�	p�� ���g�~���썻^t!�$^+	g�!�4G�dj�T��]�*]!�B�]|9�Pk��C�ՎH7!�d;�D�SDK/SV��HS�89!���4'{8J��^:,��#�!��_�Bɞ����Y7FPU�fb�+	!�䈬5�⵩uEԇqP��
�����!���.f���f��TJ�y�bM�|�!�D��>�^-�D�&3IVԀ�N٣b�!�z�8��%B�!�$�@���zV!�*�xY��GZ�_���B.\|E!�dKr���#�k�*MsH�D�9V-!�C>��h�͖�OeP`�Te�*!�d�1�zy��g��v����֛y!���44��
Hr2�)3C7of!�$ކ K�5[�CA�zt����"W5#`!��P"�Ì*hƬ��q�M�fD!�ĕ<Z{��G��[�T�dM�XI!�D)��0"��/�0�
4j�� !�$�)od^�i� ��mȅ�ʕ!�T :�B�iÊ���<��ۣ0!�D�!lC�ܛg�G�T͐��6�!�d%����S'ߛ� I	���H!�d�L7�`��m� � P{c�!S!�$��}d�a�фۥz�����D(�!���#!���/,n����#?|!�ӫ^�xMq�\�@V|m�F�3v{!�ă�)d"�%!�UMT+s�Ė#E!�$ژ[1�X"�Z\H%�q�M�?!��1�P�S�Q�=0��QuڥL!�ě�����k�d ����,�p!��Ôo$��0��".� !�P[�"OP�:'#I�6s�lY����  �L��"O`�j���������F�9,�"O&L�7eΥ)�%�P��=�JY��"O����\�>���mZ�.r�i*p"O��p�k.<$)��B�~S֨�v"O�pjD�ص8�J��1��h��\�4"O�=����hj|�8A�/���`"O� �ȉ�I�J����
�L.�X�&"O�`ĪA�%&�y�6G�M��*6"Oz���Ӎ8�*`��U�9�"OZhQ�'I�����䎘5��u��"O�C��?TR�Y��]W�ˤ"O��a	<
���!�4=8A"O�+����f��M�a`�1 �E��"O�Ĉ����AP��S@FWA i��"O��T��Px���N"O)��y�"O:���+P����X����"O@=��J#j��-��O�~Dkg"Oj�Q�`ãDm ̳q�5�Ι��"O������^|*582d�d����"On�rA.��Kø����ߟ.���S�"O �0eNF�.��hP��sw:�3"OF@+2L���A�Ƀ4@R ""Oօ�#�U1]�� CbI�F�d\�"O�	�	�&�^T����u�i�"OP�Ar�P��ⴘ�CK�&q>m�"Ox)�e#�Rȸ@�R�[�~���"O̤�P�2V�a�T�E�Jl�ۄ"ON	:/�6 J�����
�O��c"OJ x���7)�&����|��ɋ&"Oj�(�,+Y����*����XG"O�@sb�ۨJZ�{R�=&�,QE"OHQg*8LH1�g���ق�"OL	�'�L�>�����"Wܚ��"O�#'��v�p�DG�'/����"ON�+2Y��9UϠ	(|��"Oh�i�A�5���)���$n�ű"O�%�Q��1���`U2)+��@"O��ڥ�%W�̣�,E�zo�h�!"OD�j�N�f�(}a�KI%�2�Q�"O���'��rߺ��KۋN���z1"O�l�(A/=zĀ��O+���S�"O�9�6N�H�\-BQ�Z0}����"O(�"���/T�����96�j��"O𡅫�^ʤ��-�1� � �"O�����Âu>P�Tl���XZ"Oh�����
)� Ѣl�# ��ٺ0"O�SG�B;\x�ӑ��Q����r"O�����	������|d�b"OH��]�@W�ISH'o�4j�"O�E"���L�i�F'�d�]�"O�<Ӳ�I?�Z��ǧ�52�c"O d���
^�Q�2F�
eٶb�"OR��*_�;�������/F%޷�"Ov����̠E����U�M�Cl�cr"On��'o�
�򡒷�[I����"O�AbI1X^Pc��@�����6B!���=�ڼif��`el2k� �!�Ěaݾ��tf�0Jܸ[���A�!��Æe�XB��pDD�X�ƙ�!򄅎E|p�)�'
�U�|�[��7a|!��QP�x��ϕX�8)��3t!򄌮wI,�`�
G�*���wU!�O���ТE�l= �!W�� |!�$ޘ0�̡rTI�}�E`� w�!�D4����G!�HAE�R*!�!�d[��f4��O�l
N1s�-��!򤁟zFZf-6o&�m��mA�{�!�D�{��r��E;2zұ��B@�V�!��޻m�
]sH����M�H�=}Z!���s�fx�h���y�&ʉ�!�� ���w�I.:��1rEn\�,]BIcV"Oh� �CA�����V3"x@ ��"O�|�e@�5T5{��$ma��"O��  A��V�"9��%��$UzE��"O�P������0�EF/5�MPv"O�Pj�B�!��Tqc�@/�h�a"O�H��ǆ2oV��UkE�w i��"O����#�gs�[���2�� �G"O�I����� ��KӃw͢ـ�"O�Ё
�Z�2�i���h��)�yRI�D���B�hJ�q��0f�.�y���hstm$�J�ezN4"��F=�y��.��B'Q�[���Jɶ�yR �%Pl D�@O#Z��$;En]'�yB*��~�� �o�c�E���y2����\@���[dp� ���y�P�8��!��
M�T����y�/��Z��Sܮ|z|�!�H���y"�;t`z!�p燴z�)q��-�y2*\6�V���ND�a"���y�K�k}�Z��̶?�nY2�N 9�y��ґAM��Bg��==�p��Ӥ�y�@��~�|i�nG�2d�		#�K��y2�l�	Z4�N$�
�b��y"��6��\ʓ@�&Lt�@{B 2�y�*�SټIJ�#Zp�����y˞0�@}���T �JE��L]��yr^�_�Ҕ §|��Q��N��y��C��d�s ��� ��y�(-z��(C�c>�jefk9�y"����b��q� �xEB�I	�|Z��ŭ��sɊ2B�I�F��a�� �0@&�yw�
?!�B��.0"9��(K�d��p��%�0B�	�J�u��	t�!�!�H�&�^B䉼U�ܬ@�,�,,8�	`��۸r�@B�I�B�*,A�
|�:=����2%�C�Ic~.xAg�? nMxg��)�C䉐tS�5��O)<;�-b��	;`��C�	& � �r�d�<S�p#�(�0&C�	=D����L�xTR���8|�C�I<9��Ը��n��)�����B�Ƀx�<���%Az�]C	�� B�I9E0�����U�|M	�'O�E��C�	">��*�F�0��Z�bM�U`B�	;��Y0�KU�h�4�M�;Gu4B�'1�ppC��6����"E��C�I?#2q�G�q��0ѡk��85�C�	�<�H�S-6��`q�Iں;\C�I.it�\�
��4隐�ׯV�b
0C�	�:�
�B�@)��dI�HS�nu�B�I�?B�5Xw*�͆p�dE�� C䉩�Ҽ��I��f�X��tぉ*�C��eJU[&*\�3:����� C�	�d�YzՄ�LT��z7%ކd �B�I ��)KG��1Fb������x�B䉧Cp���d	��^I�hdዟ#�<C䉖	��G��� =b�3@�N4:kC��%J
������Ql(Ҫͣ[�B�1x��ӥa\@)Б�̍_?tC䉽K�&}�CI��8�0�d�;V�B�I�:,�Sd��A�_k]�B�	:_(|5)'���Ns8���D����B�I58	fE�b�@��j�%+Z!�� fd��L��kV$�2ů��}�Tઑ"OR5��� 	�������.�*���"O�C!�U%L�b��[�L���"OZ�p�f��P~��c�C�e���"O�h0�'l����Շ"֌�A�"Ov��A҂w���$��>�ʙ�p"OH�U�\���� �{v�L��"O<�@C�ɲGy2��C<$i:���"O&Xx�-8F����J({I���"O�](�ˢ  ��.��/@5��'�p$��ʀy/�Q�6$$o��0	�'lf���g_��X�F�s.��p�'�f���Um�l�u�R�t�V���'����G��&��Zl��b��X�yB���¥Y�j�8NX������y&��<����%�"ȢHR�=�ybbK�9
��f	�*}��`1g���yb�@�0�p��'l����1c)�y�FY�F���j��^B�	�4`���y2X�Gr���mB/G��)GO��yr�ыB%�g	AC��p	I�=�yR�?d�������.$��ޜ�y�ȱu��@�!�� �t��%A��y��*�"�`MҗG� i+��y���oHxb�Pd�x����y���GWf@�e���2�K�*�%�yb j~�|�Ӌ�>/�� ���y2��F#�@s'=zȱ��+�yR�=�@�
��93���!����y�k�)cK:�k��0=j���fƐ�y�E�rF&t��H�2f�@ ��T��y�!BG�a4��x�y�qn�-�y"A2~��p�4|Svu��l	��yr*ȵ8��0Ud�y{Ƽ�V���y�/�4E����&ő>io�kCmQ�yR&�!ƒE�����5 	)#戎�y���%��� m�
.����.���y��[�F�*|:$o��w�Fx�u���y�%٨ht�@��f'`]�1�љ�y�k��dc2����ՙX:�\R1� �yBB��T,�˗/K$�2Y��^��y�2mZ��w�V�|(3���y�,�1׺�20�Z("<)�".O
�y2��3h�|Z�	�=E&�q���yBf�0��ؐ���L��Ue�'�y��V�f��l��=t�%�T(ɩ�ybC�2N���w��z������y�
6�r��J׷3�=AT���y�NLz����9}�ڬ�F��y�l�&���
a(�?BC����V��y2!E%q�@�Ɉ6:|X�B�R�ybޅ(� @���axD)���yr��0w��,`@�k�sfe�.�y�`�8��x��ۍ^yc���y2�� 4}"j"��\3~�!c�H�y2��vJ������BB,�x�	�'z�)���S�!`P�c "a��]y�'���;����8�>q��oa���'��h(B.��Hԑ��DC�V����'���#MFJ� �n�N����'� KA�D������ȹw�$�	�'.�ʔ#ߏ`JX@QDQ%n;(P��'�H@� i��:q� �h7���	�'Xܨ���/� @ڀ�D8h:�	��� La���^506���/�I.��"O��B��mh���D>E$c"OR��U  mQ
y�f��KZ���&"O4�� ��s���W7_I�Q"OV���'i�ܻ�-�a<��� "O�\8h��+�:X�抸k/���"O�l	�,�5��ٶ��!A�*QQ"O��c�߄e��S��W��QZ�"O�I�Vh�F4]0�y����"O�50��Q�px ${�#�+��ڲ"O8a �)̂W%��Y�o��^���d"O<S��$>�ı���zU�U"O��Q�"K����TN�U��p�"O��@�	جg���������ӕ"O�B�oמ,� �Ke�H
�<��%"OFPS�^�\��-ɕ�ښ|q��g"O���r����v֌� 5Wi�"OdD�Vǚ:Y�E1'"T--���"O:��P,Q�0�8CD����R���"O��b��v1
��.¦&ꉀv"O�yJ΢.���qOOI��͸"O�	��� �Z�heX����l0���6"O*��M�=�v�8!K��~*���q"O�����0��I���=�r�a�"OX��Y(�#�]8t��7W!�d!<{l]eKE�
�q�ϻl;!�U�ʨ��59�\ipʌ�,�!��E�|�ڑRqa�+���H6���CS!�DLoOܰ`�E48���H:W;!��yH��	�%	"3�d�A�ط5 !���q�b(��i(��1b�n!���P�ĉ�A�J����Фlg!�$Z�*/�tcցG=>�D qU��,!�� 3��Sq-��h�(Pì- !�D��7�dd�D%�?oV �E�R�`E!�d3<O@Ip0ß�<l*<!�J��h[!�N�x�p��k�"'-�j����*F!�d�75�t)���w��`xUF)x!�$H,^+l�t�[(Q���hD[�!��gY`ኖg��|�.`�"�(A�!�dنBV^!�g-�>���A�L�t�!�DH�z���z�# �)Ҁ±�!s�!��=uP��ZW�,r ��n�g�!�dW�s\u�����DZ`�{F��1!G!�F+�ڤ#P藨|2I��J�hB!��t?�p��`A/J���D�P(yR!�$WY���d ~B(Fk�>A!��Th� @�$�!2<)��i�:=!�D%'L(Tq6�����1.��L�!�ċ@�2���!@�>�`�5�'�!���Ťyo�6\֬Q�v]5�!�d bZre��-� �.��#j�3`|!�ՙQ�Tm��@E�_��x���Ӷz?!�D?(D���e�Ծ_�,0QY	6!�$�>Z�U�0M[&��/�!��S3�� �A҂'�&qK����!�!�Đ
~�s @י&�4���-q!�G/7� ���� ������6r!�$�ϰ�c�/�!o�ਠ�W:�!��?s�jx�F� �p1�Zn!�ċw�(�!'�<j�D�@��!��ڍz*0	����80���]"!�Ę)�Ji�g��c�.	���
{!�B'�t@�EAܿ6��@�&aX�Ss!�� R�@��,m�Ć(&���"O�S�GK; Ub�����.�
��"OX��6)G�
hu(���H��4�G"O�T����Bu��r�AY��T"OQ���<W�t5���i��G"O��×D1rڊ⇬�.��qR�"Ov�Z��ٞ�0��1.,V�v���"O1a�_C9�+c�O�NYr,�"O�]��$����,M�D�&!�y���Bi�A�FX!A0m�F���y"��.�1��G %w�����J��y��0v'$*E��x�;F�E��y`P�zkt5s�NS��l@u��>�y��}E 8���H*UzL³h@��ybk���%��fo��*�(%�yr%N�p�x$����d��S2d،�yRb�R�0[�VA AL�:�y�� V�l�eɐB�Zĺa�S��yRΚ�4F �5
I� ��y�M�Vc��#�צT(�0��,�y�=/:�d���TT��E��y"�t��8�Ί�(�h k�(/�y�˅A$��d�Z�$�`�SBn	�y�ʂ�8�Ru����l�4B��y��<wp|j�+�SL0g��y��G���Y��摜w�$��eO�yb-E}��@жjZ��Mk�(S��y"��#~�&g��j)ھ�y2��;nE�O	�O^h)	����yb�{Ԓ�8�]SP�
%��y�l�+j�c&��b�@��?�yҭ��gf�UR���\��ď��yr`ӛas�0�%O�D}�Atl�y�BH�`�X5s�CO'C ~������yr�Ѱ ��XKƪڤ-�~�����y��Qp�<Т5۔O��y3R��y�i�1��&��7K�n�1�΂�yҊ��_�Z� q$*L�� � _�y�
��eJ}�D�	5�4q���yrmY=&�@��|QL-�N��y⣑�I�aA֤�+p�&�F�y"�ϓ>=X�R n]�lv��J���y�_��|	�W���_d�&/�,�y�N�=F�(@�D��W�z�����5�y�I�v&�-��MصL��lz��֕�y�l�ԡ�D)CȊ؊Tʓ��yZ�6���U�ԗ8�&���ω��yR �s��J�C�4�<�:�F� �yr&��0bX��Y�3�*���M��yB�A�6���x�䎀'm�
p�?�yR @5O�v����L�1�ҁJ  N��y��3Zi�%
�������穛�y"f��(�l�cMЍ`��[��	��y�)�=�E�fl�#4��3��_<�yBe�1 ���蕁��l�����y2�;�x�Ta�"*6������y�i?)L4��N�ÈU!�"�y�C��\�3QDԕzb�a�Q
޸�yB�K��M��Bw��D���E�y�Ē�~�	!�$Ń]ޜDR�n]��y��!T��w̙"�9qw�P�y,��Z|�P��� �J̙�cʭ�y��ߢ\�FЈ��0	)� �����y�jՔ V�hy��v�\ՓTG�!�y
� ~�-H�a!�Y�LK B�xxi�"O�A{`K����ED�Tp����"O�а��ǭ7�h!`�/lQ���6"O��
�Um���7O9V9�M:�"O�a�aeǽ:&��#E.#j�"O�� bB�D��=���5"O45�m��@�Rm�%�dv�m� "O��� XH�tP�-_�_S
QyC"O@er ��2$bz���.ы4(h�"O��!�K%�(!.�6F2��hD"O���ud^�6[���mA�Q%%Y�"O��ʁ�Z����P�I�5l !�"O��	5e�(���&#y�Ei"O��8T)Y8��ݻn��p�"O*�¡���u�&����M�Xk�"O,袦�B>q�U+!^�w+��:�"O~�����?M| ٲ�ʌ��:"O�!����(D��(=n��C�"O6��pNV i#��'�d�8�"O�$�7i͊:��a���	�TU��3�"ON8Ig`��BV��A+P�4U�"OR���ȝv7����o=k�R�"O�`��� �l|#q/tG�D�#"OА���[=��i��^0l2�y�W"O�%�G`H�Q�mʆh6�&�ӥ"OZ���@_UyQG�#[��b"Oj�3A�ɫ����s�O�wV�Y��"OZ�Z��K�ɒG��4Jڶi�D"O��Pd��;3"h=��Éu_4�[�*Ox)Ӳ�˖sv�%�V+FN��'������LVU�$��qk�5�	�'d.�8�KS�Pf|1���-i `���'p>��#B�	R�P1e(�q"H��'{T���I�2��4�:i��A�2�)��A�$Xnn%�'ߤ5�8,��4�y��ƠW',d8��:��q�e҄�y�]�K�00R��_�z+�u�4EJ��y2N��Z�x`��wu`�xT����y�mN�6ܵ!qL�i�@MK$ƕ��y�LS��n�Xfh�*m}(��S���yB!�&).�B�$ܚx����0��'0ў�O� ��C�w!�|���[86�.I�'�<iy�K�-M�"�r6#�([���'s>�c�h���D�B�1e�5��'.v�14��g�ř�Nێ
��$A�'�$��L��B�����kʿ9Dm�'P�a�4M��cИ�I@�*�s	�'�dАM�D*�I�v��V�j��	�'��= e�� o�1�c��T���i�'s|
�j�0��1�EaU�#R�`	�'h~�Bp�A�8Y��L������'�\�ńs���i]!����Y�<A��ήѺA� �;g�m�Q�Q�<�e)#�[�e  nvTU��P�<��쀲06@��'�VʄH�-�K�<�3�Z#l���{#ʛ�z�&����J�<����%�
�y���0:��+�bYJ�<�`�L:3T�����)�:�!�'�0�y�I��P���Qʍ��Д�G�N��y���<"�2d�gʔ��9qv�8�yB�5�����_�5�P��Z1�y� G�1�RgDN�A�"����\��y�E#'�q�����A,�@�e��y"!��~���:C��5��PUΆ$�y
� ޕ�!��"#�e�u�E���f"Ol���KV�PN%��B�dV�"Oޱ�">R@03LP�\x`""O|�d"��;�%k�H��-��P�"O�ذ�S�r~\][���nk"���"O@<��e�.GK�ܡr�O���"O$���T_�v����=� 	{�"OJ�(�*�.o\�M�0F�ƀۢ"O�1ibgِm6�5:�mH/B��t�D"O𘒳�Ƃ=~V��k�,k�"Y٦"OpѠc�LH;d�����qw�� �"O�X����t�T�qW	ܗ^k��5�'-���>"��`
���(��ʖ.d�C��.tQX��v/A�i�ʄ�FG
?g�C�	0)g������Wn� �B3^�VB�I�{gb�#&̝0�^X:si�k9tC�I'gƽR�*ߣ4}�-K�	<wv
B�83�֍�G+ƃ
^x=�����X6.C�I;�� ��уg1���a�I�s�B�	"fQ0h�s�P�;��a ጟ[�B�ɯI� l[����25h�����t��U�E��#6O�,����bG&s!��C|�@����I#=�J +�oP6S�!�$ț<̈ɀ�ܗV|Z\pp�ܷs;!���"9� `�kT?��`
g%8!�dZ���.K��8��lA�p4!�P�}S*)xQ�T�P�w��&!��F��<X��˛Y]<����ϲ2!�D�T#:��A��oAm���!��\k)� %�ȇ.��%y���	8!�۰2����!O�#�J�`�a:yJ!�$_�x@*�;42�����O&4J!�$��&��q���33!�s��P a"O8�W��>zئI��u��l"O�c��ܲ&d��'`H�iVV��f"O<�4��3)e��/՛IM�}+w"OXA����2j'�u�Vn�aB��iU"O��JUm&tflL�b�ԌF^,1�"O�M��B*L�z�N�A��"O����P��[��ty��)�V<!�Dʉ?�����֛r=h��bjE!�dH+�©��@D�0;�qٟ?+!��S����(W�M.�YHe�]n!�,3���d'�E�D�H&��h!����y�,
�?�����*NT!�D�@���Za�Mv�L�I�^!�DP��P5�$&�-M�yf.�
�!�$�w��qZE�Z�!�H5���Ī2-!�$9��iP`�\�V��%��F	!�$R�!I�xPe(R�,�"�dC�6 !���Y'�	�5k_>z� 䁓C�7p�!�Ē� ���*K�Ll���F�o!�d���h�G�Q�sN� Q�Ϝ�U�!�2�r�16�Ɍ7�2��um!��F�8�@��&*M��f%3k!��)4�\!���n�|	��9dN!���,T�봤XOqᚳ�ْW<!�Dۜvˬl�g��0I"��	�71!��9QV�����#�"�!ȏ0]E!�� �������;�<�b��7P!��ɔv���'�2`��å��\!�d��%򞔠�� 2&�Q��Ǒv<!��4�<k��mƠ�Ғ�ȧ{&!�d^ }��!Ô�B�5�ҝ���0#!�� ��s ��W��h����W{ޅ�"O��A3��0�^����Edy�ݸT"O�C�̌V405�ȥ��{&"O����e�[���E��K���S�"O���uOM�w�Y*#��]��DS�"Ohѱ$2��Ђ$���&��h'"O�PQ��f�0B&�=`��6"Ota)���j���� ą�H�rv"O�ڢɍ8	E|�E�Jqh�f"O:����H�k�b)	e;��c"O�H��j�H����"�/$�"e�"Ot��--O�qR�
fI���ϝ�y"��p�xl��_rX!�v����yb$Q),&�4�J�U�@�&���y"h�9h��IY�,]�S�
�{�����y� #<2lH���uP`�$	�ye�:q2�����$b��`	$�F��yR��'*��Q O?U�1�_��y2�Բ	�>�EC  VDءx�;�y�H�!3�x\��Z�m�(Jí��yjM9wC�5�BW�r�y�R��>�yr��%@��X� OS�����r�A��y���:wn��s�k�"z�.髲�U��yRg�<@��Ip'�xz0	[G�Y��ybD�L��G�,	�ժ�ǵ�y�H=�.р�i�w�6��eL��y��X�8���Ɩt�pq:�Y��y2��vt�@ )I49E&Ȓ�C��yR�
U#<��!h�8�D0����yr��>ax�&�L� ����1�y�f�5T{�sJ��D}�<���+�y��ߙV�a��+�$����gǥ�y�MO4,H�b�I�!�z���*��yr��rI�r!�q�����Q��y���옰�Hq��]����y��$;j@��IK�\*<��b��y���[����4�X%nq����.�y� ֊(�X �0"�#2��C���y�&[ ��9p�Ԕ
��X�LY�ȓ%�r�I%M���fkՓ.0q����PdlCC�e;-��Q�T�ȓt������'3�Xp`�*�&lx��	���P��(fId�d�V��d��ȓ2,�z�'F�VмH�&F՟.��H��e�6�C�C�_ h��.�?�8M�ȓ4�����Ѻg �p�]�z2����>1�v��.5��IwG�VE�@�ȓZ��ٕc+?���!���I��Ʉ�9�Y�WkS
 �qb�Ű?i�a�ȓ8	��Pa ��Cڴ#� �$։�ȓ0�v���L ��}�r�X�'�ZH��m�F�����<P(]�Ģ��t�ȓ)�p�"���6q�6�	'��lpf��ȓ�^���Qvv�k0��^�Ѕ�<�HaS�!�IL����ˎ�3�6X��\�H��զ�X���AXpՇ�dLu����1FZԊT��r��̇�Q;��jA��M�6e�7���"�2���{y�l�d�B��d���7N��ȓi��}�FF�s��(ڡ�ȏ%"
�ȓR�v�`j@ʠ�v�	X'䱅ȓS�<�"���	pxA�$�́)̴��tL��h\�lR^Ĩ�g��_eJ���uԁq� Jt��
�Mxp|��S�? B��f�;fl��MNA�fH0�"O�U��@�*@�zj�B |B�"O1�ƀ_�S�� � G���"O`=ђ �/S�H��#��F�s"O����۰C�,xP�#�*��Q�"Oܭ��ϐ�j�`����ыزA�7"O�qj%ӑ +*Qb�O20�v%:s"O,u*C��*Pmf��BN�j��dI�"O ��� E7x�UC��S#G�q�t"O��yCjZK�f@9{@�x�"OHU�0Ń�:]t�����$:<�x(�"O�-wF�?z�L�����+�4H�"O�`�ӡYnT:��k<pCp"O�t�c`S�YJc'x��=	"O�� ��;*���+6:��Pv"O$Ѫ/�v�u '��`<���"O�@��� !񲰹��?d)�IY�"O�0z���vo>�8GE$O𑺰"O*<����5R���c�3"�|I%"O��XV퉤3��a�锑7\�1"O0�x1'����B8H%�	J�"O8�&<�^�#��S�6��a[�"OLiȶ�$ L�a��-�؈�f"OP ���R&��(��##��	�"OV}Yt'�@0C#ۙ�B�w"O���SM����1w�F��%�Y7�yQ�v���)�?I�A�D
�y��֨~�N! O�	1��%XF	��yR�0~�<c��ŇQ�l�pj	.�y�F XCR�ʗ�I|�50�F��y�[�Q���I2�X�:����& ��yBF��f� '��9��,�C� �y򂏀n���cH�*.�j��1�y�BS<��1�&��)�d�ReӅ�yb�V���QL�6��D�!�,�yr���y�e�BD��D �y� ��|0��ҡV%�IS��(�y"I������� ��Ezp9�ᅲ�y2�X�_i�@$o��JQ
Y3�y".� 5�.�ժ�Z��U0�$��y҂�1,A A�QGD����;�y��	�j/>��b��S\fE��*I��y"�]
34P�P� �+N�Yc��^2�yB(ܿh�x�5��0K���a�V��y�l�q�.q���.d�\;�I��y��
����0䭠Pة�y"�\@���y���	�xP·&�y�F� >�$h&�y��`�ʛ�yQ�0��b*ė.� ��ƕ�y��+A�@��N���Ȟ7�y�V0%�4��Nx�h!3#/
��y�k�DT4y��Fޱh�r��B�N��yD֙sZ6����o�ZT���-�y��I�h%�0-��jpv9�qɔ(�y�k�9-����*�d��p@����yR��;0�e#1L	V�̬PlF��y2J��6�����fX9L��ThA�9�y��]�0�gD�;C�4��-F�y�!�N���z��Ov&Yf,Q�ybN� ���"��0tt���
�1�y�$E/Z$>�"���lX�+7l�(�y�H�����R��&j����fE���yr�aK�Ph׸^<95c�y��G5g�p��ߌ^�l��$���y
� ��06��)�!F�$�"OT����S23���3h��`'\y��"O��CT�� u��@��i��D�r�"O�Iې,Dw%�}�vJ�|lp�`"O��:�D�#4^�M��?v�f`�q"O^�ȃ��>G���f"N�7ռ%It"O8�A�:v���P����PИ"O`�:Q��KG&��FY#o�X���"O�{0���_����E�[�.��"O�!��θ|���T���6�B"O:�:�&� c�6��@� �Q��':���S@4||����A��e��8�'?vab�E2}�pi0��o|�Q�'iu�o�2�)өa&h��'�0�J�!̄��pH5��O�$c�'��'��x�	3%��p�J�'�δ˂K
yo6��E`Rz�h�H�'�V 	�靘d������Жt�"���'.̉��/��f����AK�C��m��'a�b��>�"΄4�У�'�ԹE%��M� �HT��A�@ �'�2�'&&JvZ�p��Փ8���8�'p�5�O�,N���W��zJP�'p�X��_�ȉ�FƋ�y!`��'��5	 ;[�4r!&�9v����'P��� ��3��q�ڨc��� �'IRX�0K;�H}�p����؋�'�(��uյ3$��e �� ����'�^`Hg�3_0�+�,v�6;�'W��6�ۦ����,X�kN�Dx	�'��ص��$1z�qTEF�>�%s	�'<C��\�$��M�3�́gy��	�'� D��,n��<Cd��:1.= �'�����-�}c��9�Js;� ��'�$,Dđ����:nQc鈫�y�/j�@:�$-�\��,�yrE ��Bp!瞑ya������y��$;{�x3�!وjZ깊C�y§ݎI"�K!%��kp�e%X�y�C�?T��J��ĭ*�qׁ�/�yrD�l�&! �B�RE�3W!�y���D~u����5P5�P�α�y�._3$R�́��^�;S� pA�Y&�y���g��鑪##���[�c�
�y�唝Mz ����P2j�CZ��yӏ!��d
v��֚Q
�Mә�y"n\-T#��cL��ȴ\ȴ���y҆ۧr�tQC�P�3�ۆ�Ц�y�������ei�*���y��Xx�]���H'0�(9�p�ص�y�Θ ?t𬉵��b>�SЬǹ�y��0�*�F�R8�jq�����y£݀#R
])�[#-�%��	B��y"-��%�,����Je����yR��t��dp�E������Ƈ0�y�:>��)�������C �'�yf�9H�R��@�*ݜ��w���y�m�s�:�р-Evꄚ���#�y�NֆKh&���E;i���;��E��yb,ƹw�B��6l[ �,��y�+'N�cd��S���Tk��yBK8m�����5rb�I1�P�y��7�~r5GZ7�pY�3@��y�-�?t(�#�眓��ܣ����y
� � )6��`x�;��� �>�0f"O
�x�Iº!R DL
�,�Ku"OF(IQ�2~��I	��̦bҞL�u"ON�H��5e�PJ�O�G�JUse"O�5jG�˧5�(t�Gi��v
�"Or&�5S����@#ә:�\�"O�y���+Lp�#)
1P&���"O>X� ]>)n4(G
�h�Q�Q"OX�ׄ�yT�9s�EZ�ao�!"O|���ʞ�	�z �c�	f\Щ؀"O�pw�,S�r�1UL](O�T3�"O*����?y4��2�B�k�Ƞ"OI��DTO�d��t �>
����"Oh�3�杜�ZE��\�Pi�!�"Ox�C�E�}����Ƣ���C"O��R�d��e̸���5W�XthW"O����%��2���Ж���Ϊ�P�"Oؠb��T�*`�4�4��x�Ib"O �p�� ~O ���T2j6% �"OPh;,;/��������&�f��"O�ls��Yfd�	CD
�G�T�j�"O�-c��3&6�:Č�����s"O�<�6�[<`�2l�41�b�*"O� �f8W_V���I�&d�&Iڳ"O��rG,��cAJ�AFC�,	�"O�M��G `�X��!2���"Or���5�5:�B|/��:�"O��yf�˅!)� 	 �T3�Py�n�B%���@��D�����E�2�y���>~w,�wfhR�ܫ�+ ��y�#��00�2bK��gL�a	�B��y��,4 �9���dJ�qF����yBM�{�jL��HVt-��ƍ�y�ƒj$��s��<;'NA���/�y2��%^@t0��/���2q���Ɋ�y�Dza0D�D�ټ{�,y{2����yB�U
<�hL�g��*R֘2ポ��y2��3���#+��@���"���yR�м9: �	7�̺�������yB�2[�Pi� ���4�1��!�yr���oۄ �'��ؚ���G�y�Eē<��0�/]�AɮH�5!޵�yB�M�g���/ڹ=vde��L���O`#~:!Z�;��af�A\A�q!@�8� %��K��G�\���Lf#�ȓ�/D�� &盒��\b�(�Yk�X�\�!�D�6�6@R�j������0b�!򤗶}�"=)V�D�o|��
ԅ�H[!�$�-5��\:�-�'vD�aP���gz!��
��q !bPh����S�_�!�D9. *�h�a�TI�T��Aj!�ũ�
-��.��WE��ҡ֖3!� &6�^=,y�.��Ą��:H���'Y���n	-t�~;�
�T��'َi+�(�Tt�3�D�!!ː�	�'���#�^i�XB���o� $��'��{��0���J�F�g��,��'�*��C�]�i�8�a"O9Sf`8K�'-P�� '�/plh��\�EO�|�	�'�F�P`N3+��ط��:/T|��'��؂ 
E��p�ㆬ@t�؝��'��$��� �<uP��ㄟ-a�x"�'����'$�!v������].:���'�*�������i��nG�B�@���� lD�P�N�!245��'i{&��'"Of+�O��Ȅ!ׅEl��i�"O��
gm
M	Z��a�C�&�xd�Q"O����N� ��]��`߱~���3�"O�� ĩ@"s_��gm�a�Z�"OP�4oīO�|���mq�"O^4�q	�2H��ahA�E��٠e"O�|3׬ρv檈��/�%.���E"O^D�CW%�Z	W�B@�
}6"O�8�E�z�a/�?���ѣ"O����M/'o@� #��-���W"O2��f���Y��=G�ղ<���"O��D��0|�R�� ES"F����c"O ��@@M��:Ac�Scr<a"O�ũ!oH:^�Fd@eґ]]�� �"O�I�"a��]�V�&�M/nVzU)!"O�1�uT�V�i�u-L [D�I!a"O�̙Db_)��gl�!/�E"O��ZUl�4O��C�k��E,޸�6"O�jU�̒X�H�
1Ę![�0`�"O��:��_Ne����(�W��`�"O@���o��x�B��5�
�}_��[�"O&M��I<<�6���5OLIY�"OJ�q���2���T� MB�@�"O���D���L��X��±=�\J2"O9K1IN�B����`�T�N�"O�,��nޅ-��!Sâ�n�8�"O"0� �/�Fd �'F�|n蒀"O0\��K�~'`#a�F���l��"OYKU�T"n����߇&��1��"OR,���#q���b�-`�إ:�"O��bV��lpB2��M1!"Or�B�W'O\i�A܇*�~���"O
�'u�J}�i��J�~t!c"OJ��'��G��jE֗w��y��i�����p�¤ua!�j>3W"O�4������]�-"WBl�sq"O4q���Lr�Pǭ��.B*db�"O��y�O�N-�J��E���&"Ob��G��7�(��։�3 3�8��"O����JP3_��[�
�,q$����"O��QCf�'��51@��&�E"O5	a��e}�}+w�&A���"O큁g�~Z�5k��4���ˡ"OzH7�+T�l�rfD�:��R4"Ol}x&iĊ(�:Y6��RqFz�"O�]�g�=B|���A�4>>�I'"O�x*e�$���J��O4��*�"OF!�W�u�1q�,�9hDt�"O4�sSTj@uC��4c�N��4"O��rw��?1\����<Y�7"O:5���.q}�J��%�ҽRv"OA2Ui�#���9�Ɵn�Ġ�"O�4���B�!>��B`6%��Ds5"O�$��C�#|��u�@E�9a�h�"O�1f��S
B@�b�h�e�i����$%5,0�0��?��1PǬ��E!���B�c���i鈵��;�!���`5� Hš�a{`�ր>�!�S��D��g��g�D���B�^!�'q�ȈZ ԪK��������k�!�dԐ?����W'i�d��Db\% !�Dǩ3��Af�O} ʣ[7)!�d�&&K�U��$��%\t�s� ߯e�!�� ��8���d�0�Ҵ[b��"O�]������A�׹{;��"O��7	"BRd$�@$V�I4"O���o9Z HZѨ��'�\`)T"OҐУ�r����tbĜ:��X"O���e�	T���b4Z1S�x;&"O������n)*����v�x��"O��{7�U��ȭb�aR�p�Z`"O��D���T���ы)�܁��"Ot�t�^��<�D �Q�r�@�"O�T��ʅ8_�z����*�r}{0"O@�j�,E8�\���;��ف�"On��D��V��a�HL�e��8�"O�ݙׄs�JUxw�58�\�P�"O�D�� ;w7�A�6hA�Z�:�r"O��ec;4�v���ܚ�R=x�"O�=٢�K�~j�B4:����7"O8����)��M��kI�pv�`P"Oȕ�b��*i���)���vBT��"O\��1��o��'�U�"ObU(S���$�T�������$*!���=8-���S�}�z%x��0 
!�dB�^b���/f�~��`�4Q!���&1̈I��X)6 ���(-VC!�DH�b%��fT!�Rm�gF�,9!�䕦]j�w@�>	��=�1��R!���8҅�F2��ΕdӼ��0"On<:��Q�~f�ҕ�d����"O��9��9��Bp��_��U��"O��B��ųN��"��U�~^�u�U"O�q��ć]X�4!Sn�[Vd|p#"Oz���t��5{2-��9:R� "O<��ƚ�w�x��잘r8�|R2"OD�n�}�䥰�lچv(�Y�T"Ot�D�5PxS��u�J"O(� fa�B�z5�.�"�9i�"O4|�,M�P��`@g�4
�0*"OtTUl /Jm� �QE
�x1fls"OT�:u���uh��Ѥ���r�"OX�9��U�l=0� ��� Vd����"OZ�f�Ԃ
��U�g���ja�p�"O�ITF��#�Fm*�F@����# "O��9f�����s�£}���"O�h�*$6pQ JG�hV��f"O�!��i��[G�H�L؁"O��B"�Ԝ8����i4i�p�S�<A��6�:�BS&=�2]����R�<����8v-��%7h�m�d�Z�<Yab[Y���¦�J���D$�Vn�<�b`��0Fa�L��̂D�d�<Q�%XU�sUON%'��۔��T�<�E��'H�@�j&���u(F���N�~�<	�K�;vn|E����"	��q�R�<Q�����,*�"
 u�m�O�<i�/��9�"�#�+T�F+f\�
]�<�T�d�� ���p�h�k�Z�<aV��0H��t�&)�3L���cDW�<��a@9fR"��ui���z�<�t��L�,,P���"0�=���1T�t�QH�;l���E��0c���J:D� �	� :T^��E� >�g�8D�$�EH�`�"�J�.�-�V��!+D��:gi	6�<i 4��� XjJ+D��Z�mB�j�1�M�o����*O� l�y���K�]���W�7���p"O�����$�p-ȄN�:���B%"O�\2UFS�tuC��F��Ґ�"Ot��B��>�X��+.����2"O�Y�Ќ�	j�tR d�
9a�x@�"O��?AU����d@n0Bhò"O�%q4�CX�`�0��\�IO�)K`"O4�P�ԅ 0�����B�DG ���"O�8��g�L9��J7o���"O�!����+�p�맭 VRP٫p"O�@�!�Bxr�ub�3P`Nla3"OLK��܈1�b!�6bɞ?�@U
�"O�ѡ���)P�=s@?5�΍z1"O�i��E�6M됡��E��S��"O�˳ ��q& JG��C�0�"O�ёȋ�8Nl�3�T�
~xA"O� �W���l�1��R'>�� ³"O�z4E <k��t
U���Mj�C�"O��I��Q�jش�#LP�`)��"O�+�,G�.��)�gj�N�:��p"O`$��B��<�c�ߟӲ{p�'�1O蝹R����(��ù�J��"O�0:�>
�T���ǜ����8�S�iȒN�`���²2[�X�v�Þ 1!��;h��˟�K;��q�J 6+ў���I�Oۺ���G�&��.(B�I4i��K����:�
X��Ӏ=�nB�	47.�zH	�ik��27BQ
S�rB�I4z�1�Þ#��l8���H�B䉶nx���B׫c���U@	.4��B�	���\с]��ց��	�%Z��C�I�Y��	�6���F̐*�H��yE1 	��V�"G�z��1�Ѡ�yb/C348�}rO�?M������y�jFg?Y�`W�4k�(@� ��y��Č��=�CF9}�}r�"H �yB�U(L\8����7����/���yr.�� ����cjI%#R��be�̹�y�gL�rLn��dMɘj���\_bC��;}��h��|�6�P"�,B�:B��&Ǿ}S���L�PA�f�)BTB�>s=,��3ȑ�1�$0C/6ZB�	�1:�A�@�pl�]��W*7�6B�I�bRx�˥�\�J]�d2�B����C䉪$e���P�њV��,S$eŧufC��^�P �4:kҼb�e��A��C�	 �ԋ�c
�=p��0��_
XF�C䉒��2��׽ܜ�(RH_�x��C�(kPt¥韲1<`P*�	oC䉌<��A"�p��nФ^�C�	7�&I��D�z�Nx�S�P ()�C�eW
dpqF�		���MK8N4JC��%5tH��i��%�l��'"ҁ'�tB��*p�!�0ybx�)���_$C䉈&�FTC��Ì}�*���L$-�B��	-���a��|�dJ��ȴB�7bd�p�E�Ì
ό���!;�C��(M̵PV���y|��@g�dC�	�e����s�ߝZ p����zxC�	H�j��.)�йZ��	�N�0C�IQ�} ㊅�*�L�0̒�/�rB�	�Y
��ᦂ�#�A��g�?u�FB�X��LKC%�X��a����B�	8k{ґ(� ٭++�Xk����Y�*B�)� �պ�@29Bpk�f^��A�"O�\ K� �0�7$ ��4�"O��C��W�>�.|%H���T��"O��7�ڔo�*<q��&>D�4���Q�a����7Cƺ1 �������	>24Ju��LG��r���1/���-��E����餻�H���Y����'�J��eP��*$"�d�^]���I?>V �,ʓ�hO���"�R�	U�k�X���Hޙ,����cœ@�?Y���B�j�D�0�2xE�)D�Rd�K�W�4x�_={<u�g@ @ݬ�0�{�T���A��L�5ŀ7~��F�0D�H��*J:@��\�G��1k�zg��O��[�)߰>�'m����ɷfk�0��E o��l����!\] ��Mޅm�čr eV��P�V��Z$���'��U#�⌬J@,���aZ���}�8D�t�zf�2�.	�����|7�x��ɜ�o�Z�ǌ�h�!�DΛ6�&��`�h�:Bl�2~�Is� x
q�� ڡ"�V(c��<ip�e�"lRAdM8-� �b���_�<!A�7Y�Ak�ҏa	2�R��>V�|���5$� �0֠��o*�+��D[�]xf ���M�N\)r�º��y��#L�FH"aB�������� s��i� �؜^��0�bb�'��*G��F؟�!��"'<�
#OS@�.����!�d��dM �+�bPn#$:�*c/�A��dJ��Pb����Y��V�Ҙ��yV�+��($�z0�T����(1�׀�=qop�z�M��LQ�Pi�KR�'*v���)i�;6���%h���#�"*�q�!)��r/"�T��n	"n��	*A�H�G ��U>
� �F�"S���1�� ���R��4d���W�B�LPC)O�)�&�.�5��
��fA`�HG ًҎU�� ���2F8UŜ��pm��_����4 ��`�ǆ	�s����0#�IS��= 4��eO$Ц Qi���ރBV���OFɩp�S�{�B����w��PZ�';��R ˽7ٚ� ��o�i�6�,P
��#[H�H�m���l:�O����Y�y�OGjF�\kюK�y=���ψ��x�/Gh�Tѳģ�"]L�+��L�q�`սN7� �eA��D"����і
�X��T��<.ࡰ�O*@�`�m��B��Dυ/y^�8R��9j�`8��ꈃ�����D y{z�Zf2.����ڹK�B���'�Oʥ��9g]t��B����:�����W�D1��ņ�� �CW��x�ND �s��h�V\<@��$��!r�Tv���yҤ�N�N�H�M��j�Q#���D��,E�#����&��5S�4�������P�>���w��ȠKӛT��z�aS0rp�'���0gF>����6"�,�4�(u,I�&sbh��h.~ɹR��W΂�QR��:�ў����VS28 cF	tP��u�&O�������u<X��@BN/9H�׋X�&��"C�Ē9;F��\�>���R��-0�L�D4�S�'%<����1{F�Txd�ǤWF�u�'������M���`FE���k��ɟ	�D��Z>�k��S�i�A�a����o#���<G	/dŲEy��)$�ᩃA�?t����L�"`��jb��:��O~*a�8��ϻp| �r�b�3��!��J�d{L`��p~��d��2Us�ku
¬e�lZ�*žOGB<��O�S�4�
v�ɤa�^��4DD3�?1�r�����	�Y�r��$͖>�0<�M�����m�����?�lb���6<
\�ZB,6'z����'t�Hd���hO1����-�m���L�8�<Q��>!�i�3u�)@�����x]�h"欃���IOzt��i�����Z��QB�2]0�V�d+<O�����5��5kVl����#�`�b�i�2e�jQY0!AB-�O��.ʃ
�b�'��x��9F�&4�j:z�C
O>y��+H�@ Py��IB�B���1,��$ T�6?�*��a�<bZ4�ҫ�������ɿ6�<��b�,:2���A�J|d��D-9:�:� ��Izh�C�jS7fG �ХL���Й!Hˎ^�veCFDP����.�S�'.jl�B���.��Y�E�. .��<Q��&���fV�v����Ҋ��j����&�+2���Ɲ�G}Z�Fx��'���c��03�,�z�g�=8�dQX�;��CLB+Fx�ыCk���(��I�2�<|Bb�z�$)�E���+(���\�t�S�f_"g?IJW.��]��oڎr���SԌG�H�̍�+c8�,y�K��<�J��R �:�dh3�;�Ot���ݒ4��cR�AY��$��x\0tc��$C�)� �i�J�P�9�׌��!!��ۦ"OYR�LT+l]�6%�� ��f�<�bDP8���� A]P��[wĔF�Q�7D��"g�S3a�@LH���	���ء�6D�hd�JH�|�q�@�+��Q��7D�h�`P��r�i�l�$v*����3D��04�	�|v�1#��J;�H���uӤ9��)���$ r��l#R�T,FX	��a2D��iƤ��`b�� Ri��A��P3��/D�@cf��;J�n���$7R$�<b�h8D�p�Pi�?8��;��(�x�A`7D�lqA'�$`��`\'��,y�'D����#�q�<4k���l�rXj&'9D�8h�B�(�j����̹78 	��9D��!�E�1exTXCd��$D����3D�d`�A�;�4c�HF+:`�$�"D����P )I� :C�
�N�~��"� D��#���'�����.�F�lu!B?D����%@�p����l��U�:D��� G�fi�PP��d�3¨:D������P�9b$N
H�f�ڳ�9D�tA@�A1�Y��H:�nh�"D�|C��	�j����@-F!�L|S@>D�pѠ�_�5�s��L����w?D�����ƶD�D���B�&Ԟx��.D����
<4�4����G5 P�#s6D���A��J_�"$��:F"�|X!�䀒E6}���F�+����L��M?,Q�A�JqO?�ʷ+�X	�^.��%H�i!�D��-+t� ��,:���Bǔ�Ya}B�Ωu��D��v���Z�旅P�4���7��awn].�HO�����O
��u��=>���N�>@��"O���i^3�t�p�m�<�E8�"OԕS�c�T�X�;��`���"O��ʃ��3%�ne��*�hL�"O�`6 ����q٦ꙸ �-�B"O��+d��:�Y�ǉ�z����s"O@]0䪋�V�zX*��f|�xRQ"Oxp2k��M�4y&�߃.5���"O�\P��U'=�N�j��b&Ĝɖ"OH9r	S�]
\ a����v!H"O����!+Vh�'�D=`_@��1"O�HhT��`T�7$�"%���1V"Or���I� �sWb�(~�Vi�"O \�G Z7F��aZ'��4��"OSsB�r��k�7A~����"O<��B��C|��,N5���"O�*rc�d}���,4��
�"O���GY+$t�1���!60�I�"O���I�[�`���(A)ҡ�%"O0�xR	[�!�Ա~F̊""O�E���0D=��J �ATl�$��"OŰf�3`="�\I��T"ON=$A��{��D�.6�1�"O>0*�J}y�/ȯQ��H�U"O�E������"N�3TH��Q"OZKf��?b��aPW���zb�G�D�<�LQ�h)"�I5�N�L�,Ae�Z|�<ɴ�!�T��"ǒ�i<f �GDG�<���$Cɸ�W�/6(�x�D}�<Ig��0vt쳗�MD0����\a�<1��3A�~�#⡎L¡��^u�<yC'�T7��j��){�w�<9�"E�	��L�SF�E��R�MJZ�<� D�ۆ@O6@�����0~�����"O��eFV4�8,�c�*U��5y�"O2�:�`9pa�qK�:h}�3"O^-	��_Y��ШF�I(Z�p��"O�y�,�j�|��R�MlE�9�B"O�tH�[61�~���S	P!
Ly"O�d�#ł;�JT !a���lL�B"O\e��`���f�� J���1@�"Of�)�M4! 0�6�ێiq�0��"O��Y戓tо�;��Nd�i"A*O�LhwG�u�rH E��Z�*	��'�6�ٳj��8ܠ��L�&�$\�
�'Ll�i��� S
2�8P��.�IQ
�'9���E`�5+�~8Ѣ A�� k�'��\{�ҪI~���-V�H�#�'��8J�E�!��M�J��1ڤ��'��B�+҈QoR0�q� 75|��(�'d�ԣĕ^�P�2�H7)H|��'u:�)$�8 ٸ�aE�D�)�\l��'RBhKQ!G�@U���,�B���'�1JV��h&��{D�^
i���'\H�r�؈?1�ѦjR�f�
`I�'`�q�f^��t��ֈ��7��#�'_��2#��w��ܪ�-]���X�'h�$8%d�	��P v����60��'�|�Ʌ@� T8���T�L�dDݫ�'�`è�,0�觡�<c���'���"�I�1�ld@���#/t0[�'48���J�4v���8���:1Gb���'�>�8B�J&o���1�Y!0�`s	�'�����#ʳ)UBi9��_
]��Uc�'VaQ6���),��@'S�_�`
�'��8wB�R�d��T�L�i
�'=�)�f��Ơ*@ J�@���
�'m̅+4�� d���+��B3�-`
�'B�]ptj}st��f ��;�Ё�'k�4�V�;TL��Z�m��0�&1J�'-��Id��.��p[ (�PF�9z�'��t2�I�8u�]��Y�~��X��'(��S!�ԔJw
�
Gr(�${�'.�����p���b�a^�+�'�Sg���{��3j"0�'�
I9q�1�"��B�� ��'t8:��ӼBB0�jq@��p6��'$�H9���%��Ѱo�0F��z�'.�;�dY"l+��[(>���'�d�0D�aдA�c��?�μ0�'�"��	7�F)U����Gz]nC�I�B��[�IX0.� {��\�B�I2��a���O/?�)p-��C�	M(N�����Vƍ!��;o��C䉆��)�cP�C,��`'`�=w�B�	9{��=X��Ȗ$��Sk �`a\B�	0��yv�������^B��p&F� E,J=d��!�W�]*J(�B�	�nX]C�8>�����2��B�I5�qc'����9�-�z��'��u��̏/k	f	�J,�4�'� ܈�ş�H�Q(�j�;2#�A
�'(�y��'W.z.��X#�����<�	�'v,�"%��pjj�	�h� �`���'�T���`M�nO�i1�=!�D���'�j���H�f3H�� " � �L��'B�M�@f�b�0a�D�
��� �{D��5sK���%.ŗ�Պ�"O���$`��N^��8Cm��>��
�"O��@�jA/<�"A�L�1K�$|��"O�(Ʌʼ*��LC�N2 ԈF"O���OX�+��pRTjŬz>NpC�"Oꀉ��]�%!"U�DX�`��"O��a�'�4^�b!*`���h1�"Om0���E���a������8�"O8咠bK��:aB5
ļS�d��U"OH�zÇC�r� �S*٥�x�xb"O��R�M�b$������E�&�{�"O|XbЦW:��P �[#S����u"O��bQ�:A�Ó�T�(]
�p"Oԥȳnŋ���� ��hQA0@"Oܑ+�ɪB��|H�o�:�� ��"O�,�	��J�&(2Q(�-��qQ�"OL4�%�[�>��y+��B]����w"O���B-����C	l�}"O��b \ FlXU�&S� +rq��"OxÒ��:��1j�K�04����"O6��EC�y�0HѠ����hš�y2&�����w@�!~��������y�LM�f������aD%�y�J�!z��c����M� �B
�y�AW9���K�ʋ:�̩�p,M��y2-�)m>ZQ�DS�,�N�Z�M1�y҄�(Y���a��˯-�x��+�2�y��I P�d-��fN0HИ���X*�y!��r1 ��'N�� �Z��yB���v
�	;$)�(_
"-��G�;�y"J�|���ybi� �������y�%�z������W]�8j��]��y��РyD4�(SȡJ��y󌐱�y�I5��q�%+�2�p�òe�$�y��	f���
�D�9����[��yr-`�Z�8��[��^���o�;�y�K��y,�S#�cT��&iS�y� ;/�������,����\��y2[k�y#i�>��Hԥݨ�y�x�B[ Mni���C>E����'�$4�L�(.D����43���S�'�,�I�j�+V�����/���'��&o���|px����ީ��'MB	ҭ#pO�`��N�ԍ[�'��[2@�+SN��`�A�bG����'4h���X*r�$!P��Π6Ҽ���'C&ԯ,	�f�z��P0y�P�8D��P !߀cl�|�����Q$�-D�P��L�*>*��s-�� 1 ���*OJ,˗�8\@���E�2" ��"O���ee��"�8a�@8�p��!"O�K�'��t ���J�T�3�"OT�R�M<I������:)PU(B"O΀� �		j���S��X�:�"O�u� ��9+R01 hB�*�)��"O���F �"���?x`D��"O�@0�E�<�r�*�b�3j�t� "O�-rRB\����aa�:~�~e��"OZ87��>n,��!�1 ׀�("Ov�5�i��Tq�ͤ~�^i�5"O2���ڋ[�����Q|�l�J�"O�%�ǔ�k����'ƿs�B�ɷ"O޹�hK"8=���'�b��-H�"O���/5c���I���:0��D"O� pU&*�4�Xp����'#��yɂ"Ov)@g.��{�t9��HŊa�"O
�ȓ�I��ZDCp����4�	s"O�!��S� =>�C��$��"OօI�d�v<��8���;k��|�0"Ox�#f��;K"�M�%�1��i�V"Oz�����9��(p�)Χ
ü�K�"O
	в�\��ݹ�g�2&��0�"O"A�I�rth|Ҷ�	)�*U2�"Oz��a��z�f�`�_�r�
���"O��╯�-�~��d뒺(�V��c"Or�[1*�*6~��p+5Q��r�"O0�t`�?� ����~=��"O� a�6 �Ll���6-�� �"O���E���T�PZS#�5�V�0�"O��#�a<]�t84$K�M�`+�"O섊@�6�$#c��5�r��"O��Fk��2��s�� ���"Or�ѭ+L�����aV$A���v"O���m�D	И�|(���^%�!�䍌d��uYg�M�X\��@o^8
�!��ժc� `��̊�v��!h��O�!�D;5���Ϗh��!k �%O�!��$5 �]���[,�h���J�!�d݇>��̺&���W���ԼD�!�D7A�.�1�.@�X���ǬP"1k!��'�!*�K�>5bhL{�.�'�!�D3@]�1�����,:��!PF��S	!�N�,HLDZCH�=<���uF�g�!���B>l��@  P"�xӂ�"�!�$V)�����J<J�pɉ#K�g�!�D�@����PO��+`d�
A�!�U%8�TA���#`�PdS���'^!��.�MPR�TǊ����M#b!�d��R��F (K�FL��N�� Z!�d>��a���.
~�s�� �Y�!�F�6ʬyr�._<o�¬
'KL��!�$��1�@�E�N���U�ˆE�!�D)�zՠ�� �H:�ı�IъO�!�Ć!p�2�+F��^$ܑ0(�2e!��H�9���jU�3|	�M�4_!����D�F5�$�a*&OH!��.vI�H��D�;Pa���΃VO!��R����",NH���H��9!�$O���"Ce���sEsC|B䉍V�\-)�R��j�����PB�ɶ��q+���? ���%�9NnHB�I��r�a�e�?,�Ȇ!18B�	�;�P����@�J�>��B�0Q�^B��z����@��>��K���laXC��NŰW�o��D��;W\�:�'��[v���"�,%*ꂺ)A�5Z�' �`�&�X�#�>����A�.�&IK�'�u�`�/
^EC�+��&v&Y"�'~��\��{�F��2)�
�'���!�� �&9C�.P�H	#	�'��5z��%
��H� Fت�'��:���Z`�CW@�h�'0�U�'�U-i}���U��-`���J�1�hM�c/�@����'LA��6�����Y����UR} 2Ա�'TPy("-4�)�iD�3�	��^� �z�������v ��8����f"h���)�$D&xP̤���~�$ �O�>Qrrn�%J�ΉQW��Bp����B�'�TX�����E5+��諤�.:aؓ-�d�^P�?�?�� B��6o�>3�X�� W�Z��؂���-Len㟒������<=����%�%�!���>1�k������O�j ���@�W�ꄐ�.�2k�*%;�'`��D��S�5��$��Q�r���5O��p��uS�/������s!�G���i�)��G���Z�k�|��_Jx��K�O֕1D�Ϻe�Љ���r�A=})��$;b�s�~�SD�ӑM����_C���D�!OU��Ʉn����� '}��h�l��ek�,���C�([�s�e�G�ƈ^��l��(~�S�OG<��S��1������,t�!r�9�8㟢R�͔Q�z��D�&+�fP�@P�E!�O
Bç0_�|7N�<o�N�y#�-o�d�=��ַ�?��i:�6��Q+ɼhc͈��	?��y��8�����\�[l!��뗴$��A!5�ê�~r+�\��O�>��	��/�\�5�qu~�g��P��lr���i["kl��qg�ȫ��U���" ��!�?Q 5�T���L*M��ay�	��sX��W��9 -D⟒��b���q���)��ۼO� ��$�>�C`7����O��p���	�P�
� 6�ɲ �|�k�'L:�BE�%��~*&��2 �~�cc�Hi)��:b��&�$}ru&F�}I��
�'M�a��C�V��1�*�v�"Th�'��[�LŎmY�X�ec3�L	@�'�X�r�3��-k�f��y���'��A�"H׹L��t��k�4[fPj�'�4*��-K��prT�H�Lt���'L�Xb��@��d�-|T�颦/9D�Z�+A�r���@��IV�a��2D����X�R��,X�-�yBV1H �0D���¢K�	UA�8j�4�R�*D�,�S ���M*c�E�dD{��#D�����E�>f�#���.��s��+D� Rg��x��|��eNp@t)�(D��Z*@�^����(��v*J�ZC�&D�0�oW�5.��rɜ�p��`�u�%D���AI�=0���Q1B��rȀ,i n(D����k�"��5��Gv0R����%D��X`��@����WFʰoKH�s�-D� ��,�9C^y���9�k�&D����ϓ4�r���]��!�d*D���D0	�9@���6S���A�&D�(��jQh1�Gf��逹	B�8D��냷T$�j_�1��8d�\&8�!�d�t��(JW$��7� �I����!�dBU�\)��J�Bܔ�֧EH	!򄎽
!��0���dˤP�E�F:	!��
� 1`�_�Y�1�1�ʌg�!�ě�y��}갆ΘQ���1�ԇI%!�D1M�i	�+Ǚ.�H��@�"*!�$�#��
��6.��Xc��7!���9I����>s��� �
�k�!���=�8Q�$j]2�c�GܬJ�!���d�(� �uS
�!��\/%�!򤁈 ���ბ��:����!�$�%4F�H[��T#!�|�V���	�!�D�H��I�1JՓqgx5��JI&=�!���#��H�@$Y ͓���!��$.��yKs��|Tt!Ec¹3�!�U?8�ZAsDC��u7p���B[�:R!�ę�0X��uf�^)$l+�˺h8!���Z�T��m�>2�D���	Q!�d��y	�@�5�#�U�$3!�$Sc��%k𡁬t���HR΂�{!��Q�-&� s��C�}Ҫݘ5��C�!�dV�D >�ㆢ Ӽ��\r!�dԏ_�� �1o"��+�2pT!�� DP	G�6Hl��W	P�p$i�"O���`H�%�|����B��	�"O촪��2%�5�&æ ��=�"O$���n���� (�<p:�"O"�#���o����AeفH�*�R0"ODYR�$�%Ip9��+�0�s�"OD��$�:K��On�"��#"O��-E�2�I&��-3��Ѻ���yR�=OeD�X���=,y�u�R6�yҢ�R�A3d�#iX@��ֺ�yRG�8�f�åjZ����Ԧ�y�V%M�*`���S
S��W���y(�8b�H�@j4LL�br)K��y���/�&���!��Cڤ�������y�$=�<��+ ��	`��!򤓺P�&�ðCL�k6\��n[�P�!��R?3�.(�DHQ�0���gK�n8!�Rq��O����Q���1	4!��U;,�D��C#&{J���w�ל32!��]�5x�������T�V,�Q@��\�!�$Y���T�Ur
�)�O�5�!��:��p���2n>� �C""�!�N�8*�pxU���n����� �!���m@�%�3_&ĩ���Z�!�d�7|1���͉{������R�F�!�D�����դ��{н���e>!��d�U��+�U����P
�P/!���GT�(5�8�J5�2#�4!�$W���,��{����(�n!���W���XD�8�d]H�E/c�!�R>g���v��'`�X��/?�!���	���:�& *�}R�N(x4!��]��9!�m�8�,�W��	1!򄉸hg��
��L�i�@DC��!���^����[�0(	����P!���[����*�;\��Q��J!�DL�OZH2��/N�A�c(�4M�!���x-�<�ÑW5H�Krl�5f�!�䅆��0����:q�d25�O�!򤄄SO�y�Ƥ�#������1�!�d�DLT����y��%�ϊ'�!�$�1��!`0�S7d������'H�!�}��n�6@�P���F��P�����'�����LC�i�@��S�F���'d����G� H���)��^�<�6�
�'aZ��#$@D�\F Y�%�60{�'�f���� �5�$	���۩M����'�<|Q/Y'+����$P<v�x=�'�(���Ζ���{e�W�s� ��'���iO�}� �R%���9�P��'̙a.�W_��K�����J�'�B}�󨌀,y�AЍ�VQY�'�~�J_$N�{ËU$~)`фʓbD�hq��iZl�@b�H�|���^���#�e�9�@m��ҁD���ȓsOn,�F+ۋ �Z�{���x m�ȓ1V!Y0�VX�֐;���1-%��ȓ�tH�ҡW_�TCA�Q� p歄ȓ">(X�4f'XG��e��#S�p��B��Ev�ͶU���D��v�P�ȓ"Vl�f�ǘs�p�
c�Q ����5���Yb,S���&mܫS�Ĵ��
��a�$��B2�!`d�@� ������,��QMF�� ��!]�|)��S�? R�ʅK����A�D/��Ӧ"O@�"���&6�؁���!,}�D"Oʍ�'��1s�N�PD�t��H2"Of�BP(R7vh07!��.���"O4	�/L�`NZ�E*1�P@"O�)`)�B�.�@$V�j۸%:R"O
���ZCt�Q�i�'�x�r"O*aSҨB�7 `e��-۷�:� ��d#�S�OLP����R0DV ����̔X>r�'�z�h�O ��8�bQ�<^c��*�'����Jђ�h�+`�F�Z�'Wz��Af�#A�����Ȓ[����'�Jѻ�H�)l�iia�[����'�r�i�@K2.�����K*���	�'z��8���#�3� O�ܰ		�'�n��&P�,���$���p�f,h�'��8a�e�rS�j����'�Ѡ�JT?���KG��<`��9�'Nhi#,��l	�)9�F�06���' P�r�!��������{;|�C�'wHl � E.E�(�Să�N�A�'�f�Tj�*(=�`Z2i ""�t`��'��Uc5L�΅R�#k���*��yD[y��*�3ޒ�;�K�yr Y%a��xA��tQ4c��
��y�F�"��h����>�~U���y�ۉ�Lِ��"����+͐�y�hϋ1���c�����(�����yb�p� LC i��~��� �Q�y2 ��N84�[�o@,<A��O(�y��N)&aF
aI'g��	�&BQ��y��ȭO0
���K�nj�L9����ybň�
�� �̒�5|�5(���yg�3
.� ��B�+���pB��:�y��M%�Z �tiX?2=�002���ybL�!���Q�ʼv�N��"���ybM�5/�x�bj�$v���P��y�
W�6��`�0V�u��H#BE��y��ÑtQD|q Fmu���ro�6�y���R%ʐ#Ɉf9(��4B��y�gE�l�6:"Ȋ[�θ9��ӓ�y�HO�����$*�[f*ٰ�Q�y¢�:��`փ9nh`��$�y���j%Q�B�0 Ҟ���K���y�K��$����1��1}�V��/�*�y2�@�7�0�y��O4_���3����y��;_�<a7�$vX�t(���y���S	�踂�H/: z��S��y"e�2 ����eԑ
ݖL$!�y�/�,4�,xZ& �{|h�kdŔ�y�B��F~�U�&䁪%~��E��y"�>N� X�K0P.*�!
� �y�k��(P��� �Ǝ9>�B����yNL�'f��1�f�*� a�p��Pyr�E-K�����T�}�D!�#)X`�<�aS�@s�8��ʴ&�P�J�d_�<�b���o����KV�p�X�"�mT�<ac�&��\R����T9d�VM�<9��)%�$P!�ֈ�0�H�*P�<�*��U�Թ�f4�L��"�`�<����R �b�İF{>9��g^�<ug�D� 3��+R�
 j`�	]�<��B!�Y�g�eh$�!$��N�<��h(K4�����&?�ċ�K�<� ĵ{�L<�li��꜕G���"O�u)��2�4�wJ�+c$�Ċ"OJ=�T,̶7� ����]�)rH[�*O�Y`�AZ4RKą��ŠV�8)�'�I��jJ�J�1��R��b�'6mK��X�<�Th�n�;����alN��FEf�(�� ^�@d��/H�YȖe%3~|q�'�2;����X��к��?@�,$�������ȓp*�4�0"+2c��1"��(���E�]���#�lyq@�jE��b"O�i���R�#��X�Y=-�"O�@�2�� j�l`j�S�"�� �"O4��"&��@�S�S0��2�"OZ���c\;,
�A8
Ӥx	n���"O�l�T��r�)���\%y_2���"O"�P헇>�`�3�h�FM)K"O&��E�Y� �W��1-[��%"O���$ �[�Y�'��bJ0�"O���	�)Th�2�&(&��Р5"OXőM��qC I��R�P���"O�4�3��. d.Idk�����"OL쀢Ê*��!$%�6���(�"OH4!�    ����8�tB�;`���rkҶ^�:��P�&\Oxb�؊��?zha�"�!g�r@��)7�hO���A/�x�!�̖VZ�<*&�7x,B�ɊX6�8�%\뚤(6@U�|~�C�	>h�V� �aߪ8�(1x��)it�C≠UZ�|#�a�:R9 d��>w�J,��' ���C���2C.�rњ�؞'Xў֝t�'�xر#U���h��9:�u��'�`�i�FF�8�<��aZ/X�i�'Q�#=E�4�x���%�Y�%���[pfY��y��<���xqw�ܖD�ў"~Γh�����D	C��H%���(���B?��'�a�U�Xz\��P� �[�x��	�'~��s/�LP,%�p
�&[�	��'�jIy�j��BJ� PN}���(�'�v��$	0)��=��Ȋ9r6����4�Px�� VT�H� 5TS*����y���9<�h$�D� Ge���%�8�y"ᓩ~Ŭqrq�ɧM����kޠ�y��F�i*�@F	
L�V�J��P{�����<���F�
�V  ��	A4��C�<��mM�/@�\J&#�+c�~�0��g�<9�L�FՀ�X0� &A�1${�<9��TU���&
��Yjp@��"�m�<�K�b_��s���lд�ĔM�<�US�-�}�鈄t$�8�D�S�<��ƕ9k��Ӏ$L�S���HC��L�<� ����D�q�\���@͸��k���0G{���Qe�v�j���0��5�՚��Eyb�l>���i�>n���C��Z	+N��F9�	͟��w}b�ț^ń�ʷfE�^�&I04B��(O��=�'��U�� ��z�U��cY<n�@D9���}�	jyb�'
ZX*���,b���Q.T7*,��\����)}�� ��s�s�@S��8�|E��!�lr���	���C�eʩDI�x��������)<��Y�OV�S2�#נ&��V'��z��R��s��\�';�I
P&�Xa5�'Y��3�˞]~^��F{2��t�	�+w�lD��)'��H��o�4$��[޴Ϩ�f����Śj�	�s�S�>3�=Sh��<��{��.�g}2I�Z�q����?Ԓ���ۍ�yB�)§�?������k��QA��q�d\֟І�	P?q�G�^��<9��98�)�c[g?I���Oȝ�<�IZ,c@2�j�n]�|��y	�H_�'>��<��4�M��4&p0@�4MN������{8�>����dA��N��䊰��w�x��!f��(O�=�O:��_�&��j$/ �<	Ap�#�S��y2D�y%vezvm�O �̏�HO0��$ƫ\�^yR���TxI`ch\�!��	}�
�ٖ�1N$L��[w�'$�'%�ADy��Z�R�r�l��*�4�[��H�/��|��6��|��}J��u�}_��x�'�ؑ;P���17�5P�iƼ%h\b�'l��l�D�O�'��'{�����Xn�ti��4l�FD̓��'��\�'�P;V#�<jJ.J�H�h^�k�O�]�I�L�꤬3nv�� �B�,(Bj��M���2/���bdK�>	A�A���r�'�a�t�N�,+�����w��@��lK/��OfdA���8�������x�4#X��!��΀�腪'�Գ92>��A�8S�ўX��ӹ d��/��Do��!�&H�C䉅I�"�Yp�Q+�		���n�L��ē�0|��\210�K.1�}���]�<A��-x��#a%ΦKn�ȹVnڦ��?�	�w(�1��玨��raJ� 3�!���O}��� ?&��]�t���J���FQ��Bx��Yw��#h�"��r��0%*��'�"��ɟ��?%>yQ���p�^Q 4�A)R�A�3� D�� �@�3|�Q2eC{1�wJ�O�9�K>�'���`�l���؅��G�Q5`4��v���!œ��Mc�'�V��S!887��0�cF�?�:���Ohl��'܉'f#|jDiĤb-Dx�f ��a6�p��'��	�b
�rL�gc�f�����<��O�O�g�<A����Щ8�6ɚQ,
eI�b�hG{��䯌,^Q.a�q@�}��qN�<����'5.��6�ƻ�fLaGn=c�2-S��HOn�����W�V�Ql��1����$"O�p�a!	5~�tԡU��3��	H�V������aI�AW9�4�b�Ї&>�B�ɪ���� U�F���f��,~D�B�	���-;�*�P����0�]�lB�	?|��i !!м{����w�Ș<_jB�	���pp���gôx`OH�WLPB�	�b�JT(\��|�vN���B�ɗ@�NI��H�HU,��ek�h�jC�	 ���@K��=��`�-Q���C�ɼCshdk�Cb���`p��&~o*C�I5fM��Bt�п�~Q�&5|JB�I3^2b��V(�u�ݢ -H-Z�&B䉻Yg0Yi�E�7ya1JŴb2C�I1B��P2R�֚?��+��B�W�C䉤KH=�����z
����8f�C�)� J���`�L�|h�-f�$��4"O.�#���r�U1q�@]��B"O�0*RFN�D_�Xzk��vOR���"O�8cAhԀ-ZA
� �
5^X�"O��Y���j�:���J���X�"O�4A�lx깸Cʖ6�\"O>}3�!U�x����L��|Rw"O4�n��xE��+DN\�]��3D���F�8J����n��?DtaD0D�hA���,w���P%�[�(��)ۇ -D�X��' �.I26^����3�-D��36OԉJ�p�B"�]:d��iP��'D��@���#�]�q���h��%D���m�i�jqxq���kR�YDe/D�X��-^)=l�Q��K��1*-D�ذ���8ITP���4x��e5D�p	S��՚�@.''H��8D�;��]:��E�T�8�R�G�5D������%sFf�H�Ԓe��9Ya� D��q�HE!)�h8�Pc�	?��=bX�!�d�u���0A�)"�iboģ%�!�D�=u�z%���84����}�!�Dَ3+Z�26L-Т5.ƧC�!�I�iRg�b�HD�=a�!�dǌ-�|y@�Ҙ� �"�I�!��Q�L�1$G�4��	P%@�;n!�پ3��p��*���>|�֮�*@!�dϱJz^�wG���P��l:!�d�?=��58�����I�M�� R!�� <w��m���V)�]2�FN�0�!����&�` B<m!��`�(k�!� ,��9� qa��y�"j�!�d o|Y�/�sH(��L� B!�W�q��P@�#V�����%Pt.!�E��$Z"��!��<����?!�DZ<��9Ȕ瓱~�JW���j�!��O���hD��7r�����R�!�d� YVʥ�fR.C��t�P���!�ĕ+p�����Q1ܮygJ��9s!�$_>{��@2��	7$��IC�(�!�$��R ��3/bs��V��!�$a_U��E"���F�$�!�.�d8���T�L	@�@�@u�!�ĝ�Z�E1����Ph$�
!6!�$�Wr�2�ܐ`|,4QN	3p�!���F���:l(N�F��#ϗE�!�$E{�p�%S�[(1�b!�!�䐅Qx��H`�:`��@��!�d �:TƝ��N�N�x�;"W�!��N6G�\9���4n+���A@�,!�$��X!��N13ZI�4���Py�Hۊ�X��F�
��&����X�yriR#YD~�'�Խg�]�`/�2�y2�qoČ�5��w��I�WH^�yr�C�c�� F'ӶlWv�R@�N��yb(1x��m�G-�`&�I�ú�yrI5=��p���o�: �.�y��K�����p�V4�NE;�%�y��Ǿ���"-��/OX$��3�y�#�E��Q1��[=ZQ��t��!�y��-T谱��EU�Di���Q9�y��a6�r�mڣ}�n��Df��ybM�#-��=�!��>���J�a��y��Ƶv�0;"H�6@�j �0��/�y
� b�m�"�P9��R�>\nU�g"O�L3b�I	2B�Cݦ*f��a	�'���R���Yk�!q"�2W�yB�'����&�6s��Hj�._�2���	�'�� 0�r��}��T&$�����'������t��5(b� ��lb�'>"��pL�&a��	s��0@��8	�'b�Q��7�D�I���1fL�K��M:�Y�ṟ��X�=)`B%"OJ�ٔ�#�D���έl��6"O�y�"b�{e@���5b���"O��+N$jC@�(H�bB"O慘�g�/+t荃F��e��(�"O�-�s"�0	Ӡ��A�̅+�r�"O����#�%'ЙɓĄ.�����"O�2���dQ'�^�(�P��"O>T8�f$C��֌�/L��"�"O���te�g�|�� 솖GA��y�"Oj�X` -[1�Q$ʜ>�֠)�"O,2��$������E��d"O�UYp��3\���p!B^K."��V"O<(���������ǁ8��9�"O�QRe�&��u�ġ=I�(��"OnhV�*��ܡ���.&Xp;�"O��񪎬&s6O�7r�H �"O���#!��T8���nM�p�<���"O�(ذF�h;��t/�:Ah �"O��S����-m͋3&6���"O�ȡ�5T��
j��G"O�Dᤆ��U*���V�R�lR�"O��aЎF��"����*�<�u"O��#'EP/@o�e�&��=u�i"O�[�hAj���g�'n�؋F"Ohw��}�D<��dب���"OL]�G���idp#�b޴3��8�"Oi�
�uf6�;c�^<C�"O�D�de�&�p�����N�Ȝ��"O�<r� �Fi�����90��HЄ�*|O~��TME� ����B�Y)ƨ�E�i�ў"~n��eB��)E(�Xx��A�b�PB�I�H4�$�W�H6t�Q7�^�"`�C�IP�t����Z~�`��e�~-�C�ɴu�qqNX�~]p�醇N�o�>C䉓r�`Ts4�-R\���$͔4�VB��hF@"3ΛJ�ࠂ3��=L,B�	�\�U �z��+`��.��C䉝
r	h�hJ�@��§̒��C�	�6(p�#e��y4�[`(�)��C�.>Ө��	R�~���Y��-D<C�I�`��Y3��3Nq�J��T*;��B䉲s8�1�u���C����`�S���B�ɓh���%�R�\A�L���<m�B�	
qdY�eA�,
<�$��'CNC�I��PmA0��$>��� ��LB�I�oQZ@��
�� ���ȁ�<i�B�	�"^��PA
JK���W� �*ٺB�I	Qu�A� @/E���������B�	�HX��p�j�?��&��Wz�B�	�%0�)����J�s�$c�pB�I�Ul�
*#f�P)�#aJB�IA[HD8��I8EP����l
B�(�"�I�!_�T6*A�)W#a<B��pu�f �`�X�(��U�XB�='��x����O�@�6dT�|��C�)� �3��
%��v��1�;�"O>��c�9���%	�j�\��"O�)�*@{��QRAJ�m���Q"O2 ��	EO2��d(M��шU"O�ŚPO�d����P'̵jK�;�y�fD�$�y���1P49�wJ��yb*�������+C�4O&�x����yRG8b���^>!�H�J��T��ycϵJ|d��4�A�I�:�B�eK��y�H�8>�r�za��i�pup+�&�y�'a̲���[���3�i�y2b��x�3�E۝'T�\xq�Z?�yO:�d ���.*���h����yR�E�h+�TQ��5�� � ���yb�Y5�t�jG�T�|� �����'~ў�Olp��S&QF� �
5D�}�y��'p���Q�J����W$ި]	�'���Pуߞd@���@�1k�8b�'6ؑ�2ƕ�~�YDM�yLl��'����%�F�Ӵ��J����X��'�!�q�� B��hbe�pL�q�
�'��a���Lyt�1vE�s��,��'�HH��\�꘍{e���
�'� �"���L j�&W ��!TU�<	6�L+cz�GdͿN	��Y�<���71l�H����9@���hz�<��!��k_�(x�/:d��#�x�<��J.�C#-+�1H��x�<�'�N�5��A�$��N��crɉx�<����3QH�۵N�+E��#�aLt�<)�K�)R$��@oA$S�ʩ�P�r�<��B���l���!����5@[m�<yG�C.3v)+cLȢtt�!A/Xg�<���4l�A`!U�L3:A` !E_�<��eְo�<���_z;����W�<q�&\CHz�s����\]6�:�R���hO�'\�Ra��C��("��#�Ʉȓ'M,�
Bb��&7>�(e�( F���)��2�@�PNZĘ���a�6B�	9�����.��(�A�mF�9�B�Z���@'蕪SE�8�섀z�B�	3_ܨ�%�w^�����͗[\�B�	�P!�m�"
��a��׬?�B�ɐ���KDU�3��b��ր{Y�B�	�)��lBDC� �@X`G,�".�B�1"T�X�a�C�F���+Ѭ��ƈC�	=8v��B�Z����g�.ҺC�I�o�z�	hKp	P�*&fB�9`l�-1#�+n�N�����/<	.B�I&=�Q"ό�	�pBY76BB�IO�B�\�e�:E`��W�(�:C�I��[���j�#e�T4P��B�I�G�����JS���C���C�	�6<�ٸ1����\T�3G�7E� C�ɛ@���Ο݊mjՏ��m��B��-M��yCƐzf]P����WO C�I�:H�N�N	0�+�׿u� B�	7T��5�sK�G��X��T��(C䉭(l�Q�6k�C���1���+�B�	�P_��a�E�0L=�`I����B�I�]��X������,޺=�>���'����� E�Z��\)��F%i���'O�@[!��L:vD�ԋ �(�F(x	�'{*y��%ۿT�� ��)�̾�x��� T��
E���"jΗ��$9W"O֭�'�?����A�|Lv�1�"O��%�O�O�Q��۹BG�c�"O��`SGP�@(b%�$C�%a�"O�х�@.>���@ea��dx�h��� �����x�!�w���������� ~Ӳ��wEu*L���E�t�����Q��m�E�@'z��ȓ5
��0�����pg�@�`�Q�ȓa�l�u�U;[�f�h$�� ����Zk2�a!ÓB6���ˋ��|���j��\���N��(��*�zI.̆ȓp)ȡ) l����y��ȓc�,p*5`d��zB�dhdD�ȓC��|�#�	r�r݉���RE�ȓwj�8"4́
 J�l9��G�/U��ȓT�x��0D��:��5��6!Ҿ ��5g|W�qd$a��#���
�"O��+�r��Љ�	���]rr"Oz���-�\JR�Z���T�*� g"O�`� ����	�V��}Ql��"O�0�Td��y#@� 7�2H�8�"OZ��o��o���3礊�(H5�b"O6�A�`ҢZdHa0��/?!�0�5"O, �T�'����C�W�\���"O��!D�;m$��r ���
J	��"ODD�P�̭w(�ճ!/G�i�`�4"Oȭ�@ �=3�5��ㄐ0ێu�Q"O*Uh3*��{�b�wC��&%	&"O�y��m���P�!W
*�Btٖ"O�mC≑8u2δ�2N�/
�$��"OV�	eY�	&���!���w��ڷ"OJ�렫;u���E9�ؙ"O��j0F��2�	%�\S�*��%"O���!��m� J��o�ܴ!"O�	j�-VRƜ8���2��4�"O�Y��L�m&}�'�ɀ�"O¹;��2)��,CÇ�8~�|4�g���<L1�K�.0��u�g�ؙ9��'J�����-&� ����F��)��'�fD�w�$t��P	C
8,�ʜ	�'�Fp���_q���r�}$�r�'0p�b'-�A�\�ɢa��)�'tz��j�:Z6��b�:&Q|��'���arFj;���/�/-ѐ�0�'	D���ES�g4�\V
�0�90�'\�0(fi,#��D��-/ڄR�'�҅�3ŕ+:M���3�z'�4�
�'���g�-#٦S��	9#���	�'ޑc��^�b�|���(�#9�i	�'�2)i�-�Ƅa��kO�1�"OD���$X�a�"�Q�k�I'D��u"O�89�#S&Lѹ
)F2m)&"O�����>ژi2�i�W'f�*�"O�"�̋	��=�V錪6�V"O��;󧝱,A�E�wIX%��A`"O�	Z�VDK�K�w��5��"O\���(��BKN� 憐�^����"OZ�#����HY(����22����"O.be��"���Ir(�	�$\ʩ`��
��\��-�8s�� ��M��p��eT���x�Bk�q�v��.T�x�H-��' �r�ϰ��I�Z��q�p����S�By�����}i"OB��@��`�b8pA+�JW�* nD=P��)6�����@�d��Q>˓/�% ���
7Ξ�6!�Q5����S�? �=���Nq�f!�4�0<�V;��]
��17�V�.-���C�:��O�0�5���c,0A0�ȝ:��X���'-4I(P#�8��@��N2_Ɣ�*e&�-<��my���� ��e͉*Sd6܆�	������W�
�D0�ɝq$O؁p��]'~4�'�t)�V�F�e�
��~&����x�<YҬV*nI�\��l,J ��Ɓcܓ%��c��1����¿@z�8bt挗;�h$��d�>i���ߠ<k0��@��Ce\�VmE	Z��ʵfS��Oޢ}�3����ghT
90�A%"4O5�p#2�	�n��zFH�sV�T�a[2b`r�(f&����ɺe��d8�F�;1��<0@i�����w`4Q��O
\��T�ػ�ə""`�Mِ�6q�fiQ�@;D��+W��(/��$�2��=>df�6�;�=?gn��� =�쫗�@�n-nLn\)�����@y %,����������4G_%w��p�'��y���p�(4ia눖Kz���� �k�r�ٍ,�<,(�* q�y��ᑖ�y�7=�X=²D�`���5A���$IX��"|�5��-$�%�)%����Ƣ@�<�u�ߵp�f�Q,!Zg�%�ANJ�[d�1�	�J�	�G����Q�Å��,����I���B��x�����@�Ҁ�D�Ƭ��xbb�PYd�rΚ	J$�X�2��0<��ؕ��'o�YISA��U�����Z"
"<��'�Гb��$�P��P`̅��O��g �)§HӖ�T�B�a*9S�F$(�F̆�IA�5����f�;.5�ǩ��C@��ȓd��s��):�ɱu�ӗy"�)�=1�����ό�c��g��g��@S�iߡ�y��F�E4pm�A�gv���6��2�(O:��d��Sn�T�4��-�`�8��[9�!�d$]X8DiËm��}����ƕ�ē~?<�F^�@r��Bw,Ñs�.����\�U�\���@�+c>�i#�H�=�<��}�%�J�b{V䂁�tՅȓp��d��=� ��	�8{�4���h��Q� G��udb�b3o@�KV<��>�L��(V�2B�br덌S��5�ȓOn��x2+E
#����N8�(�ȓrP�,L�{߈,!IuV�ل���e	��:�B�*%�H�݄�WB�<�d��+e����c���p�h��ȓh�$�`�-�0��\�j����
��Xq�C�-I��ɪ��%��ȓ��H�M��/�xI"&㉪Il�1�ȓ[?~� �BU���E�ՠY�T�ȓ�8|J�k�@��5/ �����o�3a���
ó��>y8^d��p�&�B���\+��F��(�\(��N��p�Wb�	rh{� �+k�6��ȓ;�)z��;c���� a��"T|��w4��t�]�"{�|��]!S�z���H��u3�[�H���K�E����|Z��;b�1��⇑�y~�)�ȓa��V��G�-���	#G�P�ȓR�މk�P�_Y^؊�LP@��ȓ��X���C.�h��c�ש��4��]���%b���U��3 ���?W��Vg�dДjw���:�܆ȓ}f�EB�#��|I�@� �J	�<a���NQc��%-�&Ł���
T�촆ȓ_?�����
r�E�vO@8�y�ȓv[�yQl��O3@�+�À�^F�ȓ*�Ղ���)_$��;�NF�V�`T��S�? �}C���3qh���=��b&"Ov|�ƂY�P�c�"O^�0!"OV5�`n�2p}��J�%șe���"O�� �t�� i�Z�l���"���6{xN���<�>	�)X9G����w�Y'0y�$��	"=�8Cqi�)!Hs��S8��-��+��� �� �'s(e
�懜kC"�(���DB�����Ӑ5;�H3B�D�T��O�6}���X#E&����Ml�E��'q�	9sJ�|1ЇD�;��'{��A�D�'�H�!��p>�/M<Θ�tƇ�K����:�!�DM;sK� 1%&A=&���V [1!�ؤ+��O~��n�К)aO?�d�b�/�
T02��?R��)��?�O�ӱ�ۗwb��s���8��YY�#H�[��!cuN�#&�c m=�OP��ʆ�O"�3"�2V���#�Ƀ�V��P)"L��`��BX�ԇA�Q�f ���Q��\(&�yr�CK�v�re)U��0��h��yb�T�6l9E(ϑk��4�U��`��X1��C�q�A��6��q �'־m�eQ�,t���JPy��� ��7\�!W�?�������	n�0�1 ��P$zJ�H�eL�"[W8���	-*V��(��N�N�zზ?Y�����J/g�̀D�U);n���hO�O���P�śe�v�S�K�h�V�����3��(��{�nQ�"-�|*�/å?��I��KÚ>�����w�'Aay�^��x�����6-�V���Z��y��)�H�2*ԃ��j���k�up����p\�E�C"�~���'idYU����UiD�G|���a���A�pM"���8L�O��Ox�R��.~���C�M��:��'��!�a��i�A����4AJp[%f��w
L�& _9�lL���hO�O�����%��{S����򉠈�D��*9Y���K^^�OE���f��F[�[ray��p0��+,O�-�q�5u��@{��A�	���Z��*#�	+� �/��)ʧu���1n1h���i��Ӝ�"O.%h���O�H���?԰ȸ����kZ`���r�L�a#�(p�hT�Ŷ\����<���a�O�oN ���h�:Upfц� z���vH45>݋p�5Fʉ�ȓpF�ps%ՂR�:�S3�Z0!85�ȓo��4ĆU;-PJ��'	ı/em���y��`��{K�	��/4����&l 0itf�&4ݲ&"P����z��)!�$V����C�	�fmF�����EȤn�*�&�JTl��)�F��ȓu�^�i�bMgs<�HA�"$x����f��'\m�hPh'	H�K��E�ȓH�� Bj˿TWΜ�#�C�J��j[D�w�L0�P��c�'���ȓ~U�Ъ�`y�t��#�:/�I��.Xp��s���%)�D�a��ȓB^	�%��$.�X�����f	��ȓ8:~�0�
:�v��'�W�%:�>�%�I��p<�f	Bcw����dy�JAr֊b(<�TAE�\��VE	���vI�
<8��I��%�L�2̂�49:�"ܻS�Ap/+OL��T��
�'�T�T��zHd
! �7�L�c
�'��0���ĝ7H��˔� �g��ɸI���'���1�qO���f$]�glL��UT7R����"O��E��`n°dk��`�!�26�XQ��'��������E-\�c7GG�>�z�x�'�d�
6j�kN�I�޷U� E�:c��%��(ЙSR�J1 ?U�%B&Uf� ��	cx �=�6�X�1�D�͗�Z�ܡA �T�<��n�$F��� !�3�p�KI�<��n��CJ����ġl "O�5��ɂ.,l�9����W���C"Oy�ԫ�C!m83�Y9�n�I"O� � 1��C�#�>��1�LP	�)�"O&m֜O�|����-xx�"O�Q�v�)e�:�D��cg�}cv"ODu�cQ�Q �e�%��X�C"O��y-mA`|�&�Ĵ@��Ȋ7"Op�0B����v��C�(�ܩ��"Ol�
Dk�7��(!�\�
�H=W"O��A�
<�X�b��T�lI�"O.�:��,��:G�Q60�H˲OL�B��d���Acj�Eu|�	aD)u!�J�1werlM���|�b
Y�3�ayĘ`c�Cb��'Sd�x�3����F.0�əA�N��$Qa�xm�
ɖb�<r���y�͘+<|���Ж
��8j��T������P��1ؾq��G*؇��WH�ȓ 8@Ѩ��9ݘ�j� ��}�ZЄ�*��a�f;RB�!�ׁ�
7,���wx&���+�<m�:8�taL�o�݆�=On(ʓ��
cK��qQ#8qQ����}�����Og"tၓǎ�$��X��j:��Ƌ��9:�)w�U'�8�ȓ]*�)�(ܿS�H�!�Nѷnc���H��␵/�(q��Y���ȓQ&��@���y>h�P��A��M��&���9@�G�1�`���'A�js�ل�((�)�#\>!L ��y�*1��Q�H
�$ ��l��A!�2���P����׮:��*@�>g�P�ȓz�D(K��ԕK n�ا#BS�$m�ȓk���+�F��/ ����I�<  ȇȓ	��N!j4
იt�PH��U.�EX�b�ޤ�G�|Y��s����Q#FxaRG�� �0�ȓiPI¦�U�����3=Un0��&&��d�N�]� �Wd�c�ن�G��5�Q:7����LYn�ȓ6��Sď/j���Q\�q�ȓ�(��L�!{0Tb�m�Q?8��`����������u��;�୆����Pt@�8�|a��o�8@���ȓ)�@�����@��]jQ,Q�x>�x�ȓ<�B1�D��	:A�-�R��1>цȓc"p���N$2�V���㉙N:���ȓ^f֭ �I;/�]!կ�� ���iz��Bf�G�Mi�ظ��^�R�����[]!�t+[!;(�$VK
�Q\���ȓ"Y��Q҈��K��}9��3Ku2��ȓB�Ǐ�
�Q� ͕3[��D�ȓ$^RuJ�5zj�`��P�����ȓ4�֍`�iD�Վ `f�M$"�h��zlpKÉ�!�Աy@(�(\� �ȓ!��@�mE_	> �R��'Sx��ȓI+D{��2R�#sY���ȓq-t}����y��V�<ze�ȓ������ ���ɘ$p�l��!��@�O�$�0�#���-Osƨ��f���a�ƕE(�E���@�����-:�q����yK�c�1֪��4��!�C<��UG�@}0���dO�]*�@̷w߬%�,��0̇�n�l��5��%5�*m!F%�Dj*H����]k�@-J2�!Q�l�>cZm��3�`H��i�5^�1��
K�R��ȓ\��Ȧ�@�f"��B��0x���S�? ڐ�`�Cy���)����#�b���"O�����)3�� !�N�%-9It"OZ���K�K	�h�v��-R�D 2T"O� �qϐ�\�ĕ��+���Hv"O�0uN�d����H�y��3C"O�=��єQg|���W�vL#&"O�����90�! g޴O֨"�"O����$̪:��k��ĩ�����"Oؖ>|}n�*���&!�vQ�v�V��y�G�Y��0�)#h�j��N�y�N'?��@�!�K�����(%�yB��X*����:ř�&���y��ɓ)�d�P�G=�I�4i���y2B�!s�dJ!��,hRhPH$-���yF��A�p��3�-V�.x�d���y�'�52���S"O�@5����y�OJ�|�iL�`��-_��y���H>"����ָ�e��y�-��L��C%�jD�P(��y�.O�tUZ�r������+'�y�C�JUj��K*4���F���y���+�4��'R��r�[&��y2��,k}�5���L����$�yR��#ΒA�����zg �TK_��y�nP<
f�4+bޟg	p= �/7�y� GwƱ����R6�0����y��Щ'� ��&`\$F�����ĭ�y���=h��Ic�O�?������6�y"A܈~*�E���H�`Ɋ������y��T�����;QJH�O��yrh[
Z��v$�"I�̙���D5�y��F�D��k6)Q/G�*ii��.�yRA�#�
3͍0![>BU��yB����D����Bm���Q�)��y�e �5xl��C�J5���y"iߙ{O��ߔC&=8%b��y�ۮa�nSO�72��D
L�yҠ��~H���E��|G�G,�yr�� �z1���ܾ	��)���y"��9~4�����	��@z� [�y�'E=lx�X��  
���E	\��yR.�2CG�����^lX�X!����֤e���˝L�p�"�TpH��5;qV��]5�	�̒�mP�<��f��+��x༺��X(N�9�ȓ8>���
*^�"��3�H��ȓu�@�j�Õ0��H�w�^��n���L����MK-\̸Armݮs���ȓ|͚`H5��,?w��i����U5���ȓ)��%ЀꕬL�N	��K҅ �D�ȓr��򮇦hҘ���$�݄ȓZ����$R���[5�Gvfe��d������G��iUjef�ȓ+�����[(
�!��)�ƅ�ȓIܲ�	Ԯ�8�f� �NWiQ0y�ȓ^��y����sh:�hb�֎vD ��.�RMH���O�d��4����D���jiѶ�׍3���LX	�b��ȓ&���χP��Ēa#�oq>��ȓ=v}��IC �]!$ٺ.0ⱆȓRT*��B�A����Ѝ5�t��(Z�q35��� ���!�2Fs*	��_
��1B���:�F��O.�b�ȓW
>�:t9p-�����W�d�\@��S�? ����*L�j���+Z�hhA"O,Qj��*�r���̋�
�S"O�h�k�]�P<�D�%��$
�"O�Q����}���Ę����e"O&� B&C� �RdϞl�tP�"OzPj'�GPT�͹1HԒ�)�"O���O�(cX�UH�$V��I�"O�X�H�_}����C�g�$C"O��h!�H�w8����8p����"O�d)��Exv�֏Ã'�D8�%"O�����8Q����S���(U8�"O�2�Ō+#�t����~h�\��"OFI���Z�x(d��5S*��F"O�FcF$`|�T.-\㨼B""O^Pá��n���.A�_��`��"OT���C�:.��0v�^�4ݸ�"O��!�@�#���c�5ҕ�1"O�L��ܱYB��  �ٞ!)�"O؄zW�C�
�V��V ��{��U��"O��IŶf�Τ�r�A�)��q)�"OT��1�O!\>м`a'V<F݄a�c"OJ�c�#ܼ9	L98B��)��钦"OD�
!d��,7��딅���,��"OмF̒�z.��P��J�G��X�"O�Г��J�+���)�B��S�V"O�e��9!�u����xGƨ"��!D��q`
$G����p�HG��T'"D�dZ&
p���@��[(^��1у?D�Xzrb�+�~�A�V�BP�<(.;D�x�է��>��a�/��bL��D8D�@
0,��H�H��`�7WWj�ѐ�%D�I��>F h0���C��8�QM!D�l�"��3>@�((��lSި� !3D�����h�Z̪�ĠX�lAF�'D��+c(1Y��\Tc��82��k5�$D�0s��O=}��8h�H�vx�T��7D��6��=����-��T�r��F)D�h�s�4��uЧ�Jz�x$�c�-D��(e�X�U!&�U=^= ��O=D��P�ʴ8�� ���BQnlH�G6T�((鐆:5�`��oT�(���U"O�L"`%�BV�鴮�t��� "O�(08n���	�#��`�Z�	�"O �ҁN��]��y�&#�8u�$"O�-�f��&�|0�A��6���"�"O(��q�?���{$-(��`��"O�� w.I�!U�,��f��6]��"O�e1&�
qZ,�%^�2����7"OZU���Z�5���D�O�y�G"O� 	���Y��d�����n�ԣ"Ot�f�J=@h-���T�-�  ��"Olb�H�Q�(s�C�"G�J��q"O�Hy � Q�m�#��99�,�3"O�Y`"�I�6���"/�V"Oژ9��CKIz��P�O�@�0�"�"O�9�@/{���7�+�f1�"O((���dKИu^h���*"O�i5k�t�����/�B�(tu"O�%����\�#�.n�y("OR`C��k#�"�")NH��"O@�`r����r�5/�/;h�"�"OX�[s�K�v"� �΅�%6�kq"ON@u"��6����Pn@� ��T[�"O,P��jԻ���B��ej�+�"O� �X3�C��Nh�M�`�V�]G��a�"O��Q�L{,A6H�R!�)�"O&��E�	68W:݈e�����8�"O�e���Z��$Y�_��nx "O��eB�"r����'�@���"O�%8 l��Z@qQT's��YP�"Of�
r��ƾ�u@��((R"O@p
�03?:�����;�z�YU"O$�J��F�~ۖTڃ�Ѣn��s�"O�Y� �@sdB�i�ꂴKքRE"Ozm9�E	1�0(�s�!#�N���"O�H��L0�J5��m��@E"O�]��X	P��P��*"�VJ�"O�Z� �.����#��:o�U��"O>�"�	z��Aat�=5Y�"OZ��w!O�b͆l�3"L�Ti��I"O����qb��s+¤\N��24"Oέ"BJ~$l@'j� :O
G"O�M�6�\6����*�+?&$��"O�h�5"Q2i)��X�r�@"K��y�ɻ'�������.}��8AS��y�
Q/wZ��v��kc�@Pck
6�yB�N�pa��&�a�@������y2��*GVPT�Lv�`:���y�7y��a �k�F��ѐl��y��֝m��cuƟ�%)�\Y�'���y�,XU�$�ئA x^�1w� ��y���6�2	�D-M�o��&ꜣ�y�[=h&3���,j��˧�y"O/S�]X׮��y�R��#���y�-�zhM����~ʞ��g�ϧ�y�ə1���U�J< ��P9�έ�y�k�	9�z%��v��%�A7�y"l�
ezu��Ƒ�δT�D_-�y�_q=ޙ�+�]�����>�y2��_�d$�T�H��^	Kb@_7�y"@T1W��x�ѮC�z�J$�q��zB�I�^���PK
5O|���E(M�XB�	�!8�I$&۱R�k�D�)�C�ɭ`�"ɀ@�$'�`�
\�1��C�	�1��)�q�YG;�����^77{@C䉰hs���ӜuR�Q�$B]�W�C�I��V��c�0y;Pi�6�P���U&BĉCLѦB�"&e����)�ȓN��=�����Н���0jju��4�lHU@��i��*�V�T�=qe�ʨ{4����)}rq�HL�	�Ey��G(� 8��Pz�C�Jg�C�I�4Ȱ�[+m��XQ�]0#�ʓl��{se�wx��
M�		�}��LĕZQ�Wz8��ƧE.!in�a�d<����0|�f�U�ʨ83)�;��+��[�uň���J|��B+F:
o�L��m�a^s≦4�l��?�~����O�рIȜy�=S�b][}�ȆLC�O�>!���H5u @�ddG���0�j���6�.�)�r �xp�`��Ĝ�R-��3@�0!@.�I��0|2F텸9�\�3��%=�<SÑx�#�V�x�J|�����`|��t,�:V��ES�!v�	*u�"��?�~rV"��z��i��5���j �r}�lK(F�O�>�RE��z9Ԉ�/8}��hԷ` B'9��O�?Ue�K�U�(H�!��H��5Q�O����|h�Q��.}�t���\c�p	L�@�S�Ӣ}�̜ˣN4�N�
e��bvOd���$�)z�'Wj��T�rHU ĨH�?���OƔ�P�"�)ҧi ӬU�8t�X��A�#=�LQl�"e���?E��	&�����K��,!$�ОPP�?��π Tyc�fm
�Ap�^�h��i�CehX���`a�ĪgNa#*G5�zL0T�x�fk�O����S�	�z-3 		X��t
�_�Hp�K�A�S�Oq�1��i޿z�>��#�� �)ܴf�2��G����'l�����!w��q�`G�H�!�#T
h5bSF��5D�(�n��W�!�d]"6}�jŉ��!�P �6S�x�!���xR�E� ӢA��A]Uw!�Z�v�s�0�Αq@��9H!��/�u�d$Y��X�bqHU6;!��E&9�n�I�0�͉$g@606!���0��T)d(�U�z	`tfۂ<)!��T����L��H�Ϙ�&!�$E(`:��u&V��*C5N���!�d��n1:�
�)���JG����!��a�u
�US��W��!��oy��`!D
W4��,Y�e�!��ʝR�f����n�V����!f!�D�A��5:�nD�<�앐#ꚵ?d!��O�h[B�yÐ 0��!�DHH��Ua���Z
Mh`�^�y!�֗X�ڍ�B�P��.ș�lʽ!�d��CFAЃ�7?�Z�� M?[!���&|�V�	�ė! �rU�!򤐑}ئ��2�G*;�4�K���2T!�D$U\p�+L��l ��սlZ!�d���0Ʉ�A����� 擖R!�B�L;0���([2Q6�1I!�ױK!�d�R�q�"e_�M n؂�K�m�!�E�n��Ƀ�n�5R��`ʒ</�!�ɢ>�"ȓ�,(�����
5�!�$D�
�F:ԎA/h�����B�m�!��R4AIR&H*v�����n�!�d2z�u��v����T`-�!��=��Y��� 8u$�[��O�y�!�ċ	D�h`5gD��q`��!���>!^H*$J
�w}¦$�2\v!����n�0������j�C��JI!�$S/r��c�G�R����#!
6!�D]�.�l�ҩ]:|��Y1��d&!�D�5�HI��A�zv���J�/d4!�dW�xDj�{6��ud��"�	3�!�$E!���2��E�Kti� G�!�$�,ql�y�A!����(��n��!�d�*	N �S�σ,���q���!��t?8�*�`#F0b�J3(�5/�!�dW�N�����-Ԉy:g�'w�!��Zsl2�N�l�*�sq�Z0R!���y��А��:u�(e�Gk��!�$�M���i$k�P�K�JE1Q !�ի��I/t�j�:f*���p@"O��e�4�Jq�D˨g�2I R"O�-�`�߽~�h��ň����à"O@�Qg+�0(R��ʆ�&!��G"OFػw��=�Ma��ۑx�켳$"O��Xd62�����KG�X�z"O�P`��9	z=p&'��`����P"O<Ԛ1
I%e�FE��g܇`��f"O���( %�XvEX�Hx"OX ����;m�u�!���p�6"O0dAW��'j?l�",[�<���"O(�闈�(=�<��!?1jb�"O��[hT�BKN�<�d�ƁH.5'!���S.̼k$�K�)����뇵Q�!�� ���aF�!D��M��	�'I��A6"O>����:u:̋s��'��x�'"OP<B7-Q
cP$�cC`�-��8 U"O2��V�h�ܡȲ���5u��[�"O�	��,%���x�`\�2|��""O�(��ŮYv���Z-{� �f"O�����3����pͅ c �(�"O*�У�D�o��� ���^��"O(I�1�إk�䠢	�'��� "OYKpHN�O�(|��GG�W~�x�f"O�� pFF�-I�Ē%�	-_���"O�`4Wj,v�*&�ۺoa(�H�"O��2s��$R�<(��aCCNt�p"O
e�f 2.{��rA�3]�) "O��8/�A_.���]�@��@Q"O��j"(�R�>ő��0/9�%"OH�� .D"����t�H�R���H�"O�8�@$E5Qj`bt�[���`�"O:d��EN��8l�ӋH`tX�U"O�!AbC�jBzH�SK�*jnDAf"Oy�c�l>f���jX<;Z���"O����wO ������\Dx���"O��6�A)$��P����$R>|9��"O����ߦ$V�e9Ǡ^8@��"O�-�I��-~}�D �N��"OHH�i�� P�\:���h:�ԓA"O����ƍ�W>B���7 ˺qi�"Or4�u��`f�L�'�]	r�f��"O��Eĉ�v�s'c��k���v"Oh���F2w"��waߙ=f.؉ "O�e��F[V �@��3d �#"OnU� o׶�er��.v:V�i�"OB�jS V�#���)Vˏ�+�S"O$a��FΕ(�:@j"E ���"O�<t���X%S���G��2"O����[�t�0M�!̦&���"O,����'(: TB���#|��J%"O�h��Z�c�����DF {X��"O�E�%x�2U)u*�!^m+�&�yr)H6Y1�i�Ǚ.%d��r��yƍ�!�L]XCpIXs�3)�Їȓ$�>�9��	0Ad}�`�]�a�ȓ{N���&�i���Th'�����RH_�ah ԛS�6QEp݄�.<�eB�8�ΕS��4|[�h���n�Ǩ�<RЌsQn�-��ȓCV�C6��Y�2%��eS?)&��ȓ>��es��
	q?r`�ÏjG��ȓ)��L�¡S�
O��C$��?��D�ȓS������ͳGJ2ખ�DXL�̄ȓ5'�AQ)�:|P4ɵo��?t$Dx��'���(WnU��$��P�C�|��1"�'*��I@Q�LV8�@Z�s!�a�
�'R�P��A3H0D)z���ThPq
�'�
lf$
�+��,2G%X,#�5
�'�a`�	?eh���	�fuȚ�'�J����٣x/�P��[Hx�i�' [�)V�?��8��ˣO��e[	�'���Y��å��0��Yp��8�y�e2"���I���8�I����y�+)��S��J12J+�����yb�-Y�	��^>�����Ã�yR%�3�<�p
�&����n�ym�.X���䨙(�r��$�L��y
� N43��,R�(�S���#�~�IP"O���̗�E�肦hF'Fy�<p "O�� u�ݘ�V��T�SIq��T"O��S#H�|���ōxi�Q"Os�a��[c% "CM�K6"O�)����A�ɺgK�T�T"O(#��9��tم�%3<�}XG"O^ћ��T�G�N���\�J�(zp"O��"�X0,%���vϗ�\2p �D"O�(�FB�a���Ƞ))l��P"O0��Sr�R�y�%eTzc"O���҈U�A�����L��a
�̳�"Ox QG�D����mE{�p5��"ObdK��Gv`�"���n����@"Oj�BѦ�=h���Ō	w�4�d"O&���k�7{������ ~�	�G"O�\��n��5*0Г�E�<6i4���"Ox��mY�n�|��6�J�kPp��5"Ona�sm��qڥ���:OC����"O����d��)x.�y'���Y'Y8 "O�A�0(R x6��KQ��A�\@�"O��k�Aw�:бuCː�8"�"O.	0�_h���2m�(GRd�t"OS#G;2+�E���07���g"O�S�ܔs�D;W�
*�(�!"O2I�V`3c��H��yܲ�0�"O9�NLr�0l�6\�0iyt"O��`R��.�tQ&�ȧK�"���"O���D. �|��c�i
)��1�"ODl*hXQ`���II�:�PP�"O�p��A��`�*%O���!0"Ox!��)�1q���0�j$���C#"O.Œ�#�c�0l��I�� �`x�"O� ��U�>�HG(�rK����"OF���OhHd
e���9�� �"O���S�9�M�U��#�:�
�"OR���V��n�kDf7qR���"O�щ��Ăq��i�'��9d��"O(�S�hQ�5(��F�]1:(�	`�"O�X�{Ф���V�"	:�8p"O�-��bO��0���S*Et}Zg"O~�+��;��D� C�6^&1S�"O���K��Bo��P�ƣ6<@D"O&y�j�4N�w�N�pP���"O��kA`7X8�m�%��Q0"O�좰%ɕJ(���[D��Ȩ�"O��:���j����"��o1,0�g"O�$ C�qx Q�aaP��˓"OD���`� i�өU��@�"O"��2�f\鉤�H�p�$9��"OBq�A.M:S�XX���V;��,R""Of����ZHY��i"�C�"O�@�*�oO&u�"�P.i �t3S"OP�k@��Q�tjH�~w8x2"O�[A�� ���s�I�#i�,"OnyH����#�6�p��ס,P��'"O���C�3�4Q�G�R�gר]�"O޽#�`Ɉ+�6إ%M��jD�"O`@��c�,�t����Ȼ"Oި[祜;t8�Y�aJ.! �E��"O����[�{��P��e˱/�ظ��"O��5,E4:HL����`�.�Q�"O�4�1Z1
��$���DA���"O��1�9�HY�
��]>��5"O� ��3��ڸE�o�#���"OX�Ñ
���D؂�Yɳ"OȬ�FmK�iN���k-K��e�P"O$T��D�L���9���:��t2�"Or�A6kޑ1 ����g\.3���&"O8[S��R��M��%�'�>`C"O�`� \�
C�n�v�#`"O��V�	�U<�a��(hrQ "Ox�x�!Y�7�2� C�(sX��"O�!j#	�!m�� �R7LH�X�"O��o�R��I��a�l���O���S�_@���ݴ�?y�'��	
O:��"�T��h�`p0��՟���ٟd"�J�Kn,����o�:�!�gd��)>B\�a��O�p�y ��gK�YFy�aR>{hP�k.@k|�	�卶]8�ͻ� X��H����/}MZ�#`T8�n�mr�}6� �Ʉ�M�Ƕi�bS?e��BD�Qĺ�zg�0D]~)(�W�?������hCP�s��I����x�"I��'��7M���m���<�C�kg?zp0$����O��*U��M}b�'`�8O�L���Dm�+/��"dBC�t�F ���;@wN 2���Tn��b�*޲u*�4z.����I�]��S�?�1Y\n��bf�l�mPX��%4�i�@���`������4�^t�1M�#�8���N�����h�Y�断hFBx�7N�[a���t�iI������F�d����.�$��ܴ���򋙏/�Va�w,��;�����?QN>)���OX�ur��վt2p����R E��(O� mڎ�Mk�PO�6�';����dt���@%R�(�&Բ�VՉ�NF�� ��\�٣��۟��	֟(����u��'��VC�70DH�2@�f<��'T\j�n�8S,�s��v�4(�D���?���㎌H��O�]�T�U�L�.]�7�Z��ТԬ�=s�K�!%�X����Z�:�j���4�P���? h��o�c,��3Õ�.b�|	��I�M���x��'QQ��	S��ɀ,U+:��ukf�&}�)�Su����ω�P���P��B�dti��ix�7m4���|"/O��R�C!�nDا�@-!N0=��ܡs��PIo�O$�d�O��D]��~���OT��0D�a���MM��� ��K�<�c�bÔLdb/Ռo��W�&a*��P#�C��c��ل"�dYq ݪA�8��qm�<���'�G%`a�ק*�@��"�	�)R��ď%1N�!i����BIR�Qdģ�V��4�	P�S�t�]�P��y�ABA�JԼ�Z$	�y�ż4��y�flM/ZN��� ��>�~bdg�f�n�Ky򃞈Pf6m�O����~�"��*)�^8�B��Ҿ����B�)��d�b�'T2�'����q�C�����2�<&�p�St-Ϩ)�0�b��<眭���-m"d!�S"�*�(O�e/�:I96HA/f,,]��%��n��N�>m2U�1~��E t���:kФ�&����O`�nZ)�ħ�M��J�d�ҩ��B�-��Ip!\�Z'b��M}����{�a�^�qF���p>��iM�7�bӤ�uK�;��EFT��8�@�O.Y��%Nզ��I�ܕO�p���'�B�i� ["F"}e��Kr��$��U:�������F���$�d�!��>C���*!��J��'��XcoV����f�h��D�!	��4~L(0(��ش \Jأ�8"�8���%�1��>��P^ �[��Ș2d��c��-0�7�K�|��/`�Hl�ԟ�F�ܴj�\4�ņ�q��p��tc����?��鉝�Iw͎�.�"�o��&��<�U�i-�7�=���P֝t��<���ע�$y"��s���AK>��k,�e�  @�?�     B  �  �  :+  C6  >  UI  nR  �X  _  ee  �k  �q  -x  p~  ��  �  5�  ��  ɝ  �  O�  ��  Ҷ  �  e�  ,�  ��  j�  �  \�  ��  ��  �  G � z  Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�� |d��"O
`�(�;���8���-0��1%"Oj4��ND^[��"3/9�0|H�"OB���H��*�ʞRy=a"O�味V�!X��!&F�:J�$���"O,��a
���C�Ą�M�"O,$3%o�-���p���+Ն�:1"O��ݢ1����`���y14]2��i�<�6��{_���c�H�`�fX�$Kn�<��A̼VI�xR[�)�Ć�pඤ�ȓA5��('nߡ4�� �)˩%� ���,��r�؊b#`T�eT09���ȓ!�b��g��}�8�F��-? �ȓ
K|m�ș�VṔ���2�%�ȓ"R�X�j�4JN�1�˘X�i����̹	_�jZ��1!g��zܶ��ȓgil,*�J�
j�Ne��i�J%b���f	�(U��:���G��$Y^م�~r�� S�%T"���k\�jx�ȓ|4�1�îJb��@ӵ�ݩn�V��/[`�"�v4�R�!ʎ<��M�ȓ`:��z�ؚh�J�Z��$HY:	��H��p�m�C1��!��B:��0��EnjZA V;9����J[
2���	��4'J�EA�IVW&��~�(aZ��ӹ�>� o�Y�|�ȓ�f�A�
Ο7�H��M�$�����mޠP����/���ANXo*�ȓTv�����{ ��-7�*h��I��sB�8�8���3����ȓNe*M�悡;������X�o��!�ȓ'lj�#F�m�+R&;�|��2)n�C��0S4���T:
b���:�0!��e֊��)��ͷV��,�ȓ0�&�8#���� ع�L�����;�P�AFd���,w�6d��r�EQ�( �gVlɦ�M,H��,DP���|�I	$G#\���ȓ"�)���E�B	yt&B�^�LɅ�4�� ��eëF�ڙ��n��R�p�ȓp`@}bŇ�=�$�AUN��P����L��p���_�a�)�Y�!��-��u�5���o�`iF�@A�p �O�"<!����P>\�7��i1> �����}"��P�Um9���ȅ�J���a���O���+�S�O�"�nGv���Q�!؁wސ����(O���@^7+V�Eܒ��0����d}�D,�O�`0D�C+g��ԙ4�+(���p��'��O01���܆n�T8@�`1+��Y�"O�0	,�#?_��2���/S ,�"O,�rf��U�]B����:3��	U�'����y�#�RJDe������y؟��F�t�	�G���ᒏ���=��{B�X;:T�����@��J���<��d�O���h��Ĉ�91b��7d�(�x4���NL!�X��΍�aúi��	R&��2�!��
sd![�+e��e��`ƾ.�!���ߴm�r
����'�!�NV�8���E�g�u�ǕCxO��Ue�]�rQi��Ж"cZU�2"O����C�#L\�UAW'sZ�9�"O4��d��%+w1���ݬ��r�"O� ���A�������QC�n5��"On
�@��(�v�(�� ��9��Oh��F��'�	2t�NdH�<`�O�Y�<��'�AK���%%�`���\�ͺ���}bH5LO�<KF喽=�DҴBC+628���"O�I�d;*bp�@�k^�w�P;!"O��1���>�3va_Sx頧�	n>I�p�G�FQ���@e��_f�y'r�
�=E�ܴX��� �ESb�J�E匒_A`Fx��'�|�!�AҮ|=:ɢpm�-Ғ�c���x��T��i`/�|>`��!]-�y�*�wv�ѠM]�r�j��`�,�ybS0S�|U[���D������	A���Or\{b�}�n�҇%Ҵ,�F}R���:�Ұ�6
�� ���!�qO���䎺 2&����A�Q0��'A"O�a~�m�>9g���i��{� �i��廡�h�<	��6�B�JO�t,�"C�\��x�<1���.%��G͚2��IE�[X�<!Fǌ�WUB�c�kQ��`���S?��{���s�=ǰ]��4FCV�(3�9D�<"&�L%4�	�F;)�4�G�5D����7J`q�b�ٔ 1��/�p���'*�"t�C�*�l|��`�Jm��.%�<����!2 ipc�T���x�����q`�
R0D Є��E�%���L�� �9�
8��kۄ)�$%�������Qx����~00�dLH����\������
�
S2VZ�)� ��c��@3��&D��@�ΠZ��X�$,���p�n)D�x����?`�$���7r0� g(D�p�k���4��0kש�v}�EB%D�0�r(ø],�	aV�:jJٛrn#D��ҡ� #��L�UF��X%'D�8�E.� w�D�ögq� m�qf%�O��	�.�̸�eW4%�N��wI�4�B�	#Io��A�=�������W�:�	6��X���,�=�u$0Ӑ��e���s��0ă�<��iC�y
��<}mv�"R�PV�ϓ�?���H�Im?����O��ț�t)�p%��r������+��>�Zw�����_ќ)��5�B�!�E��'��>��`�7.^��6��O�>�[�oF/T�az2��O�3y�	+]-����2��������VX�X��m��W�l�q��P�6hD%� �Oc��֧���$�(`�M�'C�4�ౙ�(Y��6�'+�ɻ���ǎ5Hnu�w�l�������6�'�ɺ=Cq�H��[�j!(B��91�����"?�/��fM��j$�H�I_"Ę�Vjy�S�H�<E��(��*�Sw�V�Da�9)�̝<�~b�x��'�?Ңe�MK�Y��l�o��ҕB*ʓ��x⤔�Ǝ�X�bfI��)�H���M޴�Mc�'��~r�2nA� "2�����V�4i��(�PC�	b�j����=mBv�yr�/c}p�qX�dJO>��c?y�IS�(��(}�����L����>�b���� �M�9xMpwHt�<i�Ȅ/��3!n*; ]�k�q̓���%�'_O<�q��W'f�&��bK��O~���'n`Ň�0���!cmC����*WKF�Oԣ=�}"�$��9�F�`0Ŕ�bg�T�+gx��
��?���xYj��� �qW��K�� h葞�@��d�>�;g�@C�MڡY)Μc�ŉ�v���d�3�ȟ��a��R`�A�m˹)����"O4���QP�0��p�/<j0�&��hD{���D�O8�h��N 2ڐ��T��H���`��� �Y���U3_�q���ُ$�B�c@�>��3�OJ\����2#�] ����<P�1"O�=J�	]>!Z�E�W�X14U����I7	&�3\Q|�����P� {���y2��+�H�iu�� �Ԫ%f.���2�O8���O�/@��H�3(V�x�����D?�	T�'s�9���	3�����$SE�ȓ7vʀ+L�+��Uk�I�A&�\�'o¢=��EX-q�@��rKx�C�d\[.,�ȓ>$$��̗� ��kQ���c�'�abJW��2ъ��\(O�qCw����>񅮲<A����H���4�b���)��<Y�'ZL�H�O��	%�����ŦO�ѱ\���Ƈ	�j�F%(v�'4��m��	r��Q���`~ƀ���-�06-:�$Dz��$�$K	��x��[�4���!�D�<A�'J�Oy�ɒSW���d��*
�\d7�˓""C��#'�PM��dݥ֊đa�^*{N�|�<�V�:�S�'+� (�M"p7���6f�0[,��ȓ)r4����*� ��#��6
��<��{s C��K�Pʍ
SH�@�BDz2�~�V<k6fe�� �l�n�	�)�z�<��HO�<q�Ct��3��u�<����sL�S�$;+`��v%�{�<����2
�j��:��r�l�<Y
�#HU$���)�t�L��n�o�<)V��-l�<�1�X�%�2<	0�b�<A���7f�+$N��@B�e��a�<�N)Kn*#�� d�l����T�<a3�D�c�Pkba��r��Qv�<q�&ˬj����A͔~.�$�2&]n�<���^+4�=�3�� ���RMT�<)RI��$�jl
FfD�t�0�heGWS�<�v�Yu�RYń��.�:�X�n�e�<�􅜁,l��x8�$���K�<�a�SW��Q3�F�T���hЃm�<���EQV�z/߹+Y�e��k�<��M�8��D�!e ��Dx��h�<�+!w6�xS��VY��#��Z�<Yp!��P��$�/r��AN�<�v�\�b��]Ct��_�����K�<�Sl�7�2q��!X'U��kШ�[�<0HŘKN��*
���`�gIs�<YÇʡY�\�j���&c�̈q���Y�<I��R�.�T�rO�<�nݒ�V�<���@�"X���	ܗn��:���M�<	��Ej44Dd�0�q� I�<��*���d`�#\\��J�
_A�<�b���[��UK�H_0oX�(�B�f�<ٷ�Q��J��D-�� �a� Ub�<��@P-1��I1f%W�E�FPQ�(Pv�<���ڼLOh-Y��ߟO"� �_y�<�	�Vv,���66�@p�
q�<���:M�R��b���o�<�u��|$^ ��"�'GB���@�<A���EŊU��3F���D�d�<���nf�X�&�ƎDu�AK��_�<�.�X��)bpM�KV)�B�ɹ~
t`$��:�E{�a�2z�B�	.|E�Y�E�
(:H:��+ξC䉾n��B"�Z)KT���3뉅@^B�ɧ���`�Z�:ղ]d�=qd.B�I���2� қbzժ�Fɪ��C�ɋ-�$ Ї/��<�X�$[�-�C䉨�D*⅜�b���!�܁z�B�)� ��cn^�<���y�'Y�v�z�A"Onm�$��f�(tf�3H A�"O֭Ru���xܒ���[����"O��ÀF4,�!ٗ��M��4��"O���f�:���ӓCX?;�0�j�'l2Y��������	�,�I����ɉ$�H��"$�jd�؃������Iğ$��ʟ$�	� �	ڟ,�����I�`�,`g�M�@����7����� ��ɟ���ٟ�����X��ݟ���ğ���"g���h!Cކ(�,�(ń��=FH�	̟��͟���ڟ ��ܟ�IٟH�I	<�t`�' �1"|��� �x��I���������	ٟt�I쟜���\����!$7
f�ڢ"������ޟ�����4���4�I��ܟd�I�[<LA�b�Q��MZ�@�].���	�L�I���؟x����@��՟���#U��L���*�<�O�>><���ҟ��IƟ��	��ß���֟4�Ir0؁��E�n`�����X�I��(�I˟�����d���h�IԟX�I3$���E�͎e���bBQX��'���'���'Q��'���'l2�'��p0wL�Y��a��A�"2�Rc�'��'�r�'5��'���'��'[DH�vGW
�|��ؠGoT�0��'��' ��'5�'9B�'�"�'D�d�Ҫ.���	7�Z�M�5�1�'.R�'�'���'��z�H�D�Oؑ*���: 0`�{f�#�|��HFiy��'A�)�3?���i)H� ����t�e�Ҧ��Ȑ����$ ����?��<���yи�ҡ�*�%�,�$h���?�,��,�~��'M�)�?���x��Ǌ1�XA�#/(� 1)%��O"˓�h�l���gH(Xw|#I�o����E��ۦ�	�h.��M��3B��wt�0�0ޓ+�|;!Ʋ6x��!E�'��:Od�Ş+}d��4nN�<�(M�u!��ٱ�_]���;Ɗ��<9�'���$=�hO���Ot,D�9Js��3 |�0��ܖBF��<�J>��i����y2`�E��Ȑ@'7:*��@�n�O4 �'��'/�D�>��,;�i�V샗3�P�G�HP~B�'G������OG�����ݭ	ĺ�����*�F�p�Ƙ��by�����󤇾
u�S�H)4<T�kS�ƭ����Ԧ�)%'?Q�i��O�ͽ:��E��E�#B@}�וm����O����O����м:��I�|���OthE'Έ4KI\�KPbZ�Ɏ�a�#
t���4]��%?�����D"���`��t�<�	�b<?��i�҉ӈy�O��O����˗h����hƶo����� �>A���?Y�'��O���'Hq$���
Ҷ���C�Fr����ױe��|C�O�5��$M����������?��y�P�Q��01�3��59��M��wy�\�H%�|�ٴsrD�ϓ #b0��	޴��Tr���,"���t�f�4����O����O>D aiT%�ѡSI�'�0{��̊F��dQ�;O�y� �O>H����T�OT����ab���3N��_�rh���p|F���B{����Fy^�"~&��%a:�B��,]��`25�u̓tƛfi�/����覡'�,��Ǜ�q�TMU�:������<�O��Op�ĕ���`�v?O~�AE��O�����:��/�X$���=����:�O���|j)O���Ҁq��T��!�H��]Ѱ��>��d/�đ¦��M2�Iw�T���D�x�c�%��7"ZAH�K�
��d�@}��'�=O���d�hX���G�i���I���a�J���LF
�6�����"mXp�I#m�E�6ي�pq�ᛏH^�1�'*�]�b>�o���oT�j�H8��-��b��cC��
�F��O��mZ̟0'��s�0�	1#�<�&��@"~A�B�M�&����؟����m�	ɟX�'A#�T�-?�Q��/���X�Et��!I��FW̓�?A.O
�}���/8�Pt�_.\�X/��h3�i@~IȊy2��٦�]!

��p�߷s���X`�! �����(ϓ��4�$���O����S�
��$�y�8d�FG|a�u	��'��˟����i>��&�eJu�N�&�D����H���	fy�|ZʛV�����'lĥ���3+��-ه�ؾ-Њ������O}��'��8Oz�O��YՋ��t�r��T�;v�%��?��O>rq�1'E~��'�~��	2
��c�ט���6j��ئaO�s�'`��'R��ϟh��IS�D�~|2�.
�pq�$���8޴[d�p�' 7m&�i��!�E��(���1���x��8�|���4:6�vc�^��KK0,���ORaP�ˏ��� -�57m�F��#1&)8�*I1dߌ��?�,O��D�O`�D�O���O�a�b(N�]֨@��G�;�����<1�i���O��dj>��O��	��;DP9�H��E� Qƨ�0����fӒ���u��?}�Ӗa�^�K���<�N	���0��Ru��0v d�'�8���O?���$�2wODs����(� ��Ǖ����<�(O��O��mڃ+&�	� �r�7���(��(��҉e���ɻ�M����y��'g��'rH�Eo��'H�tQC�&SϨa�l�z����'��'rN�Ӡ���q���q�? �k�O�	wH��G�4ż��q;O����<�*O?1J�'�R���e�$\�jaz&�"�	0�MK�D~�xӂ��<	��Щ3xp�)և��M��._�����d�O��D�O�,��@��$�OZ�ג+�aSČ��T������"2�p)a��E���=ͧ��$�O��ҧ�W�&�.�6M����2G��6��ᦍ9&/�I�?I�Ӡ-ƨ���r>*Q҄�� -���'���П���<�L|��Q��}��.ܺXz��C�O(�����O�4�2�G�i?1p�m�ti�O��JL<���͏<��r�^��]j�hλC)�͟H�����D�Ȧ�XEI��*geW�n$��U���W����'ɧ��'_")�
�*�� �>��q���i���'6\a3��y"�'��iQ�?q�O<��FME|�����йY�&[ ���O$˓�h��iRWK=i�,����	t�� ����i��N>�I�?�'?M[�����#) LXch�������@*�?���yRX��Sޟ��Ɉ5f��C�~��K��
Xz�8! �0�L9�Gh�͓��C�����'�D=��o��H��x��_�H5$���'��	n�I��M����B̓ron9P� �-&�t�#� ��Y!����
���ڟ0�	�<ɭOkA�ߡW���j솰^Qp��V3O�J���O,�FXmh�i�mZ0�~�d��?AƬ��/.Q��`Q�1憩�ҋۏ���<��S��y���4=��Ĺ�o; �)�D�Ю�y"/fӐ��F��8 ߴ������C�B^aU$�z���fɋ�y��'5��'9! C�yR�'��	��?�(D�Vjivu��ש*�z��	Ǿ�ў�ZyҞ��#�'!����Rŋ�x~B��k��� Ħ9	%�(�	U���<p��λB���W�3j��� Y���I�����'�?��J_�E;�g�8n(<T������Īu̅`{���'���˟����	� VZ�w�qڠ`��	���	ay�]��$�,j�4
�%̓�`���S���)A��+8�ϓk����'	ɧ��'I��'�!Fq���Z��J���v�~�!��y��'q�A��?��O�������g�	�E"�#$](� ��O�b���I���	ߟ�����������O}�v�(KfR�j���h��Z9o��?�ĻiM��Ҟ'F,w�8�O���g�0Pu-@���'��a�ݟ�'\6M_զ]�7��r�"t���	�:��`�d'K9;���� �T�`CJo�D0��<1���?����?i$�R�谈��2C@����96��:g�4��Ǧ1"m��?A���h�S�߱���%;��8b�E,��-�%+~�x�I>��d��1SݴCu��O-�i���Ո7�X�0O�����9�����R�L�>��rgȞk%�ʓ�:#���<��yR��m�ɢ]��L��J��y2�ۅ�0�yE�P��,��".��O���dfU4A�2���V�+��iF�G<D쁣��ɢG���B�1�� �G5`zƜ�HX-^)�`�P�N	(l\�be�´k�|%V+7q2$�@�}i�As�IOy� �� �;VE9m�����Ӕ=� �`��i"\%�E�"iԙh��A�7��j��ܑ,Ȗ��'�J7��M�!���x��)�$�O��$��O����^L�gAV<JJ�ic�*o�_����O����O����Oj��OΩȵ�\���6��g:eRQ��5δ�`W  1��D�OJ�$&�d�OH�$HQ����3�*�r#ٙ{��XVc�9zט�o����	����Iӟ�	��ҙ����D_'��Y¨�f-HݛWf	�M����䓒?���hJ:qQ��?!��n61��j	�~����䁌�p��b6�i�r�'�"�'d��5�	�O`�)�+*N�9d㏦r���w�{'d$�h�I����������$��� 3%���㴰�p͞(r���3D'��h��!��5�e󤍅'y	��J�'�r�#7
{P\e8&���P`�'! 4���_a�1I2�l>����]U�� g�.gV0�gA�u>@���'FN�	��DN�;&��A5��{���U����[�-��"��ע���16Μ�{�U:���.(] ��A��y״9Y&�^�9��U�C�,�8@���0OQnx��π<0ӂX��LS���򤌆�DF� r��'�"�'�"�`�E�����V(�xf�5�C�%�V�@�忟�R��&R}�1ED*<O���ҪDt
E��H�\؃g�O��aS���JevH���'OB=)�B�5���󆟇ZFB$���'P,� �'��7͒ɦ��<9���J+c���a�jW E�h1:�T5X*!�� =�j�R�,�z�@�0¥�R�-Dz���T?A-O�E��"C���f��b
µqfk�9ydS*�?����?1��ԝ���?��O�l��Zw�@Y���ʴj���ht �4���䙪#�B����	����%e�%~G�<����(t�	S�H *Y����K/�p=1��ϟ��ڴzP���%ό�YN܍c��|\�Y�i�b[����`�S�d�ƜZ�ܸ#�G�X�d`b�ɴ�y�1gC���@2N�P!b�.�y�
�P?A,O�SLT|�T�'?哊E4d���c�64�	+&��Ʌ��zGx�������ɜ`7�dȴ��k���IT=R�P����aP0Df��dG�b�t�5�#mA2T�b��)T[�H�g�N�(��zf�Һ����r���1MJ3#�Б�L�'�|����:ܛf/:�3� ���gU�a|H��5:�52Oz�'�O��1�3H�����q��s��'�6O��r	�$B��8���8=izC4O\�W�LĦ�������O$�P8�'�b�'p�T#�nL4hΌ|���$q�����-[��
�/<�|�� `��s��d��]#�p �A�a���7�Hs�:�#��,2�x��ژJ]L�~�ɰ�<T˅�8{�1ڢ� v��A�󟸡�4L^�)�)��ʓ(��c�%/R�hDk��03���ȓ7��B�*׎����\G�!GxG*�G����'/�(ْ�ע,]��K\�eL�A�%�'�Ҩ�aHXm*��'W��'�Bj|�5��џl���62����D͘];���^��ڂ�bLH0�ᘖ:�:�k%����)~�����A�6Wt�,`s���\�G�W�Lh�t{�c��H���ן|6m-`TF�a�,�`}�@�u�Y�r�?,F�P&��~����?����hO�˓NA��$�T(u��cˣAo��ȓ	^���� A�j���:/H��f�i>���sy�.�w=6�L�R�A��w�l���ʐ ~�\���']��' "�T�mc�'��I ;��@� �+F���U�!�Ç��L2�ʖ�iҶ|��	�_���(B�,�Ց��:�r��wD��6�P����}Ӯ�ϓo"��	/�M�C��h�HD#Q"M"�(<�gƔ�'K��'�O�S}(�,a�oA�LR2PůĉA#�C�ɐ殴i��قC�l���kA�XA��+�MS����$��nM�O#�Y>!�������lY�k���5@�����ݟ��ɺQ�t�b'-��5��M�QJ�X�v	�t۟���F�V<8��d�~Ā�9�	b"p�EꐾFt���*\~�Rm �OT"=�#a؂��  ��e���@��d$U�'��rY2���N����"V$r���9O��D1�Ov|)"Y�&��դT�S�)3�'Z�O|����$_4Z�A%�:u�x��q3O�+�d�ܦ%�'��S<�x��ٟx��?r:1ˇ���MX�U��A4`Ȋ���ݨJzaꇧR�nv���F����>���2�s"�ï5f�� "� =l���`%î��L;`ā2�����`�7$�4F���b��8xT�M��aJP���(���?�%�i)�S���?Y�'Y�9	�o6{\�9��F�Y~��'�^�ۀ��$�� eeޤg���a����`�'�6��Ox4a���E�s�	�1���U�O���Ŀ � ��O����On�dJѺ��?���Y �>�SM ej*�x�r�̓�3��=�#�6A��O����+QX̓+�8A[UJ��}$µ(0�ͪ.u>����4g��p�C��8�P�["�ST2Wiɢ%���1�$�Ly"b�!2Ҭeq0�o�|ܫ���!B��r�g�Il�?��?y-O�)���_����F�v.L1"O���e��&m��A�!`�U�uSG�p�'FzD2��'U�	4���Yw�v��#��M�VE�7��?�`�ڥ�'b�'�rΙ�Z�B�'��'<�D٪���0W��d
���8K��x���#Si؞�� hX+V���+d�p$��H��"�n���b��������8�?At��;,�n�I ��/w���x4ϗ��M�2�1��<�ԧ�;r'(Mӳ��f�j�
��E�<q叕�' �-��ċ�)f�\zp+M�<�e�i��S���W�+��I�O�ʧv�q�HS��E9'nߡwr鋥���?���?��D"o2(a�NW�%��HW�i��nS�	@�e�V���цL�;gc)�(OP�󣚊K�ZeS�א/~�6Mh���q-�--��5�Q�Dx\�`�@�l�uFy��X��?�����O��(V.L�f�X�oO� EA�'���'������95�|1I��P<��̋�O��=ͧRz�'3����ϟb�JUXԄ�\&�Ҝ'ul�6�wӐ�$�Oʧ<�
���?���9�Tأ�]���!6ʂ��t�jI�(�JH�׎T�P��<�L��1��\���ݘϿ�&����%#�"(&&I� ֛16a��!�R���Yn@Bà/�]����
��$?��<Z����I�	Hv�H�	E?\��ȫ�(�O��$�OR�)��L9`(?t� I��HPnU3�k���IYx�8@P��2[�e�V�g�@y:#k70���8�Obf���m�4�(�i��<O�lҵ�'��\lQ����'���'lR�c�I�I����X��Ӳ���<�Q�Fސ4E���D�P>+�>�Aq+�U<�>E������!P4� �~y��%u�H����d@����r���j	H��&��\9A&�
D�߼ �u$� �M�K#,ʲ%ٜ�?�pgB�?A&�i�6ݟ������'r�K�L��F|駢мH��q�'��x%o�Dڤ�R�׽?��2��0�hyz������D�kg��;/j�H�"�%Zؤ���|(����?I���?a��S�?Y���?ƭ	�Mt8���bN����t*� ���2��=/�=�s+�|Ξ�
��2:��Dy�G��A���p)�F��0������@�bM ":.�J�ÿ^ �6-�4c�F�A�ɩ<���$�O���#l]���4�el�>sK=f�JOd���O���g�? l(��i�P7޽�0�]f:��H�A$���hO�, �L��O�n�R��º
^�;3OZ�n���M#)O}�`l���	˟@�Orɉb����.=���y�0�Ya�X�/z��'}Lك$㛆��%{ �S���
�M�F��Wnb�P�aN�c�� ��ޕx �m:	%ʓZ�� Q��c�D-r��=������_"�X�/�0?�h�UW� ��`�=JQ�ȳ���Oj��>�	�O�5�7럊'&�p���߫H��p��O��"~�l�Z�;E�V�
��!�^�q���'ў擳�ē}�8�-��A��:��4W�>��<1����<1D�N�����O��^��+�K�n�<�b˜"j�Ni��d�;U�(�qK�f�<i��]���뀀n��IJ@
Pw�<�N��^�~@������H�p�<��c�Z�ޑ�C��g�^ؑ��m�<i6��R��YGE�;�$��h�<)�ˏ�!^�M� K�?t7N�Ҷbp�<q��Ƣ5�Y���6X"4��oBl�<�%e��n�K�ٲP����d[d�<7��g?��c . V�nг���`�<��>u���pg�
N��4G,�w�<)���0<H�b`N�#?\���Ý[�<Qp��Hx���-���qu�W�<9s�ƣ%�<�#�!������U�<����0eĩ	"ʞ\����T�S�<a�Kd綅��L�;1֝#T��O�<1w(�:E��<#�F�-* e�gm�L�<Q5�P�
��h!A�8%'|�r�m�J�<Id'U����!�����,�1�G�<�F�	R�CBI�$@�(p���Om�<13��>.�����p�����Q�<	!�S�R�J�3��a$#^u�<����/
�b���T0.v�1����Y�<�V�ۢ^$d�a"�ɮ`��H"N�[�<�[�y��ɖ�
���,s��B��aNҹJ���RF��AQ�h��B�I�<��	vHM�,��C�N�K �B��(&���H��ףj'��qF��	t�B�	�(�&�;Ռ�:v���Ȁ'm�B�"��ț�)T�#���)�`ߑj��B�ɽDM�HZ�H�V�­�nQ"^�B�ɗ	���ڱ��%<�pi �(Ze�C�):�D(�q�.T@�k���]��C䉽'����e�T�$E�+�
B�	�Q:<���"7��x�B���C�	�Y2��WÛ+m�Ĳ�֠xB䉧C%�4镃�O��p��s�BB�	)A���x����@���C�	�Z�zdi����9�(P�Nl2�C�IT4�#�HU�t��DePFB���ʐ�7�^RTI��֎U@B䉿LJ�-k�e9b`Ne��,D6��d"�Nd��T�6�ɠH��2!�6�C�$(!�A�0Y�b�(#�I�p��u
H�O�z���/I(��B |(&bү 24��'xPM2��O!$� ၫIrP
H>��cK�tؤ(�mdDe2c/,D�v`8J>1g'v�ݲc�6(�n9�'��Aؖك�*�2�l!��Q�P����e�H,����8��(�6e�Wv�0C�ԋ��q�(��rat�L�����1�ׇ��|CF&��Q���"O=B��� �F���-H�4c��ZgN!O��q�`�ҍ��b�EP`��)�+e],��n��h��� OW������'@�=��-��l.�mz�$S,�wKQ+6���{ќx2熂�&��󪉓b��`ң��'��2!��d�t�"U���E�>�iP%�S���D�EqO�%I�����b�6�9�:Z�f���AX qKZ,#�`S�Qp��!c6�!��D��"�Z�s� ȎGR��0�CR-t�)��EW���zp)�<N�8��Ƣ��!]�dٲP8A��/0��3��I�O��J#C��8*��S��< �P�'��:vb\=N��m��R1E;�� *�Rti������4��OΣ=�'>¼��$Ϲ&T����$�� r�i�	����V�Z�Au�Of8s�ĕf�)�L�=N<:e��ۼJ���F����d��ކo�o�����;��X�2'��`q���Xw%�O�ؓr��O����25�rh�d@�i�80��b���-E�Q���k@�)�\PU��b�:-k�L�8*1�����%�J�+b��R8��ؔg9(	�'hͯGk%�ub^�4P�>y�'�~<X� �Ss���O4�A�NyԈ(9@�T�:�x@�'��P!���}
��a�d���)���;պ�Q7.͵V�x2ᯟ���tW����w��Oj�6�5��m�ߴD�Vٚo�D�iD�g
�@ۃ�x���{N}���
s�ۇ��#�'y��D`ܛ�
�٧�Z��B@1�<Kƽkݴ�?���](hƀ1�c��ئ](Tg����B��PJBIS.x��uKX	+Pa�d4�P��?7qOb��Ⱦ�D�J:
�hV��:b��*�ެ"3p􁦫��&|��'��B���(6��5 �;u���3��F`(�h��ׇ��Bh8�(�' ��>��S?��v� �Ѻ�eL.>f�	Ч�
H8��"C�Ҷq9��C#H�:j���w	^>.�<}���jO�1��i��~��O���_�g�]�+�pi���>�rNn6�)E+�[/ Q�q�Ď2�\�I<����]�*�7ʖ<v%h��g�@�^Uf��C!��_t`BuH[OU2���?���i�T�P-S<�f��G)���u�%��J}���QkΙ1-��؁�S�mp����\5�׊�j�'i���  �`�S��_"i�V�H����{� ��E,�$�v`�$,��i���AL�6x
Ճ�CPm�|�%j>��~R�\����~:ӏX�8Zd�᪗CEJ�(��K��p<i�ᗋ�+E���o���!R �@��|Y�I>Q���7�	`�tO'V:l�G	X�<	z�˒$H	���B\�T�".�F�	���TMLMOb}[�+�$iVc��xс��,�����m��!����ᱟd�	�� �нM\���@Z6����2G&��D�6���ƎWł��!��Iqv�T�vw�� G傣�t�'����j��x�C�ͭyRhP-��Vii����y��ݘ�)U�FUY��i��� ��,VX�@��A�m0�"6b<���'DF�S�}��mS �ċv����f���-�d��	�R�� �'��.��y�a5m��h�b
�SqL�(�D�=��q��'��㞴�+�L�*�T�}W�p��4_LݡRLN�=��t1W%O�$L��G�xb�Z�Nɘ ����{Ԋ�볏����'�rHc�)hp B���NU��r%�q�\�d�qO IC��ĭ��JSH˧H��� @k��!o\z8�0-��<
�	�U0lO��A��&x�|��S�Y����be�\tnl�3��?z�H��)OkLG>�p��^�w�:Q[�@=F,!�D�7�n�a!E�k�< P���r����4!p���@P)2�ʼQ��U��D�SJ�&{P�!�_$Jh���>D�`���ѡR�"���ͪ�t��P�lJ�i� 7X؉'�ؕ���>.0��[�	�."�h�}b�TVH��Ta�0{q4��C�[���'���F&$��@v���J�؉O>�T��)Q�6��bn�,6:`s�H�	��`�?jf���f�3\O�	AgOR&[�^ kX�01��A�04v$d���ŐA0�����'��=�L�m���I!BR�\����O�m�&_*Q��8H�"}
я��X̸{�� |x�Ix��y��@�x�K�P}�����>/���\hX���[���k�F,�p�e��4p%���#b55���9Ѩ�ؠM���7�Au��@�v��D�.M?t��O�<���D���!R6A������`PHp�e�ў@�t!Xrg�rx�'�����in�C&�E=F2��ٿ~n��b��$RZ����:?g� �
ȫ?>d��a�$nڬ�w�+P(����K��&���6s1�ċc@3�@%"r8;�"On �s�����@���}�����6O���ͯV��t2�������A@l��H��+tYP��Sp����M6T#<�D@&A���@u��,2�t��"3g��"��xT&N(��A
ÿV(��An���'d��ȣ;���4�J3B��:�{r�	�O�Z� G��$���tM����Ȝ����)��f#�8,ۀi��܉[��Ff��,�a{��)�q��
()tpH�c�H19�
�|, ��F�4_��xZcm���@��r�H���G��2����D�	��ɯ>���~�S �Y�D�4e��m 
�(,��	'9�ѐA� (�����f0i���;���Cs�	n,���'l��O,��J?����3J�����,f͘�@�ǋq���?�5Y��x2 �/^�.,h�*�T��y��*^��'YDa�N�^���{�&��j�ɐE&�~���5�A�P�]��?Q#���RO>I����x�x���F�L~Z$x��׺T���À�8�n����'I@qp�

$#�h�`�M,�D᱒@W��B6��I6�%�F��5��H�`�l���D!bQ&���y�I�^xΜ�!����"��xr�[61�V�7�}A֤G�k1��Ɂ&�0<��*�;%f�����yDD��F�9o����
� �\�T?cz�6�Z2B�=��x�e�$,My��I�KbdQ���'�8q���:�Ve0�E�-4���d�6Z���l�Ѐb�"��m��'1^T����}���)I�Y��U5YL������Ԓ��d��.�b�p��?~@N|�b�ɢ��� �)�p����k֚���t��ׅ,ш�����4�hQY��|���T�'��QX�B���Q�?ve�A�:a��9Qu�[m8����&h�|�L�5/5F�yS�O5�H*����
�@��R����O
��$�9ce��Q)�w���X�*�nx�Jb�%brf��Ԫ�9��x���29��Twb�-/�B�G�ρ��'FV]���J&T�8��L�e3�'~,ta@!֙S��U��FAs�V\���Z'f��:��|B��P�6t�V���5j��w��/Vt,	AcS�*%��[g�6lOX�0^�py5�Ib��`4�����,���7Se#��9Ok�Ϭ%<��	�<(�셺���1~�Q��X֘>	qŏ�C������	<� ��I�JW���F�T������*\�cD�;y0R�x�՛e��U�B��@r�DD#p2�9�'d(y�O2�;T*V�	$HQ� w�D5 3�'e�T�6�YG�꽰����rB�Ό��e�pR�D�Y�1)��D�Wv��>�����녉ۮE�&�J��
8H������~X8�Y�eT�����N��������e.M��P|(Bc'
D�Y��4aI ��O�T�a{��Q)l,�$ѵ�DY��W�=h���j\2��u��C���xZc-62�DD����Yezn��	.U�#��6C\M(ѭ�+�N�u䎼�����-O�M8e�Ʊ{r
��&w�Ju	f�V�v��T@j,==���sE�`�[:.�Ț�,��]��
�*�zY��A,���M��o�v$jæJ%�v\Y��ן�ēL��캶׏k����Ϯ��U�>)g��+��qIDH�xy. ���؆R�X���k�dĴ!��� 	
�l+c��k{�pK@@���.��K�]7&^�"Gڜ7�Uᶡ_�t��dsg��0j�a{b�Kq[���T�-|%.b*P�+f���	ы)u���Q�Z�Af�xZcX��h�2M�4#u���w��X��S�KC���a@ (�\ڐ��3���b� ;�0͆㉊L�ٗKX�9���0��v��YwA܊.��Q�Z�@���0!ќ�XuEԚ4.��U�&@���5���@`E9�A�E�I�i��]%�@�A�Y�)�\[WC�/�VE��*��O��e�pk�2܍"��9�� N&+�&-�"��Oz��KJ.�u��ҍ)K4	r3��~�	�+��Re�,{��QCu��*�.�VAJ aզɰC���S��{�O5<����3ϙ�
 ��JVCV�|�U��AM�~3x��K��0=��M�,�������b��g��B�<�p���%Jv�5�ɩ1�TW�<�eg���]���A�MA��&[V�<���:߆���Ð/�HiDU�<�#�
�t��A_�s~�	!��z�<!bA_~�Ʌm� >�0��UO�<!%�X;n�� �GBסx2Pp�`	\N�<�� ��mF�l�E�@cz���r�<Ivl�pTڬ�ACBq����g�<y��QLP�X`lS
�f���nFm�<E��% �J�z�ŒK-\J�n�D�<�ڼ1D� ��X�b���V�<A��A�F������jy���QR�<�%3U��	�S�.u�8����J�<YU�6R�re���L�Ok���H�]�<�D�ǍO*@��p��%<t��&Fq�<�aF���#u��o�:͚�g�k�<A���n��pN,L�%�Fi�<Y�� y��q���<@���Ci�<Q�O�@|��Q\�T��Y�!�f�<�e�R=h�g��`�X�_�<�ȓ5�2H�1���oP�A�bۡnqB��^fm���wf�bC@���$Ѕȓ+���1�#�$Q �h��ޭf����y}8�(�$p~ 9sU	?o��(�ȓV�����
&z[N��W�P�ȓ3�BJ�\�v(��Ƈ��F�~��ȓ~
�jg��=��!>R�Hԅ��b��&+�BX0���%�X�<���H�qn�T`��+��I��Yj�<)uk��@Ʉ!CC$Βh��Z�/K�<Q���s&ٛr�W6fpEHSCE�<� .C�V�p�b�0�
�g�^5P�"O��w��7J����Ʃ�$`����"Ol#eGY�AV$!�.7/u(�c�"Otdiv�M1(�(�i���gb���"O����B�%�ȱ�Ck��\=l��2"Oi8Gժ�L�ԪC�#V��"O��bf$H��>�
���GJ��"O:<� nʳ?Kt����,C�4x�`"OJhõ�aGr��5暃 ���"O��QX�x�"$Ȕ��a[G"Ozu.S=!�R1��ފF�Fy�"OD	c+W�=�j��F�K6��k�"O�db&GΦ�J����M</�p�3"O�򇅚�l/6�����yƆ�*"Of,�bN��[�.���iG=f���:"O�1)��۬'S��)��Xn��"O@�PWl�)��( t2f)�{b"O6(�c��h0��DE�J(Z���"Oxh�Iב_�����˺Z�-7"O^H[�'U��q k���z�"Ov�h!�Y�m2R�� c�&�ڸ��"Oܠ!�N��J��H�"` ��"O0ٳp�^�8�`TP����"O@}	E�A@�A���_�@=3"O�8�C��v���rt ܔC~�x�"O̹�f��>vmS�O�����"Ou*�պ82��	먝��"O�%�	#A�6K	���"�&D� !�E�K�b ����|����0�0D��p�ʬk�N,�B+ˌ[���+D�HQ�A<~ܲ�v��q8��h�5D�xA�93�L����X�x��9� 5D�<�w$_,d,��s��ּ`b̄�"(2D�p�H]$]�\e��<��,C�2D� xr�MRA��)ԩ��h�����c2D�p�Ҭ�$VzH�5��}��ʰO2D�� %Vl�t����Vym�)��c.D��)��?�ډ��F�%�]�4L*D��2d�֫6�:@�4j�"MQ\�;c�(D��3�@�8Ĝq�R��{6�u�%D�p�1���D�D��A�K)^��#�#/D������rhm	��
�Ҁ04�/D�8��&��'�u���Ŏ:��Ę()D�$ӑ�� Bļ�6�+o��p-D�\���̓M������׃eӾ5�u+D�h��/K6Twh�)����$i<D�|�M1
�p� gAS�Z*��r��=D�xJƪB��%ѳ~�dUj L!D�`ZŌA���� ���L�׮?D�p����`��{f )C�%�#'��C�� [J$�
3�=<\�|��C�3A��C�75���	`gX���d#����$B�Ib��I�n�*p��#+�U(�C�	%s�0��#)�"b��E��l�;\� C�<|�R���4�va#^ C�	��\��sM!}i9�5���O<C䉛+{�٫�jM�(8�3���W�C��8�^���`��,��"ayi.B�I�'9�1hq�V�o�a��.<.�C�	�'Եi4)I��ѐ4`G�z|�C�I�xވ(����N*p��b�G<�C��;2x~ h�	Ͳb�JX�TF׫soPB䉘;?��:�Ś�0QVlٵd���$�ĳ��J֥	12zI�O�$F�Z9��;D�� T�AL��������A�"O�P'�1m&�=�ō�"VfD�y�"O����$h�L��R�?z6� �"OXP�@K�0V��  AC�)?xD�P""O���5����l�Pk�Mv�D"O�VS:V"$���o�.C�$�q��[�<y3	Q�-�������0X�`%��ȅb�<"�ǿ���XŠ�8���S,�T�<��YH�!� C��M�Y��R�<��)Y l)u�X�23��	�Ux�<�S��(V�u�b� ?N��R�Av�<���26*�2q/x�V�0�Ep�<��7}�m!���=N])SP�Q��`�?a�̑�rI�À�=����NIc�<�2�:C[:P8Fo�8*%$ibPeQ[�<�gV�;��� �D8dH�� ��l�<��'ѹ
������Z�BI#t�B�<c�L�hW����yB�R�!Y�<Y��Ý{JR�#�o�A^�L�w�DX�<���Te��#��֟%�����O�<�ѯN;/��1&��+P�@�$M_M�<�B�F�3�rp5�����@�<1Ŏ�[@���nÆw��[�|�<1fA-ht��X86rs@)�N�<Qֆ����a/�l ����<�#c��$�Xe�����-2��FJT{�<١"�8�d�;�D�y��j[y�<��Ȅ�K[ ��R�M�RdB5N�t�'��x����unW�'.X�*Te�%!��H��(2b`;���vL6/W"  ���=Aۓ���Q&Zs�����C�{����ȓL9`��aU�Zz�Y�Asr���V�ՙ��̐gk>��D ��^�~��ȓ8�pA��o�QV���h��{&�ą�S ��D�+��dxE�(YYJm�ȓ	���EmϱY�f(wj�&#���R��)2�_,-xZ�K�			v�ȓ8���1��/
*��@ʉ�iz���'1�<�5j�Y�R��c�-n0l���'8��h�
��jq�#�h.�p`�'�$�'�\��1�c�Ŕ(�E�'�6\ز@Z[����͹'�t0b	�'w�|�b�.:�x.i���PㄘE�<���S����/�H�*}�r�Z~�<�4fC�;Ѵm��HZ;T��Dpv��q�<���Q&�3���g��� ��	j�<��	��XS�ݨeNF>6A�Y��c�<�_�5��(���Y�58� �`�<qP냫�8!�1�K�O��@8`c�<��ŧ!^��R��AV�@r#^�<ɗ��}^�@)��L�^��aR�f�^��0=	0��9^�5Q����.��8q�
O�<�7M�?F Ĺs�T�W��s��v�<Y��L'62N�����P�8�C᪄i�<Qt�I,u.L�ٶ�ҩ��$e�mx�L�'	@`�¦�t L ��3jB���'�������20oL��	�1-SjM#L>����iX�H���`EX0�ʜ[��0hj!�ۓX%����_��d�S��MF����'�S��%ʰ�"<��H(��!��A��s[!򄓚m�����)��5!	�!�DH�<q����t�P�q5�z!�0D��H3��
v4����!�dO���ZT��H��Л�i�2q���~��H�� pp1s
úv�Hi
�(T��� �"O��:bA�r�\�S啔B'�r�"OzjC���q�F�P��"O`����2(���!�k	9�X��Q"O���'����\��@�8�.�YC�'�O��@�ӄ��K0��. 7bA"O�|BT���P���Qr�E&$%%+D"O0��5I��Zj�SE�+U�΀��"O`DXn�
e�5��'Ǟ=��T�d"O��Q���z�� :��͹`}U3"O�`��[�/�e+��X"Ds�d��"O@Т�A�s� qj!id���"Ox��Dc*G1�m#�� )K"A�"OZ5�S��Z�^����ʝ..�i�$"O�,��G+s��
����.��"Oz��3E�,-����%��v��<��"O&����$QŲE`�!n��x[G"O����[r�Zh�G�B�A,pˀ�ISx�<���J4zP��j���U�`��!�8D��jB��j쬍KF�' :�R&4D�l#vi6�p"�d�"fv}��%/D����C /�^h�&f'7ؐ��-D�����K5A˦��?8N��P�.D�𩦭�_�0�b�A�%�NT��-D���ӊ��r:Tp�B i~l�O,D�x�"$�8��u$��j���%>D��j�Æ+����_�]"�3#&:D�TxpNS
-�N��a�ifD��+*D�4�I�
YW�A���>��ը�e'D��y�Y�
������
�p)I։#D�XC�ھk�2����L�6�A%f D��"$�L&<x�Q�s�J �H��g<D������V��Y��	!w*0ST-;D���h�mGx�
�k	�g&���<D� �FȖH�	�@O%��9��>D� �v�`��� 9�1@r�;D� �p��%V�(���� �t5�p�9D�L9KS�a��xi`!�<�@Q�5�6D�(�1H��[����l�f�Hy��4D� �D��D(��U	�W��E�-D�ܘPoR�=���4r �$C�)D�<�ҋ lj)�
)JV�PA#:D��A�n�bS��;�o�����p�N8D��xs-@|ԘS�"����c�7D��X�e��Ga�{Sf����I��C6D�� !FN6ex�P'B�ljx3�H?D��{��R7	�������!\����=D��Tf�;Fא��	A�!V�ia�(D�X�3�S2��2Q�o�`ԫ�a)D�\�pU:Ls��A�:(�X�+��#D��1	@�����/Ñr9:���?D����
'2�0��	P��	���2D��!k19�M��_:ϔxjr�%D����J�g�`M3t
Ȯ�Ę� 8D�t�F䝼*(i�U���"����"D�XB5�Г/~z 	F5 eN1�#D�(+�
M���#��W� �pi�!$D���H'g+�Qn�b���Ô�<D�4��L�n�0�3��܄Gȸ���6D��P��U�#0<B%�ڤ5������1D��gg؛Oc �sa�ա-�F�aâ:D�pBoR��le��[�B\
�$6D��+�_%r̪�J�`jpUj��)D�L�.ɫ:j0��>?�&Xkr'D�� �}2��A?�����kW$�@�"On�j������Q	� U��""O*=15
\�a
Y�d��E���"O�x`�D^3BW�\9u`٪c�hA��"O��K ��f]he�����{�v� "OfQ� $]b����.�yt�6"O<D*�*Ro��`x�+���s""On@ K�%[e<l������8�%"O��f�łw��P�ԁҒ=�<1!�"O\��p�ь^�)���DJ�"6"O�T��=\�M���F�!2LA!!"Oz����]Kz��`Uw ��!�"OHID�y]r,R�̉�T���Q"O��v�,X��ij��Sw����6"OZ�'��&TA�E�˔Fk�|�"O�Y!�;}�&�rV��#YXT��"OJYE+��M���S�� X�8��"O���2�W�Q}P��҄�9e;l��$"O�L����B�aPF ;����"O���7iX@X,A 6��;4�����"O������F�q�R�>x��u �"Oz����cUTa�Vl�3!��T��"O���R�J�lU*���� ���"O�u���G�YX%��*\6�6j!�Ă�?"d�I�����P�-9W!����T�f *1E�/d�N$c�*��!��H;N�gڎ&��0IQ�#Tm!�=Ty���ËV2XNu�w(�'l�!�DC�,�$(���F����1h��_W!��)dR)��#�`��p3FE�Um!򤐐WW0H7f"-Q�5�Ԅ7]!�Y�(qn1�mQ�>���(�!� �L �0���&��R�P�!�$�w�PTHU�]�yWd(Љ@�:�!�E&��M0� ��o-�Xe��}{!��@#!x,0�)Ր�p]s �B0�!��%#+�(��o�IąFB~!��LC<2��U�-2�B�y`d[�[d!�·oyPE#b��z�l�j�+r@!�D��>0ɸ�#Zp�Fx["'� Z�!�DK�o��|bF��y�:)��U6V�!�Ě�;1��F�,jQ�ǉ;r!򄅛p2zYa�aʉ1��a�f��=�!�O�E�@��쁎�
�"O��!򄄎eM֌J��=�4��
�7�!�G�GR�R���)j�ޑ�'BQ�!�$ܻwH����8X�P��U�	 !�ӳt��)�-̄�pD@�M3+!�$��l�bVFHfl�-	,)!���4���ᖏo(���fBԱ !��
�����y3�iZ��
T!�ɞSҼ�J�+n��L��!i�!�DD,���e`U�hZ�%���?!�O�W�=P']�r��`	V��!�_>T���'+]�ru��P��#�!�D��m|��b�e��^jpa1o�=A�!�DN~V��Pfn�7;9�<��n���!��;J�)�d䀍T�� ���r�!���.��<
b�Y.wEbP�lܖ�!�+w( e32bIX^4�peR�E�!��)M���D�٪ e���T�N�J!�79�.4q���9�l�P�Y!O!���W���	W.V�0i�c�W,P!���0cX�y�%�R8�n�@cB�8I!�� Hlҳ�P
/t-"�
�%���rc"O|q��1���4�Zs$l6"O�E����Cd�y���	�Dv��B"O<�S'�£�J0"c��a�ƴQ"OTZ���$�b���T%E�j�"O���C&OpL�(%N�4�
��"O�11�T�)���aLܡU[�d2�"O�Dږ$�Ɔɹ ��>kd�[�"O����&C=� ����uShܡp"OҸ�S���6D�-��-�
JQ@z�"O.U8"nӪpU��iuϘ�-���)�"Obi10�)WX�$Q5Δ+2�� ��"O84@.�&k��3�
����"O����(�67���Z:a�>
�"O�e�v.��U6D�����U]8s"OT���0H��R�6L����"O(�+w�S)
,�Cw�U=@�U�w"O��j�2���4(87�� 5"O�8r�iɇO�������b���"O�a〽}������M��
"OB�x��K�2J��I�HH�`<�R"O���h�#&�:UZfꑤj��XC0"O�	�"�U���X!��j�6+"O��s�[�<�TqҎ�$T�|%W"O.���G_
7`)(�ďL��
T"O�����A�$h�����`7
�k6"OR0CD&:�J�ؖ5M���"O��I�R�\N��I��˒@.u: "Oބ��5/�Ԋ4*�<��i�"OBDQe��k�H��CHՇU<�!�"O���D�
4��� jD<\�]9"O`}둈Z%��0A�	N(+��[�"Ob�Q�I�n.�X:�j�1"�>"�"O�V��2)�UqS�	,P�lF"OvQ���'ZM�Is�H�*P�p���"O4��5� �&���`b(��"&d�f"Ofx�D넏s�2 `Ȑ4;�6�q"Oҵt��X��g�Aܰ�6"O�����/l2��I!y��M3�"OhtJ�D�c?����"K6o�,�;�"O���.�&)�l�""��3��$�R"O���e@	?K���aȏ����"O���2
��N1��� T�.���80"O�q�Ucq����k�\|�"Oj�[vd9FE��nT�oh��"OF�j����(�^=2Y��� ��"O8Lb���:+�8���I�L��Ѳ�"O*D;� ��)0��5!�}�Q"O�f�R�HMj��wGS�97��K�"OF�p��@�T%ry�RƖ+��
g"O��8�#�*��(���2J=x"O�H9����]2�C��I��Ĺr"OP,t�"��Q`N@�|X�"O��i��96���ۇ�5i�p��"O�E���> �|���D��ȪS"Opyr�3vX��l]'P�� ��"O�u�@�!��3�Ʀf�8��B"O�y���%�zp��e�V<�Đ�"O����[
#�l![a��hH�"O��00G�K~|݂2d�4�Z᫴"O
a�����U ��&&X!"OEq*!|sv��Fh�PH�@0"O~L���10�d����)�"�'�*)�J��;8Y&�^5\g�%X��� �H�EC�㔥���ޏ_�Z�3"O��s��E]|$YD*Ken@8K"O���$��8���4�!6W@j"O
<��OúIಹ*�I�X  9 �"O� �E�E��P�1	BF��Z�"O�J�Ɂ7�HQRg�^(C"OB�ɖ��I5F�@!aT"c�x�
"O�Es�XD"���oF�)�d@""O8�����r�jE����k�.t�e"Oʸ�7E��D���y��T&�v���"O���v
�#b�k�J�N}�$"Oz�jO܍Ir=�R.Z!�,��"O��7	 ����̀:]��p"OX\Q6�-,~���1��#�3�"Of�*ԅ�&wHu4�

��x2w"O�|�!c�-bL@�%=��U�"OF�0�ś$+t��A�G�KN�8�U"O����!

�iз�W��5��"O�0)&�D:*S"��'Z���"O������#ps�M�sl�Bz�j�"O�젰���>�VQy!,�c�=��"O�l�`�0�2�S��1D���!"O�X��F�&��1W��S� �4"OM�դ$a	�I:a$��'Ϟqc"O.��w`:`���c � �d�4"O,5�`�Q����Xå��Z�x��"OX� ��?fUJ��
	P缘��'Ub���3�b�@dKKe���	�'�d��֫҇
������Lb��	�'V����B�m���p�ܮUj4��'��|a o�t1��!5IA���'՞$�"�ѳ(�8$� b�5C�h(B�'�����)�6	R%�`�:r�}�'9�uE��*<>�Ԙu��9þ) �'�B��叔)M�t��S��-/�<�j
�'��P�Ն� zd-���;+Ve�	�'��K$��,5%��P�O5)��8(
�'5pр��,af&�e.�(�B0k	�'�Q@d_�f:��y���$8|�1��'��`��B���A0%ʓ�.3����'�H��\^�:�.�-+�
�(�'Ȉ�K���r��"��*&�`dq�'�n�����'@��  Ӧ�4�.� 
�'WЭ���R<npn�Io�( _69c
�'�y��)V �LC��ޗ�M[�"O�tȓ�nE��#�a���f"O���@%Ū@�
�i�K��	��"O�!bV�^��(!��NU>d��"O�MB�oyK��[A�L3@�:�rc"O��I��zѤ�S��1���"Ovu�u��O0�B��;�Z)e"O�Aq��0P�dK�G@�f�\\��"O @����5�n4���܇2���"O"	���.cw��s���.���1E"O�R��L�[� ��5nH��A��"O���M2U��B��3�Ii�"O9�-�@2L9"gD'�vM:3"O\d2� �p�0�3��$6�^��`"O�(y���] d�CЖ:$���7"Ol-:�	R6���#���yJu��"O$�ffC0|��i�a��3X�ڥ"O�Y��Ɨ�l4��D랆\!�5v"O��I7
O�Ad` �. H	q"O���W$��6p��z��ֺ p��"O� p�XH�35p\����,
2�˳"O`x��hܲj���$<�6�c�"O�����ҒAZ�,Aml����"OLŨP#Y�N�q�K��9���"Oح��f
}ʨ2ф�I�r��"OdpbӪO.����5�u���bs"O��P&��4��(����+%nh�2�"O����P ���F�` j�"O�X�3,G,5�8"���#~W��0"O�����Q�	"���	��i��y�"O\�+S*�	>��9bH�l�l���"O���E��*4ۓ-F�;���27"O�jC��>q�<� a�F�6%q�"O�W�E���95��ve"O��NƎ)W�m�1��b�Ј "O��kcn�SŢ�H&d�.{Yvd	a"O���W#R,a)�P1����|s�"OP��EɭR�tH���̍r���"OL�Íz��3�<v��4R�"O��82ER}3��7�Ex���R"O6-���ê'��X;�^�5�:�ڵ"O�Ȋ7ȗ���Ÿ �@�b,�H��"O
�r��� R'�Dh�&%��z1"O��Q��l8J0K�'�{�f��"O$�	M1�R������!b"O��˶M
iR0�E^p�"OHY���њV� 8�n�o�����"O�u�b]O��Ad���m�ju�p"O����D\E�h�z� ��<x�$R�"O�����/�}P���,ՅVJ[!�N-*�b}s�M�u�P&J6E�!�$��HZJR�7��	��E�>�!�d�J󮡃`%���h8aC�~�!�=J��Ie	<"i ������!�D3cL�X`a+�:v�!Kw�֏w:!��S�_W�E[�c�Sk�I��=�!��{� s�Y�����Wo!��*.&U�҅�jM�h�MǕt!�$�U�v8E�ҬFe֍x5�րz9!�DD�2����E��GA� ��?H&!�dLc�TC� O]���ʔ�
	�'�L�M�_�l������`4�'.))�
t�<��,��L0�'7X)���dđ��T��0@
�'���)�'��1i�YB�N�Y@4��'}���B�ɇ2�:8��.65��2�'QJ	�e�73z�\�P�߹vo�\�
�'dZ�A��	K|!�K�jte�	�'l��0��c��K��c/��3	�'�:x
L����X�LgTPm��'t�ƣ�!̙a��O^�,��'� ����Y�#�BօD��,	�'R�	��)�d���'��6d�"�'PF���]V�]A���!?; �[�'=�iz�X�#g$�1G��=�ܑ��'����b���=�r�����/�vA�
�'R�T����e�e#ĉ$՚a)
�'?pdRb�u2H;�Ő$:|�
�'�UC6�(u��	%Q>���	�'�e+�&�7��5�cJ�sb!Q	�'�`AB
�z�Ċ�숁g5 �3	�'����iÙ)?bi�cHwR=*	�'�* �7�ؑ ֒�NN =��L��'����	
"KO�|�U/��H�Z	��� nI�H�9	����'�_�N��!q�"OnL1�ʂ�J-n�����!De�7"O�	���@<|�6Lp�g0�8X�"O�Q��)��p�
�F4n0y@�"O�\q�i��^�R��iMz��!"Od��$��\F��i�+H&9��"O(�է� ��Ј�+�M
����"O�F�`l��۲^�(A���U$!�Q"�IP@Ԁd��];�ݞX�!��#<\��	��W�� xҏ̪W�!��+X�����6�|Te�T�,1!�D�53����Mɯ}�L��f��x/!�$�B�D���`�5)�4Z&�8u!�$H*i�hQ"��3y:�!C�B�!�_�+Av g"�"8�뫙R��ć�D���bbKɸl�(��� 8갱�ȓ?��e�@ �������:9��u�ȓ,!P&O��;d�i���b�4�ȓS�L���Z)��	gĔ�}w�u��R�j�*�GE$��)�"�C�g����7�X�����=1J|H�ν#�8U�ȓ?��}RA�DOf�؁�LK0��ȓDϚiJ�D��OW�Y2Ī"<D��'�Y�I����1i\09dO-D�,�aρ<�����2��J�C�	"E���p�N�y�����*9SdC�	%�� �dZ�� �dB�O�RC䉨]�l�J�'P�eC4�@4j?B�xB�	�y�,0
��AM��Y,&4C�I!`Ԃ�PAP���E�$"��B�ɡ=�0���ff�)��L���B�ɉ@�,���V�`M��ʉL�ZB�ɪM�� �d
��49	&�̚**�C�I\}>�����u�MiY�C�<����8n�L-!j�ObC�I5�x���g�&'�E�7�F�m$&C�I/���')7,�`[��B�_FC��3kx�أ�Mn��bґt)ڨ /D���wCGe��|�Q]�@)q�.D�(�� ��ztSnN.I�ҩ ��+D� ��NȎTј���'��a�Dl*D������<��`����u��Qc��&D���ڝ}��M��aA�}�p�(e�%D�p� �N�L���^�
ܐI���!D���"��,e"����<D�@q�eZ�8�Pb�K��%2��$D���R����HwGI?ab0���'D����k~8,�h��04�g+'D� ����2�Bb�"����$D��IG*B)8�\��'�׃t�i"1�>D�$C���.� T*�S^�᪆�<D�R2釚3"�� &O\$g�>� $9D�t;�B�$-�6�5��<u�2�Z�5D��t������uᑸR �S'+1D������7�ũ������e�%0D�����
�K]�1�n�8�Aȏ(`!򄃓T�؝��a�?5a�1HP[;x?!��$��䛧�fz ��OڳW0!�dߛ?����X�\iT����\(40!�D
��642�m�"]UJ�E�	?*!�.�܄�
�'T^L*7�S�<�!��:Ί�����+O��rU���
�!�ޠt�"�93MVA4��k�%B�!�d�4I�Ԁ� *E�\�N�Q�*͐O�!�� ���""h�r�=W.����"Oh(02��I-��Ó��o�R�sP"O��V��`:d42T��K� �p"ODDk�ݪq� {���<
4�w"O0@@� ��I�F�A�x�
V"O���E�3��Y�&-OK��"Oje3F�M����  :L��"O��+U)Ӷ+͎�3H��q�"O��D�%Z&��u' k"�P5"O~���菼-��(�E��g؊-k@"O�����;D�-R�J1�>б�"O�|E�ڿ ��ꡊ�+��5�B"ODL{� ^�].<8ZV�$r�,#u"O��:S���<�R��"@&�^1"OH������~2���'��g0$ѡ�"OYC�a�����s��3.p"O�9҇�%����֥�F�!�r"O(�jB �)�0c�Ĺ1���Z�"O�-��EԂk�"�ɃBX� �~p�"O�Z��_(G�t]8w�E��<]��"ON��ԁ~aI�A@: ����"O2	H��T�t�c��I)����y҄�%L�W)\�9�F���S�y`��m�� ����' �8�@f��y���7���q��qoz1�%E�#�y���F�3C�b� RD��y�ΑRZBщ�"�X،��!��y���%V1� �d��K��p��)��yr6}{V<<4�`Jw�
�yR�9���U8g�p�8���y���+Y���3��4֚�zQ 
��y��/zY�"�㊖w�`� Nނ�y��k�����G��%��&���ȓy�Ȑ��E[�Ƞ�E�8�p��G����#Ƙ
�����_�h-�ȓF���[��"[.hp���:t��ȓ!O�0[��L�&�R��rƶP� y��-� ]!�К
���c�.*�L�ȓB>
Ѣ�A�H�x�d0�ȓ.Ԑ���]�%�����H֘�nɅȓ{F��'�F�mKшH�+]v�ȓC^t���IWRvā���6*d��4�XH�-J?X$� �l�!򄜼$H��;"��I�19�!�DT#5
�ih0��+<j�}YԨ�Be!�d�|06]� LC/)ZڔI �Y�T!�]�.����% 	�`L�x�qB�4K!�$ *�43G���h���U�v!�7x܌t �菀e���+T�2k!�0�ʼС�{�@�Bk�!!�Q����ڥ�=b���&�R�O!�$ɎK��)#�I½l*���6�!���?h�4Ai�.G>
��c�`�|�!�B4}�>eز�V�5���Q%o�!��20+�e(G�
?�j ���X�j�!�DPQ�V�ap/��l��IK#�1"�!�\-@HP��!	�u�Lar0�դI�!�=�Nq�Z��a����ҹ)A"O��4n�G��(� ��z۞Q��"Op-9���N(0/�R�Vd��"O�9�%�J}@ ���҄-�t�W"O`�ua�}d�Ks.Z7��,F"OL3�T�+�6p!�ĠB`>�"OԠ����,�B��X1���"O� .�&m�sp�򥦖��v��"O�y��ȏXq�ڲʌ�]w�0c5"Ov�S��a�R�C޾F:�q#"O��)ɖ.U���S#!x��z�"On5�6��^<Pca�Q�>�r���"Oy�O4^��h�!��֘xz"O����K;��4��ɇ�N��\yc"O��%t-^�rBbN�+�*ea"O*�LT�R�,` 3Duw�	��"O&d)�%���,3�"L?;i���"O��(��X!��K� �gEX��"O�cH��ih��Z )���"O�;ql�=���%��V����"O99âD	l$n9C����Љj�"OT�A�B��[�vQ�G(�/'�*�"O����J�'(m����q�t퐤"O>���b�$<��I �%,����p"O�����֡;<���f�	��s�"O`�81���zL	��@-TR8C!"O~�P@�hY�4�/]��ٻ�"OvȂ	� 6��5�Pm�@,P�cq"O2��-B:Z�@���,M���0f*O
T�7NL(u�yؕ��V���'�I`7B�0H��\�4�V'X���'�P5�@v�<rth�w�ٰ
�'|�m��8Аq���}{����'��#sg�QN@��6 ��h�\�
�'\��i��j��͋U)�^�D��	�'L0����V�f�PH�� �X�ThA	�'���H�fL�)�8�0��'�qP�$^v�:�K��X�{�	��'	���T(]R�v����@�}��L"�'���2���8$ ��طy��th�'����B=�I@�3{-`�2�'{0|D�K�v�j�˱$�!n��'���@�_�	(j)s���+sd,��'�Z= �J��y`�
vx��'�D����8U :e�烂�@d�, �'22P⤬"L��UY��$��R�'ܽ#p��Z|�ነ�'\�܉�
�'�,-9r�-���g�V�X)��	�'���Rր�6p�&����H9�
���'�>����R�XiO�'_x- �'r��D��F���i��6$L@�S�'c�X��m�*xHZ�!�.$��)��'�%��GP�^ �P� `�I�'>xѶ��$�V�U\�w���'�D��q���0��*��ܟz���'�D�"d�J�^�p���`I�{����'s�	Y0�Z.T$	B�؆w��+�'Y" ʃJ��r"��A"��q(pp)�'_��s�-!��F�,��9��f�H�<a@#G�$=��U��82��S�A�<��A?R�a��)F{.M�*v�<Q�g�@ݛd��h�頊�F�<a�-U�2c��6;��My�NF�<�Re״���B�4kf$я^X�<q���'i�d���/4ؼ ��y�<����X�����(`�,���as�<aGK _lȍ��ß�/��U���EF�<�߽~˴�h&�Ǜ;�b@$��I�<�aJ?-	(���ks�Ȳ	o�<�3��z.����ōJ�vuaW#j�<���U�	&�U�T��1�h�W%�g�<� F��	P�p@�pAɩDj�s�"O|t�SN�>(zz�ϋ�}*��{!"O�CӮ֯��`�&�p#rq�"O��q")V�qdM�VL#:��p*�"OnA�"�V[
C�	�#9L�"v"OX0��jY���I���Q2�(Q"O`�q�Ú�f�f-YA�[�8zj� A"O�q�gMΧ8��x�� �T�2�"O@��G�Z�!����f-��s��|q`"O��Z3�0z�F��,3���`�"O��9 �0Y�bPH0
I�b)��!v"O���΀i��\���F�hJ���"O ъ��5YII�viG�*P�P"O&�M�z���RK��+��Uy�"O.,9O���,T�a*B�9���(3"O��+�M��-҆�*��_���"O�S��b"M�G��&
�ةK�"O�-��+9�U�L<�|}rW"OBd�Ό�dq�� �#�w��x:#"O��Çƅ�D�*Cђ1�pE"Oش#�
��n�&���b[��<� �"O��k�n
�Sh��`�������"O\��v)� �`L���K1x�"O���b!�<(dQ���á&Jf��""O�Ȱ��6d��#c@M�d��"O �0�I%D~�4yb���&I����"O0ir�@>:MH�;���:FP��J>U�[�fZ@�ׇ_/(���G� �Is��H��ؿ ���dh��$�Sd,D�+#I�2�1��A�Y>>���H*D���2��~���r7n�D{"X��:D�XipoW8oT,���V9GC$HT�"D�L�B��dC���DG�ZQ�"h!D�	��\�ws����/< DFUyg<D��ڰ'��Y��1�Wb���P��9D��kv�_{O�����"v�i0 D;D���p&�����RE���SX�I�;D�x���@ӑ��$��}&%:D�����E#�@��Fj ��7D���r�ȸI�@�E$��$q�X�j)D�l4$T^f=�s�qa̐ң,+D�,RT�ޢ)t.���o�;��!�J<D�<pN_W�x���к]q�"��-D��r#�M>�ա6��Ιq�,1D�(���Fz@XU���"2����0D�@e��K�H��U��!o:��@g0D���ȅ'9�) LȌ4bABe�9D�Ȉr&��H�5
�ɣfЖQ8�*D��4��7U���CG�_^v:7�"D���Q�C'OBd8f�G�q�^���"D��A�d��7�^�f�œI*��+D�,��Ȟ%F��\(�<I24�v�+D�T��.B?�ʅ9��!��]���*D�I@���Mcp8Ql
(c�m�­+D�paA��
��ڶMC�N�녆&D��� ��{�^���xI��C��%D���S�:"T`�GBHDʖxX��#D���w�׺r��|92�Cn��@B D����G�P�2�Ƀe�*m�b09��9D���ॐ#c`�0�_$B��! �,D��2p�R!Q�,�CK�8r���B�.D�����sA�d��O��w�r�	Q@-�O^扦&C*- U��8}n���#F$�B�I�9"�U���%^H� ��a$NJ*B�)� �hِb.;�t`HŎ[%p?����"O��K���#}�䀨��ؠ/%\+"O��#fJ'7Jثfl�^k����"O�0���ߔs �K�EB���"OQxCJ@�U|mCscР[?��0��'��ę2Z�mc�˃�dqr�ǁl!�8 ID!H%�G�#�6`���7^i!�_�U�(�����g��8����3 T!�ӛ?)\5R%�R�)��� �,�);@!��;L��ta�����Ӳ!�x-!�d�1�`�%�W#uya���6!�$ڂ
3␫����M��F�SM�!���V]��q�M�DCE��4�!�$� )�U�D@@�E*���l�_�!�$K�[�h�t`�S��F�S-R�!�$?�419�ω'g��y�.��0O!�ϩ�81��5�hq��� >4!�䜉/�-��.Vs�� ZwN�4�!��.]��8��fM<t���jJ!�d��>J$@q�Оe&*|Jv����!�40��`@M	*1��bG��!�ye�xCtEі��i5��!�d�+�!���V*X��G.�!�$�# >����$O�%
��!����!���[��8 &#ʔT)t�20NGI�!�d�d��@���RR6Q.B-!��i�~%��S=rdp�a��{!!�ُ ����/� W2�8�EႤO�!��C�yu���Y� ͢�r�!�$�
U�5���4U�1#c!��fz!�dW���̓���6�PgFL�LR!��N[�`�S��C�5$��"E<B!�d	�z�֤��2:�죧.д"!�D�/�@qȀ��z��ر���&!��1k���e���)	��Q���h!�d�s
(`c��t�pDK O���!�Μ[��E���T/�:�j��&F�!��_1�Y�"�
�����I)\2!�d�7F��m�$dE!C�d
��>#!�d>r�S�
���!R�CK�,�!��hqN��Ǚ;��+�AI'�!�䗢P2J�ʇ"p�J\�&�Aw!��BDR��X5䃉n� ar�A!u\!�d,+�XH��\�N�D�/A!��|H�ep2��x)d(�sh��	!�O�*:�٣oG?]�diC�g��|!�X�K�T�
s� �xH�cu �!��7)0*�)��uXm�DϜ�R�!�$�%�DiS֣\�0A��3�!�䕥$����u#�b�|D�@1D?!�E�i{���Al��jД�J!m�q�!�[<C����#�S-2�.��P��#A�!򤇅6iD"� қE�L�Ӡ��6T!��i�|����$M	X��ԍ+!�ɑX�xE�`j@
=������D-!��� W \�#t�/B�Lq�ꓶT�!����t 1f��B��oݞE�!�D�2[K�y���\�2�.�.�!򄔟0�$屡���H�U�D�P3e�!�$G&,j��DP�*Ր��Eѱ+�!��Y)i���B�OwĬ��c�9?�!�d7P$f��c�\%5�!,�!��̚�p9@ѣ �6� ����ܰ:p!�d%�c�NR�*�Y�F�M�G2!�� ^q!Ro���V�`Fދ�$��G"O�i���ԚY�� �d�v�E)u"Ov%۰�P�\��u���Vjc�Ł�"OD��M.H�$���
�G���e"O��+�	�RUXq$��4=Cf���"O��k�$�0q�a���*B9�"O�=(�G�#a�ĵ�q�.!$���"O��Q��0�l�Ca����3"O4�֏=}�x�iPϝ	9N܋"O���I���2`��M�![��U�"O�I��ş�d�����-YG���"O�X2�M�;JL��jPM^����"Of}�t�,`x��Tn� O7Dy!�"ON�e@�"n@�MK��?���Z�"O�邶,
&�r�Q�JʇI���S"OX%��'� j���{%�ȠQ�q��"OFI�+֞&P�[�	�<=��%"O���$���/�*� ���57��y�"O������/k����&L��| F"O�i6�Z���S�(�1�q""OLI�CX	z���ق��Y�$�2"O�ay$�H<m�6���#F_�8,�G"O:���d2:���3N!;r�p�"O��)n��6)���2(�Qq� �"OT#�ʀ.4����_��e*!"O����_�u�UاJP�!��5)'"O�f��uB��"JZ͌A`#"O�]�u�Z�<O�90)�,Z� ��"O����c_�1��@%Wv���"O�,�Q�[!a �u;�A�_���T"O���/B> ڄ���D�.E:��0"Or}:U�C-d  ��( �^���"O����d��u�㑂_���Qa"O�]#U�Y�w�FE�S���*w�#"OR���	ɓ� e! �
&
����"O��(� 
E�g� �^��&"O���d���S���r�ޙ�
\AP"O��A�O�;��9hH��GЄ�y2�D7R=��@�5�e�&��:�y��
VYH��� -���� ���yR뀬x�t)�,�E^%���F��yr)U�%B���f2�r|`תX��y�M�4��M4�	ѫS�z.�"�'�>|*�G��B����0�Խw���y�'�]�פC�6����&)C�8(�
�'����&n]�Y�-�5�^7�:M@�'�Z-����I�Z�R��!5��<s�''��� 	m*Rt�uF��1M^��	�'��P�!�v��u�[V5~}"	�'�^IypC *���0�d�L����'�p�RD�
x@�i��֡I��x�'~@���ϧ �!Ee�?�j�'2TDy��<|�y#���L3d9�'}d�s �Y���h���-����'��͙ i�0{�J��G
=�z��	�'R�JT�ۆn�����ܩ7��Hi	�'�`)X©H +�`R�٧~�F�������G��1t�ƖA���{Bf7D�l����H�&15&Jp-��[�$5D�8 NT/L�T���C����%D��*�I���%�;m�����g��!�d��|� ��U��+:!��z�f�{�!��ۆ�䤠q���D��`ĩeY!�ā���Y;���#I��K�OI1p�!�� ��ě*�X<�Ǉ]�ל��"On5�W ��Q��� fV/�XB "OV�1�@�3V��%D�0�z�"O�	��ƁI7�qBe�,;���"O�pb�n[�Q ���6��9�<�"OZDPVʘ�dĢ�O_� �9�"O.d��e�NX���1	g"]�w"O^a�K��,�b��=jR@@��"Oh�Y ��4'����Jϖ93 �Q"O���U�V�.2l]� ߁`,B��"O^�r�� =Pz�8��b0p�`"On�'�@�f| ���y�R"O�X
$II��������)���H"O�A��	/i� �3�I	z�HP�"O�@3��N�X���ځ(H��v`i#"Oҹ����6���ggۏ}�A�"O��{GG�Z7}+�&�B��h""O�!2�KL$��ܡw/��J���y�"OL���G�\M��Z�냏��:Q"O�p�«�6�l��HC����"O0l��"��%��+�Hy�Eγ�yb!R�XpJ�x`��0"&�	z�e���yB$H�j->$ig�H��؉��Q�y2���b|��Ίvk���!Đ��y�eB9Y����B�"�QL�y�հ{N�;S��!@ �i(����y�e�@���*VP_ 1�0��y2N_�@|x��㩟Mh�yZ��=�yH��p�����>>�\�N���y.��P�#��3hL(c��yB#Q:iш1a˶��H�U��2�y�J m�^銀�Áj�Pa�#�U��y����f)#&�U"j������y"���+��8� ��I�����y"�E(l���ɱ$�8r�JA��@��y�j��8�~�Ca�	����I���y�!��\e���e�z�b�3�y2
7/� ��a��]�p(����yR*A�1��h%������07jP��yb�];|�� Ѩ�Y��چ�%�y�m�5��Uɢ��$�8e(�B
�y]d���)A�êuI�Ο!�yb�ۢ0�u�Y��|�J����y  ��Q�Kǐ�洨�K�y�	ȯ&x�Y�f��%/Üe+D�J��y"�G9Nt������(�T�3�W��yB��=x@ �3暬XTuB���y"g�B��SO� Q�,�Э���y����=��٩��	I�Xhjગ�y�&$ &�@@�,�')�vL���O,�yb���PjR}P��ׅ-��3�f��yRi��	ŀԨ hӬrg~�z&���y�K
p��)8B���ڴA"�^,�y�c��}����u��<':��`�ì�yҊ�>i��&�	2����GA��y������3s�ڵwx����N��yB��ܒ����qFI�P���yr���sFL�A�&�,i�R����y�I�$�.@�U�<VO,H�[4�y2�@��}���ѯ@Q�D�F���ybn�0|`,��g̱5K���1�yROJ<�~Ȣ#��:)�P����yBŪo�0�����Աf���y"�
 rQ�O�v�&�y���y
� ���Eɀ�dr�P�ń��A���r"O^M��Ō=C��@2�)?��Qp"O�L*���6
t�(e�؏s��0��"O��a��w���P�'6O{5"O�8 "�8����(��'v�0�u"OZ�2���?�؛��O�hX���"O:�it���Z��,��A@+^�i`"O"8F��plȽ��*^h�	�6"Odsge��h�I!��#GeHDXU"ODA��:X��@�����j D���ċ�Hդ���-��+�4D�諵N($�|8"զ��'�u->D��Q�N/�pEʠ@
t�����/D��y�g�,i)t .�^H��r� D����*��/"R5��*�x�)D�ty�U�Eo��	0��4zv]b�%D�tz�#2��ux�Lعo
V}�0N)D���f���j�"����� C	*J(D�@�%Q5{6���!?�uj��'D�\ۣ˟�P���z��ҥ� [�!#D�h����5��e�t+ޅKwG"D�L�pE�%�V�j�&�!M���`C$D���!+J.�Լ�!'�m�(��� D�ص��"�VT+�nȡ$�D �j<D��1��2�2�Z���c��ݫ$�$D�(��/��/�BIh�,EF�m�l!D�@���.(x�W�(Je���� D�ر �]�"�4���嘧lPr���+D��2��ƛu�T�BTH��4�š1)(D��Y��ü3/ܭЇ$��W��T%&D��+A�[.� Ta�GѬB'�?D�0X�	Đ?Z�N�p���D�<D��+$���L�� �1D  ��,D��飍�n��i�KĜ(	�Y�`�)D��e��*@8�j¢)w�mW�%D� �2�/,����K�d6 �e�7D�$�ѣ�A�t DG��%�����3D����W#�~��Ϙl��ej��1D������z&�����L�{�0D�b"�Y0�����6wF��	,D�|�&(��bdmj�FϑTFԸ���(D��{U�ΣmE�`5��}��D#TD(D��b%\1O߬�S�bԗGcrA���!D�W K.^�b]
p�0:D��Ue>D�,�P�S�h/�i�'������N;D�W	�@�4���IW�d�"�4D�LY�#�90���@��Ɔ>_@@zG�8D�� 1i �`f,�rƤF$B��:D�HjC���{�`M��ė2Y���>D����iV,9����VL�9]J�˧�<D�Q�
�',uܐ� �A!Pu:��9D�\�vFŜ)�@��.�?<[�8u�;D�҂���|r�d��X |�ah%D�$۱!��ET�����44��i��&D��-�5�$9����ބͩ&K%D�4�e�+��q�!\�:�b=�E"D��Z�k�r@�ag [�kh�+r*?D�Sȅ?uV��q�X�8Z����<D����Ć�$����m���  D��Q��#�ĉ�G@*8Q�,��<D�xh��2	<	 ��:(L|!Ӏ0D�\��W0$H�q,C�T��+;T��� �?��̃�� ��x�"O����ͫh�� �-�w\^S�<� ���V
K�s��׋�;� �k�"O��@��XB�Pc��S�c���Q"O�Q0��(7�feA��4|>�\j�"O�K���]r��XT�V�1A�"O��s��8z�� F_4O�@X�"O�̓R�@ i��8����#����"O�Q����M��	�#�!=?x�w"OH��B +� ���֬P2R5a"O$(�ҦT��T�h�Q )�$њ�"O6d�I�+nL�v��M���B"O&�KbH�6CA�=�v(ט�8�"O��&�t�<8Qw�ƀM��!��"OrIi�̉G&��eǌ�,��0"O@j�[�{�,��� WlT@u"O�8�u,�?��t��J�4�Fp"O4��#�� }D ��V�a�lQ2"O��P4�ӧ~W,���+j��U�0"O��Hq��e���9X�F\�!��PbH�J�S�H�i��!�J;��89B�1M�P�F�q�!�$��~R�q1�'�#5�*�5�\*&!�d^�E��mڶ�W�R���_�n!�$� R��X� m�(��Tzg�BX!��x��x�AL!'���F�^4!򄃀-0��u I1V��cC"i�!���?{�<���ҽ �v�s7��$m!��Ɏ[��E ���&s�E���T_^!��Hɞ킶��&/=�9��L/&!�DE8F�dՓ� I�A526*@�#!��ɌW��h\�so&�iC/�&G!�����Y$��FP"�I�,F�e�!�0�
)�d�F�@�pLQS��1�!��
BY�1-\�@n��S�B	,\(!�D������\�f�x��� ���!�DY�#�&����jN�uq6/�(i!�&��UrWI�%`a���:�f���h��Li�D� ��u��m��b�݇ȓK(t]K�����������^U���ȓi,<rp�BN�:Pj�o.����>����w�װ>�v��M������L�HY��O͍oP����g��3�����<F�Vi�: r�!��"_H5��nC&�P1l,�5
4M�RN�}�ȓfM�e� ���r_�y�"Š��_LAQ���X>q��z_����J�C  �:�p�+���LV�x�ȓ.�q�ӏ	�8[dl�^e�]�����6��&o�F<���Յi��ȓt�� �I�lk�d�'��$��D��O�n�#�`�>o�*���8R	�ȓ?G\���̠�E0S%ؘq��P��>�D��C�\)jv���A	S�Vx�ȓ;\�"7,I4f��e{Q:��Ʉ�kG:%�)G,%c�[�x�������j�.H5�p���&��r�C䉏J��m�&U�MXmy� ��B�	&Ȩ��)R(9S�����C�I}�-"J �-�j�3��͉�B�	6��%Y�ڨ/��U�EX�g�B�	)CL%ZA��-2,�x����y;�B��m�D�녃�-�nJlFffC�IBt��P�ٶ,�T0��.@%nC�IZ���u�H��6����ܢaTbC�Ʉ6���%o�:�&j�]�_�XC�)� \���� ��ٺ���$��YӀ"Olٙ�S�3D�Q�!"ڦ�P"O�)�-S�0���
uv �*�"O�xхC��W%F-��f�<>�H"O((���ښRs�ͱ�%Q03ک�"O���D�D�|����5n/2y��"O�d�o�9FL���Jӕp�p}�"O~5�m�s �i�%*��%���R�"O ���m8Rx��ri�4QZ2Ec2"Or���	E�0�{� =2�ْ�"O�ي�o��Yb(x���/�2�x�"O�lh��.�f8C2� %[�\��"O`���Ot,1	�`��9h�0��"Ont�ά"���1�*F+U�T���"O�MpL�
g[�툔���@#�"O�p ��,[�|���IP9�lc$"O83�a]546f�9����m-l�c"O�(�V�P0p�x{F�/Yt%�`"O.�9���^¤�R�­>\��"O��['�1the*����q-Р�"O�X��1l!6�r.�;xuh�"Od��a�$ShPH"!CY8=^!;E"O���D*�UN�� F��qh�u"O�H����m��Y�hۗt�l�C0"OҰ�2Q$4�@�g�Ոo���u"O��I��ȖkO����E:_�p!�v"O(9dlB?[3�P�v�U�Z9N)�g"ONX�b�;���!�^�z�5�'�����f�]��*�c޹���' ,z!dT
&����v����
�'�~�ZEڪLC���b싓gS<\�	�'���Қ=���0	F�b��@��'�2�[%�L&'?�X�鈼N���y�'�`:!�^�/
�0Q�T1p�*�b�'ޚ�6-T+�fl!Շ�&: �'j\ U̟��@����<Y@�C��x�/��$�ha`eR4D\\̘p�BӸ'/a{�&�.���u�;@��HΫ�y�IsN|w��7`&���J��yR@&WL$@�cf�[cT�0��3�yb��.
��1�遱*�V�:��M��yb�Z42��!�D�$W��d�m���yRA� [��]��dϱ�X��٤�y2 E�%<fm0�f٩e8��g��y�A�N�
��TIR�x3tt�eC<�y��3/����,�m�� @�['�y�)�#E���	�a�z%������y"펫'F��!V��]u���%�?D�`�����J�;���cK/j�2B�I+m�T[�� V°Z�d��|xB�I�/p�U�_<߸�����$�B��+'*\��"��8�\�$�C��v?�a��e�N����f�9k�B�	�,f���@�
9Ҁ���=:��B�	��V�� ��D7|��1��=e�B�ɛtvPx�̊?���9���1f1�B��%��ݙv'(
�Rd� ���B��:�8A��#� �K`H ZB��)*ۓAI�ge��(6B��<�8B�ɭv!�U������Aa�N���"B�	
ʴRcH�6���a��w�B��N ��Y�)�A���O;X��C��	1�R�9��F,L�Z�ॡ�#��C�5�TSs)�NYx�X� o�B�)� �x!B�;ڨ鈕+����k "Op	����= ��\�,G$�z1�"O|��u�^W��c��W���0"O�1R�e۳GO�h1���p*��"OJ$r��ï)�l5����X�,aP"O��R���ހ�����	%fل*O��Y4 ��+�+|R���'�(�YR"�Etڀ��_�8]x�'Z(�ڀ-�2;��Dq�J�oHv��'ɒ�h���,��0�`$2���'Ld�4p4�`g`^.R��I�	�'�:a�cDH�@`�&�E����	�',j�J�
_�%���K0�S�O��=E�$m�*5���2��R����%���yrG�$���Jd8���n֩�yBN�P�� z���QӴ��&L:�yZcb�إ$ܸu���z�����y"�P�<�hɒ4O�l��)�����yB�ϛV����񇅋_�qa�
�0�yRaW�Yx(D�'cȬ)(���aI��y��͏N���D�V�U� �����y�H̞2r�&O��;V�@���y"�@���)�1h�>7瀱	C*G��y��+sA>5�sF��.L���'�y�h��� �����5y�V�aA!Ǻ�y2��.6dT"rʢ&��HZ!�J�y"�ȶ9���hgP��4��
P��yb�^��Јe+V
D�V�����y"�F-h��TF�:��Л�W/�y���	8=���*�0.��dApZ��y�K�1�12t
F�*n�@`���y�ݖ/�Ps�ė�[�T�@���y��Rvx�pe�%f��(&��y2�3a	��BF�"pգ���,���?�S�O���k�U�y�Љ��DI�f�DP�'�\�
T�G�ij� b���Xg��Z�'@�}���j�N�9�gү{J�q�'��=�%B�#e�.27�V٦T��'�]��fʶoZ�2$C:ب�k�',��3�3	�e@�LH�	��%��'�,)���n�J�Dj�P���']�aڕj�44�>1гh�N#qy�'�
tZ �� p�!�#�����'��CI�+Pp("R�Z�ݐ�'��@Z&OH3t��ja��-u� 2�'� 1Y"���{@`����$\�܈Q�'ZVh
B��+��M�&%S�W��8
�'	����&��A{XQ
F*�%d�(Ap	�'=�ę6J�	&�tuSu	�/	���A	�'Mn!�DH���e�AL��� 1r�'p ��U��-Eg؁1�'^�Z��b�'�bl��(2y3�mH U�Ƥ�
�'���QP��>�2بw#ܥ0��
�'$j�P$NŇA�����xVz��'t���Ѓ4� x�R��t�]��'T,��"N��h	�8:�E�f*�8��'�*��Z�U������[c����'��;�N�&y\i�EM�<LL��
�'�a{���-c��"�_�H���'�F�!�|f�`�s/
�;ּ)8�'/f�jgCα!���	�fS07P]�'�:��dH-G�❑����!�|�C�'�v��O^�l��9b ��Ћ�'Szt��L6I�\��O[�K��	��� ��'�ɜx��!QA�
niq"O�40ea7 ��� ���� �#�"O�2���+y�B��B�HZDw*O��`$
%�J3�ޣ'|f�
�'�V��'�W�A�~�v�v0��'q��A�(��x��t����'ڈ��D�m��Bw�ߛu���'<C��;��a��8�4��'�X]�oG6F���h$��-��'G`t ��ΏV�Ppcu���T`�'�N��C���~ʐd#�IN�	���A�'}V��g,��v���zT� �ļ]��'��D��oX�d�T�Ӄ��$10�!��'���a�8b�K�h�/v�Q�'><x�Cgc��2��+t	��'`pX��	1���:�
�.�D[�'}����F�J\��Kϼbr��'�ܨ�B̉#�$�C�j �ī�'y� �Wh\�[6P?c� �
�'X�i'Iބ@Z�Tqf�ɮeh��(
�'^T�J��ɋ@�v�ytK���B
�';Р0���"-����Ğ�(���'^���ѧC�R�I�Epo���
�'� �r��Re_j�څÖ4a��\8
�'{I�`Q'�ݪU��&`ּa��'X�e�*� |�9jp���
�6("�'Q����d˞L2�#@#T���
�'��b!iS$H����}"�z�'$`���8 G�(�f�aX`2�'}X��&#Ct�P�w�^5�Y�';�Dx6 K�mИTi��S�1��`�'D�hb�U�W�䬠�[�1Ԕ ;
�'|���T�_�C�<�RA�"W��[�'�,�	����_!�\Z�"I� ��'c�	K�?���Q�`��r�'1�LI#�\Z��0b)D>T��'���ص�ރ$�\�;%�*/>�p1�����E���;�C�d�(�j��:h�!�dT(Xyޑ�_�@��$R�i��L�!�D�K�n��e��I�^�Cv���?�!�[#XX�0!ZaѨ�	��)���'�D��%$�/�(�tG*�x�'�Q��O�1�������Z�p���'��]��ؠ2��k �JT���'h����W}�>%��+�"B���
�'��$�����'G�Z���'�,5	��$g��ڔ�=����'B��1���
C���@��u�B��'gt8����Ka<X#�	'��L9
�'������"c� ɷ��*���'�Ir��"d�0HA䪒	
WҨ��'�r�kƌB�3��*t�v_n��'��9z�!�=���tG̅\J�'L>�PR�h��  ��V1�. �
�'U�,R�شEo��s�9 ��'�a��	o����V�U�V��q1�'��AZB�=t�֮�N���y"➊.�&�����3X �X�s#���O�X�dF�N�d	�s/:������X�LL�	 Q��j�<�ǯ��t:�b�q�*-�&X?Q��S!x^�sf	��4�����iM22���LJ�x��"��m!�(�b���I�7g��
a��2VF��2k��/���hS昩�9C%�?#<q0�H�]�D�̖=�$$�3�{x� ���;���`âB>$f��w�K�c^`�#��4) ��ֈ|5�Є��(1ޮ��T��|"2ycbDߜ?�"=�p$Tm�^E�"��?��%���GD�� >X����'x�"#'ς�@,`"O���dˀ�(O��� ��&Zxl�1�(H�Q���D��d��5V!_�B,�ePQhW�*Kt�Sf�^�y�@Uy�D�؂�['+����e.���ybĉ-:�qFx��S�8E
<0�g�޶<��˕+p������^����9� ]�/<'��j �U�n�O�z0�'������w�	Jr�'2,YЎR�E�
��>y{��ƎBu�9�zvd[篗�)�T��w�HaeE�%��`C!`�O"Tc7!�U�����
���'R���k͟:\p�����6g�&��"O��㋎�ENd\[u�K� ̼�xb�'��y��'9�ic�������#	T�\�Y�	�:�H%��O1{� 'j8�a�D m��RE"O褃��ɮ(���S���/�*����`Ǝ��F�v���S+S�G���2"�i�!���m�`�C�� 3�ra@ä�����&��3�g?�6�L�^�49j��Y;Ra�p��GZ�<�gkO�zc=��ۭi_�,����ϟ��w�Qr��xB�0>����%�פJ�z��Ӡ%|OzA�$j7?7
�<�6���Q�I�<���:{�X��4�ݔ>�E)���B��)8�bç) �Q��L�y٨�XW�Uka�d�ȓ$b0�
�	��㑤J#�8���a��h�����6�>(��H�{x��h�	�;��D��E�U�8�c�6X�����Ҩ�yr��>���4BՈ����y��)�]�
$@BT�[��8H���"�����r|���cmO�\Y�$���X�Q
���'��}��O[����V��\�l%�����0?Q(O��/U�ܘQ�W�^y1WE��y2�E�"�1��^5D�Xy)vc�ՈO�z���m��ūĘ!�f$s��M�<9�fχVx� �B�b�x �(NM�<�g��4 uH��'h��NܠI�$FH�<a��½@F���g֐�*��.�H�<EI�!��=���_��3"F�<���O=Q%歊�.ޅel�%�A�x�<��pb�A���>m ���h�y�<�ҥďb����w2
�c��q�<ADL�$;��)��ɂ)3��l��B�g�<��E��)#qB��H�H�@�Ɠ`�<y'��q
�iS%
�#m��Q&�^V�<I�K�;c���I�B�nxX��S�<�� �c��*bod	��ʽ��B�& f����E�0�|1�+M;E��B��7��%�L		Up��3Bɳt7jB䉍B�be�p��0�0�k��M2��C�I�t�X��E
<�z8#G��+�NC�I+Y����
/ h�0��@�C�ɟ�T�K�N��R|�1P!Y�[��C�0n��`1��b���$մ9�FC�ɯc"Epw�S�]O�� �=+�C�ɮ@�8Tsr�\�G<L���	o�B�I6f�}��F�1�X�v��;W"B�I�:%r�y�D�'L�{�Lϙ�B�ɪ{y���F�A���9cN�y��C�82�@��Ԉ"
���)�HV"H �C�1(��	� d��)d�C��) F��$��%�V�����GF`B䉰6���X����b�(���ɔe�zB�ɻ1�|�W��:���̚�b8B�I�.� q��`���z�"5��*�HC�IUb���E�kh�y�tԔml:C�I�*�R1��
E�	��)Ԯ�3��B�)� �x㒀\�ƒ����b'���&"O�@�ӻZ>qhT�K0|�^��1"O"�MT�bYE�O 4E��"O��{Ӎ^0U��z5� pQ�0��"O ]�'N 3�>�Y�hF�e0�<q�"O�h�Ҹ`�T�H�_�>ȹs�"O�es`/�7>�6H	b�ϰ~��(�"OP��`�
-�.1CH:��]{'"Oiѣ\�kF��s����+�J���"Oe�J]�7�F�Q1(��I�೔"O�=����w�EW��jX�ls"O����jI0�Ԥyct0e"O����`�30�4�C� r��In<D� ��ُ6G舙�ȿBVЕ��,�O�˓!�F��`&��0��@4��x�ʰ��a�����c����7�P�
��F|2���g��ы��^<|!c��7#$B�* �Aᭂ�.74��Q��P���IT����H�"#�
O@F���[�p0"O(��"mă7N��(�J��Y��"O,0�_?P~�/��<x)�E�ɡE��Pp�a��� �z��u����$�ՃA�����CL�<9�O
J�.��%	�Q}d)��,��b� ��4��[�8	�g�O@�D��O����R��n�(P �+ln��0"O��'!��i���s�Uӣ�y�����H)��؅1<ax2/I���� ���8��0=	�&ʇMP�W"�{M�lp���5��4�$��P�ve�d��F�:�X�Y�UR��Q��qi�l�z,�%�ty��&СUj�$F��1�j��ȉO�<0U��5D��ઁ��?V� �)
�'T4�K�M�5Ӯ8	�������ӿG��1iS-
m�0��!��O7J�r�O�U�W�M <@�0���.�F��$
O���2��!'9���M�Wn�zVES.8� R��k�z�x��dS>��(����O�p�)ѮP�q��.��Jq@�'�FA���κcF�jE�9Re��!D W��l�*�B�{���8�0�(�j!�0?Y��H:��%)��U�.�2�)s~Bn��;��E��R�b�1w/^� �^ȋ�Y^���#E}��Z���%W(���b� PC��"d�ݒT�5Q� 1�B��Z��_/L�yC�Q�)�r�� �b�S*�x��Mu�y1��Ґ�A�ѯdV(Y
Ea2�|!㏎3d�F�����¼����U�9S��Թ4`���J).���'%�2g�H�G{�d�kW��ABS�=�Pmq���0<�"�Ύ�́%*J![��|��B7)ʜ4`�8Y�RYA�� � ��",ɂD�ƍ��P��Xr�H�r>]Y�+�S&�`�'�l��"�
�X����ڞM���A�(-tu�PZ>�;�Ԕw���ҭ�<STZw,=D��S�E����T���j�g��>>D �@J�IBTc�J��7�&?=#�A+5{��]38�9�����g�T-��b{�4B�ɳ<��{%Nt�t1����Ν���V�r=��V <P	�@��-��CUNWS�'�|W(j]b�@���Q�2ť�X�R�@�Qմ�pW`�4�$��O��?G��)�`��#U��0�$��C��3�H	��`D�c[� ����`��M?}n�Ȥ��X���'�:�(�4Z�8�QC��ʑ�7���M�5[>��D�>����VgD�'+z�x�b3�hF@�Q�)�JqH�ģ�.H��C�cͧ�H��gA�H0B�� ڽA7�t� �T���'E?�l�`n�뼛"��*`;�pP�ٹXlb��vS�+刐Zƃ1�)�')����b/�?$+j�4D�eD��g�,���"�OXV�椛+5v�0��>�hO�9�5A�]��
}�
lV�$��A��{���U�*�ف�<J�hH������OܦtvH$�g Q0�Y�����I��aZw�	�F�^�[D�O�<)�GVb�t�дi|���@����l� k�� ;e��#��b�l�M�
�͏q�D�޸US�2Q�S�*D M#�0�(O$ �r�>�T_��E����8<�AғI:@z���_�j�os.!i�D�eܧ:���h��r��b�/�h�Es�F�!-7���$+,�4�7K	�N�4��k/�����=��X�� /J�f������\M�+	� K��"�K%|���Ƃ.���h�� ,OH�Xq���_9�탡,C \��D8ǉR.Ix>�"gd?P[X�d,Wq� 邤�#�O�d�Q �:�"�o�U�&}aO>��/̜W�,iIg)·*����.����L2��O,A'@�K�C�	V>>�#"O� �AN:b���0��(��px�E/���6
Z!�6�Aό�\>��'c�u�	��}@:u���\�CO@!�	�'�8�vd� j��&@Q>�1����hEP͙A �hI�s�3�0<�ϑ�RfH���(<3�����f؞��'�~�RT��I#lkPU�C-��4�,�w❧L����&e(<�e�"z�Pe�EB�!,sHG�'a���cJ�D����D�	�G����� ��-��3�bB��|����d��JȕJ`�(^hu
��ҥ)+!��6K>H�f�R\6A��͖�tQ�\C�!ʶ˨�D�(d�(dmΌ��JM� b���:O\�J��'�00�� �+VzL�9E�Ѓ)V��B	�'y�G'̮;���S�&�c�xTik�}u���&�lم��B0����W�*^A�ȓ ��rս"N�Yń%DLj���g���c�0�J%�G,��bh�T�ȓ`�j�4�Q9���Pe��+)ḣȓF�Z�+É�;k��Ԛ�)֪<�9�ȓ!�̝��q�<咄��mI&��o�Ab�/(XB�ZtdG�0�x��ȓH\xl
'�ȜQ���XA�Wl\-��Vc@���̚st��PM�UjlU��>�Z]����*�M�+�e�.��ȓ&`��C`�rրs$W.{6���>�H�+�Z;~u"����H�}��ȓ���g�������J�ȓAq|@Q��9y��s�ĲZl�B��":e���!N��ta@0(6 =fC䉕
&�d�T63x���咺�bC䉇5�(���hG}k �fk��S��C�$�4ı�mL�O�| ���:Q4B�ɣ$���"�C4�dE�!@C���y�g��#'����A$
�����	�y��'�J�3Q�F $@���y@H�A&RM
)��n� ���/�yBGH%�^��"�O;d���č�!�yB��?��@DI h>�r��#�y	W�g�P+�.3K�-��N��y!D�I��p��iK!0)�����y"�t2����fX�� NN.�yRi�o����fi�Ӿj(	��y��ptrtQq	F*~?�Q�� G��y��T�$8�c�Zd߰�Q�
��y"kX�[��y�V+V4P-j	���,�ya�6�rh���	8T�L�w�T�yr�E5��
3���%n��K2����_�q�4 � r�0U{�"��koȸ��i]j$J�'܍��E+kn�1��3�a@@|�!؇� sS��ȓ3�d4RrBM�<��A ��
#�Ā�ȓu������]���}��۞K>��ȓ�>8�eS-��Փu�Q6�(�ȓX�	�`Q�5�:�s�$M�S1>Ąȓ;�A��� 't�dS��۪mipy�ȓa8h�f��!IfV(� ��c�<�ȓ0�4 �V�R3^�H���l�i�R���Z�l�@�ʝ�v��( ��p���2 "pf�n�։peKB�Q!^���+ϔ9y`��R�i�*��yh|�ȓN�<q0��4kS���b�I�I��QD�"���HsK�*�F�fL�ȓP3"�B AM�0D(�e�����܆�V*��Kw��4�.,���6΁��B��R匘ylX�&n3��A�ȓY����놂 `"]��A0C��L��S�? .���eɚq]48�.��#]`�T"OF��PA[�PZ8\0j_�b���HF"OZ�,ٜ>����=Ά ��"O^h��I�S�B`������`Q"O��c�'�1�����F�?G D̪d"O��+r#�� ��
A� �,ͪ"O<�REo�F�Xt�'��>W�u"OP�5#K�u��5P@;@~���"O�L�g��y���!�*�;) ��Z"O�A1�偷8 ��r���5)Hb�"O`��ń������î{~^���"O| QFo@	�^���'�PhF�*p"O���-b�8jS�%*�� �"Oj�&�O,J�
��ጲ#��� "O:a�&�D~��ږV}6"O��"�����
�%ݨ*άK�"Ox`���� �(�A�A�1
�"O���*��-QM�_��Ж"O.�iF�H(9wdЍ$j� D"O�M�V�����1�� C�"O�,S�G�0�2����"�ke"O�xb�CC���+@��<𠠇"On9���w�}�A��;u ƥ��"O,�{V
'_�4D�4��!/Dp�6"Or`C�Nکyk������K���t"O���B�m�ԁ �l��^Ұ8+�"O���'�	.a\�	��	�X�"O�9�B��3#�`� ���q)�\��"O�;��}��@�2a��� K�"O������Q�>�[F�������"O��` $A0M���;�*��,n��ہ"O�)��tp}�	Y4	DV�V"O�m�����q^�A�Gj�Z3"%��"O�X���+`Nl��&)�	w7�2A"O����Ѿ0�z`B��$ja@"O���u,�'N�d�c"�U�`��P�"O�XG�4Մxi�㖟)�����"O���K�n�\80BLK���;"O�]�`)ɺY�l�Q��(kSL��P"O�`�@�-�ڭ@�-;adЃ�"O&�	����0t�� VKR$]q�d"O���7NW�~ª����{��՚F"O���M$6��)ǩ�,}���4"O\0a�L�ޔ:�b���3�"Oj�k�$Ҕy�"d 'S�:�ݣ "O��:U�)3��̋�Vt��!"s"O$���N�  �J�A�ٳ#Z�`�S"O>�����8p�Jh���*_4 �"Ot���$�zS/P�r>*HСß��y"�j}v!�pb�4'�j������y�4��$`�L�>r�tۓ����yR*X?B8��Z���wh\3��=�y ��&����"B��x��a�$$�y��@�B[r5c3IM�y����R���y�m��i>�:�c�L����G�;�y�S�P(J �B�"�僀g��y"��@pq��%�Q)W���ȓ|4P�cL�DH	�5	=C�	4)�	h���l"n��B�I(� ���۝'i�}���'U�B�I=���#Im�y�FͰ �C䉶A�=E��(���Ya��u	�C��2O<��`Cf�,���@ThF� O<C�	�=��%j��hNxM�$��A�8C�)� �)jcg�=4P�*��Нw52�"O�m�2^�c��3 �h\;�"OD(� ���4���[gN5/�
�8�"O�љ��]260X���כ�x��"O���QL !_������c����C"Of`rP�[�f1p�W"�I��"O�D!��8-��Qt�3F�(��"O���� �|H�}q�+�	=�� �"OF� �A�m��%�B�w�\#!"O�|A�i�"w�X5B4�\�7�� �0"Ohh���'g����ЎZO*@�w"O�I	��27���إ��;�"O@#��T�J {a��D�d%p"O��!�D�t�XIs��Yw�Y#p"O2(���<{�$ȆF�5M8Yv"OF�k�$L�C��QQ%Y2pT��(A"O���b�ۿ
�P�4E�N^�,�"O"\���1EN�S�ʦX�l}��"O��"5�e��A���͋h�Q;r"O���$�!�z��䎞L�n�a"O:���-�!+���� ��3�,Y�V"OP`j��9٢�
U�T/ʊ��"O>����9�j���*����v"O*�cF�;>�J&).|��Y`D"O4�ƀΪ�*Ib�IҾcd�LrC"O�Y��J?�H�"n_�Q[r�Q"O<�L��L�v`�<-[8}Aw"O��PO�dg0��R
v:DQ�"O�|�F��x��m�߉B��q"O�A�$a^4y���.�9z��ii�"O��`�m�Hڌ �t�\�U� ���"OV�kSNI3S6�#��FP�B�a'"O��`)@q�\Q�!C�)�� 3"O8a�����6"0R�oN�g�P�!W"O�����B�C�OFn�XX�"Op)�/��6N���-�4�Y`�"O�-��G�n�L�c�+k�
]�G"O�P�0DT`B�ˌ-"�F�S"Ot<���&m�(����`�i�"O�d��F�Ͱ���E��x"O�4{�ւ!�V�ZfƇ4s�� V"O�-�q�رW��1WoԌKU�(��"On��ҫ�d���
��(3����"O�P�B�����I�4*J��0"OL ��F�|��y�&Ԛst!b"OJ��D`� r�����J�5�¹��"O� ��g�>$�鳆�ߗdiT�u"O�M[�l�,x�L9m�>vS���&"O0* %�t�0�'܂PXAh�"O�}�w��J���4�U�K%d!C�"O���D8�@�I 2���"O���E㌫O�8QH!B��\@�#"O*��)��BE�􁒦e�He	�"O�!xtO�C�l,�g�#�qI�"O&q��&�]1F��
(>�n�``"O�݋�Ό�h�@8:�iW�i��D�"O�k7��m�H�h�h�;^��Sd"O����>n�4��ơW0m��qa"O�Q�Wf�<^�����ٷg���K�"Ohl�tjҷc&����Nb��8`p"O�@SA�& �Aad��B��!z2"OP�Y���9!��̃��]�L� Y�b"O���7�_� BL�C@�/}�0q�"OnQE�*��y�n#
@<�0"O� X��L�Sм�q�����Tá"O���F
K�|�r^�L�<q�"O����i�4�
�Y��}�7N!D�LH��D��4��"64�Xjv�>D����O-��%�A;�ޔh4�>D��3�ƛ9�$�ˇFޛk����D:D��K�ć����1#�J�j�X$L9D�$*�����x��,�))��:D� �Al��5L�Q�H�=b��y�5g6D�X3' ů4z���7��	��&4D����$7f�H��_�4�����5D�l��ΔB�X��j�1h���,D�� f��)j�Jy�6-بRc�l7�(D�A6"�#9n �b R�.��v�=D�$)�%؋<d�r�mP�9���(�A<D�|�"ԓ �2)�� ѳp�b�`�4D���FdSXzd����NH�f�4D���� xTPR5�@ �zb�0D�Ђ�L����r�'_>�>�Xt�0D�Y�g!f�k�B�Q�F-۵�,D��"4�n�*�B}� E��,D�4R2���NnHJᄨ8k�\C&/(D��U��>;L�RA,&P��Ӱ�:D�k��T��$zUj��3�Vt@.*D����g�Q����U#�Ew`)��K<D�0(��<ԉ�5�T���x�*:D�����CZ�<�+�lؤom�xC0,;D�pH��U��a���UZ��"�+6D�D�4K��h��\z���*	�8�P#7D���/7�ȁ����F�R�k2� D��1�ѽ>�j���c��W���2Ī3D��GfɉspԠqBG�)�2�"D��b+�|�����T.�a�%D�@��̎|�y��ӎ7�����.-D��%o�7w���(A�Z�\���2�`.D�8d�P3����L�@��K.D��aQ�ڟ.�V��W6p!�lJGe8D�p���ܒ��2��W1�� ���6D��ԣP7|;��C�*S#X��Ъ2D�����V��Cd"CѮ-	��$D� ؒM,h�FB#q<T�3�D"D���/�>!䑪҂��j5RT��$D�8R��~�P����I�*T`�d%D��s���c���U&��.��9�y� Hf�Vj����_�F1��qI=�w�� �JF�)�����U�T���[��|�SmR(86�l���E#��0�%(��;�$��s���;9�vd2�)�ӛy�H$
E	��L�H�s��­{-��'�\�����i��$I���}��@�r�&~q�dJ,m�⟢}�@Ȑ01�Z��g�#dL!ڱJ��C���r8��D���J�J&�6^iڕ#��{>5�D�Ȭ}�	�����ʄK�M&�	qd���?%?�I1��L��;��53lA@��(}bď�6k�O���S� V:3�̼�aB��="��OН�u�5�)ڧ28x���uoj���/�՚�*���|��O�?AR�E�>*��W�@¦�T���'�����S�t�\�#ӧC#�<D [�;��*���]�S�>� &&��5�X��NՂ�'j�����i���v����[9%Lѐ��%���U��㟢}�u�[ �t����,L(���B[��!���?m�~�c�\>5��b� ^�J��z���:g�O�Tç`�:�%#%Xg�t3VO�(�H��=��jG�����'a�~��
�/3�~P�5͉)i~D�O����K&�)�4GEc�ǘ
94�iy��C�9fd�I<�V��?E�t��29ZN�&�ކY�X%�ŀ��L�^)���4�)�g�? ��;�k�v�Fyi�k�-p�$��m�|�����I�+;��,�m\�U��yYp�M��qO�(l�ا�	�(Ww-��*�8d���b�_5-8����#D�L)�ə>�F�	q��`@�Z� D�T���]\1����i�聹�:D��B�׎(h�7����鲴�9D��t@�C͈k�����p3�8D��d�@,z���ě�:_�â�!D���ы�R��@2MXX�t����:D��i��8n�8d!X" 0i5D��nӈ�3ʖ0c-���'>D��I��E�C|���i:E/~Ԣ1k;D��r�ʇ`���gF��{ɰ�#Ŧ9D�41V�/n`��A�e����E9D��
� M�C��થD�4ʎA���<D���΄��pqI�
�]!x1s�8D��yTϊ�w"��*
�dz@�SF�8D� �'��j�v��o͠O�؝��#,D�T� e���K��ſS��EIGN>D���C�Ǯ%�L̀v���x�J|��<D��� �P<#Ğ�e�#F�<�g�.D�X��Q/om,�Y���'\$	fL,D��Fϻ@n3��L�A>��+D��Qs1(t�����~�(�P��.D�@�����8�#'a�Lw$�c��*D��Y'Ę� ����Rr�<���;D����ۘG�n�u��<@d�7D�L���̩
= ��E�;r+�$�%4D��0Q�^�t۔� �DS�I�d�D*O.���'�j5�%�).�t"O}��O���I殐�c���$"O�j���4�T��';X�#"O�<cF��vq2UQ����9:�"O��G	V�lV��0ā�g�n�0a"O��u�ÿg�|8x%CO�$�r@3�"O~��ԉ�OD�3A��<���"O�1�ҘbǪ#��ҏO�BqZ�"O!Zg�4" }(��X7����"O~�3匓"�,R�M�;�����"O�"�î	�����,��R��5"O�-�Â�n�$�D�!��p3R"O��9�#�5c̐��뚣M̘4 �"O\���/�;�2����#G�4Y@�"O. ���Y�n��q5� �y����"O)�'���#�&�a�/4Y��"O�1'���g��� CA4n��@p"O��+uJ���c�j�U񪭰�"OB�6�%gQV ��"�ư"OR	:�F�g�h��$J�
�lc�"OR��S���.-t�i')J�R1Z�"O�m#��W�(S7i��5����"O�t�R�ܪG4X �T�G01�d�{�"O0�sF�A�i3\�����/]%��"OT1J���SI����X�;�}�"O�i� %ـv�[� �_>
AR�"O<�rp�W>��Tk�*L	��Q"O�!9��ۿ	Ԋ���($p���R"O��X�y�p'�P�C<�P�"On���K��=Q�d]�J*`���"O�=���&q�2�` �C  ��uK�"O�Tf�܄���"#��S"ՁA"O�x�-�;���{$*��XՊر"O���B��>�(��*c���R&"Ot�9��c���r��5���"O� ���b��������j��ix�"O��F�اtX*�"�E�#S���B"O0U������.�P��4�"O|1:��ߝr�f\*�W8/�Z���"O ;��>B]J�@��<J����"Ob���)�8",�yR6!T�kĴ��"O���g���m����נg\0�YS"Oxqz�%��Q$�3���DR�E�"O�I�тD)O�H��cC$Qj��"O���Ώ�=?DR#��vC��3"O\YI����$�ތ�Q"O����Q4&\�����
8"O��$�BY��8��FaL���'�`�����w��8W8+�����'�Zy�S�T'i#�ԉQ��+r�(��'6p�AF�
"y�zi�Ð���="�'6��r�n�!L��8
���vxq��'A� �"���5 ���'?z]�m��'�N�p������,��o�����'k�ű�K�%�[�JD�T��	�'eĩXeU���y`e:�'!��rSarH�'�1gf5��'������<��8s�bJ��R��
�'h��5U�Xz��/y����'愄
�Ş!d~��u2wSn}K�'��}��+R�p��+�#Y:Wh�+�'Va�G�\��
�M[�p̔��v"O�(�s�M5Z�c�X
W�Ȁ�"O�qǕ#�,i`%%ڣoH�ԡr"O��I���'\6�`$�J�hM+�"O �[�	��^��땨ĭ:�P��"O�p@�iCI�=qҘ��"OfqI *U�n萶�G8^
.�w"O|sGI:I�����F�T�����"O.��e��fo���EѤp�Zd6"O�(��)C
<�zaO�5҂`�"O���C×u�$C�nY[>8r"Oā��ݲ9= �M�y��P"�"O���aN��A@�L�N6�la�"O�y���
99�+̺U@&��d"OR�+����	 ���]:�m"OL1��@����3�ݼ �d)��"O��N��?��p!��ʓ? ���g"O�|�j=�hd�� �4b���"O����χ�j�t�K��ʛ<'T�3"O� BQ8U�,����W=�J0"$"O�� � ݩmh<�B�F3]چ@p"O�9م�_�/g��4��!3͢9�&"O����]>T��\��[�,��aYV"O�EZ�`^�=Tm;rL.K�
�"O��U琈2�P���F�Q�� Q�"O��h3��t(X%���A����"O0�z����j4DK��^"{��0�"O$��r
����Qq�FR�;t�x��"O<� *_�eJ�s]�	�x��"O\ؐ���]��ؓ���|��"OԠ:����Fp���e�0Z��G/�!�-Gh�P�@ȌW ؉�l^�!�D�4� q��];AntpKĞDR!��ߌ#&�Y��L��u����$�ǑEX!�1WQ~l�DD�!���G3z=!�܁:7t����9/�t�E�[.!�$WtU`�˲��c��Y�TbZ1y!�X�l�H��$ۄ&�Rq�3��|!�� ��B�� �~���l #l���0"OR��-�����~�Ju"OHP���33� �r˖����"O���W�	.N��SD�L��I��"O���D��s=Fĩ���� �b�"O6����:ܲ�JC�1�`Q�"O�1`��@ۆ��"N	LpC"O��B���`3�p���F��f"O<�%C�>>R�����
��Ë�y�
:Y��̱|f�=@�.�yb���$#@)ڥ�V�(sb��di�y�(�#
�(�`*�!s�H�!��yr"�;X����
�q�6��rf���y�h�:	�TU(��	�j��yk�$���y2��*�0K�	E�c{���` �����p>��ٖn�s4
�._|��U�<��al���kր�#�-K�R�<A�$�ep� S��q�xKac�b�<���NH���kK�B��D��(Ui�<d]"��1�Qp�)cDc�d�<�s�G�H�j���$L�I�Z����L`�<!tI�;?��2���@ Th0�F�<qQ��7(z�!d�I��i ��}�<�1.
H��9���
�PvD�qQ�@v�<Iue���8�dB~���$�Eo�<q!�ŵ/�n����&Ȳ�A�Bj�<���'lo��H�̎Zj�q���c�<u��0�|�YN0+էƿ\T!�1!!<5Q�́�j9�X��dB*s;!�$��w�>�Zq��#N*��4c�7t,!�dT�a����QC��Ϧ�Ջ�7<!��֏c����n*E�J��\8!�J3kL�u�"�qC�}y��G�R�!��׈)-.��J�#j'�C&�u�!�A&F.���}4��q��Q�!���8�p����8��Ň!�!�D%]���Rꍡj�6u��X?�!�$�f�6��E(S�vT�tC��!�d�z_�T{��(y,h�B:a�!�Ԧl2 ���[���à�0W�!�=M�������$$�(�F ϡ;!���E.��Q@,ݥD��h�e�@�T�!� �}JRd���|�p�4�X�!�O0vV�Pf��*@oڷz!��\�7(hzv.����� D��|�!�D�$���P�ď�C�A�]=MM!�D�V�ve��`�0�8�Q�K!�N��2{�o�
2r�Ӱ�� @0!��T1v�
	pAY-3��Z�̼i,!�$���%�mۻi��H%�^	h!!��"�d�����@�HEB�h�%_!���&(�X
"E c�F��$��/!��	u��P����n���@?9!�d�?%<��'B��G@��P��^!�DǇM�Ѓ##W:j���`
�!��:qz�k ��0��=x4�ހ"�!�D]��P��E�$��T1d&�yv!��8vv�(5����v� ,�%�!�d�+8�t+!����>�AII�{u!�ʓBZ��ƩA4A���n!�a�9�Sk��11���p螻,�!�$[0n�ъ"�y��!CH��!��KL���I#��b�&�5r�!�dJ$K�j��
M�k�iYk�:�!�� Lء�fl�H�z� חW�:�"O�ȫ���#�X���,���ӑ*OB��w�� |��ܸ�&ϓ:Z�!�'�J�1G�W�w��e�	�3:x�	�'��v��.C%��c��W^؀	�'a$	x�F��y�f};6/ϊ'��S�'�=��8.��.���2X�'��y�"���l�0��y��0p�'�H�
K80��S��>[4�}k�'zz@�  ���   �  �  k  �  �+  �7  �B  �J  �U  l_  �e  l  cr  �x  �~  *�  l�  ��  �  2�  x�  ��  ��  =�  ��  ��  R�  /�  z�  ��  o�  ��  g�  f�  � v � � �  Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�� |d��"O
`�(�;���8���-0��1%"Oj4��ND^[��"3/9�0|H�"OB���H��*�ʞRy=a"O�味V�!X��!&F�:J�$���"O,��a
���C�Ą�M�"O,$3%o�-���p���+Ն�:1"O��ݢ1����`���y14]2��i�<�6��{_���c�H�`�fX�$Kn�<��A̼VI�xR[�)�Ć�pඤ�ȓA5��('nߡ4�� �)˩%� ���,��r�؊b#`T�eT09���ȓ!�b��g��}�8�F��-? �ȓ
K|m�ș�VṔ���2�%�ȓ"R�X�j�4JN�1�˘X�i����̹	_�jZ��1!g��zܶ��ȓgil,*�J�
j�Ne��i�J%b���f	�(U��:���G��$Y^م�~r�� S�%T"���k\�jx�ȓ|4�1�îJb��@ӵ�ݩn�V��/[`�"�v4�R�!ʎ<��M�ȓ`:��z�ؚh�J�Z��$HY:	��H��p�m�C1��!��B:��0��EnjZA V;9����J[
2���	��4'J�EA�IVW&��~�(aZ��ӹ�>� o�Y�|�ȓ�f�A�
Ο7�H��M�$�����mޠP����/���ANXo*�ȓTv�����{ ��-7�*h��I��sB�8�8���3����ȓNe*M�悡;������X�o��!�ȓ'lj�#F�m�+R&;�|��2)n�C��0S4���T:
b���:�0!��e֊��)��ͷV��,�ȓ0�&�8#���� ع�L�����;�P�AFd���,w�6d��r�EQ�( �gVlɦ�M,H��,DP���|�I	$G#\���ȓ"�)���E�B	yt&B�^�LɅ�4�� ��eëF�ڙ��n��R�p�ȓp`@}bŇ�=�$�AUN��P����L��p���_�a�)�Y�!��-��u�5���o}�`iF�@A�p ��F�\�0��[���IF/5���k>bTؖ�;K'DT`�^��@��fnV���Y�b�lI��	����ȓ,nٛ��Ć3���kC��8�m�ȓ'� I ���x<=���޳{��	Fy2M3�S�d��(&�dY��N#}��Ձń�%�y�޵odx�H�v�����,@��yB��+�P(J�h=qbJ�R/ʃ�y��R+xd�
'�r�(�w���yA3�����9^)z,c����y����
I-��n��Su�q�
Ɉ�y�ʋ�G�m���GZb��C�ў"~ΓB�����C����%o!D��ȓL0q�w��)@R=8�瘆�t��}C�)vCA�j�X�c2i3hi�ȓ X��T��<us�Ӊ:�E�ȓ<T��0�U�l�j�W�
���Fy��$$��5;��R( �E��C��O�I�!��ðw���)f �9(��H1cѵ�I���Ex��� �r��x*l��
�`�`\�E"OD�EY�?���3�oH�D��eB��X�d4쓩4vԩRES�l����,1�OZd9�4"m̅�g��`S� J ��)ζQ��S�I��4|H����`�\��:>Bq�&�+w}6e��$�'�����)�|<�ѡߤbY 4��O�'F~T0�ȓ/	��[���7e��#��')����ȓب��ҏ�m�(�oA�}E ͇ȓ~����7+����ER a�j�ȓ�$�"k^�0�*�H��ܠa��ȓY�� w��QA�8�$ֲJ}.q��I��aPEg�L��AK�G�p���*�b�qR,ޤl�BH�ak��7]j8�ȓs@Q�e��o$�`��]7� )��Dz��"�ʵӅ�6F�M
�X~�'��i�0ˆqټ��q	
W@D�
��?�ӡ��@u�U��N�; �xE�VIĭ
%!�d1Dh\h����j�f܇�DF�d���/�$X�����i�R#�'�y�k�U�QJA���"�Rw��y��i��"~bED�i��y�P�ԃH�$}�KW{�<2�C�a�T��a
Q�C��� s"�������<���'Y¡�!aW������B"%S�'��i�E~F�H�g�^�O����ڴ�PxrL���*��˭w���G����=��{M�;XpNdIWp�r(t�Z��y2���p\�0��߰M0.O����~���Ou&�qG��!XD�0ě�?f�;(OB�=E���<0Z$��� �h�|�-[���'�ўb>�{�L*�2lʅ��S-����:�=���I�|$��9e+9OR�k��>m�C�	,@E.Q� ���o ��C$��.��d,}R�_�y�f�&�>	���"�/�y�����O�^QD�eLݝ�HO�����TZX}�fn�2�X����6���hOQ>�K�U+"��tH#i�2�,4�E�w�x0�?���O��j�>���Bb�Mc�X��9�O6Ov�Y��Y�u�ba���Z�y�!�'���hO�Oa|M" �Z�2H
r.]�$��X�Ǔ�HO�Lh�ǈ:6���LP0F��"�|��)�S,)CP}�bO:,6���*92 p��hO>Y��Ŝ�$�L9d�[�^��U��OHlEz����B&��R"�׍ ��&EXo� �'�ɧ���I�������\�i���4\2Yq��d~Ӛ��7DYh��u�NL1%N"1P� ��Ű=�{2��O��6�ɶ��
�e�<z�!�D��f;xI!���	ҥ�9qe�IA?q	�c~��V��3���C����6��$�O��=ͧ�ē0Za.?DA�L�qm�3n=�amZr�����vխV����p̘�F�j��V"�y��TϢE�#�]�D�H��]!�y��Z]���2��!�*�ˠ�=��=E��w<�ă8(�fU�mҁn^d��{�'Ml���0.��ȣ���@P
�'����� �:8��hO��©O��=�O�'o L��a���8"ݜX�b]��'�l`+�IbBh QsJOa`��M>q�{B�OPb� +�_�i��b�i_�(�9Į5D���U�J�=� ��'@�+Y�P��>��'�fb��'��pk��Iq�A(N�b`� $�������(���aJ��.i3�┨;P�mx}��0�FBt�*7�� i��jV暧W]~9�Ɠ8c�d:�����=�R�fB�OU�C�)� @B1�Aq� �1r�W�D���'�ў"~���\�
q�f��r�"@���y���zB��E�dt�\ZCG�.�~B�'���"��6�p踕LS2�I��'�u�S�!<5���%,��'�B���',N�q�Ȏ"l���&Y�	�'}�Q#QDމ#��r1�ֈzAʈ�'y�!!0��X�$TQ�O�
 �PJ�2�)��Ax����*�6�*���Iʊ�yB��g�H��� ����m���'�����ð�H�)�H�.1�i��(� 
�!�d��]���4�F�w�Ȩ�5�N ��b�ԅ�	��h;�d�v!��!�'�+}1��Xy��)�C�)hN�k�BH�^����?�y��B��yJ�,B�,��ȹ�B�1�r�����me�"��x9��(�A !��W%qZZئU�G�@\c�n9�ў���	���lze/B
jb�!��L|�#>��)^�v��	�6�es�d9eK-qH���z��ؠ�A#j�`������"BMI�;D��#��p#�)����) H��X��7D��� &G33�"m����=����c+D����gM�S=���n�*�%�&-+D�P��M��5�3��q���y�-*D�`��͵uE�V	��4D�U��5D�j�FZ16L�R�	,���h�5D� jtQ�hi�ٛ��X�1W��k��>D�ܪ�)�e�P�Sh���4b�b(D�\�&��s:
Q��sO�th0	&D��(r+�
��h���,��0ڄ�!D���t��!i%>�"���3�Vl�/?D��x�	@]�P�fB�2���i)D��J�B��f:�����,���C�"D����� E�z����^'���-&D����D�'�81�t�u��y.1!�����R���&�I�.	�Y�!�D��F��M^1af0�p���N�!��-X���Θ�C�h�!e*O�q!�Fxv�vE��I��̈�G�ga!�d�	h�v�zר�r���t,!���+��si��p}|I�ιT�!�d��9|5���Vub����Q�"�!��0�h�U��T���3�,B 	e!�D�O3l`@��ܒF���Ⅻה(d!��9c<
upUM\�dB��ɂ�!�d^#�8�٧號�Rl����#o!�_��h�i�
M�`��FL��lr!�$K3�F,�"eN*�
� LJZq!�$�3S$��·p������GV!��� LG�U A�
A�F�S���8L!�������4NЊ����CtO!��00���de�6S���{&d�;�!��,
�بaW�M�d#����,n!�d#\��F!�#@�	�"�-RR!��ƩmM4a$��(Z����d;!��BZ��x;�n�#A�cA�4/!�d�44"~iSЁգ�.�*�O\�P!���,^�2�I����kь�%3c!�$��T%���O�r�t�2l��K!�d�&\�2�k���r�̘�P@�s�!�Dͅ{�vy��i�:<��}�#)J�0!�ׅO,0��Ů�)i<�kghB>
!��؇V�Ѐs�*��V�4yp�=8�!�|2�}(�)Ѱ �T��� ��!�� �la-��D��b�C�}�H���"O�I����Lx8m
s�)k��Ő3"O��1�@Ң
A&<F@�4��"O�%p'B
	F��Їd�s)���c"O6M���86�܄�s@Ö��8á�'X��'��'�B�'�r�'��'f@�(���L��U��&?M�$���'#2�'a��'�R�')r�'V��')谡��
� ;&"נ"KP����'�"�'+��'���'���'7r�'��=J��Q=�0�F�3����'���'b�'{"�'�B�'���'ޘm�-��`� �9A��7n���P�'���'"B�'b�'�r�'B��'�fi'HȦ*0 ��1	4���'���'U"�'hB�'X��'_�'�!8c-� 1��Q5-H�}2��'���'�2�'���'v��',��'� U ট! i��b/vQ� ���'qB�'�B�'B�'�'["���߱H�Z*�$Q�E�DD�	��2v��'��'��'��'<B�'|�ā �� s��|4�q�'b��'B��'���'���'"��'�ĸ���i�� �x�Ai^kE�}�I���IΟ�	��0�	ϟ��	ҟT��!srF�B��G�d��� ��5�\�������ʟH������쟜�I����I�^�$RQ���'T��0��f���	�����ҟ�������	ٟ8��4�?	�*�i�56�f��L�
t�0t���Jy��'*�)�3?�p�i[�h�m;<y���SnǺ/�pb��N���[Ǧ���Z�i>��ݦ]�㉖�RvF�XG�����=�.�m����gEϦ��'����U&�-	����\���eQ���L:�;HE��R���O��h�ƨ�D)��LP�%3�A�TIbj4�
���*��?!%?%
�����+�1)!�r�Ӂ*� ݠ'/����iG�D�<%?5��$ ���E��e���_HV��nŢ'���͓A��LS�U<�0,r��4���>,�m0��50utg94_��<�L>�U�i��1��y���;�,�*�M�n� ����z�b�|"e�<����M�'�������UFT8a�~��Dʋ�!��}���ҕ'Ñ_GB�|z�烄�uG��O$���1F��D�
َ1R�a�7a�<�+O���s�$93�S�m���%ӴT�T�b�`�,��4�tt�'q�6M�Ob�O�Iy�"�c�aSu!Vժ�/J+����O�6��Ov��|�$�R�
�#��,ox�!"��љBU�M��m���0y�����䓌���D�4����=�@�k�J
�`���+�M�@�J(����O6�?qR�'�k|MH����I�N��FO)��d��Y�ܴ���|��'�?�1nT�DN4l���>[�vHBb��_�����D���$��uĤ�+�c��N>�.O�mj�,S�x�*<�ehX^bZ�)��'�.6�S^к��"m�$eSS�85q�VM�s�2ON�oQ��O��	��Mce�iZ��	�v��Jg	8~X�Ц`�!	�"M�6�is��O�� �n!��λ<)����c�\=0�<�1m���Ժe��<	��,�Ӵ �!��q*v�ʝx&\��(O:�$^�3q=B��i��'&$=��L�>��)��#�|F�|�(r���nǟ4��%C�}̓�?�!iIj>\��mΈvj��.�[\��u���Hߞ�8����<)��?����?�3ŝe+`PI��]�3���\#�?A���������������ϟ�O;Z�:�D��j򑂐��`����Ot|�'��6m�%����?���A�h�*AQ�.�2���
��]'t�yG�Z0G����A��ugo7��ϛ9-Ȉ����V�IRpI��mQ����O���O��4�u�G��O��$A��f�'#BT�B�X$|ʜ�rퟶ&`bT���޴�?y(O,�$�s}�(b�r��c���/5@�3Co]%ZM��������ɾW�Qo��<���*����M�w�5�-O���9
���K���4aH �hP=Orʓ��=aVfҖD��Is�����XgL�}K���>l��'���i����L˔hkV��-��Y�1�Ŷx$����4̛Ɨ|�O���'��;B�i}��(v�,P�P�	:D0��3a��99x�� 5"�N@ʗ��6nV@:����N���J�	�vp1�#��	���U�;)��E�g6\x���N	���U؊��C�v��s 	�ov�pak��M�J�ء(�"=�p�'�&8;)� @R�Lr1}� }#)OnM�I�	cO��D������ґ5�l��6Ŝ-G�8��n<���>s\0���F)8�z�� `̴v��QR��T|ac`(	&5t�
�� O$�,�E@3���2�eG!U� @D�S�RNĀ`��%�e���!J��Y�CB9慳��8f���S�b"��'�B�%P`��($98��O
v��7-�O �O��O�X �OT�',t4�FeEF��s�U/b��|�ߴ�?���?���-p��p��?m�i���O-�Ab"�Q�}��a�ū�)|���t�>��O���P�Tr��:�Ba�/��G���s턁8o蟬�ɉ��I�	̟���۟L�SLyZc��PI�4�e(��D�*QN$�0Ot���O�Q�)�SZhI�C/E�K�)B!��9 �1��4K�$�h��?���?�'����O��d\9�X�[Q�	:2�0(�
��%l��7�-�?�|���?��7Ua���v�I�<�^�CQO���'���'��P�P�d�	ޟt�IH?!���i&F�z�M��8�����S|�&k��L>���?1��v� Y� �%Q��!s�D-qh��ia�ib�c-�	ʟP����4$���!X�0T��;M\|X�e��C��˓��e%�D�Iϟx��YyRE�cB��[Dн	(v�WEKB�YIV���Iԟ<�IP�	ԟ8�I%�A�E�8G�r%q���&���1�l[��Ԗ'o��'�B[��Pf�XR���w������ Bc�X;'F��a��֟��T��֟�I5t��������R'e�:KX�bM�-Vz��O����Oz���<��(��)�Ov���!�� i�P C��pS|$�����	Z�I���	�AI���IZ�dI
:�ę��L�kEth�C)��f�'9b]��Q���]�$�'s��OT@u@3���U7������Z���c�:�$�O&��]�>I��'L��)EӜM�L����z��o�Ty���yr�'V��'��dS���Ʃ�"f� �*q���	�k�86��O���φ?ɴ�b?��	����lb8�1����I� ��MS���?9��r�x��5f�,f��A��2
 !���زٴ1�x�a���?���?��'��9O��d�+p�BwJ� �KP�I�_r�n䟬�	�(���@���|R��~��P�k�j��#�>�j�ا#���M�����/*� ����d�O`�ɫP���B�'/>
A;�V<X*6�O�0��<iPQ?��?	T�V)����j��@a��H(|��ɸQ�Ƭp��5����l�'�b�./����DW�נ81��І=C�u��[�4�I��?a���?����/-ߌ���=j��v�
�h�Ȭ*"w̓�?�,O��d5X �S5���ZĈ׬_k@ Pǡ̢�P7��O6�D%��柬��Ѧ��"�r��E����IҴ�a��\\���ŒxR�'���֟�Q�h�O�$�'P�1�
��A�"�JsB*H����c�a����I���c���W�O���M$�����L�ZaB�i6W���	�Q����O�2�'��\c��HZ'$D�'(�P����9�Z��H<���?����6zy�<�O} lveäz���� =O8}��4��$�.vg�lZ7����O��)�K~b���T[~u�D@�2 �~�rQ,���M[��?��]��?-��'�-���c¹s��Ȓ�G "Xv�R��M@L3Q�V�'���'���H*�4�k�ڱ S����'���BE�V��=�R�'���'��]>	�O3�x@�|�u���B�@;~�7��O����O0�B`�<�O��_�ލ�tϜ�F�;����=k����$R�`$$>1�I�����qJQ�+��5�*��ToY5�D�4�?1�(�l����t�'��W�Q'"؏enT��6oO�tsv�3@��M����> 	�����O ���O�˓},&����/���w�
N��8��^E��'b�'�RP�@��ٟ��MF�LX`8`�� }e��C;w�����HyB�'�rW��	�O�(��'^~�ȕ��PT(�C�fl��nZҟ���Z���?Q��r �<��dHঝh)�\��Ӿ�(y��h�I���ן@�'�bS`&�R -��X�
T}��[+�H���oZȟ���vy��' ��.2�~��*�� Z!�>���5�Q�a�Iȟ�'KT��!5���O����rY��ub$�c�(*�Vu�g�i2��ܟT��6f?�|�ID�t�'��\c��P�GӅ{�>P�2. �*�"ش�?���<�f�i���'��O)�$�'k����G�t���P��&r���� �>����J��?)O�)5�TaN�L#��A�@�)�t��a)�9�M�ׁX9%6���'#��'��$�O-b�'�"*�7|slh���-���iV$�Fq�7m�����O��$Ev���'t�	ҟ��сQ�\h��ѡ�_� �l���M���?Q��bZT��i���'cB�'�Zw�J�aq��P��l���;bȰݴ�?�(O�<�&2O��؟�	���a��A�
X����u�H3L��MK����L2��i��'���'���'�~�-Ķ� #�p�܋ ə0���S�	���O����O���O��'BR� �J_�mr`\��Q'L	D�X@��	����'o�'j�µ~�,O��+P/r��H;P�r4���hH��E6O���?����?)��?��Ff���#�*4�H����ll�S !��:5t7��O����O���OB��?�s��|E���^�J�1m�>��f�'I��6�'��'�2�'r�\�d2l7��O6�D�& �ܘz�ڻhp%���7$$�n�ß�I� �'2B4����'��V�z�@W�B�R{f����H_9���'�B�'z2��!8D�7-�OX�D�O���׵nl�Ӑ�G�bn(sq�p��pl���'��	��O�iMb%���}┰%K2gu��4�?)��!2��1�i&2�'���O��t�'vf�2g�R�[�`+%O�	�<�EK�>Y���5���?�����?�$�Ӆh�>d(���p�����⟰�M�s	Is���'���'N���O���'��"��=������	M�X�#��
��6m��C���4�4����f�$\�sX5�F��~JD��%�����l����Iʟ������M���?��?!�Ӻ#�a��>�e�q�҇h[u	d�����cy��	:�yʟZ���O~�D�$`v1˵BE�U���P�81��m��xX¤� �MK��?����?��^?U�RW����HX*;�Xt3���j]���'���K�'p��'�B�'�'�bH�$�<�x ���I��4a$h�DE2�c�&�d�O4�$�O�t�O�	��\)⧂�&�~訠#R�Z�h};R�����	ϟ��������ȟ���˟,
 d��M{�� d���kV����05+�c+(�p��ikB�'�b�'�BY����o8�s�T�+��_<�@��IՈo-
��i�2�'s"�'�2�'/Ҏ�[��i�r�'��E�
�6
ް�Tk\�?���tӂ�D�Oh�$�<�,����-O��I�f��5xf�N: Z]s��8�F7��O|�$�<��jа7��Ox��O���p�R�Zl���R�<,�\H� 3���OZ��K�VҜ�D4�T?q�0h�
}�� �G�CW/8X�Ho�˓N�b��i����?��':�I���TB���<������T)~M�6-�O��DG4���)�4�4���Ok,�$�2@yQO��)ېXswƏ���VB�?/��7�O����O��)E}�ǟ�p'ф��<���1n�8`u�F��M����?I>E�D�'=��`E�r�$�玬@^�tBv�^�d�O��$�(1���&���	Ɵ<���2��ć�F�8�#Y4Zhn\�I9~��L|2���?��;���V���j��?F���YEH��k7�'ւYJs�1�$�On��"�����r�X5v����
�P��t4Z�X@�N'��ڟt��럀�'b�M+Ѡ�vZ
�0���
gv9;V�L��<O����OʓO����O6���O?tH�ABM��h�:2
X�@R���<����?a�����P�P��'D�P�;4&�rr�S��$f�Ld�',��'��'-��'���Ҟ')��ʐ�HU�����W$^8١��>����?���$Y�L��&>����Z�U��AD��=c	��B ?�M#����?)��.��ϓ��I�||���_-=ڃS,	��6��O����<p�׽x=�O[��O	|�9uŊ>L�qˁm��1��BuE-�$�O�� �#��������稌$4��%��ۧ�4�o�~yr'1(87��z�d�'����3?iRj�=�b��d�ŭB8r�*�Ѧ)�	쟸rG e��&�b?�3ᔋ!4�}�s�NDH�w�f���Cք����Iџ��	�?Q N<1��
�p|IWaB�+B%N�7[y@����i�&	r�'�ɧ� ��X#_����2X󆕐b��,B�o�ǟ��I�p��C����?1���~�C�(+�J��ͪr�5�����M�H>��ą�q�O���'��!
$v�x��Gɞs�<��Ūf� 6��O ����B�I����	A�i��AaH�"�BԸ��4u=�%�� �>aa�_�?�)O�d�O��d�<�����` �y���1����tHԔu�&�ȁ�x�'���|�'�2阤?b��LF"شQIU��w�
�'��	蟜��Ο0�'�F�K�)|>��d��"Ү0�1 �
�H��զ�>���hO��Dڄ����ψZ���5+�5D���� ��t=�'Y��' ��'�B�O#%�z7�Of��^=0��i���G*z��a��6��m����	ϟ��'��������>�KB�R��񃑌B#&)J ��,Φ�����T�	ɟ0�Ŗ>�M���?a���$��@*�$��W�`=�W+�T���'����� �o>a��ky��M�憖�vϖ�����X�R�'�צ���ҟ$���8�MS��?	�������?Y"���i��!爒C"(�I�7.Z�I񟄩���t�Ity�O��'c~|Aa7,��S=�X��+;��l6j�Q�4�?���?!�'����?q��BPf0h���_�(XDB�<��#f�i�Q(��'��W��o����Y�㈬_��  b-+c~������MC���?9�B_N�S��i���'�R�'zZw3r��'%ܕPVm	�`H�#���ٴ�?����?ٴ���<�Ob��'��B1n�XB%bU�=.��Jr��'nO�6-�O,�3R���Y�I����ݟc����ɌR>��kb�̰ЩBs��^j6��O 5b�4O\��?1��?y��?e��=@�= b�]������s�X04�i��'{b�'���'����O� ق
��d��PK�-'�Aj��Ʊ��D�O����O&���O��'
j"y#޴8�x��3 ��UB<j �0K�Ms���?a��?I�����O���2:������Y�2a�G>*�]h' �ͦ�	�0�	��d����y2RG�����I�0�v��	�ʩ����.n�n%�l���Ms��?������OxA1"0�������j�J�5.�N��ُ`ȣ@�u����O����O��02�H֦%��џ���?��2��'�*=�Q�T�Y-�4�p�ȁ�M�����O�=�w0�����<���Ã-�D�H�c�
7Vy��cӲ���O��ˤ��O����<���������D�&,�Nq˓�B�UyjQA�iU��'5DBŐ�՘��O��J���^ͨ��f��]��4����i�"�'�"�OzO�IP*3�%!#����a�D��(���i$�E��4�1O~��X�mT�5iS�;wE։��mE�C%xEm�៤�I���kf�ky�R>Y��o?q��ӣM2>�bs��bl8��Ȱ8�1Op:PO�џ��I��pz��׀^�ةx�'�"�z(���;����O�2˓����O�O���C'+ziSp�� >�h���KW}�jѦH�j�O@���O2���<Yŉ�1�
`B�3o��xS�%8A��'�x��'�'��O*\c���L���@E�6�Hr�l/J1O��$�O����Of�>d�����N�8�ī\B���W����l�ޟ��	��'���I�LR���fb�7��1d���TAC#i���eX)u.�I:6g⡪F�߭��q��5�')���+�F��#;v����J�@��ȓS����w��#,Y&�;Q���'����2�m�b)�v��PX���rG�� ӓ ��������6)� d$r�KX$X�L�0g�d�8("�E']����FM��;^M���F�ĳVLW:d��[�a�P��q��N1q�0i���=����nU�!��q�CK
�\�q��2��5�(���� �٦-��lC�	�OV�$�O4 �cI�)r����h�<M�y��L��	��H#�-�� �LH�!��M#�瞓g��!�|����N��C�M3s7=�Lj����2�X��4��*H���`�˶ ��a�pl!����Eό�qe� �^<Ee<C�	.Y�����m�ߴ�?Y���'EB�Y"�U���`�4���'=��'���3'и^�݁"�@ dj�yb�'��#=�`U�?��/E%=����d�ޫR���% ��?���%�C�Ç��?���?��R��.�O(����G�j��$fL
N�*E@@9U��9��x.ɗ�Z�v &C�ٟў�j"-��{��H�L���1�C�Y��?���9X�4{#\�,vB�3���X�����А�Ba���l�p�u)��@�vmt��Y�T��zy�+��U��e��iqX��$O�5�yR�R5	 �B��O;b�`5��<z�"=!���?A(O��G�Ŧr�I�8�|嚦�O�x݈=�!�䟐������ɂ�X�	��ΧP�`����;$��y�Cn.2��*�@B�~1�a�?	��E��'t&-+ņ�HtJY�@�fZ���4�n��5�;��A(��?,O>�"�'Dr���r2���MZ�G����T�1�ў�G�)����=@��u�c	�"-�te0�'����
�2X���'��1+"p �'S.듴�d§%�"XlZ��D�I@��ʜ�Q��I�l�~U���V�.5��1u�'�"�'��a�� `6�� RD�Z�~���Q>mi4�	�aC�1W�ˎ2����A*�nux�h��6XC Df�զ�Ѵ�M�-�j9Y�n�7����6�R���@��e���q������sK����O�r���3B܀@+��g? ���:�B�|2󧈟���Rʞ�C��\�z�ീ�%[a|bOzӠ���O�@d�/J&8BKq<X�3O8��$��m�IٟH�O�p9�u�'$�'�@��mR�f:m�$g�?x\� aj�X���A^
���|:��� V�@�7�U+]�n@*#ڐ+~�R ��@'�k��}���Oz�"��X�3<�P�bhY(d�^�;4���j���Of���Ov#~�	!@h�2Dl�[���K�&�d+����܄��m���*'ď#�`�B&ӝJpT"<A��I�?Y�ɷh��юE-I#�1��4~�����ޟh��K�:b@�e�	蟜����9[w���'n�q�LV:a0����֯O\bM�1��.��
`��JP�}ʖ�ۿ����G�w�Ԥ�V�G��J���HƧ<*�@�O��Y��{1O�OɎ̫�Пў�ѳF��<�L�xd,ܴ	�������	f
�O���(���O���<	p��q�����b������^�<�DNDA�|�P�*� r><���S�4������H�'6�q�|�X-�tK�
��X�g,�#z�1�!�O���O�d+Z���OJ�S�X�cX;[����T
�+DsXq�*��|i�-["�A���8#��'�4mt� 0��P�ϊ|�ЪF��0�ش �o�:6,p%L�j����.×�O�i��'�,6�D??(D�����>��+�d��b@�oI�[��>��p� ��Ϡj
*�â,��y���D'��d\����5�x�cs��Z��n⛦�'7�	�P<Lx�ߴ�?����)�rz(�J%�7�}��DM��S��OR���Ot(���O�r����H�4�|�^W�<�yw'�;D"��C©ܘ;�Q�İ�T��|�0T��sNV�����'�	fI��a�=m��8�剁����O�����dCF�I���,n�`t�[�~�0��;�)��<)LI%�E��Z	@�}��T���J<�I�U�ZذqC/gߔ8;u
^�<ū�6����(�O���%�'���'�����',>ޖ5�u,X%��ri�!X	ZAz��ԟobq˶��+�l ���Ͽ3�O� �>=��.^,X�
ܱ�S��ԑ��7b�U��*�fXQy6�.���UJI��Lo(��ש�q��<bC�D%�$��I��x�I�LF����U��
dZ@"ƾy�¤(�'��'S�� ��~P��9�l��X�1����t�'�$�'��Ɓ�gYգqa��c��t��''�HO�=���f�'e��'�RA�~B�� X>ӏ޳^�Bc�nP4h��l�|are��%3hl��������DK� �f+�E)DaN	c�n�pj��jK�4>|�
4A�-�d{w�g>J�$
�s�	csJ�-@�$m�(yӀS�hm��a�#�gк��1��$�ݦ-�t�':�^�� 7��.w���6�#� ���"D��A�@̼.!Lt SjW�.=*�He� �HO��'���@�+.��l4p��h2�9_L���hO�]D
t�	������ڢ@����I�|R�.���@�2���(o��rv�D;��x���úpč���D�T7���d�?$�<iqD �Ft�1��Î/�<iAM	"��<;"�1k�n\��
�Mk'�U4��;����'3��3��?����.C�cf\�p�L���ϔ�?a��s�|��B��(��@%K�I�%(D�� L�#��L���XԎ_�	��I�r3O.o�p�'2�8�fɻ>������%.�1��+�_�\(zrOZ(.�H*�b�O����O��d��rx
�*��[f�@�o��{Rc��"���'�ޭj��sT皮x�"��DH&�8}�US�<j>:�v�:�Z�0�[1`��Ji]x�Ï�n)j�ˁ��N�'�x�X���?����?�)���0g�H8+ڂU���9G��u9���O��"~Γ*�P�`�B��x���3��j~`�'�ў�S.�ēj��H�vLY�	3L4�q'E8��eb �i>�'��S�i����I����	� F���CF�'<�� ��E�=8ВP���	����C�"���Cm����'�	��o�Mxny�U�	|"йJGZ�.�u!�?�(]�$�+Ĩ�|�ٓHUdd��S�@����g�'}V7�}yJ~�����DΝ+�����D5����	'CQ!��R9&�	C6��('Cl� E��-�tJ��D��Y�ɸ�����&��G���D2�*|�Iϟ�k��Y�� �	�0�����\w���'�d�C/�1%!�E ������qA�lZ�p���&`1����I�+D�	A�yr�26���sv�.(����]�Ln�bC̞�j���B)æc���O�8�voN�G�(�C�ψ N�*D
�̪N@���D��I$�Mk�x��'�RR��a�;g���ҤTt�M3q�/����T0�ÕO�FR����؆�$�������:�4�p5
�$$79Y3d�r�$���"O��(�&�*-���Q�Y6(�6"O�x�'΂#2
��e֜L��J�"O����N��6���B�U�w"ONa�S 2-��	�f�]�_v�Eht"O�H��ē^���eۤC^F�qG"O&Tzת)�"�c�e��b�ias"O
yۗ��<GlKց�8O���0f"OBH��ƑE�
X�jܥx��=Z5"OĀI�7m��} �*\0���"OD0h�G߄�6�jq��>���x�"O���2�ҞR��(��J�e�x�K�"O�uq"ψ)y�$��E+��9��"O�� �НkP���4�VV�ł�"O"�ei{�'(�R�Q��.8䤇�2[68R�-��(q� �Py�ȓ"]8-"�E!

e۱I�jeRX��p>P1�cǿTt!;⊒@� E��+|�ү�'�.�cB��qP���3�n �&�
Q�*����WW,��J,�ș���
�l�c��p �\����aR�a�E���N ��ȓ)���#�/|F��jԍ:r=���ȓ?�@}�U'ʜ!�`Mr�*�4~� ��ȓO6��Z%Z��YF_���ȓ L��ڳ�3k`M��l�p
 ����BH��C�=rh��&
lΤ����Ǯ7�Ȍ��Ǒ
7I�؇ȓ.t<�D��V�4�q��[�E-d��WB(�5�39�X!s7�N8̇�o�(A�)B�:��� v�p��@���E���P\�7
�=T�4��ȓ~��T��� V��a��ؿ8����ȓ>$�(�;5j�XR#��k{2ل�q�T5WgJ.Q�F�:�K��$F<�ȓsL6P��$Ս�R$��1p��ȅ�4C(���f۸G�b`rEF�7W|��Uq�)���N�}nP�J�/QQ���8��i�V�C���A���+V�"����i"�͓b=>�`Մ�,jGP�7lG*U��x�ȓi7�Xgc�8r
^M��]8T��Fz��Ŕ[��E�$C5Iu$p�&'�&�8�(�OJ��y��R�j-���ઉ
����^��M�Q�U�5�\4S�x���i�x��p/�3<�Dr��ۙ-����'3v-+5,�;N�֠O�7�(I�O��t�ЖF����ϓgh�6��*��2�U��\%D��ːg��	�^�2�H��� �� ~�8�"����� j˵8v�u�JH<Y7^�1��$���$�%[PdT{}��Q�l$��m�L��o\	CO8��~ڢ��o1�Aƈ�3\��W�@�<Y$��� =k�ʙ�D������YӦ%ڶK�'�HH�8^p��?9Q�@-��4K�2���eŒ�;�5HabY�)�K�h�dܮ�5��,2.��CA�_?�r-��q�f�3�\\X�� �W3VL���
��x!?�T8��`��xy��<<�Ѐ�QOţ:%JIpׂݍ �6��Ԡ�/m�DB�7=�*�"PR��i�R>q�>� ��(�F�����E��
|��B��5�Ӏ&�ȅ`'f��	϶!�V�Q$v;C䉥RwziX��V�f|�h����n�Y(q���E�n��a�������/���ؐ���bH����2faB��a�%��mx�z6�&1�u�H"iZ��"����!��	;��,5EN%Cۼ���Sl�V�>�G���U0��˸m�<�R`�uG�ϫkAP���BJ�V�Z%	cB��yRc��-�R��)MF���>�y� ��ub�(�)1����PkЛ�?E���ҟ?��J�̏�Vu"���8�y��%hR�%�w�W@�����,]��\�"I��?��D�Z�l���g~b�|�ōN�sbَ(x��eʘ6u9a~bD��\�n�Z$�߼ I�4�b��oN��d 	���	��?}��8}Ҭ���P:՟~BsGos�$�dB��$=�2Ji�'��Ɂ�e^�$Li��ʎ��FH"�8�b5�`���v���I#Ü�S#ޥ��>�N�	QgƽHE���}R#�IV ,� S�n�`��N�ybҒ;�0D�R��/v����W+ ��?%?7�^S�@��ë69`��#M��r;<���j�0��䊨w	��؅ �3�BŢ	̇ X��x�(ݯ�B`87"Dj�}
���^$K�o�0XN�O��,������6��<)��*�C䉀V��(��JГUŜة���8K��	j�G�i�����Zό��OP(:2�����lx0�S3�9R��	϶!�鉉YԆ�AÎ�cӀ�hشYH�Cc,�)a�|��D'	�|)�)yO��31�V 01��PL|ΓDhr���'j`��ʇ�g����-(�J��y���hBJ�S!�Rf�	�8Up�c�Aݷl�r�� I�~�\�0�QrUD|Ȉ{B� �n*Q������'\R��W�euD��,\�)ʘY���[n;p�XRO�
7A!/p4yj@i�z�ꈯ;&a�Ό��p��F��A��5��-��iu%?��@h	�3Nq٦�,��?iq���7ᠰ���85�F�Y��!g�
�8l.��k�e�>q`�'a���ź���[�f��o��ͻkz��x���K�R�Y%��/�ܽ��OZ�g��O�S�y��h�Bګs�Ƹy��T��u�t���x�F�zq��]�^P�G7�?��b��wGL�����t���X�Ƹ{�4r���$8�V,q�_�@ݜQ�O*"�>�J9O����1ul� ��ӊTV-s�����?�֤��n�)L��p�T-4`:ar��,]>:� �+_��C�:����@>rq�LT�:`�'_�j�	�#L��@�ǴK�T��D�?��8Ƭ�0Ox�O��9Ĩ� k\�m��M� )m��'rV��I1K��A��H��>�����-p����$l
���G�2־��'C�b)�m3�b�����yj1��'�f1b-��	���%��0|�B������#���B�V�{�ldLY�b(�|5OR=yr����y�Ɲ�l��	�SBH�VO0Ez@ω!U/\�u�=��	-������GFԼsc"�gYja��*���n�0���=`|�	�}/�	yE�*S<�����'�j���ԃLur-㡬D�T��8�"_�Q
��+�">����=ɑg?�z��'�!Vyz��V WG?��jƴ!d�.�3��y��V�l.fM�JF]�y���S�8:L��6ᒮR�6	P�p��U4d΁J��'i*h��+G�XDaD��t�6�{*��
����C�� fDs��� A�>?�����"|r��{�`���i�!Oo|mH$ƀ%w�`�6�|J�� ��ؔ@�!�y��Sh��a@g6|��Q���'���)p�ɿB�8i����(D��v��=\�M��d� ;��̓(7j���Ʉ9�F	��CA�h�D�E|��R>E���D�;s<��� [��hO6<��G��Gy2P���&�1�R�O Y���;�6 !@N��SOhx"f�%nX谑e�'�p��T�D7�8�;f얃 ��\b���Ju�u�Þ#Fn8
F �vSp��=�O�܄�7��3P�EZ��0>x���"O�b�.W�,��
���[^݂S�� mr�Ɏ{*��9b872���j��JL<
s������LF
=Z��-�O
<X�p(đ�҃��Y ����[�x3�y�h�!@	̜0���Ϋw����֋+�/Ґ��p���!�-Cwg�E{b�dj �B��Ĉd����9�~�ĩ>X]bL�O�6�#�c �#~J���ŕ�0?��&1� ]���$bS\9Ȁ����h'�x.I 2ͅ�Lh�����*�|�$�6z:��A��;�М ���yR�ԛ/�E���H�V�)��ʸJ���*Od�S���Q	
�2WN�1��d��lc��g�V�(
���%n�9
��}"f�J$��2� "�r���1����)~�d�2O~��'�o�� �O^�a�"�v���y�M�uxtd��������CC���M	�����=[�S�OW�\���'Zz����<�����\����Y�5d�)���ŚX���y�iU�f�B�"�'P��'
���?i D	`R�p �'�1"����aEk�S�Ԭ��~+��TJ��LHJ�DЮr��O�	�QF�OVy�1�$�ɊO�@��0�P�C�\��N�^����T�LC��S�H��]��F�J�1P���2p�Tp�Ի1L�
;Y\�h��D)�Ӻ���E�V���0t�@8;��pt
=$+�B�b�5/1O�4 j�����ht��rS 	�W�"ƞ)S:�b�8 ��z��� �B��6�	v������O���^�,x�[�X(Q�!�,p����Ȫ>�J��Oqd��W��@��h��M��Ri�0KU�i�u ��!z(��'�˲� wX��gk�q�%-�3��Eր���钓����T�K)��pJ�'>U4���t��m[eg��t�b���1SF�!.�XxT�!L�L|�$얚cX�ԫQ.�Ҹ'���*�K	0x`�`�!7��N>��mA�z�>����)�zL�6�
m�[��F#җE��d��f�
Bä��5��l}R�!}���C������u�B�hU��c�Y4�~�K4���y"@�>?� ��m�;m�	Ӡ��&�M���$X��,ze��!�����D�D�'�YqDL�xv����NXb�' n4�`�ƾ&g`��A8�fE��V�MF�����,W��!a�ÌH9�N	�J�y �	۸1�,5q$�R�|%a}�@�nyJ)�U�ӂT�DEJ�U�������g5x�O��� ��'�x,JED�$_P����8DY�¶X��tB��\�&���2u��.��-qFiK�,�:�{p&�>����vKҝ�"HPi0L�F���?i�,�)l�+1\O,A�傇*F���$��!! �$�'�x��e,�?
2��
�,@˩O�L>q��4�"�1@Ş�:e)@%���y҃5r���(�	J6`���_�M�B���\2@���s� �	F�Q?�S"v�؟�E�g��0�UJnH����}�'�x�F�8\PV(�%J73w8x��ᇐX�d�ʲ�=IIͩ�p��'�̫���O~	��FF�l�nБ�{R�Y%@�̠0-_��XM�s�����)(y�l��bZ�#��(��=摞@�2鑘U��ŹP�&'���	�Lğ�[Q�O�K5Lap��'�*4s��̷4:(q!�dn�)£RW��}I��"�JD��Ok��?b}*S��1�j��ɥ �a( �~!��K#>u`�A�L�hj�"�IL�4�I��	#0V�k��3M���I:H���v�їI�%��G�@"��F�����O�M��$Q'~ʄ5�Lz���װi�1BR�݃Ύ�y�D�W�v�:�# ]��a��'!Juy�O ����/'ǱO�8;��7M.VM �h1 X��]�hp�bh��A���.�Is�+ғci���uN	�qV>�yp�JȆ�Xv�O�QZ�풹C_a{b�æSdh��9Jx ��(�9V8m�5M��9�AFzZw��Bd�P4w0�Q�1> d�"��]�D~�I��gÆp� ,�ȓo��`m�Wk������"F��oZ�!�����b�O��Z��'1δY��{>�ÅW��+-�p�c��P������`����$����������@�b��5�$���~B�טG���Ѧ�vx��ہ.|^a�IǒrK��9�4 q����,c4dR&$lv7m�/D%�l##�
(D!���3g��B��=�TDs�b�>C:",�$4��˓U{�,O��CU�V#|"D��$`�P8G�����|�<��M�5i����G"O,���F�y�<��ꏘi<���ܬpv�Qj�t�<���F�J�B��7`��0S(Ii�<i��߰J���@�b��8&"e�<�0�Y��\�^�"�jk�f\h�<9a��s���{� *b��A�a�<ѡ
�*��h���A�'f�H�b�i�<�⮆O�V ��A(��i�% �a�<A��!�|xb��8H�����^�<	'BL)qL�EB�gv�D���]�<�FJޚ.���@���u�ؠYn�<����65|ܨ!�ޕ=�M`#�k�<9�g/�Hi*Lϛ�2��f�i�<��"�)V������ 3ظ�Zr��e�<9��� ���xu��>Fk��AV�<yg�.?�~r��^�^@Ժ&'I\�<9�M�8+~�4�w'�:�v���[�<A�)�USt` �Z/T��
*D�� |�;#!�*�.m��NϺ7�<=�3"O��-�F���'�7���J1"Oʙũ�Nj\�1���4��I�"O���ax�]�v L2Bֈ�3"O&�#ĈF�e{d��3�4�vH��"O|�#@H�� l�p��J0]�Պ�"O�p������M�ܺ�"O>����Dv���Y�!R��#�"O�y��ϙw
�&.�4P�}Kr"Of)��ե]���Cl�@�ҍ�a"OF=#���z�, ���	<n��"O���G�P@��!C�IT��٦"Ò�d�,|��C!�J�sKN��G"O�1iS���,IEz���q�\}:�"O�x��D�w\��Ϙ-��d�0"OY`�mUP���m�&B�@,J�"O�LW�7[T�+󋊍a�d-��"O�@8	_6���;aiرR�ҹ��"O~e;DCK� 5CōU�nRY�a"O(z�(�m�PyO^�8z��U"O6aKg@��m�V�{�F-J�>;&"Op��H���:�R��D�"O^ �� K?j��E U�1wq��Cg"O&�h�j�}�Р慊!U\T�R"O���L� Ag�9ӥ�Z$��7"O�I�Gީv�F\X�#òGE&�)�"ONܳ��A3�(�1���,yR\���"O�u��i|�����$i����"OԺ���Nu��8�(���C�	�?l�1�`£$ ��p%¢b�^C�	/z{Z���(�%f��@��'��C��F4�ĉ��ay���f"/:[�B��%S^ҹH�D�4s��8����B�	�Jp
�2�S=fu$�*p&�=оC�ɖc�z',�%%�*`S��:=�C�	5�pP1���9 �����C�ɺ |��n#v��	�f$&B�C��]��{�`�B���2OW  vTB��t%,�gד,�䴹@��H�DB�&t��H�,}L"ic���I�JC�B����q�)��	O��C�IE*��f��E�"q3�ÉS4�C��-�Z	+�i68@hyVI�$ɌC�I~X��A��}eR���d�<B�I(7<p�1Fۨ$1�,��	Ƭ6�C�	5X��PG�YB9���&V�C�ɣAϲɱ� �N���Yc�D�U=lC�	 -n��i��
Kt���A�NC�	�\�	[�b�=F�%B��*C�ɷg|��FO�gQZ]��B`	\C� �`�9� ];bx\k%��%6�`B�ic$��Ȗ�%��+PV��"O�i��J�h�aIՋ�k"�!��"O"�ʁ��.f�%�� �&|����"O��@Q&͹2�,k0@�&~����"O��x���V�Xh���)N��H�`"O��J��8o���:�.D��2�1A"OR�D*l`	�D�1�Q� "O\�v�Ҿ���+��^.H�hB"O,�%��%9��( �"̍X��;�"O����  B�\�I�B�9In0�"O�-@�5e���D�Q	��a�c"O���	����aܪG�T�"O��pD�4Pnh��T�@�Q��["O� r�:Hӭ7��إ�!)�� �"OtP9�eO�'����g.��fP;�"Of�S�͋�0P�s1LƲ=R��·"O4XK�fQ�6Ĥ1��k�20&�HT"O���̱:������1z��p"O"���h�k��[�LH�HĈ��c"O|z�KZyZ�1�5S�p�a"O���ԇݖFR(E��mC"Oʐ"�"�@CLD� �՗=�j!��"OjL�������A!� �z���"O�x�t�M�)N8�a�!���p"O���A�@�$Ȧ���?��"Of�ZW�ӬY����ͽn!ҩ��"Ov�ȶ	r;9B$�{�"O Ċ&��J?h�W"S-]�:��U"O�Lhv��`��Ģ� U�ߪ�W"O�����%o��h!��ȆTq�"O,���Ķ9\��ْ���*u�"OP1X�H�A@�*ALܧ<�8�;E"OTi��-lA|�&+y�(�0B"O ����3|���!(
<<v�T"O���.��s;ɺ'L���)�"O�dQ�-Z.Lq�
�b햬P�"O:�ⷉ��+��p�v)D)#�fmB"O�4� j�%1��pWh�/R��q�"Oz���D�71l��r�ܦe�d�k�"OTD ��Z.>��[�����EqT"O��f�A����� w�)�`V#-F!�d̍9!�� ���A�Ɩwr�x�'4�lדw�L ��X����'�� q����:��e�[g��9h�'�I���~P.�[��^<d@&�+
���$C�|�H�V�U'@|�H==��M?A �R � .8=yR�в�yb@B�xT��w/p	��	�y�L���"0����3=uD��P�õ�y2n�>	��4��^�(�$�O���y¥��EF �x���r���T ח�y�N�'by��.K�jҳ"ߌ�y2��xr�ˑ��2NX=9�R��(�O>|�V�n����&��Oe�����#�S�� �2�����,�cf��5O
�?L!�d��]}� ��È�7.F�hSm��?�!�$ůY�ȴ`�A��lbm:�I�s�!��&V�F
t�ƈY
:YC׭Q/�!�J ;�����P�
���� J ~X!�$�F=�鞛���ߨlrB�	�$�#�iN�}��`��	$fC�I0�>���H�U�UBG �
�F{��9Oh�ՂP�cI���Fg���"OA	�刡#���1�V�\�nU��"O��w/ә8���Аh�?�����"O�5Y���"#�`eSs��BoH��@"Oh`�#͇)n�>y٢C�/	p)6"O�@@u@�q���"�B��@�tP�PF{����4�p{��A6$��y�)Z�e�!�$[<�Ȱ��L�9 "�-QE�N(�!�$�68v��x#�X�L*G�!�Ĝ�MJ<:Ä�+`��9 aC�R��'a|��$᚝"sʚr��ِ�g��y��]�����ى{���'���y�E�_�B ��-�%�L���"�S�O.�j0��<#���Af��-�$��'r�a f�]*�δ1E>#(U��� RD��J�!�T5z¯G�(�&"Olͣ7/zEH�.J�Z̦����'���n:��8&G�b<<i�CF�!�<Q��@sM�z8F-&9n!�d]>���E�o)�]2T�DG�'�ўb?a��mP�^f�{���굙�d,D��jfD;Al@	x5ʛ=�pL�!-D�0YPoI�u������X(��4�D�)D�T���AH��c�$�?n��'D����X�D�V)Z !�'k~�KE%%D��3D�P.�^� c���`D`�3�!D���D�
�q�BY0zYBBm>D���C/B�T�8��ᓽH<Fq1�L;D����a�z�b��ШAK8AA��9D�$�^e pba�͆@
Ni{Fh#D�P�UnN sP�k�LXp�|љ�� D��Æጏ5Ԕ��d�h�  ��?D�Y2gV6Y(�`�PY�Y�0#� ?D�`)��� /_�p)p��XP�@�k1D�l[�k�q\��g@�d��@�r�2D�,�fN�p�ܐ!DO��.9@�,+D���.��#-�eP �|HuG{�<I��%W��Xh�b �Z�l��_y�'�ў�0 pqQ�OSB�C@e�)3��ȓj�����J�pY���EԦe�rU�����weǥ�H萧K_
�������{׮Y+\$����&B�/[��=�g����	��w��C�I��� �l�E$�rMD04'�B�ɇF�(4A4(բ70as]��XB�I"E�
�ʀ�ٝ��8����%hy@B�	,%�v5�#@\�C�����'�-)rB�I�5F��K!l1T,T��%MT�c����4}� X0e���a�F9S@d(aaN��yR��xz*0Y�k�Iehy��`S4��'�ў��,Q�B!�.C�-+@���8�h� �"O�eے��Z42�S�-t�D- �x��'���JbZ�0�kD�Ih��	
��O��8�H��LDk& 2.��{'"O�<i�.�?�0����nX�l�"O�����i�xa"S��^�}�v"OHcH��?�"�
��U�;4d|��"O�9� J#~|`8��8"���5"Oʴ��K̞e(��
���bϨI�"O��:i@	9t��ؗ�P�?�%�v"Oڙj�h��y��إbR.�d�)"O�=�aD݀*��� �[�1"O��+�ď�J�tH`�EqE��p�"OHm2��R�8 ɂMJ4u+ m��"Ol\��m��_���C�,����3�"O����(�>=3�L�C��u�ĩ�"O։���H�j%�d2R�I�*p8�"O.�t�T>5{R^ttA"O��1�	s�*Ea���
�̽ "O��z4�A�e��m��e��yk�%�!"O�y�A+͗+6�IB���.�q�"O,A�U�@Y��9ǋ՛z���9�"O^i�wcZ;�������L�A�"O���AnT�-�`�
 e4�Q"O�Q��˒�����ҩ&a��"O�e�D��e�4��(��W 
у%"O�Y�ޑ=6^p�BJ D�~�P�"Ox�9QƊ9��s�A� ��@"O^���N�'�GG;O| !0�"O� H:���)y�d%� �1bz��"O��� �"l��y���GB��q"O�5�P퇗���"&
�E2�UP�"O�̊���#J���ʙ+6���"O���qE	,�L���GL���$"O�\;"�ɮ8Tp!��:��"O ��R�U�w���T+�&	�阃"O�x�Џ�+tɜ�'J��W�
P[�"Op��&��w�VL���_�yNJ1`�"O� �e�F/MW���
�<1@�1�"O�y	�F\�j�L��hK�	J�� s"O����"ƃ+sx�����!!(B���"O�yH6 %ݢ�ó�ԹW	�(!Q"O^��3@M��~�`���i�LK�"O�
Ga�V��f�a�]��"OҼ8�+��z�a�e�0(� e�"Oع`W	
.��僂����"OЕ
��C%c0��v�U�&�"O�90'H;T� �(�@�X\A�"O�Ec� ;��AWE�Q�F�aT"O�e���Bp�	��kdjU+7�!�k�0i��ߦ81w�	�:�!�$[oC�� �+( ���Ro!�$�
hs�q�V�ɏ �����{�!��%N�N�0�fT�ez�2��H�!�� ����2�Ee�%�C�o�!�ĉ�G�$���b��G�*��Q�I�|�!���'p�$��ݩu��I�7�O�!��L���i�c�,^���"�B[�!�TLŸ�Yq�A��x$`#!̜:!���5r��骁�=U��	��d4!��
"�����p����c�!��\�G��4�C��*F����=9�!��?��5�.��g p튁��S}!��#yxb��
V�b�8T�$
\�lZ!�@�^���(rn�cu���s)�/J!�ą�?R���%�r�A��퉰h7!�D�)���B�ֆ7�v��D�V2}�!���'���)& �b���Ȃ&�1#�!򤛫I�d�5�	 1����%Z�
�!�$Z�|� %���4�\��b��w�!���8u��D��}�#Ծj�!�$W&ơ�3a\�n	��ߏ �!���)~%"��GS�t]2Dk���,�!�J�vV����.x3��q%�F )h!�DH�B�@�G%8mS�a[6 b!�R�{�4��E�q@�IA��_M!��7/�x��ι;8�ˇi�~`!�$L�Q�@�F�-wIrup 鏮K!���!���0`�I28LȐC���U=!�d��m�Z�W�R3rA
���-�!�DH|��	Å��=% a��F:<�!�$C�@��A�=e�����\�!��U�=�p�l�Q%8���>p!�$�$8>A���	.G�y�獿>!��La�y� �D#�x�&EX!�d���8� !�ɻW��	p �ΊpB!�D�j).]�C�B���P�K�I8!�D�&D�(�bS�CdH}�dhP(H!!�D78�Bu�3CCI�>���&��f9!�D�*���1JB����G�q�!��L�/n�)� X��dC!OA�\]!�Y0N��ȃ�9rHu�R��T%!�D��L�@��2a�B7<&!��  ��U�g{~m���_/nv��Rq"O"��d�X�g���`�K��0y�d�"OHypbi@�!�*�K�ʓ:*���"OK�_����%ޘ8�.�2��;�y�o��*ᱥ�E+��ujv�Q*�y��۠���Alڤ��߁�y�U:-��9(T�͖4z\�H	�y©�.�j�[cg@����J��Ξ�yr�M���B�"sHک���T��yrm$L��Hy���;cʂ@�ҎC��yB�1�F|�Q�ڿZ@$G-�yRJ_�h0�M�_��y�é�y�)�!B�usŋW��8��'��y�e�7K00CdK�N�Rl�D�ӡ�y�HLU���q�e��OV�dD��*�y2�W�T�b�KC~eJ�fY��y"�J�dQJ�k�o�%9�r@����yBi:*��qwR�0�r�RĬ��y�Q]H���d�)6p�à��y�c���L��G����bc��y-]62�l���l��ktr��2)���yiK�
�y ���u)`Jb���y�K	��DI�q��u�TP�B��y�Ϋ�8����eR��æ��yŴ)H�I���ׯ[F\�:�L��y��ͧJ�ڵ��8c���4�@��y^�w5����_�S
�%�Ҽ�y�@�4x��� o9V<�p�H��y�k��Vn����u�D��C�6�Py�ğl_z��g�$�l���-T�<�4$
pE p���N�L�2$��`)D��A�"�{�<���KQQPyĦ:D�h�®Ë_��i�hɢ^��e��o:D�t5E��KCB]0���k�q�9D� �A��7��u��5c��`%D���p�#V��B�G>
���x�G$D�H�K�:a��YW���yz,;5#D��ѷ�ͮ=��,����e�0P��4D���4ˈ�DL<�X�!C,.4(��1D�d�QA�m;��B`�r�b��0D�H[Vg�4]��p�ð3�V����/D�t(#S$R� X��>P���1�)D���@
�9����$	�}��a�3�)D�,c�Θ�	�" ��J�u\�1�PH4D��PR�W;��0 ��HBt��i6D�pƕ*��隱�L<;F1�D7D�l�TςD*�HX��N�1rge6D� !b�N�{�M��@����"�6D�Б�EԷQ�ZѹQ��z��8#�G0D�luɕ�^���p��Z
0�� h3 3D�0�N��3�t�Qh�Iy����2D�x�1mK�)���@�7���B�2D����'�;#��h����D�P�¶O1D����r+�\�$-H�U4�S0D��jn2$*N��F���)7�rS/*D��`�҉o*i�G�6�t{p%D�<�T���Z	��"�� *RUps�!D�p�
ea�H�v�^�B��9Oh�C�ɊN\X�BJ�:C��k�T6+:�C�I���wd_�!g�xP�MK�tC�I35PӖ%��iDZ��3(I�hq&B�	2j>u
�mZ��H�iVK���B��./��v��Pr:���)m7B�	� ���f۶1�d���B�)� �=c�M�5Фi�`�
c\�1&"O&}���֨�.�b�J�A@�t��"O��に�9e�J�y���Z�X�)�"O����G&�@5�#hQ#�����"O8" C��
��;�e�$l��#"O�Pa���,5��QAd��eY�"O���&�x�~Y���ĵzZ�p�"O��8�Ȁ�
2�hY$g+)&�2f"O��s��I�1$P�ڒ�D$���a�"O�(� B�\�X�{�$�Fx�"O�U�w'ߟ-���͍;y�!��"O8�cB�/~@���@��>\�lA"O��I���ҷ���$[�u˱"O�a��̟r��e OV=oF��"O���Ӭ:$\� �u�x�E�	�y��>H>���&jMbq��,��y2㜇B������7�Ap����y	B=^��
eD1N�$rQ#��y�DŤ�x4+�%(�r-�0Mݺ�Py�"Ч�T�3Uc�2a��b�s�<�F�'L؁9����е#���o�<��GHnΪ��a�)u$n��in�<����=��c�����p���U�<1�DK�a�D	QdR'���9�B^L�<�#�/Z�t4�֋�x���q�LNM�<�l�_��lc��W$}ɲ�L�<��$��	F�: ř3q<zA#�o�<�'�^�>Lr���	9ոYPr'�h�<	E��m�z|�""ż�"}�ЬP�<��b
+�hPj�AW5�:e�v��J�<��#��=$X�����/Jˀ�4il�<���I{�:BC�׬�lCA"�h�<�P�na�ϘQ=8�
�c5`⨇ȓ��@ �.�,�b�닛$3�I�ȓ{�������:�0��^�p�lY�ȓ2�.�[��Vo�\85a�1u�̇ȓ�>(��$��)����,$'D �ȓr��0��jW�
Y d(�u�
Ԇȓ>���2U3���%�Jw��ȓ]�l�sŒU����.��\��!������"b*U��n�.�F!���p�R��Ɖ
��x�䏖''z���E"U���N�,sR!�AC�0=�ȓl���B�L"Y<��Vȩ��W�JcW�"2�fy��ΐ"�m�ȓiĄ0
�,��bC��r-މ^� ��U��i����fw4�ņ�?(ȡ��n��kG����Бv`Ǆ@<p��ȓ~!\��LqPxlA���O� Ņ���t������|J�E AR���c�A�oمI�t����4~�ȓo�f���XpB}HT׸�n=�ȓT�r E$
+��Yp�5xl����U���)�Ў'R�@���#y�ȓk*��ᴊ�$n?��pmؿ)k�a�ȓn�����W<=����S��%�,�����|�"�@`��o�T��ȓ:JĴ�����X�ۃ#D�9�І�̂Ѻ�jS#)��T�Ю�-��؅ȓČI0ƣ��tv�IB�{V=�ȓV�>%�aLN�����(��ȓ*Du���92
�D�fW$Ί��y5����p�@Kw�T�/yi�����$ru�!�M���!D��R�<� ���������#b��9J��m#�"O�c��_�^�\1�n�)b�I*b"O�����W�!S��	k 3^V45H�"O���@0!�,����+�^	P�"O���1
�
�X6.X�jL�j4"O���t"��{<��E�Bmh�"O�p��؇]Y��H`�N^�iX�"OF��Kޮb�2=3�UF2�x�"Op�^¦|��ס�����"O.`�B&A3D�4���
 ��$�"O؜x�A�YF��⪈O��L�b"O�(B��V�n�%��G�zMC"O�;�h��:xp��!�jz��H�<a�l
=U�
q�3c?	�
�ɦ%G�<��ٸiK�
D�6�RQN�D�<��V����1�ʍ
��j�nD�<�f��?���)�Ky�ĄQC�<���Ʀ\�főu��n��C�TF�<�S͂XҠ��%v��t)_V�<a7��,ꢵu�͠+/��W�[y�<�(�dg`-��N��U��Ey�<�t ��p*d���!Q 8���(�%[v�<�u'\��&��qa�{ $�ƍn�<�� �N)tY{r�~���Fb��#�!�$�%:�@�$�ԋ
��kU�Y4)�!�_�8�h@�Q`J6R��İ`D�f�!��T)k��=��2v{\`1C���!�Y�G[`h�!dґ=�d�ٖ�!�N�
�

w�BK���u�`!��i}��Iu0�ʕG׀!򤍊^�R���h߳h@���ЍX�!�$�$ vm:`l�~D��%�ݔw)!�Y������{( u:P��*V!!�X
C�켹Q��	( 9 `
U�05!�d�c�~E��	��3
@���b�'~
!�N�Fzx8�������2�!�DE�UX����W�] �b�K��/�!��_�AӆGR#t�2r�-Ѕ\�!�$M9i(�����D3��H�+@;'!�DP�08fŢ�`[-ؑ�(ƶ?"!��\b&J�����D�,��L�*!��Y#j��V��IXRٳ1�!�����C�W7T�$ҷ$��s!��a~��.�^B=�0d@�!�	�di�����R�$�Ò�J!�D��S��dɔ�N�h�2�գ�u�!�d�!>;XY�ҥw�	�#�<p�!�M4��Z�H�y�uT�ۆw�!�Ix�L��	��?8lh�sMےI�!���*�*ޓ/P 
#��	h!��!&-��a�F0vW,4!�&A_!�$�n��ꛓ{Ll`����@Z!�A�K�H]����9u�q��CE!򤚼v+�݁QG�!m���&	.�!�DR<.	j�S� .. �EىP�!�Čj� pQn�*�sw$6�!��P�I�S���Y�"A+��N�\.!�(3R� �D��1M\��sb�7!��J�&�fjL%����>{*�<��N��2f�v�$d��H�_=�\��*BiA����{]�E�!���p��Tb8����F+,e�x6j,����2��YQ��鳔����ȓ��	u"��4Ӡ  A&U	,1��S�? ��p�f�+�M�%�Ή=����"O�P9�]�~�R���D��lp��"O�᳖)�2H#"��4�$�"O��2>Zy�I����y��L��"O��bQ�Y�r�V�ׯ�^잘�6"Opy�6��22����mҗcv���"ONq#��r��s�-��z�B�"O�x�2&��uܥQ�L)4I�"O��s�B}�Qg���5��"Od�!�R<�V�gi˪d� }��"O�P`}:x���9<�Jq�`"O��aé߸V��h1!S�]�^�8�"O��ؐ���1�B���A׫�FP�"O:1a�H�+2 ��@�y��1S�"O����[(k�RH;�����I#�"O�};��X�&$���G��p+xPbF"Oh�H�Խ	�!���լp��Dy�"O��+G�K��!�N
~nkW"OnD����k���uM��g�$��"O,mh��8>0tG�U�ݠ�"O�\�5��;m.p	ɀ,ӨyC�dѳ"O��R�� �e���+OP����"O&�ٳ�ǿEF$��Q>WC�=�c"O�Y�l�-�2�Qg�֯`3��E"O�����
l"
�jdH�4F#nA#�"O�P�dNL�IX&�QF��U
��R"O*� ���w ��r���+-F�d¶"O���"��$#>>%�@E(蕰*O�����E`6�gD���yk	�']h
����F�Ӕ�l�p�	�'d�q)5c�����QoG�`0��'&EʥI@(4v`(�7bT��"q �'����2�U}`��I�1r(!�
�'�,U�,�{<��!H�e9�`�	�'�������7�:T�$�\�B���'�(�A��/�e �F�%R0��'��p ��ng �rD��V�{
�'s�Kb�gF�D���a�'�������a�� `�Gؑ	ΰT2�'4<�#�h��A)T�9aL*}�t��'�쉐��.x�b@�wg�u���A�'�&�r+�u�0@�ȍ����@�'�Ja���+-�������dS�'8���"�
W��k�n�4M�<��'p��G��0��ȁǊ?,:�T�'������!�^mC�L�6(_�ly�'	L�Zv�A�rG�ق���$���0�'rrPID�|�4 Ն�:mbņ�O��A�t-M�v�����J@�^��ȓj��e�R+Ώ7k|ݰs�=g:y�ȓ!�V	�}u��� ��>w�ȓ���k�̝�d�J$�z �q��| z�c� S/LxE��B��4I��r�z��a�'3�x�A�<:� M�����	���{�13o��<�:��ȓCO�	@��<C:���+нPOڀ�ȓ2��G��5�,�� �|�8���j�faT0@��)��B#&�2a��+�4A���	UfH]�P&Ǜd{&$��a���S�ɺb�T�Q��R�b�hL��Y�<Yj=�8	�$=4�!��E���u�_�A�`��kV9N �ȓKo��#Q+��o��p��_�MnD���E�ތ��j��6�Rd�"̷|�⠇�S�? >=��χ��ȳ�C�P��u*�"O��(f̓@�`3�Q�{����"O:q��b��| M�� s?�ʖ"O%2`�Q5\��)��e�6m#X���"Oz9��֨���w��U��]�"O��g�I	Z��Asυ%P03�"O�d�5�ޮ\bi)n�^���qV"O�ehCiEL(`jr,��p�lɯk�<���4 ��ի�0� ����Py�<�����9,e\��mSqe��d3�x! �OR��ZT���_`�
3D�3��0$����������2D�h�-݃hRU��%־%��j�o0D���"�C�wE:�[�m�<�n���3D��"!�/�:ya$��X��]��e6D�\��̇�_�R��g�P7��1�w�/D�T��S<od�1A�P.X��qhf�'D�И���[pT��N�X-½A��$D�ȣ�d�	.�l���_*���kW�5D�лE�G����Q-�	2d\����(D�@8wa�T��Y�H�EJ~,H��(D�,j�J��m�,�z�(V	G'n��d�*D���4 P$$c���T�S�`�IS�$D�Y&m��g�����cޚT�:$���0D�Hk��-�hM��V�M�"x���-T��H�L��u�f�q�II> �J��f"O0�`�<i��c3�_�p#��f"Of����#21 4�į�"�U��"O��A�͗�z������$q���P�"O���h�Vܹ�OI�7���aP"O>Y��`J�=�"�a',�"r=��8"O�Xa��� �`H�O:�m�C"O0u� ���^�q��H'H.T�XG"OT\0�¦(�y[��R�)�<$b2"O��kT+B^�+�gN5S����"Oԅ#��L�/�	�@y���U*O��:��J��xrd���A�l	[�'ך�[BmJ$���S�7(���'8mhu䄰=�*���75��'�����獜�����!H,$�
�'��<Y�b� i��,S�(Q�%�Dy��';��ڦ���-��F�<" ���'I��ӵ�~���2r@
f�9�'��H9�Z2S��hӒ�����
�'������7��]���2ì��	�'sƙ��dB�|���xViܓi/��	�'��X����	q���E���u�� ��'\���A͢:|��U�] 7��|��'x,��'`��&��H���B:6!P��'��L0�l�e�RX�t!�0@�9�'pH�r�M<v�
�T��2�����'z��p�'�GR�4�J�.Ol-��'�ZH���J&;�$��lԳ"���z�'�P���>;��hyq!C-��)��'-�QN��)Ҽ`s�/�����'*�DkF�D*7�90@��{����'�j���lŒT ��I��~� �(�'����`�\�*���KI2t�~�I�'p�(�mCd��XxuN�fW��y�'��؊3@��Fj$��D݂6�fy�'�.ztL��ycm�46X�Y�'�TD�'�L�Y��arL�,�A*�'�勶g�u&>Drщ˼Tu�'}�B�GO5l[z���� �0!��� ��B��a$�Q+�f�P�`l�"O>%�D�9]"�=
���y���ȵ"Oܣ�J�6k��tj�aָ/��
�"ON��mixܡGg�N�6Q�"O6�aJT"�@���	V�S�"O��U���oؘ�0�2��<�"O��R�f@{�(�D��D�١r"O=($�->_�,x�%]�	�x
�"O�-@e�Ѣ��@�b��̚�"O��`3$����f���P鞡9�"O4m"DB�&8`V%�@�n�rDk"OR�q���d@9b o����"O�L�p�O.JJ�Nؐ=�J���"ODl��-�9BR�	�kR�W���"O�dr�h�!1l�a"U�˒Dr0�	�"O�HJ��H� ����IJ&v@a�f"O�ӯ�?_ !y�(�-m�,� "O��rq��.�\�R;+�6�R�"O���#)MM02�)�.ݵa���2"Onų�I#Ÿ��.�Q�d `'"O�m��gV�d_� p�M��ā�"O��ŋ�r���,O6�����"O�9r��[*P|3s���9���"Or�k4iʠ=�61�L��+�d��"O>�CdGĶ�=��ɛ+w�)1"O�ȄD��Ur��H���!H<,AÄ"O��Q��1M�h ��!ì�R!"O�W˛T��K��(�<Ђ��KY�<9aj՜���G��7���ƨ�p�<��dJ2���:y�����h�<�`JE,��S��@5b�R|r!�f�<yťH�k҂�1单p� ��2 �h�<Q�R'm����n�3�b}�LI�<9��
�bf��B�Z
K-4�s�B@z�<�Đ#:b�����x�����n�<	ƁǍ5���N�(H�V(JcgIf�<��,�Y�̰+R�
<�֙ .I�<��$�g��B��X�x�#��~�<���� ��p	3�=sE���/�v�<Ƈ������*W���a�C�v�<a���ENhq�DִkV�Y�f�s�<�A- 9.���kA�O^z�01�o�<a��\:�
�Y��I��8�	g�<WH@�sA+�,e��-C'G��T�B�	 
�ع չ�е�w�T�tB�ɩTj�,q"Kʞ-��|��Q�4�^B�� _�ܩ�PS�	�1��T,B^dB�I���	�����J��ٺ�Y?\B䉳ְ�J���!t,v9��͓^��B�I�d�ȹ���&8�������C��;aR�ۧ%�8(�B���pC�	�g�����*z����7R���B�I'I^�����;vHdH0 ��>]xB�Ʌ:_@�3T&�)G��P㈋�.dDB�I�H�8�B��Վg�"�Xd�[$WlfB�	����Es���I��Dd�C�I4 Ǩ��$�۞|4��_SJRC�I�����޼d�۶rC�	�4��F��*';�X�k�6C�I���X��܏
V��h��U�K�B�I#?JD��� �\*�pK�o�1��B�I�
!����,[�zՔ��S,�&�B�	J6�SUeS	
�6��'�K��B�	2Q�@r�@�-�p�1�`�|XB�)� @ +G�FJ9��ȴ��!j�*�"O4�� Gq��	r�*m]�0{"O�\����dn=9����r�"O�$��A�/1zM�5�	�r���"O�H���S#oM�)� j��R�68+"OP0#��T�I�r��ԈAX����Q"O(�h��2|�x9��I5s�i[�"OX�A���%�V� (��z$�"O�1KLD�,�B��h؈0��"O�D+`L	lv�)���6Ě�I""O8=���'���aI��\R���"Ob�AP/�L���"I����3�"O� )� X���J2��~�d�A"O0�� �K�z ��Y�[�����"O-��k�=OіQ��:qӀ(�4"ORT�3`�)����h�#Uͨ3�"OJ4�C-��y�FY�$��l�rı�"O�DGN�>E=vD�Ҩ��{���q�"O�Ÿ!�~\�S'��/g(\�U"O�s0�A BΨi����;O���"O��Y��=56��q����"r�rS"Onh
!����8��IZ�S/�� "O|����k0�塴⒤�"�F"O�x��ɷ7�tPb�'A�F�H�"Ob)B&坖<���{�?ڔU3�"O�}ҧx�����J�~A�"O����׫%����ڦ?�j��r"O�5��;y��g�����d"O���6�N��4)��P�NZ@p1�"O�lH�G
����C��ǣM�u��"O�2 Is<<jSoێ\a��
�"O4u�S�� XDz(9`�Z�r^�(1"ON)���5
���.��49"@�A"O�$��b��9yr����d�쪥OHZq/� Z�z�:g`�8H�R�x�a D�p+g��P�\	�e
�o�6�#�.3D��f�)<���@�f��p)�f0D��"eېO0|�QЦV-Ӫ8S�,D����ém��T"�l�Y�\��r�,D�<���1z��;��H,��*D��[B%�2��P��&, �d��(D�����0Ю �ǏN?+ȫ�H)D���Ѫ3�L�"v�����P5N(D�������U����HP;X¢|+��1D�S�14 ,ej�P	���Ū2D�T���N�J[0���G�V���2��0D����B˥f�T<�!��WѮ!��a-D��s�Z�!�NH��k�7 �r%� %-D�0)�+ԧlj�0�N41�B����*D�@P%#��LѢ"iܾ�yV�(D��3v%�Z������ֻx�xو��&D�L�DhS*~l"�O�1xA:u@#D���,4ҦT�6�w�9H�?D�ܺv灠6 �P��^3t�<D�X���΄]$$�NR�@�+9D���b�̝ ��Z�E�BȪ�9D�$Ar-W�,y*�)c�p�b�Ia8D��2虡C�t
E.Ӈ!tX-r�*:D�4��I��5c�A:�%S/~D�8D��s$�$aƬ����	v��iBL7D��X�/�-E���d�~-༚�K D�$cŎF:tءwF��=����)D��"�ԇ¥��qZ�Š!D��Δ�S8�I ��6�(�8Qh-D�� ���L��`
eR�G�k��9c"O�(YC��\]FI���_ �0"O� ��Bʝ���(	:P� �"O����,�7�B�x�GX�pͶ�QS"O�5�]U�V`3(�|�:8�"O��5�ȮK*X��Q�%8�]1�"O��)TAU�{"�y5蛢Ny!��"O��*(��$�mڤ��0�"O���ĸ��!m��4���'��'�!�dV4�rqhՊ9!�p��	��T�!�� ,rT�T��6k��2)C=�!�d.QA�|z�LG�Q��kQg޷#�!򤌤1\ʥ��g�!������N�!�>��P��F�'��xČ��!�d�,6���a*A�6xLd�`��0U�!�L��ԩ�wߏ[n�q���ħ0�!�$�W���*ڭw]�l��&B/!�dU  ���cT-�ԁ5�^!��@mp)ѳG����C!!� M�J ����d�ȩq�$Ο|�!�$�d:Z�b#`�o7�=qpI+�!��8c�V��"��>1\]AB�']�!�ɠd)vذ����]R�0A0!���HR"0��*^,?��=�`m�!�d9��#�h�p2��ݤ\�!�$G�&>X}�1����H��LFm�!��Rmz�B�(ӧ��uPaO�!�I;�"��r���7�ΨA��Ǯ�!�ܕ�l��@燠��)�e�ǹ �!�ݼCǬ��@�C�jw���r�ȝ|�!�D��w<1�q К7�N�k�*�mo!�$�"2���-O'Y:}�gcߊTc!�$/���eы-B������;CG!��D�ډcA����ph�5!���`m܌��̄�5��eH�(!�|��5!��*v���q&Gݱ7�!��00�4qzb�a�^(�f���!�$����Ƕ&��&[�P!�Ћ/�0���R�l�u�W-2�!�DW:N��P2�\-d ����"\�V:!�d��V.�S⡋$��ePJ�6�!��B�'�Xk$��!A�)��EK
!�D��P�������u:"��1hL��!�d��Y&�B$�#|Ћ'ɚ�r�!�d�9sQȬ��aJn�J8)''*�!��X��&��!�x�pg�m~!�d�����v.C"}��� ��d!� OE:}!$O&O�
����V�!�Ĵ\5���hW�,�hd蒢P�!�نz���V�	� �I U'�v�!���Nwl�AA��62��ys�Ռr�!�G7�*(���	-��}��oף�!��1��YUGA,Yޜ`���B�}�!�*4����F��k�Lb�&�!�D��dɨ��Z�X�"ɠ��|�!��'�=�a�Bb֨l	6��

�'��!c�N֭&`�,BF�I
z�*�'o(��t�ʚ6D���"K�o���#�'��8*��Y�l�R�
νi>�8[�'�M�5�9��虆��1Ҧe�b"O�qQ��*@4z��u@߂�4U��"O� bϋq���� ����b"OH���(�|ܒA�.���5��"O(t���sr4l��̈��ڽ!"O� H9d	q&��+|�0=��"O��s���
��ԡ F�P_(��E"O`��ī�I�5�W�N�:$ p"O
�� E3s_����L ��eCp"OZh���Z���k��w�N�ʒ"Oz�0`�B�4FD%)PiK�x�"O�e�sF;�D�ZD'��
����"O�I�A�Ρ~\�aJ���*�!e"OX- �]�xʚD��.{T8-�yB&R2�z�C��
/���Ѩ
�yBI�w\�0×��,�s!!��y��ֻ)z�䀲�I'tI�l�"l�ȓH��)��B/�R�8U#<Tl�ȓGU�q��S,(�Yb�?(%V�ȓ<2�X�Tʋi+��J� ՘م�R�n9v��0\��#Õq3��ȓF<�#U�Z=cP�jeA��|��ȓ5H����F�1�����AS�g�T��	� c듩/0V�PEJ�"����%��hDmU�q*f��Ql+Q�,���F���Y�
�e*f�"�Bڣ���ȓx7��s�a�:�bl2��F,^������gj��00\�`���M���ȓ:Zfu���Z�L�6�0b� Ԥ��ȓK�<P�hQ7!F�Q��49y���W{0�ˁ F"��!!F
�2"���ȓNn4 uof��7@˶���ȓ=WL�k#��:���[3P|-���X�m;	g`<��+��O�H
�'~�Xb������ &L8�q@
�'[f,rB-Z-
4K���%�P(�	�'XD���q��}���N�@l��'���XB	�t�|��<�L]
���B�<� HH+Z"�H �LV�����|�<�SHB�=d��rᇮ�\Eb4 Lx�<)�j5h>����Ф��2��l�<��CU2qT��K�� �^�I�_�<����GĄ���G�%8Ra�C'ZD�<1��Yt�Z�ʯOw:Ѓ���}�<)�!�#Z^-p�#i�ޠ��Nz�<q�+�L�܉3���3A�� �PƐ@�<Q'*��?���j�L�����y�G�~�<��D�8�r���a��9pZ@�'��Q�<m��<����B�9^(�Qo
R�<��%^�<�h-@� ؀%����F�	v�<�K�'�hDIQ,�?x�T p��q�<Q�ɾMɤ��Gș�RT�KcFo�<i$l"�lP#▫M&ĔK��k�<�G�N4d�����+�
r%�p�<1��� �D���y��씔{Y`݆���aR�N�޼��(��mT.�ȓ2c����H"L� 1���u4�X�ȓ\�P{f'�#v��D��]	B����C||֢޳l$���	h�̅ȓn6�)�)�*t(F�t��};���ȓ�����*�h9�f�O�dQ�ȓN�HB���q,ly���X�v���ȓ*����%C:Y�q
ٖo�lD��WH`X֬�%Gz�b�F�9e����q���C�K�'F�i����2�
Ԇȓ2�,�k�oZY`��Y�>\X��wZ��ik�ՃR�͵R�p��ȓD�<�CAԐP�2iK���7� a��i2�j�'<?Ε�`�(����S�? � �lNJig�
6�4�9�"O8�`qjӺi��RȞ5F�`��"O�q1��F9{�d�2F*(r:V)�"ON9�%�X;q��1S��oR��r"O�P���8X��isGF��(�C"O��@·8�Ҩ8%�'f�K�"O��'�ҟ���B����r"Or�猉�{-�E�i�h`�a�"Oؠyl99,%X�ǝ�.bvu�4"OP��ר�n8��@{�,��"O�� ���
�<%�0s�a��"OιK�)6|݈�97,��}\�X`�"O�7��[\��ҧJãDH��q3"O����պK����A)��e�f��a"O���\Ś��G�;�ؽ�"O����W�_�)��ßc�n���"O�U2R�Y<iN��O�3Ƙy;"OL���ݶH,8�`�3ݶI�"O�ӓ� ��L0	� rf$yE"O�����4l�7�� �2�c"O����(�9I�.ڦ|~�)��"OF!�U��D,l�!�V)Xi~e�"O����L�:�"ܩ�f�'\ZZ�8%"OL�S��I�tm`88&�(k��-	`"O�)3���$��k��
"z8M�`"OnI2��4l����lxt	�6"O�e	͓v�=���C�!�*�"O��BR�������n��a F"OBqQ�^;a��g�s�Z�"O~����D��|�A�^+f��*6"O
�ÃF����#����T�	��"O[ð�B�d�1U>NM""O"�(�A.$�2��Z�kI����"O*��I�v|`P�G�6]0Q��"O����r�F,�0 �~%
`"OP��"�1��R!�Px�Хs4"O��So����I� ���o��ٚ�"O�e��cH2��+Q���5ؔ�0�"O����m��'.0$�TGXt���˵"O�dcG�ƧR�m	'H�U�dL��"O�8b�V�e���&��j¸ӂ"O�HJ�*ۭ�(q{���%���"O��#�( #�%�%�v�u"O�Q�qDD�tM)S�N�d��t�r"O��� �<}r����ه]X�#�"O"�`�KW&=k��f.7S��2"O��󲥄�QfT8AkJ���9�"O����L�*1D�ªӔ.4�5"Ol��� Q3n��p�D�h��se"O��"@�#|�9w*ƈ+L,Pc@"O�����/c"��ƕ868�t��"O�H����:��a��$O�,:1"Oxp{�h;F�9`q�֘��"Ob�$H�n��� !�	���"O���7AR�od(T�� L%-_J��S"O�$�!�F+�r�Ҥo�<zHh�*$"O2�ШK+$"hAX�n^	C�(��w"OT����$,8����I/}�ڈ8�"O^��"h_�8�4����0�p�`"O	Z��;4E�%�BǏ43yD�r�"OlD��*�PFP�Ғ>��b"O��P��C�D�t�%���b݌��R"O���(FU��jJ�:����d"O4)�ݤ0a&��i�*	�@�9q"O� �H�I�3%>x�����|z|��"O���u�x<0+����]�
2$"OΕ��!h��K�HD%��H	�"O�=Ȱ*�zh(d"wh3���"O�I�$}��Z�ԦutT�V"Ovb�g]�������4	m��j�"ODA��E�$-�Q�@�L�5j�=R�"O4���+E��I��M���aP"Ob�2�l݅o?�MC�0E�ƀ��"O^(����u"��y�H!�N�"Ot���A�(�-��g��V`)��"O,)Z� L�p�ىt�H9ZD^�i"O�I�'T����& F��hMh"Or�*O��@�"�
e@��bĪ!"O����F܍j�H2 K�躐a"O���w�U@+�� !�S����"OJ����ˍJA��ّ��%�2|�""O H	̂�<n���voX�z��qQ"O��	�]z�֭SM�	�E�"O�u`Ϟ���̳vbE�c�v� "OPD�X%bB�x����2�Hs"O$��v�O�*J|��D|�`e"O������(��u��	Y�p���"O6�Ť߃6�ʌJ�?l�V��"O`xq���jb-Y5�� {��]x�"OT�%��P�z��fl�r�*�9"O�sg�36��e�,
��Z�"O`p�t@ټE�.U�C���@��IB�"O"@97�� qRj��%��M�Zu �"O����̘4���H��{�<��"O�a���E+䞤b�e������"OJ�s`صb��i�˛8&���"O2##lS|-8�ϐ:���"O����*@xڬ��r�No�#u"O��'L���0�g�;�μ2"O|UP�	 �~�W��&Nm��"Od����Fd��䃔�� -�y�F�>W���@!���Lj�c5�y��L/4���g���	�"�Js�˪�y�O#37,��q��s�5@����y"ʇ�׶�Z�ߚemF� �V��y��S�gX����b|�m��	��yB��dp�кgi��Qf�Tj��ȝ�y�ʈ�Nf�(���+^�"E˦�y��:`�|�kb�B	Y�x��(�y��׏My��3��̏R0	k3�ի�y"�Ş/@�,�!�L�R��r&	�y���A�Հ$�ٳI��ĩ���+�y2m�B"-��ɴH�t�A�g�$�yR��7C
.�ۡg�)> xA�o@��y�/W�P�Ǐ I��Z� N �y2e*X��݋2	J=,2�kq��yb�O�X�	u)κ"h�5�yR!6R�$�]$�쐐BY��y�́<y�·%�<_�X� I���y�I�Yۦ<�%���VN�X�&G�y"�@��*�dG4~4�t�g��	�yrET)#�.u�
ț"g&aPv�ӱ�yR�P�����7@Y�%�P5�yb)̛P�
���R�L���je��yr���l�����ߤC�brᄫ�y*�60l*�ȑ09��4�'Y��y��NQ���ğ%�884���ybCZ�V$��M�p8R<��F�.�y
� ��
S�^~>h�+���G�|"�"O�������6�|-	Ҭ	f�l�G"O�왧��<}�Hj"L�0=�`�	�"ONH��ϼ~�xbq�!>�6I�"O�q{ @���I���W�L�1f"O�,�"���`���X>H߶��"O����(?��PJGl�v�:��D"O*�x�@��z�A��>�V	T"O@�q��]]����5ʌ:N�jL�t"O�)�_W����gL�:j�=B"Oey㔱+���q��E` ��B"O^Xd�_	ߪ�Z�
�
A�)U*OHm�Bώ*kb]���_�c����
�'M&i!�e̙pzH�ʵI�$]8�C
�'"�iY�/���U��nA<WZ����'�4��"�~x!�֡V��x��'��kDI�*����
�L�&1H	�'Z� 0acK�(+ ����@�Oz�5s�'�6�aQm��C�*��O�"DSؠ+�'B���NI�&�G(��ISd�Y�'=�h���ׄA�hu�6M��W��X�'9옊�ՆM���3�
1]q��
�'���cW�q����u晸X#� ��'�����H� P���PO�ْ�'��Cؖ
�L f*^�E����'�t%��h��j��˦�Qs����"O�i�A��1S�>�(�'̖z����"OHT��iZ8	�M����A�E��"OZ���G���ಫŋ8G�a� "O��#hƬd���i�70���"O�}`�茑sI�1���̳q �ʠ"O��X�Ξ5-d��#�ӻ26��sD"O����JВ� )3� ׀_��R�"OB�9�Ɨ�r9
p�e� .<4u�$"O\�+0��4���D�*ND��"O�zU�:+�ȹ�NQ�@|bт�"O��X���7B�D 3a�I>R�(e"Ov�	E�C�hڀb+�Ge��4"O��
%�Ѡa�����2X6�; "Oz]�D%K t\��Wf>
���B�"Ol@C��:�'O�i�(�P�"O��Hr/�"1	��ۅ!�$��&"O>�@+�qt��#�=72�3"O<�BpH$:G����+ �y
�A��"O��!P.9�lT���G2Hq�S"O������V�AQDCJ�h��23"OZ���j�f�Ԩ�H%UP��e"O�9bq+7���@G*1� ,A�"O,U�o̼4I�|K4'�s�h��E"O����]'����FДkϪ��T*O��3'�;M�}�G��fGV�8�'<u��E�>�*�k� �b�~a#�'�$ I�@�V��]Svp��'����B��48́�E/��C.y��'�t4�w	Z(w���!&}Da1�'(�-тk� \�x%�I0~!~�J�'��8�d�׎fq�%ʊr.VI(
�'��E@��_C��"Y"�0)�	�'3H�	�^R��-փǺH���
�'d�h���[>A@�	�z���'+bE(S-�� �����N�5~�\{�']��F���T��瘟D�� 
�'��8�J�>!t��c¶O��1B	�'b�dA C9u�X�����wUJ�C��� ��h��d��P�7 ��vvdI)R"O��haÊ�$ab�BDh|`�j"O�%	�Y%��ƨZQJ�U��"On5C��!f���qi��^=��t"O��2��/�F^�����8Nc!�D)[̺���K$�4���H�� E!�D&�,� �Lڤ�L�y$Ȁ5$!!�T7md�٦�5!���B���Gg!��F�p������9a�l��
JOb!�D�1H�
�R�߉P��V��!,+!�d�S�x��=K�����<A!�D��j<U�e(lw���R$�87!��>[�fU�t��J�`5�0&!�П`�½��./}�Q��T-!�%?��@pT��.m�,�4HՄ1!�D�(o�����ƨJ��԰1C/6!�D��I���c��\�����(E��!�D��|e�x���Ht��B,
m!��v���т@7:K'2	!���B�̭G�-X�`�=	� Ȁ�"O�*��C�D��Xb4ORq�hm�^�xG{��I�GW0���ĽvؼV�N�cn!�P�M�B-ZE�#Ծ\y�.�.Z�OJ���
1#��պ&�SN��(W�ǭ
M��d�y<h4�ʨ"/���C�#:��c
�'�lst���w������:\&(�	�1&Q�hi*wq�����O|�p@ե�yB�Y�`p��V�@y.������I��HO�n��ź�\���@��w~�m��"O֭(R�)o����Ѡ�ZW�$"��V�zhaz�F�l����l�k)�������y��z����i�� �R�e��y��K��e�Iӌ���@����yRD����a:��~�llz�դ�y��9]7@(�/�
 �
[`�֩�y�]_ܭJ����(H�B�W�y�cN�O�xC����(B@F��y��T%y��"�'��6���I�7�yeO+{"tc�l^�Pp��N��yBd�-G��s ���;��)��?�ē�hO��*<Sl��e�e�"�¢!͌�"O�q�'��u��-*[�[��p"O�,9�jB�zY�.̀\�:�c�"OP��u�]����'���b�\"O��J%��r7ʩɀi���1�"O��"��${�P���14�"O8xj4�_�)�\����	`���"O�y8��;X\�xU��#0��J�"O)� ��+>�D�e��7��h��O��=E�d�����B�;:fJ�9��>�y���L�җ�\�.��̩ìB�y �0�`=01��!$!�� Ѹ�y�$=��k"��$i��1�kG3�y�W/i��9�n��vP��!L�y��$��ŠR*]�������y�K1,\ܱ�Z�>`z�3�Û��y���m����E$0z��S�-�Px�i��8��̈́13�LBs�)0ք\�G���)���/ģ���񐪋�jwB��$2�n�X,�F��:)f8M�Q��m^rMF|b��73�<�'a�9XݚK��H1lG�O~�Dz�O��s	�bj��\$��@qeX�[M�u�ȓA���&���sDN9�c�\$GR=�>)i�<Q-O6�"?�K��l�ҵ0E
?���Yp R}b�'Q�IF8�� �yP �D�s�fOOJ�P^�'iў�S��^D�$���T��H�:�B䉓oS�� �*�ܕy㠇P�<B�n\�I���[�q�֑B��E�@W���$�<��- qF��b�2B��:t�]q��~r�����O����
��F)���1�2���rVCQ��!
Ѐ J耖"O&<1�L�aN�ѻ�B�qi3bR�0�IE�S2�y�B�s��2D�R*:>Qa���$�y�	�d�Lؾш�eh@���'���@��jr�18g�	PD��ZX�Q�4���<��4�O?�"��ˁ"tl��e��'#�d\��A���D{��IS�	E���!�Q�sYX"BQj�\G�tnפ:������9'u���O��M�'qa~ �!o�&t��̓�6��âIM��y�	�>r�������x���0<Y�I?�z� ���U{�����6�����Qp�A�el ���a6��58�'�hX������V�^�E��
�(B"��8��'ƚI�����i���CE䊿��9���D8�O��("C�M���d���,W�\��Ɠ �a`�꒾k*�H���]��p;���,�S�4�T-(b,R��^6?�Tũ�����<�����4V�4apt��<�t �g/��L��{������I���+��U4zG<��t(̔j�B�ɣ=Y��(ЂtGR1[��	:Q����hO�>1H��w�5,�:ow��@%e)D�0ciW�@�����F6Q~jH�T,2��&�Ozx�d��b�>�a��OKJ��@"O� �a�y�)�'�Y�f����'�'��<�s�M9 �hr%��E�虡�'��}����8p#�gH�@#|}�}2��G��ħ+��4�w!�`2b���T�g�@���"s:�P�y�ʉ�g冞AOd��ȓ�v��!�יsLh3)H��ư�ȓ��&�T���YxE]\>��GxR�)j��V?ԂHX��Lti����V{�<!�nC�SaL�H�V<����$]s~RR�P��I��ȱ'���F�0�OZ
zpC�I�L�"ǯ��_z�](a%G}:݄Ɠ`V���0BH��i�±)��x��]T.Ր4Ϙ@�X�Y�B*e��ȓ)���%��#n>�فÔ�j�VAnK��������!�չ��U�&�� �O��y	��!��(ɤ�
���Y0E�$�y⍄=Mf�����ϱ�U9�����0>�L>A�	�c����7��]P��9�Va�<1b�S#W0*�k"�:)�*L�p"�[�`���tW��X�K\�b^�E���	~ZP�(�+D�41'�$Y[F� q*�Y�H�XTl'D���I�K�z ����4Pb
�@'H%D�JT����T%1 �G�f	�*)D�|rc��4r�P��"K��H���1D��bD
^|� �l�2���-5D�<��o�%>L��iB���h?��8UF �O�扈	��욣�خ]�Lx�R�I�a��C�9�f���_���g�I�ui��'���HCb�I�|��B�v������?2�Dͨ$!�e��X�?�a�A,aY��z�C��:� 1T�b���=�� łq��$�"A��8�>�`%�_�<ѵ��,s4�JC�U�����L�Y�<���ޠ���L�%vf�tQ�<�§]�}���SOƍ���3�WK�<�"��?�D0�s@m��c`F�<� ���pI�0y�P�U@�_L��"Oj\r�	4�J�;Db����h"OD�Z�â���Hs�?Z�HX��"O��z��ިl���2j�����w"O�9��3K�*(��	Cd��\�"O6 tjH�o�jt���"��}��"O�b$B�9U}��HƠG� ��i"O���!�P'f��ո�W�p�. �"Ofi�¥A9K�65s���v����"O0�r�U�TP�#���E��D"O�9��|ä]��CD��'"Ol��e�Zh<����L��,��"O��[ԉ�S�0����|1�@��"O�Q��R@(�y��̾&&n8�V"O85��a� #��Y�``�<��Rg"O���S	��vh��1 HJ�X%"O�!0�aI8z��XhW
�6�U�"O��Sn� n�ԣ��9&��!�v"O0�Iv��("މ�B#�ɂP�"O�"@	�Sh�;6�@*rl)��"O���sC�F�@�S��r
~�7"O�L#��_QY��M��F�K"O��c\��R$N"U3�e�"O���)�(#�Q!�$�'z-b��"O�
�ٟ@��l��C��K�`��"O(��
J;�NU#�!�9a��d�V"O(���i@��Yc��z� d"Oư�1�͘n׾�Ib/۝�i3�"O�mSb�nG����oT�y����`"O�l��@��4�
M�*�hd"OD9�˗hr |8`	an.\`�"O��2Vh��#�~�x7�\0)�$���"O~0�ċQ�k�@ ��ӤT�f��0"O*-Fc ��P2���#Oމ��"O@� غN�궠�EX��X��"OV!��&A8���� X! ��c�"O �{cE4 �޹�O�n��W"O��aK'��`v-�}¦e�d"O�(
��+'r��@�L��IRd"Ox]a�戰�>(� 	�>��s6"O�	!���6!���ÀW}z��l D�|yp&�j����)��(*qn7D�̓��"yw�}��%�!�l(gE*D�lJW >W �|���U�<K��٥�)D��02��d��:`��>��k�$)D�(�0��A|6� ��N!3�⁣cB$�O��IѢ�pՂaOW�-h��e$x��x2"OD�Rd�H�lH��F��	�N@�"O�\��aÐ_�T����	b�~���"O4��姏�V�Υ�N�mՒ�"�"OF ڧOh:|:�.��@�d�"O���Wg�n]0s��Jx�~�Q0"Ob*7R;���E�- ֜���"O���F���~!7N@>�h8"OJ���[$C4t4���
��%��"O��C�
B�r{p��$�˝]�&aX#"Oء;��P$e��A���^I�"O��i�g�!ݰ�0�i�4g��)�"Or�"	��[|�`�5,��E�"O�x���:[rF8��A�d��M{�"O��b�ȁ�	�CgM[�
�*���"Ov,j�G�e<�
�=�(��"OR@� �ïG�j���Ǫ=��$�"O(�9S*[:�n�9��ǽG��!��"O� V����?t ��%II.:M�<Җ"O���L?�����Й���@"O��9�ό�YN1�&Hݐ�H;"O�ȉ�(�XXE��{jTi�"OxAKba
g��ps+�1	��"ON�#d֧U;��0&��"�"O�-��ЁGڔA�C�E�7q��"OV��G*_#>����͓<V�"O �A�K�kvQX�+K�3B�U�@"O�)����U���Sj�!DDz��"O ź�Mڿ|��h�)R�_G&\�"O�����_)����!N#2�2 "OP�:ce��C)f�;��Q�F2"�Qf"O.EK��ɟq�<��KB�`��"O�)"�@$5�N	��7���Z�"O>)��e�+},�d�\�x����"OJ���n�>d_t�j!��$e~�$��"O0��;G�r-kq�� z5�G"O&��3�ո��Ԃ� �R0�({�"Od����/g���&���xˢ/Go�<i��V 	2��0�DG�}��GfC�<�f�p�>���'H&f��	e��x�<��͒��B��@�ÏUc��@�'F_�<1�T��` �*�'��"QX�<A���|��=2���Z0��1��[�<Y���e�F�i$�J |�8�Nh�<�gLƀnb�:�΅���T���g�<��ڀvy�J�VYRn|�H��{p��3�넙[f�Uᅲo���ȓ)}�����z��`c%N-��$�ȓh��I���]�1ne�Ń�$8)����+C�K©��pR@�O�S���ȓV�(��Y1�)7 �����ȓ}	�p�dU6:�Tt�!��	L�H��I�8A3�26��р��)��l;� K�T�}�<P�!�V�'�bP�ȓL�D 	u����A�w��x���ȓO��0�!�hP3G�%]L<�������ZjG���7zͩC�B{�<�&#�(ec
 B�	3�<��'�I�<��1(�bl��Ɇfe���l�I�<!����p�~���@)7㴜1	c�<i����j䃲͙)�:��3�^^�<��F���֘H�F��3���Z�<9㨑�#aF�x"٠\����L�<��AUd%
�cdP/��i+ZS�<�⡈�[��I��F�؈��4^t�<�//�R�	�$[ C����E^�<�/N�w�*H�B� G���R�X�<��*X9��9��Gֿ)x9S�a�(|	)C�=O  �g��L����C��2��騰�'�0L�����[V<i;��8���5S�$Q1o^��܃�'�?�RxY�ì&���27l6�H}d�+!����`J|�K�,޲���A�l��qp�[q�<)U��2L�\y��.�q�����]�<�D���?�L�1qǛi����S
z��a�a�PQ��#t�	vMC�'o<\;R�ׂp�`!���>G�i��O����
]���?#<�rf�(L���"d�/Zt���`x�p�`ġ(nr�v�!}5�= �돑 ��!�p��eΪ	�7CA��Ы����dп��?z"+QG~e��\ppi@�˖V�'[��z��ZU0�i�F^�˧d8d�H��8(����Q��h�c�O��S!�J��A��M���$A�tE� �c�����4(�+"��X�_�IHԅq�bEW�ӹMEօy��E@� ])vΊzr�]z���I�����aP츸7�'\����143t�Ԍ�B>(���T���SscAMǐ�P4CC�	H�I J�06?|���ID30����� ��bW*�5]p��	F0'��pA4�'��l���p��ģq.��8��+��7w6��[{�v�{�"��Z`m̞h�T��Ǻ2<V p�� Wh2���=w��S�֘D>xUE{r� ����%N}=�d�E�O�Dm��\ך%"GO���p�a�+�Ȍ�u��q��ʱ@݌$����hO,����Fat;�\�/<r�`��'f����@��Ѩ��3N&�&?�вc�0E8�ʅ��Cży��	)8��k���6OLQ��Z�z�a~A��<�zt����r\�g���c�����GI��9 �lƗnLYY��9�vd���jl�熔��y�!�
� �� I������F1��>�晰M�Q�����|z��BH�	�p�ȳ�W9.v�ٷg��,������?/tu��B}��b�?�I���<����J�l�4ɝ*(2Te�E��^�'��ɰ�� /�,�{U冫-���F ̮ �L�*1Wf��!D4��|�lJ#Ɇ�2#��@FI����ɤ�>Ճ��|�*�Ye�7E��|�4H�J?1w�O�Zž%��[�@�V�=�b��(�?A!����If�D���]���[��H2�۝e4J��$QK�P�AݛD��P#+]A��6��(!F�85��c>	K��:6���ۨ6�� 3��[�A�!S���.T�!�!y\�P�C8|��`��^5�W(��I�4���1���|˕:��q�f�	�E֖l��Kދ�Px�E�S�Z��wOD)J4�|��ҨW���`5N��{�N���	L��� 4m�8	�=��i�-v���Đ5n�<\
TL������,B$�ԑ|���T*�+2�!��4P�I����@T����_��N��8��l�����IÈ��qC�L#[g x1�H��J�!�8n���@�m,q��TdܔSp�>)L�;���>�OXh@P��-ZJ�P3�� �j�PO�`an�Z��#�ϾU2��j���5S
����5�OЉ�C��x�d�Do�]�NK �'y�l�d/Q@��x4��C'8/�8Ȉ���Q�����8.�<����9?Y#g�:�8p0V�Z*4��`�g��m�<�Q��H�4{��Ǧ+ƠI$��b�ɏLS�U!��HD6�?10��׽i:�S=ƚ��3()D�0���9e�4�� �#*�����jWb�[.O��pBlO�ȸ���&�zs� ��,x$��]����n|��#���:�|�j�C_��n@�gW�?Z
�c+����?X�C7� �)la�kA�Y:�-��e�N8�d"�떬�~�(ǄW}"n���A�U�+5�,��A�y��5]�Z�B��'F���/K���=�����(&�xI�(SER�9N|��b`��&|4d���C��M{Ej&]���H�\���.�G�<i��8'���a��^�A��T(��� �T�[_��ai�T�O$����{��hPm˚vQ>i���&M;�%�� 6�<����y��pж�ӡ �l��-��F]�����l
8O����d*�}���!/J�E�p��T�d�MU��p<�6�C�o%\��oƴ��'s�x�u�8d��#��[�X�X ��_����Q����$�	>�J�)��L�g����#뚳w�'�Z�å疴e�4 &>�����m��}`T�i��Ԣ�T�8���KR<u�͈�'����I�m�0ZgeVcFZ�	GoׯvԂ풢J��tTd�O���J��p^j� �O|��V�WV���W	�3��ȍI��p�!ը=�!�K�**��{�,g�J�`�`H��ŔC�{�����U�Z-.��0��Ij��� $�?CbzI��	G݂��#'D��yU̖'r��`!��1�"y�Q��T�x0�A�����'���	��T�>)S�R�N$������а��G8��c����X0�2� GhZ�!��ᵃ�=-'�w��uZa"
]؞*�ɛ�.r�}8v� 8N!�Gk |O�۴b�,v�:ܴG�tա�K��ԛ��WU|ه�m�DX�/ˍ)�����,�%R��d�?��ѐj� ���V�OJ8��� N~���
�MIt`�
�'���rʎ�Oq��Q�REu��
7�/����t�\���d<�g?�(�R���+��p1:��Gb�<ђ�͵<1���҄���֮D��T�sC�:�>e�J_������H*Phd��A�PZ�l�t-9|O�0�̕Jۊ�Ӑ�Hp��*0C���r�^D5�B��9'Ϊ��ԡP-Q�e+?K�����	R<tB�e	�a�O2�"dBI13�2�3�+�I8�'4�k �@�^�`#��z�,��� �ԊQ����/�g?�ŇI�"��k$��	xi""�X�<� p�2Q�Ø��8�w#�/}����'�0��!��|=�����'�����m�=lݰ'�8Y�PB
ߓ{`B��e���'�����c2<��%	L�sv���@��y�,��6�����
��|3N<C�ê�O�}x�	�!h���).>�Q�C�E�"���C��!��S8����6�Z�A�^x{�O<!�+Y	oa�A'�"~�	�y^�pvMް��$�:��B�I	k.����O*J,����+*�B��<m�p�d̨2�h�Ӣ煭8�pB�	�#����ϦI��O�$�A��-{f��uOF�zF�!x���>4�VI�ȓ2�d�@��(N�f��E&�����]"�xE2��a�	��$B������SEO�T� QlǍM�l��ʖ�ڲ��C���C$
�x���ȓ!��@م�kurd��\	OЄ�r	&�1F 0Qޚ��eF�tT����xl�q�Wc����1�ԉoVp݇ȓ(д�&$9"aW�ԇr�Y�ȓ,��x�q�!d��as�?<v���>|���TT?DDZ���x���ȓ7���&o�N�hd��h,aH��ȓQ��8�AO�.��q4c�54�l�ȓ(�n1�ӽc��yz֠��2�0���_h v����.%��8t0���h����_����ǤX�C�"P���ƅ���F*�\�(U,4S]Z���u���$�� �\ݫ�I�G��0��i�z�SF&ѯ��5�p��1�����t��,r��^�pQ�1�W���fTp��J�� S��92�2IU%A�	����Kϲ��D�K��T:D��&u��5�ȓ1��Ӕ�GC�T� �_'U֤ф�0�,�S���#�*��Ν"�����v�P���X�pJ��aCl�y�\e��D-��)Y�%�Q�G����U-?D���Ǝ�n�"���KB)[ڱ�ƥ:D� XD� 0=�3����|��e�$D�xOGm�@��]1@?Y��B#D�pz##��S*���/��pPp�"D� ���74t
�[�O &��<Z��=D��(�?��!aB=m΀Ч(/D���R�DGv����KH�PY��,D���7 	�8*�ԁu��x�W�!D��"��w�6JRJܔ0aP�j�&;D���
��Yњ��$���FdM�2&-D����X�-b`@x�㔵%�t%�i,D�P�r���)��1��l�$7�X��� D�X���)c�:�)'`L	Xi\�h�L8D�d�s
�~�lf#���>��1�,D�<y���3TJh��J���Q��+D����&�!<8�)E��22����'&D�<�W�Q=8�)�l�5``��#�o+D��9�o��CA���Rw\��FN(D�hh��'p��R /A�¨���#D�h0�T�+ؔ��M��_�DA�h D��*���V`M��d���)ؗ,8D�J�N K�Q��J�{a�IXpf9D���`ϕ�D{<48��$#ۚ�((D�lz���![�E`0�
�%B(� v�&D��q��VG����ej�VD<�ԣ+D��Z1@����y��Uf�1Q1�?D�(�U�_W,���ׁYi�p�:D��@Ԯ�:�V0{b�ɵc��C��2D�� |(%#?6�lI��!O ��P"O�B󮞉& $�
1���tu �"ORt:�#�n���6:4β�t"O��צ@P��a�`_+-�؁
�"Oڡ;Ch��)� a�Rb�c"O�|I�"�%fH�7��XH�q�q"O���
V�Im�0bD���U�0�k�"O�5g��yv8�ȇD��|�H(h�"O���d���I���/X�4`�"O����j��b��s��tI�"O���&D�?6���N�z��u+�"OT��/^���A�;b��!)�"Oʸ�[2�����ݲJ�\��#"O������V(��93c�-B}�-�"O8���Ts|��d���2o����"O�#Ԍ�s�DC�-��3z% "O(Ԃ4%Ǣ8��$cħ�=I8Px�"O���`8��u�f֔Y�IB�"Oؤ)�J,��=B��"�
d��"O&(S�d��<;�Qr��G9z�T4Ȃ"OB�ʃ&VL�lq���]�S��`�T"O�5 #�T�}+,12�S%�BT�W"O�)u��p�pŁ�Ek���"OP4��G(*D~p
��ԹD(�d9�"O���e���;JTt��$8v�a�"O�yx4�Ȱ1{2}aT�H7�Ȩyg"Op��vB@�~Hu!�<}�z� F"O
�0��C�7sf�D=��Qʧ"O�@P!���k�L�2q	�
���C�"O$$�Ϗ7��)�Ҭ[:~���jC"Of�P����r��͐+�X	��"O�]��k 4`ڂ��� #�l�"O��L�f^�}S�͇(yiɂ�"O�����D*1�^q�$a��l2T��"ON��%�Q�
t�:��*DD�i�"OX)[2'�#lp]Jr$�j�̱�"O�Zt�[�|�(�R�c�;�"Oj��g�� B��$��!."b5ӧ"O�D(�άe8v�0f�ۆ	��+q"O��+�^���� oőEm� z�"O��9�����a�Ҍep.A"O�	bs�� �d<qd�.]f�tp�"O�LЂ]�0P�Ԯ�86:��+A"O�ٶkǖC`$�k����<=9��"O�Z e���f�����+��P""O@@��`��*��A�������5"O� WG˓U!�C]�L�\`(6"Or�rd��!$�C$��Oݰh"OT���G.ksHر�2���eIXJ�<1B#Pz.��4k��p�Q���_�<9S�]d(^���C	��<��b�Np�<	�-;;�Ny$��xkL�x��m�<)�f�5lZ\j��� ������e�<yꖐ[}�I��ĶU�2A@G�X�<� ���<��h@SKK2 &b��5 ~�<)���^$, ���FJ�9����<YЃ� �l�b�@;KUZ$��Is�<�͎�MY ����L=���˘j�<ɂ���>t��+������i�<p�T�b���q�K:	��� �B�<�6�B(L
@�R�OޯY6�a,�g�<Yg��A���*0m��i!��j���0�*�;"�mR�剑.2䋰�:LFz�i#�&^�b����D�X?�҄ȋ��O_ 4b`�J�kf�-"�#�9S"\��I�G&Aa2�L�D@z'
�K�� 8�b�� �b��d.X� &è�?	� �T[YA���b�3ғ_[��p��Е��j+ ȑ�	F� A@��[��<�r@\�^Z�O��4�r`ܸ\^�᠄��4��	��HW<tF�M��d;I�PP�M�`���x�l�� AB�ЈA���G��2�Z��p�'��Ht�ޠxHv�(S,��0!b�P�G���Ǥwީd�ԬRv A���N+qC�%��2�O�1��@�G@u�PΛ����RD�ޫE�9pF��H nL�GQ�:T�Td0a��N�����BL~�	�IyxԠ򢒘�i
�ҿl���=W��:���t�$G�ѹ�o�~"�	ɡE(��1��\� �Z܂�I�9w��Z��f�֥Z�
,�ʩ�g�'*.ɈԈJ'�Z�hF��O�B� ��I��\"`/�e��e�T��㥔�T�B�A�d0醥?mZh�"�`=�Ċ���(��D�&�%U-H����;9��mQ�������Hy9Rk9<��}A�3�
�۔A��!�Ι�3����Aa��N i	�+|��,˓TD�q��B����'B&�O���G���oƸ�: B^�+��F�V%�6����F�$�!��!P�mvbMz��9^�j�`��(���O���jG3O�Rw�֯
� ő�E�.?�]���	"]���V�9��Ђ��|ZW탲)ʀ���)ٟ+NX�¤��,s>4��X9?��鑲ŮLд�bg�3��O�����-e"���( �w�j0��Ol!�0�U�DZ�u�����%U�H�n�O� Aj�.=M�-�e��=h6�"�ቾw7����]�ް?A����4�E�n��)s���M��92Զ�f�K�0|ږ�J�|xE�#j|�"���I�<��K՘�,T�6o��!E���/-.�^��O�x�^;ܸ��es�}
b�FTuJ1��LɛOܦ݆8�0!b3�ӛ�:��G! �иCG� 0�"����#�Ol�0�̼P�Z��򥁯d�X00r�'�H�:E�ʔ����'N\�@�9uV(�b�=d!����'�\�1���{u�G��t��M�0 ���6"�R��O?�ySׅݩB[(}�����r��	�'N}H��?�4��㊮Pep�AT��\���:B��|"E��e�Va�b���1�А3���ѐx2)Y���-+vg^t:��2��հpH߳cv�~�"�2����b��.pЌ3�����<�B���/r�OD-�kMEM�5�Ã�,�$���'L�=���,��Ik"j�����Q.0���:_�B䉗(^���҇.4����( T�O^`�CY-S�������7f��c��P�蠲k��d{!�D�%:~,q�B*�
V<b��K#&\�A���RGy��+,��l�}&�HA��+���aܓt*0�$�����XHF<��@n���q�D?>�����B:	���%���Ą�:���8���&~�u���^�f� �,O��!wa�lH`���C�>	V��R)�a#� ǳ).
�c#�<)��^� x4�
ߓ,Rax�$B�9t�"�/Q�e�O�0:实�5����%���`H1 ��C˦
&b�=<o�9�a�7.��0+A:D���$��g�PtX̕S��<�FE�
L��h.OJ
�f-<)rb�x2��6,��n�$d����D��<�(��	��-���� �P�j��Q�-�u��D.r�nTc0���E�-���x���P�$
4#Er�l4�H��
C��R&��x�>���+	 U�w�Y�Dz�a�'�0A2c�D#[�|�#�V�+�̽"�2�F�uMV3�l���4,`�њ�/]�	 �H	�'��:�_
:�'>�3T�=&0`�i��h2��+pu��q$���~aV)��'�X���E�c�0yŪS�;ᔸ�W��-6�)xr���V�8�O�1Xҏ��R�6��O�d���xܚ���v��PY7�L�V�(�"o�!�$\�"��M�
Dt1F�RAj�%	�Rg?��Q�t�8��0�S鼛�!X�522O��K�2I��h�<�0��&=���A���is�0��	�XA�S��T��Ę�O�Ӟ_M̴�}��؏.J��@�"S�М�g�p>ISbD�j�I�zDX��'�9�>iJT��)G��ą�~X���qӧŰ=����l��HP�D�,X5�O_����1��R��9��ixh���##���Yc<e��,Z�'x�9�eGK�z�L�վp�%�����'�N,#ӄn��5S�O6��)�O�<? Is@�C�R;$E"�'A��"'R)��!WaCNi��qWDL�)x6��wL����=�g?�!O��z��l�9�6TI�n\�<�G�F�n�	��6�u�������k��dI����W��<���;�AQA�Z2��=і%%|O�����kUJ��EĤ�u�Dmмc��Q AM٩I�B�)� Q��KݳL`������6���{��DS�p��$/8d��"|*4�\�Y.غ��?0���k�X�<�B��a�#V��	FJ\�MΖ,����F�=g� q�'Y�>��z�z=k�i� [�@�q��D�AV�B�I� �r�G,-�X����Σz��dy��I��Ȅ����1&s��'�O>?*|2�WP �{�b�& ft�9u�H0'r4��k=_�-�U`�d^1�"Ol�5�U�Aq^��Η? D�5���I�G���Ī+�Q>m���__$�9�5h\�<8q��(D� �G�S�o�8�ɲ�:${]�g��y�8������S��?y�hT>q��M��&H�!��i�⤇n�<�5�	�U�t�q�J��BB�O^�<����,�|��o��/�f ��@�f�<iG�T�1�0iaF�	.��P�3.Ib�<�3)�!���M�i��jT�Q_�<ap$_�\ڶ�*�c�$���K!�XM�<��@ZO�����K��\{��Cu�<I��6.Th�kW3=���ք�w�<1 �9���(�.@�t�& �c#s�<����K�e�	�~��A��s�<�AEnİ17�g����(�o�<-�x�AՁ�-Sm����A�C������@�QM|�p hY�w9�C�F�dh�Q���a:�j����C�	
T�v��W���:���H�>R�<C�3T;f��6�۽*�`5Z�,��6WC�I�`@PB􄟪+��,��EG"��C��#*
�,��&�m��aw��d�C�IW��!j"L��=A%�7UB�C��7-5^����7��A�aA��C�I�1Ƶ�c�i(�	�GK	��C��#hC£G(Ʊ�2EpC�8M�0�ҝCź���eƅj�B�	�p+�E�k�?6E�$iG�FD>�B��)xyĊG�u���膕W��B�I"�fx+&��0c�n=�c���jB��/߮��q�J�a�J�
�Bڅ?]hC䉋{�"bU#۽l+J�`�O�|C�	DS����@ɘ:�P}x��/�C�
8���y��	o&�;�G�]�8B�ɈN����)� 7��ر!iD>?��C�	#E�>���B���p�gď5�C䉩K��5[� 7y�DMА�B�[��B�ɧ*aq�.�l����+[^�B��7MX�|�ĉ��Xl#���`3�B�0PE޾8�B4C�A
�`��B�I$o���8�	"y:LA�%�S%�B䉏X��*@�� [�0���L�?R�B�I(N�%��L�c�J��c�=pDB�ɕ6�V�� S(Z�d�1Ng^B䉤	�D�!�����p�ʥ	'�C�ɰ r9�3+:� 4��H�R4�C�	y�4]��a /3*TK���iE�C�+��8&I�,��F-PJ\����¦)�Zd�@�=e�2HQ��".�i#jK�j�!�F/U�d�c4�Uʡ�fH�.H��O�Z�+2��?���)~�����J l�0�2F�ƚ*�|%Γ~ݬ ʖ,�c�l��*O?�ۖ��>pgAh`���[�Ȉ�$O�8mȨ�gFP(���0|��hU"&��Qq�T `�̭:��;?�T!jI_����L�@�a����UU-��@�%h�P[�#��B^�EQ�O�T��������g���~J�ɖ�	������<�P3��<��)�ڟqЃJ�S;���"W� ����í]Z����CQ$z-�O<��E��}2�)�s��'���´���=qF���͉>a�*@�'U��۴���~�S�'4*��&߈j��	�gi$-�fAme̓�0=� @����`���Ǳ�D�Q#"O@u+R���m��X$"M,"O�����^�pVxPzt��>Ed���"O&����*Q��0�o��.>pE8"O�,ʣ&�/^z�j����K7��G"OT�J�͢G#R؁�dO70����D/�Ş\��<��
�'m��qa$�&?{�]�'ۚ��'z�Y�EM����|F��kؓsk`1ઐ�u�HTd�3c��91�&V ��ODD�9;çK�8��Y��PC1��5 �B���_,�6��j)乊��@ ���S�DI����@�3��U"`��6H=�I�X
�9� i�'��Ӻ[��E\|�3��+_
�D�G�]]Z���G!=2�i�╟�>�����X�0�҈ђ*.�Ձ3hK"t)�Qs
͘-� �IAZ��O� E�"���t��@��w*|�ҳ$�+f���1���>B�L�2�!S��|>iÃ�8P �R�B�/b+�T�p`/T��Ç$�0 ��u�B0t"O ��dB�c�@����#?�|�"�"O�8CR�ƻ)���ღ�+V��Z "O�%G]�dkbD��D�������"OL:��߈\\����ă�C��E�"Ot����+0�@)�A;s���Z$"O���M�;8<��%����h�"O�1�EeK�!�>�!#�Bo��p"Oʡ�plY�'��|��G�JU2�W"O�$��� 
�,��Q E�sTBq��"ORy�C�ف]���xǎ\H���U"OƄK"�^�d&��ql '#�H��"O�p���X5hUK��5*�*�"O��1���	zƸ���\��tCG"OL$5�Kc��h�߰K&���"OʅQ��Ȁ&���W	D�e�Vx�"O~�I�%��m�"lR���[�B���"Oҹ��̜-��x�0�еqZ9K�"O�īF<|����#��a\z	:�"O�=:���5$ލ�wO^7^UT@CE"O���H�!,�pj"ES6�r�q�"O9�/W�rJ�1Z�/���"O��5��,G���S����('N�S6"Ov��D�W�^?$��_�N����F"OέKŅ_rE�u Faϲ1����"O:P!U���	c�}�a��"O6�е��k�f�K�=�L@y�"O�-��bôK,Ty5��3:뜸�c"Oe�%�բ<���wĂSD�Qђ"Oz70��r3�8[3�*q"O&I�5g��ac" ��C"O�[���%1p������#tHQ�D"O����� �BE0@��4E�p:�"O�y؁�ޡI��g��
���3"O�8����kjܠ�'��8Q�|�"O:��b��(�D	�c�рf8�졳"Ol���F��B-��� ��m~y�V"O�u2v� j��y1�o|S0�Pd"O���+QZ\���&lO���"O�%�F��%S���Dd�>���A"O>|���$+�j�VBޑG&:���"O��1�ʱ{�F����F�d\h�"Otd�ʜ��P�{������H�"O��B����$�2�e�dCU"O(x�0��%@,��SpΉ+W�n�B"OF����R��1�툯	~�j�"O��
��&f� �%,�!\��"OH���&
�%�Q�9��m#P"O��F��}����^�Yߴ1�"O�|S��˞���P�Ɗ!,"|5��"O� ~�H�Wzy��j�EZZ ���"O�Dq��n��f$V96{�Sc"O�P����u>,�����g�
�i�"OR�HG��*;��($"�
�jp"O��9KL {��3/�p�(�"O��*ug�t�z��u��|[�"O�PY�-�*>~9R�m]�����"O�th�e�>M��p�lG(�ذ!s"O.l�Ah��?��A�F�q�L<jU"O�L�֊ɹP찪(�%0�b�"O~����1?"pzb��"IT+"O�42��00����ҫ�;r��"O�Tct�K>$m�Xc�IK�.�@u[�"O�����L�4c���$�1zh��3"OLƅ�wX�d����e_��؆"O��p$��$��)g�����3"O��3@L�O'�	��S��"�j"O�)�B�ӢDAn͋ X��r���"O81BTc݇u5la�G�E�Z�[�"O� ���̛�����_�N~2��"O�y�ā]�l ��ʛ�e��ʴ"Od� ��P ��P��P�:P�}2 "O�<�2�u��"��[nl��"O�!Pl���m���^��H!�"O��O�I	����MP�"���"O��qq�]%)��YW��)�ٳ"O"ݒ�Tڐ�ӔLƖ��y�"OZ�q��@�����i�+��,a"O�ł��3�8U�SO˾7�2��w"O��Q"@(x HQ.v��)��"O����'�.C�ՈQF��\3�@"O�Y�S(�0C�B���R�n Fa�"O*H�%b�V�[��5�f�!4"Ox�ӣ�^!c^y�f�^�u��P��"O�(��˙)���З��l��t!�"O6 �]"w���[R�I!2�j�
"O��*QD��`�<��1�B�=
��"O���-��N�v�C$ɶ%����"O<�i쉥16�YpP�@+~���n8D��P��0m548�/V�h��4T���c ]���W���"O��s��u8 ��6a�]r�"O�9�R'�=D(q��O��@�`"O8(r �U"���#��=[}���v"O:��MH�P�Jܒт��%f XC"O�y[&�#C�52�C�d��آ"OAr� ފ`� ���b'�����"Oh �c<n@�@�izyV"O���+ʙ-GI9O�j��2�"O�q�ءZ8���m�:a��=2 "O������2>0�wM�0�*Qrg"O���$)PK��	!�AV�_�|�x�"O�͘ /_�o�$,3䀁�:��g"OBd[2ǆ�{t<<�B��&T4��K�"OF�HS�(]��}��[�?6� ٱ"Oʜ�����eP���j��>��� 7"O.�!w��i�Z��LGxژjT"Of	���i�~(����Q�uȄ"O|�*f�I,|�L��(���"O\izU LRފ� ��)6��!��"O>����ޜP�
H�'$W�8Y��"OB��NOQ �2GӋeN�%"O�y1DƄ:�"����Q>Oʸx"OԄɰa[,K���B<O�$@"O� ��W%��;�-(�힡;<l�9�"O���w��?b荀��"}>�x�"O���
�!|�
�P��cK-�y2O^��t\c�LȜ#J��ᢆW5�y� ��~=����>,y��)2��>�y�n�*�h�2�\%<��K��Ȭ�y�5\8��T=#��d�����yr�H*V���y�̕Q�r����Ϩ�yBJ0��\���Y�ظT�6�y�'�'(����N��P$�i��l�$�y�9�p��Ƭ��P�r��`P��y�S>'w����̀K'������y҅ě�%b���4V���F燿�yB���B� ��>a���9��F��ybN�R���ĊN�8��3�S �y�πQ\�Y��@�B%y&n���yb	�q%Ĥ��?;�J����y�D�6q�d��YAG|�Bpe���yR.�;K/:�Iǈ7��S�n���yr)�虑�S�3�H�xw�H��y��HyP(�8F��/+����Jݴ�yr�	�Bv�;�X�$���c�@��yRGH�<I��U:n���s@O��y"K�G$���?eg�(b�"�y�숥Q�����(cLۆ���y��8Xư˅I��TfESAB?�yn��z���a`�ʛc[JȘV���yR
�8&Bz!B5*(,!�6�6�yrJʜ�8M�����HU퇕�y�F�d!q#R�Q(����Ĝ��Pybŋ�&�,A�IL�/���K �k�<ᅥ�3\�$��ɘ�0���Bf�<�Q��/f�����˶ lP�{���!��3oo ��n�p�����7E!� Ho���7&�g��$C�c��J{!�D/�W���x�dOE�w��B�ɕ^xh�pe�'�Z`�Ðz��B��aI����.�Ր�c���B䉁1��(P	B{� ����C䉔^F�x	���,0��5���X2SB䉫t� �`�W�p����UA�{��B�I�[g��� �N^���HemT�kn�B�I�<��ȫ��ͪ]��}��Ɛ�FW�B��	0�j��6GID9�M	f/�oV,B䉯h�����MRՃU)�w�B�2U��K�^M��0q�	�:B�I?�9�m	�8u@���]m��D��l,��z7�S��:f��|�!򤅝m���`�G�_O���F�E�jt!�Ę�TZ ���?e5p��e�Xt!򤐩A���Ck
	UILh+Q���F�!��0I:fMZ�g�4RF}���A )^!�D��9���ˈ7Mq��Ay����;L0��S��Z��#�־�y�P�}�4��������y"�6!���s�C2߼eQ"�O��y"�C4<�.p�.5`u�"�]��yRS�@�HT��k~�v�a`[�y��B!!�hi�D
r�LM[A.�-�y�Y�{����(^`��0�I��yR,܌K�����ֳD�sc �>�y�3�"� �%?�z�ӏ,�yR%ȯ,�D\���8���D��y��x�Ԑ�͟A�Z���H+�y
� ��K��"V�t�c�J:].��*"O��X'
�A.�	q�U�L(�Y�"OP���'�~!2�Ze#�a��"O�y�B��LZ��B�1�"OƠZAg�2s��H3d�4k
�]�B"O.<�!�U}j�d��a{�4��"O�J� V8"��8���)�<T�@"O��ھb�*���F\�5z�Ճ�"OB��(Ӝ,�@Z����c���+"O�k0�M$�|�Pc�ȳN��B"O�- �4��2w�Z�<�f�B1"O�\�E�\<Y���VZ�Й��"O�y9B
B�R�ha��ɔCFL�S"OĄj�$V �z`�d��B8L�+�"O&�R7+�6W����*�+?�^�9p"O����_�hn���d��P�@�(s"O��xŪ ok:��S����2�"O�pkf���(d��)E��*�%D�<P�$B�i/�q�鏯8 �k�e8D��0PA   ��   �  b  !  �*  �4  u?  "K  �V  �b  �l  �s  �|  -�  ��  ��  �  ]�  ��  �  -�  ��  ��  �  V�  ��  ��  �  Z�  ��  ��    a � � 2 '  �& %- �3 �: "A �I wQ �W 2` g �n >u �{ ȁ ��  `� u�	����ZviC�'ln\�0Kz+��D��g�2T(���	#Ĵ��*�?YV����y�抋<+�x�ebW=t@(d���Bh,y˗�/d=��#���kh)�Ĥ�:��R�v�	����i_�B���x7'�`��G�V�T��M!��0s*�kQ��bC�HId���-���w�"�����?��j^��9�Ѐ.�6A�3+�M���fM��"B�̋FK�L#��)V6�ܠ#ݴ���O��D�O��d�@4�5��w-�2f%�j���OV�DF����?ه���B���?�V!?T�� R%.ҍ{��%y���?!����'�R���M����~"�YH�OY�j�E��h^�s~�P�8_�)��~�@�(Ola�$ʓ�pl�7�Ki|�8RBŭ,v�C�%���Df�$Dy"▖�$���L�<��g`\ʙA����|�6M�d��<��ҟ@�I��0�I۟���K�d:�"퐶�@�OO*aC�0���1�'�(6�Q�����M[��&�
6�6��(:&iK�i�>G���Q��@ۚmhBEG*X>\�Fz�7��$�D}Z1
%|f4�b��P�(IR�ԇ1j��G�ӄ:��x���M���i��4ڟ�ݭ�v�>̐�%N#?�̩���ך
8\(sC�̦EkDC�u�p�Y�#��e�p���J4FR>�Y7��7�Ms��i�b6-�&G�M(���F�,��&��e	��1���']P�2�ˍ��Qjڴ2q�fd.�T}�e�]!A̘HJ�,�'%>.M��/��4�ǂ��B1�j��8;�PF�|T�7-��%�ܴ9�L���!�=
�p,J3Lő������	�*l����p���ZT�R��f���o�˟��>�&Z2�����D�?�e�2ޠ
 &v RD�Ĕ��?���'�r�'�F6�4RPb&� ���B�:�\Q���˟$�'CR�'N�	��|\�a7�D�e�46�ě$�2�"&fZ!1f2ł�;����A'O����mT2%4^��R�aӦ(Ce`ڗ��e �G�2U��L$3�X��i���D�" T�$cq��_�>��&��Hb�'�|��'("^��	� �y�g/ֹk�P؁v�G�+�F��	���@A�=���&�T�s��4�?	�%�;|�R�D�3\ܒ�hRlIПܖ'�����iӘ�$7�SӼC���67q�|�e�{B�l�SП����59ZM��"�V��� ۴i:�x����Ch?rY2����˕�AƧy�p�'�v�#a�{�N���'�+�l�hQ�����O�j�pƄ.;����
18���O64��'��7��N�O��?JıG���Q�j�B�FX�J��'�R�'�S���|�ӊ����*��Y&d�q��'��f��!l�ߟ��۴���*I(M�n�ۥ��8.��`I��X�m��v�'#�c�<��埈�	ϟ|�'�fC�D��S���2$�m�`�i���f(�7ڇv4��8A+�K�˧��=� �L�7V�I� 
S6-�V���@	�5�(XP@"��;���J�
bX0�|B�������'Q�N5�ů^ x8��3�>vІ6��cy��Ĝ�?������|�-���kV΍�
t��a�
|ў@��I�dw��� �,^��C�f�,�P���On�n�!�M�M>ͧ�)O��T'6զŀ��*�Q�T
R}�d�'�2�'�w�$8�� CPb��w���B��S!�!x �L�p��iy'b�a�7I%2k�x�k� *}>Uk�̏�9�v�1r�T�^|^��g�$v�8��i����a�0O��Gy��]�`*�ڣ�EC���:��H35�����e�F�?���/?A�#W�.����%+_�-F4ly�Q֟����b�j%��b�D�c9������:F��I��M�' �6�bӶ�'+��A�i�4O`� ��ՋSO$��s�o!7H�)nJ�Z��������'G��0�Ʉ����ڴ!U�ХCE/~��l���Ή./t1CC¤�0<�&A�%}S���㬕!0�ѐ�Y����;��Э*	v����\��1 �����MGxRa�8�?���R����'������C��F�cC���=��b�_��a��N�Ӻo�H̓)@��䅓#�`(�2�;G���'�(��4�hO�IXΦ��c�۩[�\y��E̮9+pcZ2�M��/�6�K3{�6�Ʀl"\˓����^:ҥ�.�,IK6Ɵ�G�`�k���O���!S6aze["D�Zѧ��-���r���,�J�
��y�eQ�*O��ɰ�傱FXw�0�bD�d�t��!���lXe����?-#���1&M0�� �w�:�V�,?�1�Aӟ<c۴su�O�1�ԡ��LҰ�̜"ҫN���BV�|��'��'���'���?$�S�V�q�6A��G$(j�`���_ş�m՟$�ڴ�?A6p���FL�� ����@���'��I�L�����(�Iȟ��'���yq���E����l� {�P��FQ�$� 6��j�%Rㅃ�lWʧ��=�THR"�YDJ'yf�p`rCz�d�#���8x�2���*b���|5@�~d�v��Ǔ�ʪ�H���		o2�yٴ1y�:TWR�d>��Oz���Of �EC�
M~��p�D�1?��B�F;��0|����z�	�I�/����� ���b��Uզ��	��M��"�'��]�5B�x�p�_�Q$�T��
֡k|���A����	џ@��ky���k�6-*�{3nL�t6<i�╇g����"!�'�
t%e=
B���剪{=�] �U&Mx^��I�!��Pj&d��<�N��c�5�fh�aKF�_'�a M8�>�[s �x����3�Q缉 �Ōҟ��	ӟ �?Ɋ�	�g��Ɋ�Q*��b �#<��{��Ă�8�Ђ7�Z�v;z��s�H���'Ą7��O<�y�d������	�
<'�Y)��")�ظ[Ћe[nbS��	�<̧M?V�hvN�+΄`K��{R�� ���X.mQ��,��Q�v�c0�'�X�@��ƐPO�R��e���Y��B�h�BF@�i�t�p#��~�:�*Dn��O��A��';7M�Wy2gE� !<�
�FRU�~IC�!�����<��(j�Kn��[�T�*D�^%*�`����?1-O��=�'n���F�hBm�Un@P�%;u�R�#�P6��O
Ul�+
��	��4�?Y+O���<Q�M�77?nR�C�k^0�&���?y�(����f�Y���Ӌڪ3Y������SDyq��"V)6����]N���/|մ�a��+� !B�BG/�!,���'��-� /�4U�H���N��h�'�����>���#�'��t���t@�^�5Mb���K?��>��O.}@�H/-�8T9@L�(#��%�b�	���ܴ)5�v�|�ȅHV!�V�@��$C�Ņ�G�^6��OJʓe`���'�?!��?�.O��r��
	�+0T[�ա�j�2W�8�ӧ�)>�\QVCU0�H�'��=�G��!C��BF�$.b�89p%��M��2qc�5��C�fr��|��1w�]Γm��@Y�_�+�Pa�0E�rߊY�޴t��((*���g�	Q7�P��c�<]�XE�)_�Uw:��?����~�����l�#�L�Y�=	#���h����MÖ�iMɧ��O��	9�vճ'�$lGzD�цD�3��JԌ�����Or�d�<�,���2P�u���I�C�`�K��^%|��eRU��P	DL;���3J<��~��$���s$���'��?F	�Ы�O�)h>�0�DE�Nv�\R�� `�2T:ѡQ�'!<�I�i�+Čhkd�		A���B��?9�i&
"=��ߋC��@�-*TL����)
��I��HO�%�	�gd��Ƞ�VlJ���@�O�mڇ�M+Ol�D(A٦I����l����DI�� �ۗ&"@	�t��ڟ(���H��M��ß(��m v���MQ	P�����B�KGJm����eT�y��@H�tS>�k2*ۅ��H����<�F�ȧ}�@UR�)�
����d�b���*�O�YlZ���Ē7s\��H>Ya@Y��'�z��'x�yB8O�����Y�T�S&E��|mm��'��6�ȣ&�B�$n�Nht����{���<ɔϘ0?��'��Z>��&�O㟸P��I�8�۶��R���!�ӟ@�	9D(���� R>:����0~�������'&TH��TM(���4 ����'���)��P�^&P���#�"fD�b�iоqT½��Z�:��99�l�=%��4u���O��}B��)N,[���"�8��V�����'�͚&��z��f �?��d����ES�OT�k��Q��ˠ˫~p��P�ig�_��Æ.��?�E|�&��iC��ܔ�%�����<��U��d�A���a�@.��h�"�� ^
b�t��
*LO�	5JR�eG�]A�g@Fr�[Ċ3��@@��G�1���Z�d�)7s`�Y�@�n�!��!2ᮉ����(59�=e��ɍ�HO�)"����^�ˢ�P�ȉ9�B�����
����Ol�d�OVܯ��?����Ċ]�'P,��.��K]^m���*���4cq�!$.ư��HkǓ�TU`EB���A)���	f�,����򦉋�֮�F�X�j�]8��!�Non��Y�dm���kE�W��Ā[���z0��+���#\�!�T��u�-D�L� ��6$Q�q�D�44R���-�_˦�'���Մ?����OB�9�.S�;�\3��8��Q��*�O�D�	wv����Ob�
��,d�S	(�T���(܀:��Mʡký;x"�t��_�h�����'�((����X\,0�*��8�3�	�@2v�#��b)����x�џ��%��O��;?���T+h:A̜)�����u��Ɵ��	&sq���D�A�?A0���(�@ڎ���ٟPhFdH!	�E���7�<%�we�O<�&�Uۄ�i_��'�哤`z�打W�^���(Ԙ>(����G��VH��ǟ��Q䅦^�|�[c�Ol�<�ԯ�����0�b�8}sF�q����l܉%��L~�JޔA�Y�pM
-{T�d逵��&5H�ḱ
����XT8����ұ��Oйl�F�O�|F�U�uDς�l������Đ;)�riہiݘg�����H�lT]h������5p�Axh�))$ ��Ņ�_{�Bٴ�?�)O��s!�������O���<�b(R";U�����T]�=�NN�}�b� �<OM,7́�Q
y�G���:��j�K�!�B4�abڻ t���lĻ,�p0m�WA��b#�3�əI����V�d�,a��nBa���5?�%�ğ�������?Y6��2w٦P&8��)��j˞�y"�baW�^�[3`t3Ή}%��-O�0Gz�Oc"Z�t�sǇ �$0H���Q�����.6� < ��Bß��I㟠�Ɍ�ug�'��>�V��sEǧ��ЪFI\q�DP���t��#���\�i��*<O�|�`� �$Q���nRp7f�4��"�	�jq��T�2����Ĉ�jlÐΜ� �-"�X�<=���'����d*Kt�
2!
*1���C�-!��^=�Du
��F��õz�'��6>��T���mZ����I�3�ʩZ����MzڑS4b:z�P���(�@����	����&C�	��b7�	$*��2Љ�*-����%ӥ*޴���ײ:���I;��Չ�C��N�N`��׎E�$K�X
	�*�{�+G�Z���Af�:OXDp��'Ѭ6��YyB�g&0u�q�
+��ЅF���䓛0>�6'�>,��e��·�X��C���8u&$�S�Od�7MƤL�LU��Ɍ� �YG�S+;s���<A��!M���'��Q>�B��N����:'XA8�ɾuκ��3��� �	 `F|Z��O�֜��E9�?�O ��@�zx�����/���	�.*K���p0�Q�C�h�0]�3LY�h�d%笞�=��YA�-�1'�x)#�������O��&�"|"TAE>g���ӥ�N0,1�4B�h�B�<���
�+�
�X���h�JŹ�nB�'�P�}��b��\�"ё@㋧H%�@g��;�M;���?��+&|xwŔ�?���?9���yD��Q��t��	V�^���H��ǩa&D�b,A�A����mPנb��d�|Bf�Y��cl�hʄ	(�N�26i�bB3^���U/�������|�M�p�X��E�q#��c��?A�OH48q�'bR�'��O���'���.^�����a��B%&D�<��0�f�7�B�N_@��D�<a��i>Y�Iy�˸W���w-�t�&����*� �yGꞨs���'���'��֝����I���R!гnGZx�@�%sb���wA�V{b}�v�O
sL���N`	!w��8O�tr'�]�G�X� RAp(��=M[azRɅ���($L#`ǘ9����.n��`���6���9��O~u�@d��>���݊&"B���|��'�V*'FV&E@�ʃ^�t�f�0L>1�i 2Q�\���� �MS���?9��	�`%s�VE�:� �P2�?��.�u	���?A�O����ٴ>��Ѕ�út%��H��]�)#�؃d"�cy6)`A
� ?Max�#?�M3g��
5ш����2#ʰ
׮!���!6��O+f����'� ٰ�U�'!@<��ܜ
LYI�(K`��	�',��`º���y�/Yl3��0	��l�"���6��T6X|�ej�*��|.|��u�i8��'&�/�^�I� ���C�W(��X��%]!`��	џ��b� ���;�NQ�`$4���2bD���&��KcJ�^�	�5*[B~�b�CT`k�mP�0鈭��F�
F���a��6ʪ<�G���.���9v��La�/�Ob,m�y�O���4,e"PR'��6>Fݸ��N��OcJ�j�n%#�,@��\�J���
��6����B�'W������]�y�w��?:}$�y�4�?�-O��;"K��">����a�R	hA��R j��tBK�qO��鉺7±��IeT��EE����<�ËV��0���$v����F�*|%FT��W�I+~%J��2�3��9�.]� ��?36t;�c�8C��w��(�ƥlTL��Q�3���eh����I�	&[]�.�����!�Y�8,y5�^��M{
�tl6��2�>r����'�L+ਆM<��A'�T�+�
�d��A)�`�-�U����T�#�-� �$�2�E��\t�B�
N��(�	�xʸA��^�F�Xp�D%�TH�ȓf�8`���>w����`)?ތ�$�|xߴ��Bd��	�ic��#i�6��O�i0�f��8�����H^Q>���˔�R�dܻD�Y�sXX`��'��$���D�LE�eC	F1���G�)+ax¨���?�Ŝ|�&I^������?��l0�O��y2<��1b��(�hh���	��?y��'_t��!�'�~D8`��1�K>a�0�&�|bP>��� �2]Xc�8�&T�&叁XY���ݟ� ��_<�����!�r�P��J�O;1��(!<\���e��&
�O(@�#Fml��F��:V���(��i(��ᗊn���(�U�=��	��~��'O�>y�	7�A$΢5����FB�>d��ȓm�h�Ӵ���2���lֶf� G��,�'e|}x"�dQ��D�Ux>�Z�4�?�+O�A�,�����OJ�$�<� (�JF� cBę���j��I�k�( ��ӁG�h�j�4bT@Í��y��β�T)!�K˿xs�A&FP�dΪ4�2Ș�d�hx�7b)U��0���y
� ��2 #���6�X4CY�ɠ����'��I3�~��'5ўȰ3b�/�l53��Bl���:'�M�<A�F�`,p�)�
��UQ��FEy2�3��|�����I��ŌX�/�Y�����&M0ș` �c���-7��O.�ŞX�̚&�R7DcT��W$H0\��p�a�4{���;W@A�L+@��@8������c-���$*�R���7��K%�\;T���Q�\��xO��`�<�#�AZ�cl��U.�2=�Ҡ:��?	��� r�������:��J���|�����Y"p*c��	2yq�L��r�0�&����OT�K����iU��;�4X�%�C�R�.(�l�>mO��$�4?{�@xA
O3`!��4F�74]hd�;O�jR���Y�Y1�a�a
�F7\���+_���(�_�	,�8Q��F�hLRgZ�!�Gб�s��2�lx^�m�"I�O,0+�jS�XA��&^�T�A8d�|���~�c���O{�
�;q>	@r���R�����A�/q�'�>tq�c̅K��`�̙x��aq�J�&ѡv��Z/ƔSn��[��Kڀ (�`кE��|r̝���|�#)��F^f5 �ޕ�x�ꥣ�T~r@\��?�1�iӊ"}Z��<w�)A�虯d�j1x�`PP����	�'z�۔i��}*Z�*��V?ب�0����Y�O��y ����`�n��lj�ղb_��'i\�9��'2�'L�W�<0c��=mI|�EȚ�h�4� �/ ��Y���W�c�d�Tȍ�U�r|�O���䈦Pv��PnՌT$���bP%B�b���7��}iF�Z$DD�Mq���D��7Qc��Sq�X`���?WSⓟ���L�O��D!��z�`
]-�4�Z����0
�'�=;�Q��c���8���(*O��Gzʟ�ʓ s\=�w̥W���&A��4D�rQe�&�?y��?I����?��ɋ��}���W#gH���cZ( �h��I	�>�Ss$�;X�!+��"O�4Z��O"![D�S���"�|(��*m"�C�Ȱ;d(B+̜�p<�@N̄5�J�N��Uf��꘸
���	���E{�ቱ!3�Y��̔�T��B�یfƲB��%@� �%@Vf�4�C�B��NL|�O�l�''��@���H~�r��R��g+_�wv�Ub*ԟ�'�B�'1E��nF*a��.��W�ː�:@Q 툵� 9*���0�eD�I�S�'W�X4���E�y{�>��T[s�_iUT�@f�����!��$ư�0<��b�����IR~��݉^��[�DI!�p�.�)���0>I�L'� �)�F
4L~�Q�OCO����*C����^	`u(����m�6��Iyy�d�A^�)�(�f��߻R����e"Ĩ ���IĖhbD���Ob�s�|����bH b��A�&$&��%#w��kA�U�X$j	(��H�~��4�'�[���9�^�`��B�HH,G���ͯzj��� ��|X*��PJ���%?���'��>��Uf�Xb��	V�������J�΅�ȓ4��( L�n�"�#�mɾì�FR�?ڧN�,{ E�X�t�e�NG�!�'�ɟ|.����D�I�'�F�G�r��z�-�V  �H�Wu�l!�f��e�"m˦ǌ�O��|�<�CB��x�	"A@T�Ac��7 

^݊�aٺ h�՘Ơ��Lm2�|�<y �ƦY�%����[Rɨ�@�����''������?��d�,\��3�i�- ԭqQB�+O�C�	�Q ��Z�_&B�h�X�&6I��ʓf���'���N�-�ڀ����K� �.�lA��s(�O����O��$�<�O�lڄy@�yT���$)Ȃƴ;x|�q��W�@ѓ�ߚ,A���ǓOg��z�Տ8rjm1w���la4n��i@
!�rA
>�쬁q-�O8�1��
�|I�\/MHh���N P�����O��=���$�e���a%�"_���!�%ރR!�E�(*�|�v�W�s` =��dơ'#�'�����D�+#�&�%?��M��
�d�/��d�9i��d�<I��?��)��DCc�O4cotp��(H5^蚢O3.����O�9�J�(����I�bY�ǆò��LI��'o��Hs�a��AN� d� � �VP�ǉ O* rR�'4���8Q����$8mq&�K�g&F�jAo �D+�OR�#F[9kMJ� dC_���탴�'�����>Y�l3	#�*(p�#ʁN�T���ů�Lyʟ�˧�?��H��6�RA+�I�]Ip�p�lX�	ßT{u��4��d�to�=r3,��U�Vu���0��M�|�<3�DĠ~��[�O����&�QL0��.T�>pyX��)��|%H�@�-���3���~�I�Z����O��}�� �pKWǔ��	25L�h.6��q"O�Y(��χ�]��404������h�����-Ƽ*��]�j��RU8�C�b�@8c�j�<�eCE����	\�ʱ���[pP��	�j�=I�����u�X���B؏F�Vy�%�3�I�j��$J�nf���%��%G�9K3��=G�J0x����['����;��Ϙ'V8x�큇bƮa�E$�k���F�i��˓!�����?���ڜ냄�K+t-�C�%u+�܊
�'g����K6,
�prD_�z��(ON�Gzʟ�ʓ<D�P��>qB8��j�x�|�rS�ۦu�֡���p=�Kޝ|�#d�؂
w�vM�3�R 
W�8�I��An�`p�ù�p<i FY9f�A�殟���8`	��f5y(�/�Y�rmS�R7�"��D��T[�Y��l-4��ԅ�4�.�� �'C 6Y�'��d�p…�*HS�%�al���<D�#FK�k���3��>u-`I�f`?�dKA}�Z��c1D��M{��E~��/4q���e��O���;��S�'M�䌇D>Qh�i��q�ȡZ;O���I�{W��t�Cr��89c
�cC���dG�C��+�$�<tl[F@u� ��ę%f!�D� m"x����&^@N���O- ����O�x��<=��,�m�
~�AIԟ|r��B�7M@�0.Q?��Q��4���RP�$��:?1����pxaIU�L ���:ʧ6 jT�sN�+G�x|����G�<�'��U97E�^��iU��&MG���J�7l������O�0S�����DC�"dt�^�E��:���aIW��y���0N���F"OѶ��'�2�W�U�^�j�R��	�h��)#"���_���	��ܐ5��$��|�Z�Hĺ<���B����61�h����6��4!�4'�~c�����4LO�-�F��A��V�T�F�$�7�az�Ĕb؜�ת?^��f#��E_�'8V������Ϙ'����J�V��0(�N+d����
�'g�tx �s`E��,ȓ[�"�!*O�1Fz��	 !{b� Ar�Z-$Δ9P�Ա?����>�@f̓4�����OYĈ2e�Od���YA3��7^��!`�%Y0�\#D�_@y��'Pr�'p�CvkZ>dw��!�_}�O�Hi��^�e���!'�(]P"Ҋ���27�l�E���5R8�%>�2�T�1��1��Z�:A�a>�P���	쟐�|*n;p��D����,�feOD|yr�'��a�'ĂU��բ�
Ǣ4M$eC�K��	�M�T�V�#G2޹��E
CE��H�.�����?/O�˧�?	�eDj�*���\Kx�����q ����:�D�FB
o?����!�Y"�6�S�~e��G˂�-�0y1!��p��I�F������o����ȟ΍����8R�q�T�@^�(�<O�=�S�'�"������P�z,�֏�%ߞ9$��Y��݆�sS�)`G)ѓQ=0��dw�� G{r##��T�*�(�P%M� ] ԰���?I��Q~�����?a��?��"\���O�h�&H�(+�i2ਗ਼�R���"�U�1�aR���#�$Ҳrh�'ei��n�I���Im� �cB&7hz�˥n�XX�])�@A*O�d� ��?~���ד?ɸ�!��N��[����Ǉ<��X(!�T��0?�E@]����I{�'��Q]���a["p>�*�f�D��$˖{ݤ�i���E����뇐dU���Uc�����';�	�1�	1�,�5+C��It�Y]��}����؟�Iߟt��Sy���%X�U
R�J�+��`��X �M^3^2b�c��^�cd�`�(ц�Ɍ.T��*�q�f�&/�VDK�L��tblA�I��^�@9˓|��D�	8{j��R�,%�tP%&Ӯ~טA�I]�'s�;%�޽�i��OE�wr!3q�<D�2d[�Ò�����y3Bs�B�<��i�[� �⮑���O�hi�� �Y��$�	�Fߖ-*�^�$��̟��I>r�ƌq�F�	A��Iѫ��V�OY�Qa1E�B������I�T�ʏ�$A'Ex���8Q\e�O�t���؍n�J��DI�C����4��OX���'�B�	̳i���1�,-j<��7��W��Im���d��s��v���>i�8a4k4�OŖ'F��&Ǖd%�dȖo�4]G�-,On����������fy�\>����x�V��I� )�F3(*<(�5�J�|GB
5�*��� �j?����`U�{q�`�m+��V���ہ.J�|�2��@�Mzv�I-*\�\�w/�13സ�%]�c�L���L�}�q��P�eKtú�K�DWef�ڕ0O�xA'�'p7�GlyJ~�˟� .4KꙩM�m"6#DVr���"O�9@�	c�pyR WWS�p퉳�ȟt�h@��'�Y�0��+��Je�Z1y���\-�R�i9�t�'��Q����5(�ŻQ��M�r�x�e�}�,��B�()_0�rŊU�4]����G��LX�* dL�Oh��e�n��laT/�({���PːLt��Hō��L�ΈRCa�-��s�����f�*f�@h3��j�v�b�H�S��p�*O���!�'�=&�3��`�����l��AiOg4���+D��g�Nݬ]r�J��}��B�O�Fz�O�"P��nÂa.�H��O˒[_���*�i��t�I?4J)��ៈ�'�ʟd���+ H���'��ydD�2�+ϊl�8�(ͣ?4�A�DfY3U��x�	? �"P���C�)��Ev!%5vZtk��ܣ0�z`���W�Trj���	�r���@���DGg`M��KI7g"���'ړ��O���gʺ
���߰w1��"OV!�QK@$u���f
�� T��Y�d�ٴ�?�)OZ�C*AN�'Z�<��#/h�XA����4dN@",O��$�O����8PPA���U'F�U�g� �M�'ZV`)��OÉ>^��� �5qxTE|B.�1�"�@���IN�h� �~�AEJ10�I���N=� ��N�':�H���?I������-8d$��g�f�,�{B�����.�O�!Sn_7�^��`�ʬw6�12�'��	b�|��Ѓ"i���A�K
��ɗ'��'��'MRP>��'_"���j##�<���'@�0��O#=��4�O�͢5$�LS�d����"�����d�NOTL@H|�4d �y�����>���x�!�N	�&�'�t���?O, +#�'���O��0O��"�J�R|�AE�%S�Щ���Bx�7��Oꈩd�O8�	��j�s��.Ei�\c޲T"��	�b�f���&$x����ӟ����j�p��u�'2�O��3OV��	ƨm�����Gڋ	�>A��*)n��'^��P��'��DF)l!���ug��<�aϛ*%�����^J� ����&�?q�O�̟���#�Vx򮟚���O\�	�O\)�� ���#ğ-<¨��˟�1��O�������m��k $�?7��;�1�O�p,K�B��a�<�lZ�<Y4������I0�?q��r�H�:�YBL�����h5�e(rYB�'�B	C��?Y�����i��z��?7'Q2x�)�b�X��z��X�;E�)p5cF٦��Ubx��4mD��#���I�����CRhj�G�X��A��!W��in��Al,��8�4�I�l�S̟��D���ϧ@w�H[d�$���� ^��G,���s���̖'���	xӒ��Ky�'i��H��X���`�cϋ\fxAw"OJi�Ƈɜ2ZX9#PIZ�JF�i���'3��'���'W�')�:>�0�J��~"�46��3:�H��4�?A���?Q���?���?����?��U�f�!ƄA�:���@�%�ѽi��'�B�'br�'���'�2�'4 4�2��.P�4<YŌ�h���q�hz�N���O���O�d�<A/�V���>��/E��=вMJ�h��?���?i����*+}J�!&l�[����Վ�nZ矬�'������$����O�deS0'��a��uA �H'R�H���4�?!��?�M>�)����kf�Cn<v���Ճoi�	����J�<ٷ�[8V8�(޾Gh� Y�k�<q&K�9d��@�l"8y��j�<yQH���쉦�^%��}U+�^�<��@
?z��2$
�DÊ�(v�L^�<��E)@R��)�>b�J9��b�P�'[��'B�'�T�ig�40����
-x� IV�7M�O��d�O����OX���O���O"��hr\�@2"B.*��(@ ��\mZП��	�D�	ݟ$�IԟX�	���V*t��N��X���a��5Zʰtj�4�?y��?���Zo���	ɟ��	����T�ż1�$Y��eT4�6��$�+�M���?���?���?y��?����?�6�JR�p����>K��3�1%��'r�'J2�'���'���'\⋕�d&~)�o�P���r6M�O����Oz��O2�$�OD�d�O���ί��� ufS�[�Nq&(�~y^m���@�I���I�	��I��H�I�-V�X���O:Hi1g��@5{�4�?i��?1���?	��?����?��C�=P�B�&z����f#�)n޶Y���i��'���'O��'�R�'���'�\h�%��?q|������d����rb|�����OP���O8���O����Oh�$�O��"��ݎi"<��u�	D�Tʀ ������Ɵ�I������	ןH�������R0����^�8p�3b�MS��?1���?Y���?)���?��?�aM^y���@�(���23L��������py��Ӡ/�z����9d9��թu�.�nZb���O��Mk�w�\(�ՉY.7i��c��"X q)��'���7O|�S�%�}o�M?QuN�-S�h1��yX��re⟤�2hН���Ч��k����8O��Zrρ�	�,��a�H��1R�'��F�	��M�f�f̓�� d RR��%uR� �p��?*������'��'����?A�4�yV���ǦT��`Vc41$U�1��<�r�^�X�R�\���i>q�����C�?O�����hLl�u&�0�Z1wP�4�'�b�<x��ܥ|/~���F�d�v��O��n��"��,;���'ɧ����#!�B�	VL_�4�/���Ӱ8O@�d���_�O�R�l�;��ޓG�xםU3څ�SM�;}�5�wi����=A���d8��PYm� L���1��K:\���6�����'+�$����|�l8�64 "��C�<!���M��'�>]PR :p%�uU�W����֓k�-��c:?	�)^�0���{\��'�%��'/:0�B	�+W�dp2!J/�2	�'��@��Qe6�u�QJ:|�j�P�y�m��}�`�h!J��q� m(f��3�^�{ǋ���ٸg.��#� [��.vy�gF
�*�@�k�搁!�<LB�tQ�(́u�5�.V��c�K+��L�a
կ�,F	� �}:6�Y27�x��p/A7R��S�'S<T���`,Y70��"�/8x,� �O�7�ۤTn��J�Wv�+Dǈ?e�i�	�p�gH���������O����\�3��'=��|+�H�hpR�����G��	 !j�۴v���?Anگn�*mi��ޘi���aE�S�S��_�M�hO�Y~�����6_���dLՏ;��Tx�c@�G�F���!y�XȨO�w�00[4j��%o�#tP�� �� vt@��d��m���VF�[o����1���/c����Ԫ
k�Y!���g_�������
�n�:�g�X�Y�6dZ� |�(��l��L��a��sw�ekE��b9j`�GG���օI@ƃ�3,��U$E |X��_�pH��A��VQ� 1�B��7�%	�Ć�'*\Yԧ�>�1#ւ�=1���$�[�,r��
��S-_Vp,�PΝGɼ7��O����O�)@wyRM��F#L�hB�N�,���p@�S!�?a,Ov�Q��i>-���۠D�. �@��% ��:5H�eEğ�k!ŕ��M���?�����G�x�%�ԙ3��℁��J�J�̅#�?�d(c���O+��':��TL�jd� �`xh�0��m�����O��Sch��%�(�	ǟ��XU�UCC�`���+|���?᧡�T~��'���'0B��B~�����Tyl�>[���'�0��,�d�O���?�D/8Jr��ގ3�]{�+ԯg|��a����'��'���'��S�	���BF��[]�a�EcM�hLT�E؞�ē�?��������[� >�<1��1[�>IC�N$�������O����O\˓0�\	z�Oq���C����	O$�fX�N>	�����D���~2lɂD�0�`!����� b����D�OT���OX�F������hOO��
T�]�4"�BӦ�2�'�RS� �'��˟�č#$FX�G37Z��`��D}2�'�bS�ؑ�ƈ��ħ�?�'30xzqeQ��x���j9zJ>q)O�9@��?yQ�ϔ�6]ld�ǅ�2���!/�ON��Y�%�iD�̟8�ӟ��$_��r1���7���uEɷE=rP���� ;�Sܧ20: Z �ȠR����jS"hƠ�I��x�4�?����?	�'K#�OBQ*EB���� ��3%T\
Q��Ob�)§�?�ǋ�MpJ�c��f�%�WDQ�s���'v��'����r.��O��|�lS0��%l��S���{�
��%�'�i��6��O���OޜIqV�V�ʸ3�V�8p$j���Of�$B�C��'���I�x%��Ңdp�҉���"I�� ��|y2��0˘'7��'#"�'�£ـZ,�x�v
{<�Je�-r�~���S���I��$��K�	�� �	?P�qA�J��
:���
PS�]z�ר+U���?���?����?	Ceģ����?[H4�`֏sk4D"1H��?���?1��䓉?9�"�(�Cl�(=��q�+D�I�}�S��^����/O��D�O��d�O��d�.����O���I>A���a�ʎ���� ˈ
S�����O̒O����O�`��qM���d"���HY��Ώ  :1��Ɵ ������ɡh'�l�O�B�'���$��c\<Q���U�`]���'�'�8��t.�������ƯPvN�0 ��:j*���Տ��?-O ��D�O����O��쟦˓P�pc'�W�X�Z(�1��?q �#���?��2=������NQ�DFF1��j�-7^t�1P�0�?i��� �?���?Y����+O���Op���i�
� �A�+��ܭ����O��s��0�)�'�?���CE�H��@�v*��p%��?��?A�2�Y`-O����O���q�j�&�;��U�5L�1ja�2�<���b� �'�H�	����	�L��͠p���d�7�P,G�Q��͟�1��~y�'2"�'��'3�I�Q�Pt���Ol1~�\�𨐫T~�I����	����'�n=���mR��:�t~�H6c
:y����D�O���?����?�RY�D��  q�J
m_�\"��Y�BH��mhRY��?1���?�.O ��e!v>�H%�>�eJ#'I�Vقлv��O(�$�O��$,��O��d�&[�J�I�t8��&I�5?l��k�
�6��?���?�,O�h#�|���d{h���.[� K �I����".D�h��?	K>a���?�P����'�.�R҅Ґ^��ҧ�Dr��0���?q����D\48��ʧ�?���Rc�ӝ"��L���__yƐ��?���?�zxh��π FIa�O	~<�`Z�f�6W�.�y��'��	�<@��I����IΟp�byҏ�	O�8�˱� W�f��aJE�< �'���;��Oq��"�
M��,S�ٓ:  ���'�5�4�'���'"�O���Ο,��a�:Q�d,S�}CT�1�Z�*n��	,8Z�	�lR�S�O��(N&�����N�ES^,������B�'�b�'l�$ۑY�$��ԟ��I�<�$`�s�\Ԋ!�ɑr�I[oJT�p�4��J>���?��+�n��KX%/Y��n���Y��?QQ�B�����O��d�O~�O�ȓA�˱ wh ؐS�N׮]b_����P&�$�	T(���O��D�OR�4��=aV�߸VD�� HP�� ��;(�'���	ğX��Hyb�'���J��� �	_�5LH��6�΄!%*�f�'��'��'�副w��4��'>g��KaK��E
0�㓀 ��՗'u��' B_���	ӟ�b��P��Pks�	b��"��W�j�,A�s��ԟ���sy��#X��f�AD�E�E��y$��W;)I��O��d�OZʓ�?q���4e����)K3��왲-��z,Ic�拻E���'��Q�t �����ħ�?��w����V#�=�"%q%F�a�@X1�����O��DZ=���*��t�Y��E��V������9KY��!&.�O6�~�\	B�i����S���$���$���&�vzA��̧e��'n�iI��b����O���>=��*/ƥ8(��0��(���!(~ �	ß(��쟬�SpyʟT�(�o�+{x(u���C@Q��,�OD�BsiW8-h1O?MJ! �U��!	A�Z�$�6I���؟���ԟ����p�l�����/?Q�叽��˶�f��ڠԧ:� c�����X���?��'�*�1Sʖ2���SRj5G>���?A��Ż��$�|J�r���LRt ��
]��l`�e��5�	y��eDn"�؟��'2$&*A�d�+vr@$oɺSz�qR�0�	��H�?����?qfg�>u�Y�����yB��z�b<4g����@z~��'R"�'���[>�"��mb v+��M8�H䉓W.б�'�r�'`�R�0��џP wj���L���>&�LiaT͒���)���_y��'$bP���ɝl0K�|*��{k�p3��ׯ����E^�.�y�����'b�' ����T��0sY�B��8������8��D�O��d�<a�e��A��O�4�P8r���x���Ԅ]��]Xa�'�������	�[�'6������; V�Q��@x�\3V�ʪpET��	}y���,�7�|Z��^�\���^+\�!L� ?ʈ7��O����O$�2 �O����|��#P����G��r���H#�¨�?ɳ��=w�6�'h�'��d�.�4��E���ή}�����o��Ԕ+�6�&B��s`b�'K"�'t��T>��<y%�4L���HIA1&���d� �M���?	��\XP���'�?���?���?ɀ�Ψ{01ڒ�߄G$P{�@�?II>�u�Q��?���?����?��VيХ��tp�BZlZ	0���O2���/�`%n���	ğp�	����p���Ш��`�҅���1�<�q!��<y�fS�<����?����?�����)��,�P��I*���a�I�77*�i���������L��� ����ʓ�?���*7hj�:��-V�8*%g4�4��?i��?���?	,�"�""Ħ�A�$��wzr��k�2\����5���P�����러��zy��'m��a�O� ���Bjm��q�T�H� ��[�P�����I�d�I�O\�1ݴ�?���(�xa�1C2T��C�ʱOp�y���?����?+O����/u����~�[u�J��h	�#�n��׍_��h�	�����ϟೇ�Z��M#���?��Ӳ^w]�%�Pj �U�g��J���KP�'��_�h�	*!��������I���:5�N����Y'b���Í�#A9��Iٟp�I?^;��	�4�?i��?I�'����MGV	`�댴3��Ԛ2�50mJ��.O��
����$�OZ�$�GJ�),���«M\Vѓ�.S�X|���V��������Ԗ�M[��?����'�?Q��?��I�x�9`,E
X���J*�?q�o��?�����4������ڽhͦ)�Nߖ,���Vb��8I��o�����ן��f��?��	��X������	>usԥ�v���@M�JDNF.t���I{�M���'?a��ПP�	�P{d�ҡe�2`jRp���TpR����xB����MC���?Q���?��]?�ϓ!ʨ��ڞ#�mЌ�t�'�:���'1��' R�'S>��R0����SU��X��ǷSB	�ش�?����?��)��@y��'����R�Xh��7n$�0c�]��yr�'���'�B�'��P��xq�4O�ب�׆̓.J���hc�1�R�'T��'!��'��� {Qij>�D)�3�*�XT͟�ly ���#���I����	��4��� "�1�Mc���?���ǋQ�H�¯�(Ϟ�e��0�?���?�����d�O��`<���D�Ox�)@f��I�@��;�Xl�2M�&}�����O8���O�H�Pi�Ȧ��	ş����?-YqQ$��(�6TS^�������?������O�8��<���tD��ϧH�(���Cu
��nV�r1�H���?Y��_'�̉ �i!"�'���O���'� 6�͎6�.�&���R��CP��	+v� �I��ȗ����?ejC�[�$d�K�d[�Lv�DS#�O�Er��H�����؟��	�?��S��P�I���+��B�6�0;��-*`�a�L���h"cN����Zy�O��O��� �q���#U��\���+(:�eB~Ӥ���O�Č�.��i�O���O�$�O���t�K.w��#� ���h��O��$�OL�� ^!*:�������O<��˫Rw�D#B��pG��9��1:�.��O� 3�$�ަ%�I؟��ʟ�ث�<牃mo.:Pl�p�|�����˓sD��Γ����O��D�O���OF���"պv��$���+B�.�@�!
,$��oZџ���ǟ��I���<��i��Z�M�ZU�e�`����zã�<�-O����O����O.�d�0��l�"*�.YJ��+�� �`�4k����	؟��Iȟ�	؟|�' r�����)Pr��ġq��1�N� K�>["�'�b�'��U>����M���?Y�	�S^�l`Bo�<6����G��?1��?������O�,0!"�<��'P��%�~_�ʅ̑�u�z���?���?Q��H$�#�i��'�b�O�^�ebݬ@*1��i	�|�4�@&�''R]���� m�N�u�i>�q�����4[4��B��=��Eӟ��'_��wcz�����O��d៞A�'���SQɃ�h�����ǆ�n�Qv�'��'f*���'a�s���|B7��/����)��!#��	؟T����)�M���?Y�������?����?A3ㇺu�ܱH���X��ύ$�?9�K��?9H>�'��'�?)5g��IjjX�VL�����#Әlp���'���'�p�i�O�B�'�'1�
ԞzA�EP㭊 E��-�5�OB�|��]@�O�B�'$d�,	�|�poڹ8CȔӄ�FYd��'�6 ���l���D�O��D�OV��Om󄝲hH�)��N]�U�]�e�3d�		O0�	埔�Iӟ�����T�'��`V,00������1��{E#1a=TO���OX�O���O�-�C ��~
0hqmVD:�D�5�G.��<A���?)���$�,M�9���3�ިj&�ڭn��5�$�N�Om@��?������?���>�PP	��6sZ`[gJ��T�N�$�,0]�!(OX���O����<��F��<a�O�<��%)�d.p�&*զY�X�2�'�R�|"�'���T�V�����c`�Ŗ8#z"�CDl��C���O(�D�O&˓~J�a3���D�'i���<��{�R�~�DCf �[�'�r�':}Q��'8ɧ��̈́�nF��w/4Z�.aC�9�?�.O����d�����O��O3�0�,�6%${t����>%3�5��ҟ���2c2��	s�)�/'f �{Gn^|"��T!P�2���$��hl� �	ӟ��S����?!�
�ee��c%L1�<\1&����?�2�İ�?K>E���'��Dx�O��p��0;�d�gVZ��l�T���O��^1H�%�4�I��̓P�i��ƛ|�^P����7�����G�ɢRBr�$?I�I韘�Ɇ"4M�m�N;�:��Ƭ�O����v�&�H�I韬$�L����c�v�`m�"b��aVqy[�4bR���Iϟ��Iy�*��$��ծ�fiz�`�(�4�҄/�$�O|��+��O~�D�Z�cd �#@q���6�r�T5O6��?����?�,O�A�,��?������5e�zD�U�d鼵�&�<9���?qN>1��?��κ�?	!���J>��I�*^�bp��N�����O�D�O�˓&@(�k1��4)Cs���i""��>��3��E*h��'2�'��'B. ��'��ə#�d��ੑ�sQ�����+^wP�D�O@�D�<I'
$-a�O��5�p���k��n@�-27��6&l
������O]9�.�OڒO��31Ą$ ��1|Ѹ "vT�`R\�@��Fٯ�M�)�&�������'�r�����Mf֍�3�N�wM6��(O4��X���d$��e�R�T�*��Kn�5횝���'@�<���'���'��OL��'��S�2M� b��|76IJrKų}b���'� #����O���4&�$����u��~V^�J\����Iݟ���6U^���O�ʧ�?I���V�9I=*�B���F�"�����3�d�O��d�O�a*T�2r�QY2A��R�@��G��OD�Ğ�V��$�O6˧�?AN>G��l䰱ӧ�� �����z��kqRU'��ӷ,@ jt^I[�[}�tKv�[�\}�T�&�G���]AE�4V�I)����`KN��PH�?y���?�����V{�)!��5J�U�7oG:�Y����?����?����������Z�E�~$����GF�� p�t��џ�IП��	U��ޟ�+2�͉pm��ࡋK��܊l�#D���6+ɏ=J�d��-� )�+�/����ӨAd���	W."lO�1�׵0��a��7��q+��R�p��	�qbҫc�~T�j�8V��v�=~Z'kE�+���kC�W�d�fi�gٽOƛژY�n��'d�6��''S��X���k:
eP�����gFZ��%E����-p�f�9'� =����-38 <U" �̿-���hfj����X2��Ɏ(�y�Iɟ`�'�@P	B�-�,9a��-;���F��
tc�X-F��|�'�i��l�1��Z�' �e��8m�Xu����>J�6��(���M�����؄����/��a��M�'������@ʛ꾟�ɳퟐihD �D�E��\L��,���P��:($8�� �T.|�B`���Qd��<9��4�^m�d�Τl����ܗ]�h�����3���d�<A���33��D�O~�F�i"2�)���+�`����!�)* "�O��/l�<�c��j�Haҟʧ��i�$O�Q�fgA�n�����˔(��'��%0v-��6��(�b�$���	��`Բ�B��0>@� FTq�A�&f�~��f)�4�N�!��L~ҭR�?����h�`6��qJ4��i�0h\x����L'!��G'%P��T�C�Q$@�ЈFE
�x2�,�"pj��E��$����RL�F$P"��>A��?�u�:���"���?���?���\�UjG�ҿ�2�p��88~�麖�6F�����	lӖ,��!*M�1��'�*�[p%�� ��0Zs+[��4u��LߥpA�:�MkÄ�<Y>���'��.E�u�6ذ�-��+���j6��O6�lT&��i>�Dz"$N�P������̀����y�'/�؄A�����T��g����ɢ�HO��z}2@7MZ�؊G�ޏ{��1�'�@3��y1!�=?��d�O����O�ج��?Y������Q>2���`�85�0�ɒ�F�`�,X�$xm��Z�+�i���$ &2�~y����.�|��Ab�*H�㊗�h'
�3 �T	).�vN�&\A��@�Mc�AS�)?�6�N�r��"��'le;��1+>���	�@E{b�d��dkڕ��"N�]���KQ��N�!��I��D�����$\���L�Y^qOИ�'T剧=a��1�O�6�T�k�lH�T��%���1�Dˬ0YJ�����P���ٟ��I�|�ܖB��% �F�1 5�-���5]ۚ;>y��� �;Y9����J��\(Ӌ|��Uɐ��6f5�\2���!Y��qSD��tu�� U#F�QH�����	�xz8���O��L0����OFm��Ň�&��@�=�
ۓ�\����*R�i�ReY$q��Gyr�i>� 
N�\TZ J��0.� ��W4x�4�Icyr��3K��7m�O��D�|�OL��M�1%N>5���(v�B�@'�м^��'Ǟԩ��Z P��y��c�%��T>��O�LJ��M�O�p�HǂG����O<�)I�2P�B�԰qf�iD�����z�4�)�*FY����d���ē�y�ɬ�Mk���d���'��0��2f�� �L���'vb�'*z$�A�x������%}��	�y�Q�T���ԯi���A�jIB̕�!��c�4�?���?ᢋD�R����?���?Q_c�HX ��V�@� �O�\ٚ@��i��#��]3GN:   k�k��_�Jb>٦Ob��BҬ4(��#ͨ����˱9����SkF�R6������(�'���Krj!:{hI��kF*Oh�R�i��)�	��X�	������Iޟ������z�kB�e�d��K�2[>��%+�/Ɛx��Z�"i�{��ʡeɺ@�#�ȋ��I*�HO�xnןX�'x�a�FG�E `����6�D�Ɇ���t�22F��O���O���ͺ����?q�O�m�Ԍ�H���%�R���lk�*	�M��P���Wh��	�C/�+�N�y���n�'��(�DLْ�`�' ӯNA�*�	B�B������I"�AS��0v���"_�%Dy"kݛg$����QY��Yc"�]�&��A�����{Ӟ���<Y����'�,8���#����Qdה:qy���T�8���TE��4� i6X�i�=�CB���?,OP���CMɺ����M��m;F�F�CU�C�Z�����]��'�Լ�5�'|�?��PJv���o��$�!��|�>`z��N9-f��%��x1b"�GZ6�?@ߍ+l �Dl 4�ո��Y9Y[K���%ہ@R>68�$A���w�'�|��Q���'��6�%$`@��$݊��kr���v#����O����O4��/��,��6��,���\�p4:�PAm��.���D�A��%�󏇼2Հ,��˅�Z�R��1��O\�OZ�n����^yRcK-KۛF�2b^�X���3���*�$Z�D�t���O�5B2�W6`:��O��gy2dɃA�kvX�	���""O���ēN{�i��P�b��C �P���ڍ���R#�E �%�T�8�VF���M�X�	8�M���i����ĸ�s�&�g:�1z�O�	rˤ�A�Ic���k�8��R��2A�y#�n��І㉲��Ľ<yܴ2e�a���,��*w�:?�R0�O4ʓ�<�� ؇v��1�2#��0�xxۗ�3T��{R��d:L�u�]MJZD�pm�= ��,0v@�]h��TD�Gx�Aƈ�P~	!"�N�L��� 4D��I�mޜ(׶�зȸ1������(D�\:��E�N9�́(��)�E5D��9Q�ؽCۀ��%�PX
C�!D��{�ہf $�	�̖'>��bn>D��٬)��|rb�ɉ�|I�N<D�p�R��6̌0g�I7!�!� 8D�p��̒ ��q�ǴCި��g�2D���@ WJ�UReN=}��r�m2D���� !�����`�3�~qa �5D�[�ș�j'�p�["  )B�^�!�D;'�����Fr�t���j/S�!�� xmYT��;�v�C����I{�"O���6��},��sG�Y���t"O���3��A����T���"O
��̶r�6���K��c�|�{A"O:���Jvv���D�T.ϐ�	�"OX�PE�1 ��X�kQ7U�}f"O��3R
��B��P��MH"{����&"OH��,�ve�J�,%V�,��"O�4듩�r{B C��	����e"Ot
&��._�ny�����[�(�sC"O2P0ӢE��t $��o�X�K�"O��!$�+���«>%���"O�xyd �V M؁c�89�؂"OR�B�$݈Tc��^<dY��"O�X��)�^�dH��Ђ,�i�a"O���e�=kI0 �Do�)�d|r�"O���D��d8d��3�X�1"OZ�1c�Y�O�0HD�% �K���yr	�&F2I�s�ׂh�f����y�F�l��!�M�6T��9��G��y�i^��
��I1��1�/���y"�&_��}�2��<K�p0���չ�yҦ�SB��.KP8h�.��y2l�4!�>ѻ�n�(dbx��ʑ��y���n���H�'�굡�F�%�y���:%�ň�Pv�u@GC��yR ��_"jtI�̎��MCe�)�y��?E\M��n��n]@B(�8�y�S:|,��)��	�5!��E��y�ˇ��$4s���Ȟ' k2��'���Aޜ
� %a������3�'.��S	Ƹ�Gϟi��
�'Y�%�b
�E%Ċѫ Yz���ic8,�g%��.��p��i�<��x��IN��xHT��+(^�H�C�4>��Q�ݪW�l݅iX�P&�E�*���i�4X�0�	'��KoC�+~1���+@.J`�R�D��G�p81�"O��8�(�
W���ԥ	#"�܈�F6Opd��-MZ�(
��<E��Z�N�8�3�m�=��T ��D=�yQ�Zk���el�
%���`B;]C�	�-0�@�G���|�g�'i���l�2�Ȝb��V�}<v��	��X�(���(n)�D�Z�oG�Ȩr�j�N@�" ֳ��?�s@E�)	|ˢ�Ʌup�0т�d�'u����hU� ����t��`Gh��#K�2�Xy����y���"�QʰF���ܙ�
���y�OѤ	g�(	С��)�'!� �mUtiP��p�P�}M��� �ʹ�1φ�_��yCҨӷ�j7^��B�Ϛ�C����6� FxB��*UP=�5� �(�Y����0?�@�R�XX��&��BH���_u`�h!�Oۖo(���Y�n9�O�G�Ɓ�`NM�`W�8E}r��s�^iX)\X�'�&�b��1f�tT���+u����ȓ}G���#HV'����Sm@.y�6ʓY�����5��S�O���V�X,J��h�ӏڕ�h4@�'�x�s�7Tr���ȏ�1���'j�a�o۹s AٕO0M� ���'��a��F��(!�})��ãF�p���'D�"��� fwt��+݊l��k�X�Rp#���4�¦x��A�O�B.��b�,D����47�W"��_��l�M)���LZ�=��KD�O6؉�Ď��a�n���b���V�x�'��`�LL#E��4P�Y"i,���9�� B�>6�>A�,X$p~d� ��1��!�0��V�<���K�TxԈȚ@[�c�ۦui�
����ys�'��C��MrT8c�j�"i�`E[I<y�fU�DФ������z���	�4����M�5��� �T@���!}�nMy��̼~א��"O���@�_`��xzդ�>8!0y�Vd�P�Q(Fj���BS$oN����?�'�D�M҂�]�4��Hs!�4Jd�%��C�L�pB�	�5���
�e7!�F�r��_�)�FdTg�,vQ�TS��$����'w�2ץL6 �J��?9w�޿+٨�Z��\<Q�x`G�t�'��t��*Еv�H%s`��Y��M��/��E~h�ۆ��O⌱x�a6Ǜ�H��v���S��q���9�I���0��ۄWB��>!F� t�>�rr@ O��,�n���r��B�"
����0rq`��u�^��V恾(���"O^�@2�͚6wl8�Ks�6@�a�'���	�'��s�(�a7�yT�P"Y?��i>���w̶�[���"�6ŉJCZ� l
��,F�E�wJ�!�vmk�����2�sH2� ��������g���~bE�_��)DyR.��x�]
N	0cX��.��O �3�h�+v@�9���O�r�H�B<_�铓��1*�ޅ�$xp!�@"O,�[7eωf� �c��v[j�¥7O��x&��>���R���^|"�cW�O	�(����%�qq =�"�qo�D��"O "5P#P�����X�dB��O S7
!"UK�!<J���$�>��S�XHc�X�D�B�s�)�v�×t�	'�:�O\�)P�ܹiS:͒�lSJ�n1� ��*K��Dn	�k�:��4�V��	���'1�=�3K�'�Pmk���;������D�phC��
J������9+��1�n9q6��C�Q�K!!�M��ZE����0"��2�'ީ��0��,��|X6d_��s��#���\��A�ݬ�ik�6D���H9���x���)P}Hr	�O�ذÍ^sB�i�╆&���$P	#z�x2�9]����	��{��C�2�ұAq�4|z��:FE<�H�%�E�%H^&E�J6�(�O�T�`Cޚd:Q`�Ȓ*��&��|ڦ�;����FS�4�F�~:SI����V�߇O�L��5�H^�<�4.R�UՌ�+q�A�P��g^�L�,u�mI:��@�a���{���O^}���K52���T��hMV�B�"Oʥ:TOf�:�#uN�CH���%�i��!�l�y��=�h��`���03��īS,D��-�bI<	{����"N&��� �X58ۧcG6K������B�	�*�09t6�"�O��Iөп<�~0�k�t,@ؗ�
�|��3��#{q\�@0v���O�N�b�aܑ3 �e"��
*	����'3����0���A���>+*\��#O:|���a������ɹ툟�dA�sU��X��D�s�;��\�y2��)"=�B
�	X�	{Ed���y�b3(�4��@E^1UG"��I�7U�x	1�J�%�
��4����<k`\����7fL�CT"92X���B),rX|�cA&$�����	�b��装lI[��ͻ��/�\z���G�K3~{��?i*sP-�������h��)�0D�\3�c<elTQ$$�u�H��k�p$��LA)���N�"~nZ�
�,��#l�&<��䙲 ��B�	#H`��0�W�H K4ω�P3Hʓ0<T�ѬQ��0=�j�OU���5,�^�dK oX�� �I-Q� ps��(?�qbd�H9����R-8D�TBXJ^M�v�	)2;�Y�mY8+Q!���L�y�'�y��H���d�!�D��.��K���,�*��ިf�!���" ����&yj�5��N�!�̬C��؃���A�̃��[k!�D$o�z��ԩ!;B	�3#�5f!��F9uʹ8j��9FFh�3(ڥ`!�$ƢWkV�{�+	,�P=����}p!���(�y�"Y:B��� ��~t!��<i��`��B��8��e�Y�<S!��
KhH�"�,Bl�Ը���0!�dP?x���S"ٚo�����K !. �飗x A@Xb?O��� ��-}U�aw�5�M�
O�i��'�<�r A�%Tt嘶DZ.��Xr	2.�}�$�s����G�'�tH�m��p<arO�h������tyB�J�&i�݈���fȄ���J��y�懼P��0� �W�gF\91�g�����.+Ē�"���zLԢz�`#:0��G�6��3��V�<� ��*v����lk�)�R��y��c��g���+�����%&�3��N_��U���.��Ip�!.,"����.\�v)��͚&���c%���0p!�+�İA�'&Љ �`[Jo�,�#�	a"��	˓;���a��Ԩ��� �4�`US�H�1&Mc�C�	t,���")W�-߮�2�M�R}$�O��#�MS1Oq�f���T�D\X���Rv��$"O28K��<SI@x��' Ft&8"O<{�$�B��mڗ�LdL 1�"O����F��up�8�*��PXbQ r"O6��$J���y�gI�H"�i�"O���w�5�
��vLA�F�@���"O"`1ӏ�
"� ����8�n��"O���k�&~re*
��,x�"OL�h�B�&{-tqp��˽D_�( �"O�U�t�&x��بG��pL�=#�"O��Ǌ��A(���sYR��"O<yp�$>Ct�c��5_�p�Cb"O��@�G�N�l@�c�ޙ1��p
�"Ox��4�<A�Έ�׮_�J&��["Ot��D�[;&�4�Mڟ:*����"O�@�`
��&A�Y97�x���ˌ&�y�ؒEh�#i�|��&N�A	�H�ȓF�������bvJp�e(ԉRx �ȓ$?V��w P��:a�aЮ
����uRz!���)r\YY�N�Ե��c���{�-\S$�a��O
�%�ȓ{�8KZ9L�M���.QL�r�"O�k���d�ZFhV/C>AJP"O����Ɖ����b�>K��!�"O���!T< ~�A�הD�ġB"O�� �Q�B�p[��W�(�X�"O>�A��'e}�S�'�-M�N\@�"O�uص�.&�X$i���4�f8I�"O>ى����u�S(2E�m�N	��!�2)$CU+���B�ҥo=!�ߟ]������E�� q�Ȃ9�PyFÒ1���C�'�(�$�c�G�y�Hї`h�� A_(Ρ#��C"�y2'B�F�4��@-�RZP1)s���y¥�	P7.!*$�)T�\8��Eȴ�y��X�H���a��TѦ��D��yr����8u�2fJ/@��*����y��¹fm�����:�Ԡ��ϗ�y��<x�� Z�E&d����k���yBi�+W"V)�v�j�*����J7�y(D�	:�ݑ��׏XR�1zp	��y�	�"R-�yX�.�<e���ф��y�eEd±�ҦD�Հ-�s�T��y�P�p�E��!�{G��b"�U+�y�)�;���I�(��r�l���H?�yb��5WkN٨恼m�*=�%-^��y��d�hrVo5e�N���yb	6)�V<��i���FX��yB
F�nC@u�q�˨w�j�t�B3�yrEL��p�p&i=4QF$�fQ�JX�(���`���;ㅅ!Fd�y��_��qvjˠ&��4 �y���]c��K6XMz��҈+=�B�	�eJ�|qU�6C�n�q��d,�B�	9M��I��H�X`L��B�tB�I�B:��v�Y���AMJ4wC�I�H�ڔRbA�WJ\����<�,B�	�ZBP%pFNՀ{ �R��E�hFC�Is�^��R��"ϰ�6l��|C�)� RQ�
]�)�,�Bm���>0��"O ��ǆ��1��`J�I�ߺ<�F"OV�;���p�(��A��� �<X� "O�=�T-^�@��80�GX$�,0[v"O��3%���E���KuF�:/��X{�"OX�!E.��W�I�"ŕ*cK����"Ox���Ƥ;��3�-��`�LM��"O��Zf��
{���)�c��o�)"ODiI�Q�i�XQ��	�i�(2"O�4Y �/]��x3�MxH�"O��`N�m�֘�����l#"OYC���a@i��	�<�"Պ�"OeC���wr��J��D�s�Lq"O~eȂg�0gȴh&��9@���&"O��Qac !��u�a�#I&D��"O���N�`8���+U�G���2"O$�i�?��9x�� e�a�"Of cAO��f�hP ۧO�1�"O���X�b��@������"O>m"GBݒcު��g��&bR�\�'�ɇdH�E��\*2g�@"����}���q�]"n�ʤ w�'�>u{�Nɯ  ��R).JN�*��7n���2�i>�$��
�'�	�RD�6٤IyB��
bI��'�6a#��֏q�
=�A�!O��1.OƬ(��'<hA�{"��B�$y�1b��W#,&�@��֫*�p���ƋjjpH�ݴ/T�,��!�$l}|�� �� )8P��F�D�4\(h�?�'^p<�Y1]��:�ƕ�"�,:���7\ϼ!c���pɜ� fHB�T縀�p!�=�Ha���,��?飈I�et֘�oϩ+�d�G�����[Bo��@|qO��'�N\#K<m��[�� ���!�Nؘ&l|�<9T��-YҤ��d��4��tx��y�΂��?)��Yd�$�2���	C�cg���󣗻5]� ���'ݺ!��f���)_�EL�s�vL<�s$ʸ'��;���>1IRx�*�ٶ��w���5��N�'4&��e ��Xp�T�������L)�X��ބL�rݸP�
�
����T�q��ɣ+8<��0�/y��Aq3��NF=����L�H�#�6�~2���D�h�Ft2��O<$PҭͲfr`ja�ܳ/�H���-D��Zr�&��5Is
-)�\�c��e��'�L�C�'G`� K�t' А�'<��F.G�YH � �BAӿ*��{R	�4�4����V�
�����=�F�´��d⌠�G���<�weN J"Ƹ<!��|�
�F.��	ch�@h�����J���Ia�k��w�L�r��>] �sc�mD�OTeRhۥ$�dC�䏯k����I�<!��|�X�-�IFx����
����%:(3&��~Y̂�����Њժ�#�μ'���U�s���w�DФ'�3�I�RT$)�'����E�_r�Dr5F����Q	RMƩK~T`8ע]��'vD@x�'c��j���\|�����"��X�t��5�4� %���0=�ǆ�:4�p�^c�Ĥ�FH�$b6V�"s����CVa��I�Mc�O41+0a�4A�2da7�~,�I! ��	��<[��G�6^�0�P���Oj\�G�8a�>({2���B��c@�>�eF@�.!h�I�u��x���h~R��gb��Qp��;�	�Q��D�0�I9AO�I1\~ZQ*��:<������p(J���2�Ь���2(�*
���_d �$������&b0 A"�N�UZXxC *S�N�h  `r�!��@*"�����	?aka����N��06l�#,Þ���i̴�I(g˖���?����%�p� w�פL�b���[���E/4�����'��-c�gLq�$�PGH�MXL2���v��5�CR(5�I�s���YSD�M)�N�0�XM0Zwr,E*��Z/W�~H�l��y��� ��D��%6X����/)���4GKz*a2:�6\�A*kg�ԑ�`����K�@xy��f?ه�������D�݂�8��9 %�Jc�����CȜ�C�r9�Q��3�#� x��Y�����ʗ��ot8C�#[/i�TES��<I8]�F�4�����BEe�*��W�'�,�ą<gq��V�@�
L)��ђ{���$�6��Dgr%7O�b>������P�-�Fk�&�F�	R�y;��A����O�i! �y�K��v��rf�@�]90����M��
����@�xJ|���O|�Խ�(�����:�&��E�ON ���	i�)�����z&��A�+� ��O�4��%F<�
��*(A$�[S�|��
h�$�Y���4�$�P�����M��蘍O��0��-L�P�:\�f��h
���`�#)_¥��ӵ+������?��=� ��¬�KʚL�'(n���	�Q��?����_�r��2�� ]�ĤQ�'=��(ƨ�;A\�q���zp���ӋO�"�8��'�Z!��S�'6ҁ��IF.;�L��Plcg((L�e�I��H@�5�����8(���v�R�Y�M��<�&����I0-ļuf��OF�q!j��o��9�`�X?g�^�;`DF�WlY�ɕ�9����H�"}� ��?7�VSS�Pj5��&^���Ƈ&'ў�n��i�(�DJ3o����K�6j7MD�v��zw���$��-q�k���D�h3���7��J��2g9��ԟ�O�i��Fx�H�g&H�Be"�I�_[���?�b�%DbМ���m����HEz�ŗ,~����G�pc�i���A���(��O��x�I�2C2�kӯ��h����X�L�+7,S�v}*�F|���1my�u Äɼ�CN�y���b �$|�l� "G~�HLxbY���<��>2��E��e�$_�xٓD��E��@�$1��D
�c� ��oK&���Îjh�O��ж�QK�~��D�×)���is���L�*�ZR���a�-v�T��(�]���-Y䌹ta�<C)�4� ���A��\ҖM޸���1�JZ�H�*��<qJ[�L�:�YK������� 10�ʭ`�`����QȘ�9�n�Ԯ#l������s�"m S�z�d�)b(�J�ZH�<i�(�N�Jhz')�Dy�_>�]�q�nQ����m�P5"�D4x �C�1ȣ>��E2�@E�#b��`s�S�j�j�hS��iX-r�*���Hy�i��T���i%�����86�����G�(xz7��%�'�<�T��u�����@�4��90K>ɤ'�W�ժ�M�'l;�s��\�r�@9Y�z����t~"/�S����UM�(��q��L�<���^0�
)��e��vZ�H�DVNN�1���[�v�hc���Ę'�f�(㩄�@Dtt���F�Y�J� 	��s��| ,�,��ɛ�'`�:�dާ @�� ����9 JG|R��0�^��cc���Fh�V��j51OVH�֬�n=@�H3�/v7m�|λo�,8�IÔg�R�)Ro�Q����٢4MG}�"U�bu���&���*T]΅	B!�b�\��/�.�U�]�$T��(Իi�꥓�O(�O�ꤑa�!��8��Sl�F�pwA�F��0a�{"������Թ�a�1�����]�)��^��fe��"N���Aɘ�dw�e�%oWuΰ� ��O�Jr�o��숦�	S�u0�'*�٨���lfF��jRH�f<i�*��J1ș�bn�:1/&��`�d�85'6���gױB�"ث�*Oq>�Q�+_,�b���rDM� Z�G�"	���$�	�x�^W���!Q}��-0V p�<�R-4^�P�U�Q%�)Aا�ħ@���*�I89}�uɢIX����
��_�r��E}�M�l�ě���e��(u�l�ɐaĺ!BE%P�lc����_�,y0�D�P\�#|B �[�Va�t��%t"q���R��&�S��Lb�Y�#��-���茑���	FbJ! ��};�=�F�Сz�<�!&���ڵ�ңH��'�;"�� � ��.<�@���<A򌊇r��h# Ǘ�se2]��L�5dO�y*3�B�|H:S.å���O�����T�k����%o�u׮�-K��J	�E満�ŏY�Q���Ӷl.K.�!X`�(|�t��d(5�4S �-+��c��$C��z�V-+G�*B	� ��FJ����a�p�S�OS���C2{�X��#��C}N��0m� J�T�>��+��I8��d���!���c�1"#m�
]�\��Mō;�H�;��Rƭ�֍٧?�D�'䤌Ze�'����uK�3#�	J`)�MV�K`!�|��=4��>��F@"!xm0�JNҟ�'Lb,��S�y�`�	Ϳz#$�AA,�,l�e�D	F�P��5�'Dr��K����c�Տ�$��{36���:D���h��6O�\t�3k�.��A��_�>^`��S��O�`���M���2HC:juq�ŋݿ�\p �H�yRo<��yT�'p@�e�4@SZ�'����Fd�5K5��@f؝wÀD��g��-ĦX�Pk,$F����;�l#0�r>7���͉5(P2� Z!%/f9�0F���R�*3��x�`�8a(:!�;����Uk���H��a�]�0a�ųi1��%�A�d|���)F���d�p�4���$F�i�t,H8]"\ac��ˣĢ<y�I��dƊh�p$X�\`a��~Z�_�U�R��bhX�i�y�u��֦��2O�'W��ӏT��]�)-x�q>���ΫO�BLr3�̺?k�x+���*|�� &�w�έ�����R_��Ѝ�������O�h黗bU,A9CW�E7x�v@!5����?I�4%Zu�C`4#�3ʓ
i6EPf-R: �|K��9q�$���nC$eV"�tfڗ`,�3G��|R�����J�8EN�gt���,f�J�S�����x2$�6L2���;*��}R����b�P|Yf蛐�ڜ��c�e��*� շ%�[���I��O�Ӈ=E�IP�%YYLE����T�<��Gէ}��HR�-:�LD���!b1l�vr-
��	?�. �&VK����/ǂZX�',�m�7ï?����B  �J`�Q��hk���my�z��	1 �"��6��ے/߁'J���`�)N�G��� �B�N�9�dms��ТpYЭ�d��<�C�'<,�ͪq���C�F�Y�'�V|��ʒ�;���C�O��w$�L��d�7i�,(���T��:��>Q�����:!6a�DM� p�	 �Z�w���j�16��xR,��+�ޤ�;�DACC4N��P��J��%Z�cq_�p Q��O�=jQ>�.D9yԪRD@I��3$� �#Q.�<br`S��BR�'N.%K��Dt �!U&�"�raQ��_�1�WeǶ4�`Xj��/T�0�aFO&;]fL��x���v�͚,��5�������[뚥2c��C����m� {۬����I
s�:ܣ5LL,N]	��Ŋ��O6��E��>�4����yʀ�cS�^4��A�A�i{.���q��mħ� ���P�  �T�P��x�` �P}�!���3x��l)R
�?|Κ����v��8�CEݶb%���$� ^��\@WGس|�d��bG�~�R��D	�>xR�a�M�P\[�狏��ݸ��қHn���I�+��}�H[7�Px�}�<�� L�e��1!M� 0(rt	��0�G��+�DGfĢ( U�n�̓N�0�n��
�H����)*#�)�	+3n����
萜�6
��B�N�>i���ID�e��� �C
ԸT�<�@�K�2�P����h ��^�';�����z����P"M�~�82�+*Q�����I⦁�Ɓ>n��eҞd�
}��O���4�'>T��7�z�b�G��7F\;�_�THF�	�:rd��5�ʩX��@6�ذp�n���˅�-j����ʁ@�B!�L��hO��p�k������v(��ň,!�O�euBрEgts%�o^��A^�z#Ù	9�Xy�%(2o��8�`Ђs����=ن��E\����'Ţs�i#dڟ�S�-[�I�R-8C�����ۂ�<�~�!��#ߔ|��*��jr�:���Y� :�E�;/����(6\O=R�oІ[�������E�����C?y�O�80&FκS�g��/�O�b8 DϣusN���ֻ{�ʸz�j�2�:���N�r.^�0�ܒN��;u��)yK�`1�j[��d�ƾ{�Ꝑ���)V;�L�6%@�H^x�[w��)�:O�L�"�7���u5zP�Ł��:hNX�`۷8�qO,�[��K<���Ջ�N�4�Cw�'S��SpǙ�^�tm�q'�K�I+�g ~AZi0N֔]���D�v?	��X�12��>�&�Ƅz#KB��1�2G?Ejvc\���%#pg�1`�)q��b?֥8�+Z0��_"��6,>���]8L86��:�ĒO(lx��'�ъ�G��M����ݮvE�$sf�'v̘$��"���hSlX'�Ј�OЮ*����N���
XB��n��fEf��'4��X�1D �4a{7�F9WTU!�w�(���7�h��tMU1P�1��S�x�(���yjuk牙/C^�)2����b��O��a�H'��ѥ�&>x��� ��I89P���7�P Pyz��.G��y�M-���kɣI������[�~"�\�L�=E�(͍?�q{,�	HVZq��/��yBk��96�P��O��������ē[^�ד.�Z��8dYXŅ�'?U^��Z2�#bZ��萣��
�F���r2���k���-���J*=��ȓZ�| �D��Iv*̓@��)��݄�[�P�aC�����Dӧմ%�ȓ���x�ʎ0G�,���
D95��U��c��+%0๷���MKh4�ȓEp|)� ˉ6Z�;q��tO�y��dO��{�FĒv�����O�מ=�ȓ4p3�"W>&��� [#mj��,�zbQ��3i 
w�	5VwL�ȓ5���k��Ĺg)���7FK���ȓm�d�1�\}�B+��̸�ȓ�a�6j����!�JY��M�ȓu4>ɀ���� j��HMLV��ȓq7B�C�M�'p�<��D+�{��@������MP%�W&���ȓZo~1ee�}4��# cM]��|�ȓ���x�oO|�RIr!�ٽ�Ή�ȓepE�
N!P�$D��M�/�l��F�\�	����,�B�V�q>��ȓXе+'�a
,M��h�b�P��� ��M৫4A(��Ҏ��.W�U�ȓd�&�:qA��j�FA �#�+�6(�ȓ45ԑ���%9�u�$��n�|��ȓE��Q"b��{������/��P���wD,��,�rmIfbOJ(!��:62<q�fo�w�����L�.!����&I6��
��J�vw.���"Oh,�TR�w�tM�VJ�S֨�X5"O*��"��s設�%��	]����"O(�q�F�.x�,╨�A��S�"O���-��eԙ3�dĽ}�xZ�"O��b�<_�441PD�kK���"O La�B��C_�Y��"H#C&	��"O� b��0c��v��0$�>|*�"�"O�Ґ�����u�'K���[�"O�03���<�4 �"�zH�"O��b�I�b�.Ac��+���"OT����C�_[�%���B���iH�"O�����M&aPh��B�Y`~l0"O8��V�\�8��uif�R>d��"Oda�� �'
���(%S<�G"OZ���+��1{�݀fH̀4Q���t"ORS+�"�L�C�DW9 ��"O��I@(@&v��l��
-����"O�D�1��M��Ր�E
;���"OvP�4�I�z��˒E %�й��"O�X�!�Wߜ�#7��|W���"O�H�s�@TbԘ	�cE(j�Va$"O�
��M5Wx1�A��&5��(�0"O�������>4
�0��(��&ښЄȓ�����^�n��{#�¢vG"������r`�%e鄨�W�?4��ȓz�Լr��?�eB�X��Pp�ȓ@�(�H�A�cӼE�!�W>hb�$��}5��+��U��P�KB;L�`�ȓ8@�Q�+.	�p���;/8$�ȓ��٪'.O�� 
εV�x��o�<�6�@)C�\[�-�-C}�1�ȓc�������dU���KH0t�ȓEt�9�G���n�t�������ȓk�ʩF��\r��ᜌ
9��ȓ93J[��X-5��X�*��Um�܄�G�T��ӯ�-Q�h� ׇ_��!�ȓ��P8m���[�&oNЄ�FG0��S8�hc$DZ�sP2��ȓg3 �FC#\�����!3&��ȓns, �֤Ԙ��z��"#x2��	0�E��A�c�B��F� `��ȓ%P���/W��\��NX���hb'[�V�b)*���B��e��.� ��T@���蹣j?k�$}��]�J�`F��~*m��#O�i���ȓ,1hi��;׾�p�h�,.�&`�ȓ�¤�a.�[e�h�A��1�$8��^���&�@�����!i�9��*%  �5�C.~��z"!ʤ|S��ȓ�´�+[�8��:��ءL�L ��V����e���>�Rd��/<�l����AH��^"I��-�A����5�ȓ�FD�#R�nD�PR󰩄ȓ0��̢2�Ԧ-dYѓ�ԔZZ��Ӓ�睭!��AE�Ɓ�r,(�5D�D{fF�kH�� `÷pp�Q�%D�H����~��c0C%!"D�� 6 I�2���'b��lx�t��;D������<A,9+�j�=P��UF6D�,�w�p�"Z5����6D����J��)�(H�%��@D��,�HC�ɀy����k^&3R�uه��C�ɖ*e�,�u���A�z��B$6C�%Y�2��.UU�	�ϔ/.!�C�ɨ�8���˿;P*)��"u��B�I��Z�q��Y,�H���'s��B�	�d���j�%ǣ��)QrԽ8'
B䉒n�X)����+[�`�τy{�C�I�?ܻ�Q5>6�-2�)L�C�IoC���P�nP�M � A?e�pC�)� 6M��	��dm��v��9�N�e"OV``5���<B1��I��B�"OZE8T��!\��0P�� �`v"O^���͊0fYF��q�Jk^2�)5"O��"Fψ:J��Y�H�?QF$}�"O�=r��<`���d�(-���"O�D����5��:�����4�QT"O�킔@�/ǐ��aŗ�"��8c�"O�z���7a�`UkW�.Hnh�K�"O�-Y�k��{��ꦁ��CZa�g"O6 �Y��8�C�����z�GO��y"$��1��4i��%ڴ`�V"ǳ�y"�ȺC����D�L(�+Aዮ�y2�K�}~�S�@�;x��m"@+W��y�����h�0v�$H�&چ�yRNg�y���L�W��9�����y�l�(8�JQ�c��~H�� f ]��y���������y��!�`IȺ�y�%��!��,	���&~'�lە��y�L �
�f�3�� <o=	�d���y���hEp|�G����T�Ƥ�y�J�9y֥��n�$��K���y2 K�����A���:���� ۾�yr&��L��-��TAկ\��y�ʖ�8*oʖ��[W�U��y��#3���;'W�FP	RBO�/�yBG�]Q����Ok��t*��yBg[5�����H�ʬR$�Y"�y�a�=9�����'�:5pP0�'�y��W	=�ٸ@�´~�:��ӈ�8�y2�΄z2�Pbu�&b�"\��,�yBE�L����!գ������yB�,G� ���q״��E�Χ�yR,A�;"T;��K>l���)��J-�y��V� A�L9碖q���(�aܹ�y2㞝j\�����C�g1R!c�����d'�S�O�8���.�R��߽0Q���'��A���U6ά�Z�S-IV�s�'W�\�f
V7P+�e���U��n��	�'��uJJ�)O�zԪ�" �&���'.���LQD�Q���s�'	e��!J����Ӆ\	­��'�����J,bvh��� � �N$��'|F�2�G�?&)Pt�xMt�S�'�"�I�+\N�]z@CQ�j��P�	�'�0 If$��˜���״^�����''|�yo�hi� � �K| ,��'�졔 M�j0��	��T�D�$�'�ԭ�>j��ܚ�nU�.�X�
�'����
,9i��a��	y��a�	�'?�aG�kF�Q�p��&-#D��[��>.����E�iq�9��&"D����L��)�UkrO9�q�# D���o�4.g�ps�%�4re�}��?D���ӡ��n�Є E�H��U���(D�,��[�5�p����΁\t��VN&D��)2�C>W\b���J�vʹ"'�?D�x�+O?dE@i��$��R��֣*D��cB��$hD��f��s�4x�%�'D�xk���������&����&D�x�����j��;�Y�S���{�:D���dm� &��r�nDh�9(  #D��h�L�Ow���D�o�:dhqa;D�x �(�L���O�|=,h��+D�� B�!��^�{l�H	E�!N�L!�"O��R�DŽ?�L���N:��L��"O�}�c-�14�5�Q�ΊD��-QP"OL�%� u�0��WV-�@{�"O��+��)^�Y[�-h	����"O�e��RgDy2P-I�T(�"O����ha�A�B�`�$"O�	:���7��Qyb�C�F.D�@v�K��T%#�癥��DKDh*D��B�/�?4�n�gD27�VH�*D���b!խ,����S:F�*=k��(D�|Z$)�0F&����)A�×.2D��2߁:V����$�3:�0
7�0D���C& |���w,�!-f����-D�L�wh*��M��E�h�����+D���R䛂>����%��xi6D�@�Q�={���&��6�R��)D��gDԛVs�����0+���'D�l�@H�.�СCS#��U7����'D�����͞k���i��
s�䙘��)D�|˗�I�E��@T��%l��I�,D���D���=M����Ҷ�����%D���#"C:=(�qJ��Ҩd6E�L�<��Ʒz,����+���Æ�[G�<yW��P�F�0�)-��$"Qx�<�B.ψj�� ȒC��	9����I�<��n	&UD���1���:&I�j�<!v�X8#?��&��apnT	��Tj�<1��<Z�-�(,^e0�M�e�<Y�C�'bN@p��HE#r�6u@K�f�<4�׿?$��+@�č
�"�e�<9t�T���r�a���JdB���{�<W�B�T�p0��F/�T}���x�<�A�X�OȮdh 	G�� hk�ǂM�<��&kF�5�NL
 ��Au��J�<��V>���؀��I���Z��Xk�<����2j;(TJ�0$� \�2�P�<iQ̙�j����!�ԱV4X�r��^M�<au-�pQV ڡ���g (I�b��H�<����Q:]@p�^'	��]�d�}�<�� -s+��Q��$@�A�Hq�<y��/�\��p��*:��)	���p�<�A+N.>>�Q#/ڢN�Z͸�%�n�<�
�={^䵩WsxmpR�F@�<a�BɌFV�+���=��Ы$!�U�<	�FK#=i½Bi�o�����O�<�����n\��0x<K@�]O�<����l"�� )[R$j�J�<1r�P0zd�Rʓ�M�"�P*�k�<�J��F�H1�#2��*/i�<�W�Ȅq��4膧ڢR`�zQ˟m�<a�j�l�j�϶���q%��`�<�ˁ_jL�B�ٵ$� �)wf�c�<� �>D2D�FʨA�p����e�<y���3�f����O	^�4,�4��J�<�@�6\B����c�Q�N��)^a�<O�*iY$�i8�m���S\�<�łݔ-��БMX�a�JM�D-�]�<aU�@�+C�AdBʛY%��eJT�<�w��>�jm:��џr��e��VP�<�-=2��@+
����N�<��_0'�xr�KPR�K�#�~�<���~��YE�'��:-a�<��E��<��J�,E%bx8�3��X�<� �%��)��"�|i�R(��G��D�q"Opi+ 5 j���2q�=��"OD0���6����p�B7B;D����g�"2{��i��6N#��2q�7D��#�ۤ������"Z����6D�����
Y����+�$E$�1D�ȁ���|�=xc�@� U�p�.D��	�	�-��T+��^.f��=�g1D� ��➸�,yA��R�lpE��g=D�`���S��P�#,TK�:��5�6D�,;7a,G�Z��q`\)#4�6D�,���+.�����ND��:Vd1D�����]3�RUq��#g�<��	%D���ψ�N�Be�­�Op�m�E=D��7MM�A�zu��bCI�0�XK�<�Qe��p��E�[S&P��MI�<���Ԍ��81����)�IL\�<I��&C eѣ�D�(W����Y�<S�N�_`����0��!�w�?T�0���.{@r�\�Zd��F&D��e�
)a�]I���8��I8�E'D�L�`昃��	P�#
�}gʖ�#D��YU���0 S�bA�"f@"D���#H��d��b�'eB�y{�$D�h3�%λ{������W�9|�B��$D��җ��SO
�R6nZ ��ip`-!D��`�(�
NE�F�h�*��#D�P�ST�z�ôoK�pڞ�q�"5D� H����*j�%D�V
,$�F�%D��R�̟ nYc Hݸ�Pq�(&D�,k�`צ
����٨(�`�g�)D�������d�1���wMT���2D��1�[	� d�@ܟF���G-D�ZV�]Ԓq
�͕K��sT�)D��� �N�"q�SK$ ԍ���,D�P(C�ח-ʬ���$�r�ХXE�4D�p�B���H�S���+R�1Q$�4D�����B�,<;$"/���?D�<@D�ջ��h�3J	�:�Lm1i9D�l��k.Z/���r$q� �c�5D��A�-?��ic˟k��3A>D�l���~~�b��.Y�ڐS��.D�0��# ��ɷ#��� ,D��k�G�0����D����V�)D� �6�J@zJ$"C��'2�T�d�"D���a�R����D%>O�h��?D� ���Ȟa�.Xq��͞c\D�*D���䤚�p(�	��:b�D�w)$D��*��/Z���)�J�;H�ڼ�QA!D��"L�*W��a�3��N��H8�>D��+�H�r�i���\w����//D����[�/��mC��B߈�f/D��`��O� ¢�\`({��-D��'$J�}�^�*�a�'a%�9چ�1D�ম�{x��Cn�5s�$�0�0D��1@��(�Cp�T����C*D����"�hX9)�o_�`AC#D��(g� �(s�\�/�&U��J lO�㞌kEB(D�d����#	l޸�TE3D���!��ku��rA	n� ��<D�\�҇�2�`�Q��n�If�:D���HH���D�H'@|���7D�TXP?(bl��D��GDژ�p�0D���dC�	2�����k��x�6�.D�� .lZSE��[���3�a$ee��P%"Of����5&�΄���6K��0"OƬ´�Fڶ��v)G�0i�2�,�S�ӽ)ص[0��"<���b�ː�$o�B�	|��Z�
8=�}��	N&��p?�W��q8�@7�қ['f�b��k�<ǁ@�S���"�%O�6}��^M�<��F͜h��I���ȚH�~,֡H�<Y���AH��rB�E�C!@�z��l�<	���2��p��Ĺ\��t�1%b�<�FH��,�T�3b�u�R1���Sh�<gb1`�,�*��j��R�#d�<�i��a��d��e��VI���\�'�?YP�$E1z��HP�I͂0���k�!D�T��#�O�<9Ұ-�싲�+D�˧��A�|=:�Q�30��	�C(D��i�K�}�~}�Q!O����y�"*D����bŏs��)D�I*nM�ɹ�'D�`��
�[�5ZE��H�0���%D�d���xЩ�GRS��#D��Q��*B�Z�C��
�}+��3�'E��E@�b)�
�NI�E$��yR$U4r��!`�lr���WM��yr�\�v�8Ys�e�f��cӨ�yR
��g5�����
,��5 ��yB�\�N/@��I�o��Ȩ�L���y���0i��s�	�mT�D�CD^-�y��� ���+C&a[��#@���y��V��e��IS�B����I��y�e��n�r�H��f\��:2@�A[�=E���|,����B� k5��
�D���=��ՃbkH�s����a-�B��cs��FDT/�F=h�BݤB�ɩ!)�y�×=,F����R(~��B�h~���\�yE*!���]�C�lB��0A�4R!�#j�vH3�C�I!9�Y�F¦ �8r�!�Y�*C�	�g_ؐR�����rG�1�B䉺e.2����V'fn�a@��I
�B�I�+�����B�\�;-i�O:�=�~:�%��b����P��)�* �q�_�<AA�F�P�#Bb�j�;�^�<��E���b�#�:�NkdH�V�<ien��\��s�V�5�����O�<��E���(2�
�*^:�z0(�N�<��ġ� �)��S�EM&��s��a�<�`jZ�1�&l��Lz�h�f�Ds�<)�,J<O�|�p�	Z�sqT+��^l�<�W"Я D�[���U6���I��<1���Q�J��`fR�KD�`#�W�`��C�	}���x��T#&M^�7��~2B䉶&
�u"��V�(� �'UtB�I��0�C�JX<+h��F�P{�C�8+�8� !�Q�`z�e����l�0C�y𢙓��ZD��
D�'NVB��O�Ę��C�Jۺr �ȒBB�Ɇ{@0XRA��lBX-9����6��c��G{J|��'�9	������ʧ]��v�y�<�#�
e�xW�ߊ~����lx�<A��-�|��*�opKcJ�t�<�2O�7$-,�3eM��%E, ���u�<��.\�V��[v�"E�:T�x�#g�)[���Æ.�8p�a�*;D�����16>҄�1�w�;�.7D�� ���X3KYb��I���m�"O$�&�@�p�tB2חm���"O�p��B�3'%���&/˂tV�h�"O�IQ��@�A�uJ<|S:�"O�4�s�[�Ww��)%��
RDn��D"O$$�֡Y%'� ��GK�1̀ gU�p��I!H�PЫ�A;M\8R�߶e<PB�I�%s@�[LT9[�HR,_�t�d���>�A�\��2V�&�vI��K��m!��?��|I�g$g���K� ER�!��A8��ۑEѺ:x�Z�L��>�!�$S�\�.�RU�ڴP;Z�`�6s!�$(A�q�qF�� .��r$�.LW!�$�({�|���X1"+^��v��?�!�D�E�4
��^&��J��@5�!򤆉4:��[�V�P�|Ш��� g�!���:Ҝa�W%��1�
6�!򤅻%+��� �7�	"�B�<�!���A��jG|�-:Ӏ�$w�!��5I�
i�$J�B>�@0@�&�!�*>�J8x� 
=j���{��R�%�!�d�?1�Ps��#u������r�!���r:pL�g��"�����*'!�!r)X��4��E�^�S��H5�!�D��$��@��r�1�@
J�!�d���(]����Y��!��T�{֔@r��' B�ћE/�*"�!�d�('���"$�6$,��0S.	� !�d�_�q����g����1!�dT�}}(�a�"j��
À�51�!�D��E��#���Yl �� ˫<�!�ː
U�Ř��L
A@��01���g�!��X�1��� �+�.%+@�>�!�d��g�|�V*�t���ZP�&8�!��*�-k�%�yg�0Y#j�!�!��F<z��Ye���Yl��	���!��ܥQB�|�Z-ApY)�H�
!��jj�m�
h vћ���N!���g�döȴ*b��fc[,6�!���*�X�k��]nr�C$�39�!�d6�4m�QVaY Y����|q!�	+��y �D!�"థ��9 b!�D�A�>}R��D��9f∜_k!�䖑1�.�X���%Cm�h��0k!��_�5��k�D��
R��%O1N!�Q�΢�b�gZ���"@�ÞM!�$�-Rb�K�L�����)�NC!���S�܄P�f��ێ9I��	s=!��D%R> hA[�~��vj	r$!�;^���@�$"���7�~�U�ȓQ��#S@�5x9$Р'%h� ��P�p0c��)zUj]C��̦l��ȓ~���B�ت�x0�cυ�	Rd�ȓk�ı�Eҙ���W
D��������F �*����Ƌ�S�.�� �䝻a�2Ș���GS}���ȓ4�j�1�kɟu���Ӥ��<��i�ȓ.�5`A�P�!�Āb�<-w؆ȓ7����$P�4Q�`�# @z���}��J@��&��1�����x<a�ȓc��2�+@;�@@�V8Rl�ȓf龁f�D�������A�ȓ��t˖=_� i����1D?�x�ȓ;��ШP S1)Q��"*AfŻ�S�? >q򕏋(�@��/��0-�1�"OjٚcM�5�Ȍ{�.2P3�U�"O��!&!S�@�8�i�F���4D���cF"b��b%�*Ak.X�D D��1 i6���HF̹S���&/)D�8���	*o�>̒�j�iȩ�fc&D�����@���W��R�th	�%D�(��/�&mZ	� f�+vl4t��8D�����6/j�)'C�th�H��5D�l���gI �t�.�*��6�.D�p	%aށ(��C �*P���F�(D��c���'^c����Ձ:������"D�H���� |0�1���<����!)3D�(K�-ޟ�
Mb"DX�֍j�*.D��+�a˩HG�m��/TO¶Q��	-D��	Di*'^�
d!ϛ}:�
�)D��csAb��3�K^�d]�`"4D�@ Vb:R�}�	G}2I��g6D��Qr��<+�u�A@�� �����.D�L��k�#(Cq�ҏ}��x8Fd,D�#�ə�?`xa�d;x��zb(%D�<��Κ�3)���{���"g$D� ���K#eTI�����!1$I"D�h�A,B!KƊ�猈�����#�3D�|X"@���X�G!&����5D���� PB���Y8�V��F'D������i'rp�
��&m���&D�������|&	��+)�
-ن
?D����(����	�T�M4���%)>D�4p�P�o��ne@&L���'/D��c�o�?��|H4��	|6� -D��!`��W�x�)ԯ�PE;��+D��Q�$'����5�}� )C%�*D�\S����g�2��E��UK�P Մ)D���Ɗ��W���h;g�mKs�1D��SaJ�!t)��[� �J��.D�����#o"����H�m���d�,D� Ȇ(G���ݑE�G����0�8D�H�#OB<; ��,���ܚ�2D�X �&R�R�A�t$�,X(��j�$;D�쉄-3q�ܨ
��۔�9���:D���v뉈1l�@e
Z�;	�uh��*D��`v�n�$� G�#l�~���*Oȕ�Э�k@pi��д#�0� �"O2e{tKK 7�*�4�Y�	F��9!"Oz5�惈)7�m{6e��XTT�#"O�%����l-�r�5'|��"O ���+3ې�Ô�-��u*�"O.�B%N�?,��d�ӀB#�$C"O�t���O�𖈫di]�<���ٲ"OH\i����WL��≻#��Yq�"O�Lq@�*\��-��ON_k��3�"O`Yke�'@*r�eh�ldU�a"O�$`�C�[�l�uFYlM��Q"Oހ��B�"cK^<�t�*n(L��"O^�2Eӊs�tE�f��o���"Ox9d�֫E� p8g�qӾ�"O�=0fj�k��q�kJ�Z�x���"O�*����YH ��
Q�~��;"O�J��}�6�bV=R�>�S"O��W�$=B�9	�
� �!#�"O��a`�|cD��/��z�� ��"O�Pʔ�P�HErs�U�j��Ф"O`�I"K��v$��Kw��T�L��4"O� �48���$*��9��ݾl���"O���s�Oy�`��$KPC�9�"OBT 3�/e��uI��8>a2�"O�ȡG��2{��T��� s)��"O��v��}<4�kW���ћ�"O�I+�a}��]ҦG 7��� �"O�!�F���s��vĢ<��"O:�"�J��(Pf��й($"O��*�i�(PѤ�Ӷ6ȞY!�"O IR4nES�± 2#W1I��)��"O�l(t�6)�������c`"Op���Z5ya���[�9����"O�\���U� c�Jp�T9��"Ohи�dX�`��83D�M-���ٷ"O���HĶ^��dâ[OU�a"Oy�׋�1uQxMa���s�VQ2�"O��S�F�6Z%��8���ZA"O�J��ěb֠����KM�=!r"O����+psf��6�O:�"O�Ӡ�d]�su�њn�H)ё"OV�yrFG'�-���	�7(P���"O��Z���8?H0�3֩�v�,�KQ"O�쪧(�9�\�sP��=�D�0a"O��H��?��%��j��Ұ��"O\��uT���-���ѕ&Z� �"O��J�١DK���5�D�8�d��"Oj��\�}�*X3%���@�G"O:�0$B��1��mK��l��"O��{�	�� �,M�LD:4�~(!"O���B�.t���1��#trH�3"Ob̐���:�UZyf��k#"OR �,�4H��0�rd�aoH,��"O@�sEDH���Li���"�H�Z�!�N�2!Љkf���Z�P���(V3b�!�� 4Q�6��s�-G��,95MR�+p!�Ě�#^�i3F�4Z���Q라56!�D� -�ձ��k�4<���C�!�d[~�<���mZ����Q�!�$�)'�2��C�#u$�pza���R�!���<�N��CD 8Jh����#.�!�M� ��]��ˁ�: �Å/Z�>�!��-0&$�2�ᙗQ����L��!��ϸ=��H�F�RU0.��5��'>�Lh�O�/b9`�1f�	�9�2P��'���I��5'�XE뎕2����'���W��f��Hj�A��'���'L.�o�2y7f��)��'�|Y�'NB�b ��&�.t[r��)��dZ�'T����=�� RO�w�����'FV�j�
I)��D�?�� q�':�-	'ƀ.|�<=��,��� 	��'���s0O���.��Rc�7�P��'�c0��O�yB���<� �'�h5B��N(nD�C��n�]s�'G.�,2Kp��c��1���'�@{�Ǐ<ؐI��J$�4|�
�',��#�&���pkW!��f�X�'�^�p�
�4h<J�X%
���X�'^n#�d�#sLu�PHA�j���y	�'�TӁn�5V�xЂ�"7O��'~q�IB�f�V	�'퍌}�b��'� ��#,S�h���І�����'��=)�+b�8@�Ț.�X�
�'��xP�Þ'7�u�%��"K���	��� �Rc)g�0)á	V�6/��)c"O��
A�L,H,PzA��>@T��g"O�y�#�|�|�C���b�0�w"O��AoJ<���4�I��ր;�"O��DL�M@؝`�E(r�n�D"O*LKE*��	+n����Pq�`��"O�h����)�` ��Rg�:ĘD"O�8J1"ŧI���q�cL15�t�Z�"Oɨu�F U.��@�i�.b�4�"O�X��Ua��X�"�Kj����"OMӄ߽z��(�G��{PzEy�"Oư�A��)dUYp��*p��!'"OT����Ѫ-⠨�Gry<�a"O��b��]�+O�<{���: u�A��"OV$æf6Qv>���D&irA{c"O!���M�.�� 
A`���"O��{�d��Bq���ׂ׶g_���"O2�{6�(gZ��[��G�Y����"O ���G3Ҡl�$-��\ ����"O�`sOS9>,����	�^��p"O�@6�ȅ�4:ӌ�,!��!{T"O��	�BX�l�M���-��	�B"O�AC@�5Z���5,��L��"O	���C�Y���u [?ELc�"O���OP�Ƀ��@  -��U"O̥P�~|,�Kd`�n�P�"O�92���0�Ƅ#��È6�@�#�"OVJ��\9w`!�V����i��"Om�I�}R8eks�̥ip�s�"O1ɖ�U�i(��Q�-y{�"OX�3#"�/MBU�C���r�k�"O `���Ŷ'l����P�V�4M;�"Oz����5.�ݺ��E�؈(�"O�����%J�( }�#5"Or�[���5��(���
�pup"OT�H�EG#ƞ��D�*�Ti��"O��Yq��/A<=�1n�V!~l�a"O��J�d�
H�H S�-�̊�"O�m3�C^?��Bp+�3G�lke"O$��ʻ"�>$kҏ�;�iQh�<�"��:^X�F�9
54�@vNg�<	�OG&7~��"-�7�����
y�<9�&Q�J�T���N,9 ��Fx�<9tg�� N:0@w &rw�T8t�<���F5�����:Dh�kZX�<aƀ�qo�]�@\A�ċV��N�<Y��[,
$b�P'gQ�v:����e�<�5��%l�a0̘�-��]��^�<����/fZ*�ܵV扢��_�<���/
d>,���ɮ �q �X�<����\�P�c� �)Y�չ�H�P�<��)����=(/�'F�MY
�I�<)��2������S':�&�YPjG�<�
�����$� 6�F���VC�<Ӧ@?&���w��%VhQ@ �y�<IU��<+�ReDةj׆���B T�Ȼ7I^B��*hF*'U�P�?D�d
��Q�x��M�6� ?`�I��)D� �wm�!��Lp��_�>$� H"D�0�R&N&�p1b���3/S`�5�#D�)�Bt�.�1d�޽Ah��g#D�l �@ЯpaI��ћo���Z�,+D�$�`��C��9 O31���wO*D���֍[><z] ��^,Hc赨�e(D�� 2����2dp�h��U��t3 "O�� �r���+q��1*�x�"O-���^��,d�T�s��]2p"Or�� ?�((�.҉I+�e٦"O�����M91�@���K�=qȪ���"Of��R��ee��(�����Pt��"O������2�F��� �Yy'"Ory��� �D���ĆMy��@��"O�eA�EQ.&��P*g�8B��)[c"O��pA�s̐-"7O_�>��� D"O�03b޳I�B�s��\u�ڨkw"Oм�H���}�tm��}æ]:S"O�س�uȢX��B,U97"O�ja��-	��qA�ڶM���0�"O��N��U�&L�с�\��i�q"O�0��C��hؔšpA��r,�=KA"ON	�boK(^	ڨ���
�r�hv"O�mQ�?M��A�nCQf��"O��W�����,�P�Ќ�w"OT�%�_�'.��b�Z~�L;t"O���2� \7�$�C�Ee�Y�c"O�ݪӊ_�P<�"��7J"�BD"ON���k�@j�D�C��(&���	Q"Od}��c��DqX)X�gQ!sk�*�"O�͢.O�@��ԛ#�̓tg�C"O�����"��P�F���� �+E"O�*V�b �V��	2��VGZ(�y�l�>kO�m�l��`@V-��y"�Ќ�r������m�0D@��y�#�6\&�ՙf�g��*��D��yR��+|_�ԑ��b�1QU���y"	�-�HP�n5%�*��(ٙ�y��A� ^,����"�*yKd���yR��q4�i�͓8I��EF6�y"J�iC4���dҌ�>E"r��y�`��6N�e3���u��H��y�۷>���)f��208Izֶy8!��H�����DZ�*��Q솁�!��أoZ��!lʌP��Tyc�I�r����Y-:~ �e FN�ps���y��Y8Y4[�M*G; ȷiM��y�GX�.ٚp�SA�nP�Q&@�y���CO��A~4��5����yrh�k+@���ڒ"�&S%oY<�y2���BA�.{���k�BP]ĥh�'a�H��Mת?]�D� GVST��
�'Ɩ���/��D��;�hD.�|@�'��%c0
�+��`�Ü��lU��'�NL!,BF���,ٺ`(Q�'xL�3�#TlfuS�n��p�$,��'pN�#� E��{6b�.h�'��dq�^�11n��#Lg�fL��'QX��U��^)j�*բG�Wɸd0�'l�A�E�T�*�Ҝ��N�V��mq�'���JC�5�:aò`��Q����'8αy���yfź��_ ]|�%��'�����f-Des���Y�JX��'tl-��D2aT��k�%[I��P�'2L�Z��
�袀Z� ª*WrC�	��8YH�k͗aTp�ڰg �=.zC� z
$ꁗ~�3�	�h�pC�	�IUh�a�#]�ip�M;��zs6C�S`��d�x8��`�C�	�|n�!ҧ��n�t�8ţ�0?�C�)� ~������Iֵ�5
�Rk8���"O�`���K�v����&��*c��Jv"O��V
Z�&��)�-*uQ�Ԫ�"O�U���2)D����ڄx<&T��"O`1�R�P/BP%�t��2
G�uY�"O���ǃ�r)|��Eˎ89U����"O�	ФB8:Zؖ�R�Z�<*�"O��[&�@7}��,���lP��"O��2�G�#�ڴԤ� /�>-Q�"OF�J�N(`��h���@>�@1,�y�i+��A1�����)хjĩ�y��,l�(�e�#y�^� b`٬�y���8����e�5j
��:1 ���y��J�v�P���-^�x���+��yr�Yi�
2A��e�|ЖD��yb���$8l�1LG]����E��y����F�j��eYFEʕ�տ�y� IH��S�P
�E���y�J�J�T�B%Il�[����y¤=]�(1Zc�57d����
�y�mH�8Q8vǒ4.݋b�P��yχ5�Rd��I]�.�� �H�>�y¢	�`>���Z�V��Y�ׁ���y�N�R�9Z��ٯ�D��g"�y�M���Q8����窭��'W8�y"�2� ����@r�
�*�y��O.C�����3F&��ҧ�$�yb��Z�J�+��+H^��C�a߉�yR�� 1�%ڰ�X�L<�ꑀ��y����A؂��DI��y
䔀qo���y� 2�ZQs��-w�(��P��y2c�:�=:Q��	k�ة�B� ��yZM��ٲ҈��r���a���%��B�IB�nUR �vlhq�	9b�^B䉴jQn![�oٛkL�b�**A��B�	 e#�����L<�&�OTnC�	�a��%�
!h9��O,-�B䉯|]��k6�S�4�0'�0[*B�IN=�HzG�U|�L�@��6��C䉕c�b�p���"�P���
9�C��&wN��@�K���8��dNC�I&z.�ԛ��B/���B7wJC�ɖ*�Г�ŕ�#`P�uB��WPtB�Ɉy�h�D��
\4Yq�_�=j�B�I9Z8�R#T���ݳS	I'C䉇M�FP�PC
�񲦂�� �'=���b�N&(���%¶>�
�'��R��A�I`���Ds�h�'�"�a�-&e�,�z�hQC��h�'�����A��B���:�B�)Q��$��'X�dcǪ_/�4��v�E�J_~���'�ѫ6�58$Mh�"ݳ@�*�q�'C:p)��H�^Odlrd��a�x��'���@+79�����\�b]��'A��j��:r@
����h��	�'mH�bB�=E1�WE0*��|��'3"���X)����!h�"�'Z6Y�\��x҅�^�mldx�'��!����2��G ޝ_,�[�'�.qHp��"��2���	��T��'����"I�W^]Y%�^*Y����',����9�f<je/E�'�`�;�'��1v A�<@`���!Q���'�
�×�ƨP��h�"�I/*X������ ��J���n����`K^Mb�0�A"O:(��,j��:�)�8�b�jA"O樳g/�����3锇?Ԇ��D"Oj�;B���A��\�@i�S"OVD��e�'4z�<�`�6���V"O�� p"�9gX�A�1��0��D2�"Ot�s#����ڼW��!z:���"O����DD��Q��K�K~��s"OX��'0x�Ԉ{��M�oA:Q#�"OfA���@ƶ�z�n��s��QXt"O�)������ñ�Ec2��"O��pU$]H/� CV�*O�1pP"OR�����]s�P��N��M6�Bu"O&�3�琳.x�B���/I�̨�"O"虗��-� !"uEЋv.Ȱ9�"ObMhӢЉY�r�c�ȭ%AB"OVp@".�_� �#�	k8�0��"OE8�N@/�>h3��D@�ة%"O��J6 \�V�)�AL)n%>`��"O�HYp�άE0jm)�eϵ ��� 5"O�!z����.��9�"�/Cn�#5"O�0�"��9���P<*�!�"OP�G�C0���փ
�MN��"O��X��D���9iV����-S�"O��c�
EP�����@p8u��"Oڥ�"��_�����lW��@$"O��Q�@�gJ(�c��]/cE В$"OD�1���ъ''H<	;"��F"O$�X��	R�<�z�'w���b"O�pٕ�W�j�(��eǨ!{|�S�"O����/	t��6E�`Q�`�"O��U��5|&�5��6B옠"OH����/�؅�Rd��T�<��C"O4qQ�+�	Eb-����>ܦM"O�;i*'�L#7)�#>z�Ѫ�"O��Q1ʤtZx�J�M֒y ��$"O��[��ΩV�$�[wOߒw�؈"O�J!�� Y��MI&}ku��"O����nX�N�t�j@�:eA"OnD{ #�vLr���Ȁ']�e��"O��I!F�m�ͩ���� B�UD"O𤢵�M,W����`��>M�""O�RůT����S��t��9�0"OH����Q�b�Q��%r��S"O�u�7j��u���z 
<^�豀`"O��+��@�D��U������"O�A���@�=�Ģ���-Ȃ��"O4���Δe;$|BV���^-8v"O�	�Z��F4��(��Czpyc"O�!���ʁa��)���Վi���Z"O� �+�e��!��oڐ7��!;�"O����	!R%�r���T�ȷ"O��"�	{�R�!U�S��+	�'�X���NMx���e�M�T.|ԙ�'�$H�   q�r�y�C#[=����'�hm��k���`��<j(��'��<;��4c5h�tn�'��$��'°زDC�_]>@��ĥNY��3�'_�!q�
��j2��rhɋNQZp��'��Y�B�Z
"���Q�蓫B�ب��'@���D	� �KB;[dU1�'����`�P1��)���ѕ&��=	�'��;�	�W�\�r׉$)h���'Q����#ꝂD�,����� ؈�檆�	TVE�5S@�Q"�"O<-��F$+T �@�ñ'^B2"O&��!��Zܸe�	�#@)��'@��B�ʂ@OZa7@=vFl�'�
�!��*�i�U V�ovv4��'aF���~c��Ӹ4�Д��'�������<OTl(�ϯu��$:�'�.]�3�;D�з �
:=�"�'v��'ֲW�����	Эc�'�� ��Z':�"U�F�����'�f��Yʮ�J�J �"���e+D���Յ�,bF`��D�u�$��\"!�D�?f�̽X0a�6n�BhQ%"���Py��
7$��H&I�}�5���y����!�]��c��(?��T*Q�y2�T�M�3T@�w�n�!���3�y�%�)2�����8��Z.�yR�ŹS�$��׫�<�nU�E�X��y�+Md�tl�sO�-E�j�W��y2�M5��D�'i��G
 ��*J��y��;<���ʱț�񦁚f*�4�y���Mb�p�2� A&�?�y��q�>y-%�h�Ӷ,�"h�ĄȓB�,�$ޗ c4�����S,����(�2	�6�ۅE�,#OҘp���ȓ�$�v�)��P��+�ч�K|��'��k�̹3��3ߦ	�ȓ���പV1~��<{�A+P!��	�~��r��o�nx� �3���ld�u�����I)��ЁEW��H�ȓ@������'�0���]4LB����K�ݙR�=#(db3!Z��&��ȓS2�)�cY�9S e;s	���ԇ��:1��c�n��{r�wT�4����Jc��)����b0Їȓ&�5��J^�*Tddc�%̐QOLe�ȓv�"q�Q�J��]����{܀���V�`���{{7_e��d��']�HC'�E 2�ȉ��mܫc� }A�'��]�	�h1����*Ҙ^��#�'lڅ˴��8��`�h؏Z�ֽ[	�'�Ќ��@͠Co\�+�l�T��	�'��5�\�w2��k�7<�
A�	�'Pf%�!���(�Z)�g큈:7Z�8	�'�&�#S ��v�]�w��_ю���'��A�W�3�t�� @sn���'v�3�
�Z��!ó2|z���'$@��'!jw|�2w�,*S`��' X�5D�8GuV�+��&*���x�'�B��R"sm����Jøj��l8�'<�F��>(.dB�"�/P��<0�'��Ah;$�$ 1���'N�$Ś�'��p����=�p㪆[D����''8��%���^�>P@��X�T&��	�'-8Ⱥ�>}�����Ιۢ��	�'*��DH�6ЖeA�d��|��	�'���"��2|��4�DS��3	�'�"a�X��͌�K��g�H6�y�ԋbmxDaq��+�P�L��y�!Yx�m��B�  �@Y@roԎ�ydJ?����Oɳ)aܸ!���y�+��9<�5�+/����-])�y�̇�s��A��'�.�@E�N�y2X�"ɪ4�f��%�ѣ��
�y
� ���)n�:��_Gs4��"O�St�ëB�n��	U(]�|e"O$��T�2hBDp'N:h��%�"O �
����\� �e�����h�"O6a�5��E_�����.gv5 �"O$�h�(��z4@��b�~��&"O �����Qvb��'Ĝ>I�%@P"O��XFb��b��ڟY� 9Pd"OXؐq�H��l<�F�$ހ��"O. 9ڸN*������t�`�#D��ZI �4�4��B�ah�@a#D�<␍S<��x%�үy�����K'D�rK%-�d�Q����j1�2D� �D���,�q'U�Ph�*#G/D��qMO:ox��q���, ʴ�-D���!.9|�B ӓ�Q���
�	6D��"��הm�Tm� �M�'阍��	3D�T�1l	w�bѸe�Qw��	�6D��	��Y�;p�����ɳ�b5#�� D��a��$[�X@ ���]#��>D����A�T��K���s�y��<D��HpfCh� � !Jy����6D�
sBV�NH��A��[���W5D�tJ4CR�C���9�䄰[.�YB�-4D����3It)c�@W�&DV1�Ae=D���Co�aRZ�ˇ
�U4���/<D�L3Q��%L-���b�&x����>D�ȨsI��tҾ!2�.J�=&�9�#D D����G=�T�ӥ���3�x}R�<D�LB�/�� r�R��'����0�6D�������N���\>a���2�3D����g1�6�@�&�3}�fQ0�k0D�؃�m�:h:� �L��B���C1D�@�옞� �S$"�f����#D��Q�f! �����
s���%C%D�ȠEJ�hg��K�Y����$D�t[g��O���A��D1P���`$c#D���	QJ��%h�xd1P�<D�@�Fۇ6����qM��crD r�D;D�8c��H ��"$� �@$��c<D��$3p���A �.��M�&D�������D��	B���' D�TQc
5UKX��nG)L笐 �>D�XVn�������MR"rT�7+;D�09�H��f(�7hS�o�����8D���.��_����u&Ww�~ ���8D� Sp�/� ���S�!"L��5!;D�����ҽb��ǩӟjlJH:�,D����)�$5��@#a�M��P[F�(D���5��n!�rC*L1V��<��'D���ab	�	���0UMJ/,���I'/'D����[�.>�(cf	�P���0��9D��� ��KN�l���ӣ%��+�2D���)B)2��Y4�u1��
!$.D��H�Q�?�I@DZXMl���-D����M^�g�0S7�-�d���.D� �d������!�0zOR�	��,D�xx5��B�vU ю�>Q�"MP�@+D�t�rL\)2�2HI�]�[��8��3D����
Mj֜�t?+[�e��A7T��y3�H�g^�a���\�t"O�)@۾ �޽B N����"O6��ń��]_^}a�!�65Cv"O���h �~���s-�K̦p�"O� �(2+[�b6���B�����"O�x���Et����C�6�`]�"Oܹb��¾ �R�Af�T� ����P"O��g�Z(J��w�V0Y�9H�"O�a�B����a	U��1�`ARv"O��{#��(��t�T@
�.�)`R"O^�+�iͅ.��i��ݗYB�b"O2e/6�4���`Κ =��r"O"l��_(K�t	�o
A!�r�"O�8�'�OJ�4��D9�:G"O���m�K|B�۳
#��1��"O���F�8hn�$�I$0�X���"O�a�!:�+�ܨZY��@"Or��u�Ďp��G`T�o� 9
""O��TB��FL`�e�Z�`���"Ov�1��]t�L,��B�t��m�"O�|�J^ 0�bLIg��T\l��"O�}gc�+gpL1�RZR�IA�"O�5��_L�"xk�U�q,�@�G"O
dr꟬U�0؅n�쉲"O���1�s�TP���V�u�B�B�"Oz���K�!sl�AK��V�K����b"O�d�r��5���A�Y�A�r�PT"O$EaW�[,z�41���G&	�u8D"O�����2J�Q �H�jQ I�"O� Ƒ�mr���t]�֏L�<wd]��LEY��M�*�H�m]_�<a�ȟ��m����D*L�h���P�<9�p�Nl�T�fA�[`"�K�<!b�Ԋ0;� k�$� >&�5,r�<�ua͘�r|së�X�5�4�I�<acH�<$���P0d�^�H�c�D�<)���&3.�p
�,~t�aP�K�<�aH����:e&0KƂ��gGXC�<QS8h�`|)�_h�| 0��S�<�1(Z���W�@�Gۼ���C@P�<y�lܳ4�3nK�$�x�!EV�<�V �0
����@�|�I�-�S�<)7�Գ2]�� ��>��L3�O�w�<�$�]-��Aq�*�
�-0H�L�<�u.�� ���aY>K�LM�v�J�<٤��uH��8��x[��AD�<�����3t� 0A�=��c��u�<��-ۓN["�ӦDa�x9J��v�<I!&�S�t�P�&�1#����e�s�<y�E��f�v��ċ�7Wq�(`��V�<�u�B?�"(��&�N�|����Q�<�$�7'l(�c�Q�D�\y6�L�<1w�</ǆ�$��O��Di���H�<Q�FY�*����5��*`۰k
E�<i�,˰����.;�P;��g�<�`3Q"<FD %%8� �GE{�<�T\�t�=y�-�!s;"$)G� w�<�&�����1�#��!^*D��It�<���LE�	��� <�Y�#q�<��@�-5�-Y�`��%�5��k�<� -I�<'�E B��턀�q�Q�<ن#ίM��P�f�cR��Յ�M�<!rhL�:@S��K(��x�M�K�<��A\�2��(�A�ɨ'�.�QI�<�B��w�@����X�1��z�<�5pU�"#$��@[��O�<q�'ȆAV�A��8p �BfN�<9D�D�&�N�qR/O�~Gؑ"f(�b�<� PQ[ȓ�D���GA�&��� "O$����q��(3�Y$D�.�h�"OмCf�K���)c�]�m�`"O��T �.vxJ�UL�;`�]��"O��
��F f"�
�k�x&���"O6�#��<TB�	�ꀇÜщ�"O�5"�A�t�(m��
��B���"O^�$	�.H��Q�D8~���"OF��%�©sԝ�A�{�~Y�"O������a���7�4{ bps�"O`e:q�P!�����(����"O��P��B4�(�81#
��U"O�q��8@�`Ы�2�Z�r "OB�F��
��1�E-E�I~N �3"O��sAd�H��z2�U�S^��3�"Oʽ�CnN�{!�M���k��)3"O�����*��hA#� �Ʌ"O�!n&C¦1#�Y���1"O@��	�.u��-	%i=dѸ8��"O���$�#9lb�D%��v"O@i��`c�0���0�.E0P"O���d���m�=�J�DH]�!�$�!}�@.ں3-vx�]�@���'r����6"������#�Ԁ�'u�97�&t��`��d��'����'P�~����?|���r�'�B�a��%�$2��Y�H�j)h
�'���Zς�>�a NA�S5��
�'� =i10q�ܨ�@ʖ�QCX�
�'NȬ9�
Z��q�B0:�(��	�'Dș�E�N�[ R5)0�1(�	�	�'������ &�8�yR+k���'�>�2���M�p%���_a ��
�'Y�����=e9N�"�eؾN|�}
�'������@1��Y�DLʑD��L�	�'�Y #�����{�h��D��<	�'�������4H�|� ��@����	�'�� ��V�V�f!���&IC䍈�'�0h�0M�Lܓ��?;�$e)�'d�)�v�U�J_,xqd'�^���'�I&KJy�jD��9V�ȸB	�'�E��k�F2��TO�h�[�'��R jH-S��̨�
�W0�c�'���'+A�i���pA\�XW&�X�'||%1A2�FL*t�T����'=����)��\]�-���EAPP��'�����]M�jl�U�@�)H
�'1fP)D�^=L+�,,S�7؀i�
�'&���g��	���oM>ڍ[�'��}�0�B+oږ��f�Mc�t�
�'���pfJ[I���BN�q �UB
�'�дQ��<`0r�1�/�j�,X;�'q�ۦ�Z%JM�n�'cD�[
�'����ob�HJ�:Q
�'�������-A_����J�s�=�
�'�j�'U&���J�%`G�)S�''"D�3������
�FӬ
�'�"���6ݮ}�vGה9|�	�'ߦ�h3�3P�F�z�J�?�� Z�'�x�!�GV>X�|5����GY$��'���C�ٜ`���6͖�7b��'�FŻ��I�V�z�kV�L�C���'m�9�)�&F�i13���C䉙E�H�²�Ƥ?0^�Ҥ�]�{��C�)� ҭx�L�/ij�#��K�B���B�"On�!s�[J[0��a�Ӡ^#H�C�"OR��cc�[�B��Ӑ&aQ�"Ol����,���b�bh�iv"O��ҕ*T*Du\xz��!3$=I4"O���C)U�p�	�e�͡��pi "O�H)m�>�(�0�7�NL�F"O�ت�KD�)j
M��E��Kp"OB����U;�9�H7l�L��"O\�6B�h��`P��_�Lr�ܫP"O�L����'4S��㓮ܱv��5��"O��b�Q!|b���#�/�,�Jf"OTt¦�*G�x�A!o�0!T"O2d�g�N�7T8}cGn�2�Tī5"OD�	��J�ͻC.���&y�"O�s��$z�����y5��qs"O�)Yi�*#Zl�J�<d��l�"Ot���d�� j�"����|��"O�Hq-^�%�0L�2dC��V(ӷ"O�i�+�1ވ��(�:�h�"O�T�ա�"c��zt�WXyZ�C"O�Ѱ�� �rR��2��5� s"OP9铍]v|tqBX�m�"2�"OR�95O�ޢ�b�F�;��"Ob�K/M�g��AG���,U�"O�Tя@
	�@a*@��[����"O(y�P�M�=�,�;WiN�u�!�"O��BukW���t�&H�'J�ltrb"O0붠�+8�
%SU��-��p�5"O�Qr�i]�AL���
�_ۤ4��"Ol�����l���0�	����2"O�E7.� =H
�!�o�Y�$�%"O.]��W�?`6�)rE_�P�X�'�\���jNev���oזT����'��I�Dþ=X�$8�̙�.��'�p�����V����K�!"��m��'�� Ǉ�G+�3�D�Q�NŻ�'2�� B����$�B.Rw��-��'�,�f�.��@q�KB0�!+�'LN��ʿ:�-��@�I%��@�'��}1�ፀm��=��h*
:C
�'L>0��kIe0�8����W�0Ԣ	�'�$Y���'+JUQG$�%-�!"�'���oQ�@
�8D̈1o\��'��}⇌�)�xac�hL9�����'�r!��$ ��c�:�y�'Y�TBc*\�S�FAr+�5W� 
�'�><��k^.���#Z�zr8(�'vJ�CW� �5]b��wc���E��'/�c�*ǒQxD�؆�u�`5i�'Zf ;��=|@���dn͔�A�'ْ���!A����CW/�PC�'����F�n�PpY�J�Q]:Ix�'p[�E"!t:���[
P����'Ķ���^�WG�̑�)G�P����'�bI�2�
���0�дw�*5��'Nb�e���X%.��'�0vO蔁�'A�U��@�v�����4s�2��	�'��!+�bU�͸ ʄH�4��	�'�,��,Y�Q���ծ�7b���'�4[���}n:l8c�U�
(����'..Aٓ�H�\����"�ڴnax��'T�hV���#<V��1%�r+
���'��	@����2�p\���Ƃ>�:����� �<s��N�50rT"fI�'p���ò"O�r�ND�W6L{��J�8�b�"Oz�H�j���t9��ϋl"I0�"OL�!�6P�fQ�#��6�dQ�"ORcVD��5��iH��	�` �"O�pa�o�(a�\x ��Z7^p�5"O�Ab扐��hp���.a��"O��p�_�bR�5��n\j,�u"Of�(#j&�=kD�`�B��4"O<,�3�rl hd�D��Ip "O>h&̊4����!�O��*�"O�X���S�4�m�'�5y:���"O-��i�nh���37N���p"O*X�5�[)H�H���16P0k�"O����N��@`fy��m0U0�`Sg"O�j��-H����DL8"HJv"O����r~~��d����U"OܴI`��+�R��E������"O���<��[�H�1�`m�"OqRWB����B��#7p���"Oj�o�+?��5ؠe�(Шd�"Ol�B���$E�0���'��Q
�"O9ʢa�54�Ĺ�^�0Y8P
"O`��	�1St�)ਈ,?M�9r�"O�d���åO���p7'X�JG���"O�i+`�ۧ\xeh�փa<�("ORP���:
� ��Vf�/���"O>���ƹ6I���@I���"O�XQg�X�m_���b�(2:�"OJ�0%���h�~q'��v�*�i%"O�1b�k�"|��D��KPd��K�"O��*�:4B��i�8'��-Q"O���`���`�N,;��Z��P�e"O�9��i�-L�8��ij����"Ob��`EȦ�Դ��@H%Q�~\{R"O~�
^������D�b�z���O�<�gE[�!��Y��+�1~�  wa�s�<��,��`i��|[2P��Pp�<��N?ڶl�E��%3������We�<Y��͕Uyu���#ng�is��]�<�`�U,��"m��?>t-1
�[�<���~�^0 �)��X
2D��GKn�<�ǅ�?v�-�a���O| xYe�O�<��∞I���c��-~t�����N�<��jY!b\N�"$a�q�Z�����b�<iaEA�C7��I��҂�D���b�<�a�f/
,05�тE�>�HIRS�<Y��[�q�\}�N$8�h�%PP�<�@�G�@��#�:=�N$����S�<�C��U�
�Q�C�/�H=zjQ�<��Ob^��j0sEZ�!�w�<i�k�'_M6�@�E&_X��c�o�<c��[�ԅ���#�D�R)W�<�Х��2��d���+�
9��~�<�a��p��0c��,)���.|�<U�N=/�q
d�	�c|xJP�HO�<Ied�s����)�OEh�K�-EJ�<�!">3�u)�&
9!B��d�E�<1�g�89)�d��Ʉ^���6A�<7GƚPB6�a���6�����	g�<q�$�z���SU��T:�!���a�<9�h�{�p$J?��q�\�<��O,_�~u2�A�ww|h�b��[�<�	l'���k�!fz�E.�M�<� j����[:� �(ļo-Mx�"O�h��@_�Sa�t����J�V�C�"O��Ҥd��bG�X��'{B@g"O~��b�&��責� Ru2 S�"O��r3i��Bj�qv��	j�Di�"O,ܛ��!\��p�㌀:7>MQ%"Or�+��]��#�]�rEr�Jf"O�,d�;:�d�c���9:���hs"O����I<@�,�Y���Ue*�"O�!�@�*kցi���K�R�"OX踵*���-�'V"%7��R"O��CϏ?py �j#�܏C6 ��"O܀�diE�iҸ�µ*%�<� "Oؙ;���~'2��3]�Z�<L:�"O�7��{k8�ÅG7�H�P�"OhiزF�*+u�e��q�0���"O腢�M3%$ ��DB������"O��ҧY����C���	�"O$	���*���% �)��y8v"O�)�¡�F|�4c�1�2�"O��Qʅ�0Q�`{�![��"�r"OZx��/H�A��9�G ߳`��y�"O�U��Q�R� D:2i�z����"O0A	�+�J(�h�� fBXa"O�UA5e	Vw̼z"�H����5"O9rsI*2R�q�>}3j�в"OT�g1���c��4ZF��"O�,۠��8J�8����9�"O���F <Z���4职u�`z�"O�i1�OV>d�0iX6�t��"O��W=uS줠@��h��t"O�ڦT�U����V��o�����"O�%��oW�q(ʰ��#T20v�J�"O.��`�4��%z�" $�� �"Ov��Gh�����`�	��A�"OBMɤ�Y	6L������{�np@"O ��WaT<R�K&1}	�u"OR0��  Vq�Z�^�c�̜��"O����!�47{�1���TXe��"O�D"N��}BQ��*S<��""O�- ���0�ָQR�?pHn9��"Or����_�����	+\��y��"O誐c���
!Z�N�e̐���"O@@��
A�Q�Ш�l��@�#�"Od9�G����IR�������ر"O��w<��%�*��L{�"O"I���.�������dɺl�"Oh��e��/+��ɔޕ;����Q"OF�#�W�db�
)A�Щy�"O&ȹ�V+�ye��D��1"O�x��N�dy�A"�b�g��أ"Oz9wO��Q�H�t�K5{��ɓ"O�Dx�OB,)�l�q�@@�|w�@j&"O
�H7�.dr�Ф�P[��@"O�{�?8T4���J4��z�"O2���Ё=4�P��-�ʁ$�yH<q�&�-x�r)���J*��c#�K�<W���Ll@�q�^�Ͼ�w)�G�<���7r7���$�	�5�.�K$�D̓�hO1��	��A�7�TAI�O�^�������8�w-�$:��x�aƄ5_z4���n�8��9ze�m�Y�1�~h��2�v!�gj�;�����i�K{ 	
�'��7M����Q�,L�C=z��f"O� $�D٣���:҉U��0�@"O��+� =.�(��*J$+�V�y���r�����1}Z��C_��-��g�!}Y���++��yÅ��=M� m�V�4�b�|��I�n�p]�b"�LͱG��4sX��d"��c�tA�R�ޞ��H gG�+�C�Ai(@8ch�L|P;^���b�'��' n���Ꝁ2���p%״I�p��ON6m?�Od	��N_5T��a�����(�[��Of�'$�S�3}���;;�J�EE"T���fP"�y��: `҉��f�!d	T�{��X�F��Ob��3T���k0E�8d�Բ�GД5��ȓ�h��E���$92�!A�%4C,�'ў"|�Ҭߘ,N��(1 ��i�q��@�<���FvB�b�)�(d[�#EPwy�4OX7m4LO��V��8=�m�τ%%��q��''�-`�hf��%��Ɛ7�p|�S%4Q|��"O@]�T �!>�F!�o�6qJ�H3�'l�O����J3t"�	�EΎa7�IW"O �j�� e�ma��I�.��6"Or���UP��9�*Aw� L��"Of�kB�S�!7�4��n�0u�l�����tx����]�.tKG��հ���&D�x2l��]۪�jG۷n�N��w�'D��Bg�\����&� ($�h'��O�6-?�O��9/R�/��ǨQ	P�j%Ht�'�J#�O�%;JŜ*鎩@��_;`��?O��=E���E�L߬��g)ƗW�Ba�a���y" B�k�:ytlD�R�"���ȁ��D4�O��Sq�ۀjn�����zT�����x�O���A�|���NU���d����"��x��Z0E'h�	�L��G���RW��p=��}R�R�r��M��F9L��D��h���O�70�2��y���Su]�(�0*�$*)�)͓�hO?A�a��o1: ��eM?Ym2��e���O�ҧh���c�+6}N�l�D�	��������<1�	��D *��@(�ºuPe�Sy��7,O�=�'g�Y���ѓv @H@����M�q�4�OD6�_�k�`���/�$��e1�oֺ1*az���G�s�4�SDi$�H	*��0!�d�U��r���:!�����O-��	�q���(�EڜS�v-�vC;ib���hOq�"��[�
h��H������A�^b�!�dÓ�ȣ�!Nr���2��ʊw�!�$�5/{rmi�M_�N���%AX�Kp!�Y �����Ci����a)�az"�đ�:�x� ���^Lz�sE��	9�!��'~�"��3G�>��ڭ�1O2�	e�ŞU�,� V
^<�p�"ҥ_�[u���O0�=���=WԤ ��'nR9��LC�<��C2Z�*���)_%J��-Xv
@C�<	�h_1�Y��h��w3����FH}��'V:�h�Ԑ��H���P��a����se����zH�!u�c��?D�T�o�	�����k6Ʃh�
>D�$����#ҮPJ�g�Kg�\2�hO?�dׯz�*V�$ҡ&�n��	�'����]$d���m,wz@�@a."D��
3%�W�Fa�T��x�nL���$D� "�D]8\�����I�dlp�� D��zRO�&c���S�;gn���#?��MS�����O �S�G�s� ���:бOR��I�,����ɑ#^�r���m�1Oě��)����3&�-J��Ab����q'L6D�� �l•�H����b뀤P@t�����{�O�xaTE�Z,]y�g   ܭ@����D�=/~N�h$LU#	'�%�R�*���F���(
[
X`����ye�x��Å�hOv�'�����wIJ��1a��]&iT�%ˀ"O���%L�"�`h�p�K2�z0YpU�����اH�:����`�V���JL!�>qJ!�|��'�-���2�<���ΓҨ��@(7�#�O�a�@J�6A�E�9{ˢ-��"OJ<��̅8?���z��	:H~��"O�Y@b�Y��84�3�&
�5K#"O�<jǉeb��D�[�P��H�P"O��z�� �A �q�5�՛�(Mۥ"O�� I�?}�8��N��f������bx�����^/+u���܍Q��H�m:?ɩOX�>Q�O�us�ʌ
�̂�פ(8��A�'�d�- |E��Ü�ɨ�q�Ά8jnɅƓ��i���)bL���V-1J|�r��p���m�&ذ�W�25�m���hO�>	�U��Wx�'	F�!'q��<D���O,z��( ��Dpc*;}��'��`�ӨI���4�C�#1N��
���	7k�ҹٳ �J�X�W(<��B��$s3ܥ
��ıQ�l���P�$bT�ƓsGlP���_��-�')){B����ڟ��=�w�{{���2J��\t@9�����<����/z��`fޒ40&�;eN��mH��pD{J?]2��:b�29���	�(�3�:D��SȖ�%�D��0��]"-�U�=D����%��Gߘ���
:-n�Q�B<D��)w V| Le���6Nn
)"qC�Olc��E{ʟ���ЩR�d"�ѶDѵk.�2"O�ȋ�d�/y����@ɘT�y�"O�$Qu�K���S����&Rnq��"O��1QĝNټ�	&�E-a8��Z�>O���$��b24`ˑlՈ#�IH�HʾB�!��ZP����9z�^���-
�>�!��OЀ�"T,n&��l�'$E�"O���&� *F�C �L�|(P�'��|�	�nﲘ���O�]E����9e���hO�>�AP�Y�u�08*�"3gը�: (}\��'��?A�fjʛ^������0ˎ�%'�d=�O�-����&z��eh�˦]	01Y�|��'iz   ��w�Ƞ1 @�${�� �'�~���cr$!�oC�r~�)�O���g؞���EI�\�L�g�]�l�d @,7���'rq�84cP���b�����Q}�X�1"O�(�E��"��3.ՠq?^ �e�|BH9�	|�'E���	��
5�U��P"R�^݅ʓ/��Z0���qZ�ɶ���B�/7��� nE'N)#b��ZJ�B�	�ة�7��T|���C�J;1�FB� T����-��� �+[�O �B�3vjT���'qOv�@шU�s��B�?7� ��QhJT�b9��F�\~�B�	SWʘB�T��4��ʂ�ubC�I�] a:㬄�A� �m�]:B�ax80V�G'U���,��O�C�ɩ|01JUA@�W'�8���XC�I�'���kA9{#|�W�M�y%�C�I�*r����xXLt��f�w��C�I�F2T���4��s��͊yi�C�	+g99D�<I����)@+�C䉊JȀL�٤lLF �#�]�
�B�)� �P2J�,��_1 4�"O�M	�m������ ;N�.�{"O0��@����	�􄚀n�h�2�"O�1IF枉Om����D#m:�AU"O���HA>f��1��"�D}Pp�"O���Z5R@�Y9��5Og�[a"On �6H3f;f���F��<[��"O5���.�n[sC�!`W�l$"Oй��m�2�&�1�>e�Θ�"OJ�0"��.Q�Х´v�d	��"O8C׉Hiz$ U�V�
H�"Oe�L�H�`�ACB@˂U�T"O����Z�j�4�s��!�T"O��r�ǟ#%�u�f.e����"OD	xc �1vZ>yX �8�@��"O��7%Z!n^�2j�t��JT"O�;���>��ʑBP�H�<%K"OV|[�-��gt5���<M�J=�""OR��
�Ґ���@�8�=�"O�	�$���5*�:>��M:�'��$���b�Z�j��X%-P�'��@P�I�B�����E��=`�uY
�'|��!K�
[ڊi����2,� Q�'�����cUm<�����(�^���'b�)1Ws���g��=�V�P�'�
�㑬�'0�݋֮��I����	�'[�5��`��" �6�̍B���'>x���>s,(����<f� �'�T����D�(lcEX=�Ի�'���a���Dx���N�K��(�'����Hݫ&��-e|A���]�<Q�o[�� U��ʓ
B���W.
Q�<aD�ѤD2��۴dϛ,:��yÏQ�<�҄�=׼�"d���@ �aDAK�<)�*�	�\Q�c�ţ	n�0A�H�l�<y%)��hC���fO�9X�H�gC�<�7��M�����(�I|���ř|�<�EOX�@G�Ehc��3z�͋�B D�<���S:#��쪶���1A9Y)T�L8$��0-���'��L�.��Ӂ0D�Lx�Lx�Щ����~�%(��,D��P��Y.''Μ*u	Q�v���Ul&D��c��ܳ@�֡���0�)�W�1D����3;:L�!�a�m j��ׄ.D���b�Ѯo��Qc.I7Jp��y�� D��P�!CkR�!� 	S��
31D�li��I�;�|8łУ,Bp�ۥM$D��.3"��ܡe-�!�>��!D�lk�K�!Т�*@OVa]�ʷ�9D�t2�e�7�Ըr�數-�L��2�5D�l���R2�+6�U�[H>D(D��I�FI8l����1EG�a��i0D�(�d���K.0��+0�ƙ�E�+D�`�A�����Pu	��t��X5D��z�j��z�pРäSd��he� D�(�0`8f���3��/�heA��0D��Q%mA�aQʌ��=Z�p!'�;D���&߲�N���C,p���-=D���#K;p@�a��(F�4�İ��;D� �q*��z ����<�Vz�3D�S΀�V ) 
�3w���>D��
H�.)@�"�jB+vZ�$b(D�D�@K׷&U��3��ߜA��D�:D�()�+E�JpC!��!V��{e8D�� ��$%��@�����gDD`[�"Ol��1��%�ژx�o�=}�Jg"O*���FʅrX��&�p� �"O�j#d��p���K�T�>���"O��1�T��!I�1"�b#"O,�[��G)W�\�H� � ��D�"O���gŉ�}q��5�9B4
O�7-�n��j�U:84~��q�H�*�!�D>��L��-�$z�&��wԟ0�!��aV�rԉN 6�n��0b]��!���~G0��ũɦ]�`��*��qO��=%?bΖ}k�!*!C*L�"v�<9�]V�UxU�������P"
A�@��W��z#"^�~���a�f�n��0�L5[�@�7����3�6���I	*��TH2"��Eb0�!��$� &D�pr�R��*t(1c�?IjD�e�0D�H�LƈR�HI���S
����--D�)��W�P�S8L�T���(D����#��ALF]��2-Y>lRvM'D�XjFn��9[�R :[��!qGL%D��q��P:J�`I��+R��M�3+?���t@r�-�8����2�6Je�'z�I�hU�eQ1N�W9J]1� %^듙hO�>�s�@��*��EiS3K�9�wg5D�1�m��Z���H�	c
m�3D��Iv�Ҁf����B'��u��O
�O��S�O�܁�CQ?s��5Zd�Q�>i��(0"O
�FbJu���IMU��QZ�܇�	�]�b��pf�S�ġ��@C䉶~Ք� �D9f͊�D*��@^���hO>��.K���끁K���Q�?D�h��ؚ:���(���$cj�P��K<?1�6X����5��)Q��
.�2�������F3+�8��f�p��!�[�a�!�ɍ*P5� �9.3�(��b�/Ǒ�L`$�ӈ(�V�k����u�'���B�`�=!	çR��D)r��������^n�F{��O�NX��!хOF����Zل�k����'���Y��*�@Li>�r$Y6M$�#�3D��hӫN02�h�p�\���l�����ԇ�I�9&P���=�����f�6ja}B�x��ҁe��a�c\�<����w,Y��yr��#=Ƹ���� )���)��Ol"��L'QE"5c�!]#j���J�Tz?�H>�,O1��I)�(��:!#�M�#�є/��IN��h�j��gˍ2�j�z���)�j-*F"O���Q�YP�٣#��oa�!�鉀��	C�OH-� �{6l�!uJ��,I,t��'bt�b��×X�Zp	�bZ�8���ܴ�hO?7mN5���#�f�p'(�Q�ԙb�!�$�5i!,@ѧ�z`�������p?�Ā�!K�!y&�?^����Ux�px)O)�e�+Xx@y��8���""OXt[��,Ne��`�*9������I�HO�S!��(z��= nE:Q�P�VC�Ik�$�&��N]%�̇4�J7My�h�>E�ܴv�bԡ@/��w�����xJ��E|r=Ox#}�	dl։�V��&Bt:�!6��<�����>�E�Ό�J�X7�ϼi�*1�]R��M���O���¦·}q�}�i�/� ���,<OJ��sF��5���kp�]�NC�t#5�D;\O
x*��&h��Bƌ�\-	DF-�k�9LYr`T�VZpL��k�y
� ��d晇4L<����T�j���Y�"O�]�t�F+I@Г�ɔ������"Ob�0��W�\��{��_ar �"Ox	Q�[A��P��;����	~x���N�Uh���E�u����2�	Bx�X��a�+�l-� ʔ%�,�HR�=����2��+?0x�l|��|�wJ�)'�L�
�'�����<5��lӆ��%tJm�
�'-��S�a���%k��Q-$�+�$���d�'(ɧ���T�V���4�ܹA�L-�q����!�A�a�Z�!�)ݟ`���X��Z�H��|����D�P�;F�%x����0�r�E5�(�OޭP3�ϧ8F�x�E֘YvL6"O�!�P��?v����p�5�>=�F�'��O�4��-@�h|��e�)�2�IW�'�qO&���X>E� r/	e� ��$=�ŞԪ`�t�%��*�"�=|,���=y3�)��Y>ƶYѯ��:C�+�;N�!����!$����*��Q���I����Âw���Ф�ΎL�\C�ɇ�(�:��&�(IV�Lob���q�8G{���N�XEz� ��܂������{��dP�O[`i"�� 3�L��c�>#�1OԢ=�J>Afm�0'�����ARG�,=�$Na�<�AOܤ(`�c�l��A>�}�TR]�<A1�(9.�h����<��\����'��q{UFP�Y�z�Rd@B�L��t�	�'�Xv�N��FA����'�5����5I��m�B�	2Ą����'X�\����Y�|�Q��z�j(��'{�E0�)OSz�cQ�k�Ԑ���d>�S�4(I�6لe�P"P��0i��@��y��ޑVٜ,`C�7u�\����J�&�=E��o�><)�bZ3v��! ��ըZ��Q�ȓd�L9 �eg�<��&ɮ�֑�'1p���O��S�?9�Ot����&��Q�g��'S4�%
��yg�SR�q9�Λs����K�	Ry����3�	&�as�敔bJ�Yc��dn��į>�O��@��)�ph�RRo��Q�"OR�k�MT+$ܜ�����1(���a�"O�	�G+��w.<�2�Y�t�h�"Onx��ͺ|f$s @�����>�y2�ޝd�@�k�%¢pX4�pV�3��OH��n�O:QYFL?X�vZF���K�b�	�'IN�җ�qo��dH��?����'(h"=E�t/�D�`�e֭EjD*�a����zX����#�*=�p-�DP�H:HHÓ�:�� �hO1�t��Q��6#6����)Ήu�-��'��d		c[t��\5e~�2����!��o2^��V�A���<0�fG d5!�P'P3RPi�L�v(�p:���)�!�d"=�	���TD�q�դݭ'�!�$"*����O(oHp„%!�!�$ɒ	��T�1B�CH�Y�w�+M�!��	~�=�� ϳ�@|��c7"(!�ܧw�t�8�#����Y#�l�"��,�O��pm�,j |sb�@���E�P"O�0S��M�%i�8IG�Y�D�f$  "O~͡�."h��`ҳ��W�\Y��"O��Q$�	+�P��[�JT�"O�I8T'N!<Dl������26"Oj�a��G�X�p]r�`I�T�	�"O�T�Pƕ�O`��Ů�y��,!�R,�yA��{��8�ݏ?�!�� � ��$�x���bz<!�"OB\����'>4�I��R���A"O�E#ƪ^4l~�S�ڝ��"OPX
&�Yp��aI�	�8��9R"O0Ub��$R�<j��E��J��"O��"��͘'L��BAJ�9ή���"O���|F�uaÍ�m�DA;�"O�q���=�r���nT!!��"Ol̂�&U*M�o�!��D�E"O�p���H#�X��]8�e�"O8�I6k�3,�1���Q�|���"OЈzb_=+�(�Ł2-j��+%"O汙A�[��� �6E[�-r�"OJ ���̑.��1p"�/Lj}�"O�ih�'�f�h�Sk��wE��c"O�	ZCL�X�<���L0'(��"O�IK�b�'wV��!Rb�){4��p"O��BSd�B�xQ�A�
-,[�"O�<�t���5H���@L�
���"O�x����3���S�B"F �R"O���,PܕQ�/V��r"O��ŅC�.����aNL�v���"Oh4��F�+�P��5��p�0��"O,���@�)9���v��,pd�"%"Of]���D=��e!�얬U8��#"O80���h�d �+�m=l�{�"OL��vAX )�B )P�	�pǦ}��"O60Ђ�	�P����ڟue�!�Տb	:�bE�q�bd�95��y�OW���e���6(h\�y�5�H$*1�\T`���/��yh�K��ȸ�$�F�E`��E��y���^���("��$��ـ P'�y��ѕZcT݂�錠J��j�̆(�yR�Z9E	y�`�;VMQ�+���y2·�?��ۀ��EEE�׏�y��>?��0���.�P��tØ�y�"ξ=����s]mӠI
=�yҦO�6�����e�������ꜱ�y2��$O ��B��&��ȫ$Y/�y��9z�D#C"S4'j�ِ�)Ǔ�y��$|�K`-�9%t,\���7�y�E��Y[䢆�5ܭ����y�@�>Q�0z���xތ��SoB'�y�Q�H�I��G�z�ZqR���y�#T�h[��j�Ψ"���K��y&�D�Y� +�<��.I%�yB,L>u5f��µ_�Ȱ�g�J��y�G��n����p��-T�~������y�k�
Lbƀs��αf�Z�;��@��y���Q\Y2T���_��x��*M��ybbվ�x�C�M��8�J_��yRk�!W�u@`U.T���T�y�G�Fh�uj��2B���[U Q�y��
�b�0�	 벙 �N��yB�͢0��;7c^'���ia��y"fB0jDV�HͲ2ѱ�<�yBf�>S�^v��q�t���D�5�yg�%b�
s�fM:F�q�Ї���y¾Y-\X��!�c"�Q�+C�yR�Ǣ6RRI�CKV$	�6�'D��y򢎐o�,��͗�i��y��S��y�O2I?��+�ʜ�e�ح�7!� �y2dۂa��m�'���X���Q
Ѿ�y�![�Z�yg/HXn0�!��=�y
� @���4/����1C8��#�"O��$Jͩx��q3��J54k�Y %"O^<�r�]D�	��O��l��*a"O>��CV���`:8�b"O���gX'bn �8�N\�|�p� �"Or��0M�|d(Lq�M� �����"O<�P�S.+bN�0����8r"O���2.�y�8@R#dĤ{@���D"On��"�R�p<���%[��<�"O�Ñ,s��\�`d]�#aTQ��'�� �)��=�����(Z�r�F�( ���.�R`��
O4�0"會/2`Hᕨ��AL*mc%��"f�-�r��_�1���1�OӋH��L�!���`Dt�"O��w�J�H���R
 -�j��4;O����
)������<E�t��
����K=���Eg��y�I�1+g��aW���Ǵx��d޹)���Xr4�BMR�}��g�'�,��%BO�n�4yS���)@e�"
�3�V9	�)],�pM
2��5#G<���Ƅ-�<��ꗥ��?!ED�1r�p�[��O=#��� A��H�'���a�N-r��G���G��;�.L+�B�<#i��@�Ώ��y�.zp���H���pL �y"�.%��aK������)�f�ab%˖l� �����P��A�ȓu�P��0�U�V.U
gk� Kz�J/O^� �i�4	8�	D�?#<�F �y�Ё�W�5Wl�K
�n�� U��9�8�$� �C��4�p`��U�M�ԉ��əq�P��p枻B�pM��8E�$�>��Ub�$(7�;��Ũ�XbL-[d� e�$C�	�W�X�!��L3.�I՘9���1^h�Q).��S�O�LtۣJ��G�FmI����K}�yB�:+<�"���Tv=�b��y��ԀXY�F�B�:����y2�.Y]����h)�:�ir��y��(m�L�q�O78�}#�CA*�0>�Q�o�~'�;M��$�"C	�	k6�Ƞ���ybg�q���	�.���M��'ad�a�? �?��F"A8*�����Up���XC�'D���W���l5��2���=4@I`�n�|�Ƶ�#�l��]F����\\d����4�����͋,!�DB ]@Hª�lmf��R�P#CU�& �	CL���-Ml��,X5�Y(#:p0�C�B��q&�*�_���lΕ��0��'>���ऎbu�$��=�j��7�
8#�b�2�i�
PR�B�#fH�=2��>�,�ЕD>
 J0j�Ĝ�Qe����]If�ې cO�5�O�����DȼC �Z�V��S��p�,��K<I ځU�(i`Q!=o�HK$�13�PX��-����5F`���AV�&qHq�����'a�\�D����і!؞R����9
%&��'��D]�H+�H�1�:����~�:A���No%��z�P̃B�%�PH#	�����-E�X������%-��'(��"�1 �1A!G�U���ڶ�Og�@���pDl�(��pi�+Ɉ+%�M��)R� B�	�z�@�y��˟nBY�q&� v�7N�p$���֡m4�Y�g@�x�B맏y���=�nK:v��|��E������g';gaBG�q�(ex�'��"u��XDO�3,?r4�QA'�#!s��8�N�.=���;s���$�
0�ZB'�dPe*�B�&9v�����j�VP�`�Ә ��sŅ�h����ފ4Qԕ	�� �4�����'���F�y Z�R3a��5Nd� �'n�`�w�T)3�h�F	�� 3��V�O@d�R�n#64<�A �*)	����'��@ "Ɖ�J�Ă|�r���^-7��Y��̈́H/@x��l�~&��Oh"@�>�$�ĕS���R'	�F~X��}8�|�Qi5�.�E��T�*+[�6�a1�	K�ι�W�b���1&���{"���t�v:@ ����t�V��O��2��̞�@� $��1����"�Q�|QV�E.� (!"O<��e=7;l8bf� e�j4Ц���	[��33Ç�e�H@���4'�C�W�v��`�T��#�!�)C�������}b88��L�i���Ⱦh<m����nlʄ�f�'6��h��R  ����(!�p�ߓ9��˂�̅}=��(	� �=ڵ�Ҍ�-�ALZZf���ϟ"\ڛ��'?` K��&ZEi�V�7J�D��&�+�j�hF��H��(�ƿi��'9@�)k��2S� ��ᗘ��5��
�E��G�
E8�����^�}�
ջp�Y�q��8D�{}�m��h��Ĝ�	U��@��u�	���%�!�D�6��O�<D�p[#E�8.0�恆0��!`P'��kd�40�E�Q����L�$�:�`E$f����)��=�1�S M������1(,��I@gȇ,F��P��wT�D��[�M����� �d���LI7-�����?9���:��C�NȐDx!��4��S�<���Z)��	��*��{��C�I*yx��*ᄙ% ��A ��{���ǇN�B�iRb��q�B�1��<���Y�b34T�eM��a�reaYB�<��E@&vN8:v�X ��t�cC�<ig��"`�92p( ?4��$�+k+YPT�E�Lr&ea��5!]�|���ޜDiE*��@�L�g(����QF� v��DOV����Nm8� �Y.'t��	�-H�Quݦ4�����J\0<X�B�ĺAb�S"O"�	���]��=��Ŋ""��c��i�U����$�D��O?7�@�ki�|Y�%�7SŎ��	�/,!��"�
(��\�s�
��^�$��ɧr��5t��F��`���*Y�
ͻ��
���*�)�Oz��D�d�Jsc$������R�Gs"O�0��ő��L��A�r8Ό�2"O�\#SMش+���s���i���7"O� �S���$��B�SC�N��"O���Q��V�Zf��2)��г"O �� o��^�*dj���u��P�"OL����14���:$^.0�p3u"O���Ќ��{���aD��N��&"O�����>l���:M��v5�A��"O� RJ�cX��'�#��!Y$"O*�"voV�^;␡u����x�"O����LP�$��,��m�oyX�y�"O��S	B��V��������09W�'
�3��-�3�d7T>�d@�O(�^�����)s����[�,v�0P�;!z �2ο/��c��ǉ���0�'7\�S��O+�>}�B�UY`p+
Ǔ?����I�;R?Nh�'?����X�"���+	��M�	�'�(��U���1	�1��V<��� I�[R��?r��1"6�'o�L���'L�A�l:īɞI�@B�	 �����;�N��D�8�ȡ��~bi\�t=4�}&�$PU#��|6Uʃ-�J`i��,����@�^�(eh�I������\�͸� 	�S������F��Q�Łjf2"t��H^ay�fK���x�6?9�K�<B�1q���*�ٳҬ�I�<i���k� �#��<�n̻���\�I�=�h����2�)�S��Z���I�_I�l�ck9*:C�	�a�Hra�=ld���N�22�B�	�j�~�h��	M�����>Y�B䉒>J����Ϸf=r=��mZ3)�C� �h���S174x�	�!�6��C�ɫ���eO(i�R
"mK�C��CfĐrs鈔��u���H�WcdC�I�7�@;�L�7ߦ�-F�u+�C�	x�L��ԝE3@ ��d#��C�I�i�&��l͡&�,pS�#���C�Ɂ1V�`��:SFD��FKl�C�I���ٛ�kÓ)b��k'��Qt�C�	�2���@\s���Y��\('�B�I#kO���S"�,E��qJ�A�5B��B�7u?��'�C <���ۢ��a��)D��:���*N(ʍ�'�Z�E�Q%D�D����]"�u�ƁX
�q� �,D��*�m��`��C"MV����F
+D�� �I{BbJ1br�� ��5l��!��"Oj	+3�^�HD������<��"Oh����3A~<�tصU��)�w"O6�:�E�	��<�A�Z��"�z1"O�m�����:`�nj-�"O^�y ��8j�<=�T���ҝۤ"O����E#Lv���/N�4P�`"O.T�Ô���|���f�(�D"OBb�ϴji���%Ơ� P��"O�D���ݰm��I�CIFh���"O$����@�
������Soh���"O�����+h$ؕ��AH�IT60*b"O��i��( �A����5^`h��"O�[4�F�@)�-[DN�b���"OB����fF,��T��=h3"O�i�E+�)'D��ЕL��^xJ� �"O�qz��V/�4 �wM��e�h�"OR]i$M�3��t�gR�w�D�"O���D-T�<?J�	�Fo�%�1"O���a�@� � 0B5C��#v"O X#�-� 61�}k��JB�v"O�Ph�'P�	q���/ѓ�"O��Q!�v_�T���G~�"Of�����\t#�.�Q]�Y{�"O<�#�ūy�~4JSbQ>27�@�c"OT�
u���V�,�q�!�6���B"O�}���x������!�&�� "O�Lzv`S�%y��W��q�!"O���EaC֖}{�	<ŐLH�"OZ���.�z�4af�׸>���Ka"O�ͫw��,�v$�ҁA$B�����"O��:Gd��]���ɣ.ҚU���б"ON�
�e�I���Y�K��d�PY�"O��0DFV�@eˆ*�J��IIW"ObUR ��.L�4��IςLr8��"O���ȵ `)�I�7R�Z�"O��J���-X�E���p��M�R"OI#b#F�:}�yb)J�H,9#�"OH�8RⅩi�T�C�� 6���"O:��d�>b�@���(Q�l� "O ��̈́,
�Z`�'�G	m���"OF���\�[�<��w����4�V"O(|��f�E��hP��ѥ�J�;�"O���"� v�D	�a$L�-�p���"Ob��ԯS���!�b��G�ҨP�"OpP2b�L>s�8��Y;�衑�"O������*mn��Oɹ�Z�
�"O]�f���N̓��P=6�|	t"O��A��Tbvl�@M_ M��"O���DBD�g�~�lÇR�F"O(�� �?d7���l���"O8l;�G\1�<�2�����& y�"O"���/�;C��M��`�:N���k"Ope���Qh�l���R
k�8�p�"O���%G��Y[���7L��w��Ac"O�B�b['~  �I׈a��P��"O|�H����` α��ʀ� ���x�"ON ��-^�<��Xa�@J "O� x����<�#'K<>c�q�"O�%�pl��!er�AG�%��� "ObY�p$ԑE�����V�x��C4"O�x;c�L>��i�EV�O�p�)w"O���ai֚u5���f��.�qS"O|H��ȋx]�>.��M��"O� l�2�'2p} #�A�h���"O>�� ��5,P�3�͐��5 4"Oج�@ݓv�l)����=�N��"O�	P4�-zT6 �'���@�5"O4����.`dX� ឰ~�R�s4"O��3����1VR������ղ�"O�����)"1�mCE�X�� ��"O��ڄn �~g�a��ۄ\�4�;�"O�D�&�ɦ@6�;��(�p 3�"O�y�p���-Iޜ+��.��l�v"O0I�♗93��B�̞�w�(��"O1"UD_L���'���6=.��%"O.�DڣX?�A���:2͈r"O���"�%7n�ͳ�烰"�
��' |!����$*&�)�jK g���3i[�mn2A�r
O:���"SԂd�%5l��L#3�I�=(8���HXC1��aC�O
Z� �򲊃(��l�"O��k��k�QZ�C�<g�9)�3O�`R���$f:z�[���<E�D�]8l`�Y�b��`\%:7��y�J�'�4�q�a��{��D�剆C6H�#��6�g�'��ؐ��T`C�qi���78���+�C��ivG�/u�YЏ֑t����a`��-�M1�KQ���?Y_�T�Єn���Q#�Z'A��{����=J���\�)c�|�*d�ZM�L)��H�7!�B䉁r��Q�PÕ�~HT}[�AH(;Uf�5	2H��G�ԴP�������fM�^��1��Ϲr�R9Y""O4Aa6<�
��$�;�r����<9$[�%���1��z���[r���P��#���6�O��a~�gm�̌&+�r*X�rL��z���  �H�i�Ny1��'`���t	vGZ�ڷǃ'2N|���d�OBz�H'$�.��O�\�+� �:~8�2�9)w8�x�'nֹ3p�])��Plş#>Έ:�O��Z1�͇c)��O�>a����G|�v��8G֠��+D���J3B���R��\'���أ�4D�@$ƀ�uR�3B]�erV�*h?D��r� M�Y���QPjT3U�Й�7�?D���BC�Iԁ���J����D'�O�X���~��MCPx}bf��N�����"��y"@�%��ј�E@
p}Dђ�E
)��'ӺX	���J?��B�#���à]��l���!D����Q�In<��Ѷb�X9� Z�L٪$��C��t���DL�L��LY����;~	"�Dָ
�!�˛S<~q���݈thHQS A�:�V
G.J�D�[�i�����P%\!��k� s��� %?�DW�@���!�>{����'�Lb'��W����ur��k5k��(P�@V6��C��9AѺ�ˇm�*V�k�Tgjz�4->~�.���6�L�	6��:Dְ��Ol$����M�Àfߏz��ST�˲s�x�r��Li<ɠ�_Gsr��Pf�N���F�_O�Pr�GV25�
�H�	D-�h�$M�Dt|3�KЎ��'�X���,#'��Y���',�L������F��<
gԓ)��@b��.Tk~}Y1lğ-�0a�W��'Ud��\~��D�)�$I�7b�p�� Pc���;�o�'�Y�1�>!�]�a�t(�Z���W"��ʗ��D�"��(���]����#t&Y����F|��4"Oxi���;S����a��D[lT�cN�5�0�ۓ�Z����?�hy�_?�̓(:��a�w���� ˊ�v,� �H�%`&��	��?=49;1�S&yp�+�F�7R��,{�#W�,; ]���ab�ICEϋ��~���9?�	Gy"�O�-�Ɓ�3KP�z��yK1"�0��O�y����_���#�[���#�gߖ"��}C���$'��Ш�Y�ȓ�D�B�KJ�48Sc*����'].s��aeI��sKd� T��3^Q>�zR�� Dġu��/�ҌТ2D��	ՊֺFTpEr �A,��[���P�`�(�&=��ǎ"tʍi����}R��߲�����:�J��`����?�Q, %�1�����)B�yÕ�4,v3���I�7]k���d@	kͤ	�k�#�){�K�џ0�r��.o�*��|:�!��Y2�0�ł2I�]9���z�<� X�i&C
; �Jx�`х	��
���*�,A�
qO>*T뙆y=�yK4
�n�H`Z��8D��rƦU�.N8z�"����6D��ɶ̆�JNԽB�͍�� �2�6D��iA%L�q���P��R"�I�&D�x�g��6@�Q삝4�-E�&D��!�|��Ec��Y����K"D���4�VQ5�qH�P?�t���|��u��`�qO?�r%A֘C�r	%�S�"���6D�I���@x�"�	t8�ѡ�.�<�
\�:)��ӓ3q�+�Lڔp�����ڎ ��=��ɵC�N�`�����
�eۖYRc�I)\�r1 OxJ&X|k
�(0*�"�|e��ɵr,à,��7��8�Ҕ��6{�"ݱ�)�"`]�҄"O���@Y�Z^�؆�V6U[0��F�i4����(�ZԦO?7�˙Z�=�ᐱ:D��E�xe!�Xg�<U+�ow(U��F�#z���!~<�S��C�6��y��"��$������Z�'�]�ְ>ia���̵Id�]12���lW<!�B8 Җ��B�I�1�����p�M�$�� u#=��h�e����'�ӧR�}I%K�l��D9��݌#�(B�.a��(`��=��PB�N�7�8�a���C��)��5��� ��\a��� ���if�8D� ��ꊢe0V	�V��;n\�J��<Q�(\�\�yӓ �$9)��H"B�r�#�H�	m.����6 |�4��	F������MbQ�!Y�'@�jnC�	�ow����<M�ԉY#J��#�|C�>w��!���E����@�.C�6CmjI�U h+�H钣�	p�VC�	0
J*47�ȥ_�b���I�{��C�ə8Պ�zGOZ�f�K��ѐZ&FC��9(tqFj��lq����� �VC�	�����F���d�u@��b�C�	J���5�D�b��K�����B�l�vD8�B���13�����~C�	��8��oX7 �T0��ό�2,C�	�#�j	s��+<^Ȋ��P&`OC䉜B�`[#)ө%*��8ţϐ��	J&�ć�#(��~&��'�%���C�́6��ꑭ,�����A)k�PT#�%M��DҦ�D3{����腴1Z���$�E\lp�K�9U����	���x�!ͬ|�Z͂�ҥ��$��^Z�q �`G�P�P�:Wu�!�ds��m*Ƭ��r��b��)����Z0��XP�F����2O��3�؉z��%!��y"�U�EK�	��j��it���7�Z76�H]`�����#�6kgq��'�T�P2�Ĵ(��(�EG�iА�
�'�Z4�e��/P�&)��C�̘�q/�_}d�AQⅸ��>Y�ÛXivt-H������UIX���Fʚi����Ox5�5Q��|�{��ƗW�i�"O�M��R�"�$���Z�~	�G�|2와[�v��y��䋘�~op�ҮA�	�P���"�y�S<m�<�d˷uӔy�kC�y�f��7Բc֊���W���y"���'�&���H��|�� � �.�y"��L�n$c$〱G�T�eaN��y"�:����`! 
<H`�o���yR�E�5=T�:�%�� �%B���#�y�kS�F)8)� ��)��Xp�jJ��yB�ջ-	�uAY�9X���z�|9�ȓe%T�Q�*μ: ح+�f�9T?�ȓi?nR/\0��7"I�O⥄�=��$��"-XC�*�̦8�z���=���ڱm�~�*���/5\|��!Hգ�ƛ ݬ 1B��%B�)� U�.ؚz^�i6dK6~�H$��"O�li�M�>�ΐq�cQg��"�"O0�H�ی_�	���uRQ"O`%z���,Q��8e���N�1"O�U��
�?�Xu{�@U/-��B"O�����efјWmcI�`���y"��J~�Y���(�h3�ƅ�y�*�7aO�5�@��"��%[R���yC5vj0)	3d��l�(|)�fB�y" ܷ<ؐY�u��aP<��Ƈ��y"*�ht��ꦇ��-���ì�y�G	x�.�5�9Q�>����yR���YE��HCC�!Q�:��C-F��Py"�2~��eaW&ՒU<zLIAi�<�#	��.�h��s�ܒ0Ќ9��@�L�<q�f��
Z���"�1��HT�ZK�<9�c��I�N�*��T^�e��ȒG�<�v�C;Q�>�`!8}&�BD@�<!�)V9�Y��6i?0x��b�<���M^a��bP[-_�� �B�Q�<�5K$0Q��%w��q�u��z�<r�8Šc���H�	�cM�^�<�4�I>0�pxD�'!�<�pb��L�<9A���c��m�T�+_X.����J�<��
*[�8J$�C�9=���R�<�͓@�,y���Z�E�=w�B䉎7PM1���2��!�Ǝ�r�hB�IN���"@G�,��ٲ��]�!i`B�I[X�r���Dk%�2Luz�B䉼=��B��>���qV�HZVB�	����Мym�t��	�2���"Or(��6bx���	m����A"O���%�U���Z�(�/
���q""OnU�cCƥswj	[%��_4���"O�U0�%S�(�f�ң,?����"O�����&KFx�b�{��$ S $`@B�E�((��g�o��h�<I��C�"�� �B���NN4��ta�e�˓B/8=��59���'(�d�@%�2
�$UR`�C�X�L���#��bLZ5%V��?E��W�?��U�3X%�H��D�/�\"U���^�~4�Eb˄�~�JP)"a��&C��\���ܞAνhFЂ��U�mA ���W�AKXx���
��s��ד&��'��{��7�)��8s��`�t��Ay�¹S�0��_6���=�	�i跪�!H���n���UL�4Q� �)ҧ������dy2�잍S�>oZ#?���� �?�֝�\=�Q�q+Ȁj�|�r�
�Dy� !����`��%x�����+��q��hd����O��vQ�V�q��aavD�"1�<�1C�>����f���O��=@���"eϘ�%�c��q��'�-s����,S��8��dO�,>�in��o`r�:�(�s���셓�HF�`=���T�`U�Z!�>�	�B�T��ᓿjI�)��+�h<�#*�B�6�'�(|�g�����O��u��e �X�����B� j�p�'
���NN�ɧ��|�O[�,p|�/W�	ya�:�ҷ��8?�7�:��So�	Y��ڑ3����B�>:�����U:�O�?e(28v�� ��D6�d,X�E��'ʾL��Sm�R�sf��x0�!�_:!k�������ا�S����#Ҥ�`wI�95����O�M��)��1v�=��H ��{�m�$?Tk׀��?��>���<�N��h��Uɨ$�J��3�0D�����Gf�e�O��BV�$P��S8=7�����2]h1s2�ЊC���cC�r-{��Vs�?���5��%�OT���[��'D���q��{�����X�+ �̰4�7D�$�5���ZQ��1lA$i���;D�Y���T}i�o٢!� ���m.D�� :�sRi̋i��)g�@@�%"O�I�,��z��8@�.�,<�c#"O�=�C�+q����Kw�"�"O4� ����vx�U+�M5��y8�"Or8㎡cR�1Bʍ'�ݓp"O�a�JV%�����I�/@N~a��"Of�� U�nK>9��h��L� �6"O��Adӓ7i����5P���"O.����=���h�!Q8���d"O���'2 ����f�@����"O�����'ՀEK���|�BA�"O� ���ݵ͎P5�_�P����"O��k�/'w�� �"V�V��v"O��j�Јw���!>���H�"O$ ���W��d˴$^�B�(B�"O
��a�(R�D  �K�<��HqW"O(����ߋr��(��	u��Hu"O�У4�A���c�H�1gdZ���"O���Eo�5,��1sG��(�>�P"Opi%탫�ԡ�UfK<K����"O����.�-�,�*R��Fob\j�"On �kJnL��� ω
x��$@�"O���M��Ob@ap��O:XR��"O<�r��6\��xh�,ީV< �H5"O��2%׭��A��3�r`H�"O�ܻvG����d��݃U��"O��Z�iEl��~�@�X�hJ�#�!��a3O��QY��r@GW��!��=o�4+v��kS��P�gH�!�2x�N���+�16n�P�0�ʨQ�!��_�꘨W�V R��W�!�Y m/�8C��	���B3�L �!���X:�BEoB�%���Q�*��D�!�$Ȣz�l���	�p����Q�p!��^�9�����=P��6FǗc�!��	<w���O V��4�cOJ0N�!�$P0"d� �6�ߗ/��IJ����d�!�$$sb"!�$��'b(����k!��|�����.X8i���c�-_!�䍤T�,AB�!e^�1�bШH!�$@;hi�����IO�zR\�1=!��?s�!�;��o΍,!�d]�2DU0`��v�<8�Nɏ.�!��X(�難/�'�f�)%.?�!��*��z"Y���̊WGM�%�!򤌝H&4�Z�
�R{r���K�!�$)�0u�"捋O��<��a�8�!�䛗�.(T!��W���K�@�Z�!��_;1��5�P�V�X���  p!�S�P~��3t �;X�lZ�c[\!�$��Ob�k"�;�QP�%�uZ!��T��ɉ@,����r�c��!��DgRИ�� 6��Hq�� 7!�DN�$:T�u�C>K�2 (��O3L!��Q�{8L�y2D�5/�=X5(^#Yl!�֘}�=��T�)4�A�&�o�!�$� �ji:㠝 :���%Å+�!�Đphn��1.�	P�20ZG	�]�!���3X��S1oC�����A��8�!�D�$Y2����Ex�hzOV+�!�dQ&.o���
Ɇ.����m���!�D���\cgȋ'}��j�&e!�S�&S�*�
o:�{���=h!�d�=qORh�UK�8�r��E@�

K!�� Ҁ�qj���J�	t�8���"O�!����&pr�\('��k����"O���P"�0!I^ �W�[�4dP�"O�id�o�Be+�$H�\�:�!�"O��Cq�	�\�T�p�D"t"O4L)&D\&�n���@�*�
U"O<7Ɗ���C��'�h��"O�l��?.�e��E��5RA�1"O�jbeG�`��sn���v��"O�lѢ�	�Tq�߾0���Ò"Oz���� D�T�ߞN����"O���ubG�_^�`qҤʎ%�ɁB"O�y` �35w2uy��_!;s�(�"OD�4i��9Jh·$ƀ:�L��"O��Z��F���`v��7޼��"O�Q���%*���ۣ`(��hU"OؐKࠓe�$�ҥm�<�Z	�%"OF[�M��&1.�+��!d�t<s�"OB�aB��j�
����I2I6<�V"O�Ix��G+UT�����C6��}Y"O��B����{o�@A���F�:��t"O�q�\�W*H��
>J���"O�}��e3��Hr%@}�B�(�"OX����V�蠈C���?֝�"O�@��"0�A9 %�w���qW"O����&6��
��z����"O�$��-�&_�������(�`e"O�D)��r�JԂ�L�\R���"ON��
��k��͋�+��s6\l��"O�,�S�=:��i��c� 4�L���"O�j6A@�O0����C�~���"O��T��7$�+3���9���r "O�7�ƛi��p�3J-p�U!p"O�Hs�kN�2}�6�@.v\֬rA"O�!�,Z7=VĘ�ǧ�
*e.�G"Oޤ�Ĉ�~i���G�B�	���"O#2	.y}j݊��({R���W�D{��Ɍ$�l�����=<.����bw!�d��>Ahs�E/_,q`�.�9f!�d@�Y��-�����iˠ�ȵ�V�W^!���4ky�mL�s���ʠ�٪��B�2dej� aK�ݻi�$��B�	�t6�Yه��8_���bw��C�	ZV��kV�o��(�x`�B�	!e1��I&��G���W��,K�B�b�A���)e�Gg�8`��C�x���҃B�X�%��� �C�I�V ؉YSΓ�pg�M�5�L/5'�C��/n
���ۈz�j2�I��C��6���Q�c�d�0%��Ĕ'k�C䉠q�!t��'F`�뢧
S�bC䉂�ք	vL�'sn���"K |C2C�	�9P��x�B��z���H�#�!�B�ɅNpv躓�W�Qԍ�Ph B��.Y��̃R���佛3f(:�C�I�1�|�/E�{��]Y�F�8p�C�I \"hA��ǚ�y,V�
ԅ�6h.lC�2A&�Bw���hX����O� JC�	+.��r�;9t��箌�o�RB�I5Hz���@�	�XD3A�M%x~C�	�Q�|�QP=�Vp�կ��{��C��'��zeH�q,��TnC��C�IahA���_/%F�i�v/�d�C�I#h`���ʵ
Y8�P4b$;B�)� `����*ssS`���ݣ�"OJ��FͅOO򝂗e�;o�xApE"Oi�냍	Fp��D�V��CS"ONȁ �T�Sp�MiTGa:	�ȓ��1G�m�j����Z�@se�ȓ{a�h��E�%8�� �%i�h�N�ȓ\9��ˏR3B�SE�
1n=�ćȓ}߾�`v���%�� Q�J�M��݆ȓCQT�Sb�������ߪY~��!pxx��['A�.lA3��'!�����vae"�8�(�*COy��}D�|X4h��R���k�'\�_�D�ȓ���8Jօ3%�rbNE*8)�p�ȓ*2�!(��H��0A���ux�(��'�z͡@�ѕZP��H3晡'����#$�`3�Á=�v�(���(<e(������X�<Թ�fA_#�ȓ~��s!�J[�8�YG��Mն5��E�T)7�6��4�̤���ȓX�h�3�NS6=�摋h"l���ȓ2N^��Tk[4s�N ���7�*܆�8C
`�f	��rŢ�,� ��{:��㈖08��M���[U D��	.D�.�?%�� ��Њ:xpD�ȓF\(��2�SM�	���N��Y���.��_�8D����"`�t��`Bf,O�R.���A�eY����n/�5��l��P�8A�V�����9p�%)�g�"ip���O�0��g^�8���2BT��&g^`hL�ȓ$9 �*�nN�6eF�������
 ���P� (?�8�$��&M�0�ȓA����'&�5��c�b��x����M�ҝ#WF�X���zaI΋vv�0��`$��vh��(�K��޾p�T����|����A��M�%)L�w1���#3�ęi Q`5㔀�/iZ���ȓ���e׸a���%�Y!F�l�ȓ+�Q{A/�~B�q��L�f����=�P�م��4��a6C�
m�ܩ�ȓ/��IF)�"@>\�J�6��5��J�d�"v(;o��%�
��S��a���b���A�8Ƽq��Y>P��F!Ɓ6I�Q��M>�$x�ȓ!�}���G�2,���F�7��ȓ[$Zd��lN�*�zвV�W1[�~���?�X�hK7H���J�+��ņ�?K$���.�^Q"0rJـ6�p��7g"݈Bdз|��CD*��o���ȓ�X%�q�G;\���Ɛ���#(D�Й�E��'��Q�L["}P��iլ:D����Q��ĜX�hz�A��´t!��ů"F�L�ԌW�~�t2���$!�d���!E��&k���8R`�;�!�G���A	�=��ST�̀F�!�d��0w�dx��4'�(X���Q!���(ϔ����Z�;Z�Sc�
l�!�DX�z��DȥGˬKS������$!�]0H��4�-��D9���?!�_�r�Va�&U0ި��,��.W!򄐷Z2���+M��*�߲t"!�Pp:d!��ʔ�]R��R�!�dQ�	���"�T�5�L(��UM`!�&��,q�JT�)�<��`��<�!�� 4, ��U1yXȢ�oޥgwv]hA��OnY� �*�M��O�'K"f����?Y۴b���ڰU�m��-��ڗc�~x(�)�4��E�T�"젩��,ʟX�dM��+����I��8��t�01��/4��i�#���@6����-=��Ą��?O�h���_H���ѐ?�X�!0N4�S��s�z�"�Dp6M��f��@w�L]m��LE��4q	�)��Q�=�v����ک{�����?I��?.O�"=9���"*4�=�r�P�6s�= �	I�'N�6�����ɻ�M����Xw�����%R�x!&�q�/J�C�^=k#j�<y��ۺ6#���?����?IR��\�'+PA OC�p�T�[S	�-� A�],;�r�x�o�49���1�d�+Q�4ϊ�G���H>a�EϧS����%��y�:��p,�
F6*��2��lJ���K��l<�O��j��'@=��A�OzP��n�')�Bt4�[K@T�C��Bi
�!r�R
&D�������O�(��I�=��QsQ��wPRm*"O� 1ċo��U
�Ē�1ۆD���-�M�F�i��'V���O��	A��Dqī�%	,V�y�`�OH���4gu��۟�����@���d���'�"��GGW�t��$1�I�^����Ԁ��b��Z���S넽q�A�~bL6���i�Q��
�씜��ۀ�^�K��QыA���svd�D�}*���,�ƌ�L@6]/|�bCR;��m�^T���wVXg# �J�yؤ��;;�Č8�ē�?�����'���i�2�8vƅ�sΨU*�܂^ĺ]�I�OJ��d�2�:0#V��;y�´C%M�:mD�����9�޴��$�{T\o��'>� U�_����4�V�:C^��S��@������?���5Yh9g��m�>�7i�'8-�(�g�z���FȎ�ލ�w���*T{D-c�'���"�E��)��C'5�j��g��;$``�b��b���r�DMO��u��%J?*%4�U�|�eJ��?��
\�OQ��nҧҔTIU�F'&2�d��%��D"�)�'����nR<�;�'TtF`��M��ME�|��z��Unͦ�;SN()�>�I�K�?Th}�$�ź%d�v!ͤd7�O���*����?����M`�zW� �c� 9� 0z�lN�`�(��#	�^���@�|�:P���i��D���Ok�V�Ǟaue���@D��	�M�VEԨ�p�$�yT�� 1��8xι���(1X"ϟk��$B�c�(.�B}��pԛ�$A�?A�� S���#|nڸf��)S�� �w~}-.�["�Oh��%ړ��'�|:�` =��Sꐑ�8����榭r�4���b[w�X�rQznT���(�� ϣ<q�f�w산����?A��?Y�����nl���Ę}�B)
���Jc��I� �J02��$�U1{Xm�d�݀o��� M���bJ>��CW���h��G��6́���?��3C��\"�{�������O&�l���Ueh8�Vr� S@k�'VJ�Q ��V4c�Z���>I��B��h޴L�'�b�'��� ����dɄ�=ˤ��TE�2l���퉢WTT:uF\:�.x�+���(�"�i'�6-?���L��7��s�&Tp��  ��   %    �     �+  �7  �B  �K  8X  1a  ug  �m  t  [z  ��  ��  $�  e�  ��  �  )�  k�  ��  �  3�  v�  K�  �  X�  9�  !�  c�  ��  %  � �  G  Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�� |d��"O
`�(�;���8���-0��1%"Oj4��ND^[��"3/9�0|H�"OB���H��*�ʞRy=a"O�味V�!X��!&F�:J�$���"O,��a
���C�Ą�M�"O,$3%o�-���p���+Ն�:1"O��ݢ1����`���y14]2��i�<�6��{_���c�H�`�fX�$Kn�<��A̼VI�xR[�)�Ć�pඤ�ȓA5��('nߡ4�� �)˩%� ���,��r�؊b#`T�eT09���ȓ!�b��g��}�8�F��-? �ȓ
K|m�ș�VṔ���2�%�ȓ"R�X�j�4JN�1�˘X�i����̹	_�jZ��1!g��zܶ��ȓgil,*�J�
j�Ne��i�J%b���f	�(U��:���G��$Y^م�~r�� S�%T"���k\�jx�ȓ|4�1�îJb��@ӵ�ݩn�V��/[`�"�v4�R�!ʎ<��M�ȓ`:��z�ؚh�J�Z��$HY:	��H��p�m�C1��!��B:��0��EnjZA V;9����J[
2���	��4'J�EA�IVW&��~�(aZ��ӹ�>� o�Y�|�ȓ�f�A�
Ο7�H��M�$�����mޠP����/���ANXo*�ȓTv�����{ ��-7�*h��I��sB�8�8���3����ȓNe*M�悡;������X�o��!�ȓ'lj�#F�m�+R&;�|��2)n�C��0S4���T:
b���:�0!��e֊��)��ͷV��,��IJ��5�t�cnE�b��Q�kX�y�}�ȓ;?���Gf���A����C+�Յȓ <���u`�>vqF`�f�Y�k+^��ȓ#���#��\2�߻4�:��?Iӓ2����.�!h聻���Q����SU�D1Qm�.o��)��^����sh 	s�l ң㇜9������X�'���+�ǒ�҆���gL.�&e��'��L��I,0`���ÀڒcD��	�'����Aˁ����Y&O���.Y�
�'���;`�"R}F���+]�YX�W�3�hO?���"��s�(��i8:h��E�ay���s��*1	A�[��U*Bbld* �7D�pjbKۋ@�0x�����ٶ�"�"4��=�SܧNO�0e��S�F����7bq��L6T�q磉��.@s%�D�ZQ���?A���t�A�'h�T[���3�����	+T7��J�'��yУ�	<���&+�:6S�]�dc??�p,.] S‬�x$Ca!�JB���ILy♟�:�f��NL��m� �p�֢�>4�'=\ؓ#�'+�((���7&?B���'��%򁚎�Z�*��N�*�1H>	�=�^��ū9�A��oT�QX����	�<�ܴe���Ҍ_��X�MHw�DQ�"O@(;��Nb�l��C!�l4h)s�IS�������D^z�+8��rς)�!�Ą1KԐ2$�K����n��-%1ON�=�|�Ճ-eI8mpwH�S�����Y�<� LR��O	6��h�f�J�
C\R"O�]�FX�D9�4��JL�^T	��O��9�)�6pۤ���(�0lH$>D���	
�`{>d��a�$I9(8ѕ�'D��*�.C�F�� A�������b1lO�60����h��F͊z]X�E��qs!��bBJ-�1�.P�����$�9U�OP�q�)�$��2�򙡦A��B�2R
ˍ���&�O�aِ#� i|+�� I/N� P�'a�'КB /۪ ��аJ%�-k�'vL�w#�U�B�c0d�w����hO��;�I�V���"Z,�<�����C��	MPDtveL��H ����IXhc��F{��׋K�����!?
���  �"�?�ݴ�O?]r�d��&�@x�6�� o�D���Chy��'�tpP�}z�(�̼,j&��O0�'%�����`֐�-�#k	�*����t�]*g�a}BA(?Ig�ʃTzfa��'�N��T�b�'�^���O@j���F {�L9Jt��D5��)��hO����g��v�T�	���gk(d�s�|��)��;C�ܐ�E�G�p��X
W��	/�B≭��Ȥ��>k�.yc�L��I�#�'�PHx��ݜe���6�ġj΄�H<�y��ɓi/|tք��S�N9���+5X���DS�I3�䏧R��!۴�Z�R ��ȓY�u�w��'oNd0(ä� <�̇�V, ��)�T���p��29-��'�tG{��D&V���5+UD2�V���
��yBP�Bф�Ӌ�5���@�/�^�O\a�)�3}m��E��qc4o����Ue���'�{��.����c�Tb�K��y��]��m!�.�}r�X�sN�p>�H<�p�D�6��%�6�6:*ސ��#�O�<y��-yZ�	4&�Nɚ��a��hO�d5��:q�ǓoԐ)[4!�b�ȓzPj�x2�I3lvu���O뾰��&�r-�%(l�Ҝwť_�����?A��2If�sAjْ4���H@�a�<�-̈́l���p�������^�<-���ٰ�N�Ґ�aq�?h��B䉖.���0�(�8qw���sFU w�B��	jmZePg慣K�b�1�ՕA�F���4�O?un�� ������<:�e  T�W�
B�ɻ	�`���O�f$�Y�D?8y��I_؟\r�%��ZS�|�j�
R
2e��-D���S�_0N�4j���36H&a�Q�>A����9E�y�)ש_�"|;��g@�">Y��i��A���&RRb9���'P\��)���$����afH8w.Q�$���4���`��s�����Y�kL��S)n9K�"O��xa��Ot�|��ı_�T�@�>�S�'�џ@������N4D�x��Ua�"�ڈ��Iz}��_X����+W5`�B�0bK���y�Ä�{�0�A�*�h(ڱe� �y��^�y�R�`Gn�2*
N�Y�Ȉ��y��E>�M�%`N3��\P����y⢍-TRN��f�A#���F�ڂ�y�V#X�hH�S�6���Lʭ��xb��*f�8����L/@�[ģK�N�}�S���I�%8��T��+�~AS�N����Od�: /�S����"׉4�1;P�U}�'����J�O��H�CKU*ppF�W	��1�'��Z�ަ"Z��� N��L!�''���I3ӆY��ِA,��Ol��� ����*qw�� *��e��w�'B�ɔ�J`j���c��m+�ꍛ2iZC�I!I��Ģ^�B��H�m_�U�6�<i��T>��^/l��h�&����t�0<O�"<a2��U����"X/;c��" *R`�<i�S�9�C/J���"�C���O���?���Y(�hK�Ee����#�<�:d��A�a��|cԥ��,E��|�Gz��'.Ie��b�����M�	�'%N�Bf�	7�D����b���	�'8"��f�b��Х�[�ܐۓ��'&�xҮ�5A��E �N���(��?O6M�gJ����(�Q�  �"O����0)�t���*t4�2"O�
!-�V��R �;w:�1d�'t1O(I��@JP�a��Ø�\���Р"ODX÷��	L&ؑ�� �4�jQ��'X���fN���|Ak�uۈP@���?��6�R���{�a&ӫk�8��x��E	�)��t�n��C�/W�"��'��IS�)�'R�б&��	F�x	�l&N�� �O���d]O�a�'��\H� (�H�5�O��S�g?��O�0��%�C�;��6�.e���'��D�0��E[D��s�O��!�D6T9�U��;&�0���@���}���E�'�|-���;l�BA��EɕRQ��'��]Rr�Ô�R$QҏJ,|0�8���>E��'bL��2�s������\��'4*DC�fN-a,�d��F�i/T��O>��4��O`b�H*���AY�(Cf�G��u� 3D�0��*�k��is�L��1'��+�y��M'[��h Oº|ъ�O�y�R�M��-p�G�G�H�&$��y"����a�rJ�x]m+A��y2�L��l�H��:�Y��k��y��P�o�D*��((���N̒�ybO0ұ,��D� �W;�y�D�n��x��c�(�ď�<�y�5
_��z o_�J���h3 ���y��9h,�R���0.g��9bb�ybo��2�� ���!�h����Y�yb�:|U�	0V ��
=pX&��y2	��X����T�v���	I9�y"o��T�@���߬OoȤ9���yb�ϪF�1�1I�M
�y�ac��yR��A�1� @�,Kʎ�����y"�-H��q��.��\+ ���yR�q�!'D���Ywh@��y��F!rb�Hլ�5-FUY6��y��K��Ձ7���%*��@d�>�y���0_�ɩ��O=F�X�lV��y�T5:$����\�MG!k���
�yR���YE�㔨F�A��$hwc��y�����=�ʑ�En�1�y��ץqj�h����0��u��yr.3̊P�7��
������[��y�NT�J���	�	Q ���oG��y���WN��v�_&�mCB��y2��*��z���S�����]��y�ªc���j0L�x�C��yM�>,�,���חh����T�.�y�&��Q�*�	7l��e#�詣����y�ꀅ(��U�3�L���M�C���y2��H���+S瞦�@��(R�y
� � �`�J�RP��)�P���"OVl��cM%��!e��oے�q2"O"��G�i�F4E�N'����S"O�(��$��@���w醧~�X��"O"���g��djzdnԇI��S��'x2�'���' 2�'F��'"B�'t�P瞏|Y����b}ry���'r�'�"�',��'9��'��'p������8E�r�l�hl�js�'�r�'���'x��'l2�'}r�'�(y�gƘ=~����& 	.XcF����'nr�'�'*��'���'oR�'h��G�{�[@����m{$�'
��'!R�'�"�',��'O��'}jA��I!;�J0ۧ��(c���A��'���'<��'�r�'�R�'�B�'�����k��d*����.Q���'�B�'!��'���'R�'r�'��5�4KU�1�93��9y��!x��'�r�'+R�'���'��'���'�<,s���R�R=�d#_�[:���'��'���'6"�'�'Q��'���q�X�d�"�x��kz����'���'��'���'���'pR�'�A�q)D�@&읓0k��`p5�'���'���'t��'R�'���'��%�p�[-#�t�s�e�,[��1e�'��'C��'��'���'��'��9"w� 3#J�@�N
NU���'��'��'���'���n����O���W�͆���XCڗc�&�xUJ
Ky��'^�)�3?ᠼi|�`�¼:A��J7%�2r�ԋ����]���	J�i>���][�n����QF\{�@���5�M��w����ش��D�.\Ɯs+�<��S�N���LA�%Ӫ��!�*s�b���Ijy���B��,Rc�ҵ>�z�K�*�r��ݴ]j2D�<	�'��'[��w6.��qH��	��@<Z<P8�`��O6�z����& h�cڴ�yboO'mIܔk	�.�J�,�3�y"�M2�ZY9�n¢D�ў����Db!N;β�˂k�'J8H}i6z���'��'�6-X�sg1OPCb	��\ȘG��"�^E���O��O"��'�2�iB��>Q�k�
P��6�بn$���T��I~�l��M F�\ *�1��\|ݱ[�NZJ�B��33���� Q�t����,O���?E��'FM+���Bnޡ7qU�Թ�y��}�`��֑��ܴ�?�I>�'#r�9B��&^�(�)r��Pt�����?A�4�?qd�1�MC�O���Q��m��i6�T��t0���lBP`Ұa8��P2MΛ{P���b#^�a���/Ǽ�&��5@���1c,����n Rp�0b%�Cd,����Ý\�!�႙":�Y� �1bJ41F���� A�c$1O���I�Y�ı��J����ߛ%��L�˘r���`eY'5��������"��J4f�(��/��xǮ�a���2$Gu(f��PPp�"��g�`��1�^�T*d�E��)\�4A�&��(�����Dx ib�	{�="�CĹ-5��礒�g �/�~�S��J�L�!4c�>q�޽c޴�?����?�����I�]S���p��e�$q�☣��6M�<9�I�E�����'xZc�ȁì�be@�"U��T�j�!�4]V;�M���?��jT�x"�'T����N7
X`d�&lR!��if�p	#G�)�۟��I�;��̹s�X�*�#�	U����ش�?����?v�H}�'��'��T�_˴u�Å�6nV�Zf�	)"�O6������ϟ���ݟ�Z�!B�[�"!!��3Oұ��ʂ�r!�O�=��Y�	ş��	h�i�e�S�@Ipf12ңʸ�(<�7�>҃EO~�'��'bX>ESQ.��N�#'�2U5 �R$��Z��H<���?�H>�/O4��-T�E�p�S�\l�� "�ħ�1O��D�O.��<�'�?g��i@�8a�Iwb��t��u ��-l�'iB�|����h�Q�tx�e�8�a8�дP}<�*��>1���?)���I�&>y���;��i6a��?NAh��M����?9,OZʓ�I����B-h�����AV��4aD�Ț��V�'��Z�h�o��ħ�?q�'x���k¬c;6�*W��b��1贖xB^�l��4�S�t���]�@TO��R���R�M�+O̳w
��������� ��'�N�� �1d����E[� �I�4��Ă:��b?)r@JdQ�pk�p�҉�,gӤ�f�������8���?i�}bBJ��(قД�v�Am�L�L6MSz�"|��qp
�1��4;�@Gl�T\CB�i��'���S�l�.O����O@�ɧ��hB��/�K�7L͢�$��b�1O����O���ޗ. h�bB��dRIz��"I��l����B@��ē�?1�����C��JN����P������'�	"M��c����t�I�����G�z�����t�$��K�m
RY��`~y�'�r�'��'�b�':j�)��e�
�f��*S�	�B��*�-��O���O��d�O��䁈P�T��X�pmR�LM�]*��i����6m�O��d�O�O��D�O���@ �vO�v�Ю@F�B�IG�+�T(it�-��d�OR�D�On�D�O�i�Cc�O��D�Or-������l���\�^V�9�)�����I�	Ο��		Apa&�>�$��P/dU� ��t(E��+F̛&�'S��'�r��.��ϟ����?�zq�V<���-�&%���Ɯ�ē�?A�����u�BM�S�� x� Q_4|y�C�	[��@%�i!��:9ER��	�����ϟ|�SvyZcݺ� #o79vL��/� L��4�?���D|����eB�S�v\���35!n,��%�M�D��?����?�����)O���O(����3D�:��J�P/J\�#䦑AO�]�S�O��O�h�Yu� ���$�� ?W7�O����OLE#��<1��?9��~ք�Nc���Q�e9��.��'t�s��|��'W��'v�ȳ�>hdԬ@� ��O%�ݓ�Gc�|��	fFTʓ�?����?QH>��V_$��C:Xv��T1����'>��(��|"�'(R�'��[R�Y(�G�h�<��
U �@CV+�7��D�<�����d�O���O�et��<0XR���Ι���[*58����a���O���O�ʓ	����OZFus�-F��*Q��A"���4�?���?�H>����?��n���~��$�`L����!B�g����d�O��$�On˓OB��/�f�$P�Sa@ Y�#cӚ��T1X�RmlZ��'���	���Br��\`�՟�^y8�KN�p��oZƟD��ky�@�6}����	�?���b�0KP	h硛/�u���ګ�ē�?���-��������U9B�d���O22x*S�i9��.�|��I˟��I���gyZc�n�2 G@�"��P���{��H��4�?a�������4��4^s8X1��1u�戣H��M� ����?A��?���(O��D�O�����#��Y�I�6F��!{)�ŦeX��R��#1'/?E���'%L�,�>�J!GҒ ��� ��RO6��O���O�����<���?���~B�N�\����1ΥA��Д��'[��'�|��'q"�'L:d��#��O�8�'��;�2����m�v��4s����?����?�K>�1o���%�8�(�q%����Ҵ�']D,���'���s��'�'�����Q���4M�D�^Mb��I��tie�,���O����O���?!�\��i��ӬQϪ\au�![oNX�bF���?AL>���?I,O6���W�|��P�^ႀK@*CdV�ہ��X}"�'XB�'W��Пd�	*_����ɫ�$��4H�Ou��(�iO�q~�x�I<q��?�*O��䄙i��?O�؜ ��?�|����z�
���4�?�����$�O��������?*���j�0 �vI�F�¬1s&6m�O
�$�<�H�N�O0��5���9荡����Y��P���M�-Ov��O�8)�O���z����I��7m&H�����|�(V�i0�	**�ݴp�����`�����ިCR੧�g{�e��*X0BΛf�'����;��9���f��=*�Ə��u���xQP\���vӊ��Q@�O��d�O�$埶�S���O�kg5�4�U�t>���� g�`7�ҢiĘH1f��ӉC�`� �b��J5��,	j��ߴ�?����?�vߎ��?}�Oz�BB�]y��T���Zl1�؊�A�U�8P�ru�	�O<��5A�X�1���H���1&@ }@�7�O.e��I�<�"]?Y�?Y�b����t �,@�e��CVL�$F"�	�G����s #����'��"[}�x�f����@�W�y�v��W�<����@�?���?�����&���*a�4&|8�*�H��*�(�5�AQ~B�'oR�'$�I�	op��O+8#v���hҡ��n�g�fmp�O��$�Oh�D�<A��?B���?�@��7]	�E��œyw����}���� �	ny��'���1_>������hWgN�:0��s$���H9�۴��'��'�Z@�c�.��L�V4I�u�X�qw+_�l�̟h�Iky"�SQÜ�����k�^HݤA�&�ӣ3(�P�S�WڛY����t�爌�ЗO	���5��۲mC��Ca����5�׃ݿ�MS.O�Y"�E���:����d㟊��'~�I)G�~����g���ej��ش�?��Q(`M��K�O���S>7-X�F�����W>#D��Z�k�*#��6 !~�87�O��D�O����g�i>9�Dg�"P��٥A�M�p�Bb!P��M����?1��?a����+���Od�JQ
��*����R��"�ϦY��ß@��5��=�ٴ�?����?���?�鍵$_8y�J�M}Y� ԡ�M�N>��P>�?1���?A��?y��kI�,��G߷o4�*����Q���BR�i���_%D�7M�O|���O����b��O��k1���?(ĪD��.��ɭsG����t�	ş��IџX�OV#]d(�r�ЦZ��qj��	u٪6��O"���OP�$YU��V����?%򐡳��βY�.T� ��Q�؜)6�}�0�	ş���ߟ��Is��B�1��7-��@_:m����` �.�
`�p���$�O�$�O���<I�q`�`�'K[�}R"!�LDP�aנ#5ΰ*a^���I����	ɟ,�	+F��pش�?a��!<B�g[�_�6�!�N[4��=
��i���'�rY���	![��'���N�LxC�%{�j� F����']��'��@�#q6-�O����O��)Q�
��Q"��F�jm��NȈd��Eo����'C�	 ��4�'������4?Hf`��P�)�j�!��΀\GjAo�̟�	.]#&�4�?����?a���
�f����(������#�	0�1`\�����Q�,I��ß`�I�$��D�i�jT�$�� (52�;�ϖc����$-"6M�O����O������$�O����\��qF�Њ#�~���n�R$�nZ���IΟd���D����'��� � 9Nү��8�&�
%�Q��i��'����m�z6��O����OV��O�N�!(�n�a�d,�*�H�
߿��F�|bM �yʟ�d�On�$��%�� "�OP4&�0� P��r�J�m�ߟX˰*��M���?����?�S?��U�vp�3" &rʤX�/��MW���'괔0�'���'��'N�Z>�V�H/^|�c$��.Q"2���F���ڴ�?q���?���R]�Sly��'`x\�!�H��!"g�h{��v�O��yr�'s"�'���'��ӓ!Т��������B���`��c�r���a��M3���?	��?������O��Q:�����U�Y�X����na�D�ڦ��Işl�����	�`HC���M����?!b�xT�$��Ɯ�!�rQ�f@�V��'�"�'&�I䟌��oa>��	���Y��ɟ �t����]���(�$�Δ1b��	֟���ҟxg��%�M��?��z�R�P�P@)J/�Q!	�*K���'Z��ʟ$+7�>M�'��ܡ��M#�$Y�c�T�󱠍�:��1�����!��ꟀQ")���M#��?������?��\%��Hi`�),�
�T��B4�	۟�9�A���Ry�O��'Ev=KI�~�T��� �a�0�o��N>}�ڴ�?y��?�������?���A�L��Di֍c�b���i�6���j��iD�@a�'��V��q����TLF
���t� R�n�I��M���?I�6�2I�i��'��'�Zw��9s(�PQ�S�x�"ݴ�?���U^]�v���<�Om���'���L�:���S!�Џ~��=`SG\�V\6��Ol8�6������	�����՟����7t���F�hɤ"�JX4~� �E:��ϓ���OV���O\���O�x��$��z���� �;9Ω�E�UE��lß�����8�I:����<y�=��#�<u���:R*�	����<I/O�D�OB��O��dA�q��9oZ�}Ψ*�.P�OĨ�[4��&�z�R�4�?����?a��?-O8��=$f�T)I��q��؀SNq`a_3�n-n������������I�2u]�|lZ����I<NOtc�!��$M٣i��F&��Aݴ�?y��?�/OL�$N�3����~�$\:,�� ЕoS�c\@"4@Ч�MK��?A���?��ջ [���'`��'���KY�Zh񅂇�%Ä9�e�uӮ6��O�˓�?�!���|�N>��ѫ�S�TL���.,�����hӞ�iоXAr�i�r�'Mb�O���Ӻ3 �% ��]ʵ�)}�� i��KϦe����T84�q�h驟��!u���bw�L�9�j� �*WV6�U#⠕mZ�� �	ן���?�I��X�	�="qC�&�2xq��Ε6P��`�4xx|�Y�����|ZN~��I~�A#��B4�D�ܭ,):d�ib�'���BJ6��O��$�Ot���O��ԪZ;b��ҁ�4l.����Er'��|R���yʟ:��O���֎
�*��s�E�e��E�,БlZǟ����T�M���?����?)�U?���_t�����p�N� �C�'kN��'��lb�'H��'���'�T�8�@yŔs,e�
�U�N�K��KI<��?�O>���?��3&��}i+���F%01�Y������d�O��O��iT\�w8������QP�-��Cסk|���W���Iş'���	ş|���PݟX�g�K�p�F�p��?|��{TC����D�O����O�ʓm3�i����D-\�F1�tR!��{� +�ʓ�l}�6�Of�O��$�O���H�OR�'�6��N^ľA��G��*ش�?����D./Rq'>E���?E�F�x �(�L�6za��W��ē�?����n������S�T��{����nB��V��s��#�M�)O�Q
Aަ���|�����'ˢ1ҳeG�5�D1�׬�.�4�bܴ�?!�6`����S�'B�X��Dī}���p$S��]o�5�0b�4�?����?A�':��'���Z���UeKr���#clF	(�6��?[����1��˟�K��Z2;_ �;�	�^�؃�C��M���?��	"TX��x��'s��O�	e"V)mz�`Gj/+��t��i��'��d�
;�I�OJ���O@��rh�������Ԋ�}Y�@�̦��I���}AI<Q��?yJ>��ˢERs͔� ��`Q�ӟ>PrT�'��q��'���������l�'U�l��g�:���PM5p��@쀏~��Oh��O.�Oj�$�O0��$I'h@P�&k�3�$API +�D�<Q���?	����Ѧv��̧_��#/[�,	Ad�I�vŮ��'[r�'_�'Zb�'�ae�'�z��c��Z��0�d�D )�����>���?�����K�t�|�$>��b�<������/"6u9҈R��M������?���muB����. K�6M��}�}���Ԟ3L�6m�O��d�<i���QT�O?���5�O�+1�<���,A@QXq��
��'W����r�|��<t�t�N�}V�sE�M��4
��i��ɛP�0�	�4_��ʟl��"���V�3R�ą��MN�0��c�'Z��I������,��'x)��#�,��v�Ƚ $b@
h�4�nZ
ℽ�����I�T�S����@�DG�t�H�1%F�{3��� �N�~ Dx����'�H���M�;��)�b16��̻��`Ӣ�d�OP�����'���ßP�	6�Y��B�Xa Rǀ�*4�b��d4�$�OP���O�d����s�2���J�GL�2�\���I����ON�D\y�D�'W�'���{AT�K���`A�b1��*�9��=3:�InL�7�@�$8�j�� ")#p��-_�b `s�֦
U�I�e"O���@؁NG�<y�G	5^�H��	"@����3Tn���\ร��V�GA�I���&@^>@%aK�1��UM�RP=��d3^�T�Q�S�kt���<t6��B�gF�.I��@�Y| @a5i��w �\�'�?T�l�0�di�����
T(2�F�qȤ���A�f��8Cf�>[,����:�0u����<.�L���-D����>x��L�U�'���'��dT��M�vLCpKIѦdoZ}��E�C�J=B?�R����e��[��]���	1�tdB��9��aӀ��a�ɛ-G BZ��:R!�:5�>��D	U����	)x���$������E�%1k��Ǳ!E���n ��yB�'�}Bt��年!�0C�k2@����#��|⅚x�ǎ"X���(!�Ϗ�A@မ
�y�G��1�X7��Ob�$�|r�HN�?���?��Ʉ�$z�`3�'�2D�X �L�Ȓ8Q�>bA��Y�2�*��b>��yT�HcD,�'o� � �܏6�`���E/q�,Xzs"A�9Kai3
[�i#V�RG,�
����p>�Β�~u�+"@"9Y &���&�,��W�Of�6?%?&��5)��}l�=hӏ��V��s:D�,P�bE�WZ,��NA�Ls�o6Q���'\0��1������]Ȅ��	ʣ�?�������d	�?����?1�Y���O@���3���j���B1�J}1�۴
4�)�'h��Q��?�=IB���&� �
��Yv�QA ����7�޻b�H��3(÷i��p��hO�00q�A6���&D0MJI��O��9d�'��ey�i�]�P�Q�98�c@���y� �0Hr!�ed�D5�L�`�<Q�."=�O_�	&WE�=@۴{�RT�歆�r�0ey�FH�j��9���?���?����?Y������E"\n$���*x�}�bI��8d�=}֌8��h�7�V����"@�r�p��0IS�H�0&ݑk��|��I�+x)FY� �'=i�Fʘ�6G6B/�5?qd��g�!?	��˟ �	7g9�Vy�e¯�(�d�G{��ɴ3���`cT��m�2KZ�C*BC�I�r	KYRZ���m���j��7OzX�'��	�/
����Oj�$�|چ���'6(u��5��Ѥ��[�R����?�����v�'PhUa�/��$�)��襀�����[6Zw�ԛv�I)^S�T��bA	�ȝ�,�/Z� 
%ādx�P	�=�0e�R�]/r]��qB�#8M����П���Al��LI�H?��P���<	��?[F��eq���k��c�X�'�ў擔�ē2*P
!��Վu;0�];U��t�"��ٹA�iR�'%哯jI�-������<�,i�� U,��yb��%�8��n�.&/����X�	a�S����'�JhW��s|��Te���&N�B$��p�GZM0R���8O?�D	-l^p����Ŀ?s��p�`�"Ȕ���E�Oj�oڔ���O�>�9�ȡ� �̔s�|��OP
�D�O������H%�e��AN�݀Xh ���I��HOH���O�UhƏ�<<j�*�$��8�dF��O"���rT����O����O��������?���T��0��C\&76��i$�\ .٘�!��A�^X��C`vp��'�HO�l04%C8<\0`�醾A�e����b<�c0�v�hf�ݚ)8�I6ғ^WP����	!9�`SR,@+zanY����ƛ&�'���'sb�'��w.�,cu@ݾP��m[�,�Ql.��';\��`ʎ	%2�3�&�QVdհA,:ғ7�v�'��1:�xٴ��sv�+Xj��F�J��,�8���?����?9a`ێ�?�����t���*r��Y�ƃ����z����=�����C��h 2ˑ4\:h��n\C���Fy�lA�z�`)qL�����5 �z�Τ0��J��r����d2��4)A�c�h EyB���?��iВ4��nS�l��)��J� ��{�ci����<��������Ҙ � �:���)@lz!��B��Z^axB�	2o�lx���df��{@3���8h=����\y�$�M���ޟ`��]�T#�:���t�1<z��0Lݻq�Ջ�'���'�rmt(U5��rg�9uh-1˰~J'�!gh�!*����^l�z�Yw�'mx�zD�K:TH�K4�-2��r$U?AB��Q7�u��6 �>��aG7ʓwt��I�M���?I-�X��A�ا<߆	Q3	ϸ�>Ly���O����O��D�O�I:�/��\�����pZqlA��\\��	5��-~����ݞct`)j��M!~"���'��7��O��$�<�V�ǣ�?��?Q��LC�`9 A��7��mCBf�,���W��
�����`G�M�cZV�&�2��E+F��h���`HN� 6.ܢ:�K�	��h���ܟh�t�s�ʍ� v�`ᥘ6]������'|�6ML�i��h��N���W��1��	E��H�k�����'�Oأ=�C$ߴ�f��jƩ�d�h]j�'������%��M<g�8�G�S * ��BK��B�I~���p���Tw��S.�
*��B�	��.��a�m~�x� �^�*�B�)� �3̾s1���P��0Ԋ@"O�p��Ǖ`�D�C��ǔx)�"ON���l��	��YȠN�y�Nсa"O^���3���Y�ҹd٘h�r"O�	�n�)jj��a�9)4�1�"Oxi�'$NV����h�_�U��"O���-U�p���'b�\څ"O���"�Jh��8�U�V�n���"O�(���1i�]��"V/B��8D"O�	�0i�j7 3�O��a�@�h�"O�Iyd�%J��K���tX��"O�űR��体F�~y䘢�"O1�gB&cE�w	��E[>�J�"ORY2GhR�B��*0b�x"Onm�� ���Ύ���90"O��:��\B. 3�O�U|�w"O�t����X{d"eG�b�� 6"OxiC��D�0�d30쌳h����"O��p�H.�u��J�
Ucl��"O�i4�/:���0�	��sp�EK"O�� �h �VP�أ0^RXRG"O�q�(��T` �`,��Tpr�"OU��I�^�1�^�4�Ȓ�\6�y�m7~ּ�!ǃ8=�&�bW��!�y�gMx�	!�g�%:F��Lӓ�y� 'K!^P1�ş1srX�v���q�rYɊ�OY��g3O��`�X.E�PKS��
@�R�+�"O�zgM��*��թ�1P��h�O(�	'�4��+zqO|��;Hڐ�2���2P��Q2��Ku����$<2�9��� �|I�p�ԩ>���0/����4�'�ɑQ>7m�E�p9@��#[08�"@=ay�*�%TǶa&�� ���!�P K�Ƒ���cw�>т
I
 ����Ę5fw���nЛ��	a嫘�[(�'�f���GQ��|�������WsR��	;���K3
� H!��%Ut��d�*\�\	a��6�0➰K��O�,���D��3ץ�=N���ۦH�#�6��f�aH<)a��5Ft�9�c�2$�Є�4��X�ɹ��`2��sӆ|a�H�a%�$)��F�%l@�p��'BJqKV"�m��SW,��2 $<�*,�Ê͝U��A` ��Si9|O����	�S�I�e��?]fx��^�`p %�=~t����Z�3}�$��n�&2D�W攱�HN1K`���'>*`1��� U���8��g9J�s�4w��֡@^�I%l�6X�"��xs����y'!��`y,D ���4�RX�"ذ?A CRA��GkiG@�W��R��4zb�O�h{�:O��`Q��3K��족�O�T�I>%jT�+Y��ZFĝ\x���V�z�'#�\˦$�bnl���ޕ:TЌٴp�X�pG�]�6��⏸P	3�U@����'bJ�Ovl��ϗ���ɼjS���`�Y4M
Y�G ޴�B�cL�h0T��Bp�T:�jO�i�JE&�tzj�O�84��T#0�JTg�8<4�2/1�d�4K�<5�Ǔhl�բ�Y�.q����}�]�B�K.AZA�q�|��J�yr�<N,�Z���<�rBN�^����OVM���#���h���������P%���E�l��-�f!�<��@B?���G�<	��U���(�
��]"b�Q�)W\ԥq)�!c��"?1�*�>��&���QY�o�*r��|�c�V%>��p��B���x�7��7Q�H����֍
�pp�����RA��<4�PX��"�ޥ����L���'}�&�v��E"���H�(-�K>a����G���I,4��� X��1
�&�84�(�t�S�8;0�a� �����	�,#<A���:���� �2I{��X1V�P�k�_*f$��'R�I�bx��� `*��Dk��Q�;�rH;6����Qt	M�~��g'��'+�������!L�x0��Z�-.>Ma�n�l��#�M��Շ)��b�x�1�ĥ-����K�6������r�������Dx���������C� �X#��G�Pq0UAG -��؊֍E2�x�]����#K5M��]�P�Pp2QY>u��-cԨAT"�!&�R<��\L�b�OR= ��L6-b� 4F�:�2�gy��d+.}vAD�{ļ���,N.R�)2�Õ%T�	&�r0�vF�?]��/�1O�s�kª9H�Hs#�B��yg.9&���Ԫt���)p��qy*�����yR�-����FiB'C�p�
��,� d�VAK,&u0��� �џ�=�  hs�!i� G�Ia�ay�mأX�L�#=O��?��wC�t��!F03x��a�/D��0�1���XAl�J�-�m?�hǌ�s�n�`�%�F��#��Z�Q��3��*Fډ'#2��c�s>%���'D~Y	I~�J͢8- �����09���I~r)D�Y�
}cvN[S�V�[���?�3��ݞy0�[Q��2��=��+j��6�&>������G��PbA�Û���ܞ��i�0
I�ܩ1o*[]�`�r�1K#@����������N�9�yK��:��B3!0ntk�,�#5�ݘ��Ɉs+,5�V�K=P��4�2��t�V
~V�@��2z�l��?��D�<Ya���������&^�k��`l.t2ț��O�y�æ��>Ӏ���i�`��!��iZ�w�x��
Q��qFI�Sb�D{�ia��]�����C�' ���SV�?��ώ�|q�a�M)1���!�B���Rდ-+�J��p%�T�ހ��o����|��)@6y:2#	�kM��c�	�����Mk��<�Nġr����J��Js�I�"�dx��G��Bnx��	���u)F@�9�����Px���y2�̬!1J��샿!�B��/���D�NK>��[0`�ў���Cp��!HG ��y�lF�9~��� ��pR���n�':H�`tHY*&�"�P�iU�P��d8��	)^(I�B[�:�h��L�����&Yj!��;��1��J�W����S`�O~���'otehÄZ%�\h�w?��;&�S+/�v��rhJ`��'�<��cW�m�su�&k���9�y�$o���y���V��� ʗ)]�X��䇌�Ot^�*�Ol�0��99��`Q�ў~�@�0�{��_�$FV��c�� �VR� N\��dIfl����'��D	�l��yn�I(Op擛��mbeC��VK6<B�K��\N�k����h�l�8Q�������ȓd!F����тB�.� t�f�$z!mߒ%8�G�<�-�(��b��7��8������8V�(؉DO4�qx=��6]��Uâ%{��2�er����˱^��x��'xr,`��|�� -��$�"&�b��W/!.�R�!��p����A�-�ʁq�D6���O8 �d�ۦ�8�He�d'��0L1OXE��/��4Ħ�� i�QX�������l+�nK9	��	%s��o�FI�0�lI`�=B�;3|^ibi� ����iC`�^�1��v�d�N�qG�4%6,�'�󉚁;`���V
ml��EOt���{�`���.�&��OX�@�w��B-��x���ˠe�?d���r�'��\�Uj�R��VX�P�O��OTF�K�c؞EW|���?g�Y3��ɨ2�zٷ��@bq���+F��!P�y�ץ��J=!Z��D�mur�;u��Ѐr��M���|�RK�Ae\%��/����7�+�u�+EM�XAK�Hׁ�y�F�/>R%� ��t�"�ϼ��I��y�E՝}_��
KȮErA�Rg�,�]B�̍�d��i����4w>���c��д����H�*{�x@c	 jҰ`CCg�A��Ũ���<��	�9p��s���<j��� *�f�],;�H�P�/l�l|����i�6�Oպ����֗�Q���gC4l���+�E�,[�@0Y��W�$)WOK�t��	�e�E�L�O4�I�L�g?�
9�Q@q��)P��С�S|�'y@ A�'WJ��;$X��x��'�bmz���7�>ܙY�qÇi�٦m{���W�����@0J� �p�O~\��� `@��G�-o���I��T�vΐ�C���=O����Aՠ*g�;0�� Z����O�U8aDԑe�� �@�M�/�n����_6|��u�v�<+͉��>��`�V!������O<`�t�=9ƯY�GȦQ�+E�w�R-����#|�$x�d
e?��n�F�<�Q ����O?��':����Q��cM�@Z�OM�x�4=� I._�L�9Ҭ�EyQ���sEcޭ1BG�)�p��'T(8a���h�4��C	�8�)O�N9�矘��G�#��9�e��^	ع"�-�S���*t@6����#�����m���Ť5���vE	;��X���z�p��.��LD��Q�x�Mu.�"g��3�y��3H18��(^qX�(Ơ�y���S�l ���Ub����?�'to��;�o�'<�@ɀ�x��A��X��=B����,�'1��y�l%��Ԡ'�"_����=�!�S!��(G�ΕU���e�{��]2��\[� �m�-�53��+M|ڞO����S��ZX��GV�rI~U�'i�� ,>4Y��\�d�G~�Rݼ�!��F����,�}�BES�fّQ]҈�b�9��mZ�(��-9^w�D��I
Q;����э0cȭ"Տ
'h:8�
�n�Gf�>�8@a�ɱ�h:�`�$8�,���(��6D��l��s�VL�	�H"�o�V�Z�d���(U���;U�*��S��;ET��AW�3C�'
�����Z)&��!�G�?��c?�I�h��PI�+��z��
�e�
�'�7�jd��(+�e�,UP�>��'|��VeQ(K��¦N�M���ǈ,������a� m�p����'f��g}Zw�hT��&V�@Њ�+��s���a�V�zJpa`�X=��i�r��#4(��� ����*qoNw�=@��R)�Mc�i�����'�:�3tHǏ"���,�ݘ!���'�~���H='F����4o�8�ܪ6%"=����e�d-��! f���hW*�#JN��S�AƲ(�"ҧ�' L�T�,{Э�#%!d�S�,\=�I
~Bɚ%��8z���m�p�'d�`�h��VZ�S�N�5)�8�	�mC��j��>�2[�%)Yw�بK��4'qOh5 �HK�8�x1[� U�*��V�F#R��'��P�e�)x`U@�?-`���lg��{���7���1���wH��t�[�7=��{`�`8��]�uΈX�	�4[���Ñ�K��Yㄈ?��i�'�]�w���� �i��M7��Z�ጅ=��� ��'�j)�ǪN�,�#� &Z4 [�(x�X���*}&�|���o.����r����x"�5!�U�OU�8��5��F�%v�ɠ�ȺD�l������E�I����3��)�`��O�[� S�I�@�I o�<̹w�۴(Pv( wB�7:4ʓ.S�Aۡ�)M�����O��\�g̓_������,1F�
G.𡑁�t�t�[D����%~42q̓��!��
$2�r��SFDa�hY�U:rڬA �'��~�D���w~�Y��/��	�!&r>*���'1r=rӏ���8��-WCNn�a��'��1X�ほ>����PHC�`/
0J��p�	ϓ �
1H��V��� Z�K�^�S�], �HT`�֙M=^9�H>a�ƹ�^8����
qE�� &�Teܓ'O|0��̅9y����R��Y&�����"~�Xx���!#�]���!�ɗ1�" �h��U����q ���}� �A	�(X"�ڰ=12V	X2���cJ)7I"((��?�!�}V��p�,2<O`��a�[�mg��J�AդV%�a�Y���O���� |�Ĭ*Q�v�ja�`��X��[Q��3GlB����ě?��pJ�+"\ZDb�̙A$>]kuJT���'���z%"̲�\��*;X�� ��J���d�~Z�8�R�	�Z ���8��'���B���1�v�0�G�2G�*��}r�Lg��:�JƱ2�nEK�Ͱ:?��s���3+d)7�F���-�w�<���5�7/RK����FF����N=s"ĳP$A!��)�'h*��*0+�=2���څ��+6H\h�"

�F��{�̕&h"��j&K����е�N$j�
d01�{?�P��u�"P�S(����4����čo�xa�D�*a1�]����- �i�g$�9�h����$��+qڝ�(mt��%s�ǋu�6<�gO4j�F�'��S��l�z.�D��e��e�"��1A&��
>�s��<��NY�?���s�@&PSʵ� 7O�����P�We 1�L�J��=���'a����Q�ڔ�OB��t��9g�zT
]�8�j����8�ЫB�X0��HGAEA���DαS5�i�4j=N��6iX�T��9Q��#bD�m���
�I�s�4��>g�`L�0�E��yG�¬.N�܋7 H`{
��פT��M�U�S؞4+Q�!K;�a/Lޑ&�7a�Bx���#�A/PαS"�!By� ��-ga`���9�HO�!�dl��=��<J�ˊ1i�3�I�쓲��pX3"e�>����x�j�
E�A2�H��<�Ё���
5����1~dI��D�I���r�&ߺH�����JLx�̇�wy֤Bf%�8J�����i-Cj��D�w��A�<1h!���t�F�Rf�)^� X� �y��H�{C�����9��yGL�/'�VqqTg�8�tC䉃r���s��&�DM�Bܝ6�B9(�Xǰ?�d�Ƿ�l��T��n�04la�<iq�б)
�ɫ�d�a�%⦣V�<!a)1qv�3#�����9�Mj�<ѣj�箥{g�-~:����K�<a��[�|Ȥ��R� e!�lJ�n�}�<�0�ƴf�$�*�F�B���bFN�<w�ҭQVP�Y�V�,d&�����M�<����%hW8+v�M2'FfA0�OL�<�7	T�%ܜZ#��b�œ�F�P�<9U/�;sr���!������Ǟw�<y��D��kd��"��L�4�y�<%�J'C]�:$���m��9�Λx�<a0Z	Z���{ ��F��XT�HP�<	� NLS�h����N�*`��lWu�<��FR�/�����C<�!�a �m�<!���:J��]�Ql� $@HD�<a���< gi(�[�Xd��$|�<�B",p6�1� @_u��-�y�<Y��L��q#��U@X����O�s�<��	ܢ@�N|q�*_@���T�<q��o��X���̉�]`�[
�'EI��'&1ȼ:�e@+,|4c	�'�!�$:�k2��ZB<<��'�P�Ya�[!}�.0�����^6*ѣ�'���b��@taC� �9c�.���'/|	桔�PJ���3N��9�ʓ�d����l�A1QoK+-z���v��� 0�Խ8Z���{%�4��G�2)�uL��h���(�m�����S�? l��1Q�p���=pT,��"O�e��$�1�(0�Ε!
�FU#�"O��q7�H>fuT��Pc�&s�Զv"OT�3�o�nS�c"�hކ1�"O��z�	�u�r���"��L4�h(�"O��95!L�;3D̥u��`B"O�E�IF�qj}�Ё�� n�(*�"O�bbhFkґq+��}d��`F"Of�R��^x�9���Z'1I�"Oz(e
X�E1���=]���"O��	� d���P����ʰ��"O�Exq`��/-<z� ��(��H�"OT��(�"����8�Lic�"O���QF���\h�7/�,�x�"O��
�O���-�t�X��n4 �"O�8)F�Ì �>yJ�m�t�@c"Oh��tɞ�~��ХSLn�PA"O�1�I��t{�	�ӣR�Wcl�z�"Oƍ�i�4P�<�P���uF�4Y�"O�����»w�8G�`GDke"O8l"%ÂW���IfF[�w9h��"Ott�"�����S#�@�$��"O�<��-�/��b֪b�&)�4o/D����Z�_�}��+�-_Nhx�.9D��:��6a�|U�$�VM��B�	#�h�j���|�el�I��C�	�wN�!��O�x(�zFl*L�C�	f*^�Iq��'bH3`��Zl�C�	�ub�1�ŀ8H�]Y�Y�sfB�I�l�ڥ;�èP��5��V�A�DB�I�(,m���0e�XC�*�xB�I=B��B�D�R~��X�ԣ�B�I$ �",Hr��6 j���V�P@m�C䉳m�&�Y@h�pP�p��[2N��C��s�е跋�1J|1#���Z�C�	`�T 8���H�"��iC䉒4�ū��!�f�9g�U�gf�B�	8�K̖J�
ɡc��B�	/j>����)߳O�R��5^!"C䉯k�lA:�BI%�ơ �n ��B�	9>���C/T�a�bɩ��ܨ�B��  c��15O�$zh&m�$a�<:�C�	�RST�{�'4TaY��$��C䉔Bjb��-@u�&x�ƞ|��C�	_#s�ʛn���o��i��B�I�FoH�1� �O'��蘁b�C�ɟH�<yB#_3���:O� ߠC䉼��ǂ��ȣƮ��2B�	�tA�@������њ��L�z�B�ɮs�Er�G?DV�ݳ-L(F�JC�I�Fɋ���?D�J!��H=8T�B�	�8D�����\	Jn5��84)�B�ɅF�f|���=�>�� &.4�B䉜
J��zG&��n�*��+����C��J�������i�E �㔟#��C�	 ".��I��]+"�t`Adͫs�^B�5^�*�b���#��=�1�
�V��B�I5feT��Q��V#<�2�GEe�B�I�]��a	D�֤i��t��
ǵݨB�I�qX�qF-4�B���B!J�>Y��	/3��a��
G7JT�W��8w�!�$�%{6]cc��)7��GB3q�!�d��.�Hr�����q �� >0�!�ƀ%<��H^�PA��S�Py
� TҐ�ƔM�\J�푎L�t�"O��cc$�B߈��R
�&��U�v"O�	�����^bA�efG��� ��"O�J^x0���j���"O��)�2@�tv 2d�Q��2O�=E�k�)`z 3�g�,UG�i�sO��Px°iiVQ���7Ndr�"F�è%�(5P�'��)
�GN�t*�@���@�	���Z
�'�"\"Dh
�uD0 K	�?p^+
�'�r��;�r�qL�c���	�' �qe_n��'~h��+	�'��Kw��j��0���D)}S�@�'ڼ5�0�ʄ�G耗n���'w̥���V�X&�ɬp
8��'���⠯W�����l�1��y��)�^KHx�@5g��� �Z��B��N�᧎�5k"��k�哟&hC䉁8�*7�QnPl����<�C�ɵX��KAH��u����ځM��B�9e�6'W��� i֌ͻJh�`�ȓcS�5s2�D�Hj1[�4l�:d�ȓ1I����Ed΅�pʄ�=�vQ��c�ay��P>��j��O�([f܄���qjN�IM�2���2&J���#q�i�tċ4]�(}�S�X?Jnp���jT�PC镔��Mb¢�;l����ȓo�0�Т�<
��Ӡ"ۍ@6�)�ȓ>��[��X
��U�1�t1�ȓY�Zl���]װ܊�)��̈́�4�^�9S�܏��b'H^I��$���b-�3!�\����>���uV
��"ޕl�ܨ*�� � 8��<�ߓ�K�)cdt�q�R$U��XPl9D���6$ÅN_\�aEG+d���+D���랾t(�Ț��O6K�B�*�))D�$����I�Q*M�?\<A�Ǆ:D��H^�Y��1HS��/�Q[S�9D��{�Ɓ�p�rQ�H>\ؠ��:D����ؔ<&H���>nD�L��9D��0�hїyD�!.���0���6D��N֤p��d��?E����p5D��4J��l��}zV���O�X����hO?�$G�@�Q`U�sU� b!�P�!�dB�Wz S#��=:Rp��o��!��G�tL�a�R曉;������Q\!��ĠS0<���ۢK&йħ���!��L�d��dPD�J��@�GX��!�D�+i�k0+��K��̠����!��2�x���Jo�p��ڸ
�!�$Y?e$�����*o�=Zk�\�!�d�����9Z�!"O�h��O��dU�a����5��Y�P��ڡ�!�$Ãd�.0�`�WxV��TfЩ�!��� [d�4j�"V,nH9v��$Vw!��Ϡ>�9@怵#2,$J-p!�D6p�^a@�F袤�RgjG!򤌤6F��3�!O\���U ߅.!�`������hXy��o\&m�!�
�xȁ�Y��țbiРj>��,�S�O��]�Q-	�e�rT`�ɖ#v$]c	�'xvu"�.ia����Hr�X�@6�yBǇ+r�D����@P�и��3�yR�[G������N!M���U'H>�y$�x�*���*D�0���)I��y
� $y�w�=���Y��WA�ڵ�D"O�	�E��_��g�?R�^���"O2)p`(8VB5� G+s�z�ٔ"OJ����R}H�J�t�q"O @�E���Ƀ"�@�}��)��"OZ����R 	<} 6�D�(�8ɺ"OTl+S��B�,��:tV$sdO2�zd&�4uC�nN,��B�͍Y�<)�N� ofЌ[��S�r@�19��Qh<��*ҲOk�`�B;,p��B�Q�yr	��W��	��=*F�JP���y2�֊A.:h	�(ɋP�d�`W���y�L�$X�M��1E8�H�1�*�yr*X���4	Q��jWR�1�H��yrʄ9>����D��]E��
�����y"�!^�,�i��lu*��uś�y�=FN�0�n��h�d�c���y�� s�� ���<`ֶd��Á��yReFM��S�;`�2� �	"�y�$�<v���q��
S_,X`"Z��yD]�K��q���Ұb�q���@��y�,�߸�i0naV��p�G�+�y�e�1:��y ���X�����E;�yB�,
�D��&��[�"�I��ͷ�y��50D�x��D�<$5D-��y��w  a�%��e�r!��!P;�y��KG� �c�i�PfIs�B�y��ȑ7�<XЕ�	~��|�rhB)�y��Y�J��OE�|why��	�y�eA!fS�AP�lt�vh�a��y�Ȋ�^Qjwa��<'p9����>�y�#=���rd�,28"Y��è�yB�J0wd���+�/�B�z�˸�y��Ҡg�Z�Z0/T(�Թ��(�y�꘨H�4a��	��Rd�A�>3�U��8*�@��B�4��Tˀ #ب�ȓ)�~��.��T����.7ԇ�Q�x8�#+�- O��S�X9C�]�ȓt-�����ϨX��k`��[��|�ȓh�^x��됙:�ʍ����BG|�<)����0��D��]y���|�<���.���p�ή^nh(V��\�<1�Ԟ��\��.�&�ڵ4�X�<12Gۯz��H���Ynb���'�V�<�4B4.A��JC���y��'Y�<�DǄsTU��mCf2�Ҷ@\~�<9��O,t��E�Rx���WM!�$\�)H^IqH��uv]��%��p�!�C`��� �̭C��5ƅ�_?!�$��k�Ш�7#Jp�!Ô�EG!�%,Y��`�H'\E
��
�v�!�$��-.�)�D�0s��aq�EY<r!��Xr��EskL�B!p"�N:�!�d֥Cb�x����Eq�TSՈۻX�!�dI" �|o��`p��C�&�	
�!�I�x>X��xo�R�eξ)�!�D�8�v�5KZ'Hmb����>�!�DŬm~|�bW�Դ[I��3p��.r�!��-I����Iċ^+��ѕ�N�y�!�d{�lq�̟�c)B�# L,P,!���.<Jf�dd	����	!�� gȱc�'^�E(��uB�;�!�d%�3w��8,�)��«W�!�d��Y
�8Y9Ό`dy��-D�� �0#�#�9>���q�ܺ XМQ�"O8dpr��J7�=�5��
^O6QR�"O2-`�B�cN8�:��>a*X#G"O>�;��[\�l���NFq"�"O����!ՙ	_�)�#�ˉv���h�"O��rf��$$�����G#i�.��"OfH9C��@�(�cT��I��\kr"OF:�i�Hy~�TjH/Y�
\Ȗ"O��S���9hǐ#0J܍2�2�v"O Ah#�
GNqQ�X��Hۓ"O&���dSg��.B|�U*'"O����-��$�@����"OJ��"o�)�
���-&��|S�"OL�޳X�f1cu� ��d7"O�A�ce�	X�����	@ �x"O�8p)
�F(�a�BL4�p��"O<)��Oq�:p���,\�dy�"O��T�D�3ӌ�i�k�>Qb
�˱"O敚0'�/�"���]|�E"Oz$�p�X��
�o:A���"O���p��G����-�#6i8�"O��cǓ3ctq����}�L�E"O8����0Lx��hL)�H��"O����K3U! `��)����"O ]���W	m��H�e�N
��Z�"OBE�A����+�[�^lӰ"O
ȸ�S( ������7b�
�"O��3��ɰB\6��<U�����e2D�أ�	�&J�J	{F�ױb��i�0D�0uг<��`+%�����$-D�����$ǪE��͕81R\L���&D���$>XC���T�x�DX��/$D��&eԹZ�(�P#:��uЧ�"D��7̒� f<m��P�\�a��J%D��r M�,4,�G�<~�B1�&l!D��[uG�_L�yS��6t���>D��QC����$�?<AF��FF:D��K�"��*���gC���*�)9D��8t럮D��D���Y�
%��BSl*D�H���ܘ$4��iW�u1�BG�B�I5#N�@�B@�iS*ͫ���H�LC�ɭ��1�"�$5\��ٿ
�lB�	/.���&jQ.
@T5�+�.�&C�� .h�-#7fق5u��V�.��B�I�DѨP��@��,�2NR-45�B�	���t���H�B����҇+>D���6�Ɯ=�n�"4ݨ"/<ŉs� D��h���GS
ܪ ��*JjQ�6H<D�L�a��v��2� \*��$��;D�2P��"p��Q�� �M�`8D��cu�ܳGy����,�8mj�hcա*D��X��<�e�P$B�3Eo(D�|	���b�sW��1B���$D���.�+�$�c匆s���d�.D����Z%t�b�j�a��_�hXw�1D�T�WF!eS`�s���	x/�t�¨1D��ҳ +D銽���[�Y��swi-D�����8��]���V��HCV�(D� �R�ͱ�(E� ǂk)��AW�%D�����<X��z��ȩ?ܾ)��1D����gL8^C���7+����`��I-D��B��90l�9�1hF�H�ӱ%-D���Wk.>�)�Ԅ�N�Au,D��h'���<��k�<a����W,+D�� ������Mfz܂W�� \�$"O֝k�����b�T/)=�`��"O����B2��$酎L[��aI"O�੤K���
���KRr@|S@"O�h��M
u�p\�e�ݓ��y�"Ox��TM�rz.�5�0ݺEau"O�����!4������7�\���"O�X�phN��h�#āf����s"O"��cڝ���g��9w�r�"O���7J�-ᮌ�햓_�,8f"O&љE�E0&YW-%��T�"O��:$i^b��u�G5_�Dk�"O�4a�ɚ;.�������\a"Op�ʅI=/3j����w��34"O^��dOW�<�L�z��į;�^�Җ"OX<�$�;e�ҩX�BZ�v,��"Olx�#I�����D9�XIɆ"O�u�[@�������"O�a�:`��s��Z�G�Ti��"Ox��7-��$I���7҅=�6E�"OT=Kb�@��ةR��W����"O�A�%3�|	����A�~ �W"O�m�BK�?g,�$�1m��g�FMd"O�XӔ�Vs��Mx���<~hpT"OT@fL�L���9�*ƀ��� G"O���4�TNҬ(
#
«z�� �S"O�1ä�f�����ج,xv�8�"ON	�!�2���j�'�q��Mr'"O2�{�.ΌY������-w� �1�"O�Yr��M�X�4�À%R{�~�!W"O ��e���j�2c٤{v�V(�y��=Y�d<������:��1�yR�_ov�Qb4
ώP(�e�2NƠ�yB��Q�� �lXSf�� �HX8�yb��m?��8�!܀��q��"�y���*��! 2IE��F�� .W.�y���1G�s&g�T�줘c��+�y�
�/m�H�ʖ*\�N��=�T��y��ϛ$ؠ����6�Xik�Ő��y��@�J��ف6�A��ك�
�+�yb���u�`H�@�['B�r�х��<�yr�T%.Br�ytf�@�fE���y��:���4G��=Z6����C��yR�G5n��윫/�T\vK�5�y� D�6!��)T+#�(�"5�5�y��Ue�����A	33���U�yR���x@\T#",�2|��	c1!ҝ�y�_�`Ϛ�PfG�w�����n���yR�L5h�\�X��6t�T����<�y��X�G�:�٤���k�Yے��8�y�囱4P���k���Br‣�y�
��s]4Uk7�ͦj>�Eqaa�yh�)|*�KG��b���	��y��J640)3i]>b�h)C�JC��yn��	g����B�\��@]p��QRpt.����jv��&}�$}�ȓe���'�Bvl�"���p��\�ȓ��s�GҬ(�@݈�L��8|�ȓ*�l��K��4р��P�f�d���)��q�%�!��I1'�����ȓR}d-z�e�1��B �Յ�)��~B��a��n8���D�+R���yF,�4�A�m�ĭ�� P��ȓL���-5/Pi��?8�����S�? p*�kX�pi��$+���tY "O����%!4�ĥ�U���y��"O|M�'�6�d�G
Z�!��DK"O���4D�'+F�0:0���Y�@��"O�p�)E6	� C�/C�pd<;"Oty�¤Z*_am�&�H��
�"O���6LI�B�8�kwKL,qЊ]�"O�H��n̋s�-�2.�|���"O�P:g�C�i��5BfKx��8B�"O�+� _ f�p����-< X��"O�{7*�'�$s��O�k��8��"OДC��/Dd\A�@(K�V��p"O��a"aO�e�DAa�ӫt�\��"O���� O&����N��ԃ&"O��:C��=���3���iZ�Xs"O��a��	y�ș�$�&gYah"O>�˗�K�b��5�r�{�x�$"O8`���
�(�Vl�R�t���"O�@tDLL�ׁ�(�:a�"O.��Fm�P��i���YP>4�g"O�\VbWcY�ڱE�4Qz�ؒ"O.L��,��A�t���� 2�a�#"O������\=��sʵQ�p���"O��S�+�� ㈒v`*���"O8-�v��+�l��q�ˬZ�]��"ON��Aی;~>����tt�@��"O��rV(J�1�J0x��W�S����"O�%X��Kɾъ�JuV�!"O��.�X��hg��=�uS�"Oz���hݥ�L%��j]7!�m��"O��s��88�f*�>K \��"O�T�gDm����*�NduZ�"O8���+P��Hٻ=�
�i0"O>�p�C�H�EP�zE��"Oj͒2�Y�<��N����M�#"O�kpȞ"r�$��0�Z�B5"O�H��HS�`����H��D�%�%"O�H��&�ʐ�gJ06��A�"O�ұ897�hK�H˭-�<-jg"Oj�u��[te���J,6����C"O���U�
�:���n@��^��!�X��\ڠO�=���Ω<!�$�в`�R�{`�冚r�!�$�=3pr�H�'!d���E�!��5yG��ZWlJ1j%:ɓ��)�!�,%@��a�.W2o*m�cϮl!��-� !�ID�TEKB h!��:�.�J�F�$���!�!�/KO!�$Q5��
��E� �"�Io!�$�`0��"�ŇWjl���L� 8�!�$WH�A�4��vb|"2�ϱm�!�$��z��Ijū[?6�F����@F�!��?0,��D���	��`KP
S�!�Wx���Oݸx��K���s!�V�H�ʽ�ǍW�1�WD�Y�RŅȓtYpV[�X���]�=gz��"O���<,��ts��*Yd "O�l�!��u�2]���Zr����"O�X�p�T�А�I���6WX��"O��I�/P~�Zf)Z�V4�飒"O�ٰ�KE�p�ֈ뱡��%5�b�"O�8R7%�a�a��l�X�K�"OƝ���r��e�.c���(�"O����P�h��]j�%ХZ�\+�"O�  ��.G��\`Yp%�:�V�j�"O��P�S����X�^cd��"O
�Ru��;nܜmb$�K�aPI �"Ot�j�DQX&ݢ�h�0G4�2"O�E�V�+O�h��(�;6,kT"O<���Y'�h�j]�C��z�"Of�c�J�xV���P�B��m�t"O�h0׫?_��*r���ޡA�"O��� ؄OB���G{Æ8&"O�q���@�p=�CU�Bp��"O6d��o�U���J_zi;A"O���wĂ�f?N����բM�9��"O9;å�lf��J�*`�"OF�� �u�h�MNj�Թ��"Oj���II _4+lȒx�b���"O"�j֎�&r�P���j*>龜0�"OzX+���[�r��c*� 3�0 �W"OhaP��;`�x�wHת�ơX&"O(%K���JH��j�$_���ِP"Ov���ᗃAJ���Ė�j]�"OT@��͋VXƠ�`D B��"O��3`��ht�$�w
�t��"O&��C�W6�c���7'\��"OX�ˆ�W !i�s��1�����"OFł��qu��z��˹TF0���"O��y�`�9�1��_�i0�"O���d��jj��A��g�d��b"O@��S���GX�y֤�%p��-Y�"O��k�oj���Kp�2l�P��"Ox�)P�T���92�G�vpR��"O��8�,H+��#B�H�3S�	Cg"Oj$
�;"��AP�4A:��"O Y`7AV�@9��SE!�)Z6"O�a�wĈ�aKHxs%@E�и2"O���g_;��$�d�^ Z�ɠD"O��B���dБ����C����"O��QR�H�L��Ҵ��9}5��8F"O!�2���X�YR	5SV��d"O.��ň�<cD,a@	Ok��"�"O��I�� �\昤i�jK�)�&%�"ODir�*� Ky=
vIS�-T"O����IX,�b��:q��l�"O�Ȋ6�Wx�(E���<� ��b"O��)#��5�v]`4�:ws��I#"OP��r�_�J� S�@�Vq�X��"O����
�5K#m�Mk yy4"Od��"���Hb�y�ś�GW8�D"O��y��Ш.�ɒ�!E_)��#3"O$��7�:{
�X��@X�9  "�"O�dif#_24l {���C%��3�"O<���Igr�J���(."�YjS"Onpp� �LDx���4~��t��"O$�۲
�AAV���&����X��"O|'��0(��kR�Ʌq�4�"O9Q�(T�t[R�[фԩ pZɻ1"OH ��M8[�$$��X;�P�"O�y���C�$��t��
5Js��B"O|��`.M��2��4
�[F��@"Od����0�JؖIԎ$�8��B"O�X�uL����0D'Y�,A`"O���"hN�"�Z���'[%8��<{�"O��U�p�XT�E��jĔsf"O�8�V���H*�9��&@%_m��Z@"O�x`��Ǻp�MHScF,j����D"O� �����ʓ>G�ʡ��{��8�"Ot�����	�B�YvG�fdj���"O�E�s�	��895��v��|��\�sTiǢL�*)��Za��5�^#�,��*1�`�o�`��u"A��\�Z\�\֬H:$,��ȓ[`�X+֬֨NJ u��_Ѻ$��/Ǧ���Ƿ5Ф9� �^���0�ȓ>q�Ѱ���`E��h��F�@��хȓ tX��K % �9B��\�8p��8��Y�����3�Z�OM�M�� �}(����AI�1C�$�]����h�gF=�����Ƅ$�Z@��!�`�	�0�8� ׷_�T��h��${`��A���X�S�`=�ȓE���o-��9P`χ�	[�|��@���)����(B��O���ȓW� �W!
 �H`��w�֩��QF ��UNPj(�3%,B�$<��?��ᣤP>l�#RʤU*�p��,�K�9g'd�#f�G ap~��ȓa�h�%LZ�`7F���&�V�)�ȓo ��`�I��u�<�UM4bN�ȓv��jM�ZD d��#�k�����& u�H�,�l��X;P�q��K�jL���΄f]��SDAE#1�܇�=~hH`f�2�ԋ�,�3^py�ȓm�p2r!��iǴ �V�1�A��A��ټ}G�ٲ�)�('���ȓB�:��lV%��f��/���ȓV�j�q����5	Z���F�%�b}��<�r��m�E�J�9 ��=fՆ��lt���R���H
`���H�ȓ� |���e7�`��!��2c����eD�,I�`��bVbLɤ��i��ȓR��Z��X䂝��L��&Є�)���(��X&	�$5��Ê7J`~u��8�XҦC[�k� �dם&*.e�ȓBhz��GcЀK[t��fɊ�N�(�ȓ���@�%j��sW
T��B���$�V(3\IW����\�+Gz�2�'&z-I2�@� �Tm�&�[�i�E��'{� #Վ��3KZ�r����y	�A�'��uY�㓮N�|P�U��w<.�H�'�ļzQ��� �6�B�ǋD8�P��'���cӶz����'��8;�'��A�旷-�~�S��L �K�'E�5`3�/K�f��@�lha�'�Jp����1l����EZ�>��S
�'���G�Fj�{��T�;��x�	�'�\u���4S<H�hҝ3t��	�'������\N�9J�A2�Z	�'��pHrkW�"�@P��.߂�P	�'�ȵ�p$	11�~ 07̔�tYb	�'o�H��-�9�B�eߛZ��	�'IF�2���!|j��Yvl��	����	�'=(I�%̗�w Nd��{䨰	�'F�����]gdS�"N�zu�5��'B�(��mT�3��}�Պ��zg���'�5�`➅Y�U{��Չw����'%�P���M'+9�����x�,#�'b�,�R��&JZ��"��?v�8�'��%���zVP���NlH�K�'��Qc3NG�~���σm���� &��a�������K�k��ś%"O:QA�9H(yа(Q!o��-��"O��@R���Zs��hb&��F�$��"O"��d�Y�.8�G�B���`�"O謉�N�@��7�����x�w*O
,	�`�
{�^�����JۦM@�'g�щ2��&��c�!��l)�(�	�'V2�Qpd��^���ØL��*�'F<�0��C��J4 !ĄK��}0�'?U!�B�4"*�b�KW�=N��*�'�ޝ{Å�"l2L�4��?6�Ժ�'���"�\�Lk����o�+{ްJ�'�bu��.�+��F(:pae�T^�<Q&�7&A �T��<k8�3+�Y�<�1��-�~���1"��R0ΝY�<�҆�+,��$C��0^��y"���W�<i��J>����S,#� }�0)W�<�6i׼u�щf���\@
�B�G�<ICZq����Uk	�F$2��$�Z�<1��:1.�u�F��Yl�����Kb�<�R�C�8I�vC��F� ���\B�<�4�[��԰D��:���B�>D�8�f$�0*hk@b�#K� Ԓ�;D��R��4D�u��@�yb�U���:D�� 4��^�F%�@�\
���BI6D����K�7�u��K�,:�����2D��*0�J�7�$���M���z��.D��Ka�ܯ^�^T(��S:W@E�-D����;I�J���-��C���D?D�`Si�r��p �v�ʹ->!���!`;��5\ ȭ��)�!���I���Y�ѯ:�ŀ� ���!�D+FE�I�D+I�p�h�&���;!�$��Ƭ�Z2���'�!�Su/MJ!��<,"�Q���@�@s!��M&mI��Y�@�DY�j�)Z!�$�!�0Q��`C��4��*ʭ=!���
����Kk�J9�W"OZ(�)���
�0���_�L)8"O$�z���I��c��/S�(&"O.�!2��(w�9���NԶ�u"Op�+�pG��1�/��$��&"O�h�U�Y�q����� ��yi�"O�����	�\ll�d�ͯ4^(� B"O8U�&A��\3%kT�!.�ij�"Oءsb�j2,R�
�vT�C"O�� rKXV 0(s@�S& mxԻ"O�|`�,�H�
���(7��k�"O�y����	0�)�V�(ۀ���"O�����[8�p1Ja���J��"O^\��)�J}�*�.Z�ty�"O�`ǩG!eIܙ���5=��"O����b4\�P�h�-�ld˵"O�C�jսSް���M��#��ͣ2"O�hP M�D[�(p2�S a�����"O�4��A�-�h�.��L �b�"Oh�.�a��h�7'0���g"OV����ًC3�E+Rć�$H<��"O�Ո�ӡEGn��d,	C��p�"O�xb�[�Y�H\`!,�{<t:�"O�ЪĞ:NiCt��$.��5c"OZ�j$~t9���_F�0y�"O,L���F{����,�1:�te{p"O^l�%n�%�}PQ�"G�$E{�"O� ��C�"0P���5L�-I�"O2a�^Y�^�@e�еY�"x��"O�	a�BJ�M�9���G'5w&��g"O����&^.qb�±G�;IF�C"Ous暶E�.	p敷"�ة�D"OF,�%]T���t�߃V��Y�"O1(�/G�5s֩�2,��͸T"O�-av��Yv�����$<�"OPu�u E2i����F	4�F`�"O�(p�G���a�b��;B�|X�"O>\0q'ިn�����
�J\d�:"O��Rh4HX�7�Z�-FD�27"O^Q��b�2v�P&��8by��"O0Q&�@�O���k΄�7?fy��"O�G�Wg��I�C�o ��3"O�� T"�9��p��Dτ:
��0"Ob�q �މ<^ru��$*���"O4���a��T�����H;D�C
>!ҵ��F"&��g8D��زE��L"ޱpq��q��h��4D��c$��4
����,43�<k4 0D�ĚTN��tN.E��GE	N����3D�����¿
�~L��,�;VPpp"�3D�����]�*��=����37Dh@j4D�pZE��Z���X`�U,��X�h1D��Q�
��89t�!D�i�&T�T�0D�X�2H�jO�Pr$�ÖP�|�D<D�T	��2�0=҅�æ3J��x�<D���3� ���yq�b��"s��H'�&D���� ��s�d�DbϦ��R�8�VB�	�6ܱ`/�U��<j钖~�C�BPH+Q���UX�c��hcHC䉩QAɶ)n"���Q�8C�	�qI:�r��x9܀SE���B��{!��:3�;�ة�Ã'~ՌC��|�h���;� ��ӊC6Z�C�ɱ�I %�O7q�����8U�C�^i�L�#��>
H�!�)��z��C�I�b��x�p�S� �x�D-3c��C�	>N��U�]�ݲ���:c�>C�Q\�ɯ@��}��OU � C�I7iFY��N�ny|ŀW�X><��C�	�M@��H�3 *�9¬\<��C�	�1��)8vM�N�9#���w��C�6?�d����?��iR����C�=�rI��e�����U�c=�B�	l(�R�hD}��<�^+M&C�����烗M���b6�'F}C�I�@�AЕ0�Ȉ�u�ܭ7(�B�ɢ9���r�4f�Mg��%�C�.4�R�� �$��z3��\A,B��!k^���S�U�d�V��$a̪�B�I'5�0�L\#U�&�Y�L֋o�B�I�w�$�Ca��Z���^�)PXB�I�O�|�ք�9A����d�\�|�C�	�ML�5��G��BY*�Bj��B�v�HhV�Pv�	B�e���pC䉑��i�%/L�Ze`U� �B�ɰm�Ե�����j����k�R��B䉂x����2

�:~�(e
-<"C䉩(��0�Q�� |�L�C��T��C�.?��hE�I��0�刟ak�C�I=W6�|[�B��L)��"�#����C�If#e���<CĮ�������C�)�  ����a+QOB�w�v�"�"O�8	�M�,]	B|X4�X|8���"O�H�1��.>tx�r%��.L���"OACp'�z����)D��"Or���-�0���Sg�$�|$ۂ"O���"�-|*Й���Du���"Or�x��F�*?�i�1+�P�x�a�"Op|�CbО-�Ԫ��N��d��"OH�(M?�p��F�߬#���ZT"O\�1�& 1,�\��'OY,_�����"O:���폡@ zY��=eP]�R"Oj��M��D8).�SY���"O, ���Ѹ0�T���ݜ ��"ONY�C��mԍ�%,�i"0H�"O���AE�Q��I��؇m��2"OP����8eꘛ�^�E^x�R"O(!��3y�Z��0M�	3Tat"O�i� �X8h:����H$�wG=D��FP�l�<}p􊔸`��4$9D�pH��]�j ha ���so� !�8D��0#o�xI uI�Y�^���i�6D�x�!l�x��[��J�6D�<x�[�G2e����H�M g>D��A$�E+M���'ۅz����¨6D���1��'}�ܡ�j�9����C7D���������QC׎I���C�b!D�T��G#��y�U�ӹ#7\	��=D���T*\%W�� �I��T[��f�9D�l�'���>�����υ)����L7D�x�Xe�l8����3�aX�.7D���%gC��F HC�-J~M8�4D���5V�t��q!^�70hEK��2D��� ��Ϣ$S�˝;0�8��GF%D�|:b�5^��pυ� ��-�Ū"D�Tjeg_�->�ʕ��]+܉�ª?D�Pa5��i>�@z�"��ĕ���<D���招P��Qu�@��=�F�%D���wH��\D�X�Po��I�VY�@N(D��kf	I$�r�! �> �AQ�<D�Tz�����@PC��|"�m���9D��qveӹ>�B�4���� @7D������l�q,U3
���O2D�Q�
J?z�The�F���@@r)4D��`�)F�E�UyA��/��Ԑu�.D�L%N

Zt�yn��p4M D�8h��m���E�ݬ@�r<i�f1D����P1��m��nP�C29��b0D�d��$�?!�f�bƎO0����V�;D��C�m��oM!B͠-�.,sI;D�l�Bn�w�lZC
�{��d�G�.D��Ӕ�L�Gd3��Ǝi	� 	��,D���倇�j�P�;���{���-+D��I���S~���蟮p,]B �%D���AӪw_�E��a�a/4�� $D�D�C�����jR(\,z� ���"D�X�0�5m"���)�>M$`qg#D���P5J�8�l�� 7�aj?D�d����9ec��y��/c��i�a>D����
�gӦ�ul�������:T���6��.v܉��ϵ���"O�\C NW�*w��3Dn�/?��8��"O��94,�1	{8����,`z8�Sb"O6(�/ C�!9�aZ�8�"O� �k)q�9!1Aب~�Zr"O� ~��竂�0����iߚ9�~��"O0�d-��t@j�Wc�;��g"O�p�#�3m�i��S�/)�a"Ox��,�����jw\���C"Ot��cj�1AA� ��%,�t}	$"Oɩ��[&^�69��B��z�nY�"O�X�d+ȫo�x0���!6�\Yy""O(�xP��(n6n��%�2Wb�]��"O^Uñ��~�6�`���5rWHJ3"Ot�UJ,.9�D�4?(�r%�G{�<y��߰}<P2.Z�^�pJ��]t�<��lԙmEP�b�A4�����v�<q5���(���e!�;�]��Xq�<�b��@خ}k�Kڸ�x�pҁ�i�<Y 喇%WLp�	�Mlx��AoUk�<���#)v� �@ߴ�v�ī�L�<#i��+��}�"�۲j|�87��o�<1S��#iA� ����1���l�<1"�<q�JH��ѯ � 0K��Q�<��bX:�nP3���|�d!E��B�<iƥ�I�<��j�9\��{V$�}�<ifoT j$  2Bƶp1j|�&�Uy�<Ad���o��1�4Cmn���L�<Wf̒s,������c�� ��Kb�<Y0e\�u��ݻ�'L'�5kdjGS�<��/E�$y�BȉlH�H���T�<�$nO?`�x:���Na�0Hu�R�<Q�a��}���E���}�I��]B�<9��SF��h���Am�)#�B�I�#�a��O1Ur��B
�/3PC�N���NU�E�y��k�6ODtC�I������5vˑ�u{:C�I�D�
1C��rʲ�y��K�NW�B�I��a��KU.������T7�C�I�Y��P!Ҁh�^ѨBoІ�C�	�j�x�ys��8~�x!�gܶ&f�C�I;fujy�2��WҨ�R!  6}C�ɐCUT!Kc�A5��%]d�B�IY���Y�BP)��[1��;<?DC�	3�F0A���#UŔٚ�JX"U�nB�I�^:������b%`֪e�@B�I�U�$)it�L/ ����'Bd�C�I0m'�h�'A�y���9pH�]�C��S�µ��6V����f��C��,l�\$�G�� ��F%�o�4C�	�P`��
�%�Z**�����%7nC�Is�t䃕`ҝ�"% ��ň!�JC�	�GǢ��'\��lfj�YRC�/
�#V�
@w��S����xC�B�	)Im佩W�NƭH���;qC�IR��0�g�V�7�qS1�U8H�C�	�5 �1u��L�C�	 t���cv�6b���0�?<0C� �p�����2�)���(]��B䉺8�8�:	����L*�%ݢJ��B䉵 -6m�� I�Eu��c���eC��%���C$�� R8QQ��j�.B�[{�͠%)�GY8h*���&XC�h�!&I��B\�?Fh�'��y+�K&�h��I��sI��I�'��E�$�Q7T���U�nrM2�'�M�+�:�zʷ��m�n���'	��:�BU^���j��'f��C�'m��d(0�9C�R0]Z���	��� ����c�d�B�Û�� �$"O�dI���D��HJ�;n��{"OB5��f�?]oU�d���^��c"O��c��F�3�Ԅ�7��'�n��"Obzr�'d#�T�! �^a���"O��I�k�i����4:�()�"O�as���>EE(�9C�!T�ެh�"OXp�Ѓ��*3�黲��4 �g"O:YXb�ŋC?�YyB��7�����"O`4��9���ָ)���"O$���������&aa�"Op��U��9fSv��:�ơXG"OX
��Dw����Ǣ��仆"O&����M� �B���7E��<�e"O���%ʯC!.���\�%�x̓F"O e�r�& �*{�`L�X5�\3u"O��#W!A�d�M@"�N���b�"O�	�%k��>�t��ΐr�!�$�5j@(C�[��MCb��0P!�$#"(�V��8��2�ÏR�!�D�Z&LE�&�V�$�lC'�!��9!6�˓o���m�[!�d�-�2QY1B�.�����l��t!�� �ޝH�ƅ�:a����@�  �!���7˘�Yc�&z,Θ{�f�!򤙚H��́�ׄ1j�j�U�V�!�$ۣT|~����
�i,X�U	$?=!�Û���5hG�AٌP�3�*t$!�d�0R300AG�<7,d�s��A!�$\N(P����X}&���I�Wv!��Dt`���釠hb��E�,!�P2|Y��� �xN��s�$40+!����o�`U������eݘK��@�ȓ^�t�[���k��M������4�>�[0N��d�ڰ�Ү
Y����ȓf�
���P�Ԏ,)::ф�-��ZU'E��|�c,+:1�ՆȓZy���RdV�;�j�RQ˽Gp$؇�i�� ��)ؼM��H�,���"On9����\��b(��(�h�Cp"OXz2�βq�.}�&JE`�4 �"Ot#0�ۯ^ �W$_�_A��x�"O@��-TH�6�a�S�w.�j"O(7
��XD����m!(
d"O��P���
��"So��*�S"O�I�D����h��H�r��Q7"OpAE�HAL9:�̓)vrD�0�"O��!�!2�a��b	,`��5a�"O*���ݶ �$m�!��fntM��"O�	cрKw���R��s�tp4"O�]��ݲkp���b`�h\�Lۢ"O�ôd	�}e⁒���'���q"O�� �"E��q�͜&͊ ��"O�tXa�٦n]8��$�]&r#�y�4"O�����<��DR�
D�~�`�a"Ol�y���u2��{�)�_�Y t"O���q_�qC�4�a�­cN���"O>��f�\�v��+s��2::<�rt*OH*��("zp*�#m�8K�'�,�:�n�]�&��f0���'�H�t�!�^��5��,b�X��'����dǨM�����:I��'}��)T�V��q���!Dz2�;�'������ �~���iD�4|J��
��� ҕ1 ��l��o\b�y��"ODa����!W���ZOŪ$J$L��"O(�
tIצ_�`T:�M_�>,�d!d"O���W�ZOP�z���6t�xF"O�!�f��Q�� !�	�'"O����D��iIGl�i����"O�\`��Ζ
U��	7+�2L��"O��6���"݁��Ć0��"O8d���R#��Q
M�ZԄ��"O��HM��]��pfHP�b��I2"O���,�+53*=k�G
/u�̴[�"O$hC�l�'Z&���>�:���"O�D��EƐhN��$�]7 �\�+�"O
Mk���:� f�@q�5"Oh�
f效<x>�Z��� �p�["O�� �K�;0���m�"�sC"Oh����:nZ���"V)c�P�g"O񁐆�5B���cY>��I�"O�d�b���T�2���s�,I�"O0��AB6Q7�ɐ�&���	�"O����2[�`P(���P���"OT� �L��W��Wd:�x�"OlЁ�08;N�f�� B2�ykd"O�=�$c�8b�ؒT/$A*A+Q*O��1��	 ���ad��x�'��U�$o�V.�$r��7hf�i�'���Ģ�qD.`�I��YI�'9l-��Y=��� L�*�jI��'�j����]�ti ���n.���'�H�;P&͸=l0*0l�jp���	�'���q���3
"8B&B�eȡ;
�'���W��%Y�dQg,��\��T
�'�4@�G�h��@Q���h��Ѫ	�'#^T+��v@���t��52[&xH	�'���FI�,Z�@�D�(�� �	�'36��Yc�c��D)P�d�	�'��LH���5FQ�di�w�|,
�'�\�٣&ٞ�ZahD�_�ok���'|đs/��xP��G�;ao�E��'P,�Y�D�>Q`�H��L/l�pp�'� ���H�?�`3f�\�`���'�64kI��f�T�c)�'S�Zc�'�8��1N��<X�#f�P�p��
�'#�y˱!�p;��9�F�)C�Z\:
�'U�p)c�*hn��X�(Ԑ�\Ղ	�'��-@�2w�R� 'V3T�&x��'%F\�'�
�o��;�-4R���)�'iְcҊG�o��q�CAѥ�`
�'neB�/�B����&+5r �
�'�("�`�0'~h(�O�	 M�	�'��xㅩ6|�ܙ�HfJ���'$r):ӄF\)"TZ�LK�s�'f��c3KάEdܣ�-��7Μ��'2�=2Nܩ	&$��e�9��	�'�����	Շq+B�Ö"���i	�'ž����r^V���n�-B�
�'�Mj���1w� �ەeV�/���
�'�"P�T Z -��)�(ј'K�i
�'�� ��@�����Ǖ��"��' zM�p)��%K�/Z�~�%��'��T�m��=���|_d���'���� � ���yJQj�'��������r��EP1v�����'[����"{�'�Θ@BJpZ	��� \�I�:�tU���#}t�bQ"O�����ɟ&)�5�fS69�La@p"O�[#�Z�:Xc䏅2q����"O�p�+A��b����ތe���"O�(2"��4g朴I�d��l�*��U"O 4��/<��!�S�מ?�,s�"O`pQ� �cB�H�㌾/����`"OFm�u�C.:t\ሂ�8_f�1"Ol��w"�g�PHӀ�X�!�"O��)3��6�A6�(}8�@kQ"Of�� '��:�����@�E"��G"O�-i0kV�C^��N�7p&L�ɶ"O.�x%�� ;�9�,O�0�0�%"O ��R�� Y���ٱE��2"O��
DA���z��:\��"O�`7"�G2X���ʊGᶹ�"O� n�#f�,��LWi��sU"Ov��!��<���Z��V��أ"O�="5�&�,�����?���"O��A�2qE^�Ie �	���!"O޴�dᇧv���,����"O]*��L�8R$m�w���2��02"On̈��Og�
\�&�K�X��"O̐B�!�	X�n	{�F� Ii����"O\����I/D��0Pa�I�<M 2�"OTx8�MZ���y�CӊV8�A�4"O�Ej�l���5)c�0��� "O��Pׅ��Le�0�u�@ ��r�"OH9�ߖ.z�*Ն/A��%"O6-�%
a�%@[������"O X�IҒW��p��!=y��
�"O(1�` ��lĀQ�㪘�a�Fl36"O��A推&�n�C��E��bc"O� !b�;'4��	H_(�J}I�"O sD+ۚ..ܜ���	�n؛u"OJQIa�4��� 1��!�J��'"O��1��hx��K�K�7O��p��"Oh��jF�;.�����~���a�"O����٘��x�"�@�V*H��r"OX���B܋@:� q���Ǥ�Q"O��B�#�=,�t�+BHO�Q�ZJ�"OtHCӌ�
w+���I�+j���A4"Ox� g%��±�����@�"O�d�R��Va��3Ď�k�,Ya�"O\]��,�bB|�$c].P��`�"O��r!�^�|�`��Q�A�k��sD"O��;c@�/~:��t"#�ȹ�"Oxm���[��˓���~<��"OΑ��
T�a�Fl�pC�V�<�au"OP��9�������aI�"O� BB�_̨y�A\0W��1C�"OP�g�5x<��[�o�@�{`"O��w��+�ޘ p+	�1u0��"O���P"��9!l��g�I* v��h6"O$ �2@�$gC�CP��>�0�"Ol0���>Q������r����"Oh)�C���5x���K��yr��v��q������;��Z/�y��n�D��B�
�������y�aGX�]ڇIӈ{��}22�W��y2�T>5��V���l����+F��y�ǧ3�x2R�F�9��D
�-J�yr��B5e���Q�^"�aCW!���y�F�Gh�j2DQ�Gi
	�VZ��y
� � iD�K�'#rGR?N)�@�#"O�����
j-�QrW枚t����3"O���q,�-y��9c��;�4]��"Olp��JQ4<��{#�!V�;B"O:���O�����]|`P"O��#�E �n��qY$�_*W8��3"O���S�D�O�t�C3��m�1;�"Oܽ:g�H�g%�-�ad��?j� Ð"O������"�����^Z�{D"Oh%���ōp���ASW(4K "OJ�jg 8'�0L@� �&���"OR����C�%�,סV<�6]PB"O������/�(���ƪ3
 eC"Of|c�f�!=�tx��Z(�Fl��"OtI��M�+�\Y(P�S2T�"O�}(�%A<W�ѓ`��0�^���"O��k��!�^;�!�)�V	{�"Op �Mľc���b1bλY�0��"Or4pQ��p�T%F�=m�哶"O�a�CjVzpԨ 5.�gl���#"O�}ٰ�]"�l��Y̼��%"O��@b*X�-'`�q�lK�g[ �*"O�-Q���^��WES-]p��"Ofl���#!(�1�`��7)���"OpUAU��b�LԁWÒL��d�7"O�d)�
	s���I�\�6��U"O0�!F��Q��y0g�	�v��pi�"O�˂�A�q�98�ڸB%�	�u"O<)�b�jlv=z�%K�9��x�"O���B��k�L �bK�=��"Od5z2�B \�v\���M+T�2Y��"O�M��&��rW��0�3�Խ�@"O �q&�ρx���P�Юa��I�"OD{Q&\Nt��!�sa���'"O���~>�qk�N��(���y�
��
Q��"��qQ����fV�y,���屒�֣s�]�b�(�y"e͎
+���F �^|������y�Ö>�*PH�N��Z�t�ӕ�P0�y��n���p ��p1JuA��y�䞌p�`��T�Ѹ)�\���`D)�y��*z��R�0]dU8����y�
4FM���b�ʴ�iX `��yRo{����A9�
<) ���yҁP��U�}���xp�A�yb�
NKJ���MS�{j�3�	��y�S��d�a�J p�B,�-� �y�˜	]�EZ�lިQJyxA���y��Ϊ2�^Ȃ�G�x��UK��yR#A1r��dm^�#����$]��y�/� �R��%p����a�L�yR�������\gV�*�fJ��y��TJŸ��JM9>����y��ǐT7�D�`b�v�2-:���2�yRO��Q˖L�G�nReVD�y�m�G���h��n�(5�E�\��y��Oo �D`-e�ȩ�tn���yB �`��h�p�O	c�p�P4˟��y���f�ؤBCD;p�̡
$lM�y���n	�)��e)d2�c�[0�y�K�rkz|�%��p�΀������y��h��X1��Tk�|H4�@�y��@�qg6��g��{��e���!�yҪ��z4��s�Ɖ�V@P�Ճ�y
� $41��=�^9�Ŋ��<X�"Oa��\�.��I���QM����"O2բ�#ۊYD�k3���a9�%�w"O�pҳƎ&,� �%l�J�̋�"O|X��-|�ZL����5�p�'s�'l�11p!J)0��¥"��TQD<�	�'����]�L�P(��H-Q�r�J
�'����I��a @̪�҅6JŚ�'�T�0�ϒ�_�t8z�m�!+�Z��'�ў"}:`*�5�0T������~mɠË2�!�d��d|m�%lV��P��Bӻf�!�Dʕ`��$�G FD�j��cAԯN�!�D�,�|���cʍ[����C�#���x��)� %��
4�Y5x�Q��hi�<��-r��	� A�h�$���[�<٣���c�h8@��Nm:f��s�<yUɈ�k�ީ�Q�Ç J`��P��y�<��O/<��j]�EB�A��`�<yƾup�DH�źW��u���\u�<a���^�N�yf-F� -�Q��Vs��hO�O��}��@�6VۊUy$��'Y� �ϓ�O�Q��n��T��B@������AX� �!O�~b��:rG��.b	%�5D���`�`�h��J�m^� �a�3D����%@	����B�Kv��bEn�>-OȓO�3�� �/�q���;#5���t%L��!�dˋpƸ�qc r� .ٺh�6مȓ3�2e��;�ĝ��!�6M�l%��L+�tq1C�q�Z�@R/@��D{��'��ܨ�BA�2�К��M
Zժ�A�'t� ���-E���8��V� "OTЙЏǪ[��a��A*��g�'��<a I�$���%�� 
�b���Rs�<A�0E�#˅&LAr��J����(O�e��': 3��K�5����x"�)��3p��1 &���2 �.y�O��=�~bw#�HP�m�s*NVJ�]�@�DB~R�O���Pay콰��Ń8��z��9!�$�O��ˆ����i��-"�8ۗ"O�ᰤ	��*v�Ż�BX +q�� U�'�ў�%៳Z�|݊� !#Ǯcc'D�v��zA/�F�I"W��9V9pb� D{���ˉ�=��`Q�fRw�Y)�E���d�<)�?�^1AQ��$�
�3s�M,=װDFx��'���2�ta{v���L�p"�'5��蠣@j�𩑵+B!L�r�M�R�\�|$��?eA�`�&Nq�ܠ�ԖB�!�/5D���/�qFzd� �P�4Z��:�3�	D؞d�p�SG�pi(�7�Z��0�Oe۴8�㇭G�!��qa���6N��ȓhڬ#S��n�N��P�;�����	��O<ei�(�4VǶ��u�҄!&{�"O"(�(M�"av|����'�&dB�V�| ��哫V���ӡ�;E��\�ӢW��B䉳9s���b�/T&-��C��>�
� ��p<)���8���&�̶�r��5��r�I�<��}ʟl�DU�#v��D@��K܌b�Ί�$ hC�up�t�c�U^����&�T	;j8�����O���sFW�`|i�sLe�
 ��Y����I8��=j��F��~��W�n ��J����'+���r��%��"p�X"	��
�����D1CHD=8򍠆�"����n�xb,[��% �i~��ĄȓH���YT	��V���׏L�J�NP��S�? Hhx�KJ,Y��r������"OnM�d�9�,���3����FQ����Ɂ0���k��aʘy�d�"��~x�ȋ3˯<it J+4�1U�\Iᠷ�N�'�1O����y�'�9C~��Z�"ڂԜ@�"O(���@#bP	�A½/�)��"OK�=q�*t)�@�{���@H��MkM>iד.�
!s��@[G�)+S�T�+�}��t�P�)���a�5c��W�r�x�"OV�§.��eB�d��D:hc�{H<!��4�t���!�MX���hH�<Qci�8@u8=� �\$8�,��fIKZ�'�a���Y�a�H���?}���K�ݨO#�j�1D�����Z0�l��3$\��F{���X�qY����ސ&��!�&b%n�	��HO?�� ��D���#E�@-fд�f�"D��q�\�7�f9�U��a5�h�$M"?y�Ex��� @�4]�vL	�`��`Ψ���	s?��jjΔ��WT&f��wF�Q�'axRF�&�^(� Ɯ��Q��cٚ��O��~:e(�.%vh25���/(�pV"Z��XG{��I�*��(Ó�M�"��'�-u�B�	%lJ@HӷM�5�"bH(��B�	aj<����,�
�R ����7�I#�]J�$Y�i9�B(��C�ɐg.l�V�[�-_����L�/��B��d�^xXgj2"�Q��?��=�	�'z1D���
�t��,����2ʁ�ȓ.���V2	��H�A�ʥ�'�ў"|"1BW�v��)h���
Hpmڱm�}�<qS�ӣP5�a��-
$��2��c̓��=q!B95+��cW# 7St����[�<)C�470Xy�ǃ�Nd@��Cڦy!ݴL�''��O�����+٠@�����?���fgǂ_a{����?	h�k4�&��I����a1���M��wKB��n�&x��PnF<�a��_}���׎��S4����סC!�Ќ:$4���Gy�Й£#��n!�D^�x��4!T���w�T����E�	I!�D2vV-B��p�)�0H6!�Dل,�F|��/9�4�Ñ�a)1O��I}�S�'u�&�{��P�$RШj��mpy��s^ �Ҋ��L�Ё*���q;α�?�`�'�j�8�T����7��^��
�O��ѐꛮ8�Ќ �4/����h��ў"~J��ʄ D�S�AD'L����	��p=��}�D`���WLٍS�N8Cw���y�NdCb���\y���F�ǈ�y��3lH*�"ϐN����b�"�y���	]nP�%J�?�($ ���yB���x����fY;F�J��gIT4�y�CL��kS�ON:�(vK��y����r
xu�狌 KL@������x��'�t��6���9Ql��ɩT-�M��'��q��Ǿ�ĀɃ+��S�(dz�'{����K\�u f#ȱ]΁��'�B���\8��hBK�6+�����'��@uA7k$q�i�'��]��'`��і�D��ҥ�A��:yx���'�$��` "c&T�d
=��*
�'�t���-J�4M� �
D:���'&0�\�@�-1#�K�k��X��'L��zԈb��9	�6�]
�'��q����G.\����W�9��� L�:�e�1-[,�H�jPYN@�"OXX���ݢ)r����<�����"O�r��ڀS@� �` �.FF�&"O�E��R�f�a���]�l($	�"O���^tA@L8	'�2f"O2��c"E�L��p�`�-7��y6"O�)��?R=v,i���!a+�"O��b��9޾��
� ҈<i�"O�=S�V^��PJ
+�X�q�"Ojd��!M�1pWi��O�>Q�"O�!8��K�G�A)&-R�֬3�"O�0"u��G�"\)�Bʄ8�n�{�'�*<Q��"h�@�gƎk���'���
��M�[��$�r.�S�n +�'v�l�&l$֤]�` ^-JƬp�'��� t���+��#`� �:�b�Z�'wā�Ac@ p�7ɑ1$�ZDs
�'��p8�E\8e��E��Խ�樋�'2B5�Wa
/D����tA��+*���'%�u;U��G˨M�#iԝx�V9A�'=b���W���w➡k�0+�'}d\�/G=}�Ju�7�5b�����'���y�J��v)t/%�b��sLKO�<� ��R�
��890M�S
BB�	�a���5%�(�UOLxB��q�L�#�)W�������^��i7*��l���B�b�IHƃ�.z���(���!��[����s���TD����B�!򄝶@_8Ԑ���@3J�q�J�"Y�!�m,4 ���!/$��a#B�u�!��<1�{umѳ[�t�g/��)�!��Z�Ar ��[<<���M�-3!�$ڙd�h�B���8�\��m߀F!!��x�t�I`�	s��a��&$!���9`p!��� ���R��Py
�*
�{��I
�,���ܤ�y��F�(PDT�3m��4B�8Y6D\�y����$��'�2��r���yR�٭Q�݀�
��-#�:�E@�y�$�.��$��&�j�CQ�4�y�M��w_$A�k��+5ZMٳP��y"��=s7��'Ü���+c,��y�!R�H6t�#��(pB�A�����y�l�	?z�x�EK�&�%�2(�y�ļn����᫈��&0�3��W�<���E�^x����l��q�D�P�<Y����Rɜ���^'=S<9�FO�<�E�+L������O24��Hp�<!�c�&K��yȷ#/ubz��E��F�<)!O2������xp��Ӫ�}�<��A�)/�T�Tb��,��I���x�<iG�Y�:,*��᨟�)�Ĥ���Uq�<�E�9�>�BND���{�Cl�<qӬ7;��ABL9v`���f�<9��	?W��`XFnӔ,1Xs��g�<q��7J�k�e���<[�)�z�<�"�--1���2��-!��^v�<��n+v���iKm���0ǜO�<��	�� @��.�$>�0�"TH�<q�A�캡��	��X��3�y"��h ��a	��s��3B�˓�y2gȉ}���(�P�Y���� �	�y"�Q�}'�r�G��]J�-ڰj	�ye�M �q2c�߶M'�m{��J0�y
� �p@�ْ]bZP�4�5M�ti{@"O �����/�Tu3���V$&�q�"O \�Ȟ��ܜ�4m�@��M��"O,5�q��7J����@̂�*�|lQ�"O
p�.�����M�1����"Oz�ҵfΰk����-Y=?���"O
�sq�	E"h���H�,�(SA"O�L�c�!Bf�I5��4uf\ٵ�'mVx��V�	:H(�JHC:�捹i�<$��C�I�>�0��-[�*Ǡ}9�nX hd�b�x)���ja����Ӳ%LV��-ީv�l0hUT�o��B��4���rnO�OCV �0��+N���yC�_�u���f�2�B��L�$�J��_���%0Us�5XP�)4����α�v��;/��I��m��k�P������i�d���.p ���#��H�ES�Z���H ��xk3��Y��	�t���9DĎ�j(��h�fU���C�	X���B�W�X�zQ�@��<&�H�O~E��b? �PX��K/� ��P�G���	��A��}�����^0�,0�BN4D�eMF!\E���6.�L�'� ���>	��M�y�����`DtIb�Uh<�feSE�i�T���~( �A��.R:U��D�J�vHk	�7R�c��P�b�:1%E�/�����Q�n�AŅ�,����=�� 2AI�#�P�sǃ#`� ��2�j񡛇4a�Ջ���$S�$�<��]&V�0�� �'`S�̀ǣ�*d�a�g�ޒQ)|���l�`(WkԞ>��E����9����O��s��'���E�,O�`�(�n�����9�%�"OJa[DMܑ?���W P��U�b"O����O,.%� �g�C�[�th�"O����jRs�⅂ ��*a٢h��"OL����1f<��3Ũof�%�p�I.�@��P�音9��ٳ���'D�`[���lY!�,���E
��K�P5y�ɀ.f"D8��z�)�'=��h��	�&A(�2v��z���ȓ1�v��)��(`��j��,5�ɧO�Y�4��>_`���
��)��"�EN��y�@��8��	:7H8d��O��А1���
7�����W���pOp�9A��<�r�p�C�??V��2W���*�F?>W�č����h5K�"����rM8ä	;�,�!�-�� /ԙ#"O�@��F�4ل�s��ߛQV�S��OFL۰��r3�5��9W��iD4܎�S��_�S����Dиf*�zt��l�P����-E�1�f�$�J�Y�c
%P��.���ɃA��F;�hX�^�d遡�1\��d�O�����0�����f��+�O|�y���,9,�2[�;�x�B�O��ؒ���!bb�����AG�ɡP��"q	�[B��}<q1�x�C�]�x�h`	g�6�p��͖�����7��reDys!KA�v�sA�^:���1�G�D�=���sg���!��4BV�7D��ۄ ڧX���"���4/e����ǺM�]�u/��v��H��&H*Kv�˜'���BW,��,o�d�ܰu�N�+�6U��f�%채�7O����I�~+�%Ȳ#[2F+�l) `B2��K�� <��3��OV?aEHފM���T>o޽@S!��)�|0GΘK�qO
���&N�6�I�.��l��� �)�X��C��iq�ы�-J�!�$ �����/
�lX�!
�HdpbB�>J�^� (F4�D��4�SX}���s�,q�gÇG�0��S���yr�WΙ�\�Jm
���������T��5���Ј(>�q�I�P]~P)�jī��"�<1z ����j���b�� �@}�c�0V�K�9���!��I/`9���	�'��W��(@)�����@�%�}���05�W��~�J�R��Y2��s��IBh��]�H��@k��l�.���$D��R�N�@@,`8�� ��> G�$��"�xPh�:O���HO0Y���=^7 �T�� |l����'t� �7`�+8U��@��kOXtI��g\��`�8�!�dA�R�taz&i1ܽЄC�o�O6���N�9�DI�ŉ��M��nE&�����|YB��f���lS<��|�U"O�����O�Bl|�{7
m��H����:<e�dkD&W�u���fMʴ�ţ��� p�17AU�U;P�PA�Յf�BtK�"O��(�$�$���q���( �4��VJ>Q�0L�"t�P�B �;@���8Մs���>����+k�5��,M_g�4���_��$S�-���cGұ82� q���*x�0Kv�B
F]�*3%K�%;x���k����	 ,�ēW���Y��U�/X��➈2�".IJ=�e�>QH��2�$ܪ7(z����{U�j{j�S�NV	hS���O�<YlZ�pEvp8á�(��ŲDc��1˾s�䆅7v�Ѣ�_�I0v\�'��'J7|�ݷs<�i���`80W#���C�I7>���2茝�Ȕ���ɠR�x]���ڽ+�������;	�$JV7?��	O�` �D��H�\C*]Q�!U7Ҋ��KRXH u��7g��!�ci��Z�2;T�ҧaZ�,(���7bI�eiR0Awa~�n�!8ܥ���*	m�e%����'�6��v��p�(�����Ny8�h��k�<.�\���:M�X	�N��y��7!�t���Nի?6ڄ�S�X"mSRN��X�����?�P��	��<qVa
;q��	��<z�@(���F�<�$/Y��iQ3[>!��O˅M����e��B�-���S���@�;4B���I؏!|L�����B��� ��<|O.�2�O�\¡�6	�#T4U`䇇=~sTZV!F�"X���SG�~�k��ax�rF�\�X@�$���O�l"��Z>��(��Թ :l%>����p���(��t9*ءb�"D����K�&k�$���P"�  �hz�b}�$ĸ�������Q<��A��D=�%���E(�y�fЩhf�����ʭF���GѤ�yR��Z=(���_��||P7�\��y"d�($�~\U�E�QD��S��0�y�S/G��0���@D(���f���y�b��7>>�8V`η;�|�S���y�q�(�3����4.@�8�Ϙ�y�`�'�Ru���U�3c��zcط�y�/"R�l���.�^(��U8�y�W"6L�)a�h	1/7nໄ�]��y���n�Zȃ�+_8�Ju�p����~�"%_���Pg�+\O�`K��*U���'B�3}+�(��' ��c�`8Mi�1Z�G
�v��T�Y6�L5h�U��y⫈	���iD`e�$kQ������$�	h	Ɂ!S8�>a�v��~~�6�X=/F2��#�*D� A��ޕD���N��6�|ipwE�u�q���
�U�|�S��y�P	d��]�R�T���qHR��yB�N��B�P���PD��rAiǮ�yR��0���y�Y��0=��D��@�ڹk��3�h�T�$g��V�zVB�8�R5��^�l�j��'�XC䉆7ƴ�`�ꅈ�4�R'�˭)f
�<�2FP4���H�哮'��0�JM$(s!BfU�X9�C�I�"���Y⍎'',a�dHQ/
b7��?H������s���v&^�~�fi��'RwN��v"O\$ GɎ�C2Hu�1J��r&"O��:%՝q��ö�O!��i�"O��򧫙(Kl�u���N�5&��82"O�+o	K��и
23�DlQ�"O����f0f����*��i����*OP����"@�P�ǕGM$t��'9v����9d�aa5J��>nz�I�'�a���܎G�h|���(H��
�'�&���/� 3t�F����)�y�Jܹt�m0� ^�<�\D�J��y�#�7{en@`���8��T3����yOڼ-L�(���\Vx
K���y�1DI��V��B�Х[1�.�y��O�)����!]16ަ�U)M��y�JO4��3�S��:�D��yR
׏KHj���"��BC*�y�'�>4�f�Z$���H%�"�^��y�,��#L�"D���P'��y�%б#��5�͋69�(��ꇂ�y
� FUG�&ci�E���^!%�T��"OLIi��҄kW�H4���S��q��"O����F+����fCڵZ��Ss"O6A���� ���G�uq��bG"OD��iѝW�\��A�!jB q"O�k��>llLx��K�F��A"O��1f���Y�(�� �á!��i�"O չ����5,��ԓK]�mb�"O\�Y�>:�8t��.`�`�3�"O|� c�4�Y��������"O�\����1	0�Bό�$�
1I1"Op5C�n� u^1䯎�����"O��2�ʖ�X}�e	�,�d�,E1�"O@U7m�2LL���*؆n���"O�U���w"Mq��Ƒ ����"O@����N�`"���OId��أ@"O�xC�I�4-7��B�f�Xd�%"O�yՂ�)�����É0��H�"O�����P��h��|D��@"O�uA�J
8A�ı��a׫X�՛�"O<Q�%��Y��@!��Et��tb"O<����������5ETv��u"O:��Q̓^P���)C�z5n��"O����� �(1��o*��0"ON4#`I�
7x�#���<*�c"O:����r�`YB�j��q��"O�<jdN��~���m�P�puQ�"O�����\�(�����@�"O�z��C<�}I���	>*V"O�aH���s�5��-#.����"Oh���eگaנp��8�����"O��e��8��u����!j�Dz"Oj�+���>-�T�ikS�Yv0�ȓIY�4���BNp`}!�+A���h�ȓS��=kR�e.TYh���6�����R�/�<�\���c7~�6��ȓ\Y��s�K�*�8�`w+��N��i��Aܕ��$^8O)�`���=Yc��ȓ�P���>�R�0�7P��ȓo�z�<iatUh�	Q ]����ȓ'�t�����dM��`hXԇ�E�����ȰD������<�&H��d,�\s�Lɰ>���3,_��ȓ4a��`��� %�� �,b�� ��C��Q�h�"V��ep�߯_R���b��%�&ύ0��3���*u� ����"ӧ=Ui�����G7��ȓUƑ"'J!X����+ʻ}X�����Z4���
b2X���	�#mL&��ȓ\�X��ߐI�Y�k�3�H��IH�A��)ھa�޵Ac�_9l���ȓlR������J~����J0)vd�� �n%�'W@����LW pb
���K|H�T��5�K�0�Z���4�<!�p�Ҵ~�b�:Ѕ�Wǔ��M|јd����3$	_�LX�ȓ%� \��L���d�Ba��lVj�ȓ�<ف��Ӧr���k��w߀`�ȓb��t�IhDԌs#)�'Z�`L�ȓ�t�`�`bj���$�mu���^ ���;�[�ʄ��M�ȓ@�f���#�
,<�7�Ek�Z���I�b��c�P7Z��8���4񦱆ȓ�!P����D�*%��:j#ل�S�? ���BS.���b
V$ќ�8"O�Ыd�F/��)���S�$�����"O���${�D
f�,p�"�K"OH�"`@ըR�b�6AaQ�@"O&!�6��\s���t	Ea�*�kc"O�\�C��1Ѐ���ma�)�!"O�UH��4����Κ�$&��"O�-�k�~��)CЮD�&AHS"O*�I�˶Q��� �-X�I�z$"O ��[R�)�I�s��y��
$�ybKÌ,��E���͸t�����M�y���)N�~� ��F�;'p�ZG�<�p=�1�N	]�ҙ�O�I�7����<ބ6"O�0� ��_n6t��mغ��|��DX� ��h�V������x���-|�,JUJݜ^�d���"O�$�'X<QN�e�e@��8�iӁ��#���T�`�pf�F�g��U-fQ������B�}a��[ ��d
)^�А�#7Sd�Ј���BaE�l7�@s�!�O q�#�="��P�t�Q�^pq�V�'��L��nP�Xdm�v9O�9�Q�X	G�"E�$�P�=�"O�I*�>F `Ua�'6��A�|��&3� �j�a\%0�?��[ ��󀡅�UNA)�.#D����dD.l�2���f�>����L�,oF^��k�<Q"`�1����	�7����0#��!���2�FI�B�I�u0"L���>r9�6!։=Sv�xg#CT
@���S�h։�#���6�ɃO.H|KP�;<O��V 	L)Fdcp�{��BVc	�tiJ�I5�}+:\9!e8D�7�ղMMd�R�K_�8|#��9�	�9h�h pBQ?�����*1�dC�d��	*�b�b:D��)�+@,�u� �V1cV�[�#�T�
L>v�;�gy�e8o������ȧ&�t ��L��y"/�xl:�f�2���iđ�y�̂�=�� �����i��@��y���-��P�J�;1�1��l��y��˘��*e
)2;2���"���Oh�����OD�����Z>}�P�#��%c�%�
�'�Ҹ��d�V�
�C��@�YFڪO���H^�f��O�>��7f�0{��D)�!��s�f)D�H��іY�R�h5O�z����&}�*�!&�"�S��M� z'�M<q���1�hϗy$$��S�$�O�
��3��1Q�h
,�ЩBC�	m�e����xba��"��J'�
�%&|����;�
!t��IB���~�o�S����HR��wC�(���U�iɖJZ? Xj�'�QxDW�~�6�S�)Yd�{d�'5pѨ�	�f�6A������TCW{�&�S��D $Wd�B"�7Eͮ�swdL�)��{¬�<t@Ȩ��@%Tc:u��C�W&��
��)*t��G��L4������x�b�(|ax""�'y�����%8bBQjԊ���'�dv�Xf�^�|��͐�Ɏ�������e��A,ǜ~�Ht��7zA�fA6s�vB���tTXF�	+�ڐP��Z�}��x@�F�Sj����-
�����ϑ��~L`u�Y�)��������\%:�N����\�.�-h#�ҿUh!�]�w�Z�c�A�WO(�r�@�EZ��Ŀ3�
�դ�2b�� q���<1�)@�RH"�"K�Je͈<B�����*�u[�����&\O~�2�ܕ,q��q�7%mP�i��G�K�$�:b�¢,>�@ �DE_x��m�!�'g+̬7p�a��C
�4�VN�j��*��F��j��s��1z^8�N|"�/G>P?h�J$��)w	��H�	F�<��N��X���z��S�s�ƀ0 oK8Y�|x�%)ޯVH0�g�L	�G�$_�X�t�\9~�,Y�%O�pVJ��#o>D��0� 74�2�iC*~�xrd��	"� @ ��#@�2���ɦE���D2
ʦX� ����K�{.���Qj���p=�2N�!�p�� O��(�f]�R��gm�C�	V�v�>p&lZ�-G�C�I�7F� VC�9M�l0�d�	_�Nc�0�4b�-Q�E�D
�qa���NY�)]r=���]2�y�"�8~gVD�$�,6�H(�BFѩ,���WF%�	C��~K$Tnpу_���`D�y
� \:DoI��
���\�3L�*"O��[�oL�dE����D��\n˖"O`��f��5w8�3`Ҋi(�"O�m���S�@$��X$�|#"O�;�(�a͌�pW�xی	4"O��k�k��`9���6��y�@�|ܓq��4K��L�ԛ����p���`(��i �]	�� $�l��N��`�&��(��!V>w�ni�P/KV��0g-�)i5sե�����$!;O�} �,�mT(�C�OT�B+�uE�,9b�(5��;�"O��{�/�5R����60z��>�G��3i<t�(�I%�.pQ�Ա1c�	; OY="�	�"O:h%5)_��
��P��V 2��R T �1� �j>�3��Z89-pX���-k��B���s���d��85�7��G�>i��ǧYZ�g�{I�X`�H?�!Q�Jx�Arn�$$׊��ɱn�>�yG8O��I*vC~ �����u���kg흍"cxB�I�qF p`��Z	��DAX1�N�'<��"l��f����S?97Z$���?|X�p������B��A6��*�DقB�.]�Ŭ�!J�8D�.}��@���}&�x3��TB�č�iζ]b��B�>$�h0ED�'[����!(ZZ��$L�p@��P�P{��D	`�:��A���J�����+.<O�I����.�ēt�JJ-�>-u�D!����u��d�$t�5�A%��\�f݅ȓz^da�7�p�,1߲x!N*D�0J�L��R�أ�n_:�p���*D��h� �a`2�@#F\�\P%c��*D��'�� [�`5H��ƹ< ���5D�$hDAC|���r���?A0!I��2D���wD&XI�[RG;
_>=�b.%D�LHeD���b1i%��:�:�(6d%D�|� �_� j��a��g�a�t�1D�0��	E��5XwO�:0�x8��,D�x�agI8MI��Q��r�@�a�*D���SƘ>���d����cO�����`Ť!PdP�ɨ��b�S�qܱSnRbiv���	"r��c�#\g�ּIf@ءq��%��D1M�l�wB:D�(�LO�@�LQ2�9<fx��;dL��5�:�D��-�8���k���"v�:�*Ɛ�y�B��c�,A��Z���`�S�7/*�@��K�Q���O?�I6b����J�'��y�fΌ�VކB�I�'%�C�u��i�LȎ"�n�;�&�����3͂��DX49��M���%w����Yqa|�FO�e�L�҃�ڝP�́��hϔEK�x��Ёm�}��'I"��f` ����f%�13�Ɍ�ON,����@�O��re(ɸ3��r&hÅ�<���'eP��h�9YІ}��*�5V�z@8�4�a#gkZp�S��Ms!*�D�0�s1�ۖ�Š�D�<����hҜY�IEm�Z��#�_�<Q&�R��8,;�G�wLlH�ua�X�<�"�	q}�C��zh� j��J�y��3��a�O,G�<D�݊�yrKI�-�ǡ�S�=�S�W��y��ī������:dP8<xt�A�y��@�q�HógQ�SҕD�ُ�y���`~|�z�M_��x���y��Or<�[㫕�\e��1�I�1�y�oC�~� l��b[�O>�a��O�y�dI�#�%˷,��:LDt� 1�yb�&c_���ρkˆX �B��y���>[>�j�aV����@�;�y�u�lř ��@e蒇�y��X<+� �
ɰ=��u"�珍�y
� Bs���P\�Zu/�=%J�2�"O��8��ԥN����+��t�� bA"O����	]�^���ղ7�2�i@"O(� Ѧ�=L��}�GT3��hPD"ORHI�̻`L>p�'ҶqO�cD"OZЊp阤t�N,��%�+��"O�(VfH%�a�p� (*�1"O|V
�9 p�S�dVa�v'�g�<yTȃ� �d�'(���3Bj�\�<�ѪF�����L�*>�`I�"j�Z�<�u���K8��⵨Z/cڪH�4`�i�<�Ϟ�|q����G>���a�<�f홣z�P����}�I]\�<�s�B��|�@����"����Fʘw�<q& ��R��@$*�M�����r�<��dy�T�sv�VQ�<h��Ӏ�y��	<3��+CA�~;4�[qÉ��yB�U�v��p�/Ev>�����y�ݣ&��SAx�V�d�C?�y��Φc�]�3Jؚp+���Ӥ�yr�A�t� ��fh�&��U+���yBeX�8m�\ @�2�� �VÅ�y�Y�s��Y��+�p�s�yD�� Tu��Q��lqD���y�ʂ�g�đ7�ǮH�V)�ul��y��iC�\B��16���e�+�yr
�4 �~A����#-�������"�y�@�6|-�D F*��>;�u����y�*�2J���a� ��[F�L�@kN�y��·;��( ���	R�<���'���y�iД�c/~y���t���y�KN�A 2����W7w��$��j<�y�j��Mh�aI�m�TX����yr�֎w3v��n��R,�ؑ�C�)`�v�ף�M�E�ŝ��84�E�4��sN4�1��|���'�X��	���)�'A6���@�"0ȃ�,A��$pJ% �B<Y��Dٛ$�l�H�~��=�A#��{"kT�y�9���a�4��Y�pɣ��� _ �7�O���L�/]F|��Q0y��J�O~��"�K`�S�O��)K�	��4���[Ca�p)��0ܴe�2E����ӫ!�, j_�-���d� �(��B��u���Ob���C@� �  ��΍�.��l#����'LVl��Ӏ�Xa�F�Z�`C��Q�3(Ո�,�@�)�i^Y�]�2�Z�)�R@zfeϷ}��Rԣ<��F��7M����.׷/�)�L�m?!��'�h��r�������`'L�Xd	Ω���𩀝Y]����]���� нT�� ��J0�l��jڂ1n���v'�?��I37�׿��b>1�&�Q1{�v�j�O��# �Y�"d-?qň�V���dq�+N&���`&����p(��d�O�`���ODiڰ�K=(b�U�1+d�!S�`�&��'�%[��ӎt6�EN�=�L�D ڽV��$��	T �=V�b?7���ӊg����!è`Q3���U�c�;��DA�S�'=)�@4��)��ޫINI��@8?���=���� ��E-��	P͇1�t��r:O��X�"�_�S�O�M;�qL���@�=��ԍ�4�O�R�xs�s>���l��׍�H`9 F*��I)7�<��S>��V��|�,AɎ�'����G�<�$E�;�/N�9n�����F_�Ot�r$�doii�g )f�@pa� ��f�H�J?qs6��9�PH�w�
e�Z���� D���1�'��|�)D�	�&���A D�@���'<P�Sq��q�@� 3b<D�dYC��43ۘ�POA,�b���:D�p��*L#�Υh*,Z�x�#ci8D�G�&2��=jw���}�LX�4B4D�� JtY�ٍ']�7O����E"O>��U�[�[On��,Y+g�谑"O�]���b�N:BK� 5O��C"O��ì ���D$N�1X�E�"Oʰ9�ź4TfP)5�6\�W��y��H/�r���E��d���"��yR���akWe�ȂA�܍1ؘa	�'����
�H($�ďr�9)�'������Wb���4o������;D��� ۳-���J�X{>qz0�8D�Ȱ�f	7k=DXyv"ܳx�u�v�6D��1��9	�x�$Iم7�b��?D�\�pHB:�|��5 �&H��e
9D����(ҕY���'�^=4�l�1�8D���Ы�
.v(��Ei۝q�V���6D����Wxl.��#G(qF* +'D�t�֊�5q옵Yu��g���.%D�h"'��q8X⣂D2Y��a%�?D���]ʲy;S XL:�a�M���!�$N=mz蕺#�F5''N<��B9!���$U��� �6-��c�F�x!�D��6��I�VfD��P!�WA�2�!�d@�`���O�8'S2S�@�$\!��%B��͂�.W9.Q�SGfJ(f[!�D�wY���B�G�l�F����ɞ/^!�'1�(�r�ӹ;� dK�CZ�
 !�d�26p��Ξ�~�����̃(v!���A��[�i.��,�
<�!��z��M��L;M�v8��" �!�D�-N����F�\�H����5#D!�DȜ"����C3NpIDG�X9!�K�p�
1"]5 3x5�&��]"!�D�.a���,�cXx4��`8!�d�3T��0��h��?����"�;�!򄆡x��b�+	-60�����ګ!�$@0i��S+��QK����c�)!��#fI���4)<�	x3(��!�$rL�����FTF�&�dy!��,iI.Ā֦L�f;2��K�(�!�$���,�)��J0*��6�б'�!��S]~hh@QS�:LU�(f!��U�Fp�1i�f�(�n�����,N!�X�N���B�A~N��*j!���,)���e!�&^cv4�w��S4!�$��7��|��	9^�<���ֿm�!�$�,fx�Hr΄�8M�U�Ţ��U�!�+ceD<�F��If��R�!�O��%`��1b��X���!�d�����S` �a �q"���A�!�Ę*y8�9S	�=����װ{�!�H/ZX��A�8�*�BA�W�Ur!�J�9)�X˓aHV�&�bbI�;d!�Q4|�1A��(�
�s���,�!�D-�`�
�C'ٖm
���"{!�O�nfLyZ0卥R�2�ↂ/+|!�T$ꚭ���\�W��l�6KF)I!��%x5Ѣ͚��](���: B!�$%԰bE�ED����&+!��B9�R�A�#�dR�S.m*!�$ߛI�Ѓq3 �z=���V�|j!򄞾q���F�W/|�6!��̓7X!�d�r_4��,���ǥ��VW!�'%�E�g�S�L�JZ�%�*r�!��J*c��CEAǿ"�����FC]�!�� ��Q��Ș?y��!$�V2jz(�2"Oh���#�92�%��L@�] ��(�"O|���*�/p�h����
z�𔩧"Ob�K��ю�=P��!{@��""O�Y�5�޺(�X���n6 !�"O�h��D"6��u	��C)��i�"O�������C:>��OT ����"O�9�S��Z��\1���6�r"O�X��F�?]�x)��mּ ˀ:�"OdM�`Ȋ7(��M��g[ ��I�"Ovi�P��3� �ɥ�O�Y�`$��"O2���A�;q;h�*e�B�4T\�d"O|�� G	�@$�dHH�>�X�"OVm#@���p�\��Wݣ3��ܙ�"Ofu��J�)Z��a�l��!��+�"OL� �1~Jer���	FҀ�t"OT����Wm�XєK�U@J���"O,� ��Tr�}�&��2n#ȣC"OBT02⇹#w�؄�͎5(�)�"O� 3.U>���B�Z.iFL26"ODԻD��7��+�)̓6��1s"O��sW�V�;�Y�W��'&�2r"O��ׄ�"����S�\��iA"O�����'Z*��%)���@i�g"O(�pH�.����'p��B"Otd�S&ׅ%!���$W �0Q�a"O�s�ʇ�Q�Yr�~ؚ�"O�5�2�C���N��uI�"O|�cnx~�ع"�3����"O^���@�S#��l�P)�"O2p�H@��\����NB�i)c"Oj�y�	Φb�f�3P��
k?���t"O���H���hpK�cgܡx����yR�#G��qg�J"H����_��y�N�E������x~4�B�+�yr�YF˞	��ևwZ��E��&�y2���:�N@8�@ʗE�eԎZ��y��(^6Q+1,H�o��8�c����y���V�ҹA��f)�a��*�y`��2�e���*]!��b��y�O&q�	��GA	gL`�3Z� B�	�ʝ 7�г?�ڌ5���Y�C�hĚ�2d����%�d&��l/�C�I3�d!Dm++�M�t��d��C�I�US�I��咪So�t��N��B ~C�I�FH#�G�\���GOU�:!�B�	<D!�l({�$�^�d�2B�&LfԍʁE�6/6<���/o.B�I�R��Ia���)��M��	N�B�P��T�WN�8���J`eD =�@C�	s�8�¶����䇟K�C�!I�$��]��BC��E��	�w`,D�H�De�#c|���͟]����>D�� M� Ψy 猬L{h"�K D�8�5�գ��uR1��qL�3g?D��� ��yv�#P/��VR�<D��JHL>�L�2TB�
����M;D�h�7�F� #p�xf+֮a���9�;D��bE
$HN,0�dQ$��\YQg:D�x� ?Sd0�`B�>ٮ��R
=D�X �q52ܰ�뙓[O�h�wm7D�0�e����G
ض=X�T��	+D��af��[�ʅ�D�H�ިYf*D��{¯Q:|a�pkE�L�� &)D�� H���Y�V�$[� ��50q�"Or��T�\(*��e���h�J���"O���`��]��Kt��?��{�"O���d�1VǪ�wLl����"O����[��F|���@����"O��8W,FMـ]�A 	>hb�	�"OH��CNO�;ܐ�.տ?{=��"O�d%���9�Nq�RC��xu�@"O��vkͶWY�9�!S�gЎ�s�"O| 4e@=L���R�O�	��Ū"O�L�夑"T.�EK��ߺ"�|4)�"O����'�3��Q2�	gꉊ$&7D��24�U�?B^,��	Ӱy�ȅ���4D�H�Ӡ
d8{e/FDe���ү2D�ԈH܆z8����hqKe-1D�t��ۧCJ2<�/ 1id@͋��/D�@�k���z=�ƈ	#`	^@{w�,D�l���2X�������e�W�,D��ǁ(¨�3E4U�ZA1'D�@��JL�s�:W6p�I#D�X�CW)T��h1�ĔPy��"D� �̊�@<�лQ��P����E$D�|���P?G8��Ti�.�a��<D��
���R�.���U�� �L:D�\����{����&�$G����7D��ёC0)a���q%H6���j:D�3t/R/?ty����6���D�$D�t�UCTjCŠ�/��%����1`=D�|Kg���>5:�{P"�	t>�Ya�;D�( ��!�`QH�	��:D��2��:vؐ�zQ�ǫ~Kxd��=D�lr�H��I��?0�Nܹ�>D�d��G�}�u�	:Xx��r�h7D�T�"fC5����vH˦d-�5�#)D�L�˥a�2�b�M�	��u��L(D����T�oN���ء�tESa
&D��PJ��^(-��? �=�%$D����X:�8����_��yz��7D����� �\�;�K'0Q�2�L+D����E�N�B�$��pw湃�'D����P�X��#��SK��Q�D"D�8��MI�1�Z���H1���Z�!D��ڧ"� ��Ɔ�o�J��!�,D�t��#Y�\��k�4Sb�/D�t���	`g¸�u�M�uH%I�'/D��0����l#nQc�# %@U�b@ D�PJ��܏}v�๕C���t9�?D��
�!��TV�ȫE�ǟ :P�e+(D�x��V�5Z�����w�h�'�'D���2�ԯ���pW� 5j�j�ۄ�3D��Y3�	\~QpÊA+'��8�2D�����+d���iު4���C/D����ʆ/3�j#ێ.�v�+��"D�,�BD�p��M��ℓ:�8!t@!D�8�pE��`��W�c�"ZR$+D�����Jѓc�,#�f�:�/W�yR��s>�8���"�,�_´�ȓ~~���V�j�@i�6�ɲ�D���d4�+��!5���H\�I�TP�ȓ&��)�Q���� �.)t��ȓLP��XD/�
A� ���ME'�t�ȓ0����1* .
Eʜ�b`��*� �ȓsF�e��ne�t]����x��ĄȓWT���  @�?�     }  �!  �+  �5  �@  �L  �X  �d  �o  j{  k�  9�  ��  ��  A�  �  �  ��  ��  9�  |�  ��  ,�  ��  ��  �  ^ �	 � 5 y �" %) h/ �5 < LB �H �O EV �\ �c Rj "q {z �� k� �� � �� �� 4� � ��  `� u�	����ZvIC�'ln\�0�Iz+��D�/j�2T����	#Ĵ��*�?YV����y�抋<+�����ݗ�z5���N�qd�Yq5N�2u�~H�f)BDgH�$ٷ��N�ysL��� ���&�E�3m�\�!�� f|	�`ǈ��tĨ0eݥ_��T�œ�[r 1W�������v@mڏ:E
���%Vz��4/��PjH�I�!ǿJ,^9���Ri�O�PӲi� 	���'p��'G��'LЕ0G
�8�i��>E{�J��'�Z���c�B�*P�O0��蟦q��"�����O�HQ�c
�9<�A+�<c�,�w����'�Od�$��;O���L�G��ɉ��G�|�ڣbտh�XZ���d�����W�<a�V���FGC�'��Tx��6B!6]H�Cߋ-�hS6֝j�I�<���Dn�����y�О^xP�AB�O8u)!j��?����?��?���?����)g�B�/ ;R݂%3�ĕ��02*�O��oZ��M���i��6M�O��o�� �aڴ&b*�
�L,@2�
4�Xz��j	�9�� ۅ���qӆmo���X���~��ޏ���K�(���(0,L1kbA�l[�i�Ă-�p�(3Ȕ$�2�~��Ul�?��'(��N�$�D�11N��v���pƣM�b� u�i��a3ѥ�
x���C�(9XcH��m�W=�v�cӀn�'��{0်~�lH�!�f� !Ѕ����sQ���M�ƼiP
6�˃`
�`�gQ"� 5;7 _|L�z� �	?K��9�C�J�0Îίҝp�Ĝ�+��nZ��Mc�i=N�2bgM� J5a���2s�~�"+]�Q���r�ʺiJ�y�b&�P�7�:dYP!qMֲHY����C:a����,�	5���j/�c��b��T=]�M��L���?���?���iF��0�l@�S�D��#��H�`����<q��?1��F8�A�EH6W��Ѽin�0�u�,���A�D:�"Pk�� ��ax2t�!$�j�VJ���'�Đ0��5���=uM��@��'#��a.O�@�'�N�˦�!��:�Ȉ�6h���?�����?i����O��k�X:�t�y���o�$�5��O���$Hg! �!���4���ɖRV�2���*+���z�f�?'����<Q�������'*��i	�@��w	�(t�ޥ<Er���O
�3t�]u��k ��Ц:a��vZT�zÇK�vjLX�"��H중�O�P#�K(�"DHҏ��g2����;���X�Hņմ3����f���мp!��H9G��OĬmڵ�H�6�$vx8j�a��Qk�"��O����O��d�<!��Ĥ�BQ�����^�BakU����hO����Ҧɓܴ�?i��i��)�:S<t�4�ΗKɀ�:q-�. C7-�Ov�H�����'�?����?	,OzA��$8��x�+� r�5[�cGN:�m	(�a/(8DjF��F���ϸ'�0��ޞE�2Y	f@�"wj�0 脯M(	X�)�R5Z :�����OT��K�T���6gO�9���e"[>3^�cC��ڦ��)O����'��$�?�O+�ɝ��QҲ�H�]�T�8�	��hO���$�>5������S*��0�� U���'B7���&���?m�'�D����I�:�� z�f�t�P�-N%+>�ꓶ?�����D�|��O0���B �
~�6$
 bK%r.���D�pa(��f�;2L�v��p<���*0U�E"�,^l�\k�+�	-p�\ZC��D�:�`�D��=�����'��<@B[�f�VE�bLL*&��d�s��[�D�I��M[��ITyҔ�Ȉ��V�j���"���9+��0Ri�Op��$;�I���u
Po��=�bf�*q���R���M�кi��Ӭ,��%�ش�?1�'��UC���:�@%��JW`6IR�����O^�di>=�G��%@R�1�æ� *V�<��cm��~��L��Ǚu�dL��		R�ra:dc^8�00Bԥ^�S�!�e� l=���S;��vaV�NQ �녥,x�� ��џ��۴�?!`��'k8��#?2�sc��;���4$h���}��b���U�L�$)2K��LA�
&�$��E{�Or6��(�2�p�ƋZ/"���fm:�n���xh�4%nF9���iㆸ� Q�`�O�A�5�6qRp��M��x!�iD�/�'��h�l��{���:�D�.���3�(JܧPZ�u��D�qm�00�aA��z�OD,��揮�lef�G�<�@0r� q��R �V�ccx�I�)M��uZ���=tTE3$�gO���z�����5#L|:��$LU�*8��$�	��D:C�Ӧ���?�J>����?�+O�%0�J�V2�
r��v$���K@�'^��$`�4���Ʀe�I�v�΅�G��1`�(7 �3��P`�4�?a,O�,8�����O��$�<C �?E_I���-�лBN�h�aR4�i!�R�%�M0�� U>!�3�	 %(8-�%��o%z�C�������1�`^�OAX Pe$I�O�^��i*��v�^X{1�f��!p�ĵ?O&|+����s-[o�ئh.O����'1�R�'a�F�U����H�#�=ȃi��oў$��S���~X�I
s���j�<���O��m��M3�x�V�'��d�O�哖\��(iVjN�ZH^1�'U�.Sv����M���?������)�;Q^N�p@�d�h��MC������I���!"���ש�bX�$`��"R�0k�Վ�a3*�;׉+O����R"j��Dv�"A�`t ���$V\!�
���¥bϤ�ȋ)<I����OR��:�	O�O~D��D��TÐ%q'���$�$�����'Yj�J��5y.[a�&�9�M>���i=�^��������Op�bb��#��K�P�D��L�����O�dt>��$��Y+ŀ����Y��)� ���C�R����l�EL�ۧ�'YH��٠R���إ)�6yx�A 6��:#�bN�Ę�V$��c��=�O����',�6-Fy�	F)HQ�4����a��H�QbR���<���@���X�ќb���ʂ�,���?q)ON�=�'?�����4��)�����`������!V7-�O�in=f]�hܴ�?1,Or��<9T�L�9^�U�KI�L]�Y0K͗�?��A�N���_2ՔX�jA=8xU��4A��w�֍�Ef���,My��6��	 
T���1.��[{8}p�.V##� آ�d�8�x�'a�f���z��hJ�Z.����h�Ѥ�O�Mnڎ�H���xp���H��K��D)���%1<p��$1?A���]���xG������RN�'?��h��o\�Ɉ1��887��z�2��MI5h�۴�?�-O�t�n�����O���<ypˉ"5���	��A2�cԠT����lp�`l��0=�2.�����)�ء��)�l���q��T�l��-�h����6��U�J$�)�+U ��w:O�����ڄ(������t4�@�2lk�D�'f�����̟�'��,p"8>ʱ����L���5�*�S�I
Z�ָ��`ϟZ�R��'�;��'7�Ȧ%���?i�'�6H@��E�~��e�T��(C��q	\�{X��?���D�|�O�0��K�����5m�*�v��!� U����R
�*i�1�qI(,O61�r
M�� �W YB}(X�!$�>p3��t�A�BiX� DAά6� *4�ƌt��̀���C�2|ka���1�̢P+��&�`�$���yJ��00 \S��Ϟml�A!r��O>6P�'��#=�'��'�B��%HZ�Cwm0�O�(=�9H>92�i�H6��<I���"���')R��0tA� �5�O=@����J\��'���	��'��'@�����9: ��O�x��HҁC�ޘbr ��sb����)O��s��Ј0�9��Qv6�D�5e.��i��gbzySr�t-ax"	�$�?Q�i� �Q����̈��M)���u��'�(���<g��8�d�2��q�}�eU�����4)�q �w�"�����.V��������D�
`�P�o���	k��E�:���	[����ΐ&1�R50���>7���'���sоi"�چ8$������|�˟T��W�܅C��X��LZh��� Js�|�r�Y��[=cK��#��<�'eH%��69f!�;NhV��'�mB��3�ɧ�|��s�R��PHq��<t�Z9ʆ"OX�3'HQ� D؀�����	�����<�tn���D5�&j�?hv|ё�i��'}�Y@�O��\"��U�In�����}�`"P�'��%J�����^� �x8Q䍀�A���"� ���1O aC��'k�Y�N�\) �Y��!(�"چ�|�/�!�?����y��F�
r2}�)ܜ5"~K��ɥ�y�>PR���֦�0,'���B��$�d�����|��=(T~`{"��Nb��ဎ�=����F�~V���Iӟ����D��� �I�S`�J?D����)�6�0� &C$**��"G��O��`#�'�X���Ɓ�8�L�CB_`R��b	���h����A�i��!�&8�MD} ��;�(����X����������?���x��'J��D˭5pX`���R5|0h��D�9q����O���'�O��VN��q�x{�-Îw�8Q�|�C`�,lnyb�Ԃ[%6��O����'u�����`����Cɒ�\h���O�zb-�O6�}>��4���.e��^�kHp����2������Y:~�.](T�� )؜F�ZP� Q��T$t�$���� �hU���p��$��mފ:�d�����/z��$�Oz�=3��r�DU>��᥍���q'���I]��<�G��h�&�P�aO�+�l��+:�O\��I`儭�c�\h��xX a�T~,��<�7��=y���'�rZ>�ENOǟ � �ԍ4P"�(��J4&�P�Q���؟\�	'p�brș!bVm�!"َ�?�Ob���r!�U�KwP��5Ĝ!>���c�60�U��1g�� '��h�`��aIRFJ��&
,|�$D�C���+ ��O�$�"|��iϮ�n��&� �i$T���d�X�<���8�B1��+��t\8�����|�'�}��� ��M�d���T���M�K>�T�����?������Θ8�ܨ��aH�B��%Vc�h�f-S�(�<�F��M#�,B����|�<i�H�8.neyZ2/[��9��]�E��9� d�D	�� 	k5����yb�M�"�Yi��^	����$C.�?	�OVI;v�'��'��O���-	�6���@�#�,ৣ;D�D �B�9fJm�S�K�4�,��tL�<�B�i>}��sy�":o�tzu�׏<f��r�@�S�41�s�Uv��'���'k��]ߟ����|�6�N�!�ǒ!Z�����V�8A��,���d��<�VGX�?  ���MH�M�Hxcs�3@�b� �t��T� ������!�l��e�ԆkxQ���	=mzڰ:G�'�j��j�񠂙�6ٔ���<�!�d�I�����dN�@X$��
P;@��'��7-5��%zIo���ɱ9�.hR��2j��#'	�Yh�����b)�ӟ$���l�h�(.���� ��or(	�Pώ&G�$ zr$*DD`{�,��o��Ն�I?^��YA߱U������;^sq���8!X��$��R��qį0Oʽ�'U�6M][yB� F���P�CB�%JN`������0>	q��&q�$}��!�I�$h埐逤-�S�Ok~6m�4�@��!-$:	���c��3P4�D�<ԯ�	s�f�'�Y>]З�j���Ԁ8Cq�-Y� �:�) �Xޟ ��5`���PFA�1� Yp7��tZ�8����Z����jE�+��U���
��N�'�9���ՎdM~M"l�1*��}����ܾ@j�" e� ǆ��]g��)�OZd��'�6�^}�O��)Ĩ<:r� Ǐ85��!;�JQ�p�"�)�'V����Ƕ��iy��G�|9��M`�i�1O�)��鎨U�  ����P�H5m� ���Oh�d�!���8+�O��d�O���zޙ�7$Ơ~��=� �V7.4R�)�h
�����W��M�"l˜FF~9�|�<٣I/_�VXK�����*�x�˘��a�6�˯w����^�.O�����y�����Q����'�>�ѓ�. ;�'�6����јϘ'D y�l�".꾀H1�ӂ4� �(�'�ܑ�%E��h��0iݚ2ij����?!7�i>I$�L��	{�-���U�}���r��^2q���TOz�X�I��d�	��uw�'[��'�F}ڃ�P�viX���䕯i�RC���0��d@�+�m�o̦����b�Q�ĪEHL�p%*�A�)B�@woɓx��\;��_*r]�D�a�G�p����I3Q�؂4����s4�S�5w� ����#O�\�D��Iъ�)�I8YHU����
�\A�e*�g�ֈ�'ў��*�i18�N��{I���WA�7�bDP6�'��6m�Ohn���MS+��iXTHঽ�I���[ oYK0024jF�E'������4�	"3-ld��ɟ�ϧbS�S�v%��,2�~�v�Õ$����'�f����@Ȝ
^��� !) ʓ9���b!U�YC�Θ�i�I��ۯOo�8����,�RQ�@�r�tE÷!-ʓҘ��ԟ��'�)�#@�+6T4[#H�3�ޔ�H>����0=�a�7�(i(��r�9゚���hO�)��4��Q�$�dJ���Tj�!�O:�ɬE;C�i�r�'q�ә:�>��I��<p��Ꚋ]�j��"gZ,B��	��@���1�}w�J/�|���mԖ��	6��cHRym�sN$t�|*�	[Y~"����4�7$#i��-f�����n� r6X3��(C�i!I���۔Q���'��>����B��T���>�r�!wO�{V���ȓc ���6��X뮬B ����<D"�$�'Y
�M��'C谘2Ra�+V2z���4�?!��?!�1RR�����?1��?�w��]����ĭ�7N�LBz0xf	�l̈́��ҧJ��y��"
ИO��'�h�3cJJ$��F�E�`0y���4Fz4�R\�]�<H(����O��'Q� �#a��&��h&�F�Un���������`2��'l��$	�+� TRx���/�I��C�>{��x���ޓm7��j@�(c^˓����П�'6PJ4�T5BL���@-yPP`j���_yNm	d�'2r�'�R�t�)��ϟ���'K���t%M�޼Q�n�tڀu� a�e<y6bџBHЊ��K4�ؽ뤦�#8F�����=��p@�Q'~��p"G�ua�<y7� ��i�CǏ�J�9����:bւM�IşĢL<����?aM>��O�lc���A�$���gK~���'�鈖��Tj���AR�43~x����?Y��K8���'F��5p�F%��4�?��'6����'��_~��4^��Lp�$lGx�E3c�q�&��2��ҧ��0<!�n�'Ҝi���Ž9chE3���
Ól*����#��2��A��HO�J����A�=0��<vH�V�Dc���6
ɇT�:������?yƥS�EI��ĕ���}҆�s�I<e�޴�䓅���OH�6�L'f2iԎ{%,�O�$�v��P��Q����5L	#|���H�B�EC��3���W�t~���S� �c���S_.��B��x�O�\�(�m��f9<�"u$�oѓ�O|t��?!���z�XC�"\WG�l�B�s�7D��Y�G6�٩g�70�:�O#��c��>M*լ�G%��3#C��x40P�C��1��`y��Μ5����'���'X�	�j��ٳ��ʣ��h����.��ĚU(� E�Scn��`v���Q��w�g�#hL�i�� 3
\�v�wG�x ���P��<K҅�@xv��bK\�g�S�? ��q��M:r-�:�ؔS3���'�'���0�~B�'zў������Ҵ��bHg"zJq �u�<q�i ��D��I=+��Q��Gy��)��|�����s �q�l.I�� ٣���qkBe���O��d�O:��<�|�(R���B%��1�P#a�=�T��tL�2B�)�4G\Յ�ɥz����X 2�I���|��,[#�R�'!R�#ҫ9�����'R��pDg�f:�{6E���,�cUN9�?����hO�#<�nΚ�V�#�6$, unKc�<ABT�
���R=KYVM"�^򉂴�$�<��K�8h���?i;���!"��骅&!r���Bp!-O����ɷZ�$�&�O��1y��G�0.��d+��$`���H�dlDm�/7�����K3OU�e�'�~�O2	@�N�qHp@!g'S,iL����"O��P�~��,bFH.��0���'�4�Dd� ԑ�ޙ=x<=���37:�'��('# �I^�t�'���B�B=:�M�4(2I<��4�'�r��y��f
y���F�N&�>��$�	�U��(F� �N�pl���;?��j���a�&�/ϔ��u�1�'SO�<�(�(�h�se��l����'|ъ�P��3�'�"�k	�?��U ��W�D������y�6%f�RE(T�d�qG!� ��OjeF��"�G.|����+�B���iìv2�Iwy��P���'�r�'1�#c������U���"&�� �L5�-�W)Zq6-�,J}�pϐx��2�1O�]���Z�>����$�����Kӝ\�v��3j�RK���R�2A�1�1O�Y��R����ԝt��XÀ�'i��(:���D�O��=ق�2F�V``#+�G�d��!�D&�y��6	�q{��E�)Ϡ�b�)ȧ��I�����<Yf�˟?[-A��k	�$(5�Ұ�0����?����?q/O����tǋ�KY@��H����zv@&0����FT7lp��2Uk����k�#DC�0圁jaf%b�
p�ϖ*R[H�BT�L�ǓX�H��Ή1s���w�Z�`^Ƥ�SI՟���t�'����@E�L��i����^OP!���;D���Q�fG6T����"�8����$�k}S���MD���'8P�b���?��%�ݠPe�4�	jy"�'���'�x��cL)�	5� �*�x����D�d�N�+[^�
��&	ax���~ܡ�l�1 l��`E����I���2��96d�
�o���	ݟx�'����CE�6���4�Z��O>�
�	<�	{����X�]�� �����	�?���O&}.&8P�+�.qS����� �'�8�\������O0eY��3Jl�C*�,�41e��O����"��m�1h�
CK^�P�,S�{j�?�S�����JPz爃|�~�h�,n~�+���}r�"�ld���G�[P�Oz� F��P3�ar��D�Id��Oh\Ô�'B��<)%��$G��5�eI��+�@y��k�<�1R�>�PqQ�#Xl P(��o�'��}
�dfRA��>e|ph�cy�Y����������	�l��my5�"8�ņ.j��������8���;ZrP�5nJug ɐpY>��g�"�tQ�D�\k0���0�	��	"��hG�ǵ.���B��XK�g�H���Cso� ��" ǜ'�����s~2 ���?��hO����e&��u�U0{�ice<D�`P�倰X�����7E�-�4O�<A��)z/O
��6��A�ȱ��/i�~��Ѯz%H���O����O��S���'�@l��l�l�X5�Ħ�;`����K�d�8Y�GIY;iV<�L���p<a��Q?=�>����ǸLJ�ڒ,�,
P���2/��
Ң6�*��D��_�D:�l��f�$Q:��U&W��<k��'���Ir�'�Q)�Q�I�*<#����@�|s�'^\�u�47P,݂�b]-�p�!H>yv]�t�'{�ĩ5�:�	ޡGZ�  �H�\��!C�
���T���Iğ��ɖK�,[�)S�R���ё'E�J��m!PjF�S��bUR2:�B�{��q�ܻw�۰=�LI��nP�@\�Iv���hтe��S�A�|�hD�0;Jp����@���'F�	�~~�@�gO˚)�� �IK� ��O����.Xr�BpO�Ϭh��AX5d��.�O�Y��O��`"J'r� ��'y�2jj4���i�|b��0-�I��DyA��#'�\����?qg���p���
��QNC������OiLթt:�� P#��eLP+C�� 8�a��� ���2
�\����9a�@<d�pR��;\���{�(�Iǟ$G��?O� 
ET�#Τ��H	>��� "Od�03���.�q�HLF9%�	�h��DA�ȟ
�`��G߶A׬]c�ed���6Ϻ<��/����IVP��E�G�&�@ �ȍ$��a4��fA�`ʡOAD�pxYB�2�3�I0>�"�YP,ٶ&#�4:"NN/V7��r��?�v�ʡ��P�va<�3�8D,2��%}��)�K::g�$l!�򤍹]��O �3��U���r��Òe(��jq+��^2C�I�z�0�Y��ޮ5C�@�ɟ�j5�ʓD�����$B"�8�4�~G�L��E-�4�ehB񦩛7 7\O\{�f�'Z$۶H�#�R!��m����!fI�O�	/�p<� h�[�l����*�N�8�u��f=mX�Q��������5���u��^c�rת���T5!��w�z�Fz�������W;����j�>�B�	/��W��EJxE�� M#}ҒO���'<�\��0aٴKr
��'"Or��`��H����0�:F{8O����ӂ�����\�j�j����W"CS���5	���ᳬD-���D�^{�r5�1O�x1��'ڒO(�s�1z�,��M0[d��U"O��0��O	�^��@
;?��=j#�'�d�d_�)�-�˘�a�M�%ə3%�'w. 
��qӴ�����+HH
0���������9D�j,�HP�" S ��1���}u��|��B5V���πi��cED~BE�#���[e�:\�y2@C�Op���2��sb�ѿoKƍ{�OjTѧ�'W�6��X�O�	C�Ԅ+�Ȇg>q�&�L�!�d >�4{��	qb��&X�Dbџ�(��)p.���g�Q�0:P0u��R�7-�	˓Э
(�Q���IS��u�0Aެ)?��
d"+�	=Sl���VKvB��I <f�QP��ZL1O�Y0�'���7E��/}|��'"�:b��@�d�|R��:�?����y�9e����H�~TB���IR8�y№�*�Ö��q~4|%������m�����8�g�<>���#Ǐ�h���3Ay� l�K��0�A�ѴWr@�@�GP2t�H���1�u�-u��O�p��@
#lVT���,Y�Iǟ���ߟt �E� rdɡ�c�"t�i>%H��T�<^�E��s�<��7�,F~4p��_��ѕ�tc
�J�񥉀'y��p8�n�ЈO`@�G�'��)��%2��S�F�F�nD��'P�>���[���yg�[1.������[��t�&&�O"��'6���퇕��v.�9)��!�*O�|8F��OX�p�<�)���)�Ox��ENZS���$%K*����O�I�ʌ~��Sc�^@8�@�t�Ou�(7K߽@zҐz@#]7rL�!k�'�*BW� !0R�A*$�22."��ʬ|��!���?dr�9���<�'�ҟ0�	~J~B�O��B���Tr���/ǝ9�zY9@"O(���jI[��KMZ�ɅM(�hOF�E��"�w��Q)*�������a6�' B�0o �����O~R�'0B�|ݹ����l)�� U3!~q���<lҲiثNm���bY�\}�%o����ɲvf��O�	'�%$�T�Yge �������K�r�な��O^d5����4���>�~ps��>I �I�e@�]9�rrj���h~dƙ�?����hO�牲3��hA-C�`d@�&Y�?�:C�IeN`��%D��H7���Ⴠ&=������HO�i�O��#y�$;���;+��9���@Ba��CK��Gm "�?���?�����$�Ox�S�c����̓�n�x�FA�&~Pd�"��9����� I���� I]�'�,Q -�}��
R���;|�H���(b��92681�)�џ����Ỏ	��
* ����ƅ�~��,�!/�O�D>��g�O�Hq�I��� �
� �< �p��F"OH�[rLX�Lj���`��jyd��r_��Sڴ�?!)O�|zTn�Ҧţ�IEԟ��'Ұ�H����0%�+�<d���Ɋ@4L�	��H�ɻ5�T)�BG=ј�y�-��Sp8�"-חJ�p���B�����CԠQ��`S�$ʓF��xK�q�T}CE�4f�^�P�{q@�X1�ɞt���a�S#S|�%�T 9�K�����$�|�"�J0C�R��5�ܠwN(r2��Wy2�'�a|b	�M f�S"a݋E��4:D�P���hO�	�Fy���Y׮� u��>$,���U����	(�lڡ8Qd������� Gu��'��@S�eV�z̙��G0et�a��'I��:tF�2*ȑH�K<t�n�|ڋ�lߝI��ڄѢ*�5
s ��y��M1z$ȭ�!��b<��bJ0�'Jrt+����Y��X���+:�b��A�������(���?ᛧ� �`�HN9%?Ҍ{r!R��vT�0"O6���ƀ0vrvtf� u��u���d�O�Ez�Ok@����;`��Q���N�44���fH剗m�,l�ڴ�J���?y*O���(P=��,B?j� =⦊T��~<�g���� �f�S�n�]ːK)j��^:p��'Kb���<�0�(��CS�0$�q��Ip ɇ�I�j`��aE�K8 �O��QaeCNQ��T�e�t8���yԜ�p�Iѿ/�H˓\���I0�M�Ο�'��ĕ2	.�<Ð�Lp}�P���8S!��ÔC> �x�Q.o�-؁�J1[�-��|������3�\�f��<=0A2�f��.$ Yyd�Oh�3$,�O��$�<!�S�� �:T1Y�lO�j�B$����2�p�Sg`�u�:����	* Z�	Ǔ	<%��4���@'��.���F�ξf�U����CC�L��2O���&�'y�1��	2&� �d���eܰ����'ўD|���+W��E��ܜC�!���yҋ��!<��-�1sa��{qB�?���Dɦ���My�b[<!H6-�O<�$b>m�6�4R��AӰ�ؾ6���(�O�AS1m�O����OPa�5;O�OR��h�1��r�j�JU�Ǆ ]�#>�sEØ�^�iB�6b��9�s&Ů$B������]@��Ka�r+ΐXׁ	�;���<�C�矠�I���'c�F	;��#�,`�K^��@�H���?�J>i��霬"z,9�
�n��5��B��DI���� ��!�I�WBd����7N�ڍ��L�;n)���	Myr�'�2�'&r]>��'4��Ť�1
��ʑ�`�>�B�O�#=!�4�O$�	$� �J�"�봅F�+���C��s�O0u�J|"%���56�6̛�QG�a�R�����'̆}�q:O�(�'o��O�R5Or�V�C�֩C$�ͭ
<5�v�R%:��6��Of��Uh�O��#	��s���	P�\c�N)�JU�id��B�E�J�~�a�������*�����u��'Y��O2b6Oށ�%EA${��8��e��$:AbCA�Y�b�'|ƌ�R�'@���z|���ugiJ�<Y0MuY̼{�C�%/���b�l��?q��L͟���.&�.�Q����d�O6���O"�ہXb���-	um�s$��h`V�Ox��U9�,��x���ͬ?7��d����X�"B�y���"��
{�V`oZ�<ٔ�Ɵ�		l1���?	���rc%�A���j��J�)R�P���	��43�'7�$b���?�ѻ��$a�(�c�?7�P�h5 p���N�����%��n�j�F�ǦeΓw��{�4J��@�������b�)���811�n�Y�����>^��o�$'<ΓC}�5�	ڟ�����ϓz��1�'&�@Ő��9{��0�d��^C�4� )Z����?en9�,O�㚭��+��M.(�8�Qa�H�`C�	7J�LXE.C-
��q��\7��O>�D�O��$�OF���O|�d�O��D�n�"Mq��91of�Aq
�/V�nZ�X��şt��Ɵ<�	ҟ���������)?Z�c�S�g,,�Sb�W=X�|޴�?Q���?����?��?Q��?���Ib�0	s��@#b�q�O�LT]Q��iUR�' �'KT��Oj����9�ޑ��ω�R������l���֟�I���G��P-8$� �� �pK�iv��j�7-�O����d�O\�O&�D��6@��dhĶ{�#�m<l��mZ蟄���(&�D�O��i�Ųr'�&T"�f��S��AI'D� �6�|�n�t�ۈR�%K:D��
��<|�x5�rGιk�#D���G�	A0�D	�?)����%D��O�%�D�-�'D�Ã�#D��Qw�\!��j!^�7�.`h�B"��?)��?����?�t��*`�q���IF\Q�`�=g��'RR�'���'���'R��'�R�Ê]q�❾|��\y�[�h��7��O����O�d�O$�$�Or���O����LY<trt5G�Ƽz ��5cnXo���x�I�\�I��p��ş��Iҟ����NF�5a Y�Mx�aXH��h�J�ݴ�?	��?1��?Y���?9���?��� l@`���1��8
W�4i� �Ò�ip�'���'8��'"��'�R�'#L�E�ĄattH�dO
TmVѓ�es�>�D�O��d�O���Of�D�O4���O����A$)��-ݙ��!@��ߦ1��ӟ���韜�	֟$��� ���ȋ��9��`w'�&!���-��M����?����?����?9��?����?A�ᐌ,�,���a�%��(��F�'b�'wb�'	��'9��'�BڷA�����5
tXA��9k��7��O
���O��$�O����O���O��$����jP�S�\�CdO�4��nZ���	ҟ���ן���֟$�Iٟh�I(W�Pxa���T[��0j��݆�xش�?����?9���?A��?���?Q��,�p	s �:y� �D��0�^p�Ѷi��IٟH�'?��C␳?�i��F�Jw¹*���Ц�r�;�	�?&?�bߴ�y��ױ�2�[� ʔ��]rV��R�i��$�<%?!Ed�=R���ID�DÐ��$��A�-*,� c��O�DC�EI%}V�A��2��|�'�T��N�02x	ƪ�?谍"���8�$�q`D+��u�? @ę6FX��eҠ"�
��g�'@�'ێ˓�?Y�4�yR\���g�B�N�Rx��e�0xܚi'	�<���������g~�OQ��)u�H;NQ��~3|d:DnA!�&��ңQ�#C�Iyy��'B�>��(u�N���"NNu#��F��$Q֦}A�E)?Y�i��|�O��L�lV�V�@U�Æ�J"\�`�0Od�$t���d�dH�v���a@N�,r5���
�S*��:�%�ԃA'�F9�g��ş��'<1�NЀ�-����BЖC�≣�P�,�4��<)����L���`�@��d5�!:��S�TW�0`^���I�����H���j�֔i��C&`оrO2|xf� �*Yqp�����= E���P�My��'[���T�
!)F��h$�L�U�B�'!�'FR�'��ɟ�M�DƜ��?�u�O/���S�h��~�l�b�?���i��O.`�'��6-�Ȧ��R��&cH+��%!�]�x�F�;T��k2��	��L��cU����`HZy"�O{�Y!9\4Hs m¨E�8�zԤ�6h]��'���'RR�'B���C)�����/qP�dL��Vv~���O������b�nyb�|���'?q`�N]hh��Bi�h�1j�����&eӎ��D�5˜`��:OP���+�<�!Mw$Ē�G�L$CdϷIK�4@E)�į<I���?���?I�d�вġ�%j����$��?q����A٦��HL���������O�#F�P%�xʅ-Z4?<i�(O��'�6M���13L<ͧ��+���zT ���j�^�S&#$��mAWU�SͲy�'\��.����F�|ZI�ڼ�#���i�ͦ;�@��'���'+B�'N�Ok�I��M[0�޴\�:�(/	Ej�Ӄ�;cy����?	Ƶi~�Oy�'��6��jMX��scP�l*F)�WH�7���nZ�� ��M�E�������*���r4��Ny��� u����_o����e&{�\���	ޟp������	ҟ��O���`��ۊq�"{S F_��R��i`��(�'l2�'��Om�cӊ�	6H,�(��چ ���N��%��|o��M�x��O�$�O�Ȉ����yB��;&�̰3@QR�\��% ��A�?k���g%�*`@�'m�i>I��?~EP�J�^�X�f��!����	ퟠ�����'�7S,F�^˓�?�uOߺ\`���#&Q�v�3�dہ��'��^�&eg�@�O>|JpN�^�,�q�f����1��O^��Ed�9���Zʓ�J7�94*D�"�'t��C�PE�b��ƆЭ,�D����?���?Q���h���ɲ�*�$�E	g�A����gyF����u�PFM����I��M�M>)�����e���ퟅy=�ܸ�f�>�?Qu�i��7��O�����s>�d�O�����ÙD�<��C�V�D�%�2E�Iá���O���?���?����?)�&#\��F�,s�@�5!$3by�*OFxm�	�:��	՟8��B�՟�w  �kt���JR�R��dɕ�B����Ǧ5#ݴ���|j�'�?9 �dN�W@�VYli��
��aÿ�򄁊i$��%G����O�ʓp����N��p�����r�\�c���?	��?���?I/O��o�]���̓W��ez���$0K~Ѓ��E-O������MیB�>�#�i587�f��`�ӼQ;�����d��Q��^h��U3O����|�z<p0eӽO;<����w�괙c��S2,�!�(�Z��$��?����?���?9���!��
]��z�$�2��hS�X�	�M��@��?I���6�ς*ض�*ħ�l*����d�
�O�|oZ��M���Ps�m�F@��<i�xvqY%�!�8]�so¿�0�P�J�B(�1Z'Wl�OFʓ�O����P)�)9FDJ�M�|0A���Ħ�H�`F����	ҟP�OFN��5���>b!H߶S�T͛(O���'G:7mѦՒK<ͧ�:w�V>4�FQ*pd��\,d,� ޛu���'K��]B�/O��).n�~��7��.n̖����d�9����:}����������&g��99"�ڱ���"E�8��}�	ӟ0۴��'�B�jr���'`��$-��0��5�L�v�7��O*��ヺ���O*��iWN4@���<!@��)�p�˶_˜)I��U��?�*O|���O��$�O��D�Ob�]l�<�l�p͕�twD�ܴ!z9!��?Y����'�?���i��DR�M����OM��Bf��R� 7��֦}$�����?	�IF �R�bu�4 I�5��+��-El�@&�����[���f����X�	`y�����7J��E!A�<�H��!� �?�VI��b�'	��j��i`O�$Ot}2rϗ�`��Ob��'Ԋ7�ئI�M<��d��.Ӿ�C��"P]K���?���Q�sN�J4:Ȫ+Od�)A;R�"�x!�g���s��`���"`�,{�H|�C�O����OZ��OĢ}��'�6YS���=O�i{�n��z䪉B������ɜo���'�7� ���OH����q��	e�U%�� bf�L:J�$ߦ��4Y4��{vE��'���7}�Xz�׈8�T-��H�;-������A��	�|�W��	��	۟��ԟt��c��ь��Ǐ��3R-�qy��zӆ �Dh�O����O������O!'.��0���fg"q�Q���9~�'7-JǦ��J<�'���'e�����fS�V���y�E�M�|�$j߹[oR�*/Ou3��z�f��4�5�Ľ<iE��?����ӔJ�P�Q4F�?����?1��?�����$Uউ�s�Eޟ�� �<@$�$Q���)HŒoj�h��'{�66�D�O�d�' P6M��ϓ�z�*��Ԙ>q�XPUM(u+>����Kr/V�Iџ@R��R��м
7��Jy�O��N��U��ɳ7 �4xbv�%дZR��'R�'DR�'�Bᓌi�R,�7��-��Ae써gTP�D�O��$\Ц}e$
럈�ɺ�MO>Ia�S�e����w�S*q��a"��{7�'�d7-�����%/@�u0��t���	9�Z��C� �4�� )[{̈3�L<T6@ca�|yR�'�B�'��D�F�,����	c�<,+�l�C�b�'��	8�M�d"�?����?qΟ������`j0��+�Va�V_����O��nZ��?iL<�'�����e�$��Q�]s"�����O����s�цXU�=�/O����^NjEa�H7�A�U�<Z�CT��DEа�ܨ�����On���OJ��+��<�C�i6ni�ue���5��IH����X��V]SR�'� 6m1�	%��ğ�͠�	�4H>ybW�)�h�������M�T�"+����<���;i�]�G��4PR��)O�� w'�Q^��Q�#9Ҩ�	�Of˓�?���?y���?�����IQ"6��;*�9�J�c�ŝ��N7�Z�}h�D�O��d:�9O8�n��<2�Ú|~���C@
�t�A�=�M[��i��'����O��1Ҽ��'kx|����28�ȩ�OL�fX�H���'���ic�@��\j��|T����<�s��3\�xyyd��;)���)F/�ڟh�Iǟ���LyR�r�
9����On���O�q�r�挤{�m�z��y��hY���'���7P�� {��O�I�ch �0Цy[t K*R�QPn�O4�D��ΈVQK�Vʓ�j�FFT��'҂�ʅ��9M��a�g,APDu���?���?��h���	�l��`���J�/�q��<1i���Hͦ����@��<�I.�M#���OD��W�R�i�6�Z'kZ2�va��'�47�@�u��4Bm�W�<���SЊ���
U%Ќ���S�-'.�sXn�x
׮�C�B�O���?I��?����?�����h�;R&��V�K&��dsr�<ᥴil2%U�'b�'��O�劓0�&,"AGT�$Az�# �D*�z���w���O��Mq�xS�l�$���D�
WA��6�˓A�"}a�D5}�TN>y+O��H����>��2�'[�$#x�����O��d�O��D�O���<I��'*.i)��+z) �� ���{�h5)��lb��t~���O}��p�d9�	ʟ(Q�?&�������&6JpR2�� [��c�?O8�d'}��iѡ!>�<��:�w�������@�	 �������?����?���?�����'t�}�`�?s�ja@F���4J�����?)���?���iQ��x��'��`�0�O�j��ζ/�"���f�U�.%�'��a�ɨ�M�C�i^��LT&�E��<���0��P+���0*��+�/�P�� �S���7�x\��(	=�䓴��Oh�$�O���9h����u�
%��hA�<�\�$�O(ʓ8a���ܩ_����H�O��XcF�C$@]L�c愊%�li�(O�}�'+�7�9'����?�+6*��?�X&�)\��R�¨b'�+��O+g�'����F(ДI�ʟ�d�"A<xʠ��'4TXl)7"�"z�!�dC,�(��2�l9`�Sc�C:$����%�$Y��� M/qd4����Rt]��f�lP��[c�B.8��{�N�(\^����?" BbY�M�l=Sc�@hX��OP~%�I�6?$�m�v,D�*:��a�S+`�v���ƫt�*d�ca�����F�Կ*��[�IO�d@��B�_�R̸R��ʰ��L��I
��p��;�
���
��?���s�
��Q�ηJu����?q��?ͧ�MS�(.����Ce�l>@�� �q"=	�� /��3;�&M���0ga��jE�2�ʘ}$�����0mh�	��N�B\@d��I��A��G��G#Є��� Rz$�:�o�F@�Q �Y6�L@���$v|���3N@��N
9/D�Ä�O�}����V��S��>Z$��ڐ��'p:y8$F	d���@\��;1�I5Rh!0"DF�f�KI�r%�h1�X-�H�b�G�}�`T�㛁 o��1Ɇ5B�� H�L |�s#<Wq)����<�,!iGE� iLz��G�DŲhi�O�xH�Y2�%*{P�����(�5s!��k���6U�xq�( ��D�b���n�����.{�1q��'���'+r�O�����
ƚU�#fD�	 �V�[��؟��	�:�0�?ͧ&r\Ee�l�|�i�DR�52P���r۴�?�7��!�?����?�����*O��F�)O�ͲЀ��]�Ƽ駊	֟����ؓ�eE[�Ş^U�͈2e��(�q�X
.<ԬY��?�T��?���?������OT�DN0p�xtK��_�Y�̀,	{���D�em��b>)�I���1��\GX]c�j�2
��h��Q�������8�I�� ٗ'���'0b=Op�p��Z^���I�ĝ�F�ź`�'��''蔂�[>��Iߟ�I�t���U).v����n��]�!��Ꟁ�I�p�'�B�',|R�4\G�
u�Yu͔Mx G�&���d�2!'����۟�I|y���T�N�*�'+c�&�¥��uh��8_����㟤�	t��㟠��?�4Ejg-� �N��0�;?�ak��e�	ӟ��I��'p�LS�=����qnQ'>���bB�\|p1��'�"�'e|2�'d�ܗ/��$ˈs��A�l��5tD��������,�	�l�'�"��`S>}�	�?y��R��x�6�3�ş�bA����H%�D������g�EI�1��h[�f�5k�lL`�
&ҬD����\��Dy��(��ş��I�?�;�)�[�d1A3��=���qɐ|������ Y`���?�'ouf ��aҝv_����Z����IBy2m��l�2�'"�'_�^� � ���f����0Տ:I�#�'7��'�ق��IQϊXh��]�=3x��L��?�2Q���'���'�D^�$����3'd�mUJ�%Y%bT�R����(arIe�S�O�bc��؉℥@�)��X���f���'\��'�HVY�d�����I�<Ir�����=St�ʅ `v�u�h�w};M>���?���Q�Y�ɝ( �+��+t�B91��?��!��:���D�'�^�(._�Sc����J���K"j������8.��uy��'x��'��I�F�(��*��*�����˱0f��� ����?I��?�/O���O$Dq��� q�I�`	��B�J�;���@�OZ�O����OX�X�:q�Oڨ�Z�
r���YSmM8x���Y-O��D�O��D�<1���yB,՞�?J�1f�A��IE}�9[�e<��D�O*�$�O:�J������,�(�|����5��DS���@�B�'k2Z� �I񟈀e����O٘���@���恁5mh93���?����9S�i$>��	��K�gC�B�jö��!W4���Zʟ`�'�r�'wΕjs�'��O+��P`���dL� }}���'ȯF0V�lʡ��/�M�(����矬�'&IR��ܥ� �I��Ü�\q������:E&��:�I-�I��1��M0� <4v���IMz���f�F�o�ٟ$�	�������|6/]�:'bi�����1�q��?��B�?����?I���b-�b�'>ИAd"��b
�p���$pr���ҟ��'�6��a^��'����#k���kMju��ɧM�3�5��y¯Z�*��`��x�0�צ�/�<��$t���Oj���p���,�	N���V�
�
��a�@��6r��	�'�Tq�t����'��\��	�;�~D#��'������϶J��b�'dy�'�R�d�O��D�`�	�Q�'��?��M���/n1O���<a��n5,]��Op��`��U���V@]�O��L���?i���'�2�'�d}���QJ��yU��V+�A�I9X��Õk�I֟��'�"\d��ģ���7y�h���{�X�١O��|�?��?q�ƌ�C	BL�O���VZ=��ԑ�%�,,j,�6�'"�'X�)9V���N|J��y��^��Xb4�3Mdt���J��?�-O6�$�Of��)�ON��V�]/X^2�b�òU�"���ݳT����<��Ċ?$̛�^>y�	�?�z.O4)X� ̢S&!S�'�,%�tZ�'"�'_�����'�ԟ��a����҄�A�I<a5|�<��?W�m�"�iq��'C��O�"O�Iq�,`�0�Įs����eb(?J���=�d�O����O(���|�'8L%�7!;��ڇF϶EvD-�%�tӬ���O��DZ�0�4�&����`���R.>G�F<[`̉�+��)�ć�OT�D�O���7&d��|b��?��@H�Bi��O�t��A��������?ّ,j牧���'��'P�'��x"\���O�96�u��[�x� ����l�' ��'��Q�{�o�9��ř�D*M��X ��	=X�8xH<����?a���d�Oh�Tc�v���ɹ6�(qQ���mp�8`��OƒO����O�ʓKb@�2�O���w���^ Y�j�r�H�8-O*�D�O��Ĵ<����?���ל�?�6�мOs>EѤɝ?����!����d�O��d�O˓brN幤���I <Mzϔ4:�4=p�ڑ���'�R\�d�	ߟ<B�������O�^}J�(W�x�|m	fX 64M����?1��򄚳"�B,&>�	ܼ�ň��L�ڧ�ҪRK6T:'�ByB�'��ɻ8�p��g���|����-'@��iƦwx����F��ؖ'~�IjR�Ӹ�'�?���v��	;y��l���R�"��!�d�%h����<�cFӇ�?iO~BL~j�.u٫�`� mf�����Ui*X��	n�z���4�?Q��?Q���
��?���eo���ɕC#��k���@�~�	�Plp`8���?,O��0�i�O 	��G,t���E��p�*��1�Ѧ�I۟$�I ֚p���`������	ӟ@�
�� 
��ڔ�r�FEGџ��I`y@32E�Oj��'}�b��L���GޝC������.B�'�vlJ4�h����O����O��O�������&�8b|�Ȱχ6(
��L��I��,�	��I՟�ORT4y���<���ә+�N�R��0�x7��O�d�O���o�T_����w�����u�4H[wHϨk�Z�.f�x�	����Iߟ\��ǟD�	vF���4[h S���RR�!Ч�m��%#��?a��?Y���?-O��I�(��T$nx��dl�9rdUAFhʤ?�,���O$���O����O~���j|�Xm�ԟ|�ɍAhX�AM˴>��42F��-I�@$��Ɵ�	�$�'�_����'��ת+�0���	<cn�	ɗbɜV�"�'���'(�&��,D67M�O��d�O����;)�8�m��M��(��ᖠ���d�O(��?�����|����4�=����EW��  �RU6񫰮�O^��O��B�����u��ɟ �I�?��ןDvc�/��-	�<g`�,��Hy��'E"5ˠX����O|!���+13dȗiF�R�i�,�Op�z����m��蟈�	�?A����\�	��4kT���cB���#�O�o̔-2�ς���PE������I���O�R�'�r�'|���GHϦ:
����i�&����yӨ�D�O(���-�����O����O��$�O�� H�: ��u4n�"A9R*��#A�'bS�d�+a��⟬����Lp҈	"(��bJ�4�0|��E�ڟ �	�
Ǻ�R�4�?����?I��Rj���<q�(:p`��C�,h��y���PXy2!��y�Q�d�	ȟ��	Ɵ��	����5S1 ���*�o�8or-!7/
�M#���?Y��?A@[?��'+2N�oP4\`��i��Mj�ό�_)��r�'b�� �I؟��	� 3)V��M��GӍ0i��֡�E���L��?���?���?�����O���w0�ĸ��)_}a�9CqN͋q�� :Q�O���O��d�OʧR��Ĳiz��'�0��؉"Βd�`ǒ7<r��9e�'���'w�X� ��k~j���ϓtUt�tɅZV�܂BgmޔX�IןD���t�� �hQ
ܴ�?����?y�'6%$P	p�Y�[�ձ&`�"r�&����?A*O������)�4�ĉe�$+��`�/DN��!��O����O�y�s/��Q����t���?�S՟����f�����VMz!{�IVTy��'�����'P2W��Sr���*��q+/�L��\��)�?iF��4'��'�b�'A�d�O���'����=:�2�
�B�a���d�����|�O��O���ħT�� �c^�W�r��7���- J6��Ob�$�O�1V��l���O���O��䆸c�̡�D�W�[C�`��gWo(��d�O|�0��H0K~B���?���s_��2 �c���5&���$GS�D���8|�}��'W�'P.��"� sj�I@wW�\�2Q;aZ�d�(p�|�'+��'Z�]� pi\�`ĚժR��v�Q�%�<2}�u�}2�'�'u"�'&2�
����o`�5$B��b(pgV��'���'�V���n�'��!FL����q��J���by2�'�|"�'��ř��E>W����P�1�` �fm��Rx�	ɟ0����'�mk#a&�iYS4A�#��7H�u#j�\	��d�O��O��D�O�0#`��O��25��k��<4��.S3%���ҟ��	Cy��8C�������: ۤ&�^#��"�*ޑ+7 ���o;��O"���2$�h�' ��%q���CF�#�d�m�	Ry��n�^6-�|B��j�R��B���&M&���t��Hڶe�OF�D�O���C��O��Oq��P�T((J:�ɖ�!;����t�'�z)�$�s����O�����t&���I K�n����!^�<q����!���:�.�?E�T�'�~@ؠ�K�@@�𻤠$<�
�:@�g���$�O��\�+	x�$�,��៰�Q�9�4爮9H��G`ԳF���Ic�k�j�$?���ʟd�ɣO� ` �+#�8�v͘?O`��ǟ�r�����ē�?)���}F��b��4��U��]$F���b(O|�!�O˓�?����?Q,O�m�P�T3><�@ݠq��p���шx��H$������0%�������Ð�W;]A��S*D�~�0L��e�6{c�T�I���Ipy�ʄ�.3�����I�8,B�#W=S�6���g�'��|��'��*Yf��5A�T�hwɕ�u$δ`���71�	�(�	���'��)ǌ,�)_S�H�k�d&���d�^*@��D�O֒O��d�OQsU��O��n�uYi�)-%�Y��5\.za��ڟl��ey2,Ā`�P����矚��5Ό�Մ�B��&u��I�R�5���O���I����8�ԟ��Ҥ�"*J�@�͝��~�Z��'L剒	�
|��4����Ol���oy���S��Q��8aǲ-����?9���?A��$���b��p̧sZX��2��dJH�sE�E,���ɾU�fP�4�?����?9�'|ɉ'vb�ʼ_��PX�!þ�N��Ǝ̆���46�=����S�OU2O�F���'`��D�P\
�M3_�7M�O�d�O&e+�b�i>I�'�!��I@��pzC#�+#1Ε���?q��?��N��������O���׹�
�q�]"0�\ir!�U�*����OF)`��Hf�i>�Gx2�Q=i�jx�\=�lm���5�?���7��Q�����O����O.�oJ�ti�M3Y�����-P	u�H����הR߉'�r������.��i�X౯5=�dS�BG�y^Pa�IԟT�������Cy�OU��1<���x���s�.���4�̬#��'�r�'��|b�'����]V,�(M�r�	�$J:'\�0�dl��F���џ��	����'�� Bk+�I��\�:4I��E�j5�|9FBܢ�f���Ox�Od���O  1u���/W�"�Y�o��<9����lƊ{���'��S��`PT�ħ�?��Ds޴Q�Qg<^%6�\&��8H>���?	Sd
Z����fРs,��/��.xl5؀��"�?1/OI�2����u�O��O,�˓@v�������9!'�j�����ȟ��	8��"<�}�S
N�@�z���\+_ %���៼Bb�ȟ0��П���?��'H�%�|���X�ܨ��%B͚��Idu2#<1��t�'���%Z� $�U�vEU4Qw�U`��'�'T2D^>A���'%�ȟ<�E���rN	6p�5�ޠ>V\qH��#扫Q��'?m������}��H��B/=N�$a6��� ��	��@�'�I����|����?I�Or��&�X��N�(��	
�S�䃖A0��������P��ϟ��U\�H���J��Ĕ���*>�L=�'�b�'��|r�'�B� �h�!��q�*Y
ţYS�����m=*����O����O
�d�<���ɾ���õm� 0��J��>S����E����O8�D0���O:��U)�Dе@��HiÊJ�?�t ���E��	��h���(�'H|��C�(��ڱ&��}Abe
���	4
]�����O��O���O��Be��8L��	��d�6؈t�&r�'��Y����ҝ��'�?���GWr�[BM��4��I�B�:Nb�IM>A��?qrl�w������4��H��X-C�2z��ϸ�?A+OD���VΦ�O�b�OOtʓJ�BH���/D�0�1feN^(�����	�PQ�"<�}
��"%�:A:K�Α�ß� �A�M���?y��*v�x��'��d`S�����a�ʊ�X8�@¢�'&�H���#��70�B��0GJ�����C��M���?�>�@�@�x�'�0OL��+R*KP�X�B�["�5�!�� x 1O��D�Op�$��*� T�����M�f�`��OXR��_�П���g�������&A�?�&�I��ۻ. ��Xi���<���?����ڸ7������[	��Db��4\$(TN|�I��<��d�	��8��.S�"��T"�fd� �M;(à̀% 9������Iş����d���۶�M!��"0�����H<h����?���?����?)����O�h�6��<ʡ�	K�^�s�)�|�r|H1��OT���O����O�d�O��)JŦ���ß�8�ȴ)����iQ�ɱ�������	dy2�'���� �$��f�&�GcW;h�\H�-�#s���'�'���a2 6��O����O��IIP�}�戟6@N�|��h�J��$�O��?�t���|"����4����WB\��H���1�<%H0��O��$�O9�VI�¦I�����	�?i����tx#@��U���܋r"[�/�HyB�'� 	T�'$V��Sq����i8MZ�D�}�e��ϕ��?� N�Kc���'���'����O��'��.x?
,�W��+X�Rq��5�� M�W���|�O��O����B!�����AE��B����N�X7�O,���O��P0I�2��O����O����1��9Y��\(Ϥ�±L"$p����O�˓)��LPJ~Z���?��l�B�X��t�-ɥ�Q�9�������?!CLD� ɛ&�'���'%�~�'��J��"����Q��5�Х�/OԜ������I����I����	��<�J�U*�Y�Əg�b��l\ _L��Kݴ�?Q���?�s��SMy�'Đ�z�Z�[��P�c�R@� Ӷ�;�yR�'���'�"��DAj���ג�9�t��	#�n��ӧN�"�'�'��'\��B��j���c6�W$��)�?иX�w[���IɟL��my�~�.��?���<:�ܤ{"�C�t�r9[��\��?���?A���'�1O����,��2J���lM*h$ґ���'���'�R�'q���\>9��ɟ���켐�N�c�f��4)�>:��h$����~y���O^�a#JE�X���7��E
���<A��1����?	���?a����D�F�2��=a�c��8 l��D�O���MFxJ?ݪ��G��@�k�`�e�����O�hWN��u�	������?�O<I�D ��ׄ�d4H�"�ҘWԜ�x��?Igc�f��&��/���"�>5���'���'��m�g�&�$�O6��x���&FKƜq#b�����K9��'�JLq�y"�'���'[ � t���-z�w�܍H2�1��'��}_�O,�d�O��O.��F�Q����cӞu"�8�F�<�	F̓�?�����d�O�`tJ�'�4��@@�&J�����3����?���?��y^�D�3��l+��y����i��S�
O\ �0A�6?Y��?�+O|���c��	
�^��h216�̘,ar_���I|�PyҌR�T�^�rR�]��Ē���E��qQ0����	ԟ���ny��'�*̟��DW�rܮ �ի"��hY�K����O0�O�˓.d��9d�]�V��"�p��GN�.�A��,�O���<���5�Oh�'Z�tĒ�zl8�F!+X��+U� i�'Y�ɔSY��F+�?��T9_���QL�ψ���(B6Z��P�ʤl���
+��¤">P�F��m�5c���y�j�C�M�DN"@�<�1�Z)��̂Gvj��O���|Γ�?!��R̚��9(�x�#Q��q�!R��M37�i����OD�$㟦�����=M(Ȕ���� ���w�,"��$:G�B3��4�1(��N3�x{A/�'yX�Ì&���3��F��!���"�Жu�΄�փ��69!�$�1Oi��&C���X&�?ef|:�$P'Z��MR$M͌mC��U�Ģ=V:e�!S��|xw�H�A)6�z"FY�F|���F�iD�5zX�FXb*K>z"(���)��q쉀*����`��*&$ꐪ�-������N���:%�Ӈ/���1 U�.�f1A�\�i�ܡR�]�&y�%�̛�u���T��OV�D�O���\�i+\�z���Fx����%?M۶ ȰW��GF�)����Z+^b>Oęv.����% �^Ȕp��LX"S� u���ö3Y� �TmK2� �|jw�G���f�<�(KLs��PZ�Ƈ#�����E~���?�'�HO��t�[(7lޑPIP_
���"Op�bԒ<l��k�g��i���y2�O����d�����'t�)� �qH��ĉ�$�*�ҙCD�P��Ɲ�7�� )!Β���۟��	��uw�'V�0�~H���Ҿ���)jJ�C��IP���"��U�`�G�V�d�s�-5<OP����G#����5���`�ҡ*��z�FC�;��Ls�Iԁ3���2R$��WL�T�P�/����hg�!8��L���e�	��uf�O��>���'>B8��Ԉ$��y�nU�S頼��'!9��H�#�aC���K�~p��{���>�,O� �S&AS}�i�,��ץ�9�$5+���8%�����O���%i>���O��ӈ���!�$��(h����סE�Yӧ`�6� "m�*�T�����9�B�"tb--���՛AY�}q��9�@Ě/4C�'��Q���?��O� ��`ݨS�P��N��F.d3���*lOhaȲ�N)�*����X5@,2q[5
OΙZ��Γwer�P�C�bxv�M܇�~R�|��hX���D�Oj�'G�l0۴7���D�!8�*l��jZ�xS�'(��4�h�G#L���	Hc��O��V��B7[梔3v�	�h��c����$����$`�.5�N����A�H��3��1I
���IU�:8���P@_��VK�p�\ P/Z~B͖8�?���h��6��+w�Ϣ4r�uq��4�>j�"O��@�vB��#
J�k�+3�'���<�Ӡ	�\X��{���$��q#҈�K�7��O����O�U�@'�o���D�O���OGJ�]���v��G���7&�@�*�Z���x�&��hi QjAj-��|�GނX����I�ڵ@@�ݚ([:�mD�/�8�/R;��c%�ȩ2ir02��u왩#�Y�p'XUg A�!A<�M�i�f�@:��,Or7mȀK�	�W��7#@�!w�U�����	r��h���SS*W�K����-�1*�t|�W�O����]��4���2�'���ٝ-����!N��z�4ℭ &��UɅl�B�t���L�Iџ��Yw��'3�I(-w@�l
2M�0�A�A=Q6�D�Q � �H6���D���d�4�"�	`�&q����Å�ޑ3�̑!�6��P��䌑%n@�Ge�Y�N�cp�J<)H��[��'0R�'6�T����z�o��%�ԏ�(NX�6�$W������D��#�5)��A���#� �=Y��i"T����J�;�M#��M���N�Hy��[�n�S��X$/�b��%d ��?�����4�]�F�F@�D�\�bq�kC 8t��1s����Dѥ ���3��E�����s�Z:6L�4b��+�.:j�Dz4ǚ�=,���!�f�'l���#G��즟��,#��ɩ�I
&��$�wɤ�(����?���HаK��mS�mו:&�1dk�y(<��g��^�ڙ[��0�XI�3iɽI�������Ē�G�H9�O�W>�z�f즡x�g��b��TRTg�7@V4ha�
�?)�M&�z�ÎA&�Y��)b�*6]>��O�|y�CKж]G��)O	� YCN<�4ɝ�~����.�5V���u��;V��aXǱ|J� _�j�8���L�3��=@��c��gg��D���ȏ��c�U���_.\�δ���W�l^(0�GM%��xBcۀfw���ڒP��X�`�H#~4��=�'D�Q�X��(H�/�	�2`�ZR`#�%ى����'��'��}����^S��'�r�'?$yf��DjR� �Š�q�@ۻFfvy � ��w&��T)z4�z�� �St���:r𔀖��1FY����T�}��(�Ԇx�D�nZ-��-��h7��r��I�!kT�@����HW�}��A��,	ڴf����'�dy÷�����v���r�Q�]@ tI�ʍ��� �*^wH<�qᜇ:�`��JL&�Zlk�Wh��Jg�'��`�'�ɗ$��Å"Ɲ?+�����L��2}����#~ə��?���?�R?����|Z@�:{C�������>�I�`Q�I�6I��"G�o-���ڴ=FƼ��	6 ���&��$� ����F� t4ر�	��_��@3�j��Pl`	���@��E{���!e�yXbf� !	j)��	49�2���Dg�a���į<����'�d���.�� �>{5Ɓ;7�R=P	���AG���P(]����t��T��!�I��M�����(�&�m�㟜n�'"@Ѣ�)ܓHQ����	�L���)��?�mO�?���?�����x��Х��}���DZ+be�
d�2n��ض'ȬIl�d+���@1,�%�V�0��%��
Z;�|���8	�$��"mXMu�(���~�'�"����91��U�Ҍ[���X��(kL�,a�b5�	s؞l�7��/�����
�?�ά��Y�'5RMF��'&P ��bn��"�̔oNvɪ� ��`ג�yꊔ
{�6-�Od��|Ҳ����MK"�J�6O���OJp�B=���Q�$?��'�xĭڋn���)���-X�T>1�O�<�{��ٸ&��]K�l�}�|�H<!�Tt�J}�R��>b͈�n�#f�D�&?�ä��,4
I
�閣,�,�C�j1�D�-G�b�u���m�Ο�~�X�FР�ɜ�A8��AҠy��H��wX�`�U�ai�h��C�R�㥪;OxXFyr�Y�Ƙ�A�U�Bhv9[A��#D�`� ��O���Ob�cq�Q�f����O��$�Od� � ���g���,K��p����U������%DBp]˓ Bg"��m=8�X��|bGk�����L�O6���,�Ju��%�H�gJ Y��N�8�|�D!�I�T@hBB ��V*�8�w� ���恵[��Mq3Κ"h�]�a�6�	� h����x��2���!_2@� re�y2��7 ��-�S�V!(�zċJ�~��'H�"=�'�ēH�c$Q�_@���'�8`3^��tUU�~���'TB�'�B'�~�������c�0�pR�0�d����
��1Ҩ�A�1՛V녴�p<��@�U����Ό�E1�V�#�JzW�/v/U9d$Y� T�8S��L��<G{�]0;R:��u�C�P[by @K�]����?Y��?�(O2��$�ɯ~7����j	�I>5����0�^ f��X�,����jC��*"qO�Hn��ؗ'W�R�er�X�dt���9w�U�	��e�1�@+n�S����$�I5� ��Iҟ��'(�DU3�k
�$e�$��4���R���Wքh0�Q�4G���V��q8�PP���T~�P�t-�,��<Yb����-�G��2t��a	��v2��s`ҞH��"<�3)�ȟH��J}�JV���� ��ذ��>e]�����?������O�<��Ċ��D�8@A�q<,[��"��|
SDS�O���q���m.<��A�����������OH ��Oy�P>�㇆���7�N�I�\��o��-!6�r��\/�?���	��D���!/�՛$h�N�*���mڠ 7g�`]�i+�O�J�p$���u���5�hy11�"�:�F��h/c{ڭH�J Z8��i���ēC��t�I��F��i�X�Y"*V4e �ٻ�� B혴� �%$�4���D�pv��ۓ��w����B�hO��Cb�'���eժ�n\�A��(RdۓMo}2�' �hJ�f�m�r�'mb�'��� r��-ыZI6�x�̐�bQc2'��������^�=�r�#�1���'�t�sNɷ:]PY#��̙���9~�J���ϊ��1�gу��O�&���Ѕ˵Va�@��W�`���i�'�"�'�~�������b���$�!rn��@Č�.
�5�!�wH<��3+��Jĉ�A'`���X�d�b�'�� ���$M�U��Z�lԣFS�3��G-C;�$[�$V^GL���<�I���R�����u>%8QC��q�@��$��:�P�'�V�5��`���0x�R��8}3n5�A���q�Q�x��"���2L��Fb,h��P(D:Bhz,P=��`b'F�|x�Q��%�;��#<y���v$�+����!x���v�n��	9�M�Ӳi�S���I[�~Z�a%ɔ>S)@p�dG��@(H|��\��e��H�K�5�윩�%�!K5���������'t�i��nt�A��Ϧ��E�<,!p�	�@�(�������?A��~����?i�Os�A���ē)|�5aꊥY�l��$R
=����I�|��c�<���K{0��sM�(M�>Z�//,O�hW�'�P�`�3o�BR,jӦ��~�������Iٟ��?��4aװp��R�D�}����a(<aGd�g�����<+�R��� 0����`ybHݮ.e�7��O
��|"����M��
��raXV�^#5�f4G�Լ-�b�'�h�[P�jӔ����'9�YS�f�TR?=��EL�z΢���"�gf��"`b)��M��4�G��R^0�P*���>	�#צ;�P@r�H����&F+��ޑ"!"ll���lݟ �~em�3
b	�'ȉA��"�]ܓ�?a˓io�xPe@]���i󮍆mH�<��*�(O��
]H�$eU kK�e�1�$DX�U�O|�d�O��agU�UW�D�Or�d�O^�*a�D�EoӱgZ7N�戚��S�R��<Z⌬��$$$�R$3T�xCU�!\PD�%���3������U��#�ȉ��Ĝ�Q���~&��r��� Bmh��&�V�(,˅��+O�	�<�ta��S�?�>�0#U[��0�r唪|�0p��h�<��E�'G��p��0*�x%h!�j��b�'w����D[�V=� ���?!� ����dQq�^A��A�I۟4��ԟ$�Xw\�'��)M=~���2�"q1D�F��z�Y�$�пS�����K��}��ɱF�xU�6�ʤro�S�Q�b>r��mٮn��TK�@�'uJҽ ���R�'��qq ���X�g�O=/�|������?����䓨?y����'�B�(���=G���Y�X9�,X
�'�؉jF�(�BYRjڐTE�8�{�>�.O dMEo}һi8�:G��v��IӖkLy,� ���O����*���d�Oh��.G�fy��)�iK�A!F�s�d+Ug3�rt�I¤j��5(	˓7�Y���W�z�Ib�d�_�����'P;S���
�"�>l֘| ��G�
y�F�r�'�N�H��?i�Ol���cՀ?���K��
�RZ�)�����O��S7�n\��f܅g_�<��5���DP$G�&�q�$"\���za�эx�i��'���+�H�ۮO���|b��8�M��$�@;�4��&νU�Qa��jB��'~DP�F��{ڼ(��!t564ӥ�AӁ	E�� h\r霚�xa��ȀQb�LB�xb��,����$��9"@�4�u7K1/��;;�� G�T�79PM1f�Z�ZO|��r�'|���ئ�����N��S'�IT�P�+��x��T�
��q�m_:NC>Y��
D*B�=ͧK�Q�L��@�M|`��/Һ*}�t{0���,��f�'"��'�Bx����"P+��'5��'_,���X�}s��:wi
#~V���C�jtDE{����c�x�C��x$�ԫ��	?}�͕>�����8Bǔ��&�K!�貂T3�0�7k X ��Џ�Ė>����%N,��jqn�S�n��܀{x���<?�!�S���SΟ��>��$������hW G��#C�}�<A���p��,+�MH�4��	j@H\N�$Do���)�>�`�׈ �)��8M�iWǑw,ub���BD��')r�'��'�?I�O��YJ�	ɵ:��h�/$/��x�7g�=�N��`N�>'����#h���0<��ƹ�x�@����JP�0���x�����	����.�+,���ɜ=2N):!��s���:w�G?���&��O�4l���M�����Odb�X�IS(�@ ��j� q�<D�x�m�����D�Td� x��
<�	���d�<�N^�
�	�1@���CD ��e?�Y��i��?��p�2�9��?��OB��yT���TY�A��˟�17�7L���� ��G��  �4,O��@f�Q2v���q�&5�?	�#(n|�2`I$>�5����{X���$E�O��oڶ�~"�ǅ"6�@wHֳB��m)Fi\���'�r�'��W��
M�;�+@�a��]�
�' t�CׯW�D�𥋀)�(w�F��SKX?�,O8��b�ɦ�������O��`'�i����'/�'�|}�U���U��钮�O���U�l{b�0'�\C�|r���$��b,!=p��E�ا.�ب:v�x2�_*|}D5��|����>������A^��'��	�ēs����I��M#1������`%oV��S�&W���yF����'���'��q�([�O����"a�}x�rQ��;�@���r5o�t��4)I?<����P�I  R����˟t�	�D����hO�q���!�
	E�&�*5	�A�:�R�o�;�N�ضk��A��xr%Ǔ"Ӫ��c^8>� ��Bw��(�iײ2J:9�Ɇ^���H��L<�0'�V�j��l�"G#�<H����Ta���O�	�O�c���v*�`���C�\�vE�;WF2D�l��$ӥb�Z��+;xc��0}B4ғuL�	T}¦I�!)���c	ۮ<��={��=l�B�	�_�|�(i̧%7�8`�����B�6m�JfK+G���,L_DT��=@�Y�ꍢT��D[W���}D��ȓ�.lDMc��O�Kk`]3�F�v�<Q�	��;,�x�N����M�p�<�m�L��x%5G6f�a�@�n�<y��)O�ּ*�@I�e�.PabdOo�<y�F����K�.1�4!UbLn�<��HO.�bC��)]lΩ`eiNh�<	5�;#��a�%^*H�����h�<iqJ^(]�����P�f��ěR�Xe�<U:�60�HO�$=0"��h�<!V�U���H[ n$m�ZH�σr�<i � ,Sb�1S��9M2�1x[>�C䉯l  L�Ve��#����T僖1��B�I�V�:�3"�V �yH��^+˄C�I1�<�;�������F�>�DC�	8Sr09z"�#w�倔lܽ/{�C�	E�����Խ��A���ڨ#&�C�I'S��Ë��\��9�&�u��B䉫,"԰��+J1B)С�ʡ�fB�!1m�l�'C@.N*
qw'F�DB�I3+��M��f\�A�řp%�E�nC�	�/�4RA��iQ��9�o�q�6B�I.	32�qg�١r��! )pE�C�	_����e��.�B(��#U#6��C��[n(`���$k�^t�uϟ-hI@C䉗H� ��!#�F5J� �/K�B�	�ҸS)��U�,���EizB��8"�)���	�)�wat=��6D�� Ĩ* �&<��0J��ǲQ���Z�"O2�h��W+L�,
C?.u(��u"O�`C@�"}��@�p㝇s�L�"O  � 뒀�|:ՄW�����d�O�P�+P)�0>��G�?�P���Fp:��ª�G�4��	��Tq:��	�Z������Y!Ǻ�#$W)ff
B��(JV�dL>)u0�!u�Ҳ�0p��R�0� ��Ӎ,��Qݹ3��`Ku*���bB䉙PD������
7�xA��U�p�9Ť��F�H��D��'�������C��S2�%��uz�'h�5�"%U-���xpG�&v��uX�*W\]��.�r ��DD 6��c%��e��p�G�z��{2.�y��x�'����S(���HH����=`��h�*1D� p�25 �ҁ�N�c�R%�.�	�A�p�a fżfh�>��gՃN:�)��>��TE.)D�8BE.W�ܫ&IA,>,���Ɇ�(@�"U�����	M��~�,ڄ��T��$�&S��J��yr�C%j ��I�LB��$�*�bڟ�?�&��g�*��Ah2lO�puIɑP_T�*���*�ZP�'m��8IԃKMr�K�#����B�~�Ts�]��y҂�()&�x�AODF��)b��=�(OBѳ�������BH1�8��� { AI�$�L�<�C�?]��\8�
�l$���JN�<���Z�|tFq�sl��q�n�[�mXO�<�4&A�u/�y(��tz�a�a�O�<!P9a�0RɎ�)p�s�]F�<��_�(>&���	gTfa{�lC�<��nѲZ��A���T�,4���C�<� 
N< �(	��	[�8�P�Z~�<a�NJ�H���ԅM)����,S�<9Ջίx_��:�� l��U�a� @�<	�N�)���p�b<X���K!��~X�����Ey�r�'�|�p��?9Ȕ���7?���"O� u���B�&m�G.F܀y�O4T�s�W�l�4��',Ϩ�cFI�M\��jz� ��M90
@�����Xw�pU$L�N?:��)O�=�5�P�F1�1O��#�� & "�0#�av�j�x@�64�O�Ol��ђć�HT\Mg����H��hChP���T%r�}b��|���y�mw����(�n��L>���݅)�j�Χh���v�	���I�*O��Z�j�tnVhz�Ša'�hj��';���;8�ٔ��$Y@+W��l�����#�M*�E��E�2uIؙFk�9<�Ʉ��i����O߲@��Y����>B\b���Я|���$ʍg+h�O�6D�S`�3N���t-F�o�y�.�?T���HJ�h�����$����d- �&A��6�v�KS�CB#�ȚRʬ4���Y�
ϖ�q哮wlfm02��YG�!��S�o��A%#� �>ݻ��^7 *��V(�dx�x��,���`I�덒,$�`��)������U��0�҂�Y�Q�,����xa�͒+(�P��x����*͈P����k�4 ��+�O�	p��Qb"ܫ�+�����7��+0�䈲
C>L�d��h�{o��"S!O�)�4��D˗����WK����'A^�����b{$9��N�V����d�V$���̎�"�l���U����P%��C��Y���rD{uN!T�^08�Mݤ,�|[���Q�� R�?��0@rZ�����Mo�j4�,i�� �L)R����G�2ʆ  �E�����Ӄm�~q�O����c�N�9����67�Q��-]=�Px"!:`�rd���C�lb�:v�P:XR�S��F90��`F�*e����a�8d�fL��!�:dv6-�"q��n�		�,��M3�`PA*���a~*�N\d ���'i�r]�I�>"����tr�D궎7kS�(�bN.y��4H7'�m�fm�F�H�;%��OV����&\�>�0�ʦ;V��a��2�@��_�O�\��'�;戅h�!6B�P�j��Eq���"���%/zyD�i�Х ��pRnA���' �A�Ί�E�:x�r��1��yJ�'T�9����͜�84NR)�2��] K8��A�8�0`��K�Ūċ� �&Dh�a Qi����'��}r����@�o+L=E�^�%� U��@�}rP��"T"��S���J��J ���Q���+��"�x;W�2�O(P�ՠ,b�J�b�1�袖CG�NvL�V�$w^Kn	,l5l��4�$O�x1n:�pWĨs[����u�'���q� #��}4c!ܨPa��³Xڢ�`�S+maF���‎H�&,���� ��  $;r�$ؠk�`xI걒�HA�W0W�� ��#ſ�=����q�p\ ��تv�.�2oBq"� 6"O��8���d0�*�Ξ0=L�zv�O�� �A�v�O�>)�7��>�!rD�?a�B���&>D�0�GeW�w�.�
�I�o��-�v.��g�r�Sϓ����,%��H�k��mJ�ȓO���p
�=�r�C��(|D��B���3�Z
56U2��$�(�ȓ:�L�� #��k� �I�Ί��̇ȓ)NYPt�F�*�iD#KS���ȓZmT�#㞯u઩[�1rjpe����YE�ϧ� ��˦��i��"��@cP�;1	|MR �N��ń�+v�@��_�`����-΅)q25��S'�pQ�^/Q}�		�W�2B^I�ȓ*���&%˨�D ��.�/�$��ȓ/������W�ف��IfZ���J>����gX���|�<�6*.�nH؂n��n��۲�w��|�v�H�}�Ԁ�bԂ&TI�t�ìp`$����z!a�EB�(�@E�I:d�������O�L9���qI�9k�>�d�	-;��Qi�遰P�b铔eT��y���x�@�7Eڤb�}��']����ؽ*�2=;����<����[l��f�y>\�`�IO�ǦB��0;���X�m�^�p��+K�C���3\�$�a���*��BJ|�>3ȆOm>U�(�m}��JLE؟��@&��6��i8T�H���Y(2��.V1ڠ���F2����ɶp��H�'�H�ZQ,�5p�^#?9u�g�膠S�\���x��]�+�$���	���iԎ�yr¢\RZȸ�"M� Œ���LC&$�	�/RX�4K�.}>(ь�	���3��ŖHZ���0�}�P�3D�D�aGK y�.I�e��;��tS�O%r��ǬrӮ4�'�m��ם���O���4	�F�n]H7��*$��'��+jߟ���*�%
z�H��k��ز�O]����a2cڎ^�2y[ҡ�4n�L��D߫ʸ'�n�#U�<ѷ�[���y[N~�N5 ]~��a��8M�hKE�g�<ɶȄ�)��`!&�;f���r�Xi�B�=! �/�gy�IQ>=��UP�"�kl��ER��y��]2�z���!�'m�XyR
=-��Q�J��0?y��W�M��x�w�V1`��Ѡ���P؞�2F�t�D}��=p횘w����� )[!��Ɛ`.=h�̕����	��!A(!�$��Wy�ɢ�dRS�j�k��ǈ,�!��ٵ\�F�U쌅'�.�x&o O!��&p��@�a�'O-��;!��'q !��;b`5�T��7�<3���">u!��%+��-X��O>*�behn�iU!��й:��D4��+�OW!�DǢ���C,y�L��L&y�!�dA'^��T�gܯ}�t�J�*܌X3!�ПM��&�tU���X!�,��U�P�L�qOh����Y�\���h�^��
��ĸ�Q�0\Ov���Ļ��d�((��9���|)Є���2��X�-�"}z�0��v�lٓ!�Օ-�d�).#�
��<���\�!��k�'�XM�������"�Z?IA�1D�2h�PjL6j�N��֏;D��Z`D�	/6�!��iy1D!O�T�:`�Ħ�1�M	V(�P�Y�ԸO�D <�#�F��A��9u�Y�e{`IP�O��I%�#(0QR釐o�,���؜Qp�z" �M�M��`ph)��J�<UM@�<�/[�^&�ًG��	���P,�mx�У7Ĉ
��x2�iT�y{s���
�ꖇQ D��@LN!e�F���*��jM��ɶ2�����l�0�.�&J��O$���W%L�y;۴^Qܹ`s- s����?����<���2�>9�`��9D��W�P�"��T�R;�ٸ���| �;ڴ~��u
�!B�����.擵��λ8�N����t��!�& 	4w���+r§J�O�PC�G50,��4b��2��C�%R�fg�1:8�����"y@�tDy
� �0zW+�-8l�w΀�{��!��'<x�.@�~�mG�f�Aǩ��0�W:P��l[ E�p�~�a��O���|�d;d�l���iT�b(`b���'f8)0J�䖼�J���F#B��'f;�pV�D��2�X�+U%N@�ȓ'p����ޘ,Z�1��AL�,H�k"�P}��Q�g qabX���OI��;G�t���(D��4�#�)����ȓ\,�u@5��;�lбtf����܇��f��F��O\L�ą}:Y@�E
9�,"Oh�#,��TC��bad]�)�u"O|2@�IoT�E�B����"OL}�ЦM��z�S����Ł`"O���󏜾X�^�������n@pq"O �X�Jٚ#�,"�i�%�*Ѳ�"O��ДJ��6u��h��u��� `"O�|q���W���9���/����1"Oj�+�+�`)�!�
ŰA�F}�v"O޸{�,1y�x%��'I�7��!�"O>M��ܲ7_9���>�@e �"On]�Ơ��TƖ���-؞��q�"O�m��K�lK�@����	w�"O� i��[V��rޫ*Q�ɂ�"O�I�G�����C�a?|iVje"Op90&�#a�8�R�\����$I|�<y��Q8J�l� �"j��09�H��<qDR�774љ'Ł�2�HP�p��~�<iD zL]X�$��mG�s#��|�<����@�D�س��� ����q�<�+E� �=�h�~��� n�<	�"D;*�j�����A1�
�dX\�<I��
:�]��٭>�i(� �s�<I�CW� ��|�B���Ys�<!�� [�<�*�0o���i�s�<ɶ	�9^ЭX%H�-B�N��$�G�<�3h�F�`���㈧���C�Z�<Q�U�z� ��	H[�4[hP�<��BD=x��:ǣ[��X@��VY�<	�N�V|�����X�8���Y�<I��A�OHL���(��ua�	�N�<1Oɏ��X!�	�a|Y1
s�<1 ��8M�X�Yc� ?�2����Ѭ��x�J�3&��p�14�"I�v.
�y�A�r�B��4��?$n�����>�yҁӸ��鰮��D����!�yr.�%t/
���2�T%r�lU��y�K�a��D+���)�~E�Q��yr ��ݠ���8U����p����y�Mn�x`C'	��E�vd8�ܑ�yr���Ds�;���,��Z�g�,�y�h��08pȀQ���QB)v�Y��y��ם� �Ff&K-0)��(��y�C΄;�����قA�.8���yRN7 -�	�fe�)4�K�mK�y��MXf�@ *�y��ǁ�y��>�����l��fv�sFL:�y��݂%\���ϟ aF6*��yRM���QbIE%T{����#��y��<aM�@��-"0�Z!H]��y��5L��@&�C��j����yr
ȏg���L��XHS��J%�y�LV1}�ur0�U*��ɠ�*J�y��T�tN�Q������)!��Ɖ�yҮ�]�N�˃I�"z���B���y�]
-����G���x�q�BE��y�I�U����$l�T��LB��y
� �E#%Smpݙl��(`�¤"OLx��	ȮJ�JIc��G< 3�J"O�܋V-Y3�4{�mβ]���"O�� EM1>��ze'��) ���K�A���gIO����	�O�3�������y.���(�5�Zyq3���hI
����=���X��؃�F��%d�D���z}��ٍ{��~��N��e��E��4
��b�
8z!�[i0\8#�'��5s�Хs"�)��ŹC�j�;���{�ġX�dQ�W�ɑ$?.�)!�'����́��ֽ��Z��r�#�F�2�v~��"//��]����LWI�d�1, \l��OJ�!��3)���U@C536Q�ë�<R�|1�&g
��$O�I!M����@U���P���C��!���Lr�8���Z�L5Jh:g\��%"c� .�����cЫK���
&Ň!g�%hE��˦xI>IԂV�W:|#?Ypَ|�&Us�gӺ!�& 86�ʻE7�̈�hS7׸'H�aI&:2��ۼ���-�h�p��+p���hF0([
�`5�'`Zp'D���y�-�';���2s)�
ɪ + �ε�����O1�t� ��T��샽������@�N%�0�ٔF��ȡ&֥ieQ����DJS�LkP!�X�r|�Ҏ�O�A�Wb<� �禘�9�l��4`�x�"�K9�Dp��5�
�mC��	�)�m�'n�6��YCӋ�l�I1S&�K��
��a����LU��P��`Z�.�� M4?8��u�\;�'R�A����!�XPZ3)ݕ����$W�8��8�F[hK�! !ܐz*r$�wL�G�������!�O� ��Ô�� u��k],p��c�
�L�+��'\|�ݱyy�B��ܺ*�T`�Ɔ/&Z��ƽQ�'>L�jqdN>?]D8��};�c5"��~(��ד*DX�Jt��fq4u�D��cu��r� P��Ӯ��">i�)@�#,�tG$
�`�Q���<1�H�"��fI�5 y�sf�u}b��J�]��˽sC����,_���'K���G,^s_��k�/;��i�
>t���_:�����ʽVY��ASiL;3��#>I�N�h���ԬT,��K�&ӿm$ �����'�D��/<h��g��[v40(�H�"b0�ˇ�� <����	,~B�˒�E#AH��a`�K�.�.��	F�HÓx:M���<��t��鎨g7����h^\�B�F}§X��xr˚�^����"U�<�6�F�y]R���ђK��e����F�'^��j1�[�^V9Xv!B�,�2؜'��i���6Bz��4E��U~��s�']б�c��i��𧆏�c$l�{B���5&m�W�τ X$��1Lÿa�Z �u#�O�M
�MBYC4���m�S�	��4H���%}"ȉV&>���$ ]�P0��Y�y� \�T8���}nZ���5��-�n�UF���y4�M�0=�pM�%L������P��,ۼ%�۱��I��t٘b�ɐTX�Dr�� FtH��"#^�Krڕ����F��e)���I��H��&#N��ڔ��4 �j�҈�O2����D�O�@�����!�I,9���av*؇��i�Z(Cc�+Bq"�	f1���#��+�*ȱ�)�1gb^�b�ڪ|��oZ=^ �pb�OL創.��Y��F�1ek��g0���#`>��1d;6֙y�	C(,��8 �K��'��9vꇪ4�Z���'M�e�˟��y�ꖈpZ���Op0�w�$�s��� Y<cs�T�Č�&�4�5�#�O���t�O�&=J2�8v,M��W7C�Q�3�J�yR��&f`T1���QGyboj���4�$�JME)� t�"�A�M�'p��<yo<dSJLA!� 4~"7-ϙlG�,����(qq7��?j�RRF!Ѵ0�	���x"�C�m�(�Q�'*nƘ�CeO
J(%��O�(p{q�	 n<[3-^=mc�x��M���n�r�֓uS���2���z�dh;��������?ɢC��?) O�I���`��Z]�!� Dx4���
��}����E��'Z���ӄ����6���.`��0!@ia ��-3J���#f�00
�&p��yJ~���ɢ �:����&��e�*C3yd�H֧R�g�H���W�#�F���D9#�Z�c4$�Z�>�À�H0	�`��M.��'.D�O��A��,�&@� |�R*�aA�����3 z�Z��-n э���-d:�}D�0m� �B�R9��4�����%�0l���BF��lq�	ïU}�Z��Or�ff�	�n��Cd��%�6a�s)�+��iE?f*Ę ��Wn��3�^w?��`�J�)`�|��2�� # n$r�K�myR���~��<95�0+ʜ�e �;x��t)CV�W�:,J7��;�ཁ#�]��t�81�rݭ*wN'��|�4��5#F����ho:�0��T��ٖ�NX���P��??��m��M��X���%1�~�	���^����-�;0nqR��V^�'7��F�"o|�LВo�\V�]��a�I#F�۶坩��g�2}�i�	wK���$�.6�p���B9����B3�fz��ߣ� j�J'�	: �^����z�~��������O��8�C��9#x�"���a��-�@$��wv�i�1����b�ˢIĢ�{cO��Y���!��1�	=c�<Lf險7�J�Iэ�' fl�1b�Ӕ!��x���T]xy dΦ��rA�)mt���ϫ<9����Sd�<ɤHυ�Q��3zj�nZ�g�4�@�
���	����9P�V����%B(+�0�$���l$�(׳���p��>�O�Oq��av��c��lhsk͑1u����/?�p=Ywl\�:�0��Ç�3���3`׻E��<(�G�(��r_��@���y�2�Rȟ�R�@�]r�e��ȉ��� ��["��"��yʶ+�4(v��ؐ�	�M	��Y&��?b �xȲ#�h����ӏE��S��W�G��QL>,�ڠ24��,%	��y�'"�AT��9f(K�'�:`(	�
6�剹u�lqIt�	}�`@se
e��[S����Q�#�!t׶�Tn���Jr�%��b5?��u��@!˭i$h�Y�Pȣ �OZ!���Ʃt�4�.�P��(ߚ/xQ�|�� ^<Z9��l�$+�@���̷{��ġh��?��L�@	,�T?M$?��+��5��uc��8/g�hg��X8���.O�x;��Pc������6��P0���+�b�"��x݉'���E*'��l�%�q�U J�`t�ê�M�T�w��d}x���f�P6��?�
ڦ����@�[H��P�ԟ��'�i�f�Q�(z���f��)2iЂ1�|��+6a�±�(6����J*)��� �nXCҦ)���YԆ��V�,  ���'�:��e��xHi��"0Z���	�	���n�<$��)v/J�C�`P��ڝqi6�A���"w��z0�Ii��E{R�
#;�$
aKE�H�V�*c� ���1��	A�ɓkb��KΣ6����e [T��5.�1�F~�'�CYB���ȏ19���ԫ<r�Rx�&)ʐP^�C���k�IK�4eY�۩<h�a�ӡ���x�t%&���"*>H�$AD�)k�����Z.n�< ��5}R��!|��G!�? 0\��-M���'( |��%\�\��l�O�.:��a�
ӕoX��U�'��t[�/�z6��0k��c�6l	�]�e}�(�o�/H3�H82fӶ�0<)��I�a�@�w�MU�8X{v`�vvF9��uS!���#���)��Dׄ���V�OL��`Ţ��M�tLJu��n\h����9�DUM�ѹRa�T� ��dŷ	FD���;�O��J!��/���4�F�N��y��%ՌV��#<�ՒxҦR70V�xKٴP�y�3,\���}� d�Gr$�H�Ǆ�i4џ���a��A�ȓ+E>SR��
S�S'�`��=K�`!ʇA�B}^�rN>�I��^�p���*&{ر��<���)(O^y�`Й:� �%,>bv�R��� 
"�[���ʥ$�+c�8W�+}�S�02$���3 �c�ِ<���D����:�	�f���gf>LO,<��\�,��q�DKޔL���'.�dʖc7h��p��E�iH,=N��'��Ht@�C�j�"6�PIY��hw�8D���nD/n6 <�ܞ�8P��&�	���G�x����l�T(�5�Q߄Po�I[*B���~=~�Kϓ	�*@���>�~�I�E#a<K2N�� ŌQjJ�3�ɂ-Z垱ac$�*L�O�<a��8��O�|�U�

�ZeP�n�$𛂙|m@�.$񙆡ۇ�`p�$(��1�Ԩ�g}r���S<d����e�:�D,=�j�8�KF�,8�XR�Ӱ�0=QŃ�7d>�Ѣ�@ $�J��xA��S9m��B��ߢPs 1RM����}��
6E�N�Z��cE�D�%m֢{���7��8zr˟78����E�&V��0c�C��WH ��O~���a,�� ��F�;�X0��Ή�"�H�%+�� ���'��J�-H�!����{b���R���0)�L�S�\�es�����,���J�*�O�4[2�.h���֣���u7m^}�}��� k�2R1�ȓ.W7a�.�<ɗ&G!!. Ѓ��+0f	a���x�b׽<��@�\�Ib���_��� �^<`
��-��d��y��bM����qO�o��z�lќ|2"Xģ�^w$}���[�7M싧#������O��GV$��)��4N0��a�I(<I��A\!&*�~R����?y�
J
C� ������l��TF�G+��2��|RN��򉛯+�4%��&�|R(M1��Sq�I�dĘ��e�E�'���'���9DN�9?�6YR�)@��ҭ���@�⃄	Ɩ���	l]:����,�H��dd8i����`�����iV;�P#sǔ0���3Z�[��{&l�+����L��'���q�ӟ�Eލ!J�	 v��6'l1K%� ����� "�m�u���0=ْ�>9P��e�;}H��ˈ�m��-�:�~B"�ZN���<�_w��'P֔�a��Zt8����&n"ԅ�I3w�ꁰ����Jb��b�I^`�P$��Oɜ2���Ƽ� �e�Ɯ?��U�}�V�;Ĺ1��OM��"�j�$
.�%�VJ
S�'F����A�\��@�U�$^JHc�'I(qA�Q�^P�"�$ވ▼i*����:OV����;\�QঊOJ*|�����RAł��o"W��hfkD��R$H�iy!p���&6FŻ��B/��� �QE|�X��|��>2L�<0�FҠu�m���')0�!Ǭ�#3�$�����HR�E�h�����*QY<fmµB�5J�y�"Acy�n���	�`)=�D1;��ϲ�0?Y�oI"6.�)�П>��-�j�DT�`�'��'[�A���P� e�V���Hx'�<,}�x�E׿�"�Z��D��7R����/��4p��5"��%r�]>E�j�{�O0+&� �u�M�K>��,\���ɣ O7O��b��x��s�M�Wc�����Q�j��ɞZ+H5qŜ��(QA����yn&�=d�LI���7D�Z��d ��ՒІ�8�tX�!I�y�ay2�;�H��B� ���r�l���{RX��F㳟���ߝY<�'���O ԠDKʫ��auʊ�$�-K�Pm���z�E[��yZch�8��L"^V=z֩��i@<5���Ǩw����h4�5��CS�yhr���o���RE�>E(j�@ A�
Ju�-�m�V�Q��OP�8@��12���K�۪I�� !���w��hHc �)��X�Q�i��'�N����d��u`��5M��QL<�v�D� lFX�t�~�����h�ZD�'���Kѯ`Ӳ�)�!�QV8sG��;��4��:O�%��W�$4�Xя��~�@�M(P~�o�U����Q
�ox����F�E�踸1+�H�裗�˙�MC1�ߟ$���;9|"Y{7��
T��suk�O�N�Vk���On�x
�+:�<��vC�2�ԇ퉥�~�y�O�5��/�b��"�8D�X]c K1X��)��$���r�Aش+��a+#�%V���ONXʓ�ތI�/V]- l@��^�VKRD�?)RjH�l�I	����t�4nPf���j��4�\ջu�܊bZdcr�̎F��8C7�E]؞ @��)ה)7�J8U��c�!+LO���p-��AEҰ���O�a`���>B�����U>���"O@l3L޽s��m�`� z"O>5��Þa��E���T3BX�tP�"O
Y�I�,:��5�6�� h�5��"O�i	dΌ�eړ���^��͓�"O 5h���M����ƍ,� "O����N'%��1�����⁛�"O ���� �T���"у�)�P! 0"O�53�J�~H>���"0h��=*"O8�Bc�˳���H"�ț@�d�ç"OP�#
��.:�K��2r8�"O�@��;jA!0֍��h���"Oؑxr�߇\h&)��L�@��%"Ot,�׆X�_�Xh��.
'o�PГ"O��Q�ʄMa��mۑ2/<
"O����]�[����Y<a&��"O���'E����l�>����'"O % � ¾ bx3��ū�Ĩ"O*���ƎD���*�T����"O�T�cMDF���p ���
�*O�	���\&���o��&8�'e�X��M[�J��R��2�P��'֨1(���>=�D)RM&�����'R
�s�Y:ڶ�H�!E�@z�'�T��$�X�!;�j�ʎzhqS�'+�I#��+��ڵx6����'~���2GY/o4�k`%�t�"��'�w%�-N��wȜ�_�<m��'l^	�*K�85Nd:G�N�Q'&hK�'=���T��Y`8��A݂X��ɡ�'\$`�g��JX&)v���@��t��vD
b�H8n��h�w%�#{$e��^h.��d��ܤ��6ݤ4�ȓ-��1r�EI��Q�@U~�d��ȓH�p�"�Vo�"���?�f���.��'@����a�	E�/� ��( yCEQ�Vj`CV=r��ȓ[м��s���Al��2�C7>�\�ȓT� [�*�n,��{�#�wT��ȓx�2�I�`T�3"�كG�>?n��t4��`�BG�$�$M�7�Յ��q@Oa����UJ6s�L�ȓ9S2Dc�
ٰ*"���'ڴ]gx͇ȓ\u}2U)�&1"��PC�~2&m��wfx�{�.Pj�K��سW��܅�v�����f��#7�T�e!���ȓ^���["�❒£��y�ȓX�q��O�#F� ���M/P!Tx�ȓ7j�bb�DvY�dZ�K(r[ �ȓd]u��m�Vm�3K
�6��Յ�JN:iR'����*xb/D}@9�ȓTXd����N9&`J���!W��D�ȓA��<c�MQ�d>`E�a���U����P�j�pJ4IpV���J "���q��[�O e����^�t���S�? �u3�ϵ^�t=؆$Τp¨cC"OJY3q���5��̓��ӗ|�sd"Ob�����k�r$C���4/�.��"Oؑ�N!RL	j#KU���i)"O���4�<��ء�5  "Of9�W�6�������4\F@�I3"O�d+�_�F�ll���HO@����"O�P�$m=,�HP�W�	�� �"O�(�w�M$�3Bc��
��s
�'*`�%i�	$z���M;eq��r�'w,��gK�d�l|ipN�a��( �'���Q%I��lI�ݠ'S�~�
�'�tx�櫍'N�@F̪I�M�	�'ì��Q��CӾ��h ,u���' p��"�]��U��F�A�Ɉ�'fɰ�H�3qx��EƊ:B&8[	�'�j����hkxu� fťi��X��'^�0��D�+�4BЀ+ylZ�'O�Qp���]#z@8�m�k:�͉�'�����:��@2�$\~���'YlT��l�-D��堖��^�#�'F~�+���x�$��E-U���'
��ڴ=�N�P����V� ���'�(0�amg��S��N�2(�'�[�L�O�)sD�5Jb� ��',�yǡ�$8J�d��fɨr��a��'P�-�Vc 1&�r�ځ��c�p�(�'����U
�=6���^�\$�'�`�E���ဤ�kRPk���'n&PƧ�51/��0 /��K��p��'�&$ǊʫE���(����Fc,b�'v(�z�h�]�B�@PJ^�E�L�X
�'��MɄ%��Uw��B��[1E�e8
�'�`MP o�8!�$��6Rި�'ز�I���?0X��E�|xB\�'BxRA��kv� �G
�n�|D*�'�� ���&т�
F��4l�ta�'�V�!�����\@�D�S0U	
�'�����X�j�0lۡ(ȌuǊ��
�'��ͫ�\�1v�	�l�{@��Q
�'�� ��
ͺYn@�d���p@@13�'A95�I��Nժ�aCW�����'�d�"��H =��'WO�d��'d��Y��C�i �r#Ɖ<�@@i�'~��B 
X2c>Eq򭂬]�Fak�'�ą��	J� � �[Rɚ0Q@J���'���v*R�T������As�$)r�'��YU�� �*xb6�_�x#Z C�'V��J̤S�����b� �)i�<!�.
V�`�cN�+@q��TBb�<��_�AS�p�7��&@���V�E�<���®+��0�4,�K�hD�A�<�Rd���(�cc�9}�fX�gF�<Y1	�r{:���=s��SaL{�<y4�Z�4����􏔶/E"@f�m�<Q��s,K�bR�}R8��m�<y�#�_�Ҍ�V�s�N��RGMc�<�sCA:�b��ehV
����W�<Y�����HQ�tE�P��3s� ��hO1�$�*[,8�6}k�!�!�V`�"O�x� �*�,�3fˣBl�\���_x��iAB�*P\ �R�˃Q6p�@�.-D�$K��ձ�ּ 2�U)kj����0D��3�F���-h��k�`�XA�,D�� ��kv�h4�CgG0N�h)�"O�1���z�H��EkL'R����"O�ի�f�4r��M;�)ܲ&q`-A%"O����+��eP�0����7i�+4"O�p���w�������=��"Oj�Xu$G�bI� J��V�kE����"OT��b�߉�x̓ JܳYD�p�"O�@�T�95Ҭ0����8?Z��#"Ov���W�7���TGU�	���"O�Yj�CK�� ��E�,��R�"O���!�1*��X!�j�'%y���"OHx!�B�!sr��j�'AA��j`"O�<b*P&�t��s'ĩκ�97"O�0ہ��-/�k�Z�`��@˳"OQP��[<l]��!$G�M߲�"Oڨw�@�BP�ȶ�!f�v�d"O�iaF��GB����Ӫ{�̄��"OH(	�� �v\Z�tdU��`�5"O���s��,Ŋy��c	���Ps"O:���዇+� �Ⅽ3(hi  "O ����jT�< ��!]?�L�e"O���@"�rU*�E�[�b4p@"O����+�n���"�+�*|Lcr"O��O)j�\�+:Q�BA�"O��Z��н��=�꒳y��aP"Od�f��w�����	)vl� "O�� tL��E�r�A�iTp��"OX��Bj�6QWX��F���fS��!�"O${2J�#k@&X�58�� �"O���4�C���0�I�|�dK-D���l�� �
��N���"e��� D��[e#�6�M�bXc�l��"D�Tx!��r�H��H�Uf�T��$?D�9d�N7M}F��쓓�F�k��<D��H�dmxt�䩏{ZZY��6D��k���.��ph�o���a$3D���k?�he�Pŋ����#�>D��a�$�z���(�"!4��*�k(D�d9���D��1���x>R��sL#D���
�e[���׬�7��@�%!D�H����
$�
AJ�	�>;��90"3D�y! �	q��U3v��qd�0D���ŭ&a�P\�&G	,ʞt���.D�؃ �����0�ȕ$#�ܐ�i.D�${�oŲp�ּ�g$�K2�0���*D��d���\9�d@� .ghH.$D�h�pA��E@�ʔ)��}�`�#D�49��'T���"��
%TY�!!D�8 �!%$5\��D�ɑTLR��&O D��'�>ExrMM�	^X@q��?D�t�Vh�����	�y��I>D��ڷbI�^vb����.g<�lsQ=D��3$��=33@�Yf�
���$� k:D��FO	��P�� �r�ɑFc,D���QA�,"�ֵc�f��m��a7 D��r�,�O�(�a$T�(��#D�$���7[� AGA~� �� D�(b�͟G1I�g��'�*-���;D��Ѐh\;Z�A����႑�$D�x���?� ����\�`���!D�d��l6~A�@�Y�lF�x	�f,D�<RVHra��W�A���񧈊3��B�Ig 2dH��U7X󲅲B��J�B䉑T��vI@5l�DTJ5g��)�pB�)� N5K&�
$�Ref`�O�	�3"O�� �'4�9����T2�A2�"O8-�ƪG��(��8S�t)�"O�I���^�tQB�a��:t���`"O�� ī]4I��%+���WD��ju"O4�A�$K�i�Z�*P �>d-lL["O:�	����Jr��ɉ�-���j�"O�M�UA�uL���F=rٸͱ"O��:GN�T⧬�>S1V���"Of!IA��D����6N�ە"Orl����v�x�YRd(d`�#"O"�@&0K�C��/O�(#�"O��aj�,�:=X�&بGE�U8w"Ox��w�X�f��ٱ��s�&XpE"O@J�*5{>n@�^8^�zJ�"O���SJr�l� �S�7��̡u"O"(�|< �Zt�R�{� �Q$L�@�<��G�ObJ�� �.i�)1i�z�<9��4t��9�M#�a�.F[�<�֧_�Z}�zFf�5(�r���KXK�<��gH~�����s��H��Ip�<�gk�+w�4�t+�ADDxiQ�[u�<��� )1�9ɦ�fO8��t�<��B��tQ�WeV1\\�u�䊆k�<�Ҥ��?⪈�SLշM����	R�<�'��2;C.l`T�5k���#`�O�<� e�r<�2���	���WH�<��נ_
ܴ�#�B2�(��%�m�<I��V<iђ�a�Y-?�l�Z��j�<a��ؙw�����ʀ'�$�E$c�<1D�E�m8�Q�'�f-`Ѩ�%IW�<�U	�,;�B�CG��2���Vm�O�<y�Y�y�,�ZC앚8}8���P�<1D�5�8��¤��O|��!t��M�<�6f�V,$����q T����H�<�1 L�Ph���ժiW�Ĳw!D�<���-h�b�!��S�6VTԻ��}�<�Ӆ)3�D�IT�X 8��v�o�<Y�=5�bY�aƲq������XC�<)�� M�Iy��;�(4҃���<�ïE6���FC�03�=����~�<��I&�� �)�)7���s�(�O�<��(�O���q����N]{�OO�<Y�:.T���v�[
`�ڵ��Uc�<1�o�%�t��D�p� SE��J�<qݞ+x� �1/��Fkt��CAC�<)�aR����i,-�yRs-V�<�Um.	��	��\)���+�N�N�<���ҍ{�>��йj�p�K��C�<��!@��4mR0n]�FfXY�D*VS�<a iD+��K 6j����a[M�<a�O�%�\��n,C	�L)Q��F�<�g/{��"�OH3#�ꏴ�y҉�$�;�F��,�^�+�"O�W%�,�y���£&��x¥"O81hP!I�"qk�.߮V-1�"OF!�aA_�i� ����	b��A"O6��2�ؖ(d�em��ܑ�"O-��HB�`T����#s:���"O�,�#r�d��)F��$���"O��
���y}���5n ~����"Ov���]�/,��$�B�yh�d��"O�p�ńҘ\N��VjƎ:[����"O�;����&Y�-�a�DWR0S"O� "�&A22�P�A�N�J�"O�� ��7$��SGK��8�'}�\c3L\�[;�����I��Q�'��H�o�s�豳W%�QTJ(q	�'L�����V���*G��K�.�Z	�'�B���O��r��"���{ͨ`��'U2Q0E�v�8�*#lF	1��x�'�nq�	8X^6L�'W��I�'������)����)�T�&I{�'�̀�aJB�Zp�/��Ζ=��'�6 ��"փ$/@i�1cآ=#���'J�q"�D&WQ䩋�׹h�X��'�nH��#��=+�0ɸ	��'�`\
�"Ҁٴ�;0͗(��E�
�'���R ���H,P�."��(�'���Ȕ��8���'"��}��'�x�;r.�7i�1��e��l%�	�'<�лC��Vi�e�:7����'%X9X��ܺh�������`&qp�'ў"~�����*��Eɳh46��(��{?�'.ެ��!݋ ��a���@����d*�>��1+�~��f��p2`l1�"O���w!?
�[-
�KVU�5O���-��!�"����@ O�|u!�ė�G�^tyb�l�&��r�Uh!�D��L�z�j=X¬D��mףC!�̈́r�Da��ץ&��=��.
V֛F�)��!��f�0C�-*��$m��Ų��7D��C`�*��r�I7Ѹa��:D�8J�(B�k�x�Y��G�	����`�O��'|��y��u���A0@:S�*H�<AX�	F��y2fʚu̺��I�T�T�h� ���M��'����ֆw�� RDeV	Z�:ě�'Ȍ�a���y����F�L�PC΍i�'XX�Pi�< k&�)7��0�'%�躃���<
v��to
�PLB�	�C�%"�OK�A�X�f�Tq>B�I��qr�
�-S`��9u�TY��C�I�G8���.�nٴ�:f��w� C�	+��R�oK�3��0;��Q�D�6C�Iu�R� �,�8d�zX��e��^C�I�.��(�����\;��S�S�����!��ͦ�DL'n��9���!;x"	�I;D��S�X VR�3��i�"���
8D���P�E�W���`�,~1��j�`;D��"�ˀW�`4�0
� 4��"�:D��
�bS�F�N�q�M r�jpX�b8D�X��/m�~H�� Z1+ iB�5D����� A��b��� �1D�����LMSb)�|)�b�2D�P+tI�? ���Ƀ[�8���+/D�X�� t z��b�ON��c�k"D���tNJy$t���A�	o��ɣ� ��0|z��&d�2�
�fۼS�ց!�og�<1��e�u��e���`�B�j�'��x2枯v��M[�C�y,rBG��1ў"~�_�����-N8)����0�\l,��':�}b!�6��ğ>9Ό������h��'%�P�jE84LD��嘨wt���'��T��*�TO��w#W<rQ&���'߮�k�U�6�L�:Ưڤ3a�@��'ob� ��3dq�U�bC3{����	�']j���Ӟr����r��y�|���'!4�T��+%T�(@�;m�Yb��� h�YtO���@eȤ�#҂�jV"O�:jP<Q���p�i�`9@"OV�4EP�r��S��/:����a"O����}"�hՊT�>���"ORh��L�<K�i��wS�M[�"O,))Qf�����USl|Q�"O*T	�h�rs�)s�!�|@8�s"O���� �I���OE�f@��"O,}�V*F[���
���;�)d"O��H`�ٲ|����K�+ ��0��'�ў"~2u�T�qj�#v��*X�>�`4g@��y�ە �`M�%h4����O$��D�ne��)D/�/�v��Ѝc�!��-,��3d\�l�ҌR��C1,�!��
����"�$R����"��+B!��4�r�襈�i�|�yt�F3,�{��
1VZXg͈e�@�k��3�OP���̻$�����'Фx.|)��Ŭf!�94�P)�B`E�<^xP8l�d!�$ɼĒ�C5F�I>�����W6W�yR�|2O@�񪃌�@�أ K�{
�X�"O��{À�ִP�N@�:'"O�%�&W�S��LJ䬍p�j���"O�)�3��<�5�F :&�AS�"O��3;V玈r7��>!~��p�	E�����b��Rf+�/Q�$�r�*�/�B�	C�U�AÏ�[+¹4�_5OeFB��!v��,aЃ��\���IU��2B�I�z�������.!²y�cAԐ!��C�	٘��Q	���R��[$B䉴]\N�1 獱�V��mF*�C䉗E��3�^�]z�)u�V�=ˀ��'ʓv�Q�$�@�>h��@`��E�̍�ȓW49���طk")�׉Ш����W�@a��ֵ C̭� �J.D�<����4y�� �0 f���*D�@�ц�3HG��c�&�:��$8>D�$�5�F"A�(�c'E˟ �U�V�7D��t�tj$I���J� �2t�7D�$�RW��9K��
�X����5D�����CϪ�j�!
'3Z H�d�4D�0Ƀ�)�r`��'ƀ5yڈ�(D�|)�i�:d�@i5�B�K�^MSD
(D�����˯z�ƭ�D��<u!mjAA+\O�c�<
b��e#┊��7j��r�J*D�й���7�"�+���=��4�)D��cb��)cWNa�Ӣ�*E�����(D���#j��+�Θ`���;�l��ք%D���E��d@,:D$�>�� �.D�\rTX+"��@z���D�<�L��`�����:A�F�K�O8��'��D�A$+P�E���&��ȷ�8D����V4���El�;x06�+�A,D���.%L8=�d[6cW�)v!)D��Zt�ѓ	o$��HF&Nr�d��%D��#1��//FA���G2z^6�[�n$D�|��$ق ��|��i�)�>\Cqa���	ix���4"�<����v�C:*����"�O&�OL`bVK3R�<Δo"*ai"O�;�JK����Y; �y�E"O���c��������	(
R��"O$�H�F�	��!6Dư
�n�`"O�Y���
�gx(zwB����8�"O޸�u�=c`����HX Z"O� �`��5=r
Y)T��h����"O�ܓ�*Ҩ	��0��=2���[r"Op8�2�xې����_22���"O��	�bQ�q�1�u.�$Aֆ5��"Ox�q��/�<��vm�8&,	�"O��Bы@�q�E3vK�?w�(�)�"O�hC�SR��+�RdF���"Ob�"
:f�+ �O�B]�#���yB�)u4��C�D��P���ybE�Ĉ��LSO�b�	�Á��yR�Y�DXI�mܖx㤱ʂ*8�y�CX�e�5�Amɶo��@y��E%�yB�ȳ"3�6�[�ZhD�`TJ�yR�9����¥^�PC���r���yR�:Ҽ	ڇ�J	��3�y��:h�`X��ȂFp�q����y�����^�1a�M'�F�݄�yª�6!Nv-8s�8|��=�@�Y��J����(���˄a ���i�ȓJh��䄄%���V����|��m#@X�7F�+ v	5*�6[�F��ȓۊ�a�f^����`W�2JV���ȓ"�v}���%�D���`�6�vՆ�}�Fx��10�ڵ�%Z+N=R���}�L��I��	��}�lX�Z��1��8~t:�BX��%�!C�$!Ӽ��d�Z�R��u_����9Z���qu����O6j���Ə��G:�x�ȓ	�v��B�/
���n��R�z1�ȓ~�0Y���(�Lz�P���ل��~}�5HI;������V#\�Ȅȓ7|2��c�RX�0H��B�I��[D ���,ei�� 	�'���ȓT�bd�Pө\dҐ{���su|��[��3�ͼ2��Sn��3�����v�6��c%O�^����HE$�hI�ȓi+|DYw�U9"W��1E��/$���]�48�k���r7N�^#
�'�~���wy�q�!�ݖ�Q
�'�8�BNДL��(y������}0	�'�&PP��� �d�Hm��"4EP�'s�Y�G�jt���r�5G����'<�Y�r����0��8,N�'���U�z�`��f�/7 ��
�'�^h;�m13�=�"ʟv�J<h�'q~�2�4x���4˟�
:�2�'<��`B�4Q@t���;�t��	�'�.0q��K[YRBɅjiH�B�'��@�U�/�;!�(�0W)�8I~C�r�N�*�'�C"�Ti�NѨ:B�I"Z��̑qfN���H�DR�X�C�I�� ��2��z�(�Á�+d��C�	
�f1��/����N���C�	������"ԯ;0��J�D��x��C��8t�T鋶���a�6���$�3e�W�n�x�+à7i+�E�ȓ�t	�*�J��p��
|����ȓ=-�����W�Hq��(B9��i���X��%a�Dؔ%b��$�D��ȓN �9HFi�A���y�Q�sߌh�ȓ>�䕲1�0� |��У�:�ȓEbpy鏟f����Mt�e�ȓ[@�p#`�cj�` ���7=ؤ��+ob�3���v[p�33�}�@ȇ�S�? � �B�߱ �p��DHH:�d��"Od9�tD>�����?I��
w"OL��$��H
�9آ�٧.��ѣ�"OF��wmCG���Y���ེG"O�삠���rZ�QK������U"Of��˔��a"���q�"O6�J5�:߬��*�=%����"O�(EG�>�J	���8_,�k"OVU�Ԁ����0��kg`A�"O�y�Dd�Z�q���]_� +�"O�9��&����M�8�< ���{�<Y&�;�hak�ߡ#�ej3�w�<9�b� �"�)^���#B��s�<���5*��)%�D'+�rDR�b�i�<���&+:Y�Ȏ%Y+^!r��\e�<9T�_=�l�c5����K�<�c��M���z�)ҟT��D�L_�<�'�W>i7�İ�dɓg`��G`�<�����pEdM[�lR&'48�)A�`�<��*F+n�*(�v�ƺH�����F�<���oh��v�Ҵr�P���ay�<��b�(�-�q`ë#0$����s�<i�ω	H��gI��6I(m�f��q�<� �����#bJ�OL��o�<!E	|�&13��3Ia"����Zk�<�&OA)g�r]��%^7
�<"�COk�<��W9Y���ԧ�tT�r��b�<Q4��4@+}�T4�v�I�<��톗����٨T����]H�<���^�օR�V�L,�`�KA�<)�	º|���Z�Ś4.���o�w�<Q2O7X����*KR����[J�<q��*@��}Є�ܵ84�y�1��B�<�N߿0OR ���m�y8SA�<��L�o�T�C� *{��M�d(}�<Q�\"#��BGf��I�\U��d�<��a_|n�$�f��|KH�[���h�<q�&� �$'*L�G�0B� h�<����-$|y&�1$��<p��Mm�<���~�N�A��N����҈�h�<�A��G7ʡs�/V�DUr8�oP�<	��L�uh�43��S*�"�*��Cr�<���пWH�I$��;H����lMr�<	���c�D�K�a	j���9"�v�<��)P/r��a���D��
i8���{�< %�!\�:��w��Fn�2�ABa�<iB)��n.�h*�h�.VJ�$3��R�<��j_�W�v�P�,�j�[�!�U�<90N�
��M��H:B��1uG�z�<Q�/�@ˤjO�Z���i�u�<a�n��"��G�����rF�s�<R�W�a=n� ���<��r���m�<i�GY�%_R$��C�aP��x��Rm�<��$50d؁+��P#V=� �g�<)#�͌�����/w��)&��b�<aՍ!'|�;�.��M��#�\x�<���-\�$(��<Cb>�#"��H�<��T�r�$M��GH�Q����PC�<ɂ�J�#d���ѡL�&����~�<�V�/*VQ���%�QQ�-<D�8��+[3�0��m�	�F�	�!9D���E(��&�@��f�<^h2O4D���h�
j���4lJ��(�)�VC�d��Ұ�G���ڢ���NC�)� (�y$C�A���xf��>[J��˖"O>���!�`�Y B�c�l�0"O����	�i��`�N[��rXjR"O��"� X�z�Z�pfǏ�4)�k�"O04�6��x9�)1�&}�Mh�"O|����@�z06d�d�@$�p"O�
�.�a����d�	�$�:H�"O\Y��F
s�M���G<��Q�"Ol�[s�D�fRV�CT�uaV�+3"O`�1@I�F35tA��SbP|y�"OȲ���]xι�@�$��%y�"O4�� �#wWb ��oiߐd!�"O��񀊁4x(Z	��r���"O��#x��)�""V$g��"O�� Q�ƅ�4-܈�"O:��ǀ�p�$��l*�j"O�|��fT�o7Z��!-ϼp�H#w"O��w���Y~N���@�[h$�"O�L���1��1��o<8�"O�E[�.mܰ��D��1����"O�̡�KυIr�8�GZh�VՑ�"Od!�7��(P�8p �[�t�H�"O�i��Ę;=	�)B�/�6�X��"O��c2m�6�r���,�s/�H�"O�Ѡʈ�n0�@T&��t��"O�mh�'S��EKP�Y-e��(�"O(�k¦T���"2C^\�Z�B�"O(|�$IM�� ���q��]�"ObEk�������4����`"Ot�V/:X,� Q�y�``r�"O|-acW�khl�%J �zpI��"O`ur ��1e4$����t@��"O�9A��-~�l
s)߫gn2� R"Oֹ�1�;C�C��B�lBHD�r"O\-c�-8KHɦ���6�<A�F"OJ�@��D���a���1o ��"O�a���#�6�3��rS
D��"O:ck5~�~���"ג
8�<8�"O�����r:��Z��˕��i�"O@b��޸K��i�����y�"O���n+IR̨c�H�t�����"O��ⰦF/�(}����V��hy�"Ol�������-ڑ���ns����"OrqQ�A2v<)i�L�.jX
�3g"O����ʟ�%�>�:t��x[h���"O���(�z�ڭ�eɅ�K��"O��鰥ܢ&�|��	�'c<B�x�"O���@�TI"��g�"��"O�ʴϊ�0�L��A�D�ڱ
�"O�#G�]"F7ze��<v���XW"OB|{�Ń"2�����eU� �$q�5"Ol���hU|��u�GcД@tek"OX7	�*��7#�3YR�r "O���i��b�EÌ�oڎ���"O���w�P�E�tl2��I"2��z�"O�+�c��E�A4��N����"O~�DE���VIB�M� vf9��"O��X`#�'(�"`p��ԫPl�Xd"OT8�ckT �ZcF�	?_���p"O>�R������u�PO��}t^��b"O�����'E����L�Gc�$"O&�8s�#D���K�v��T�g"O��*S�Q-H��p#�Z�I�Bl �"O��Z "ڊ(����#˲^հ��"O� ��j'�Ӟ'�a��P
Ҍ�r"O`��O�9KF��r�BϤ5Ѩ���"O�����$>�I�@����sA"O^����R�2O�{6B��"Ot`�e�E�}��`a�c��
xPB"O@�qc��h�#[�_<�C"O40q��%':iá��:�.�pE"O�MhR1,��Q�H(��1�"O�`��O�E��RHp�đÇ"OpPY&u� ���Ě�EL�9��"O�Ҵ��"�z#.��W2��r"O�A�J�Rs�@ �'ɻBм"Or�h�/���:�ZA���V��i�"OD�ҵ��,{v2�R2���l�*��1"O:h��ŉ��5j(�jKF�sC"O�Y05'F66���fL�0لX�"O�����T$�q+�ji�v883"O$<;W��P�8rbgʩP�F}�P"O�D�T`^a.L)I2G&���d"O�E�b4���藈A�&����"O��F����4�F�_�<�˖"O��j����Ry�E�R0D�v@ad"O����S�P�#�-�]9&1��"OJ���E�+0b�	V�ȔD��R"Oд[eΈ/^��S�A��}v��A"OR` �k�DK`0!P`K�[E�|"t"O�l��o[� lp5&�.�	RB"OVDK�.ѝpz�<;aĊ�n�E� "O��(<4l�0���a���Q"O.uH0! 	+�f�P�#Ш~C���"O(yrЃ�
~H��ȇZ�J]��Z�"O<�K���dQ��K�AB"O��:���7�XYPAӃw��8��"O�Łq���K�`�R�	�u�Μ�"O9[��S �4�w�Ɠ|��Ar "O�*P��?{�U!�S#bbs"O�0��̑�&d2'��%��,)�"Olź�D�>��LcgŞ"L�����"O�K',qI�@iЁ;��-;�"O���&���bvvP�� 9[�9��"OԹ��|(t��.z��U"Oд`K��b�0'�փd���b�"O<���Dҡ<ڬ�s3�LQq��hQ"O����K^D��a���zED�:�"OL�CKU�~c��a���"��"O ��q$ԷMD���w�\(M��|��"O�'%N`t��d+_�^��ف"O�l ����:��(*#���8��C�"O�i0B ��,ٚ�����@"OXi���!Z�N��]�Xɬ�b"OdA/m�f����`M��C�yB��%I�*�a�W�Uy4����M��yB���>shLʀ�ՅS����aa��yR�!"HU*��A�Q�9����y2
�̪��D�#a| ��f�@(�y�N� �(���fW�'�,������yY,�*��#H�t��i�"Ç�y����
,��#dI.oW6�y��J��yR�A�^Ɉ�[V�,g��Xj� ��y�tg�5�D�;Y��T�7aҨ�yIE`��R�a1^X�%�7���yr�T�&!�E�O)*��:�d���y2H� l0�S���  4Ҝ�V���y����G��;���r��AFK.�y
� PppU�X�IR�z�L/6Հ���"Ot,a���01��0�)w�$��"O�J%�2\�|�Qp]�[V�p �"O* s�.����YpDT�"O��C���P�HTˋ$0���k"O��3�jS�d$��R�P,%��"Ob��1i'8�A��ɔ�j$��"O^��3��,A��H��Թ]vZ)�g"O ��&�ɳz��\���\�:^� �"O �P6,�2]f�H��K@Z�1�A"O�e����LA�a�6�HPq� J�"OD��j9#�h(��Ҭk��"O`�ꗢ r�X��$��.[�Xp0"O����j_	:�����L' �P�"O2<H3��~���Q�j�~�ʹ�2"O���oʼT��1Ã
�.��e�"O�e���
�Ѩ	�c����b"OJ��+�K�]�pƍ�PGJ���"O��:EB�*&�*0B�囗'E�{�"O =�R
-B*QER�F�X k6"O���4�� �ܵ)�$K3�Չv"OHH ���@�D����:j� �zc"O����E����FDz�TK�"O��� �>��Tj!Ǝ7�` �`"O~�z ���2 �ɇ��D�h!�C"O"�����b��($�VA*x��0"O�`�B�; �R�r�,˸x$����"O@�ë/W�]�!�� )��"O�����R�#�&���
i�= '"O�	*g �L�T(��+d�.��F"O�$�֧��I!@� �H(*���*�"O�p�Wx���.w3Z�B�"O�AŠ�#��a����$΁ "OD�S쒕E�޽� h�-Lr "O`�:"�ˬӄE;�$W%(]I	�')�1Z�mԷIͰPq�P���:�'�`�H�e�	%J�耇�,
��P�'���։�#(�0����B!F��'͎��a�kc�a���I�q��\m����n=��4�aă����ȓ:c<C�`�7oȡ9�HB�8��ȓ�VTQU�
����Q��y���ޔ����tћ��X�7_���2�}2 H�p��Y��jH=1X��ȓ7iL�s�XS,�¶	;.Tp��%��.�$Y��T�`i^!��f^f�<!T%����мvI����F�<)e��oBlP���x�B�*AG�F�<�C�Ӆ)q�Q��ǃ�=��k[�<���^"/`����f��C�9�.p��hO1�&�k��$g,�cԷP4Y�M�!��,T��a��jX�������u�!�$Z�qjI��N��n
�c!� 0�!�dY�apVA�6D�51GaV��!�$Ҩ�t��kI�9�:��/N
�!�D�-�����@�K�px�eN ^�!�$ߠE`lhR3��Z��P���[G�!�
	K�ܐ�oͤM-ԅ! J���!���6bB����?08T�0˅#kl!�H?a ���H/���k�-P!�$��l���E��+is��T)!�d ��j�!&l�$��(�B�v�!���r�"d���)z�e�Vg�!���W�Ƶ*�dnE:0�3��o!�� �����aވӲD��_3j��!"O��3��zb���,��V��Y&"Oz2�m�.n}��zg��v�����"O�@��ݭ9�P�P��+$�i��"O�aSe�-.�5t�[�<ԉ�1"OB�ѭ׊I��3ƪ�)ȠRf"OHa��ϑ�1>�#��0@ 	I0��(D{���K�x���d�0��ÀD�1 !�$�f�L�ǖ� yR𦊗.i�!��P,���ԧ���y��*��9�!��^�H���J�x�P��rL]�!��n��x9��Y�-� ��s@>�!��+7�:yZ	�dT���rʔ�#�!�;�]�Rb�9A\�0���L]!��f��(X[.��(a�@4r!���&�2�
"��2>썢CEV}!�D�B����/�.z$��1e�aT!�D���ȳRʞ�K&h탢� O!�[�B�J|т�љ1ln=�_+[�!�˿]*��IԾV����f-�d�!���%�4XK��Z�Bx:��R�*�!���6p������*M;���u���!�  �2� �lC�G(�:��!=!�Iz!�\؆(&H&Y��|=!��4}r�4��j7(���	!� �6��;eM�6`&<1S��
>7�!�Y���1L��8B��+[��+�"O����A�1���7��S�:�Ş$���K2-�?z9vɰ�.�-gK�ȓv뾁�f퀙Wܨ����ܨ��ȓ`T��s�
�)�)8�Gޛm�¤�ȓU�-�d�ԣ"��ؠgM�X��͆ȓ6�R��'N�?��]�N�fY��r:,�cQ���'�Jp�$��⡇�xrT�GZl SBԝv�V��ȓ�p�����:6�|AH��יVn<���P�@a{C����a[�'\�s�t��SU,)B����+'Rpc7��3:���ȓD��`#D�4<�AD# ���,�	ᐎć'%���V��H��:;R��I>L��!�Ïz�ƥ��V�ᨇ%��x��%�
D�D)�ȓ�́S��D4r	Ӆ%�an� ���<��셠s.�����}�t��_rD���.u�@ĳ���~݄�I3�43V��=%.h��@��N�����v`�h�1���*T� �ȓn���À�_�u���Җ��m?2Єȓ\ex�gM�AJ��N�4JR	��[be���ިb�L� �4h_�<�ȓ��II&�ѐ��y �/�1.H@�ȓ{�=æ'٤Q��-VI+\t(���j��q�[2���	R�$���ȓ4Q��&T�U����ϒ3��х�`cA�Ed1:��·IC�)�ȓdOp��$���w鮑ʡc��%��ȓM���Є��7(�n-U`�/B�F��ȓZ��h"�����٠hX��B)��$���!��1�ԙ����RՅ�}���А��)U��%@��q�ҕ�ȓj2�S�J�?���E��=	�����7�����^ B�}��Aϡ^�>4��xo�ex�'PK�X��ҝ%�dͅȓx��u&��o���x���l�t��S�? �02A�� ���
����f"O�PU�Ʈ�5(�!�~�:�ye"O�TiP�;E��a��ʟ/f�N9��"O�8��%�<t��'��jJ�"Oܑ۰��3��9�g��KI,H�S"Ot���ǼEpܩ����f�"�a"OV-{�T�PppOȤ/By�4"O��R�@'�Za�gɻ+��`"O�L��g�t��9a��%�J�+!"O6��G�_�9��s���Ɓ
�"OmJ�H.KmN�2�W�;7H�"Ox-W�ʕ�I����A3(@v�<Aæ�8<ڢF�1�X��kWp�<�����l�%��-H^�(�sΙa�<���ճu�T���_-qt�`R�]�<ɷ�c=t�(���+O�����.KW�<ѵ���:P�y�%��/���!�BS�<�S�I4m�l�ǉ��G�d���f�e�<)�~���S�ކ�=A���^�<�#�G�<���ٗH:9�ĐZs��Y�<)�$ɥM����1��+&\@�2��\�<	
M�9f��H$xv�UK�t�<��i���(�������e$[s�<�'�ZU�<Ygk�^��U�Q��h�<���� \����O��(U��`�<�2��9L��7*N[e��P�RV�<���_r��-��PH6������x�<��-B4V�p����߅AF��1Ab@�<�dЁ(�XЇQ�:$����t�<�'��b.@[��7W�Lyi�FL�<9FE����b*Y�^�����m�B�<	u̎;ZP͠ㄳTGš)�U�<��Ld`}Ӡ�( >u��QO�<���' �!w`({@�"�H�<�T��(i��CK�$2��X�]G�<�#N�m�\���hK�D�q�U	KJ�<���ܮG:��t��3��@qRL�<��J==}�xq7���B�T����JF�<1F�A�#�4�BC�}��D[!J�h�<y`�R�\�zw�;�m���`�<���N�vd��ǰ8Z
 '�x�<���7#��iZ��F/4�����i�<���H ��{1d�.-o��1GI�j�<!`�V�*�6e�,�)qr�@�G��f�<�¢Jf^D,��F��a8U,Da�<������Q��<��A��Au�<i4 ʖn+Μ�,I57�"5H���s�<it��#3I�t��j�t���W�<11$WC�hq�i�.`����V�<!AHsB\M�H�8e�,@#M�U�<Ѥ@^)_�ؐS��'�U�H	\�<Y�b[1W�M��oTzPQ��T�<����:ds��h��K}�*�c��v�<p��:e�Tq��I9SP�A3e�r�<���\�o�"x��_���l�<�΁� �̛!�\�X��Q��nc�<9סV�"�ի��3����#Lb�<)f'lF�8�$ˊ��tS� �^�<9�� #@i>�4�u~���#]c�<�'�Ǌ/�ܲ���n� �E�h�<	��7��|y���>N�Q("#�a�<	�	P2Wg�ͩ�.�=Y�H����e�<Y!�\V9�@@�0B<���_�<aëA=o9x�1��!8>苔�d�<� nm���ӭf��͛��̀�L��"OLu ��M7.|�APĬܙd7:�	w"O�����ȂG��UikݦS#�!zt"OĢ��C"YZQ��6`Թ�"O|�
��f����L\#8б�"Ol��"՛#%�p�/LY����"O�a�4-O*��੤̓,[���"O�x�cѬ:ؼ���% �z!G"O�u��N�	��h�ս3��X:�"O:,�4#Zx���:2�J��R"O$�a%�HI�th�3%T��u"O�x�C�ReB����D��N���)"O����/_����8���rɱ�"O�t������I:�烧!��1ٰ"O85Ҵ��e�� �I3�-0`"OT�j@�Z X��6e���5CV"O��kLB|��ͺb�T-�L�@�"O"L�$��=X&\���Ùa0��5"O�l���[u�)�A�I

p�R"O^ �1��6oV��Fg]7=�xE�$"Otepf���צ�L�L�bS"O�Ńu�æ_�"0:V��`�=%"Or�qC��|��;ׄ�	>[ܽ�4"O�Q
�lOSF8 �$T�Ub�e"O��#"��>OZ8t��P�,_Z��"O��p6��
zD�������k2"O|�jt�Q>3Ȁ�[`�T=u�v��"O�y3iH�`lx�ɠ�]!$�d"O����R���s��g�(g"O|�Dc��Qi��Id���"O6 А���W�|d��m�*�ZP�'"O��R"�Wc��p!�f�/gWJ"Or�a���O��hH�D�wQ����"OzYo֦!j�=���̳9�0�K�"Oxä�H1&�2�����Ω�D"O���@��<a�8����9L�4�x�"OR�f����8B�������"Oq���`�걡ʔ�O�X�"O�$����,��\�e�9K��W"O��h�Ɍ�@�p`fB
{�$@(@"Oȡ�uϙJZH� ��'�`�W"O0PaP�W�l�t�4��.��A�"O������@�"Lh��1��"O���GW�G-�D(s�#�n�"O��	��V�Y���c"�Ԝv��1��"O��	���X�ݢ���k�4"O���%2H%(L񂅋"9����W"O��#֣�^ n��D�3֤""O��h4�ٵL��:en��]J�Ӡ"O�h�`��p`��aD�W�E��ӑ"Ob̻"���
G��5�H!w�,0K�"Ol����'%Z�KP��q�� B"O~�H���L�! <����e8O�=E�DÝ
�>`�@'B���ćĂ�y"���R?�|{4&Q�h����R�y(Ц!
j�� ��*������y��8HI�ca�	 Ir�4R�۫�y���.E�lF�m2Jh�B�,�yR�N~0��P�6�D�R����y�Ꮴ)wڼ�Ŏ(͜��q��#@vў"~Γ=�:')KĐ�H��O�6��ȓd�����S0���"�lUu������|�a@Dkw���cb ���K�E��ݫѠ��Ra,x��S�? >��6d�$z]�}��/��j�⡚�"OH�ɀ�ǫ�P-k1.�B�b�#"On]Bqu��yH�"U����?O�=E��lđjJ���'kQ$��hBE!�;�yr��7N0Z��\��*%i����yl�x0rc]�G��j�G�3�y҉\�:n�Ѓ;Q�j�=�yB��o9$A��д9H��:Q�H2�y� O���2�\0��%I��$�y�m�[�xm�r+X�-�7D�����'�ɧ���$�j �x#���IP4Q��Ȏ�9 !򄝸T@`�bdͫ
N69��(O"e!�϶o6�IX��F�O0 �siײ$N!��P���%�P�S	�,	�*P� �!�$�Y?�	Xt��j����P�M�@�!�$Q��ؓȇA8��	]�.�!�D0w�I��&P��ԉ�\�Ix���O��"~6Lې�&j$"�2�r�9h�u�<Q5e1���;1�M(2��E�I�<��ޔ� 1*rgԢM��$���k�<�Ӆَ���i-P�w*��pOFj�<I7���K԰}iu![(b�u��XZ�<�7)Q >|���㨓$5���R��^�<��MSq��$�چ}��/T,���hO?��K�=na��Qwˀ�T��]�,D�h��W+j����G�D�=ɒG,D�P�E����2�R*o���K)D���&͓*T��i�φ��UX��,D�L�JM�e��z6B w�bY!'�-D���g�>jS�;�Q��(I�Ů+D�dʣ,M�pBU�Sc[�:
�0�f�'�O��O�	i�#ʔ��`OPz�L�e"O���̕�u���s��Ǒ)sJX#�"O�Tҕ�� ��p2-]pK`�k�"O1f�
�/@&@c"/���۷"O��x��Ƨ�R )��$�� !7"O@�[U��l�`������ "O��)#���:����f�~FFH��"O\ ��ɾa�z�3��$FlEZ"O��X�)�j qpM����"O��;w�מa����Iû1��af"O8��􂐈m�4���E�>�}�"O~i�UpRXyDj� 48H��5"O�u�+�(X3u�A�+�e�"O&t��&�pcX�c��Zh�<(0�"Oh)�'T�1|䍪%א'?P��"O�92 ƻmXr`�%�u:l�H�"O�ĉ!�{f���E�%��U�r"O�ȹ��A�n�p�.Sx.�X"O�]�ulĆ*ߜ(���ߐKq�BU"O�����&o��k���kf��A"O8����;1i�A1�I.�t ��"O���E��6��eQ!��;m� aU"Oa�� "�ܣ@��8��2"O�HH7�@2Hؼ�%�%�R�8u"OHj��=*)Z<X2����t�ف"O��'F-� �Ғ1�Y�@"O6$@7��:w�%���CQ� "Ol}p7�O�zZ�ѴLX�dʴ���"O�L�Ɩ$�<I�E&nf���t"O�,�Pő0��{��X�5<�h�"O�	�R�N3�<eA��q-��r�"O���ᕾ3|�Pk#��'t��Lp"O�����s�eA���`�()�"O� X�#HL�='��xFDי;�ޥ*�"OT���$O F�x�5��6{�nL�"O.���(��J�~��!�I쒝��"O8��5�,��1E�A~�!�r"Ola��٣p�px�VS*wn�ۖ"O~�L�!:�d4���#dh�"O�x)�K$��5��N,WV�T;�"O��@�nM'h܉G.íj)LY�"OB�v/+ P��(s��V>��i�"O��Q�F'7�d�pg&\�.��Z"O�0a�*-%�,Q���:�K�"OUV�_3 vt,*�g�M�d���"O�PӃC��C�~��GD�<j�B  �"O,���.5�`�T-\%|� "Olq���Ru�ٓ%C�\j ��A"O��6���B���oDz�����"O����鉃��jb�^�)��ٵ"O�TyFM�+?P@�R	ܴf����"O l�'m˧<�Z�A���8Y�4�1!"O��(E/9(�M��3bF�ó"O�!/���ɱ1�˘E�|y�"O̹"p*E�B��3�j��t"O�ݰP�T#d��s�	Ps�2d@`"O��˒l�F�J�8'(����}K�"Of�
dN'W'PK�얲1m�iP"O|I7NN�:�Mx��@�FUL��1"O��ZV��	'*]�	N=r,�92�"O�1Vbݪe��Ƞ�^:o��T"O&�{6�� v�B-�Vg"0,�F"O�+�%͙�zH�3lY	$����"O*�����u� I�넹!��!"O2|�^�a�����.�1³"O$��eO�2�h�b�h�	N�P��"O��)�?"ʼ��q��]�&@��"Oި�4�Lj]fpY�a�?5�����"O�a���'`���-Z����"O�@�3`�,t��ɻ�,��/|�T("O�!�H
�D�DeA��ixT<�"Ǫ ���-~�`@���1���;4"O�"!-��M;
�
(Q�eh�"O&�c�*�(%C�K��Mj8�"O���N�o&��!���"?���A"O&P�Q�V����-��9F"Opk�-�"v�cb��t��"O`P�F�9nD\���*ãJwVH�d"O<ݪ"��ca�X�fL�,s_��k"OPm�S �=���� G�0V�\�"O��
��-?Yd�oJ�Y�PňD"Ody:�� ���ү[����"O�h��>E�.AJ��˫���9"O��0�ܢX����<�0�q"O��B�H�l����	�Č�C"Ot�sF�̢ �!-K@��B"O�-i�B�nejP�i� +�H��"O�XRO���~T@�5X�k`"O�q*�(¤���(%��PNި�"Obݘg�v⑪Ab+�V0�y��(l�0 2�B��?�D�զ��y��<x�S05�����˨�yr�D&&�"<��.�1b�@��T0�y�"�*)�-xG�7"N.)0�ą��y2F�1@�,p� ��q�FQ�y��8����%K�Xm!�O�*�y"	�� 1��V�JTR��ʚ��y
� b9�r/�b��A IK�g��͛G"O܉8v�&n%�h�>,��ؙ�"O u�ׯԨK�t8��ޓU��� 6"O\4!� �$'�t��Eޕ-иe��"O�1���	'�\��cT��
@H�"O�a�"!
�g�T��#��-J���"O�(�a�ޛj��}Q�'�X��@"O��8�FȚ*W��y��@;�d��"OR=Ȣ��1��]`ҁ\D�JIx�"O�!��'��91q��G\4 r"O.�"�[�Fj�& !#j�"O|��Ǎ�w���Ҳ��ag"O�aPנ :WKU�Ĝ��W��y���u�~ i2$�|�бRfjT�yR�:ʊ��ʖn!�v"+��O��3?I�GJ�4,��٩|�ֱ�6�Q��?��2�����*LD2u G5y�d��ȓ
d�ػ��Дc��t! �ʴ~��Ն�	�đ��n�>f��z#h��T����i6*U@��� N��:T�1r@$�ȓG¢����Q8a:Ι�g�̮.����MY�$�@åp��I��O�e�D�I>q,O1�1O��y��\mr����I�"%a5"O"��#ƛ�%.5���bcd�A"OB�q�噩L�h��j`�ZMy�"O�}ӲZ�c�h�S�]�s�>z�"O^��R�6N�$Q�k͞�2��F"O��7g^.� ��m�$��Q"O<t�f�?E��Ё��P� �@��6���Ot����C�K���)qM�M�8Lq
�V`��/�O�Q���@e�=���F),c��"O2![�=V���D�9'�1R"O\H�P=K�Z(AnƵD8���t"O �f��ܼ!�lټ%�Mi6"Ot��D�=_^8�+���{~�(�"O-��h�0q����5GN�B!ܰڥ"O�t�p�&13F%Qq��b6�hB"O���r�)yy��[4�%�����"O�4��c�Z�hD���I�
��,I�"Ox	�
A�T��m��M�d���"O���g�~-��p�.	�&Z�3D�P���X�����!�P��hʀ�0D����Ǎ����f��#a"�!�F<D���p��\$��NػL�&!CD�5D���͇�m�����G�ڭ�%b4D��`��U:Y��첀O��4U��0O1D��1���_�xP��eQ�);n��U "D��$�]�~����%�!\�Q�?D��F�@�i���z�F+D���6C��Yjg�Ћa. i 4D� 0���$/<�P�lʸx��
w�<D���q�	v��(�0��6C�r�<�6��"�[����[�Ё��l�<�R�	fh+�j����&:хȓ9�]	�%M-���y�R5(���ȓi{�MʕF����y��\�u�T�ȓ<t�H�����9�r�)�@�7.ZM�ȓ
^x�b��l�~���"_)�0Є�h�Pd(fl�-]\t	���L�l�ȓK(�P����nt��H���p,��$w���SB��2�nxq�Ó�6;�d��HP.���u @iq��#<z���{"�2�LA�Ϣ�0D6>w�Ɇȓ8�-P�Ρ,����$��%��S�? &A3�I��-N4h�앤>Z9�"Ot�����6�.��0�8?����e"OMrpfѺ��)�G�m��M��"O��"� A�O����J! �o$�y2.�^g�$ytǛ�u�,��RmI��y`��"0�",F&	�Må�O6�y�j�H	d(a *�7bE�%�O�y��
�o�6��$���Ku���y��O�}22gf��
*2��4AI�y�	�?��-1Q@�,n@��qoA��y��;^Ej��'��4��qA�+�y.F�G�@9����ckD���n���y��FѴ�ka�ԟle�!��yb���#�iSg�K���Y!b�V��y�'1�R��n�$n]���y@F�lh��)�� �9H ��yb�_�|j��a��|P���Lݞ�yrhI�V�:�Q6�_�%R��$�y����<�2<	SΙ�Q�P�i�(���y2�ҝ��@`.�#@�X��蓽�yǏP�Y���׃;�:��CƂ��yRźir�\لE	�/��mh���y�͢4�\l"pkLZҺa�p���y2��-DW��0eE�.Rf������y2J�g���5Q^h�0�T.�y��&l� ���cG	C�H���L�y"���Z����43���r����y��� B6�X $�T1�B�	�!�yb�G�cV���)��,�|�s�۠�y�c��14@��⏆7\:�S��yO�#=�r�ڑn�:9Ԛ�prG)�y�쐯�a!�ӑ�b��y".
��zu����2�*�O�y�~J�3��Eؤ��u��4�y�  3u����� �.B�']��y���yh�B���z�R1��y�+�"�4�@ϛ/;��l��T�yb�9,j퀆B�E�
��	�!�yҡO�t�w�Z�Tp.��DA��y"�Sb8�E!X$b�J@���A��y��σ1!}C��')����ޓ�y�EV+�Vp�C��o���V���y�fC�x�Ys�L�v	ti�˗��yrf�3�2�ɄĖ�g|b��[��y�M��28djR�M+\�T���X=�ybƁ�6!��1f�Wi<�@{4���y�F�\�g�-.vu��+���y�I�+�ě��A}�MZ�F�/�y��<4!��!�p��Փ����y�L��J��
cC�mR��(f��yυ�vv �3%E6gzؖ,lH1��9H�] ���.d��6�ۮ=�M��*�x��W�|�\dqŪbȄ8�ȓ9�.��t�}Y<I!�Kd�D�ȓ*5�`0��Y
	g��;��B[�`Ȅ�7+f�;���CZM+ba��+�����V,�s�ب18 t��Lܦ
�`�ȓA��)Q��
R�R��7�#pM
��|I�)Q$ p�ѫP�0�tQ�֪f�<���
�� =���d�T�d$W`�<���ô �9; a��#ϤőIu�<q��ˊB=���Ɉ.���a��s�<��)��<��Ձ�����	KV�<q�ޛYm 1yE��-���D�{�<� H4��.T�L������E���h�"O<P��������X�,���R"O"�Y�C�@+���h��y"OZ �2��6�ʴ�c�$R�$��"Oj婖#G�f�J�ݚKVn�h#"O8��2(4O+�`sq�� 6��Jq"OԘ�!ǖ8/iܙ��	W�Rq�*O��!��Q(��#�¡z� ���',�U	���#^;��H�'���
��*X��M��LӐ#�d��'�5�Fi�(!��G	���'n�9:E� gց���W5@���k	�'���$�H;�4Ys���?J�U��')&
��֮w=A�!�@vd���'2r}s!ЌBh���D����	�'S�刖�>tX���P�(k	�'��jp�M� $��`�7F�t2
�'a�1h�\� ���B�H33�D���'k����0H�<R2�ʫ*�D��'8(��U��3!�`�A�I�! ĸ�'"�P��n0��HȔ� dƀ5j�'�5y�����0�j��Q\�i@�'W�p�W���F}���x
��i
�'��p�!�
?�:xck�4q���	�'�X�pm�2�i�ǦL�iO����'sf�)���>L���A�a)~���'�8�dK8��L*M�����'c	�v��ULI�5 �H����'BT� i�:/sT�f��>@{0���'X
m�q�A'KW�+��I�;d�yY�'�8ثQ�v�,96�^�=4��r�'�x�1�	��tM�|e���a%>�#�'�5�Ҍ�;s�VB��Y��lh�
�'���4/_.P9�*g"�3v6,ѫ	�'��)�Jځg�Y� Y�s�t���'�,��1�O�5dP��b�v��
�'�^�DMWo;�����>J�8 �'L�p 檖�
Z�bUe^7@V�#
�'��[4�I'>l�G`�<%�)	�'�6������-z�� �4���	�'�ƅS�h�1󄸁�E5@(�c	�'����فF�ĢS��#+| ��'f��V��]�r�����"���'��m�`BS)9�����(E��|]��'���%nZbX� M
�N���'�zM)deB+u/J���B<V�4P�ȓ.N�j�l̕|C��9���:F֢=�ȓt�j�P��ۋ8"��4h�4���ȓ9�0�����n��i	�JC9c"L����Xݸ�a;��g㋱q�0��,�A�`���9�E."�$ԇ�&D��Y3D	�?�d��.H�H�*L�ȓ	SP0�B����h֡ȹpf ��ȓ��1i7,W�k3��yvN�Y�ą�5�:��,O$��8Ф��� ą�	In�Ӈ�T	�p��5m�:�i�ȓ(���q%$9���BBM�7"x�M�ȓF|T���k�D2Ҍ���PH�ȓz����M�]�⸲��O)4h�|��K��GIF�PT�@��.���ȓh���r�[,���A%��[FR�����6�A 0|�9��N7k����ȓB���{GM�}'T���Ѱ[b��@�RPQ�ЩO���hq@�-!��]��S�? ���c {F)S�!�F7Dh¡"OF�H��7%2ح��`�.-��s"OrUcd�̍)j��ӭ9:�X7"O���e�U�`�R�c�%�T"O�A��!\�zo|�B$  �>�I��"O2�+� @q$m�`H�Gw��c�"O��qg��j�,˵N�mc(�2"O���V	]�	d]��*�X`�6"O���A?�L����-F��p"O��i�c[V��crZQ�"Oj5�� !s,
E�`� ~��K%"O�ب�L-@�j՛4����"O�0��`�7i4��h�0��Qa�"O���1�
�T���' 2��@��"O
t�fۋS�Q��5VrP ��"O�PӃ�A@� a@
�!X��@R�"O�p���3*�����W�Z|�}��"Oj�)�ܖz������:%oT1�"OZ� 0. �6��9ل κP��y��"O.]���~��/M  J���S"O:E��/A$oǼ��7ϝ�!��{�"O�x�`�tټ��קۇ%� �t"OF�)�#�i�
���/9�"OD�FO�~��h��ƳyQ�}h�"O�Ӂ�ۼb�Ně�'J%6(�P9�"O�� Յŧ8U8}�񯌕b�|�H�"O�1�T�̔H��"��O�ɼQhU"OF	
��ƳtW~ J@Eȼ�B�*"O&�����5�*]P��ǑC��"O�qfn����aA�� ����"O� ��h�-[��5���������"O���)��04J,��Z+C�����"O@��P�y^�]Q�O`Ȟ5W"O֜@�ڇ$��q��Ѯ;�t���O:$Q���0>irF�(�\�����!w�cBNE�<�&�ǶP�HƓ(3\�:q�
{�<����8�	��>�ĝ�P y�'��?!xЀP{n881)G��y�P�9D�̡3�F(>QP��l�Z)��=�{��@�$��է �������yR$���d������x�B�5��>���*�S� X�]�*�,HD�aA�/I�4�C�	15���s�߿^����m�O���ēO,��.7U�"�a4\ˎ�#���Y�y�����a�O�3'����LՈ����
:>�g�i���$@�a���G�īb`|\Q�G\�'L�'��	ryR�Ӻ2(Nٺ���
�����Xy`B䉉y	�d�C�K{K���1@̠C2O�����2�R�E�T&�y�!�2�2�IW��	21<�3�Ǌ�y�/;>��"��$F5Y�m��'h�5����ݝoo�@��,u��{���=U����D�ğ\��M)EF��1�L5_����!*D� (�K �BP��F��UەA)D�$�!RW�@��E�3�%͈�<Q	�v3�cn]7�,A�֬7�p���I�4�O<�I�'���!%
�:.�(��TL�
f4B�I\)P}��*�1qh��A�K����Od�ɍ��	2`@U�D��8� �w�!�dQ�W��r���
l�?�t���d)<O$�
ҀVJj�Ird�0�$H'OT9s��
`����c�ȥ�1fJ�D
6#a{BhIܰ�S�S��ȡB� I���?��'� U:�eU�BNN	j��+t�+�y�ӓ,2����`��0�T��y
� �\x@DV"����%�(�`1�"OH�h�$2��yv%�S���W"Od�С(Z���$ϫ~ Mb�"OR�C�>ɮըf^Y*!i�"O��{�\�+oz����ƣ0�:@���'1��	�Vz�Y�gğ� lѫ'��"f&B�ɏg�`9 d܊!z���
�Y�2�?9��IS<�z�·�Y��Ϻ�!�$��������O�}�"EsE$���!��C��(pT���-��C��n!���O'�m��O��~(X�(�C
�|k�ġ�	!O��z�h��Z�\|g"؞D���O����s����#�>E4�D8P�z�\�	xx�hy6&j���D�!ת���8LO�d�>��aE�8�*��E�A$H&�]�a�Nt�<aA ՞J��೥ߜn��D��=��'7ў�OrN�����8+Q��ң!��K�>�C�'��yh�'g��H`6��1�,P��'㞔a�,WR��6j;��1��'���r�Őf���r ء�2i:�'m� ��X8q@����M��0��OZ`�d	c���E#N�d�!��	p���)Tw ��'��s��x�P酠f!���yd�4�&f����Ys�=F�!�䈩w�<��Å��4���D6�!�Ă=	������6-:FのIwa~�R��릎у�~᪕�ATf�#�N)D�`@7�T18���'�Ej�-�2j1D�[D�"ՔM2�՚ 9t)Rԯ/\O�b��23BM�T�(���g:�X�Sa�"�r���Og��J4��x5��-9z*�{��)�	��X�v�c���"4^�q 킗]��ְ>�7�A"� ���dD FM�!L3�hOQ>��8O�q�`L�ǺUG��q2T�
T�'���i��1&���.�|�HI0<r�q �'����e�CaV���^�.u2���Xt�����ɡ($ꄪ� '�����D=��=;��`���9��Ӂϒ2[�HB�IsՒ����ېg^B�;��ƕ�
"�(�Ot�֩�' �-���iw�A�q"O���VA�\�ZLx(�jn�!H��=4�����ðfM[S�M8- ��cF"��Pz�'I�>)Z,�7]M��R�ꖮ>�=0�� D�8�NXi�h�(�DӚ ��H�U�=�ߚ�(Oq�|x�B�p8h�gCߙ7W�a�"O:�;�'fnaƯ_�G���2���O����H$<��v��iT�=�Q�O���<��|ڌ}�ıL$��k��W�.H+�NU�<�DC�e��I�f��;ra$�� ^��'sa}�M��Tʈx"I�t����^��yB@�7�R�+�����|�` ���y�A
�w���	 ��(X���O�"
�'�~��=4�^�+��P����h�<9�,@�gHD�3%��6��*d	@?i��퓶fX����L�<a~m��.��l��B��,�=6�\5����,�2���'�a}B�FP�n\�#�i�j|C5�V��y��H/;r�tQ�NϒYk�P�F���yr R�:�rH(!�G�Sm��	!iգ��ODD'A��?�KVV:u1�d���H�vIR���)D���s!�3"�XM�T�H
y�4�a�D>�yr?OB4姈�ҢY�B��
�-V�GI
�5-�'�y��^�ؤ�� �B���Pe�TY���|"�'���O�`��lJXV"����S�? j<�5�Q88t��3� �*����D"Ob�T蚀(FZ<��F��+��:�	J������8�gL�+z���/
�!��J�R��M��rC �sTo�U�ў8�ቛt J99��uu��KC��*OX�C�	#3m��p�"^0�i��܅L�FC�I. ��0��+�/.���a'�G+���=�"t�Y�2I�,T�L�i�1Q
C��M��h��B1��@�w"
U�D�ܰ��)���	�N��d��!&_�d�DX�y�*�+|��i�ל#:������hO���d�0�Tpj��*�]ZТźV�!���I�P��4!Х8������9���u�ԅ��cx��
��]��:4����# ����K�<�I�ЀAD#	*D�X������K��$D�$�����}�v@�Yx8偦&7D��T]�'
U���@�ѐn?D�X���v��rş�T��#�<��<Y�I�jkj��u�:%�PX�n�z�<Qg(6~���sl�C�8|����wy� 3�O|�!a�3����	J�.]���'Z��-wO�D���P3q�d�0�8D��;�HZ&l����cc��B�h4D��aD���)t��5� n�a��/D��" �V�%	
���խ`��/"D�����(>t�c�f)~��wi=D��y!�5�1�T*]�x�r:D����̊jh����n�����6D�Tk���$ˊt��F'#�PY��6D��n�xXR��#š
�m"�(D�p`��@��)3�C�6�����$D��8GDEp�܃q)�N��E�-D���@��b�6`�tg� "�n(Q�m-D�h(#�4N�BF6hB�5"*D����+ZU��k�`� ##�&D��TLx��ib��v�J�b#D�Hs��'Ռ%���.*6#T�5D�<��eր.��5��. ^����1D�,���'k� ��K�2;6ZMH`/0D����+DF�` ����q����u,D��󠃈)_`N����K!
=4����?D���B�y�Y�C�k/l��O>D�|c1��HQN�	Af�3C6T2��/D��ˁ�N-Ru�ALU\2p:�d)D��� g�:L8H;# �	S���#�%D��Hb>b��XZ�	 L�Y"�l!D�0��	����[�Ę%Ee<D�$�����T�r	�'��'�\��a;D�ТӢ��x�! �T*T,^�x� 'D�S6�ӱV���iQc�8�(9��&(D��!�R�z	��N�
u -0U�(D���Pԟ>즅YW� 8:�܌��(4D���WI"�,)�B��~/D�D����r��:R┎MQVPj��/D�0���=�x����8�<Xi4�,D�������� ���yrb<��.7D�L���
8	�d�� G�2^8�B�4D���5`�)-X4��ԤÕ\Tx��4D�@q��Mm�N���*B�$�֍�"�3D����Q<S���2��@6Ϭ��qL0D�,e�;4�LC�K����up�&9D���Q��pʱaw灾R��M��e"D��C�����u#c��W(��Ǭ%D�DJӏ�3!q4`˓%�4d��=Y�#D�� ^��%�'^<�,hfC%�D W"O�E���"�Bi��Ԟ���	�"O~	�˒���5a�Be����"O$Q1��M;�R��
%eR��T"OP�pbM$T����DJczx��"O�1���<S�&8�C��/B^D�8T"Oգ�节n����a�?	Uv�qq"O��c �#QĽ���]�x`L=`"Oԫ3��@tc�D� F���!"Op`#����͊g��j�`|!w"O��(D�
2��0z4E�2a1���"O`�9G�{ ԁ$��`Lh�"O�1� �H
z�؇C�+S�r�"Ohe���RI���M'}��"O�1!�~� �G��'�.�"O����^�	²y	deNc���u"O�,�v�N�ȋ���T�LS�"O�;���7$"�"$�L��q�"OV���k��;�l�������� "O^\���8[�JL�MCڀ�(g"O�����\�Yp���Z�๋"OV��� ��QQ���G���"O��0ao �j�
DA�E���$�v"O��R� .2�(�3�+��1A�"O"�Sb�U�0?p����p���Y�"O �S�g���8E�*�� ��"O���V7�|rҢ�555����"ORbqNY�D��0ض`O�p�p� �"OX	4��7!֬Es�O����8�f"O>�⁆�V� ��4C�t���"O�CU�<nYKW��A��yZF"O:+u��{��� f�%�l���"O0e۶�ٞZ��8�*��Wu��2"O�y�Ĥ
����*�	J�k�X#R"O�d�۲[�4�Xp蘝/L��1p"O�x)��FM4f����թ.�Ld��'"�$�4T
��U�߀�4@���V!�䄸~v��!]=(��i�k�$8�!�K��a�4�1	IX�bi�!�!�D�/x�4h!�D��X:|8Y�NV�c!�d�|�|��Is9L�%�[�
!�$@�_x��!%K�2k��Ҭ�!�E�N�����+!(y�v,�$�}☟Pf�CtX��WAC�.���B��?D��"�Bf��`3�iބ$_>iP3�i�DE{���݅W�p熛#R6�m!���'1��B�"��ՑV�ͦJZ�A^6,y`��0?�V01ްYhȂiy��z�eG��ԗ'Y��F�� غ�%��R�,���']�9y���0��L
��Ve�L����'ӞmBfjO�3�]��%λH�F��
�'B0�(1i�3����C�?E/��'�ў"~�6`�pr*5a�X�?�ّ���v�<�cF�*�\��'�nAr�#�X�<����f0�9gזm�jp��Ƈ[��h̓Bh���?\����W�f�d�D{R�'A�@
��� <I{�b֌O����'P���n0�8�����	B8� �'������њ��Y:EhLM`�eH��)�4�K=��ȔNV�b3�����B�y�M	��*��[h���_Zİ��4�Px�H���õB!0�x�2�6�O���M�K|*��P~��	��;�4[p�s���0=1�&Ƀl�1`�-G	�����FD�B���OV� \`A�$ˀ�R�L��.k`1bҀ.4��@�O�A��u��� O�t:�B5��~���� ^bu:�C�?@ۚu1�E��;.!�$ޙ_<�pbG��~ڐ�ӧ�F�o, ��e��H� ����+6�2�c�M��uKB8�"O0$�$K�/^�
T
��W@�<At"O��4l��7��pW��1,/ H!Q�'��I�E�b	��3x%������|J�O���D٨:����̑8,Zfp8��m��$+��ȟv��pK�NS�!��$�WdF@k�"O�5��ǃp��&C�oS�[�"O¹cR�Y���)��@8�X��"OHR��Y�G��x�	�-/L��6Z�T��Ajn�<%?��B-�N�V@�U�����@5�1�ݨ�r��Tn�S5 !�g�x�>Yc@(2MԦ��?E��'mv�  ��@Ä���(�т,4�p�w%��El�"4��m���"����yxP��D�����+��|���H���(��q��	O�<��'nH��&D p�v�#`�ȼPy`���'?��P���<jX�ɷ⊒t�$��'���[ �^W�y���7�� �'��r�^�'�L$����-����K�,��T؞��#H:�~�!a���x����ԇ��<����VF�DU�&�6`8C& R8�$'�(�L(]���&\0�W���Dy��R�<<ɐ��n�v�;� 5M&���$ڎ���U�!4%�����	�~d\�6�d<LO���ŕ�l��e+�i��r'(�����(O�5�O'�����؛
P����K�9�"O$��"'�t��
�k��j�b��O8���a�T�g[.M�3�؉	��E�'9D���( "oKv�# -r&�i��l,}�F�y���O���$�j	���'^`�Q
�'��\��	"f�,Z�fʈG8��9
�'�V84�+)�L#�k��*3�\zI��G{���IH�L���Ό4J������6�y���&�p���eɒ/�J��b� =޸'�ay��'��b���q�¨�2+[5l����'����	�2 ����&:�Y+r$�eӶ����y�%��$��֝�m�B��%�J�eԹ�b$�-
LC�I�?��eQDn�*ip�Ap����a�2OV���O�a11ώ1m�̺uI@3��|b�}R�)����܉��<c����5 ����|b^�b>O�����n��T�5�Z�gdD0[��'ޱOjB쒬kP=��	�VH:T���'�.Y���1Y�����޴X�p�z�HM
+R@�=�y��Pf)��lA�=?l�@��A?+
�B�ɡ#���%��/Yy`¥1�ON\Gz��D�x��K�K�G6�d/��0?�-O(�d� 1��&9&�$ҳ"O���D�9~��	�MC�����^H�����'2"w� )_y@��G����y2��&+4R-;򏈞N���s�ꄋ�y2���R���`4��Ld(mq�hƢ�y�d��h]�0B� œ�z��$�~��'F"�@�@C�G 0���1Mf����4 4	J�"A�����Ao,K���ȓwy�ɀ��*�� /�&QҠ�ȓh R��v �u�DH0��ˤ
�T�ȓkR��uOUqly��M[$z�~͇�R-�XX��.&�ްX�J�	�p������8)�U�H;�
0�B��eh+$�`�áU9���{akP�Β$간4D��(P�_ ]0���BI��B���S��1D�� �\y�ęp%$�� _*m��幐�>�����7?�hቲ�J	�2�0�h�v�!�$�2q:}�E@�!zf��!���'0ў�>�1�31�0��95� a��5D�Q�B�U�U�WA	�,d��0��4D���j��r X�)ȗ`@��3�5?�)O,�O>A�1޳4`j�{U�S�/�Xำ�5D�(��5b���Iu�T0j��h D����-ߛy�օ��GU*_�4`y�c"D��;7�;e8��s1�,"�B3+.,O��<!��^*}6L����F�;���D�W�<�TiB�k�`����.:�X�;Co�T�<����.�N0 ����bφ];��L�'�Q?���g���kcǈ��%J��0D�Ƞ�H(e|(,Id��R�nm;�˭>9�'\�O�>����l��l�8E�:�6A9D��R�
O��I�	B�E�����*�	vy��SC��Q@Q�#]0�b��V�B��3`�X!���`Y,[���$�B�I��T]˷�1J��@8b�zB��?�q���E�%����L�#�JB�	,p~�t;Q闀X4�� ķs�.��P���~*u�^.!nb]�֛&bFy� �~�<��Տ`�J0Q5���c����؇�HO��}��\ni���\����C�@�U��3-��$Q�z��)�G%HW���ȓ`�Ā��+�s+Jia#'_���`��MK�I��U��q�$�̏t���o�<A%U>v�ec���j�s\�<	���.ғ.�9�_)yy��Al����' 1On�sD!]4=AT��a�0�y67O���d�0D�jĩ����b_�K�qO&7�|�Z˓a��b?CPn�Jv���"� +2D���5D�D�᧟_D�MQ�nN'zv* ��N!�	 �Q��O-n4��,J�..E��n�.��e��'�p���#Z^��K�5�^C�'���N�`b��b��1&ah%�R��y�#�5#���0��$P�L�S��y"� a���CO��R����GZ��y��DT��t�V�C3fI����y�AM+�L�"���>Jf�cg�2�y�Q�)&����J4;s�R"L9�yB)�<������1�.|����(�yB��=��"�ُ'[��Cר�y򯄜zZ�ك$l}a��2�yR,MzP���F
,d6�8� �-�y�%��'c�H3�F4Cr!�o3�y��P
$���&�*=��x��ך�y��)&�0A�K 2�<H���E�y��	1;��	��cMa����$��?�y��F�zF�����9]����ӣE�yR�ڍE�r��F$��a��O)�y���#sT�A5��S<PUY��yr��lS�xӉ�*Aw��ɗ	��yB���0��)�q�!$�b�X'���y���a��( �j�)1��	�� ��ybIu��A���X	���V�J�y���h<��#�I�ԡ˕GD�y��,���ɟ���kU���y��O7u88�%W�u��t���ʸ�y�fږK��d:L�{�J@)�Py��Qq����#R�2l�&KA�<�5.��\Ir��l�ثB��E�<��
I+ ���bP�*ڰT�P�RV�<� ���` �}kV,�5i�A��"O�� ����^�U�5kT�wh�0��"O�y��l�����{��[Gz�#�"OdT*�KW����V,"5٘�"O��`�J��,P�m#�! v"O��W`ȅR�"tb�)ߗO4|�"O�\K�%�&6_h�
@���/��5"Oz�Xs�S�p�& 8�Ѭzwp%a2"O� �F�F��A�a슐-^���"O��&`ʩ&��,@ӫʉE�衕"O������ZH��k�=dP��`7"O��A�!x���ѦA�.K�̈*e!4��!���PI	�E�4.�t!�5�+D���暭*|K�'����u��i5D�H�ǎb�
ܡf��IH�p`�/D����l�fz� E�mw�`�r�,D��� ��7�R���H����F1D�0�k�#"��ٖaF�ml���#!D��z��O�J�%X��G	'Y7�#D����	9g��3m؞Ҿ�*��>D���@��:�dzu"K}p& HB�=D��ӗ*��%�Zai�-J���L;D��T��,`}Ӷ�r�ɫI,�C�I�F2B��	�58~�
An�8�fC�ɗH��)S��1�r
�I��C䉵AdмfkӠs�h1�Ǘ� PC�	�M�D��6� z��M� ��"�4C�	;c�ƩifiU�P��e�2�P�R��B�	��V�4m�}	D��hnޭp�& D��4IZ�(*thc� I7A�QJ@4D��ȳ�_�*��`���s�Z5gC0D��Ҁh +*�Ĉ�%��-�0=��
-D�Г�$ ����d_��J4g/D�tp�ˮ1����(Y�&��$�Ҧ0D��4K�57��]�4O�
��Հ�&%D�p7ꔊJ3r�a�#A��x��� D��[잕a (�eK�/c? ��dn?D��"s�)B��Rb��b��f�?D�,�3�r�`�"aւt��`�H=D��K��ȧ>���C�$(��D�Vm8D�t*�
�(�,8C� �_�\�3D�D@!ө!z�<���3ft����-4D������[ZDa��T�[yjI��3D�DZ�l��K��Z�̓� ~r��g���X���U�g�a|bj��:�p�2��V�-{����
���0>�S��T}T:���QQ���>���CY�m-���NTx���	Q�H �j�;��a�?1C���O���Z�0�'_�l�v����>�#]�����Z�AG.��O���H�&3�<�R���q�q�t�>����O���gGO�O�vU��B��|#�"O�(�a�;ʄ�C��.�2Dav�'d䤃`��:!�ɇ�	�*�X��\�>W�DBH�}ߐ���G���W�Y��M#Ǭ5-��4�&��)`baA��K�<�0'ݛE� ��7Id���˦ �6�p�ddӅơq��sSY�E��F��c��ٌ��=�ȓk���{��"0��(��
K
Ig����KZ�r#�8"3�>1���O����D�+Rc|YiE,4ہ"O���d�ǎzVh,��LF��$�'�|��e#n�е�퉦�Q��$���h&�-0�����33�b��e�Ov�iKvY�A�+A�7Ò��a"Oh�#v�L�q^v�{�I�'A�����ɹKl�3f��.9����O3Dԍ��B��|�~C�I�2�e����-xV�Y��F;`N*C�	�= ��0�Ӆ{[|ز�S41+RB�)� j�*�
R�_$��faҊ8�x�ˣ"O@�Z`	��t�Ĥ��2��x��"O�șF�� ,D%IW�A��Y*"O@�$�%p���r	�>�<��a"O���� J-%�lp�hR�d��d�b"O�8b0IM�c�����n	%(6b�"O��s�lP�K��<��&M�& V�S�"O���� �̩��.Z�ٚ��'/��C��\��$����.�&`�Y�ժ^r	��"�BO>B�Z)�N�PF���OJ�r��ݵ=����çEI8pB�+�^{�m��J�S��ȓ,x�p��ϹaR��0&cO�?�����O����?�������d1 �,��g���%x�hbE��2D��'J�������
�W1���%��Z�R��b��t��"�C8[�u�'�lpZ�R�Dc<��7o��1�$$��|"/ 0�",�OS$��F8z��)sY�`P����|h�IU+[&�n!Z��1�O21����Vo>�U �3=� Ū��ةn0<A�F�Y�4ã�Ю|@����#�Uj6��u +�s�
|iw�7O�5��819#��;:۶a��hA�R	68���u	v�@mP��W������c
�Б�A�/Ep!a�o�9=���:X\eqsMZ?�n �!��=�X��j��Y@���b��Q��"�-��ʧ 8�-�w�
v?��J�@E�e��ظG��44����!@	�鈌��>a�����ږǺ� ��Q�$up���(l*x�{�)��^L2��������bG:����+�����N�[��4J��Vp����TT���� �
Z|$ݻpe��6�:���C^b��y�f��Z0u8s.l2L�e&ʙEi����ER�5�6���E _c�9O�)j�0z�\��
ɗV��"S�	�D�S���(v5Fɲj�!Qnzps��Q:?r�ps��4M�*%{4��0P�콰�#G�5�x��S1@��+�~>#>it(S�UA�d��d�čk$��<I%D��FNE�1�]�B%4h���VD�l��'�ʥ�"��8�� S����ɴ���a ��J�X�s�'���
�/�>04P�m��Lip ��I�E�̰��C�$�`��T&Fk���J$o��:>(hR-v���X�=��I2'ٲQ�J���� ?j��Q���'�.�J�̏�?s���6��	ad
�
>�$��凝�j�����P@�ʱ��
��_�ݚ���91�\K�SM��D���[�Xy�!�� �x��d��ԑL�&P��+�7AQ��O��+�T�� �UX�(� D��	͞:��J�< �I2#9�ay¦T8b��t���M)6&xEz"��~��C^hZ�yQ+�
Md��ʜ�\W"����� 5�P�=7���eG2<&LR4b��X�8$M���x" ��=���!b8���b�`�Q���o��G��&`>��������S9G�h�K�,K7��5^}j�jJ�R���%�O<�@���#W6�Ie��,tgt��$@=ά"ŃV $�z��JM:Y8��,OL���Hc�
��ޞx�Ҹ�U�ɯ7#&��2HL�9�]l��jâ�[�Y���7D*���$�4Q���!��P(<��D��>ںY�D僸of�l:e��`~B�Jp��t�d�ޏ@���ã��6H��x�}�5*F�9��s@��?.)ZBU�<郠C�Q���k��]���[?b�HP�O>E�4J��|��f���LѤ�y��'�R��iץ[-j���!��K�^�0�)<O�IKʅ�F��`��/-�pՊ3"O�j�悩]��a(P�ZdT�C�"O��a��ɺa$XD��Բ}T�j�"O��A1+�dq��s�ƃ`fF��q"O��5D��>ݣ�V	i|��Ӧ"O�(�@)�` `!ɇ�lU��b"O�|p7�u�hI�H�*N�j�"O����i�% � �N
�"O��"�B �V1 �Ƕp��q�%"O�0"5�Q�1f��
��L�Vy�B"O�$�QI_"<P��e�N�E����"O&�����&b$�#R(^�<a�1�M"�޼=c�!���$��M�T���E\.��[��Rk�&O�N�K��f2z��WJȪ5���J�>�ԅ��I�,��Sq�۱7���a�߻X�&#?f�@ـ�)U蝍����2	�Eчiۑ4V^�`B��
w�C�� >.�Pe	�"[��}�捚���J,��įb�����
-�l�QE�6/�Ly+��R��r�
�"O�D�F�<0�(Ѣ�>Ć��Dg����
y� {��_�3�)� ����:-\I�� K�D��!�'<�,`���g�,x�ֵ�|���AQCD-��U��~R([�yX�ؠ&�R!$Ȁ�B��O6��bF�6���2qI ��.�;�|iV�:�����yB�XQp�UK��7���a�I�!��-�ɵ&w|�(i�2��\������Y���jb���-O1�J��  <D��F_�� ��	�{L����!5b��%�h�2i
σj��e�&��H)�r�M/I��lY=�>L��I�vcf�'�� ��w��Y��	�t~�ʤ�B)�(�R�mNX؟����"��� gk�P�E?a����?O�q�� 8i���R�I1/�8yVt�Q$̤���Z�"O�É�"n2<0cT�X���P�/�=�qOt4G�,O�Y
"��r9D�0E���,�2$"O�Q���表���x�L�jr���2ݑ�'d��rp�E�2���2��#A7���[nQkL����D�*�d���EQ]6X��1D�L��lTi����	��\ �-D��	Ѕ[n0�I2����$��g�)D��8��[�@�r���M� u��E�Gd#D��T�\{�x����_�y�ܕ;D�#D�ԣsF�:x���C��t)z�O,D�l����%1�2���N�0���+D���dIs�a��dջ���cՌ'D�p�������H(1��!�ĈXG�#D�`���R(��l��钤n�}��J?D��5�O�z�RT��"��|�"�,Q��H1�<)'c�4v�6p+3��;A�xٸ�nKH�����7_7�� h_l��Q%$f%�a�%�H�cЅV?PHQbp�'��@�"�Y�P�ȕ��'p�)y�y��ڦr�9i;O�a���_ޢe*G��~`/Җjܑ(k�K��&��y�<�S()/b��4�ʌU vQ��ϙ�9��r�i��E���Ĭo��{�0�S�^���ϻf�0CŇ%ɚ�����B+���Ɠ
�$#gKO'궵X�N�e��y&`ɲt��PR�.{����0̗1j�	���(O
�cH�?U7 ��T�ܞ�����'5*�Ȕ ݝ��m�! p���O+��h�� �32�U��g��hв�
�
�|R�;x~��2cƅ�a4��FjS��`1
���Ғ0�6�2\lԄ���7�Fy�O����I9l�Vx@IJ�`(i�'�.�Y��J��i��c�����oFe�7�T�N�d�P�v��I@����p����HlɑG�r�"tQ�'Y�0���D	�4D9�q@B3�b(�����{���@Ԑ($��4z��A�"to�"��!������R lJ���t
zx��	 mF����Yu�v`�x�(lY&dΦz��� @�3)�HJ@�C�`H�D�)�N8�Hc�둕��i��̝?X�M�0D+扝>\�Y�p��<� I��e�����e��B�iCT�Ā�/P�>j�У ���!�$O��X���1B�t���ڇ&���AX���&�$F�6(�� ���'���C���)cE���H����Z�!�D� M�P]��w���RcF){Ҡ�$(5�D�)z�>�'����P� �`YgC�
A����3�8��j&!Č��g��Ҙ�ȓ&��	�Qh�!ȼA�FЯ�\�ȓvTP��u��8F�^��D�\�8�,���<�P�U�U 9������)FŅ�?��9�ρ[Ȟ��"��0tw`-�ȓb}{��ɺ,�T�+QNP��d-�ȓ=开���[qF�	 �V/a��4U�}�/ޏ!����FE)�I��YYܱCƌ�^_2��ž�h �ȓ<՘�y3��C��,�`��4+���J�*e��̹N�f���"۶����j"��?߼L��A%h�\$���lxu�R=w�"� DY6%Xلȓ6�0ԉCfE�Y��t�&���9X4��h��P�������&	1f�5�ȓt݆1��n՞YÎ�@TF^:)�}��S�? Нsi�)��H�QBT�a�b�1"O���D�3
��-�c��W��p��"O^L*�Ǚml�����1�a p"O�hh E�����%ō*�x��F"O���ό�ju�M��Eԅ4�ԔP"O,����?<�����Ց7�L���"O�� ���H`L%���D%�q"OP�P�]�~ժd3Q�L�E<lX4"O����eG�<�t�!�e}z&�R�<1�	(`v�T�ӵXt}�L�<�@���,xdCG�n�pRj
I�<�G�R�?~�`!J2L��� w$�@�<���U
��8�L(~�8(hA�{�<!�0_G4���萑@5��s�h�j�<��!E(Fԁ��	5I�z9+��Eg�<q3��;.�RuR2dۯx���G[U�<y#�;^f� b3D
�B�F!+�Bu�<�R-=D�x'�':�bA�abGm�<�2�E,l|�1)��x�Q1�F�A�<1�K�&��`�u&�퐠���x�<9M�J��=�r!�&:6F���l�<�b�� x�8���]��2fd�f�<aЂ��&af��;��z�{�<����?��ѷ��D���MVu�<��H�b~ m`�#�v�~A��H�<q��ՎH��8
G$�(w��pD'@G�<Q3�@���\��� �L���Iv�<�[6S(՛�x�D�C���H�<9�%lTn�a���:{W�RO�<q@���5���pb�y��w��K�<��F��,�ѡi�$���дXG�<��ީ8���;P�O#5���B�<�E#��~< Gn��$+<hD��A�<yp�@)�@ƢK� q�d��x�<!��-����%̸|��XK�hy�<م�>G�͉6)M -��Ce�t�<Dd��w�r")��!>�� &�TY�<y�EA+>�nP��fS�_a��T�<�T�L�1� ��`(A�?d\衱��[�<A�M4y3� 9���"M��t��R�<�$�"H7Tx`R�R�+��ٕΏE�<9�ɾQ;"Iq� {�Q�$IA�<YA,�;>Z\%c���8Zlj���A�<�3���x�T)�ҡɡ���IaAV�<�DK�gML���'��g�N�<I�a�?�r𪕢�3�^�h� \K�<1qD�=KrH�2�R�{a�C�F@�<q i�*Tf�!a���/��phH|?9�L��-&~���Ԟ �q �ѹ�P�+�.�a|��\(w���G�'�(m!���*6dHy�I��j: ��'[&�`wT &��@���b��DÎB�Ԑk߸P2��\h�Oa��)����5�(��fĚ^ȨQp�'d��lR(���ᡏ^�PC��[�%�2��	;}����-݃'��0���|��ac;D�#V�!������3���ز��Oda �Z�-�^5+ۓX� S���Q2�n��980Ć!�L�CC�-Z��bZS�8S7��s���cq��y�� sE� �p�
+f��E����' �|nB+ �����	G����apA� L�(49����6!��X�l�1�
�,�qAbj���a�]��X�O�}�+�q��Q�L�+D�&W0���� �"	3,�m(���]u�m�I"/��,����#�a{�C(�X]�"ED}�f���F��0>Q�W�Z2����6~xsS�2~�M�c�X�gOP|��S�? ,���͝u�2��?YG�T��	�Q�$���� ���*�J�2�v�"�Hئ_�C�	�LN��Ip�T�Qa2�9ǂ֓��C�	<@i�H�(�)���i �$@�B��)Ev�j��H^�ň�O՚8��B�	�(�>-z$.Q!m�ղ�I��~B�I�+�`h��ܮnְ%��L�$[TB��
`��{��+DP�ݨ�$���B䉘@C��"Ƨ�5<�0�e!^��B��6kr
|� �CO��0��M�3?�C�ɧH_p����1D<D=�EI�$��C�ɪX���%�� (~̩ԧ� ���d�OT�s�/}"��)����G�(z*D�i�%���yr��4ܾ�k)�m�<;�b���	��B1P&��?!\a���;6�DS�d]�}�z���k��yB�V�u4���0��=ud�*�#G�d�IWS��Y�j��c>c�ls�)G�A���-D��QZ�C5�dS�)�*���˳$�h��b���.��R�O�8M
���ɒG�
�Y��S�Xg�\�����;v���d��&���Z�e�?w˓(I�� ��=6F�8	�֖XHp�ȓFa@�:�j��# ��#��UmZ�U�\������h���@�#(�Q?7m�/�=�3�9-/0q���T-!�����2iA*(6=�ܳwrahaNܪ/���b���|��џў��S��"Љ��3r/0� B-ғh��9F��<yfN��EN���G��4��;C��.LI��(櫜z��3.ݳ6�����y�R�j�˃ f� $<sf����mU-$d�,rV��S>h�rYC們0�Z"�I��|�]1 �!�s*U/6�s��IfB�I�b��`7���+�0X����a��� f�Qq�r��b��;K�8f+k>�pgmV(�<L��ԟ�d��2G�q������K4Z�{r�I-Y�l� ���3G$��&P�\���*:��HR<l���M�/U��cȊ%���I }����,	_�fT������}�� �5�GȊ3ζ��ɕ+�XQ��O�,Ⰾ�)2,l{�@���{1B�#�Px�x��4���г�!��p��}����,��6m�!69�НcX�j.��t�;8��;e
Jps��K�
�s�V)�ȓc�\��KH�3�P�gc�q���#��Z���Ӏ�
&{3�59�����#M�,'�:���i^������"Q?��ש��'� ���G�u�"I�T"r�=��ނL�.,��Q z���Nán�7�[�'�!*oޠ`����ԯ1WJp��̓%X�|d�GkAZ�O��b0�V��tI����d�$��l��+L�m��*�쐑�x���'\$5�x	��'�����#7�h�H 8:X��S �m�Pa�#���x��9�H���1\ `  ��P鸱�r��|�C�	@� �CN�~bMhB
*}&�6�V�fx�ux"Ϯ�Z`y��$O(��,�(`�yA��Sp�'��a�GĜ?�<4� �
?af@�g��(�R��9|����'���2��ʈ!f�=�CoR_~�
���@�TcFu�NAE��s��$�]�N{ZU�cnR�F��Ӄ���y�H&ن�����3��0��H��~"�^&D
|���|����j� �h�vjД�$�*vx!�$�`�L%�n�5*��|��C���'Ub��e�Gx��#5!ܿM *�
Ak�� "�hj��9D����\�L��ޭJ*t��ł4D��3'ӓ'����@.��-4hE*��2D�4c(�h���I)A�\���1D�x�!��B|�5�1��6��x �.D�,�Q
=IT,)	�j�76����RD*D�����H*� }"�)Ȃy�%k+D�4�� [;[x2��5�]_��e8�C,D���f�qv�����w�t�i!�+D�|���\e�� Ƃ�:S��Q�F*D��y#\,nM���8v7����l+D�,��#2Ŝ� �� Pp`�EK�b�� Qrd�e=�3�I�
l�:d��-ڞ]�3N�5M���ٽi�d`���%��p�ָ�%�1��t�2C�hc�b֏S�Q�0@ aʣd��F~�P�}��:�a@	R�g�? t��2��)�n�B��]Bf"O,� ��jXg��W��	*�\��p�A8n���t��	�0|2�⑊`I�`� �˴J@xa��&@�<iu��5_�:�@P7`nj�1��?U"��@؎��1GQ	Q����'��Dq��&,����f�5#Tx���}� e��L�!��U�cf޿Nn��P�*�z{ֈx2��p?QR`��s�z<@�V�X�IU�\A�')N�;c !p���~*6aT	l,�US .W�ۤ�+�F��<��L�}>�:��":B ��!��p}�)W�CT�A��^n���I�|c�X�4�\\�h�mЈ?]!�DT[S�X�bH�%�� �� �N��-O�|z�(˽5�&>c�s�.�,��Cӓ:T�M��,�O�S��F�W�����
W���H	�C])X~�QuM�/۰?�&�^B�윢��ؘ#2�j�$�v�:G�����%��hѦX*h�r����2�lp�E6D�	�f#? �s�#k�V���D6D�,r�kS�H~��R�1c�"#�4D�0XF
�&mn�1�dᑀ7�8��
2D�P��̿_���#"�d��<1�e<D� �2�L-OŖ!�Ҋ�*��\��?D�8;4j��I�d�v�\.y�����)D�hH� A)m�H%)�%ڈ�J��Rl'D���!�9a +T�s�� ��kG	w!�D��J%��'.K`&l!����;c!�dsLhEZ���l�����qK!��NJ��� ��FhN�(���#�!�ߣR����� �Ui�����&"�!�D��������3/VN�� J�)C�!��U�)
��VA�6WS ]��g\Yp!�䇶SX.�H��_(,S,���Œ�AZz`+���G �(��	%42񂇌��G � �1+�prP��đ$JjĂ�O2l:3FĹc�� ��Ne�\��ůN�2aL�F��0��>Y6ǈ�3,I��o]�]�.�p1̙f�]�&�XaL&�y"���{�ډ�-B	��ӣa���4��b��L���V�s#C�	p@H5Щْ}�.1��T?@���8g$ԣ�MS�OW�%�*���(�0�q�B�+��x�Q(uB�9(�8I1H/),$))�64� �Q��(.��5�3g�>m��؂.�(����ނ8q����Q�-z�cB1TV&�Gy�G�u�\�xǋ��F���C����<i�k�@��ٲSrӄ�p� �nu���(ee"(C�W�f1R�W�
&`�B�o��8��Ю��Q�?	��&���!�����ƿi��1���V0�L���AV�"+Ѷd�0�E��/G�N<cbGKq�<�'Ñ0^�����+:6��bጒ�{>���i�H�!�Gǿ^%�I���c�'Y)�y�we�h�!U)fJ$}Bč��S�DU��'O8��
��-�v�H�<�Њ�z�z�ѐ�P����bBa؁ϔ�6Q�<x�U�ːX� gI,m��䳂I4<O�P�`���n����4�� �^n�9�q�ǒF&����3��Y�E���3|��A����R"N�i\����e�1O��Uf�g��	)$�^�����_fքY�O�<T��O.PC $���[�)�:���'*�2i>̹b��<@�%����DN
[Ĥ�A��)	�B��wL�2�Ɠ0%u:a���ѳ<�0� �'H�@��C�:|��iL$?z��qv��5�'{��a��L�*� z{��1.Z�?wf�p��4D�8!��ɗnt��"2h�$����5D�$Kæ�!��Ruj��bXƀBK-D����̍�Q�|EY`�;G�ހ���*D�����Q�h2V��<Eut�� %*D�Xy���LKFъ���)�"쓥�)D�4�@�CoRMr&KX Z�����,#D�80T�R8u��(�FY�e�贻��#D���0��8S�p�WgݒP�H�� D�,��E�gp��f��=u���1
*D�DbT���aY�圳�괱�i%D���%��Sv�sE��d��<(��%D����肓P�V�if�$���Uo"D�� s �ȩE� ��&d�?"�f�0E"O��q`��;KS`�Q�.H��V}�P"O���e�X�5�L�!7��5l��0"O�e�A�&/�<:BLH8 �i�"OX����R�}J��TK�"O�a@�#�a�|��j�)j��=)�"O�����̸�	T#�
1]�`9�"O��)��@(>� ��E�,CVe��"OP0:��J�(�d�JDV�Y?}R�"O̸�3���I ����R67{�H��"O�$B�����������<�!"O�\�w���P��×2��䋕"O^���z��;�$Kg�AJ"O�x��G�3+u��U��	|G����"O
m�׍�/(�h�ơ�b!���"O�����X�y ��Ң�׉A�bQ��"OrEQ"X��5FT����"O���B��+R����ּs,��v"O¥:���)~���M�.̊!��"O�<Մ�|��	�mUG>1�(�>��mЈl��6�S������?1�t��3��k� ��V��Wf�O�8�O:� ��>��<%?�À��>A ��ʨml{�-}��Q��8�=�z�IC�I�ab�B6_a�9�C}?Y(S�w�㞢}���]�X'R,k7� �k����F�n�Q�e�r�S�Oz��K��[cɐP�l@��l�Ӵ�/��-w�a��F�JYC���kǮ����$��N����K:���?��~�vViڧ���:���q����faQ��<��}H�j�dU�p�v��(D8q�Bj�s�,���<���)�'o�&�3��L�?I�D��I�b(i�ɸ�HO>m�O�8>�QsGN�i7�ECEA%x�D��}B)����|D��#ǈp�r��N�!h�`��V��ϸ'��`#����DA%�R `3��`�R�!��W)��I�$�>#<�*��
�st&=�`Z+0_�kE��V?�#�V��h����B��)D��=�'@&g�lur�"O�(e�J̜s�$%���v*�13�x1�D+k�ܻp�@n��̕'��R`ςE�4F&§_F���+�	�<�`	�f	�\�u�_?q�؄3I*0C��:����cMAj= �b2�8�40���O�T�aVYQ����0|�A�ZH��O$}=�b< t���X@��d���L<��f���X1�?[��i�a�>pt�h��	"�'}���JE��v*�(��Q���ܦMn~�D�|��&Mo|��遉P^"i �ʫz�-q1�L 4��'��]S�B�@iJ�~:ٴ�h21�L�[�ԩ�b�X�`���঑�eKߺ5bP�+B��0|RubX�� ������}�3LU&�a��+�+A/��sQə�<Ye��O���!����v<Ӡ�!q@dр��:�C�H'�O,�BQM!^��C�C5����"Oz�0���:�����3��x�!"O�\k�
'G� �c�C�7�r��4"O8��9�$��tB����X��"O>azs(ZsD0��7be� �"O�x�
�(8y�8"N�@1�!�"OD��)�$6�\	"�2W�{R"O����O̤�h� W"�P���"O$h˷*A�f􂙙��XK�D"O�P$"�9!n�2�`K�RD>a�4"O��`�euƺ�A��;U1ޙ[�"O(T��M\!18rϛ[-*t�p"O�Y��_w.�:��T ]���"O��� #;�̤Tf+�e�P"O��u �Wy���%�38D��p"O�2@nK�s�l�
�KHY`�!"O�]��13R���Ė�N-�H��"O,A��A�?6�i��"�.@�)�"O��#-F*1Pu�4Z�څX�"OB�Y@���:��`aJ�)��m�w"O� ��{��H9LX���*�+u���"O�-s�MTv��%	�*4"��l��"O�H�&����Eq�I��gX�"�"O��Hdlȹ]֪�R�&O?:" ��"O&1C�nӒ)�(�"��)�hY9�'�V0�RQ�:i8|�*Q<x���'L�P���	���*@
�8Y� c�'f�0���Q�&�i��+E�6�Fp��'�(��A���_[�A�bւ":�ܱ�'�Ҵ�I$G������h(���'��S�L�#��H��+��)�'�J��L�[���ـ�щ7��9
�'�ҕ8V��d��<��dIH�TQ�<	�Ν�T��;0,�;N��QcDU�<'i�0H�m�g�N7\�|)s���L�<qA
=ln>��S�3��� Et�<�%m�l��'D�X�>A8s�YZ�<�n��}�����O[:����`�V�<!�5��!	�/�?=j��q�V�<����7��*7R�R�P81��N�<9�jY �.I�ě)4�n��C@C�<�B�]�� ���էjpD�s�A|�<���>��l�􎉣;M�l���[@�<���N�3���'�[aT�!��B�<1eFC�c�a8��T.F��P�s�z�<�'DG	Pݾ�G�+*�^ օIm�<A`H�rx���A�9A0�u�k�<�G��y�����a�l��%�d�<I����h�5!e�����K�f�<i����`x	�ڲ'��cǺ}��yp�� ���V�(|ȓd�� ݀�ȓ!�j��P��no$ܡ��W�,0�ȓk����Rkɒ`y)5*Ô_�䉅ȓ���, 	А@]j�h� �YV�<�0�N2��P 5A��-��&LU�<�bȊ9_զ���H�H��8DoLN�<)GFG/-��D�g��ZA�SH�<iff̳S�x��bN߈<7��Q�H�<�T�B&x$���o�4��i�L7D�@�D�{�:Is�`�j[��y��8D�`r��0 ��x��S��,J�$8D��p��J���soʽjF���)4D��b5�QP�����
g7�x%�3D����_�"z��a���P�ȋ�"3D�)v�#�XDeJ�[ �>D�H4 ��@�N�V��X��+0D��HD	�8n}�,ʴ��
F<���d�;D��B2���QH�,�̊�v��|#(?D���䐀4�R�+����FAs$�*D��+�"L2,�zŋ�"�0�
)D� �F�n��I�3�!m
ؐ��)D�� V3E;hmag�|���'D���qDX�{���T�:v4-�!'2D�! ��Ҕ��j�$m`4}Pt�/D� �e�_4�J�A�{��!J��?D�LB%Dةl^�[��/?�
�
>D�L㵁�,
��y�'n�j�S��!D�u�çH��l�7���bEc�k,D���@�

R�b��T�V�W\UaBG)D��C�暪g72�Ɔ�;D!	�B'�IQ���O��[�K@���E��C�A����'�@i{��*L� TjrH6<aX��':���q�V�Z�4	��
9a�r��'�$��
UNr`Iѕ�ŔHAZ�	��� e�aɳC���堑�l�4p�A"ODE�4�A�P&AzD�ʣV���g"O)�D�M~o�E���wwҰ��"O� � Ɨ�C�<-�T�ͽk�@r"O�!8��ʻa�D���VLYKr"O8H��Pnu|i8��(HdI�"O�y��QH�e���
^װy��"O�m����|��	7ŎŢ�P"O���,�a� ���߯�T$��"O���LJ5.�v����U��|p"O�ݛ�,^}�v	����X(n�T"O�����2�X�xץ�x|��"O0��*�"I�P@aC�G�LQ*u"O����*;ݖ|:"ŋ�D+.���"O|�� P�n�,$!A$�x�<�"OT�Y�Õ
d�f�s�&b�l��"ODX����%b�	aMO�{*��"OY�^%����F��a��n�<�.�DT��B��ȴ�����Cm�<�ڇp4څ�����XP�W�l�<�0��!(���4i�r L�sRG�N�<F�G�Θ)��I�X�@���dUH�<� h���5�5�h	#��]u�B�	N}|�Q�������ϟ$"�B�ɮp|�ih�M ;�M��e�)2yB�	:�D�h�� ��<P�ȥaϾC剽rV�[S(֞PP�(򃣗;d�!��T%$��H!�3_]���r"�-�!��<Lr�xk#�&U��ՋW��Py2!Q�yv]xE#,O�� �h� �y�ė��PQ��%x�Бt�Ӹ�y�ˋ/���p	иZ��T��y�	�=�j9dDU*=���@QA���y2d�.������.IT�jS���y�	�;\{�A�"i� �d\�ҎH%�yr�"|��c��A�� gLպ�y���%b�&$�S
�i b�4&A��y�l�;����3ƛ>]H��󇂷�y�G�8��ȑ%�<���N�>�y�V_���I#~������
�y�b��\.�K�FBY�p� O#�y�ϝ<��]<���z ��y�@�[�$y��X�ȸ�K�NQ��y�z�= �n�$xιp�n޶�y2��X)�(��CH
X�������ybCK�py�9�0�M/�����H9�y�F0��W��\o���1�K��y�� V�� 0�+OP��8F����yr��y0�4C7�C�4������y"@ΦH�\`Ⅽ�)'X�1l�yC�V�I� e5$�T��$IT�y� M�a�`��V
! �y�#�����*�@.ҁW\�mP�̙+n�h�ȓ��E�ɗ{��m#��R�~!�� ��Tc�E_�!��M�(�P���٬Y`�ncs��2u.�G��ȓL��¹p��Jf!@]Vq�ȓv H @a"3lءӂ�bI�U��H5^�{��O�KnU"�ʙ�Otq�ȓ?\`h���
;%F���X�1�f͆ȓTQ]ۄ��
��3U2lR-�ȓ�p@4%6/,�<P��+~���ȓBC�d�̡D|��jՅ̂2>����D ����\Q��?���S�? �8�敂((�E��b2=<��"O.2R�Wx3����2+*@G"OH	X�D�0B Ѐ&,Z��PDf�<���-p�ɰ-A�bPԹ��d�<�&"W�oc2	cT�:w �����F�<Y�l��pI��ܶ���H$B�<!!c 'I��L�ֆ��"x���"z�<�1_��Ї釞#mڨ�� `�<��&X���J'�Q'���d�\�<i���rrz�ip�>�D��!��U�<�G���R��ѓE�рj�}ц�Tk�<٣eI��BjG>^�TqY�]g�<y�)N07���Q��R�BA���\d�<��Ǚ��0ePdf�'����]G�<�P��,֚�(#Wy`�t)���D�<��e�-\ڕ���
&"��Xt.�g�<�/�Cð�q D�he$dV-�z�<1�"� �T�1��09��[��u�<��k�"�h���kF�p��@�0�q�<�r̘3,kbl[ՋӨu�0�(WM�l�<IU^j���C�C�<ǰ��sbe�<�!��u�n�tF�:|��Un_]�<��)�8�b0�'��Oi���tEW�<�bG�f�DQ���@�AQ�UG�<I�n\+]*��Fŀ�$@y��N�<I��:�H����*�����AJ�<Y�D(;�^Mh@���T��\[�H�<	�)�>�@g��p���#A�<�7��&Y��U��DA0|߀ux6��r�<�4X[��h�H��?s �Ha��i�<Y�aB�"�:xP�[�jH|��)Xn�<a�
�e��tp0E�2Z��J�g�t�<a�eI3a�TZ֝S�hx�P�LV�<��#��j $c�Zh�����M�<A'b�,q~5�U�ѽ{	<��TI�<�e�٧G<����S�0^q1J�A�<9u��4��x��o�F�$�pANd�<�W��?D�6���l�46�^�R�_�<�1G�;	L�	���0f������Y�<	��va��{��\�9N� 4��[�<Ad�O�
�h7C��q��Ar�<A1��x��{��ݛ�Jyv-�e�<��]2\����B
"T�(�4+Td�<��gH=k���
�7:謘$��^�<�� �LDȨr��D$X3�9��d�p�<�td�3ٺl�F�˖-{f1���
w�<i �7���s�ݐx��[� �p�<Y�o®�رȅ!D�z�쓶/Mp�<�u���4�d	a��V�\*����<y��:o,�R�c+<��'���':��D�t�~мxa��>Y�,{f� 2�� T:��G"��gz0�s���ҌqB%�'IJ�'+n�d�&�x���1�A�N�Il
�Ѕ��R;�[r�N:���'l|�,{���Ke�'z���"�%���Æ�P������O�T*��O�9m�<{R��<��?Yݴ̈́�����.G� B� ޤ��p�]�L��	
�x;�cۂe��T�
.(Z
�ї�i�P6��O4�m�՟����?іO,vT�cN�Y�=�5K"N��!�!�f�����'�B�')�Y��Sş|h�C�� <���N� Hl�� ��<Xg:��q���mT�����6C�h����"(�ģ<��+M���g�+B���;��С{� Y��PtV�(}�PwHR�4/)C���/�1O-CA�'�ԉ
���8C�r�9��.umڰ�s���`��6��On˓w���Zw��im�����녱Ը��I\�v�!�AESC"K|� �#���W���X�	o�dy�b��@"������'>�cIL�EN�@�f���i}�|s k��# Z�1���?����>|AIS<��"�I<&Ȋ��f$rōi����o��Sh��c��>9Q��y@% y�ZUC�Ɍ#jh|�`M��.V�0�n�EZ� R�̨P�h8��7�����͔��>l ��I��MD��d�i�L�Њ�&8�YXUO��BE�:��$?��՟|�	������� ��!U��W���# 2��帣�'7B6-[֦�m'=li9��۲~M���;_���I�4yZ�+ڴ�?,O��>[*����O\6m��&��`�eaK�B�"�`16�0	��k6�b��_�a���+���ؖ�&��'�5�hu�t5p�� ��9��M{���5?�΁���$Q�����9�Ë pT�Z-�kL�>fv`�)�`�p����̸��֌�?�g����"|n�5*X x(_�(9b���/X14��͟�'��D{�'+��=)�&[
l������z��Dy��lӈqo�ڟ��۴�?Y���u��.a�N� # ؊Z��u�sm�3b�z˓C�ri7�Ǵ�?����?��c뎺~z��WP���pWJ�
�<�g��|����A��M#!&���{��O�PA�L/���zݳ%�й����5���H�l�5a�V����o�J|��H��LPlz2x�G���3gfD�"$��嚛o���4"���$�O`5'�P���'�JD�ϖ�r��)ხ�<R��{��'^|8��	�����n�1tʙ��E�¦-�ڴ���b�'��$H�"g,\8gKU�Tf2�Y��P2V�P@1C�E.L�^���O���O<�^�˧�?I1�@�2j��ƤX�#�f�I'b�I��؀�.�=VH|�Q�XFL����r��eFy��<`h�-`*�- �Q)b�ߣ|l�	t��^���R��S�"�:��S�F�zδe��S�1��O�a���'�TŃ��1j�)����H6@�$��&8=(O����O��S˦��f�:���kg�ƒ;�%ӗ`3D��+6OYJ`�]J��E�	�Ō�� ��44���|��'i��x�@�$ \  ��   \  <  �  6   �,  8  �C  0O  ZZ  0e  Zn  �y  �  ��  �  ��  Ǡ  �  J�  ��  ӹ  �  b�  ��  �  A�  ��  ��  &�  ��  ��  @   a ~ P �' �/ q7 �= �C �H  Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�� |d��"O
`�(�;���8���-0��1%"Oj4��ND^[��"3/9�0|H�"OB���H��*�ʞRy=a"O�味V�!X��!&F�:J�$���"O,��a
���C�Ą�M�"O,$3%o�-���p���+Ն�:1"O��ݢ1����`���y14]2��i�<�6��{_���c�H�`�fX�$Kn�<��A̼VI�xR[�)�Ć�pඤ�ȓA5��('nߡ4�� �)˩%� ���,��r�؊b#`T�eT09���ȓ!�b��g��}�8�F��-? �ȓ
K|m�ș�VṔ���2�%�ȓ"R�X�j�4JN�1�˘X�i����̹	_�jZ��1!g��zܶ��ȓgil,*�J�
j�Ne��i�J%b���f	�(U��:���G��$Y^م�~r�� S�%T"���k\�jx�ȓ|4�1�îJb��@ӵ�ݩn�V��/[`�"�v4�R�!ʎ<��M�ȓ`:��z�ؚh�J�Z��$HY:	��H��p�m�C1��!��B:��0��EnjZA V;9����J[
2���	��4'J�EA�IVW&��~�(aZ��ӹ�>� o�Y�|�ȓ�f�A�
Ο7�H��M�$�����mޠP����/���ANXo*�ȓTv�����{ ���-7�*h͓+ZL�$ �Oh��o�.�l���ژN[J@	�"OF�K�2+T�<)���80"O�+�@��>mZ�B�-_ƺ�9%�	U>Ub���B֥XW�����(D�\�fB�A?��b��8g�����(\O�c��!�m�%5�8v�^&sgj��cD#D�Bg�	.t0@i��X+�hHhre�>��O������������9���a���*�횤�yŔ�%s2@z'������C$�~x���|8��S��M�=� �b���8�(�r��$,Oz��C��	� �Ȓ���C+����d��o��`��O���̉)���� ��W������x�_���'G�>y��	
�I��quD7{�Ē�h(D���A���*]�%��?.َA�r�x��':����'>§68P�N�l��D�eW��Z�Ȃq9 P�ȓ3�B��&/��2 �R_�7���=�[�8!���OJ|ca�"gY��Ѯد �p)	��wF�$n��Urd!X�\Q�:u��!�$S2*2(A6���ZD��Cd�,>��dR��ӪǬ_�hЃ�P�}��	|����֌B�[�=#�H�Ws*m��=��?�J��O�aǇ��LB�����<+��'(�I$ha�	�ʌ8�9N<!"J6�S�elj�������N����,=�ȓL����P�Ŵ|�H���#?����?Iӓ�*IS��U,#^uR2��8cKV���4�8�m�f#�I���K�	�x5А�>�e	n�� ���֚`9�IP�l�l�h1�OL��F�*g@T(����bI(-�x����5旝rg�H!&��"Q4:��ȓfҀ�0�A6O_�!#-����ȓF'Щ�ơ��R����K�U`���
0�-#ㄖ�^�`�6�֒j�ʌ��S�? ������V�E��,�+ie�PD"O�1S���:fD�1�"_7G6��@�'_��� ~s���F�|�.r�
�5��C�	<XV��X��T%��ψ>\ "?����W���ȚffF�$ޭB!�T(�tkŌ�7lq,+��m�!��2�R|*�HѪ.�r ����-*!�$�+��H���j�
 б�ܓxl�O��c!�'�(�7e�X3�a� �W��s�'���2#�C�n"��#�*��E_<� ���O���5�O.�k��G5k���  I�L��=���'�8��z3C���m������F�)D�@������ZtA��M@�+�	-��H��ħo���@D�úxf<�R��a�@�ȓa
@��(�d���3�hԮ �&Є�@v���\�&�2EK7�'���ȓV�V�c��M�bĠi�7y.�Ɠ1��;�jC�q��F
7`\�0�
�'4�T����nn0X�ʓW�h1��2�S����2;l\X0GC�^�^d���W3�yBoA���iu��8#�*�Tg��y�*�19I��rHİ\6q��
�y��6E��́�h��)�e�B���>��O\h�A�(�(���2:�� �"O��C�@�1d��ؐd�d�n�"O�Ѐ�=��pWd�%:gZI
��'u�Oi�P�н�\��e�~r�D��|��)�;�rɳroכ2��t��L5W(c��D{���F�<�*�ō(*�>�������.�O��t�B�PӂQ��':M�I8���b�'�b�!��P	B��\>�YcT�W~Ņ�����	|��l��ޟ!j���&ʫ`e�B�ɹQv(�����T#8Mp�g� B����+�I�a�"Q���6xmD�@�	;���my��|��i^,����@�Ifx��Fc͌v?��N���X��M�3NVĐ���j�� L�4��I=/�^a&fT(���P��h� C�I�@�T�87���{>�@���0D:Ѕ�' 84����ڒO\1��ĥOV<Ey�5��,��"���3��+��
�k��B�ɾA�XTkqAK���TRB�Ƈxf�O������	�d1��꒎ҫXpx\��>�!�d #O2\���+�f�T1�1O
��8<O>�b�K�7�@� Sl��O#�=�<O��=�'��'ppa5�<C}2�d�Gz� pJ74������%E��!7DD/w{�4��g=?�	�AUک���� ���0� �W!x���^ː�th�$=�T)ᨏT7�����LS��B.x�Y�QOF�'d:TG|��S�F܀�u��X�q��i��yV�C��&vj�p���S�U"�M�C�N¨�I^����V�!GnT�4/�,y�lG�]}�0�"O���m��JR�d�-Z���1�w~��'����Q�е(x}B �Ɗ0�*�a	�'ʢ,#`�R�b��᠐��#=*x#	�'�0iJd��=P�x+��)Ⱥ�����Ƥ�y��#�'Ql������XX����kFL��ȓz'�Eʗg�7<��M�¥J�&9����'��m~��9O6$rV���r��	�U�Vm3ON��%JMP���!́�n��@��g�O��OD����C��]y�ILL��X7!уi��{�d�m��H�b�K�tͦp ��K��!�I8]��8�.6�T�s�)���O��=���e�E�A(�h��	N	Z]���"O� ��2��
W�<��IP�~B�����IL8�Tb2d�i���S3�K�J��[ �;D�xZ0�� j��y*������I�+6D���2@�
 <r(:��-=3Ь��6\OBc���Θc�x��ʝ�|P����2D�<*�h�5h1x�y��V$�԰R� %��3
Q����+4�X�7	n�k㈖�
i�eC�"O�L��m�$k�J8`�WiPR�9"��`8�d!�E�)n3Tq	r��>l��Id�.D���M f�>��!��<Sa��`B��O��IQx��@ōU�i�8�%�!-Y*=��L0<O0��ē#d��y�e*N��B�ǻ?�� �ȓ|�n�UG�r0YX�n�#Yv8p��1M@Q��	��l)�	P2ZJ���V`
-�Fb�_��Wnc�"�GxB�'�V<Ku���)�0P��g� 9�
�'w�Ā��8�xKw��;-�.H�O�E���V+A���i��Ra��)q���$ }�ʲ�l!���M�q f\wf�y2��'=��P�Jw�������y"�H2�޸��fѹ{_��᫜*�Py2b
���3Ň 6`|�`! v�<I�Ť9��1�I�5�
����x�<)5b�6Y��y��&����Y9-s�<y�铋L� ��.a�Ɲyì_I�<�p��c��� ��A+0��Y�k�<��� �b �(4	qf+�_�<��j�9,A0��Ib޽H�#�_�<�a/�Nl�+X�M���p��Z�<�g�/8�����	;C8,�aV#�q�<	�j6X�*R (�2L��"�m�<�"
�$�\�����(H�)���j�<i#�ҧCJ,˖�ǎn�蘗E�}�<9�!T0HMEٴ��/�����Q�<�c��]���Y!*	b(��A�|�<!� ��4F���'���VU�5�O�<i��͚>)�e��a�"n|M�ӥu�<A爀:9�Y��Lp(T
!�q�<Y��HԖ������U��X��fEm�<�$C�&�1"�} ���d��e�<y�n��*���˶�D�;d���*H�<����p�t-��`���TB�<	S�<=����t�$on�1QjY�<�1g��B|�4I�,�q�X�<��C�y+(rG�=�:4�$�GS�<�lI(F���	#	9�!�Q�<���I0��詁dӑQ	*�\��M�$Uk�W9Vh$��E�*��ȓ8�D�aׁZ�f�9��2{$̆ȓM��$`CB[1?FAP �H6pXĆ�UH�P�ҷ[߼����_	j-�ȓv���ga=U��iS2�V�d̅ȓ<[���$�0*>ĹP�C'b�\��ȓj��`�G�HuUا ̟@I���sD��7��?Xw.4����W�D���c'Vx!0�ݺQ�⡩b�Y�1Hp��"v�a�l��9Yeǁ�'���ȓ%
�fgV�"�uSCP�R3�a�ȓCz,)�cCҾu��X;e�/D��1���	X d̠S���uI��uJu�ȓ@�=�%�@�j���!3r��@�����X�a�%Q,R"�Ϊ-���ȓ�L��j*B��EYdl�0\��y�ȓ/xU��&���E�O�o5�S�? ���ES��l�
D��#�d�9�"O�4���dH��a5���d"O��4��I��0)#ÝP����"Ob�A�h��M�b9�A/*ּI""OV0�V���%Ȃ�Յ����'���')�'2�'eb�'Hr�'�.��o�0z"Ȣ�ʊ�ureص�'6��'���'H��'�"�'q��'82d	c�E�/���S�&'JJld���':��'���'O��'V��'�2�'���q#��3���+�+o�P��'~��' ��'�b�'�R�'���'^ࢱjZ�M���3��er
���'���'j��'���'�R�'}B�'� ��&�A�����
~+$�s �'[��'ab�'���'���'&R�'�D��g��?ʺa
P���j���'�r�'���'�r�'72�'���'��yYg��pwb��S�ȩS��lz�'!��'s��'�r�'�R�'���'l|p��	����ׇ��3�\=r�'���'w��'�2�'���'���'��qQWh^�K^��gŬ"=�|��'�B�'e��'���'""�'L��'[���`L+m�v���
��-�@@��' �'���'���'4�'4r�'�4p�ʞ��@�0U�x� ��'q�'er�'B�'j��'�"�'���hhɃs��*�.x��'�R�'��'OB�'��,i�X�$�OLY�@�X-��7'5E�x*��TyB�'��)�3?��i5\lkg�۰Z������#u.�B����dXǦ��IA�i>��˦���$g C$�"#@�|�b�� �M;�=е�uA~��ٰC����H�\��,>Ѹ���M8Fd��3�$tC1Of���<��i�2V�0�B,@��(�nȅR4�o�&�jb����U���M�;|n���,K�c6������C9�6��O�7Mz�,���N֚4����<ySe�pS�ۧf�9IL���6���<�7E
>Wl
Ȳ����hO���O2#���B�ܜ�щO�@V���3O*ʓ�� ����̘'w�LI C�'I]2i��e&n����e�'1�')>˓�?�ܴ�y�Y�@�e�Y�44�� 7
^l�qQ�J8?�nν2d�$�.Si�'b�p;�NU��?��3p� �%�D?E��c5����<i�S��y2�A�x���@�,D�rZ����S�yr){������0q�4�?�O>�'���۹Y��J֪��r�Bs�'��i�ҧ]�A���OF�P'�])`�D � �� i1N�c�6���z�M�m�n�O���|���?���?��(��H�E�	%~���Fb�2C����(O�8mZ�Č	�	ş���R�Sş@22&׍s������?&<��D"������qڴ���|��'�?�t*�3S'ND�B�[Ŭ0@f�JT�|�&b����$��i�=b����O��_H	��H-gϠXB,݆ڈ���?���?	��|:-O��oZ	m�T��I>zu���U�
�R���A�a���I"�M3����	��M���'��6�`���z�Y��"�s`�QGC�|��b.�y��'��;��J���{�V�����ߵ���C$3�o�kޝ��u������|�	П$��ӟ����2<�$؝$)�}���Ҹ�?����?ᓱi0�i�O{�b��OLX�LA�L�~h��f�h	�@���M+��i�tȔp�6Aq�'n"C@;c�$s�N.fSz��R��r¬L�����-�\b&�|�\������	��4��
����@�U�N��������	}yR�d�F ��<�����I�p���X"LM5	���C/׶0�I���$���i+۴���|���xw�H��>w�B��
�77x��vǙe�(�C��"�����L�3��	��>�OD��`��>�X@��HJ"Īɚ5��O��D�O��D�O1��ʓ	���M�w�� ;w��B���˱)P��w_�TRݴ��'
��HD���^/R1�%'�5�����$s��7��){�H�m������� 4l�YR| �6(6?ё��jl�@ړESY�x2���<�.ON�D�O����Ot�d�O�˧ĸ��F^��U�5�Z�/�S �i�����'�"�'0�%mzޭQgX���5+TG�	g��������M+u�i�ɧ���O�2B��2Ҹ� �'�~�;S��j~��� �|#�'T��
P�V�q�T�y��|2P�����HA@�*%m�-c"b�yc��������I�L�Ioy�Ho�Z1�b�<I�����tc� f�����hH>��L��I8�McU�i��'���Cp�_l�$8�u�_�I�	ڜ'N�"X4��I�/~��	�?��0�%c��-�	+L�A�Bmw�L����Z!y����ԟ����@��{�O�r��(	�V���,�"#�3�Xj�rjs�T�7��O@�Ϧ��?�;�x��+�$`�i1s���H����� l�^�$��Ø �q5OP��΍lJ� I'�G3 0��p5	���H�WR�p��3��<����?Y���?i���?�T��.�$�aCE�l��ذ�
'������9�`�ğL�Iԟ�$?A�I�tȨ��D��X��h2��/J��Z�O��n���M�M>�'������r̔J���;�	�,���`�R�4E�.OZ�rf��B83�2�d�<�$En{^B�/*���A��*�?a���?Y��?ͧ��D������������$�c883W Ұ_$$�`�ܟ�#ܴ��'w��Q�����O47��3Hﴀ�oSz�&����Z)n����_(.��d�O���tƘ7P���� o�<A��ؿ� ��j0����8qč��*{�E@�<OL�����h~tD@��>1b�4��&�b�$�O���Ԧu[P�8ڢ�iD�'�lq�`��NSL%!f¸H��q���6�DPĦ���4���,ƻt���?�e�����MX�k!s��!�-Ip_��Z�j�����J>i+O��ܰ��¼_��*8��	Q��=9��v���b�'��T>���_.s.-C1C]%qFv8B��0?��V�8P�4]?���|�O���Q'$N��xRiH�h���QH�(f]e f�%*���e_�0�Ӄ]L>�R��o�ɂ���"�Ȧ/rT�N�9f}����<�I͟P�)�S[y��`�x5�A�43��d���r�`����Q'����O el�N�i>تOX=mZ�[��+F�TB�>`��}��4�?	!ϗ<q�J�ϓ�?�šF88t*P(����d �[���&J�V�{�Ț]���<Q�V�8Qi� 7����3���^��t�i*�:��'tb�'��
ioz޵���^:�(��𫈒m-����Z��MKƳi�.O�)��J�I �B&�v��^���Z��C�j8�G(Y:����)0�,��ùi� �O�ʓ�?	� �p�P��T$s4����(e������?���?�,Oim�	�F��'bN�����)U���T%ó��;E��'����>q�il6�j≌	{�1�v�D�s���� K;$����;g�3c�B��a�^y��O����3c	03��Y�6����J; #��s�Y�'2�'ZB�'r�sޑBrϑ�<�����/;�&�����xI�4�p���?���i_ɧ��w���*��L�V�i٥!�9, �'��6]�����4=v��2Ζ�<���p|9s�@@�""!IQVQS��ξ9s&��0�Ɂ�䓺��O�D�O��D�O���S�OiT��N<CÔ�+�͎-	^�˓ ���Ϝ�ir��ɟ�%?9��&q��!tm^�Q�J�Y�^�( �Oj�n��MK>ͧ���RM�=�&	��FC������AFg����5+.O0�z���8#fL�׌1�$�<�c灇|���JW��!J�t1��߂�?���?����?ͧ���ަ�D��ݟ|Ze���p8�͢�-��@��
t�埈�4���|�^�X�4O���Iu�lx�.\|��핦p?x+�MM�6�t��1O4���ְP�B�E|�˓����La��1f�.^�L���QQs�ϓ�?q��?���?����O�: �؞;'v�����1D$S��'W��'�6���$�X�\����|�/�j�h�H�K��w26�A��E
I�O�Ul��MK�':���L�<��w�pqC�E�$6YȆ��{6QZaH��n�:�i"�����$�O��$�O��䎩 �.d���҈k�Q�H�8H�j�D�O�˓aӛV��@��ЗO[0YZ�@�ziR���8.��A�O4��'N�7mG榉'���?�B�E�V	2ĉ���VL�!�Q�&D�-I�5:v0�'��"P�,���Q�|R��*C�b�GҖF���u&X�
	��'8��'!���U����4���S�J��@��j#��I�!p^��}@����@}�s�t���,���D�8Gk� ��Я�����I��*(c�s�h�	E�Ni�q��0��� $������f#Һ\Vn�ϓ��d�OZ�d�O"���O��D�|��"�����!�ɘ;W�:\;#'K<S����(<���'j���'�`6=�h�Sƭ� ��Ҭf��qi�VȦ���4���|J�'�?焵H]�Γ���5��;�J�3R�s/"<ϓW#�I��V.!xPurM>�(O^���O��Xva��s}�P�6
�����l�O��$�O����<ѧ�i*T1��'���'��!�M�G�UzD�ٲ2
J�p����y}��l�>��	s≖_}��f�;i21!@B |#�	͟TÑ��vH��W&�Dy�O��ňw.߈4[�B�w�8͛%-�9>w�T��� �'���'���sޭ�6�	5' �pj�E�fX�1Rs�ٟ���4VR�����?��i�ɧ��wT�	ƈ����h"�3sۚm��'\7������ vO�r �t���ILK��*�H�N�E����%(/R�
�j�0a���ՌF�IWy��'�r�'B2�'�.zM�Uqv�I�#\��+FO1K�剕�?i�ٟ���џ�%?��	�H��A�a�F�H��q�_,z�m��O	n�?�O<ͧ����y
$Qt.K(H	@��r�'M4 *%#]5�>�.O9P���lhܘ�b,2�ĺ<i���'����"�ߣ8�J���/�?I���?���j��ͧ���˦m�CHWڟ�[� H����]!E#*#և����1ش���?QvR�9ܴ���iΎ�CV�d�p����r��p�g�ǋy
j�y�'��J�x��d��d��	�?!�ݲZRf�҅( \.|�B�<HZ����T�I�����⟸�	P�'`� �eh�U?v�"�,Z:>�#��?1��NɛFH:���FߦU&�L���$QG޴���~4Q RM]D�	#�M��i#���$��C�'t" �7�`P���^	~�i��D� V��)2�+�*f�iPT�^�?Ա&�P8)�܂fl�O��
1�6{�bus3)#8�ȡ�c�Tf������2	t�����y��a�AmR��!=�8���`N�y��$%,�!!���t�֡S̆2��M�ՇU;�B-Yg�];f�|�pc���Xrx�1lԗ��Ń�M�=�����2�>���X 
�8$�PM�%=Z��:ЌP6`� ��sM0�<�3`@�9���b�P>6����K�?	2X��R�[ L�p��ȇEK����ĕ<��\�q��L MN99��� Eăm1�aQ	U.�+��O����OR����΂�XL�B��r�LF�y������	.t;I�?ͧ	���@�4d�!��ɫsU��R3�is��'�b�
�'Dr�'���O�剜�� ޑ���ݎJfĔ�dAF�>���iSB�'��}����)�� q�(I�$�I�*݋7AC�{�b�n e�����x�	͟@��fy��'0E	"As��cH�4�P$�5C�6�K>��b>�I�t9��M-�����n���@]z�*=�M����?�������.O����O4�侟�@��Y&A!4U��+��[��(V�`Ӫ�O,� �SA�$�'�r�'����$�ЁPkM;h �aP@ �8y��7M�Or�	�m�<y��?�������#ɝ
X�Q2%�E�)i��z}��8D�'y��'	RX��s�-|�����D[Ӗ��jͯl{\�'DR�'>r�|B�'?�iη75�AR)��Qd<y���`�9(2�|��'6�'���)b�1��Q�x�ˁ�N'gA��i%c��]Ǥ�lZΟ��	���&���I���b��u?	G
�d枴���U�c��<B��]m}��'�"�'��ɐ3�ⴖO�Ҿ@Y@@��q�h9��n׏3b!��g�
�D<�d�O��,V����C�'Br(8e��).�
 ��iӖ�$�O�˓bD,��+����O���K�"��%aB�ȾV��xZd�� t <%����͟�Ӓ+�y�S�D��N �	 nۈW�T����2�M�*O>��C��O��D�O��d�h���CNԂj��f��az�t@'���6�'v���O��Ɓ���>|5Iŏ����@�i����7�'G��'�Op��Οh�I�$��EPK#P	�ܨa��+k��)XߴVr��k���I�O�	�6$,F���
:8R��M��-�	ߟ��I�\r���'y��'$�O��K�	�te�QB�r�p����D�<l�OV��OZ��p"jt���'V���噀%�o�͟�,ΰ���|����?q.Ohtжjȶ&�N��d�c��k6���I�� ��	Iy"�'7��'%��)r8*���HУg(.�����>j{��c#mÃ���?����?q,O����O�PY%��<�0oS������i�RqJ��&���Ot���<����5[�ɓBи(g'N�8���b�-T�������֟<�'�3O�%�'�������J9�#(�v`F��ɦ>����?���ă&2p��&>���!Ln���x�J�T#"!K��Mc��?!)O����O��`�O��OB i��[�@�޴��E��5��I��4�?����2T�V9'>��	�?�X�y��T��9�5�B�Lc6��<����?�A�E��?�K~
��!��<J�&X�U�]P>u��lJ��і'�>@���k����O��O���%�V���sb쐐*R�d�>po�jy�(�g�"�;�I&��i�Nc�#N�;�����ڿ�@D�ش����@�i���'RR�O��O��6��������ֿ��\
R�ip\�2�'�b�'C��O?�I��)\�,��x���<Q��#���o��V�'��'��Y�]����I8	wV�X��HN� q�/�7eLyh�y��U�.��b?E��m?-(R��g�#��Qp��>}��l�ȟ�
^F��&5��y��d؉&坘k�xQ��B%"R�T�Qep��c����[yR�'�RE�5j<"�0d�d�j�
��_��	ß���j���?Q� *$�B�7U��Ղ�N�Zc�����'W�ށ�<I���$�O�aj�ë?��"�&D�����Zsqx��Ъt�`���O�㟴�	�,L�-��7-�20�Fp��W� ���SJ���'=�_���ə1T �ORf��=6Y�ԌL1�,-w��x��iw�O\���Or����Y+Z�'�25���Q�jk��6
R��Kߴ�?�����53��p%>a���?��-<,y��䊴`(�Lk�38�7��<I���?i��?)K~������ƒY�������",�@���٦ݔ'hƼ�lb�f��O���O% �5�ia���.�D�c��hG��m���T�I^^H��	����O��I�|n�:�uj��	�Bz�	�$�:K�h6M��;#.0m�ȟ<�����ӿ���|��3���+G#��3r�l�%e��D�8�lZ0����	ӟ�Iǟ��r��O��CF���r�t��mρ(̾��ʦE����ɾ'ٞ�XI<�'�?�(�(�w	�mǲp��@�*5l�$I�i���'�bJǻ	G�P>��I�4�ɿKQ���H����J��h����۴�?)VbZ���T�'�'�dLq7nA�'�-"�#Ty��8�I�>� ����?�*O���O����<9@�/E��,�!P�T�����0F:��x��'e�'1�IΟ��	�Q} ��8Ix|��/�-f��f�!B�|�'XRV� ��!�����Z
[$��5�烙����O����O���?���>�N���$>(�H�E��r4`)��$�X� �I�p��Ty��\�Ef �z ʅ�Ԍ?S�9��
�&^�i1�[⦑����T�'�R�'�ڵ���'��'��i����RP]���Sk�ZDn�����Ijy���F,��<���kC�5�̴��MĬ.�mJC�DZv�	ߟ��'Sfe�v�'V�O��Iɇ�)y�/�>b��_V��P�d2�F�&�MCgU?��I�?�	�O��圡-�y�UoB S�]�V�i=�ɐ|�(��ɼ��'����"�%��E0jH�l,�#�f����C����m���h���?=��� ��ԟ\�'CW�U=��Î�p&���d��M�eu=���O|��|�K~b��r�Z LM���|2���.��i�D�i0b�'�"��*n�7-�O����O����O�� �� hv���QaR:��:��i�^�@�����?����?� Hά2��s�͜?WK�(�"�'6a���'b*(�giӨ�D�O��d�O� �Oe��\.QH{U���KG�1�䦊�.F��Bk�	�p�	���	�D�OVH�wMɗ"�j<����B$�4z�l�?}/�6��O����OX��GR�TZ����;�!����9�:4�`�_�.��I���v����ӟ��I럠�	ȟ8��J���ܴ�hA(4E�Gے5y����:]��� �isr�'�R�'�X�<�X�V瓢)��Aa�bM���
F���ԟ���ݟ���П�ׯ��M����?Q�j�#@��@2�	7�:d9�CZ4���'X��'8�	��Ԓ�dc>�������T	�6��ѶL\"�F��Q$�:�Ms��?A���?!1�,<��'���'���ǎ0.;���:�KF��e��7-�O ʓ�?��P�|�����4���k��G�JCIŒr@0�'@�.�M;���?�d͓�-����'���'�4�O���*m�	z��Ӟ}ev01��.a�l��?�F&���<�g~Zwږ�����>+��T��>sGx��ܴ^8�lQ�i��''��O���'��'H~��H�$,8����!M.R탰arӊ�����O����O4M�O	��'/"�'��P2�H� �H遥%L °4�+oӸ���O���I�P֒�mZ�����֟��I֟֝�.����-��gɢ�%j��]��6�O�˓(�"�S��'c��'��X��U�>%�I�R�� "7(4b�Er���$�Y�m�͟���۟ �I��骟��G���af�1���Gs�r�f�>Q�D��<�+OZ�$�O����O��O#".����?"�ӳJ��/�(���٦e��Ɵ�I͟�1�����?�D�[�(s�sa ]���E�"$ߠK�ؔΓ���Ol��OX�D�OD-<�n�9*88��M��-@cBƓ��$�ܴ�?���?���?!.O��d?4��'!`����O�[cd�q���\⸙n����ğ��I7��I�-m��m��T�I4C��2ɠx��03� ����ܴ�?����?�,O8�ć�YJ���O�����(�0n�ys�$���Z�JO�7-�O��D�O�D�y0�m�����	�X��3�HՒTLT�.��D��
)V����4�?q-OJ�Dx��I5�4���Dl2mb�^�d�Y` Z�M���?�'#�;���'R�'g�D�OIr
�CP-�bb�="0(�"O�:D�|ꓓ?��՞�?����4���Op��1f��*X�޴
@�$l�`qܴ_4
3�i���'P2�O����'n��'R����?Z$Y�u��?|Y�'/p��(r3b�O�O�i+�i�OĀ��O�U#�@�e��Qg0�!&b��A��ӟ4�	Q(Xݴ�?���?����?��Izؓ&D99�Z�j�H 8
lnΟ��')>����	�O �d�Ox����M����&H�.������	�G�B9ڌ}�'�ɧ5���:�@q�F�	v$���i�.����S��$�<����?����D�Wb9����,O'*,���Tx�)��NC��?1K>���?ar"F���HaH.J�c�P���<I���?����"��Χjr9��_�	�ʀK�d	�r>�'�B�'[�'�R�'<�͸0�'��ؓ��\�m �ܪ#�ٜ/zM�6ƴ>)��?����E�.{�4'>�+'b�S���bCѰu#T��-��Mk��䓎?a��@������	�)�tRB�P�3_�����݈|6��Ot�ī<���G�(��O�2�O�taq�<����M"9L�2�$�d�O���E�����n���B_�����<�Z)lXy�؟K��7�B���'���D>?���nȌ*w�]�b��!Q����1�Iٟ�P�����'�b?�#T΀,qD�<ᄟ� ���J`Ә��®\ܦ��I����	�?u�K<	��p~��Ʉ%1Pt�Z�)�=-��iG�i�٩7����8�D�3� *q��A��D�$�F��M����?������c�xR�'|�O(p8�b�+�D(� ʍ�N�ā���i$�'Xԥy �?�I�O��D�OL��w��"H�B�U
P(sq@�֦��I3u�T]�I<1��?9J>���޴;�@C�Q�!��R���'r8����' �Iڟ������'�*�Iׂ�C�Ӕ@��DF�P�"]�s�~O��$�O��O���O�D[��UX���lL"&�}95G�H�1O����O��D�<�s�Iy��	:�ƹ��@P�1tR�p"GM%ԉ'�|b�'B�ЍK� ҅P�ȅ�Ġ� ���!����듅?����?A,O ���D�W��(r���K�FͲ#)�`��γ w�(ٴ�?�N>A��?��ĉ
�?AN��p�N��9��@�ir����� ~Ӹ���O0�J������'h��O܃��h��K%8��{��
<v�Or�d�O�Z��O~�O�S�&P!s�Hc`��ۢF���7��<�BCZ�����~J���b"���1��$]I��1�f���<��dNwӖ��OB�R��O��O��>]s�B��!�h�j�a��R�R�	u�f]n^��},2�'���O�hO6�ą*�rDF�aY4���M�ݴD76�����S�O_b�Бe�\��qOY4T��i`�*A�wsz7m�O����O�)jn�o�i>��O��1�����e�p	����f�i���'"�$��X�d�O���ԫO^�+rϞ+����!v;��oZ���j!-л���|ڏ�dP4*���p�
 a�d��\�V�'�b�
��'��I؟(��۟T�'X��0��W"/�@� M�Q��$���0F~O`��/ړ�?�2� ��R�C�t���W��"�2��!�?���?A���?Y/O���=�H��_(7�8�  *R�)i��W^��n�ן��I�4'���	�`&Ī#��7͇uKX���ȹ��$�4d!%p�O@���O���<���U�H8�O�8�i�)�8��ƴ�hIX'�o���d �d�O���G�^˱O\ ����R��0(7b׳
�n��G�i0�'��	Č��I|���:���2�^9Ҧ��6��L���%1�'�'- x��T?�z4�F��D$B�鑫Z���Dfӄ˓ e��6�iPd�'�?)����ɤ�j|Q �Z9��\�����N�(6m�O���V�x �b?e0�٫�<���ޭ0������2a�O���O��D��r�$�Oʧa��['k��|�J$���"���f�iC�K��=�����U"{��X�0��+���n�=�Ms���?��!�4)/O.˧�?��'���E�1�r�Ǚi��ȡ�!扒�n4ZK|����?Q�`\B�⁈@�׀ ��
�;=jX�"�i>rA
+'gTO���O��d/}r`Y�vm.PC� ƝA�B�"�ON���$ه>s1O��d�O���O��$X;
��4*�e		��iBk;���W-�O����O����OҒO����Od�!ņ�(qs��s)ݔ[�HxC櫍�q������IΟl�	`y��X�B擒]2x0���Z%;Y�L�(�7���?������?��_�.��'ꌠscl���2�����H����O����O���<Y�ȅ R�O��(�d�ÎQbm��`z�ʵp��p���$(��O��d�`z�O�qAiN+���S�L��nC�ivB�'��	17f��L|����A)�yNx5����p���Z+:i�'���'��M��T?2���6��L��呔=�d�fn���}ep���i����?���SL�I �X�J��ز3��HZF��j��6�OT�ă:P��b?�*�	F�0(��Z(�S�p��s&HTצ������I�?i�J<!� .JMG^��T)yuCX-xް�!�ip�b����ܟܢ򊐯tB��k͂=X ��!U��M����?A��=Y��
ƕx��'�O.�R�H�h�K�f�((�������0�1O��O��d�#B�T쪖�]@��R!�64��lZʟ��ɧ�ē�?)�������a�,}�j�v���u���B�D}�օ��'#�'BU��"�/����e��4��!���	*)�&�J<Q���?�L>Y��?�����2��c�&�( Ŵ@ؕL��5����<	��?����?	��'ήp��id��Hw�K��F�A5���&��0��)p��$�OD�D�O<���<�[z^�'>^.�3`%�������AP,ĺ3�iD��'�b�'vR�'��1��c����O� �Q�J0v�t��EA6��ranͦ����,��kyb�'ۂ���U�|pt�2@�<I��/
� қ��'n��']Bi�/��6M�O����O0�)��VT��`	j�@Q�֡$���n�ʟ\�'�B"^����'7�i>7m�,$����ƒ���z��	e���'�B/�+R36��O����O��i�����(_B��̪(@n�5eT5y���'g2�C�!���'�i>���@T�4l�jAz��mɷѨ��2�iP����Fh�T��O����� �i�O���OJ;p ]�'왰PL��R�Xb����a�WB����$���}�S��d���T� Q�>R[�l/K��lZן�����\y����M����?���?9�Ӻ�7��*_�LX9���'Ƞ�+LǦE��Iy����yʟ���O����*WX�9ǯK�TP!�5,Q~�o�в�Ǒ��M����?i���?vY?���k^`�G��'t�l��k�7y��'C���O���O,���OD�d�O�}�B�{Q �	��߲Z��X���^�&$DUmZ��,��ٟP�������<��H���{�n>`�E��.V��I 6E��<)���?)��?aO~§�?q�N[%/�|L�%��7�:i ���6���'���'��'��P�HRWBm�<�`%&�%�Id�(W̐��VR�L�����wy2
�6���?%F�8w ڜ���2*3D��p�����'�R���O��`w��0�UQP闋�B�jD�`�N���O(�d�Orp'��O��$�O�����ƍ�� �;V+͂1�ޑSg��W�	ڟ��'���������&P����n�!S���i!U�4�	�"���ޟx�	џ`�S���'C 9�"��;R�&���Je���5��y� ���O�O�*4�'�G���
V�H�4S�4mb0�xC�i��'�b�O�NO�����]y\(�1DC�jT��rdE�	���������P��cbRPf�%JNt�ĥ�M����?���,)Ƹxc�xr�'8��O�H�C�^	�Ç-�''����%�^#�1O��d�O���PY�t-8	�(�� M�d5\�l��Q�� ��ē�?�������`�\s`��G��7Q�H��W�GR}rP=Ø'�B�'�ϟ�	J."��y���ԸgLXŠTkE�GK!�'�"�'�ʟ�d�<�q
��0�
�� ۙ0&έRi^	v��dC�t~�'2�\�����\��'K+���SMS�{R���R���T�<am���D�	���$�@�'
Jh��T�M�A�<��jP)��=)XA��Q}��'+2U��ɬF�6�?�F�=4�D���T�C�4k���)����' �'R�I9D���Q�'�� V�j�Er6���]Z�6T�"�i)BU���I�@d��?����ꑅ�*����ɞ'ǚd���iv�'O�	�#3�uC�G;�~�cfܙp����M5����'�$Q C`��/�0�!�ڨ5a��H|R�ER�b
lښw�˖G�-�:$EOQ:Jd��r�'��9�G�����#��G�2�-��w$����3�К��A>{ź�)��T��aѢ��S�BTӖ.��^V��c�v��t���%IK~��$� ;N^ �	L��D!rte�F6��"f�Z����0�R/Rcd��!n
Qq��1&> �e Y�3�z ���,���$�Ai�1C�'	��'[R i��I�|R�E�{�f(0�@�,�`��䛲6\��1E�Ș`�p�O:$l�3�u��E�BŔ��h�q����#�͘�qv-P�Ubl9�oMc"�̍�rږ�&�(�탬_��e1ʇ�4��CQ���઴,�O��$>���$l�)�nN�+(	�eM�AJ!���O0�9�e������&�*n'v��e�e���$�'`�I�W�lHߴCZ��g�@�=xZi�!�P	{V4���?���?�d��?Q���$]�y�rx@7��m�v�x��	-�B k3�ՃC�����ʕP��y2-�w�4�������q늁g��}&�݂T����lސЮ�95��W�-HD���!�8���O�)�����ɻ~SΙ�р�D��� �.~�ZxG{���<�0��Ab�7y���8B䉑/��p}�$����R����4�{�4�O�˓{���q�W����Z�T��H������ xӾ���LM7Q1|�4�'�2�'�tȲ�MZ����*�8x�r l�|�fn�in1�qP=)�p�6��_�'æ(���
)^s.��)\�"O\�O�4�qG��(*�`�&�)f��0Ɍ�dΓL�b�'�^Ԫ2.��O�P��'M\�P����8O���,BAƜ��˦��3I=.�����[c≉Uf���e�A
�jA�"��xY��"e�<���O���|j@�R,�?y����m�> ��!�ߢ/�a� �M�9Jc�u6�ℕ!n*�
c>�$��E\)�g�T�?����F�9p�8!'�X�N�=����_=���|u\��d�P��Q��z>�NΙ���NV�0�^�D$Ʊ����O ��#?%?�$������d��JHΪ=��i�`>D���A� N�(4Z&N˨$`U��j=�u���'VlH:� Wd��y�n&!�>5����?�VI�*{�uZ���?9���?I�����v�5;an-\�L�+rY���!�/���d��F��(:J�H���$���	)eX�����/*�ZĲ���#=*�E�S<��H+���.����'�?ŉ�BZ�d��O������<WhDTځf ]`N����O��{�f�O	l�?�M�gy��'��	�1��ʤq�̈Xd�	�P#<Q����O� �AΑI8hk�ǃ?�`�oe�Dm�G��?��Sfy򎒙Qz6͗>y�XQ˗C?G(�� �f�`���O����OH����O��$d>e��Z�Pʤ5n�F�` �bI�Y�%�4�ks��{��}���0I��):,anڕ��<��K��,���3��]�6��Șr��n��B���O��$��I� ���l :6�J�Д�E�TS��$�Oʓ�?�ʟ�́$��1�Z���H� 8f��"On���ND�K�����1G�܀��8O�Ym�����'�`���j� �D�O�ʧ�J��V�\�H��1�1"�@�I�o���?����?�I
d��ە�l���e
����Lv��� �m�4��3@Kܢ<9�c�5l�t�#� ?Q4>��R�+����8�`$ٱ+��"\���g+UQ�P�R��O@!mZ���'�?A���3`�#��9 ���?!���9O�	�	ѳ/ў%�3D��c]���W�'-
O� 
ƌݪ�d��⒨$d�6O(�ǮP�Y�	ɟd�O�H�c��'
b�'��H�1�5awh���!��{R�E%����A�-t֤�sl���'���?����I���z4�σ$��Fo=ʩ�G'p��$���lp�%@]<y�nd�}��YCF�Hum�2A�,z�^�z�C��Q:bnp�N9�����(O6�;�e�:�n�R�À�<���"OZ���D!��u#��[�ܬC��D�O"QDz�~�X�$M����2���>!�Z�$�OؤB�dׂ
dB���O���O>����?Q�>�uڠ(��H��X�	�Z	[�4ywZ%5�Ѵ!
��A��߻����Ze�l����)1��<��	/rP�m�[���f�
W)(��F��Q:���H
x�,�+�)�G�&��Ua�)_���$�<�,��_ۦ5*�t�'�Z��Iӧ�>F)���V Dlq��*D����E��4��`��a+:�0ūǴ�HOdxc�l�O��\<Q����P�Aބq��Q)#�N `��Of�$�O8�d�?F3���OB�9ڴM��<7�`��ěZ�,ҖF�("�(m���¦1Qp�'O�����N�)��Ac��;O�y�uB	�N�.�Zr��%f�x�$�?jBVx��<ړr��X��9�Mj�f��{��L�d�X-� �=P����'��I���?�O��U8W䒡rU��R�A�R~��Ó�hOF�����HJ��8VJն$��M��3O4�m��|�'�1k�KlӠ���Ot�g�? D����#*�pq��٣s^�����>H����O\�D^�~�@�D:~2� ���J*$Q�OՖ����+-��re���X�j��]6L�\h�AG
En	�P�5������奛�f�py�L��Fy�l�!�?���i�H�����(b������X.]�	��7OZ����i�F�8C�(�Tݩe�÷i���6�2">�rU�����G j��1�8>��I9ѥ�F&r�ɗj�����4�?Q���ɘ2_����O��ɉ#���9$L���1;��2])B�y�̄�S� +�M�R">�|
���$NV�Jǌ�A�P]�&E��Z��`@�a��M���Ǎ۾\r �޴>hz ���w��ٳ񧜷<�BTH�c�,�P�#���=�RedӤ�o�㟸F���Z��t/Z`��@y4��#~mNE͓�?i�RyL������\�AB�V�n�Dx"E,ғY�
��JeHX��ַr�ȅ3��ļ�&a��������7�@�����������;^w��'X�١W"B�Qyе5��?1��Z��@Lr�y�&�8F�̐@e8��d�³���<Q񦘏�6٨���,R�jpqWe߇.oH)�L�x��T*-�Eur��'Q��D��>�
:���"0�2e��-H@�8E�ɀc����5|O�}��N�&����[�h�
�O��䇀�X`��&p�Ѡ�B�O���Gz�O-�'I>�x�c`�4da��=�\Y���,�x����OD�$�O���2Lk���O2��-Д���`�\ 1���<ez<��@��-��H0D�ئݪd�#O��@��!�lz�R�ҬR��KR������Y="~�5�R��"�|\	��$ړ�d<�	�����n�(0�x�JH1~?l��d៌��Uy��'��O���L�ڡ΋4�`$��a�)89���$5ړ7�L��gɛuQ�x05JW���L�9����'��ɐU���!�4�?!����	~�0�# O*7\����%�(a�k�O����O�]�)����@�N�zd�w��DW�Ev�7�R"hTz,rV��5�(O����5|.�9T.^�_2:��
�,Y>�Qr'��(+F��5�-Xs��{��ݣ&��kԤ�OH��!���Op��Js>�Q@ǔ7::d�h#$�O��"~Γ`�P��H�4J�ei�/;���'�ў��ēN,jX�T��+jX���L�M���̓d$���iP��'�哔|��t������-��v�0�l͸T�B,j���?���j#b���4r�S�t��'+���"��x� ��>zƹ��"�]�X0qA�{"P�$��O?�dߵWr|��0Oė)Q�Uwm�.M��Ac%��O ��9?%?��IDy�o�4�0|���U<!��L��W��y�BW&��a]`<ˑؤL��}�y��'h"=�'�?с��,\��4.�X�1���?���i^�@�&ߠ�?���?)�Y�S۟���Y'db�5�ϱ�0���@@k�r1�s �
l�>�:a��!D�SG�'���T�3om�`k���s2�31)]�u�����+v�: X�g9��D�I'�B��f ���e�e�[�s����m ��I�d��?��?)*OF����HU�I��˞�0�&�y�"O<���F�@� ��h�&xY
aX�.�A�'�����>z�8᯻6s
�+���+J��� 
�~h�}��?q��?��%��|J����Z�;��0��+8��e�6�:�=+`cQ�l|zy�LP�_W<�3ǝ�8_��Fy���^z��L%)�8
�L�8z=~䃔g�	�U�����z�^��	'H������QZ��ӌ�����:�<*f)E>��`������IRy�'��O�:y;�C���4,����oӉ ~��d=ړr)�${'k��#����OO"T �eϓM�X0���DL�,0���?�����)�?h/D, .��?�>T�����zp���O(���O����O^b�ʧC��{�\�4lM�q!�&c`��Fy"Õ1�蟌@��A-K ��B���^4�剓-���$�O�����X>5�щ�@�h��)�5IW�]���$3�)��<�Fި?��2,:������`�,I<����!J,�S�㋖zl,�Q����<���A�':�F�'�Q>9k���x�	ԟ�+B
'����>t�r��K�Ȓ�[�4H$8���i��}4���R?��|��46�J��l�#_T�u"�"Y~Ls!��'�,���ۙjI"�Q�b�,�h����,;D�$	IK�r���ڄz�Ȳ��'��6�ΦM��\��?���C�T+rA���	�	� ���)�<�����>i�����	hK�:f}~]�GCy�'6#=9GƠ���SNM�=[D�Aud�)zp��O����ɼa6ҁ��ρ؟T�I����	��u��'����>���ML)f^؁�TC���~�%�Z�����4-t�����IE�p���(���SN�6���A(]r��yfʊ�U�d1�㉌w��!2.��&�� ����(p�F��pa��BϦ�*�4��'���'8�b�+ǟ%��ɨ@�-�
��5������,��� ��?g�ͫ�鉚���<��O�+6���V�d����D͝!OLi1#.X�+��'e��'^�ܓ��'�R0�ʡH���=)�5C� <�!��9�4�C!d��X7���:����˓$ð0�4`�Vt�yA4�/8|S�GaaqR�Čv��u��e,��O��Y��'�RXpT�iRan�6��#����'���'5�O�
4�
��W�P>�r��5.\5R�bC�i�c���O���jMd�2�:�')�����%B^L�'�BX>�����z���'�q�6�(ӿ.vQ�	Ο��	�H��A�!f��>��t�!@��?�OEZ�JƄ�)V�h�Ke�Q" �B���D6*�1K7B�!r��m�b]"8��]�`�[1V����%P7u�)���L z�h�P�I�l���O^�?!�!�=i���;�E̮0.����d���I}x��q���Y��	/$t��z�g!�O��&��bč�z��J4S�#�5�~� �$��/����O�ʧ^i�u"��?���,�d��,K�v��y[�G��WǢ�K2D�<�j���Q�-
*���u�g�(��c>��V���@�g� Z����-Y�� �sF��Z���$I��u�N�� �~�Ͳ@��D���m��[�D\�� ؂ ���3��6�p���ǟ��'�?�/OTa�����1�T�.>��!�4"O�0he��<�$���xã�r�1O��D�R�'�Z7m�O�0KQ'UA6\��P�H��`Ӷ��O �]��
����O,�$�O��$�c���?Y �\�j�A��.��f��b�I�-(�����}�ڸui_4aD�'�HO
�ٵ֐f��� *�Br|@Q�ڄd/��C��$<���)u�
#��	"�\~̐�`F =+�%���!��E�0��	ҟx��o����)l�D��(U�M<�{ƃQ�-�!�ҷ�PP�oT�! �d�7͚�ԀDzʟ�˓[@��i���K"��(}�"�9`f'q�d����'���'v������'��	 �Ay�=8dn�%v$�Y�N&f�z �bk�1y�Y@�N����%�'`VM�)�0u�897�	�3;��H�,%�c��ȼJDP0;�'7�0<!ah]ӟ\)ڴ`�HM#�,٧	�n0�!�⢷�� �M+�����ON��$'
��{n�E���J�z����]k�)�B 1V�zlK�϶)��Hϓ|��	_yR���ܪ듛?Q+���� 7�ґ���^²�Y!l��V����O��$�$�h�	�Ό'�	 �O�O���5c��HQ���`~�<Y2�Yyuȹ��B�S�Zb>�rDj8T�hѴf85���C�k0ʓ���	��Ms��i����c"���\b@MZ(Eh���O������P)�9`�m�TBH�pAN�nka|�e;���C�؀0牔,IB"�y�,�R�'��R&�t�2�D�O��'T�����?y��%�(ᦃ�#G,���`�U�o�V=��$�]�3�|*�c>�ĉ�WW�xB��L�Q5�-(�B<�M�a,_Ŵ9�N>E���n.��*�	l^�o�
O���&��>�?��i&���?	F��e.�șbNS�8��`�l�o[��ϓ�?)�MC8h:��ȀVC��a���+}:Gx�J0ғ��I�,���E%*G�q��.Ɍ$4�d�OxB�Y��$�O����O�u�;�?a���IsQ^�^i��Z�KD+@�qQ��'�&��V �%r��s�ƓKF{"��1:�[!T</�xuatdV8$��ę�|~�u�3O[�b)����hOpȇ� sd����MV�b�H����O
�#��'�b�',�O�ʧa,z8�7cU%td�����U���h5\m��.@���GY�����r�'�L�蘧�+�Ζ!��e�D�ۜ]:��� 	O�<�cJ�%�΍Q��Q&�p� M�<�s+_'& ,�c���s:�)�IT�<�Ql^
��İ%��W�$Љ`FP�<�āW!�b	����%�� T+PK�<����! ��@Dg�4�D��+�~�<���W��p��K��X�#�|�<I������k"�	3@Xt�<����eJ�@�
Oa�d�(U�W�<���|\���GCNب�a�{�< ?q� M��O�O)�9�bOz�<��GڃbE� ���
���3���a�<��O
l�L�����>��1f�`�<y2��S_,=��ɽ+��)0 �[�<Y��5w�Yqf(���r��T�<�#�� !l���Pn�Z�6A�x�<a0�X�;�l*�i��r훃�v�<��
��X�ƖN���s���r�<��X(I���M(V���*�n�<� \;`Aڼ <�Dڳ�I�q<���"OL�R��`�й`�]5$�v�a�"OR����-� ���F������"O&�i�.�x@Q�D�L虠t"O,X��M��a�|l��΍:ـ�4"O����jЛi� �1.��R� �9�"OduW�X*�ċs� �8���B�"O�`����'8p��ٗc��4;D"O�ȈfȌ�%t�i:�Ҏ9�&!Y�"O>$�D'��ĥQ�+�j�\)��S���a:��'?੒�%�DL:��I��ˤ!-"bH�@s,�q�x���h؟��AS8�f����O��(��*)z���{R�4}�����P,}x!N	��)�BʠYVĪ1�@5�6��C���#�ɒ
�&���A�Q����eF?9���ʜ.t�@�!+ފ7��s���_)��@�]2�zW��g�^��Bנc��̻jc�(St	�X� �EN��K�M�'h����Y2�\eB�q�(�Ϙ'��퓢D�8f�0���k�,dE���`F�<�ē|�G�2Mc�`�?��"Y1e�REHՎ�u�
�ڄ�آy��Q�!E�m� I����0��y�P��&T���bX�T>"Yi�^�@�v��VC�x��M�� ��@Ӵ��$�C�)�X"�<X��,џO�,��-Y�X�i�'5i�'TCev@"5&��0-x�	P|�'����ĸt>Z°�A q��K���'�ص��� �u*�:B�>j0�92�'�Z��Έc��'Q�'����d�ؤ��0w��9	��\��n=h>�U�<��f(��T��O 3����T`�g��(���(���ʄ���1J�D|���P>d��*Eyܓ4T��Qw�er���4�� ��tԚ�Ssʁ�%��р�$EL�y�x`�>I����]�"�1�`B��ՈD_@��ϕ`�rq�@0\O�TN��(�4a��Ɔ�;�����DЄ��i��I��X<@��~���P��+-m&���4ա�B[�	� u��  �X�⃶&��0{�b��yT>-@
�P��4ۑ��T[�͡�a20�Vu�D�&. ��q�A�I9xa��Ċn��cF��5��<*5!,��6g���K��^CH��u #b��'�H��q(")J`q2c�^��{&߉yd��ݕT�F��3)E���OF?a �|AbŪx1O�\K�b�h�$�$Z��iWeA�n�0��R�R��M��bκ6���.�p=���y�tqC��pL0$����A�"��:A�'�ި���ģ@@�9��] ������'S�c�&�%��Ez�N�:h�(X�r���BL?� ��f�@��a�/�42���� �p�-"
�j�4�0���L���4,S̓~��0$3"!�r�ZN+��j3fʨÐ�B��8��3��9x�
ƄÎv㦍4I$�qO� �S*�<-�t����էu�VEe�y%r���Eם"H\���O,>���OvT�Fj�Jg���2BX�_����oW%-$�̢p��o��D��ɕQ����ݖ �(� fb��d��]�<A�b��`���>���̺&�va��Gf#ֵ��@�RW�'����dԚV�	�[�*����H��F����:��;�p���9���m���ێSm����'需X�l�+.�T��k�k}�4q� ;?����qV�mi�$QP�6͋�%������dY�c�THY2*�ez���4F�j�'�����'�(��hwĈ*i�F不��)d���+u)T(�`L6L�Q�<d�6-U*	�*������ą!4�g?A�L<U�!j$řC�l���V���Q�c�Ҝ���iޙZj�� h{#�[�K'�YFL��u �ɗp^�񴄉D�s��󰌙�|�\�`L0���/9~����^��k��}<|ɫ���(n̛6��Rrǃ�r]�55얛+�b��i�e��x2�40MB���Z�@�u�'+V1?٦������e#bE&z(�	2+����B��tP�(�i�V� �m@�|�'Yҕ��_��t���KN��H�a�'1襩�@֍<1�4yЂ�Z6Ҕ��O���$��a��� _[LiI��U�f����$'ΡE���̈́�_Z%(b玪��X0��?��E�&~�$?O��^�FJd�ٱ�NIc\c�&��X�i�LF�]��Ұ�Tr���A�i�������#�_x?�`&DްL~���eQ�~?%>y��L��%�}�IM�V����g*��Z4��an�:��D{R�E�" ���f�&M�b��d�&1��d�BB�(2�Չ���1tx��7�>�'���~��J4+L0Eʦk]�<�<�E�W;>�e�F�Y��H�pB�|F�Q(�@�7���3b ��1ֆR!FҼ�b�R(7$F��|����¹'*[,P~
�R�'�&7rڡb��GΟ�Be��A��M0��F�x�#"K�
��;ymP�shT�U��/I� �3&d�Lk�9�JM0EL���W���`ट��K���f�:%���=:��QPl0H�A�ϱ]�ځ�'k]=AM&!�0�3p�����w�&(C����,��[����Tm�"D?����8P�韐��6M��FC�MB�,v�:c4��g%K�ش�� e��#=yC�q�Pѱ���(4��d�f�Ҧmb���C���2�D� </Z�Q�j��8V	�:g4��]�1�m`���#`�q"H�\�ڤW�O�iV���pm���L%k�Q��Y��ʀc�'��)[��=��5)�̵>)UKѨ �xIq6�Aa�? v`�&�D3����j� T�,��Eo6_�2�H0��+�fB���t�a��d 
���d޵P*V����]0v�Ѣ�CЉ��\	�O����79�Όa4�<��.��g^�D���@ǾP�ʙ���>��$J�h��t��4����SD�%�v�Ѵ�ŧ�8d��fW)���m_m;�|�I=��T��$�B9n���W�ەGǤHp!RX��T� pTax"M�+9Z���"��:�����ڃ#� 2�L�0�Z0����	J�8�e� b�JdIU��:��=����Z�,b2�T�TE�����3i�9�a�wS�i����_WX����i��١�O��@���fѹc�_�H[b�Џ�w��7lQ��A��d���P�],0�D �%Bn��I�4v�+��S"f�@�]�{	a#��P��Ot��o\+#��8��@�&wlM�I��~~ƴ0f��*�Čbv��4+��	��cDCf�T?E�'��t3b�+eڈ�`��unj�C�!^7p��M�֮�8M�ay�w�{q�T .Oĵ��
]=/w����F�7'���@T��~��L�?�&?Y��M�}½"�ƛ:�rȘ���O0E�	�~�'j8��%k#�8=�ET{���Q�[2��a��
4��$I`��ee�!+Sf�.@A�B��yZ�D��+Rb�.AC�R�d�~IT����б�RY�DAqVf���C2]���.�;0j1� ��)�l�Z��O��4[$�@4��O0��-�!,"<,T\a;s�K�>Ub-�%$28��s��e�WMz^�a�*ң�1O�,B��7u������<Tl�3��$��pQ���L�dB�%P�Lϧ]�(Z��1q☨��Y->Pz<�͛�%ܰR�/����F~��i��ITf�/Ha��y�(�c��m2����C�e۴'P�M���l��PY�PKԫ^"+7������%&���Ȇ�J�uX��d1ޛͅ�:��I�*�6 ��R5����$)��L6R�p��.��t[�"Bň~@�Eq����jU6������)�ƖE��o�m�b&X�}��}*�FQ�j��aDzlގq��h���v�� JB�L$�?Y��̃Fp�(�g�d$�E  dή1q�j�����'H���mb��1@#���Re�D[����HY��#�G	c��,ϓT� d�V���A2�wg��*@JAR6/ʈX��Ms���O%=�z\���d�֍�)ʨO4�O�XV�p���TN�&�@1R�Mm��B�Ÿ��=A��� ���u��m� ��1��4x ������_�ܱN<�go
$T�ЌoZ�G2�!���̾x�l�J�'F�6���J��p0�<8C�Oq��0x�"�h�by�ƙx"Ô�b�>8Ж#]����j�`���?)��!)���+`���&���� ˄�"T>9Ҋ��h��\���ӬsՒ��.�X��@�2��5I�8�8S%ɜ|a"ъI�p$���Zf��!�KV?pF�l��
 [� ��an�<";d��Ă�Q}Ȉ�f%��	��`c3h��`�,�я�*�"�$�V��/�d�]A��*^�b	p�H��3쟿h!���䏟(��)��酭l#���f�ğA�B�`u�7I���c��'Zld�e�צ��!�*'q�p�O<Y�'�L#:湁�IӺz8����	�e,�D��1]s���a�)y�Vqf�OBZQ#!G C�<�ل"S�x%�E!�U�U�hqJ����dD�	NL����x��ɸVOƒz��6�ҩ	�Q3GYW���GǪ�>���g~����Q)�E�qY5�N�jx����WPE�MA��p?i�M��S�l��G���Ma0#�vQx!F�50xE�O�(ppB-�4�ѬH��.H�Ud:D�DP�
��Q��*݄_a}�%E�I��K����@���ST�׿_$�Q�AKG�"Ě���V���b���.��F��� ����Ɲ��p�YwU��d���ӆ��C���V�ʊG;��Dz�%��h�D؁#�ii�mԁYX`^w�����M�plɳ��N
v<a��=0�e[��|+���h�3f��D}2#43׊u1�B4o�z����O��?1w�H7#� E�b��*;;�eK�+	wߚ�=}�/Z�YA���(B�v	x�㒲f��8*$�� "ui#D(�OH8�"
#G��sCA�0�vm�P���U��2�.����?Ec��|�cç"$��r�J�~@��c,D5k�NARC�W��0=1���<!�ôj`��S�Er�\�q�E3W>�����Cw~�B�&.|��i]��{U����'G���ܲ�����." ν�F�0d@1Oμ�N�O�,y�O!��� ���ӘS�ݫ��g��4�U��.�h�[4�ޝ
x��y�%LeP�붇f>#>i1�Hw�b|SXq��9���hZ���X_��FA	�O�d1�+�?˓F�&�����gц}���*J�ʕ����O��ye�g���jd�AQe��h��D&$����Ȳ(¾�d$p4Y�<��h�Ӥd�8����Hs��Y���)E��,�Tኟ:�����	�-�P隿zk��0O�Sơ��*T��(2Q�8g�z�;�'!�7m� ���ɞ�Ơ�ֲi� ,એ30N����ekȄKG��#2ٓ��A�fq%�ۗ��6tfp[��\�4�h9 (�<�Am�8vazիU��is��� JWa�"a�5�'U80�2O[H�tT�#�Szԩ��d!S_�i�".�$W�l��a��Z�0�͎lb�Mp��Fj~��)�qO��)ȫo�؀k�>�>@y��.���������>�1h un�.���
��D1G$���I�A;�I���BB��%�&`,�tP���1?����	?tQ���(��{�/N	e�A��L"&�̄x�j�:�1�O���O$�{ɗ�r	�7-��~��4�i�ȒV��6'�֩{�#��~/���g�*扙>����c��)�mq�c��g�bb���r�{�b$�OG	oi�,�ʬ���+�7=�JyKgl	���h�� �S�? ���oÄ%�����j���� ����6MZ6��?-,Vx�'r�fjB�9˦\Q���J��QHV�_&&Ś�d�5_az�+�-�r��b*������'��-��=�U�%�~"���I#��x��|R�.&2�5၆)�����݅���R��A�'H��i�\J�g�*!aL0���&`$��p��!5B(m`�'��3|bĥO��OH��`��Q��$_7��Ŋ�'��A#�L�	&4��D)�^�]S�'�\@p!���pBsMP6u� �
�)M}*P�b�gӮ(�"
�?˶�	��a���S$kϕ����/`	��$�Y��E��ο%[�D{�*ԃ��m_ �x�i��Z(�?Y�/��F��M\	a�E�G���&(���ӺT��T|&5�mL}��ljňB�"�9I�oB��p=��IxFR���n�� 1L��2*��b��AB��h�ެ(��1�V����(0����u�jܗU��4�/�k�/ϬM�0�E^�z�9%Eׇ!=Q���q�ۆ��D��Kj��I*�6I��"Z�Lk��1@k֦)����g�$�M˓a]�y�h��0��v��**P�L�@�X�S=ȼ	���^��'�
����,?I��
0���p�!GۈL�jsCI��<�8F�^� ����Oʦv���h�r�@ld��E�n!KF�`��E{�P���fA��1�|�j���Y�j��EHM�Qٵ"O�T�s'R�uY.M���
�yj�@"O�ꇩ�2]V�@���Pf@�"O�M�1�D+U]���7#Dd�!@&"O��*�dصh���BA�9x]F��"O�|q��h��f�"tT�Z�"O�ةe��;��@�!��  B�� "O�t�6l�q� l�!��<Gڜ�`b"OX4x���< ���CJ��x����"O(<�+�{�����iD�F�,�A1"O���+\�&�ڲf�NMbe��"Ox|����^00X��/�#,�z1�U"O���2��/��%�U�d�X5Js"O�����.3�M3S�]I�}�B"O��C&NY�f�����T6���0"Ot�Aj<ӎ�PB	@%��S"O��{��Ow�À��E�8�"O��ks��C���mH�G���؀"O���K�*����B!��ԂR"O�a�F�g���Sf��F�<}�"O����2H���mK.C��5"O����+��!�lU�t���"O�QJSI�"t���1,J�?�xC%"Ozx t'O T+�E��j@*F�~�k�"O����hZ
h4�PUC���]� "O������5��4�pA^��(H�"O��v��	J�T��q�M�<���2"O�H��$�7ME�=K�Í1��*�"O���)GB���A�:i\�d"O�%
�ʑ�"-��`���! ���G"OF�"�b=Z��a�T�SxA�"O��@^"1���k��( ���[�"OXly# ���H@�#��N2YP&"OxDPu��Se��j�"G�\��;�"O�HXg̑�z(��Y0b�:-<<�yw"O�ɔ*D�wen�ؤ@� (lȪ�"O��6��+��<r�F�|�p�d"O�!�&�2!)�Л0���&��"O���E�� 8�f�y�#�N�u�&"O>I�7�"�S�Tn$8h�P"OmZ`��O��j6�
7���ȶ"O`�Pd`]	/g�9�w��/l��x��"OH�g��%�6�	�f� �pc�"O:�bD/�xT@�$D}�ؕx�"Ot���LM!-�>ER��ֵ���B"O��*ŎM�-�D��B�
oX(E{�"O����oZ!:���V��|E�u2t"OH1[��1��S"P����ZF"O��D"��)���
�C��Z�Pb"O� �`!���b����`��z�0uz"O�ɚ��W:V`��Ji��"OZy�f�4b邁�ը^���s"OrՂ$�6h��8GkK�!�J0�"O�ٛ��OL��2S�ރ|P���b"O��AA��r3��i%��a8��sG"O�s���w���2�>FD	8�"O��Ҡ�C��ѠG\�8;��"O,%�'I=z�<�Aƌ-WG�lpw"O�8�e��!��@�b�:KFHey�"Op1Z�B�'e�:�Q�%�11:ژ��"O¡P�?�ެ�E��W3Z�
"OX�B�M�$$���dh���"O~*�K�W�6�j�>\��"O�T�5dI*�< �(^�%�x��5"O��h4d\�Y� ³(�F�^u��"O���PH�,�8a4��'�-JG"O���r-ƎD�^8k�N("��s�"O<t֨�9~=�G�V=�x�h�"OlI���q<�ؗi��I�(|!�"Oj4q�B��[S	���2�a��3LO��`�h	ZQ(��Ѥ<�:�a�"Ofu��U.>~p\�F�'���P�x��)�S�:pD}$fB�d:��@�
�Ŏ��$e�܋rOP�h9���1C��l
�M&D��Y��޸G`�t��웈H��T��O/D��b��Zr�V��R� ����+D���
ƦnnTr��!m��c�M?D��p�Ɇ�}��A�bI ��)� �qO���?Z$�b���K:���l�w�!��u(z�j`!צItC��\ �a�O2l �!�hH�XB@�1*I�@�<O��hO�O�8� �	0RZ�'	��*����Ĉ&C:����⍻Q����AN�sD!���O�굪r��M|��ӯV}�!�D 851$���R�_nH�0/��y�!��� 4�N��#)�9.j1�U.F(M�!�\�>�hT�v����+V,N�P�!�K�f4I�Nƞ+̅ʃ+\�h�!��U�H>��d���dB���69�!�� �L�Z竃2��2�9Y!�$T�-6(�cB̙y;�a�oI!�DL9H�XɁcl\~��`�T#�ea!�M
j�4��6�֠��ⅣNMў��<	H~�⯑c}����DϰV����g�P�<�pܰM��Ӄa��M>2��KLc�<)F�oߖ�k�� /Dː�W^�<��I6h��C�ˋw�t��!c�[�<IW��ET��X�އy��Q�*�l�<�&�L�\���#FP�PI�)�i�<�eE�9>��6n=dz4-�f}�<�D؝P�@��B:g�l��D�w�<A�B�Jn6Ջ� Z�A�@$jq�s�<!�X?G�@�!��P�3���c��H�<����	~:�X#��+."�тa�O�Q���Oa��Ѳ�˩8�hl��!�!1��	�'�&j5��<�fm5�õ'�B\�H�h��	L���C�,\/����B��ƓO|����3���إ��  �r�� �$dHC䉤gA|�����#�a�kC�EHC�	���a.Sz��胂@c�C�	�;Dl�fJ���$�sV��a�B�I��0zs�V
�!����B�	-d��X�e��:�8��[l�C�)� . �f�@�J�S�G�Q�� "OHM��A�-��`&ʘ(B�bP� "O"ѫ��פ�|1`/	m6\���"O���O��U�Q!.�DI�My�"O6E�&�b��lI�x9`�2c"O�aI����I2�{�,�*�d���"O�p���j QP���9r�Z�q1"O���ԝ/Y��&�A�(�'"O,J&5$4�6�Q�
D��"Ox8[�N s�@z�d�.'��X`"O��10h�� 4�pm�#
�d`"O4U�2�� F�4�����P���)\O��$��hYT��:ˤ%Ӗ"O�ث��Q��\�AIҢ	�"_����.4�(���o��RS��&W$C��=? �0���RԲ�[��4 Y�B�ɪ^������! ������pu�B�I�*�<��c��2����0��V��"?����J0>��Rd�
'�8���'[00V�d8�O,T�C�Rxd`����XK���b"OL+����
٪!�� :8�|�"O�p�"@�|>�x�ť�4p�E���^��sܧr��U�$��4(�4!U�
�D=���ȓT�)��NL�kf�!�qAK%TȆ�b/$-I��
Fx9��B�� �ȓ5�iAb�AS�F<x��R�RJ��ȓJb8K%a3i���D���!�=1�y�?��'. ,z�(�#K���0Δ�v�ZxJ�'�v��s�ץP,0��-Ù?i~	H�'?jR��� �3=�l�p	�'���s��)��x�%h�+e	��'~9��#2�Dy���-Us�9��'+��q��
5Uv�����z�vD��'s�����F�s:��@!��
��]���3�S���E�k�^U Qiz[�S!�Z��y���I>LIY�b�_~��� �Q��y ��F��z��,� �SU��$�yRm��_b$u*��vUHH���y2)J;(�X�T�_H��P��	>�y�c�b�tq��<\�јC"O��y�R0	���s�늴MC��(#,O�y2�D,p����̂=%�@Hb�C��yBJ'm���Ȳl͓4*�졑 L=�yrl˫H*mµ�@�3�RYA�K��y2��+1�~��1)��$��!���[$�yB�(S��!�.�0oV�!��O8��Ak�TҶ�,@�K�2D���_�<Y��8}�Y���7Qb�2,
X�<�S՗�и��,-��c	�m�<��p9z�jeZ*x��HۄeD_�<�5hx�y�j�(]1�����U�<��f�<\��E��f��27$�"��N�<rK@�GӾ��i���	D�Er��G{R��>��4���6��H�'M�d�
�'I8�*t�>.�$؋� ����
�'�����ƌ�0����1bX	
�'Ė��eA�G4 ��D� ~7�p	�'�����(N�|F����^�{Nhs	��?)�i�cEH!�F�/�i⧁���y�E�(f���)I�wvDx'�=��OV"~"�m�A�viB��F
F2}C��Wi�<�M��µ�҃C`�L+W��d�<y���0���x�ą6X�=��E�]�<���[?" ��2i�Aʔ�I�C_`�<� ��x�F�	�9��*� <]B��D"O��٠�|
�'�=uT<�"Ot5A��)ZS�L�=F����"O�3"O/!A���U����8�"O@PQ7�K�R�0�z���+%�@�S"O��iJ�Q�Dd
���<3�BI��"OV� �c7���L�
�x���"O�a���سl�� ���߰T".8�"O�|[Ң	��ik�i�]�ԑ"O��@��2]���0�H�
�C�"O�����?�|�ʂM.�t"D"O|����G� ���e��~#~�"O<�1�R 1�=ꀥ��h0:\h�"O����^<6��ۃ'� �"O�;A���5�D���
h��	��"O���͞<�@��wc�=o��+�"OdX��ȉt���"�vM ��""O����Q�z��S��KB���A"OD�PK���۴�<I��4�"O^�З���:��ՍL��hR�"OVq؆���JC`�ѕ?���Pd"Oʌ��#щi���:o�8Mhۡ"O� [�J�;DMX�(p�g"O�s��C�i�l�08��`["Or���E�5��u��*�/���i0"O�=)�'"�)y%ꇐ)��	(&"OX�"�hUR��8�ĂE�q,"��"OR�1�J�v��z��qNys0"ONT#�*�ilE�F�X7!h��"OP(4� Q�T��oS�[l�:�"O� XV'B�I��q �C�n�Ty��"O���u�� bP
a�
�����"OԸ۳���kgj�s��02LL�"O�q2J�\���Ð<.�AQ"O��rv�GN�d���%�v5�D"O���GL@.D2���@�bR�8A�"O@�B�O>m���6X����"O��Q�B��sh����H�A 	�"O�e9�j�5E�ؔ�u�ѬT��"O4�� �3ذK� �2c*��"O�)����G��{�M�-�t"O�����S"̑I2��2w �4"O ��hR�\�� ���^0{4"O���j6`���h�42�e�2"O̬�gk�
@:d�#'��A�Uð"O0 FA6cw2D+A�%gj�`Q"OR��`m�(**:C���\����"Ox%�2-ۯ@�d+����\���?D�8ňǚNٌ�� v�P'<D�,��O��R�O�m�t̛�(D�@�dKC�)*�s�瘥h9��_!�d�q�t�+6m˶	�q�"䘪!C!򤅋U�"x��J�#-TT�!ڲ)!��,] �D\.+t��$!�7Vd���R�h��D�֣\}!��ӏlk���?W�a��T!7l!�dӅL�^��U�O�:Ԯ��PUE�!�)H6�IHC"c�28�񠍭U�!��k~��"OV�C_�e��`�_!���B���0읎}����e@�u�!�䌊X#z]�5�)hv6�u��&=�!�߮E9Dea�(W*o���ԫ��!�+��\���Q�:S�p
Q�!�d<r�h�cpcǈ?+z��0	�>4�!�� �9ç�����IA�f�,��p[e"O���!�3P ��oB~�<A(�"O��ж�6�[�EN�X��M�7"O�`��>����i�����"O�kd�Ф:JՂ��h�K5"O0��b��b>�����	��y`q"OB'�x�PP2�@8"O<qJ$��iPB�[SGΑ:��r�"O�`a��]�'㜅�fZ<I���"O�\K��������B�H�����"O:�����	t�H)�D�$gy�Q�"O�������q!4(��<^X�"O��+@�F������6K[����"O��2g*�0!�Fe�(��e"O���l�7^�&���i3j�0�"O���O���yXR+6`�"O����ל�Ztq�*^�w���1�"Od��A`S�?X���"�$/���e*O���Y��<S �U�Ri��j!D�t��M�d�����)�#�� "f3D�Љ�ڻFg��GiA0�(�1#�2D�P����(J��=8�bE��8��e)-D�H�gg��(�I��$�CSh6D��Y��`��XQD<�d)� O4D�\(E})%���߫zf$�p�6D�Dz'	֚�J��aF�v6����)D�����Y��@�zv��W^:9�"�(D��Z���"<��q�0��oܾh��`&D�@�-�2jx���ڜe�Ј���!D����=f1����)^��+ *O0Y����mٶ��������!"Oi�����P~$�Pc��+o��Њ"O� ��!�-�(`��d_g�����"O�|�/״T�<h"��+nމKv"Oڈ���[��9��C�hl�E�w"OZ�q�A�UG�#�!L�
1���y��ֵՌ��� R6ر��H��y���=u���7�� #� p.��yRFV7�`Ub��Q�������y�G�~-6%{��� � !A����ybO��Z��������e�#a�	�y eBf�C�W�N4S�$H �ya�6GM�H��οu��d�I&�y"�?I����� T>l����&J�y���T�䒄�C�;�n*�C4�y�����1Y��>����R��y��ŷ[�"�j����4��pW� ��yB��(N��}�#��vr�y:P�3�yb��������k*�0*0�N�yҧ�o1�(j��H�]��9�T��y�N��ڥP��)%��i���
�y2	T�a4 ]��D�!N���b�y���n�x�2&b�	$�ecRJ��y����0 ��Ћ���0s����y����S�递�-2��ce��y�B�.nj4���
����!���y��3 W2]�bN�6�~D�PK�y"��/Z��ڠL�x����'�B�y���4���.E[�5:7F��y2f6ICXDK$��Dݪ����.�y��hj<����5���E�ߧ�yj�3Fg>�c��
1�����9�y�-3�X`��]�iBA��y�c�C�4bR$,*�T]��'��y
� p�q4��h��
�0[�Jh��"O�I�#&EDⶈ�;pƞ\;b"O	��(��"&T�����LN����"O��b
i��0ᕋ�/[H�9�"O찘�:�
l"f
�Yb��J�"Oڝ�C��&B�4��c��kP�<��"Ob�"��M�X��J&1:�h{5"Op1H��ڧu:�z +�$ |=�"O��`$)]2?8��hJ
'Jf�k�"O�py茜<ڊ|� +N�6���"O"���H��"�h��N�u�a"O
�Cvl��4�Z�� ��$B\ "OTؠ�ϩB<F�:��@�Y�	�"O����(0b���{fOç#T(�"O�����&~O��� ,B�4����P"O2UR���fw���)p�""Op�r�-h�$R��Q�k���"O��&
L�����+���8"O�s��Q�dVT��� }��H9�"O� F�T,SKv|�s��_10� "O�$��&Z�D���å?}&J��!"O��qE��i=��A@�@�}lH�8d"O}��JR�*���Kc�[�c��"O�1J���/`1qw-�%1�<p�"O��ȑ�# �n����
���"O:�0ӬM1Z�@aK�K��jJ	9�"Ov�W�%	�lU�P�[P����y�$[sD4}��a
�R"0 JeL�-�y���m�T�yp�Y�=a4H��y�aؓ���z󪩒c�Ŗ�y�&��g�,;��֚����Ɨ�y�㖆�~5�B:f,�1#D��yb'P-�%�4CҤZ{<l�!�K*�yr΀�st����Ь	�<��	�y҈ѿ! ���� 3qD� S�&��y2D�$m��mz#�	�g�49��ǚ�yb�O�yO�Ջ�$�>s�j�Xa��y�l���aH��l�f����&�y���.DR��7�΍:_<��A��y��xq�e�67���ϓ��y�w�����υ0�H�4c�;�yr�S"�f�c���:D�	�yBaN;���2Ό_���j��O"�y���y{Pa� #�n�ãO��y&Ԙp`*P�0o�8�|[�,���y�o\�Ql�}��MN�W�zq�9�yb��(�:�:6jU�����P�y2o/v ��`@��>I�%�# ՠ�y�V('�x�k�3� X�̦�y2�bT){D!L,p�����y2�U�_yX��g�C�"�T)B*��y�g]tqx�X��ȗ	)R�pP
�$�y��\y[�բ�dy	� �y"lá~����`M�~#$�G�-�y��Ƨ,��$����v0Ό�6+��yr�u�&�BR�l,��#Ǘ �y�M�->7Ni��Ib�i;�/���y�
�4"�l�5�ӈ�4Sj�B��4!'l�x�_�TٱD+H>Yo�C䉒Ip��r$�l�����(���"O�q�b�?k4��6���w��
�"O��;3a�>HD �v�<l��]"`"O�t+�q�܂d�ަyʴ�G"O�ԸBB�Ko����X�,F`��"O� JUZ�GJ>]�b1��KA�i"��zG"O��:�O�=��͠�	�:A�X��"O4�{�� ���Y����L$�|8�"O���b�պ2� 
��
	6��z"O0<���<�P4��L;~A��1"O���a��7[Xt�cdNQ��;�"O ��cC�5/�PA��P?U�"+C"O|�̕ ��[aiͺ�^"O���C�
\��P�P'@�c�X@R�"O�Q�#�ߖL���(6���n���r�"O*i��i�H���O�X�8�(A"O�d�d��:�����Ƈ����"O�"c�óCа[@���4�g"O\�"B+Z��b�>�,�0"O�4#e��BJ@�9�'�?1��U"O��R�)W8D� e FL��2���"O49�bd�U�h,bхU&�U��"O�dj��ŏ.�|�B�e��6�UX7"O��:s��8��<1�����4��"O��AǍE�l~���5��/d�&�#�"O�=�G���NQ%��0B<d��"Ot՛��}RHh���ȧ	��Hu"OLd*�iz�
A�w���a�œC"ONtz��S�F�)q���a6TC�"O�%��.9ut���U���|B�"Ol,�`"��4)dI�DL�&u��pB"OZI2�XҬq�"�5I�2���"O�d�v�P��H�aO�����"OP��A /qf>�`GB�b��`pc"O�|;��3
�mX�R2SЌ��t"O�ȓ���4� ��#�7��-�B"O`��aa�`w�q`Eϙ�)�T��f"O��ck��.Sf�0˻�f�H�"Ob�#I�)ZhP�0n�7�H�"O�y�BZ�&g	[c�-*z���w"O�xD�?51�5�k�Ke�,�0"O*��d
���Y2cϐ^IJ��"O�H�0�Vc� PG*H��"OP����ڻN��(����6 ̄ir"OFE����Š@ˣB#%.Ţ�"O.���	�G�ny�e!мN؜I�"O�����B>�c$�M�f,�#"OЀ;T#��qrN�v��+���g"O�*�	��:��3"�x��	�"Oz�ĤȚ|.ht�D��L, �T"O���Q���x��V�U�:EA3"O��p�O}��$A�2!轰P"Oxy�1.�/�z}C�O��_��0�"O�x;�Ə!�n}��J*A	��)"OfA��
N;d<�������舴"Org���>��C�L���"O��i���V/)�g���|l���"O6D�c@-ހ�1�[< >�ȧ"O�Y�HЃow*4��B|�8�p"O�� fE�%Aa9�H��Lߖ�B"O�=Ȇ@�.X�^�
 *E�VŎQg"Oz�Z���
�Hђ�H�3%U8��"O�X� ڷ^�zy�ᇶfM�y0�"O�,��
?v�P���96�*5��"O$H��C*��ԃ��2���"v"O���JC7b�vhے�@>k�����"O���j�z�
�00%H!E����E"O�[��Bk��A�E�+v�d"O�h�Tf�@ ��3w H�e.���"O� �Lk��O7+��囶�֘�虪�"O�E�

 �9�-�|��s�"OR�3�+h<Y���2X�:eKu*Oeyf�NS�t��E?�q�'N�1��^ I1�ˑ�/��J�'�4�����M�v�H���3+f���'F�e9S�V�.-��`�K�z� m�	�'�y�����,�`PP�ᅿk �=
�'�5���:c9�s nT�i��`�	�'2&��&�<hK2y(�Z a;�U
�'��%��kG$E�~%##"	l���Q�'ڠ�BU�Ku�:�C��Zc��D0�'�t����7V�n18���]6�T��'���a�Y�)�¡�'Ǎ)"spԲ	�'�.M�� ȯ8~pz��OD�Y��'�9�.�Y,���
��d4��r�'y�p�A�ʾ��yv��p	��'Q6XA#$����yE"ҡw�����'�n8�ǎ�v�m�T�9:��|��'��,�ׂ\���
���@"O@U���=�LĈ �Y�E�޼��"OX��gC�8�8�2���$���"O����[@�x&X�$�.0K�"O:��#�R%�����H�i| �)�"O���whɅ3����w�
�rL�U"O�+pB��T͛t���"O!ʵ#i��a��5ۖ}h"O ջw�$j^�i�L�%8�|��"O�'_=��)�G)�/����"O��`�Ʈ5m�r�n�2/�*=[�"O ��2g;C�͘��\;r����!"O�`a@�K�t������=���"O��gM��k�������""O<�¤��?I^�! �cw��G"Oh�z�HR�4���O��Ja�AY�"O�	�1*܂m�8�3�/2ȝ�1"O�R3�[$@��Q�6T���ʲ"O~�JF��@)�IQ��;!x�S�"OZ(��N\�t~�}q��� �ޡ��"OE��I�Aq���0��,Uz�Ix "O]"An�pQzy��.
�7p���"O�ዕ�N��)fMÚn�-A�"O��c��U/K�ШU�ݴU`�@�"O@�9�G�a�0dB��I�0�"O�ڑ T2u;
e;�ɂ'&7�;S"O�8�jH�O*6<J��,\�:ɒ"O:THaC�-�������&�&��f"O�`O�8�]2(�-3|�""O�p;2�$��u�p�3x&���"O�٫���'7����ڣ>u|�z@"O+�[�jޮ<��	vY����r�<���O<Il.���C">����� ��E{��)�，C�Z3wJ�L���geC�	�o[�`�6�K hHq�k�m�B�I,C�5��j/��(C��M-�C�I�)р�5��!7�����\��B�Ir���9[������CS�B�	uTJA ��.|ol��0bٺ	pC��&3_Du���^5m�2����*9NC�	���de�����]��ԱZ��C䉧dn����
�^v�Q��K��4�pC�	`(q��&�-�Ƶ����]�:C�G�|��k�,YV0*@���C�ɍ|�2�XхҕjK& ��n�� ��B�)� ��%,*����o��7��m1�"O���g@.9�����ނ:�����"O�|���F�?�2ԥ��~j��R"O�4�!�6 ꐧ�<*m.�yG"O��Ku㔎�nQ8P���j��I"O��1$��Z´�"1f5�L첕"O��0��آR�����nU�UԚ0"O2�9@�Fo� PGkLW�zT�3"O(���`�>�I��85��t�C�	v�`��� >Vy�"�
�����:D�Xd�Z%jcfxS� �<�59��:D��M����T 	o@��@��5D�qbd݀H�pA�s덒��L3��4D���7�]�;�~�)&�ʏ}����&D�ȡ��Ĝr��8���;
|�s7�%D��JWAüs㠌k��R�6��5�!D�8z�ɀ>5�� %��UJSg>D�h��G��Bǋ�ɤ���&D��Q �:qi@J���l0�|�$@ D������5X8�$��l�>�aae>D�`�$��=`��vF�(F(�A!�
;D����	�'�4�3`e�jL��&.D�D
�	^1Ŕ� %H�ER*�$�)D�8YW�_�"�2ŋ�1c<�ZǍ3D��k��ߜ
�b��P?vn����A&D����'wX�K�MK�.���4�"D����/��8v�֡�mЊ)�5�+D�bG��w���suʺB�L�o+D�����P0��50����-�xD�a*D�h�D\(h�B<xD�A�fBxH�On�=E�.͔*lr`A�+�L�0G�^<N>!�d�0W��yZ��:!b�M�>
!�[LtM�S̓=r��ha�X^!��ɫ/K�qj��m������"�!�$X1qk<�B�G�-e��2N^�!��?βE��k6D�8ر1.� q�!�am���MQ$����u,��d�!�D2NV�ܒ !�,7�J�8q��#ru!�FD9��,E$b����+*gm!�䜁#&>�yH�3��Id�/U!�T#(�0)�ᄼ=۾A!���? 6!��|V��fʆ�~�� #�=N!�Č�6��@9��؂G��q1!�$MG����g�+��� �M]� !!��[Ϊ�JnN���Kߤ1!�d�6z�.}Fd��T���e� �]�!�d��{A�P���9Cr(5�#�!�$��ce�� �B-`��h�H�!�d f�,40�f�,�1�0E�s�!�d߰W�B�i�M�:Z6fyP�F�x-!��?��UP�F!/1�j�o�5B!�߸(�)���_?I��C		b7!�$S�_�Uigӊ���Q�B�Q!��*E8䚐�m�0e�!�� j�b���-��xp�=9/�;~P!�DӐ/>p��W�$]_�4�o=!�D�7��ɦ�'ą�������'��8�る-��@"����~�<Iv�W|�.�xm��>�s�$A�<A��[�z�2� 8��X#�z�<�j a�� `�ʐ�LC"�Aw�<��)�\���#o�&Q�yR��w�<9��Âb	� ��K�lifiRN�<!p�܈$��1P �$g��YW��u�<� ���T�C�4i�O8W}�)+"OxӶ)T/�RtX�#P�5y��"O�L�4���>�
!�!gf��r"O��wJE�`��3w�e_Ѝ �"O�l�ï�=2#�xz��N�.|�ӷ"OT�f!�)nhbG&	l`6�R�"Op��_��a&\7VG)�"OvЁ�@(I�0(S��sd�$ "O����ɖE�x�-əb�|��"O� {���k���i�M�F�⬩G"O� p��1t��u�0o	�&8J�"O��4��uqR	c �H$�h�("OD]P� �1����tAO
M	�"Oұ���ܝ~���:B@,Y�,y�"Oh��R�!����Jя,�Z���"O�%�e%g����)	D=x�!�"O�aa���	.��2㧉�;�,�T"O�rn\�"Xԃ"��Yj��f"O�y����9�}hs�'TМzb"ON�9�̚�v,�ŉ�V5^�s�"Oj�C�us`�3JZe3Z��"O��Seg^X�
	 4��t/�� '"O}��a��F,^�Ѵ]��2��1"Ob��*��q���'-R�1J&XC�"O��ơ�4�@)a�۴[E��0�"O�Q�+	�HLp�_�r�1 �"O�����<g�ȨA�(W�c��4 �"O*PruC[:I�L�9��/~b��2"OQ1���!�z̒��Hm��S"O,9�$�ωG2F�8�B0G���S"O�c�٬S�a�����z?8ya"Ox��Ɏ	r�X)�0� zx9��"O��`�@��`���Ŷ4��"O�|�͒�L{j�tEгS�D"O��X��ۆ+Q~!xGN&J�̙�"O�Dڐ�F&L�����(�	�C"Oģq�4�T$ñl�7U�Nq�"O�����~�mQeEK�p�4Y��"O��P���q�0�r�%H�F@���V"O@1�d(�*ײX�e�O30`dq�"O�$aq ��QF|ɳb0z� `�"O$���$�&�$b�CH��{�"O��� G�	b²3�!"�<�i�"O*�z�kJ=URBH���ԋ�p�2"O��h�YԌ���-�d�a@'"O�dB3�G!J����#fM"B�"O���� �JC�U"f�� 2�4J"O��hr�G�{���� ǉfu$p1�"O�\��L��U���9UD��#|���"O�ċ1H�C�E��#D5#Z�Ċ"OLp�Q*r,J �Ͼ1YdX�"ONMP$�]=Q�����/.Mh�	e"O&,B$�3�Dd
5�8�H-z�"O��#j[��`��FDg�ܴ��"On�3�aM7�6	�$kN���D��"O�P @,��fc$���jO���"Obm��S-BN��
ە:����"OP;u�*l�n	����p�P"O�MX͝�O����U�����7"O�Հ�C�+��pZ���4�[�"O�%c5N�k�2�fcb�ڷ"O.@A�	W-JQ�qv"��_r꼲#"O��h]Q��-��� �UL ���U�<�m�*V�B�q�]t�.�Q���|�<� �,Q�G�)dw��CÍ����F"O �;�Ô�_���s5-�6)�����"O��×;N�Ε(��� {41��"O�=�	x`�i1nN�c]��4"O��xǦ�Z�z��O�M�{�"O&��ƪِR��X%���EI�Q�"OPt��i���>ժ"��=8�	b�"OXQ�3-C�P���$Q"+:��E"O�Y�w-�4{�]�S��
I����"O��#��l��i�6ɕ:v��X�"O֨��W;A���X u�D�{�"O��с��@��ᨐ�L���a�#"O0��H����0�U�	�U��"O<]+��	��)��ḣH��x�"OV�OԷ�0�v���� �	�"O<�#��,���=hL1��"O(I�$����Hz7"ک|\"��"O\S�b�k%�����,@Y�"O�U0�f���`%�C�Ԑе"O�[@&��$�pEEˮ��$!"O:T0��.�mIt��	���\1�y���;���%��=f�*t��B�yR�
~�~��$�ʘS�z�aW���yb$Q7Bhp�CE: �(͓#1�y"�P(V�)�oR���e���E�y"�"CP܄
��Z�]���J��"�y�dZ0`Ht���	��E4��yr�ݮM]2�v�Wv�~���=�y�T��(XEM���X��D']��y�cA�a��L�"N�I�V�C$K��y��0B����¯F֦�U��y"�ן{��l&��F8�|ren��y�C�W��U�˖�E)|���$��y�E�v��\15��)6U�PIǅ�y�&C��L��ӎɳ�,	�S�y�J�:EW��Q��H�N$H�#K��y"m�p,`� ?~}���y��ǽ���U�93S,�y��W.�t`��V�?*�+�	��y�iY�9�nu�&ÙD�dY���y�I�0�Zg��0�P1�+W#�y"�Πt��`� ��$�� �#�1�y$/o�|�0m E�"8S��P�yb˟�&xQ⧃T>0b|�el^��y�Ώc��i�C̛m��9b%D^��yb�
4�6�����O�ms�)�yC_XٜH0"��A3�������y!�;~��B�FIoƸs�$�"�y"-�4H�p\��OG�!c0�T ,D�4�q���v<2h�0�v��)V�)D��(�[?�rI�1�+~��A�E*=D�A�ƏrifA��F�4�DM��" D��Ԇ�+q� =���
P�e��#D��¤�A�w�2hQ���Sv���7D�����P	7-V5�JĻ ]�eh+��a�����V�=�����n��Y�ƥ���4D�'(M_T$�"	Tva�5S�*/D��h�Hų� L�w 2W��}���2D���M�~�n�1�mT�#(��fA=D�\RB�J�]� Mѻ�$q�;D�b��\'��5 U�Ms���1.4D�(v�0κ�ȗ��(1�9* �1��*�ONyBAa�Es��֍O�~hT�@"O����	n)�$-?G4j��3"O� �D���:º�����%!��;'"ON1p�7r�p�2�O�G�*�p�"O�lp� ב-P�r�M�I��p�"O�P�%@�m���c��/v��"O4	�,Q)<��lHT.�6uer�j���!LO�9��P�?���B�l��\S�"O&ŨԎ�(�4�vnKt�T�"O��I��V�$"��r�ώ#�N���"Ovp�監e_D�TiG"�T�"O����N�����t)�#���C�"OVӢ@_
l���$ɉ�m9�0� "O(5�R�D6L�ҹ���Z�	�P���|r�'5"�'�|YG��]v� 4i���n���'�*���U2 o\�;s�IRl��'�ܕ"���{ݲ�����4}��'�\����� p�TL�g����"O4Y�NKc\��B)6yA�b"O~TH�(�7��Q����*$k�"O�����(D��b���)��I���'���>,�i�����$6����OFj�<A���[Vћ�	�$D/��Aŀ�i�<�G`�;O�d:�@I�/�R����Af�<�"�Y�O�.I)�#IԾ��#��_�<A7�e�R�h��͞|}�d��L�Z�<)D���ȵ+��{Ԇe�ĄW�<٢�5 @�i`�E��(b`K1�S��0=am��+ $�R�#��Q�5�L�<�!l�
b����c�0$޴|\hC�I6�
�aWǀ; 2$@I���6B�I�U ����"��U��0U��B�I=���1!�0j�<B���rB�	�
d@H��&O*�޽���V{VB��^�Č�Ա03D@��(��j$.$������Q��Ö�`�*���m��N��x5"O<aR!eƾMlq��ĸU�|iR!"O�$Y�e҂�l��I�6J�tU3"Oƕ�2��;mxL�������c"O�9 �]:&PE���,��p"O��Rq
��G$�P7�!j�La��"O��)1"��4���¯�$PL�8�"OT-v1�P=��M �H!ܰa�"O½�-kL�x �[���k�"O�X�EI։�.���+�3Ē��"OX�PA�T�����Z�HY� �"Oj�  ���1#2"�*b���A�"O�sAŽDL�r��;$#"O>̀�G�W��b&O�n����"O�p1��0���.F�2�`H�`"OHYh�[��"�`d��b�)� "O�:�a��Q���bW��)(��-Yd"O��)���m��=�ТO�e����"O���Ve��l�fBY1<<QB�"O5 3jT�WL�"%��])����"O���өT2K`�ЂEF�y����"O��c\�G�$tx&���V����%"OBh�!Cf��0�R\�Gr��W"O`��`�����OT*�욣"O�5�b�S(0�m�`i�����"Ot��s�� ��̃ƍ��u��`�4"Oh`c1 ٞ ��i˃�Q;k�r<�g"OlY0u�J4�n�uJ�7�����"O�A5NΧnhx��&�7ik���"O��8V)��xT�0c�gL�3�"O����!&!F�p�ʜnb�ّ�"O� f�@�L�V��2��uDX��!"OD,��ŗ =<��St/M�J.8���"OR�vP��<�Yu�0`!�,`�"Oj�$�
�c:p0�A�3�B��"OtP�v�<���j�Ɛ#�z�se*Ot%�c֯,2`8�$^�Opnmc	�'�>۶��>�� �Oe����'�8u��E�}`�r"U�M�z���'�~�(�D�}�d��Ms�E��'m�(��C�Kd�Ah�(Y�����'��G�X'} q�#�z�D%D�踱+
�a�.E���*I> ��'-D�� ��2.�R5�6G�.�Ɖ���&D�����;h�̠k4�Ԧ�i�:D�����K6|�O1!��X7O;D� !@aΉ{�P��%��B�ވ%LhC�	D� 	��T;@+|HV���hB�I�0��f�J�H#P���L۠kC�	�i)|��uj������eW�*B4C�N.̙q�#Dti�	D�F��B䉏,9(ᢂ�J��I�f�V$��B�ɑ	"�	���h�-�0�ұ:�B䉉{�n18G�+��8#hO�'F�C�ɔTr��z�Zfچ͋Dk̛yl�C�ɿW�2\4b֘�Pq���H5~���D�!?��mC��@<���$E6rR!��t�	xw��f}c�bR�TO!�$�p��aă�&��@����0!��Z�9��ڦS��oй-�!�ƐV�Ƥ5�L�|���d[�!�d	�A8E�#H�v�(�k��y�!�Xe�XdK`o�6uՂ��f�/D(!�=(���i*�D�t톛c�!�ĝ9U��)E���)���&lY�!�d������^�o�E� �+I�!�ʩ7����m�1��xr5��Q�!��A�fQ��B��D�`��cW�M!�d�����a�&Xb<Y�3n��
�!�T	�Y��B�n��r,1V!򄞤E$V�3EK��y�t����!�$�)��$4*}�t��MR&|!�DǽC�!B���2Y�&�</�!�N�4�����n'� (洤�����C�~8���L+\M&�n�y�D�*H�T�v��=ܬ���E�y�ƌ*_��YS���h�Pq�3B���yB�L;���8U�Z����A'V�yI�'Fפ���6����E3�yҀ�� ���ԋ1x� .��y��$,.�BJ�� s���y�B
�WN��dA�" ���
�y���-�����xFxSw��y�a�14�ܜ���H� ��*�
�"�yb/�-1z6%�gއCWʕ`��y��*K���� ^�D�,pb��>�y��������Ƨ'���*�h���yrß��|t	�c���q�O��y��W(W��p�V��^�����2�yI1:P<���i^>u:1ȸ�y�G�{/��H�@�94DQ� �y2��"	k��j���$d��'�y�`J�!�dx�S)�1|�(��+���y��r�:�1�蔱"�����b���PyR��g�D��
�a�M���b�<� ��(��ʍDnl��� �;�Ib"O���B�9JҞu��	�C��{5"O��3!&M"V���E"b���"O�h( �'
��I�eڂ��a��"O|�S'�=V#lDJ�֫(� ��"O�����m����� B�@��|��"O�󧎛��)3�d�(��&"O"]P2�n�`	�d��{"��#"Ob	 =0VX���Ct��5"O��@eӝ\�P]R�"V�>�d�"O����F Z�2�ˇ6��U�"O�)@G�<;`�UB�I|���Z�"O"�zc$�	}^<!PhR�X�2"O6Eb!�E�+�ي�ƀ�1��c"Oب�t,�?��3E˞�~I��"OiÃB�=#�s��Y-7��%�"O��k��BP�r����L� �v]����W�'��7OT�TB6���jX�R�"O��� $˨	�@�� �	uB �"O:�����O�����
�I�\�C"O�ے�٬^V��z��ˇDO�0��"O�<0�MTXc��0�d��Lغd"O�E����1Hp~�d�9}�"O�XR�'�-meƁ���.c�Lt���'��IH��HP���p�p��Y�!��2D����ؔwu���D�G�t��T�.D�@Y�f�?S�1g�;u��y!7�-D���C�"i`������Fє�P d+D�������lwT��A�j�&9�j)D�({!�-���V�R�e�5i@&D��1gU:o�F���	�HTɁ�O�$�O�?Q���y2��t0��,Ol�aj��+�y�,xB��iZ��*�z5a͏�y2@O?.�@3��Aj�B��d�G��y�K)�F�C�Bڵ���0���y�Ei2�tkH�.DZ���y"H��"R��Q%*�4	U�\0���2�yj�V��:�B=q��^�ybiprF�s�Ƿy��F'��y2l
�I>�b�s������4�yr(8"�3# ����qA���!��'Q	4�O%]�K�>P�5b�'U����&\
hi��A�C�9#�'���(Q�E$����;����'�n ����M�`1i�i@07I2|��'����cbĮ|�>)z�EV.,k ���'����0郱G�� �@�;rRbE��'��5�&Si��`���]aB��' F5A �v�b6b��2�'�	!��b�T�م!��	nvx�'
N��0c]5g�r�%k��Tĩ2�'$��;5E�={Evx�K�P�rm��'�h��S�!�(�RC]JN��
�'R"8�Jf�|T����WW�m[�'�\$(�eP�$�Ur��	�	�'}�%��<̎ ����N��	�'�r�� i���#M�8m6�b	�'��,���G�lƠ|��30�	 �'� ���,O��j&M�Zfн��'�F�RrEe��BƘ�Y*R�z�'�y�`�?�\YPw偭*��`�'��qH�aU6�� HWI��	^�)�':鹇&�NO�=�&D����q�'쎱�6�E(f�ysvn��d�3��� ��	QH��}.p	w��3�*��"O�p`%L)<	6�3d�~�8��1"O��@�I!������aI3"O��;�� 5���[�}��)�"O�`A�Hۦ0�2h3�J�4N~�X�Q"O����ɚ*]Q�@�kInQ��"O�H#��,jf�JW���Bg@� �"O�	�k[�Uu���B+8I�,�'"O����R5В�imV�+C���"O�[�$ڮ���7+M
 �
'"OPre/�O��I�hܔ01�"O�Y��݃O.�U���35̎ `"O:@�vb�>{&	I�(G�m�P8��"O^1�R��<�45J���
]�}�a"O�踅�9�>�q�O�+�N5�"O�,�5��;[�XP��Oɇj�$�B3"O��&�^�5�C��#	�9��"O����ܠ�ƊZs[6��2"O��b���?oXҴ�I�.@fVAc�"O��,�3f�q�sKZ�Wtٷ"O&�X��ܧd/��L�q���S�y�=�����G�H��SŃ��y"�A���!�hږ9����k��y��@��f�X�Q:yp���$�0�y��.~(�*��B�����ǚ�y2�M�,������,*>9��E��ye��e�ܝ+���n��<C�K��y�F��/�e��AW�4�� ����y�E�Hv�!SA�=p{��jh��yR!"[dnɒsdڠq���I�	��yr�׿\����V �<eJ!٠�^��yrg�Ҡ$ȐL@�T��ٱ�y�A
�+\p�\�L�Fx�-қ�y�C��캔ou��m���ybZ�xz�]�B�C*j�$=����yG��#Yp!cP��_B�m+�E'�yBhL��iC%��T�pu�ϛ��y2��k~�I���S����E��y��>�歃�IJߪ��F�K�yr&^����.OEq<�A�����yRJ?J](%۬6���/�yB�ÂE��5� �S�A#d{���(�yBkً)9eH���Do���y"�ӵ(�����k� �]��gY�y��,w*8�vEF�r}�A�SFQ��yBKD+(@���뚐g.2�i�@��y2ހIм�R�h� /�����y�#X�����ɊP����E%��yBd�.0K~�0D��K�ё���+�yr��:cEF|ۡ�Ѝ?�������yb���v�I�g<���D�T�yR-Z
QZȓ����I��o��y2G��k�~�ʒ�\�t�r��Ό��y���_n �KB[�o�R`�N� �y2�/`R(���,��c��p9"oE��y��R>WqBA���%�y8�m�#�y�I��{N=X�+#���Z3oC1�yhԣNf���C�֡B�,��L��y��V�@�~�bM�>�6��p��&�y*�,�6���$��/F����(�yr���ST�Uc"���b�	�y�<�|hʳ��6O1��zD��/�yb���( �t@��ѨD��Z�l 8�y�
[H @� �K7�����X
�y
� �A�r:Ԗ9�w�=#e���"O8(p��K:y�=�B�ޱ#����"O\�[�)�)!�R��=���Jp"O���dϤa��$S4�T�[~���R"OF͠7F;?Ά� ��"{ցhp"O�����3#�HP��o͠mn}��"O�e�6M��TS�.�/j4��6"O U�Ɲ
u���@,,�!��۴1�X���nȓJ�����6�!�Q?6�!(����1�hXǂ]�ji!����q�)� (բ	: ��G�!�$Rq��+�F�9	�:� �
*�!��ʍA娕hS�2:�9�T��%�!��ۇm��0m���[0�CK�!�1	.0(�4�ާ��`p���2
!�I0A��0"U,{z��-�W!�
@bqSF϶ 蚨�W�h:!���sP�,)T�A&c�"k�l�_!�ٛcR��퍛W�-JU޿0�!�dEl߮�{T!��� �C�@�u�!�$�L#XE�`˙_���S��zY!�/eU�1(K:�.4�MC�f!�d$U��U��!G�,*A瑘O!�܌���!�V�� ��>Q;!�B�w�L��P��<��coט\�!�dV5�:Ě6��� pКCoZ�Q�!���M��p$U%i�}�!��=�!�$z�N������x`�l�:�!�dH(G?����V-`��a�0N��J�!�d��E�6U��¸}��P���b�!�d��\�*$�ѣ��i��K��ƿa�!�ET��wɐ�V��VI)|!�$Z�{��|kȘ�
Ű$J���>�!��;�<��P5dJ� H�V3�!�d�&y�HZQe�7%]��IBU�!�DB&��A��d�2YW���ǺD!�d^�)H�5Hl��6E�p�v��q�!�$�$,K�Z�"h a�e�k�!�dVto�ȩ*T-i��(ae 6Z�!��S� .�ь
�4؉s�#�+C/!�d�p��!L��-�\��#C�MG!�؆r�
XᴎH�S��	ж㋔u=!򤇸�u�@� �`��@��ɶS8!�$@&�Z�]"�U�"�Y�b~!�ą�{޽"T� �"���ZPc١fa!�dX'P�
`��oA#0{�}�4�ɯ[!�$��J1�Õ7)Kb�SpG���!�dO%5��B�L�N��W�"nB!�$�!� ��EJ=*��0�+��H+!��B�g�����x��4a�	�!!��](b��y���ns.�����=|�!���0w }�D�� W�<��*Mt�!�Ĝ\x�����_�D0T�]x!��ٴj�� Cң��@��9��%si!���ԁ�#B�P���[!�D^�-� ��ޮJ)ֱ�h˴@�!򤙮<T�E�s�ӡ.
�09V���}�!򤃬m�
�Jh�����!e�!�$֋z�>H��l�G܀-�U�A�E�!��\;��	A���}��uc��n�!��10�����B�'!�n��c�76�!�d� r��#�#��Bj�*ľcC"Oz��N�鑰l)	v��"O([$�I3�����P�v!$"O� ��� ��vؑ����!���3Q"OР�� ڗvz��C�O�7hD�l*$"OD�x�G��Up.�Bv��"O�p�Q�Q_�
�G�7&^M"O�X���Z�v���!�I�"0�"O,@���bM�����W��+`"O����c�sru	B`�}�L+�"O�Pk�۟B�:�`Լh@�i"O�`����)#��t�46G�2 s�"O��W�	2�RU����k�����"O���#Fé�y����A P�Q"O����f ���l�/�D9E"O"��ǕI�~�k3��-����"O*�Pä�+UpP�ؕ��F�Y+!"O�p�4����TE
\�D� "Oz���
G�*(ΑÔ��;E�Z�@�"O:��E�?��P'��PƲ�A"O�� ec+��D��g��
ߊ�A�"OJP�$FP�;i(�yP�;��=�`"O���M���ك��2A���"O�A���>Tqĥ��]("O�,:S�Lf�J�i�N�N���"E"O��s CR�6$���I@�=�(S�"OtQ�c��9�|0J���)]�R��"ODy���Fʮ�g��5Eq�!3"O(�@Ȅ-�
}�q鋇+X8PG"Op�� �2�p��SR���"O@,��v��3I	;D��"O�9��ָ%�.��g�X(��A&"OD���W�.p���7-��[D�+g"O4�(�C�bE��M@�-!d�Z1"O(M!�'NF��ċ5��*+��Y`"O.8P,�Q�dY�i\2J��c2"O���g�h<��F�U�RB,�'��O0�#5��8t���ŤC�w�h�"O�i:�	������3^���"O����^�2~Dy�Ң�	fQD�b�"O������A���CaL�CK-�V"O�����̻Z�]83��8Pͮys�"O��[GOW�h&y�������"O^�J7)ʃ'Ɲzf�TC�\ZT�'nQ�\Z� V�	i(D:%��7?�F���&#D�+#iR7�0px@+��X4��E5�	E����	,P~�i�)[�\ b�8�O�˓��)q�N	b�RYZqI�U~�И�"OTp�CO�M���0e�S������'���h�#�+l�h�	�D��L59`w�5D����-z�Jև�J���)M���O��0a�����ǈ�J�����L�<�&`�3T��<��
$�PYhBC���0=��OO>HT��RfI�֜�a�dSy�<a�̜)nN�	����(�))�$_�<I�)�
8`G�8,30飃�^؞��=y��=�� �r��,��u��D8����]4�2,�1�\�y�PU�/:D�<�eN�uR,�%�ۤ*tJ�P�6D��s �_�S'�|�����l'+�>a���S�'�||�A��"\!7�i�B���>1�e�j=hH�W�˃��`$�g�<!4��W�y��K�/BNp�LY����kӺ�}��bU ����U,fr�`-X}2�'o�m����./�r!zТT6R�&�:�4�hO1� ��'�N��`�E�x<��P�M����'u��S��٦"܊TQ���(l���{��O���� ����\_�:�k��mnƔ ��'��1|Bp��0��3S�(pAO �Q�*�<�˓Q�z8�v��;%�"<�F��8)���ȓ ]���A�2B�vyG�G2Rtą�`� ��	z% e{�Yw,���I_��10Ѱ���q��	B�bJ,�O.�C�eU�	�kW�w"<�u�y�("<�M>��^�R���3".E%c�f�!G�ZW�<�!�0!s���ȩL��I���Q�<�'�p �CEA�32�`�҅SH<نc��/c�!�G�؍YZ1��)޻ G���(O?u��-X A�-��`�g�&����&�Ih���n�=+o��n������<�+���< *ó�.�z�OX� �v��.AX�T��q?aW��%��{���-\���*�@�<�D��(`�?\��m���MG�H�`D�J����L��߲7a��h�l ���ȓK�f���h�D�1��F\�C�5��q��q3Yǜ�(Ub�0�@�ȓ|�V����k�����(v������>��M^��f��/ 4�,�[�\��f�]4&uK3ț�
��lkd�H�4>�4��E�'�n��g��*O`��I�Q�����}�lv�'���rpG��$�U("AަR��E}R+GD�O/@�!���i,�1��+�0@�h�O��d��a��d' U�;�v�DUL��+�(O�(�OD�Q(<���g�R���`�"Q����<�@=�B��oČP�� {�*��Oz���U�k6�,���@An���V�1!��H�F}��B2"�L9Bh	4�6*�^�R���s��s�1��\k2"S�p�q�">D�d���F��D�6쒽���[E�!D��;%o���HA�O�Ut�\��`�]������(!�epM�+.��"b�Y�!��� � #\,fnM�����F��D?,O�˓z�6��	l,���ώ0h`ع��� P�!�$��u�,���o	'z��]��J��a�I�<��#� ��$&?�gy�(�T&�\����I��}^"jd��.Ml�z��A�KXРrQ.XO$���bQ���<E��/�cJ�,y4,Ba���hO�>3�fV>@| J�#A�#���bCk����'ba{��˴o	 �!��}h�< ��ߜ�ON�<ِߦ�@�̏g�liS��ޓqS�t�F(D���	�2~��x�aa@.Z��4��&g���<a�O?�I'��)/�1'^�,�����@8D�� f�6 ��������5 �Oᑞ"~�I3�~�%)<~��9���>R����$-�H0L ��\�rȨ]c2��.]��Նȓy~H������#�ȡ|L�<� �
Тu=r%$5!gN�RH\(��i�
�C��X� e����*�@�M��jQ��b�!��stD�Nu�Q���?��C� @\;"�A�v`�8�N�<Y�g[A� �+�� !����@��I��G{�`����H'�[�gL�3�l��y�#A)G�ř�H4W�][��B8�yB�O :a0D,l�0їŬr{Z���'�Lc!�ʵ3������%`fqh�'����a�#K0�rp&Ik��#�]��ʓ���qTmʉjPa!�Q�B��Їȓc񮘨co��BFv`1bD/��e��R����������0�C]
z����y� Y�V���
`H���]����s��j5�Y>C��-��кwaD��bf*D��  ��3C�l��}�Ռݦ,q��{��i=ў"~n
��RɄ�|'�Uy l_7M�B䉶~}�l`��Dv�u#���i"B��&R~�q۷��m��YRে�mZ�ʓ�䓆h��D@���T�
�����) l!���<�KF�����)@3��64/!��n����&ԆL�dh&�Z6\H!��,YE8.Ѽ�& x��8nWQ�F{*��X�*@Zi��V�L��@��"O�����L!�#���X�"O�H+`"�4t̸��!���tdY��d#�S�r̡�4b
�D�2�O��3�|C�ɗ嚽x'K:=��@n� 5��6�4�I�<��'�]�EC�$�X}(���J��H�'0꤈�)�i��(� �>t�e����d!��S�&�������9~�ڼ��+�<<K.��+&0�7�P"m��iV+^�|J|�ȓ!LU��.�6=	�H���f�\�ȓ2��!/^�B�.��v�C1 =����wvч*��z����Į�)<"���'��"=E�DCK�&�� 5�A9�B��� ���y��D5ڥ+�̳WZ��4��	�ēM�a|�`��s�A�G���rR�Z$ C�I�~k����H��/�b�+��k��B�I�Uq�����9}�1����4���d6�$K�Pq�AN#^ô�	�n����=O����B@����жʔX�܈K���[���IHV�j���С?<lY��FZ *����Fxb9�L��u�P���!!-�/zOB71D��A�hD�v5�Sl�=b4����z�<m馕�'Ӫ�E�Df�VZD��A�/��m�$%��yB	\�,���褻�aJUꑣBX	�' :�Fy��D���[�cJ�Q"�zu��!:��28O�22N::F�qf�$ t���"O꘩���:����NK>t����"O���RA������}[༈��"O�d"��X.;%�i�5��@�h�0�"O�4�ୋK� �ɷ Ŀ5Ƭ�2a"O6���Ⱥ o朁v�S	�Y t"O�łS�Y*�\�ɤlM!l�t�Y"Ot�"�K��ܥ�&&���t�!"O�]�3�"de2)і���&Q�e@�"O�(A��F,�Jpz��[,<��H�"O0�;�D�)b�0��5w��"O�$�3���_����I�(\�á"Ov�㗩WI|��0�!vG�A
�"O0`
�+�U�����Ϻ�q�"O�)��Ff�0�J�I;�`Yz�"O��3^�a�j���Ą<��\kC"OLT+�Fq<���:*�b�
@"OR����$�z��f�/Wq�<�r"O���iԉ�FQ��٧6i2h��"OR`ѕGU �$A�/�5]h1�"ON��FP-SLf0X�$�w�2��r"ON�� �J��ҤB|:�l �"O�!�`��F��cv�.y$�8 a"O��;�d�&���
 /1��`�"O�lh5�ΈMƾH�0h��U�z<��"O��sr���kR�A�a&Rvda�"O��7J��H��x	�%�"�m��"O�%�d&��A�%D�:m�~�q�"OVT�HB,v���d��:ksT�P�"O��SA�1'����A��}:��!"O�X���
��j4�$�Trd:C"O� x}���^�:���"��_�� "O
x0�;<��5�(�*�:��"O������	H=�S'�$ �4��4"OP���$��sa�@�$��=���5"O�e�A��1�0���T,*b�	�"OX��"AgFH�5��l<#�"Ob#��C�x2ʽ;��˞TO����"O6у�ک\C:숦��)Y\i��"O�b�W.+�\��w�F:T�����'���a@�O"���B�*�y�d�+d- 	�'��Tá��#�����΢�L�� ��D�F�{o�*��m<pЇ�f�8	�FKE"*LJd<<V��X�](�&K(�.x� ���;��نȓLh�R�FK�f���)!�H0p��rHD�F�ʯhy�|����?!F<�ȓE�� �aP�A��-U�9_���ȓI�Q���� ��T������@ڬD����N��� �,8�U�ȓdn���� 1i�h�Y��<n��ȓH�m��KN�F�)f���jt�ȓoR����$؉Vﰽ)"��~�؀��Y��qTHy�8Qi��NQ�V=��"���AJ�!,fxdi�)��dQ>��Y_���B�U{J�8O1j���ȓtaq#`TX�U�筈,Vy|�ȓ��}�3O��E�Ry��Mđ���Y|eR��&}���Q�|{�,��|���`2��>���wډY�i�ȓ���`�Ӹ=�x�A�dĄ�䠅�ml|���O߾5�d�U��;-�:��z?�Y`��W*]~��$��B�,��jS��P���L<9� ���J�|�ȓvH��� Ė~@���Z��aV�����R6p����:��чȓ,ײ��
]�B�m�`6
-�P��r*����B%r 2�wh(�֘��N�H��Ӓ3*�٫B��7#ZŅȓ>���p�/����#�F�y!�=�¸(#Ɣ�p�\���N�0l!��}>dPVo�2^�ȱ�g!��B|<L�)4N�%:������4�����Px��84�u"� �p �s��Z+��O�8��)ZA�c>�[���6j���,q���`��1D�0�O<U��|k�m[B��8#�f�>aD۲nܔ���9}��i �tlZ� ��2�Z0@�سJ&!���.`�4�	FʞO��R�c��Z�' �`�dF.
)���Ov�*`�� n��YRE[!.D�+#�'gN��@�B�HUψ� &�h T��.���{4A�����S$~�~�1��&c���ƥ$�t�,�#CL*4���� !�!U�`�����*��0HE"OfxяթOi��#�S�{Ŷ��Y�tb�@�o�>���>E�e�D�l�a�qM��؅�y"�-b�B��#&�N Є�^�G��M
�P I̿����'��48%nP��>�C����W)�@���hz�Q 
9W�H�W�h�H���U�2.�SE-�O8��V��"]sH��dG�<��Ͳ��	�~�	E�P̧GeBAOB�\��gf�&^؋=D�X��dD�?�"�K����*��0`;?�D�2W
�"|R��¦Y�YX��Jz"c	q�<IrNK|Ρ�"(L|�@ӓ(Ro�<9�ˊ�i�z�2�%�aCh�����A�<�C2U2�Q�6�Z�?6��Jr���<1��<�V���jO�2��+�z�<� h�!#�
 v�xh�g�G5܉KF"Ot(����R`d��T+��3v]��"O�𨴂ٱq�Tt��y�"O���$A�&Q�� fDIl,z�"Ob��cIR%,>�
7eGZ�Pd�"OpySt�-2S֬�P$�2Ґk��I�W�tqCT�Hm�Oh�!RPDA�v�*B�K�V�@Ek�'?b�f��(���3ŢɣU�N�x�cVlCbE�b�~��s��� ��K���q��78_��,D�xY ˉ=\���A��;m@ ���O�����\�#6��&d0LO0D��DGu�!aCC&6`~� %�'�8|"��FU� \����/#g�y G�M�8|� ��mG!���7�8��W�fu����w��O��[An�8Vv1 f5�'@��-��!�>}�mxb�,0��Ʉȓ
  �w�ԉ<��	 ���o�,��@�~�V��#/ 2�j��&OAR�g�ɷ:��m���Bf83F|�Z��&�|7����M3���;���i�Cس|[�ū'`�g�>��.�;�)��]�|^�H�3LO����K�WW�h	�3g�X���;��McEe
�!=�� c6O��_�TP�t9���	7m����:���3r��(�ƱP���!o(5�S"O*qz�b.�P��ִdE�TI�r�z�8 ,�kT���VL�-%�IڄH�T��ƅ�,h̀��҂��z�B�6D[�-�� م"�~iBA<lO(��_!J&�#��ߗO:�s��0p$p�jS��
a�t��d!R�D�#g",4���pv�:L6�c�џqO����
[��ةa�E�_M���1����k�nl[�O�<-|��ç4O�)��|bP[FiN���pAU@�pГ�6�y�3ҠGe,T@u$0lO��p�ݣ}p[��'RF�QSc��@g��-r|!Rń( ����q@�' B�]� hM�g�Z+�2����?P�xB䉻<�R�JqGT+N�]�HL�����s�E�~T��Ф;�Ȑ� ��:=�X�n*S����G�7T-q��i�!����Wr.�rƊC�+|�=�ד
������Kf¼	�G$�<Xo6�2RDV�L����⪄�e���5&�/ Cn����*/�D4aց�?^e8�
�����(��c�	xdh@���qO��M�Z��Yp�ERzh��r��]"vΡ�7��'������>T���x�bTz'��S�+�}x���S�$c�n�#!�?~���a��;H|Z֋�=j��gl�X����c�j�aW?���	Qa��= SN�,=GZے���I6$���"O֡�:A��!�E���A�t�J���Jܢq�м�F�^1I|��`v�����
 ��:4��f��)!G��+��zR�4eZ�AF���6,���%-[4X+��{�=�8!7#�]զu�u��8eBa}R ι`r�0�!%'�%�iˏ��'|PꂣS<��a� ��k8d��`���iS�EȈx��C�)
��A$P!��N���!��O�:�E�Ds8�Ʉ�_�a\��Daݠ0[��pD�CZ�O��� a�9���¯v��q�)G�#zB�z��C��?0�m���f%,\��I�/��+�����xb��G{r��+NU`�@R�/Y�q��G�0>�B��N>Ą)��wLR�i3��"&�^�x�(9_tmq�d�7QZ(��	0�Y`2DY �x��p��&n"=!`Î�.�}Z��Ίo�P �wJncb��!J��y"�P�� �3}�1pA&��yrΎ)�4"�oZmT�!%��y2��Q�@|
F&Ǥ[$񱑌���y�c[�\v$ �Q��R�
@��y���230�lkc`-V7�UQ�E��y�mH(<��2�ƇR;:]��mђ�y�n̋'��W�ؕMH@d�5�Ы�y"+]�d�$�B�O W�+瀌$�C��y�Y�w�ÝH�|��'��K��C�	!�d���
	 ��s�HN�d��c*��� 0�O�1�#��<��UÇ�U-�<Li�'����b�+����	 c$&L���''�a�B*X��C�ɥN�X�BlD�N�p:�B/'�X�a�MW�s� iJ�bWZ�O����1	ށ\���seύd�	�'�-P��k�v aD��$�� X 0E�}��*�<�I%�gy�%J��̒���9��*�\=�y�FT��2!�`@ӆ0�%�g*�h@b��1	
,E0c�1lOЌ���55�X��S�[� 5D4p0�'�����I�i�ivH}	V�O�2�x�/�.?P�H��� t�D�Z�9��i0��N$>��D���dR�Et�Qd�Q��#}���ڇjid���I%��p⁝U�<�!��t8&}�#̊C42H�q���h'cS�>0ļ d�'�9��db�H��A6a��$�A�2��H�")�O�`a��7�B���?�(m{���C�� y���+EԶ�Si�o><��	%=��=��B��K�T��C�O	0#>���P�"uX�D��H�v`३���bFk��Be��pO&#,hH��\�<qv)����zG��'0l��ۗ`��<!��L.r�f�ɼ|��aVi�]�O\Z��7��(; ���c�zR>��
�' f�����~|>��C�èk�Ҁ1�O�`(a�Q�p=!ª� Bv"qk6E&SC }��hF���SD�ÐT'�z� ʲqp�+��Q:$B����B-D����I�8�B0����%(��a�-�X�́È�	ʌkt���C�(4��(�C `t!�dA�
�4� br���"��Wy!��V�/��s`j4V�D���ͧ!��Q��τ_���s��6?Y!��3p�R�xN =�V���e/U@!�dF>"��<r$�+0���j�NZ�;l!�%Z/D�ɴ��s������]6!��up�!�#q�𴃀⍤#?!�D'p�LK6%�9�����a7k!!��J�&����K��Er���r(!�JH%�]���؞R�*I�r��ɱ<�X]8�'A��Qt�E�^�TC G�LXb9+��H�;�걀�OrLڤ��2pD��Y�!@?~��)P�N�	���;�޹�y�MѬk<�Yr�NВzpri��b:�?��ݤ�%��')�[Í-h;�Mb����'Fr��R�+�E�ZD���@"O^�`�K�����7��t r��	5��0� �z�hIakgӌ�'����GO+�D
6.��[��;N���0J� �a}"��-Jta����DFl��W/A[jM[�eN�'o�o-W��M��J�o���Y��'�\�
�	
�윩���j��؋􄅟P�b�a�+D�M��Hf�����T-2�D��b#+Eh�#�b2q0�a�4$�P`�Hˌ��8��/B��Re�}��!Txl��ݴQ��!� +?:�ʲ .�s�1chT? �8ٳ埶Bb^���)D� ��ǿ-踑R D�;x�n�z%m��S�b̻R�+Fr���N���O겍�ė8��?�
��*
��e2��Q�K�����d���C�݀a]�b�݄l��쑴C��Q� ���i.h��0�ђ;�n8�Ej�DX�l
�Ͼa��{���EM����.ғuv<;��_1��7̈́3GK��S�O�e��`����!��3��1R��S��'ݐx"���qV�1 �~�Ǝ��?�  �e ��'��	Cg�+�Yv�/�S�Sr�$BLѻV�,h AȱH*
i�ȓ;"ҁ����:�c�J+fNɸ3b��9�]�У�����S�G t�'��]a�D�c4 �x�B�&�pŠ�'rf4+#,̴`U�EJ��!��H{(O�]1�b�) �����ռq���[6��4��D���3!�!�+���֢Z�0��@ �* ��!��¡4�����0w�!i�o�S�!��
P���1��gf�}��[x�!����tk@�{d�M JQ�!�ge�e�!��*�(}����ik��H�D�J�!��1M���[Ҡ�8tV*D{�̓�Py��l[�TrD'G�P��t�q�=�yr��=�T�"c��[�${��ӫ�yeZ�W�P��!�IWn�x���yb�]>~�X#��[�P 0iǔ�y�W���gD�"Q�����yb+#-լ|���\���#��"�y��UlĖݸӥ/x����E_��y�H�@�$����	A*l<��o�	�yr��?11� R��J)	���<�y��,͈=
�a���ac٩�y��6HƉ��`VwN2��yb��#�����fѭ	�lKњ�y
� xh	�g��E����c\�"O8�Ê�{H�p�
�uЦ��'"O�-��N�"J�QgΙ�`����"O���Oڀ)G&�Z0l�l��"O����o]� ���h��Jqu"O�@ ��4G���R��]�1�~d"ObA����"��@�¡Y:uU����"O>]��%i���1�*�7^�! �"Oљ �C���&�M�!@�R�"Ov)�1L]	��,��e��"e���"O���EK�?jp���[�U�\(��"O`���N�F��aҤ�ڤ�&"O�e* ���tPB��Q��84-�9Cs"O��+c �),:��'�"���r�"O8�	A��=J|�x��C܍/��X�"O8j��<sڝyDkM,�j�C�"Ox=KR�[.T�8�p�K@,0���B�"O:��̀�rPq:�*T�Q�m	�"O��j3-ͥ+zk0HYlR�2f"O(ꂁG:�bm(�H���"Oz(����?~6�1p�X?�0e��"OH��D����x��'B.?�čp"OPH�W
!ub�U��D*$�rQ�"O 	�UJ��RE�� 4CY9 	t"O�E� M�R��ؠ��# ?R�x&"O��zԘ�6q@��M+F܉$"O� ��N��ĺ����ip"OXH�����Z�ˀ�z��PP�"O2��DزEf�����/@�\��P"O��*��I0l��8�E!��C�>�8v"O�0�g�'hN�ty0`�0Tp=��"O>�g\�+�<�8� @�C����v"O����ҝqĲD@�!֔B����"O�YЃ�
*h��b 3#�By��"O*�:Ĭ��G/R��w�����!a"O��N�)Y3j�!�'ѓ02��g"ObPس O�t�DKu��8�� �"OZ�k�d�+?Q���E�	,�P)�"O�=��M9G�:��� 7����"Op8��k������+�?s����"Ob�I`��(;Ъ�4y�x1�"ON)�v�Z���窇�����1"O�������`�O#_��lJ�"O, *F@�Y:� ����v�0a�"O�$�rΤ��[M�?S�kRO�,�Rĕ1_n���!aҨ �c�S1f�DT�'��<���A���Rv'��%���R����n��j9��Vh^�Y��@�X�1��	 �B�I2L$�0���[2�U���2���lv��AN1]>�ӧH��D���ha��
�h=s��'z�!��x]��A�L�/�|��L�߄�'\�!��@d���O�E˵�&�z' 4�D�'��}�V����R2���d�b9��G¥M�� ka!Im��TCEG�oda`�BH �d��)�+?�TC����G���bw/�,W�lQ�f��=���X#"O�Ј1"�`��P���[.D�BV]�[���#4��Z�>E��̃<���

5c(�� f���y��� �n�a�,F}�� XU�җ��#���-.o>e9I|�>A'#*k�.�#F^��C� �x؟@׎ޡ13�\Qo�9a�d��DM5s��U0FC����"%т+d:��b�A:N�f�����<��O��ɠ���:c>��☞?�2�S�%��Ѳ�>D�X���L�8$xT�ϏUg�5�>?A��L����"|B1LC�[9~yX�+�u:�;@�	t�<� �zfM�0�dk3G´G%�u"O���#
.%!�A��T�[�"O�P!��݄h��h���=)���"�"O�I� n��0c@ ���uꚸ�R"OVP�䃇;�>u�D�жb�.]cR"O�D�"D~��ҫ/���S�"O�DBN\��)b�St��e�E"O��`e��<=��t�D��V�T)��"O^�3^%	�� `5��+"�Ft�""O =Qs�W4�(����~�T�( �I�b5AS�t�OW� )�Y��@݋ Ue�E8�'W �q�9
F�
��ĀD�|��eER/���`!Tn��s���GIC�����r����f5D�$��Hײ}b�h�b��J�����Ov%�GM�+AЀ�,/LO��2t�˯C T	�n�=��{��'�NՑ#hκ���TĔf�>���݃I�ԉh�Ɇ'!��G(���a�@"l���2�O���f�� \\Ys��!�'BC(�2ࠐ) �G'�&����ȓK��y�k�ǅ،R�q�LI��I�Ӌ�B��(%@N��<�}&�\��)�v�6\�����1J \��k'�X���\�P�d!��Ro.`�Ď��j2"�ه�I4L�iI5f��H���Do����f���UnJYچ�Y<ec�A�؜��-�<��dl���P�4�"MWl�4(�h��/�*m82$Q�	�<*\�i;&�һ�y"蛭 �E���O"���/]Q��O�4ӓ�	=/�Te�"�H!l�7�n>���$*���ݷ DT&̐�l�Pt��*Զ/����I7"J����(o��FD�+v�2*S��Җ��aE`��g�#U�v�˒E����{RNL�&��S�D�_���U삻��O
h�U���/b��OR�+�R�+�\�C��X�SN�'}9���<n��Pq�տ��=i/K#�B���Nͳ[` ��]?y7��u`�%����!V,���ΐt�z� �O�S�- � * K�+-�P�I�`� �C�I�]s<2R/Ӭ6 �(Ta�p�u'��m�u@'��E�VL��.��S �\<z���3i�n�11j�
/O#q���/Z���~�
��<�ܘ	�F۰l���ĒU3@<���6�v���͋7j�L(Ie��"}k����ܑ�����Z�$qx�I�"$"<F�$�^���+����	2����M����4Sji���Ui�u'�,� ��f�:�P��n�F@�礀�r�d��1�T�Y�6(�& ��c��WB�2��Q��?yr��9q�b�t�2�0��>��I�d䙤FB��sV	�w�<q$��w��@+� (�
|Sp ̮@n��SW�'"����A5 �ܦ��On��UFR�h4 ��FΞZ����'9`�����> h�5ϗ�n�"d�6j��@h�كG��Z�h�¦�'����MKb��0�M'h�z�*���؍hPLp��e*Ys�[?���i�<<���I�S�X5@B�;D��`��W2a����[�*�{�̴<����nO<�(��Q;�"*��F6�,�[,[�<81��Xg�<�0�{ܨ R�E�e] ����h�O>�.G]���$ I$h�T�Wn���+M�!�D
w���9R���F��ף�Tݤ`�H�"�a~B�Ńj���ៈ��-��)�.�yR�Mu��c�DB��|`0�S-�y�
E�\�e �&��?�p��b�S��y¯^��©����2���y�	�y�NC����S�C!5�L�*�+	��yB������ӊy��(UB+�y�*_Մ�[2'�$is.���Ƙ�y�OQ�MG���6 Y7�,�� ��y�E�s#fjG/D3*�Rq#����yr�X�o�p�ూ֦h�����4�y�ǈ��)�ģ��afr<x'�yBb½�X���
@,B�KQ釒�?���E)/���9m��@+���<* ��RD����	�F��H*H�vs�ˬq!: ����45�`�����y�锸[��3!f�21��e3��'�6�)^�u����ّ>:bN�m=�$��Ǟ0U�|A��=D�d�&�Zc��uy�h�%n�`p���Z�lغ�`&^�����(��)� �e�s�hH�(�c��jO�W"OxD��P%>s"����Tbpk��Ǵ-We��E>�d��	\˶���"ĥ?V(ⴎ �QK������ �C��U�nit7-�7j�����z�r}ao�
C=!��ۖH���@��>��Ȃ��	�qOp��	�^Ү��j,�'r����S�M�@tAP�4q��T�ȓ~�0�AI��m��Ce�G7tZ�بwJ�A����V�`�<�0bX�Gn�
&�5@�~��D�M�<a�=j�Ri���ה5?��ё���$͓��UvYI��'[Z�XU ^�S�Ĉb�*w��ۓQN�d�E��@����1F��/UD4�a��B;}�!��(�%�֌43@i�'
5`�OFɰ�AL/R"~2�,�&?�9Ư4�N����KV�<���4L���x���4w� zpD�^�<�a��B���;�E�C��̩5��w�<�2�YkĔ�G��v"0���p�<��%O0e8��H�v���cWn�<���ЦG�h�J7!T�j3L�j�!�i�<y3f�a�ڡ+���N�\S`�]�<��N�}L0�� c�fR
dģYC�<��b�	p�Z���6��%��!�d�<��KK�� �.ъn�@ìb�<�F��d�؇_o YZǜP�<!tm��8)��ý{�i�S��R�<�! �AS~�Ӏ%�5�re(.SV�<YF�	�<ҸD���@�4X�IW�<��$�H����剓���C� PW�<i1)E�n�X��\eJ�k���R~�&�!�ΐ��ɛ|�������̜c��Z�'r">q��]�Ua�&��Z!���~��A�J�qԌ@X�,_$jp� �%D�$X#aV�bht��ի��Rӈ(�2Od����\����"$>0hS���amp��~�%�/~�qg��o��� ⁗0�y���X0#bA	X1Ș2��2(�%�%���5-
��EC�(*�U?5s���[6�'�⍊&�Ь�&�J$���p�:̋�h�VUȷ-V�RժD�g#�1v|h��܏#�d��G�j�h�	F�H|.��D��<1�I "0��ģ���?x�6���t�'N���Vy�Ym�z�"��H7%�8Ң��x{�(3f��ժ��'�0/�!��b��t�F�bY�(C�� 7��vZ�k�ܘ�3��ԦeAw�L�ܒe����7y1�kl��mF";W��sDNe)��w�!�dQc�! V!X�M'�4Zデ?��@��d�=��BI!6;|6Ͳ~2�ؠK+�&�ԈrD�f�%�D �	�bQ��2�Od�
"�X�Y��;Rh��l4��x�J�*��h��Ħ�M�M��H���V�n|��DB!3��(˶�E*�j,q��!A���BtaPdt�qK��i�n8AǦ�#D�0<r���o�b��T��@�v9Bv~�x�ēQFl��1!�_<�<Ӊ�6�Y��X҅c��<�A�ٔRAb��A�E�^=q�t�҄Z/
@@3�'\���P�B(D�p@wOY1�扛4	��*9�D�F��t����ɞ9J�  ��S�ʧq�"	HH>I�D�d�!*�~�0�Y��H�<��k+��C"h� OF
�[S	ONyRO	�4 89��'�J��'ː)�tQwt�I�
�'��)��B͏<50i���Dh�q
�'k�YڧO̹,;�GWe���'G`Kpǎ#r&6\y�A�,�ڙr	�'6<�0��f�D|�@�^t��0X�'�Ur��S���8�fhN�\0�'�Ќcfh�,Ti�)���@k���k�':�)�(�<N��`J��k,n���'D~ �$��O�B%'Z٣�'=�d�'�g��0�F��Z�����'9(	Bʎ	�R�aB�)�t����`�C'3�T�z�bQ�K�r���*aFҥ���*k��pv+�"?�h ��FB�!���%��I�� F�A���ȓK��0�P�ԁ7�����LA�>�}��S�? �����F�:�lκhY|�z�"O���C*b���ѡ��Die"O*{�Z�r P�#!`�}$蘂d"Ofe'BMg�|��P� J�0�2"O&(���\�1E��� � A�x ��"O�XRC��6kՔ�k'�	@���y�"O,���[�py)p����g"O�����ڰVN�x(��A3`��QS"O�Iid,�+HذAY�NZ���"OnA�ӈI.� `4^v��q��"O�5s�(�}�9�@�
6�p�`"O��ز�:K��t�R�
jP�i0"O= ��	vO0ɓ4�ӹpR&�q�"O$�x#,�AsfD���H.A��� "OlѲB1��-�M?] ��y6"O츊��8OHH�r5��Z���0"O0��O��i��a����!����F�'XfH�f�.y����jѩJ�-p���X��E���0��&c	1/�	���S�O
��DLIV�zadš?
�uR��HKƀ��O�Y(O?y���%*[�qW�E/^�I�Cӷ:�r\����O�Ƶ����9��d"�$7�tU�$J[ܓu�(X���z��r��$�>)���0/c�!�̉�.qO�Y����	փr�2��YJ�-*2�,? Eʣ�������Qh>>V��As�P�. QDˈ����s�:}������	�.�&�cA�>9��BB�\����b7����i#�� cg�������TJ劕_E�"=!r�O�0mz� �	:X ��_�>�j͉�}B�/�IXa���h�fK6|������#\�FU��K�ΘN'qO�>Ɋp��(PTlȃW�:���
�$d��
U�&�S�O�-j��MME&++�b�[  �"�Oa���I-��;`���MP�iE���O��1�O8�j�ՌK��� �*��U)����>�h�a�P�#�OL���/F�<e����@ĘQ(��Q�'�`��CFJ(:F��"K�0|z��s�p$s���h�����U5Mr%1�(�g�5�˽����Z`�D(i�aMW�t�P
�;Y���6l��?��')�͢ç<�\t'ޗ^@F�hsnAnc���3�5}�Ɯ4��|k]��ŞB/�
Q��%(��x����r<4��'Q����/�+�zO>9�"��20N��u���+�TA���y�/K<�Y%��}
���*F҅0��U!I3��iM�PK�Ġr�{\�O�O���I���T��+���R��["	��]("��1�,ع�(�5X�!� j�Ŧ�;��ON�u{�Ϗ�4������W����7w�����Mk�ʗc��O��O�ND8�:f?�X�ϔ�F���z�"OV��gb<;I|�j'�RTǺ�� "O�mó��-"<�� 2�Ǫ"�F"4"O���R���C��u+uL���l�"O~(0��޲aQ�9�`�[<"�:Q�"O�Mbh'� �e��`f<� 4"O^�	Cb�P^J-�ԣ��	Nl���"O^�A��0���Y�Ю@C�9$"O�� s$�X.�I��*��`��I�G"O
1:$��5y�d��@�F�V����'}���3��霈"0�ӆm�t"O~逢�Z�q��0のQ@�Ƹ�T"O�+�L�ɊT"3h+��0+�"Ob�Q�ؗJ�!P�ۤ�J�/�y��W*��ɤE������+��y",؅X��p#��6��}����0�y�
H){2���!Ƶ1�2=��R��y�&'n��d1EK$��b�_)�y�힙WO��×d�I��z�OѦ�y���6��<��`��i�t��@��'�y�H��[yޤ��+�!i~Q���E1�y���[��	Qԡ��cT����3�y��X;0����T�Tǒ���)_�y
� 0aUO�+b��\�'C�Kqd�JA"O��PP-�&g�� �$��'\@b"O�䉣�_=��厒�-Iԭ@%"OT�f�ވ�F�B�,��:�T��w"O\�S/N>�,���K  ?ْ�%"O� P�V2 L5��ߩ[�.��3"O��	m��&�� ���1��8`0"O��&k��<1��:�°o�m�#"O�)X!��;|��&��K+l���"Od|�`	�4lbNxpG;g��As"O��#M�G�{����1�D8��"O��:c��K��1�Cܸe悕�"O��'�ޠ�F}0�B	�~E9d"O��c��Ey��KaK��.��"OX�C'20�t�po;y���rw"O�	�$Ê48|���@ȬyG�{�"O��۔aΞs�M0�`�XAza�"O\p)]�S�D"�&(��HOk!�d��-&�P�7��5��m�+�!�@�6�������ި�8@�7d�!�$2E��TrP�lʂB�"�x!�S�U{�M��~K�� �3o!�J-�v �f��8���dD۰2[!�*������c1(uSF�uF!��L5�8��**�7%�"9!�D�&4�f��ݑ'��c�L8)�!������B�R�kf��{gOC>nt!�$C� (�)V�Ә5����MN�n !��-O]&5#Ud*��m� )�!�$�`�����Jq� ���~c!�(Z
�Y� �6v9 ��坠8�!�d	N�[f�Ah��Ӥ���!��Ŭ�&pa#K�(z?�Ԃ����g�!�$T�z�����q�9�1�K�i!�I�Hx�%I�#^�|d3��`g!�+_V����(C�`0{djE�GY!�d��й�g%G�$���+���9jX!����8$#��*h�؍GDR-SR!���-"]�t��f����}��ȅ)Bn!�D��|֢ s�a�El@lZ���1!��N7 �����
�m_�Q��!R�_!�M?N4	�3Z�ūu��#Z!�$�z���fU�-|ha�+	N!򄗺'a��0�4R�(ͳw��>
�!��&H�\�c�'��(&R|�!��&fw)fB�3���Q���]�!�D�]< 	�#d��n������@�!��A�p��0��*ot����άD!�X;J�~t�%�@��i#E��g�!�$ɦq.`�b�,^�Tb �#�d[�j�!�<04<H8�_E��)�b��!��9Y� L �k=?8M�C�!2�!��ݰ(<Ep�<gn��]a�!��0iO��C�[�\0jY�:t!�ć� ���C�$3"ش���%ZX!��0n;�Q���.v��� �"@V6!�!ҕ��BW;ހ��r�W4H"!�Ѓ7�ǃ";6�X�jؔ�Pyr�� };huI�A��Lh�C'��y�/̿q��|���[
h�#pʐ��yrOÊ.��ԉDh�?6�ãR��yr!ݜ~�^,"���G�|TP'L��yn ��MiA��5l���A���;�ya��9e� )�
�kv^��c��y
� ��(s*�:�`rl�3m�  �"O:A��B��"�e�Ͻ?���S%"O�<�nF4��U!�Kڇ#�����"O�L��+�>���IwK�|�4��"O�@R,ڮp���c�+��W4��b"Ob��&~����?|CL� "O��JRa��p�PK$�˷.+�Au"O�H�w(��� ��-�yiE"O��ҖM��'P��S)ŀ/:�Ö"O�5p�$�0Jr1Y�J؄;�� �"O"�2���f$|���=8��-;"Ov��BkV+�B�8��ڬ<˞�Pt"OZPٱ��W'�V��46�� �"O�i��m���[r�CT $ s"O���QfΡ�V�ǃG�4��6"O�5��.D. ��&e��b""O*�u�H�(\�PY�%\9E>Tc�"O ���`E�]V�1c$K5AD��"O�⁭ec��C*��Ek#"O�=�T*c�MsRJ]�:%�E"O���ϬwA�|�� 	 9"O�a*U�# �|�p��&3 %8�"Oġh���^�$a�aX"$ ��1�"O��8�o,%u��S��7g�:�C"O��z�ͽS�4�#&.��E����"Ov�#@+G(]x`�'P�X�ݸ@"O����ʛ�m ~y��FP
_%���"O�h	�Of٦LJ�HR`"O�q�c�_{��@�s�==p̬h"O؍[Ƭ�d����	�#Zm��"OZ��2aX�R8\�T�TĐyt"O �`�'˜�����n��xDP0�""O����A�\ �� {����"O�Q� ��mx�<0�(�5��|cQ"O؉�G��v�x��I/1H���"OX�{0dV�h"���<a�z��U"O"���2���'���n�¨+E"O1�X�@�R��bEܬN��}(�"O���T�ա>"\�����Kڤ� �"O�e�����F8�(A
�?�8�i�"O��Xʂ�gy�p�-`|^��"O��@匩�!��& ]�8��"OD����\�d���b�X�h���"O(�(���"l��!i�j���1w"OT����R�&(���!�K*���@w"O� �A�<y:@ �^�.��j�"O
5i�d�	Wjy��)9Ty[q"O-@4���A�ʨ�d�Ny�]�"O�A�;T�6��%�W24�F��"Of���Ʌ�.�A✱[Z@�Q�"OZ�ؕ��7Hx*$��bYh=r���"O����C2ٲb���I�V��"O�<K@��e۞��dk�x�p9��"O�Ly������|!����0�S"O�TY�JQ(R)%@L��Y�J)�"O�!3�g�)}�m:��H�k��u��"O��HEl�&�X@�������'"ORY�Q�ٮ^H⭁��A9c�q�"O�X"LX�z���e6X��;$"Ox  ���1x�:�KE��(�b�"O$�����n�`��ӄß^�\��3"O:cgl�� ��p�5�����"O�P@�߀Q�2�H��[�h��c"O���5F3B0�b�F�F�+R"O� �D ��֫rQ��a�&v>>�Y�"OPȆ,� ܋ҡA.U\���"Op$;�gE�c��ؖ��)����"Ox�����z< �#qpA��"ON��0'[�q��D1r�D�
�
f"O�0JA�AB-H"�%5�YC�"OLH3@�i1�� �B�{��H:�"O�	�`k7	����Y��d��"O�0Ȃ� 78l��N�i
�:�'�j��n�T��oQ�}��TC�'�Z��5�=<��Q�FT�q�:Ū�'���uE\�y�,𐫏 _U����'Ĉ�قBZ3�XX`g��h����'{�aR���>N����[�X�̝��'������@3K��sPkӡO3.e��'L^��'i�:q�z��D�0}f����'��h�TI�$t4����!��]t�5H�'�F� �)�E>e%G^�Z��i(�'zȸ�j��i:v�@��[1Q�� 	�'}n���_��v����ƭ@*�Z�'�¹ӵ��3\���GS�:�S�'����B��4���IrFE�f*I
�'������/)�}@���_5L`2
�'�5�����C��]H�aS	�'��,�g��H��8�$
�U�dJ	�'������,���៵L�(@�	�'��1�è��=2 �1�A����'&J�G�?'����0;����'u���Di�n�scf_�+^V���'��p�w�Áx0p��RLx���';�Q�g$��,�VfXN���'���zf��o+T�fD�=��5��'��I� �'?p����P>g�0Q�'�6���MS�+CV͑Ai�O�Z��	�'gt��B�!�JA�p�ܭ6!^� 
�'u@�+��ڿl�4H��*��|Lj���'���������a �l�Z�'#�S)P:���1W�� L�e��'	aӌ
$8N�d��e��+�'z ��6I�Mnv�#k�6E�	�'�Q�U-��E�t,��`W r�~��
�'L�B�a�	B��)RB��A�A���Z�9@��� u��D&lD�@�ȓ*r�@bD I��B�).�%�d�ȓZ��(���¬jQ��@������܆ȓY���)��_�B-رa ��M�ȓD�� @�?�   V  "  �  Z   ,  �7  �B  �M  �V  �b  �m  �s  /z  ��  �  &�  i�  ��  �  2�  v�  ��  ��  =�  ��  ��  �  ��  ��  �  ��  ��  ��  � � e U �# �) A,  Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�� |d��"O
`�(�;���8���-0��1%"Oj4��ND^[��"3/9�0|H�"OB���H��*�ʞRy=a"O�味V�!X��!&F�:J�$���"O,��a
���C�Ą�M�"O,$3%o�-���p���+Ն�:1"O��ݢ1����`���y14]2��i�<�6��{_���c�H�`�fX�$Kn�<��A̼VI�xR[�)�Ć�pඤ�ȓA5��('nߡ4�� �)˩%� ���,��r�؊b#`T�eT09���ȓ!�b��g��}�8�F��-? �ȓ
K|m�ș�VṔ���2�%�ȓ"R�X�j�4JN�1�˘X�i����̹	_�jZ��1!g��zܶ��ȓgil,*�J�
j�Ne��i�J%b���f	�(U��:���G��$Y^م�~r�� S�%T"���k\�jx�ȓ|4�1�îJb��@ӵ�ݩn�V��/[`�"�v4�R�!ʎ<��M�ȓ`:��z�ؚh�J�Z��$HY:	��H��p�m�C1��!��B:��0��EnjZA V;9����J[
2���	��4'J�EA�IVW&��~�(aZ��ӹ�>� o�Y�|�ȓ�f�A�
Ο7�H��M�$�����mޠP����/���ANXo*�ȓTv�����{ ��-7�*h��I��sB�8�8���3������X?����0W����(=��
�KN�<��,�c4��0�N?,�R� P^ܓ��%�'Xg�a��^<Z&�kEOƢٮ%�ȓ\TF�n#��a:��D
B�
f60�(O���M�O`��yB&L�6Z�3v��/����A��y2�0q`���A�Mh0��A��Ik��hOF�x��-mվ��NȌ2*PGO��a��VU� 9�ノ*��qc��O ��r}��'���	2�LvM���PvXF��UA�ZS<4���v?Q"�|RMT&V`��hBJZ�1 �ò�̏ט'%��)
��G�(�l� 7�/�D!2ch��b*�<��2%���ؘM��;@C�2,J���k�'�џ��Ыߣ"�Vd�D�7_ʬ]���!�eH������y�π�r.
����f�䡐�.��nb!�ƥ�ⴹ���>wTuJc(Ņ�"O�৉\��(hb����|`B���"ONX�!(Χ4ό��V��h��8�"ORp&� �vQI,H'4�[�"O���O҇bJ4�v� P��"O(2�
�04V��u�Өk��h��"Ot٠�f]2Ԭ���IȾ_\�I"F"OVȺ$� <����h�=�� �c��<�S�i���!B�FǛ\.��7�U��!��v̜ѡN�5+��G�ǜ�!�� t�t��@K�z�t�w,�ud�{��$��U�P�C�ϼj��=(��S�PV!�M�w@�`��� �he���Q��'��;��\-~�mZ�����	DnӢs@C䉃��r���VÔ���л,P2c�@�'<��/x�"���,��e"�.\�M������#D��![�6�H�0f^?>�,Q� 8��'����Q�%T��0!��Wʹ:�4D�� B�yU�1F�6��g +<$5E�iK�𤇝zӘeac��	��`�ޗ0�az��;��"O��9�f#5;�Es5$C�$�7-4�DQ6I	�q�z]A%]5'��M(�!D��)u��rK 8���ͽ/�����+D��R�H]�C�����+C����.$���~���-W�{�b�`���5��L1�"O��Y�(�0 U�)��	P����8$�'��"=E���ˎ5���P�el9@�k��~y!�DэI�c4'<��l�31i�I���O0��yr��u�8@D��	\��b�	S/�y��T;������.�B���y"O��.drA��9s�ta�a���yr(��Y�@ܑ�-�9]��r�%Z��~2�)ڧeF $:%WW�!8�"\�r!r��ȓ!d�m���4|��c��cIR� p�l��	�H�����.Q=J�����	n�B�I��&�C�S�>J����D�qC�)/�T�k��I$kȅ���D�0��B�ɩ"�4s���7.bۦ��5��b�xG{J|z5�K�L�a;�iG�H�~�Xa �X�<a��<zZl�3r��16�z�2�����IF����}",˛biTٓ��a�.�Ʉ���yR@��N�x8p�gFT�� Z!!�<԰?��'nt z�H�8BЭkt�T��D��'4ډ��*��t�����LTڤ���6�{�I�QlH�Vo��V����# I�?!��Q
s��M�b�W�0�ۄH�-!���ϓ�hO�]W�$5���U��<���&D�|�T�V�<��T:�%ш*���sH1}"(s����FT�f���h
'* ڜ�Gc<�O��ɡ��I�w���H�ˑ=z��̪���ʋx� @�I��0V�	�c5@�!��>�=����(�g��6�!�$P�v�4��q�� Xd2�x�KP/!�d�6mu6����I�2.rܒя��/Q!���ɂ!xfnE�I��up��	~:	�.On��ĕ qٶO����U{��d�{�����7OV#}�u��s)!�DO	Τ��U&�ot�j#DP{.џ�G�dD��(���7nI>�=��EQ��y�iO�	|2!�׈�"T�,�"B�y�����;T*�*n�~�7&���M�J<��O���#��ip�P1Sz\��c(ÎN(��?��.���j��'�j�[�32�h�ȓ�^m9��]�|�H�K�3�P�I_�'	��T������3�
[c��(Ћ�,�^�*î;D�08�/�4�9 �i'�f�(Q�9�IJ��,[��;tf�����B�@t)�m%�4hشA����j��4���O�����h�f� ��>,�jdcB��1���D~Ri0�'/���óq�q���޵|R��ȓ:�H�b��6�F���qQ�.D�T�7d��v���1�lݔ��p��*D��#4冤:�jE��'��#�C,��0<�H.`����k�q�<�yaSx�lFx�E�D�2�Fߩ9���/�0�PyR��h���fM>9����B�c�<)�/�Yy�,z�˱<���� ��x�aS0Nzq�� \���+�n�yr�� j0�����`_KjN�"��5D��� ��5*�N	�$���>���M?�\�a���:dh�R4��4&^89�N�yBe�$QK&��/!���0�o��<I�{f.�gy
� X!I_0��)��]<*V�9�OH�=9���K�t2���ǜY�a��I�  ���'$�D� &���S�ԑR�BjGk�e'��j5�O1��V��Tq��K�`+%L¨#�кD�=$��@�Ǭ-�'��3�M净�Y�qO��I�H��ğ'],x�J+Ïz���!)��Wp�+�_�1O&��	1>�h�Q+�.j�Kt�u�B�<M�`xx���;+/�%E�Li��'�O��d%�'+^��7	�cYt�[��<z8j�ȓ^F��F,.E�ة3�K���5����IZ}��L<Q�H>$�x��B�̳W��t�1��L�<�Aa˹
8h�#tb��р���C�\��M�Ǔ(U��0R��Dz�T2��΍P(����$�O��S�O���ؐ�?�:��pjн	+�9��'Gr����=b�Ӣ�;7��q9pD[w}"�|ʟ�O`Ȩ�cw��Q�Ŕq1|�1��'��I�z�^}��f��`��,�%!�l��B�I*l��)F�.G� ��� ��>�K<N~R�8bѶy�%Me6�l�� _e�<�����0AW�A{���0	�d�<Q$OB��L��uM �s%JEX��L�<i�j��f��AB'�JȎ���A����:�~�?aA�Q�N��E+��֥��a	�SN�<�0`˦w�H�[a#څN�!��EQ�<Y ���D5�T�жO���ps"�U�<a�C�&/�؊��3��Ę�S�<)
	>����*dr�*#cZP�<	���	 dǩ�"�z��TT�<٣g}��<Z�g��>�F@��F�O�<)�I�(m8�zC���fl�� +MI�<��a:⌫�JO5R��<#`��p�<a�$ �F+ڸ� ��,U��-�w�<q �7'Gڙ"��,B�bd��v�<��%;:)蒈ˆs�&�����v�<ɥLӅamT��h�73�E�SDp�<�b��T���-�;���Zm�<Y'��*���Y2����ڈ��E_�<��ꎚ�7��%�aJ�	S�y�Fҩ>脈�
�%H�]������yҏ����3�Í&��`��	�Py�@�r�h9¤��o5�lj��b�<Q�ʙ�6Tr�M���
'�\�<���
�zeRUz�I&z��ѵϑV�<3�C4hc��`�}-G�B�I4DҀ�v��֔m�$i9:��C�	91��3JE9! ��Z�C�I�1h�ś���$f9Z���S�^C�I�\�9D)�M��Qy�	^��C䉩I������(5OĄ(rE�Z1`C��b �q��l#��B��!ZJC�ɱ"�NĲ��&�ڑ+��U�3�6C�	Gp�ل��D�vDʥE�m��B�I48���Պ(	FV$�@)�&6�C䉯  �JӁ�S��
��
���C�ɔ|����� �d1dM
9m
�B�	�5����l΄WL�qS����o=�C�I���csfۨ@�(�` E�6.�C�R��Iq �syڑۧ^�qz2B�9�̋�A\�+���1���>u�B�IC �%z�G�F¨saE�	*B�	/�$"����RA��kßZ��C�-[2�}z�z#����Km�B��e�ֽ鶫�`�
ḣ�ۍ.��B�ɻ��u��o�H�Ic�ō��C�)� t����9'�puC�٧@8|p"O4Q�7�R�O�aD�".�6��"O ��!H�a�v �#.�2J��9q"O�ɀ4ß�.I������)w�䠩@"O�	g�Ӏ!x�c�)�
΂����'12�'�R�'���'��'���'�|�P('!�P����S�\�2&�'���'��'���'���'���'� u+�X&!����$7i�pa"��'r"�'8r�'�"�'��'���';���J�\�J�Ҷ۹.�8<a��'���'N��'��'���'�b�'����Q�C� RdIꓫF��*�p��'���'�b�'m��'Jr�'���'Nz�y�%�'Ʉ���7sL"��a�'L��'���'�b�',B�'��'��l�s!ܕE�R�G��a"�*��'r��'s��'LB�'���':��'�����ʹ
t\��'�� ����'�R�'��'���'E�'ur�'�F�{2h[U��`��k�ր×�'�B�'&"�'���'R�'X�'^���@�v7L��B�N]��t�'8"�'�'���'��'�B�'�`FجCrBt�ѳ|Ø�q��'���'�b�'���'Dr�'��w��ܫq�<U(�d�Sās
NMI��'�R�'^��'���'>2�' B�'�*�"��)F�����L!/d�pT�'-�'F�'r��'S"�l�H���O��BC喩}'�$.	8��'j�wf��?�(O1��� �MK��׎j�L(�!ǆ�t�r��4ʛ>L����'~�7��O2�O��O67�O�'o�\�E�-j�$dz'$]�D���lZПx�q�V)L�^�-W�a9"K�1���O�U����<k$,ڴ���f��U��y��'��IW�O�h�y�eN���Pt+>T�vt��`��L؂������Ҵmzޝ*��:u����ЈC�4�J#��)�?Y�4�yRX����p�A�Q��nwV�H�*�0]U�0[)�;:����L�x��2��=�'�?� m+x�F#vN	#/r��f�<�/O��O�Uo�sc�C��O�&Q��0V�2\�N�$� �.Oj��wӪ�u}��@9�d��O�E�TX��ޑ��D�d�����P=:t1�8��RbP�#tr���$��h�r�]
 �:4տɪ���$�O?�I�H0��Ფ����R����	�M�qc\~"�xӊ�D&�4�2E��B�b?�Eb�fXr� $���O��rӬ�d�q�F@�4��4A�T�fX�u��ŰI"�4b�C�!�<��Fܗ<�t	'�(���Ϙ'$��(Fb�;e ����Y!�8q�O��l
g랴�Iɟ��	X�'!YR�"S#] ���h�|9�uW�d�IͦM{N>��?��� h%����;�����(��C�#k��@�'v��RWG@��P��"��T�b%���G5C,4���V&2j�+jN�)&� �P����!C��΄;�CQ�]A�NC6j���lC�Nl����2�D�c'�"@e�%�K%?(���	�*���c�~G���k�Or(�O�.@��.!�Tс3�C;3�8���i�QҐ�xP�.w��@�m�勄�1Q�@��N!��y�Gn�m�`���dM��O�Xs$A���I�P\���/Ԥ*��B
��}y��HS[�5/&�M���śS�B�Ɔ�MK狶E��b��u��YsN�7G<�	џ(�	^�Iџ,�I4trl=�ɝp��M/Eb�`0gCD9X(f���4�?q��?���\	?Q4��O��ɧ&NT�Z�� (�Y�b͕4
r6��O�O<���O<=h�皇t��'�i��)@�x�:HZ&��}���@�4�?����?���41�(�,�'�RP%G�A5P`r�@y葥��'3��')�iS�G�������O60n��H@_�d��e���6�'�R˕kM��'6�S�?}��5��ԇ)� ���f ���r+��M����?�v��9+����<�|�0�P`��t����
8)px����/Y���)��'��'��Q�P�O�~�S�R�A|�CTa�4D�d�`�o��D��^0	w1O>E�	�J\�L��<C����2�ʒz���4�?���?��e_���D�|����~�冱nr�ܱ��A�H�l`@V��L��c��B����'�?���?9�M�0��}���My�B��@�7M���'�Q[�X��i����$3���?���U�F~�l��U�Y���'�8:2��;��$�O\�d�OR˓vA���f���<v�Q���p�Pq�F⊼����O��d�O��O��D�O� ���<;/R0�&�ӯ&��)���W;Cq\�O���O��<�tg�������*tVR$�5�3^�LM�����Ms���?q�����?y�L?�0��'>F��5+��:�`�s�Gq�q��O����Od���<р����)�O��:�1Z��]��WZ����K�ۦe�	~��Ɵ`��1n{D��>i�`��y��T�Ǔ_¢����hӾ�d�O�˓Q;@	y(�����O���Ŋ�͂p�ԚzEH��C*H/�x$���	П�;�
�`�S�t��j$��RB�$L��JUJ���M�)O������O��d�O`��8����.�'@�~�E!L)Z�������������.u�S�'^�6�H�s����7͜�!RBUo�&�~4�I����	韬��{yr�'��"FfE��H�.JRQ��{��T�Dp7���v���"|2�:��pN��h�z�i�F�{J�B�iSR�'H�aO�P��	��0���,���qx�ɠ���h�'�:T��>1���U̓�?I��?��� R�IbD43	^�c�A��L��iL���._C�	֟ ���%��X�`�\�5$��`��(GU�.A<�u4��<����?�����DݔR� �u�I�i�P,��N�:#��D��j�<i��?)���䓓?!�~�f�Gb�7�*5�Z�Ds��8b)���?����?y+O�9҃�?e���
�i��DINְANhӐ���O��D&���O��$�/k���.��p4B��s�6U㇬���듉?I��?I-O�\R���|j��|��J��5b�0Zg)ՠH�X�5�i�B�|B�'��*R�H�qO4�餯�?&*��/�7QD�E��i���'9�	�N�x�O=r�'D��Kߦda�,���G�]�����G�]�O�$�OV`zFl,��~�压9&��� �L�W����K\��u�'9`��'���'bR�OB�i��8 ��n-��h�+H�U�"it�rӦ���O����O8�O��4�ہ�ڷ8�ɈӃN�i�#�iul����a���D�O��$8$��,��5XĬ]�3�ر!g�9v�@,Y�%D���֟��Iҟ<�R��Ot,7���%��u�tI��f����FE�צy����x��m��h�J<�'�?���oJ��z�)�5[�Z�"�A���R�qѾi�r�'���22 ��g~2�'!�jS�kJ�U��#�4�0�Q�7-�On|�W��f�i>��I՟�'K��0�Ch�)�HѕT�T�
w�~�D̩R#@�&���O
�$�<�c瞬]R�sb~FycQ��/æ��b�x��'�'q�˟|��)Tr�)���(�-�U/	_!��`ҊIџ<$���	۟8�'	�x�i>5r@-��k%L	c@��*UTrer�f�>1���?�������O����lΈ��_8r���(ǔ{xੲTB¦Y�6�':R�'8�Q���1���ħ^k�@�fM5yx� x�����X���i��'N�I��L���J�:���H�i��*�J��C+`T��٦���kx���'g���������'�r��5g��=8,�� �=
�V��C#��ē�?1�l6��G�Xz�S�4F�0EȢ�!Q��B��2gV#���Ox,����Oz�$�O��韮�Ӻ���{ߐx�"��%��$�D��U�Iҟt@��![l�c���?9�i�;0i[: ��@ۡ)M�[d<��Ah�N�Z�$�OT���O�d��p�S�$i�1 D�B�b�A/��r.G�d� 6����1����p�1�τ*����%\)(�4�?I��?a1���?��O�� �'r���3a&�?U;.�y'���v��Е�t�'Nr�'d;���1ޘyu�ޣP����Dw�V�@ !�>�'��SПt��by��գ,#^p��l�v۲�b��6�6M�O|Ds��O�O���Oʓ7A�4�.�ؕ͘�,�DH
�d� U"�'Z�'��Q�l�I�Pc�V�	L��c��6l��Y�$^ &�Z��IuyB�'1rR�d�	Qj��'���B�)�ڠ�]�=�b=nZ�x�	K���?i�x��r����I2��w|��i'��q��$�>���?�����d0���%>]���SN�򕯅,��F�5�MK���?)O���O��:���O�O�n�(wچ�"��q�Z�Y!�A�4�?�����D��R8��'>i���?��N���{�)�;^$�Hf�4x<6m�<)���?���&�?�M~����vf��$$ �[��Igh���&���)�'���B�ft�hL�O�O�@�{�"�Js?=A��֡
���mğ����1�bm�	��'��-��F���d^��[RO�|��Y����M�uJϚH���'B��'��4n)�4��%[��' 6T�P!юJ	�օȦ���NK����	�t���?��O��ӓO�H H�HNȠ�ϙ�z�X؋ش�?y���?���Ո��?M�ObyR��Y�5t���t-�X��P��IX̓0��Ԩ#��T�'#��'�$ �Mǅ��Y��Q�� �bӴ���2D�'��S�����By�MG�]�(�;shH�>��3s�O�{8&6����6G�O���?	���?i+Of��!t�BH�tN�F����6/�9=0�$���	ڟh�	Hy��'iR�V�q������C�\Y�`�s.��?�)Ot���Oʓ�?q�͵���D LP��x ��-�@�ۂM7�M����?y���'nb�T#��*ܴ

�� 8H0v\�EȖP�T�'���'v��'F�F�Ө6m�O���	7�P(Jҭƶ/X�A# �	30 nZҟ��I��X�'HR瞞��4�'���S�|=��T	T�)I�G�&u���'�r�'H2��O
7��O�d�O.��!Z�t�deo���
�9l��\�'���^��O���=K'��C�'B� t�;)��oiyR�� ��7-�OX�$�O��i���DK:RK@d��ƕX���zdC� DI�l�'7§P1�"�'"�i>���,�*�(��L�f��DjS49h���T�i@@U�c�~�^�D�O(��������O���O�)Z�Ԛ2�na���R$A2�L���G��9x�E��D�IZy�O��O�iM+4>X1:�j� Lʸ�!Ů�3SJ�6��O@�$�O��k�JV֦��I՟,�Iꟈ�i����/F������64�s�g�����<�㦐�<�O���'���X>��3��I�gv� 3�R6��O��i���ޟ��I��í��	�q�&�h� ��:뎔0F.��}T6��O�L��2O����Op���O����O��C�4��2�͏q�@� ʏ%4:ب�����I���	ߟTz���ʓ�?�`�U��pJ�T"���.�?G)V��' R�'�R�'��'��5�gFe�|P� �)yG+@�t!y��A5P�X�Աi��'N�'�b^�<��!2��8Z������-y�������m��̀ߴ�?i��?1��?���9��i���'�p� *��UxTBTC�7{��@gwӂ��Oh��<��=�D,ϧ�?���^��i�d�y��1�Tg�	�����i:��'�"�'BJxQR�i�����O2���:<Y@���Y<&����A�5D�5�ڦq�	[y�'�Q��Od��'�s�ai�&��S��x�Dl	ER)+�ib�':�]�@�h�����O\����x�i�O�3�t��i���)4�m m�[}�'�np�4�4��']�ը%�$H��\���-q����4H�x2�i)��'H��O����'I�'��"����`7"�/b��S��٦R�#�����y�O��Oyr	PVX�&�K�Qz};�� $4�v6��O&�D�O
̂u�N�	ԟ��	[?��Ėv0h�jS�O��t�֧�ͦ�&��uI�ħ�?���?�%$Y%B�VZ�CJ zK����c��R0�v�'��q� )��O,��#���. ��G@�W��h!%HU<��c�_���N˟��'�R�'�Z�$C����ZȎt���ī(�H�1�՝tofH�M<���?L>����?q#Ί�'󊀈�HW<YQㆨċ0.*��<���?����� ��'q��3֨�) �11A��L#�4�'w"�'��'v2�'��,k�'D�E�#��1)%ĭ��Ɓh*�rv�>���?����$��\�$>($���w��b榄�X�H�r�y���D2�$�O��D+����2}��3QY*-4@Q�i[���>�MK��?�)OD����Dh�S��x��7Q�J<�1'F��0� �� ��H�H<���?�dm��<�L>�O���"��&6��y�0l�r���ߴ����q��o*����Ov�	Py~�O�rT���"ɣ�H,�����M����?��X�<�I>�~RS	_��hY�(�6%l�@'�L���А�MK���?����e�xr�'�Z�`ƢN.,���&X�%��JjӦ�;�'�O.�OZ�?����:��C̒�i����U�Qmb(�4�?���?ID�NY!�'���'���z=d�ԅ��g����N��2�f�|rꂿVg���d�O���^�0n~<!f
SΜ=ˠ��Z
�mZΟ�R+����?1������^�i�f)��j�0 C�m3!aN^}⧀ZY�\���	֟���syf��vv��*q������ٖxۺ��(��Ot��3���Ov��]�T<u*f�WH�q�I+ZA<�Ӈ�Ot˓�?)��?�-O���^�|*'`I�|ʆ 'K4�����|}�'9b�|�'8r�ȁ8���@�gTd	�5C؋-R܊P
׽ o���?9��?q+O��A%�J�YL��S��	�� iM�S+�I9ݴ�?M>���?��Nֻ�?qK�\� �F�%�YphT�$9Bɛ7bu�,�$�O� �t@c����'D���'T�X� u, r�v�"1�U�0Of�D�Opuɱ��O��O�� fYd٢��L�A�j�7��#q��6�<�U���Z��Fɭ~���jB����e�	m� �U�UM�`jӎ��O�-,
Lb�|��4k+~	;�N�-B�<�(SOԵ�M�c,?�F�'(B�'w�d� ���O,X�O�3_�<dСCf���T�L���֋�O2b��?M��gXp�QD ��q�"�'�T,j޴�?����?� X�1Ή��$�>�!��.T#rTH"R�-�r}YNU����'�jl���J�$�O����K_�[@ � ��kW��	t��MoZܟ�jb����|z����	(�M3��[�v[��
,3�&�'� �'��	ן\��͟t�I֟��%��ӆ���~�zQ��l�Bp<)�'�2�'���|"�'�r�^O�-s3-�� ���[6�:e��x�y"�'���'���'o�+��'N�E3W�,%���u�ǆ_��	¦y�����O��1���O����3.&�p��iѬРĀ? �AMr���O����O�d�<ѵ��6ىO6�9�)]�-��e�tN�?C�ɳ��b���d�O��cB�1�S�2�q��3\�d�	 v
6��O����O"�d��4��'�?����b����%eI0S��}�`C͂�]����?��	\l9��m�S�t097YT��(s\N�Z4��9�M.ON)��⦁����d��-�'���6=}��L0gnY+/D��4�?���t�l1Fx��dhQ(F]$��iب3��m0@�1�M+��HA!�F�'R�'���G$���O�1z��K-��kd�Z�Lhq�G���V 4�S�OxB J4/��Q�,�&�D�:��J/r�&6M�O����O<�#��D�����IM?�� ��7eh��ޮc��z���}�*����<���?9��X�L�5L �r7���GL��\�`�2��i�D�9 �Of��O �Ok�!e� L�t!�����z��IK:�c�D�Iҟ��'�b�9��{r��!mCB�P!��7qM��\�$��şD�)Γ��$�4�U�U(ߨ_$M��`�� �}�w ��"z�	�����Xy2�'�t���N���A�'DL�<@C��i �i���'���|�X�T��e�~X7MM�	[��b���&�Xu�t&F.8���ş���ty"�' Ҭ�ȟ��DÖv�<�b &i@#v�ɭNX��o����$���'h}�����h����-�S���
��G({��%o�Ė'>��˼��)�Ov������� ��� �F?Q&�A�+ f���x�X����K��~�c��8���\�р��f�'b�mZǟ��IB�2H��ߟ`�'a�T��X���g�:x"6"T�0�l7-�O~�$ֵ��y1���I��a/�( �3��(̰F˛������7�O>���O8�I x�i>�{���dp:@q�.��W�@�ؖ"]��M{�&������y�'L��a���e 8H4��##Y���o�2�d�O���L���˓���O��I%f4ha�㇊�_�U�7�\�9�̩��y�2�>���O���-M�9�0aч}�
��@f�3� yn�����%.S����?q������m�b���S�
8*]�Â�\}�gJ���'�B�'RW�\��m�O����Y|��|�e��2���L<���?�O>����?�P��yqD�2 �>ȖD
kW�W ��<	���?���HQʎ̧���0ƛ4G��h��+`�|��'���'��'���'�޸a�O�5��A�<�s���M�T4��]�����$��Tyr$�v���ШՐp��+*��F�����	V�������O�(c��9 @����Ʉƙ�w�4A�8��8�I��wv�-0� UH��0��b?�{�w�9k��ߛ���:&DA����'�Ƒ����-V!qdŃ
BD�;V�\�[�\U���Q@Y���[�i���YuKW�"IF�aUG�Q+�e{��Y�OL,�pmۻc���5�����0�B\-2�NM�e�Ƭf�`�9Bn�p4����k֡W�2|
�� 4Ѱ��`٦$Dp���m�
%Hq�#�Cf`x�%"�A� ����(�(ɗ�L�M.PU;T�']��'��i��B��V(A���`74	�Fd�:K ��@f��g0�6�
�V�P�(��L>	ԋ'�NPA��UN��bG�,w��P!.	� ~�7͗�048���L>���Y���=�Eĉ$Ic�a�D���?��O��������'��Oƙ�`Lm~�����JabԁC"O`L"���ݢLa�%S7�	"9O���k�����'�I��jL�&�5�`՚1G-/z�����㟬��ğ\�^w�2�'��I���h8 T�Ӳa^ �A��@D�9{��P�򭻄��NH��WB0������"�gO�2b�O�*8��� \U�$�^c�>�E��7#�8d#�%Z�*t<�0Ƌ�w�v1:��?�����'��ؠ��f�v<�'��8�8a"O�����
|fYj2F��m}@D�YĦ%��{yB�B�7� �'�?���+�����\�UG"��?9�]�\}���?ɟO��̪&O؟m�Bay�U�����*��M�.��Q�Qy�R5çI�H�џ��s�J�pa:�JD�e���plٚ8�B4�5G�&x8��q�׿,N=D�֜�?�R�i��d�d9*�ň��-H2)G�����<����<�w!R�/+-���3b��p2 ��n<Q��i�JЊ\2S�Qy5+.I�xؙ'��	*P*����4�?������/E>���`���5&�3*�`���G��=�����OR�q���:�i{���A���|Z-����
6j�V-�a+Ol@�P'�>E�*\i�ɝ�pl�l�E��<�|��C��(��P�)U�Xe)WfXY�$�*S���'��O��O�V�aA��=x��8��>Z��y��'�yR�ɍ\0m��/ځ.MDc���0<qw�I&��Q��T�-�P@���,d��J�4�?��?qC[/&�L�c��?��?�;X�*a`C?@�,��ȇ&�8A
��ތ46lUr��RO�h��ؘ��v"*��d��=��{���
��1��N��"�*A�T�7�F�W=o�1���D' �y�ݝ5���d���6���`ėI��7��Cy�	��?�}�I�d�	E`�V���H�{��
��Ɠ&BX��e���[F��"��Y�3�n�͓�?A����?���IyO�Mxy����NTq2��.��I%�ׄU���'""�'���X���|�r��"�� �錿z]�G]9�X؈a��k�JD�R���way"�ɰ1W ��Ӂ�v26�J6��A݄Ё�dJ�o�Td3To�R�E�#`�Dy"b��e��"LU���!A&v�DL��?��Fj�v���<�����'�6`91�95D*���ˑoCx i���n��E ��t���Q���6I�N�<�soն�?i*O�L)tD���~��'TʵfW�g����b��m�X-B��'{R���/j��')�)�PTR(a��	�_���Ct�y���!�f�u<1eO)V��p ��'(�h��n� ʼ�r#�"�y�Uȍ�g�<��M�~��@�5�j�����N��������D���"�{�b�oZ��4�3	�xWr��C��8A����mN@y2�'��O>�g��d��u��ԑ:(��{�!�i�4_�b�X�G�1�&@�УG������dѐGKjhn�����J��*�0��^�4M�La����T{}���'����ShL���7��%q����|,�h�0�k�3L_�e��ꗍ~�����>�B�5-�
ah��Y'�yqe��'8q���C4�6%�BBT��*I\���>1����h��4k����'���x !Ǥsa�ۅ��@F��D�Or��$�e�<��+�����䈓��ax��u����8�� ��f&ߥ��\Y��@���������� �IQpM+seL�����ٟd���ߑ����V5�ܺ���z_0�{�����F%
�/Q� �Cͧ���|2M<i$B�3'�ڰP2�H
꼥����qDz���^��ӭז7^�֝%��d �e>�n"��]�U*�p�QnX-��c6@H�~
̔x�42��2 Bh�4��I-�IQ�:� ��Y;<H��rc��G��C�I !�p�0�� ���K0��	���~ݑ���DT�9b�8�LI�8^�`�G�g:��YFEŠD΂�d�O��$�Ol����?1�����B�	vu&�����#\I����	YY<�@T�18X���G�-g��V�I_�\=b����]�����%?JU��@�+ M�H�&�E�,XM���l�'��4�g��F8jؠ�
a��<+��?y��i�O�d�O|���G��'-^ZTAAO�S/��8!+D���3B
�~��!6́�u�"Q��y�#~�.���<����(�&�'�r�D�v�����[#W�Ɯ�5�
��b�'3�XE�'��9��!ЅTf�`L�ƩJ��TJd�Q^Z\H�l��Zrn�Q6��3�p<�g)I��I!#`U2� `Q���\���YB���:�F�h!L�cf�h��Þ!�MFx��;�?i��iS�7��O]; �Q�_䶬�J,d
�#��<������|�RVF�o��M��Ȁi�2��I\���,jӠ���ID`��)"-E�S6
��)�OL˓[٨��4�����'��&(u�I�g
��j1-C4-��}�Cυ*.��0�I�K0�<�Ӂ���Tx@�"
�+��i�|b5G)*R��CŸ\֑�o�z�DM�H@`"���*Q�* +&b)j7�b?�r�φ"��t0���X�PqB1}`��?)��i��"}j�'^NZ�!�c�b �䇘$7�X���'���{r����xQ�g�:�f��Б����Ov �ХFّ��D��-��M����?���5�\90�N��?)���?���#��2
Ű�X�߽C�\����]�8���ѨǕ#,A:D�H�=	�7擯
	5� 3O���Dh�=D�����O�2U�w '_�<]"'�C>����ҥxBq���sg/���yӎ WҘ�d�? �h}x7�_�R�����N�O�I�O��P��,�hB$��$��(��U�N7D�D�ej4�}SW������ %
i���	��HO�i�O��K�|�3`���������寉#]Z)8��(��ğx����uG�'G"7�҅�f��" HVa!R�� |�3*�n���s�
�>,��,<O��쉎�z������e���Ȱ`S�Z�FXY@n[ ªU�Ӎ8��V�	�*:�`�Vn��z�N��Ԍ���O��d�O�⟘�bS�'H�\$���6iW�����f�P'�LS a��R~m�0:���+�(1���Mc�����Mn(�O�҈Ӆ�x�Rv`:���Rӫ�)���'�i���'��=����施(�lQ�>��]��8�0l��G�90h(Mp����p<Y��[���7�'��D���"w���o�kf�|�$C<.8�;����hO���'�"\�d����5�z}ɥ�;bl� DG'�Iӟ���I��d�I3
�#mj�bd`ʐ(�#<)��4���o�.�ַ~N)x�
#�4���'��	b>�۬O(�d�|��
���?�7�R�K����i�4�<�@�\��?y���h��s��c�U���^�?�Ey o�,7��\I-��=h�M��ݢF��s2�p⡟>ٷKی?��xp�E߭0��pX�EL a��QY1	E�T�� � ��4�}펝s�@��I����$B����ٴ�?I��l*����v"�]�4��!��'<��'q֜E��_@��f�:D�>8�R�i>m�� %������L9g�qYC�?$:��2��O��d�OXQ-"6Ze��'��'��dݡ`4ʏOTȸ����.P�:܋5eX�t�$x�TS�����9�Rb>�O�Y�Ń� �X�h��Ŵ;"~!@�,`)�	�阗;��[� Cq�>Y��OT�8���@����^&HJLx,<��lZ �M3�s�")A�S�gy��'�*zL�-����#A�	��+!O����XN�5QÍ¨4�[$��@���$��*�$�<����*F�*`nK�\8�s�J�q�x������?I��?Y�)�ɟ�ͧ�$r�ݖ׺]�g�G�1%8��wI�
NՄ���휵 5�
�xYp"�?J���2�U�d|���2>����,� U��!! A�Har�C�'7��'�V����n�K���&Г��((D��)�R���+Ԯ` G-�N9�S�F�h0��<��[���'��e{�hw�D�D�OkcI4J}�гC*�c4���$��?!�y��UZ���?�O)Pl����>WQx�c\�� f%G�.g �S���	,�~��Ń-��\����H����
=���{Q�9����'�D+V�(2��51G)�K�'Z��c���Ni����]�8�[2�Ңdq,�K��!F�ʓ�?���i� ��p�mZ-kRpl�㈟.�!��	說'`E�x��u�"B�<>̴0��bw���'z�؂�b�D���O�˧`H�*�S�? �-4G
v����0-?^�p�I�O���/rO���0� ǂFv����O��Ӥr�Υh'j�7��8�S�ů0�'<�@���l����"�D���<���,�R����Y��VR�(�'%2R��`����'�B����'�b��h�S�����@��'P�M��'���'��'��$[nz�>(�g�ӄ�B�b�$����'Z ���ȶ޽^LlX��Ň�M���?�l�`���F5�?����?A���pM��G-�?J��i���5��� ��'q�L���!v&H��+4�s�.�ك�z�X��e�M�VA�ڭB��
B��8}�Ah����N}{�nB�._���|2�i�<7x��n�`�b1m�Za°���#_ln]�޴u.�6�'�~1{������O�E�"-�+1��I'��mTj���84�8��푓c�x�6��e���S�`�(�Ʉ�HO�	[v��O��P\���m֭T����� 8��ɻ0��N�z�*��?!���?��]?-�	�|���ix!�ƀ:sfՁw�
�t�BJ�2༡ `;\O(sD����{ Zy�8�@�^�T`�lв$m�=��&�D�3���!׏��b�h0���۟�I���Dy��'��O�D#�
�
)�x���͓�m殄��"O |k4(Ϻk���-P�T���BR}2W�0ID
 �M#���?�&�(t��|X��9e�n�j�b	�?���/,r�3��?q�O�t�ɡ$��P��	�e@�F��U��Mt��
o����a5�p<�uj\�=
b=R���h��@[eMf�#�!�/4��Z$ ъ-}� y�b�#�Dxb�7�?�#�i*��',X�qS���dU��n�3L�ڕ(��'���'�R�'$�O��'`<�Ic� �eհD�b�M��	
�'��6�.,���G^W�!K�C�N�D"�IN}��,O����aɉ=f0�q�B��1-���"OZqȗG�	+���֡�<CpX� �"O)� �:Ũ���82��Q�B"O��Yd��X�Z{�F�O<�q"O�H�hܣ54�pP.�e�� "OBDh�B�.����g.��1"O���WJ��Y)"F ����"O���*,�"�`'%�`�"O��Q��b=@:E�w��d(�"O֙�Ch҈�ސHT) O8f�� "O �U���0,A��
L�2�"O���C2C\6)����i�X �"O�I:���͔�)fa�?jf�Cg"O�- kD*6n�;g`O7{��ڰ"O�Ђ�5���3��%^��ܢ�"OT�A�� zd�]��./S�8x��"OD��	˦'����e���&��x"O��y��� #v��B�k�3!����"Od�����ED���q�Z��)�"O8@	v�Tdd����)G�C��\)�"Oh`uk�
Y�	T�w�pDB�"Ov0;�j��Y��4�"�V�~�!d"O�X���H�l���z�{M�(��"Ob���X6 )�䆀S�����"O��� ����iY"O>#G�֮B�`��FW���4"O���^�!a�)�%l�Tiq�"O,m	��_�aƆH�cg�
�G�'�f��@�ɗ����- ��k�Y���2BO�-�|��Z�0I�'����j�
`(�i���53J�?���Q�6�g���� ���}h�y�y���=��x �*]f���=�2���D��/���a!v>��t��)!u����Ο[�b�b���w8�V���)�Ӝ*�2����e��!�f�{�̫& �9Y�J�S�g�9"�&��Q�To�4#����G*^v��n�_�dL1F���NJ�8?j�F��Oȡz@FJ� �� ��'r�4����OZQ����f B�I@d�h�����h��
	Q��i�gZ�T���
�f��Q"A�V�Q��i,Z��U���z�i3@k�X�]��A�R��8}"��c̓u��I%��b�Ƙ����
��,S�d"�F�A��%�<!�N�.�$zuA��n+�)�6MXF?�s�$Q����E�$?\�z�"}�g�	C�� �b�~���dʘ���Gށ-�}R0L�6@�[B�9:���Պ�EC�P�eT��y�g��ʷ�:Xd\%Bp�΃[�.���y}�"�s��`qؗ@����J�HO4T��Fc�b�@�Ǻw8 ���NS5z�ı12�	{�π �\�D�"1���u̜7U�� �K޵d��#k8OTԘ�dG̼#Ċ	�w�)�k�0/ٮ�h�$�E���&�p<Q��p�"h	��L�P��@�B�jE��5�g(��H)/�v�xs(P�&5��9OqCmO�0��)֌/q�����0wT��'���"MH��H�(����&:9 fA?cI��k�n��7�r��#"��1�Lɝ&k&xy'�~>#<����3)��\��0@�F8ǈ;z��ɨ-?� @2ʑ����g�4 ﮣ=�q��U��G�t�Q#��4���:Y�*�*��'t�	����C�&�D��7�!d�e"�NF\�a#�삨4u�Wy���Ǘ1���B/�##W���S�(��~�'�^�����@��	�հB�])D�i��z�X�X,����Z�`bN�zF���*��@����R�&��/��˓�~�P�T������:P퀂v9$|����O,R��]�^AH��E�2�4Y�b�����ɫ� h��͞�J ��C�<�O�xDD,�AC� �̴:�^��yBL�]t0e
&�\�#J���H����$©w���іh��w���a+ct"�xs��=-	v){�P��G{�O���Ѣb�2J ��Ά�&��e[��'������еA�QIf��l�\�p�-֍�?9�)�I��/1n]�b��!a)�b�
�XȐ� [1%��	XW�Q��J�8��و� ��Ty<��%x�;0n��*���򕪦<I�И9��I�G2��bG�|
&���~�aw�部Q%`�	��]|�R�'@ R�~x¤贳4�뇠AE}*��ƍ
t��	�n�,F�)��#�-�?A���@o��`@ဒk��pąy�'chha�M�8z��e�� �:��	�y�(�zT��'c�x��%�<�6��6f�j�R���W:�� �.��/�-���	U����	7A�|�'3
���d/~eLp��fΡ\�l, 3�Jy���yr�K���S�4�i�uHӨ�9��i��� ozD� (;��>����=7$rq��/g��a��c.��?<��H�	��P�g�E,*�p�'^c�qkÅ�;R9�`qaɜ,9b ��ԃWRr���%6W��H�N?���c�Ă�{[���ޜhsH�	'[�\H����l���ɶ��`�ˁ̚�;����μ(�Hb�`�4nP�)���N^&<`��3Ew��H3����<c�k��o4�a���|c�0��n��� �B�8F�����(�O୹C,ڙq�B5ͻB]B��ç�)�DY�"ŷ[� $G|R�[(����&M�+�R���C � ����(�H�2!Y2MғK��'�����'����oT�L|"�Ȁl�T��RH\rbIaJ"�g�NR�Q���r�� b��)� m��L 0�jXC�O	aT�K&"�>%���(���(�0�e V�C���čx�O ��Qg�'7ʥ��#��������N^.�u�L|������=Lh����¡��S��1O\y��A�F}Ѳ�t��V�i��8�ӠS�oڶ�c�f����rƜa��|�Bn(=r�嘢
жK�EA��X�md���'�I�-�M0�]V���&�LFj�]2]���i���8KcP�2FK Qu�$ҧ��G^��0E��4Q�URzrj����DT��5���SN �Qˁ� �4I'��*͐b�4K/��jM�yh4��Y5�	e�O��K�I�4�i��S;k�|���.(���BK������b��KdN�W�Z�Z��U��] wB4Nq^h�'z⠘�q�\	��z.݇_��ȣ#�XW�T�d@��wa�|���|�w�D7mN��y"ŷ{�����'ZX1 ^�Ҙ��C&�R��p��O�`�"
��=��Q�D��#��do�6���{E	�"�>P�.!�A�ɟ4��)�����$��'Bʸ�)����EB��,X�1Z�X�q�H��d���d�ʆ�	�% ����T>�ڇ�^ۼ;�kM/iHЛk3J��á����V�s�R�P�R�!glc>�Oz4R�,|��i�ˌ�#I2`��:扞c�2a��Je ��0�?���%�(s�_�a�hY�=�XpT,@xѰ�
�n��EydA�R��Zt D-l�xв��P!���@W�U�<��
]ьQꏮI�t�Y!Bг?���p?�M+&'�5���r@�~� ؓceb���I�v�����f�{�I�6=����n���<;R.�1��H��J)-��(˓�O��P}�3%�>�BQ�?�ч�Ï	����u
�<[n�9s�Fj��j�'p�÷톼s�h�E�&�|v�,�ywŅ.��hKc�[���l�OO6��(O����%[,!X��1O�= �D62�J���Ѧk�0IK>�Ɇ]�1KC�#B�@e!��ċ��g�Ё�D�A'=o����⊘WtƅC��oT�t���}�'t���&��1a���7�5g],���4.��@Cǟ d_>��4��0z(�aC�
�,t��B򝟰��y�h���>I f� 8��j���:8L|Q˲� ^��x�|Pɶ��D�	P��Z��J�p!�k��/�e�휚V�v5s@#+�$�)�^�k�{�������ұ�CfY?U�T1�aHD�uj�K4%�|��QqES�S�Dˀ�<k�Ύ�5� �DC^,}�X*4��M"�OfYA�M,�O�.T� FߜE�%kW������yR��]����%�R�O���[��L���'!.�ё�@7 ��lQ�T��b� � ��dA�W�`�;]
P���D).���*�.T9%�erE��IH��#ˎrjB����9У$�;N9�a���%I�0$�`���	��1�C�#}�¸ᐫ.�#Dt�i�h� !'�Y
u/��ӚC�	Ul�����	v̡�"j���1S�nL{�zȒd��k"qO������{�? ��� +_5V��q�FM��6fz�`O`h	��J�e$����(	�,O\��B&,�	�l�\��F.��p��uXB*9
�c��p�c�8/�Rp�I%?k>���9<ORt�Y�>���I(w�F�35hŹ&uz���<l�2dy�V�iV��� >���%3LOd=ڐMC�.�*h�YyYR�b�V�i-�;`AM�y�d<ؔES�nf*i��{R��*&�҅ж:%�|@�&��?a�h������^�n�P��<؆�˪&g�	J����+~d���У-x��hvo���'_�0�ʚw֚ٸ�A�6Тd���m m0-O�A����O��j��$�)���ՙf>�t�bb̢w��/~Xb�Tj0�B}�Ǫ��sM|���Ըo��yb�Ce��Sdʊʂ���,��+a�#��'���R�� �.}F��ª;�N�C��$a�B�"F���*����TzԘL�%T�l�Ԉ�5џqO��55"�Qsb�K��ؚ��O�$�PO$x�1틿�Ơ�Z!�Pqf�;��'�Uir��2�0�e��*?�"h��O���'�ZʓF�O���I*%\@(�4�N9+rV�Y'ٟom̤P�����y"ɿ/���MI�KC� ^�
�1%CT�@���'x((,O��АL��tD.b��ݠ&a�	��p��Y��@C�f2�"=��m@�pڅp �9O���۶k�����?��1 �O�`�rE�<�˓d��Аe�W�aϟ�z�I:^��q�0"_�D[�� ��X" Q)B�'��H���,"��D"Fu?I<�Oq�L��X"�AA�BK<�H���?ɥ��*a`��S�t�P�����CE�$��'r&��Cd-sI�XїhQ�v��!oRZ?I�͚ޟ��/�|"���Yyʟ����Ց?��:�J�2���P�A��^�W \�7���k�%?��;]��xh��w1��"G��渑�EV�@���*��-6�8q�a����|�-Oqr6۟`��%j �pɕ�.��f�ą�nl��b��A߲����M��y�g[�e���㟸5�xhÆӣ�?Ȁ�$���Y/O�ٙV�~���P;v��Րk?p��̑(o�M�c::�����.H���ϴa�����|�'ۖ�ڇ�?	rA�I$8��aS`BD�]}��A��O�d��4�T��ѯO>[t��D�Yxy�`QdJ4�ɑ�I�]�xe��ܓo/l�DP�T���wG������ƱS8E%NR�^y��IVjۨ	�qfm@�j4����`����`�*�	� -���d�1'VEX�N�%/��0"EE͠���<s��x�R:OT�c��<9[w-�1	&ME=BE�����3
�Y�޴nrM���.�E�Š�T#�H�<����=��I�.�Y}@����Lğ�s�PZGk��r���Vc��t:�mQ"�O�xi��)���	'��a(�PXCc�wy"/��*۔�J�'A�	ALT8XT�Sh�=7>��i,� QDD䃇MU�x�q��$_��l�us5&TF��@�
"Zl���O@�B��O�-��Ŏ���O�`���1x�dP�"�9�\8QԠ�!V���P'Jq��τ�O�Ι��yg�oB�"K���C��Mcb�L�Xlax�ɛ X(a�3K��`����H��L>�T��L�'�=��*�#f��(��?��}ؓ1O޵`fJ7��`��$��i��	y��)Eĕf����o.b�.��hϛVLL T�Ջ`�`��7#\Ux��v"eL�J2�'�r$	��Ɠ0�P$k��m��
�%V�$�xK�U�vl�Ӣ��0[r%�ֳ�?)W�:���w�f@2��7����r��U|%��'gF���JnuI�ɩYR5hrn�<ݰ���']��?ٕ!T����[:*�Ҥ�ى�R4j�'�|������D�[�l=��dJ��x�㘶1��9u�����{3/݁A8И�L�W�jQ���ɞws�Z����;q�g�'�
D s�Q0e~x8�����P��D=nHJ4ʄ��X����tc�����`�V(+�D���WZZ�|��:Oz����'&�`r�j��`�|�Q��-�Șgc'��Kf%ѧY�p��i��������n�9E�Ȗ!tjrF�1�yr���q���c��)��K� C7ژ�Iu7�I�b@���2�����9�Z�rN0�G�/�����G>��;�
J�P�t��p,ߵ�^��C�a�p�A��OG�~r�ɯE����i��8�������0<�QЯ�e���4}C&��t�4���Gґ��.���y�	J���"ۚ��z҇٦��DU�u�������)§6Gh�۷��qG��Sd���0�ȓ� <�tP�%�*�Cm���0}R*Z�pZ`����yR�Tw��!���� %a'N�*��x�M&H���"V�T�*��W�]bEle�����?��Ί�:�p"CʂfĒH�0`UP�<��j� Z�]s�
�%(�:�ƝJ�<���u���&C^L�1a)@�<��3�%k�3r!ȅkC��B�əb����=Be�pf�X�zB䉯R�hj"nط��`j���	v�C��/6�@�"a�,B��*w���C�)� h�#�*H���T�ŵC-<�;"O΄Qd��2mT���AF$/��I&"O�Ă#a�dΰ�paP9^�Ps"O|A���M�n{���
��9�ku"O�;�, �q�0�z�j	�o!L-��"O�9���*YQ�b)�*b,��9�"O�l���S�6��f� 3)
���"O\�i#f�mA�h��$�"R�8�"O�؃@o�������-z���T"O\T���"!q��̎mSL�ӡ"O@ѓtER�g�8*��0vD��r7"O�i���_Z�����.  + J�"OR5b6�Í? .�H7�$0�!��"O��3#�X`�Dڧg�|��� "Olu�G��+�z�HǈK��A%"O�a�ʆ�L�B��f��a�jȨ�"O����ƛ�/O��'U9۪�{e"O���1%P���*��J�"O��ҡ\M��U�W%� ��"O��eO�:���sW+ְ*�2x�"O���>�Z�[%J�?xB�A"O�YyЅ�6�zM*4)�9��=+�"OQ�bgvd�b'�*uu��{�"O�ѡ��/9"�* �g^��W"O>�q��Np�"K6��ة2"O���'��6l���'�=I�Pɣ�"O������5&�����/�<\�"O$d����o���"�)"�n�"�"OXq�r!MX�0I�čN��} �"Op�x��\2�>!PP$~�*A3F"O�� ���9����c@�)����r"O�,�B�
�9�����\{~��j"O|��e���$�bJ�R�^���"O Ӡ�X5�0Ⅸ^4���0"O�X�A����LL��|�� "O��@Wj�p6���֫F�N�H�`�"O RsH�3Q�x��͝��)2V"O�M�"N�M�f4h�.�{�2�{P"O��XAFD;��n[e��@3�"O�M���%[���֡UD�i�"O�ᛃL�hC-i�-�U� �B�"O��s*�:��̊@FQ.-�>({"OΝ�Q�),N�HAgQ�E��J`"Oh�8DJ Jx�,���/0%c�"O��@��R� Dp)����M8��a"O���LЧn6<�{dP"�f��"O���wBC&	3�  �сB���s"O	�Ԧ��1QF�r�E�,n̺4(�"Ox��3T�x�B0L �`��"O�Y�f�۱d�,H�d$��%2�"O|���l����m�Q#O7 � �Z0"O��R�5/�܀�O��Р��"O!R�U�=m�۷)��9��`v"Ohyj����	Ҙ�S2��M5]�F"O�\k�

�<b���#=dɀ< �"O��Dn̛����|�,U� "Oh<x3BΓ\�N��� H,!��D��"OpsBb0 �>�8�͌�<���"OYb'�/�2�[��KƁۃ"OJI�[�VI� ��� B�:�"O���qmи�]�	�	+�zis"O6�J�M���I�"��#^�U�#�'�1O���#�2Gv�����5Ok�1IT"O�Yy�� q���`�Xb�m��"O� *�#�]}<�hW@�>Xa6�Ad"OtJ�M�ɸXSs.�<m{����[��F{�����w��y��*+l���禑�4�!�۝i��s��*;~�	`f��P�!���+�v��Q/B�ABJt�TEI�.�!�ՕG��$#�#4�T�@��_�o���O��=E����B�LX��j�\�lЊ� [��p>�J<�w��c�DI13�O(���$@^�<�uj3��bD�Ѡ?�mqr��Z�<A)E�3�����9$TYt%�T�<�u�ۭ(J�� *�.�=�1�E�<YVC�|:�`2��F\hQia/�A�<��\d�q�� 8z�����r�<�s�G>���Õ,\�f���C[k�<�1#��*�'�_�/ޘ�����z�'�ax��ҧ$)���d�!��E����yB��.=̔�MH+
mT	0�E���yr�қʄ�@�V |���P	�yr��zz�]�C�W!gƀq�|�Py"�
��d���TTm\p FIRO�<i'�Z%z��"A$Ԁ~9��[�
ZR�<Q1*�<c۔�[#lο�����@N�'�ў�'7s�d�Vȁ�&�;����a��J��c�yE�5�B�]��|��PJ���Ø� {�5�#�ŗ��M���t�H>�`EM6����ȓ+АYC��� k5�ΛYS`	�ȓQJx���̿r�r����FYhA��B��1y0kĳr�aB�c@�^W���EJ�T3ak 3�Z�t��^�V�����8
��J�I�"�E�)��@�ȓ%�X�X4��({� �Y��܋F� �ȓO�v���Y1�������Ѕȓ=D-���H9+�*��&�tRL��ȓj����󨗽g;iᱫ_�g���ȓH8@CI�\ ^�QP�ǐ����Wy�,����50�̠� �	W��Q�ȓ�ح��ߢ}M1���Y!>����k�z5ɲ�M3�J���7F��X�ȓ2G�D � ��(A �ʧ
�4�Ɇȓb0��P��hѾ�Ҁ-��nRQ�ȓ2�:%�G�	\�H=p�n�S��%�ȓ7��t�U�L1T~f�����4hمȓb�-b�	�cx"�CbZ�g���ȓ�f�Ð̈O�r�KG �s�Ȇȓ7�$� �G�7�q��4{f6��ȓ�<x��us��ڔ�Χ�R���F}*}i6���1z��9\e
��ȓ�B��t��v=@�C�8V����[ 6��C�C�=����N�9kW䭆�(�iy �]�E$rUS&�ʰWӺ���5n�Ѳ��t�rY�/L57������LR�O��#o���|u�ȓd)���D�iR@���\.����	R̓!Aؔ��y�p��AI�Z���J��r��²�Z�j
d��q܄3C(X�g��R LU�cn����p4���_�MDT�C�
�feb���\��	���
�?+b�gIT
����,EOG�2� @0 �'O�M�ȓF;(hJV!ΉiNT�3R"@7a�D<�ȓ�d��e��#IL��H�=9p���l8��HqgўT�)I���	���;�&�CL�	a6i%��>�.1��S�? �P�,�[��)S�>W���"O8�����)p�(U���k��<�&"OJ��4怣�@��
�4|�D"O ����	і�h�Ψ:�$�pF�O���J'WpAB��\$d����4Cay"�	���(���e�a'M_(?�B�2@��0�2�Ժ��|"@*�
��B�ɏ:J���U⏭E����睞?q�B䉂&E��Pd��-� IF�;�v6M'�S��M;�cZ�+�A��D�k,HiçL�Jܓ�yZ�\�<�OJ�)� Z�Mq��!�ʆ_Ƥm��'�Z��l�0hd&X��
F�W�}��'�t�C�H�'��c�#U:aTF  �'jT���W	5�0��F��C�'pHA��-φ*��&PI#�I���y�� 9i~űc��i�����)�yb�J�P�3O�7bH�qU�U*�yRi�6�"�z�hM3&��q Ĩ�?�y�ˍ�\��lQh�P��jQ��y��JP� �G]��Y$��6�yR
�S�Zᩆ�[�"�рʝ�y�#_>�钀�4 ��|3Ge���y�FM.��D'�F1�&��yr	�7+^��uN
���5���y�ā�<?��A�����d�6�R��'a{�cݖ8��D��G�t
%��@��p>�O<���8ibv,5��5y���{�/�^�<Q�bI�=��E���-%GX�SAFN\�'�?�	�*�jQ����!H���Y	a:D��h�	@s�8h*%���!K9D�lzv�?N��`�2CȝT̅ �,9D���5,� ��M��ɦ�h��)D�v͋���qã�7�)�U'D�ta�),��1r+�,a��h�"?ғ�hO�S�s�E�"�[�b���*ϸ-t�B䉗%O\ȱP揥uY�����	�B�I�9Je��Y�y��#�6q��C�	<u|�p�X*,P���/UdB�I/O0�9�`ϟ�y�H����`�8B�ɞ?��y���:TbԘ���L�N�fC��#��w�v�A����*iu*�<1U�i$��Z$M��a�5L��S��12�QW�!�$��0*Hh$,��8����c�"!n!���Y�6I�G�E91Z��`#�yR!�$�:ɘ��4�TG@�<=�IT��Dz�i�'�Dt�D��*z>X�8D��C'��-�`�8�f
�f|0�[f�9D�`M��O_����GL��,he�5�����`Y�>�M�3"ܸOu�h3"O��3��<y0��YA���n T��8� � h�Y�#l=.Z�1�"O�@�Â�V�b5�rV�<��B"OQ�g�O�j^��( �ߛ
����"O~؀�8�U���:-�bL3 b�<��TX���>z�%RwFKt�<�u�[�2�B<�j��rg`"�AKg�<ѐ/Q'f�����?��\����H�<�e�Y6�H$�*vJ����ZA�<�E��=D���$D�+�.(1(G{�<ɣ�>E��)�lN���|���u�<i�JB�@�<L)ˎK�D�Y'NX�<�V�^���r��x��(�JR�<�F��h�ؑ3�ȧ	,�Y�'��J�<i�i>9�󀌚!o��X��Wq�<� >�qe�
�d�8��K:tY!"OT�8�Gʰ]sdL՞$F�+a"O�I$E�0t�����N�^��B�"O�����n����@ �lj�"OLUAD�� xS���eZ �DlB"O6�ڑÓ
�����G\��@��a"Of� �g��U��x�'ŉ]���"O����bS�"e���Px�� f"O.��aoP- ~�l� �~�@�`�"OB���4�0b�
���L1"O6��ƬHt������Q�.��s"O�<j h��J����Q)B�B���""Oz�ȶ�H��2�p)ƕSP��"O�񛂎�*<���]�7=�,�a"OZ���f�#6%�p�O6R�p��"O�%ѱǀ(,fd	�O�$�r�C"O�usߕ�j��Ӳ^��Ȁ�"O �B�L� ���X��]�â�kb"O�E�s�a��3R"D�]�� K�"OT�(�iZ�J��ih��H-9�~A�"OL��V�ҏ.���ɧF��)��"O���rH��2�} �k�Y�-�"OP)�a�I'Bn�iVk<v�����"O���!���,�h���j�e;��x�"O���¡v����bJE�#Ȥ8d"O�Y����_�����H*���"O4��&ǆ0���K>���v"O��H4��4$��£_�E8�qx�"O��'��#�!bF�+x��X�"Ol���蚶b#�	�2�/w����"O����?���z�f�5D7h��'"O�u�DeQ�o΁�4k�+���"O�B0��ߖt��GЉv'���V"OF�{#��0*u��fϧ9�9H�"OZ� l4z�yd'�=��%#�"O�86�t��R�Y�og" Y$"O|TH��N��,�1S�ħ.Lv�h�"O�ɗ�7 �����E�ZF\y0"Of�1��>4긊&�#�*!�"O*� p��J�����f�ubq"O~؛��Qm@���c��i�V"Ob����Q����6��^.��q"OtM�e��G�����`�qaS"O� ��]�2��d�J7:�ܑ�"Oؽ�bD%��|#���ȽK�"O�);n݋"0R�B`"G5�`L�"Oz�b4kI�/�t�Y�`D;ҁ�q"O���D@W�R]!�.��_��� "On��&�6*b�ѡ�-ѹr�`�"O(Ps1aѠ:
�!1�I=F��� C"O�����(�@�լ����x�*O�ܛR��?>7���L��B��ɺ�'F�B�t �����	���'�"0�qj�/�2��q�I1�a��'� Fj�uϨ��q��r:qq�'��C5H�A(@�
��m�����'y�0"�mh��2 �Yb}���
�'�䌛*߬��4A�7-��
�'��Ѕ�D�q��R#��ż�P�'#�p�����#P9q2A�-�s�'L��#O�>$< 1'��|q��y�'��-qcdI&	�^�z1C��@h���
�'����c��N/���0j��#��t�'@��@&)�T�l��#�&��
��� a��{�4#�H\0,M�d�B"O2���΁�=��Ӯ08�	�"O��Qn[�m��u���[���p"O�q��A5`�&���AЁ}�R!Ru"O�x��U����  �72J���@"O�eZP态 iB�p�a� 0��%�0"O8`  ��A�dl6��q����"Oޤ ��K�7�0��w�Ԏ7���9�"Or���J�-Cl���|	b"O�IE�D���M�֋�=@���z�"O�,�t��Ar��&�Y������"O�1��[�i@d]����M�XT�P"O����ڛ���*'eBF�$؋�"O��i���]˘��A���Sׂ��"Ox8��L6$v�DW���\�F�!��	��^M�3��_G�1��i!�D��3Jp�gC׳R@�L����f)!�C�dN�Z���'	2$��& �" B!�Dߪh	��Ȱ@�"�B��ٶy!�$BP�H��n;8LcPHG6S�!�d�C�@�ဎߡ+R��h#�Pk�!�W�wL�l��V�v��-�����(!�$�l�lɣ2�N�igaT��i!�d��|����I�@����*�!��ߞ/Y�����o� erwjD?A�!��O���*P	Q�(�!�B�4�Ra�'N�	a�v�gN�1E!�dO!��d@3-	�D�Q�Cl!�d�5�t!	@�A�Ka��bQ�!�dФ*�VՑwf <�-��`P�!�L-)�	Pt�@b��	j�,Y�!�D@$�v����n�.���̓?�!���O�B����$F�p��ҋi�!�d&Mt�q���^hz�2��Q<|!�D�m�.��sJD�}K��K!j�!�d@�=�I#�f�}?�;$��P�!�DQ;�ԻWFB0�x���^e!!�@�1j�	�n�k���S1<�!�D�J4��`N�O�����J��?!�d���{Eǅ�4٘�aQ�; Z!�D�7]�t��
vײ�JQ��;!���;88tx��v�|�%ʋQ1!��p$
t��@ʷ7b���d׹1!��^?����h��r|q�C8x!�2N��r� g:�T#E%E�4!�dF�6H�Jv/���$^�!�<"䡺�ީ��:�nA5q�!��	+��@��ꘈ�X��Mɥ-�!�
���4yP�N�5��y�Plنc�!��&Y��0w��1:l|"u��L�!�$@(V$��s�̈́�6�t��G%ݤ�!��ǷL@2\Aw��}�r����g�!�6�e��,(#*X�Հ�!��KO����ӿ e���ԂQ4�!�@ٖ��u��n�Q0��֤G�!�$N�{#"���ˎ&fB$�;c)�I�!��R��Q$L6c1��3�a<M!�Ď3u.l�c䎃
�b����D�!��B��}�"���.�"��EAף;f!��1�N-��
�p��Cf��<SL!��88���A�'ȗ`�~䓰k�M4!�D�������4$�bX�kE"cO!�Ċ�c��!��f�3���$GI!�˞Q�]ʥJٖ{A�u����"<P!�� T�% #'\�y�b�=u0E�"O��Ô��#m4�x��>rH���"O ��U���kC��PuAΡl���I�"O������9��̫�aҖ��S`"O\��u��WJ�b��k�h��"O"m��A�<9���2a�Y�"O{�`�1<%�00Fn�*\�P"OB����3����\�v��m� "O|�A �3����F�*P�X8�"O�����8���{T ߫G���"O�c�K�\@�e�3�گh�-�b"O�R�l���8���̔,��s"O&��' ���,˩)��:�"O�y	�E�Y��	��k]]�ژJ�"O���$a�:s�tÂ˘�.0��"O*�{��<������D�#C"O�=X���&�J�K�<�^H��"O�����Wa�i�O��w�\��"Ovu�w�7m��(bO�.8�����"O6��B���t5�Zc�X���s"O�9��O���D�r�m%Z��b"Oc�.˱� ���J�$0�"O�%�"Ţ0��X�BM��5�`"O�p��%P�R�<= q�����y�E"O*���#�_�-3ԏ7�r(��"O������2�E�����<���"OH}
��Z�x(���
�4ר��!"O�装��6�z@8v+��Ȉ��"O@�����:%��S&-ߖG���"O�QC�7m�˃IA�&���C"O�$y�U� b��&��)��a�1"O��"ӯ<Ns��J���q�}c�"OQ��o��;10�)�d�&�1�"O�	�'�ǕP��C�ٞ�R� q"O�%ѡ@
M�"���c3Nrt@�"O�� ���M$X��;�&d9�"OE`��D$��IX�o�p��E�w"Oi����7�D��"��]�&�*�"O�Q��h,>H��㗅_�,4Qb"OzU�1#^�a'�i� ��>��13�"OBDp��P�<J�9�B��:3�У�"O2Q�'�1������8qf4d"O:]��X�.�%J��Q�k�ls�"O:Ĉ�J8z,�$��4*�Z ��"O�8"����t��Qp�ΙR�*��1"O��9eC�q���ǁ�mIB#"O2��5*Ҽ	C�ˣ��)<`LH�"OJ(�f�����kZ�1(i�$"O�I����Op�!ʔ
%�ɚ�"O�ExA��Fe����Y���"O~�#�f	 !��s3(� $�`"O.}ۤ˛�|�mkU���X����!"O6�'%�0(�0�JN�!�JT E"O�y�Cg�#D�\�y�)�wY�I�"O��i���X�6�b4�\IR@k�"O��X�ًi9V�J�&G� R|XI"Or�0�\:����dC'"-��c�"OP�٤V ���7d�B5�:�"O�`�ύ&s4�}c�� ���I`
�'% H�#?��B%I-8P��'+z���BO;b���	c.Q7��@:�'A������>��*�?�* �'$ =�p	�YӔ��'#�@���'@\�+d&/Wv2�AD�f$6�`	��� 
ѓ�i��b�~����
1�(D"O�T�[��L�A6	V�X1s�"O�M��G�0� �HǮ� ����"O�y1do\T��k��Q'-ْB�*O��C��\��ѥ��!`I�u��'�(L�B͘�|~��pj��,΢��
�'���Q�I�N%�7"T1��4�	�'fBu�Ņ�

� ����'����	�'Cr �
�&���P��ٓ)[h�	�'�DQ`�, n��,޻o��M��'�eV:g貰ڇI��`��(��'3y��s�*�*��Yʆ�i
�'�ΰ�fo
 O�B���Ì�L����'V�#�f�H���1R�<Ex��'��e��nW�(�!h�$
�F���'B����Y4���y�	�-qȘ�'��͠�	4[���+���i�y�	�'.farB�-�΀�$��a&����'  U�B)X�y���	X�����'�>�����	R���-њz�����'�D�Sa�r|��!�s���P�'�<ZG���b�� s��b��-D��{P�Ն-2��e� q���`�#8D����鎸!�J�c��Ԗ��� U!D��H$�T�S�V����/vS��s3�=D����(� ;��(V$R�^sH)X�>D�����P��<B�G.\F�/D� 7��B1D��"�56 
��/D�|��t;�L�Qn�>>�h.D�L����R5�`K�n�lT�f*)D���@A�p��۵�[1y}T��(D��)��2G��a2Γ�^��'D���I�rR�L���M {�YX$�&D�����G��X�L�IzQ�?D��(�+.h�1�3,� wM��)D��ED��L 䱒 /C=IA��:D�(��ޙlchd3 ,�'o�I�57D����D�%If�1ks/_�&�J�v/3D�l���(Rr�@鑮ߖ�Xq�G3D��
 %��t�z1A���5�Z��c/D�+)ؙh,�a�I�*U�X���J*D�|���Ə{��M�)X�)-����;D�D��)q�Ư��*���� %D�T0���|��i%��/��d邦#D��3��O�9�jM���1��j��?D��+��0R�Lh��	rS�ѩ@E=D�!F�K�|�0�Q/�1Kp$,���=D���Ʌ�*���H�P��ڀF0D��#ՠY)�NH�Ձ#���6�8D������1��q8��H�w��U���*D��)&K�zz���kI6BG�a94�*D�L�6d�<w:�A���%$>>!�*It��˵菐5(Z�;'�A7D!��q$�%���L�ڱ�w'U*p!�T� h�q�$��1z��2�Gݽ^!�Dg�	�A��m ����aS!��S4R�
vC��X�`\:��P%�!�$C�L3x��Qc����P�c�v�!򄌧W�<B��4Tb=p�D\4�!��ÉBP\8���ϘM��5�*�!�$�*c��H��.2h;�T N�A!�dֽB��.Z4�]`�b�K�!��U��V)�g(%������k�!�Ĕ�YW�U0���+{,ʲ���j�!�� ��1ē5��p����u8"O� �A�6I��� /C/SC��#�"OF4��gޖ!��5��ž�TPh�"O�E�r���M6ܴ����Sz8)6"O�Y��d������$p|��"OH9�T:<8�8J�i։V�)�d"O|����(0�3�	��c߲K1"O���d�E#s쨠b�"�$l�˧"O�q����>(I(�wDн[H���"O�j�
�=]NZ1e�e>��k�"O�t��� ]���*S�(H���E"Oe"Q��P��%k�G�
	|���"O�d;W��rR�eb��ٍr�z�c�"O(4��AܞfS�q�� S"��s"O>y�w�� %Ȕ�o̻Id���"Ot�h���+���B�R�vl�A"O�ӓ�ѥ+"aH�b�d���"O$��3�E�5\�%3G�W�LͶ�2"OlI�e��oP�kDHW�-ex��"O��p0e͝~&:�
m�%�r"Oj�#�X?H.1�e�>�4|	D"OvHc�(��{i����)Z�����@"OPx2M�hs �@���0�&H�"O:k䁑����v%v����"O�\���L��E�X?W��%G"Oz9��a�3r�8��\�b} "O�����K���c��Oh�,�"O�� "�*s��4��B�-J�8���"O��1OA�tVp�w_9k�.xQ�"Otq*D!*a�fTb��I�9��D�"O>�b�f��_��pc�	rxu�"O0��� �t���	d�J�{`�\+u"OT�*�H]�v2���^�I��"O=KƎ�;�hI�RX4>&�[�"OJL�a啁F�B%ڣDO�ebd"Ox�FHU�RM(�`ӽGv�"O의u��`���q��s���c!"O\�Վv�}x"O�Os:@Y�"O��)2�&1��A�L G\�ȂR"OF��d�/�dM���%`>t��"O�E�Ţ�;51��ZeɎ�4��r�"Ov�jr�ȻW�hx[�''����`"Oj��㧝��x����K���kt"Oƴb��GB�9�E�D�h�"OP�)*�[Klxs�Ae$��u"O��x�iG�[�0�%bZ�h���"O,�s�KI� \�F�H��f���"O��1I۳c�E�5��2:�.�ۅ"OT�7�4d�H���/.�6�k7"O�]�X2�0A�:w}r��*��y���*0����u�ݯ$9l9H�#�y�Yo�|�c�?$G�٢5+L �y����,y����+!�@����)�y� ]�O�,j�U"&�\��C�>�y�W�n����A�p۪\ɟ�y�A�L0�P+"L_�hG�٢��H4�y2g_�� |ѱa���Ei�fD�y`�j5")� T�*9k̋�y�2Vk�qJb��7�d��a.�$�y� 3R`�p���Ђ�H��y¤ƌ;62!���8\@�Hg�$�y�$ҖT;���;9��]����y"��%0���Á�(8��]H@Ú �y�	��a/T�ʱ�C�-�
��"�A9�y
� ,ɺ�D�~���C��6>$�a"O�A��I�dT���%,P';(X	5"O������6 �؀���!!���7"O�i �g�"u(��bV�>�;�"O��p�G'U*�&�>ؒP��"O~D�R��M�P�ՠ�� "O.��%��$>q8E[���!��Q8"O��-��~^Խ�ȇ# �P��"O�Ԇ�D��!��܋,� "OR ���Cye`�Y b٤����%"O��f�^�yY.���c�m����"Ov��ɦ/d��e�5�8I��"O�����������㑞.�� "O0:�m�1㰬Ч�&�@�"O���a �tXʐb�c�d��R"O�����@.%����"Ō%R����f"O�Б˘:ɐt���sT0��"OXL;�ؗP <e�2�	�=�~��"OxL�@�#��TzdC��O��"O���r+J���l���p "O��2Ä70��z7�E�}$b��"O��s��^�po>xq�c�-u�R�*�"O�l��g���:�G��L��pr"Or���L�$-p<:p$H�|���x"O���S��rBd3wBR0Y<� �B"Ox ���5>�d�`����h 4��&"O���A��%OB���M�*���e"OXPiA���D�bY( �c��!�d[�i��0�bө`F����S�<�!��6V��<�נB�P�(e�R��,je!�H�}�8��n��yn:�f�
�!���q��]ja��/[��yr��q !�dA�E`:U���#k����֭�Y	!�D�oł���$q8�(�V�P�	!��
:�xşW9B1���?�!��>�� !�����$��6c�!���<�����M�>{r !����N!�ӆΥB� gaUEF">tExd"O0��`�g��!����1��U"O.D�'�Q�l�pE�������k%"O<�k�ߔ9ȎTj�K6n� �4"OD]	sW<�~�*�i��!ز"O���rH
+p�V�13kգ�Pp�"O����̚Mj���&�J0u Uy�"O���`��@-����J;|sD@`"O�h@Q�>�4�d�	��dR�"O"U�d�N�h6B�*�!W����)2"O�](W�
n��5+�7�Vԓd"O,��V�D���`��ֶk�2�"Oh��ŗ2? ��׮V#�A�"O���d	{�ȁ8F��b��U�"O( �g'�mYX�����-~�43�"O�;���+7bTd �`ę���s�"O ��2m��)�Xi��SM���Q"O��B�bƬd5����ǤM�ɚ�"O�XP��[���C��ء]��L2�"O�8�ѭ%v�Zd��랹|���"O0��+�"X���	ńBU��"O&���#�`g��@�G�?iP�r5"OLxA�C��kD�"�
JV��"O�5�EGyT
��� �J6�E�"Op!�!	�ed2��j� �h�i�"O�a�&�5%�f�i�T-~�t`"O�1' ��z�WHПE��u9a"O� f��r!��=��r�&ٽMy(��G"O�Ix �'"�ʐ�G�"\Z�R5"O�r��J'Y$�Y�z��b"Ot9-ȒT9l9����C�"On��p��W�����˚e�tS�"O��9�ȅC֐b����~�5"Ov$� +X���J-�HD��"O�C��
X�"a�#*���VX��"O|��Ŕ���aӂ��#��"OX�zG��Dhv��F"�;�u["O`��g�Ϻ�%@��D/*�B���"OX�Y�(J�"H�0�F�4� ��r"O
9�&
R��d)�_e�<"O��A0�ɐv�DE��	�4�&\a�"O��Y!-f�1��Aۑ ��\&"O`P�3�"0-& C�׭)�(!{"O�P�/Q�uZ-���V��(�5"Ox������M�a*N�c$x�"O���QnN�/�����*Z��B�"OF�٥)��N,�	�	�����w"O��KW�^�=RS�ͮz�$	 "O�AHG)YyLh�c!��xުTʠ"O:x�D��e��y��P*!�)�"O�,�%䄟K8  �T�;3v�J7"O�`A�^�ft��&Q�UU���g"O� H��W 	���Z!+Cn�"O���t`�%쭪U�H:B���P4"O슄HųM�hl�Fo��W�d(��"O�qsue��	��lrp�.�x�"O�kT�_�ؾ�Ȇ
;}�i�"Oh500c�0J�bM8�&��fh�0"O<�(�Tѓ�%W'\ʘ2�"O��B�l^�c��-���>pZ�"OƐ1v�C�I9H���TV<A�"O`�eMX�}S�Q�6̌I�&q �"On���ؼ-��4b��A�
w&l:%"O�Y@df�.w�%bGʇ9C2�R�"Ot�e�Ub2���IB�U'��0t"O�p���Y�'?4���O�u�±xQ"OqyO�;i��Y;�΁K���s"O,�4%:(�@P3�L�)m����1"O���QDU� ���3��^찼��"O�<i@�ٹp�\8�bhY�=|\U �"O�=�&m�L��4�vF^�o��TCg"O�����Y�#	ye˽n�4�E"OR�钤�/�qju� �: `��R"O�4�է�9WА����t����"O2az7�� PtD�L�g�r� "O���gʒ�n\A�2�xxg"O� ��!�H�������W"O�ŸG �8Q���w�Q�4����"O�����c;�M�6/�Y �"�"O�]��j�9,T|Q23O&n�>Q�u"O�;�[��<�b,�2'�Uʴ"O���0��|PaM�2%/��(�"O�8H�(� �t����Y����"�"O�Q��Q
/jUA�|h`e'���y�oA�gRn�фQ�����C���yB_�,��0�F�~F�E��摆�yrA LĢ�*�ɩ}>1�-U�y�C��k��H��JJ'"���-�yҮK;$Ԃ�iGj�>;6��)'���y��d�d�6Ϣ>A��s���yR#�h�fT��![8:nyVFĦ�y
� ��`3C�>����T �)���ڕ"OX�"�;ʼ�*����/� �R"O<PK6�E��p��#�#yJ�["O�+ᯚ_$P&�؊zu����"O�l����\��a��#N���"Ov��f	�Vd��Q�P�0���W"O�ٻC�V�_b6��)��o$���"Oބ�5<T@+��3
��"O�-`#��@�
$��`ʞ9� �!�"O^���lY�8{��B��9阘I�"O�@b �"B���1�e��}�$"O�Yh��S�#�
E����8t�>�!"O�b�ǁK}v�	�L�9�\E��"O����G�?, L�����N�6��3"Oz1ZF`׶*�h�ǘ-����"O.�� (ޅ2�.���E�+�H�2a"OV���D:�.�+䉕'��u�"O�5�4ԣF�2���i| 5��"O$��eʼ D��섯�d�"O���a�,zה�3�¸	�)�"O�a��Lp@-y�g�Ml�{�'=<���*T��7�	ƪ��'h�M����"@�y�ȇ$6��#�'�6��d,���(��u�ؚnzBu��'lh���19��T"�'~RH�*�'��x�tӤ!aF���w��p!�'�H���%z���������K�'��5� �B�@8쩺��2h�z
�'~5C���_Pf����$A��h
�'I���Ojc��.=#���'yt8�r��7w��ҳ����v1;	�'��b���y���jB�0nU��'��#$�;i�<�'�T29v�z�'��b-��.p�q��,�9b�'46��A� l�n�C"��N���*�'{��1���9�lh�hW12��5z
�'���K�X�.1���ׁ�(VG�t`
�'�.�YG�Mx~	�H�S>Z�
�'_��dOj��e���\�Mkސ�	�'��Z�B��XDr�`&ԭ>g�x�	�'(�-X�!P�%�0�(��4CD�c	�'-��S�ɈM�^B��*.54p��'8��cW%��@�h*aE_�U�4��'/(	�QG�3f�L���f�Mրq	�'!q��@$����{V69!	�'���2a#0N8�"�Ar�|�+	�'��R%녅	� ����_�~$�y�'m�u��1=�v�H�T�}XЈ�'�ƀ�v��!=���sg��n+@a3�' t����(�I!�L*8Ԇ�G��i�p� .N zD-)'�����U��\�E��!� 2e��,�@��4�|=x��*��P�\�W���ȓ`?�T�P̒ �R��� ����ȓ3"#7��:?^��!#M�8
��h�ȓ0E\�a`��u���(��E�����l�(VH� <�D+A"�2)�L��V�X�ʴܓ(�X@K�#�:��ȓB�.5�%��|�6}P1�ތ��h�ȓg�|؀���ŋ`'ӇGvz�ȓL�Ps�@�Y�|=y��S:�����%ʦW�D��J�@��J=D�8��Q���k���l�H̙��:D��xP%_+A0�Tb7�G��2��2E#D�� �A�MC�5(��*���lD�"OL��'�B4�����CI{Qj#"OV�q�Ƶ^8"ɪPC/;Ї"O���a
B�-��g�*;Н�$"O��H�ɉ�"mxpz��Ė
 >��&"O �+c��8	'��b�4�&"O~H˦�,��4S�e>��h#r"O:�	'�/	ZlI�J@���b"O(8��� G� ��D��%���
�"O�Mz�-�%�����F�,�Tu��"OB��ƪ�+q%:�X%lD�k�"O��H�
������K�;�XPU"O��z"�P��ԋC��y���"O>q@3hW��$4�&I =}u���y�M�2..����3b��i��y�k�&c/�8s��0b�h$�yBN�l8PZ�� �t�tCS� ��y,�8AL��JQ�f�vp���7�y���.I������ӫr��4��n[��y��/T�a;1�ThD�ҵ���y"��(r�'�e��H��>�y��#�� �'([v������yR��
D�葅��Zڴ���y�f�6�\8��‡TP!�"��y�)[�,B����̓6H0��ۡE�'�y­�^L��n�/:4��P!�4�ybDԭ�Tٶ�4ذ�1�L[��yV y��a�u���9oD���,���y����I=z�+UbԭJ�m�J�y`�)�0A�G�(qH�!٧��
�y�O޼yua���;V�Q1ׁR%�y2(
1������P��B�J�)�yBO��
���v�v���;匔�y����Xp�E�q��`j*	'�y�dʱz�� ��e��E�S"��y���+4&];�`ڃ]0T��h��yrе&$��Qf�T5�C�J�y��?RG�<��O�_�Z��BO�!�y�D�"������B訨�2�P��y"��'5*4��H���MK�c9�y�D�
'��ƌZ�j�a��B��y� �<vB���Â7�%@�^��y�l�:^E�1���:6���x����y��Fy*�x��'hD ���y���>��08d���h"�EL��y�b�A�� H�lM}3��Qd�2�yb��I���
�h�.��Eo���ydV�Q�}2�*C�3GȠ��(���yB	��݀o�	_�R�"�V��y�.��^G�|)�
��N�J)	��"�ybo5�>H�c@;��=J���'�y�a��9è�%Iw$�1�-˜�y��.6l��ܖz�L!���y"BB^����Q�C#�jd)F�U��yr^�D}�,��k�$l���f���yn�7vv�h �c}��!q�Z��yr"��5�@����C�*�d*J��yM̦b(�홰e$c�t�����yBfѴ+wz���9q�L$2�j�ybJΏ�9��1f�J�3�ܫ�y"�ٓEX���g�_^�8�@O8�y"�\�j�HQ�qP-,���Y7���y�����&d˛,����;�y��
��H��U��F�:�(���y
�  ��S�
#@��س��y*��!�"Ov�k�ć�aq�$rF%��^LA�"O �#C��oJ�RA�I�\ �6"O`��g+R�
���3�\�E"O�2���z�2Ћ �%^��H��"O& s�(/|&���/�#I�Hq"O|����;j+T$Y�m�k�����"O,�R�^'����ዞ���p�"O���fD`m�,cB ��f?�А"O@�J�n�C�T̰3	J8 a�"On�`d)A�hxb(G4ʌ��"Od�AQ���N��;b��Þ�z""Od�0��X�T��"�,�.��]#�"O�0�j@.=�a��K^�0� } A"O�[�O+c��H�j1M� ��"ON	:S��P���*	l���"Oy3�ڞ
��q�ӭ�]�xy�"O"=�� �,q	�a@UG�#W��H�"O�=r���??ҜM#�	cg�9
"O<�X ���5��H�����>̨�#"O�e9�1Sf��G�U*)�;U"O�X���	,��(�A�`t5��"O���.�?��I��	�'(�H 2"Of�)d��~�r���a�>��٣�"O]��Ƀ�W�F�Sb� j�v�2"O�=Y�a�Jt�aHC�����[�"O���C�d(]�����#ʱK�"OHa��C9}F��Y�+�Z�l�v"O�����Wp�镋�/"���Z'"O�u0�l����f˃�P����D"Oj ���M� �J'X\j1#M;D�4*���o�t!�F�
EJ	i�%9D�|{�k'���sm^/�P�r=D��T�M�K���f��֜ぢ>D���vi�6R�<J�F�9XpnQ*b�<D�Sn)d�*�i��=\�����a9D�`���(�d��6l�0Z'.8D�8�t��	Y}���?*]�}R�)D��Ё�31˖�ZA��� �2<D����X�@ly"t�˼Q�,Ӱ�8D�D(B�
'�Ւ�l�:u�Fi�UN7D�X1�%I?38������4$*eJ��(D��ǋ�*�����T��Ы5E&D��Q(�R;���v��X�h7D��Q�L�,/�qҡ��(7+`u�f6D�lx �D��b����8C$��7E D�����Qf\���G� ��X�B/?D���K�uxr�k��K��@,8�C�I),Ģ�f��p��ޱL
�C�I8Y!����:��{��]�,�LB�ɺ�i vk��b�����2.��C�ɄYt�Hc���1�(��Z�U��C䉃.��mS�Ӳ9��JG�r��B�I�3w8xڅ�R����)��{.�B�I) 4��Ѳ(I�h
-;��~
~B�IM��haÇ�9���qL޸B�xB�I�E��)H3�Ěs�<� @�Ƴp C�	�H��0�+^W��H����e�PB�I #��R!!�;l��9��GU�}�B䉕}���b �8MN� ��d�B䉯@lU@'߅9DR���#�
B�I3:(�@J]�/�B<8�FM�}�@B�	hu�PH��m��ȉ�DK�DB�	��<r7���N�"�;����� �Yұ����U	U�ؕ:Y:�k�"O��2��>d�uL���hP�"O�y�N$"*H�`�띪\�4��"O�ТrH��\��-�%ѹ6|�M�"Oԍ�x�"X��E��T��R�"On��BdY�2�TPpoג?�(���"Ob�P�ϳ�481�D�>�d��"O���tB�RZ���M��-�v"O��Ǫ���+�-َ ����7"O�L�Q�J�d�B�s�^��"Obh���o�r��*D*K�hYQB"Or�B����A�j�$k�-�`"O-�&$�l�����/�8 1t��6"OJ�P�o�2{�t�Q.: ��"O����V77�h!�f�~"rh��"O�\Z IPᢼ�p�{�j� g"O�X�$Z����@�۷nj��"O�͠RKɴ ��Q�ɷ,�DI*�"O,����̘})|ؙ��^�q	!�7y��=S�&[!t@��1��P�!��D��@��H�a6Z<)f� "�!��0Y�\h"
��35�Yc�DK��!�ЪG����F$^�m#��P�B�	'!�2i4�KF^(�y�t$
zx!�dO�q�$�`��-�Jl�C]�H�!��ыud��WJ/N��p�H�D�!�\Fl`hE�ƛ-�&=�6��!��:	i�	�P 	�Rp�1�B��}j!�D��*��K�/��S�
�ًB!�$C�X��@Z
6T�qI!"�	2!�-sr��L�: �la���& y!�$ۧLT����ЁH<t�2���
Cb!�d?HKZ�B .�*]�4��k!����>ĸQ�x!")�UB�aP!�$A2W���`��a!�a0T% �b$!�$�1��yS0�J�>.�S��!���0�����l 9��JrCE�!�$�,i��䯁;s���CȚ�D!��^5��p�D��=�*{5(��T�!򄟔$ �m���)ztd��g3�!�V�} Qӣ��;�jb	�!�䙦L$(�Y��ױ
je�W�ڥ	!򤕡
%X���d[+H_:�۰�D	6�!�Ā	uJ��$:XB7i�H�!��FRp�0`[�Ys��	w�	7A�!�$<a�겥ܷ5��AB)�	
�!���w�^]s���.e�Q(_(Td!�DE�:g�$�v��)����0����!�g֎���+���<�!��
�!�$�=d��a�aeX�?�00��C�h�!�$_�-�A 3h~|��hȸI�!��[X�L�X��Fr��U� �!��q1�г� jV��F�L�!�΄#�r�)B@D`�[3`�>�!�� ��x53'/�T�D��ra�0�!�9i���y1���vg��[c�p!�d�T�n���'�>\�ei"�¶�!�P0vӄ(9D��C5Y �.2�!�DE�N���
J%���x�郓7�!�d:SM��cT+М:�f����!"�!�d��U4L�0�LEsh����d�!��!v���F_�ԁ�E��!�D8fyx��AB-4�f)�!�$،;���"��@�=\�@���!�� f�kPL߁ì�STĀ ^�M�"OVEr�L��O�����B�<fR��
�"O6�raSBx���n��of��y�"O�Y�HZ?m�b#M@�9.:�-�yr-��h2��r�@�eԎ�X�@��y�	MnH��( �J8Xq��·C[��y�Y�1~�r6��
SG�)���L�y�#�p��=g�W?M���"�C��y�O@ltTR�� OT����.ҹ�y�c:}� �����J�T�����y� �Ze���ЍȘB����Fo��y���:{..�XsY�C	����.�y"ϔ;i����B�7MF�k%oĊ�y��c~4�3o�xq�D(��y2N_�\��q;6d��.��2�ˊ�y�!�-��	���\lzŢSA���yB�P�u�ؠ{�^�<���(�_�y�挧z2ఉ�0(v� �*n�!��,d���	��5p����'m�!��$3+
,Y���B^�� G�&!�d��Qv�ғyQ��P�]�b�!��ˌd����լH�X5D�0ç!��Z�c(I(�C�$�
ݑ�B�,S!򄗕�,#�'ïo�H�I����!򄓰?s�\Xצי>�-hAA^��!�D��y�9Y��\�)%*��<�!�P,i:���D�0$����W(��!��@D.�#q/T/K;�2��^�e!���$4������$1B-k�e{"!��P�2��U�Sk�O&��q�m &H!�d���Ӂ�Ąc�`��FK�|�!��%S3`0�㈀��Q���E�!���.� �q�o؍�&)I@	_ T!��ֆ=�y5O���U�*��_G!�d�?'���4��j���H�
d!�d��Xx�
����f��蟹?7!�6��hi��_����ك@_u,!��˛b�$����yD	C�	Er!�dQ�A��ճ��J��5���UL!�䜜m�d����#laS� �;L!�T���y�)�R��xr�$�j�!��@�x�
�T�rmC�M��K�!�X 0Y6�;�	?5���І7�!�d�6z*�!�Y���9���L'|!�dB�y�X��g(�56�HZ��cr!��Uc�I-ԆD8W�Ac1̭#�"O8׃�'5v~�{&hO#"��H0"O`�q�j��^�lXb0lA6/e��2"O���㣔�\O���b%'Qj��"OlI��X�z�pR�ƃ�Xkpa�"O*�y��@*g7vq`�@-|Ɇx�"OJ���	�>V><�`�U�A�X��"O^���kj̘q�� .1��"Oȕ��u�(�%��a"O�b�A�&{9򢯁�[���S@"O��kg� 0���0F��$v6�� "O\=A0��7[�,�D��$�9#"O"#�|\y`��?&o؁1r"O0�`r�Ƚ%K:p���Ǧ]̴���"O�� ���c4>E��94$�:#"Orp�7)�/s��9d-�#~�[�"O�!��V�&.����ڃ���B"O\�䪄�+�`p�k�4�0��$"O� ���Q4\����˒Ў�Q�"O� ����Ըy�J�:�톝cc� 7"O ��u�R�g�]#�,ӊJa�<u"O��Κ�`��W+�7-���"O��҇i�H/�U��PP����"O��"�m�*o]��2�)P����"O��j�NL���9PY4���"O02!]%:���	D��nTP�"O�Jc�܆��#�Bm��"Ol�O��А�c'Б)"Ohq�i�#�����៨����"Oh���-]/8@���/��fhȠ��"O�
$
��1V<e�D��Y܌�f"O$qs���ԛ�g�K��'"O���!��J�*)�C%u�,C�"O��"��4U-lp��P�E�
���"O،�����ɣ��6=��7�-D�k���'w%@�(���`Z��	U�,D��#�l	r��+��w�� d 5D��r0K�"(��=;�3!\��q�/D��1瞕z4�����-c;�t�W�+D�ؚs��(����]C����)*D��zqD_�"�H�9�M�����G:D����%�,���@�f׹uQdu��b7D���O�%i�Ӱ�)Ș�D5D��������x���%W)I �1�/D���2��}L��c��%��}�$D� ��d��aM>)S��[#8�ڭ!�*D�l8�AV�5I�y�&ԊsB��y�'D��h񍎖Ċ�Z���"IB�ɡ #D�  aF�=����
	�P�"�-D� r�@p?�P0�3/�<I�tG6D��"q�H)>(�RM�;]��h��M>D�x+cG
G]~e��F],��H�*D���� ڧ0���BX	ϚA� �=D�X+�L���%:��	�~�v���;D�()�nQ#2�a�n	Dth�ѣG8D�`QP�9a(F&D7%<	�W�3D�� H\!A"���&[�\����2D��q-�<;��h2�-I�	Z~pId�0D����4lTzc���Ht�7�.D�`��� �>B��C��žw5�ݸ��>D���ʚP\��+$HB�wp�S4�=D�/Dc����<,8�8��:D�,{��D �����`B�rĬzE8D�L��b�/]�q�-� >����4D��82�_�Gv1�)Z���S�=D�4S�hA�@��0�5��	�����.D�XA�+��F�b8��B��B���gF+D��%ŀ5����d#�2Y��Yl#D��Z���ei�����3xź��.D�lBm�6	�NZ<�d��-D�ؘG	�2�:�2�h֪vV��l,D�4*f��A���*G�S= y���*D��D�?�����A�t{��y�(D�<r��[5��`;�Z�!��s�1D�8[���.
V<�b�	T���1W�9D��
��X43�-I�ԢS��|K�#D�T���1r��x�(�x`Q�.D��i�@�0w �C�Q#0�{2�.D�Dڣ�E��.q�!�͆2��!D�8���N3��p0#5+m��� D��k��zr\�T�� �٘��>D��RQ�W;���V*�h8~�hb"*D�x��� ���5�ĉ��v�3 �'D�� �8ruLM?R��T�̞=����r"Ot�������&��Ĥ���n��t"OtP���p�
��Dأr~����"O�P��b�+���C�=nh>��"ODM��X�-L(��dMʿ	_��B"O��b���*a�6$�"� Em�"O.��r_*{u�YU'���V"O,�J�.�e����^�<�.�`"O���K�	L��朁5}��J3"O��r����H�$�Y��|{6I9�"O6�墘�>Ƹ�%��9Ag�ӳ"O�I`� ��fm���)8^|S�"O�1��l5wM`(��&`I�*O���A*��lri`��Ȳ6�d���'WDt�"���!��U$2}Ј��']d�S��6�a���څ@�2�8�'|"Q"	���<X#�
�����'�.�S0OL'<{�h�1MA)W4p��'B��q�6j�����b�x�r�'�Ɲ�s����Pӷ/P[.Z���'y�m�B4bH���`�]zp���'��	� *FY^zg@˒~�}��'� ٓ�c��NR+�f��Zy��'	(!؄e�2v�6ǈ�-^���
�'������
�mr�'�La��'���А�=��@3#�\ɚ�A/OR�=E�� _<C��ܑ�)�1���r���y��P�,�&�qqˌ�
�䈸g����ēGa|������	�N�?F�ЦX���'�Q� ���M;���1�@LaF�θhr͚�`!�DF�P��@��ԅ1\�q�+�;!��/��:�选Z8�YV���Rz!�ć$�.񆍚�[(V�	�ԿpO!�$�7phZ7p����W�Q9!��_�c�0�d`�5\�:�kV.1!�ڳ2�4��_�1C��S	�tt�B3O�$�!���M���I�t~�""O��+Ф^G,m��D�fX�"O�e*��N8�j��-�"S��WO<Q!V��h.��R��,|�t\�'D��BGM�al��3oU��j����$�O�˓A��I�3�ʛs���;1BĄDc�E�ȓ[��8���Q�8<0���>��<�ȓ	;,�:e��[o�sS��
c�}y���s�4 �-��I��C�BH�*��=�'�(D��R@FËKp`	p6c��<{��j6�%D�(�@"N7T�����$j�Ihc� |O,c����
� �(��C#8.\ڔ	"D��O�sv�c�,�Q�X0�E ?��O�b�"|�giv ���6鋷1�xqkץGc�<Af��Z�����_�*���a�<�h�-`�Z1 gMR�k��웦�Y}R�'u<� �#�#z���{��K^AxHhJ����IE�$��"�08��	�5� ���B�\;!�Xn~J�g!|N�(�4 !���r��M�C&���6T�`-��e���iSj����i78�:4����	�!�Q����:���(V
Ε�7 `v�D{���'��r�f&VŒd� ���(��	�'�f�zch�$f����靊ڰA�'�$�֤����_�4ޝ�
�'6�|3�jBRS ��t�L/6�È�d+�h|��i�$vbՓ��؁V��5P'"OB��Ĭw/�@���H�d�8�QD"O� D��K�++����Ǉ2@$}�a�8�S��y-Z��jQ'�=r�s�I�yRΐ �*��/ׄ.2��p�O���>)�O0Թ�0=uH�:�e�/ؕ*T�i����s�4�[��Q6#�ȃ#������Ie>I3ӡ��s�$�8�R�I��`j*Of���P�`�ĉE�»ja4���	a8�D�d��-i*I��O�gO��[�+D��K˜2�m���_�mP"� s��ܴ��>��O��<�RJ�V�RŸ�L�g�����C^�<����n6��W�φ��5I���Z�@m�Ʀ��g���$�1p����E99�ୄ�`��p�ЊP/�'y#RP1��D�OZYFz�O"$t ҍ��k�Q'&RO��p@���k�(D�$�i7���8X�);S�=W���'-ў"~��	�/<E��H��Ǆ_����T@\b��ĩ���<���8|�qCl�}�d!�u��0֔���<iN<E�K7z�����,Ӫ^�dh���O��HO��'�B�TJS�jT�:0l��D���	�'6"H�!�ҴQ��ڷ�ųs�V��	�'�,�H$�`��,^���8	�'�.<+���� Bn՛c�P��Ѫ�':*y[G�N%=[p �vbM�C�@t�ϓ�O������bS����ݧ(�j��&"O��#-�!�\�(#��i�D�"�|��O����<�. S�*%��j��S�֑2�n�G�<�40!� �����a���!d�M0��,�;�S��P��@:pC҂T�X�Z�N��_k��<��4�,?�G٣eE�q"�`N'<'R�8�/B�<�2���/x�L	ci�],ИI1iHצ)3��Fy2�i�DD{�OF��
���Bs���2�H��	ۓ�?N����J�b�L�p� �|^�pq�%���O4�=��ɞ?�D�P�8����K�<���j�n����%��!��HSI�<��g�����e&��cpKC�<��b�82Fڵ�T�ҡ9�`ػf�w�<I��݂,����� 8�@��	�K�<�"�\.���o�	�&Р�[K�<�(��"�e���ȁ("v|@G�G�<!���4b2���K�\D>�F��B�<���'��*V(ǝ"�X���z�'%� F�t��+u
��P��(;�P$F��y"晕F�p��&�_���S����0�S�OF���HT-:GzM�V�X��S��M;�'�����Q쩻�l�$Q:5Y�OD�"a/;�O��h򩖫.q��WcS�shH}Kӫ+�S�O^bS)>;�h�b!P7YX8�AM4�y2�T2CX��c1�
�
�(<��0�yB��j� MxR��/{�D94���0=)�B�ڐ4<ԥQ��+v���T��hO��$�9���0	�G���:c�+�|D{ʟ�,@VgP�oGr�FbF1 _�xj�'~�@\��cnևO�BE�f�K+���ȓN*ب��kI�hI��0�V�\t�ȓlئ�!0
�l�#��-AllZ=+����܎d��G�3����cI_�N���j�����7D�F,[Fo�< ���D���y�I��(=>��خOz(��s�-���6��O��$Z��F�+� ���\%����N>D�L�0�΋d� � �+<&u��^_~�xJ?�8�dd0+F�W��	�|��'ғ?��@m�K���"��%�a��U�6�y���y�EO���03h�J� ��Rm	���<q���(Y�\���F:�d`iRMe!�� ��`,��T���㉝{_���sW�2��'m���p��AE׉$tPD!
�'���*�eH%Tym� �]0�T��	�'G.������8���G��{��k	�'z%��#�-BO7�0�:�"O� ��!����3��t��1!"O�X�eM��	�p�P�/F�q�PM�"O� ԭ �-��uҎQ���"OL)���'2�rL�Q�ܭAL��"O>�8��:f��kf��[�f`""O�d��Jʾ"7�	q��
�`5H�H7"O��X$۠Onv�y�	�*	36��V"O�E��e�3.Yl�p�� ����"O��ȣ��	x��=D�1#ێ� �"O�ة���W����2�Ȟ-ΪH�"Oܕ���	�pZ��F��&V��A�	�'� m��� >�Ri��ǗU����
�':l���"Z��
���(T��\I	�'HRD�%�M&l�\Q��"T�L���'.<��B="\��X�BΏ{�-��'ڴU�������B�^H��'�� ��n�0���[�^:���"�'��-��.xG�(�1�W�t!t��'�<5s0e��,{b�@�jB,}�H���'�����f��mQ҉�&�^�'I���'��!��H�-v �͋Ia���	�'���2��Gra@�x£�0�>�C�'��d��̎��:Ǐ�z?�	�'b��ù��A�(ۧI�rA	�'O��;rO0lR����P�<�dA��'���)v�	B����u��]�ĳ�'��	*@٦�4@�V�ϔ"���'�䲲'�tI ��Z��0�	�'���+�JJ�D��b�nG��b	�'�}R@�H'T�Y���݁I�^T�	�'7�hã�D.
#��cG��=�		�'~�A�3�J��:G���}�(��'�(
V���e5B�0^8x�y�'Ǿl#3��% ~$q2WiC�:�rE��'�&��F�,�67mʿ-B~x{�'�R�(n��@됆�r�3�'��	�ʌ1^�6���E7�j%��'� @��\�Zf(8�a�J9��(��'?r���lC�]:�q#�h�paQ	�'6 ����~s$�ؠ S�j5�y	�'���۪@�!���� ���	�'zH��pA�"Ap���p�K�u�>\C�'���0�ۑ4"����E�. �'��<Qs�T�8��])	�g��Y�'��`zȝJ2�-�G�\�T�^��
�'�h��bf�*9� ��I�����y���
��lG�)iX��s鑏�'$�T��V���A�6|/�]�
�'@���&��7%l�S��͵o��Y�'��	8���D��A�P�u}��h�'H�b�hG=t
�AJdѝv���'[�Y�/)� A"�$��F��'�zĸqG� t,Y�c�ڙ
e���'��1'%�()���-�7����':rE���Z� p�Rg׺�l���'�ޙ�1�
n��m��G��HH��'ޤtJ�K�%cVB�y�
�(J�@�'��aP'�B�jLsd���+�R(�
�'���A!�;hT�.����=�
�'�A�$O�#E�a��h�$����  P$�aCZ"G#�M�HP��"OH�SEᏗp���1"����h�"OxŒ"�	7wy�BΟ�%)�jF"O<��%hݱNA�M%�Ñ  �1""O�8�é��@�	�cI�>�� q"O���̌:�<���AĻ%�)�5"O2��F({#vx@QE�ah	��"OTMs�Ÿ{��)A��ҧ>� �{�"O�x2Ul�4 ����CܞeP��T"O��IæP�O#��+S��u� "OR��� ��(H�Қ���2�"O��)��#a���뷤��K�"�+�"O���]26u�'�+'���%H���yҋ�-�Ey �	��X�3Ҫ	�y��6_�(�!��=��*��X�y�B)y���C����ݩ�yrC����x�"��	f���f�G#�y�� H�1X���;o��
�jȍ�Py�βOg��5[ v�Z��JX�<��̕~ j���:���3�U�<	4�ݗ{��E7�I_�N@�di�E�<	a�/3�:�a�%�+FIƨ��n�<�s��>���@�R�]݀u�E�8T�L{�5��9E
6'6DS��4D� K���3a�a�A�+(��T�B�4D���fвQ�V�`�#��e<r��Ԭ2D����,������m�����e3D��h��I�;jB��f�M�vl�!���Ӌ��'PrlF�,OLb�))� -�s+ٱ��� "O^H#S��S�l��"�̊"�*t ��ŵ1�d� ��t$��D�W�4��@�7 ��1��(V�yA��>�玜4�R���ǜ�O�b���L�<�,()m<�rd'D�0����OI�F�&�ʲL/�)�S�_�"峦�Ъ3�"�����!'lB�ɰ%�b��:7h�s+���%#a�� ��>�X^*
��j[�5��������'x�Ⓙ'X�<��c͢�c!b׀:%*��d�"|I�93�A�Cʢ���%Y�l��zℐ3il�'xܼA�$b$���G3P;.ũ�'�4�)�@� s���"&��[:����'"�]��Ǐ�>�� !�N�S�T���'Rt���&�2�ڥ+�4H�pL��'*tR��Y*)���#��^�H����'�P	�3/(8��� �ըD
����'t�𨄫S(@�.��ߞp�
�'Ϥ +�B�Y�c�#QV�!�'qj�s0� T����e�(Vfh)	�'J�H�Qa�� ���D�S�M�H���'K�� R�Y4$>
4@�)��7z�Y�
�'�,�&B�(��R�ݧ]�Yh
�'zt��T�Q�c�$�p���'v�
�'��b�A��[ �A�Ր~�>��	�'gҹ�K�{TFm0��vR����'񶄃3��2gP}�PCۥln�9�'R2$�ČҶ6�6ؐ�CW���0
�'7L12㴕"&��2�	�]�5	�'F�P�g#��!��[#�ɶ�X�	�'2�M
A6~e�H�2)#U.��r1���*k`��~&����ǆ�w�εc2�?^�di#5���ħF�Zё��4}#�<�d �_"�y�@�����$�b�a���D.U�J�6H���RC��,��-�.��O(��`�B�H@峓�.��H,�	�nH�{�Z�-A�	{��J>Q��n����U*tZ"�2��q\p�%�¡H��ɕ��Q��b/:I��j�:,r�|ڲh�4v4�DkYx��d�o��;�|P��!N����� �-����4���p��������Y8T ���O��A2Ak�"_�响?9>�ӧɅ�7���=CȌ�HN���cO�
C&^����U�{v�T�S�0p�۷^�x�&bP3M^�p��˂T:�aÕ�ǟf.넡5}��U�:��S�v�>���;`�6����ܼn1�>aGJ�MWܝc-B�OS���P�u�:̚��ю6@ЀT����M�F)�?��xK�����S[�g���mM�We1t�<�`�du���(���c&Nߤ����F�v�4���*�ӛ^A���R+�x�ZQ��ǈ�fNR��ed+���5?~a{�K�<~O|�+��J.<�d��FH^����WDֹt ���N�k���(��9�"�:'�5���. ��e
[��e�
��*rd��I����$��*�����Մ4(��ɑ��|,4��B�+�@y#���S ��GC�(����T�2$����z&:��ʟj� �gV=P�p|zÏ��&���A��	�yj�K�n�$2���9RO�a�z� ��%6M�)H7X�R �B�R�4�p�Q�k��l��>O*=Q��3}"�W�\q�@�2�E
�\YN?�s��2'@�(E�ɸ3w�����/:W�"|B��@�A��T�Un*u��
�N�8D:
<��2r��`h��d�73J�bU��v��X��ɻu�`��A�T�pG)
�|���ї���iR�IP�NG�,�� �@$$\N�s�`�&�f���C�X؟�C9K�����Þe��!,��0��kҁ{����O2j�컐�'�,�'o��,�O��:{����c��L�����E�_�ƣ?Q���&�%�VZ���@X:�V/tD���ھj���ғd�x��b�>E���<_B ���Y�Cf<��e�h���'��pJs���Ҽ=�O>�ԍǆCeԫ/Df�2�S�m��:�`�<{&f$3��'��cQG�+R���� ȅ�h�LX��d�C$����6(D3���cȆ��Х��oװx'~ � �y2�T�����ľ+�0�QQ���hO�E(�D���H����ß
f���$ЌO����"O�(Ѝ^���9ؕa��pz���"OV�h%��0��2�ϙ;���&f�W���A�'������l�~p�W�W=V@�[ӓD:����K^��D�+�ⳉ�xTcu ��!��30�x�J֭��C�F�`���?I�'�L�0G�ޢ:N�1G��J�#�� ��O�|�
�q����y2�>��Ya�K�y�숚�,��A0̓��=}�ټZ���6sd���N_3F�f��g�ϩT#�Q��~G���10�p�fG+���Q� |[%[�7�OL�A�,�S�D���]������'�h�TB�Z����'B �����0[)�-��H=^&�j�y�p� ���MSU	�P��;'`������+NA�I�����BKσV6�?�b��E&�������L2ؐ#�	v�����=MQ>�j��Y�j�G^+E��4��L�/5�� H�<Af�YG�g���#/v��:�ׇ_�01 �	�!L٘)���/�|i��]�`G��'��ɹ��$f�)6�T�:�0�K�O���pRB6OLm��I=丧�?�I���!!r�`�g� �}�	�|�4B���-v���	.1� �6���"5�P%�R�:cK�P�	$�X�����M"�@�*sK7������ҷUB��B�/Z�[&ZC�IZ�k3�_�D��U��ŝz��p���ɾ5$�x�IU?95eK�B�A!�����~�4%Q�8NbKL��X���K`��aR��c�<W	W�t��.�������?x�XR���!�:��c-��a�X��'��>�I>u\�hd��h.�Ř��D�=0��&���f�^�����=�'L^J=�#�Q�]1�h�sÞ���I#?$틵#481��鉌8�����Ä�]$^mrt��2}�\���H9�~���Wƀ��&��ĪS�T����V��C�8�S����H/��s�DPʶHc�'�2�A	�8<��6�"o�
 �6P	(����3���k$)�'�NPIE�;	�Y�O���LȂ��ΫD\�@q�FH�Q�*�!P�,	��O(��ĭ��*d�`��
�'&��:���b�����6Noj�!R ۭ*��:�H�m�)��@�#[_�Hq���m��tB��s�vl�k�)"��rmTI�fd:��O�\)1��V��f�<k�K-M1���I�H=*��dӅ@J�!Jb����7�W���J�o��V Hq�HA�-cbU���h?�B���C�EyK~�=	0��	M���q+JT�DBFkܓ!�Mr��ԂU,\���� �+$��&AV4�-#C"K2.�q2��S#K`�05#\rX�̒�#�3v�!Eaل@�Y׍T.6
�[Ç���d��u�cQ:0|�A��؇F�M��5`X�S9X$)Dʇ/ ��,�DK�y�U�0`�Y��	'x1�pe�5:�^!1ӡWQ�pڇ��Q�x�C��Ox�9!��{4�������.���-��Y�6,Sv�'�l�c�סǀ`׳i�	��0y��Iփ��<��ARB��9j.�d�g5ћ�k�&��3�)� X�%��,�,��h�&6QD at��+*����,"�����$�@�-'�0Uȥ��?{���C�D%�4�"�ӇZ��ԋ�)�O�DJ�ƍT� �rd���!���8c�%ggb�xUK�myR�L�"�����/�1�Ef	�l'�;'���	�i[3�Ҡk�"$�6�ȓT�< �]08�j��f喝#i��l�Fڼ�S�5ޢĊ�M����:bu(�:C���I�Vd� �"��Yzd$��=����FDV���'+���@�ßW*����ۯ��z�b	
%�^��պ�+�!��3�	�upc$	�����èC�HX����FV�z��O \���;���:g6�b��qO�е��>�0?1�dP�j6�(A��$�B�k'�B_�'��E��iG{/q��hw,S2+��9� *ŧ8�Y�E"O �v��ifrH�3/_,��\*@R����O�}�qOQ>����!t�~ �cm��L�&�xc�#D���5䘍[�Ғ��S��0+3(?D�h��B��v����.q��0c�I<D��ҳ�ے3|�RO����`��&D��2��ɓX'h��`�T
	f����%D�|���3�h� �e�B��-��� D����@�՚��P�D ���$� D�𠲈T���9�L
RGv�j�%?D���εG ��r4����4�3�7D����
 �D
���UA'�4D���cE%z��0�f�.��l��&4D�P8 o�ac� ���7^3�P03l>D�x`@�9����a�$R�>e�u�=D���w�� >���/!��A�k=D�{�My����ULL�c��VL'D�òH��b�ر;��#v@P0{Qc"D�Ȩ�-@�t��ɻh�w�t+!A2D��6I�cV|�h&-& ��c.D���SJ��~���҈�w�ĩs�2D� HPEZ<n�8}#�O��f�U�20D�|i���3ԁ�JY�G��ԛQc2D���G��Nh���*wf���`2D�|j�	�S���dDȢ?D��	%� L�"�f[$^�D���;D��iP嗣?��P�h�8���S�6D��C ���̡j� J�b#��y�-(D�@8�Z �4��S�Bx��Q0�(D��kg��#����pL�Q��x��-D�\��g��?ޠX�"�Ӯ$�d�A�A*D����W@��#�Q�1�4��g�(D��.�#<aԒ%�&: �V�'D�D���5\���N	_.�Ya �.D��J��R�RQ����� �嫐H9D���T�h SG&���!�*3D�
�oJ"�V�)A�Xd��%��'D��Cr ^3Xlv���$K���2�$D�6E�<+�^xǮ�)yOJ��S��^�<y�dH TR�_ W��\k�iZ�<GN�B.(BJ	�p���i�<��O�/0��c��� =��1�@I�<���8bm��pd��_e^�y��D�<�pb�5�mR�mU+5�.�A K�o�<Q׏L5u�b`0��נlW6�YPp�<Q&G��j��V%�:<�Ԭ��AVg�<��[{>DiB�M�m��a�׃�`�<��&�lc°I�9y�r��x�<Q��ԿTj�,��K֞H��tR�)�a�<�g�WyJ� ���.H�́e�\�<)��-&n�(䧋
zG��Q��V�<���̐x�*@��iY	F�)i�oML�<���R�{��򥛄F��}X��f�<D�Fd�試ĂQ
1�a'�I�<� Hˡ�N�`Lt��`[�<�Z�0r"O��Ae���[cl�S��S�R�x5a�"O`��@(Ѣz/���ƣ�?u����"O��K�-$��`�DQ�����"O�!kQO̧P㊅�s�ܸ��I "OLp
�j�J�İ���̮1&����"O��K4�͉fu�y��놁c/�*$"O�����6�L\����M��y "O`��b�#��Y�R�^|���"O�C&�"Kچ����M	e�9p2"Oҍ�D品����.����(u"O��`�2v�\4	�LvD,T"O<(�7!��Px���yRZ@�s"O�rTj�
�%cqr6�Ib����yr��!J�ē�.��kBT}�P�%�y�Q8-/��H�[��;��§�yr!��JQ���5�DD$�i�C���y�Q0�R�ag,::4�@�#��y�'��S.�x�S�0,A�� �yBFW\���F:( �m �C�,�yB΅		N���+N.�~�4I_��y���_�ځj��F�)]�+c�Ü�y�%P65�8���NX�"��5+S��yBɀ�w��5
틐��K��yRK�:p�
Q%�!af��y"�ԅ��$J������� �S��y2�ŉl�d5��ԨE�� h ��*�yҎ�<_�
�/,��3�,O�T��'�ؘb��M)F��-��.B�(ؠ���'�D쐖�n�zA���;PFBT#�'P )�d��?���0˒
Z����'�b `tm��ih:�)U�,T�x5�
�'������L ,�5Ct��U����'�p�b���l"`��%�C�~���'���� ԫ;)��+Q�=~(�3�'�^pK1C�_��cܙO�����'z�ё%ƟF�MӃn@�?�y �'����"�^�2�	r[�]�>�H�'�dKJ��1 Fd��L�:?�H"�'�,�:	Z���'��.�d���'���q�j�'Vt*\�f�;xq�`�'-�mF1s��QI�"G����"O���8��u����fс�"O��9"�2X�Tp11�@�p��$�U"O4rː3J����j�n��c2"O�D
(E��H�u�K�|V��A"OT����>tD�)�UpY*��t"O�Q��뚾	D �%e��^0@�V"O �hCL�:Vؠ���@2p��G"O��R�tż�s��io�@:G%�[�<1'�@�A�FU�ЎָMsZ!��@�U�<�d�	l��R$?�0��KV�<�sFI�P� Y���;����$W�<�gΜ	`��Yc�`�=�$]�B]S�<	`#M67�v�1�j��;�&��u�r�<ɱ�k����E�:�����\Q�<��?0[�x�5��!c��P0×L�<�T�j��!Ѧ��r����N�<�� �z�yP%ΔlA�}��!T���D���b� ���ME�e�� 1%a+D���������vA_eG�P�U2D�H�Dمz�,=���%'����n%D�zӢ4Ę-!���6��	�'7D�$�Wd����ևĬC8���!7�!�MÀ�π  �!��-F�|�ZC�?N�,q��"O&`
R��r��p�!	�Ҥ���B�"���OЬ���3?���V�8 �yJ���mK���v�^��W���ө٭-s�|�E&3/�M9�g�,t�T�y��)(
R|
�b[q}���d�4�!�"$�8�yZ�(5P��`��Y�)G�i�)O�H�O@�y�!c�Q���'u�R�&ý	�p]r��N�ָ�
�'����Q�t�6��,Y%z�kbI�?(��rw�SI͖u��"�>%���'��1���?��t��
Od�"��ӪZ���롫&\O��4��6}�n���Ӭ#���f?�� !��I�.#>�)�B#k��'_L`(���>�R�S�h1�@Lf9X��a�oܓ"m�pf֖4��� +���0.���cF��=y�1����c4P�"��>j 5�G��a{�f8v�D W�.�F�"��I`~�����t�����'��P�O�b�%�P�%�R�2�M�p<���q��1�DH��!��W�� B�"OpaȐ���FLN�sA�!g(��E�z(
�U�=t�"f�Y�|uؐ`ǣAA��#e�Ӷ�,��'Ó�0$@v��4&����d���y��30����Ț�.� ��G�O�!N���Ǫe����"JQ~��I�'�t�r��h��g�F��Db��9�\`q0�2C+�$ ���w�l(C'��&+�(�e	(�����L"|�m�� � [ȸ�2o�.����$�pp���3B�k�v�P�_/.�J�!W'=&<��.O��}��b��XR���CN�+�>Y��n1G1�m�H�xL~C�I�C>`A��S�T�J��Ȁ�~]��ă�:=[���>�?��%ɬO$@i��3}*��+T�NnD4�IQ�Ջ�8|h�"O� �#n)}謑�BiؽDcm�Ǌ�;�F��'Λ.��S��?	g�Z�x)b=Y$��jCXMy�	S�<ɶ(�*L�J5*�n�y�D!�,FT?�u
рt����*)LO��sd�V�s�ځ���+L�aj�'�넎�y�l͙���-K��%��%AP�`�"D�8Wk�/*�0�B�\)̒(+w�&ړ��݊�+"�'{�t�[��>��7&\1DX�8�ȓN�P�JD�ʖ1���u��.5�L��"�4��R7w�@BHG�P��� ڀrB2L��_o��a���,}�v����� ��	��t��.Oy"�3:p����+@��AQhP��y�(�u��c4K�D �`䄀��� A.�8D�*+��#�B.�#c�m�s!��
Ǵ5Za
OK�<a&�̒]9����@�j�8�Ձ��c��-X�F�.<ɏ�L��Ӈ� a�|Y &�6Kw��5� 4���p��0O�uyU�����	��e^�,�!�Ԁ�Ta}�,a�P�@ڴ&.�Ѫ&���<1� 7#)���VG�>�
^��D������u���u8��z��(� �n��S��b�JǞ{32Ble��O4Crin�E"��	�,Nxzuk�AĆ���QJ�fc��C��L[������S	)�N����2}`I���(DbԈ��V����Oι �o�fBn�;T��u����e��
��!XV$ƻB���U��~rI�/��ZV㛳,�٪#-�.T�����[,d7�d�;���J�{J~��,՟~<��3֊�,M2`�!�e���ɧÉ?f���D�[�����	�%hb�:1"!:H{���UR�|2����U�2� �-�[9�m����y"m��fV4M� 	�$(�*�Px� Q�S����ϘO	~��b'۴-�*�)U�>�����O�y!�a��Lj�逶��<���DT��'rBQ2G��1ԼЄ�'�:�;"���<p����M�>q�mY�;9H�!��10�̺�,ΐ%ق��S�7L��'A�>�I*2b��i�/	��d��ҟh\p�$>J8��1Ns�Y���,�'�p���90,�"bw����y� y�P�ђ��%��Ɉ��9��P- �aPŦM�/@�(��"�~��+2g�U������C*1`�I����r�$�$/��Su�a���W8i�QPP�'78��oܫɄ���ܐX��p�%L�+>ލ�Q̉�+���'`�M١�`J�X�O�;@�>h)q/�2IZ9���w�~�$�����O|������J3$ē%�(a�'rͭvs���m�,"{���(\r�q��P�ɧ��r��'��!�e��^1C@ꕄ�M[���2�D�C �(cV� A�o?	�����O���h�4(�h�vI+mS�Nd���"�-�Uݨ�(B��¦Q�z<Ic�dV�����RGPS�F�Q�'��%%,�?��ϸ'�t�reŚ}&�T[?PG��(�{�-��'�d�a@��))q��HrIJ�|U�J�L�9!��}`Xg�����ޗB�� �!(�O����F�8��u3-��b7D�;'.��9�r�ۃ��wy�O\���#��=��EcЭ��g0N���� �%j�K  ���j�J$�>dY�"O��(v-S�El�餋�y� �#-`�&0��N�Z��Q�=ո��IBr͹�+�K� f��!"�[�":E^�6#���$�	E��p�/L�c��7�V�eXNp�T�ȡ1���v��,�v�E��:�ݼn]깘��~�?I0��P;�����v-���5�kܓ������Ԁ4�D��I~�#mՀ7�P����B����L v�� �e��FP@�?��>��;%�@�Q��(+",*�0C,��k���(��	�z� �����T�b�JB��I���|���RL��z��@�D����"O@%�f�ؘ������+Z�z��i�h#ع� ��Z)Z�B�34���ѯKz�ત�"��H�1���Ǌ���d��X~�ء�|�ȳ���'�<��g�̈l� p8�hڽ	]D�ΓzB¬��I������'�u�4o�~��C���$Dd���Y�����LYXu��_�gԢ�#��[�Juj����'.����$R�Arda!A��9R���S�팾d����c�K��ʕ�}�F*
ax��0=>.M ���`�<�!`3(9��)PE��H���H$a�ay��� �&��=E�ԧR�f��с��?qK��У?�y���7}-�U�Љ>h0����e�4�y�iX8?df��'Po�d��0��yr��?�.Đp�؏c�L �W���y���#q5�,"�+S2e�����+O&�y�[�VUȁ�cd^���piH#�y��K;�0S�	S�R�nk���y"���^<��#��M�(�H7J�<�y���8t4Hd�� 8���!厅��y�+[�9!\���MZ�PHՋ�y��U�Z�!�H�R-T��
�yBd�4
L��'ŌR�B��t"r��'���4���<��0���H���Z�'{u����Ri��i��W7O��{�'����V9����W�W�GS��k�'�ޔ��OրD���ЌΞ,G���'�2�qϚ�	A�M)��'G���e�I�mZq�#4���
�'P6�9�@Ӻ0��A�B�!y��	�'/4�*�/Q�h��v�	�p�C�	�q��u��i� o�ř��0l��B䉀.�h��d�S�\��	�m»?�B�I`%�	�6!�L����W"L�EnC��A��h� �8X"��W&�C�I1h.Tm�G�T�cب
daTU��B�I��|�b��PV���=x��C�	Z��t��#�!*C!��)��B�ɊuG���ԡ�;5Ǿ]P4N�kD�B�ɼ}�.����#�Y��!Q�P�*C��7'qzXcC�
�`1i3��5<]C�I v�,���(�-s�|�3��T��B�	�?�<-b�#D-ZI@��2�@�;/�B�I$`�ƕK��ؐ�6�I)^�O��B�I�l@"�Z��1G�*Q;�Κ�~h�B䉮�8	Z��˪u��ga�bp�C�	��R ��ً`(�����~�8B�I!���cG�;wȠ;vD�#.B�I��իC�W33C���uk=9�&B�I(Q�2���H}Dt]K�%O>C�B�I�-Ob�:�H��T`"��J�:dB��X �@�ƳD��9��	4;�C��5<HXXyDER�J���+G�x�C�ɹ^o��`$�zG�Eq�75�b�|a� 0;�����A�,ؗdx��#	:Y`���#\��Z|���ʚ�Ǧȅ��dK��H�f���LsP(��9��9��ic�#=E�$Dr�H�䏓q da¶�ƘC���c�Ogb)
�Jۂb��:��[�/��I�`�?/��M��'1��uP�Pk�	yve�D�Ω�O���̊� �1O�� �]05���(ԙ��cˠ|ar��57O����`�i���$\yz�f�Լ( ��b��N(Ub�	v���(��		='�e���O��$�U��7E�<�'O����P�4�h��޴;��͛�́s<���?�O>)�C�[�L�ba�>-� ���mD��u����ȟ�)8�o��xh�b��	'D�D�"O:ȣ6�Q*�� �+aHHСb"O"9�`�?2J\�Rn�-#�[�"OT����*L4���CR���h""O&�)����J�@)7kK �fÆ"O��wAU;�K�i�H�|��'�ў���h�ȕ�)�m�(*�,I����TH�'���+�O.dT�b��9eU���������.)�R�y�$Z)Vj�ؙ��1T�b��E{��T��c|�q�<��!A��N\\��ɏ�~�c��Ĉ%E��Ѷ�ϩ]�䭂L�V��\Z�'~L�Z6��"GA��T���
�D/[��`��)[�$�A�M�*O��(I�m��A
ç0�|���
2Qe�b�#�0(�:�C�Ǻn?�$E��&9P�O�>�f���[z�ya(�,Lt�9�BA����«��C�qO�>�@נ�I<l�Iϵ1�^����O�ف�#�)�&l\b���1#B���K��}}<��'TB�R4��U�8p���@�@���'�,���D�,�,uh�k��?x���
�'���n�\rCW�*�̘�	�'������G�v�x��ag̯5>��	�'���fg�[����ܸ3$�s	�'}�dw�߳@��IY�c�"(fbIp�'�^�y��Eִ
�A͡#��q�';|��@��5(�������L��u�
�'��)�T%�'eB�+%L�*��	�'��Iq���P�N�5�!_6f�;�'��H%O!�@�a��Pm��
�'8�Y��`0V� ��J8�Y
�'���"��iZx�����0���	�'�4e��C�{ɤ�`��O#nm 
�'�ab��4v��h���!p	�'%l�)����]#��jєBG� )	�'��i�����<\1{�' ��IcJO	B�����Ֆ'=��'d�P`)K�1��y�"C�����'��t���#kA����6Z0,!�'����H��(��d�+&<A��'!�{��p�>A+����a�'?\�ee��V���1���>�ht��'N�!��J��d��PJ%˘:e񀠣�'�fԓ"΋�%��Akg%ȓ`�ZU2�'I����X%%�RUáh��\�.%��'5��ӫ�4"�$����C�^�4�z�'��$�����A�,�Z�����'uj��T�T�J��S�C:P�P�'��p8g,����I���,^� ���'H�c�78���Q�=&〘��'��E�u/�2�ްp�kɪ.W�P��'��,�"*qY!b�*VF���'dtDIef�9�:	J1!��Y"�p:�'��1���1vZy#��M#r��',th5ku�(�6A
R�2�
�'$Zp�bf��:gt�x��S4IWJ���'�#�Y�vNnqh�E߅?X�	��'wj�y��_>�  �Q�0Q ������ ix���w�ƵA��ua�f�<A�mN�Xϴqp#�ܳ�l���M
e�<	f�+h�R�+Q�+C���  �^�<��e�1 ƴy����{w�!ä�<��*؁?64� #FX#o�e��c�{�<� 6}RļS��0[h�,`�5��"O��)q@ֆj� h����r�Z\��"O��h��F%B� ��2��2����"O��9�'�%Ȳg�������"O��yB��(7�$)���J�tku"O�	c�e�	����	U�[���0�"O�$6�؂^Sxa��&�.a�Z�HD"O,I�7��)�l!4㑞�\e��"O�XT�DM��]S�AіP��qjg"O�< ढ़*[xd�� /O*Y�"O�(�"�H,���B��}ӦU{6"O@9%H�10J�
`�d�����"O�Q����?.V�I"ub�	�TI�"O0�����"=ZU�B�S{~��R"O�x�6��|�|��ueS?)���s"O� j�Ç$<�<�!���>��w"O$��Gi�	yER�c%U=kZX���"Or)�7듗Wuj9��ۊdV0���"Ov|YD�Ǔo�֤Rp���&�~�JC"O^�a�^�TI"-j�l^�m�X��"O�� "�:�l��&�N�w����"O����"P蹨�k�{���x�"O�X���5(�pDh䊃u�TP�"O�㇬F�f�JŠ�ɘ~uX�@"O�X#��֡5*��Qo
6?Z��F"O>	 �вcK2	KРR�RWL��e"O���O��8�Y� �yB#"O��1 g̯n��l�u�K�"s��H�"O����/��;��L���W�Sf�XB"O|���m��|>)��o�1	[�ru"O��7�ʺQCo�#"V~	�"O>4���A�ƅ�aX+�D���"ObU(3��4�Vq�VE�a�I�"ODlX`Ɖ�&�r �Wi��OFu�"O����
7B�~ 11�;"#�b"O6 �&E�:Z�0���J�q<d�"O�M��	K�K� ɰ�Х!���"O�h&�����p��%�,�����"O�I3�>T� ��To֓i����"O��� ��=d{�B�H�0G�8  R"O�dђ��Pd��H�0L<1"On��͉*`�pK�m�,_̺|��"O��bBŻy@"���
'-�Li�"Ol���o�\�z��ڱ`�Zس"ON8Õr���ag��v�J�[�"OH���\�Z�� ��-r���"Odتe#�3eq*(����JU�ݲr"O�xj��L{���N��4N�Q�`"O�h�C�����UR�fPLT�x�"OBR�I��*л7�޽"|�{V"Ov��$�׽7����F��x�q�"OHu�+C�4վ�8 `�=>(��bd"O^i�D�z<�ʡ���\7�Ȉt"O�dA�Ӻ)�̉��Y� 
A��"O�T1���/�0��J\g"�9�"O�4)���*�đk>c ��*�"Obe�e��&&��,�b.*)Ѐ"O���Ǥ@,4�P�ă�e����D"O ¶��"#ְ auA=K��u�4"O��9b ������BR�#�"O�D�t�Ϋm�ZE�e��
���"O���ãe[JЈ�����3"O��-��#adKqj�(45d�ڷ"O���B	1���v��|@�@�"O� �p�ͦ5j�ZpD�[�u��"O�5��i5�$��ǥ
��m��"O���I�7e�ƌ�aӉO�y��"O�u�B(�
~���z#`�~p�Ja"OZ���L\,
�����V>E{�"Oָ����1�"WJ0>�8�AUE�<�q�M�&�z��!|V	1���<��F��#֕��B�N[�|�db�O�<��ĖrjDi� FF�3�NM�<Q6�ɗ�������k��#�*H�<Yw�¿$�$Q�
0>8[��VE�<Id�W�5D�;!J�t�)k�A�<���H�Iqŉ� �������<GG
}߾<:;C#	HR��O�<�
�QOz�iT��D�|=�$�Gp�<y��B/@Ɗ�Sr��"��=��$i�<�BMU�{j�e"a��4+��*0�Nc�<�3�G8Y�1�B�Sk���b�<�CmT�2ޝ�p`چF���Y��IC�<a��-^�⁠����4	��fOY�<���5 <n�C��AL�9 �)��y�Č�]� �f�#s�2�`�/���yb�8g�j�c��[s=2���!Ո�y���D��԰���l�¨3��y2�\�&c(y�i�`���D�:�yh޳zaơ�%BƁf����)�&�y"hE9-�d�dE�`���sBΤ�y��P&"a��KH)F<��1c��y�M��a� %%Ů{��P`��y�㖦\00��m�>i
!a���y�O�Lش3E�_�Z�p�b	�yB#��YT.\���9:'E+�y��ÍS�~	����w��1�+�
�y"�S�xk�|0!�7ov�4�2��y"�v��=�o\=b-`�;�Ƙ��y��y4�t�T��A��X��y�N�dR8Xu�Qx���{g���y��-��
�G�m�v�r�K��y���y���A�r*\��f���yNT�(�Dq���9��h�/K��yb��9[��1D
�.A�)ڵ�� �ymW�F�'֊�P��yR�o �48���gN���蒲�yR"���������4Pɠj=�y��7"M*��M�,^�N�rp���y���f�Z�a�d��O����y��+��1�?{��9�AB?�y�BL}0ܨ�
t.bI����y�?���Jq��"d�00�L��y�@�/<�
���oF�T&�4�׮Ќ�y�I�!@���GO5�� G���yR��:��=�4���mr��K	�y�N�1:�Q	�K*9|�dDH��y�N�@}���w
%��=!�`I�y�I�
vj%��}���ɰд�y��l�����O�5L�L z�E�y�J
�@%�u��Bg��mߚ�y�-��T$�(f�A��HL��ybbX	0�İ L�T�(]��б�ybI�:�`��L���!��y��˷W�pɠV���@������y��Y;���EA,e�9�a���y�虅�z(�fA��\N��[ ���y��p�FY1�F��Zx�P��V��y
� �]Ѐ�El4hطiG.d�Be�7"O�UYr�Cy��	"G,U�{B"O�!u�X�`���F�;EI2l1T"O����}cBXab�
�[G�Xց5D�daA�99�p��KE|cj��5D��	Fg�5��[���:�6��4D�@Ѡ�.������L�JФPP�%D� ��'��rgv�Do�-	�搓�6D�$� . �a�B�3��*`�
�H�.D�����(@B:�U�N ���#�i?D���H[43�D�QaA�W�ԥx��/D��@��t$����e�0�
i�S�+D��"��f;`��c��W�����,D�@���@��Q�Ö�+��(bUF/D���/�&8� ��鑲I�z<RP'(D�pC 5vpȂ�O�[�b�+�D'D���⣃�U��M��M(5�D�Xp�(D� �ga����BcϜ.g�0��'D��h3/�L�l���I<P)�My��2D���H_�|��4iM�n��pL1D���B/�  ��58�É:[7�,z�f-D� ��@F�R�y@	}�pDc�n'D�P�!m��N�Q��^�W� ,p.'D�T��#�40d�Q!�B[����1D����   ��   �  �  �"  C-  17  B  MN  �Y  �d  m  �w  E�  �  ^�  8�  }�  ë  �  L�  ��  
�  M�  ��  ��  �  Z�  ��  ��  $�  b�  � �	 * k  �# * �0 7 ]= F zR Z �` m �u �| :� {� F�  `� u�	����Zv	B�'lj\�0bOz+��D��g�2T����	#Ĵ�v����?YV����y�抋<+��{e��%d5�y#@�iTR�Y�	&j�i��K�h�e G;3k������!@�)]P��up@k�'MC��Hf�H]�ڀ�J ���7h�z�\9Дe� 2�"u�;>����!��b�U�D�[r�+/��њ,�<� pa�L�g-D���V>�1x��޽h�&�l�(����I�������A:�%��e� nX։چOؘ�����4�(` q�®�M���?��' ������?Q�L|�!Vm����E��1��,����?q��?��?)�x�.<�E.ɳ�� ��'�P4  �vi֫E $(Մ�R�x0#���yD�<Q��(O�5� G�.c�\��ǺT��1�eZ�n"��y��I(F��q+�kT�#g�$A:&�%����=�A�F-/��'`�'���'b�'�Sżóiϙl&\Y��	sb��t���؉�4��V�O�7-�O�qo��W�<�Hߴz.4<��$�o�L����IXN���E]�:�V)	�R�(��4�*ș�p)�H��!ʱEY�'�M[�Oɐ͠��Š'|ڤz�C��/����̉
�P9:�g)`8����fț�Myӎ�	�?=���f�)p���CAB��Q^G��7� �w��1�h�6,����0y��K��O��l� �M��i4	A��=:�q��I��<؁GS�@qړ`ۊp�,7Mݦ���4u�퉣F8'�*H�Q��d�d�t!�+ע,!o�a/�pjǀ+i��z`���1��i6M�Ŧm���x��{1bR-�\���A�#��Ir�2lB|�@!Xg^�:�4N�����s<1���zF������'.���c���kcZGq����'��O����O�������O2Z`���?��4�稙�|l��@���D�O��$�O x�w��7+�u�5�������9l�N�=I.!3��];Ab����"G�4Y0]4��oZ1}��RiM������/	D�|�A4��f�$`gƤ<)W�0�
G�YդQ�@B<c������OT�$�On�O,���O��?��h�;O6��0LY-N]4�{r�Y��?a�f<j(�P�L������|�%�'��c#���	���� Cߔkxx����$� lJ�Yl������wk���kG�؎Mz�̤^	�`���?1��U?D���EB��F�ە*�����̭(��`����H�0?	C/��&QH�Һ �>9�g&��T�I~"-�>Y[N9c�.��
Yd��g_~��]��?i��i)j#}*�O�6��PMľa��Q%�܎H<�PK>q��?)���d0�S�g�7*��@�#�c������ʟ���4sK�&�'�7�g>Q���3#�<��""�I/U�����ayb%�f����'���'G�=uͰP���p�̀�(� ���ʕ�G�M�A(����} gaҎ���qO^A��5| Q��Q�΍k��?	�b��Rcz�\A��E~1��h��<ٱ���%:�`�S�ӇB�ԩ��"�"�MC"V� z���O��i9&�H�"�O�v�H�蒆� Y�j��Af�Y�'wax2��,s@�q���`50�T<�?�����Dr��O���0�]�H��88b���@N�'�:9��Bf���O ���O�ʓ���a>u�c��z���R��� 0���	����	�?O}��mZ<@p����:v��Iie�:!���x � ^@���tW$urA0�@��f�@f�h��ֈFzH\�������%%ڜ{L��w�'-�6�\m�'��IZ~�'��z��}@�P�#�2ٻ���,�?�ϓ��'K���ǔi�"q31����Av�f=O�7͍ͦ��O���c|���$�O�1h�c��*��O��s��[cc��?���ԝx��?��yP.qK�I=0=2��i�҄�2oƞ�v@S�ق��&��ax���(6�\p�'���!6�=&h��I)@|���r�C(%JT���D�.#��䝥`�r�'��6m�O�KСגe�0�q���ےd0�<	�Ɣ����u�4٘'ܼ1�a��.N�TM��" �L�I>�C�i
ў��M��#'2�v)3#,�7`<-�Ћy!���'&�7�ƭO*>HlZo�ƴ�'g���?���+C�cJ�P�2`ԋP�R���^����I�l�)��I��T�6E�S-GQ+��A�����rM#�V5�x5@����U9��MB
UK&�6����5)S&^��U��21d|�r�͊-�2`�ӹRp0#��F�:�@��G��t~R
ˍ�?��iQp��c>�kG��)z|*��M
 j�y��4���O�OX��OD�v�<�G�0&�xqU)V���X�A�	��?	�4�?���i7�!+g��re����Ŝ����޴�?)��?��dϋu7�MY��?����?9�w`:����ҏ;$Δ�Be�!��� >���sFȱ"����&���Ò�^CҨ�ゕSjP'��0D��;��b>c���EN�.�~����GN�H�)��)�*O�xr��'1��'^�É4^��@&��T!�MU��4	!�d˚[ذ ���;���T, ��j���X������'�l���_4��$NW�+[Nh�Co����7M�O��d�O��Şz`bm鑦.<���vR U���9r/̞[�kF��|�dI�Wg�8��<qYX����!#=�ECƉZ/ڱB�A*,�1� .G(`L�+n��0Gx��ڟfI���Vؼu���5G���0�b���?�����'�>��4�_��D1��2].�0Sb |O4c��:�+3��8���H�*P1��?����Q��iyi�5[��?)kGn���zݨd��( ���
 �O���?q����D<m7�YjR�,E����Ċ9�� *L��A�y�P(���ˣ���S�'O Ez�EŨC0�}K�a�ns�Af!�aj���ʁlܦ٠��\6McV����O6̢��'1�7��my�*R1T2�8��d� e���L�����<Y��\�$�)�
��a�`��#�"��eY��?�.O��=�'0��ff���)q���!m�i����,`N�6��O�-n�	k�p��4�?�/Ob��<�׎[��pp%	�[�l��؜�?���H�۶O�x\��H�H�_i
����t�Ж@du*�H�T�@�Ã�3��I2�z񉇁C��{�"5|�������r��%D�;%�@�@�6I[�-Y4%4�'��m���0��&B"�'����K8w���!�C8hh�h5�&��>�Of���V�& Vؙ�lԴh��I�2�Iş Y�4z���|��W:c�\q)����H��`��Gz7��O(˓R���"�'�?���?�-O��0�K�V�����YQ�⩲�jSip`f�Ġ��X�Β*!�ʧ��=�@�"C伸���(����D=8�j�qC��(��\cAL��'j
��|�b뎣�p���x!�F|B�rB�L�w� 
شM=�ɒCe�D�v�g�~8�:a�J�|�Q0�L:	mL��?����~zu%�HH�\���Z��C
��x��'�M�v�i�ɧ��Op�	L��e`�ϓs8 ���[�5��P�-����d�O����<*�p瓈[��X�!oK )I@�n�(S$��֍ϼ!�h���؇�$�I	˓[1&})R����H;�.D�h�Q��6*�*܃"�/ȘMs'�ք/0`!�d�'&���ꐋL���iу��cq�;��'�?I�i��"=����7{�󣯘������s�剞�HO��6�I3)f�x����9D H���c�@n��O
Yo��M�*OZ��6'���)�	�<����U�)� QPҙp���R��W�t�	�����2ث�F��G�0��(�7Oi��B�7A����(�6��dK� �0<� ���N�L����ּi��K2�i���ѯ	�ߊ�� ǢD9��[�}N�h�	՟��'���X��[K}��Rw���Co��O>���0=�£�	��(2 .j�d��Gy��h0�J�<=�0@����c��]-5� ��Ey� �z��'	[>e)�Q��|��j�bt�HC5���Vߊt�&���0|����̼]�re���i��.�8�t���F��g1l]K�.�
Yc�'���eDP0"Ԇ,��b�h�X�Eאi׺d��?�KCܺ9�"�*l
|�T�d�8?�e ��`�I}�O��g���[��	��� b���^.�<�[��\�䴚�Ĝ�hO��O�':���s��1E�hA�J�� �S�'v��'��/(	"�c�'L��'��<��-#͍)P�l��ʔ"t�S�Ӻ$� o��X�+���Ptc>c��+�hN�j�~S�)�&�~]�ۥr�$\��4R������5F��H�|B'"�5|�>�Γ&R��[�ΧV��*��M�S���p~"���?���hO��Zf+��q�pqҮ��c9胕�2D��2�P�(v��Q�]�x���.�O��Hd�����'�剻+��AY�B �.�H�"K���9{��]v\t�Iȟ8����tQ^wQ��'�򬟩A:�!�@f��p���k�F3���(�ܩ?D0x D/`��L	��'��M !����b�*��q
\�2�hH�,b�| &[6E��1SdF�C�@@E}r��&$H��M�3s^��/�%:0a���0��fm'ғ��D-?YSL�R<5�1��L�G�\ܟ ��]̓��pڲ�=Aྀ��l��kM�p�	��M��'��v�{ӄ�'F_�]A��i���'�l�1�)�"u$�0.�<��5�'��	�"�'S��Ͱ5�X�����tDxf9�^!+$��/U5�֮H�U,|��T��B�n����.1}�5HD�|I�5A�ձx�DI�d���+�M�� 2�t��!9�|I��̖4��(#�S��� R��Y�v�*4����9�!�$ۏs������9{p�a�Uh�O�=ͧK&�D�Xˊ�a0�݆
�������X��=J��?����Ɂ�ǌ�$�%Q���s(��&>��2E�!�����O�9��sh)S,G��MӰg\x���?�іZ'��s%N=ټ�)�(?��Ҕ-���P��	���OF��������I]�I� �cg%�87��(�F��JC���uq ���O�}*�'Id��&�3&��2F�0)�N�J	�'n>9r2��1ub��h `
�XN�Yڍ���Ob1Ez�d^s�T���4x@#I�^�2�'a��':����u�r�'d��'���s!���́AH�(� �ߐI��Y$Vզ��aI�2h�Lj1+<�3�	�=�\�h�JΤ�i��F/b���	�MCC��	!�~x�r��ņ��xQ!��<��(��*(qy7��?���A�J �� �'x��?���D��NV�%/�8e�^T�@��A]B��=j���A�ƅ:I\�����r#��O��$ZE���$�'��	�Y����E�ʌI��#�BQ�+�HH4�z���I���������̟��I�|��l�45�Lɺ�O��3��!ʆ�R"�$�*��P�x�^�J��i��ȇ�Ia�h�  ����-�p�t(�3�9x�iu�&�����ƦYD�!>�>�I��5�<
0%�� T@$�E�+�@�C�����I�'��,)W�	��t� �#D���`)2|O�b�t��'C+*�d���*0�Űq�0��S����	gy-)d����?�2�
,|���p2��G��ݹ3�J�?A�Ql~�����?!�O�<Y6 �xֲ�0Юf�hQ���
��<J�ɂ`<\�ɴgX�+�ax2\�zy耛�d5��7-&9r"`($���P�@��T�)u��懌p����b�	=?[����O��-i�%,�e,͏)���%����ɗ��yrA����<#WF�Q���D{�O�@�$_f��s�ȟ@Y�i�f��.8�Q��[wDP˟��Iџ�O�VP���'�Ұ� "|=�Lh�[y@����'���,��A�t�$(}�oD�Z�'���چ!��m@բ�B��薄L�X�I�#���τ�|����۴D�eA�/>A^��O�D�'��|e̝8�H�2)nD��OĔ;�'`"��<��L7l �� �:as��@�|�<Q4	�6}�T�m0ey8e�L�'4R� �m&��0MH,��cԀ)9?f�2��?���?)`$��`0��r���?a���?i�w�`�I��_!c�kD소C��$#G�V<7��"G�(a1���t�1�1O�p�V�׈;�p���6q��d��LԢ	mڷ =4�;6�0�c>a�e��;B �+2<f�����Nl�XS����Fr��$ ?��l�֟�IM�'30�����xa6�J��V;+O��Y�"O�h�6Q-|^� x�����6QQW�'uJ3��|j����Y�۰�"��^!.E",�!,$����_��$�O��D�O����O���r>e��NW�:������2Y��i��
�n��ٰ+C��>��޴^p�����gpL+S̛5���@�[�i3�	����<1ACԦ���H+8�؈�UD#2���x�Ù�Wgr�el[�L;v�`�I�؟ ��M�'1��8v���&5��ԭ]3�9��g)|ODc�x��*	�7X��䑺2�`J�&�NŦ}�	Ky"�@ c(�'�?s/� e� ����A�����/:�?���L˗���	�|:�#�Y�悚�J��9���f���&5�͹���+����ɥv��� p�&�C�
���J�OL%w��8��O�`���ւ�����Cs瞔'ڼ�s%�2?���k�'֔��ւ	����E��7�^�:
�'%��b"�-;��<�$��0�����3�҇&z̹9����c֒\��Ѡ�?)/O����J���ЗO䘝s��'��tRM������B�+��}# �'�b/��)DD5��֬0���͑� ��S|��n��|P�����W��8�&D���D_>`�2I@C5����4
��KL=����uZ�8��E����v�8��I�
�do�)�'p���k!�P�jD�	��� �^u$,���̍�"�^���i�J3]g��E{��'H#=�m�2�D����%39����:fۛ��'���'��dc���n��'r�'���<��X�@��1m&�����7�VQX0I�.
JF��J�K����J,]N��w|!���'|�C�D2�D��P�H}�U�"FJ0�@���ʴH��iйb|��=��x��.t/z� %]�+Q�)�9��]�+T���DЙha�h� ��DQB��d�!��<2�%j�ԇ0<F@#R吲8����HO�'���-U�Jl!w��.C�-RT)��m�iQ�M�E
����OJ���O\���O���h>)(��H�i��H2�*e|�" GC8[j����$��F�rR�i�P��=�X�C뀇P/T=�MU��>�xf�L#3��	$fY��M��֚(���7�Z�'� Pz��m��RQ�Yj�	�AL��?A��hO0"<aeE��s/�����F����E�P��<�<����OsvȨ��HUTPm`�bEK򉡪M����Ą�YwQmğ��I/=�q��*z~$ڰ��g0e�	ӟP�RA���8�I�|��-y$��EA�\g�	�J�}��2�8��K�0U�D���BA�q�7�̴z�j-�'7"YC�iǝc&��%a��H��9!ÓL?��	$����8[��JJqB�钟Ӟ�ȓc7$Ł��H �0�Ӭבv�����I%�?yvH�c%9i�Z�D�U�ɬ3�R|��4�?����
�Y���\n�񙲂yU`��jX�W�r���O
��c�-�l1zT�ʇ\��Q���|ΟLS ��s��&lЬ����(�t��>z��Q2dQPc(I��s�Б���@�P��e��9�F�]�n��0"�������km¯o�v�m蟸G�d/X1����GʪZ �bJ���?�K>Q��$�I��<�tc@����YR�A�`Aџ<ܴG��|�mN�L�{��`�(�:�`�l��$���'�'tG�	���'�2�'����-t�H���G��Y����lbɔe&`\p�&7d��A��n�g̓@��J�Na��I��x�:��M�c�Rq�i(��J�8BT�7�W��M�O��ų���y� �}��@إS�N<�o�3��L=���6���D�K���k�!X�2$�f�]7'�!�.W\��(�fF�l�\5+�#T�=��$�HO�	4���(z?����:Ljb���&AE{J�Z6DȽ'(��$�O����O�ݯ;�?����?!e�Q�@JR�� tW�I����kʑ����4h�kT#�/|�����_AZ�*�C@��D���X0^���d�(;j`���-�D�B։��s��6mC8|�	�w�>?A�-J�*$ H���v�t�c��>B�i�IğxSO<����?QN>ٜO�V�PK
�-CB�9 �y��9N>	���U:��X���x�u�̤dΈ��I��M3�l���y��'���ƺi�r�'ڂ�Y����j�)���&��Kڟd��8�4��$�	�vb�&ʨp| �YE�i� �X�$4`���DJ��b�f����dٲwM���@�+���&�_�8nΝ����(L�����B!N�TDI��Pr�v��U"}���'���2���O*�m����DZd�ѷ�
�\[��J񈐓LA�'B�R�'M�DۓEb�!G�p2�$
Ȗ5�!�dx��F	͘]��h�Ä�X�0��%����	��M�Ċ!�?��?����`�N��?�k�f@|���*!�ʁH�	H�?a��}�|[!o�s�� yM�V&�6]>!�O�B�i�O�l�Ѝ�Z�������bd����'ʓ ͘-��_�H���Q#�?V Xy
���e�.j�i��N�K�n�^H�	џD�3O��7���@mF|I2�m��y��
p^Q*G�O��a!팙��O�=F��蝠w���ğ�/ ��e��?q��?Y�����A�(̡�?A���?���yG�y� �X&a�hB�nB)��*\
et�7-�	w!�	�S>)�g̓[8ք��I�9�H���R8N���� 7��� �J4$L��0���aP���|J�PeV,ϻ��Ʌ+И|ܥ��C�	X��	S~�m�?Q��hO��#ӣ$Q��x��0/�)y��8D����Lza",kB�O }9�	�i�<qG�i>���uyR#W&�y0&,Z5#m�Tg~����Q��a���'�2�'��4�'T�<�N`H/��xyj�F]"�`܀�M�VL�@N�/@�m���<�W�N�,l��Ti�{D`}���l�#A�F݆iy���'pJ��S�X<$B,`�W˔L%`��'O�X�� Co��uF��|���B��?a���hO#<iC���*�(4������ ��J�g�<q��c>t��	�>
��x��i�I��M3������'?��¨MYxIi@~�F��w�O���?���?aӣ[�j=����!6�I� :6l��Q�JЩ8�"�Q���L[��a ���gꉩef��),�҇`�P��L`�žSyf�kAm�f������O���8?�2�/53r9�c+Ťt��;��If�Ie�dP7(ȕ!����狦Z��U��0�O���ɗ!Ҳ���nJ%�N|���زd5���<�� ���?��Of��M�V�H�dV?_�0�e-��Zs2�'Y�IR&�J�.��'_M˜Hi��I���v�J��{���ۀkZ�6�����PT�M���g��c���|��E�Pc��st.N�|��؂T OY~��\�?!���h����:\���L�	NO�h��b�U�C�$Yp�%ꅔ����P1>�n�?9��S#"| �0�� ������	�J˓��L�R��O�d�O�v�Ţ��M�����A�@� DR��j�q�g�ՐO�iHW�M���Is>c��#�E�]����7����P12cX$2v�ٖC�JGjȃ�(�8Xc>c� ��c%7 �a.�f�-Z!��OB��4��	џTD{2�!2��{���\eQE�ݟP(!��l3�򤦑�`l:�̰u�I%�HO��ay+	�G&8 8g����b	�3b7�,X��'��'�bR���?�q������E�$09�$�ԌE���SFD�*�s�$�#G�]��	�&Ux���-�4���ee�/%BHM���B#>�\�ܤoV�m3a�'���K�5n!�!�k�1��@����?q��hO�"<ɦ�I�F�,2C˂�@�b<
S��C�<�䏍6LqT��'�(&��2@E@�	����<Q��(��OM�P#��ṟ���K8yL$�������O����O��!�KD�T<��J��y7l��5f�J
�u�gV����hc,I��|��Q,ڬ���cH�E(~�Qw-G>7�9b��դq�eJGmP�HIĤz��'� ����?��Od�Ӱ֚a�����b0���C�|b�'#����L��!F�Hj�a���1����%1���K�.��P����;�?)O��!�<�O��ٟ�BfZ`�n��1`%Z����)��� �	1ln��V���}�Q`�RЦ��
0��r�8b^�F��[G(���ܧd䪥�FH\�"��]�ш��(�B�3�n�h�ʈR�Q�Z�@B���	!D�O���6�'�y
� x,���Z�"�2��%Jq�	`�"O� з���4ɤ+Ⱥ�#%�	��h����\�9�r9��)= ".�iMb�.e��(�<1�㑺����$T6������t1�A�ڼ`_F�C$�ĆF���ZTFW�-}Zi���9�3�	3(�t�(g�[��i��G;)����S��H#��voٗx���5�3�	�]ÈqP��A�5�ͦ2��� ��i̢�*o6�	�?!���"����H�!�H1�K�#���'�i�V%���U�'p�9�)O�iGzʟ�ʓDȦ�SCI�<�XS�5������2���F@��p=��U0��Q�U�V�c����J��4K.޾j���5'P����I#L��4����{>�d�0\`=;��?!�4x���s2T��Ǔ�� ��n	�F>�E	!/
�b��5����ܴj2��dGx��ǍH7�P�*��lX[�E��y����P��D�#�\9����\��I|yU*��7˯h���� ����@�������[W�ў�Γ���E��k۠ ��mA�� �45#�%���0<���K�'wF ���6�tI@ĭL�wb���T���I���>�|�p �݈_	�eAq8+Y�ć�0�����5����U�3
�H��I��?a�F�2ϖ����K77;�%TgJp��2DhV�4�.�F�T���*R���6A�Z��	,Q���Ċ������T�D��$yrb��(�`�s��K�[1�0���BlѠ���J�!2�����N���ӫl2��� �;s�e+���#�
�t咵�Ʌ�Mk��S�|�����:��K8r��Pa�<�"K]�]il0�i�z��=rq�	^�'���}�bл���#S �)�f�ذ	Ŗ�M�`�N���d��'��g�'*�r�í6�HAzgJ�j���Ïy�� �0=�b놎WҴ۴艻�J��)z�-ǒ���ɜJ��yK�GӭR �=yr�=�p�%� Yr��O`c>c�DhjT� s
 Q�ؒ6pHA�2D�Y��Y�b����Z�"�J¥<qB�)§Pb���!$/oi�1��@��u� � �(�~?��CU�@��3�F9F���v�R�4,D��W+E�?iͻ{rX�ChAi)t��iġ> �����@�I͟��ɿ-�L�RȄZ	�Qa�i���O*�`�o$��A�.�W��qh�����{rM�K�1i�n1`2�9B®��9EBY? lPe�ǣ�]u�<�b�!�d]̬�	��h�|*A])TOv|Iр�}h�0�Q�_Ny��'��(���B T�1�d��"A�@9I>���4����'�.XDCI�0��xh�E$Nql(H+O�u;Q��O�8JV��O�˧`��pj�'�?Yg��:x���Ĉ�1z[*@���I>�?!� ~�t��ԣF�-3^6-	d�S}̧=�T� s���a�.�� ��
]Q����P�c�V�;��)��i%�R�ZM�6���d�?9��$K��y�61�Q��<�yR�K2�?���������tr3��8�xC��[�\�0E��:D��ᡠ�6xL��'�e��)8�I��،�4�����=b
����<nܨ!�vr>�$�O����&Q����)�O��d�O����O����'!aS�٫�kP	\v�w��2�M'�6�u�N	>TDx���?#<�2�V�4�kp�C#+Q
,��l^�����U>G(�= �Dɕ`����ʟ��RC.Ǐ���M��䨰e���Iɢ�V2t>�SR�I៬F{�:OZ��5��/��3DK�[n鲣O
�e�j-Ѥ�;�0
r�O`�Gz�O��X�t�e��[�Vy5`��<�2��v-�4e�m§�T՟p��� ���?�	ß�Χ
y��j�
��)�3I�#t�Q�*ŕo�&4���Ҫ	��d�W8�<:u�̎c���a�/˔G�@̫�fC�=��hS�j� 6�p�p�4JU��@�W���Gx��ӷ�?Q�$�" �l;C�Л9�\H1�V��?Q���9��Ԭ���ތ%���B[�wl��IM�'�<�J6k1>���C`����3+O]mZX�'�Bհ���O�᫅*�p hkGCӜ|FT����%F܎�����I���+�	�2+�X�;7<!*�ͬE�T#c��[�YF|�C��p��<�֧�X&�����֝�WlԩP�ʙ*_��@���e%,#>��j�ğ��	ķLiYT���w0@����nNH�'Ta~�蜂l3l�h�J�Q�N�Ȱ��>�!Z��&�߄Y	.4Xeǔ�4MZ9s���<I����<a�����	l.�M�1,�&��5��
��n�j��+����k�
)�ڤ@��\Zr��9�&}��G����֤I����U0O��Jg��#���
���a`d�R�_l�O4���I�*�	�V�qwD��'�:`����?��O�O��)� $ˆ� ���C��M�6\3T"O\��nN�[� ē��4�d�C�ɮ�ȟ��Z��L�H�\�s��X'h鹣B�On�H-�H��I2�d,"ƀ���f�sׄؑ]��l��J�Rx�r�K&@mV��Ԯ%r���/'>(qub�.0����L�^(ñ�
mN��b����J��"�?m��}R�W�Z�Ľ���;'Gt�y䡓?��$ߏwkr�'�ў�Γ)Viy Q5<�%3FM<�.��6Q��B�ק!׶���I��`m���� �HO���O��
Pb���ٸ 6�JV��A!��@�
ޔ�0?�������8A���E�6�bF�
�(<�N ���	��6Q��B�I�Gf�P�'³9��Ю2�+�&P,mW����&�5<�Usc����Ole���'���"ʼC^,�ɂb�T{��P�'Jў`E|�!Ԏ-x����T((TI@�S��y"���#��x�aҚS������4�������qy�ڳ��7��Op��n>�iR�t��Y��FЂ3*���C�O^�1���O���Odx`oI�tɬA���]F�*��|BV�Ţ=K�0c�@�9iZ	0�&�E�'�4y���v���N0�M� &�!.�j����	=X�B��t+�!�Paڇ/o�pp��͚�y���7 ���u�i>��(�h�tZ�ǖnt���<D����.јJl
qQ��UR6�[D?�Ob��'@���	պePL�QF`A�j��$�O��Ī<1����	-꣧G\\��
\+M�蹂��\r?����O�YD����`=���b%E #vYA��B���'���x�%Q�ӱ`��j�ύ	F�`K�T4�Z�4�?�� �(�y���?	������Ă�5�hع����P੘1!��P�pa�3�i"� �<]52j�O�ݨ�؟�^w�܅��yG%CV�x#R�[.>����ٍG �������"���<	\w�"�'����'5�$Q!1娘��˔Pc��Y�#��c6���'���[9B3O���1ԟ�^w ��̓*���H�����K&ǚ/�~����3����I����2m����O�������*G�=�u��3(I I�G��\'�p�I�[�f���O�؋e�O�!�ɲ,J��sӬp�r��R,D �ʒ��*	�Ɉ4ks��m��?��ϟ���8��(����D�O���Dn `Yp喛l�0ɸ�EӰH�P���Nv�����O��$�ߺ����yc����4Y�`�q�`ԳD6�V�VEX�)��G��8O��:�-c�6�l����!��u��ON�t�����`�ޖy޶�6
@2h��6��C$�	�{�BQmھ�M{�'�?-���X��?1�h�a"Ԡ���Ǯ![��4K˙DU���D�?XT�p��'�M�r�OX�韆��⋆�Oמղ�a�0@��&�\�<�!��<A�Ԉݨ,@�ta ٦A���t��ݟ�����	��P��ʟ�"�,��+���0�NM7P�
�L�M����?���?���?����?����?i�4f�@yɃ�(q�,�K����<tV7��Ob�$�Ox�d�O�$�O��$�O��(YV���!R.q��2���� b6�o�ǟT��������,�'���n?��*ϨU�H]�5lݛ9P�0�4dSu}B�'���'�џP�E�Ni�5�5M�t�ՌB'�M[�����Oh�$�O��Oj���B��0:�!�z�؃@�Rq �n�ߟ����̕��4[>q�O����FK��8�t$�MV�X˥"O4<��o�$��rD�sP±p "O蠉���%0�� 4&���"O��
u�H��DX`���)dx�5"O�I؄�F�N�)��(4�zQsc"OD�ْ�D�}KJ�h��_8X��`h���֟����h�����IĄ�-�d�����[VR��6(Đ�M���?���?a���?���?���?)��
#}�����_�HS��xFM�4J���'(b�'���'�B�'���'�\��B%�rU���˟��I0�i�"�'���'oB�'��'2��'�]�e)@�����&��|� C
u�����O0���O|���Ob��O>�d�O �dC	RB�`$)��nz~�cJ���]��͟��Iӟ���4�	����ß�(�-��g��-�DǱaS�� [I��7M�O���Oz���O^�$�O����O��3H
�Jq�������7��Tl��4�I��@��ڟL��ğ�����	%V��X����aό<��ǒ��0��4�?���?����?���?���?��y��m���.+T����E)f�	p�i���'���'��'FR�'��'��=RW���zZ��3�C��O(`��y�<���O~���O
�d�O��D�O,��OH���K�hb� ��ץT�Ɯ�� �E�	����ٟ��	ß��I������, p�� kzAyP)�=��w��M#���?��?y���?Q��?)��?�@��&-�D��'U=q���7��՛���d��\y��0Z3NtJ�eKt�P��nLqD�loڅN��b����I�S��Mc�w�j�KhL�Z/r%�dH4Y���i��'��:O��S�c̽X�簟��qΞ�A���U$��s�@�Oک��G\BL�D�(��|Z�'~>y��T���e�k�.�a���$4���ѦaDm6��k�? t�ⶃ�.����0�A�Wш�#�':�'��˓�?��4�y�_���W�Q���Q&	�Z��"�<��/��@��|��J�V~�OԬ�Q6�U�-��$K |�JH@�ăƈ�Fa��ISy��'��>�	��䀒HA%:�Tu!T�Y���Ȧ�DO6?q��i|��|�O|�Вū\��<bЫ��X��|:�4O��n�P���(Kt�������*'�*3�d0!s�� ��$�B&҅(W-�<ʄ�IƟ̖'�1��H�1�!f"@h���?��Z!Q���ٴw����<�'���d�[�.K)>���(�o/��x�\���	�)ϓ�H�
�R�kًU�N͐4��+ҶE�"i������ �B��� u��r�5"�N��'r�K�bu�-{��٩�x�K�M��H������:D�tZçD;`�L�hш;V�����&�	�V���ڒ�F%1v\�k6)��˕n��#uV�#FǶO�`�H�&���f4:��^�[�L<[���:tZ���D�5w6�Lʬ{��y	  ��9����3�Q�oМ�����I�B� ��8r 	U#\e���pe��"e�HbSσ8=������1+I֮�z�0���پ�?��4!�	Ke	�z�Ah�����������T���S�ō>���'Ab����^�֘1,� �&�>H4q
�*5���=�սi�,H�'��6m�H}��O`���7_`����nX{i<#�ĔF���ZFA��c��"���4h^t��D�]�o �[w�,(Β��e��z��X�����
�#G���G �9�tC��:1|����U�x����e
U�tl�[cG-gB�?W�x�wAս?b�a�Q-j���\���m�a��9с��4+�D�n=r�Jmr���#,��rrDE�X�N���)�!I�����"1s<$)l7f��2��?����퍋;f���r�_�c��h���QZ�,Pa��@N���i�R�'�O�:˓+��B7G	�B��C�������	#v2�#<ͧ�?y�w1�:am���Q�
nL�)���&�aIıiA��'���Oq>Oj�O�|>�����M��{� G�dVR�b>)��ӟ�둬u��m���,zn��'�R�M���?��M��֓x�O_r�'Ym!���Vcb��`���W~�3�\����ݟ$	� :?	��?)���?I�
þ.����MN�+k��+��8�?���i�$���x�Ov��'D�	�|�R$���-����o�$�t��I�xEh:?���?��?i)���vbD�6�(вh�<1_�H��+��~7�	%���	�$�IeyR�'��G_!_�X��O��B��r�,PE��Ȋyr�'ab�'��I�i`����͌y�2|! ��C��K�tyB�'�b�'��Iݟ8��:Tn �*p��ѮY2�Թ��W!xi^��?���?q)OP�qPI@KⓚI.����(��n7n�� ��3@����I�� ��{y��'�bm ǸO�I��W������2?$����?�����^�R���'>��	Լ����-n�~t��Ռ	򜳀��ʟؖ'2b�'3�tڊ�	eލ��I):���s䊖E���kp*�O�ʓ|�Fq��i>��t��:����b�`�8v��,�(;��'7rON�1��)��g��6+�;և�*^J@aL��FHR�Ÿk�n6M�O���OR������O���#Z���؆�%S��S��&f�H�D����$�O*��|
N~��k���I��(H�d9f,�N�ƜrǺi���'���[�d�'nb�'b�'��iT*�!3@�c�ϙn�H�`�'��'Ya� ����O����'�B�$`]x�c��[�ے�#f.׬&�R�'`x)X1Bi���$�O��$�Of(�O��D	:�l(���u*�U�&ć,g���i��IП<�I�H��Ɵ �O|4�y�.Ynd~�����)5��Z���_�7��O����O���r��P���IS�06���;@� `��Ö)m�d�I��T�	���%?�E��M+c/F(=!�+C�z�q�&��?���?9��?Q������O\|�D<�F8��啒Q�f��'n��U��OZ��Ξo���D�O����O�e���̦���ӟ��MOi�Y��@�j!���W�������џ��	SyR�'�>�H�OJR0O 8Jr��?vN6�Vc$j�2��@�'�"�'4R�'�����yӞ���O:�����w��5Q���-h�$IIS��O��<��ӦX�WX����Th'm<�]�%�*OdmuL����'s�?X26M�Oj�d�O,�I��v�dX!s}�c`*N<����1�#u����?���5�?)����4�8�
����u�GXZEz�$\ C]:�	[vXt�ݴ�?Q���?��������?)���`kPB)V��yq��?gobMb�}%~�j���?y.O�5���O@�{��Úx��=aP"�j�x@Ӷ
N�������$�	4Y�v!��͟��	���	��PVA��*��	IS��j�%b��_�D��Py2+��O��O���'�rA�":Ed)5l�?��IP�*D7u���'/�`����X�d�O����O���O�󄃋]gpM�"�&��q��s��I&H�2�	럼��ן�������O�TA��M��ؑ�S�j�̘bٍ9P�6-�O����ON�[�[���	�O-&E���T������/�@jբu���I�\����$?����M���a��qs�қw9�\��d���?����?q���?Q������OT�:�<��AscꍁS�����J�jl��Z2%�O��D�Of�$�O ���O(��K�ɦ���Ɵ���V�\�=�����!*��o�P���<��WyR�'���OY�0Oa�v'W�u�<Đ�	�8{�l#D�'7�'���'��0�Iw�2��O������Z��O_���	T��H��Hf�O��D�<Q�Nb̧�?�,O��/� ����n�-*{T��b�	e5pE�'���'��T@!Kq�z��O�������O*$��=9�n���r�p@Bա�<��e\ڼ������|�ɟR,�6lƷK1��3G)�.WPpe�'v��;��j����O��D�l���OR���O�1b��#��0�%��5�X��E�OZ���j�O�ʓbs��Χ��'���ƍ����&?x��JE2+m�f�'�R�'�Tm���Ow"�'"�'�b��v�L�A+RW}V-iP&�n�r�'��I�[�|�&?��ӟ��I�2�tl	T^�0��q��"�k����ԟ$���M����?���?�C_?1�f��@t��Q?f������P�@�'�����'���'��'$rP���E��VvUh�Gі5�z��3*��lN�s�4�?i��?��p���Ty��'{�8�[�x�eZ��ÕL7����_2�y��'K��'�r�'z��'��!`���q�3M�gQD�p�c��R�Z���O��d�Ot�$�O��d�<��Q��}�'$ -z���5����Ջ�:H���?y��?����ă�jb��&>��	\�-�>���i ��ڄ��П��n��П�	,Z���	o~2�M78y�dy�#�8f��Hr�P/�?)��?(Oҩ��^�ҟ��=j�ٲ C�5X�;���%��$�����Tr�,��T'���l�^����Z�6�̩��)�{��ĵ<�4d�>��W>Q���?B,O�9��֙E{iҦL�)2�� V�'���'�R�8��'Pɧ�OX�m���L��t��.h"�����q���i��'"��O�2O@��K
��1�֟)�2��!�A�v��p��#��������ۄ�����b�p�@����M{��?Q�zi�QR�x��'��9O�<!�W��`�T E!A�(��F�'q�'r�iHE���'K�;�>}8@i
�\H6�dK�a��	���'��E�BN�O*���O��O(Y�'�X�{ͲB�(vwx�t*�<I�E��<�-O����O��ķ<QH�.��5 �fI� ��X�0d �&ٖ- e�x"�',B�|2�'-b�Ň5*�b`B�0w#[� E�Y~0���'%�����ԟ��'!�@u�矔i����0#�t<�s�G�8p�r�yb�'�'�r�'� �P�'X�8CK��rɀ
Mʨ���'���'���'��G�<eXڴ�?q�_X�<�"�>&
9{�$F�
)@���?�H>��?�%�έ�?��Ov����pRi���\13�-�S�'���'{剷7j&P�L|
��b�/�B"D�A��
4���S�+Հ�䓴?Y�#|d�8���S�U��i^:D�q�E�6�*�@
����'vr���p�P˧�?Q��D�剹RN�3DCJR�\0$��o�J��O2��à8���D4���ݔ{��uh��T�%� Pf�/��u��j؃_)r��rL�yx���`�O��UV&�|[` -�<�;OR:ē�+F(��U� ��Bs،
�J���n��M{g�'G��'���]>u�	�$5s�� p���
��hcP���58A�����;Z�H���5�?�B�S�|"�d��aE��㦈�#H�6��bDT�<	e
H?2r�ũ��+j���a�JBզ��g&�7:3��*�<>�@	 2�tr�C��J�X�q�⎑8����m�=,�nY�`���K���M��i��l��5��X7.��Z2�j�#ݞ��㊉�����a�F �^��f͋�������w��YJ����8
M�v�P�;v��T�{��'��  ���F���'.�i3   �?OҸ0z��"M�2s$�E�`�)G�q�D���ѵ����Y�<�s�
,�T��wE��}��9�;x�!�QOQ9K6��܈	hꨳ3F����O��	?�zu�F��:{�
�A �U�O~ڝ���?!�O򸧟�c��K���2@Y���$��s��Kѭ<D���G�G�&)Y�k�3E����Ũ:}��'u�"=�'�?�4�$�*��m�|��j�:�	5�Bl#}�N����'���'�2Nyݹ�I��n�$W�|��	��CF�!v1C]��O�{��`f�����Q�'hġ�i�6~�`P�G�V3�@�AQ8��a�'�Ov������u�
9A�$��FɄ.ט�بO��#.��5�l���MV��h9P�ig�E	���?��d'�D�-j�@�:� ���$l]�K�@+D�C�A��Gƀi�� 8$�RL'�3�m��eyrb����	��Ĥ������X�
�n��q�1h���?y��V��ܒ���?Y�O��`#�L�%N�P�����V�a�#R�F'�)�#m�"�����'wF��Ы9��4����	�7`�8^�2�Vf]#j�4*��'�4���?�۴P#6uk�]�	�<��#�5D�F	Ey2�'@i��d�L�1�o4t}��
�';�|�Gɛ�I���@��c2X��H}bV�,�F���M���?9+�"�{;�*��$�>�n�Z$��[���O����O��ئ��$܄]�����T>ٮ;X��u��$8%�\H�IL�)�>��>q!�G�������?��?�a7 Э�!Wo�66���%K �I/w��� ����ش�?1K|�5MG?��ʠf�!c���	YZ��O��<�M�U���0�$$��Q�Sb�{�����{�-�$�2�xn�Cj܀!��X� ���L�)�`�$�O��4�vT��.�O���O�6-Y�&��I�Åg����OT%�JEj2�J�wp��񲀕��?i`ٟ�b>�}�r4��ƫC���� 5�V}��,G�^o�<z6	D�7���l���� �,��D�!�n5���R��rW���|J>I�>�G�OZt!J�oěn�8|�Mr�<�����FX��l$0�bgܓm񑞒��Ÿ�m�oI��b�OUy6�Ɵ��/����	şD�	͟�j��2��w�J��6��< �*d	+eMI�R~$A�b��b�t-�#ƚ��uw��##���X���K�@,[E���B+֌K�)�SR��4��:|�Ҵ	�"cݱ�pŔ�\�c�d�7g�l�*�"�A�?*pļ+��@�uq�������nӚ�d�<�����
H�2/��g�.Ĺ��ӕP;V��IO}B2_ً����}��� bE���(O�mZ����'�(`�h��7m�r�Q�p"�08� ����\*�,�I��H�Ia7ԉ�I���Χ���Vg�5+�܄�ҡ%[���ÎѰ�l$��Q��4O�Zł#}8x�;E+�#]r�	TE�;OL4	@�J.Q� j�G��@��h���$D� p¦���#`�*����-ȱmL<�#�,D�X�G�����D�ȗG<@ P�)ꓶȟ��ƃ��/<XezQ�V�@a�pCc��M{L>I���*-�	��l�O��MٳJ�_^j�{����*jAh�0;�2�'�2lZ� 疩ʀLN�i6�(
��_ :���'�u'��$U���ݕlbv1�-���'J����[�I����eI�F$`E���ԉ�,p�zX ŏ�`t�0@�f�{���ٟ �	���%>���J�4E����g( �>a� 0eS���'���Y�pzaMR�A��xB��,?%�H�C6\O`��=���܂j��1A`J��k6�3�[-8x��7	~�X�$�O��4�DQ��O��d�Ov7M_�U�:��7܏��y2l��C!,5Z���J��@K���Y�ԟXb>�Q0��p�oD�f<ä���4�|qFEޅ.�(`'j�|�P9���QCIY��i̼���-j8���_2`��{q��o<r�D���D�U��ʓ�Z�t���)�Ġ:�!��Ʈ@�b��%���o/铦?��i>u�'����p���*js�����H��X=�?I7#�m����?����?�c������O�l��Q�����%*�h�����M�Ŭ������%,�Q��'`(���%�kc��{r�
=�i�v�϶[ %�$ T�����0����u��wnQ��"�ŕ O��k5)��x;d�Xs.�/7\^	H��"���g�����<�����"������>y���!t�]@Ϡ��Fm��@R�S�b��8Q���n�Ey�Fl�_��zS-L�$n��E/ ט����2&�Z0��ފ	�^��	��l�	�������Χߐ��#�U>��6-��D����&�6m�UBH�=9��U8��J�G[1���\9D�4YP$
W����G��3\�i�vH]�~ǔ� ��I���?�"i�០��4)r�Q;a"�^���ɦ�,x�\�)��?I-O��$'�)��T�z6�@�,��P+b�I�N�=x!��88���)��E5d�y�.͟*Z=z�4�?�*O�
�)��9��ٟ��Ox�]�G� `3N��T(����7�"�'�BdZ#�npRK(�Z�a2��4%����  ��nخy+2a���>n�ا˄7_n�M�>	K�z?�Q����05* ����6%޶�tb���sgE�R�q�
�b�0)���DX1L�b�=�'f��H��ۋФ9ڤ�ߴq����OY�(z��N�|����0#K/A�B����hO�	�@�k�T����Z;& k���>K����$ޔg[7��O�$�O󩋯�n�d�OV�$~�ry!��D0�^1CP��.�A�Z
5�
��J\+3��Ffq�Ę�'�����O�.�|�� �@L,q�-�FX 8��"
�-�mp���D�q��A�=H��iW���{#�̧g*�X9x�)��E�:G��1����П��'4 s�����{W� ��c��΋+���O�w���'Z��P��%pȔ�J�,�#L�U��{b+4��|����MsׅI	�T葢ڊ>�Jq��,wuҡ��� ���'���'B�z�����Η��0`
�!%px�Y��ɝ˛Ff�rk�a�&"C�o�z�D3K�|�#�!6� �qN�M[�ϑ�"ĐsW`�p=�Ń��m0^� �
ƻE���w�O�C���O��l�����?!���^\��)��7Hߜ���/[v��������Q	C<K^��p�K�{N�Fy�k�d�$�<�CܶY���l��!#s	�?�	+f��c��a��������8���I՟��'$j����Q��p�-�-^�*����N,G��U8�/��7�H�ɡZ�,;7*0ʓY���x��<S�Z�+��W�̸���k։
V�^�+@���>����0�^~
1�I2�Ms�
�+H�|!�U	N Y(ag\ 1�B������$�OR⟒��93�W�������A�@�"O ��1���lF��p�	�g���"!B���$�<�v��ě��'��^>�#4�Ж �k�fT�+�(�Ĭ�.
�`0������ɖ`�p|��JV��*� Z%Z� ����ݫu4� �(:O��UA���dj�b���m� �0Q�%��]��9�#�S�v)���ЖAd�9Ш�2
u�J��gtH��}���?�üi���h�g�? ��c��8{ɠ���K�E�����w�Iޟ��)�gy��+y̜��vJ� 4��)���-�~��i>���4˛Q�����,���W���
r8v�	R��@�i�r�'��O���@A�'%2�'���B�G�X�A��r����8Ad��W�<]2��l4Ϝ��џ�����*4M���Dk���8�#у�)o��pC"�w��dpC��>!�%c��M���z)̻U"�zA�m��� $[�7�Xu�'I 7������c�>�nZv�h��E, �w��U.N����'�ў�Gz�H\+Nx�X��׾]�.�kd�Ɛ��	�ߴ;M�V�|��])k4���iln ��D6ghp�DA	V"���'�f�i�*"=ьy�T�P 2@��S��1صC���ē�p>AȐ]��q"��8ZP�]�6cK�s����r!X�*�.�`YkS��/-9Z��ȓGF�q��AQ�B45��,
�@c�i��p-�A����,8��j篍�6C�5��'`$9Rī
�n�v���+^�>(����t�ڤ1�ΆS���q�3_����|%�
�lB<�5�w��`���ȓQܹh1
��A�A��mX�*���c��8����1�^�S�ϕ
�p�ȓ}5
HA7��3b������dV�)��r�����)��yz1�Y������U�<�{��m|䭫�k�9^�Ňȓ5� ���z��蛷�S51���ȓv�Cg�? T�sJ��j�ȓc�$���^'V|��/H�6 ���XV��S�E�R֠(�7��q��/�����R3{�Ne���N�l1�ȓGt.qe�k���R�s|���<K���F	�?E��0'�S �Є�b�
�@$�w�򜐦e����ȓt�>)sbʑ�]̈W�!J����"O�2l	HfL���
N3�\P�"O�EHSI��vX��˒ĖzD�S�"O�����$e)v�r�'�� ڀ�h�"OZ�I�y�R�sW'j�b�J0g'D�<$Fϟ�LPQ��&�H��`�3D��!6N,v���zT��FFf���0D�Ԓ3�^$T�B
Meߐ����/D���piQ
��Gh�[����+D�Lr�D�B�HU�jT"k����5D��Z���*uz*� �P�` FI�6D�\�q@�,qИ`1$<�N�kף7D��C'�V����`��P�Z�r�.D�x��Q�^ %Ң�O�&�ra-�p���� iі��O�PM��ؼJ�2��n�OT�
�'S(� `C
.�~y�"�	<`���'�T|�K[�(6L�O�>��-Ūu��t:�e�����)D��q������
��|� ��XyRj�A��3�B����	�Ei2�ǄD�L6d�0�&��td����va�c��C�@�Xթ�n�7C�D��!��}��:����?A��X�'��P��C�j�aچh�}�'�V�&��|?D�Ȁ��x��%`E3�k��]26$�t?�C�	UR  a&R�KyP٦$���7m�"��dB�i΂.Ӛ| � �r��M#"��Bj�4K��	)\� ���P�<AEl�N�b�{ց
o�V���ӐVǴ��;e�����X�(����<S�fm�tD�1my�!�4�
sC ��a�X�/3��
�<�O����+�
w�6��(�m��� e����,1�@͍z�r��Fi�<���\44���{��0E5��(=��ظv�X5Nt�Ӂ	�
� "=i5�T�rqthÕ,�
#=Ą�H?��5l]�Y�(x��kB
zsRD��o)Z��%����}+��A�¾�(��	xwz2�#O�Gc$:�윋O66��A`n�q1ȍG��[��F��M����2�D];A~�i�� H��qO��Lޡ;�瘷[�48��$�^b�H�Bd��p�8�lZ��l��,GN!0G�R(ʲq�@]?�	8I�Z<��	��p���ź�T���N�6l��SIF6X�V���'�l��D#Z.A!���!�!�:�X�$Z+!HLŨg�Y:�r��'�^IJ�� �� ��x�a�Jf��\���	�@|��� �DdH����$bC7nZɪ����Q���A�BU��'lZ�z��O<���
T(a�{R�ɱgn����'�F�:&AM�$��c�V�"~
Ď%��mL!J��1�$h
��'��-�g?I'�tMr�S��uB,���̂��D�5f;�� ��
@�3�+�2�I�]�B8r3�S'%�@��	��ԍ!דP7�p��4��@�W�EF�|BE��4M���H�O;��SR��z`�B0kO�ɑ7�
1\��|a�O*O�]s�m.�ɘ2��0��'ŅT�0`æ��h.�b�4h�f͊j-��!���$S��}�U΋w�pٶF�t�B�/f��*S<S�Q��Q2�j� Ɛ X�6�F"�<���L�Dy �T-�,Yb����)���A�'$� 15j��z'6ؓL��a��4Q����ܠ��Ӏ>�^�V�'��AB��Q-cc�L��g�*tHภ�G����C)�V��=��.�M�G��B�P�iV#���fH#���A�<���ë0�"�0��]�5p� 	�{~r�źIl:Ā�!S�s�$`HU�d�O��(k�69#���7dT�~�>�Y	�'6��2/ֲ8	��h�(iX�#_�	���2M˓ �\D��S�Ϙ'�� y�H��T|R�Z�Kq,�Q�'��AW��5d�)aa�pT�k#F!jL^m+֯�PŃ`�E|������TzB����񢐸d&"O���c�N�y�����%�7^�奘�C�tyIF&�r�ݳ�D�1n!���0U���J�mL8@�8���m�)v��I�r�VUbSOT���B6�P�Q>ɋ��ԿY]�I��@���I!D�|�0�H�dgr��!.б~��/�:A��OIan|��n�x���O2��ĝ�"*�����7��QR��x�aO�:vB<`��ޡ@D��� �7#l	��eX$[��!b�/	(�i#�'"���BȜ�l�z��W�Wr�yэ�^�E�֣�z�,��s//��y��lL .��P�nГ'v����f�<���ʛ@A q��j͵
zlPxP��]}"Tb�e��c |��H�e���H�p�Ȃ�4heQ
eiG�:Ը�"O���ㅵEwZ�ڣ�[+W,D�ï��z9P@{D�ū<���:ub��?���'M
��f"J�aϜ@�PN�����j�jmh%X"�L�Q��Т��]8z���r��;3� s�)ɮ�̡+��H��
`�G�]�Pȸ�/��U�!+`$,ړ1�H�q�ײ?��3�Ŕ�s��O��x��nl�03Lܞm�y9
�'�q�S&&_̃!��Z�<4k�4/{���� �};�dۥK�c�¢�s���7#4x��d���{�����*5D�0���,���FF��8�n0s��0M����B.�mc
����A^��pc��*׭�70��@�
�&\R#�.�O�XPV��u}l��v�Օ.Ӽ�x)ˍ:���U
�'\�Hq��-r��Ĉs�'_�)ҦR5{B4�:��׮8u��X�2�0l��S�Č'o��DJ� ,Xx�Ñ6��p�' ܌b L}�κ@��5j��'��x�, �>�1��|�����Α�Ei��V�a�|�t��O]�Z�6�)��d��NgN@��Q�ƕ�� �$bR���8�;�����\�(	�@&?M('���Q2q���^9~��`u:�<��tu��e�vxM8R:#<��M�1L�"љQ�境�I�<�nދ:'�yp�_�;*���OrD4
� <YxJ1OZ�d� ��h��2c�r㮀�S�f�	DꁌN��cC� .�0>�*\8!\�!HA�W�j����G�k�ĉڴ
>10�
ѭ>��@�͕;wM*�0cQ�%����yG�2m��Iҋ�%�(�&`�	߰>Y��@�:86-ݺ3:"�Y�l"fD��-V�ҥCS�pĮ�h���4������96<.�q���|�,U���{�c�i�P�3ōX+Y;�\PU�2��������6@#Ƶ����r ��b�ٺ�-��i���p��(�`<�1��A-�)��0���2���p(�đ�k���(�(<u��X��c\�R��;|�,��b"r��H��C��L�p�}�'Ņ�v��P����4;��)7�P�xTRx"�i͖ʼ�"��V��w�'mvp��1,�/5"��P�!�O }�a�G�<C�u��2�l<ȡa��r��3ĝ�*}�cPF�A��.�:J�M���^0�t �1��3��	�PD���'F����8JU�'�I�O頴3V���9Ci��,�śv��:`��P�sP�q�����?n[�K�/ϖ?HI��M-���慁��M[��Q�<��e�%�^X����g�V�'����UH\��j�OJ�*^�I�É�_�6ɉ�A|ku�Q�u�����nf
�`��4Q� h�n�F��f��Q����4.���G	��l�� ��Cc��l�^���ط�.k��<� �%r,h�	�|��f�L2*�`BGBu�XT8���p����ADL5H�6G�gH� (gI?�O��r��&K\$�'-��q<17���@,XA�G�qy���Ms���&;#�ɓ�·�����w�ͨm�V�y��\�h�5��D#�@:Z� ����ᚖb|Z��u���1��9:�7�ϫS�m�CC�G|��i���*��B�k��?9�et�ܜuy*@A��ٝ:���	�����:�QЬ<@L��]�9�E<W�L�x�m� �vt�,�,7i$���.�P�@-Ǘ,΢�*C��W"}a"�&�lH�r�Z�0f�;5`T�9�� �$�{W�I��v��zGg�o�X��˲n���j���+qx,��?a�A۩
����S(�Y#"m"��"P��N_6��	���\*����N��s�#d�P���
&UF���n����'�H�ݴJ";5�f�U��LJ:5��\�!C"�Q�!�O�5�2-� ,Z�u����<=eD�B#�&�p��[@�	"�6MӶ{�P�WGM�9YvXz3���I3.As��~~�죵ɗ2P�T��/O-L/�:��D� <���4��+ `4h�GwᣧԢ:s���Ë�
�bxa�I�w�la��&I<��� JW��7mו��\�#J�|-Dx"#A�&였�F� D���-K8�Mc'! ��� �d��uQ�QQw/� s`������Ċ��M�!P�l✡�f�ņKg�# �U>�	��.X�iPt�T�'L�x���Y  `��L��^��a7dJ�X��%���ô;�x��wA�L�U�#
6HoZ�p��	�>��%uK�p܎���mT�������'����M� Tܶ�"���+T�P:�L-#�b�'�i���s�J�LK�ũ�'��\��hP�<\��d�_M��@�/Z�Y��F�t�xpCaJ� =j�<�*:��PN\�
i2p��S"Dj����L�!���C�%�| 6\�ԢG�S��oZ�z�l:/�/�J��AKrJ�� 
&�Oz�ɷ�;N�dP����L�"$B��O�}*Dc4k�JPZ�Ш4��c�c�&C5"/��q�J��?�<�0��&hA���F,?����+ӎ 7"��!�t8���M -\�v ��ST��3���F�(�b%9cx$*U�L9�X3� �/Z�;6�"RW�4��Iu�Q90N��0�(� d!H�|T��5�OZ]P�5����7H�N|[��u.�1�.	XG(H�tH�435���Ӛ0��5B4N�\X�@�|<��I�e���b�M��$�8C�\�r"���D h���A�e锡Kq��v�Y�ff��קGo�\8p
�}Ǟ(	w&g�h�թQ'
T�b,_�&H��E|bbڼKvex�#JiܹP�����G�11��Q��+8�Rx�Ɂ-
�fpA�C̹̾��O��UZ��\CK<@A N�Y"�=�'���B f<P��t�s�G�gP<�T��o�{E�:�j@+�@1I����������a��NuD|�̅	1����`�eO�Lx7d�O�Dp�`�(b��3�V�+~0��A�qh�ZրI�8t��ZG�(a���,5a�y�q+ϐ������j�����ÍY��/��2B`#T��6Ș�Ѳ��9d��k�X:i��)�#��*���k!&�zX���I�w��I�êM�O��� ��"}"�U�m�v���ԇ;�,E�Sq=�ƚ�]�l��O,Z��ו,��"£O)9�l��'�
�K��o���¡�-�P�?@WX���H�G�e�ge�c>YɲG�
�y���J���ǅ�xUj��� ��x�ሲS�h�1Ń
����3c$>>=� #��F�P;�\q,�7M�Ջ�H�Q�d�Ez"&�Q��c�ϙ�4h���)��0=���6�^�t��&2���
˒�3���(?h�h#�5�:ujI�q�a}r�Ĉ6��l��&���<1Aą���'"��tmB�i�����e�eRF��K�M�+�L !k�){���"�N��y����s���c���.�`�8�L�6�!(�*��:%���B�	 ��tp��s�����G����u�Ub8I1��+D��js��6*~Hy!���YG��4��<4"��E�g�n�Ջ�ɰ4�f��o�$>���������Mۘ]� 5!B膂 �4� 3�ʠټ����''���&`	yi4��!GV�N�u�˓0��`�Wc�l≓\��ԏKl*,��$�>,�^C�	
�H@��W��>�
��ʵ}�*C�	#���)���W>�	�,Um5�C�L�J���ޫ_Z�\�'C�p�!�d�=����)׷J�h��Hl�!��˸�N��]�2F�R".!�!�T��$ܘ`ѿ2)��� &лa�!�D��!��(�A�>M���2�ES�9f!�F�4���l\#M�T��%A�q !�dZ�+_V�`��1
����MZ�!�d�3���e`�- S�УCL�p!�d:V�ܻg�lY���G��!��
�51���(��*1��;����!��4���Ec�2)���Q�]/)�!���eA$$��	�� q�T��H��=�!�ݪ�.�:"J�H��Wi��!�d�8L�Ds �$]F	Zq�Μa�!�Dx���O1@�-�	I�XA!�� 6uB��9i�����D�L�2XR"Od���ȉ_��4��!��Z�x��1"On�	���i�n5�b� �{x�i�A"O�h�"s/:�fnOu�A!"O��\�6�\$�� P�BaȤE"O~UB$IO�,�*7��!5�n��"O��1a�dC��S��u��41�"O�͉a(��yþ!�ٲ;���+�"O����f�D��2�R<ul�Z�"O�]�ӏЍJ���+�0G�`K�"Ov��#�mɘ���3��b"O4��	H�{����*��.}z5"Obe	��?�������"OD}���Qot�Ben
�e
a�"O�����[{P���D�|{DoH�gp����bi��`m[N�Sa�L�[�!��M���Yp�@�d��E��K�M�!��T"�aF	�_(-��̏�O-!�O f���k�
6Lx��c�X�,!��۟3�Zd�]C�T�1邹�!�Ńi�D�rJ '������{�!��Y=f�:���6y�|��E�A�!�����E��փ[���*�G�!��P7;6�����_��;���!�D�<L*[a��;W�Dq����2py!�ݱO���&W�rܫ���Rm!��+[�Z�$�:׈\��U�)R!�$�����������<j�cO�C@!��8w�N|�_2 �2)[Gǒ\3!�� $\8C�E�a��|���eK!�$L�z�h��h^%|I٣�a&Pi!���*�2LR"��g_�D#�H�zg!�Df<�`�qK�'6^�h!�� M�!�d�&_���:���=EM�	s��J�!�ĕ�B�b(!B� Z3��Aj(�!�D\��J-��E:C����)̮�!���\z����P$p�@Q�
!M!򤏴Rw��S��r���)3!�䅿)�R0鴍�	F��+��6E!��,}`�x�Ĩeys�.�!�ێ� s�͋�$������rz!�V�2�T|�Qi^�1�!�T!,	;!�DU�b��ᘑ
�-b� �XG�7&!��	��t�X/?��B𫙥n�!�d:W�L9C�ԅ+xze�WK�j!�[%*����7�?\~,�4k[�|"!�PGX�����+aSf�:�K�b�i	�AJ9�O��1��� 7��QP4�M<^�T]��'�`����O5�RO����-Q�%X��4�i�Z�`E{��	��g�|�#�1ET�t�'�Z����Ȁ�F����yaD%$^�*�K�u��9���xR��.>k��q
��Da�Scΰ|TH�c���|��C4~��ɋy����v��f��G��@t)ʨ�.J����Iְ����L*�41%��v&�ϖ'�h���T3�M�ӆ��&J���h���9��u�'�Zwڼ7�Ơe��(y�4�rP�%;z(�́N�'�d0Ѷ�Y ���%� G�,=����9���CK�6Yr�m�q��_Q����(y��GC���l�M�<��)�iGXjW�[�Y#�u��<aw�E�M���iG�ϲqHD`�1V����`ƨ/��̓)&U��(~p�)	�!�l��jB�nh��oY�20I2*�f8�q�`ޡs\6�١�Ҋ ��YU�!g��8�mù]
����@�u��s��I�p�%xw�V�z�p(!d!�]��Dh�'墵�����"���X�>8ȹ��n�*Hic%��0<��I�|e�q�RIZ;k
�Ѓ�F��{�Q�B ۢ*	�ih���(I�~�AI�K�%ʢ���lt���%
&�����b��?ǈ͈ê:�	�Y�XT��[0T�TI��y��'�hq񤄏%5�X$���E�0�)O�4#�_�wՐ��Ā�	�<(�gA]V�j�{U	�?jL��#� <<Q�(��y��Y�q�2bİ����3%2Y��!�5Y7�)�$NKX����O@;w0a�jE�z�=��FT�jx�AuA-Fe�"CԳO)ĵ��'���?�Dg���Jv��1Q�bQ����c�Qr��'k�q1˟/.C&��I�V��A��?;�|��0`�>����BQ;�Ǟ~8
����*�b�M�c�E��g�u�'�n���կV	���ۿqWB�h��?cL�8Jq�T dJ�i��,O�b�8�7C�3 ~�03� ���,*a���I�2���*��K�>OL��$N��x�v�'��gEd����ѭ�̦�Z�-C�g�DY#ƥ<AaFԝCXV�FGQ
^��Cq/$T�D6۪4B�)H�c�;<��D���hOp)�U�$x=����4an결i=*<���G����"LȽc�����Y�(o�/n�΄[����)���IU�k����\�5��~R�`R��cC��)C��ڐhl5� "m�vtX�0ش����>��'�6%X�k�������`pucNx2^�b&�Of�š�&a$ц�!2Ǣ¯`��=Q@�Q�I��@�)�5̰��#�D?qì�H�ZQ�U�Ւ/�Z���-�y�'� �iAMF�˾�h5��,g�1)���1w���v��#:W����N3q���-gJ<�w-�yH�5���7�l)ٌQ=xl�ׅ!<��bL�<�i��	��"�![�@H2kDo�It}b�ќc��QР
�<������աS&�;�Ì1E��}�lե> %`�	�p蚁� �±aNV\�(A"q��G}�:O,�w��88���@q,�X���I���	��_+�9:ã� e��x��.�e�B5��f�̈Ox����?o���#�O�&}�퀓1O�݈')��V��dJ�D�a�\
��D�!��@O�[q$z�� �I��I��?��4/�8[a��%���b�<cb2�̓UF81UJ� ���1".�/oB8E|���$Wo��c�N�=����l\6�|Lp�n�Fm��q�# X���� � ��gDϦ�:ך�0�i�	^X�`���D8�iqq��)9�&�z�D�a���a&퀏.��� ��E�sx ���)�6���� <Ox!���i(6����.2�X���,L��ƕ��#�/u�,M��;�[I��Z�eL8�"�P������I�4d"���kOW�������~Ԡ�O�� ���>T��JG.�=>�ur���??44��d)���^�b�Ø/��dѤ���b6s��}�ሏ?Zў|�^�.F��f�_�K����T��PM���f��1(��T�0�+,O���rŎΤ�	�+
�a�ek0��lGP���D
���>�w�E� 
�(5�s�2�6���0?�߾{�J����Čo�� ��b�%��D0AD \O����bْ~�L$��SZnt���%_�6˶IًsPY��O���>�l"�e��W����0OfTj&���i�����CC)kK��*�����eO^��4�B1T�Lɓ�T�d�O�x��F:u���ѭO��l[C6OD�Q��@�\]�5CUCٖu�y����)E'�|���M�A�l����f-��Pp��7	�e����*]i���|rVbX�o-�³DU�5�hH�tN,'��d�Ҋ���>rn�ՠ���)B��๥툁ag"=�|Z�iZ�Zw�x(���19Z,0��>t�a!�'�0�҃f��s������;�($K5��j ��#�1��I��z7��<٥(V8��PΧET�H�^��9OR�ac+ğ>|�0�<���+�D}��)-�<v6B��|�Ӻ3��M��x s��]9z[t\�Ge�&k�E�@�\ܔ��M�=Ԗl�g�'0zEkg��EMF�h��P0D���G�6���Y�l�<Ap���80��|
J?�)�l�
"&]�3T��1��rJ��2%j�e8���5 RL��BK~���[р��N1�\&͔@yrfU��Z���F�|r��.BB�J��D�hm3�Nl8�[�#�o����Ŕa0\1A�k}��^�z�,�r�M��4��`}��N�:
,�fT��O���h��U����R�6��Wi��,�H�º:�0�OY��,��5��ƤD�f�T�e$�a��k��� �IL!<�Lxh���0|�8A��g�>�+��)OMTu�G�5g����E��
�=��#��',m�eg��M�d�	�c��M��U�M6���i���4���S��囹�%)Ib$0�E��k����!�����(6�O�.r�1�K
�r,Yi'�N#B���)7��^#��i�Y�I\J��	��#�|UP��4}��AUk�d?џ��QIَ���k��E���a�Ab��A����g�ZEnZ�}���ɒ^�	�{,E#�O~�X�F�F!�ՠj~�5`Š�~�\ Ir�ݞ�	�d�q�,�	�?A1���*�X���S��7mߡ�ybh��7L��S�[�����A��~r��2p_��z���O*��1���;�hOfd�w* 7{��` ���"���xTnv�N�b�5L�DX����!/�T>��[f�R�Xr`�x��:P$�9iM�dc�&U�e����DJ� �ҫh-��h��}	~�J��)�87��	���y��Ip(��s�әiX�����)���(WC�'�:������Y�<0Γ}r4���#8���[):�Lzub^D��G|r���t)A��	/N͉F�4�y�]II��XT��0�\���~bԂR�<���j�>aSKBr�I�M��'-ؐऄ�9�)��[!:p��'�XAZ�+�+��%�y�ؑ��� ޤ�ՋL<Z(L���l��s��`��O��@e�4}��]
=ȣ=�$lR�[m�॒s�ty�Wk�B&���� ��=9�w+�q��"[/l�m�nۗPY�%R�'����
ד1	T�Bá
�1B�)teO+u5j�i#HB'%�j�?a ���}-�Ԫ%�i�:({R��8a�BD�j<�hE�/+�	r3�	~V�jQ�ׁX-���m��F�I�*n��A, ��R���&E�8�"A�����F66�C�\�n��M>Q��O!���`M�L�qnL�z�\[w0Oh��,ڴXg�ū�ޕ5�#�ɲ6;�x qG��1���)�0l?,m�4O��Ўy�n7�qv���K�0,�H"$K�5YE�%o�9~?�	��I�6	�لT�H�X���ܻ<7 -#�V�����2�LJ�l�b1�o�y�V`�ևJّ�`��(<�H�)�
��>Ԫ�ʂ�~�&���Pqt�A�I)~�6i ���s�h&�!x�<�!��M ���&�cdOT�[��]�U�e��c�\�E�%��bfh�vD�}�I�<Q3��?Vўْ��1`r>�@X&2�	�(τm�B�yN!.�����IW�Y�����Zt�Q���PrAI��i��qye�U[��z"�M%N�x�V�L=�i��3"�U�Ѐ ua}�i�6�I1�*sd�4�ɨl��~2"��	�h	JA
	���8t��B�DQ���fx��:p��f��-���B�̌\�U��E	�#)Lxa��O�ѨO���NYޔ�9�ʔ7v
���'QTE[0)'h=����
O(n&TIM<����\2M���(�&�� �y~R-E��x�I�R�m�k[(FՈ��>�1`�[B(�4�V�(��Ӡ�8ړ-��$H��ɐ���h�( �������O��	�)�ēD�P�S�S"m�6�C�ã"�	.�zx�cX0=�����z����&)�����ʁ*z���_�����Oz���gK�W��y��Y.z���Q��A�Uhs�'9\��SnVR�|;R�ݥ:�F(��AͳUv��C��UjmT)+�OG�'��=Ya/TYX���N��R~�q���3mRQ#�V�MEP���mV�kn|�O��8��ˌ4W��p�]
*dx�ȳ�D�3����eG#[�P�B�#ǅB���n��&�4�r]*PA�:s6�=���;�"�FKd&|���"Q�ޠ�'�N 2��E�iu���{�p��	�W{��ecAWg�����X�J0z�����䙋/ H�@��9�\�����m������)�(OH�O�hڢ0�>U"��*6@D�B�ǩs�|�y�'>�=�	P�ڄ�5�̤�)xm�{��Aï�<J>i���-�% �D�̎�:����>|�x|��+ڸ!N��QdvZt">у'�/P~D3�ٴ}j����F��<��f_/{��� Ɖ�e�z%�J@?��-� pΌ,9�#I�h��j���]�'x����:.|��!A�,	��ի�+�����ʗ��?�4�I�z�x��O$	�I� q���@,JH�셕:B̝�c0�]��4�ON�ȗ-�81 ��s�ɇ#JH�#�넬<Y���~B
Y~���3�Ԝ��eҚr� ��D�L֜�{F�'V��yBK�)ݎ�h$@�`n�Ð���E��� �X�����4\-#d�O�N�>��ݔO��a�'Q`-c� ՕV��
ñ5+ؤ[��dU4K4Bqm���z��td�j�$` ?0�آ�)��j\���-�U�A�˞*�٨�M�@\ҹS��hO��O�+Ҝ�JVAL.}��<��'Y���&�I�$����� �z���I|&�dAFE�)1�H�#�g]=m
�%���$�ĝ��)$�}"lK�҉R���/i8����VB��R�'��`H���#.?��uS>A�2�$%�@�e�$��u�&	=�h�g�'�46MBM�H��� I6pBR%��jU�&-v9ՊT�<#�'.�d�-����MK� +��i;�}�'�8o���4 ˺b����6扸&����
y�*��I�$� A����!���M)N,q'ƍO�|qZ�%ټ�OVtGzJ|�h�,z�&@�GJI)|$��H�C�<y'��QLi��[>`�z�E�s�<�A#1�8�g�@9(��8��DD�<��+2[�+�Ϗ4X�JdHb�	C�<ㅥT��*dǇ{�Ja���Wg�<Y�!�
6��m��D��	��@��Da�<��R�4Sju�e`��b..|H'�F�<��d�fb� 4�?=���x6l\M�<��B۠|+1�K^/�M�G�b�<1į�3ƨ�K�={LF( �e�<�A/ӥ1�Hm�s==�fI�B�Ed�<a��4�������H%9��"O�P���ˉ�2��D�E�U,x��W"O�A@�!��İ��GY&.�$��"O� �Q�e�L�e~�rǤT�6��"O�,p "#~�α�惐�z�,��""O���I#(�8�U#@�w�j�bf"O0��N�? Hh���!S����"O(�gf\�p%d!�%b�R���iC"O��K4N�=U���� �{�z)3"O�� f��CК�Cw���V+v	k"OP�C�DŴq�"M[�E��G9�o,D�@X�ĉ�h����qjk:�t�)D��;�,e�E)�KGQr�j7)D����HΕ=]L՚�E&i��F�$D�p�SHT!\N��"-�JD��>D����X+M�ls�I��i����#:D�@5��5i�X�ML�7��(��d+D�PS	�	9����-�+kآXeH(D��b%$�$ �i��)��َ�!�G!D�	tM\�3�����R�x��f"D�T scJ��LTq����,�p�P�*O��Z4��6���vC�>Z*���%"O��3nǛn%�1炐�9&�9�"OZ4D�P� @�/]bs���D"O�5�T�6�r00��8\���"O�P`'Źk+�Id#֨���Z$"O[C킴t�0	�34ߌ�#�"O8d�Ԡ�v�Y��CL�T���"O`��O��*�N��(��"O��S�2̳�*X�B����"O�!��}*�0�jIPθ9""O"%���R+U��Q�i�!9!�)�"OҵS�ϝ�
��)���.]��C�"O�Y[�Y нSğ�F����"OnD:� �!�bI��T�#�0�c"O(���Fh��ʷ%_")��A��"OPx����%|I�OZ	[s��F"O���� dm�8�M�/����"O�!�#�;3I�<� ѺL0`X "O4䰆c�
�����3�:q��"Ot�(��1:��a!b�8-�$"O���.�-Yp��j�nӺS� ���"O�j���1�Xu���ƜQv8��"O�H0DN��S�ܼ��ܟFj2�H0"Oh�����;��AAP�>6\��D"O(0� SN��Eȳ�ڵ`E̴�"O֑�@�$Ѯ�b�ܭ}��YIb"Oa�`C)z��2E��"Y����"Od�U��>���$8U?T�A"O�94�)a^��㉅%%!��0e"O�ܨ�L͝!�L5@���h�b"O�p��#Ǹ)�z��a�| �%�G"On�wf�"4~��EƂ*HLh+"O�Rl\�\���N�}]���"O����
+���#��ND�Y3"O���AN���i�@��7]UjP�P"O�Ѐ�v��{�NQ��EPw"O����1D:��x`�?��M�"OD�Al �-�X[�eH�I=N��"O8�$�B"�@��E}:cw"O��k�+�9W~| �U6-�a�"O�1ǵn/(eY���!�x�"O(�ׇC�R�L4�5L�1`�l�t"O�ÒJ��TѴ٪&�	]����"Or{K��-7��ے៮U�0�q"O�m�5�	��@$:@�H���ٺ""O��X��P��o
x�r)pO(�� �xe�������Nכ�A%"O���"\�T�fM��Ԣ����'�Q��j�F��Y>��e�k����!D� (N�h�0$9�)��s>��sW�>D�HR�I�TAd�ɳ%��l��H��D!D��CC�t�
����)����f D��I!HV��p�3��j1�t�6#D���,H�(����`*��f�x Y�G D�d �m=kY�9g/��Sզ�C�>D����
A�lߺyrr���g��%:D����*N5P���<S�\ ���*D�ȹ�߻Co����-��	SN��'-D�pH�!0B��an)X�2�QP@+D��w,�OE��`����{� �X�&/D�t�֠HG,`g�]�8uN�R�-D����g������"�X[B�I�,D�|bt����Nи3�ŉe�JH��+D��ȕf*t u�&F�W�)D����ذp>X@b��	C����l-D�0�cl_�!��TC����pr�>D��K5��lc0l��_�Y�����:D��0����4��5BC�D�x��3D�l;����mD<���+5{N���3D���G	5e#�Q9cDO*~	DQV	7D�`����X��A	�J�1mRx�gK*D��K���$"�5���P #�J\���4D��[J�<q,>X�pa�1;�ɱU�1D�LY�#�/<.�1���S�$/(	���-D�L�����5����ޕ��g D�,��b�8L�t��?L�,:u�8D�dRP�I<�J����T�h�e�)T���1@��^�>͛@�بz0��q"O���
V[N��w�ѫsdZ8�"O�y�׃^�P9�d2$�W�M�<��"O,"����h`���r��-��"O��S��	ȺC"�"�rԈ�"OB���*�qęk�i'{�Z="OD�h3�)Ln�P�+Gd "�"O�@˴cJ+4�� ���}e���"O:����� ���a�F�#]0��"O,�����mH�(�� X�1T ���"OvTۄ-� �T�����5� �"ON�����R���a�*� Ʈ���"OZQ87琛P��	8&���h\�q""O�Qс�?-�"�{cĻ)��̱"O���E�:tY&"O�o׬�K"Ox,�e^<3ք)��ŮJ��{�"OvM�Flǰc��*�._=B�L�"Oh5�`d�Y�R<B�#,���Qu"O��覮�6zXp�Lߜ ,xX`b"O�<��Q7p"��k�����"On�1�釐O�d�`�9T����"O�=�I�'vҩ)���3�t�""OpT҅�<����'T+e�܅Z�"O*��j��5dE %�>d���1"O����
)�CS?`z|��U"OR�*`E�DQ($����:SH4+�"OpA�B�-��+�l,HPػ�"O`��eD;3d0Ö���˱"O�c�	K9(�3���4x��Ur�"O.���je� �BlʊK<���"O\!��̚3f'x�"S#K�8��"O��0�1H0�x�'�R�y�͘P"OnY���H�6�
�p�/� ��w"O� �1Q̍�X�(@z lS�"O���
�C=��QG4 Py"O8�d�ҏ����p���(�ԕɕ"O�s*ɀ:��'�r\A�5"O\�٢-S0I:Ԩ�E�6cLd��"O�� �	ς�J�o9[��8R"O�Ȼf��7,i����t㎝��"O�}P�Ř[����2�Ǻ��e+A"O����Ĝ+�<9���T�PA��"O�t�6d׆i�y(�a�3��$��"O�Hj�M{���a������"O ����F� =b��T���"O8��-�F @ �(2�0�9�"O���Ǡ	�>(�fæR�8M�"OL�h��.%��4E�<`�p��"O��UmD�Z�)&W D����`"Od�R��|\�}wˀ��<Dv"O�U�pkJ�,���#���.����R"O45�*.]�hI�iW>y���"O�,	��3�%pW�(�@�"O�#D�(�4HcF
�Ul��P"O`3��V�qSbi��酆]�%Ad"Ot=����g���S�g�BR5��"OVe֯�w^��Z�`]!�:�"OFY�c۾K������ZM��"O��iK�	H%rX��戎\��}"`"O��%�� ������T"OH��VN׏M�X(�rC����+�"O�PAw�?Pqa#����V4ѡ"OF8{SL�O��P�ri�yRI""O���r�F�&Q��F���4�"O4�Q%; Q@K����	�"O�=��HSlj~�)6��
9�&d�b"OL䏌#�Qc�lX	�=@�"O�܊Af�5O�L��K�&YC�%P#"O\���*Ԯ7<�iP$*5��"O<�
T�̈́���9r�6��""Obɺb��� ���e�r���"O��qte
�2D<ͫ�/R�$w�m��"O�0@���.r�lA���.M��#�"O�(c˗�E��-�G�ϕ18�y��"O�5:fC�3��\��eӺ .�a�"O���QnV-Z���*�36*|:g"O.$RPJ|�z�"vG[3�6%Y�"O
���KF�^f����G(Ob:�*O*�b�A
 %�h�bN_�> �'N�
�� ��踒�6�&��'J��%��#��Gȯ( ��'�,�酫�����ِ@Ғ�q@�'��rrJ��zCDd��P�s����'�J��m�J�Qh�Fʢ���)�',
���)�LJ������Lb8��'i��J&�HW�0�I"��x��',؁�V�=�2Uq�cJ� X���'@t�s�eV�{b�;e��	w�8h�'��q0���6v�QYD�	9t�P�'�L��@�8+���'�?_��
�'����@a�(  �3���S-�
�'�^��d_�i6b]��	��d0�
�'?8m��G�]�茸wnĎG����'~b���A�3}�1�'̛�E�aP�'ND���� (a����@�
.�@��'�B��A�:|�ـV��)m�1�':d|� ��c=�u�B��g�<q
��� 䥠!h�9e��y�Dǹ�ع�"O�A�7�܋`���УX�n�z1k"O ��.��8�t8%�ڟZ��pX�"OR�!AH�A64�Q/_���I�"O��a��W�'��a�%Y�>J����"Oĵ���4;�X,�7��n2J��"O�aAL�H�h��8"@���"O ���%<XTb�,�k�Q�"O�hS�H��S*2������H&"Ou�!bR%?�|i@ ��6�3"OŨ2i�?k{ڰ���S�TVf�st"O Zug�9}�2!����B�!��"O�%0�&�"l�0'S[+��)"OZ����	>>s��І�$+�F䩳"O<M�Ѥ�9i�>��҇�>,>(Ĳ�"O�x� 	�3����E�cNV�{"O0�w��y�(,c���U+v\��"O�(æ\G��"�	I@��s"O2a[siX�i��Qg. �`�=�1"O�|�E� :� � ��Z�Q�0%�A"O-4	Y�<�Z�Y��B��NDK�"O�A�F�D�}Ȏ��!�x\c�"Ol�e�Ny�ݛ�g:�BX�5"O�l90g�4����uGq�ؽa"Or|2#�I��=Bp	w� ���"O���g&h����_ A�({�"O�h��]<#��#aD�\H�D"O�����A:�ء؅�Hb�t(��"O�ł��W��([�`��\����"OY�ḡ: ��i��� .���"�"O�|.���c����ݠ�yx!��W ���H�i��l1�k5�Ҝ.O!�$�d+J�:��e$d 3
ԏZK!���n0���匲~����u�L�%�!��*�@ÀI��CN��{d!�#K�xҶ�#���h�#�HQ!�d\$:� ��HׯG�ޥz�A�7!�<$�X��b�SmZe���b�!�ĖRS�q  P�.�ڦ+W*�!��4/���+/z$cV��?�!��5Q,�� �"og�y��@�X�!��Һ5�q�DE��~��q`�y�!��?^U��ԡ�^�6�I�(�4E3!�ŀS!��Q�`��e���!���r�P�c�&�Sv��*
���';��*Uo��\@p�S��r ;�'yrD�.��Z��8�A��t�8+�'a��"��&uU�-� �W'j4���'bl��R%	�O���j�L�5R����'��@�QkB�_�RQ��k?T��\i�'&��1�HE�Bܠ ��韶q1!�'�FL��؁}�Qd.f��<��'��a+q��<��M`���+L�(EH�'u.|��I®E5��j�n�2DOVq�'3��c�k�m�8a�2��$>�����'x����ɊH��9�T�H�CW�d[�'	0`�0�,Lф�ǔ'?��'�R�Ԯq��s�̸%-�'LP1Q��%%|
��r�� �-Y�'T�=P4�C}��Bc?�4��'��WH�"���X���.�0۵�$$���b�N�j�#%Wrd���)D�h"�X+>Љ�b߶\Xb��'*D�X%&���[RE� ������&D�� ��K�HKU���Y��]ti�"ONĳuFP9unRx��(�nsj�Jb"O��I0�p>s�O� ^���"O.�YwI�7*h@s'� bE��"OZ�[3$�<3�� �d�X���"Ox�F�Amʍ�abG��>��"O�`)�d��q��DD�n��B�"O>E�Ҏ��`�P6ڋ��D"O�EAb�˕a�ƴ ��U�JhP"O���aց:D4���
�W�Ҍ�"Of$S�G�1Otd�u��]-�yG�*R�TE
L��H§�y����~�����K�~ţGJ�y��\�*v��y�PI�fx�����(O�=�O��R�)�	r�F�z�	"q��1a�'�8�ғ�;^X��$���n�����'�X) g��q�J<��E7�T��	�'�R�eלL�~!'�H�	�'�δ�j3<:Hy�e)�
��� 
�'���[%�޻8n&T��	�65-��	�'	"�[�A�x�D����.?��,8�'�jTڠ�O�M��q�a�+$ �;�'u�!�C�Yg�VbsA.8��XC�'7���DY�t�������A�fP	�'�X� �E�XH�+B!9O�y����x��\y�A���E1�,���&*��O$#:�ߕD�pk�l�f�Hh�1mGf�<��o#�81N	<w�.�B�!�i�<���Ȱ5Mv����<�����d؞ؓ��|BN̟)�8 �Qs0"�{A�U�y���6���jZ�}��`F,�p>9L<��!��.��� m´bXTx��I�<ᷧQm&��1H6����uo{��Ms��hO�.���FF��O[hVB��!�ğ�5V���%۲YO�)�Tk�$�qOl�=%?!P�هF� BAL�^�hw�9D�d��S�=�"�+��!A�*D��
�J�DU�ԩ�c��v����Ah*D���C@M N�l����C5Pޠ0��m&D�<J���`|9��bT�
vh(0�� D��b��=37��h�a�?C�,�@(>D��SA*���`C� @�*1@&D�� �d
? ��1�mD�<�$D��B�_�Y��|H&��8|� �  D����W�f(��q��g��� ?D����#��a0)Ǿ{	�X�!D� ����?2shQҷB�S'�P���+D���q��!2U�����(��̚ �(D� ����XL,z�C�����@L,D�4��	J�f
:4�@dA?vp� +D��Y�٦��y����-���*D��蔧�ND}�DEڈ8�Ɯ�N>D��3���q�Q�4�=!Ҋ�rci6D��b�]$��` �&K �!�d4T�e:�,�v[���!��@����!"k�����z�#ܢv�!��BGbp��x���R!���!��G�yMĹH3�\�I���a�� �!�(|�ઊX�d(J"m��<�!���8*�	A�b���ا�z�!�D��bn�<q�>]B����yB��$?��bŞ.B�@��C�S��C䉱�� R�O��B2nD�+Q`"=q��T?)Z��0p�mK�l� )��[�e9D�� �ҡO�Ϛ܈#`T�Z�*A"O��p�1A|��ЀĔO���S"On%�&�H�+'�HA�8x���3�"O�4Z'�|���f��V��D"O���B��`��$�&���=��"O8�I�L��=�*������V�d�����-�S�'{	Lq3�8@�a Z0���Zh H. +?�F��G��G7�(��B�R����|����F?nځ��A��x�
��2D����8%zɄȓ] �(�D��1�1�F7�䝄����)qi���h�u��	)�<4��}�{�� |*"1!T	��Dg^���hO�>�2�((8W0�Պ_'�3��9D�|Y�j�QQ )�GDӄ�J�9D���稍�1?����UKf@*��1D����Ǘ�W���*�kv}X�o���y�l��R΅�v�y�4)ӆt����g30�Xq\&#VA"6�Ad1�ȓ\��� O��D���������.W����S������tW��vcʂnp��ʉ*-��ȓj�$�r��!i��Hs��.-G"U�����.����{&�/G�^��ȓ4���ʘI��*#�K�h�&��F{��4j�_�y�E`
��z�s��@#�yR(,-�@��$aĳd4)�gD�y���?+.��a�U�0i3)�%�y���, ��I\Z�i�/�����0>�&G��f�r8�&l�=h�Aee�<���JJ�4H�!_%��FFa�<���ɓ4�p)3Ą�aې�+��A^�<ar#F�w��lr`��v�~��N�O�<���<��j`�Q����I�yb�׻|^��+��w��Iq��1�y� ��dm�"��9@k�ѐB)E��y�E�7����.L�2["������y���	?� a��$"��S4eN�yb/ǒB��Hjw�1�rDq�ṇ�yϐ�A#PA�  ޗ$V�����y�o��QZ6̛D�o`E@��=�yr+�8yc2��ņȻb�����Ȓ��y�(F��e�c�J0`�4�K���+�y�	�B�4��N��^i~ubG�D�yRNF�`x(�"p��Z X@���y�͜�!�����O���*�n���yr/�E8Dٺ5�H�� ö�.�y��A)�0� j�8!F���
��yb
� 	#.�6	�H)�Kۊ�yBm��t�6"�k���~x�!W	�y��
l��)�p���д"�Ԗ�y�Q���6a1a P(��
�y W�Ló��D��+d�@��y��ق0�����7v ����yr�-zd(tM�-TZ�����yR'�+
ZY١�@��" �۞�y2�S(��(��֧~��Z2L��y���yj�3��E N$��9�OU(�y�3VxJ%��C�D<X��U��y���C�qugK�A6pp �)���yB���fh�g�2I�> Z��S��y£�����ȴmF*���rP'F��y`H���1(%I�8�H�Y�.˘�y2D�)LF��p�h3�8��	�'�y
� ��ɦ�޾��*���K̲�2�"O"�	�f~fRiH0W�+�hL�a"O
 ���D��Y�� ����""O1�b싌F�� �P!����	�"O����#TY��ٿN�i�!"Ob�r«��,����0m׽Ey���v"O��l,ni: 2 �R�JN�Q��"OBX����K֒���l�7o�H���"Oh爆%`�C�X�\�X�"O�l*�DL�n�ZPP�DG�@�Teu"O�i(�C��2m-[f��J0"OP�+C�=J@��A+��{F�0�"O��+ fۯf�P���͢?���"O݉R/��Pe(�"�W*"$)г"O�,95��
W���X�L�bq
�cp"O���D&y�E��+�mZ����"O�t�G%H�HdbЄ�	9)�1$"OH	{tᏁS���a$�[V��s"O\���CʵrPtS`^#go�$B�"O,᱂�����͹W��L\$���"OLa8��r�ȱ���T+.��%"O��6�Q42f�DY0�۟]�4B#"O�$�$Sy2��S-��sS"O�(�B�R�#���.a�Z�h%"Ox�2!F���HQ���S"O(�׍W��Z�莺o����"Or	2�AAsX�WC"/.�@�"Opx��.]�=7pm�rc>&}`�
�"Of�� # �DT�G�=Ad���V"O���� ͵KQ*U��`K
uR�0(�"O.�b@`Y� �Ѐ�B	��2uC�"OؕY�dÍ'3��h�cj6�)� "O���
��A�P��M *2���"O�I )�h>��1�	�r&���"O �S�ů�u�
�*�ҔRF"O|�"T�Q�|4��p���qǤ�8�"O���P� l����cƸ���"O(����+��5�fR�[��D"OS�n���h���KR�t<�(�p"OԪǉD�&�
�S�*ײN���"O،a'�T����Ȕ;l� P�"O�+p�_0�}�&(��<X��T"O�T�s˃�%<D{���-uZ�"OP��v�L&�
�b����mc�<�'"O�%`���w�I��O��EL$��E"O���dȭDM��S�xnL��"O��`��2��sh�#�.��v"O�"Q[��p�WVc�
q��"OftrB@٨>�I2ƆЪ�ht��"O*;��Q�XY2)��'E=�,��"O����Y z:��ʦ��w�
a�"O�!Q�!��A�/D�:��ջ�"O�y�RT]����Q��C�0��"O����7α�$ ��#�H0F"O��´�E15��Q�a	a�IW��y蘕�R[�!�L�>�@���y�hI�<|)�ի5zb�j�Ɗ��y2�c�ɑ�ԓ;�JyХG[�y&�}���� ��:#6`k��>�y��׊��H1��h;����c#�y�D�]�*H�&��0beL�24�H��yr+��0N���2)ߦ+���S��,�yCϭt{��vV�%��H ���y�,/z���h.�jY��C��y
� �%�5�M&|S�PyAj���X�"Ol�;��+fTD%p����D��"`�<���AY�$3�d-�Q�%�B�<�%��4@D̠a��#�F���
x�<�V!F V!��ԎU�.�>�� �Hp�<�֬�w��i�l:�����SW�<��M�D�P��׾}T�Hc4*�U�<A��)[T��% ˰E�y�@Vg�<�AƔ�PW��1��5�`�Kc�M�<����3k&���a'H��UM�<y�*]��� (w�U�ȴ��d͖N�<a��V��
��Յ K|iq%K�<�JR&p����� z��u�3��m�<�VTz�9��l��TnZ���o�<a6	?Opc����#�%{r�@j�<I j��� �c�63�̉�s,j�<�EE7`�P�r􉘰v1��{"��|�<��Myt65J���06�Ջ�K�]�<I3CW�~@>t���ͩ���sN�_�<�wl8��1����]C|d���_�<�u�<q�����!5�Zek��w�<�4h]5VJ�($�Ú1YN�����k�<I A�����!&���gnh�<ascK�i�4Cc�Y� �@�hDe�k�<
�=M�DPEN0ږ�{��Sb�<����lwf�3RMV+A 0���&PY�<�D&�e
�2�ܫ}�!��,�}�<aVKAq���`�'Z�p�J�GG}�<I��G�v�:��v$ŸV�B��x�<���i;��H�)
7o�A�#J�<I&ID8N��`e(	_dl�@�O�<�2c	�v��	JU�ɟ ���B���H�<����h�"�kς���FAEH�<I�B9�yanX;�ؼ*��C�<�S,\�4�4�Q�#`�����}�<�G�̵,|���#_��P#!��{�<1Sɒ�V���;�.#A�|�a�N8T���g�)PN����Щ)Qpԑ��6D�����8_p<5b�k�� p�m3D����Dg�8頧�S%Z�#�B-D����ȉ��6e������G�*D��S#c�%�� v(�+o�<�F�(D���a!M��"1X�E�����j)D��x�ע�$L����y�����'D�d��ϙd�T�UL��B�X�2�$D� ��f�)�E��B��H�!G D��:��²0�(�
���F펩i3D>D�D0'�܆"��BroɆ`&TuQ�)=D��p��42`rВ�I�7>\����;D���p%�;Of�-����C�f���,D���ϋ
i�zP��La,5�$)D�t�vM�\�(3��ʒ/14�q�.(D�����Ûw�hj��'u3`5K��:D� ��S�i�� gE�8D@�,7D�����-1!R����$J��@w�0D���Ь@�z�|���IR�\�XH1j$D�@��͋9i��A�t'O��xX��#D�|Q�W�stލATA̡����g<D�Xw*��E���[%�_�gf)c�&:D�����"���y%-��!A�Dp5�6D��J�Ʌ�R?ε�j�
y����5D�8� �J�F��x�A��8H����4D�Ђ4��K�n|	BiH�`����2D�8s,�v�D���ǀ0:"��Ӂ0D�� X�C" �, ������]�V� AJ�"ORY"�' AH�Ę��ɰ�f"Ov�I@D2<�X��F�84�<�p"O"Y8�	�7k]����8S�‘$"On�8��>J(9�K9uĈ�"OvL"��2'<�;�ܣVe��s�"O���_5Y�j��ʉ]�8{�"O���!��0o���J&��YA�"O��CG9O�T���
1^��q"ONрi�0>!�Jb�i�"O�(�6腺6��uЎ�)U ^詧"O�$����J? qYT��]��ˁ"O8l�«�a�=����2�"O��9�ꅱ �H�6Θ=�.�"O�!��8F�F�#̾l~�Ur"OX4J��].sgfE� ��(B|p�"O�bҎ�6q��ee"y�̑D"O"l��J�5\@T�EjV0�"��"O�H�d�j�r�iׂYӒ�Bv"O��{�F-j0���Ի�@q3"Ohi��B0#�8��� O}lm	�"OTQȄAJ?B����� g��3"O�g�?���jq���4Ov�"O��K�`�F�JQ� (��A�� Y2"O|�! m�0[8�̪�8e��X�"O.��@-o�h����u�1"��y�J��V��2n +!�HX�!I\��y"
�wX"lS��(*P��c��y���w�NUi��\���������yB�C�.9���<�^�1D��y� �p�����+|�<�vE�6�yR%Զ^�)�È	$x%Α��
��yr�X >��򐇑�d�b��c�U�yBi��f(�B'��N"���,��y� ^�C�`X;E�@�r\rp�p��)��c(QG���+�ƚ�M���ȓv��A�2�� a]$��N+S�%�ȓn⮠y�̓v��Բd+�?'(�h�ȓ{������'�is��;Դ�ȓY����!K�kRf=҅��5�|�ȓ˾-�q�ռ8�uJ�@�7x&�8�ȓb�$����xd26fI�Sp��]��Y�!�46�R��r$>:�� �� ��;CJ)p��������K���ȓN�be�Ba��k"
�����3*L5��F�r��P��+XNr@i0�
%�����~o�$���̕L�^���D����ȓcpq��I�+ ��U�HU<��ȓg�������@�t���H~�ɄȓI�p*Bꛃ\��թ�bҔRN�]��A�Pa�æ_f�\�)M��)�ȓk�2�Q�h{?��
��V=}�I������Ĉ�< � ��@�D�_�`��1�L����R��d2d"���Ņȓt~��h.��cy���)^�QG���sVa�UK�"KΡX`�Y����CZ�)"E��Os(��P��9����f�V�xp�G��и��R�.�n=�ȓkl�ƈ==t�ɤ	,�E���b4hBǉ��Riq�M�,���ȓb����683L���-#?J���l���s���fN!8�π3K%�ՇȓZZ�(�	0A��|1��ԩv�� ��B*�=�e%��~��#Ķ1��S�?  l��!^�bf��d���.*8a;�"Ol�Z�
�g��Ցb��D=�g"O������jјpx�`F#X=�mg"OP�3��ݾM�}��OWC	X	�!"OF�ׯ QZ�����Q�u��4�d"O�@��e��p|%����x�\%�a"O`9�G�UZ��
;����i�k�!�>BR�X�D"
�B�\ kt��c�!���%��M�q�(�i�Cζ!�!�D�?_o޼ �G��9�.��w���T�!�$
�]�Hh��Nus���'K)&p!�D�;G�r<�NU _\дyU���{^!��Y����i�rK�Ai�$3�!�l���}A*i�C�N/\?!�d�V�`E��ȪbΠ,�VS!�$R�|j�<R��ѭ� sL!�Ė�Y'�1X`���[����K�.�!��"�b3�	z��#��~�!��V�;���!��Y����w�C�=�!�3d�Q m�a�
I����@�!�Կ�h�ab��<���F��!��.��u�P?4�0݃�a߽�!�d�M|}�&
p� `G�T�;�!�d<M����Ȩ����A�ؓ@�!�d�6����"�_	�jU�/�Y!�dK�6�K�*�?�޵���S1G�!�K&	�Jܚ��O�%��B� =!�Yj�bY{��vj�堖�Y�!�d�H��7-�S��i��j�!�d:ި ��׊z����D�!��$ㄘ�]6D贋b��-1�!�D�#Hm��P.?l��@/h!�d���`���FV�	0�yRQ)�7L!򄕺K�  �D��>gy�T#�H18;!�DƕF��i�"ɿU�hM�&�Z�a:!򄀤$�>�؄�M�Bp�K�� 7�!�D������a_�0$ƅ�eD�t�!��;/��I���<Bf��f�r�!��Ė%&������}1�0� �Jp�!�dD&`�P�'��	|zX]
Tc�,�!��3��Pd�֡4Bl%�W�ӂ:\!�$Eg��9p3N��A�ҳKL!���:����J�,,T0�*i!�$��k�h�R�䓸�t� t��0\�!�d��=�Vd�#��
��,2�˱/�!�d��t���L�!$�4�G�#}$!��Ƞ���JԦh�,�+��ڏ_j!�[W�{7虦g�|��%`�.8M!�̡eD!��Μ�x�A�-�!��AD2q$�7W��u�d�ݕ!�!�6I� q��$Q�y�g��]�!�L�fA{��_�����eF+,�!�d�d��dz��9��ȣ�/�!�D_�Z^r�x@��<�	�#�J j�!�Q�m�0��(N2��`ZS�ϐ�!�Č52P��FL_)�d��aM�/Z!�Ğ%C�r�(��'w�@��� Dr!�V�(�P�*���H���dE#z�!�P�N�z�������8f�ך%�!�N#1�� �F^�]���� ��!�Dͤ~4��8U� (���(o�!�A�$0��K�F�a�A��<w!�$=,��k�"O�J4ʃ�؏5d!�Ӹ"Ʃ;`��ʝ� �O�!-!�� lY{�f�h[P�$�Ɠ^�@���"O┃B'�bJ�h��_�7�α �"O�	i���l���I���""O@)���
�+�.0'��_�\�@�"O�-z��˳b��|z'@��pŞ��"O,�BQ"N7�l�2���F[�d�"O����F�0Z���B��;B���"Ob|��a�/����E`(�$X�"O�Q!4b/!�Lʇ��-N�L�h�"O����*TY�H$�](=VT�"Oh`��vR�çܷ+�Vl�P"O�İ7�Ș+�j��OӐv��"O����:A^�`��/�*���"O���	�&����(�;Xb��ku"O���P��%�NlQ�RIt8@V"Ol���8�\i�e'�/~�#"O�	���Ł"�l�����?@��E"O��'F
i�hKcHA�0=�G"O\�!�-�"�:�(�(�qk�"O��s�������IɆE���"O����+ǋU���ʕ�.z��0��"O��*�Ʃ`�a��N F�b��"OQ���\�\��F(i���"O�h��dR-⴨5��
��$z�"O��ZF!�oz�"��E�DO�e3�"Oxe�XR�~ �c�M�NX�7"O�	���n���(�3 ��H�"Ol�q7CUDv�ђ�I����c"O:$�`�XE�w��R�:`��"O���O4d\<���U��ay "O�@�R��`�hDyQbҢbX�TY#"O�4���:M��X�Ǉ֭S'�m�0"O�=[�� BPV�3��.%&|��"O���削�r��@Z�i���s"OhX:7ㅬqzԒViI\\�I��"O�\
� P�w<��]".�`�"ODȓ���R��a�ڥX�"O����+&4������Y��D"O�mI��N�)����"x=L�(s"O$4r�:#����wg�0x%DU�"Ob��O;T#4��%����*q"O����6mF(��A�I"O�%�G$/p�H�J�/����d"O<��`fF�9��A�&��I8�Ĩ�"O}�@�I�*0*-���LLe��"Ò�͏�L9���q���m$\h�3"O�aYR�t$�d��F�����"OܽT��>+CpTі%ͯ�"�څ"OL�k�'L*J!�� Q'�Qs��;&"O%�Р�5�R9�']�2�2Tj@"O��z$蚈 Ĥ�� ^��1hP"OvxW"��[K��i��)�܌��"O�|R��\�K:1��≟E7�� t"O6mp�O˶VfPd�3!�)q�"O\�q����C�h#�ʦ{��=��"O��9�f�(��E0� D�"i��"O���w%�I�����@;�F	+P"O��v�/*g�,�`܆]�R�h�"O�	*������P7��*���"O��Ł��f뼹�aB��{�,�S�"Oh��-�3vwJ�K�P/g��y�"O(s퓅lQ�4��F�M�|��"O0�V�E p�\����M�P�W"OB���,�9U��{��^�4-� �"O� �EKW�]2�
�lĊZ�T�[�"O���Y"=�h��L����00�'~�7@ HN���"�Kg����'�mz�g˛���e�.1*�]i�'�޴�sL�c��I�Ͷ��}��'ft��t�
� ��aJ �������'X,��e@�?m�T����	74�'r5�U/��J��pr��q�y"�'�
` t�
A�ؓS�Ɔt���8�'@�� ��G�����]	�� ��'-����#Gi���)��!�'}��q�U,���A�!D���
�'%͡��ʷSi�H����l��P1	�' P	�W�*X���0J �"	�'�p`�q�Q7r�B5kݕWJb��	�'w"�Y� 1Q�@+�kׂO/�d��'���P�
��-!��'L���'� z"�(?��1e ��Q�'!�������P�5J#7?�r�'�PB��ԉ�@�U��)���'*�(�P$���d�	%C�vĵ��'�$�c���V�-sA�+^���'X���	�52p�Y���\D���'�x(����Д�ƉD��)P�'�LЀ6m֧y<:�Q���%��l@�'�J-�G�P�.Țc�P$��h	�'���q�U�_�)�"�^�i���Z	�'�x,a��ux���ľ\a̝B
�'�rHi�B�g hi��(�0d�B
�'�)"�C�{���p�aO�$kj8z�'��]9`�x"̪!Z+��|��'����Z5:��"�ĩ0Vj���'Nx�؆�O�z6�p�3�\Nz�	�'��ه'�13 LF�^�MNj�P�'��1����zW���-R�4�x���'�z�p��[�Z���uB�!]�X��'i�|ipnñ4~�Q�"[Q���'wl`��J�p,���e�OR����'�x�Z$�[�;HB�YU�]L��EB�'�4�3�ⅎ�"���Q8��P!�'s4Iq�kI���&L"�� $�d�<�%f�S�N�	�Ӝd�P�+U�Eb�<)�N�7��`(���/6�a Y�<��iݰop�a���
 R,JD��<���3v�d��g�uMJ|��S�<񷁎�^������n��@�bgAJ�<١�"���5eF����j���<Q��� "W�-�U`�Pٺ�n�C�<���c`��2�$F�����H�<��I�*v���ن��y���! n�Y�<����>D+�9�"	2$�6�Br@�U�<��aвs�^誷&˭GK�h�_T�<��±@�ڐ� ��-g�AB��JI�<��c�&N" Q��"%�Fb���k�<����0��� \:�z��c�<��B�A�J%��CX�Y�C"�j�<��>�8���1"��H�JZf�<�S�X��A�AQ�yi�hc-c�<�a@(��y4A��"�!��D�<� �[�)c��6aH�}:���@�<��.��x�j�SD�fh�~�<��̌�%9�PH���O��b�_F�<Q�Ɣ�"8��!R�[�F�A�(Fk�<q�J�"N��b����Y�$"j�<� �M� O˛km�`#4�Fuv���"O�<�pg F���"�#�&TFi��"OH����d�$p�O��,���"O��`�A�9�:%��H̨a��y�"O�l�� @�h
���[�|At�[�v:!�D��'��*@�s����T�{!�agD��=g\�A*��|!�DS�"�h�$�)� a"�=*s!�Ě�~Y�� ��������ON�g!�D0V,��u`��Ai6<ۃ�E+wS!�d��	�΍K��M~J���D.э)A!�H� }�����*��aqO�4N(!��ζ$�Zɋ1���������=r!�K/[H�q"��$4��e�Э$A!�䋾`g�8�sdD7ܔ
��$	^!���:/�m*� ���C ��>!�L�b��d��h�\Z4ó%��L!��!urP��B"ؐS<hA㭋\�!��.
��Y�A�[A
���MBH�!�׾_\dQ�.'$�l��f� �!�$̚ �%A�bԳP2,RV��!��$�P ��DiY��͑h�!��B�b.̣�g��l�56!�$
LP����4(�̬s�j�*a0!�.!:�	��ʗ}� ���$.!�$#CJ֕0F ��d�,D�u*�!�!�HH$.- E��ܢm� �E%HC!�D�p�*�xB,�
�T�L�`!�,Z�i0$2�R��Iܕ2�!��B?n��eZ�'ͻ[���4h��z�!��۲E�`rA�5�z쐁�g�!�$�.� � eN�<�1��+�!�d��^��!-�}M�`�W
=z!�d�)����(/�(�PDٕ
!�d�Dh�����T1�q���͔\�!�Dʺst�0qHA Z���ʹz|!�dW�lhx2��"�!�8q!��ƳP��{j�>���2A"ں#R!�dO'��`�D���3�`�AΨ|d!�~��t���6T�����,:!�W�C16��Ҥ>^����m ;fX!�d%��@a�;wCD��┟O!�̈́H�lj���~$�����U)J!�D��i�|̂�%Q�#l�����q
�'K��!�ΌD�<Ԑ	�! ���'_u#
5��:�*MB�$B�'%BD��L$ x��(�;#����'e�t�4͑�%Le(�̂oz	��'I$U����!1zމ�ꇳ�` j�')�)����YZ���D�  �	�'-��K�Ȍ@�Ey���,��S�'D�۴�G�@��]��B��m S�'<�l���ŜV���"����'R��:'��$d3S� 3
d��'u��T�ͩF~�1 @ǣG�s�'L�� ��]�mZ8�%D�<�XR
�'�pò�Z�i�|� �03[I�	�'�-��f�p�z�B�nJ1���K�'K��	٢i�is��O&�`�b�'~ ;�L��	�fj� _�$�'H�Fղ%�~���S=���	�'�ڧ|zr������i��'T���o�	Ps�CX	u�f�r�'�t��Z�h�p�����o��!��� Z���c�
�0i���! ��@0"O�C�NB�V~��[��#^�H��"O\X U��
B*D��N�=L�9�@"O��H�.@��-����:p���W"O���O����<��%�"OJ�@iK"],@�l��@�c�"O�4�����1
�5
��
��"O��	dʔ����Z4D�5z�,��u"O�$�1o����6��'�}�"Op�REG�J �R����L���2�"O�ءq��<�p���L�
Y��P�"OB!)��٥G�,y(@�ɩ)B�-�""O�9��!���]Yd�Z�l*n|3�"OnL�v���3�`\�VQPtd��"O��R��P�dY��h��Q�c�"Op���ٲqy�d�"j�;�0l�"O����o� �\�eI� �8Ae"O�ȩ��1~���(�.E-�|<��"OV���Δx�@� ���F����"O�r��: �����+0<]*��5D�L��C� G:̩�mؼN�pH8D��+��ɧcul���J�0������4D��s�[����
$���I3D����h�A���P%ţcl*�:ƭ1D�*C�+1����@�(	�qQj.D�8 E��JR�բW�^9u"y�1'2D�d�c�
0�6���JP�X������<D�(��g��]$��Qs�MQ7�2�7D�p�GH ���I̍�?�H���4D�|���W8d��<`��Ƙ/�4]��=D�����r��$
#�
�Z�ɂ�9D�8@B�����)t��k��;b�9D�� !+)�� �jU*b*P��N6D��	Go�6��}����%M�3b(6D�����I����fkT���A�1.4D����%�$��pB�� v�8��g`5D�\�%/L2�p4���+z~V�	%8D���ƍ;n7��/�Y�6�K��"D�L���)Q��j%f��MBvm%D�0x��"KP�3�E�O�)��!D�����Aݤ�� E�WDܰ��e D�aSd�M�.Īm�q׼�h	2D�� �hC>_.d;��T�d"�H��/D�ؑ�aT$Ut\*��1
_f@��J/D�����'t�iv��:xٺ�e2D�lP֍P*(���`�(p�p�6D�<�3�7���+ӎj�M��+&D������ y�j\��fR-�2#�O%D�@���E��i��d�b岰h�`#D�0��ύ�PS�*�J�'ض`ʱ&#D�P���9�ܴAG�k�|s5�!D�$�W�����3Qd�(: u{��!D�0���J*֊��G��w����b D���T��L���c��}�>ȫ�?D�8��
�qC4�����'�2�0�D<D�T�q�]0&�ve�փM�=��,���:D�\p����tZ -�a��y�����-7D�D�AF����M�p�e�$	iF�0D��y���Myཋ!��v	6UH�,D��j�͛N�����]�H-p1�	8D�,�� �6XȤ�ARd�z�J����;D���&a�"��lx�(� rMPU��$8D�\	�C�r����A
N2\���&K5D�;
`���,ʘ-�����2D�� ��E��nX�ٰř�V��p�"Ov���+�S�x��PʰQ@"O:TbG$A9���3J`1�S"O�� fB����P�ǎD*��z�"O^ipg����AqA��5���""O�!���rZ~`�$X�k9�tr�"O�����e
eCFzM���U"O���W��\6��bΕZ�t�
"Ox$	�/ֆ=faA4�E��6�z4"O���`G�:h��#�U�J`��"O(f�G;TV�&q-��3�)�N�<��J�
����r	B	"FJ�<���șh���&�K�=��h�D�<a3m�n��c��v�𐅢�U�<��	,(��,���ߧ�#�F�^A!���+G6	 ���?4����)L?q�!���%�`5ZǮ�rK`��BQ�!�K�J��H�"�mX��� 1�!����ȭ�1�\��@K����!�W��!F ��'fլpJD�"O.ղjJ !�`	��R,cRX�{�"O�$c �M�G��1���݀UpʜYS"O��f_304�aڑO'Jch�A"Oҍ�h+E�� �n��oGjA��"O�-Z���	�̤�`��!4�`a�"O�	�RoU<g�vd�ݞ|��"Od���˸
_�Ӂ�ņ;␹$"Oh�d�I�a��4�#�%E�Xr"O�%ekG>b���jeS�d	"O��3c3Y����L��jl��6"O��b����Sd�ҏLxx�"O̵�WEU4d�r����J�2Tb�"O��c�/\�yM�D8*

l�c�"O�ACR� ��q��KH�:�"OƵ���]�4���:����2)�"O41�FΪ~�.��f��h�\"b"O�H �E
�*�V�@"ĀV�ԡsE"O���R��!;��yxF�	�t�(�yR ������R���v陧�R��y� U<�ޑ�U��&�5��X��y���"z`�B`��L�A*�`��yB$������#Ѥ#2&e�����ybh9�\�c(p���Q	E�6��B��;a���ׇ
�v��ҡ�C�!:C�ɑh�
��R�8w:A�� VX}�C�I����ud������mS�.*�C䉩R)�8"GgUȴXY�Č*��C�I)5b`p��3{�A`�]�P��C��/_[)�FM��d�f��?L7�B�.M���� �7@L)�"(E�FHB�iK�����ҫ:x45c�	Y-�:B�I1Y�j]��nK2|�&�ۥd�!U�B�	�X Hw���IS��p���StC�	6�V���$�	TBDe����=.C�	�-��,[`d�3E"4��p��]��B䉣+�Tcg"��e����3VB�I�NX�ŦT:@�W����C�ɅM8����̒f )2h7n�HC�IM���!E�<dx��*f�U2r=lB��z�@dc��>��@��H��ԢB�
Nr��R��r=k���)�@C��!j��l�(G�.y�S�"O�=a�c��f�`�gM��i�Q*OfMp��G\��
�g�2v")���� ����)��O�4!�q
�4w�P�a3"O�	��Ьckn��g������"O 	��$]<�.���d<f˺5"O�p�ti�'k��� ��%�(�a"O(�R���@���=�<��"O$Aہ��I�I2'NF�cN�hj2"O�iCU-G��~,J�C+G&jM�R"O ��Q�IP����6�,KD�b"O��M9��؁�^	P��2"O��K���q�ir'!���"O���v�Ǘ$>�BCo�

�
�'*�zsm��WflA��<nY�	�'�<q��زPm���DӮz�:0r
�'0T`��b��1�|����
�,�*
�'[�]��蕣7)@Q��TB��'T5�w#S�6�=AfG?���8	�':�Lӄ,�%�mE��<��ȡ�'<8@I0 :0o�1CD�<�`�S�'|�� �S�J�{�@�1�@��
�'���v��v�6��f�H�,6�� 
�')Z�C.��0y�PzF�>}�T��'b	�C(ð3$��څ��[�4���'!���Á<+�A��	#���Y
�'�0E�V�@nΝ`�疹)`�D��'̢\`s��Ӽ�;����"|f%I�'>���,�E��	]/d��Q�'p�)A�D&��5KUĨPk�'$��$BM/'��#�Y�7N��'v��j%`B�w��2ů�0}���R	�'<��a�(���
�/H�����'j��ca��b1�2'ӿ;VJ���'�P�`�[-e�\1�"��,7j.���'��U+w�J�A	쨀��<.�����'�0� 1'қ�F@�C��v�<��'���e&H�>4�$ءn_�q��)��'�&�U�C���]"a��gۄ	��'s@ 3�M�RӖ� ς6d.�l��'�pA��_"F�53��XF��a�'' `�r.�#ў�P1�ߩ<�\s�'�~�SB�(Y�L}k��8�(�'W�=XWK�"G����.b�ma	�'��i!��<-��;զ�.#��<��'gh�FM�"�l�Ԉ�2N�`�'��r� [?"1еS �тg�y��_I{��"AT�9�|�8� �y��)j�@@5(-,3�0���yBkH�!�>��v䐩p�٤HX+�y�K��nD;�ő�x�q{����yGX�x�F]�r��3�6L1�n_�y���,�0	���H�B%e1�k
��y��4 q�:C���E����o���y���}'���鞢9�$����y��0yb��Aa�/7
��#�]��y�e��5HcuJĐ/���-���yr���f�R�ȃ6p7|<�
P��y�eO�e�6���.f��I"�ς��y�ıv(,��^5ds�|�s�D	�y��T�65�����G*c劄�"�K��yr��m*�E!T��.N̠ H�j2�y"�I� U�(�99&��R���yR�=�l�I�I#1�^젥d�y"�ٳAqX���H�+袰��eߤ�y��X�Od����u8�]X�)��yr)Ŋ6����տW� ࣐!^��y
� ^p�v烂i�p�DU��1�C"O��q��n�P9�H\7u�f��7"O +���-	K����.X�"�$| �"OV��쟻_�6���	r��郂"O�u����$�bP����G"d䲕"O�Չ#��<{��,@m�1�"O�X�,˛4���q�!Ώ_	���"O��Z �P�� `�("��p"O�����̓:���h�1�`�7"O��r�H(��4v�F�97"O���r��:����B
�\�a�"O֑���V����V�Sࠀ�"O� �e Uy
uraE��t'�b�"O��"�7O��Tt�D)i�=K�"O���j
Pe:�`DBȟ��0�"O���F��AkV@%l�!{s"O<��wo�x�>d��	Y֍��"Oj�����*��X�1�T�B�n��&"O����.�� �����a�5X��8��"O� +#� @�f�ȓ���p�j�	p"O1RǞ�S���ᵤ�4k���I6"OȜ��B�A���آ$�8U���`"OY��L!M��IZc��1�jQ8V"O�q�"'G�
!��ӓ$�P�8�f"OZ� M�<�zih�I�"|�P�"O�D�w�M��U	��@�#AlYs�"OQdbI�읱(N�`"���"O���	�`�t��gƋ�r\��"OvɁe㇓o� 0a��*�Q"3"O�Q'l�2&��✱e�U� "O2��G�>�@G��<6���+�"O�d�cV��<*R�L�=�Q*�"O�l�#
�K*Έ���(ˎ��"O�x8mE�gֆ�0�%\�Q�B��"O�a���	�шhq��0�dIC�"O,a���V�Dӊ%�q&$�bYq"O�D���J!f٢�8��S=Ec��"O�h����pR�#�h����"O��0�	��j�Y�BùF�T��"O�*5�޶f�J�0aG�3���x�"O$�CP��$bP�(i���q�"O6��Æ��x�0�O�q��`�"O�i0G*��0��̭::��"O�]�� �f�@��=�
���"O�T�����B�T�*�팁�jIiW"O~-R�䉶fK����5bv��`�"O$� bwe$�j(X�.Ө6F%D��("ϵJM(�ӧ�ڹ-3��1��"D��a��- �)3��E�G�©�TD-D�y���aIz6Ə-UN�e�*-D�x)@�B�2�]y�	��$���"��?D��s�$��]@�k�)�F$�{�m<D���'�_�/����F(pp�ixAL%D� ����s�fty��W�Akl-�r"D�[$��zdQq-�8JLNm���:D��a h��%Ў�p�B�;�!�d�<a�"p��^-`m��q�I�H�!���nCV��4�^�p_��J�h4!�$7	���薑X�z�k�&B�E!�$̪q�8}��L?=P���6�-L!��I�t4�􅂦*0LRqG=K2!�DRyϠh[v(Ũ^N��b��6!��*i�,)(��D�s��D�Ch�h�!��2*�J�b�J5�XF��2!�� ����R�8�>8�(E�]����"OP��,�(L+ɔ�G:`�0�"O���m��a�Ƙ"�O1-z8q"Of왐H1t�z�`@-v����"O<\�G���3n�R�<	����"O����âp�a�Ӂ�>.~2ت"OX(� ���횤�9`u�51#"O���	�HЖh�Cl�RX�ds�"O�����
�u(l�wʚ�EO�)8�"O���4cI��>��hϿ&5!K"OX`�nS]j��Q
͚�%���y�A	�0B�hЏD#Z԰Y�S�0�y�l�!R��iІY�]Y��G��yҨ�U��P����T'�XJ��
��yBH\3��t����M.�q�
�8�y�L��ub&�j�.W:c|]��E%�y�lҁ!3ʱi��_�.S�u�����yb��6 ���T�;*�̘��o�<)3n� �P4�R��{AD���E�J�<�䧗#��`�%$��0��H�<q��m ����yxT*��]�<7 K\
��� d�!fpiU�\�<1�^�]�p���ÎLـգUF�~�<Y�-C8܁h�@��T#�1)�m�z�<�TN��.��TIE%�	Q�ܭ�vcZa�<A�GQ�;�f�A��~n0�R��^�<!@	5H΂ �7���u!��Ҕ�Y�<A��ځdz0򆣉8l�$!���V�<�GF#K�樫Dg8N������N�<�`gS s,�p˾f��|x��q�<'aU~ސ�3 '�MF<���p�<I�oQ�q6b�S�A	�RC�:��\p�<�Ζ+M!���4$CXv����p�<� �P�du��;q�U�}ԙH'-\s�<	�߽�Mʖ����|��.r�<�A�>�ݓv���,�5�!�m�<��/�>V�0�ؘ��=R3cT�<Q�V�8�V� 0�=H���RC�I�43�����#��8���=6�@C�I� ��lX�I��(ÎE:r�ŉosC�I(K���x��Ć�b�`�BC�I�3�|J��)@4���g�~V�B䉕M�x�2b�ֿ{6��Rf\�Q�B䉉#��P�X�2�N�T���t0�C�ɿEȾ�c�
T�8�nj�!�4"hB�I�Ӷ��&��E�.�*`!I:�C��	R�ʍ����8��W��T�zC�I�r �z�ēh�$���#�V��B�Ir� +2��-%�)�W��,٬C�l�\��g����&PQ�,��J�rC�ɄTc�pK�bG*�2tkI$88�B�	�{��b EM��#P�R�?�|B�	
\+��h"E�/�M�$�4R}HB��;L��U�Q�����¡ЫX�(B�	�	I(��b�G�����SeR�B�	(d�ΔqvH�/�T#т]�L{�B�	�D�Ԣj��Y��$�2�[�cʢB��3<���x4)��#N�9 Ӥِ3IRC䉝��͹�� #Y���!�EUxB��4b�4��J� 	r�Y`���S�zC��4����o�\��k�M�>C䉃<|m��+=f"8���Jז5�LB�ɂMG���$���܉y�B6ts.B�#0=����u4��eҚf��C�)� �� �pk4�� _�$� "O*��"��׮��˰K�Z��"O���B� ��Rk9�� �"O���.��SL�Rg�PZ�nĘ�"O�%(�j�����	����c�"O>eA�`O��`�
W��o��X�S"O��hFC�;Q䠭�A��M]H]�"O\��E���;�6�H�F����R"O�q7�X�:ކ!�R+ך.ؾ!Pp"O��!�M^�>$���ɨ��c�n�<1�CQ�KݐIQB*�#yU�T�vgMh�<9���]�ū ��"R[��q��f�<c ¿ޅՐvO���`Ö��@�ȓ|��A�GΔ'<�\#���DR\��@*(�	�Ï	_Ci
�X�BT�ȓ
R(es�L�;9E�A�3Z�*ф�w�FHƧ
֞�y�A��.���ȓl䶍�֏½y�j$��l׮�Du���HZ3����dK7'��&��m��[���IT���X3$�O�|Ŕ=��59���w�D;���j�Dۘ�� ��Bt�qᰣ�(!�ఢ�OT��e�ȓT��lPq.P�]"Uj�@�keZm�ȓ>~:Љ6`J�R�ƴ���7g�8��ȓ`y�)x��[�32B!��04���ȓi�@���B�):����K�+]$<��O�P��V�z�p�R�e:����&��h#F31�=XUFѯ	[ʩ�ȓ@�@�&�
T���+E���F5�م��
=Ȕ#D"�!���O�vв��p��Y�MN<���Q�L�.܆ȓ<��*�I�+7btP ��8��T��n��a/�:?�xY;��	�U�ȓd�(�z���6�Z\�FM~V���ȓD����-O(�zs��8r���Rb������s�h�NP�V\�!��_d���Û�u��
FK40qj}�ȓ X��@�C�Y*�h3����;�<��u^6%ˑ�Q84���N�dć�=�%;�A�
<���#V�j���)/��y�(`��ųS��X<h�ȓs���S�D�p��S�Ď$>t��ȓ}��yЃ֦e.:��ׇ�w7��ȓ��HtJ�49蘻�+�=�1�ȓ4�H`QQ�,�{���P�Մ�$�Z8�T��U�\���C[𨡄ȓ^{~��	^N,Ra�ـ4%����N������B�9�c�4,�Ʌ�phR����m��T#
�l���ȓhC* H�掤3u08A�E�/�N��jα�G�<=�$D`OýP��ȓ�Ջ�#C%N�M�Vʕ�|b��ȓAu�0٠�?t(	 ���n���J�|�� Ro�t��ağ��=�ȓQ�@��啷���&��#Z�Z�ȓ]��c�b^�|.��	�\�Li�ȓ?zX��� �HĹ��N�� ��djA�*��h�V&�������Ĭ;�NdkЄ�3�\�S(2��EL���Ŝ���+Ud�z��ȓk<�) �Ҟ�dE3�U�*��(��5_��C�-e9��x B\a�'�~����:b�*�1sk�i$�Us�')�Q�;�P�8�/I?w��9���  1;r @F�Ts�р/�.]q"OZ=Z�EٗN��qH@��5vu�a�A"O�K��<^�<ݹw���D��
A"O<�kde^�uD�����6)�#�"O��`'h� \�=`���4�ٗ"Ov��	!���G [��ͻQ"O֤�!i�P�uo��E����"O�*�K�72������B=UҰ S�"O��q�˄E�ڴ�E�]�:��a"O����J� ^��"S��$x�ʸpD"Onţ0�/y��Bd�_�@B��A�"O,9`c�Z&�ē�h��i$ҭA�"O|��r�)c]�XH�����&
F"O��qш�9$�i8�Y�x�B�c"O�ɩ��3��}kRS�U�
)c�"O��[�.�Ĉ�`�
2l�{"OP$��
�0 t�×�
(����"Oh���N_�=Ѿ���VE�H9���I]}��	�,W�IT�DB�c煕K!�d�$���yc�
:��m��Ƙ=T=!�V�8��@�� �r��86��%�!��Z����f�#x��J��,�!�AE�@��G�j�ؔ $�1:�B>O��r�動,~h�X��?1GιP@"O�y�M�gF�1��\�-�����"O��c�Őq�X!�.�ؘw"O=ðk�=� �g�ؽ��zg�7D�@��4Xd�ydo3Zq�!d5D��P4��9�$��	�O7�X ��4D�\�DgN�~|�1L\�Q�M�5/�O���6+"|�._&(�����i�
�C�ɮ�Z�sS��nt�)��J�*J�:�=��O@�?=9A�?�.1�O��,��"G`!D�P�r����|饇��𭋶/���D{��	E�k�P��ׯ0���k��;/�!���bn���b���Fܚ�#̡�1O���Ā4]M�%��Ɵ�����z!�ߨncFa�7YhV�$	f̞+`!��{�i���C�dL��2p���S'!���&S�D���X������Q� �!���(ML�9ĤϚv(RC��`G�OH�鉞!6͂a �Y��j"GF&�4B�I������k�,27V=���	�P��O��eaxb�ʞ\rX4	��c�,-�VL���'�铘h�l����!G0Ej� B�Q��A��ڼ�Px�ޮ4�Z�%�I�yu����-�'��>�IB�I�,�r��@���r��ց/�pC�Ir�R��!��	Ѭ�oT.!�51cM��!_��|B��(���)��͝�Ō�B��""O82���R戸!�
S�9�f�[�	tx����$93�dhɢBC����"2�e���>ͧ��Iӯ���s`�C����-P�B�I�E����7k)M$]��o�%x��K�{�3O�44ONb� �ŭ\�s��[Ҫ�&/(pB��hX�إOB���,��U;�&��&󆽲S�O|��� QU�%녪�)��5��c�R.�$�O��|�C�7Ɋ9��eUI3�� F�<�W�H�T>�lప'#<�8h�n^�x�ў"~�I'aP�@9G�Y�$��UH18q�B�I*�z<I�A�g�0Is��� "0p��z؟������L�����;2��} ��5D�� �
ԩc�$����+���J6
7D��s��C"IAT��1��9�n�Ôh/D�̛f��!�ܐ	�Oݤf�jK��-D�� ��P�s���MI�F�N�w"O�� l�hM�qJao˲N���7"O����A@���Q�m	}KF��"O�yH�IP����f
� ��!t"O,fꀣ�JM� �'Ό��"O�\��h�$@�IT�۽/F�0�"O�l*���7y�4�a�������'�v�q�ˠs�@��5'%�$��'���g�ՎDZ�!Hҹ��]��'��[@�`�,������Vd#�O���dƥ2D.����Y�-����т�cx!���:	nT(aÝ<f�����	g1O�7M8��u"�h�0z���E�X+%� ��ȓZ�r�4�I��2��aҝ ������tBөF= �R���*[t<��L���@DK�e��!��jLL���-O�	�WG�%(���c��> R����S�Tx�F�FiIA
�;Q�Ɯ��b�u�$��<>~����8	ɦt'��G{���$�!Fny�ϛ|�~�A��߰<��I��3���aP�i�u)�
���	����3ra@9:Q�	ò ��O��=�~j�'ӟs &�!��G�dLThsǕQ�<���ڰ�y��I�'L���6��sx��Dx��վ�|��(��^�Q�a���yRE�/v�H0�G����8-iq㗖�y"(�
�&���	�!B���G���y�ǚ0�V�A�`��
�@���.�(O���DW#R�D��ԏL0�{�@�6lazR^���'C���@�
^��h��"OA�p
�'��qp"O S�P��e�98x$"J�(q����%#@���ez|D�5e�
@?!�dA�zy�x��&f�X�ѪA�;91Od�=�|z��J'6Z6�`��w�X��6�c�<�V�"j�5J�k�D�Me~�o#�O¥P�O����kWCY.ZL����O�S��̙>��lCP �"��mr+D��Q�[��. �A/D�y��xr�*D�p%��t�qˀ��
���ٵ�%D�P"G�� �Ve����9�b�1�d(�S�'G��e+@)ˆ9��	�')įJ�(}��M��D1f7���V.M:a�<���ϗO�<a"��;Iܼ�:Y؊��0�Gf�'[�hͧk~h����]��D�ξ��@ng(<ɳ�C3^Ёa`̸Nʌ`@$��<��tG��㕂{tzxIc �7�$9�Ȟ�ybeK	ssbmY7!ƕ0prd�߷�?)���9FC���"K�O�p(r�B�,v,݄���i��g֣_Ub4(т��c�Hф�u��͢�M�sΐ,����-w��`��G�T!'c�0B�Dl[����ȓ-Τ$Ŗ����ڴ��8����ȓo<M����^�:�b���[J����p\��	���k�����.�L�ȓ.X�,��R��Y���2`&"�D��S�,~�3 .�P:P�;[�a�$B��#T�6�*0�r`U���� �T⟴$��:��)�#	i�� ��tc�)!�$$'R|�N�%M���vI�3'1O���z�X�"J�4� ��+b������H�<y��P%M��`2 \���Aۆ��Dܓ�hO�O�P��!�0��@a�1�4���'�>}�W-M4����"$�M�tя�$Y�0<��f�5����2��Tӭ�E�<� ҄rp	@9t�:@�Aꆷ ބs&"O�e��S�$}<Px�[�2e"��7"Oj��,Q�! Vd9y\�p!"O���S-�<W}P�P6�õ\>"`��"O܅:���j$����` �~X ��'VQ�X��X�P��b��ۻ$��l�Fl7�	K��[��_1Ƃ�� �د��<qq�5D� ��F)-C�8�gW�{G����i3D��`�˹3v�co�	�J��-6D���"���"�(p��-�+'ҕ�T�5D���Tga؅�2�K/mg� �(D�9����f�2}�� I�&� ��(D�t�$g�t���`ȂI#�9�`�$D�|�@��^��'H��P1�)�j#D��y�ID<O�¼�/,���G�#D���6�&B:�펟��-!Ac D�ڒ��+D�i�$%M�3��i�f;D��sǡ�
) j���K�[�vQ���3D�`x��+A�YPi�KQ!��d0D��(��FT�;�a�mJx���9D�,q�D_�8���mD	K�P��wj2D��h秛L�>��u�a^���#D��R�K��5 �Ɔ�P���+<D��xV�ȧ:�Sq��Ws(-��9D���B�b���(�M�T�pr#A5D�xC�*4-�s��E�4���6G4D�4x��[?Mb��M�m]���-5D��Cs-��\9z���zX��1�i3D�4Z`	�H$� �p�P�:�t#�;D�,)Э	/(4I���>	�0s&�6D�X ���52�"��f̗("�ȂŠ4D�ȨҪL.��!�n�#%� kf�2D��:v�'QZ���Q1l��`��>D���sg@<����.7���wK"D��hbC̔5T�zA��)l�� �(?D����#z��)g���'�>Ṅ�'D��*%�� ��m b �,����H*D��ԁ�$'�hi��f�10�⭺f>D��S�� !��d��N(��q�a D���F�qRD�1���^=t�B))D��6Κ�]���G�jՀYH�'D��	��K�~B����Z3+Xh�% D�$�`DS?+E���DF �*����<D���q��'J��d�%.Qe7� ���6D��B���=(2���ō7q:��/D���C�АT�R���O��Q���R��.D�P��ꖫH Z�0T��21�ȘI�/D��x$�	���A�͆6EZ� *D�2D�����٢9��Z'E��!��TAwe0D� cU�X�E��ە�C69'|l1i9D����@P���y@�*@6/�J�*%�8D�yVj�-	�<�G��%�ba8�g6D��8�	l��q	 �ʚ4*y��e0D�d	p&.BΒ0䊝5R���-D��zd痂$�����͕M��!��+D��j�K��`*}C�jˁٶ�!$�+D���PB�sz��Â�0Dv�zv#(D�`r���=G��i�$ĢZ�~��&-)D��%%P�
0$�dM�Os�w,+D��B\0
hp�P�
�~X@ۦB(D��B�J�Q#��:��
0TŚI�6�:D�|��U5Yj��A@.��<�2e`8D��Cd� �\ى�2[��r�5D�(b�I@�4��1wǙ�0�$HcP�4D�� ��:%D��#�́�4�_%�R "O�0q7ɃY��0�I��*%�w"O،�2�G3B����運�z���"On� �Y����	�6�XT"Ohɀ@=Qr���1���p��L�4"O&m ��3jqa��7.}d�""O�YF��6�.�0сR.3p��s�"OV�yG�R�Tf<(�͉ ^�	�"O8]�T��9� d)��U'[s�a�"O.�i�n^�i�� !\�`�9�"Ob���_?<�c�n�c��v"O�q���L:+�0x{�-ʔvsO�y��*[l\�6�ق\X���k���y��FJ��M��F"I^�LY��t��ȓ+L���키ܑ��;_՘��ȓb�p�@c��S�Y�E���%�<��n0ԼZ&�X�~#�!v斠l���ȓ<�$��hƱE��XæԜ2����T�&Mh'`��YI�q�î5��$���A"7,S*eT�Ř�$֠R���ȓ7�� ��s`l��OV�0$<ņ�^kfM����=����֊K�vQ��u�H��F�Fr��`��P�Ґx�ȓ`iPe�e�Q�ڬ��hJН��sl����"J�c�����'��IZ��:c>�Y �-s�|u34b�8	8��6i*D�|����E)���$KW<i�0%	��=D�ȸ��A./�I��C(a74���,!D�LY���y�0U��c/�R�N+�]��D�@�O�T�8��{\�9��*D�����_�~��t��BP�`o��!Â$?��R�h�#Uv��l@�C�(�P�G2��&Z,px�L� ]Խ�ХN��!� r��	V(��IK�<Z7���xqў����6 e����m��?B� lL.d�B�	<�JhJ;!=01�%BB�7Y��B�	?v ��2��h�jC�ɟ~�hx�u�8���Ҫ��V8JC�E�#B�������}P�C��"����&= j���j*�C�	j�J�hP:vA��c��1w����D{J~:�ܫq��-�6[��j�r�<1����,��3��֘HWhGg�y�<�-֤O:�1�kG/-��!�z�<��# �R\��P	�i�_B�<1�+
3]�D�O�=:�j�p��Y~�<Q�*���	q�Hն̐T�'��c�<ђ��WW�Y����2\fm�WŊd�'Vb��8k�Y3O�+~�,Ԓ'�.y��C䉌k�vl�5オ_�`E�4J׻S B��+"N�I��˖�N%���ں=�B�ɹk풤;�.E0k���!۔(@�C䉶=n�A�Q�C��q�����D=�I	Q8!r����fa*���|�	x���0'n�̗:-������g1Od$ډ���c�ӡ&�9�"k��V�&!��Q�*�C䉗�,�{��H*[f(�`@!L,8`#=��m�OV��;3�>,x�A´cw ����5LO�� ö��{w�����ʁ9�P�7���M��7�矰{'f�F��i���'J>R�@(�Ƀ�HO1���1ф
�U�](�l�)0�P���"O�,��Fô!�z��k��i��8�"O�1*T�H�@D��VT��"O������#r��mʰzK2�H��i��� �d�4�Y�",
%3��pli��']&�D�y�L�6!Of�89 �7-(!�$�$2�tE��$8J�\٢ o���@D���<m@0��䒔 �h���4�yr�"J�L��G��f��5�Ҿ�y�`B<Mt4 3�/A�*��DbeE���y"�¢E�NaxT��"�H�Tc���y�=| @|��K����4z�_"�y���}���Ӗ��.UX�]��˖4�y҈��(߰I�%a�v��iB#��y"�:AfT�a�	pw �Q%%���y�B��aa|9@#�K*<]��p)�6�y��/S���5��1���%�G��y2�M�JV��5�ϸ<��Q�$���y�bY.q���	����2�ް2�7�y�O^�
�ެi���+S��%�5�y����̍�J�3Q).`{��R��y�BF<�6�Z���W�Uڴꖼ�y�"�b�n���.vy�`s���~|�_�b>˓�L��f/�1?�`�3pj�a|TĆȓ+�`A��*W:�	�U<B� ���B�+���O�x'�:o��� RFYP�OT�*�����U�TOF��>�דMepU�h��{��他��pd���=f�y�f3H\�-��K͌UV�X��sd)�5F4C(�]z��?z.TX�?1ӓO�������PU�	��.�u�y��?�FޜM"��H�[�N0�
Al�<�`��$B?�Q���N�`(E V �d�<���G�da���6�ǐs6J5H���`�<1�$f�9h�-QI� ��ZU�IX���O��U����/���p&�9}6��	�'���#�g}V��*ܮ{Q֝j	�'�@M�ꓤ,Q�YG�I7ml���'tq7�Թ�V<�v�"V�8 ��'�}BGA:�r4!����'0�9�g�±?��X����jHI
�'����>	RxI�I��B�h�B�' d){b�ɡp`�SL�9�~�j	�'<��SgDY�R��9�a�-},p 	�'���bM0��1�ݟ1�~���'0Pܑc���@��N�(����'� �
0�9[�)�p��:�k�'^��#E�-f��`�ɟ�]6�xO>Q��3lOh�$� Zph`5,���5
O�6�Obzy���2H�~X(# �JK!���&��y��ď!� �Qt�C�|���4�S�OY��h�N�b>(e{�!߀� �Z�'bF�2���+�UAS��@���H�lG{��o�*^a��B㏦4FjA�bǋ�yR��e��)�D
ج(�D	�KY	�y2"Z�m���	q�ĬR�ʎ��y� фD��`�#�Ea
8#����y���/aO8L�@��+�|�Y�B�#��O"���>s����镬D�H�XW�<Q/����3��0.�xXB
_V�<	-Q�'ټ%34E.<2���,Q�<q�G������o�(�"���L�<���3f�>���l�
#Gc�<���Z6Ht��bbKV�I���.b�<ǎ^%A�j�b�$S�v�)zW�_�<�fn�wN��ʵ��qbv���CB�<Y��^R*��΃e��i����w�<�C`�1Th>|��-�=i�2IڂMt�<� >��M�VX����`��s����"O�̘���"�I��!��m���g"Oj���B�;&�@Q�̼[��:�"OT��RmQ|q��qf��\  D�"OB��ԋ��4"��B�m��-Q�"Ob,�D�G	�z%�6*dt*�"OD���C�m؎���K�*"O�x�5i��ʩXp�>;���zA�O���Ăep����^�t4H�N�=�!򄂡_;!����;-�t̋�!�,Q����֫��W�2KҺ?�!�do
�Iؤ�V�>qS�Z�W!�dC�q�T=I3$�#�BM�㌩	L!�d�%|y�0��4������"�!�D��!O"�bf`��h��Ӓ�Z�Rz!��-O	�<�"f��S�@�H�cM=@h!��?[Ed�����/I�̌س"T�<!�$���FP��h͏B�"L��^8!�dS'w�<:PG&l�6�1/\� !��"{�XxyT���|����%i!�D�6+L�� ��B�u�K�"7h!��ud��C�I(=>�0�@? !�$ �\\��W�ǭw!��6�H�!�dیY���@��� 9lȃ���F�!�$D�7�*Aa���X[T,f�`�!���q� ���V�h �bE.�!�D�$a5���F�$7� �@�p�!�]�(�Tg�?7�� T@C%!��ʧ��4b�)P�,	+�ٕ
5��MEƑR1��G���f
͕�yr�ߔ`��l�慑;9�^Mau�5�yrmO�a��d��+V��dGU%�yd��Z���ӠLH�/< artEG��y�a�ހ-�Ǆ�U' %�����yr�\8�THs�&��6�%�4�6�y���+�Pd��a�2|��}�A�I��y���4�f�1�F� ���뵋E=�y�m�\��<k�.�,WD4ؕ�	�y�#���u���؈W|:�(5���y2��:�l-7��N���% ϛ�yr����v��mY!I8��2�N�=�yRC�7W�\�XկX�A,=ؓ�ݰ�y��żw�a@J33�V}1�`.�y���$��l[�E��=�iAD���y��Q�<��Ф�gU��Pd%�5�y��C�=-J�6��6��T!��yR$ �=A�%�wk�Y�"Q�I��yҤ��=�@2���.Y��%�r���yRCݓ0*X����K3�0*��
;�y�[#5en\�l��J�@1A�Q�yr�Z|��M�tj�EP����J,��)���'!�AR��?!�DP�*׾v�h	�'y��#� ��
�tm��f��{8�h�'��I�)neՂu��<qC����'�"yu''P򂭲eŐ&q����'7���Paػmrt�&�,�RIA�'��H�TC-^�,�g���,�}��'��a@G�8L�P�I-J<IZ�'�j�ca��+H8�f�#���S�'��(U+�,S`LL�v�رL� �'ޒ�C� ����UA@��~��'G,���- �Be�=	�/F -Y
�'��\��#�(k�P�)�l {��A	�'z ��$�ʕK�5� �K�,D"��� ���v���H�r	8�
�E?H��"O�-�1e��R��q�I �S(�Av"O4��E^�]@)p�܄5H�c"O�)CwJI,^��d�����b�ƑҒ"O\A�bn��4�l�2/��N��I�"O��ac�Z��J	���w���"O��Q"Gɿ}v<�F�£N���E"OB%r���7-}�9Y7��IȾ�ʁ"O�@�+T;gqX��C�y��Y�"O2�a�#� h�"H�p�	%��E��"O(���T�7��Xj
X�eW�1k�"OdI�R�N�X������K �z`�"O�dx䫘"UL�1b7i��0���"O�؛��܂,,�x�f)�����"Op!���[��Ԋ7O�x(#"O��q�G�<P��3�0���t"O&�"�!K_��* �Ϊh� %01"O����c�8�𡹤��b��u�"O����|����CMS��8X�"O������������7fLl�%�I$N�ǠOT�'n��v�H�L��T�V6���ȓnu
��b��^S�MR��A�&�>1�������R��ҧh�j��daڗrF6�(�)�{Pz�� "O�\AB���)�&fg��I,�P�<�t$�c�,�HS �\���ی8�HYS��&km,Ba�њ	c�}r��e�Ѱ3kK,)�����AbN��q�׬B�ܺ"`�x؟�g	�`�^���Ĳ!B�%���Az�$.S��j�'�ٺ>�&T�C�˓|�"�J'E!�D�+7�`��?�����B�&��F�?�4�'�U><�T�sǤ#��=+֭B6l��aǒZ��`�4D���5�Жr����(xı�C�^�r��2�2��B�ݹ=�`�g}£Kv��8����,B�8G���y�עޛ�����'mp�"A�+�52qdh����a�5p7��	B�GC,���`�<�7g�
�`r�k���A,�'Т3�ռc$`Ŋ��L�g&�#=!�/�p��!�_3�h��J?�у�[6L��Q�1�ɲY�f}�@�O�<۴u��$p�$��Mַ	f��|�'xiY��"V�"cƇH"j��4,(>�dj£wMr�p�-#ܑ?7K�+p��2��~�؁a��F��؁b�*7D�w.DeL�{t+�D^L�I�/4h
�@{ȒkԾ�b���O0L�ƠK�B�:5��[j��'�=D�6o�m�gX������M<���p L#2�e�QI�o��T(P� ��4O�m� dh� HZNH�2G(4!�d�IF��bbB6}���ax��j��R,���wOE��hO�,T��%��`�D��ħjf�X�Q���C���ѹ,p4�?�E��0|zv��68�8�a�[�&���V�Y�<q��˲p�YBϑ����6�����vռ葁 ںs'p� �1��@��~2��/ ���#����!`ɑƢ��W�6ɎP�u��|�Z�g�'�µ��o1����ƨ���RJj��&�'.����\DL���L:�����ô� �U�'R���A�<a7�M�"f�ʣZQ�`��Ɔz�9�H^��lA*ɀR���G�<\� 9l���<���n����2�F�*4	f�B9}^��q��K:d`�ȓQ�i ��j��E���7b����P�
��L`�'ގ�����>qD�W�R�{1�YI�T���IH<�%M��9��M1�b[�bV��)��2���kY -�!V�9|O*�F{� 𔊗2SfZ"w�'�=J� ��]�B�QH� KD�&�09�@�f�V	H驒EV��yR�X�n��) 
X�0g����� *�x���N�9�C�9�(����/ÞX��rpo�"5����'"O�p��FI�Z���3��.�3�
�%f�,�̼s��%Ȣ.�&�1�1O�D�C�Ju' Ѡ%�H�*���O�T�3@Ār�bn_�G&�j�nbV H������Y2���0�p=�W��q#���q�"<xmJ��}��;M�>�&,�1��:��Ջ@FͲ#�б�bA�*vJ@\��#��};�C�I�+��`DL's�\ �`�&���O⺥h� 5C`!������|����V��U�@�l��8c�J�<� 6��Eȡ=h�AjEX*�`��@��\)�0����'S��R�-=��ϸ'D
p�Vk��o���r�rP����T���m��H�I4�@�|0ͪ7�W 0����hEA�\�w�,�p=��-��ai��f��hk��z�'@�c0
�U�6�e�H��a��^�ڂ�sS�H���y�4�?'#�C�	�dL���b_�m*�yE�'jB���Fq���.�"eK�l�3%���D�4�ǯ5B|9�U�d:􄹶ꍓ�yRaL�"+�ز��B;J�C���>gܨ`��,)�� �CĻ$`�N|�>�Q�OD���p�C�"�9"�I�r����Yaw40)e���ݻ@J1b��I�WE^��P������D���u"v��:C�_�L�ўhJ���&~����UE�n��������|�ī$8�@�� 8�(�k�<qի�@xt) ���o��{�
��]�@�/&ZU!1MPg@F���jW��H�k,�1�@��w�Ҥ	�k&�Z �!�d��p��C�a	"� ��u(S8��#��K��<�P�Z�*�[aޟޭ�����L:���P�[��=��._1S�a|���t�����eB$�� Z�,�Uq:x+�G�d=��C�N#b���eg���0>�ǩ�$'2y"�û=5Z��l�B��,��ϒ/CXH��Nptp�xT�H���J��l��i���a���Cd#��?i�e4h�2`YT!�(N��U)�b7le�t�S��F𤂄
#<E����<?8pqd�I��ZQ(� ƏT��I��G:����D�'f�h���f+��`L~*B%�An|�w��c��LycbC;%[RDdǥ|l �I�0)(�+bE�F~TFx����U�DQ�1�2���cي�y�(4��$��8�� Ο�Y"��)n3�̒�d�8���Dr�>|�$EO8z)��Aci�XB�x'CNPa|R@� +4��R�%� )�<#�� �b�iȼ�(T%�&adl"�AFYKܬbSP �R�359���wf<�x�\Q���Sn��>rHa�!~�8�B��%F٢�-�%_�8���f��L2T�Ŏ-x�|�u	�<a ��T��\������]�>��'L~6D����/~�z%$Φ ��	�ņS�Pu^�;r�j��B��R��"�I��9���;B��葆әC8��@5�n�A�ٝo60�Ad�\�S������ќ W�����F5�#<��L�Jnb�ԓ8���Y@��)7) D����֞>b�B�c��q��40���)$xn��C�A+`4��a�+Y�i��$��A�5#�L��Y�J��ɡV��#�T���3N���+d�P�C��	o���Y;,/p�Z���9 ���6��I���B"F(c�J�0��h��݀O���\	�E� ,�(MV��b�P���u��n�<����8Y� �A�+?�l,�$�\Bج��E���(�M�$���d)=P�(��H�<�~�-�Ȧ��G�S��>���_�w��,=ғa���kW��f�z��'O>���0�N�>v�V�sDG�(��$P��Q���w�?Jj4�(��rr޼bŌ|�@���$���(Od��a��Z����4��?�t��]��ِ�(O�Y�LAb�)m�T���\�_���$g�$��v�Rgn�.M��a+�Y9$�1',J5r�$KX4F�y�#�y� �n��3ˈm��f� Y��y�7�ʣ��`#l���ߡ)��F�c�,Tr���-Z�,�{�5��|[�_�p�zT��!8��-�D�'r0�c �	h�*H�&�G�(����	DFP�!��h�|n�"R����H�=�(�а-[E^Z)�������ӌݺ�xa��b�����' �V蕀�@@�'h�����SF����`�(�T|	P�	>>N���h��$���Ƌo`B���FU<�zx��<w�r���ƅO`J�� �F��:"<96-�c�J��@�<�dp��妍p�E
T�`�P/�%ۄ���3�إj�RFCs�x�� �J�t�$�E��*IwhnX���'���#J٪*�б�&����S6�	�6���⢏*o �O����i����/�����$=>����ٙY�Y #mX�(Ҡ�_t�}�tg37D��P��4/�ĉ@�A��.��mzm0����-X\е�۔\	�xX�G<܆�a�M>w�lQ�a)�z0�9�c�QQ�'��(�CF�8R�6���ɾ��Y(�1=`��a�����U/�e��ĨcɰB$Halޭ^��L9��-?�0��dS���#<	�@'"�,�[�,Y�g���M̦�ě'v ���ݔ&{:�ѡN�KN�mJG �q}�aϦ5��`ˊᜥ��e�;'��T��녔����n�8Y��c
�iN<��Q�U�,��i���N�q�"��6�«,J��*����ɉoC&���� (��7W�.�aB�wU�h�ɍ�T���"�L�#*9�S	�+:�	kѥS�B(�6�W�#H@���#�.ɂ�4f�.�j��E
n�v͓Y3� �C,�H��V
�� L�qʵ#��cѰ�9F��FLs�ā,*$t���5�d��`��l�P eDm�t|�� -i5Ƒ:��i!��y�6��!"�2�p��1)���@ Ξr< BJCN�'�\�d�ղv\@�v%K�@�'����Z�y�Be�/[P:��U��m�	/^�r倦F�P����Q�˘$ؒ�3�CI- �2e߸r��Q��'���)��G�m}��%a��d{�8K�W�n���ͼS�MKVN�u����.ǲn{��3\4eq�k�w��(��H�g@�{��,_t�
��Q��0"���eP(h��V�ATnD�Q	V�Q��F'� 2�rYr�E��z�J�́?bpJ SN�$E]|`��))U��LX2�	Q5���=�2Z�E:�0<9T�H+M���e)	B%�m"�L�e�����(��gcai�1�OI�JB�5�"KQ z7� ���`���F|
� ��9�Z(��}��O�|p���۲ME�'�*���?=��dc��^9)�B,i��C���IëkI�x�ҥ�Q�r�8�`H�;!�$Зs$�yF)�2J�@����}�I��`���t�Ulʈ��W�PW�(׎={wo~�y���Ս|�TD�Y�1�h�8�&�|��fU�7c���TH.���3DUZ+�xa���Mh��z��Ъ?LJ��EbK�2h��ʌ��w�hi�ѬS41|x��Ī��'axR+Ìe����S�G�P�	,H��� |����S�Ʀ,Є���+dn0���߭:�h����d*`7%��U��15j
�1�,�(���h ̈�ፇI�P��=�J]񩟾��F*ŵJ�Z�;�e�L�| �"O(z&B�32
�D"〇n�f�q&`� c+�k3�6$9D���W�g  �|�f�d�uj���H�=)jl���5��� �3��
V)E��0�Y�"|ıkJO)b�\xr�	��B��5@��92���2��DE5&����
 ��W�S)az�#� \� �,�i�k(#��E�>2�"C����ْ�	�^�h����~[�e������&O�d�" ����AU��b��K���X+�KLG��I��|��V�Bmp-At��x8��"O�� ��E��C���nO��� M�
��U��	�%W�lP>�缳�.�7`zՃC#S��L1��r�<�#nU5,�<Z��^�|'�0A��J�;�P]�'�H I�O�ߘϘ'֬%\�('�,��e C�l�	�'iP����rA�U�ph۟h٦�Hߊ^��80'D?�O��7D�C��q)u%��u}�%C�'���r�
��ē2�bI���M�|gv��aZ�Ipԅȓw�4�K�0CJ`I���no����=���c�*�HIRR�ќ��D��w;j�Ã�9+r�+w�#8�
|�ȓSŎ����Ⱦgh�d0�Y�&�I�ȓ96|�ӆƍ�.`�`��9����ȓG���V�A
J����`d)�݇ȓhJ298�G�6m*�"w�SO3`���=6���mi��]�%�	�$<�ȓ���0��`Y����C�+�*`��B���[�A�2HC���&�z"Nم�?���±���YS3G��Հń�p,��7��7^�zTb��"=(��U{�����*(�i%	�g��1�ȓ[+�
É�=g}���Ǆ�P�ȓ�Љ# �G>LP�����(I��y�������hd)ԱQ@�H�so����g�\�z厄k/jh���G=R�X�ȓ}v�Ti��X�_�5!'T!.j�t��$QЁ���;�!���q��ȓn�E�H&I���2l�7�Ň�bh�mpN�6ReTi��S����:
�d��ėC`x�ÉӾ^݈��ȓ$'\�hQ�H2:��-��F�J�e�ȓ>��1m�>����ƂUR(�ȓ@�@�Vg��R9!�8h5.(�ȓH$�ӢC"S�"���8;�l��ȓw�BŻ�
54M+C"���sE"O���7�N# �����O(��չ�"O"y)�Ȃ,M&�,�@M�аC�"O=a�GƮ�6!��:юAhf"O�,��-�l�����
���"O��"6@JZ�L)c��EP���"O���&�+O�Ru�W(ר�:��"Oޕ��[<Z���x��"Pn�H�"O:��¦X�D
e� D �@"O����'L��i�E���T"O褱dJ� 9��	rC�+>V(�34"O\<�7*3Tͪ�B+&Y�!32"O�-�!@@ :V��u/��X�$x��"O�1�Al)x�d0#�;�R��"O�A�@iH��rX9&+�::�D[�"O� r�p�/�Y��ͩbj�x@�"O�9R�� $ ����j

d�v���"OX��Á�$7�r�� 1^��:!"OTm���Y6���i��ċ�"O:xzg��a0�a�r`P0bs"OB���k�������5a��`"Ora9��M�R���WM��e��"Odi��J���)�`دs��@q%"O���3��i�p$�FNJ��0���"Of�& ʀ!]��n���E��"O��)SǕm �֭-7}6;�"OXMQ�kIOlL�낎�9>=J	��"OB�(Q��%���BG�����"O�L�ì,52e���"�ꙉ�"O:ȨS�	=e�3DE
�Hh)�"O��Q%�� ���K�DT
}YKS"O�Ih�/A�`��ٙ���7R��"O�P$b
�ֹ1�DT0�r]��"Oе���N�z5�v↙0��}۷"O��$��(W0F�V�H��"O������w�DE��&P3d����"O�!`J�z��ը�E[�XEa��"Od*���;0����թA,�*�"Ob�"t%ĝqھ���Ņs<\t"O�谷�8Zq���% )��xq"Oj�A��
(���T�չg�2T�&"O�6�Ϋ �LB��IE� �"O���
�/��`XB�F-�e��"O`�Kť�5cl����PG"Oؤ�#�I	��6"�#ǚ��v"Oh4�t.[����e#ۣ�Zp��"O����\
y@�Y��#�-b�v,�Q"O����R/Q��(BBGP��s�*O"��ǜ,�@�� ��2��C	�'�x�:0�84.����P�J�V�r
�'�ĩ�蕭lA�d*Q!�B7�e�	�'m
�I�΁�q.`A�۟�&%c	�'l�s0��JHi� #ܣu 4t@�'M�� �_����mR�z�V�x	�'���aʤk��pQ�@ތ|�p��'��yJ3^�x\:���7CA���'I�����+�
�v�K�C�
��'��iva]�7�I+&�B-G�����'3��f��e�$�0ƃ�5�����'�4���	\��P��M�8�����'bQ�w�YO����P����I�'����>T@� ??�8I�'������w̢��g��%84")*	�'� 1�6}�����腼.��R	�'��!�-U&[<�2�/�ta�a�	�'��8�.�8:��s���dQ�DZ	�'�ĩ:��¼!@Љ���[Vne��'0 Q��^dxČH�.�q>T0�y�Sp<P8!# Q�Oa�x����3c�>�[5�jK�q��'�
S��RF�ib0ߚe���-P3�z�;-O�uK�4�3}Rjǡ,.�%�`/��v�B�ˀoťŐxRH��r���$�@-�sLѓue���b�#�\y�ɔ#<����^&|h��5cW�s���P���ca�x2�֍^
��jã�l$�����i��|�3%�3Pd�IEfV?Dj��
�'�X�P!�FV� 4��5���X�O��@a��:b�A�!�)"(��򉎤=�DȹEB�s�A0��;�!�$V~��Ӈ)�$ot��Fψ#h�t9�g`?y��,B�f�	h�ڦ�����)�� H�^'R�q�!S:�x"��J��wg�5@��Ź�^�hBNa���(}zlmktIXO���)� �9k��'5�A��jT�a�bHg�'M4�!m�S�|0���pڔ�0��?$���u�;I�Fe�H�	�y�g�������֗wa�	#�'������,�Д{���"�@xb���(����q.ӃC\젱%�U�g�r��"O*�:�j�3��`�@��fO�A*JC)���y#�	'�)Y���&T��ϸ'r��j�%@W,�pGk� ������9��XIUnK�d� �Ѓ]�jǺ��&T
yӤ(! N�6������p=9�cǳGZ���[&!�����q�':�)�d�B�,�`��Gz ���?c"6�v�R։Q�Yn�C��6D�\�qOP<zV�!��O"F�X�3�>�B�Q�Zs:$Y%�<Π��gH�}�OL�u	�'T�Gl��" �hA�|`�'��9��_�.w B�f�����`[Gj��RG��#Ҁ�8�蘚��g�aH��'�sv`��e��S]����).��{B���=��ZS���X��r�!M�͡���,3���(�O�}�
҈���#c��F�����	�x\���D�Ŷ5�� ��P)C��1�'Q�>��A�\tW.�`WƠ
I,�ȓ�|���G
��v�0T�p�n�U�9 �h#ݐL{vjӌ^,J�R����dUY����*���GLZ�f��/�y��7�(蕃��*���KwoQ�Q�BQ{ �M�]?@�H�?q�c�Oh�Fxr�=�>I�08-�z0Г��>�0>Q�7����
VR�Ш�(A�]�.d�v�W�i��:������h�V�XB�H�
��H�FF�(}��0c#0�I�g�n��c�m�F-MV��9Y����|��h'd���"�ݗq���`�c�V؟�Ӣ�QOa��c�k��qPe!G��Y�`�q&۾r�`�r�e�t����5��d��{����Ƙo�ڹɐ�DH���AG^�8:.=#w.�z6Xa�$ߩw��%?%�d�7R��q��݉�>Qz�J�Fu+Eh��ơ ��&� %�TN��Q��"<�u���W޾�a���5u D��-��<i�m��xk3��e�5�?�x%��>	4q�F��,Tz�� +�S���#�e�R� �r����X��81_�����	u�Z�`B��2�)��49�H��u�@H���0����g�"��*��A2&�Mx��ڳiq� r����U(�}���I��FX���&:��,H��7g�����7:$cw��#&��svm�"-u��s�s,
Z�H>`����'�68�Ɂ# "��;��!h�|(��͟f� (���gT�Gz�X5p6���R���6a�7'��+��\�d�0����*~0qk�HI� ��ͰE���o4���w��4q���`*��_�8��&�L��O�Ԁ��W47���A�N�K!�iR�vfC {��Ⅸ�s!Jى1E/ij*,��O�]�� g��_
 K�'}�аz�g�h�>4 �B�0p�d�w�*V|�|�f��p8H p엉0�\�B�L�:G`�1J�C  �x�hCȔ( θ�SD�]"w7V,H�,
6�N�@�Z��yW&�0b�V<HG`�/"�\�2�@���>�b�� |t�xc������:�I��}OB�	�AP���90H�A���G䅜Pٙ1h����b4IN�~IH�1a� �m����t
7MN�x吔j�C�
^�"=ᢆHo ���ǃ?uGT��5�]�,i�a��_Uz� ��XPԭґ]�x��2�^SwN�y�)H�B�4!���(D�	gę�(O�Q��a"3j���o�0sǸ|��iu4�{�&�4��Qi��	:�Q�������Qɞg�E��#�x&�H�B��U@�}
I�?��pg�
`%(��_�B�����_%{>J�#q�0�hI�e��d��i�7Å��vM�'���ߴ*��p��i
�0�2�B1�y'ʐ?D"��9��5�`��
�ư>����75�^%�w��"w�n�2bP8TK�uÐ#�=^ژ!b'�v�B�J	�l~����A�:�r�Ņ#v��D�A�|��+6�zɱAař'�~ԫ�z�z"=9���{����@~0�����>E0�g�h<ؐҰ��'}&���]�B t����L���A�W�C;G���S���o3Ƭ�@�I
���@�`0� XХ)ԣz16љ/ jv�ԇ�*���
��1"�c�68�9�Ԭȳ."����(a���At�Y�J���R1�0>AC�_;;5��p%ʄ-< |Ѷ(�2O\����-U.d�>����զ���E� ]m�.�6�IZ��V3%}�q�Ua}"b�?���v C�B ]�p�V&���,7v#��O���7�i�N$�C#I#lP`3*��V����6�=2�<�1��.e��(ژ�(��V�'G��U⎌y��p3䍍b�\̲��J\!���LI#@�hH#��0F�8��w�܀[˘dx��J3-�8�j�{��1����$O�"<���K��un��)Væ+3	[�J�r!=;�8�2�l̳6�����d�`}����%K�͌�}!>PZ��7'��-2��Kz��Ԣ�B�'a�ic
�G�����:b�8�-W9�L�H��%�H�K���Q�p�I$A���H)��f�7m��&x��w��U�q�I��ݨ7˘+h�V�p	�i�^�HAo��uRl(��2y�$��jĲkyU�ش�z9Zf��B�^��
򜨰�V!`=��q4�T
`�� �����Q���<^����Vb߸Y��Kvx����Jr�H�B��� Lޜ�g��T+�𫕀ɒe��|��@p�6MŖy�"��K���s!O�5�Dp��@Q�'Sp�BB$�WT%�c�@��X#�'�݈�ʙ�o04���[+-1^=���?�@Bhr����ԓ;(� �ыp���CX�r���S A#�(�� �O��A��i=���C��I�猝q���Vرm�9OPAt��qw�j;���F@�B��!$7�� ^�2�K� gV2ђ�e��Fj��U�'wX���D��J�O�:F
 (e�QD���*P�гAT����	�B��"e�	 ?O$`���@
���B8emN8����%3h��:,�axRB��%~��k+iO�MI�A]03a�@ bܔ
�c�%d��`��F�e+�QA��  a:�TRv��&hj�lX��$��6� ���%�Y����e���9H
�I�ɖ���Yx &��F2�����O�~�R��� H���X�6�1P�G�4q"A3R"O���7L����1֪�y\�a8x�zT��m��d�@��0�@���'>����.8�睯c���cde�~�m��K��'f:C��/b�����g�(��ԄQ��p� B��-sL�QɂIB�#A�F�%��ĘB�?�HO@	�4*Rب"E�#*��c�'��`���-�-9a��e�L:R�:��b�����r��uE�5[�`ȃ�(,��$�/�܀A�V &����kF2��O�٧�׎a�ZGC;��r0���zZ~�X��6h�6��%͜$�P�L�#�v�(�"O���&O19�):r΄�S��T��f��)h�0�#n� '�V4RuNL�}l���|*�.4~j�NY6*�
�S���#e�j%� ��B���[�ft����76O���tGۓ4/:v�(��a[�ğ-O~�!#�#gp��҉��6�̤�ue��I�~����az�iL�n�����r˾I8U�M$�*ٳ��#X�����k��h
P�S�y3n��ēVx�XXg���9h ��Wh�O������&-�� ��.��l8��K��د���yz�JU̍-|�
8��\�Fi!��}�D!��JI8�b1(��ݪ<J�ʷ��H���Ӏ��!
е���$��C3 �m���C��2�]# J|�<I�GGiF����$_5qJ��b�ZFr��'�� �Wʴ��Ϙ'[��`��<zG�!3� Ľpی1�	�'lr<�nƗ5�!j��I�S����C�nlA�9�O
�uc��k�lx��
؟K�F��4�'ִ��f�U0�ēN�\3� �"�hR�`�/X/��<n�HZ3&
p��ܑ GP�T��Ňȓ1���0��q��Z*7<ȇ�����7���[/8��Մ
F{Tɇ�d��9igK�;qzj��h��0��
��Ι:��zb�<��W*�p�!�(Eq,	
c�3=dP��yx��	���[�hE:�h�!@e��3��I�#+MY#F���Ɩ	�fy�ȓҘD��	 Ya�)�L�6���.����I���8����Щ�ȓ\I�9��
�f��m�e�V�����}�ͱ������-0���0R䠇ȓX;�$9b�R?����`\7��<��/^�[T�Rΰk���^� Y��;�v�a���f}-�c�8:<��ȓ3��A2j��R"Q9C��:f�$�ȓ)�r�Q��m��`B�:/�8��]����`_�OZ�����/)��p��y4@�ES:� �u�ګ����,l|HR2̍�t�|�p�^� B=�ȓpǔl)�� t A�v��ȓ}�*�[�OΜ2�0I�BC�%�ȓK�J�)V�W%~2�pb����]��Psd�����b�B�pq�P�`�$���� �Ɣ�4m�=h���8
ȇȓp(u���;^Q*A���M�[]*M�ȓC��i:�ݡ�ȫd@��مȓ`�>`@�oXTx#��&=�)��2�L(3ꟹ������H(Yat��ȓ@k<� ⏔(S�P�wђ:dJD�ȓCHH��t'ԿZ,0�ՋOJ5~��ȓ7T�,J����d�@r�.��*CD$ ��!��<y��P~2�[��hES���8 ��Q��
��?A�����	���5W�X��5}��teхV�9aCޭݴ8��JB�����<[�myF����)§�)���U�s�K�	0�͓O8��P�����姈��,I��2_�~�� M&q�%ڲƏt��(��G���S�i#�iiݱCg� �i�~	�ŧ�"��B�%Y�t'�������(�,��'Z}�-�H|� �@��W�[6\hi��RՓ�+M40�|Q�u���?�1e�)���v�O�b�iQĕ#ꠠ&	������xRmR�3&d	��O���8�<-���&�
��	�/O�@:�'ؘ`*�&�����%yp�3*\D�'��Ҽ,�	%8��$}3�S�O�0i�sf�O���xC
S�enx�)�?f�8�d8}"�~�'6�����-I�!�00��&Í�)̄9b�����?1r��1O�O[�Ѱ7�Ȩ!�$��J��5��<#�}�JM=<Ί��Q?���|��h�-5��!pIN��Ǔ78��'��!1H�����x�ᖇq�E�b�:5���`�N](�?�/7�˓�~����o9����7�"��r���&��d��� ��~Y���ϸ��t,��7Y� �`��?
A{`/ȢT�`�8�Dj�O�����;	똝B�1�4�GE2��P�1�0�We��O0�h�͔�Tؒ8(�L5{��/OPeC򀐣2��OQ>�A����81L��C�: �=��O譂�T�*,2�OQ?�*��C!H|���o�+3��.'�J��ŁP�>DbOf�O2��sM~��WH���,�ezu��ʟ%_�Ty�D;����U�.��	�,]{��CƩ��j�⴯�*Xt2�ڥg�>�GKT'}TTŪ��9O�Iؼ��`&��9%�*����u�����)��-��'J����g�O4<��dOۋJ�� �# ��D@��O��(��$�OP,"�Hގt\�Yr�8p��P�"O���kϔl�A�S�T�iw�x�"OL�+EřP����C�!bԼ�"O��(�Ń<`�����$�\��1�"O�����B"}C4���"s`Yw"OT�ki�3u3�rtG�8ވ��"O^|�F���$�:PfD�3��Qq�"OB��G͍;�3���,<ز�"O܅(0�
�$�]����{/�h1�"O��Q�䐲[� b�܇R��!˖"O2t��FU��unU'X<���"O.q�`f�p���U	����"Ov��g���*d��́t�Ȫ�"On��IH�ȆU��|a4� u"O�l[��.�.��S��.O��2"O��3�f)��J�p7�Ũ�Ƙ"�yr΁�>>��R�I
�{�I�&�ޝ�y��Ч(�ldȇ�R�nb�IV���y���4��*�d�,gxإ!uG ��yB��S���a�#�]&��lU��y��$4�t}�����b��@��G��y����q_8��V��(�ځ+� /�y�f�/{4�3�#�r�B�(�y���9J*�P!��{$e��ײ�yrB���:��p��A�Rd��yR��?]��E�tw�dM2!	�y���~n0 � �HhY����kJ'�yҪ�&F���b��?e%�Mqg`B�yR��y�$��L��+q��yg��yBfN,R���PFM��%ϟ�)q����A+4�Z�,V�i�J�`�OHI���%����ڬd���A�J��ȓ��"#���O E���˂d�2�ȓ#��X����<��S�Җ2jy��4�AJ�B�FB�3!���/�zE��|"��x�hPb�l�r'B�
�&B�ɶw�ܑ�G5���Ã�A�B�	z�ي�@M%2�x��(@�B��C�	)=��Ij3a̭)�0PK��a!tI,D�Ȫ���l��y	���/ �0�@�/D�\�@��G���ɤ��Jp�`[��3D���A߲(�h�o�Zg>�p�2D����EƆuf��A�JaG'-D��pC_�'�`=J�a�S�K@!,D�䀶�'d�T(�6��?6���+��)D�� &=#�N�1R��p�oEci�P*�"O�%��$��Lz 	j�נgdB|"O��a��
�e
�ҧ��QHXɻ6�'�Q���Ţ.�k��l�ظVc=D�8�)��z�	��&ZuZx�z&D�ps��Y�R��٣��X65�`&%D���D��$H
��)��Ո ��YuO0D�$P$�F7J���(Ä�*H��5��'*D�p�DLɀ8(�	���58���b��"D�l�e�J g��T��KMhŘئM D�ȱ�ʅBX�Di�j�Z���!�<D��ZQ�ݓ[o:�@�Q9A�<�ip�:D�t�ѥүX�p��Q`Q�|}D(HD�7D��C���ߜ�{TKĂ%�24�5D� W#Z
Z�<`��) .D�q�h-D����Aʔ�zP	6��9��tY��*D�(�ү@�(��htKɤ}Df���'D�����؉D����S��.@*b��&D���H<R'.U�Dg@�}XZ�
d&D�t*$ɿz����� 1Dޜ�ѫ!D�8
T�]	W�.�ᴬ�k��$Zg�,D�D�f��J��#ff԰]��ā�d/D��C�U^y oӢi�� �6�,D�ГQ��|ֆ(ې-��Py��l&D��#�ؖe�U �
v)1��U�4�!�D�$R^���H��
K>���`�<�!��8VPV�0���&i�+E�4!J!��Y�$���7/���l�T���fa!�D �
ʪ��������B��G�!�DʥL�(A��,|�]�p!�$5S!�ӡ��(E,ցGkr��W��'UN!�䂫h����Z
3_�(�4�E, D!����.�W��8D����\2!��`����Ĉ�S:�Qv�
G'!�$Xr�N-� A� �t�%�A4^
!򄎥|t���"� ��R��!�dɘ da
���ڄ
$��J!�DUv�hđ"�=�r8�g���'!�d	j����V3[}��s ϒ3F!��@Y��UY��C�e�ta����F9!���={.�6�� }b��yp4!�d*D����{A�4[�lX�N!�dH58
�ӏ��>�ڃ
"�!����a�t�d�.^���d�Ȋ+�!�dS�t���a�̧2��5��IX�V�!�D�z�4�Fl�?D����%
Z�!�D�d�n�ap�N��	�R�|�!���ob�AIV��-Q}�P����.K!�dD��m���ʇ\b�ڔkY*J!�dԡrMڀ�b��u{��
�N�7<!�d�#V7xu@�e����Z�N+"�!��Z݀U+��S!���R�#�=I�!��O�-����'��0A� ȣ���s�!�d1PD�ĨCa^�;KZ��T�4N!���*�f�v#SM�W��(!򤜓�j$iD	��N)�x+U̕)�!�k�"p�d�ڕt2�	�1J��aM!�ėaO,���a͗R�����hQ�q�!���(<P�E�¦^/ߪx�'�� �!򤉅RfXu��J�x��H��$��6�!�d���R�2��G��`:��ܷ7|!�$T#1���saS&�9I��\o!�޽@���"������F��-q6!��U?�TU!Ν�9ؔ���n�Z�!�� \�
����TR��%��9�\��"O�LР�>�^�0FO�a��4��"O�,:4�	�1Ŗ-k&aˈG�.$"O 8���#l-����2�R���"O��j`/@�IZ��C��G�v|Y4"O0ఋߤPqRhY�%^�_vP`�"OVQR7ƀ��l�I�דs�P�b"O*%ic�U�}��P�%�$G9�ݠ�"O��� (Y{v#�=#Z��"O��K���(N�������!�b"O�M!�
�]�r8@���^H�p"O 9� d� E�պ��T'�d40!"Oi(�a�Np0�CU��'\��"O�(oL�!��X<�
^!��ķ@:D���*�:������@�qb!���c�����V./��<�@�OJ!��G;Xt=õjW-(V��W�.!���?f�d}����
��]�g&Is%!��'�c��� �0yrfo!�D��=��쩳��4$r�2��%�!�$DdOl`���;�^\�ߒw�!���$l)45"u-�"*�8�!dI�L*!��Z#!?�i@�֬4����6�'.�!�$[�p�:���*��w��x�E�!}!�D�=۔�`�ᒚ3�B�R��WjP!���J<r�S�,Wz��9�Q�da!�d�+(w�vL�y�Bj�7�!��~���܂E�B$��1!�!�$���%��F�{��2l��$*������nZ�╊�!�$:�jy!F�F}Z��P D�!�9l��0��ር
FB�"@N��!�$L�`A���A۹.���pvD�l!�dө?�|�k��_�(J"���l�!!�D]C�Pi���77�X� nA�*!�ě.kxD9p�<C�, ��N!V�!�+�"����N,׺dv�ע �!�d���"��t��VÊ��4
�'�`���j�x �2h�%h�s	�'�x�J%��/+0�2$΢R�(qQ	�'Y����[�=�Ԩ�@Ĵ^��Pc�'jp ���U�b��㗣�5P�9�'����G��
�蛂Fm��'r�M�7)�uvH�3���=��I8�'�RU[h���F���(,����'��Tk�R�V�8s��_%��X8�'�z�p��D�A��#��"�<pr�'�vP�
�y��h�%��T�E��'>�Q�D�*�9Y��)˦ �'T��U��r�0E&>�T�0�'ט� F�S'%�n}���ԢL2�p��'Ŭt� ����E�U�'s�t�
�'��}h�\
cQ���uL��bj ���'-�ɰ�KΌ>Bꕠ��Zմ���'@
=����n>��G�JO�
�'�aJ��D4/O ��"6|�;�'����� !m���P�P�E� �
�'�:yH���NC����-m����'��BC �7s�8l	v�K�^T�A��'B��eƌ3~z��0E�CaVdX�'�Ju�g
>y�C�@0�ؒ�'��	���m<��K6C�+8�3�'¸e�`+��{i�uYf��d�2�'؄����
�g��B�<� ��� �<Ò��!0W����m�q���"O$ɠU��$X�(a���Zl��[�"O A9�iX�{�Ayqn	� J�l�a"O6��Y܍��b��p���!�"OHҥ�"9�ʥˣ�T�6���C"O.U��k�u��MHVA�y�@"Ot���$˞$vH�A����S��QQ"O��:���6[����d�)�.m�"Ov�چ�T�/U6�3�V�W���p�"O���u.I�'�
�i`f�B&`�$"O����i�hU�yB�F*s�P��q"O��#g���\(���?�z�+�"Ot���b؜%˅��_ib\#�"O�!h�8@��@��%.f�X""Ob\��/�--<y���N荹`"O q�t��;���GG4?��("OzX�a��z�P%�w/1��"O�E�킴o���uO�:$^�l(D�$�/ǧ9֚![ũ�. ��!D�$�M��,҂5�t�l0e�?D�l��13B�	�!S�U�R)�T�=D�dۃC(�����dФ|�D�* �=D�����*C�V���B*��	��.D���W#�D[���&����������d�Ob)�U�`	h��	����֟�c4�8����^���R��Ǿr��Q�=�`���ŵ���Ӄ�(@�I�|���R)�剭~)���#%C�T`T�顉Ǻ̮��D�?4r�	����@4j���4��	œPtMi��μ�ÃU�5�ჲR ՜!9q�^�>�|�J7 ��ǟ��?9���?ٴm��Q�L'�xp��� r��Dy�'Ԭ����AtH�a�n2N���'��6M�ަ�%�T�S�?�'cNu�1��81r�aƂ# ���R�
e���Q�'��'x��j������I�h��D�h�!00@�sFڃp�t�CJ�E��X3�M9K֣|N,�{��$[������U	^�*}�d��6\8u���J�~V��5�؜y�0l��$ЬX�v6M'����n4#��a� �p��y �#�9��@3 �iO��D�O�����u,�r�H�&�8����:FqO �L�>���<�ꥡ�('0t��r��A�D�ʦ��ߴ���7��l����'��pPvj�3���$�@�`���O�9r��O��O�<IelL�3�
|b'�M�5��1i���R�=�S�Y�b:0�2^�q��a���Q���#	T'%z�c��W+5'����'ه�(�#/
N@5��n�
`
�O�(~|����ɟ��P.�0����M[ �~"�3\��3�J$�&�P�=p7��'�O�i&���Xn$T�S��o����F�+,z�����ۦ�#��< ��m�p�j��v���?�̔'��-��Hz���d�O��'X�������M�7 #3������B����eeD�|b��S�mo��)u-�p3� yd�P;	cdE���߄u���غ�#	ظӢ	P#��5��Q�c�IG}"	N�r!��D�o�x�7k�]�ب1gA�J�f�Gș{�l�q�
�F�:@Π������5�~��ď Qfĉ�qEܧ\�����7��IǟĆ��S�qu��� ���9d�<��,��f�|�B�O�����b��L2��"�)��,���OR�D̖�B���)�O����O�����yG��S�R]K�
�E�Ų!OB
���&�Y.~P��GV1��0��O��deO~�H9�XYrlG�.��}j{~|�ץK���d�2lW�s�0Y@A�n�Ӯs��oB}B��c`P)�p؅aDr\��Z��Dm�x� �������,O���w¤N� H�em�U��7jӱ5�!�dW�Vp��w��J$DEO  Jv���2�M���iY�'d��ty�]�hy�D��n��PH$���]� d2N7�'"�'d֝ɟ��۟L�E�� �||`Ui[��@а��}��6!FF�h)�P�A:
9�3!��X|��<�7E�q��H��#j:?R!��ѐ��
��8�n\�SS0h!5e�9j�Aу(-�<��TmZ$=S��A磌P��a H_�}� ERE�i\�6-�O��?��'�P��f%� MΕ��S7"�����O$b��&�
�`�S�ȉO�5��c,}���7��6�<��T'�~RW����   ��   �  �  C  �  �+  �6  ?  qJ  �T  7[  �a  �g  4n  rt  �z  ��  >�  �  Ó  �  J�  ��  Ь  �  V�  �  P�  ��  j�  ��  M�  /�  Y�  �  Y � �  Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�� |d��"O
`�(�;���8���-0��1%"Oj4��ND^[��"3/9�0|H�"OB���H��*�ʞRy=a"O�味V�!X��!&F�:J�$���"O,��a
���C�Ą�M�"O,$3%o�-���p���+Ն�:1"O��ݢ1����`���y14]2��i�<�6��{_���c�H�`�fX�$Kn�<��A̼VI�xR[�)�Ć�pඤ�ȓA5��('nߡ4�� �)˩%� ���,��r�؊b#`T�eT09���ȓ!�b��g��}�8�F��-? �ȓ
K|m�ș�VṔ���2�%�ȓ"R�X�j�4JN�1�˘X�i����̹	_�jZ��1!g��zܶ��ȓgil,*�J�
j�Ne��i�J%b���f	�(U��:���G��$Y^م�~r�� S�%T"���k\�jx�ȓ|4�1�îJb��@ӵ�ݩn�V��/[`�"�v4�R�!ʎ<��M�ȓ`:��z�ؚh�J�Z��$HY:	��H��p�m�C1��!��B:��0��EnjZA V;9����J[
2���	��4'J�EA�IVW&��~�(aZ��ӹ�>� o�Y�|�ȓ�f�A�
Ο7�H��M�$�����mޠP����/���ANXo*�ȓTv�����{ ��-7�*h��I��sB�8�8���3����ȓNe*M�悡;������X�o��!�ȓ'lj�#F�m�+R&;�|��2)n�C��0S4���T:
b���:�0!��e֊��)��ͷV��,�ȓ0�&�8#���� ع�L�����;�P�AFd���,w�6d��r�EQ�( �gVlɦ�M,H��,DP���|�I	$G#\���EyY� G��B:F���2�)\�qxLIY�nݣ�yRkMH��e1�k ��F�����y2�RT�0�;�5U��0����y�l_�i?�y�GM� ���W%��y��8Vnd18����}`��`����>�N�(��ӸbT&}i�T�\Ips�*D�h;��3&�tm�7��X�"e��'D���փ'���\Jԑ��#+D��
1���6)&YhEn�>y�Q{��$D� �f�B�
�� %l'�4��t�"D�,����2+�R<[$T:i�"���$D�T��f�AR�\��L9�\с�!�O�Ov��с�H���22��o�>5�%"OTC�C�:- 1�ПKF�!5��6?���	R+�vx�doI1Y���t�!�D��rb*([�a�2RW���k\9т�=E��'�\�b�˒�?D��y�`Y	]�4��'�Ȭ�V�|ޠxqu���HD֍�-Ov���ʒg��Y�iJ�L��%���$@<!�Ě�;Ŋ��@�z�-���a�!�Ւ3F��jĭ�M�l��3���3!�Ĝ&c�D�`����e1�z7dW��!�_�A �2�˔m��L�=��f�|�)CH�Rt�זGty�)F��y
� mPU%hϮt�I�=�-YeX�L�'�0����3U�(�&��)~��a��o�!xy���N�O��n�O���P���TAR��k�B�-S.eJU�t�0Dr�P,6v���y��%��#Z*���.8�D�`�N���C�ɽGp!Sd�צ/��0s�\�z���E��u'�8n�y�����]�6��������X�nH,(�!���d~h��N3�~�$� ��'�a|��	R��x��Rv�p�1j�1�~�0Ob��SM�D�Od��M�a�Ra��眱B)
��d"Oly3���A�����Ϥui&�!Úx�1O�)s>Ob��'AV@9r뚪L�xs�R�<hT��I^�ffZ�R �QZ%���Y5/X{�'r�iP�)�1[�FY�pݸf�M>�M�<F�� �B� ̓@��.x|p@���y"g��RH�`Ӏ�Z�8��D���O���!z�XZ1�_�>��h�s�!�D�o�阒�0G`�|��"��ߐB�Ɂd&��h�5��W3I3�C䉡u򘩪&�ݑV ���Ш_B��C��'?�Aq�j�w�8(s ��VݒC�I�[�X�QB��# �8 �σ'�nC䉼_��S���SZ�ٔ���~�PC�	8*|� �P�NNnᰂI�N�B䉡)*`�F�v��fŚ�t��B�	�i����%�5f:��9�B�5qs��A"��)M&��hê��B�	d����c&�`ڱ�kD�B�ɣ^�2��g�]�L0�@s�4�6C�	]�|�A�РN�������f$C���i�G2S���i`�	��B�	J��l83�ʰ�`����B
~�� �h����N�<�S�a(BY��h1D�ە�$��ˇ�jz�e{�A�mw�̦]Fx�I--���"-�����ꍵ>��B�I�F���A���,��D�`�
W�B�I�Z�,8����o`�<��n[:<�TB�6}/T8�!F<;@ua��6\*B䉛��!!����V���E#"��C�	�/�jy�3���D\^@�U ��C�8v��L����0�*���I�q��ꓵhO�>�����4R�De����[�J]G-�jzQ?�0���B�`��
�*���p#�)�D,�OՁ!([����"�;k�zp�O��=E�T��&�z��iգa�й#�§�y�^�"�)(�B&0��y���4��O�~J6�G+�V]�d#X`�LxN�o�<��l�@��H"Ş�
O����g�<���^*pF�0V�,N(Lk�Kg�<I��'��a���& ��R&Ra̓��=���I(F0T'�K�Z��p�1�Y�'7��o�'CRN-`�C�Tn�H�fN �<��:b�A�ҎI<H)�h�AE՝9$�5͓\��"~��IY%+Z@)A�
�=�ȅAb�N�<��/	��)��iC
Z�plyb��By��)ʧ����f��u�����'S�чȓ!�̤7%�/u<Pw�	x&���ɂ��?aUI�r�؈P���z]�<`��XA؟��\?��PIƫ0j�TA )��هȓ�*�(aQ>T��;�` �7��܇�S�,:'e�g'0�+���6R;�]�ȓJ0����nȓ�����߮0j���hO�>1qBN�!c!���0*:)!�&*�O��%�^����Mz�e+��O����S�? �sr��!.�:=��ˇ�&���4��W�'��Ц�����2W���M�6MS��iu�!��	q�nly�A׾B��q{��ڸw�<a��T>���ВXZnM��WWN���&F!D��)��D.;�֥��S ./�,���<ғ�p<�7L��kU�1��Q�[\I���u�<a$���%��hQ4�(%��X�<y���q3�h��1Pȱ(aʅj�<y�_!j�mBs��#TH`�#��n�<�c/,=hD%qbA�
�.8�@�Xj�<)�k�3YBL:�IY�|H�Uq��]j�<ɢ@įW�:8Z�E�="�����MP�<��gD�WPT� �,_�c� ��WM�'�ўʧDhx�B�Jަ|��(r1�ɩ<�DB�ɪ|@�iw��9[:h���\��OpO4p��� ��L���<4�B9�c�L�_�!򤚼|L:�z�
�q� �Y�* <��n�爟$q![!C�ț�.P? ��2"O"�� hǀe��5�@(��6��9)3�� E{��)��r�R��T&Ϡf{�� &��v�!���(E��*�C�H~���w���1O����O �s��O��L3�/���J ��Z0�Y�N=�h�h�N(,��5����R�{�Xh���r�܉�ȓ	,��ؒU҄�L�� ��=��m7T�y�7q� c�
t�ȓp���jU���0�;5o\57��E}"�S�:+$�)��\��PY�Ѐ�'2�ʓ�0?� ٽc���#G��9ؔ�%mo�<�t������ΟV@�qi���k�<ibO��4�J�
�9�:���d�<�!�
L.�
ôk��\f`�Z�<1��e�A"���/��Th#�_�<!�'7V@�5͋4D�~azի]�<Q���5�T�{d$U�"T����IO�<�DÎ-���U��% 栕 6��J�<�a��^	�]��b!�8�g�E�<3�D�1^��dʞmR*X����f�<I'D��R��3wə�&{6�IsGl�<!��Lp��g�����!FLVf�<���?]���i�D�hi �^�<�B�'7v��2��J;BaG��q�<��CL�PC:�cU�\$������s�<!֡A$>��X�wB=�f	�Kn�<��#ɴn�����E�ѰF�@E�<�U
�[�*<�VL�PI���[�<�ġ�6a���"DD���]��W[�<�E��6)𑬈
"=.)pp��U�<1q �.��I���,/
ɳ"K�O�<�ϐ�΂\Pg&��5���W��S�<q1�{Q���WnGv0t��JR�<)��>b��D6�"UJ(`
�S�<�GB����I؅Œ�`�0؊�[R�<��*�\	��L�vu:E�K�<��3;���HЃ)��J`��\�<���U�D
"�q5)	 xX����R]�<iP�
 �3��Αw̍��MAc�<��Bް(�'B��� fAFt�<	`����И�ʟr-P-���i�<�FgػQT`�;�CəUr8����De�<����~k���b��0���X��JU�<A���	Za��:�F�@̾����G�<i�h�
r#���7��c�ß|�<9�$ո�8�aKV�$�h�#��z�<� �:A�[� �AI�߄=�0"OLX�d�%4�X"�ۮ1�����"O�<1���R+��iקM�u��0@�"O�XQ��ߜ(5��O�I�>A"O�p;�gq�1b� ,u��hS$!��?���?I���?����?q���?Y���?�BA�v�daB`EM���#�T��?i���?1���?����?��?����?i�.�kjaH�E�:�����/�?����?���?���?Q��?����?�"mXi���Z(8���׌6 8a���?����?���?���?I���?1��|�v|��e��M�h�[W���C���?Y���?)��?9���?����?���e.��m��������ܑ��?Y��?1��?I��?a��?��H��\��2�6	H���:q�|�����?���?9���?���?���?���d���q��	�=�#�M�	d������?	��?���?���?i���?���/V��{�!2�h�Ag�^�<@��?����?����?���?����?�\d���懒>�8�Ҥ1f<�j���?����?I��?1���?��?9��f��ބxO��(�-:ƬՊ2��O����O��d�O����O����O����O�����ÎA�0� ��� k�'�O ���O>���O����O>�D�O��d�OT�!��6�b���OCa�^$���O����O��D�O�D�O��Ħ��	���u.�o��\��I�BT��¢�����O�S�g~�J��4���@ Qxti��GG��2̉�J�O]����M������|��M��$��`��i�x�����iQ���'[�m���/��Ĉ�Y�Nx�хƤ��S�wR��Ş��Ɇ�9c�b����^yB��:F6�HT�ta���)S ��U��M#��Ti̓��I~���y���R�Z�qƍW�6�-�&������uӒ�IyyJ~���F�V��$�~_�l�D�!.��Cʗ-JZ���C$0���J�;�٪��4���DT�z���#���*yo�dr��4��Ī<�K>q�i6V�i�y2�"L+숃$��C����ϟ���|���<���M��'F�Ɂu3�@��!��(r�˺��O8y���2�u�P�)U3�eRQ��O`�3��ƮS� ���E�<}6��T.�<�*O4��s�� �͛WXH��h�1��9��Ď즍��O(?�ſiw"�|�Ob�`��"L�zy(����ҔB��H��'`R�i}R"-��`��O�T$H�
B��YCcЎ�|�ˤ�žF1��� �#�5�s��'t��T�B5�a�� \3���"f�N(jiX�zrG�k��\(�����Тo���-�P4c"OL�x#�i��
�Dzp�#3�.P/\�q0d݅@�DtP�E:<�x���Co��U�B
{RK�u�$a�`���I�1B#��6d&,��M�O�<!x)>���2���':��DM�}�ZQ���� 9<��B"�H�[�l���*��.�I���>b�X(����F�:�b�P�8� ��'h����O��4�	�'��قcV�`�BYS�M_� ���ش�?��>�IFx�O���5ƫ��T.r���܋wa���1�Z
�Mc��@�gZ�F�'���'x�t#+��O2�Ze(�%oRL����'�X)*��P��U�3�+�S�'�?q�O��%��n��9{��Ԑ����iR�'����*<��O���O6���;}B�48�?+|�ڡ얥,gD��'<��'����O~���O
�d�O�4(�.K�\�T�h #�>���Gئi�ɵ3�0�{L<�'�?I���K�i�ԨJ�jQ�u�0N1*rΜn�ڟ\���6?!��?Y��?*�a0�I<)z0;�d�z�UA���(w��'�(��ݟ ��Ay��'w"��(��ȪV�Iْ옅ǑyZPa�y2�'~2�'��IEo��Z�O]B0c C�|i{!,R?�`�+�O,�d�O��$�<���?�6*�f����%4Xp�`�^5%Tu��������O���O�˓<���둔�D�D�$�j%
݋Eh��#eg�:�6�O@�$�<����?�e��l�'C׾�A��8����D�-m�ß(�I[y�"��c�����$�k���w| ����->uc�OB�GΛ�^�h�I˟Xb!�.§�nZ�M8��A0fڎh�Pӫ�1�v7-�<��́�2��Fi�~���jT����BB$ �P{���XV�G�nқV�'!�� ��)��g�I%��e[E�S?0�l�e� 3wF7�+��xn��d��ߟ����?)�����I1f�L��"�1x~��gM��<@����4@�40���?�,O��8���Oh�Ӏ���3�X�`�^4�l�0��D��i��۟���6��7�M����?����?a�Ӻ#$(I p)ฑ��*K�=#�h�Ц����L��%�V�)��'�?!�$����5�Zwk×r^,�!�i�r�\h7��O����O��d m���O�59���4MҶ���<0���pT�D�%cs���Iǟx�	�����^��*�+Y�\���Ӵ!�V\Bq�O*>�b$��e�P�$�O��$�OP��O��	�d��a��B��#!a��F�C�b'	�L�	��<�����e��Fщش]��Q�Ci�>��%�d����4���i�B�'�2�'�W���ɐ{2��Jg���4��w�x��"Ɇ�X$�ߴ�?�aǐ�?���?��s8L��i�'�4]i�P?ǲ��nE�T8�w�a�����O��d�<���Z�|j���~��Ěq�^7�J�`6v]�p.�,`\�v�'R�'R���7��O��$�O2�iϸ-i��#�%ypR��4�N6zI�am��� �'u��[=���jy��M� V@C�&ʯ;���z�G�h�کd�i�b�'�<tQt�Z�$�O���ꟺ���O�AAM�O��9�ʜ���aF�ZW}b��M�o�O��d�<ͧ���S�<�4m8>}���̃:kX7�R%e��lğ��	؟h���?E�I՟���>O�}*�aЙD��P��2-@���44��2���?Q.O��,�i�Od"G�b�K�-��VH��0�`�ߦ��	ߟ$�ɦ/a2,��4�?Q��?����?�;)Gf����#4#��QT!%3��m͟x�'��䣛����ON�$�Od�:R�Q%��h��C�8r6I���ئ��"�ZH��4�?��?Q�!Y�_?���1ݬ�cAW9kYL�d!In}B����yR�'H��'�2�'$�;R����Zf�8HF�˚�R@�į��M���?���?�t]?�'���ܻY�� �hڠjފAҦ�ߙR{��k�'���'C��'��O�:�5�k�)�'藦8�H���+|p�����%�I˟P�	�����myR�'M��:�O�4	x�m�.$��M����MI��ˠ'sӾ�D�O^�d�O����O�%��!�	ܟT����6)���f扉;qv���޵�M����?9����d�O*%y�3�<�ĺ���u�	�bN����$��m�����O����O.��6��Ӧ=��ҟ8���?�bRgYH�1�� l��������Mk�����O��yd;��$�<�禙���dq��â	�6���n��D�OQ�5 �a���d�	�?�S֟��5�=���AX�>�[��F<��D�O:� ���O�O�=��̕�	��"r�K�;�Tر��̝�M�g3%G��'~��'s�$�OA��'v"a:fqB5y�jE.����ǖq�X���4h��ua����ē�3�5�i럎�Z�$�̢��e0 �F�  ����������  ��4�?y��?q��?�;p|���7[:w����'�8[�,LlZ�h�'��������O��$�O����*o�d)z��P����	ʦa��t�� x�4�?����?����Q?��kM�%g4u"�.E$>M\Tȶ�I}��!l+��'�"�'C�'/�ɹnZ���n���
7�P'��n�П8�Iɟ�����)�<1�x APJ7a��Ԋ]����5��<����?q��?y��?��M��T��i	J�r�d]�k� � H�87��ցp�v�$�O����O8���<��KiL@ϧ �(���;|�T�m��W�Ա ׽ir��'tR�'��	�<I
�N|���Ab3�K'Z�p�Ĩ��/����'��'^��'�n�џ'�����kWES�7����N� �n۟���byF�I���n��̻R�̒p֩ɇ��c�* `�.�M�	��P�	A����	z�~��
9A�>��t �O,-����E�'�
�b q���O�R�O��(Z�K5�M�iNTY�+şf�Ȥo럴��;m���IX�)��a\���2��a{�d��HJ�b�|7�ŋAڜm�ٟ8�����S%�ē�?�b߯XΒ�#'Y+�S&ۻ9���U6�yB�|����O9c�G��
T�6��)@��'�Hʦ��	�����3%�D�RI<����?i�'�tz�
Wi9��	����;��4��,.x9�S�T�'`�۟�|ì�3}Ent��.^��QƱic�E�F&O����O�Ok�^�#�|�C&�WF�֥�g\3V�I�e�IPy�'�B�'@��pQ��pb��W��E�C+%��`��
����?1��䓅?9�;]J��k،M��@D�gz�86� �?�,O��d�O�$�<'�R���iW)tRdݲ$�Ĥy"D��g�?`Ɖ'�|r�'�2#�y�N�?T�"���	kb�
E戄9��7��O��D�O���s�4���d7��O��D
�{Z4S���s?�Tj�L7���nӟ�&���Iӟp0d��۟<�O�$:T԰`0��
X��Q�7�i���'��I�{@2�1J|�����Td�|%�|����1aB|,DƔ�l��'�"�'�2����'tɧ�	W���)�@0��b�e@�]��fS���R̔'�MۇX?q���?���O t�7��K��R!@	kR��!r�i�r�'s,��B�'Cɧ�O9� ��E�X�H 1D.Y� XZH��4��Q&�x�x��AB�0<���ټ��+�-mZ��ඣEx�<9e�@%A�D���ݥC�p�`��5Z$��O��D���R�4�E/i���1�ګ_�f�Y��?NWt�"��w�b�x���O^aCR�;T;�������0[7f=2!`�t���c�t0�-�9dr.���
� M��Gw�\����[�h��b����tU��i�<�.�D�O��D�ON��;�?����Tć�(!!�Q� S����E�+������Zu##cV^<Z��㉎A� �(�;�F#w<L��֯�*w���rϓ�#���T��i�"y�$쏌��#<����+dy�l�CGY�!���w�Q*%8�I���F{r���->V\�f¢�%fg��a|��|�U-D<�|���V�6Ps�[���'��7��O�;g$ 6W?9���M��xDߞ�$��
�2�^���Ο|�������I�|���
�\��(C��^�q�4А:6�Njr�U�7�p��ɐ)��R��4R�d�	�4�ze��bV�M	��`��!(����?i_�5��"nvT`A�,?Q�/A��$�IUyҍ�L�}�a� �(���)��;��'��{��b��(g猒\���bf�
��Ol�n�+	� ɪF�؂^K����Ó  ���jy2d7w ��?�(��=����O�)U�ؐiE�t`0cJ�f`�Bo�OL�N�1G�<�'��/?�\�H�ɟ�'��� &�Kb���Fq�����.^���E�>����j�Ra�v���H%ހ���H��@�����̽_��40�	՟�F�t�'P��b�I�F����J�9J�f��'�21�G*β�P$�<ƖER�CՑ�l&�3n�̝1�Ɵ�{Q��
��M{���?��A��q����?���?��ӼTɊ�6ޅiC�~�(��Ğz�t,yA�E?Yb���7e4�|&�܈���7�V�����XD<�@�ߐ"e"�a��������[�q��'R��E	�J<,��/Q�N�h|B��a��,o�ǟ�[D����>��?Q2�
;Υ0O���Ab����x"}[��S,�F�G(,���JX�'�<5�����B?l��'��5l�Ν��m=1��M�c��!G����OT���O�ͯ��?9���Dɂ�[(���p��8o
�"�3'*���b�291ޭ� ]�%�y��)s8�PԊR;��Q�HZ.�mDހr�h�JkP�]��y2�ހH�+�� Chl�c�R8랴��Wa 	;I���#۫U�uɥ�-�y2%�[�����8Q%��ң�´Ә'�
c�h�B�U2�M����?)�&]�I?X��g��
v���!5I�"�?���Ԙ ���?q�Ok�yc�n�B�`8�G�>5n61ч"ɘ������l	Fk_�$џt��,_2�椱�G�0J�Z<p���<*R>��o vѳ׮ܚ5� �r��3[�,#<iv����ߴvl���':�T�'��Nl�P�d�C��j*�֟��?E�t��-�)1���&C����E�2�O��=�'8�viK�ssl���X%��$J"��7��P��R2��M����?Q,�����O���q�Ul�H��t+Y=m@�%��O������Z��BT)~����Z�h�'�����0�,�+Uv����Ez�/8r|�5�͖��\��EO�"���C�'�ӗ�.!C�LN'/ǘ�{�D�-N��'Y�1)�E�ɧ�O]�ˡ O!lq�5��B�-}�P�'��U+� @��=��/�.v�2�)�i>)�����9��8�s�X�0%0�.�(|���'�b�'XV�a�mk��'l���y��@ uh�Q���J�I�LP"��3Ԡ�"<�ܘ���r�ԁ���i<��O�I^�@�	��e1`<��h	5\? �'��0�JU%F	n�P���))���D�\�菓 '�!k�̎�<�
���O��D]2fː��Y����#bF.}*b@u�J��n%�@i�Ɠ'��PЋO[��(##���'`H#=	�'�?�)O�� ��6-�ʷ�2�N���K��j��1��O��D�O��$������?��O�K�%�4����G	�?\I�JQ�V[� K��Q:4(2ŕ}8�p0���+0���-��n���Behٍ �|+q"5�"�S�)7T�\I�B�+ B�"<AEDU���xՠ^� � yL[�o����?	���!�z-ZV���裎�~��$�̲�o��%�qRPGͬ��@�!3�	�MI>Q���/���'�rΊ�V�`�pc�\2Z����a��-���'" Hc�'<��(P#Pl�1#R�p�k�3<�t�B%�
1X��
ZuB����3c����bR5�|i�lQ�0,���G�=4�M��@Z

��	�E̡}j�=�u�П���4q雖�' ��s���d�ȱ�@3	�!�P�8�IN�S�O9�٩ ,��;*8�d�|"�[�'� 6mA-W�lp��)D !b)�ٌ֮���'�剋U�r���O��ģ|zp�V�?yQn�%P?~��5�F�Z��K&+_�?�S$�Сf�[�_��mZ�����dZ>!�O�&�[�"� �	ö�)V���J���KS
B��t
�cAK��KP��V���X�-`�t��^���	4j�6p�4 ʽ��I�7l:�d�֦���4�?���4(]<p��lK��.�HL����'�R�'�`Q�� �&u��M3>�!kÓߑ����
]�B,SW�ʍ9��DB"���M;���?��nԘ��X9�?����?�����C��ԧu�V� R�[#P���s!�!#�
-#D��
�Z�8�G7~�!K��tAP*�ΓX�@���^�fJZ�BC�\N�q�VЊ�4��T����5���Uܧi��ps��g����@��a1����ē(����V(F�������)�3��Á^�!JW�ֳ��M	���<!�D	�<�1�����\�p�>�d�O��Fz�O}�'�� Ue�)j{�<c�DX�R��gÕ�TS0]��'z��'&rDu����ݟ`̧v�u*e#[? �X(S͟?Eba4c��e6�I2�/�*"����',O���
#���A� �}�QpD��-L401���	`�2��� �~��%I�Ď
3�6=)��M�}h��fB�p�G�#�*nN���5��O��4���O&��1���N3�I��%�H��%����]FB�I:��$j��f�ą�#f��&'"b�xJܴ�?�.OtY0n��	�(І��i3R�]�,����Q���,��A
����'<�pyX�fؕ�>M�OD��h�#te�F
�'J�K��'�"x��}���	WY�� �� �)�)"�
���h��"
!�'�� ���{ܛ֮�>�sJ�(dv]����I]B�6���<���?y���%y��W=J�PF$�/H2!�DJڦ��@�2`������g�ld���̔'V��Ѱe�>����򩒫'�$�,U�N�i�%=�����q٘���Ob�h ��._$d50���b�F�=lni�Eº|��NE)z9���wІ�٣*�i��A$2�0�"��Y=C��a��'#h�S�)+��i�f����DɜG��X�E��8����i�I�M�1�i�b��RkՎ�R�� ��a�L��2�1O��$0<O�}�!�H�1�f2�&��.]����'��"=�N_���z��R!#�(�Z�AH���'��'C�a��"��'&2�'�׊L��ꀈ�.5zR���K��9��Eɧ�7�z ;@��E�\������G?�d�&Y�KsH��SH�X�g냅��D��
�6��n]%������K�~��P��揥�y��ˊ
�f!3*��DWg�6mUGybIX�?�}�	ɟX�I�l
L9�C�T/���Ȇ��>_��P'����	$ߖ��a�F�BU��+2����� �۴Cۛ&�|��OT�dP��+Fm$��4� �=[.���r��b�����X���p�ɀ�u��'���'�L�+_(�ؠ] )�[�	Iy�`�:QF9�+A���M��"�e8��Q����nXp�� �dߎm�#���T�4;B�H	�ȁ�-Ԯ}�a��$�gF�}k2HB�C�vM�U%�qJȈ���֟�+ܴ|����'��I��P�?T�����rA�ٯ�����F��<A	ϓ��+xM�)��b�F�"m�@!�J>Q�GĢL����|�b�a�i�m�u�NR�4e����$� ��I0D�Ј��N9c����ѬdE�Y�L-D���bILS�<����J�r���`!+!D��9S�R/p����.G�p(8�!D�|r3͐'��"FL_4@B����*D��ʷF�.%�ju!$�#�x8�"�3D��w��(Q��e3a�׉)��Q�-3D�,��,�N�<iF�ԉS:���4.D�����.>\�{�oR�l����#1D� #�E�7�N�IfG\6^Y��1o1D�\ɑhK�90Px�٧hgZ�"�*1D��ҤI
"vIP���.�,�6�KS&0D���j
500����b�.1��/D�����Ø4*��2�,l�58ǯ-D��1� �6&�)��I
UG�)�*D�h�!��0��L�fh�5�~r�$D��*֮V-E�L�	4���IUN��y��T	|s��L�Y�8r���7�yR�vJ]��,�Y���U�H,�y�(���PzKְX� #�&��y�*�7,�R5+���>M+>D:ed��ybL�0�`��	8L��Y$!��y"&CRJp�g���8\L�JΈ��y�@�����`�ȧ*�9�`h���y2	��28����r��A�����y�L��C��tbwc�8&�`C��,�y"��E�����C���C��'�Py��Di�}P��%�,�Eˉ�<i�)��&�v$fG� R�PC��e�<y��٘w'T��DS-傐��u�<YQdJb��<
A
ȖK�u�s�<9V��Y
�I�4-Է^/�A����v��lKu��I��)4�heZ#	ݛo�(�Oڡ��C�\z�$)�	�rd��:*YQB�㞼I��j�S�%;�B���i����U%)�듥p?�3)��vԊ��V�M8e�l2���c�`��Iƣ�0��a�'�(4ql�����bE��G����'	�����&�j׉�,GC����(J�l �O�}#c)Ap='��'m�d���W�m�D}� �@ "_<4D{�H��M��#͖*�TB`( q}bB��}Ժ��6G�0���O��3B�{�h���?~7�*{��6PN�c����_sr�Q�UO�hɆ}��Ar����dF�j4�Ȁ%ɐo4I���i��	7�Y2�ҲpeX���G
 n����sk�`,,	S�պڰ=	f͍^}�kT9��႔��6��[w�G?)�ty���M�? �=е�W&c�xh3�YdABe���'H��Ȅk]�gz��s���4�`5�@EĴ h��+7,O6�hb���)����#Ga�NQ(�(:����WCc&�����r�'ƖI�-?�䩇��S�rhi�'���2i0B0��6�o�veYG�;�db_��ȶ�>�&lB��rV�O�0�a;��Y1�,N 
��6�i�2!� K��
@	#0Q�}c2'�f����f(I�<�OV��ɋ�M���bD�29���؀cU:��۰��������a�&���4Ps�W��p��rN�	Ÿу�	݌W��ٚ'g��طvv����.~�w
ϻ(4���������0��>0�r(bT �>g������2����'��	����' �;���$�ؔӓD(�@�6D���Xx��؋]�����#ғ;0AX�h�<4����C�ՎC�h���	�a��L��)K�{G�Ey��>Kϐ��x��G�=� �E��i�>d�r���uה|���B���ZGJ�!Cm<x:2m���Ms�Ȩ>+Ȩ;b��'Ǧ�4'S���������韛V�܀4P�X���>� p�*��Jm�Uj8�t�QA�����k����3��2K*�sa�A�\�f���4s�F8o��f�ܘr�O�3�,h	��ˡ������6���K�.!�O��H��'>�U!�]��dYR"��y�ث�'m�@�e��o?�p���@�|��T�9d)��{�O���ǟB$���ɿ��A�*N�s�
-q�O��wQ�p�!I�<$�D$�'��D��9Ȣ�JpFB�e�����&�4N�$O��
^��湨C�-=Uj	�w鉜C�V�'@�7s\U��Ȇ�j5���TEb���4S}����9c���AEv�H1ѯ��+��И7�'ƨ����9�(;�H�s����4|z�9�G*�>%'�Wj^�12�PG|�KϘp��WV�F�t\+uA�9���94.LK(<��
O,l4�R1e�HZ�j���<{)��ƞxҐx�?O"j!���s�.٨I�����z0)sg�(_a}�&޾sо%�(�s�	z6�\��y��_/@�ؒO.�I  ؑ�3���'sȴR��*!��MW�m�&�±,�ּ���DPZ��Gz�%͆kQ6xc�H���P�e*���ɹoD(��e+�5q��x!��dО��B��6�X�G�70^�H
Ǔ{E
��W�!g!��+Bŉ;�楻S���:�Pp*y������hO�i#9�6��R�U�/�чV�
L&1��J���L�N�i`F̉v�<�`E�\A�a|�!
fj	R.N#g���w�J�S(Bɱ�}e$qҌ���;��@B��5��)'���
�V�
�^~d%�fZ9d\�� !Ӥ��'� e�0��5d=��H�)ݔZ�ȹM�NU�%Ä�^�1(��XsnK�^��<tB�C�Fֺ3�r��4/R�jt�`Dzr�S1l���D�Еz�tyjf�Фh8��≬ �\��A��&�L�
Ó6h~�5�M�W�ޖ(d ���hX;t�֌�.ۋ��>I�k�F�l�Q5
�4j��Ca̋t8V �����Ą��y��G�0d��a%��R�'̉'���3�Be��х	Q �їew�i�n\*�0<��1?�-�'�_�6cRp�Ɓ�$E&R��Qf@
-QN�4p��Ex��=}
L��ѫ�b *X�*�����j�Pxs�ހ-�Ll"�͏_��ɝA�$��@j	�_?�|ZD%�:Jon"<���Bhxΐ��%0O�0 B<,�(����9߲���A,C�4��Y�U�����0���#���5Ԛ[�i��!NܧO�O�-�<�`"R�ab�9"�LC��ap'%D<J�"���w�x�#�Z�B�d�K��V>�%@���RW����]"T�x�!�+����ɢ��<c��T#C%�ax�G=}w����ǀ�MSf&��Wz�<�ҎI�RP���֏< �q!��s≍�Mϕ���ֆY��P���n��'�,��i�.��;�.�d(BI�Zs
L���R��'�<�Q��M��<�'i�x�H`�#�j|���A�l��t4�G�D�l!3���9����XW8� R�F�Y~t�f��:�yI��I!b%j��'o��҅�{�ʧZ,�>�Kv*ִ��; /
�e�rH�2�
�$'�}2���b*�j�s�8��9����!L�>QÉ���̣��.!��Oj�'�V�1#�E4
ǐ@)�F�a�䰘��A�'�XE�t��l��G�I��Ӏ"=6�#���40��;􇆘@>�*�k�<�W��?Zb���OsȨ��l�,O�͂�bH7e@lk�f^s3��Y�>O�%rWԖF��423���ek��$>��|��(H�!�B�M4GY�,"�L"M�@��o��Eq���2`"���በ��|(�,R���aR�A���eۧB� ���)/�&d(O�2�' ,� �� @��P�� �����*�0>d��ϼs�B�D�z��/��k�托��+7:�I�M�#jN++,��'��]+�tA
ª4NC�LJАg�Y9qȣ�hOR�(��0hF7m�����a�Za��o_�\-�d�4�%�p��!ڈp�t�ъ<�dS�Q���ϧ,���,�9��	J��+4���p!٤c	Yr���㺁��O���!/5�?i��
�����>�d!G�6�F Sc$V.P�I�g�
�riwgu��A`�
E��v����<��l	���5��$+ƦL�L·�ٶ�?��iO��M�h%�T>�	ަ�H�윳8P}��#~�3P�tJ�����/3�
��{�? p�T�XB��C���ٳ
�y��G����>���1���������h±GT�J�,'N(Cp�D�����`ґԛ�dI>��-�5Z H`ѧ�L��Њ��5Q����'�Te��T�VD
1sSZ�\*�O�U�EIA�-Ǽ����$.;�geO�5�v�(�y�k.1��'xI�N��0 �R�0�R�A�-#hU�U��@�r�$3n�5�6�F��x� [�dɄ� c+S�w�| �A�͗���IJ<�i�#<!�^�<����252�Yv�+<�Ssf��a{�钧1�΍��%��!Ǉt㶴1��
=�z�:R�\
�r��d�>=f�r6�`��G_�\����`� &�I�a�I,s0M˧'M�<1��\0Sd$�܂ݓc����)T�rV�R�B>�*X�y�%�y��-.KB�)c�/?���F	���g$Ҁu��!4ڦ�@� �;=z�E�4C�ÃNFH�����d5P�L��E��sa���@�1�DF#5O�9Y@Fp�����4O�<+�f��2���3�ߧ}�D�0�ړr�&�OE��I#:���抭���`�^�p�4�w�'�,���%�%���c���E���[cF>5kZ!RD!��?&8��DݺP
����X`k��b=4�rE��|yw#
�OnE�g��uEzi���}�P�����Æ
���Y1�HsV���'23�E�5x�P��"j��pf�q�'� ���%]n�1����2(0� )>|Q��oѸ��$�As��N}2�>�g�S�+�:�ˀ�L3K8�%�� �":�84�v�ӜL��5��O�*�R��M!<R�p5(� 5�x�� N��'-O)r	P/Od��\4V��Z(!A�!Mla��t�L��>�p�w�,�� ���BL a��-��eR�'R
��A$�H�`����s�hU��8��s֢\��O|�iC�
 N�X�2O��Ve����i�����UT`��s)r��:��䀞g
��-��g*�����(d�I�j(܍`�HG"B+TK�O����XE�jӴ�z��M�*�܌b-O���O�lR�(�J�4�p�x�s�Cʿ'�6�X�8�5��8�%��s�3d̕�4���O��pM���F\ȒI^S~¯�M~J?�n�Vl[��S%�|[NW���a�V��`cfީ�T��P����ČSdE�%�v�
}��OL#>�u���6D�P���̠�uL|��A�0�L��V��"�9>�(@�GMh敫�*ڊTФ�ɪi���P%T�UF��r ��+���r�h��S(��A�Z�+�])�,}r�G�C���옻%砜�ǯĸ�y��ݐmL��Yv�)>|J�)q�W���O��@���EO�ɪ@�7Am�U�fj�*$��[����J4<qЎL�/&ax�h�N�l����$X��h	�!V*H����9�0<1 �x"�ҮIϨys���B��00Oð{B*��MC��;"�bu�rb*U�4i�4>�lA#2��_��'�ZA� �'P���mS-)ǐ����al��6�Ǐ?Ha{)�Q����نҎ`�pkW1-�������!o��,���Ov�O�-���&N7v���99��b�>���z�0��-�9)s�@J6�DV�I���?P�`2�K�3��	�OT�c�ϟ�n�t����H��h�L&x���A��;~p}��Y�vIaxңC'^�t�s	ȔD���c�ؑc�:es�Y�x��MK�Z�y&�L�\�'��ənnB`��/WL4P���7L�j���.4�l�������g�'b_�m[���6��ɜDQ���[�-���1TUȼX �B2 Mɵ K�1M��B�'9a4��(�D�f-°����S��
�C�J���O��N�*��ҬI�p�4}�\w7��>�O݇P'�yᢀ٢m�*�A �P�J;`J4�R5��&�7ELʧa���ߵ)�F���lX*��pCB�Z&�\�VfԿ~N����D-w�t��	ǓqW�劆�˿Q��9H� 'CF
s-M�(���e!��T�RqlZ���i�<1`\?���%�&+�������N�@�1�C@<�B�	=t�dh6J��B��{U���C���A�#Q�&#��)P#>��4�E�J��_�u��0+l��r��ڦ]}6Q�c�֌��=ٰ��&j�l٘U�K�!�+�L v��12!?�V����4c�bA�'dY �	)�Db�3?1��	9'�`8�a#C���*b�v�ś��'g䜉�����L�Xe$>�Su���ə�J)�H��G>�Йn�ys��	����$B�i������[H��#�
�T��	27�DD5��S�Ov��dL�:E�X��@��P�4���'T�$�`�+�0�,�B&�X�{��2\O�%�4�شq7Ԍ�4ċ�g�ڱ@B"O�zs��,cx.$1f�ǙMVm�"O�	j0�B/��M��/ێ���*OB�+�lC=�
��=9�9��'rD�Q��!AC�D&���D��'��yx
<S����E���>+�t�'=P��¹1O�����C/r��B��� Zܐt�'i� ([$	S&^X|)��"O�$!�/Z�>�ó(�9rM��
�"O4m	� �+���&;B��3�"O\�ڤ�Rru��b��GR�Ȋ0"O"��!�+I��Q��
�xO"O��W&�9�<9��-ԟG0V-�"Op
��H� �p�u�y��ͫ6"O(Ҷk�=�p�A��2V��g"O(QeO���]@�Q=TxX�"O�L�0c� ��q�`	�l��E	�"O��5��jYyR/ޙt�8�#�"OʑR �~AL͢��95�>( �"O�%pE�(��K 
��i��"O�Ht��$�|���� �p���"Of��'��!U��I���63�D)�"O��!t�֚a��p��%{��-I�"O65z5G�%�&)y2�)w�
��"O�y�jJ�r�0�Ǐ�	O��)s6"O��w���Lh�;o�� �B"O\(���?;p��H�fս)qL�"OuJ�\�zPj�^b4q��"O��_�=Ef�"�ȁ-FJda"O�ͱ痡v햀�ѡͫj)�v"O�H���<܈�)�oM0��7"O
%�5�ۈ9x@Y�bn��F:�"O�d�G�]88��;���o���Ѥ"O(<�cj�A2�9k4$� ��"O��)h�-S��1�Ä 7 ����5"OI��.5*��1���GfL�A�"O@�#oȎrHu�L�����H�<9�cӦX��9����d��PDWA�<��bŵL=.�#b��|	��GTF�<�a� C�
8�W^�W�Ve���F�<�d��"�R����Ըn��"tF�I�<���2-&�$zFHt���x��ED�<�#�Q� zބ���r��(�E�@�<�D��1E�����%fp��AB�}�<i��Q�� P� ���
�N�<i�l[]��q�\�#��ِ���s�<�t��AV* �.K��0G�Or�<���\*��T��=U�4Q��q�<�2A�"G9�q���;4�"(2B�i�<A�B�LA�-�*R�Y���c�	O�<�V�З� ���i�/K(�P6C�O�<GfN)f�j�� �2�1��AJN�<�TB6L���:0��(�*CP�<9�m�4x\`�@s�5.^�}�pI�K�<	��Z�f#U��&!v�b�G]�<���TYH-��j�"+�{�c�M�<�"��&�B¨�>@�+W�P�<y�
_�<)te��:��s`�O�<�ЋV8x>i���Γ(N�D����L�<�r^�v��� �ǐM�<��N�~�<�4C���D=�p%�}�n :��D{�<�s�)9w`i��d�3/��5ct�<1�\�(~P�9�N�H-*�
��s�<�pM�al�Y�n5%���dj�<I��Í?_H�h6���|��]2�LDe�<�pIA�V�N`�F*-J���&�x�<i����j���
Dn¢4d��Â-�O�<y��ÝY�>hQ�-��3AK�M�<�(@>05�أ�B,
��y���#D��rK�8⾀q��A#`~ O �=1�#�;5��Q�������X�<� �8���Ξd�����4=��
"O���'�	T\>��OZ� 7ƀ�1"O���u�È+%���	��%S"Oz���FBHD���Dj�iu"O��c!^A�,�@���
�p���"On�:`g��Jwʥ���W1��A�""O ���4D)��9쑛_\Ƥs�"O�m���۱Y.�K�*݉3W��(�"O��a2�ʊ&����`˃�N��E�%"ODhC"'[W|JS��=p,�AK�"O�8��ӟ	����/ɕg�S�"O�H��֕9��l[W�&x�$1[�"O؀2`�:� ���lr�	C"O~�R$�\!z�d���7,=0p�"O^͡��+:8��6�E�!��[@"O�� ��"
в���*ߵU� I!"OJ�Z��D'9,��C���^��e�Itx��q`n�F�z7���)V8Y��-3D�|��!�����u\��M��1D���щ #	(�2F��|���5�<D�������@q�h�� �?c˺��ҭ&D����':W���F��kD�!�G$D�<�.D*i:���eDs�@$D��;W�F���i�'#_����CV� D�X���°2��S�h9g.�)*5�+D�\c�Ҙ>��%S�O�y�P�*D�p���֏R�n�aT��x�
(,O�<!�+�� ;�)r���]Zr]�S��Q�<�3��5#U��e�\�$�\q��
�hO?�	/|@��hʗn�h{0��}
B�Ʉ)o:�Q��J$N���kK�A��C�I/2��PAM�>2�
6��$خ�'d�Ey����N�w��l!�ˇx������y��BW�
tЀ�< �@��'mўb>�CȒ �>��4c�gO�`Ն%�O:6�c�l��#iɄh�|m�׎����a��T����bn*"�N��e[+{��q��,�y¥8Ι��Ë4_�8ѭ�fI`b����0W �K!&_�c�\���(�O�xC�I��"�H�'��x7ji)��X$,7�B�ɑ[� � ߣ0`��0�PnsxB�	�4�ڥ��$~.�� �eв�B�I�n�"!�,��%�~s�ό[wB���,uȧ@�v��Y�����@�$B�	#���	u�O��'�-�
B�	.8y�͜Q��Y9��	�s��C�	f�Zd�Baŕuꦁ���Ȑb:.B�ɶ���ѭ�,vޞ�C%��	��B��&V�̒��P)�0�1��ϫj��B�	N�v��v�#L �σ�zB�I8&1�����C�v�,���͌�w�,B�ɉ*���S��C3�P�wHL�qn�B䉽��	R�ы6��e�ˠ7̎B�	
�<�s�Od�<�re�� vB�I=s(����n� !}l3!F;P�C�I�9�a��(I��� ��-ut B�I_�V�2��V��a{���0v2B�	!1� ��Ǯ2')J}�W�D�t! B�I=L\(8�3m��
|
)J́@~�B�ɵ6:�Ls2΄�'��Qb�@�B�	�"��[�A,���k)C��B�ɃY~r��dH��*��� xz
�'#�i�e'҅&Gh�/U�IWv��
�'�><2q*��#���9 _�3ipQ�O�=E�� x:�o�!5.�)��!��1A#"O�t���[�%X�q���0}�8���I\X��BX�>.z�"`��9z0��& &D�x#eP�I8Th�DS)zVQ
1-8D�<���Xi`Ё�˄%��a���5D���s�C=G("`�6�֫@b"D'>D����E)3"L`��'�E�epW�;D���s&ȵ|�!؄��d��P{�$5D�l!�Տt��XQ��k�	x�� �d �O&�r�C�A}�-��O�4��Y��"O�#��ÖT
���͕�U�읈e"OLM�5��-��Ҷ�\�r� �"O����懿K��݃�#2����"Oj�P�K��$N1�DĀ'V(��&"O�\��S%~'�ܰ'��>
���Z�"O�" L��nvX�G�@�:8�QP<O8��$�rTv���	�
��p
�a�!�D�*k�Q�'�`� [#GD��!���h��H�?C�������
 �!���:ᦩ:ah�Z�49�vo� !�!�ď�()��"ʯnkv,5/�-s!�D�wC$�x-��Q�Z�(�^�N_!�01��yb�àz���Wb�!�+F6���g�������ȷ�PyBEԾ�Z��
�.G�>�[%cҴ�y�/�]zf����ɼ:0TM	��=�y�o߷7�
Vk&mV�BD��.�yr@�:��!�uF\-H5 %DJ����dX�,"A�_��H��/O)=��2�"*D��Qr��R�h�R�$����BG-D�43cC�%�X��6%P�?�P0 ��)�O��'d$jW�:-�H����w7��	�'p�8��IK!�8:���lٲ� �'��XۀDޠ\�c�C��i�d��
�'wV�P���2�xx����)8���'ٺ���)9� h �B�".!pLy�'�pUQf���>�XFß4�lx��'��9�ڱ=%�|��)z`H��'� yZum����L)�i�&���z	�'n�b��/C�8����t��(�'M���Mձ5�vDB7���jI���'�����h	5p�������b�Ly�'HZ�#���#	�*�R�#d�b�'Tm��g/8��p��MH����']T�E��j8� *�2G2���'�.��®�-K~�@�U�?�ny��'��}٢��/#�]�GÌ�'����'�(�T��Q��ȁ�)B�`�'ez��r�ݹ߅>+"��1����yr���:�j4Ч��!�f��aH��yRM�+H������~`�IK�y"F*z��0A�D�a*V=�y�
э;�2��@�9I|�kaF�+�yb��Z�H	���40�X�B�F��y�!�%=z4�G�O%*N�JA�߯�y�AR�=��13�*	��p ��y"oͮe�e��\��*�8�J��y�(ƧDxT�a
�&&�����2�y��U#yn�7�=�n�����y"c��d,��ڐ'�Ǯ�"V�B��y�^9'��m�X"T �5���yR�P��|K"Ip%�"dT9&1���ǄV鞽CcAf�����L0!�L�T��ݐw�,�艕͑�.!�� &pвiX9
��,q��GB����"OL�B�7U|�ѧ�R*4��5:�"On]0����D� ���T�8�J�y$"O�H��?k�bTP�/��6�6���"O��"DOy�t�C�nH4)�(Y�"O0]��iؓMG�2!/�t����"O&�t�G/&\��$C�zxkr"O)h
V�/e|���ҟ(b(���"O�8X���m����T���e���y�Qgf8ɷ��0ArU���А�y��*G�e�BJ��Vm�b۰�yb��;X;�p
��]~�D�DR.�yB�ƺٮdj��_�#���a�y"�U�g���YwfK�G^�A�B��y"fG<m�`��R�mYH0�;�y�hA�'��*� ը;D�4�e��y2k@�b��fL&N�q��/�y2��>S�Ta�a�!J!��I���y"dXr��1A'ˢ@�0!y��2�y�-�K�*Ur��3$V��a���yr�݀a��ȲBm��,}n�kF���y�A��\=sZ��~<�����y�e��~t�M�>Z.�{d׊�yr.'�FQ�Se�?=�\��˩�y�k�/%���4֠�ӥ(���yU�y�M�=��mke��y��čD݂�8DȆ���QEOI��yB��=�.�9f�H*zt[��0�yb�X:�n pH[�T㤠��(��y���$v�d���Q˚��bL�6�y�L�A�
�yR˖�5�&)� �� �y�e$H{"Y��Y'����4�yk@�E�m���0Q%<}!G��yr�݂:k�-��+E��!vO���y�(9@ƅ���Ì88�[�圴�y��4@hBIb�N�7N��	�ɋ�y�Յo�|�F�T�.�:��')Գ�y��E+#aT��� ۻ!�&E�Wd��y��-SF~8ȗ   �G�%�yRi�X"�;�B.e�m�a,��yRoS-� � Iц9b��  �y�N[�f)Dd&l��97��uŨ�yBG�|�.qJ���8�6������y�̜sݰQY��Ǘe��e���L��y���b���)��X�
�R@➶�y��I��˵aŴJG���
��yB�Z$j<��(T%�-�"�
�#"�y�*�����
��0����ȱ�y�&�	�QM�)/�JQX���.�yb��	��+F��"Ԏ�͂��y�@ɪmv�*7��	BD�Dx�g���y�G)����M-39������y2���h�r'���+����⍤�y2��fA�V�A�N��0�iӪ�yB��9^�V��T�B��
�� �y�NÏ[W���5d׆.�xf�,�y°y�y*I�B���2�"\	23!�J�@X$T��#�u}�B��!�dKy5A���]t��FAJ�!�D�/$�I�l�<������!��H+J��� پ(ވ���N73�!��,�6�Y��_.p������!򄘰
�(�k3�w���ӬW�!���v3aز�M�e�^$��K�,#�!�� P�@G�PRd�(p։�@���"O�E�C�ݬ[����+R�?Kp���"Ot�j��'h抉H�--X"�K�"O\` ԨK������N�>p�����"O�SF�������/��	�:�"OPDv���	ݸ�sT~q:9B7"O�ɰ��
OꍁƉ�!fl���"Ob9!bJ/a�
���O�M^��X�"O
���r`0��ѣDQ�x)"O��Ywj�[8:H� eܑ~@J"�"O��3D�F#l���X�I����@"O���dg�'n���ᛙH�ܴ�"O���K��'�I����Z��!P"O�����<-��+C*S�"w����"OV�P�(���p% � �+c�U��"O,ah"�̞]���c!�
mK�U+�"O��9��Hw�p��dL]1���R"O��;���Z�
�A�h� F^\"O|�pG�T4E��3��'�Н+""O����F��8,ᱷ[5~��a�"O`X!l�=,�#�%�Wa���"Op5���E3B*eP��I;�0�!"O.�*C+Q?U\��4KZ�B�ߓ,!�D�G�<���.v�lb�V]	!�͍u.����F�I!�e�����!�Xa���i� a��92�b�2z!򤇁R�x� �	���  bD	u[!�?W����7o�����"(:!�E@�\왆�;��b'>.!��T0�l4	�G�~��T _��!��{K��z��O��((��_6�!���SE�\S
�x�5@�6rE!�ͿB���"k�|��	�m�Gb!�ÿy��r1$^)o���v�АnG��]�+`�$[���A������yb L�b0HBƄ�1�=Uͱ�y�⟅O*�(��@�=#����T�H)�y)G�9Nz��	�*��	��*���yR���|����ˁ��.-��W��Py2�F�Fʘ��Pj� ei�b�d�<�͟�e���FJ	?A�*�^�<�g�'Aa�Y��Z�2ĄT�mc�<y愸""�1��H3L��tQ��W�<�Q����{��J�m�ڜ @*��<�FOf��G=��\���Gw�||�ȓ|c�2�֘��#C(9�N�3�'O X!��u|\�hU-{u�8��']�Q�a� O����7��yP:��
�'ώT 	?u$"��#�O�s2���
�'k��c��,���9CD��p�"��
�'t -h����"�P�_X��	�'���R��Y�*��DM\���	1	�''X}�wVrF�3���=4S�E1�'.85��E��;�)����'�ty�G�Цs����w�S�%���k�'sv��Θ?z�C�%�1��	�'�&m�G��tT�iC�c]��8$��'�X���i\�V���E� Gb��'P`� +��>�遢�	p~X�'~�03O�_�,��P�@f��hr�'P���W�	�`��e�f�r�'��p��B6���Kȵ%WL��',!!�kBTĈp�Gj=ѣpo)D� �$ P�l��LT.DÕ�&D�� h�h�3�:L� �Ăq��h@1"O��@�^7.6�dlAY�d�	�"O,�x��.�.�8l	�K�Ҵ�""Of9� L0�p�EkZ�D~����"O���T��9���x��`"O��*q�&Z�a�#�L!�dӒ"O�4(Ċ5V���U�7G����"O�[����U��+!K �\mҀ	"O�Q�'������P���L�.�i"O�jl_$mV�R%V�#�t0�D"O��	&�	�J��r��:F�B� �"O�#b+�Dk��3f����"O<�:�H&RR~D��i�����"O�p
"�ϥ"CҝB@U:f{0��"OR$�7�
P�}���k_��i�"O���Ô�k�B�CP�US(R�"O"�f�C�53v�c@`Xco2��"O��H��W�<��x� �VH���%"O@)@�:O��G�.0�x��"O�Uc�QzD A��V�m�aB�"O�a�����(袪��j1�Ȫ�"O.ݘ�'�1o�yҳ��"I���"O4A�&���]�Q;�A_�L*i"Oz�H�.��iS�b�D�NI"�"O��䄏Z� �ce@����w"OX�;� �2ڸ��3���	�t���"O݋r��O�H�֮B�nzL��@"O�� C��8}y�P�2�l��"O������4Q�X�g�ݰh���3"O�RA�� O���(��7&�^!	e"O�0��*1ĩg���+ "O8��˞#s�<I1gV�P�{�"O�]��dǬM������2n��5��"Oƭ���ؽK`x�����q�"O�Z�[����P�L��$�Lr�"OФ��)x|����!p�!v"OJ9C��I�X��C&B�dr��c"OB�٤�]��sg��
�,�yc"O�� #ٺ4\�-�Bŏ9+�l��d"On8���I�;*����\�^w�8k0"OH�x�F;��9�Dɝ.l�#�"O"h"�G&:PJdj��Xij�F"O��8ч_�"�ԋ�)�
0T,y��"O�M(p��7��Ir /�|d��"O�I�C@fN~�k���/N�"OR�� ��8�*�I�Nȇ �rB"O�)A�����U���]H"O�L&��c��ؐPcD
�<�6"O��a�(Azì��6F�-�3"O� �&(�Af��U�@c(��R"Oؠ�� U*��Rr�	H�th�6"O.I�.D%Bn��E@]��b�3�"OxmYÂ�1"�x[vOG9���"O��`FK1��A0uE�![�N�2"O�eB׏\?��t0���,y�|���"O�8��L�vjYj�b�:r����"O$	�סߖW1�,9��G>P��Q�"OJ�r3���#�"E�>��Ӓ"O��*�n]���	�@�Ћt^8�6"O��:VBV�)"T-���5W��
�"OpeX5��:p�$��O|!H@"O� ���we�Tp��D=�Y)R"O%��Sm�)��CD0w�x8t"O����\!>Vv�ձd�3F��y
� �]ےFH.<�*��P��w)��K"O��I�&�Ǩhy�@�]2��"O8�R"��c)DD��E�Y`�ܰ�"O8$�snN8N��*7�Ψn$��
q"O�0��L�	�T��ȁV=H��w"O��r�	?�$��NEA" h0q"O�� `hT'SD���m�� =�]#r"Op�1FH۰:�a��LF�ATn�03"O���"����Y7��'~\�]�"O"�A4b�?|���b�ƈ('f�$�"Oh�S��M��x�[�*Y8���"O�CcÆ�:�ҧ�Y+<��!"OH�J�*ٻG�6X�C �-l|�"O��hP�ȟ<���yB��\�,��"OzE@���3c�I�T�ė'H\�'"O�u��l:&HAap���v5�"Ox�	G��,4Z�c@>/�L�a"Oܭx����8\bԌ̥["�$��"Oj4�qCY�	`���d��[�2"OB}rp�C�T4z@�tLX�L0��rP"Op�8B�օQe�ͱ�j�1�����"O^�����<-�,iW)�'|>��@"OJ���A@�u]���bIép���f"O�L�LB��� �m	`��;�"O�S#'�v,�x�榖�1��"O�0��Ao�^�"�f¨!��-��"Oj�(��5%*9J�f�y����"O@�9V˓�n7����!�*x�V"OB�u�[��RA�Nу"k��#q"O�}��Ŀ�d�� ���(V�r�"O&��&)��ĠaEf47.y �"O8����q�\Ɉ���K�rH�5"O����Л?N�;��ں:D���"O\�J��߂`��x���>S���E"O���j��4Ĉ��'�E;>O�,��"O�]�S��]z��*�mV�[N�"d"O��� b��|ёLJ���"O��j# ͋a�RU1f�̀SN���"Op|3��!�4��v�S6&Q9`"Oz�ZR��<{#p�x���=}��i"O�I�׮��
��k�l4�D�٠"O(��r��b���3��Hּ�"O*���h{���F��~jy��"O�qJ�lX���D�*a��J1"OH���aT�o�Y�S�F�.��S"O �%� vb,M��
&�nx:�"O&�H��Ҭc	׭J�[f��1 "O�0��Y�Y"�5�*�lsV"Op,�@�Q@3��As��N?|Ly�"O��'�+B�����7T^�Q�"O89�H�+iK�����P;.l�"Op�C��;=�� ����(���x�"OH!&�G�KGl���#�:r"O�A��-�(t�qFN�m��#�"O����.V$0V��A	xѺE"OD���T�.�����ؽ���s"O�HJ򅐣?<Q-Au���ŗ��yB�U*�|ô��"(D�r�ߒ�yr�߭HD�`K"��)r��k��ݙ�y��̑H�H��@/���X�,�3�yR㜗z蠀!$�
�)3�i��y�*J�v�. E� /��a�����y�JȂ"���"��T,~[���1BX�y�/@.����S��@&va���N�y
� ������Z j��^�u,�D �"OL�/���%�&@�P$@a�q"O@y�!�MK���כM�tE�"O��ʒa 5`\������B�"O��JB��h@��/E�,2l`"O��HgCJ
2�`9[�D�rP=2"OШ�5�ɗq���0��
~Z&8�W"O԰��MG'Ds�p��)	6TT~i{G"Ond9@@̣r�X��(z��`+"O��Bv�ϷR���zGP����W"O֠A�W�\6��z�%�|�d1�"OZ%��B�	Q���х�t�t��"OB��a��2�.)s�	"T�(X"OB���)i�l%���Nfk 0ʶ"O���B"I'h���	1�W�\��@R"O�)b�cT�}O��{RB?J��"O,��r�8{���^�30��"Oԙ1݅/t�!w��d�����"OY1�e�=����#��3/��H��"O&�'��0�&�_8t�|�1"OH�PhR�a#�1"կ
C�(u"O`y�e�
d�`�K AD*2�؜��"O^m�q��'^�����՘{c�bs"O25��H�za>YP����}.F@Z0"Oҭ�C�:[d*Q�مW{��q"O���&�F��@Bo�hb-�4"O*-�&�[ղ�N��>`�A"O�x�UH�Ztf����eQ�Lh"O@�9�Jǋ���Qv�]'Qg�@(�"OQ� �Fy������i���`"O�s��$HE�R��e�8!�"O�H���
f�D���K���k"O�0r�H !��d0�'�;w���!"O�Tg�_#���2�c�|[&���"O��b��L6!m����K���~̛4"O.�q`�e�,���� KE<=��"O\��$��;i���%�t-c"O�AzTD��@,����O�W����"O�����I8!glX:�&�!8�ܰ �"OP%�C,^	az���Z�6D
�"O��r��ٓ#����6jES�� �"O�,aB������\�κuh�"O�d�r.�,�jD��΋Xf�"@"O0h��bS?`H�`g� F8�K"O�dA��t���ƆD�%"O^Q�W��^�ȠeN�o���!"OBU�$��kv@ۤC�p�.�x�"O@H��ś�Ym��)D�˽f�e�7"O��"�����i��
E@ԔX"O=��X;��&�X=G3�(�"O�Dj��6����d	��q"O�A�"���)�� �a�І"OhĒ��5<H�<����m�Hܓ0"O�1�N�,	3aW�G7l9��"O6$I I�?H��ɋ�ߌ$3�u!2"O����m$f�"M�ŎV
K�� "O�!W(�UOh��������"On��#
؝a�8��j:{���xa"O���S��#R�j}���M(m��3"O�I	!�QrH\�EE	�	���C"O����[�hd�u�L�f�<�j�"O�c��F�NZ2�C5Õm��2w"O�A ���Xԭ�w�B�uJ���"O~���-����+�??��0Z"O� �q8�YKɶ���oNS�ra+"OZ�	�ȍ�Km�����̪eP�e�"OV�QD�G%b�f�5hS�\��"O�h!�!��M�v웤8��;�"O�L;���6;UL��ę�'�-8�"O0�!�EQ	s��(�m��� Q��"Od-bAn�m�6Q ҫ�N�����"O歲tHִ{!6�)� ߧ	۸`�d"O`{�ĕ���A���E;J͸�"O��F̏0x���#�=A���s&"O�15��*�4��䓍o�|��"O<08�gȣi��2E._
��C"O��qDd]�Z�ҡ�O�.��زg"Ov���#S٤��U��-b��U*O6�Qa�J�I����S�#��8
�'�`���G�teU�m�L9�')z�!ׇ]w��s��E�IH��'P�%C�(�������=�`��'�8I�Иu�[�R)2��D��'���x��ۡ"\+�C����P�l%D���>����B�T�:�cs
���yb̗������h n��bg���y"怵vEh��&��xa&�3�y�c;k[� `��B�*"���y�(�-�N��t�#�tz����y)M)@��#U"��ɂ��=�y�bʛ2{��1��=%za{a)ם�yr�R@3�|)��$c��p���y�m�3z JEڗ�꘸e#��y�k�;%F�%^)IZt{���y��8L�islO�86�A"\��y�-B?)�֨��cG�/���c�%�y��Fgf��cm%*��C���y�JK(1� �ȴ&�d�cr$9�y�!� \Y����,� ��Y7Ε��y���T*�#Ђ�"nht�q�`T:�yb C �))��_�b�}�'E��yB��<B���a g��_�P��G-��y���G6��[`�������y��̻X��%�R� ���K��y"���(��[�蟰D8���ի�y�ў#"`��lR�;�� J,�y2hE>�£�Ҿ7`,�3��y�̕�0��X�q&Ŷ{��I)�h��yBӰ#�a:�$�w���+�.[$�yB�0�pə��Z� 9ٺ3·��y2�āi0İô�)����q���yr/� i�2�c�	X�
��I���ڐ�Py��_�t�v�z�jJ�E6����UB�<�t�]�%�Z��B�_:��5��F�<!�E1	9v�w�Ҡ9E�X�<9Į[�G���q��P�<�`2EDI�<t+�61`�`	��6����RV�<�g��4rj:3�}�|��F�x�<���z�Vx���$&X�ԸA�Eo�<y �N�%�i��!H�~F����i�<�P�wk�] 5/R"(�.̓�\�<��R<���a&V##�8�!�@O�<�1G��@۔1eB6)�P$*�HW�<Q`���|�sL/ּ���JBR�<�����b��'��8�H�w��L�<�wS�."���1���%��S�<i���"jɫ3 E�(����o�M�<���1@XzLА-�,nLtp'�F�<� �e���i� ��P�H޸�c�"Oj����"`�"�B�~��A "OV�sC�
}5�pH��;Xȴ�!c"O� CBJ��
��0���	��8@�"O���w�HP�Ƀ���+0q��"O<t�DÙnpu��"((�JU��"OH;J�1�X1�@'H�yD�"OԠ�n+<҂��׋�L��7"O���]<@�ZQ{�+�_6�1pT"Oبp#��@��m�֩ܕ*j��&"O���m�oL>����ӉK@���"O~|c��#*��BT��2����"O��Ѳ�T,�����Z:��v"O���Aۻ] ZX��J�`�Z�"�"O���bC�Nɪ�{4*ϳS�u�q"O ����p�̨�5J��p�;c"O��bb@��[^�(˖�A&-�Y8U"Oz��+@(�R��Lk���#"O$p�P�L��B���	�3�&r""O�J�ԲL���7�����T"O^\P�k�5�y�F�Ƃ���2a"Od�:��%��<5.�S�^z1"Ox��#�Z&.�ت�FڲK�eKQ"O$��(�,>ͼ�;g�G�z@��"Oʕ�%I!!�0.{�Q)%"ODx�5-�1��U��GĖ����1"O��Y�L�?�ΐ�ƊZ���P�"O��6fD�!�*8�E�bun�V"O�[���9A�)j.$��8�"OL���Of��L�en �q����"O<���mx����5	���a"O$�c��C�i��u���U� ���8&"O8$Y �2^r�9�c���Х"O�;t�Q�����	�Nw��:�"O�b��)!�Rp���Ⱥ'��9�U"O>	��#C�s�24ص�˹;�<ġw"O2q���I8I:�b���:Sn���A"Ol��E��7o�p㶨�4jc��"d"O|�r�'��b@���L�DO���Q"O��q3�͋��(��,ե>]�|1�"O��������݋g��<94"Ou:���<v�~\Ȅ��P��-�"OrA� �z-@t2u$Իcb�r�"O�=c�m�����Ƣ�)�9S"O�L�b����=�bB��2k0"Ozs��\x�	0 �//�(H�"Oh��f�G���Z%�;�z"O�,��+{��d�\��B�H�"O�Y@��P�R=���,v��E��"O��Z���K��Rq�j��0iS"O����H�I�0y��cS72Ǽ�sf"O
�q��ٲT��j�c�!�n��"O@�C���� P-��_�R�"ON��b�ҍ����7��		�@qu"O���֡/{���,��cb"Ox��ș/�bّ�R)�ԉ�"O�2�̚+	4�b[��b�(�y�'�2F��x��� @�izA'��y�m��CpRl�k��e��Ạ���yR�A�v=�S-��@ѷ%Ƶ�y2���I�R��C�*Nm����	��yi�{.虅�
�<��� G%ˏ�yBc�H��dB�#4�X{�D���yr B*T��U����z����oT1�y
� ���j�5[�t�1rn� Y�
��Q"O��w*O�N~�X���.n����"O�X�� k�D�3��E_U:Hi2"O��p��M$����ϙ	N�#�"O&j�Đ�)5�À��hJb�"O���+J�Q���A2b�2!P*�"O�!R�- B(I�@�r	Ѥ"O�|��9Kp~�Z���s��� t"Oxa�4��U,�b�/\$�ҴR�"OZ$[���%&��s�2Κ�s�"Od�B�E�nn�s A�5?���e"O��4�/"\�Dc��[?i���{�"ON�� ��(xp퓰Bq��"O:���у 3~��눘Y"U�C"O9xbB"�U8 $��1oh� "O$�*wOY�M�x�"�%f���h�"O�3Q%ֲ&��r ��/, 8#"O@�f��?N�P�+ ��.5�]B�"O���ئ{U�4���Z�؆drd"O2�i��Ơ
e�us3�W?r�ӄ"OV|�`��0q�*�C���:b��"O�)�FV�(Z�`J"�Z�|C0Z"O��ɑ�#W>�qd/�<��"Or��Oԝ5��!�gʴg�iX�"O����|����F	8{
hu"O�%�тA6��;�e?�p+�"O����h�BV���bdQ�A^��"O��rW@�{`v���?"z�j�"Ob@�U�9sQ:���~+T��y�_�s�$h2@J).�h8ɇ���y��d�0'̕�V�*��@	��y�'��lzL�%	�d��Q󧥚�y����v��,Y���
`���"��y��\����q(�<��c ��yR��_	x%q�B�"�JA�bm��y�nV�y,d#�k�8�@-����y��T#2��@--�0$hU��y�L׾n����Ĕ<B5.��C�T��y���2?�ʰ�����#�Xu��GY��y�L�0� ŏ��T��3���y"���my&��u�uR�Ο7�y�E�w
�أ�M՟~X(ŉ�i���y�ہ/>�y�$B:�h�3P�J�y��ޫ4�����.�t�r6�H��y"�M���:b �7�2u�U�;�y��D1aR8�;F�t\�"r�A�y2Ή�a���sc*W�	/|T�!"��y2��a_�����
�\x!!Ԑ�y���J���
��/?�j�D�#�yr�ϥF�~0�բ^�}�L� q�Ɂ�y��ʥ;"P��	W�hX�1����yB �<\\%���$7(����y"�� E䰃�
��7�K�y�N�����H�&�($-P	���ѵ�y���"v<
�	#!y�M9��[?�y���:	���k�\�Y����y�C�1A����B�b�^�QD��y�i��L{��R^�X|
d��.�y�`Z�r��`�IQ�"��hC�7�y"8E��	���C��]q�I΋�yB���Z3~e�,C�u���_�yBJM�{a���'#��B��1L�1��'BP3�e��?����ADϢ&�"|��'#,XVφ�$̼�
T�  ߖ1[��� �y��/�>�d���M=S/��S�"ObiBf��Xs��"-�p
qf"O�M�ƚ�Q�q8��؉QR& ��"O�x#��?�l�'e�7pX��1�"Od�r�J(*�bGm�4$A�1��"Ovx�V�^�:O��QAn�**6��A"O����	HQ�e�D��(Iw�U�s"O���E).8���ρM=���W"Oz��]
r��3��)�&"O��굦�7&n��J���0����"O|��B��
~:���%��!�:�"O�!�7�ǵJ��"���8�t���"O^uр����j�����"��"O|���`7��Z�|��M@"O6m{rg��0�"B!�2)+�s�"O����ƨ|Ʈ��oO�R: ��"Ol��R�ߥr��\�An�){�D��"O����.�np�c.�>�*�A"Oܑ����`���80��y�0\hG"O~!p�֖`�\ղ3�ů(�20�u"O�w��~-��j��#pzDP!"O|q�%�p7 �W*ʹd�å"O��
�L	4O@L:��N�H)��"Oj(Ň3�2�X��B"��y˗"O$<��*ۓs�M� �Z�}+�Tr�"O��D�_�Q	�1T�J:+&L5p"O2���IGJ"T4��
�BEp�"O���[p؂1'
��|�"OPa�2#�)#ᩍ�u���"O�bfA�	24���'ܘ5"Oİ�L� Sh�M���W�H��D"O������i+0�c���m��q�u"O�)*�τ4��t�O�#<�N�[�"OR��dAHB9S�Mڞq��=�"O,��j&Q�8xZ��^�0����"O0�L�<������R�  �S�"O
5�v/�"2f<#�S
6LX��"O`�!��Cń5�Ʃ������5"O*�H�aM�`⛠.��(�\Q ��,D��S��+L26�ޏ,5p��>D�t�o3j_�����&&X���;D����ΝLm�&��?v�*t��L>D��k� �$S�0�A��"mN��!D����Ń�1�\��TJG�p�@�cc>D�X�RM�;tB��"Y�T�4�<D�p�2J7$.��V"��"M�3$<D�t@�e_�<u
 �C��Kl
��щ:D�([$�H��lIƁP������8D�Q�˅�0��8C�A ��AI��5D��Z%NB�ZwlH��ʌI����1D��G��f��m0�M	,|���;D��W� 4J�Dm@u�E�Tة�,D�d�ggR�x���������=�k4D�p��@�O�F��J��G�E��'D��Q�� 
=�V93aÑOޞm��$D����-W���Ѡ�����j�7D��P�Bx�H�K�8.9C�0D�Kt`AAƪ�r�H"7��Q6)D����!����;���S��`� g'D�l�F+\Е�A��g�a1�)0D�,ó#	�(�-Kc�D�j� D�"D�$	�h�O�d�)�Zyh��!D����Ði��P����vX���4j3D����βA)���Uh�-(�U�%2D�� �`��<��B"�� E�Jh�5"O���@�- �.tȢ���9F"Oݑ�F �_�h勀^�{JH�ڑ"O6q:Ц*J�V b��C+T�0��"O,��3��S��q���]�y�"O���@�IVi�P@b����j�"O�azB֋����&K����"O�89�,1*�8*������B�"O�X�#'�i�4⣅��~�ZbC"O���u�]�4�0!
��Q�j��a"O�� E`_�b�H fl��np|�h�"O��F-�
,�2a�c,�l�T��"OE���Z��+FK�J��h��"O��RbI�l&��0]���*T.�%�yBף9T9�C`#c���)��W�y��V!qJ��G#�o��r��5�y	�)$\|"��2]��A���X	�y�<i��iKOt�9���:�y��@�|��!E�>a�!
D�B�y���b��Li$n�/pҘ d
��y*�<�ܙ�@�^�0).�{�	O��y҇F�M�bq �Y8v��*��ǃ�y��Cn��幁�D�m7���B�y�C�L��e��K�=T6�p�����yRN>(LLA��[=j|y+A�O��y��/Q�t"lЯaap%�����yb�ƚ ��umJ)Sq0Ɩ��y���r���թ�9Lۀ,ZF�I��y�AE.K���84NC�<�j�X�GԢ�y���!SP����1�f�Jح�y∓�2����vJ;;��E�h��yb$�\���7'(-k�r��y���0-�q�dCɕ<9bȓ�Ƒ�yΐ-US�����%j( ��,<�y�n�&�dm�K�D��qqK��y�
����
�#�2c)
%ȐjE�yB/S�I������&VA�1%CO��yB��7%I� +���Q~f)��*�y��=ttI"�׽Oj�=��)M��y��ƟG�f�8 	9�x8�(���y�-��-�&�h�) �6���!�jU��y���4�D��f�	<Z��-�j���y��Bܠ�aK�L#L��A@H��yrMY�	A�<3��.>n��5�*�yr�B
��@kw@X�)#��Y�c���y���B[`��t�<Y-2��T*��y;Wi.�@�.�%�]KuϞ��yrJʟ*;Ġ;GeՁ��Jp�*�yHۨ+���(�$B��r�͋�yo��<_,HC�[$섐%Ȑ��yr�-�hQ���P�)M�ـ$���ybf��Z}E˶���>�!�K���yb�G�p�Q�d�rу����yB�
��ySF� �* *�$���y�e�8��D��O�A�6���L���y���7E���:Dî=e8����'�y�X�{8���v W�<� ����yb@^?v���ߟ/�*	 �D���y�$ۤ.�1�A��Ux�����y���
1��1��ۻ_��˂���y�\�yk��*���8SI��0�#��y�c�A=��R"c��JcPa ��0�y���>\ �H�JY��jB'��y2��<\��!�W�
?���ǝzcZC�)� P]4�)z�ڰ`�iΉ"�8�a"Oj�ZPm���අ�(�0k�"O���s�8�8�!o�8h� ��"OJ���" �=�tj��QT�L�s�"O�9�mS�s�X�d!��s�\D8p"OzM��ھt.a ŠŗG)	��"OĤ#�猐�8xP2���Lrl�y�"Oh�����5n&�툶O�>`@Q��"O���7�9�k_�U�ܡ�T"O��"R�R	PI��E!�>���u"O���E<rM˓@вn>�@f"O|�0$�:݄�����"||%�"O�,���A�A��`b4�Ǚ<󢅘�"O�D`�A�Mءqw��4{�n�A�"O �P� !з�S�v22yJ�"O���n[�%��Eq ��%-���"O.�X3d�<X0Xe�&?$|�Q"O�T3t�; ���c�TRp@Y[�"O�E��͟��32��=x�XC"O,�'`Ҡ���ɍ*���"O�ض�ƴ����\��j"OZ���6D�X�I��E3k�>���"Oح���]�4f���ʍ�.}��"Oތ�g��7ͦq�G�I ����5"O(|��DR�AfXP ��SzdE�"O�*��7c��% �d�'l@�x��"Ol$��]�5�x�!�"o)F��"O:q�D�B|�:E��m�I�4"O|y8��#T��ٹ��2U��s�"OD8�#T�F.q �G[,�p���"O�E�t��%8J��R�B�@���U"O����n�'1h݀A녃z)����"OP��&�Ip�dӄ�O	r�z��$"OD�)���ԂA ��-PX0"�"OP�b	W'Jz�a�(�j���9'"O�a1�
����5������yBc�+r���x'�٧4��{Ӡ�%�y��G+�Z��&y�x���'�yR��9S���Wݤ��}��̵�y��_�u�)�"�S��@�#�T��y��T#9��@	� C"AL�,��y䙛y:<|1G�S�$�@�c+���y�F|>�e��Ƴ!^��B�y���)͢h`a>.L�`�a- ��y2��N���0X�uP� ��ybNH9`D��pA/R��Am���y2f^�eD�H��w��ɐŐ�yr�LL]�, ���o�hT�^��y�`�=8����df�R�0�ۏ�y"�U�mǺe�&���v�� 3��]0�yr+�7q*�-�V�˒W�'�ω�yd��.r(=H6�`T���.�y���kCh0h&��V����%-� �yO�Tsl@ 1h���x$�s�S�y��6":��W�-xU\���ֻ�y����zD
y�0)§�$h����yR�1��Z�A�?�XR4�J��y2i@)k
°b$I�xv&|��-�y�혘"� &iنd+j��&�D/�y�C��64f86g �q_H���'��s�͛�Vu�Eőp��=�
�'�6�y�a; GF�@��@5n��5�	�'�b�ХN�!x*��s�kIl$p�0	�'���K�n^���͡��a �L���� b�襥��$)�`��!O�6��t"O�H�vhǆ\�j�7ϔY�!	"O�-� �Om��۷��)6��i�"O���	He\q҇�ϩbpfe�"Ob�3E��%�&43��Pz5�T"O�<�#�ٛSQ\��s+�:"O���ۿj�~�:@-�:��,2'"O��s�*��"(�D����Y5"OZ�B�-��6��t]<(Ǭ@�s"O�qڗ,��/��(���>M�����"OX-��Ǘ0`�<�`���le�Ј�"O<��T	�}��rΜ:tb�V�U�<���٧�b��QJS���[e$�P�<i��2�ؙ����3>���1 G�<᧊�3�m
%o��~�"7�LD�<Q��B�d��PG�~R���UW�<�2(�S���ɗă�1F�9!Ai�<�V��}_�����k�4&�h�<y��(�`�9��ɪf�ER�C`�<�Q�S�m#r�6.��6~�	B1�r�<9���$N����aG�*-����OV�<�qe�8ή{p�s��i�[�<	�*	17C��{���6�@�K�U�<�����#\��[p�(��&�J�<���>Zh@%&�]�A��l�<�3%��3���eX��^)eJ_e�<1v)�8s0}C��bJ�� ��d�<I�e��I�j�a�D�q(�v�<I���t
�]��!�3�|���j�<��:vR���B[8x��ʂi�<�f(�
&^�<�"��<��W�I�!�D�<T��$J�9UȎ`8��Q�0�!�1mĸ�Ԋ�$v��}�Ba�p!�$	1NdA0W�D�W��q�mO
q!�d=k|�,z�@2s8�$*�L��R!򄏂A~�#�8Z�\���� T!�$ύG!4�x@O��Tj�A�c�ܰz�!��V?9I��@⨊*L^�j���a�!������Xa$�~?
:�&ne!��� ��%���M�_1H��,�46�!�$	`Zl��NP�(�`��Л�!�F,I]�0cD�*�4bT�d!�d�"7X-'FT;��0�+�p !��ӑl�Ti
�=��e�u��CJ!�$�r�����fY����3��B!���<���� kΑy�'T,%!�d&A�@,a�"������ &!�d�5k��4��,i�&�!1��3t�!�%k~�1�faU,m^"Dء�Z�U�!�D+4�]b����Cة����']�!�d�4/�$董�Z�%B
-HU�Vc�!�٨����4	��n� uJ ѻl�!�	�Y�4��\�Tw�]�"eۃh�!�$R�er��j6O۝2����\"�!���7	p��#d�lD��+�[�!�P��(q�.��H��ڗĝ.V�!�D'�K��:4{zi	Ɂ�Qs!�-r��1(��^��z�H`c!�[4�8bR�8��I�DHۑ_!�dU ?����
)'�pi)ч�3=m!򄊷zF,�S�� ?gB\@�:6�!��{���r�Cܧ+/%�f o�!�#cx��݀#�ф��!u3!�d��,�l�:'G7b��	�F�ĜoH!�� :��Cƽ-nN����,��s�"Op���֛�0�A��] q�8h�"Ohܘ��L�)"��1�nސ�P��"O��JB�φ"����&8O���"Of�!Tk�{�a'ŕ{1�u��"O汹�F!0�b`�U�Q���"O�����-
��T�,,��"O��n���3�&; �b�"O�lpf�j�&e�d���,��"O� u�\�)����t�Z�[�"O�c��h���Q��U�2�9t"O`�x��5SD�qMJ,��4:�"O�MR`0ec��M^"���"O�eu�^7D�qK��^�*S���w"O��gϮA�������4Mj�"�"O|���Ӳ�Թ9���
F�{�"O���l�>gl�MѤ$�2Ή �"O.�pW�ƄGY�R��&m��k�"Ox�	�b�k#*�C1kSZ1"O�XwCħj$y�$f�&��@�b"O.؛5%ܡ9��d�eB9���"O�X��5L�E�W�M1j�dqab"O���6�]l&Z��l�.1�t)xR"O�$�$I��}y��� *�Jx�9#�"O@M��$�
}N���i� kQ�s"OʝR�%�W�1�ei�*g���q"O��Fֺc�b�[�S3QJҷ"OD@��u������)O���"O�A�� �C{�����lHzL��"OZ}���#t`5` ï/4�@��"O@:u�ռP����n9=uT�r�"O�q���Z-B�#��_>7f̰��"O
}�2cF�#�I�բ�MfJ�˗"Otܰ�O�g���	�G�b[B�3�"O~u9�-F�ei"e�"B�1?�A��"O8��@��'�J��惂&5,���"O<=R���)_*��v!�</��u"O��VK� 1w��Q�W�A�$�C"Of�2Ǘ[.���A2L%�3�"O�EDI+2�p�ن5%l�0"OEI��V����,V�E��"O����X�"Ӭ�"��1`y�"O�,U댨Ac$���ʤ&�8��"O(�(0�X�Rd1#o�1�CE"O��p� R'E0�]j�͈q_��K�"O�)A��9j�����Fy0�C�"OV�C7�Bߊ!;RM�n"�³"O������+�:�Z7�O�3b)k "O�x�A��F��y�êPVh�"Ob ��G�vO�����ԬhP���v"OU�R�$QĤ�cq�G�~1��S1"OȐ��f�6Ɋ��c�@'���r"O��6�b,8�e"ݍ,	��Z�"O��`��
&I�	�����]��"O��#aO�&ƭ����>}H�P"Orԫ�&�;u���-�T��#"O�����[�k)��q,V8NN>��S"O8��i	�2� ���'p�ܺS"Ol9����d�����]O~�� "OD h�ҬzHf�1�*A�Yʥ"OHI�r��$70HJC�*2R��!"O�2��82�,#��O�0�F"O��8�����Ǉt���	A"O�e��T�~�8�'�eט� R"O�  ��ņ;G����� G�T@��"O� WOE�cl�5c�hƹ�*Ij�"O�����M�Y����ö�׬.����ȓA�$JgCJ)X�&Qwb´�(1��HHAP�dE��`s���Tu����E=�,@�m܃F[h�˂C�l��̅�2e��IF���P��m��#B,hyj,��Q���A"�(z�Z�)A��(B�� A�!�։�H�z��o�(Z�X��ȓQ	�q3�Jٰi =��c���ȓeh\,�GM�WʙJU��Z���ȓ\�D��K6)rL�(
׈�ȓ~��u�n�@�N�s����-��*�,��0\�3�h�(�|I�ȓu��%
��,b|�p���+��=�ȓx�\�TΞ�R��q��Re|Z �ȓqS�|�#�U9<gX�¦2��]��8XĈz��
y�p����B?�̄�f*������z�J�u��&R`��ȓ�m�5���E�ݩ�m�z����ȓN�P g�W�va��g߲�>a�ȓH[�(C��о~A&L����5e�����3`���ǟ)i�8)�N/|yԅ��<��`HV�i��aq`�5P�h �'�60OPc�|�=�v˙�l\��ɲk^(��@(�y�<��'D���1"��2�QQ�Yy�<�T/T,���B�43�v5�7Ywx���'� `���L�B�^ly!$�2t"T��'���cӫ^1}�҅���#�l�ߓݘ'�R��%ΏV��1�"��<�\��'�f	)4o��WmD�!�/GhF$�ڴ�hO?7�Q;]+�ux@R|ahL����c�!��1Q���VB�� Ȁ�K��8"�������m�b�Ti� 2BaU�^oB��2 �RL`��t%������[XB�I��t��fL�{dV�"�-k��C�	?#�ȰЈ>�>5X�D�2;!�C�ɢd�f�胪�-{�x4�_�(�lC��
��,8��;cќXۓ_Xn�C�	j���eI*s������%�|c�X��I�4�� w͆ur~H���N850>C�|������H�	i#�.w��C�I�b���*��SWI�v�B�I�j&Uy4�S8��h"r' ŰC�I]@D����U���2�Љ)C�C�ɫ�>����Z�K��@����U�B�9۶L˶m�=9��h[� Q�! ����������bk��T	�1���X�5��p+ԓ�yB�КZ5+�gB ����;�'IIA�- =�QgȞ ��R�'���G���<�7)7`2�1�'1�}A���2pF�!gc�7��x�OV"=A��)[�rl�p{ӊT	xಘ�H_8#�!�^#aB�`V�S�V���pd�7��'шIEzҚ|B��(��3���_�}�!F��yB��!-^n�:���I3�	����IE���$�<	�`ʜ{B�3����ǭwy��IS�O�=sD��V���Ж1�$���i�����,n�TE����Dp�ؒ����'t����58k��kv$�U��Q�A�D@!�$��.9ht�6�C90��81��S&w7!���r�R�	�X<�#%��ZW�x2�		)�=J@JG'Br�`y��ӼH��B䉡Cb(���dB�=vt����1 �"=�#�π �$�F_w�&p�"@
NOB�ʔ"O�(�@��P2�i�TA�$�� T�����*�j��X�f��,�"�)�F���y��C/J�����	�,|�B̤�yr/J�I�n0���8ȴ��K�	�y�H�7�8u��cȈ0x� {���yr�Ǭ!����ED��D!��o���y"g
	L1V�B�h����z�팔�y�j�;1T��3�#@�
�p��瑦�yb9�R%�`҃�`*㍜��yAȝj$4Hǌ��ZHa���B��y�KA3j��WH��q*qС�	$�yr�"P��T��T;����`ݏ�y��ŀ�f��i�E�� #đ�y�AD�m�*8b�M�C���"
-�y���f�|Q	:I��Y�朔�yk��|��dDܿ���Ň�x��'mv� ��H%|�H�]����"�'�B�е]�~ŀ��+R�Nj!gۡ�yr�Ǽj�Bu�!E�6��T�����y�ݸz�f{�R�+A�ՁD/�"�p?a�O�	+'$�v96Dّ��-"O��c�H�=�\���E46���c�"Ol���<��U�'�k����'�����L�#�Ҡu"��@϶7�az����X�z�j�'8[2�,)�.�i
�'�x�g�2Zph*�D�DL��'����A�֙U�¬�v�O?"t����'@±c�ǅ�<W|�F���x� �'��Y+����;2��Y�|_~��M<�
�i�qQ��%_{��@�@8����}J��o�<�Q��K�=X�U��`s�	R*9d� ���\:C��E�ȓ��d�!A��{��壳%	�5�m�ȓ+v����ي[�hE(�T���Ԇȓw��i�r�ͺd#� #�	5Y�ȓ�n|s���?�X��1	X�^=���	L�غrDF0Ab���n�,R���3h�8�P3|��) ��E JՅȓ/|$��f��C�i��=8��ȓ'�pRa� =d�51�m��r�&4��ThBy 1��(|��S�@Ҫ���I�)���Fzx2(]8VU�Lk뙜L�6B�I W� ̰g�('���$@V�k^*">)��I�
���!TbA�9g����<5!��<n�*ps3.��b��)�6'R�O��pG)ǉNŤZ���1��k`"O�0�7D�,B�rM�ec8$0ra������I7Cw��򊇶)��gA�I��C�I�[��Uk1Ό�s2p��p�N`�C���2�+�gĵ0C*�c�N*�@B�I:bY��)��Yl�*QQw�2B䉻j\x��©�,X���M�&��F{��9O~�Q���B��r@@2?�@�W"O�y�@"DC`%a6��-�&�C "O�1;��C�flنL'M�"�3�"O�]�M$Ĝa� ��-/�}"OΔ�U
bsȽxWH�)c�r��"Ov%�C �5 ?��IuĈ9;��!�3"O>tP��
{������)�"O�` g� p7b�S�`��xQ�U"O��B΄�/μCO�.U�nŹ�"O���R�c�^]�rL^8mb�Z#"O�Ix!�O\� WI�_u��ѵ"O� �����މP``];�b��aR�7"O�H2N΋.���Ț.��%@"O�t{BmC̜I�JL_��"O���g��,Ei�����N�1w"O�MC�L͋""���pcX;����"O
�a@lס���)�:!*�'��O.̑��E��F|5�҅a��6"O�j���3B���x���j�v��"O�%�L�=�� �ʜ-�j!R"O�4�۴�t���H6���9�"Oք�ӊǺv�Xq0�P:F�X�k�"OLH,VI`鱦g�#��И�"O�	��X�@D��s�'Q�%����"O�Xk�ڠ|C���rjFX[""Oh�%�C����*�ʔcF�=�!�d�-T��<)�FP�)Pw�,�!�ۨ�v���-�<)`� �ԦI~!�	�W���	4LˀXV��$�Pk!�$ĈI Pe�$`?�H��%��1�!��oN� {A'��%����!���2\��rh�2X�-`�vB!�DZ?&>^;t�.l�%:�!��V&!����6�ʄ(����JC� !�$ ���
� ��sB��6�!�$��&Q�]�1"�k�^該�_]�!�Ĕ�0hQұAˌ.�2��f`��+�!��]^��LxmBx�m"ao:<�!�d��H���הgr84���D�!�$�7<�"I'�O�Cr�5P��V��!�:F|.�i�_���))kޣ%�!�$ 2~L��)�\��d�Lђ7�!�$	ECj]3��#X�8��u,Nc�!�$R,Q"��ř=c�) &l;!�!�D�~��|)�Aѫ �^aI�Ր)�!�$��|l��(�l�乓�IX�!򄆕t��(�`%K��hI��ǒ�SJ!���e��$S����jtDc�O��V5!��.CP��Bb�5W�\	1��!��Hʆ#�zn��[#�O�#!�L�!�ٲP$�-	�m 2�T>�!�ҩk��a�甐B�`��_�;�!��úe�"�:���x������G�pj!���"~����/A�T/(�	��lg!�D�0.�IÜ**��[r�eM!�54U`y��B�h�L�s�k+!�G*uLu����Hx��ȳ4!��Y;4�:wO���Cg޽ b!�$�|��!Z�$B4u��h��d!����ɛ��
bR�ȦC��_az�芆6�DX��%(a&�`p��)v���G�	&&L=�����PyRa���^\
�]Z����`��[�<yb�ٯ	P@�H� �	��hJ���[�<i�+V�C���˃��$%p�rǀV�<Y �عg1긙� 	�&��yQ ��R�<Y6K�*^"��-��en���"[e�<a4 �*G�0RHQ�'4�0���Da�<��EX�`�X��랱'��i�Bb�<�tLl��1G�� j�t�&�LX�<��k�w��C�"ӾR>��O�m�<�����5n6a���AXw�<)���]�f=;��k��uH��E{�<���B��D;��̇�:�:p!Jz�<� 5$I< �̓37�%ڗfZ�<��Ϟ�Lw���8�<��G�U�<� ����7] {Q#kZ���"O�i�Ԉ��t`����M*W"$��"O�t`�A�O�ezs��AJ�W"O�a`)
1JL�(�d��tn�A��"O}��Y/g2��������(�"O�����F��do�(�9a�"O����"��Eh������f�i"O�aX� ؙ^� 
2�#3���q�"Oȳ�� �����NO�y<(�#E"O�P�����i�.Y��� �"O��V���!���(��%D��Ç=8��t�D�(Jm�A�"D�X��Y�;��򵪟�i�=���>D��r���1k��x�J�)b�����3D���r�ԕL�����X 4�\�*3D���s��%Q~��dKB{�>�pr�3D��˂�/y��i�u׃�Vܻ��/D�LR(X�����*՗8/���k+D�Ly�JR	ͥi�,���NG!�D�*Uor�X��� r���A�C�_?!�D�2yԸ�з(��A��!`AŦ49!�D� W�L{�Obc�����S&o"�|�/�N������)����X�֤�tɘ�0@�m�ȓ[��ЙF��!]�dy��l{�f0�?�@���H���,ҧ�����&�����9�u�ȓ&�,	 "�<fW���T'sD	s �'x�{V�<�>��o�>K�����W�b��H��Pr�<�w�N�H8j@+r* X�Y���}V�x��c�5!�N� ���Z��1 m2�蜲�lB� z�X�(4\O�4�p���.2uD��T�D���O7rj���DR#$�*N>��d�! �:vm�Έ�� �`	�p��0@�OȎ8"$Bf�dH�=,
ƥ�2%��+�)��q8�\��Y	�hD3��I�8솜�cO��q���#x�̙�(�3��	�8�z ��C�v	ןR@�dأ+�u����`�Or�e�s�<�0g��^r�,���)c��хnη_
�e'�ji��*��J\��z2*�Wf@k�䂸2���U��d@�F�3 B4�{����0��	�f�xh�ƙ7d��ʤB����/U�*b��΅S(����܎�0=YWG(^���F�z�$���רu�>(a���'jؾ9c�!��	�MѺi�,A���:�NV$��^=��I�|�0�ag�F<�<���Ć�>��AI�I��=�M3�9.��"B��p��\�u�øV��O���b�)�S�]���!E�ϹM�f�����"9 HV�pq^y��/Xo�B�����$S� �W�ܻ?�ѱ2���b�����F8�$�G�b ���&L;����"{��m`�@9c�x�SYl8���N�'8T�h�!j^(# ��TI�c�}��I<QB(\�U�����q�$�#:?�+'J�>��UG�1j�ay���	9~b����`<�,�A!�x��`�65�I�zD�E+��ܴ�8�u�pExD!3hɊ<�8�R�d�+&�2O�e���z�S�5b"H� o
f� D���еy��@c����x�*�<�3�>Qu.�!�p���툵V���ʎ�U��k�`Cq���g�L���1%�`U�K��P�	RP]&A��ax���&ye����¢$�~�i�#���|�ao��le$ R��':�D��<�G�F�	].0ÍǉV����M�J�'�h��%�0�t�@����t+��#u��1fk�%'�B� wh��yR"օ8n�Q��ֵs�]�v,B��y�F4?�dAs@�l�.T�r���vl�}�2(V(�t o�>TVB�	�r@�t 	P�t6�hK��vgD����j�4 T�8��@�|Fy2oBLSbհU�V�0<F�bA���>i2���d�0��BK��
�S��M�����A�Ȋ	+��@!���g*����Z�^AZu�'J�����C27'ў�Xc� R�Li�$)S�g����\?Y�ǈ8N��x����
@�c�� D����fJ��L���G	B�����O���W�
��ԍ	d�E9j;�����i
h�X��b��w!D�4cC�@�C�	�kC�]I���*O69�V ߮[���F�ڔu_���DR�o
���U��|FyrG?:c`�H�O���bT��ڰ>��(��-�شh�$i���p��� b H��!�y�m�D;���)� �ѣ��H� ���Xv'B�M8�x!�&���F�	#'��� �gC,N>��O�%�v�V7m4i
P">s����	�'��ѳ���r+����k��=��ٽy�P�I���2E,��Y����}��?`d�B�`��͐r�Ȥrg"O��;g�T?6mH�mR7P�,̑a�ar�da���a�<A{�m�-��	
<�`���8��Ȱ+�{1���dï_<��w�5/�x�׸�� `���]6 ��"�ʥ:Fx��	�W[��H�ʙ�;�
�!lI�w�D�?���K����a�T�.z�1�#�XR��_�71BT�c��{��RfY��!�d�!J���K&%���+v�ɤ3��b�Aԩ;]�X*B�^<f �\:��SY?镏 	}�l���ğ*� ślt�<�2���XNP�p��a�蔛E.��(�
,��%��~5`�n�:_�@��� �j}^8��'��*E��N�Q�HT��I?_��a@��)J/2`�"��VXh�Tg��1�ƈ,K������~D�7F�PT2��`1N�i�����a2F�Qw�[>vI�P;����$=��2vc�Z�i˜s��L0P�ߵDj�����3x�!�D��<���8D��+����$РҟtGV����]=w��@1��\�*T��"���G��=�<q���Iȣ<���\#���W��Ȅa�\ԋ�.�6e�����K�7Q��ܐ���?��];v

�O�Eken��Z�R�G}F�3zC8$���B��{F�Tc�0�wC#b��;�O�)ȇF�5���P�r����c�M`�������;dڸ+��U�U�uH�JV�9���Cs|�r덦3<�R2Ϝ8Iw��	�,��tc�/"�ҵ�G�D|b<�«�$6"�R"\8Hv���0�a �/Z�X{Z�@�ꆎ�T��$���T���^b(p�(=aR2P�⍎ ��l��bK�t�
�kօBf!��p��"��1�H�}��C�(28���'wƝ��������QbV�T�yp�{"KI+�,���E�@��ŘdO�������9�@����\��i���az]�:��U���_�LO�H��$R�����<�R1``�@��iFx��ć�`�F)�C�$�<öaE�Mp�fԓS2fp� LR0lXD�P$Fg�Za�#G$V���b��0�t�ٌ�,�Ac�R���B��,�O�!pɾTՎT�F��1p�Ј%d\$���;���n ��`�ʌ\K�8��H�Rޚ|��B��	y��E�%��P����EZ��<iHm���'��ݙ�a�U���3��<(j=X���/>�q���ј!��pS�B�V<���Y\|�Q�ʴ"z!h�e-8�m�'���Ĝ&z�$x�U��|����d�j���=9'	�5UZ����Շ)��8�Ԕq��M!c%ջI�R-��)�%�.l�T�B��B����܌ R6�\��G��Vu�Daȍq-�P*W�H�4t��D�*o��p'bζF�l���-�%iF��faIt&�|K��N�*H�䐨i�� '���r"�e�J6������eE^q�m'�O�����:MX �"��,��@�2��	��ą�,�,���ꏔ/��ٻ ̎;IT<��ɓ+��t���\>�(��-�<��q�g� P@��'b���_�x����M��D�3y��8�����sB��ܦ��poՂD^���SzF��������HP��N:,�7�k?�r�1C����H:�3�ILT�%ą���<(�%
4f��g"t(��[yB��!���a�Asd��v�Ru_2urRό)�Y���i�<�h���g�'c�,:�&��GQ:� ��g]52��Q5��mw
���郌y�aK���8nl�!��L��\&�}Q�N]�z��Q��/2����b\W��x��<�z�ү)c��¥	���a�C!;�I8np.l#ԊZ�[Z�$C�e��!"���B8q���Cab�
b�*��P�p=��BX1� �P$�L�z�ڭ�TH-� �2��n��]���>yD(٦����=�䑰��̖*��Z#ُi��a���O��Ƀ�ʤK6nQ�6�BD�nyT���}����O��[[8aʁk�6V��ǋ	 �yr)��{}R11���Ms�8�GG��u���'�ԐDDP���I�|y�a��XP�'�v�AA	�r�6	��k2hNn�jAO���P7�R�H�L�6*�l ����>�E2OV��G�i�4���E�gZt�R�� �_�� �P/zP��ə=Vj|��(=H�G�"Z�,���Eǔ>��ࠩO��ݴ;Z~\��40v�@t/�B�tu8��
�1s�=��c�<<&t��V)��xIZ���ɉ\l�I�qA_P����
)L�z�͖�6�:���A4W�h����T�u�`}m�w,$��[�[&��e�Z/)`�A"g'£n��$�,��49�@�Ht�p˦�ڰCƱO�e�V��y�fԫ	�_2��͛�o�5���o
v����M�w�@�i�bM4FH�& �m���+�jEs �#aEj`�>��J8���Y�[(�0���@�	��\��� B���)�8h��AjL��?`��,�"�� `W�?Q�].|F���C�
w���u�Ƌ1"���W$,�OH} 3�ɓ�l�A���e�!�S�Յ3�,!@�'Dfi�k>�Fa8C^��9r��_����w]�L�Ѡ̇����҅��p>q�/�Vc YyÁ�,���yE�Y�meB	��Кe��Bo۝Q���F�] ��0Ǝ�)��)�A�-nbLّeP[yr��g�dPFC8C�Tp��.W��HO�虇g��}],��ݢd!�E#w��	V6�Lu�6hYb�{ۗ _'Z�<�!ۡgu���2lM8)ax�H��8��M�b��)	�����?��l%%$���b@̏i,va�G(_&=��aJr��(���BVx��A�s�Z)�� ���+$מ�ٵa˛s����^�a��
�. �=C��).�����\%-��5��@Y3%�޼�R�{��cƆPK�j�<� Bqceb�"v��蚖�ԥ���ۀ�'����L�P+&Xؤ�',͜P�˛5��0J'��JŦL�",�&6���8��Ȣw�<�?�g_5HB$y�$QT��E��]�'v���MB�1��Ղ~b-��{��Q"���*Nm�Q�ƃUu�0�5��$A����D��ko����ŭ'b��1d�z0��>XN�2rA��N������mb���C��$f�ތ0 &Y�H掉`ץ�>*캥k$D���G��5F�;���m3d](F!«�nAI�Õ�%� ��&��g4�rD�mBэ����d�	~]IT�����p�DQ2C�~�� !�U�Xf6���/X�� ��\�4@P�NR���Q���Q.V�F�UσD�'0z���cR�~@��JT ���ɏ���6o�����J�V�ݨedM�0@L��'��M��m�4j	 2��y��%Z�x~H��s<�[뇶l�")��xr�(�'۰�k (ȥ3L�����J���-�������x�KS��lP"�]�woLp��"O��ڱD���0�1�ѐ}ObRQ�O�D�a�N�[��d�!����1�)O�!j��O�pX5���]ƨUOBA���O
 `3bK|�>,C�aZ�I�� !� 7 �J���C3����­8Y��j�@'_����C�z��}��C;x�$ĺå\5w�N1#�ʻ\��=�sk�:��Yc�'J�y�r��Y���(U�m]&E!��ɱ.U��b+@��0��,�LxN,�P�޷$=�ȓo��tk�k٢#:x`���ʰ!K����^���#�}�S�OuByH�LRL���
g��-��3	�'���j�^Hƞ��O�z⎨�'Y��P"G�]i�����&q�p�'��yՀ�3H󪐫�*ˍp P��'�4a�u�^�x���ҔZ'�}��'VX���:.䈣�U��IY�'S�y���/1�<�/�/J ��K�'�V�3g ��v�RÍÀL�D��'��C�cӢ0�S�ĠD�I��'��407dR�����Ӥ0SJ�J�'��H�$rH�y�雫*��(��'�c6�܀gf�	���v�P�3�'S�1Tʇ0`W2`�.�;>t�UK�'�6Q��
Ƙg�l�vC�&����'�.A� �B�z-9�L_�)���'LDl�`E%-�~\xFeޔ�����'}��2��͢@35�D���jIQ�ȓN j�񎖾���0�뙭�<��ȓ
�n1`��{>x��#+U��	�����o�4j�9V� vx��#��q��)08��5��7};T�ȓ?; ���'T9<�\��`j�R�L��	¨(�N�y��	�E� �	պ0�ȓr�*��RE�'zI�q�P�S�u�ȓ��J��K�J��p�'R��H�ȓ��C�Y-A��X!4g�"d��l��!����
8:=A`��������L��t0��Z���-��@hw R�<i��?%&��8�Y�p�:��F�Uw�<i��\-f�0��>G��S���j�<9���\󆐢r'�KN`%jd�IL�<��靈8h�-XDE��k��Lʑ��M�<�(Np��0!-�U�A�S�<Af�s�� 4��W;�B��D�<�7,O8V��ؑo�Y�(���J�<�E��I��)�C�٥:� e���<#H��P��K�!����w��u�<���Q$L��E�֝V�q��E[�<���o�kQ��Z���2G�[�<��]-�6�I��;�T�Sa�XS�<)�fՆ�&�"�+ ��\Âh�J�<���
8�X��b %�>�A"&�O�<�5E]�'�$�� �.��|9t#�G�<� r� H�vJ]#4�I5t�ԹK�"O����W>$�^���hY.i�кP"O�\V%ɇc��Y�Hʧ!_Ԁ{"O�xW&�DZ~�����/�ҐC5"ORѸ$璃;Mp݃hĎ5����"OL�����O'P0��.�3w���"O� �#&�%Q	�99���]�����"O,����J����a��6�j��"O:]�b
M"8V\B�%E.e��	$"O���s������~�(W"O�-�#i��<��Q '�U>\���"OZ���k G�Y��YG2ЬI�"O�j��P�%��cWCؖ�P��"OP8�bᔶNmZ6�H�<s�"O�В��N���� O��'8P�!"O�A�g��Tr 1��J�l�[7"On	�NW� E�)�� H�rZh"O��ؒ�vx�SAN�D}���"O��#i�.Ej����ΧLSJ��&"OָK�3TоQ+ǯИEQ$Y�$"O(�3c��lBt��|D���A"OD5
¬�#4��L�����!:���@"O�uj����_��Mc�E֞:=�+�"OR��/�,6�D�DW2c�|��"OzXqV&S(I]�-���T�.pr�"OZ�����	+���aJ6�q&"O��R�Q:F��K��UP����"OD��%��)-b�*�	=�R��0"O��d�O����:�/� �2�"O�ģ�MH�rqh��F�+n�*R`!�$�J�t���[�g��i�$΅%h!�����������"v�^X!�ė�K��@��ҹ`�-�.A�!��=E�d���,)����p�^�!�d�*�r���%R����w�U�!�D�4��Ի���&%�4�1�FҊ �!���)	D�7
�0V��7Ǎ��C�I�$�Qh� 4STt!�FB��x[�B�	~v~ �r��>E�*��b
�T%zB�	�|��	��;}\=�2*�8S�@B�I-|/��rq!ڳ�,��&Ƣ	_XB�	E�)I�֬@0>��qd�!f*B�	:c#P!@��W������P�!�:B�ɚ(����JXl����;dԪB��EC�f*�'at���v(��8��B䉔u���xe�O��8@d���]�B䉠D���1���!�*�R�a�6}��B�I�{(b���.�$S�#׬��nB�p/�0�ю��&�,���h��S'FB�I�$^�-;gՑ,�Z�g�V8HB�	�Fb�QD`��� ��$F��}��C�I�S��8���z::% ��S%��I�pB 5�N'?� ���[ @M;�&� ��YfK4�Oh�Z�c�7����b �_@X��C��c��8X���.���>].�#3N]�\Ί����E'�Q����E�91�������v���E]/Y݄� ���?��C���\�!��S�(���K@l�Kݎ�I�#�4���(Z;�����XV�O|<� &�;Jje27�@�;��Q�'�R�$�� C���p�����5s��B�8dˌdP���K����I�c��S-ڛ�f�y`%G4����� Լ �fZw� y��
߸F�Zm�%�@	�(Gn~���c�������K�MAO'd$E{$ �{�n+�N,@�R4���D��H݀SC�A����P<�dq7 ��yK�?V�Y�%ǻlAh�䘗�?�#%]4Yij�c� �`G�e�F.�'�� 
�x� �H�Т�ٷ�!�F"O�\���N$�H��Q�Vd�C*��k��Lr�ԑz��5�G-<��3ʓ>v�diԭE;M�@+cM��Z.✆�	��P�qeg+�ʬq�.�8`\+Ah��s�!�1��P��C&�O"�i�	�*�Nْ7�'4��7�	y.�)5iЩ�T�ʇ��$2��O��dۧ��$N��F��)D-8�'I��zůFi6��
��O�7�Ř�D(U�z���#�(��@1�Oڍ{J��}��1ݐԻ�)� t("$�#o��B�I�p��5���'��財��1(�h;�ޣ)�\�9��_
(T-B��?�=Al�?�L��OC�l$"��ek8����K�/�<#Oζ5��7g��2���B�jy�@� P8{qa~�	� ���b��5R�	@U�\��?IEJ	�1�B�b��Ϭ!��x�'@��Ӷ)��P��ω?9��\����#R\!��L,��9Rؠ_(A�G��4h���ł��C�l�ubP7}Yh��+�'�~�iU!~���C*�u&�ڰ �>�y�&Қy?����)׸~h����#�#o.���[z�`��w��(6�y	�fZ�'R@�i����;�����/�����_���;�(@�C�VQ��j��CB%�d(�3j�3�-T�F�8�S���O����d��H���3�O�	0�a��H�.��'2�q8��	 *�4}�)�TA���p�����^��#U��VK��Y֎ߍa�\C�&+n� H���N��HWnߨr�A�RF� Q�L�@��q���:gN0��9|�Ƒ��:������R����Lƽ~��#=�Ul�t�����	G�8�� TBl�9L�9G�Z��B*��D.�t��a̞��Ʉ�,��0D}�KZ��D�� �O��R����P�C�n�O���x�&�h��� '����e�V��*8��\%�`�sOݮCy��G�����=� 4�/��N��в~G��ɣP�ȽC��Ġ6��P�:�> rUo]8�P�a�F���Z��Ů��p7���;O���dS��� ���!؂��t@5��%Ξc��2��(6�2G�0Q��A�H�.e/�x����o��������(�'����YG��I�!�AG��H�{��� Vr ����$� Ҵ`����ƒIp�	񫋈��aA��f҉������ �(ؕSf���F\
(+�=Q1*�j�$���J ��lJ�N�0�&\����l4�(�!�j�J�a�U�]D�ɵSԨ���p �9�!7E��Y��V�w���BѾqȠ#����b�cg�'���R�HE�d��i�Y��kX+'�.i�ɤ+�����j���:"�� O�H�"Iؙ]����+&���,E�%�Fy0��O�\dl�rדP�<�c�֚\��e�"��S�x�1�MP�6���
��̬�ՌƘ�aC��,�$]a1,[�V�v��-P�5���r*RUy҂�7/�){��=���A�����'������;�ET�W
��NN��|| ��ڕ�4*�cW�$���!����䭳�#e5h�2b��5$@ٰ�:��OfA�&��x&����DN%0��C�V�k����M.HC��	��ʹ5ha��gJ-}-�����"?��3Gוmu��b��/�d�e��*r!���K)5[���I�5)쐃Z8(���ӋnR��E�0$��d"X�8���fE�Z��0b�:(�<1���`L�Ӆ�L�4-�HwS����0 F�	%@��n+\O��Ec���j�����K"|�ۗ��z8y�T��.8�J8�ܴz�Z ��"�'O����'P"�Z��O�#$�T��IZ�(�'x���u�7H~Q�$�:b���R�{�0WvL�����,Dw��9+�GS�=-O$�Y���$#�iӷ����|݀�/�EFtJbNZ�{�bmcaK��>�1��L�t�jLy�g���.�i`�G�x�ΠwM s��Q	��b��gM�z�'���qg���&�:���+؀ ��]� ��#np$�0BNS�:��~��.lΕ�
��U��j۽��̪6G�x��X��w�� 5|8����mL�KPYR(˚a�vA�A��q�z��.^Y|$y���6b0iD	T%v�8��k��E���z}⩍��MÑh[�^�s�镦q�"��ƒ��y�u/�>�d�'��ջF��4~Z�u�4�=+�⇊ݥD��9�M����c�,|�󄚑Q ����!�95$��w��6Yɺ5q�B=ܤ+��	��@��l[֨O�,�􊜘X�ܝ�0˘�w��n� K�ҽ�E.��]g�N�D���j][}��z�(
7�`Ӽ<���ۮ���t�5C���;�m
�]Ͷ���+�A�d���HD���J�n��	���7L�b�ˠT�|��i'�i��i���S�Vo�x�K�Cűj�頰��x9�IbW�1�)�|i����IM�bNP�Wc�#x������> �t��D�0�҇[�XF��۴d�F���X%3M�\����=q, (I�+���I&P���A%�8JϠ�� ���:W|c� {�e[�V��D�3�>���B1"P�p�%�'r��7��c���6b
�"LEh�'��~�a��̓h(����UUy�E}��4��=�`@E���I��slT�l�N��P��+�w�����`��(	A��vfbď�uk�qBC��, �9�׌<wO�j��Xg�� S��Q�b�TAr���2��%A�/U0Q��`�O|xc,�R�N=k�@�>�'`��`����:��Q����r���ƈE�)�'xU��D*u��[���.n���*�b����� �9� �L��U1�N���1a��"+~�����e���(O)(�	�y�,�cD��!޽{F�I�;���4�N;n�Yb������h ɀ �ѫ�
К���eMӪO�N|	�A��x����O,^�<��Dk1axb�q'l5P �B>d�|� �C��?7���6�;v(֏W4��y��ǃt,z �)�e�x��Js�l ��]�5��bR�R-f� !Yƭ�>2��Q��g\6��ϙ�&����&.D?0���[�%!���*a��*�Y�D$I-a�.�1s�<��+�|=���ŒŦ(�Qf�Ox� �1���['�C1g�,G�pi@���:m�b�49'�P�Hѭ
Ǫ]AI��+dY�S���x|$[�M"dh�đ�"�Lj��=���� h##��;~:���R�/}�E��H�$Sz8ȱ��-��S�̳�JT�'/�P�e��B�@!�Sm���h��Z>P��Ռ�$1��o`"��8a�I����2�IŪ#��;��I8��#E�%�0C�	�G8E8&b���3�$�6�!���f)�D:�-�8cJ�8)0� ���5���<a�G��7af�D�Ѽ#���t �K����"���$�g�Ę<}PUd]�.�4)�� ~�^��p���PH���nR3X/Ģ?�`�GG��t�ҌG4�k�F�M�'��4�F!x�h� �ɜ:0�v`�3��<Nb�a�VΒ�PQ��1Ci] 6N��Df�V��D(&(��Q�$0���]�9�B��<��
P1bl1��<�!RT U7��8U��df�1H��)
�b�F�V�zf�	��y�@�
��Y�NP�<:�;�E<��� �q�a����S[����Ď�Vy�br����1B��T @'��xR,R"iX�u�t��'Z�PUI3�݄(J -��eܧH��a���7$�]���'��0a�lUXl̰;��2
��ı���Ё�ʊ�T &��AȐf�\Pj3�7i�ICA �](<��'	�Gr��J��E� ��%[F�'��(���N^��c?�˃��+�p4HE�#Cپ�8g#D�x�F*<@oH7���m�՚P���rC R� Ǟc��}��0%�x��ԻN��R�p�<) �ݒ>�ȧ�65Kx�R@ Y�<	�A(@�	�.�R\��S�<�ƌ��=�n(Jᬒ�P*��0o@O�<��O6F���*�AW����Q�<Q��2��m�dC$t�Q��Ot�<7��7�N]S�iȵ?��L�.�p�<���~�+c�O�Nbd���_#!���uW���¯��i��a:��S�U�!�Ď4,b����Y�g�H[�6h�!���]�8`��N�N���0b��!�䊮;��p�+�s������\�!��5�0iH��c'"Db��ެg�!�D��T�A�
-y:�� �2i!�d�:�P}��B�3irh0��L'T=!�D�0h��C�$6 V�QK�cs�!�O)�n������U�z�W�]�r!���9�!:/Ө$zmB���i!��Y�M	��H��4Wc�?0�!�E!c� ����.0�@��Pc֒U�!�dB��"�G��$|�xE��6�!�J$KHa1�V'L�Ȣ八S!�_s������~�&�r4囟k!���RB A�P��m�ju�7BH�8V!�ɠydʁ	�OY/����cȅ�!�L�wQ��2Tͼqݒ�X"�7q!����-9ڐip�
a�j�1�ݮ}!�d\H�H�H��1(���3#C'#!���ƔJ֤�hHA��i	!�O����˓iP7Ѷ8{�RQ�!��O4��E΄�E*�8
��X�M�!�X/ur�����VJ�+��azr�����en�	W�d������L8H�bQ*�Q�D����~(��>Q����'1�xҡI,U>���F�(n��C�>���ͶQ���;��i�~���@5x1,\@t�W�/n��cT���`!��_$P���>%?���"رr�� *�n,
4+�
f�Ԍ�I�w����φ"@���S�O��)�Uf>]��D��s:�5r�#ۂXd���U�O<��S�S՟��O0
8�=0�
s#wdZ�� *�$٣ +06�dF!�0|R���K׎1�6EɺQG�pHW�Y�U��i�d�X�nR��ItԞa�g�)�� ��tb��v�p�0��:8�<i!�xr�-uqz}�6b"���ǃ��YZd�S��D0(�BU�-Odm��o���HM�"}����8(� �J&�D���]hs���5V$\�Ɯ@f�>E�T�g���/��`��907�@�V���x�(���D�v���H�O�t#/ʻ����Ʃ�
iyE;e��OA3��DR>�l${)�}*F��;S!~���@ۿn)��g?���qק��v�1vDX��� #���0|����T��P�&Y�7qO^,F��E������B�M0�y���M[�!�B�>��~*�*��s}Zw��4��[q�؃��s��ϙ�KqO�����65p`��6A�$�=3
��=�r�ޙ�@�D�DNQ��&Q�2�M��(u��ē9�6�A�V�5y�>�	)<&�������̹3Ap5��^���G���S�O���:�--���"K/¬j�4^�A��C���S�i0�S�Mdq�"��*P<�ɠ"F+rt, �T&Q�.��
��>�s�O�n�8W��?#�a�s�{�p�)�Ɇ	sx��O:�{�Y�O��t˙<���+p(P	lxбc`�U����OHd˓�}����?&P� �@@ v=X�$X$h`.�Q��'��	�O EcI��H�;��8�#��f������5R\9`!,D�hˆD��%��Т޽z&8Mqנ>D���޸K5�D��ʚ�:���Š7D��!ʖ*(�n9�v�[��I  ;D��1cKJ�n�f��6uJ�,K�9D���'ɥ|+��Cҥ-\g^���7D�ȓeC�*-�����l� k::�k��4D���pL�:~��@3���D*��k2D��Z�Q����Z��`K��/D�lC�댦p�\9qaš[���S�-D���%Ά�6e�(D*M$t,��)D�dq M�i��yY���x[V(6�&D�L�b�̟a��R��ƻg����#D��6��6v��U�P'�y�B&D�\�d�����3 �/}ڱRt�"D���H��d�ZHqF5*"�i���>D�X� B�5&��X�Q�MפQ Q*D�<�c�лx8#�ɅA挍ѥJ*D� x�/H�AP���d�\te�d�+D�@�ō�D�ep��G�� ���+D����C�����}��X�#�*D����e\�X�*��R�PT���@#'D�lzQ.�=*J��XPd֔b&�qA�/$D�`Z�́(�.,�rj�>|���Y��>D��4�=�X8�fRcG*�Be�;D�d��Z/��l/���0'�9D�H�܆�.��w,W(Q�m:�:D���eړx0��V�$]�8RB+D��@�B�5�V/�3�&�c�	)D��+@,�,�0�Q%�>C.�U���(D�:C�ʉ#���{�d�Q�t��@%D�$���I�� RjW�k�(hc�) D����)DQ?~�MU�Kg$$
��(D��@@��%�` �'��B<���+%D����,���aC�&P�u���"D�8����?�څ�a��?�ȡ@�;D�j�d�!ָ�r,A�j�N�He�4D��×�T�]BpA7 �Q6�A�.D�|��@�/��I��J�~�� -?D��22��X�Rr&$�;�d1@��=D�@�C��S/ �R��S0�BY���-D�lj��E2*�Bt&r�$�3`,D��2 �K��h�֪H�cB���)D��rd̎�Y;��U�5���3�"D�l(AU%N�1���BS����E.D���`"�5%�L�p��H~t����(D�9�M6HH�KY�R@�A�&D�� P(j�K� �<X�#���q�e��"OH��g�6���Fh?l����"Oh�ɳb�_�Ca��5-��X�1"O4�&�Y�K�Z��iG7ײ�p"Ob��D��0@=I�
L�� Bv"O����ڰ]Ml(�&���d�\Q�"O"\�*�,*
b̉�Z
��0d"O������r��\��`�	M��$
1"O6i(� ۽]W�4���&|�x=2%"O�����j�Kf���'�Lc"O�L�Fd��Hr*�"��!(�\���"O��"A"���
�J��I*[Z�K�"Ol�a�F�1��1ul�A�"O�5H7�P�|�r�{S�.08��"OVQH�^�[�>���_�LA�"O����\	d�F��B&F��Ɖ@"O�Y����8g&p P��ģf�I�F"OB��$I��4N.$ۆ�O�PAZ[�"Oظը�;&`Q���Lm��"O���aHP�N��\����0=�"O�t��)�����W�W�_�pAc1"O�q�`�:Y�f�lJ�2\9�"Oz�ӲJ]�x�F�a�k��F��	`"O*!�#�/���TJg�m�7"O��Kf� ������7-	1!�$�V� ڳ���8�ɋ�E !��ej΅����2����g*f!�B;̌0H�+�
�"�A0�c!�d��s`�����$`���V!򤆉~��YJ4CNoY���U�ʮIB!��A�ʵAS�3K
�{���~+!����jCb �c�؉�&ˇ�M���'{�6��"aӬ77�Т�����y2�@#BZfDK�n �a��jEOQ��y�(ܼ1��xb���J|v���>�y����li�7I�0n�ӯ��yB,G>g҉��!�*	�J0p��і�y��н'ôdC'� ��s��^1�yBjK#@�Q��Q q�R=y�]�y���,u������f`���L\
�y���){� �K6J��L��-�Ǥ�"�y����O� ���S�:�ϣ�y�̕8?��1�pLJ3Z�3��>�yB�L�+�\�Y=y����͓�yrlL�'z����ۢt�`ö͟4�y2�ݻWdE:�%W�n�h6l��yeϒMk�,[P�ƶLj��j�����y���'<ك'�ןKs,c �W�y"#�!28�1�
�0 ��q��#�yR䁋Gd@����<lX��VhF��y2G�iS>Y"  *;�θ(sA�y��Y�r(�Ɗ�7HDp|�I� �y��� })D��W̭G��4bL�2�y�jԋ.tT8��/?������*�y��	<W4L�ֆ�GjT1���3�y�����)r_%dq��EE��VB��^E���"�M���;�j�� k�C�!nq�I@� �F���P��6��B��/=6<�seh��n�zv�� M+�B�U�������Y_r[��F�"8�C�	�n�dЊ� ѭf@���7�7Ja>B��'w���Նӕ*::[5
ѼV�pB�	>X�=�'�16�h�eh΅|$jB�IU�
����#<����ʢ@TZB�)� 4�xf�?sx�؀Ɍ�NT�,K#"O,�i���x4<ls#��6��V"O�t�Dn) �t�[�b:vy���'"OvUx���-�,@F��<df��3�"O�F5^R2��f�X�JY��9'"O��PkS�H�Ą@�-·OL�C"O،C�ID	�&�cG�T�U�d:s"O�e�0oڟc���H�g�32�"O8H�ס^��k�$�=,���"O���� (��I���v���"O�L�ÉΕg�5x�ӭ+j��"ON4qe�%%�e��N�4�Fœ�"OT�e4��Y���(?�k�"O���R(ӹe�� s��b�(�"O�5�@H0��$�+r5 �q�"OTЁq˟�!\�i��k�2"lS�"O~�aC+D����j
59�b��"O$��mS)L�`�p��Gr���C&"OХ�GMGX<A��L��n�z�"O��[���J$���b�p��P��"OĨ�KJ"Mh)��C�>��5"O�BÂ�H9:1�ώ����"O2`藇ݭv�J�a�k3J)��y	�'	| Д�B�:�c���]��'�Z-���h���;P�K�`d�q�'��,+�<�4�H�ʓ+V����'{����Ą'$��	g��Gy�1z�'��4q!B<<� @j�`��Ca�P�
�'�P���?�$T�R�6K��`	�'aXx	V�ō^��a납0�؃	�'3�1!��8ٲ-��'7R(�	�'``��Ѯ�O3�tA6�GGE4�r�'�6ph3j׻��q5
֥;�N�'��L`�N_@� `���1B�'K�]��I�	L�Re���41��,��'�| zьŻ5
���V�[|��3
�':����mT q��*� ��?vђ	�'dj�@w�,CaZ��D;O'�e��'��TI`��	�(�P�<o��'�X����!�=¶�%7�Ek	�'��x��_11(�����+;h���'(�37�����e��J�; ���'t��X�lғll�Y8iI<�>0��'#�|b�])a��T��̓�z��'rو��6G�,��S���8���'�A���+L�\� R�4;�'� ��ξ
Cd�
#�N�AmDz�'��dr��9=ú��B��>=���j�'�H�sS��x �!� bl����'��8��̝-gԂ�&��+Vz�ɺ�'� X��� ����a?N=���'�ĭYpiF>xRz�j��[q�r���'��-aY.`AA�=T ��"�'ې���[�dP@�N X���'�h�bPǓ�UPf9�wg�* ��
�'�]�0�\�P�@t(�b09�'ՠ�y7#C�<��p�#cN�6<h(�'���p��AS
$�o�#]84���'��!�&�
o����� Y!4��'i\�H���J��y��	�x�'�p����	�`ur5�32ȶ���'g<Y�����( yK�2�FH�'�H��l�s����p�U�0��iR�'
6آE)�\5+������I��� y�%-П�V�3�ȖO��"O 	B�L	"�����#4�P$��"OBH�eaU�%a�-�殆56KR�Js"O�ThT�o7��8�{�B��"OX|�`��4��!t���O�.��B"OD�����;X�֑�E�֭\�05�"O>UB�$ZV͠'`
9��!�"O� KAg����� �i�.!��"O�y�b�/�`y��X@r���"O���@ڡ  �����(q�ڱ"O"Q+1ˎ#S$AStICU\�Ѫ�"OD�(�ˁ���0Ҧ�)?���v"O�-h�j�9f�4�SDہ*ؑ�"O�
���6"���L?}	$"O���tIZ�^�z�S������	�"OJ��礄:{m�82�]9~֪2�"O�J��P7���r������"O��b��P���P2^��!mK�B3!�d�>g�i
E)fA-�C�H
�!�Eup=`�k=C��7`��!�$�D!�P�5(7vנ��ST�!��Ŋt��x�G��`�b�h2탲1`!�$
%` �  ��   ;  6  �  �   �+  �6  �A  'K  �V  B`  �f  �l  5s  wy  �  ��  ?�  ��  Ę  �  I�  ��  α  �  S�  ��  E�  	�  L�  ��  P�  ��  ��  7�  S  � �  �  Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�� |d��"O
`�(�;���8���-0��1%"Oj4��ND^[��"3/9�0|H�"OB���H��*�ʞRy=a"O�味V�!X��!&F�:J�$���"O,��a
���C�Ą�M�"O,$3%o�-���p���+Ն�:1"O��ݢ1����`���y14]2��i�<�6��{_���c�H�`�fX�$Kn�<��A̼VI�xR[�)�Ć�pඤ�ȓA5��('nߡ4�� �)˩%� ���,��r�؊b#`T�eT09���ȓ!�b��g��}�8�F��-? �ȓ
K|m�ș�VṔ���2�%�ȓ"R�X�j�4JN�1�˘X�i����̹	_�jZ��1!g��zܶ��ȓgil,*�J�
j�Ne��i�J%b���f	�(U��:���G��$Y^م�~r�� S�%T"���k\�jx�ȓ|4�1�îJb��@ӵ�ݩn�V��/[`�"�v4�R�!ʎ<��M�ȓ`:��z�ؚh�J�Z��$HY:	��H��p�m�C1��!��B:��0��EnjZA V;9����J[
2���	��4'J�EA�IVW&��~�(aZ��ӹ�>� o�Y�|�ȓ�f�A�
Ο7�H��M�$�����mޠP����/���ANXo*�ȓTv�����{ ��-7�*h��I��sB�8�8���3����ȓNe*M�悡;������X�o��!�ȓ'lj�#F�m�+R&;�|E{��Oh"pPC�}2$�����x-+
�'D8���$9���0�]V����	�'�6D
�/�/%�a��jA7Hb��	�'����R��/����.��@�P
��Q�ܙ􇈘�HД$K�_�D|�q`,D�ԑ�� |^eqQ��\n�#e �<a�4�OQ>�S�GEa a�v���`%�tR	'D�<�E�sY�u˥�7�z�[�#��w���	����3��A�%Ι����F�$D��x���u�,�W��p���#D�D��fG�k�l��8�FQ0T��>I����P������0�&C�,�ȓ@R1�ׯ��I�F�3��EǪ�Fzb�>�U�	�"�rA��?;��h����0L!�D��.3Py'/Þu�r���I� ��)��H�0u�ӕH�*}D�Z1t�0�i�'�ў�}���
X�z4�ʇ�RX�&�R$�O`6�<yc&+S̊��s��)���˦��U�IU�@FP6W���Ї�B"	���3g�)}��'M�D�:o:�2⋒)�ec��N@��y�	�0�`�H���YN>EKB�ԾdD���� ړPU`@��F�c��IZA �$G���O��س@��n�8=�E�$j�du�$]���<E�����K�t���rr��"�Rćȓ9|ڬ���5R^|ĸ �S���~2�'p���B%��tHD3`2U���wL�C�	*�e0f�D	c+� �e��� ���hO>)ӕC׎7�>����IOB���O'�������[W�^�_�r&f��x�80;��d�)�(O�O�I�ǣMAn\�B�ėG�A�
��� J����0lBʙ��OG%%���`����Ҭ�mn�qB(<:���f��y��Z�X��d�0�D �T��?��>H�d9F��||����]M���V�#�㨟�H�N�����U�T���K�"ORh �E.JYЃ��6S�O��=E�t�Q�����M�
ju���,N��yB��a��ӈ\������T�y�A��?�ڭj��BZ��U�ߘ�y��Ӕ0���Rd�֏􅐷J�j���O���DP�tAV$i�(�>r0P��Z�j�{�';�	�&��2�T�C�GC<BZh�5"O��E��9(��]�-�Z<Jv"O����-�*>�ڗ�N�+<0LI��IC>U:`�V�Q0�dI��j��� D��	s+�{4@D �/s�$ّ�":D�8�i�4}��Xf��C���#7D�887���mH�7᝕v���;�`�4��	lܓHl��r׮_�r��g/�b�rՇ��y̓��x�B�G�(UYfd�&w����ȓ8�va
w��I�L9F&,-B��ȓ]J���R�J���(jNS�%�^�'�̆� ���8]
c�\[d!�|�x�'� ٩����	$R�0q� m��e�b��7��{�!򄈸t�L�Kac�: ���'�P�����<���'��'�噆& 6���$�c,��	�'���[��P�5��)PF � b?A"	�'�n�����,R2X�� @�p�`����ēM#�)�'<Q��Xn;xaNBH�&j�.  	�'t��A�.�����Q���f�LM��O 6-3lO!AH�=����Z)`+�0-�І����yb�Α:|�=8P��MM
�R��&�y�/�7?���SeՒW������O�0G�$�þ3w����	
����d���y�I�7��B�/��7 dP�c���y�/70��q��FʠG�z�B�,�6�y���.���1g�V��
懿��'��ϓ^�F�{3*�.�X,2���r���'���9�1JŶՈd!4[9���7D��*�W�6���ʶR?�,��K7D�K�a�(��������XXЂ'?q�O�O�gyBg�(z��)���	��b\>�yb(�?��-�ҩ��ļ;�jč��$�O���d�/	 ���ѹ2�l�'g-kI!��T�&*�L�5l+`���G9":���'p=�����:2�3ᄭJ��`�'azR�|����0 f�^t1�U���O�'G�%?qq�qC�Q ��"\q��edӪ!x�xB�O?7�֥l6����O�<,{���3e�	H��H�(	�!ʒm�Z	�V�E�&d� 2��yb�D(�0�]����L��%���4�'��n�P��x"l� f(4⒁�	��lA��'4�$���Av�҃�ӳb��l
ŇXO����<	�5M0P���b4n����T����?٠��Q����j3xzB��dh�<i��X8(�����H0>�E��[b�����OY�D�F�޽MҮ�b��,YI|�
�'��@K$�F�A~��c�$[b��Ɋ{�k�m��uG��D��N�)C0�xQ�� ��L��*D��iugH�o]�5�q(ُF��0"J%ʓ2��x�	�3=(L�+EF�M��Z�L���O�"~�B�˔R��Y���	�@٘��Ѧ��]Ĕ�f���L:�OP����ȓC/�4*�}#�DZ�hv�T=��S�? ~�"�.M�	�H��R�6;��3�'y�'�>L���-m�*@:Rn�~|�9�'1V�����T����1�U�{�����x�B��i�>e��I,�v�j&l�!��=��{����|eb$P���V�F$�Rʘ��y���� �I��ןD|J��B�]9Ǹ'ў�������3 řl�~,��'W^�<yT�_&*�t�A����C�rM�Sj�D�'���D���kd���1ڮ�j2��$CbC��R�<<��H�4���D�#��C�	���H!���*��t��2uZC�ɳ��0͍�C�BFU�VC�I?.W�{V+��(�D@V/�}�B��1��~�	PD�"z:!��lΈY�ȓ!��Р�>}���&'�U�~��hO?YД�E�|��e���U%��H� -:D�d
�/Fy��89G���2䂸8��4D��!�cT*�� 6��6O�nh�f�4D��´��O�1�c �(�:@�D�2D���a
�nM����(c�H�)��0D���1�KtT-*Ec��1����.D��a'-�l)V�� ��8<I�e��),��'�S�'�T!�Rų\�(�a��1Z�j���j���p)_��n�)"�W),��x��9<щq��i�(X)5mM�l(���	���7���@�,RC�蠧F\?x#��ȓV�a�Ԏ�9 �����lO %��">r�:�jyr�#�رr�*�����5�⡆�b�	�R�E�1�=�ơ�>P�<�ߓ!֦)�T��˜X��c���u��ɯG	: �ɒG��8���ԟ,ȸq����(�C��=l��C�U� P!�W�Y���=�V�p���}$�3@Wf�B�*z�|�*1iYV�<�"��gg����-
wTi��aWI�<!����p_��
ՍI~�r�ه��F�<�U
��ZN�`e^��ά�u�V�<�T��^B`q;f#/]lL��N\�<a�ګrd��+�A���H���Z�<�A ��vc�N�C���0-�O�<!3��7\-��ag��q�ziX&k]L�<�5�4<��P�2Mfa�a8�!PE�<yU�̔tjYВ��) �=('�I�<���	~���a���<�|��&K�z�<���SW |<��a:xr�%	@ϕa�<1��*@ ��
�ϒ�\��Հ`�_�<��H~�M����-\H���S]�<nڄ�)a�F�V�2d!qZS�<��&����R�Z�$N��tnNP�<Y��M>#�D`��G�1����W�r�<��S9H#��;3��pw0rwn�y�<qRc�b8DQ�"e߂
#����d
|�<!�l^�Y�L(7M?.|0ȹ��t�<�@ͳk5�<��i�?eI.��Љ�t�<�͵KD��3�ȽU8�M�&n�e�<��Þ�쥨F�O���Kr ��(�C��;�vt�E�W�`B�����*��B��.1ض}��7�Z�9������B�I9sঠa$�S0ɈV�)ueB�%128��OO�+���� �(xS�C��i��My"ĂNيQ��0��C�ɟRS4��-3xe ���C�I�C�IYڔ���+R�1h���"!@�ejC�	#�����ݬg���i���)=PC�	�F�������[���BS�\���B�)� � ׀����14ꐠ� ��"OP�z�g�H�i����31�.ˤ"O�t�I�(D����肚A�e�6"O*$Jt#�?b�(@�uJT�X��aa"ON�a�cV�u'4����Ж4��8a��'>��'���'���'2�'�R�':���]����h�i�0Tb	"��'���'���'�B�'���'?��'�.x��O(@�����\�s����'f��'RR�'�2�'���'i2�'+1����7���*���*��+��'���'���'���'���'��'��R2�	�FQag0^���	�'���'���'�"�'���'���'�BpP�M��gR��E�Ժ$�*%XU�'���'}��'��'l��'�2�'����W!R�H�P�Ej��`W�'���'��'���'�r�'��'�n�(U����t��p��2{�h!�w�'T�'Hr�'�r�'�B�'���'<V9�(ɐ <����\';	���V�'�'+��'�"�'�b�'��'	2��k7�aC��SXy{�'�b�'���'�R�'���'��'�t�k���R(\��o\j+����'�R�'���'��'��'!B�'�N9���:%8��čU�����'���'��'(R�'3��'�R�'�2�z#�֭&�ٳ`!�tK.5�'���'m��'4��',�
r��D�O����ؒ$ut� ��r7TE�A^Xy"�'��)�3?��i�*]Y��Q� r���y�*�񦭒���
ͦ1��v�i>�	�)�g��=(#�<�u�⅏2�M�r���@�4���yK�U1ւ��ӱi.2�"�]�,�4��W�)�b�0�	Ty��S�S�2�0V'Ҧ�P� #/[�T��4�L�<!����'
��w��rn�n�r╃.0�Iҡ�O47�c�����s@r$y�4�yR�Ĕ3���y�H��0QJ%�"E��yr�K)tݘ@�Q%�> *ў�՟9�d+g�Xt�U��p�Y`G�`���'e�'��7��/l�1O,L�w�߂)��U�ǯ��HtQE��O��OX%�'
B�i��d�>9w�H�����Qzh�K�BX~Bʋgg�Y�N�	ҘO2�A����H��I�'cdl�S&�PTA��*X�,!x��'��	ٟ"~Γ+�.�8��s\���(Z��X�2�v�!���[�����u�i>�uF�k����P7:^0����X����!���8�r�l�[~2�0���+B�U(�����b�T�)#��+�bC􅇒d�$t��؀��x2��6JKPx�&�G�L����Q��?�2��r��C6E�Zd
�)���fSf���C!Z/l� !ށS<�<�����#��APy!���?m�И/44��O#a>����}d��B�B�(]�̑Rg>D�q�?8r�*�&�7In1C ��a\h]�`�Q�ԕ��&����7�Ɂqޭ�F�S�9ji`��	s�LXPf�}�d�82#�	�民��̏I�MQt��U��$p�/��[됤S����&�V-E�Y�F�����	Ɵ����?}�Sɟ�;BLُ<5�ʇ��'����
�#����OxA[E��O���O���1�����O|�)�G�� F��{խO�sc�� ��SƦ�aF"�4�M;���?����Z�'�?����?�$�^�M�t��B<����u�6����V_|�O_�S�ɐ&�����t°4�M��7r�E)�4�?����?��B�T曖�'F��'_���u�`�y Ή����M>J�84ޮ�M;J>)t,��<ͧ�?���?9��!��ybD!�N�J��DPX�G�iD���Yq&7-�O���O��$�d���O��$�("HP'�D��Ad�im|9�'A�y�'���O;2�'�哙7�%X����M��Y�EE88��@H4�\<�M���?I���?	�^?}�'pB��P�;�n�$P�^� 5�J> �
���O��D�ON���O�˓x8=``8������4P>�xcw�^/?���e�iw�I㟴�'v�'��g��y��C�<q����9M&<�!햍4~� 0�)���?���?�梏g��6�'
�ʓk�N��L�?0Q /4fϔ6�O����Oʓ�?��"��|:(O�`���� �p����!bg�����R�WG���O��$�O�lP��Eצ��IٟD���?Q�r(Vd��4�o*7\�芖B��M����d�O�LAV<���$�<��a	�%F�y� �td�SU�C�NdӸ�D�OuR�*_��	՟����?�럈�AgnIBp��jDP@I��G����?�W����?�.O���S5�*�O�<��E�^�"}� �1f8�8Q�4u���sv�i���'F��O6���':��'~��v� 7W@XT�f��n���Z�%mӸD��(�O��ı<ͧ��'�?)D��*w� {ql�2w�Ј�`8/����''��'%D�{g�uӴ�$�O����Ol���h(r�f(����f4a������iK�S� �g�m��?����?y��8���N
! nz�H!/Zқ�'Ȃ�X��m�P�D�O0�$�Oе�O��dC. �n�s�)��uiz���L�~����q���	ԟ��IΟ�Iv�=J�$i""�B`���3Guеi@,�M����?)��?	�T?ٖ'}ra�(|cf��v��\���c�	β ��1��'���'��'LBY>������M3c��d~Bሶkli7*A�.�iq۴�?���?	���?.OR����e��I� �d0jc ;D���0$�~.p�':�'�b�'3rOX;Hj6-�O<�d�eD�ҢY@<�h3`ԑV�ΑlZş`��ǟp�'�������'��P�?kܭ�0*
�b�ۦô""���'<B�'���A9��6M�O�D�O8��͚*�Y�f�pWB��`ۻ���o��0�'��C����|��M� �8�p�
F��+w%עg��{ѷi��'(�p#��z�*��Ob��������Oܝ!6+[��ވk4g�i߸|	e��_}��'vJ�i�U�`����O�N�%[���"��%	D�X%o�j���z�B7-�O@�$�O����P���OV��� wﲠ�P��l��5r���n��)mZ%~�VsӺ�D�OԊ 1�ܓ���	�D�r ���!P����fE!7��l��������Z���M���?Y��?��Ӻ{���I��݃"[�G弤�H�̦��I|y����yʟ��D�O2���n9��X�N�>����,�5%J�lZ���J�a���MC���?����?1�_?��"�
��(��"4Bq��H2Eb��A'�O��D�<���?�����$ԭV�8aڴ "	�E�c
^�l�>�A��f�I��|�	]�	}y��گ9dPВ򩉽 *��d�
{����y�'��'��8,��8�OO�1"L�0q�nlѴѱ(��\حO��d�OΓO��T>,��'� PR"^j �d�X +�1��O2���O>���<��c�T��O��1��9C�\������ c����?�$�<!v�Nd�F�"0�d�ΗBv�I@��ˏQ)�el��L�Iy��B:`�������b0CH0R��أ'��
�%A�IZ�	ry��	��O��>Q��1X0�At�e��.w�6�<I� όE �6e�~����2������}�Z	�#ȑ*<5&�T�l��˓ s�YDx���IU4[����[+I,fyqw*Ö�M��ӝ5��'_��'t�4J �D�O�٪A.�/�H@!��6�d�c�ͦ�`�7�S�O���A�(.�E���֯g�])g&��k��6��OV�d�O����^����	N?����@x8Ai�)�/H ����I[�?����<����?����=�O�t�h����(Drֲi[r*RO����OJ�Ok�ؤ{�,�H��f�	����I�:H�	��t�I��`�	�@�O����$��"�&}���;J��kT�M�I��O����OԓO�ʓ:�\ʰ_�OJ�L�҆I9M��b&�c̓�?����?�,O� aîW�|b���,x0�Y	bH�:
��ǂQ`}��'��|�^�l���>�Q�̝s��639r])d��X}��'�r�',�	�E�| �N|:sGF�%M�(#eD��U�l�)䞦l9���'��'���&{�b�trs'�(5bA���Q��JL��+e�h�$�O�ʓ]$��������'�t%φ~�-�6NѝTi9�(�t&O�ʓ!��Fx���<�2��g��ò�E�}L@Q���$�$�D<mK���'����)?Y�lİi�T쩓,����F��榉�'�:�Q������4�Q�A"8E���δ$i��!��-�N6��O��d�O|��I�	ҟ��!#ƫx{tq��J���D*����M�2k^p���t�DW��J-)5�C�!5��8C��3hx�1mZ��x�I���V뎌��'+"�O ڡ	��Y��C�ٻF�4�B�d�	?1O����O�D��f(~%���ྔ+�e�F�l��p!��%���?������C��G� �q� B/4f(곢	E}2�����'���'I"S��
�&djځ�/�6R��7�AZN<)��?�M>!*Oٻ���i��F�Y#hV4�1�̑X�1O��O����<q�I�GD�1YÀ	Ѣ&+���(��;44�'�R�|R��v��>9w�	#;�$y�U��s
���ݦ9���P��ʟܲ���ɦ�ڦ��m��߷UP�W�C�>�Z	���Ϧ��	b�Iqy�]���'�5ж ѐ<������Ɋ�qj�4�?�����=y��e'>��I�?����� �Pu�n�~H$�pM���ē��ٶ���'HA<%q� ��@�@!D��VdR�l�gy�f
�mG6M�I���'>�� ?��ˌ.���E�S�(����Ŧ��'at����4��'{��Z���'�Lq+d�)�R۴4��B�i���'���O�XOL���2)X��M�6BUc���|�m�_����?�g̓�?�t��u�fH��6�4����Q�F�'���'"TZ�f"��OD�d�O�ԉ2� p��"1�X�sRt�0TA�{��*��?����?)��?����8V����FI����c.Ϭ���'tY��4������_yZc�� �DÊ�V�&�S�eQ�B��
�OL�p&���O`���O��NC�=�en��qxZErR�0+�y�.�9�'T��'S�'U�I�YP�,���;0�#=P�P����\�b�,����P��}y`X6X�t�%Jnz�{�+/��D͖ ����?	���䓡�$��yB��[OzT���H�f	А�7�I�P����?i���?�/Oxp�',�Z��@�5ڵMB;2�d&�<�5۴�?iN>a,O�Q�������x ���f�
��r!��s����'�\����ѵ��'�?������S�Ȟ)�̤��/0Z����5�xR[����b �S�� g�6�I�"�����8�oM�M,OD�����������������'�9�g���j��k@����ڴ��D��{�b?�a���jA�p'k��Ɉ�1�j��4��-ئ�	�����?�K<��U�8��*����� ̏>
b<S��i��s���ڟ�x� H�'�+j���,��O�Z���i�R�'���O]DO��d�Ol�I3l�@���g]0dv�lEk��M�Rb�4�C�>�՟��	� !J�2��`1��!K(�+�.��M��0�n���x��'�"�|Zc���x!`
(D�Dm1`�"+�� K�O$Z���O��$�O4���O �$�|z��z�Be��o#��zT+'kڨ�G���O��O˓<[J\�u͐��0Ƀ�a_1�J-�˅��䓡?���?1(O��	F A��X �"��n��3C�4��cдg�fO���#�$�<�4Fy}+�5�"��	�*0Ӣ}�@������O����O��e���2��d��@��&�%.����'� s+R7m�O��OT��d�6b
��Е�5JN��S`�2Û�'�RY������ħ�?��'r
�%3e%��t���)U��G����xB�'�(�J^6/�81��ú���4��$��Z~�oڲ��	�OZ���~"��B���#�61$�I��J���M��'�8��!�87�`|�5��\�����48�)2Ҷi�"�'�B�O��O���XA����կj�)�+Q*<2&���I�,�,A�\��Xaj]<j�I+��F�M����?��s�<�(v�x�'fR�O��2��ӱZ����L`�d`��'A��'Er�-n[!*�n�z��P�?��7�OJ8᱅m������	Y�i��3D鋈��+��oC�ԛ$�=��?���?*O@��7��0i�hC�ڑP����[�N\�T%�<�Iן4%�8�O̱����6u�9�p�O VTh�����O�D�O>����A�<��$[q�E.���wfč;6t��&\�,�Iߟ\%�(DyRL�PQ�Aԯڊ/��r��L�����O��D�O0ʓy2iƕ��+�`�L���m��v���"F�`�@7��O��O���$�h��0�N�j����	@�����'�B]�0�Ӌ�ħ�?��'x���#T�+|;� ��Ε���� ՝xr�'�X�YG��Pkp@�G��8D<=��4���H�}�m�����O��	N\~�
(��D8�F�eU@� �.Y��M[��?���P$����L<)��<A�l;�*[�o���ߦ}�pn��M���?i����5�x��'�� �ɑZ�,[����sr��V�i��m���/�i>c���3G9��A�'�S&ʡ%I��tA;۴�?	���?�EmS-d�'��'8��z�;!�ӗ�H�c��A�	��b��U"�I���I����������m����J�M+��:��u�d�OX�Ok��*�ԭ��D۶����5�����	�f�`c�D�	ݟ���ny��\P�U�e��8�<���X'{��a��J>�����&������p!��߹
nx �t ��6���8�m۶q�ܙ��sy��'�b�'��	�R��� �Oy�AZ�a�e6*	Q3����C�O^�d�O��O\�D�O4I�TU��8�O�&>��;s�O�)W�� gi�>Y���?I����DX9Jh��%>��� z;
�����A�F�1��X%�M�����?��1%�����L��a��4X�x0��*sJ�7-�O����<�I��u݉O���O��s�#C� �%X��"p`b<���OF�L)`�t��Y�(�
��\'d����fɑ����nZEy��C�L}�7m�n�t�'��TH:?�&�^���j4��QB��o��!����̉e
؟$�b?�xā��Nd:ݳW�F==��)�d���$���]�	�0�I�?q�L<q�d��qF��1^���/ϥJ�r�J"�i���'�ɧ����͙^�Re��c��G��\[���,�0m��H��ߟ �f�ē�?	��~RL�-BX<����i�p�6��M�M>�wMۚ.�O�r�'Fr�P/m�p�X��T����0!�؞X�6��Oˠ 	q������IV�i���T���e� 5���d@�>ѕM_ �?�-Of�$�O��Ķ<Il��xߖ�2r唳.� �p�G�A�~uK��xr�'���|b�'��Gx��U�F:�*���CV� 	�c�'��Ο,��ޟ@�'�hQU`p>}��rLX�P/�� �R/.��OГO����O�yJ�2O�ۤ�Y/
���bΎ�*S Y���J[}��'V��'U�ɜa<�yjJ|z�˅�s�!BV��?d�$��A<F����'��'���'?��!��'8�y�5� B�Q:�sӈ�
d�*$o�����	Vy��ץWg��>�d�>5i�d܊s�BYh���U�\�@�[m��矼��"e����i�~��$[N`��WI�Ӗ�i�%��ݔ'q���l�D��O���O��>� ��׹d�B�)u��
\'@%m�ߟ���~�h�)�9�t`�f�frf�����u��6M>l,4�&ꀒ �J���);O��H�O�zd$a�$�1L$�"O�*��¥ )�T�&�ߘ8"i��L�(*,�RL�dV�=�2���+=��kc�ǯ4��+��ؖ$7R�Z�I�<N�3$�0̤-p�)3��s�d;I�Ƞ���mjr!RB��<�As��$����ǤR%)���0�.]���Zs�@'�zD;4��J�(�0B@H���2í�Od��O��������?��OO�-�F ٹu���!��N�ҁ�Z$6=T)U�~9|l���q8����� ���垸mM��<
�~d�5��T�Z��М��|��K�msL,i�3�%ob��E
�;nT@�PGINkX*PH�"�П���4P�'M��'��Ov�I�F�;�90�G��3`�1w�'��'�$,���] M3�1æG6Kg�i��yJx����<qv%OB�������M�����n�1�� G��I�-]V��	ǟ��'e�"@�1cQ]������"�M���9M�"���I�2�\<
e�N8���#�� ��r �e;t%�3�]^�Dzt�S����u�P�#$���iE�t��pf�No+��}�!��џL�'�IZ$�1t�bmS�`P�&�a�y��'�"���*Y%�@�C6�u;�'e�6���Y�j�D�[�`۫GS��<1Ea��F�'R�^>}�����4������F�8\���[l������Nh�*S�|�f��%C��-˛.��˧��h��5N4�(�*_�tM2ͤO� E��*W�~�����w5$Р6O�_�eSՉ�:��$��e|J�yWc�9[ϼ�ӂ�_��s����F��1+�4�?���DED��X��׈!�x}��X>Ә'�R�'>�	�3�L��%��˙�8�6�J��i>qˌ��Z7cW�C��+��Y6ōm�q�v%�O~�$�Od+Ҧ�^Z����O����O�u��4�,�� �9-Î@��/Os@HPgƢJgp6��Ϧuj��^@I�b>�O(�D'R)bC8	(����"ƴd@��^%wt�-5f�P�= ���eh!R!��U/��S��f�mz޽qt��22��Qd��p)�	���H#�MKV��[q�Oq���'wRMH�K�mH��
�|KB�E�j��<���O�$�	k�I�2��I!�HO����O�˓`�4�6��EA���g<g��y7�ނs��\)���?���?&����O0��Lfy�1�ף+�`�Jb� 5E�1@g^�"j�����K�����9*l(�JM�Y�t� B��L4@T��3��u�C"�}�r�J�t���Q�m@&k��D�Ywy�	�m(�(֎��]��YIZ���Ek�sB}�Qm��Ȗ'g���U�L@�H�UIm���`F�3{z!򄘞w�.��6�Dq.a9�AZ1O�z-�O�ʓxɊ8�c����d�O����`E<T����`�	%.D4���Ov����2[����O�擬d��%Y���<h������ym�l�낊.�N�rp���Y��|ڧ�'ix|:�̙5$&��0z�l��	"�ɚ��ŵw�	�1��L8���'�O���<�(�
D���H�)Ir|��<����?����)K�c�0��T`�y�<L���ٍ7!�Ĕ���K��Sv���VHDh�iE���ԕ'��Q���>Y�����&b�����^J�pb����|%ʋ��r���Oj�b3�[�H�b����,~-q��|�*���`Cݥ1i@	��B]*�ؐ��>!P�H�=�	 �!Bw,��� !�'5�v8���5<���0��T��4�OVE)��'��'>�I�ZA�tr�ō3nA�!�e���1O��/<O���D$��*381	EA�(lO�@�'>*#=�i�?`���R4g�Mly��a�#��&�'�r�'D*���'��y�B�'�B�'^W���;h��cC2{�½��$�4kuP8���jF6�4�[
=N�p�G�I�=:*̣�'�N�s�����v����ܫi :US�ΉW�4("ï���OuȑA����q��&r��(a'!9��x��L%�M�c�i9�	�+���,O��d�:y�(��K��p�䟛PZLC�=k�ށcǁ�3o<��DH?w"����ʌ���.���d�<�U�K"T���q�k
*z��ҭU�A @��@��?���?���X���O4�m>9y�φ la�)cZ�7����b���H�d fFӫ!~�{sɅ5"�X���H�UQ�� V��'�P�B�/<�U���G�i�5ʢ�[2S~%�s���������?�HO��Ф�Q�@FX�	�h�6|������H�$��uӬo�埬�'����q��djU�)�4� s������X�ҵ�C6���q��1>+�@�<������?	-O�2�Zn�t�'��!�A]���@q'�LW�V��s�'���q���'G�)��$��1o@t�x��'/��8�k�z� ��I�JڨJ�lO�cl�?b���a�-`����ʖ��y�1 \�N�8����)OL ��']87�m}B�33����g�f��U��B����'���'�DRĪ��/^p���D��l�	�';�7�ǔN`��D�9��}��@R�*x�$�<����DA��O�\>Y��̟tAU�w�,��iA�i��ԟ���#�lq7�}�`���O$�.��ʧ'�Dd��PY	T�8t�"٥O�-#�.�$`�ła�Б}48��1&���ra��S�	o5��!:)�1���?s�l�9WM�+7��Ɏ~��$�ЦE
��i��"��Â�3�H����*y��s�34�Ȃ �� TV	s�k�H��d�)Oj�Gz2�&tU�p��J�u�����"iF6��Ov��O q��0t����O*��O戬;� �!!h�CR���`��^0� cD�%�<�0D�p�*��2m=1��'��]Y'���i��J��m]r�'��V:I����R؀��&#�k�\�p�)��)D�T2�T���� k#��|������ձm�Hpj�Y�m�,O�a�T���O��O���ei>csn(����$�61
�"Olq3%]B�FE���)T��I�.?����(�M����D�h���RǍ�Te�I�KG�e!�֍�z�j߹xI쐫�)�=YI!�?	6tH�$���hqo.i>!򄗅0=�e�� �5B�>�y'N�1'�!�D�-0Ƅॆ�m�tѼ!��.<��9��o�	.�DYW��(�!��o�yX��=����d�!�G�D��#f�<�~0C�X1c�!�ē&EFdkЧ��F���o��6�!��ڄtC|Ur`��yD� ���fi!��D�%y^���'sJ}Ђn�#=?!�Ć�m���j��V�!�D��ph�a1!�X��¢�˒m(��1.6!��zj	��W�M'̭2�Mƨ&�!�d=N�t�{T�ۻ]����ҋ]�J�!�Dڣ�2�Bb�Е.�Z��KO4S�!��V@����c��y�J 'WJ!�$��7N\*'�T�$A��b��;&!�U�⢽:����r���U!�ϕ,�r4���T�x��e,�!�dЁl��!��d�9�#*u!�D�	^Ny��Z&=�,8i�"�7f!�$:Ҡ%�$hց ��E�fH�!�ެ*�,�0�ȁ�	�}0Q��]�!��Cg:e��!J�(�r���A�	"�!�d�G��a�gI�q�`�RoV)�!�$&� ��kOg�6�E�^�!��A@i8�_�$�PV^5!���D��u��,"�"&~��Jv"O���l�~���	i^�Ka�$�B"O�H*��F&��0��Mx_�TB"O������o��E�5���^��<��'�z�����=�F$	=���观#�Xu ��p=��@сCFʩO�M�Ӎ�$Ψ�y��	��*ذ�I%B��U�r�		�Q>��.��R"N����V�`a��&�	�m�ac���.<`Q?�+c�K2�4r�"ؖc�6A�e��rv��#��Xw���A?!��PW�b��4D�b�b#��?HK6�z%þ<��O~��eG�7�� Ȉ�d�/l����3	��bc�J�z�����Op1b"�u,�\&��'������ S��s����l]d8�r)pE�,2�G�z�'N�tR�I��l��.}XR!
��H�Rx@Գt&�,n��!Ӄ-�<)�L-k'���$��L<	��og�H
�*FXߦd�p�ǡt~��>�u ��aþ��&!T�X�`|�����<4�éIR�E؁D�/!S�����"Q�<�-Q�=D�6�[�S���r=�%A�}��Y�ۿRB]���U�RJ)��)�5o����$-�5�^4�%��X�Ïl��\���-���;D�D��B"^���y�A4�<����H�,^�hU�u�X�H?Zi�?1���8�
<;�P4*\��@�oR3H��EP�G�"=�ā�-9��Lh\w�Q?I�F���z��		��Z	Va96Ɛ$.d�9�c⋰P��Gy�'I�V`;2�`��12��VJ�ܘ4�2AȼKF��c��cٴ;�0C�'�S����ϸ�*��� |�Ը0�K8]�B��
[�9)Ф�Ʈ���HQ��D��u�'��,i�M�Oĝ�!+�$"d��i��RV@��L̹_2�O�)�b���k���@��AG�/�4�dN�`���TM��+�t�6@ÁfT�r���U��M_�OC�<��B� ���|r�í� �c��������q~�@E'/�p4xS'�-#� u�1h�OT]1v゛EF����@�k���0K�5#���X�e�Yu�t�����3���0���Z�#1uZŰ�"B7@_�e�R�W�I,K�"u�Fz������[�N}s'˄�@(Q�*_�_�~�	���F�"u��g�I�>��"@�.B
@��Lk 둮Dv�'�Ҕ�B�V)����~V�I���ó-�/ �
	�5ʞ�{i~��.��)�B������OV�k�iw���)LY�6���X�a,�"�J8xwh|1'	�R��d"ɒ�l����s��73`X"��Ҭ	�$�R��}2!�'.��yܘ� 5$K�J��t���J�|��I����va˵ y�0�0�_ Q���+ٴ$��#�dZ=��yJ���{0��#�`R�6yK���O����ʧ$�v`r�ԙZR��ab�H"%Y*U�gH��!m�x�'�%P��B��yF��'�PAvY-d�����̡�?y�$G��ӌM1H�,��'�6�!�9� * I��8G� �M�;�����	�?rTB��%0� *� ��'J,��A2�A�eq����./��������4�';�e���K�c�lI�Dp��+N?��H1X�҄� �2�}�R�M>+���!']y��#�Fȷn%��i>����5���q #�V�R���bY!'�]qe3Or!iQ$�:��@u�럴�s$�I�&D�	2g�k3�h)�OW_�UkFl��\�%\�p�'�(]�~�ҩF�=� �҃@MX�&�Ǎ��mj��� B}�ԣ>�gB�?\�ͻz�&�׋ظ)Ø!jb�3-j��	Ay���!hO�)�ɠ����d9ֺ�8��.����򦎺TAL�Gx�"��=�t[u �_�5�]=�~�'	�E��&n4%�as�T�'��	.X��Dr�K�;	`Y���`8aj �
�o� sH�<1�p�-g��UA@��C����h�8-8ԗ�c�!����'#�66�s�� �)[j�Q��L�2$Ad;O
ј��֮P���ɰ$S����Iv�'=~�0��´V������C�\���K���(3�.Mi!�x�\���GO�'%K\�[raŪ=g.��VH�s�`P��E�e�V���� ͓�9��a���H4C��q3��V�	r!�E�'��	��&-��ħ�?A��\l�r�"f^�Z�@��Q<��u�>ғwN�7'Q��``��>u����ݓ���+�.e"�_ U���TY�Е'U���i�
��F�B|�R�'
����xWbmh�%M�3M�?'�L��s-Ʀ&��P��L�#Q��q�¤�ֽ<�.O���r�ȫ}��8` ��	E�p pN�L?��#94N)����3�da;C��^�'!.0�B�[�/n�͘��
7��A�#jt��dy�X�|G��% v4�Q��4�A�snX�J��eO�=E���G~���3C�T̻!i�=�4�Ē����0�E��!�O���?�*O1��$ưtl�YhEH�8R�d�
܄&�N��H#c;h�Ԃ��1$��f�I͌��'�M����H!3ïM�pp���X�(�'��.K�4)"���v���b��n�j�)S�%�a�D��$�]鶇Z�F2�YF�	tЩKV���.����I&T�0h���/f�V��0♗ 6�">�|Y�oӨ'��B�� L��Ey�h�$��唤%tRP�b�(D
�<B�'���f�'v��{�*���lh���J>!VZp`�!�P�'�,�aK�����N� �����mK�$YJ�A��Qp؟8��LY�U@�F�倉��N�pN�؉�D׮l_*!I'
K�2@DKa�D�B'�ɓD�Ă��>o	(���c�4vR�>I �Xh}0��	�vpKg/��$��ϔ;Z�	tU7_�Vd���pӀ��v�P�yn���CɪLT4H ���\c�@�r�>|d ;ӫ�2Jq������$ɹ��P��M]�q� �=����`�̉����Ҁ(��c��Y*�2�'�0y!���	8����@��=�Dhz��72,��7�'<����e���Ql��f4�pp�7gs�ш��?�O"��#�W���1eg�w�8�(�,_)9��Ȉ��W��򙰏���;23��hs�Y' f(��.Z`��O �����N5��W}NMRd%�krfYJ&�i��(�GӉ	
��seE�IĜ�Ϙ'�N%ZB��Pf�-Ĳ%ke��*+P���r+n�"�%I+�TX���auў�r�m	*V��ዖ�z�6Aa���
W[���h�8Y>h�PG�Ԋ@y]�mEEI���B�$�V-Փ���&��x ѳ�Z��#^��� ��l����.��O�8��]�'ݜ�a�jԋY1�DɣoA�N����Ν&C\�Ez�݌Xʢ�ӳ(S�X���^�a.�	�a���h��4 �	�q.̊S�Q��2'�F��@��0]g­:��OhI��{���S�F֒r*�PP�� �����'	U�d,;$��.E�h6ݟ�O`�bM�8q.�8�Ek\�����tƣ>qe�YcR�
Q�Άs�P���E�X�'�����%	@@��aXa�����D.�?����(��Q���5%;�zT�ñlA������(o\QQ�k���O8���Y^�\�(������:K�
m��D�@�'~
l��4�`d"D;��[%&ߎ�* "�_"Q�AŎ=�O�ٳ��ח
̾AQHT*?D�f���g.�x���������ϡ���<�-O���A��>��a��|���ċ�	w�~�[TJ�8x�ȴ�h��)8�rS◚%䈁3�\�) 8���O�Y�,�'bm��k�7}D(�֘}�
�;,O�[�h��L(��8[t���	=@�]�F���T��bd��:0��'����F�<������E�;f{�}P�B�e^���[{�ĸa�/�A�,�X��dՆ_��)�w��#��X�Kzv��S*G�
kf���?��o����
WY���'�J�I�/�!�bݰ�A��[�+�xe����HOfA끇�.X�!��%��<��O��aʠ��OZq���T�va�-O2�v��L�|���+ϐ9�2+F^�H	e�Ⱦ"��z��Ŷ�M��ț5i!��SL��P��R�?˓�?)5#V'ɪ��DJ�!��6�� PQr�y���O� [*X�!�^-ǽ�uקI�'x�uA#F �l��e��M�4���/I��@��8���OЉ����O�NE�f��7o|ٸ`ɳV���e�D-f�}q��'O����U�y7ًM	�F	�y�
��LD	�?���a�	8��d�<���`��22ɫQ�N`4f2r�<�I7�;;��8��DR�Z�@�0�`�<$d�x��f���3� V	Y�lB�E�a��B���aW���'����%�*-�� �o�`��/{+��S��%|�$,��
mV޼#���r�8]��C�oxЩ�b��B�z�#ϟ�	����>�¥��AZ;7�1a�l��M�E�Ozٻ���$Cm��`x݅I+�T�'*� Q��S=j��!ṆI�\��J2e�8�ӷ�����O�����OJ���.If��bE
S"�Ԅ� /n�UcBGN	��O0�B�(������N��7kR?��� ��""��'3&��'��Ipy��.�y���NA^�*1'�&]�lAc�'U�k=� ��	�W�|��Qj^:�؀_� W�"�(��Ff�;ӌ�7f�37l�XJ�"[�<qǾ��d�
�2�M1�F̸���&R\Ñ�I�}�Ĕڂ��8?T�c&��\��%�B\�m�ڍa�K�[쓶?Q�Ovr�)sGۄ5�ZTb�'�#AN�P�'��M��FO�
L�q  �	PB�� W�(O�T��*
�$z�������"u��Z��O<��%���|b�'���MK�U�
�������5��pҠF�P�P������o����T�w��T��c����ǖ�2��p�A�'�|BS>��_�ڴΓ{��[孒fp�3&˿@��!@��c�'�x�c��KmL� o\�?h��O��j�@��d����pg�^o<`���'�bS��� )S�<��+��$�6ݛf��;O"$�R�#��c%O�G�0�3i�H���dF�&��ExP� ��f�A���d��.�8�S��L�JnD� ��F��F����'��5��N�. �j%�tg��nE8�Q��$P#%Ѣ��`��.a��/�"�۰.@eQ�O֢=��MJ�
0ʨ	gg�~��� �D1�N���<�ua�-�˟��y'&M&� w.�?Y�
I��ı�M���3�S�O���]<77�] �.1�8 �C�d6c��(	�q���s���,��Q�� �d�
EE���L>7$�4��Ü�3����$B����;R�A�eFչ:kT)(�KS�w�@�/,6��c闡f5��ÆCC�7t@�-06��gᇁ&�����t�#lP�bq>-��hB�
�jHP�]�9��	5��U:SK�
&h*�S� ^�x�⟌�af�{k����� �K�Tp��ܘ��'"���O����󉍿*~YIA,Y�e��Y�'��N�����臵TD�Xҧ!��?�[�/л/����f� P@���!1�_���jUg�i?���~��ÏAM��JT�V�_Zq�Q�	�4�Op�i%%q�4�#A��v}k��x2�����M���T�u��w��I�<�\��'_̥��������־�I�G� v��!7�Z�V�*B�)G�e�^yIX?2èk᥂Dr�ZB具��O��O���U�<W�Z@{���7g\t¦GZY=��	�'8�yw�U,������Z#<�ĩ@DX�WΥ ���CԦ�L>1"��56$@f_�]��¦��� "��c��50`*"?2eH&'P�7l8$�����T���6?r���	I�	�<�WE)?wT &�ج.F� ��F�'���T����F�dgL9��L�#P��1 VG����'4�0"ROѮA�ƕE�$EM6��ǢA�9�i5��%|R��e��1��O?�%���St��-o;*�+E��?baASV��Y��"�Q>�:aܑ�r�E�y��(rT�@;]����r�����̒I8|j�V:Df�ه�ONh���ו��#��9uNX�ȓG.��#��G����v�|�@؆���=0#�ʷ?q�๶l	�&nF���hX����G��<ٴ U�G`p����乐c�W>b��c��i�fe��tƨ0U�6kGȐ׏�)zBD��e�0��㎎�q*8m`��#(����]+���7	F�'
 ��ԉjY�H�ȓ�b���7y8���T�y��&�nh)e���j����5O�����oD 옦"ֈj����K	/ 
=��	��z�V�"*��k�)zޤ�ȓ�����[�,��F��j	���ȓ^8�C�NW�V)г��}5��ȓ&�<д��DT&�A3L�Qzd��l�z`iw��u�<ՋG��#��q��Z�����SH��k����=���%+Pݒ�l��W R�k�&^ 46}�ȓz��P&��+O9p��QUfDp�ȓ7�XM��FƜy�Vp�V�ڸy����ȓ��r�Xl�,�fǜ�a������Ԓqa�/
2y�I��b���_��<i��^Ѹ�挥AV���;pZ�Q� \2Z�N@c�B�� ��S�? \��DZ �P�rGLmi�r%"O4�+T�O=_e"��G�
�6`(��"O������?����i]�]�ƀ�R"O���ðjE�Ԡ�.[yN樠�"O2��#�Q%�pu��C�R]R`8�"O�ԐVj �A�̫����	]�U"O,�����f�FQC!���v9uCW"O\ cbң@C�ab2`I�o��8�e"OZ���.���T��) @V�0c"O"�Y�;Z���EH/6@z	�'���)�~5�����Å|k�<+�'��%T�ۑXJ�Q�
�z��p�'������,]@� ^&tO";�'@@,�f	��ib��W�␺	�'�����X'$(L��NJ�����'9���ƭ��PȂ������'���b��G p �1�1?��$	�'�
�Z@�<Q�����m����'���)`-��O�����i���
�'RV��w%Y�!_f�c��F6b:f��'��$�5�I�M�BT�q�ʱ^�4�Z�'�������u2�	sa�܀h}��b	�'�rcآQ��hqM,_M��P
�'մ�A�"�i��}*��>a����	�'�H����۽)˖Ļ#옠V責��'br]v�
�X�$I �V+�M"�'46�ʱ��&8���O_�\�Z���'�N��g�4K��xh����`(�'�����_0x BE��_�H��'D���'��o�D��D,�!XY�!��'�`�&o	�k�L��ÃN�Y;�'�"!ȧM�7i��$��&'I�  ��'��H��Ȗo�D@a4㙚1����'n$˦�U$^������� 4�h�'�Ř�G	wv��l��1�:U��'kH��/Д�H�2�A4"�����'�e��
�=rH��gͣC��q�'>��=�>H �+ �3��q!�0D��b�	L��$Au%މv�D`d�;D��	�Q�tX�@A�װb2aؕ*8D���!֜r�x���)W!|V��!	8D�L�� N	&mn\�`�S	cV�R�
9D��E�^|��\��H�H>ěb$D�| W�L�� �� r5PP��.D�<�Ek����`�AY*<&$�D�"D�Љ���D;QBb����}0��?D���r��4V<i�/Et��"�I?D�d8SmN�c��x0C�͂/ẕ��<T��q&�L�C�ʩSE;]t�}�"O�mh��R;M5��2��7&�bK�"O. �ukɺ�h0��k_�T��"O|Q�'N�2�|��!�*xȦ�"O��S�,J��X*s���I&"O�٦O�>,�3Kŏ�A"OXY�4hR?nsB����ٱ�S"O@�3�	�g�2��#�ֵb�D�81"O�[�C�#&�x:1*Ӷ5��IC�"O<���@O3(��HUH�kd.<��"O�`(C�δoN�Q`�� OR���OFݣ2�Y�s�)�!�0'zp0r# D� 9���I*� �ό}>J��G�>D�hy�i
 =Q>m+&㈹_,p��� D����.�["��*Co
�y�(X!%*�1�S�'C[��GS�"Ja�d�CU�`t��S�? P����ɝ3���0$�X���9T"OreA�A[�$41 ˏ�#��d@�"O�
�\6'�<��$�Fy��uR'"O|`��H*m�����`H�"O��k�M�~ǞE��l�\��%k�"O�eQ'O�|�b&�~�X��"O*�۵ ��M�p���7t`�dR��G{��i�03���0�.�9�0����<%!�$��N@
w���T�ʅ�S�� !�d��+Z����1+ذ�	u��!�DѤNyP٢����h[�����0J%!�_w��Y��<+S I(�j!�D)SX2աӍ�f�(�A'�ʪD�!��ُ}�$(u֛y�*�S��N�>�!�D��go��:3�Z�B�p@٢d�i�!�;]�Bi�4-Ɂ0o�����шd)!�d<	)�,a���X 庀ƛ=/���T��
���<@tL:*�\h��`$D���4#�$Y�h�Ǥ��3�FDB�E!D�,�w�6	I�Ȋ��-NLzg  D�0!7�,8�*��E��r�����>D��� �G�'��㥩[F��*+/D����䏽H ���@^EpȒs'"D�T��D�W�:�@��{�4��M2D�TyJȀX��ը_?�R��.D��u/PEbִ���/1�D	���,D������Ox�q�&ޑ��b�/6D�����A,�]ґn]�.��`Q�'D�|i�/�,�r����2	���֡&D�$3����a��t�1h��PF
�u�#D�Ȣu�+[s~���K�Q(@F� D�p�So���L�Ӑ*:P�S7�?D��Õ �s�ZB��=ja�?lO��xy6bŅ7Q�l[� W����;D���X�b��-���g:D�t�4�P��!��'�
Ɋ��:D�tJ$�H�R F�E�Tml��%D�̻`��I��(�! �;b`T�7D�ī��4%�Ȝ9���;L��A`�6D����:t�����8?��,�g4D���fG�wo2-�	�#����`�>D�:�'�1�
ur��ߓ:�d���<����S r4<��oG��A�A��mg�C�	�o�$��O�u���@5iB䉡7*��vH���T���{� B�	���帐�ˌu�.A��*O�K2�C䉑F�h�sPfW�A�j2����Z�C�I�\@��S�X{6�Sc�S�MONB�I,=>d:�Eɣs�ܩ�WA�b(6B�	g8�ђjX�-o��F��13�C䉯O� �]�DԱ֌UR�#<A�3/B	%�]"�£<Z��ȓ	��݊f�G�>z!����n�ȓ[^z����+0ʨ��@;�Ȱ�����E��1|R�`ѢO�<RC��+x�Yf��N�FSR�ZK�<A�MZf�0xe��pnТ���J�<����B�4�;���epP��l�<���e�
���H�nA����d�<Q'�M!����i��a��I`�<����/K��|�R�I�4�����c�<��o�^/N!cq,�,B	պeB�_�'�ў�{'��kt�P�R}v#���+L�X���g�������b�3? R׏	�lXQ'(D�� 8�+h�z$ɣ	��e�u��"O��A��y�,l2U��9 ��8��"O″�
��8�>!�6g�=�\�`"O"���l���Z���� %�$"ODt��:&���G��R�捙�"O�t�f�)=��q��'���!�"O�`"����H؜ӐeM�+��-�"OLѡG/�;���棅�X�ƍr�"O���Θ�L�R5�0BS�]���2"O0���U�H'Ԉr�N|�10"O�aK�A��&3كs�W�\�Z��"O�T:d�2�MߗK��i0�"O6�����W5��ؓk_�r���D"O*課��p�T8�F*9V��"O\�B��׶�{�)}�Z����Z8��j"��1ID�S���nF�`ʗ9D�h�&�P�6����].��p�e6D�Dr��#|�d�G�۵6瘝�Ua)D��H�m��{���b�c[N��R�+D�8�!mژy�!Jt��;*����-D�d���,R!h万��G����,D��8G���3hz�5AY�QܲI��)D���Qɛ<2��%���%
������(D��O��=6t�PN$k"��؁:D���" 	'5ʉ�A�̎q6�Y���9D������A_f��W��7ea*�(�!D�8a�Q�yNΘ��I�-i�(��"D��NJDm�w�ډ�#W$?D��bթ,��̂cm�82��'D��aA�
%ILh��1yqjdׄ2D��X�/`���E�-M����o�C����0Wm��PDx�*b�ǫ`��B�ɨb1P�Z�&�$�v�``�Et�B�	?q�{�M�l�B��0:�B�'M�<yc��j�x'(9b��C�i���M�G��|JS��
�L@�ȓW;���3�.5.����ȓu� ة�|y����
�r ��,B��S-� ��b-�'=�T���x��m�:@1t��v�2��>A����4!Y~Q�FI�y� �'��2�y�J%7�����B��+����y���Pkh���*\�xa��y�c��b��I�	{�̨�߳�yҁ?O�ȑ�-I.|Zĝ�bm ��yIC�}("��Eo�-n�@,rq��;�y��{(ι! ���e`&8{cH��y�������GQ�a}z��"���y2Y�c��I�GĚ�|���?�y��ާDDA֫��O̘�s����yªX�FJ|h��< �
\(@�'���Ƣ���`��"��e��
�'�� �3Mɵ^�*�k�
��m�tU��'���U�X�V�~��0e°2���'t�<8PBQ�7Oh|���V�(�:�#
�'�8��a�N:}봙ɀLJQY|	�'l����ONV��@
�N�*T`�'��)�D*J�c���nD"(��� "Om�0+�E��p���J�4a�"O����^�<礥� K��HGh��P"O�i��Kݞ0�A�̺Z4���"O��('��`톼��أh�p�s"Oxp;��6&��-���,�h�v"O$��AZ�e]�A��/��*��0j�"O� ��+T,�;D��E��0��<�w"O����ɤ.���R͟@hN�P�"O��`#@�qŖ@�򂈝Ve�0"O���P�lg(܊g�%/>���"Oj��� P%Q��%Reه%�Bs"O��炀�?�h���;��U"O,!"�̇d��d���=OFXa��"OBH�Eo��Q)�`򔬆�[6L�F"OZ��JX"W��h�l��g��h�"O��*�H�!���KR- |���"O��a�/Y;TI `�5l޼�`"O�eHPŇ�$I��H߳X���"O��"hI�b�,���=O����"O"K0&�,kzh�&�#�i�""Oȁ�c�UsBB�UA!J��"Ol5���^�t�� ر݈G�uj�"O��hf"����p�^�Rw�KB"O���1�Q�,��U���G�vp� [u"O��&�#Pt��q�_<mRjIy�"O0,렉K�L)���gȗX4�H�"O��G�O�j���-�7X`�u"O�����[����4�9.(�"O.@BD> +J1;��l���"O���!7]S�-:��4"���"O�E�a�^>MDӰ�P��X\C�"O��z���%K|��c�/. ����"O�8ѵgǽc�
��W�*:Dd�h&"O>ܙ֩�<pZa)!��K1ta"O̭��'�QxZ�BP�M;;��k�"O�i�EM�������]R,Q�0"O� %��#&TD��J�2|GvY��"OX��O�|u�ph%�Z
~EH��"O� r�A�v�EK�g:��`"O�iYT	.K.�y2�K�d�R "O��r�XXjz���j��E�:���"O�i�7�,�m���T%$�h�I�"O��!K�2G�Z��Q$#�Ɯ�'"O���ݛ~�J$+PC�����@2"O� x�C�x	bᘲ0XY��"Ob����|�x���E{R8�"O�Su�ѱ*���&�T�7Ԓ��C"OV��`"�:8�}p�πt���ӧ"OFxH����p�Q�ˡF���5"O@�1MK> ����p؟$6B���"OZ���	���#���68�H��"O:�C4�М	�A�8��2�"OQ��ĲzJD����D2�A"O�8��k��2��iC�&���#"Ol�[Q��t�DAX�(�[�ιke"O��CL�p�(Úx{ ���"O2hP�'��ck�M��I�,�"���"O�1�oW�+�� 5<Uw�D�s"O�������飗���V���C�"O��Xr��.�ܳ$��)�p�"O�����
y�,9s�L��|�2	�'� lP���G|��z�CϿ!�N��	�')��ȱӞ?"�1�ψ b����'�$��Ё`�j�S!O��K6�{�'��a$EAͻ�bD-{.���'p�(R�fF�cu.|� �7yΦ9
�'px�K��c%z\kS,��i��8a�'2�̂q�Gd���J8���'cbP`%ΏN��Ёe�O6K��8�'N6���+ߨU�h�����WF����� �03s圇C&�8RዯbRq8�"O�A�p�ۼB�C�/϶4q���"O<�!��n�z���+�XhP��"O�UCP�9%G� R�K�UGT�"�"O
Iw���DQ��Ɏ0OEX��"O<t��ÍM����VYOr���"O�-��
Ѫ"����qI�_�Q@"O`
a�ӡ-t|�;6��:�Ç"O��2���k��XKħΫ:Q��*p"O:@2d+S(M�9�dũVO�aY�"O����D1�����?�h� 0"O���o [�dɲ,6{h�
�"OĬX$ݿ<�
��EL*w*,+g"O��R*.9T9[�*ߘ/[Tͺf"O$(b�J�~|J��ygx�bS"O�a���9yp)2�I��yS��e"O�9�
CV1�� 筄:gM�$��"Oj5��(`M�$��![��A�"OPH耄�;}� �����D��1"O�)[�ˠkn�e�� R��4��"O��;��_�o�H|��W�l�t��"O��RuE
�e��pK�to��J�"ON�{����~�4"&o��%�F|:�"Ovx�b���F��1.X����"Obp9Ӌ��kf|�b�5_�H�"O4��ggb�`Yzt�?=���ұ"Ojt*�.	�Sa���ό���z�"O>��'hЀ�4yVfE�<���cR"O�uj��J�NpC1�Z;��E;�"O$�S��$O�@jī�⨰�"O� ���H���� +�3|�84"O(��"Cْ&�6�k7#�)M(J�"Oz]�d�*B'v%!��0{!�dY-��Cbl�>G��8ʓ7T��A�u���
�k>d�2�A)+D��fOɬnM�EÑ�Z�r�� �$D��rN�9&-�I���&�Q�V�"D�����##P�	ȗ�Xf0���&D�$�A!�ƺD�t"�K�Τ��2D��S�	��%E~��o��v��w	/D�ȸ۱�^�����?k^����h.D��zV�uVQ�D�
����.D�L#�	`�Jm�G��u�؁��g>D���A$�%FuX�*ؘ��(�B>D��� $3(�,��[$
�|�8��6D�D+�)ǌ��}�eģp%Vc��1D���vɝ)���A��O@mp�o1D��)#�r������{�k��/D��[�1���r�lW	�θj�e.D��8�d�v��s�o�0op-��!D���.6�NX6��#��U"�� D�A/͂;�$�83/G�EJq$�1D����U_�����#-z╂�*D�0H�V��W�W�,z���h*D��[s�طedF�I��U) l\��E*D��4�/`,�� A��tVd�"I,D�X�Bk��^k��bQ�ua,hc$!*D�Й1$�Ī�u�I8E�j�JE�I��y�OG�|�v�Ħh��E�%c�8�y��D(@4�B�1]��0p�/H�y"��-�^��f�B!YR�v)���y��K�ApV �lߊQ6��Ư��y�$C	:u����� �D�)W��y�n�@	�EXUkՁKkޜ�F��y
� ���D�P�FcX��<@�x��"O�`�2��2;�|m1$��o��:�"O���I�4>�V�Pv�@�J�� h�"O
�q�/�xDSW���`�`P��"O�t�u��)��4�W�!�}&"O&i�,�*4��7�uc�yq"O�`���� `���F��B�x`Q�"O����Q�9��e�S����"O~5�%Uk6 �ru�B�"��la�"ODY�U#�<���7�D�K�(��"O �j�l#.�
ř/#�BH�"OQ��_�r�R���Ĝ�6	x�yw"O>��FX�lhs�F�*���R""OXyj[#l��4U�/�܈y%"O��$GϿ'r�����gU���T"O|��$+�,ٺ�,
:B�#"O8�ta΅Al�0�Ùe��J�"Ov�' 
t�չ�
ĕ�Pu.�!�$ơj@��G�>� ��_�!�$�"ruN�2a��Qva�0��H�!�ĝ.n���qB���b�+@
t�!�D�3��[uč�X�GL�Xl!�d�y�;n�uƦ�{� �(�!�$�}W�<X �,Q�����E>Q�!���^8��@�<V���o�S�!��ů`����fظy��ia�	,�!�d׍'�|<��L`W���A��Th!�Ē�Pu��R'�OR0�����\H!�,Y8��¢��|X�S���!��8r�M:"],#��q��R$9�!�ā#zB�be/".�XjaE�{!�#E�jٲ���9���i�ܪAd!��Mt��Ĥ,��xY�*A�~E!�0]JX�����fn�KV��#+!�]�$� ��)�?ZDZ�i�`!�d�k��`��
N6��k2!�dȺY����@H�@7&�k�K�6!�̙fx��t�y!�4��Dd�!�د}{���a£A4�@v���!�հ9��5"Ӣ\�^�����L9�!��Mʰ:0 ��9�b�p�
ǵ#!�dj�� ��#�11�r��Bp"O���G�1T��zt+D�m6��J�"Oj�q`�Z(0<�����l��!"O��
eJ�>A� jA�
�]�"O�8㱥K�w7�58&IW}�y;�"O��ICl'8�(��"0�\��"OZ��+	�"�F8�����ˢ"O��2V@� ����?/�섡S"O~���X4=� B���q�X}��"OP��		�q�.M���	�FD"Oމ��ȗ=2diA�"M��"O�<�!��f�-�#���.¼T�E"O��6�V$ ]�t�!�p�d�r�"OB�����&@�j$��n�h�A�"O�0�B�/�Ĩ����W�Ÿ�"O~�U�V�y?\a��&�K�Ԥ7"OBiH���?z�\L���w��P"Oh�KҀ\��	�fk�4h���v"OLM*GdA?j֥Q��%Kd��
c"OҬC�kX*�,`#o�5�J!"O'з}3�mb�X�@��zf"Oh<���#�P%��Έ%�Lh�"O�p���5�l$�a�еN�d�Ò"O� �P�ԉ��C�:�b4�\�#��q�w"O��b֫�3��Ą�6�\�0�"O� a�Ş}�j�A�b +nHШ�"O&]�R�~& ��v��~@�Ȼ"O��C�"�#�0�9g/Ӧ52L��v"O��b�)7�D�z���uv�q�"O�$�A�{n2�rSc��fpx19�"O>0���WB�.Era�AUE��%"OJ����Q��K��4d3�Q�"OH���G�1
��8�͗�+u<��"O�-��!�[?L�p*W/"dBI�"O��"d�N�n~��ѬZGt*""O�TȐa��1]�H#�i�� A�D��"OPT��J/rJ�����	�F���+�"O��X6�"�I��Hխ%h\KG"O4��ԥ�wi����� �kr"O��S��J���3�$���M��"ORѣ�e��������ڷE��Msw"Oµ+c�E�W���p�_9�$��"O��W�>EY4��^��$�r�"O�I�CLCg�����ٗ霼"O�)���R�H�Փ�[�S�z��f"Op�;& �"SW�Y���E�~�n(Y�"O����Q7���!��̱I����4"O�-���<&� Y���$X�t�g"Ot@�r-�/��)ttH�"O*��� Q�B�p��4Of2Q:r"O*�Jc��n�z���C�:G}�ˢ"O���3OL��Y�"V�Cd�P"O��)��>�����o(cT$��"Oj���xŴ�j��!;�� "O�A��K]�Rq~xwP�p9�U+!"O~�x�lϏ1�������$"OVI���ã>�~=���`���ȕ"OH�X��>���4&�1��mA�"Oh�����CQ�0�TC��8�Sr"Oʩ;&�N�P:b<p�P�+�("O��z`-
�7������ܟuM`�y"O��N��qXFtHC��vl�%�"O8�[�Α=UJc��$\.P��"OBHaEW[��+��٫SP}x�"OX�rrG���(��׶p!`Љ�"O�2Pg=+@D+�o\+Q�6e��"OJ��rm�k�h��PN��y�01�"O����'^�)�$�R-V����"ON@���1�p5���k@�"O��&$,��IS
��/*��(�"O�-b�Y(i*��gI�zd�*q"O�ax���26�j�0�&	�T����W"O���SG��"g$��'g�1&DT}+�"O��r�+�"͆����k/h�;@"OvЄ]�=Ѵh�r#
7{*����"O�T�q�V�0��ϕ�{���0"O�`�5j�?��8�PA�Sz$qE"O�tRQ&˦Vm�� 	#M��  �"O�������b"+/�xH[W"O�p�tA5&��Hɦ�\(3"O������>��5�%HӕM׸`�$"O��G�81f�EA 	O�@�@�[�"O2�k��-.i��G9����"O�E�%N �����ѮN,��I�"OL]���_��J��%7���#�"Ohiqׁ�
 �P�9QKR�Z���"O�jw�� x����J��P"O� �(S��yx-2q	��.e�"O�ds�G
>�D]�i��6h2�(�"O��C�G�OS�;g��
=ZA�r"O�4��d��7��M3F��Ոd"O��`�C
�M\$�P�1@c��"c"OPl�4VYY8hj��Dp�2m��"O��HR6N:6���@#UZjtk"O`G
V�(����DJ��+Sȴ��"O�1p�ɕ?qi6��7���r6��3�"O�2S� D���! G�.@1&"OL<����>0��arga��a>P �"O���)�t�:������Y"Vh��"O��F���k)N��OF�)���"O&�YF�]=T�`|���7��M�q"O�x���B���wa�;S�zt�""O��á��6as�h�o��Ĵ �"O���Ȣa�1b��.|�Ւ�"O��� ��W.�'��Cfޑ0"OuKu	v)� �V&L�?F���"O%B�
�&b�%+a�g�X�:"O�<k"����jm(��0Q(� B�"O�{Dbx��cb�8"> �"O�("Jǳ9y *�k�d8��"O�=��EA�Њ��+��0m�"O�#�ԑ>�:�;�J�fɄ��"O��c�Ι?
��1�dۡ2����F"OB���HB�tCR5z$��'U7
�@�"O���EH*<� ��$��BJ=��"O�1��A�!Z�ZѨU"
>3P�#�"O�X!�f����pB�/ډ9Cّ "OH��2��K��1s�`�\7�-;s"O����ኗr?lС��N�1SU�"O�ثr�P�̅���̹fEA�7"Ov�sf��0���b��<:��"O�)bp�Z�Eۀ�C@#��"O<��AƠf}����\$�J�C�"O�uq�̗�(ߖ}�T��'��x�"O�L�c�6z2x@ږ�K�t�Bh*A"Ov�ۣ �?,0 �ӗK	y"��X"O��q���+V��"��ŵE�]�"O:(��&M�+�(������쪵"ONyz�儸B���Į͢��Q�"Ol��EĹC���`�mJ�m�d�!&"O� sp)ҭ1kh��a��,F���" "Oޤ���%��2&i�9�9q�"O�T����C�q	K�:8
"O��	����6��fg�*B��au"OZ���c8t&]��ܒ+!�(�"O���H&M�M����"O�-�i�
0	d�HGl"&�f���"OJ���`U�)��1˖�Óa�X$��"O�i��I�. 
Y���3KڑPu"O�)��!7x\x#��a2�-+%"Ov8�5��4w�b	@aKO��A�"O�k��
Q@���
�?v	�L"Oz�#���b(���S)� 8���"O�5�����vD�a�ɉOd��"O�ᘆJݶ�R �5.�70� ��"O.|H3&C�N���[�4�$ z "O�L��Y']���LG0@y"`��"O<X'*�}��%�3B�	i�03�"OF�QCB<�Fy31'I�[o4��"O�Mqm�<���G�Z�w"O�rW�ܧN���B#ƕ�:W ��"O� �%����pp��!6D��Km�XA�"O�љ2�U \��,t�ʔ	��E��"ONа4��(�0��W�߃zԞ�2�"O�����6�#�D�,�!"OX �E�OzB@VNֽ�Z���"O�T�aQ��U1�C "\����"OƙSP%D����(aM�S"n,Y�"ON0�Ţ�f���p�Js����y�r��+7톑��5j�σ��y2kT�[Xm)4%��z����n���y��=,��}rF�-%��8�/��y���#���)�.�
p�0IC`��ybj�:Rz,!�!޹b<r����7�y�A3M(� XG"�7)�|i`�ˍ��y"�%o��k��Pe�mCԩҝ�y�Ɨ�8�\X��<1���CŅ��yH� T���f��z���)݄�y2�L�0P�EĊ	$�8@����$�yr-��@?"!��!��`� 
��yB�A�!��ZPۚ�Xё �	��y"	�`��8	�� �p��hk�"�y"��&n�����i�`�I��y����i�8D8fZ�Ā��/��y�.4���PЫ�?#���gW'�y�nK��ց�ϑ"9$����y��ěq���0`��#�+�#Y�x�ȓh�{�g�v(wf��M�ȓKA���M�4���Ͱ{5�܅�/wP����f��"�c�����Y=r��䁀,\��@�v�Ï[^~х�'x�c�7b0Z��sc\�m�0���!N�!ch�wB���
h�݅ȓ]�T@��D�
Ht$�ɍ����ȓ\BVL��hݘl�b�I�,
�\O���[�����H5/���)�*�mJ��ȓ#aHR�N=I�HI�fn��y"��ȓ7<���D�w�M��R�'�<L��]�ȼ��%o�xL���@�j+v��ȓU�Q����8�zy"�=,u�T�ȓYNv��cB�0 �,�BM��5�A��EE4��#��8`��Y���
� %��[���L�<��d@)�0�~��ȓ0R�C���Jta���>&4ȇȓd��	Xs#JlU����$^�.܇ȓ3����FC]7\��S��@��ȓX!6�Z`ƽAC�Cӆڂ-�61�ȓjZ81�����2�O;@�����<|�� ��vVh���:G[�ɇ�t�$-���.]��U�7\:[���cp6��8=������[��Y��ߢ�p��Z�tT���"��=�ȓL
���!x
u��i�6Nߺ���G~~��t�;����h���e=L`��Ǉ��-\��d�4I���V�9+N�[O��S`� ֜��q	�Mi�Х0�ak&AM�A����ȓg?4�R��%U��r$��1U��ȓv�Q/H8a�kCc7�,�����b��D��x	��:L�ّ�'Q���J�g0���=d�Pq�'$�H�%.`}�d� ��e��M�'�b�����m�0"\3i�dt��'����p)�TRиjS$�&_��ݫ�'��}cEjL%@k��jBV�"�x�s��� l,�� ��r��`�����-bl"Ovt
U�ّ?lh�2�˗7n��U"OJ��+زh �h%�
Y_�A��"Od�y�m\({T�	�R=^�� "O�Rwm�I��Aa�%��=�`H "O��Ґₖ'dir6&3O( �d"O�Z����O�&ۇ�׷1/\sq"OZ�"�)b�dr���d���"O�m�tbԯCZ010[�G	���"O� IQ�UW`��J-a��"OL	
����,�S!)R�>k(�B�"O�9���W, "�g�
b��"O�U� �6�>��f�$\���W"O� ��=*�&�حiU�Bp"O��Q6핻V�E���0S���"O8qۗ얗cn|t!��R@@\��"O怛���=Ynd�4Ƙ3]UT���"Op-8B�E�-�e	��Թy\4$��"OduY����hZ�T��)B��p"OQ5���X	�c��oE���"O���h �<����&Ì�B�`�"O�HE��0b�i�s�M5T99"Ox5���{�-���7/*z`�4"O��
"I+V�m�0A��mx@��0"O�E�+�<)H"��[w��B"OJ(` �^�P�A"�8{�!B"O����O�����r`S�O�L���"O���wf�R.�%� �B,�`�Q"O><7���y
m4Q� /[2j�C�	�J��ף6F6�jr����C�	�V:D���R�@�gm�USC�I6�p�"�N^#� ���(K���C��1��ȳ�	�P��M���G*�B�2ZX*b�Ж9�(ᚁ�D�F6�B�I�]�ȩ@�#-="�c�j�!ONB�I�&cD�A-�&_�饪��
B�	�cU�+O��%��' �3JB��J���� '	�[�X�sR�{�NB��.h��붂M�`��0�g'*B�	�2j�Y�uk� 7�^QЄJJ B�$}f�-"f.�?�pE�0.$�C�	��1��/ֶch�p���ŵW��C�	7nUl(�תC)�İB��P�C��6H$:���S���Ff�*
��C�	�.����sfl9BA�z.�C䉁pJ�2 ES�$�f�(D�ϿH`�C�I,�.��r�˾v_>��f��0j�<C�	?\N�pC�덧*rH�d���C�ɀU�Г ����B89�/��k�B�	�L�洪q��:{��p��BN�8~�C��?��������MUƘ����z`"O�q���K�� X��D h��j�"OxD�Wё0���#ƦVV�X"O����&
�V���irI�t=��b�"Or=
�^�H�N9��F��^(��"OЁ����lV�ݢ��؍�x��"O�,���A���Z�@ܺ�X��#"O�E��"���\�"E/	�#�����"OD�ҕ��D-�E�2)��ˣ"O���d�]="x2��Q|F�� "OQ�Y)c��  b�v6�S��^�<�NT�-��C�eϬWV��� o�<F��V}�tP�&��m��4
n�<q�hƻJ�6DP���C���y� g�<� \� D5!�L��FL�Ϛ���"O(��_	\�x=iEB�k���J "O�Ô��'�zы���P��*�"O���%��'@�F���ba1|�"O�4ɥ)H*�tH�O�X��1�f"Od�'�УO�Fh�p�_E��qk!"Oje�s)ă< $�[��������"O�@0D��31��(��	�37❒T"On��F
�>C�)qwK� Pl��"O8e���m	ڰ'G�#uH�w"O�A���I�v�X�`��,rhPS�"O0��g#��^�R���)_�-�"Olu� �\�\'~50�͐�He���u"OjUҷFW%t�h�k�oΖpd�p��"O6�&�@e�J@��o�Z�\(�5"O"x�� 
�6*����K��[��,�S"O�A��ۡ3��8y1�D�<�����"Ob��k�2Yn�9"�M3uN�@��"OF�#�c�7��e��ť%��ZA"O����S�5�,qk���1\�th�"O^�qD� V(��3ۿ9B4=)r"O�m�r�C!��H���S�i!�5"O:u
�ΐ5���FS�?��"Or���5��;!�!j�Ѵ"O:s���Xaxh��!� P�|�C4"Oj�9A�Wu�	#3��+�0��"O������x�r�W-\2(�(m�`"O��9�d�Z�����B5`f(���"O��	�L�t�t�lPc��k3"O�  ɉ>����׋�%6�@ �r"O�Tಆ���H����Z��"O���U
�������n�<rC"O��ԭ����I�H�+w�V�f"O����Ђ$rXi���1�X��r"O�᫷��6���Bp�Ǒu�Xrc"O^�����s�ؒ�C�t��"O�m��� q@}K"
�!jl��v"O<�3H��;e$bE@��>��!�2"O��S�_�/���w��vܢ�["O$�k��]�^�4͊�#�.!Ҷ)�"O�HZqIU$o�|��dK�4�^���"O���T�A`J]
6��)�����"O�=8���hh!遂	����"O>1�D�^V�� ȝl>Jq"OL�*"-ͯ`G�T[#�ьY�B=Y�"OT�����D)r	¤&�8}�"O���IKaV�e�_;iδd�"On�h��,��)C(C2��P[�"O�Ĺ�;d�l,����8����e"OL��/7�����VJx�y�$"ON Z��"m�dd
��7Cr%��"O�|K�@LU���K!�*Gb&i��"O��Z'�(VYB���<�2���"O~ �'��b"��� �μ��"OB4��aP�e��M�I
N�R=�"O�=Pg��nf*!�����` �"O��`�+z�)���P�p��m�"O�(�a ƛIA�4s�*CO�Π[�"O��Ƃ�J�X�'4o	\И2"O�Xp�N�.����Q�͋i��"O�ͺ��Ŕ^t`G#A�2+�qp'"O��	f��|�d!Pńō1����6"O�*)P�+l�]�J�%�2!�6"O���cMJ�8P�	��\��%��"O� ���a�;0-�����%B�2%� "OT�AVNM&9KZ	�/D<O�t���"Oΰ��FA!u
` ��� �4��"O�	����@��,�����0�V �"OHQz��Lhhұ��/a�Z�R�"O΅Y�H!
Z(�#�b�H���	�'��5��@�HR*�k�!�x�D��',r�j&Y
j�v�#@�7l9����'5��[�O5`�D�G+�ex� j�'2����C�O`��b'B�c7��!�'���2ׇH�G�b��V@��V����' �X���94��[A�еI��(��'�2�S�@CF������n
�J�'�0���¾S`�K!��dD�\B�'�$�k'ЊBl$�'R#`3��P�'l�J�h�
=��9��g��)�$PX�'2�!XB	:ƎPA�	(5��C�'��U���:R�Н� k��0�@��''�5�tLۼ^������*�j��'�Z�7��{c9�0 qLK�'T�xK�!ʦ�t�h0 �9�ب��'�����_)�l�I�C�"RR�x��'����6
Հ`N������5NN��b�'�H\�P��>�b@��EД3���'��yaІȀ)��x�S.��,2"p��'�"���nߌc���S!�4�v=H	�'���B��% ���M̖/u��#	�'�����B�~�"I��8�ء	�'�53 	]�:�Õ�_�@r�]��'m0��RO1� :%�>�F���'������l�<��"U�Z2��'IčAsg��^xn��3��'�(h�'@��؆��"+n\���ڛ.�m��'��y�E
����ICE�@x(��'�
xڧ�ȩ_ ��Ə�H8��'� E(e��[~z�i"�Й|.�Z�'�p'\�>rL\��ӧ{�Is�'�ī�H�!lX�Nݱ]�b� �'��T�f�\�E���у��:[�����'���R��Êr)\82D�=L$���'c�}r�
�-r`����S�2P��'�Ũw�F�>�"�0��ف%�h�'��
F�� �A�3)�la�'rh�GAPd�`Vl�+l2��'A�lPp��.
����P�Ǟu��i	�'Pp:�ʤ[�f�S�~
����'�6ȁ��ŸS��*ө 4{A��c�'s�hygСQ�>L�%�T�g7|�'ݖ��@W?gh��)��؆d\�H0�'������vq5*�NO/M]�1��'�"���2���x*�Hj�i��'զ���KLu11P�̆CP8X�'7�)�C`FB�6D"��ȋk����'�)� �8@��G�]a��?���["=r�U�
j$ri��kQX�C�Sn��zf��� �ȓp��}�ևL�k�$�zE-VH�~�ȓ����M��R��c`ή'[
,�ȓ 6!롬�yc�PI�M(M<Z)��f��H��� h��� ��;��E�ȓC�= ��OY�����ڳ9�rT�ȓ_Q�c�	0Mo���éj�(u���9)Bn�4D�0���$P����p�l��@eH��y"k3F���S�? vqʄ����:�B =���[""O�@[�O5�~��ց��)�$q�r"O�S�����@� �"�0m�"O�}�EV�S<��1�\�z���"O�A�]�l(��LZ�o��4��"O�TYU��F�fU�0!�;V��A@�"Oΰ�GܽDK�h��@݀y�N�K�"O��,��@�~Q �	>O�0�)A"O,�AC��M�����>Zĥ�"O�Cu�I�\#֋=;>$�x�"O�������\����e��Jd�"O,�1�*�hKfğ>�<i�C"O$��p��c�Li6��;QylЂ"O��aq��C��ea��/pd��r"OJ��a�R0��	�&����@"O�!`����	���*A~T�"O��BK1/�����"�9"�x��"Or��f�S؂1�7�OB�~5"O$|H��>/�}Yw�ȶ\8R�"O.�{�]�$�0{2�ɖ/�6�µ"OH��v��%@�&�a��o�J���"Ol ����/�e����p����"O^[hݕr�<��X��D��"O�%����T�ب7S�z����"O��ui�_����"0�ZeHA"O�<�w샎D����ǡ��V$�u٠"O&A�ULQ&CO���SN4��e"O܅#�,�)��=��4�B�QF"OB1�͞�'?b,��KL=7��˒"O)�d�FZ&D�җ�"�>��"Oօ���C23���GR�Ӧ	)e"O��ö�[6tj��G��S��tC�"Or�3!�-V̜r��ȩdr.��Q"O�1JW��b▨�!d(Yɀaҕ"O�e�!�ӊw�\�'�E��\p�`"O`� g|�n;6�(c� �90"OR�9c�Q�4����j_@�@�k�"O���%)�*�.��t��P�Y�0"Or�� הv�ت��V�q���0"O��ԦX�jd�xU/ɗZ�P�R"O~�jԠt��,�3.ƍP��"O�q� �x�����_x�x"OH�a�ʄ���P�-*$i2�"O
Eց��y-�Z@}��"O��a��G���lĊ[�HqP"OnhHENR�JLEˆK N2ae"O��(L��bw��+c:���"O
�{���Cd��
�j�Ea�"O��S�C���Aç>E�5ʗ"O���2$_.d :�9|��h�"O�y�!ٿc�TI1�^� �̙Y�"Ox!  .ʸ�"� ���t��%A�"OF���g�#B8�s� 0w�d$�g"OF�t)݌�t0X�"��t�^h��"OX�y����/�j`�
ȵ1��䲕"Ob�:`�[5mM��(\{XD�ѣ"OhD�5�Q�Oe8��'ƞ�y��"O,�(Vl�3}�4I0'�мF��qi#"Oj��`�h�������_��ە"O�U"���	1�^EҐ.ѵT�j]�e"OT���F0Hp�Ui����"t �Z&"O��Ƞ����a�����b�K3D� *͜`x:��E܁Z �Q#�>D���b`��:��8/��%G�=D�� ����~\����\C�("O�9��ԲM=��sl��H�@!�U"O�iر
گ7������ q۬<ba"O|���X}H��Hȕ.��`:�"OK�jK��{�!4<�J	À�V0�yb�E, "����	�.��4k'�y�nC�Rf���/W*\�@ ��M��y���(H�,�Bt��V��X���?�yb 	 6|<��A�4`vX�����yB	T+B��%k���T���gі�yB��	VeD�aR���O~V<3���y򭁍p::�h1o1K�B}[e�3�y�"��N�
��t�7=�(E�%+Q
�y2L/�]�`��4;��m2���y"�<� #�ř3z�A�Bފ�y��7t���Tkѿ==�X�Ql��y"F�Ob�8�.�2H��!JP*͝�y"�̡W��J���9\@���	�y�B��=R��*p)3"Ƒ��y�iə�Q	ڇ e �RF���y��<9��A� �5e���ab��ydL��BdؠD�)h�9:bM@!�y2�Ĕ`���t��2��4�!m��ybOָAl�h��OA./s|K����yr��#�hx����(1�(2��[��y�e[�kxl1�C��v��=:S��y�J��?���򍙯i�켒E�F��y�^1�4 ��g�Tme-Ζ�y�g�(&iR��#c��e�j�#'Ț��y�o� 
�%33'a%��A�O�y2*�*H�8Q�t�Рc�DCgۄ�y����4���L�Zr|)j�h��y�-Xh���hB�IS�̈c@��y�&вzG��#���m�����gP��y[3�����*;d�<���U�yRnS;{0j!IՎ� 9&�LH�e\�yb
�2g?$|�M�8��=¡]��yb���+��� `J6�\� I���y��O�s�d��!�D�x��E`��"�y�+ג�������\!��)����yO��ZT�B�L.f}y	8�yRN�e�ܹ6荺HY5r�F$�yb$�0��Q��<̎\��Z��y��xCމI�ܝ R���S���y��5��\��	 Gq|	���"�y�O�)�҈�3�����Y�2��y2F�yv��p�Λ~0�s��P��y�V.Y�h��s���~��ؑ��1�y����<w�i#��C6vWm��cݜ�y�D��iI�izNg��=0@#ˏ�yE�H��8@CmQ��J}S2�� �y���5�ʌ����?�Ԍ��gF>�yң��b; �
'���ĭ(�+@-�y��dy���P�S������ݽ�yR�ڱ	�!�AF>z�zt:���	�y"��1c�/k�v�r��^��y�)�V�x�8 !� cZ�X���;�yn�����Z��@�g�y��޲�Zթ��[5|����"��yR�ˮO�\�P�B�����yRJ]�l��1Q #� ~�H����,�y�?x ¸X�BєU���JO��y��A?U,%#&��Jf�]����%�yB��7�4-
��M&0�E���y
� �����b��xX2GC8.� �&"O�a��D�]V�j5�ƝLN�91�"O�hr��Z,0�[�C�4' X�"O����EITK�IԠ��s1��� "Of`�P�F�+�*PYwBW=P��%2�"O��yg��?���cF��!䔅A"O�%b�A�j��Y��`��0���{*O� 8��[�RSJ� $�Z:��8�'% ���RJ�(�B��;H��5��'�ȅ�͋%�&]�2D��A��s�'u�%څM�-Yp���U�@��$��'�&T�r�_��R��`��&�L�S�'o:I �C-Z�9`Ƃ�#����'r�yz��K�<d�f*̵�BT"�'HR=b5a�;�|�v��"���'M���7i�� S��2� �'C5*�R�@�����а[�'�p��JE�3:�"B�ν�'.$��D'3�U��-y_6Ms�'T�ћ�j��7j4\{A��u��	�'�:�U/�3+�D��h�g���2�'� d�QJܧ]�l0�t��]��P�'m�=#a�5H���Y�N�B���'ILY��33���Sǝ3v�T`j�'��ySb�K�t]d�"�Ո"�q:�'�����e��Jb~�xA�N9f$�0�'��u����p��B�\���r�'o$m��� rܠ��_�kǔ��',qK���9(�1�E�4�T��'��h���~�n�[�Ʀ ��tS�'�<�w�\;s�ժ1āk�u��'���#�ңf���ڀ��j��M�
�'���Vė�J���/������.D�,�M�K�R�(`b�,m0~���o'D�,"#Α0��<�@$0�V��g�/D�h��'��W��uQe�[\.4[�k/D�0�0�4+�1��ـx�^,�p�,D��!7"����(�4e�2B�<�� +D��kU->�D�C�Э|���-+D�H�q�
M��ᒀ��%&���x7%D�X���t�R�"�o� 0�)�5D�<�G��}��t��*>\!�5�3D���L�hh7 �;@O4A�H<D��BwO9�"�V�B,H�a1*OȺ1�ܑ��s ��CMnI�g"O�r�A1j�ؽp��6EI��"O*@q"��
�<�"�-@M!Q"OdZ��P!)�r��J��Ma(-8r"Ocʄ�m�x r�,K�#\tP!�"O����OP'\��m���Ӕph�Ș�"O�P�΅�+������B� (�"O�,#�H
#���q7I1F@(g"O�M���$!� �xV̀I֪3Q"O)�áR�X9����!. HB�"O��2�!�_b�����>/>I+�"O`()�J� /�5�ՉA�3@�:�"O������4�p����D��"O�;����c��I	f.I�>�@u�`"O�*�g��}P����J�9���)�"O�)��)�\����4չw��ARv"O|��t�7P[T���a��}[ya"Od �#c�O�rL $F��0�9"O��o8���ia�T�^� m	u"OD)s�㑣k��T�aĐ>���`�"O� ���H��m0������E��PZF"O(l��ν��ɀ���"��e��"Oh�zD*�0v�AP �]nY���U"OVL��AD����P'��/n*��f"O| �a�Q�#�v�C1��3�Q�"OQ�b�$h�&�4v6Ry�G���yraB"<�C3��>m|pu#Fj��y�$��F�
i�P�T�x�,�buF��y���L1����D�q�UA�BQ�y����%&s�ƅ�8�¥��Ę�y*ɱ#�\Ń�욙4G@Y��a���y�V�Lw����'̼�*� ��y�J�29$�uh� ґ�vL�5M\��y�۷]Pf� �k�*2��烘��y���7l��E3�����^7���yB�46~�Q�k�?p�K��-�y�ሪv#N}P%˵uB�a�5��y2䕶p���zg+C�j>a�fL\��y«Q(��R�$ô����`�<I��E�>�����R- �L���\�<I��<G:T9!�&N���P�D�<YcN޲-
��W�B�� 'b�z�<�#]:	������G`s�<�¥Z���e �ߏ
I|�f�I�<��ߣF�m+�LA�@�$4���^�<�g�S,Z*��EVc��M�Z�<A�%ڗ�.Y;���k�P�C�*�X�<a�E�-3���o�cK�q�	�{�<�r��.�u�`�[�
�!B��M�<	`���d��L���C��(�#��d�<q��U��\d�J/�P
�]^�<ѷ+��%w*���L��_�:`zbN�X�<Q��]�T��蒲�U�ZH�#"	T�<)V*X$�
�����E#��EG�<�R�Se���u��;B��ݒf��J�<��/_(T��҂,O:������]k�<9�,�m���aٲuD�GFZN�<QӆտCҘ|�0/��@N��z	ER�<��GF��R� Q�Q63�r(���E�<��Ј|�PD��H�k���YP�I�<�q�y����֯Y�k��Á�@F�<9�S�A��	i"�ŷ$���3��JH�<q5���Z�RT�QH˗,�P��)G�<Q�<�xp���ɪ1�Z���c_w�<)gaїv*���,��k�"a�V}�<IM̳E|���Ç�&j<�u�Q�|�<�"M��WG,��0(C�r����A�]�<����Hi����=������W�<��*H��`v��)Q�� BpB�U�<!U#֌Ciny�V"_�ҊL{4f�\�<�JD-Q�x���y3���N�W�<�GI�<��I��������pbX^�<9�� �P��a�'X^$̲��W�<���&Z,���˦f/�5�U�<�#%���κLN��AT�@N�<!���,r���;$o��UC�U0�BT�<Q�ꟊP�M1�n��KW�`��]R�<�
���:%a^/\�h=p@K\R�<�b�K.d�аsb"Ҩy�$P��c�L�<���JNq8���b��-� �b���n�<�R��9�X� B�Џp����QUS�<��%\��)@�2_��K��J�<1���"����A�ñ1W�xS��H����U��U�r``�(����NJ3h�����S�? ��CM�
O,�P톢T�&�6"O>���hE�d�pe�h�z��1O*��ѡo����C�R�{@���2pQ�D���,���Bv�|�!�����B�"2w`E� 
�?W���2��
0=�B�ɹ3��KR�	Jj�ȃ��@-��o�����ٹ��JW[��.Վl��`c@"O�,ڷHʾ,�~� �&óT X�"O`�-Y�|80� �AgE�C4"O~p�Rkaj�(�A/}A����'�Q��yu>E)$�����*32t xrl,D�x02%K:N���G�ĎJ��p �%D�(KäY�sT��39XJ椻�l#D��R�Ƥ~�jd��
�j����Ƭ4D�8���C�uT�*�!�&xC:e��/D��Z#�������oqW 8�O*O.�`2�#9Lb�ƓE�n��U�'HQ�8�w�I
�*��qg(E�x�+2D�{�#ʹ�J�8Ceϡ3oD��s�/D����JG���cj/;b��1� �=�S�'U���K�ǆ�v�
�0{�L��ȓ������O)S�,�(4�Ċ�謇ē�n��K���Ժ�@ܕ,�I�"Ob�riב2��`�#�&4+m���i���P�$?�x��f����Bh���4D�l�u���c��Ds�[{m>��e6⓳��w��ju\�y�Mè5��-���@k��y��i�>Q��&d��AaQ��5R
��U�c�<�mO�g�nlBq��Z75ۀK�<�E�9�̱�
t��d��!�}�<�f�  � nZ�
����D
B�<�G�\�:��WLF�h]�̉D�<���Z�v�H��jؕRG�p���@�<��f�-sbx ���9|Fru`��{�<ɠG�=u��X�L%���a�I�t��p=!bh>D�F�Ô�4_8��t�@K�<)�dI5(X��B�G�G������o�<�q*3}�h�G� =��8�Dm�<a�aT�l�8г�M�8D�l0�$��f�<���-us�=��o�1$���j��Kb��D?�{��4��7#x4�;B��&^�|��զ���p?Q�O���%N3A�+E7L�	)�"O��jfM)C��	*'u:
���6�S��Gx�"��ӡp8M�$aZ�;��B�	�6gXYbǄ ���q�J�f�G{��9O�q"����q��z�+�<�
�"O&��sEH%}�<�p$�S
n)Bt�'$����IF��Ha$��7b�n�:A�*�ZB䉱_g�Y�D�'퀥�'>C��	7�ȍ1Ю�m/�H[�
�T� C�ɾr���ʜ33t��1 '�;b��B�I7A��iB�ן	6�-�4�O0���Ms�'�'��<!Ձ,X�h,�w��3?3�)@mJH<�+��"���"�&�J���+LzD��F�<q�"bZ��bE(J�" ���c�a��H�'qO���u "�s�V=)� 08�"O,���b�z�="m�'N��U9�"O2���T�.���:��0����Q"O~\���Sh>$a�	����;0"O&��uN�6�6�ɚ%��sp"O�D��˦ygv@���ZRɜ�� "O�u��o�O�.K�[�]�����'q�1�=AɎ>p3��BU,�8&�B5h�ۦI$������Q����~9^��teO�7�C�)� BU�� B/N� �A�=fiH�"O|�^�ڭ:�S�U�bL#��OI�'���Oz�t�D'@>iAƘ-�xq�'Fv�!���;Fr�<�!#� Vp��P��-�d�h?�O��јO$�@y��A� M�U$
J�����	{�����$w��)i���> M����Cg��Fx�����z�x������͐B!*D��s�H ����C�]˺1�)D�0b�iٯ4d�Q��&ڜ)�b��oyR�)�'.l�y��$zZ����Єȓe��m�Aa��s��M��V�1Ӯ�$��F{���bǺ{e
�� @E�6�ּ��ډ��=q-O4�I�`����8G*�@�B�"	k�C�I� ��RR��!S	>�r�L�p	�C�ɝ}�f��q��)b���@�֪P�hB�I�{d���Kפl���9C@A>�.B�	�T�Nij5?�ΰ�
�$�">�L>)K~JF��W��ٗ �
t뀮d�'�ax��
��;%�%(���Rf��y�D5�b�z���X�$-"�?Y�'��؈��ʰ��
�H�A�J�:	ߓm��'�:|�eE���؄�A=���B�'�$�1Q��r�Aa��7&��A�'���:�S�gybi��<'�1#�ΧR|�z�I��y��P�^�QZ�*؋,8p�� ��yb�ێ5K,t�%�7���'��x�r�|,H�Ĝ?f�Z�;r/��EB!�"ONdyP�
R��]��[�U���|��U������0�BK��J1]��ɗn31X
�'�Y��g8��H�Bd�� 
�'3X%&�J2%݀q����5���(
�'��	�,�3ZXB�j���<��U�J>	���)�5.�>QĀJ/(ցj�'�Q F{J?��=�UF�	=vI�큾w�����^U�<I"�	'jjl  (�d��j���N(<��4G^��hS�Q
��"en�!	(̄�X��4ʕ�7?}Hp��z�(��ȓQ�\<��%��h�5�V�/r(��ȓ�M��IӤ@��vJ	D$��i�'Sp`KU���>Q�zc

�3 �Ś�'�R�`5�-F�������	��җb9D���k�a�<�qQm
�Fy��E�7D�,���A���h�F�@�8�I�4D�КP�܍=��a�D��?A~�ap��3D���3a:h` 	Zե�=F��u��+&��hO��d�H��0+�L-5� ��f�r6=�S��M�F�יK�44��' �p@b�Mu�'ў�f?���􀊽4���шՈw���F-��R6<v���@l�����M��d�/>°cr�^tp$�3�b�<�%O�g�hx�M���!⡒^�<	0º ���!��-�	�sf@[�<� �V[�S̚�5�ĘF!GW�<i�)ݦ2!�x3���O<蔠��]~��)�'V}L(�`��H�: �v�	m��!̓�hO?j��ߴKC�H�D�'?�"��
?D��j���U*�z��b��!���0D�l�$��A�t����CU�z�r��2D��@qU.�8 �IB3rt�	�+D�X�U��ά%���޵)Ӥ]`��(D��s����y�b0�>)���!Vc%D��[�p�V�rV�T�Ry�4�Xr�<ᒯP�{�@��S�G�lK�L�n�<AկI^�|�ʑoV�`�!��ER�<� �5CF����� DgҾVR��q"O��S�oSܚ؂C�� Lp$��"OR��w
Št�&���&'�:E"O���&D\�R��q��;t��"O�qC$l�$h���AN�+��1"Ot���䝃�p5I,Бz��pk�"O�lS��hd1SR�
Zڤ��2"O���T'�|l ��!���)��"O�)�6=���ҡR(D��"O����G�Ov��v0*!��"O6�ʇ��H���r5��*1�	@p"O
A�č� Q����C�.9��@"O
y�pmW�}�E�6�F�uHQY�"O4�����5@��Ƭ߮:|Ő�"O��*d�دY���&�J�*h�A"OB� �gQ�A:�-�� Ad�$�"Oؼq��*A�0�������"O�;��БI�Z5��J4wh�
%"O6���Ǯ&�bH�#+��oL�q"O"��T�߷<wF�����&k!��W"O��Z��ґ�i�b-���"O�xj�F]F$T$���M�N:��!�"OTS��U�>��|a2��`�N�"O�q��jI�D�urm�~-��$"O�0���>#�p"��N;�fi�"O�9���N�y<����L���"Ox�:t 4������31 �9s�"O��Bf�&��J�\���K�"O��U(J�mXa ү�3ʔW"O
���I8  �4����z.D9�"O�XA�!�Y����í�^!��	"OD�9$F2p�>��$
T+Z��( "O�ر���	q&�ږ��M�r y�"O���E�f1~8�����Ұ"O��1 ��b� �Acяo��#�"Or�s�BV?:(,4�s?���;%"O�8���S{�	��B�D>F	�"O����q��2w/�&�Y0"O�P��بLV(	"��ȕ@ �4�	�'Π� �ֽw*�%@v
��zE���	�'U�ac�A�,U�`��}O�E�'����V!շP� �AE�.���'�+3�Ӏr����5��l����'�$�WGˏn.����`�l��'S��`eo��h�αhu�\�uz�5b�'#R��2��#t��A����<O�<q"/J�2��E._C��V/L�<��.B
Q�d�!nQ�3�����L�<A'�iU�����N,	q\\���DO�<Q!`��#����(�"��  &�n�<�
�h^��#���>B�Q�t��M�<�RMȚ<�PXk ��� ���BWF�<�F&H:
@-[�"�>4^X�JcL�C�<A�H�n��H��;�F�C �x�<�B#:^�VDK���MQ�����y�<a3�
p�C�B���Yès�<����s�,h�&ԕBfd0XR�<1��!�|�H��Z{���;�K�a�<���@�>���ހ!�D��'�X�<��m�]��*��INT�C I�a�<aZ�u����`.P	C� I��DCW�<����?c(�r� �=G��,Q�<i�@3k�8ecR���74�̀H�<��,6k�	�PԈy˵n�G�<� ����J�4(� �D�W��Ű�
O��{L�`�����9\p����,�`��'��P��=,ΐ�
7���������z��4[Fk\�ħU��=�q�݅������|A��e��-�7o�k�^�D�;>�\-�':�T3��^������j1�䵒∜'N�RI�P(�S$���"O5G
4&����ߟ$�ԑU�p���<E��<�pF-��3�I��$-;tӨzX�試f�5Y\��$�U;l�d��(���a���,9Ҽ`p����MU�������^����w�'�L���ͥ<g�">�+Ѱ�ܑ�@�� ����,���2a��$�~���'�h�j�d"O)�#�I�Z��h!������@C�=O����7SB����������Q�m@�LH'�/��|��MPp�<���\�(5��Y��C�\I�
7b��
�ٛ��T�4(�5Ā/v.���O��{�'˿t<���*K� s�Ic��'����:���@&B�C�.Ũ4��$M|=�E�	l,� 4�'Ĵ���Mҡ&��-y%��Ba�����X�6צab$�2 �t��eh�|B��4s�����M=ͪAC���B�<��˨ys lS%�ѺYJ��t���<��B7Q���D�E����)��'ix���aΪV�D��1�&�!�$	�
^z�󃮉�;����6�������O������h���1�?#<��ҝ5��&�� z����i����"�V?L���I-%:��l^#e�4���I��h�H�J��'��ia� �4;N q��Q��9���d��T���c�=)ȟ��2�_?���5�%$�,�p�"O�,���ֆ5t��ЋŞdǔ��Q������\)�0�����0|��'�5B�� ��o�/^�����X�<�gh��(����T�|���j£�{����q)����g�NVj��B�i�
 �5�Y_Շ+4���D��=pN�e��bނaS2��D�[:H��B��W�x�҂�]��-�R(%pC�Iv瘍XW�\�9#����L-i�XC� �dM�Lӎj��M�Ħ��p��B�I�vȲ�1���������e'3�B� u�
�a��Q�L�����ǫNLnB�(}��1'-�*	@�P�"�B�,��%[�%|w@P�l��%"�C�I-�n���'cM�0���ѧ@!zC�I$f���P��+��j%��%y�"C�ɀ���R \1P��\���
a{�C�I=ɚ� `HS�4�v�ye��)��C�	#X�*��&���\�y�`j��WP�C�ɟs��3�Ǯ	3p����Bm��B�C@����#�6YHe���5@tC�	�R�B���
�=-&�K0^�,C�I64t���K(s�vIHũ�#y�xC�����iB�m^ �S�"�t�VC��X�BD�$�_�����ܼ)�C�9	��0Ж*&a�)�D�*RDB�!1eŇI(.1��f(ÇW(B�ɀW�z�C�  �GJ�5�T�]vB�	�$
��#���T-��;c'ԁ@�C�I]�8��_Kz��AmR,TC�	��0]*�L���m�4�STC�C�I�S��`nV[��Q���K�`�xC䉜 -�� Rn&d�,�W ���2C�I�cc�A�vAX'�����Q�qsC�I<T)3�[t����J�1��B䉳r>�0@�R2�r)��E[�5�C�	�j~uB�:c��`���<a	�C�1g- g$τ37(�J	�a��C�	qwf)��ۉA8"�J�O�< C�ɳ05���g@�E�0�ޘE40B�I+~��ɗ�F
31uk��P B�)� ��(A��t��	WǞ�@ۄ(�p�'��O$a��[���e�͆a[4"Od���싥]���"J����CĚ����\�S�On����H�O��)�mۑO�B�'HX����бE����"5
B\��y��'�y�%_�+B@��Gn��,��,�B(׃�x��'\���'oO�#�L����Z�"�B���OXa�v燓,�=��BʦHG��@�'��OV< ��%��0���"b6��a�"Oz6/�	�|���3\M��"O���5�0 �9��]�x睊�C"O���ڧ[������P�g���`!�䕇k��l*1�@�D0ě �O�xm!�ő;�28� @;*!�իcKzJ!�@�x xԎȕx�+� /E!�L�-�;ũ>%��+f��+!��F0�<�@��&|x��#�!��Z��AC.�C�>ͳ�*L'
�!����������3Hz�<�P���!�X
Hx����Y����b��!�ʢ18�H Ǣ�{�`�3�P�*9!�ϧJͤ��G���ؤ��o>!��3T<�ʢ��NW��G��!��S$���8��>E��y��Ym�!��|���%NN�{� ��A�A�!��U�K\��A1(Y|��a�3H�6Cr!�d�`CtjKI���6�Qu!�_>$��IθCl�Fœ�]���°bY �B���D}�D�u��5u���E �ă�Kܖ@�R sn<m�<tA1�8,O8�8D��� q,���N�΀��Ã7*��ȓ/9
	PR��4�4�P�_FP8�&�Q��=	�qO���I'$�j
�f�7#+�eQ�"O��+�P�raz�:&&B b~�: �)2�p1���L<���D0`)F��d���"�aH<!a�a�jL[�MPh��R-P�Y�|@6�&�O&-3��ܪw�ĵ��ő�W��آ#�'�z�S�c�	�#����D���š�S� �C�	"R��$��4�lW(+�ޒO�8�$,7�)������gI�p@t��_�B�%J����D�,�́q���q�B�	^��5P�瀪L֌i�ì_1�B�	�J�T⁦��r�z�R�`!HHB�&g~��j��S �M�gm
��C�	3w"���%�r�ҥ���E�r��C��>>F��`H�R��C�	̞C�IH�Lt�@L.!]�չ�'4B�	<;�H�h��k}��1�ݬJ,B䉚�hɨ�nܒ:=ލʷ�
�B�	6Vb:ز�I	t1F��l=�C�	�RC�a9��Ȑq~���I%:BB䉝adP�SȀ:�,�3'G3[vLB�.����V�T�69h�*���C�I�EIR9Sq�ױ?.N�jd*&NB�	�eN|xsHW�$�L�b�B�	W�"�a�L�LL�iA���:�B�	0~５鶩��ą E!I�0�B��q��l��Jk��qyuB(l�B�I#�D@:��]!�����nC�H6�B��9 x�-���-p��/@�&�xB�	��"����dQ�Ҋ=�C䉈|���`��$�4m�C�	�e���L_�ո�(��C�	>�x���A�_e*�bv�=tڸB�)� ���f�d�-��7�l��"O~���f��bW�]ؗNܴ>���"O"h��E	1I�Ѳ�k�]�R��W"O |�e�5Lx�u��M,(�}��"O+�T�;��q2o�NKܬzC �y�'n�*��ӕzF(���<��I1$��d�BB�4p<U#7Mϑ'��4͌�l�^�I#�ӵ������݌v��B���>Np}�"d�!�y��)yȮ����S�3Jb��r��>��D�-$����dɳ��za�,m���q��
j�a~�JE5�y���8dw"�7�Κ{>�D+p ˀ�y"�ԇ7t�}P���?A !��`���yr�%iFZ<ِ��Bt��ㇲ�y�O&g�ҐPcd�
n�,e�����y�F��"��mcCB1`\y��)Ş�yk�7/���#7!�T~�"ÏK7�y���QDB]�#CZ$/l��ǡN�yr�FW���W9&g6�W��y���|���K�"C�wEӦeB2�yG�p����3�����!Fύ��y�N��L�f$�fˑ�z	��E�J0�yB#��c �� L�{Ob�+d%�y�iQ�U�D!���.t
�,!�+��y"H?>a�Q{�͏�k�6i�Ad%�y�[(�A��E�l�E�@���yOΰ]9����*ށnX�% ee�y���.0j������V����臬�y���P���%�?v9�$�_��ybO�,�6�p&�T��T4W��:�yrᕗH4�\Jv��W����ɔ�yb΅�I���Cr�+A`��:7��6�y^: ��<���<>�|��o�2�y2�J�]b�)R���4)�B=+F�Щ�y�!��^��qx�$�=��)�k�ybnݶ{Zx��T�=�~Z����'�v�����G"T!�l�sHXP��'u���` .�����r�t��'�Ѐ��#� �$4���B7at��x
�'��rUD��0Q2��vK꼹	�'a.cR�V�T�|Xɷd	�JaX
�'5X-;
��@�p2@�b����'��xEnY" �,as`k��Q	��'F`���צs�zd""*�1K=��9�'��k��Kj��vGD�S�8�'0bY��
:\�܀j�,)N���'��d�F�zf`�����S��A�	�'�x�3]���@�ΐ���{	�'������8
EV%���FIl�	�'?X��!-�W�2�;�N�2?2X�0	�'����{	�����#^@yY	�'�vѩ�C^(I6�xB�Q�		,8�'kRѩ(�/��A����7 ���'�.i# �~C*�)c�Z.<�Ū�'��93� c��A�2`�x��'���5��87�5!�!�z�.!;�'Da�aDA./�VhK�ɐq\"�Q
�'���ǩT/`&�%�s�� x��p	�'�ޤ��b�/u��D:�%�T=i�'��q��B�-7��-r��	��X:�'/i���R�A���!�$э|�����'<z� ���1���P�<y�>0:�'��j����w
h9��Ѽ	~�	�'��x8E#Z1Y%�%Z%B�9T��0B
�'�����:�<�
�eĽD���p	��� ���$%]�ɓ�:X�~�Q0"Of�!6�D� vM���n��Q"O��WV�O�$�z��5Y6���"Or��p+�$)��*�ȧZD0XZ�"Opa�!�]�Dq3m��
��0"O,�2�ͭu���%&{o��&"On� �2�F�gU�4�"|�P"O�2k�#Q,	����@㰘�#"O�86$�3�����z!&j�"O*�� ��y�I��̓�\��"O�XC�FD��j����1�J��6"O651c"0q�ꙈУi�6��"O\8��]Q��T�!v�~	��"O�A��Ma�2��*#u�dMӓ"On`� 	�!�*��(H�j""O��z��!+�Z� ��2�t��"O�	� Mx�<��'�)<�:�@a"O�Hv R����Q
�=�%5"Ox5�Â[8]����P���Er�̃"O�HR ���������� _u"�B6"OV���j�&!@1�woK�LR�)p"O<�W@�P�J���N��6�D�p3"O\؊�$*F��L�$+��s�\�"O�0�'�%f޲���Kɼs��9�T"O���W�@]��H�߹b	�xi�"O�1�"�:p<Y�ڝ�Z�#�'R�-�e�E;s���2s� �ti�@�'v�e��R�(:��2�7\�H��'�Z���Y8TB�aҠF�|��'�ش�p�Ͼn*1W�=Ѵa�'됥Ƞ�ZZibD
�	�4�:�'�XT���$.���f�������'�H\R�iB�&���0�����䅡�'�j�z̀�M�4� �%�-���'��PA)���aA�� ^Y�02�'Td��P�aА���.��QLj"�'�P�!'�9-��,��a�p��|��'#X�P�b*���WfzDJ���'F��j��� �΀*�%X=v���	�':���A	�������M�'�zh�n~NŊ���	�rX�
�'A��@"�]R,z�uc��<�c
�'�f�YN��Ӭ�Q%O�-T�*��� ���@i��*�b�-�8�t`��/��y��*��X�e2.F� �Q���TUa���n]J\��H��>���ȓi�F��nڳ��@ʗ/=�]��9��	�lə'~����xՇȓfp&����r.F ��[9Ad�@���P4u�
~�]j�
�5p��%��O=�����ȏU�p��e ��Z����0��Xrʍ�\m��*���%�.��ȓS�d0��!ӨX�4oE�hb�ȓ�0��I�. ь@B"`�J;Hp�ȓuJ���ֳs�&5z�`�$�ZU��	�!�p�#	��%�AdǢ?�" ��Bh�[�ɒ�zJ�Hq�G�L}b�ȓm'�I�A�¬;8��ъ�JY
���Wm4�Ra�)]��<HфY�d���7�bWLI� q��UNB�č�ȓl�zco<"| ��NF�FY�ȓi,�`��Dlv5�r��KM��jZč8%d���[�*�?)�Ɇ�(ք�j�Rp��#�b��%��S�? �I
3��8�yb����R0�T"O��G��~�@�pT�\�9��y"O"�ڳb��zpHE�ޣYxd�%"O���%��E]��1C�=J
��"O�0���!���	$��$HP"O�D�bċ�ͩ�*ݘP��A3"Ot��q/_�)g������3�0��"O �R�λM h�	V�B�)Ѵ��"O�U	�*F�̅R���ע ��"O��*b��JV���u�\46����1"O�uSW�]IK�`��#	m\2Y�"O�Œ�G�5,Ȩz����FT�c�"O~1
��"��D`wD2P�˰"O8���N%�f�@e�^ĺX�#"O8i�@M�=�>,�0靐T��H��"O `��
	K�(8B3�Z^�<��"O�	Ӳ�Б,�$���d��$��"O��x-��9�Ԣ.A9 A��"O��k5�̈_��a���=��ۗ"O��Z�+֪Ep��B��4Ft��"OL��"����ba�P��W��hD"O��r@�5�x�A0�	>�h7"O��!��9L6��iр�*dx�|�"O�D���^xe��Ц(,xdX�P"OD��Z$=v���d̺4�ey�"O&l���% �E�'m�B4@"O.4�� ]��@�b ��q�"O�%���B�`1�%L^��r�"OX�ەf��P����##�(�P"O�vG�?�>Q�Qc����H�"O�����������2�,�8�"Oة����
�p����=X�`�"OJ	�6� �S�6�(d)v��;�"OФ�l��
��=Ae�ۙ:�f�)3"O@����C�Z���ϑ=7i��i�"OB�$��}�o�u[^Q��"O��&o̦����t���W^��HE"O����޸%%��i�)F��h�"O|�KdA��]��H�q ��"O����CH�f����B1��"O�H�!Κ�B�$If#ÓR6 ) "OH\�J��(�h�RӃΤ$�H�"O��X�O@5��ٲ�i�Ը�Sf"O�[��[ rHa�e�?�U@f"O����MF�e(��8�kϓ��{%"O�X�h�.wV��@��M�"O:;��К% ��E@�^����"Oj���!C� X���H�h�&�+�"O:q��Kƛ::�H�ECA�z�\ 7"O ���+��9��|HcI�_�vق"O��)B(�>|����&�Me����b"O�0AޛmĠ�)�ݩ�JaYg"OZ��#$�-X�<93'Hˤe~r���"O@�x����Eɇ��B�L9R"O*ܚ"	�a�����B�g�l�'"OT���G-n$j����M-4R,1�"O^ىWg��G��yW$�v�|��"Of���hI$�#%L��XhP"Ofl��(,<�BT?�#�"OD�X�RI&x�7��H�e 5"OJ�¥J�]KxT*�G�$b;2�� "OԤXw�B�m�1�Ӆ��?t|�""O~@PTl%�� d�h'� ��"O�IH�53��|�F�! ��""O� �0��/��E<�;S$�a4E�6"O(���m�N�4��㙳��p�a"O��	t�T���VB�U��+t"O����L7�&�Bw�>|)7"O�-��>D�l��CX�
�-�A"O
آ�+)�4QR��,�N��"Oܡ��K*�-ʦ��-����"Of���W�[.��4FY\��D��"ON��'X/(�}����*U��Y2"O��#�Q�n(´E�����"O��ڐ�D�*���P[2=rjE"O�]*�� ��Њ�n��^rZ�J"O^�"�n^TR40��NA�9��҅"O����nX�e(�)�fb�hpʰ"O t1�E%	<݉�C� ��1�2"O�����!E���*ţX<w\uY�"O
��Vۋ/)Zhe�?g|Є 4"O� �nG=PD�����DiY̸
�"O(��(W+C�"qǅ��AeR�"O։� �Xy�tEb�枺-<n%س"O~p�%�K\׾)Y���!>��A"Ox���i�2Q�ܱW�R��)��"O�HB�JMV��Z�ğ-(ӂt"Ob�2g�O�v�LণD=t�aia"O<(5@ݮ1$yU����I�"O�T���D>Z�$���b��^.,�x`"ORt�-K�.��M9WA@�]���2e"O8�x�+�1L����e��:.�l��c"O�k� �-!�Ӈi�P��q;v"Ot��%݃SJX؆�O�l�v�(�"OT�9�k�'b���3�	��-��xS"O���pĜ7�����B�/z��K�"Ozx�9 ���ҋ�2x�����"O<E��ᘤ$U8X�5O�A0r"O"�b �ªo��#r�,mƘP"O����4X��Pr%#�;mVH,�Q"O�Tq�b&W	�	�a�e��Q{V"O��(b� <x��20��u1F"O��B�f˜�����-G�0��"O��"@��XctKͲ>_���$�/�0�'��(��x��'�Mk�O�7�O��G.pD>ŋ�f�ZY��2O�
/O��=%>�"Ed
� 9P�p�i_�;��� &�9D��2a��^�P�{t�ǥd�$��
�<I��Ez�)�43q"� Oh�����TCƄ�	��HO�>5`�K	�t�<�I�q�R!=E�Q��[�';CT���dC.�p����w�ҥ�>!5�=�S��j�x���"�"<�P1{��L��O֥j��)��%׊YP!+ϛJ:La{��d�D�Yx�"<Y��)�<OQ�e� bG;,ECԡ�*>���	Jy����p跮W�;�@hXv�="H�F�ɤh��"�nѩ:;p��	_0���!g�Xi�+u��?�O|��-��LȜ���΄��1p䦈h��݉!**�O�=����R��Ts�X�M9"������,��F��j>�=E�$Ï�|L�D�R�EƘ�J'�M��/�I'�0|��M̋p�. ���̠eK� �釂��'y�c���eJ�O(���Ȉ3�fU��^;g���"�Oɢ�v�D�O��>�Ɇ�v4��ϚRc�x�ǆ���D3�?!%F,���NFp܌A�X�闎�i����'�dFy�����l�dn=W_�L[ԁ 8��6��U��ȟ���$��7Z�S�F�G��գR�I�0|*P��2&�.��ժKl��*sMU�<�����4ؔ�V��8��,ˇ��P��hO1��[�B*yA K"�ˈ��IQ�d~Ӓ�O��S�B�7+ZvuJ�`Pw)�0�왫3.�x�>q���K���� D�����2Pv�סN�r��a"ObA#ԤH^�$1��P*7攥�`"O��2�<>��0hֱ���Rt"O !�dnJ�}"�YS��>�}K$"O,���o�Y͔m[c��n�	�"O>�+�gVk^�t�Waڧ`Ԫ�J�"OJ=��F�=e������Tg_R���'��2-F�<[H��Nܡ"LE�'�j�@qD����o5�a�ӆ�y2�1�Dk@���r�b�yqE��y2DN0	�!KcI��q�H��P�F�y��Q���c@��5�8-B `B1�yR�@�T&걑��
�,�LPЧҽ�y��O*<0����ą�)�5�G&� �yB��/��u�Q��`s��'�yBM[�tV��{Ci�E��TI����y"���`���!���	���8�E��y����fC��{��T�rD
�yr*P A�p�C+ٲl���iЦ�y���_��ő�!��aB�5i�gL�y�n�'�3Um��&rz����y"ýs�ĭ��`���p ����yrdS�x�R��r+ߕH�ґjK��y�C5J���8���v�C�y��A�I�	ӁӜT�,�5��y�!N�(�8�����;�\5�%���y�ŗ-p�h0f�G��%".e8E�� j"`�S��EY��I<T!���h=���'��4<E[��\�!��3G6��!�%��?�x�s΅2j�!�S-\kV�P����e�^-��,���!��0c�ш���W��S�+рg�!�X:,ÚHS�ÄM�6����W�!�$�N�đX�&�74�|�2�,-v!�D]&I��P�0k�*I��%��HV!��=dͬW�a�J�{�	�369x�ȓ=����pZV雴��Z�"9��3�
�tA�!�dpS��'^��ȓV* �ۖi.7B��AG�	P�����J�D��_��@Q ���2�yz&"O`�P5)+7H��7옲s�yb�"O*y���F�Lh��I%S7D���"O��T�\��v��dj�"O@eD�B��a�ȽV�� ��"O�A���$;B�[��]���#"Oe(񀉾W�z��hؿ?�5j1"O(�� ��*�)���
K�<�z6"O��j��7 J�0�'@�[j���"O�y��f.��H#��.P�$yv"O��9��K��27�ȷ/B��b�"O��Ӣ�9y�Yh��_!@�1ѓ"O�q���0q}�,R���,�Y�"O���u�O\�y5 6��i"O޵ш�9}l���Nލ�b�q"OZ��iM�r�vt�w�Ԑj��ɠ2"O���J�؍�F�ɠ{�x�"O*�b��*D��Q�@"N���w"O<�[F��<&�8�3Ø|�eQu"O:��a�S/`	��`/ �Oc�i��"Ov��BcU@�������?G�-�t"O�-{3ɍy���)#-�05�� A"O��o��p�,���͇�%��:�y�Eg1�z0�S�� X����yBF�1�$�u�����i�����y
� ��r�>-��P�q���h����"O��)��Ք^�`��f��<�ڸ�S"O8I��+�
K��m	�	�+lpѱ"O8�A�Y*C}�S)^&[g��2""O�I9Bɔ�X�� "ӨƾyV tQ�"O���޲b���DhG�B��I�"O�(�4H��8�H�BE��r3�%I�"O���fǓ�?@6�I�%6lSP�#D��r�E'N
m���H�@�+��5D�\"�"�fݤ5�7��gF>�{F�4D��Y�L�@�� �!�ەK"e��i3D�����))�x3���!��%0D�� Э� Tf`[��F�X�����#D����ϑ6$��p�r*48�HII5#?D�R��2w��<rt�M����I0D�t�$̟�b��g�~b�`��g)D��8�-_�|���*T㗳Rtvɸ�+D�dkT-A�
���ʐK+c �Q�/.D� �1MX�o6�1�N:J�&E	�?D�8b�	R�|���B��8;�DP8�E=D�8�2 ��x�#g��r1X�3�#<D����!֯
H��ڷ �[�P��@<D�ء���7�R����ج'ˌh�� .D�H �+��dw(H�"l-a�>��-D����Ok�aC�O�0�<x{�$,D�,����.�}	m]����f D��Sqf
bt@d��%@*1t�s�k9D��s��E�W�|��VA��pt�}Y��5D�����1�
�[F�B!yq �u�3D�P����t�T�����nU�Aa��/D��J�эhVL#�=�J����(D��B�͂6���'�?�� �-,D���r@��K����a�5�J���d.D�h��%�/�*��V#�\��2�&D�0��H��p��Q����"m��	���9D�p��B�@�LVHcN�2�N<D��q�g[���p� L�=�L;�9D��8#j"�t���VZ�~�@p�7D����x֤��!�T�!�h +1M4D���霺)U�-R�$�$`��1D�d"�<6��� �Qa-ȠcC/D��ʲ��(�:h�,��4��,y�.D�88�h��DzȈ�"�(:j0�F�&D�4��SM���+rfV�ND�#/D�(c�H*{��5�4/�#\�����+D�����.H�	�c�gaBE��(D�0�!d�Ve;J��e��`0D�P�䊝;KD�QE�P�]c&)D����ǘa|$��P2�!#wI+D���D��:�$Q�T'{z�i�4%+D�dP`��=f�uAV 7����,$D�,��N,9I��!�J�rY��z�>D��y5`:0	� 򶈉��xF�1D��a�ҹ8���	���Z��;D�ظP��-xљ��ݯrtԐrN9D�p���2_R����N�R�u�5D�S�ŝ1;��h6�̛"ۄpQ�O5D�T�w��:q�h2T�E�n�4��4D�<{�
�Pm#WD�K-��(��0D�Z̛3j�!�@.�� ��賦C/D��PdSR&j(��J���h,D��PfX�;+�;�I$�����/D�p����B��u��i	��� bg� D��A�%_��hj�x���a��!D�� ����m��S`�0�1"��0�Qb"Ofä��0,��X��+����T"O��Q�k�$E�(��' �?��=��"O�@E�7{[İ�d(ۯq�t}cD"O,����!6�(H1��G,�\}��*O��q�5�J���aV?8\��'[V�y�J�NxֱIe�X��2�
�'� E@�JX"#82!
M��_t�2
�'�L�`�'&�&��Kڑ�J)J	�'/ށ���^9&D	r+�p��p�'_� d��=^h�it�\7k�<�S�'PL@���=����^M(���'4���e*Ёm��|!�-�-�j�k�'��&`
oP.��(�l��'�V(�6��NnH��^90P(�'�ι1��4U�PD	wͳX
��A�'����@�*��qA��d�8�H�'*m��
����s�A�)�ƈ��'�`{![b��р�%mtV48�'ߐ�qR�21V�(�B!g���P�'VVK3h� '�A�$��-H��	�'��	�S튛RT�D�̓,zN��'��q�dF?*1$��)�$$d"Ej�'�dRvJ�>� �� ��3�X<��'���A��	
\��!�#aʏ@�r��'��%AQ��C����[(I�Di�'k�]�cG��V�x�WC@�DD���'���N�+�*]�0�L�t�T}��'�t���M:���`�hREI�'T̍���)G���a�O��| �'h��H�,/�P%0!O��v b	�'���H�]� d�=�1�	�Z����'����I���S�۴Pc�8q	�'�l�Q-5N@� 욧u���8
�'�����A�T�Ѐ�ףl�"D�	�'dxXR.��ځ:��;5V��ȓ|e�Lxvˀ�2x��k��5#�$<�ȓV�����\�mSP��/sƀ�ȓ0�d��
�6 ���3)�ȓ?�@��
Y��.­Ƞ�B�<9�M�#_"̸!�̒m��(�ac�<� #U�����T�Cu����D]�<q4.� g��Svi�&ل�Q�m�n�<q�CG� S5;j�\�/�m�<�7#K�b��S5m��-�*�m�<�5욒r�BP/Q�&� �%�Kh�<	PI�5��{�-H���Y��Ta�<�tA4j���mI=t����i�[�<�3&C6P��˰��1D�+���S�<��(SZ��p�֯ͧ~��
Z�<�%ER���Sɕ�{�2M3�@WT�<aV��
(
y�$%�(rΨ �O�O�<���OLƴ	�f�Z��T�O�I�<�R�L�i��:�I� F	�q�f��E�<Y�ךY����M�sD�Aׅ�z�<��޴�~�"�B_ �Z��}�<�1e�2��A��K�I�zDB�/�Q�<AH�Wt�Q���3	��e��aJM�<	t�]���a�Q L��v`jI�<�!H��)��_`��
WA~�<	��ݪQ�&d�u�֝M���T��}�<Q!�2s���҈�//\HRÌ�w�<�#IVM�"��`�,���r�<�a	¥U1P�6�D�P�Hyr��q�<� x�re�H?��c $UD�Af"O.�2��N.����� `���V"OVtzVH�]�y[�E�,n�\DH7"O`��4�Q�0����+��"O����   ��     %  ;#  �-  8  NC  	O  4V  Z]  "e   l  w  ��  �  /�  w�  ��  �  U�  ��  ڳ  �  `�  ��  ��  '�  i�  ��  ��  1�  q�  ��  ��  � 8 � �   f& �- N5 �; �A H VO �U �[ oe we  `� u�	����Zv)A�'ld\�0�Dz+:�D�/g�2T@���	#Ĵ�'��?YV����y�抋<+`�2e��M�\��T��IYn��qA��nmztJ�H�(�� ԇ��_��x�l�)R+?��	�5�ص��"ӧ=�d)&,� rxD!�Xo���0|&� FC�`��;O�H�8�'2���ծhJ��V�I=@a�$�
V�.�l��5㕊�)��ɞ�`U<��`�#̴��$�O8���O��O����$؂z^�A3�I*��:��O���Y�۴���O`@����p��O
���#��W;��T�H�)jv��O:�D�O��D�O���Ox�1���(�Z��َw��堔�Ӎ@�+�/��H����_c>����)��p���JBE
��W-]�S�
�>c�����b�>��'X�O���j��U�`��y��Cb�6zm���E�I.a�D�B��O���OD�d�Oh���O>�D�|��w:l8��� tH��F��l�q��_r��a��l�?�MC�n:��näiA�6헁��!�S�Bm>Lqh$l\�/a�0R1�[%��u�'���'�b�˶�:0f
�0)��WǺl��'� �C�B�Q��1�H�Q�4�{��C-1F2��0��S]1��#�M�3�i����t>Y��κ�%�$�4��[�U�)�߸�Mӄd��>�@�6b�d2�[�cӒ4���nyD6mW٦�4Aɼ ��B�0ȇ��8f���l�-�"D�1�T�@ɛ��c� o�,H("�)@dl���)d��(k')tK�m�Fi�"�~��Ev~b�KG�ٌk�����4f"��}�P�{%l�58~f�#�ψ7��sZcH`���A�h��D{UiC�5��%0��i�r]C�-nW*c����K��'�O�ʡ�M$"��C@�*\�0��BI�`׺DR���O@�Dæq�S�?i��)����`� �����YG2�])���6��"v�ٰ!�2R�����D�I�G2�h�-��B�ݴ\Wv�q�D�:t���NR�l������0<��f����Tሏ�M&/I�:Y`U�s�߽^n�F��5΢��Óy��ѕ'n�W� S1�Wt�$D"PK��l����\��}������ryB�'��*gʝ5֍���` $Pʇ�'C2��t���a�|���y�O7�=/>* �&�
����b4쁕B�S���C��7�M�����O��Q�oK���#�ͻ9����W	g��'|Z�O�x��E�$�|ӄ���A �ӊT�hi�$M�)�*�P6�v`�l�'N���kȡ2�t���h��!�/��OR��`��R�*��1:R��2���O8�c��'��7��x�OY�I��@m։{���-?l�@�k��r"�'02�'-"V�t�|�/�#@���3�l�T̂�I�'"bhs�P�nZԟL��4���a�8R�,����59���6�>	���'剥oa������'��-^@t��釁,>�5� /͚f������i~�M����q�h�^>]�3�	�(r��3
�ƌJ���]v��p�� ��բPl�2Z�͓U�Q��O;Y�fU����ߠ@��!I�������)O�IB�'����?�OL���+kA���Ҫ�Ov�"BC:ړ�0<ɣ���y�p1�

�_���&����ɨ�Ms�i�ɧ���O�8}�R!A0�ʚy���o��t�%J-���d�O��<1+���^�hг�oǑ�rq{��?|j�H���P$1�6P�"����D�!O�-����-z�n5��'ӻe� T�@���bq(���K�m�=#u�=3MRIcAO1�(O��FI��p��Z� � 4"�p���  2Jh�ЉGz"_���'^r��O�~�&$"���b�(�����<�y��	�x| GЊh��n@��?�"�i��x��oZP�$n�(;�7��O���Z^�����#4 
��E�ߩ\5T��O4�8� �O��d�O������E��F��1hY�1h^c:ტ��2R�R��-� �6�3Ó{�R�dlK�]0,�`�.�1��H&ǈA��(r�Ă=1kؕ"p���x7o�*-"�X�@ �p~�Nޞ�?������'+J�����/E�%�LܱR��
�Q�(�Ix���������L3426M�t��((�`i���'�6�-)�~)#�U��6��S�7b���n�Ny�$� ��7��O��Ŀ|�',�?A�J�[�A�Վ�)B`�d�G��?��T�fLc� E�v6U{�
J�k��A��H�1x	H��-��y�ӯS�9Ԁٛ��̨��A9?��hd�����Q+Y�9K�!+I3PLP޴	�S#��ؚ��� `U��v� :.Z�Aª��I>�Ms����
�R0qU�[��!1�r��'g�|R�	�>@�8A���>2�dH��7���?��i��7&��Ą9%�Ѐ�L�*�>(�$��x]&HlݟH�I͟���D
OP���ɟ��	؟4�;|ud��d����A(����]P�bA^(���I�Al4�Ѐ�u���P��h�jT���H@����в
N���#+�%q3Z4��,TD8c���<��ʧyĶ�w��ۼ�g�RHX$�D�(:�� ��f�)�M�$H�>����՟�|��ş���$�"!9D�§ �t��f�P��d$����]���WBƸO��� Ι�v3vL*!o�<ɂ�i�z7��OF�oZ͟���?��O����FN�,����,Q�M:2\��S�B�&7m�O��D�Ot�S�'UΌ�{�L_�4��{U��237Fղ"nʠ8�,%30��e�`�zE;,O��ەfF1wB��5�̷eH�ҕ�O�:l��rF�X2y����@�qX�`-=u�Żʂ���C7�F3qF���'���'��OP#|J��Ǉ/W�j�拨Ė�!g&�t�<���/7"i��Dڗ
�$+�Gn�	(�MC����5�`�oZ���	=(�48©�Ht$�9Ŭ�(*>���ǟȱE��۟��՟<�PoX[F�l�
X�	E�Y��� �!���m��`���;�*u�c�'����*�'I���tM�+:��nׂL�.ac�GI*us^ +d&�������7J���D ܦՋ+Od${�BH;�����P�zJ0�|b�'�m����Q�:D"��_��${����>1��i9D=� .�?_n��f�ʹw�*�*��u���%Ϭ�E�i�^���y.�.l�4��jF�(�4��P���%Fb�'��p Q�߆�Ʃ �B5V�������'^�X}h��D�_|�u�'A�P�!�
lJ�
 q2هlR�<�A��,�4� ��OGƌ	S�l_81Sֈ"����O�|bv�'��7�\�Ok�,��y���J�:�րڥ R�Ng�}R���`��r���K0�֕�1�8��?a�i�T7-2�Č�9����	>��<�E��\���D�O��p�������?���?�/O����i�.ְHf-��\ ���$]��^5��e�X�pP����j�'��=�G-ǹmn�'���Q�ZEjCT�M�2 ����L�h��M�e��|���/�q͓J쨢u��a���@1��X#��2�4��I�����f�g�*87�P�AJ� Z�D1JTÐ9*�
@�'����uش�0|R���3�"��C:>�`yk�ٟ ���M�4�i�B�wӄ�'�J*�zt� 
2"�Z��4JU�a�$T��C�a������Op�d�O���L����?���u=V�
��R�d�ruV�P���bBM�D18����V���j�2�p<q�Ȇ�$}D��e�_fN��J��gL�$�pƖ;a�$!�6�%JϢ���F�4�-Fx�&�C5�����5r�n�c�`�$��<(�V�(���'uTb
�A�� �D�E�����'���'Fў �<9�'�5PL�ٛ�L��>��9��_�I�M;�i��,��=8�4�?��~�����3��X�&܎�B ����?��@�6�?�������2-e��� X!ך��Ei�1iH
�]�M�����G4��+�?��ȃ7(S#w.�v""J̅QWN�~#h��VB -r��6��Q���'"����7呜��[��	�&�M�a(�$)�O����W�A[�	3c+8J��s��'2H��]�n���	��N
��ף��?�B[��1%J��MC��?9.��[#�O��`1A֋��,��j��hך���O��d�6]ڄ��uo�3qפu2㓓 ���'��)	P��%B%f[6P����>:~��"[P�{Sϔ&m2A�ݯs�ĸZ�7:�X�'T8l�0U���x�
��N.�RM�'�6��˟D�D9O����T����_�n�Nu�"O@yY�֊`���X���z��@�ԟ{��G\��xd�A�+cx�B��M�0lZ��p�'�(��s��>���?�-O��uƠu*��^�Y���.�إ $�>~��q�F�Ѡ0�˧��=A�o���쌫DŘ�'?ꭓV�Ѽ4�l���ώ�y1����#�aw��|ZЄ�[�M�-,��vfڅ0��0F]�:y�ڴe��	0�������g�{�`٫r��r�I���,��\Fb�+�'+
�=�����¨9���&xt��Iҟt�ߴu����|�Ok��Z��a��W;�$q0��V�]:ꠓ�H��U'��27�ß@�I���ɺ�u��' R<��!�$��=k����fO^�F��S��
F+f`�����L�<�j�Ԫ�p<sO�).��R%Ž ��B��ĲC�Hź�u���fJ�Dq����ЦI���E�<j����M��밝x1d�Ov��-ړ�O��p�BK�0	��P6OD�H� xh"O�Ȋ�+��v�Kp�[��X�|�-d���<�&�֖f �F�'�I�<����]��d0��?z��'L�u�'��'�"���A z�d rg
$ WVp���By�!XE��ƮQ��Ok���'��H�([s���V�^�<xND�Ek��W7l 	��7b@zhb���Ɣ��Fe��O�D�!�'��<����T���vq���T���0��ğ��?ͧӘ'�
�#QM��S�|�QE���g��/O˓�hO�)]���9#��?:Ƅ�ЏT��5[A(�7�M3��S�6�;h�P6��O���O��)�z��D%̈́�S���z�������æ�d�O<U��닚NB�'��Y>�O��s�A�y����(�0 �T`Iu���D�R`��q�>E�dD�3I�l٥�D*j�<uŕ����T�ҥl�|�o�柬&?���!,I��J�$E�/c^�#�G���t�I���	ꟼ�	ϟ��'���'9�)^�cl���	,q���1FKpў���$���<q�9�኶�;B�iڶnX�MT�����i��V�܊�K��?u�Iڟ���iyM�_�,�#ƥJ3*�� PQ=�x]�wh"X5f�n��1X4-S��?�3�Imn���œ0��Xa�]'U8}�wb9J*�q�`+�	�
q�2�$�ţRg~�������Rs���B�^+s��X��O�O��U������d�	^�;�����:8��#b��01���q�<��bƵjY�yh2e�L;UB!��D�I8�HO��O˓-9ģ5nY7}7�=���� ��Jw��" }HA����?i���?!���?���t`��f��!;ac] Eb�J�*F6�
I(G�:$P�Q	�zӐ!��	)a�B� \���S�X�:���mtPr�ս�p��V�u�Iq�a��N �E
q�uʄ	�{~bLR =���e���8�.�鳉�/;}V����?)��d(�0#@�b7n�yyR|���S�T��ȓ5�臋�^��1`r�CX�`�&�̛�4�?	-O4�1���y�	��(�6��@yr�	2��;����Eʏ؟��ɶ�����؟�'c������	�����M�TgD:Lf|��L1fE�Pa����$;6\b�<Y1�nm� 8��L�ia*dB۴B�h����|��[�y9���7rd4��&�Q��qB�N~��P�?��|�ɘ�%GB}���S>e��A
��yB�A?�~���(]_�2���D ��?��'f��U�7Al���孉gKL>��d���|�[>��.)��rWh�>%ƌҁ��pD4����(ZD�3��m����M]�!�ZV��h0�5����6���z$��&����`�U��*��6-W�\�Q>���@
 "ڂ��/n4:���J)?�Jy"'2��<��OC��EK�$x|8�.��	���)O��d�O^��?���?��_�Xm��S�"hk�'P H'�yK�� ���7��̓�?ѥ_���',���zd�=���\�jq����6&�6��O��D�OLXIF!�@���d�OB���O:�ݩi�f�kq#Ŵ;��:A$��Q��'(҈�i�U�a�4��Td�/<�8)B��V�h�m;�'#}���(r����y��^�x62�s�
��<&�b���*�fGs���$	7�|�$���i�O����O��DW�Pf�3Q&�E�,�{�����U��?�(O�d�O����#4�a{��$�.ൃ��ퟘ��'����<9��
�����.=�&MZ�.J E.���u�8����LB��D�O
���OM�2�ҾY%$1ҕ�[����*�(����Ș���8ni"QQ����8�֥rӴ]����ӎm��-O��H�TE[)P���#��%��5��,��IUf�2�LdӘ�l'�M���C�
`4?��ٴ5��e�%�������$ �L�X��I��M;��	{�'���`)�������,,�T��'�PP�B*M7x����'�!�<�bH>!вiC�U��s�F��MK��?�0(5N0APd�֝Abp��ř$�?��r��A��?a�O	��"'�r���C�>1�6 �
��h���b{ ��S�O��t����(O^�x��ܖr3�%aA�]/y�
6m\�r����\�@� q"	U&R�6Y[4��gT�A�P�Ώ���E˨��	?��v\8�Ԣ 0rt��. 
�=�ȓa����"�/���؄#U� ����	!�?�q���Hq��Dִ�D%�a�X�� R�Eݴ��O-|�q��'=
��r���hL,-�Bm%G&�x��'��%)���s��/V4�J!n˺R5�J�>���,#Y�|�D�����c��4 ��a^ܥ�G��5I��6�ōX� EZ�EP.I0u���b)jИ�ո=ݪͲ2f�1:,�ܑ�F]~�̀�?���|��I�#H1y"ES�T�T,��-�!��Ǻ3В�B�%Z.�l�e�*zџ0���i�*v���� @�*pܘU@� !z�6��Or���O�d�t��m�n��O��$�O��])T�zXS�m9i}�TiD��kCa�0Dא�2��Q!^�V4E�����y�MT#]��l��+M$��a��[�,�-{������@2�U�R$d�����y"a �(\��2�e�NaΝ�T��?9�O̐���?���$
�r����¸8m�D�Q-�C�xPYA Ԕ-7Ԉ��S!}��˓/�����ڟ4�'J�P��ډ�����I�z� �b6`^.*��\Ѡ�'^b�'�~����ԟ\ΧX�v(!`G�L]��� Ў��q�� h��F#Dh�]m	=�џ����2o�P�qƁ�a�� J�$�ڑ���p�<j(n�����:u]T����|��]�'�$@Dǁ]
��3�	�n�ʉ+C�A��?٧�i&X7-:����Oa��a!U���iȩvzBq�
���'˰8�6������ȵ�;{!r)�I>1*O��fր�R_��I<>;j����2Xp�Q�m���	ȟx�IX͟T���|�P�=F��mis!�[�D8�P��1�n�qjǢ!�p�GHӜ����dO���ꄜ+{����F��mV���	���!�.Ğg�X����4'�0m�s�7�|���Ot�?�R%Z���QN�) KP�K�,%�4��	��A�R�R"�QiSf�5dx��D{�O����C{��I��R9�U�EA�R���Ʀ�M���ȌbgF�O�݉�H�n����*sb�'����d���!Zņ
~fp}�q� ƹ�J?Y��Q��葳�i��cg��*�"?	��ސC��@�VL^�X3z5j�ES�EX8UI�'d���UCֺ��C*x���S*R�0G���+?Y���$��4h�>Mͧ���')׃;2
�q`%��rz�,��+�*��[Q I��ş�A���	��h�*�B�J  A^U;W.�$����Ƃr�J���O����n�,����O
���O�Df��&g���ZW5`f��;��!����F�7m�,@�T���D�']�r䡗�g�ج[K��
�H�J�j	M��pm�z'��
rD>�S�CB�M�Q�r�� 2�J���*�DX�˝�Gm@P��@a� ̖'�Z=Z��̟�'�1ڠK�=}5�4�5
�_( )�"O�DrF�P����SB딸rk6��'���!��|���򄔷NmM��fo� qr�L ;�1�gY�`<���Ov�D�O.M�;�?��������w[d�ċ�#�Tl"f�ڐ6Z�ɶ��}��e2�i>bxA�e�V2��Eyr�A]��ȃ�:�\h0H��XDׅ�ؕ��n�����F�MK46hDy2���*V�h��)��aV�^���
�j��&E1ғ�O�$�A0H�4d�ƃZ�:�(�r�"O�!�f�6�<��kņ���a�|B�z�\�D�<'V7*��S��p�s�Q+	j4�a�ŉ*ɒ�S.����I$%D�����'0f��+�G@��X�@(�*
U	��eҌZ|�)!�� R%D=kE����OʱQ�@	�:m�x�jDM�d���R�$5203��0x�T!8B��2Y?��?��̘ݟ��u~¦�?TPB�Ϋc��A����0>��JF7���!BN-��lS�!VJ��X{�5��z��ȼ_ �̐`�]�NUJ�	gy�&]�z7��Ox��|�ҩ
�?A��_	$a���!H�9F���?��R<�`Ys����9[l��#��<�2.���طL8m�� MC��d�� h#?	��W�\fI�ǝ�F(�%��Uqv�i�W�mn��!�il�QydC�5n�D�[�ǧi�ܝ�'�ȉ����v�<ҧ��b��b^̰��g�=m����t��6�y�N@J$ɀ���;u��y$�ҫ��O��F��K�:h�DO�D|��Ñ��z�6m�O��D�O���w�� b��D�O8�d�O0�I��� {���Sл��;()Y�υ)w� 1��4Rx0ei���~�g�D�D���k�+fX����S�C�xr����Ƭ�b���((I��O4~��uQ��|Qd�M��w�P�GQ
�����	7�Rm������(I��'dў��kT���(!6�S�M� i��H{�<!G��H䘸�ҹ7CzD!
Kyy�;��|2����Z�m��ԑ a�	(R 1 ���Vt��S��1��D�O�D�O��I�O���|>��oA�S?�(S
 � �t��%X^�rhJ�a��"��(a`A7��<Qfj��<ѫu�RB��B���!N��a�׮S�x��tN�%D�H�1W%�M�4�V6����O���ū�ZIv鉶횗@ji�"�B!l|��'�ў�Gx�m��`�l`c�
{���U�Ӡ�yb/����Y�b�1 ݊A�͚���_"�&�'N剼#�����*��F<o_�S��Qa;��SpJ2,~.���OP��ec�O���n>]*�(ؒnZPR�'ĩ~��b%Ch�B H��t+N5NĘ6+�R�'X�$	���$��1�E֬xDqr��$D-p�p'cJ�Z�.��ψZ���C����O�8cZv�v�'��	��it�W�^1LI��吣��O@���� ,�j�1�*��u�|Hig�6R<�O��=ͧa8�cՒ+7�y����7*R��KVBJ��?q*O@I�%��O����O�ʧvHFp#��#���SfU+1zt�YwB�^ې�B���?���
AH�����$kf��A"��o���#)�؜��C'#l��;�a�"���ɝt/І�� cw��p$��E5�`�gCD���L�1J`͚�J2+�g�=Ú�����D��0OB�Qc�{�|={+̵5�&6l"D�@�s��=`��h�oӏ""��G�?��?A���=<�� V�F�����g�����	����'�ر��'�'^�`�J�>o8ᛃA��3��0z���-�ԛ��$t�8���E9�Na�O���$�z�����F��<=`A��|E����M�� Ʀd��,�ġ����d� ޠ:$εC�,��L�,�D ��O<�;�oC�T0�Q�B��E�d�<Mu�ջ�'�R��i1M�'�܀�~�1/O� FzʟXʓЍr�f�<�lI��-b��T)'�Y=�?I���?!���?�	9)��p���zF��F���0���c�K�`#. ���M�^u���¥&O"1���:�e�F�%ep�X2��\��$���P�Le�S���>�p<!��
�.��9�J0eb��MS�Ox*��	՟�D{b�I�z�> ��[ J� b���c�`C�I�t�2��U�:Z�R�d���:�O���'�剴|S�i�K~r��D�1��X���D�7����Ȝ���'�R�'��nF=
�2U; /�1gD8�3wo4!��Xj��L�p�/	z=>��a�'t~�{���K/����G�%�RgP�ek��@���j�4�1���0<a�/�۟���@~�o�L&�]
r.�;k:�=y�������0>I��%�H��s�1u�����jCF�����HPL�3��׊{$8(�Fl�';�~��I}y"�L��)Z*�����/H���$�ʓ ����P������O�|p���������k�;H�T�g�(�Sc,��RB���Syڍy6I��v:a�'�,dR ���X�4˅�I2`/�F�dAT�:b\Bg�$#e��W/KP��Ia�'��>��S�? �``-߾r�i��D�V�z52"OZaph��Y�lłV�� ml���h��q0Q�X�B����� Q�a ��ˣ�rӴ�Ц��<!Ƨ������>z�ȣ¬3>~���EOYG;�u�&D�"���Bp�Y��Ȣ�o�m�g��(��tc[�;���I�!���cJ#pC|=�P�ѫblN�3e�s�g�T�j����*E��ɺa��p�u�ݴ��	�B`����Z�g�I�H`^�U�O��r 	�S������xJb,:�`ʻQ��� �厰��̖'�"=�O�剠;�A��K͸ɞ���S���B؇�M� �l��P@��L1�@ �*�;�~�qΜ;{ ����r�H\B��ɚ ��x�F'-$x"�_c��m�`B�i�1�@��%[����0O�e��ɐ1�� @��P����J��%��=��Om��HO�"<!�+˚o6���iZ��ǉW�<! S�k.]���B�P�U:&�S���$�<iAmƋ���G���(f'�����2m4Ms��J:�hOv�	��4"|��`ҁo�B���r������E�`Z��<*9���k�7AԬ���-�1��I�]�"�D @��7)bV��E�0C����8Pj�C�ɋ5:XP��ܽ7���xO-\������(�@IO?`���!�BQ��|��k9���%4�bo�z�֢~�&b�}��%R�X"o_R��q~�d@�x�Z$�vAǤP��X�"I�d�O
���&!�h��,#Ģ�P�A��O��ůȏ1�"��PK�%��T*��)�J�`)U#ryP}�vI #���+G���CĦ�Њ��v>}hR�=:�HI5�Q�*$� +TJ3D�8�v̅�b�F�3���u0�S�?��he�>�H"�K��uc�GJ�)Ϝ˦����dy	����3ʓY"~�kS\��i"[Y���d*!yaz¢^#=���ó� �u@�\��&ؘ'r�3ӓ_A0@9�I�CG�髥��*{z��`M>���G럸�|�<�#V5MlI���>z��� ��c�<��E��uu6�s�9F�������xy!*�S�OЀUh�N_8�j[3΂�=��P��]�'�8(T��O�Mp��e��a�8���w�I�Wȍ7E�D�#�-���p|'�'��:��'�b�'r�k��M�S҈HK�����mz>5)�M_G�,12��0)�ja
G
)�J\M�NY�f<Yk5�ٱu��`q%�>��4�'F�&W*���&����N�B
��Ё#�s~2���?q����O��=�P5�X�Z�l�
EV�)O���$߫/t=K3E�oYxq��A�'��s�x �%�:F|��#�/⺴�'��-�p�'�Bu��'.�ӮMHH��������"rF�[��|�ZEfO���l��b*R���W���3f���)�|2�O�|1�G�@�2�����85��Q��'`��@��Α<�ιZ�MQ���剏@������!%�ᱝO�
����B�`)J�%����'����?��O�OM�	�~��0��Jvt���bR�g��C�Ɍ_TV���uAv��z	£�$ړm̑?�Р��c`9{`��']��PzQ��ru�@����XR$.!�&��S��џp��˟�z�L�::�3��ϔ
d��Dў`J���3�i��,�a��$A����'�����M"�Vl6#��9q��C��\d �3�˖YGp����@	|~�؉T"�95��)K���煃z��ʈ �F�iB��r��i"捛W��ɢ �6��O��=џ':��#i��8H1#��R4���'��{AeάX�xh@�B4#�X���h�����ĕ'l����D�\�.��Ɓ���j0I��۔M����E�'0��'���O��'����w��ʴ��̘���!h��-
��Tf��3�1KL��eI3��%�= �@�zޖ�Q2�Z:"��3`y����PB�%+ K!�@14ǁW�'��8������"��ph�P�D�+&��!���hO�">��h�R.fE(f�H=R��t�"dx�\Dx2�S S����k"�{��(���Ц]��My��$��&��o>%�ƪ��#��)�6��-7f��e��O�]��k�On���Ond��,�*����Z�f� ��?�2kR�i~���̏��,ʰ@2�x-�����h�
}�sd�ek���&�ڤ<1��D,1+�Ё��N<يUh@D�d�'
����?���D��X��G�Kin`;* �_-��0?y��R�cA 
nq9�+�{�K���4
�<)��I/�,0j��B�}{HD�7d�gy�l�=�'��U>��� ПX�I�EL:P(��1L{����zU�i�	�j����W����Y�D�>e>ହ��b>ѓ���춥��Í{��L�w�|��I�I�!I��D���C�O��BNV��uJ4N/�S>^�&}�
�Q�`���N؋"�|�	!P��D�O��S�q~
� �D*g�ZD����3L�lcC"O2�'���:@��c֡Л �ZE�����O��Ez�O��I#�,H	;��H�Q��6Ҵ�!W�'�"�'��b���t�'���'��D�'�!�gl���K��;W1����H\
�dx����~0r�Eƥ;���e��T�Fx���x���h��U�8��l9Vj�w�B}�ɉ{v�����N�
�
)�8�O�h��	�#�q�#N�Ґ�W��P����O>�$*ړ�y�k��Z���#$Ӂ:X� DhN$��x��E3����҇F�7|�����	QB� ��|������&,�!
��B|�����+��8�&V9HǠ���O����O*�)�O���e>y�ҁ߹G�^�趤V�gV �2K]7'bt�w��~�=re?:�
�E�(�(r7&��E�B9h(�ಉN/�N��Ӈʱt�j��e�P>�@���T�=	B�b��ā�Z�2ȇ�c�8h�	��vID�Q�@�Ysr�IT�'��L�`,�cJ���&C=,!P�ϓ�Ob�{u�'��T(\6v��[��UyҍpӰ���<I��ǔa��&�'��1����Dn�*spkć<�$��'X�\�q�'�B�'I��㏽/k��r�M���6�(C�Xt�7���E�@)��J5�$u��i�K}Q���A�|�Э��D�)��o��M��(Xb�}���� &P�/�P`�>!O���DiҴ5ڝ�'E���gɧ�$fKc|�b�� ���;K�ze��'��E0�� 7�|��#M�H���k�7�I�)��J�*���v팧8ʓ�?�����D�O��'���Z$���O�h�x�ڦ"9O�џD(ش����(�	��:�J_5[t8���Dc�O��{M|BbW�2����,�$S~N郡��E}�&�',���P:O P�B�'_��O��'�O�����	
��!s���)A�M-�6��On�C`g�O`T���5��s��NO,�yr7���P�@�>C�<����Q�^�?��?��T��'_���Ox�$�:��k�p"�Ij����� ={x�cኪ%qf�d�O&`�#f�O����i�b�s��N
�yBǙB�xDP�lՄ.OR�#�^�c��lG�?Q��7��fY?��ٟ���J��!(jL��e��I�x�q ˙��?�"�Tş��I�~p�	��?���Uxnڴ?&��r�(o�|1� #;��@�����M;��'+D����?)Ӧ	�Q��S�����?��F��;�2�
��&aъ�{wƘ�2���f���I��$)[w�b;O�u+ߟ���[MT��a������c$�
 �-!��1O��҃x�R<mZX�}��u��O���%�"��+̹`����������7m֤�z�����mڥ�M#�'�?�d�'w��ؕ�O����"�B���*2g�`Z���3�iKNmP�"}ӂ��'T���|�J���]y�'.� l�Th�G?ܜ�Q���2�}� "O��vዼe��\۔%�=j�l��Ľi��'�2�'���'���'�B�'�.X�d"����xԈ�8�de2��yӪ���O
�d�O�d�O2���O>�$�O���g�f� ��E�I�W>�,�Bڦ�I��Iޟ��	˟D�	˟P�Iß9�<�c %���0#eL��t�J(mߟ���Ɵ$�	ɟ��'Q�SA?��^�c��MqpG�+�<hp�b�Ӧ]�I䟄��ʟ�E{��'��,c@�,F�	Q`nA 5��'x�IğԨ��B��n�D��]_td�� V���	�a*c��l�Φ%h��?1���?�����|ʑ�9Im�h�uK�&��9I֎d!�$�8��}�E�5�$����*!�Ͱ��ɂ��3S�ȱ� �ek!�$E�i6�0�E�$���& hf!�d	iD� K��N��jX�i^!�$Y6<�`��m����Di�t!�����şd�������<�p��n�!G���*Z�D$�)ٴ�?���?y��?���?���?���2��kU�K��Q����@��w�i���'��'�B�'�2�'�2�'Ъi��C.	�)� ��	g� M�Fp�\�d�O���O����Ot��O����Odu(%!��=|��#΁G��򧤑�������џD������ܟ,��ڟ�PӮ~*���P�͡$��a �ː�M����?a��?I��?Q���?Y���?����m��+Õ_�d-�c .B���'�b�'r�'XB�'���'H��z�Zy;���9j*)�&�� s�n6�O��D�OP���O����OR�$�O*��D+DFA�@o�>�-D��:aʦ��ß��	ȟ���ߟ�I���Iߟ\��='�r��ʈ�=jF��`�ɔ�M����?���?���?���?���?���4�ҀA���.ar��$@֦s���'���'�2�'�2�'���'�rc��O�0P:4�Ŕe%�D�k�^�6�O����O��i���'���'M��'�0�ĕ� �ġ�O�42��I`����O��D�O����O6���OR�$�OP�*
�HJ�f"ڊC�S�i^�����?Q���hO�'o���
���`t�RA�	�t��j�4S�܉�'���O�����z�4�yw��
7$|�� �
Rv����:Fb�ii�<%?�b�VE���I5�MP�@ώ���`���TV`���m^�XP�]�x㟠�i>�̓C_�mp�&�7=�tۂǋ1y�2DҥcӦk��<��D�? ��g��{r@�ɅKt $+��'��I��`�-O��g���	myrϊ�5]�Adɇ�$�֕0�۟��d�%w�RY�$៲wH�i>���H?gܐ��s�*�҄�u]r��D.��)9��F{��'�ڴy��ܿ3�z`�$�>Q�<���0��fD*�y��'��6-�O���|���4��9��� Wߢ���^�_"L�'��i��	�D��!��O�m1aM�	P��%�Yw�~xsNȤS���_�D�K���'���;m��&������͹o�VH�1�cy��d�֑yD����I�?��O���^r�aq�4����-��ʓ�?�4�y� m����FiE�(�l�1V/L.+��
nN�n�8�Q6�3w䜉�(q����?���?���n�n�٢LWJ;���F��C3�����?9��?	��?�(O�]o�E�h��+J�QrѭM�`O�q�H�Z�x�	��	��'��MP��O�����M# �XJ���kĻJ"x��Jز��X��P�<�޴>�B٣1c�.o<���P��i�'�~�� kĂ|U���GBc���q�M��y2 �?�8�S��K5���6(�0�0?ɇX����IM�l0�q��Z;3�1�"��S��t�ǡRE��Q�<7661ZJJ�p�����_/�����L��-L�!~,A�D�ʙQ�5'�)v���{#E?VP�LiІ^�kF�IF.K�=F\�����	<i�զS?X�V���AR���.��',\>m��b�x	A�C���ҟ0����"���ݻ�	�K78-
�J�1rdb���-ʽ�?9,O��ěv��B��� ���j0)�I�!e��؀��Yݟ[޴j���ƗB�ؐ��|�O��'�V�J��:�V�A�љ1f�Q��E��y"�+	�]��1�,G��Dx�Ĉ��8���D֐U�r	�c)ځQ"��!	P�B��Ua`��-LK�	���At��!A^°�bt��5�b!��!$�5���7x#p���}Zq��S$�2M���";!��(�D�d��d�֏V,P|ӣY�,�`���'@;h��5釥K:
Eh=a���(��P�iޘ������C"�{$f��A�S������L&�������{���˟d �I�C+�t�'�&VM�Y1!���(�I��D�Iܟ|����pㄜ�M���?If(�B*J��`�R(Ee6��K���?)����?!���V�{���?���c:8eO08�ћ#�A1
�u����?��?���^�!x!�)쟮=��� �I;�����	XJ�E��<���O��d�,#>��O,�D:
KҦ�K��j��(ksÚȟ�����hba� �Mc+������'O����.R�k�D��,��*U���?��PE1��?����O���)�җ �I����x��؀��85���Y @�a��
�g������v��Jm�Pbɼ�GX�qI��R�ܽ[����E��(�	0�IA�ϟ���ǟx�I�my8��A����+��2����H�	ԟL�	ڟ���y�Ɋq��])1[�a�����%�Cd�5��զi�I�?����?!�����?Y�G9km��k"�	5�m�Ѝ�}�a&�O۠�΢������kv��vOX���I������:/ �p�3Ά�t����q�ߊ:{$���"�ȨfK�æ�r�438��˲̃�`�l�8�Gܚ_g�e6熚8��e�U��Yj����Z#jg6��Y+EAxYzdEِKO��·䁔$ȨɊd�U�M�8�T��8��17n�h�d��%̝�f�jd�c�'���'��#�~����$*�(.�J��N�e:!b�j�����Z�`�=.�L����L;z�C�IY.I�y���?J�x����?�pu��I�f��j0�Aa��Cd�t�Z�Ɓ7^���lZ��M����d�Oz����N�́��.]��	@�D!򤘅Ut�M�u��1���2��.
�}�h��pyb$ܦq�;�?����MS'E�8��S����H�QV	M?%`�k��r�'�G�袳�P�I�©A$���t�;�,ԥ[Zd��z�'��AٴT��m�a O�u�6��L ���T	X,@x�ia��-% ���QG�5�O�@�v�'�r����'uv�����'�&<�!+�+\����O*⟢}ZV W�K��e���(&H���E�Cܓ�hO�)Ts?Q3K
v��1��%u0\Q��?5��I	QXh���4�?�����	S�3.r��w�0��!4rt}�i����Q2r�۟ �%�Ο��<���Rňl��F�7F"�ê�N�zD�'�`�����N
�\򒎃?1�u:C�%>��u���	۟ �*���MIO��|
�賏�	 K"��I� �	{؞x�Z7�H�v+�7Vu���$�(Q?q�W�Ժ.WT�V�,��Ź1�'�?����?ᖤĔR2�D����?���?I!���7�#fA��Y��w/PxH��P%sð�EBs���H�;g6,���5��d�)4D�@��:K����e<,��8��4"ȵ�҄E�ы��tcdӸ��Y��s4`N>�͹�%�(A�ٲ6H<6�	�5�����1����Iş�n�}�ja�`����M�� 8 B�	<3������}�� ��:Y����S^������|�'�`t:d�ؗr��LWC�5J۬)��J~�b�@��'{R�'���x��IܟTΧW q)��(o�q�*��c�Z�#%G�2F�5��CQ�ҁ��`�@a��1ʓ%F���%EϨp�eTƅ7*r6m��I�?�h0���LfĨ���]�B\ĲH�C"4�x��c~���M� 湂5��.�ڄ�$o�m����f��PxR��)��`��W�~M�ؠ��?�y�T0#b�}�W���s�B5X�,԰��I��MM>��\�s���'��iyxq�b��L<D�p��,tD��Ð��O@��#�O����Oxm���
A�}9`�>�;iWx��	[��d�8R��7	^~�F~R$�$~ؔqdl��Zb���C�<md�Z
��D�$#�/Cl�liA�������5������$�'���C��1������&1ò���p%lPb�枿Wp�`��T!(x��ɽ�~�&�oz�5۠��P�����ƭ��*1���۴�?����iKº����M��(O����f�L�4�QY1�6�(��\��8y0�"����	���˧�ħp��lZ���W�ʈ�E��޴�'h�CT�5zj�I���,J	�#~R�䙑-�1k�*�"i,	i�o�K}�Y#�?�s�|����h�UPT.7~j�@2N!�[�q	�M�K�9�mK�ɀQ�8��Io"ą�cƲ&~��Q��T��c��mZ̦��}⫟�_�lA�X�5kգa�T��#�#&|�'��IS8�� &ʺ'/Ƅ�`�{��i�L�wo�����8H����T�@+v�8\��	�	��B�	�b�<`[��PG�L�8��Ǌ�hC�II I�7�M!Xp� �°IXC�	>C@���*eT�p:DK�6�pB��
:����J \`�8�d� zNB䉙��=)���wB�(1��Ѭ@� B�IyBf�P��;y-r7f�8l(B��V������C����ΌDL�C�	�F��H8�腧����$*�k�C�5_�2%"�DXa�DZ��B�	*k��y��t(qҷ)D�\��B�ɔ;��c ����^��!�6=J�C��9�p=�P 
���Q��+>�C�ɡxS�����>>�!��C+�C�	�Z��s��L�D��%�@���C�I�h��i�
�am��Ӄi�#<ެC�y{�8rg@N�T�T���k��C�	�-�xPƉ"$�<D��ٳ i�B�I�5*�Ѱ��5"]p��b�]�fC�ɖxYhA'J�Ab\�
T���\C�	6%!��0��Yd|H8fh:<�nC�	8w�d�#&��o�Db�V�3�*C�I6A3�%1�Ǣ���"�I�_�B�I�t��&3d�������`�C�	(Xhhx!�P�:���aa��
�C�ɢ^I#�K�[2��+Ũ�4OC�'J�1r C�i ��ӥ�\�
C��uHj�� ǥ[�耓�"�C�I�?�,(aaCż q.q��dحW�,C䉷b�����.϶ �����&`�B䉭YvZ���:�>]��J�,4�JC�cd@#�%�2V��bHN�0�B䉗�:uS��C;V��Xs�<޺B䉑igz!�󈚈55�h�5C�cJ�B�1k��� Gc\;i����B�8!,�Ɠ$�@���Y5��
�("� x���L��@}~���E�*\�Q"Z�^��p�ȓR&t2��B�L��hؕ�I��(�<э��I����5�\�ѐPj��r�!�Ǧ
e�Ue�O8�}RU��p�!�ПsJ�y@�S��1�Ta��Z�!�d�8s
H� � [2;�����Q6�!�DW1R�)�A�'V��mx�!5\�!�V�f(��KR�-��`�GmW�T^!�DE>Z&~0Ƈ&�t�Bf��RA!�d�*@P����ǝ�m�"��`kE�!G!� �%�����@���j��!�� v�r̜�qX*�b.ڼl�b4+�"O���L�$d��"��D0Fɺ4"O�$ZVI�-:t�CR��A�޹��"O)��� s�p{!ݵq�y�"O����&V3I��]x��ǙF`�!�"O���M�gs1(0l��+�R�`$"O�)�)_"A[F%���,h3%r3"O�M�֊FB���W,��ՠ�"O, s� 
�zb���W)e��"O���FK�U=���h]�R��"OPt�c�
�cFB�Ke��T���F"O�qZ�G���q(�'ݼ5k<��"O<)���¾e�T� Tf��}Q*8	3"O�	(�R�t���#�&Q�@@E��"O��0E�	,�y�%ܣL��̪S"O:�k��g�f|;��؂%�49��"O&}�VL� }����J*K�x"O���$�4�8��fÙ6a*H�"Ot!S@D$@�������~�
p"O~HK�Õ�X�zT��Q E�b���"O>ͺEIۥ;MX�����6�`8�"O���0B�$刳J�,/�F��"O��p��6�T �@U�?�v�x�"O ����HHLJ�y��x�xT{�"O�, ��۬<#��S�@`̬P0�"O̥�Må9�,cA$ש^�t�"O��v�Ǫt��ٻdn؜�ʬ�A"ODyŠ/�R�Ɂ�	
�֬�"O��q���ZݸHŬ._�9�3"O�����!�6E���XԲ�(�"O� ��W�D�4BTS`|���"OZx�V���S�z���/3k0�k�"Oބ����,}J���1��x����"Oz���/L*(~|�e@�U�"O�LV!͟Z~�AG ĶB�ܥ���Iw8��+7�^�D�c����\c��.D��	�I��b	��R�v�8C�ɫ_I|Y�,�HD�æ��SbJ�����0<��{�(��u���ơ�� @6� �� ��0=� ���#�x�'�49
�f׈l9PW�s��r�'�D}�$��P"t`�aJ^p�y��ʛT~�=�|���C�7����M�W���2��W�<�N1gO��tiZ�jzp�0��ۨj�\�h`�5�g~��5���$�\�i�tYP�D�yrC=`qh�SѪO�~��h��۰*4��[�g�;����M.lO����\���-�#�*1�ĥ�$�'��9�S[�0�©�
�a�Z-�Gi#�|�i�n�0�����"O´ ��R7Ts�8��/�� ��M(ǞxK�BPI�]���P��*Y�'Us��br@޶9x�qca����dD��tEv��qH�"��D+���6\�� c�Ǫ�l8�q�̴
�e��
sܧ�ēE�JVh�,����B�U�N��A��E���*����9͘��!���/1�����Y�p| h��L�����R��.y���\�od\����sR�ː�ћ0}џ0�Q�S  p,}���[��f��vٻ ;�	 �2�tRa�;W,�#�KwˎT8W+�>�@)�i��:%�M��7/W�i�Q#^!>��,�0	5lB�[>��g"�^���0��f�O>aQ!L��(O�OSb5��A�/X宅�!�@�@����4D�A��4=��[�"��`���)u�@ <�Q�D��'����B\=tX갥V/az�8���J8l$�#}�􍑃hFIG�XO��毂�<��'斈�V唫-�FD l�6����'�XaYe��?I'� Y����f� �`��ybF��§2D�RPɍ����zp�_��y��0D�� ]X$������荪ܔ��b"OZ���	b���1Շ�4q�欘$"Of�ѥ"s`��PKÜ%�:��q"O������Vc��#,N�)�@u3�"O�t�
[���Ǫ�V���ʱ"O�`� �#��s$	\�x�v�P�"Op"q�L�obxch�q�V��"O��)�kA�:֠�I��g��<K"O&و������@�ěo�l���'�����D����,��g+s�0���8D�	E�ɶ?����%íO�|z��(}�)��+ {��T3/�H�Y&%�&<�hB䉫�(M�U�M�O�fM�b�ޒX��h�퉴n�
�z�A]�X�H+e'�S�4C�	�����������ؙ��:D��yc݉zk2�����6-���C1O�#=I�#	76X�A!��Ǎ;�@���AWX�<,�fژݫ���^�V�*U��Z�$����=��}2��"*Y�6
�;Nq�P0�d���xB�Ņ4�
���c���L���A8-PqO�����H:��[�y��+ȝv��˴�>��א:�t'���}�ٴJ��1���-(�F��O��:et��\|��b�߮'��i�R�W�#֨$��??���/#D�]Q�O瑞����NR��a��U/fp���A �O2 ��^�XK#A-�Z�
҃��X���+��ɴ6Ԓ��)�S;Z%S�Q&�
,cxأ>)��U�w7�Y�k��3%T��O]�(��� ����9�K�K� ���{��'눔�.��`M�%�5�6En�U�'s[�.دEf�	Js/���蟮Š��X�0S<����#u�Pi�"OJ|5N�8p4�*p�7Zr�i	���S琌oڦU�\��2(kD�g�'��iB�
�p8,�)�87��8!�G}��Ұ=����aB ���k�a�fu���*j��xr'����OڍB6+�u���2�c�	Bҡ3���;P�heB.�W�n�zQ��:���0q�h��,���yca�I=�4"O��i��#5�hq��s��"�8OT4z��A��UQw*��!���E���a�	@SM�5JSB!��@&�y����5� o��EN^�i����/A@�(AN|��A[��H�7�ʁ�A�?�@�B���LVDS��,途�Ge�	b�P܆�I1C-bE*B�����	�26 Sbٲ%�dp0��ٝ
�:�)����1PCH[���CX�~p�,F|����6z,y�K�?2u&�/�~��� 8�Rx1�V�I���� �]W�<� �Q�BI�E�{�v����X?�$�J�)����7KΩfj��F���5�Ұ�E�M"1����aH��y2��v��E�̫I%���
�5�ġq�9Oȴ���LhK?���A��2kL��RΆ�D(��P)�OH(d�ïu��8`��gc8��C/�:7�.�p�͢�^i���6x%���@(�Q��02QlT�:��?�FO�!�@q��q�)(~~�� B[��  C�ΑI�!�ɂ�h�i����H��Q;_�6��#�dIc�S��9Ő�0�M�_��y���6:����4J`�ϧb$Fu#�g��{�i��xl�u+W�A =LEi⣚�C�ʔ�����Հ;���vK�4x�$��_�����(U�$���`�,~�J��dA�T�e���t	҉�-IZ<����nT���Β��9a�7��!��a��
Z)(�^�J@���!��-�9���G�\�����=n1vX�>�g�2���b
�9 ��x�hL�Ef��`��F�<!��A�{C@��!^�3eH�5Gh�<!��U�n��Բ�)��te��bW�`�Jm���Ѕ��.V�<`t��/~����B74���R�"Ox�s4M&	~ Ű�!O��8r'"O�����^
�f,��x�|P�0"O� 0����Z2`���ָh���Q�"O<����>Jkl��g����vP w"O� �'���n��[�EV�q��B�"O*���2�l�yP��(�|<Z"O:���	����Q��Y�Rtp��v"O2�y����&X��� ^�Q��"O��'߱*�����!ћN��"O��D��l�K"����:X�"O^urS����T9�$�]�_�ht�#"O��z�`؋v�p$As&�-�Х�"O ���O�2��H(P%U�����"O&C�DJ)8�z���GN�o�D18"O.\ْ�_6)@�m#�܇U�0�I�"Ob���CJ^Ghm���'�>-HA"O6�k��K��4���j�H�"O��!4a=~�b��s�V�gZ4�"OXA��M�d\χ
%VY "O�DL�-tm)3�ܿZ��$��"O���&�Jg�@��f��)�����"O�A���>P>`��Ƀ}�T�:"O"�Q��K�o_��h�-�Z< 3��C�4�؁%Ҝ���[(@b�0$��2"���"gEܼq;!�d��'"�)2�����B0b��%"!�#��y桎�}��`�Sr!�û, 8����4&=����Xa�!��pH!Ǆ�;������B!��&O�h��BN�)#��`�DʷL�!�QB�.D�%�Bp0�K���!�ĉ J/��9�`ŞTS�1�GH�+7!�d��D�}���)c~쪓�a!�$ܓl�v��E�ڗM����gKA!�DS93c�Y�@�;w\��(�k!�䉔/��p@7BI:7_�!�����!����=�Ƨ bX���t��-�!򄌺[=-"��څF���ߟXС�$*`�<ݑVa
g�ʔ 2�y�H��n:(4�FjȊ^(��T��y�ٸs��)��Z3'��2���y��E�O����$����s���y�D6k�]!���5]�<���@�yR��NP���B-X�P蔴��Ե�y��5h@��1�S�<L����	�y���'5�Y�񪏧u�|k�(��yҤ۫$R�: ��1~�	1rmL-�y��H?1dBd�#�U(�!32��yb�
�$�������^*�򁄘�y�$���,IQ���N���B �y�-�� ?���	C�Oy`8�DĖ�yr�L��	2�\�5�8$�`S�yb�R{���Ca {Yv�Еa���y�E("�i�)�)b5ZI���R:�y��C�rI��e�O5|(�f㖶�yBA�6+70�v(Y6"P3�N>�y���_@��(b���N��٣�y���A�V}�%�ŧ.��P �,܌�y2E\3E��|�j
%��r'�W��O����k��&
0\�2��4\��ᖟ��Ț*S��W+�Z��0#1�7�R�~� �غj���S#�7�1�'G���E��+{8�(�!�&�)�u�Y�K�D鸶��b�"�d��r8��ؑ��$ $:�-D�Y��:�*iӲ4B�������4�͂�\$���	���#�@�2��pk�鍗7񞀂�
O$	镯/n�bI��V�J44�Q�F��y*��㉞M*���NU��[��V5������@]:�kzX���p,�4�8؈�)^�TP���d�A��g��'��́d�C�N�����E�I"	�J����C�w,j�NGRn��X�0�N R��%a�{��B��	w�b-ק� ��X�mʶh��VkòD���)����uY�m�B��0!56-I��^���Ok�'}���w��Y����F��j`}�=	��V�����ɏ@@� �bH�PgΡPTLH&0��
 ����Oh2�,ʸ3680'e�Н[���sJ����	�T���@sf򼛱 R������O�)
�x�Eox�I���D��:���Z!��z��l�H�Yz0��N�d������3su���4$�.B3<�b-}�%�M�8��4��(`����Z���'��lƷX�4 �D�ØZ̢���Z�����d��ȳ_7..�*wƚu�ZMB⨉�|��t�&��27`�[�����	`
�&�n��g�*%|��űi,B {�,����mQ��_�@08�����2b����2�P�l��dXG[��-!��$:ʓuF4��P�[�i<b�;�%�>T1| YcLþN5�xr��XzP��<�,�*bG��5��"�fν:TXQ��xB�OXP���b�DI[/��Q�'WR�Z�m\!0"�E;�,�[�1��bCq����F˘�DM�r�I���`����ȷE�"˷�R:8�X
*O�������4<��t�c�k�"ɳ�B'���̢=C�ݲ4�N�E���a�ԥ/ �-�7l�3�E[�G[�YVN\���d�0jJ ч*֗RuL�Fj̯U�R�o�c�P��V���qCH6mŃTh�(G~"h #d�Ӆ@շ,.����LO�n1D"�O\ӧ5
	@�`�8�k^�h���i"A�ZР�@&O���箙$9�h�YJ��6��n���P�hוI�HO��u�d�|b��ڄ+����VB\$Y=�}����J��d�	�-��O ���͂�2z%��3_n˖�>�"c�)�i�P�8�>�s�׋���ݟ|�I�W�d�Q$�m�J��͇2Nb�C�Ί#H��b�H����r5l� k�9� Ā�o��5�e�=��[�W(G����t��5�b�Q��S���Gn���N�s��}�(4�8�D��ğ�;�6l�ał.R�h���D4��~��:?��� �i7KY>3{n���
�>y�,P�ҿ63�xr��4z��D5�����8as�ӭ>q$]z�x��O$\x���d�O���	p��2r+O�HNi#J��`ٚ��!�$Kr��a�F�h����0N� GA�Y��bt���5����z�p%�$��ɟ�6#��n�t�V"P�6��V'�>9�K�
v�0r$g }՜i�3 �=ĩRe���Sŉ�z��?�J�MʈKa���۴��W<�ƨY91��ᓰK� ���������O����S�(m`��Xt�)����OL���F�����@'�LQ�DX�s���cЃ�-�p<�6M2!��Ȉ�wx���+��m\~�FD�%�p�I<�"o�~��� ���e>
��H���/Ar�*ўb��OT$�W��$<���m߂�:&�>9򂒐ET���b["jtl���"�E���֟�Rٴ0���� �T1i�7-�uW�>���*�hQ��G;1r�Ej�S=>ة�U�Y~�'H�L0�?��pH>i� Bɒx�T���+Cw�R���$�>���?�'d�UC���	��+bJ�*ɞ*D�IU(<��˒ � ��Ǯ�)R����^�}?, D�''H0b�C
:u�V3���8s�Y.h0� E5Qka}	�*"���fNQ���E��4$Iօ3"�p���|Pf�f���T�)Ȓ�	cL8}��W�d?n���HB�:�|�P��(�HOF�J�#G�_7X�R �@�0վl��W�\��G�
;���k]2�����Ƶy�Ѫ�K�>;�$1�\�*�xB@�/hY�1�0���jH�
C B�M�%F����K)�A�F��r�'i,5d# !0�ܭ�0��z܍���B��xe��T�e
�⎱=����%Q�?�v�H1ާyWA#Lq"�g��,��qfU2��$��e�@�8��|�unEJ�0�p��Sְ۰ �5T-�@�����ONZ�fӢ<VP����+����+um������2Q�@81���l��O@tP��Ej�#%ß���'E´`��w�8�j߄�}i�O�)s�ĞI���֪Xx?�M<��A�M��CD�P',��W%
�}!�aI2'��~�D�	q��
8բ��$30��s
��fP��VF�I�bP2˱>1��>�O��&����<�T!'M?-�5qSM@4!��;]�Y�t%пX.��pC�'�ڼ�	�u�䖐�(�?�';��u��v��9�"���L�.sÓS�Ʊ�b�7i�e��Ox@�U��/�҉��mB�� ���#}rS� ����E�0�� �h��g+�+&�l��'/ L VA�'���1�C��@�0�Z��j���Df7>��4	���W8�m�E�x�p�G�Z�Pެ�r���f؞,Abυ�l��\yW�A�^�f��S��2dv\�Ȋ�ԟ�]{S�$ҙi�Xa(gk5>|HB�jH I!�$¹)*�U�v#�~��(u��$�0�Z����i�J9B��4�(�ct��
]n���U�z�u+BGǷ%��
�e&����
�+��D��	�R���/���'t���AE��1���"ʖc��dIF����EM�F��0����FJ剀�*@�6f@�*T~]�
�Y��	jt��-��F��*�(���� H�b�
MB@���F@欀��i,`!Q�AR(T|A�� ؼU����D�i�h���I�)�̑�`�Y�T0�
�'P�1�q��z����I�=N��Sm3Z�.���I��9ӲF}�P�����jA"�"=�1�OEx�CjP�a�<��5�@d�CE@�
W��~�a�T�3$Ҍ9�r�iR��O���O* ���J�*e*2h��k�4���o���B��*20�ƕKʚ�w�4�3�-Y�����Tǉ�g_��p3Fc[���$`��	x��+Or��"'�A��� w��9s�8��аi�� 7�G�\`n�9c�
'�庍�D�?�t�t�G?�hE �_�%�����'���J$ȵG�4����t��5I& N�4����Ϗ.��h��,i�	�dJ2%���K&�Y�J��� (�D@���I�iI�'e�f}	LXƦ���Bl�(�DH�k�v�P%1��X*�!�#D	x�jU꙰RWh�'�t��F_�ԑ��`_5~(��O����'�|���d�]���y�5�f0�����$T!441���$,ݫ�놴K�B@G+�[��yI�j��:8nI�����tl�g�~��L���-�<�c�i�`Y�gϱ�?���S�g�L�ڌ��!vVtR�<ba�!'M� �)�'
�����F�)�<�ؓ�
rh�`��H[�h��d_o�Ƞ��c����ś_�:�x1/ ]M��s.#�O�!k�$L��v�:��b��a�"��5Q�18*�F�F@�t�UL��9��BU w뢝�O�т��N6 z<���. <_��U�	�oh@�d/0}X�h�o�T�&S�e$�*�y��&B�a�jj6���Ƃ��夁���6�I>v���d�U��J��kgI4��=o��l7j�F!S4;m�!��'�<"?1��5�n����;r��a�M3Y��0ʂ�'�T��b�9UR�Sf�)�����F�
A�6��D�����w���ц9�4�a��M�G�d#��S<_��{��Zr�:�����I ���bk��9���"~�⟼S��ʠa��̑D,B/oE���w�1}���s�U�3�]/=ƖA��a��y��Z�9+�X�y�5j_��V����S>��'R\�����+JP2VFB2�I��T�rq(���2$ 	c!�È{����Ɉ]�2����9��`B)	)&7���4[fjI;M*!)ՄQ;���!HN5z�n(�s�خl������!\qOT�W�1�d_&|H�Sz.��h�6��!J
b%�����p<AL�4((��wep�n�#>/�e��֭{C:����]��$[ן�Х�ֺ�5#,�t�ΰN56���4ֈ�qwL�=۶ a4��
_r�?AV�[������Y��lC�`Q�d[�hL�r�:H=���Z�6����#c'J�	50��� ��Ef��'H$�	�>�W�@R���M��k�<Mc�e��;p�P(ը<_T�����v�?��z�d���T*�Qd≙0v�Ъ�
�!!���J��'���g��z(���z�s<��v$�8�����҈g�Q��y�ΖS|&�t ��X�ଟ�����W�fZm�CH�2 ��8���~���	YK ]i礏ڼ���_1,��P�� �T���H�<��	�%y^i��H�m�
�����P�O�����O�RƤ���P&���u�)���?1A�E |���K��#H L��u��	��A�&�s��8�DD13����Ħ�bw
�"��)d��3���\
6'�L"v����$O99��(8�B�26�����4�򕑗����d!*g�,��C����-T�r���'Ѫ%���/�"�Μ�Sm��:Ē�[�F�:0r)���9xU�8�G$�Z�'�l�87f�?�d�R���d`���j�'�ԝ1�\r�)�tD"��韤 b�إ#ɷz��bAeP/�HX(k8�H��=Xλ��H���#�2x8�J.<N��'�������	xZp�s�%���v�x�zש�9I�4|�'ƍ#I�C��N#1���b,V Q��h��G�;��;�`߽��ɴ&-)Q��P�,�3�mǤMj��>fm�I�Ph: aJ�V��	S�N�!V�����F}��_��A��`Q���2C�<|ȸ�A��/��U�
�h��|F|��	�Y��Fíp�*��s���V�FhrG��H���	A�B�|��i�d�7�$XG~�n�+d�ֹ@@fKgD�̪*�n��@��d�$$6�pD�|rN�*�h�AK�!_�@w�A�;g����'���2s��yDi��ds��'] 8�9�d����]���@�'
�uRP�C'0�U)���ZȚ�b�'�`yB!�1LenL �,#	����'���h�A�""�j�kҬ$���'2�h0���s��=`!�u\����'q�����W���ó�n��PK
�'�<�[���۳�O�z��`���BV�<�t,��(�:��W�'����dOR�<�cɈ:bv��a�^�UB�/YG�<�JP�(f-��$u{���4�NE�<iH�]g�v��<��g��U�<� �� �&Di Arń�?W>d�P"OtAx0�Df+^iaE��/Nx��"O�s��E�,(���5O:�qH�"OJ%�G�,mf2�Z��j�~Uu"O`0����yʔ��+ì��Q"O�@)W��.��:���1<9��"O��!F�+.���0W/U�/j� �"O����X/� ��§C�F{��$"Old��W���e7z��x�"O�����&W�Rd��+|j�1;`"Ox@�p޴D��#��VM�a�7"OT��� 4�{`��63���"Ox骵ǎ
E�����$-� T�v"OJ�Kj@�(�!�@�G'e9@"O�I0gC�-=��1�ċ%�@q2�"O����v�������""Oh�3 ��aXFP@Rh)0��F"O�d�S�TB���S��L^ᛰ"OԘ3dJ�:0�|u�gM�B��"O�x�>�H�Ԣ��fe�"O$���X�3��|��'@l��2"OF�@@c�M�v�Pa� hp]�"O�!K���J�R��ב
^(l��"Ov]��oO������V.��"O"�)��i��ʄ�G*9��q"O
	�P��(	�R84-��	 ڍ��"O���D�Jx�Q�5+ �f;�W-�ybe�x�TZ�"��`L�Jf���y�aS���0�� �b��Nǡ&�!�S�&�aBAW�q����b��N!�䌒t�@ ��)!l0,Xe!@�gW!�DM*7t�%��'ò�p�o]&b�!�Z�'������H& b�kb�\�h�!��L�P��!S�ST�3D�J�!�$K�W�ҡ2��U�P>a1����!��T/]����Ȝ�+b��:m!��qd���#	#2��R��ԍ*!��ej�p����Mь@�!�dزf|�ZR�<s����^W�!��	z�p�b�"ΉX���S�ꆟv�!��>�6)C%d� v� ��@��!�$���81a�)l�ܱB�;�!�$��fN
I���،l  ���˾S�!�$��@K�f_$V���sh��M|!�$:5;X4X�ώF�ɀ�hW>M!���xL�#�Nz�˅n %@!�DÉC��!U+L�U��(1�@i�!�ò��k��lmAEKڃ}�!�Ø5P��,Ѣz�(�{�J�N�!�ď�ywf��3-Vn��$���V6"!�DXm�X���Q6|���+U��P�!�䌨q�����T�:�<A)޿:<!�dZ��l��֍�2#��ՎɐQ:!�$#VQ���t/�y\�ʣ [�bM!���K({���g�����oI�TG!��0P���t��,X�F�Q��'U-!�D	>y�,���Ը}P%i�#"Hv!��SqH��u����v�W�A�M�!�H�킀�č?�qY'�؎T�!��F�Kޜӓ�R�bH��e��?e!��۽U>�AJӌTb[��j�,�?^!�dnQ	`��+Q�����rU!�dGiht�� j�Td*�I&��[&!�dĆ&�0pX��T�ASh8񤒗>!�� x�s䧆)B�zو����&]��w"O��C�޿z!�SGLP~ٳg"OR�ˁ�P7-t0}����pa��"O��*קȆ@�nC��u[8���"O|��.�>���RrkISx�A�"O\Z�M�)>�`�����(<\I�"Oq�g���DZ�`�'�!���["OX�A��L�*����Z�R>bd�q"O�=ᦈ�;iJ��s̦1�D)�'"O6��E�O%&M� Ŭ��uZ䄸V"O����K�M�C�ݱpb�B�"Ov}P��׻������QQ�9b"O�0�$����a���?��"Odl���:Y]���SD��WѴ�$"Oơ���G��a���¸#��}��"OLP�q��AՈ�_[ Y�"O^l���;M�Je����7��(xT"O�P���O����4��s��y�'��0C"���#_���B��;nNz`
�'6*W.�
�29k�m��e^�Ѹ
�'�>Py%�T�EqMh���\C(T�
�'�"�
����W�xh�HA�Xq�ܰ�'�x�P3� �M���3�G\�d5����'0FX�+ǢM7�*�H:���'����`W��Ј��W�g���'�;�k�94�T�J���1�r��'��@�FS�%[l����� .�*���'+����&��*����E� �Mav"O�La,ԮI�^��RJ
��.l�%"OĈ�t�I��d0A1� �H;�Pa�"O�M�Ui҆^0�I���B�� "O6tb�T&�0�j%� �3�(͡`"O��K�!܌5���Ao�	��T"O��C5MR��� �_�X� "O�=����)f���J�,G�"����"O(Ar%.3����M!��s�"Ob���C��F]h
��f�5�""OnU#!�Y=<���@>���Q"O�+�cS

�^L���;;��(u"O�@�A�5�m2�!Ѳ�i�"O�H9�`^�[@���m�L����"O���ԬԄ#X��[��< �`�""O� �6q�@X�%��^�z�Xc"O\`�r}#F
]<!��S"O��0"�� *}�Y����(�5"Oڡ���мS�!���F��`3"O�6�աy�(���M-G2��g"O��%"�wl0	�F���b�"O��"e�z,j�h3v�4`��"O�l�橀�ST��k�'�ut��YS"O�1$�H#^]��E
DW�|I�"Oy�ӯ��X�.���%A�c|!{�"O  "�@�'�ljA�3$��(�u"O
�HS�F��*b3���x#"OfIiqoٿA��16�ǹCZM2�"O�����;(��;D�鈑��"O�Mp�cD�Vr����T9>� �A�"O���/�ҍ��o�l�2��s"O��"%S0;��mF�ٌ��T"O~l,-ўE��]!U�J	`vč8�y2�� <An��אL�H�dP�Py��5 �9��!=	�E�Y�<a@g�:s.���e؇{�5�kNQ�<�o�ZI�B@��kn�u�Le�<� �(  M��e�J5��J�@�<Л�"O���@���6�ެT��AJu"Of02�i��� :1�/{gd8"O�=�6U�u�ح�@��_�`)�"Oj�ٱ�V�'���So��T����"O�hK"�~����M�;Ot�"O�Y�W�B�n�h+O��"��XA�"O [��G+w�Z�ScN�f_��BW"O���Ta��9LDXa�/A%Z#"O��U�	&R���G@4/��"O�)c6#оd��b@'�]���"O��۴g�5?ڞ���F�v��)j"O�����ƭCOֵ�e�2�ੲ�"O���3+�1���i� �*�tt1�"OZec0�ǻ�U�$C�}�}�'"Oj�����z��p�"���`�%-�yR� J�v$�&\gx�رT�y�%Q<-�D�$" X��0�Ř��y��4D~��'�M-W�L��!'R��y2���#�|���"N2mȡ����6�y�FŖe�"�͈+!�.lr�����y��X?B�T#�(Ⱥ��i�����y҃թ[ ҁr�F	ʞP�a��
�y�"��PaR���J�~�q1f��y"
�Ą8�m�w^h(c��\�yL:6�Ќ�3ύ7^V2X��W��y�
�(�(���R���+ nڍ�yCD�)_�Y�1�P�\�97�2�yb�D|��7�R)H%6�٥��y��
!#�TR��I�(T�i���,�y�.�%]줤�5Cר#�� *Q��yT�H֚��F�EC��I@)/�y2e�I�6d�r�O#F+�	@�п�yR
H�������C,$���C�yRI؜`��[��C�lxڤ�Þ�yr�� Q��2���7�r�CD���y�C95��i7㍯g����V�yR�֕,��Bk� eŠih����y"	&`шQ!2��B�)�8�yr�6�ZiP@l)�����\�y¤M>?�J����Qo��x����y��@_�ɐ�gq�e��m�=�y"OJ#��h#�͗a�����I-��'�ў�O��H��������u	E�?$�	�'u����ٹRC@�a�X
�N���'7&!	��ս��(����'��f��W�@���
��l�~��'��Q+��٢nK����B�2a�Q
�'�ۃ�ƏG���R���53�(		�'n ��(12���O��+>a��'E��;G%=��M�rI�8:��}�'ĵ�f��J:�Q��,���	�'��<� ��Zb��*"CT�*�t �'�\q�V	��E閠�ѡ��-ۄup�'�ĩj4�I�$,)k�.xh����'b8��]�{�$����nB����'&������_x��ӭҰg�^���'�:(0GM�T[�psb�uDՀ�'�*M@c.� ����f�6%��'�d�tKE�@��5a�n��cQT9	�',H���C:��<Y	
���'@D����1��`Q�*A�T����'2�a�fܥ}�,�cfE'Ng����'g���Q�J&T��n�v�(
��� zP��c�58G�l0�C����"O����S�Uj�c)�^�q6"O:Щ@ �2FТ8��另Z�"�'"O\y�!(O�I�YY�E% �a2"Oe�u'
d�zj��9�3Q"O���3@�x��Մ��bAX"O�p%��D)��)gc�=0�����"OvSugɂ|�감��nO<��@"O�(q#  �E�g�2GTeHb"O�5�d�K��p
�"�t�S`"OV�9� �[�t��>.R�|�"O�e2 �
��H��/��LDZ�0�"Oة'/KD׬126(S�FB�M��"O: q�IX�,;꩐%Y�38D]Hq"Ov蚥J�$�P�B�[��Xi"OT��1�C���6�Z�U��C�"OPA��*�eL�4
���"Ot�!�d�<\�R�!0���~�h@�"OTɡ�K�cY����\��;"Ox܁���C2l ���.�.t@�"O.�{rIB*W���)�N��h��"O2��!�t djR�ߔP�"O���W�M�>ƾ�D�]1l��"O4s3���y��d�d�@ZH��P"O�9#��+x�`��b��? =���!"O��(�H�L�D�s�I�^�DD�6"O��J�M�(]n��W�@�dz(=�D"Ov�x�[�3]P}hb�"l �!�7"Otp	U���mh�C�-�t0 "O�����*RTp��P�,��"O���f�V<y!ڤ��D�+�|e��"O������r(e���A�(��T�"OXa��sYZ��Ăßm��P	"OB J5I��nbzy�qa@j���"O�,K�iÜ���u�ڮQ���a"O�x���\��8$s�`١}��Sc"O����~KC��b2�
9zn�"O��@p@�TD����Ӄeh$Qۖ"Ox����;`�<��k��6i���"O�� k�2�60;���rT�Q��"O���D	� ����Cj	9>�MJd"O`<)�/U�,f(a	��k�BL���>D�eE5h�n}��
�0�r�8��>D�<Y`���7P$òNS,_n��EN(D��� �W�M�C4
��.OX��f�!D�T(UhK��Z ǫC$t���+D��h@8�+��-i�@�F�(D��3t!E/x����`�7�`�am*D��BҮZ!i񖙰ubA	{>��&D��[��(#KHY�BkY=+iኀ�"D�@!�� +�L�w$يw����b"D�ܒ���/(�tI�0(�\�ɹ`` D�4���}<�,s"��"+Ϭ��T�9D� ;�!�5(��\t/�9?r��un6D�̸��X�H�bA� �3B��Z��2D�,��郐ip�a�Վ�>�����;D� ��6C�� �d�W1&� 9��.D����[�v� x +Ñw	��C�*D��*��@L�>Y	u��m2�A�"g,D�8���	o�(����JpQJ�&.D�x(�(��h��8gcE=�f#�,D��u�HW<��`��F� ���-D�@�X�E�B#��Aΐ�e/Κ��B�ɨN�5�C��8~Zq���țf� B�)� ��4���e�F�u�@��E"Ol��aL_�(0QC�+��z��.K�<!c-)�b]�`�A$:�P�@%Ck�<A�*�$ &pD�E��J�0l���^�<����1)����Fk\��|�JT��O�<��o�3�<q�tǕ A�&݊3cWt�<A�(�9�������2�RL�cʕm�<��Ŋ!F,�Y��2_Ȏ	����s�<���8�|�9��3T���q�<1�*j�:!��TW�� p�e�<� $6,@͠C��_��(�$c�<9�&�{:�I�5,� ��u�<����S��{2�E1;8���R��r�<��N�28�H4MޭW~H��kSc�<9�I�o����ҿh%@U��Z�<�@�4���o¸��S��V�<��#��7� ���MR0b�h�CĎ�m�<�o�?f�21"`�[2% ��S歍i�<�҅�7�����-q(
,��*L~�<�v�߼o���!K4�:-J%Ir�<A�Fr|�	�cՁh���p��]H�<�u勹j2�3��6��U��]�<�F.)v`�ؓ�O��9��ْ�d�V�<92��.X����杇8�9)�g�Q�<�7��?��B�CY�41Ѥ	E�<Y �EU�ܹ�K�4�6� @�<)fa�"ɠp(��$}佐��Q~�<a�1B��(��Ot� ��u�<�&�tL^�#c
ذ �F�k�<�"��hj`�vH�&pD�p�i�<�0Iǹ$�(,��	Jْ1']b�<)E�M�I*v��%���KE�t�<�Oס��x���L�l) 1�Ls�<�0胘'ǜE�����}�c�Uv�<ɴ�!ڔ�1qb��BU�t0�+It�<铆٬e���bB�	W�Z�s�HRq�<R�T�Kl�PӷŅ4]������H�<��k�mv�g쏄s� pCE��<��B�4i����'+��-$��?츅ȓAμD� �eYt�)Pj�`���x�9�f��c�x�(�L��
`)� џE<�0S�P�q����ȓ �
���Ҡr{uH�����`��Tab`Dٺ��/h���ȓw�b�ِ��Z����𭃶'����M�&F�q��"t藮)A�$���D�9W#`��XR������ȓntF5��cP�W9�P�P���)�ȓ,j0a�/��X��ɣ�uR\�ȓSV�S,^0MD"4 �'L6]����$�i���A��`m�4nC�Y�ȓ~WX�ҧ��)è0j�b2����ȓMB���fP(TCGf�%��4��I�rD�UC��\xZ��:q�-J����vQZ �V ��{�ą�vԲ�s��Pz�b/9��M��u���`J�c�j�"P��O|e�ȓ0
�p+�gG,|�� ��OX���=������eA�d>(Y��@�G榼cb'���y2N�E�<��^�>�LU2j)�y׿��	³�ٵ>5L����y�[,]����ЁW#_� HQ�����yBEã��;�R�P�(����4�y� ̜9�$�s��G]��y
� R�t�ڂ$^���*��TQ%"O�d�0��4.�-k0	�"�n�2�"O� j��hl��������ӕ"O�<s7k�8���Svǒ'v~��#�"O� 4Bş`.`�{$���6`��"O��!�	ʾ<S��s@�T��ơ�b"O��9BH�p^� �r�؎W��9�5O~��� ����Y��o��0�@Z&!��OT�V�@����֭Ŧ?q!�Ā
�A�(��<�Ѳ��W
,Z!�Q�@X�M��j��`�BiQ�F��!�$�2$#� 
E�D�U	���o�!��Md�-�U��&Q0Y�a�\�id!�$UI�T��aDUxّ0��4�!�$X	kp�K3l�4-D�����0�!���(9�( r	Y�b�x��&A*�!�Ď6�	v�_6niB�f��sl!��A����.<^1��{!��=n�a�ҍȻt}�q�$��h`!�Ę�L����l�tԵ�����#P!��(P�R-��%S9K���K5�_3^�!��ظC���/OD���Hߜk�!򄃴U����ȟ$�d�����!�d_�'ұ�".�2��<�F�<l!�$�]<�ŀQ�E�¨��j�Ch!�d� rlr�!�Κ<x���Y��P�S!�$Q�#������F���T�nC!���L���S��m��8R�mY�j!�d�;����&�s�B=���\\!�\�`��M��cQ)n+ `W�[�B��P�����/��g"��1$D""ͤ)���:lOp➴�t��3k��}��W
�j��e�-D��p���l +W��+@y�W�(D���� [�وt!&6pL@dj'D�(�GDA�d7�9)�f�%l�J��$	$T���M
e8�yD*��V"O�� �L�pTl���Ӌj��0�"OrE�Ϝ:��Ġ�CG�}@|qa��0�	L�'3ETY���å>7DՐR+	\qB���mޔ��!�AZ���QW��_}���z��`�NP'h1�J] a�Dl�ȓ,��X��@�&���ХM�~�l��o{��Rb+�&�N�"a�I�Aˮ ��/$T E'�l~2u�"ՇO~��ȓ�X,!6 ��n8@rŀ�}�̄�ȓ=�\-�#"���iGJ�* u��ȓX���ضC7�2����_�!+6��ȓy\�:�!u���� "
u,8-��@N�����?�2���M��J�� �ȓ"� �Ȗ�DF��X�c_�`p�� o���q%�:����\�ȓq6
48u��#S0��af٣_������l;WAC�,�h"���HJ���?��W!)[����$)	_����V��"h�5F2�M��)HT�v��ȓ�|�d�NM'� �+E�VrхȓT�:�Hc����s,�,1��H�ȓ'N��k��k��%	��Ѕȓ'騵;"���k��9Χ0lƙ�ȓ[U�����R�T�,aA2��
$�l�ȓ5tTlZbmR�"ypq臃�~5��g�� 	�$�*ɞ�U@ z����;ޮ�c��Ӵ~o"���j�8]���,j�8��#���(�*� W�9�����S�? <05gK �ޥ!�jB�S֒��U"O>��_�a����!j�]���"O�	�
�x�|UX�ɔ�S��1"Oh��@���ȇ�ݟA]D��p"OF�@3+���P��B�vRۣ"OH��ĩ�9.w�0�aa��c`B�Q"Ol�@d"@�o�t,�e�1,U
��"OD��&h�"I����U.ݣ3E�u��"O��G��(=�r�j�F؍f5Ή��"O)y��!C߲�"�^HL�PR"O�5iGoL�h������6͐-(�"O�cP�?,�d�! !�a\B� �"O�@�����<D�D`G�)���q"O���%�PL����ݱͪ��W"O���� (.����&, �"O���  �犌S��q�$��"Oڑ��K��%���g�Ҿ$��"O���h	Xz��'_�Y��}�B"O~)D��6V���LӽF�LQk1"O�1§�ـ�\�	Q�7ɀ�+�"O�! ��4
��zw�A�8�6�ڐ"O�-��
&Ii�!!��H�u����"O��A��;P�d�S�(��P"O� [W��1'�<\�E�CS��"ON�*B˃ or��tJ@"�v�35"O��t�νaod��J�2ٮ�2�"Oj�2��'_�]b��3���U"O�!	�<��AQčȩ(�t�"O�@P5�͸1�R�`g�62!�P�"Od�Q���\��I�1�J#ymS'"O:}BA d�s�$��X�� "O���I�� p&�VE���"O�!��2~�ry��ķ+��-�"O�<Q ѕ�^i��E�fgՁ"OP+�#`��
�k���W"O�|;҉<-t���N�c��a "O���70a�u�v�M��j�"O��s�bTi�E���x�:l!d"Oͻă�: �2�̘="|l��"O��� �W7B|�g��M�FX�#"O"���B@&"�Jq�����b"OR���G%<i�<���|	r�$�?�y��")*�;�̅L=Jy���y"㋰�J�Yaȍ�qY��yn��Eӕ�fL�P� ��y�E�'/Z�.�]�Tp����yb�6c8�c�R�Rp�AfZ�y2D݉J�8�-&J?�a��@ʎ�y"�X?t"�!1K��j���jZ�yBE�o�@�H� kPq!/^
�y��ҳ@���'���w�f�'#K��yr
N&~ 
�"�MFr D�AЖ�yRA؅>���!
:p(P9 ���yr�@�V"��E˴:{PWm/�y�eˮm
\�W�.=�v���yb��<G���1ݵ(J�jD��y� X
#�PS�'���#"F��yrcנy�J�@���P�>�R����yҡ��
�|�hջK��y����:�y���$~.L���*.2��v]��y�ە]�~�R� [2|�@�I$��yRc�%=ȃ�1K�VjM�&�0�y���m�> �t�N;EjԀì��y�Y80���E�V��>X����y
� ���.R63� `�Ou�A�"O�1���A�lQ�0��/<�~��"O�0kЈ஼�3�ڼ�\��v"Op[�
�`��0GI��xC��iW"Ox�"��p�z%i7�h�B"O�ճa� 2pD�E�a��Q1f"O�l���T�P.�$قD�U"O
�A�44=1���)��i!�"O��3GcW�{~ry �c�$��"ObTBdG�����%gX�qgZEx0"O��!��������lY�_Ԙ�7"O�``���$��둘;X i)�"O�� �ޜv���Ɗz�H���"O��I�#��/:d��`j� >4z"O6�ib�JH9����;`}8�"O艃� ��%'�"r>���d�í�yr��;!t�I+v�Wj^�T�C"��y��n��9�'�J3��ĸ�K�y�)�
ku(�7V��4KC
��y��j�q�B��H�b�%��y��^�q�ڥ���:�J��0���y�l�>/�x��Mۉ���
�J3�y���$
����� ��4�����ә�y����ibl��n��
���yb
J�W�^�0%)�w�Zu����y"DŦ	S�@a��J6c���3%���y��O�
�Xe���e��;e��yL�	��e��Y(��d�Q*�yrG���P�ʀ�"���Z��yC��P��%a��}��y�lA�yR�߮~Fx�0b��rZ�i6���y�l��?�ȉ{��X>qb0#�O��y" �<0��!F��d1l�H�bY��y���A��xY ID
a�f\@ H��yr/ЦCx�+�FM�h�T��R���y�P��)r�X)f��e�ӊ�y���j�:����_��
 _�yiO�h�q��U����'���y��Ӵ*�4�T�GNL����1�y�j˕k8�)��9�ެ&hY��yRŃ�3�&,�b�S�#��,�t�B��y�9	FS&�L���-_F�����N8IW��E����&�Tl�� ��c"�P`ʂ�$�h� P�@\����pUH䑓ǒ�:>��Y�� <�ȓ)���з"��
��y$�λD�<ńȓ�֌�F:c�&����Xz�ȓ-HZ�#��dXPW+� ���-J�=�0!�>�@Xt@,!�0�ȓz��v쐬G(�k�D�/2������,�#f��($J(I۲N�~��	��8n]�$@J�"�D�B�&ф?�t�ȓ�q��f�0z��jE�Jv��O���z� �Q��-B�"]?|Xl��fm<�	���mB�e��a��#�t(@0���zqlف�%�:(�0��ȓ:�Ҩ�cJ �Tn�9 ��7�����u(�)�,��I�xk�0CD�ȓ[����0�Kb��2�l,i�\�����*#�Ԩg(Qj�A�4�8ń�(��yV��?�ސa���#�X���v����'�$�BxA"��>іŅ�!׮x� �Ss�4�gA\���9�ȓeh؋��W�Q؜�`ug� ��i��S�? T���ꔏ?�r�8A�V<�n ��"O��B��z�P�ƀV�C�RP��"O���bㆴ'�����ϊ�a�fup"O~ �2#�'CXܐ �n�.H�27"O��A�H�5 xY��B)�ղ�"O�=a im�4<y�"�IN��"O0I�e�=78>�x���*��`�"O �F�C���`3M�-�z�s"O�	!2d�(mL6�Eŉ!�A��"O���"`\$�XJW�����a"OFKD,**�������~�LL2�"O�UX��wdd�K���4)�D��"OL��`�'GR�1��՛jhܸR"O~4;5鍣i��{gH��E�P��"Oҽ:���(5Vb�� �N�P4�D"Oris"�Nh&4!��A40��A�%"O�9
�� ���"&V�}-��3"Ota�C�p,@����J*`+�"O8�Xr�ҥO&���f�
(��2"OP�+���_:~Ib�Bɯ:"���""O�Af�������#xL8�"OJ���/X�D�L(�FlP�D��#�"O�Lx�����ي���
�(��y�M�=u���Ć�G�Ԑ� H��y/�<x���g�B1���qN��y�Q��֨� )�5F� �Q��.�yR�� T2�HB���7� �X B^�yY�Mi���J�E�<�v%��y"I��X` b�·�qR�`�!��Y�'��-9�/C�A3ZAzEgO�y `1�'5�}��h�n\dy0�h���8�'M��x�%�A�h��C,Op��'�F�:�	�U�h��"�6��3�'���H�<~ąPc���4UR�';�5�����|��ч]� �<�I�'j�h�b@D.���B��0A>��'�$r��\Tr�"*�t ��'���!�h7�䋡�[�X�D8#�'�l�Z��U
U���g֘I���*�'DҬũF��'N�o�Д"�'PNP��ҏb0\ e@\1X�4A�
�'Ԝyb�l�⨨�%
%PQ�M�	�'����A��GD��"3��|o�]�	�'��e�c�MY;^�1��N	
b�r
�'�4���"NEǜ�� �D$u��i�'+��i��A�&=n�2a�_lNtz
�'Y @��ZU�A�	2h:��	�'��`��ξb�z8�Ԝrf�̑
�'d��(��N���i���j
�'��d *M$#n (a� e�͂	�'�Dz dO2'�<`Y��\�+ V�)	�'_�� ���H�PR.�qi= 	�'�ܥ�.�0%9.y���v
(\r�'hR0Ip��J�)r&�v�&y��'sX�Ir��D�c�@�g� t2�'�@E�"��j�~�Ht���]�$-0�'b��ã��"]!��Qw�59�'V�%��I V�� 5)��P�����'pу�
�<��`�L�Ab
e��'[�)K#+�62$+��5j�Y�
�'� ���
95_Y�r!��[pJQ�
�'X6d����)R������>D�	�'�L$� �q<F���!O�@)a�'�0U��M�,�V!���#:�H9���� � �։Dz�L����1Vj�a"Ob����1�`Ite�?V^�1"O\\���Нr�zi�M@�=�<�#"O&�
�<}4j���G+f�@D"O�tq�����iu�����"O�jW���¸��G�/�L�"O�����>_�񰷥ĳ7��$"O��{A<<±� $C%�PH"O^�S���&�Щ`�䎞?ȡ#�"O����զj �T3։J/;}̵A�"O���kt(��G�A���R"Oz y!d�!l�.I#�AݘO60EE"O������8(�]"��U�;�&|x�"O�O�W�x0���B ��|��"O6�* 	���b1�rC� %T�,��"O�Db]�O��x���=��ȕ"O�� �SSkVl� �%i����"OX��O�1cq�P�`W�%Oʔz�"O8��פ'N�5���0}�n̡�"O�y��;�*����F�	˶U
�"O��sr�M�[Z�V��x���0"O@���@B
4�>uj�AC��4��"O��h���?w�̡Hu@P��!�"O���h8�0��$�$��=��"OH|Bg�4FY�)@�xm�2�"O�|k�
I�3zN���:f��p"O�)��#ݰb��(�B � uAlQ�v"O^9�2lP7oe�f'&n�!"Ot�Ӏ�͞t��P$[:O�(�y�"O� �)GYr��`Û�*-�y��"O�X�c)�� ��k�!#&��J�"O�9bŃPc8�Z���G ���'"O y*�Ϻ:.�Py����s*�!��"O���&���3f��l��%{"�s"O�9��#�-`s���WK�G{F�2�"Olغ�䞪3Yf)�'l�s&|[�"O�[�gQ>60�-��� ZU�$�"O��0�HҳU����Ve]�d�e�3"O�aY��8v�����c�b�&�pA"O:9 mӷX�l�e�$U�ɣ"O|X���Gڨ:v�J�ĭ��"O,�"��	I��\ӓH
<B��A"O�q��=�09�3�wg�@�"ODkr� #V�I��S
� ��"O�|�lD&�R��Z�T�U"O�q���=WbX ���y�2upf"Of}�Ǥ��W�xHs��Vߞ���"O���fG�0<�tY�tg�_��5Ȃ"Od*�_[�|���h��1�b�#"OR���D�� m,�ca�v��P"O6�RT�Wd��Ҕ�±a�x$�q"O�8�F�N��T(�ۤ{��}�2�0D�(�@ED� �����}��A�c"D�\���5ز����6k����� D�<Z��:��5!���j�@p�1D��u 0B9���7Ɏ�Pys�,D��e��)���vċ�
��c&0D�l��ဌ�XȫwEKMyf"-D�h�G���I��D��ɑ�tr"��)D�X�U��
�@#)O�=�̩ځb<D��I���L)h����fU� j�<��퓥FN���<�pկ�{�<�թɜp��`�rO�.BD��JS�<Q� ]�	�2�$,υ(�f���O�<� �<ccA14��S`�
y�0"Oځ"��%S	.��t�(Y.�%5"OJр��u���$/ӣB�t�"O�2iV?,Ȳ�BNؐ$��t+"Od�3��˵�Ԩ`mT�~���`�"Oz���I�s��;�l9!��MR�"OLp�/J���R��$�%:s"O���q�Ϻ<�ؑk�5~���"O�X�e.Xj�A��:V��}��"O0h`�%[t��u����a�$"O�ը�H�r� �P���'l���b"O����9}�=	��"��Dx*Ov�s�Q�f"�a�(�6o`��'(���@�ӜNp�e㣭}��h��'�"LIe�̢W��x�j�^�J�'Q�|�V̍9_^�}�2-�xH �'0d�	 KGO'����Ɲ ����
�'X޴��āצ�q���%o����'�~!��<Pj�p�G;X�Y�'T�!�2I�q�j�;����m�ʓ,��i�F92!11��
�� �)J&M�-��Ё�+�Z��ȓl�Xh*�!�h�H�7�Ǳ!]���ȓn��O��%B���d�ȓk�Ѣ�)Ly�`����gi\-��[���˓��d`���2�>����ȓ+��	�E(׋rH"�{珎%,<�<��o����뗱ݴ�s�Q?�Bh�ȓ[��%`p�R=��d�S�o�ʭ��.2f� d��b塀3䪔�r�v�ȓa�~с��^�r/���C�4:H�ȓSu�I�u[�@���WL�.q�чȓ��h(�jY�����N)i�vՆȓC^���	޲}���cf˦S� ���e�@bߘ'Z�0t���	���ȓ+6�����j�8�jE�V5~��UH��x��4v��+M-�  �ȓ%�`|����W��Kbb�`Z���S���'��G�.I���%:�X���]�V���0 �ar"ʑ�`��фȓQ��eb��v|�ʓ��;���ð��7A�?t�
�)%�1O��B�I3SF��9�T+������o�B䉭>�ɹ�ϙ>�*! ��ϜCƦB䉳Yo�,�"φq��4�����s�B�I�Ic85��!>���G�Ë��C䉁L$1	TD��_��=ap���
��C�Ip����gl��H��Y1&�^'w�\C䉌[?��g��-Eh�x+3k�"[�C�I�{�z5��E̜A&�D����e^hC�I�G/��*r؊0��8"���J]�C�ɽ:���R!�X��\�uiB+��C��4 B�E�A$׍�~u�޴vh�B�ɛr]0A ��_�~�+�$ܫ2;�B�	�a^��tFV�R�2A
�S�B䉕p`�9He݋l�V�2���-p�fB�I�)�U)6@�$}2��ƙW�PB��|z����Oj[Ɯɰ
�",1(B�I+W ]���Ǜ^�v�Ѓ֤%�B�I#u��:e��H?X��#jU4B�IU �5hˌ';B�`���N�C�	6rD�yc��E8;��X!6��5��䁁hk�H+�B�"6�ȉ�g��D`!򄈽I�n���ȝY}��D�y^!�� ���&�V�C�=JB�1x����"O�@!�革�HLP��
:AH�x�"O̻�*�14M�S�S?آA��"O8�f��D�~�c»QҊ1K�"O�8S��H�T��M��ɥP�|�r�"O�Q;4K��)n>�s"�͈J�~}k�"O��
�逕cwЩ���=t&�`1"O:xC��N�Y������7~&%�"OJ ��ܒ?��J�Y��8��N&D�Dz��ӑ�L-��+�a� !D�h���2C�xq+�埙<�c�=D����7M�}
q�@/g����:D��k( MR|�&�8!�px��f8D�XCam]�`�qK��īˀ-��K7D��AW�B'!4�!Cf� "s%`	��3D�����5C2��b�ФI�n-D�DA�ܱxU������Alt��q/+D���#B�&X�����0�\�c2E<D�@���$y�%$]�R�a�:D�4����;�� � nY�>U�=D��§��* ��I&��+q� �bQc6D�p#�f���@tϙ�&^���H4D�8*�%�s�`�!�0���KMDC�ɶ�F=�,���z���ܰwzC��baa��_J�ɐ�Հl�4B�I-	��M�X�AV�ТԩF!SBtC��(Qx��@�G��g�ʬ��nFB�B�	<P��*��a�	��	��B�ɛm����E�&����aB�L�.B�	���i!�B�(슬�%�[�7&PC䉾Z|�JW.Rĉ(ul[32�C䉼)��#�K#���$0�C�I�٤Y�4d�-�$����՞��C�I"Jޜe��J��o��0	� �B����h�1�U� ��x`�D�4Z��C�ɏK\��
U^�8��2 ��C�	�L�4�	�"ٍ�V}yr��~�\C䉡7q�b�V3p�6qQ�F�C�C�Ɍ`Q�IZ��7Q��<�r��|��C�I�q�*�����6V��y�䈕>\�C䉔^��9h��yv��S1c�%
Z�C�M*��1C�Q�p������C�I`m���� ��!�S��B�I/C�^�@��R�C��]kP�ՎV�C�H��Y7J�cO���� O+��C�I%�2i��BA�yR|�{��O�Y�C�Ia�
���ʮC�Z5c�$��B�I�Y���z�@� "�[Á�3;|B䉈t��Ҁ,�>Wuz�IG�h�C�I 7U���&�2:M�4c��D(��B�,|(�ё��$l��$Ã��-o��B�Is,L�٦�%v���r M^�urC�	Yl�-!f�?7��1S��%&�TC�ɴ��9�5∃xbjH���8�@C�$_�$��jڑ[�<��Ő4m`�B��8��T��f�1sl�J�'��Q��B�	�/y^��S�լ=9Fu�&ʠT\�B�I�v���X�g�y2t%+�B��;f�����C۠y�0�X�f��Pq�B�Kٚ��H&`Ch�� ��s��B�I����z�LMF8у*Z�pC���� `Ҳ�
9����"N�B�I1*���?��$@�I�4Q��C䉚y�� �4��yDȨ��kY*(�B�)� ��e݋.�B�A�E�'+PSe"O��:Ro�.sXإe͔Mq�"O�}��EA�6��@�p喑^�p��0"O=
���?�p�)VĆ*��@"O2AZ��C.vH V��a��Y�"O�܂2LD�C��$Z�˵i�����"O$eY��ElH���
$��09�"O��pUF�o�ʨ�T韷3����"OZE&-7T$�Dzf�S��3"�-�yR�7Yʪ���`�%Su"e�����yB	N1a$����>H����"��y2��x�6TX��I���ҡ�y�)=xj������$���C�y��Уi�!+�K	z%�mr�C�y�`ב7D��F;`�0��l��y�g�+?p� $ :[g��U��y�\�p��e`wmE�VԖ	���O��y"
H�;�T�""S`ҭA5G�8�y���5Zx$Bq��b����y�Z,"���М:G�*fE��y�O
�Vy���J�C�$�:�yBN�E,�h���<J�\��'���y��VEt����(��,zu����y��Ń_�i�AΑ�!�N�s0�P�y�3c{B���N����r@A�yҤ��w	tuy�)��P��7�ߪ�yb��>xy
��%�	!,��!�V��y��6"�4P�II�|2D��j��y"��2,�d�+��'4�����y� |�&IKH�n�����y2��@�JDwl�&�:)i����y��N�GwtuKB`����5�]�y��\m�M�4㗰}�ȡ*4����y�G*6�����s��KF*�yBAQ&��d�vw��]�h�"�y2j	_������0k׺8�dA���y�-�.�� ;Є�k<�Q�S���y�D�_���zW�ĉf���cB���yr�-��H�$�Gt׊P�G����yg�6{*��E@=pF ig+T�y23\5�栆�4VD#W����y©�(�
T9tb�!/�@8@S��yR��^,fвЯ4.E���E�ǌ�y2�E�<�H��FѐpS�]ؕ�Q3�y��8T`�|[���=%�i��H��y��2��x��KȦ5b,�D�M��y��m<����n^�&��	#�J-�yB Y�{:�����)Ǌz2����y�%�==�U0K�	@�����y���$s�݊D�	1B )um��yr�����P%@����BG�] �y� �5�f�{��R�,IFO�y�	ɑ��} $�Fw� �����y��Y<9|��F���8`&���y��T4-O*dH$���+BB��a��y�dS@f
T��%gv�!�*�	�y�
KF�f��!�/I���D-ʙ�y���,��`�h	�H���6��yB�ѣnS6�H�I�B�9�Ŭ�y��,GV�ZP��[ �$�B��yRkKL&����F��Jm�S���y�*�1kQ��̈�/Fȼ��d�*�y��1p�1HP�ݭ�J��A��yBH {U�����9��au�V��y
� |{ �9ni��6Ș�f��	��"OZ9j7��5
6n]pG���!x�"�"O���3�S�Z�Ҭ�*T�g��"O���D�9A)D9t,_jl#�"Ol�[)_!�l�6p�(��"OD�����im�)Z�fG�n�$0�"OR�1DM|ڒa����O��+�"OR���M-:�c�g�禙  "O�����UK.��ƍ��Uٞ�""O�$��߸<�*h����-Ďe�!"O�}�1/C�a�����JI9 & �`"O:h����%t`�x��(h�5k�"Oօ��G�E8�U��(
b2	�"O�x"�'�$-�E��XD]xC"O(42�)	���2N�64HQ[ "OK]Sv��S�+��Q ���#h@8�y2nۋ=|^ECՅG���S#�ֿ�y��Z&Eg0��*��r�s�yBh�Kr�[�N��01��q@��y"��!_��%Z�؁%�t�;1�ʘ�yj]<4y���&8=|葁��y�#��r��+�I7�x�K1B���y�A׺0ǎ��ej3*/n}b����y�&β>	� ��U*�ЊG���y��n���'l>$�T�3���y�,;3h�L2�L�B}���V:�y��C�
�E�'&�{�d=��`�"�y�揙N�f��Tlʕt�dA��&ȑ�y�e��R�RzZ�t[��r���ȓjE
'CO#~��1KQ��d��>�l���۞$Cv�Ց/V%��qc(G���8���X�Dt���
. �1�Y�$���{[�<�ȓ@�H�BR�ʈJ�h�k��;�Ņȓ.�6�)0��3�Ҳe�7 H��ȓx�l���ա�5�6�ݴ:; �ȓv����t"�f��ghU;vQ�%�ȓpvK���|��I�2oV��bd��\�0]9 �Ňhn֔1��Z&R�T(�ȓ�8I�� ��H�ʅy4�"	#���S 4)�M�?�:�R�!��t�l}�ȓd��)`�A��IjCbJ�t���ȓw�Y��
�����Q�D���t4��
�)��^\�<�K�\m,�ȓ8�4�@$	��R�G�)_�,��*�9ّ ¹�X��W�D�m�V�� �����	D�ƕQ"#=@Ąȓ6�&A!e"��tI�����_�>]��O�1x�i�g�2���2b�j��ȓ|3���VF!7P�a'�14l���B���Vf�`�B<a�Y�oM�L��a(6u�$��#r:.T 2nQ>Sz�y�ȓ=EX�c�)y���;Q4�}��>D�2�c�W����).Y��y��u��R҈Ŏ~�r�ء�а��-�����?F�N�;"N�t���ȓy�=7��'x��rCD�6�=�ȓT�8�c,��q$�h�ѡ�)? �]�ȓ
���C!	�kX,�a$j�"x!�ȓ^�����٭;I ��fB�o���<24)�V�)+�,�Y��!pm�]��![Zi�Ȟ�e&�]A1#˛2^L�ȓDu��z�a�/J���Y�!F<S���R�~�[wJ˩J ��9#�
5����S�? �)%9�d9It�F<��5m:D���� ϝV�p�g��?<�ܑe�6D�,��k�4h��L@\��IEH5D��ӓˁ- �����cK?W�X��w
&D�lq�
n�F$*��BPE�Qo"D���QӰ5��D�X-�h3� D�Xw��=x���e� ����@�1D�\I�WE�� �)�"����)D��+�&�M0�r�����dA*D��(�@Ď-�vؐwi�L�teA�'D��!��_����AĪ$�p��aL"D��:�	�dc��@�x\�:b�$D��b��Ѫ!���9��39'%D�@���V�)-:��I�/����G$D�T9�I�z�ꥑ�(d�>W�K!�$@�xA���r��uk5N�$'�!��O.Wb� ig���V��k ��!�$�CÉd�P5�ඔ��'Ͳ�b̀�\\Rh �dC2s�ؕ2�'J�%����[�̝�v�=;�'�����9ˍ�*ǒ(��ɑ"O�y��J�1|XHc��_dޅ1F"O���rsı:iZ�/Gĉ�R"O���
��w�p݂�Ψ!<Z�`%"Op}a5��`0(h�َ 
,2v"O�1�NV�pP��4@��ѐ"O�XQ�&\4]����7�!��bR"O�3oJ�cg�UqB��>���"O�$��H���!�A�I��5"O�) vL*D���*�d�24��ԡ�"O�ѱ�O+9=�a#�@�*`�"OЛB�I�V&�&ǌ!^���"O�(���-�r9�0c��nmx`"O�a0ɚ"Zh���a��<�y"OX�u�C80���)��̗sV Yؒ"O&i2���:��@v@_3F���a"O����j�>GP������K�z�"OzP2�R1���
�����}�"O�� ҇�e+|��*_t�x�C"O�M��)�����=䰰�b"O��&�͉CZ4�f�;E����"O�F�G�nI�8Z�A�Æ\��"Or%�W(0Kq��w!��~¬Б"O�Ie G�h��U��/W�Dv��"O�U`�$6w�}S3h�F�Ԛg"O�E�2��d(N���g�sD~�E"O��;�?\��r�/$)��˴"O�ҕ�G�u��JQ�!r!��
�"O��e�
+������Ҹ4w�M��"O�8�u�B�>}�-B�(�:m����"O^���.���$Z3�u��Q"O�<�U�}���Q!J�C`�Q�s"O����E����T�͡;BBT(B"O��@�Fw� 8P �T�+�d��!"O��i�M
("3���	X��@�"O��k��ł	x\�
�D�����"O6�G/�^9`e	�5��8�p"O��R�ϟ�ؠ{e���X����e"O��J6�7�����hi�p�P"O>`j��4L�UZ�'��,C�"O�}c�,��?�ʥ8�oT�x�"O�5�ȞtJ�Ũ��SN��3"OD���B��Z��ȣp�C3�����"O��_�P��ȑG��;舱�e"O� ��qSh�,]����+J2ٲh��"Oh @�α<��邩�y��	Pv"OT�����r���Чn��20����"O�x)���RⱣU��V @PAu"O��c��i#a�ՌЌ�����y�D�y�tI�&]r�H���@��y�`�$h��KP��9{f��Ԅ��y�	N;*��R��L
7J��W&ܐ�y��݋m.T9����0�dA�G���y���K=���g�;0�j�8w���y���V:�[C�'-"�⦈��y2�]�NI�B����ը�A��yB�K�?��d�#�|�c����y�i'
���1�7=�� S��y��������h��`�'���y�E�@�X��$�+zޜ�w
	�yb,չe60��C Ż�t	����y�#�l`�I�1ER����V ���yr'R:?HL�@���E�v����y��"�ۆ!B;h�nu���yBF�c8�Xdd�(M��(� �yr ˀe 3&�V��1�*���y�
A�̝�V��-J��\�r�[�y�"�)q5��9v���YQ�`ReA<�y��v"��DĂz���(A�M��y��-�z͙�CS�;;[2��,�y"C%-8�y
G�J�=���q��'�y��5yR���\39��!��̈.�y�GũE�8����1�bu) �6�y2o��\����f��`D�I:��"�y�,�(id�����1R��FeJ<�y��R;j��kO�r1L[&c��y�⑐z� ��� d�����X=�y�D2]U��
\�U)`���I	�y sהE�B�-C�p��-��yr��I�)��J_h D\�O�:�y"$x�r���B/a.z��b
	��y���'3�d�#�OďY�ꅙB%�yrP�p� �Co�}lu�aN��y�jK%yk��CM�7B6;QBC��y	�r����54<�u���P��yLt�ܪ�HK)W�<!+E����'�ўb>A�u�׌k�j}Y`�@�|�H�0�;D����J�u�����ٔ2Xd ���:D��� B��b�!�$�ط)�6�rt�3D��`f��+'���pk�9����2D�L�2CT�$�Ac�(� 6+�貕m2D�����Cs��PO</cv84�.D�x�(��D�+�JN�IZb�7D� ����2�x��!؇+��i���9D�0�Fd����ք,=Ι�s�8D�lȕ���!^vp1ej/-�`�`8T��"���H�� A�A���%N4D��dc�$�.9��'I3(^�Cj'D�L�T��~@2,R/}�jQ 9D����=�TK�	O35�i;�5D�� t�8_�P%d�[��R3#4D���î��E�b������3����RB&D�(�SCů ���ѩZ	� ��
#D����伐�Y�����?D�8�gA;O�����ٳ&J�h�7(0D�p��DD�>�Q(F%��T�qm/D�Ġ�.�[J* ��X�W�4�6(9D�l�p��	z�X�hUX/gn�ʃO7D�� h@� ���.�Y�#��&v�RdZ6"Ob�HǉZ�Vbh��S�r���"r"O�`c�o 2�69{��E(��h�"O�,�EX0G�NY��ͫZx��"O�9J �C��&�I�>��0�"O�`��#G��Ģ��և@� !"OPӡ%�'�L����1z� ��"O��@��&��dr���XE*""O^T��J�2Q�z����K�(rV!��"OR-�0�Ph��M�2[ƭ!f"O\9�q�%P���!-��R"OB��!4|J��b�*�N)�Q"O�Ų����E� U��@�Cچ�[u"O��b�aN*�d
&R�q��y��"O�|[�II<�@P׋�f�Qv"O�Ijl}JÂjӻU���!"O�D��.�>=^mB��l2T���`~M�4"ά)�"�,�h�,t�ȓL-j�rjU� �Q��̑���ȓ��H�"�@����oʔ&�ن�EDI�ڗqu\�g��8���ȓA�~}��H^�Ma�gD3=
x|��m��Xra@'��ʴD�/.�Շ�B�z�X'�Hq���膅S��5��=4�QJta�,>.�5��,�n��x�ȓ+*��uCö6��R!aј0�����^��Bqd]���	e�)����'H�[��@�;�:a�q*�#xϖ1��'��qB�(D����"��wYVMi�'��a���ΙdP����V=��'{4��"Ԥ_IxDH�%[�=���'�N��?A��Y�H3%Vp
�'���CFOG7C��Q�����]l��'��W�!(�W���E�`��	�'4l��1aN�5��t���U�G�	�'m:��MK3TӪ�	�#��:��5��'�^1 :#9$��a��$���'�xق�*[<&[����
�@(Z�'V�l{T,��>]�,��۴��I�'F�5���rX�X�a(�Z�:�'$��gZ ��Z�#Y�#D��'\����'�jy94��N����',�)��_,q��x�I�/�N���'Bd�y��O�j� ���Y�(���'�������$7�ňf�X�tQ	�';j��a�ߥ�z�@�ԮP�Z|!	�'Ǌ)��n�24��%)aNV0��:�'?ra�5��>.sp�CG��8��D��'��M�bl�'=QjP���I��t�'�>��B�>�8���I
'(��-��'k0��Æ�^��1:&׃���b�':D;�j��B�p��U�ЬjԹ+�'�$$��d��tz.*,���0j�'E��� ���K�4#�I�:uzq��'��d˓n�;M�]�S揙:Jt,�'���K��	[̾�hToɟ>�̓�'��'��3��%�&Nmha�	�'����O�0���5 ���S����K]�)�d|�e��Jh���ȓ_�-�M�/*U	��\��0��r�Ԫ�.R�;^���UÂ�n��ȓoz�ٳ�éR8�Q���? ��ȓ]�
��,ŏ�
�hV��:4����ȓT���DC׉t��H��T�r����S�? �����N]�=:��-	�b"O@}�D�Ħ<����I�h��[S"Ot���bƜ%���$�ܵs����"O�z6���, �dKU�<�!�"Oz�1���0�f�A�ʚ�z�<��p"O�)XV����p)��6��-�q"O���WP1FpP(փR�RS"O
E�găEC������+��T��"O�\�!�L�
�3l$��5;�"O����`��b��I�i�r"O:����Bd�%���˱��و�"O������7K�1�6�itv���"O�r�ƃ�QǼ��M��GfN���"O�X	t�<؀e{c�I�Xi��ʳ"O�吲@��t����)GNNxi"OblA��.
+B�(���?RP���"O���F>G��m*�̋-6�X0p"Op(��Iu���0NѲ"���[6*OU����b}��`V�/mE�D��'c�py�˕���Ʌ��._�pt��'v�@�"������u,L�Z�t�)�'dD!M�M6
(�%�S�T|��'���(�%��Qzz|��"T����'xV�`l�>Vn(�����Q�~�3�'��x�&+�
9�J���<����'���3J��Nc�+!)�5�"��'�6� ����+��-)Yw�6���'f����+ O�*@x6bS{ʡ�
�'���zDg�;|B6�I��=yg�<0�'�8��4ͪ}a�-�VȚ��q�'�<��i�=u��.���Dk�'��L�R�ΰO�:��4I[�����'�4�pD`�C,���$���j�
�'g�����x
����
/�4��'8�̓�G�4d��.k�t���')�[�P��@��]�V>D|3�'���i�,W�}b�c&�?Djd��'{H����	����DdX'6,���'h���j�' l(�i�j�,m���#��bs� \A!�)˚���MG��`��L���90ɟR����ȓv���PT�H��8������M�ȓ&�"	r�ǅ-V,ı׬e �ȓ.1b�P�M�� p9�i�����ȓ;�>�5B^�3��m�槅�b�B��,�r��U���zf��#�i��:���k�M�c�HF@I�dJ@� <���OMh�(������
#�D�ȓm~��V�A�k����s ��,� <��A�r��%T88�,�
Eʅ�X&���ȓt�&���/M�h�,2��7R�4��-K���E	/��J'��2V� ��1���D#�RP����S�"l�ȓc��y�W*UnZ���߿>�,��q���!�A�<u�=���U9w��\��-�|�BcO!�>���m
 L�R���b�ݳfj��-�+[�@Y�ńȓNP��֎�19由��(����D�ʓ��c3J�$�jY�J�@C.B�$L� �v)I��6�{V+_�j�B䉀^9��Q�L�%P
�Z�L�v�B䉱-�����@�Eʼ����D^��C�I!LTf��,�=t�~�X�+C��C�I<�mR�H�#2�|{ӆK��VB�)� �0)L�2�*b��8鲁��"OZ�:�&�r�Д�&�݁z���"O�q#u"�%�v<hPE�/-˸-�"O0}��el�i�IH7 ��H:�"O(uJ�j� ���	��+�4�r�"O>�b�c�8{8e攮~���W"OZ�{&���@�֪L�3v���V"Oi�K=qFt����d�}P�"O`5�WA�}�r=Ņ,Pֹ�"O�E� fC�t!E�g6b���"O|�z��H,/�Dd��Gz&�q"ONDSc���Z�r�� S�\��$"O^�/�P���BA!
�e�t���"O�yC�n�c���`7ǒ"*xKe"OX�Q�$F�&��:YrM��"O���q�4MTmB���C&�� "O`��aʺ7Ĕ�pÌ�& � :�"OȄ�'��m7�q+j�{R�=�&"O~k2��(]l|��"C^<�@"OH-Ip��Q�B-����5"�!��v�<�A�L�Jo&uk�c�	�!��{H�Xy#��$�JE0S �7G�!��Sa�t����9N���I��!���Ig��!#LQ�Gq��S��A�!��n\sB`TA�����L�\N(����rAʣI -(� ,iċ�&� �ȓB��`�#\�HI�$A')��A|�����]	6H�b��{H��ȓE��p2,��1=����9���X�����HX���R��w�J�ȓ3�,��c8h�1�!Q��ȓ>uR�	՗T���+	 �􀸅ʓ<���:�J�Hpe��� E3�B�	������H@���G/g�C�ɀk� 
��H�3Fp�P+I��C�	�s�
�ثk�^����>�B�ɗ=N��Q�҈&�Ne��E�R��B�ɀRSҪ{.mad�|�C��-=L:�$	=F�V�H��R�C�ɲq/�+�Y�㄀�Aa^I��B�	�?�@�0���8�
�KB v$ B����ȁ��[>7�� �^�-�C��p������N�!�}(T#�'t�fB䉪,c�L[� ߼	���A%,!OvC�	W�f�;���b����3B3�B�I���c�Ȏ�rg"��b� i�C�2���� ��M/ �Cǫ����C��Dk�M�Dj��U�<t�P�C,Gp�C�ɑ&r�ux��,��<B�C�
YZ�b��뉙R��hPhS "̎��`��%k�B�	-Ky�S��ЄJQ8���aAm�zB�	��>�!�,č����|�NB䉒��R�^�i ���G"�[o@B�I�EO �3Ǎ`�ڢ�5�:B�	�c�"([D���Hڷ-������&D�i���&�v��0ZKz�࣮7D�ȣ"i"Hg����h����3ad2D�T�Zr���m�"��+&�.D�x�Vl̳V�LQG�ƅv��h� )D��a��=8��X�IC+ ��A�I%D�� �/:C`�`0�l�$-���Ƨ.D�ܫ���e;�U{Ǉ% Ȑ�+D�lH���RM8шjo+A��y��W;�~`�qh�0B3�4��݀�y
� Fe� �J��lE"��[�G�3c"O��q�À9y"A�`�,0��"OX�W�L����%|�Vy��"O�b�^������׿��q5"O��E�T�B�|���K�;��}�"Ol�q��:v""�&+�!F^�({ "O4��tNB1P�t��J��g6t5��"OTe�'�%�\hJ��è3?�@"�"Ov��"c��l(���2J����"Oؐ0�hˁ(H�e�~/��0"O����z�(hX��t�Hр"O�Lag��w!Ԭ҃*�jK�5 w"O$����1$�lX���]�Q��X82"O�Ĺ&��~X�ձ���w9�ط"O��R�lЧ$�hy0#i	�g}�x�t"Op�[�O	`�¬��$mB�<��"O�tɄ�6 �����C 
'pu"O��q�Z9�~��⁞c8!�r"Ov���m
�,����#B܆f�3"O��UI �5eJ��ᖊ0����"O��)�b�2~<U�tVZ�P�Kv"O�ps�- �p-�ek3 V����?��?��x���0Ȟ<x����Y	=j���ȓ*����# � -�\b��)%���<qM��Z��	��a4�����L=4j�(#n�!�ɧBf�e��К -,y��M�N��'�a|B��Pnܥh���<qWEa":�y��.m�N�P�(�mC(�Ī��M˝'Ha~��ǤIZ�]b��RaE\Us��V��䓐hOq�6�8��?Q`$��Mo��""Or]��^�1�yv�O�US*u���|B]��F��'QTH��l��%j�aP��)v�|��'�lP�r�G�M�H2�ԏf�j�3�y2�0ғ��fp�r�Ɛ����wIK8KL��	e̓�?I��̸q����%���Z"�)Z���M����		".�u�c�3������0b��x�|ΰ�d����r�y���Gƺ���3D�Xj�J�iU���PV��ȁ�&D��`�A#u(eeI��Y`b-�#�"D� SbԴ1���V�/+-��{�C#��0<����"��gcX�&v�C���|8�@EzbĀ2=]T�ac��,-`t� E&	��y�,�M��WK�$)|��A�mҺ�y)�.w=6��'!)�<���U��y��D�䭢s�6 ��ED��(Oң=�O�Z%����;"Bxh�����R�ȕ`
�'���'C$a�"�:��Pqr��N�L��yR���� ��i1���0d6�Z4���OT�O���<1�FUVW��:0͖D�Ճ��d8��af`V�E�N� '┦6 )hFo,�����=�~���
Ep��Z#0�xA �	YW�<Ig�ڼ>>�����%"����WU�'�yR����r��+Y�H$�А��M�\B≿N�ȸ˴#�8Z��h�r�z��b��'����䤟\�~jg�L=V�8���� ����妉^�<iF��hKʉSFHR�D8Tz��X}b�)ҧ_�Ʃr��"iG$H9w��S~�<)������OJ"MY�) �|�n�I!a��k߂��'����io�|B-QNp���k�+)0����6ў�>&���OW T��}B�m_kJ&�R7΀�x��":�v�v"�;^���DA�#���Ħ�D{��.�%-'�`��ɞd�:�D!U3��?i�'|�9��DB~�x�yu엾77^ R�'S�aI�]=H�*��q�C5��$���ا� ���E���#T�hB��+C�IqX�d��"Y9'��tH'�h�s�)��hO��26Mj��ABȈg�"٨���u��B��=wը�j�۔ra0LBWǐ�y��b�X �R)�y"��D�?i1W�Q����Uv��cUi,�Ofʓ�m�@�Ә`�}qF����*�)��@�e�zT�8�V΄0#�d���%���O4����������$8�b�!���Zd�7D���4"�9Kt��Q'@� �4���4D� ���Ds��G�>��H`�4D�܃qdW68z*��J��~B����"7ғ�axBD�&2���b��Ȩ	8��gMG��y�`@u�@�������&!�3���dK�� #��P�v����!X�O""<ю����f��� � ����Je	M�yr���s+T���F �> �Q�ܺ�y�K�sꨄ(�π�)�2�������y�HN$t�	 �sք	���:���XE��'��zP�� y�	 k3ve�Q	�'���g��~�~�2�gW*#�L��4�PxBɤV���E�Z�m�>a�Q���=��3�ċ�' ^��FA��⼺� H�G�!�ͨc�	���(-��	�iK 	���E{ʟ&�� ��ia;� �X���IF"O�����d� ��   |�v�@��+�S��y�,�H8��p��d����G��yR�Yl�j��D��;�=��4�~b�'��	�SN��GD���e@�U�^.Oآ=�O�2:O��2%��,xzxy�)�
���:O���$5Air�d�4��u�0&ȷ%�	s�Dl�Nh����?�
`f��a�xY8� UJ"�hh��-�O��'t�Q��� L����qi� XA�U)s�i��'0��"���<���䐐g���W�H ��Ď,�݆�׶Ě�䁻H����*��r?Z���hO �=�Q),,��t-L�4k&d�Z�X��$0�al.T�ѠW���d�߂�z����جaR
ţ{��ͺ3��ج]Gy��|��CKw�DJ@��'J�Ș��+�s8�$8N�H��Ѭg�D���A2u�ti3�j6D�1�p9�8��� Z~@�(
3D�,���D�7|�$�P���t}�8{��'g�X��xl̴0 HTE�
���'m,�zSԮ�!�,m��	��'g���ï>*�\�U�B�`��A�'�d6�	F��~n�#Y$�� ���!���y�F�uM���j;u���Q��$�M��O¹%��A��d�E��,[�eéh|�1�f�66����$!�D�<��\}�v��"���.��B'Oҟ<�?Y���OZ�)s�*�*|x��Vu��3C�	�<9��ə9e���J�7��R�
V��D4�Oz�T�ѹ�]P$�G!B>�Id[�tE{�Op�'&RuP�k������� ��Vg�<ɂ��z�.�������k�x?I�'�&����� aJ�0�
 .u4�#���.�a}b�yE�_�.��m�a0d��'W��hO�����&r�xX'���'�������+��xF{ʟ� sFh���r7����]sL�2g!��K5H�i�4+33\�Ȗ��=����>�������� C�7
�"p^0 �'��v�Ҷ$�J�kTD�Ka�ȂAi��yr�Xڟd�~�Ӻ[��$ nH]@�C�<��j��Qj�<�聡'���;$H�$\8���ke�<�s�K�w9���4N�"qüC�C]i�<�5$�R~t�H�V,�hap�~�<� �Eƥk��0Vg� O0xؠ�IR>�Ñ��y ��k˸@SbP���&D��I�X0�����N�T�4�"�e�$��O27���~���i�j9C�`�5t��ң�Օ}����'��(;��)~Q�%��zɪ���i��$ܯ��V�O�Y�S�y"ˉ�f���	���i2����	��<%��_�A|�YTz,25SǦضA3
�mZw(<I��F�7hl}9��'�T����S�D=�d!�i�|��BY:20���t��%5{B��T�����X�v���,ģp@'���'%ax��6hn��IGOs�ڼ�C	�y��S�R%x���uP������ybhQv�j4ӕH&YgZ�]��y����@�&��(��;��ͥ�y���AhL��ȏ�֦�(Vn��y��Ѧz4 ���}�f��e���y���gT��y�E�{.,��ȫ�y2*M�:Ւ}�AO��n[���(R��yRd�3p�`��E�R`����%-Ǚ�y�$ُ2$B Z6J��tK��� �y��#�uCÅ@3�����y�@�
K��ػ� Ϣ&s�ɑvh(�yI�:B�@�F힃#�<�1g^��y�'� {�^)�+��\�7L6�y��ަG\��"�]�P�&��yB(�#'}&���
F4H��`�y�M �3�h�P5@�x��C����y�����eM��"[d-��cߐ�y2�� f�P����h(L��Ã��y�Mn���`����L"�y"M�	j�vd8c��3FbؑK$���y���
x�*��a$��6�z<�ң���yr�[�EM�6��1z�x( �)Z�I�!��@�=�;��7B�ʝ�H��[�!��ߡM�P���F�%����U5mC!� e�vԩ�êC����'�\/N!�$S�\\9pʝ�2�7�	o;!��p�D�A��+"o�)Je('�!�$�(c����3��5|���ƌ�[�!�D���бy��R�x��Ypw%�D_!���'R>���O�2 �l��7d�}�!��mP\�p�O�#m��q��|�!���!�>��LF�kR�0�Q{!��F+5��L�7Y�r<`G�4!!򤁽X,!��d�+(�h4(��]r3!�˾y�ĥ��`V)oTeh��V�4�!�$��(�ҳn��a�`i��NVG�!��0S ��Mz����P�!�dښZ�"PȂ�'a����!�D�J@h�8S�a�.ĨC��q}!�Dҝ{�,���f�+�� �w䃤ag!�č4m^<�4c�1b�p�r��αp�!���,]t�+3-V�T}P�K���!�$�L��a��[`��{G��ht!��ޅ=z�iG�?rԄS��@(Q!���2$��`�Aٞ �H����2I�!�U
T(5O9W�aX�bY�.�!�D�;����d��a��!�0:h�)S��U��u��{O!�$T�h؄�P����F���А͍|+!�$�.�|5��O�:�X�r-�*!�_�En�B@�T��\���^�%�!�dς0(&4���|����r���"�!��4x"<5'��L�6�ct��^�!�� ���uW�^��Er%
N�^��	c"O�MatK�8J�����H�#.��"Ol���M� =�Pa3v'�; `�
7"O�㤜>���p𥐻1a��f"Ol�p�eUB�}��&EB�M�"O8	괄�n�jI��ղ5<�x�"O��J�6hD0 �b[&}J=�C"O� �� ��r�a,q6N�1g"O��ږ��ji��s ��@4�"O��㐎n'i�#��!ry�E�"O�P��?w'��Yg(�.�cu"OP�I��ZXV�C5�����"O�`��:f]ޥ�p�R�Y�H(��"Or��2���-��P��H%p�~С�"O>%��	��N�(@Uǁ)���c�"OpTIw&O*>��VI;���a�"O@|c$��J\�ES���t�n��"O�m2#�Ĉں�U��8P��"O�Ɋd'Z�EB�n_�=I�"O��z�n�-NҀx9N��n��j�"O��`�X+	������X��4��"O5��̂?[b��P�O�����"Op��V��4�
2�X�NG�e(@"Oz\P ��$3� K�&M@E��PW"OB �`��=n�PJg�ð
Af|��"O&�#��"Y�ը�[�s=��{"OL��ƀ�3(L0XR�d�bÔ"O��{�HT�G.�;u"}��dف"O6����x�^%� ��1;�"Hf"OZ��.o��"d"U��E�"OHt&��%6r8�@� t8,q�"O�P� NL3�f����?����7"O�qH�"�8xa �����[�H�S"O�����Q��!'����ެ2d"Of�qpşh-LD�V�L(�4q�&"O&�`��U�FD���C�kh�᫆"O.��ӭ$�0-Ja�T42�Viye"O(-
i�:4;�YQ�'0�x���"O��A!�V8E�̸���-�μ�"O>չa�I�0�h8����>�H�S"O��clǷe�}rwE�`�l�ӱ"O�}���^�0�Ѣd�*e�$E��"O�q������HacĽA��Q�"O�'R.n
���b���n�I�"OؔhgV�4'�H{��� W|Y�"OLc�cͫM��(F��0C�M�r"O֡��&�1O��;���m(
�s�"OjD�#���gU�(`A'�?h,M��"O��k��#3���D&Z��!���'��I�GO0�0 �� i+�0J7	��8B�ɉ=�>�#���0C��r��л36-=��ƌ��H]ʥH��
�d4�EK�;D���皏J|"f#ʝg tE��`4D�i'��H�����H�n�V�3c ?D��#$p�*� ȭQE,��
9D���u��20�1P˓'aa�5$1D���	� 8���x�o�$FGJ���<D�(����x��2j��48ׁ<D�xsQ��H`HW�$���f�;D���r�G�=\�Z�o��Ww~}Y�k8D�����`�$-�����;D�D#�ˤ>0��AA� �T�����:D��Q5�Z��졃a1=�f����4D�|���ןz�Ա�a2`�K�h=D�� ny�e)�50#@�8�:~Lu�"O�Q�`���}+ &r�P�e"OR(r���%��u����#��;V"OB!�D��?�\}��Md�X�"ON%�䈦D�X-H�Ș�e&�"O�c�%�u���Շ(���"O�T��f
= ݊ŀ��0Ԗ�5"O�ӓ�/bm#S���-�Y�"Oz�5�4D���Xv/U�? �x��"O`�q��X*��s�����t�J"O�X�$(F)6 �IyR�ԢjPa�"O��`%�C���g�E�)s��2"O�|�Ң]��a'��(c���1"OU�7�?Q��!�0�߁BJ�M) "Ol�C Y5�|�"`�!?I��"OhP0��T)�T�*�@̺@7��r�"O�s.�<lR�C`�+Yy��D"O���Ŭ�� Ɋ��� �%s���"Oz�U�!V���z�H�B�Z�"O�EZ�C[�Q�Z��0�_h!<��S*O��ȑ�ΐ�t�"��2�ʱ��'Qz���[��n�"�β!�j8��'ٛ�ۗk������o\��A"O��k��RwL�k��U-��XU"OV1�W	�C��R`FF�6Yq"OTP鴨�R�h��E�O���"O}��ڳ:���#P?dP�H�"O���D�?��e�Ņ]Th��A"O
�.
,Z�� 3����	�@�)�"O�0�֫]�R�*� ��^�9��uX%"O���V,!N=��b�ʍN����"Of��1M��L��M�g�F�j����"O�R����7&�H��7�8�"O�]��K�8��=(��+@�g"O�i����1ӢR5`┩�"O�TqGl��~GFU��U-'y��e"ON�ȓ��;6L�!��ׇyd�Eyd"O���OU1L�2 �4a��Gb�q��"O��Р�ǚZ� ]�3!%o�u�"O�l�$�3�=�щ�y�jG"O-�lA�E ��rI���U��>LO�<b!�J�xP���qA�:ٮ��"Oj��Ud#���bj�:��[7"O�lf#T��`�j����؛�"O������.<�z�r�4�l��""O�$��U>]c6@��T,0�`$I4"O��ajX5@O>t�����J!���"OX�HBAĖ58���W�u�0"O��D�}}}X�����yr"OPȣPV7L��0�����> Z"O4���Q��MI�"H�C�,j�"Or�3M�$@���`��?j��rD"O��4/E �����ɰD|���"OI�n�$i��}��`ND�B�c�"O�	��B�L��d��A�`8���"O�� fT����� ���lD��˃"O���D�ο	�}���9OV�1�"O��ea�a@@X�ǀ�u�z��"O~�	��-bT�ahG�]B�jE1�"O�ġV'�/ ��d�e��$c`"O,�Ѥ	�:��s��و>�jP)�"O���H�<溔z�IK
��8Q��D:LO���M�M�\�6�Z�h�p$�S"OZ,�׋]�bȞe��+~
4��b"O� DK�a��d6FrC�ɖ`�D�j�"OJ�ˁD�-�Ќb��'p��0�!"O�آ��7��@K�CE��X&"O�!���&v�(�J��=`�N��q"OB���NΪH�&�J&�+�8�A"O.��R��pBu��K��cv���"O�X!���2� j�d�Ky��E"O�:��9�@����&*a���"Of03�_{p�0�CTAF"O�t�7�ڒ)>
LY����3?Xxd"O\����G)<��O#�M�"O�y�͚x�b s��m:��"O����$�K2�q��f�N|�"O���dJ;z`*�厚)����"O������r06Y���-����W"O�d�d�D�%ᴬ����>�T	�"O�!S ��ĦuH1�D�>=��"O��ґL��RS��c��?���"O�L��*�$Dq�(� ��P��" "OV�q�f[*�҄��O>$���"Oʍ��.l��0NR�N(����"O�-����k�yVk�+� �	�"O�$�0�ѐP�8q���7`�s`"O�1�`�6tN�˰��i.f�8"OEKƃ
�bA�Ug�0�0*�"O��2�È	2w�����%"O����͌i��9���>d�r �"O� (ŋP�!�.d+�)�'�h"O�x;�Ü�l���P@��#c��"O ��P,� _���闾c�J�!""O\�j�D�`�輚��B�p�fM(�"O�a8s/��w6����]�cQF	�"OPD��)̀.,�4��M
n=.�I�"O�a�&�ʛ(��!��ܦiؔ�G"O$�s ��+Q5�p�z��#u"OR�{���?wY
9Pq]�5�$*D"OijȕS�6�R!��9C���s�"O��HA	Űu��d,kl%q�"O�(piߜ ��q�+�L���"Oh��@�݇{���!�F�h3��¥"OF7��u ��A���<;"����"O��
@��5�(��D�3v
^<yc"O|UC2��(/#�yzv�^�B
p�;s"O@�z��P0�h�4�_
�1��"O\����Z�`qX���'/N(s�"Oh��"�dI�����a��jA"OܥdA�4��እ�� �H0�"O~�ucۉ�@xa��1x��s"Ou{��Y�n������\,k'"O(��T�ȼy��u �$��`H""O<�*$#� �va�AI�P��9 "O�X¤��_b�����?a����"O�ذFIV�bVV��HI)D���!2"O@�u��646��Ň���`"O�����A�mI�B'��2��4 #"O"9��K]  < �"�N(eL+�"O���a�$i�<:��^^Z�t�`�LH�2bf $����$��Wn�8����o��@C�b�{�!����
��R�g�:o���O��!��#z�}yg��C��1��ǭ�!��@� L�."jdY6'��A�!�$�}�B�G�FX�4B�G̪]!�D�=G�n���N�#>�L�"���
�!�DO
l�r���$��%����ފw�!�� �!"V���D�����*���2Y��"O<X��o�T����CЪAx,則"O��q&��5��P���M�q*V"OE�k[&A (щ�`ل Ŵ��"O�Dy%A��c#�R@�"{UF��"OT�¡��&��I�qn�17��{�"O,�FB�[�r(Zw��=;��Z�"OVQ@���CaȜ`�될�ٙ�"O"�� ���+/�Q��#|�A�"O^�R1NG�GʘE��2`�Ub""OR���%E3�<�y�I��z�ZY�"O�0����i�3f՛$ ����"O���G䏅|�Q�� �<2y�"O����1�X���,Xg:�(�"O@�ⳤ��!TB��a,�'A	�"O�PГ��
g\�I� )��֜���"O���!GG�m @ʙC��I�% 'D�$h��H�pqМ�� D�F�M D���pED�O����2KY�X)��#D�K�[?\i�����3*�$��$D��H�`�zO������-��p4�%D����fL*Qo�����"�`F,D��[����#�&ba]R @��y� �
g+�%�g�	e4TR �3�y�_^�P���X�Y�s�L��y�I�&Mܹ�1�X.Q_�����%�y�т"�\
#
�{�؄i���yҫ0U���b�O
sa�t@�B�b���$ȕ ��82���H	��`j[5Waz���(_'���V蟑Y�I��J�={!���:�� �(]yf �&B�1oy1Od�=�|B�b�/<࢐)����j�㢉M�<�dԮ!� BR��_8
]K�J�<i��'��J������k#eID�<�6d��.�j����ƥfRP�Hu��@�<���_,��cY��9�D�(CB�6>�)�E�mv�8�Cf\>N��B�	�w��ec9+�j�Z�$�5Jz�B�	8 F-�v� /�L�P+��p-�B��P�8S�	%,6$�%U3�rB�	�-%�PXF��h�4e�r�R�MvB�	5y��]A�"��z<ũB���,�hB�� ]�|ђ��
�+)�.[�}C�ɠp΢s��N�$gј�k�$K�B��t�8<�tO�;L`�����K��B�	�9��p`dW%a�~!*C�Ӣ<��B�I�~���#U�Au��0 �~�C�	�@��
�T�3(R������z)�B�ɺO��c�Υ=X0��e���B�	�/��`�Rz(:�be �7\6B�I):t�-�e�,rJD�qp`�xTB�	*� aH�+�(i�gR�A�B�I>~��k$㈪�<���,\�^�C�ɴG[�؁�Ľ_4�qRb�"j�C�}p�{ebK)!���+�M�0�C�I��ӥ�0r=����܆cw>B������c�?w� bG[�%1�C��+^�m��&؋:��(b!S)x��C�	�d�P��F�H�R����
��V2�C��N�~mRE�?�lR#Ǜ�
��C�	}��ᢖȏ�	J*�@oխ\J�B�I�.��#H�_<�G��)\Y�B�	*��#u�ؿ*��q	�f|�C�ɰyH�m�!�P�e�1:�fʌ&��C�)� �����1���1��LB\x�Q"O�uA�.�7RɊ�@EL�����8�"Oژ9� P���U�엋<�-�"O�C�FB�XH����ۼ��"O�}�SiU5�h�� ���m��A"O��mR"�2�ӄc�6'�(�[�"O�e"ƥ������c��Ơ�"ON��-]�h��0�G�&	r�"O"�� FB�%� �AAC;Z���3"O���C�=&V�У��	2x |3�"O�ARb��'�n���;]җ��~8��r�+�Nc��0%FG��%���9D���C��O�4��6Mw���q @x�
B�I<�|c� �֨M��O5Buѣ�7�0<!�{��/'c�=�e��W��qʖ���0=�b��]�<�']�U[�ƾVu�1�!�aP\��'x�cTcSC;|�x��A�.F&�Љy�%�4+L(��=�|��&�AOZ��%l�R����E�<!U�;f�\����X9\����-��WB��l�&�/�g~2�T,0���-�t�A�R��yb+�f4��*�4S�(��Q�)���3^� ��j�S�����5h���i�j���91�D���y�*_+��-)6��T���́|m80���H���I��Bf�!�X�}T��5�Q�Mp�ؗf܃U��'�� h��͹�k5�O*�"1�����$a`�0��L�%"�ب)��_�<�BDά/>VD0��Ъ�,� �_�-A��Ҳ�Ea���!�B���5�}L<a���`��|3�+:bA� ��y<i�AF�b> r��E�NN�`j��<:΍`FC�~V�x�D���tك�<O8�&� �Z(D��
*���ɸ"�>�e��d)*�k呣� D�����Pd^C�ɭH�`�%C?|�
��W��&���/��Gx��}��'�ة!�&f�ʘ����@5��:D����Z$��9JU��-���YQ"��+^��ۋ�����?��$������� �(����dǠ:o7�C�7"�y@A螐E%8�IdZ�m:�Dy����CU"D����I�t�h%o*�p?R5j���݃_���Cn�"	���[��/no��|؟��u���ww�`��Tr�Z� ����S�@B�S���xB��j4H9+��׆e 2\���@5�y�g�4f'T�VcP'^;��@o<�yBfP yаpA���F������̸�y2���,OZU��
�OXq"VgF�yr�\��J(0?��[Ï���y��B="�^�I!M��L�y�	�y2)�T[d�X�¾�m�b���y���u��9d�Q�pI�F����y�
���Fh�`��&���vL	��y��ݨM��9Ys���_|�5GI�y��ю.�8�r���Y�%єĀ�p<��D�q}C ��A� 	�7��MS!�M-T|�Mb�CY�R��Aҭ�GH��hO�|@S�U+Q�D����5x � j�"O�!�آJ@L;��@2e� !Hd�9lOdzr�I�$v]� )���Q�
O7���	����GB@�0�O�-k$<��6��\�gҵ!\�m3�h�*j�\����Q�'
��B�`��zpf�W�GB*��	�'�~t�U��'_@�FÕ>)^وI������' �O|m[!,
�t^F]��ȳmN̐"O���sD�sy������q�Ni�;�x؞��J��5��#�[9.l��%}R*D�s^�8`I<1��Գi��30oC�i�8Ek��$X���	�'+2M���Ͽ��2(��R=8�b�D~�%Є�b@ԟ�"=�eK� ��KgO����y�#��Z؟CSK֋�� ruD�DvD�v�ټdk�7��C�B�qG�N���O��ݺcd��5�h������t����^-:B�b3m��a�Z>�BV�Y"ر�靝)�Z ���<�T؞|Za��Z#���S�)<�~���/����lW�w\�u��}�:���ϐWHtc�b�\Y|��@�Yu�<1��'�b���$Y�G�.j��2�a�i��4ÆH��D��˟�܋�*M� �f��������-�O�� ��PbP���d�4�S6�,Ɇ\�`eA&4��z�/}�Li�#>�5(ފ(��Mr�.�����e�'� �c��:Oȑ!�@�� ~��'L�p��GO�$ ʐ�g�
+y��ȓ ��Ҋ\ �jPk FX�H� ���A�)G6m�aХ���?�9���g�(���'2�6��#�$D�H8��޽}��d"\�1`��bJ�7���+�4s�F�+sC/6]TE���W.����/u>D x���%�%a(T�H�P�(b\�]?�-Q\�)3b�k���Ä­yҼ�se��>Q�V�ƙ�4��-�����*G5��OV͉E
E�W����$��X��O64Ȓ�R�K3IQ���>t�,\
�'����S98@�����m����'���9` ���M�t'��$���=	%8qH��?R�d�P"O�`+���BDe˦2��DsPd�g���	)EW�x�-��C�g��^g���;�ݸgd��W�P��� K���g�O<EZ��B��Y�j!��C���{�eɩ�0?��-�ot��`����dh��h�A�'o���V�7��qO?��'�ݷ4>�e8�k�Ij"!�!D�8��gH(+�nd:�,@6^^����?}b�ـm�:�j�y������f$���7k$Ի����y"���H���M��1Q�	�y��BDJt�0O�c6m့�y�nO�5����g�0[:��kAbؾ�yr'0/Vz���dP���ʠa���yR�-4����	d�(��w��>�y"�C,�P�(�<�N8AǉX�yb�H�R�R� �R))�������y�E�.RAy�.ùU-T���RJ��TBAJ+�'7މ#3�M �(���̌�u�ȓz՞�pɔf��ѕS�/���ȓ.k@�rR'��]�|t�ɠDO�A�	�'t����mѸ�	��>{�����·a-��!���!���a�����fӀT2,����۬+C!�d�v��5 U,G9 �-��>F!�dQ)�R����%�T��b?y3!�);YbE#�M�� |�Y��1!�$LVUx�eZy;�q�P��K!��
H�>mk�o�0&Lx�"!u�!�dĵpB&�9���82�<8�������N�ui������h sB͋�yB�҂�^,Y���eq�죄C�6�y��ǫF�� �bA�3^5�`�.�.�y�)�	`�	�����"��:s&^��yb̚25�R�2c�9A[�q3����yh�z�� B��;�x�Gϓ�yR��&2��̩�.D��}I' G�y"Ē={,L(�e�
�<U�|����y҂B,}�) ��04`89ђN/�y2��e���S!�"4i�� nD��y��Ê'b6���Mԟ(, ����=�y����V>|R���]� !�g�y"#��3"ưZ�,D.`,��f2�yr"Y,;����@"�!/���ء�D��y���rn8�gOR�N��0*E�yB+��s���������0����y.�b&.!*����p�*V?�y2g�J��j� �HF=xu�R�y��7W/>�x���Y���e��y
� ��M�< )�h��G0F	Z�"O T�vH�gK���3�\k=�} �"O,��w�V�R`���9}xvdR�"O�-���Z$�����h`�	j�"On�A� ÒCTzdj���1Il��QG"O�x6��5C�b�8@n`qq#"O�0
0$/Pd���\~1�g"O�@8�c�!	|ɘVj�8p`�J�"O@��GB55ot��&�_c�"��f"OX�RM/Y�|��jD����6"O��PmE6R�"�ȕH�"M�NM�"O��� (@%W�N%t�M	]��D:�"O�dц�F�I� a�!��x�h�P"OB��%&K���\��kY9 r�a3"O�9�̴J1d��+@�C��i�"OV��U��ذ��G�Y�K��Ei�"O�C�+�-P5�U � ���r]i�"O6|񶧈-�xI&��$$v�� "O��4+�"���;��.A��:"ORU(�.�%*�
�в��pm�5�y�d߿bH��	��Ė~R�<�&����yj�=]��(�EV�i�B���!���y"��l:�j�#��b$�ìS�yB�[�PJ0���<J6ż�y�.ԜG-�DP�%D4U����#�?�yb+O�l�rmiq�p����Wa���yrGU�xg��+�a�91b���[��y2 0�F P�(�(A.%����y��^��ތ�Q�9�&@sE
Z3�y�%38~�i*Ĕ�5�֌�t���y"��V���A�l[ 7����N��y�ݧh"hZ�h�*ژ�I<�y�W�UqRe�H� ����#�yBN�9V�N���͋2���u���y�E�A�4 r��!{��A�?�y�ӫa� �D��� *�Q����y"�0N`lF I�I�B�y�QITI��[
�Z�'E��yR˗:J�S!��R�6a�iƝ�yR�/Y�VU��`ٹ�\��
���y2�A�%r�W1� ,a��y2f�����D*I�1N�+!��6�yĞ�g��ԊU�X#1�!�y2�((�Q%��K���Z���yRY�Z̽a����G$�A�����y�Þ�z,6 �pB�=�����8�yR��li�����*IP�X�,��y��ިW�x@sb+ɮ~��X&&�>�y"�*B�oE~����yRC(�d�9�ת� x�N���yŌ�5�t��o�n���҇�yb��o�a�FI�Z0z4��E��y�H�yQ����L?��i�\;�yR�̉'^8��P7=.t1 7�Ņ�y2/S����0Jʏ|q6���y�H^�_�>Q)���4�%�H�oE�ȓp!\�Q�G��k7��j%'upr���l�Isi[ D<���ږA�1��;[\�� ��:n��PVO��w�~��ȓ	"B\!����9��E��,����ȓyJę�e'�Dnf��sM�^H8��*Ԑ��Y�:f\IH�KRI�)�ȓ��3�g˰�F�XS��?!����PtvmG�:��9� ��@��t��S�? .��s.Q.ZU�)N�c�"OxI�/��Gf����:f/*�"OLu�u��G�0k�*�J	z|�"O��CA�bw$�RC��8V[!+�"O��t#�.!�<�@�%� kn�m�"O���ԧ:O@�K�a�+!\��3w"Od\�fFׯg�&���Á1�~p��"O(�d��T�\�����Es�"OJ}s kĴip��Ud�W��h�E"O��pi�h�db��&����"O�d2� 
=  ༓r��L��I��"O^0�2FT�e��U �
z��iX�"O�;���p��D��	��jp8��"O^���)R�	�bf,���"OvIQ֯�^C8y�F#(��p�f"O|��7o�v�P&c�_�~�@"O�Q��"lr4�c�� ]�^D�2"O~�I6 �%z��*q@��L ��"O\�a��[�e$�]b��]��1P"OI�bB�lƈx��)	S((�� "O�r1�W%m��:t���dJY�r"O&� ħU!�%�G��� ���"O�d��ۊ^��ypB���*�"O��k�
IQ2�� ��_�����"O��c���
��ƭ�E���"Oj�0A�gMZ]��,�.:�Нk�"OA���:JRb8١ń�H�"O� qԧ����+��-�<�!f"OVQ7g^0P��H#��vmN���"O��S���Z�5��ɱc���""Ob�1����*S�$˧�A�~|Qs�"O�	y�+��(���H�,�咶�ϙ�yr�\
%p�pF�Ŵ'��٧G
;�yb��U�a4k@��H���KJ,�yRI"P�D�x��E�H aF�M��y����a��c�i�2�sa���yb��'�(�"e�T�>�����yB ʢ�*�ۥ�&�����]��y��
���M�!^�Dh�n��yB��)nxi�-B.7�rQ#�
�(�yB��#a�9z��#"�R���A�;�y�	��12д2�j��(;nLJw�T�y"Ƙ�0��t'u�Ԍچ �#�y��:v��� Z�bD��S���y"A�H5�@�tB�gu6�;��U�y��F��(�"�@�M7z��N��yRMI�z]���Ɛ�H��x�A�V��y�gK�#ÂD�v��
5���"J6�y"�!�>\��L� F!B�d׽�y�X��|�i_�TH���B����yeM��ÇعO�K͛��yRF��NhF�!�b�@���Bi���y�-�R �lF��5�,��.�y�R*���Y"���0#�'+������L(�/�.C8����V 
Y ��ȓ���!�`�87Cޝ�ᬑ�WI���N�jd����Ô�
~�$C�I>FXz	Gœ�^ǲ���H.�RC��M�hԹ'�H�s�|�d�y��B�I�C��Ł�`G0I^@�Y�@tB��dϬ8hf̈́~�0]J㍉�@q&B�	�a^ܝz�ɖ�MP�p��Fſ]"B�	W@���$�8� Ȍ�'�
B�	�}4f��P�"mƬp���$B�)� �9���,<�d� jw�:�"O� ��!D�J^l�H5��1h"<Rb"O̰rb��[mP-�)�ZY��R�"OI����R\��g]$p`����"O�ݠ��W�}�&�Y\L�b@"O��Z�.f�xd@�K�b?0���"OlYa�G"&��q��E�s�HH�p"O�eʒ-X��AyGhZ���\"O���B'��jg�p&<�x�E"Ov�{��;0xĂ���N���Z�"O��r�T�ұ�fQ?��U�s"O��Z����n>� �ĕ:N��)�#"O��c��i\p��*ӵJ�8�"O�M�/��Q^p0ؐ�4^�����"O���R,�P����%/�Z �"O��[�BQ�OXP�6�TX~��V"O�,��(1�@8�%V�-��"O� �C��D8��Ӄ
����"Od��K��)Ex��J� ���b"On�IƉݖ&��Ir� ��&\�"O���&	�	�A�@5x�d%pv"Ol���̹fZ̨�́=~���B�"Ox��m�<9�aJ�-�0��"O���gߩ��4�E(t��*6"O��q�J�:%����ș(m,�Q�"O�aR�
=.���C'�i�����"O��s����-}���e�ә���t*O�(:�#
���(G�A>mi���'$l�{!�� 6䬩�f�]�u�t��'��ԋ�+L<��h�e]/?�D%X�'�^�ig�A�S�����A!]�L
�'I��ڳn�Xvt���
Z�Ex�'��Yx���')"��FJЋ��A��'�>Њe��FQ�%� 튕�j|y
�'��E{���)4�&Ř�Xi	�'��̱v*A�`¦��P�U����'	��A���G��	��e׈6���X�'�t8�$N�%|����I�&r}^i��'HL�Ħ�G�"1pcL�|����'��Z��  Vd7L��"x���'<��  �qX��!�B!|���'�@9aX�g5�jIڨF�I�'´D0�\<X!����7aF	�'�%фڃ)���if
))����'��Q���S�y@尵�M�U�\4��'3�9a ��,��	rc�A�`��'^��%'�)�<�Ѩ��>0Fa�'ؘh���O	�*Iڱ`�74&�
�'������fLq��� 8ja��'{�u@g�^p�)�g_�&����'d���3K��5*���G��&�t��'y0`x�'��H���F+�6h�%��'3��g\�tb��*�r�T���'xUYa�	�]�pz�k� �B�'O |��&$Hx��y����'�&L�t � �Y�0~oZP��'��\�"ؽH�5z�Uv]�8��'Of��F�9��A^0_��
�'�˧KN'���e�CB6݊�'0�����7K���C��K���*�'�����V����d昶9d.1��'	�P2��?�@��O�N�8���'�0c��9e�8A��琰;<$M
�'l�:��&(���iܢZ�F]���� ��'�8>�~��㋁	�ṉ����|R��SF	|>�"?ieCέTĖ���Ƭa�a���Llc�DN��~ROH�e��b��}J���j� �k�d�:Tn���@�ʦ%�A�UD�S�O��h��˧]]�}SGm4G&�[`��f��s
a��(��0�k��#p|�@`�����'�cp����$��T��S	�]��a��Α�ē���ˎ���#��<���i��lfp�փ�?��$+���"}*2��e�aq�K�߸ ۓbTѦ��Lv�S�O�������nW.Y��W�d��L��H[�)3a���L5fʕ넭�Bу��ժ��'�b�q������J <�����8���F%�>�ēp<m��O��	'@R5(��0|{�h����9������Ӄe���	C���~
��
&j ��riF�4=�`���<��i�&��/�fpC+O�ᓟP�@�c�U�O�0���ML9�X��T�$�s���g�S��N�8
s�s��3F�,����#��'9�������ԩ�88u���6�&<ƴ�"R��ēMy�m����D�B.D>irQ)W�8���F���d�J���"}ʡP<*������U�"���Y��Ŧ�W�|�S�O`H��᧊+�p����71��p�T[��/a�d$�'��-X�
+wSPbǋ���'����2�����_7XQF���H�Kʨ�ē7:`�����`<.��!�	w���E��Y}b�U�q5�O�>����+M�|����Q�l {��h�r�k�� �)�'J|Z�¯��Z.U@�	Z"EDt�ԇA��a���~ɲ\xt�O32��4/=�y���[�e�s��.5	T�]��y2����ǭ_	
c�4�#���yb+D:u���&\-��x�芮�y�;i�VEP�!�f��r@� �y���	��jCG�:���7 ǈ�yBK;^d���*R::���Sgԧ�y�I��VM����%-��z��@7�y"g�'U���0M�,m"�8���y�h�?��e�t�E�9�:�i�����y��	*a\H`�X�,��es@���yő�B�ၠ�,z�%�G�Y;�y2˔�43v�Y��ʗ,���@-�yr'ԻG�z��.��l4%3w�A&�y���Cl\��$	��&�X��4�y�KՑ(D�!F�U*�X��O�/�y��<<�
���I�!X(�K�ٵ�y2�ۿXlL���EA����$���ybJъ~B��Wd�&���@���y��1�M�KZ�rg^y��L��y#�^�`�y���h���;�b��yBÔ�0����2��2
��F�0�y�� P��ݱ���9���H�fN<�y��6(�0$8҃��8��4��-A$�y��u&b�Ar�L�&��Y������yR�Y
�h��l�.TxB�XR��yn�	�*��u&��Y�Z����:�yb��gxV��W@ǋT����τ�y��W�Pg:L���E�G&�q�k���y�䗓$9v� +ǫB���AC�V��y�(���Q4��(���k�yBl]}�\����� ��:`�Q*�yB�$�BqGw�� W�H�y��ͷ�~h{�d�2;����6�ɤ�y��]}w\����	�<���F��>�y�O�h�Ĥ�fgž.���f����y"�T(t@�`�߇!� ��F��yrCT:~l3��̓0 ��̞7�y"���2 ���	9;l*eHUR��yr�ԆA��x�Ƅ��I@�#O��y
� �!B�e��(r�Cg��U��1s"OxQx�l�)rM1	�@ə,6:���"O�;d��[Rb}��(�%)" ��"OK%�	=\�x��)^��P�"O<���i��X�|�2"�.Z���E"O�\ @ReaL=Q��.�(�R"Ob ����i&n
�$o
��c"O�D�@�ɥ$+�	��ˁN�<�C"O\9Y��ˢ:�m�2��qK`��4"On�A��/��p�a�:S�\a��"O�A��Gl��Q�E��6Uu�l
�"O*�	��Δ^2~�P#�W@q9�"OPa#�J/PșPEǉ�sB)��"O`�q3���p��@.4���p�"OZX{���16�>xʦA�� ��"O���0���.���@����>�tḀ"O�ׇْG���فO^'\*��ʆ"O��!�+�/���n%xH`�*O���pA�2"6xhx#��9Eҍ��'#����ɏ/a�b�"s癑C�&P2�'cx����~$j�� ��oaVt�
�'	P] ��N-�1��#��t�ij�'G���$�I�;�hxf�s�Q�'"(���l[��<��%$�� �D�H�'�B��teC�/�bq{[�k8�x�'
lу֜S����`��($�vJ�'��ذR�[, Y@�0��ƨk�'{h��� ��QA��E�8k�'9][�#�V�^���e���쨢�'�fm�6f"b�x��S:2ir49�'r��qg��&ipy1�Ǌ0$���&O����hم�dyZ��Íe�^��k;4��C���9�A�?�͆�L����v���a���q�X4��؆�>ΰ(�
ˤfD��F�W�v�*�ȓ!�v�PS`H�9�`5!��B� P��/2��da"x�x&���s6:P��/�!珼/vՑ�4����jG"MB*L ��1���1Fu ��cO���Ŕ�@�V�q�m�*;���ȓC}t4(���9�t�R�>8ʸ���q ��k�$�6��e�<@\B��+s�g�T.|�:���T�lڼ��ȓ<b�H&#SZ�h9��"�̈́ȓy0E���Yc�p��0���ȓ�L��NV��=�RmމNLڼ��Y�6� �MӃ�:���H��Isp��ȓ`6>��3��(vN�bR㗗B �ȓn�Vhp%�Y�S��"�)J:&,6����h���1':��*a@:s!�ȓWh�		�i��a %��\ ��}�$�{��� �����ɒ!�t���1v�ijQI˫6a�Cu.ʴF9N��S�mxt��E�lxc��wF��ȓ1���VC�"Q��편#,]��r�6HBI�k�x¢�+NS�H�ȓbf���G�#<H�����{r"͆�����R)ŏ[���$M )�` ��n��q��H�$��C�QKhp��^
�Ku(�i�����ۏwW8H���X�لe�4b�f��JM��$��T�de����*��yh�@�9|A4M�ȓj4h�ɱ��28��R��)R��VDX)S�W�.�
�w�%1�.Ԅ�S�? �TZ�� ,��d���f�^Ѩ�"O
3�πvuXyyFb���ܔ �"OD�0�M6��|ɲ��5BI��"O�q�3��0'�R�I�+~HZH��"O<$��:2K� �'CU"NΨ��t"O�ŋb�Ѥ&o�M�$���d0F"O��#�+<-h���gF$H�=�"O����:���&%��^��Q"O�p���4v���Ò|����"O.�a��X(^��� �bɵG���"O
��g�Pv�HA�A�2�h�i0"O"]���ŵUO�pF��P��m��"OlP�'`���z��?T�@١B"O�<"b!H�+�VD�alK�R�}@"O`�r�lC/\>�X��ͭG�Ҡc�"O�	 �.�Pc�YtǞr���"Ov���m�+����@�Ʀ=�H,�"O�P�W��0�:��Y3&.6�yS"O^)�q�� ��C��Y�bĈ��"O.L�g �YtP��@����ժ�"O��3 % ��9ٳ�$�� "O�̊�M�%�L��Ĕ�<�J�X�"O��IT%�/�.xC4!��|����"O:�IkY
O�R���ۦH�T@#�"O��ڄ���3mv�JDd�:t�P�)"O�p:�#ʐ(.��p��<c ���"O%�al�6h�ehsb�
�z"Oj��ȵ3D��!#�J]��#�"O��ӇԵ!]�	ՠܝU��"O�(�G�E���2�Ο< qr��P"O�J�.վF���赎�%�\�s�"O�L�S��|�X���k����"Ob���:P�:%*&�^�N��5�"O�A@$��h�h��!-�0Gwu� "O>����cX8�:-�.;n@�� "O�-�R��"D|�������r #�"O�d�s��-%
 ��v�\44�p��"Ovp&�[�"b��j�;Iv��"O��Z���B�����GxU��"OF�RŊY0 >`�4'H� �"O�H�2�@^0	���p��Z�"O�ѱ�M	+�*�RBcȟ3G>`�e"O,����O#F��\��Ϛ)i=�2"Ob�`�ǉ	�Ti#��bQ�EPE�*�S��U�,i�e�dAL7@�!�dW\!�d��A�����DX,W&&�q�#DH!�$ f�@���"F27Ƶ u�
aY!��F]ѦL��k�5B����n�Ab!�^�l����B�W�f�nM���,EU!�̧VxL ��é��Lc�jɳ[!�DHy��
����q�z�z�O�
fJ!��V; ���'�-.�l!b���1D�!��-U,"Т����|���Q!��F�K�P�J�ݞ�ҸH���!��B\���e(q�&! �'!�dJ�U����	]�R��Sv�\'!�d;j&� �#��(����/!��B8�aX�@���gk!p!!�䈡#4�"��\c8����ɦz!�dH���� c�W�"�Z�{�M��se!�d90ʜ]��� d�6��/�!��.%EdX��Ӧ1ú	 A�A!�!�D�W[���w�:�L�s�?�!��$ܒ�b2��'46�xP�ح%�!�� @����͵j��EB�	=�Xi�"OX� �ѻ3�ڔ#є_�=x�"Oh�
�>��[�(P�Y�|Hq"O����X� ��}��fȻ>x�F"O
)ʓ�G@.@�Ҕ%�=�m��"OL�תw�t�Z��F�
�I�/g�!�͠c
����D#b@a�(�7~3!��t-�]�VAV�䌼��glK!򤄳MSHP�m �A�l�t��A@!�Ą�2���h��Ù[������I+9!��b��Z1$Ѱg���ا��%!�4Q�D�I�Ƃ�s����T��30!�%a���x/لѪE��h�!���rP��1�ϵi�j�X��:b�!�dY�8���L���*K�;]n��'=�$�%��U\��
�n��j8|y�',�0z%�O�X��6�D�P� ��'f�)yqş0 �" �5�H��:
�'\؛P�"�X2��>�|�'��q{#��H�)eDӔd%�y�])�I��ŤP~���y⅏*$-���&Q��P[UC��y���@4d���F� l�A����yR�σK�ҙzV�/)�jDHR�y_�C��q�C܏,�j�ڦ�A��y�#��Z�p�p'�<9P4�R�$�yr"��j��1�6<�̨���ybJ�?n}�h[�X==��i��L��y,�/+��G�H�A��4b�͏��yr	D�9���Ԏq��	�`X�<�8�Qa�Ræ���ɦ)h�trD,L8�?i���?��4��I�F�7���C��?E냌�"�!x�n��b(��C����	pƭ|.�u��Z�G㋀V��(��NR�Q��ɨ�/�A@t��͌��duRF���\�l��F�a�d��Ѭ��g��)��ǝ<���S��Ե/Ap�h��*Z��o��y�'�P������C��9d� �i��}�v��O�$d52�'�j�'��H���pU:���&�e�Ƅ�{b�h��Tl�T�I�?���Ʀ����Ow�8s3�Y�v];2�J��?�&%�?n����?��?����~���O7���R�d��ъ�
��	�Iy����%��H��TY��@-
t���S�l-���-b��O8X����WX�Qb���h��q�Fޜ<�t3��-�&p)uo�i�.O�=�݈�r
6�I���'c
�qp�f��MKq����p��4V"���&�tS��T�hn�kG�Z']��%�Y��<���|Zԥڡ�*'�ӳ[�>$bF��Es�7-6�d��q�SHy��R�H�7-kӚ܁GH�}E\l@��W+<6�s�	͟���vƒڟ����h(�MY��S@@N�4���jC+,��1�(�4E'rt��Ƃ�6�2�2S�P;j�l�Fy�*�3w ����`��&���)�KJ/&� ��a��:gZ8y�%�nt"�*�.�^7m ��:W��d�צe�q �}��!��H'��u�0Ƅi� ���_y��'!r�'j���p�IΦq�`ށd4��%�Z�`uX��x2��l�T��'ė:Lfh݉�^-jS��l�+�M�J9�Vc��x6-�O��D�O����[;�,�ĭE�wp6@:ӧӠ:��pc#�ON�D�O�(S(�o��2T��4r�6���% �uw��; `$�$땿t��x -,��'}��BɐX`� �RF�,e���Hh�����-�QQ؈
&J�6��4Ix��i8gC�V���%���d�O$>�O(^��GB_P�)�ƇNۚ�ℂ!����b>)$��h�����TkL�Ni���$\O6)mڤ�M��O4�R�#Ϟs�A���u��k�O��Y�y�4�?���?�'�����?9��M��	3#�m!Cl��-��	��]�,�0!1���Ft��H�j��ͺ�.� "���?���=�Ns ��	��-!��<}v��0#+ډb�a�sn�r����;��Y��0�S��y��!�L4M+"g���$N%7�0��Ѧ���4�?�e�-�g}b�Ⱦ�HQZr�_����.S*&��$�O��d�Ws`��F��!B,J�O��qOYnZ	�M�K>��ƙ����48`v�3�Ȝ+#P}X�7K�Ё��'��EQ�3$��' ��'=@��˟��Iئ��a�-4���h�#Ε��x[���;*
2ess�O
��C,�?�Q�^6����?a��.(UjBB�[8��sR�,%�4Xir�ҼAW<���R�&|�;6?T  7�ݕ=�)'*�\}� P�t�jP10O�gA�!H�(�%m�C�I�Oh5mZ.�MS����$�O(O���\75�`���cVPY G�IAX��U>����E�����K6nL>:ě��|�B_�|��$�|B@�ؼ�S�[ :  �^=�'8,�@D�8dM��Z}�����'q�lu��-XgF]��$�e�j�'��)�,_�X67/3c��}��'̄U�ځO��� �H���'kh��+���f�����
�''~�Yu�X.U:���:7�R�"	�'v6(	 b�$X	�B�6^�4��'�z$�D���:�x�a)/@���'��}�W���.q�g˚# ?���'�p�9J��Hk����>x(*�'��˳��	�X�������D���'A�4S�@��I~"�[�JD�f3���'#�����mB�%AQ���V �h�
�'$
�"!��e����ԕ>\�8�	�'!&hD��y����Ǭ6(t!�
�'�zpç	�.Y��h�Y���	�'>p����LF���d	�P^��
�'��<����6?���s�*S�6-��'A��)%���>͘����Ck
ĸ�'�f��2���q�2��$7>\,A�'�q)�º �$\B�$_�.}(�'�4a�Ĥ^��a����aמ��
�'P�;`GG�|<d+�J�LQ\�`
�''p9���A���2D^9N[����'Z`X G�!y��RꇟSȨ��
�'�\|򑤍�gPN!Z!��)Č�R�<�Rg��MѼ�t�O'=r�t�%_F�<!���[(�����-{ӈ|�-�[�<ǎN�o�z�21��&E�Jd�AY�<9���"�*  @Ϧ#��yQ%��Q�<)*��*C�Қy�R�(&N�<y�F	�C$�[#��K
:!B�@r�<�D ��u((�ǂ���Б,Sd�<QR20�
� �޷F��%�]�<Y�_c�&\��Ň7Bt`�bM\�<yRND�ds��'g�T�٧�Fp�<��W,4������#�\�`l�<���<%L�,�4ꂝtO2H9���g�<� �J���r�+T L
�@�Ĩ�J�<��>�\h���1M�YցOF�<�G˻8r�����B�H�T�X���D�<T*��x�-���ؕO�(�p���C�<�B�]�}@4D���Ω�j�&K�<��G�3� &h:f��*�H�<�)qg�H`¥,NH�WK�@�<)f@J�9Y��#T�(����)~�<Y��	q@�И3@�st^����w�<��%�K�(��s ^��,�狝I�<y4�I�*Tj�Tm�!z�h1���SC�<� ��NP;s*�My�G4V5��"O�-ipգzQv��m��]*�q��"O$���-+���ܴG{��g"O�i;��$z�~�����Zfν�"O�a�ɳU**�h�!�+ĎY�""OĔ�b�4*�hc@��(��X�"O,�BR�M�r�1 ��'��Q�"O�`���	.CS�ܸōə"	�`{�"O"e��$W��P=1�I�"O��zj��lx1V!�@���S�"O�ɣ�8N�ƕ�境�?�
@"O��߯uD���Y�q�h)y"O(�w��-rT�Y >n�F�x"OH�kb��niؑcY�e؎�A"O�̑#� z)P�3�����"O.��7MY3K�u�s���T�0$"O�闢��hyI�U`J��&"O��%A�%m��H��M/�<D��"OXE�!m�s�t������*��b"O0h�0
�)5�nLZ� �����"Olxc�F�-v��X{�� e{r|J%"O�c��,Oja ����ʁ"O"�j^ fW�p���>gT5.�y��.{�zY1�Fۋ[�V ��ƍ�y�e��kv��J�� FR�]3��'�y�+I7�b(���'
������y �O\9b����fh��G��y2`�#W7vL	���O)U��0
�'�� ���6a����
!% �@
ӓ�?�4K�,�D6�o�j%Q�("�H����]@0��e��ޟ@�	۟�������I�����JJ&C[j��v/�U$�|����0Y�L��k�[�8� (LI۠�"p��)^Ҫ�<a�,i=4��q~�����ɕ�1�>�J�J��M��шx��a����-Ϙ�<�ҌI����ڴx��:c@%n��b6�X�e�:�P^���?����'ډOL�YB�h�X� е��7L������>�R��I��E� "�Y���H-C�)*��i�|�lYy2L�}|�6�O8��|2m�29��wA�S�P��Z����@���?9��L��"ύU.�eg�c��P)��֝�KĴ\�G�:W�hADJM�b� �%��	�nB�g����ђ#�{Y����[�d���Z1�D|���Mι��,tU �O��s��'���+�I�~j��!��`������؇$�`㟠�)��<!�4/�§�%4���`G=^�ʡ�'ʑ���ܴu���'���r��pL�'��M.�K6 �+ 
E�$%z���d�O���矐`���O��d�OX6��0tp�A8t\�a
"`�O�\�N�jew;��R��6��c��i�>��(� ��_:�y箄,R�ڜa�Ƒ&$�v�RglܔL��\#4o���"!�Z2u����.ʶ�U4��W�N��O��]4g�9��X?���٥*�EK��oZ����<A�(��?��9�x8�*4.`��ȀK��ʙ����<�b�>R�8cV�y#I3!���� �Qܓj�F-wӼ�O��i��,7�_�L����*&Y!Մ�#M����9h��be�՟��	ןh�	-�u��'�ҳi�:�`Od���
2�V8�C"(�����/��a^p #Aȋ(�ĵ�Q��;��,a����-�5�o&htꙡ@�ڢz0V�H�h��"��0b�;��b�����'<�E�v
ͅ|7������ �hA��4*�N��I-�M��^��Ty�� p�N�dƺ|�a��I�,�<���|2�,��Q�
������LW�5��'�>s��6�1���1��Gy��K��7-yӞi4���������T�Y��l�Iȟ��d�[��T��ޟ���`�צ͊E�;,���(�Ș�g��,��F��Y&dr�\��em�
�lGy��F�!���i4�̉b��%�M�uU�]i�a�)D�����^z�>�-�B ���i �O�d���'��6�W�O�j�Fʋ|�(Pc�� \;V�qwm�O���?���?�*Ob���Ox6�u�J�Z��P[.�`��=�`<��<�S���v���"�.L)��1a�p��\o<{ٴ� xиim��'�r�OM����)�t�KV,�%W�"�0C�£G���'�2J����jv��4�2%-@�m��I9 ��p�뎟q{����A4q�6�`�A�R��O><�C0n01p�aחA�,y�C�A�=Q�)��'0=�] ���C�d�˄�9`(�>��B��LS�4sh���'��O2��z�gI0D$�`ǭž��Z#�O`�O���<Q'���dM(�cݭr��UPRaq����4I̛�Q�d���	�l�!ӣ��BG­?�6���C����	Q�	C�����^   RT?���Q=ã�R�ds���D�?9����S��?��&W$q�t(�q��8HƁ��l�}8�(�شPx��i���AV�M3T��d�rN�0$���I������П $��>a A�=   �Rw�'{�6mV����IUy��'���'@�v��IIrlp��Ǳ�D�c��S�~b�'1��'�ayr+X9+Cv �D��5Ȳa�e[�Y���o�˟��ܴ�?Ag�i��$[>����O0�M�4wT�@D����� ^`�Er'�'i��'0�ɉ��'o��'�Ur%���yV���J�[\]s�a��y|�E��&���@¶�Q�h�A��`�?�(O�}B�����������?e��ȑ��˄"�!���q�N%Z���;H>�!��9�(OΙ���'#J7��m@L�iT+E#��q���?9+O2�d�O�O�O�\��g�8|<���U�G��S�'��L
ѮQi�]��ȋ��t��	�lZ\��u��'��'@�6�^ T  ��m����#�F��˜D���w���;�'�2�';�����!%�R�'���'�ϻC�d�"�'��h')�3�W](@Z�JҺ
�a %�<D���y��'�Da�,~y"ӫ}������}�1`�AR�=ʅ��+����W��xN�O|��I�g,�o󶈁�BM�|T��c��������Ɗm�\�d
�x�\��ɔ��gy2�'ޛ�H��$yAŋ�i�1��$�q�vB�I�	h0�5�S;uL�: 
 p|���/�M��i�'��jw�O��':��A$��/��A�O������c.$� ��D   ��@��@�㐎@x�(���F�d�OL�Yxa���?��M
���ۖ��:o���)��E�� x�`�-]��U�MB|i���B�H`�]�����W0��l���}�1f�i��7m�O
 ��G�Oq��I��Y1��}�`S��Ci������?������b�O�5ۂ�̠r�<Q�O,�mZ-�M�N>Qp�ߖ���O��KR�ј-��5Y��ӳen�AG�O����O�"B   �ğ<m�c�;�h	�K�.8��X
f�*I���?)�T�Zl(\������Xj@���b���aӞ�m�ӟ��4^\E.�Mk��?���ߑ�EE %���P���2HD���9t*t52���?!�E�H-��E�3�|9���.9H�X�WJT!NC�!iGeݪ_�! ��\z82��I�'+l@a4�Ѣ~p�āB¹fά3�G�v=�bc�e�xu9/F�\�Iiu��p�'z[�����x�t�D�~�����:è|�T��bAi��˄K���'Nɧ����ƀv�0sG00��xW.���p>��id07mgӬ�;��� f�����G	5�f�;R�>��?�K>y�}��� <  �T<fE����6��x1���;H����NV�R-c��n֟��O-�Y��W�O0n8�tC�c=���B�O���O^˓�?���?�-O��-EX�T��OȄ;�����p>��i��6MaӂTIэ�1~���̂$����$H��M3��C)Av��'O��'
�@����'�Fh�����	or���Ȧ�"D�2f;af r��q+^�;D�����i���O3kLG���5J�X�V���r���oЛF%+v���;�&Df~�QQ����j�ת�(�q�kL�'Z�l���gH(@*��h�:J �f���?�$�i0�7�O2#~nډ:Gr�م�׷o�  ��ː�v��������@؞��v�<A��� ��<X<.����!ʓ^f�f�i��OBe�K{�y�d��^��Y2 ��x�Б7�'���=�5��-   �!��J_w4*yb�Ւf��,�흽GϚ�SEc#��;lO>�B �  �XZ!� �I�JC�ɹF��!�HI�r"�[6�ݢc�B��"}�d@���D���Y�C�Ɏo;�hЃݤ`��,�]�;i�B�'U�l ��)?��:.y�TB�	:D���ƇǍgH8@Z�.	�$B䉡C���C��(@����7E7�B�E��D��I�#Z�a@gnT�v��B䉭x}� �⨒-Vݖ�0���?8N�C�	>�\�Y��e��"�fD&�C�I�@��Eʩ{�T�#fE+vm�C�ɡ~�X<�E��O��xPh�rdC��FBn<Z℉;E���(sاq�C�	�f%1ƃ�j�ƙsA,���C�	 N�P%˶$;�y0c.�5��B�Iw�|X�'*N�i��ɒs�ģA$fC��1�<�R�\2x�&�a$�þ-��B��4/zy����2?����B�'2ǂC�I*| 2y� �]�1q`�a��M�7�����Ol��A�M�=�E��̱q�A�4��s ��q����	؟��ɲ�u��'��'gH���
 �o\P�����gm��RP�22�)�Ā� J�}p�c��?Sd�bDR��(O�%�'�gF���ćB�p����]6V�r��y��tl� p0	a#B�5�(O�U��i�~�;Q��+��9
с7l��A����9�O<����?��iA��7�e�L��Pa�kI��y��ا� ���o��}D`��Έ\Ϡ����>AѶi`n7m�<�b�;e�f�'��i{:����H�}b!����Z��鷧�OD͐��O`�$�O8�kT�Z98�����:n} \ �w�h����A8�	��!��V5@�s���6�ΰ�/ �9�5.{�4�"��� d�4:���[���2�O�̠=s��i�T�w�!65���/�����O\����8��H(&�����H��x��៰�Iw�S�O��kr�Ɲ[v��AbM�nrZ���'��Q�''�7-Ȣ&�T�b�2�\��Bk0��To�O��mZL�Uش�?����?)��G�" ����M���Z�,A;w�/�Y�/�-�2�/C��p�3mM�e�2a�!)�+f���n��i^d�'�ue�6䵣G#W'Z/�͊q�������*��Q�hR�'����A�8�i�ь޶ �eR�-��R��t�c�	��%P�ᇦ*X�IzN��$�֦�`��~r��T��^Ʋ �(ڧW�"�	P�T����h��	,T�B��H�1F����6
����I!�M�c�i��'F�.��*���,Q��-!b�Ǳs���Ο<���0�2��˟4����X�I�s󎊪�*�8�
 ]��p��g؁�$|�VQ��hdJ˓m��Y�ܟF�):d;vȂ�Z��:%NE�����):��J!b�C��}y.�#6��隐�ΫV���J6\���D��I���x�+��I��kt�&��j-O,A��'ߜ6�9&��nʐ0�hd�v&����Zp���x�	:ʓu���Gͻ^�JL"	C0�H��Au�&��He&��S�?%�'� ����@&�x�b$�J#I�⩡T�FU�\���'q2�'UB�a��I؟H�	=�anZ�9~�ł���
7����eE�n8��� U�nj�q�/�28��IfND�'-8���b��YF =�2%�\|0����.�@��7��(?<~}aF��.j4k�lj�N�,��p�B�:U&�8G��1C���V��[�!D�MS�i�rR��	�l��Ly��iF��g$\�� \�hC@[�F����OR����/�^90�E�< �.I[vF<��|��4�?	��i׶7��O�ID���MlZ������u�wHFGsP`Fk�%5����oQ��?�� N�?9���?�GM�Py�l�L|J�/�A�X�uj���kɵ'*^!y4��=c�1Dyҩ��/�`�{��ǵ
ڥ�w,�$s���1&����;W�ہd�,�¡�cK�Fy��*�?Ip�i�7m�O���|{��6�u��k�Q!s��	����E�)�'w1̼SS��$*.�RS�Qv��@�����M���]�TJ��� �@�@9RE��D�.KT$AI>��Ǯ�?1M>K<���E "  ��PzaO�p�������ȓ8``��-��~ ��t�D}2� *D����J�s�8�O�0���)D�$�#*#dt0�3��-o�<e���%D�d{�\q��1)�,�;2�Y��k1D���G	��"`�ȵd7'���Ѕ9D�d� eۢt����w���xx���s'%D�(2G��.��I��8L4nEH�a6D��3�A�5#����%� �$"w�4D��сM�Cj�r���%ݶi��'D���P��l�>���C�!�HX@+D���b�0�bb�d�~�"�$D��(p���g4H����T `䰩��N"D�<y��,�(��M�&Eھ�j�	;D� �.	_��p��Q��l�X��8D�x�Rh2kP�Yw܍[A
�0�f8D��!��<j�R �\?��|��#D�ĸ�d�?QD�c�Y7z�f$�# "D�\�`iC�|4�(j�+�H�N�۱�#D�ЩC�!����I�ֈC5K"D���p��?=�&�k�&�b9q���>D��pT�Q*C\]�C�^4`.��c3a=D�����J8�����L�]2�`Q�&;D�X��O&{{�)ٳEݨ=J��#�E6D���q��<g�JЋ��Y�)�T1��(6D��賏F�%�v�(�/V�y�Z Sbl3D� ��E�#, ��E�TSKb9��5D�X�@D�A�dR�@�
�o)D�@�b�B�'�.Ya����{�@���%D�x!�Ā= @�ͧ>#dŨ5C"D��3V�7�.$��,�nK<)�!D��r�Q�)�.�B�kDu��p�5D�� 4r��׶6<�!q�OU2W@ }��"O<áM��5�hP�".T�3%�-z�"O���͝�&]J��w��*{ܴ�_�<�4���N��xrcȧi�JE��g�G�<���M7����	����9ATK�k�<�䦏=zJ���#/������@k�<A��P�GG�����G�>��a�{�<i�͜&s�m���x ��9��n�<)g!�}��
� �-KR8�NC�V�Gn�\߂@�C��!��B�;Q ��h� ��X֞]H�F�.cȎB�	�h��K�����=�1.�&~B�	�j����#��e�V�R�!H�	��B�	�q_8�a٫n����a��Y�DC��%6�i�O��_��-R$Ȣ72C�-lx�JpF5;���1_�C�I(������9��p��+WT��B�I,3Y�y�&�?�A箂�.B�Ɋgif�0�ɖ���Hg�%&a�C�	](�
a�U������(��C�	�%Al���)�P�� �W)'!�B䉹sj��lR��\����$#�B䉱6�4�c6F��~��X���&�C�-;��A ��?R;`�"$U�,��C�Iu�8�CeWB*8��՜IخC�	�u$ld���6%���AGJ	g�C��f�J�ZSB�'ڶAF�2h�C�I�eT,��Z�V&m�3$�
	�"C�	6�`���0p�\���O -�XC�I*{�Țk���1D#N�A�&C䉼5l8@BA�r�-���_�[C�Z����8��i�a� ��C�	����l��J-�iɵaL(V�nC�	�i),�I$�'E�*-��-ɚ fC�I
��������}C0e¯$��C�I�%԰�a��M~X���fA�]u�C�ɹz�4��'�J�G\� �g^!>�jB�I6_�D-yD�*PSB�qD���<|2B䉺Uf!���K8<��J�RE�B��5L�Z��&ު7����
�4vi�B��&c��]Qv�A�1����.��B�I�+��խW~0��P��B�I�k��Aj��Մ)�D6,Q,p!���m .�bpDʄ\&��g��7!���b�`��B9^#�h��GF�!�d���� �Ҫˬw��e�0퉪�!�ĝ�L�܃g�I(��J��!�x�j�FA{u*�y�����XB�7ib�z��#1z��C�O`C�0�ֽz%�]<$y��T"�C��: ��+��7c����*ǻW(tC�I�|2��E/q�4QwBF�E�B�	~����.KQ6f�p�B>E�,B�ɶu�6QxGA�M
�¯^)�6B�3���7�����3��B�	�I"(y����8F��֣RDB�@���ˣ1
�С��3.B䉪Ycz���ȋ]��y8��R�m< B䉥I�e���c�#BJQ���<D��80���WW��"�-
�e�d93$';D���)�0\���7HE-�&)
�E7D����Ρ&.$y ��X�JX"�3D�4�������� f֝0U�5[G�2D�4�`a�9�|ܛ�a��#������+D�� �P!���g]�i���,����@"O�d����4��� �$�����"OL@B��>�l��3�ӛN��e� "OF\����H�#C�.�
���"OJ�9diFu,a"��r����"O�ؤN�?P4~��e` l1ˆ"Ot�1��84�� �f��-���+f"O�[��ǝmd(d��g�z�z�ґ"O$�C���*�Q���^���K�<0��d,nA#W"m��ժ#I�<�%��.w�H8t@@p2��BRI�k�<�NºQ�%�e犘{���A�g�<i�
B�{�EB�O�e�h�"���e�<Y�oN�{u�D35�O/i�$�㭅k�<	F;m �]��)���E�i�<�S&3�Rdc�̡O��p�QmH{�<aGHO|6�C�qT��-Iu�<	�H }�NB����(`��t�<q@�O'C�EP�/�\�BuP�[z�<� $M�����,�q�$�}�<�qo]�G��t2efJ�h����U�	z�<I��P�<�P�2@cQs���Rt)�t�<����\T�� F�Y��2!��n�<y�儫nn0�,ʂ']�Hp�<���\M�D+k�(i�����Ej�<�5iГ�~�£ɐ��p�i�&Qi�<�V��_/��pD�yo��Qc,�\�<!�K��JG�:^R��q���W�<�����%�[ X�d�5�J�
��B䉿[~�����ɾ�T$)ň��^�jB�6�D=��$S� �Z�*p� ~g`B�;���'��4�tH	:
�0B�84b�{�a,(a�@)�"�.B�I3ngĔ���<��p+U�Q�L2.B�	�,�˕���9+&5x7aڱC�,B�I$R�E��- �PA��c�*7�C�	,, ��T��<��QE*RӨC��<[�@����_<�����)�vC�IW5<�4���+�0�ˆ�L9&C�	|��R'T!���"��ȾpQ�B�ɝ<Ф�{ ���b�~�"��1_��B��4=�N(rEe���;%	V�%��B�  ��D�@o�$P�"$�U�ޱ{��B�	�p�1(��M��)�A��
*W�C��52~*�F��,��U�����C䉤t�p��!m<l���N��nB�I��ZH���	�G )�� �jg�C�	�6$$<1'��(mTFx� 'S�eŐC�	�n��J1놭���@T�L3�C�ɳTmZ�2W�� .��- D�!x��B䉗W:�@!���%tT�h�+�&��B�	%}�xU���&$�HIVo �C�,g�@�"D�'Tl W��0D�C䉪?�*eCR��@�Z����.R�B�ɌrL]� D��|�>D�PO*V�^B䉢YO PI�G�x+ �TlD�.*RB䉨'QI�$�? ��.o(\k�"Oڑ"1��a�b�k�@B�Wy�]+�"Oi�d�kǶ���@9BCz�h""O (�L� h@	e�׹G,F���"OP9
�\�n-�R�EW%*�QH"O��	�!��S�v[g�+5&�h�"O6����]23]@����)�Q�!"O��2�D3y�>�RN�8�T��c"O� �	�FG�=;�ة�PL�@q"Oh�ɠE�!~X`��5��c"O�b�S�D�J,Ӆ?.��"O"��'EP"0`���o�|qK�"O^����  �Aq��buH3%"O�QuX�8���Se��T"OEJ�Aށf9z���ӈ(�ѱ�"OVIY5�
s�Õʈ!���"O蜙I	Nz	�Pj <�j,�E"O\c��2�Ԝ�#�&^���`�"O��E,� ���0�,,N��Ak�"O�!�N�&�h��F��7���x�"O,��Jf��a���Έ("O:@k`��4[R]0�kS3!Ɩ�x�"O�؆�ڃ&}��v��h�:Q"O �k�&�j2"��7hY�0 nY2F"O�}�D�	{(HQ�G*_�Z`@�"OF�2eŗv bdԥ�7�B�4"O�l+�'��84��{�s*ONu@�1mD)�3B��*����'�L���¾ylhC�U�:d��'4�\�1�sJ h�e��Q,��	�'���a�$�>Lc�m1�-@ LKp�3�'"�I��a��<��Dp��0,ʑ`�'Gp9�'i��p �/��e[�';�y�g+�\ zB�J����v�h)Q�* j�E�ҋ��v)t��ȓ"���(QD���|!�ǜK�8�ȓp��!�a .*p��kWBU.h��a�HEA�-3ɸ���]�Z8P���1'2]�e��ie��ZtA��Y�����{n����>p-�HX4Es�q�ȓ^�䠳��	E��eC��7%�$��/�t; k'>���`�1I��T�ȓt���҆ U�VIrGIM/D�H}��w*�:�O�1ɨ"�ʅ,z@B��ȓ�6Lp��Q-8��M+!,���u^��@�0+m�٢aRej��ȓ��;���3|"Rċ��١��|�ȓ
��$�r�ߪF�e�P����ȓZT�r���<���x�� ���ȓ,��!����&@<���FC�v��ȓ"4EPecӏq��x�2dϘ%ºԄȓ)�,�s�HZq����6dˌ ��ȓx\�ģl�,~�xd���Ry����!J�ȩHlؐH�k��W3�1�ȓ-&$�K��B����y�ʛ,m�8�ȓ�JԠ��ݖКwn�A~� ���)Y��H=��9�b#l�����;�>U�ܰ ۖi	 ���)Rҥ��y>\ u��$_!�	Y�O�
,j戆ȓ+���J��M+�81��F�Ƽ�ȓ�ֽ󆥔/pX� �NV?NtT����V���4���熷F*���ȓD\���&Ow:`��%�0^�L݆ȓS�bea��ڥ z�Q 3`�%`����ј��"�"47"���-SU�ȓcX�XK�$X��D�"#�ؑ�ȓh��m��%�|+\8�c��"9�H����C%f�PS䈗u
|d��3l	
 �
��K�N�Ȝ��i�`s��H(TB0(�G*L-�ȓ:������
%�b�J3�T�e޴�ȓ9�a�"�N�~C�U1������S�? ��Y���:6R�S7.��
^(9��"O�$��f�6�yt�ϩz�8"OR� �ź|.���D�$0j��T"O|H�,^r�:���5h���"O�aMk������µ0��=B�"O��҃���#��Q�f�& d�"O8@g�#Y:0I����v���"O����o͚4F��9"M)p,&�5"O��)RO�4�FK 1MpX�"O���\�M��0d��
��1�U"Ot�+¯у'H�)8t#
 ��i�"O2�j�/G�MPHu��Ҝ.~F���"OT��'��E�^���A�'c�h{�"Of z$� &F���#*�
u����"Ov�`��1�0�KԈ��4�٣"O>�iTm��	�~����%���"OhT��oK�afL�(�	��� ��"O���P%RT����ȊߦU�F"O��d-ۢ/��`@g��sl`�u"O�q G���Z�l�c���"O~���g�:�d�R&Ό?YZ���"O&�K�&CYA�����uAJ�b�"O���*Z�9dЙs�L�@���"O�9�`BnsZ�p�"^�J���"Ob��%�_�0j�q�EB	>D�Y8#"OZ���EO������!B�܈2�"O^�zVg�+hl���5e�N2�"Oe�w�ʲ[*��K IY'zlЋ�"Odlp$�ݨ b"ըP� �<�b6"O�$ꔯP(szL�`��.h��T"O6��C珊
̵8k�&�$��"Ol�� �5�p�(�*�!s� ��'����cM�#pt8�K���)ۼ|��'�Ej��֨�L#�����'���m�� ���b��W��f���'�� ScX8 tM��ĪH��'�\ 	!�D1�*]�ë́*xL&��'���7�l�p�1��L�]4M��'�R�1�-F�YS�d�f!۟O����'<R�Q�H�>�xX�3[�I? �Z�'����Y�
T|���
E1Qg��q�'��kw%��+}fR�AS�X����'�V`a`A̱�:x��ϷMipxP�'�&4�F� D�k�Ā} ��'�qy"�+L���b**x�&���'��٪ ��$k�ڑǜuS�Q��'df)����CaB��n�6��'x��zum�>h�JQI^7b�nQ�'@�躕�R�SֵQG�A�*�lQ��'\}yU���
j��k�Ș2W6U�ʓ0�C�ͬO����[(���:�RY�W#��%��8EY�~�Z������Z���&��q(&���(�T(��;�x�GN *|0r(B�4�2@�ȓ}��[�
3 ��SF9T�H�ȓ}����V�e L���Ҍ����=MZ�B��	Nr���5��t��C �x��)V$+�4�A)H'FՇȓr�F���+��NfI[�+�0%����Z�j�(���0P��*�^3��ȓ�p����[&oj�(��aI�g� \��&m肆H؝6���{�k&�R�ȓ_����@��D8�t�:o� ���4�`L	1���G��CK����S�? �aW���
��E�w�Ҭ��"O����x8�\�ߕ\��,�f"OD����(Pp)AH#^O�08"O)@�u�� �Ӏ��FAxl�a"O��J4�2i��*0�ݠ�4U��"Oz@���Ⱦq�h�0��u�P��"O9XԈ�1L�NT��NA�0�;f"OT��E�HZL�ɑ,�Ö!�"Ob�c$W"D����lJ�4���xF"O�Pu�B+4Y��z��$��"O	k���6\������F�u��8��"OZ��+v�$b��Scyvh�"O H(�K)uii���s;^}��"O����UA���YDح/ά<*W"O2��cR�
�4����A¨i��"O0���ϣ۰ѫ�[�H��"O���sK2-stP��ʟ"��Z�"O "�+�1�e+)��,��5�$"O��h����hɞ��ŇD�D�=�"O(x+ud����P�y��\��"O `��кO���Ǚ��\�@"O^yH���:�LezAA�j����"O��0�KK-�
��q��b-�, �"O2�����9A�s䟂}���zu"O<�XG��Q�d���A�1�(eB�"O�@K���/:���sA�v$Y��"OBC�])VE��!۽�T��"O��H`�jjܠ���`QF��"O 3����!���"m_�,I^-��"O�iZ��D�#L�@"+A�oF�5�S"O���䍛#o(�	�$ U*6M�� "OB@@��F�z�R��sH_e�t��U"O(lAï�<L-���$@��%��"O�|ȑgI�$nT2���J�õ"O�]8��L4!$����VTN�	�"O��KR��w��)�S�['L�²"O8�­Z�v� =����&x%�s"O��V-g�.ESы�!p���'��8���Q)'ä+�$�4`����'ڪ(�1�и,d�J�[4�'GFm���9k �"�S�L�Q+�'�|ly�Ʌ�y�����W3D\��'�\Bw��|B�Y�P �:���'�p!E��C��.�*��S�/�yb�^c�����)f��9"�Y��y2�ԝI�(ʆ�O���)8�W�y��_&|�Nx��ϥ���d��yR`C�ZE���W9 @�t4Cƣ�y��K�*y�`�R*�gZ��y�m�K�*��W%g=�i�e�	�y£�ty����Z�]���B�yR��a���k�� "+�}�G��y"h�3x'�*"f\�^,p����yҭMT�Ԫ��?PbB�L��y�$�D�sc�$%����8�y�b�LWt�PB��� ��# ;�yR/�5�,��w��B��`�a��y2��
�v���E@���bɥ�Py�(Ȃ&a�5�S���X\<�d�x�<)րE/-�d��\h�r 
\�:1��ȓwV8�	�J�N�P��H�0]�q��k� �c���*�!qݸه�&!��k�F�+��0N�&4�!��"�9g��i�DE�u���&�X��S�? �5�������| Ӣ/����2"O�TA�F�i�Ey7aV/9�p��"O�����;d=��϶E�\�ۅ"O��3��3��Y�t�jXT�"R"O���j���tab��6d@ ��"O��jrB�(��	#�T�Ga����"O����i�>F���+��c�橸"O�Q�0b[6���IX�>G��:�"O�DY��H�@�4H�I�p)|�I�"O��&��&�e�f�qp�%� "O�bD� :lU���"O�mKF�E C�ȍI�Fߺ&P&%�r"Oi���$Wb`�ef�')6�'"Op��ѼH���
���W����"OX�Q���'7 8��L]�g�h["O�W
@��8��Z3P�l� �|�<���-"\���/6oL��|�<�FAB�pzJ�)��W,/d~�Sck�}�<9W,C4O#j�Ru����0C��y�<��Ɵd~�D�P%ӎJ��:b�u�<)��w�R��B�HLł���g�<�U�CrV�	��J?*K�V��e�<!Cc_��1�f�(�Z!�%KL`�<i���mJ���oHS��"�h�^�<	��T3rM>$�����J,�ep���Z�<���*�%m�? ��D��O�!�B�	K8��ċ	} Z�jq J�g�2B��;D��hzrJU
a�Zԋ�˙��C�?o�U�w���}O~9�h��n�C䉶ѼE�fƔ0i+���p�+<�C�IN]���,��z�����B��B�	�B�*4���)z>$���L�G��B�	�e��a�ӄN"W��)�`�7-�B�	*�aRCƎ�L�u�5ij��B�ID�0��n^>`X\:W��%�C�:%Qf��ӄfD�#ThE��C�Ii��fH�JjzY�š�h�C�ɼ3�����Ή?)�DY�b=0 C�/����$� b�@Ѭ�)�"O�2��%MXёpDc�f�#�"Oֱaώ=98�Dy

$T�xc�"O�(��TxJC��/w|�@����y2��2k,
42��Jw��t��/�y��X%�1J�zh��[3'�!�yB�Su��%+��:�����Q�yҡ˙d�`õ���I�$��`�6�y��*z�>؋�N��Q�r88�i �yrF
�P��aȩW!O��y2�=�����v��I���y"������4��n��B�♜�y��ĳj�$�A�*;�T-R G��yB�J8�,��f�0E��ق¯Y��Py*A�VD���Z5�R%�C�Z�<�����Z���:eaG�|����L�m�<�C�*[�	jW@�-H���c%c�<�v���p:/؟XFF�Ř]�<��0H�e�AA�S�8����Ft�<灗)S�ƍ�!oG��I \XB䉐`�uX�ϵ>�^ h��,c�"B䉰X�^�+�d5C[ �8b�_}j�C�	%XA�	�h:�Y��(F-B�	'V���	զ߳5N6A-xm�C��6���蒠\X��c�χ0CB�I�Z��h�+�5�Ni����qR�C�)� �]�@��	,�q���*�8=A"OT���*��  �(�[�8�s�"O�2��	�*���PJ�*-鎥�p"O�M����*h��[c�F ;Ϫ)z�"O�����ٲ5��zW�	�v̄�J�"O6��"��:��M9��f��ّ"OĘS��!%��2�!��0�"O)���5�t,Q�E�
��9��"O��0k�%�U��	��'ξ��"O&\s�*�) �쬈��]�E$@q"a"OR����@��3B��i���a"O|�1EU%�܍a�2
HU�"O )vN�!�(� ��C����y��6*��@b
�Q�Jl���'�y��u;�mA�
V-7;8tq"$���y2/+����(�9�,#R#Q�yB F ٞ�p#�N	7�BŐ?�y�n��f��4���ђ ��h��y2nQ/(N���̆�.�����S�<!gE��0�j��\��1���o�<��
��}��z6�_<v����h�<�'[���Q*�`	�i�m��Al�<	�ƕ�nsR,I4�OFe��HMh�<YqE��N��aE�!��u��kZd�<I@��6����,�1@tj�kTa�<6�ZM�NčT�ҍ�%�c�<9dĄ<
�c�̔9�xBvECs�<���P<hlD��j	�F�6���<��p߸e�2���k��u��(U�#Vu���+��'��X:�I�62+�R�$�(]��и�'[tqp䋝0<���V*\���'+����:oΊ��
8u�@	�'46�K��.j�8-���һ%�$ӊ��?bax�� �E{WO�<Eb�`!e���x��&D��+�b�rꑱ�`ԖQ��`�ē}{����c�Fക0&��C-ԭ���y��XAC�j��P�]��c�-dH]��$ �Es�DK�
�ʸ)S��T�f��>Ɋ�����J�x���T)0���A����>�HU�B̉�H@,P�D�Kf!�DA(���9�&A	D8��g�
k!�U�s��H0��4A�]��#I�kT!������ZTB�g1��� T�2�!�dԣ�����L��0=�D�Ӊ���!�B4}�:�X���Y8�����y�!�DW&3R)��&\�$�UA�P���)�	yHj�I,s
�R����'��귃�P��t�&"�,�'�H���U�w��\��i��$u#�'�N� 6nC�8Ⱥ�c�@G��h�'A�9S��$��4���<H���
�'(|K��:E	��V�E�(����'Q��q�&4C�Hiv��<���m D�Pxf�܀Y�t9��C	0�|���*�����A�F�N�[�a�A�	&���p"O�1@ՋȂAHA�$'S�X��DQC��BX�ܐQ��b����+������'D�����
��P�we��hk�Ȓ��x�����l(�$,��@\��%�S�MG�U��	~̓#�Ju���J�p��� �%ެ�ȓ��%)6ATLF�	�+^�R8&��E{���(������4��5B+�8�yeJ�u�:x�E�O?*��P���N�y�E�=�Ҩ�Ǣ�ys���3K����?Q지 NMё� 'ܺ� �R�YQb�1�"O�$��۰-v��U�џI2؝)�"O|��+Q�e��8��0͘��ֵi�����0�b�5D /_e>T��,Ϟ9V!��#A��9#G�9]M��BG!��1U��p�Owqz�J���r(!��G8I�H�W���O[H�s�O�K!�^���(��N��c��i1�`	�!��ZF���!JX)U�qeX��!�d]�_|D�
�.�A����̬<�!�$�H$²��"Z�,����e!�d�2lM��®]�@bYK��6F!��Ȯ`r��##��F1ZY����!�$[3JJB��Ou������:�!�$3�����:��}� %/P�!��Ѥ�j�j�L&8��Y�iɌt����E�����	�eH?p�Yԃ��y��[e~I�A�B2m�z�"tLY"�yd�jV�������]��4�#���y"�x�zp� �(S6�Z4�[���{�ʢ=�|��9	�z�XՌţ6��<i0F@�<����A ��f�ޡ������`�<�х��M������U�A��X�<�a���r pg�2K�`�v.[~�<����5Z�T5�ѧ޶V*����Sy�<�ݬr��m��ˊf��|�ӂU��yRo�A� ����dy&00C�́�y����Qy A°$��5���gΓ�y��Ӳg>���f�"�LPyO��y�NSe(؊Wo�&S�8=`R�/�yb�>Br��r��LR �����y>P��HI�X�CqD�3a�T��y��Y�mj��B',S��C��M��yr�Y�t��q�����b�y acD��0<���$I %���3v]8,58�{��1C!�dV%\�|��`B��E)P�Pk&!�dW�⹢�(m����lP��!��"=s�#.�[�@�rêW�5�!�$�),�F�AEC#�pQ�$	��ux!򄞚A2�{!O�)Ĝ	S�)�32u!��Z(U�Z)sӆ�3���Thɉ8s!�ˏ
��k���a���3�!LO!�d�2H}:,A��]8p~��Pc�ٓ�!򤕾t��a*��ג^_�u��iގm�!�d ��F�st�SAA����W0l�!�_����A�*)�8��8G�!��?_�K�W?h!���"Ǳu�!�d��.Y�4 n��y�bHx�/\
GsB"Jl؟l����:蹆bɱ^��1�9lO�,1^ �'����R�_H,ppl�(�n ��'e6!�VQ#K��!�E�+��ی}b�'��1D��g��M�1��͋?3pv4;��̚�y� ܢNz`���+)����%�=�?ѧGJA����:y���M0BV�T����W�d�q��6D�T��n�*QH ��C��h�LA�#`�b=��٦a9I<�g�'�h`"�쏪94�x!�MZx��ϓ�OB��%!\�uH%�DzR	��^�m�=�0>�5HG�>ƮA(��!��HԪEt؟4�%4�xH�n&_xԈ�!�ѓ2������s���'E�Z.zX���4$-R��D5�������s��mrYz�AW�V��"Oz,x�ƕJ�,H�a��V �Aq�\��G{��I{��9�bY�j2y���N�!�$7aYH��PC�y��#*�xJ!�� 6P�W������L�~���c�"O\��B���=�R�a���X'"O*���9F�a����4-h>�(A"O��s`��N���cuN��c"OB%1/�;�&���7c?���"ON��a(t����S\0>!ka"O�pu�F~�Yۅd��W�ݩ�"O��h"���YT{�$S1:N6͠""O`�@�GI���s�J�?ۢ���"OZ�`���@0��^<\���"OZ%�g�.-�lIP@PO��9�"O"��o˭m�D��W���~ό5���'Q�O�1� ��2Sy�M�Qa@;�ى�"O�Eq�M��*��`��R�=�6�a "OhȢ�DQb�ır�7(�xb"O�=Pr�Ӓs�v��D"ۄt4��"O
d
�L�3GM`�Hv"O�����ˌ�\0���䒉#1"Ol��R�֦uV꜊`�U�^��Ѩ�"O�k�dѕQ's�팟*��P�"Oڥ9�K*>%�[G"M'p�`�"O��"	I�>Ȁ�!� l(Eb�"O�C�%Ȱd�|�f!�*C*C�"O.�['cۘm� E�rSN��"OPUx6�3�FE�E&�/R8�]2�"O��� ��-g(3��?�-pf"Of��t���]~�$v�bX�"OP���'`u��V.g{<`�"O�(귡�n6X��6`d(U�S"O�u�#LR��v|��aY�2[���"O�Y!�d\Y4F��7*U�3X����"O�`�G$�0pl1(�Iſv;@	�q"OT|�1���c+j(רˑ�J�R"Op�������@���a"O��yq���6d �!X"*	\!aa"O���"+�00�B1�%@�3!�}�1"OʡÓ���Եw�Y�4-A"O��#�ʌN�z��߿y$���"O���/(G�@�d��D�Jakb"O��#�&�;38`q�(����"O
�C��G�H����!;Lf��Q"O������+�j6A��p�����"O�9��� \E���	�/`L�e�B"O����G���b��0ae�:�"O�+��ϮW�,�c���s<\�"O�ᘔ�2&�8��V�B�s%����"O�i�@I,�SWD��_4��h""O�@2��X�w>>iҰt&8��t"O�,�(U!@-�0�&(����Y�"OXZ�\����`iFEb֪M2-�!�R�H�h��'D�!���i��z�!��� H*��V�(E�i1b����!�ěQ�HB$�_�h��He���!��l�4���ų"+��2��(!���D�Z�`E�_�mBqؤ���5�!�䃥U"9˅���
C
��n��!�M*S�rs�Gװ:3� ��H�!�$��k�\mP��ؤ<M�##�E�a~�"F!U.BaƪA�!���趭oѐn�;b!�O�G��24�N�5dԭ)�W!�D0/�ܱ��ZzlN��s�4!�ė<cw�1�n�UL���K<V�!�d�q���a��r5���
	�H�!��y�� �@#�x��)D�H{!�� �ȁ3�S*>*���OĤvz4*Q"O�M뀈����8����;~,�	3"O� #i��k���;3,T#t��:%"O&�["L	HZv�j��	o��P "O���@�
M��Iz�+۵b���R2"O�d��*�Wb�%��Xv�D�q"O��cP��Rn,���T�/k8Mq"O���畂�X<���X%��8�"O�EbR|6$9���v�څy�"O��p1!��1����+�*%�"PK�"O$}p���b���J&�: �"O"y�AX�f�������rtTM6"ON@��@,bd�2�
xoI�"O�9+w�U|����c
U4�8�"O�t��L�*F<�K`֋%L�8��"O�	��ǃ��,�U!��;� �"Od��$�۳��l���W)J�H�w"O5sRa�6�t�t�S��H��"OX1)���3 �V�0�N�>C
�D��"OX0h��%F.< �,Z2k+,�1�"O���U�ZPŶ�S�lP1h�1�"O�l#��N�v�8���2� ��&"O\l�C�D� 
p����〉"O
I��A�uP�q��I�k��X"O�A�@��6 �8'�ü=�A��I�s�I�P�,�'%mԘhӎ�`��ѱ/�q�l��wO:9+$�)E�Ԡ�Gi��hJ��c�ē�PEڑJԙx��9OQy�(j�	��� N���2"O8��i��c�E��*�K3�R�'� ��aإ(����)݄PCR�ѨD�JckGTǘ8���3Am`���
ؒT��v��=k�49ڄ�Vn-1�éչ�y��Yn�s�)PP�t��=x�"��Ŧ =V� �	u3�4�˗.ø]i�k���w )�T�Fr#>�c��3̸��'���d�$N9��رcռGP���S��>H��a�TC�̂<FS��|"El��n���y�f�i��HvL)Z�!�r����$g�F�0EC;=�!����gP��p�� �\���Kƪ񒡆���Q
	ϓ0|��x� M2%�V9�&�},Y�>Y��_�H����6	7Ϛ|c�da��Q��͞n0Lh:0�
v8DY���2v|����$4��"�\�HY� �$�tTxrmC�/�\���Œ�h��o"�$0��U�_�@ �OM�}�;N�R�F��A��鐗��� ڜa�ȓ|��9�viژ5k�f	8Ty:́gO^�h���y1��02d��%��}��!��)3K>����42Þ��@΀t+���"��yB*�(ɐPs5gE$���8�m��'�(�+፠1�&5��&ސ3G��r,C�$�4r�M��[h���O'O�0�b��B4m�����G�'���Є�ՀJ�H�ԯR�C�8p�挙
H�P����&L��q�7��^W��zE�B�k����>4��z�ŝ�Q�&�!�I8pκQ)A��P��a%�Þt7��k�VL� ��R�.��Oߠ���2�(L���	H��Y�հ'�\�A�O������Fت�ТO�!�p僝�:�6�y�-Z)��Ȩ�BY�Q1���s�B@״��R�L��}��,ه�5k�dR!�;����6l�H:��Z���Q�Gi�/� 9"[�#n�jR#ͱ\�F�Z`�Ӡt��@"�-%3���,���>Z��:���y:��_e�X
���<�<�%�P*ph�!9�"�y	[$$_�����L&����K����i:�`NE� �+�%=
TxTT���pt�@�p$J]�ߓ]+R!(Ą��	�B����I���e��DA֥�g@X��&��T�X1X D	h�$�|�r�K��H��)Õ�ƚ ;6��+q�D�SM"$�8��O�|y5j� �����7p���P��Q�֙)2H�,&�QSW�N�:qq5�ܚ'��%�Bٴv��y�NӖT��9`3M2���Q&�ԐI�D�C.<O��aV�O�pA#O�0�j�{¨�$E��0�@������P�ٹ$��EJܴ&��3�ԕwXs$�;L��AY�a|��$�'Β4_H�5Rꆤ
0�\$�<rd
�&=�`���	�z�2u�u���A�`P�`cH��k-�Z�&�3V QnX�Ҷ�H S�$�%��f>�)���i��ب�基��[�LS�$�,�y�j_lW���!kN:#�*�0���7��Ɉ��8��3�"�2�)cj_�i\� �e͸>j�u�sD��;�9���34��	4g��.g:<�&ဘUb��y�N�!Fr�͒��i
�y6OPR�癯(l,˖��Po��F�D�Bu��Ra��>'ل< ;�@@a�ȏ^�'��l�� �[u�Dz�%��;sB�SO�����׉�r�wD��!����$���:�#��d�ĤA�&`�!R��:�c�� t��%*�;d��1c�{5����]�(�Ч�)T`����,k�l�Z%@\1	sب�%F<At��V���(�(�(�AZ�KψwX�!�o�	��y�r��&1���h	ӓ{�]qC��U���iQeEE����7a��0}�iE��XLt ��q9�gYS���	�C��Ȃ��Hx��P��0�5��A��H���3�%���	�@��������r�'��,�D=���C�`N�H�?}�|9E��&�d�R�~	���T��D0P�#Z4�c#r�H�u+Y�h�P�C4&�Ol�8 /�2*(wkD�T���	�
�� �у¢q�F���D���B�9�}b�o;W[^���Zj��0͒ yl�R��$�ⵁ��$�O���Q��x��ؗ�W���;w���!��.�xRV}!�j�9w�N���m]{�����Wy�Ɔ�qi
7䖜|�`�+R%�>G��-�U'��e�4#E��U���<B�n�$w�<E�E�M?z�H*2,P=M�$hJH�]�����A& ����'�.�&_�w.����%R��U'c�(��B�9f��E'F�X#?��h����C�?:.�5JλC_44
�mA6�2e�R�e�P�+�cӲ��`ƸG�0h����<*�-��F=�U!��a�F�C$��77�q��A
%
����tMԧY�~�'J}���+I�ɒ6�T�(�&tٴ�5�����+.mm^9z#X¬�á�(	���)���2ƌ����0V�ڰ��5s�B�lY�ϲ�`3AT����'�Z�R��.Ib���#W�2�P5+�H��2�����fK":3h9`3�ղA�J�b�k�/Je�4��O��'�F����K�r���J׹z*�d8ፕ=i��؄�֟+�f����*�n����&�N�n+h\*3/��|���q7�_�m��ܫ&��&4�8�gi�>�V�i������?�K�l=�5��BТ(��(���O\������)�楀?B�z�bd[l�يG�@�G����C6���V=Q�P��>3���7�d�[e�J�"u��[sA�+'Lv�R��S�����癹i��͚���f���q�LYÅ�ʈJE H"d�Q�f<� K�-T4\:�������Gt�UA�IM�Nʤٓ��1��9�G_�y��<=I�(KPI�6s�y)G��Iź���$r���[̀���n)i��}pr�BNT^���ٛ~����_!�8L�d�şXɄ����_�l���C�MRVܭ�T��D��d�hR$���a�:.��!����>@�����C�t�Ӣk8��7�P�+2�݁g�y����r��-Լ$��-f��?�04�!8OF�kB݀������z�3��<%�h8�� �O����_"y��YE-� �0<����$n� Հc�(l<$ poCC����s�C(P;P��m���M�BH�^z]H�*�(gX�ͣU,^�,�H��e�VR�p�:E��^��Q���& �0-�k��5�cH�1O�9��>���b���`ؖi�<���� ���CǱa���[1���W������2-4d<[�OI:�č"���1�2�2f���#�.\h�	'���I�jà9td�D�-cP�e��lN7�$ �C�NX��bF�ۦ���iӪ!=l6m�\˼T���Xj�l��VLC	d�)�2 "yx-��9o�8�� &�-:�1
ϓm�!�*��"l�U��(Y�?���f�0J ��#l�m��y��9�E@< B5�r��93'][��K�`�[�x�1�z�a;����=�����B���yv@\
��S��Vȡ�͓?o���y�@N�C�2M�L�4���	�R��S����@��D-S�l���1��:Db ![�̨ ����(�)Y���z���QB�إa�
I<C'���W9;��9L���軠��Cؤ��˓�Q����N<� m��(J�4�
˓g-�Ѥ#��' tA�a��
ݰym�"�x��Rd�+#&�˦Aڵ(�D\k2IƼ.D�D��m�Q�bL7!�X�xvDC�����Ih����O���V�̒|j�\����F��l���WHj,D�͓Qz�����M�m�@����\�y7�P��&A���h�oM�T��j3�'�T����Q�������
l?�A��呿5O$�s��N�Yp�-Ǽk��7�H&r����ކ�`��VO��zb�'���G�R�D|��.�:�q��$�M��>WЬ�Բ�g�͂�"Y�޴(���yr$I�[c���)�z������ H����-l���ӓL@�B�<0�`�Hv�:F�b|�p�A�g ��{c��c��t�4	`N�DW��m � �gU��Q0g�X���׈��y�'�
#�>�
Y[
�lc�酅/tl�@�	+��
[��j1�R�SF����j,�� �wG�9��K՗qh�H�0ό��P���'P(�+3�?H4����;e񊁿bhX�o�l�sQ��ː��f�����<j9x!*����'�V�
b��%�.H(��D>��})�y�C����aab�-&�`��C7X��q
�!�F�R�������B���̥Iʈ�����YY��0�'t��Z�&[��.ܡס�����[(1c��`�	�}T��qAP.>}��j��[�<��G��ѲS�w$ΩJ�Ɂ="9��&M%总�'��3c�?z@,�9�'��|᎔K#��;2�6���$S�Ww�Ɋ��I�0
�s��S�J:�A�Z-{3� �6�\<
���4uՈ�h4	E�|Ѳ2�'ц��I��x�j���- �p@RF"��cz�l�Iƻ�<��#S0Y6��'ݲg��V?o7>K�C8�Op �%^��󰂐.r�6��ѝ|�bP�u�8؛am��eV�L�5��	 �bGʃ��t8օ�`?ZQ���9Ft��II6z�0�(�#�g�p��c@W؞�!E��p��+v����"Tste�W�ڭi���8d�Fe��-�6F[��9U���Q���ذT��Y�p-ecL7���RQʂ�>j�����,[á�d�hbl��tK�l(;��@%LUp�6��9I�4x1`�2g�p��V�h`j���'g>1Sf��KXf͸V&�B��`��|���C7�
!T����>Py豫�EĒ. 6x�⚇Ѭ��qo[���9Æ���m�'�j��u3tBپg�v�*�a��	�}a�c^�|&���6ʄ�6�D!HVc؜THb�s�`$�u��0#��f̥ �G�=���J�O�@��e)�'B���� mĳY?�1׀N^�<]j�+	-�H$��c^P���B[d�.�+B�6Dx�)�	+ '�Aq�
B?&(�I�F�Q�Ƶ�e�$��b\�An�aU霪#'�� $���@�a�x`��9�Djb`"4�܈s��Vh|��jq�d�H��A�:�d7MM/z�P�h�.�/�j��.\����G�U�%�ժ�,¼�0��Z��k3��\��T�J�xx�P�2*��	�X���2y=Jq��B�7���K�#�� �W��Y-�]{c�O=w66����3{>N��[��mAjE���	�5�d�Ƀi�hbP#?bK
�J�1�^}�![Xc2����"?�b�#����nڠ�A&�I���3K�9V�l��'Ǩ��O�!y��tP3,���(Or���SAϲT�'�2��G��H;���@)���Wp�����J��B��,�޸3O�01�.�,�B�ڡ�R,)!�%�v������rmY����v��	�疋D��N��P�N�,��	��ȵ0Δ8�$"O�1�f!V;_�\$�ы�#�R��$�1ov��5��Xh!2��:I�1�Z�O8;�տO- �����+���%
O����D�j>4%J��XU��)_�P�L�vҠ1`=���	�0=�ȕ�6Q�H����]�=�G��p8�@9��I&T�vhހ!Ǝ$b5�C�e��
R�YѪ]A�O�!�dư]����$W�~�XQ�砚�WՉ'���������(�k�yQ>���gda0��5���ؗ6D�t��AK)/T�M���:��d!T"8����4AL/��C!8c?OL��#�� � =i�K"@.Q��O&�ѓ��Y���Q��U� ܺ�@T<�jm�剘�XS�J��;7��`��NNA��#&�k��`�3�d�N���:OP��&`��*.Y���ϛ��hy�"ON��3�+β���kA�Kr�uX��dN<�Z�*��)�W�P��p&�xR��E>!�D".��+�fT�)g�5�� �d!����a!�8�R�z�$�<!���$�4�f�Г*Ţ�( 2�!���t9>�)��"l�t8��G�/!!�d�>���1G%���YrBٸw!��:*00�Α�Q� �5T~!��ޱ_J��K� [�=��=Y���-@!���:$��+r��43�
��6MM�D!�d�8����$kb�S�>h!�d�1D,v8��K��\������4�!�d��B�?�40�%��,H�pA�"OJ���F[4��WEQ�L �"O�M��O	6u�M��R��H$"O���Mޮ`gD %��'Jt�'"O*���	W������D�Qn590"Ol�rw�ͣ&���v&�%4��ه"O�	�?��<�RE�8o�8���"O@U���1I��RG��䥒"O��2&��LB���cm�a�JB4"O"l�r�3l�^��U)U'�=�"O4�*�ثe����Ȏtέ�"OJuJ�)KS|P�C�F�G<�= �"O20Q�G<W9�E�GJ�
lJMS�"O���P��K��і(�!g��'"O��y��ҺT��Ȼ���MŌ}�V"OҬ#��7(#>`�@�͂9y�"Od�S�(��|M�U�gF�&'We�!�DH0$���Eh��{X���K�5&�!�^�'��:Pn@�K�mYg�=$!�D!0d��AW
!x�F�W�A!�����V%�9;6,�P�kV!�Dف-1��2&�-2DP1+2!�d���� {�C�67���(B�pJ!�D��:�v'X�u�����͇5P!�/i;u��ІW{��p"޷3!�DO��
��!�Nub�bd�ډG'!�!:�:�z�k�S�R����Z"!�DÆgwla9媞+t��Qg��&!�dS�3�����g�^�s��1Tq!�Q�+���GԂU����%ܡ7{!�� `���� �I���Di^8p"O���ē�Tt��'��C�S"O�0�,@�V8����I��6�x!�"O���v�I�_����UJ�V΀M
p"O��"f!@�,�2q��	ٹ.�N���"OԄt�U/vc x7;5����"O�a�#�%D��1i4�־!�J�#�"O��bE��;p+6a�D�<����"O�e�AiНP7�,)����U��0y"O��v��#z�y�n���� ��"O@k�ܩ&
����X(f->��T"O�Q횏"BW0�qA��H�y���s��`�����^<�h��~y�ȓ$05[So26�jՠ�M�@�ȓR�%��n$�P,6�P1V�B��yy<p��݈�0�G�ǤM]����j=xeETcI��d_�"�h��ȓ^b.��� �\��� p��>%䥆�3���4F�;y��H���D7���ȓhF�`�E3\fy`��K5�X��Mrl�� �ې]hcɘg��Շȓ Ԏ(�',`� ����Q�`��ȓ5~�}PCJ�hX�낆YFA�ȓs������V;9qً�Ϗ�K���ȓBLLj�@?�T�k0b�$T^8�ȓl,���I�,#O��;2�JQAn��ȓ���5/ܱ&LD����R�6`>8�ȓo��u뢡�>�ı�gM�~��ȓe5T��!��<L�U���^�^AEybʕ�d7P����I�4��Q�\?��H9D��<uN!�M�A�<��k�T��Hѳ�%W���L�� H$�"~Γ,4(�s����c�p�����MvȄȓ.&:M��B��n7̩�r��)�Q�I�h+���;(TZ���N�iB�7����鐪"�����^�:j%$@�tT��"�S:Ut��%Ћc*L����{�<)֣	.2e�E��P�p�M�F�M�b<��2s߄hqP!ڕm���bF��1c�I����; ]�LB5O��SV.HaJ���BL`8AG%3YvpC�dU= g�uD���`lR�EǶvLP�0��|*qlG$1]~`cO>��A�d�0�Aɚ2j�dtR,�s�� ���&"��$å�<M)��Y�jR9Qv�zPΈ�g�:������0E���F.�j�Y��c��N4G�"�(�"=:P�>��H��jQ#�o��9� QDj ]�"Ȁ�i�B��$ad��=�J([p�K�d|j���*4��rv��4>	�ՙ ��-.�h�$�C�d߈i� �����rB˄N:*�
�͘�=���O�b`̻����A��v�&�RP�0�e�ȓ5b�tQ�,	�b��dR��;r�����1Ϝ�8�m��!ᚑs�@�4a�lil�g��H
J>�5����X�B�H;,N�j��\ax�\��?%X�` �[H��;�.Q�c�h ���B5���"7-T*��R�	G�;w0Hì�-��<1mޱ!m.59�'��K�uҠ^y��J	�U�n���!sb��vvD�4��
���{q�ްT@H	P���K��}�Qn�? �M[�'� �5��c'Dl�w��[M�x�AW���A��|Ɯ�eD��e��,b`�+��j%)��x�QB���T����3�Y�� !� 04�|h"��  ��S�B�u�6�� �!#�HB!@�? ��9���[ .!JBn����+p�I���A0� �d"�8E�q��T	lLr0��I8C�) j��kClb���U��B�\3�>��F��	s@K9\R���Ɵ$7��@d�1��c�eU:�O�ȫ��`<�����U��h��|�3V��\���?mV@}yf!R/D�3Ŋ�%]�ԛ֥�TohA$'^�
F���`��v��0j�5Cv굳Pd.|Od1`� g�Fx�v���a�@�PV. �)�4
�E�o8ԕ`�/�c�Hi��̡e�J`�c�b�D�@�.���W� �2$7��QE��/m��C��K�@�j�?2�څ����{�j��űP�z�s���
=�=�g��J�@ cE�V�4����Sj�|�p<�4�3!�����/�&HhQ�
�l�!��I/�(l0��?j�J��_	eR�@E��iC�}`���"z�
ԁ1���W�&��
�ԏ>9ԐZF���pԈdÈy���1s\����U�K���H����J��� $Lń-7��R�gT	TF��D��G�Bh��+4R����M�p|�7�
+��=��KnD��ñG@�|D���
ӓM글.g}`�1��V����V��sS^�3:�Ԭ�vn��J\�x� �;-�d�Ë͚k���%L�/8��"� d�WOG$� YS�P���Ay�O�aJ�+�$j�I��R2���PcjU%t�hu�ƮX�K� u1�'�^Mg+��o�}㔮��4���(�
�w�`�{��8mR4��ᢎ�P �"�&�W�A��BG
>qr�;Ѭ�6�D�u��ʾ���@����@�+�MsV�Yf��0B��9��_�`�a9�_ !1O�"�S�&J�5�m	6�ҡR�<IҌة3��t iW�E��W)�#Ú�BChL7�b�1$Ѫl )33��3bi�AX!h��a��0�ѱ5�KF��:[ӓ#u4����P��$�X�"�9r�~�`���?(�PK�&x�S�'}$�bM�8�ɺt�z� �<y�5�$G�=��}ڤ*�/u$9�ϓ<��m���.q,!�'�����)���y������.k��|�����'�lr���r ¤S��Y8s�գ�@�7_F.�h��� O0�͘�
���i���`�D�O��ICa@�c�H�d�A�ZҞ�@�0�Qf��L7k��,Q��pc�\���G+r?�v[�{��ݒ%��_s�)�תn~�������IvA�%��F��Gnl�x։А/' YYgD��l�!T��b�!���sH�=�ц�Di|�'^�9�&G؛v���3��L�|�fD�5>��9Wȼ;�}�qͅmC�XG~���8"G��[���4A,�)�A��vF*Qi�[�g�|ukb�D>�[w���4󅫚!{����O�,�V� l��q���o1H����3OY�Ҏ�dM�P�񢕆 ��U�&Q5Q��\+2'Yl�9��.! ,�щN��M���3D����%�� �~�Yf���dܮ&�a)�6$;Fyq5nPc.]��Z(�H�T��鞛\#X�8����)��9�&����EB�	!|�҂�+vH�-�1D��tf�0��ᝰ?1��R�d�O��x��
�5��#N�sD����]si��H��HDN<+�z1��m��Y0�U�@C�*�˒Kր^Ҩ��_7��4��*�v-�eͪ>!�<�L���kӴY_8��烄!$��`+���(q�%¸1R4
��J!��O@Ű%�����@�]0�`�a�� @ڔ�2�懚����C͔�T�O�t�|�ihv���A��̺�1�@	<��*\�A,�E~��0^X��ߛW��8���_D����L8{{�}��-�Ta�'f����#e~p�Js�@j�]><�6 A�FV�A�*�j��-Rk3��6d�@Ȇ��bq8�'�:M�#��L�B	db�i�v�ݫ֊1)"�&.R���͊l1s��ΰj�dA��Ż8E֤�v��,�΋�C�@�Ӄ��	r��=̴��J�(�7�_�q1Pt�a�'C!FŲ��G~���qף��VXAB��.N]~�Woߝp5\h[5�u����eG��u7� D��  �c�'Q�"`ң�J�Z9��M�t5IzUNC�>젌E� &�,��x���J�nXD	nK%�H���,���ɔ"�81�2�������jP\"�J�2�|ɠ���j���G!:~�`3��'�*� $�%7��#�ښi��e����)1�0�g��M4f�B��i�Z�aQ�F�C��TgIU�0��iŜ]~�I�u�d�5�J1k�D(�ά��E8�M)D`t�C)�ɩEdx#��I#��Bh�TS̸����b:�8
�`�J����3f�ZԂ�	�zV��`��$�#��Įl��A�'��;A�%�1bͰa�D��N<y%h�0I���
	W�@;%JMU�Z�,����e��6W��H@U�1J�
���jʦ������Zf�\Of~`�S�3g�ح�-ܐMcrx�3&� �Qj��'��4P�S�:�q!o�*O�;d�� �KJU�:�����@�l^bpEaQ
�'0%��"�qag_k,�ӑB4N��d��kۃs�����'��58g��<��%�3fb�X��w�b�qc�F�l�!Cf�[��<|w�ǘ5p`�V.ٱbk�=�r�r�I'��h�;��һ$xN��O[P���JQ�Z�\�ў<���ɟt�勖��!u�H��Ơ��O�ā��Òp4�2�@�_m��6�B�\�(Q�㜣.m��&ϝ`1ay�m�<I� ++���
��:�M�P"�$�8��]n��*g�-��)"@`�����H-su*�� ��#tj����$��0�E�S>C� 9j��A�J�gd�DNǦS,~4�S�O�*	�V��y�bG�<a��q�� @�a;G�nXR5f��!��b�uC"��$c�����8�O�E�b�ҭeHd4ztƟ�T6��C�RNGR��hɂ�Mc�
2z/�pB�	(U�!�M� �r�w"�&"���O�A�fl!yk�k�I�-��QB%�%VԞe���J�~d�!c��.*��m*�-xӖ���D@�@��)&>Y��B��I@*|y����G�<+%:��$B"D�m��z4�Z�'�&(b4Α$\�^�ѧ��(R�~E��!B� �'��ʄc]E��s�j�3':�0���f#�b��yB!C�-��r d���$���(,����Ю�ē,T:x�兖#X	��ڥ��#����wZX�Bc��egdc"��'�ع�'۞�#I<}��1�L:%�z���-�3�eK��6O�B!����k
�y��E���E��U�Y2���@w�B�NY��"F�w�@+�OD�pmd0�<9ǯ�sjjztIզ]!|XW�2t�RQwFǢA�Zu��U�^>`8���1���0��և}�H��Ucׂw�@�e=z��T#�M�����?
Bhf㖋K8\@�K��	uB�c@�a5t7@F
�n1�Qa�	|����wy.�D�\�Q�)��o��}C���'�:p@pL)&,@�"[0�ʌ���B��
"��� �%q��
KF8H �,Ϊ#&tcq��԰�D��Ȍ���K�"6<��S�S'8����'2���ᒥ 3��.I~�Ƽ�Ԅ�ҠXq`S�<.S"L�KE8�Y��M�0Eѡ#�0&�؀�ß�(O�1�V#�)�-��-Շ?(����|��8# ��3�^�k:,\�B��o�DU��BP::��=��̀S@���Gg�o�-�`/]o�E��yw����R�P1��.7����"�K)`w��� aD	�p��Y�,_������n��[��4
��
�/���1�w�%p��7$�4�f���d�	�'@��$E�9���a�N�#Wd�S�jL^����͜#�R	
e�ף=�\����z�'��s��6_�}����L)
ӓ.�6 ��M�0W��p�? �H���DWvȀ���݆j/�	p�ȇ+�^�@%�,�O� �d��QX�0��F99g�d��	Mz.09v�H� ��<9R�qw�,�O�N)CiP��Hy�o�1$��T��'D��[�M^
y� �;�J��@�Z�W݋I�C	��+5/ r_U(���'�Z"c!ACQR�C�_%=���	�',E�a��(�6U��Y5	���b�$�M�$�ѧHԴ=�V�ע7�3ғ'^�Q��g�qh���� 3�v��ɀ3�pQ���4;\���[�q���g\̽�E�#9����L#&1n�Ҥ�V�+�@ =d��G~�D-R��Q��J���'`X��0`A�7�y`!E��0�^��ȓR�P��S���m���Wg�䴗'ϴy
3�[
]x�OQ>}�F:/�HDzw�@����H;D�ؠ�I����)�����%끣;D�l96   N^�8���}֡�BO5D���ꈩy\XR�gV4	!����2D� J"[ "/Fи��R��p�ô,2D��Ç`ޣwBִ{�e��Z���-D�HІk�b?.�h!�M� ^����7D��8�C�7���w ]a���%�!D�`�a�Ь}:�{�fѵ��P�T$<D�Pц/�>��0� V��z'�9D��ɣ�2K��i����&T�A(5D��;���:>)�t�E��#X<�C!D��!��e�c��9V�)�-=D� G朶
�,�uҤZ�hr�'D�4���L8?� ��&��L]��ID�3D�(	�LG'8.�x*��Q0����`-D��A�ϞV��iu���^���n6D�!��ez�� ,ٗU6 �E�6D�(U����8c�Y�n��șI5D�����Ǯ^Kf���P�V[�\
g1D�#RGĀ-�pИ �c=�KCc��y���O�p�)�J�/n�B��� �y҇��L0�%
ߴa��]��!�y��#��ī5�I�c`xhf��?�y�/۔Q�Ac2�<Z��E�ѓ�y�"��W"���@����N���y�p<�@q�f�t�eƶ�yRő=G���"�*Y�M�b*���y���6v�И�琁<��t���y� ���3��óa��│,�y��1^��r(\�r��h1$bܚ�y�׼}�f9��+_ލ'�=b�!�d��\ߪT1�[�C�n��q�]>u�!�B�#~�ä%�-���3$�'C�!�đt��	VNM�j
�{��O_�!��)>�����T�||ؠ��4mr!�՞�Z� �`�:(��4  ��'\�4J�+�"�e��a2�X�'X!���'()~=P!�T��
�'��5H���0o��Y��.F ��	�'7D��N.S,�m���� |	��'�R��U@/4����Ϲ+����'�����g�: ��۾ NP�'ۢB��U2�6py�*Z�L�yC�'2�Ԫ�e]�T�\�2k�6U�$H��'����E[n��-y2�@%�|� �'�:pS�N_˜P�@�B%~�k�'��`h�nK,"�@:5kV����'��	�,�3Q�B�!Ӡ�3�2��'� �ɐ����(3C��:m�'��!��B�A�.M�B�Bp�$[�'�V��%Ƀi	ܵ�#�:o1T��
�'K0�s2F�A ��`+HS����� ���ǯ�i�]�c�"M��0�d"O`4�v�S#K���Db�$Y�<��'_ =(�c�,1 �t!ɹ1�Xi:�]h�4[#A����,�a�:�,�}�Gj+d������4��E g�'��I�7h���P��SdܧV����� |��(���Ӿh}�q��!�?N��ϒ�y�GX������|:�ڹc]Je�Q��+x'�Qy�ğ"CP��>	V�ɓ�a�T����g�/d� ��̫�?�O|%�%X0d����uj�9gI��=� �!����K�~�	�W���S�O mѧ�OyR��[ �@=L��4-����2o
x
��ħ��'I7r}Pd�+W��C7C�=%���d��EG2�z��>9�-8�ֱ��!�=�|�Q��{��ٰK]+PE�'����4���O�I�?�&J�@F�i��I =��E�`TA��@z����M�h�n�'���BtD(�B��"n����0�'M�`���8M;xOQ>-�b���ʡ���P�:�1zG��O��\:�1OQ?�UDV|2�Fn��&V#���QDf�ɏ{rF�h��R{���!;���3n�tC��٤h�k�.&��ѴH��k�qO�O���aWkD�6��(�Pm�$I�$�ē6������Άx��@�K�P�p�	֮O����J\��ӈ}�'��O7|<�5!ܿS�"Ms�MǻF�1��4�$��g�� o�ʱT�� ��mB����zF(�6�<�ɑ���(�~2���s��a2EӵA��1��I�(C���>Y6�Y%O�F��(��]9R*�	+��+2��9����>�GDsv@K<�ʟ�A��jӼpk�JZx���ĞO���`4O�`Ȱ�G)�?��j��M뮟z��g��˄�1SbDʮd���Ï$=A�H I�)S�_�H{�"~�Zw��<(CEǭnҼ(5�P��s��e~��)�8�1H>q��i�<Q�|�`H�>{�2i����R�!��D/"td�샽m�м��o�bl!��,��Ѷo\�f�
(��E�5LV!��
}: :f啻Y�p��EǤ=?!��7!�n��*��.�LP�/X�M!�$+	-�����S6�L��Q�T�I�!�D�SsZ� I�"��uQ��m�!�ę)JYJ=Xw�^�Y��l g�̟B�!�d�/x%�]z��l!A�R�P� w"O��{��ÝK��P�b�C�f��`�G"OP���NZ:RTY�\I�̬s�"O 0�C�H� ��!��:��1�"On��O�>5��dØi,�#�"O0�ìDK��hy��b�^�x�"O������W���Ϯ�`�a"O�e[���.��H��/ǀq"ObiJ�����1��hO�(�轩�"O�U@��^�8��ur���T�F`��"O��Q`��6K�fQ@�-�n��0�"Ob�D(хX(�P���v�V� �"OX4�`��%Y�@�  +H�E��*O�8�ʂ�z�f,���t��X�'��WKT�YD��S� 
����'��"�E������@�,�����'���ԍ3�b�;cG6U����x�<�(�4�68X0��W�p���*Yt�<���B�X	����������(Aq�<��-�+^��5��f��<3�+vFe�<���,��9I§��2�p����J�<��ėn��ٵ�Z����F�E�<�b7�N��SC�ޜ���U�<�&���^���*�K���32��F�<yq��e����N�4�`���M@�<9KҩwT,%��&-h�-QB�<�*�=�L�p��O|�5[!�y�<q�H?���b)=��" �l�<��M�/�j�S�bvO��r� Ee�<Yfۻ7G�p��f �2'�0�ǎf�<�C�;Cf�� G\�,@r���_�<� ��$*؞%�aw�%Fa���&"O@�X��ǣv������ YJ�p#"O����f�Yqv`��/����"O���eg�PA6��4���x)rt
�"O��:bHT�c"u@CIX���"O��bE�OKC�4�Q�
�b(C�"O0� �
�l�%h"�N[�"O�}�"�K��@���J76E�E"Olx��ȃ-z���)��i$X��"O��A���>�QRK�5AD��A"OX`�%�3_� �qJ�L4�ez�"O��Cd�,$,`'�G�
ΰ�`d"O"������V<i��
�v��"O�)c�k:�\]��!�
S��$Õ"OB�kPh�+sA���/�%z�X�"O�M[�26��!/�<b	�٣�"O���u��8<�V�X��Q�vV��6"O��"��=#ΐ�+����(��"O�W����8�1��8*Ӳ�Rbg�<i�@�u�(������1�NY��k\`�<��	π�|p`E̙n��bK�Z�<р��V�F�c�/Ǭl���8pc�|�<Y���	Z�x���[KX�Mc�<	TH��5��1�eЦP ��cl�\�<3��G2�5`��c�З@KP�<���O�Y�,i!���?hU�0R@�q�<�0�܌[|�-�H���-��OQk�<�em�F�b�٢5�􀂄g�r�<!� ]�7]�Ѐ�ō4|`�Q� ��F�<i�����W�)_u��9�ʌg�<�&a�8xs��q���V���B�kKc�<���4�;�
�����SC�<�Wk�2s�v)�f��xy���%DJ�<AR ؆K
�0�-�Ҳ���W`�<�=i%��W��H�M&ONv}��=W[�i�1��[�'�F�1�"O�<���ɍǜ�QǆF���HɄ"O�J���2e 2ŇB�$�Y�"O�(@TVH<�3�F�4(v�d"O�8��ϲe7�����KI	n�9#"Ox�A�B!{&����P̰�Y�"OD�떬��B`�~h^dye"O �����^��h�ې[�$��s"O�(��	@�:r dSn�K�*��"O0m�Q�K\�e���N�x�� �"O�5�4�K��ڤc���.2�z]�q"O,�6"�tO���K�+��)7"OR�31�ˠ7	�%�K�6r8�"O�;�B�_���]����A"OڄaD��g�ztB���$�lq4"Ofx�
��N�
qJr��2n�Xm�C"O(�Ȇl��:�W3��x�"O�P�C��xHV,��Bŉp��1�%"O�P1&NL� X��s���W��!b"O�4#H�&| dC2��=���1�"O0�hU��?V�ꠃ� �6)�ĸڗ"OE��g��~M*F�׬{�H ��"O��K�V�������̪�"O��z�(�u�4�IJ�s��0�G"O\��K� h��2�΂'�`���"O�� �O1}|�A�R�5`A�M"O��Qj %}X���:�0"O�L�W��S�R�V�4�J���"O�x�DS;f�\�Aq����P;�"O� ,q
FK��J���kЇ�j�*�"Ol}*�N?�l�҇�0����C"Or�#fE���}����&pH�"O��0M�Ŭ�����+��Q"O���n� 
8��@(^�
�,1��"O��w� �4��6�G�/�h�HF"O�hH6���f����&�%g���`"O��8��T@�*T��eX4�y�6"OEc%�(,�j�!��Yr ��"O����߆v���x&�U5bb��"O�,���Y�I��z�f[ ^>�S"O���f! �f`�!	ą�'y%XJS"Oڥ	�K6H�!��^���"Oj]�b��Y�V!�2n�t�@(��"O���g �� ͠R�D�R"O~q�'I40�|��a��s�!@�"Ojm:��-5zac�g�&]��"OP4��R-	ld2PU]f<P"O�
V��=�R��CE�:Lvʡ�p"O�eB/Y�c�)�����I�M1V"O�Ġ�Af���cC�cD��;e"O$3�F�)v����k��k1��P�"Op$�s�Y6��$�E���b1�V"Or�R��?n��tIa�D���j�"O*��g��aS�p��J�4>�,�r"O�4���R��f�ۡ���2�"O �q�J��L�1q釄_��$I�"O܅����ZX��%�_�,��HQ�"O�	3b]�
��0�ᓣR�`� "O�T[�%�-@��)�C5���w"O �c��}T���E�ZW�p�"O����)�%b��ҵ�t���"O� d�	4t4���k�m��"O$���*�9%Y޸P��ѐV̤a�"O�C��M�bb��I% �D��"O\1��c��aGv,�����Nl8q"Ol�bWÛ6c� �zP�O �B�؄"O�y����k�!q��';��u3D"O�sT��>,��2ag2}Ì�zq"O\1١"�t�^���ǁG�2t2�"O^,p֨�W6j��!2��{Q"O|� ��>)�\KL�a0-Q3"O΅ !�Z{�t#rdM!^��̢�"O��!@�ܓY� �#3O�`"O֑�5�I�q�E��4vY��"OfL0 #B(�� G�@&�y�0"OZ�����:Q�� ňG|��"Of��i:&"$��g�p���
V"O �*�	Zh�¤Ɠ�~=��c�"O�c�hM0�$@:�ȣO&����"O�Qq!ư,�r��� Чc1
�h�"O���l�/;zI�pW/KOBX`u"O�-��.IiAXq0D��0)�p0Q"OZ�-٥G���皪r$j��"Oz�yqI�D�$A`%�8*"1�"O�1@�ˋ+��y�d�
JD "OVmS+�3��HQ��R> �����"O�遤"�>V��s�GEc��I0�"ORDr�#ȢZ�eK�-�Di��J!"OH�ð��x��Ґ,� ����"O�9[ �	�u؜!B J�8�m�"O(��D�T�x�~U���,x��G"O�x�	��]�4Ts�ㅓt�@�"O�Y��+ݏq$�$�'�¿W���ۂ"O� tk���&2�Ҭ����D�8���"O>����#Jh��G�%y�>�e"O����
�:�,��$U!y�84��"O*���A�V��H��m��h���R�"O������w��� �e�:g��"O��F|e����)h@S�JYc�<�p�.P�ex@��5�!cS��H�<��m̽Ee�@�BTb�Z%�j�<�?A����*?D��Q2��Dj�<���+�xq��$>k��)7f�b�<�$�c�N��d�Ep��u£-��yB���|a:􄂝h�ȅ24C� �y�BI'1��i��֒jd�`T��(�y�'�}��ݣ��	c�*|�c�_�y��X�A�Ta�/��a�T�QcG�y"�)C�4�u��,
}�Ǩň�y�k���JS�bQ��OT��yB�;4� ��7���0i�aBد�yr�65��
$Y�s#��!1�@��y��6Ȥ�h��V1UB��0��y¦49&�����H�_���UE��yr�t6�]�T�,��*�yR���8*�xA�H�	y�H|i3CO��yRg�� !�d��Z�a)����y�2E�6}:V"�C��m+�͂��y���Ju���A��>A�h�Z���ȓ�@�e�!0!ܔY6���|��ȓw�pI�OV�8 ׯ�'����ȓ5�8	bF��p�.}�q@
�z[�Y��3Iӓ*ٓ:e�$2B��)o���P\����
�Vs��I��];n�^u�ȓGr0�� @�?�       �  !   �+  �6  �A  K  �V  �`  g  fm  �s  �y  >�  ��  Ì  �  J�  ��  ϥ  �  U�  ��  ؾ  �  ��  y�  ��  ��  *�  m�  (�  j�  V �	  O V  Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�� |d��"O
`�(�;���8���-0��1%"Oj4��ND^[��"3/9�0|H�"OB���H��*�ʞRy=a"O�味V�!X��!&F�:J�$���"O,��a
���C�Ą�M�"O,$3%o�-���p���+Ն�:1"O��ݢ1����`���y14]2��i�<�6��{_���c�H�`�fX�$Kn�<��A̼VI�xR[�)�Ć�pඤ�ȓA5��('nߡ4�� �)˩%� ���,��r�؊b#`T�eT09���ȓ!�b��g��}�8�F��-? �ȓ
K|m�ș�VṔ���2�%�ȓ"R�X�j�4JN�1�˘X�i����̹	_�jZ��1!g��zܶ��ȓgil,*�J�
j�Ne��i�J%b���f	�(U��:���G��$Y^م�~r�� S�%T"���k\�jx�ȓ|4�1�îJb��@ӵ�ݩn�V��/[`�"�v4�R�!ʎ<��M�ȓ`:��z�ؚh�J�Z��$HY:	��H��p�m�C1��!��B:��0��EnjZA V;9����J[
2���	��4'J�EA�IVW&��~�(aZ��ӹ�>� o�Y�|�ȓ�f�A�
Ο7�H��M�$�����mޠP����/���ANXo*�ȓTv�����{ ��-7�*h��I��sB�8�8���3����ȓNe*M�悡;������X�o��!�ȓ'lj�#F�m�+R&;�|��2)n�C��0S4���T:
b���:�0!��e֊��)��ͷV��,�ȓ0�&�8#���� ع�L����'��~BB8���(1�_�5C��a/���y���#x[�d���<����^��yr�53�r�뒩D�E9�8��P���<���d��89�*:P�d�0A����~�S�8Q�eI0�>q�"j�2�j�S����hO?�MA����5dF,��
�#oh!���oO�����Ũ(�a�O�baqO�<��I��U���R�"|!sk�"��B�Ħ����"l~Ջ2�=rm�PX�(�O��(�'��4�V/\�)	���'c:̑ӓ��'����Z�L�
�`��%���'�N8S��N-�*����@�,���8�S��?	�#�5*�"����j�N=��h�<�aU�C�6�@��ɣ�"�5��Y�<���$��D�QH �s�L ��[o�'�ayBH�1��Ap��-�. S��y��P4��q�[�,�XY��E	�(OZ�=�O����sbN�1������"�D���']��	�\8�����!!���Q��)��<�2�3���c�S�v�t-�j t�<�.�#F�	���Ck�	�d(�l�<Y�㊱f�h���QEhI!��b�<�V 
8���k���O^�(!��Y�<A�]�
����E�(� ��T�'ڑ?vиM[ŌΦ��4d_�S�H#<Q���?��BŪv�9�F�{QԥŎ3�E!���'�|����1X�jD��	��tH:݄�S�? fQ2D�Ϝ�,h2��P�]�nHط"O��P5�ާ�$Qz@5О�h�"O����O�0�� aA�I�z1��"O6I���SEՂ `� ��2,���S"O�x(��K!Q¥�� ����@�0"O���Ю-Aa��`��M;"O�`D�K3%|$02ݚ2ψXP��'g���[���e��챆nc!X~���!�>��ton�y6-Ζed�П>]�$��8�p�Eh�c�8�s��5M༄�ȓi����,d9���󠖸eT
��<n}�����r��ܱ�_3�B݄ȓx����ۜJ�2܉��	l�ڑ�'���D;�)�S�ETt�s��
�!~���R�N�F�Z�����I�S�ҷ��=�^5*�N�7��<��S"�ԩ0�š �T�o��a�$��{er��G�V�ֆOuF.Ѕȓj�2E�Ԩ�V����5͓Z���]?y�O.z�E���U�
���r�5R�p	��
�yb��l�x���ˀ
Dkx=�R����d��4ˑ�b?��3��}�6�*��7$�� ��7D�����o���b]��a��3D��3S � NV`��K�.�d�A�I2��hO���XJ����[	a�F(�e	�[���ȓd ��b,Ɛ�N�x!�C�P���OV�=�O��ɉ8_Ԁ�ccR���	��4��B�	)M􄩚��ס/��S�)F�M���O �	��Dx��R>�F�JÉƂekjL@�)�)%��\E�$���Q԰��"E�3�`}bC.O�y2j�C���8w�C ��H�R'�y���Ez���'�<ZA�G�d�RqW�(����'TTd�`>:0* Ě���,��'��U("l�^0��	'@�6č�
�'�P���K�`�	d�=Āq��'���xף�"u��b�Mӭd��T��{��B���bN���A�V$6ɹ�0h|4�O����`Ѵ�[��-�@u� .aL�	��I�<A��F�r�H�P�� ft(JD&�D�<���UB�bp+�;UJ|`Јj�B�I:,�.i/e�	[W���AT-���'��>��nL�4rb�9mɴ?)�Ȼ6K�z�D6�S����4` #��9@���a��n����<����D"Pxq�;bF�%1b�T�&�!��+$��|R��I�rZ䉪�^�+��O���DM/eP��b�1L�L��mF^��ȓ5�$Q�O� !)��S'* 	��	~�0;>Zy��'�5h�\���[o
�<���T>}���s���Fh� M� }�)�ӆp(ƑB��H\���R��[,�C�>X���F��Ff[̀%"��㟐��I�[���a#�e�`��� ���1VA��A$��H�hƁK�<��i���z�A&T�8x&�� �H��'�qO��O��`0C���v�l�C���,�x��'�'i�,
�&�a`�ݡg�úJ��}��~���'_1O�S�-p�Bf0Q�;b!E�EPy��=�0�x i�6�KF�TO����s�O2���K�.]J0�� ����-0�e�	e[��)�SO~b��'O�0 �"X< �q�K �y"/Q=l$�gc�HB�:����(On��$Z�d�|�� �)#'��H�����d��Q�<8s$
�|�B����@bܶ���a�A˲DȋP��ɪ/\�465��a |#��ր~��D�"�8���S�? ��)�|��鱶�݋	����'��O�h.�oŠ���"O��0"O�hgM�
q�����k^��t�H�Y�mZX�,�5QL��B�J���vqp�1D���4�Y*�u9"��9H�.`�"=�hO��,T�I���$@%��� � �x��C�	0,M������g7܌0��	s�$B��6
��h�w"�Q���c����C��i�4i���P�:@HN5B�C�I��	�5�F�QӞQ�/N>+�B�	���@�R��3��0�$�"r@v��D �����#K˚>������^�y�֤�ȓnKƅ�6E��L�87�q����U���a�O�;x]XG�Mw��L���fUS��Q1[9����Y;@B@���8�c��։ �yr��Z9(�����O�P��ӄU���3���R>�I�EVH<I� ڰr(��0wI��[d��g�aX�����M[�'m��J_h�����J�hPs�ET�yb��B�p�C"M�>9vQ��H���?0�ļ<ъ�i�v;���H52^�X�3�5T!��*rNZ�X!��Zsm�\�%� �Ob����<��S������a���(�j݊�0h�a�D�ya�O���5���n�:	y����M1P| ��'�!�1׎uz�-��v�x�Ȃ�G�@z!�R%�l3�fϰe��ipr��]	!���<{�*%��JD@a�J��x�ɼ�TI���#J�ȑ�"�Am�C�I�(ub��ʜ�Azڦ(M��jB�ɁL����
/~2h�Kb�ƂV,�B�	�C�i3��S�|�Zq1Վ�7?z�B�	T�j����hM ��?݀B䉧��I�$��"z�.�
Y+c�tB��M7�i	����ĉ#�-V�kJ�C�56c �"��$G1���c�R�l�~C䉼ìu0�l!9�pI�Aʑ�ݦC�I�AvL��Ăk�p�5J��hC�ɛD��`�ς��C�+�T�C�	'dƭd�[4t��K"/ʀy�ȓ^����
ݩ�F>:�Qe!D���a05>�2����2�#>D�4�#�Q%��H�@-	8���� D���.@��r}K.ZR~�D�!+D������XS���DY�VD���)D�L@T&R�*\��d�k�F�h��&D�pY�·;0z�bC�1j���	%D��IU/i�Dӂ��j�.`�D�0D��C-�f�|T�@��L/H�y�/D��p�%GxYs���HXE!�C(D��PuELj���$
��i?���DN1D�d�rI1(�
ַk�bI9��/D�\�EB�Rp( q�R�P���o.D� :��ӽrV���ӧP��V�1D��ħ�t��(ғLS�nl��XG�9D�8�Di�7�nQ"R!S�Dq�A�r6D�$ d�ǒC�^}r$L�6U��B.D��T�SiN�2���7G�Z��!D���2D�y��`.�SPfP���=D�Ѓ6�P�5�������2��P���5D�(�p�5 W������`�P:&�7D�x����}�Z)K��SO���C$"D��`c�&z>���$IW[�na�sF=D��qW�s��i����*^��+A�=D�̢c�ݜB�|ِ���8�����L D�� �={U�3qE�����W��0Q��"O�e��(�?�i��I��P���[�"OB��͸K�$���Ŝ|�$M�b"O�@�Q��U�ʱ��'ʂU�*�� "O]��)��݁*z5��'hr�'�"�'��'r�'4b�':�0r�k� #�i#� � # �C��'���'��'<��'���'T��'��T
W��n��8rf�Dm7
�)��'"�'b�'42�'���'r�'Q渹`hO�2��x%��c�܈j��'���'!b�'Hr�'w2�'���'�~��f/a`d����S�����3�'-r�'���'�2�'1�'��'(VHB�[ S�:ي�H5|=��'�R�'�R�'=��'���'r�'��P" !Ƥ]�ƙ�d�E/'ظ�ː�'N��'���'�2�'�R�'�"�'�2j�d'�U2rAI�	zU�'�B�'Mr�'�'"�'���'�}BD�%�R��R��[{���'��'~��'���'*2�'q��'�6��D�Ǯ6�x|:���2ZW�L2#�'b�'�"�'e��'���']��'�*�FP $�5a՗�����'P��'(b�'OR�'R�'"�'^���O�%)�>!��ƲW����?)��?)���?a��?���?����?Y�`BE"T� S�(j�0R���%�?����?y���?���?���5����']rC^�ư����ܟQ-|-�g�òhO�˓�?�-O1��I5�M+$�ͤ`߰�y��u���j�C�Z��\�'�7�=�i>�I���R�
��(��doТcC�P�sdY����ɂb��!6�;?�O���I(�D�S��DX#�3>Eڳ�ƫ�'�\��G�4e�-�L�E���7C~A��]t|7�D�T�1O��?m����B";e�T�r��C^���@���?q���yT�b>; a��x�0ef�����I��8{��Z��0��<���'+��E{�O��&I�@�7�՛ό�H���y�_�8'�p+ܴ!����<� ��J�qm֎;� f���'�F��?��yZ��K�FJ�nҜ,���D-q��)��<?9�-!޹{�QP�'- ���Q��?���$���'J[���@�����<��S��y
�3҉C�mB7 -�Y�e�<�yy��M8G��h�ڴ������nRv"�OK�}~��UB��y"�'���'�FP�k����l>E���݂����ۑ_���L�
<�$呰�5(Z�p�M�+���`c�Q�D ��#Pq��dC�� (�tE�1�;R=�%nD*�$�"���)[G�	�2��,b��tS��Ͼ2Y�dZ�'�5�����̻]���X���/~?�S��9=�@�4��x��Ȓ��4,��ɳ��#At-!�΍'ocsi�3�ವ��d��<0H�$�(�XƮR6��ԩcM�}��H�
��S����iL�4ʌ�q�N�����D�W"��t��O�a�� ����.�`ciX�>XP�vlO-tX�h�	RՓ��eӠ�$�O�$�
��'i2���I�	~��҅Ę.
�2܉�4��$��R������i��A�~L�P+bC�<V�����f|�쀳�٦��I埨���?�9K<I�U����N�bK�m�"
TL|�&�i��H�G�4�1O�X�m6�m�T ԣJ��x�Y�4�޴�?)���?�fe�%�?�����O�ɮ-N�]�&K�~��X��B��;)H!�y�j�3��O��'��D'h��(��N�:E&�h�l��id6�O`�jt��Z�����s�i���nճ�^ɉ�&�+��ԡ�(�>q��e̓�?����?�-O��pa$�*�����d��i�z��s H$K���>������$[1;����$/٪�mc'�GBq{���Oz���O���O�|��d�?�����"El�x� "G�Cr�����zӰ���O��D,���O���K�#T,��6�is��Q�D˸y6y�4fR�v�Z�:�O��d�O���<��!{��Oe�H���	e~
�"�oQ��UЦ�,�M[�����$P;l�Ohp3�U6?8.���h��n�U�ix��'Pb�'�Pa�V>U�	��X�����IJ��-^���#�́]AJ(I<Y��?�'ϖ�6�"��<�OQfD2��IiҔ9s����k�4��D_�h�H�lZ�����O���]O~�O�,��%.0�%Q����M�(OX-�s�)�S8iR���3A8:�f����X:?c�6-�����O����O��)�OX���|"�� �d��b��R�X$�4k2T�6�]S�l��y��	�O�u��b]�m����3(���K�릙��ӟ���lIcݴ�?���?���?�;?��eY�$Ri8:9�����4�o���@�'2�%h�����O&��?���5y�l �1M�=����
|Ӵ��^3u>V�n���d�	��P�Ɏ��ɴ�Dr��|��x���
~;W��3%D�ϓ�?����?9��?�+O��h�%��5%|�CdF��0Dq#�D�>WR��';�џ�':��'G�̚F�z�(�+%dfЙ�(�"-���'���'���'��[>�ȧ�
��M����R�8%H$!	� ��mU"+9�6�'��'���'��Iȟ3��q>�ҵ�V;f�D��Ǯδ&��9f���M{���?���?���?93��N���'�R���h����#<�*���S�iR6�O��$�O�ʓ�?��M�|��~e�3O'J���M@*��T˙>�M���?���?9/������'1�'�����
M(tc��\y��X�(�y�h6��O`ʓ�?y�%�|�I>��� �pt'C挘�a$*;�G�i�r�'��(�o�����O�D�l���O������ G� 	Xl,م}��'r��s�'hɧ�t�~j�H@^`��r���@^9Be����}
ĬM�M����?)���
�'�?���?ёd��37�M�	�d<�������/-���'�i>�&?]���I���@��.b�{�$�4i���4�?��?�`#�c����'4��'wr��uרZ'G4���W�B�=��!��l	���'{ �+�y�'l��'�mR�Ɠ	(=d5��P��ؽ7�l���$��~��n���۟`�I���I��X�`�^�
]\�Yr��5��Qj嫨>Y���P~��'���' ��'�����"�[&L4J@�TQ�M��IkȹPGbӆ���O��D�O�H�OJ�����D�Q��M��%ez�)���1=v��	uyr�'���'���'a|LS�"o�P���$�+�x���<X�c��Z�.6��Ol�D�OB�D�O�ʓ�?!E��|"���t��l��ƒ�J�0� "���'��'ZD�~:DΈ�a�6�'InҾM:���P ��r��j8lZ �aӶ���OZ��<��ujΧ�?��R3X��Ɉ4Xu�)�"K�8�a��`ړ�?���?���)�r	���i�R�'{��Ol4u{�#Q�|�\P��"Z^�5�BG�x���<���A�0�'�?*O�i���%�P�P��i��-@�a�4�?��ye�HC2�i}��'�b�O����'<h)���Źm��ЊIN��,أ�,�>��]M�Q����?�+O�	6�T�:@�z�[	R� L�g�0�M����H���'���'����O���'�"��9��%P���yA�58����t6M�G�p�D�OV��|�I~���l�� s �"��5[w,\�u�aQ����	ӟ�����,�1ش�?���?���?��&�����	��{ff��R��o����'�#���	�O���O�ɱ��1(��T�C��02YP�a"F����I�N��	޴�?!��?!�:���~?�D�|% ���fC�����[�6��I��8��{y��'��S	V�}Q@\j|�x�G` T	�y��D�O0�$�O�9�Ou�	��8�PK��$b����~�PL��Cd����P����T�	�,�I�������:�M�w鉂p"z�!꜐h�|xҧ����v�'*�'���'��I쟨QG�e>�)�J.&�ڐ��p��J7���Mk��?y���?	��?�0-IX⛦�'�B�R6~����1��RU�=�v��e47�O����O�ʓ�?�Љ�|�K�@Ig�"����O��]��
#Br�.���O��{�x��F���'��d�X�&״�A U�7�llR�d��I^OV�W3DDx���]�P�j�ڀ�LF�4:��i��	02
X�*ڴ�S�������؜e7�E��!�(� 6a
����\��r��$�S�'h�(��B�Dvn���Hǽw�N m�80Ҽ3۴�?���?���e�'&£GW��})�k����P���A 6̈́�b��"|"��k�Py���E�; |� 	G�K�P����i��'��X��O4�d�Ot�Iuɘ6�@|�����W�.x�b�(ɶ��O��D�O�1�'�M�~
Ԡ�`K �u�W�FѦ���2u�AL<y��?�M>��i�P�L W%��qc��8}s& �'ώ<�y"�'���'��	�%��#���)R�:3�ŉZ��	�!�ك�ē�?�������=�^	�`B�-^�ZG(�(���k��$�O��$�O$ʓ*tzH3�?�:]�a�_�L2�\ҒF�B0�%�e^�t�����&�p�'�����O*%�r-Ǔ?�����!�7v/��0�V�l��某��Yy2��z1:��\��h�#��@rm]�h�+��OҦ��IV�	_y�m;��'y���gǡo����2ʆ�CqܖĦ��I󟤖'�T��/���O����ˢ��`_0?q�a	�hF�Jh�&�l�'���3��T?%��!�	4>�b��=ri� ��ml�:� k0���i���'�?��'4K�Ɇv	V��H�@��	�ǋ�gt�6�<�0��X���Oc��xPj�.W�Ne�F��R�j�ڴyC��ӺiK��'/��O�\OT����+Np���#��H���bXv�FPm��H"<E���'�Z���@�1��Uij���#�M����?��W�L37���O��I�p_�C$LԷ"Pf�2���	O�b�T�D��ҟ����4�	ٟ���<s^����O(�l�!���:�t��ܴ�?�g��i1�O��d>��ƀ� 4��'��0y���7�>I�@S���D �� ��蟸�'X*8�D��$O�)�.�(S,��ǂ*M�.O����O��ĩ<�*O|\{@�h�t �4���H��|���Ǚhn1O����O��d�<����kd�)�3b*��Ն�F&Qq���"/H���4��˟|�'��	484��'@�RQ�1�+Fb��g-ݪ[��'�R�'�2X��� cI���'T���7�
uj�9 D�G::|p��i}��'��Ixy"����Y�L�"�ްt��C*6��l���n���D�OJʓ�\Qf���'q�$�^%���
fb�F4�l5g
Z6ͷ<�)O����?��|n�5O�Q�R���9H�p�S�I!4� 6ͩ<Y�C�WM���~2���2㔟�X�-Ì	����Ǫ$#8݈@�pӾ�2���Ex����#8������	0�������0�M{b�ܴ_֛�'h�'�t�:�D�O&�I���6˼��a�N$�\�P�¦�hCm7�S�Ob��)� p�I�@$j�v���+E�~�Ʊi�R�'BbQ$>O����O|��* 9R��ׇP%�d*�IG3dSb�X��>�Iß��Iџ�H�BK�$���0�| ��]>�M���
ż	�4�x��'�|Zc$��F�D��p�gH�Fb�8�O�i���F���'��S���ul��r��
U���R*�!b�8<	e��D�	ٟp��A�IYyʉV�
8�gCN*"��mҵ���v\�y��'�R�'7��	xE&t��O�Er�ƚ�%���w&��Nk~%�O���OܓO��}u���'M*,Uԭk���qBO�@pd���O,���O�ĭ<YP�7O�OJFUCs!�(clL`� wZ���{�.�d(���<�FN~� ��P�7gh�۱�X`��m��t�IMyR��	9j���$ퟬ�@��s��d�b�¸+cН��e�Y�IEy�'Z��O�S8?����a�fz���쎧a��7��<!�"t��I�~����w��8� L3%:T�3�#}��,H�kp�ʓ_�Ȣ<�~�P��;L\@���_��lC��ަM��Ɔ9�MC���?1���rq��Śa����go�8A;0�	q �ndo ;B#<E�d�'�d@�^i[f��*�5:Q����M���?��t2~8T��ON�	���LJ&o�3c��\��$��^�c���6��8�I�$���Z5&|��1!FN0��DW(��M��#���7�xB���ش���C�X.9�T#B��1�$kKo}�E��'��'��X��Y1`��L�����/^=Br�X��5Ye�y�L<����?�K>�)O�ÐE߸?^`br��o����+1O��$�Ox�ĥ<)W�����ID�s6p-+��؊=�XÂi\n�������	^��yy��	���B?H�is�%�#Zq������	�`��򟈔'�=�E.�>�>�e�rdM�^9V�B�l�ǟ�$���'3����}2�V�MJ"�1��*#iV1�ET�M��?Y-OA��+f�����S�M���$'�k\|�Y�j�H�}�N<�+O:��w�~r2`K2h��� ����h��4z��ئi�'* ��G�q�z��O�b�Ol�/+A��W�$( �
M�o�byR�V�O����ǂ�"�02��K�T�N|��i���y�.v�B��O��D��J�&�D��ܦ�i��IVL��b��]0��i��!2���S�dP���#
ͺ�F�W�\\�J���4�?!��?a��#"�' ��'W�B l&q�&$�+D���7b����&�֟p�	ʟ���-�1���A��GOrq[q�C��M3��L.�\����O����<��v{d�HЭ|-��+�*_���'�>��y"�'���'�'`n�U;�!Z��d�BÂ׺[����q�I��x�	u�	zy�M�(I.��BV()/�RQ��g��]P	[g�|��'vB�'���Vl��O�"��b�g�(�{d�?��	[�O��$�OܓO���O�}A�k�O�ݢGb��E��E�+kt�P"@�T}��']��'��� wu�(jM|�DO?1�;��	g��� �ҘwZ���'��'���'kd�A��'��J�B5s���T�P�e˔�I��lZ�L�Ijy�lмII��@�D��b5Cl^9XrV�+�7s;}1D�`�I���I8/G��	K�~��,�"t��E�0i�,���b�ަA�'���|Ӗ��O<b�O���#V���t0���!�Q�� l������4&�E��DĒR^��P�]�=�(x2dA͘�M��{�v�'��'.��@ �D�O���S�����ō� >:��dIަ�)��⟠%�"|j��o��|q�'5+���R Fɜ"L񋑵i�r�'呲xɴO��O��	{���qӶO�n\��2[��ݴ���0�X����'R��'���+��[�ܜT��O�"��`�Fx��ٵ|���%�$�I꟤%��X�b?xӗ��p	$��D�
/&1��|�
�[���$�O|�$�O�ʓ%%j5w��?bպ;AP�88Tm!C-�ԉ'vR�'	�'wB�'2� T � R��2��3�P0*a��=x�'��'2U���������sh�-Y��6���s �K%��$�Ov�d=��Ot��O�X	���9#+B����C�����hr��'B�'[�S������ħR��YQC�
�6��Sb�:u#2ASüi|��'
���W��>!��˞a���ӭ��j�\8 ׉Q�����p�'/PȺG/�	�O����*������U�u@��L�Y�*i'�l�Iٟ��Qޟ�&��)Z�l(eɊ)��]H����Hl�m[y�D�'	_6�[���'��tJ ?��)��Ȁ&�B�s��r&�ͦ���ҟ�Z��B�S�*Hb�H��>��	�Qi�!�xE�	:U��",�'�x��q�'�4��@�E_r�3�K���`���&� ���$%ە��$
��,)�,N��`!�P�W$��QOϟ�v8R����T���*�̌i�텦C��0�E3��KdS�%��re���@�t�ɹN�h�;S+��:kN��#$l0�,W"Q����"͟Y�hM�0F�"8"��2���0��Q;Ѓ�`s��B�O���O����º����?��O^hƮS
-�0I #�4 1t9
�bNe�杩��� �`�raEW�tZ:� 5h^B�'�8�� ԝ	1흶'�(�ÒK9���#��ݛ'� e{�(^&иB�+"5�!x2o��L�� � ��tS�JB�UY6-V�L�`�	{�'��Ox�۷����I����=xA�W"O���2X����f�b18�+�V�i�f�'��H�($Cߴ�?Q�K�4�%-R8\%q�#�5H��U����?�����?������	��N��`���5z���u�ޡ���"���.,�N^=e��E��\4h���Ey�nR�4����R�Q�$͠2�Q�"���0R)B'�Ni���-/��c������Ey�o��?���?i��nX�8[1@)k�$��G�āqGl�.O���:�)§�p�w�׵;ʺ\�rg����Gx2�i>	��4,����M*( �����^;������d��F�nz>��IC���!yH"$�j��Q"�阌MZ���/.rR��'�.uyCB�!��abu��^�ZQ�H=9���_>I�T�N�}��QY�� �je:,���9}���6�� A�ǡ{��}��i'*.ʕ��K��%����I���)Rm�=�hJS ��V��'|�	����?��)�O:԰�Ě�R�����l�x�~l1F"Oz�+��� ,�D^�~�h���'�J"=�0g�:X���H7T�*��@ؐ�6�'�r�'O&a���G<#��'����yG��	�^eɕ�L�S3^�KbMV�n���"�Yhwd�&e�����W��?��<Y�9FkX"��鰅�Ӈ^�NT�$��U�Z�!b���l,�����I-���-S.hR��ɏ[v)u"I�$�(��$?c�Dڟ�E�'2�	5*�=�)ӊL�'\�Z�'[t@L�c�� �a �R�E��O�Fz�ObQ�|����/j��1�e��	�rM�m��{���[Պ^��0�����	��u��'A�?�HS
́ �	a1HY�~O�&bA0 ����f�5�p�A$�p<��`H-S��Z����O��yva^'5o
hS&I��fX6�k��W{>��Y$-~kq	0ьx2�?6,�v�'ג6��Ѧa�?	r�i̇?�j�)�-�
6t�i��ײNV!�U.Px`Y��
@kR�Kw�P0�1O�=l�ؗ'R��J��~*�\B��R%.1?��c�@e\������?�ā?�?9���d@��(-�xsv��T*��6`W�z���a4� <)R����XM���tȟ|��xFy�,� E�)���ܜz�́�e��!�քI�Ô�n�fғ�M�
[0�jAj�~V�A��$�2h��o�x�'y$0�4�[�b�5�M�5�$2�yb�'�y"�݆WI����3ø��EG�+�x�+b��9��Sa�'(ȵi��A"���O�˓�\���i���'���t�(�I	~��P�6�y\Aj2'L�<|���	͟@��c�6?�i@�n�d����|� R�|�g�	*����z���hld��˱G�BD;�do�Oi��q�$1������*p�L�N���A��O�Um�*��'��!]N)+�LW�u��7	'���<����<Q4�T�|����S�ű{L!�D
�z���D�=wHzu�{L\�hf�)S�`�o�d�	ß�zc̘+#����I��8�����j��H�"$��Kx�l'*
t1���D����T3�y��|r.=���E��()p���AL���lҳ	e���*�C��g&^���������dB>"E��'�A:`5D�a��
S���nZ���D�+�O�����X��% V-��KQ� Q�� �!�$�Ln�M �F���TC�fV�S��I��HO4��'��I&M��L�F��vP� H�A���;��� F\`�I͟��I�� ���p��i>(f'��;�E�5��-W���ģGr��9�S$h�>p�QbP<{Xz�!��)~Q�����?P���<>tf���sp~ Ѥ͓8�h�{!G��*=x4�ʙ'M���%.�@�'f�4!U&�/��֯?V�B�,5�����9�M���i��[����L�~��PRf	�)\�;sBMK�x���X�y��F��L�i�f��.e�b� �4�?.O���Gɦ��	蟘"7F"��Y[�-V06h5������2���ß`Χ��2͉6o���6�@lQ�tm,���˃�0��%K�z���,��ȥHI�L�´0�uÃ'Xܜa�Kۺ�`��O�'7  TB&# ���O�a���'v67���IW&���D\�g��QQ0.I>2F�'�2��S�`��L��ǲ yT��>c
B��;�M�'�é�ʬ��ˀ�x֎�A5H��?�-O�i�B� �����Of˧?H����KEB�g��db�l~(Y����?�&�.~�!����.(tB�T�.6�:*���Q�R	�S�S/E�vU��C�_z��'��Yӳ�'�th1h��s
��æ�78�@��O��4�	Jh� R�u|�	J� AD�O��n��'��'p��ak�Y�$jĉ���D�N#6��<Q���<�ѭ�t�,���n\&4�~�!���j�\X�4P�֖|�
��E��ՃR�/qL.�A����C��7��OR�d�O6��`����d�OX�d�O�.A�8�T�h@'�5@)��^�$����NbXf���v�n�qU���b>7�@�=F��	�(|V1Ufs"R�
ፒ��^��@�S		�4dlbUj�R�禙#緟� ȅ�".I���AB�� v��BȦ��ݴ�?q"�7�?�}�'�RkP�~�q� 6�@ �������!��@�HĴ?3 �a&D+��O��Dz��OBZ��cR��-K��l�oEM�X�IT,T�|a\�Jǟ��	֟��I��u�'k�3�TUx,�+�ڍ[Q�N88�U�c��|�<�K��Y�#$$��FЮ&��d�Σ�(OH�3`��_�^e�uLU�c���1�C�v�=����h���;f� <*�yf��h�����Iq����	Ć�D��3iN�H�$�����럼�	��ڟ���l���*H�P�"䇶I��P����0>�H>a�jR�mc��YqdF�[5��)I�1O��l�ݟ�$�p�H|z��� ���
`K��)ʔ	Уq�<1��E3>�z�B���s�.��C�C�<1� K�	��;2C*m�	R�C�<لG�,����%�̓���(S�<V)�5�8������7[ڥI��Xu�<	vOR�~(͋�nL7#a$eA��Ji�<����>�,�PbZ�gM��A2��h�<	!W�9���B��k�T�q'��M�<I�Y5�P-7�����(dh
M�<��%̄hzV}+�� #�<�H��I�<!����O���!�� 1�0�0��YK�<g)��_�"��C�$�B�{�#	L�<�T@\�F��	vίQ�Z�JPOL�<�p/\q铅ת}5���D��M�<1�JS�5��:���|�m��@S�<aT�qF���%A�U⸩���W�<��Ѣ ΰx�d^�`<�Ly��W�<�w��r%���ln�s�h�O�<��AO�`!ʶF
�r�����Nd�<Ѧ%�<6 �&n�?iltq�EEb�<���֮-9�$CZ�&�!) o z�<	�F	#H�4bd,!t�ļ�Q� s�<Y���8@����Ϸm�X� �	H�<�DLV�� �C��(r&$8�n�Y�<���Q/\���S-�(`�
��p��W�<�ƄЖ@����]�C�!(��\�<I�D:&�l��Vd��-CW�\R�<�BҒi��9�"�U`�j�R�<9��D� S�!Y%i�kV��V�J�<�R��#ee�t�DW�.(�l�B�<���`IS�f^0�����	�\��C�-{����	�B�`��IH�6(t�K����p4��V�Xb>�������&m0%9b�Uv`�(��C:	hc�C�cfXD3e�O�����U�L��N�7�a���H,6�|�+"bC%$!{���}���`�ć�b�6�'��O��x�8�(��X�(RM���48�V}q�>�@��?)�v���W�IQJ��=):0�A�"\�c4�	�Y�0Yۗ�|2��m0X��GMF���U�[�L5��b�#qT6����;n=\4���D#=��<C��6����
�y��~���a'b��h�����šO�Ph�H86��˓W>�|��?�"5f!�V��	H�ܐ�!0��$j��h
p`8 ՚�dJ�3� O�I�jT�q� A��f�Kώ�#�i�B��0FH{܍�<�O�.<92���$k���N@wm�RZ!3b۰!�LK�� 4W�I$�S���=�O�^�ɖ.*G�4а�!F�TI��'�`�G�o(���6� e�����&
	`|��sS��b2�Hit�9m频�<ip����ɉ�@�|4Iw�E�	��i����3;�	��W�4^Ś$�'�̜۝w��A�1&H `xr�YE��.<c4��PC	\�J>���o����D%(��0��C��|�N]�g����'t����Z*\���c4ɗ
?yМ�H�`yb̃3e|��1�g��Z�
�?��D	?8��[�yʟ�W�x����̈A�.�ӡ��`_*��Z N.9��]j�M�B��D��T>]p�'!J�Q��&_�$��J�%Aĕ�L�H2V˅�)!T�=�����#$�ɉp�)���%ZV�qP�
\�V�Z�yR�*HVם%��>�rcD�n��"��BIt�q�d�wF@5��ŀR�(uGzZw�(��ȼ���i�%iV�_8�XT+��%l����A�E��I� .�,D	�W�VU��O�<Qр#J��L,�C��dhX��}"	�$ZV 8�@M�h�^�0���F�H�g��j�#K	�
�8�( $ܺV��M�-�$Tc����ק�	���'��5�oD�Fw�]���11��i�zF�ip��-���9K�\��y�c\�&���|��8�� `б�X�K�a��ᖸ}~�豟>����1����k,z� ��i�P��A�	�6僘0�r��ЩG��UZ��I���O
]�֡k���ĥS�$k�U�;��)A�/F�*�:0��-����žX᪣<��M�w��O�}
M�c7\�s�-R��� �̗4t�{��#O��I澥ˤϣf�O��'O�Nr1K�ƞ�_78bu����'X�asϏ�|Y:@��+��2#d^��eC�OT�IpF�K��Y���
;�����'���"Z�U*�&���٫d��d��%:ê�.���`�u�v5�r�@�M,
� �Z=A�`OH����F��t9�U�fc>�@%"f�r�saH��7Ϯ�
d-%}�ʀ4	��I�XH�e@�E.��'�x�: m�)��5��&�)�B�jÀ��'�f �@>O�͓ ̛�u��0��4i�½+A���CV~ᣒ�L(X�ITŠ��(3�4<�r���+z	ʣ<���V�Sb��O*�h��J�`�R��1�J���ݸ�R�r>�K�&��8{�I�
i�L�P&��pnɧ�E���UN�`uj_;a�������e�t=�`�t��&�V�d̙%�U��o_���Y��t����T� -�lc�B ]�{���Ka�R�|n�$�����B��|IǈP��H]���I2Q6H�0�ݷ44�e�'nP�,[H]
�4OH\�O� �Sb�Bl�CsvެA?���'f�[7*�OV�GI�m�t)��2e�K����^�c��h�l�	9�63��3.�r���X��������'1-q�c�&�z��$
łNܶ��� �A�t�x!�'"P-��e˙)�a|b �au8������i��T5!�`�RЋ
�(���r\�3 놢�H�@�ĵ#F���c��?e�D`Ƈ
�R5sb)�7A�\�p�:�IW�d�@h֧J1R4qd%�!
�]�v�b��Wk�+*�!ŞVc�bCN)�#^�ZUI�-I����� ;2���m���D;G!�L��I�[� #Ĉ1z̄�q��$_Ĉ·�3���pm�'�~h`$Ảk(�y�$�9��Xh)O���⥂$(��!�f��_�Hw�I�N[��2��ןtM�*���Ct�	%n��E|BMV���)����A��΋S��cQ�K�bXj`F}���:�wε�	��gP�cD���� �T+ڰ��s�'���h!�	h.6��gk_G�,��A2�؁&@�RP\m�_s;"9��l���D��)��@#����ah��v)�2�џ���̯"rJ���c˅KpyP%a��Y9��8IK!U���F�ˈ!:I��ˏ�3�P�N�,����ˁd�ࢄ	�]v�䧌�G�:�+ы�<�uH��r^���Tz��)cFme�'nn��h�"�fd���.C�����x���m�5""�hz08G/�.[yN���`Ab�P�F}���3t谙w�E9(ŖmfYPU �0������hO>離 �	7��S�*�yn�`���?7���Gx��;��H��E
kr0�Jŀ����D
�HઽC�H��~>%K��SY�IC�0Uޠk$AD_
�$��C��l҈D ��ӿ^���t���hF��d�<�����)��X�d�&!��IB�"�� ��ۧL�,�Qw`P#+�2�s���<��O͡���0�ўN��x��!�M�'1B$��&Ѿ T���Z8S�̌�+T�I�qO�P���T?}0�iO5{���$�ъy|��+�'s�Ua�oO��>���r�����ߗ1�h�`�an!(�i]����$C��g��?1`�J�{��A��5V��H1�1LO�!rĂ
����'�DH�#])J�L���72��T�J�4 �Ҕ�@�o�)�矰��&R��`D+&Ə7{Vѣ�-�ɯw�Vӧ��i�e��١�ڣ5��]���P�z��	��8,��'l�b���6&�fh� T4S0�CɆVI�O�a��	D��[����F�'a�h9R'u�C��D� D��eh���í
o�I5B�)$^a�T�OnTz�U>ӧ�i��'����7#�1�>)�p%|������	*��<#���Y��(��A���	JKވ�g+&G�x(Q�����)0�,{'��4�LA�"�~qF�b�J�)���)��1)��Q�z��T�T�b��p���[�1�G�%�O��~b0f&W�i���"�C�S�}�'�L�ǛN�N� ����XL��ˉ�$��-
.� �Y�XP�$��b�ڦ��0�S��nHμ�s�J����d`P�]3KoV���W/�>Y�^&Fe�4ͻ6D�+���@K�ذ� �vV�0�IX������$*�
j��ҩA?.q��IW�3e�"<iu��K�*��7��~]�D��N~r�߁��X�%� 2�<m�����OBg��* ș�n����s(@���3N�3ݨ]#�O�@7l�p�_�xc�A8ׅ�B{�Xp�6O6��QJ�jjp�vÇ>,��BvS�����-_z�	� ɭ,t��b	5ʓL�"���W�HT�PUY�0$D���!h<)WE��`��Y�T�� ���A0�L�2ՄY	��%�x�>1���8DC�E�;0�V��7J9T8���H�2��a��	pmV�3���KDh1!��_B�j�	P)YL�'�*$�e���a��`FFU�h���O�$���Ev�rҫ�>�$�(P��?�l�A�Y���u�ЪP�eI&8��C�	6l�ۥ�ٰ*�L鐴�ܡ^���b�Nў
��f��.	[���ɜ����7ERMr��������	�4D�5�JVe�3��#b�LGy
� �;gI�pቓ�f�����34���U�,�
�۰D43Mbԥ�Vj\��v���M�4A��I)o��dQ��J�v�v��tڄO�����Z6e���O��'j��ءf�(�>���3�u�Ə�F�H� �\��6H�?���&i�2�'��E�	X���= �u��?0'� s�]0_Wr A�l1l�w��!��)�Ɂ7A|\�uСj�9[w�U!ȼ�9�H:C�hI�Ή�5'Z���s��1@�|�Ļ|�1<Oy�`#H�[�Ё��Q >�� �>3"96#�IV�l+s�Z�6Q�)��H�.�pK��9>f�`�|��9[�f��;0J�'g哒v�B�[	2?��5�D6t�h�lZ9�"�"D�� 8Q��i^�,h$����'k����ֿA�ճT����.8���/~�l�H>�^?蓐|��E>�8��O"a~���A���}�D��>��l�Q�j����O�����Y�I,yش	Bn�5�ܹ�U+Oj��]�`dV�RGŝ���S��4,�Y{V#��Jl�H"D��v̢�͞�:��$��h��a���e�O츨��]R������<`��,*L=�S��
Yziї��^��5U2��}�l��aI��G��Od��B۶-p���K�=ZER�F�J�I�H=ZDP��&���O�p 궆J�K���Ri��2�Y٢�i]�Q�Qj���*Fy�'�d���M����&X�������'�lk%#9�l��?�$�|�&+��OZ��á\5�������>vP���}��4�,i��*0U`�ಋ�'��T��*Q�אWƑi�mN�s����ɈR�|�tmy�S���˼ng�<q�B��Qk�i��$J�U��\A��k��]a�.�69΢�[#�5d����C.�|��:OU	�K<H*b���V�B��3��>	��0����cn�ja�t�AUl��$���˶�ӟ~�R�h�`��HT������T�&���O�q�|�2���W"d5��I ���˥B�m��{!JF#>�<�7K��ɡ:�,����]�a��CN'X���K���*-�����~�O
��]�:�h�B��Ù8�@�+v��p��cb�A�0���`�N�� !��%s�n�'�XQ�IN�p��aaf�,"0۔�b�0��fc��홉yʟlA��dC
J��X�����Ϟ c�C␝>#������.���6�t���{*�FΓjj� �+�N�*A����	��O�T��m�\8TE�:@Av����C#Pv(���*e���xT&CY�:5 �yR.S/q������|�
֝3�ҠHwF�o:�x$�\�P��8qE!�4��aI��#O��c>�F,���ԓ$����@��O]��[�gԂ_�N<K�|�oĠf^���]�ޟj1
��������x���D�9o��`�f��q!�M��V��d��(���s��� �O�uI6H\�#p�b��' >a�]<0�
�B�^�d�rcm� c�,M�����G�	wV�2��
��X�{*�����K�Z�ь�B�D@�Ȕ�O�8(��*��+g(�;��U�p�$�?n ����FF8
5���E�1L���<���U�q��Ο;ȘO���b�����"$B�'�T�c�#_�{?��Em�"�{�C&��<�S�;���=��(tÃ@:LѢf���y����<yp��Ty��Mr��y��&�"���锐6F�u�d�к��\�>)�&�r��E��ʇ���ҁ�q��x�x�H��j�
�����2���S���dQ����:��S�	�j�4��Q4�cF>y���Av�33F�xXM�q��ᑣ�M>$��81g�|J?��\�MC �mll���S�R}&(i��@�dч
%�MR��Y�A�a�r���7�O`��H<	JF�h��9�E���6�?��'?��z�-�'�
D,�<�SVnڜA���Si�_���dB\$A��`"ȟp6I���9�O�KciH0�<��J�8d� �q"OD5)�F@;���h�k��P"O��a�ȕ(E�xhvG(w.�"O2�s"
́g�.��@癀2k [R"O����D]�MI�,Y�F��E�|"O�T��Ʃ.�]�Q���E�
��y���e�2�ia. 4�-��M��y����|���#�5��4��#�8�y�$#^��0&]}��=�Gh��y�n	�
H�<�s�Z�TV1r�9�yB���$��rΓ�:�����y"�M�  b$]}��h� �y⎈�q�����W�)�(|���ʉ�y�G9^�;�i[�W<VP�5�[��yrN�N��$�+VYz5��/ԛ�y�4��wk��7���RjR"�y2E� .\ ��RcȅV��`k\��y�AI<s�R���۔co��j�m��y2��:���z (Z�)6	�*�y��<4�� �F��<��ŦP��y
� ����7q"��CoT�he9G"O&�����+Z�Ѻ�m�3�2L�"O8(`+Ī%K00���zU���!"OԐ��z��v-��n>�ux�"Or	kB��s����LL�+!;R"O`��Sf^/_��,�R+��踒�"OT����[��|��U�`8qrw"O2�+!��x���I�N�8a،(p�"O֌����D��mC��&B��A�"O�ip�������u�TR��,�"O���kضlP^18A��umD�""Oơ�	H�w�(5q��2@f��Ѕ"O,�H�O�(���V擜YB.�ض"O�\��jR�hS@K^X�"O����"6-~1{��D�v"O(�zp�s�0p����N�L�;`"O5�`�Х�z�1nP����"O�-0"#%��1Iî�j�&��"O�˰ƌh	>� R��zjY�f"O���~�;��	mg:�&"O�Rܘ(]�(�%f�=U���P"O�r�+�(\=��g$ֳ1FD�U"O���L%�	A��A;!,P嘂"O�qI�$X�D@ƎҷX�B�%"O����	�j6)� �U*%D��j�"OV��Ԯ�b�i�O�S��2 "OX��0%�?gG
y�33fB�+�"O�)�b�E-e,Vh��+�4tr�˳"Ol�	��g^�Y�w���j��zS"O��-P��p#�$n��I�"O>�@	��NuܸqD�_���Ts�"O�1�ͥ7�l�� �dg"�9�"O�P��×�jId�xp�I-vaZ1a�"O��3���$U�xM����J[�=��"O�Jp%��]3*%�J�+GfIp"O��P�Ϗ>E ,���+tZJ�JU"Od\�V!�R@�؂,3LP͂"O�����Z���S���5f<��"O����㓤 I�؊1��4F&A��"O������Zֶ�dP�Y��[�"O*䪇��
 ��$�_�#�a��"O� hU��2r�� K悜+4mFգd"O$�ƫN?Nw�%��ݷwDv�x3"O88jozRl0�J�jNr�%"O����݆ �\������j"O��)������� ��K"O|�j7�>*(MB  S{Ov0��"O�l��F��Zh�bP/X*P8:0y�"O����%�
V����ˁD���"O�	p�^~��Q2�c��o���"O�EcTƋ-qo(����7�ޥ#�"O��0WE�.,�P���+tj@��"Op��D͈�6��E��aQdh^��U"O�(gJ��#q!�S��9X�"O��Ä��=�*ĪF��x�<MZ""OX���~���V��<�.( �"O:]���}��}��R2/�r� �"O$���,"��#p�ȮM$,!R"OBj�Ԙ|!Aa�)�/N���c"Oz�ؕ䃘LM���6OQJ	9c"O�l�5�Pa� �I��F��qA"O���G��;����,�"�$ 	�"Ov�K�-ZV<m[��ނ-���4"O���A�{� K5�R-g�,��t"O� �	��S��$�i	�)}�İ�"Ot�&��<` �QM�;���8�"Oi��I���ص1�K�0hT�r"OH1���~����/�0TWD��Q"O�����5�d��ŶEJLjc"O|1�&���w�tx"U��';����"O�p�����u$��R��W)O����"OLe@ŨA��d� ͅ�_�Jl��"O�`�A
Ҩ �Z�9T�غ/�̨�u"O� 厗�xCv)��,�71� ����@���	(�`E�bnx�j��Y�C<!��H�i��.U��{�x��	�'7~��p��l�(��N� �����'�8�
�O��\<d��VQZ�'�(|0C�ٓ)˼�Vb_���4��'=��यL�k<ppB"[�G�R�'��H�bϟ�)G&x+��տ��;�'l,�����w@�� �F�3����'*��]">OM�+@�(����'�28���Υ:�YR���pm��*�'�F��`ݗ<��)�`�ݕa�X-��'Gx��j��N��AK��TPb�Ҍ��>�'T�i���)_���+�s�H�ȓx���'����Nx��Յȓ �
�Bc`�E�z������D�ȓB�Q��Bߩ��,��L�&���hO�>�3I��`Z�a NKp!4TS�'D���P��
���2��^� 0��&D�8��`[U��+G�ʉO�*0��9D��1��	��F!XD�ē.��3t�7D�`!����v%��8�@���,5D�\H���*�D�����!�p\��5D�����k�tYr#ʜ�U*4�H�a5D�T�Sm.?ƔZ�ơy�bP�uE!D�P��� �U�R��5���~a��#,D�0x���w�.���kE�z}�tF*D�Ё��S:sL�ha���G�aiw,D�XqfnY|���`��([d��k4D�D����l��|�5+߶Z��q��=D���l@(`���Qk�7`Re Ō:D���gJ��k�6��3nD��%�dJ8D�D�P�e ��'��-N�؁��5D���ff.��G�I2&��m[��1D�\� �ܝ}�&, `[,��v0D�����|��˞d����0�-D�0�qoPU���s�^�"��hI� D�@�)��$�`��W!�Ʌm+D����&,�B1"&�<H��S��.D���B� �|���a���1�Y@��-D��H��R�
M���V�_{b���`,D���PLԈ)nԀ�b�
:T1Ha,D��rə�#!]���'"* 	ȣ�+D�Lq�)S�K�������-t�$)�+.D��­Ʌ�p��&O�nT�,A�,D��4㞮q�PM�!oK�
��xy �*D��S���v7\#գ;�4��C�)D��{� (	�0a��OG2LW�z5�'D��j�&[� MXe�A���Rg%ғ�hO�S"]Y���:������x<�C��71�]��@Y�G��HwȚ�.��=y�}��~2fD�4��@"H�;(9�[$l�v�<yEOƐ�:L ��Upv��$+�g�<��7enj!�E-֥L�*�EL�<�g����P�L�`0ʱ�TI}�i>E�=� H�e��5/�̫����rf���'{�O�y��n�x��I:�o�^��p�"O�(@�K� �#�n��	T��@�"OTD�"�Bhݢ��0R�L�	�"On����#0�� ë*���q@�''剜}G��"��) �=;��VxDC��:" fQ �'�$8���c�<C�ɟR..��2��7:���§�Y�n�B�%>�੫uFS8�0}r�/��j��B�ɤ#�v��dM݅9�'�qz�B�;X7������ P �+� �o+�B�I�&rś#&����e���MZbC䉦(p�D��FI= ����k�!|�B�ɋve�A0$�$t�\݈�l	@���'�a}"D�.�F�p�P9����'���yB��4�
��$�6\,+`H��y�oV-�|�8Ȟ-)��1��_�y� ��Ӑ��@< `  #�%�y�H�<h�f�ᒌ_0	O�m�%*���y�LY*b�bt��g$z�(�p�/�y�d��!~���ϗ�~�v@���ƶ�y"I��7�T�``J��	0n$ʀ	I�y���8X��Ӛ������y�E�W��]1K �x(^,K�eϖ�y�eIH��i� �֗9Ң���y"��:
��xqbC-p*ř3���y��9Cc�Qq@�$4�-�e)�v(<I����0��փIh�5�5& t����VU��
�/��J\��tCŲ�N���Ι9�'<`H؉��U9Q������<��+S?NxY���)1&�%�ȓ,3L-�� Y�}�P-���	&XJX��e�H�{�o��&V���fd	(l,=�'>ў"|�SPB!s%ߍ(hĩ��J�<���M�+����6�4����g�O�<�C��mF��Pm��l������M�<Q�+Q�N����*�->��jRM�<���0/��R�}L~0E#EK�<Yw�j9Dl���D�F.N5�"J�<Q'�Ka�p"�Ь(?ZpڅC�<IR*�gJ(�3�H/��h��)^W�<�kO:J��D���JҒK�O�<����pД��f�yu�����G�<�4$V8p�؈9G�:YZH(IE�Ni�<�ae<u���0�XB��� A��j�<�wf�l�R�"l
� ��Ni�<��	͜$�6|i���Oƪ���b�<ip�ֶm�t��Y �0!�e�<ѥ � J��J����C�0<j2��`�<q �;i���6��2%z��a�h�<�e�%�VH �ް;|i��.Z�<�s ʧK﨤�d���Q+G�q�<�3@K$4�4(����+<l��gp�<9���j��-�E
�#2�p��Hj�<9n��~�j���5�t5P�G�N�<yao�xU)����9��z�n�p�<��ę1H4R4�t�Tz�IZ�g�<A��K�g�M�6j�mN�����M�<Yg�$4K�s�'�$MZ��G�<� H�U;��Ԯ�w�N���>D��!&nL<w~Ԕ���1�8h� .:D��C�z�����X)I"<x��6D�p�F(�PA�%���Ұy���Ł1D��(w� �m�N�A(���a�N.D�� t������>�����t ��b"O2�" IN5�����8$�~��"O\�a��LK�4�C�C�$8��"O.VDP��.��1��^*�;"OHhH�N���B4F��M��"O>�
RƟ�����aK
>�L9`#"OzX��j��9H���U`0���B"OP��шB�U�z\���>]�"Od�#EA�k�*tK��A�2O��A""O��#��TdбpT-���1%"OF%u�J�2���ɀ�5a��u��"O�P;�"���,z�	VM�Uc�"O.Q���,"z `�#K4s��|Bd"O,�z�B�Ae�M�gRz��̳3"O��A�#�X�|( �J>$���s�"O�7jT�$��{��h��"O��+Ίw� �2�R{�L�U"Ota9s R.��a6�\=Li��(f"O~�(��G���j��sRb��1"OVQb���3"��2��DU�-��"O��`�] 
FYa���Cf$ȷ"O�h�ݷQ��Bvj�: .vdG"O��J�"��%��Ä�~B	��"O������,\�R���!ob�3"O�	'㑯It�(��郇Fe�5jQ"O@��Å1MM���^�SX�SV"O \PF�Mc&�ӧ�|���!%"O �swlR�[�l���D $s���5"O�yp��Zt�y����c�"O���,l�rB�֚o���	D"O2�1d���	gB����W�yT��"OLt�W#�#8��Hs�)ЩsWblRq"OrT�4���n�jP�H�7U8 ���"O\�C��]�2\���6|�2:�"O�`����Pꄈ	2�EY�`@$"O^���n�~�(8��<GF����"O^XId�SH����.0D:ɡ"O���3Ɠ5NyJM��M���ꨛ�"OD�p�<pP[Q����	�W"Omx�M͛)8
dq�ˉ�j��aS%"O�\y�A~�Kt��z��eK�"O���e��T����+�uθ)%"O���f�t�Ĉ%+�0f�!"O�1ƨ��PD�(���Z�-K��q"O(h kܾ~�80BA�.CG���"O����Q��6�	�o�\x8PC"O�:�I��i��]S��Y�wH^�X�"O��R�l�@Z�� ܯ��I�"O� �`�m�\�"VD@&#��dz "O^U�"*8�p娍�.��E"O,4#��I_5^0�G/)�2�xS"O���7H�>\i��;|���p"Oޑ���͔s0����P�X���""O�abC~� ���Й(�8trQ"O���5�ĺ0fQ����i*!"O����K¯q��%8��D�W���"O��d��b`�uI]v�cA"Onɩ����{���"���0cȠ�"ON����K/2 	с�2`1�u"O<�
��J_��Y��,ZfHs�"O��9c�j�Bt��gX�#d"O
X��V�<e�����rN��r"O��AcB��D0Rf�Ŧ6j  s�"OJqS�i8�<�$�84��"O� ��Yb��r��� �L��`vX��"OlL�&���z��x��F������"O(�2˞+-ʀ�V	�X��F"O�0��]X���%��B�x��"O�*��\�}�L�$EJ�56�xX�"OF��ҠI�wJ���J.Izb�"O�$s剖6=6��i������'�<c�O3Z~0�����l��'K�Y�w����Yq�L
��'L8�tmL_��E��HZ�Olp���'�25c��Tt��h��^����'�V<�RK�6E��[��-%���'i0��1 �y�
�X�'P��;W*ZD��rD�3~�D}��'X0pZ��-L��t���ɷr���'��e:P�Q%5p�d%<n�j���'������%$����s�ȇs�vI��'����-�NN�Z��
�f���yI���eҷ`�)0�9�bD�y�+�X��7*+�Ȣ2�ͦ�y��G!UJ@���������y"K�7��=Ч�"b5l��G����yRI��Wd���l�	Hs��	��E�y�/�J�$ �$��A�H��g+V��y�&]�)�б���'?�.��'���y"�	<�SJ�27���6���yb2g��˴S�(,��3�)B��y�3E��Ȩb�L�T��X ���y�eQmN�!� Y}�<I���yr³?�85"sGT�d�`x�B��(�y�NArՃf��Z��M��B�8�y��#�`�6���A��LK��E��y��-�qrU�нj�������yR%�P�HD VJ۝t�Ea��W3�y�,������� �mU>=Y�O��yr�I�>� ���4R�5��!ދ�y����cHmhc��\op)ғ�	"�y��RV�E85�*U�m*�B�:�y2
%J�v%��kY	ǰ�4��	�y2E9Ef�KJՐ>b�5)���y���04 @�J�7d����M:�y�o^MZ�kf
cY�ԱQ�K+�ym�n�2 �5l6c��Ip�K�+�y�9[������T0g�`�Ύ�yB��YY�A�3�zj�y�p���y���IL>)�Qe�$s��,��yrJ�1q������)L������A�y�U�|���3�$-�>�1G�
��y�/Z�*}�t�À"�<�6�ڒ�y�)
�~�9��p����-���yr�\3v4ʁ B6d��8����y�	�"���q�Z.&i���t�,�y���W.��`:������'�y�d�+hqX��f��\������y��N��zIѐA>#�$����y�.��~@�w�ߡ&� �E���y��iT��hZ�P~0�H�)���y�j^�R�-@�Sf"���+|hC�Iڼ� ���(N9VM�dGU:^(,C�I5��@ UfJ�;�2U @���	z
C�	�\@�m��� i��p�S=B�B�ɍ@������6�����C��B�I�t��I��g<Z�� �h.�B�I[����AI�4>Hx��?x��B�)� :�@G݆Fn~��G��7����"O�QGFGw&�(Gfү=�����"O��K
�;�:00����<�	�"OzM*�gF`D�� �o�����W"O𵨗�ֺ%˔�����'U:� "O:��#��W1�Љv/�r�z�"OdE�����X�K�MΨ&nfl{�"O��Y7MB{d8��l�LU����"O�lR���y�N!� fcN�r�"O+7�N�*���2��4XH���"O���m�(������)u�݂p"OVqbP�ѹJ}��Q�])h"|+�"O"�eG�b��p��$k|���V"O.죳�B�\D>�!�gϨ#��F"OF隐C&I4\(�+H{�	A�"ODٻ���0h�2��T/x�`�'"O`8�B�<�PZ5�T�1af2"O.e���=	��1��½5����"Ov	�i�Sn�:AɅ9:~ ��"OH���[�G"<\!#Hkg�=��"OıI��ſ7.P!�MU,O�y�"O�� �,��n�F=��h�-�y�ȓT��EkcLu��T�4��1��ȓLq�,XR�"�l��Q���:�<��ȓ6&X���ك/�Bh� ��3Hq��'���g�8~1J� �
@UH���H1j��g`��aJPc���d�T��3p伻v)X��r��i�19��ȓ2�{�g �<�sg��dF��HE����`�c�A�䭖�u���ȓ�U�N@�o<Ĉ�kQ� �lz`"OH1*e��e�t\ST���
$��Z"O��0��_�^#$U9̐�E��J�"O`0��Ʌ�$"����R�l�"%��"O،�&��~hl���8~��À"O�U3�J��`�ǉ�#Ke���"O��aŃ7PX�y���:~_,d	�"O���Q�`< ����V pY���"O�Y��_.Kt����8a�di�7"OT\�b���M��0 d�-$��"O !�8~�	�u���$��%"O�X���G�"��a�Ҧ΄o��8Q�"O�l1j|9���&��t�,z�"O��y%,R2�>y�D��-:��"O�Ѕ�W<y����@���Q"OZɉ���}�D��bŗP�Ȍ�F"O����+��n*�=�g�Qf����"Oȴ&, �2�v�
5�V5�"OTl
��6`���kg�^�B��h1"Of� 1!� �X]k�WӴ<�g"OLI�W�Ѣ2-8=�� �	y�Z�j�"O$�r��4x�x��?�!:5"OJ��D��437�8��n�8F��q�"O�;C�͒"鲵p��ݟ����6"OE���ˁÀؘ`�
���IC"OR��1�H; P|���8QQ"O���@��L� U0�λK!�e��"O(A�bU�f����f�c�}i�"OpD{�G]$��iKс�0p��"O��+	��	�@i�UC&"O^PB���%y�r41�����l�f"O�D�c�չ"�t8�m�$�Z!i"O:��A.Y�h9	�K�C�(�b "O�Z3\�V� ��*�����"O� 	���Q�	���!�X��`�"O���,�^(�Zd
��k���5"O$�2��?N��Q�B��"q�����"O]�t�C�/b	�6ކ=�\q"O����K9O�-9��� /��q�"O�W�ZC�訐�5/p��R"O<�s`��GkX���c	��͈B"O2�C�Ja0�y�B�R�8�)�"O��p�L���P��W�]8�\2!"O6�"��
������:���"O�D�dd�؞q��nK�W�z͛v"O�<R�I))�<hhpn5�&Tۃ"O���04�ze�@�M�J��JF"O�3w��mhm��ѵ)�0Ñ"O��v�M_�Ͳ��4pU@�"O�$b"��>	�
�xFk��f���"O@�P X'��D�h��\�@"O �{p�E�`Wt�Ҵk�i��"O,�3&ᜥA�$�
����c"O���r��b�`��)�����	�"O�p����K��IQ�� X̖��"O�$kQ�A����K��P!g�0�*""O@U1��4�r� #u��-�&"O�� ���+y�&��0Ȁ=->�KP"O0`g�ܒ8����Eą��"O&P�&���^m�6���>Q�3`"O޴����rR��Cc��xI���"O� �/� 4�fDIw��>C@bM�"O(����W-Urt��( �@$�ah�"OTP�b��A�ăp�̊R?A�7"O$�qCeD	W�e��h�P2(4ZS"Oڜ�#��,z��:i��~C~�H"O�}@��<c����B�.A]���W"O�u�����@��\kf�	�`�ĩ�"O�mrRąpd�Zw�&mtv�p�"O�=Ӄ��4:���S�����\���"O���YhD�hF�y��%X�!��v��8"�4R��]��A^4!�d[�OZ:,pcd�2��y �e�*!���W�@�9�-�@�2�ÿ3!�$��WX�h��Ƣ6y���C$�%!�D�Z�` ��rH0p�d�8�!��gDp���O,&�9��'�!�䋕Z���*ͭ:ji�/A� �!�da���E#�͒� ��G�!�DZ�+ֵ#3Mһ5���
%`��l�!�d\1�
�Ih$;�L͙��?{!�D�)��svi`��\p�NU,>!�$��?[�1����ڲA�!��MT��z��_�P}B1�D,W�V&!�$W�|�tU�̻!b���$吩 !�@�9��q�e���<U��+�*V!��C%x2`Jq/оZP��\?Ӭ��[�<h��c+9� ��/ĠK�,��w�r��2-����B�$$�&��u�8����7HD�)
�o�i���r�r��b +C�T��ț5{�4	�ȓC�<8Z�I�K�\����N�Ʃ����-�UN��Gvച�C61r��ȓn�V�JUc���r#��J��M�l�B,��@�h�@V����ȓ�Px���]�=E*N8�ȓJTș$ĉZ�=+OUG� ��ȓ!���P�BUJ��=6�����S�? ҅�'f��[p���Hԡ1���U"O�eYP��o��	סǿI��ñ"O���W�Q<L���^�bvu��"O�=����ׄ��p��g:��"O�yb�M�|��]��o�:h��y"OdɃ&(�44/`���	_�]���E"O�H�(�J�I��*J)���"Oΐ���X>^��|��吃$���"O(����=)\j8�$�;V# (f"OhIJG�Ӭ=@	 ϑ�]q���"O�X�3�̞!���NF�h�q""On�т�ɌJ3ֹ+F�CK���e"O� c�@:n�� I2j�_|�"O �X7L� mR2lK!A�W	��sT"Oh<K�&.u��<�cT�P[ڱ0"ON���:m;���%(N����"Oh����s�d���`��!���C"Ol�s��mZ�`n��F<0��"OА���Yj�dR��ԓkx�"O�}�F'̽i�>�XU���7����"O ��$j�+}��t G�D�z���"O������0򺔚c!�'|���B�"O����+@�1���F��<�t��"O�Y1���f�́�b��<�.��"O~�����L�X+v��	�$A�"O�,���*4�|�bk1%x��W"O��1`gT.`?@yc�c_�!&Z��#"Ol�n
�jJ���$��%"O���K� o8� ��A(J���"O8�Jp�1����y��c"O�@�V���@�2a[�I��-(�"O����q^"�Y��]�@�����"O�U!�m�=*l�J ��-�D=:"O�TP��.eDlBs�[�T]�5"O��Q\&	0��B�!Q~���i�"O������7ߪd@7�Ke���	"O�=�qJ�:i�@tmǼt� �f"O0�a�̕�\�`���+j���"O�����"���R�.U����A"OPj3�P�o��h���.
��"O e����6 ���k�6l\�"O.���4>	��[�jVI�AS�"O� �r$T�j��iD2J�d�#"O(�p���5]Wn�j��X�eS�)"Oh��A��ూ��2~�z{w"O�XЦ!"+�p�Љk�v4�"O��#V%N�Q�U���S�h��"O``fN�%&�h0�6o�1<��y9F"O�]3Qd��m?��iSMėC�`]�"Of�+�<�h�`���"OE���^��D�EQ3�F1��"OR�r��BB^��i$9�A4"OJ$8T&��e=�̋r�K���s"O�Բ�HD��P1ƭ��|��"O�;��z�:��b,HsE.��"O���!�P$&�j��a?�݈�"O*5�biGA\$z�̘�N����"O���aH�'��d©��T���"O&�¤��Z��+W�O �QR�"OL��Ō�~�tP@'�4J��K�"O8�6��oA��[�a�l��"O�,�a�ގu>]� %���"@"O��+Fm�4*�xx���
�`}�q��"O ���#�8N*���c�?{~���"O� �s�eN#J��m�7>P���"O�h��F���	%�N�9A����"O~,�K�-D_�9!S.Q1V-�D:&"O�0EJX�����[2B��P�"O�a8�_38��Sv��n�BU"OZ������ `��-�8C�$�b"O8<JfHI.�jq0�윪P��}�B"O�e ��Ւ|��\�kԦ1��d�"O&=ȃ�/(����ŉ �j����"O�Pdh�
����u�J#��hb"O�uӖ�NG��� j߸lpJh�U"O4�7��b�x{Ë=h��`��"O>��0�֑~ 0�2��w\��"O>���a�\ �¤B�;ibݸ�"ON`r�F�J�6���]�`�a4"OH�#�A�)d�M�ʣaWV��"O��bզ˴ ��y� ��-i�"O�9cÈ�r�xT�r G3J3P�I�"O����ADI�4h�/�:/���"O�!��`N� �:�`oB�u���"O*�3���I�H�8rM�+ �PT"O���h�_ƌ��@/*|i�"OL�,]����*" ��7E���y��
�ޅ�ɪo7|�򦉥�yҌ�%v��yp��yD���H�"�yR(��I�x�`��%o��l�ê�?�yR	�W��K�*<iA����j���yB*ӟ����Ei�����.���yR��9�lXhTLK�^������y��+

�h�����\z<Jg�D��y�FF�\g.���.�����Q/�y2͟�@�Н�@�лu`T����y�+̌6��؈$�X�s����F��%�y�#ϖ��DQQ����#��ʉ�y��U-+Ҹ��m	S4y����y�_�g*��K�	 }�1a����yRe�� y����X� B:���g:�y��ڹ<IL���
�/U������yR��6^B<�G}�Hz�c��y�k�1u+>̩�+���
U�ه�y��W��L��cE������O?�y҄n4:���dT�=�ȃC��.�y�CK��!��HӔ��>
|���'�N@+3�_�r��$_\�!�'�����&-d��ئ�L�R��y�'��\0b��
٪k�ć�PʂT8�'g��	���4�
��t�T�\�h��'���a d�-p�maD҉>4�k�'�B�Bp×T�-h�&�0rz�
�'�-"��4'=(��	A&,�X3	�'@���ç�s��q �uKr�9�'�f�XU#�>SU��%lpؤk
�'��$8��L�����]9i�H"
�'�Y*�BPD̡e���Z��8	�'] �#ə�@��d�%K=��'�2���䍵@$�æP�Cv���'B��*4�.�� <����'��)B��7�iZc�Ę:'¨Z�'+z�8�&EU�r�1���1$Q�'�A���@�x0B	�C#ǌ-�|y8	�'�q�vd��eFqY&��#0~�
�'�B����	;�x�ɒo>��'~!2i�
X�(��DU*KzBР�'���1)���Pb��0W��s��� 4�(�A�V�u���ջ���i"ODLhQJ\�H��}�H��"O�E(V�W�X�����;�J�d"Oj�Jƭ�2g#h�H��:n�P���"O��Ԅ�y�j�B�;+���W"O����U�-L�]��E�{���#�"O&Q�#ύm�4�[�c�'K�:}��"O��r!,E*.)z��� W�VI�S"O���!#q��+��As��� "O�e`�
�m,n�k���;T�^�+"O�͹�,ڪ=� @Ǡ$9�R�	�"O��PЎ�1ڄ�	QMX=>����"O�]��BT����G:�|��"O�M�0�<%\�*��o�<��"O��;"K�&\p��I�h�*��"O�TYU�0^'��Q�c�Vт�"O��C�����1��<�^d�"Of�P�L�u���õd���h���"OT�+�)��Z����m�5��}`�"O4�%��/�����G	`j��"O԰A�m�K5v $��`t�3"Oj�pfd�ԩFe�=�"͑R"OL5�/�PU�ĤQ�rS"O�a�W�׏>)��《A�~��"O>�ʕ2]���6���=��l��"OV�2s��{̄�C�(/x�IrU"O�	v���ʐ�#?e����"O��4+U<��D�0#Ί7���r"O��@7a��>!�e����U�p"O�eZ�A�z���'a^�O:r8��"ON��DI+
��˦��($���`"O�Uq'N<h5�ˆ�Y�*da��"Oz��c�!i'�(��V�[A�t"Oj�d��hJ�!� ��H�"O������y �� �Y]�lsw"O�h@ʧ>���(&DO#�l�"O�r%������P5x��D"OfLK�A��=
����
(W,�!k�"O�=��ڭV�l��ՠβ_E���G"O������S����%f��[�"OH�#��5*l�����J�Re"OD�P��8t���O~.m�S"ON����R�\��S�+�e ���"O�(�����iapkk�(�{$"Or�3�oK)9��"���R��8f"O�,��}��-�G��`�`&�D
!��.O�T|��JXpS�=����16�!�$V.*���A��-b�㑥�Gy!�DL�0�(@Z�N�&���W�ѓ_!��m3ΔB�l�
���B�!�$)j�v	;`�\~(+r.��!��31%�Ū�ɉ������ð:!�$\�a��B�e�vr�L�c���!�dB�'��8�d�Dzs*	�#�R2�!���u�^�S�� h"�3�(!��K+	�ma�DP�1�և:�!�䍭T�`��*A�F��څ'�8�!�$� oEv0���*OB��)T�V�b�!��9.��@!$�>7���GѤp�!�d�R�lq�)
�j?DUYD���&�!�
(�h��2-�=*P���FZ�pb!�D/KpAI�n�9��5e�:`^!򤍭��@O�1N,�A��cO�!�$<�ʩ���{>P�L��E�!�� �@�C.�n ���gQ�"O�q�Ҧ�v,�\��(r
h�k�"O0 �"�B���s��O�4]()!g"O��hCnT�L���C9URH��&"O�4n�!T��M)q�	<g���` �1D��P�*�<wLY:���
�	P -%D�p�hD�G�{v�E��a�5�#D�L0G쐳U8Qb�ǝ>R�V)�� D��3��4l@��Z&�WI�C�g<D�HyGb��9�Xy��m��O��i��:D�lx��Y�:pؙ��ɞ1s>�y�R�"D����H�L
\8�k�����N;D��8��׵7�FIi�腔6C�m9�9D�l�VaیC��CE�zV��G7D���u���3�d��6�^�Jt���8D����(�9�V�ܟ0d���J*D���1�4���@�%�Z-Z&5D���d��ALfP�І��^�t�3��4D�\��,wI�}B���>1O�����(D�l�7�<cE��ys����i� &D�|��Uw�}�3�E4�����!D��I&n�	�`I�p��
S"��z�)?D�dR�T�BR΂( ��9E�8D������l�,H����G0�8Sg�6D���hʉ��K��T/Arh���?D���NQy��!��S+R�4\�2�;D�ؒf�.+(&���]�*� ��G9D�(��-�NLx��5'�
'�#�c6D�( 5c�[� ��HٱU���A#4D�DQ�m/�-#��2ل\P2�-D�T�Fc�$���#ϔ06*�Mj�o+D�<٠g1�� T�=�J4�V�'D����ɕA/2Esm�O�Y�g�%D��hŭ9��J�ǳ$N}juA?D�,�W�b��+�x8�eI��3S�C����pS�@�h�����$Y.=lzB�	�m�v���s8JMd�\�p�`B�	:a����n�N�@1`q�[kD�C�	$o���LO+#�*�q�C�,^�zC�I>l������46	��С��U�^C�	OS��Aɋ?�����>3Q4C�	<ed�ɇc�`��y0a�,H��B�16�ةP�֏JV��QϞ�`��B�ID8���R���vkA�8�ZB�	 G���5���K�U�V��=�B�ɤt��1pPD�Mtd��T�ݼĜB�ɟ4C���1K�?��z'�@(o�jB�	&�;���U���+D�P�ZlTB�I	yα���S6��X��`Ϊy� B�	�U����B�(���j�d� L
�B�IK�t԰
N$�bPХI�!0R�B�	�rJf��&�G=a�yE��8`�B�8ZVX�G��[d��i�`�~^B�I��\�  eLr�A��5r< B�	2f<桒�$t���#�GG�a֠B�I�xih�AZ!J�I����'T��B�I(���c�'&xAh�+ȩ}m4B�ɡ_蹱U��:@��kG�I�PuB�I�I�d�A��>۬�9@`��.��C�� ���a��4]zA2���w��C�Ƀ9C�l����{�&$��
Ųz��C�	�@�:����^6(���+2)�C�!�t���Ĺ"#�|�TH�	�C�I�1@,hu��Y�j��s��~m�B�)� İ����A��d
�j�mpe@�"O�4A��M��R�1�/ �c M��"O����Ξ3;I"$���;@�~ݛb"O�z��BxѤ�S��ׅI���"O����7:�X���DO�U�v"Oڅ�`�:���7M�>)MB�6"O����!�g�Nh��+�o]��6"Oh�k��*02��sKB;)Rh%c"O(��u(�f�T���	E�DDRh��"O�x'-�z+��#qn� =�0E"O���sعZ#�غ �-<�YE"O�<B6kɖd4�D�̘�/ ��"O��Rt�̊o)�ٰs�}��sD"O@dS�F�m��L��X*S�6��R"O�<x�A@*<�^���J�w a��"O��Rb��>A�f �&��M~��c"O�ؐ��'pc��K��N�����"O��W�ߦmW��Z�'N#B�y@"O|HR$� (�XTM� !r�K"O�����`5^��WL�nd�� q"OU����, ���_�$]��"O*K�쌔.A�rH]Bz���"O����ǒ��0Z�ƀ����E"OX���ԾO�M�%���Fi
q"O��@�%�$���j1e5[���H�"O�0��3g.��"�T����*O^�
�OO�Sн�A�@�T�~X3
�'�М����)_�|�q�O�:�Y�	�'��)#1c�$X=Z@  �R
3�z���'4�U�ڐb�|����S��$#�'�=��s�("��z�Z��'3��%Ab���aAߘ��
�'��1�a��rk���TjOy|�-c�'��3����
х��m:չ�'��i�R˗53���ڠIƀv��I��'6�ɅEҢ[rΐ��AJ�h*��'j�B�d��
;Z�" ��;,<�x:�'G�a#ab�~ 	��) 5(�T��'��l�D=�r�T���O�֭��'b��Ɔp����ĭ<]���Y�'9nu�T'L�P��i��j�.$�>�	�'r�Ha"N$my<�0ũ=_�@�	�'*B9�fL�H�p'�_��8!�'�.��f�����Ϸ3�V��'���.�,�3��2 (��
�'_f��C֑*�C���(y�8
�'�j���Ғg�A�ƍ'�EZ	�'�x��E؇p����7IשsU¹ 
�'݆��ц�>x&�l���g!���	�'��5Y���*0	��!� a���'�EYp�O�"�,�"��&�n���'aԙ�p�E%<>D��6n��h�'"���F%�7Pz���.��(���'4(\Ҵ���!��� O����X!	�'��{G�Ё"�L�/��1`V	��yR��9l�F������"�fǃ:�y�&�ff�@3>>2�aW��y���yC/
�M�l�x��(Ge.��ȓ|".4���2S�2�[��S�vk>P�ȓ]��B�60�6����Ņȓ����2��1��+���"��ȓW��k�&O?!Qh��n�7Dd��ȓDD����'d ��cQD�7�>Ɇ�G�[7Q���pe�Րn(��S�? B�Ќ�$'v��Q�D�.*��P"O*)S���Qy�'�P�?|jh�"O��R��^7
�]�c�/ ����"O��+4JD�C_^eb��I���آ"Ov��G�9e?h���
��m��4S7"Ox�����=w.|��ԩP���	�`"O�D �g����J��zX���"O�,�c��u$L�)"EDڡ��"OqS!�;6�hH���X^)i�"O �����2ai��	%=��=�&"O@�g��`I`tг)ԅ`�z��u"O�|��#���C���N쒁"O�ܫD�&1,t `�*"O~�ϐ�JՖ�CP2�d�Q�"Oࠐ֥��VF�6�§d��m�"O<�R�O�l]��@w��s����"O>�¢�X�F��=��E�t��a�q"Ob���C���v{��նk9��Õ"ON-�Ĩ�fΤT�V�ٷ8�p V"O������Y-�䆂���q"O�4�i�!�}�ť2[DX��"O:�����K@a��cQ�*�N���"O��x�0E��Q���rMX�4"O�آ���g-}�W �:(KL(�R"O��zt��(x&:�G�_>��`��"Oe��)W*@!G�0�-�U"O��pŉL2T�LE�Q�~~b���"O��&Eհ9	�7�i�l�b"O��bc��)���Xs�>\fv�p�"O�4bt&B7,xe�&/Ƕ"kl)"A"O��q�`՚(z*�>q��tS"O���!��}�afMĭL@m9g"O չw�$�L1-Y1	bY�"O�͘rK��(���̅�,F�K�"OX�h�$ʌS���
�Jը3��"O�Ԛ�ʛ*�M�s�B|5p	��"O��q�'Y�R� В��'&̲�a�"O�a���W��Z=~�l�"O�y珈6X0(T(_)�l�Y"Ojp!B��*�5�Gh�{��)A"O��fj��2��'���Ct֝��"O���NS m�8�iN,�N� g"O���'��CI�L��A�7�
d�e"O�hq�HB�6H(�a��8�D��"Oh��$�e(H���G���Y�T"O�Pc�JևV9|,P'(Vt�)3�"O\�'��I'��Se'@cX�a"O�!T6=F�	I�@n$�#"O�����L�:,P��@�)h�4��"O~e�d,��S�^)#A�I9-��%"O��	K�JY�e�T�O� +�"OHI�1劽Y�J�QUꗸ0R([�"O��;�X��H�~T̬��"O���1�h�0a3���msf0�f"O~8��,Γ9p�7��3_Li2"O �(0��Q����e�%gU��yV"O��ME\*�qPf�;,Txg"OrH��Ic�<�av��$>��"O�%�o��琬�2�K*��u��"O�E�CÄq�� �
Zۄ3Q"OP�!Q�'R���(���.���c�"Oĉ鳧��:�*��t���l9��"OV5 Ư^�am }�U ��y�H�"OD`im����ɲ�L,\�Uۧ"O� N�s�N�Z�L>�^hJ�"O:u���o�љ!��e����"O  ���<���Au�I��ty"O����Bg�0٫ظjE���f2D��r���Z��8�( �lɑa�=D�́ )�xi�@�t4��ge D�H��ƃV���С�߈$��}�q" D�lb����U�� b$�����T�;D��^"A�֎�1<�b4�Q� �!��M#.Y:#K�9&ر�A[s!���{N�Zf(�i�$�ЎѺT=!�D��gY\<�E�����'��[�!�dϙ!6t²K ��}�uÑ�\\!򤉼k4��aAN#L�&���I�>!��J5a&*��L)}0�I!�*�&.!���4MA�PBJ
4$h`;T��R(!��RRL���Cq�Ř�H���!�d`y� �T�G�+�Hy���'!���B����&M?�h���Ӝ!�$��Pƺ�S����.�B�i�@7�!��ݫ*������ǜi@�jvn٥<�!��-^UBW@�)@v"�˗,M�m!򄀈eTD��j� ��U��ݯM!��C�A���c�.��+�u�%cJ9!���F����DL�,G� <�"½O�!� uV���s��(��ͩa��=!��0I�>�i�,B�Tl��◤��M�!�D�>y��M)
3nd�4�V 0!���<μuheM��6����� "!�Ĝ:|��
])��1{��S!�$΄!b�! *�\�XaGo�@w!��P�!���Γ�s,�J�/!:�!��NC��i8�H��5�����Pgf!�$��rC��)2�؉>�E(B�B3IW!��2�����&��"t���@A�A!�9�ҡ�E�^��|�ÀE��!�ĵN&08$� ?�&�B���!k�!�R#Y&��Vb��?����s/�o1!��	<Bm.T1�pBl��N�\-!�L <�D���nY� qEZ�!�L3�HN�\�@���#�-�'�&�����g�Ĳ`'�=:�z�*�'B��1+��TN�5%H�:�px�'��q �eT#f+L�D�B�1� ��
�'}�	ޅZ��T��-�.�=H�'qH�#-�9 � �2�)�L	�'l�"b�( ��؂��:�� ��'Hf�e�6
Lx�CJ#K��r�'��$�ʡ-���#d��B�dHb�'�r@��Zm�A0���>� �'~V�!-_|�c��1+�T��'.ؠQ�ƴlA>�!˃�&�|�
�'3z	��h�	Z����ĕ!3�P�'����Pa�e�niy�oμ�����'��1���ߨn]m@3X~4  
�'��c�B���r}����.c���Y
�'��RwbO�	|�Q�un@�o1B5��'ٰ�{��ӑ9��yZ���m�H�	�'rZ<���J�3�B(�3���d"L�'���u뚪�j���L��X���'�� p���I���pbA��0'�	�'�h��elϾ0�T�`�e�r�E��'�R(+�N�d����A�X�~��
�'G�t�BU�%�mK.�,L<���	��� 2�r�P�B+,]1��zt��v"Ov8�Bc>Kj�������C�"O�1e��](��@U �J{N�c�"Ob���6\��p�Mxd͹�"O�АC�Dt���Q�AtY�ȉ�"O��G�^�r�	� zKµ�C"O�%��g_6Ԕ`�B�6a;��`R"O�<�Q�)\C�Ի��Z0��}�"OJ!�#c��Z��ѱ(O�ݲ"O�T�/-F�8��D��<¤��"O�컴
�6q˺t��Ą"��6"O��lI1N r�@í���|H�"O�UQ U7��سkЁM@D"�"O�ŊR`���V��#` 4 �P"O6 �"�j�f�"d��,���"O$��4�
+@�j�dѶu�H�"O�3�āT��Ug�ҕ[�"���"O�����q�J5z2�ʑ��А�"OZ�SaKX�QZx��M�(���"O��GdL�2� P6�G��A!�"O��A���U4h`'�>g}�ų"ORᢁ��$
�YB�Ғeζ��d"O����M
\}P��F+k"�B"O!h�R.=�@�e�D�]��Y��"O`����EI�e�Uφ.��=ۣ"Oܑ�d�df��(K�_�F���"O!aFe7�^��ߤ�t��f"O�,� �U�2�pX�@����ѓr"OIM>
��(Js��(�Ҭ2B"Opa��
�R�l�
`�/~��ly"O5Ô�M�*���Qδ�"OP���N��B�"�C��$�bК�"OZ���dP�4圼R@R�OM~٣w"O���۽P�dH����$=��"O��qظVߊT�n�[�p��"O~�@�j6�x��"N�	��� "O���
7Hu���;���F"O�ܙ�e�����I}	�C-�6�y2�6=��qWKz�dYjS���y������x�$߸vO �����y�B-�"���/E#J���BF��y��[���I�ɀ��J8�".�y�� 4�Л��In|B��1(���y�	@:%iЙ1S����a��$�yb�F�����ԑ<��A覥KE�B�I�=8�F낝N�@���o^(C䉗=,DX�� �-\��]� R,L�6C�I�7"�wʖ�ڑ�*�&]8B䉦7'U�N_�p�Ga� С�U�2uh$0!�]4nN�QA��_=\�!�$e� ��A8}bd�c��ѻ o!�#?yxй�,��k��1ZI����ȓFrD"M�)d'���.Q8��Y��,fP�)��X�`�i\1G`�ȓ�p�xļ0��9F�����F�<QEA��(��̃�IR0^3Z`�dJV�<!`W�N}2�[SC�ډS��{�<�e N���A#d+��ZQ��a�<qfϑhm��ᕅ�V]@ �5�x�<q1	ӌB�Խ��m½�V��R`Iu�<q�oVF�� ��193���{�<Yc!�)_�Pl�5�îj��	�Zn�<i1�Ӕ@P��r!Ӭx�e�6Ql�<7oÉ
�tOB�
dmKc�j�<� �QI�ݎ��5��-V,O��Uc�"O���"o/MD� @���kxt���"Ov�aU���		&�D�M:u!HL�<���&*6��dL�8��	1	An�<�OJ
f�n���W6�ڬ����N�<� �^<Sz��rƖ����7��H�<�F�W2U����n�#���0P!�B�<A�^�v���	�̀�|q�`�GY}�<鐈��0�K�� >᧏Wx�<Yp�	�$�U�M\<:ƒ`���k�<)��ݟb�h���J�t�t�h2'e�<ᦡ��� �3�(�sH�@�!�c�<���[�:��Ul[�	��|�@�x�<��*S3k��5l3K�:�b���{�<9`��)\_�l𡁀
��jr�y�<q�h�pɜ�3�Ŝ�R3�qp��@�<���*]�.��S炄fF|���^u�<q�ۘ2ĨmpA���<6{�<��@�s�.L�'Lp�Ȅ1�t�<���;��0Qa�75;dQ���w�<�g��1 e����2vV� �j}�<A�-��bQR��������WÃ|�<Aqǖ�y2�!k�vn�v&�x�<�5�%ER���B�n)����N�<��C#),L�qc�B��#�* ʄC�	���u�o�:r�� ��H�>��B�Ib� q�E��)�|[���V�:C�I�cV6�JW�3HMJ�pĠ+��B��)qf1ZV�Z�j�f�"b,[�[��B�I�y/0apAP ;�zX����<g"B�	%�*U�s�c�� ��n�,�f"O�@0�Ԟ9����@�p�T`!D"O2�S��O,I������0�t|Cs"Of�9�`ǖ]����ƀ��7�`y�2"O���ơ2s�xJS���a��}�B"O�|��hʔ81�� ��i��C'"O����n|����0��$ZNr԰"O�$�A�I.��Л��MI9K�"O��!���I����79i�"O�x����Z׼ h�YY��]�"O�a�ufH�r'g��0���i�"OF�qFg�C� 	�G%R�"�8�""O���\;�(1�f�M�8^vlzp"OH����i�.5 #�$dm�ɡ�"O���L[.7��1�bЭ}c�[�"O��������S�\�`>D��A"O����EGĜC%!��:!bIc "O��Q�'L:;&Z��`��r�vq�B"O��y�k@7���S����j��!�"O�A�"oL�h��V�˅Y�Fd̰`�'HH�R��֛dn����BT@m;�'���(� E�"�Dy% A�x �
�'v�h��1�B(����2X���	�'jAr���m���&ɕ�V�6�
�'[dŒG��S^���uD[� Q�	�'&�z  �P�氱S�|fj�K�'3��&�5���3��oӘA��'����r��Yf\c�(e�Υ��'�pl�P�N�*�E�G	^�j���'���՟>����y2s�'N.�$�Y0L3�Q���Q�vI��'}��$�L5D��x�ЄF��V��'
�J��[�5�����]�v�����'�x��t	�e�rM�0Ch������� ��$�J�/�`�iDe
�*��;�"O�"gj\�W��%�7��i��"O,���ݣǲX�a��C��E��"Oą8�싓P*Ȱ��7x���h�"O�5c�j[1���(ԫ�<W����"O�ys�j����ɫ'��H�Hm���'�<�n�v'x��Æ�zg4!h�Y� Ӽc�(E}"�>�4��@���N��,3������k�'+�-}B��4,Z%	)�ݳ�)ޚXf���)_%�O��+�[E�bG:E6�DC!KbX��V���iH�y��9O2Հ歒�k�`��iH�
S�ظ�]�����
�4҂��P ɡ�GM��O���d�>1"凖y��H�6�Ht��<b�@�F�����i-� JMHp4��+hh}�'���%I���9*�R�Ǒ�+�'`$Lapl�2{F`�$�����8:�'�
�)G7&���b����"���'�Bh�$�-L���XW��-3K޹��'(
��bِl�Z��]���'�z){��E"~S�i<��n:$�$��-^�Kfaр��[I�@&�?LOP⟬I�3�����
O"?;B�`�=\Oj�z�y�&P�z��q�H�4 ���,3��'O^6-2�i>��'QH���C++��RQ�9n{@�i�=�S��?a�#ˋIb�̃"��>3&Q��][�<a!����� b��4&!3���}�<��'m����� i$$	.Qw�<I&���u �����ZG�H�<)�I!s�T|���N�e�n5�@�A�<�Q��zW�����X��9�l�{�<!��Y�6EjL�$�#�4@��M�<q��ؐ!�z��&��L.ND����E�<9�n��ld��M�k:TtkVe�K�<i`��Y��M�*����f�E�<�!C�E8,a�F��~ڀhBD�~�'y�y2�O�Q�D�[a�ȨͲ]��)�p=ш}R�="���č l�PB�K��y#Ϭ<{�H�.֏F�ڤcq���y­@�z8����[�C�H����,z���$�Nوs�ĹCs�����\�	ԉ'���]̓ø'{@ �H�'��az��EvO\��'�hqX�)��Fm{BA�qQ,���'���c'�,ɒ�����pE� ��'~\�sā��pD�`��,;�2���'��p=�3�	�.�cd�͂QS�<pt��R�<�W�\���{p��)ʘ
���M�<1��Σ6�����b�T��K�T�<)��=2?��I�`�F��2�P{�<���N�p+Jc&����XfAG��T���#tkp����a !�s�@E�ȓ_3i��h&)�E�@	�r�����P�I�4iQ�J�N80ab�#�Vm�?A���~r��G����-,���s�<�s��3@P���hػZ��U��Hn��hO1�����d�:i�%��XY���0"ORME���*q���0`�PAw��X�<9�j�3=�P¨�@ �m�k�iX���O���u��Y�h`�&�'gat@A��ZHH<ѐ�����!�*���� �w�<���&SV���je�L���Lu�<)�LB�O�(���_4>_h� %O�h�<��N�F��Q��O�o����b�<��)H":%1�i�49�q8 ŞD�<�� (K`��t��UϚ 1c�y�<� ڐ�RȎH|ҝЕAJ��Ti7"O�����i(8i��Eޯ��8��"O$�@āTG��в.�T�ū1"O� ���1Ÿ$P�.��5c��"OVx��g�� h>xK�΅�a�I�"O�I+s�ʐ
ұ0����Un�"O�)MS�رw��rX��"O��0OG]Zea4LU:o@���'4� 0@m�8�����!I�KJ��7�$D�����Z&"@��25�,0�J(D���p(�%@��PR��>GT8h��$D����mN�ƕ@��� C��ͽ�y"���j����gݖۄd��aӤ���6}>�O���
�6���	� ��n��ȓp��$b�{9R�1o[�R|�Gz�-1��$���LW8�@b�q�4��O֑�tB���8�z!�%>� ��db9D��r��	9�b�C�G��wb:����u�X�'���������I�C+���8\�刁"OB����1N���{�%M�C�.U����8�(O?�	�aG���N�l��ya��*sm�B�I.-f`X���K�\�d�UƂ�L ���"�)���+am֥O��Qg/63`1;��7D�<�P�����D�PD�k1D�؃�'k��2��{:t��q:D�4�Qo���P@@%�H��dK9D�Px�M8Ŧ s�h��v����@`7D�2��¬[�AS��#0���m*��m� V\ə$jΞ~�T|��+^#-�x��џ��?E�M� c�@�3�`R���%�f�H��?Qe�)�'c�B���%ŗu�"�*�
��hNP#	�'��-�PL�<4ꤤ�p�\%Z����'�0Db�ǰX�e�����!�`+fʚ<r�!򤖘,>LQi�k��Zt��j<!�D|`B��-I7r�<�V����`ӜQ���9lV�˔cސx�2�"O��3Vf��*V�(�A�T��@A�D;�S��=��@q�i�[�rty7��^ԤC�	 U��|��2�z��U�41�h듮�댣|�'�z��,Ӈ1�Vt�p�D[?>!�'Ld�b$�"�t0r�JǊa�ꄒ��>I�O.��$�=
2%Hc��.:���'�-y�!��s?ty�`�Y����T�B�D�!��,���R��kݰ�;���G�!�թ{ul�XF��%]ט	*f
A$T�!�$��vd�P�Ib�u�bA�Ap!�d_V� �����na������W!�d[�_���S�cB�^�+�к
�'�������4�h�G�>���i
Ó�(O����ޜ׋���3�n�K�<Q#D�!�<��甂Br|cu�N�<��5�0�ꁩ� ��k���T�<)C��_��H/���f�|�<�P���x�M#BMDZ�L��G�`�<�A0 �%�B��$�4E�^�<QF�+y3(֦A	G�����]�<AVj�rpH���)Vz��2��� $������| X/JMȠ �EM	�dH5D��Pd ݣl����ʍ���uE7D�d�R�ν#h$�Ȃ	��ZI�)D�ȋӨܛQN��rFάgO�a�0D&D�P�2+U�o$��H��7T9f��PC��d��I\?�)V/Z��i�)P� L=����K�<Qrʗ�54@y�@�O45|\�k�"SB�'�ў�g�? � 	B�qo�XyQ�����R"O6yz&&d�'E�/' \�"O���JZ�v�&��r�%<��	�'��mx�cš`�<��ꙇV�V���'f̉�Q��`�hR%��.>_�(Z�'��t��Ĺ?�v�cф�62�j��'���XFDy�`#+A���i�'�)��k�5@��3��@�R��
�'=&̒��74���  �'%�f��'�y��̸6�:���ς:���'fR��	����rbO����'�m����rQ�� d1��$��'$XؕH��Ĉ����/��0�'CD=k��Ш
WR!�#kE&!��a�'@�e�n�<餐HD
+���
�'�B���	/K���&���mQ�Hi�'��x�/�z<���N�m�~���'�yA��2,�����ٛ�z�c�'��e�Х��i��	��ؙ		@Q��'�Y+�<w@*	`s���IFP��'���Mǰ��	
��[i5D�KR�9&������7��u��c5D���k�$8U�6"Q1 ��z3D���&�P0N��� Gh<"&�R�$D����@ՠa�5PP���K��,q׊=D��+V�C.;:9S��:J��Db�d=D��A%��s)�u�f͍�L���D/D�x�Q�ܨ��W�~��@�-D�@QG� HM���\s���8D�$��F@�)u�u��0z��Y�"D��ڣ�R�}��!�i�L�	�vA&D� �5!�[�NI�C�1M`y��9D��R�I�^g��r�@������ �7D�����2/�ʜyƆ�K�j�z3*4D�(c��ǜkP\9����pzua3D�Lyt�[@H` ���G�٫eF,D��#!܄(<5H)@�Ԭ�сE6LO�����m��Ը�ߊ.�B�J�/� ָj-Q�s�4��"O���F�,���ܠh��p�"Ox�Z�ƞ�%{��iv�H�T@e31"Of)���D�.PP�:�쟾~Z$
f"O�P��)]�	��Sv(ހf[��;"OR�9�D�4��`IS�Q�9�d"O��"�g΀s�~Qih�a#��B�"O��@�T�%�P�8��D�Yu�"O@,�f�F�`�~5��c��*��I�$"O�p#���i����;L�:���"Oj�˄nٓ$�$�eB�=H�ܱ��"O,� �*/wI�1��X[7
�c�"O��Bo�ض��E H����	�"O�H��O��F�ȱ8%U$�8��"O*���9*.��1�!cgP$B�"O�Lh��P���c�$�AϒW�O�<�Th���Ą_�a�2�DS�<	T�� s�}�7+�F]�٨�g�<���q��:�Ɯ�<D��hpLJj�<��/A��9����r�#$�X�<a�KV
�8��Pˁ"ņ�:��PT�<�#�E��aP��x� )���Yo�<q�hۼ"�6X2�`����գw��s�<��&O�`��2F�� K������r�<ɳ�Q���h3,�25t����j�<q�V9�,Xc�a���{�Jn�<��R;Q��S�D
@�RH���d�<� �#q	ΖF��h"#D�d�0�"O�P����S/��s" ���u�W"Od�#��8 ��A��)jĻ0"O�q��O�4t���w�� $�Y"OhȒQ.C������
��0����	sܤD��� "Hd>��DB�J̹�7c���y��le��b�NS|��J�-�#Z��8(��8��/�)�'Sph�Q��!:��X�`I범�ȓr�,E�w̜�&ѲEY��D�bk�H9'�Ҵz��Cb�� &B� ��T����F0[�0�4!�:E蔇����}�g�p�8�8	"�0[��*ͺl��f��-f,��B�3DCꔱ+|O*�h���/E�F�X�9?<-!e�I-DhQ�Q P �N�BHL��t���a�@���P���s��ݯ
=2��"O�$av��a��谄/�%u
*��A�'dv�H�L�I��Iz� 9 �4yF����Έa7�[%�$��v�'4  ³$%D��Jf�K���`�t]�7�4R$�V�g����!�J���(���Gt`�'<_,a�y��� R���:�˃B�"@(0Î��>1@�O�Z�z�+����0!��Hu8��W�	� �.�!�� �<�烋��yҡ��@e�s�K)G�����G��hO`�mсC���"*�*��%�1BA� �E@3'�f@��$c9a Qr��҄��x��S4n<%{�.�k��0��ݿ�?��3D�츃��Wp�ݫ�e�5m	45c�.�7%����?S�ڡ��!)����ȓ
7u�a/کLjZ�:$H�&p[F���#����Ħ�A�8HB'E�Z��Ԧ4)F"ԑ>���^�(�c �J�HJ�iRQM@|X�$Ô"�z���!F�>{�^�0�m�Lvn�:w+-hhp��7�����G��q��Ն�	�C�T��F��N� #��׼#<ѡ���������(���&Ń�e���Q�6y�vK�/N�����ݧYYj<uH3����*K��� .�>����P
(������E�Af�ɚ�W�F"�B�
��`=F����nE�jR�0����s��P�"H�A!�Dy)c�	�#* 3sID��e�r� �t�h�B�2�R�J��[5���	�".8Ii�$N�mz�y���Н:Q��:/��;_a|��VyM��b'�48p�tJ�뎧P� ��"��j�娱G
�C��Lj�K�?*���s�F�N8���RH�9W������5)k���� WTp�eP�K{�l)�ɘl\�<0�!��v[�pAI	w��cÉM�N!�C�Z�	�B�	�"~���.�&p���ɋ�p��	*�'^j�uBW��j��z׏ݢ'w��f���q�缣R��b��D�v�3s�
a`�!�u�<q�]x�u8���1����盜A5���g@�R�K!��*u���'y�y�L����'��y��v㌱ �N~&q�
�at���p)��oΔ�mU�F.��X�(�3g���2㪘z�N�$B
#�FKf
-1�����F o�R���H0k����V�H�wW���
��Ĺ�)ݓe�x���_��8��f�(�rb(��\�` p
O,P���^�h�>r�E��
�8�%{��ՠ�(� S�H�+ ��V�:x�7-j�8zM?睝�&D�7J2W���!b%�6C�ɺA���s������ �F[��S�꙲8>|PQ��?	P#$%o>�c�@�������>I�h�Рz!%��WSRtjt�w��n�G��`c��Çm�ҙ��C=<z����� T���,�E�*�#G�.i�P�'|�G��V�j�a���(����{�n��C��/44�c1K>QR`�d�9DDH6O�*��%�G�՛g��!k��Z�xJ�7A@�R��=UT�����yr@D�!qH�3�:�8jv��6CF�B�IǑ{\`�{�aɕ$~Ĩ��i���!�́h��"�� qe�l�T�ޮ�$@�1�E1s �83L>T�3�W/��� pg1O�q���U�(��R��BM��dG�'�l����tH��Ր&'vXHV�ق/RB����5J�XIB�e�z��D�]�~p
�뛐:��@�����Ot���I��mF��cD��ƞ�0Yw�b#�n��i�mP���?>���y�'|Р�S�O�\%����28����O�ZdEBfv c/uB�O���H6��O���/�\aα��i�X���p�m����?c���Q�.@�my���@,�#f�
���d�w#�ؽ*zҨ0/[�?q'B���c��8EOv=�#@�{-t� 0:�O��C�8|6"cߪ6���C�y,�wb�l�k��[�ud s�% �jH(NF�To����~�b )��qB��Ğu[ ��X�b���I�j�T�+�']%&��'�V��6.� G�*i��A$
��@�'��%�d�Ú(5N��6�C� �l�h
�'�p��G+�)z�9���9x��X�	��� 2��/��7t��@�Y�7��y�"O���mX�^+�<1p�lw�-��"O�5��&��̜IX��3GD�J�"OT�	��='�꼂ӭGZ����"O|T�ƅ(tU��B��;o�X��5"O�0 $BڥI*�y1��ǂY�"O���B�g�Z��0��iɜ���"O�9�w�ŝr���'&:��x0C"O��*�b�,`䥻���?4Y�Ab"Ode�s�ȢL��Pb;1V�	[F"O~�`e�_ayT��a|O|Q2@"O�Da�C�.2D\�S@�d.摘�"O�p�`g�X'ʑ����f%, s�"OF�adg�'��#�( C4"$+ "O����O�\�z�q�&�y�Պ�"O�����p�)��f�_���"OtݫQCύot," �XN@E��"O2���HE�xr�p[�5Y4�<9"O�$�j3?��㞯XuU"O���3!�� C�0�B�R ~����"O�р�e�hCp5�Ah	�<����"O|t�E�� H��(5��='��L�"Oz�#X�m-Fy`4ݦ�ޤ��"O�-`t�:&�x�E"�z����"O�U�'B��q�ƍ���� ���b`"O�Q&��oK�X2��fL� 0f"O��`���iþ�r2���o#Y �"Oq�Q�וZ� 0��į:��k$"O޹��i�-
x���"k�~Л�"O�U,\�[��\HuHZJ\0�'"OH9����?e:�a�%@�(i. !:"O�}�Ъ �|�U��NB>*X=�W"OD4��މ}��{RG�<r@\�2"O�x��cϜ.��u��ԇ>�>��Q"O2<���דD_B�31f+���Z�"O�4�a�p���/8D�"OQpd�����h��	3T�	w"O ��'6�Z�CJJ��ˢ"ONdB���|LhX�`Ѵ}�����"O����I�5_�TH����<|ag"O:4y�聭��i4��)�`�q"Ob��T��S�X��W(|�8�6"O܅��m~��h�c�s<�	i�s�<Q�%�1�\�&@�C(�8E��[�<a���F�`��/�yO�� �A�V�<!�#Y�"\�֥/Bƭ`e�D�<3	\�R��x��ˌ"y���"��C�<�`ėi��шP�8f������<)��<"�QB�݇N�0��P�~�<�%�ũ�j��� Z�da��Ow�<�dM�	S�v�!N)()<`B�ms�<i�F��rĴt
G! �<���*�C�R�<Iӫ�c�Ru�͈��I*�N�<YP�I� <� Ήw{*t��`�<!vC�,(�ː���0O)T��HHv7~����
��ŨU,D�x���!J�0xD�W�R`� �+&D�H���ؽ3�l4"sG�/���"DH8D�Hr4�Pl�l� �[�W��葃�6D��K�ϋ�h�p�!��8Œ�2D���J��Dyhr U�'�*C��3D�(+���^ڒ�;�@ٴ/n�(�D2D�����/1f 1#oB6?ܠk�
0D�쪄�*,���$@aT���".D�� �Є`B(H�JYH�O�wj�M��"O���O�^��BRD ���V"O��ʷ�Q_u�fK��2��"O�*��KC>4;�d&"�DД"O����%`��{�mG�h�1�"O���΃�t�~�+C{�0ͱ'"O�i� X�!,8��ɜ�*W�D(�"Oı��I�/U�m�f�E�7I�ܪE"O������<�0!%ݶF0��!"O����G�2�A[�Ğ�f|��"OJ�c�j�%�<�X���0ulJ��"O"5 0)� w�=y����X@����"Oڜ��N���`y��@�:3XИ�"O��Y�G�j�T��̗�S_NEAP"O�EC�kă}�Zܩ��g*�X""O�ĉ 
&�VT(��N#�!c5"O��c��-R���c�:-��XU"O�m�f�7*�Z)3��6ָ8�"O�zʁ�Q�A�B�KDjC"O���� ��&��B�G$SBtM��"O`����8+n�D �*I�\��dȡ"O5����_z�9)��AU�8Ѩ$"O��1�/G�v���@���6_���"O�LH �٘x�]य�I���� "O��3���T�4�M�maU"OpHc�I��#��iq�W�d�R��"O���7�>{�/Q'X�|TZ,Sv�<aыY8�q��+B
2Ԩ�I~�<�aBC�I����6c�%�܈��z�<�6k��jqf���˻a�qH!̆Y�<ɢ��^�9q7�<h���^s�<����@�^�Bc��+��M���ER�<aN8GG5����64t�	�h�[�<c+��i������L�F��ԈG~�<����}h�aZ�J��A�S�x�<1���#�8"#��>]�|8���r�<Q�gx�ṭ��0o�j�B,�u�<�B��_ٸ1�N�	vBݨ1J�H�<��M�I��@��_�����J@�<�aiG�J� @ `��"�F��VmF[�<1CGO�ef�*�%߈<���h�&]U�<Q�h�i�� �"�Z򐸲ˑx�<)��1G�4�c�Nێ��"�M�<��!D��Fd�T�H�R}��T.�K�<!�k'8Z��� ,�
$�{�<#Ɉ����uY�T�x����C�<a��F�N0Ր�KMuD�J��T�<A`%) �IA���p��Ǣ�l�<9�d�W|v�2�i��c��C�����8����f��[̦H�T�_H���7�hL@��$�����CNgم�L���BD
02��c��Vć�3�� G���Q����`Y�P�z܇�cm`��G�ѩf�,��ƪ�*-� ��ȓ.�`��d�>w���s5o���!��p"ؘ��#9����E� �|��1�l%
֎��:��I �Ht���<)�4ڨC���+GBGu�H]��1|,@�k&��	{�ڼ@@T���{���ҢS5�����^j���W�Ԡv�A9V�d�kg혘(h]��Vu�tc2L?:Y�R�Z�
���M��	�c_ ����F�.tQ��:v�8B��@�.�A���̝D����S�? ơ�d"C��Ҧ��E�RbS"O u��P�b(�Å��/���p"O�)C��^TF��13C�@��7"O���d�̛L\��6��?�Q) "O�E���#O'��;�b��<��H��"O��M`f��Y��}s�`W"OJ�� �!S43r���ҁ+�"O@�ʳ�L�J+X,�Ei0up���"O,Ib$��TT(ŨO	U{$!����(��D����TO(l#G�݆>Tx��h�y,�b[�B�XJ��T���yK�1f+JԘ�y���Ŗ ���wTC4�ýs�!��)�!a%�����t(N�fv�	4X`B��wja��쫴�͑s6����	 ���W�.�O���=Ol�H�K="�\x"�[�=�<�%�+D���R�S��D��7�2�J�5�V<��䣀����Pc�-ȳzw yq3�LD�M�"O��r�E�7]*��@*�आ�+���X ��+w�|�����>TxGF⪩�d�@:<��B�ɶL
J���S��Fm��d�?h�:ʓM��C��0=����g3�� ��|���+A��Dx���O�9:th+���pR���$ȸN��4�Ү�D�<)-Ѣ8ߴ�A毞�%:]*�$�@�'@YsHO�no>��#�>�N�W�"¤�Z�C?D���3n��4>t��3n�k�Ȁ3��s��P���=�Bc�"~:D`�#0)�p�4%B�v'np���t�<���O���@����4����"Er�	�Mm2ه�	/f�ҭC"C��z�$���<DC�ɿER4x1�N�b�.��CE4~�C�1���:S���2/P����A�B��k�\�p�G�Q;�9�����+��B�ɀٲ$ R霰}�n�ǋ��~��B�I�bU���2 �V]q����[�B䉪q���	�@3t�!�k_3_�B�	�4��	 ͚tk�T� �7J�B�Ɍrն�p��M}�P:u��~��B�	�!'�\�4���xX���.B��2�h�9�Dk�V\SR`M�'��C�	�~7�@���j�P`H�ǖ�/�C�	0f|`�5BB�\=t���U�=+2C�	/.�v��φ�}J6��4.��*��C�	-,��ڲ��2Q�.�ccN	�N�C�I�V�hX�]�7�9V��f�jC�	丁҅(B/,�Zh��%5�vC�� VR�Ē�kX!,�H�E�.� C�I ��*�`UAK>ڵ	�&C䉏.� ��E��v�b�F�85�^B�əb�X�q����Pa2����fvC�I�C8����&uh����ͧnN�B�	�+0P� $���NxT ���&u"�B䉨B<��L�\� ��hZ?(�B�%H 	)�/Lb��C��),JC�	�iy��B�J�� ���w�1Q�PC�I�:]l��/	8:����29:|C�I4��8q��E:{.jݹ1(�q�B�I�N����*@�tz�a�'�TB��$�,����T�G�D�	2B@��.B�	�x�Ѫ�H�/E�"9Bb�PdB�I�>��`	}�Xx��ϛ`r�B�I��� �wM��_�d��q�����B�ɨL�$ls�
�ԪA�#C��B�	��Z8�#�C8���r�h�˘B�I=@]�d���_D�`J��� C�I G���@� �`؃Dƒ�'C�)� �Rc���L>jT�$BƗq��)s�"O,��sJ�Lq�e	"bÊ���a"O ܐCOA�����۷8a{�"O$IF�� ;$�0% S):1)U"OH�(w�C��Lu�H�{y�e U"O� 3�1
Z����ѿ�����"O��x`U�	�m���ٵG�|Б"O���&!Ѯar�Ɣ�G�\���"O�}�h�a�$���Kz���"O�Qa����b�H��7j�On��t"O�)3F"M%X�� H�=!,24��"O(1�D	��EVB$��ϐ%��Y��"O�Л���y`��RSe�}v�x��"Odx��͎'BYr�k���\3n�h�"O~I!��3���
�dy;xz6"O��RC��R6*5V	�D���A�"O2�k�!��wMބC5'X B~�erg"O��W�?p���g:4[����"O�0�V�A#,�i�1`V,v1��A�"OJ�yA�HGY��;�ғ%D�[ "O�׊��Il�pr!+��S��L�#"O1�%,�0�� �@��l}� "O�y�k�=)8��$��P�8�2c"O��R�=M��B�\���t"O�8&�˧tJ ��"�4[�2 ��"O�5@�,��b�H�&��?m�R�C"O��;��L	\D����[�L��f"O2H4���%���d� ofT�q�"O��ò����L��GN,A�ɉc"O����ӈ9Cf,�t�'9��"OP�ˁ*�	1N�A�wͱ:#dHZ�"O��b�G�A�"�r�B
";X�1�"O���ш�
LV\�'��/%J���"OR��u�Vf��wEȑM,�kR"O�9�m xf�;�N6����"OޑA#@�`bL��C�:�F�[V"Ol���wН�!��$OѠ� "Ot	�m #���8�/��բ�"O�\�#�� �9�`�ݙ�(��"O���(B�\��h��@���T!�"ON��'�< +�9�o]-T�	��"O4�`��
XD��0�eG�ą�"O ��w�
�A��qХ��	C�	� "O�6��1E�B(�+�*3�xSǌ2D�z����J��R���{pL8*�*O��Z%B�<,h9+��ƙ~X��"O�-
�cK�J�H��/E[�e�"O��+�+F^��S�X k^�Q�"OH�blӵe�,ykŭ�	r��Y�0"O��Y�E�Rm u���R��b"O��]�6l�b)C	t��p�a"O�L2B/Ul�,���S�}�(F"O��Q��6a킗��1s��4�"O�ؘ!���I`�m��\��z���"O ŀ�!�$��H��EֵO�rh�!"O���P�˙(��PI�CӻXR��0"O�ىէֶ_�4�;v� E0�ɑ�"O��A�^?$De e�,-r��"O�ȣ�[%jJq��k
���T"O<-ʔ�Xkx�I� $Q��[�"On�0�(ƟXV�Y0� M.N�:�"O��P��� �� v/Ǭo��Ȁ"OTl�H�"��������8��D"Oi
��U�$�d��E�1��<�""O� nq�1�G"~�⭂ü5_x��"O�� �I�*7*:��t &U� 4"O���!��� β�)Fl��i)\�;�"O0�3��,*�4 �Kն����"Oh���H��(�H@ �#s�ʍI�"O��x&� Y�$���J��@"O|�ib�r2�� w �ѩ�"O����.fq< )C�Kd��)R"O��c x���`�lR�s�[�"Oj�I&%D�v���6͐.~�>�*c"O�\P7i��J�J��p��,�$M��"O@��E	G��GT6G���"O2�Y�h�63��w�u�J��"O��'g�1=xp���\�<� P�E"OȼSŎ�y��*g㝸ݶP�@"O�!��iJ�%Z|��򤎹N���A�"OĔIW,#�1��@�\�#�"O��:���?*��ä���G�~�!�"OHrvkG�1�⮚2P`$D�u"O>��L�a�804��8.�("O�͈�m;	�y�#7j�8�1"O�-Ö��;9^��T/�BUY�"O,=Q�A�hrybS�J*: @AcB"O�,@�-�2�Z��\/-LQ�"O����O� #v��y�L#/��Cw"O����Yy�f����ʭo����"O��맯�+	��=�2B�>QL���"O���b�F~}�uK�$_FЬ�A"O�<R���C��K��T9
���I&"Ojȳ�ġ-y�x��	&��4@"Of��u�B�1��%��	���	S&"O��I(�4N���n��_����"O8��TCV�%d �ǎZ�!`P �"O����ϲ��1�kӱ_dL�s"Oܙ �nʌ0�<JAgJxt��G"O���fO���{b`�$&v��R�"Ov��Tދc|����O-wP����"O����dL)OF2$����	V��*�"O�8ېM�f���7L�`C����"O����L����b�5"Op4#�T�:M���&k݇S|Q��"O�E!wER�l3�`��*�2[B����"O�9�uH�Pь�ӕ�]t;��J`"O�}Q� ��!�����X�<K�/�y�#ڇ<P`|���q��S!@��0=��JC;Y��`��ǉ�"�������*�v��	�P��;��c?�)�B�t$�1<���4-S�a2"�	� $<`�|ʫ��� �V� �z�i��)��C&�$C
�(O�OO0�"�	� U:s�0vT�J<�t�,�S�U�N�c��U�L�EEJ9t��'�p�Dy��� L�BIpo�7����lT��	h��ȟ�!H��њ]��t!'�"Mln�	�:��a�4j����TCf�Ow<hĉ�����'0�#=��vzF�i��r�	�`y<p�D�x��PS���O�`�� ��Q��S�o�~9I�O4�����1�VO�s *l�h߯+��6m[��(O�?q���D��A;UjN*Q�5�K'�Ote�; �� j,O�(cZ����-�+�|p�P�#t��sd�Iy��Q<C�ԉ��)��U��j�EB�Fj䝛�D�x	�'���Gy���.B>dih]���I��a���ƕ���ڷ�(O�>�	�܌.	�ℊK>T���z�k`Ӏ������$����cJh�|��W*.��"=��Iٟh
PF��U��y[��P.01bѫ��.�	�X�Q���	�1g�y��{t�:~0(��7�x��Hi���π V�b�O�J�`-�Ģ�(TxY�R�P��)ҧR��],� �(!��[9���l�K#Q�"��	�m��	�U�\I��92#fI�(O���S�"�N"��"���"OO�C�hb��Ӄ�0�S��N�pz�'יx��`b�L�aѪ�'�`7�!��?��'Pn�aQ�Z"&��@����9!��CE����!j
��l��Wդ3��A�������! "O��bT��2�dZ��ӠNd��A�"OL�BoK��Jиw��'L�༹4"O����T(G>�x��d��~�0tC�"O���q Ño�ʌ1��������"Ov�pf̭i� ����Pu��$"Oj�:#�P�aPgaE^���d"O`�"�J>Z4X����<VR�p�"O4h���;� ��u�Hq#�"O�4���C?t���`T�Q�h!��"O�����ͩVӖ�d&�����"OD�*�-	E��\RЅ�=6 �
�"O��fj�VX����R�A�"O���DĢd�^��˾ _�Y�d*Ofu�.S�>�T�E���V��y�'<�Ä��@�U�$ ��.X��'�2�Ò)G�L����� �X��5	�'�|G�6๱��1SC�2�'�ҝ��,��P�<3F��E���B�'B`U�C�1::d��s`P�:��Q��'f�d���Ս'^���D57�ڱ��'��A*�MA�yk̐1���[��)�'d*�qMG�'l���ŰXvrE�
�'e�`{rf��50e����P�mc
�'`�����\�b�0���0b�H�'�~|�b�HI@Pw� �
�'�.0�v��'C��E�'չ��|p�'?�ģ2Ȕ	��L	A�
���'Rq���2Og�l���ī3z
�R�'�(���É���ͻ1.���
�'$���쒀�ހK�* �)c	�'�
U
P�d^��o�|ʜ���'tp�J3�8I�|�đ_�0��
�'��e鄊��h��PPK��dJB��
�'�8��5JO�;���r�Y4(T< 	�'�\U��DE���kؐ�\���'⌁� o{��9�����ڡ�	�'88�a�E�2C�*�B�+��� �'Zm�1F��0BaP
���d���')���Qwl[���;De��*
�'����i��5L�	�珙H6���'OZ]r"L��[�jaɵ�.i_Z
�'��0@��M<��f��e�ֈI�'�8����*9��@3��Q�p�
�'R��3��>4������\W�����'�<�-J�,Ǟ ��ÓO�.�r�'�@X�Iӝq�LQt�y~�S�'<�Ty��\��P��nmp��ʓc�L�)MJ+rB��/Ǳo�Ƒ��κ��삢dZ�#Y�e�,$��e@>y�A��"�4�z�j�&3��ȓ/�l��ccVn�q��#^����dZ�B���>�ı�σFߦɄ�R\:�HɃ7���X��H	zn�$�ȓv�X���蘺C1���"؋gn蜄�b��}�ǡ��WFv�I`��1{���z��z%��hZ<�yQ  P�e��E�u[��A�
�=�e�%�@܄�S�? ��ڳ�9V%d�s�.���\�"O��3�Sk�Eh ��0=��Y���'��'��qh1?X.4����&v�2���',~�#�J]�F��1PaM��|H	�'���ZѠ\44��8�̇�C��'�J�h)A:��� Q� 	̌y�'��(�R$�<�B��U��*즸b�'�>8;6IŎ0�H�p ��Y�LA��'�Ih'�1�H�� *�1�U��'z�pRb$_',����.J餘�'8��'X-!v�}R�	A"�va�'�L�Jc��.D��8`G�r.$�h
�'���r#�Co�KD��]�H���'�j���o�+H�X����O0 Q��'0��+Յװ{"B]�""��h��'��D��)ӏ�*a�������'K����O��B�2����Q�v��'�]�rvxU%�Z	Od��'���SF��x���xѢ�6C����'ݼa�����01*V�P�и��'� 豨�9.���NA�E�ʤ��'	ȋ��A+�*9j��64�&��
�'��(�r�U�n�[r����0�'�P��8x<� � �,,t(�
�'�28�@\�qhV����'ʞM
�'^Q ��
$���HP�׻��iP�'&B��b�'p|` `J�;vv��']"%�%Ä��4�#菥;N|��
�';��AZ�m�FY! oY):���
�' ��J ɦ>�r1  ��,L|�!	�'����Ɯ�s7�88F.�	NԱ	�'�T�8Dć+%���$(_� ��Tx	�'�Je�v��� �i_� ��d��'jc��T�acM(����'X�m��#.�
e�)��%�
�'�$�#���$p���`�^�!R
�'2� �!�a-T��O��>��	�'�츀�'K�+O�mRD��F�
	�'-����.0�Ą����"X(r�'
|�R�Q	q�X���,��@�`�'�9A�+��"X$IiԚ�L��')�(�����3��
��(�'�rL�5aG9G���x�Jͷݦ	��'<�r�n��&�=2k�Z ��'�� �Z,aoN���S�M��'���Jk6x��M�!N�q`�'�&�jg��
A{r�@&Ao���'�}��nP�_�|��R��h$��'x6y�7�~� ���E�yZm��'����3"I�zH�)�"k�-�`�*�'W��J\v��X�	A&<X�'�L���+6�쐴���+�� ��'{H����vW��cɛ�8�� �'���� �c��˕4�<�P�'Qn���ܰ'�������v�����'>�b���+�\�'��Xr�'��eE��$�͎1G�tT3�'r޽�T�"h2X�gnU�v�6a��'&�R*�b�(���_4p
lm�
�'z����f���|X���
e����	�'kNX�j=�ք��A�aaL]��'%P���ᒱ=���㘡ZO�2�'�ʝ�%meɃP�Q�����X�<)�)٫>^f�yc��N������O�<� M�B%و7Ē�yG��n*ճ�"OEQ��&�<��Ε�z9� 8�"O>���À� Լ�s����F �P��"O� H���%�Т�!C@<�"O4�i24
l�Q�υ-����"OH�٧��(}(
(	�,3xȊ���"Oj��7���M"���f7��Б"O&����L-2�v�:e���$��"O҈�j\�U�xY�X�1��qq�"O�`U��,�vAE��
?�B䉶"O���IU99�z�&]�����"O��Y2#H#!3���E�9\�>�Õ"O�\���$j�y�sƔ9s����"OxmR�a-e��]$��ё�"O I�^,�B0�d�^�=�XC�"O����ap���R�R�v��v"O�)��U�"�Xࢁ>T��$q1"OBi󳈘�>��}{t�H�F�Y�"O$�Z�.��IX� �:@x"ORI�AA�� ��ySf/Cx�p"O��*��
�1T��D/û7�� Y�"O4m�b��}��0Q��_�%;��j�"O�ɒ�2P�H����8*16��"O����kˏo�,��(�18���B"O| �D���ܝ2S�� !X��"O��A�ՒFz�`Z�.����0"O:��a/�2x1DѲ���Ft{�"O�<hÄF��Ҍ�gݢXH�"OP���/{�}��
0�4Yzs"O<�����j6 �Q��>8��5K�"O�x�6I�\P�� C�p�!R"O@,��D�4�)�4�c�"O0I�$�P`Z2�0�/'`�~� �"O�u#�d�r����D7�J��"O�	� ͒{dD�%� x,YG"O�C�lY,i��z�O$YfT��b"O���C��G2,C�,C�n��x3�"OT�:䮑�0���X!I�|�d�A"O�Ia1
�$_	��ѡMޣL��,H�"O�h�g)t���i7K��0�w�<��#	�nںY82G�*$PHʒa�U�<9�&ݿ�������o��X��-BR�<�Dfك$2�:��ڌ͊(�ZN�<�NbMA�H�E��W��o�<a��� ���P 	�y�@�h!�k�<��^�M[���a'ua4KQ��n��ȓ	,����[mք����:yr�ȅ��2����1C��Ӣ�̴tϴ��W�Y{�(��Ik#��*�u��p"�s��H/q�qqA�Կ0�f1��9~J	S�B�%̂��BF=\.)��pƤ��# ��c� �B4͏�k��)��n� ��u(@�9����D�6F2�5��'2���- ���5C	y�ȓ:o�)�f	J�+�8\K��/U"z9��?�juq� Y=���	��B33M�H�ȓ :\�f��7_m���à�+H𺈆ȓ �d!��Ε+.O<�0��1;{ba�ȓ74	��?3��#��]_6ҝ��DY������s�0��B	���Ņ��>��R2n�D1�� �H��ȓr?��u7X���%�ÿT��5�ȓp�D�9��!(��c$��#=�X�ȓ2��H�hڕF��(Ɇ�7��A��S�? �m ��]
o���bD�/�>08�"O�8)��kJJ�C4_�=cP"OȘ��o�^�x�&��0TH6u �"O6�уG�9lZز��=�""O�8���ѓE=<0S!]�;�C�"O�5��ރ@�,�`�/c�!34"O29�͐��d�j��5b�ű�"OxDqr���<�(r���U�!��"O���#G�[���b��~<��j�"O�cէ1]��0��P�D����A"O�i��   ��     �  �  R  �*  3  <  UB  �H  O  IU  �[  �a  h  Wn  �t  �z  "�  e�  ��  �  -�  q�  ��  )�  k�  ��  ��  ��  �  ��  b�  R�  ��  ��  �  j�   Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�� |d��"O
`�(�;���8���-0��1%"Oj4��ND^[��"3/9�0|H�"OB���H��*�ʞRy=a"O�味V�!X��!&F�:J�$���"O,��a
���C�Ą�M�"O,$3%o�-���p���+Ն�:1"O��ݢ1����`���y14]2��i�<�6��{_���c�H�`�fX�$Kn�<��A̼VI�xR[�)�Ć�pඤ�ȓA5��('nߡ4�� �)˩%� ���,��r�؊b#`T�eT09���ȓ!�b��g��}�8�F��-? �ȓ
K|m�ș�VṔ���2�%�ȓ"R�X�j�4JN�1�˘X�i����̹	_�jZ��1!g��zܶ��ȓgil,*�J�
j�Ne��i�J%b���f	�(U��:���G��$Y^م�~r�� S�%T"���k\�jx�ȓ|4�1�îJb��@ӵ�ݩn�V��/[`�"�v4�R�!ʎ<��M�ȓ`:��z�ؚh�J�Z��$HY:	��H��p�m�C1��!��B:��0��EnjZA V;9����J[
2���	��4'J�EA�IVW&��~�(aZ��ӹ�>� o�Y�|�ȓ�f�A�
Ο7�H��M�$�����mޠP����/���ANXo*�ȓTv�����{ ��-7�*h��I��sB�8�8���3����ȓNe*M�悡;������X�o��!�ȓ'lj�#F�m�+R&;�|��2)n�C��0S4���T:
b���:�0!��e֊��)��ͷV��,�ȓ0�&�8#���� ع�L�����;�P�AFd���,w�6d��r�EQ�( �gVlɦ�M,H��,DP���|�I	$G#\���ȓ"�)���E�B	yt&B�^�LɅ�4�� ��eëF�ڙ��n��R�p�ȓp`@}bŇ�=�$�AUN��P����L��p���_�a�)�Y�!��-��u�5���o}�`iF�@A�p �'�ў"|
 զFz��#���4����jIm�<!�M_(R�����(�M���Âdæ�hO?牊)Π|�7b[w�j �F�' C�	( y:��6j��U-Йh��� �'�"o��Fkν���;�L5c�a���O�6m�>)H|:��<"W���M������zھC䉫a�.�Z��ީ������'�C��Y�±	�b���8����C䉈?���.�64M�T*�b���>�'a}R	�|g
�{�@�HKΘ�Ԍù�y�j�4��ᚣ�K+$XLcW�P��y� U2O0TY��G�:y��r�牃�y�[6~�@)��*q8��p��y�*P:u���7���3e,��G��p?ѩO&��@C ����ժ2l�x :�"O>)�s�)h��ޭ:�����Oh"~zGm�	 ��X��T�3:�4����I�<�uBÿ`�ذ+w!�kR]qO���t���F۷R�@ ˶��?&�ߎb��ϓ��4��� y:�I�?fp�-IbYa�4]1"Od��Q�M�w@*�`D�'����7O��� �yY��n~��������I+o�8�ŕ\Z@�9&�U=Zz�B�ɮ	Sv-���/~X�{���
V	�d�<a��T�'��>�OB��0ƒ�7�4L��R.O&���6O��@)_"D|��U �|��!H`W!�ĕtyPL�7�#/�t�dʉ�U�a��Of�[���.�>���Z�2j:$�s"O������j͘�Z�/��Ht��0"O�"F�h.B岔D�Pv�lBQ"OH]���پ�YS툲jo��"ON�
�*5�p�B�bV�	f0;��'�P�H����l@�в�h��<	�r�Ez��'edeJGj�#)Θ���k���)��d+�'g�z�3��9��$ Gf�
I�4,&���D�ˠ�2&�R&֡	��C䉂tkj��e��]i�QB�����C�I�A�@4{f%L.���gR0 ?�C䉹r�4��&�4e�JT{u%</�@C�	���-4k4R�s�$O�G�ZB�I�S�,8��488���Z��0B�	�(%Ia晇&�9"�B";�B䉔g���rhC%�4�ȴ�PA�B�I$]�
�;GGDy2,�W��V.�B�	<N�-�c��2A�XE����1P�B�	�Y> �иi�������lB�I�q�!��$I�@���V��IN^B�ɨgX�x������Wa@�$\,B�	�W�xW/%T"��w�Ҥ18B�I �����Nˊ����2Q:C�	��.������ES�O	g�JC��#�Be+�N��y��s�
!�:C�	t�4U�"���~Y"Ģ0NG�"� C��(%�H��	I'g �������*C�	 N�:,*��\��:)�3U�DC�I>[T�0�e�O�]~�q�TeH�
�xB�	(n�\`*��M�����3��K�vB�	`̓%� �H��a��G%�tB�ɔ~"1�,Z��@BE,��C�ɡWR�0�@�
:�U��_w�|B�I;.ր4��M��G�|��W,;W�NB�	1T���a�PH[�FɐBf
C�	e�x=Zd��e=J���
,D(�C�IR��4�S�v&�,�Mr�C䉪��!d��7:�F|�7��k��C䉣c2��W��r�<�`�X<�C�I�2�u����moL!@Y$V�lC䉌~zf$r��ǃ���'��	�d"O4԰�	i�ݑeZIT�j�"O�,����&]1X�!E��z.)+�"O{"n@N����h�r@��"O��1�	@�*r`��"X���0"O����-F�h�B�i3�W�?E�A*�"O��P���C�X8�d�)[np�"O���E�F(T)��P��F:PH�a��"O��a�)(�Nx��Z+QCz� "Op�)�� �	|��!gN �*;�	�V"O�0:�����Z ��C3!����"O24�����k�]�6��S$�p�"O�1��#�J�B�ɦ#Y���a"O��$ )�1Q��%*��c"O����p�V�kDI;M�.�a��l�<�c�٦$�����ɟ�Z>0�j�<��B6u��$�F���S.�5�fLo�<� �}z
�Զ�ا�S�T�s"OQ�5�K�$��Q�4�"ڸ�97"O�P;�`c�¹��O-E�����"O��B�/	�qS��a��O_��%��"O0��N�`#@�$l۾_{�X(�"O@�s��WL�#"�/Rs|!�"O8�C���ha�-�׻g|ms�"O.i�B�S���!���P^�R�"O���Ӭ9�ڡr��J�H^�"O(�QD&�#d�
��Eȫ5W���"O����`S-9�8�lڌa�y��"OVy�T��25�<H@c̚�t}�8��"O(bŉ�&�4�i�sȨ�y��~�:\��$���f�S���y�`Q&\t�	U�ˁO�2�[rD���y"�˻,�ra^�K���1�cÓ�yRD�"H��Y��5<����NO�yr�Q�i�4��0.��4� �����y"�I�q2�����+��t��%X��y���m��l����8�����I�yre�K�0)�AHN"��0r�����yr��>�Hh��[�e���EAZ��y2�Μs��cv�sz�tk�$���y����+}4�{W�I?k���	B�C��y�BғЩqwa �W���B��[��y�(V&]a D����%a��(�0�R��y"cĉ"S�T��ڵ"nȽ���\��y��Vd�h���ǩ�n	��@B��y�aG ~�����p��aլ�&�y��U�d�Rqg)��"��4� �y"D�T�)�c
M��B싳fҒ�y" T�CX��-\I�ڭ`�o�5�yrG<%?±[%8�� Y��ȼ�y���>.�*u-�#	�Z!k�R�yRE�9Ć-��E�v����1�ybg�S�QF�x��?�y2LK������h0rZuq�@��y�C�^��i���\�g?��Q0�C��yr�Y)�:4�D�+_�c �/�y'Ǔ)Xv�ӊ��&��kW�ӂ�y�����M2��[�oU���ȑ��y"��<[��@��{V4`;��Ԣ�yR�ܙ\
��2?5.�%C;�y4$o`���BB<Ŋ�Y���y�-�pq2%*D�!/�Zq�甭�y2Oߦp������(0�.1��*��y�����eI�D�<����	��y���1R_Bڣ�(<:n�� � �yb̂�x�2,շ9�m[��X��yR���P��1Q�'�.���SAc���yүG?fV���NY�TX3%\��yr�H+"*��1Z�R��JS��y�hU�m��$��9�ne�2�W��yb�K�gD3k
-AzI�b��"�y�� U��4�ͼO�pH��B3�yB�*u�X%�A�v������y�/�	j��x!w>�q�1*�yR`��	��B�ܝpF���S��y��D�D����n`�x�Sh2�yR��8���j�c�X�[�yb��v�󷃎��<hWL�y"#�3J�����԰$LQ�V!�y"�M�	�0�8��|�8i�"H��y��##4�kF`�o�ꕋ� ��y
� ��`%Ͻh�8�s�"�n(���"OdJ��/4�������	
�a�"O(�*�?tLhA���Ӕ]��"O��㴬�;4LyGm3d0��"O�� 2�ȾF4N�`,K�l������'��'���'���'*��'���'4X�r�;.���a1�.5a"$3��'�r�'�R�'F�'���'2�'���E$\�e�%�6wj��A�'6B�'xB�'���'�"�'v��')�E���$#��I�`�ehb� �'��'r�'��'�2�'~��'��,C���&:���!�ڛIE|�9P�'�2�'!�'Z��'�R�'b�'��$�&�[�{d�9�Eܛ7/��Y��'�b�'B�'���'��'{�'�(��g.� n�x�Dd��reL�h��'���'�'���'�"�'o�'��I#��*�^�2������
#��'-��'���'%b�'�r�'��b^$�,����_$P�Ѕ	J@�'���'Xr�'���'�r�'J�h	�
IرYT�H�%���$� 
b�'���'H��'S2�'3r�' ��K�DK�$V���S%
��%��xs���?����?q���?���?����?!��:5��qr��"ڌP��N�(Ƽ�����?����?����?����?a���?���/�D��M��k���C�°	T���?Q��?���?9���?V�i���'@^� ġ�w. (z��=��M�ʥ<	���󙟤iش[:ܒ�ƞ�{��6��+f��A��l~�AgӚ�$%�4��DkӴ�Ƀ�οZp�6!�#R���I'E�ۦ��	 |a4�l�i~��_�;�3R@�e�I ��;0��=��8
7�O<1O��Į<���I��r�����L<&8`Pu�(� oZ��c�,�X�S��Mϻn��ɚDm�*��Qy�0d�ܝ���'՛4O��S�ӑt�~�o��<Q`�-�.�B���)��
`���<	��>j�	���*�hO�i�O
J7h�9�F@� ��j8�"41O�ʓ��Ǜ6R���'e�t�R��4ᰐ�N�#�y�C�'��' ˓�?y�4�y"Y�ۑ�A�(��,x��Ʋ<�&�0?��"4��'-
o̧!���)_w���$
g������4Y�0Ph��G! ����O?�I2�ʹ�0��Yy�T�U�ڴmv��I
�MS!k�V~�o�P�d%�4�`e�s��,/�T�7�ΐ^�X�i��Od��z���D��HL67�%?�3��|l�|�թ�Jۊ���
L�D�K���9fǴq�
�f��I$�n�E��|��� �J-qt�A�T$H�䮑��yb�^2n��D�qN80t�8���?o�	�Ƌ��� �@�U�-$�HP�g�5~��ȸ �$Ux��	#W��CGƁ�C�䌫ĩ�^�V��s�/L���g���|���J��ǉ1�F�b����o�T�jF�	�J�l���%P �[�.R�F
��k�L�k�����^ Z��ͨ7���(�k�*Ȑ�M���?1��ڥ�����K =H h�T&}/P�ȶHvӺ���O�m;��O�O�I�O���������^ɹ�����ഺi�(�Q�{���$�O4���:t'�t�	�GߊH�ÈL��L}����)���9�4%ԍ����S�'�?���{}~`��ޣ[ �$�Q��4RU��i�b�';�C+mA�Op���O���8~zvy�O@�3 �P`cM������?)�d��xy-O��D�O��$����IF�E@�w$	�c��	psè>ag䈼��<a�S��'�d�X�!i��:��׈DH�%y��>!q	�(@����?����?q���?��Ȑ2p/����l�q�5�D9�W"�*����O��$�O�O���Oh��U�ܟ,D�0#�s�v��-	62 2�����	����\�ɱr�����{]���9X�ZuSƣѹ��mZ��H�	�t&�L�I��bC�R/_D7�p�T��-������(e�"���]�L�	����IƟ|���Cb�@���p�Y��`�-�ˠ�B՞g���n���%���ꟴ�`Bދ!��Oh$+`�c�u,D�H�հ4 ��M���?�*O��a�]E��͟��S*hT;$�S9(!BL���N:6���H<���?)#�AR����_�I�hF�[8Z7v�X�%Ж'˛��'�,���r�'-�'����'fZc-ԩ�N��GL@=H0oR�n�(�ݴ�?��r�Hͳ&��z�S�',�0-��`�#,`R�C���f��lzA'�����	zy�O�B�'��	�^j��GP @,�qg*�-��=��4*�~8S��Wz�S�OF�D\,D�M 7|Iwꅹ8x0�4�?!��?���G �?I���i�O8�ə�򒋅
E��Q'��25��`�y2�Ǟ7&�N���O�$ÝhrQ53x>x�®��Jk6�o�H2W/����?�������%	�����n��@�H@�� �1��E݌�'2�'$�^�P�IV����sBV%Z���N&V����XRy2�'X���9O��\��P�4�`���J^����������'�2�'�R� `�/U���,���ᘁn��H�iC���d�O~�D�O���?���gB��O#\�kP��� �d �*.��,i�O�9gV�?9��'')���$�'e�H)��V�YeZ֡��"��ȓb*.���nZ���	_{^���'��=`�)֤L���0Be:�X����Z=*D�A0�@�~��)X�AJ6�Ł�]���	8\�<|�㣖�K&��"Տ�vP�vI�<2*BZ���K5z�x��.p��� -�ԯ-ɤ�H	����4�҇u����U�I�`�8S��1O���m�i6Nŉ�l�ΟD���K�BK�[��8�!K�[r\C��B�=@p�5B4jzD�V'�/�.�|b>����'m�]%���T�-�2 �P ���
!���h��q�O>�����`�ܳ�+V;w�h@b�˺n�@��'�⛟��,��<�D$�,R��Z�5@܄(#3d{���	hx���'��,r��C:;���b!=�o����'g�0���l��;, �����*�b�����?�.M�������?���?��P?���_��!��⇕++�8�Eb�EH. ���eA���`A�lV��YG¯?�=�q)�H�:��g�&91�.Q*p`@S��,�<�D(�3�1��O������#\�©0¨ؼS���-mZdhW�*��88A���?�eƁ�?a���?�gy�'G�	��fD��/.n	z��D%��B�	�:IbL�P �PJB)���x�R��D�|�,O��F`
ݦr���A�@�J��%���,���ȟ���ޟ0	�J�؟��	ן�I7� ���<�X,����R��_�$�1d�Ȃ*.���)�������مf`p٧�K�i2 �'��V.}��M�${�+�+M��Dy&�R,H��8؁�ɖ;���ܦ���ҼҜ��b�k�t|�R��M����d�O���ٟ�1q�>4֔�y׌M!NYT�5�#O��=a�'�jf`'��"�|�����<��i6��<A���3�6�'oR^>݂C$��q�mꔫ=F�@ ��ь,�I���P����Q�ӅթK\��fM�u���a���pF�8�)�7
��`��@;J�D<!��#�3�x@�/��:��p��@�}��(bAΕ4�"\��E�/&~�e'��T����'#ʓh}2�����M�4�i�RR>�0a��	���ZGC$2����k]͟��?E��'�h��Qc�I��
��E�s1v�Ўy��I-�M+�i��L��J�"qr��>jy�سV�[�y��"�X���'��]>5 �	ݟ�������"*�|,�Jٟz5��Ě94���(C�P�J!�Q�Y�n>v!�������.�e���ˁ�OЀ��e+��=�r4Y#A�"�����բmزh�`,��5
x̲�l-���.҃�]�JY`]_q�Jq�#��K��`B�w�6w��D2�� S��F0kVݱ3,q;���#�O��d�Op�ľ<�����O���CeȈ1`���ݕ%T
�؋y��'�<6m���i%� )�a��?	�gi Y�ǏڜC�|�s*X��<�I<�ԭ��J�ß�	ϟ����u7�'��,��+o8;�CWPM50�"Q�
���&�+^tמr-�h;�x>#>鐭�1���v�� ��9��e3>��6MU�,��S�4$�T�p��hO�a�w�$*���DA�^��i�O.L��O�O���]���<����?���k2���2��t�ƹ�Q�U2�|��'�<e�b(/��8�eo�Z��<ɢ)lӼn�|��?]��]y����>7m-��Y둮3��-:H��;G����O��D�Oy`1�O����O�aSN�r4�r�� @	��[{�z�k�hI�{��aG]Yx��"�N�'An����L�0.�� ��j|t*d�[.c��H��d*\�B��Bz]�c�D�?��'6ҝ��d,2gV��7��4!|�1��Ӗ���<���?iH>�'�?�D_�mr� ��gL��2<.m��C�ɳc�6]{�`8>K|�c.B�t�-�I5�M;��ip�j|���T�����Iϟ�iޡR�Gߌ΄9!�iE�_��2�4$����ПT���2��7��({�b����*�<�-�� �b��=�%V�H=���	ߛ��,$B���,$@2�]
n{��0c��G��Ḗ�A���҈��1�0YDJ�"RWv��'g�aj���?O~������'�Y�.����V2jވ���������$�����\�	)\�z��?�a|e+��t>P��fɯD�F@A�g��Y��$Ԙ k��n�ȟ ��L�t�_�b/��'w2��	S�h�hԤ\����lK�{#��ã�L���'�T=�dX��d�~
����z�,x���A^����!S�`�g�Lƴ�c�Q�?����cE,M�,�!ı�x�96F3t|J����}��шQ���'�Λ�v�jf��m������X+O�Oc��R��3��"�-�P �5��8G�;D��(猚U���!��Y�=�a��%s|��`��O^�+��+3l =B�D�;?�Нy`��O��d�\�+���O����O�D���S��?��bJ�D�����
Ǧ,�Ѐ��A�^[��J�n�5<���k��@1Y�g�'֞�5�߻Yz��p���g��Ti`mW=dF���5�wI6aQ�����P��O ��v)�X��c�ܣ.= ��%�OfP遥�O0n�M�gy��'Z剓_d�c�C\�����Ʌ�>��B�	ҟX:UOH8l�]���_) �
��I�HO�J&�O�ʓ =~X�d���QRB�u*B��+bZ1/�?a���?���Wڔ�(���?9�Og��C��9eԈ9ElG8+"H�A�D�d�5��d��0��-,O�uk7mT�P�Y&Wg��1A�	<x���DE�b-F�x6�F�* ZD�/j�� Հ�Q��ɩ$^���O����!I��j��v�ĀI��O���<�������� |x e�`�(dK`۝Z9!�$S	:��p7�ɖ'�>E)D% ]%�D�?x3��d�<�-����Oz���|� @i3��0�<�UN�R'���am �$�O����(o �^�`��޴��p�OjZ�;"FݒK�$p�1�� d `я�dȎM�S0`�ɦ��SD�!l�	��A�B4<�`�$��6`�@^
�p����=��}�I%�M�G��d�'$ %���\ �V�#P�
c[�$�'��O?�ɚq��!y�aI�&:�I�.��~�T�hO�)�m�ɐ	��X'��G�u�r�T�NMx�ɴ%�Jqش�?Y���iRߢ���OF��?+'�m��gK�z2�}�%��h�"!$�+x7~4�$��k��h��|Ҋ��bzFԨgB��X�"�B���*h��$#�#
JRt	�f��\@z��R��6���w��c>�������D�<�p�B���P���OjQm%���Oe>��Fk����B�` ����������OL��K�u�2-����80X�y��J"L�1OT��]�'e���'��c�ę\,��p��)���6O���H�H�\�`R -x��@"OT�v"K�Sֺ��i�Ep@�"O`��aa��?J08;�E�!�&���"O�qٴ�:Wdp�J���$�4��"OFI0���z��լ�3s��c"O0@�)�",Ϟ1�i˴Hof�cB"O ���E�-F	�%"ڃ!YZ4�"Or9�Ee&>��#T]4s�t�0"O(�p�%'-S��[A�G�&}RY�D"O<�ڱIӈ(BA���XnP�e"O�a�F#F��ʈ���q�P�ڧ"O�`c�&�L�h���� ��K""OZĊB�ګ,����kK7A�$5s�"Ov鳬�P��������	UT5�q"O��:񋛻g�$�0�N0 -\ZF"O�}���A�E\�UE�@K�\�"Od�r���t��т�,vt�-)C"O�����
y���^i��7"O��� �I�CqN�Р�H�{,��K�"O襘f�ċb����@�ǉ�,��"O�Y�eTY�5���
#����"O�<���
�z�!
�Ǎ/m �j"OJdX�n
�Gmp
��z���z�"Ojuˑ�M`�<Qc@���-�^�{�"Oa�2�Ɋv�6*���	��Uٗ"O�5RC(+�xH�5�ɿBK��r"Oԉ	�h�>���%�J<��"O��H`6n����k�5�T`�"O����)] /}�A���^B� ءp"O��t���J��:��(Z�Zq�r"O�JЈń�����&4l��c@"O��*R@U)F��8]^�r�[�b�T�S�jD�:P�����h���S!��@���1�����u!��H4x!��*-)�`���)U����@�D�X�-�5,���3��'?���a);Q�f�e�'1OZeZۓ ?� �Y�k~E9Ck��T||�nK�e@��qv��7bJ�*�'
���w� .4l�ˑHX�TR�:�}�!š+�)��CΝC8pѲ����X-�D*��_$�Q	�sA!�9o
]ŎS
�I�7�88����5PpP�:�h�4�?qu�>ICcɢv0��aw�� d�z���d^�<ADa �M�fڠ��)�丛��Yݦ"��̬�YA7͎<7��1��I�b�,8I �W�8��a���M k�����L�Աd%��lEpX�r �?*��X7DU'�$��%k��B�ɟt,buI�&�3Y"�hj�i�8��b�`��� g�Ұ��-�`Od��}ڷ��0������G/���d�P�<Y�� �3�q��կ`r�r�ʕ�5Y
��4�	�^�\�$�
(\H'?���xr�V,<u�E�d��B��Y���G�?I�H����y�I
E��lA�IGY�J(��,�W��R`�6Tt�!��"�p<D%P^�>00�oY,*���u� t�'�P�?KbP@�O�k���޴1W�-��`�}��@L�S�&�w,��ʐ�E�8��1-�-r����,�>�aܯ)�l�!CU�&��a@�B?�}Jg	�;9	�r��q��2��D��HJc��? �hc���S��)�. ���S�Г^��O��I=��j#�ǹ! ����\�=�;��E�'���d�+�&ȹ%(��4�* ��a�V�T�3IT�B�B}#D�I%Dv4��b¢*�&�HU�DH?��G#~y"�9�J�%@`ʵ�h}A�j�-�@�eO@�ū��HO�ȅ!ԬiD�L�љV� �W�L!Fl�� εx� |l�D}r�G�/�2�@��<G4�C�L֐5g|���&�.$Y��>q I#�Nv�9h2k/X�Ȍ��LT��ųd�����=Aa6�^��lS8�ڀ ӆ�*tAT��d�I`?C���Sņ��W�v����W���gB.��B�Lw�'^q�T;�r�*��"|�HqڴQ�@�С�F	|�0�
 lK$��'w���IA� l��o@�ҥ�V)<M0�$d[!dp��	7{�t(c$��Đ�y�.OH�r�c���"�d߳5��A ����}�:�GzB �$V��
��Q�k��8���ר0D�Ie-�04�@�#j:��	E�D�'��5�U��%���˻,����L3U�I�T�?LOx͉q��83����*jA��)�&��a���X�$���&2|O�I�1G+@���ݗf~4 
4�P)]�E~r��6P�>4�X�A�J� �  %��͝��=he�@<�x�ɰ�)�/n�Z��Q�*��+\�=̀dlZ*%�P@2i��q���X��I��˓QF��gI�Z���B�%z��Mcm�x����I�H?�u���R�`�CQ�Z�x$%K�I}R�=z����+�L�RC@��HOV����5C�A��U�1WX�l�j^0�R7L�;T��Du�� V�����ܻ!����s$��
O:A�&��0zμv#
�xǂ���I'^����G-���)��5�-xS�U�o>Ls�q�������g�΍�,�A�=��'��n�ZɃ��S��Aa��ӏ<���i!�3c���@��!QTq 
�*{^�L��9�Jw��F��#pT��6mʐTOHD��8�̐؄헎Gd|P��
A�ؽ�>��'��#��]�����4`�M�Z ���-�<��"M����ɾ~�l�����5)R$�Z�.\@"=��M��~l��á�lr��3/MN}��8N�HeY���9�r��"�I�>7������I�@��/�^�w�*�(H{�����ēyL<mT��*!4f�a�(׫ʲŘ���6 U��$v�1��.-�EH�� �V�i �i�i��27O1��&��-.%���ܸl�������j{���d_:)�*]���0,�d���	&<�rD'�j�N	��@�9`�d�C����I�E�@je!O�S��Qh�(p��,��BK���ء�P��~A���g��x��D��_|��k�`O�n&!3ဝ'�Px��{�PqQ���}��C�9����� T����_*Θ�GKҝM�����X��Y;���*$���Y�8�!��аtn4���޼8儵BG��	E�V�)��̉��T8K���TFHK�|.��'m��V�by,x�����$#��IӒ	$=B�x�B�a_!�"iG�Q�⊶o��]*5DUZ!�$ĽatJ0y'����6����H!��r?��:1��3	�v��4I<!��ږ&�t8��m�|B9��.\!��3�PDP"�˂y��t!Q��1WS!�$Y��F��q�\�c�F0�PB�- !�["Ad 3$]�-��,���̆1!�$�
s��h��02� �a�!�<?!�D������b_�E4y� �o�!�$��_�(kq�[%:�)݆%u!���l^�����9���h�c�!�D�)'�z=�P�� � x�UMF�|�!�$_x�F��b�2}���:��Ӻ]6!�+I���wF�p�"�@�I�4!���(;�<82���u�@�k��+!򄅨SX�����~��qPK�n�!��,QI$�BƍJ[������
�!�D�=��!�Ɩ>�D��щLY�!�d�B"����]q�Ȱ�nܕI�!��[�e��%����'R���@5P�!��3"cf����F�p~X�y#��)�!�DO$W���Y��8d�$�ԤJ!��C�r�
����"{el�H�J�J9!�Qs��	��Yi��	se�	V!!�Ą8{2��2%C�'x_��[����!��4r���iP!@�qU䆖j.!�� 1�� �8Xb1rWl�u*����"OB� 3�'5���HC�Y%���"O��PO�&Ba�y��C(@�"O4�c匐����3E�O�-Pg"OLu���!7\��ً�hM��"O�A�W��{�Č��̟�t�hӶ"O�L��U,Fm�C �;n��x�"O��@���Å+/3�PT"O�LZ��_=3c|a�C5B;5"O��SS�ч`�Xes7�(aiP"O��b���t���J��+�D��E"O.]��%Y��8�3giۨZ7��3�"Oб{����1�d@�g�9)����"O�	�O4�0�H����Z̢0"O�va�GN��/ʣ'���"O���MU5[� ��C�Fg� �a"OX��G�=A�b����	�w}b�@�"OƝ��lA�?{м�I�:g�- �"Oʕ�$��?,���&�2X7b}��"O��@ܚU:\ܱ��x1���"OtȠÍK�^��Q���$���`"OX��c��wX�����Y&�0:�"O�����M>��3C���"On�P��J�)V��҇ҾBJ(2�"O�07�8 �PJE��;z� �Q"O9���(WLa����V|A�"Ǒ"����$O؍6����f"O�z5b�
�0 ���o���7"O8��#�r��1S�4���G"OVA�SbW�p(��!�Zj���3"O(5��Y�aH����A�0t��A"O�Z�0�e�K�p�(T0���\!�䀋l�h�B�%@
~ā��J�!�d� .��L��N���Z�r��+=�!�D�x�E� ��2����V)	4z!�d��z;��L	��|����5�!�H�%S�u�TND����W'��/�!�DB[��EB��
a1�0F'�;ji!��^垽�F���.0��``E§L�!򤃜`,X�����Id��b�U6�!�$��@�0� �߶ق��Ej!�$�91o hV�Ԡ9d���2m1!�K�0���㕾c�4�眼8-!�$F�6Xpu���%��)�̀�u"!�$�)\e�7F�/��Q�r	�V�!�DB�x�N���;o�t`� OM4"�!��O�a�ZT; �&Y���fdߧn!�d��ה�{х�������V+5�!��6p�Y1i!Z1�#H!�$ȥ!���9 ��h8N��_2>�!��"~~�ɲgQ�8:iX��
�GC!��(������批c�Þ�C䉰>�r,���N�SJ��6J�,z�B�4,�(� ���z�ۄi��>B�I+���:�d�^#0�>B�I *�XP��*SG�}�^	s*B�	��r�أ̆���̫����^B�,���8�cG.1��<�1cZ��FB䉌@�B�� �ǳ�4����@�B�I�gs��5e�C�vh�S�T�UXZC��?B��P[�n
� gT��X�MK^B�P\��Ӏ	*e~(d1F W�V�2B�ɷh�z$��d5 ���a��U�"b0B�I8t��5��<z�!�@�[P�C�)� >-Z�-.�|A`��8�J��t"O
 �4��>�މ
�Nڼ(?��+�"OT��T�!% P�+Z/a(4�"O,�;��;{�@Rd��D�셛T"OBi���E���cR�<��`"O��@"��7!�%�eA��7�l10"Oe� eǜH�h�h4Ό�-e`�� "O��TEG)*� �Y�,
�`�z(��"O��yՋ�^�������[ʢE"�"O�%*�ƟAK�D��#�9���"O�15��"u�H��^pe�ѩf"OX1���v
 qZ�i��)ęؔ"Ol��P�x/�D�%�P�n�F��"OД�Iɀw@�vL4PTJ�"O$�ȗA�T;�}˷ˆ�_�I�P"O.�R���#�hJrK׺Q ���"O�`�����/>��q3
ʕG�R9�4"O=:%N��H�4��ш�P�(Q�V"O�`P.ތt����Rg�3"On*G�C	�@[��Գ(���Pd"O�X��a�nP@!N�������"OJѸ� D�Ȁ��L�j(��"O�iٲn�P�zVZ��<�D�S!�y�+�+l�������2N����Tϔ6�y¡_�:j]�UZ,3J���y��"+�DH4$^�T&��K��Ň�y� �_~1��,Y�M0�e���y��L�\KИ�ℰF�Yx&����y"����`�H1��g�0���(�y������#�I�a�h�2��y2�ۈG��p(����m//�yB��@\$Hr 	׳9��"a�y��):R�1�ǋ
��E	��1�y2�.i\���ݓ,J1x%e
�yB�@���i�n�{�r���L��y�&�8%qf�qS\����C/J&�y"A�|�a{�-�K��Q��f
	�y���3D���r1���F9f����] �yB�ծ8Rmh��נ(ڄ(��J �y!�!n<���鉗(h��B@)�y� 3����!M�R_<�8�J8�y"$~)��3q���EV|@�1���yₗ{�2hQ�=6<�yi����y҅�%6����#_�y���:Qi�7�yR���h�#Dq���U���y2��&Ƕ ��*a�X�A`MD��y�̀!d�rl��L'd|�HT�y�f��dѶ�bcJ�Y��u�����y��3e�ykc�	�R�)�"�A�yʒ(,�`�J�K@�Lƀc�̴��d�����'�J<Q���QøT�i�!r�i�'RF�`��EC���c^@X�
�'DY��n�(��he�(_���!����B���I�^F���'E�U\�`�Չ�1�!�D���P��	T�x�jǃW�M!�Ą�F�����PjB�]�(!�M
W'ԑk���D��u ȉ
G!�d�^ӄ�E3@XvL�g��F�!�$0=R>Ÿj�6/KZ�gȋmj!�Q���A�[�����&U!�� C+Z	�"K�i� I;aK�<�!��/��y'��4��q�0�^�!��Xzu^��p�P^p�C���P�!�d$�T�K�h�'7a&i�@�U�!�� ���$B#9�}Jŗ���"O4��`�2.�-*e��?��4h1"O@
6���,�ıhDdޡ�����ID>�{��R> �Jɂ�(چg�>����?D��)R��/?���C��4a�(�q�2D����d��M(]k�4>=dT�dn/D���p)�8���pV&�5>���Ԭ.D���6*�$�*��j�+�*��+D�h���JRL��t�Ý�؀�W)D������7�a� ʁ&3��B��(T�4�E+�<WA���r�_�_\��6"O��F��O�U�n�Q�8�6Q��D{���,S@,�����hE�V�R�!���)���s��"rQ栱��R- �!��#x���C2%��� ��- x!��YD'*l��T� �ƈ�#�Ȑj�!�$�)!J�5k�a��J}��e��&y��	S��<ɉ��'J\�"��ܗCȚUs ��4����"Oi1�&�-f��!��ȑ-�n�C�^�XD{��	��a-�����/_2�p�eƀ0q�!��9!B�gbW6=#Ac��]�4�!�ћ}����9��j�#X�;�a~[�4Y4�	,vtX����"��r�6D�D�B.j�P�y�(P�D5r�3D��x3E�Z۸�J3FO�X��.2D��[�����`b���?[�`���1D���'*	
;��\�6�[��0뤬2D�k�/ o��[d%
�O�H����/D���mJ4Ύ���ʊ8#R��*#\O�b�8x�ܱ:�$1*����'D����/O� �u����^ɪ�@VO%D��p���Xk���N^"N����dl#D�P���@�`	�2��ƔD�T��e+"D���Cf�n �ȑ�Ʊ�X�f#;D�Dh��I$s����� %����A7D��"�	+*�P�FފpO��cB/D�T�C�M !��Ab�M���0�m.D���ޤ���h��0���(�,D��XDJR��r�p��-��e�Dd(D��t�ڃǺ��hײ�ś6�$D���4��Udq��a�"ޅb��6D�+�H.o����T=L\����o1D�x!��(Z�*��ԻbKP� D�/D�\B��<B�>)��H�	A�` �.D����_^�~Dcń@Oa��+D�L��dvXf ���Q{@"qʲo+D�@Ae��8�H�ċ�=���Cl+D���WCϗ�DTHa�G�3X�	�� *D�ı�莪54r��oQ�Z�� �=D�4s�HR4}��@� �H�P��'�;D��h�\�b��5�իV�2�y��%D���QL� �PِLҳW�Z�`I&D�rq�];v= �XZ�	#$D������b�v���F.�D��d�"D��饌��g5�:�Ç�1�b��!D�h � н�*Q�e)B(c}@ �`�$D�pB�	�b��<�#��W���7� D�(zDDNd�qdH��U��Q�Q(?D��Q� nD�]Adڵ<��Q���;D����Z:%]�0��k c����Ѫ8D�<��nQ�nDb&�[�Y�|=��9D����/ȋ)k��c��٭ 6���E9D�{���=�F��zl!P��5D� Ca��,h �0-D�3͚��a�3D�� f�yb��t{������,6�|��"O��2��8{S&�j&V5�D]8�"O~ؘӤW0L�R�:�.�#�Z���"O�б�Z�Ŵ�Suo\z�u�"O����iC�H	�Us�@���x�
r"O�I)�c��	]�y�3Z�nZ5�"O�-d�=ת�VlJIj�K�"O�t3u	��z̞��7M�QQ��@�"O�x�F�6C�B��t��YG��""O� J�:Z�N80����;>��J�"O�����S	�����`[���"O�DK�̙�E�B9��B�0P��d"O|��#*P;����3���Ga\��"O���'� 0�YU+�?���90"Oڠ3���!��E�] �&]c&"O�h��Oy��x�H��>����#"O�H�۰^�PU�CJ�V�,y�"O*��D� cB�]�3��[�bI"OH�CČT� cN�)`��v~P��f"O�"#D�B�y��X��sc"O��۱�7 ��A�3晦p�h��"Ol�@s��B�4�j<���8P#!��?:L�a���Þ��! !�D۶K��#%���V��J�V!�Y�(n�"��ݟx��xSp�ڷ^!�d�$�P*E��9H���ᶁ@	\!���{�@@T��$�(H�'���DR!�Y�+��U:6O��`�p�Ճ�#AJ!�$��2h=1��	/��ݠ�� �t@!�).��e�S�Iw���d+��`@!�$��;F�9Ɇ�$g��AE��9	-!�$��o!�B��f�b�f�Py�사fn�t�� �[GV��E�
�y¥+y �m@O@
��	��M]��y�	�&��U�b�\Mv�R�`K�y�.�,HR}p �A�A�,e�	�y�B��@{���D�:�6A�d ��y�"�:j��qB��.j;z�u�ۉ�y�OI�E[�Y��O
�$�*�y↏���rqIͫ7�^A�.��y���53��M���	2.#�1�7�G��y"��-n�L�Bf�8�8�� ��y�]9r�@�7O��8��	)�yҪ@'t �� L�o�m��	�y�!uO$\x��M{���h��P%�yr.04����D�s:�H&E���yR�xՊ�A��:�~<����y��5i:��w��0I$(t���yR�R4�&2U�Y.1�J�DdY��y�[Ri.��c ����R�ى�y�̹)�"M���ˎw�&<K#"�yr�� _?Puh��\�;	\)����y�C�7��u��(7�@]��G ��y��N3"u�P�A��rs-J�yr-�)Dly'�85���Sf���y���8B�� "�ӄ)���ՎM��yrg�h/�1��Y*���:d���y�o��Q+���S��$�8a0�� �y2AʊL(J`�WkF4P!�+�y��%~f~�ʣ�����è7�y�.Vr�&	b��Y�"�ȫ����yb�Ԅ��+Cؙ^D�a͏�y�H�"ȴ� ��:H�E�Զ�yҭZ����Z���,�3�/\��y
� P@��O՟E��Y�O�/Z-���B"O���gI�"q"ԑ����N��)F"O:Eh�CL�X�|}��oאs��<��"OnH�-U�p�	��8=�uH"O2�w�6v*B89��I'i��0Y"OR�b!� 1x����*a��"O~$ b��f�R���!�N�HQ�"Oz�rȞ6 �jeѴ͉nd 2"O>��r��Ai�`17ѐig��a�"OjePI�4^�N-3�	K��Ӷ"O�,Za	N�v_��Y�#Ե0J8�"O\��BEE�	E���#�- v��"O�5r���$�AzCIXV���"O�Qˢ��*t��\1�Gb
-s"O:��4肋�ޠ�5�Oc����"O$�IHôA��C"GG�y�.QhG"Oh��F�Ӌ P Q(����4��-�D"O�1�E��5Q��i!`� ��CG"O���V��HPd�����"O,)@��I6xTm�w��:)�Re�"O�Lӗ�O?v	x�&� �����"O|�����t���:6�,T`^=8�"OVxѭخ�JB#d8�QȔ�yB�"v�<��J�z����Ŕ��y��X�U#�i�QNxsF̢��'�yb�U.d�x�`KO;k>���,�ybfE5^xtd���Db�ꍚa��1�yb�D�6�����'\�Xp6�[Ҋ���yr�^�?SP��D��9���k"L��y®Ƭ<��q�!�+9V�=ڐ�U7�yB��*_� �b@���4��X0�ݹ�y�.�
fn����,�	:0oB/�y�@[
�}A&�߯(��IswKW��y���1>
��ŅN������y�'L7+S�[ƀ�'M���D%)�y�-�3�$dB��G�B 'Ǚ$�y���sV�kq�Xn(�m�v�0�y��0J��q���c�̸vdB7�y���1��|���Z��lKd(Z��yr���,�I
�k��	"8)3����ybe\�3�$��V�':Όc��H��yBJWt����؄Jl�U��%��ybd�+_P�A'ځZh�	R�yra=�Q�D�
�Nt�VoJ��y"��%1��@���*|�����y���O_n�Q6
A�6�h���*���yr#��Z��;S��YA"`yt�ϸ�yR�E(3خ�����T~��(���yr(�&E���c׬�7|#�Dh��y�e�e~!y� �4{k|���Ϋ�y/Ҡ�~��a�c�B��N��yb(HK�rQcǠ� lL����e��y�)Ȋdv�}ʡ��e�*h���y�Ij|�@@���X��tR.B�yB��	u�(@%!�P���[�k�yB�	�kF���a'@�LM\HY�kR��y�\<{mz؂�dwx���$X/�y��ݲXm�1�S�U�E]��g$�y��� o���R��	i�UYƕ�y"K&iY�y��-B�y����y���6,�b�xA@�uY���b��yRm�7��]���ԀC�F�*⎉2�yb�
���S���1,L-�A���y��n��z�/&R �A�Ĩ�y
� ؉hd��#��p�T�Rt� "Ox���4G��s���sL0��"O��p��l~@D��+�5�|)��"O1+CFβ��u��>��5��"OL���O!"���Dȇ�|��"O\���X.�L*`�˭��#r"O��%�N�hv�X5S������"O�*��\�x��Sa���"OH��I�|��@9D\<��� g"O�m��"��L\�#�`گA�::U"O=Pwf�"}��aQ,vj	��"O��r��k���A�NR�dA��'�D5���Z/�ͱS疗&�Z���'�B4��͏�x�6�ہ��7!�2�b�'��XQA��*!h ؁��!�I�'ԙ�CE��MA�e�(� ��'��$*�g�T��-б��#"]���'�6Y��ԇ�����S�Ef�`�'�JU�%� gDh9Cb5����'I���w�ZS����I�\�RYh�'h.iR𧄬n�h��
Q�V��8�'Δ:@�q��n�^8�t�\��yr��?L�&��2$q�m����y"o i�T5���J{2\� �P��yƃ�!"B�:�(R�F�H�Ä0�y®F<��@��G??��	B6,?�yr#D�c�Ș���$G� �
���y�]1��MqīY�&���ەN��y2��]C�(􂛪�N�YŪ�y��A�o���
3�,#:��:�Ƈ�ya����^8N!!��A��y"eD�}�=a֢݋!hi���%�yR%�Q�����U?J.��plF'�y�'L%p�U:��
m���k�o�,�y�B60��ڤ�R�]Y�I���9�y�J�H��BD�U=bQ����y��)Lƾ8�b���T��i��`Z��y"�,���`�Z,J��m2啗�y��,!:��*�o)�+$�Q�yrOS�9�*���9l�v������y�F��v��z��5��Hj��]��y�"Ņ����Ʉwb8��F�y�m�2o�h���K(es��ZC���y��G4�h��ŵ$��ҢX��yB\{d�����=S 0�"���y�N��8><�vCC6������y�,���Yj�Y8+F���]�y�H¼#뺼J��U���E�6�yҧʚO�0��/9Jj�`)ćƚ�y�T�8�bPˍC`�!�Ш�yb��3\�,m#�Il�H0&�y��]n,bY�3j�y{hQ�bF���yb��
yLQ�� \v����L��y��._�8�� ���i,mj���y2h�?V�À&�0nP&���Ⱥ�yBB?L��K*<�d���ۮ�y���w��uIdn�0(����ݿ�yb@
� ���@�"���`���y"� � �R�*��x�7i���y��@x&p��d^!���T�B��y�O��C@@�b��H�\t
�����y�
5^����KӬ�P=��LX��yrgC3g$�A7�����H�����y��(k��(` W�yo>��p����y
� �t��Q�wѬ0xBn�B(R�"O�|�E";r�HD-�x�pL"OT%A�嗲L�q�6-H�}�(�"Oz}ؔ�[�r� k�읫B��4��"O�yH%�C �
�R���$��=�'"OH)�f�3[���2��J�o(ȁ��"O0��#�Ú�:�	�#F�p@'"O��sBiހ3��|H`H�" ��"O~��a�3p��rsgW�8+���"O��ړE@�)��m�1�K~��r!"Oh�� B�B�� x��Jʹ��"O��q5N3����P%O`�8�"O�S�)ˁa(�A!4FZ>e��w"OZp�&�%p�g�ˢ#��bv"O8UᢤCo#�x���D+E�ـ"O*��+ҁ]�h�@�:%�B"O�0eǾAQ<�ԥňa�6��!"O\��A2;i.�yB�8\m�E��"O��!kT��x��A1m�`�;r"O�@H�n��n~	��Y��P�0�"O�]���ep��)�3���a"OH��,l�S��Ľl�HYA�"O4����HG�@���|`Bt"O�P��,�0<n����_���"O�R$��@�N4�H��g���Y�"Ohx���>@��&��'�"6"O�� ��A�o�2��#L� �ڥ�"On�1�Z�����ǂիa�\�8�"Oj��l�,��dr��H*R*<�k#"OX�:���4Q��` ��Cɚ�"O2�0���o�N�b�,אl]�x�"O>���KRx0-ӷ�^(NƔQU"O�I� �!z�d)��E�S.�eJ$"O���FO;��la��'-�l��"O��;�#� 9|�beɊ��)+�"O�q�B
"7�F)��hЪjբ1"Op�
�@��L��=��僦�q�W"O
��Fb��h�P�����t|���"O����]���j2C�r�x�J�"O��+��W=V|\�����'q���e"O����,��{�%�/F�*�"O���つSU��筊 �:�{�"O��"F��[<t1+�@�C�"O&E���(X�!8�.�L�h "Oe�����ɘ��@�ؽH�"OpуF�8���K�@K
]i&�*q"O�90ŤՈ'D6�
 N�B�`�*R"O�xA����2I`�Nަ3��8��"O��;CD��O������"Ohآ��+�a�͞�\�z%*�"OZ� i�3��Y�`�YK�@�sG"O�����a"x9�5戴^��\F"O�!;�͑�he�	�CC�+����"OĔ1A�{A&��h�0>�ژ2�"O����wI��x�?���y�"OB��0#�"`l���&xT0-*�"OƄj7aL2P�7�
PJ�S�"O@�)e���j<�uQ�ϹE�ʭQ$"OJbT��y;֙;C�	K�n��"O>Y"p#E�{�8�c_(}o�%��"O�P�Jϻ=����=5l\��e"O���♙C�L1S�P&<ʔRd"O��v�ZIc�`s$�3J��p�5"OL��`�V!qp"��&Y�f���¶"O� ����YV�{b�_�}�
]`�"O`� ���({=�Q��D�da�,A"O�����*��灂/tpv|�""O�{���!�`ѹ��A�0N���"Ox�B��V)f����V�W@����"O��@C�h�0Mp��/6��m7"OZ���إ?ޠp�e���C�ۑ"O�Py�+[�{��غ b�JWb��6"O��I� _�+����]�u?��
�"Ox�a`(�eTD9���_�y<��H�"ORD:6&�1&� 8�qo���a��"O��+��Z�qnNq���X���"�"O�}
u�O�.MԹ���H�fm
�:a"Ox�P�.OV��,W vk��k�"O����DŢӌ#%S(x0�"OVb�C׽eT�8�tj$���"O�ؘa��<5�b�3`瀈"����"O䄫TFȠ!�d�3�F�9��1p�"O6
��,�s`eQ$�J-8"O�9��ƌ|�V��Yn$Щ�"OtC/ɉ?��y��$B(]�00a"O���@��GԤR�c��s��X�"O���r�u��AEb(o��2"O�a�4,Mr��b!T;XQ�Ԃ`"O�=��CW:{��D��%�	�(铃"Ox��Bk�M1���C�S�.'ּ� "O�QbsG1T�``*X�lx	Є"O踛3A�5̼�����Ipl�;�"OPy:R��L����NC�����"OYɑ��>�ԓp��2N"I�P"O2|�@��>9:j`�W,[M��"O��3b�9a��Ip���_1"�`�"O��X��<%(b�8�%��W�%K�"OP��u"�*DE��ZU��{]�q�*O�DhBO��iʢ.Q$$��Hx�'����([rXC7h1�f��'�pȅ�32���ϊ�(�ͨ�'��A���*�B� 	mf��	�'�X���uea�� (t��Qq�'d�A�'C�t�P7�`�,I��'	���'�Py�;��Dh�2ܛ�'���ra�R�NQa���e�X�
�'L����`�!kM|,��hR�**�<	�'R�Ɋ$Q
(��5@�'� a��'�������o1 �CA^�ڍ��'8�%Y�=@��C4Θw��3	�'�\uÃ��!	�X��@f�E�HH8�'���%�5��1ۖ�E�tJ9��'P���բ$��rmI/ev���
�'����"Ʉ ZI)�ߊa�����'Q�Yb��3&��ѧ_�#�(��'���yS-T�	:�@��E����'�<�Ǜ�!%2q���	;� d��'��S�[T��Y�Dڜ-L��'A���U��!<<pFW�&�jP�'��eӣ�ӝ8���d�a48
�'��al� :��x�AK�X�b	�'�Jh#�C_z� �P���K���:	�'�!0��|jZLS䅖��ҍ��'k��®�:>�*x��>�:	�'w@풵��q!Č� �۟}�Z�'nQj&�Ot�T;��������
�',H���FNT���fB+����'�����R�y�H�W�ꘉ���� x�fe������KM"�@T"O ��Q��vm*�;P�!cR"O��hT��cE�ٺ���*B�����"Oֹئ��M�c�L[��m	�"O,iAd�J�j�b��9��6"O@d�eX�h�B2'%�z}"O~����Zg\�����IB�p9��"O�,1'��.q�uB��ƴ���"O.�y���2Ўq�p�F��ڥȄ"Oޤ��C�Fn1��͞��a�4"O��ʴ�<8�4�C	�%Ju�8*�"O��IU�՗Xݒ�&��mo\ɛd"O*H#�NX)�@qjp/��:N��R"O�-!2J�:a,�U�c�R0/~���"OȤ҅)
#!�ԥy�UC��s�"OV%`ҦO^z��3�M!c���6"O�i�j'4�,�s�A�o&��s�"O!b� 
uҡ��%?X�!d"OB
 f�0b�v@�m��K�: R�"O
��#��S�X܃�R 	��a��"O" J��P��ZXVlX���ҷ"O���0*��'a��'�L�[h`��"O@���$S�A�N
(�|�qw"O�`A��X�|�e�з9�^��"OV�@aK�/�0���BO�8�
�"O~%�6D�oT;�`�.=��|f"O��Qc	��H$�:�o�n�*}�V"O�eiqΆsy��C� H;z���"O<��mA'WUPh��̬z<��"OĤ�E����V�� �b��}�f"O\͢�Ȟ�Z�P�R�o�m�R�2�"OJ�FD \v={�-�<��(��"O���`�6Y@N��+�_�jђ�"O����]��ִ"�����]�"Ode��%�+D�F��#[��p�"Ot�ஆs���3M�+S�Bqҥ"OM2��^$�Y	���(�Ԫa"O�e:4�U�Ev���� � �G"O�� ��oS���`��3�b��"O��ءd�5�F��J�:bǰ�$"O�!U	ɭ9Z0���i�.T���t"Ol(b%�#[~��iC�d!1b"O$Ly� 
����+1Ji�⑑e"O��B�^��}�$Ib��.N+8 !�$l��	7C��,s�x��jĦ<!��*s�1�aX\.�ц �o�!�D�9LMXx1d��	{�oUB!�D��ke��iT�X) ���A�Y�!�V4D���n;)�	b�Z=�!��;3��Ԃ�e��o�t�@�M�9�!��5I�t0Gœ)���P`�a�!�$��%2�)Ճ(U��,0����(n!�$�9��[����a�����DJ& O!�ě36p�<�gJ���{��R�Z:!�DS5GcV���͂�o���V�!�M1.2Й��@�(�\�Q�[�S�!��C:aCfkR���е�ɡu�!�$�o�vD��G���QQVi� W�!򄑡/V��(C`��l�py���5|�!�D19�y"$c!H�rA I��e�!��ƚy����Zz~*��GƥC�!򤃩r�D#�#�TULl�u��YZ!�$)�T�R�lT���q�C�&�!�d�I���#W�W>D���Q(3}<!�� $\*�Ŕ1H!���B���-!t"O���U�1f5�b���S6�0W"Ol�ۑO_�&��I�d՝�B���"O �֗=hY8Ʃ�&'���
�"O�HZ�$�"4�8%�X�Z�2;U"O^Ų��#�*D�&ĩI�  I�"O�l�B�7��#Ƃ�(��p�W"O,$�3��D��<)�֨(~v)("Ol�
�M3:d��8 ǆpݒt�S"O����ܗ'�@ك"'�(Ŕ��'"OXܱ��^y���X�fA�R�bv"O��a�2h�"	�%�JO�y;V"O��:EF���X)��=��ɤ"O�=���ӭ{L�,#��C(�P"O`=zV/חi���cʌiM"!��"O�P�����D��$@r�ɹa;.�3�"O�M�����x�"˦G��)�"OT�b^�Pc6	H�`�@|&=X�"O�p��Q�H"��悈Zx�IC�"O: c#蝾�:��$�*BY���"Oȉ�'�=��a c֫<D���#"Ol��Dh�%j����'���h*"O���Bhı,Ԡ���+Z�O��"O̡3�S�.
 � �N�YX�E"O�`��$q����.t��g"OJ!J��2���۷nş^p�:�"O�d�e)��w��$(�bׇ\��MXC"O�<���I=*�P1��������"OF�����7� �� �E��>�""O��v��ohH��&O5��QQ�"O��`a\�	LΩ +En���Rw"O��je�ޑiߚ	��)��u�^��Q"O|�ˢ�D,*�z� �!2 Pi�"O�$���/{p-P��Q�U�M��"O�TqTiիS=��A�f��?�Yx0"O������')fn��ł����9�"O�lw+L�i�t�#��BBαr"O�Bf)��#�b�X��X�|ǎ9W"Ox���8`��4�G*�~w�� "OZ�P�T�(�j����ss���"O� b�'���B�ÇF֫��q��"O�k�-�"<ؕ���+���w"O$��l�Y̰�e��S�Pu�"O��Q�^�Р��R%<����C"O�|��' �IR��)�D?1��1�"OT�Ð���E$AP $�%,h�L��"Or]�5!��W�`	 �	� .�"O����ߧ\��	BK�R���)u"O`+��ɬ�l#�iб~�t��u"O�=#�*Fq|hg�	��`�4"O�=E�QB:^ �ˌ�3,LJ�"O��p�hG�l�ƥC!��]"�	B�"O`�R:em�Ĉs	ݐS~B�J�"O�I��܏c�$�pFϵxT�d"O�p0�E$
n`�$-V�q"O�p:�I���Vm�A��ԨO!�$�*ˆ<*2F����`�T�&�!�DQ�|FH�+҃״P�a{��Ɍ8�!򄒝'z�x��O&�J���#��!�$�>?*���	j�e����7N�!�DA�Y(y�t#@ Ab�T�d�k�!�H�6rj��U��CR��#F)�!�d�a���zր��#K����	<�!��[�]�4
W�. ]V]�Gȓ�P�!�� @���l<?�P�D� ��T"Oh�x4'�1Dnv��e*,s���˔"O
�����<}�H�{��=���JR"Of�!���?)������P�#���h"O �n*�����_�1g�[�"O�Bf�D>eRx�C�.[Z�p�"O"���� Mr��k��E� q֤�g"O�m"桏�r�q)&�:&mj��"OzT:�!��|T]��׾ kȨ0�"O����E	+gpعQq��N���"O&�K���P޴M���\K��"OZ1���H�	�E���6Q�ĭ	"O��H �^�[�dY`������"O^�����!^2j��N��I��(�"O�c����w���ѱ��s�L�9�*Ot�AVj�Ju�q��#�%4A��'��� �e>��
�
���'�lZE�N�S�nXx��D}�����'�*�7�ʭ�t��2+0e(��
�'��yJ�ʀ����yRL�+_����'(�ese�o�Ru8�7kS��'����&0E���P�Z�y�t�
�'xq�!�=0��߸~~n�
�'��a)2h;�z\�Aզ}w�e�	�'�
(2v ��q��)r���cP"���'Ė8 ���&bl�"A�օR����'��+eF�*A��%��Z�}o¥ �'G�5JB*Z��W�_\DP��']�m@���>�Фط	6H]�
�'�81������@w�	�����
�'$�yc�\�hǞ�y�Ƶ��A[
�'�l�ʁ ��6R0�uB�!-Nm��'�,�r@"	��V�D�	AP�p�''D�:F��
hq���c(��(���'��uʅ*�f����eI��,8�	�'R�)��À茔Ȅ!�<�Bm��'�i�m<08�Aa��13P����'���P��_�T4�b��ǿ�ʙS
�'� :N4o|@�صÕ����
�'� 5�@�G���5n�! $�b�'�F�[թ$?��p����z/�}B�'q,�H �7VD`�������'��; �N1ZSl�!Lx��c�'Pt�ׄ[�+����"��v�9j�'���q��ʐg�QEO�=��@�'��a C�;8�>8��(>��� �'K�Q�]�H4"dK$5c*<�h
�'98�����KĠ!ITI����'���9P�A�h��ͩ��3	�� �'�$HC� �))F�cAŁ ���q�'�`����_I�M8��xALU)�'� ����d����mH�t(��'}���,E�(�ZF)�,v�P���'��P[��ǣP �H���o0~��'Ӣ!��eǑ	^Hc!�fC|(��'����dܭ) xt�ϥ^�"@��'ɔi��D��HI��h���A��0�'X�4[�۠u�(a���6kv~M#�'^��kƤ>�J��e�>���'���;�@�
s�6`"N��`�]�
�'���� ��9 h��՚0�Bȡ�'�f��ABA,0�:Ȣ�k�U�`P�'��Uz%	��v>x�ʠ#�G�H|P�'�8kRI�oP!��ђq%�(��� ���J-flB
�"�S�z�÷"Or= �h�R��SB�Wm�1�C"O���#��A~5����4XY���"O*T�rV)K�(8��`� �yV"Od�ْD�;2�HF<S{(M�"O�D�V�@>�q3��%nN��7"O �鱫\�$��r�$�({]�Xr�"Ol�(4��7����0) �j6НR"O��G�A:�>����O�	�����"Ovx��ܖ4�(��|�ZY"�"O�⡯�
��ɒuI/��i��"O�1:af��M2����nB�"4���"O�Y��B
7=4��m�RPt<�w"O��Xs�Z%d羈1b�\�=A�Cd"OL5�d��"|����E/��"O
D��bǨ|�
G*_����$"O��3���iB�@�1)EK��U�b"O��a�ᙟ%\���Hƌ2�V][�"O
�` Ƙ~2 {�hV��p)Ct"O��ff~��1"�8�T�a�"OZ`!�^T�4�"�Q�;��ę�"O����&�|�4H��I�z�vT	A"O�l󓮄6s���rE+i�}�"O�@:��yz@���C�`�>��&"O*���/(pn<��V�M�>)�"Ov����ǅ�4�c�*A�^�RPK�"O�a�E�%0f��I:��k"O4�8g�Ш\�6DPшLmAs"O�$� ��U��}�JIZ�erR"Ou���	07�B1@�H�E6�k"O�iC�N�T��#g	4
d
3"O��
p�;AmB�B���c��I�!"O�3s�^U� k�Mӻ`�,��R"Or8($!�1)���b%M+U��}��"O Uqs`��T�"g��=�0T#�"O�s���Cv�5¶#s�j (�"O̰I���8���٢+�*\Q"O�%Z�F�E4�i%P,g?��C"O��+Ѭ�!8/ܜ��B(?*��W"O���a)�pi0�(��t"`"O �6�Т�1�d�H)-XP"Of��T�I�T^�4
�kəy�dQ"�"O�P��@$}���a���V��B"Or�W�yڌih��˴K�.��"O|�'���;h2�'D�T�I�"Ot�F�#Y����U&\!4^��2�"O,< vkA�w�r%+R����̡"O,�3�V�p	�E��_(&�I�"O\��gG.LZ�"%bG#"*��aG"Otije�"�i"�%*&�Za"O� 4� �Q?n�9�a/N	L�
*On 3���c
�b`/�3s� ��'U蹫�ީO��a��@!r���@�'ƤPBG���� BWB�As�'�rDr�*�-��U���(`z ��'�����S��i���*~�z�'�l��q����=��k��֐Xc�'іX�-CֆaÕH]-F͉�'���x�$*�F�u$ŕ[�����'=4�rq��:_� ���&�CĢ�:�'������\�Nu2H$Μ�	�1��'k�\�#��SK��0"��O�F���'U�����6���+"$�7`� ��'#�����G"���p,����	��� D��Ǝȝ[�����ϲmx�""O��` ׆)���`ױBn�#"Oz�bnN>�\�!���
Lb�r�"O� �3cW� H�H��(J�"O8@Y5)��9�I�4�ȏq��Z$"O` �!��+f �8!�# i��3"O�T�"��/�Hp�^c��ʤ"O*�R,���X��@�|�>l"O`x�� �1#��B�I�A1�4�'"O�=R4@�{)�l�D�̰NF�"O�jUgB� &��")�+-�%��"O���m �9"5�+ �4<|��"O 5�B.[J�đ�	��I��!4"O(XFű\)���U��+8V1�"O8�%�0��$����'���"O��P��B�+�|�f@[�z �h"O��dD����R����2Ux�"O�@cB��(���G\H�٢"Ol���(�&x�E!2J�	+]����"O�I��(& �&�ԃ*\�\#&"O$@�"�i����'䆗JZ��j"O�Т��($��B5]&0�S6"O,u*�P�}O|!d��1m�re"O�A�!F��~��)���4P4"O �i��T�&�,s�@%mB=�a"OTXӓG�C�*�nՁ%H��k�!�$�8C8~��`�մ�NLBvI�T	!�K	�
%Be��K^.�;��I	_!�D�>՚M"�@GpV4z�E\�!��3���v��6J�!2ÆY�*{!�$�=z�(]��ja��Xru��>\!�d��&z:��bU%���w��2K!�Ě�H|I�$Hq�����!�-p�!�^�`��A�e�;m��%�r�R�!�$К�IZG*�Z�L�A�|Z!�d�O7���O2Q�&������%A!���Nɖ9Z4�ɕE���"2*�1!�Y�k]��#a��n�����9�!�D��.¬�D�T+jD)����-�!��E��D��ɁoU�q��Z�!�D�3=�:k�58���\�u�3"OTy�a�ؚ�8�#%���'�dm��"O�%!�I�`m�H�e"��p踌z�"O�drB%�;4ԡF(��}l�(@"Oإ@_�6Т�M�^S��`"O�I�`� j`P�g_�&O:0Zs"O 4��&u�4��Gl
92���"Ol�"���>�h���'~Q�"O^��"셪t:��'Γ1&��+�"O2�g_����@%�"U�%�"O��1t"��x�7%TVd��w"Oȼ�O�;F��(b�S[ܰ�G"OHLAfc��x8�1�
�SQqI�"OD����	)xt6M�#�ν;J��9�"O�|��˩>cؤ6�ƹ`��{�"O���եQ�
0~�:4� 4pIP"O| :A"F%����˫y�$�"O0�B�-E�1����Ɔ�5$�*�"O*�+2 ]�r=�"%N�%� X��"O���Ƅ�M�Z�鵤��>�TTq"Oh�{�LEb��X���>��a�"O�|���ca����5I�ѹa��/�!��X)N�29���7e:�`k`�Ԣg{!�dV$d*��h�$|H��n F!��  �r&�_�a
�����]! |(��"O:����،B�$-9� �3�		�"O���"ĽK`�Hӡ�C�u��e�g"OP��ĄA�C^�m��/ߡ�)� "O�傅T5f��l�D��+%���"O� 0���[�,]��� <ih��"O&I�A7#4i��%a`x��"O��)#֟��4d�j��"O�43��L4����Ě�SUА;�"O�Y�)�%"�����C�:GY>�p�"O��P��\PX4���/&XPX�"O�XJ���"��
$F�t���"O6!03�R7UY�x0��Y�H�r��b"O�-�	R@T��/�8>��Pp"O���e��k�`c�͋�(��r"O�E���Bv�91�L�H���"OT9�Ӭ6��ex&��y�$xp1"O�t�7�6��X6dC7+�a��"O�8RBT�+$����H��rǤ��"O� ��,�*��5����Y��p��"O����Ƌ�'�b��Ƅݳ~Z�@;4"Od�S �ֽ!�R�ѱ"Aa2�"Ol��t.֢1G��
C�.���"O��XA(�tO�+&՛R�m3`"O�LS�)�?D�y7�S"���"O����ݘ \@��a�FЋC2�y��K�ow�E+�}��1f���y�)څ@�\M�'&$N|�%H���yr��,WH��ȴ�E�*�IԱ�y�oW:�b(C�G"y ��)� �y����X���.V�|� ��ۼ�yB �2\ъ���C.m�h�����y���#�B���5h(j
�B��yr��c�����,Y,΅�'���yҧL6lQP{��_���7���y�
:$�� 蟡U�x�'$��y��X�XPⰤ�B� ��bW��yRǙ��>E1���75{�*��U��y��	(L� ��Â5$�2��DF�y�%�7e� �3SiX�)��РN۱�yB@�RU0�Ȇ�M=&��u��h^:�y�i�!�H@��"�:�eA��yRÇ�@TLi�jԾ$��	e@�#�y¢���1p���[�����yB�T�$H�)�=*�b�X��	��y�.O�aT 42�ˀOTu�b�݆�y� V(v����78�ک�`+��y2a�lN�QsĚ�/P~j5���yb�Ӆ���,9g��3*K�yR�&>o(-���F�t�`t=�y�A� :~�1!��Cl`ţ�JW��yR ś~l���rH�9�4�e��y�g�'N��[B�amD��G�&#!��v�X ���S���p�-}�!��)	�Փ1$�rn���T-CN!�$�=�y�	ڰ
q�|@�O =!�D�&F<0����l��P��ԋ&�!�䝙J}XA���Q`
!Aw%�!�D
�E��$�5�Ζ)Kj%� ��a�!�S@�8 �6*�l���ԯ@�X�!����Eг']��P�_|!�$	�a���l��>�5��B�+�!�D�\�܉��ǉ��|�g�u!�$*2|8��䉞R`��POwm!�� 
����M	�|��u��
4"O2MZà�3[�	۲B�:ԠP"O�	*%8h�Z�8ҠU�B�� �S"Ofib���N�yKՁg�b�2'"O��S����l���4��1�"O
i��N'W^AS%n��b��"O���!�3�
Z�LE�n��	kq"Ovd��	��������3�"OVU���H*l.d�S�- -�n���"O.]j!M��6�	��+E?\����"O���ō��	4V��H]&V���j'"O������D\J��)
�<�n�[�"O�8���(D���C�j���X�"O��r�E� Y˪h��FN+Y*��"Oح.�<Wt	�6h��,�T�w"O��K�K�5�rSWf�R�|�C�"O�Dc
)�L�LE�Y�� �"O�y���I1���f��L�
x�C"Otxhr�^�,�dh�ˍ41����"O0 ˷�#T�R���Vh�0*t"O�����'֘:�+��B�p�"O��aF�8X��<։��!��8�"OD�WlJ+S�V!�R'ͦE��,�"O���
7�f9B�P�\���!"O6��amIB]ΘkgfȔ8�ɉ$"Ol�"#�Y�aT����L�z	� �"O��ꔆP3J���c�J���h05"OJ�C�օj�;�	8ކ�Q"O>�ItӅr`X'		�Dq �"O� �� IF�-�E�#�`�x�"O^1���%8��e$��@�@"O��P�L�Ts����!+�:��"O�M�b��0w�陖I��ݸ7"O���3��,��E 4H�7*��MB"O"�ST�Ԑe���ȝ6�Q��"O�+�Ä��8�D��#43Z���"O�*c������C*?\�#"Oz$Q���.D�T��إ-~���"O�@�C�)=�d��,QOw�k�"O.xh�>2ؖ���Ȕ,����"OtQ2T���9� �a�Ǐ�AF6u"OD��gGк���@��y?��S�"O�\KàdlP6n��~��"O����Ǖ��Ny��L�Uƛ��=D��!B�K:RܞLʦ�ך]da� A=D��J�J!}�p���'H!�@�<D����H�5�t��i�9c��Y�:D��H��`����K��4m��Z#�7D�L�� �c���y�	G
H���i��3D���A�-b�T�G��#2"�1��1D�T� ɂ��0�@O�(�D�.D�,jG� :�A��E�O���(D� àl��H�F(�F�0��W�&D�����>c��8���4��Ct�$D�8i�*��>]>���k������-D���F�I*I�PŚ5���R���ΞT�<	�`�A`P�������r��L�<��,���Q�У�)P�MA�+�c�<!���>9�L�tC<"��=Iq��[�<���U������V%'��#�fCl�<��ˊ:xs}�HTA��lSV��k�<I"(˿|
�rQ��[�䩚$eg�<����?+�YQ�l��(��5J�`�<I��Z��sHܒ.�L�Dm�X�<� ��j$������ )�<��iBQ"O�d��"���qpC��[x��"O��bҤ�=]�ܡ:tƕ0nP"O�cŉ/5�p�a5�Q�J�Q��"O�I��!�,$$�R��þ3�U�G"O110�:"��	�f$B�{��@�"Or�c�l\��f�P�8�x�b"O��2�7�p����L*j�ʑ3�"Oܡ���L�&S�ۨ|�F��"O^1QBԬl��y:���(�"��u"OT����WPrD��>�N�9�"O�Ms1��n�9h�I�.k�&D�"O���ʎ�V����H=Y>�
"OtԀ��E�F㈬Hᡜ�@����"O�Y�'7X�AC�g�,?4l�£"Oz��ה
���ã\4d)���"O(@q����FC�	U&f��"O���DM��I0V$y�	#Ld�'"O�D�5H*T��Asm��p"O��' ,Z�p�:���9FW�i3"O(��� ܀�7@8đ�"O�8�� 	�$�Ҵ�%�%��٠"O�-�e���u�Piԍڈ_h���"O��[�`�	f�*4�G�ܡQA��(�"O��I�.~ڄ1�E��q%<�	�"Oib��đ'[�	1�3R`a!"O�AC&F�`�T떃U+��]�6"O��F��(
 �;!�F�[V�5"O�YHaF��^ ������P(�uX2"O����l�j�2��y�\���"O�e���pB�x�T B�ܘ�"O�\��-��@��I��R�{~<|�"O�̐�f��*�ұ$L�\a]q�"O�E�dnה����"S�H�(�6"O���A��*c����AA�H��"OF	�@ۥQ���1��$.@�v"O ��.H#AE����@�:(����"Obp��K�w�<���k�q "Ol�����#���[>�J�"O�,���jmn�0���E��e��"O��r���6&���X
��Ii�"O��!"e�/+����hʂ%��p!E"OԹ�(�F�v]1��2O�H��"O�ц-ˌ;L���>72�=�c"Ofu�@�7c�Zy��عx;�i��"O����ٕ��Ӗ-��I(��"O�D� ���0�:9h �H9API��"O�TKFg��RB�W|��Y�"O�hs�5j���шI�
�j�"O�=)�I�6I����� �=_Ҟ��b"O�$�d���:�y0��4gj$ɒ"Oj<��Ȅ"VL��"��E��@t"Ov�q�fY�u���p2�ƶ0���c"O	��dK��4u��1�jX��"O. �H
H�X��RL
���"O��n@�8M��k��M ���6"O����O�H]�r��ܜ�y"O��C�H(;�6��@L
���z�"O��V�� X(���O4*�Dp�W"O!��Vꖸ`n>A���"OT=�Ԉ�Y>��GO��ΐ33"Of����S�C;T�`�A))2�-R�"O 	�Uo�U|�@�L� ��+#"Oh�����A_���c.P:�@�t"O� ��S�a@6MX~����C16�T!iD"O�-��Š@�R%ۥ��<��x��"OBehr� >H�P[� �%��;�"O*�+uK�#1�mY��P�;� �Pr"O�y����se���@�2�����"Oȭ�J�7@FMrR���k��� �"Oz�0��2j|�@���vdFQі"O,�j��рI��P���E��!�$��C9�J�$��6�li���jZ!�D΃u��p$/S�9��A�D��Vq!��� Y8 7��%h��F�>�!�*"�Ȋ�Ǘ;�y#��Q�&�!�d��"��ǈ�`��a���dO!�$U},T8#�NܪqRM(�MLQ9!�Ćr��q�dL��Q�b���̇C%!�$R� �a�Ǎ*^ܑ�AE%	!��D V}& jwJO)[�A����m�!򤙎^CFp)�$	�,� S*�98\!��]�P�pM�P�4�(���1\!��W7jj]��eD"���'�%�!�$ʐt7�9��1{�%`Ǩ���!�D�!JEh�Yv"W�zr�BH(*�!�D�=8���B����Q��.Z���ȓ��pCU,�>B�h���;Z\v]�ȓ�F�b2`R�Ho��H7bK�x�P��26��P��1ky:x�ѭ�
#�
�ȓ�*\�$��'\@q���5���5�,���a�%/����_��L�ȓ>������˽>�!8C��+;��@������%OF�M��"���R�ȓB�(�A��N+_:���(T�D��/��%���=OQ��:dO��^=�ȓˌYPko�NA�)�%�ȓ0�~9!�n�>2>P�0u��b�h5��AD )�hǼK�6a�@�˒gK�)��p��9�U.H�ҡ��'�7�
!�ȓ���SEA(JShIң W�c��X��m)XٛK�_r:\��-PaĆ�RH�J1��F���B�jlHE�ȓb1ts6�	�K���a�H� G9*	�ȓ9�p�`X����5U� M�@�ȓ*X��gĸ]V �茿)2�M���Ĝp�����L�R�^܄�n����\6�����ц9: ��8��mQ�D��M��I! *����ȓG�t1��KA�`� ���ټU2��T܈1��A�&z�\� �G�5NH���8l�@ؑ�W�����
�G}�X��Z3�L��솛,�rts5'Y�U�^���a�©9�-ɂU�X���
� wJR��S3(T���t>�1µ"@@ ��g>\���Ѥ�*őD#��Z݄ȓlT����,�@!�-�>1�d��T�AS@ hW�i�D�dD��ȓo�X��G��s��^��)�ȓi 9r� �$I�� O�V��ȓC���P�e��f?��H��;��=�ȓ9U�D�X��`��чQ� U��dD�y�DL��.�^x�t��F�zP��~���HMV1I�YjvnS�0���
���I�'/�X�1�ԧk�Q��M�mBRb�M6Qqv�[�?M�̇ȓO(Fp��i
�5�^��"l��a�p��ȓB�����K1N���Cl7.�0u��S�? ��'����)ˡ�L�W�|+"O����*V�w d���"O+e���
�"O$�%EA�J=[EdۏU��QI�"O��I��73*�`�O�͂�A�"Oܨ���XO��b��R	^#��X�"O�:0d��!��Q� Ra���R"O\=y��H�Z���B�>&��Y��'M�	̦�+�BJ�o;�h��7��9�%�"D���0��5�vP��%�{V��f� D��cʥ>���X ��voD�S�<D� ���PGTܔ���GB���@0D� )G�Z!i4���a��M��ABrh1D�T��A�U�sgјV�z�sR�3D���u9+�$:Binz�0D��hǶl'NhSRe�9W�2y�B�-D���`�׌AbR��1�
VΉ�n.D����!<w�MX�9J����j-D��+��%��!c)ԠAިȉ)D��" ��I��d ćVφ4��,D�4�gO̞Pd����ҶNx�h:�/*D��@�G�8���M��(�Y*rh'D�<5o�/�T|�4`����Q��%D� {5��_
̐dT'_���;�-/D�P�E��b�̴���ͅ�v��7�.D����늾vc���b��%BY,l�vlӀO��S�3���+�8��C��)2�ܨ�@�Luџ`�=٨����1��)M�wb�$��A"OJ��rGC�N���v��r�^���"O�0aˑ.U���b��D�|�t�"O��u�,DB:��}[j\YA"OFUB@VG����G��Rn���"O�`G�x�H0kt��%Wv��h&"OL�3O֤x@(�RkI'��Pc2"OƩ�Pq.C �֡4Ӛ�Hu�d"\O�5�pB�%!����ᄶh�d"O��{5V�84�'���L��"O��j0b�Gj�,8���+X����"��3LOJ�;3A�D�~P���0"�����"O6��%�;#jǂ�Y�6	R�\�D{��)�A�qA����L�+�
#�!�Ė,W����/ٝ�f$�Х���!���($��H�pIɼ0�/�&s!�dB�s޺����B�D��s�.2p!�D7������3(�4y���(�ay��I"��9�c�V1�d}	0G�;a"(C�I�����3��+3w���C��\C��o���9�蛳PR�p�f�B�@B�	�~0賆M̯^�t�A ,��*i0B�	�$�����Z|�pn�=B�ɣz،��d��0(h��y�e�4/u�C�B��5o�:-R�������	q?�{"�	�/�M�u`��v�
��?,K�B�I	�f�뇥փ(FL���77n�6�3�9?%?�O��wIN�w�@��pZ�Ī�"O��(���(� �>:��1"Or��hV)-� 4�v�A�SPlqK�"O^�2��?��m��G�.J8�!��"O��3c$��(�+g���d4f�[W"O��k#��%U�P)�?/��`"O�m(R��m�`����V�	��"O.ň����f�t�t�Hmd�EB"O�=d��O>Y
�(I>7_�ixe"O��eH�x �hX�aE[��L�"O
4pg��=u��_�R����2"O� R1�ȭ)arŐS��hm���r"O� K҇� �lk�T�.X>��"ObHa�.�bC��9Q�%lhF��"O�٥��rj��!�Ъ/U�p�"O�ɀk�T.qz"��@M��"O԰�� H��M�C��$Z2�9Ȁ"O&� k�;����T�Լm%����"O�	 ���""Ĝ4r�&�G���:�"O���k��@׸���Ȅ%��rT"OȀ5C�2X��J�'��Lj��Q@"O� U�٢�"c���Y5�I "O8�Z5ʈ1;�t C�Y�o�w�yr�·5�L��aĸa�V�R��=�yr��'{��D��ZTܻ��_��y�mլ="y#�H��(�<�yE�T̔�c�HO�@�x�y%� �yB��Gt$QaDǫ>Bz��� �y�J�)�,0��;=s���T"���yB�P ;hH҄�׷%��S��y%/
:���dI����LE��y" �>�|���Q:F��	��� �y�f�8'?��X�F:0��%i�`,�y�W5V�u��ŕ�&�^���B�y2��nSD,����)��A`񆍪�yb3'Vi:���Ԡ��$×�y���{2@T{q@��q,����,�y�i�q8Rdh0`0��0Y �]5�yb*�
� �1ы��[4�S�W��y2���X[�	7��"&��r��y2*�=G\L=91E�j|��Z:�y����Pe~,JA����5�$W��y��{T���؊^��b�E��yr"�<\`	��ꂓX��0�DD���yr��Y Q��$��d.�#�D �y�GE�4��H*�iK�Y�>0�E���yr*F�VW��r�c1N���(Ā޳�y�ID�*���I��JҮ�裋V��y����[�.PsK���s煄�y��ދ[ 2�s+��o�&̓�jR��y�l��� �p�9�t�k7�]P!��]�N�Pd��� �Ԗ<b m)!��ɉ2ЪuZ�蚎�t[)J?+1!��M�,�<p���ͱ�X��S�ʽ&!��[�7����e� ����$!�ǥ8bj P�\>3|�X�5A�Q!��ɹPU�*ԫC
J
��ː D�o!�Ĝ���y T�L�k�VD�7��l�!�� 0\>��4"�A��f,J�+�!�D��l:���oGz�F��@a\�I�!�$	�B�ʌz��v��+�)P�l!�Ȓ<��(���t��Hz0nY�'�!򤊋:�N��(�+w0AQ�㐺�!�$H�V���'�i�ǃؚSE!���LVh�&��&���6bB�4!�ת����!�O�������<!�$��d��Ȃ�E��qw��X�A�z!�Ā8gؒ��C���$f)��C�$X!��$p�b��LAa��ڳ)PG!��%#����e�f���b��*\\!���@�@a[V��L����Qf�\.!��`R�L���G�P�BiBA��<Q!�DC�[a��@�l�,���!��!�D���#"��D�W�Ի"j!��(9�Ĝ`��߸�2ݢヅ3@h!�� ����hH:i�:��a����#�"O")�jJ/o`̉%ծU�@���"ON���>�ؙ "K�%y2݁�"O�� "��`��@��*̹7%�!�"O�$��:�R�@����ĲD"O�4�̓�.�b֌�9)��}�6"O�Tɢ:p�p3nTv���'�(��-P�s�60�f��&zl�'��le�:�8�ö�I�zː�*�'oH���A�7�����|���	�'�fM�T�G/ T�ptN׽K�0ݱ�'�t�� f�P�4��NM)NG���'i�\Q����jy�k'BS�v���'�� K���\հp
��D��D��'�(87e�]�F�ˤ��AJ$�c�<� DA�)�����Q$r��	�w�<�Qd�6R�D�$]!E�pP��Fr�<��R�},�:u��"���
c��l�<�P`�2�\*b�OPک2�g�S�<q�&-b���K��4��l�B/TO�<)����K/���%�4S|D�	��t�<�l��kq`)��, r�)��s�<�!��$S�
e:1�Ů<���%�Fj�<���]�"��x��,%	;ll��+�`�<Y�I�>�bN�$]^�*0�t�<�P�$�69
��7 ��q�m�<��B�.���"� �%�@q�E��O�<�hʭm��`�-jK�P�EK�L�<	!���&�Z���]_ 5!!��K�<� 0)���
���"<��ib�<W�09f-U#H"��re�<A@��>�T}ق�y��d�^�C�ɀ_�Hl�W��)X녯�N�C�	�u��%��� /�
݃�])Z�C��)u�q��;R ��*]���C�I�UKN���왼Pv5��_�NC䉠	i�%S2��+z��r��1VtC�Eh�	�c�o�։@���.� B�:����[�E���i7��b3�C��6d���[T�9�E��	�4P;��Y9B*����/�Qp�ӹ�*��'_�!�$�MP��D�Y�Ywh�j%%�7�!�����R�H3M�4���؇~|!�($[RYڅ�ƖU�4�aW�J�Y!�$�}+�8�p��>�x���۞\)!�D�9:�@�K�3iVp�,´!�I�n"}3�Ǝ�MGL'�ߘ�!�Y�e_l��/F�b3BE���!wS!�F�rD��J��]X���C?S!�DO4҄ ��T�Z5�8�viQ,s6!��x�])*ó!L�zd�ٍ!(!�Ȓ.a&g�C;��5� �H�?.!�$Hz^8S��I:-DX�*ΫO!�Z,8�,��`Ђ�p�P�K"ij!�T10!�7�G �����Ik�!�d�A
Qk��U�\��+��B+%�!�)Ѱ��5(�e��uB�f� q!���7w���Q닅a�^�x�E�\Q!�dQ�YS��T$�'L��Ms�U�"T!�7
�"� ��������'!�d�
VF�c��A�-kp�ꆦ��r!��d�� �G6S�qs$"y"!򄀳t(@Cs��'bO6�:�C &!�DQ.X�<SW�-d$�p�����!�� r%+��!�"��UbӖ�l�x1"O^�k��ÿ��ic�����(��"O�h��ɲ��jW�_?+�q��"O�(p1�Q<]�:lCR�^� L14"O�����Xax�mS��M��X+"O�0��"hɚ%��@�~U�D"O�Y��i�6r�P�	U?��t@�"O4	v��o
��qN��4$x0"O$���`�i~�q�Q��.sX0@�"O��2֤˴yX���v���z�\�S"Oh���'i(m�F��6��Zd"O�{U��F$�fѲ@�b4{G"OzE"�%	�Z+
� ��|�2�"OƤ�d	ӎ
Z�P@aP*6�re��"O��4�ęBF��(4�,%8"OtU%���.��!r%�DL�`��!"O���dJ�'k�̸�� �lv�]B"ON�1��p�:�DC<�Pv"O٘r��.S6���P+Cs�"O$����F-͐Ѫ����a#��_0mF�@���	�=G���c�^�_ l5��(R�1�a~�I�n2�=f��/d���sag�UB\=��C�a�v�j&�J;t�(H5�O@�O�Q��hտ"� �!Ҭ��U�9�g2��i�/��~"c�!��-����2="e I�"H	i��VQx]y6)�#S�������a|��C0�2�h?{ޚQ蔪�M;�È�Z��G��O �z(� 8�h�]wy���v̛�D�\λD:dꓩ�/mX��AM)~�0�ȓy0��xqJ�9}h��hʈg	�Y�G�
��ԡ��,���8V ��|7��;p ����4CUN4�s�]��֦&¤J����@1,��$=�OfL�s�H�mv��zP풙&��} ��D&m(wܵ�0�)�H�WB`y $rӊ����OO}����-�O�e�oS�u��R7��t�[��I�V�&\�wi;C�jûܞ��C6x$��*tn=@��s�P�KZ@H:D�K)A���kd�Y?'z q��E�d~��³L�&��1,_�'��8�7"Ŷ ƌr lӆ��Q!�H����Pn����<J�]�/�P�fe҄2�����}�g+[(7�� vF�pp����O8H��n�02٢��Ó3�B�(�$M�,����nxL*��ԋF�r!P�� ��f�0�J�hشSW*z����59���$F)�bL#�Q0Rp|[$*];*����4#q�z�Ί$jq
��Q�XN�3T�j���i�㖋)�U��@������8Hx�n��FSf1Un�5r�����I�?Ic�w*t v�˸6)Pcd�o�*�+���
��I�����ҡ��}AP�;bx]�DՆ;ZhD����b���	�|G\y�%��xAXQb�HN��X�7U�:XbX�gD�g��I'8o���pgD	L	D�D�R�)���I<uB�ЄP��;�IN�3�1���w�Ϙ4S���g�?D;�٧)['n.y��%��M���G�<�&M�D�̧޲���F�|�|��KΉ|����b���Q���7��<��藿i�Z��@�S�\%��eJ"/��Y�4��)~.\���0KQ�0�B�'���X���/��%!���"t��'���H!��/
ĸpl�7X���q._=$���uAW�I��.'@�8�ǽ}�J(*`@΃$�!�ĝ�2�@��$��l��@�% �B��v�\){�t$��H��"�5�Ĩ[&5�j!������ �7f�lR2-���i��p�l`C�H&$��ߊ��`�F̧Gz���۸M��y3+�q��ػbG�9�а���~�f��QnT�~Z�԰��ԛt�P�>�BoJ46(�q��_�#��I8�)�/��TK�^�q��A�2�&x�bϊ53$�E[��ԦY� �S�*U�}�fJӍQ/^M�A��#�D[#CE�.�&�(���Dx�Ks��+-�*�8�L�wij�8C�G��L4���
7��k�:�M3�����F$�O���C�=0*���O��1�],wM����0��Dإ"V8D�#=1R얹#��zǥ�O&�b��'�n�{ҍB6EN!�f��2/\�q�
G�n�(`� D�m֤�"�\�g�f$˦�'@B=�M�3-Z�YJ6
�r}�£MNĥ�ꃶ7Y����b�
�Mk�)	�2�DU�f�OX�c���A���[[w���&�^D�q�R,\M�Eo���� UZ0�"D	���ğ,�S�I1󫂔Q)��([7�PEq���+ş���7�2wT�)����
�L���Jˬ|�� cg�P�Gv�� �i=^u�u�g��򄕘���YdL�y?bѨ��Ԑ(K^�1דY1�[��KTenM�*
H2�)Pj$��A0d�ׇ-��y� �R��\`Q�4	�BԒ`E0�Xn�+Y���5鶡ӓx@v�*�+�j�^ !��͊\�p��="92��4M%�8��,ɷ�,�ҍ@"w�
�ؓ	*I4�A����)�W
��=��➈#%�F^̧9�jz�@
j�$A�/XD,��l-C�Ty3�%);���tl����ԺcfɊ}�� RQeg�uZ�^�]?|)����8dHҀ�a"D��9oč��!@Z�`D���AS�N� �Οp��!F$J/8��5O�����bF�����@*wI�5o�ȝc���#��9t�'N��$F�K�R�2�.B�!�Ü>(v ��U�#W��dMs��$�\���)� �AiA�I:m�~@A�0��d�"O�@�@�WjJ��rf
s�iG�' �`��\X�la�Eu����O�o�<��b�9D��Çe
R�R��K�L5B��c1D��T!�X���`��$z�N��":D��J�#�h�Zu�Ș>&�$BF�&D������r�bɹ��.u���³�(D�pi3숲T��E�!�I���hA�:D�|�"�
&Y8l��Z��]�8D�s�TyN�²�H&4}̌���5D����f�u�J�8C�.J��b�"0D�K��B't�u�@B�|FX�"/D�l)%��/���C%O�j�0@K>D��z�kT� �Hk�_�Ihn����!D�p���-��g��"U�P����3D�<���7x�ZhB4�Zr� ���*4D��a ��(�&q���o�i:I4D�v���[Ħ	L�xa$�]��6C�I�D��e�e��_�(|@���I��C�(P�֙P�kSO�*Ӊ�1�hC�Ɋ5~��u��%8a& ����<C�I�*��r��J&e��a�' R"C䉇s�<��q��x�� f�y��B䉕YV����AR 	{V�&���m��B�ɚ,j�b��67��@ �����B�9k��	c'��M�Δ�&.K"�B�IPi�k���5\���"7�	�_�XB��,{s�H�b��^ـ഍�(�JB�I!0��ձVG�#tā�E��(\B�ɬk0��e��̔E�t>�B�I����4D�]�|�'��B�I�w��Q
��5&�Ly�����kR�C�iɰQ�T�kZQ���9Pj��"OB�@c��hٺu�e�P+Kb��A"O|�1AD�l�z��"!��ճf"O� �D� �tX�FހC�N��r"O�����X�U��屖��p����"OĨTֆ�|d�R�C�HY����"O�|���Ύ&�H��&b�5ad���"Ob�(q@٩T��e�L*=:��"O:���"����Š� �'Ba	�"O�E��t�}Qag[����L�H�<QT˙<b�J�����|��ًu%PK�<��	T�T��W��3_�-��N
h�<���A� �xٺ�{Z�)1\n�<yR%ϻs�"-1�T�B�g�<�`/Q�Gg(�3��м(�0�6��a�<�qK�X �����V%JA��X�<I4��<���31�]�|��A��O�<p�֤ڦ)��#PV,���K�<i�(W�["���E%W�)>��ȓ_P��P������;w��Н�ȓC`D�1���-����b�����Jh��M���c�]J!�ȓ:���"�f�
h�d�Y�	�p�:���Ch
D@`�[��Я��-�$�ȓ@��G�ХOw��TF�� aD�ȓ.�f<���U}��_Ȇ1�ȓag@�����?�m��Ϧa����kh�p	"c]��Ak&O�ހ͇ȓk����V�W�#> �kP�zCر��b��t���F5l݆�2�h����L��~"Y�.�9n����Ċ�m&<�ȓP�A�U�Ք��Bp&�8�N���S�?  l�g�;O\�SO�3x�$؁A"O�qacո7�����Q'�J�҄"O���'_1I����F��VN�xzB"O����EI�5��iw�"WO�yb#"O8���q5�p#A�9),L��V"O�X8F��gB~���@4r72���"OU��\ޘuuZ�Z&4��"O�J�=Ђ@� 4}B{�"Ot�����<����� 5P���"O���"�ӈ6` ����+��u"O�5;���RN2�I"&�+r�j�"Ol+�˓G���0��͛Kk\8�"O�q�U�P�C$��f�	u�^��U"Oh-�C*6@zA�L�%�fP �"O�	�m_U,"T)&J��
St��5"O���ং	^��R*ͨ@̸:$"O�@��$ժxh�a��2V*���"OnTS�Q>�)�JT6eg�m�"O�!(�P�J�Y��E�[a��"O��Y$)�*�ʈT� �mIX$`3"O&���)ϽoUz�bL�!���g"Oj�q6����҅	2`�7<�8�"O�uc@+1��TaR`�&���"O.���@��)S� x� �|���"O��L�9r�2��A��CG"O����&����ͼN^L�"O`�VFYcev�K�~L�	�"O�(���w���
�2~Qڽ)�"O�UbF�(2.���Kޡ1�6|q�"OZ;fhR
/Q�@ܸ/��9	�"O2<T�،m(`@�
sY���"O� ��D�Ma�H��ӣ�IV"O�@��J���@Ȩ�nE�C���sd"O(:#)G�+X�8�MÏB���"O���h=њ�ڝ��%��"O���6��+CY�D�@�!@�~-B"O��)Z�r8|��ԊF�ㄩ�"O
EpÆW�zo�1�T8G�aq"O─h��0����?j0�c"O��)�!؀��ِ�f]�p�"O��T�R�i)p<�n�.=�]��"O0�����Vp��nG�K�d�)A"O VQp,�A��2,�>Ek��g�<��k��OJf\��.×ad�	c0GA{�<�D ��'�䝚UDr%�U2�)L�<��A�	
�bǈUDK�8r�VM�<��l��G꺀[ѧZ77�ι�.�b�<qe�֧IR]:�P�V����a�<	1�W��.��B)��q�O�X�<!��H�	���7�AF�Z�@�[�<��ϑ1��)�����h��j�<���M�B͸��Q�F2I�"�x$�y�<AS�,39�1����Y^d��&"O`�d@U�P�)uȋ�+��A��"O�xr&�ƿ��MrtgǃPC��ab"O�a��5D���(NE��*�"O6���
O\
��hӮe6�|�"O� �r� 0o�Ms�'R=y=v�3�"O¸�w��Y~�u#1F�3FV�"O��c�+T�ф�� �|ʐ"O2�Q��`A�a?x�Hg"OP�BLD,oBL1k$��F.�`"O���hڬM�tX���g��8�"O6�[��#���"�'V�r���"O� �@cwi�;��BB��+n��DP�"OV%q`gN�{��z�jZ̞d��'	�d0�� hG��4��;Z��]�'w�� +�m;f�Q�M@!"�Tz�'fJ�3s�v�T�P�T�4�LK	�'��*@�	$�s�a#���'�6�x�m���˂[���'��@ۤf�f؊��B��_8n��
�'`�e���4j+�m�,T�e8��J
�'�~ؓ���6~�����H�:W�&�:�'k Ͱ'/	6Q��0���/\̪�'��1Ta���8���b�-'K��c�'_\����3f�hb�����Q�' 1r퇮]�Rp* ��U��'%�xEL�;�����;-m�=��'����Ce��A3����D)�!�'ˈ�*��u���e��
6���p�'ABM�A�+m<���DT�F
����'�$1��^�#�~z��R$4BL,J�'�NM�VK<*Nj���ڗ*nzr�'�Ј���U�y(\�cB�
���'ۤ����7�~A�q���	���q�'D4E�+?���irH0��
�'t�1-�� �:��`�(�N)��eQ)$R*D���ݫP��xPuH9[�H	������0?Ad�W
4�\��wN6��M��� a�zHI����t� j^�o-�	�'�0�'�(O8d��	�7�:M8����'IV ��]>hj7��b?Yפ���>x�Zw`^�rU�f}���W)�953�< �ŨUðTY��X��0>ij2"A���ypi�O�����󂆥+� �"�'�����9/`@��	��#��|��� Į�ȭ,�is�ӫPh�C䉞0qƢ�qÏ��S������_�A�l[2��8k�4�]nBX0o�}h��9��p;U�����#BT,b�X��'�d��	k����cU-����g#�	B���w�G+2N���+��|82�� �i��8��_tMc�O��'�.,����BD~	�`�Sj0Y���B�B��M �?Q`iK+3�4�*$!ѝ636�b����Z�<�AW�*p8]j��)T�����K���(r:���Ԛj,�A�ӡ��"�����F#I�v-�1-s"�#d� JT�ݪ3�L�ҷ���g,�/0�Y���8��a��Y�L-G4:p �ϋh>��i�'��� a�dT�Q�4a��=S�T[W�����*F�MT8�s�4v����iǴxӂ)�
f��9��1AI�'m��%�B s�����'-�HAA�>&,U�l�OP�$����@����r�43ȬXmZ����GHTߦ��@�OR8U��@23����ORm�$�DA1�K��/32f�ɅU�"�CGQ?����A�$��\ws�iꑋT5B!�02�^���-���L]34I�`j��Zo���0<���H)E~+D�GH1r'L��<Y���cC�˓Y�682rj1��[�& B�*�}� A�@���fI���S�<�Fu�wO�l+���A�v�)a�Q.Xx}��I�@���Hdk���1�.x��Ȟ�"D�s��Y'I4�@"O�!���ʹA����k 1/=��p�O�"T(��]�q�I��}ڒ��<�q���ׯ`=�XNGs�<q�PL%��K��զ12�I@Ih�٪NkpD� ���0<���Hf�z��gn�hR�3vA��<iv��/~�4ʓA���12�9�S�C���A��(O�:t��銃)�P)RL��x�4���Oj83��8J����V��
*�Tmh���0�V����i R���U��n09C�ĻM����&�'���w4�)R߶X�lB0�8LC���q���[�kF�G�%���K�4�����,Lt �!%�3i}d7��%Q0
���n�JA��'[&��G��2��'`�!�N��ĵ���\�3H�aٌ�D�'3��*'���?i%n�!��L2�(�s �x�/܆2���� ��Є9�@ЊT��q/ȾX�����X����HX�^���Ia����k~�����UY8ݰ��0t��293��]�O4� Xsd̈́\�t�XTlV�h�J�<!$�k�ÏA�j�OlDAT�W3s�ʌ9C��6O�ic���GOf	Cw��4�p��5@�xXitd�p�̬Q�4k���s���� ��ma( 9�6@�$�O�y� �e>�Ջe�դd��A僑�'�p ���ہ\zB}
�XS0�SIg��d0�O�{BJ |H O�Jg�����pC�mAq�X��HO.]��1	�X��� 㺀h��ӆ0~8���>�8�A��V0� O\��� ㍠��y���)I��Y�$I�c��;����o�6M��	�*գ �P��?���P�8y� ir�3�Y; nd˥0�� �`�@�	P��kq�(�jA�"Ot1cCn�q��!ϰ!����@W37�,|9�a\!=��W".	x%sS�O��ɱ~ ��w�� ���fI��AqEW������mf�p��'������1+�w��8�G�DǤikP_���ea�k��~2�~���=x��e�i#h�֢��G�!��_� �;�A@����A�i�RH��2������6�qpk\8.�T�*.��qnB�I�=\M�T��"8_�$C�	��"B䉆d\)Uj1�A����GGB�� �`�c�OQ8�H�* �&>��B�ɾ(NP钑�R?0R��1l��!�B�I�1��s�)_(����"C�	?/��uhE�G
uQ�R��[^�NC��)
�`1����z�ۑ�Tlg�B�	5�ֵ��&��x~�@��/�)G�jB䉮`tVe#6�1:]I���|�C�-���)Ƀ=�u�v��#9IHC�	"�li�G)�> ���V5��C�	�=�"��VN�:@��hԢT�Tk<C�	�jϪ���j��`t�BaWd�
C䉔#dJ5�ӆ۠L�h�Se�o��C�I�c���qBdH1f V���KU�M_�C�ɮo0�#�d��n�h�����EP0C�ɟg�
��A�1Յ
5}�X��5D�ěB�]�j!6����)y2$D�DkE����R��ٚ$��@�Ц?D���u��$�0؁ª:.ج�h;D� �j����a�hU�M����9D���N�5|8̥[�-ѫ-F�����(D�dK���0 "�4��a$D��u+݇Ei����Q*2�yB��'D��j�
ď1��� �,��8�� D��Y%��q$��ʥGM'ݰ؂u�2D�ܚRb��=�քr�.͒x��l�.D��(��R.-޵;Uˌzxf��@�/D�hxR�$%�r���"�+iRV�y�O�	-������
L��h�*>�y£�
){�=)҄�	O"i� ��7�yR�^>�̥�t��FH���&�y��͂`zڬ�7��O���Y��_��y��VL4��2i�~s�8�y�T��D"��RE�dKceQ��y�S�\X�R��V�61����y��-f����-?{<PC�G�y2�0
vh�e��*}	h%!�O���y"oםv؎4(WC �A	XJ�gߝ�y��C�Y� �d+��b�A��y2��K6���c[T��1��y���Ha����T��Q�?�y�#,�,T�3G�~��E��6�y�C�&/��-CN�gM ��S�y��3&Ι"Ċ�>Q�n�P���y��bwL�r�&y1F���
)�y�e
�@Yh�2Q� �$���IF��y��%�頑�E+���&d���y2IH;U.��@�T�/�؉R�y�G1��i���J}��)���y�mR'E���S�X
��f���y��$X1����I]di�����y�������)OKrx��1$��y��@"��	�m_4T���A.�4�yB*�2t B@R0�čN��N^'�y��N���3�F�|B:ɒ��"�yrg��A�nJ��	�p�.u` f���y
� J �ϸX�dg�v����"O�tpw�F C�h�ju`,Bє��"O�|XW@A@E`�<F��"O����h��U(�-�����"O�3G��j��*؀Sѕ"OH����[�nzM� �X�"O�E��'�q�@@(��A��"O��5�&��P�w��.B��u�"O4�[/_�ff�t��IҶ;���
�"O|t�bɅ�'O��+h�aE�1�E"O�A�gOXM�B���	;G�p�F"OV}��5�|�gE8l%\X�v"O�ݺP�H{f��d�l�����"O~T�g�˲ �`�z�Ş� ո���"OHyۅg�ЌyА�֖ s�"O�<!�ȝ<�FqI�o�/y��P�T"O49T�Y�SYVd����$^ܜ�{�"O��2�D��T���孒3l��)0`"O&%�RQ]�u@�ނL��K"O��v`]J ����7�f���"O�TS!�Į&3t�2��a��zp"OB��˔�fUt=S"/J�h�P�s�"Ob�Æ5
b�2t�
�Z>jX��"O�P%�9e(��snU�R%B"O��ۑ�bc��[��Ѓ�p�@"O�54D�$���q���5]VX��"O����÷xl��6M�<!AW"O���-��9�*�#	�h�ȑ4"O�y�BO��\�	DБ�ڈ"OZ�JBk�;Z�Ҡ���L3~i!�"O0�Rq�V<b>��hPk	R"��"O̹tn]&�2*�1���"OF�
���
�l@���=Y0}��"O>�Ȗ�3u�he�*q9�`�"OVUi��ۇ��l���}yB �"O��s��ɴ�(�6ǋ�J�%��"OZ�@�B�h��4z"��>'dT��"O�5��.>�"3%�.�8[�"O�1ScN��d�ہ��<+����P"O�IB����E 6c�=d�6�h�"O���d����Qdܝ7ն�Y�"O��Z��?/6iC�䖀m �i�"O�K'l�-)@�E�7�;�"OZԻVΐ;�����g�:@���'"OLU�Q���460�15 M�4*@
�"O�eѢ��C� �aQ�" �1�"Od ��)*������WHiH�"Op5�o)*�(���>9�ɡ���W��ࢁO��-!��1��e#§~$V����."!	1��6Y
D�WB�{Q�'��ç����%�L X7�H�o�lmѦ������Ҳm�A�@�(��O��T�p���cZ2�(�Έ`>ƍ;�'Fj�0��R�l�C�>�|n�8s��P���1)<�P���H8�t�#�y��C�u�����y���E�h���ۣ��|�͡'��q�\ ��_;=�1Oa�����"���!A	�4@$��	�X��� �y�)���0|��3��DeOR�8�3�Qg̓S�<�#�g>5pu�H�"U����C8����2?��Yq8L�<E�\r1���W���k� ��pF�͓8 n%piKy�S�O�
`JبH	z���,��q�QZB��L�����JJ����[�;Uڹ�g�m� ��iH�ѳC��{؟`@qJ?&��9zr	�#?��*�'�"x���z*���ى4&zd��'{�P�� �9�6� �̀)U,�i	�'�	�T,C]�����'>Z�0	�'
�:��.s��0AU`8!R�0`ۓ���� ,'�	�J0+��Q�-��h�`"ON���ʜN=f 3 �����@"O�	� l�v]䨲g\�� p�p"Oh��Ū�79��FM�ܚ�9�"O�.�D��@��HL����J�03!��Y�B���5��<IBlG+Հ *!��éNΆ�0$� *GZ�:�*U�y%!��%HT%�5OF\*��re�/�!��ԄK<���ϒb%��c7�ȤM!��[�9( `Һ+z֔�� ��b!�$��L?$���kg�,Ko�"�!�$�Pu�mJ�"�3�8��[=g�!�D�q��`�B�!F��;�g�b !��W5L]6y��Aû4��9F�F!�!�РI�|DB�͢E D�{�FJ�Q!�d� ����rJ��%�T��T�4!�d]8]��3Ua�\�Np�Q�ȍT0!��S�޼��Y����UӾp}!��G�b6D�C7�	������ 4�!��#7-<�(0�@;�j�lL�U�!�
�U?f�0G�J�r��٢��Y�!���� ll����$Wb�9jm�9�!�đ%[@��Ȝ�R
y��̒�!�d�[�� �H�2dC~L��+]�Y�!�dտ@qX�z�
�(β2���!�ć� ��y�����J!��tʗw�!�=I�	bc-J�`�l���I��s�!��!FjTl��.T0s���S)�/�!�D�-~� i��z��,q�H�3:�!�d?��|*���Pn�,)p��8�!�~�n܃&�F/e$)2@*��x!�D�0r�xqjP� �
�xH�'!�4���F Ȉ	��H[�&�c�!�6JM�� Շ'#B���J���!�DB�/�\�6��#���:w�^�7�!�D�;W��r2J�9{��D�N�!�$H�sXB$�C,G�mq����֟0�!�DE�8�� ��F�!н��V�0�!�$��M� #(Ee���f�׃v�!���(���
)y�h$��O��4�!�ӑN�vy���� �R<p&ɘ*I�!��D ����$�	'�=�ɐ��!�$����ʑ���<[����S�!�$�S:�����	i�LX h�-!�ٟ.4mBBC\�UzQ��h�&.!�ݐ%����⡕���"ϳ!�L�f0`H�b *�M0 ꌞ~�!�(n"��B�֥L&���ƣQ�%�!�d��ef�Qe��HlAKpC�d�!�$4�b�r��$Od8�s�Q�+�!��~O����[R/vi�`�!�$�d������]<D�rW(�//�!�䅢Ъ@��S8p�x��L��!�D�5w�m��z��� !,5�!�>T���zƯ�!������F�!�D��fsxD{��B�:�Y�!���h!�d�0r3�|cCN,{&.����J�$�!�$E1q0�&v�T���6Ml��ȓK�ԩh��E#C�F5J'a;h��P�ȓ;�Bh�d��l�\�Ӓ� O����H��Q
C�ԤPoXVbw����6mt�Ҫŵ"�iq1同݊�ȓ6��Ѣ�վ��D
=�d�ȓpF��H@`�O����CN6$%r���S�? ���Q�B�dL���4I��@��"O��y4
-p�4���-@p�pp�"Of����#I���3�J�!��mc�"O,��B,®���
�f�y�Nak0"ON�Յʠ&R䓵�tЎ���"O��Sa3H�|���HS��bC"O�P�@E�VQ�d��ȏk?(��#"O�����C��\8�%�n/�]�g"O�����ۥr3��;&�S?#0\��"O�����ΈdF(x��� ;l 8�"OHp3"��[ƬxY��,`!n��t*O�Y�V.ǉ-(�5�X���@�'^ȋ��VXT�q:���"�t��'3�<��D잰J��7��4�'��@���эf�����w�@Ac�'#8�e�����կلe�-*
�'�*M�DU�uG�9hdD��j�:8��'Vд��L)5.$�sc�b����'�Α���p��@*ca� [��B�'2��Q�Z�(/@U��I6M5ƈ��'QRy �IYBj�!")�W-r��	�'|>�9R*^R؀���d�n%��'`V�I1LA+6^d4��I[����'���(��R�8~t"�"�=��h�
�'�����BJ�n.T;���	���8
�'Ί���B�<	I�`&ǬP�vt��'�,�����$��i`JA�Ozh�J�'����`��W�$����2��#�'���H��Ѿ��X!����x�'��i9����I�C���N1��'-!��bXv3X1∌��0���'ɴr��if�)p�M���"O$�hS�M]��2�Y�(jM{ "Ov�(����n=뢫Y#$�p2D"O�xBE)x �ɸ�@�*
�-
�"O���E�M;�z�a�O�:�	��"Oљ�o�[.dy�H�##�v� "O�8�#��)'����U(k��H�"O0�kGH�"?�q�hK&Zr�p��"O�Qr,��.!�F�VdX�y"O���_-m�$���
=&Q��c�"ONqa¦�0|��H�$b9j�v"Ol�JV+Z�6E�A�hхAx�q!"OL!�v`	�/+$���&��B��*O4��4G�Jz��7i\0��i
�'avI�s�ްE�6��@I)��U[�'Ґ��ׄ�)^M�ݢ�˲���'@�t� ��,&,�I�tM�<��'��A�,\�~��$�N� �����'R<e���?"�	a�$G[v��'�&�c4Ȑ�4Àei�aJ̐��'D����"цP+T��@�8n�H�+�'�&L�DP�tJ���+R�sv��'Y�r+J�/�^{����	�H�9�'�Zu@ᜠ@� =���Np�9�'�h�
���%�
�X�D�(��w�<�f�K$0��[Q��&$n(�F��<��	FI���P��!�:ɠFoD~�<ɴ�B�Kq���4�M��y�ī�P�<I�I�,PjIiP�F��r��c�<�bmPC��1zP�y���1g�J�<1��Yb|$E���j��8���_\�<Ѧ�D��=g�ȝ���c��Y�<�ݩ2K��2.��X�dp�<� �����	)��&x"��kc"O|���c��]yxŒ�%\
>x�"O��7�ł6f���M�4��q�"O��ҩ�f�0��1�\[�p���"O�m� �!�.	�K�=�TLr�"O8P+O�cO�	 ��čs��l��"ON�Zs�՟��(�iN�=;dQb�"O�cb��iP	�Wm�
LN�[�"O��r�mԆZ������ ��Q�0"O�:�Gέ>�Є�AI"]��[D"O�x2B�ӵYZPȰ��\�d�� �7"O�`�W�!8��`"� �.t��t"O�$��n[i�X��)Ѕ ^,q�"O�XQ.�#6p1#n@�T�"OX���K�����B��Y8�"Os��X,ri4�;v���lr"OT0b/�FV�<*'�Ȱ>w�Q"O����*���D "U�IGo<	�"Op���öM@�;�'��ɸ�X�"O��6�̅*�u����5Ra�%"OȘ�b`G=P��<�"f���$X�"O����� ��h�K�IBq�"O�DBHV.Sz�)��
X57j��'���b��U�5�,�2*�,"$(�'/	��l�f᱐ D��X �'<��y���m9���,F�GJ,��'S�8���Y� �f�:��^9*�����'�2�1�����)�)��y���'ބ���dωk���XxRB�'t$䡁�ܔoᔸ`4�˦kU���'�Q��F[���`��*00��S�'��щ��ݣG������#��9Y�'���pSċ9d�r���ܹ]f��'���S��֮@����t\��'�Z���� ՓAچw1H@z	�'�rm6F�*4�Ȓ!. /r^�	�'V6�" ��$'*��&�m�Dc�'�����P7fU�J��DK
�'�j �B�~��!���A"+C�h	�'1��	CCX8U��d�#�K8M��A�'����� ���i:(��'f�%��.�^L�����;�L���'����  �x/L%b�K2H��h`	�'K���֊�P��qkrFP�����'и$a*	�e�~��,���XY	�'غ<+�h[�"*2p��N�w�-�'�������&���P�T�v�6���'p����O"l���p��5
�'�D	�g��u2���� +����'���`�#0���q��wФ���'~mE�اW,FqIƨ>n��}z�'P�a���R�@~�s�c�)9�'�^����]W��rլ�Zy�x��'��J�k[��v)i���=X�~@	�'Ȑ�ƉD�"d�c�(�C��lj�'���+��[�,"d�����)5~\��'j4)����Hhj�	���e��A�'�6PK��>Bz���q�B�= Ԉ�'^=�6�A�	|(���E��&&�X�'DT��(�o���pfKw���'��[eG�
>Ͷ4{`��>���
�'��]�Ec[~F\l�/�|V	��'�"<0��O�Ta��ħE���'Onŀb�F�G�d	% ��D��)��� XM�&���)0"Y���ۄ"OVp0GJ�8i�]�jD��P8H�"OdQ�n78Yh���X�L8�"O�i�n:�ɑ�L7����y��)e����Y�9cA�]��y��\L�������LbqZ"�y����%>l�ص.H0K���Fӆ�y�*��)""<��l����	��y�ϣE��""
��I�Glͽ�yb�E>P(��䌂j	4��a���y�fϯs�@l��oG�_S���I�%�yBm� $��  �'v�U3��yB�VCR��b`(}�&`"�(�y"K�=   ��     
  �  S   �+  �6  �A  �J  LV  �`  (g  vm  �s  z  ]�  ��  �  '�  j�  ��  �  3�  t�  ��  ��  8�  ��  ��  �  ��  ]�  ��  ��  ��  < �	 7 x `  Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�� |d��"O
`�(�;���8���-0��1%"Oj4��ND^[��"3/9�0|H�"OB���H��*�ʞRy=a"O�味V�!X��!&F�:J�$���"O,��a
���C�Ą�M�"O,$3%o�-���p���+Ն�:1"O��ݢ1����`���y14]2��i�<�6��{_���c�H�`�fX�$Kn�<��A̼VI�xR[�)�Ć�pඤ�ȓA5��('nߡ4�� �)˩%� ���,��r�؊b#`T�eT09���ȓ!�b��g��}�8�F��-? �ȓ
K|m�ș�VṔ���2�%�ȓ"R�X�j�4JN�1�˘X�i����̹	_�jZ��1!g��zܶ��ȓgil,*�J�
j�Ne��i�J%b���f	�(U��:���G��$Y^م�~r�� S�%T"���k\�jx�ȓ|4�1�îJb��@ӵ�ݩn�V��/[`�"�v4�R�!ʎ<��M�ȓ`:��z�ؚh�J�Z��$HY:	��H��p�m�C1��!��B:��0��EnjZA V;9����J[
2���	��4'J�EA�IVW&��~�(aZ��ӹ�>� o�Y�|�ȓ�f�A�
Ο7�H��M�$�����mޠP����/���ANXo*�ȓTv�����{ ��-7�*h��I��sB�8�8���3����ȓNe*M�悡;������X�o��!�ȓ'lj�#F�m�+R&;�|��2)n�C��0S4���T:
b���:�0!��e֊��)��ͷV��,�ȓ0�&�8#���� ع�L�����;�P�AFd���,w�6d��r�EQ�( �gVlɦ�M,H��,DP���|�I	$G#\���ȓ"�)���E�B	yt&B�^�LɅ����$�H+q�O�����(Sp$��&D��)d�8Mʂ�s�d��<Cb��@ ���F{��)��5��1e!_�UU� ���� �!��	F�<�qmNgL
���1B!�dȥd	!1��.G�ISl �Q!��ɚa�h �"�;XϰM���N�a�!�$ݛ>8%
��05� IB��
�!�B�M�(�#fM4	��uP��!���Z�B��iT�x�cGM0�!���(�P$���!� '�p�Q�<���Z����-Lm��9q�N�Z�@���	��4H��ցK�25*�@7h~Ry��-�$�j����,�����3-�Jɪ�͑,C�ڕDxB�'�R`c�%[U*5;���`t�HK�'`hPS����#���+ڛ~P��zT"Of=���3La��
t	��G��6�	z�Oi�A�+ZB�X� ׃�?na[����0=�v#��P���y��H�6�V�3�u��7��?�ϓ�����n��y�`ܡ
��0 ���!�הG�x�'4|����� 3)�!��5/�$�r��0X&�Aƅ �Q�!�$_� {Z�����
=�e�T�ݸJ���x��)�	\f
�� %^#δ8ba�6H~�2����?� �%��D^��Ճ��Y$<�j��*O2ac,Īg�ܳ�L�.i[z��
����dK�!�:�5�J�e�"-H��%�!���\z� ab�Z�����N6[�ay2�x�U�(үӥ#� ` �ӈ D�g�,D�Tӕ�R�'L4��U�R4eM 6L,D�0��I�]J�bԭ0-��tRs�,D��1��/6�ļ�2-�<(���:4%8D��pV�~\��s�6YҖ����)��hO��L�x݉��N��I�%G�(X�B�I,\b�a!�E��z�R�����0@�vB��0nt�:��۾ED&�r��J�",C�	�3-�0�ˇ�2�.��Z����hOQ>-(C�\}˶L@���	^����,D���7��F����(V��
R
0D�[�c@��V��S\Ӭ��L.� n"�,��U�S��X�&/et듦�=q�O$�W��y�j)�b�Î]T�l��'����O���O찡ժ�p�h�
Ǌ�:{� ����<���ħ@�n[ժӪ
R��sjK">O�O��I�����O�Y����[T���U�F5zX�X�'��:��$�'<a�ј5�	A�l�zR	W�7 �@�=��d�zС��1�8e�t� a-�M<�O>��'�>9Q⃼z-��
n�k^H��G1D��G?���3�-��0�d�>���<�L>��y�&if�D��M�2��E�Sܚ�yr�:y۔��6�`��y��+ѻ�yB��'�����G7bl�p���yRD��4<pg@�A8m g�3�y����z�ru�h��HO֬�@��y�$�3s`zL�@�Ŀ/H�@G�ג�y��wӾ���ˎQ��%���	?�y��ެk�2�:��(NthBd�N,�y�Ƙ�u��Q��43*�A&�y��T��\�5��&�x�r,�%��!�S�O>�0�V�A ����`�2N�T���'�xj�	��H��
�&��8������yr�B�CHre��KA�rV���y� �
8���H�Eo�݈���y��:PԀI��A͍޾�����y�#Ν.6��bt��(L���bA�QqO�HR��Q`�g�	 ���qꗕp[B�XB�[G��D,�ɶc�b}r�V�b|�(Z6*�m#�i2��0��˯(�� B*e_t�O0�I|UQ��O0�$�#�sN���Wh�&�Vak �A��p?i�43����@�n5n�s�	4?)������'45 �i9)�^�Iƌ��	Ó ���H�]��V�b��BR���%��j���S.-�`}8f ���1+���=�"�'b����+bI����Fڳ
�\H�S
_�w �l�˓+�z�ŕ6�LX�Ý._�h$�܆�	hC���w	�P�^13ƍ�V6B�	�c��ص��4h8�;��Lm��"=I<����Aҵ`�ά�7e	�[�ܝ+���y��9,1V��!��8B�C��F�铪hO��L�@�\�t�Z���ϐzHĂf"O���,["y�Ek�#3H\�b"O����s ��R�A�h��'6�O��z��U?a���h$�H�X�+D"O2�@g�|��x��<fN�9�T�?�S��y"��Fo<�i��B�D��ۑI�y�$�jz@� ��(qfR �G ��zK�ϓ�1OB�G��)�fIb����8 /�pl��ȓ`$0`b�2lЁH3描#�J���S�? ��H%,G˔DВ���>�-c�\�4&�$F{�� ="�oT!N0�@ςk���B9D��c�EO�Vc������CǨ�[������"�\��+8��}�  ^%Y!�DJ
^���#���b|\h	fOͳq!�V�uX)�;Cm��A`��S�!��47��i`1��}d� �p	?�!�@�C2���C�U>d9Z�֥2�!�DCy���mļ@�}���EEz!�DQ�4U�)�Q��d�TC��i\��?aH>!�˃cM$9"�O)@ظE�Ǖ~�<�&M߅D^QYpI�e�샒�@�'ўʧjb列�� !�L�Q� "E���削�O4Л�@����Xc��)��-�U�i�ў"~n�ZH.x��K�݂��$b��R�JC�	#J�rw킽HZ�� �'Qzh���0?!&��  ���A��IfQ�Ry�����$8,O8ReΈ"W{@�y!��h��8XU�	$����3S|����Ŏ~W0�)�JТY"�C�	
2��`�4�&gY��ّ-��2Ĉ�',�O~"}��}~�)�� �8�T��Q�<��>[�,x@O��v�)�C�P�'��x��wn�����%&r	`�Y��p?Y�O�-rv�]M��"s� ���"O�=բ���Z0��.NRQ�'��_���'S���C'&X� 6v���@7U�!�$�	<k���%��PzX*��ǗmH!�$D	g���c�
=NF\��ċ��:<!�$C'%7�J��Y��}���ǫ|[�9���dǹ2'� �vdϬc�QB�O
Ha~�]�LSQ)�zd։UR�h)D`�pI2D��P�H�d�:������(�܄r��/D�DXv
�]�ӗJW F3��M.D�dJ􍈂�~�2�'��8ƺԙb'D�СD�V�t�Jdʇ��";%Nԑb�#D��@�I۶BgF� ��E�o�0����3D�4��'\��=�&��{��1��5D��×`M/{�y�BJ�XYD�h#�8D�s�C�.:��I�![bn�X�O$D���k��-���[�ѴI(�Bů<D��a$Ā�n��R�
�B�%��(D� !�,�M.�Uz��G�>�Ĩ�J#D��#���E�L�E%I����!!D�8�!+7ip�iAǔb-Y�'/>D�l�gi�z~h\�w�9A���!�!;D��i���)�,��֐fg���$D��(©�8b��4����^k�A ��.D�<jg�îs\�m���[�x͸�7D���@��r�\�r`+Ľc�Z����4D�Xb2/��~021��4?C(y�T�3D��z�n� �іB�g9b�e$D���D�M�$E(pz��_�T��z0*#D�lr��c72W�;N��Z��[9�y2,�i�$h�D-%L��H����y���$f.@�Ąב@T���$	 �yRo��p� ҆Y���ؑ&�W��y��/�^�I��qtm��Z �yL������)�5��bx�M0�'�n� Rhɍ}�ZSˆ�Z�����':@auᐏkD�	N)T��'�&uA!@xP�@�$ڸ!�$�+�'F��[t	Y.����<�P��'K�L�	G�b��� ���'��p��c]1z\إAE̍v�(i���� ^q�R޿#�{ܼ��B�5Z��ȓrw��wK11��,	�/'����ȓ��C$�6 �CD�(4��`�ȓe�Υjt�z&4���¨?S��ȓ]zz���A@E�RA�Ld,�I؟\����\���������p�	�,�Ɉ6����(����43�V�NGV������	蟈��럘�I쟐�	Ο0���t����j�*"��R�8),Q��֟��Iϟ��ǟ���ğ��I��x�	wAz��F��(��F�'�����ꟼ��� ��ҟ8��ğ �	ҟ8��<}�\��Q˟�n�ƀBt�J��	ʟ��������۟��	��	џ��	�3\��P���}���8B S�)���I�H�I؟H��ߟ��	���ߟ��I�Jȥ���Q��r@F�J��'|��'R��'�R�'��'v�'IL����&	��Ւ �Y�@�,j5�'k��'�R�'��'���'�B�'~�!�Ջ�+ ���`KF�� �'8b�'�2�'��'���'L��'6�y��Z1�j����c�&���'���'�2�'7b�'���'���'���*�)�_��e�S
=D��h�t�'���'���'0"�'�2�'���'�<e[<;Ӽ�*w(@� �]�S�'���'���'"��'��'���'� �з��E�Q� ��6S��a��'���'���'��'���t�~���O���#��-=�@�b&�lV��٥eYy2�'N�)�3?Qb�i��e㲭�:P�@���_>�����-���Ԧ���n�i>����[�@�s�ٛc�
h2 ���0�M���j�^Y�۴����9*�F��5��/j4Y��)B�#
<y�᪀�`b�b�|��[yr��-}�Щ�K�P΅c�AI��$=�4"U�h�<	����&���w�r-맭�2Hմ�jƯEN�d�O�7x�����';X�ش�y��vXX@�eY�H�2l2t'��y2��S��#�*Cvў�SП䘄	M!D)����k֒e�]�g�j��'J�'�&7�j�1O��yӌ�2[�6��! �2v�%�գ�O�Ol�'�2�i|�$�>y3J).�pi���$N&�ԙ��KN~�i�J��������OO��@���V��I&E� �
�KG�I���2ӥ!4%.`�'(�I�"~Γ|�,帲/��I"�a��I�vh��Γ<��&����$Ҧ���h�i>������� Ô��v�{R³�(�IǦ��	�H��nZI~��B^���XƏ\��*DbP) �j��a�jiڝP�l9<�48ж���`u���<6��d�B�ͭF�����q��pҦ���œ4ߜ���-!HLE�Á�W*��2K?1�j��BE��ctD�A[$7�\CB��<q<�	4O!He �5ch��r�ǥ,e��w��� g �$cD,*R S3@>���I<D~P���¯81j�c%��,F�� �@95���hஓ%}sfț�Z�5��$2 ,
��)2�愹3D��9��K/��(a��/i[([��]�υD(0�1dh]�4yp�� ��tAPa�|M�2�mg����O��$�.��'��A���1��8Q'Mϫ��A:ߴ����;��ꟈ�i�)x�I²DS6!�aN�-��x$�{�x8 b��I������	�?��L<��@:����ı~�
�eK
�X��m�u�i��d`��4���쟄���w��t�3���R(�Q���(�@`�ܴ�?Y-O�d"�B�<y-O6�D��l�D /� ���j��=� A�V�	��'W����I�~���?9��?I"c�O��	��C��r���f� 3R���'L�"9���O��!��Ƣ,q��,j�ؙ���O0;Vś`P��1�1?����?��?	+���S怠2�n���
�,.���X��<|j��>9������ҏW�(,r�MR3��MR��l�*,k&�D�O����O&���O@�"�?���I'5x �"eկW���3.w�6˓�?�N>���?�"I�F��o�"�2Q�@�$�L���%E^\��?!���?�*O�,b�Oi��Lq�A�+����k(6tHt|z�4�?�I>�,Ox������12c<�@'m�-��)z�l:r���'���'�򃚽df��'_���?�C/�/HV��#D�[�=<���/����?���X�
�&O�S�F�)E�#,nĐ�S$dInZPy�,ֺ6�6�C\���'-���.?1���W�������I�	������Q�'�
Q�����H"H$\�BO��0?�p��/f��P&,2�'���?!��ԟ�'b��bF�	�Jdve�ee�7ꁓ��f�&�prl3D1O>���%&+��!��(�pY� I��D���ߴ�?���?�5@�)��F�'�r�'�"��u��XM�֙��.�)~H�
I��M�*O�x��S<U)�?q����	Mm~I����@�j�b�ƾoX�ش�?�� �./@���'�2�'1��~��'���p`��kc�|�1��f����O,�c5O���O�d�OL��O��䓡X�*�`�V�gK�� ���.@������Ϧ�����I˟�������?)�L�-t���D .
d����u�l�Γ����Ox�d�O(�x@�:�L�{�`�K�Hh#���4����e�i$�	ß�'%b�'B.S����\�G�\̣#�,��Yk�*�0T����'M��'��Ħ1�	.&����4�?	�B�&m�!�� ��D*�.�)^�r�1շi=�'2T���	_�H�SQ���]'6�Q�&�vHcfHJ�nY���'��'��b�iSH6M�O����O�iՉz���`V��,��Z�$�&��em����'��E���t�'|�i>7� |͘����yv���/CLy2'�i���'��xshӨ�D�O�蟞���OX���&"LT���4�;-���@@fNA}b�'i��ҕ�'qɧ���~2ޠn�@J��Ms)�� ��ď�M�Te��ꛆ�'0B�'_�t�O)R�'>⣛�)��|I��֚X-��g�>/;�6�ڤ���$�O���|BK~
�lwDi�%�zc�1y��ׇp�V�1w�i���'DҢ	+?�7M�O���O����O뮕���Y7�_�#S�Y=��F�'��]�	b`�z�����j���O8�+��U�yn~I�A@]'Q����E�릕��,�H��4�?!��?�����v?Ac�I�a�2=s4b�#S�PZ���}}�Ǎ7�y"U����ʟ0��ԟ|�	�}����([ T;D9�a�B����0Cݿ�M��?���?y�U?�'_�i\ bRN��)�J}�̲d� ]���'���' ��+B�'xBY>U��G���M�r�p$�v-QU����cQ�n�v�'�2�'���'����r�lj>��O��2��'���A^p�T��'���P�'���'��Ў��7m�OF��܏Gq�$3��m#`� �Ń0ʡo�Ɵ��I�\�'	��4�'����1�<�#���_�L8Cu �!Qʛ�'���'�rHd�H7��Ol�$�O���Ʃt?tAi�n1�����$i)d�nZ����'��͉�����'��i>7-���\"@ɖY X�C���f�'bD��qs�6��O<���O��i��!+��W_)5�`
@$M���'���V
��'Q�i>-���)��������
z��
��i�VmKa	cӠ���O�d���)�O���O���2�ZD��իF��
���Ѳ�Lݦ��#���%��}�Sן*�l��2)V԰��wnY	�٭�M����?��}k�{�U�Ԕ'���O��pEM+Gؖ,9�.��t�zq���i�X��clt��'������
��ZPy#f�K����{�Ͱ�M��9N�E��i�R�'2�'�\�'�~��Ȍ�� �C]�^��pB�����?j���$�O��$�Oj��O2ʓO��ȫu%�hQ�yq��7i��m
�`Y�&T��'���'`҅�~*)O��D �[u<<�F�E�nF�I��Г0��ě'5OPʓ�?����?I��?Yq�\3O���IV�E���9~(q�h�7dx6m�O����O6���O���?����|�2�@5#q����O�*��$�6�%\/�F�'���'���'E�#�7� 7m�Ob��I1. �Y�a�CN~��Ae�5J��oZ������'�򏄋��$�'b�D�j4��� KΝ}��"��"����'>��'���&<n6��O����O����;����7T��Z��3��=m����'�"&����Sy��M���N�0�8���c%<���R$PӦٕ'����w�v�(5�OB�OOl�j���ٕ�Z�XR�+W�O('���l{y����O��xE����GA�'oC��!x4�i#|�itDh�����O��|�'�r�O&�L`%i��{�,y��y'�7_�M��"|z�S�)�E�x\��څ%�����ic��'�O�=�dO���Ob��p1���`N��xqGR�UTc�܂� )�ɟ@��ܟ�0JH)}<���}��KC,ٽ�M;�m��8��xB�'Zr�|Zcu��rHXi�@��ȃ�c�OA9G��O��$�O�ʓc�$��d�H�{��M`d�زlN�!��Ҩ/��'���'�'���D縭�a�
8o�"�"�i����I��0����IП��'��}���~>���M�(6u¤�bA��`aNБ���>���?	J>�+O��Z \���f̉�*椙����_����wӎ���O���O|��O7f��a�a�����O�9m��q�2�#��x�ȍ�c@�$�M���������O���I�c�L��]�����it��'Q�	�gB�h�L|:���ɜKmؼ��ᄿsp̕�&�"bщ'��ɂ�x"<�OR��h�B۷+?8��"@�66�����4��$�C��mڣ��i�O*�	[~�n��TƲ��t�/T@��{w`� �M�+O�S��)��/�����-���T�(�q:d7MЧ0;V�lZ��8�IΟ��Ӹ�ē�?��E�I�y�� ��K���ss��6���'���O>���:J�S�aG:�f��1�E�~����4�?A���?)�É�D��'�R�'���X3�HQs��x=`�� �\�@�O��`u��O��d�O��$�O��$v�i�M��j�6{��P�4���0�mӴ��͖ ���>q������J�
H�	�TLJ�B'�,��N|}��-ʘ'\��'RT�8QG���ix��IYB�my&h�#�+I<����?9N>�*OJ�Qd��?*k ��H�*^ʖi��*��1O���OP�$�<���R�D��͏$Yp���]�R��@X�+� ��������j�@yrL"����0bCr� 0�������JJ�VM�IƟ��Iן��'�^8��,3��^�،"I�X��QrFwI���u���D;�d�<���Ov�n*|���Xe�nm��n��o�����myB�ەV�����<����00��|@C!ė5�t �[u�	HyB���O��#���=zļjf��_�7�<�懄�}&�ƹ~
����Q��H�����rX��҈	8N"Yfv�:ʓSqLqDx��d�*�FD`U� m�| ݺ�MK���p��6�'��'5���5�I-]Pͱ��c�A۴�RmZ�4Z�Ex����O��� ���'��8}4cwnǖb(�R�i��'��/���c����n?1�+0�a�o�1\�n̚�*�G�g*�<���?)�z�����@��B5��*L# ����t�i2�a�TO.�d�O2�$�<��"�41�Ɖ1i�
j4��!�!�'¼);�'r�'���';�^>��� ��)<z9�&a�9��xSlބs�\y�J<����?�����<��䖸x(�0֫�6.V��OO�v��D�O>���?)����DT�x.
�oz�9�+ڵz�`d�OE�.s�h�F�>���?������<y�o�T��l$I��ٍ		"�J!�����O^���O˓z$������<rD��c#o������P�wX7��O����<(OHA1��?�HN��`�K�$��R���s0��nZş\��`yB�V�#���^����cmS�[����;Q��	P�}�m8���e��6u�!lP:ּ��g�z��1���ӵi(��'�?��'\^�I=&�p�3�e�C@��F�Ūu�p7M2�|����/c�����үI���H#%`�X0)%�I�	�D�	�?%XN<��HPr���
�i�HI>>b�=�E�'�2�G<zq��@ԧ�
���8R(�8h�7M�O����Or��q������	`?��&\�x�9`ɗV0���n؞��	����	�`��ep$�x�œ�$ڲF�(�ݴ�?��n�q�'��'ɧ56�L#R�nX�$kX$/���Z��@��OX���O��<IפÀU[l��RKդ@P� �K''�01����O��O��'�2���*9��)W�N��!�}Z�M���?Y-O2�Q(��|
��ү=�x=z���OZ�aR`�i�I�'��Fy��.� ���%�"}rT+����D�OZ�d�On˓�j��S��ԃ˘e�x��TA�t��m��6S��6��O�O��$҅Y��<B0�U��A���ΐ6���';�R���FÖ��'�?���I���!�H�&钅�1L��>O�"r�xb�'�<H�vI�};arEEž0-�Ɉ۴���ۑh%p�m������Ot�	^X~2�F*���� T�$5���MS+O�i�3�)�2J�,���0]�4Y�Ն��d��79g��o��I������O5p�m��;���r�\�P]v�p2�䦕Y`":�S�O���ۊ$����	
t�����۴$�6��OT���O^İ���]�I韼�	s?�U��(s�h�$E<@M��OV�-0�<����?)�0 ,Y�\5v�f�*%�ʤ�%a2�i�� �-Ym"O��O��Ok,T�	��S��7)����
��IE�nc���I̟��	Xyr�@�>���]�-C�r�"��g�6��Q�3�d�O���*�D�<���I�u����h�+J�:`��Ыd���<��?�����̑ �BŢu�h�%�M� ��a�0��/��-�'l��'�'m�IR>��1v�����1�,��DX�;�B��'�b�'�Z�d�d�����'-,�QB�W�7�6h���Ez�x��i��|�R�\{q&%��nB�{�`��^%q��*pQ�7�Od��<1co�4Ut�O�"�ORfJ�=��D0���'.L�����bӎ˓�?i�NU�H���4���bh&�0fG�>E(9�U�	'�M�+ObA��J�M���h���^��'Yr�{с5+�Ќ*��?�5�ٴ�?���t���
���ē;#�Eh �R�B
�5k"]JV)ʦ�{��M��?�����V�x��'�"챵B�=?��$�5=Pָ˷!`�&�ʠ�'�i>c�`��E��yq�C!@��X�&JR�0͚�4�?!���?i�呡%��'���'Zr��r���rQ���u�H�`�: �����1�1O����O��Dԛ|VzAèP��X�F�I��n��dp�"�����?���?Y,Ok,�m�x�򡉉)K�Th0�d��"����c�,��ʟ���yyr�<%�ً���C�nP9R�7#Z]��-8��П8'�D�'��i'�S d0�(e��!^�虢��Ș'["�'ZRV�H�������N�%UN5q0��$�R]�Sf\�����O��� ���O��$7��Ē�V�~	�2/�B*������sØ��'<�'��\�ԩ�D	��'^B�yYQ�A<7��C7!b`u� �iJb�|R�'K�eO��yB�>�b �BI=b`͋dR(�������	򟤕'�|qK �!�I�Ov�	݃>�N i�"R�t�G�Ց.p�'�8�I����t��&��8���RJR�`CB�:D�؉��o�@y���H6MXq��'��T�$?�rn�

�<ɓ�A�Du`�RCI�Ԧ	�Iӟp!�D��$�b?A	 �<�����E���(��r�v���cEܦQ�	�����?M�K<��;���y��,7h4��$���M<e���ie�E�'�ɧ���V���2!ϰ=!��s'�F�v�p�mZП��I՟h�a&�ē�?���~���l���=f���A���M�H>q��37V�O�"�'PR��`I��:C�1VJvM�%h�a#.6M�O�k2Jn�	ҟ���h�i���w�I�
D�Ke�ת[jBU D�>A� �t��?q��?Y+O�)� �x���ׁ�čy+���	�&NY�4Z�'0��'y�'1��'Gܵ�s�	!@�l �Ԙy��R�V�]�8��ğ`�	vyr��"Ɗ���&hzE���H�:htB~���?Q�����?Y�Y�މ�]����5_h.��G��"90QJ T����韐�	By"E��u����Z���$E�f8���ƒ)@�u#Ц5��H�I֟0��-d��s�۞"K��v�,8ܶ���fքG���'�W�L+ЅN+�ħ�?���*K"4i�C��m��-r��ВWX�4ڷ�x��'�BF�y��|���|
pD͊f[rpce)
w�
� Ӳi �ɫ:�˛��i����d��N��'��I�D�����B�F�l"ܴ�?I��x]@���S���	67,t-j�̊�$�]lZ�JB����4�?���?I�'܉'���+��C��_&UzDT�!��*hoX7m�\t��/��ڟ�#�mL�ye�@����%�F�\
�M����?	��V>N��v�xb�'��O�$��E<>|��!�{�T�(a�i;�'~lҙ��	�O����Opx�A�8O��9##I��k\��`Φ�����:	�I<I���?�J>����D�Pd�R�T0��9��@}b��6�R��8��%Vwԕ�v��@��hC�a��u��c c�Mi�M���yb�޽m:�!5mX�u�A�Em)�O�˖�QԖ��GX']����V&��f�z	��d�AV��o��]�D���bÕ�_׌��0G�Pe�u*��ąB�y�JW�3̱h��R�x�f��'МYlt��IV�o�����شEj�gC�#�P�6[�aX��� �҉e���Z�]�D=�U��4(����$D��㷨�T ��C`�4���I��`��k����;w&(�t��'T�=᨟Ε��N���%R �x���)�c�^�����P��O��D����2��C�UM���i��dK����' �̼8wDZcl��Q��kkR�X�>O����9tvLF&N���t�v%�h�a|�I<�DZ�e*���n�J���@�[����h�oß|��r�tm��r��'��	 �i+���g�s�����aʇ5���;%DB�l�B�qu���-sh�T>]�|�I�R���� q�����-.��e�'�U�$�!��Ss�e���P<`�^]q��K�fQa'Z�|�ݸ&� ���gMN���J�	f��QB��(��V~J~ZK>I�Z�.="D�]�T��2�$d��l�0���#o�`K��7(B2}Fx�7�S�ă��2A�A�	��d9�}�eKɎq��'T*�y�,_�B�'!B�'6���ퟐ�ɥ-�䙺pޛC{x#d�ٹ������#8@W�*q�
	���?�=�4�-&Z����&�#+��D��ɨ}����2n���)L,D(�g�'̐��r��c*5f��sW,�K�'�n5���?1����<1���X| ��鏬1�RU�b�f�<	2�� d%��%��[�����_<�������8�o�	�HD�
��p�����E�x�Ԥ����D��ٟD�d�Lɟ\�I�|�H�}�@Ic�L�z�Y&��)|��4�@#�f��H�B(��D��H��I�-ť���R�T�������M"Q@Z�mN�Y��B%X�&����$+v��5���Ln����.?9�k�����4y��d�.T��ŖD�(��aj%U����'���˟�?�OR|�OM�wB�%�2��(xH����'9�᪂��'L�X��X�{QNܒ�'^2�b`�'�剰�t�����$�|:s�Q;� )ya#�5r�f �I�����?Y��g��ȢRB0)�`5h��^�a��P-����V	I��lD@��A)�XA��I�%�x�U�Ĉ���3�FʾyZʧu=�lyBd3N�`X5,[�rǌhFy��&�? �i�Zc?š�+K1)����ۂR�R��q�L��xx��`�4\�h�s �!JA �'�-�O�%���DDZ�;g\�"w�049E�w��)%���MK��?Q-�&Pт�OR���O�}����X?�E�AԆf2<	�t+X�,�l���,����4E��J�R��R ׺Î���EY�A���H��A��7��HX�!ҏ�9�U����ɓ����R�����V��MUG�@�`(��*T�a�'�z7M\yJ~��'��ċ�W%��ႌU�����)Ն,!�V��4%��L�vX�N�,�Tb��D��I4zeH�W�t_:�`
TD6���ҟ�D�8<{|���П���ğ�2Xw)��'��x��׶wz6c�C,}�����D60Y���*5�D�EgC����W�
w�O(�y N�\����([^�q��Cf0h�5J#^�l��K]/z��Ʌ6e��c� ���7�|u�7�T8&\q� ý��	��O�l	�Ms�"�~j@:	�e�`�S�DvX,�Q#y�<�e��S��1��h��>_��{״.������4�?�-O����W֦��)<xf����O�&q
�e���X���ß(�I�Dݖ5�I���ͧX~fMz׏��y��=1hW,�Ы��]�\�h- d�
g��Q�dI�,����M;ʓA�v�1ge�w�x	q6�DZ�b1�!t�]kP�V	S�L�07��0 cZ�k�7ʓ'|��ɽ�M��b��O4h��+ȧJ���C(�?Y���?����?���?�O~���v��u@@�
r���j�o��U��	k��� @�X�͙)R�j��R�2����7Ob4m��'nL�k�l���O\�'- BdBb�A%���
&�_BX��W�	%�?9���?q��F1�#A�� ��Hk� H����+T�ƈ��'B�x7d�;�S5pQ���6D�@��ÏݦyqtaξjJ*����:6����ۻa^и�O���5FxrB�>�?��i3X6�O�ʧs�f��;Z|�tk�9[di����������T��1Ѣ��j�
ݘ��M�3���j����9�@~xh��c���@��si 1 ��U 	kLl��n�O�$�|���8�?���?�vh9�t�fgK3��	��d�n���Ʉ]V�Bcj\�ժ��-��c>�d�5C��\;У�I*�{Q���)0���KA�Rf�8���("&�5��#�m�<6� a�Ed��ao�0�x�I-�M���?1N~:���?���B>��ʕh�5������B%B㌜���?��o�b�"m\#p���'��2���<I�M���A�4�?��#P�lNLܨw)�
4֝9u	U=�?�����P�Gg��?i���?Y��5��O��$�&9�聐Dͱu�������T��F^9R��0����)G�Zt�Ǘ/�E:��&<�$�/��Z-	����^�L�� !��9��/���$MB�i��E$��I��l�'��\i�䅺)���8�BƘ�j%��'��@ѷ=�v��SD�(CXa��.0�S�d�d�0B5��"�"u�틱�8G�!�Zo �� ��9aVn]���G�!���{l�M����7r���G�F�H�!�dں!e*���8t�0�E�Q�5�!�D@�_��4gƊGn��)�̾x1!��u0ԉ�u��4TjPysɌ%!�ěW�����+Ğa0PA��/ ^!� u�V�)�gI2d��ʐeӰEL!��)t�쌈%�o�4F��l?!��3�(�`N�h�x�!D�='!��đP�h�Q�2=�:�DΔM !�$������e#z.t����Tt!�$Ǧ?j�
���o7t�X6C�>�!�6�s�;r5zAC �~!��~�0�����6G|���#�!�dT)M��+��X<D�𕯐�!�FJ	֐7I��`ؐ�m�M�!�d��4�ޕX�-V'l�]I���*>D!�$���zd�e��9	R"Ȩ5���T!�S05�U�D4����Oәp�!��*���H7��$�<�"4oP*:�!��W${��0t-�Q� K���!�d�fs*�sv���bq���/�!�ٳ�l���
B,�j��K,u�!�é\ؾ��b �MaʜQa<f�!��93)��X¡:s��k�b��!��	O�Dd�17cvb�5��,�!�$�';m*�Y��;��y2��7#i!�F.Vb�����P>L�T�po۳o7!�D;Q�����%	:K>ܠaѩv!�d�e���4��+nԾL�/Z�Z!�dI�"���$�!j��;��%��x�G�<�(aS�x@�b�����d��\)��$��O!*��؞a�c?M����tB�"��9)�x��C<?�A��3҄��ӏ.}��i�K���QQ�Z'DNȒ�ѨU���=U��t@�����)�~	$���LD�<���+��I	j��H�H"?��'����#�������}�=*�X���X�(��_9Z�V�jԳT#@?r�>!�ӓ�H5H�h"z/*8W�?2I��;3�\�T�V �I�آ-������d�熖���Qi�j�k9�����!>�h�u�	�&)�\�Ha��s�#��f��=B���#��/hr�1�#��B�l��
L�١B(7�	s:g�W9��7���=P$ ��z��EZ��#�*�x�1�KJ���W��O�1�14�t�a��O	�*���A����\u��#�h ���;���D�(�d��/��e*�/O�<�W@˦A�|��WؼMZPȂ�ޓ<��m �Gɦ���@.��:��f�O@��_�̓d
E�8�)r�^�@�у��&P��U���b��T��������F����(w,�	^8���¤��O��+�d��R�B����L�`�'+�c�t��Q�qrt�0���=2R�Ey��#et��A�1�t�2������ F|"ª��x��CF�L.�=��`�7������,ġ��*�s�S��h�FdI���?C�Pes�	'1�ʈ�uZ���"��8�RNď��Z��h2�������y��O��aa@�S�O[d�sG��%��@Ȑ�-��>H��#R�|�&��z�-3)O`��f�I�"T�EY�W�
+�=���9-&��*FMH�����2��ZV��Q�?7�	7IIb�p�	>	
��4���/0q��,.g ᑤH��s����i��'�ޠR���@�>�p��3X
z-k��I >o ��[.�?�'�,�u� �E,�2��r�u����b�'�qX�J� m3�m#[=����_`��)�+�:��N٩�ʩ��"��V���S�0N���T����Q�U!��F�;Gy�q:�T!�HX�'�a�p"̉P¢��&lL�B���lZ.Tޤx�NQv��(V�N�A��UH��M�6nY�R�I,M��0���L������T�,ݰ֝>ɤ	�-R��$����"dD�EZ�h�@� qcY2XXJ6�@�h��`�E8;d�,K���'[���2��H.� p��S��Mi��s�����Ȁ.@�h�9�@�tԧy�-���H�`��Z*0W\�!��g��{C�\v���'��&Ǳ|b)��4��}�f
�'����>V��C��*�|ডz ��An�aAݼۥ�SSb�mȅ�Ns1v���ȏ��?1'�І|lE��X�����!.v�𐈚�"��A��9XUJ��-��!�	�30��(��K)�BQ�S�Nw��gyb��vCH� ȇ�B����(!��I#`�Bu�*�/ �ѩ��0G�����D�+}(�@'V72�IqG�߬\z$��֏ҫ@�bt!�0O��ȡ_�Е'�Zw�+*@D�r���wa�q�G"v0  @�Q	W+(r.9�P D}�wU��j  ��P9�ۦk{��U%Y����<�Q-9�����KP)�tX� K�z8!EL�F8�D}R�Чw��(���S��e��;�HҀ��M&"�"vfW-ym��[�M�ة�(O��Ӻc�'D��!���;+�(���Ⱥ-e.�aa�
)ǚ0�ϖ�U���5ZҎ4c0��=+�[���y�����IX�N��Fh�q�T�`��&��E�'����u�vX� �ũ^,��J��ѧO8T��EՉ?9*����ע8H����S�^�T�����iz�H��INy���K�-�4p�@XhW�A/+�P���תvQRHc��6�����[@~���Zi�u��/� A;��4/PQ�3��6��	ry2��v�Ͽ����ب�ˬd�ȳ��K�p<�f�
l3��I$�Bo��x`��r����4��u�Z�h@�]��^8��	YyZwa�H͒��c�/�b�� 1Ï�p"~){éʒjڢ���Rd�I�eU�D�%�˅&`��F�%�8����D�)Ϥ�y�j�3-�ZQ��bˏM�ʓ)N��ªm�6�ADi�i�ޭ�S���'3�ზ��37 �����T�j�7K(�l=q�	��Hq���]y�V���)�ht�A�Z�:4�����$��);B�V�\���G��;XNH ��R�yw�L�s����-��i�H��=�?9+O����ι��ՕKRMdM1TV��Z�k��Z�Q�\�@)�$��Aa��e<���E����*g�W�q�@ȯW����O~���Ĩ<� ?>]3�cq��#RJ�}(*"͉�E�
���O4)RPL�32 �#^4�JѥW�,�'D�Ѣc�D.,�6�p#�Q:<�SX���'�:=�W z6N���o�/w��CL�ܩ����JhdY6@S4^k<c��ӽZ(���NQ�%�4��$(�j�p`[�Ag�r�埘<�B ���(G��$pn�7���ˏ�4�Zr��V�OhعD�TN�MQ"Or��񦃵~�ny��C"��T(�(����O���rÛ6_�8��R���{�훦,.bQ��g!8 �F����=7L'`}�	ђ
��Dk��B� Rr��3UQ�a�x����!�˂�"MB�bU�E ��'�v���P�	JN�!�?d��)�{��>�����O8^�MRv*���F��c�	W(��!p�y=�Ad,ف~�`�r�J=BGa{��Y�Ol\ؑF)�l�~�b�3`ʜd��Ε=)���2���q��xZc������S���%�B��0,��di	�'�0�B�'YТܨ%���2���'d@�v��$;lZE��r̨�À�8?<5���7V$�#��5\O��C`�5	yis#V���H��ںv^�Y37b߆{�*L<�bfԞMwf�b?A��Ϥ��]��n��XX��R��>9C�B�7c��"}� )7]~6f �Pcgh�R� ������ �԰=i��Ń?�� �ng ��H�v�\=��G� ���rP�p<�1�ֵH���I��� � B:P!L݄�wLcb�	,3�.�J�ǘ�-���2�f0�9��"�>#ƶ�����=SDސ�Ԥ	#f�B!���b��'�zuz������yG
B�S�p9ᗅ+S�H�bg�!f��%��0p�ޞL��;w�g|��aa�$�Ɉ#�8��R�g�8��"�I�Q���d�,ш0zF���؈uR<���7��B�%8�G�"PLa����,X&��	��8"$
5|OD����?y͠�KZ�rX��ѐF�,n��	�,:>��*�M	~�y'��)�j�Zq〱W�����C��yb.
�kK^}bV���vI�šŷbf�E}��&��F�V��~pj�����X2��L�֩!�ҲL���'3|O*,�`����2�Z6�-� �A�Ě�R��A �m���A���c�, @[ @��ԛch�Y�Q�<,O���ূY���*�Ճ*Q�Ȱ<*O*P�� L�*��A��P<�%�>�էW']Ȥ��-lu��!���8�zt@Ս\l^�P�'b�Izy�?-�tG���Is�'�*��t��!�"�tݲ䢎W�b	���]�Z�Q���YT^����� �Z��⮗V ���<i-Oƣze�����Sj�� 5��C�-�4��F~BȎ�K\�E�-�Ф�]�[���B1F0b�H��+��h�.	�	Tc��'B���:a:B	��䂠>���Lpj����I7-GF}BH_�ɳ.ڎ��&��~5X�K�
^�������$�'�|�Fe
�`��H�����]��˓iD����6vvT���YE�P��y��'�$pT�C7W�`IR藗ې�vB�!%8uq��d~�ɱ��ĵ<��~��`�2�.ıV䁖	�rx���Z��0+��R<+�i�d'Ǡ�p<�1d�`��L��x�h���<�!@Vy�Z��#D���H���Cׂ[��yh iˠZ9�m�4O����S#���Uf�5&$`��%�ȫEa��R��*~�viTi���?Y���d�<�;�y��O�ZU�a��c/�2��+L~�·&1g���d�4?��g�9��)�!��	!�f��g��o?��<!S#ٟF���@B�N4g�zA��A�
���~����U�j%�נ���$L��36�x�Qv+��F�h�b�"	�9a���:%7�Xj����Ԣ�P�ė'���O)f!���X�� ��ع���Öj2}q.�Q'J!z����GYԧyG��>|A8Ł�S'"T��1��n���+O�˓.���}��3;�8�B˨EP��$b�_v�<��ɞk����S�*�6 �a��8!�� �d�̡b�#W�	��Zr��O"�Ĭ<I(O" I"2Ort�T#�eW�!��(�r��z�M�]	�y�0,[ ��X;E�iH&n6 u��I������d��s���G�J� '~�b1�D8lhzʓj���1�Հa���e�Lx�𐧟�ɛk����'�6�X��1���b������:�=c��~��?aI|�1Q~�&�оF:�����([`��(B
�i��P\���0�Ӽ#IڢG�f8��k����m��MZM�ҟl'�8���I�1a"5��ӉdWfP��@M\D2��I�|�<�Jrm.���A,c�YB�*�"�EA$���Tk	V3�'"Rቒ`j-#�b�+����Wp�.��%f��56���L3?QC�<E�$m��ǉ����n�c��:�%ɝ,ĝ���G;�BB�B�h�'�X�q$[�{�X�9����6�
��OƑ)[fj�p7˝�}�5����Icȕ//�p�����^��OT���,�xF,8)4�K>�QP�O��,OBL�c̒���Q�E%��O���hb�dZäQ�<Z����-]�>��'�ў�>�Ra��N!��(SCĚX��a���	U&����!ԳS�j�Z���qlp�������Ǒ& �W��D���>�&!����"�LN�G�P�#�@K�}%�HI��K4}3r�CA/�>)�NZ2Gߢ處�*:�ʐk�-�^��?u)�q��y�*@(#��� !a��n�O$�\w�+̀"|�Z
al�\��	�h��5"��O.�Q��*ټX����bGJo���J|
�/�1�yb�!P�8s@B�hܰ�5lޡk�~-�G�����1C��b����&Fr�y֎ƙ+2@�%/���	�s�$e��`��A"��)��_�p����э�,����EO=��1 7��?������U<,����U.��"��]ɵ�[�?���ʡ ]/-��ݗXc�dF.Eiz�)��6�0�3�2^���I7v�8�8p��9��$�/xκ�q�	ס3�̐�,Y/�O�ħ�N���%��]�0:c煿O�
��4,i����W~>֝#\�����-����18g_��
õ��33� iF�l�T V( 0]	�#�s�O��O�L�� w��ro01��
3օ_�N�+����iwG��p3`\��ℙ2:
#>�;D���E!X�B�^T���(_����'�
���H~Bc�8A��"� ͣS`�h5'�@��"?	�9D�� �L0?�'-�:���Q֬¡Z�0S�&�8�hO��Oj�)q��3,�H��(�㘱�>Ѡ�c~2f�#��|�E'�Q�ᓍ\������^]�"o�$��	1X�����5or�S�O�^�R!��>�B�Y��%<��]@��%��||�\B��L>9�hQ<&q
�SB�U�羹¦�v���F��|q'�=,O��ҕ�M@�Ƅy��P�x�墂"O���C-gp\�#��ب#�,��"O�2�� C�N��#�P)
�X9p�"O���v�FrG��qe��qY!"O��2E���
H���!S�(���"OBeą�P�H��#ڛ.w&�:�"O�Xi5 C,~�`���M<TX����"O����]�gÎ��G�%!=�A5"O��I�^^b�i�D,ZdCa"O��;4F���>���e�!����"O�ݪ�Mթ�`�S凿_p��	U"O� �]i0ǆ;M�.)��@�v��ID"O���F�wR��X����S<	�p"Ov�#�l�pՂ)1#²i-� x�"Oj��Q�����a�n�N�Yd"O~�)�.ʟ[��}����CA����"O:�sP*��	�������%s(�|BB"O�$�1�.U�����~{A��"O��@���U�Ha�M�j{�Y�"O<�wK�-M0%a'(�\e��"O�-Aa@�:���ReF�a_���w"O�Y�d瑅8���aq�R�|N�]b&"O<�rd.��.�%�[�H�t��"O}cMPOa�!"#�
Tn��&"O�h����\�����-�6c@N@�&"O��	Rʉ=%��H��l�d�(���"OҸ�&٦[3h��`�~�y�"O�d
�텗*�X��mB9qب��"OX9S֭ q����g�ܽQ���F"ORE��ǻJ�+6��_=ν�"O��y&!�,js^��c��+Q8|��"O-����Z���ߎA04͡�"O+��H���a\W�x!� E�<�$T-L�&�����(#^���K�<��+�&l�x�J�n��H�a!u��I�<��G�3e�}ҲIK��rb�W~�<�TlA�l����9��q�@�[v�<A���<A��٤J�<I3�(�qo�r�<Y�ʓ�qsTu��@:
 䍌T�<�Wf�.Qj�P�mѸV~u���z�<9'��f(0���4b���2��~�<��e8s�r���g�0|�)�WO|�<��_eq��ے-�)L ��ՏO}�<��4x���5Ǎ�W��p� #�~�<�&b��h����BA�WgFPW@b�<!�LF'.��[fL¹m%��K7w�<�t��&2tP��a�2V����7T��h���7�i��Ƃ�pҠ�0�n0D�hs�dY'��n��V|���m.D�����R�||P���(ۧ6".ሇh.D����䄉��`g�X������M?D�Ĳ@ȝ�]!z�`�ճl���W&>D��iT�^�fY�`+��5.	*=Ӥ�<D��(r	]�v�A��X�MG"����:D�Hk䓶'�,�BĈ�+g�����&D���Iӂ=<ɲ���
u�=���#D�P&bY�^�����097�`rg�%D��	R&U�#d��A�T�P�Tx'�"D�ܓ�!��)��m�Q�Ro�2�3��!D��P!��6e�E8wIрU�D"Ə!D�p�����b#���k��at� D���W`�d8��s���	�ĵ�"%=D���O͕E^�u��X�E��9D��7��l=P���K/`k��C�8D�|�n3&�z��ƣP�j��b�4D� j��?#�:��P�E?/�mɠ�4D��r&�?,�b)�1
-'�L�	׫2D�����/1�%H��]$lcQf/D�I�fV$I����)C -9����/.D�����R]����1�ʕ��-D��(�!R-}����RN�7~O��qw"?D�0q��<$�h�e�ܴ���f�;D��GJ�w�kץ�
5O�$�!I8D���E� BVy��ſf�t|�Q**D�z���'=��z�ɂ��l�#�,&D�� Ҹ�$$C�Y�ʭ�oG�W�) �"OR}ӗ��nW6�QU	��3�L�r"O�$����.Vd����*��C�T�
B�'�l���T: l4�H�s��Ҧ"D�l���'V�6��ǃ��m�J�0!�;D��bԀQ�S�,@I��[[4L�l7D�p��ՂoA�aB���.�L�Zte;D����X��xpacB��� �@9D�x w���� �H�v�0��N6D��!I�3�q��K�/��1�'�3D�<`�������I�7�Y���5D�����C�$aQ��g��J�a9D�PㄚG&�C��
x�\�t�,D����O�dT��� ��XxYCQD=D���#�ĳ`|��voܞ�"!qR�:D��K;N�ꑻ��Yf��B�9D� ����;b X1j@�A�=c QX��+D��+T�M5"1�a��E�|iؐشm>D��a��](��(D���Iоi�>D����;��{儂m3��`�(D���#		�;�@�e��W3��R��'D�\c0kwh�
���H�z�0�#D��`��P�w���@�5�Ȃ�"D�0£I�o�$�!fZ�5�<�
�;D�̃&��Et���5J���B:D��p��Y :,�ԃ�2\��(�4l8�Ic��ħ��\�� 7H���d��!��=�ȓo5�Jb�40v`+�G�z�TH�ȓZ<�\��,�>2��qSg�s��݇����G(P�j�n�IR�؁Y*}��]��B�d�D��ǉ	 �0��ȓ�船�&S��l8ʠQ�}�@��ȓ؀+qjD�N��(21	�h��	�ȓ�vp����
B�&e�"�;1[�y�ȓ%�V8���%C�0be&N�~�*8�ȓY5�h�e,�$Xa��I��,1x��g�� �d��i �|��%ֲ*f�d��Ah�D�܉]�d�c'HdU�ȓ0�,
Ad��F���k�� �>@��l���
1���P E,�;��X�ȓe쉰��@p�
���L�+f��p�D��#OD-TJO�Rs�}��/���~w�ԓso��GP�����Rf8�5)�i�&�j���1��i
f�P�b��,IƊƦ%�I��-#�޴��T��ؐ�H!��Y�n\�t��;eJ)Ң��V���E�Ԑ���7!�o�0�d��&�4�{���� )ZYs�A�&:���~c�!KD(e����H�+p�pI�ȓ.$v�C�'K)f0mcE-@�m45���n��0I���y5���y���)����qDZ�P��4h����%��-#��=�P���Hڕ
� `�ȓLF�Ы��ԟP�6��!VJ���ȓm0��RO؝mL����$R;�Vu�ȓ*��Z�eĥA�
��a�i��[!���ѥ�I|8���IPf��ȓ` ��!�xf�w��q �D�ȓH�,`J��O1]����D݋g(�E��p�j�rWNՂpF8ܢ�0-W��ȓz��`� NX�hƈ�kӪH&1Ňȓ7�䈩⣔%+�,�ۄ��+2ξ0��]��l��juz�3��0�T=��S�? (,��T'-������q ��R"OVA#c���50����kA�2�J<�"O�1%N���$Բj��ֆ"t"O�#�i	̠u�(�����G"O�ՋgL8s�B�r��F�LM�v"O�1���0L|XI/�U։8�"O�I��:������kL��٦�Gx���'w���H��1&l�!���"$����'�\1����G�*�����,��a�'�,q������i����ƼY�'��I���#RP��bI�.�ƅ��'����Ϛ"=�=��h�,�AI�'w����d�#�����Ɏ�L0�	�'���Sį1�&�#e�ŝ�H��'�*�;�C,>��m!u�׈0Xl `�'A�IyEDK�$,�<�ԎP')��$x�O��=E��1e$h���	5��!���y�f�i>�0��
?�B�oߺ�y�C\a34 ,��;��F�y�M�<���[w*R�`h����.
,��'�zRL%j�[wdJHWT)��-Y�y�׬y�Aǋ�/XHp�rd��y�Pv��3CP�s�R'L��yB�Y�+X�8�Ȃ�f����ꀱ�y¯'���ÀWͰ���H��p<���2ozzt�P���T� pKJ�mA!��U�z�Pkɓ-�h��e�M�F^!��"u�Ҝà��.f`�����|m!��H��J�u�ز5}>̐���N!�$C�	F��r� Zpr��ITK�A�!��2DJ�ahC-\�Le��ǋ�t
!��qv�!����X�~�"`E��	(!�$�|��AX��@���򱤝�r�!�J�A�Tq[��}��t�5E��!�$Ɵ]n��a�Yl̪�{fď3�!�dÔf����hH�kR��� űR�!�D���$X0��%��,�C-��O&��R�x���h����d��ث�"O�9z�f_�\-ѴB_3~�\C0��d����/�޴@��E��`k�)M�}c�C�IWҢ�!���>�H%��ʚ0Y ��hOQ>��DqQÎQy,���#.D�����(QۗbӅ}�Th2G9D�,s���t�4�6�O�\��H�:D���ھ@���bp,�F�Uy�
:D�$!�Z�,X�qGg��\!��#"D�܉����2ϪT�s+�&W⠳&J+D���􀌞!^�$qQ���T����UA*D��Y3Że4�Za8p�hK�,3D�P��‭.H�lJd'�+��P;�D/D�xj1�S3"��%sG̹P�d,;`�-D�P�!�?eT��%��&u?�x�V",D�|c�˛�.�����t �bW�(D�D���ۚh�~��3�G�)J�4I�#D� A��9n�V	K�k۫l�H���?D��
��.�����F�f�
�"D�X�uA+6:��ʕ�l�p���,?D����)�ڬhuÑ�8�9[��<D�tq�fǾ;^�H�*��b����;D�x9��J��8�ԾM�TY�q�,D�؂U��2sF��gM�_"V	B�&D��0` �\2��kR2{�liec.D��s���^��:��0�T,D�� �]�J�,����	�4�l�.^U!�� v�p2,P�w~���P�K�
|[�"O��Q��,��!�V�.EX"OnhE끎t��*��^����"OjXбbT>ȡRg�R� ϴ��e"OB�9���U� d��N�5�l�4"Oܔ��ͪD�u�.�.d�ڠ��"OH�	�	PY+i�TGM��"OZ�0pm��Oa��T���_F�i:E"O� �K�l�w�D�G/�D�"Ol��C�H��bXyE�9-E|r&"O���%[KI�I@���(*0��x�"O�̠@ꖐBÎm�f�v#��� "O@��+�`�Y�g"y+��Q�"Ox�T)M�;E���TFAj���"O*���! ���Q>h6�a�"O���Tg�-���R�c�n�{�"OT�0d�1�tb��>ASj�""O*��(�hC�0"�e�'G�8@�"OМ!N����isf��0=�`{�"O��O /���S�m�<6u��"O(� ׇF�0�fDY���jh씩�"O���`ȏ+�Z�R!��AB��4"O��CH&K�B���)
<�TL�"OJ��/Z;Hrf	S�Z��"O��tN�9KM �R����`!�8b�"O>!:c�3z����61�0R�"O~d`�XR����K"U�\�4"O�]�FLSI�*x��HӦLF�$��"O �׋��1g�ȫ�ɀ�8�xm�w"O�Xb�EZ��HB�Y>�EXv"O��1U�CTu�-�5��90����R"O@IkG�J�4��#���_�l�Y3"O�$p�H�)*���v��I�5�E"O��X��ΛNf꭪s�ѝw�(`�T"O��#�✠w*��tg]*Zl�q�"Ov�C�S1F�X��D
=f�ṕ�"O�(��HX�'�bh���6c�,u�"OP�#@L&�}��l�[��l��"O<5�d�v��$��Df���"O��Ѐ�\�Kf�-a���䃒"O���2�$&	^�ч��\�^��d"OD��1	�s洱���{���0"O�dZg�&=s�@2*\1�~Ѳ"Oz��Y?`�z���H��~��X��"O<��'���p9���^�d��"O�V�=+��x'�B�W`��"O(�j�f@��,Iɰ�I$�T�`"O����l�<=F���E�'�9bp"O�����Z	j�Mq�U�m��"O`�th���
:G���E�ґ�"O��#Iۚ+�Pw揭�h��c"O���ؼ5�@(ǳ)����"O"�0��0rD�������3��a�"O��!q'K�l� qƂ�d�6���"O��b��+B�L���E�+3����"O��h���&�i�(%�t"O��1��&���桘3I�BE�"O`� R�� OLby�@a�g�x4�E"O\���3��W�ܐx�d	��"Oܤ��fC9H׀}@�dL��T�)$"O�� /�r�"\I�B�9'�ɐW"O�l�4N��I��#a���ԛ�"O���֌J&5�	J#�V�g�
�g"O�R���XhR���W�J�
Y;u"O� �tr��O�7=�-H�ʶ1o�D7"OB�!! 9��zG�u6��"O��:�U�,? �+T�Ny��["O �s��L��"�3�bP�a��$AT"Oj,
`!.J>@d�F�� _ĺ��"O�-����W��%��hȯ8�}9r"OBhQ1� U	<�0	ߙl<��v"Ox�`��H�P������w�0!�"O���6hOHdI�+2�����"O��P@ ȏT�X�'>�<P��"O Tqe/�)%�N��a&�~9�&"O�eɒ�rq`�%
HM�c�"O�p���Q{oN0W$��"O�EYT��@�()�6Ç?C6�;V"OP�:�C]#B�3լ�p�iku"O�x	�C����="ŉ�0f�Z��S"O0�D�]�|p֌z���f�>�	�"O��G�1����K�zY��"O����c�*h�4)�&�;
�P�ك"O\pS¯���zYX�%�&jr�Ie"O4⧈�+%�R]y/�-Q�x�J�"OLA(���F�=p��L{���"O��_�kwDͰ��5Bx:T��"O�Ya��NBH!��'�I�"O���s�\�0�<AD�K$&���"O�t���O�Ą�b�d�!�"OʉXqHP"qV���%�2Ȧ�;�"O���AM{$=YV T���9��"OΠQ ��$w��ʢ�7yL���"O\S���1G���8k�5�8�c$"OF\���S�B���D
�C���J0"O�QI6"�$Q^h�'�)
����"O�з�T ���@��>0���"O�ءC��8&���sb/��E�Ě�"O*��W

�S �Sn�[ٴ�v"O��p��[7Dk���R$<���"OL	��@�8���PL�2Q05��"O�0��֠J�jh9��y����"O�¥�X,_� �bE&K�sw"O�@3,ڃA�J��g���:B"O&��d�4PYDp�� �#+&	qq"OlTŁ�j�\8St한e���2"ONu�B���\� �W�&�2�"O�4h�	�9��l��왚5u���F"O�[�(G��R4奇�u[��h"OH��ƖLOLリK=T�j"O$�w��3M��J@�Z6,\��"O��i@�@�xeC&�\,L}y�"O�%��?3�VL��()��"O> �"��R��+���z�"OB�a���Q,����_�J䉛2"O\I�L�5� !�Ф׏a���"Oh���nO�x��Ŭ'��a�"O��J��X𱗋D������"O�@�eG��d��$ɕ\��]��"OXqH����LcBI#�(�p�"O�0r2$��Lw��u��;�"O~��P�?H-rጪ1��S�"O*,G��+-�)�Wɢ\M��B�"O�����O��Ap#�$7BD��T"O���f&;1l���hyG��K�<yr��~������_q �����G�<Iǃ�3�vE2!�^L7f c�E�[�<���7�=���J f���|�<� .ݛ�HB�R\8}��`ͤZ�n�8�"Ov$�ʏ�7� ���E�e���"O��������X4k��:�"O>E�U<O�� ��`_�Z����"OR+D���0z��X4��:S�Zc�"O<h{�c�b�ͳ��B�Ec��ja"O�(V�9l�M��,L�dGH�@Q"O0Gɍ"^��y�B�șN�\:�"OD��A�
�2I���	�� i�"O@����"�81�@�8/����"O0�$K�,K�.8���Q)o�"�s�"OLh��j�,7Wz�p�/�n�&Ń3"O6Lx�B_ =��eyQ)\����ʑ"O��
���7w �	��T@3���7"O�B'�,}|���-�I/� �"O�T���,Ob&� 􊂇j"	Y"O؅ �`Y0w�m��Hk_���F"O��kD��a�
�Z�a7�Q��y��n�`s+��KF��y���y�(@��v��<%+@��p��)gLA�5��9E�n}YF
IYܹ�ȓ;�����܇sߚȃ�ߟh� l��@�$h�w矰I�~]#�*R�\�̈́ȓ$p�)k�&E~��A/�1u�^4�����f��n�˕!öU͞h�ȓ?�b�*2!�!A�n���ȓL��i��2b�L�8wd�2 c2=�ȓ��<x�ˍ�="�:+g��ȓ|����Q4I��`Tj��Zy��ur�0"S�-����6�V�K�ȓ�9(��8@�0���JWjh��-O��#! #� p�ꓨ-�Z���~+��Pv�Dd0��/�"3�����3�]
}!�]�W	W34ê��ȓC΍���@G୙�g�, �JІȓ0�1ck�������V!K�V�ȓ
��qa��F�n��Y�U��$CiX0�����r��ߙ�.��`U�?`9��D�n<##GVo����sa$4q�`��<@l�璼
��ɕ
S�O����ȓa���H�V�I.�9!*P�C�z�ȓ	b|��CE���\A�#R��-��r�t�«�
>������R56�������v�	O����*�@��ȓRA�m9ÁȀ(bD
��;��E�ȓZ/���f?l����UE��^�ȓ+`pY�!����L
T���ȓ;�<!SD;n�
DX�.�H��6IzE�BJx��O�
W/R�ȓZ&��"�"����0���ȓvgT�kP͜���up��MFP�ȓ�<�y@	�9���R70�f5�ȓ�t�r����M�N!���74�D-��d.ͫ'܎-�4�E���Q�ȓ1�J=�E��	p��殄"\0��ȓ|H���E�<���Q8t# ��jXj�B��,��a��1d���7p&,Po�$#h���n6=nلȓz'D�ZW~A��/(�ȓKF�i���׶#������[jNU��462��ѣ�f��Șc�S+k2
9�ȓ?����D m^���	*G���ȓ6)�Ճ��û w"Y���J$Vi譅ȓUF�@�� �zm�[fJ�@ְ���S�? (\�4�R�P�hP,�$=^p�p�"O�Tb���l��E�!�U8x@B�"OTx{j&D�&X���j)d��F"O�1YeL�D4��p��A12&��"�"Od�U�
&P�)c�^�m%z��"O���֢)�:��(��F���"O4���o�-�}�����!$"O,�s���wY��;�'�e	��S�"O|�҇J��3���;�`�XK�A�Q"O�� �⎙#��, �	K^���B"O�ɹ��/)���YW���.�=��"O�\�������@�I�<*�ƍ�"O^|2I�0PƜͣ���v���"O2Y�B��=�.�j�
�	2�^�q�"OܠY5_��|�X@���?��T �"O���& �4A�]Y@*�g�a��"O�ͫͦ>*$(+a��d�"}�"O�!Q���76 �"ׂM�
��@�"O�I��)t�����號m�&�h�"O�Xz1NT�b��G5y~�A��"O|�� �|�`�ʗ�ۓ6?�Y"Oz5��,�lcf���9VZ���"O���FgǄ#D���S"���"Oei D�!�6M�"�S� �N��t"Op��CJ]���ta��T��s"OF�4�Yz�~�����9^zT`��"O�}PP���M�4)qc�I
��H�F"O��j��D�m;���Ā�sq �Х"O0�b��S:T
�����jJr�!�"Ov|"s�ݰJs��8���/gF��
P"O�$���=k=ȼQG�� ́t"O��0d��F�!x�>S(� �4"O��s�=%�*��g�˴(ԝۣ"O��{���7,�	aR�����l��"O�L �Ǽcb@DABAS?b�DWf�<���Ű;f|r�C̾�X��G�e�<f�S/�*����N�d�	b�<9����@�$�� �@�}g�1 ��[�<�!�Ɖx�޽�ǌ5;���CC�GV�<��#�Dt��J&@0R�@�GR�<�Ѯ�*+���Y��F�<=�&��h�<�c"�L{t	����(��| ���J�<����;�2hp2!Ʉ�iC$S|�<YFFQ��A�c�%l`hؑ6�z�<QEc�[�`��򄐟1)[Ɋt�<�C	�I�:Ix��/�L�bb�r�<ya�W�,G(,R"�T��rt	y�<��
8*t���WDSX�@TK�<�p�;:�� 	A'U`�4|11gE�<�`oɾ!>�	��D֪>4�rU�A�<��ùW��02%%���f�:�&�B�<���R@�F��u�K�N��Hѭ�~�<!�&l\Ha�O�5ib�@�Ђ�|�<I"�K��i���1'�f���Zw�<!��d=���Dʯ1V�\��	y�<�Bj%0tNE�נ�nU��h%kCx�<�ЯOB�bᰴ &
����3�@�<�f�J�GE^ �V+D��~<��FMx�<is+i'$�q�)M�11B�;WnQs�<A�c2b��hj�M��ҥS��p�<a$��<hr°1��<p4KR�h�<�Į2I��!V��1l�����\�<�d��;
t�i$h�")\�BM�U�<Q&
F�Bx�P��N�!c�\T�<� Ԥ
��bl�0�'Π]��� �"O`0[��<`s�q�$Q�b��$"O�`H��:[8��"B-�2�&"O��@cL?�$���"�˦�a�"O��2�%�&��T��-"�xa"OX��^�i��1��A�:�%ca"O�e�J�
��K �k����b"OL�#�E�F�p`�X���"OR�ѥ		b��� d@�V���"OZC�4<�L�ABp�HI`"O5�B�Ĩo7�� ���L*�y�"O<�!Q��F�2��&)"����"O��'�ԕ ��]��
�G	�-�w"O�h�ao-�I�u�ѣR�"XA"OQ��D��m��A�'��:�� ��"O ��E/�?r}�e����x�\�*�"O<	A#G'r>Tp���M<h�M8�"O4P�AdP�|RFa� �4e �V"O�8s��"[��X �p��!"O�ա�,~�.8Jd @.~��t�b"OV��Gc^��$�E@�vv҅��"O0�"�%	�q�tLJ4��$�9�"O�8����ve��1
о9 @9�"O��(��	~�!EI�PS�yT"O|! '	���v��|-�P�"O�q0'��u���*E���q���@"O:$g��!8�~���kP�L�*���"O���h� 	��Z�늯u�u��"OԱ��Eq�pPP�[*�h k�NLb�<Atf�0N��cʒ�{��t#��X�<yb��Np�C"�[�U	���-�{�<�cK��<�7(ݩ:y6bF�\�<) ��/v���c���R�&�Z�<��Ҙ"�`@t�W?ь�A5+�T�<�QK�9p���'�u!�4Q IM�<q0#D>N����D�5�`S�RD�<	�!سs� ��*2v�RXX�h�C�<�u�҅|0X��eOZ0-|4��IYV�<��B)7��|Q�ɀ�q�]�U,�R�<1�P	llf�0���;Y>�tp�%T��#��脸y�
�/R�@"�&D����ҿv�Z&��bm���#D�ʤG_�!�~\�F�'z��8��&D�X�)
6S�����,Ɨ &����G"D�����= ��]iP�3�f�0�b D�ȩ�"K�Z�`���hJ�:� $pG�?D��+�H@<���r�+:!d��P�0D��3 ��l0�����|XR0��0D���Uj�1���)���v1L���,D��a.ˇDi���#Br]V��C()D�#�C?�Ԕ��Z=���'D��b�c��+	41#��aexGA%D�P��#�?�֡��O��9�p8!T�"D�,3��*]ɰ�cV%�h���#D��pBԝ.N�y3�_;-b�9�.D��8�� �\U�$����08"��-D��H�̓��t���lF%?��999D��ؒe�  �FC�2ۘA�)D���v�\Z�4�"�;m1\9Z�j$D�lk��
��D ���	2�V��s�#D��3&��&}:�"�� �"Ѱ֩4D�THU��P�jŢ3���)����3D�<��J�:Y� �Pg��$q�$D�P���UY���z��K����"$D�� \�he@��y�b��&�9}�ṁ"O��(#C_r���q2#�8�ke"O��8H�/dw|�7<ɸ<�q"O�Ax*�HҜ��H�5����u"O �P� #c�����ƕ�	�`��"O`i�� >;U��J�E׀^�
� "O��rA�
1<FX2����O�^�b"O�����j5��倾�f��"O�Ӆ�� !�B-R�NF�"O� ��E� ]�]��	�3"O*E�C'E�&�8u���4mX�C"O��r�	b bh ���ϒ��"O����`�a���#CG(��-�"O��s��:#�N�{�'��>�V��S"OtI3��S;)d�49��]-Ey�5��"OR-Pd(�P��"��vę{�"Ob@*�`�xG˛�[Di(�"O��",̂��c�c
(���"O��c�a��Z9R��V@��D]��!�"O@��UW�=��DQ7��/Z�ٙ"O�ȂEm9(GRl��79���"O`�3�VS��4,މrev=!�"O�)�� � %�i�a��:O~}�"Oԙ��ꅊdl��D�!?�L�6"O��*#� eX(q5��_�LLiR"O�\��D�!��P���H�<)vQ�"O�,1wJ_�(��`ku)]�0)b�	D"OX�C��Y�`��	L�h���"O%XG`��v�r��AĞ9N��8Q"O����E��p��
o��j�"O,��!��tl�\y%��"H~��1�"O� �4EF�	������{c�4"O�9 u��B\j�+^�7Th���"O�l+���i�,)rd�dt,��"Ou)wL�y&2PI�C3q`J�A�"O$�p���$�Z�у�˿BP��9#"O���J$0 ��k� 7H�
w"O��k⠌�X2��W$�8c8�](U"O4y�U)�3l}` �鐵7��@A"O��S�&��Zfə���7%�3"O��\ObР"�N��L�y"O��/%�@@w�74��,x�"O$�+�m��&�.S��n��qZ�"O����	����3�O�o��""OH]aB�R'x$8a7�ɉ
!�E"OH��EB]0jw�+��.?��9S"O�U

ĚA�*%�D�V	-��	P"OƜ	2&X�Ar"�S�	9 �%��"Of�zdP(}.^J6�F�(s���"OJ����A��D:	F�X2u"O�]@ �^���Rꍱd1v�1 "O*m���K}M$AjfjP�!�U��"O8 �,��#��8����X�`��"O����18-zX"w�`�"OxI�SA@�<\:D8��(W��q�"O�-���%����N 
��`��"OT<�����&my!/�xDIg"O(@��V6Q�J�͈�^^��J�"O��m!O�N�Xaq�L��Z�b�2v"O��4*�2O�ؕ����c���ѷ"O�P���� g���c��k)h���"O�\��� 	���Н��h"O��۲E��q�A±G����`�"O:��2�6SX�,y2���(Q�P"O� >���Z9����h֋y뎜��"O��p�$U�=:���ю5"Oܔ�#�0d���㷀Q!V��P��"O8}���ST�]��@�S�.p� "OT��M����:��.��W"O�S4�V^L�Ɂԡ�$C���"O�h��Kר�^Ej����U�bŃ3"O�m�eF�������h9p"Or� 2nL5t�u��{�A{"O|�L�4���Ѡ!^��N�;E"O����e�^�d�k2�%f�A�"O��AMO))��RhP=�<]f"O\�hT�8q�5��&66�6 �"O�8;��ɻ7�p�ˀ&� V�ԉQ"O�yR"՚V9
H�!F�9�D�1"OD��c���x���R6��~2���e"O��X3��{���%��o�<�+W"Opd�qc�4}�x͙e��H�4 `"O0T�C
�"�0�ku��:���q"OT�	r���u���"#��n���"O��ң�+pf�aLJ�0wr��"O�x[0
^,)�=`Dȱ{AtIj�"O��*�	�HΚ��rA�f.��"O>)�s�� �j8��a[�F)��i"O�}{$%���jQsN
�?x��"O�Sk���z�[x,����"O,�:��ͯ�	�Ѕ�Q*����"O蕨B�o��Cf%�L ����"O&��ĕ��nt'e<�,�hR"O�I(��2j��K���	t"OZ��V�\<Q(ڠ��΄7�&�"O���Q�\�R[�AJ�A�:7�Aр"O�:��mBx���6�-�&"OP˂I�+���nT1,i"	r"O��4��l�.����uT��0"O����O�g���Ȥ��auD�zt"O �sMѥ<��P�aF�#����A"O��8g�I6�$���=m���K�"OJY*w�\�U �9�F�+��0"O<5�D͂l�JhifCߧg���� "O��b2C�rM�m�硗���l	�"O�c�)�xm��1]c`%��"O�Щ@�W�
ܤm�EhϾe0N!2"Orp)��
Y#�i��d�oD͓�"O�`�U�,P�G�ef�k��2D�k6�91����AǸ>BX���/D�D)���+i�����C�'>���
�-D�,��ЀM�9v�B�+����SN+D����?E<��l�,�Đ1�y҄٭XΉJ�G�9�������y�@�Z���)��b򩚑l��yR����	����QM�#V81!
�'�����@�fk��$(G�hyr

�'v�م���^,�H�L@ c(>X�	�'3Xy���?=�Δ�bΊ'?���'M��7GD�YJ�h�a�S!�q{�'S�r ��6V(��t#1G��Y �'���q@N_VND��!d�#@�e�'{�!�@f�h�֜���J@�����'����G<n!���Ł7�NE2�'Ap9pC��X�~I;�	��*L����'缸�JuuB��&l���H�'a�5�3"_"2���Wd��T���'G�	�=
]����c�O����	��� ��h"%�2^r����n� a�-�"O�Żte؏ў@rЌ&C�!�s"O����G=~��@� ��A@pA"OZ)q@+��}��(�@�k]�%�f"O��(��ɽ5V0(�S	U�*X|"�"O�e��	ʐ#�p�1�@�;4�"O���Kw�t1 ��đZ5S�"ORu�T�ą"��h�%�H��,��"O�y A��U6�VzGZ}
�i���y��,zx=cW���p���[��J�yB��1Q!��R���b���Ҷ�W��yB���K����ScηaY�8�f��yB�G�Fd�H��9[_�MP/�1�y�MŶKEV���RTQ�q���ՙ�y�-ŶpYb9y'e[
G|�QU�K�yb�P9RT�ИT$]%F\:��F@��yR�1[�P�'�83�x͙dhK �y�̀5�6TIg�׀&�^]j'�ƣ�yR�������u�(��ǜ�y�٘_t8�P��L�� �m@��yrϑ�J�� ���̤I&��X��y��N�Tm��U�6����Õ�yЇ%c� �k��+/L�{�n���yҪ���rcF$D�u�����y��98��r���o���G@�"�yr*�!W�ti��Ծ�AF���yM���Rv��/(Z)J�U��yB���C$��0�؄krI������y2�����b�g�U��1t�B��y2N$ ~��j��ӓ	}*�	d�W/�ya�#JpLԉ`^�}+��s���y���?qS� �ʀ�ha���s�]/�y�'x*0�D�G�g-����Ã��y��z�pa�I�"]�P�fĄ�y%j>�=S�C	�T�`�L^��yBW�'pb̲�T�����:�y��܊Q��(���4;�&�i7�G�yB�
�
�xIwJ��\��q U��y"��&<��͂Wlv$���� �y��H09Rb���]Ԋ1RE'���y��3H�`�c�ӃX�� ��KM��y�+�
�J�%JU�����V�yB��/�`����K�diT0��E�y�F�09��S�BZ-�	Q�G9�yb�4����Q�޻Z,zh)�d	/�yBi�|�:��$�GM-��Y��&�y���g���bg���H��e���y2��>��AS`�#��Y�r��yWS��!�����t���1�y"��2y��p�	~���H��y�`D�@/���e`��~c����y�,�"am�(���h����C
�y2#���8`��ڄ8X܁q͒��y"J��{���'�nT�䛰���y���wf��A�$G�`´)p@����y����=G8���7Q8�� �˕�y�(�떴� ������RȎ��y��F'
Yۢ&Z(kz-����=�yB��F?l�8Q�ٞK��-(b��y�ꃳ��@$\(A<h���B��y��-z�ؚ��M�>��Y����y�銜R�@��$Z>�`hr�l�.�yb�̞��h�$I@�<�(�����y�h�0┙�7n��4�Ш�0B��y
� rň���X���*E�m��f"Of����	od�����;�b�ؤ"Oڕz4g�"V.W:j�&��S"O��(�jI�	�����.��v)��"O2��ħ�?dLt���xSG"O^tB�A��H܁'B!C�BTP�"O�����.5�j A���0����"O�0ƨ��cS>�X�l��;�Je�#"Oj�@�O��o��� ce�+�8���"O����N*8��
*�7�Hq�6"O��c�#T?<��([{�,�i�"OP��dΡ/4�9� ��=m8TY�"OL,R���=R�\96�^�Dx�C�"O��7'�fu����2K��`s�"OD���A
*Ԑ$��通@�0&"O0HY�AӨ�r����ِm�z�"O���ެd�"y���L��Dc�"O,$��"��~���ѷp�©0�"O�A���z�eá�#C��
�"ODU�l���0ga�02I�0��"OȬY��
.�R%Bs)��}U�q"O����62�0��!D6IY0��"O��ѧM�6f��ል}^ �"OT���a�F�LaH�㓑|K�	(d"Oz8X�e�:d�.ps5(ĩ#J�-�"O�4��P�)�ޅC�B>Z�R"O>����z���p�֍X�4��"O�,����S~�Y���E���`"O����L���ʢ�2z��"O�h�>n|r���Z�~E�"O=�����*F�l�J4�)c�"Oz4W�	<a�~R6�

H��&"O0�Sk"3G
IfK�%MJ�;�"O`�Ps�ڸ|Z=hшb�yAC"O(���ȁ!�H)�˨�|��"Oj� ��+n�j�F��U��w"O$�!��8/�`t��2�ZBa"OD����VsPJWo�ޚq(�"O��0C�0�v�0pܶ|�@\(�"O�ݹ&���*Sr��G��U�8�ҵ"O4��$�V�ڌrUDޥNԎ|1"O0X���ūO��5{�[�u����u"OVQ�b`��l�< �qsd�N*�yg1�xXB��/bd X���ў�y�DI�F����C �X���*�,�y2���@�S�[�Q�"Q���yl�� &V���?g�BO�y���^!���g@Y⬉�K��y"�S$;l�B%eH�q	��óg�0�yr�[�*�8�I��s�$�A�����y�H�&�¹�ģ�d04	������yҠ��T|`�Ha��X��Aq��� �y�W`�:��P��Q����V"A!�yRJk9H�S���S�����y��8j� ��\�<�X����C�y�J�,tSج���Z�5_�"�L��yҦ�Z��\TE��-�j�"k+�yb��\�Dp��0%\V���AA�y2��Y0\�2FD �ErPh�bӍ�y�̽�d�7��:��`X\��l��_�������^��#�
}C�ɄȓQ��!�ȕ�[^��$qٓ�&D������G��%��>�|$�i#D��k�g] LڀAۀ�Y/f�^#�a"D�� ������ul��3s��',�""O��!䋝��\cTO�l����c"Oz-*�**����$�E�����"O$`���6��H�U��Z��98!"O�-�C.�%t�`$&S�.H�X�"Op�Fo
l/�Ӥe	#K�ZYZ�"O���ܠ ̮,�edS*t��ie"O�\��,ǑA��H�`
�!nWh��"Od� d��HI�%Ke#F�H8���"O ��DW($�	;w�ȾiG�ebp"O�LD�G���CEB)y#�P��"O0�0g�v=��#2��j"O6a`��4)��`pw���?�~���'�6I�s@۠C���1Bq^v��
�'��x���p́QħY�_+�U�
�'��Q(oB�]yh8j6BV�Y� 	�'�:m"�bP�"���Q�M4eɦX@	�'�*�3��b�]i�K��O��Y��'8���$i�=$�`��F��A����'f�j�@� (h��GnF:i�
���'����/G�q�N���%�)e�.�X�'^��Aa�3E���F�Z�`�J���'��1�Gw�h��*Yyt0�' �CF��8n�1���c�u��'0��hf�*8+l%�#e�
��(�'����R7+8���ro�%~����',��'$޸~���7�6�'�<x �P�En���@?9����'�~���[�4�J��00`j��'PMkP�ŒL^X��AF�R�J,��'�a��ŏl���04�95�\:�'�R�A��&T�(��EL�V��(�'���H�#�(��EZ*7X���'�����jֺ>sE6�����'����5�D=2����dHT�Ƙ�ȓ8�:IZ��m�Ю�j�<�2B"O��� �W�
�ʷH�Tt� "O�0h��i�T��RF���(�"O��CVi�9'�������u��dr"O �S���F8z�A��?wSN�
�"O��tk��y� ;�K�<PR�s"Oz�*Pn�����T͛�J4�uz�"O��i|V9�t��5<>��e"O���iʥq�I���1/(Hr"OZa�)�n� �r.ʦD�0��"O~�:ч��c���A�������p"O�Y�V�_�Upt���.1�\�`B"O^@��"��0�@!�R�)b�x0�"O��[�Q�/���C�-aD����"OA�W�=4�`{c�1D`�@�"Oԑ�wˌ"�J�B�,�yTp�[�"O�9�foW�1�@t���ͥ-��@�"OнA��	B��)Ģ��O-��¤"OFT��I�cX�<�%�=!r"O����\2g�B­�%��+�"On�kD�XID�sI�?���D"O�)��3W�!��d���m��yR�M�P��_#qfe�pO� �yb�¨iX�Ls�O�j�`��6�y��`�n�{�(Z0�]sȄ�y�ح\�Z�)�I	6�L�zB�ڇ�y2Ѧ*2@�Xg�ӯ]Yi��$�yR��W6h 0�+d��I���y�ߓ T8�
D�W!Q��yt�	�y
� x��o� ^p��'\=m�x�"O���t�
�Q�F���؟%d6��"O�%���N�h��	Bdc�&]ڄA�"OX<��rifAs#DMāM!���aV�S1��,#(��ahŘ2a!�`�ę���$H������>�!�D�!W��Z��W�Ǽ��n^��!�d�@�&���5|��,���!�dH8RA�]04�ߕD�������D�!�$��H�܄�&�T�g���R'Eg}!��H�5�X�p$#�,6 ��e3f��$�Kؘ-Kqa��~)�"X3�y���!M�t�E�Β`�Ц��yҋ������s
�)�hx@0	���y��-��m��Sx��mZ-u!�ֵo_V�@aM��.� LSB�5�!��ψ6P�H0�"�&�J�իZ�1z!��$�Y�����")�Kڼq!��Y�������O�H�t<���^�?!��C*9�<��PA�6��L!�,K}��PU�Q>�z�q�M�?% !���H/@m�UFM8�ޡ��M��1O!�D�C� �5΄d��d�@&`<!�-�Z�c���u�0���G4B�!�$��M�� F(@!Ud��B��=�!�DTQR���$X4z;��A�A��o�!���&�åG�*&�H���8F{!���[�:j��Ō}P�󲉚<7<!򄌵$�怙��)
�l�$	ױa$!򤊶+(}2EAO�ތ�U�á.!��"M�t} 1"�X��	2!�$�((��íM�+Q���� :!�$	L�d�r�)F4[���0��;!��N�Q@�1�E�!@�	�4�!���5���ڂ&��4��A�I�*�!�Y,o"�CGRm��ɹQ�Β�Py���yB@�8�Ƣn]4 z��
�yǓ0v��%b��-!��Q�yr��6��]��ʥn�!�O��y��\<@ )�dՖlG6�Y�Ѩ�y�gI387�m	��F�9�&�7�y	D�3�P�sgA��b-@�o���y"(p����M��|ܲc��y�
էo�:#���9`���3TA]��yB휅>1"�X�c��k�0Ы���y�� P�U�e��]�.-x�"0�y��b,�9%�[����OG!�yªQ�s-�mP�킚��q����y��@���,Á5,N��G��0�y2��:|1��� �,-پ�h��<�y��"0eic�\�.���ǣז�y¦ΦsJ� �%z걈&�0�y��7=�M��R>0�I{ы���y2h�� *6Pt�V�	�䂧�;�y��ҘAUH�� 	
�?�NL�7�^*�ybo -e�����*	�ѳ��۴�y�("6�p;G+�vj*���ڱ�y�$PYfub��6o]�a����yRh��p�<*���-a�
�Q��O�y�(��`+�ys�"&ɠ�P0�"�yb�5|�����!N�I &L��y����;���cDE�*GH�3��6�y㉞d��XYWf�2m�L�i5D��y�.C��s$L%l}�Q����y
� ��[��˖
 �V�W<���j�"OĀAŀ�HG�!�q�Y&c����"O��Ӓ�S�Q~0�1iL�G��H��*O�AKb �rGD�s4x��
�'Z�yKA�S2K���FA(q�hc�'ɪ1��W4A�JD#c���tr�'־uK���1K�B���|�<��
�02b9qFj�9Y)ޱ��XK�<OB	}��`Ҏ�9mvha�7��E�<��
:X@5�q��1 |ƕkO�[�<W��vZH���0<i���D�~�<q���:�̬a'��-$"��f�~�<��@YQ!z,�DE��|��A$�Sx�<9���~��8k"�(=O&����w�<�B�W1RX&�ڒ�%=����bFw�<	F�P�s����CK�o�
Ma���t�<��%IT�g�V!Wi �y�Ιt�<��Tf�,d����Qc�a�͕s�<iƒ�-���Fѥ3y��2���s�<��"��H?�4�Œ�}$0т�Eq�<�-U;HR���@�Y�$	�b$\k�<�S,�Tv��f���Y��0IS���<� �S�+ŦS k���J(�tDIB�<�fD�xФ��1ް	�PD���X�<�oX@�(�
&,ߪ%T:v��`�<bg�P�($�j٥N�(��t�<��I>P��!,�,��٩ԥq�<���Y2��1��To+�@+8L!�O��(�7L�>V��!���5<:!���8{��a���k��OGC(!�4�����Q�i� Q�L�!�DY�P��XG�J�<��l����!�
�^�TX�G�qŸ����ɞH�!�d@,Z�|�@����u�� u�K!�D?W�;w��(j��P�
I�!9!�Ĕ�!b�{����#n�d����#5!�R��`���Qt]���&��n!�\��(�`V�P�bG>�P�%ПH�!�DK���h��L
*A��Y��yy!�䊪Wp�u����~Ft�b�#׈c!�C3���b(�6b�b�ڱ"ja!�U�@�и�bh
7��;�]��!���QɠH �5jP���4�_D!�͖J��d@�1��ړ�I^"!��؅"�*�Є) ��Y H� >!�DF�-�(ѱ�

~�l-�@Hŧ
�!��SȬ�R��p2G�Y�!�$U6���*�D��X�g�!�$B�(1F���W[�h��Z �!�)-��c���]���t�+#G!��V�t7"ѡgA�r|�xaVZ�x/!�$�8s1L��+��es��m40!�$C�x�]�MÃ{p���k��!�B�X�԰���U�hA$��1�A>!��\gQ�`��d� 28�˷F�$�!�^�| 4�Ҋ>������!��-i��b��x��b�ի�!��j�����5R��,F9O�!�
� M���; ��@��Q?o!���EX�	@��9�hm�wJ��.!�d��i�����d��f� BS��3!�d�eΌ��\�N�4��q�P:m�!�$L'Y[���uA�8��I!;k!�D�&R8��2s���fQBe'ٙ{_!�� �t�'�"	�ڸ��K�/BnPl�q"O�P#Ћ6�����OP��"O�m�v,P'V	|�i EB��i�"Ox|Фa	:_������}x�$:a"O�%�$s��]y"�7~�)+"O���GM�%\��a�!�԰��"O�X1�ɶ<�ؽ����v�����"O�u9�'�����N�au��3"O�$A�"6 ?�,��"B�]�9�"Ojr�]wݢ̸wύ&n'p��"O�������5)6E��}5J�"Oh���.E�|�1��
Z��Kb"Oz)�`�Z;���0MC�f�S"Oj��L٫f-F�
6���{����"Onc���J68R5$�7�j�{�"O�H�d���d���-}iJ5"O�
��=>(!X�)�VQsB"O�a�v��*e6�`�>~B�!"O �;��ؗ��	3R� �MB& �w"O���TD7L$=#ua�#b�e"O�U�"��Ht�#�/
�"Z"O��bw��<c�d��t�ԌQ+�!�"O!�����aq��7�p}B�"OJ���o�?@���B6e����"O2�xd	��vVn���*^�F<ܣq"OH���aů{�8���z-n���"O�\�� �.x&�ēv��s-�!��"O:�
E�V8�b}�K�}`�ȣ"O�i�TA=�
L�� �/L�1K6"O��{�EB�y6t�0��գz<f�2�"O x @gҞ/=�t��G�u)0��0"OI�`���L�gD?�a�"O@Ɂ
Τ	?,����*1��� "Ox5j�oDٴ!qfD�/��h�"O��h��ʏ	�
�����^Z`�"Or)KW �7V��RR�¤$��˓"O2�t8��5���=$^�H�"O�izāU�)*�Y�aY#�u	C"O���B��1�� ��B�
p���ʣ"O�|��<e�2�2�#Q��چ"O�5be��Hm ��  ��Z�r�H�"O��!��P�<�Q�V)bz�0;�"OP��<C��\@�ʖ�AE�hT"OV���)§
1&��R�W':i� "Ovk׼��|%���hh�t"O�L��痂Zj ���Ǎ!hi1"O>Ă�M�589`t�D��dS�͐t"O��i$��	2�����&>��"O!
w�Y=,���1���L���"OD���-�X�VL�E�
���z7"O&%q��G�K%�Ё�C�5���%"O����a�q��,�l�&:U)"OJ����v0�8��C�6vRe�w"OJ�ru7ª��Bl�
z��u"O�(�2�ųs �� j�=k\`�8a"O�Ic���N��T����04�|x�"O���lһr�"���H
�2��� "O��,WK�XQy�H�3�q#*OH�����	�S/F�9&v���'� 1��3N b�MV�*�p���'���ۄcl�!�? -J�)�'�డP&�39�����JI�L���'���!��A�F��h��LB?{��'��x�g���=�lU��bn=1a	��� ��a���c�^4&d�3jL��"Oڴ���62��T���S^� �"OJ���oפ'��ݐ���6��� "O(-���88�U{&�F.F�!��"O�i���6b���A��K�<᬴�"O�}��a�<�c`��I�")Y�"O�{ƪO= ��� "�Y��!��"On���N�XBT�@��A�ppt�"O4*��^#b9*t�ӫZY*�e"O&m��hC#'�fL@'�0|w���"O�M�v"^x-ΰ����pnx��"O+�,�,��4�QK��DS[#"O��4�Y��>�-IQ� CA- �y��7g����%�P1ʱ�!bA�HOr�=�O�2�1�㕼g��	q�埌T����'�z�8p��D��δ3&���'�zP`�D��4�Q���"p`�'A��0q�X�.L����,��i�'�ў"~b��	p׺X��Joa�x�#�~�<aK�5�����Ḃ`�`%٥.�Q�<�w*�:!���Q�,рVb�`j&�i�<1�j�;\�1��G!3_���n�'�ay�N�F��+�
L�*����о�O0�󤌩9���@��y����G��&�!��/=�Va�#�5^��0�P~�!�P��`��L�=}\)���[�!�$6�
3�O�<=���d|�g~��'��Q� �&���p�M�.��"�'�ў"~�è �=i�)�p�R��e15�T`�<iǧJc�ʬ�!*� :D�w�\�<�� �:|�b���������R�<�2논A��2�����q;���K�'�ў�e�p�i2ΗI	: P�'ֶ�@�ȓlzH��4��H媴���*��8�ȓ6��C#	�7κ���An�ȗ'��	r�)��O�`���L2�D	h�Nʾ0�����>�	�c �d�"�F�#Z���*Z8[<���(�� ;�f�P�����j��n���A~��� f�8q` ۼz�~�i0�F�y��� s�1aJE�_�tQ��K��ydK/<�.��fҷL3�����'aўb>0�H�xy���j^6JSH �Q',D�Dڤ�]�$>H�c�[���h"�$D��{G�ɄY"�!-rޕ��,6D��q��B�o/�1a20���X��5�O|�'J�=Q �R�SR1H�D�i�d)S"OXQ��+��jb�{�,�7_3���"O�;�,B����a%�P4N:��"O�dQ��47bx���;
�)��"O�U��/�c��Q�J�%_�,Z7�O����=a`��t��j��$h��pX�EKI��؛5�x2�KHƎD�b�
%�u1�L���<���׿ d��B ��\ ��UO��g џ0l�L�OM����Tzт�
���'(zx@S��$?�S��,�K%F!��R�x�� �!4�~R��X��O�>�ju	�0f�Ĉ���"px	���y��F{�����|��Mg�U9�c�	���Px�ؒ�9B���w��L���4OV#=��	Q�		:f�=pq��@�	K�<)lͩZ
�)��H�Tp ���I�<���n��頳��6Q�xU�4��y�@&�A���nA
�b�X�=Lr���<D�X��� J�D㴄�s��U�&�IW�O�Oe�\�Pfӡc(�����	yvd!�O��
�S�? ���W����*TT	(p�B��<$�x���!���ȔO	�ma\�¡6D�0b7�EjZL�4�Y+W���>�RP���'t*\3�`Ά8�	�wP<��U�y�����X�Npa@�џM6P�g^���J<E���3�|Т���wr"懆�+��F~R���lpdhb��*;��Q6��C�|�|b�듡0=Y�`�X�Bt���*Dܼ����tH<i�G	^Ze���,��D���̫;�!�$�)m���"y�)���ų ��y��6a$|�cO��uS�YӲ�]C�B�	�a�ƹXg,�!\�1G�b;�O\�=�~��LYm#��a�	�Lh�F�Em�'��x2)�	1o��hW�T�zT�8U@��aJp7�&���%Z
�����C�:�1 �6� o�(h��-ɷCf�)f&E�+�<�K
�''Z�(h�t�@�6+ $"=�i��O���G�4!ɗ{�0ȣ��ԃe^��!�]��0?�*O�9)�F�S�����,��y���OT�������(���bs@ ���c2IS�t�v��8��CܧA |$���]�`:��K�O��8�0�>�דz6Xx�*G7->u��lSE(�D��0Ӭ���Λ4u�t�Ѯ�3��e��I�<�4A��%���
1U��$
�� O�4$�i铨Mۋ���9\n�aA�?G� h ��E��y��4�� BF�A"\�pơ����Y���O�m�T�A�iI�"�-d�x�����"�'V��|Â ���ȝxq�'bp��ȓ|lv����	�p�����Dr*̇�hڜЕd۔TK� @�aL#�^��ȓ$�%�� -��:�)�7�j���/k�E���17*�Y 睲z���<i���)��
�$iGh� U�µ��
E"!�䎛pP�#�NL�r����hF�f���@��H��1�ףY�hH\d����Yx��a ;O���01�،jwj�}�h2�'T�n�!�D'(��5x1�U�N"4c$���a{���ݗ#E�d�ŉ�,<���xBkJ,y�!�	�:U���9_��d�'�]�8{!��6aW�eX�G��~������@[!��Lm��@�ЇBM ��50�Q�8E�t�޼)�tA�mO�O�(�C��,�y�&˒|��D�%*�A'��˲l@��=�{Bk��k��#�/.1��dK�,ܰ=�{�	§6��#�/R�l�ybA��R����w��2��d����?	�'s����.&f�+��4�	��'���Ţ�R����c�ƉFf����{"�'t��Ѿ?hV��g��fr�I�Ah:iC���l���� 	�V7@��
e�X���	~�	�r�<�KZ;5cZ��`�I�C�I�WyҭqŎ��z��YbTEͻg��F{��9O|(i`F�} m�r�ٝZ���'~�ɽDMv8a�gӬ��	 ȷLaC�I�?ese	ٲd�xx����>/��B�&SV��`��>rv^�g���B�	�J:>�YA�ѭ�B�s�
?i�C�	�4n��#lع2�BPÛ�q��B�	5B$�%�>QH�����=
�B�I2u~R(h��=�:< ���mZ~b� E{��4��"v��r���9ݦ�j$�Z��y"�8;�y�f�v����o���ē�hO�����D�M��� m��h�l$y�"Ob}x�&dklд��
mص��"O� �@xpjڷƌD�Ɖ�LD$�R"O�E8�+4FO�8"q���J0d�I��'��ExF[94��šKhz5�fސ�y2��P��TBQ�g��Ё�y�CX�-�(w�wUT�3�A��y2�#h��T�u��p��Y�腉�y"+�%7$�ZV�U#lO8�c��B��yG�
Y�t�(��'X�8�j!��y�o/[ظ��C7_8.�  ��0=��Ҏ[��}�G
b��`���y�a�Ę�w�V�^Rb���e�$�yR�J�9����tkЭW���S`�T>�y��P0h�ht�S�b�+�9�y��ϵ3y�$����I�ڄ�a��y(ܴU�bQXW�߀F'���JF��yb��	�Z�hWC�i�"�M�y�I#�5p�D;[������y�o�.(��8��N��hpa��y�H:A�ށ��IX�|�px�+���yB)�,Z�&�S#�n���(g�A �yB@B ��D����g�L��F��y�M��8M�� U�e�	�t�Ş�y��L�e�8���d�MR�(O<�ybnTX��M�eb
=%�>���� �y�*��*K�u`�%Q���̌�yb �od�1�gF���(!�F�5�yb��W$bT(��ԛ��u�&��>�y�ō+������A�˨uc6���yj�:��Ӡ'�ر2�T��yb��9�8���@��`�&�yB��<-s6]"�R�>����)���y�(��(���!��%�:k'cA��yBH�(v���¢��$�:��@�?�y�ğ(rn�r�Y."d~y�����y2"[�n�P�#J�c�B�+2����yrOŰ!8Z�YR�ܿ]��9�Mݶ�yBK@����#j�v� ���yB#	�M�<��K�	z"+�8�yB�B+��8ũ�Z*Q�ȗ�y(K?1<J�ɀ`��@��a�8�yB��-D�2���I�m�fp�a/���y�D�/X���6��T�l����y⢏E��� �d�1L�\E�"LL�y�A�;� 	q
� mM�A[r���y2�ӡ>[\I�.�����Tnˀ�y�I��z������!a��֣��0?�!�J�r�CD�J�4uɄ�K7z����P�<�!�?|�-�P-5]���ɕ�N�<�'�׸ qB�d�)R����
p�<`M�o���)�ē�|ظsF<D�p�iK>|�L;Ɋ�u`�����(D��� ��?oJU��!� �hٺӃ5D�L�툊;���!��N�LI�<D���c�V�(�(p�ԃ� nd0�'�=D�г�/T%]V(��o%Sn\%��&D���οW���դ�& 0	���0D��cŦ	C�(���]7%<Ar#=D�T�W��7gZEx�d�H����D8D�蹗��"��zRe �1D��*7D�<H!Ŝ$�����+E1ǠT��(2D� ���ǖv����tM^>�洱�D%D�<�ʊ\͌iQ6��>R��#D�����H^V��2	 e�� �E�=D��(� �7D�Aaq��t���Vf<$�,�� �� Ǉ�>5Á)ѭ'�(� ���
px�1���p>i ��t�HP���_�geh�"w��M��+d�J�g�413s���B}l0��$*Bv1�`ꝟ!��h �A�V�8C�I1�8��r�������^?0B4ʓ2Hx8����;y���`��(��"}��.��q� ���.���5���o�<���D0l.��葚Lc$m���){HF��i���&җ�2�&>9�=Iqʔ�q���bGĭzV4��$Ɍr��L"�L�(Q[f� 5���kH�p�$*ѝ�|����Q�� ��dLI����'���+�I��[^��D�O��8=����z�>��'b�&�Y�@\&%����w��
E��,a��:Bzfy1��ցH�\C�I����'��p�;B�%-��dO�Hz:Ƞ��W8 C��i�B�����g��Oz@8{�O�wX!���Ȝz�
�j�"O9��
-��9�`]Ch��RȐ1x޵�®X�S�i �`�-��:`qF=p��xb)�����`�.w���y�΃���>�ӆ]Gd =����3d� �ď0-V�ac.��~S>�+��JI�(۱��4�&����H��� ֜q���ήU h�DzR�� M.@YrQn�,X*�'�(�`��Ă�E���av�S����+��Ȳ9c�EID
O�Ap��&�xe�7%%>�hƵi	���D�.��)�T��Ƭ � �.I0��p��\clfD���4
R ��bԕ�Ҡ�	�'βc&�W������>�BaB!�
�c�n	30A�h�����K%��i�
�jTsvG>}rM�p�t*^�{Mֈ  FQ2��>q�̣g����� :a���'���L�)
�s�k�=f\�Y�ϿI�ܔR�+_dy���(&�Ů�W�( ��(nR��ʦK�?7ZT ����-s ���mr��уOG�1�P���2H�d�Y^(<�����݁�NI;|�Hp$Ȧ�z�/�=8w�y����a��-"�ݓCgR�s�a��U���!C�
L�`hQP�N�y��@�fpP��1��pC�Ủf�2�0�G�����ۼnan�X����8�N�9"���'lV}���(�`x�M]*���!W�!�1o�(k�����!(x3Vm��{���%n���)z� C5f��IP.�p<�g���T��e�AŇ�V��Bc�z�',�����+Q���"�X(mL��A�<hpW
�c�T��Rf�	�bÄ���p����(�R``�����x&C�8fЛ��
��D��#Y��rDC�"Z���(O7��5��^_C�����L6�*|�d���y��Io�NݲWF�0ӦQ�Cld��ؑ���/~`�	c�Z>�b��l�3��L�j�8�'zΐ	a�Æ�V��'�!1�����C`Ju��O�1)�A��,c�+��V�V^��b��06h萒&ɳFbK�H�p<A�FA�~�� ��^8�t<AQ�@J�'(��q��$;N�藎� G@��	n��ӓ�� 1m�|[l�I�u ��[{H<�1�S�(��@JC�x%<mZ�a^�� ��O�6�p�'"'V虣Qm�*��HZS�)��N�� ��03�`����B�B䉘sC����°�2�Jd��-�8�W$A��&��èF��m#փ���,oF8	W�̃3�	�[U����	�h춬9�@8�z��c
 Lx��/w�
��iǙ<��5 ��+~Zaz"/���p���X�,�C��O�e�+�-���x4�;24�����ކo�Tٰ.-L��h���F%�ȓ7�|#�o�)��=���'e�U�'
�4z� 
d����M�݌�G�����2��1p���Z4A�Î���yҋ�7�.h�T\5x�5��J�6��Lb�6O��N�9�reK���y������h3�x&t�x��x҄A)��Q�GI�[�,9���@��򬟥�����'�� QtA-BH��W��0ؠ�'b�tK�'V�)�>�@�JجvTl �'�J�F���Y^ฅ-�6�� 	�'y8쁵�ɜ	Z� P"[<,�����'�H�A)X	����S��>���'z�̊�	øze���$+=W�)��'��eb�_�#���sca�93� ,:
�'\ޝчWF䔐����8����	�'Ҽ�{s�ڞ��u�Ńa���'�&���AP�v �Y��N�c�B��'7�� ���<x���.w��|�	�'�B���(��zŐa!AOT�h��ձ�P��u:�O��SfJ�s�.�zA���p���4"O�YZ���^f����«H���D	��d���3� �A�b�"��	�`��-	�"O��h5�_ |�0�УhQ�ԃ��؍S���O>���>���Á��2L�9s����ٹH6!�$���9�f��fR`	E�E�i@��б"��
��'�P�O�M���FQN6���6���b)F?���&j�A&�3E
�����[���=i�/ 7�p�/��L��q��U�R)d0�Eپ�H����5~��2O�N�%[�΃�+�&B�	3�lZ� �'K ���F>f�&k`o@$V�'�(��j�g}R���d��ä��/�fm c� �y�(n����+ڇ)ĺ��gbE��M�m�G�hY����̑PIN1�ƥh�&�2aV����I8�ܬ�,Jt?)g��7����>���:�*h�<	��S =>@��5?f�L��Ef��HH��d.g�O��0�1/y,�ّ�HZ�_s��z�'7:h{a�X�@`��k��J��	s�C����"~�I2,�c噌bz�J���r]�C�I.mDj��@$LZ�h��ӂ33B䉨{���5Y;G��A`��Й{�B�	(�b�W�0�h���@!a>
B�	os�<񷇆�(�|��5O_�[�B�ɏQ�0�0��
C�A8��Y�S�B�ɚln� 7��@���H�Y�xB�9��@x�B!�,�"� �V�C�	v��$�UM�.M�$�1 ��R��C�*br�	�c �����Δ.��C䉓iT���W�I���;$c�5Kc�C�(\:0yto)E�k�$}�C�ɛu�Z��'R	
22ht�̺;��C䉕`�� �D�Q��,���^U�C��9!ѻs̉"Erq&&�:�DC�I�#�p h��ҳy����e�B��O�ZI
6�"�� ��)���B��,=�l��+W�ޤ�ǁ3�B䉰�l]�1NĤ���C�X�9��B�ɥ��8 wGV5 ��9���-r�~B�	� Ҽ4�d��
N�(0s
��Kb�C�	�T]"QN_=!�y�Ќg�C��Z��\{�o�"�$j�cL
R��B��%Y�4Y�b���lB�P�
H�v�C�y*I����-{�]y2@�PQJC�	�[��!6"���|�P���.X�@B䉇dX����B�H��g�K�!EC�	�m>�x�(1�D�p����B䉹\��x��b�����L�4D�B�Iz���'���d����6��=#��B�I�쉀�J���|)t��52�C䉁!̎���H�; �bȂ��\-#�C�	�4�	�bH8.琜0$T�RqpC�	�dQ�a85CZ�7[F�@@��	�DC�I3p_Na��B������E�zB�	6]3����?n+��z@�Q>�B�\%ZX�D����M�q^\C䉻uz�|�Q��p�eI<��B�I5\�T1����
S�E4jǮPX�"O��`���s6�	�n۝F�`���"O�ش �o���q��Ї`x���W"ODe��$�*N����9S>t�a"O����NO_vhCD���j�s"O���b�.;c�uj�e�.�� ��"O���p/��?� M�<BP����"OXl�"���x�:������t��"O0�{@	Ak�@;��*k�\] "O���F�ГQ�����[�?�����"O� �<rQn�<���*�-G�*��h��"Oh�)��.�*]�rK�S�b���"O���5���~�R���5�X��"OڐpT��Jɢ�Z�X+��!2�"O��ꅨ������ډ6�|�c"O޴2g�!}2`KFf̤I��|Zq"O^�R�ȳ__td4�ӷ
!,a�"OX\(��78YP�@4�E�0#�%�""O��d�İ|1�ɑ�du(y��"O 8�S�L�zeLpcB��3Z]��"O9�ƒ��$���X�J):X��"O���*_a�&\1�b��j�|�5"O��� '1 �b�ˇ��М��"O♑��E�����o�4��A"O�x2u�Uep��e�
w��A��"O̼I�-� ]�:���X�߰]s�"O�H�P��dw��)0G�g�~�y�"O�I�3y��d�FL�Ǌ����|R�)�,c`�urҧ��Ac2��bT�A.PB�	�^��#� �C����dPRObB�I4\�x#uhZ���)Kt*X	Q�nB䉄z�t�q�� P��
&��%x�B�I�ge����K��,�c�07P�C��OkBѡ�'=$q�a�Z�~a�C�	?D|�����u��]�/�1I�rC�I�(^����	Jr��0�cH,4�B�ɵv嶡�̈r���t��J6�C�#$VVL�A���Br�j!�ZMb�B�I.gM�%;��C�Q0���=ǌC�/7 ��o�Q��7��k�C�	
(f��"�+k.b�{g?�����7 � ��Dԥ`>v�e��#�!�Y/O�b�qp��s���Ðs6!�$ϗo���QE̊R�RׇF>!�?T�S��	�}����&3`)!���-?5��Y��E<�p:��Ͼ�!�D��\c
E��� �طK@3r!��0�I�Lc�(9�IB3<`!�DJ����t�\�Zh��I�Lp\!�dY8S2x ��lA�BRp�X���wX!��'p�R" �1.PCf�>A!�D�5���c�#E\P"E��!�a��!zb�V8*F���T+5v�!�d
�,�9xR*W0[�P��h�gf!�d�(R�#a+Z�g����A!򄔹d�$��F�H4$<f]0$�cC!�^U,��e#	�y;>rP	Y,x*!���0yR �7e/�Z4ȍv!�? ��嘤DK�I�Ĉ!Ǚ�|�!��\?9��B$��T���f��!�txF;L+x�8�M�(��p�*�e�<q���G-%z7�.j,q�[�<�A�@$!��]Ѵ$�nٶ�Ѧ�Q�<�q�ǃ.��
��I|��q)vfAN�<Ʌ�(;Z@��.�xw
�Ȣ�O�<����K��1�Fl$(DL��(M�<I2K�T�`���U!t��X��	D�<�� �7r�8e���1�B��ΈB�<���.4E���!IP�y~�$���C�<!!(�Q�a����}�8�� }�<�N�!U*<c�^�G��a���L�<�d�
=
ƎL���U$9�I�0�H�<�V-::��Bˈ�pB��Ue�O�<��L�b�(A�0C@ܡ(q ���S�? ���h��um�}�Ѕ4�}��"O>��"�]�]�aCBU�x�$x1"O]�4�a�`�0�1J�f q"O�y�aW�t�6E9-W���$"O,}���@j9��e�R+8U��AC"OR�KI��&K���E휸SC"91D"OJ����t}bۦ�W:,^�qa!"O�ۖ�tud�PQ�E�Jd�xs"O��#��̝g ��PDN4@Aı*A"Ol�37�	I�،p�)F ��"Orpb�*24f�$�S�^� 8.e��"O~�8�BY��T@*E�;/(�p�"O��� �
� �P�"V~ �M��"O�Iz��	 _�l�!�@�,q�F�jc"O�8їW�]��@�P@ʀ(���a"OPQZi�9a]L�P�9���"Of�5 �?0r�k��јC��XQ"O\��������BP�םL���a�"O�%s���1�@��3��2���S1"OBЋwoX�	��xp���.=����"O��ҩ�$�E���[��Z�"Oؕ�#!M-;rn5
��*�ĝ�"O&���]�^U,;g%۝t�Pd�G"O�����pȞ4����M�6I`"O��9���*P7���CE�9N ���e"O�U�rC2�d0Ç�K�d}�F"O\��dkZ62D`͋��mqvYg"O�5�ꐚ{ �(���
�i�r9�g"O
��$�͐^�Qt�NO�0�y�"O�0�� ��,EpF��/�b0��"O̘�0$�I���0�%��w`uQg"O�PyR)
�)�>884�X<��"OV-�g�r�P�
d�>�"O6�c&&K�mV��˰fU":���5"O>�C�kS�jTJ�dO]5v��l�"O IC��F &�xd1G'B A�9�"O�AȢ�  g X��O~��ȁ�"O�m��;0�V�3�&�x���z�"OB��������^�g�|�S""O�0S�g���*Fm��+�2i�"O���'��VdJ!�A�O5"�jz"Od��gT'1ڜjA (��"OH�2cIw��Ոw#h��v"O��ZW�>d�5 �h��3	��j""OB����xB�qSc� �9�P"Oz,y�[�"����f��vˠp�"O��S4eX.0 �W��Q�T�C�"O�]��� #�X�G$T!s�e`�"O�sJ�?�P�s��IJ}��"O��9�ʡr?0l�!'˞-d���"O��PG�I�f�H��@�3�ڨ�"O����*�#^���8�hE� s|z"O���f�ƪ	o�(KSlN�1x"Ի"O��� ��&KZL��,�%p]@�"OexD�énm&�R��w�`�"O�E�S�V�]��IqE��z�b�(�"O�aC%2 4q�4���%w�`��"O�h$�Xjv��$��Wm�0J�"O4�1wO�q�l��I[*P�"Op[�bC5ܔ��5[\0�'"ON�;�f۸c:0�9��®[7(<)w"O~Ъ�fŢo)�Qʜ�'vQ�h�<�E^c��SХ_(6+�)�0jT�<Q0u~H�X���OӶCfd�l�<� ��y��J�(hue�'�hac"O��+��'>��A�wĆ@��'B�7J�>QR�E�8�z�:3'����:�Ř^�<b	M�}H�<�qj�f���:4B�q��^�LVd�Z�O<��A�ϥ=���M�K[�m	���ZQ
��0,�&� ��g�ΰ^�L�I>�7�>�D�29��:K��@���*���^�<i���]^=p��ؘ<����HۦQ��
# �x��	�*��A"��y*Ԅ� :9F����EU��:E�d] Z��E��
4@8!K��ɼ=<!�ی(��	���E�kH氘��Ff�O`��!�؄m6��~�u�W!����&�s$>��Wb�|�<qKլ
&�ɀw�4+��˳�D�2�B���9�$�y���$I;U��!b��K��d���!�d2W���'.R�u̒�C��vJ�<��iR��'݆R�����h�dՈG�i��lE��JAȁ��~"d*J̸i�n�i��"����yR�Ǔ��܋a�QW���Ơ��'B�� A؎���N�fBOF&0��?���R"O
��T�����c��΍>�@}�ѧ�O^��?E���Z�"x�2J
�}�mz`��?��ȓu��{�ƅ�8�&\��4C�؅ȓw��5닄F��9"҇kD̵��w�R=@`�ٰ���y�DV�%�����2�du{Ԍ_���b����-��O���%�!�(�1��E�Q̸,�ȓa�0I��A�x�z�I�&�S!�i��;�45ke��"yFAQ�jP�e�$-�ȓE�arA�/P�s�˚��Ȅ�S� �5��"�XԮÑ�؄�ȓ0
"��`x#FG	O�����G�ެ�v��S<��"��  �\��;S��X`�ƎS:��(Y�
w�?D��Q��H ��P����R�lm9u&D��b1#1�hB�!L-\�y��)%D��kV,Q�*��Tr1�,��4�@1D�pд"��P �y� ,@��,D�����X���r��"��(�-7D�������Ȥh�9�ָ���2D��ʐ�,s��!�2"�Kq���$$.D��!�fL6�T�:���Pm��,D����n�4��v�J�2X-�Qj<D��*�X4 ���a��I0]��Q8Vh<D���IJ�;A�d\��Ѐ�:D��(r%Or�&�sGmļY*��K;D�0�KLLmr��$�CS{��*�*D��p�Zxd�� ���o �5`�+D���*_*ޞ��3e)�0�PE�&D�Ĺ�)-���ã��f����ek#D�x:�O�}U�B��n��S��!D����*��� )Fm�!�B����>D� pT��
Y�vˉ�BĊ�	��3D�
@���K�L�v�ج���.D� �۩Y��3�P�RO��{��9D�i"�*���{f��F����I6D����8�>0�R���I��0D��
�NJG��k5a�h� �ץ0D�D�vF#���+���;2Q��#=D��(uŕ 9�>��� >?60�"�4D�P�5g�&Y
PA��g��^cL���>D�<:e�����4���!jVES��?D���ͯO��G�;%��qAf<D�3�a�~�\1��Ȧ^���'8D���� L ��Q�MƂ}K���W)7D�� p�z��W/�Ջ���e��HcC"O�����&%��A��/c:�"O����ς|\d�S�Hл-Vm�T"O�H�[�@2!������,��"OD�y�LL9R�P�ڸ ����"O����ڲ}�p��o\�7%��2�"O~1�a��/whp%��v���5"O���K�)���Q�-lP�0�C"O�9�a^.[úX8��;[A���"O8���@�!Sl��#�-u9b�� "O����AɥQ'�=�BO��<���"OR�� �ԁbں�x����B "O�8J�둬1�V���*��K�"O���#�䃷�8��|K�"O^��5�`a���!�=�b"O�Hbݢ`J�Ca�N>P��"Oj�(5(���j�`�*|��q�"O�L��A�)k�1��Ŝ>�Ԅs"O�cD�]�e�Xy�Ĩ&ڪ,�$"O�qY� pIl� È�Ʋ!5"O����&��HY2ǡ�1r�&��"O�T����p�f�I �S<L���"O�re,�V�H��i��k���yBG���SQ$ї+H0eA��]�y�A��PD���)�a~���
��y�FR�P�u��`����Å�1�y2G�����S�_�
֒�x5N���y����Il	9�!7k�<�4JJ��y2�(FU6��#���\Rz�p��E��y�'�1]Y6,ac2]I���u����y� 2)��s�HO�EB($�4C
=�y��д16Ū��'GY�ZɃ?�y���9?�hd���e����B,�y2(Ĺ7P���@$�"xHEN��y�M+Q��3,�&�楂qS��y��ʸ$���i7��:���BB�y�L�:_��C�D)-��2� �y҈�c�0��e^
�� 02KC��y�PVQZEXQ�H(���B��y��U�:��E�Cn ��oV�y�Κ3I���哀P������yR�M�RNQ!��=^i4 tL�+�yBI��S���Ð�V�j�ʓ��%�y��B�f�١@ݷJQ6Գ�cǵ�y�FH�
B����38�L4�����y�ILq���{0mȷ- �0 ���y�),lU.풶��t��[ a�y�BO�oX$� �i�2�:�H� �y�+Z�C�N8�#L��n	��k� ���y+�.L�t�C���.�B孊&�yM�)i"X!Z���qN@aE�4�y@�*N�V��C�j���C킮�y�l�币z��7f�H���yr!Hk��`SӍщg�0T#5,�;�0?av	�O�dSg�-b�{��O�>����)��tЂ?�y� ����,n�t}��i|�Ӻk�����IЈb�&|��'E]}��)�'>��E�e܈xb�HeϏ�C�X�ȓ1�j\��M%(�|���75I�E{RD,�'yx��ks�_�:�]���6^��?	��IV���G���f��uc��j��2�'��DEy����U0~bi�G"s��$s��M��dS8�(O�>�ڇ �ј,�O��ޔ+!"n��1p�)�']Em��`� ����00؍��@��0|R��4+^Q)���z�Y���C�Fa�<%>� � ��C^+f!��HS�T
��xR"�3�O����±	˞j���2i#>zD�fZ�PK�'.��^�O���`�.>=�6Q�Ki�bYB�H���㟢7��"��#�<@��tϋ%�O�}�ç�j ����7K�B�ڕ�X���>9�L&�S�S�D�T���ȜC_*��IK�
�O�P�7�)�{8xA{/�;�(�m,��(z#<q��)����F g ���BD�Y���_��ȟ�a�E�܀]�4�3��N&CNJ��;��a�D	���QK�HwQڄ��n���'�l�GyZ����p���BeՄN��qI�M���'��#=�~��ᎇQrȬs�,6��b�(�v�<	�,��ea9��(�1�m�d�<Q���Ӷv�p�RC�=�L�傑 j���Ŧ���N���р�y*W(n��5)�Ҭ>7r�!ÿ`���Y|l2��'�D�gR��T�XS�&4)�'�$������M�Z2��{�h�
�'��\�P���;��� �ۖv����	�'5Z�CS�F09+��P�tD:�'���堌�U%^1�CΫ}����'7R�Z�K?����Q	Z���0��'[�)�pꈩ9�	��^�&M�'��+�H�8��`�����P�'B,▢A�k�H��%�z8`�
�'�LT͌?%�Α��^�,X*�'S��C�{��"��"�-��'-��1���3݈�@�
�)ب*�'	�(«��gW���#xz��
�'V�$����	j>B���=v*�)�	�'��}�c�3���kVrx��'�}	�#�v���l���'?�x�	��Y\z����4\��'6�pq�o��a B��&AҔt����'~D\�@�\, ���I��N �T���'���S�gK�@|��!���mN,Q��'j��"b��I�H!���ʭe�
Ms�'Ϧ������(��C�"�a�V9��'�Z��,��4Q@�3QK��Qa.�)�'`�-Kw! �7k�Q����/�"�1�'p�"!�K�	֌�0��&@���'��$���3AN<�GJ>��Y�	�'��("�t��R�U0C�
�
�'[���v�'�-��i�`��L�<�eH�!����[Ų��A�}�<9�!�\�xa@'Yg�!�o]N�<14�+Sh�e{�#�H���uϙK�<�'��=�D����; 3|�0.�D�<��j��=s�Y�e�B>s2�X膨Y�<����6�s��u�.�����n�<��m\d<IL&1��-�T�)D��x%�̝��pR��i֜r�'D��L�3Vu8�ŮO�b���d� D�lk�J��ڍI@H�Ub�cg�9D��Be����-;AH�JĘ�s��7D���Q���c�d�1�.5�k�H7D� ��1��I� �Ʀb�ax�6D��q�H	�*^����<z��yE/D��qtG��_��ak@FBX���Ӄ?�hO�Tܚ8��eX:u��3U+�<��C䉌r�(��ǘE)�;Q�X�5��C�	�n��К���9E֡q!�lbC�!�J,\]B��\�#8��@�'D��Rf.�j`r�
�U�:L %D�`���[�fhd���� X�|�We#D�� ��B�k�$ f����!c�6�;'"OH�UΗ 2�>x4Nñ|q�H!"O�a�#�D&y�-:I���'"O��XAŚ<;ܐ�L��e�R��E"O�9GJK*�h9���ܪ2���r�"OR�� �dm��XT�ڛ^pBW"O��$T�&}�i�(���8h�"O|U�bR�I̊�fؔd��$2�"OĠ��C��}j�X��Ɛq}<]��"O*��ɠ��sf�cxLi�"Ot)�Mֿ2�~�(Qf
h�&���"Oā�0#�:}rr�0D�L++w �Y�"OЀȗ�I�*��-����ZO�<�¤�7sP� qI�np��s��N�<��MK�9�Sw�ȋwr�tC���f�<��O�5.�|�ɰ�/b�t3�o�a�<2(�*THT"���GX��.Gf�<y@����H��;A#�ъ7(Ib�<�w�,
P|Q{p���Ԍ� m\�<�c坑Vh�ѡV	c"!���E@�<�63gw5�s@+
���d#}�<1�k�c-��/J�o�<��ox�<�&�.�]��+-�>)1��w�<���>H���̥,��]S��_�<����#�����*(ҍ8�U\�<�&��=UB�X��Ҡ"�6Dp��o�<�Dj�>u��]��ĜQ@9�u�`�<qv�R
���D�ug�@���^�<Q혔q�p�a�)��5Q�o�<�u�)X�%��a�h��0��a�<U�_9\�T!$j�j�  �e][�<	Ƕ4��Y��>0~p�c-�T�<� ���b�l����_>w�t���[�<A�m�-L�� `F��9R1��2Wl�l�<@%W,DȈ�@�H�/
�	���r�<��%��3n�;e�U"Oװ�k��n�<Qa@�?�y��G&c��P!�q�<)f�Ø[�Z�5��$D4�c���a�<a�ч#��e׹p#�6C�\�<ɓ��+��B���)�R�scB_�<���u��}�e���jlRP��\�<�#%4UuQ`,D.*C��9�b�Y�<���(	��9�+U`1��GYV�<fcڰ:[x�{B�B-Rz�x�Gi�<�6ڿ7/��r" -@�>���jLP�<1%>>��q�jՃ`-[G�M�<1����3|�tc���]�
@��E�<a$Œ�*^pj�'Ӹ=���z��F�<�P�F =*��$�4e���Ʉ��D�<)V.^0��� ��'tZ��m�J�<a�(	�KF�g�,/�^� ��}�<�DG�3	JF�(�`ݼ��Q�x�<ig-H�7��0�׭B�
�P�Ɉ]�<��cJ5Gs��!A���l��4�s�G^�<�Q�^0� �)S��,r;Z���Y�<�uB�*O.�:�'���*bS��X�<�M��0� 5���	���1�H�i�<i��^3�4B �[�1�(m���g�<�FE
$os���RZ&�e�s�D_�<���_�mo\�8�F�\	d�y�*�r�<a��
@�\�afʉH�����(D�<)T��d���*r!J�2!u��A�<��G�":�.����.�Dub0�X�<4^	���
Y�W�r����S�<� �!���Onu��#�nI�P"OjY0�J�yE�ٱ$�O�g[r�#"O���4��O�ެJ'�K4E>l2�"O�� �"kE|��/�w8��w"Oz<Qa�R	r����,%V��a"O���,J���ȡb��b�a+�"Of�@$k��M"��gĘ<	!&E��"O���n�#@����ޕZ���b"O\ii$���-
h� �$��2�"O��Pn�' ���Ң�̇r���[p"O�K� ͪ>-`�Ӂx�p�q�"O
9�V'ǑJ��,P��Q�l����"O(�1�L��18hl�
�#q-,Y�"O ��gH�p��֢��[o:�sa"OJ��v$
.3;�1�GWdbe �"O`�sd��C2��׀�!p?�X��"Od%��h�'\tAQnL�<���q"Ot���K��Kl�t q-ƴe9�!Za"O���f�]f4���KJ�Y@�q�"O"X�KW��2$l@�M~}�"O���si�.Z݈r��E�u�E"O(�#g�	>�j�R,,`�p"O����&���j�5� �4"OH5y�a�$}���#d\�D"O^�X#N\<*�����n:i�"O�e��E�����q�MR�
mA"O�x+�d9O�t�yF�
#<M0�r�"Oj%
�Axw��9�U4$���%"O�$����?3�����]?B��թu"O6��T�2r\uX�AN�����"O6�RB��r���Y��._X�R�"O|���s� �;#�ǹN6�=��"O|��4��nʘ���J��n�Yi�"Oĭ�En˦	2��aꖕ k�Ր�"OX8���C!B<c�h�"��}�"Oj��$Ab &�!�'/��̒B"O��2��f�J���8p{a��"Oƈ��+:��{&�Q�g]bR�"O��S���n�e�@���R�"O8��@�.e��Pl������"O�<��)A=��1#���^P4]�"O���Ѭŉ\Z`Q c�(.]P=��"OT,y2�ƫ7`����*qI��Op�<9���+�I�V$_�v�J���p�<�$-�6yZ3��6N8�H��Fh�<ARiHC@a��:j,����og�<��K�8θq�ŵnh��E�a�<aB&
� .U�t
[��0�.�]�<����E�5�d,#j��c��ZW�<��*[6w xG �D�bѐ@%.D��� F�&�"	@�	�I�>�1D@+D������g8�P�"�	 ~!�B5D� �怼D߲$	Q#\�=4p)1�5D�x v��FϬuPq�F>W��Ѧ9D����!�4�����#�jXe�#8D�\ 4�T�FF�c\�����m2D�,J���-Fn����9�(�!��M1nBE0��Ƙ ��;F�^��!򄓝&�(����M|�I���D�5'�����*I�t�R�V�y� ��iM��sW�(5#�x�q��y�ͩ&b�U/Μ.\h�R��M�y��ݕ����q��<�zL` Y,�y�!�Zv�ڑ�8j�0�a����y
� ��c�T�9�FD�A }���x'"O����;� PHA%�&F��� �"O����������D�aw���0"O�X�q �*�e�!��'9�Ȱ"Ot��C	*:/$h�D^�<�pf"O4�pf�
d΅����\�j���"OЍ�&Mݹ� �B3]!n���bU"OZm�O�+�\98%
ĳ`�*@��"OL4�U��>�hKRo�Mؘ��"OU��ɠ,f���sh�#G��*t"O����K��bQ�m���(t<���"O��C�ԉ6t����T9�
|)�"O�S�ܨ~�ƔqGkM�2�~��t"OМ�A��-[��Y5�Ӊ;7��X7"Or���)܁ ,��:ዚ#U&�]�&"O�qi�a^�OPTL��	@�>g��`"Of\�E�B �ԓ�h�Z�4"O��)�S��ic猃I�J,��"O`;Ge,I��eF�|�ƌ��"OR�+3   �